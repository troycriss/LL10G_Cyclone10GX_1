`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
i1IVvOo14iSXthIkPRGOHklN2I0LPMCqyt3vIQ+3xNztTB1sLGNJ1JMWgGj8RQuU
LM6zH5AzPIO+4zXyYlUmt5nlT8s+lQ9VqbFik99hFsp3C0cWbXBI8C1DO9YuR+wl
V2OEtS7Yn5lt6xw3yiCqWv4bnkXaootqYmDSUYktQ2s=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 35376), data_block
i/9hE4F6/77tIgRGLMc94JcMTj1hJVsbg497/tX1YG4YwCP2XuTzjFW/+yIYQrkr
RCaRjrEW7VQkgMKlmFTlfl4vfP7iGnckBesmcLEpnc1gfhH5fEQ9ORANkm0SR1Rr
Et85eu+8hPOa0Dpibq/1Av8F7MPMM6nrm284fCNNakugm4jWY/uhcBh1TkZ5R1iP
IuJYqpgh2WtDhSJIfe8JHJr4D57QWZ7LCHhRCdr83XfPV5IEo6DMkVNH4ac137VU
6s1l9k5+9aYzQvLP5UOZ9YGaZnK1mUCGwSTNpX29YJWbQV07vN/xNWlL/xlrJZy3
/A/Q13F9CIsZOnsFmKPEs9PLU4yV3CC8mN88inH/ZBg9/8fpuNFgLgi5zsgdQWvM
6fefQvm+g2/6ezDUzj3bac52Zj7r+WypRammE3WqWLD+uKOycl2gRIQq9ysjh+ns
lWlHNNGyUhUQQnrB5G20O7Y9dLjVqbviZ6HFal9eQg7pPphDOQV/kAqdut8PQOpR
okHVRqS/g2i+Ij5X7HvbJZzt0nnVCNhvcZG3Bx0CdodVorWkowPCI1Aavp+NYN0K
JgWi8hHp1FI8n3jGI5GXoZ8TxYerJH1MXB7mrWY37DTkz9nbUy9LGWA7KJbhNxTJ
n8icuQS5dmRx77dxnHCTM8cx2H7Gaj+kKaY7DFcWHcLGLIAuTI6Od7JflFm9Y3Kv
I5/nOijX3kQKYV2Dw5sparrWMva7bngTqPZScA7/pRB3WOaufsRGaWSDYdbhbVnj
V9GZLhyZy/L7lRiPvIj4FCNF5YuZNxC0zWYMJMEI6jXy0Lyi6rvytkWwScVTMD+X
vZEge6oPxdHwSMopX1EJp+TmXFHKHBcwsjLQt8/BHOUWjlsr/U6GXHn8e6twnEDi
+XW4VVaexEvNPSgnQ9T+xhHH/WBSZkivNbyUE6Jn5aaHgoDcwgNsHc3oH//LdqAN
0ih+SCqb3HpR0tFl721/yOk4ydb4Q5nzfyC/42anADOBYW22+iUIHQG5gng2R90X
PAZccMCd2GWl7yP096kAXiXaybRn78Cz9HRp81Rv+OgVdZEg2ailT9JheoX2aVYJ
KsCKnoShERJPwJz8U8fYfNmOWJWlBka6y931S0pYrvqjOuyjKK0pQhiVLHpqAf1f
yW33eLpNP0irbjZuEEnkYeDYE+NXH7OX4O/iuvZduz0z8Ja/TEQijbJYzpdCFi5j
nrErK+FpAzrkIHRmk8HmAdl8tYSEZreFZlfCmmqBha5EVQDYOUlQ3y1HtglcbjzH
CAXq56shlAa0QzvDbrsSvqKd25kMMwsCL8jQ8Lz+tyQUmnvTtPgnaaS9dF8sH1U4
KAiYM3g7NaKOMSphpL3wmq8CeLu5+BjTUZNvmIOu/MuzG/hHIZx1o5xDrdZxYP1I
0ihIMkF0MvLaPQDKVMHK5uUB9lo/oM0B2BWdEsnAe0ssjR+KW8xJ6OJkpO+W33JW
iCV2MBImkf/QFpgrcbpJ/hGHzvVQ3sx6OvXfEaKq2caT2QtfZ3TZZiEaRKKfTszZ
cJc3DYbA6VbSUA0t6JLbNQ3mrS80Wyf2xlTP/CphE1cq7vbllIcq8g5NoF7NPEuy
Gm/6rQs5/ZzOh1dIqvqHuZpKzZ4C6Ywa58Md5xVE73yJowLiXiQ2ezIZt2vaRH+p
sBQmD8BMAYHrAsjf0On0I4nadJO/uW6BY+eQFBcAUhmFSB8oWL9JCx+Oszd9h1jN
eQ6gZLuROgfeS2X1q/PtxkYdh17acPWifBfu1zAMsWpg3+IrfYmmW3PgadJV5pOI
L9WOWw4SYAAkC7jm6mM7mmfU9fDGMR0jIHyOlMWScE8WKf/LNhRTwOghIC03dlTl
rbqNCxE0dKrtmFHRzV3kGQSmuqD+904zK1atu5btDS0KKKsFdq3ZeavfunS6Iw2+
tGeuxAvCrnWxl+ltKbzGcIuWI2jOHJPG1NAQtGNy83cQ3xQzftfjcbCpMaPJubdo
NPoYOiXJbOvIPKXzwe3TnCEYZxxoota1tFbVs2M7WbN6o8QFt2plqGrJg1zrJJfO
Xu1OmexHhQqWe9buMeCb++vjt2qV01M1w+iwAqUUsgqRulvv6Q1Wjawo7m/HsZhf
c5DEclvSPKSpFWQLlILz6QrzcSfHDnMjTg6JxCQ+W+66IDBsYJODYjpaOaFt3uPp
ziCQs71IQH5AbX3t8YzWjexO34cdgKM2Si+GPq5L4l8WTyENK+yztoHr5OrBzOLb
hTmGO9Mj8i0PN4qf3z9M2/PX7oUf22MkWcl3Rcrv0KkQjmXpWYV0rCIba0g0lZpc
A3HcM7Xijn6kVSniEQgOCY46EnFKpp2li8LJr+Wb0rrvwXtF56mxP0F7lzBjGqbQ
t+WTyRN6N1Br/MKAughBguissvWY9EF1z40vHTIDWdwXwZkSaJNPy+0EeJNqpQuL
+W/8jT0FGbOKbcgr6Cv9355FjUwH5F3ldBwf2GzrYErecvpui5LIDwVSzxIxPNqu
kR7d/Rfa/YbF46Kuc0S8L9Q3huv8vrj/LnB6r8Ckgd8F2WZiq2JAA9RV0rwt/6qy
qqTUbZHuggPx0dKt5ydVIEtP/sLqVemVLblc5tzsV3yfdDK1Fnm+kmtoEr7RUIIF
7YvI22yNjaOgPr+XqdXeVNQI1gDY/bPUoI/lwzItM+t2SdJ3+qby30ylQLoT+Lz8
r+9lqzrmGl47OLBWwShd5mqNyO7OVexbdgyezAQ56NxSvPY7z+Qyjwb0RUi/ZGLf
Mtt8iltxEWiEfEIk+TgPJNQz3MTQrkcDMmjCN0sVWfVOsuOjss2vGvulmK4FT/m8
Cd2C+ue8MK+zIAC8iUnXab71MfcVcSqI5YhQF/JbUdp2+RdWn1q2f50bFAXIUl0v
zCqWNFncwxInBTR2bPyDJ01A6IVyoBkvLRlbpGSKlQdPP6nfMCD2QAlvtdKu0Hnw
9/9vOUFxQY6y94+OeIBptb+7IU2xSXM9Lck6LDujCHr1VfZvLMudu29RzsVD3zP+
ZCMa4ZAUBdezaIqKhdtRADuWjHys/eXDZZjXSLBUBMPKi5wzGpMPfUDP8LA8mAxi
IKClTFptgqybjj8JvHT+s7ZVY7kiJOjrPGOSrzmiz1XXfsIvy2uHIRGIuIA2LBez
GMuxV0yJSLaxIjQknPZuefh4cvU8um+YX5vDYznr+zq/geH7kVNnOlFEccdHWnLl
q4KRmJPeuGm98blo3b8Hb79/fCLT9TOHPoqixsjmzsSs70r8bTk0ZcBW3c6Jxy8C
Y+EcI5mBo4UBsA52qt4ngoqiN3PgY2I7eDqDg62ZlwoMFox/N7jOHaWt1b3SNHX/
lEak+mZJJ2Xw91G/Xx2VmWB2YCC7kvcLe1H/QjWqV+XGYlu0w+FwnTyX1faHe/XE
pI8dne5Xrt90znQqQ7vQmaCXJn4tPNWqtzoc6tPLlRTsp7X0DlKdchdMtms7Wtfa
r0GGuOs2E3Q/v+DimVIxbN+vNE50cLT058rrO5uWLpQiRrtZXXlqn+tWXYgW/glY
0lbmsiQ5LKMhikNYWvDTdCHDCatEyNDmBZoUg5o00ati1LPgz+Z7v19fOISTbFbU
PLPa6dh8z7DP7xijTWDZBSk1ue/Sm0wA8C0BKCZxFXcoL4AeJ2Oco9z+QBFBDdi0
7CtayOEr8K7IO72Kcx/5v/9+5DHesvGrjX+kQGdS9xjicd+EFD62wzdQHTMacClr
qOYSXA86YP6ncv5bsTaZemicy3XR2d7O1mscLKZvU9f/fLOLihG7iYPv1whzUYHL
5xnJ4oDU+sHhyeHV9cPnyXFSdRTnO5DHP9qVL+YEXjCjA5q+FT+xQXfmF0IvU9Hw
kwE5SHrTIqjtc4y3O6chgasj/kp72rMeGWQANRSwLebjBKt0tgdAQds+QKD/AAWG
JmQSd5W2zRbH4MH/56wTeyYKzKDXpgstLGapFQkWnkBFOF3ceZ2XUu/ot21FulJ7
SCfSv5VkCY2EoHRi/MyJ2leGIm3+BhaugZwgUbBShlzzBG+TQeI9BhLgzaSFGQxv
VR9IgaGlihNgalgbVy6hxgVB+CQkTHwjDPEUYwVlNsv2c+A68Lomoa+/PIOpAkra
8JsLP9qd29rv8Jmc4RGEWWImpK2oJ93r5R0IrpzkEJwRw6r+hE97MQkqevQBQc0v
K2bMf4Lac+uysYK4UoJs6LCzCLrQkSPd3ZRenJmdgqbK4TGSDH9OxfwGgMdJn+ut
Xlh5mH0b/4qe10pj624ZlXRj5FFHLGGxgHGffD6Qi9OGWHXV37d2n/d5fU9E+s+E
Nl8GS+uBZQq6PHF6pDCbJz6NBfU/stD5OtSgr4S6Dxs/7+vBw28WOydqk5AaH9Tx
O/lQpnFBDZZUZda0Ae6oGyjxG5NX0egMdNrAo9GlyKXd1LZ0Fgt3pXrGxx8Zu5+T
mdthRKdmpkMOv3UslZccTZuumWmke07tx6Qql0CarnRzhKs77gaPqYXOdvAGffvF
0thjUbtPK41LG+0o4QzhfzRirzHfOht3fLcM62gE1eckAbMTaQXg9Tkr70DE8Ndd
Dge6fNtZ2wvbw3+YkGA/8TpLjMq0xyV5qLAGUlc01IAclJ1omKrHf/ihvKto0JjM
1LsDwamfnSeIOBAQuX8YJEYAoX4TPbao0DHpih/Lwm+HlUBgPAOgOfyHubHfCUvO
gg38wWIJl20TllKUVxzYwwSFFhzc2tmxqMH8HrY92bAFr+ckoBIs/5E/kfG49xW3
QslS4afzVSasbAaSXO4wKUfHVUyX/jutzxphGM9TYUVjtpK730loTPcQF1zZC6SK
sP+aGMlfP/4CRKV1pLO0LoD4CdOoFznWAf7VnRh2hhaPAm4EpdnrTU5wngnb1CtN
RYXg3+5yrxto0wYZNWOzNtgaY8vxJuC71tgjc2R9o00hG9SCyBsnkwyTzE0YzQn4
RNUoEti6W+GB92Nk1CRpjerYJB2sMUZZXpLcypRAptsUNqtny1tsKjwAJpyipBg+
3zIFJfRpZBOKNrgs4xU+JCc5pl5IWQG7F82eax8Q0EJaRv/yVGF8sDKByZOgHNMw
EFRRvzTv4eowJheIaT2LAmHYdZQrOwkb3xeuIMU+ewhhQ9qZnfjOj5IdXFnqGp/7
87CGCCniIX8g7j+WMSFIdJzl7uDYQuKlHD6YVt659vb1J6RQ0caHPaPsS4LZlVBq
9c8dFmHr1AK1D4O2d/12m7dfQLIy/0KgRsG57mf0s/93YHFu0LHFifwmFdqwjxJz
XjmM1+s3LezODnYm2w2qfE8BxXAZLU0/4MtF5DYsGXx9/gbJX0nS/HnOOy56jUC4
RlmR/FyeijhH+izJdfiEIPy5qyLSh5sunrfHVVWBpM6e1hro052e665UfW/jgisP
OOJihwbZRxmU4wbv7Dc4ic88r3S0ZrKeDuS5kbRDwJi6FSXDPYYhYRY/dYlxGRpP
Sh4dRr5/HBpjemeL5Fq4WrbH8k2WySDT+pkQh7aQlrlfhTYMY86qCJsC/c95flmH
paAGvtfbcdvhtCh78yBpcwBLY00Mqy9KIQFjPOhDjyYvo9Bu2mmeiXZXPT/I8Ti/
o52ZCrKD8t0dtCDkdfBU81qpDFejjvdN6LCOVk4aQ6KBBxqLUEW4Ki1u49CWOiOD
Nz7fjgCJJG8DHGh+beiNEHrzbH22LW9HmcfpJ5YhW/h3J0N5fk1NBJvC3WzZPycu
wReX8bZ9l0M6pctjP0Ul2l7xRLFiEFNYyt3x27tqDAfz20XmhLO2hPEULDuIwszV
r8VUB125dA9ZPAB2GjxlHFRE+9mBJdSb2QM8MViNrTF8r0n2e2zrYo9CEdD9FtIM
GfRUX5bXYz3rtXahchvU3YvrKAG+Ouvq06c3yrffsX2tJW+OCQaN8qx51lOvpKCm
wH89XIGAtLVQL23NjFVjXgYyIwSQad8f+ZOXDKSMZw3Kcp5dnrnrI26QywnWcnzS
vSYIKT2IOaPsyDkiw21K+vA7myxbPc6sN+31qpMub6ECdY/KUQSkHvJA9LYqk7QK
7Lh/FF6YGunRT+on8yVSFl4eZGAIWlxeU7bbg7lRytCo910gM6bgzIbCsmcMt+ny
yqlb0FyU2AluU6FMTNCgc7DdG8w9F7euUOhySestKFZuoAj+9SBAOj6L56zpfNua
QMVR7YXWEH8SJo37Y3K9S+miSeyxdUjVtoIxc3sIS5Q13hUVI5ZTjoHE4yf/OLp6
UMNwodFC3bIkmWRu3KHvy8SKXKcUbNZL0u0/i1roWHT/V0dNTvTftgBEO04q21vZ
sSAZatbc0B/4jFVijZ4gFh2G9IsXmdm6D6B3/Mc8STnN+StzFArtLFyv5vkRLMvW
2iS039r65U7/DWriGYxYeidrVdEg78WjwBoKVzMzc6oIWuTe8ltJfkP3KM9XsAVA
9wjlRXJWcI4POYSbKe/pd/3Td6bTOi5M8/YF9LiQmZ53Vneg+y+0y08ftrRPqfez
AlZyCyv+A3Z/LmbrocSqqxWWpzf05ZFiOoait/IMYirrgtRl+9js3pkeO5CgZXdj
seLE21QihSwNc8QWvm+tGAWadSZbTKWskH6fVZC1t8C4xRFqlvN3uoIBiE069dsm
LA6OK1rqmdQjTVTu2UFFfYCg3kNUaUPwDBKSwTHCEx1MjkbTL+YBrrQxNQk5Vix8
szb21W/00kmGCk2TAxEPLkWaQfOKOfnU/pOxzc2lK1bjXOcYxxYZF3Z7ipRjFx4E
BbpZjojIdMZXT+OdvV6EWPpzpxR+pz1dk9fMRsx2b+ft6FOLxF5G605mGyWfGggO
J50A/FG2htJtKktl/dgoWJxZ6BPr0OXAlTJyQ8F6xPtufWD3QclHMQOiG39iNTAI
MUgyah3WyYs3e9GZViaYBNl0TJXbDAtObCTngHjXDt7buqDLOGdP07xyhoMPUX8k
B8NVjsOEI+uDkFgFuIJM+9Je7aAjbeFaLThyr/gOlA3NP0mYyxGgxwJYBTjcxTkN
JuP3K0FbJ7VuejlWO34HF0dnRAszStvhgKffAJfzQr/eGg64TbH0TIdQmoKdBXQL
B34ptFpsSNJBHelTgmXQUZ/4Fs/wZqE0u7yC1EAVZRNOct4WCANERk2hGaoVx4OC
UMAJLtFP3CFBQW6Up3CJcDOj2pZ02dfkxNJuZtrGj+6s72E4N+v/9DX/ml1p97XX
wyNO8dvGe3GjEUK0Fro69zD91Fa7UAmDZgZBCGxiw3syfBwqEvowuvM3yMEve5kw
qVT3OffDbzpHL4GwaRgmjJ9cq14TOQnK6RF+BmMCLPSRIdY61ndW7gvQ4nRvQcw+
rLvuWzKAfeOHJ2ZW9azrxD1LfGHOU6uJNy2oL0ipWbWgUv+o0j/IUDxuteearsaq
Sz5nug7iY+81tEZQF9dW5FniGnHsEc05xP6EPsyEqXyYCtmyFA2TMRsg9O85317D
aIrKvoRKx2Ocv4YNQvlNAIMNOm9RNYYvLfNF6kYZnCK3Mgmm6W2FxiGOiCkRMhS4
cwCGMacA0KFVnhBRYrxHULNFuzNMUp1JQol6GKZ6aM9wER1RL9/IBcT26OpHWs6N
8tt8Cse8O2k0XdS7VmWtX1TEqtA+Erj5o/kFbdjxVDaIuFFbHoJ9fPqmp4iXcZSO
9Dnm9CfhyaW7Ai+Cm891mc0DF6U+Y5KeVKuR2qgtyIbITQfUgzRKRZiyXup7izlD
ef5GTWIaxfwH1y4Lu4lQuLERK6CKDtZikkJij+D4twe940GoVaqDW9WSd4d5tZ2j
6jwVAidXFIkNngAu4Kpj9Jqv7nILXbbAN2aV7xMqHpfTZSv8XGpVKmqpbVmSE9fQ
I4fzrbpftLzzzsitVKRe7gv587ouKSHzOFmLcA1hi0FARed1j37J+5i7E7Gfo5jg
bevdzbxNV929xPLtQnLaWoa2ahMGuBefptklwSzCcxVOQKagkC2q6+nG0DFvscko
HVZTYwU1HcVk8E5ciM7EjOBtwdazxta4d6wLqBr1kzKtWo0G6fSiaxOKRljSzm0q
WY4AC7k+itNjZrUseIm3Kl15oxEMnyiCVFE9cPJt3VtsCTpE5368y8oR7jtu5a2q
4x146n0Hz6kV5be6LZYa9RxBq5eC77O+tlNFtUnD+zbnXg56ZKv0vBdmdOspRyGn
rT5ysGkxEBZP/O6im+6idPervrtF898QluSZQxhrVbC4jxEBCaswK+xOAgAELeVW
ySZz86OXDOdCCkcDNAzFukFZcRBXlIYQVEsQTdcpfJZVm082knEYaN6uUI5fffE1
9qbbUV3ZdzfLz5l4sJqMV9N4N16lKYw8TSaLVW9AVrwybrKLReM1y3K5eYGmI1o7
KjtukyL4BV3UOr4SSh8w0PdCX5imC8ixVwee7yzxF5UfHRVcaqH9KqodZH7aXtgE
JyRcYMy93z3WBjm4l9aeCUdxwYzTiX0/T6/wDlfHkysZJ3AXklXa+zDPDriqnuP2
JYGR98yvs748oyGL3p8/eTuRihqlQgAt0K6qhHx3AGjaJEM6o2b6VVqKtvz4V6gA
c1t1/KEnIJ7O5cVS/P5Z8Q2M42wezJhiOLUIWiuSlJnhc5TV6WUbaUANCoU/jnfl
3Cn/6+Sg2Zme9JifmJl4DPBqI0XByiN0+S9ABokxhm+m/3e3S0bDaq1MkolJshJH
rqJPiaTlWZqRFkrkixeENUjkCWfA0rAr8JbqnQLor+QYlYkkpfwycyxjzvgLC9gZ
+ZAm7/9DElP3lKRynrF9LTLadxtJ5oYcSOtkMYegWNcDMaP/efnbK2k+5boIoDFy
hZLEFyGa+V5eXoy1xec8/eaESl3IP6cGTF8QVva3jDGeeSAplF/Zv1n6Tl0ZTlKS
Xc6AYneMEeU73tjZHftHTji6xDldXFBRdkn+aZIGoqtIsisJCBo3M5M+h5DHJgY0
VlIf0nInQISLzKDUZntjcEX4hy0G8XwoGJsvwEGQsBB/Fa64y59PjSEy9YCk45Sr
b69KCASwaNYmEx0eIGEz3XuB8CgiUXrj6cBefYFfQSqQKVbCCUFwYof/T+AJmHrd
vS4/MB/kTmgOqDSTofqlWd2F2GHCVmXjyQlL+MFbqSHoe+Vzs203uOc2IDU3LB1S
1DrQQXp2x/b8n2O/XWn3gaLY2iaXRrTD1rPA5qBpiBkAp+p8YpBZciFNYM9/n4Ue
aN2bbg+Ft8Hu/Io/Y9D8kfBENeYZEJ1lS4iZh+coQXOI8Up6CMTwDltK545adS90
hc9rOOAdDoZEA9mn3PsxzuGKt+csujp9eEKKhN/Y+ufFQ4/fskhDGYSs265SdZhr
rtXd8fOkQeuQ+lFzIEzsq5BBvOsz6fhWOPRsYOvde+8clVbqPhYyUBjoJoL9hI0W
ILIvVhfb72USqpeiTNOuTweseoK7lvduOvrWIgBh+sfVM+zSWs4/7KCx37sSFqcH
3yBSCh89mzYrkaJ78c5sQ3b5Vikeb43N0V2Tv2/+mp/4ieteRZlY0b6dq1+09Mjk
GF8z4BHvIV71wE+ohCRUDhZLDalPMIycpfISmklfpTLkIFhCe6YrGrjXOxvKntC8
gvGCvYQH5OxKyMkFprgiIcZjMeed0Ry+Krw3jZ6hAsmlBZfiM+aBfOfXvN6Du0W1
Cna0q3tIazAbRxcBIcdGXqsvPf16lbzBgo3IjGb1U7nosqMPozXYJw8IAV/DJGuJ
5b4kFiJxCdgsA+z4svaz1zirDETV8qNnXU2pA/KdtYROYJejWIkfPFBpQBEx/W/v
Jmy5HiHTcvl0atMGFXzDge57rLgtBDFvwYgmsnH9hQT5UhTcSDiD0k3BufhkW2lu
A8pd5BmySuPh5Eze2qKqFsNE+YpNpbrJxgVC8y6zc/lW7du8gMIm/XLMPIO9DfK1
4vjBrpNO6IVYx23NlYP8TkOYPcSl1J9jL+g/N62SFu4uaU+bSOrPD/znlbQcAhYJ
qzdwoFLMeTAR4kl/P51/Mqg63Cg8WvZ3gzw3UkAbiHRc0sL0ISgUondTXLbP4lYs
64b3FamaODDP5bhrXLQLbqgibRqEJrIFisGU1vmV/WQq0HHLsoCynay1k/kG3ghl
ih2WX3DXQz4qD9oZeTPHtP28oxF596od8bgT6iWQMAXS3VDeYgsuhEGR4gm6Gh5z
+8Z1A2jhTN7zs2RjmUKWYH4nFM50e4/oKEeKnlr8xnHB7PKaELFGgWjPZciiRb/2
p7Nbo64XrOU9oO8lrDSzFMgCQCAv8iAQVIB3D9gdSe31R00KJmU8tecaJD7aNFJO
4VSbf9u6KohSR31/fClrcqFHIO1BKO83xEsuyORqIm72URE4Gh6AJed0MuEbOBIl
4lUNdF0CUFH6z3ZiNcu3aIp9g7CvgiDmJGb25AKtGm5eqmKMIGh/MrQPhgal5CHB
lVmKqsBXQvdwdDthiNmQ7UfMsYqKToo1evFZ1/xKx0mQ+kqll5KB9VGYa9sG3rFh
BorErkwgaHemalg0vn9YesEaRj3lJRG+QrKGTChVl5YRu2EBtqfE/WejKviZuzQD
lwkrWF4La/8DyGBPRkcHFPFirrc/0+IRuqbogL1l2NLOTXlQAoV2fVSg8ZwTBFv7
NN5DS+TYpWngIXniCCTfBGCJD1gKx6Qn6u1+iRQRWmaOfbtPvPN9ATDNRs0+IbI+
CnALU3UQY+x2Z3T70N+J5cSkpK7Z0gkJE5ACsui2QZv3hYEoGs0+xJ6xokoWI9ej
a4NXnKGeqTpIrzHHcYKYtwN6K6IVsT1nPG9gul/MTcA7yYl+tFgNCNuklXcsnTKA
A/Ry5hh178ICWY4N8It9kS9lFGl8+a9D+EIMUmx7L48Jg9VXzPg0kH9wzmekIpl9
tY+sI8FPYcX1USjvehzWsuNlbkuzorK9CprLCRPylFNwBpbA5rn8zaR+wLbvLRdo
R/FYZ/Iq6Ov141q6x/pWK2lK+qFLuURojG25U8LOah8VjF4jsP/qIxHQoSajeruC
nWrck5uHW6qQIhDijKHrLW4JSuX9z0mOHn8KbYK7KGUtlISrZJ7m3e51L8iVC09W
Q1aTaqw1GUQ2JdoJunAP5eER2RjctRM9lRol9+SPIpCDn/2FpuZ8sYFj6ATceRTu
7GueO1F6372ABHJKJjNdyRCKjalYP8AUZzm9muHK7sog73TF2toFxKq/uxosYRqJ
yD7fi/YPCJzXJvn3AtFoRbngU5M/VBESFKEo26m+j9EXM9tqRYDI/IoYK+L/fRXI
w6QhGt1piLnYRMHGcren0ITOkz0jOdYEdpBLYKG8VrA9r4hWlx7cW5SIP9NKOjbO
iHjfOyLfBsvXyAI7fJEpsm7LMz3KC8FD3uZ2EUZSyykjCxVG1fRFblYXVd7pf/ro
Ys/cBT/QaFHNePmKqKHT8y32S8IoEMq1ToYjBdfDqBqVKZZ32622XGmhw8kzPnlK
VP/n0ZorusvekMry6QpmwrBZVh9hOmWgMQuPhLY4Ec0CYmirsR6ikpKJ+FwtmPCT
87WBNBa7ISCgWEb+2pL3HAd+n1c6VXVAIiI9sLC4H8FjID0pvIqfUB1iYIajgjfc
I7UBMygnnWpeeq8ccKTspAJY6c0Ly/KS9pcv0J+63B0mG4d+bViGmbwWt64zHvKu
wWPq/ran9mGDUtMtibf2q4RcnRjoIB3xIVIegxL0dSxcQiJhuDkyd91FwOdWleqJ
VXse83+SAW1STX5ZJZsRF/teJxe4IbpjajnWsyEmIo4JZ/Ohof9PxsdWrp0Rt2RM
aVR6gxPb1V9HsslLYJlPQpJg6+VfuqXCsZw0kNPIrcSzFEyyu1fX/CJK7uCEtWjT
9CrtckeuV/Bgkf/McCZbkUTC7V5CGn/R3eBM0QFykxoKYLgFld1MvYbDO9fgEdRa
YfzoqIb7n1CpKrAWvhZ5a01gtEGJxAuNbERlsS1HhKVs87QryGSR9+8z7tBzUyRN
YiylaqimYtXxTRzWQMyIJ8emwRftvQKJDOzyMX4vVkkDQEirqWWgXmAPYGCwkfKs
6B/EbcWDS6g3IhYhi+JIQlvO20fdGYRRUrDPoLcu2G4xb3Wju9V8rHaF51Ixa/HV
J6a1u7Y0aclpvAiojzCu/uqizieptXbiVqMYZUWe3XrznWON0MhP6uiubostpdeo
ep3qrP0FKCbEha3FpWfCsC3CVeCIpkR/MHmroSZx2C7FIRKvZ92LQszRu1ARYpVe
YWweeOzaatJ9WepjUNmA8msWDFY4F7OcxU34RG7wzIO9MfT9RFOM/0lsdfUcBKMH
45E5AmQ3hemo4WnUAEhjBaTi4L8xhEw+faj/gf1+kt5cqF7Y2SRPo5z5wlxSfm9j
R3IDpKK/FnnRmZEi5exCwV/SPzr+kXeAKYsFZu5CL7vHUMwkXi74EWnUgyLkHdnI
y7RwgmCApBgcxJNH7LDXFsqLTpo4TxWCLGbzR1nHTZMiCc631uZ09gZ1Sy7YWCLl
3KXPC/+qzbQpGVsXXHwlI7Y2GYzf2d0mCWmYPQZ3Qq8WXiyl4p+EYyFGqyxX7mGb
sWaZoG4ZWsKciT5sEsLH9cpqfVKJ/fWLrkkeA34mceQKJt494p0hzi+zZzqCUCNE
alsC+C9PDombaj7LwqgjImteIlhm3+DmUkja9W53grZ/pUAj7tT4BcI1S/uxqRJD
Rq3tSq1iTMADEiDp4p/heBdC8bEpHNZ7vQ96qrsIzOYDwNiryb0XEutPCNDnjS5X
Mm5HMrkRvrCZnNKKNtcw1ct34LcKSBOUHDDHBow4fI+5dIhK35DFM5DRWUg9iDSj
c9XTyNi+GCpollmTHXZv7BD/pmE9T7mkXaLzd0k3dP9LQeDx7B1BqXqiQnQUPPkU
ch1wmd1NEn2j4n0c7PNeT0pGoQ4eAt45V9naZjAcxJa5ibGA7agB4JKIEEE7Tg2B
8NCnl0AI42av58XHbLShaVO1HZ7cnLv3O1ZD8i4LsoCac/111PyRjqTfeeIXvglG
YgWszt6ty34+w+3i4i0NkkRoncJaFjOMnKZRrekYo5YiVGGiOFF3Y8C+8LT/5rgw
KUQ6TmUF6za8Xc2rlTI5vBPntq3ShuhkRSXSmtXtkzvmRFptrVcNbtEklmEphWJ+
vYsIEpArmf2zqlk5XT5T7JMAWIYY+MaYgzK8FY3U4ybb9SApaiq8D7fxgnETTq0H
FBgVVus0W2iSqmGTJAcIjVxaCJ0lcXK+jHqReBZL4bj4q4B4fAmQ2fAW7oqEHDnq
/b8FVCjTAN7xGLtIrUajzYKz76XrGJhzUj2mohXTjTyp5fM68w5GMZDaegpnzbRq
rJyHqjRFQoR9JN/BvD6lPKiq0+6t5Py/Xio6bYW6MXMBqdeD/rYH9UZQ/zRxc72J
s6DH6bJVsUQQVg6KrUND67x4FIfCf9im+CaVb6OWXPb+L8vLtZtNg4Z9yCeo0/CP
jPBY4pQeCxT1IptKgMWsekW6xKYeYnt67M93XgJAO2z3PnQeXzCUz7Ky0jJArHhs
V2JjRQ0xJBkbmOMVEdyhpCdbPBeXDC+eSLn4NkWv10q9v5TWOf4JrVhwURlaTcyH
/EIWvSe20XLPJAPMFDAOQwTrAYHwGS2vk36VP+E3UMzDidiqdMM6lJ4ue97Eecsn
HnnUyelChEWSypx/LMh413+m3lCZ9iB0ISS/mudNGoepZ+Wmz0L5gBvOoSyGbYHv
38rhc0DP4A6FGpV4TUGtoHqHZiwiHuAj5QtnOyyJBtI6Gb4vuBE4PE0rAyb1fN8F
GYPIgvTdZ0OZJ3LZr1qJfo4oMowlbuJQPgWtg6a66DOdz3JrTEiodZ3TWQusg/47
aBN0k+j5/SCtcvzchg9gbJUFGwO+rlTdIrtU8xr2R0xyHKUTyUt/iS3GWST9+bCG
dTeL0j3eogHdjm1vHQYySeSIdLZJ5OHCLqKkJ0GBQAF0cmaCni3UATEyXFPENuBD
XywrueXSA6f9zEQjhNj0ay4se6rO5JaONVmlTVxLdI/Ratc3E6nOiAWJgy7dshXm
RQSgmRO0AROSq9Fm7PDWcIVYZw+yP0Eq+ytaaM3F3sZw8d9dm27+ThgfcfreZJCx
pJGpK4wgbwhRi36+Tpy9Q5y2YuYL6etssFXUwlIAcv8twUIYlFOg+CYyAP4fK78u
BWfNA9r38ek2K28SWjD2/9fgdPHnqpRiyVcjXQCbzB5W8bSazQ8qGeMHgBgCFY0j
jjj8vKuY1qnNOlyJVYl/NEqUgZ9Ikh3OGDbNdBfTiZ54S9QIO7qVwEMEhxGnD5Aa
GPJm6Lu4TDdLQyOh6ZgD5YjYizUkmEmSAHbweA/FeXujrK0IoUr2n5VOijYPUJpK
j8kuBlvrpv7dBcgM5tdt4gCTBtoYz07jqVdGbg9TPHECK0soZbsDg3CWzH0M3be4
Kql3JHYPElZdgbhoTd7Dx+RAlcc4gYy1MHi719q6If3d0Yhyu6JTpoLQEs6H0ZpQ
lyE9I8wRG/2bL38iWC6AytKX1RKk1yjIpqs5AX5IG7MVEYQlZuEnSmxZLbSQT0XR
/xCxrocz/53Vb6J1kp4GvU91slZMbZtnjlFcBeyzZVn5SR46vVyIrtlAo4W/cwip
YA66w+aiTmQxIVHpF3uuNYoehwYJCaZe1B5fpmxGdyx3OjMf6Wp+6BQfjykXb9E3
fc13znbCt7p5fJxI6Kv1eHLqf62bMvlTeCR6LgDWFnMV0Vj+4dMGbPS3jM/UgLJ9
1045n6XwpeVnpmM0GHshU+shrKf7DR9OcsR6B6WGENApu+QlQMv3RAj88l/9JxyF
0WAPT1cXn7l6LW4M3T7HUr5LetEggnWQ6zcYZ6yauZAOU9UhBgWfdAr+oWNjgkpU
uqPD4h2qpDR4lbKLOhOCKhnd3DsbUipsymC8DOl/n8NZy6upBwS0JsDHg2AKg3E7
7sdxvgPS12ceOMZli8EHV9PHrvj1yZdKnIvA1H9ZW3eFInTJ8pqXusFpDFt2MCXc
fTfMVobSarpnCM1nOw1H8zMEPQmxDgmdRgOtVytk2mtweib/Qf9cg5UFqYSPHt6N
Ae/jyflQ5Dt27Q6/uU/HgNAR8R/LhPIPvrYI/DTsXqonUUT+5uOwvanwxuCA11gh
+ZwTBvbpiuPv36wYfBjWmJHqidAOQaR5PXmwYrVHlz9QsboIb4Pnx1uc7ObseOfc
EwiEH0EUywnHwvNcjbnmqN81s7m3V857Hz1NBmbpuEy8Vfs4xFBzgYlA+14ufNFc
sTzdRWXzJJFvU14KAE9FJRcloRts4Zm2V166r2SN2QitzwJKdAV5JjI5IchwgFEZ
LYbBB6jzXhPwbnoXDuHsHQI1SGojBBH3Szh6OXpvC1oxhk8jY7aywkKt6nrTVNW9
OEmdaecuvZt/fIfEmoYMgi+M4o/O8UpakqXCCEBd5SmGn5NHOGwBD1Yu4pOoolGO
T//JCmwOE2IArQCWQxJOzwPwd+Uhtvjmf89rRCiYB93qRVY/x0vPREDiA7Giw6Ht
OlRHwu/H/qkixpIg6TMweHwcLzBztwZZ+s4GgHeh2GDx2mPVN+0KXw55danmuO/Y
6EQ3t3Dulvph/kO/c57QlzZs58/Mu/ZlS4Cp7HOpTCdC9OUVJE2BCw/lRf/Sv3GT
N7LWg/HQJFoi3KeXd129A8q+jcXuvPaTP6vxCHRTaviqbkqe4jTUVa3HuzV4ImW/
E1NjzFYpNsw0pxlUXYGlemAuHCJkklFe1PvbkW72NTVkCAJTbtdaKHkF0WpOR5PU
FhrtYw9oJEi67s9C7zwbD2w2zVzcjzh487BxsLbCD02ht6ltCmNUPSB6QnZI4gji
DRXQ6/aRLgEhabHqEaR17wSm0AOkih/J2vS13xdX1nOsMRc46X5dpf10pRAR4sEF
CD8v7OStubZG9D6YMhyV8oFIHCJrgciQgATRuMGqJqjEQyib+AB8Oz/05/u1PTcw
DDUqmV88lR1dK2Crf8Hvbb5N9jAZl1CVxYFhMjAIMu4vfasR1iZOK/lysM1YRTGW
P9m1zmn4gWKid4lEpabRRgLpj044A2SyYUA59rFPdY7MZRVIwxkKiwGrhQJYZGNA
Btrw0CMbfPFnM2ERT6CqXZAZDSqrDhoYX3ry6rQ+qy0f4LaRKmHYxOUpOVImbfGU
K5ydwlnuG3tSldYwNU++7NUjuq6JBfJu0nPLLkL/iU9qUisj/LXup9Vbbznzcb71
qHqU8YFvejtTAr0Qh90RLgjvm0ovlkhlYvJU/KtSuXuH/+/UqdXSV317Sh/xosTL
8DPtjXqQq7ipD/tJRoIR+JlnTfSV6Gmyz68r5DAgD/BsOoMtFRWH8VltsTzTOcDq
cNCF+CxLLb/MT5/6GlF0mag7g+zZ14WEpkwKp1yR0zaMCwi7t7hC0cvLchgQt9WN
JIhhe/Slppq28+uIqjb3meTIX6v6I6pS28AJieCY+UBI5NBDZsFN8R2FlqYoVTHM
qkGQvayw3uxshGu7yLEILvvQ5pMyUtcddH3e/c76JNIbHqum7dRj6r2LUsbrA9RK
/UD5/oFnBndeHFJwKu88Rm5IvxqW4pOjyhREkp48kSn9eCdS4+yPKez4NHJ9NEl2
X9SIiZuKVxQOTXQPsbS6j28Zj2jV3jYCBDin/2ClEzsm2G0mr7bl86ufJIAZ5wmK
etUee9LBtAaZdFOXmetfUJLFTPqlJbpdyhB9/R5seNMIM45br67X87X9b/tGjQoD
2qISd3bR1ObMN48RTexaAKvLyc5Xwcuy9Z0d3tAjY3YZy/ZcsI1TlYeUE9lzVdTU
YPRVBlrTDXgyOm86wNltU1Nk+HSMQsqsz09IwW6YNKlGbhbeO04RWgfIHFZlZrRp
zKyG9swjAP608zTD9sXo9Z1PMGohs1WIHUSdt04DtlI5z3dUMn/5+5xLn5r2xspb
TyKCFvPtM2JPl1LuAMrcH28xIr9Q/nLB7+++U4uYX3gHhHR24/GhU1Psjj94gunr
wdiqqHi8kAnvo4sQYAGHNtXAF+Q6yVSz/VKizL0lMFtxBy7aYgCdRF5S7t296qmq
JgLK/hvPU2c+qTb6Wd0Ngq7hfywmNpHyC6oNybPnaaeSJh+AFZmyPnrBMhKVhEo5
UMhHwTrMKB3ix9dNpPoMhe8LlOO3cmzC1cjDIdBq0SW3Y7iHyzi8yKo/F5mD2Vlx
tW1fnRa2Z6ERdOyOvV4rq98sNDt8ZiL2b0+pD8TpsDbf+hS+Se+bPoqBCsQC2/TX
UOB1QCxrJziANQ1Q7AP8Q3kG4wTYq+ua8BNYPBaxNdNPx08x94xiT1u0Qz/crnvn
rF683zyNS88nal3YLVPtMmWbrsbh9nv0fycTzES6TZ+VwIn4LPbHgqIq4yp5KruT
4Frojn8JJyOcKDg+daE393AjBd4lBZxXroko4cPVwCl4dVBByUN9dCPu+iIssoR+
AarQChLKUmtepPYbtE5jA93RbKUM5liFDj6Z4kDavdtEVcTF5l3dBb6AN125Debk
RqwX9ZVlBw2FfOZfgdSivIRNjrMDWWMOf17tW9Eg9dsRu6KqDRTs3SyiSmDpXcS1
rwMeVSsTOHP7rdvQMEltBMLzvddyzEFrGkAkEgZgPRecYqktP796+u7U9alfTYV0
QGfpwinxm4x1Sg8CEPUHnNKP2PNzoI/o7EB5X0kJmFyBQ1PjaU9aCtSsoSagy3HT
djFtxmGuSsJAs31cmB5o/9txy/5CJV7yF8f3V06EksqvLnn4H6FBIi+rZQFcN5s0
0jVjRRXiU+gncrUgLSvcatNStzJkBEaayV9T1MCACGFTDVI+OzJCmMDVD/L87KTY
YL/Vp9F2lNvQ1Fn/78Rwco7faWyiXAWkYI0JFiSZCEO2SDgxVIDzlQd4DxJBVxt2
cKm1E5HOmpjsgd6IPejl8h2D1t7jKyf8L3PW3FjafUXdwmYtDOyne8z8nBEjTQMi
k6DCMuEh2OLbCPbIG4dTFEgHIJWQgPLogejLyVOd+l4yeX7hsORTKLP2LwZaV3WO
KS/HAMBLpQVAk+pvejvjTYgvVKAG6OBFEWMigsLjzWLtsEbNX9KvOyikep5kyqz9
ald8Zg7jbvEJHgNRD73GauFNFSj5J6vv2QIwU35cVl0qqUW7MpMbQ5XaOuXeBFfn
TIZMmm4c7BI/m6xRDhkbuT4mhYKznYvtawcRApiTXUy9AsWoQtCIRx2tmGezkCvh
uQ4EASAOLQouwL8GCRmHrmU6JDFTswfkS4eF6z6LjZgrxEO00882s6jhqRuDNGuc
/MGNlnxdswOduAdM3m5sGxkU2JjBcxGVIXu0rlhH29PQL4sCf9fQVYT1CCkQXtrz
fjlD9P842nZ+8qxeR/OVtcw1ueW7M0S05q3MjpS+UtMooLop504DwHb1wwUbQREC
s7BD0DqIAHlH0XAqR5rhChXNH+zCuDU+ZXbb76Kzq2d0349Sd49k/q0os/fm3jjj
VD7ou4DlLf/wv0OxNVUPe1/FNLq+c65xigtzwbBuKHe4umb9WWh/8b/+dMtZ7w0/
OxlljU3K6+r7nyG2tgEwBEgxvPrgnLnnYL4DsoMyaNiiNqyZiBZDCP0lRcerpp1s
BAeWu1S8x+SuuN8oOjHunWmdEj3weor6JxBuNGWFGaRpUcpR5Qu89gMXwb7dwR1E
YWBPmYSMbwnBGWEE3I2M5KkTgtbXP8bchBb2ajlffnd1IG4YHGoAQaj+YRWB+5JC
/wc8/l4ojQwUD95fkkvwDViIC1T9sudcBX5fi6IkmKedwZAC/vElREfCNoBWHhjp
8mwcWAJ9+QtPu5xIFmmfszBaHT/EqO1+M4Be+XMAjFAopgz1Ioz4EABkozAn7R/S
mtMS/83wknKbL38NykHxkciA1CvnVDxmYX+G0zpCoiCddebGLsGHSiaNIkq3UCew
F5dh0vLrqxsmthc+GsBAj7ITwUH03nKiSDtu8KlmWVdI7w592N9s0xhgRUJu+kqj
5+0UaEgUN15oEAYdCY1XmMeOU7TUEeMKy1+IUDhAdm8ysJyAjC6yBea+SlrWh294
/BshzHGK5bbGSLKhsYXncVvZ84g9ahhhdHgAi/dsWNuj6K9bmSj8ZEgjBINi9/Xn
iz6zqZRjHQmnHYPW+OBOFUfP2lVGEInksrZc9NQtM4CIBwP/r2EWYptGYOWNc80E
rx6HNisRd4LcKGbkVvNhQQhLtqBD125NlJ0rQCboKYZLKwCf1qv4cdR9bycPKpN3
Tv6KKnUmSUrQeueecsOwzQW7BOOxeO0+oZEWsryl3Sm0Xk1ut9MvMzHvax/0j7I9
ONnhAXNGfUMGfbreVfGt0/fiNk7BukEDqZ+YwfhjxabszoihLHhOgJQuzAersOqQ
dRZAqSE410jzBPC3VszfHuHdj6+DuuiK0/EZ1d5agmSp24J7MDxL2jMcDW0pIZ1a
6MLGcZh5sWzJGFOwD1S4AZjN3f65eBWqZRU98ZrYg5tSd/61v1hHJdF5eFr2LCIf
hVvwv2M59F7wHIwxqzpOmSoKWKc5T08IIK9zrbqN5bkQQiFfRKMtFcpUv96jxJ0E
idaRlcTPgVOhH784P4hLb2BZAY5lMwUz0GP/iUgMGcY+QqJWnARe3YlO7Uc5zTDM
3pl2ljGt+2V7y3aN+ssWIMLGg0ce188ThulX7z3jSuZYXcoI8tA6D5OwHlQ6/tLT
D2IzZK9KXM1JPN+0bML5UbZAofMMFYrnz1EtP3QjKoC1wIb726zc6W6d6bcO0r47
rhZG3rLOBrpefkXIvtpO5lB25Vo3A2cdL9xLxyz2txnbtl7Az8XbDkJXGvhHQnkB
9kPqSlBgeSLdvwqhHUxRGLPW5UJfCuvimCjMUyNyYqgPO0CqRc6z20VgSZ6hXxrb
3e8JHvA2raT0FIB71dPhWGu8m9goo2IraY1duE12bblRbZiQLg/ddefVHbg8h/W3
BEm7Nont7bVUQTsYFPGqgZ7aiv1DyHD6+sfZHASTBkTjlgmS+2eQSTuLYIc2vPBB
uV7MnzWVphtNQSuFCmdkQ9a5l9e0ZUB1XX/JwOpOE/RRLjC1Ia7b6JoGSHbW34aY
gBPF/2t5Nbtx9IYRGmqw8maF4mBHi3zdAVfkldlO7WVsBWqu65oiMoifImL20C6I
qq8bCsWATuAU46kQTtD/5XAlIBcTJo/Zbjjp92XReYONi5C3A/lL5QpsvqHAMo+i
w0T2BFwn8AYZk9ROX2WS9/XI9Gh1GvA5tZLZ7WF6X4mSqKNvN4lreorSHfqKj/Xr
yaqxY87EJWMqOJvZ17DUbrI0KVGjntIwqGM0adWnDYNuVlf6ZnhH2ducRB4MiOyY
8OwkIdThd6G/aDXFFGSFxDlK2m+tt9Cleczu5KPN7QArbju4TrhkcrALfWtS9f0F
buQNaJqMJeJffIO//D5q/laSDilono67RRnEkMvUJxW2Fj2EU1qOgaxt/VgTh6yr
z1+Ai6xx2/iKUjYYaO16Eh8dKtZ2nQDjaprtJ35cPPYp7zNH04oEt5X5+RlQgF1i
0Vi21v7sOeMmMSH+3GXzGz5ISGt8XH+es5if6LfpBctzi6pHyCQag5s4cbRQuaPg
EncyzhaQpcUYsJJvjPeOn8CnurJV7oZBt4SxcK5u9uOWNppsews2BZDyWhlc7y41
EgTt4N9iftgT6o8obf4kEKMAyJ6qdHt4kdPgRC880ZIEBRGEakLjVEfo/sIT28AG
cD+sVD2N4V2Vhf+EJWyUyAs/yyllsUw+W52XPjFrJjPbfIUWpZunflpM2ZQH0T14
n3SsPMBxTe79+M/TDWdZOMEf0C42Js4PV1Z0UAbLXHPeP2DnKqOGymSNXwofQfZU
y6qO5Ks8cpyGxRQ4bYXr4waAvkgU8EGxOHjuTayavSAPhLgEjFMz+Q2twgKRSuUr
+be4alZcFzS6gogbNpfzi+wK4OnAGjrK3i05Ytu0y0QRY2nk51EG4rSpPD6arbrv
IcFAsum57DNNl8r9Um4I2AIr586muxSshO1BH7HIsiPi5Ldjwe4ZUwiw+uNVTShm
whDKyPK8Qng3gU20a16ehNJYvCdVEtxxnIFnI5NiAmVvAWOReRMoAWgAOTAHBvmh
tYvF7jQPUQuD9KFtRxwD8Wclg95K+Q3HbBs3Yze+cZ2HVnsyt8/NhDAitrZKFnaw
fvzwz735uVhs1aJ5Ch5CswCXOMq0J0H6+3G0e9Ph84ak8aChq8bMeFhkgjyGrwYq
jbq9pB9jFq24KnizEZYmQgDSUF2Yknek/IbvlxMrKNP1oBdO1yZztXtmo1M8y7jn
h50gwOVohkru16EdlNCAGZ5EjX/oflMnESbz+VWZxeklG8tFWeRqed/3hSwlTbX8
qGmFo3O8B5IJOlVPqAOrJuJpiyVsDGdOiFXE+O1trgNelaMRuoX5TrOIwsLhxF9m
7CPXYsAIJZ6SPNluDZ9AZur7lI+07/OovRTdZJblTjjNUmFMNK/1/mHf9e8n9yG6
aUIHUaFwyqN1cIkOGBaljRD9jwMvM0riQwwHK3+tnh4eTwqbHp8lZUOsFfg5g9Pn
dIILSdtcHx/7n+60uCRX3oe6HByZbOmTyH95CYlW/vEvrgiuh7ioJYTsWAb9zhii
jNCVIkFgSSzQ6ZfWWR8pYfiyFkrY12urW9v/DZFkmGs/qSp8Vy7pMP1DKG9kR+GZ
+JHKCypHv89lDugKl3GOuijscstgfPNvdM9v7F/UAryY+rju4NU1U2orVlCvkY3j
M3l9nt1cUK62cctBNQ1hx0mtkiGkOFw692ayylrvKjIJq4vtqLE0N7nGtZvpLvsw
QgZg5ZtVp5OgW7ix6It8ZzoL12e5+PXnbeGhHq3EZHH6NVHfErjfy3GtHKHw/qm0
4wx1IExxfr2tpy3dX7CFDH8Uih+8hmiUPfkNFB+ZZ8Lsv7iRqjdfbAy8/LYt42oz
KtGNZhoAnEvggT0fJ0F/cnpPmeOEP5UZmBqAnurnQy2+Uel5aoeyCYSiXdqOYHKq
4mmi5VDCsb4IHrqjwPBOc+gdmBnOVhTDmkI9lhmdLnx+GpMfP9KhUpICVCkia9y/
H6LP5cI8do4QrPDovxizyFe+KMpL8xONh4Rd4Uha9WNJSxKQvjyTDkS2rU4iv99F
eNRvOZvVTM2wIhPS7Ozfg5BkiXPQ3L8+L/vhwYrUBNbR+p1w+NFS5r+kZD7zmDtz
IhZE7/8DBKy6X5u3Y0Wo7EPldsUE2QC27PQgQCYpEpT6qiyJd2asd6qdwh7HvEx/
mBGgjIIfcd0WlOhomWnmTENF7GEiG1TpK4rqvu2nZfSVbsf1/L8A7VN82+Jur8JP
KXqnEvMDEpLaksuSncDbwM7csJWLoocpa8BRGZZLdcKt2uNREnNg2XfBlwVOWBA/
ioIZlrnjG/jzLvPeyU7heuLfCQWPK/FKsUewzFM9PZ78EwGrJJEXSUbs2rfZogry
qeNdcedYAqAO/5CgZR/GoYNZI0xFyK+2cfubNuHR8rXhFiBJqsYFFyTCe+ab+Eal
dV0lCR39jeL6LjpwsFh8Ydjv7PNMN7FPbNldW0bgJE3m2YloqvnthYcANIs5TGY6
jzVSQfuP5NBUyqhG6DoFTDIeGGXAXAbg3DXcUTGx94NHXLeW3rErB/nzzLBVXjV/
kh/8trt1XCvrfREX4t6wAEAqgCSyA3weinqS8l99gImwIHFGYTsv+1AVgFrQvjfc
HjfQIHKrizBak1QW1PmPeutBpzvNC3MnyxCP9lKmqNUbwP7gPNl7zLJpPRgAqayX
hFuXaO8GfG7psrIUlSj04hH4fO4Y9F02SonPEQYLOM3VxdMwvdUMLeqanvHC1U9L
43GBU+LEJxwrDB7gXBK2Edkp5QTNvxFlroPaXxliUMP+DAbPDKm/dX7jo5AIeQ9f
YQhMvBJElePdYi7jJuomWnRSpsvknSe0xF0Cztryn1AQ3Us+UGoO+LshHWJ3QYXk
lQw6zVQqELIof3Pia9JH4ZsjIsPL1U8bZSUr4a9DUDt0eMQ/HbR3eEORodGnCTRm
KYe7eEZvzj9ew69MMWrUGJ6E0H8h0SCsU0qWsVytSQG/DkVHVEiGCQ59IDCkyEls
3suEDtxM31HRWHkHpkzD7sgWKpMgnJ/guTgVYEOno+nJbBeHSo+27uD3W0cI9dFY
jeXXAn2N+qnghjyPQzqFPRySn/jE0yu68jwqOTWs30YIDBL0dZe7mOryx2qnQWrA
ZoWkhK7y50Qlad3r7vBVrjzijqGJ11BNZ7RMmeDzHTobdx0c2pKH/+un3Nn8bUS7
ATjycRh3uGEz8xiBQ/Pja1Ntb9P0QfL4RBPChBtRCsz/YDRqCdAfgdfYDwFtncVd
dxZl1SSM/ibbW0fIyakgsHJAsEGMNFZoz/uDQCYrRYzq5TZqEzXMEyEz+IW4zAH/
hR7vWC0flUaaf2zk/pDbiMBplsHZAb7+vVy6OLZCXB+Ws8lefjJeTHjBOF65PHmP
eEuZQQnUBAWQOOiBp7tNoWsGKtPMCZhA2SOGJ3T05+X+VGcD+09lhYSZaMar3zB0
/fDWM6wmNYgcBw6QBwhz+zJM46TdfcsGQOnrLZ+D1vzohzR1mhe7qwnsI7GXs0p+
DlJgtTSAxQwUTg/gRpyUvRalGxBhx76xxq04mY5od8Owz0sgU4Bar0HB6GMFtqzY
uKTKIvWTJaAGrElDw9BSFdXuicMARvkOMqMVnC095gKo7AKemIjR/V2+3WnsAjO+
fgqXHEu1v2pK8G7f+SxfJ5fHM3A394Us4zmeJVjd/VPCwXWk3DftRCbMofM26x+3
g+xm17QNvnoroLweKUp1axS2lZvh7B56bjdihSNjZuQV4zKDx09VtgtVG/5veIHQ
uHyieR3P/nD9I8V2EDgF5SiSsTr7IU+PHgw/ZDPASTGruTilDK78/wKP/ypxXlWg
/zSCr+ez4vBGu8q9AoQebGEbpHKZTRshRjxJ54VXTDTrErUjeOZbWpj1SSkAOW3D
JY4zMgj2ewP5iF7KvXaBE5LlI3oPxubFYAbCfLMp1YR4x+lTDYQi+qIHqcAs4Djx
NkC0Cm4wZEacjKC1L7TFHB03syINGfAV+FkZ6iH1iKJbMETywQoNzplsG6RSPzy5
HgOd10FZRIxXlZgTMXNlBresLvoLkyLJuBCHSFhycBZogXGKUJpWIPxC7ztht/PN
MJc93SM7OJmq3sGfb3FBvribpfLHdULiNaDVtva42cLwrJeXwBFErZ8hWNMPPgkh
EPjjwVTRgFHTn23fcUx4RwJOq2MUfjKu+J1e6Vjrr/53b4rgNWslK2SbDO4qevjT
BUORgxajTl/JLdQRlonB/6NyFjgONyoxbOZx03D6o/1ai7JZ5AtndffWioKifsiM
Y7pIM4dx73I7jbgwEW6bznu5nEB9KLH6kruh4CDKOpinr+hpLI0of3g5szCNXpSg
7jkxNuNDm3UZkcIyIkQZkgpb1nY+jjpWasveU+q6t7nrGedh6Ivt33Y9NDih1vr/
V6ULueJ1vsxL0YRqaZoaeRV45cqZQP3UeASp79f+eTQdmgrnYUIHXQSJrmyR1BOM
p72GjZkHK66T3RN0cGh0YrKWkjEaWiGSDfG8NpgYALD5rZ/oJusIdrpdlEnvSgxG
tCiAYxCgeR+wGtnyfujJl8mACW7MGDrHPh7JX+DXWA3da6i+AYonR2uLqCTta0CL
AzdEbgEJlbgZ8pZLHH9Qeq88Ml7MYUpRYGjK3/1VG0S8w1IgWr8qMfWYYRRDWHq3
msL639AV4cFic0wvYNeZ/uiq7cNRQA86HD7bEtawnN25+9to4JPdRGOYtJVFDJWf
OC3kzNxVnxJxCxMmw1mxufaTlbViK/c+dqMP1NdSVW+IH0dg6SCeTSR9fUeHaGnn
LG2UfmF4dXy1mTEmjfUVrHf+J4Vj3lspGp6nkvD4DjBTE3FKTQma7es9cklGREq3
N6EVSKrs6r5Jn0lo2Onm5nK1r7rbsyVNw49GC+10zHUtcrIYmitr+lk7SDhaJPAq
BKOii0RBdAi9nMFW9PB26sdy8Yb20MxMiTo1Y8Pw5R6lMR7d7fW9bTMfc9Ng0lQy
kedzBx+ETnmgS5yPVUXpUPBpdV6a2h+dG7/uxgZFwostWMwOY4Ai2Jgyzcq68rO+
jbG8n4KngxCGqQZ5UzCvMx1c1xXOQnTC7eMaSH8OjnW2o+K0QfPLmfaYRLlDcm5L
eY8WaQRJom2kGJY8xLnOiY7HMX5ozvfSe2f/O5b3Vv8qchfLMkdmmAlAVe5Gmi6b
S/2V20Bklpdg9tXjpqm0TT/DqL8PP8/3larXz7MxxglQC+EpyRYLAREe4EbymmLG
mpIHqWWr9jcXCMkC0SqN0byWrmNQxgnCHs9QgpZZJmp2yzHMimpBU5OPHS6iYUIc
vv8QDtfprpStNRs8cqv4hk6hh9EIDEseJKXlqA2I2egZOcY8yq2OvSQ/PIE/nHsG
zJpZbYKQAcKX6uLSOR2GrrxxFS8s+OE9MX4+Rc4Ve2KnX7pZxEdK2xtrPcjzHM7U
Dv0Rc858lpEOp18bl0QnXjAPCLMayfBnlVFVP+nE+oqGhIqFm93Wqaseez7VYkGx
VAK576lZ980ovWGDCpF39MyUyOp3mpZmzzS8vl4DCrAr4xuPsfFIqBbSVTmkIFk6
92xQmkOnQeKXIsV/QoxrEMdqPvOd7aouwQBxks6l0HL7az0yABI09aIez9XC9cps
E4TEX7EsYYMSxYemECTHi6bcXBikuXFcuKf69T6p71J7glgUj2tVzauLm/EvOZVW
4op2u0vi1nwZ50cp60AOynacQBYbLd72S2UopLcTwoRiwxvSpIEFiX/sB3srnfwZ
WE/1WXjVCXaYP9TlOAxocx8mK35AoPxKsGQJQRmFYthqaN/UOlbFFjrg6lbJ5e6l
Rhggev8svjaQQgmCwWBLqVLtyRN2utLdCB0k3wIPH9DlmWmLbjr8+r9LaQLUgGb5
iIEPQMDHFsaHIkDA4vKx+tJoPueSvcNa2/4SJtfA9U/fq7HpDHEtceX13RgqsvR3
jxT64n6dmdW4N7FYIDZ4P6rAd2eHRQ7D+xStd3Bs26s9eD2ZGX/87rviWysdR9SX
GRsvd2+eknvMibh+1qdHNldTDUZRSoIYtKU3Ngd5sCEES/TQWtedSSmLwc4mVFme
nuGEhQnZ/BlXcuBTRvrd+iDRFEAL5/caF+s8IkUhkceTjBMoAaYt0XbG/7pJ4JiM
+NlJalM3uTMy/j7+oK+x5BUsmvNFGCVC29vgKxZ1VcjOdiqRuT5yh4C7gbRB1iZk
r/arMXcA/XB7bo+LtXUX5R3iUTNvT6SeV5VLe3aeHa/hkEiQACaWr3Wr5qHctk5V
2nlYqLP95VfY+rxJPyv8ddbXKwFevdq74KBoIXtukj1ezHmn2czBGVXgFWhDpnW1
+gstr3iLY8X2jDNUDZSSUnW3jjS9wrOZvZLqLMDyYPMh9ztiOA14Hqj1GAj35P80
xDV3LuanBJ8kMOp0vzySH2ELDwKkVmvbJvKMdrTrADXVq9FilZQ0ieScSGSDdUPc
UYuMDeyd4PHejCVMIi8kcequhzQTEV6OlliCnma4lMca0ICu2i4lXKPg6sd4YJf2
q3BZLJdLBIpf080xrxYAO5LEQMIjRtFbc+v7Zs8KjG20+PPQ2muTL468zRbqAG96
Nj3P5zNIs3ZMGuXW+kPeDbbP8Flvk4TTcWMIXm8xGSk/M7WO7SvbKRZP+TvFjFpF
tl5mSxN9ldzNiLsOOjJPynM3EKXMPQWbBLN3EbELotjO1mK8S62FHksTxOp7KM9q
SeeCR0bwnBGxYAu/JWsgGxjS/16HNEbRGRgtAGMcFr4fKC43uwpR8Jrq7j9i6X2R
c0L4JTawpPAP1FApswOm5Y7AFkI7SFNpZywCpwM/y3gvi6rpb+8qbiEaLED06YRQ
9V1wdJuZz/VOAMS4tVhMdnv8Ann1fWUenIdW8Jri/OBzpE290bhLqwEs0pBYqpOz
d5psfUqE7gpOqXFZLvp5hxWyRsbfB2YfAD9eTRfvmuMYcIozGjedrKYgoMql+Y+C
amXZIssMdwsZK0RJVvfp6Qbd1dahsmQng2Q7WKHX+kR7VGNrq8QKo25qzYBItRk1
GKucZfvBzTZwREmhFTMKNVB1Z6CgLusngupuzdcuIKsqbL0HQNBqGK1N/7CxtHPr
/P+4OzvJO1ujJMcCqoomXsQNBWMe/JxlDoxHReFp6guJvwloJcrhcAl2pL/qdS72
tX8TXJjYHT1fJIXYPANhO7QzJYejjOZyiP7ZRmkg+mK3lgZLjLSKA0CGa4Jlj+05
Iitxd25R1VZEY6b6Mv2kV7QDz2pmOYdSEca8w5ip2qM4vskgG93a4KFbPOwSxHCL
AkOiFyitGeAgC7nwjpzS1EYlXh7u6jpFGWejOXVdD1QyIcsiNEVpvPVF2OwdJlfa
GONH82s16yDIoirZQlMOdTgVblMZujBkXeIT0P3qRorOcOry8ro0d7LOuXg2mCA+
WffPgMteWsDjcSqR7ooMuAT9p+Y3k4VkTHhaf+6UsaXqNWwI3ash8nC+mgYzyxKQ
vlD1KvNdaIULYic9MjpokIIn1/z8GErJ/y0HRG/St1zJvD6YmmLMfHP4nu0igSUV
FHWd9Y1VJS3cTX6TgjTxs6uzKAG1UlOxO8YLEHkXg3pdLzYC0HTUfJBrmAScqOMY
5+BV0Z5aZIOoUz98XsMQWYfNeTBekJncyLMme/cI4JrRKWl6wQIyvQsEKMvzYyEm
hBk8FzKo47P//tyfp3uRmG/whi4EK4ytaKJ3u7BH+M7AMPERtCYKD3ri+7KWC6O0
OSb1mS84BeMVicD7Azt9OrS8Avb9Rh2Py23EhHO/4Uze87f6R6PC/oJRl575OCJ+
zTAsVE8J6gVCyDvPWJ1SAU/+QAEyn0D105ucLoeXbK0kBIT+5Uak/zTCaBBPnaxz
YjRqb4mqHHtI4NgpFFb/uA3wScd44zmYIb+f6xfIckNAZeTCjs6Xn/j1ltUEJ2T5
PLl3QUwX+/iKRyB2kx72GjHlJv9losSW10e7iSpe+MXnpfOOIeZy2bTUOPd379Rb
48tt5+jZ+D6VKj9WAM4o+621wNGOUcA29XQbVbTPWLryEHRQZ/ZykzY6HmnI7rXn
a7v5SIhQNdtND02sOL5HDnflCsvnzg5U07oBYObtwa9/QYJqjWFqXMdFdpdV5ZXC
fVYO7LAiqrpJrDMDis6V4BucaG87uhzOrgxh5eXPVigQ8yt8zq8jZL3q8ccbOfj3
rGN9XEQP/RPvVoSc/fJ5O+/BeeuWucSvl6xDJYjlFiXwQ2XeZNDxFKlirrEI7+aU
U8PyaFGXi5sf8xUoNnmcK11OlVFs41txu6JwtBDdkMJ54MDETyOYiM7unzpa6Hnh
ITgjSHZSpchlFZQAyJVEr51kDK1tuSPPQNQ3dHk6aeN4VHg0k3f5zOxO53Z5VFHk
Vxg2Z8gvSl8G8j+Yx4ccMHCcGn91dW2PjmJcxUdPIQr9hEQ1xEAniRKr6phYyFi1
zgrFiG9a0uFPKqNy75uV/fD5e3WoocnoAorbzUUvCgnpTi104TYlOFxVfLUvFPhw
78Bspv6n2wIJN62gQhkOhAI6qNGIdP/soVr4eemsyug/O+Ydfb+bwVqPbAsDXjJS
wQOFUvEawx+MitFAQUt/n31Obkj+FjvUlv/iEjyV+DMfHWFsCcFkXfWOft8Yw2jf
Z4FjzWMEcg6PDtm1iwpDGX9/PJL0XiBfoxcoIzRWapcSAdf3wLZfOwGQXtnJK0HW
7IoPOxTMIQLxlhqHaVycUcf48qeEUyeWO6rcs7Ucb/DpWWm6//IBJ1jnaOmRrYIE
hiC84oKzjFIN1qDjTxzN+407GzU7QhYv+euHzRvuZJ5ro89b9bxgDOCfi/HCX6zW
fI1hVcDmjVHBeXT3lQREeq9gzP0byheYRZH1fKM1mywrElcjK+p/p8GeRNq/HIis
S9c1BQr++HM8xa2fWwIjZRS4Sm66raZD+kYTurUsoetXhUB6PiCq4eu2sKUX/3nA
lT9tAc+ndD/06pLPdDjSYGh4TNHVCaNlveRlkkxIzgEbf71uHIbFHZN127FVK4dC
+V9/PtBBys4kTunYIlajvVSiqx0v8h5RJVHH6CfJ8mOdgKoFl7wvJzk+4yyhtzLl
woUxIBkk6MZHBMIGDVgxyLl0kNwCNe205nj1G/0JzpPmyRQEFOJd76AWczkjcyEi
qamQnhrkhUQ6iECHdjyQV7tuY9x3M0f6MaQ6iuRt7kLvRe1CnneJVosFIjmM+F/G
V6KddZRr3auP9xLvayZlMfnr2dwzUSl3XDhiFl+cLq7H9dJZzv0u6AmOXNyBH8a1
pO70b/rJ5Q4h7dNTER7DpT6EMfQMMyAzIG45TiUoSxNnC0x2pjUkKDzmoVDHoQxb
z3Du6yDfjSitC+JKRpwLt6shomyxr7NbHc3utzMznqK0l2W7ZWgm2bbvwiNcvpIj
YrNBQLxicq98c5I7O0UUs54n4hgPwq1ly0HpG/Wfd8xnsrBp+hZWaYuKOE/hRdcG
VlmoiTocXdgaVMHiP7a8BE+tvQ1VP/Ww4umCgkaEiiCTEQ1KYCdPLsQTbqjLiC3q
PVcKyvx1zmieZzu5BYDN4OwBo8/c4sSp964RoCEXfQK1F/KTHU8h4EM7uxVOdWUE
j7Ik1WYcBtbne3TXMIUo3PgE+4EfxJY9bPsUWLCMgBESovhh+vdxQQ0G93STdOnK
ZSE4v05mhZtDNYlFzFBFKaiSCB+MJlltrTykqr9PqCLV8ll4pAWeQVM1cwkfFdmE
3FU6bQ5skS6viT6wluPNqDw/itiywEgGE9bgRRB5URoHwbwFJg9skjrSWFcix2UV
U81QVhyl5UQ9EcSkyh3j19NhFdEhz63EGttEbnPp5/hkls9BV/jlvISxRwg0eA80
lXBwWI8C4i9GZcEGl38yy8UYJyOpctj2kFEVRQtPJeQJYtszGvigZdoN0W3FmB7w
Wn9evtMEW0zLEcFi9HdSonBgeqojONHiVBizSQoP3p8y+/gFMYnQ9DZ+06IypJzV
WUxbj7x12AD4CoBqKhM23cS3UwSpiyZjnYI+ajQRjYYiLigoxV5z7DhAiuJ/5q2Z
760EJ3p7JHChzgBt0/VQWTyH1iutznCv4G4hwxrOBX4g6KxcFAzsLVpI7NkBz+aI
FBfUavdebxEVj1d/2vYFA7bzPTiRZUxzoRpDnElAbAxsVrYEDKukt69D+06HptlG
c1OFpDUVa0MDEYSx6NhJ6MLjY+VuNTeMzpv0z5yg9sbOdTU1SEzt7aNMrpLnpyQJ
9qGLoDUMvGLx2o/otb7Nr42/1uIWo2YooEpHq7Famje7BKI5uwNcoFIshAtkDRhj
3hu+d1A7az4lu2f5ACtzf0FHaqC2QvNaCGEM0O+vHkNvGmEXo9hldB8TJWSP+ttk
dQ48K6gsf7bs3+L4PdMjq1v6u8EI/KLjXhGCeUD+xRZFpOl+K+Hc7HEQf+R0MJxp
akBO+HAVBh+2MUGDCLRBRx7Krs9V81gOYJsOpmQI06Y/68b2UYqYyCcf+d4Z4I8U
MLkXh3Jjkx1GfgonCU1i0l9A5AN6Qv6Z82zNpBmsX5fbeyNQzKKLMks9FppFk6V5
m0N4bHd1ycqzDuULxYdDeofQqd7pbWEk94KNyruDi1i5x1mf3zosCYHBI5gx9ID5
r22jsGLUVxScBVlinsptRXMdaQaU7jQt/Je9KCs/EEASSzpvqYJHiQBztaErVvpE
fJwQQdAAx1veXocObTmy+2wjUph1puwiasB4il/VV0+CFCpGXyXLunvIxQTgEzy2
pWuFOkXjNIQO7kRteH9/WiD3L/9ZPpvRY/mp6WEnAMFnNXisdaFEMx6/H33Pn6Vr
Rg0E7VyVBtqvTJ3q7OLMJQf763nIALZBKKGVwDRJq+SMuREo652XUsnTW66ZunlK
5cVM/QorZEFePrIe6+R7OTqKXM34lWtFN4oRLr6RDEeJ/kpo/MUTTTvLfYXK1AEB
htx5QlF2eHjR2Mc26lPVz/v8BIWogdJ4GzIU9Y/uzcV23xXm6D4ztuduL0P1Vzvt
gfLSBUZXKeLq6TmadmRBjVyhRFHg2LJpWj4FK+98DUUQBbO8zXSWAiydYk9WdtN3
dExi0yk1LpN87/Kll5arIXUcCqsoViP4uUX8uYtg2zMg9DIeeiPyN/XOztyiBie4
2u6jJUUsfL5+pD3xVkWwm+ZwFi1/cE2dPs1mht392GlxJUpdcmcjgNhSHF59YpHu
5yNjBJjNu1fsFZaUWb3w8zDVVc2Zlve8YyyU+SRmQ4izQT/5eFwv6l5TX9svyylS
pfZvFZ4EruPgKI+7jELUYp0UIs1Nchrc60a6Vb4/spdkx42Ydi7R21JRRxS7plX/
3flsC/AywZojK88ixSSSX162Hgv7PNJlzcQu27VIdcu1GhC42lycHg/bwNcS2pbT
H83E+eVQy5Zq8u+ZaGm6uGuBWnIlAWGdgJJIqSxa50CtLiHYWacCc8gKNgolZrBS
BOB2zes065W76Anm2tPagK2jy+7EqTwD3wErj49dmNzyMWe8JDGgs+CJpsHBE99W
qDWQXsFQiqAyATB4zTencjAx+wKdA8jtLuCTtEC1HwK7jnywxsd1Hjw1EbD9OiBt
aoOsj1RbXwiMOKNjjfNmOfx9FIApFvOXQN8L1fA69IUlInOndrSZSdWRFPuF9rgQ
ErJJumTe7FSsRDTdSfHTyAmi9qjRY5Fb85ENpQdlw5aPNyySOVj2jU8RjeUx9zAU
gsE1n6w+CE7oAbqwlBIwtgRWaKbnnOELKqS6AAWZknWoMnmUJgmbu+eaY1krEb/U
pqNdPaGkqakGQVfxchOjlEFFHU9plgfNSz285RWw6SmoigIQJn16MCRo5qEUmfDq
twU4Yvj9QXNcWb3O8WMuPnTnlcKmxydP85jqNQWpAi9nW7iZqBIvuNWJaaPrtbr9
6vN4HXq8Hof84BL1h6Z53ThLbp5TseKrFG+aeu9ZQ2HzdJ7H377fLIWgApTDsruV
uBsjw7kMYPUO1QKgMlAB57/hA1l8jQ6QnFvsN1F+6mJyIWF4B/hZ92jvSqaGTMqs
XwY2d3hQt1v06FguJOUl0bFYiBQmmYE8wS4iXAkyJ8Ftl4f+keopNTIXhqkZ/a11
5u7WjxHYs8JXfXsgQjTpDRvRtqhcIuF1Aiw8OE9w9oJSzQGNU70qqaNPMdCKC/Xo
WMtfpb0WJuIzOSlyGYGguqss0J3zjXpMEyf6H8MfjfxQAAvAo2vzA+R338nzhI1c
78HPlXqUJpw5geXe8iIF1/1VXi57RnkgOccYsqXQ0nE5UtkaSfFpJvmH/KoTPXHb
qXat5CVnMsT+xHWOHeedh2C0um0BeaC758TxT2fu1n95lmi/YVje7y4mQPZ7LulU
nrntxmIEj8cAbdTLY03spOMcZiiEfpaMyy9ox1wGNFCGqXeo2QZSp3OxHMGiU8ON
NaQn4jKR1FI5l7/BLISkSqH+V1oEc2p+fzmX4oQ0aunIofaify9UEoLSfVhnzBUr
34yS/vzuPuEhw2+1VlZPYbcaLeKR6sluon8DGKRyzzn+NvzpgKVUnsQxCvK/bgdG
qgLqX7XnLbOUauSgeD0rsR2aG6+TLy43zgG4QpFGaFhN3H8GIjKDHeiYFKnzXSSL
X1uOSrE5ErBFwmdZor70Cb6anpAO95Bg74SMn5ixIUde94au3avv5E/pa1GlD/xs
+mSAhatDHA5dbqZBh6MOqVucpEX6J+F+pZQtXzcQ45QkKSxIK8Qm5ITfl5AeeD7K
9h4nmL/rCVMVKqaEZd5x757nUHctrQke1bUGTQnqVvXUY1Wkm/BytfltbJOTPKw3
jA8Eur5FNIukdwF5CjaijFGQ2uJyRgF2oaW6equ3Bz1Dgx8pkVd1bZxBdj3BJQfx
Rq7k/iJVUWPfy1d0/DY/eNw3ggSBzJw9p9U+Qqys2Jw+wvenfMrG5XP+/X3JXSMt
2mYjbUgMkTouulwe6mYnafnqC7P/qTYwBZ7ckjYDTb9t1SWxGv+LobRl2iJPDB0B
3qjzXodHz4TcIgexkLWtfhLFEXlwXvK1P47te/Tnt0W6vvoTGCXRzYVlp1+yQoQy
XrRfp9a8+WKNYg33eNvgI3hb3XlTA0Nrm4YOqfnjI4YKNe6BrKHYQlypLkZt/O7O
uHKYDftPHdEwShGr/wpIiKocqndYx/YdiM4JRXXjNVZxj0sYAtmtNg9JmoE6VhyO
QmFx4kuP4D54YWlYPaFYpZOJ3qNti4/7Z33NFeqde2AA64ZdRHby14Ax3NjaRrnZ
rIDAEAbWpxAJV5uPtsAXTMn3PizCZ+4R7GgpY7whpyDy+3DgDkoXX4rAwH0M22um
/RhXoNv0gUgdHuiwQ0BbWx9U9YB2veAjODy7tZJh7RLMc12I9mEu7Gg2lbNcuio4
zM7vMROeFA/2vqiFdPbZ2+CL2ZBVQBqsCfO2Qc/O2ojR8z+VaOawRdKhDnSIiFPe
RxPQAw1zI0BeCWRC7yXE9Ar7TWpkGSy56u+Lyn8QQcGCK9eS7sCgF8t5qdgag0Yt
04n9nUDKlDNpzsNUbbTRaeGa1XgpQY1oa89nAB4QjICsitK47XL1UwQ+s6bDEPoS
IzGfrbC+vvmIYDM8Hq8rbfnwb/fdxzI4cHzRRj9IQV4ni4IMoip4oq5tWbzX73io
B7+dqb+nncrNA+XVpsYLtoMlc1P382FHwt4ZZbTeQOQ6gRPCYpJfLLhuZuJUJ93y
7FkV+fAcHHm4zjEWpTRuEXFxUx1R6EjeTkJXRVtfG65Uv5gz55Qf153hBhAvz/3I
Ibh8aUlEpiwnFLbe2bg7aYuaIxTjxu05XgKSAC8KLcUtPygIcaDprcwh0XOduUC6
t4zSWXe2Q0ugM2ZohkIatDz0lV2MwJG7VoYrse1RCgZC7A2aQ3APWWVdvJjJCwtO
lK9OCFAArhV1g4ZcYV5yKoxLtedSHjr77RJqVYypbL+GqiU3Ya95watoElSZkbIF
VIymyTrA5+Ou/2vAhCdLBZB3tsUZNFa3+6cRyZZGOejWxABCmvj4rwm7H+zOov9J
JwcUiUPH7YcL2G65RT0c10pvLlPjBWbmMBvndTqfePpIIWabxNA/IpCtgF6zKjCS
uLhbRAWlAY9ntzT2tbS8OXl3EjEU4UmU5lTBdWuSRyMZlI2VpDferyBSi3vhss+M
4K+RhxuZV/+SfynGQTuq8erdf/MJaA1WX3Jqx7/C61cLbW5peXN0uqG2W4ZEgVt+
zIDW225ixz45VBp6SpHVPZBwKnisMIYsJCwzpL1jznHlPgEwbppQRJm62025DlJ1
gJGqyvjZKw7ejmoe5BpWzYFW2dxyFTbWVj/clIay6cWTKYu1Bc2kYIjW7wk2Hdf9
OyV8XwlEdA0VXH6xdWxDSFYKDvaNWxod27u98Akboz21opB+O563Fk3nElVEsmmZ
3Zzg8jHKC+nC1G7PGbjrYTxP4T42m9fMSB6SPE3XbYuZtR9DG1OH5WucLLa+7wwq
lOauYKzhdKACd7EiVJbE+pAcZu52M4pB4YYI6saElX7GMHLjIqfCRBXXGaLQd1H2
+UPWm87NsQjP/vwE6WgYXBjaBAB5SKHLsi0/h0iiLJW8gzX+OBs2wP61o/obRAWy
ztaQCyEM3ICYTZrXwQ7fSjizxWwh7HaKPsGZNtIxp5h52zSplPtNpb920gMtHrY8
0ZJ82at/ynrHg32pUdkXzxj6RolI9BzqrMjxgYXpzQNMBV4bYijeg7kkIJ3kgi+g
hXz/rSoyjIr8mMLYmiRvo6OvaI5Y20MMCsVcbypAyULRq3ulgLy8l4CPmgXDFG7v
Ro3jHRna4SGL/LrWAZtoQPtu1LG45V+iQWUEj7IOdsWwQOH9hykj5NOJNyWUDkD+
MirN4ROa1E19SuUc0mWGp/vTWcH3EJpXcKCkpds+XMfIF6XmA6whL/YLJ8lCr7ql
1OSqUM9EhvkIeg8lsRSsZnJqDTmJQhnAq+Cylai5jbRlW3dDfSZSB5LZsK+KChvJ
CXFxRWiNoArstFHe+HyJkeg2UePm/WJMSpUG/WGoX+8D5y7gJ3vzFNlyveeMMX61
s1fTipptuh71DcmizNTdw0IONycagu0gWFwkN9MCA03Vavj7I2tScI/dKDDeSraI
xRbWh/p/T3Ut35akRkm6jBx8uVI0AkVvSigMeOmW2UogkpzQF7vdUUxFBvr0FIyr
6/EnTR18QC33ysYn80ABT262UxM0xOk+219AUTyUFfW3nC1LEqSVU93TZi2zlvjp
R7iLUTSn1vdo0+Z7qJ8lugeyevkKRaRmZrBNYXlb1rJjG6GWN5AN3fFXeGVSAFd3
us6WFnAltuRkUX5Y7V61VHESAFYNbckWKD9m/W9yOIzcWUT6eATyllzc8PebIU02
QrqEIx1oBZ6E0RJBGjUCFaD48QBSEvjA1Ej4Q3sibCtqJTcRxY6sKiCgJh/+oGbD
Qq4D+ZsHJrpeS18pyucM2NdGlM98oMF+L9succG+RoW3vQuKyYcoJF4VeWDN7xvg
Xgj1iNz2ncp/MPXNRa6yKYOUmPG4hPJ4SlFBrjUyg8SLotyAg13z/NYByE3MzgxM
q92nLxNaQ+Hc7WpL6rX+4pSvs8PRMSu27Fwa1rLc20O0Ezq/BTGHpR/32iv0B2PU
5JChLJKXiGkV0F7ZIy5WxrVlVh2UfkUzmuEjfpCw66uxJkKCa8CbUL546TDXijS9
eeh1gWb7XttmYirTve0XxDJp1qzqYNqIxrTVipGQ5v55g6QxwJ+m/NUEV3iu5sPq
j4P/5H3fPtQFPQMRbmIqTOhxXPwasDg+ohxnp+lDOxO1reXq/hyB9i3Vyn7OoB7y
GnSMPhXaba0W0V4Ol//eLxYfhjjrzEIt3cfdsCgY9pdgJYtxIaZY4d3Is3kCCcZS
l1lOrrQatCMS61/dZvT/9zhsd7OfKRP13StwqzfnB4J1SUaSHF8j+TuwO5sERdzY
XpWUNEHXJisztQM5x/t4S3pcYM9QyluhEm8zFUIoOlhLpv3HqyxHZaSmkpmAxTvv
zfqgXnX7KzEChsKF4HaqmuZDptWKk57e1jsZqrvx2dmKxL6q/Q+Uk+qxfMxbj6f1
Bk/rKGAZfb1TPKEC2YD2pGK38M/G9b6H2iMAqQ7ueyGWPXLVuXbpD0IIPSSoiYu+
9VhauLLaZsLwxS75fXeaCy5RiBNCH7aqXaU6xApV0yn7PHNQC1lgDsLye3FO+gCQ
JcodtQ0ynXByDTWy1l2xgQCpewj0B9i2RHfveSsG+7cDIfzuYnCbsXMytbUU0Rq7
oeNWqyGa1O6XFXK6rRRu8tiGmvqUNXATvC5n16u8/7NQiosRAnwpQn7etIlHUG1E
KaBl42jDirVCm461R0/OdhA/CDbRKH2hzpGblTa+sUbcJwoZm9i83YXk1j1RDYon
Ab+D4RM0dtzA/O08R1z8PxPAIUvqpnTZT9tpo76wBImkFK0EiaX6rbfO39+fhNS2
9jiPsjk1uGaFrw3C5/S2+7BztUIYdDlJwibonQ6dBFwtxyVByPFgZgTPY0f77NQT
06DFbA+KEjsDyTRFzLllU0XUDJ7j4BMApL11RrkRmbhf0rPlBZl13NdGa3uyOsP8
BmGfXephcEtrHIl2xGx2NyLWUs/9PeD3io0k9gIPfcngREnLBcXJY4Wgu9UE3mYJ
O1ZC0/GtBEK3nufYwxVZ9uKMB5opkBMkFehAdrj97hznscwTrD1+OwZk/+Q7967K
vtsqIdUO4MaIO5auUhNMd3faNL5AS6BNSgukdbG3S/o3N0T9ouGZf+zBmTkHgAxf
uMGR49k4ShkfwM/ji8aYZRidLbXk+f+PFBrBcaGNCBzYAOVKO3F1EvLtYGhJ8Tmk
dfxXiYr0/316MYDxO2wMhqBsD3VfVcE64ZBATZF7gZ719wbsBxQMhMjx7HVPBsjC
j8tUX0TZA54JlGzlp35NUvJaOVjwKBpyXPHCTTGHOtZDlJWxdjOIbs4zCbyq1kcV
sWdbFphFxZnglTvsEXDxlx0+QakiMraslL44YoF8jaigFQZob2LcNjqHMNR98caq
qSCtPLStPzVJaS6VhVpPNQkIe5mLnK6YTfgSznllu968jJfvraEpt3Xdimudvuf/
EQXOaFgEQXklqj5fbspHPVlEUYaqY/HO/Bct93XQAaQsaulpwsPWJTaq+hoy9pBu
5nfbq6lkfN4o0OmZ0njMTdfyCcuO1NvJhXLjGJqzdGZOl6O/GoX/85BX2w6TRg0Q
qPdU9eimJZbOLN/sOBT6T26I0irqXE6iXNuc6lukNdjP4Dcek34mMerRvFnjjgdC
uMgbBtdeui+NR60cHWHDIo6pNp5cK7R0/pQXaeH4NX8qqW6Rl3G6goNYluCsGpXk
BIBgrYc+4gMICTlRnnzpnrkGxTjZG/eDCU1cYtlg1bqPLHAy2k/gl3PTaYWr8dWi
ElX6o0gcasm70P7pfIwngJzt3PaF3OoCKovRmvOyCYr57DUquevFnMtPrZcpNM1u
EXwibApLSL5RZ3avz6SDVnvJk8NHedNahFFROBLZUC2W4NPPMr2wFq9k0ztD5JMX
A+VoIMahH1bn5WsO/u9DmpGb4GnJSYi6U3ysnT7GlTGH5TlB3npnI6eSaeJjIwMf
xfaU4A/k6F0BHALXpI+2S4a/BUQdU6MXd969Aq/71CSoUjGAWw00pJ6h3/h3aW7f
CCXWa1gR+SKjB2JZzY6ekAIZBuxKFdommQzHm9unowfyzpebndPfRSBwP1AUIDgk
e6FuwuX2DW7jPT9mvuaLgrjxYX1bldFo0VPDfVgqTqmY6odQfqjSMLDRv3h570DB
FOQYNALmZ/gUJNJlcqRnujhviP/dsn2FyZ2As8klDSBnSO46nJ+HalMXOFhVGFjn
iKKxA74ClJP3I9g8JCKy+ljea8vRplmSzmYimTZSuQpjrimM/nQDpTD8ZSnKsy94
TgQMgrUPiodqcFvB/IaQh/vxSyaMCCNob9R07YZ15FWQQ1oSwGsORz4+dyWWRNm8
QyBhOzpsoI7PGesBmULAiMt+0dVsPH/Nqp5aQMmieIaq26pI8UxJwfGPJozL9POJ
E4LPZ8aUDM0lw9KPyhEMzURd7MJXOk5m/xjQwYakCvSBWMR35KHrkk4BTvltbhBR
Hpu8RmEhbaG6tenNYFsL6K7k1+9vzS1ah5TnnZkIR8MOpwSk5uoHpy95sHbQ1DXX
SymgZ/erNOG5gFejMOYBkPkkyw+xFZP75JICcGoHa8zw9nxdNZuIF8T+WsUE9K9U
0enwoHGrKZCfLEI1osmPsgseix8ON35CtQAiwIwkSauDSCCZ19BQ0N+DjQ4cS0VR
ikq9xdeE6AOp4TkkqWSnYzHo4/VqY8uMvr563gzQ8kRsoZ+qUf+AOqNon+/roODH
MseAJPJt9mCHbbW5y9FNsborXQEPSv3KegF9GvDT5nqtHutREFpUzmZmnyr1FL+z
TMJb1IuCz2nIzwmjt2vHyE16CrhrWhj2Bb8066ui8pCR95R3XnBC0zxMZ+2SUCpw
TQWlt+lBcOVeNq3g0nEztE00R8hyNXmS0kEd3mR8FIFT1l4XSSUGypRom4RYgOTI
2Ts1GO0TtMkZKw9e7EscGv5F0eY1GHK5zqDT7m1Yulgh0xM76Gp66XPwKFDCp7KX
dLAiqAxjpTd2pOgNWrrbvvmtBgpz3fZNzJvIfUehc9+/VkVCtA2wXT4yhDkm0a3+
fLFRUlCQJDXagHBCH5/tOFa2SYlJZgwWbX9eqlfmdR6WL9hd78oMuAmQKxGqr/ss
fns3+6uH0toRysZWJIehg9E1qP17kLgZsIS8Hm4r/irmqmvfI7f7LFUksSIAe0Jg
o9ujQ/CeABKlSdIdMu05XT/iFPgEQr2ZaNzhl9qANHoPeGNXvUo8tRITvq0Ck3rr
NoyMvTdxh73uOoU/7lywvLqG1uM5idJsZulDxnVJHZ2cywnqu8fTH2bj9mokEtj9
+n/XxZqM4DNN9uaRor2JIGLDLzZAc2j3he1v/frQtBpyAKyKhEbFAM+jsvD12OZ7
E0v0EOP6D/htNBt7KiaUIIVajY4TRel5zFenODZ7xQqrm3AKRtechkXZYaG7i5su
O3U1ApUwnFlSqrYTxg4BzyskYN8dll0yYquuOIvLiJ40zuNJRnGSPhrQlApwkGCt
BkLk/CTsCU53m9bWfAt9u/aHt47A0dPMChPSh3FSznFvkaq0WmAbBJsvJMHi5WtL
6KaGFj6t6TC6RQ63VK+KwZdOH0wgf+D/0kBFsDAuKQZHvFE2umBjFiV2doM/Y/M8
gq58nt8/1SbNPuecX6+CUAQtEVVWDGgrHj7hc94dk4KSuuhSViJN4vNAfL6cws6u
XUntA4W5w6DbR5k9OTNgCDFBxF8VZNcQMxwqKctcnd+eNoviY+voljEKrUFi1E8c
48rl+QZ6DBMA40w10Ghby0RTQZIYCJWptIPYxkNnjMXM1IKijZIdkNGuc2KhMiFu
ai9EAifqP5P7HasTRihEfOiGout343gxyQinJBwxsHMH+LWWdIlAybyR+mZJfnUI
aQVk77tEA/0fXKlbqcydA7JxMiSMuNJnD/vBpotN/CkOTV52e2TI7ozcNFWsPLtY
gEk8ybytVjz/SyKTqphsTKLImAezB5caB8JaTqVb2TQDhXwW+Q3LSo1kdxIcEkT3
q+RsgS/3+z4H0SyC9nadUgsFSupB+6vUMiCLKLiSIZzhyUvc1PFsxM3xV0nhybk4
xZpiHAVfsFyWpT9EFnFl/KuCZsBxqjlzmcfEqNRjJptnPXEBG7CPVV3udPhHy9NH
N8Q0KONfFdgPa6+ZWRb9ACkpu/47RhQq9JwhftGYRVTvR+OwziOaBoWhfWq+la8Q
FQMtBg2BPfQXFyo74dul+wQwq8SgL0OKat+P5uzWJaj1Hx3rSk/BblVoacXdEv0u
PGeQJr3ZN+hDIkooMclT3JpvuyjTGWy7aZy//7961EQUh3tJ1VVmIgXoe4vLRejT
ciXqGstJFIu4ncK1c/SutmrSZQcQT5yjnq0V7SWsJTh+GqdKeO3lsb3DZDWOsqap
Vh6iukz+S+BYTKuneFmN0BIdvLeXk3NX6n6NkZDQvkGAObkpgswMolMzaXJL8kw2
nR7FfgfiElPq1njrkvatZNQ2pRIMtJl3RdOEXhsONkHuqhKnpnHs+GhrWk9FrBrP
pXBjRNB74uTsh6t0UbpSBy5Wh5KMqYjPAoYXIUnaUrsYQKJHmoeij/C57Xmjgu0G
GomwaC1suqGCSXPP4VmmKJs/+PSp+NiFllBZpokiBRUJNuFQ9q2HFrUj8aYvQ2CT
3Dj873gSj/YSRhG+yolNiS+L7it1sFo11dtF/5ZSeordXhZnQ6Vp+WBXMb9egWN9
BtKWMs1ShJ0uKmKoxpuOiSNdMAgi5Klld2VoCHf+d0kPYs3cdmbj6rUPTzJzSL5H
cS8kLuZ7ka0W2k/R0aYuK5Yfp/m8WUYhVDlVp+NtT1eZLnH4KP6sve4Dory3f7fH
aZmLqumtsskVpmk2N0YcgsfEysNTPxzY04Msbp+vX+XlyGOD2mePviSeJfHTSQxp
Bymt3JlNKUT5A2FVP66PVz59J8KWTsYurijB2tCa/meu1vrbGAmLZ/wlbdkvS951
hSFbrQTa266OAcY7dms1wNhvd1/XBnex8BtCVveosO11NYqu99uOBICEhUk2BRc3
eTcNMod5gfT+MuNSXtu4fmkm/QwoLSDwE+glzsWoaSHjVeQRlPA0nD/oxsbRbF5X
X5ODeW/cTCA/nxULSW/SOi6f1makUuJyittJoT3+LCSZRXu4KpiJPofF+pn+DpRj
Mi+mea/5vFnN7/3KqUzdxtob3HT0AwDxuU5u34S2kT7pm275nS7D9wh8gJ3d0YPb
TjNyrwv109F8/gcBT3D/4zLceVhm3laQ0750kOD5AO42bXKd4KNT/dygxZWrxklk
IYY74My0CBLvCdjpuQQ0XOcP7Zg0zkjrNoHe0uthc1xI950Aboe1C/NVWNwcFyLU
O8DjHFHzPOdkLu9Y54sfO+BmEezrVVRxB7xrsibCMyVgXae8k0TWEPt+mAI1UIWK
WJ+ZYLPUcQJGwEV0C4tgSVfSne4VkFNtLb62M96YsaGKOrwySfmmaSoy82gJXNw2
YZP3bEhjEA89EfzjEoU6K35aMk+MFQZf8lmH5pYTMiJbc+bFesUILdLLUCsolF6O
RDWo5jG/kKaNFuUlIe2BUstR/iIFleG/5oEXOuDcEMQ5YR77ZSRz5ZrKw1Wyc46E
sxHTccdikZtb/tt1ZsGuDFvzdPyfsaRdMQ0GiAAdFp2OqYLGSYQAXwT2RnTwyJZt
gwkWyzSJwm1Ckt7K2SAu9PooLdQYd35+9yKCLwTToluVwePQ27E0DZapGCJyLEpY
8bNkWbKiNi/+zeDg18qJv6HzDC4RpJejRdCb+Bia69lLVVv5GL6zdc+35y2Kdee8
moDZtoAjsByV3ZucSffJwECqFczAkkyIExvEiJmCQSFGW3YEETtvZ8Ei/ibeu38r
gMp8otQwMPr2ICet6IBZozFVHKxJiq5KgfyzbXGkfAMC0+LWg8gGyzY64fooBLLH
vCUxA4cHuZMUFO+zQA3C02ixm6vWrslqfCURniMCgr7gDyXmU4U1etDf2CCRsMJS
gv8MFxTanFVju7yGlMq31nODmq4E9vTfjkgtzMUE61TgvPBf3dQI313LbUnchWes
PaeZE+EhpY+6+dfqAdEYtAu/2n4/0DP3jJg6XLO8wcH/HvtxY9i61qtqrPpgviTK
pOQxY1fa/OgEZyuQAW3BV2CxMBbyxbv1EzCLsjAGV55quecvYVDkHt/L44l846xf
TXqifPd0FPos8XAzShkeiNeTKqQewILEFT6u5LQIeokfm3uBpHad1mp/9xWkDF2K
anxCs6VBrF1LE8XFn/nroAI/BzMXop8ivn1wDgo4VL+EfytqCIFLRuU3N8ra3z1A
XB69B2blBJG92sIbF6B54ZT5d9TdFpdNMl+nlTGU4Cwp5ibe1vcvwMM7QfmbDBm2
UvvC5t8uhF3IAGHQqBa429pv1MN0Hn4Tee/s/S0jDiQD3Xc1dRsuyDBYbd952Wf0
x7+oR2zAqtIguYz7xn76zv8Rkaa9WW7MRDXI8JyWLxi0PMBHYivdel9nAXYHkYlm
muDOIpLDvYqUh5t2xNavEXR3/y1QCeQEKMI0bMLY0vby6Lgzk2MYmRdtqcdk5Qw6
VEQzAeMfevUq0wmpPNP72oUq2dtAZns43rdOsaE6KXFwTHspxYDyMIntNClJtUe4
P5K9sIE+/8xUUQhZrFeOVQT8Ew6OhCIBcHBT00MJCksnV6joCH4EAiyuWgiHFKSL
UdnB//ATkgvg2vU0b2ep1c/wE+tIroPyfCpIadlVp4p4uVAFcUAU5qUzUuzf9Ang
mEHgM1yK1h/0uorjTHDwPJYkVnqrUaKz0DGFl7vhH2nOFFgMjE2Zfv6qdIL/NLOj
KwBmshacDUGUx0YpFkso9gZtOOY7AulQDRYfDNgcDwvBjYqBKGd8TW+TwjRaVFMv
oel6W4o+ZUE7aDoLthyZ6Vnc7cBv4JUGfCgdLudoq6nX5fcP/XyZ2NZrgAZYLmwu
azLtabScsp5etmkVZvVMGPlrEPyfVxv6xRM1egVBT1hbF6eBoWAj+oJC7MVYhCLK
CZqfaLZADv7poNNx735sdkUOlPX3BcoGA/+/e6MCcuXGm53QpMqCWDntJ+dihbeA
zAtAYcdiKLKBjb7f4UgnGtOAAZdQuxCrGeuQ0K/zRFBgdb0vqHF0trhXjwBSekyM
tkmlxFN/VgqBKP56oiqZITGgujINYxzPKSe2hAv58LejsxkvfTif2D6tX7Iyt8q0
K7xGDySKBXF9lcat5JGZtEG6qgHU3SFIlYzy9Zd8ciQDXHIBvRY6uG+rWv4oEfwc
GeawKC516o1u83s1FuMMTAL7V2bo4X7zoz5owJA9x2NzV8dSuJveKKt00G9mBhOj
WWivJFoUJcn+6gecjgHpatCTv9+b7y6j/HmhYsLz5w1E2rLFe/mjiGbnvhIIWO5N
lOOwEWk51bYyEA9dXrSbH0gWoBui0L0vN0APqiiOh3NuWSdMapUILAQkkjF+F5Vh
YBNJ/joDZ/SVUxOWjIy7iZ3tebScBsjPMm2r5q/CsHnA3o2tUjJLzpio7hmDNiCW
bejOWvkCfsf5QI4o1v1D7A6OR8tuQDYE+uC/bz0Mrm9/t5x0P+leKy+ebLSJC3md
SAL0cXpC7ik2AiNayvZzqrv680Ahybxn8RoRquxHgnX8EcqMHOYaP1OiGlXwdxAX
eu3g2lLAlZ6EX3yrhROaNMaJb368Q2PehDGIhP/+ry54EJPkVWrnGjGlVzjwndOc
AQdDUc1gjsbDAWztWLA1V88HokT0iXxk9ckhZL3qoGmY95/0tATscdbXRmndwaR1
a9RS/lDfdx4iFZntcZMFf334mi9TULwHL8WR1QE2NtsCtQNXRwRRk2j/j4Sh83O2
PbBGsIF6pu8eja9+f9DFEvDzN/beu+PcpxL1YxO/PcWr6ZLFUIjl6t21pzpVm5Ov
i43nC0ky0jau2463OK9aHPk30oHNGL5Ul92EeXPeZW6BaVO+FXCg9WqHWcsbfFEL
BZZCXJ8RylxrzoQ5wxh1LsZq7GyKl/c/1dSJJEwGwMI1GSaTBz9FOfSfiTC5qS1s
cZW9iqHN3i2ctMWXwc6fzGtecW6vCFp03st0NNvrMKgcF/sGe4lOcWtqKivmz6hv
49gIFSoOOZMaUXxCRaYV4AuY5NfXzR1/fg8afl1Qz9hqsZ4Jm5gXMB/6gRxbHq4l
Wtl6UVEOoFKsnNv+LAX65iksz1pOR4sqrCrut4OX1qSqsXabTkl+9Fx9VjUgbGGC
BuT0Lqjx+KFQ/SE4HzwYyK/5dQyFfQio2ev831FZRR8I842ABf0IQAll583Noyy7
ii08mHEGtWxg4FRmHu82V+r/TntsbAmK0xqZhqIwDV5FlM32QQNTlsuiMefAVhh3
V98n7rOSCYmxzkuWyLLko606LP+G0ZdeokWgG7ULdK5vKajj15x1T5Cz5FqaYupi
D8kKdd1hqVlRqVGgpiqtHs1hlnZcL2rf1ZAAAPidYTrW+jLXX1I6JK4lImAKQdvK
/sLFDJEHgYT3U7/VCK6zqdX2KqYzbuo26pOa+8TpMdjTt+L5CxVuqwU/gAzKp7M1
0cqvL8iwEUj8cYyMZb5aCn9RVa0WUrpBD040NZr8xiO5ccGUfP4CPNYOAyNihp9h
Ed33EJ5d4Iy0Syj9hERHGRGxNfjG3uRhor3YRt0lqH4FqEKWAHcteOWOLrtODFA6
EE9bmUZgTgB5QBO5Ur2xYSYldLhxKj+3YpsCT7TTnxltBIMVIjxC/FJsteqRoZr3
4cbrlr7ILFHed5vpUcrLJV+Gn93itCoRVqX5sNqxg0dlZ1s8y0eBCLsspNsxOReG
cQmqz2NwOR2f1XizN/RzxDMEi8rLiZn9rwKWvrq8YhdCpiciRn0mzSOSccTbzrVI
k7MgX5EVw4U9zfIRyAFtXKSw5vkmFfGjuhEa/R63yvpD6tsLFS61ib2+XXzdsEWj
mKWIWfgYyDfdppvioRUpEAfG8WFg0ziebS7WKBW9FjI9vWIYskUQq4yhoorN/Yix
enZjzzOfeBRizxxF/N5JW8p01jjdDOG+jtAuRBmiSmuEH8ZZEs1PL2V9eGFA/tTk
JkF1A7p3Gy+MsPDA+ALLPs3Qqesu80KTL/c2+9ThGxdkS4WGkwiST6nE2j4XLpch
+V8YYF5JmXpdVIFsFLPEeralCRyoI+0cbhvp4Yn6hlv2CbBbzZt9fPHsoQB9SxUk
OjjlGlmIuqKojFvi+fVN+hFxLw2NA2mQQ2ZLUqk8zh4MX6PTF7Z1wZrSnwg6Enmz
3DGrdQMp+Etl+B9yPEDhNjlrCUphrnaxHDotVt5CLwIJ5eguq8kk08HczXU/RxHb
xVnFdpv2ON20SYsfqmqWpkxrdWKGUzYpA4mayQC+yZqXVhtq8CXiQXXUJA6D4vvp
HtJ4yt/Q+nFiwGIk9y0ydmCReLcy5obVBG6eUwyS9zzZMRBIwTuJ0gF5unet+WMF
PXv9zwWAeCUAKHWvOYvIij7bKZv9gc66jxv8KDXqVV9rvNHVjc42l2oaVMVHGBbK
1yIFylPxwPhRZ9tv4JXpU85tFDp1GzZyyrbo0UFiF2zyS/w/t0/kFkkUbH/UrNZn
o9+VJRL97AdD1c4IMJjgf9vvkyzZ+UKWJcNnI7rx1iAWivw6qkGiiTKhN8vGxlLP
jnJ2Ygm7wBUtM3fExjxLkLxjtfP7io8lep5yKhA38ATHAPGFFT/i0nixSxCh1aMk
c3eNkP/0pxzcw24ri8bnPwfDpGfxaQLdLgrt3yrrLMCKMJg0pRyfeMmXpeXNRX4U
xQsGFV9Td8vvbuF8rRBZxYDtFHQQelUv/ox4IbL9T9Wi6hwbUPj7XeASJL5FP53v
/uTGd4dYcC+Y1SIXQYFeXi9rlRDSHxwX+d7DXVgSP6T1fOmcVUgHFxmdWeEBxDlC
0ju9eRAVoOmX05oUvL/S/CLN04BSMJZxw/+dE7CgHHICKjH9TsITKHTrB3RsUI9K
gccZBD8qetY2HOoCzMMIlIy/bdehZjs4UjZD1HvhBBxsWJ8YkfFU5ZSD+6vhIog5
Cskt+z6/BhpKdJgUYIKOctOngp8lSlNf9JkPhmo5liC7cv4IXvCQqIxK+d4c8KgS
DX/h7YZvXB11tT7l3ju0xZiPOVmKh6EwRECI4o2fOWaF5vwvwo4X/v/0NuXvhKZC
9tFXC1HNUBTeUdaaDXM4xG4yhlaX+jdjx24WKki8o4uQuTEZ0lQZE63cSG8KB1od
Oypbtg3yWroFACOKmz4qngBC0GoAD2arpNGlfNuQYc02f9nGEMqZXiV1Xw1c4lyc
/RB5OZmK4Yim9xlzlU3F/c4jfkWY+1T63slIfJuNnEXeFufNDdzz4Pv87sCrYfxr
vIPD8m6rZn34AL0QgdmCL/Ut2rBayyLaICMQx/eJL8W0YTDPYFDICSzZwS8JGGUY
V/kif5k5T7+jSvPOf4bFCENoeeyxHIu3wipuO7BHoHWN/hCKXCVrm/7wLCbdl9RE
XLxnDNwdBv1UN7LQn+BHZc65ZbQyMX5QFGe96ROTsT0zpZxwrZyDMfZU96hWfPuq
MTtdYjFyxeeJqs4M9e0seuh1PMQRGKG6nT3/Ok5CVywrYyuCglQRHLiBMK/SVkSI
8gbArBGHPf8LbLBoE74cajGUxlwDrfdNBEIgRyZr03rkI1HCEmPGYxPsAmtEGfkV
fwllWBK0A/f45n1U5eFwvdqiJGUhR/Tqwgx48tRXeWw+n5dCHCWlVwlUlzvriffW
GMJWQrouC3vrDY+RlwoU4u5T2QDp+4fezqA3Py+h/F4NgD8Ci6PbUiwfvOBaCttE
HSV8sLtiFXs+pVE7T6qltZBwGPHagZx4y1qGGSlJjUVcEULg9clFBT4UHbEe1pQz
Atn3OfCfzPgZqw0V0f/vNWvSDR/Ieido8AMoZKWTq5LmMW4oG9XGn6gvWngCmaCL
en5ghaU38vfAB3Lkb1suagFUnjpAsJjNtZNoSCl25Xfm28yifZAsB+bQU77Lr68/
yWyUUOq9Zh1Yw37FPgYMGRHisdgm3m9aiWBaqQlVG0NiM4m1LHjwh79gamsQF5OB
WZZThF+HopRuAmq+SxYcTk2Ydnjmdx7Jcpv7nmL7REWOVBrAb6uUBGSV8HIFwPw3
qHsjwksbLFqZ09TIKq8GUO2EeLti/MAZjyriTHvAYL67ZFNn6m/UWwyThTnsEjQp
fTPRU+TYT2k8QbNR5CF1t18LMGgw0Na9nHtvqY6Ix+O8PJV3bInbLOvPriXQVWg9
1u44mJXuMktfH3J4fDWGjFoMTabIUXBmG/ln307SFgMgo17BL4rT7MOIK0cPzYAf
SezZkwzqLRlszSdT9EAO0GrqWAGFSqtIjm1CfEfeuHmnJVSpk/MJUHN82BxWYmCQ
ACeTOYDotCt+Z8IsosR09B5lAzxFHGRP6yvT50czeFfYS98D6JCUcigwPeUW+kA5
ZoDiGcATTsmEyFjYI/rsk+hVytt8QnKPBzjwyeyeNOSXmOhzLTMmYDKVLtSpcNQJ
upw7jdAA2llxT49WE35mFnqiwkztiCpOz4qdzdftwfvsGpfoJuKoW9YYNTrdPdo1
`pragma protect end_protected

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
o6HVEaOPO4oY5R0jI/gw+vovpuSJ2BbYGwxGGWYJQMePcrW0coE5JUNk5sEIyhl9
gMByBs0ODYg6g6SEJu8QbKSG6v6vrFxQwY4tu4QBpNGAcKxSrwv/2nF0isVamJY2
fnZZFy4vFh7K1pk9sMHjCUi4sIrOhlo/0L055S4VBaM=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 10768), data_block
DjBrolB+k0r1Z7TrYxoubVu+c94QkNXCXziNUHKpL/5rAWanQpp5NKcOw9V2dVMs
yd/DDwD4hQmJfOLx/S1bLU8jltaXMxuY8vOMK8+RCx6MwRahoN9BfJjOeS0kfdLs
gheOkce9ZJRsF/RDozN+1E3cnyjKwd/4/BWwpTA6a77oynlaevdSUyIqCKfRAxP2
FZE84cDcpiMAxs21cbAKQ3JSCR87S3FNW/Fl2sTABpIW/YDhqlF+xNQoZG0UW+I4
jJGofdcQjpt0hy/JuOLz1dBE6WI7cB01Xs6XBZ+ke7fHP6oltt5W+ZkErXoLHDO4
90J62kM0WXWtVlxhRfLvvzWfIcBfK1CyClHYIW5phmovHxsf9YgsQB1+qylKiLFG
a7/wSOAuutJRj7QtNZjk0y3QHMuWZZY+xuGP/p9fOaBz8Y1AU0jriPkPwsl1x3jO
vZB2qKdm7c1Sb+D3dsZbb1Du81uW/mUELlrOcI7xYnh3gJAoueIx91tXd4prKWw4
rIPIStHRSpFBqnwfhx9UtkX1U11TvQ+hVBY9h0iEy876lFFuRkp+1T0Cf52OLoOA
6t39QlwuOmQVEssN/WULjNrh7uQRF2KWgZk/pYOiLW1kcSe6RT6nAs3YSJDU9ToN
vH+0wZkiCicAuyHvrTEHOXfC0Mh25Pt0OqD8ff3Dp6mqThLJVvMpY3YHL4fm4pQY
FduCqMohZB/O/q+l2oR4rco5colj67ewe1jdyeEcgl+/tumvi5l6dGYaPCcjQyPZ
jaJG+md0abXEXx/mpytnEyh21ZIRs56hKGAPA5N2NWbi9v7o+MLfBWum4Rkolx+Q
z6LxmgdmIJNca4nzdldkVKSt6zyE7MyMio8S88SPsG5qzJJKKWgbtCj9PBiHD/W7
+J6LNNVdtakKCZCZSXJSeFbZ2QWbtNV5EOBb0D1mbo6GKXt20y6UhCOG2rpFpRnn
+P9W7JF+n0UGv40fkmkhe9RdQHoZgoAH0F03lBDSgXXwurXLpfVL0sm5TcAetg+Q
XazJxyveKDCTBCYAJm8JfoHWq53NKiXNGRnCEQA+GfD/WxPXIn2W9ey5bav5q5O4
q3PRDghGE8dLOSrslmj2SwyuSEGTvn7LXjhLUu88WBECamXAc8hTdrl7t7WBExXo
8ekCC0SWBo7J5dNtuejzY28uku95s2bJe2Mg2sEIrkNTnVhjrJd5OxqRW36Bmm3G
VAX4M9oMQP+Y5ZtawStgMIY5eZYBj7TKjjoNDbtlxNqynhmbMW8RH5+wvSBZsml8
SBQWtfMNZnH/z3otdjMYOBiojdHXiFwyYJxVURVTsRtDzLKQadrWpvJCKZUsE/Vc
wkEs6SBCvu/hIkfkj/hJpZjI36xDBBgsZTiwnvZ/wuyD94WJ/4MC7pz+pT5hGlEt
EGaibVWnqgXyHSM9UeP8/ZyS5IuGbae5z/nK7UUkRFRFichdGWyIUZ39ZFi3WujA
mRVeUAy/zSqt6UNMBwmQgKEcodaUtfMP/Mqnuy9I99yvGU6gbX3DH4KkIZ4lFRTn
WrTMVCeQwbUZ1k40p2PAc2ec/CW6P9ed1UcIIOW3N8UwPG59ingb1csLLi+Kqolh
uEworafjS5iEP2YjVxhWOO6/UiMvcuB4uDE6iG72rm0PPfbpslIOjm4vNGJs1Dow
ifkZMc+kOxUmwXg+00A9WlPE4ykFcFXkORqxf8S3qLVoEp/L2cyGA+LSuR6AAFYb
WbS+KrIaCVWQ8vMVWDl2M0WYv422jx4vcrdJ2YZkdMZbaTlgih8s9GP3Ou6evQif
3znH9eIg9hMKzKbmjts297yUjWd9RJw3ogFK30g5i6lUd1uPRauNPE4BSOlPTgn8
aqtQbXZMIrdphnXoyl3XjK2BAhC8H7thUpLq/arfI8AonoepeVqnGqTEg6zj5IiN
NGRVaUnfMzb3N+gYitBq3i9BFvvp/QCWDlQQtIlR2ahCwSL3iM+8vBECE94dFeMl
IcE7QazCAyIUNl+jP85rCCkg/sJ9fyuUj9PMbQo9fmjkpG5FqIDxGxvE4wuvyDiW
71oZ+LBiSE+m1jFHIogXsGKtArmcCFeP48yZG0R/wdsikxCY+uixe4jDqAgM/hg5
VNUA/fzspyL1qmux7I9Y2P2GrCarHNEXDaO+EZ9ue00xny7win9P48IjwqgibrWv
smgXL0DxOvGQn4opksENCthi8HrQFw1rGAkcZewkOnAOb7jW8NQjkvUbDgUYXPqu
qufkWKl63ok4PyTBA+t3WVay/y9Bi8OTY5l8uAqAvHzqWxOiLoUmy9s7wEVKMyKw
ORcRw+TqEJF0zUsV3SyL4pX0udpCzbm86eHgjA2jaLx9wiLU6uL1StKqwxipbBVz
XESCGA2YLVKJPvvWOmghSLtTPnnOXWhlgv2Dtu7UOyCpqqg/Hum425S059wYmAkQ
HjY9v22QZR+t9i7UYMxSIcqT+cyXfjAV6yqxnUG7aSf8WuAIM41rNuGK7422Efgl
mJv/hXL68R4ISsH3ZoYCUIKadA1MpUZ0I5KGC67RdKbfa7lNtaNuBnT07jWNpvpM
GFLUqaXT859sgnIfnwuWxxaeFTBVyhXBN7hicfoZrhkuPpI+IRrlwAv+yDzP0ka5
xLnV6u8FWDghjSEsoj+z3lm+J2sL8Efsi5k8Mb02xI44P+8o0ebhpLASV0x99jH2
cJyfU16erWJc5lGhFKUgaUxJCqu01o0a1vb/mfGJxFw8K729o+hHdtY04K3olRmE
hbgyaspkEF4y0XtdtqPiwS/Ux79GI+bbcrcl/mLI3pPNYgVN98aRZCkIg1u6D5us
izSWmnleuJQRuTMbhQjPtbEydxsZVkSDkhNibMiVIYcdN4Ynuiq5LXL6Apj0/0a9
8P1terlJ1kQleBaJ6GG7s5jd0Ukp7h0B6Gibosq09ibgEEKOO1TOBZz7TaU4/lnC
kgIWp3tEm3uLi8I7WBhZsqFHGba6NMOX577BfOi1MwffRGA1a2snyOtNRkV3cxxK
Igmc2dhvgXay/3fxRwfIC60r2fxl5h4S/No4DLukoyPa9gm/ehZgKRUYR3vDs1nD
QxExLAQJ2Dybdmyoe4ig5cHDwslYNCdYa/7fyrwqEhHHX7yLAluJ2vrSimUKaexM
wmo5Qjt4Sov41GzY5xh6CIK0PLuMwSxBkttG9MrpjWkbkwsqBxaZzFpA+LIo1pi3
+oAQwIbZnqMFrLO4VjVbw4rUbVm54SdSCD9kmKeL71rjn6Obg8ZEVR8HbOe3AXjX
gSsCxr06vRYLBnMkG7nHp3AuV5I6v5F2E1WSqbqM5VkJ0nhGWbtMNZxaXLeG05xd
JhCuqX7RE0tnmUHXRHEZMd2tINwtU6Yc+cSiHvyh9qtleIxJJnrobIE0uyVxMTdX
QCIUGXcJDusck6emozPbs+NbfPNYTHimZftuSh3M8u4BPEWJtq47kkxzr7zge4tN
dKe/fUk/eAqbl8L1hO9XYMBDTHj2V8TcDYf71u73iUZjX+Zz3xwymCZgziDuWTGx
irlscRyc05Z0OIr7tsi6d/sUXrkoAH6+rrTIfxjU0KsPdcIqZb9av6d+BDYdRecW
CW91/EcQj4TAoPxlnwoiVahn1mLgFMQ2lfvy0Z+yoncR2/itL4SfPCPAcS3pNqmq
TYxZZ0p8BzZxrQf7JpP4RngXKJce9wfROqqVKLk8wfB397vuVNNzl0oB6XxKfejM
+ledse6epBQaRLZTVQvSb5100N9zvsa7D3igzE7oaNZW9xqqBrOKEIwMUXdT2mai
mgwofsg/PQ6yQpQ3DVHQTaCRTDaAV8n4Px8aAalywOsyqiG8DuW2nZdqFN5saE/c
RCf7aIvq+6iixklLWTlB0ht2MVwlT97iuCFTb3vI/+FX/Ns2IpF2mRT0Z1ZYdLne
eKu/Vo+4uVwcKFjFVWHHHZHjfkLrEO1fVJexQp79+zr6eOH4ythtHGDn6OtC3qjo
oDmUOB09kFh4WfhDmH7XmrysrXBNCRPdXwDa8SwhD4dxMHQtaWzIOQAqZC/iZAYs
R+bnK8wCn1uy9gpDW0yfe+pGICs32iEJ3jj1AAE0CCYI7En6sMExxGwGF3OZMs+5
0hEQobnwyLlEa9GjjcgTjb9KX7cAkYm1Vqhm1pJLHYYDrZPNl+nMHhrBiFnhPumu
agZWRZ9RjSwl6PhB1Dqu2XG38fQSkLr+Zz156ghNnkEvNZ5GYlXzJvAYNYlt4OTh
T1kYYBeE9xB8SP9AP9evQguJgTqXgbowohOmtWPZwr1/ssi2waYGi20WZr/xkpXK
mBQmBsE9YkDu0gtV2nZn+o9mI8VbvLGoUwVJr52rn2LmbHtjeaPRKdNmFclTMuLR
2TUCdgxIUFzxk++M77QlvCBzpopEGPJoqF4IC8Y4mKVoyBY/P1k4EwUPHwetEVP/
unNqMgiKKw1TvK+sdScuGC8NcB0k75bFE8fttZfbC/QjXkzWXOYggfElP9p1Tpj5
Vks+hDz/MgE3tzXpdJoncK1pitVeLc21Z8AeulhqhCVHVCyulfnw93QaSfks02v4
qJYXqQlzZjZTOv9hrLnnPjOXGpNQ2/eQB86XUZKlcmTvyWkx/yKbR+d7R6CqsBNo
4qM2aR7WCQBiRBK7rlAC9L/TMqCTcMqpy2eLAZw9MjSslflqMhpvA0b0/Z9Eoljl
wRtirwzITj/J3yAe97sifwdx1sL3NY/tC1HTvewwA5PieqERpScw9i3VJ2ED6phq
YsoNEc861MNuJ80q5t0W2hUbdODaZAkRQ4eY9KZkPkGY1dkw3wlGdRqds+gYNs1B
WNXBnrWwkuckZjaQeDvJUJEMMnNDMmOfn8oSzd5nD4Cg2dWlIU7GYMuU0twcXZRH
K6gw8U1gBcu30La2H0DEmbByAiFkGaarJLhdAN9BbXfF+6PhTMd1udV8Jgfs8lZP
4N3R0/2XCUrNAXVPvul3C2fjGG501+qpxt9F1QozT8zk0NBDrJNsJMF9B8iveZL7
d25fB5o4z7fHYbOoHxCu02uj2viGiOd7ur4WVBVRrqS5PDXGsyN5RQHyIOFBgYOc
s403SiKEPgMNFi4SUIqdyBF6phyIVxNexGnEEmxNjKaGKPXEPX3Eg+Y4VV91Vaia
XEUtvoEpnSWJNF9z93jvJd1N66u2WaaSFfp4bHnzfVjFALzV9hkNJSgUsoztsgWb
sNNqCx26loJSp34w3W2u0du971O8GfIAfH0Bi5ufgwS8ZdynNsp6prCU1HwaIbK/
Gp8RjIDQKv4nV1Sx56F+tL/FbCzadj061aj88NXeQ9RdRcxeZUxwd88s1tDgRBIt
gDNzifdL84TO3RJlFJjDUk0tBvRrDou4uDjxTPbNBwIytRRt8nvukxxXNJkj9j3/
lPwfEBy7wW4Mh8WG3b70wam3U6jyT938PxssmvY2zCpGuNXQfHAkuNZ2Z2Uelypf
4I+7aWDkCl2OtD3GmGRaUT9JWKlGS9n0egdbvRMcTaKV0JZiYluoMhLxo5xixqqz
84fmccPk4j06fEcq+godCk/I1yJJT/SPLyJZbdJkO2CrHj93cKjMlO7G9bpg8/Gw
0m8CgOxtJm5NEdm0gIWkEpj0j4vLCaTYYcAS/QK9TeUUCFkAXozH8An1LLkdWh/A
5SP1WWfV4McdBUJqCPydo97Lea7dqcdiylUfLizVTiuhHM5ccAWo+BMsc0/9/srj
T9qqOuRNcf2BjRtRY6CUsf9pDiUJgdLGT43n0Gu0Dm8CyaWvx9ntpYEB2xp5CJ0+
pVfTvLRhRAKBpm+Lswnoa60jRGbz9ibcucENTU8fl106SqG5TMu7twsKWtM8E0vy
u2zxDswGMTsJYomn+Hj0Ul7hJuZDylNnsOEaLkP64leC6NJPe+2fDp0jQCoNzq0O
OHXDgkHnZIPQNWJq7HG0tzlBq9hK+mys3Ce5Z0zkNYi+fjlMbCPsyfrWgzQRUos7
PgFh4/7iPQLIqeFHojkRkeAnqtad0II56B9vfxHHDOQr3BdQqhUlrMPzwj/gSMVQ
2uF0jD6YfTxlgLz+c1Q4LchAJvZMvXJ9kwQR5BC2tPEHxVUbhxD7qjzw3lTfNedf
zH0DSXls+rBacM/nBQztXID8gEgfPTvHOFG2VaTfQ5nRVUDyUpYmNhUkw0XgPJKv
rP1DrLRH+k5qNdDPVHRYPanN7HXoE8jQd94I1GyY4paq1p+VZaWVbq/7RszYBN9E
K19xLOX4zxyEZOOZ2uin71Gq/PO0oXSym6euVYVAkVpYasia7M+ZHvvGVB3sKrpS
Bw3QFy2gMmeW5MHPyFz4BJG43Dckt28kYqPETel7M8Li0fZAjjuEufdqONhitUWW
wvmFhvnt3Z01nMloVXnJeY6NqucLz0bLZwWZiQcDRksnAq6YtNrBsQPsIHkuQBgW
rPHsLTC6pwleoJhlY9EHWrGUC4vlWo9ZkdTbiyBx+3bPAyDwJ/LD1LDTUZTzNeA5
50k0Ugi67KiELMJk3hVPVCHHS79dBsAW0HO1dh5AV5vcG+8F4S3sBlGUMREkHKXX
1i4t79qj3czzHN5QHsdXAHy07xf6vbl6WMLU8svBu4pwXidoVgzdc6Xh6NHEojMM
L9hEEGro+jNm3AgW98wQSFu45vXw9/c0Ft+yMiHlNWw9EhKwm4vUli7f2zXpjEgF
lOZfKPUfJJnxM9Zo6wktINCZERxsSOO1pjjM+oJVUuYYQ3IrD04KP5B1SVuWrHJ8
8xJfUbCFlyhL/fzOyd6LJXYPKZjOIQ3sgmiPmNtyDCji8OolVrDonVycZ72bF/8r
TwDKh2BZiSUEDMM1QQj7EeQMVFPaaq6FSF8XisS9I8z7U3V6/sxOzO3dElQgxB+R
HhHGGzjNYZ2ra+z/MV11zs6wH/yq58movggewmDk2d58AWITfa8r5Q17RRDm4RL4
reVW31pZed0I883fTgXl1P2fHHu04NO6FetVo0WhLaOpZoZnxs6iNZUSA9hhFnoo
IPhr8k5ZrQxPblIgMyG1G4x5bcIWQxGbcA0KWnr+xixOKcbj1RQxkhwqA47Db5XG
EFsHTzZdDItkwlm6nO7lXZ7yDjnPNEOGqJstKKqm+oGsl9PbuNIkhF78q5zbZhfA
vVIAsqFOc7JbOjDKgw0tQUEwCXPuTFIlVbL8eqzqnP1E3+WAnizpN/46T0Nq8Dwp
H+6FXcKV0repBI6YuPnoqY3Q4pPgQW7aOZHaOhwHFUDNP7DNq/BfJAxD4KUyR7qN
D9dyjcyvNuMHRKmfyGQ+D5AwH6Bu0emfMLmHH4HT3cv3ywMylpWWAwYKIC9YkhCa
40kwnKzhBlHc3FCGmaczrQCgzx2UDpYWhquK7DrD/Bl3JW8oddZI5HgQlgR6Vjzd
iTkcLZQxkeHJvUIfozkrKznA3zIc2vIgvk73QRRMkhTuRN5AjCxF+BrGDK+vXMyr
MXQakiM/ImEKZfeOfHBlx31rrZwapO/M2HmnrM90gQuoLKjmjaaFQnx9JhL28iXO
eqj/QLyUEohF3tVsY6cbrkZz1mKzkoQIWw7VowsjFKbtrSXMNA3iODhWFFIaGFSZ
OBx3jGbyfi+kFA0m78/zoaIEkGFwBXZryPE+aeW1eouj0d155viCAdTU/XoDE8JP
o/U4Nixad7KPzsP+mRx3cglJyBE790G0zB8l9BEhp/wpWNTnuoJ4AsKY/Od2/Cpa
7IzOI8tMXnPXbnIiumwXNISHSAH97yul3OCkv0PlWXGbavf6B7TkxHN4rkhpWkY+
qpvFxrSWbkHSZtGAifWPtnN17lP5gc1Sges46rbPBNspmGX/UT5RzYmr4ClfCZkv
hQs7CAf0+Arf6fe/arSS76mcLiLhkvIiiQT/i/HXbYbCBdETNU0hF94zFILiJ5xi
jFsLhjYnQlxbJAbCbUMwVyHLdn69V84gtIdsa6hsSv/7gu9RL14fZ7WUxeOmWNkf
dnmMA2OhijAN+lUDHEUVPyfhYOupEobP1qUWPNm+QjF4nyTLtssO/CZ5/t+KLOfl
Nm0XgT2A3BmtwTfMwispJIugis5j2tFwDXW3NzqKBpfBAxx8DRqRl+G/G4FI36KV
m1bS4r1t64RCSZQr9tA2jtAsXCNsvKocx5pfKHBTZUERR3opgVF458pKzKtoxme4
qLHCa/RwxNovhUQQ5zhWh19hMEA//B8HeJCunGUR0bbI/p+u3kFCzYR9K2EHpnKC
0nsQ7y138JBkfoiZoTsNQASySBQ2kWZ8/azT2Cji01bKvkw3ARnt0us89qp3l27M
n64pQWAUTE4XiALFlrEG/29+JUSPOEgvcKqQpAjFOFj7Y5ZpRoutfQHobXndMW2j
v6FMf9IksHjWG3Fn8Iv4n55CPgux2F1CM5NMc1IM8TZSgcLHvNQySpeoCIXXubz5
3iLwlDaZoh0bRdQPisQHXcMLqFG14Mv9nrXIt1ghJuvCUWyC8s9RmMGQjo6EP6SU
ebEJ20ukmVEEz3SSki2f3lR/0D6LvITO6XOXVX1k1UpZaLQACGBjfh04ber7ntGB
LIgk6BG0CH//n9WZ1IskCI3FWf+cKtmRlXgpTytN6rikwI223opA9y6/y2CQ3FU7
PoLQk4thUeC27KeoLoCTNau3dFJqht/6D4KgBMJUE9HcQPPuBWBF4sTpFfb53jje
MmekOA0aumBl+rUHhukPnYG7JB/OugbpvmJ5JpUnCM+BHaI/awkhkVgfmCTjayML
Mtjt2d7xF5PkSKl30bNHgjJd9w45dpwd+uqrBfFQqV7d4sCyBE9wuBYTJ7uor3qC
LDZkSf63pY41w95EkSXCNJkMyUn9FabJk3msBo+hfoOzyrcNI5nPDT9c79oXJhnD
iZRH06voJq2m3VDcoPKvt1hCYfHfQjJaRKD2XFGZckx0Ff2w8OqwKvwIQH0wa6pg
pzvtaJMndVD1O1a8Tj/9hsn2JlYC2RL+SZuJxhS4PwIA0qUU7njyJL51mHI1YGk1
OXyX9VLSyjHjiSPQTn62ECDUQazlc71rW+H9bdX5NhEVAoY9z4+wje9P1mI1gOs2
/YZo0eyIw3MgoM/YNVC08SArGRqLKY6YDdw66GvtKH9zfOLjU5KjaMjWvWIEzMC9
X0tqHbMD9bLbVfV979kbu2H1BNbNxllCIPJsyBp2f0QNoMuXJg2DeubDquBoeObJ
Pz+/yQwbLbkywpSIqsS5Wgqm2pKYuunEO1gGU6VWtpBfGPwgLVRbrlGUW7BGFS3/
p7ex+5NZ98bgtInsyTmaxTv1MqZWKW+C9sDP/ONHjL5lew2Q09Pf06WKx4f98GrW
tIhcd5GbY8TMrB1MJF0260s+2T60G1zPVEr7BY5Y2db0sr8icHl6N5+1ehmmpxxI
J7P5+k5aTnbIlxQzR0pZSKeboOA+kx1wQkwT7jmGSI2XAawJWEkbHYIkyq8OgOfC
oZG1Glhved/R19FumTWZv0ezQNVcIFJAS51Qj1gRzbOE+HHbQFnjzct2KOZKqIaQ
ZFrpJ6+Y0RzovsEZ/VWSd3e+TjG3SL5gS72fNlExbmWoSYuj9bgHZbnR25JllQ3P
QZP5hYDwcLA9f2pb7ihUXBh1nr788mNZ3WAswAUmaJ3qRdRBm7z5l5+zSJiNb7Yg
3Vj17ndkpqp3FUP7vxnWtUlBcPu2R5X/BukyggeBKAOgzNVLFntx7+aTtxjz34fD
8DdbzRqgkts6T7rKvWlYTTfAaN9NCUpisMCzjCyhZHeJo24LpcJEUw8Rki4cs+wG
a+93EOm4qBRy+oE0lSkPjsF1hK69goS923mTuvrPQWmefGuw2c1GQNL3pf44RkbU
PGMiu7p/0VrQ2nEAT52ZOPI6m3XhbYHi9fYQni/fHgvebmyeiKnZZWCKihFcGU0M
OFOL8QCCg4h3IOMpyMQZKMYp8L9MMa0pLdyaU4TpG3qw4FaN3xkayc66USnhTQdS
S1th0tiXGBoRd7135inFpAK+apvjfh4+LRiXlRkpeI4xMjm7NJe2/wnCGj85gPf4
7NykqRkFGAGDIrvBN8CFkvofiPkfM6XY6p7haziqH9H7axSUXGU09pu7PAEOZs02
0LzHlRq9Pz3PnidmLfPhPXlvi/sK3wf7lWfKj8FdZUE0aC59z2W7n+P1GhIKCy0r
wUY40LaylvagECmRNCaEm3agirT8VC6lXfkKakVmolkVcOAySKkGCc4zgphDYTjh
D7P14FP2NKeMmqt2shaxFXnyOlVNCkf+FpjqLi4R7ZWzaVh0HD8cUz1iwe6EMwnT
+JxnoFZCYcsEh0bzWQdV8KzrWtB6Iv8b2YqZ1IisTgb5K3OYoOYr7eNNzlaezleg
6nOvc3UK1GkSUntvQ2p5OOx0TT8lHb5BEIsj6XuOYLPrwHdX2VrhWuGH6mUMjX4B
GfalaCOMXN4ah3eP8iCXo5Z4bqLTgawByzzXM0FpO3H3w6XMtIdWl/e0nk0VZCbL
Wji1PgVB49S38RN+UDwFCzjvsnWoNh7Bg3GstUpBUlf8XhINxWz+H5jxOmsQ5WY4
8pl4twhNqu+H/jU9UeNOEJ/RrJyK9EgAccr+rikNvm9Wpv4eVnU31hNTFAXdR66d
iHhdxHBijpsivD2dxJzT3xve6iqZo8kgWIfyR+UODLluQ9RP1Ywt99emCBIE1Lq8
mFaVhITniVaZiRD+ToByDAOSyZ1Tp//zADc4HmiV+rvuXw6oEDdarFQQNIqzjwVU
hzJe8MEIypa4yMtV4b4hEynRHfetFrD1kFk8tOwhuUG7/KGifJD1HcPr1NtUihvG
8ScZsV8diDf700iS5iwAr7aNsYOSx0BGjSpYeFnOUKSoEf2t6TiEhwnQNqm968TX
xJ2NC57BkbilELgS0hTuUfNLHuZhUuRGC9ztciWuZ508cem/MGzxc+v6egKCFdNr
Q3Wuew2OB+tRYVI4AwGZ9s8bv1giGg5d8vUqzZHdVrlrqscODXpomN8d8qpmyJ77
Itwi1siYRfayPNkNFgBPkw85U+z/FNhPSNQ0LnYt7NGeWq8prB5w2hWImlsrbsTw
4/9V09QPiK2bahrzpip4d2pzni/QofHjNinvAdKyX1Vce1yD/XzYflkI1zXEWq0D
03vWxItG2tCYuQzQvBjoyfnygGAJsW85JoLIirNmSiETuqU932djTVEIomI8F7f4
AH5czrMNhrqp6Dxan9DjBiTGby0IDjb++/j2qeMDouhnwDX1zF3KeObLVM8Bqo60
ef1h5XV6EU5CWwLRtDBiBaY/LL/cpXCaeQUrAaro6lHMZaHVliiX+P4l9yXBWuqV
WUIXlXodcW3Zqg9LdGroBVObFUo1NkcuAMFbc+b0QrqrNVOBdBbtJHTepr+QiiKf
8RIxtM9Olxk8XUktrBzRPF9i15ffcergG32Er0TdUD727eURN3d89S87MqVUFy2P
FX03zRgWb9vGYOOLuqignxvyVOmETJOBdfi7tPSTvJHljWZVHHXMVmGvJM822rls
Z16SLX1H86RjVJ9I3lT/aGfwjkhWFq9N2dDtSpPPYfn/hplBz49MMccrBaeOHCj7
HIehVZtRU+ZiOZOTF0oyHHJwih9Fmo/Dd+FI2hgpq3YeFEH1qLaaGNlOBM7w7NVC
yrpOKPefHGdB5JnmLvrCYZ8Fawe/h9KQL1bnb8G0RstaE2Un8IugSGlTP/weXuqD
5BBrzCk2a1tOFAozqBdPKqqOmWDUsWLUhGzP7EvOGfXRJNacwBc4A6oDTYUuTPNQ
uaXe14L+UlF6/j27g9U2FQt0ctecBbpRYuSWETnN2ZOZPuWreh2ija9yY/T2wpae
ddwurVhSa7rIOnAfGWjsL5UoUs4WHyCEB4a4ZP1s1ojfYdwpXf7hnSiH72YDLelR
wcVlpmtX4M6IsIVTtJMRMS0UoaBCjZ12+na9m2WzovikfDkjDm7U1wNcEz0fafHS
sNY2csxdEAGaZ8/D7GwtvZqmYTw5rtaXDJaOs2IaF2OORyom4Wm4iJM4xWrjF3Ze
F8HM5JKAKryAFJqQQm53mojIGXgGaA19KtHfz8v7hRrIIs5G6DEhl1rAa4MZzhT/
yQsabEwMPT5MiN++Vzkr058tLFwHYJmCQGOYapxtplTrDK8jxRaSwbBIrZIiuApz
f+dG29XCC8RepumLm6UvX5Dv8MnTDfJyyEgAFeOZhI6sPR/yg3Q9ZvpUlWOZu3bw
j92P6U4A9Lrca36fUG5Rsukrg8k87l6KYsAKmmoo+qqONMoXEnecWKWdJoFAK4ba
fRGdM0KZecpHgyWp/IzuzDgssvjLR4vKqlTV9y3bS4j/EnUFjzQ4W+M0w429xpAw
fOBqzmeLw+dcM+O+kqvQ95VPeduNDmw8WzI755yydH0iknzcoCJ8BdNSx4yV0t/k
oY6h6806XRw3J2vYuBcjnTVnJVl8kcpZilKmPN7gpa2nLvxA4geZA+H6lp7S2+xs
00JIi8i/MIivfAdHGamwR4lIgj2zVwl2P7vAQIfU7B8ZMnaWeTatWcb3i8PwQzLe
jHCAQBjflOJmTtz0xh2TwRZ9jpqOtqMziwwM5W9aWWw5zq2lWZryRI/BqAbLIEB1
OJZgAWNUT4Ex0gDd41wQM08BO4v/eNLwZFzyV9ZYYFNq/zOT8I4eziQI+ZdLeqP7
xecylBUja8LPNGTyeduOinkG2WKhevLSL/d7ftb8ttrjeSR0qrH98ZnHSBIze8ih
zDjPcczsrrQKv8Aq7aWFm57nHXwC8ZpCeN6ybQDS+Lg23U49a5LHI6jN/eHhL4wn
Jia7mT/rQFK0L+C20yzCJlAZKiDUA42P694Q0BKPL5ODJI5iUD+l/ItIPFwSNVtw
4Cp37/tP5TLB6jPgbFj3QMrmvOiJyGy3M7cOZN8VDz3xwfyDxTfWUFig4sUrZzr5
LaWR20wlJAtDsLj0yxiNK8o9J69DDOi7KbEUyDDZ/kFFacNjiVWgMd3tzJi+u5z8
4s1RFfXzgypX5MQR7SmKoeAIfneMnWddpJ8jKheIOWFOvI1P/gAro0o9zlLr3Ovv
R9CPZUfSGjtBerJo/s/b/fN63EtD9YzpT86Jeqy4evHAdlK28G6H39h81W5Z+/iC
7rio2Eu4bl5U6ORyKT95P9WmaFveCiSq8hXkEJr7i+uiHzwlhRit7TQymgo1x33N
9A8EEU2KQ91HxPmrD0webkD58XF45Pr9ORRftRSDOWIGCYRQdVk1xZGYfn4MMKGT
+lKlYt0c9h9SHXqcM3uOUOHr/96Pkg2HrKx3eLw8VM3tMIHtZpqqnQsiRJMjJQFV
yYD3SNcIDhs20QwejxrRlpAcwfaz5Xa8qTAKgE71fuu8bMjoKQWVMmfcdBq7qagD
yHORlSvtn2joi1PzhrB3OJxIZPBKUeDldRPxS9Ws1p/Q6uv+oN4EWdNRRBcpAP2E
sLZLwb+TJ4YmnUrqMCg1svh4BQtUgKbHgPxF4NMaX8JcqDqc9jtq/niWGd6NBacT
p50vfCf5F2IRnvdXHHwvJ6CuOGAk5vpTlQnJTYWmCpee7wO8GO/W1BRnCLPM99ex
sHTWDCnCuIZ9Is4bJsCB8/n4zjQ2vOqw4U9gFQbrvBwoGMOm74nhebRg/IyKjb96
D6snsln4cmH/McMlJFWxJwbfVt6sKacqVqVfvhEs3RqLefwJXDFVLqnEL+1qUpZ9
0J/MH6qh1pyCHRU9eb/ksFPuvASTriSYM3yemZ9gyGlgZydTgPw5VeHpU+pGRWQ4
p/Yo1TSU+Rf6yxhs+cTmhfcQtbrrj12LrJSz7jxeDBu3ycQhYp0R5PYc05qRwlXp
Q1kjA/H55sBVbQzxQot4kV3unh7y2sHeEM4yDFTSeM1hFsTZF6hBvZ/Q2AKahbIV
vYrvV/WBs5ANhW4nbbIzaK1rb118tKhzeepc8er88dncPSVPRwiR5H/DPf9+JdgH
mdd/ff7LoFlTpG0dmXco+s9803bNC84938SEaYvN4QKqEAsVuNOxxE88IltUKU68
lwgUaU8XQNy1l6y0a2gPt678B1efBvcwzprI1jzsWz10eVpPE1J0Zjp76qpARQXo
rvT3VRGcXGpOBeCrqeTOSBLfkgqibzgW4xDCyCamtTFKm0pOhk3cbL3qkrr6Fd5v
vkw8qz4OV5qvuyp+8tPdsOWhTJHaKJQ0XrqNmNhJpW+yRgGf7M3LvRZthzBGKC45
CEEtyazF2SInwXn8xDOvRd238iqNj8t364FytP13/arAZzz42QDqzMXMWF/0lKu+
bZ9Sbpjve/FBuzSgq0FQWWyvAVZnicoElrlmuTOg55CYJuPHaaqo/9pMPL88/HEM
m7qlHVraJvqTiq6wFWGBQVuQ78ar0N3MMtQJGqIoBXx4y7dXhY00CT05LvRsn84B
XzGUS4c56BqVP2MbvfmTTA==
`pragma protect end_protected

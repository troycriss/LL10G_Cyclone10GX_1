`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
JK6k9Rxd3NHw2MbRI6Jl/lb2FWjwfFkubmsUS6XyKmUaTfU1VNUzn+mfwnp3VFLB
0U92phY5U+jE7XsRoD7+SbW08+1I/omFk85rstPvRFyvxZ5LT56ILVvqDgxE/JxX
562LIZ0qnX4YZ2+ekUvY0wD5iULiISAmPrrnn5SXhlQ=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 11552), data_block
btVJoGwVlR8j3qF0om+dYEBhZ+BYhrQT6+doIyasSEWpVYYA5KvYIiz4mpqb+Bex
yYlRZ6E+qyrgZ/5x8n477Df9ufSNSNxBh4fHtj8twaYtI3kQtveaCIxQTGpq44Sl
DwcUMl+8HoDwvpvNbfTgsexq9sn5KygcDnWwReRcy87Lbgb4qWZGNIImnKDDwpIc
vVRi/LfF6DLs0y6lSu+NmeSo7EGUApYaNPb0uCdHh0sc7aHaSb3QBdYtEPoBLuHz
BYoQiTUhb7KpIXjaua5gUN00Tz7wmM+suvD1wZQ3NcsV2IQI4FWLso65S/c9xtgP
/k8vp7sFcUqsG/tfAPNAYGTncZOizV0OwUX1GrJdmq+Cq7ZzJS+DbrQG0j/PpkeT
1kHWttcPW6DyaKAaXWIrIQ/RmxnAMucxFzex/EPn8XfHQlrug/F57uYLGvZmPdEb
FhNBYSCplQgYwnRLLAZR8n48prLbJoA9OkUHC5oqyufWs7tPDmLfFS3AELnu47bk
sfsa4iwfbzhWL3TF8dyKtsh2cFpHj6RlEAQxMy8MKyvFteUqeRy4NF89el9R1sGr
ttgaqwuvCYtm6baak+rppSG3BCC82TAGvuqHzepI0vjQnOkH3qkuMjldv/P9c134
qhEnI4GegT7HTY8rPwk4MfCXAI7yY3TUjJN4AZe+DI77yJpm3Ak0MVvxW8K3a4DX
n26aNT9GxrcTrBa6LX1/4tKliMxnI7l/BbkeYRBmeYCVWTHddGqSgfKQDFVZw75u
DFTL2wuPtsvfwAkPl0qqqFjLd4MBAPOlU6W/Ep94bRQEKWfVuFwCrkZUJG87r0So
eDTKWhSBSnIzB0Pl6t1DNy9G5ZiwAdI/4eCaCsiBQtt/7UGC3XDQp++Qtp1XLb8g
qHBQrSPEenWOIvdqlmJsEBkuQblqg49G58iDEONz7ICvLBxvVaFAQ+bl5Nabnr3Q
zDtrbHkIvt2ic6Kq+glYySzLJkOw5d//+JEc5DQnKVgwXzXWmzsd24vwTVnOcQrm
O1BMfOYO8FeI5M1asjP1WCxqpFacahiiugQhFKPhOsClwgtUCVXS4Q1O3C9Pelde
HL/x5fmQrBEtmLyY/hGpVxyQGT+nl8Sno5g9K7BPdTZnMvqSMDI2d0XDbgB+qPTU
8bVNhrsd9l3RblDhE+kN2x7+TOlg53LZxXI3gyaMSuzsAl3iNu8ZuhKtwFXP13IZ
jq3dUbXmMq4hWZ1lJgzyasofSDH5rtq6h0t/XPJIkwMg0wV58AC0G0prin3BbZV3
64K8V4e18e4tEPudKk5gPTiF1Fbw7eBgrkgf1zNo2PQ6LPWkeO/iv43fiDTC9zq3
J0JvZjzlw30xcEkOsRywZOc7qT3k8DeA5GZ2REQhX/8ylLK02sjz7k9yotctBwBb
xmP82f08uWSeZ668NOAEBoQJ3s8B8TjjYD6MUtgRfnnqkNfi1mLuQ2J1BElLu/bJ
NJi4dvBG25isrmeS7VWDr2Ezyx4N92hGh4vp38y4D2OU78If9p5UduNT6hCfNUrR
efFypc8C1sTP/vwyE6E1PjS4ZxLAAQcCfVxpZpLvW6WtBniSal01YmD1SJlqsYnW
H3F7XAzotSZd5fWOuqJ1koTD9C5+T+WfWXTaTGXI0XOM6bSwRfKyg6g3RGlfucly
dec/CcL3U2bl4w9k61fSqbmf9w8C2I1qTKVLoE54QpJWQAQe8kibgC+JadQ8fGNK
5Qt2nTvEhAQFhP+VBm2R3WQuToXDZEE3sBRFXeE+ehjWjOggcywnf9UtXt+tfYLh
ybQywISGTPyHJugKFBg36d5KewGH2II+cZZ/j3eJV7EKx5hdsrqdf0P71ZGvqjqW
th1f9LWHfoAsL9JxDsLisWM19PILyjjgP86XkaHQS4OZBBbLopX+4F+ui+BGwiQI
8gBrJ+4oF28Z2+4lL//eVR0BqtR+4vAnLsCLwcTPyWjDN8lVCyHlOYV5PFBB8xzw
kRSypSNaRXbQJYD/27yCtqO+FJs39s/GziTGtjdj+1LSX5G1lLLrNEvnr+Q/tskW
GVaIHFLs+UespnVsJj8zG8RuaAmT/M1RD1ZTKMLu9patC0v0ahqCo0GPwzxHCAid
kPeAagPuB5qlWw63UqX4jxWGBSnxUQcwKuXWegrcOnlfaAmgGAoDC/k4lmLT9cfW
pygMXymAzPIGd+1keubBKAXnejcBjv3w5aOggUmW+sLaIHfYguRcjkWcfsP1ppsr
TC0gWnSbU3cFx8aUnUpt2BK2W2jyYWab2gkQlTdvWZNOsUj/3Aw6UYqFB0Azg7uN
IPaL5kI+1gmvLN0oost10zyUGoItT0ZCX+Eg624ho2XgTkH/SbWpp3sxCvtqYLAW
U2C/fcyt4Cua4af5+CjbPLslDQ4alh7QKm8KE+9BMrBVLVPv3CVAlnBSq0r2E/Xi
EWrwpN5j5yJfkGFZv64xlGbqVlpQQegj8QZSPqKTK12o22Txs+kCNjtNtHHMP7ee
AaPHpsjRS+R1pmm+w6XBIirPTJbNai84GlHU1+Fakvkbwp7gnO7WEXS1tYGWbFQu
1MzXNxCJ298BYRIX7u6uWFPl7A8yKhOsHF7fIz41VVczO1VJ//1JqwbPXxuJUqya
mDWPXRZNTOdID2xsb92sFhpouI2bgJz/6isxGF9Z5myTxrRVRU8HLI68QApVWyEb
nlV2GjTA7WTprhhyF64rmaratiHIZI+vUW1lLK882PJ/tdxCoGBBcMQKO1Mddokp
Zi9T5Q7kOpmasbcyQORl5kpm6ZBjV1hqYSHmO4rESuRWLql8/YjbBDmAE6xmSk9A
Sx+fVaIED/yVCLGwvixTN3KMHPneCZORhf5OZweLC5cC4m2+79HsWX1xGDLR6Ncv
YMHdA5KrSuCeLF5Ci6dPYvm0Wj9YxLV7peQKCRC4wsxh1UWUck9Fg8dyHLcEJnG4
s6s+s883W+2EkBIc8c9a04QykAsAlhHoVGHcfQ2G47pRueqES+qhqhRQuD9hiP2Q
8kHD04z3eumEjcPS+TnK2GYKBJ1Fq8lsDfFm6X/Iq7bL4eS8SOcBJGUbuEmXfG5C
ic0jdlCs7ml18odu9PbnLYP+XcDAzyCBfStoHClCmfbeu7rJuQXAg1FWl4qLyqC6
hIs7UZ5bCNBfbKgEt0RIxxKYp6ObXEZhEQRMiqmbRMkNltp6kT7Rmpl3Ejzjp+fF
lJ5F0TrCqWdXNE+2QXUsVtn0f3lVSWMFvmP/i4kmYNIrAcs0cPU3S3AebHzoCt7k
svbPiU4G2xJnFLJkLkmnfgNRtFB4r4b69K4w3YNckkHczJCwZH41rCPxqVHLONRB
MhKp7LC9EkZIBz1m3R+yM/syu8VUtzpMJ8623oyZqvbiximV0nCKxB1zkTHSMEEM
BxiPN2JJpSTPqqnJoImT4uthO8xyGcUkO8Jp14+wmXZfhYWo/IEkeo7FxVCMc0j/
eQqPKyrfXzlpF0ulmiM2lM2mTmLDPbeGcg2wvloniufEkhZ74jfjM6u1zl2/3Tfu
hmTjEtjQMZA1gLpsqsy50noURXuTHeI59qucKCSPQB5myTrEqN4jjRSx8LJgQ2Ht
bc2x++/T1p3CPD9bgqa3fuY5r923R7mHdK0W3/BFbmncqJ3qD1g5H5pT2CfSu5j7
6OsyEti+13hKCQQ6ol30najxY4E3gzFfAOgCCWS0hvOpIxBvouzwyN1el2dWkjIm
bPu58Nvxmo3j7pOkxUJBTTy81v1qJhTTPi1H5aRgw6MnEOxCOyG8TKxUYg2ovFkM
LO844w66rLUUyS3wVk5FsrhKdYEHnxEt2CblCgd4cjUcg5vt/DJyQKfRxF1FtEpw
bnqNwNeiztfjvFWFvjO68Ci/L/Mg40Xrcgn3B10E1ScxZtUbr4iZ1in5PTvo/tWY
EUBkvAQKNn1sswAHuKzV7+mFh0QodSg0pwPUXb9o7rff0HHxzrOUXLcmmA1jfNg2
mvY2DMIYcCbwmAPw9yn387mqErXcLgmPru1BIKYeS8I/JEDpfpQLKaI0iapOD/ee
Nh6W7o5dYx+0LWDXQLfig7at+bXJ6njuudTRwfk4zxasCavuC+rUQDFtm14xkd3h
d3RCmn5RdphHSecwKlOOme2SYbkr4l6lTacYyg7HVlxZE2omgqdOHu/2RQX27+Ze
cS0I3NWbBRM+6+qRj7v92RZVtgkEn24tkjsbs2VZqbDrlpQckgNf+F5m261uDVEb
zpIGXyiRpBYCo0B9X/Z7qQkcPLwEGT0RrZ42abPbqHHEmlATZ4tay3fQA28KF5YB
MvtZ4JI6C59qSxR0aDLYzPqjXZeO+3hhfR5mmw3UlHYm4uTpD97RUSP01jZ5DWVu
h5uHg/W43wzbE/aoJ6Kj1ju3KazfsBFTvQI1fl2c+As84XDGz1bFI2DjZH0LkoeC
GMbTveJgJ9zF6za4YNRZzbTTtvYCvZbqOGzeV8apJ0KjNOXlsGcKIk+lCzMnEENs
ZIproqGU/zDoZsnHBkKgZotcTy8/fcTfvYm4oOtaH24Rm1B6mlMUKzgk2sfPUI0g
K33HnDN7z5w6zZpelKOzRcimiObsaubo2zqYaC9kO6nWXdGr/iwYdWg4C2n1k4Fs
W9uAuz0nrpyx3bfY+u2cw3l1iqn0+3RkmZ8VOxiMo5GmkfdX22yQ771n7a7U/9kj
/itVunE6bJOD3hlHQA7P6stGsKPmbrPZsrxKQfaKNx3asq5tXs6me6KPOw6WIlF7
HGcDxZqpv7lqH/dEz2ZLYhJBCQuqTIOrzRf87hwQeGKT9FCBWS24qGjngXKuuQT8
sJH2fPyLVk47+V5Q9CwqKE5TcmuaF5dc02Ucu2c92d3MrBlPXfTBNzIJB0boUYlv
+Eu3fgVkccQGYBRVpKloqExnJlPfCrRrV9W64D43k1ujMvJo06GtsQm3jWULW7iR
XT+cOornF2KyXpMSrqtgURcfOuxSeqEhb5w/4k1Gqicop9Gp5wtbPyae+h78rmN2
cO1mUpoqfLG0XTYRr7ZfKJKbYuAsatIHiNw6f6gCHd9a70pDcu3X9WxrEINOZmr6
QcFmw4puH057437QvLv1loUeuuhPTOx9UVzJLtrLfGIoIhGySxZ7GbT0gE9da3yE
5WxDanY4Ysy4ND8TP6XmY/R4OMLlbF88UpFfcSO1cda9e3xzWo3SQYuksuc69ibS
vaelwSMP1JPbgafMPpC7N69tvHjICmJiw3oTR/piCDF7x0oRXL1xCpjaAOcz1pVA
/H0OZxhTXjpiH4PoS/5TLYSn+0deNc0czpaSWV3n/d4B06quNhBbxxtNLpgsoz7c
IFFU7D8uU9VZ+NH83sGAZaTaVsF17kT9nAqJwAjVn+B/2zU9T4PsdDv7F3MZEkqn
S3S07IyyUvZhrzo7cyXTkj4huvxg8LkZFPJ5/GqwOryYY4jTdNJ99nZEqREd7qGR
oU+2UWPNB+vSo1DQs4iVISEucIT2KidMmbVy8lFThq8Y6l9EKuWuRAYizDakv0lp
4fMx+D7qq0DzJaYy1A9Di14C01RUu5RfCSoOfOf8kerus0uhfdz1IFH0qjj/tt7K
KvEHUVBKpMSRGyDifTU9SJmGZTjuTnuSujOj06988SdSlTbrNeLrBIIysIsPPtfH
zToEcKU3k1Cn9U1r9EwS/3a/Ic9jlGvj69SIvJUyu/zyXT5jFQTHn/c5TfF78WcH
R3Zh6LqHArkbbMcIAdzItuIut4D5GoOMLM4R3Yz9RFkPoQuOsrQWgefWgcAWJCJN
DX+UKUxwbLJq4d3LVbHbTvJ7/YdtMEcP+MiXRm+DSAYd4Jq9Md6NDcz5Aqawl6WT
CEe69hLc2KaWat3JIT+JcAkzXnbrsPfYopLR4YdRoLTnl39/dnZauv3gvnaNniS+
4hMQkNvs2H1AFtgggcLCNTCnzh9UZsG9YPDXKlPKVJYzmEqbHdiYlqJ7amOXnUkn
7ghEdmoguRlnWp28xTlo1Q5qvghrL3XgYfbJ+k8aIB3/YGcziXhtCrePWwaO/87o
oHejTGh9QhcAq6lhS/jCKiC1yhSUrF6TQPfGtRFmMEZ2FjlYvsPIR3GdohHTBMmY
94l0o088Yj13teEB6QW+zsg2L4uWpKH5rbnSt9h/VQ9YTUZbbdOkRNS6ULvmRvM/
d05jrdxlPPFXcNg2v7J1IDQQxxWxEoCAc+A8usjgdwZpo+gufWpQK0caYDdndESJ
/L0lFuY1OVtvT/ALi+vu1ivdu8NiY27xPfPG3DbdirRFzByF1ALuhay10lwSbMpe
XRbAiyNyn6ijzLofhqgdDc5F6SgoYbU7ohWSrZirYOuxLgb/YlThy11i7bVFM5RT
Rx1VphQojUdmatKRPlWhs6p8JPMzkOchJ6rnqol0yqGp7OpWyBsgmDpx7OAyt3o+
YT4O27mDIGr1HF4Ff22h06280CmKvjxVdW61mo9z/aH2f0+k1zF5ot0hZ9K6AWpf
e7t1Mwhjq3TMjBlNWK/l0mIYzCNDvrBW8AD65nYeU4y+3rjFJaoxFR5uCyYAcHet
Zk3khS9dW8TNspHI88GZVVkxV4RmGCayJsSEJQxn48UlvzO3esQVqEB8Dm41R7cc
vUIBxzKLHzGNpf4TYtusjwcjMH4a/oWvqIImV9ZIqOSrby6OjuicXwxPGs/sFgkA
LrUC+6064XJb+NhD7IsiTxR/TYIf2Q9GdYdA5IM/iL4nfvBKYpDXtv5qo/QWMqdL
zCugZTP1/JhnJfmwdXAhaDxgNDE90dLSgqua4T+X05SLtGzot4Deb2TgbM9G5KZO
/3oyLmEaxnRwkmoFQ+5GX+ZFd/6t/ZPDGD5r4PoGj8fPM2jB25zY3UnwmjQAToD3
C3jOem+epkmgJpmEOfuHTKJ3dqRZsclCUF8h12Ymcv4bg7f933PR/6yh2MN5buZG
DJdO+nvf1kuYrS6HEOvrNcppg4J/IiNTD9Y8bOxbSdFFhiW7jVqgLcGkY9n4AaQ4
P1NUrqZMNtc2HBD9GpR3aBLD8uss2gxTdl4oxTriwLEABq1lWk/RARCzyGSd+vm+
b9XEJDgkl9BteFcUoCuoDbyRjNvgVG+NSifrQuln1ZK0lAAFZvwD6V3lP11VD2Xd
6JXmoGnCGlui+nqJsRjspP+5Z8F/6Dtg83QIdZUNiXGhsuf6fPW9qm8aaCcXzVq0
wq1kQzuJaRRVdHpienB5m7CAYxMxd5z0YCZDLVWClVglMQvME7jn3M7RCXPIsKcg
qixRkMnbJ/bN+vTtPPNzPJaswCC1vcO4ARIn8YRIjMayVmMGBDibd8ZLhW0H23Tp
OyRBLPT1rSHURzR9g50DG5KHH+MLCbrFNiLNlRZGkgQY5YRC736ej00sc7QMrbvX
y00/3eu1C7CGgzxSKPlSyRTSAVe7oubcaIanPqaenV4XJvIo0J+qg0gey63sElTm
H8J8Jz5uExTNiKmNGersiTr9s4fnPARINvsO9KINOY25LxAU4QEJAbqYSqC5uniR
dTteWNW3q6wCqV6QfeARzqfMja9BulcR8Zd8nKIGHhqs5fg+oBRbiBcVPdmT7x8G
RmQuRxr6LNw7yPrR4ALo7Cvk6mHWRXeEvfRjVJxquef/Z752S9qvL/coWShNYTfy
z0eJwtZYEV2Jt6dqEwBIxq84eocKYQDhM4XhLT4rvNPOJgrinuXB+QWPNfc4WJCA
G1IQIa2TPdbMrexHxZPVtDxOlJJEfgxEbseAjcTIPQ6G0byfwTAeTkZ+wgY99osV
XntTwQV5zwmOTsSftiSGmcBNVs3CpuhVfSz94lfKwtrJWpqwea1ZsA8AXUkDsNzR
pr45bIkb6mszivhWgqEgWLMz90DK9vk4FGwbzVYbCEWFkvE3JnJV3aNcjU8MiCON
m3r2LgenzbSGcHNhSVjBn/7w53QJYsSySLTJAI0hnMRSTtvcYs5GDkPUrAhtHAd5
nXO5nnxK2CyKslds/ERpsQb2CaNUFQlP4skuhND5fz7j0BCkas8TFPOhxw6l+yQF
s237qXWD/2RZ07w78gmvyQiovCt5mzBqF2qgEywMzsgBR3R1h9WhTH4aVOyIRuob
dn4sUyOJ3zc55BL1hD6floXhOhGnLaN0mBJTDk7mqQq+RPUNXnL25WOgb+jEfpO2
4+lICw1G/TnlNKNeYWoaCNgxCgNf3J+lp7UtQmJK2zxH1xhdHoJDJocbuHaFb13d
NJu+VA5vZEZ3c+o/+osaMnSB8CKmMVEWc7cTDOfZpIK61ImuKufBzltATDdlJAzc
E4nDvlxyP2O1Q7FFHU0AdnXV2HOmapad7MR1zc4cwKU6JFmebXITEhHuf8fOJ3OZ
6aoK+0z+qQBqtj81gBt8MfxFWDH06cRaOhbPM8eG2FynzXjL+tR1VFWuP9yysvYN
ovwzU1ul0ZBrpQxksCil1ZeGenr32rhhyZkkn3LRku+xTiDzjb5V42y29gysw04e
Z6zoMoOvW8wLFr0jQBYRzf9StEA+xTlxE/hiaUO5Bse9OX2rXQQKPh4K/N9YrlhQ
py6LevUfo7Dz/cyIP/8nNAo4Pm+NRuYhk1EvpXjTd9qEfuKAga2Yl/wzxHu7wonE
o/+xrc8FRScT9YnnOaClMhRtGigrax1ys6XIA6SFTsuSxKiYiWts1EJtnD3NRRGT
AsatGyfb0aepo3cnGtuzqlPln+OhW4zl/p5Jyq8YjeFZTJWyyX2f8rdTGuvjwf7l
DDVb+4ETRsvzSsyd6dAznWo2lEXgtkvh5ObFnaDOMO7JJ255YFUUK5Yfv70edoxl
xOMW1dPFSmPiKd8wu/1jMM9BuxskYME4M0I4fJ5aCmyucGumWa5zQ0kLvJ7ZSRGD
Vyo7LyH/cUjC+wpiJXqsMryPkCUUaSPPavcfqNKGs+NjOaz38yt9Jmbc3rvnXmqw
Gzr8vhQBwHSm6xzzgfqKUYOdZJP7eo8kRo9lvujzAPKBm2m6gXCy9FlvYkoONPbi
mupS/Te97RPXBJeYKyR8BKrj2IdvVlHDFek/Luup+DiMn84crtG0frCx1i+wBqup
AVEjA+7bfyrO2XuivKzLcdIyz/wyi3BPu1z1o9KGBBelTkJqDLRAjbweY5BJeCW7
HF4rEZ/l/SBFMXmpcC46yT4Qw3SKv3NnS+x3cHlhmvnBv9VdqxToOCmkAVMMEJxZ
Vkh+5c/acyJRKs4uynENYkKa6tRA2ipJlPBBPaFS8FZpJ+7smc0lg8mCTMhiwP2/
cwFAxllW3kf2lh38mhly5iqNckPseNAhduMlx8NVWWabPrfZ4WfDj6hxyUtDKztI
JSr4DTfbmAKmEsjXhCn+0BYp4dytS3k/HhBIH+qj7n5oGrm57FAUApcN1N/xvLJR
eLkdVH3pw7pvZRnDHr5aRQePnOY+N7MmVYUewO+LcdQUEa25ogswS6iw3QiD4Msc
jDYQSeAne2ZpU4ju6CbBuOC/aBvR3UeM0CVGUDRtuXoABxmc4fFRo5rItHIec7LT
CitPnhiXU0CWPgp44+tIxY1Yt1qnRP27ug089XScDQLVYG/j4mKq09kJ3skm3SNs
YuyQt6GM4wcOipGj6GA+9pMQGYaeG6c9nLwRtAD5FeN7wRlgkfos5qEWisWBvnZQ
u+B5XeF5FWB8M8w0rSn1IdozOj0Kovv1dGpXRWDL5d3H41IPeNffeaW9yqhAiPrT
bHFmb8EYBgX8VuNMlXXJSHWx0sI6eMH0dvjAaT/joiDXovbzBkVLBPds8tjnMr19
m6W6tWYwa1njoSEhlu0AxzRHTo2XG4Gsn7x9ARBDAA4847mNKDcs5C9L3JR7rP1g
L+domWsVQLWvpQfe9jbeUlMoVJYY7x3zn4u6hyevJLcenPXdo/rTJhazidBshawF
rRDldfRqciP+XFubBQZzAEECkzBePFMYOW1zKM+IX9tV4j4NQ6pttPhdmlp8mHDO
GMzCG5y+QDhGsYhaYe4rYGWUVJ2HQSeSNSK2ovSl/0+P+wWgoCZeniYka9ipxDWt
Ah6XY7YJyJIDLh0Cdx/dg5yK1xlDLXZ+E1GLzoIKDdWB7DTlyuHOUm1CzGNlOP9Q
1N3xb2xPaSe2TTFtu8m/X1XmuqzpzzrkS8WihXz34jq/FTkkMQuJq1u6SMuDgWcP
tdU2okGpDwoBoSgNu6+vVgbHvNRfcAb/E39iDq3xLInvhGlLPiBNhpcTg+jCq2GF
VILh1+qs59UipqKIHVrTnU2E/mwDuKCj6MvvVIg81g+7SO2CjL1QkONY9U+qJLpy
OANBZy7/xVnRRxOnLFu8idhV0cyLJdorw3rZQayr9Q34MaZEtTXB+x8VxFhcarss
gOVi5f+v8OnwDVhWFVJIDBAJBYl78YVEJg9v+NHIYe31NRU392jBZ4hn96WoIUEp
JHzm141W1Dy0cZNFVLb99oRZVirHn1Ev1GUzfvZYnZrTSrdAkh98S9Bjxp03QWyu
VFvkVHHzvr1AMEVCh+fOx0En8MSbZAyLlV7ZgEDXU4K1RWqs1LxicZ+APqtAWp6C
MmtoZ8E8/Ujm8zJpwCwPxKC7dqHDBddQ2Ue3R/DYZejhrLJGWO9aKICx4RMcS0Hk
xkvUwq5VJQBKVQVB+JCp98Wi7sw+5HQolOuUXvCP/IhkW2VgzlP8C2VxaNcSJP0c
jHChUk1qGpt5YN61VC+V9Ex2d7Njc9kw/0Az9Q9zMoyB31grRk4R7d5qXI514PvM
i8A7aj3fo+m/v0K+ITc8ie/NJ7woldlM+iJhk9G6Y+9MZ2u1Hh0XfrXdnRb1hqCb
6Fr6XGvx7tPglaHQeX9hwmyxY7nZO2yFGdIBFL/YERLjBvOX8ochHtF51PR+mMYO
ucMytycYdDGNivoB6nuRBlP/cybkTMY79J0u6JeujHfEOR3XwZQ6pF1Bi3OtpYHa
BXKbToY2duQIv6S7AHeU/Tj7jL4cDjbvIQQfq9Gof4TokwxM+oLmvjC94fnaSl7A
Pdp/HxiO8w5VngESEruGEHl+wwZD93cD/OWCAdXaWzjWL4Tzr/VS3dPLmRYvsYbV
YIWRTQoLjRImQKBSZ7dir+0RSa6se4HUQfuxALRNiJKuxCFSgSbJNWMvqFBG+9fO
1s9VkURMTY1zrwbLK2P9rUtDcMVd6BpJj5fLX4gB3rrEK+GxMXlYqrYY6RlmFh4y
4cnJPDypv9bRdWAH0ucmjIzVo0b1ceW/jMBa2NagpCPbexP4QFxOa80uachMVpF9
Gh7rohIXjuQYX1KBvzd3Jwozk6r+YVvpXhBnrN5FkkIbYQQULUWST3NzVqFRPbjl
i92UYgjBxPKRIVg5qtgXVHWtAyY2DMbRGtFBw+BMLfcZG3YU00SqymlrYCYBMbUK
VTh43KSe+GMYZNYrLshEMOTWdvieK41TVSmpUusyQtzlmaYi9k5a5HNDvcSHqWH/
Zg/6dUZ5TAKUdpimG4zbGab8hTECnsUQNt7gPS9fYW0hDoIAjjt42fpUHF0FCR86
P1U9WBKE5Rr/mpwQh3j801ellXvDkHRIjiNEh3tQ/dCSvMrCH4UAKU3KGfDR4Mso
BMKiIXZT6myiDdGfhi6JqeHw4CNYL0fexvQI5Al9qGmxdgQjZHehkV1ZHFg4TVA5
k5ndKli8OMy2PkhYAm+E0mXFvdCAZGviHPuYXOY0igC3sY50gUE0/tbUtVZ8IxZq
554rme/QtDjJ8WRBvdTqa8NStOcdnZZn/PYVaoRbx1/3ejcGHU6jZXMr90bhMv4x
QVy9WReN6AJltBuXvZEmxpphyv/6tYxMo4msK3hvWp/10hgEuChjzL9zUN3QQ5Qh
/EsaMfjbv5fsRKk+XfiF7w0igFF63VN5sKixExfCev82EoeMu3pIZYYw4U39fcBi
Z1fXfN6iHLvJR2BQpAhQSzWJE6fJwJabAQ7s4dtQA+rw8/5ARpyGObu8Ur8b0z1y
HQDposukYHxayDyIpPmBCqUjfhsQ+gMkG69VJKlBxOAb+3C9A/CNhaAQj3tqulMX
7mRsz1083jRvr3x7jfGQUQDc2eXrRu21GUNqaV1V0OCHStULSV7rkqGehI20nvbR
s8HmDnWCdnvsTk5U+3lOQr4UljoYqwq2HNXgfinncR7TNx+yOR1+XOSgYHUKVjDb
1xzt2AwOfkMAFMf0BudqXYcNO/1JY2kM1aSlWOuHCuT02jhaEQQVF0/nAPUTdhm4
/o6mXMLWqLLC2uAvU9rcavszhJkygfXjn4I6qryKtfsoliSnVQEsh92Q9MOntptD
wg4ChhgPpvlc29YxnuTNPC7X4seBGpCjGcZWu02FPoHB3U8IoCPLGS2fkJJSPMFc
WzuNC21wauQ0vx17K1ZrqLWZ9U9jAlT664jggyXjTxDxRUEFEzwZ0k6k8M0GvNhn
+oQLr8LOSS1LfnFiPp4kYKj+Qp8KEjE4BD4f68oc+3heY1s34k7c6higOlJrXomA
/CJuW8HAgjI8Qr4ffQBQKls9LAz7uE4KhQmxA/vocxBOVcLnkETKz3PAamjWM4qf
JYhNFJcQHmdNO1apFm6U6r/O5gkf2SMnOOZJE0MdN875eJYAi9PDK/vFh45AXSKn
vK+nwq1IvP8vu8jZ/yTelaVXXi1kM+Q5kf7OoF89n7UoREEkHvFOCpZ/5rxZvhVH
Q8NVm4BZ9iGtxiXp41HMd/57txKoOoqlNzwABTA0rVx74KF2Lcc0xelikXdND8L+
cZ1wc4gKz9UUjt/2A/eWIRS5xSlwffAcOQiRvMGBdI5YmiSjsNghhdWgQ7l3HCn8
HnLe4JvhT4BvUjRL4D6a3UjoT3JVW4R8974nnt9np7sw1kQMO9c5fMRAvqGwFN+T
GyGCB5cxr9QtttWSKcQaY2xYnEuf+JOa4BbTmJTDUCxvvSXjKcHy9DT32RgQb76f
aGsKer4n//noH5Kr+SbJohrhO/48mvTBT67ugI+FDXbab4w6ZxwlY+8J1lqZIrVU
0CbbVBZOgSTOo7UCRlPdK7eVfAHtmZ8EptAg0mQphGJVn9t5dsdzpMYc3sgNMG6Z
cDU3JSt96mxQo/U7sMO7xOOHt4OWzYKHVOWZZqjeboEpzgndC3/Yt5sdKLZ82fkp
LFwrLf/eyK4GneSv/Vb53UtedwTOWh6+eZFk57nqh7x17rf/I83P0GrFilhraGya
6T9GRTVwZ+fZFCMwy46liWss09vbiaXYFMHql5nD33gunUC1psTdU8Smz0P0G8Z5
jaRDCbSnnmpwfjb0zdEFI6JcxkdkGVRrdOgn2rVnDkLsGnlIO9eIX2y+MAeoy1sB
F0iv1SX3LnmUnqhXjnuJKFv4GvUEgOV0+JGgkKx5NznfRV1c3QXQIHglOROX8EqN
+4X0KGDgrIRTL5bLFSaSuNJjwYz48W06FmeoedTsD9NqsdbSX+97H6z4qtQz8kfJ
oLIFmrVnoRetapfax/4H4Ql5yCaQcwcC7fq07KCqO+JKBPJXqPCVicFjh1o+LHjj
nPK80sQi3sfWxWM3vDxYqGkJA6N9HmDN8oAhTjKd0g1LkP9Jyi4vMfKETvwnw5NW
FkEDJl6+3W8VFsXXSF3iZDH4sSSeZOP8cNNjDqkD9DEfNrB+A2cAGI9CSqhFcWoK
fOzSEaBBpm9uZrOi8JZw1D7/BTf+mZg6JPMvB+Me2ahAEXtVkIahkGZwut+StSwv
rjtrO+3F2BXWDOt2O47+eWwTKb+jZT0D5QEC7sbbB2MNAHva+VUBSXRXm6Pf9/KI
HzyKXkqRe4lmHhz3LMFM/hVNFrTcC+iv90O1t5vIkLXayKSs1XSkhQaaFnwP4Ali
JnEtH9xOwt81VOlIk/VEUOnpUHGCte//t1P4zbSXFeJa5RBylo2gU02UhBYAqBGE
1d50YP1kbnPyTvDlG67rvwuqBOe6qsXFZcAhrc612+YO1xgvYVG4q+BMdZVgdbGf
2saHNGr93YBr+aQZUPPXmD1sUnx6Ma73lMEm36pRnWhOl2lIIoHCbA4oTRfcMzxJ
D10Z9HDtdXiVjNkWbFSfjGLvBMG0RaTL+L0ihFyvybHx3KRjtAO8C/tCTLn8PQsd
IosWGLOJY18zHnTk26vkTlmUaR0wB3Yajk2ADR3T4r/uIYOLhKq/nB/YpCGNoh5A
Liy2mXR+xlzpbiMhry60j+QGtTXGbYqDU28Hqc644qmJE0HKPH9nHt6aq9Mzny3o
f2qNGqrgVmfXCYrHnDzdFR1xpQdVx/s/CHD3xT8TaXCmtmo56x7sblitf3wMsP8X
6NFOGChr5di4oGSLifL03JuaFJm4xX/fsnLtPJuTywJmZKObsjRG1dtdj6iW5lss
4Cax5/Uyn/0rmWnxpVGoUzFhIQiDh60xd7rYlvd8ZLZ4RC77S2IeRhRXWRt9W5SZ
0Z2Psv99hB06ZARJd6c1vaROWvVdR3Xa7LapEI2WRp4CV94I/hjjtiZGCEVrP4BC
fq6ta2Cff5fzj38pOowcEY94ttBv6RIVbDZGMDetdiPA3Wiyv/bZuGGJ0xMJmfHn
qTJZ4HQBKpa/NPnwMJd1TSrrLNhJSTs/97lryti4Ut5c6RAONQnpBd3a5APOweVc
EPnEGVIgZw59H/w1X5r0fZoNKBJJE4UDv2i7quYSqboTKWwIPif1SjByZOAVvpt4
ao6QUANlSpL7Q+aCBDff0OsRIgJMbsZ1CLnmdOAgI7mfFoRPaY2aeVq3gEmN+gmr
z2w+ycLuQ9ZmtAndQ3+2iIUO7y0ydP70IN6YJAWR7iJ9Iuxzcy4avYcrMAuHbg4U
Qfr18P7yrl5EOGl2NZf2nigzOSYaw/iyswuETcToGoBiVi59A26A0DWLvc7DqgAK
ZhB7Ghs58HTV/ZxZNhe6hdrOjGvQWbACIsziHCB7IF8rzsj0q/I78gHptyE3ahs+
HyjJZOLyBgkZfHFbcXB+pysyOYatNu2Y2S1xU5KaB7/JiFsnUdKyhnLXzO3QRIKz
ccZ69EWym5GCoOVj+eVRCVK9BfZBfk5CmI/iyXeqL3oaj76zqFzPEW6UD6eS6Nyr
hDATfCn1tTp0ez6ZpuzLT3Lg5RxwXecV3RTndHhWIM0OgR/98EI/Zv/iKrsst06u
gvZ/BM/KOIbPAI27EIuS2z4onNYScMlSKXOPRDJw+a6oepFdMqyrZSeUz9FeFhxa
a/g4bn1zXLmT3jPRqwv2/TqMsaVD0GaKV2KCN2sy+a65JvW1L3+98lkaYHRc37pn
X68eCpqUOtvY97/ayYF5qXK+kkpzNUCVBVHpeNNz9J0h0Dia9Uog3GHAkjMFjQIK
BnnVp7PQEbmoqiR+67TIDLWNVH2Jxg6uUY1wsGA76M4GW8NH0tj9hRrGdqvWGMaM
ibjd4SDp7pShBIYbOC04D6vQa4XISga+zFpADWd9j14j8fRoFV1nkuJuJtnwOb4b
1PvVobDHU4KZGNDLlQkSwNSeN7QNGUsruaydGd960FU=
`pragma protect end_protected

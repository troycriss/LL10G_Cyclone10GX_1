`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
XBCnSHgXtS+sNi+Y71YQVAZOQ9Uf9HBwzn4djcDf1aKrsjyErzCB5KCtyJICHLNx
7oGB+xU0/EyzEICjs5G7zG/hm0JYPGsVh9Q/7i5itgOU2afj65P+3su+Nc+XHB30
wnGKM3X9oj9DyrZTtzu365TSUPtMsSC9CKzhe9GySYU=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 9088), data_block
8VM7nMOJ6hBX1Gdvvq7t6HjprTEc3d64H58wQ4vIZjn8XIufeeTiYy9kNu/7CBQ1
Baj5R/fAXAvZSwUwtsNS40KhHxytpH97MyxvEAOruPq1F3HlLNIs359vyjF7ZioT
u0lHkNT2eEpfpV8KKpIbwxqzvOvqISSawANsOGVxImmHw7+Jmo/4lElK5XRxwWG3
xSEbVrIusr8wjRc4LPoIdkQUid0UmUKEb9ciGEzvfPIbH2oIh8zFOwg2CBygoT7m
SlUnqWuXegXvSwgcceZh2s880zO8WtUeiQnBpGKPTFTnSBJhQCacuMWMVsY0ZU/S
Nm3FANzfAIuhd/tQLCRicZR5MPad7YQSAQlJVMeUROJG5ihJTWD3X6LHF+NiibHC
v1ned6JjdroEsomiKWEQesVRczH3yby2O/fu/JFNjH/5huYBHIiB9s9pDoc5LiJ0
fhQcbpJLPyr0lgQ7dWlEtkWvTBU7ohu4SKnKvrcq5T6f3lCcxeNFPovTvnNnrjT6
M5v+jiplGZTZTRZJJKCVZ12ut/iIucskkHrsncYsuunEecWPXlZPrVbbE0+PwbgJ
POXXfGHkgYkYc6tI29Rb6eyrBCcnqiJZfiZIAQQOXMybmKFLb8ZqJGFmL7MrUPjU
DR7YZ5yDU2VS4rVn4EO6yTrxZnhfEjPwQ9e2NIDF7YirCm8j+wXdCh4qL3QcE4IV
Uqx/FI7grBDLPkqD+rKU5XKuOshTR8vyBbvrDQ17frJQAPlnThQtOK5bAsJuygr6
lq4lYOIdez9HPK731RGLEZkCwFiszzyDM08KQMfM3ZYuRpyy+8ZZkdVFVzpthCut
0Qc29sDoKajIcp6Qa4IsxLEvTv8x9d3uxOaygeGOOL9/XZzGKuXUk0RlqCjHnw1U
MdJLTSg6+SsnpPqp89WuDeb7CTYbgjdn00yz3tA+bfJdYqUzMgw8XraF6K2/IyzV
nkaf+I4knU3hgTJ4ohSujQwrUbSCmq8OqpzMgqyCvQvZn4o0684Fs3JD6mb1a1WL
fKvybGfnW3ZYxedsE5WYqwnm7JyNAB/veJ0HjcRqKIhv7kCyqdeVEXmKpEK0xVVh
oNpTVklIJO+/TF9vM5Z0LJGhmM1e4l71EHZCazwJZnW6cZvYhr5JGGvjyZJv9bbk
JtXP2yVKp7dkM9nQi9aHOxxdXMh4Yc7yeC2holUDu/s5pj7ssHdQc9ZX3dNmerMX
FHPB2O2ID3OGAEVUlTYhKgUOmKB95PRuWrDvnDQBw73P1oyTw6jLyiicbO3v1/YI
WfqFIF5Sy0C99q4gk8IMG9Kpypw4BRE07RycWsw3ukR1xSdJmGOZAm60hr3h2cYs
502+OkLTZTem/gV6YF/sBqcD7ID2ddgeGZIXCm6Ln8YRftiEzHVDh2x3Eope+3qt
VZ3JZ1xTRvBSB1qTs6FVh4B2hoTZdb1g4SeXRwMEhgJVwj32BhCPMB7GYagGxuFt
Spc7eA8LP9oRz1j8cGT4jDzY5T0Pd5LJ84Tlk/WibnaEACdOyzrRzXuEKFM4iMml
i6E9n6an+5tvVqj8KEeIYwR8GZb1JbHz4mkeSOWyfmTRW//cU/4c+JS8c8SegNWA
VHz+zIlN9PF30XzTitygW9McZ3Q8QrgCxLEFeGRKOhkVaFAkCNvP4DE7WKIdbLK1
rXwGONFnTEC5Ezjrp1X/CHOK4CvLr5A1YZeusz4BdE2ZqukspHe+hBN2oQRKEakl
NF6+b6hlHtK5cXv0apAF+QmOoXiozZHA5LE3FDZ7ucu/uWll+fv+KjcX71SsQFLe
wm9OAwUZlOpCjtCAenTopkVuajAj25AFD4SLdBL7nSkd3H3LCKyCOw9oVl/Z39VU
qa835LEupGz/jgwn5gZes5yqanmXt/s3wMEzeeVKicc1SjxAYo6uPZx12OOBeF1i
XiByudnTxJVLZkQEiLH9718KlzxbKFN1zJMZvJHe9yJqlIzNFofodWz3Pbii/V1t
kdAmr6E77m+wGMKFoMMG2fF7NencqxGHdqkTmgOs7+m9hXCKev3g/DvHQT2JCIFv
Ke3WberRV2VV/NjaLiOP7YcrMH+zqVPQqMD1I5oDyf6qfPrBwLrOdUj5gNLH2kho
yKhb8Y5SHvz9FvEiOS/v6WCvYQjVHETbsZ3spGeMV70L5j8P3jYevQAxjRv6fbZ9
zeUjP1ys4MwqzVZ2cgf2f9GfgqYbUyVZicUlxRjDxIwMuDs4FHwbu211NI9kyfg5
Jdh2antaYESTSln2ME+a6IEX0YPcqq6+I04jNaDjovadq0S0bC0OAAh1QpyCE4fU
cC8PXMfbGXrQm3/0jdY0TahCn6SIpyY4bYGWGg1kWGTRXEr1rH1Al1eUUAAVANy6
cpg+xMt9SHHpveTbXU257aHTslyBRZg6eip6GID1j5IZF9+QIDClcnSszZws4vCS
X2unZSSjozG3lb9FcJHy5PuEA7Z3NsyxILb54vH1KRbc5p/GRQFTriAdcaT2KsT4
l9zwuKOJdb8ju3YXdGCFj7o+tdcB21phGshUXcDpeE4E/7KuSPOAoYo6NxhpSVcV
neHRtoF4TsMyhwAevnL5ntMjokZinnGvBfJp16hnSh8/zjv7RBwUOeU0Rq84sMSE
dJP2mWii/cstdf45AxBixSfU0vUGGBUEyaE62mn83FmeLf08e+UUexriF7TTh858
HvKAmsfR3mEpk0w65E67ppQz459SPpKfcR25NFQdyExtsapLTjTz20YMWt4t6u2F
M/T97EGcUlkQrM12qebJXOMCveCxT1ERlHMrtDLvRVZWMpkEo3Bjv0xLXmo6q4FY
m2B2cFKQJ9rjrJGAuLpJiezVYHQlQeYgtjjSPZaVrEC6z007IKmsYKVTb2y4o2Hg
g33z8hl+w+QgNQ714qP4a+PrbYPYIjtth3G3UouwaEc2ar3dOomEsoicef15wthU
mQ3nhQmhRx6coNi+XYbaM6OoirYGV4qt/R1jvSA8w3M6SP0NBwIPi8QjKZkjhaKb
raS/UBIyK2pBgd/yATcdLP6WE7QDEX+sl+yfSOMSLSC81RLsLNTtZ+G8yeoB10yx
BKWAExNIYfWK6qAIMmIhtaLl9g1V/DyTOky71NFnRMl1u5+4W9AlXiYu7bZOrBP5
qkOicl97z0iG5eq4HwSaoCtAtP2YEl4CoXbL7nPYm4Iwp+hRahcFALGAeN0Zv0cr
Bjl9f4HXeUmJsAyF4UQUSb1PSVoAmpOHZ5oeySt03ERnNOfwlVExidfcRPz8eaht
QDmpnVqOhsxE1ncaqszgCxYlzp+uHHUOjyCdB7ACvSNAUVpwAfmoSNoFw0srbnNK
Pbb/I24oWs60CQaQhHwv3O0cjpUH8V4d/YRrO7QcodMC0rI6o0o0uoS3GkwUf8R1
3Wypf424xpDMh0Uu5DYDpMwotemt65MnPtda/JWKQBY/rUo/pBTR0sAo2KvKCEqk
1GML/uSiI26kb++7gwXCx5ywZMmoo4A/wcUcNBAKt0y/Qky48VsJxUh9v8mCNdOE
2+EKF4mqI8+Rt0Oi0gwamqa21AnV5iWILzS86eVbefFLCMapSITLMvm2uFLMYPpO
9qrPeTJdMeRgW5o+B4nx/HUTlVZSrRxyWEVbjQRRLtO2jTP9+i2X9+OMFbIJfsaM
7l+NFRGT+Uksu0NGSwlVs8aYVNWYiPvwWCoqkQgs85tn8i1s8mI8lpruKzhwersV
ZwTCWlzAnxAfgxSDb/IKLJIcjf17GVcZizY/z9RZNkPiJ3CHjip13myrBpNfQbIo
Cn7iJA8Jns3OvdT5dziUW/386AttxuDonMnOM/09Q/9XUgHA1usQMe3XNJ5Ko4oP
eC5Xa3PTv6AEDvLxbz4Kfm6p21ZO9mIDeb7qvdJ4ERbo8CbfYYV1BlzPr8QyrAyl
4rE9WdL6xnDAXMTkPSREWtA9qhIpBfux+YreN3EiMnA0udN8ZPIovIGUw2TWXWEx
lcTW37VhGptEwGO6pr6vcmTMwiSQqA6PIwMyMD++cQgoNVpkrSdxJhBm3V8W8D/Y
OQ2+kmWBNQIXHogxsQLIa+Cz1c4sbzoc80IPqDmIVSKiyPzrszOsbyxq3Kr+PBJ0
/VngVshPEtbIluCcgGDh1h359ytKahMqAw2K1XJER8gAbiIr/T4J/U+tTd8HYHzg
izY0sv0VYBBMhb4ww6hvcZDWCH1ZhgvI2d9mKXZzkQiPwQocH0+eTX1i1D+stjOE
3Lkls1oFOujmySrrcxHE2Is3nYus6rXG7Nwz3/4HfRirPn1RRW3voElrCTL4FKSL
sTUvlOisnS418rJnmJY/+0tuB9+WXqe6czyMvU0unNYA7ANvXnesKF6z9A2DUJGU
Sl5KP0RE4FRNm37g8GYrC1TCgbPAdXco+jYjXyyUZKFgtH5x0ljGJc6ToEGr+3RX
xnk2HUDaXBoyteXqXsXVZVwFGb8/BvZLwjzDPOZ0k5ZFVXYo4h20C2fhNd+tKSaK
5gBFdibdLcfAopzDrmDaEkYYUlA2bBazLugKCHG9Z9qMgj8saPuAhLR7Oe8AgdDC
6xXO9Pu6cbYaykdqcL9DWV+QvBSfHlpfAcJyph8tZqERNO924lf5bwgHDv7IOsaE
L5ijO8AoJVI5sGLabfl5JIlOJmnAquysa6m33/eHKQTH6w+RAnk3ZyquiYxAu1s9
Zp/XRyxWqM+BlZeuTR2HSfQOp7vIF0ZgeDdI0JTx+7EIr4AGN3piI/SrvKgxQagt
KAg9W/xDdtPeOGCSbf6UwIqG/2wsNi2YK4zYvPMsezKl8eSlB7DZJED4xd2Fze49
ZYBSLecIqOI2xUjKIReYXw2nbyDDi6Ijc7ND4U2u4yALlsOWa6avmIXWYPg4S7oO
HLDZZi8m1AApDlfsUq75PHoP0Cr+caw76Dff+Uuz4YVev7YmveU49T4pMCW2c+op
sqRwBIyDj/uF1PhVk5kdKWh5Q6n4efiTRPv2lvZjEV1my1PwRybSLnuaBURrCSiU
ngnrbmdlgB25w3HZIj+ZchiZcQAsALxIN2XusEe5FXfCK/5YVp/vQxtLuMR6SQXA
ZpCAAy/egEZrD/ziOJG3nmCHOAeAc7S2PsH+5u4C2xopXOvkQ3gVAmxNhdHm2bOO
UVIr9Auz9nQciWd1X2bdyWunMUvDbpXIFEY8AKeuRnbJPh4kKfjlRBbZ7a6DKznl
Ei8N/diRuDNeRaPMflUd8SQozyFrdC3dXkip6cODthrD0mBs+7Dp8i0BePJaoAfW
kC+lkRNBPfTe4qGmjfvKQOgdxmQk2+Y7Nk6dLqDUY40Bz7J25Rl81mSjdr5R902D
5dE4UbFq20P1g1eEBAZNZr+c75y2Aj/J3RCp04mSvROcURBZYx8DENbN1C7Q16qi
V44PANtvUHq0z/X2licfMr1ibBnk4u7PflAZB4ildrZpjSLsg5irwFQDyoyg/wsM
Z5ytcT0WBdQXR61tZluS+2H7dXrYVgsHfhfN+0cw3ocRVm9vDJf6iyJ1eGXIKNGF
FJNCloOZjaA9y/XCIIJ6fKjXIMeQK5o2dh4J84Khd1RdPqsm2BgiR8uSD1whEcqp
8K+1eaCUWUCdxNH+/V0tfX8NYTyOSmH9d6Qp6AfVOtwBGq+vWDp/waiRHlv0HnxC
OSPbXlG1wA21QmTNsXsFMnaISr+XV0dsPeXMpwuGZbdKgpOtY5zGMy9+huXwiIhu
fxHfgIkiHr/jJtQAHz2HPu2l1t4IvPv2yia/VWBX1QzeZhzGNGkD4d1ogJ9wKi6u
B36oQsLpKXbLhl5DylS+DPZ/wOFds3zgD9lS8BaVNFMeGfdoZS5ui2kxlso3O46F
m5Lp3vzgezT7xrdcAp/gsi4lmrVeVm6cL+Lqin8ML0IRmWVGx90czUbHJVm7+Joy
TIu5kUbfzp75PEmJUK9rFiud4k1MuZk4hL2zcZe3X2WCFVO08BnzSwb1canNeHIo
Oaqqx9ChBsTEQYfaesM8t6LYSYKbPVhmCgNGIB9F/solXGtmhvvHg2tYaa5Oshj1
d6k5xUH+O87ncqC1iRGBnyap+w2M1Z+u+N+gJ3bUiF9nbjmOb9FftVn1IMF//hHu
1gCirwNsUqdpacouF5mlmAYhc3sXEsNFpqAGtLDcaL1B35MlFa6pgTDlWe5uKQsw
ktHOSZw5Wx73b5/eswmVnfCf2I8rBIS8Tm31cZeG9mb6I3C7nXls/iju4DbuuVvN
abF9ghkYKJEeCTP4jrvI8tQrCKzi7k7AlEt4CyOGVJOxWl5moORhwtOQzhgKpsSJ
GzkbQpnaoTHTxWNkdxP+oiFhXhzjOlmps1KfYpUFDxBjFMbH6CwoD5/Hzsjg/G9i
GJsAzcMNVP2NO4g/K9813JXQlkv1yq1hH/W3oqoOifomFMKN6bmTBVzxUSxmbZIL
+sozpG+/biyZ/GSzsB1qI3xBzLUqLZJTYQJIchCze1bBoGASkuHCw8d+O7+tt74H
zY0/Ba4TykmeScXrfBcqFXW3FiT+buus6C6SofpiSFPGaYN+841sk3HEOwrAskUw
Foc1PAYrZzYCtlD86RUCT9Epq/j6mnjoHKI3JWxuXr4r/XYU1iwDnImeqV2MUcP/
5HQG9QGEXijZcfK5h8PyeyEyGWG9ZSI7NERVb/RJrGwaMYrFBeR3fJZ8TX9+DqK6
7xmlIER8GF1PXej4PyVCfFi+HDp9TnaBR/k07wU8cKGdgXx+Z9FtXMkXKCmm9ck+
aWvGf3+3w9KyC+AA01X1ZJ6fXWPnuz/TP7YQ9TWiMEeV0bAN2XsL9vGewS1j8D50
GjumttLxC0ivZP/U66A45w5CPSReoh9rfuuawoq+0ht1rDwtWFB6GO2t8X/CjHoW
feJSjpO3HaV2EEwLnN+HSQBm/mBYwJ8gJHaxpqhzld+5TLKu6g+83JlJKBuo0pB7
aNUmU13c//T7e4kmRo7xtVkwRG4ZFfVEwwPUWd0hdhlKeLmcNo3rl378dXsgEA0R
Hv0NNzf0HXEs9zYI0B+cdIf5wE1HrTyXwoOWdjSPSeHyN77cM3alMT91oQcmvIHh
FaiFemKFjvrJz3tBq+HYPG5H+xweMHs28lTXRJILc0EO+U83M8LY6eYHMtuQhicT
lzvzBhyVVHoX5h+qAPfpjzZdB9lXlmHFpCdbAhk1hItCYa+0Q2+ghSe8LfetUuMk
dqlzWgjfcFNTlTnTUM/lyDWhFDACtAsr3dC6ck/i6gqWZ72cQCjkcPAvDE4nnBIh
bMUOPQlWcNwTKQIkbnpGW3UmCwFtdQ8CdjnnG+d6AIY61CLbzfURjPWLIuQ0Ub0k
dMEezUl1OV4JtnqfzJBdev0TbPpOhfU3P22zKYKvzn2l+YWKWsYRCIYQrEze+96X
OqN9vB4zbiEVcFvR0hbfuNQgkXldU73QZglji6/25MParMsgOIJJF6CeP9ioLnPP
B6ArrMJJ3+TrTv5eMlLALYTIV/cFKexwBuGPKiw4OMUNeNvosYmdSgmoLy8Sxo4i
uQAfAKuK74s7K29PUaOK0lZROj1I/9tLF+OGxQ5WTE/ZqHxfgpBYVswrGOfwAN1O
rTHW18fNk2eKiyxYY1gwwYd5ntVfO3GYsz44gBdsjI0YSAi2YCnnv2alJyffGe7k
lYdnf47sLK5HckeCTICXgBOCrJaOBZONPWS5XvJdGd8CwCzVg1zx/IVb9+YqBRdv
TgLWHP4vjsdqB+pr3bUFw8CKFHEoMu8+dK5mGx0F4HG9yiBxQNXdAmGtwa0Z1Wyp
1cg/KKdN0W+835N78hOwgM2gxURC8KR2CmyQb1xthj5VfGjxxZYw1YDrlL0HzHcq
7YnKtLUIUS2t7xHuJJSYiiH0UUFh7a6XZjHKCIPfUf2Ik9i25l0QBSDMXdE/Z9bM
lWFhQueP3mjqMkZ37dSzJULH9pHElZOSz2n5Wg1W2ehkO9eOFzXo1w4bv2SKDjEq
alDNzWzW1WLjTd4WWa2+HPy3XtlAr7WlSd4CamTYCPj1ZyBiGbcqvF4M3p3/XvX5
qslcWxKmnb/6FhVEvALZ9JgYa9HK2ZR1g1p1F41gsVksJRHE2GQqHL9s0VKgknTw
T3yIus8XQlKYx31c0qiu3kSM8NKmuNCrrOVTBYhJKAa7BGyolB5owqE45eBZMSXY
KFEVfJ4OxXKz365MAufOD6P7BObmOUK6Cq4fnl5dmvMI/2pVzAz0iptqwsnN83Gb
Gau71aGeTXeoCgS3sP7Gc6+YhZKge4/6IYCKhnDgUvO8t7VXl8s2sVJq3MGtZu4R
71z3i/rn3jxIqFsXFZveXdRrn/YLAsnd0NxDhfRcwDLbIzXPjJ6SZFwD42RF3KiN
TUO9gp1NOxqClZleC8SNuPRYp8g8kfH1yNHD1bkOS0DoywtMN5PU9bJp1oW9WhFd
IRNLW8BdoMrFgF4GwL3HKvz6phXm9NSi/3nfjHL5QG5gesp+zQoMvhF1jaghjd7m
gQUcUn5x67r3dlS4kQrhQiH8adG7N05F+EGP1+PfMwnqp4mXL2000gbmZd1j1oBb
NjRUzuuB4LQFvBeM2Qh4eswNMi0dT0ycKRoMKjTfCJSbCJ6pv4nTyCR9o1QaDd5H
MAxKP+WpuPWhpmONefCkRMAmpE2uGESHqoLwCe9fkGhEmHhI48eyQ9SbsXJx7YNt
dznnOdh6XiVqIFb9tzznmV5qVP5NDzmbL21hWS772zR2yQN4eVsKTAHF/AbDQBsQ
ze51QPKeNBB6ypp/aMeryjZ4qQUnlpwQeufwF7DzqE3ufTvmpcxDMB//DlRG2fID
7wm299zs8BAGfJfCdziUyf0GYxmeZb4iinfB5BIvPrYYYIAJ+JrN1dJbGoxXowPj
En8k22FxFsPOd+gZZ7EToKQ5el6VQGvragpQgdhvJwq9IMI6DHsY+pytDu+2sUNq
3aLR2v6tceElALnS0xM5KAblUCaiBTKtsr3ldY6BqtDRaAVRlOMGlnAOSKhQqnyI
EjulLpIT8ytq4CwJnVt+ZiRzRviG5w/K04Bh+UyryJzDxb5xWnEsb9At4RvaHUd2
+aOJrsW4Bg5om0CXnUKzh+/Waxhwq/6k+R/wtzagwGsSll6MgRE9sNx93w6t4bQ1
QcWcijrVvuJWqiT47Rru3MaAL2LS/tpaVrcTMWS7qAQbXmNFG7uPqnMdJqkytoqT
SjBQbPKrCpkjACHlKaEhBNY4CA+p1OiGLclMkRsvIejwf+f9bIMJ8bmSGOHzMjF+
BsP/QUzErK4Yrq/IuDxDK9gEvKHXufIpX/j8zTPGqdzsbYu2PxP9XP9ACIFlacOq
dYQhUhsoUB2G8pSWwh2hP00HJz6+457YvqAcA5tM6h6rn3dpneAVHwMCnNPvQwwJ
xqNrNkqtt3xpqsRLmVo+hb4asjNLLtFzEWanF5WUcEwabCJoGr/7EAVfNcjbNVmL
E5IuO/G28W8qMTlCYAufGO49FXcALYbg9bNcwCzUx/9l9zJZZkojhWv306QLp4yN
DO090Ks3u7ql7emKCu27h59fCLiM+PXccJpiKERAdhfKO57mY3DC5KPmgeh8Qe5u
8BLByoVrTHzxDAMajp/0KIfHXoNwi2/Lfz3X7zr1avwR2tnESTbUjpgOne3ksMEp
RlpuFLetT/o8w2k8pbC2Ou1m25Cz61/1Gs2MgNoB4Y/EfLJkuh1j6vgmL028jvqA
w1JE4z9BZrt8sKCeMrVFQywCR2FcV+jMn7455zHHaV5SFNlcgJ/lZ83YViloE6MS
kR2BsP+OMJapcn+n7yYKANPu0pOlfkibYQLAEXqmkvnwjHsBetvfjY/2mcTEtwWW
WE5lhRCKampw6a2qAAovecIUVgWkRH9cBmyNFz1PCR8yoQPexkmlp9ikB+EpCGG8
TxoDgKGsdFmdEXxd69ea8A/RxlHYroEsFbMGykkbPNSOthxG96X28QDhoPpHyO7T
zmP2p55/xGD9rJQMVwEP43oaHdB4HM3y/hWKivG6ih5aoZhZ/xP4Bm8CogmVMF+c
OIRxQ7X/ATdVforJvqxFmkrGf86qUIJV2K3xKXCfiGUQyRQ3HUKk74KCmzWv6V6o
QX7AXSl59Tk0JcC7e99V4Caa7bNyBseska+Zhxa6V32MKc4//7ZmxQkBCoOe+8sS
nZPnus6SSayDYexsiLFfaSLk1jgHIUSd4uqNlOk9TO0uk4HakTFbTeDkGMGnK/B3
8+5j/rJcmTs2W6QW/YsK2xfMLe0+i2Hk5n6x9AtZ/6bxJHhTQ3xYbgEMxPv2Rz4U
sUOY9oSA+s8HwIkqUxbmGA2fTitMcUHS5pm92ZC8jN0xqHWJbiLvEKLj/lc/Egnw
jSDq/7iO1HjQP7v1AicqVbHsE+AGwdiNpoS1Nf3EOwty/mAOQXwTEf3Hy0EzAIM0
cXN5IrWSck5ZsFTLIx0zDw2jaskT4TAXWHvDNu6pY07yuQdmqEEOdx7NLkI8R8nx
RAFyb/pRQA6lcQwqmNxIgYW6eUTKSPSmb3o4z+EMZa/w0EbNpSPBHku1sckosRtq
V8+HYA/CQox50cKh9KXlOhhM1voLZINeqmJKI/JGztjUSBScd2tyv+/olofJ65xa
ecQKkrCznh1xNoOasCxFPMW9/ZKkU0f5m77aars5osz5hFMeDho5Ehf0T2+E17MR
7o8X8YwH21q8dMLXxY+7mrKRKOPBG99mBEKPlaTto2zEWrXvaXTLwjcWxDXNYSaI
nh8wdQnAK5CeYSV0AU2+0TskcSuea1BZ1I/ftcVzJeNBOfWB4UQ4LOC9iJb2XCFA
6DXK4/rRGPTcpxWK1osr2cIG38vcRaGj8N/6i2nXlEYpTf7t0aVw8dMPLSjgeEOk
Yc0Zvx0bqhp7KjYk7FsEv3i4mCRcrwVJzRdZrYFDsk/Pl/RGVDsE7yEaE/56AYXa
VSP7bbYi+riNaUwZEo+LuuZRUSH1h5P0GJ0u24JWy2o240noZjZVSI5WLTljDAvD
CysJrVg4X6ACZ+7OAkcBO70h/l1x1fPxZfg/pArr+bGH0D9TtA6rv7XF/CZSFrkH
71mK92HZew706nZ3n12rMHykgVRkq/Evlco18PFYb6fnQCYbtOgEgoMA/jySuqTr
MPNjuEuJkK5mAQ0fZyCQt9PuqmPKJEnhA2wxXs8WEcgmjLGQsnNUsWUa219Zr2Oh
dfKwetKJp9WxA4Potqb40eh5jvT0GmrE1HGT29B5DHHh/c0zQjfJxZeGwjCflKxk
yxXa4Gk+QYCZdb45KoXAQxMPuNh6JLWRNC0dMr3JuwyRpbbRZ/loq5Uz+PcktQwN
Eq9ExaAQ+6TnMtWSTx2MsMJ9BP2YXT532wb5usTmenwzotMvCVK4mAYFLIiDQ2yi
mRyxQzT+Uudv9SNdeejCAyYtzSHhkjuIFIRjtD5Z/IEWK+BSXc5SF5DwRwt1QmP5
N/i5aftq1oHzCiTisv0oxFX4rJOr4tFhauBU4RRNihXDVcXKRn2B1p6dFT2/Ak9r
GDWLh5ldPkZcGn4Oya27KGo5bcNNKdIPa3WlDjTWU6uc4aTK5E5MV551SRE2JrkL
de6pT4B+PlHBEal9WFh/otxbXqpEwrGTu+ty/afUMOEoZcmj4o0wg427GOXlnWTB
+Ar9zTRKrR3LQZfO+Z0HBeb+Hp34kxcApa31zJu2sSAirufeca9VQOw4Og40IsqC
HQnWdDcyG7x1VnDjchllo58YDsVKdSCKqqQs104LEToWnbiSX1LCZBGKNFfHDlre
ZhqpNoXl73zziFdAJqTC/K9yhO2pTTv35T45GDqlD6LEZnrYZ9XBP8cDpDHK2ZKX
vk1CY5Dcl01FHaarz5DsasJlzw52O+zm3N4iU57/MGFOinORacantOgoKNje0D4e
2P8ZWr4uAgyrrcJU8puqmyNcDCHK4ElhsqYnI68nAu8b9cOkGn2joFW21pTtfHJn
LTvDT/LBYBBsFuxT0syTybAxc+fx1+sQbakfd8VzRTeLNJd4jRxjCbIgNOzI/ZKn
VuwKYeZkpg0LLp/7U9aYq5FViFpHqnRLG6Lc0mwgmRQ72ElICIdfpPkMuSaUCFSQ
VRaPdbEuO9cga/xgituZZKDQzokvqbcb2SClt5/przfmaaivQUnOLJnEG0bUBbTI
Kqggz3py1q7CnvWebNZfzQ==
`pragma protect end_protected

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
eN17G0wxNGPqILdgC427ezNcdPLRsK/aQVyABRY6k1lIOYaYKFIvW+3zlqrFB79n
p76GuTp84E9H1l33Qu/dFMfjToay7pTRx+4yQkPmafcGLqk2ONeoAM3krXT2n4m9
bn3aBYXJjRQawsl4b2KMF2sqehRn4j8xK7lRD1kdeNo=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 36832), data_block
PWSXW+bvGNhbWn5+4FMhX8kuOc2E5YRL7HaEOb90Y5cg2M51cqOs94Gi5ztND929
21ezMJQBD60hBLns1iepyBMyVGgHWn89UmhC4+thYSoH32h5fm3p/rtgIWdAknl2
MzEajO32DVseCnQTA/MATpDXDMFjayTXPHhDtxboS5u4dYJa+tMtVNNrN5z3fGSk
0XQIGEjmGeyG5p8z0tGqv0YrcVg+RIExHHoz7/+V3ZbjfDCqtX/9VWZYacnu5qTN
0bPdd54XfTVnDImNgwZ/VnpXMygfcFpJeUL53zgCJvIkuOym8Yh7Lv8NxnoCEZmW
bO4tWnyNSmmJjQdbc9jpYveQgiR61W5kgho+vJoUhfn1LSrjpeBJuFwuUwYOXJSz
LoAkWXKE3aYIndbYKoNnAsYFmBaz+4+XXaYznFNRYdKkyUewARKMX+RgARmL2Syh
/0hrf64xnGWOUhZ4DnNZL/OYVHAM+qrQKWhD5mjxBASIFfW6m7TVrYpsQSo5NOnx
/cdPjF+eJHOfFFn0SDAvn2eLldrcmV50uwDC8WSRKWtlbWkmGVNJjOTy4zgI7Xc/
WpQ+kiP67yolbf/1b49QADiqFcvgmagisRlvcoIy+76XjVt+eLtJHxSgOdHSshlW
rFKGUMFdHwiQ/uDCeg+yo9nTGkBymXLyV4K+o6OlTgcEAwRWK7xnG5QfDsxdT86x
V4eXD5xIey2U/l7P/CtMRYpiOt7JbchvrJ/INxNAitbQ7Zowxfx89LwTvx203SXm
Yy9bRM3DmCgbtYLyS44Wh8VFIV7rzmskqvXppbCmbuo7Jj5OTiDO4lbE3iiQ2SSy
Gp8ckmjK7qF6lkZT4M0GI7W1Mu1pVk0xwHYkGgT6T7bvF/8zD/P99cg3upD15UTq
o8PNjlhITw9tIJePmdQjDqNO6TAD7Eqvk2rb6W1gs1Cw2LQpuG/0Bw4tXZR5TdEC
7oRlSttyYnasFDiGvDyX0SzUyjVPldEo4YYjF7B/rFj0ynNKCW4KVrQd2JVUya4m
zaWioyjP2572AxqRNTclKsCgxgqzXXP1LUM+Q7HcV7LX4fw3uzcnvY22Yu5Es00A
2h0hSIZLlT8VxY0xvCV73DcC9JrixiCN/rItHG5QNH259qBKDeVovEeIA3BHzfLy
ni89q1U1V9jNSNRTe744onoJerIYBYL0BQ4UhYIPI7hKcDR16+ceQ1nyOjF6ygEQ
6eeRYfvsievWs1hhWi9J0diVQrhYn8mE/5j5W+rsmqH7ODZzAKpQUZpqQKPyrtji
oG2wi9yfYCPd/FfFcmtKu1UbYKxAMoNXk7rgywoWDnS98dkWtj3wChYIZIClISVZ
JkX1Ron7hDpkgGR/kRc1v0f25ujUsUQ1emRPZmYeC+vDHpY8yUYl/NSQKXeQEniS
QXQVRwn1bF0UXqPsli19iquCcMjoPd1PmJI4r8nlbPYNEZEAobiQrIVIfD1FfU9f
Nq6ftLBTCO++HDDEZa1Sa8pSyNSqkEHkMWJIZGWTvPQsJTH/rCVrBW8+za61ECMm
JPEm48blxIS/bnQZQqjUKHJw2tvOM7hZ2wpYGDAOYpKsrRDgqtldcygkvLAecXff
crmJdaY7Os2FF4aJ1EOWiIL9RjjSLnVFw0FM6NG/a32fY/MRc4GqFe5BoPvnTum1
83qWd29h3GjtlomR2CnJOa7KnkdH50qWs2ldeMVBaV9rQ24YFgzL6tt8XSaNrhZB
WwmNt8DfxHKVeAm/w5JpHd92dyQmJNBjqSON6WORRIrF1C8qoZZkI8+/Qqe3s/5w
W7KME8qtSz8B4NOUvM6pW/M67ZoeAkPy17TivlhrddVbYjayW7uW8NDg9JqiK4tX
tzIJZ2AzodrJXwce3yBK9ZYG/rov2qBb39dQGOpPzmhtAPfBDvU2t3/WeYhPdRFh
ibZvBVVvjbIDaxDgDoYnjl9sSJRNDN6MmO7VGWaTG1t9kK1Cyh82RxzR088b3Dsm
2xWgoqhpnpmdO1+u/5tuwZpDQOuYMNOFoPL3MTKepmKyAj35autjDwvfeNHeO0+O
jVjgIe4tIFWJjqhF4IgCKXx4Ygl7Zen7rhuKyFrIaWXlwLi5SLFmP6sR0sVQKAi0
1GYM9N7ITg9CmonPImhC9OrsAXQPrZWIBmRnJ+0jKdJvgdfd8tlol9YDbD3fRB5L
VqgcTFSwNxKT06h7GENbUHkSRQVDeEfhtgtTKUGnW4V5fafrPTzk8YoPFVTytb8v
oyEGnU95wPyfwzqZlZW/NKdVICVX8uEuhWV8D9OqpyDt50MD26gDLQ2G4XqPEE7w
Aun5jOZiIndwLmlzfuWFLLJZFeZPRYAhqauTAc+70EMuiO/I+l0rQjgKYSiC3nED
0xOBqN+GYp5qHT9xz25Odm7wVpYW3bWmzRURlswKEsKw2fJKX6l6ytX0UhGYtMDn
q0i5pW6NoMzuvcIKmJzEkSMJk884Z0mjgh5qoTuw9Rd7BVEp9e6y3S0Jd3AFmqLQ
1xknoVQesYpBu/c4JoRjYbmyOYTQ/+Pku+++JXF1jpnWxbwIMWSIJdyTMEskYWSr
DCtdw0DivXruy6fQF98SDU8pItfeVcukpJ7okz5WCYc12GGGdQ7Q21jnKtDKSUbx
qOrNpRzuUgW26uAWXX/rtGORGkIvHC3ZIHk+Dytwx1eOXNtDgywoGnoFoVdBTvmw
pfy9k/XtdmWQ4dNXKh5y/iB3wzGiQCzjSAx9x4rEK4EXfjTGH+XFWcohUZXs6hPY
ChvIa7s52LhjdA06xfZftVfIkiUJmDNChUglMSvDc2WZlZzKHwmC9sZT3/SzpRIW
MbH25chy4sTwwdrsXcWwTIYWUkbAHYoIZ6fEypZrHx4RzMOEm9P5uI5qRibv4seZ
jAIqFxi29lDh2q35mvorEO9+DJ9W+4QKE0ESHfh+DFxQw6v8GM/OYIlq09ctfV4c
hC5dRgYuOPi7dxnBTkWRqbzFaWX/LeHal9S3Qb6TCTupaHrcFndMrxHtznXHcFhv
yjUM6+GNQmitnRhVahUNSQRyXFJLT1XjsLFegwdL9RAts3IAC1f9Ax159bR33I9V
9juK8oAUn4+peFXR1GsU5EIJOqoRUujEfQMndKWEKjqFDeE9Clg2Hv6kNTHqIlph
WB+76TTxqECHlxUZ1byQjEY/8BGKUIWCkdIPitu0PKWgb2YSlYghl7cgzFd3UPTw
xqN+RL43aXEDDVSAgwo87ABCl2B+KwweKn507JRjk/YLG44nBJ2pnb2TQLJlCi6i
30wfHPcCFLrvuL54rDY5bFbX0XrxWn3PMAzmYmmm5WtEdLR0TwdtjW5qcDx+BFzK
Z7QmET/q8GZkEwZ4DcYmnTn9qNJmhdt46Vcv/TKMMjBhDlTU8b8FW9QGvdA0X2i/
HltVm31Qe5sOC0sbLSEJ8iyHlLphkDN59bGRmWw3hQZpuGjBCNl69Gc28H9DPhJk
Cs7PcHoXVVTpJi5UHMv1vgZerYmdlW1jl668BifV1Sz2fXIa3KOKiawsnonI0mrL
4iQcyhOxK8/bXZbgWAQZX+qgrOHQnGVdcO/no8CpOwVd3kKhurZz3pFZcZ3ia0PE
4bwFnOu89iLkY2Yh6yNgLx3hW/yKxx00dUeKe8UH0vpH4hG3cuzf2h/3pVPrEM4K
kXpYdJHJbRbl41b/LOPTfz5LS+GtaGTY90rwIJCvm2usg5P5RWQayfm6rsuo4hT/
36VR0pAFtQ0D8sXAyh7XY8V6Vva4hVl+Dc5DkNRiq7QL6fxTsnWgEMuwiCcM8gQL
d2nIQ4Wv8Igc8CB+u4EU4J7DyN3j62ur6dVeDY+8+tWvMZ75a0ORJUOsBlb07DQx
fYJDvnHRa0SgtviBktmua4vZi6dQVPgBoLMIvEfVU+8v/5wqKOaJ2eDB4yIDjo64
GWxyoIy8yMOOTuPP53oqoPu3pM89ezId5IxHkz6z2oTst1C0Aj84et131jGtBua5
3aTXLU9uZh4MUazi58FSBrD8EqrRq84E09E5nYZQqvZXqwvHkQ+2YvNsZZ5JkEnW
bMHtkRu7jqk2/9R7Li7mkIh5+XMMKDNEDzrRvZiQFA+mwUzygw7iJHoC7aPbA2pZ
+FZUFPW9pG+3fuU3XOSrsfFqqak97hkqBRNV6SlW+jXuR2ADqcC4Oj7pZobNDSOX
/gYisRB5j93M6KSu2DyvXb0wPLATXaLnO8KTVhQoub91fIPhjU9puoMdooi9URjW
UpYy1T/xfYPbDVeq8MkgeViPe5mw0NZth3efS4hC0kmbjX54AxDwkf94MsnRP1X3
QIp075ib8cTcEIwWn3y3EzVBl8o7GuK5jPbjhwOXpXFHXld+mXnpt39oUsXRRWga
4zR/uR/LAFrZEAxH8RcxFBFwsvL11+YUxeGvjK526ScY3GdD0TDuoAL1+dJd6htc
sfWQH8Sb+GQuQQdTqVxOgxeeDBF99DjPxb/ZiWRpVj8jBuS8Xhw6Rm21kfm2ojTY
36WRJApsqQ/CoCame1rHR3gvk+GIBGkoV6jQdEEw1Vcfs63MO9Wwe9xAi3GJJBPD
pPZeT/dOCZR1AC06HdOpxy4J30I1GWXqXkbjZNXN5ZQr1ATes6oeIWbaQQ3AdjZZ
f3ZV6nPOfn0fke2XlukFtEg+DFVAF/voT/xgn0R4uU4Pz9XbHw/fcv4H9xk94oWE
xIHk+bz5MygxI6VCSpk+Hu4S7LEiKriX7sgFHacVy8YwOwI2WJ/XHTxMKNOlGOQn
PZZsdtcBmujkq7ZrjBJZx4Ieq/9qw6u7Kq0cLUkpQHXhruQfo+8bDw8LHOi0gI4u
JfsJsIO80W1lUaR6gt62z8tmDyGu2c6BUXfa8Io6TtGcklnpb3TxbbTHq5gRFTjy
IxgURE0ASr5apS581ueHgmnHVlGOFL8Hi4wsxg6C8mOosGMXa3Uohm0vtg0MmcV4
clXwxnepbzhWEJ7wrqD+BTg2iCvi4kh8UCqneIgzu7ngx0cwVF7bUBFA4hMvvGJm
f8EyaMwB5YI/LrW0aFQoPiD3XHXhJhYWNQuWCjDvVnhGxdsTc6jJJPtdQyw06rN+
BmYJYsAAEpkJrrXTgBh1uWbvMGdD5ja4+zFPRDUByefoJAkREjpMfvGrAmRMy1Qi
AM2gayUl+4LHJykDzY7+3N7pSmJkbWmQQL5bk0vKjc2PJswiEKFgONRyZqAxpYno
G6DzJjHsZmyQMqCsjHm0+gjGNkKtWjE3pFZ79SXTEJEW6Yrl2YrSSwwjFF8ZGmQ3
fyuuqM9F1L917wIkdyxuaqJ7YjHsFMnDfFh33AWpb0tuD79VPGQHHdP5NwKxsJ1S
AGEodWNl3m4LmCMWSxqpyU6x6zws9DefcefNUD3FlAO81+7lpgQ8IED15Y2KjTIF
DyFEdHlz0X+SlDT8QMLoZX7V6i3mwQnE0CP+KpGCvQkH82q1wZJxE+mP3FwhT11N
ye5DbEYZY/EMcOPbRFH+YJEH+CiPp2baFKoCgfLngZ5hP+Q3MZta9gPw+f0+Go4W
0GARyQ+cmfF6xV55mfRQO0rJ7OPC+BzANZk3cws+nyOs0OkZvouFPni7xli5lIWF
PygUOPJo24wiaJMLjCKnSoYqi/PAWVwYVFJRSYXKHMJ/E2NHK/2qI4I+SNkzP55C
hvzfoZVHxMG45qbY6Kd7BGhx6Cjv4EoP0qZhqhuF0UrGxuJnQuz5I/++X1aFyOVS
dNeab+PRpa+EcTJS7S8zsHMgRIE4Y7edDNZv6co1Egp5tz9yctvPgerRqHR0xx4p
AE4zxq7/xKVB1lnx/Hn08laZYBDrChpMXAp3/sYI4BzBwuSdM/+rrE7/9ZgULRK9
kbNR7Kq1AbP0HvBs0vZ16Ya8JxhUSJjUKHSwUDAxZgBcsJOsTe9eGOerh7u4Kiq8
zDj/i0EE02Kaqd085Mokobgp1bf5tZry78xw53TB/FfaHdbsJG78rJ7FxS1EF9vC
EIc8KVDQYOOLcOmeJ+M/5PdlQc27JPOeOYCq/EiqRfb78TT+QyabnoQR534NCSj7
znojRluAQw95JD2EZs6FmUhGBMKFRyeXrR+fQg/bBjf189xzhD0n5ZFlZMVbPZyv
19rI842sUvaH/I62KUjXEUOHVyfxN9rTbyay/aAcY5kjhK/erMlHa9CWhIa0EI9I
/IbzG4/PBA30+M8wP5hoagRQNwRAbm++EAx7L7lrKTvYGIx/CjKZ8zKkF5JwjQD+
e+GtSK5lZIE1Cw6U6tsyCgf1w8XQFeLD8EmB91ppJEsi7pCI8GcWEKoMicHAC86Y
nlpZjAPWSX1NgbXbvXQNbavgGAGP1iLqleAEXrUSQyFi+2D+Ng6rSARDxxvBynF7
NGXOXpNtzQgyCZALlYEND3BippdqKehoYiFqUdIUaVy8PL/bUSmajueOn6wBQk67
VoVIkSijjRSLTpSAvon0peMQCMPCW92Cqpg6yO5YNuoMnPcFrj/Z4MKuLtAM3/hX
Vlqe6BW0Z8Wcts+EjYUjAwq6vB+DdXR2DslVqNbazSfEGxIGDmX2irhcHxOcUTmS
1eAx87t4F+nQrj0kS2ucPKmxsO7srMkxMdL4dyX5GQ7uOiIznnivaS0AfsdRM/Px
BhFC2FTwVYVWjX+qD6V4hFp9zjLHOK9C4bFL3zUBS31e/SEcjII+Wx9O9xfBzgY7
CWJJeOgozKdY1ajluthk1Mqxc7FI+6D1Iw/9aPcIzk/PO38JpfMAy237RS3X7+SR
QCcpXjVTltnwD7JaFQdK2wDA+3+0nC8DTIjSvOzXD9Mt9lQvmpm+xRgjlSnLRruA
TBRvFf97mrFdUaEBvlkkdHYZRIr7Ut6c3pKr0uLYuvZQ4Fgbet17I1SNUmLTaQJz
MXSPQZE9YC9m8+OVCddNmrJOxfFcSGnb5cVhGhfUgRl6IRqOxK97TtQlqjxI0E5p
z5jYiy4zWySKhaLvfQiG9RO3Y2wTFKavkv+GymmSoXGE5A95IDtdOkO6gPU7Gct1
2lffOd9EGRthgjqjSGCVWxGGI244HbkOoliR1aBY8hWs33Is/XVOtd/r4UQIF7pF
npEBfKcS04WoNtNVlvYjNuCQnIiTcRBpop/skwZAfo90/hkixJEjM3fBO89CLiwH
bLu8t36Wu96DSUWXVSiRU1KwaCWkGVz1PNfmxPKT3ZxsjsLPjv7Pu2/KKSgvv+Mb
FFN/+cAnBRRUmYvffkf+vmIIzLcm1amR/zCOHV0DckUdHrpSe5vvVnnV9tY0gcQ4
aUA7EyhTJuYAJoALM5dC6FcF+BSsrjqsAqxlU1IEAD5vhw48j+V0WLMBbsVT/y6T
qQ1GaordkPe2jL45AIDTMy/gvITPPXWIT12GSCeHYiila+9X/fIdjFVo2nr7J8Uq
I0WGfnImCj8aFghdzCXoVgb1Dl2EzlAEjkOXke8WN6bZqNcK7fhsaECs8XbWS9I5
lcF+5aoTpa0TD0b/KAFvP405fgXptMZbJT3QOZhVUAcds06GdQ+J69JEzZzCu94A
d0gamRnYxoXh1KUxzJ8wkCmGFaB5TZ3MwAcFeRvyePF/KHlp0QRvp5rkaogmW9Uq
D1vRokuTp5Wz57s/qKOI5WMxgA4jllxGM3drsSyXcuP0eXYBKbsj+m/vECPuLSek
76EJ9x7VgVy4g/QAgZpP8O16Jx0UhkzkokHZ20vbFvtnfrDJoGgienx39O+xGbLU
FyO9Bq0Ycvkd3NY6uOT1Dvdf0BaLuzl2cEekoApZuUtjus0fVoXQ+imtSl7BJgew
Wjx8vne4DXxsAbeQfBV9Mf5jARuzMBQNXX6Tgz5o26d3/PTzevUkRyJQC1rXFRk7
gWCpKhJHQS44SXoQclL9iUOiXrLTvtwX0oQgw+J4TXt3yXtIYHgRLhwRPib3XFxu
a/FVO3/5TKYtLCFll4LD4PvWpB44o89wMxkENhz8o94iicMpDio1NE24D6VGGul0
oz/7GO2vE8U+RT6RwBmBdfC3Q67WEoqP9ftK+HFepJYd9sFark0cuBtgvTzz9Ro8
Zkvfb1dRp7yF458gksPrbToaTybsih4m2SGj3QXHdaNJCDGVaDiMOX7S7O3A2AMc
RJ1K0MUKuKt8cPYrIsdnnOAIhnuYowkbCx+SLGS6b/0niQil35WLdjlO/6wTZYt/
HGQ+D5HcjDeUJNK1awRP7YtfcZqySS3vcGXQyr3/hkMbBH0dITXbtr9LMhSJ9Af5
wF22vFbWQifF2dr9T7BrDMyuoSAcDEPXTMdynsrs7UmZVCg8RHKrdj9a1YRHX6N8
4127IOCBfkCQJFhWj0aAcHR83t6cNRIc89ybnCxOlA7uR+WGuDpVvyJjPZa5G23U
ueyQQF8yq4sEtUkytT5TbUU+y/DwfHE+IrCnb71rZlYJIXL5DBQpP/PNStSHBe3a
cKjTZztqUzg11DYGksi78dpFStbIG7gCQPxPFh9z6/omkYjCFiyL99U8VcNxv7lM
SukhzQvxG/6/Q+6VwNM2aDTJpp4F7dVdSV3H+pOTJmliHROgzGSyHXVzNLBPdSZX
PF16IiO/ieW7+bIxfWETCH60/WuLFlAD9j2SPvcI1Km2OKFNqkgDz/CRwzQaFaYs
w1nJIKwotvFN0WSBQtMgRcjb1A0uMDm7DUc2RG9ooQTNkKfnD4SNgK/lXHci1y7+
c/FbcXYNYHJ94QX82ipIAE+pYmW4BScxCj0wwOMgiGhmZ6aFBnqbMg+G3soFH6hi
iiT80Y5/sc5RooiyyE33djH3vd33kretdhmbMA246+CyOL9WBvsgyCL/S7URju8s
dnjeDO04NaGB5WwFQKoYMnUf2w+n74c0ls3jsb3uvGLh4iCUeWfRQmqpFZCvXeFz
28DAt0kWyOosuLV1zhgiEj3SEL+K9tgTBrnCQrfgBRksx0FsPBQABZB7S7QW6mey
FAtEsNGpeXZ8JsPNvsTUC3JgumhERw6RZTZnz6+HRnC0R2++zOyOzKmaIMsjRzSm
xgyI1uw7yTkXxZvtzzskzwK9yc9ODs+XvWowoLUOtngqTQf6A8Pn5r568uTGRNUZ
ZObmllulzpuDrfibwuoehnxMpS612iQXfPKrMvctpFXAQ6p605LY3mIDjJljbQMc
yOCW4e+h2tdxOCKSZpOEqyiU2Wv2alWr7kIl2q+vVesSEMqCDaM00YXNXI7Dkv29
ufMNMSEKQ6hclvspUpoklFLpwNdMxP6JbQ8wsdGn8IgFmSM7VZgPs64+f55G7CCx
KhYO0iCJ2Qy3RT1IwY4JunKvtEmMpLNA5Sf7XRGUvtn/cDPN3KSS9Vd5uYfdD+1D
tMmsKnk96qxjDgY1sHGK1kDUZAZ8Ad5lVgSqNckNu7sk2gSCD7kDwlk+mrO0WNbD
nrbaJi6p2ieGwwh7EPTXp1/F0CMZX3peP/YlNNP7jLkeq402inT6e8QzmyutBz5H
65sysDXHoyv7seE12OEB/iXm8YVdqZtn/EOJ+UxonT13YR37Wxrgjk+A3SeZHpkz
nzUrCCIVgnJMregp62cUcouBR9TEGB4VIbtBVcVrJHjqFJVIEZtOQcgImadeIzBp
H+Mvf5R8F9vgqeE+JDa/AEBr4EJjOG/5+rr6+5dK9kX4fL/2kRDQrbuQwRdRU8n9
BpEqjKDQYFH6/c5c1VkYSSj9uk9GiuhAEqC4emGCRT25qrdJ81v5gHK29As39ZFJ
lV0tUjAG54VfgBraAFTPxx/AiqfwMwQSv8S6A99etRDl2sbHQmIfPYBhu/LOY1iH
SxyCRCEHFTD3pW4ospsKMoBn4KEWSJQ8m6mV5k36txswbp2gbfHUL5tIN2CbMfMe
0DK2VOEwEpsQ6AZwrA5sqbE/dBImXtODJG7EMwX+Yofvr0ZCxrSeMNcR/jaiBwkD
+DbysW37zn45EIjPH9LhKlnw5NQSfC8diufU/1q9jr+TN4LbZ1zsAAWrqEioh9qJ
YBvvvU9gcTXHeJYak8tM2klfoL6fDF0oK+SFvU3RamfldzCWjsaonpd8tMUF02La
XBSIdi42XUFnrRHnsVj4LUDYnTn0O/PcrBDJEtbTl1qsNnkzWu8Zxo9IvuU5o5DH
Xr+sg2kMHbyMT2aj9NDI1Vuy6pO7p6Pys3/CD2o0Bhf1FgwpNsc3GHHSV3uMaaPW
SgZALYmsxRSzJ2mU1P4EetyQE+7LvlkQJsjEC6XAskOD501HvA/yeJrNu0iVRnuL
faI8XCWrIsweX9QqVjmKRIk5RdD1N9hEcgzHxPMadNHi1JzUnmcfr8ayJfwZUQtT
WWuTNQUC3kvgi83lEbx1Rt4+pk9nYJHgdo0qV2NGPOYsFpmySqETAztravhJPWPe
4fGCs3XV78LEY7j6+gTWnTi+a7bCo+PzHeHRQ1W+65SmJ/3H41b4DfovILymgb96
lPm36Bg6eVeKLFzgQcxbKsF/8xvJR6juF+wJUbnCD6cmEZIwWQrDGc8ofQYRBPWi
GMAb2cNEH3Cz1zUelm6rcmaCVg9jwenj685SC2lXbYGj4xiMac4L2LOCldSucbky
5b7vOlOV70w2V/H7LWskk9FrfeBzy2vtKEKi2hu8eeejiyU5bUpsYz2UeEWmp5zT
wPPT0mH+SqwA0t6UuolySaTiw6eBaFANBclLqHLeurDbouqZzunogLi7T9+hYghy
IIisTzGVVvtgwboTOZOoh5Ywe5ayl37Bex0zOY3sg99gyNOZ/TxIqXiwabf2q5IH
eg+j90iYwIMcX/8aBskQiGfqBdaMweBsVngcKQRc1H0AQ+euTXF73BKyHRRvWMiL
8+2/tnimsLyFK91QMzrxeLBqiwotqsNVaP37k4PtfKMRtWluYONx4l7sNvYJ/Wo7
OT3nFkn0TI/qViwbWzRdxYvt5wMsRSr1mYD2pk6ipspXk13sGA4hcf33hr9q1Df4
iolNaMGyfUAo81yB6uLJKFPN1+15AfwDbNqvq4ZTQB968Al8dLkWL5y+hqY4spWk
NHDiNASc06nutYsilOXH7h5j2jylgI7QnWucqxl2ajIMD33oZDWiuvKEAc1ox5rs
xTuDrQnDjE8IUWs8GWi0UD7RIE0b1qjTBA8Z4neT93k7m7u1mqWEUMx83Ok75PbP
UugBJpZBasNZwAEs3+hpXlJ6tqaJXo7bD+4nppEog3MgdOkQMN6v9BQT7m35x3dG
OUnG6d/WdgHBT9iPYM9lY6LNXcClBBau5iLE6SiMEutXlVV7CEtO2YxuHMGlw7nr
VKmTDh4PdXv0hEHTa60Jt9DRMSw45qWEnIY7+DSXTcQ00Yr9gkDeaPB7bFq/G5Aq
2mf4AACxI/DRc4176vDPh7E886Vkr9tpfqXcij0i83xDxAEvhbykVivIiREqt+6S
Km6RLV1mb4lROLPO18V41v3cBQKPhA3tH/luvzWWvo5VinSTTVUMqxtIjtrudFZV
nCI/f5hz6wcW/MvzkPjfMHjdDuu3uKw7oeiYE5sG175dkv54vpDez/36O0V8KJ4q
qZyvcqIkPtyTUDbxGerGEwHUniIGq+B7fwAhxazyvCKC1i0jCATQDp5A8rPLeN7C
nJLCvhjHCu4fNWi85SDCNKPKJMWxNGij6bGok7c5iegtGUA6DnAB1aVxXv7ysr/j
yEOqA1pjdUkAXjnhQdCwbTLP7vLVR0QEyOM0iAIjaNHbl7HAQLCuUyrC5tYMEeGx
qAccfeHGk3uBtmUpSxm7pAjzjngHDQUzx9HT3rGPfIBtUdnJ12sXkUwoBQxIA+Eq
g+s0ikL8oR/l18FZhOdCw1EW7egwFHE4Wkcsj/N0MlAZ0FHSbGLLTAOoexZzza+X
Fy5UZ5x43eeunIIWMIZJNqt3yBxhKYPPstFUSGr87JlSEtvyOq6NKO2ZTzqY2COe
sivIgkvxIfVdkSkpBK8fDlIcOV3aXI0NaEeWH+ucSvDx23JxlVLVjOEjCYGsgSOC
/STsFXQ7jB6Y+QRZQ+bgtwXsDGruVcPkHwfPEHLbVK0nsUAtHIaMu+G5EQEWMHQw
5N6cZXkJTWrOq0Ta/NJn1YEYZaDpPQR+BIsd+ICXQS8wuqvoGl2Oqs7kBlyHI5Pt
gyF6Mz71ZykncGol0Qt+3eLXyy/IDgF6fqxzuQQzVj37t92hyVTLdU4r+WDLP5KZ
MQ0dSIie7z0TPPxuynPMeaUBPahkG6YqUV3XzGsMD4AOGk31jcPOT2D1wO+MdUln
DfR2gRG5fAvgOlxK0PkYWWPRPWAzm2ItSY6RNbKuciVYiE7iSkrthAqLjPNkvdWm
22jQeejKv2Z4t0IfWne1El91qRpUq76SEH/oxIyyBXsbztYMVm6nia1zzC2rwc9b
B0UYGRCw6kqwjYj7y56UD3M9dn3wO5NscUbohucyFYO62w46N8nelHmVjgUzTLDc
+1CrCp3brjqGn6flIbRg85lLg65ziWYWoObqT4U1TOabNUpH1+XEu8zZuNEfS9Fy
U5IQdKI+RIL7WfJyy0oW5U8yXm7RZm+HFGsrfziwFx9+viyZyW7otYFe/bhiLV0W
Pi1Q0rppIjyBiAYO4xTKRq9iBdTvcdqOIcp35aA38CrKnQDjvBAZLdYnLUrs8ECk
SxotRLv8kbs0aNmQGqA1vudZF+UVgW/buuyNjRNVqhhRkG+/gPTFC2Atx4ZAGf/l
aKhIssiDYZHYDP5CADXTkA9dGyHsG4K+wA5q4Zh/LtPh9VtKbw+VwnP03T7FhEaC
QNfl2RduzUhMfflYcXLzXQIAHUw0FEJMKdZq0dBM6eVkSXNylKbY0+Gng+zT3rD4
QGknMWJd+DA17ewqoFUrNQWZqHxgPZZGRw/eELjx4twBPWKmn4a50lCg2rSkB+RC
PZb2tF87NfbUkJ2ePCs4RflAdDQIbtHyvwdKmadj/jooeqkljr3jh2ob+WoBC+aG
k8nfBW01ZT0x6dQ1+Ps6NZ7gFBr7iX7s/KUnR/RBrSJzEpygHPqYfbkGQsONIsgU
pVEo+A2cNG5iLRaKTVIZj7AzVYAsCFv7nMoqX+HSgYreB5XGKITVypyNk8/JvAqT
ST/yio40ve+BXo5EmYLJSLEI9JTaSwbtv8bHVsxTBYamUFdeaMIGvy18NqDzRMZ6
+wJTrokpRdLJomtqv+crvNiX/Ql97AzII2YEMZniD96BwTOZitIOyTG0AfUwrn0O
ApW9ddyYkp4mRUr37KFoavPBmq+KTqdKBqYPo7WlJoUz3Lgndo7/Z+htC+62U00P
jJ1w/473MtLQ58aVzr0WqqTIY/LcmibkYxkIJAdbU6Ur3okADX2tPTyMW4uGM3+w
TJlj104V896SGVy0lcW30G+0FnGvMPDj413Q9hpCXkjPI3ITK/CD/vJLFqLsZrSv
EM2ZoY4RBpboxfAEXyL5EJ+LP/GqQ4gDOkdmLfxTV862BYMxMrfhr+RCP5vrphQY
cukOHMX4mFfy29c58q5vEO/AIP9/OG0WlrkXQP3s02/howkYqMHoF1DmnwcMkpgV
XOEnCuGrOEyq1oNz7L8DPQjeOyrT1I+m+tA4MkYTauxnh4RZJ3aK0WIxUc6FK55H
6bk7z9Z0YgfffvvBI047pMNJ82SOgtzsNT7TjGel8KvUTGwxkO/b43A9me+0PEel
78ONj2Ye/2RMo17RpWm+kMUWJdajBDQLCx2xF4ePsdCazRKV+1SYiBXZjhWHUgmn
bvzJZ+y9GRpL5SPEGjioD8TGyjRBX3ztsxpRCOMja4GqO1fp51xtSGfyuwBZguZ2
oiqQVmWsOJvOHJann1GPSEVsDtfD4m6AeFwWXQcj4or2TjU//3g8OzfoiObOkeP5
+NWYLuiYopzTuTs92JLjYi93ASJ+bvt8sLpegEQnEF+YiV/fNamLF5b8VuYCvKgD
n4xwk6e41RXY1inxpWCukBpC29yfUhtJz4/OBPW7j45KdNO8usbV/jRUCv/VJap4
8+1Hf63o/cLoI0U5kubIUHDe6a4TB4lKs7eX3inCCTQEjHATcwLvqbZc5/TVI/wS
orBKXSojyMcEYwkZYko0W8PUfbZjRgmfp06ECau5HqWIo98LTNQjU4BP7c2ODV7a
xYffcRTRZUPTzpLqVMlUoIkN30+EXU11zEl/1SkD6C7od3LpA9tq8vXYFnnaDaeD
snX5GjIG0Zjckpuj65A81q8GVthvJROn6h4GyqhXrPSepaplKZI4yuQm7+tb8qZN
rAUwiJomht45ut4+q2ROSW6pXK657Mjvs5oGGgstertoZop2KdL2/zRhC5QhYe6z
+GNKah/8yQqY21QeHymq2O6Mk2M4aoPWyobudxEBHU/YABlsR3TSaomHJ0Q8/1D+
iridg1SA+Jx7kBlULA31TyJZ9OXdDR11mqHIATmfBZ799mn1g4Tm+q0JFo4KMKWg
sUYQOX+tV3pM1mNtr5ME++xKSScZ2DU/inJQ73qDiSy/Fz4H0kzAhf88E3iTK13O
nAU/ap4LJtuvFpot2YfHp7rMOFbAJM0SR0+rldlyNqnvYJBryJYQRvUyjBlJmMyC
PzELeFSGRx43GLQu7mSUaY1ffdhu7gJjg/xRPC3cS2UytA9ktrWYx6DEosZmlrXo
W36askQ/5hwtLDY4FI1ceMBo70tUiKPMQO8ypBYv6/fdv40LAWAaZCPDbWUUvqbS
R0/NVj4ZEd28AKamvJSwl/AL+EWIo/uKzaQ3bMCQcUpuFYvdXj7+/+5AC1wDUiTS
tV7mOH2CHnZw+5H5CTzQUTcHdNCZ+pPnd7h4ituxZJ2u2UKYKN2Gxg6mhkEIK3on
Hybno8epPPztuulD6SIvF8la+zfk9d+9BjSiBYfSiSCP4SH7WHfqZpblntvdmr88
YJAX9L5IwmhkJ8mk9pRhH4s1qejkN4VIvsoEtmrSbxx7AxUC7LJK/jUhL7VR2P/v
dWe/il5sslg2Mg9xZX5wTndz7ePe9VxaPVn1I7PKHHZbKmtY36cKOMBWNyUKtM59
kN3BNmNiq4wUl3oYSh6R16dlA0Yhp/jHo7V500FtRtfbkTteF6GMWPPYS4TfZ4fN
v8GY7CCzfccCa6R6BciVDieyylMO+7A5PNdOZy9hJnqTPAepJ9eqsV7NdQYU9EL7
d8KUOhTHIY+qvWCd3p2xeZfwFzqivLEhljViUmOhTM+ta783bBj3ObNUlodZ5V4M
yUvbraCglaVaouZ3ij+U/Yd1C75bWxmLQVgE2qbV74uDX1Ox4oHlEs9u90Z3MCLk
ue+9ht/+z6C/vtvB3E5B9g1EBg94YgK5CHNzU7u/GQQwFXR+Jj2ycRBMS1JypxEO
/E4lBW7jQvlNL7lZ44F8JlIDYWfzXcdiVaJKvMxNPM1D931ipojn/6Fdgxrsz0hq
DU0MDtHRkGC6dsRctFh/5LcN01dfVwfOICuFAu1USMP3UaSgsTh0O6TaT1iKke36
P++JCpCBZ23s6bdKDECHk4L1XPAdzFHUjg8kP2uk13A0d3BjNdN1N8y6uBGPjEjx
zCjihKhOAa8fihuwewQYFcEjRMQzBaQ6i+bM+2k9HP0FtwxS6TzVrJs/TISY6OhX
3GB7OMoL6Q/WepYfZOUFxuMxj4pqT0W18yZBSpt/hCitku7DaTFDwIeLSLWGrDc2
fflKnl2JiaL7hYw4gXcY8S0tiZgkAzeUAYUNzl2OcIcWjHhjcNRlakI/uNx/4EoP
/Oe3xQGAUmCx1oHIH9G36xI/h7YaBCZWvUEeAVxM64LKSyWL67AwuGnI58etPZjv
+AUSR6zEOG9gNermvcm18xzSyKvfPuAr4o2EuztKNxySga0OglcHmnN+1oZX1Y2w
Y4DCOFJm7j5e2MljxGyogcpw9J4SPp8DCx9KUI7iNFYgf6jGrBl9UqiJrDXeQQ03
Z4auQbHom4PdM7Oa4Zu8wZTnDgGLhGWutFf06MAhiru/bSiYT7FG8CBivXeZJw6/
tLhUny3nhrFkGQ2rE16W1PI7BBdvZpXaFk5ts1Yrxi3pPCl5bxNiLv5cAM6AI0oF
E4VN8oMbh9SB4lJ9PRKwR3qBOmh5OGbXMsho1/vEWL17meE3n4onxutzYq6FcrIj
a38XxDjPBzPE4Gt+EhI0YSnmXkvKN74ekOf0A00NmRj3HWmAVj5QGNWPrQxfylEu
ZETWhGAbif1p+5w2PsHFF/IjuLT7nHAAvYzEZybctrrSR9oMlsLOe95Qu74KymE+
i9VYuWjiEon5jaLNHVTau/687LmVieITcmI6h2OZObRFafS/U2fjHFsv9IMo4bcy
dGVqDxmKw+mF8Wz3rw1w8LfusFONJSXS73ZJ6LFVQ6cVn2DqL25QgN/WkhstKPjP
wsZ+aOfmo5dGe6/xWuaY1Ys4ohqLPzY2jNRLDcuQbiVlsvcJhExM6Li0O0VN+Ew1
hzIXhP82ofV3+74wmKqIN8gHsctoMQolu4N23/EHWZtAKIak3xgf1nX9eeZ02xZK
n0We/iy+wu17JPlBmeRwinCietKaiv4h0I5Hed5wUfThkFOYTVwWdKCJ20l17YQV
oO898gN4RhVXaTC7KJyEg/yzqYsC1Dn/u5YuSiNG0J+v/hBaeoOq5V6pLi7MeDeT
/NEYl49UYNbNpd4tfgsevXKSrL0HC5/BHvZaeblZ4CEKlT4QlYZmBVnnm0Y1TRVk
84CWHA8KCT3hW0//nSl0aZakGMNqnJ+iliaRg/SZ3F3epkBP1iUUDnQBMpOzDOJV
qcbBVtS+EVfcez6j45L+k1g84k9XaL3ncB+Z9YafsEf0aD91lQSkXeVgy35AoQxG
otLWTcsV9wxfQM30i6GvE6xOulZsmCPxkiQtD8r0uU5bvD3zsqAqPJ2Q+8ZqSeMb
w2lvmUOlKvIVCiZnlA+XvaSTm8JjzSptFOZovwxr1onuxVIl/yOcIPkkz6r/pQTK
QaGbY956io8RfxrRxfipM796F0UqsTRKX9+htl2MS2lONWJM7F/IHJPN2uHreZbK
W2LsEY+lKBmqvqIPEmtVgFaaw9k+PZ+cdVSjrOz/hFkQc9H/8NLFvfUj3b72DPAI
mdkmPlh6QQL8zzlqg/o1Uu4kNcomEfkwDFIvtfERFFBzYENVjQ2wOs6kGhB3+Yrl
uNf4O5uBZsnGN/153G0eKPrTd+NZei3OBJW/Ar5TykdnHFjViR1HRS/UbTDVOlRa
RnUwqrgTuyLtel63mD8kMVnjZhu/GbPwPw/4kPe8rg/S3TJPU4dAdlxGcEweQZvG
NHjAyJXQcCfHcJ15lNA14g/iSYyquVQww8LtN/WZYpnMRlWS7dMDqY43prJflMkJ
DV63kP/kNacBbVEgoI2PuPTRwF/mZlM8Swj+BkYSNLplqMyfEP0Jd+7fO80P+bZT
zCVlhOqd2eG0j7CI+fizXyLehbDqA7rB0g98mr59pfi0TsAsvN6frDUVI963xEgk
+SmKrQ2ASGPMKR4zdZX55onIv5+YS/pT9ZA6CkcsDwwU0LPVlMIh5qDfHotm3dYe
iKrMWjfF53bB6w7bKMtBD5ToT3ZJ7aHDil107lsD+7md/eYQCnlex1gH2jUZRRoT
9uk29s2+ky0d8BMb5npPZfGnbyNHJV+CE1lAlWh6H1yUJWHuTViOekp6q4ld4kg4
dBIQTWFkY02t16xQsVTY3meQVujZEiJtMxiQDA+yJQ2e7lRfhPj9zaIIBiL8KXEY
Z+k6sPGVOYEZSWQalz1szniT5ubqSErRYf36+y+OpqP/sCjYozmLmTJurEc3b3J9
CLmzpx4buCzUjyjH9+M+w05GP/ikHmUX3sJMUlI/6HYQoRX/5ueduh17o/GSDISD
rPcY/s1N6VOD7p0FyOJTh3+RnguKF22Z+w/ThkVaZ76pgN20U1kYqyLhBHqZyzl7
LqVYuPRVSOkfqT3FBdfjMKo44qPMcYultSzRvudqeArEI+ZOUmzf6rSzKwn0408f
WkUMN5yuQunD40y28+KnseaMQAX8iCjr4DzaZf63HbiEabGFTM39UDSBWEZUKVWX
xk3GK1gyY7cdkugyOgxQsR9IEJhA42wgJO4lxJpsDzaKdS62BifwV+wDQ5olCxrQ
OJpBoDNRrNS1rIitlu6iBW8asl+iYJtHOPB6a834/fA4rZrxNLhhkrP9z9ilNVJb
3+8vtSbPRoVJ3xbsMxPxbyFOQus7fsoVTmXkeMLrGqu8nuXgHPvTfeYcAxoYOTgk
lYGLc16lIRvDdXl8WKqtFOakU6YK/5nDBKvqWnQJNXyoIWzdnxOMBepd2HO4qd8o
vBzQS6kVXwgZNFA5axjlpgwm7mvz+5BDIW8wQlBB5y8gGwc3EXwjFmmj0WAWTAhg
TNGiCZx3bLXTK0TfSrPNlsuFkBCHKrAYpzcWPrU2FnzAc0psNpmEJebu/wY4cIfG
Y4LRrYE5DIq00SGO8AIHRyNkkX5XOB0NHS73kmCJNql2YdyGZSaGdNX3uNEE89xP
zkfYMsk9PzK1OndNjevmQNmNP8UeL06QWR4YHe1Y6wVthPrseDt4qUp4KjjTzwU0
BsQZxkcpWDf/16bjAzFEgeh/BP41KQOuvS7xk7lxBLqnxPmWjCEbRJal4I4sfK8U
2nMAi2eF3iqke+Z0ln9SvAeqEcG9PDuz9lW9uM3O4kpLqAD1hllCqDs6/AvVfDFR
kYcx8Bqw2SDRVqXF1edB50LEaSHEzOAwkyuRPHNYXKwo69+jOiBcto2wsocyUCOA
oMiEhx1JwFqHqh66v+aZFCFbBoJ0MTW7zHY6SwSFVe24abHNQWgTRKDJIDmw87qC
nYBLltPYmj3QoIDRrIjd0RNgSXKAtnmYhepKNVarz/03+Kn5sf8ouI6T0ZKSolIW
Y/zGu4noZ2AH8AZFZj/ki4myhC2MVlfIFvqJuhtDbqfVxY7W/dO1L7WLtRtfTGXw
2oO3H0Ak+cNO8egc4HbvaetMYsorue6BhHZJgzIbokKNCkul9Z3uIEbWlOsJ8WNU
mBK8ImgIIjL4F9MbCAY3s/sI4N8+u3sUmN5hrXE6IyYAuYno4ubTf4cGxtQ8jwHK
7G5uBtH++osftT+TGAydxfloXLjPZIyqnnAn2uechwDcxJ9fxjaMbOm7hY3w/fm5
Oxcaurv423inkHDrD8HoM72goNDsjH7s5XPMDuUkEYgE6jLgZAz9xoyZk3NGvw0G
Bf440xwaIUh19Oe1b//V3Nm5X9vtJFzclXFVdBZ1VX0U+qsZ6Pzj9hUYqhlDIeMv
qDE9rCy8kNmEBocmE/OUKbF8vut5gxv9W8NDbvN27tPxYr8Bw29+T6JJhS938ugT
GVdEtnqnMShxGiBmsEB1KVGPToezhZSXLDhW7xWOS7PXH0NzIooORaqWPGSCluNg
nc4nCyW+O7NbIpiorATvNEqpT3ocP+DeES2oEg8CRZvAfIq7AZuslIIOKY0c4+pt
+/SnvOxoMlE2diVn7377et+bjcYIVWC6tZmW01SBA0sO6Gcb0ZRd5PQFI2O4VcOu
OjEcM7CKvFvjfQRBBv3shLKYeQSPpfkBNCrbHKnKuOGSOhhYnCJwI79bv0sOypVO
O56MRqkf1Wm3GOgiHX98PfK7A+tXwO7LTapXQ3Q3UelW7Os9S+jQnHmtPZ95BNJb
o2iO7H5fEEAIgvGvnvQYNWPDyZOZx9D2+pCHQ8JBt6QGWL0VbLQrvz3WOO4/l3Uh
pVqTc18TkoRFE17K3+rT/zf4Mr49UOup7Evzh2g97pXpeFf0X0QWxo/ntpQR7smj
4l52RF3iNGJMGdhiLvF4vfcScHXVWDgJkr6CQMIiHSEYxvWEJelVSGv2ytm3xH9K
ruVqKpfmsp3zZM5b1HNgAe1dpiZs0EAV29bUn+dVq+qstMt4RmGT2meAimZfUDO3
BkNpxlQLMOi7chzWXSWaJI2A1MXizkyK8T4oPI5XiBmK8qzKS57nJn7QruQoTlkA
asrwXFdA1+7LfJ5/PPKsstuZhkGXRPzp1cj2peZEpsKCWYf9i1CGGzIH1TFkudbq
K83IslmgueIUbrgvWjTYlWZvQEMKvTqHl9/JIJ0pMJt6yoGWqvRHfIfAhNj/R2DE
kIrieYoYnu7+GCxtLAcCm5FuiQv7nKHR0nHY3VMPRD7f+yquyULeUTDRqvd+Xyu6
/PWSV8X/h/0GCIPzRWsdZqxBt5iFIZys4cGpatf1kY1BYLUpS4xehS0QWtCyTKQ7
xfIUl7x8HmQ0nG5ZrobSx6wueU3Kk8bqqivDBdwVmfcuue/uDMaJrMYkEpvYHLkK
pq4+vhmX57Igd/z8T5f4Dp3I13WrMBbvtFO5wbl4gCc+7erNvy+hm5pDHfNvg3f/
3m85D9YF2GgLtDAI1CcAYxTCbwR9s2jr4kt2xbn+ztEn787MEJI/f00tZH7ciFhQ
rXKWQZ1ZUTw9SuHUJODiBShWDsqvtN/TEFiFadU9Z9ElfhYzBBKaIbHyz3BCDi1/
eLxmJcgnN4GsWhHV3IYK0egZzDaImTX7VoXmyG7BluB3UfZG0XpEI/xGQi0vMxST
sI11MD0EwXeMM5lEZbuvvvBrSzACsL8bOuXtIHVf4sSbD4Fj8sHQFNUhmzOK3b2p
n3P3v7Sjpacx+KqE2zzPqxjew5Oh2yac0n0QY7z5dN54U3jQVeem8NrJGy7fajnO
KLmwRzGWEPnbk2gqs6490Y79A9EsRxShhCWwhdQfFayxajU0YIRJqFkxh4uEvd50
3580LAUjZdcCkp7lqHf/BeM8xkNr8wZJpD4jzWkt4+gkaPh250/Z9Uxtm6GUmkdI
9g+iRuX+GoanSdhAet+2gFLNyYYYBHD4IZoH+juDfGNqDr2YWR7My9Md+8x3Njst
OHSGH77xet7wZiSslOM9DjXFquEQ+N2keKWDQBGwnovvMBodF0AW21boDafIxr0T
38NkALRsDW6Nu6hf8ctWL88O6KrwJKIRf+CurUrVc3BIb3fDydHjC7l4ujoliINE
KBetrbEMWOb9tmtr8gdTZNB/a6bzjrr9lCHUNDBGWiEPRukdwj1rlPhxqtUSQhef
WusarU8dB3eoy04rCrUFk1fjTOJyy1uE02O0EpCkt8KQ0X1Sbc/pv517fbsKBCGW
8AuQWD8Y8ZMrKFckroM7vEIDf6l5fQUMHwmFz/j3r55hQnmRjhsQj1xVYDn2An7G
CDQrgmtryZJ7OKR5J04xzkbbMbcgbsUzWTKvVtL4tnQI7Jpo8W0yZifnR3u2cSKy
sZ6KNa7YieoGODpD7lB0y7lF+t4t8vPqPbTkGKBvZ9fCYoRTTl950QK1Sm6frh2c
BHA01pQY9XvptxlRhPSV6tygVTNHTe5e9RYlPCt33tJGfP5mvz0CWabJi1P6ss3o
i/avwA7xkKhW66j2ZjHvz9aOO/aIM8XlWaFd7h0Sc20H/99Mlt94H8RudU/7qe+I
wcyIEoDIsik0/7i1mZ0fp5ur5ZUT1OcU6cki5B+JXrmukHv9AXcSvLlXx1lq0MxM
i1kFwttYzMRckHF9MB4bxHc1udIfu/oU0cP8oxwtLOdE9kEU+/Zz4Az+JX28WGop
0GZ7FfZ+qKPusaD1/Wwk9vlOCOjUvEGrJWk9d1MDVklS4RNMwu3rlgILhnxo1fgl
0ykuZdWZeeuGJnMkZKA1ptYFla1SRiK/QP5MGiQAN41JzzDo1WbiL9mdveBBB/21
wZm+x1aZFwFO472NPRi2Q1rFp9MXpON49gpA1/J9zcl6VmTgP4vgfZgUYnjpYElX
efCaLvfl6uPM0eo7z4QrUoHmxorn8sd0G0rDcWv9WG531jWlJ0c0RKZ/CWhogUta
WmoBtM7HPhXy/PYcj463rrVzMPHvZsW1E/o1vbcMK8fodpTe0u2lWKIv44iiujGC
jGp3xxYHew479C3WM2D2+HMo9t2NbGdSqP9ah8Zv2JTFsNiMG5qNJU5RxHyyQkOt
fkkCgin3ENPAZ4GTPvr20sXZBC3uf03uR6U3kLUwKwxPXvDy6COM/DftfQqhKkTV
MJx6HWoPiPKQdqkAdFToZ3jUQmRZqbEhxKSkVHLDbuQ+kyEg7O068fyvD7sUwQoV
Nyk0HdwigLRY6suu0HlAUsFBM3oLzX/LAPuwzV62N0+D6A1z4/EXTvY4BfojPPxs
WiiB4oc/C3zzQHbhZoidC1eZPotJ+sxpAxZF0Y2iBFE6Ujs8lnUehcs7z1Evsuy6
EfrUFa4spflB9nxNqylpVspdz7jqpmpqQzYUuduybwHgnEpCayzWZF4ENZLQZju8
l+FwmMPFvA7oV03QDxUB2mQLr4dsddbJydCGpzAmvoe0iBjLT2np/jZOCVnrTI3L
u6eEVEx29jLPi84QpU4MVxgK6T52XWpYum/nUsDA9SpjfLogbfnduif3qOEN1p/W
fjsEodxBh+0u4wu0V3N1IVunVEfONCo1HZKT1G2j+h4rz2kZQnO9gDgUvfV7O9PQ
Pheb5jEcfDhbmtXIhLL1RtOedLdjubg1a9XcU+7WKR/Ez70uT22EOlFfOav5rIZF
IXTvRto89EaZvacW105obHV3JUQgPzXoegMVVI/OXjD55S6+KAGDzbInIW6f6y1z
dEEFPKfVcHmbeCtavs9wDEKmOUIbxe+DwNlfnMNqAiBLM3kpIX/6YjLRxvlHJ2rc
0znIodNp9HUu0sTexnBCxBA3TtbWMPAGi3jwpr8GbKYKkuPxBtAYoWCNDzU0KEdL
0PJhoR0N63IsoTGuGTO6l2gs4peihcqJ2HhEIQ1CTLk0T47k6E4G4ZHcQDvOHqp2
mxQnqdpcJic8VSHy4VUxuGHts1G7v86DvmNvxJcgNWBcPjbhsoVcDt4pmwKhxya4
jElrB2vifdI9fvLDxyjx90ZtUUkR9A7g3eZm3Suy70aKKlo1yuAfzGJBTa2QXFmX
hmygyxwIqZhcfsu1LXHzsuBPYP2H8T4pQ21I1abEg5LUDPf/cuD/rrKnWc7UDVqp
EAiO2NSizmmC2RJr5kW4yP1dZ9G0ZbfIcBsUgibpyYF7TxkfC1RvJIXmnewXBuSQ
Ec1k+KoZjlZ4aIChaHsOOqhgq/tJ7kX4IZ3LgDHC/gunsdMD2oCzCIF5azYOHBkz
JYaFfQ0lNubpVvgNSqlREWYJmkMC8G5Ih+Tk6EU2+x61Cic704Iys23x4TOrE2Ef
7Af5fO4A5FA+tu4vXGmYe6fQK+j4UjG6L4w2nMcOURzkdO2AIPNX8nOFqIAM8Ad8
H88b3ON+C/NKEFFc9v6fxQ4Ee3ZWu8kKU9Pa3KxbFrG9NXcFXftMt2KAlm99kNyQ
c9OKDOFr4+YSc65OxL7I+V8fDFCvW9bpOWwLA9zQ0v4+fZsPsJThfhdry1HcK2yW
TVSZbA8NME2CfWDuJhJEBDdIXozbU7iQkSaJBR180V8Rdm4EmIZWZInQ0zpRflL6
1qOMorHpkxwyA0gO4Y0Xi2GFAXgTvJumCxeT3egAWIe05Stv8UkHSB6KdSzfqT39
LaIHUQiN/B9gl0NSt/RFNR8vRXxQqpFFaMbwJ3cskLKrRyBBvS0qZZHsKAjQ3P0I
1G/b3rtN2zrVlk2vYo6Ce2dqUMzH9HfSIbW2JnZSotAQ05wNbDn+9yASCnnC92zw
mzIX2gQKcxqP7udFMw5NqgNMWDd9CWzmWk19wp1jm1DxTlzCvA2SI0po6/ss4B/B
cOcmDVhM0NQcgTi47ueKCyZWQHq7V/hJX4U/KmSBxkYw/Wxo/hPCmINXmmQ0NsEB
bOYdd2vOYJ0cx0YGOQ5ZBoklIqFkE0BRt4JVg4zbHRRr8JPAUpdi9BME85QgDvoY
0h3R6Zs1fKJgnyv73yDS/VnkICv5wub4iD5J3a2kFJifNPxWcxKyPFSHB99IQGov
gKs3xxaaua4s8BPWst/ZQjWSdOZ3mOdYl59DIn4IdL30D9Y40yEci39ys8rhZFfa
KdrLRocBh6lFYwzWECqsYMQwnEJ7mxkM2Inox/numZZtmGGB+OdsbLmd83BTKGRV
zBh5ZImN8ccvD5eKaSY4kf7ICUz20cfzbjEkV4or/5A/DN0kW3Wr9qOUOs3I5M9W
7C4S6gNiGtDC2Z56cJWu6KpVPS/rgNB7YR/31n6VQWGT4JOAJtr1vZZdEdEbHncE
vmVMux0PlKpNJdTkSHV0MYDx1RjCSMmzjDmQRy2s9Q/2nFVqFhgOsXlsoTILCBiL
cmiPs7MzbW6vt3YqNbNmTM7fA4u34TBu8W2i2DfZ/aoUwPHs35fOq+BFQk3pWVPy
le9Qf2LIkME6hfhWrT07yp/WPWG8HUdyPik4uNSYJPnO9qHnmDyrVTKXK8ya5+8C
nFCQNxczsEFdlCrc9bflX1jyuEOaTWzwM1Dd8nTgKVU5CoE2j51ZIetq6f1fuf5B
L4tbBuot7JTbE8Ir76Mkvy1Hp0tTMMCDo2PapgBsIvwx1N6YSTzuZgm/7xuaDP5O
fQ6uO+mWJfmTAlJEhAmNyU40nr+x5dC61Fuwiegr86NkLAoHNiVNKBpvipcwLCUo
nrui/COhPUDFrPMzZPMKb6KYtOGT/vzK+3diIA4lO4oqdFhmY91SzPSsRgHT4AdT
+SMg1ufuVWmObGMTVcPk/J9y9RjgRlXND93whUU5i8ndhrtJSX757wPztBw9/Tgl
NLbWSSrT1GbQtpqQwZMwGSAgs3oQVeTpW3kpr3BLrkIMsqej0NZmQRXhpYNpfCuV
y5sVVKA5ZgSUAf0/tLTZGBVfnz9a/ZuaTe1U7DCX5h+QPh8L5Q7ywjnldgEnYj8p
rtxrn1lXEKZ4MLo7AWYxg+2db2nXKHjFKwttsjF3EQSY7rsXdDy+RPzY0IgbOUv7
KW4IZP4qlyrtdB6hIYAZZ2NY9GFxFARYgAwMYw9QI68azCs4UDI9M7eWfYkpKuIM
46ynnkDU8j7sbsdFfB5TiVx48WX9hfJCThlXpmtWnp2/m5gLIJsl+OdGVoUFFLNc
z3klJGmnai+0ax45iQvocmq/ha7dYgQvie7XWcGbQWel3JTO6BJ/xTudngO7i+3V
7smzOV3Y04xjfjwYSnhefr7Qcc/MvOu/0UwzGPx8uJrekIaMrdaztl6yYA5H4HYi
XXMYKN3oUtNLmGSqp0oKQyPqwTABn6HyRqWxrn0iZC/mh9cq37dbUoROoRaTADTr
4xfPgGkSLPFkvWMC5jyduasLffzk03K5xQ4bkVndfcQra6+wB7/J4yxPsP20sxnk
qqGCwHMDXRmxJ0Vm1eMhL+kKBl7W2oZEg5dzv2vuX42GZQS9oIdvrLqhcZd+STyn
EZkCbUj3fy28rL2siY8nvpLUZl7PePfBVyBOvixQrZwS2vRlvjSIdpB35w8bAeJK
QYePIeDl/ov26zs4L74JQ4eaSngCtla3c9GKyyrt/BLS4FcHpkOjctl4d8MlQcjQ
tcmBQLwYOT7es5mCal/NdOnSAGRTCkmmxuvvpFnpXL9GWQjY45rArDcfMw7ASamR
j0S5CfQwglwbPymWHi1fPvAKwLl6NUPaRfrjpppbclbm7/+0dYuvQsax1iOJKEMx
ZqKJG4sUMJttHi1uQXHZfYdD0I1uYDhKlsYx0Nj5SpsflytJy76NWHB16DgQHcxV
P+rhSnAp8VGqKxcYAf7yQ1AkpsdrEQDB1HXZQxbXFUeRtnQfA1Dv17ZkLTt+EVIl
Pq/qCwAtN5+4PEPzJOhd8hFGPN38t4LVfkaVHR1bDUwaXHf1NPOpA1Fzef54aheJ
pOiDxSd7EtgQiGMcfRwnYXh+4ibE2rsE0z8lKJTtHPHjM0aiJh9al3fZVKoLtPHo
ewboJvAtJIZf1IzZitPtUyRWZY3mddPzzZU/g4F0HSEptaZYxqO164GfF0vX2Svh
UEm1ZJrce85P07arV+PKgGB5NyRHzcNSYTdwvDnFPmhanP/iOY3haElqSLHb7/+f
vFvHnutdrUbmC2dExGx3bDpauyKBT5Sjw6syFgzQU55hD9giohIHFWt/EYJSTIcN
LhJIPohuE0ar5kEskxc0GVPiujGYGQcIG9xVUgVL+jAme3FBh3sn9s/XGCSXq06O
2naaVw36fw4P+fKzeKJkL3iRAl3zTFWbuH99gZTNRU/El0oXnjBDB5v8XS0QC2Se
eomNN0eAJrA7d8wXE48Jnl3la6sN3Pbp/kP1sf9D9/L3OC+Ay9d3awr6GTJFrXKi
7ZOo6oxzbvLJLDhsFj1Bu+WoJzw7KFyTRQAeag0afJHIXdYpgd3tmJigDdQAGxhk
vZNjchMCq7adtL9i42UOVnkWHR9eE5o4NmDdFlfiBeUhmi0nbrp3db5lkZiviWjP
Irk+BBNX9ct2v3eCt/sIC7bVfGK17FSyGKmsvYEpcSG+n246ziVJKd1xilLvDS5K
PRaOBrOpcPMEeur8ocVr9QUOXd/YgWkehIj/p0OFI/N+kiUJ2wc1xMoOM6ReZOAF
8UOBTlm/g+sCpmnG/VCI9lnrs2fV0P6B3VubGBqvMJSnYGFEFY/4C8YLDicbaqh+
IbEBY2rOXNOrC+ip3bhISrkhRA/MOy5Wr+9Cbukvvnok7/hvfdqcNBdlW1/ZfFhX
A1dh3Q6QX9m0/IQpXTiZJP+ISQywmo5hXe71mLHUVRZa2Tv85/sCXBRETVT1XvJP
mk4u8uqrItVWOA6MclnXFyhVlShSinEyOnrYYT2wuqHvL0TSs8IEXgXctFSSXE3N
Jua4U2OcsZNbW32uHLXjuJErnXEmjYTHQLlsd1a1IolUm/LotTj0J1zPuXZMyxrt
dRXPUye2UeVfwAaYiuQWxfNbJ5/hDrzuxH2G7KawjaIlOqD9X1HWsq74huNQ4nXL
cIFCAhDKAl9B/S0T/NDOtFcmHsXqi/sE1jy48MKvWP0ojGt8kUn1wlZV5L08VLvB
QspHaFesiIErWWcdaVDveq9KxFdhXREtxt5yJwTUNDcUKlvHjxJeUDgNxjA8KLws
PQmQ/N8vYXh4wGC5lGT1hU2iANUMyAxwC0YeRcDuU104fauXNjjdbSb2i/OhfXac
MQPftqYP7FBm+cJDdiejr6tbNhBFYbzmYpBftfHi4MhtSZSwEdmmzlcctNmnVaGE
I0Ie7OnS4MElL+s27gCsc0Usuop74j0n9mVRrLsyBQvTjcb++He8hvy/Rtk8N9IM
gPUL8mY12Xed1WaIPlXVU4mKGpI6FdwUu/ThgZzrlEwDsy+rFX9ncV1AVQtAXhWa
xjMpTafqGd9lhe7k3K5TEeoocKQptLg01wlgQtfQ7zcvgaRXfjRZHlvvhcVqcJfk
hwI8+SQD3/sSVEra/o9+J7zElfHyl//gKG+6+F6bEvQg5IRTIC8bZLdadt6K3Xal
ah/ow3W/XhS3ILo2xlA/kthwSL4JfYykyLNlHes43lNp8cyxc8q+NI8/WrziL/Ck
v/q1xSa9LciAz7RJ7Y6liezWPHCp1hvVmRob5yXHfS0BbdzAaoCNopG0wonQL49v
rdj1w6N7d70/H6o3UKJxa8MFo28hQn7F8PAAntWQT3u3lOAsNux5aCI77/3FrCOZ
zNGtuPhCELSglhjN2UeaIJ2kkDgC7ugU004RvXiLfloO5MxEyg93wQW302S2A+J0
fBE2hfS9StKCPlOGP2l9lKkopcuX8yPhRankJ6kSnAU2Khv85o06eKU4AhNN7B2s
6/qOnLeXl0ReYb6rDo5w+YeDb3z1bLxtOSz4Bwcx2PcMcIjDy548jZKjM0bTk2Kv
RtH6IPY/iak1nZ8dlX9uqC39qNMpVbXAIsoBG+NfnrolVHOj1O1P6P7OCSgj9+ou
mY+Y5QlqyFuSBNxXQ57tn42ivqd9SKyfNQD/Oob1W49pbRjrgjPsKnJ/TqtAPuMi
wnG/dG8Nl7t/Ho0RDeYnQWBX6+6gPtUhDpcuVem/4BeYiSWj3RlQzjQaL6rTsMJR
7+Dpgu3ShHAoSrNCzZ4iRwiMKIA2tlJofnSuwnhA4+NTVOre9yPZ0feTBUp/uq7Q
Mb+DxvfW+26IHcS7GSePUY5X31k2xkYhMtDQNTQLGBge5/FYXnw3CG2hMHZuaQrD
8CyxvIDpwt5ZRCTJeGsy4krF4LOJp2fxUkswYNz2nMX0fnqV+I3G5djOe1P9/usm
06ROEBq9TipdbOfa3p9jtdJHaT6ZSMOeYJqUuAwoh9ilDU5PUcqiIjSV0YHYMjro
BnjxgS92YF1tyc3ZA/0HdEOdQ/hTulWxXZDCmWO5cy+tZKdMIUukHwECnGgBST7k
eAnNjCOY0IW+QnIkZ3Lhyc96cTxacirPyUtvwALxb2tvGlJQb3M+SQW/5Ys3ZqSM
bNHYIaN9PIPVKQ0UB+2HINMqAf0+M1qqQGXtc2ilrZS+m+xETdgY8fMZQT2lJxMu
iJMv7aYT40AWx4iZCBoZcniYQ/mewmuuxeDr4KkADy/9j3/785vNy+e+CTVHRPBZ
eoGLu/KXmqSmJi9yLZlq5IZEv9Z4w8Y+dP3lMxnMqPDZ89GcPMuCJlv10LY2e4l4
lLvukkWV7Ptin98bgB3wXMoFy9Acn7CY0yya4JD01XmX73kWKIfR6JSbsNQ8HUh6
qdwcOCBVjHvcfxaY6NkshknWWHRdRwJnvNLnPPaqOZjeclr6K8lPwaQ9jpx2LHPO
qMqtb6n7j2f/bLjw50yaBWI25llBtTRVaEu4VRzT5GTdo7QyagqT0O1D3q7faq4i
WCLKrbr/uBlcW0KpEMnPLWRtk20Lb1sqAUJNeK3AS+JkgK+c9RbF3ZQiazY5SWyP
Uforoh2mrWSGGTBb8bG8SA3uvAdxCpe7LnFlO4/Aonl7r2WuHV3rkiTG27AoETgm
fmIX1jgSBnQtoJx0xLCeHpEoCfPtsjXXQQJ0LvloB50huRP1+ZbAeo9r2DIUe6PX
E8qV1NHeT1f1lqNTxicO0A9PU2PvgDmNtbTeYL0MSYmKpVTS7JrjCqnGwsIlzam5
xMGNfNFMcVx6iYPRJlWOYTExlTWhSv3suQrVIu3WphPj/KhXApDtLEOyUYucmtNu
3yA4zzqkIiD+5fhHytGtskGvNxdYo9mtVgX6G/7ZAiHqm+TzuhXTLv4OjKPD4N8q
szu65yReAyXul+c0miWWndL2OQZ2eli0EJjN00JfxfIus5X3vO8J5xRpq73GsN+3
n1HqRVXsD48C8i6xXg3Z+1KjPchYDg1IWUcHwiUDAkWmz/gyYfRaRVqlDuDl3cwH
2E5YJJJSeumn9ejxKFScNCqpdzuV5oVGhyeklEd8DTPoTTUad0fLZh2hG4xTQqED
RgQnVPHZw3Nt7xt4PuXqeQxNNfIjXooJ5IJCDHbrRP9QZmhgVBoASYtRobL3ewOE
fU+c4t60zhUHHxA6jAX3Iw0DIiu4e7xR/wicN1/uxlgRPop50pk8wYaHWVp5LLI0
pzEhz3ov1vxbM8BA9nOVzHPhfkzf1a1Nny35RBIqP8Hi2xIvUIJW28j4oNJ0zOEE
C4AVFDZRfNFSujKgArVMehV/ItyFT9gBemZfO2XrNGVhYxZQl/uUXKwnip7YYfQ3
eRYlhNsgWwAK/ACS4mhsxsYIYta1f+4joI8HS63CdzhH/nduugL35L+Iysid4ebM
kDWAISjSiyhlm2ey8i/V9WPElkE6oxj72sn7nrmDEufyqrpA11vYfjgbNfYohgGl
JwrdbYHjaIUCTj8DM/65BMuWRTEgjhT6/rSaQ5j4GDYZ41rmTLalt96QP/M6Gdl/
qxphQ2ZWGjDzknj7pGuH2PDJXb3EsbIZ1HJd4XnN69lJ/flB6G7AM48TlltsIhnC
WWowyQEsjJtxMEXPhY91XfGd42DdybfbKcxBiOGM5a1kYcyqfg0JpPKQMugd87BY
fWyJ6QzcSb0jGDOm8Yded9OIMdyQzag+2B0Btx4GuoHKNO/ncilL3eDCIzNkX1Hw
hqVRxuDxqKAztoxSJ8Jp6pwuZZxwp7evOZthexRpXrpdBANE8RR15Eiu4QiagKqZ
BHnj2TmMVyNE8cugS821VLtlZOPcc4kSF7vsamKnaXgn9UPFJaMoB0IjXiJKkGMw
DBM82aHHAyWjunyqUmZBJ1xwmDn1ysxjLl/XjKcXnURqtIgIKLNjlHadedaNySUc
eVKKWZ2Z3MaZnEWel3jUo2USrPcyeJMGRMradiUBYGXfR3uFg6vEMsFv44UQnrv0
7gxVxpZBjXalLwsdcX3Za4X0KJwpIzqAF20cb+Ts/2dC9x/wFHTOTXj+JSpHJmDp
82UMaUvPVjaeux1pD1OiwUrG13AOdrTDsSgz69vYOqly94CxFaU0wIf72hd7JxOO
yvZSNUfFKMLo5l5rAfbfWQlfFLE/5ivh6hIJfRyo8IdgXHLUUVDE30wZxmHpeRgT
GoAP4cr8CkJhwgFM9gbIQNVaZX/upUSM4roxUSTr2h/JGbxgFPmPpquJkdKr2Bmc
IIULjpxOmGto+mk5RRF/LswsdEr6I4w+77WSG3AyKE6D7vIpjxqcxpgYqZP3HVJV
H6bSZLO7dpuJ8z1PjbgXCAEY2GYQhVVacqFk6l4z2O5p/JX5yEFDG3Fk1F//Jpjw
Y3EpAHssEzOP2ga72/EjVnC+9aD/NRwv2g92ndc5+AhPmtUXS59x1WviKDsbmJoY
KIVxxqcY5bLfJXsL1/MpVC8+pGHIWWqm+n13MmH2j2s9bC+cVia5FIM08V3Vd+nB
sf++tlaWZPckkvrP4sxTVO8bYfEdCQcispWRvC/zoi1UPl1f1N6Xd6+HOm67Hy9N
WjPd1kA8gJY+6TrqRW3ajWW+tl2dgiK9ci2xl2UNP/6z+vPpB+OxPu/PpXMbrAnW
4+qCEF2O49ndGdcv1TEQPeD81ixIbXEZorLXofyNZRb3DCdE2xGITYqNBZSPLjWL
DV7hVwXjqb2HlkTJRFGs1LenmYySaYlS7nsEwYno2bjtcTBAuNCFwASCKz+sJP8u
Xm5HxkOPdcvk0h+JqIPnIp+q1zPSC2zbR8lwbq5dRr77O0jnzmQI2jhOO5iXFWFG
nPb/xmjGd19EhJhQkylVRiL92kG+2mdFGKpgrTmpuj/0bVrA3y2518usHee79iyP
n1o3YZZw7gNOt6F2FVrXV6dtjyKnr4EiYTzjnkA0c/cWWyMtcSPqSwDTBQtDW0iS
g2cgoa8A5Kcb8W1ntOhnqeQk7zxOFDGVwlljvx7aYfoc++4dYG2q9WrOq5Udc8wO
ny8kLj+vrfJlqLEMK5lq4Vp6QcdXjA1bUgnZ/MyFT9yCAvxJ6xDP4lm2MTjWwCva
nMu7wklQJKDKSZBQQwR4w4CvQrJFC67RnW/9lu4HXTmN3N56YYLDsD08WYq44ME5
0vW1nkk/ffzYpQgWktmfo1X8aju2n5pJ4K5wNFNN8LKUpIHwm2OCozcU/WEri/1x
37vOv4f2RVVI2c7+p1FtbkneubTknBeUHdzqVt3Y8fpFnCOX6FPwf8LHpDa2oY8z
ihhR7e/jXRvbk4ZrEgRy7sPBDdyQFopsDVD8Fh8xRQlZtwnlPJaQt94ij5CoRk82
f63BEjs4sEJtP5OmQfGlr98L1YdYIWwLZnCAzis1wK+my2zu3mSM79U2fl4XmIA0
s3C4tkGhksD3sPRtC+Q1WYGg+gBYeir0a6NChe1mlK5X2cu+itblgmYF48NG2du+
B+3LGXoXGOsOlZmzOzG8Ww0KgYq4kO3QFkYlT/M+Cy0EJ8VNPv9drLhVjjpdooX0
C5QapbNmAo8RMOsI2NK22AjmVZOIhILUxQYVSD8ilgmam8m3W/oRB6kEy07ZpMyT
rsYFEbOk49HdPk4Uq9VYEDM5ivzshPZQNYnDeCd4RakICAsoPwwZtdaO7m/9iqQt
GvSE5Jf6HpxCZoEGU0G11WTuysu/QCWBpK30d7vBLB6bNykxqLsGWa6xlyXeQqjx
RMQaFuHk3UEsQAjc9ciC6JV9gu2XUnZht6LQ06Ubm+Ag+3UA1UdySMVAcjw/qbqe
6EmVIBAeDyYs1xfDEnNswswxyZgHfF2ANTXnl5jONV7D+/Y+7MI9cC7vM4SfvVxI
Z0R6vu2fk4h4e/tK50oI8/DLCH6EmNSNLvd8UOMHn2AeHhAbf5a1pSu/Oy+165bv
/eCPKdicD9wh+rpi4lmheU/5Ayx6Rl4b7lvbWwC+yuiGzP40jJBiuR2f786KzDdL
TXNszSfRugZglNwW5N50EaK2XStgdBkaS7eJlfN+Z7KXsJ9CFVIf5H+eh+TYQH3Q
5K31OD+LZh0W8M9k5AWSSjPlsG2DeEeO40y+yw5sdUmM0p/5sSnJlvPPExLysrwG
qnJV4cZBfUnWsTHz6TbBwDTqDINJNAHEUvteWnLUTp9OowyJpGG1heuzLnvt16UU
N+NA6egQDzyVYI1X6lRFlxOcleP1jmprS4x1xZmT29u8IAeWdW6JkBV+MEY1SNLH
Lam30p7yI5M0KnNXPjFmYoiCeNpw1y08Tg5cp1JzaEyIQxEg2hcl0JbcZbCQ4thJ
5jUG/vO3iUIp72wb7DHleRnJX9SDzZebAznIg2I/049wYfBBDAPZXLTLNwF/6sdQ
yUVhr2GTIM+V1rOl2I4E29h8u+gEEZGjcSuh2F5dEFWcwrkc+LlWYHoAcPET+J2i
K23bor6llmz4v1qpm9/48T1xE/t/cOhNIB/nizAMravBHW02kCK+TgWw6a2qGz04
BpVhI6eCWCGyyOL8RkojTSwmhfmNQANqSYJB6hr1J2ls1xF793CVojFXco6Xe+l1
rZvIA7Rh9Ld5TOSTJYk3nuMn6AdPYWJcMFcQSTeDbRt1x4Fwbwqqv0uChBRw2Vn9
7UIQPpOw+7DqJwO2NT/LlOO5bovyGtj3jwy9z3j8h0jdL/AMUSz2afftavaMIORx
5NRNMlpminEKRyJW7YzkddS4FmsKZYfHkIscjpXJ8WiJ4DlVWd01FBfMC7xUOvl8
GSrFad5XQ5EkoyQdP7kSayIZ2Onzj+oZlhXayQOZ95YfkHSS92fK2QRz0FQP2kIg
1ZUvHCkPYP+kEyKHFbadGCGpc0bEUg8m6U9FPs1RojNiamxtw9UGTn5st4SbzY/n
jGSs+PSdj2Z2QsJpRqv4tvfiJqij+yQVoChc7FqgSJBGiq+oiDV4VqfxWQ4pwMZ/
jzyI10fanA4Cxj0MZm51FuTUr+PyH0kxnZkYnN2gH+vyH2H3O87271O9Fief5lfX
cHYlIiMT2qC51acjiiT0H1/PIEpNh9OMdvf5HEC0/G5vROFwwmoTXTYazY/3D2wF
0FtxJaPG/n8Dn4XoC8lbDBhz/1SoqDx0gpvjpQEDUqfb2GN9uGLffM7FE//yVGfo
XW+ejm7y/PDE6nWirmHd+gIr8Ql6sxjEd7jZR6fY9pnIUJvozddKcWLxp2NDdAGS
6/n2to7OJXpRS5GO8/TfWGx7QDBET5bTlKGvJivIgjsOOVFuhYohmQIgV3Gplemq
myK+k81nF08hJM3/xTgAXZkDWkP5BS2UOolI0+P9+pyiLdpMiLtpy+EbbcMau3eT
1TB0Oz+H5t2+n3H2Pgg4ozZBVi+W65IfwwQCM1zIfQbK4AWpjpbUFYizlZ03OBf8
LwSfw0fpS8IEO2Nu1kueTnUWXYbqcmbeUgDcIDIaH8tlkZILdfbyEgPDvrjczV6k
t+JUsyOGpaBVEKQ131yNnh4rsCJlu5AxegA9AxkVAxZhVrzdb/XoEzhYgXwZNCyq
2d2ODO787b7NSsAyay0/rmjbJusmsVuBQtEzLkvO+7DKEQcBMozw33i/SMgcAVJq
YFIIZE/cJ9fE7yN/bVzPy4NPSOks8BIMLjiiOLdzbKTrL+R/ZEb8L3jKay4zKsgw
3Ue3e9GCHso8mbx9jKYBJWDMWIEYxNxIkEw4AknMG1rNE3a8CDLQ+WAQ0M5TR33d
KIKVm5pXvqEp2pUeyGh+p9QI7tzUFHBrwP/oRkOr/sQZ8HzXUiTgyLHQ2zuJ3R7A
Jgg9bCeQeZqa9iAvLgTgLHed8GKE9tKKiKbU5LNIxrkY2AQrSPvCfopQEasnErXs
R4Nnjr1RmPUDbz1IToqsuhXCD0RzKJj9cTw7kmQOYmm6nxXomMLoJ/eVuG6nIOQH
/w/GeN+E+RCGXMfhfABY0Uc0l80vKqhBlyW1vcihYjEzM//cA7/6qV1BWrigGC+H
hA7N9vgk0KCeMkJRZq7+j+v3NLiAitd9ygxmBI2gAggNtvEBKfsLnLVvPN3/DpWn
im++OVvyQ7tvMbqA151UMRfcA4Tu31ZJIInr4E843Rp6DiEqWEYFIM2xfUs9q5i4
KIEvjR4ZSma00oT+8Z1fPQsR6kIgTjsOzGS372BNEGHl10qVlgxF+qXxLjp+Yzcu
ba3eeGMjPTckhYVb+JJOR6VB2WM7o3XVqSW0eBxBPnZsTlh99cROzR0CDkuGFrFV
X2dKkhMb5f6sxhcX58gx9drDTw97mrklCowdjwTaIMTBuTvdm3WnSJGaljDuy/YF
tU2f+1Nvkh+2r9Le8VEBXEyiGgx91+pKFPuOPIm9ea2GUjUNe/HQbrZL8zJ/jzsR
UeTel/fahPh7hJ9Cg3tOPVNFUZgnrOPnV4wrwJa3Wsx/3Owrg3ElsMVBAzOiUUss
kritd2hDX0Q8OhKV2E4YH2JditLV4P2Si6CrwtDpP+i5fzH+QhBwFetw2C/7kLuB
rNRoFkeN99txtX4BcLfR8UjKnXB0nrrjS8Q8demgEZ7CtHBe5cWdNdPafas5j/z0
nXPqTq4KEOrIu3phQ9k/sEcV53xj5ZehvMRLeW8HoTVVtmtCFzCTCnnBcqtKt/ap
UgQ3juUx67K9aGJPnad/JJtraSZSUKYwCWfthOL2D8L363zMpocfN8U4/58iFQyQ
9metRnfHE8CHLams1ilO5C90DkyfbgvnJX8uvizpmMzhtq9kCzKvsjquwp5aLzL3
tQu2mvjZ/5U1jk1/3Bhm4gigtrxHjDZj/1PQL0YzL2yjzdcjHr1urMIWyTGSXQmx
bioaqjMNZHjyihUAkkgWFR6RWVQ8ai1hru3MDH1h9az8NALD0djwii1o2lIJmLtK
XhhJtolSfsRYZD013QysE5XsMhKd9sR7qVVTeJmG5cqYzvQBXIeZG/jBg6rW7VKM
4MkOmsQMfYqV3nDmue7/fGvZeMYSLP8zeeP7DhidT5dkaWnQXxTkh05cjwiCv/RW
Ek8B5FPIpm0LBPbXJyF+fTiZhjNRfzfKfXDIrq9+diLht35/0uIeGRg1STVIXN01
k34e+AHMnUA3b3SKN40xzwBOYb3YJvRzlp7V+4tOmdnXcvjBlfzljXDLi1twmZzs
XXAfh1tfxk1BzaP78lbvE8eYBLdvpZEJcmxvBA+cRc6xX4k1VIo/5lCHVmJKluJ9
unn8luw2CDBPTdaWH2iUeknEmGQ3GBWS9najK2nBQ+JOXNlSHIm5riYW+0GueshJ
gSQOzCRqJqayoLvD946wvBd6l7uqYuU2ujS99iT6sfhrjfGdi2fuHbB9WSp8DiVv
cLH8D1bPx79YGSLjMZe4ARXWOGIMq2e1MsHMboiQCj8XOcw2HopoB8ohmoYsctgh
XcMdvpF06zB69tm/JrG47vvFTTftwdToDIMFrBSsYpRDGJbf0NvKTjyMNKmHmzlb
dr5Ma7+c4nlNQpPcoY4Qp/pRkVvsaTwbnrkYfGQB+H/9Vg75bvClEs8Tmz4Cnx5Y
KxBZCabroeXbfU/9dmBo45g2E+pYYg3+6h+Wc2F5ueWnnnqT7bzzwTiicjtVtYmn
ZpXrRf7AQJtoNg6XTRYSw3ArEa52SlMMT8wmbtyBXntjlW4biSjQp8zZRIYvdBZe
jJzsopW3DhVTdSQ9ya17/C1uv4HFBp4+mXi4ERpvvtvCkWZub8pVCiAG9cn9/kaq
rzoskAG5IUsX/+5hgHn86CejsK2diqqTgIBYMqIyDUbwBpZoT7jQRJUKxlaPO8cQ
8y+BKZhQGsATFXhlfJ83RFrZ4KQ4WYDLw2hbLbOMfP1+5K+w+pORIT9zkV1XSkd5
xC66TTB5vXMD8h7SXGrqyMElIVdxfQ/1Vvs3Bbi3QVl6GA/+Ws/PTfry4G+efnwm
dpngDaFWYYWqnTAK6EzPInYT1EYUlsEm34UPTsj1focF0GVGJpY94sH3SxAWbfOC
qUFI4q44U2ImRk2UoB2H/KSQTuvjxZHVa9iqaV7/DLqmWq26ytkpuGiUzMJrrx5K
KFyU4pUa6KYGiBk6MxE+o5LAXnNKLzNWALReNK21wCaxGLOoH5QsSwBGbP1BabZs
DjMwvvvhhxlZNrmxTLuQ7JUWTvZ5Lo3jiAxfxJ6peNN0k3725E4+nizbZLxpLLko
DJQBV0+5jR5noqvMGk+O0D0HM9DXJepoMkDUY/xJdEgABTlDvhxdtLJYiUih4AIv
4/LqwROYDVOoeKnoOitOxVUJu57gT7Iw4WvbdcoqqEpJjovAC3PkRs/PI3AKNTES
XsDXvB3ezQ6iGwqchK3S0bb9EPlLy/Gj7fNYsnAdD/UGyc66Ao2bC3i++6JY6MPO
ExJS3H+7iyb/x/wOEVqBtkFcalRQtHpip7Jb8t6aS4cnDCzV5NNlyuwMxnp3Mmv7
1zE0sn7Y438rgEQHr1m2bN+HoFpqGEUzHwS424K+R9bFKeJR/akY7rpdv5YjNCRR
pGSft3dvnFOeA0YwENy3u6ijvwsKjceiL8CWumgnzXeBbZ4QSVyltlC15hxHpiUL
nTjfLJpWeSQY0fJOVl+rgUKlTxEygyn5VWvfv7gkpQOf+0dA5SBSP/Nl2jU0K9uR
LUiXyk6/aUVppykOpUFC39k0v++t1gk30MBBKotiY52m+YQObhoajuZ4Z/rmmsuc
+ITYCYnpBWqS/YQ6wra90iSdFam0lhnn/4oGZyf2+jtVg13S2a+m+MNtE0/dF+nk
cxmgafRC2qF2rtJ0pD1Ci2E7t5P4glWJ/W7N9zz7eNI5jijKZIMhu4f03Y0dZdTx
Ic9ALV1wF9auIhONch3pIviSjVoU3NKi9XCqdXO9ecuXiZzXdHBYhN8PQgLA9tbE
JBs9PbF/9UZdG9grKmAqCHsv8hXikbMoonFL9k/jO8PUlARCn3VK2XNunsx299i2
7v/Zl/2bYvV2SUU/xD7b7cpVvRQJZe0oK8Ib5lLc26Kdjocfm1D0rjJTochJwSHY
jUbaSUeiDsbDYP9ozZ/xDHqG402IjiHW3A1rQ9r7OKPAoHVZEkGPXxQzRn1YfRYi
Ag/wpjGn8nbELMmviVTfjEiml370TeqLCBW9NWmJly5LPxf96wMXwv08acRTkLaz
73IKmZY6QBWgEfQ9geGyQwOE8xscTGJWRxt2aHSwM4x10i4Cq8EZ/x1ujo9cO/Ew
ezI5maPpkVXa3S0YTHfV24eb7poPPZGpKW0SnREz23OSUuumPXEh/CNhARk44jBL
pkdSKqfDt27DhGtharKfeHGAYNBIznYO95p6jAzDfz1f3jEMVetTrx+7X2KDYgC6
j7hJpLWQsbytBQRjMaj1PPSXVN3uerKSGusKMNPlqDyDPv3sTZVXp0+zEdDefzEp
KX2ccDYzfCyYmguY3/nMuS717n/6CVh1SlsOBoCsZg2cWQnM2ASlez1bjOO5iXR5
jtXLjy1AT3RPj+lMIZt8yPjweTFKwtQM8P5nWKrfdhT55qxM/1Yzt+ePqv+GXZGV
haTt++Zxp0nS/aznXQp5yedu1FCYzBfnv6TN28YnRljOoB1j0218yurbuFkgXlh+
t+TQYhABxi9+DLWDrf/CzpfEBEs23JZHdvEGhObbOCG+M8JjayXynGQEXKDda0y+
RDv8Yxe/M10TdUKUseSTiPTgpWqyRAuGiK3J1nPuXQfQwl6fpen2LzNPuFLRJl7H
JPB4isBPQJw+9/uJ/pdDZYjlGBklATu7qQYP24HOFyQHKWwilJ6qmyBmG5Qe7Wz0
8LGADJLkIqKV0ivqTaMpPatFx3QNW2A1ZTBkIaRU3Xotvp5VdacBrT2Nf7JDL34l
EJ5W1ZfOI/gKiA5Ulf7sEJvZJLNgjx+/Mjc9o4NnQn4VCvoUqkMDwNNzP/Gg6Pgm
375DWH6dOXhPapVUbQmrsh8wJeIHdJCdPV9xIqVbRdKA/UcyLwvFqWJZDYUNoL2m
nzJiTHt546M7ZphaMFUsKaE0AhiIyAR6Slc2iG2xTysBePhd65i0h7aXsedLvaY9
+G+wyCAjzYI9MTTqqFQDU9RAdZjd+WqU2kKeHVK3XyK5t9jVPMZgDhfV8hcieyMB
VnDiSq7rgH6psVS9gvwR42G2t2+wQIrp5OP6fs0z3j2Vq0F3zbq3w5DA5zbN9kBU
zLKZJoav0ATdy5ltWDZW4tPscG9Wzpc/bHKjbyQfyhSpMAl9+wXCXPLhwu/XST+W
jIvonkZjo61nltLs65eL7DAMSyahl5zPWP7Xscnab+Lp+PxbVzOpkaLlqjoANTsM
JQ3tSFjBVgzSNnMZBa0/G37+nLVgKXlT+TvDYFur0EkoHo8kCLLw+EvidyJD2gfd
tdB5olyftd9vhzhXnF2ROuSrIaC1si9yfdt0PjJl2gmaadee59yPUs9v/g5KZwrZ
to2wsoxpTbA96mpnsi5KQ+nlDp1AjqAXy0B7kn+iIC5gQhTDQZtkhnG2PkZC3uEL
zbw2hZwjr5uJCfRpRJyw00wKa3NCzrsg0EgXs92DH7E2u4AWMitNdlk1hPfDD4/E
qw2Yvwovc7cwmTbt6qjvTcn5CC90AiQYQPqdzeiRfPH5R87ZP+aVpXvS9s9REeUB
ynBjPJ8x9v6wy4h67YGU5iIRhzvZa31SB9zboD3Z5Nr4Oc4tY86Com2g9b1tsJ9+
DLXNpMYSH22kRDevESvEtmy86MfT6JEYmP+vcjDbcgzZVqTdoApZrdePiRgI88Pw
+dCTyg9agtHJSyoPMZ9VJ7RHFEFaGTdL8SopyKqR1AT58Qp79c5HFL/Om+YNq12W
uEZizyja9YVHBHpTQuasInPpa3gdaH6NT5WClHwqR5iZWLOQs+9T0brCkN5D66tP
g5PYmfg1jQFCPhJiogAWkwrx5WEno4LvgC2PtOFlEPkdb9XpYoYKSWi3C8MJyZPL
RHpC3QTjiBxIMJv8fzo95cxbdG17mwHrJO89OHzcLNJFYtUvhIKqn7m3CA/tUBDR
4ZKJgN/EjBDcx899hdfCfytpt5N5lrPrDCImhmtfwA/9/vJabPhV4pGSfeJLRDx6
qFxrG098CRR6LuEvlq6RSBE5EbcRhWXi2Y3D+rtlDr4oWIXEcj9Eu6Q9nDCJyqTW
UNGfX+iuGBHQYSOM8w32g6fezPcJPcTvlSIKYdfQNzvIcI4m+Cv1zMhnpqp1ORzs
AaffkFal8jvaI5R8WvnvWxF8S6mz7mEy8/JEqPCwGcKzOd3gCY7bIN+a0Hl50isB
E4Vqvz5bFhzeZzMyVyUG65a0En/8HuAVyCM78uX+IvOs1Iymq/8V/mNGspdYrgpe
QzBJMbENU0YypPCTJxc0sCsY3ZOUeZgIl6qqJxLaywltarSlS8hgg15evfOHv6zG
uI1430MT5gMt2N75g0jFbqSulVEH26khH7H2W+rlqgjCTB+DcPBGCkW9rkKE97gM
ylHs33j3M58CSq3e5eWsbqGe0hD2slhL5OGYE7WKAVbMu/2PKLP6+FoQSoX0b8rs
M4paQ1JqLsY9jvSXYh36NS/EdAYYn6cFoXl32rgJrU/dNW33+ITaxm1JUz67rI8C
46EXWx6lTt2FLDMTLx4t8CxkRn3f7d8Vp5dfpHf7LAsyzfe4R5jS4J8ccfX1HeCa
ESiiz7rU0jC1OmK4n3PIDNw9BV1ztDgFaQ5lclIg7NeqzB6iAzZHlprwEKv1J4z7
7JZcZI4z6WOJAwwf/cGBzPEkZvIH1zhRcTzR4cfhcayBYrvFRcAKHNdU9J2pCmR7
p0OZj39s1aOpWdjpUXbdz6rfHDdOWDKc82c4mmo4/Anv6gSxctrwu4UTpbZpgdwu
0yJ8RUwXtaegRg2qlNTKOlhxoseI/1KEZWk55GFRnvOP/zO3U4sf4by5vJyVxyr+
YZIeweVzwvsSsQ+vjSa9gXaVa0G8m+CpHso5eN9bgvHPkvskGTXUZBQw9BLg8Hub
QGvlAlkHoTaqMeFq8x09cldC3uHSMU70860wROqE24Er/xol5kCJiohaIZpW6CyL
9WkwYAi2a67PCX+Kjvfi1wa2gADHpKHzVv+Tg6mM8mbjNxTWgArXMWqwbnCzt7Gb
by4FyvdYLUwnB661JVqp+yz2h13uLtKx1LHroQeso4KwZo2JjLAAW25VApvhpYsN
lUeuFwOTpWNkRMmCADipYreQOqiYWrGumKpa80jHXdTSgyPX4pVWuuLjvU+OxRft
lyryJjCLqsw+9wXA282hb1kyQWhXeEpHhnyPS7SVPcvYwUEenpgpWuQJef6g3o+b
PiHkYsLRZZX+/9IuM3mtSCfAqWf9PkmAHhXfH/MWdFf44EtMdY/5gcG6dNJ/y0Hn
MZUu32905aAzRk2ezYOoIAdUtJH0KB5cXJ0CIR2x6CG4LJ7emU9429D4FQ47mS7o
MXzfbZ0sHgVDfEH37tscIUUqDOai9EVw4xvSfz4K5k9UvUJ434jOjybr0QIMUrC7
mSJtCvo0GkPyDjcTSagnVkmSBk9OvVHE7Rj8n/qEJlZ3ZH0i86/3DCT3hJe0ULhr
TMQRoH1Ci+9ZSADRIjNKqclvfCBekL8wp2bRxR4a9Y2CnZaEZCG9qx1bwM6Bx9HO
Gaa7mX+/P/41WCb3QBgvctAsIwD69C+lnIqH2NjUUPtZJh09kUxJEHq1OGQuxaz1
o9vvslFus7nRrZj95FgS+SDIhlSADT11CDX0x3ATah/flFeUDPM4BkDI9Y3gtFsy
kPMuYL+NHCs0MCeEn3a3KOR8Yr1PgOibPQDzURJqP8QaOZjwEkuDF90rnuoBxDXj
8E2Pzj+wR8Tr0YdmGdBE+Xz5aDjAlIcdhVmwywacU795bNfI12kh4pcehqb/sOG/
muLH3pnyEV81Bt/N4oA+0qCiKJKKwHXiBqHzq8C4ovRyv34+nlMCrLZO3oy829DE
KJgY5wVmedwrcMTVINU3gBGURCgntItXDt5r2hEPn6n9pDlMG4aXBDR+fJZ10kAz
xtoKQCkdpDR2gVzrCLcPfrNKyO1AMc8wKu6XRj2bPt+lTHtrPtDO1ENIg3TeYH9o
nTQqfLVAZHE2K1SnrPJXZ0FawCKHdJsqz12hklNaAd+n4YgFqQBkypTqH19nuW+u
H1lGajlTSvwIPqFXHQqGhAP3p1BTkzOX+NhCV6Lmk47BhFtVg0COUjtuBxxzoW+l
lxn51quEkr7ZxSnWPux1g/EZP9Ox+I1gVo74MRCdcODhd4wM9tS9VVQbU6AcjH/g
FSH5x/9VmO3htgQxGthBqLDzuQLVj6Z+bGqldkrOcownnpcS/VeiZSzPtZ3DQ4GT
Ik7qLr42nJFsvvVCV9sjQb/yPY6eFrtl00B7/5ne0nGcW2P5L8KkNaNOuz0QA8dA
cr8DJk5aievHCd58ppk0QfVFcHtHukhG+PTihFqZGvEx/pG4rObD82Pcv+GAUurb
4cuQduApouMCZ17OjlQskIVJAblJRer59ZUhKw9MPd5fDR1KoK3tMrpmw8RU1Opv
OjombtfRylPrpvQ/fwg9nJbe055Ygs6YYa46PcUGDnkLOQlqYioe5pMbcrsk9OZo
ciYdJSwS+TMCGXlcYqTY6Dq1fK8zjvLApwmRI+zIcRYofd1AhzIXIgWWQZyEPMaG
HY28iapGorFt23MD+uALDXHIfAcV1edfmj8EGq1e9tlAVFd3ht7OVh+AY6+djQIf
MEl2WpCyZJNgbXzD/znpz/7Hm2ohaJOL+jpBkG36O+EupdgWRDjSW3VmH5QU52sM
fQoPcdppz2trNDsvFOP9vAVPdFKacvP8473entR7pqAGCM6Oz5YvdHowOzhaF6WB
M/5k4vZICrJtGnrU+W1ydXYprjAMTXt8zRYQ0R0cA07wij6koHzsHZCA2E9MbYRL
7bnr7JJH4OcU5HhRLs4rR2hIJ+9k7oeUI28GFJY09MFGKJu4lwLxrzdkyQCWwV2d
/R1CoxAG1BXEDEm/wSLR3mIZJW6W8hQofD5Kg6UKZt5ReGCWNrYuTfDQ9J0twWW/
1rPvgoaPytG+q+14agoS3pkUQn5QYfKOnvBBNLZSrhaDg/Cv2GJlw4x1/3A26hGr
JlGYxFsvdiyxZXtCRNxdlzFkaFiXpWgow06q804e3jnWVH0qbwCh1ne9SuByVUmW
yBoP81IIOtjlEz4aAW832PpqDlPxF/vtJ/gZSCDFPDT/wTUwh9XZk27FyPBDdJB0
gdr75rYXrknAfBa/isUVMpGFdADXjmSAZXUg+LtjquBdwB1ROHMT0JUEJDzVC7wp
EZDBzt627RBxA2G+0EdyJc3nw+c7dzJUDhKczXKXdz8SDVLlbOAFrd8loJ5sgKUZ
gk16QpYj4DUZt6YOGtpqf9pyA2GaLOeMc8DAwVpBA579XoPj2WHcZZv+w2S/Wd/a
JYl4dSGy0psIsCDYJvdmNeQlHHtTaAXInQ9hzZM/pbk8tef6XkwoIXy3DILTlAs3
oaY2hd8x+X2QJSXr66ZHnEbZJNGOehkcomQ1dtmkKdbwFCPWwfyKOKoyFAGNpXM/
Bi5k9n4BAzagf749kCxh8Kb5sXwtuJCLliLLzN8aiN0CAAc8I15+/prJh+pPT0U5
ppL8iumzYlNQnov/rRdIdYh89Ux2JmvspAMucG3PEExD9Hr9x8lNypyKJqj6bQtH
vWpnVfS1C6Yzg5vLofS4b677lF3JS3PzkmjfHfyi7CqWRySFEtwDafQivYxhoDjI
m44cPD+abBcjFJCwcvpnVTavtnw+09MWPIZZTsjCGGRaEJOi8ppHsnPtYsjRTgFj
yJTy18ZkiRP2k2e30tMhfbfSfgEzps1h1eN9VzeQaYebXC4afzKI6XC1s9SCPCs2
7FZF9l79luhmUD2RYkBT8y+toTS57VLFqGJK/Cbi61enNocDwF0Ly9fnVZZN4+Pi
/6oXAetoKCDEiTd22+9sV9UuHx3xLK2vMoe5zmYZ9vZH6U3VFZ0NV7UUtF/Ml9o0
EbxuwNZmoFVnPFVZ6A4Bv3vwEYKzXvlkKZjfmOnZufVQGKvKgKthYAqnvIRDfwig
iyInHu0qJKjeP/mejGENQ6m68iKINPe7GXFKxgkOXkKgTL8Yq10Q4Vr6VUEGRzxU
i3PoVEkhtTUMW3C6qB/WwoNavZLxkxPq3qRz1ba0zPERWoW2mYG0K/puYhf2L3LV
lXG9DPRtgOctuhzVwHrL7tB6b9QtUjpKch8BrUVskXXjwVBPTRf7gDcF/hLUnXLH
xaaqG2htHMTn9VhMhA5fOQAan6PDtWSY3sswRGHZnlWQ5jGqenyutG5AdVPjozK/
8rWX1PSbqqg0/trUVPgOgpfwhHMVUKl+ii7RtgZfuB12L0fIPt1Mjz5fXrWEM4cM
+rGeXi5PYfuJETcCwCUt1D2gs0kfsTZ7zqOdyZQ2f0hiW7EKCl13avNUExuuRmWs
Q59IukmxpomA+QHOEdpoqXYXmoglf+LeM/856q+kh8dnoNUrQjyB4N0x+wvDhwan
AvB75/sglDYnl0cRbxq0eYZ4US0PAX5xwBsM0cRE8GP7UKEDpHwW4MXi7tu/Agsg
XnatR4nx9CtP7SbKX3StcXVGNb4TUozqCzeNVsan+IcLjXvrNJdVQYMW5VhvOcyu
neVVo0CFIueACSnaOSlqYUJgcVgpey4jWEMqSZC2tYAoEetUem6HvE7zgqJzKebD
CbBPMeUnvSGex5Bek8Jq81Fa+heuZSfJ4bNLxX/B2tsscygJL6l84ZmFrHxZKUPR
jpRW5rDZKEpQxwpkTYVj54T7WxLxs6R4y0bIqeKvqUtIbnMK3aI4J1ojdGCjmRRZ
CzHKk4/zn2iFbWrK+LEN3S5CDQh4MvxeC7zA7mVByGOBXs2zSUlITdylLEO10cVe
nlBnNMPnM9SGcg96Vw9bJtoSw6FJ8uUfzca3Q39ETdEDyZM59jxCG0Ct8T6CHAGZ
yT4o5rZMfC3oA4KWG86D2Y9fYAP0RdQn2k6gJMk0x1i8LHEnyzrJLGsYuZLvAC8y
t+TFfWRBvXjJP1jX8Hn9R6V1w4Sgw6Wm2eq4iAd32oDvL4nwE/Qke5SajBtYXqEo
OdRIwzOMIgZiwit5dlYU9DddazDlwXPAz0ryIt5R7utXvuAutG7yLD8Ybn1FfiVe
4svNxpKU40vauLpa3I4sMYU+vYzet2+d8oYVq8z75CHF96UhXjNrOok2s7hFd4my
Gpyuauz2DvZo6c6HJbe3ni8s24z6xahm6+RNU8pzpxlYlsMWGRo4a+hpfvNY68UV
09TR+WqwxV8jB9RtvQPhlFwiFeU8MzkmaFMoInPKUnGlgFhZaw9OANweWLt7N9NA
NnFm7r5pKaF6Z+5QTjFq3tlAfKOvqXQ+uZJeN55qreaMDDNf2SLgz/y3uuYKU4Lz
AK/gW81AMak+LaDRYp+pbBpy2a3AtUo5NBP1eNKZeXGZCA/Rq31GmWDNNoitlTuH
Z0P0L/g299Z66xk+lF6cHUPN/Dr8nzHNf1ukbbX3FXbrDuv/LH+v9ys8UH/ETk2A
C0JBWW5idxA8Yp6md2FnXgwklZPso2y+Esf5JJ8Q3FUu0BpWmbjP2tPpW+aW6STM
7AleZ2dCpfBOtvME9AxrQSNKKGPNrmFfhCy9KR2rqZlIXpnXFF6kdXs2leRM9hkL
IPEjaM4mHHpjNDcKTexA7dJqGN+SSBVwdmrdjmAVOuQp489ifb+ByZpdNeLI6ZSJ
2mQp60Zu/pUZFVSmc3ROXORMDOc6K6MoQS07hBSEYhE7XRPuUEiqZ6wgLicS2KID
SW96GjvJ6VUxr2pTFBY8G5WFrsVRwyWy8k65JZuYVoIkbyCBJudJTsxhtn/jnJbA
6tKppogxPW+ibu4s1uzx5tWxZaltRkqh9vcsF2lI18HRKaA3cOT/KAl7tAXCUgsz
BO4mroH0I6+KLVSP25XnhlsB860cNmyl53hxXY7QZ9uN7KvJbfIu/L3Y5D9wNiYN
IDsIYbaosBw6tYT64fHHFRS68XXQmfCAF2Os8y67ywzbCZ1Lp75VhpthhrMaZWKH
ZqzKvxD/IWyY/a7td25dahTZ2jNPUK+cgt6F5mB7sc0PUsyzqo7LSSU4pqDb1aOr
4RvOwEpo6nvFDyvP+Ml6zIoAkuWncdZt+RzgF+J/w/7ulYshe4o7qdMFQx+IKGAn
ogunyN/ivWNbGlQeG/b3D3nxU1dT5+8ehTgKdnmJJ137C5uouOdMuY8Ll2BkefJh
MMCioP0r7CNW6tm7z9UUu0qFeJG9MDzIokub3ouzcDmw9ngPCspX1OVdO0dfi9T0
irfoOPSE1YnJ1r+WVXvrTbR6iJKjR5hOvQRlE6EzTi6WdzPECzng++iWFae670j2
jWV4pdmcBpQJctwyfN7NXIMKDPHPvMhZLzrXoM/iWTb8MPyWUivn1W1tL0T2IaZO
i6qxDco7v1XZ+Bstc0lAQLs6Bg/nGQFMIosxfnIuk2A4c4f0m9R1u2MtbwwGs3Bg
05utpcj6R5fb9IZanJSFIDbdvnoxS7kcgsfb4oAry1yoKJ3OKg3g+IuUePAARgjC
tO+evC+srQvWt2mU4y2pyQ+Ia0RXQlfet0ryVQbjk89giYTXU2o60IKbbAW3HVRx
XBToMR8HoEyWu0HYabzgygqS8xaPmFPlUQjU9rnjeCltsPLidAYUJtaURVQu4cs/
tgZ81UWlYi5K1NUIqVI75tqjTTzwamkkYSfgjUQWqGJY5xN/6FXkipI7fgc97Ri5
fW2JFjPHcLogD050kU1iBuBLTCzzzOIYODeTJ8/K/9n3rAFnapVUOsGA3jn0vnKI
m5+GlpamFcKVJAgNxY0NbjPe1Q6Y2fXTFYNLg4WvYRoMpMj63AdNcdPs0iV6Irtx
oC5SrvtNdu8AEPTbDg9Zr8dv/nlVFUNcaMmPu/7oVXj8mNt9xXUDWCDpyM2IPmEY
M1R5E0n7tkNlM9rqYnUSiaZytMjfYB85bXP4Fs7kwliR5x5Wo8vpTNovoEnuPOJ7
oTRk9pcEmG+rR0Ye1y4WtFEfqzRZkMaTn40katOrtx6P7Is5tBGljnZTTEnDLwGQ
jC4nYTt0tFAtmI62253rZGJBaIMo+bkDY1o6hiubokcvlEDxWmCyLNJD2/8gli02
CeweEZ9bqoy6eR+NbMC0STcMVDJUdpJlsmrAeEg7qUW40PMV+3lT/2rZHJljo0pv
Ej5Qc1ZkM+WlvNhFfGOn4XhrqlcASyi0lMnRuhjpL3v+A7NVIeUnsQxEyZwkeqki
MK3WBME9jeYgjTX8gcFjJ98lk02pS9urZM3FtONV893/7Ogrv3AyGtY6lFWaHobq
9ESX4ogPWqRH/E+VR3wScrAkbcXDVc9ehcS9tBJnZbA2niqFuBHJbHNv9szzGbaO
0p/gYqhkoCtShlTgfxz3yLNT1utwguzWEMlISpu6vt9jRVpgJ/iW0+L9UTJ6Xj1U
oJgFrYFzpAr9xbrBL2fS/1GQAn5+NI//nZ6xaMxarHJwsDng/IqDVXOrLrgkxZ5L
zBugEaeJOcDxXw35tg5yAORlsEt/0COXigdZV+sM812hkXA+CfL8ByR7MSFgqiRD
uyzKyWfwNs+WhVFF48cdXj+WKUWjyaU+eodrFP0Qv57r30CqEM0kNhxAO3WXWBhg
ApoXw/tD7GVsw8b67mrBMJ0RRTTnYZdRGd95oicb7N7qgeYROM5qwGXBKAzDSZxr
tAbNn9eVjPetuXChuUbNj0Y67KbgKUU3N1FYvcFYI/MWhrDpswgoBq/3Rv7mTX9M
fIwieSW0LAC/0IsPj21kuG9LxV3oAgtfV06nVDIyKehstTp0IID2Z4KSq2RatIyD
kJtfbUKi4E6t5scJLPBIex5Oj8epwvVERzPvZbYwv7tr1MszBL0V1vk+bJmuDElw
mlZpOdu6LdHRKV1EAzFDNjE/Ontcds0g+6+14ezwiJjlu4o44lxCiPeVMrYrWYBi
rtMIKCLAAodxbZqg7ODRtLMzI9z4pYyR53JHnVtz3VmCCLkxLleybOsiw77jajTa
eXvBv2eCYD2doETsKuPYHgQQSmRrBLO7Z2/PyXslQSDk8s2o3Y4NwZjrw5QuH8La
ozh+V4l1hJCKtlLMEWW4mcR5S9OB3VpUEXko4z6JHLA4Eyf4v0dkX/nVVg7621Xv
bUimJRwtQG83n36+BwNtMOPOr3FtBmm5RKNw0JsMqYuGUIkePenYY+m1+VousGBD
cWkOfUHaFfAbnajTjkQ/NZ5qSap9vlSvc/ErU06JO7/3zqWY58HvbIPQwTRISn5g
TwfPfWSYBxOHNVMAyMKbyz7aZOrIYXtr9nvvInuCXisgHW37rqB5nucnX0N+GopA
UzAN+bSjJyssFwPIADhNESFimCoINqkG0QNBpmTYay02ZvLbOmUyTbi/Ur7gOV8V
PvCVOpZAa+uER5QZODAoTOUajMMm28S2HBux/GkhWvyn9rLE/BHDGdci2hAJHsIf
x1rrKemkudF6ZVPo/Itsw115QaPi/1LFVHwj9Dh2d/PdJPJC+tvcA0PuOxBgwIx5
ZmYlRxDZ9JldZcJF/D8CF/yvFQBdnt+Jygy82hQAPpDffcjfc7alpFxgCaKoOIb1
4f3lh5zbNfNo/4Yn4xUVdgbHENPL9Fa5uXqyX1Awpbs6glXGREBUQjlUpngIVZB9
tlY09BxwyHjHxWZgcFAym6/NbeHWOdHZ+DwMJs1RR+wYeh0GToVeYCMS6YtZu123
AyOPD9J2+it11WxwcyI3cuL/2qfa7rf8WTgT4CjSnC/LjvRZ6bCY4HwQDEcUM/Ph
FkUadCWnIWu/c3tYptmxSDZkN9g2o1JbMPNbDazfZVn2GSxYR8l3PfX7NTyS07QK
wEHNGUfK52udQELi36LH8trVRZ+/yPcQ4shL0fkvqmCWnBTD5te0yzKl1pdgCx8Y
eq2ibTZOz+NmJJkfCjuvdEzsteNy1ONe2vhGdZBm1G2hK8YHUBF8OrXUDFpQQ91u
ui1iyUIExKRelowwCy9pa7wFfsIamhX9Gcrzwgl6OQNbZ6zXLj+nKXPuNObhTSsB
Avkne+Ug4UUI/t28yUOdg0jcdcFypee8v4AsXGtpdxp5jrsZpj+1hHljk+4MqgRu
vFdw3nMw7CR+QCjjIpDrNIQrr66JCdVxwD6qfcngrYxi0nL7SX+8IUd847ln07jE
CMTHwFfy4NU2/g8WGZvNfD0BuGdPEunDrX/kUhhHtag+gMTkvUbeAol6DUB0V0zZ
kqJhxeOANRITw5Kp1rRyB7W8xnPC/delqSCgGw95oGJgXAJM7kcr4BmiIARl3Cvr
s+ivfjPninfPqkMWWsa2JQq65SdH1AVQHU98pNP/408DKpXtbqcL2tnYAfOIZVWr
h5Y1I45rBhVGHfynJDRg4oPyljQH3Pb+X5Kv5MFcoNW0dHsVr9oN45Jo/e8lgpx3
mnrMI2kveea+Uzbo2XWknCsHwL7tbcbtFs6viHhQcKODM8J1ZpDdV4sBu6XBZu0k
vq2Rk30kp4oeEzmCq3xtRggcfxJlBIRm4qQVO6X5R95f2BU6WsMiWBnTehthDD8P
+Gx2jaM4N+8L1SQUvztDfhrMoUXySdOc/4z4Ds+yuMdznHX7OBl+Yvyo7aofb85J
uuEpAVOKi6JEb77sbWL8l+4Rkt/WfJrO/WwfhTmbBG5iW+tc6QOhKhzgAabn2SYs
3A8mQpSxz5PgFdonuny1sMXn3OazdJqXfYGAu14XYaRvJlVvaEBF79m2pDCjQmvn
ChR2DS91YJbJvmGAjfLAUiwTn7LV3wF6tgFvVudkCI3IUyJ/gxSD7YF1zEWwd2lU
kzz955nYyjvx4sYCoIpsLvpjS2FW+T46RECse2xWgeRqLnBjaf1dK58mNZ73SjRG
Py+RFi9DiLZoCWu4Lbb9ImcH19JfsLPyvNAwkUmDEjog+V3JvZ35KUgh9KRGqcOC
qXnWWpyKnuPUc/OA9CX72Kgqu1LDKaYB/TQi71RRDo8xSqVfza4WvcFRFua0YRKo
suGIlgHeq+FP9YklxGVl1IQbwT3FBb3idLp0/ZTjw2S/hQlaOT8tQb4YiPylFmsp
CY1ql5/y0vbtEfZKAXevstP80WmtME13tOGsUfjz7qYLpfnQfF9QlIBRB3EgQEop
oNdZWphQsElgV+MHL5j98A==
`pragma protect end_protected

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
o95PcSJOj+83Wkoc7TZOP0JgV/OqbSisf4IOCZo6D7ezBTrpeky3eObhbryR7HNF
Q9zZAeYNb+GlVxjhdpOOVDzOs0dTt6b8iiojIgPyTALR/XUd1pKLYCuP+gyzWLhh
t4ZMDG8ZkO/tKhADTQPMXuIez+U/MNbR7ExLgL48sIs=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 3056), data_block
eq2BWcS1S6sbjPRnLBQBWtTQl12BljBYQH6EhW0Yt+nk7gXQ7PLU2LMDmOSaVRFt
63P0BqvQd+WtAsnLhHwGFfIohCidNW6hgOkgeS1dA6JObknKiHtH/mI7XlSk+ADc
pxsdzaW8OJmIJJobFtaa2Zu9yVzLdodNdSWJmLTWdAnTkxfPabFjGuZRZUXGQVlF
MgHYjk84rGfUEgZ3HKdQpd1xfAW7ZKD3ZWXjWQ6eV/Z/ICqMSXPZtKcBdBdk9fBA
JiJRNXpnADv7HsTx0U9Wy6sSmp1j7AWCSECFGGGTm+9bUiH1jXuEufgmJieum/Dv
qWH6XLZqw4W1zQ9EWzQ5ZCGcBXpCnFOc9VEVbUibfNztSxf8trnNjM98uI/obt6f
BvggjX4e3Meo+VZ3arkTtwYjl75uTuSvyxNXxEb0bZ6N2ti2yrMtNt3+MR2Wv9JE
Q2/OTKLRqY0411YR08r3p6g5oYgz/ZLYBObzKZHOrJqEI+Db0+PCGn91WUpRnnEx
Q/Q4aVpEldGjilDsaPZKyc81C7f/nyl9r2zziGeOPBoZLtMShGdZoo2zWrYkUGro
GrqV7F0xBZk8vhLiktVI5OFdnUJfx1RVX6e7n314MbqEunRzBw69EkXDBDIyDt/g
wSj0OQRj1HLhOJrrr+Mm60WAizIJz8Is5YvBl3eqAxd4SrVzwMRNmwRVPDbIs+P3
WiBlOGoPy9VDHtjp0IHo5++gvZixDovtiKn3Vo6M/xrFwE2BuzbD+11iNN/povbA
hFoWZWifzyN+oB/xkbJkoGSXXg1my8OO3i4H/bxCBnAvHtKgQ4omOSm9P4r0ilHy
D0UgEAsquitztb8Gvc+iMUBFCbTT0zufopJZ4EYO5FrnHRJT+zudj2iG1ZDh+KI8
0NNiBoyHGn+ZzmYBY+QLiwl7OuUCwwCBDWSLxdrm8WAQLhza9DrrBqNu4MN/EB4j
W1MUNfCgJgh8QSJkhpe86GM83NJuSrrDX5vgvtqFff/EwaStr0guW3Cq69SedZMx
MqWhil9nh8tUxih8EITdYCT/PB31vYHOlxy8a+YHFGF0iDNrJ7BpT4TbNNMxeQh6
AZnSi3E0tvy998PN8gJ8ZAqyJPI+7v1bck+loTQEORgHhVjmK61ifzgaVs6CLWrv
myWh794yn5fXjAJEdqIHXBII1Qgrw0MdI6BevfFgNxEKCxOajt+Z1t/EgYNCsQSX
vbYxYBg0cInHj5tvq29MIqwcaJaeCDahu9vY3oZqKMNT4zXOCaQke2YeCnlRQQqw
niYsQIbSDix2kkp3Fwjuq6SCXqJ7VsbLwKTdE6n0jAAV2qoMjPxFMUC4hMnI2XS8
7OzezqIz9sBprsKuPOx/+xz9N1oxZzBfapVOBsCmN4yD56eN5CyRdZ28UCnnhwjt
xBzstkM9wRHSC2txnjbRmAvl7JSR/AGJF74bIZ5SyCyQ75RHEUO33U4Mo0WCy7T1
rlFD+3lCo8e/PmSuKy2cfYIA5bRJvb0+86BjSyb8NKtpRYAdj1uvhrnJby50nP3+
6D6t2TXzaVH+FeeN391ajW8+J+o7G4hWPDSSoU+UtFchTpFoSs6eYEoxYEIuxf3U
ZwEEuLUw7T1FKgl8fwtrYp4pKyEcH59d3pMqVFe1xzpkH8A1xC5a6LHVCi32MaK3
aB4wu6eocmFIhIzYwRqEBDtPekYFJzFa7lrS0LETbHQg+z4tzVWYbBxt61MTQGaW
stMWVDp8jagEbjuSnFz8Y0AuZpoE2aKf3UC/7o96fco6FTYBzbKq1Ep15rEc7c3v
3AszEwdraiKIgFGjaO2k0qtBK/fxtjSwCS3vlsVOwEEkoKM+QWma+ke0/u5Ogs4x
ebEK8G6nzGv6GiamHIGM/cGJ2pL8p0Srmd4lDTHD0Zle8jFeyqBwFKMrf+qc/a98
q7PZgEqmPMGmmyUC+CvVZdNFXuarHib8r3eZU54dLcQ4Qx03G/t0oKGu+aTw+8nA
wg2No+WbGWPWlNB2+/jfeDmn5j+I4HoItG2qsk9Y6Xw+Zpi8+uYEW49E5OyUSyc5
8Mhbo40UwN3c5vLs/MihCbl7lg+NqgNnocc2JES/0Mx/CX688pRtxVDSDUB67jf/
JOop52MpfRsIyrsiY1V0SX+7+yPfbjDHc1dKtAXSoqm35OvPC+bDWNTgj3KTcnFF
APR6xKdv5Jk2KZOUiLLReR+UTKJxI1Wo5ozU+8sx0zatn7qKaQrHPm8LCGdqiwTq
FqmB1gOAy02so1vVneE/tJkB1eKoGtHZ7k4kSFshAYxwdxk2hbDKsDQmdbZ302jE
KEUcI1/R+avCovDrdZ5rNDr0WCAn8EPBaLzkGkc+LlkxuASEYq29604Ykw4BBYqn
wjBSNrE1gTlIFR0rCowxqszBEdA3ePPrmMEJMk61/qj1rNtIwTX1+Fds3BABHU8U
mpJ5VAkJXS5/X0J+h44JafVifvyPnpoEiShDt25aNCz4F2yDZLH3CTIKILzsWfD6
QqxR/CKG/xltqgP6NcL/E803NXzpzBwmThxs7P4Pzns1DAeAq+rnajuKyWkm21Jq
wOlBcdIg7crKjqDuuAIMhXEftjlXR+kWW9v0A2/z2f04+k5ajWoYuYzmFgC7IvLQ
tSCAtld/XQOI0nirx6GzeC3BDvVwjfk4gqi2aZohhXZ9IS6s9wDtLG0ugx9pqyxh
LzCcOZ+CdlgH5LYhjHgVcozteSt6TCO8kweoM/0+vpKbKWnlgjN2V0rqr5aVYdhU
VpnqvBWLMPpboMkXXVF78klKIygCNV3Q6/K77pIWTaXDTak1xDxgmM5Vg5hESP9D
AJv5qq5wYMel6vybh8aPUOEWLnrtErvuQb/JiOicPUczSas2K0H3cOW4VKfuF4ks
Avd2+Y6Qiw8n7a0IiToQLQleiGLzIzZUT1KKvI+ovSo34wiWHZlSzDwXv1UVkrkj
DbxKieFg1i6VJDjM5ds+jU/BevEH0MotgXNZII9gbkC0YVJpvYlilKn7fWve+aFa
ufPMndLjSmFpPfD3LAJpW5KP7ktueoLYHZoQx1tqf5rxI66iiar9QDoWvB4OIej+
HsR5QWmXfQAgEGr5zJq9dQajjjMNEsvv1uBLhEtJ3KUwbAaNANWg49MDStMpnNqk
g7JrQsDqSyo4loxcsI0nq03E+QR7dnp7BJFvs5iLw1GhGs6X/RptAs4aDELKvm26
Cib8G/XKX5q1HqFjsHynbvwqlLpEyJwBSoDxJuuAJ9lsDCL94P7WDJ5+UTdJoxXO
jr1oJQ2ElwQZ0Ihd9wV5fdJdUzHNgZyxJ2OSZ7JJrM75bxzMg1BFnXZmFXelAGET
p5eaoLPETdR/qZQjTIAWE0xsIQhqq/RkQk29iQJfU8Nyz9nH+xrhCNg1uxF/p+s9
Myj162HvdVDQebHVRAwIFj2TPOkiv3i/zdjjEWOTZM5c+G3XKlinagIZ+MT8w02Y
aqt5b3KxeMQL+7a0jU51C5pNc0v5J90qlDPxzseIStHATMnYYRMGazqUklDhmoku
9m/9hPbvV/j+y9vnwTJtvOT3YyCXf/JkQ+QtSuvBypPxjDV1YMgnVlS1ZnasuMY4
TjvrMgW51IvIMy8Z2pKCm5V8BUmowjAs9/yex9mU/WUL7EigQD0NY082ImrJ446X
yEt4bHJdkQcoL86WCUm3PVvztMlqogjgfO1LIWU3JIQ5iPNDmH9cLnBF7caQvvcz
O/vT7Z4DpcNn8CvaAcfpmNsHu9QP1/nW8yMntZ5dWfsrFVVcOYldm13gxoSPa0pp
DKx71itUEyLwS3GQVk4CGYP+JS3jCLwW3Lha+r9S+PnnxjLgo8zEOh+2msPSvGNv
E1AwPPsWZhIFcftZ5QdimI0eYWFF7kxSiPjCsmzncpLOXCyaj/UzrmZjyXQllZKR
jIs5rFnUasi0TmBM5XW4w2IgpQf9mRKFkphPZzv1/1rWI2dDcEvcTcFoPaT4GqDK
D5IyluKuNV3Lip6l/bekJIxJn36h44X26qY6af0V2LwS82vV4E0wAnxcjaQKseJV
9uEpRmOXGhsQ4WSOPdtKM2X5HooJf0UpS6Vf7MLC8EM=
`pragma protect end_protected

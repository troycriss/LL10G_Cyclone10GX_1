// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
Ad3sUrymvDgQjeuc7z3Dsy81nBQhbqmq7hMCs1O5CiyrF1XH6j97VMdQtdyXoAsigHcDtJAJxqP7
sHjoUYVmiYRK0rSHiX0Ny6P2i9nmjfJjR1G5yftITjfDFkl4P5IP6napDvmNgEmcpr29+dZkweXL
PUAJgqcayc51AzZ+ONZ3WyJ/PiGxEu7uBYDA55FrpMUR22xDJA6t+h4cwoDM7unpezMdhgffGGuL
/WiurAE5DvkNDJjwgw171Qd6CcmtP86wqA/nFWMBeWlmzLxIwd4klawaBat/E8kNaaLvyWN7OUx+
MmsNB0FW8MviVApaqI+ggrrBqSBQzpQ+5Zuziw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 59584)
WosViTtVQZy7eBIiF0FQioc1Qn2bRt7p6Ul9/XI+M2Gytd+hR322cLrpJYMelxFKzUn56f3ZQWS7
IFlQbnOZZfa75wK7AGn9SlPfpIiRuFM3r4/9nDgRKNtT4S9If3BZJZTItuFli5jURXJngRE9k1K6
qkzHkP2l4s/QNOJQgjxEZKppXpkEslFuZcuBb4m9vGMGITxLA+Kk37vXK/XVNG0pOqg9IgN/OKBp
lY72yu/YVd9vA4pRDUI/8OqUeD3XM35Sh/U46UBtqVFEaarx1qwKE26elPHBbiUJNVeeA/MRgKcb
thMoyUtWBWsTG8yPQj0x5NHyunHxBUrLAlN2af4r40tdH7sccsGFhUjiRdOwRDaJe9IpuYKTGqaE
4kaAjUAytcam7oxD6+AhtZyNLJE9saY/qb+HRQa5cvo2gxVrIqkaNEqsh+wp3dQLGSXrLuclsrIR
1u5/JNUajbUXmyjsGLrKUubJf9b7V1gvJS6fuMTbXzYUKSuk1k/5CPV+lsNzQdqLfZiFnjkYkcqy
qWb7L/OT/aFjqN+8Z4q9RFhlJoIFcOfk/Syl16sN/dDTtns2bmZw0mWN8vbB+CFu+l21+mcWjSnc
JgDZwD+z4h0HHbRm/28bQ7ZjfMm/xXV9t66aCzIjC0eXByeGBa1mQjYNOBrpq3LYEVXnsz+kPWdT
dkZC0vOVAdTv3Cpyayb19egfk8htUyBS56ZCCBxh0rns9TI4m+jcFbWIemUMuskIIzySLFTvmo5K
+QU0MVhygISf+1oRXd6uUqpqOahkYRhaBF8j8zGGwauG7CeJNGRLeRHeAqQ1FScXWPWDKPNGa9gq
BZZcakaUv5eQWbzdz/UfW7ndFv7RzYiUGwGZDkeL4Eg/5aVnBiDRxxCnbvQWORom9r3c5F4RDe7c
aEkm9A/Z9orxPp1Ml75QcatQa5dYvpZYJeFgzKNou+4GkFhx8aan35t6zoTCuBGGZNtRi0v6NEb1
kUYu6E/CmkkKI0ZBu+PkaK5dSz8AY8n1z4TfsKcSjaXqIbOojLkViqBqggfFAdt6jEIyTJo1dlxL
5Iv/IGKksNkr08IdCps0/d/hJ/2cL/5fMGMmOuJjBBIsxgnOWKdw/BdFdwwfrXoCI/65y0XJdKmf
BJx/cANi19EJ3khhry5dm8hAW5q2KKA0avG/yh2z6mgseY2Dx4kPTS+fkMiQJeTghPN1lJOZrG96
P6UJtC+OrGmbzIWERhoGW/JLW9f9wuaysJxZAXPc84fzvLu3QIvi7pTIH2d130com+ja6kGfx66f
ZSX9hBacmfW/I98TfUSlIxaizvIZwtXJG2l9ms0M8kkiMPOWUGby57xIvGyDd+83uuZep1L8vVHC
jOa+qOc49B7ItxLAHM1UDC80lJkVZwoPegkaEaALBOdWJSXKFNbTcY8SYhecNqsSd8cppZcxPju/
lt3//S9rH9pRKCy8rICz30+HP3asLctEPFcz2GPnzKc7aIzyuzQIXIc4XhLy8KvJLVd5Cruzp63t
2cnoKWLUxVRMYHfvD4e65lwp4KEO6eIfKo/7OOtepbJAnSwBZxfMSyDP11Uq3ew61TFbfunsBomy
mbhaj1vwepKiQGxCf7bXMPx83sYyr9E6PM52SsJuXMEumb28NO1goKXhJQuog82MQzIrl/6H1JBu
JG8nlUswcJRuoPN0MbHJWPj5aT8AsQs7erbgd9L5HbTyMXxrm5gSN3RZ/ahgJmN27uXWmdEcVFG4
wLYy/gIdNXw5qGm9uM4H22OpEQYqOh071ghKZfnDGQT4DwlT9ZBqW5ps5oToW9qJa/1hOVoq9Szf
txwpYIQ31NcRDjFQsBeFFls6UydppJX0kCMH8KYBoBhrCUBLMyAIxJ1eqHepxlo8OXwkv1NPFx1H
wy74yhEpR1kLRry1+wkgBPvE0lGKp/g7fuRY3VREWkf6+FNA2bB9i4GBlz0cL1OyQszs9b51BJlg
SkuemJf2q5T1oFrMOF4syX5MoBZNGWtOSz3GuDchnBENGHSbmH0TH/KR2PSJRi5+C/XvR9Gua+Az
XHfm6qzOEhDawIdKp32N2HL/BAedBYO870CuJCxpSv04FQWTGpcPxpwpCKIZJXJblUqMGtWb/QD2
kpVc/kk+fYQn+jLnCLWkSwssaMQgvEBLNl+2IEt0fuN2bLnNKyUbtihJcXNrth0+j/15c8fuP0at
R3QYSOF06QzjL4mtjWRkD0oybScZFMdtB7BQWrrcmoXVagsERAATNxoFkU4g1SWaQ8HqSemLZ9x5
htNVqQlM/BC4EVet1+i7tGyy76vNMGV8/f+a9hCBzUbhZoVI07Iwt0eq86JqqxUBv2ZdnZwJ31XC
IqINGwTL4Qe58okT+Zd+evRaa+cx168CsJvfOIEmAXa9x9lHylp97RVmuOIaLdWCe2QcJxXb05MZ
1BXxAV6Cyu/HKc7nwb7NHl4+glVRp2ZAn+6u9KUJaAZnOsGogQ/OhrYZmiY0t4TZTzv9QtSD54KK
eZjnIArONd6qzKBjDqdaHyQYv49VQm2qgPrE6vwqmVpVFrunG5KUwbr4vav/UwmxoXA4Y2EdHFB5
r4dv9CvffPpY2NHpfNVnbCiQAF46JhufdGAuxqhjYf3gHL4bL/MDBt58wiedzdIYc/O9RmqPRw6W
eLUar0Y04a0Eu5aw1U2lKx55rcjpVJ/QXddOTu16q8B7kD+xG2w4UPPxilbuim7ImLeN3CgZK/6U
r5P6m1tdAMup+PukOXXAardZ58M/G9ZZUu8yGC4RuWhKNr9JWZtDVq2XRu4s3qbs2EKRJlFld3Dk
p6ogm8bMod5y3otMdSu3P97j0orMJg3wWVyCsGGCbGU7w1arrrZWD8jS/pDKOOZq8ZLeuunrhA/O
wbKryF7y+9nBO6o3DfZVCc5U8XiXgBezSjP9hFbsZABV9Lx7fSbQFU7Yn+eUFfSp34sXsKDI8T7U
Vw9nEKPv9oQWKWiHNtNluMV7lFDFrHl1J251pGkio/pLjssKA7nC2GsNsjhd8TmbGugahtQnO6We
+eQpxQwoD4rA3XVnQ0xQWgtp5uUXMfIV2N1vg+YgdBlQkcWdevF0tSkGU6juzP5VSkrI4p6Va2rS
C46B4iVTjMjNsdQaU/0Y/XNSgcG0FOkwDwQev1lmGEvmvchJ2hYeNP0ttkluOc7R3lCN+uy9nZw6
fnl551JYSDK2Hstc+HNYC7Fkk5dTabpxczcv5GulIyGITMIyAap3D+IqDnzmpegKLEUdefHYhgnl
GzoYPFmO8SYQLPwCK7Tb0yE24gYiQKuBwrYM9axBJP4nIu06t569eGQgAG6fbxU8ic0NKfdHuq2Q
wg2tOQFvcc+XTHLOo788traZPncd6Mmb5FpmjEOrkJqvlQh7ItFqjdPZk8E+UpW23VDyLQcwiEWc
G5HfdN0YHGs66adkpmtBkOEr5ez1GbKypXqr5A3bJkOlsQWHK7DEvQZ3z/ZTFuiHG6rdAZrE+829
3KZwIkHfUSdjuBvEUtRJ9OF+xN5zm0BvC2UveWkX8PHOrwSHZ15dUbl3I45IqhIYp/Tf7zWoJ5+v
yeBIIwaNWvbI40YjFDiOc9dS7eiq0vek/aYJpU6IHVrsTbfaT1LMbqZ4suJT4GKA/idCJtkqtDyc
GCKesZd4yzC6/tdXTYvRj6OShjH5H1FToBZDviwq60wx10H5qJ+xs5f8GIOfGSKc6FXSe7/woRiw
KlC6jeF/IC/2oJogpemcOFqYl3MmON7+CdrMDmJNb0qLdyXhlaayo7PhIAWVTOqce1dNN5BNhqCz
XlOufEZEeDfojqIzrymikjsj0Qjr/Swl8gMKaTaFAo31ipkG/c3BOMbsF5UL7gXIqvt0vezWJgcb
q1OFBIWtcD4WMgoj+cdYDcgDb5RuzZGRQ52Rp6EDA5tQbHXj3918xhEWrT9668C3v6EcvdSMjTbQ
eDHfTz29GfcJTtetrZrt/VdJpiHo7fMMwXADVh60W+ySL1x/aBCCGBigJD1zq7gMgTlM8QPdeTQe
yypO22IGLz57TiYtcGOdi/r6kQHGL8BV1HuZTLZJ4kEv0S8BH5VbeyUwZApptvsxTJFd9QZJ8fmP
E/DauSejv9uERMEn2i9VxPLho6Qg+PgjA9+B9GMOzpl0aR6GtYwDMQd4U+KZileMS2Qx+ZC2dq57
F0qYY12AVXZgioJLgvZm+KyRSsdVGSUB4G6p6q8VZvr3aTgLtlcNcCnF7hgN6FCifnRPGyABr+kU
szXHCKMiZVVdI20avrNF8xMTwykY8PtEMb0SInG4aaqiAEvY6c7sbomy7strRK+rSVVlbKyJM4Cm
g1wCJOtj68NPgUQwlIk5F9GRyvwpo0hMxkQeVHA9kt0FBwBEFvPb+XnUh3Y4KBaTMZWLxYeHNAbg
/lcu398wvHShjAHbMOwM5nLQXPi8qhsGK5+lf23rQEGdlmjgdfvlcapEZc57hhIQ1Zf+PgEkYkxC
p+v2UAiIoOe1FlrGdrBSa/UivvlbQTbrwZ4zQ+zzRr1geyLlHI1C2U2Ld5uNO5jpdLteR0S5ahoX
P5M4pcYozKftS1HoZ0RPs2eEAw1xu3+p9Z2LYB81p6dp7TMBs8Q0d/6x0Db1VAjtUIK1ShxBjQHM
UiPhvnF5TKqS0ulJQE0s2Xm5KdxXy3qFW/3X3lmLlYX5wekzVVB0siQEB/i9L2C8pSkQL71b73jq
s5kKgM1PTa86nk33dLMuik+Tz6L3t0hXUjGqwKokR1TieiIYbHBhVw5jL/u9PC0Z1roGhC3YDfPX
tWftlpYKqWKiYet7V/otoZ4YF4Vllq2on7jPGsN2CmuH0N4yZY8qq04Mb3BkbAjMkH+/381E3sxA
4i8ziODTzERwgEZXcj8r0KnhZ5mngwWZaqs2oiYfl9b4ABTd9irW1/sZmjPl/EGqLI5qqlm29bTf
5ytXAhJWyqay0p4bBycm8hilFqBIOEAtA+9ZjIk0EKbnknGGuvv7NTWwTKQeOgaJeVJjTeWtq78B
lUvn4HA5MRoYjDk1O37iq3VLrvICClT/ZgprROQcS6VyFf62nEjPK3W5mmPYnD4zG0sZYr66K0xI
qlHXjnF8kYFdmPQn/+S0fdk/2iGJLvXfeXytEcTJa3zpJBYYx1+HLnaKDqR4rLvMZNCSygen1QGL
vSQw6UbHaU9aZwLogrWCHBcp8S7XfteD1y0CR0ZPMjhTqHWGkUqNX5gQUYr8HZRCDhY7xxCCs1KB
O+oZnTWo1qQ+DWPhkJ+ZVVOVQuKk1aBSAqgNTSRU0FenmuRrTjcl4PMIA8i9BnwlQowfXFekf7ae
cQmkWhW+AmS/L9DEX6IjsE/1/zVME0Y4q7K7oqkpX308vi/fmJNqJbcpl+RJTnVv2/I3k9IQzwzn
EJZkZugePDsjxVcTogIWBsJJN/N+9bcvUrG71wakmORdz5RK9uU9BhV63hN6SrKnyvp79axJ9eAd
4lvpPMtKLY0MF6LUFohSJ78hridi6ktjHjCsCdW1XpHp2UnLGSuu/u5ICevNzoR759RX7dQ1NaXR
8v0USLhBQ2KHFA0q6dxIT9DrWzHgG9BKimweVlZtT9oGZ/pTATtaCq+7KCmOw+ZhplRYF1KY2vB3
yh+gfVX0FdE4eVmT/pSY9pOKrHjMQsA4+QyaEGdr8HhzL4pvYFN/XaQw3JL/nELPrJCbeIc1rrv+
BKTmoGnN7654crVwmjXcCaZNSDV5OvGoRcDluDhm37/3aYBsyofA0xPZc/O+BsNmXSowfZUo08La
flcrY1DW4WEo7ptyOeszFT89WcUXwjsFBW4VNT9zJgq4qDRYcNdcTrINm6o9CRX+Gak9NJO4m6LM
Zu3m5DSLQqv1FU8juC59cfH80boWkc6C3OvKsVsE+SU++MTNCUyem22OfXyqkrO/xD27CE6xXZ4f
f5728si0FtaI7E/5QqXBETXsmx+lkylHcyZ6ziGgHDL10RjYZdWj8M2uA4NhLbSN4WCKr0AA8OJr
0S7MK3LgOeBx6Nh/SuQ1BuY3dzv79RnYU2v/iU/48B8AQRAjC58m5kzpEjLdwEZ+wfv+PXMhMfBa
iDb5+631V1czk8loYwEBJSaIZbvfoLe1BdTXcwzzS/YvI9oCc5oPD+TBzAIJ0yndTF6D878iKcpN
64lGap/yGPQQpflLjrxT+wXbfQ5Ieanrj7vu6//gji6MBaJLf4fzCk8CJRXfwlNv6wXrcc7rjEDQ
tUop4IqqJDYYjiVswLlU9EH9vFNLe2KUgwzQZmbRLh5Gl0Ee+q3ZHN4zs+oOlhlTxf5WJELm9YUk
ZtyuHmZHi/+VC6GXuntf5j/2ybTT/OR0cu4pKxnY7msWw1KPfVIaZsl+1gb2R5QWyCBhTGFcBF9+
0VI740tIvx3G+P2UK75mYspvCkwv2swSPv+lnajURqBrBsmq8Jfu0K0k+owwDttZ3IJMt5KLnluP
nRG44/fYo3ylneQSxGvvo+90mNXuIKTYp/eeURlGSTOYZArdfDNYgM898mlwO01bEnM3XZc5+VYo
n0Oj8XqPbAcin43D+MsGjPkm1BsasBgyAonKvUzapZBK3jFVbdrhqJDarI9mLCieNkI1x2BNLED7
TogSjPNll409jlWfOZHlUvdm1yQ5mKYI2H3jEYy1uhfxdNcMXSVmt+0JRscXZ8aEc3mb2/6zTwwa
jevQLGG7nq2D+8icqSUXIufWbzZZw+XOJipSZdiCkS6tQq3LhlBQ44/qn+hac1gQmtmXeAOhgAFF
hIvskKF9EsgBfhVmCO8wY628+Zjrptcfvtv05dX4c+h2ZwEh5ykPcdQPOx/WNWZPKXCSSyJGQbnK
SsAF32yVDzee3o4tYEcJMoBpUTR3IdS5E2z5ujLtr4qy3GjawSyjzCqeyP1Gab7YBSWk3aKO3TMN
FloAF0Fmy2UipKO8O+I7LAQ9XmRAR5o/BDcMEX6wHJPss6IF3XFegzkPsvq+Rr7zM1dzOrcQXynV
dHCNQon5ggU/bXp/mFFT4Zi0c0Rc1KPl10d9yVyEPQXdag9VL2JEszNhtTEDXnn7gA7gWbmkdIs/
LhWna/TnknEYgekmN9Q0wgxCHdjub6AjyLuXIreMxDjctGIQUKM2XUCcclyRmpe/8A+OqXrGC/Z6
UuknzY/WGGUMYu5dxfvgafbvqWC+OsnwDrKvec1+9YygVty1nGgmXnJvOiTg3pdL+3A3IcGSTmk6
C7/Ducgijm647DByOkgkFEY68hykh23AUfv/M+BA08vNAfRXHabdiF17nHjP/k5EcNGB3LIGTgLH
H9Zupd+IeOQEjl8L8gr3+ejB+UhSD9JS+1X7zwuxAqSBDHwJ6CcLR4vVdamWsklqcxWSF3TuHakv
KrZucgSTGAo9rGgAdDE1PEUFNFlkEjpYMyimK38OyQYXD2swXRc8+98Z8sN4CKz2jvqAnJBdee0e
0sHKrN0IivSC0jRRJXEJDYzi6EqopmPrZJQC2eDPIgGU/xPDhTLY7wGQkJQGsknZ5qPbqjMj+Nw+
Z4IXHDtLnoSN5VjTt0WHvBly3VVyYp25zlIheKxCStAy/gVMWnbATbxPkRCGClxzdNMEjc8xKytF
OPj/LdBFw51QtKkY3wmbjAARs8w2jGmH/Etul/6DJ08f8+Q5nMOu5O9FepJdbYThtf2cQe0sgksW
eIzZuPzFeA4h+3wgFa7oHRowED8ONPW2sFI7M7/5x3qwGk4Uj95mwFm601xINes3KeVS8R1eCPob
Y8ipZMcPigwS74y98N3h6ikSK8GAPk5HRr9zJnWrdnihRZ3DmhJ7PmA6hEs1U8joqVHYjVTFE50E
W/dNLD5Wn4KMnkFeg/JngHjVkGwTX2eAXDi/jBwpWyWvlGQ8Od0nqIQFbsF7toS9R4VmHPxGLSp9
WlWwvCT/s90OY1a7dJq6PivDBvvlxpr7awOSpR32TLTgdinab2DxH0wSPHyqfRmyGoihIYwJwYpH
qT2LsQotEfhTNl94lqhTP9hvgveO6HYr1LjxV74IpdAmjE3x68O+nHN+mO80HM2qPQOWIm4rzo/G
wXa12OhCL82lWPUXcc1fGA7VaaQZbCJ298A/xlhfnNs919NV35tPhL8rBNX42UvYjza70hmUEI5W
v7mGiZUnFzub2Xo72Ob82VJynK7RxBMsjjQ1HBG3qyujjLjpz6c4uZYE0AZsXQqjWaZaEVavbaiH
jwCBILf47VIl6jtmVkWbpzNLvIigHVg/5+tn4GMuDiGkk/IyiJ5KVh3+QMVxMDW78OKPPf8U4gqf
UMC7HdW81APwBA6y9HfaRkP6pAfQUa4mHNuSfvHKPpMwVH2eRMIaNsgknP8rKoXYxc7lBrq8EGwn
hZnQ3kBN/oY3XjdjB5Lk3VcLY+HelCUNRLfEFCnfiEl9y1l8Fb0oESSwSOerllAXmQc5yMd2q1cS
gLa9qa+a0UC5+WTYlHKI9IiyF4VYCyjTY/Zs+WckkUzY4yfpAiuPhc5Uxo5WID6GOKGIJ9ratU8H
FV0m3iOPSPQ0fjOKZGtAU1VTb2y7TgqbScF4MIp5SS5kUsAm9MRwu7fi9lSPaNkCxs3sa21NS182
zoJZhISeuJ1ivg5jwatf043DYP5gqLlsNeGNpbgRTQ29kdwZGqBjgnnLAMzsRkFDpsdGJW76bYl5
RmkkiOCPSCNd9PLyzNMAFfBPfq0btNXKW3PM/KlcWI56Z6ADB/BHHzMx5KygUDOkSb2P/B0RDHXJ
m7VehGkmWcEb4E8sbED7NFc65QDo9aakw9t4yAlu5M1YnsGM+lOYIAoCbG63qoJeKDvIAUStzgX+
9W6pp+XmmkykBSvGovELMVAxnE/g8FtA5nKK/y2pMQGz87r/4WCcazGKXPXZ/5DW3rYoLiUFygbm
2Igp0TvklWhHNiR+fy9z0sECDooawWssYZTiXU0MlOkS5jeWRCCjAzL61M/wKuh+TMrOYZboisaj
t547Ru+4It03dCNLehNml/z1i0jIucG/yHnSinbJBRjKBqfhnLYwvD3NXvd05UvVEtxV2lZDrMNw
bmXur5EwGSF8G4i+JHbRRxEgq8vaha+AkVOOGReqbyru8Oo4sxqBZcvtpei5CE1H54upMY6yR7xt
SUo0Q4K3ZS/9/bS980x3UNVPmbtKg/o1owKrtYXz9f2KA3hhHIlP2Kjn6hfoOXsriaraqVmgwNLq
B55B19ckJxaGdjd2SkCMsX++rnkHuS7DbLmv62cygxax67AJ7+DvqK55zOkDZQFzdtu1TzvoTosz
bDbaB+ciam/rpu3yashpsMA6CeaR2Yt6X99/Gi04k55YDBhpGjwfWWsz6AKkOgFQgZwvPvYRDB5W
ZGoRAKnaLZx+mTGPYwfSu8Zmb+DxUoVRY1zLXHEM2Y3AKfNE/1q/OIOarVMmgyQhwZYChJbN76zf
4ajzJKkIszA/SxL9jEeflrIsUXGq/7YrISB8XJBu59kyUaQVZjPf3KHu8zeJufXNU2DEb9EIRb9g
+o8tMFTuHG0dIdPBTMlkMOhSLZvTq/IX1Nba7r+Gj9AGW3M03kdndYXeEYLEyp2eAvkg5LuC5cvv
eyjbiW0baY9wLFUAobyNtC+xUI7B2Sd8GVYyiIvXb1uyrqz5d4wuV+HoO6EOCH+3aVSMNAQSVPPB
YTnxPWkoucMh5c+1xkUH1v10CMdTy3/OKf7lYiSxXObH80/Po+58ycglk7tQxHqbADV6gSF2Fke+
hIPgpw927LoLLV+yr4R0E9B9LeZ4WdRgDKSETWjdO7IdKBFMvjK4n3nQyzYwxcaKDIciEk//UraM
lEPi+9xpDIxK9FcfN0F7NtY4Wu79vWNB2JksxIjM7YMXcozXYfVY4g+W+6TQZ6/wAJq2qi4Zz5p1
Xio1yULoIMb8uFPmtZrhBgcUV8Bstk5IVxtbDfasHMxFACtaDY/che3UnGxjRy4aoqSs4x36maRW
7ni1YEcEY0baYYsgZikCJMioXyIuf7xZdjdyLzZvr+AIQoqQphuB6Y96MgtRc0KmKJBn8IP4xqnK
k9q/1J+gXBTcwqb6YIdiC7cY1vQf0jefwqyRSMn/KK4IGNm1V4zHZ3ICVaGboXRLtYIPsj8R61XA
uGTlmW55ahpQ4eXRkAjP6ZauoRrgW/KCRXPaQchZr94fOq1dprj13i3+x9NAMAAhFDX6TPqRG7kd
GTHpX2jg4IjSl9dOps9BM3Nye3tbpyo3jx2EmV7eQuLekiK2ZIzb/cPs9lsAy6+eoOszj2sKt7e/
tVfHom0JfYKbQ0n63/CF3ZzeCnKDmrBJ7O8ZeJG+XBETA+LKmf0dz6CZT8u1o6nwAbznKfqsgaMH
jmLJ6H/+1IMbnc1LIDw64up5NnnrK1mkTBL+W59wDp51jsIc7Pvhyvx857VWoeCCR0KR2i0xMuV+
QhtTWfORy43Wduo7Xx135V10VJHppQXevv37rVJzNPXxlOhTBh8a6ZMSH841wrXXKi08ulZomdXl
iEf9ejoSV/jGjVmfbNIw90CtZ6lIZyVeQNdCyPps/MgfBZf/D/S9LaXlTo7+zOlOsHGVrTRNtTGt
vb3K6jd9S+u7noTHY5eZnY4ghQY9xOIZ5+WiTfebhrAe6fjPtufFjF5WE5oMRegF80FcpQi2uzar
U8jkI1exAwj4V/UYK+qkzSB0jYWF81DvShTGPChrkioc8KvItjIx20lUhhaO9w8JKHDrKFzRwF8L
mzkF7p/RTcy2UnJ1YAMYmGgnMwcHTbfMSIBR8NRMaGgmSk2qhgbgJV8F29BvF71yO7OkQbCG4Voc
3Y1PTCzhOsjx7Qa3n5mXru/FIa2VF5fXvlf7ety/lOf/AX6mCfZ1uBWPxgWq6nAAndULDgslKsq8
3Ah/hXS0FIGQeEQ/KVKtvHbZqSViZxAVFaKAmUKiF2/1M9I2TTY7ZgB0fMY0PEgGq+SBFbEWPcvg
/QAN/J330N5zPtw83gHHUrUUNYTFHSuKPBuEeIsW3dUMfJFumHMmL05SSMGKbeM2EuHxYAZ01Jbk
tSjMaN7+X6rIJBlSioZcTer6SwAFb4PeVjo+KfJmVzW/iCMEALBuslOojbzio0125v/bALYsX46R
Ls/t/JkrDNqhBVnivVlUGCIL0JFfE182r10AwaJaWv82Vvea1H+cfkdlcKxONNNwnYw6VJlrTluc
miRM3JNgdx7u4qKHf3g6uwvzwTbuKcd5JZccWalMUr3CfkeNwGcw9Fm9BGbBCJAeuWBZggbmi2eO
6B9ewFPV5OoGeh+rerMb53Q1FQXZkC85zassLu/7euIM5sOurd+VN3LyMrz4ribLCGkPmFOKvHxN
N2E69I7scUD8sOTuEjumXZjqGeXvFNOGd+K6SgkWUp2QPQyj/Sa26KY+hhmSSdzN3Co1UfN5d8UJ
B5vk3iMjy5cdnp/1IhqMUIfE9UN/LCXdVCmTuVE4/Og5leoycMA8MtfJtQfxxcXF5rx+DhmqXxzC
rtWvItr0LmkOlGeYbXt9h1e1q/RvRuJgm6tiNO9d6DRS0MSYCCkolTBszKjZMZS1gkreVqz+4YVT
NNq9kUO2qYGZ2uVwbCThyEOGfIzjapZM0/KNMJhQKU6226CUxL9ABDaxqJmc6WeqKhVhcIkDcaIj
bq5MU+hJmDgT140VaRU0ZG0AgZl+lnmcArHXnGniYk1n9lC6VBP0LNUPdKn6HiFx/vBCWvcH+xdv
56WI6dL3PUehrrRUCg/gbDhiZq2j0qv+0655otBzZjRjth8yibeGaeI2oRhB+9VJNKH8vmm/rGH9
0MEU3/UBFaYzJIJ/joNqbkuG0cyGYnRIKgRIFKdc02OghzTlbsXVKzgsE0/PyYR6IQXllo8XakAE
ZmWM7X6VjINyyrvgyzUtm/SQ+X7lCfNDolJPHCUaCBB5vMAtjXXZ4M+S384WiKffE7S+fy0SXtSN
Xhp/4yEiUDGQ3JUuej7qNEoI9UzGvPrAhGLB8YwbWjhD8vEOJ6szBsTlBUfcHEOlFQa771jVR/Fc
IdX9AyC7eUyZ5Gh9/fRphNRe5SGVomOFR9mq3nDhqsjtc4VHD8XNeT/UTg7GJgpb+ha8t/H25cLG
fmFoc8x7Ild4JK0cmUoj16+CVbtyDmEmm+1YIoyCXTK2S2zJ87rcRmr6popot1E9SCU+YDGIuODR
o1WKcQSTpS0RWGeLlOFqQmUizPYSXvkmY3TAbzL2L9CB3j9OJvOrF6Fo6T1fd4uu/XRQ8t0PhOLN
N6/1yW1ekS4Iwf9yxbM7BMQ5B56koS5CYLMKc96ifDQEfVp0jkQvADCqA3zbbGOOjKLfr0UGGKGT
08jSIB/DqUXq/RbSpDnnjj4KgovsbC0U/NBxbRyDdieJxAXXDUAZ679CH5749q3U1ri+afgKLLa8
bbakko6m0plA5GIrd4Iyu4zzcVoFVW7rTp/uCkNSB/O2lbfdrOv9uIBHH3LSJwlsp6V+My8tMUW+
AxEv0+1hgGB1RFnqaVcX+B7l29baYC/Gvg3WrYB+dzaKUh5yIv7XNSO2J1oMoN2MSG21CKXIaf6k
wgk8NgxofA9pyMAKQXzHb4RDw8/ZDj4hAcDGc5krWfk8mM0VfBD75j82CDyXcURhWgHuA7Yroa1w
2867wr0dO32Ibn+HVJKqSWJjMSIHvJzM2eo/KEtdGPwO8C7zBtAPp2Gj2pb5KHg2lr7qyFHt2TaF
//+vEPhCsDKwbHC6KnY7Zpl9qzJXAt/BdvF8mgJ3usdfHqrFzPZUYbBQnL3j9iy0HXcbzkzrCNRY
aAz2MM5HFIBBirBAwtrFIZuk11SYMZrmmETatKweX+DzSeHKFjSc7Fsrdknc8ebog63KraRQOYL0
Vn95g4jBCwAMzT5M44HApy1iazQQmrv4GIl0XCuJ1+soXpnA+89qR88rkP3Ib8WlsngdpgKf0kkt
VVIcMlW7Pw9UzQ7XCNW1jpS6f5ybybOG8UdMxwJcjRgmyPGrZWLMLMRYLifICRIgbpq0f4pM4PxU
YBaY+0Hd13OE0ErhvyfJLSLIKHy0ejxeMu2rGRHSAP41VsXFTJvMWhNLaxGnWyO4u975d9PDt+jQ
AdHXk0k5ZRX/SbliWHTXLRsDJJe1Ibuls93iCb0rxZqrXekAOLR4Pqov098CuLbg4IEA1CYqakP/
yoO8gQVKQTP+Z+dBY5zMJw4e0c+8A3U2/el7zlwIXLdWO/uj7aCFtRYY/RsqBnnbksnhqwx72wyG
+n0EZIrF43XcXmGpwHHduynrFNXT6OQ7E3mnT0u+oqDhShk2Y6QtucftQElWNyvG47ztzEdCxAjt
q5cx3z4EtL5UGTVu4oDyXU+lLvUWDR2zAspeIs31hq+K+U0szW3SJFrNdJYyA4GETVvb0DzwrAx3
hVNxpPHPsAtkwE7yBi5HQ6J3b9q75qHLxjzyefrROMf967C5rTKsvfvh7RI3KpGlN9Awj4HUYDtE
00KDuswj9lyxigOD7TDUl6LwxEeyHnkc9lwncn4hQN4JA5HMp7Tq5OqDuuwQLLB18CIWlvg5ueYo
vrLRDt28pSSsHFZDOfSloxP7gpYqTUUZov1nufb3+R23XQf/UpUV3Ii5nfy284FgEXKW20IPswAG
fMqjGtRUFD2fv7MUSg+K987qRT3v628gySgVM+nf+ccE9UdgcYxA8ZJMIxg2VMG9cfbenC4IY0eZ
g4AGy6i8Hh4WlUDCojcdy9YT5/b1XBefEDiZjGsCTn4FARE7ncAipJDya7cuOjNOInDc1bxQG+qg
VpEh+ZbO0JbZdAQYi9Dve0a8Y3nv+HuAey5KzapNDfMW7OePF6hh/ClWmIdzcuK+42gqibiDO7op
cUpANmagBVPEt2MRw6Kf4yqMZc40GA8HLOrWhQjZ69F7jje0Rqcw2Mp9KsM6DlKzTMjbqLfdx3tT
NwFiKoMqOc0Bcjw9lOR5BYJkI0splZpJsRnJclmAVqnyRgngZmORreZZjCi6hgXez3vni49QDtM+
gf7/EuQ6JevwhLOuR8z1VcMiHiE15LBIn7poFVhzYrYCk4laNZXD8gp2l5h8h8P4oWL4HO2CPz8m
Mk2HKYGVDKQysHDYuHfpInS2QCkkWWse8OUQBmBp3Tb/72Wn5dyO1+Ln00HHtGgsl5gjs3oGO0PO
IAeFngz6YKb302ux3iEnZJ4O1HaNgZXa0O9QQfzlD6C9onN/XUCySteYDgijaLGEdPPc0+7V+HYe
hEHHA5nDNKmBuX2RBS6vaZdFN0+n6XMKbT2JCv/CO74mcZhWRZ32TGzpWrrZn0gdIsCQgrlIjFJZ
/b7Ov7bbv2Ioz+1+vr8xFPmL2cMv++Chb8/Ga1dLKy6+hZN1IrEQjwYuYoRyKzkzJmXm+yrpjQae
ZH6MOppzWzDV4rybj2MnSMMcowTfb+YxGmsQEW3DL0eiQf0OUCeHiQzhfB5V2a4Czgfku1fc+ogg
oHWqzkVpQZJ+f3EkOR+3H6QP6As7xEIPNPufQ4eVgtkv2DM805HTaqaTpEFgQTv5mAkZwYNtW3+F
c/uvngPDhlifSIzigMO0nnT+LaacGPepVSbyrgidaPlWzlwSBVtqHGdqTViuIOUJeoL+OZyQ5ZXd
gWnl1ucbVgfLABWFWNKyKklAUhNrmKcfcIDceaRUJtkFgJ4TEwlBIqOATqixmRmOjh4UNir4xXXn
/l3LIdJiw6y0J77Ak3L1ljQ/bpm2h0fvsS5WImGeVqM0WnJwRARRWGcI/8dDtkXCtXYkmSD/Vq+I
QZfkHbvpNBtuRiBZ7Ik7iqBmcFm1q3RskIBvLRxJt9I8R87WwGIwDMccUYxmqLgmzWCaVVsZ8p0N
sobcaLfDO4pCeVNQuCc2pYjCGg+YKokK8vacZFk3Ms8HhrZ/9KED7bv3nU52ZF/gYBQo68yfhxj+
FtOIIz1OsDcuyWcfw1/u+8OjK97HJXO6fNT42sjUj2Dh/2eILeQ7e7t5EaiBD+8ceim9dI/7SSVF
YvuhSmkeRXU0SqWzIzy7BsSiPncclqpIyn9PQLF7CzqvcnHgqGV6i6TolZ2NRF7jqaGZDGrs6mgM
ypmRe3KCaRcq15U4EesqRvU93xC+k4/JCDVPmF8SNIIyp8Urh7U+dS8xwTRhsRWv6wQcSx5LKiEF
uq2j+TSm+zao3GpkoU+pyUMJX8OpxYwQqpU1x3R9NsTU/Qka77PLShs9lDRP3yMojotxYLJ9QOJp
cpF05lu1zZTZIxm8w18bMbTnsmjPZ5h+ICft/6lJeFOMq6IlqiWAYxS71PT1tbtBjeJHOhSaaXcQ
y7WDw5tizyv3EwS+3knYjyLdWEGJeanCUAT7OS1YBeKPSRhB7+Aidbt9e5g0d9yjQC0EnTKr6Dkh
mwr621cPRVFxBKxcD1SK8ZtYrBJ9rScPut0QT4tpNlvFj571LjTDqMlVbfTBBdw23nvOIUwFUVe3
biFk2MlfFKFRw4C+XJHNH1YAX9nHeUUogxYQL8CsJMKA4OIq+Jypsyj62Rz53SnkakPaQ2ofuaXC
KnCc4PjITN1w1fQ1Yyx5dESgDtWhftiOceylDiv7/rBaC7y5NBzntpb/Z4O3LnzvX3VNF56qWQ4L
sbyWTrUONLGkCvoeNY6OTuMewHTq3YdIIFi4+wGMsnW2TTLmtfREUqF+l4ItKzegbc49ZEBYAzY2
5YIuZt7pEVxJ/vfhQHVxdO3fa7P3fYaS9aYfCvoyyZdzRYURTvIwdbgNrwGWOLKvmH9+1d6Uc63h
RmO4/bs+mYj2rDfok9T+GGbjk8xwZjG9rXdGcRQxh3tmN1TxSTSu9gvu9izehv5/5DxNjb3BZMq7
B+WfH1Cn1Cw2HNZjZvLZMgGeFprTKPKWL6Tmu9eqqQzAjaA0TF2SYoFb6HMFq3fisNZl/bAv8uom
LUf6gqdhGb6Lax36k6D8VaO5jRAFqsQnScGloOGCiP9CuNjUqC5vVntcLAfnF4CmNF2if846WqRo
O5L0IASgx4VtJPPbvSPbyQhQWhEmEeyquFbThV2QY7pCv8QKdW0puAc1WDAOLBojWYLgtMqINWan
GS/8YnC0VV6Sp1bh+LDIQZM+qmJHjI1USs6NB0cC6Iq7W7cjOdqm3VS1MXLizdfGfhJ6lO5YiliB
WZtsDDbg2FucEbRXp1htU2bR1/QLcP4s+wCppX/0IxDCYeqe6uE4G+cmYId0OqigCTQ0lo9SI4wA
4dEyL5mDJINfSu21AVoGnt2/Q2J8aUBlYjKEsUUm4n3cScqsPkNZPqq+eEbEGIMGD+YIUhMUh9pW
92t/tYo4RvaXbkpirUZUO3+EVGjxZg51GMgj2WWTBS9cxtlFpyuF7fW7gZ+StSt37z1eMiiTITST
CSVA5x4DtFLMe+DVL46Yr2+d+Bn1dWbyPyPA5V8Ie60C9NU3zMp3c+6iePiLfiXRwmqE+W6kW9FA
0ttLDKSCFs1sA+3Ob5IS3Pqeqj2y2iyu0XQi5q8ghsRLnhaYxuYWJLqMDDwviV8lZHLPH3dLw3wV
nKqLMXBGRMiUWlyDbrBq0HUgf95vIl6lzCbzGszk0SPa7yFeGjXp3kt4GBPQwNOdko+7T+poITc4
bewF2iMazbVmvJFbyLcRLheoPP72MaMopTjr6Vbrn0aIzLQ4AW7W6/TffXfDZu5BgWeIRzCAJXnd
KIWrsgT9uSWdv3/GyV7isbrudUI/4rJHeEjJPnH3olvmxpRTnq7hpDiQ7ldq0wyKSOJ2uIG6zS3X
BfPMK0nkXKZKp8hL+72KCY8D0NagIEFkUjI8cexGojcUOrGBZJYRzeuNV+CSegJ9NqhMuzgaluWm
ERr62PsQrlJtRA3eUj3glj8KDHd1duA7KToayd7yLvJcxZHGdmnyo1OICnbj9khnQKH3H2r7cm6j
vRqHcbMiQJ84bqxuw3HmY0R+05SQu5IDyosoxhwicN8Pf8BEgh1SsB4SmnXNuGfbJPtxgrlpPHTk
4o8PlwEflA4o6O0AUHu4Ydr6LCpltZOffn/lPva/IKTzCc2oNAqiS5jv8ohENCFrzk6Ls5ZUXsTe
3Rs5slj8MSS55g6RBbUqsg+m1Jk8UtkZdK0evXTpj7z7mK0qF+6UCIx4rLfxagJPRKXKhDd8rl38
oAbGoDWWDcckZDu2k5D4bR6teM7ieOC2IANzCVnspc9INJQQEh6txbOXBsXTPoqFPPqunoDQigJi
8pG3aZTIRnaALxAufPBX1hqa0UiE1FghIySGjDK8UZqLMrA/M63IU8YdieUbaADHMqCsQMnxBZWW
GF5zBP9in94JABnLDWOVPTX7R+TbDFgZtC9/xnATD8YDtFwkzjDy6gXkTLVcIHLTupZEo8tB3k+M
D6QttvbmHruIniSW4AoNWjEunRYe9XeYVoVNRfPcKPQcSHF57uwzLz561rtXsbzqzHLzd1mk9HUj
VmgssnARCH8wxSZfFw7HX5B3w3mk4zgikRHdiFOCg6Vn5iXwnFhT6RQrbEJwyZ4msjAlurE65Ktc
ydKFfEj8k1/b3qoJpulxwWQnpzfSm1XynEH5P3OrKKGNs0Xs5qDh1qv2xBkjf83BqJ+GiMqHHK8A
RmgJu8NVB36mOBBHxFkGRzj7aHP9auFraQNLMt5XJI84jdKUTJ1LE6Ig+1rKBNo7DjmmV1bhhlGK
hiACNFZmB8nNZsgbbAbzBO0ZGJRwZm2bqv9lZKJ6ZywuXi9F7ldan2fEp8kc1wA4sA2pmIFd5fXV
EhhOve1AwbpTgvU4T5osyavQQoXwoKYMCl4luV3FWpY0uGy4YvT+nmOqFL7fwJeMfYx0EWMx7jKE
kpa+1N7id7I2UnQ7zPqAOPLhjE7Rho5grlPMF3Ts+Ts+IyoEMamt/6nmPdBSq2KADPIdHPRGI85e
Wurlq9pxFMrOd3Z09Jni5QTUoSXDLjttS4CtsD4p92QKOQP0oARXihbn9zOLS1LTYuPSIrIb/ynR
ISOb8cw18Agj9ATBQ3wvGGmjBUDnw1Tjc5mCrJMvoTi1ph8oerw9nLi8aTPNoRyMKgb5TdS9RssC
4N2nAm3hDn2GPcorcbt9b34sboKVqrwzsj8iFEVEYRu9qxIymxdFATgcYlhNpMrMSo/eojGVGCl8
0FNtjRcCd8dYOLxkycQXxkNNnSCAaxcTViTBU4ui3KQ7FAEfs7w3yX5IBOteNZxwC2FMt5Vih0cI
S1ZGrg0g2iTl7qzDuUsRhOI9cYfqDSY6Io+RLoGjdV6SOnyczNy5rmp+z1jcn9maeRzjvTnYB/KX
k+49lHi4t+wrEIr6M98G5rQ1PgblxdcrutoG0ofz4r1Z//EGP6g1yYsqu5cWH0Gn5MkeyMoyw8GF
BqItPuL730MPUJIirOYmPTBEj2uYp55+dsjfBGyBxoHcDdlPZzSvCVhuac9fOmYcL3sTTT+J3yV1
4CLmdWkUsm/QdPbGHrixZsERUFl887+Ive6kIWHTvQ28r20xYiyb1FMXetXuqfSARpe3z3UgC4ZC
ANYPBUsGGqLutH4/npY9ySwLdY8CyoAt3LsQjvTTG46LFB7BYnsrSkFh6/9lN2iugup3j92THUTX
StGu/3MAMkOXNGDRBkgBbaJOtK5wudgggo7T8GXTyMtIe7U10gXbibz+EQcOzbbzx5J9WgUVOF27
mSShnXXEeiZWqB+46cLkegizbD2X1/ViG90sP5bCSbOmHJKSOXlvAWfAVNOYApBfHeFlCZSAAaIg
WGlobWZfZptyEw0SiU8lFERtLCCj10pFhQhwgik6Di8TYPF4csvLwdnNsr+mjVMv4VUdoNfLTYRz
Hgg/KJ1OaNBrER4Cz4uKuH8/CKZvQarJC2IvsgdiJBjCFl0l9g0/7z1xwgr4NssWaIqB7xzDeBT9
ZF90j8M5csuVsqFW4bhazCGfWSHafVfLW8IjvnwHqAuaAyEIQ73d54X7A3twcp9/7u6rE69TtcLh
LduyoTwxsSvbdsJUIsiVB62R4Z3Cbr5CsTz9DKOqS7UYNNHSyqauZ1PFrw4L6u3wff4DrH94gXrK
KHlTIIJkA9A5K87D6zDbxc3nM36s3hmpoweS3vSo+uC2xXTBm/zdu+GjwjNnh0lNI3hBsfN+paf8
kkZqM7F3yPsoUVKvI3a5Oc+tpNGMMTw6dsEfUgv6KheJFR9lLg/AyaMg9xoD/7exOr2aw3iboxZk
MH0T3D3F6bXhF25N2ND20QcHkTl1+GhQ09sH46bZ1qE3Yzo5wwlillWPx+s/+URv4v8McRr7AHaG
vHuUxOKPiH5S0gbkzG+y6kqMfzHpMIghIqc2JIVO2pc6lqD9ba5u97MLyA47+1r78FtN+Lu10SJ7
W1EpVZ+IxLOzRhXsbG9JTO7ARcJhl9XDm6B548YCwuyfCtd5d1o/Dwf5BP7CMCeeDCAp8CQ1qSMn
bCwM0HMkiM+cMBHekmaT20KTYzDXdnP12v24CjIzjkuraG0GfBROlnvG6j+fYDoVMhgKYcoDNTLx
mCfpFzPVZBQA3FRa1qi4Bdk9XFPCqjsTjhaw53wqnEncRK/iiKiuFHvH1dYSYpGrrckw9ns+dcZH
FswmHI71NRM8lVRRmT8jiWjpO/PzyD00xXJctThlA4LmDZ28vk1Zxv0oajQ58l34iYcSFciBV///
beYV17GrItrHoq5eh5PlUD+m9VonVJ/WG8haaQak+lW8LzqhhQgVoyFySSFZu/v8/ACbYBw5XX+0
4aFH/LJqIdCcghE6vN7/bbzv4R0AC5l23Ccve3vG8DGVLLYcMfsH4+9DG+Ony9kTK4R1WQFvgvFv
8EpoYd9/AqJ0FHShQVehjloss2BTryhFmAp8X0FWniJtQNaRImpzeh9o851zO/Fjn23LZOakRJcH
mgGLlwGzxHbo7j8b24NZYJ1d2zbVxYyLH9rSbnhd7qogV2fSOyyp6J9TjKd7VWBV0F0nbM4xcRCP
kj8AhumCNNODoBlHZzxL92w4tqEiOTwxuQtQJwqUFohQk4ZqzX/2Re8BjQM/lq+CIOZrM/cb76o3
xISciO74hXSw9qLPJ66SKAr7TNypN0GLpdMWLaySO/smNC/0oHt/V2W5xDCgp729GgXplgmJmOKN
vHfjjemNBlb23e710rfqCDJ3n9x/cZFiv5FzhYAv5mDrU01ZWdGfMEzlSaDYpGt9HnPyu2egnraD
iW6RQb9C6jbSkRmLoYaWcI737AFzdrTpQKKE1+1oSNKd6s6YJF1Eqib9NLaU0JOznhQRNYHG+S+g
AOV2lUeJqAEskwJoXkixUcqE9/K+494vYLH36FqotXHm8J+fW20Uo/iXfYRLgEARsyaWCTQLMWYc
YjQtrK1GtdtZ83s5WRjdx49jr1CascdUtIvidv0OwbTMXy5yE55Wjapt1oHT2RJRtGt0QMGbEgA5
u6BCC2GsnZ0IVi07oJj1vI4W6yjc1/m0XO3mAgHCdEYVq4avBtCjSdJUzHMachHz9AUoSgXhsVo+
ScU4yP+H9HiP68sgpmF0Youw5lXYsYoMRBpWUZ8u1ozkuDvBj81i7x/28fYlSl6WadzYV6mMdh/X
r/BuaTQLDMNgEddaSwJ1c0/qusc+J0cWh2tLQa+WYQB13CuXUo4ZWTRSo3np4WnHLIdninZAhnoW
C0Znd8b83w+pM/gVFdh2SHRRFlQZ2ixytKvwiQSqt2IspYuxfCfFS6YE/nJcFhFMk8RLPASIiYXp
Ukyp4gdIoIT/G3h96IereAOcueUX7AuA755BpWVLXUUd3u6J06PzMAQ+D5zCKy25EufcJhxMlSWJ
Olamx5z8x4HAff9c+Y9Vr1KeEULBI30sbOmCcJ70Hx/6PFKnVeHfRFSnZRTjIGnHEa6DKbzvpsbv
TqYFsJ7RxbPO4e1G4Vp9plz6e33z5g9vx54eAYeYUzTlKEq7FyHQVTLk0EKF9VeHVBNPC2AbGLmI
2HjTWFaQVUFS6XNzCUlDCnzzPAMQ2faHa//zWtWXk+W57gXLCHI0fDl8KxKAuW1yMyozXeArkOfO
VJmSe6XkZLnQfumhvgohWRZDWlYCKgICEXtZalSBugVqaxOtDyNPBe6lBVJqd4Z5bP0NiavS/jez
G2INOIsqSm9zmQCG1igGbwVcoTtzrPXFzG1rCsX7MXX8sxyhskHJawsK2KgDGmHdPxLPFdXc6l8d
FuoK7voESIrb73Duzwq/ERSRySsC64wFgJxxm8IIyl4SnFVZVUT0Y4+2bAoksPVbRdkNQUZCqy66
EbZaWgoW1+H0zSfnFy68f1VxWok9Rbva/Ky3q/2+/yo0Ad70eGYHasZM3aUeXFRLKjEakWBJV0pe
AJjq6eRbWv4MFQTqr8nWO3tjja1axW439edJdA6QCj/00vbSuiOpIueCpgsGlJ1ZKyYGOh7jjTAH
KTDKkKRyi9fzNJSUWmdS9sRI6ClzufcxZA5y7k4CGQWg4L+CLdeK0Y7lp/dFY0arJiiMN5o1Xrnf
SLmEKodi67FXz3SeamGV8iwHDB2WkT/Gcy6yo1lRWFwwzikkumLtoAqfP8gfkHG9f73Pre3UZB5w
cqmGY6FCbaef9WHR1oHwATV8tXIbW/Ja/+j0oAiMh5vgLnhNZLHVCaeUv5EokOteXwgHgPnKKwkk
FokjGLFRIbSELFQb33H1xz3sMV767tdH47PxFP0nV1GZZzqxXBSOyNq9CgBFm6vWPNBE4PE8S3i0
qpyew+MjGLQZ8ByDIRyj+MtSQvuI8OLKH32ylbsmJwO0rzFv9WLWTuCUbea7tw5023hjtvHzcdJb
TDxpew91m/Mondy4FRHQltSn9NrCbTVx6SZDC8AnK8k9IsQIHvt09C+SrW3mCE/8W2gphu9uW8Wg
8nN0J2O565Q3grCZ39EegEs5ZG+EdlJEz5y8/eKREvmEooonjbHTj5V6zwG5O/gAjRQsPCRUBx7u
SlnU7Yn/rB0/GT0TDfJnWCvp0tBwoHuorqbPuf3E7qPAqRWrUKJzXUBak/yAMHl5F/JgAESE7pt+
/v1xCCPk2IChAEQgSr++x5Oevn3zaNfflXV8pV0KC0jdtRcZkbDYynFpelB8i1BIDaYv5BNoUiCe
u6nyR33ox7ratFt06/M7MtsFATUosppCO7pyY/V4tlqvD0Lfd9SOul0aCbvzVw5ks96JOsg3KhVY
IJ8xFzpKAr2fzbpHskPN1eXeJKTUD/xjLNCE7QB3J+BH2ipAeDYRr7Hahy+kjx+tOgCz6FU7e6sN
uB3JFjbbqyc6cMJEYxPp27lKXfh3gX2hDTuvjUAYd1MPy4WSkXQM7YXbggqjCaRrrEC6jSlYT6GB
D6HmzaVM/Pr6+p6ZcVq/beVOMHvBduwyTCBj/OSMe07e/DJ1jisSlRNpYTgbdEnIDPbG8Fb67pCa
eSY8ezMrfqsAwMgteTdakVmA/s9TZvqKKhiDTAMge8I4jl6lvaS3E0nXEGVH3UHbFI7wadSgj0Y8
F94gX0kZ77XcniU16ZnD+P3kM2XTNuqQ/pSA4btAiLNFt9a283IFPheTWmTuFCn10rx2x3Byo8X/
C7rvznA55HqCYApZZyKe0tEOwW8UTZc4/3JaCUOP+POtqeOrZre5UE2AyONLw1yfI2b4jtCTbZ08
bs0l2zOR7rWYtRGKAQolPrZCCAIWCWN2PLqKEpzwvMhRe+7kJ63+rhf4imQaUtiqK1xfThG2DBmA
M0o0Hc6oziLdl1/5AQzMCeBj2luGJLF+nDeM/90TVfggw9EPwEVV1ipGPLerJ730F3FaA8BqUSuz
MFD8nN9I9kyTM4BvkoIWhOCTyKkn6uAmEHApoGothdJ+fl3CzcuqgZ3R5wZP7hwpHirKe10zyG6z
OpEFjLgzoquTBABrNtNZUHs+LzVlDZ66rDrv/jvlJekJWX58dXdkLBdkYjCUq5AQXMYvHMrvoEMz
um/h69Pwa0z1NcHPFGndlL97ULqfpWRkxjNfvrfx7YmpAtY9SsigszYZ1J+vNUfNghh4Buod9o0y
YgvqQRFWmo9cOV7g3e49BwMZ7fMVkFlryeiA8W5eZnYOsoJTsJj0p3PaZ7uacpD1B0F1Fa+lBzz1
uGNpS4eqpRqKSJpxB+gkQ6RhBiOl0lQ9/kq5YbDB0YJ0g9bvLJ+bFzrj/o4aalT27pAd7LULuq+k
M+adD657VLaIRhCo+zOnm9d2a9TbEmJZrCtP/ZIYQ2VHC2XCAtcIoZEBbqgq140TnUQjAIIYNLTr
ywCfDwqe+Km+q67IeSo7xyj+bpy1BqG1SreZ4P1t2rjkIX5XcAVayhIFn3a1I+BHgXlfUaX7H4bW
1UIwjD35OxP1eOwQLADZjh6i0L/P2vOh1qurlkBA81ZIrGttYpCZ+7Wxw8qB9v9B8cYnyjUY2S2S
9eyQPiuATiwiWFBC6cuMCu4iOMsh/FrUGxhCls7HHLqhtjKrvUD5AV8cqG6QQF+eclpoUtUDiLAK
/IHJwLfc+7A+LenuKElBvUCpk9NrqVZ0zUaA/yQ92Vpun5/IfkNeVXm/S6VcxPlM3NEEvSsH0jKN
wN6qcy2VD4zfyhB2C1+LCadN4MB3Wvqve285j7whBul2HZr/6BzJX+qFiy/5DuJBCwEKfwaPqzUY
QbnIhx/i0VqQmjpg+1szcVzqKv1ixTd7NHIFeRORdikqPgh67yD9g6mz7nc8S73jh98/folMr2/F
X6C4wIdvs9HPAeGhD9C9zdOfPBSsKKciAdrguzpMGsGk7yQjI7pwKxVdSYxXt0JI0MxFxWr6F6Py
dTbGribMIVtayP2I27ZrMjwlL8/7HzMG2HF6NexHiL7elsckXk0s7HYahBn0ZyCYtFItOYEBGmuS
4Jp1SAep174ze6rBJ6mqz9kwJ9/FbshC/ymZkhtn+phB3sS+9QDiQIEhdtfnDMVR+Fomwg9XC6Pv
7p+8GC71yvNjhGuOCGf3nEbFAgPzqKpccQuxTsiSf93+EeC4JmLKV9p3PZXwsZ7N8cdLwVNs8iA7
9th200N59WrylXWA+zkagxRZxIEL3D0okkRc9f6elX1cmHdIkfphp3gMWMHW6AB3E1IzaKoBS/3i
zN6W9LZN92GCldPATavaSZk/35iTgwi+y8i3vl5x6qh2enCyd6qCOOCZXPXaxaMe8Ps6Mtnwq+7q
BGaCpI8mDN3RMmqPgwpGZgeCAJZWJet4OTr4FhD6UDcmak+uaBqReek998toMZ25JenSB+5WCtED
uSAtPXBJSk7OhIniFrd9UGZwlrY2pwy/s1TjPbbOXXZTCV7BAEXHTjcoHqPcsJ/QPqTfdQ6zsFtr
IV/TuAQEdhOWj5aZ40lLWfVruWqKUhCbWhQNFllBxvyxNAS3zLEIcNutSp0TaT2IZSItIYJI5YnS
2ErrFhswdo8tcvmeHNT46MzAhOv53U9keOUIrkF5gpwsZAeeenXoq2/ei1drvQPSG0+3L0b7Xhof
2Eex2A8fI5KnFATEFdzyyeLXgfaTz12zRCE019u+uQOZlz1vWktz0Sw122LebqYkYU1A2Ej9bVHN
ApHQQTSnqT8XqVr4oGW0L3zLEcio8q5y5v6m58lY83UIC7FzokDaNjQOkFVh3VDhqwiyh6ksPLcu
mG/9ls7CT3EC+RX530bd3RSpRCMRedqOZK3PPN+dtRnnMPCot9m9sdum7wXRxhCfcADHX6rkNR0x
X1P3l8H/J/reeaTk07I6YBV53LyNnPg9e6RF6bIGH1Tbq+dZ38QPGRJlUaQJn+o1ps8lGHRaknqU
5yzx6g9OHQHZa80GyN2mNnogGCHrLGgXRTdxqf/Y5A0cYMwHROKma1cQ9p3wH9XxYUMTp7up5CKd
NJx2Le56fOJlJR4JjLzGkW+5eV/q5LzW/22jUQsuDXOtGvcyfvp54htf/ulFrltrUgBsLYMyVQWW
Wa/otV+qjZILbnhSNDBLH7wDRGWnti3L9WTkJU5FPLrd5LWSN6kRzXIlmz7q+CajwJkCd9U/Nhir
CGusCn/ojL9NQpH7JP/dgJX9J4x9IS9aHme+41+xRvthgnPURRXyUCqkr0zX7fo4aBEEr6cdewqB
owyf7hErhVdmUM2O8PjgRsythxqsOmjZuPHXdZD5mWZtCjRQ0t7dNTMq8ALfLrrs7W54t6ULtP3g
OISDav/qAsJAGgK3aE8krEPPWQJ3MV2/O4DBchSnmAvfOU/ySc1p5biXcUF7doVSVyONASCPeSYN
ewxF8aJonDleZZ6XgdFsgoXw7ZDvhPB8YtxeDckF5dRVubK5XYrfuJmpeMVdt0IMXA0Emg8aoR0Y
Sr/T7hiuD4b6YiPyId84AFwDhpgEoLK0nsplEUrd3GlfdIPaWaz7HBxJgWUMm6Ci3682xvKj+tCw
3mktEfjMjSG7qzGBcHkfSbkzf30HowLSLWYVCH8wEe4xBmjZoKqdqzP4s35RokLwvyb297PCUBN+
LgpvexPmi4+92J+7wMcGXQcoxSEAUyj+pzEw4VIAou6p+/PcWs5jt/c4LI9+9Ojd3Sy/nmR8wWb2
VduCo+ljOXAL9SLUtUzmJ1fjCT8HfHecqZvK7TKbt3APBvmeADNsZ+O8mTMAVP5uNCLsq0VjgAbM
bHM6mMTgo+gz+wcCZjl2DTC99F8CBNRw+JQE61DbTrhyWHNyqA3xOAAbq1jRMHZucSPx6NJFP6Sx
wijO5iy5fkEv03qcGkbb0p4f4sCbNZH7iU9Sta5FF2ymJXvd3/6eJPP+aAIT+FMjQPw55ZqzgoQA
3vdQ1Ux2cQDiMKfMNRpnC/DXHC0eF49qXp9gttsMWvUW7guI0elf6YW4wuWs8G2KmRa0fyxFazFt
Ej1Sa33Zqfq/WCbuwzRyP/AHOM4Qr0zjR61pBciJIw5NIfKC7AZNu9tpXRVjD3Tc6bJ2A5z54ftf
x3/dDpSnBLgLDTmd4LDOH0FkxbQt+y3gns56Z9CgxIYRh3Mx9XfTRxVfZHlaFFtTyoJ9UBJcCl8m
YMCPI4w/AJz6A1OShNvCWkqih8nRHOmoVvZZ437Q4YLGcNIRmuIh/tlNbGSwRSWIxsTfAFrVoem4
i0nv+Y8tMNimUByBVwlrXzbCxDFOvqM8nFnvsQE62Rteukbo2ovQBE4kLNlIgtLzS5FkRXLlMbuI
Vu4AHIN9OzPQ1ek3lUys/tVugETPJvys+rKLhLL7zHKAkYYXfc/b7zcKXVOGDsqgVBpog8pM5/Dh
5+rgEt5sjshsQBcEBxnk9GEFfYYwXPlvQPVt5pYIIzT2bh7/MbLxZZw08ftwwF9frcqFZ1R3kPX4
NOZQjsctVvDzvi8Byk5N6V/yls+3SokNDat28NZe9YO9uMdfWEn+BHBENqGOm38orXkZtS0v2i9a
aTYRpESaR5giVpPVDNBLaHrJERLEqwtSR20aJwgoPOfEnKzFsCX5H9LNjQ9J215KBJncRlxx0uF5
uWVMmHpfATpzUpwn+0KgTfe1mqg44rVBAnScQYdhTxzl+omiiq8dtQ5NdtoYBQcIU3dKrKBT2bJF
EzOXD2T3XRIiFtJW2elWRmIvBSqlmix4bzv8H4jtwx5ZJvuemZQDpv32FwCTWx+p/h5bxYVhXr6K
nqxiClYry7xLZs+0aKU+b9yWvEbPIs7FR1LQpRGvdgAMSu6ojJYeXNVe3W3bdLRZYqVtAeXzvcHw
pCgv/RrGoouGJBJT0d3LrtIBuwcnLUkVc7me4ZPczBNzOa8mBncWkPlzIpHsccYGlAZr2BVBGDJ9
8uA5ImFcm9aPiggWNNF+UDwDJNxOTcRXP4UNLm8olKa0TRNwzQQTmaB9zHLfxyJN3/s9s3VaFZe3
qtbXXmDHyB5r348Atli0HmNfhZkPe5LmROPT4uKi3k0C03+d4hY9Q3yG+J5k5IBMgVxjIEk/sHIG
DJIFJe01ur1Ff3brBkvWBJ+1TDveoSJvnlllQzU0G4ar8PLWA8wNkyEdmC2XCepihhqjbpvN9yOn
V2ZbjPTZz5C5Y7idU8IBT+1H/270QOmBJz2i47Erx+JDCy9duMmtHra6JBkiyfWw3FT1T6hsJWQu
sVYuIc9Xk0EX4FSeUNlVbf921oZfCHDO3LebKuz+5Bw2Ec3Lz0Wjey5DJ9vkJD5FqCFLxkEwvDhz
/WHC8GCcgrbuENk8mCGm1rHzRKBmUfP060nqsa8bo2iQgwgWnHJnkzAYp1JC0w0Wj/9T6AN8pd+w
AhWOL/AA/1ADOc0xHyj4iREUmgJY9QU1RgJqp2spsfMA2BLiPZ9ZkaHbDEwBzME1ygi7LnNNjgaL
v+ksydnNbOAdTgOKneMSzL/bi7mPWNN0d2d3CbU5CRbot2ZGcPBCazWdgwb1Y7x9OzsXVfji//Ym
bmdhfunrC0E+uJf14JVdmasFsjPvltW0g+YuhINr+hI08we+9jft7i9KgaIZzhfIPipD0+5dBi7x
7fSuZbmzcyHymDEGhF498pVp6tGStTnHg9mpB1+16CJM8RZy0huy6M5T0taE4Pk3xq4H5x7tc1RG
qnXk0U0e5aY9RccmQMQpj07InOEXGKrFcP6JcZlUgRTgscKYXa7OOQ/sY5aFHzpCs62VqoLtoBzx
Wnhf/2YMwrQ0K7qgnuXJLVLJRdwBv2pyVMzQw3ZmX5RNq/80omxUZRVaiOG4WJV+n1FZ69yF449S
kl0Ng4jofNJgor7gF2e+mVzBy1+PyGTjqWjKkF1DDTHQc+pF2gpKbceCpzn2yXXiq/LDWs+K8L1P
Zv87J/l/XJRFETu1iSdVcoBuaLilU7GDzPknUTXFgEx/4auQqHJWryDOJTwju0v4gpczP/QAk+fD
14IladGqc/OlILi+7JMXnS2DYv1LHW35DCp6pKKd4bEoMPO8VccRBY9+ZrKkaPodEcfFLgeJblWD
1gyS6wJvLvuHBTtTwJsiSW4ykIXN/lkVMPO3co0kSc0xKVSEQx5E2qn9XadXfI17MZrRSDfPRahp
hyYX6uf4XOBmdpTchUGcYsZ/xdDqaaC8mOZeLJksHh4Gup8+ZMcIRA31d1Pi7+oFhmdAMHYPZuBA
GFP3pRSNS9OVSFjwRcEDFulM7uBz6IqBrFqDCQ8VyKB5r8/BvZCLb3Fi3IlxWzG2IhczFrPnjO12
TpDYWkqZug8bLbakM+2qrxusT9ERIa5qX/PAhMKGsDPaZ5MFAUHqlXMdDL5h4KkHzhf2qa+Kkyut
bAnaLRVm2iH4P4Oj8ybzWw5TvBooHYi308dVu+9qGHCWX9uLeyHkSzZaRkEEVDAJ0ISzdS3/6m0F
Ux2kFW7jHxzv+S30QALTghafDyhEAz5jV4UFd2c63jBlAttgd9/Fs65sJZlESNV+X5COHw11Vich
noUorJJQyoh9TkjS8FmU1SiogWlIQG/8JB8VkUHp7c4QRyvk2MHDkzahVO0iGOAWW1xyRFPdKDiQ
SHqWUiq+40wnDS4817Z/PiTmSNubCLEW0a1zffRyG+ajV/WaxEPagX02jMBtHR6VcFnPMRBLogG6
lDVpsofw8qSlMg12Asi0lPcbh+XHuneYtdKP+hveQ5Ws6tZX6any9oN+6jFGsK2z2x6HI1SeDSEO
BGxHsWsU18PdtSXEcQh9BSZEl9lqYcBZMxQvgimmIfbmVbT2mTwDJwTkX7zQuohDhXuXd5R/kNoF
nLPHBsZEIHCFQZm11e6F0zE10N2XcAauozCxVV9UMekWDeyjQlAF/7Du8nC6+kRA3dSHBQ5tMraR
j/VkVQOynGiLoORiuuVitW0DC5l51TJFHVC1FSOn4TtivBD6NOzSuoNhcTq3oOBNYZsw7Mci5n//
blzJsoCCnl0HaUTgsPzjFTYSg1JV29vbx0C5GDspkWk8LBB7j40WV4PwWk//s4/TeDjZhgTZ0Lvn
NT8sD2jfE7M7wCX//COHHmA1Z4Deilr35gwREw3AO6of4aZkI+hgrNjV4hOopWlEAQ7Irjx1+sG2
NPRIu+w0n2RgBcaDu3YnJ0Mb9FecahLglrFgXkAA9rkIdGKiAKBrlUXC/kZsEOOsPeEOTa/NFFe4
hyXo+rMyWEfI2KduDpGLG5d9sWvnlfvQGbsVpdmy0cdBj9cN7xbdfvGlnUQ3rBniZS15JCiCfGxt
61daEUAR8a6Hn9GWY3czwiUzv0/oGeqa3jfd3serRV8JdjpTdhxb6YPjwAA8LWTatdl1Zob3FJQP
wpLeoOekLXQs00vQimeAsL9So/d9CoGy99zSXDk6syLo7cHr1pvA1adQBk+w1TFe5pF2206lB/IR
p//eHfD7rvUgcftIvRJl03XtbZHOP6XD6uQ3q/IFPoIXDVL+RpUFb79vqmq8Ct716T+9oTb0d5qk
mpbVk6W00soCGapO+R+CevLOK4Bw3a5UsfP9ff49tnxHEiMpcEyp/n28Qf1NkoGO33FHbNOS/ywG
ae+yJSnfAbv3VVP6w1RsXSbjBJEm55VlOPWpaVUKPW2k2wkMH3PF53AG4O5a7Vhv50hASMxdanh/
OysRWwgVDdX33dhKUZv4r2NKO1K28RhWib5tXBzc28ER5YHy57JP80erU0lVNM7xZ0ziiN0qVrXm
r8wc0GccgmaI/srrdu4ymD3tP82LBHZix7v9OWNZwELdbsKP+/newDnYYV5FmxZ/0XdYX5P5L0yJ
Uh3Azv9FxkJO1JFQPRl1s5HPCbjQTFLVBW2v+cSDU+W9o7RT1r81ux56ePxB3FsFtWM13LRL268X
0pnBJPzsKHBGCDH4B6+PXcdWc4fOw5nINjVMzTwNZusYe3J/xHON+BziluPzO0RZj1RZgKd1oNIc
95Wp/deeNxcdJmZ57J6wLcaNzoMviEdT0nRyr2zzqglWRydqaYTZoc0J7VoRReQp0T9f0h6bgaLg
EZwvMVPOlZRvX+iSwR7W0y+qyX8n6kFNe3kh1UUbV50cqOTIxzls7eXbElOy9tK5xYKga4dvote/
gfWnBoFqj9L0tQQxx5uanYS9qS6IL5/yXtFC3q6V8j8zDq6Ue/ZD6XF7s6PeU8v9F+mKx2vm/zX5
QMmnEjWhaytW8KzmMaKz3KVKLxFp5qTxWDbPBeQXcUN6GdG0lHD7dyuyia4FM4M+bHsMkqgW4U0N
6eCc+yHLl3ZvRR+Gh8ae4cG0GJR1of6qkymrU7cSV3eRMsVQDnVnED4bBatGs6MBwhv3gHkyqdXg
OT8G9MU6PuoTLQCKYgQYGydRS0nZhqyQIWe8A3heti+sSkaX0p6xZTtmtIYPcy0hYqRFE8Q3FNA1
G8oAP1g5BVdw1ryPUVPNmNir0lGO6/UJt5drXT2lVgI9/UfoWSoTRz6NLES2IOfug/Y/BMtWyAI6
0nQzpn/n+uRupKYXZR57KZT1yQlykmezn8ZN36XpyiYyGmx9dRiqy2WnNl/McRsi5uj6DF+mTw3B
BrGtWyUAHIlqUHI5QgZN8AO8TF7Z4jUW0JM1Wo0XfVvSELZK82ameilMXpIU08b41ckyZb+Cdar7
9IxJFgSnysCU/EjwQ33douTFJ71VIfP2tAdFIv3kp+qkNb8440eDM82k14kekhUny2Xwxbh3sbuF
ulsdxYBOisdITX+uAyCtIR+ZIVAuLqpWhl4JFg9nsCcDQ52XDSYiDZyUFGTfoclnnzF/W0lBa2ck
9N+pZdlZtaXmHaXnuhA6m4yChArLbOg36WbGgfNIf2VRX5DTeIUOLbVkJSL10g6mCqM03nJfqR0A
vT8+m0v95hfgxIZlit9ewqjuSgViMKuC6D45/3fLYmLgiB9QV4PJOWMjKzeV5qAMAfY3eCpUIS/q
KdgAcp341TfwARuQq8+JPd3suORZjzf23DIZlEj9UYpsV+z0sTeqZ+x96lRmWomZaIpN1tdiIxsK
+I2luOQXL05RamMe+5cY4TAmff9W9OxlpyIzpCWwFRA6gipKzU91bJlZQdVT183hI/KVNKvW29S+
7OF8Lys4Gk4G7N24U0U0lfFvVUZ85ImqbaRy7Xu9chFuC0OeIOdlvVv+itCLu23fU/kMSb9WNmE5
zwPgErtHGPaH20oJXN8OIT7TYs7xRZvqec7VdLoas58VOP7frpx2QJ4oPmJlUjlWSjBdwf6uzitd
gEXXNrTnfXoA/7AaoBMAIBGG6unypg1GzIY/uGxgDSUHsaMxa4xk6kaDv8umW7hQwut7Z98PWSfB
koO0I0DjQFeQAkhsCA57hvhZ8ncVczf2Pb9TEUhQ5jCm41SFPnb5W8yUVIlYKhtpyhxxtCiYcpQd
f6ZUa/vSs3R23bPmnEF3tbhtYNCW7jTgSD0jEyRE5Udt2BCQL7Xrf0hvTyAQhSAHZQdjIV0vA0rV
ON3cluv5OfJ6Oyne8o7n9GiRik7934Y+EMWPFT0xDm2GTB7v8F4rJE+RkTt83S9VrhQNuZ1/SD7a
z76pdOeyHcFtlPo+PahA+cbvFyXpnQcBiJgrdr1GF83GWFTTQl3QBZBRVHTtb65G23Hcoe4V5Y3/
tC20QMnf/aaFE3yVakXJXp9tgXPf2iqkGzh+hjeqfuSykSHeRL4YCKgADwZXMQucgvJICryEMvkX
MVi67wfXW1RRcIn8xJcghSlwzjSNk4uiiYRmEqEYRQRKwoHwJ742zMbVSbh1JHd9sLWptkBnZ91y
ipOYjKCjekFAGTHccIVYmdpIzqiKw3ou19qLckte/4PYRbui8wyjx8V06SRObmZaIXv2feFqPj2M
xOCJDn9ZPJsny4C6QmJhFrgmw8ZghjNPqEgZtzpzeUbgKG63djcbsUHZe4j4d5J0msB5bIfDChl4
MfisMfkNZyo6XA9qQbSJ15TM1VYGgE6FmqXL8nG+jJrL176I0hs3XjpOBnAR8b105vFip91Whd16
pOq2FQYpk7v11sBe7+bu0s5Gdp+MCS0ZVJl082fhmm5+Q7fjWDGLrtf1l8pTG001Kt2QvVvKPmps
oZye+AbyQzEcSeV79iOHgiMxZ/IQOL+mm7Kk2KzmctrJJmAVChsTbvOT+F3YCMeYz6jqSjBYH8lk
TB554DW6UAxHK7vpMZ0FrmQ+mErl803H5zJTTbdmjwcakDYR6xxKSecfy8y+d+pcGnVi//kJ96t3
jfzpTmZW5e9qtZfc+t5xzGec5xW4LSz6Pp+MHeB81WmeR4V41oOTtHDgYEYdI5yL28aVKWncb5HN
+UBjz+8fSMjHW4yNHod1tIwXPRM53zocdkUNCwi7WWBEBNHMQClzZwliIx1xyBaY1Fhl9q1/EVlw
kRg+X5y4CFdTm4ArOZB1z5LOaxNIU1dEPiUR+VVfdce8AaEjuvu1xqO/9TblSHjXVonUeEb9XIwt
pCUNDlPmh/IIEUm8KWLufag7XskEMavVFHPltf9gMAVa/14XWRsUoB/kTRzCH2nfuOgLfPjZpSdn
p9cRgduhz3r+40CCSzh2eW8Xi3LE1hbARW0NnxkfjbKubD3/IuarU99JQqDwiMqGGc2nIsRY4JaG
Ny2M70a73WfJZED/ZXfZhbJo2YiP2hPLayWYiw7IaaxrXXE5+9sbkrrg854CQXYzHxyuUNBtQu9r
vpXnSHa/ho3OsZO9YDyDXtvUD+hzex8cfPDpGIFGPhV82sI1dNklVPttkMVnxICNXscKCFNjk/Ir
2mJcB+modWs1fNgP5PRLhW0QTlnaYp79fY0zArVT+dECAZWHb1D3p7VgTU+Jv9jOsqyHY801C1/T
sKHE6A+52F9/NyCdENPPF5sSrioLUw3hFep11mLYziQ5GquAllAqiPdLO7xEAy2cssI4FTW10nDZ
MyfjAmbOJfXfs0a2FSBGhgAUE22USK3M1gfdPoT57Ykoimnxz47SdRD3XwpJdl8QNHvFz/V4nE/b
4edeHnUyJ0UT1eU34mCvCkA55PhTTv8STeP6I3rO8uEBUKSv90wzvNYeqmBHP1mYBjf27nwBcr3V
z1LGNJsk4UzSQHk2O0bwPLTX/Nd0LpzzynEjbnYuyb7e2teFQ7xTr6E3h/63tfkzKGAcYqnPxQx7
8vc2SJmsHefTItFttQkIGFUGw1A6RyESqseC5mCQFjXFHHSqhIcjamh/w9jDILn8vvzLg6ydxlnq
KcPbjtqrsCVXBlx8Ui9diwWziKO1X7Sv650mTljgGId1kCYIFc05Tj27zs+DRlpA/XBbhyt2A6xZ
8egz5fpHeSwVA47MtdDoFninEtN76mV3Yyqu8mTf8beUrQ7HDuoFrUB7CRR4QGjx+DSwxHUy9mW/
RbEPQhGZpv2U1i+acJMFNyIfKNth626wpGJn42hcJUwg1SGSzEhLtSuWpEdHRYo+RGLUxmHO4wWK
oUqQMKEbQ6ReuUqy/35EscqLYXc007eL7xWz2+mLCwXBkWFMl2UDNM0ZwMLJe5EAoLf4J1796A6J
Mvhwb+1Tl6gqglESUCVDgqFAVMheC1o2Z11iWlAnBONwGI4zwiwcnjFYHkQtjo/TMSmK7WrtWErt
FsIlSZFTGjUwnRGKn//jur+bOJ4cCs3Rh+5pDBnme9lyWTdOyBDJRzd5WaSEP/6CeN+aO25K8Z2/
K6STuNpQVlEwLq/aGUz0HONHrN68zCK8bhsPlsRQWj9Y/Mt3TPlLAxnUSnWiXcNsNn7shKajwz3w
k9z2nyBK7LGmgVv+BjaV5dPuMh5uv/bR7QEERISNU/gDfpuHcoNOHTUKltAQTJ2EMBOnzRiYkvFp
2S/Hvg3xUKdkvEF3AmfITayBdRPQDJESBKXWB6UaxvlMYYuCNb79BNDEJunE7uD5NgswwTxE0eZf
vEV31IQrn9ybGcwFLX3ZWWp88913eacOBgYQBX7AbhIpvQqVaLllC58wCrajgwzdwiIQmEe9hWv1
ybWJ0wRssniLTsSh7+zvsSfX2uu+YH8sboqYUPTdVbvL1sx3FBdDFWwdOHVIfz2vtIE3aQ5d18Z1
Dkqgrq9vAGQerROtc84a2rJOF8QlePolHBjzOzCh8N6P7LLN0OlyLALtoKKmC3n2WP6Wl1uCLn0F
6sADQVd7u+oc/34ZSUkPLrcuJoTyr/vGWfcIadwWRo/sCiH0id+PIEDuOIDyRokWux9g/ppAQqhD
f1Qyd/dKo3Ap0UvSm2H7mte8JThNVkexeHV+MAoj+BG8MopjYbxwHbzuBqie8K9uAaPHffUAnIMx
ZDs1vsniZd62E+6z9mzS0a6ELDDpJ3peuTy6zHPKAVvt8s5SrOMaDYfp4KHuRXxDAAC49G7iagLH
oLUJyCq/wp76SrL8DAAkgayFkc08yZlCv/OoG1OJKT9mwRL4tXuaekucJ3zNWg7hKla7ykQo2S0Y
ldiowMSLK+dzoLM9yDNR0j8kU27NP8JEIfGotRUfcwDrt6qpH/fFm9umItR0/WRBe5pmZnBZWfPc
ab9JRUKKRL/sRIVEYu2mR9RDgyOZFXlN8HH/czulnGH3jVd4CL7t8rXLV+2XWtAzV0JDNFisPTS5
1fr9WbQzWS1tHHXVcUrGpcJnNVfm7BirYavHezHJHePiuYx+QgOfgjSl7yI2acEq+HLUCvBgiYsM
UktgiVM7YiZDupRmFA/1YbraU8syTQLGQCJ5i5ivu11Vguv3qeSupSIrN8hgGGFWA834lQ0ZUNWt
Ul0AifyyQg9iT2jUMxBHO3HBF2JTOnllqjl1M0dyCONeeB8fdfclYiN91AseajX8qszT8Q8XKyDR
qBaZddnQp2Pm8/V0zis/k3W3oC52JmphmoXuLGzlBq71FC74piNHTXm2AXiJUDHuVFej2ZWBaVZP
+IrtpndvFlMa+Ka3vXpLIcH2+E5GXxiuWkjdcnxEzCJnOJRKeq8XcaICiuB0MU3tHgjbRddgjLXV
n38TXFV2yNzHSCC1rVFvRLBjYvUCL8HaqupstrysM+7NOsBAV0ivv/+mt4ntR0BOwFaSiQyXRtzO
PIgiq8P1t2ZHCzrgoO7OplT4ywi7hjg9w91Gnfd6MkzIUkhoUrmaYReAvZC37QBWFsmklsNPnnnG
LDh89Cx+9Sks2I1qmUD2ZeK3odieXT7xGYZcHQ0WYGS2oU1Ej3BHqj6vzdb3ARFpff7pV8QBf3DK
jPRRcVp0WhnrU62+e75iVYVZn7AaEjImnW7coJTOD9iXzkZxKIuyD+uTW7qF3QnlCEq/bdlqyFxO
r81KKXrUxCqLcMCPeUiMx+U1hozb9SeqHyYqcobgauCKEN0Rz/KMtUZL6swB7r2yqN2aGwa+9wUT
egMKpWL237w+O5o+SiuqikTSOXjAWuiODJVRr5r7IJs4oOOV6W1f1IozH3jpv6Uq0wTkDec+68Aj
YlPHN3Psh0JhgcXQ32zs01PHCXO0xdEUuZkuKy2fleHxAAUkGb/aY/K91IrR35NmWEB7BG4rVk1D
FYedp3XJdJAk5Jx2+YDAltwASrvceI/XLIpN+kuOl5u/pIfmk7EEhqIdJBlXYUJ08eO0mPdxWP3v
ZJzSce/Tewpg1DORqkshoZeq7oGUIs06CJSWG5iB66H6xoXIYVXKp+oY/NG+PfWf3v6MEPd+pMa2
QyU9r0ErL9lVkCh2PPNwNP2DFhkbhfBiLV2B3lxTbC9BSy7WKNQZZuIn6C9qRqYMBVnYcf8V6Mv6
5DEV/Pb2J+c2ywKQOBkRT5lK8vb8HnlOpBQZk5/bqjNfvcuhVebxg+IIKa0YL63UZeS4XRV+BGnO
DPHNz0giLwhqqttmGRdiZcE2Q8z1nNwia1AMuqy7UfiYAVNKVL3513O8mEBQuhHUUEVcnecC7IJp
85wYNn0JBs9JnqLQgq7DrBDPNAmdjdbmZJezK+LESXug84+2oB7Igiq5q7n1IU5C1jqNrZjpaTh4
7C6w75cEsnGADmmtlveVqILxD2tB7aNr9IZpSrj486ajMqqDwC7ylM4f+9bXRdwCzlQcM4R+SjMB
EN3M3lmCc45CBgA011+fhtQFh6XJGDsDss8yYfzpJzisVYkcs4arrghXkioNkRip9sOIAB4OEkzC
a/t/r1lPHL7Otb50iFhoM8p5RVh+KVxXBFO2hnXDHWC5j6XRSeHIr+96ta9wJo+u1phhea6JgYD2
9s2aqc5ia8hFhkLlwpzBXaCMV47TrIt64TEJL1GJ9h9G8A+T6mOfdAWI90oiP0ErpFce2omRyrVN
O+7R/ooStyJJkgKi0017a+k96Cx10GVDlvK10KeUYG2GzXdjYwNFEbMUBRfFWuXxGjIDKIFCeN/v
FV8x3GqyBb7IrdcPGhON+N/HsLb8R79VNflqb/R59oHmBXZYOc35EgEOERezri6sPyCQy6PDIEfx
z/PPXD85GkHnEwGf7NQL+T679BOi+fQdqr5yWwVltiF5RHN2m5t5Q3DwmKJwJE4FEHlbu7gxCu3S
r34SMBqNACiqLNzDW3YVIordmlb1fHx3enAhoa7/m07ooCx1Xu+jD9SiMNcei+kubY1A03TKKt7a
Np/+TIsmQwTUl2jBzktVSWJTZjYCBTuEBIOkymcPOiUus3KBoEx0lRDiIa0Fybc3WdZHkgvthJA9
WmPrKBN3M840MV37co2HVdOvAb4VZ14B+yLwDYQAHlhfHzlGgrHpCAiVLQZxXd20y8LtuFRy6l9Z
nkmh4ZJcJaQxZNMTfi2TH68rtelrZwHkS9MGaH8+hNF+iHokKOAhIIKgGpshHn3tuGAbg0u860P5
n1s8Id57tMkQhBG/PGlM3uw2MOeOdIumP7vd/JUeNFhvnQkB64gAf5/kHFs9G3yXlkS+xKi5dSjK
NjG7jUBGW6Qo5ARgFuNyTic+1RvEDrst18raDqd2N1qy1njH4A4UdeGd7qFB7DXhhw/csWKok6iY
Shbaqheq0A8uD7TzX/A+bEHJXaRcUbhNT05YrBpEZWk3X3IxFEcwgbUaBR2MC/VC0Oh/PV3XCrMA
ebSWVCyi8U3i721Ph5Nlaq9CeOQSY+jZoONBJaO9DC1D+CZDPyBJ7zJ3HeG7T9Jajg4MqXAmyFy/
wzJt9QHhM3LtvsQ583MvPFGGANHKeL1whBo1QDIesCbN/zr6iZtUvbeUB/Ei5xuLRa2uJ0F8k/RQ
a7aMcbxG3SDTNmG+Xlr5OKJTKImgjT+seR3Rm1gWODTzgyEfWyxFwbWlePafL1fYqrvaSF8dk6hh
72WKgn0ljs9gMADuaKvguuwzeY3KFocm0lzAPYbyvHRRIOrSI9kVGWLkPiAUg4gzCAW89bHd5/ig
T1duYZZlXC9CnmjnW3UyxaBQoH37m+Oc8RLyppdBw92nN5Gpgr5JqqWG2MEmg47CdgRZr85zeiQw
eAz4oUzsWL1OnN8sqQERhP9HHAe1/9qUNHe1Y0KGBPauOyIGyCDQt67an45XJUlCmjVWZS0yoCBj
AlZBz8lXZjQpR02BmFdbG40c2mJ69SFeC3LT8CI4+805r65lNavE4vjN5XhEGMhVY9sVXQigSkPY
AAW0nAkgpQ1M7nembJwYOAEuCkIaJBhJlp0MnsQ6kLHLjcx8eOJc1H0koU4N+dpmXd0vIxYirvBk
joZxRKAOW3s5s+0svjL6eSZ45oWsvxAxIXGDbHDCzaWN9xQ10laZdpnH40jwcgrCRocMCoF5ehOC
KJxZF0h0vcnkQwv91G0Bm93bLT6Zr2NYK3No8qO2RqG14cMK91GpLHvCq2EOaj4NqYWItTnPsItI
/OfllStaxrEoNTkGwfk5tniG8xiO5QUT3MY78qI55UDwFKAnBF8mO/B4/iF6BDCOSv5qeIYl3A0e
faqn8SRuzl2wqQB50sicA6t6acUflp00cE2h4ixALgaKr9/LNyU3gkah56LU1cfXndSVY4QgYvJO
c8WCpCdShDzJBeu6CjjIODsiu3D3ohaag5iF1q6v1qzEJgXiBCB2RTlOhl5AjI0hlY9P7Gro442T
+5r1RZMCl5PEbMF1CK0VkLt23x4A5SuOZOAg/iU53GW7Z/uie4SUtiXMKr/pJJ2Zjpbsx9sPFmXV
+VCmEgEKqxYVN08CFAfxM8CfktSZh9NBg7fFDzXTI/bRejpT4RVPwBVSIczGNZNoaQkLyD3zrFbg
o2rm2vehYkarK0Wk6TP3ulJ9l4se/zW/JegcaRiXBM/2K8mnS77FHOkWnc+jqMq02pFIazdXCdYg
FZRnhIh+j/5iZ2TQA7uIPmsQTGasMb8CDaYTpNQomiS9bRDhzUeCVoshEuVODHs+VI8kfXEadkod
rp5uEMRGULh2ZYSzSLUDQWcp1HX0YDm/qAi/+EorgWxQxMmafSgcbAGk3ltNJtuZzU45tGsOhX0e
c00FF2fpqpPUlkjCaf8aBsw1DEBM0SLuJncLaODvnzHBtN3f7FYDSANJtaATaJFpCYKpS+cBGgJb
TRPDrsTGSkVFDkDBlrhTaXFpftaMLPJCFgYrRX2db+ohzF3tKkLJVschjy7sFuEPb3crnfIqyo+o
WTnS0YO3Qo8nBKS+9ikRj/LA5zc24BuQuRU0waz9NoJ2PNZm2tWhg+GWR0iZSR8PUlqvVnEd7KyL
GOQJ77bRi1ctluNAfeIXYTmZgjsrGt4JzB3y1+HElT+naFDBRpK4rPVx4KGasxlg7X0lHz6+cjhA
HwVTFlSKYVD7eSKnb36nuFaGad+0cZgCtbZDbY9TVkCEnT97/eVNYIYF+8XDJTHrXLs+3oyBus+X
kupGgxI+0O6KB9DAqjf8yO33Q8EpHbVF/70EfwLGnCyaV00hKUwhbYPCm6wBDkTq4H/aeLwT7rXU
Nuh9NBf/BsB5uR9/hQ08o+omT7hrKoOvK2+VbECJ/Gn8IBvOymDdJHUmfFs/LZ6CvLfW6KohGOLh
SqMK1Xzbi7iqDFOH7HpYoy11TXgx16Y30sMYP468S9kjTS73OiCgfu1Bv83PSOKF9Zym7RuT8U6U
M9SorEtfZ1k51XYprODltSYMmaLHb11Nip03Mc1L1iFz3RvfMt+wOCZwFKdU5zez7qdxfH+fA8Ke
EHVppEGzM3NYYZJWbwkHUPuTnPatW0shS2jqgGz7GBtMXG5ApDjdHrnYwtF0lFUGWQtQxQMvwiYn
EEcZdBzLU+cLw9DgESKl2nR3wMK0NL5CbnLhPcyVwmErbQdSXZAJxnTsiFHZe//o5MjBcGMeanPO
TyKXuAb5R4ygbPnM3AuiuEw3XAJ96+Yp3JZYcUqFCnk5BOhuPY++N0qwhM9BCM/cdWz7qqafvtb8
MwYK3Vdc0+x0+Cq7hqAjmIuNzkcnPDG48SgIPiU9Li4pXKXkWKHsZ+G9J0DIrgtgVxiLUaW2BLlS
gnimN8zUTJH2CZhPhtZxtEbZu1wNIq6nZBVb30HjoaW1sog0CjlUyKtWpqSVEN+DbaIuLwrzZmLM
ZJM0Bt6XbEMZ+0NagJPgfpGshUxn2aS9ug90XhlsW8ekMdhB0ZO8gIP8Fh4MuAaocvSTH6WI/rKW
gA8uliAAtFXHb4kkyP9anStWQs3V/OW9W+ATAcP4VkxH4fZet71+qWnDRrjCxbGN15PRkt33O5Ru
lzrlD/nU64WLfKpjFCTF+6w70apUd6QHW7IC9w5oTg5dFvjuY85AT0nESt1VbwML9gGpPt+uCYs4
H6utFxh5aUY6lTyJH/EO+CCQUGlDDTVomDHTFGerPRjT8ohXvTgf5Axovq9Xgw8wWzLINZIqUeHD
Monaud8TeQWcHGczg3/IIFjplybLY0z083tc68gNpIJGKxuU/yrT+Eyd3MchfX99mSKGYpxf6OID
PnPY5DiThv/VVkwJXD/j5swhAFUkDZwrmOjfx4WmeAD5Ajckc9jmOXCLvZAsI9f/oR/2DwX+7O5T
BXVvi1K1rsnTaLnwyjsEQkMveMOP8yDXPlW5NpCJNjdtIXEGdUaRAIAPwH2eTCIfvpvDCSjX+ydX
dE29kWtE4X5s8L4/0ljeF4UwcAuHD9NvW2Q+TBWTu3xKvX5EVbO/0yhMKurebinx9GqhnzRtQaKV
TLsnLcpPLTBrmOFqVnOdC6sGE/RC607CfNVCPFu6PyWtB8HdKNv2L7UmDAY8jFxxCJcgv1kaydPk
YM8AwC42uqfpBYwxDv7dQMfyahySUjAZvKkXL2kfVEqfhxo13h7RqgSKGkJ4+oGeBXU+IZWiieDv
sW7ClWRoXao57Z8BqLNEGhRCpPUOrCGQQszyqInWVLpTHI17WTQl1E6IkKBNHNeQlpDbVAnflIXv
L7UL5mzxPR8Zz/D0/jMiU9SnBbvb1Jkg1+9Z24GZPCSCmGMdqqCBF1uj0Zx/FBeO/EvHimSJpdw+
SRwGtaMM+3GjPUF/Q3ptW5PEuQWtJnwfxD2UrOwTXalh0F5xXrwny7rrbe6xwOpXWzVhkGs3R7Tz
9zY1hBJesDcTUWCQDiUzH21l1TVNtlMTYiKYrWHCkD+QJ+Bg451EFQ2WMU2FHEQ75KZT+uicqf5f
g0gptDDMTLRh9zIEbDv3fJmp40AmUE/X5meg4e+EZwvhqhLtm+LzHvaBhmQ3aJnnK+EZWVBCy6sT
mSUa8MD3vhDKtpAQRe8yPdb6nHXoNWdiZnulkKP+aYsLy3tIaT0bX0jviPZW6HDR8K54Cl4dFaK5
i3cYI5bl1LwbNPIVVR7DbvSUv0VCyYLiWZRszEhTOyBGuIdn9+jLE8v/RButsxWGRB5qHDi5qIHN
S69PVn8w5qx5o6q4qFdJHLyK6ZKy9/SKS0nWKwPBsh8i99KvBQyEYRx1SJrx2dC+pT83qFyBqrq5
4KPcg7WTTqp8kndGbisa/cWeGtI6LzXUiHz1Kdn+OizstPufdWjJ5J7ov5wFIbpN1Rhm9b2oiQdw
6RdZcUMs6r6dImSR8iTWqgM1Qu1ymWC4yzPj1WjzhLiHiEpc2WLMXiT8VugM4Xs2E/YwAdtPmJ0T
b0TslC8g+JtIUSRy6hRydvATGkOqel3tR4NJ8SiCiSsQU3E5WnRbnj1VxVrS+veg0Jvtg1BHKS+p
y+CzNH0Rf4UUTf+GKyAZhp0vAeujWw7aFjVJDG2xHmj+p9RYboZIq0zsG8+UletdVKQfAhXRc1aa
Aq8o1LqIfXENPVqDCFENbUTc7ZjYyz87PIQzfJBG3N5t+o0pV/hK6FSLZZRVLO3Uh3KyHtM+Y8zy
zmxl2FV+S/BgpGiCaIXKkNwuQcvJwT9RHc6CevjX+EecvNKKc6nXvYtQ2U0bimX3YPeBflkI5kD2
JQOIeR/bgJcYY51a8e79VqNPxWoP4cB02va7tiCiR7OUbYIZ1zEW+fyz2TpiI+BNPtpV4BeI3rM1
pSprpCAWSTEjhCeYxl38CIOUECKWlBNt2lWwItPVQCm/8I9DxpWc8Hp6aUXfl4Ru9Pfr64iHCKxt
IVp0Qbldg68rTdF9HsUyMGk63qt3E7AUqP2LkK8FYhJ+RfUMMuCNuO3s5cjz3DouC9FeyVSAVTK0
ycHgux4mpqxLsVox2u2py1Z9pPk/BH/YMFtKTdjJdiAxB1k0+Muao18hz8OwtB0GLesMy53+yOQJ
iZjmFgyNv6Fqs2Xm5rYBx5aLZH9+W7g6DUsS+Wslmbq55sF1paV1VK3u8bnSytBAwJR0F/eOHDAd
UcDvyv1LtAdoL8uUpvuQfdwbvg68OzDRO6zxEzYIwtolAB57Iagkpo3PdLoBKHNPMMf0bEKkwb13
+W12rHGv24N5AKn4Jwz77SffY5QDwSETeoKNMyNlJjRP2KnU7C72a6nnbD7wJsym/19H2K0Xf/MP
YGwTmkGghEIdjRN9kHRdasaqarW3KgjZqr3q8P1zAt4nGn2Y8KetaVlelP42JaU11jGbwBYIAH51
hz2552W/Thsoj4gLoViHEtHesDqBBXfygOajgQEO3dnnOqGgHvnMXvgcg4eboK1XWkeLvGj4Cp3+
0xM220otz63HMJ7pzJKlYDkTDZIIPhbXeva+Ns1HI0sGUzucUJ4lhOMek2vMG1+ZB5rV9sRN4FkW
PU+QPwBA0jhBYc5eNF3QpNHcc27HEHSIi9Jn6QFVQHcC1A2TkzYO4v45/buFlpY1YxG6oDW1ArFm
fWp77PxHgO7JKdR6LUQT8TkG9v9dPAzVstvS4gLvXu6xR1jr3lPZVwnmt12MGsFU0Re1JBSJRnn5
vEMY3UvoJG7fyAePC8Pj8i6IYdn67mvucg15riZcKrPqvwRklFyFABgWTvr7F12V7gDnLoOtGzxC
Q3PvkMnsrXbcnmwd5lGwA9dyml1eRUMC5D0XgtEsIOIHq4SglPmLoYsMUIqTifPvZIiu3QMY0A77
K+VYK0cAy7ADaSo0oX48vIJl2iMnfz9up3VuL0UvHsRT+KWnlR44tMOD/PSk9cTcJ1nB/xjLv5gy
6t5LtbSkvUDNy3F8gMlvTqGNBqtqbiK2OAFGl8J81JS0JywTrsfyQqSzmASkGJELGIlVi53Bj+B7
JqwRokkBZ+hKCpwdhoH74PXzpWjQ1qsS0WKYYyfe4W0tf3GQtHu6j7I0suvq23Yj/ca1AG7tPRR6
sZvwIZZVCt3XwJLOsblnn/twTZ2vF6uTqqOtQsxOF0NaKrjySrNu1XbSKI/4mXScnrgrcOdzlNyv
d442nYxzILkcD+KEtnnaGNLucECYblaOq1DgAaquP3OCHOVxwaF1R7FDfMmNr3DmGykYe+rlufDy
AyckwpDJWF31p2Ji5+JZOynFHcTu0fp0N8QQE14XCehEupMMQ0pIwm4o2tnhKN0eSvYl/6H89rHd
/uUiWKZJHKUDfUvgRdu4HYQEVgg05GE3r/TexYk8CTgNZFgdyxREx8w2sNpYKlramwvbin2sV6Kx
izuD9Gq4b3u1lq0Bcf7ekHq1aM4Euo/m+1Aiew6ykv3zjOjJ3ZWW1nyR6E7+3QOCMnxsm8tDBm7u
3f+B9apwmS6xYRhwEx6RQKcMmPYdpZ6CVyq8B+b5Iatil6SXzFT9GrXrNf/dYxG5k8SsQCjgL6yh
1QxynU+LfNAm67MAOqV1ngwu+qbOTiRN4mRTHQ/WzHQGf1zbB1t/C8DYo52CTP7BaFni0Rdlw2tI
oL2/eqSHWDwp0Q/GaLDgUVkiMkQZcVMBJFMPvFgtRM39FhK6aL1oHnKG4F1rPcNL/B9A6UdsnL28
nXNFCEAg7PrmH1VKSSCuh7pznxV3m7cyDS5pnV+x3ZfsyLlAN5yKBM5Cn4Jlo5Fo21WOpB4O/LfB
YnIXUE6m76zmr2TX8xcP8PHuXLunU+5WsZk8BHcDJsetkHp4Pt7vi9BEa5lmA7KUE09wzkpZ5m3a
h6009XA7uWbgMM8K5nDXbbUTbdgV18Hj2yasBAQ8Po3yktjC/eTqE1/ysZtMpQ6tEidX1sS9f4Zr
FI//l+nUufWbH03/nQ8bmpFp9ymzG52K7fCAtKbuu2bxEsBVBOdvz7dr7jJpaCatmiVv1L8I8p72
IyriffeHfFS7FOAnvU8HG//LB2Cc6lnMT8om+H/ltHeSjN7Z7wekwGtlmZYZZZ7nxpQ0W6n5PkQS
EmcSLqpoT6FxsvIMwSmHJ56yf4PUDqLSBWl+ebUwMwRms1/JxTXLTvZucCx3lAGqpRl3HXFSqCWa
musHs/h1EMgi6YWKCYqkIwCDO8TWZ0arjOYq+QytUzC1PzU9vwyY6OI+FDO8aiv5mRkhqliemtMC
lqmTpTQlWDUgLFO0wFN5uxPr5V+ubZAiyYcE6wrI06IGyk67butNABwPU5LLYxOe3vRCLzyfHSRy
iIufkHqT/BlucvrHHBulJgbjX6Z8I/Ps/tFwHT2xY0JeIKZCYBmFICF2E/GjkgaCWNh15rxk1lNR
Xql7tIOZBv0u4ZrlzAxjjHtBWsNDYrujbI1C4ftgqc6z3d3Q6xh2P98O6KW/QPNiilrl7OxRTlQ0
1M9/Gt/63BCfQ9TafyOKpL5chBrQu/rbkFjp+p7jLypk9P20RS3l+25HYm4TOFUlxJtfn0rzPINh
g0QGzANazK5LsVnYpTHNGIP9zZgkEIqPuJ8V3/3PMrB/jUYMIQJ/q1kCRR53FQlgZQRW+s/qmIX0
n2wMEcx45rorzUWvvj5V9HSLXTaYyqQLukg//ZAuVW3fq6GeJ/VJhnpX4mq3EY+S0bK0sLJLCovg
Sy9+sfFlyQyRq1l+gRlGSiB5DZQ7uQnf0JVWISQnjomyAvX4MHd0ksrlgX6utAtdx/+rl+7QXQdK
EwYbYCSFaXOpoMwUhjhND0IXHGIuXqRoeWWyrEk5JY/h/0J1rrfrMOtqf96E76QsGQTeEN5c1ucV
W4xj+L76s4lKgPdQ1HSdHi9EOYJjDDSoJe16dXo2+wW5ntdZAbjgxrF+hB2vUjV48Lg1EdmCI8Sz
KInMhAH7VHUK2P0Xi9FelcFPinhvMbXqDVh6ETi6axP6VbcHJcXv/BtO7YcjuWY+pScKVx1IiWeQ
v2+cf5trLOXmgGbm6xxQdxklZlHzdVHq/DZl2puE59upbU3piVSG+0TZt8l1zt3h+4l1tOnOMnWa
0yHhjunUp/t4abzsK+rjmGYfYTcJvsSD5HpeR92UPwc9TPGXcvXfUlGIIncgNZ5AuolEQ4xOrZ1t
nY/rXQBiUC84x6qRxeHd1x2eZy/DILTDSBK6OamocJV1LHQ+XcdAOP3dffi+6jFGtFhUdBYw7gtg
aXxb8HdnXNFnK7zAeOpYl3GFbghH5tfHbNyNHldbG/pcKgi8lsoLMK8n9vLKoYWpvtAwj/YeNOgW
/vEGCurY9QCf6ut61fu0DSaHBDLn77ekho66tk0zB9uRW8tyD+tA6DhfiHwygA7xIz06X8tqtVVU
QvK3OBdk3lCGDKSRyO+o8QceMJfmrTLLujS/ZO6L6PwmNsyJRLqP04+TVI+cww0tY4tXMLgwZiso
gJ7Tb6VzgFaQvTPJNDRAjtyZL4WfKl5QfNSbyKCGuTZHjtR5G9t++lPfDZzhDlyZXjLw/9UEdTn+
1JjnAAch1BVFZ+8L6bh3+9th20o8XF6X/RtEVSaZIYv31ZtfxDoAgtosfn5i0Q6OJ4Ia6azkqzpO
xbyF8+GUFAw61TT9/CXuiY9dECNePJhl2fEbybi8es15NT2BdazzRklo+680hIXUUxyZc1d86Cv3
f1KJ+xoCwn2tmpaOGHcsq3jcttR8ka1j2pR8JKcwmh/R/SSNAQwHEkUX3XGCUdShMSpiQhhXuBzO
xS22fzskimaGo/XfZyMg0OREoXEkAgZyjwZk/ulMXeDNOHA9zivyzflB322MG5QBUP1RA1at4cjq
xIlFlqFaxRAOdjjZhNAEmPqOBLXX8t0ZnjJhVmOmYHXEUXoFF5YoofouXDAO521XfTHkwUAEhzKg
o21RnZllaEb4dtRRW9Zs6jdmyB1PVeIf6MyfqpYLxmJsvw++WOPEv6+RyVtRuJjGENL8dSdc8Xa5
gDrNHj//EIj9Nyg+dldPpA5YJIH/QQ6PcYOIwRd9plKNATFSByM3ehpa0DuLdVaAvFa8sLsMz3ja
e9SIFPxZXdtj449KLo+pSNro35G7nIhxeaPwQbOysHRswiB+OOVVdgUP3GBM7cPYA5s6Gq11DLNQ
GNao3Jn01ZHYmr0bRb52c2kBuRO/rSgw0oPJAVEQNWWu+uDo2K5dXxVi6/m78Yk6hdfGGfTV0/L3
dHuCKIo0kxp5uDC8LNOipdDNQF2R8GsfhY3hvxhQUIMbABxYwBbofnBaPCVj/hDy81y6/9f7BwSL
/9PE5F8rWsR2PkjT9uoSrXzPAJZkTzyPo2F3AnmLtO9AQpNlmipvoDMlzVji6j7wL3I0FUgRDZYH
LTVQ1o8ly8G2a7pK8tWYypJDcNfqQb2ed6JTqdtmcZxHoeOAEJccqNID2rpZ/ltOa7fe5GfBGr8+
RgQsKMp80os6OQCsXK1C4ovMhAqvW9eJKHGqLgItlJXgxgTsiABd1KQG6CCqfCkmThVJVjyeDkXS
y3epDaetC3NSjVajDZ3WFGf5gNSdII4t29nyxeX1zxlJMBXTQklxz5g72seqkW105v1x+gF/2+K/
Y4K/+1RQ23FjqZLb32FlsvzvS9Mi7KIXsJFqoXwZj4z7uv/MktgeB9sF3J6OCjjjBZO5qkHyJgTD
PkTl805V63m8/5VsGl5hJgKta2BQC5pgXA6X8sEdH4PUkk87o+uKkwNkMQm7EO+pogX5i6JKRZBt
JRwMiAsbaYLNAP3gBWvyjy5PYTIM7AZTL4/v8Gc2XIzI33ELf9XRMMF7WmoFld3LfQKI/gyj4+mH
9EAZ8tNJawBH7kbs1DLeeHJNwUnRHHwrtzLzAc3bGZm8IUNGhqJoeDldBUkyGhsYb4lo52dcW71Q
ED+r7R1zQatEGLR6UZiSoUNKn1ks8QtuEMNJUzj7bk3lb6H9XSpNEq1/wUpR1F/s5i9RRqno2zkk
nhONPGsnYY4lfX+zDQkU1td5qpbdqejw0Ndmug/E0eiz1tOohBoVSeWNvDXkYHGI49Jibetb8ETu
cLQKRBo0wBhSNs9Qx5Wxman0UjvNu/oDwsiF9/g0khI7FcjymrRMwigETORBKQMk9gNFCyczlBOD
v9/bsIZ2P2V3su4uaUG0n+b6cateBPGOE+UyTA7DqcasF6+c8MUtKljkA9BwuLlPHerpQhiosHjF
59Q5em+O0dVokPRVaTAZK/ml2aL+3kutUELKYomeS3vDfjIF6ZLQZ4S5dPOQpXxYzUcEg2jDeqYb
sfseeGTe71wgmkLo5xLsBAqw24FfNKSz0dFjBn/lES9nypaj5B+fwlfwoIRIRi3U91Th9Rk2M2Yt
oyqAsDUk39wYz8BZHcxfG1YecX9Nw+2sMriNzsUj2dK5QIwTwh8uk+cxaQd7DYuFWXTpHbxRiiQs
pDA0bg/6qV60W5ZRKs5SenZS7MxjQluIbmVzYDwuogN8jPDcKA3Ah/rHnhKZ23/UJtDi4tW3k5BB
akmowIvz3++gYoxl6hMqc1tcau/InGUOyOUMwa/nPKdp+LZy41Ek9sOKFj01mHcD3BLh4SNAomVm
fdz5s7MK0bIhTjmvlNGKg3V6azE6ASspyukggZnCHf73h+AySvOp5kImL4VDciIq5IgYBARY8W7r
m7fFa9NeH/3G8jJT2j1kRHd5VphgNbYyDwG9wcYHfxQHL8ab2in1GS7Rt0CJxOUmJPrrQ3lIg+p3
O6LzTkOCmDlIEak5gTwkjqr+/11tedSj2SNdApw2puG7HCUdSl0DmMTC4Yr4JSyS1QcKR11/BlQp
gpE4xB+4tmYLZlm6zDFeKZD165+G7Js3zritweXu6CFbe+AahnkNJPZ8yUvx8eNZtpEcC+kCmQXK
NuxdmZorMwUxHrvwu5b99CLPJNXzyJncdNlshY88PSuOql/FILT+YAqpmCUDEdNbE6ROLQwI9dGU
bKuRGPGlSws7gTB6moVpp4XbVIJq26GdHLP9tbqO9D/r1rc4AbgtkRKlRfoNlcGMIWius3q6aO5r
vT1gvMFDerIA/L7MdeDjXGdfHaNAC3MKvx8cruOj6ogq9bG0Kbr0OU3AHllsO3lZqOj4TFkzQSgy
AD8uSDPEA2dFbIOn1/81KWZVYC5xjVx+4rKVHjaum2uHXOfwah31t+HnMwMAa314N25FrWxZbRot
ib3vp7qvPNyxJ7CMRVUNRwOAXA6UU+Ur7OCOle+yM+WkyjuUHRKjIRPr52UacFaZ5EBCkKxJZW9q
3nRrilpSnOeX8bdvDdeU92M+h26l/tqMPKSspMrhFbzQDVDQYvq7wfWorZnsTr3P5r9xI7sDMSwa
6n/OGyeZgRJyYmIEl5XPnbZIBViwxtxBp6oxglnSaA8f1uDiW/rmmKhVWVJ4guNljxPYzitrZafZ
o3qYhg+aUH3moNcn1Zu4DPeVuJHDHwfI+ctWfWq1wK9hRsz22fNzmp61PigjHitUUe0FldH0Qz3B
FNgeGGvllnoQUTMHBnH0WD4KcD61xd3nrSYggf/XYMLeCSPP7GsfQGDN5jiUiaQBomfpCuPv2CXX
ktrQQC4NSqNGPtJ0L/KOZTnnw5QaCmzPluhST8GgZjsKEXK9VY1gKDTMp4iyzH4PAe3ZuL+kFTtV
SNPCFRsTeaz+j5TTv9rsUlyRZns2HH6+TCCIVGcH3F6lRWK8/t/JMpXxTXiKPrMyHH+ycTT8sbzJ
xmk0Wfld4LEiFNV6Rt1rGe1cgfib71TMD7JDRa5YKBfhRBakwruu7bQuUuy6oyUyNUADu+ZQHVxQ
FZAFQBz46rHhpdfcELtxS3WZ4l+qkwwEsjy593dqzwng/Dv4Jdp6f0/R+NdDCzuRPhjtT/Q1Yz3X
yKX9hsiyPFDsl2eCtdyk9Lu0hSVYZ3iFPwQnaivq1mcOqmhUHD/L7505NV0LFOcWc++iZEOdB1Mj
QHzU6JgZTBdjPIQdQTl5mhDOJPWo9cxW2+u43jvER5ieZ2FJz4cRYiozhUoTe7nnV+Op3VVDy+su
WII3YYrVIvBruymYoxTn4FS9QL29RNEtcqTEghznnMa7ueeSu0y0KQdypd8TZOHU0oOBvkTQk46m
apDdUo7rXBaNSTUy6gTfOGr7SDGYPXCy9JprtJewR8ZrYPL/+N0aGTDiotMLfHG1EKba2rSfLK1a
MzCO8M/e/sxzHHE4bHm0G0nLU+viz4Skv/wmqCY8iaerGEGNmfq9BRY6X5bKUAwFqWi82JxYgA8g
fYBhbXuGuELwUu6mJ/ITDdFqvW1GSOx5fJrST7gL5mOEQSW0nT5x5Td6e4IaRoKPwJLab1oouvtK
O6CB+r9XOQ7hrDXoNkGcTqlnvhyaz5CgXdMR0MczQLkV22VuAdDSVKIELzU517A1CtppdLk8uvzZ
8uVri7RmyGX77JSAhQoox91t5toVJ3YHoWSFBMNW2l6bc8AKt+XWvxuFFdZlMT4dxiqtVNA0mhje
WspKIGHrAyq2mD9ZPT63GfMdQAm2s+xHrsOp6YYwReAJmNXHr+/55yzMrIa6e8ULS15ZFiU4thOg
Y3F9Zsd4gOcfQscdZYdSOZ+knJHeMHMy6zQPoU9F2j37Rm8Lf+RQ9FEarn7kgo+i5W/g1S75oaWV
dnUD882/jRbV2l9c1jucyNt3ZYakAObVIjC+ZD25qJ3+tJ9E8USqF7sGwXpC+49bO2n10sHmFiC3
LVLm25px6SdAEzgMRKQyt+lqjH+v0+K4dGRUkNaHhVA92R9VwSuoiZCsnHgRVtrVbEETzZsGmH7z
Ym+gpMZX198/KUnbP0ysFihqZjS152WDViGlrJXdb62tn9DjNDCAPzg1AvfDd7xRo9cRGNtNkel7
juh3YtXKL3WCQF5rbT4LE09FmYrZOpjvpdpzJvqzr468NbpfqE5E+spMvux5SPMgXwtt4Pndme2J
0s9GbT4sdCyM7HrUpXgsgb7QReVRf4mdaqNsfn6fUMEMzHt9xRfMLc1tgjh6vsfUzTSINz8SQIVP
w8MNbQYyOqfLA2TKdNADYEq1hu2ypUmXkpeldmcNLuaLFTyCC7q/QYcKe5lCEKzJ7EPtaDqJDWhI
mfAyfnCQcyJLBoB0L/6g/5VfrlRMGzrB54iW9F4+MTxlrPwuZnMVsO6isb89Ejddf/5qtJKua9B2
LrFEksfWC2FjY4hshd3vEUKqDBrfzDse50XSGSoRf4ySAkj1UIAiZFQdrVaQ7bu/BOvkDZDrj957
wl4PocmH364T9+qRKXadfzfZlPcxAHD01GcymB5xHTUUAWHxXFhvGtk41v7bPhZWiE+wHFl0ZL3O
owiOBvUZcnWRrRyxjj7tcJfhOzcFjqXiJfLts5am5ppg9ubeFyA4Qp26sg1PKN1vUGVcDLwUu26F
RLBKdgFrcEp834Kv+lcqHOseHBLbIy7BALDCzkeeQbJg21Sv9EZbjo38ElrvdZJz0axrSICl1zDP
2PZgSn12mueCvjPGP8DXvBUi3y1SSnp0AnmOI2ojt3vviqiXj8RyNSJw4X99phjZfumo1IxA3hab
g1P7Ho9opUrrtwNP47iETcU0/lMtlzTwu9w/pA3S6W8JU6GcdtRCBowup7dVsPcSxvJIxdHeCF0r
MjlV+diETUhQ2Z3t//S4OawjTtAGs/ivvWKJ3jgvwUhV8FT/rZgl9TvR5KsBh1fSaD9i97srCzgg
8x2lmsjQa7grm4X/dmoCZeJKgrfVDvnlTPY2yS835mTxj9sGJl/inDEextFkweErOdk1ECbUVgQE
WVeZYR/Y9V/WNSfzTKltUMRSdRS/EmnVv0bPwuvirALYh1rMizdn0gSsPyn4CKXTemFociMO4Iq4
rEfXBUKkE5kofsAB9mECcRyNq72Q2ZmaYor/XXm+13XUFbhaM6jzevV+4GcF9NWHoB/IR5IXmx2R
YG5zVnPHMg7lj+YZ1o+rAYADTH+O1xWarAC2kb8XkkZe6UMRVRDdrM72Zd3/aoakDwKhhdJppN4N
MsIQoHcJ3pgWJTKfzfYmxi7yAlspC0/5+qcJWpN3zh1fJUrDAq6n8UCnygeMwIPeNaXQ2CKnEHiu
qJ/8z7xPA7YnIzT/qwaolngqZKvblCzq5UMnG/ELnp2Bg7lt+FggGb/HypyhvKvMsBzDR3P1YRgc
llyyIbXz1VWS4AmDbrK7CIOLzyk4fLHlCThiaPJvCVTHubsTEWX6B4Fzo4Act1BUAiWfGuLbkmlh
nk4kVLLULEEIQlG7FpViCJKR4QQTgZ7iQKSVgLlz0ZGdGxNJmsoWDCnKMUukGOaxuZckEdi89Non
J4LLQRome++JYa1Dtj+/WR6Ns4Zjk3Vq1bSf0TpTmZsQors2qsL97y2owXKGe5MqfKr0snhoNCxk
GfD1jc/LRT8wCc5XVQnIo6HjnYEwrwfuCUrPllC0/bZIdxJn+5+i3tEWV+YhLPYoI/pO/ynr7fc+
cC6fT2iR4dyzWWLIOvh8uGAM3gPW642CRsgTzWkn+xu0/xdIWzri1NjmpDME5C0yFGLAWIAWp9EX
jQ/4U83UyNY5GyY05AngQqVNQq9FcRXn5/07a6a4eeOsruKr1iJH+JYuxFpbd5VS+vSLNKSXqekV
IT3MtXQq71as8ZRl3nrljFbhy9E/WnAc7+3vNaAGjxF8xDQN1njRLiHFwvjwOP9WwWFSNSNUu5zL
PnOA8jL+EMUWQjI4wX7fehphy1wTd5dV5ejGG0GYcf+rIEuUNMwrQ/MO3d0yN7Iynsq7P8AmL9Z7
FVRTWVu97UDULZfgf1GGxUxTa4XpGWC/VgTsVxSngWkMVA2Afk6nEEJJ3/MyqAFGquvS8oqyPwUO
vT6Bxi7es1dbuzATiIiayHpHMZPfZlFiFBqDCXpTjhTaH78JqT1pxU/wXc/P2KmQug9m/KbPtfSS
qxh8tvvC6gtn67HtvOA/VDSNdnI/hflK9DQ9jfw0LPRNHZSwUY5PuRngtIoNsWuXqxspZcCMhvcl
KM2Xo4W2Zyh4+s/U6pUoGutUj5h6XI33Y5cG4kJHHhpnKeO0vKB7+kBSeIXX3uZYmTTtaaWPtznb
G8Y/eaRNt4gK1nX22izAGhH+oJwBGlrWvV5jVl6terUPMNb85qSpsGncyqk3bNbtaxvVVhFKt4Md
CNuqnIX7F4S+vR9XzQyapkqRdSjxaH3fhOneOxSaIH8HmfjZ3KjSDSBEB8vLdOVTfwhadJizs7vV
6MKGX9swYxMKwfKMGBGrclBIAPCJ5i/dSe5Lwa0ZiT3JehSbrAyz14ZU1+1iI4N++ne/xqEml8st
VKquc8sSzxZRr0CuBr+qzpLQOmkDhdD+wdRGS40jKi+fDOaNgJBCoSS+NDJomoEaWlpawRKknAbq
jqmICBcRxSfVgeM1oy1y53pRBjfAF+JolFrP4nzFcoOQBpiT+lOC6hiav+JHT9+P+9cHnsNaHuB4
VNIhT+hFZvV/Sxoe2ySiXUnmxNzx6+xwwxmJESBLzhibe6uoBziuldGnAfWtkJQC5KHtnULJfgaa
ItE4Bad3yw6p9WzT1IdUqMAn3WCvwAEYK9FKDuWgWVr6Id7IkJf2eO7Rw4ihTpXpzXUfv/JRBh3d
aHDp8Hx5p76TK+VGZGB+WknVel2zmf03xwRChF1zBFOhRQyShpFcxtEMX1fSNZTCWjXj4ja6KIF8
0xHSlqObdJClQKWVVWXK++wC73THm3ybjFdiVrxK18f/9+96liadTHf5gvvJzGYYQ+iz+xDffiLX
e1FUg6xXw5C2kfOMf90zwMCzPwEWzY1L8B1VmlxKVY2qzUOXe3rivjowunLv1GNpGGUYCElVQ3Mn
DDCEWy84WDnm62M2Q4pPtWPIE2OvQPkUJmtHfwktaIrAU4deEoCI24yuqHB8UzTZgfb9I5GIaR+c
ILVpTy8k/8k1ZtFVr53eFRR8Mjl9TB3qXeA6Cl3HeV5OpDPJ2SyTH9VE92pxOhE8BAxJtEWQ9O5E
ZTu4co5XgpEp23Ad1PXZ1aI7Amfl2oZpXoDPYCpCMkWloVFXtWCDu14lXycou7YRvvVOr5N+Qsxb
DFOGOpJGxotkLHF4fzwNNANh9paiA0hapHTYjAUlXTpFTbddGvqkE6J5+n1ug4oleoZvZW8FiBkX
vt9cVUZnc7Wa6WRcEljJiUWwkra5P4ricUOu/L1pRazvjUoCmjA3Z1A0RHjfhY02wjOSt160eXrq
5Qda8EfM7Uk/f2/gQqLGFrACpUfUcyC5gVjgpmoiqiY4nR8phWf8MUVp6L5m4wR4MVgeWbwgJgJs
nHh5ygeg8G6GRwskyVfG0O/HhDFp8rGi5tA2zK7ppxjOY7nekvwWfYUfjBAzovRWaxIj6+InKtWQ
U5BNvhm1qumNQZQAgKNAudgyQ0h+benN0TOg/nOaWg2OXCeUCnbpCoLS0Ne/HF632RXre0QLJjxm
DsLgBw1LW+I5AzVQBl1Hr7QqHSoonSULttbW9mk056wLiZ4Ww5UcJtWmNqvCuthe1R7ziQQp9cE9
FeRWshHbdPKJLgRRSt0z5/66Iqnq+XtlazG0eJex/CxsiDkKUT+GnlEThI/D7mh6sr8BCx9KdlpZ
6U69nCdPh+vuUX0147n3uL6LdvRw8qCHRYWumx43jCrqNEMrtKPwrMFHlAzdJg+5nHq1WYzJEUFl
FzH7u/U6Ut3pvgl9mnbJdLxCKwIIzvf2nMWQoTtraD6hX3Rt0ouyw+g/QZ2e6eWa7JUVdt+fNYVr
owhDuooBRkb4QLZWUWQKGvrtQnFDbSEpTlrDDXzJGktbThS1IXHcNMB5pitynd0r7rslPx0xwfFV
KhqmitLdlrAIL4VbpijmDkzMD56D2Jqi6eT4DEuDoUy/zPvSaCH6s4adslAhWCduQNW0DW8WrAFU
B4HVEB+QCko6eEsyLsS0BT005uxBGI3BUyYeg+2Aw6td2AkcDB98yBoZsKYhmEROYSjab8VpxHnV
u99Y64rTvFCZBCX0rKaZtQ15N9IRm+23wYQiSh2CAqYvgnCt0oAU9TWvOeEcVdt/9JkQzECXbLAg
7bcWS0owavPg+/ajCSc0SC75P52gs24cjSxWGFn1GoSg12lx/DQ1AhIe+KK8zfqT7MTVqwTBkMPO
x9TsRqYpBnFO764vIV+8/hZCo2cT8UrluwmHeYOTBaGtviry0fzXgpukfyGOTH9zXOs4ELisgies
T1SWrlK7BXWKKKoh0oBY3wC5XqC0MBdDcJFFeLYnrZpw1F6uAk98t+SwdRAT8qVqkjU14yqb1Y1E
aIdMAvwwx55QCywbESjL8cYZKUMs8NTmPebRRSbI+7KgKCbGOmOy8jR6qPwxZ1uzhbUjcfWOEeLt
VblYaohPZQNOPE/0a8tqNGaHMK8ok8EkN/uaWe4AUjwPZtUHZPyn1CaEZbyhrYszAXTu9XWw456M
ZPbVLtnBQRYn0Pv92sfYOYExe9Gyijw8cDhQF6j8JRtQU4YLrk9Lny0E1/I6oUT3EdHkPQJihfw5
YjwHT94rxFfjXl+lsoZgxY9kTgcghkDoFU/01P8zYldxjKB4u/VMdgfKa1Vf+EH2q6CnFUDoJO4A
Ve3WnTIR2hGUDtVhy/YnU1+XjC5BV9/gRut4Uv18yrZMyenk25MRjrKkgJ3eIJhOfWjhBYsH7KTx
m61TwZJQRBnWzvobHmacs3lVXRnB0FooWl20eSmdfzD9qdIvpe7SD813K7jVB2ydEtOrP55PfHJo
yMOEoJBG/hrpp6jSGN2qe+4rRj6fRquQWhdday5xfPGtZPOJzJaVAkY7dyFKFMxniyg+cNuvMUHD
ThnnjFNaApDm5aKpzzKYGDSUgx6niKkqu8ePbN5z3uPpzPeBVAP29Yu1/bxW+4nDQa8bBOzlzsEO
kXldmzfZONyE78p8tKlNWV3IdzNVx2dKIdZTo7OrvXeZ108nDfSCnbcPcUlmcYOqoT6AsaI5fJ/G
9g149mu8hl74L54fgqHzEtXeuHQTjZk5KjLM2y2Y3PXLbok8gU6lB7tptdEY1hsQUpN9OOroGKhO
6HmkOoVZDJcHMqmOtMcUQOWzyUqo+m8dK9pTAjRekKP/I0DF6GGEtjveOSm4AJA+3AhZI7E20mVp
uQCwnf+YQv8452D34CzesDAvSuSAnIsuYUZj39qBZ1cwpoJgQ2kQFc3N+jU+O7KzKGnDrX8eFKpo
5ixNVBcSHeTRx18UazVfFyh0FMliXZ3SySjkC1rHIdmp0hcQY0Ff9U5XFMzzV6ugtSBGsLf3FRgx
c8zAxcCUhJgj79LsACbfqfeZflnW5si3GgP7ZlWrFQveVRk/qx8fgglDK0PSGPhzIJ4uhrNQa8dR
7in3tCgG1enZVbwfyqdrE7Ly1D4sGz3KS1+tIqT81CA5JQAjdTP3WqIkUotAqPvZZ/q0MiBr+WDc
payBaz3vrz4Zt5wSesJiNEZmun3/S7iBz3bsv+ZP966kI3vye87ccnYHms8eKw7w5u5rSRr0F/KM
KC28GdOdtvJsBQz6jKi99VDf/GuCJtJn9tuqGdJSn/+TxoMBXsS3k11LFvDWl3hnTzmbHUXMVKaU
xG+y0to5dtpzrWrYCULjgn+xMDQ2NS8bCXrfzmIo0MKQ/epqkvjgnNG5nnVZDubou3bXlo1ZCqcI
vE8ZRiRzQoonvZ5u1mmq6lcjNq1jD2R46qiWaqEG7zRffo9FI7f9sT5wYaOnTUCQIe7xzwhl72DQ
h45P8FKCAzMutcSkkRXMZggXCVfMGVcvkqRkkd7iNhaFIbSyTLwTIdCXNmiz2y3/nQI1Fo4mnWO1
XQ1bPBVRFwIJ5hA9kl8eHoDexVf9af3SQOEsj3Qf8nzMEvdoe+5FFJR4bT8M+U5MkKwrlw2x2cU/
RAGaEBS9TCSG1vZA3lRRHImGeA6nRwo7oTwfL/eNA8lp5mV5RySF6SB/OS+u8bqTkm0VV/Olp8XJ
Y9Wtn2jIBr42Tm/m34+EfLLHYlEDbTbCvoeqrOe/QwhAEmhqYNybY62C7U6a4IffX2Nr+FvulcC6
pAHLWf9lvDST1ig97W5ziHxm9hGcCcATlmi1wMwwBIFU6UaORTAmewIR8faMp1ok2l48fTLtLlmr
wb764TxQDIcsmiaMrVPT5zQIley+0IbZDEM6aWALG7/qVVHVNVP75/EB3W/Uv9+Uum1dPAvPHR5R
zXehxFhwf9y9ARVUHM+SGS7Om/VTiVJE+4euZFMwMwTGP11oOo11rLtkxmU3jZ9HOIHOEzNi0RDW
SmMexXsmHQs5+wqfVb56hO6OFj4yEhEAerFDT8hKrqm/WVpnFvVajKOASjIXDwuUHSg//fOqCxOo
A+f/z3ziv0ZLGiJTyEXcMA5odTYhIR98QmvzTu7JU2WbbglZydHnslTIO9r2C2ZAEMUyJpnXAPde
2sh1/iQxzMVMSKC5kQQxei9pFu4ry/o9w0K/PnLBQHXVECwe8DdqA4O596MgUAtUhCcHn0y4xZPZ
fql4Z/zSIzpmf1hmLNy2I/u4jqwDBXEbfInkrSF8fFafg1Jla5JRFvHDziCesbhge66Xi5aWuRjB
Ts8ui1ckuzzhc4HZYVrKwmltKnbJxjFyQlnJzgtUwrzZOjI8kqirVSC4X+0KvN0Ntm0OF4KzUnOM
/fiucSPGgjgXXC6+FHHDXaZ/olh4lAV5QrYujg/IKKwxIMskUNyyLapqRG1yyv06zASkXYSF7r8l
io/kZwwjJCCLtUbK/lKZjp01nBpRupwvT+AAol77SS6eu+H6ASQFk5ktKmjXZtfwMRLHnvvcFnxS
BL9Q7HpaaQr5AJAzh2ObECSt9OUga645TrUC9zFZNlBsndrIxUv7ww5G4A8eF5c0C+unOotC3w5m
1lEzW1RrirC4h12FRzRQMwkEBFFWFVPNLsVLs+mtZEIljIYSXO2tCQnWb53f1oXdg1UjFeMzGzc0
0alRGps8BA6Iv+/0Rm445+vk+t0hfdYGPMgjJFV+mjHsoD+48w8n8QJxGwce1c1xyEINADYxexA7
ifMRLfIw0imBqUzyvl5Xb+VR3AHUMUJdMoWn9uAiBh0d9vOzkkompnidIPvB+qDHq7K3AFSthneE
ON/gXKrqlzXZ1wjsT7AlfR3R0UKwXUtoc8rw4GAfJu6bqM3FbTnmrY4McmTTSV4GgkxtnzrPpN88
e9TR5rxzlnsWGUjtd3lPWsHt3oIjhy2qQnQSKhMKgyD/ZJjbgtDeM/5Y9aRjKR9nmohMbBh+LHPb
cgHBOA7HFd/19Y/wYmFkp/FMPEOYB2nKbgwSpS07wOTZqZLc/Fy3E14GUlIY5b59YA10Yl6qf2t7
k2o5tZD6HBRlhhIhTH/3YWNSueOgUueumBU5q6weLo0wkGQTJ5BQ53UREVPYragUiedj3m7jmOCO
xUn+PoqCh14+1hk3C4gvDyPn5ps/Hn0V8YcaZWtLqwzuofboNTc23eaX11NJbuxrKNnDAzxfdUVc
N9k1LB7LGJMmIR2ZwjhaaC/oDqadBJdhWIrXqktQHzlqvN8sW9Z6KkZT9cU2qam1cOCB65tccHYQ
rBTJyCML3rHDmcSXYaLV2h/1flzX7kyzOjvZydQ8YDDHUFutCBV5r2xGxxErvDwbabaWM30ORtgV
DM3TgNVAjvALn8QKSZKdAPWzao1cZBBL0xk6VB29etyJvNQvXCqho2Le2jhmRrnDcUKB5+NvTtNc
R9+bOS/aKP+hwrH3KN/vganV9hKN6dXaWHfryh70ggnOZx238CgMEUoI9Ud1C+SfYrShyKus5HQL
VXNMlz5A2LvXmQf3X5NkPm0KkkM2XOVPZCie3aM1CNMFEoIiOq0P9HtDS+nI1oALbdJb/iYc98ek
G6G86g1Zfc5/MLbDoaYTNBXeqRgZ/d7uz0OxJkv2d39oWnjXssR2v1iV8IgxzZXnPj+W5NFfc/CE
LT5QnpgxhqQRpdS9JBgd67sr464sWmiiKAoCR0lTjXUiiuGoxwqu577H5nCPIiSRISHqkwHZ+uWY
zmhvYIrx4sFwAel8lXcxoSJQxX7UMGPd/8ax4dMPAFktaS1gb3qRUCvhX7yJxwoaTL/Af9iGm/He
XsT+kZyZ2y3W+HsnGx9KUxyGO8GpZHM5hF9+xd0XJ73wAwrORCneVhdZ8+QY7/bCcYiFjMPjDszP
S5Vb3b1JwzKgDkDs0sCiNEDXzrgWYqBsHRPr3+fwnfJxFLy8uvsmM/IPzZBevJpm+2T//9hjUhnN
UL4pGnsNGek3nDxuQFuBMnSJW/CpqgDZ4fhRvzNvZD3B/KFa3pdANWVFfayiRGDYlXAbP/yY81ro
Qr9p7yx34BocO4pq0ct+32U19xYjLsC3swabG4LGff9IMN8KjlVUwQdUguOwTSqKrx9J7KHgmDYI
A3/o95E8M5eEYD+U2Ln0OtguY4yQJv8kRPAao2ealAEDW9wbapHJSvKA4kSe6eODkAYfBSUK1b19
xgtm99urSggMBlmIa65kELe6KPmrSFHgfxQKiWgiFYVc+fYOm+CSONEgFPTk1/y8t29f1DhWOmhd
g0a9Jfe9pMPpAIjW2zIZWjaJuQSKszVRhTjXUinru2w7TVfUUdE6ynH1mZlHRLLtb62pD92JVEg2
GnZa0MMjQIasF+aQ9KvRQJ/hww2favf9Gk4tdLKNEJgvhGOj9cuBU7c53N3m5Oh7eIAuUgKidyFc
UnMEnU/XZeU5MCp/x/ZU2m/BNSIgWwYI2BpgbWUkxLKu63fFLFP9iN9UhRC+hhzTQu9RVONEG3ey
aAyfLnoNMxqC09O7JauXrPpMX7uKwS4riJ6G4O4B2AD7XL3ft7cQryakGrAQIadib7/GZhywkUo7
/+/SeokxerFHFERh8/6o/NPW8NmNus59spzjYAcAA1G22pUmmuy7WXYWPA1U0S4fs3axxElA+XgK
zThuYYzSewVY9ENwcrGp3nVOfK0FhCwfg6nWYrFyIJWQg6OWD/rXkVt9fBJU84Vy3SEbJqjxq00i
Y6Am2E22X44htjLfwAISjKK4HGe/BgOOCKCzM3zuQQyrv/L+97ZZmCevo8GZ+jywkaStec/R6IJU
lSHsYp7zVAoDPJk+bFgYdfo8kXqGFAr8lScwuTy2aRxRAOmBuxK0i5BSjYZ80bni7xetsW2D35cY
jXcxkfHnx7jSyiMPsLAUrjHWeV/YI9OxLVHhg3uvA9k6ayrBW6kMMp/ofmEAYZFYFvDO2cu3P+Ei
MGbb6o5k4OkfdbT1i2/cRyoOXRlT99IzIUgzQ6pFYRYCjlFd39EGmdSOJHnzr4Kllcm/0UHahdb6
r+09eOeL+BdV2Zv6JQ/gagv9mOrVqsE7ReY7QHKOed+NxsGimbeq8DTZlQ9wzvE2tKbTjcb7HEUP
dGgHSE4SnVCfZVhvpR989IXBN/8S9ZcF9TACwVvZaw2VD08xAr4okIkelduJeiSM0Ts6HACIrS1v
B2mS0DFE4k+ZMQzTd8qDx6zLtLchBd+JO/YTc98xLyP+txmMvRxO2/oxQyT1VLLoO/rFtRHggsXU
/CDCxHckeFLoj9GYWEruysMW+tPSgaFmvblCUMDv+yo+QyfWaJ+2VYC8JP1VZBkQZeVbSowEtKhx
5HMmGFt/+vqkBfMA5GP1yutpzlbkS70Q0ZHrVyJ9B/4YGxVH1XFIE7hG0aTXTUu1eY1XOegZnv2l
+Uc4pHv32kZhPj0UB+OdAqxMokpWsGXNKznIp+kP4J1rphntNghJLFnEMhzfrP4WFATQMHw1FTN5
1qsB6zorkeirTcgHvg0RDMvjCXb3hA9SNw6S7H+1Wbgt29HoVKiYbqiz76DwS657XqRV5TkF9sdA
U5CAFhkKuNLkC74RbCmFraQ+DGP12y5VqYns1gQor8rjNbuR2c5vhoUVK0hVWaf38dm5YOurXNLR
nG4N68QLPcnc1ygFjv32YRKEGutdv6hzfD8CwSl76hbxMrGxKyvae23cX+Z+XkLk5bCx6PlHPUtZ
vca8OhPrtug0nV90kphbEvlML+KmkCWdrUjBSN+YFsuOTvxF23RzzhgiloTLzo9h0ABfbeyMIliH
pG0XMjuWU+gkRBpVnm2og3ySf4NrT/mMgkUr9cFiE/Yi0lFbbKdSIE4oYmcGJBvAKEWGUTkNTJIV
+aoXmPQ/CUU4S+VOKBOJQqcdrg9Ld7uBS/wgcP++xzdj1dM89zrHEvBEr0l7dGpzFYyKWVTmHix4
UKo7oDGVRNjHo7TEC4aWzAEJZTQ16gM+mEGLxg5sJSQIppOaPDv/2QneecqSip/UJroCGANokiSf
CEOooAMCSN7bZ9M2uh8Gg8j5Ci8Xpgyr92nBgPRY8R56CRwgc2VzuM5aGqqEpM11Rck2LEB3qu7Y
o80x55BtAyzrj1PSr0njD1ijm0N8MKXGnOH71vqstHuGnWHfuIC8VThWS5dgLSQyvbRhb8A4Ahit
9pkmfzQXE6tyQ5ny7oTlNYlOcfZp75qkKTqdHoLoAMUvZaJUseOXaPI5UosZB2Vya/dma9JzZ+hr
zLEfSyCgAkiDOG3Op+l3tu3SpL4bEnBGCcTuHrf4W2p1kSnCAKdZJXrO54FXXWkt1pCGhAYGeOF6
QUq0cwMcomDtD+7bFT5g2iEaIAHLuLCfJndmUSDDkIQTDoxHcoXKSo36lDHaydCrzyHLZVZSWXCT
L7D1OVUiKDTKA0ZRcceNIGQkQjjyXCSR4RGzysiDKexOM5hcBAJb7kg8olmye8R5JDWNqqpzhjUr
M184BPYT6T4hu7YPnjehq+lNwBv3cOuIy616q9/V+5VhUr8eCmZJETlg2Ic5WUMHG2LgYu1auy+j
SIktFKZOP73y6m7H2VNiQ5rSu3d3MJKiwEH5YSecDS7LJNi7Xk78Ae8GtYn3+lGw5mRwinPrfOso
L4QbIM+7h5OrsBGgSWo502e3J2xHHTXC0lN0imJRhmFToWT6v/mnOX2TGoQV6fu1A0SOh28qEEHr
6NZPkkLGYEDonRG9trL1JHXiAI99dN8QuKbob8Q2YFsPWqxfA3bXBaYBAX3z/C5EibamGcfuXTP3
EaWT/lraYNbjlE7HaEsUMQnH8H9yIT99LFSaLV3VdERyRLfJQ5x7q0uj2RGC47SvLBEL7Q3RZYcM
Xvc0xFc4kRw9myvp2VbfdG89QWZhhNQUTIs6S2ZsDt95tvnmYsBzbkZsDh8KvDDvWyTKW8+kKW6c
+FOo4pOKPxOGVL7v0m/pG7Y1j9gNvNgfZoqn6ceI5M6mmL974hypIiHCU5yXGrjaIfQKIctcz/5a
2rKVO52hE5PSiFde5dL1zna28vFMYmZNMZGyUXOufLkyqvI79Xmccw09+UBwFhTHjpwLe9s3jAEr
pcjdt8hvAuOZ1UyXBJRV+d5fysuAUQ7SZ3Qs5ClmBSaOy9ZkIZJnEXg1XHrWiykTXaGtlk8/G3yG
0JF7gEKDZ/I1ea2ktKwpR4xQ+rlJHEwZH9xDYtEwr/KDF3MZlkH5P1yJPqlDSKDkU5l1+NO1b9rh
7jLEDVECDGpBeTCMSjm8knuiAivv71V4F6mj1iu/4gjjY1jIh+bAAy8U/ftsB6NYtti3OCOtVlII
UjJjiXd09r9ncAZgwn2wPVJRI0yG9lDk3wbtfvtQQEeWS9vXO4FF8Uqgqilv8ru1iUZPPKoDYM3Q
P5E39ndyHVj2UQQRylN4+bRaQ7hveHzyP2dZXFgYXNvDq3NHQed+CnWuxjUlRZlgDVMGic46ezqH
AxWUPaLqNzWdM3B5GfqSM+KQwedRPIZnzTg9njq0ci8CssXP7aVaJV8TSJhmYrHh71EtODuwWSxO
qLt+3p6K8GaUian2txTDECUNhKxMZDApJ5HQO32T7zoZbyGdTM6rhJYyeVWznb6F+wHSOgdcaLL6
1Zc15nFTfKfIPEFmBu+7W7rYHC0I7I/Jv+EiNXh+rjVUvc5RMNdk3cI0Kh8ZtG9rST2UiMpBSN7U
x3/UGKS53MRv+n8HDuDZzpNXbiwLFM4k3JDK0s/RGW3Yi6jVqU1imcOgC6Ibk91RqlGK6AW6wdOy
EV4An15FbprwSaWAGAQNDYX+TlNu4Dwznft4WCcLIFxuU8FLwSwuGLS3vXUTRdD9et63xKpa0aLh
PqA6d3AI/bQIPXwlVzIAoBI5Q1hvWoacV1/NtRWQfHhm+/SZ77G+Bmp+dlxwBP1PFaqi72Y5H6Qe
3yUNo4uEZZwHx7YrLldOEq+xLx33XvFSGybq6V9I+cElgLbBn2ygcVEDe5DfCRZ2T6cbIUWzBvY2
utEzR/iBUetZeZt+Fidnd7nvQ5O8oq97KwzhHockvUb5zeysFyRu7WSLwSwovpep1RyR2o+2FRo+
spJvzizPThEtOX3OE0PoZLPswiVQaUmf+FIh8s+XkkM4xs/TAYLdv+abGqXU6sDdi2c0NpfC7Afm
mpQCT0eJqL1CibMd844k/K95DA03rviw6kkoMtM66ELsJNgzlLwADBvJ2R3u3MTSGpjnnDAoHkQz
AsRJpv/gWPwHp5WZT9+oEP931hlDJ6JJWqOfyjwqNLyuin5Z7+EI33ciCHGYBIyeFwpM/T4PTulW
8FbqEJ6GTbpXd+4dJWmip14k9b5TXOPQ9av8n1BoKAJnm9bM4emT8lHtd8plBlWqZshn7zBEh7Zr
FD1lDyWO9+lKYM1/Ko4y7RF/Qk9ht0byClVRSuPZjwMKaecGf7Dalac0aq7HNdVeWuxMjQJaAr08
7RIz43J2CWTRKgQi9WiGQBz5hK9YOl7pNRh0emAF+aCWRwhxd1kGaogXySklXB+bNfyqH11JkJRq
zZHAsE/KKiRLfv7eof0AfsJn4Z6qQtTXAon8eXq9pYDXj7WZ9242objp5lGJwDH45BqNsnHnM7hw
42f0ImOJeS7+tk73/SPh2CG3X0MeULVY+4A0G3F15dwG3wf1sHEQMhnUnu6RKXxrCRdOyW+DkzS3
NkQ6HktoMp0ba2CObhNtDK4s1bgpVJoPXwC0CTQtvcJb4q15EE6dMuNOteLc7q47aetRPnTQqqLu
lomAHJxVhqrwcDWVl+gMeJNQW+3o5pdqw+1Zln1ARvchAaZNOD4fNUjh8Mv1Jhxx8P7KJCjDfA6k
2r0Nn4nM3OUcfuhNVLD+2eltyuQKjbHSpbI5F5hfofsE/TdI0kVWeAp9GuvinZU21FmQ1nNXyL+1
dISomA82qBlI2EY4GHJWJk6O40gA+eTdRStGDF6hDKPwIJH6Owm3DNxLant/NSuDGSSiCJsA4ZFF
6f3ztcn0+K5NVzydRJEUqplYkAJlcLc0xlml6ykLvAWYzWz7gz+11m5P5j8YkVJoTC+rTsFRDKtH
ATIkvChIrczbFLOCHGF9jNxTnJ3wcnaDWBSE5ilzDXjqs4suK/JULemRD8CVGwSsJdCDxoLMIiDL
eUfRu8a4/42A50BfRdkbaxQFMSiw6oT/2B3VdCe0uSv8xvKDuhlBkDm1tX5US4OetovslNBhOuSg
Ue6+grpkU6lQbp4oPuIeS+5yCM4DATvCJqfdV32khCXXBM7vAiEApUvLmC2S44XymMlIudf31H01
COJoTVKITsDp5Eyls4AP4TzQrcdjTja/NyJgKhFbgtLeoXzt8Ylo7Qdud1cYyAXuaw2kQeH/V8aw
NdxmeGZxxN/5hZgMBuOUrUnRpq64KTTP9kbyBTBqraUXP0GtdNAWMCvg38sWEdb6rXq4UW99OArQ
XQy+/rKgqPt5lMyZ3B4uWs2Z+VFfueG6IRyM2czwA0ONygRg3/9NXBkYzXuzF5Jcq195OrlfmTMq
2ql6Mw/M6fzJK7p54zBSRlnyPtuVZKm3nZ4NBZuVd3GVTohqZEkaFoPhwW4ShtPOSzhiAfOeu/SO
npQUxrirW8AVRkFUFAfeAdxA97FK+q99+iP/USBkFT4rfnuguykxjbOwNFF3NE687FNo9/IO9kNR
EEncpJAZwv4qxEh9NBVm7aMQwFd/VmeVfk+K+O9IBUFfR4oo3XAdBGIwM/f9tJqSXk46deT3J4NO
TwKLHXCp15QZtZFKuWaGNPq2Y22Xhopqf1JpusDRfrcCvcfja74Km9wROZT6eXrnu6iKBZtiAW5K
8iGNsilr1LNKhGcCk+IogO6EieDjOiTpeC7/tOPIoVVBUmPdtg14yDVHLbYw5ChmOnQMMIMFQHta
MqEAahm4aV+uQwqHQ+bci4NKhDjrej4MgXwL8rPeF5k7TYnCA8ej3OWAHe9avaA8S4KI4dRkgFE6
p0FzJSg01H4S1KAwz7lor229skdLm3RAker/yA5utkkPwE1tpGU6HTeh3xKRT+y1XD1g6gaBzgNb
5OMWMQ2cbSpwbIC44FVcNtn3U8gtCmw9glanmEWZfGNUSzWyGfKjkE3YONgdZPhckzOSTkVcI0Hp
VOOtFaBLNVnIlOGxPodLBxqqkpo5mtjatUom03NBARs9RBHzurXH/41952wbkmN9/06E5jJ13Z2X
EQ7+/BFieOoJMO2wua/Avy1ncOTPxZOKuzu89YtHg0vqN1HEcI6l7g1QBKbxhgo0J9VRecUv84ZY
EfQ1VrtCkHyVm3AoMJoS27DcY+XoIG8ILYxb6bB8OngZFE+kTRiG8/DjykBAPviZPtmlLD+BecVF
+tZbq7URPJ9vt/mN2sH0PRSFDqUnSrtXANe+N+JZQAYnl0y0l2XWH+85U5ZPYceSKrylt0G+C+Em
ouTAi59GmPc1qcZ71YJ1U20MtaVuNoG/JxLjishn8k5AvbhRaLnbOkzF380/dypoNNjUKLEr0AtP
zpYqAa1+mjbkglOcDmdw3Y9LMbhQnGhACqdUdViPP5t8CWfzoCtBef6JXw06SJ134SiGK1P5+SCk
nhWBZuQUkkpKnlEZH0p9QFHFu+fcxKfS0B6DdL76grtijHY2nY/HyDWFqxUOI47ysseRJUt+CojE
NWU/utC53ydubG9/gEsT55rrmjNP6Fuo/wEB49PeXoPBsxoKGMT1sN7aUw/vGQruLjlibk3Tfzgn
n3sGShkMf/VXK6axS6/xAPXs+iLUvDw4MeDvhSkzqXWfYLaxc8TAzIBZEaxykaQublSj1SbbWRaD
tbJ4FLl5vxC7KCp5KY8P5v14+aphRwWhZb5VH+bo9vEl9mcsEpXU/mhY7K1qSWHLENrqWY35pcL2
w1gS24tpoeR6bKv/rwqSdPkOOiCUV54RFziY4+OaoQnjlaBF6yJ/l9D86bP7s41fFeIAhkm9N0SQ
TxzskeW3I/pUvFXC7M2/5mZH1dLIkeeUoLnvEQjJWxN6Ah3LuGYG/rBFnXnBvkU62TRShN0kiO3g
cjVMmSbIR06YmZksejVqhUTwzJVGfvtZ9c7/YWWBoF4Z8RGK86VoyHAtCf1NQu9enxvIzB1Lu7Eg
2OF607Dbxdtm2wpUFYoGHgmM5I26cAwUJRmPvERjfmlVCKzxyogIK+bACrMyGSkF8EJOGbbQTdM7
jQ3U979tiNtiuRERKEwNyF05OvIwvWwSUAcYJjELFrw1FJqRqMBvjS3Kb3WA7UrjT+RNdw+n4IB2
atgRgFJZa+HKnBoQ25VIUMdihCRFw2dMxv0q/nHmkOVFp8tbbpM1hzkXOUmOKXBEdZQawSJgj+Bu
xcBJ3rzkBD2ZoCTiUSE+c9KdNRW50sEFJfZDn1szWlZKyEmd8/kpvSG41GNmZE90nxiRyEHx6XZZ
O2AeDewBUmqyHOcTo1IwDsBSGp7x9aocnd+yvA2dr1ALR3uvDUdU0k/6Sxj99T1wp0mMkIYZoqAE
27YX8+N+uh2XMcjotWt56ktTBKyV3NvjarC1387kisJOy0EunQu4nz0MrgyJ8XQq0VokPOLfofQg
nohw/5TdxQCO9MjO8SPNIL7RyttGljp8Uo7a83my/fJGtgxF4TpDlw9VvD1ctNxGSveUpeDOJp6u
SMWY4QhYTHLpTpehLnqNIWqgeCMwl/vg0hkXDxNFJyb5dKtiUJr82K/W9D+MoPG8PI5B5RyW/0ZH
3M/EcJvDx9qHuqhjhAMrvs623OB5XQZse+fswP9tK/5VoJscbwpc9CTRmBtYUxptO3W83fHzv1+G
95UTl5vnBY2j4YnKWxUaXSW+qIWRToUsP7n/zvEHmjpj4oO2W8MLevm+NrqwaEXyUkZWPI+g+b5R
2HDxUfsGFc/Cr/9yagZpnbnMbAS2Si6POumux8T1YuH9DWU05zUTpow/TOq3G4JNOhUUEF99iP9i
Iha2LytRLcvKe20+W6Vhtg4HnxxMptNe45LXsgDKdFetLT7UwdII2fqwDak2civ8H1+QGv08vXRa
pyk7ayQrSrbnfLFRKB811tDJyOU5A8Can3DRGpf7VDO6Ny80OZNF0t7DzJY2AvS+l0z7t13LXOXa
lY2kM1po5SRJKVEax0PpJhmQmIEGwUXKWNgXg/SOHT/2ns2K98QNJ86ziV4p0Gpd/bWbOt1b2zBY
SFHojFP+Jn6+OxiD6m2LCMlenGOXqoDSbGzPWAN3ec8BNGrt/WEiGcshQa1g5hH5M6xji7DJR/GS
ja02SIthiYhKBPYc9rzywCcRwUyqL2dKC/fWbNn5gT5VhkLHwcd9/ucSOViozv/hSde+TXIOlylm
pmXUnVPgV8ijVJ/7HyopJsfOtQE2/z9crAkmPEa9Tq+2AWlwdxykHDsjeqV+zbNT+GeMUrTMwz/1
wR65TWA4XIxiWdqUkxud3F5nLK2SnPxp8I/YZrquCE/jounif//pTwVCEMGlt7cSevjtaDeUjcqF
WtkTvI28YwiQigTFmKLlnQra1u08jr6lLQhtuuT9leBOguHjG+nqHBgRcz+iS+U+5Ol5SKORyeeL
1MMnyjt1avyf9kbLPgDUNg6UXWKVZL5kWhfw3225jcg51061o2tGYz+03e+q7Ayte0eI+juQn279
EZ+U3VCA9XTUDGMqnXtcr7aB7zwufzzFhZI34NlGF4k/woACU5isxyTJQ9ewYekVKD34iTTaY6iW
6jzP9iLDpuRxfNMe42POYzgFoojeZGuWqtdkgE9EeoXUJeekXePvQmUwJek0Th02eisvGSK2l7WT
IMKF60f6wdhTd+YPX77iylTtBJk2O/MxAv/Iac9OgpYkNiGLTGABIK0rtC3Geca0N/pL9OUXo1VA
cN68uJGchyM7UcmsfWCFRBb3Ce5fg0eeFtU8OF0zyxBatbd05Pz8qzh8tp7cAz2E2nRAWrMCEsSC
73o2eE7a7secOAz9djRc7qynfna/qqBVAp64LYIrllRuYfWpPK+zhmNhUHR99MxaNylVSjo2PTtA
20d1xpO7kM5Qsb4Ze9bT7X5k4gOrQ9yuYoBWYQhiq2kUahhX9aycT9q9H8lvfEaoL5Gwqve+pd9J
rcIkqLC4JM2S3mX3DzFbBROM+CxbVgYEJ/yaYJJlqPcCRJrl4/60U2cqL8SDWUrEsDnq+LQrQ5Ch
4ELYGfkXm9wyDtVTzJMnzwz9quxJlEmIj2H47+ACzt1ZtbNYxJ2E0uFtHNZRqvnvh7CEdqb7740M
ODps/sN2/svEbNG9wCpWiPEXEGJN680Cy/j4eeINVSWjGHneOA3HPnHMiz/76QabTyEE1RXrorwQ
9VRmJV/mGbyEbjO96aP6MH1Q3s4ar9LS6D6HBff3cb1WdWkjSOTZgMHO7C0iR6glkB8FrQLFGEV+
WfKhXx/p7nUgnHlvxzwaQk6PIQcA8SAY/rGo0Qs4FrBMoWBaRWgh0npPqLXUoeFvga9hWLwTi4Rd
tB9sHZSCBmhfi4ZfHtaWlw2phWy+LCAk6CoeIF0zQt79W0j7Eo5CSGm7bCFTkTUJQlMZ/i8kFx5X
qqPUPixOqrf+1xhiIWPvHrYvIrr3iF1fcinkzmnWvHBqLtY2vZBraGbIEavrvtnOE3Etgd7ZDQdM
kuiKaYfNKBOzC0QOqos3+wVE50uDKWRqj2A8yWHYqzy4oASy5CVWhpFKU26iwnP5J2+0tP5EXpVf
opzBXkfXg0fHT0wgEvguWrcjT5wyrBWplh20KUBMJxx41HqNjCO2Ujp8rl3OwltBSqdfQskWgupd
ngdrSuzi0wncZI8FHhneHAf7XRhJC5pQpQRtqbn4TpU7Df7Y294iXbzxn/W6q6tUegVpV8gKUG5r
rO8JJTlXXc92UhPjCNOO7TOG98A1QDv/z11SNb3kOQS34gQV877i8sDalbHi2935UEbpV8cE9E7X
kWG4q/Qd5/PipiNtGMBEzMRsQyZtuthOOLPcewsdUgDPzJC05Su1JBclbj4mTyogYp/XlH+8Umt0
s8L+6Cl6TKXQAqd7/hFiyalyU3JLQiDcBuVel8pZGIZ0oRcGgTmXpeIevOF0Y5f6HtyypvO3iXC9
/GK9BwwZCx8wFp0mMwAG6IoyS8OaEf8rGbV69p/cf2GFJU9XDdvSZ1X3kN8Cxhr47EmWh5atOCU+
64luU0cfU40a7GIG68ziq+uyp8bS8dPY2nql2aEik/En7EiN/tKzpgCzeMJRLgftbi9ZgSClzWwd
O72jRDt5AilE2OaOrTfrzbTU8Nl7fFsQl1CnxJXFVgRnZikinwd80q12Iu0H0B38VCOBsLMNrTRY
3o7n1Nq7Dz+OevjolIH2Z3eQQioISeZrqQb2ZBgqu4UgyBulrmnP/Nxo8g2JxlL7msQNCg9J08JC
0sn5Q/50bu9kRAQ7jJQZUKONLjCCiwJg8PUL8UyQtQr9NlsMc58x50Fj4CxzH3ZCge/NdJjq2IWq
yaXJnwTQD1ukI/PMQFkHYIZeX7v79naZtlok7vNtk/TRb7219wq09EnuKSY4fCCRx9ShKZ/4OxzC
BXT+1xltpYyDNkTKIlCzzIcRdFQ8ogOqOD2KktpLmb4vp70HePbf3WMt8izmMlwZVDE+8jubyVmR
ekOKrdHTL5DY4NlpK8na8mMDtEc7gg/j/FkW77BiXNkHkM9E0oMHGNxc3mtxOfmPC4LmyEPWlcDx
FkhytraQ3vf88Ubn+KhE1S1YNuki4RujiUP5ibqtRbC3Q0hOdosZAB3PrxLE5ULe7YXbMdeZURiy
XBcYXG6I+HBNbTIgCrS0M82VMDt005U4Pi4vHiuji53d3cdhGUZVwkQ3tNFjro+DFA5J2B4T+7e1
92pKnwAddzH2GnMRvL/+k9wBMKVAZ7omsaN2IKi2penzNU6U2Vc7HsQJji2MLly0RGNnjvhRadfx
5w7nlIcG/hdEKrN1oPvgGxGyUHT/np08vFC2dSeDMou53KzpEv6wqY8Qxkc0j2TN59cp7VxOSyWk
/6wzCVDMhIJtvfbUKi9r0UGTmFtWwd/YHxa/ISizcX0qTR+s08DhDm2DBh7Ip44CQ6QkRRdAPYs9
URDkGMzKCfM3+rc10IsIJpjv2jamVAFrYNgM3S1pkutg1aajk9LcwPMnvarX9I1SslOPoAjPLcs0
N9e8u4lUIrPykL1+BBeQI9TKE03s2Id7TeBMz026VFl9JFGOtdXBtvy9aVzqD9eXAxQdd6KEvDHN
mETmVsNxo1h5h2136dnGlsUoTebm1iw03mPv1yqLEVEaZiTibSHYo8U+2frTPme245ptu1QYHzHl
+WgIEij89SZNViiMs6MnMfpOCQCbM6PjSkqwhjDgTDYcDpT0kbHW5TkLv5usIhrsJw1hI3ikYt3C
2r4Se/7n27VSOJjQq+BqhqZYTv0JVnMnB1YAkjXqQM6+qkxEffWbajwcdvk0/xnn+ddltF40Gp6S
GiKojMI3BwC9Bk701GbzO81bOaZPxSxJk3MVnDsuawDt6TNJaBVkxLZRUu/dWAAdwAcsixk+pDLX
EPIpLJvkGrtQhd0iK5+h4e41IB9LG13Bc08OfCwm08904XVGIOOGlPjI8eW60YDnpPz6yXATL+Zx
I7WbIjog99BwnWgwP2jILTXiH4aoSHdjuGkYYZGs4b8qzV2zFVZB1INXK4lnSqHPdmEIKQyRP4DH
cLFZdoIrxEXQNNgO+cE5TfNDrgBQYmgF9ZmAGpAMJoolrgrFMBOHpvyDXCyoYpWcx004K0d/tNQg
wVwfOScKBC3mZ7cJt6IMk9+CuZKr7ZnFipufyYdCIU0oLmEdA+JpaPu19M3scSLBTAXA5+yeAaW+
u+T1L+TyHrmsqZz3yEw5OU8VU/qKsDNDgARkv3qZwIzJNBMzJbw0I+sH9cVEc1ZV+7V538tXXfXh
JMfqsGDY56MNwVxhxN/37ymu4szo1VS2vlV0m5PBSwv7pCf8KFRMhZiNS/24Srt2lPhdoXO4HRdm
PDjj9LF4bhREepwZMy2gfKTlBj1Q+3HgyF2TmtYxywhNKJ6FzeeftKik0dLIvNLHP+1BY7Deo2MS
ig+TLUv+tYis/CoKCOeTvjoF1acWFGG3Dh5iyG2pWRwBNizEN/p6GzB1OVmDIfzQ0EF9rNXCu1Kz
aGJA3eSc0v8lUBSj9mPk/Rrz+9GCbIcff91XdaJniR4Rp4dJ5qhJX1HvB1JbQyIIOaa7ZnUaRe2h
QuOy38I2Bu+MKfpKDPfOEYHTBgf1lhy8FqoB7QfVQe2y38YqRM8KPPWxuNPdYF9lS7jhNZPn5Jg+
8w5kySuxyV3I8J8KjluvCbRxHZ6PaMq7tQ3NJDldn36ZFt8HKCjgLFXMDE/zSni94H3JTzXj9ER/
a8kb4Jk+whygYfcqn0+RTI7AVvWL3JLC+cLh7ubdRInq8L9hXKsTK2oA4EFPzyTcwT/PbwwexlQQ
gaPsSOL8bBlt6x3f+/LTenWzn2xc2wb243zfsQjyK39K/1v3PMtlB8ZNM+Qy7e5CZKW9sHHcrlqv
Q2CJHjiV/DMyk+AcMTVxN1bbFzi7EM5zYIiAmIy6BHa5Nu6sOtgLpfDQ7xAM86KDygdvSjtp9EdN
EER4DJoq9XhEJ1ZCxGl8VscBt40vhwDwq2yB7gquD+zOsn4LbXKDhZtdnQ5FpZCW661UgbcVIO/g
R62sPtQO7d576yDuRX/+eI6p9r363hDec4gSMXbKgoKG2CWcymDcPZEp6SNNlRA7hrQhpK8NsDII
zesfYDcty+DeoVZSNmBDneLHe8+UoyaI9eQ2doduwMYE0sC6TAUbzflT0bwxpaHm0ZcBW2Ayw0+O
hJuq9q3K21yrpgCwKgAjog18EG8KZifbl5nbBXN10gO7HGxVp49P4UkcUpYaNxcG5nSCAvMBeyXL
jZ5aVSd+LTJll7pR9pSbdjr/WG1bQ3QoZsTeFzCfIxzfT1b7XITQvYqxcEX6di8X/UW5egtnPglw
wy810p54NuMKbstknsDZgb7RBn/7L3ELvKwah8oCYvGxx97wd5AWb5i+glE6GLy4iZa0e73b1IMr
p4IZov10Ng2oWDoYVih4Dz25eof0MGOcXne84HwH8ZrK3B+sXkRJpzacreTDjghQOg0JPe67pihD
RjsDN6ZiK1K1T5XCMs4utYHxNTRmPjl6FSVik0fD7T4qmtbN34tORn+Wk8po6mfZL30swoVW//9L
R4FMABmSqSLTzTgAxnDU1cTyKRXJAjCHKZG3GcBODmX8XZGLkswMc419JDnVJZVyEvcqOlwUL08f
Lw1kj6VdX3t2iopgKIzPWIpJ516vb4u8ycB6NilBk5dycNuZi36k94glAqsO88MBJ1W4rQUY5Zyx
bo+WnENrJMNDoCEB23gcjFlyqEFiCtCQto/K24LHLxO30zEh0+/N8OpeXCNBESIAXPZZDSrS8EvB
oNUc7xT8uQQGIio8NEjAWcdcS9SUc8G63L1ZODYG9T5JXY43OCBdCS1sVaK6NDA4lN25cUkM3bI3
hkf6aROOH97rVNmb4dbLk/b2Eb+bodTDQNZYA0Rzco6dtmyGenRXDjGZMNQNfyzWgnFP0JRcQVTA
0AF2TTPyzyIIc90w59iEhoumKzs7A93X6d4pAhYFQI0gTe+gm3WUSjFMJ4wssoEf2s8sWddSORau
2unl0iNsIpPRdSwJcHyvqwNJ53yp5/4EmtmgIF+mBE4W6Tuf696LpP7rBC2RBni5ldha8lDbhVXS
cCxEyeAwVSj3DmzfMTku7MumBjvLb0xZu3zR2USQq6T45PZCGmr69oOoy0Z9JroKjp+EBmZjOCy7
KRNe2BDNzHkOyWQ0d5q+rz6XLbsTlz9vpIZaw5XzaOhK5XANOZRBxQ8ObPElC0UAjx/LYcCFZoVr
8R0RXv1TCBDqccWaW4vaZMunyBVIuG8o/NsbC7lSmtlDH0OTzqSjURvq0Gem4UUSDk8vgtB5WP48
tnTjSAEivMIvhT0s05+y5S9ay9DAA73oyEJqjZiOGzFZYm+pumWGYJm3nDcSPM8AI+peUyz76j7B
QdMZgik93c/YGtzqkWI7FVEc8330/4VGjSF2Y+BHfFJ3uH2RMKfC17wffZ4Tsu89InH1CVliP3Dw
TBQMx7YS/0FVHUQHY1z2y+i1PZThGEFqSPSTEpBo7E1ORu+o4Mndb2zTZ7zmkJ7OOuDpFyJ3/n1+
Ylha13FFqOB9f5XNTfrUX0h6RqtTbhu+I15y6sOSQJ2o48HIZ6jov/pJECr5ukbon4jKfp7QrNlA
lrNDsAkNAoGGNXwH3b3VoYSCIaCkAbMa0LEpgeMX58/Ebw0CAhIumYD9/DrPpstO35ckrbD0FGGE
5numMOY7AHQeyDjbrVZGXrVX8kJ3mRK20xDfmKc5QdhFnsi8Nz9E5x4xc1QoUOpl3Gq0LM+P0kTf
YR9xkhwHS2WlEUlbUwhszbMslJFAN6dA2I54983WGoJJfZp9vBnyrLysULi2KC1t/k9As2B/NE12
BqjpT8XSGzy2QKK0pWreGr/1Clux1vIEry9f8f9b5pO/ZsuaJ0CbHPbWVPIMLt4cIvNUnwlNFD79
5hqgdUdOqVMqzXPEl1jYUhoE8PgTkVQloNiWsGGRrhDsQlHpQ4x4YDY0ce9RdM8rkB9H+YC8+ZtX
LYzNvw3iRd27keFAZLQbPs/pS/fBgpRZoZFkV9WTBC7RlOwlOTConqu1rUZ1Y2jerS7FzN/YzGYr
PknzJzCZNOjR+3yRGlAictpC6nzvEtceXBKizM7BitM7UDi7iMs+cTzgqmx/IRIWqOT8M3iMICTy
+CPjm4Hhave/71ynvIbaasHdyMMylGrDjuXaowW2I+WgJQ9QNnRMTejvpsoB11J3lasxdlCeIzED
9qSw/etNnNvB1rXRO3Ant1fkMBK8UGXhh0urDM53bNSPaAUK0BmXyOmg9DpFmNLrAqvv/aY3MRD1
ieo0QF3gydMXBRhapvN3jMbebSDURbNpL3t93lJXqShhF27XM5Zr2TfhsoxuW6m7LskbDeexamqr
XNOxFcLT1ynDHL9X7kf2A/yX+4klHTFy6r3Gf8sS7o8d2IMR1cjMg5xrhIM/AhCKULzHIdqCeWu5
XlBaScgLKm5qj8W8zPdcCsbQSmFWqAtpHqTyhRk0bJkxMHR2WO0V9YNFzb+G7yzYey6eFXW8oNij
rKB1eG6xGU5P2VpDEdpNlTqdZyl7d9HOCjVpiJNQzYdtoqm4y4uAXKqV7V5kLhTsfv1UzN/xVD6F
PdWWQ1DfXK+fHlBRF5LjzAxU+JLf87fdzxAgUe2Zt9zB9pMw9gBKM4gCtW1XqDU6yzXWRkFaa1Qe
i/0H/NaZdz1I1ViANo542c6+qmmHv0IRsq56DuEQRCFXdpSwokpmMt+3LpFLW3y1diu3nIIlQXiu
kKoxTjUWKZMWGlzH4oeuYuRuA/ZYJSFwby/2Ucxhxh2FHTMTvDqaWhxaZ2Fv4p1KXNJ50iYW7Opr
83AhdYZRmVaBx5qggUR4PU1766qf2p45IwE6b+u+zkfBUCMyfL0Em3xmM7tbi9OHMzMng3fidWWW
/X1udJyqLuCOL5Ha4wkgyPcwk8g02KGCGR6CFzjTTuRYNietCMZlg2HUMuhp6ZrzaLo9MSJiiAla
jri4re0h9fGfFDqdsvLHPx5o6IVeETdGP8xbUoIv8NcC95fBbIHNSudDmhn+cJ6/8ykjd4+z48GJ
zLQAbgYkDZb1ExtuixCDgg5uTJA6iZ4b1qLyY+i43TQXhZuI6O8ruOoIZ8sbe5aifUX1Ym79wMgP
cFEuYn7LXCCOKOwKxOJEvJ2T9+WFUpeWODzmmH8i27Hrl79jipfH1RyTi2oVtTepCYcm39uqjarh
StN9v7lwF+nxtrHdtWDf8Ib8yTfwAfrS29HeOlcHkP7o3FQ+yd+LeP6pAAxP9cgnezqSp0LkIEKV
/pnA5kbcqqYMIkW9orLPnGrSM/zuiIbB5ORtjgQ9C4rOHp7ZN0O4XNnI/CyJLXOaLqkr7jtgpu/z
+TZ89NxFmDtbnSmPZ+hTPfTK2GTbxtrBO0g4oWasG6ZtAWUWh/GXBwdfJ/cIiBa9ky5P366eC+6K
cxPuHPOr10nooWY1m6pZguOXXNS8ddCdaNJPwR/DTn3TPDnCKkbzbYyeoEXXmvIvw3IRSzPQFT/j
9FjLlW2nI/xkkJ3S3EEX5ARKAZtL/X5aZBQyfy2FMzlLBV6q9/lK4gy+MLz+pEvXaUHV5rso2agN
WSJaSrqBaxtNvZ8KGbMBXEOGWVsf7cxDqfY9opU6rZSsBekQEA4PS4nISVUi7AzTSqdCVYM0X7bL
J6PiZ1C4J5W34AybaAk/Vw1acLFVjc8gxpwxqmNNbvDsWl+AMPZ6pQzhKUNAqHw8W/X/DVZTbdBX
ZQcXoSIkJPvg8lOKyPL/ipfeoo1EsCgk61Al830g3k87d2Au7BqHKuzJXWSfY8qG0s63aVV91T+J
bPlhFjDcVH4zBsXIEMBfFmU3JXZ9SDg8+xV30NmFKHRTQY7lZQB6Kg1sTuaIL2yIalNLm/0S8Qjx
Rk9YGoko5xFDxJyT77yiYMWncSfvQ5J/HNLdsLeZLHwIIRfihgAsW/DgSbZslKVuskCsV82+Dy+A
Bwr47vgn77rvSYkT4VPIkJz63qpdsBF/84sK9SUhB8yNKEamZEGSIGlWTSGLiLou77FzfMJeUzMC
b6aFbllp1kaMijiM2zWkht3dDBJPnRLh7Hot90P55ZZ7V+YY8gcc9Ves5/cvE3zvIdDjcJcjHTv3
FqBPORoQPP6wfhYp3EgfCY3wCXQ59FL1ePqOJ8rI3+bO/c0R+BjqX/FZpbffD6eZvPCSxqhtlE2J
Q81Vl7efdy5CJhqFqief+JWZQmMx3b63cowlZa32Ff3ZGxUyMkK3M467/L2vOF4hfAGvzvUyM9Hn
qfVa5mChhi7wwPIEEXIaEEXTkeizRZoH45Exe2rU1WUaZaR2H9GPKXgbVnnK7+YKRIeSUXhVPNM5
vnA0M2OHCx76ho+iow7hNZ4AY1joh7AdyyVvuJitbVldHaGZXY92Z3j5/JXuYbSUV6uMXRuTciWl
q662F+cv5+kqN4+3q7u+JTNsaGwC5PhKKt5YT3K7qO57/EJvbT7J38AJcSzInfVBJ48ha/h0gBeQ
kD0jKMrgAh/13bCz3Zae151yrPylN886Ku5SXoPF/i5cAqUKn1CwyFoOxRVvWsruwkuwSISTEhzc
zVEuNLSG7kGwzB1SbckIWp4/nRK1Yns6DuSUHLZxulu029c23JoEjXHRUQ4k350n5QiOTSNGL6HM
3jGaF4/Eh649vklE/dO0gnrycvAz+QYfzeZ9mHsSyrNkoAqW9H0WxKM4rg9v47WD9Wpd2R/Eq4kc
vTaoUUpUttDcZSs9TPi9uLhoAJLZqdWRscv4gIxojlDwlrt0jKd8e28qf+okV4+C7NkHZKUnfV+n
nHQQiK6mBjpLJ8qnE8ekRlB40DDtV+iuPzgDhJTR3Ox3DSOsSUaahu2fs7pL9WgI/pSUILfYsuuJ
s6kX1kVDecR4VnmGnISxNer5S1jGlSFFnrCgIR6pyqg/GtMmG05wEc/tQ+Nlk79SdU1GScHzhhPV
pE3UibZLGILNsRWLI+4SVST/i5WkY2gJisyyWvIXtklR7nRtcRBxC3CHqY+xrcOzkQHMnmFN9C9b
n9UrHGqO7PfTuOhF52NFHtG8T4IfXiqw+CHdKW6LGsGRPsXl5I96kRFtrH7OddwIEZiMjtmhZkZ0
qkW0vcaWmWeDrwDKRcHT3dIuLVa2NOfWy+lzFOychucInJzqDjryXeKfu6ow6XuulXF/m1K4TXb6
fUHft6sWK5DbwImeDifd8xnVraQFBh121zgHjiFTis+MWEO8de3RYL94p8GkOXGIN387PBRTYEzs
2yHFqO+RlD6ZqcbRXBilsoi4rfZVfvSQ6sQW6qMRog1nCRGGkFValqXy2ldYqeL++3PPvX/W3Srp
rTmtleXc4+OdMqAgCWytKqhWKbgW0NNhwOooO2XyVBynHgvxlKynznBGywNYxl2Gp132nnIMwY4s
N0YaobwLcM2eNKu0ZHcMQJBRknGJEEHwxI36xSgOwCldQHTUHPzvDihV32HEgq13YXWP02uQNE3H
YiE5esAr+XYGDtjOuFxg0sZWfx8lQSVwSE5m2JrbfBkpev432Yb0S15NlbfrJiallBOH4+HNfMyJ
Vt0nlaLqAwwZC3hb5h9fu6SLSEhfXD4GjSj54Btxf6yz19CFgENh3DLE3RBv5DNXGwy1mLgWAWLo
Y2mWqNSk9Hjnwsf7iqgaTWdxWZitM0hb+r/Cnrk7NoE8WaQcgz9QGlv6Q5SK+jwJ+vGla40wQxGY
ahA2QIb5vSAzp7SSeJVEDvzyxHXbG3OlrDDd70k8YZ+letonNWvRCJKLeLqtMIl03V9qpOuIllCq
W/p/mN+9xr70DoEJuflca9h0ST0uqGT2oqzvf60uXTW+GkghX/sU71N86GFtNjWacXu52HdAMT2N
y1m6jY6aJyIlIWlTHyHVdc0rvNgveAKt0Y5e3PRHrsVo2c8ouxiTNyiVH5a3OwToxROqP9SPQaz/
3xuRVb6DebH87RSdbnay33M4yVXkfyId8a+61BmWkFASxZZDYiG9G2sTX38hLEFIIkLR0u69DlIz
OfnDeTXn5uU/sgMtzSmRjLaKsjWI/AXi7tRXEUBIykezPO46LpwBOKv6f++RLi15eTRmPb9VQAYe
mPWJpPhxXWXDLgIX4YaZxV/Ki+vA6L0wU2MEqg1QuQbIi1eZx5iQGSZW9GidCcrJG8t6FnzsBDCT
l4dO38gTw+PmX8J41j1wXg33LiIM5YK3blpvYIon4QmyV1cwQgKqNLqLAMpt8E71kJixcvrKXV/m
bVhAQLb5X7CWHsv9DBIWvJ7gUZlvjZVCGZtmK4cVJZOjom8Olwnp26YnhG2JeC6xZJdjmUA+XO2r
JFpSOdioiy5EUQWN9UM+c9YKKAjeQEC762E4E1joI9LqiQx8nCS9fPvxTG5pbqJAAueDLpKwNmll
1iWQf/zpriISV6yhC+AYbhrxEh22jio6R6lmUJjvegAiNgdlxoQtzPo3FM/CgyS+rqIlRM8Rq6X0
2tJvdHF9yxkeRLgUmlVLgpLkXj4TLqn3PBPAxjlazdT5FRSmbSKEKcsOlgOKPlN7/PljyWt7zTW0
BTbtluYlpZbYw07p0u8mvC9f3YeMUoVogg8XYuLwgPOK0dQ7Bc4M6KLqkC0Kzpc1tcqpgiLabpLV
sW0wIXG1S83lk+H8sofDDR5c5RCsiFZnukOS0Ni8bD7ZPylek+28YcAjeMzSeaOHgI1oIYbsOdQT
SljBdtmMoNN4zZqE66S9A/I4LeUfp39RfzNNgXoSLyYLAVAVaO+isH2u3ZK15npAsjbd2VnQhvfA
ZFWUWBWa8E6VQN7rXNfI75I03gguqJk5qC3jJ/+T6AVLYTaIO72k0oei0273Dqh6+GTj0CtIvfEq
okYNV+LBgek+3CKLU8xpTHz3yV2SzKShwXCZrKUcLdolRz+pE3erNmaZiX1OZ2X/kBH40x91wsRp
UQgdjG4Slg1ACujGVGGCvl9i1tUQsZzxwLehNSOwOuIRyZ6aXZyMIeRqAtLzu4ZVy2EnpenSWXhI
575RA/kkwIdbvWAmeerZAVL0Yc1Coxa09eJHvh8Oh4xUUuwf+AHxf7FepsVwNstIz2kOpCxauafw
BIsV7muzc9f9i8krjac7/9osVhQgwJ/RbwlnuFIy6AXLp4BIb3NuZEETrb9kLPsL6Noao6y+CQVR
QSetNdmwMM0GZZrMV373NcWIjBg0IPDZw44cS3uiKuQpaDOB1Rdqm78+L+/EWKgI63fmuBCDkOTm
WfdFFifEjW9HpRN4Xe01ZcfVHBUEM0CZaNfpHJviVNaRcMOHg6XM1hTpmLgBeRdWHP0hx2hU7r/S
qo1m4o147BGzpgsRB0S31o3GnG4kMRZpIfwc+/Eys+mJ/46PnDVpLUSfjmAxXBV1MO0xhx9S7f/2
lNnhYC6qFPpAAvK3wiZgZOh0eoYqHuNyw+uAhhgnQNPpcdFMhHJtpXHYw21GNUc8yAcMHNawxARx
9OBT4mOYky4j2kemLUkYFEUMFE2qvcllcPAtBISdstn4kwqodgT4bPGL5CWHeZFUqyqsM4vVq34h
upCL4J633uYHWgNUbFNyx8Jg5Mjf4BMjCzzV46UUA7UA1I7F/YbxvrGMAzx1lSOMJLNm1zW9jC4W
0QUNVGTUU9mpB7uxq2QGgAGreA76kKn2SZtS5MlcSV44CNFC1V1LC+Kw1QQra8ecd3XIiNJScHuE
vMMkiwSW1Ke+sooDlBISIlsWv/hzNl7TCyMVUKgKiwjjtbFoZFDpHJyW1KRgskeExw51Y9VLpjdC
SoJmlM5ySUi175utDdl1Qve5xVLi2l8RJoSh41l5zp03iFllsZygOrgglJDUfW0IljHXRJeJnF+6
9nvN43d2ZDUjg4J9k8r2ztf9GjoYzXAu3wVROQEyjLb6Du5CnG5MnvfpFzLOY0wScyiQJb/P/ppP
5mC3pbbinx6FgIPOkiQwMuFKGY/TWjbIBqP+qVRj0P6X2vB/Np8pia72Lg7P+w+T75CQ4WPLDav+
2e7i5D9MPMGkkM7uIdvluT72b8CWdJEj5StmMmwJ5PTGK2sDpIBMmht3qaS/h7ZHdOVrHdCHNg+K
VxrL49Rx8OxlnDfn9UYsikdfjbQ/H+sslNxg1gAISNBxUEbbuXTRWGI9zc0SkQGQvckhuYBWN27Y
6SKnD5hopLbD8TIiNMCDjCwUA+GnO1i6uXjdM5ztAhSsvCP5Ql7kmrq8gbhikjri9ZiTcicK6A+5
UsaRe68TE/0yoAZ5doSJo5qWz8OFua3Oxx/0riFRy03WkBu2zS+jfeR2BjpUtyL7H1hzdS7/93UD
SoEouWnRn+XS1CzzJRXxep7r/ay7bJUdOG17dQhIIr1IbTyJpxbwzO5WeMc1leZsrfkjBPp/w2Xr
tKVexkowdMAj9omigBUZyDL5xK15WqPx3oMfyxV8BqBbYOkddDvC0iJX6Us8bFbcz6IYaXetvkVH
/GzMYmQ+rxq3Thul7NJ+NENuF9ohhgo4F72NbgF6p1rsQFIDmZS3GpcTOV4RePa8TwPPJy/CrLRx
VinGH5qBZDXHgAuyFXy7QFRWi5J0jUHr7NdgenJzFF+7ZoxoceSj/GXZ42svjuE/BtKigzHxPQ+g
xXh1SAGU1QaeuQfmoO3MY4QWOJfgJyrNUyhdG60iH8El+/ZwuioKGn62rlwwPHI1BPMFCUv3ChYc
GbosltFBKBJZQf4/f6mWCoQXQlDzL6SL+BB22p2KgtNqmv9O8Te5I0dzPXYDPwLlarFZEwUNquZ9
Vb/zq/sPRFh+XbO15gV4w8IJX8IbzQpLY621AeOxF2BH9VgAzEndPS3u4dEvNMPqFTTNCF7Ek6/i
jLQV3UBhpj5+GUaBVT7vwS72Ohax9aLdsa42C9L84Mhw7fr4yEc5bxhXiMqQmaKOXrbuG8XGBu8J
l+XUPX2a0gJLXXhVc6BHO6cQilf4CDTOSr5MllloGz8zmhtrFblrQyAPbRooeDoiCZhs0Ht+exG8
ZxJIVNocEndTlen4tBE/FhDUN4sSdTXbu5eXThNq3kQy5EgcLSP7XBnrfCBWdErg5gAuYVkMs2k/
vKwa3gR8UW+WVYNLuWB7MvM9Jt00QWj1HyvLImI5PBGyASp77bu+J7nVDvyz5/zqszJsJYEAwq8Y
OFSJntu2qvPCTW8MXRHkfMy98DarUCvMxhob+3EXmruJWfPB2Y6Y4gh4kX8JL4I4e1rITqAPgYQH
8yXK+8X5NB1v0jcTXt8ZQHjfyfZgx3Y89EBt3ppBwDc71GzuSonoJn7CxIa+yOdXhu343Lkst4JH
I51YIuY7C/uwpp3DCdb5jW1MWQ==
`pragma protect end_protected

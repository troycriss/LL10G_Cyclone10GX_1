`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
IFwKtuaYUjL3A03OlwM9lhHpovAey+5POjgsKOffV5drD3V1AAp1Ih9M9LYyzTaI
ucU6cr7Fnje+vrEQjqhyIw+mugD3zLKOSnTpaOCum8HjGkeJ1irMLC64luj1XIBO
HgGpULR/5k+207Gxb+Ap8lCxEbg1J5V4QPS1gBHrup4=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 59664), data_block
BLIiLwdPYhC1t3G+y/aUOj5gaBu+4e1UBlV14PwIZdrVNcoDQM2P61iDYfKER2Q+
182N4LzUTRCcG5nkFZDdgfZ/4hiMEKN9ssvgTrGtEuIrfqbuawu9PXj3IHPQo23M
/f7GCuP0xXYKXzj21cbuPlryDl/dOwCIk51dwjKfBEBj7vYoXBhj9hGzKKSoZWcK
VP6+/ab40uwipKmTjgDnpuMdw1m7arAshAp4eSnvyFTlYrYhT6x/yyvB1hxogQ/R
lfKphEpx8Fo36bgyLo071MH44TKAxl9HRAYaIV0jFL8jVUvni+IeweSTecjf5AVW
VABshxQ5QXxS0xfGuG7DhheRwPNMEXcc7jDFkPOanU+rdYQPH+/Iqtlnl6hlgGNO
91lQ2CuVTVTcPBoOZuUVYnpb5eUE7EIg4N2/QEFGZRL/9wOINBSbVqDMGPxYajqI
j3BGgCxGKwaPP/14Bf4NQKQIOkFyumryE030/9FBuum1Kf7kL3rnpd4SpKcMORLl
Xfr4eWoHR9LxqnU2Qmo9UPzRsJVP3XOUB0eR2b6aRCKNoW1mrtnqS6MRjXZBmzsY
1cmcW+6KR9ghFVxG94pFo+MzYXeQZ0UD2a20va1KABLRxNyJ70DliZAN0WwnpIHZ
LDLZ9lK5lfa8Xa152ye3NPue4hSrF9xZpGpGW4vbiL5o9vSabssMek3X1jqG0vgL
C9iHzcyBaP6wbpx1ohYuYrAIDBRnKz9C3+GKJg4GEU7tKdkZd8zJ/kCjiL4Jn65S
4uO7fcoSUO72S2FIns0iWea1wMymVp5E3+Hs/SqgJ6u+5nRSag6U6wjSsRvZPtzG
YGx8EwM5chspZH42yBwlxs6k3Aake7XHynFRJH4tuQVIxgaVDTEpho4RHcljYAZH
zilcC1mC7I8htHjj6EfkkCvPhMjjjFX9Y5J9TBrjtc+rhkmyW2R9AdixLJmXZmSq
V7qd2szONJV8sj1DqW3LH/NRwx4+0JQRu6aHYuFAAyn0EwmPDzFblMOjFwYI1J7x
UEpy0rAu2XBMW6K2RsnV3TFT8aUufBFeB1QHwVGvdSvCV0jlbvtj1yWn7Y3BJ/vr
mS4uIHnqPFWFJrGYoTl9svyFr/zSBuTWZ9aBlgyn9S5e2QyxNO8RbJIaqR8E6jK3
8a1Q/fUjjPAsaX6h2b33CbxZ9gxQs8WFWMkPeoh1Ah+vFmZFfQht/8AJZ4xSel4u
lfB1S8w99LP9I0vncemQ7pFklkQE4rLKcOM0UyLaQsJ7NO2hcqA6j3aviJe0f+Xw
+VgYKW2TWo0ymH1bclEPNgF4cnG/pptWW7snsBf/hxiFgJ5kIQtSOf1fRWOiY6ZE
tV5M0UBei73ncYmfqN7veAcqrql2fLPNqwVktfJGFAMQTtBLKRGtvO1AUBftCDS9
HZsV/2HC3DnhC+InJLg6PGyInJIvD74bsHXgLDEyB1pxY6QcfpDJydF8iRMFO9KG
SkY8nz4iCkeQgaKyLefWla40wZrYNGtQcCDEhjNWr3l3LLuvlEALA5V6SwzsaeQn
zYtMvCWKDBkgKqtdLzgNpXALpyRAWDc5iOPf3Kt5OHqzYCZ3t2/DfE4VBME9Q3UC
bvYJuX5TrtDiTClrAwCzEO6vBSsl7W9c3Rstfxkmf/KSWMkBktdHCcD/MQjflI85
wqpbLXiIdtaDavrFcRK4DQRiMoL6hC5CXBiugTE9s0EuTZRwT7V1BGDVQ4iCAcZI
NJjaH7bl2eCxoE/KQ4hI9WIzuRMfFHNhnHnpk8HMOqfL+icUYc4ecb/BI7jdyQ95
h6qLM41ZLVCgwwg+xiMZ7RHwG3RL3H5mT1lDQMWTklUC8TtjQ47/vwQ4IKjad9M9
Fff/AjmA7qT0daJkUnQ/ci9WP2hL38B9rOP1fz+IW+MoKblNjyf2/rMZOvWRMJTZ
UhzabtiWk/ZGupMG7tB8r6OLvh/b3YvjWB1IwobuXmpo3b4b7w7YLNH2TISzkmuf
AkP7kZwrW2tfBLWXW+SIcVsGA6NG6R1IcXC9bQXh87OqMb5UpMrJflBTzMwZqCcI
+h3Zy1C3uemmenpjSHmQYaLSqY1WFj9+v6BlgFkhMaYVUzX4t+QY3S+yQw/hz0am
/PABJbMf/TNj1bQFX7SKy4EVkj8/zIXUYGDIwpjDtEWGyLV5yUkESFEtCjebFqht
gjNMKalVz0VGAyEd08hWC68xa/Kf1NSzZyeFYWGbJgIJJ07RgS0l3dHRbxb0LsWs
QqApn392rb6U3Db6ck4Dvf3Bd3B36IriagrIScJTH+Mk50Ww2RCAyz391CEpndIK
SoWNzWRMEPwaD5qcgR88E7m4zmvEdJa3niPLiq1fgxMhaDostt32vXZLMQ9C7NzV
25mCFCO7gFh2V/pbFGrsXraOEOXBkHCiMMH1Bd8SOPxMRzwkLipDf0CwnqrpxJPg
1i/9yCFnLCEwjTk7GGSi9x8q4iYK2kXC3MouANQ+F2Gz4G8dM+eGr+b9CNVPWWaI
zNqyxhoflUF4nqJdX3jC5aTV/KGwDz7z6oaukrSxeCqZdkkWOJX6kCj7NsNOmhgn
4cvVUvemIuPg93qo49eQ5QqP2A8spo5fP+OVnIfsfuWve7+qtxo1jx5ZIuR+FEKf
e7nEyA5KYD0OcSDEG4fcQwXookuViYTFWWg64gL1gMGL74frsiAlTt7XHdyiqDvt
GpOYULdVkie6BIrR7Sbol3y0CK4zxj1ridHuzjfJis563rC6gdTflLsYDXpHZzGh
LuMVpkt3I7qTHtH4Ih+ScCEg3n96wWUZ9rb/fGcQjio+GF50fsMck8wX7JxNJ9IY
jflxuVcrwJQmBE5SGG6R0PkRTV+oojRftXMW/UR74BW7wp6xgdZYuJ/YZN4WnoFr
ZknmTMPAN80F9AVE4NGAOrPitzvrZSlYszHyN/aDMqEngMtJYjrs1WWX+D+Tg6/9
YWsAUcEwAotjh8MMC/BLe6awW8+fw+PL7RXkY1I1Itcwo2mcGx+sC97QIOUbVh5A
59d0PVCMtKUk8RIbRgCipAcaFYFMQzDGJB6aV2rw3jEAcpgaurY20Qee06JigHYX
+W1cB3M3MonRKthiZDKjUTgAxs32HRZu9S0I3JkiFl4SArcmEqeFfBBNfF1k6QXo
cZxDfhqJSuVOahcbHLoMP2asaiCCdjcOcx0HxkLqefkfa+nH2dZUzBIrGVETVqbY
oWeMNLElE+xtf62m0qqqigylmEVb/0js71Q8d55e8SJydbU7IvpRD7A7ma5Kpbi0
0qe5NBK+yQDkx2vZWOtxu5rxCM4XVKpUtX8dhjovqrfBt/BuOFw9hpRse8sxxYho
NFBlndrTJN+PRZ91SFlqP1/1coHc2EOyBbrDoT8iGwqUxJbaGZ32lEusEcaxVA35
pCLk67x1OseCPkAchihsQWgAfH8YLmRT5K/HQA8yuIISGOUfTK6SvtGth6Hw3BvD
Y8CBYjB+g3xIyGzOGxYZ57UhDMYDPYdO3lruFl3wP4y67pTfzTsTZ3xlLJQtrUD1
WR23dxuaDT9YRk5gg1+Z9LtuvX/ajnfNZBIAl8tem6EPBnYMW1hIKTFD0vjy3Lbi
fNTIMSqGm9R7YLgpnHyrTPAZ/Q2latDte5p3xelfJgU4u0zrMomQbh+h037CjC4l
qpLZN//5MVSIHPNRUQzPxPF0c+UZK09q+3fY3Euafv2F9woA7ugvK9FeYuizZmug
P0PUGJNAVACuySmenE8pusPjd3HD0nBrXYwrZouZkSKr1IAEeSgb/y8yzRDRWi9I
smiC4HcsvpHx7BUb0FiaT7w3wXrTHvjW5iAGuZSBJRoWb0UGWjPraBY1lnQASU+f
XPA54yrhk506il0x6hOGKhCSykSoOBcuZ1Qut9ISI79h/ztF2CWuRlOx51POHk1x
V+uXNc92rXfrNf8nm7owoCM+vPINjGU+sls/tRfe02Z9t59vVfY9fBPxBQOU+D1n
RCDDngh40vYhIcs1bjMLYVNYAkgg2r7mJX2y7hu2OMLykktNoCkuZhq+OL6ohCqW
ptGx+DdEYy8DLI6uJ4PMjyMyg3fVBUePXcCZ6nbSLlyNsqkV04N4IySadHiuJImL
6l3yNahmZxg1aR26d6amZjr94OFwbYyMi7rSQ5PlgHPXqhAto9JPBlcmW4jEbrlL
07KQ+YY92AB41B7QEmFdfyTTjzJ6nER1/0SEiVphoCuYZ8SRL7PBTh+LaZ4Ujgjj
dySt/GIsxDckejuvFldJPkxnsSb949O2ldkCwkJVfTIPpeSifNG6OKCCh4StEI+/
nOVM6RBiCD5XYCd5UtisB/QKuEVJf6bU3CGYJRzTfd27JOXvUDt71JLP5Y2bijyp
Oazcmld+RTG349fsEhz/qshqjgRvUwfN0/tnt5f/7LWhtwwrrFYYqzkRzUUVwhfH
bxDeh03Sxf0MqwAEKqvvMEtoZXmYxoBBIpG0UKVXA1S21D5EfHWOPIKUxO0tBGUN
QiEjEkHAdMHUNxuSxJUoD3GSJvkxRH1T2A6LvdquzDYUmfKIXRdYhzA2QLO9Ya4c
KvSAEzRGnMTEab941jNmnJaUjex1PApZEhspL4kwO85aS89zmuUA0d5w5q5ZmRkQ
KNktvfLj984vn1Fz11+UliNHOmXrcWs4c2rtvgAeSfWfeUikKZgleAX/BgCqEkaf
4htd2s5KjY3iDej+PsRCc62uq4xQJjJSmcDAXy6napA2ntPHhLXybGPl6IM9/c0A
7Gsn2ffg38/cuXcGRe2qkWkBOQp44WE047Vi/MyGWbjsOo57Nul63rlSgecllIOs
ud7W3MeiR0BlQ5u0dNvTYUeE4e19+dOzSPmH4YAfj8OvSMmA9l03GgeCJPWiuFfH
3YXm3WXymQ/f3bu7W0mdKDyTMVRgnfyOLKRJMi4tZopIzOW/563X/76MY2mXuaSQ
cfjHnmej8fw+Ho7q7CTCTU1bMh8wAlgQO3umnS9/mq7N7CELVvPB8gn5chM0IYUQ
6AmlhaZ8R/kD6wl+KpJ2lAh76TKD7t99+rht81qKCAS1Ssy1OsznYi4P2yii9d9g
Y/dRHx49CY4M+gghbXaEYybZynS5psUQuAWi/omOEDNhrifgGleyjh5dljm7cZc4
yq4cZameDEb7TgFpXZ1Ep/CfZiJKqiLzrziWW5CnDrhkloM9VNvG5YIy/WpyFL/H
Kt17XSCR0amnw3bCB/eYjoBFwC5kGg6N/xFpMc4WSupzEprWpgDQyDtrVaa7DdWC
ilxjefEEf0LB6wexH7MvJrWjV/51ciGXVNlw8K77Ozhf1C9I1XQwPQmTXKzlfOBB
YNhZ436SpbnYB50KJU4JpZHhWKRtHrFiJvB8ihtGXHuTSswI4ivIGNiv3hEgv4bp
o+uOeGkNWskcdqLZgdhHFKrTl4X/wYmn9urNL07qkWwQqb7rX77+WlNLvpBpYeY6
iHmnYBK5D1v5nb8dYIVlopaAoucZupFjvBiOMxSla3Y28tOBK95frBsfJUOibBSp
Zb4uzjZr0lzhGTEw5BQx9ZH4pNgxriE8P0U2bwE3RK3faSXC3UiA5mFzuncJRdts
sndfuINUjnt7J7mjLIurYWIdAKWGJcM61NLDLVB/VZd/8J2J2nrv48dMOVU1UFHH
I542W3JExdESMH2/AnDhnEhrPE5iQKXIMYZvJOdURCo+1wgP230CR9EFzW11D1uU
5svivchImg7ZULbRF+9Mwvn/C1wfH4+kFaQY7wQqmxpO3P1MuVwiNk5L1WC4t/Zb
ahdCBn1zr9O6Mosj/nWtZ44fXVe/6AsT/1x/BsaFZumL2NliZ4FbTfyyARqwm51r
7MfkMuGA8G+KgVAlSm4iKSutR85miyRnugPptoesuKZgkuCbBZcK8wjpG7FFrPb6
1JwliITVmrkYPpY46TOX4f+5cXNITE8GJv+gyemz5k4IpF1//XTAkWLBBZfPxuBz
zxmZLXrpaSRP5nwU8IdRt80rHHoRbTjucX/YmUqjHpe/oxPQc3ywDpbY9tizdOCf
LEkYdtihYOnyON4acLJ7mr+aRn3Hmh7JcZIzYePcG3qMP85JThAD23BDux9qHMZD
NduUQpr2GR9n8Z0UhU6iHc51d6serWdEvQteQhW9vjVzOAM8RzVJSXcT5wmNGxZy
p8TkSCNk2iQ1jQLcZMzJaw59mbTiqO+kiFWvLhFfCq1ugXHC5cNk+oMbT0bmaP2H
JVZ8J5b676d7NJWHpROWbBkdeeQFcQ22No+hvhqqMfD2qOUG9WjtA/bQyEFpJczp
M5VKOcfeES60cYGxDhg/Jby4QrMH0tkVVBk+hysDxgehdddLn62A8Otz1piou/yK
6BLXgN/xVaHJp61JlpsX/B5DJ6WbFD2Acaluaxt9TrKZyZb1bpAQHoEui4ze6cHY
HqIlRDxb/pByFgcrUC9NcyZGmBJ5tJVePeV08z+2/WOJfi50zXx9IiKaVsOc8y8N
cB7wh8B/2fR/u5sdDfw2NGHx6B3JIU1hUAQ4cKicbu+BhfXI2wJTjmj6YDvYAOlB
7uX1Wba4kQOrolZGL/V1rR+/j0FSOvG+3zpYk9U0+cV2TP9Xe63yEwzIxJ4R3J7w
8hJR545xiLEahooH00v4hALJRdYn/QnG+EWGFFxUGszwUstfwnL34HNGgg171S+X
nGVv8vtb604BAwOOYSiQvImIEk7WP9dSdMuMlfHSjnrD5yYw1yz7Ge47wv0mo1Yr
fH9ifc3py8x2UtcrUePcIWMEyabtMg+Bq1wy27eE9Cg+YskGM6XxzTXTn3JXJ2ZP
TMHtFEwM93kljvhnAqFwBLvAjHMg0w1BPWDJO9e9rUUzj1EpoRbV/q0PlxYuTof/
zBoeuVhXggZTNtrGKIHmsNc5o+keb0eojoor60UdphEkDgJ7IrZth9aEYT8zZxIS
3DRaqnAu540ZEbm+4BnNZ3UB38931ux4+dnnoyxHSZFI/K0vJ//2Zok/PuI+Ich+
31lJn+3q/Myf2bbe+KM9OQ/Tq1raC79DkNzQrar5B0GwRk+6URst6NIwFDMjrdtT
RsFkX2dbPw/zdMIufBiO6fIn8IUc9FfDs/RSB0soVp8XozVpop2ELgj+kX/b4yZ5
GqvD6yursVSeyOOCsiRXiFtSOTw8t+Qc3mrVLZf5BBxd39lZiUiokigXN7DAxMUQ
2PI3liQkMUOOXJhfCCAbZrKe54J5Y/5JLZymE5pIuqTyBxyflaxnJMS+0VbGAUX4
7FOcEi/O/liE3N585cTzjDdNsPFqc3UvqwVdqXUTi6JgYwZ3e8Elye5d9oDiwihp
y2C4OM0tAVBwp2zNyK3J6iyk1Kgf8N4XStz25HyNMNYDBN8VRRiivsBUFo1qa2BM
gNLPPFwaxQQv7jm3zbzVZl45+g4QObA6mKf9q0Hzt6lw3t0FPzZXXPSCsIJOfOQT
rthOXeSEAhLv9LeNpUsQOcoo4PxX/4dWWMSkorWOR23HsRTxjJgMBVVCC52lcKJB
tvQ4gvNT19uh80JdJogNuY/6kEhdcWSjNVgTJIIENvzfsDn7SnHFyOnkb+zXsggm
J4q4o6wcKOwc1tEk7JaVGeH7heA8CSmFnOc8zVqVPfG4Lav/qc21d4k/klqHgoZV
1u/m+sff4Sx1E16O5ho6Cc01dc8xPYW3Grog8cIFD0RrGaU/x3IFvon3T/HEbsF9
9L/VC+M/DOxRuYGzRn2l09F1bE8pNrVWTSYuTOkNmOZXlcEWLFyLsVbMOilMOfhR
iMKAlHg7ufV9VxtZN2u9HgVvq6iZQnoW4okX6pME0wH6xV1yNpA/PY5MzzoJRYC9
Xw8gE3CjJ38fqxUoNAPq+lFSvdCG9VmOz3RfOULkKiehQTD3pO9u8doBsIl7sFgM
mIOoMCT5gbZ1O+VNLuPQz2n0HlsP2l7DABgFNtF/JYFmswkpd5J8EeQiqzA85oy/
nBJLXwnEYn+JB9FiVBIONxdOK0HvfMS88GjQGucJdOOsuzYuOOmnOFGterx+Ww5Y
yycfXFbzP8xIll48fVEv3xUWH3a6kTNW/pRrieXjscMuGM2+CfT4aCIa1eRvdswX
GQwWHXL8fsklaqJfOaJK/vyNcJMHqwQbOgawMkv4tbprxfNJo/FnrEmy/6tV6fcx
RGpqy9cubB2xgaQGGFsU2M5Un4YSojukg/hhaMCLBVB6orM7uWJhGpwYWFqhn6cs
G5kF5kio4bTGZ7qguzzmL50hvcoo7yYFUPpJPNC6ag8fPW+3y6r28Vh/Y2xg1Z85
vl/bURCUUHSKX/8DJP4oVdxz6LGT5E5QSVnvgLDG2mh/Ra6UYXl6ZlNoZRWBlBwH
TEPV53tuyguJFlUsv5kC+YYL3u31cUGS25qV4qu5f82M/y+w9wd7AbeYXodmAmU3
Gue+8Gbpu27xhvMY7qdV3QtLkl3UPqJfr/dhhbCGTKf2+DIdFQ8BXvoAw9JlZlfQ
9xAsNralj0fvsu/fg53IMqkBQP2QaOrqPb2HCb+GTOsH0+Xw+KQ2ytMYmmfXFeuR
w+pBBqMrBAc2oKZpKtbvzmuz56dbpdEU4qHyrTZKDCpF80jnSzzv+KqtFCMQB8qn
P0evy5rFzOoaQWWXlqUVAdhZsYtNRfqgx5OYuMxRc8SL8pK+MrhIBLLB+dN2g4tQ
lfTXdmR1yTTjmzATQophs6QKaphJzt0qPxSDfb0aV2JnXi1Uu1+K9Js+G5YlphaA
Z6VyA8Sur86j+q8kJWeZzDBDKM/IDk9mBYvwjZPU06r6usN41zAorNWFtjuInc9Z
ejU0FjnDvm7RSWtqdIcbcXjWiy59di0MDPYHAGEQho185e/m+vMegsJBqIbDgm9N
YT4q2o71yCYSEZH2cIT3/5Hsc6I/OJ867mdqhKSBqymJMehNTmOs4qk3k1hDnbOx
MCBbFPenYngw3M7RHbmXfq7i8m2mv7xheUmx/kuV95gzZmkFwxVMy2tN4Z5hr5AA
uOgQHV+91nG53WMxtcqiqu8Xmy1LQc7ehmmb3hE6jzu6xxMOmY0Kr5IyLde3mTil
W4l24UnqLhpoT6Zxd8FtU65sS6+GrwnZ9ep2xP8rX8oufcqGj1r7p8GAb6hV4N8X
kRbNu7tr08225gG9ZMF+kDnGj3wXRJVGiWqa0tQ8MgZ2nxcHdEpujX8m/dBlnHhg
eHDktEWpkkXtOPxBLR+tVoS3DowXI33qJOsN9PUt0Gm9cdur79omlnoJ2+tpYr1I
/l9rYQ1T1zBRXyQ6mAn3N2K69TeKxLfopxzlGI1gUuk3ueL2gnVdFIq8Jk0u/ZYX
7zu99+GmfcNck/Vlm+NznXHhMORD77ShqAbtyaF2wGgj5Y20FZC48zjhPJ7szJ7Q
0uAI1nqw+2DKL3goOeDVNYrW+9QBNemTHJVvddOwd9fmW59unGIk5ODWnC7wKSJy
yaQ4Hx3vgYqpp+3mFv4yzOZKAc3+Id+ybV0rreidRfnPwGadWyObJAX93SCttGEw
MHeta5BYzDIe5PyQmFbo3EVLbswd1D2NaQBAlg8LDhmIJXOKRcPW4gnYC3MQFSub
DZ+1jkPs/Ro7ForoVuXwPeKuXBZ5AuOhS0rv7qHjmyymc6eSjMk1lnrZwgp4VdRr
+HydOrNxROTuZE8UdYOIidJMkc6f8qNGQyKcmRyw/UIaXj+YUgu/5K3j6VjOq5Nb
5DXm6fIprUjRqpPQjkEpsPOUTjE5DC4muSutHoNokGQJRBh8a8aMmy5wQFl55SFX
UyjM6zatB5N+oDarLrHldEmikkJX8SPhTUEpeF7QxCnXbAaVOi0sXFfLbVLnVksn
OcD3ane0H9NXAqtjN/v368riylj4xKlKLxeJU40ZQztzj6kIfLXfmDq9q1WfVzjM
iZ7ZZKEzdlc2EuP7xrSo01Ym19dQB/jGuEIoEsdZCvDcBhANDunKt4AyvG2YOq8Q
kGb/gs5MRAQdBEnyIdPIswIJGcbgPCCNenz6sMJAZgq1Ws4lmWbnj2hxug4ThMzY
PQMCWPGIHMu2zW0lLAxobWXb6JQ2gKJ0UPdzY3dypUHieh2S3DE2L1YA4LUVEwtq
T5UA1ioLznqXrmtXhJZo9JoJyCpoCYtcO3qP5aG2vWnMlEEqnTAW8g1Czua1Sbkl
tk2nrh63+KD77mx8Ej/u5J7QKDqXDXAR/aqMADMDagbghrw3nz5TixTiHnUrZIES
r7WhKut/+gzjGpMT/uXpQx+oDUJCHmeQqpjoUHmQCfzF181hrvlpJW+2094ZoZ6B
Soy/8c5EcBIXXAEjWgcVym59VfOeLaQysPEOTFLRd/4N938nirsgW3YN5dXzAdW3
34C3mdQL8lQlka4VkDoq0E5suHxN3OcTt0qSJRmvdVxQhgSgtUoroc6DN4Cwf2GZ
IVajtmthSxO7dzQe2B+YaQZWJLMvD6qrrlSRFUv236wM8m8e8rqTyk0wziebE26P
eFaEDoOZp/rTNn2LS/60VmA1mo2cs0Eu/8gOn5MVBaCbx66O1p/GdNr3y4z7cWd4
B//pgqQKnpzqnDNjfvYnbdm0yR8gNiEm017WPX7vNFMwNpf8sY9QYwy0V7OTSL3M
mRzb6I37tRU7CWlAPWaBoZIMvxiHK9mTv6LAJXCKltDdh5sLkkk2UQIfRHwNwqhZ
r+o83tMFCDzjjgx2BN5HBinYUFDblD/w6eZY//LR28aRz+Ntosc5g7Xps39gfFEq
rmx1wNKb0lV7UshibepMFbokx6sjk0MKuGy5ryb+zbhadPpPN7tu0sDhAe6FRI7p
G/5v91Fk7mQm3/GZjlL2AUU880QhGcaqWFcq5NXwxBKlsYChMi2guHc72vwccMu1
FTscLHpN2CSOFZHlsMh3QaeyGkpw4JA/rgBGiVZDE02JgA6vdjutJeq+pdjvm0Mq
O3xHCJ4FaZRmptUUkNwfnltoCCRIMiQrftlXr+4FYgeP66PBOHQyAOeepqvevDGD
sS27rypBBhteQNtrueLtV5n4q7qR6DrZrKOdeh6itQfWuApEXhF8YDp0pT3/jXss
z0bm9XX1HfE5x1yGvM1pwYwFrtJZJoPWobXkO4KU1TL8Z16rmWQDwRt3rusMQva/
HztAuhqIv+1J8F0QH8PZn2Yqjulrq2PELv8DUqUzz3wUEpc65wOknleGVeVDCEZr
DUY9y46t/SqTyc7vqkEC72M7JyPEPo/ecDIIxaNJgMCg7L2aO+zS/xZLtza/5wc8
IMzEaBnBAvZF3zJmfddp1NsNE+DAmg/1JW8GiN8ptsiIUT8SRPRkg4BwMTuH9yMW
yvmRyWbWluBUoCDfUNL9kdJDkubXYS2ObtyOxSp++uXIFM1zwG+wFPmUWQUEKNiD
WaePvCGMkgxlTDP0BUTM/p+OW43wIbp4RmA4g1OEPfF4RXY76Tq9ecYBXJOFPORV
A1s++D4CXweAb12k5f9pokZK5TX11oXb5ja3XvLyknQTBTskxR9wH5y05iQRa5ie
AOziJbzOw2iHUbR9g1DuwBRsQklQH4n0KIKGSj+eWz0yTGED5NKh71OW3nIt4jNg
8CY3D/iV+9m7cePgF5blqiWcJb0ooWNauYg+PQCOST+i+vRmTRbz1ER9alLitDJ+
hk5hgcKo/EQ9/7cIxUC+duy55KmWRwZM15HSLYDe33NxWdyc3nxsQzYjK2DzP/CI
rN7hfKoVkSrBvf3kFJnN6xoNfvNbbc7zYBxabOE1xH43/qoLMnDb1L/IxTy3o+Xr
Q0X2eFOJEZ8Xc8oTUT2vD18g5IuBxnp+QGYTK9+M/dPnlsGCQte7/XwVsUqscTOm
2jpKlIQ7eGdzJmcQnQb3bIRp7TnhI5v6mCIT5ZXZNgcBTbWK00lJ67Dc7DybM/ed
UuJLxJh1xlLZKLDvrKvOX9A4ekCjFNXBS5rn/HF4qT9qy8o7Weky1hXTKn+eqhGl
Pd+djeqS0gODqt9YMjCkx84k1VHwKFQ1E0nOeTHHtws6EWYIci6qrqv0SP1U0K3e
eqGJxJVGULjvrUXaEfVjAUYsHB5FAhJoIOJLGuGcs33sHOYHUUb9JtNFtyRRG4T4
eU3+/Cpuvg4RQVEVrpl7w/z/6lYOEiKScEBzyg4VUkF5UVSmmATTDhrpi881Irgq
6ozUd67xvUKQYGIIpo+8U5VldZFH/5IdvtPRtvtn8tK/eV9Rhrfja45UdfWGV3xf
WotZzMifJy0732oIXQ+9vTqOTWMFcMRD1rOAohkc/1MKA163MbYF2TU2mws91fct
QrE7CgiSQm9HwkjW4A7toyr1AKeO96t9ATUsk7a9rcOD1kt5zQktUeBn+xc2j2Ou
QSXBHV6f1cVwMqI3ICIrMdEIPuIHrpF7sZf9nwPolMrb+gOw9+a4Wkhv8+Xf4/96
Wpk9EFeAC9k1RnsHrmjX/d9a+h6thPS8dSINTALZNbWRwv9+NWCqAA+l5CE5vSa5
LzE3a8yJmL7pDmqJIG02bwWyHzLvRomJS+ibWdxBcR7MfwoAwlk4dSbXrVHNv5My
Fvj5kjvlYM9di7CdS2Q6LomW/C5bGQ4vDJKfhRVKWt7Cd2pS768w9cNVU1F1OAHE
7XBD8iBdhtnO3syUe1uI4Sw1Etz/DCylnbMEqXACpD1eeWP4KaLmpPHQb1YfdK5b
BLuS5Wawkhlsn6x369vP2T9QVLeNFDdQ3tnvPxOSpZbflJHpJeS4J+xnfzET8kLs
BWVIecuCFmEYnycF/3acL4YV8fVqg+y3zXMyEyKC09sHkFervUK40TokSSocWC7G
E6hhzokBI+220vdJSmTb0LJfwbr6uiJkZmcdtU3yTP4d8TwID4zjhm6lqkGWnldo
ImFHmDavp0YBDSNeEBkJ2R9Vx4u8yyMqrdX7Z3PZ/FYVzERqtt5xSrFYIvt3Nrvy
/EdGJ1yw/BAFSp1Rcu8Bxwa9T+sNG1PO0iZHKzGPaJD0ZSzfxz+e6JXzsagKutus
4GeBSc3alyZliOzV4D8QsTzMpeCcmJ2RAWnSWxJilVWSjbxSQ7Lv9kU/9w1HyelG
WVt61abngQv6LMTiRpIQz3WgfDv2RMjOy9nQcLtUF6XFKe/hmad/IMF5wlj6JMvg
kjQtIaw4yTGkS/mRSi0CwMveJIjZkmH88bXKJMb4/RL43iQi9lGyuORMIpv4sEI4
P1KE5ZOYDzGkjap8naofyd7ytVUBk1M09FPlYUJHWnePKOVOruWsiDfNiS08w4fw
50Q+A7K4+mJ92InEs8HtLV50rIZJmyPt15v9O/ZLrjSUQstuxeK0zH1+2xA/l2nn
bZQhDaW0PYPVxMN9s6hi5RbOqgYOEMn3MoGFosOvZtNGGrkZOMBYSBTy3M4Ttt84
2PTwMrLE7hf/z8r4wA9Utjy5gSwOj3aRUQmJ+V75S24Th3EP118adHDeEPKy9W8t
H4xHsvJlnMzgX5RdnN38px4GF8v8G24aluBnXtH1IE3Ni5h+PIq9Be7Ax3XG7h3F
8UOeYpvptU0siFdxrqcYw/B0P5AdbqrG5Rp0/saorAxjPAHxWEirM1f43MAm9ASi
fzOx+q8x/FQlZ45ztxs2jmGI2gwaKVUvJWLRZXH9sLCXeoGvewDXmYMm3fV6BfGp
hSKIPnwqjJ1zyJ5YSTRF0wDpdBDkJucatnJndXpOWT61x8PrbdbxUwCeIotyyvl/
HENti8jG5jA1aVbXYRfWRLdM5QP42KmRyOg34jEJ2NdqiFXoS9U2b6Enc/H1aL86
ROJFSgMFQ5+cPoVCoIzUkDftGY4GDC5PpIJmEnaiFsl4y2eegWRRuFGqE3rctmQA
o2Fo4/iextDiYTPw6oCVFmlu9UIWhURFoOHTD1+K17W+dZzwoXO4DnFun+VboCBC
9jSTP06Xa2B9ID6WWHgJKd8HyP1rD6CB42Ehrl0YZAErRbQYzzFgmdR5CZUywNbS
4u2KgsZR2KShr04DCzk0djRsm7PMemJKkWiBQED37tzAizETeYpoRuhgNBFuXZHw
TPlUTnxarfoG2tgGSt8wPyu1TksepL/kcWLVK7oPqMEKD0NVNNGc1ToIMbWbsuJs
vanVhdepRYHrbOG4G/dSF7JTqclY10+DR81ERj7x7MNOodxecWtsBJktC61+TBpK
JVADSjXLkdyz3TkZPxpNFdHa3krpwaMREQxXDRRLo3IrHaaSOxMXWnI903nA0O8b
TImuZdasCdbIcD68Xy1rjfH+09cJOKeol1l5zgAF0cozsmc72PS1gE/iJsZ+fnkj
XygXEa7SBxoX6+FXZBGn4+FFljnNDKYNHHIfBKep6WgLJBHG+O4+2S9AKkxd810P
zrvplMZms412+JSCpaxNqfwZCpcZCu3q+w5Cl//42QQNFiHAOIVd8k+pMz4J0ti0
xscaP+aRsF5x0THX6AAPfZolgtqsxvUfpeh4Q2VL6mh5IukpVc9D8kVtik5B8kfQ
o3tx9hhZ4YcOb5y/UJaYsOxofZX2gka13IKj6n7bU47jP52cUIxmZ+5ckopq1b5q
XLyALEQe8L7xr9Nue9W+MApbzuHD/cEuWTPnErUIjBoLSmvLTrXnHMwYzSBmr16X
CJ7JgiDp/LeGzfY6unYlNw0ZR+r6ISsZ6ncpEIgbiJZh7Ngnq0j2WrQ1wDOcaT4V
GFMKuRsLELRuGmDHxKPNTnAyV87SF0phTTByS4wziL1aTW/lANB8fU+fKxwz/SFU
BvB8N8chLgaM0s/WLFzJUJMClFyUfx5vZ9wHPpDqjv/YHBNFpb3hFMxJnwhJXmLr
EdOrROUqVpiTrQhta26STiXoZ4fatoIk8/k3Q8eX9ImVl1KD3J2jHALEyWhJ7Km9
GwBaiQZk7z0KOl1FJArwlVbIHFijcABXgVOxjGFw88AOl2LeNlZd8ywnpvq0canG
rt7uU1w7UwE17N4+hrW4fcpa6YYAOgMj3cRkkGmH5dWFNyT9LwIiBD3oMhyOlXEt
F/Eik3a6Tm6jEUChZgp+7LFxuld4PVs68iaXzzvp3ZfBQkB3Mpwx1LGEgs4ISjij
N9b4Ub2aIHlswKfjJr5MsXvlJV5Krs4Scv7rYh6ulhatGkVghfflTkdrBJXFPx7D
kLS2nUa95eB4J3Nk4lTxpI98Qch6yPNKAnki/ZX2pnnblF8MzXDceRSbKRVb3rDf
EfRUsGf63qZ73HX2iVY0G2PM61zt55luoAUGU2h0YLfrFJUNAXtAOuhXr9VlojBq
7xeOx03dHTadMZUh2gwP1eamsH1kST7l70SD/EYvE58Earinnckp1Eo+v30WVs9a
fWJ4PxPK47CXiQZY4l1u+JvRKeHtViAm2WWwu7EBRJFnT1eUZKdfnQhreEzTUi//
/jjLJWYDV2ipvEmsI6DxiMD/haebtm1g5w1rG3WLSghUN49cdg7/2/oY/fR9kn4A
kCTQoBYAjbwhY7GVIG5FQdisU0BfZS9McGV9beMrfiWi0TACJRQgIGdAZcWxrSQ1
gLsEicJjXsqBmGtw9LflzzxaHDYbh7+I7YRa+3D79u8EJ8Nm6QRWuMpwghY8J2tc
s0fVjBfng2zP73+0NzFXe0xlneXxw4dtUnDyLux8ZMI32/kZkKnUylNZZu06cfxl
IkbbfUUdfv/Ci6hDUJB5t9zSTb7RuEBhhxwz7vIjygQWVUsIdflJAV2emFtHKkVV
U901QtVv0qHER9s/9iZioRQfhkKnwux+b86ERxfniBJVU3j/4h0eOrCkrTZ0iWR2
2PaoTsY1pI1co4xoHFp8LUdtbK7so/ep7F83uFaesxE0IpqAPyYIKs5q7pyEcTNR
98LxJCUPxDwW2+OADgfKJF8ZvMyyl+ITg5cwvr8f5oK5XhWBlR6Apl27cdxJstGQ
DSJtWs5IAJpAhvVyVJc/5DdTHMdZviIY68Cigmx4J//Ur86ZIbZ3Mx7hb+DgABaq
ruquFG29yAsgoSxnylyh57UZLWiWxAxo7OFSEb63Zmwv8885In7CF8hY9ao0p2f4
lLJogn/HPBCwKa2DofLxSd8YVBtGZINxpe5mBP7Qkd5dtsGSwvSPI1nY4BhggY4M
jwsrFtiyPH2eARaV3F1Fu9KEKBDTAu5qeGCvSnE5GVulkG2MuLkwu2pWggDalPIu
rRwp5aIoZMhwvUkZpVXUU4c7DQgq2lKYcZsEZgc1cMqpzEg6r5s1/468dkwn9RYD
qfXnuF+Pan4B9SYPeEnFLSpKlH3JkTn24V3J2qTkG/MfLObuc0vD+MS6Q9mCpE3i
ownVjOrTNsPOHGYYI4r7v/lk0sIgFrEeK/NlRtNTuKbE2KEE671CH59XD9BAOGs8
nIhaJCDmQmLotGQPparbLFG2xhdd67ogtED5/6ATBsjMprFhjKnJaU3OlSWMSwk2
s3O1vZMyhJUqPehZTfC/tN8FodPxKQv310HiSmJSNhrsqHO+YS4+ujndPe9b/bVE
ywU+FQ1pAOAemVaIdiyTPmnHVHA6ryWA3aqnEGixJ2vtNS3f0+JqE7iU4kshBbnv
Xm0K/oiyJghWOhjOkoeMF9mYuHso9sLVoe2RXvAOMns5c0gh6EHmu77xYXIBO/Z+
U2Y3vLrwWEeJJ7n++OgQU0KXQZFz6Km8ePje3RNCF8rubPyGCJwklHwutYN3g/24
Gy8uiSTU074BEVnRl8MQf3YBuFFVyc0A9E4Uie111rPSW0WoChzqPlVmiBdjoH/a
AZ2al1JUqg44sFhmFFt3Bj5CPvXNeq1MpFYmoRdPYrltTzGzcvIJ062Xlia6/urE
AMup8hWYGywHSvSCmrNRNMD2gWnUAxDkAmJ2MJvGlephETsNA9Lpyk/wdRcHjwwy
J+ily74fwrAPyTfKUVAFPHR7xFN6LktsPzGM5c4Szp/iUpVmNtxkDhK7rBpSROYM
R/ylc90V6xBtQ5Z06Ts+/GuBVF1ee6GZy78OiM89P5AyfsYcy0eV2J+b5QuD4YZr
wl2Qf1uHdEbZVLRv6cR+npeXLYI9wl1gKJJhqM5nKwb/9lj1xCyXsBbvNkSoozfR
ZiaGcckPc1VShmRn3aXw8hFlqgnaTyFFyHPxT1K5cBWx22s/6yNIn3ppdhDScjGh
wp70724FxgGElzFuQaF4sI0AAV2VrPA8cs26auI+iaoKcNl/nLXyoEyfyQQpiHZ6
YNrTL9nfxN5I4vDzfq2aqBTQK1K1UiurB5T/GErFi1ofmbf66D9iT1x5kABsNT2S
a5mKlOn7uNBkKzyT7yCqN6xQ1iPlbGEsU5S8n8qdBaRFqtUVn89eKSsQi3kPAP3F
TLYx8i7bm57Zv2mRMwDpuHjViOxHzxXacZ+R4NZKO/1LP4OCoeWP613b1gsCqj+t
mnnqDKeitxdEtxmSUPJWQeRq+Qg5ctZD2buryy1X4IvJ9oIc8hItWUTuw3Pd89Lp
lsQex19La108/dONZYgR2Xph/nu7VhzS2ZXWR4tG/MoWGHc4itnNSPBxRJ4o5mvX
HAod9A9mJzqwpfyBE7dpCUA68j3lcSAdx5WoZE4LmT9/LCrj/3bd+JGxxZANQQUH
m71OW57/yeAJpTpGljVTpSFE1PNvhym2DCpAQ2khxAwzC17Rcu/bqKtjTTzlc0np
h4dClYAIotR2aAyn6XjSkuhsM/xAoupHpWopAuPLAZGQbUWqseUk5ukczZXMRGdd
ldJs4Q+mLr+xnQBAhzZofYTF3xC6rv0i1ugUkXxUL3u5V0VZnvS1ajTA8nYrEi/5
9E5bibrTf6BoLoQwo40eBOzs2WW/kM9/vFuo3oQfFVaI/3cm0Ee8JDh9OZKgw5PA
UmTY9zp8dIAaAClkSiI9bWABdzYNh42QvPfuHYvBVWxxWEZApRut4dWQZ0Mgbqld
Of8KQTjVdSN8BqsGGuX6qANb9+2jCSxltlTX2ZDw2VBGqRyRWi2ln2AZGNeLnvll
8WlL9f/X+W/pjiRI5CFtqBQQPxX0GusKbe+U+jzM/wRSkak+lHFMY17UjcKIhlys
XLtBz0hOhGh/E51OFM/FFoLQu0I8GN2m+QvHr3DEnrQL/a6Gy+Gx4fY3LAYE/nr8
YrqQ5oCiLolGGhK8AbnnAvC7YwAS7g1loot+yLqXCHH7ISrruGJXPG5zGqPiK5lZ
T1ijVNjv2jeuaaAkoI9bRewK/evIx3HQ9ur7ZdhWy4+zf0MLbnYTZlCnPwKIb9x1
NGhn90eXILIryqaJOvajkeRnfWRcPKpQJ1lAELOU95fkLlyIJd9S3cHWLJBlO19W
6o/IBbCEjJqK5tMMBpxYMMMabrOvTfagOVqmQcux1dEXR14oCHazuEuhZ3wyKwuF
ms5tfUoTdX1piDNxMAILoyixdEV4d+C52Yn9yuGhbBOEWO4NJJocwSF87Ci7zRe5
0zaPcLDF9iq75z+U37gmAH4QQ5WiN/SGquKC7uh4IVT5ATU5TsEs1um0xpIzbQJF
/6ZXyZXN86SUV0fYtCUdGqqH0GZqBkBvFe1ZRkaB3RUzOIFUynM9XjmZePv7j1OG
mlaewKEEiOEp8R6tyYMM5XMUxficrf/BD4156E1qlUntZrbW58dnXZqlECb3BjS6
pTGrAKtb5zWW99IFIvwflazffRkxODvBdhISKDh4yaMs2TmCrLxursqJJKBKnqpe
YlqoLBdbJkQFdcZafRfPu1WZf4vBQWyQJl8djgwhtjWz4fYpMqZQdCwVg4MJURVP
rM8EALL+81b+LR1v9wAHUpzXulVT4BAtDb9LGRUnYQB67U1Oge14GrGQ643mCnTo
frrsMjAK6kX5EWKMQFiTqqqB5414D2UHooioAb5qLRNqVi4tp9EHFBLdfmiX5EL6
f6Cl0cRMdZjwNWrBbPBOFfRps01SQXcQ8F9ht5vclxEtTaDD20xW8ICOfVzYNxgT
PKi2SmnCSibz9MLB/IcGy81gLeyWjPXtQqStQAlakjR/793ka5GC6qpzUh0tQfTi
ZVUOroHFXpqU4X6SY7nHip5I4qSscJFi9lmtO9iiW7S10AyXMiO0FTHaH7aqh6Tt
nFdpY/P4IxEyssffPf8m/iKUHvXtzu8zY2XgTOTVk1nWG2JXIhOGkC7Qov+GAOf5
CiY9cDvSpbYzVx3vaOf/BYNM+xKww7iNJoi+KCVtXotbfco3DgsHJCdO0mypg+8n
Rc2ipYzuxkkrS3K/R8yEZt9pLkLGQZZVz5RlmCE/ajzlBV7+aVDaV5u7/qjy4dSE
po7uTjDqMUWcTu75FbcD8o2FzWtaZJKgEw95/p07K0IIwaO7spYQB6CdQkCed3f4
udvAsnusZdqg3gUC6+bRnn2oM/Fz/bGrmAZ/U0lYT2HT99OAPqyweTvzukYbV2HO
WqYQQla/RUQZkxHAsKOeH+pL98wM2fk3BqvpA3IcfGcH/xhmEsuuF5Tvjs2vOlHy
R2DMbNZFTEfHqTmKo1VJi5t8wAYd2AnkmTilAFNjdvgknLZ03CcDxhKYHFNdV/Px
8Xr7gMSdX5YIO1/M/vhOXpULdzO5vUxfGUo6kAxPT+t5uJNc0XO/8TFajxq96xtN
novM19X4xbXFjQ10+AvU6/mVvJGg54bcb1Bfs7ziKfdEZRlHtd1nVCHe9RGV96g3
MFvjVhs8iXfp9GOnQyioTwZqWqosuUN3+dViTXQaHMreJa6x05WJVNAKzZzubm9s
7eI6BviG2xrrYh6iJli/H7Nr0YRRagrVjB71lh0Hg872K9HhlojQXSxD9ul9Kzbh
GVvt/Kr7BmFPyeYZ0d3ZL2MrwUbcaMTnMUjF0NuoY8wMQ+D+tTFkvQm6AbVFji4k
OnoW4yhdQbT+usIgMJ8FH/I2B4IzrQY4YkaPHcjU5xCp6GvmoXaMasMIAWsx9GFg
oWkvTzDqyW6HOdP4JuSRNRzfO2dv8mEWMgy9DKM4EWwq9p31dpyV31LFJpaQ/bOh
3+jHMl4kuS9PnUoTHfvuz7SNiEXtwf/ej15E2vamqDVUQNny/Pm+4WgbBNDSoENH
rr5UWYbU9rhtA4Js6etE+MDHMVgTS5ohylQrpDRfokZ8TTz9MU8Sr7qNDBKJtteY
67oVj2IKJLCPrp21uA6Q+r0EbrmCpCB23ej++ppjZpqO0LQfVQ8rCIZ2r4c++4C6
z85mPVrMQSdd8JIAwCrbD0Niy7O+E59DflJgVgXkqqaaT76CYI8q0RR9OA1Gl9bJ
v2gqx0+MsvRKgvTd7IkO3DOsERREPRfO6eZQAcuKAxkkKAtKjKjanuvOU2zTWSmQ
+RsISwh95IN8xnTA1SbeIAyoZvHMBhW+64+JdNpWQvXgyY9gzIZJGtZgCdF/t223
PNB2ZqORbjCQuZSF/PMQljQNin+b5btSccVGXoAFAp6GkwNa+TFrLj/w+OQILmcU
vq9icm8hDhwSkKwxKXyCST8d1qrNV3q/6D+O6nnioFS2fEnhZMtx9gdKDsgbdKOH
ze5qtENw9FbYLV67qM9Hfzq9INBml/k3t7hF2o512A2PZY2w3JevLpzJ7kT/9boz
U9exyNKRRj5pDbP/PbcQBnPOoImZJDTcGSPXyOJ4jeM2sH9f1651HiG2NGPZZTHK
svSO2XwuD4vlQaeOqdfSLfmc1UI/x+WuCO1KS4CQr5km+iVgDo/e6CbVlgG/FoLs
EsNXuizHrEXMPxX0Z8JVmWj4oFH/aLhNg8TozH1yI2sGauOi6yCGhGfP008WYa6d
1Ec23sQByMbOWFApBNoCTsOX4atUh4oQ5u2Pi+1zjO0wruiKoZlA5GAnDuV4pFBa
WbnjQfuRDgpc8WPVx5T0M9elY+R9snAvSg/sWJIFQYd4O4uLrAq/leVHRal2taPb
p6EUuZF0kpS0F3159F2ccmuHzbviJZgljBy61iFETyrV+m9Jtmi7onsw7U9zyqmZ
he6ejtPQx2+YHYz5sad3vasoUaUuf3t34skZrFdUwdVIvbKX4CSs+LJc79QyH9/K
rfTS8hH6YF5ndYNbddiFnlskCE1AIDFVfct7P7EH85XoASkmdJYV6xmuY5eL+57x
1nHBvAYcTOXj13TfwUvAR/+dFSpaXowaW+T4ExkLYU/PnTDw30ls4NGKduRk6n/u
ZOt5MbtC/Y8pQKvRHTh1ZtI1yFnHCKxCrRFWhM6oUWaV6mYDZasHFA8Q+K7p/mEs
GCVhKkGJSEMwwyQ6vZq8ErY1HHpTmEePylEUxhWjqE9etj2WkoXuJUj+6xCA9jXh
0t7dwgSfPVixZA7UOir37fBg5ILHUa6QeFti8ASlERuLhr8eK/ZVOsTYdXzcvTCE
t4KF/Tlwj/1weRUcCwrCr5PGoUDYx9UAT0E3lTcDAf64jK6CMEROfBipqjm6Yv1f
N9tdyBbbxZJ8nNyvBCL5hLImbTdmNB6lCii0U9P6SD3494TxanI5IbbOSD6rBV4P
IfmY3e03OYjCES3PJyrS50K7JGFl/z6hCokYK6jfDHfnZQPcSYSwDPjpnXUf4gHC
gTRVl5z8QK6r5llhl2TcBcXvL9W9bsLHaQmjpWHzPtxVAC6z65elUcSgVAmFAhCf
1cbpnG1Sl9J0xSKJaeR0nWpSEBnv1zxuAFsU75YW74pSODehXsUXLIVhAXKY0Z2s
quy6DmrYYaYUdlf9uXywdUS3qvJKJ0Q8e3+uJYOED1UKuGx6VPwWa64fAFs08gwS
aaTN5n8mWxC93dTPT3XtZgjhfRWve1VuXLc9s2RSMiuWxoAp55/v1bfkdtysdBh0
P81qvN4Gc7znvsfEVL3oQwNoMUqpEoYVnxaExutbq6bkNkKz7WMrOggfMAagEqKZ
31Yj1xLDehd1D56l5jMb1y4gc8T7vpgYRkFti0KmHdxQPFz3Rfix7gcndeDDep9U
gVB9mcVfoXMPTCxcFi6ICrpXAe3nLOJgrYlooRAB7A4LddMItLLFWScyTW9W3TY7
Jzd1hBl2wEBKKc6ZqLyCFcGH33t6s7pVA825EoPKGIgqCW3TT3CjZ3hrwusU/hkw
ndhJSLodTw4MUViNxcQhmG8JGsBI87iRq/qlGZNGL052mxX2c9o1UPLSllYtNUtl
orowwZhVzHKJ4cEYpeD4fOubL3/+VZ7zTcM+7U1joyA9wWxVePzQ3Z2YToYFCVhm
dKfIqar23yIe1NOV3h9ps3gzBBhn5btMyHwYl9Bz9LhKMiTvVAi8lU341j39TlGe
yS5v65VQHpb7Vq3yfPK9mfQmrjztJ9qIL0ywTYUkotASPf61MzwAWSvooMHPDjls
7VLxYdaLCnCEEtfXVCiOmwO2NmAgXsVFwev8MUqEXt++RExOokDP3x08fP2zbie+
tNmT2k/oH8ddK6m8TTBs0ehfmfAwel82WixhawiG5DgmLq1q/EFhCg+zGpG3n4iz
axYhbJU6ZifHPlJrqQJvw1hKzC8q8EDhkt6dziVpm6bmLNWT10RhbtB4RRPfOrGR
x1EG6qhDRSpOp86QI8HQMyE4JNGGfxw+YWmdSsDunL0YgN9N1bJ9lZP5MYa8iLjt
XQy/C1lPI+34PeAQcvmA0eHXGV18TuQ8ae9Mi/UdJw4ipTIh3e1HzoyDl9VFrChm
yI3BHXw0qPLBxcwu6EyTxR5pAj+LW0IO3i5qLUUOeOfjb6Chq1dbUz2nAuYRDNbI
gCvDQX9u/AszGKpG6zdQ0zl7A2FVOP/5V8RQGnZ8ecghh+uOV/+nnJo/69r3NW2r
XyTc7dVQpUg/hX2UQhIQFIsxmDWTh6xUyoM9kgBPIgWrqjCnF/rEyHRcGtoAwMFg
tVEXBFkTz/rrfwDeIiu+Zu5+lR/HRruXSVwQWsz6CpMz2DYqHx1IOmwrUYCKSE3Y
BeOPcIPwpXZS4p9alW8WeOJbm3zXjufhzJ7q0U/fLNvz2r8LLNBFHUjFD1M6vNKz
EAU3l/E3pszxPyiqh5D3IIA4nfzZihdEE/oBkODDMIJTVCKuiDMoOXftjfCnnf5j
rjNNmQGF+qBpNTnF07S137801v6/zDvUAxiF/Ss2BzEaHS9nSFaQE8tvFFeVWbCu
xx8p/fEyYpcn974ulV/WPODeE6tog3Ut6q2TPDgHqTK/rF46sBKXzoQ2PtHAZUpr
lPr4uZsXI01FnMI4Qt2pvSCPCeiyDUsc0hxHOv2WMeL7ndSj6TRYlBvUfJaHY70G
2WL2qsaRUy6ZNAVyFMUeGjY7KkMmYrl9m6CM9nSZvNaICKJWubBcmLKJkV5sTsgj
/i7su6MskVLPvtKnArCOjbBVpz26EIi0HPxDzVLBtP6d+EFN4z+2SbqGujUR8qU/
u2fyc8o4K5S7X4s+1JkI8/63xo5mdp5AJn54Kxcz+M+XZmn2p5RTqaO77gg/ZQZW
uUrE265IQM+DZizEY2soPmeUb0w2OVjQEfpqtv4m6bmVw0BvrZuieQsTp6mzhZGl
GZ4EEfYa8G7PSaPj++UevRaCZAgNcHjgZbwinTIzlo9VMlzQfpn7mxaJPh8cjyxW
GGmmbKJK88Op1Kk13l+ekB85334xrLplXu59qFp+Y0Fv3JhYGquQ38GhwQXC883y
+T8NBCurkzBfmRHtw/uJwnWKBMee5Nr9qwpLb9KPCUT3ctKuOPXRqiNDvznl3C5+
Q1Xj5PfYrFcYb7+4DhkLMb2KKPG0qH94oHhntZhdWDRI1WTGSGctBHJB55JzElua
RRX4qdqqHzCEiW+tH0Q941CGx5yEXnYe4qlNI7lHOdpUh8+E0P8IaeZXQczhYCjS
PHXoRwWQmflswR71zc5WPKBU8qs/CCI7GzdpNHWAO1cq+MLusP3k5g//XEhfd3Cu
eb2qCKkZY/7EnlXsqEXrkWXBvbUAkdQNA7yYwf5sBG+5wuxJRbXNGoFPZ+hnNqyt
VM+MBn+l2yxjvN1OX8ru5CEMyjBwMpV0/nL6LMamZC+eZeOuykyqEWjH4X4R7eZD
LsumXY/lvLPt9mmec9o0v1kYWpZRv7uzMAAvUjr9T4QVshxFoHivGw9JBNGeJaKS
TqZJL2GCq01JD0yQbFnbv+Mo5kCW8UEp2EjuYkcaRarwYvfbn5OkvfYgbbKA/8we
dUDNqvHgyyNp5CYqgefQnsbDxsJMoseFa3hxgjqBzqmLF6x5aNA+UFMXp40QGa3V
v4I3OXVMew8VHmIxwqM4sEhJTePTc8rf8Iefo1/enlfYK5LDnm77HA4uUmy2SUho
gaRFdJY2c2nlvVzWZ9AV4ufBoXN+JrMc4UJQwVqenAbZTywT3lJ9Ec/b9gXqSWi4
CK/RrgpjkhFMyl0JcSdnVeEMSAqXQ3XKyYyZeKM0iiJfSj9Sf371BqE353lJJX8Z
dSV9JHMzt7FUwgNa/hNGhC5BroUQI9Dm84BL7WqJOy22LGZJRNwKuxHLDQ/UIdNP
Qzzrcw1yiqWa8vCCLNak/bXJFUQv3cKh+dj8i5oyTvx/p1IegoumTN5+apmsXvN7
rCbCP0341HPjyr6eJIPLlWLBHnhyf4qN+wn+haO/5PGUY3mT3WkL/ML7V2ksRcjQ
6YPsuTWcsedVqjHVm7HvWnsczJjhOrsmi7apDjmjxypXlYs/gCrooBJqYIzGdqTo
xQNjIlQdtroK5rVxM6ihMgNRA5aM3VqIXc6f9AOwsyLaFbJKMsWgFhvxZyIAkd5P
oCe1xtK4k7S1JTG5eHPaj3T4yKzhYUqSC5besy0yF68g5xYnuj499lrd9Dbbnp76
meHAeWKWjpg3rfFZ8aVeeEXaWrexdCjv5P7e++D8N4FAbpqyxUYqu5MFL0aMBKsd
BIKRCTDw3IHFExKTSqVzg+4tzmr/6ivHhMbSp0g4eva90tm/3o6ELK21hFll9ggn
eNQE2OeXj+vOIO1R2PUCvrp239jfgmPRuIkQZl5tYLgxq96o0UrleXdhUT1f35Jw
/brbAepQz1V34oJAaBWbKqgaRAoXxSOB9s89QuJj9LtWNeG9wKqpWuEQi20Lw/bN
1dd5LgrrBvi1lT4/nyIiXOnhj1+Aa0QwGvzgTits4A2REItO9Iuwmtvy4ul9Wb5T
6yyZmtI1XQO1qtgC/DYuLrwWzElBZ++r15UBTnqryb2gISyb2QCAXElFXhiM6+ng
sDDgfl6isa66uxUS6CEzGtJaZC8GwF+SAgfzajFouSZ3Z7M3Eu57I9zY9TIxd2CJ
KuPLaW9s7VY8qL0FUMmB5rXnIOz8Gbbn2rvDHqYJ25k4xaF9H6E1ibQ4LH95ewn8
4fV8E9a0JhQX4478ewDe2yh+ZyAvhRnhne5UWrdqvtB2XK1cUXOD4PWH2PiVmvbQ
GPDbOx0pO/H4rMnW00c4l+WtwaMS2iwAaTEf+yOyKQXzD9qmnW0E5J8Mj8OAvNZt
ozk/q5/tFepN39T+Am5IE/g/vmxBToxDAvtzQKdnN8rss7Bf7gTZis+Xt7CaOZqB
8zq/Ia9gjCdMbJ7rrYNx5DVsL2qDK5pg5tPOtKXBeYoXrk7Vpi6KGXaK+jLA6ekB
z/7oifqjqHLHOq5lps5adR2mcR9PhYSJ8l+ss/3McMR0OYnWEytAfEq2KXiqBywq
Cu3tI0JS1aTu3FqBfKiLJbfWTBIFD4wd7CyXTJvlRL3Dj3ltTMh3XB6kKsAL/K6n
dUgJe3dTnLutq4AaHY7OidHxdqGjkeYITqAYg/KofxHY5jnT+WKdtonxDLoRHFXv
fKcZRFyRPAryWfrj5/h/eWrBl9HIIsiGIrxMfamvWZXlBYULsAGiL9SuAj223ONt
qVw1hn4tFIFYvlRBbGlrjmvmV4kGcpT5Zmq48w3n+woFtLU+Yl97GmYaDptfMHuC
zkwlE/VLqX8YOuDRnKzB6EtaBPER8nS4aiQqhdnZ2me33y717C941vkzZuuFr69P
6NoBxgwdycGdUcSmNANWu9wDexTdm+KYqJm8WSRlenAn9/DWcva9SGVGC0Zz4hBw
Od1hUzTb8soxXJ8k2V0fsILvkwT9ar8l9ZkrUdgvLDU0YTeWegYAvqVfWg81Mvkv
d2i5HD8OXpTxuW9NjW//gcA6pGT7qmrl9QCgtnROWHEFuIgN0CbWE1kW7CYEAOcF
J797J301I6sKZP3WtYf7DEy36d1z9ZPNyPF2Knc1kiLEyH7vcVowYydJX8wAKeeZ
yz3Tnn0e6f1mBLgL+E6B7KRaeSUNdK07AW8M37x8NFdwNotVuC271Lwg5eavGZ2+
4eo677tYMt2oWXnp0cZl1MP1w4l3D8+W/Ww0LXXYesgJ3aqVpmB9/WKPBw/y2Ofq
y2mL9OUB5jSGNkpERRW5/O5cQU8P7WymS1K/6coMHRp+MfcdonEc6nt7FVw6yr3/
xO+pn4ldjr3rRb9hcRsi2O36PQbQZGUPf6gUo6+dJh10nfyfl+uR9riGb32/p3KP
a3uIjlX2Qd6le2nd/x4F/22XnY5ZtnEKOcYN0QQVlGHCXGjBPOzY5ADemT7gkSfm
Edasavrg+8suopYnmT/EFjeuUnYTBTP7/7IXk6+hXapu7v7QjZ7TeC/7HFeF64g4
bVzQD6tqMvufbh2HFcjEAZVm/WX2sjXQmMZST4W6JkFSbPn34ZX3eqlINlL6mMZL
aRVwKalnw6jJ7EUgwIpR86hqi3lr5BBNwJpcTD+xF517o8LjlHfR4DUH1m77Kdzr
nkzY5xZfJkCh49+MnGZHU8w0i6kjzFBM8nS6Rt+Hf64qElCY6SLjA1vH0tAm/fLB
Folx/HuLUPHV572Nol9IOMmyoGRcmBp+7pN7uFwV8WoBQ7zGsiunryjQ3A1A9GLR
PtV/nVAAIYtFSVGLHE20L2cgW9Mjku4smTL0Cxj3ym6T2G1hMZXgzALEc3vi3Yvt
/pf5EVc/C1SwB1YVaqvuKlRNeMrtkiv4lX+gCJfyIIFuXTHV2uLxBWj9P3VvYrHG
rHjWsbmf7srNrIUebbVqspgxbek9o6r4KjhN4nduSnezbSTjcpv4sCZaXDl8Hkk2
qsuVzDv0yB1rh92n4lLRnpNB2a9E0epDylmJjR3HA/W36qBFjt+QCFYl9SrajNY3
z/3oEv+IvEavCL7L8bQiv82PYV/GG9++Pha5dQ1pHu0EdIIhNwP1/HO4Y7HNfq+n
2gpBTVQIqkh4iKMjKsLRN9aSetYbu+KA5z09P4UrETiMSSwsx5Csl/JMYtb1Sgw1
CtRxkbgw1FEDZ2NTWzQUcHUzaHMW4BC+y1ZHraWZIQ08LV1Rgt9ZRhnGR1NVWWUe
DtljHrGYoMmLvN6cE0O+nl9p02Df+XG9gA/0e5xFV8rN1Hwg63razZdPJePhS3x3
rbx9xPD3Yyix0SzJ+KEbeksEG8Auh9fRxSPBuGK4TfpN/mN9IqLyEnzUDfYD5TLa
/1b0NZ5nT91Xr+vZ44ViSjc4YJ4LTTmrnFzsyJIYJ2UyiteSelgstQkAUKncKQO0
9B275BMo0tL77ZAsTB1f76oQsG6qGt+RFc67NvMzcCplSaQAIn4/QRn6MoM6xmhq
jDIAt5DkliWZgSOSv/mw2IMFg/hpZl+XZWE+hJduz1Jpl32dedPJvOWwmPUGsA32
TktXRK7NgXjSpnfvxmvl2bp4NALUpVaJHohty2PH+iBBZnS3XkjZ9cIZa9ybNhfC
lijh0m8R72LqrAfviyXNJlkmaIWm4kGTqJiGAA+K79U4N9A1FmFz8jlOH/roSqEx
5MOMQz2JmLBfv94HXKLO6HWKutS4tNndFumh7VMwQkleaUAdaIaiOqASGKuMfory
dpaV7nZCWXsGo/jaTse2y1KUuJSm5y2iL+5WxiG1LVfwXPr/gSHU3WVWXtBj3qIg
K2HhqFMTK0gXxvT0PImXgU32QSeiMwTYcmDDzp/e08uzGXToWTL+M43ByZ8SbwkO
V9j/Ix/LLUnq4MOJMd3EI2M3+Hy48kVdPIq79GSuasrj0X9MPaUioHr/AQ0VofAq
rEKqkJUJYsv0Vkgpsan97u3ffI7mdEUd55BR7e2LbdE9UoeIUIfydxDFAd6Qz7Vn
y56RmiHt8bh/1MgU/UV4hxu6DuMNSEVTCKfI1vGtlTkwIdeQW/Mt+JW+e63kYH+L
G92WlanNjVMjir77OQw8SIB6wgwtFgqJ497kNIhm2bWoLseXRxPXIJUTY/cWzmyy
tZKjn9ABUGAe2dUeGnilPcdtqs8nJox/GaSRO2BjW368BrH8WF9i6o2dfzzjyTkE
KcZyOSdfTxBJA2AzPUrwR0rwoYNVeCox22cja8e6QRrc/zSak1wcleZEFRdtt8DE
hDYiPtnE/438uEZ0l/F6DhPUE4RDy/eNxbmOFR2llH79ohVT+p/A+7x35hfPMelt
FSbAViYB74UfrU+I/MorAN6agaOJxg0cwqRRkRNk6YXklZnixo7JG+wr08RVsWYM
XclbDicXu5Dwi+toGzF3v6itPyLMo2UsPr6fbBXUpezvfv0KmbmQDkQLy/tP4qNh
CfVxEKvdN9Pki9u30S06ZretrZcJeJT29TmDGw7JzgptBWcQAKwpjI+iEIozDatX
N9Lflps540A5N+Y44iECab97HD7Z59LLUJVppLFDC0MpsMc7OqN66yYU9ic43pdr
R7WBtiTAwcDNs1XfExzuOvo/TjEy9yveVCQNkGrho8yO/aawfD2qwvhn+CbR0G/+
RsBOJ3TgWZARjImZiCWMSeS2f5N4DDr2bLQl799+gm9FQ/HU9bQ3gTxCXBPBNRCJ
Ci4WvIfXYU9GsLjTJ43U1uyy6Ycn38m7NJSpti4UmD20KOql97ytsbCWmD0Umjwm
hmLw7/IuyJCIneNLp28tATN01tfjt/VdmJb4Wu8qhdhwcTRseHxo1qSk4W4ug6WM
e3EuFVpB1movkR4A7Bd146hBInlA++wH0Mh59TEZ0fYMhlaPeptkjMULQT9kAvAI
aoYwdWffY67eJ4mjkl3u/VvScB2pnBdmGHdeZ996j7xER8oNuxurDuLcWS+W3Ju7
pXweW6KvyuVCm6WgzQeyNXZL95F6okkXc+8Mscak/2DMwbVdBi1/uddgmQiRBjAh
ROL5KfezWP2F8aU/F5JQUYMwrvU2kdkQbLC0BtqIBut2SuI+76ZtH9lshCxOMXoM
DpArtDK2aTy06Ot1/E6tBmbxXVvf4WiSl5kEisN28TCt7RU4bnhChESf2lofJbQM
cALZZayy8oghYmTVXCluY8bVXLrE9FOhw4l6IS5HpTap12DL+jQLFMQTYUeVTxao
133K3lkxD74fFjwHUdyypgzXWodyD6e77rbVqlXzMDtVCanwjv1bFstLtw/wci2Z
/2LdFIUXmfjByZFwWFCqYXs8cG54cvnCYDygBVboVPIjPfZUi9vl2oGQM1y2SH6R
ZvvHeoCqzp+b4wKFhebyoShOmhPcsf8M0B29GS061z8QUKf7mQG1L08wmNRj56+f
6jwXRyB1DgPyEvh/5i+LRcCLl82cejS5W1MYY1hz94jLYZV26A0TBpO5K3Wed6i/
svIRP9mEDsrVIbbUHC/M5tYXRmiEvpsWpWvUcXeKB4FMgkCeEdzQDBBJLd4G6A20
oVRTuTAFXix2vWUj9XG1enyuoSBXGogxgZHl3jyj1+DBcit182p7Zsh2eHzI/lcw
uFkiLf9vGCsnpa2m1hWCIH3QWqm+WwFrPSgoBdAiP4aZn8Vo2FJZ1WsHEU9cJUvu
sGMPEps8T0UySHNizZ5l2raZeme4uXL3nhh1JKn+fVDxOqa1YcNe1MKv6SF+7pPL
tCTlWH43Gf5OmcW/EqFzMEqPjZsPFBVEBOnYo1rmClr+u1fq2Ks8FHvjlA52Kz4a
/Nfcbs+QiYuX7HaKKMrj8m8irajLvF5CScAobvhkiVzf/9HHvFUKkhrJvyaBGXFF
2SToIiqQwAQ3d/iHjpmBBArn+w3t4sgtv8Enpom60a1n5lflBjKynzX8fXqwfK9k
htwNsT/D44MD4VdoS7vuiAQC6Y13Ip9I6Xal0gbPluTvIarTmHWh2EyXDNPkcsYW
bonn361h1tdvfoYPGJ1L5vm/iMfSRkkmK6h6Vfkm/lyka/55r4O5f2mu2MShuGWz
KN3Bh68mJbIEt9fOW5cm+SF7lNQOqPWxE57XaxajJNjMkh9xlc869JwwKfXGiv/Y
Lz34wawEbJnuZ3qppmcTW7msCjMdw+clFfsXURQJgysy5hswPFoVTqnn91shV4De
d5mFO+LJa7OuIaCQLKhQIlkvro7XLNXLT8B6+vP35+vyaxHvcZ1Qt8HftwGgm2Z7
agyc501ZGxCytEiL9xvnLh9rw18thzrTFxAsmU7EwVYsUd4eq6p7OlAV08yBdjpN
lyteHJ3JhGQrv4NgDHRDxNNThJ/gOkp091qOHAkYJ8BKPR9cEyx6cSU6atbeX+HU
wgcNgG39+koj9aE7YudScYVyrSYhhTevTpgvNXS09u517Z7AGkhOjKQQneT5vq4S
gJE6zlUFS3GLiMpMfDNONrPGPqU4fic/SaFIrnbnFh15P2lPcrAT1oRLy0SqrTym
dN4P3ogB2ZDAub8Y93DKP6YHrlrv25Mn4kNjL6zf6GusYuSTciS2eXRzdByZ/Ihv
YTN5NuwXZRgfA6R/CSgsm3dJwUQb+qNRDpFywytmjncz8D8fnyOMKOAVlLhkQDiB
6IpdiEJVuTrhXMqcEb1OkB0dirwe+o4m335d6vsVDwLS5nfd/3UpUhL3es0OlsKC
v05sjIjQW0Pofiw80FPDWNPTPcG0dhFKgCrVsOrFCWePAyvkgu4zSBqCpVMJdRn7
MkyfuOphNdZyj+WO5rhaT6V7G0iiJJvTqn6z4MfO1rk6ln/sjEe1uJpd+MQs1HTv
dhnTDzH+EW8GpWm5vxzgNylT5GOP8AFBO2OrpkIzhADY0ZweMNmIou8Ha5fVoO5F
lXalZh4tkwMkhefFxC0MSXAzvmvWeSqM8N+BGZhfyijZXwGuqZUWzIN2YCCrCTGi
cSKHsWPQ3N2sZJZKj9/orkBg66mqduYJjALBCAyWA8WooImM/BlMA6q9+MrlbMlk
YeN8xbZwJwgWKzk8bTFBOQDeNXAH8GzXERxEZ9RXhhFMf1hqF75urc4tsOW/cQ2V
4LeY9r/i9EtP9my1qd9bwGuxytkrFiOFFB/rnssoHU5BEhx6EGGBabWJof8+xI7c
PrVB1d9ZMrmD3jIjfoKK97pNx2RsCoLaHwafp6mSFXpDDOjvqxeOy289xEzt6+7C
N9EOm/ypOqXHKzXPB23J7GlW+xiZ4nrjA9cCEOG9/CxyxoXaQbEmcgxVqO1vyW7G
dpqJtrnrlYex/21D6yu47yQA2vrLUg2mIezgCUMuObX0lnMncQc30E11R9FRoa1h
T9m1zsh7VFtRNLKYvqaKnPsaCvzL6LI6xcg6XvyPL9So1aAyvI1hZRJySuCXDHJf
N6sRlVA8DJseE4jlnHJCuI7LFbSOZih7RpCJHt9PeNNm8/H2I2ssUg1qQINY3GmB
f023iTlsMinvqB3A2x9fXjpMZWHSNE7f9haosGFKOzVz836t+0i4iFf/ea/OQoR+
mDRNYjX+hkQsfaG7QlOn0ylVNUHahaA7QgoiZjYyC8Cboh77GPY0u9PzGs7SM90u
Ul6j8J3N6j2zQ4C3y4pBuROOrj8iaW8NJjeK4vSaLVgCILoZhtsVpGqzciIqu4Si
3wFq3i5SD3W+nkjpj6HFdJMl5MQxxIU+4AACzmg+pFGyKPdznorAXPlvwCZlzTzs
vIf0e9/Vc7wlDFhAZQxVC4Mku96IIUDOXrmL+tvBxjClTe19kxFgSrOpvQmmFJH1
iIfBXXlxxGj426iBL1QBP6FMv2h3ah6dUHlfdO6Ik0RDUlcVIuhhkdyMlclyK+Tj
paRXbjV57FzZBleHWaJBoF8jD2gA4kQtJl55CwEU1nRNAbJhLnJjonPbIUXfmiBi
s9GJ7tJ1Hhywi7DAjdp1Rt0JBbiJLaDhJZ7B1EeHFgdYWXrtq87xkQATt6YxTnjb
2EjKx8mXBIiLiiplNLlwPBmX6HEze8Ix41Olv4DEDu54CLHByy9HvLGTmD5NpltI
B5MCE8FpkFNW0xUIWF5SA1vhsW3U+mXcIn8XTGlMYjX+kkscqchdJyZBqDmQHIdz
Vr1+AAx13oQ9V3yS/c8Nsp8I4jrZxsKxKLYhVQJUHqwxU9T7pTs6ICD81xI/o/n3
0mEdGstqzK+4WsE2l2mFHLiqXuJPlHgQSo4x0DVuKMhC43MKkGXbiJ7ziHbuADYl
dH6mKp/GN8uFUNzZN/T3oTMYK9+raok2HZQ3ecq2f00WLV5pinOHktR5VBB26BMu
XaomGQY3/ZNV35AaCzgMgLmsNJtysrg/5I+Vw39rvSioLxtHn8fU43gGC3uQixbP
83FFKOZzmiqtsREAEEKRlsr3mxtIkpszfNEpBxNwkcUZbbsAQFidU0XLxtkes7Gr
N3fYXmuy7pU7XfC8jEPOhN9hZ26NzWdMm7gJv8JEELT+O0VWCbvlX0nU0uFWAQkW
icJGp3tM7oHPfv+kLCIjUx2xI4aQFJPDtxMJuZ5TuG3Rk69nm9Q07fms0I/glq77
MOrMHMOuhnEDbiesdQpXWhO6XW4uvj3kd60JdjN6DO9dwuymMkhIaT3tFzX3DhNg
CZXFVtgmobLLF5rD/GHDGwDB4R8id4bq98ezC/SYKysSK5lg1u3bJHrTVWJM5Sax
W3t35Lgil13MXufK5n9TDYK0DpjJYJvOlwKjGH4fLN4q/IrW6mkeemK41btcOUDj
v7qJlaFiC3q/3S8quWI5QM25tKBbzRP0IwGbUxj6xVJJcMOAeHL9q0+x0oOMLpWZ
Rn4zGwKZJAkXshPwbdPEkrJLHNAVavOpF5Pjjpoeuy9TojCikMKxeRiHTRkookzb
z+4Gx1uqjMmU/TZrMYtVZEEWmII3Y7+oTNaXkE70fPVtWQjtKpB5iC3B61X9GUwy
D9481GstbGUqIY9bBVW5xjZckCOc50U3kxKj19u+E3jROXulOSz4FZlIAakQWKTL
po/EnBwfJLFAoEU3Oof03hLlveD+nnXiISLr4CimYFfeufYP6+L1HL3+M77lkj4k
jJgrm7ODqCNlP3RTbtSf+Erq4fVVpyyoI2taRsn8BM80NQc+YTM8RumxQLQwlVuw
sxS4nbIvPUZpIFnFygqMsP4QvbG/jDmqvUNo/R+LQ1d4mOfjQp6hXyorDxuKcouE
PSkRNUcHabPArfhpOOIwsqvKdwKhvphQhua7yYPxUe+wHoA/xp8ahdXC5zfLfRbN
vrWUppEgIv20QsnKUUR+px/pk/bMMaRKDVHmFkvGu57jzLdcdgPWtiDOCkQEXvG6
RSX63sAQ1x4oXQCtRoTXW03cefiRFQNKlKHj3G0tWMQM28QNGguucPPEOVZcUqfe
Kg2ZUrfoRPSBWtyWMTWza0oPxNXbwoa7pQEyR7NVvt4/oioV2AoU2eskcbdfzFHg
Q5UBoHw7b9x3DlJO6cwmnODHtP+jy0ivjYTuL6n4fQ+43lmIWe37M6mpICJCYrzr
O6cE/I6q/fE2O+YRt0mRFRFYw3dYzIDyaDl3ZlD8KAnLY3K01ujQXg0Tjs+62kbn
76tFSpRMJatxfiXMgSX+kix2t/Hz8tRdl/IxKlkwBZwBDJ3fOyBR60DogvO4nVLO
k3lrECX0cBhFTjp63P5wBp5X+8rNGFCN8Ai9XNe22H4B6jBhohrOBLRSMaDJ9PMo
xb+941KoaD92DtKfXwszS3v9uqp/QqaqLxQTHKBLbyg+rZAfvU9GUcbZYQGrT6ag
iCMxk0A0sMrNfhmS2yZUWzz4rxEm36G4/G8Z3930wmi1wZo/p+YGDEbDTaF9iU4V
//fP0JRu4XpFcZ8n2XcrmyyphvT3lciY0+qpncJH/Fs0PWDCnVObZSJcR+Q2U0GV
o0lV/87r0tqg0X0LGN3JSeFrr9pY+79vwVblyWxtuFkoz/znGX5Oy9+jf7KFsGXT
y0Q3B7ARbwxn8XE6A01yykyZdTEDjVLt2pBeeT6VzqDeBtxrxL1iEeXJDQeUVmtJ
Mc6FcknR8S+C77iMmeqaNnE1jYKSrqGwoJ+B6LllMKAu6VNFMGFQYVEt8QgW3+3I
fHkcCgo+c3wsTtq2pUKGW1Ke+DeCH4GRm8mlQdhpDXvsUaxIttM4YT88xuwY9VtN
tIXX+GFzcDhN/ClfasdMQvLr2pG3Dzrn7DfTn0Dp0WqjsgTlrjanq5fjijCgONgW
RggeSWS3LP4wXRk9xZYSXQCQKH7QMEzzftgJ/VE/G7APJSJtqZJeBjV8iFhIAanE
03kew5SX/GRFAEYN9deYq/uJ6Dy4JR2rclsITnSxfczgAB/0T9CMBPBNv2UTVt6C
6VaPTKW77mRKRxREH9Zx3+picwQjraN9tDmA6BIlMzc7+5hU3Q/7aHhGtyx9reN4
zlAcbCq30ogyFfhHeNWT/TGwb6HvklXO8R9O+A/2WWKNZb6YsPJQBi/7+WnvIVXz
QmYu/CUMQSDvKd3nWUPdnNKKSeIjY4VFVKubNW3FQ+9QQsn4wCb9Kh3igk5bCPnN
P8A+SVNkU4dbgkQQpewzu1QsAkP+a0GDp34OcyteZIX75qyh4G7bI/6udFA0nlV2
Er6647TU3gIjgM2n2FjD4F7PUvpnakI+VSaJUiZ7SXOFakty0u+6jLhTNFpsxb9c
QoiixdugJIqXc3SG9F+nidi3V++LcdzCTIO62R9OD62h1Sm2vshdRV4YxPDkXeK5
HaYef4yDZEGrP7FtQ6oZdC6x8WThyILva7A1FBxYhwDdqUydSNUyVxSMFKJxeYwG
+YAtYnNg0iqa0KG3xFDtxBRGPIVe6fiJ5j69Upzen5X33NZ4/HWVKoeIpVvEJjnL
TdiRz+1acMX0W+JS9Pr37HlzIZTQ3c+hFDqENHVljF28lgAGFnXnD2NDlDFBDrBi
JjoRJLKIlo4Y4rlVhLyU3mto4SW14jz5IdKrHATqVY2hzy477zB7EBHZhuzu4Kk8
zYaa0TtcFU1aBzC/8p3O/YFEinfxs2fVTORi2irhAMU8+/nYHNlbu4g5tMZkkCPV
Fz3eOcQGTCOQwCpN4YUniAuwoYgMEhfMwOP3qpUSwTtin6fYz8L1g3SuNVjdOHzV
D3s6gOtkG/FgnQZeRoOmqYdFHdaD+xLgUlJ6A4x/4RUn1XVvrSGLGmMkk7awMztG
AzFoT8AQDt2/TpJKFh/FemFP5ZI+MF43/unaiQjM7/8S690JQitZ7aE8m6rNcon8
sH4b10CiLx+DC3wS4YZ+9S2Ko7nMLXhnqqCR+/eCOUyZSUs+WqPorFPVdKjBzkEg
+2RCLgVMYUd6cyCiDfZ98JF8vReJ8sgAgShnHITwmGsrNQnK44wKipkXwBwrjWZJ
GHtZZVKxQezgKariGw+GFk/guKma2IsJcoBrJmIVrxHK9XEea/Br6qa/u2AqBsGQ
2Bqdks+DgC81hNB5PX5RebNwzMgt8Zu3Mt4H2YKJHlAvxsGLNpdru3BLh43jOA11
11FSwborNRb10kTlRCG3Ajdj4mUkB3IJWyGU7tQcutftYzo2nlWkN1omblWCdnzp
vd6b1S2da24mNQgeNcljCX7e54jKAYACARUtXE3onfCbEYKdaVGG8xIdDAId2ONJ
xq8pxDg+JlezrKo4Sid9Al9iZ5ZmqryL7bD9y0woRbT7lPdyeP6f7pTWPeSeiGWe
Knb3aRdI9c9DoeqsTQpkH8wVXBWrI2iJs5ndSNtMfwbYQviH56f3YTf4CqcuZvoW
j5YkgmbhoXd6GZP6+aBixHxpszLQN9esGXEi1fZ/kw6uhMx4v1FNrgPtPJxvFm4e
qj3ngyaIj/rhGu0UbyMI/JPdXPyMP4menV5C+GqWi0I0lJy2U37WTgUrWRQgNvyd
SY3JQex7zK9Ob9xHCyBv3j92CBioKydnc8zqiYqQ3gCWYADjO2lYr2y3HzDw+uXD
NLoBt8mnxuab0Es87LPLD5OVhVJdXhi/eaRB0jhgFwQOIilwFYrKg+rh+qBS2lBy
sNLjCGAC2RlTH7sUqpLL7YP92xkZLKvcEqvv/HJsVGZKYPekCioStfhPPXANAzTs
BXcaX251gRulYL8CYQNnNC/Kp84NWy7wkuB/nOflLeFvZXwkfgMPax+DeqHN+zRk
G3Cgol2JbFwAiRW7ygH4y0698zotq80rO6GzN4LrjfpujlGPufZqBxSQVRf5QuuU
Oth+yXDOv4WjgRpO9wJacpRjQRuikAh++262K+wB90of9A5ztJVHLteaHsCrfZjf
eZj7wPs+P8b5Eix9AgzEo5Ri6acHw91iOy8V8tPhxA8AC82WzSkGvYJ6S27BnFo4
dwGQbYH3tJOzR7MJF2deVsnNHSaU/zMlixM8TZ4c/N/0htdETS1B4LJStdwocxt5
nj45XjE6NjC2X9/wCneiwZNcRW5HxD+h7jOiQZo/o2K8xcP7ItcZl4ZK+9w5yoYd
fpH48aVhgUDqct93G2KRRND3pj9JuDduxKs6LIHJ0c/wsAZV3Zs5K3RsQkogutSG
xbBfgXPnSzV8FFS1hvTGVrw2PwjVkPX3zXnvlu0I4zCYi5oYVGVJCAtkdBUSGsK9
ODz6JYO5PfBEyRuYnUBAXkC3lTjhq0QZ26YrvNN+QjUMrD7pUW/zBCOHt0Elg9Aa
KfgV8QkPaIE5+/g8u4rnm6Ja2l8roduLR1Uc9H6mCasbWvcNZOpm0qMD3xhs6esr
/E9I1sRphPWucQda8F2lYz+OoTWrVMLAfns0aw3smbRBfk4UDE+NvATwUDEzPMXF
/Tol0fd1m3g8iQaL/fzTbPAjhMwltK3FbwtGqraHTlP8p/xnH040T1xzY6Z26Jry
s9HMg5G3R4rlnw5fI4gQL7nDnExsrQTFeMAux32C5lkUY5PE1b2ZrJ7mIwqad3tR
wBSDOIeigy1qIfBjy7nz+WozH8hKUm5LNUrSJ5FjjHYQgneOSXVuCykA4MjYWtyA
r+6aqxgj+k1E2Dv2MfXVpcQ82dbVX1cJeYZKRC1+DN+RXLNfJcIGD/x/IFeGM7XR
3LR4iSQxy8V5JWfBppotmfuXWRylfj2eC8i+uJV0BTP3N6JkHR2A9e+R/rW+mt0N
uNL1cbmPLMW1ZNZjK5GlfMnH+nmuklC2nEV8w+E5qVR0yKX44pMsW1UKYyWv5gPe
Zl4Popal2dCdF4iM3PbqVY0PuUPC5xFokldp7KKQm1g8rkOZEjySpnwIqK3FUJtG
OPq17hqwc0KZGvZyDLg1eNyviVyw4LPCRsbnJSD3poPqcCXy+s4u7l8mrVX/p3ZP
UW7HVEGytjij6vADiI7nW8EFo9GDRoV5JpSxaPZIElFCQE+9WLOyadRQM/AEQjhL
COE6elk+K/ohjqpmO5WEjnAFdfIDshUNcK8HEU0MgD4DIos9QuS1Y0p1XaGTgE/t
ZZxLWtOGozszzK4145ICgEQjCjfUQfezI40gfPHp8owceRKu6ou1jG2QCeAugXm9
8Y7UEjp7wVUe4eod97ylu8LZNTKJLq5P/sNwGtM9AhM6TIDY7KpXCAFIP2ByVSo3
YJZiRibPrREHTGylGgzp5kN1cOJmylpj/1OT4g6ufxFk+8VB7iLCZZBsVSu7yN9D
CqCnWv2OtYE0aPmNwAITIw4hGTYLxRbpAK5nZy/o9l9rpWCnGvjwHPi02NoJHep7
Qcn+g7UcJWX2xfY6+pRNpffMWbwRbY7hHkkyr9KfQdki4yPXB6EXP1iP0BNj+LWb
ka34ddcwRBijQoKy6RaxWf6fnj2kPZ4fX0NIBkDhAsG1vHcR/DiLs2BkGGbjSpRa
rxLZPejRI4T/lwdPDX2TsuwRTx8pi1UlUC0nlESPrMWekpTgmUjVrkakw1U+9LWh
H/G7Q/GNSQM04ZczRiXhG8cx+lP8NsK0eq8g7wBGp6sdKwtFfyiydcWNjuDHis06
l3Icc6Mjh0ST9IqHPyGpDhnub3Ob6lloHT8X/XOLyLwGGHcSUjClgsQ0K5Zrb8NE
GcAush9Abr/URGIyMSmtJsAnoLDuWDNi2UTiV56MgheSm/QaRrYkLhC10Jb9FzNh
G64WH7BehxLG+mjcmncA3oYBKU/EMjRORO/egy87S1otgEtCUlYWDyKqXrzVnTxB
GddM/kDvc+Yqxd1Fp+FFl2O7HzbUo4ZW+fTVf+yahYgKoSF/1fr/qa1R8JXjySYi
EiplcTv39TJZ1zPBRUKka7xTRppyCrOcpBu94XI4jiz2vaTqXazW1OnGeCtoJvL6
jPE+9iE0Ynpkqy1kChOfvuzuhRWleEnuRxsJFVsOBg6aqslm7XIwudOaqBU4Zogx
vqercJPWQclEq+gYESa+8kL0gII/dUQCHfonS/SumHiRveGx6EhcishvpJxjPlEK
TXmbdemoe8DdkT0aFlE7JE2k8O8YevRuCAWFOS86WAdy6msDRkuq52d/1XBc7/wW
0hTnEg14Gl8HXxlQRilCoZxxdgTtCosvG4m26ub8SAKVASlg8NMgyQAwMi0bV5PI
zJTqUKzlpGIWldXA4WXJvyBvVEjmNBXCEAQ7V/dIP0SoMsJ/wddtJZuv9j3T38cN
titpO7WvVb3WZJtWSL2CLG3xiF8ZXoCaduvo4oArQRhdb84LIODZRQm0cI8XTQUw
3ME76up4TK02H+uZbAiu99adO8O01T0/8qa3XSL2PO55XhhwMRrZgP67ggHeShAh
+Pa8RUWOM4CSH2r65MJ6jkygQ5FeQqhKN9JlSLqrlx1ghrvDtvxPzLDB41D/aSbc
jN+fKC1sljdlZJ7ZRKgdNLNsXfAs9Kp6qRwrf6DirnxWIdLDGCdfNoGqG0sz+Dsk
lpEvTVYqwLRkQAOwsPY6qZh8lXiaJARMvMG9JSbOpDQt3osC/RddnbaQi7mrNhLl
Bb22pc79y0YuQ8mRy2ZcXTFgrztXufsKRiRBugSHmqBGoy1rP3xvHxcGSD83sqk5
8cuKvP23D4yDX6j1cVcArq7gYziTjnhmamAKvZnAU3j7D6yeupqWMdlNI2I+hf3d
TN+REqLuMn5LY+driMymGqSzMrqB6esHU+3zkyOGwV2syhGXOuhNGAosV7KhuC8C
SrbwKTSOXLcdfXC2JAfcW8kDJuta+GbDwWT7ETx1ofCl36I7UxALYlXHno6diMNq
/nTgpW9Iwd3fbTzXQFJjmT6N35uzgpLqQbFOKG3Lz5DOFEFOzhbKF637C0QmunWe
jcl9jge+2tIKCgyTcAwsG1UBVyOmCEX941I9mVZB8mK2wBw2rVNJCKUfSU29s6Vs
mr4BwdmPhf2EzYf9jmQVXG+wOJnA8PrxHGI5ml9RbO57GEIulvtiwA7+sgs81B8E
Ou+iIfTu3H686/E84YaHrZUQ38nM6usjgCfiNIR5/mD1+ji9wDdzmxUGL/vHm49+
OBPu3WE1RIDfXWYNigCERB4Ru7KE9fQMBiP9BFxeD3jRXdbbzdrM/NqaRQULqvvO
Kobyns7FfJJad7wYT92xGHesNqmbonZ8Y4WOl/BWhykUZzKPMkCtea88DYn6JhFF
Yt190yYNewBJIQO8QHtTWK+2jnpf0C/JMvWR0P16zmH6Zoym/1W1hiKqKVB1VAcx
51yaiUt5uSIExDqblXnrp2yuWeYyz3Z5oxXG8HaYUTDO+nl43OuLfQ+UM5obufxo
af8m9eU0wEV2Ue3/lhvvl+d6E0dWCS9+GxzC2kwfPxQ30CPu7w+aNd2LMTXA1SXU
UJPf277+UaenA2xi3DIDUuRWT5WcZQVItQv65XhCjqtCMbHmpWHzPuiEOJQHBn6U
XGo4MNAwshAVkSXPn8yVcsdGjNky7kpYJc7X7i5R2qpjR9hVfeLE/I/kEjKjYaVG
XL7eYQYwhSuSAYP8b3GzOm4+4ToxgXlKrgzdtGW0Ei4sACcLBnKHimva6WWjPDqL
GkWDppDnBHhqdsvpQhjBf8IcaQGNfFM+9zHQrPzYzt0fa5dYFYN3LwTcH8BHM76k
OdlZZ7hRqYOVCbvho1EDmVcZc4qyN9lu4XmU+9Lt9Ko0RPCPHacD6Pvf2o4G63rp
xppuBgCHBdVwI5B1+7wCsSdzPH+kguPFNjBfxiDoZb/SzDZEoL/QdJxmjz7ajRDC
Mg6N7QxopbWZMeKu11CbjJztVFFytfYlo+jGq1xoW86gtnbO1JR1f4d5ItXMEBxR
lZAzAKiaIyZbOYtJXrFsEmePKzniiPzqBE0TClLo2KQVEg/lXDA4E7DQV3KjFBOY
bhsIFyi0APWLv8OIIljyuqnz9NelRNyM+bDn5JvtHnzukSErw1atzBSX8YXSuYZZ
f0bfW2def3zJzrPPdD8cm6D8LmeZ13ZdvKjI0g+1GNtnl9ggajGoXHn1kqIPU9HJ
Er88UxxTWpEPvjMGkJoGF1+++yEFLsRYWo0gT0Kf6CUOQikD5MzVooWRnNBTYhks
v3/luOtO6M84ARe1q+m1Lc7kE7i+2HW6UykSH3CNmc04o8GNm2U3BHI3zA0cCnuu
coYnWDdofSIA5rWYe/ktgtQORAQex/MfKPEow1o4wuymk9T0DBz36iu6WMXF5s5u
OzoWrqjlQ02xZLD17dV3h9PielQQwdMUWCm3TCWmwpwR9TSkr/CyVYwPSuaygBQd
dDW8ZkJvs6TogrVQuMYqL2a1aYu9JfYmoy06S4jX+b8qiT1VQy9w91cXSwMMtVGa
w9bXPqLgmfPkaqOkYcROMsHWpNrFX3QZ3pAFzGy1bq60uQ1VGjSJ/Y6LIzECh1wZ
nkQOnoDdO+yJNxqlhZhrxK7B755qwf4X9bgmGC9qP5SaamCScdIt/2yWno7XHc4i
Y4QYYTyau4SuGtELresPvsGHJkcu2AziMVYu7rD5ysoaKASC3ENshlDqXbMY+Dyl
JhoEdojDkuNamTPrvXe7l+GzJ/2qqW72QDSIhr37ArdzyeSR2tChhCzAQJ8wjSRR
s9Y+Ih34J1YRlxQEN7QssVQ2D1xyPrlVH9gLN1ES93jHIdIsnz04tjATGkopaypr
xtgRy4iL7c759wBfj2oZCwvWmVxKXN81AojwW/XmdyqjYpGB54MbmjhiVbyQ6+vB
MZmJI0z59f699TwXhMECvjI9Q3GxzzTzQrjy45wph9K4eU7YvoxBlKTNfGFpVn9n
zoIenwPf53LrMNzCie7e9qi60FLCzlZfGxc+Uk2Bui8DX0oBDJ6nNPx7vleXrRIe
SnZHMUpRCCPrIK6qKJI+IWnMwlG/myDL/vqUS3JW9kd9i42edmt+w1QIQ7OmwpBa
4iZbnpJO0R01MB++osA1rI920JyQI4N9PiJO/QJMN/uR6Ea5zkQCL28FwrN9UG1t
zqNapW9I6KlImP7bctgvtt2pyFBBT+Wn24UJ29J59DuqXEcknviKhtOJyXvh95Qi
xMjBmVErhVBmqKjJu0U+SXUl2q9o11TNsqqazQnwb/JVtK/EYyD8muZ4fPlqav0O
FvhCtkJAJDlmfva7M735z453WwDvQFPmd8QXNvEsV51YTPFHw/Gntg0s/KqA6/Bc
LoxRqG8nVKqRMw3gHUGT5dawl/pbgfao/QP8Cu4cpXcLta4cJcZcWjkUpV/5WNPN
8O25C41Uig48W9Oky8v9BC7G83HcWc9cXsdolrOz3+1PNjSlyWl5241iQ1kbL/jv
2kwQ6L4Pfpz6EErxkT9fZjXJT9W8UvQgft9RltXZwQ3PRaXrZbunszu6PdNqgiBL
7qw7d5wfjV3Dw4H6XD2UwN6MUmPhgB/FWCx8JWRFDElucmJOzs4TuLnRRBhKePfo
qw+cy+JI3VGqOncmxlU/xcVJDZxHzBDXxOFkk2tqJPGxCzgQiOXyhCWhRGri/Xiz
WlBB6pKJmAzxF6Or5d9lB79gzfV2qR/EJRoELfN1hsNc2Wfz3O3RUUm9D80aoTY6
4INpWhya/yH7JITTiN5N4jUbaUkUq9icruoDV3bBdDLkjaOMY4K6VFtzBK6hKpAz
jmjEd2/kfOMPtjIro1ayIv7NQWwJvi92M9i2OYqEvf8r5vNRBoxYYnnvvCX8Oiv/
R01NWbtpKiKjXgOx5v/B22/Dz0KoUIf86dEdOVd6euR1ZHV1X864pNkvf5YMRNtY
RzYrLDi5leyIkO7hhuljlrqv0gRZuWbs4augrH+BSm/XjwhKKrxufWNOmJZ0bSZo
K4R7WR6cj6wzRPuOjA5qP4xZ6D+HGaUXPAo+0XL62GWj6xaUqqCFhybL77Edn6w7
pznkZSwrJVm2MFddDxPAZQujXaWM0RzyyBbeZroAR6LnmXHOnjPKV3ahDiCBXxhX
lfdcidtVAmNKgQ9uzXPjA/WcGv/YUrYnDfDIrbdeeK3q4r2QyXi+5yz7inRNU2zu
63mJKdV3aGghHQtW+cXdPn18pZRyJLfVuk0Mp1NAG+4rduUxj6N/gb8PfAnOX0KQ
K8vTh8LKlZ18VUoLub4ZVGNt4j6iR/gDN/meFSWiDjcIgbbcJUqDHEKih1kd0vRj
OWPA1CmK0sepq9NQIBpm7gz24CgwuBSspEon61YANcKFaDM3FD+5AL3Z+H7NsSb9
kg5oK9M1R1uNtQOmk8o4ymM4ScZfQFMwzcc3Mq9DEIXMbxKZKKmB4XIZfT7ppxH3
oGU2zkdFfL1pfggyzAxoW6tfAyvY+ruuTywgXnx4p9o0ne/ddH93cmZWFn1is8Az
eg+WEfHyJ18j7gB8nkZba8sHsGHAQlQLQRYnFAD0MnCWFXgQuZ9bFm024fyiaaxL
TbPyCIRiyj16QRNxMhjgD7pOGKnGTQcc0MgV8tKzvCq4C/0KPsxkhTr2G3TnZBdT
RkYSuhLl4Bpc/j3HSB2bUZX+YpNIr6apjkgFxc5UO7UfYg3SmIUQZx9r1UOxhgpy
XaiMD9liQA4zDniVQdOIbMkSdHx+kFukatWzyf4HrtPXokhV7BIlsEyPP34wbNIU
asfGjcZATjciu33G0bB072w0b8H+FRxGtAh/nKhalBpJcBOgKHY5O7wJ0AAhBKub
H0f0oqAdKL1h3+AHBqmIUKiL3vWhJtiSEyAGegjUH4gbnLbYx6G61sVpYNNEWGbc
KTr/mRortFUtWv68Hi2qg9RelnxcK2DnWDUj6H0QvqFcCpvh5R4ppN+nUOWzxmH0
vBhoTcUflg4J7kvDdDhvOl6353IajUJ1sNHmAbtbfsgaLj5sYhCiP40sG8GmfyTb
uTQHJW+++njlYptSrO2EyHO5qoGsJa+0WpAat8/atFAoo39CfDwH0cMxrazro1P0
F5yq7NS1iHvTjB9HFqOv5R016nUPA3+rwZJV/gsWxH/gPVBnswu8Hu7jCGEocj2/
8QHI40r+7cA25Exjl0ZYIlblBiTQRIk5i61Pz6NSMKbzPibDn4cJTXJACG2xsjVx
jCeqcH7Ptwp1O8/xU7YUX5ksgmMd97I0pjIGTaQ2Wg0z3vuOOSZNzGzGhcGttcrO
wZTPrQFOQwiWwsFqQBuH4MfmBmcmy4iq5RbLz9oAPuslpSCQHvFU8E+HmtRBg6JE
1q1kfNpfk59suKvfb7O09TM3+KbqKrQAaPMYH2OTrpQ/fWQ8NPAQiozeSh2ummQa
MhhjS6hECmfIlJjOICfC9M+SZjvONioLAm27d1u083eSuq31rww5l+GPNu2UfBJf
/FGFdtbaKSP2GWOiMhSH75JcO6BHIzp/LjhP0xHqluJW/1/uZ/LAgFW0kyQfG70d
hu4Q1SWSIhbqm/F5t/emPnXzR1uqZaT97baZfMl4UGvs//oP4APtlEeVMv4R/gHP
ad+871fpUkvXfjPIFxqlq/ZzScvY2Ldmx29qBR7iSjdRMZ8QNJWWsOckNEv7gzPU
/fbDL1XioAn+pRgmizcLTOfBG/F06j4aJZ1mM8xzVe7yk/iWG15+JySCIBRmxcgs
VBxQ79SptyzzLo9ygui8WyJZ6QaBJ2sWwE/7WWszQ/CC0sjZGUw2JgHA9asjdyGu
NEKkjVukdutodHk+L85mbfBocgAAYHc3stJ3d78ZfYWvdaRvLrRj7NU0Uez8BFgT
Vyj+tNVu4zsf9zo7gVTHZOPIVR/ntdx61mRgA5vAdt/YdLxXra4QxQz4Wze7UJBI
Cbs5VYfR6f00dsKUH++LYN8gggg/Q81EoLF87rq7H/JTuM3RTE20gTuUgFZn1sTB
CXqyl7iE1eEVeKSfHWMyW3A/psdBa0HqCuIXLHSwASqY1vSyWyXUvcTxCctzeKvz
t6z392GjmeozUzDmGmR2OO3QmHzva/Jdf3mvIXNoh/+URP1rwbowWkwsiNBLBOzK
/goVW6ZrKqJ1gCMPV/IW+Wk0Wc9+LR3bj4LA13lEOKxQbEPc/E/mD/42eDe0qJkU
uOhSnGx7hyz7qPp/uKi4/a50Yncsub5Cq1xQ4pEZTA0ejbQVE8SO1szMEtQPxbTU
FzLPA2gSI0YNPUYWX2VkGoSkQAABKP/SGStSQa+4yhXgTWEXdUE6XaTd9InurDHs
VWhpbq7w3rS+D/JHRyBwqz8I3/cgyzx6Jptuq0FvlVYKNLWGfX2hpK2FiIbG84JX
GJHRzfdGLZlkua4GNjHNkSXfG4Ub9+g1vXCm2ZgAZTp3LdIrP2uuSanRxMC8KdXJ
1MGeqsLdaGCZmZxtaXhJl0mW3MHkyVKQiqQAozHAzvj67QLVXK8mPtAi/8rz5J8Q
oMTkKwEKaXC73xJPlq173jtmka+562yrVUdHPXyytxxSjkwSAKZ44gxYK6kjXVfo
hi6YeonPGjeneLT4cip0IkjntVWC8HSmNHvPaZYG9V/bJ23oyLQvlO58Ha7Nzk12
mGN+SulnPWOgwvi6XbSUO3T6Sf+PxPc+MzFXdG/h+ImtbrQqvvNj6dlCIKy7Q2wK
jkUgNRCTZdIG35+yHYdSpmpEU72rKxGsJ+E7HQOeO63pngyaAU230wTdKJ2DFZAb
SOgLT1iJSO0YVj4/5lyunJ6j4Qzxo02qGbSwzKIzWCvUU6oEY2I2lLDuvpah35XV
7kIKrxJg2TFa30Y3daGJ4dl0s/fGkJH4GaJU6iS0qD8ZoCBvsdCGjPfj1yF+5ARy
j1e3YVqKGaeoaxHlbcAzGitN2u2FsUW3ZBTB7jEPF5deTs26JUOP09LzZWTxiJTD
uHSvMICutvxIIcCvK+AVMkSYPg8j+U4EYyWt2SzYU/aME3k1QhaJHVu1Xfx0pwmE
IugmFC3bHHhXWWBMsDqxtfgyOnclH5aCQ/tSw1nIUzdxAthWxRN77C3orzCbwmuo
vX5s5YLtfkejzIyA/2DJit2Geto5MjpXT+KpimH75LJdI0jFz5jK17pyool3FUfx
i7Sin4/f9v5XXogdIWComTPazg5XHl+1HAhPoRd0aSpLY1qOQEksQdeDnDL1gYEp
gZ4jCCwfRGEKLoSmUL0PfJx3iOWM1bDF0IRcKTxGtXno3e8Kb/ZDllUYhwe3ZSwk
XEHhe9+KMkZ03EW/3akda1nM+G2+oSQaI62fwfZpHmTT0nB01oI44W/et/j9jYkG
oV2oNH0Zy9AjzBMsNgVPThRIH2Op4LnkvnP/uvjZ5siojMNbtltfMeWM4nr54fjq
+X5Kezylw8wlwm9ZlreFH78GTDl6xbSGjOtmKkFpraoB43zj4fA8N6EcaEbUWOuK
hhWHHB+9nh9Ao/FDKGFu11SptWc5eEcp3FyYVF6t8Db6Hq5pQlTJUg8TPUTpnBQg
mEWh9HddBSIYdXn+qckl6gFPPzYFkTPdALocnIBGrXuTxc1FBpEY5/q3lIfRwW5x
pVqq4qjyAP3wxR+64djMHAB+7OtNyIMKYl3QAr9AKx4X3zPOQobznsZe4oaKbmw/
4wBcZbQmN337iKv644Zm/ZCMvcVTU6fJrOYxJhENDu0l0mHdyF7xKeLzsTiHPXhs
Dk5qxcTJ6JrDrZX8XWQBIxlRdqSOlpCOFQN5LYOZhl+wNq9J3DOZ8WgUsXGPH16b
zpoMrSWrwC0nPG+XncEC11fXp+wqDL/pcHwagEiTt4mPZqh+LgUBK16PPeexR1QV
QGmFpU54nishd9K0roV8w/ieuA5glHlCX2xNfOBVYpxy1cKFnrjx7dBG6eMW/24b
ScWk1Wm+9IX2DqLoRmAM1+mwx3JneHfvwDaV7zVy8LYpvtZffhphIuUbX0cinSjx
TatHMR7JLz9pALBMNHD19jw9Zs6WqSCBbee2TBqqVsukPab6285oHmFVjLQuyJcP
HVZjJ05gror4szg1t7HL4021rorPcbpln64U07Wv1tKGUc0/TbqvBjERieYIsWZk
p3PSG2dR8LS49EmMx4eXYddvSrlDlJ+Q0nFU018AWxKbif0RFt1uFMehPrazyfTr
J6F9sQ5ze/K5qibOTCVxUm+5NuQ3d4qhmDKKahRPNtxAH9/uIlxhpS+vrxKWmBMu
Q03HAny9mHFnh2MJGWn76jm1dGfvkj42XBk9RhdpJBtGk/+lRKCmcfM0CGq++u3A
rYavYQhaqFoTC44vMDD61YD1fAltvMQ3o2TLlJbBW/+p1vKMRV2rJA0v3eTfG3YJ
6xlUuOROyp7NKIlFFwygAKs9SSauftEzhWfWN4cuvUMQwPkrtcrcLR6iEZt9YSG1
Q10TTYP7lLcU5oW0826dBiUvYZOPWmdNeQiZZc/yfCgmUaRCZ1Ie6wTeVlhcg1I2
n9IbP+gePUct7EPmHZNyBkqms4BSQY5terjA0JhooFNhf4RIZ4ccb1NSUammjmuM
DOb/mVlyPIJPx3cYi5N1GqU7gCptn+12w+O8l/W2Bqbm25WFfrqL9oRZ6Ic/yBgA
R8c/ZEipUCtFM8EIfVcQ4hfJWV1sGK4mNEhUYXsSi5tuz/X1ZAZzeSAjq+TWfupN
VZ9hCAfXrafzciHmWUhYhS1NCzSuAlkLiLWRIsjiF5uKNHMyeK1QPaZpGjQ3OCWs
C/Qt0TjWf3wv2iIdRGG8g9ww6HbVp7YDUWwNl/dRPjmnQGT7VJzFozqdUgbDIn6P
5isZIy9Wh7FH8hahvCRzcHpt0SVEzqBQ2xQNCyznBehlqJF0tZez21kmZnQaJf5R
F91nHQoWpD3LVC4QPem2C59uwxHryaCUWo6vY+zF+topxxRcQWmY7gG94rcuGpV7
O4btvByz+XMFVmhxPKk8k3pVX1qny1aBH87Bx6u68ajTqQUNmVC4cE6TTN8FXOFU
uGqs/W/D7jlqS0Bsxo63N6UHn9SI9pNFK/h413GAc9WGsp6GARZj7bb0ryzKMY0d
/NRfLkR3lwoJW7Aqh3/RTPhP7Wh4tWV2V1zzOtUki91BPXD6uLPdOCDd2HpkV4Re
E7HksrDru1tuVoikyOLaQHg80T01xFqMqDmGsKZ3t3OaCkeVkOJL8TJyOpzByfy9
sa3Tk4r4Qt9tGoRlZ2EvACRjzBgyvYe01FSG6ZY++IH7x7vtZ1TUp2HmtBuwr+UH
zSROeHt5czjq4kCaAvAcfA6udXCYmwH1IIKpCYhmdaur4ib5EquI734mssgmtld1
2luX94++XpfMmgbhsiURuv4qoLZz0RxVZesdNOnc7rEvhu+JYDUlfNxlAxhQNwBq
jViNPQa1Tu4bINrdGs79Q4GvsZEOxeviLUgsDoEUUDzBQIaoNSB4xcbzpp2/440W
2rZ/bwi5JUUkcl4wWiLH6lRhSBktisDx2Zkzn9bswOUJy4zAVi7Ai9hJIqUvKu/0
j3AKSlSg0cfaygRWwuCcR4uqlQPIVljLLpyXj7nTYMuBW0Yjujt/9ZpIOfkNBOIa
AkUaJacU6NIyFLiydlaJAHN7BSwGhjvAzvkp9xEBXoyqkkT84iUic2K8zr6BtXua
5CfSIFiFwuqwtJcMWfhCb6D3oh/tPY/MCvOl1+0mEa2fbYn7i7XdFltupZU8Zenh
H8GG3EjvjaDeJefsCOndPDGDuEOfVTPdsItGE5dF3Iosav9sWH8LpmsuqRI8o8aN
obspaS4FKAUTwegkHpUs68Z4wpJBjnmGm3PBnvMc0bIhbkhTD+x4qGKIJnoSaT2Y
GH7h8QTEgrbPGxvZYxIVdupvKx8pGlv2AQ4kfORdalo1XPSWWStQgSlT8af4rWT/
KnvZfs/JAQ04tSjFg2s+ushRrgNQXqdCxG7N8umR+xTPkJ88SpzPx+7sqK61FrqP
Cj1mHobWzjOfNN1o0wAH5RpAQNdHJgrXA0xJP3vkEGodrsVA7rpqo2lIUK3zXa6k
Xrx5zTaNUc44fjJ3TLs5In7ZsKfb1sFNGIRz7Cq9KTBFkXJPPCIHpMLynEqkP0kZ
uAfGk7cxrfO7DJ1gCLn0oX9F4hA40pMAQx43j5c2oa30tT1A7qJSi/6Wfug1CJci
DgW7Rm5LF21nh5AYIOgUSNZVlzRmdpIL/06R25yXxcM8PS2IdF8uHs2RkM83WAXV
JjpPIa7C7LVquYsMO7vmrvhEsKnMGfjCvvCGBMZ+H9BPszP3U4Oom6gOV/R9AHwo
Pu3VTvCVh76qqhGyNdt/MlJqxZySPGKaC5B1cP/PCxFxn096oJ1IKyeA0ssfZCuT
se2/tKjjvQjsUhZhtNsHJOJ1rPybCcVXrwdBZ6OQ+kv20NCG23jUgJuiQk598G/Q
7k3Ccent3hB30HSBPgeiRNGXegLKJFKWnyC+/n766pWGnVIo1BdX5TD2gKZQ/viy
4uo58l/R4K3OBYDjLl3jzQskysNh2Yk+DscD67yRiFcneFiFvgsKVarR/ng/XE1j
MgybSIPbEdQSynK438zmaKY4n2VDfwtwZnc0CMRDGPZ2XiLre3HN/x1B4X4Jq0+p
ldVYbvqvvSRZ83db5uE2bPtTUI/HvAKwoIznK9GwuPtvVd0MMrzzClwo/mMgvSiz
YO7Af1u4PoVZeEpU8Ghs1SSFnsoJWOct8frRtAFPaVTG7YwTYug5DbAgHxmkecFP
UYXHIjko3dcDhLe0BUDwXmlnQ58nbYtdP0iezc7XtYe5L8gzoxUqGC5v+4q/xOW+
iKdjZw1WJimNzuKF4mv0tPbp734LrjtURJxyw5GanRkW4eyqwpfU8HXBC7xdrrfg
4M4MqcIPTPmRurbeo1bqDYyV/mjzOeh9+VZFdwDDUtx1t4CxGGhvecny1kd2ogBK
zx2BPwsU292/vUPYIx96zEDLybfUzqLPJAGp8vXrCERZfdaCOLvelkPC+Ju7JtQp
hlzy7xRKoYlH3Nn6LbuaHVmhCOaRzwxLqcJ1Dmhgkc5Pls0M9Uc8YJ4j4SVgDFs6
+DK+IjnS9BlfxJNDs2EOD/i9SJRqDuupT13Fi6wMkSYUSceSsk2cmyBpyE61ToG2
8U4jJI/C7EykoXZ02YYguzOttAWeJ5vDszmsSaGxqZNjSEAHMCrulic92hpieXBB
ZrWDE7f58STjURKk9d5SCPccSsppi9PNFxZ1JFkKaMOqpjljXZ812CNrPD5Upv7i
cipb6eEk4qy1PJBOV8TH20QGteOIimG8m1aYFLaopdtKL26kR+TA6Xnnn4KOxA0Y
2v/QX3VrWyJDQwoLOR5z97S839x8gin/lc0WixXKZJEc694lSOXwq0KyP+DAfhlV
HrzAfa5yD8qAJvWdTcyyKKtr0xnWEFcnA2Qw8PSUqIHyRPxQco3MEt5ZIERQCGE2
dX4Eohy0N1oAVqtmXrEGkqUrM3vWld39AaQAcwidAFA9b+j/HUtRPKLhVXmqyodx
b+cCDpGtufnwmDhx8/3kuPBsDYcqORTRATbLhBr6GZMWhHEFYXyipP5tsTygpU4s
PdccD/L2lHmf+JKWQQ65/Q9x7bF0PnkJBrJWfWKsagt65gAWbxqRrp3aoe6ay9/p
XKZs3rVE+CxwKrGFG19bXA+jWUjqHH0LQ99rtRjQdaQswIP9Fh9nyC3cCDWwwwVb
aDHExEmZMa+OLUwk3bNOCIzmmMQkY/bk3Zo1c7/PL7B//bfWT38FQ82oHo3mXrdx
CWWc8XD7y9wjxNHSVwisydYui9/NaGDYCqx7NyFnNmCzs5gIHu0iJaqt5JRzx4cM
rQpn7hl9rgW2J9fKpoVJD6sREZCsssdIQRAeQlGfO2y8Ot2r0yYknOfgdk1cVXpe
URUYN6+m3aSjyaw4eaIOQZ5RZzZwaXkkizGlggHag5dkBHZRRKPtDj0GNhCg/NZh
kLQvXhJ08j4e5S3TFo3pqfCIE+mgb4DlgBMibjdoFHRco1c6Yce5VNFRrn22RlkR
RFaiyDCJwOIbEWnh1anZ1bZwvvDfsHcyUdqcMmmFQfomDe18Le2wKbi+eKOquii7
vtqJ36ih8MhZ/TUN3AdP94gU6BRx43im9y/JIFqVNdiZpM7Qe1AsfEZPIt3XU5vh
10n4FJ83uV+O1joPYf4Bx5BCVQYjNgaFrV9JS/1oBDODkGAUL2eItnDVx9pvxsr3
bsgSk+aoPF1i9h34D1mwPwWf857d4QHvyWvR+BP3F8F6xz9Q8ulHiFfih7Ok0izm
NEVqoDTgw88VU1HSoRdbc9yJCQkY+xiumJl4TU9Spx0wFicy7Q7vHPw711NC6g9z
9g1VqpIUqGeVlA3YU0eAsAtjD8j9SWpc+Q7owdlGKgIeik5KjSH/PdlP2wpEFi3r
6xzb/fvHWNn0ZmVKjyxAz2zFbk0WvKxvb+jk0n6EznIygiuufI6MjIb3+ugO1BMg
bG5bbsy6zkYVstbkRgTUG0q8FIawGk2BQW5MkENU3XOMUf11i34H4Pm8zJrrMyX5
xGKHsjiZYwLmiSX5POv3OvwZGEbek+THzUHZWnHBLlplpCqNAlYf1qTzxMkn4pQX
7YWmLhJ2rB16AumIAt6ycBJFU8+zz++OhArL4Yr2v6XRQH3hIQvMvDv7KsxShsCl
vGh96pBzCqd575aB4AhsDyE6sp+8a4OkymHpFotH19sMibaA9JhGz0Wth0kQdYml
GF4jERZciS9snUhicv9aYpAxxR07UBy24aq8HOztlpceYFj1dIXlJlpfcqEGW7QZ
hdiTS273i5WY22Ud+Nu9yA9w2M39Nsdwm+ZZfsk1EPYPcjt4v5WZfFnRBKjjYOGi
yAMjT8zW8i4eqDK3pfCfv9RHpisMSFMX5CX+SLrobYYKKSbY4H/ar1YIu3kEJuns
GFrDIksevMxtz+M+odSejDLs3aktrjEz9sda00YXjoxtDo6+cJanU02As3h6V6i4
MawP09AzOg4/FaysYXUiL2Y2kDNJ3YvFiQXJ045aJ+0w8+vOxncjzZOVjC4NsG4H
v6YZmhldrDZWgm1zqAZzRUxt1haH8EdYL89eCrcq2zejWGB9WJRbvbgXVOWgU76N
Sweo2RjFhBdyN3wcfDMyn8XCVRU+wqE7LzFh65DWpInceJPUiNq26Y4OhMghre4N
PYVsv2bo9sfvMu+oQZDry/d9Gt2Hw2paSAcuOb24BHbSwobU+uKYEY5xfYXDp949
oZUjzCauwVZr+q00pu9PF0Dc/aNryTZSP3XauGndztr8dNbTL9fW6wkXesHDjln3
F5cvK5MpUsUd9nENsl1XE554VOtvM/ModgR+GQXvxZbnNi65Fa3keIG7MjSPwrbP
7SZ4SHxs/nEsFX5gNuk3C357Uou8QkUstjU3itj1UAAqmacSJ4syWbFqX5oCoEuh
z+qnVFRochgUd2Sx8ctV3YFa86c6UaDD484C8kemLf6QdPvdgk30HeTdbo/fpoRl
V3fOYZh5rhy1v5SVpIDOBmMWdNuZrtyQdby6/Pzx69/gJEfHwpY/FXQiajWz77Ga
60wPwh1IVK6VuKiNHwwpIJdJazkYqScHlXL5RrtvDYs+vyexL5G+aB9omysRrimD
oN8ytPimpgbK4Giil26Bjnxe+Y1845XfcnNNOCNnziDL3lWrS8wQnxcFW67l3ZV0
EaaUrPNVdGZ/R1RCIkI+IVVGG1Gyg7d+aMKh0dGMjf0D1xVrMIsmmYpxpf9BFMs3
PrHTSOsPihEIJkP7YQioMDoN097f7ZfRynet8dZHiuo7QWQKk1n+DsM/g9++2PjJ
okTS8tw41+UIClBpTWRNTJltpUcb0b1iLGnJPMtVwZ89IXUWdeb3oDjRq9FEPWax
HCmW7d4aXjxVIpeuMp9khcBmWgcryerxmpybcDRLluEryJHeC2wLZw035FwnWdXZ
tZ73hU2Qv14FyacBlXsuzU74hRGZNkONUwRdeYquQkT1uVxLkh8Wxry50SDytK2e
L302i3EB7J5GEmRoANu+p0J+E+LJpNR/7BLU6GGFUO+FkC8V2JifgNzGFNxPg0Gh
iMJNaFx5B5rQnGcN9p6NDvucDcbf55QVslfSE5f9czw9Wdil2ROoB3cXwnaN8kRD
WqHNJnroiZMEQVCHQsjQMIyZhh1J9rbC5yTBoUY6RfAtAWtKusZ9RlAQxNxwx5rY
wuvEe3NEKhH7br5VjbRRiS+eLhPNkj2BBMwE1xpOkXjJbtPJ/NcvVjUG0DFQsu7B
pOR1qEzmPjkW+GHDiFa6RqpYHhQT8WXenFkNPPgv1peAvnN7854akrrIgfB+nNuZ
TwISyAX9kdPouZEGRyhAwrnRU0uAuJQYK+u3wSxnL+lYYGqkpZS4lbpA2FacYqde
27A0ru9z3KSCPmYob5ozuux4MwjOqFOGaloJJiPK86+IHJ+aAaRdUVU50K9hOKFn
LVwFCGd1UQn7rYH5anhB90KrVJ0QCFViXGeA7xy3kBOthi3nKDVOJ9tEHjN6Ue+x
QRlauGh+5WxOSYZk1A3NRyEV5eb/L6AJZ/1VOOpYcHDRFAnVJExJCBcHx4D7Lxay
WE2CXsttT5znUwXpWvbTqF96tzNjUMJDTfSd5mL1Gy98Wb4R3s8T4os9hpHGj1FY
tVGp4UlqdQLHCZLbefLSuGHncJLVYaTOYrrdUVnTg4HAxeJu+RF74FIQi17fqcrE
vJPZ/exlq7zSTHLdLM/qwguPLU6linhFaVA18PQK2T4964ZWBja/hcPDsONnL86j
ry4FSfGJ2ZLE0xT7Wakl5tJFFjfaKQX9cteNKaZY0dilfY16+xC87CboC7VnMIN7
JVAm3UsEYT+11J5yshbu96m4xW+Sv/BvnO+PYMzkS1qFb60EH+VE3bz86qirWRCD
g37jMJ4Uu7vBAvNOTFYIldDIMI3q7zfrYRZttuevOYPVT4MKZRCeEIkBAqDJLMjx
mGcu57ImTY5pQN64NDPz+6DbObuRKdyfKdJYwqoNO9TO54nOFEbgLvCFj94yzewK
jRDzXdREYQoXuSUXcfe40AYJEXE7Oj1Ep5Ks/3G1FiGCunBiGoeKOfY9h9qPCyRt
pOvzblfTH90E9TCYQ3L+478gsJ4QuQhsnESUxrVonotvbZxhS+SpMBA9/i5h7tc3
3qr6y9+7C16sSq/R16/ug2/VcSerVW1XIMK51qsvxejzfmTen4fosMq1E7FpWQwj
FNCBI1VtJX1g7SwaA1vWFjCgM/JAqcmu2SRcrNdfPEon5Ufr4LBvxNpi/2Sjeb4j
vlXKM+yVVXzXR7/k8X0C2lfFc5TwHybTrs2eiUu6MjWFOjoqCOCcSKuAIHm5fFni
6eFCZW2k/Bd+WkWxppOPeO1n7GJ/VodJ61Br4oxU/ZV0qO0UZB5Ef2ecPi6qGyrh
ukE41UVLk0o9DQvYI7m7JsCNwx8/tx0Jkr+L0gjYugTAIQZ1qbQuq9yXjgPEJvfN
HHT8cOqJZKivaFH7tEz9G9HHwOgrRMrqqdAUbLb4CAWV7uCjzOOBrhaVtydppDv0
p9R8t9XuobRABxrX2o4aVQK8Gqa/xoOnRU+DsQq/QvX8pns+ixIADwxikt6NAG1O
Qa0ITGeUKhQcg4n5TYpxheaz3ffVP+gEGT4zrbWIc5lmpaQDDwnW4h0/vJOVQIx9
x5Vp334gM2LQyXLnuvOC62wgsj7n4T6U4On5PQuFF2RW0lIJukIekLNSluPb+xhd
dln60IlYVTG1ol6SgY1GmsmLcInAXL03TQAGxCKWfvzAsjTjiy5uEYCRmJdpD+xG
YEJvMH3ePTIxacnolimZvbUomSo2J93SQrC/8FUqnr1stA8CkiSIaP4T7Qdj/EIJ
GCFjX3fEhPAZQHlrMQyYp+0MbYVZypY9ViDDExwtt0nB0Ng8a1NmZVpadOEP0F6R
AdSPuJRNHLfuf/B6TSlEiuHClfENofQDgKdSGLMJCVrN6UUP5EbeKW6WWelM6ZE9
dF9KiOZF6WqQnYeVQAniUB8ql5Y2OQLm646aIB3urFduJq3ddnTni6UpDeXACUoN
YdcfzwlEl3hQh2e0lounRiik1kIhcMIG4sxiM1B5IsRlZLluDA905CRtBYg0ns+6
1vbbcZx8dAwIxwWfooSQNWUpOz0snqYMm44dhb0TZq6RylRU1Bs1DmGbFRKBCPCj
PSirIDnwDVB8HQ25uvDrC1uk/gILGKViv723ppkgsvKpKhyyNw0IS5OebLK9Cr4w
3r5k8zECnpH8yLgsNXzZATYq+vWZJJYkr18+pc+wzBcjEIuLScEIeZkwxnZ+YkSk
c5msl41utiQQOFbi2NwIKmQY2EvfS28mkHUaBXJiH0s9cGTqJAV1+xaJSlQgBuG9
Ug4T0hFumytAUbEvNfaVAs1eBo7UxWT/WSsFb33n4FrKbw0GNT06ai8961E4WFAs
VOG1chfUVuVtJEKKe6++TiZu1CAVSB8iuWGQy/AGZd2nuo1yhevueNlGfe1yy3at
9QXv8opM+lJK8pP2BNvjsuudRRnCEotq3PASuQ/hdbeT84tr32JUwG4aDGq8Cugb
kJKHRG+krHLlZnri603OKxHhSqHCvmThPnudV2Dvqf7nzw1WKS90kn+DYZgrfmdS
9IjBpLdHvX7rkcB6OMM2a6krXGay0pXQa+wWI6Wj0xuhxKa77M3p3YS90Ym58hA4
+Vx6KfFnwjlJKmHqvty0KZ3bq4tmt2lWvYRpbZwZ0y8BeeYh0+1CyFRs/Ze5yYt0
UlD17T7mvwzJYQSYvDaDiNBjf6CfkwlcFtrxrb8sKbO7LipqX4ud1zNDpl7dRVRd
r6ErtS+2us5nSyf3SltP53n9JZ15pZb4EX8aH5wBet4sObmqpvfLV0opLMQS0G5x
uIj3UemjwoCXRa7sihbC4d+SidhXb562mdZvcpbwb7n1dlMsrdoVtOTm0+HdvdAx
mf0d9GmPoFQ1dX9HNMBvNyzmO8Dyjcz2iIUhFtZdvkvEtcyIDbEvBJLAqZ97IM27
rudABoZ5CUwrjsdE3IbHF6l+5dNiw3CTsHcY19kMenIJ0C12f4w1q3fqtK8RXARx
m0Y/p5u2kN/n31zqu6CP/RbEg/vRf3/ofIjFddm2d8ponSYcaHIuijwADEc5/odS
WWXiiovf62VhxDEKpU79ddbwhiiKZpIqfN7RC8MtrBf0yCv06ipOMqZPj0PmxHFy
8oS8n3OOWyHdX6+qvRL8rtVkNTispjd4yEalnaPPzh9XFZeGnbYmdxH4azb+jHRg
vmfHwqGjHGOnQwcGLC/FhhPKSv2lBtf11RUY14GMbSVMlXXt6HX6GbgWFndJVszT
UHRLJo/5h4hf/AidiBssLItRBoYLs88Ld8PBqIv86uC03emVplJbHn+1odGOB86R
axjtk2DSJMkyXPha3k7kEv2Z3YU6+MCwfmC0+P84mVCzZhEOWnMsdLyCHkKzf4PT
d4nG4AjFmzHxnyp9ylKpAGbylOP2l+hGZJWwPdM1VgtltEwZmPIAC7aTcKQyqmf4
ntG01fWK4OEIp1ILueKZ+sxhOgXCdDHQvNjxx/rAJO+l2H1ShqgbwfcHEiwnuWnH
MdJH+1lnDwGrWuMFXIWwWX/HxLo6YHjlKARZ/WNkv+5iJ5da8NMFQT7cPNi1KofK
sAfL/gBUDiu5K+z4cE/viDSK8qGqd5Zs4k6dBprb+wr2OKd48jExNSjw1W9bxkxB
nZcylx7DiKG9LYWNqXQRQPoUYVBQOfnwXYFLNOpI1NTmA3kWNVMquVLmwviOMvhn
ailKg8O+y48pfD8ooWKxYk/47fBVNTFPbGvn9Ct0p5kLCgTwT8bMOmWMHDZCpgOd
PO/e8qiEd+wYZahCrTT6bqTSYi6H303wdnl4yC3qfDjkB5yXD3/aT77ZL7wacvxk
XvlRRcWcrfAyXtHdECvJ0D0TrvI/R8rZtkPFGErp2dXgyQSNmJcQnmv+eZdiuBeV
PotKGtD8x1QhJF3AntLCFF5s/tK5zYU4aowm6BVe2Eqhv+RHbl9KRFuYkeHcrw4g
UVw4o/wOntJu4ivAOSfyXNi71g/epYEC3j2WRMjdfu9Rvh76ExVBTRU6MM9bRAu0
rwYrWS03tgY1yApXhiCU1KKU+jElYDwOCKPCliU4S9Yx+xILlfuvy8j6r7emsgPK
9/mRKwGyWVnRKLRKEtvKlW217GcopAop5mobWXxB+FP0vrh3ynHs9D8QaJ2C/Cb9
/dmh1oTac3exd2KwLlVa9btxDLZY2fi8CZCEoA4dB6bjbAn1+99DhmWzjLkC/CkT
HhuCHlWHA4nrvHaFyQiJ/NqOYSijDUpJK5bHzW4iicd+RuLlrz99kXk8tu+ixBeY
3xkgTze/k6RkYgPEEb6n2uz/ygCdgSntU3cR4HE7+biHX5fmZJpOagzs/PmtzjTE
QanqQ2MAAYG/MyrufK76u3OM6ShQL08mkZOy9BtdoL1cV5sqJi+0yJQrILrKMI+F
3hw/qBSvjW9GOvHJf8u2Cw3rBrTPQaApS0fVc0R7DzR+JUWX2TSxtw+9HvYEQl2O
JsyvsUc1L9G4VQvZrsk5svkV/+TSgtC+vonkKxDPo4h1yteyvBYGkNeDn0QmqJAT
f1Ybq7wbHW2ywjmYD5UiZMb4tQraGs0s6k6sz5nG1ZlFCLriIgN9b+oTli6cmgtO
Ef/7Q05TKDuDkSyG5BBUZZmm2GtITBAz6Tlr2CvmjM0fSltrv4bnEscevRh4F5yF
DSxgqxi0FXA6JRb0kkPgu+7hXIpdTn5dt0UcljOIzaYbWvi0uzmGr5yFenlIHZ+j
G913oSbYovkj89oNlZWxQw7h+HvuTxiDEoVxr10a35lmPH9e5UAUzWNPSr9iu7wr
4l9D81ExzfjLOAZq/tAs3xxL9fm03IyQGJiMV6BLcO0H/S4+n+PjR+9QcMLrRHUD
Vk7uIIlkWyB09EjweayAkOHJUQB1zVBE6dJZKACsVvFKFDHdsLa7xzbDdKG1ZAii
jWIrW1Lgxx/BhYEBH25prArgi2b4wIF7bZgyjmdtS2K7oqd0NWZdy8u2hqqp8clm
9aWlAZ66aztpUhO/i3ciVDm76A+JXXmgrnTru4OCJtSSTQAozI92lT0Jp2dlasXO
LYVNDW/b+IAPpAVFLFIMgmggwddR4Bca/XOzcTE1d6wMMQtW41D5ogPEIe5Eu/U/
H2l6aRMMxOG4hUAc23SJCZhA9MCJ7xId/ozAwdMH1M/5J+2ZCxNk/3+WG+UN5fnV
VLllZqC06JYnhTC0+Kzaofj06UTmYMX+eV764ZNedV5l2AJb/6Lrm8y1OrePGRIs
Pn1G/8X6Fxps8C0odXsPZOU4DmN8jbWxGKXHgUsRONdTCa8ZLQJ5ioeHMCpvYIe9
JEd+sMUA4ovdd9WmLcAh8gFAk6guuhqbd9rZSXZ4/QMA6a1Q+WOTtc5IrifL/Sd6
qhLSUmTddFnOuPA11zinpKzc6tEqXibEmjgLghiU+LZA+HIX5ww57EYlQ+hNrTH8
gLn4xX0IH8mS2qTy5ULeadViRW0U854/S5S+AZCgCAfLFtFeZHogADUlOtGeE1mR
bzkW7p70PRYkeg9ger6hblmHIAr/S5EA6OvYUJsmbOGvQdW8vxZNUVctHGbCj4OB
dyXzqRuYAIAbCtaEixy6sr2bv9a2VtxSR4XjD3auynId7taXfQPg0urdywQIVLta
QWFV4m5I8D6tD9rn99hGTcPJznUvro/rASgvnZMYBPA/B/u8CBQvSto+CY+DCI7/
bQ9fvO+PRCGZcWGwbMpadi7jAJjPHRkjTlSf00fWsop8/f6N5XYFlsh+lpVGQUSm
psJu4CA7mYIdLRhdo9n33dKv9Gt189Pqi5Oqz+m6MIXstY5oVmBPjv9gQ11tJz2Y
w7YJ0TAYS6c59Gg1eMHIKYlPuZIl69vnFapgMSL9vLGwC/z5Lp4dXa/mhURiu8C5
vsU33CJqPiXxWtTWJPNP5Go/CW39P6PGv2vjvZqlrH61g6gzzKKZdiqJdTjwZ7Gy
OX82GL7doEB29/P4AXG6NW+tcYROEXEpFJ3TCWvILyjZv4VmDUYp0/T1u2f0ZjEr
o9evFyiCjXfcfuTHik/v0skgGQsV5YkCfrghzMFuXZNpgDH24pKs4aEIfv5Mk/gm
sLwxl7XYKX0dpvufBtcwLcM/yhS9OXS/r+/cQzwzAHd95IIxrnarDB/NoJKJGI1t
eZzt87EDjlbXpeIQFOodb0wYTi264ZUS5HOS/nxvtnou1OB9/FFOZcdPtbPAEiDT
uwyUNdAe+B3H7pUgw7weytLVYIH++sgyzbQs6NRpgHGkR38lGSy4sKmsKZO3m3nF
jRDdYbZOc+yVpUrv21TaKlvmBIC9RENNkAtGdDiEsh9BmdvMvZg3ZVTkue0K3fWL
nPsQ80xUOT8T+ttaBSnWeo6hYDqHcfhMbRFH61QhpSbyXM68a0mpBngz83dzLfeS
dY/6priuBn5ybmYt51CC76U2lmiX9acPBKOO8FF+W8k0eeEXL/PpGkJNHDE9Mfdy
YIHB1ScliHXkpIykeWIMxFlrjkPAYloaWwg+VyPHs+zTHEM5NzeeqQJBZ6szHeaa
lca9Y4P8T19PXACJ4Gk+ButbiyN8LjU4gPo5i1dNnLCEKDzuhftt8iOudsaU8q2z
iFvKsGP+axdtfrpWyU1MV2mvysC9gXzfB0psvrMKogWSOfrxuDs6hyt2/NBQnE0N
4QuldsN1yhEIEbDhbEcRBF1DnGCxW5D6d3uEwSQqU16PheQ0uAZBWirPaJVrEuZc
ZiISL/nD5OVLCQ3iqfZkWdmAiGQKXi7hWqrzXIv0fPC6uCvN85BgoFEEEKygBK+Z
lkI+hzQ6V7N0TZjLauJWIe1rHNDmaILMGgUelPdzdwR/oA5JGeODKSim6bgPjQGz
vj6X7Z0aR9oCC5+p4beOz4fNY/75GTwAkMBRJEH8u1O9KdDo/8YWjkkTxEcK9aN8
/2bi37OBzaWliPdqLId7LQ44q2b5/Chg9TMnO5KnM741sBzaUEXYxBhWixc9VMD8
XS4nHkZs2yOkFHK+iW8LiJ7FdTzPLRwMaYxoDZ1WV1Q0MhVZjFBZf93HAPiJNFQk
n/hbrHlb1zO2QuigtCM86q00bbqOUVDUMCemt9tqmh9Utz54vlcH1baQWB3Q8a11
CW/m31bLKvsMeWIA0epSqpCRuMo2SDw1wXHevUkdXTk3yX+e3raXHz0ik1PPqEem
iR0teewbYG7uruwGR7KzA2P/5l4xrpffomnpZ39O7pzMAj1b1ctJaC1WS/pUYWEh
1pFk/15C9M721/sNSnEZcJX2iUwAfvKYa88vmmR9DQLqnrJWZHRw+vqYfSH599L2
JLVB8s83oH2wpNAp1Vdw6VWUkP8Cu0wEB7TjeCMruNS/7huLHp5fQctNL4jYW2Tc
viSF4EncdZYTOcrz08qu74PMTEJKDMDmpoanOM9qPkyGaEZS3hktYPYnHSWL1U0s
Pyf2Wsjs3KCVYR1iVRKp67ENxNxoofesvMPIyqsW5ZLgxSfwPYRl3+ahOzMMXSLR
kFLqvdpkTfyg16bHfhQo9CWR8NC+dfi/A2FkDnxddQ9BI9nY2wlu26xWaG6XLVfr
HuSNug97Z7NRnEN+65q+bInZ2qwneXJxb/M/IApn4CmoWiZFQ8voIQzWdaCyknTK
+u+jlG9dpnHiqVvbK720OqXiMT71Vv4TQtWGGoluOCKyS+Bv9EXAiaKCXN1VYm5g
W/q2FCl80FT0pUX+nvID/zjHt5I2NZ0Oy1/j2QYPht4ysHTckigF75sMxiOBRt+W
ekxokSYbDejsiBGAVSpgT/ZoTx4/p2TIpKbxOD5mpdI5djggJel63T+/Rj9OJCY6
foGGksme7GGlgO4Vk/skivVb8+sTFotQwJTeTixADyzZtmzUrw3o6EB2H7fnwDY0
waenSXRTbatdjxNSKJmMGlLqekItOxufceDpKEHq8IaVqNlzliJnRZUoaf8HN5uV
zWmkOrZ1ITMr86PET0kUUeQSwoLLKEkeJcRIRcSexSbvTxqYq/T6YaZAHJcG1hTp
Zgw7BFWI5twtZOB2DPTd2ZF3ufhYZg39+DSNT2G5c1iaFKcgWaQm1LiV4I/3mQxf
4kY0KJp5WkzVeJacPRyZGSncYkkJ6ha4BURivVjT/evR5szGGmYAsGQr1wpykWlH
3rf3P49isT/W1UTDNI12Shu47ax67Ct1KyHtBW8rKUMLVwf7Pdm94zB0pJB36qPe
vgAeVE9FBJX995Nlej6QO68gCOWp1ixjQ+3LMeV+iGqXgFnq0vI/1N+dn5NBBEW8
vs7qwieW3MRPFdKwToAEIoEWp0ibAAFYS0q7VdaolbumwlOw9wLBMzVZcCjaozvg
+HkdslxYSRRLWIHk19n+Vsg0egqxPQyFxHut/L9pdPqXw5VSSCoLAyDJC+EP4Ej9
y5OoYDk2LfJRM9SiAygsvFLhwZ9yocE1dIwzQIgTDt+9CyIWZMUeqExyeS8lF5h1
S0wfL+/qYPJiqXkO+P3ZHDoM4k8sGLL52Ig/P1aLdMciGDH87DJUeG+7br5ULw4q
jjKHtf36EzJpSKpnrTyASfQuOqKLECyK0h7WuOPMxgPSTW+k6UEAt1o7eLZfeHff
sCDnpCB3gPMLKf/njcYwwdqDRcdaYcy/Up+PKmspr8NZTVyQt0LLY7V26cZs7iNV
Aib+mO9Oj95uZAx2sOv/d2lzmUVDClaZQ+yEw2yy/7u/6QhHA23n1sBq8Vdt63Wm
UO4E2Z1SZPOMZYqF+n+K1e/dyCvGKxSJQ/8Wq/DOduGU5fkPNzk5/L5eYibMIXTA
Nz+759So0OHdnXRKUiwWN90pyqA3H0X81LYW6KHWNdYo9fQzUttehzNuHGN6PCD1
g4n2uLMgXecdS9YyB9KlpEEWbAzCqowcMc8ZmONKmSYRThYT4Mav1m9ibOnnHFJn
3rE5mw2n9RzI7me5i0v/xe6wzzplKtW+41er1ZPaMbe4m9WXPxi/pb2dKemJVmuI
r0wC0ChhlTr06AE3mCR55/uSlDOcRM34X9doU/SDl3EcUJ5PVmO+Z8LkhtKA6gKW
QOJKu3whh9GtporbRbiH3FrCDTDieHsitI/zSh7cq6QcJHRS3aA9OdhHz4GRWoT5
+JRdHaj6mEfVptJcAYCn5xEbr9+ru7WdPdNL9Oy4NYRcmaZy1WLGjiNn5eEZxXwE
VeNTT3R+yNRQzGEDk58OGxvO9kJcoiQ70qgOfOui2j80aDr8XbqwWGPt7oRko1/s
qs2DGji6SnAQBTjdyiRFqHKPSjyuEO9mnACJlqMvYuV+JJSTJzr5k5PWW48I2YjI
jSmEMgBfI+21rIPzaTX+FyLY2Ld0beIybqqlMHY6wvGP22VQ6Cq1ZyVReSXAzyvJ
9GNYe89dp/V4KNXQpduhiJdqHWAKKehvDsyFLJEZfdOFUId7EdHLMIdegQT8t+s5
ttUuAZU0sX/BqyIjlemwfY1zk/iZD6OgRBi5CV5An285rGCNNAfrEHwoYjifVENz
94zQNOZ/l3nLzsLU29wNbD90IytbohcN3AISK+fo/Hu/W/oKL/P0HoUq8bmHKg5M
gxWnljl4NtvH2xzkYuIlkjpf6jmckUVvLnwjJXtWNw3ZQg6DiOA2s8OrN9ivToea
R0w0xiCSUEan1Idq8JgQBjFilK2uGO1aXGt8UfajwwX+sEB3jjucIAsf33vECxlA
hLe1kIZG52Q+cma86Q3GvHkgYoTYSNNhQkLgmpyNODq+aYuQzZyLpAfWfnsOLZin
f+Zrv1J3VIfLou01j+/vIw8BB1NHiYWavjCGyXas5hj3uk7Qh63e+aSM3VuXJ2w6
1fdVKW2IkElfcPp/l9NiUC9k4Ch6w1cGzQU7Fs1VqVqXc27PX/Y56BSKQ0bE8X6L
BGEEvaFKrMWgt/onOxnr34zK7iQspXhwsQkzFFjaKLeNB7lGxgsLLgvdPKklGTw1
OvAvfimZtWVKdEmobIwLf8tjI7Ce4z4OyZrM6LIxmtb58T08G7lm/Xv7xckuMLRO
hmH4UPTyEZpXvFhZFtdKcJznvlVm5AP0qWainwo1KM0HGa+xPCq4eAYFb1uaZBsT
vkzwMbnDn4JV5GB4rt/5tksjpK6XSY3/nRevGir/47QVo/9lNnlrcpTLwlSawJyt
zWy5MmTPYgqZbEpaM8hOfXI42XuiDJujRGJLgyM6o1a/9kzg7imIfl/FIUbcpTol
mzY7YdCw1BA8SVpBSEL1ML5iPyN/X7YaiPWsXcwkb7Sqn8Ong+Lu86uaC45M805K
9VaIx2SKqYT0HBzA31Pr5r3WwaCV+8z58QrGD9dSsiuP1kjawaLZRC0yGhyQAcWr
IvXZZriwIaMqXJb8blTQ8olXCKewqQdqdtxXdyDhxQgHcDXF0NzwRXkraKOSGi/0
CynpeVab6/05eN0v74G7/qRwvyMLKY+k/Y9odpUhmEtEnhzR/GhWS1y0GhbCZpWt
K5GPKdO64Ih57OXwqyg/3JgATRZkNanJYLFGFHTS+ZzMr66FD1ZOhn/2PDOlF8XV
WKa0Ar3MWK4YiHWMHhNMCxulLiupQRRqMZJRM9qavGClTLm2M9kfVhqwKa8sqsv+
qrd14d1UZfef6nKMpVwLv7jtDUWM0C3pScApnSOtjxuNaT81/w9vN2KcqVCnY610
HTkFKjqXRO6TnLky+/dz4CuDrhUJ31djJOOXR1+VS4C9g5UxM8kWXseqFBvX6JbP
emrkL9mExs0imphB3RUuNWNZMJcyrvDKM3bJM4SH7Qhc2bI6rbE/EwXpYJaBrQVE
9pl6nrDtPw/7ftwwWPfCAfhTJ5Rr6lgPbkDJuPW4bqgZQ0+Tq5w6ehRflYgIQRry
XV0O7mphfSqtr/SAwWqHrPi6NuK4G1DlgSt6ngtFSHmoq+/xe19m+0a3ku89od9u
4ce6KBR8YSdF3CHBArpoOxG3Oeqrxm3v5UMxSO1ewTztTEFNQrvnwg/Tf0ysiMTX
z7K47gT4wJ4fIwZF6aP7N4i6otULDdKX1TeM8Bhu8U/J3g1vKtXMeWMnon4fEyaX
gtYaY4McGT3WHvwm/MiPpKmpQSv+SmppwNZbvlvApElxtcGqwxPJ/oNgycSV17Sg
8XhJqliz8bVstocWlGQL9RHES6Qf+t1f1q0CJBDet4VrQeIe8MFYjad/yzBbyiZO
BNtPmvAIR5N/iRZBSwt7EjeorNZ2Nhus1PbWQYT+MP/EktMcgzTOP9VfuDjOf0LO
AsOUdY781LfuefK+UIl1bX4kkHQ4aSwCvUjSRuafPTe0QvMzj4y/78C2y9fWq/TT
C6PDAmFprgs3cpHNog3xa4Q1oUyXaI+N/fwDL2f/K4I5deF7Z+85DnGSVI1sJNyX
hiQxxaxmaua1QGNfJHifXLgNtBo7HF63m2L87FKKeY6+0BZMmE8TuFKyJLqrJ0p+
w/K4EyPPPj9C+Ekyv4eczvnqpKo7nBKdKJWMGrX6sBPk2Im2+wxz639bdYMABhz0
kQBuP0uB41pwQO6kku0UarG145wBHYvVsQgOCrMr26x8Ec7pK177XrRCTtafmJts
mSSCVrjVfBh+m2kog/3fojTIDB0J1JcpkYOko7b/dPwgcG8xGFRThVBZt1kI4gXS
GXucIPzzDwPxiRChcwGUtCzSY4RmT/Frq+2vGrxyes/c0upB242QcCK1TQ0LN735
qs1vqMTZNVcWXciWMTcrh4iSNbsT0SIfyfjICfu6DwvY7tBS614fuD+7ezF6ehaa
/jq6IP6hmh2aKd9KGio1kkfJyfe14Q1h0q/DkqG3vxn3bO+eiNLt2J7JqMOLqEgw
D4/ccoznlKHXznT0PWG3dk82bPo7jXpJRFE7MBG5lnPMKykg95rD/FDaHx0c+Nbe
flvAyWvMyIA6ujQNO6jrCW9rA8ZnRZmLVMmp4ZWeoT35vuIdkiyElsiEqNPFl50j
VqeAtnTWZMDWTETIJ82xsga7G5JM//9et61icAR8wAnPACiyWw+/4NoIZfXU4juf
CxxI8MPGLRMHUwING8mxJg2Ggjv0t0zAYn9VCQ++Pkq2vC8XSVOApi8y24gMjBVa
oZq3ty01XqizVOxIy39NPjfmX+wuajygLzqPaIyECKqAeSJ6ZtXz+YILI7BIX+YR
nDq2lyOseCeJKvhauSq5HTB1NE/fcOvBM0oLvKFS8C3UWNHfEP5SNvgn/qOPlkgL
jKIINA1G+Fe3nLEyczvOjEkHGPrQOXtQZImgKD12K1Ada0OMjwy1wzTFfxDFgwxk
2uCu3YESwzuDqCB4f5cQFmgys2TBGn//euNdFbkf4+EE8qoewVl7EWU7UqOAcukj
Oa8TLUMcvKv3CtW5zBhH2dhtwVfcntywoPeWlYOY7xvgu8jZz4apNwk/EnGbVC3M
PfcV+/g28yr5P/Orou1z4hkXSmaz7dKiGQXOkS/FxFzOt79ZOWUbuoMSPmykfHsa
0tTAcD7J3Ysv4/Yxe7gGEvdQCOnPUBy2KSWB9CyevtLuLB7xef0b/2OMTug4tavF
8Rw0B+1pRCRvv0A6f3mvIPNCSzd44Ey3ddIY4EIjzBCuSqENW7Q5tkgk6muPCXAw
HrFcFSjQ+9LnbQL3G5cPz/F/ejZ3FwSQ0wlNzBzUAw/P82/WtPcYAINl5s4CViAW
FuiNxVDPdJEta3HGRfJW79ETZ3X2a//I4espVL7EKIfYX/HgVLiGGcYjur/v/VZ/
WY2LE3BU0PGq8f3nmMXosuMQaK8aYa50BMhLOWHW/wYAGKutM1j71P2EqbPZ6Aki
pQ8QOXjXos1hLcdo7UZOAefR2Yv6w2XSYgPAwnpKQ8NrLMYi5c6AoGA7eE3XKRtV
faljn4Gvo1JfKvVEoMuC2wE1cKQs6xVn+JrrNxgE33fsI1iwypD210Yvs/VUrhS8
034ncFK1Mn93EkOgFmYOj8g6Abd0D4yXPW3A4ILF7suRighlBMBDEiERLFDB6v+W
7v3jxFBfungjS/aoraDEZA09AaH5TABuLqvnPSlvVBX5kRdxSncoIeBeeppyjLiu
myAGLLAFnEdwNlsSMPCOA/pnkPA6ySC7eutW2PrSYb36lu1IZx5iE2YNsJdTbseG
lYU8izg9t5qp0SjI1NGeNXZlH0iPNMKxBP5Xq1wtU4WM4FAsIZNiGhF/m21GBS/T
hoPuc8O1KsjpQCsdOv9mH5Jvd5RE1faXyxR2U9Vcr677APAHIH5ISz8+mptInUxv
V2nV1kaEzmV/rbPBUw03+636dXiW572xhKzW7CiJTnYeHM3xkLI+MEG6VawniTl4
e17SjSxMTqxVXo1frIiBAcaUPH1EtN8ObPg9ZwHfyc0q6pogmlUqzGTw2RJwBofW
PzgJ8ESVSFXlRUwD72z4bv39CynQChKUJ5/BlZaHW0c/s2yYvdvXgjHLIJDebRV5
8/Iv5QtUXt0f36BaFT3iccHUrXjOYNEvXgKWNi2auAKK/Yiu3AZSW6Fc+foF6Fbe
b0iepMdFF3b/VMb5TLaa4KZv+i2yJfAqh36RL59XJfW9lEVDIDm52s6UGfx83jhk
3RQbYNCJitaYYBO+udwuXvDZRT/cH458tVFxTMzwMcYaQUukdNhLM5aEHf09kU/Y
5a9s8LECXfdM11EcFqU0FaZnLI2lsv6wzntG283QYs9suGCfF/MTLglUJFGcET+Y
E00RhG2rYu4iCyWhCs57pz9GHHnCeIGX6g+wnYjFkzL7DEc1ZewD3umqdPze/X6H
dJT3tnQ6GNiYRcW+yYJZ1qKKi9ExinHRoosIDbGGcgyKx1mN9L5zUjSzhMkEEr+U
mql1TyaIhWaC3+fxi5nxX9iworakZzRsv8X/NzeLua3TEBG8DHtRFkbPE48nm1WG
zOGc2jCnaF9H4uGqHlb4z/8Xqyw/bwnLT0lDfiThgq0He5STejzv3S60RT64tpYT
DDxE+TXT8BFhi2AIMzyCfLf9ZTO3C/lguFR3k4ZOnwNDLX6bD5iFMgEUiPey9N5r
G/EYjn4YwgKJBgARPhkCJ2F8c8kakIlID7UbFrfPc7FcfVq+zdrzemo7nL/w/Tif
fJ1q4J1E6FXp1OZBNTollQg4UK+kplDII+SOmlztWjdChcL5o+gaD0FqNc8REAoi
w1Rr2Is2PBIPu+3PfWueOlbB78eiFrad7GbzzVQaS9EKS3nBc8nsGdQ8CJ0BRhB0
Ml7REy8cuPbh5eB0U/cZbLyBoJoGZDGM6545WoFdt4TNuAfjbG8OzjRps+ddbJWp
+0QKtw/023a6I3AXxChGKuLL+ubnYZ6/ZNZ1zLqi+OvSFBbQASBA6GPo68D5glko
yPuqaXSePVRKax4B4Sqyi5VN5l9IEoysEENuhw5Lt0v6DutXHvIWVWRwQoDYAxm/
Nom2BT4Qd+SO9kbLm/jWIFTvZts7zbBgQueXwNtj2hKYbrvqJxDSJ6ZeghkZu8BA
qjnTEcd8lxj/Rj91i3fVvXjB9XCdhYEKZwNIcz22rA/G5GVHIr+tiydEjBDMC4wv
DP2py1c33TAWiuhKH+mTWi/cjt/1Z8UDkaOHeZR0RCH7LW61/DROIIo+JV3bn2Hs
xHt1bXZljNBPPK5kT/8bjfSWGz6wvcACiywoeFmtIGINDoPaTGuv1vL9gUhVcjJ2
QUoQIMkDY5/owmZ0lDuHIfzUHlfVUTYoiTOB90MRvgdmr7SW/eoj22/OySswBNFw
H6hOGrYuPGxSJS8EkG0BY9mB6OUiPVwfrywasj+6/1nV0RDNVxm1y1sSQZfUS93B
cDmPiCDA2PsKwxiJS5X4USIL/S2lWWU4hxYKWvVD2H80sE1yQWJ20h+6EP7FOllc
uVE95dnt+4zIiWZ1cA4koRmYP2KfaaZVyoubere/5LICJZpkQlqQ1NLF/fFJ1q12
3Q6y6bajNwvF8QR36nLFbqGALu1OKzWzCqesY5AvQW6M4LUa4+G7h9mtxmNUdPpo
RU7pfxfNcPLMBwvKmwFSclWlJpTNFsaxdU7GwqnyNVCUDk0A+cRBC5efWTN31YDI
dZyr/YZfKeS1Kshy2hTXSbX51+xHUS69iEIMreYiO7a2G5Y6MJKIXALSEHjQ+1lk
asEctmQWJ/w40AdL52P4dSctQfgA9496QzOplRY44A1+ACsSAj4q284Q1Zse6QrL
GZedwhe+NN7/a/fXlehnKFBVthc9NyVmU4X9LrU35/ZoiKqMezyZYOatDQpVeS4z
9qnBXcIadUBaBzBklVnSMJOBWGDV0oa+u7g0MG0K4mRrIkMakEf7OFLC598En+V7
5aOGRFNGFtbePxjXlyh5JOrCOO8ehPTwrgECeRAoW/FlY1s4NgY/wugxIa0VaTbS
tzLkF1Dye+4UJrFLiQyfoVY90SRQDQs8coXIcz/RgxwKNupIpTzaOjTzi5GqOt0E
ciTH4gYjgBLjGONejfonHGVjZI13iMma1B8egR4XXvZ6y/x0oi1W2IQ9gdUa+DiK
mm6e+Xa5QgyDAqVjaVV6Alt3CZTk+8PFrVwaZA7HwrxiA1wPce2kqIiQ+tKA7udw
sbeLqwSPbFK/+uYgxn0rndy2YipRhLvsYMFEbdlsk31LU8lfaYSZVHH2i2ZjyMaq
amU32YsJ/kGcxNqUGRUIDI4QS1TW45kPjfpii5BoA5+qbRq2yOUh+JlR1mwnhB6q
Sgp5YGJbq7WnaDiPgcew3DxY7UF/BZEaEekdwvhLEXeqj0csrsl7c+bs+QeNhdkS
rkzqB0yZN347uh0+lzifT8mT2tFO4TyaaKCJz/G8TAxHNLyOQdu7QYfsuqDNBLLa
AgfO3i0wI6kbbuwcY7CTe7jFrjafC7/wTDVQ+YynSWGUqzVPMMlQNNxpsBRLtAKj
89Hwps4CNWje142BDpY2Y2cglNsWpMT3KOhA27Ikbb9JjYZy4BYe3IurJB01wGq+
WoncaC/FOw7rUQQaTtjz7i9bLAskRJEUx4CQBaITQYb8w6yVj6EaLQGEdI5f38eM
sKvFGLw9vCKa5TFTn5+V0drFOWLTNNcT2Y2GzLU50ngh+EcvC0/dN8u9T4dLSvdr
eLIu1kmb4WP4SYuTlu3t2wXYr1qgKm0z3dkIsFfObijbzgcSTWd1M3yj0mow49A1
z1hYzwopmfIsPBxtsvZS+BuEZOcVSg7MOSYUz7wRScR9SjvB2scYsUypXf1LiMmO
W0y8QanofiKrvwuhRl194ccSDht6KTAXSd5N0b5w0Z1KacHQIgQyi0MneFAbFa0U
6tCr4xyuWoox714Il6aV3w1C9qeYRAHfingS4waOfvLlgBjOrW9PK+VSpiAwVoxN
s7EiXaG5CcbHzB41X5Qqumb+KoqE4XElropsyYQX4rbphisQb480u1H9K0USvrAN
3VZtKbWAgChFdE+OUkmi+ZsXbtVQGRMl18W/hBHdyfyF+RjSOQHQUFKlnK/j3uA+
fWLYdNtnSLPsYFwuH3+oTtkWYffqEwX/KyUY8hJzxkVhI3NfIX+bggd1cppEoefz
rnNWlE1Od9ImxaToB8zi9RPeUfrOmNFXT3SoKEstnAd4mXF6xsIwQR3Ikcvj3q7z
KVrBzsQ6YkRm0NSW3zYdFonxRl27dX6iff3vPdWS7k/mpC2Sz/ZkIjioYPkvAslA
1xo1z6W4vyblFYaF5GUVMZXRaByy6C/Na0oKocUaR1dx64g29WVOjiRHj15qyrj8
DSVbZO9WgYX6NOhPiOczuSSma7DIvIrXJETcfAC9+4COCSoYBV/8ODblaU2hbChn
kc7DZ8cjZGEeZK4Xvd69wOh9qMijJI4FiaUURytAq00ffDmLLwWLzvkSTSbOUH0b
SkZIGQr/I6O3GNVw4IXKAEEbIgRpSo+HuqgYWq6MIxwtYmk5RUbcLmWNL7Id4UOo
yE4tYKyspySmniJmH1FiKisyhY0lWK7umU+g/b26+VMKU0DoFTO3+M95nK/FMQOg
OMkZFuUQ7BdvvHxhOXic2b+L78V723u+iqjNoZTG8JOWFI9rYp7y2Zvmmqib1bz1
1EqkiZP8decFXzQccwfG+W0c2Mblk8RMJwYoajve/cUXR5SkkQo/sNh/MUcoafUe
cFJDApjdWZphIkKsX3+hDSwb2fLaCyJsS/iTbAyiF/O+r8QxU+dZFvsPKVEUc6s1
03XPDwxwHkxGjEuAqmzxn/UMTWAmKEgG0//Lbr15zw0WWb7VFeZupOJZtCaWYznq
eVCUVpW5qjGb8fovEUJVJINlbx6Fl5QRFS59Daw8hKCUW/E7UfKlE9R35rbN3fBC
/dB2IjFSjQF9WSJwB49bjox6E3IjHB/1FjNRcFWOQB/PMJKrwqh64XYVak8Mx9P2
Oj4+4v61T7wWynHlRg509xjU4Z1dTLuvmQ3ysXhQYWZhRw11sFZl//2ZBkCVngVc
dsdt0JhefeXu10fahgHi6oA++AfPjMLqjgh3xAU7PZsqH1Z3ztnDJLHsOw8jyo4C
/MSxPwiH5fcvCWwPw6qeN/AJ4RHRGnWRsa4SUAPiZRBOrppO1BfBlRPBS0uQ2VJv
xI7SshozlKG98OORLcserKfTvR3livkndVZsuZ4iPsoorJyPZIuNKUwBTS2uXhVU
ZuDc4AxGhJU0CFD5uBtFYxo1u5usCPnI9FkkVGDhYM0ls/jab4YnHi67EBVyn40z
CBN1cBtpSqxcsRsfs2VyJdsltLIvfBMTzYVvkkDQZbRID82Is5MjYHr8BI99cN/A
WqqzXP5gFncPeMT5mwZaGBzqXAMbwLqKmr4gnHakrCZlg7LOHNJYqHFixRneHzUu
BhYQASmwt62hZrk2ktuLGhK8zLG8uapV3vWB8xYVHGIdX8Wyum+bpECfxiblAeDJ
V+xatpKqcepdZgJMgrDL0d/F/iyx/nllMdWQjUTivBMKq45SRgi3xJPzg26Bnbqs
xHvqvlfRVxFccjACUj1g4H1gyqx4pP0ETihg047QZJQv4wvKdBFkhxh5W9tiy2Ou
6i5JFZhi+B++2n7QIs0IHePvgf1CcBRugaOixa2D7HW15hsvhCX5On4UxJz8cr0w
38IK20dXViQFlBZWxHlnlBO3EHrmGi4unMkDMLIUH90hw0Dl3Nyq6oA7+EBdOa90
Iao7deiYoURYX18NIEvCrSqlnh6veN8XZmh3MHxxH0A08OglRDxAnF96YiW2Rm5Z
Lgyzyr8kB4dbKa3Zy9bNNPZuiGXHVugMatmzIUYkpdtucS0o8WZEltL+sT/Z2DwZ
i6lHufwf9Bp3HGFVfu8NZyS3RyXEiSiu7D4v6/pZU9Eqn3G2+eAhsFxdk6TD/e10
3j+cK77yHPZgfEQ0VXfCwh65yUKye2INecA7sKuyd5Qz/LTYChGiwmaD+JeNiJcF
flO39Do2ifn73L0PWUiMSsDG+2YJ3KSIzn+dSVBpxxsUf1Oy/kmG5aNRNenJkwQL
QwqL3nvA1QLh7ZwteVDDOAx1kJSyyyq9Kd8wyp5wMH5YRiigpsSuVDgpPMiVGYUo
C/67jyusfKv0Tzn+lae8W94u9F3AuWekgILTUaZwS/sO8ijjgxG/gwwqaQN8/DRY
5wKBiMCnXJ2NeqEoG7EhKMh871I544lQIUxHPTXFJDCqg3ya1Btpvi0BJG061ncL
0yeaWGMEoZV0OGWS/cF2iV34BDBNGTkO6gAbTaq3osgrt8y5Rfd6h0mTIoyR3VhP
T1pXPiKWVKMs+BrnIC0hCvdCRTuH+bgYIsHYVxEkZWqZHynBvg9FwC8+W17HAmRc
45qZNi1AExfhzyi6+OtVcGP2FHagdgHSFg5EX3XQfL/INVCWumOhVJdkF3bGp4Mb
L/p2XN8s6CJo9/mRU/ZpxSQaL7kYrHzeaB3h9fr3UKc+WP/I2aly7J5o81SY3r/L
tyHn8GUdEr0knLh7uwDMb1Ujelv81RDzLFWtuQffUYMolI003Cu7q/yWu2Qw771j
BnOytscAjWBp3Eu3+sR/fZ6pBpXAwBO/wfKnU46NNpBFxqrxmV2830zQet4i/ZOw
TMe/viRWmKAC4g79fWrVACPuanuAmB1Jo4WZeiVoBkCVQyZRzHU609dvue8NDIuG
ukWY7i5jvKdoA2QFrdYYSIq6/lr2n5Ag0Jpe44rLufbJ2ryd+gOrukjUgss4f7j2
8fVR6mCJaKvSnISLbujRoySvl1TsnFhKUU2MC2qViSmBbMBTfRmqeDSF4xYmFxre
fAvQwNBIddq5/FDOMZzL+51p0NP/1Lf2RX7J6/FegdZasLUSjcHargg90paJa7lm
r2JA1Bbe2n9nbYv1PdulxyVcT3vrbEs7NwPnyyeFy7wvjYnB6FsHXRnG1u96eJmA
AvmzGnEH7HhriGBB4SK99XJzPGAfbJ84SKxd2bberQGI4Mhys1XQ+Qp8MIp9Qu0q
8G9imzMUiVhdecwuk2/fR2hWu1S/T2b5dx0Guk7UMCKJr+pjZo8n8yTjzwDZ28os
2dmsnhUizY/bz5DhptA1UkJubDy1SWXQN8oBChq+YZUiBwdxTmyVcCfMNEf5xa5f
hvkWkS8JNJH/4ftuyHlggVpYmYNyLlE6iPrDdQSpVfSyeHYPKHYGOW0OxZ8XSX1e
iZ8Tluj42d3yJmmGq9Qfi3OcNYIRI2faygh4yJBneKyjzBCbTIP9m4J4KkBAPZwV
2vUZY5uJBbXkWV4r/k0Y2joiYdvG7174E6EtLyeooE6gP1JLy5h1CRCqtMQrdhAZ
6hsBjvpaJAvZP6LxFhpCnui6ewyHdmligbHiHF64d7IhyaA39f1ayb67fMlJLVev
mxCExWR2vZ8Haml11ppNITEyWxlAFisJDGoRSt8xfS+i5IuhkdjzhLrPkNcgMn00
reBVhNirIkg1WrnKL5TbSjde4pDaGy4q3aA4EwxQu3hK+sghxt/pJovVNVEVQbOM
TYTbnUsJpQnh/SlekXmSQI+3G4qe8wTq5285WIw5Uzgk86zBSHRHPC8KDOeLcp7s
iTdSICH2m9cUnWWH32HaTI4dw5+DEb1iZz9FKwWpCv+w2dCIJ8itRN/L2vxje1I6
yyW8RTKVnjp/H2cheN+MftFdYTtYUFwoZThr6+il+uvYwG8/UQxSueaHHvQhVdXN
s9k2wfcW2E/1agXJ9vrmC9al0qxX7TZ2K6pgKVLjpoiyyG16cjk19g6xjZpFSDwJ
Ux0QoWYn1CnwCaEA14VTIggpLMDQs2+1D/TZIbZwQkAkPc8QeG61dD8r76pa1OJ9
FDuk+Z7ycWpwGqIt6oB0BDm5z2TKX0qB+kXXv6GATMB7FoIZAd4iASHZn4Pb4UPI
sFFlhFeDsugMCaPQwQQSrY/ou8gMwiQCpJkLKYzAZOUtdCsuztM67juHTYhxhhCA
9VGh8Dx5RvNs0nVb7hw0udT3/XzZIndZ6MlkKrBwgGP57eFdG73ldnJAXNNMzumz
eO9lCEmoX6o7JxFQ1DmtL3mC6F5tJ6agHg1MtUhjtt/JUsuzPif4LFWSeeoIgQWb
XHpRx1VxD1CKp/5wP+Qnr9b8O4TjMs08pfuh8ufJ2XjtxGAmw0Marynhb1KPFZnw
QADDg8ZQMdPfG5iaihlYZYLJyImQx2c+r2cGw/a5gQVmR1coaBrLjZ8+7hu7TogE
mefiJFXoxSszwnalhwA03PxCKtbGSj3RnrccMMTlVF2k9OskHyQRpxi7IGkO32x+
HeIya3c9Opg/1ZIf4nvy7EeL8+mzVRJ0w8W9Q8eQmZ4ufoNWIYmkMuq/nViugo/a
BmLmqYWxp6mYSf47RHEaZyquzXF1L0EL/o1OloMY/LUpAmaLjFrvaGAdw4HgTroM
QykE0hFNCXSmoeDcKh/X1u39f9qIXM4e6z/Nn8LBgXNKmkrPzErJ87+y+snhp8MZ
Y8LMxq1cHY8fVY2ceSw0oNFA7ATZtBHyC1wXrDuIkEDYB+bHO4bRPknvNCFfn9uI
Zby4JcZ89tQ9BykRhwfdKCnxwb4wp/J7ClLHJHanXsYlhbPAAyVcRz0rMR1UQqaP
H9W9rt4sSOdzukGdoGVcAD6c2W+Fo9B5x6B7M7M9D1K/yS1P1Bgzd8wDMCkpmMSh
oV7i5XawKmR6FVjtsgj31lJw7WFUGB6u75IDldOyMF2XIn2eI/tEM97Q3tq6GY+q
dcZY4EP7pp1y0UrSa2qbMnXjBVi1Cb2iM5I5BPW2Rz1POSP2LX8NMq00tZE2MBa2
802HoTYPoX0/eUGEDCa2EVamFYWs0HSkBA0dec+ZG4jlRD/9oTaESrydlWl6a/Gu
dXy5g4Euin4B3HERL6g5wElLfU4mv1Tyjv7FWkgMYzPpKRUE4pOBIQU5Mayyi8y8
kpQrUdir32aF8ALT3WuroA836kocDqsCbD3NsFo4iiK50R0TDLzkVqPe3JX2O3+D
d7zTHLZGf0HLO2Ll9Jg11PslUiYHfDO7QzgOPAYSEz3kyM9ZvFxG4vFJrgol0X3e
opTqSbhiC8O3swfDhrqg3Bqkzw5l6EUbfckexa9hAmgctpCNJKsSjaovesQn7/H4
c9exT0q4VC5Zx+qBJflWTv6XOWv+Y7EhnCiDiXzvP4fYOt9UuBSotyUyxlaU8tkw
RE/mUuDoQa6zcqYL1jT2YYRAGlHW4GVwhJOe2mT5XR3N0kUW6IF78u4Eh8c4mII7
oR9H5C4kFCdVPuHIh6Oa0jpbZQgKfaRKLbGspAWVkt8nTeIbaQmWKbxCSoftNYD6
oEZ7zZr3UzsRnGBdEK+8M7Rd0agDqDHTc7UubiWVpvH5Yqe2saUBj9kHRaadhYY2
AujZ1WGW0vOzHBKS7Selqn1sRDA/VnZe19KpUly4MFLmC4qG4wzlTL7CbTaA8xsB
PaleIuRrG76w1elYi+k6pfzmcLLTk0zazXMYrJ05S+G/jcMJleDlwkOOFcXNuvsQ
TTQBLvGBRcBsu6gQeIJT8+Fid6Q90ll5yMWREmkyEV7eX17bZAMiQwpZyTJPUStQ
1zQ/Gb8ofPA25dYuP7yDsduNAvjqklojQQmONpNEFW6Cj53F2OpPv+rFsDdkqjsi
KXHi7V7FTxOs5GsGdhXlNbuhVUUtrRrJshNFe3CEUV2y5Nkfdg8WCnsxeH0LV+zH
bxlDMPiumX5TkliKWT0EHoAthGwL6VLKY3bBqzgBgeUpsqHMFcoF1R5OQSYKTxnV
7+6bCI6RB6e7JKpZ/kPuISsDU0mqOtCuiJLYt1fKDD8dwpFVRisoMSbK80T0xaau
8Mc7ArGLQz92FgTImQTjOd8qNCGUrPsVPFDlKXoWOI0nv2oRsWt0+oU2NXxLLj0q
cOemBQxyY9v7sRt6SlITFNOCjVw7fe4zcSJcSP09wNNmunqEDcKFSI0MG9j+3Td4
tU6YF8kiLbZ7g+izizUntqLfgS1C9s4htHH4Zvte1v/3t6HkiKUL518Y59PO6QrN
LndX0TxVo5InU9zAxlcou0hUWkxF42wqu2N85XEJ9rw+LlwEC2GY2h5PtpYW524j
yQE8CRPuOZwNbliJ9vNZZe3VsPRHfXN22u46Gt1f3k8O4TNo85zhp5OZoHqLvNYN
W1Lzd+jjXug6N4pktdc2rzk4Go9X6qI7Rf9W1foi35GOg+UTt/rzWDYnvIoAioU6
4vCFc0kKFOZ1XaXJ3wUJsetza1RJuvIGx4iyKhk2WmdxF6Vxe4izEUcxZMaxERhL
oby9zO0/JDjRFq54ubOX9pRY7FJTeesfvAftWNV/dUq1LQRQsYY6pdnJL7aS1GYk
UCH4QainUKTSYF+qgRKscc7GY3jQFpvIP5Qkj2EBDJFazzleb+CmJt/Hr/1SW3/o
GuGCVmImTuwpAaKFhHt5sujVJSJB0JD1hf7B1MzMPLh0xZUtqMDZSU8JyZmEfkpX
p096/cm8kJonSNMxfDF7otQ4ToWFeqowJMCzxySYILRvsSX1QnWOKo+pRBnjcmOD
7RyLPHsBgw4aGvsCmfOOB9CHwYvvoqVTnnkTvqFBCUqAatdnT7jYNA3V6Nrj98BJ
e6xBYouCNblrbKzYGOAIdnzOk3kSpd+iMjrF9wZgFCfIfHYEffjTQswxrTLxNj4W
daS45JoJYHC6qyp25toftThEg/M4+b7klDt6I3cLVJLtPvcjrneegR8Th0KZGNjJ
4+Zt+Wu8aR3i11DR9fOs1+nsi6jawvfvpkd3PFt9snHEHA4Ta/Puc1NxFY2qQUbt
vAZCrBuqW+dl7J8KLzxJ24JGVM+z1n4QCcTQDmMGRrGMV+2DgNNhXjytd6E4hfl4
jv68EKkSRiviDreF5InInr51nDsopTcsM50/mzCQ7EI7IEVjrOT/QbrjJzvYLNTx
eYUzKTctAVOTjfsK6DwwAmqQvfT89xMla+IPYd0hTerjhkxKAjn08YxOPwDaBV7z
x1Sb2czADoQDkgYVgFDaxe7wekXk09ycAfltzgs1cHxdTUSpsvYgYh+llZEfPBzG
6Om/0evkF2Va1/LJCogcH+KT1bfMHeXP/cf6b2V+w1TJxCDH4jZ/Ha1uSJgAUJfo
yVqHGj+vL4RyRNBFmmRM/OFHVInGcBo3fyyLZyP9x2JuodjPA8MsctICEAYV/iU+
tl3LCQOgiHp56pS/8hCOTAYDKFrbyGvGom9bdJKzEXEAOyu+Tg0JEiO4C7AT4FPy
B8rur4+EEvcHs24Qxgmq6BZbh+Vy9Bi1IwRJ4ag00FVTE9XXhjsaaId4rLzyaIC9
XKt0Dn24MUctxgYr7ghSJQQcWQ+hu3EhcWjlXebEmxi3T9tp5a68mhxJktOYC4B0
se1FFgaIGvGZIj97g6Ypo0eyqwIlED5lB1AcQPJvSxvtWUzsJjYjPYFAxd88QEew
cP2jA3yz4K7hgNyOsA5k3PU8UyPkyqnWDpkJXBMSr3gFoKkwqVveOrJhMMp/Pw5a
mnas7OzTZDqWuPJXciin0DgoDQ4hZi83EBR4/0DHnB13s69/OhGehHAikjniwbDR
CFS74KIvBEUp5CJzvC+9Hp0s/kdc6s3cXtKffS7geMQORroO/+K5DwmvVH1pQZac
TDUrgkAqAZFbxb7qLRBmIpN2Ag5Ygij+9+dt+XnUnAo1+9/8UlESBCbfaWBTyoQu
MAbSR0xdEghuQZBDWDH5M4emvDOMx1DmRVOZ1xoqiIx6g6EBjj7KDqfCe23/SjpT
30OJvrtvl3XpDXKQpDnmq3NKBwtpr+stBrR25/xqMNm622pv9R3m5zdyWC5xwU+6
/bvXkm6Y8aHWu+SqzsLwKsY0B+W3DSS8otgtzusabt5bFXezlLIc0IvckNFYQGeN
nthTel4WfOlqLvB5Yu8QMo0JXq9/lQsgLKPPxOSwVGhJGopzgbxizqNdBqBitDQB
XSugmoEH09/wEvULlmGS/5OyJo177ubJ3Zr6j+gHbxH+aRhpwFF71+sK1Qh5DOhu
mfsl3Wj9n7IxGoegxl7mLSXXN5eY0b4RYcHsuchMbqf8SWArduHs2xBaZ9cwtuTP
WKaRAvdlz7UENPZOhWze//F0SuHQ73IxCm7g/mjma3yEfb/6ARnq7bKQaOlHLAP6
ouo2rqaP40SrEFKwNDypnhx5iBqjkF5W9zl9EYlAKfEIZ3YQZLSYnHCrBrD3rb9M
9mF1h14Zn3LYXg7YZPdkQsx+3ZD4GaWdQMz0P9OiPjzpyJAOCR4X1VgrBZ9v//cc
wMzZ2rpdspFEhFrkzP0KaHxctOCZgg9tCKOMtbYlUUDClkTfkr6DGMp1kTzq9XPM
uQGPZU/W6gFom3zEchnlWXRoBlQZdkZ6jRgdjQoER8F0msh5w51EQM26xkA15lPo
rp4gLNERP5csAwZnAQVWd7c8jkmhZhR2EnTxrOU75oYcaYJ7mxeGnVPPEEbhlS07
CoJwbhqXkHkORpsLe9m2zlGTujq9wX67j8ZzTgpED8JeGuwCihzeUlbBG9Qh1lgk
A3Ll1ATCbu7C5r9404q/tqz3crETdbX7BZLeB+TCzNI1zmK140qGFIEW/hB6bSBJ
CYHLJWPN5xBmPjTn7q+tJv/zcq5wAEdCGzr3ZdnqoCMpINeH8KLhKvgCjjhDH7a+
iHOayGyIpYvShCwbwLHRvt8yTsUPa014oSRXxQhp6pDiBXfnge/K7I4iVfU58Ldj
5Osbbx+Eu+/tJlZVdMoegTgIqmEVRqvyBQJscd1y2LxE1721SQX9ph0b8I8/ibwC
OyJ84OJNsx57ZY39ICxl8U83WETkxCm04hMS8ctmerS9Lj9YxNpWwm3IBCg1SP+K
vHyXlFaioXefkGr5N3NKHXnzwayb7E427UV/6KsGY3HUi3+err0LQs2vS/K1msJw
IYczVoC0D6QEQlsxBrp6XHfHcXK2AlT5B3ybxrvyQbtKvJ9ZjTbgozpyYqUjKgSw
GmjfdjRk1L/th4/2DbOYYDiC0sBgcC/va3Z8SQy1Bebyz0lHjyOGmXqOYC7R+Ztf
OG/sdMZ226+yww6ne7yq22cXoLDlydWirFwqaT9fBFU+9vtgStseHHp4t8kQoCCB
uqbBKzswl46kn2/09HJHF0vsbHL69cRqoYh8HkWCuhUgVS2Y7ZtQxogkEWEEAv7l
3s9i93FEhnekHUhDO0gnfSb4I8RmWkH0/QcDKCXrfazd11b15e4FxFRdrfQovuUs
WSsYyJgyuAmpgDf6VCBXP8+JXWhPpIGthv5PBCNYiQ0279DA8f+7kudtCQ9kgOwl
NiL9GEYNRbcnbfWQ/ljwYsj94VmZc0Jqf7SDTI/Vd4ngYot9gOloyo9UomCx6zm9
J4GOh0n2ofuc3KQOo93XFtUFmQVamtSLrxNpvVKoNuXOeVi+OSgjOK19fqHD+W6h
ZR9KddMeZb92pfOc3i5VzCQvAJmxvYH80TzrBNwBSYcJFlWHMA8QWGVsHAM5MFNd
FJYw4pdiPpKvnrsph5N53T/cU1zDxSrjzg55RxFjXGtgDnD3uGOxkuZkEjiXjJCT
2x7ATcU88SLhPBOia7/0ll3aMC7WcrjEa3S4e8m0w7UYZADYqqgTYAiySyfsIheA
374nyqMOQySN+DZ99be0hqR9t8DIvKWYN4I1hHj3Q+hrSMI6ti4WzogVFKpyXync
t+1cTqFENsG6UQ+7eDEdwkfe8sAT/4ZMBWzHroONLO1+XhBNh3Yxi0ob4srh40Lv
8xWRKvzAgg0qpjrvg13ExddrTZRJr8OaYUOsZfD/F3hDW5An6eZf3HsKgMZDDp8O
BqA2zYG+qY6jGJIVrTDw0hO5GD0VQlk/ZNUji4C1pe22fpgTW9oSw2p3xSAc96db
Sa8ZOAeNFNaSLuObpKgK+cwcrqflK5pPFGa1xQNV6LTiqrIu/lN6jVVpV2Mr8hhI
fYkTjL/teRMdIhE6zSo4icTdYswQsMtMON94X/YhqBD9fDloiSCc/nsCtEKRSLCz
THwe3W7Bud/XX23KxS3SoDYPVv/DrnkU2BioEaz0EHCvut4JiVpp3JLwl9LgLeqj
6gTGThLWmdU9pmyhJ/djt3le9KVx/PDewuo2cTksniJYPgOG3Afi1RkK+jhUdFCV
aRN1Lie3ePP/42GlZFeaSwgZ4Sxpw+9fFUM5yOUvCb6rkr1pAAT+tPry/oCi1q9X
d+y4u4SNG2QywlVpJI/d2R9+l6ViLPkXtibDShsG/xfPwj7hqlDaWcfIafBmoURF
7g6rMYZh/R5TbPUqdHnx2gaOb3SHdUOb4d/CmVbqe8lH372coP+iIHMxr60N6mqS
wafS1F+uO/Ll7Z6QAV44LA6guDrhJiX3uH8tuYWfnt9d0YJRaQJToLn2kAI9M/+4
ZD/AV78zfNLEeIHR/LmNXnsVToxYVzAGcJlxR5TFNRSTNdJrSFVRhuppu9PJyWsX
HKm9E+tILym2o3lqywMps81GTPvEL9eF1xCzWOqNyc3O6/JAbbmjdawLeql2lKE3
dm9gy80DpnEQz7gXBzVWUDUkMUVrQ0FJC0y9e8/SNNF0S5My+xgfJ7NQAHqdvcYn
9NdarbVi9pYIe4JO3d0KrQ34jMvAvwV7WcWJx0MeQgDRz17SgbCIqVEHa9vVsyYb
IleBeQAYecLjOHVF/jwPVWXJJgfiVt5nOskQk87/2jnNsdWLZ8R3Z2VUIz9Kie+M
xu63lrwAhejVjzSrCrwG4OSddwrdN07M+WRrjVCiUmUVrxFEtJfEHrkrYTgZtjR7
tbB4Q4cX5DqnEHd9cK866L3oXqIohmO28yKT9oABuWqHodSBP7zXUMMjAe9emN4U
6AvFP5tybBtCHXxraOErtdmVyGirNARkm6UeiIaenqucQvxwYtwZ5olEmPalp6xW
zol1PS/eM7Uc43m/HSJRfz9FAQZVs2s6epB3b+auyFigK0BpeEJRq57+OZOMSvBv
lnE98L8i7ve505F99SieW4oCzRKKHNWjvIlwTNlZyWzHzHxBQg2QChhfosW4b+f8
nXJkSr609zz4zj/nPD2XegLaUCebYLBUTrFqnSpzhN9MlqtvIqbxFsyXxPaXlw14
ivNkFyG3qAMcgG3BkQgN0tgyCyu/67dZKuZoDd7E/ZSrLhUS7st1itchPrz9teZQ
ob8BeBzhWteBYmD59CtQUeqOYlHs3Ns72fR/Swvzo45UxSUm7Jakmj0x+dI72cmg
`pragma protect end_protected

module alt_mge_xcvr_reset_ctrl_txpll (
		input  wire       clock,         //         clock.clk
		input  wire       reset,         //         reset.reset
		output wire [0:0] pll_powerdown  // pll_powerdown.pll_powerdown
	);
endmodule


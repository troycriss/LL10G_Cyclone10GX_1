`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
E9m4FPLV5TIe7lYLJkBZwjUzyI6Kr+ZMNIbk4gdTd5dnJ7/k1OEtGygnJgji1L7M
Di3vXh99vCKPrUTYue5oRZfBsRDfVh5S0VoxpqVE5wacYqb0DGOLIJ8Kf42Jn6Hs
bC53LMZ0h4LqEaPxTMPtqOWdFBerY9LxbxeeajP37ow=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 5792), data_block
x0FleDsqdJWh/g4jh2ufeDGvn2VT3OgXF+gfqWDIH+bOETWhi7PU4VN6I7tIvyDs
y7S8PQ1DFGgfsp3PbR2RMNfwq1DbA2o8hXlfIny0pNsGEGYxLGa48vLcCRDa8rcU
DmYsW3DSwwotS9+HXz0VjlEJ1tEYFr0/vvwwH/Nv5Qbhy9uvI8AEzGDtyQtpqv/7
Fow0kwNAOKugXubHKs0S9Q9eRo1eC7W2c0G/yLp2zsgd/TWMetJZcD+3YKCYWCT9
ENxndtn4Cm5HXbYRV/E69nmJ4bPoJKrVcnPNjs8tfcuGgZ//JWk1DGDmRaswbPW6
5//Ut/VuRjQ2ac6UIXHR+gRd57VocOxBITFQOaGnEcoW1MIL4ADJbJBqmkZ0Gwyr
iRMJL8j8YSDmWQyz+DhoASobOSfKNi8V+q64IxepJu6FOs/qzZPtHxSn2HbsocaR
M5f4w3R43QzsqffZfn448ntI4+e4B2lEKLVExpJ1ovOGKLkGlouiKw2ALSzRUqOc
1yxJGD+0wy4AkkNK6yxmklrgY7QzmL3u/94aLE2MWSv9Zi13Yq8UY8hxkkkrybrW
4DiAZOy8Rwc/zhgmSRcBrj1vmTNZIQnpxhgweCwx+qa8ltwiYJihC0XbSlTgQu5Y
+h3prGWHZzBxr0ONfsXCrR282BUUhZw3L+/MhccvEI/z0B5pnwEE7rwhZEg9Uz2e
Sz8SK5sdYKqgb7NcMXRTxmdfwQJti3DVumt3IahUsRCZ4DlEn4lSp2ByPDLrByW6
iewSU5v5ynOC8NoLVqFk8yOIRcmkPTy8k9CBOhxflHi2lscD16dNeX1HBLBtCfk4
NlPHMtUEshDBGLhmKG+ALBUoBjadgfVCcdG+tSik1SHa8Ps6YPVreLAqS1xuQ3MJ
yBDWoDuvqXmiCFkCFWd8+6KEib+tQyBoLYihsGlBOQ3eRQ2MXu0/wlgFFdOQOtKs
o3c1Lm0DvqFOZp0WvNxErcj0aLZ2cTrw0kVAUX3uaIzo7231zRkLKk6YCS2FcpgK
/Bk+cnMPeAeMJ1UIkxZFLtL3THwhQm9lyTOiffSpeIvuzFykE74quZ1cEkmQnj0N
qzQFzK3JsLzYYidKanup4WbKkQyvibMXp/5aqWc2s3RkhckCvxxYWo0ULa5ubzfm
4JRnBzYlr2C1froW0y/rLDCcaZhHSta4oDV0WeLeJ8Nu/v56QraTtLzzT7aw+r0M
60Gfwe2DJu/GOXv4hNE5FFIdrluTy7n8qLqvW1cp3UPIg6XVLLXH5PZ0ctHtf/6Q
Q4FhdlTbP0v0r/0VmUpy5u7BMTGExw9QbmnikFixJrLJUHgOU1l7AtX15RfQs5n+
DnlEgJ3zgEa6UZbSNNWCTP66ykUnuDtGvkwDh1VXhOaeDEXZwNSWKvx2VpIJ8G+D
hnUpEGmcKbpnis30vyBeEIPIUIjsJ1utSkZBnjN3dcfv8ZgosYht1Qu3KwfwvMDa
3wm+Ba3bqhy5Rg3jLcHSj0ZKce4Nhm1h/kDRc73mBNWagB8CaAS8vtJQdCJ1PFAK
iOGgA34dLh75SqokAkjgDZC5kzqGZZfQty+1r98bJbcnjLt2yyNzOSryRUXnX2VY
CyRu78Y3dyq99u0je+9nvQx7366Zf1ELVMMz8ozkOyf8MFc4npu2sv8EVoK0nIth
hxr1/LiRzj7kN0kSyfvakpKcDjM4kmD/Vrwy1izUWAnwNGf8NdFc1FsjrB29sPka
IeIHIeVdo//CN9gEW5q/safNxtlObkGHfe277E1z3AYYFiJUCWwal+DosBbR+Clc
2V1/464GSoZhvNcKZCjp0cTrBTf2FiHgVIhLhUezYsM45YZr43MQi20F+8kBwu5U
hhekH46iVNpB/HiTqAD3b/GJUquXffa528IfU1dwAGr66jwKXDqlJdgYojhasD2v
FZBFhua+BhZLlCTWBUKcSvFIkE1vQUchnrTnXD1Tq7vJjwuY8yw4NUR+dgyvN/yA
qiwNMGoxM1oZxPMXyCOtYa+NqYJDZGXn5A2nL0dfcMbYDl4AExgJaMCw1HWWo65U
0fsjSncWnJe651Vi9aDWhFLH++K8044KbMGv0xHWIAuX6xvl58fVdb4w9kCvkmM8
wG0svYpdyGvgNmjxvhwfzfEz9o4C7++GoDj0F01nwym03fw0dzTlUmXRijFGsmdk
jaHKlpWpJUieEBmVMIhJqnbGqhedLBolI0rVFW84T44guDs+QMZoMpJ1IJK0jpPG
NbzrII8bZHz62DbYxDCJTqIYwie6dsb9qy7XkvaWOZVeQqgqlxxMVX1QVsuVBm6I
eyMwFgJF5J/wKNN7vwBMXU8CV0PejvWHLpRql0pDbf/cYH3UnmYvmTut97XRx0HD
guWi4gh9NKGxrMVqKL3OFEW+eKs8bwMNMgCSgCxkvdMbndA+77OPvAWLc5MnboaM
W4nbMUif7Ajcr6IsYuVrqyl3jKu1Ib4g2yQG3mEU6BWkUwPMgCDoqmXv7dK8iGOs
JVt65tqTL1n2oGeZxNVmyBGDhTghn7vAvWNvJm5TDNqHzxMdh4gXqPVvhCXpjuP/
IHUB/Nf4UsduXNFHqvPw9Y3ayFUYJCQzbbf3pcqhQLJcCX08aCqaOXghRObPJuCT
E6hDzy+zxpeAHIG0LsGzvE5+KTQnP+joWwQHc+ixTdDKnT1vf07/0yZdR9iV8ijW
DdVcfwutgHurcPsVWA2K7OBWxwEXA5kvt83dQQUPUmzFLaGuqPa17GK75f4e+uMg
93vLRIpKa438dSPjM6FDbIwenmUwbFhzyD8MK1Z1JvLLEmP6bLeuoUe2no9BFBD8
oe3JdQJnMYYbiDS5/k4WN83es0+6IyFGmMRK+btBdcM5MBu+K0A7oA01/YTAh3FI
t8D4BNaHh2eieyyOdxryHkhUN3jOelxFqMex+5NYshNyY01PqfsbRUra/JG0tIlL
y507+OB45Jen4mvuYqusRcmM8yV980RUIUvC6PHVOZIYB6UhFET2lx2zc5dSMqao
t0iW8fDlToyCKv+P2Fw9dksbRDuVsLsxVKAcA9Zvy/irDBwcRSA+w3nZjgsr1PTb
rp1IJtiXiaEVGkzYZZC9QSR/NcAtshrXJ04zOffYdN40ObyL6srRGWFKXu8/b/qC
QlQiiOTcV7Shrf6ZqnsHKQfn6iY7q9obFQN8V0WFinNrRY6KzOLl6jILS0vKssev
0uuN7fGWHO/L/hd60Dly+ZWIjVOVW82QEYkRgRURchG4aH6A31/8taXNLNFs28+N
ye//dHgznyeAvI/RuEIIDefVgkPx3EtHNHNxbsJGKHBdoZW+kUXXaC0D1mgvK207
Rhd7VGtOezFxKtfYEpr2Zt/60+5Js2UqtcdZvSZa3z134HvRsFr1Tq5ZWRESTOUA
Z/5HLhLu+NbzatTb3uMUW6LkBjIv7ykREmgA4MkLAvrPvISAIetUVSD8GtlbVEmT
Xd00KJhByZQEBs7RVP5sX4JwO8nq7bernShTdO+R5OQ6PaB8k4VHXFllN1QKsG++
gUPRLlnmqVr447f6JOdGcKeqKldHd/XS52BayRR/lRlY1DlWSqURq9sbD7o2MaFz
82ctbUnHtQHgYlWj0ruqmm3cJwSb1tPG+m4P6zWQA6KktKk9YCw2b94NATZRE5NQ
3uHoQmRR0nw0g82lcI310vDAeKnqHfRD+ouYbq3Gdte9J1TR8Q4n8tPG5VF42RiA
FZ7Pt1sCZ4XELjxmx959MPL0b1pIvZ+FGnufLdxoHgr8h7gm37MxN/OAzc3b8Iv+
F1T+KkS36vEu8/OeHNRX+vmfbQdFw5E+5eMvCj8i7rbCyY/jn2nMO7tvKzOegmMR
2vudroIgsBcQ6DjZhA+jT/B7yY3RZ7PtrT3VdLp+oXxPqo86GmfXWFib1dBb+nCD
cHYjvh2MdImXMf5F1NQehvHpsSmnnnLTth8mfBX8fbezqutxTxbgiAwLkPRg8TPS
qAH9RVHAIeMhFnJKB42WzPMJozHXyD5lHg7exZPQ+Pfb831de9lzWWYPrEzJ6VTC
xb41p6j31vH1mTnmKDhVKs8eTbz5bNCcB5lfCa+MP1hnDPnAHPCAiTGOSbEmbKzi
7GA6jlaGSmRmU2NtvJCN/mRLoqnxqAcV5ExX8/+55I3Fh3UUwMUWL1WO86hfSFhU
q9bZPPgwG1ulP/6eYNkOyIoUeXYiJT4tCQSVGraEPj5jc5//K8SABGscVZiOit5Y
9WRofHYhaPxNSbbWFD1IhDBfs/97BzWGlzDNDAA/g2CJGGZnahWf8HhC0y7oRiaF
EchjJGIjus/QfJ3MlqhqrXxkxbLMgwCPqGipltWPfTLNYNeQA7Ugc4Hu8gxJ7DvB
dufjcFPrS0wZnrRfCDCQtv15jODcpvzae1eI9rnJadyDnZOo00v3cyCiB7i+E/9Z
Lx7ZTNtv97cXlLGGr/VI94j2LgJdsUjm31a6SG3zsm+kZYAwaO3/THOl162Ywzbq
kte05UFyp7CbP3cG5EzqaQtjmkeqpyrluSpjf6yps/hphY1rAOw5ZU//xliL5xdk
MqnO9UKhc5OyO7vZb7H5c8ngAMlHYFZIYsodT8DzDXsvQ6b5OP8s9L54Hd5f2PnG
XS6WfYSEnGLIrnKl/A7vN8AfuirxlyJ6T7E9Td7uZ0X9GuTfYDJpvFf12/pWtLwb
p0sP+kuwxvwQlyKi5D3+oU+8QmnBZLeM0u7/79A8R0lWt+EOWEohY84qMlQZeixF
/WuI31LM3mOYjxPA2o+6RlKCoofggNxxW0C0sHjkJ1UH32RJAjba+sc+1UdFbKzg
qB43PWR2hm7TjVtMCInxV/jebjggyOjjn8p5fSc+u9BYaZ002ERIIQef/z8AVoKF
py6QyDkS5FzRKNeclYTB8cMUteWKEwvBsFuBJlixWZkDpfu4rcXIaKkyNHFn2e86
3RjcysTUxMUINgZGT70vCPQGNp/1H+AiQ9H5gb4BZMk80WHgzez7kx0nBJxedxH4
C5IpzCL/j/1WHjO4fVfn+67Vi+1bjow4ERPVczotxHMhpjqudYPITg3cZCmP0Q9h
kj/KtduzgUOyIUh7+hNXL81zn86QaXE22bLHMO0o4v88kG7iDzlC3M5nxmgh8OeV
Lz7k7LmLKni58RRPUhpSDN8gvAdVcQRunUf0+6mbBc5L6FrfiTQV2+aq+7iyQwEX
vs3nz3ZYj1EJv5TPhLSs1jrtJi9gMa2YrAwkUV7s/O7ggCydBcMGMTcH5p8FyuNf
qTmQ67/vCITvKRV1UGFYHhgk4MxyPokeuPq40JFH5lEocP55j9LujUzmaLnQ+yrW
ek82HFNsmkE9/mkBnEVbdsQ2dJC05LoEms6wLQdlO880K5YP9fLRjJ1WX/QBy/OA
Kxlbk6FBP7HCytcWfiw8MgjK7xY9HqKlT7ovkmpW/iZSs8Uo1iuf7UG74zQvtnLq
RTeC7G15PsLDZVsFs6yY7XTpSJEas/6AmYo+8nkCwoZsY6qbNAKnnYs9+mQ2i5A2
LBClGQvrwNk8m6XNirW/axiuxPIboXcCmO5qPYBR7A8FXZ+b8SbvQmnGSHSPcOV6
1dmC6bAGgbvcZ8zHmdJHVP99e6ZnkItBWFKGNZkKT1mT0bdHSGiLITbi9piYSr0E
f+bhybK1KUZMUQSQS7yEP88DVWGgUAylZgySFpgX1HaSHc3FJJFNC1uqG/HKLktK
FFA/h6Rvz5KfM2Mnmzu7kaoluEooqrS1uIpmqzs3USQBeBqBlQpuyWvCJmCSHTWG
VUCxwFELyBBwLtCPKRTQtRNIj/bbbkNCxDsJ9+TTVguVOk7L4q8l9KaeBYBusqfn
I3h9atlLw3M0yPKXgGHpwRuzzY3VlVlLVIoxYNo/x4TpWDI08+d1jrOFsAK7/mPC
TXMeYp8GL7V0ZzrMvd5LLdKkPQevLqn6KJpAwu2XupWHzaGWbKhBQH8gTBltqMik
gZ97sHxqR3tlBXPNK6hwTVY5+iQJwyumz2+OD1pCuMwZO62pZF6glPI/h+2e6s6S
u0gfjmQ0Qx2Da1c5SteLlzmUVRytHN5bwn4MDpCjFCoZLzuV4ZMY4JZgOEcXOkxz
i9qCy+snTlteMHIY5rKNJYaJIQjH2YOC7JuVmJXs6YjkPBSdp7UaBmhxiyM/xc+t
FFDW4I1yhZ+NxQZFPqSlCec5xVgLgf47wnhuIFbdLjV+D6hsCGROS3XY1uwO5KQT
Wd0ZZJdK4JUAKqwJZ+nEA8L3xLWtSAAsAJc6ofgXO7jqTvu/9DUkv07vMCRSebWP
pWOSqE0Wg//qLY5tzXF0QkFD5BHIkuJD4Qrv1coIw6VvsMzgjdUEdik07o/U9g9N
7UM8PHTvtKhhwxfMOtongbdTA2DPnbQtfOzawRJBOhn9GUk+5V3cjJ1ALjrBHIwM
lGjd6VraccstiUImNqx5AZZdcinUd1t4fxcQLgSB6fDptfLERoru0RuUWCDxVf7l
6qfCsfeY4pP3nNadxYdiyvgfS47T6DtRmZw1+wDk+IwF2zDwgURiRG7jZ3uvn7RD
pf3za+4HdkBHq+IO0hrTg+b5LrGYH+zeQUIGLpQLHukEOR62cQsOYGDWkc+MBjeW
Fm66l8yrLFCIkl2oAQJgQMJe64KSlvdBCIwoYRpxivHK60eWVJfe6SJ8zWEBY5mO
SM6W2jae3/9fgRD1JEn/2EvZ5CsFdrRGcOZd4zs7fUFiozaRLGFaqaHv2Mrtka3k
WQRfuFWXD90GITbSZzLcAGrpfHC37N738Di7dk/N9/GuDBNpfbYyEC0VnETuuWt2
mz1rNc/envuAz8xdqNPb8WEoHcRsjm2qbGwaCXwL/pHFE141jUT3FfTiFLRiTaDY
eRZvZYNQ+dq0cMV4RdIHkHHJsUcjpZTum34Phy8w9wwV/+c+ia4tm5BSYTfb/ymc
x0ZFqkhS5cKlEvTX9psvedN4Ip9YBIjcVtTH3Bxdqv1ED3Yogr9/sIsW2HeMLLh5
UhJ0Q4mSR2uca5IdGg++lxT9WIoJvzNwTgSwFaD/+bpCH42WDk9LhZs7/j2iSA0r
3L0Mdh+sy0G0Dx0Cw1v4OoOlOmjZgvnLI0At5OugrzLX6eHsNH09ZviBHprd+HjP
CvOXp3v5xv7HYcyqsCMlrA5xVfFbHz9NzgA1FOt4UsC/V0Z0/9Zb3MU/lnFLnVJX
J0DKZ4UvlsDUkH5xydriJO+ft1PdRX6EuTMIndgl0E7S2Rzzpx/89LNofR4qAnTQ
EfvSFYMnBbWtlVVM6ZqCGOeLzOZOCqSE8ce1eifnE4aR24+Hq8EB9x0wncAe3LTG
hCyT4ssp26f3WzdDvW+grbgaqUh/vbnHfZuB2HmlKCD3/Q0/8buEktnIYZ1Sxmha
BJZobelIDfTiuQUFZ/tYXaO+kchyi57M3r7AcxVFkLiE3sQmUlyE0vX+gmP3Ghnv
64seXNsN9EXrlFVine5WHw+vTe2XTCZSfwmT8Zxi8Ip2iWIOd8vYgAqpldJgFqva
Sf4GVn3ff4qNMnltiX3eFJ/bD4NtLzE+eAR87k5RtgR/x5gId3hN2Wo57qbDpllA
HSRVGrhKf1316l3HchVvqAB0AY3cokAXRM+w+39vDQvX48XgNV4fKJj5cCyvfIjx
hCG46mFn+LSwQO++lhgNqMclDCgAf6/vgul8KsoJXKQrbwQnOJTiaWB32ufMOsMs
wFwmDIlyckUHa+DJhvymR3dEaj/NgSFgoj+o7Mv0vJM=
`pragma protect end_protected

// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
B5JefwrUT4oonhyx+/RyTgUQaoaNHtBkJkiW8DAX2QiG4VSSCjg8XggIM23RIahDEF4qvcxCVVQ1
Pq5QUx7elRS+gZYy/otMrwBQlwCer1rTe2x/QzP7q6Kf9p1x4lrS8lHB/my/JBBdwbj+f7i1D0Uu
kkuEdWvkSRR3nj8pLEFsgRdxe2aAb3rIXW1UTeIn0Uzg9dmjnDPt9QrspZ9j1gVknL+JCeA61LSO
JOVT0PzAszSkVWYHZbW38Em7I9i1VkST00zj7iZi3X07jQGc/n6dW7aP9uIEjhkSaiuuMjLXirnp
qQ5MGea0G00AU8NyVwSFs5LS4u1la8YBvrGZiA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5920)
e3iAiXcEU6nNMEYjyKX9waxMNbzQizUBonoAwWtO/N0tRsIRwG8nBbcnm397GuX0tQF9cp+3cE6T
Ag6s9PWaaPBqaSlNfd43no17c8dIUde2rwO2DUmhJs3gkkEM1AXt9S9AkUc9HUhCJRnvzVChbUcr
dF3emLHLEs74S0M2gfJyDlDVqKCL3EPk1QZjM2dxlRiKtAeeGFeWc0tzL153kT8LerDGsUSt1B4M
k6MC5t6BTB4RO5RUUTTtfTrARN4jXveyFsC8Y8Sif4rSg4t00qd09m4l7ikrU6ZW0AB9sYgfOJ2G
/xHveTJeBmVs79M1j/i/u7qePC6khFoNVY3jCRTWGBgsHx5Um+wamT+N1AjqU31nkYoYDOKmDPhx
SRf3f7hNDrUrF/Vzmtqi9/BbM3UMrMsfLFUWEOHETan2/iZ6lFxxh7gfpqLZuKnFafSwRUTM8RRA
3p3dHVWnXZ9iN0HnyK+AQrHhNovLwCz8X3sygJq8f68VkngE82zX00EyxYGHLodRhpt7mRrKhyFF
QowpMOpiHgy8ZF3XdrkHAl2eoDEnlwSq+urMlBMmg6+qjEhABf4Fi56IRoUBFf+Mkgj7mwbue4lj
daG336kmzQyCk4sV0iDjEUZSwidPpSVKxEISVZXD5lh5vn3LGelWlZnFb4bV4IMi8qahXYLm899R
1d2ap2xsgnxHz3THOlLVzlyWpJPg8yz17yrYBsYkuRPsY7hrcKUoasYe3SgNDL2sUzyYAbwbEvHp
/vyYY2Bka4mWN1YyIbLe9EDUWasO64PQa+IRdAidxWhWx0zneuvoLiFicZvRPMrjF9vwHfcEKTui
O81OTQjj0czZ61XmmjFNAEYEqSqQRu9jK5c5ZsuF4e6GgtjCPn7N7uzWxfIorj1D0AFyOTd+1WbR
kb3skmdQoWyOYxtokUE4+X8KFYyarDn98AFAKcVv1SoQhxC2Gll2eMR9rf7HYFigmwVvIXAnBO2K
0waI4rC9g/f72vzrDOb+lMVqlgjg91urLYdktzBrGvayRts94m9CAjL56iizTgaX5Jmq8MVw9Os4
FDBkjjp5AZSfm0RJ8Sfwd2P/bhrqDfVg/vtmM8UfjNaHlsTu0mYNg67VkgIaJ7J3JxL0kjHWU6Oy
xjv7SOT5jFf7BuFxHHmdWkiswtO7ZNsTIcZxnsFOuy+3UBBbusEABXWNJWZwqBo9BxmZYmjGuu7O
MC6+pJyBEYsl3zcxoKHzryb0ft+PaVAIrIKnV5L54W2qlhZVjtneap9hkNzy4S+5IKwaOtKbh1zB
Fa3ZfqZHQsR2fnO3jNU+VpgtmgxL6QtangabXXiZhYoON3+iYBY7kWUSi6q9ugDs40CVtPyv6ESy
TALsEWhyzXAw2BaTPQA+RM0/3XOd7Pac7HiHD5OpSTGqX0p1FUuWEf7gb0EAm6Vto21LLc6IWoSn
6LqEEFxerPigZZAGvN6Uzc6bBNVFmCqaZa+TabsbNgUgsDOV53O1qp8FvoKLBR7UrJo6+jYS5Jg4
1wegCcWdhmmbrYptoANQZzKQu1GZ4x2R3ggdOIxLENmYqkc2Vl5y2i8O3B/81TIijDHlpYfuNL8T
cf8DMMLk/CYbznT4GBC2qhLXiHxpmh2zKOG1+uexANtyS+IS113eTsaH69uSG15Fen7eVpLZQVxy
6uDzzQ6/E3at4JVPXH35MpVmoN+W0Bb+GHcc4zkOPRQe3x8Q6EievuEv0RutakQgYpRxYAP0HGfk
loAwPGkg9Xr7UcB8GkFm2K0Zy4fQT2ubunMdFb/RT21k53XvzmAskNARqhzU05v24RaOinGSHfYF
jFzkhtyLSAp/LUBqDUe3GQuj+RCyBjhCCMvHn4Jz16D08fmOALRAIEm0W9bTj4H8FMX2IEn2eOmK
6eb3MRIoCkcjLxoGbd7tTnHvc9losCb45BcZxlUS3rq+z4Pcjtn6bQv0rseK/BsFqFt9EGHbFo0p
FelARV6Ru3k6Jvvf0N/ctGDsUpiXfjhgbQI7Luy+TdKEUYJxx4Rv1wdMj3VNH0YeO87yM/KXWNw0
k7H558F9FthDW8cCdqSmJ6YYm1e2azDAxZIfnVW0+7/o2qAfLL3fIkYj81ZxVpJIWljU2pxEjy+i
jkvDDc5NrX8X5iG3odNo0/v6FAeMIGd1RjF+e0clOLgJE1Q1XDipDTTeTxixLVqEAXq0ZJdVXRqi
WPz6a8g3c6ij5gopO2wN226avOXwmYxWjcz/0BneTC0m+oaGNnIQS0sp4CCE4pWSzE0sc3zt6mXV
so2xDNHNj7cA/P4vB+BwIGl3fbVso5H/dUNUouJ2qxy+IHK1OQ/AVqM45iCip5CZ78Pa0JqJINZU
QcLVTyjq+XZyyvgZUU07aoRxqY8ZEeuCVkYvJnMZtc4JojlvdzTjRuYOlMpay1uhYnHiCh+BcOVJ
CmF9p68FYIYrCI3JM43nHNvu+by+6MzRgV1vd3ulnrO1oxTK4CqhfCrliWHaPbEClpajsax+Gcf+
9zC6H1/a2o4rjIKHFu2wsj2dprjkPaj/wica3Sl46eQDgZoF4e8kRezkalsNWu1ot2DsdmLt+moQ
+5WFqXA9AHQtuwZ8D+aSIQDf93nNiVtyBvuvD50R7LDpbfn1Jdk4Fufriq/0u0cjuVAjdNx6uZgz
/N//YJ5MU31oZnCEsBtQ/qg6K4LmEMLBUwdXeJ7ls7YWXoyLaotDXcjMisss5k7jFR9Cv41FBQIS
ZacXLijocPJEnXxReViOeTZ0J4AN9nuuV9p70Uq94kqlHYSxA7KMnnERmnQWCYOgtvBGhQbva+Mo
4sOy+d+1crlWM4iYWzhkHqPx+7Mp9tJZrL87bzX7CNF27Z1Jo3GRvUu999Le/1QIPZtgwJM167lG
c9cX4LoAR/WMDbmw3rZNnXcrT8C7ip0IJWlOGL2EhSNoxiIF5rs8F8w3XEAIs8NwicdsyGfRw6qM
nuOpL6IqTpnk7eKdbsHCbNqJ5dDhbogAZncWEUDdAiimKS7JBNTJmozM2jqsdQ5aq+8Cy7v5O3JL
gkmqB53QbMn3H8uk7gjIIp+WfAfgHBW7s+C4zyonLKbHuZqb7tTiAjQgfC+7+lk4UO7HTuA+3ns0
J6ICv01Qqujcgo82Vy1rSdJyY42yRSyR0wg8cmNn0cuTkr6U5VQ5ulWoifN69sQtEmec+0JnZpUT
zw52n7d9LuPIomyfEqGllA45lyH427s2/hfXSQt46STeayP+us48msxFbZZRK65gQTrqJhe0Nxb4
E3eLGV3DHnpfCj2HowkyWfBt133itG2PGrboc7Kh8uisgGACYgQ8BGlvcqBcaV/cm0aBX6X17Cfd
lW6DeJ+KSnXog2WZIH5M9tA3RSsKyZ3uU1UjErg9u8fJIL9Pw7AiBEeP6jkggDIxjAwR4pms7ZyY
POjlFgSPtZ3x1HdSlYsVYy0jvJz7I7YhOKd5LKEaJEjJzjVDdxogNQc/hRHJm+UO6xfMSfK/pZyQ
PF0/mWvbgLd1BPmyU1qYXb/46fwscJXg/5lDe+WwpnUc8gJ7xOr+Z/AhBaVlxLywy89Uh/t/NcDx
WM+WYHqEV/J1iYXqt/I5BIG1fC5BDe3Git0MN+a7mDaZLakGgUeplrhx4TGfLfP353e6NrKicnpl
doWEmgK7gMjBVixyju5TlAjCU2dJLprhFnX8YpSs1JBF9EAD22r/QuJxYQNfJ25fFKkFoYR8hDuz
3PiD6c/qI77/S+Gy1ioylyhyhprwiFyMiNE4I48KS1xhO11RzRYx/XHJlK7vYo8bGzma5kCb47Jf
0qO0niPers2EPFPZ4VjEOhS4Ki0z5WdFofiHqQc08N2ci6iVykDren+h04opzdocxj1SIFkF8V91
KVxY81HqG+6mBvgqS6OdwISKViqBVgC9I6Z/ka1g+Sd0Nkivhk19j5GhXYff9BwLLr/VAOpP3uj7
r+La1mZ4mPEvv5P4oblxUE7JfFcfwMzJO9VbdF6lXgyboqciUaLiz/d5FiLpgKgsQGUERGIyL5wp
5shHyxgsjvSrV7IlK/7QaRiLLZX8WCZKcGfk3DFeiYwvac7WGX6/BI+h/9WsKX9xzpe5cDtuq/kO
SvweUTA9HGt/V9Fojynlu5JXis/IB+7pzAZg+ekSwgeQY9eBHV3Z5+LCq1Gd7k25d4xJGn5OoTJy
c2oee4o8xCcI1tXBpEgeVS7Ai2yf4AfSTgP4/8nzBneXCPQoc24yemvTv7OXGGSih78i7HPtO6Hj
2LUpBWFNnZPunkGsAHVsx4npvoLzILHt1WgafnrHBg5G4jSBOwQuZapy3MABao9dJduZR4w2L03G
656Gd5vtMhIddYBv5fq+CMl66obcls1sil2sqhFtKiR2kFZYr8oYhwuLK91F8NxyJgnT2UFrwJHb
z/r+KTXEzTcJ9pYeH0w/7lPo1vLxxrnUjNLzs7tEidl2z3aNSl2YfyMWt2fjz5tJq124RSNt86r4
AbqJroeVEH4Q5IBU5Ut1FuRc8CAUq9pJf1Zvl5KFK+Co5B+agJ1rlOwukALfH26CdsErsGnAw0jc
4MniTEbeyYVJAMJ7/caHADQPza5YABP8x1akzbVRzK4vX7OuWY8dpJyVu2ZvJ5sHIyRU4LXdgZrk
T0okmTlBtqXF/Vck1cpDvd31RmxjgLZXRAytMMtUrtrcslDYCdVt0WCyP4l+ygO917wcdmZw+C/B
m3TexPXqJVwr+a8N7YqzVERDMBj1K9bT5rJX/B0I3ak2dViDegUNmyIu+t61eIQdS64+ClxZcuqz
3lpq4OOcvAwHg6eOArwPN4waqscjTon847QIG8erdIrGl5kHnZc8TpE8BOL/fuh1gWCmhI9lTNsw
W36P8WQwQSQ7GL/MVkD7YIs25EkbCpCm7KkIyYjWoavGsHXxiqDCpg+Q+L/hJnoLQ399n9mku5K5
KaXyUp2Eger147VCfov/cO0K60SkupfpUyNH62n1YjC2gbsEqebKACbyAhiI7hbfsmXgJi0NE4lO
RbrNSFGlF6ffvFqj8d0FsFDx9ukJC2mMLpnmbEQQh8Rwu6Ozg/JP3lO4L3E6+zlmjc9fMnCRvgew
YtNDIGRVybZVKRP5dYRsM78rtKBQzyzgKLC8oWCgMkIn+JZYLaVTbY444ycv1RO8fjtf/6zDqICV
vesWz38aLr39m515l6fWzyil2JnaKrf9xFyeGW8u3zLEWThs2NgguGv/jD6vAeLQ9/W9pGIOUCvX
zAkMPLRTLET6MEjhSb7mxG4kYtfzCwabuBG7dGkPMdK9eZ4bOSHChTVeXZFCPKhbvyTYooAIK5jC
+u8Aoy7STX5N4EP1JqQBLkYyEse0SI8iEuwmHfqDo8T7hvib07Xk5g7EhTvsd6KynYxmxIS2tFlR
yw237EEYNanwxKnlbw8ymy4CK0YP+1ej5x94rGioPfL/B1EI8EpeAK6dzI+g6pSaJnaTEzbWlFM3
ah9sLLV2bMv8zWIJFns0TfPotB2+I53q3lTZzumnp1/1KGHI8HEa7C6dZ5Cdliz6VTCdvjSdTggD
0Sv2k2T0QocqTKbnJc5yf0gRKMpyuf2cPGUDjnlWfKsFpvMaRaHn7LOKP/6dfVuiJ+v4ulymb7gh
rcWI0KpLuPhdYa4O1UqebWKfj5SmsSifQVUa35PCyB5ZDoRW8878sqSVDJt7z/dHTsx+GLmnWy7k
1jKpz4anJvj4PISAmAWBOlLd0fMPmKUe1k23p8xWvlFBvEl1C9gkzMdzYKgKsYz11msjP1hxeldk
9E2UTDe0zvq7xPYO7Jh8cGbr7VZSBufOAumTULJC1VZNmKN15UlYpynCOtDgBcHsK/WbjKxwQ+wh
Tx51HHTuG0MznjgpKGRUlEHdHy7CpAd+FKup+r2hZ0ExreXCxqy5UtaeLzZKD/7IYN3ljhdeB/qZ
dW5B3SeKpRaR0ZonQ3GxwqHGrKjWHCxhLIvb5PCIWRGvBr7XM0XG1aoXMY2wsk+zqCwbp12p2ZIv
c0dBCqzGxjHxUSkOq4S8NIdNvnIBh6RU6XKE1pClZd8sRcoiLdXqSvCpG8Fx/b0sPVbFJyqKf7ev
+VC5vLMwpqxPdvjKHLzH28flYdYo2+F6f/cPL3bDdoaHGB0k6P0pYAa2kNMs7djEIfoasGjvHcX9
+T3NFE0mRV52S4FIj5GrLxOgpOGz2wBpSmr/zTal5Hv5CDp0D9IyJ6GzaeMdj4C8525Jftb3QkGc
3YQsew80QqHAppHWe+p+BnxSp8lTR1eb3roxn/EVm7ogUMz1ZeZDU7kcXy/boI+fLTvxOCLNj8F3
cOXHwUyV2Ln+/RDnhi3EB4VDNlHQyPGqYhnheq4VNyvvWApVl43kLir4cV0trHlcY6/ChPptlKj6
y6G6WcK12sNHPQRk+52nkDTAjFafqhEGUhjqXkoqXJQhcwzGwCNNoPtoavMuiJwCE6M8r2H9NCCB
8RMDK8hjZ34sdZF2PTdAdZFST1OVu5XLGwPwwNpGpNvsruXzFj6moH22HpKYvynf5rBML3H7HeyL
Q0Suvv0X1qzh6Nn2X2OdLSea0glqyy+ZRepJAetegNdyeHo+4sxhO+wRPgLJAXLd60iuzNYiTgdR
v72KkGLZIPiAeUrFXpsEFq0jp6ekWWHkSRncH1NLylaGDacxQxvcST1djS66u43qDeVfzbuH9S5V
72jihLlg8fCJQoMTeStBxzKSCAs+OAq/Qt3ZNfVW4V4odbgNG7CpMrHNrS5WJAPNl/jubFTx5SkM
arWGozRY4hYs4n1u/HCLBuanirMO6Elm7XMjIn7i4yD4/xbI2GQ/c+RH512ioZCrO1rPwcmIrXTU
vnNhhz9iCVBljo80l394gWDXMokj6oW0ZhaeEDu0cmztbz4nJokXjT6UiDXGMsFxRpH5m5DKPVMe
Eq6dzdU+pgCIfUJH8Ien6qUabO0ggWua4Z2cXGubKoTY2LQjtHeJ1zNAsZhCTtYJQ/1GPqOjVp5M
ARULAjn0vDuKe3cwSMqGxPvoeOeP8fVl0k9XZ8s55MOqTjaAtc4aWx9Jl/vC/z4F9n+qCx6Z9ofM
lygVZxo4ng6H1RcX8ow9r3SIXDasiI6u1paWwpwi24P8owWAln5av0zQ5gqvaL/jCeL3P2JX7+vH
4mR8152PFY6CnytE/bww1SIiwfw1ChSeyFslSlo+hGzWpAnIlqJc90COcosqPaHmLdkTo1XEvRtH
dEsNw8mHlxg4BnML58eTF99bvAIjakyo2Ipgzwq0wliHEaLmA1oN6M0x1xJc93TAfJKM/9Wij7MY
LuK5Z4lAwWiB5PLcUA35U0Yq9PgarJWI/GvvL7e+QW+MouJctNb4q0MQLWbinn7ce192olgjiecw
fxQz8XlJJq9wh+JnIQ+/1NhXDEUNWwOZjwqAJuozBk3M/o6U+qNDJ11JGjRbrTJEmorwgzwgfwuf
o+dXdq2O1nSoUhfxEGQRB0Fut/8SpbKnyxIiXDB8LEZBqwOkg8F35k/3S2Oj1VlLFD7g0U3Q4Eij
SVUcpiSkd1B1hnaIj+hWAXJ4Uv9k+e0peLLjeHvs/HgQTptb+uzrhr3JXOISBm77QJGLA+QFys2L
qPaxMYacHn79jJzfGn7F4EtLINC14TU567LZnb0w35cvQ28dHZtQ51mCQtLMCrniS5O1UBszUPKE
AREwDV0IVApLKE+yDALaSMTVkgdib38t9f4zk2V9rpOeu0hHJoJ7NllslOFsDR76JGH1rRSFJZfY
UNqemOJuG2Gq0aqED66woYPG26/MGamidv8ODkgkK+N/u6vKj1Ew8yNRvpkmaCYNnWrAy+nmH/L4
RFjyRhd6BI+yTJ1LlQRU1kKturm2hpTHpD5fRx/rUjYoHJIyH2+4NgvF+lpkcpprhg==
`pragma protect end_protected

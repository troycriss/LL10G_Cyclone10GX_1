`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
q81cTNkK+StC2oh76wuUZQcw4fmG63d+xCoktkWRv5WQNdfBRB2gYE26718y/CZ+
/y63f1VxVVDDbqstlzWDwq/FDWLU4Z7fBfIx7CFmC6Y2Di1sCpt83MjIVGPl/2YT
O78y4UzA5KhDvG8xv4qJjsDkCkm6evAYpBdt1i1HZ18=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 4176), data_block
6U9ZaKGhyAGXXJ9opTSO3w0iCjV3KSvz7+RlTfumXpv6rsoj1NnVdPrgHmj3OWs9
MWw5TjmsK6d+vp8RfWF6WVgvgODypRsHV+X03C53dnQhddaFoXOiwlMu4bc736tJ
GTDmfAaS1hEbnQ9bZbm5k0i9cVhxL45RbfGgwKrymV5WC3IyOOd01hoykBKglsl/
GaLhFA9xgvY//dysKRlAQj6rr3UhC8BUkj6XY0IagsS8qZ7r7cXQVvl8JdLl0yaH
ycwZH07tKktkhc0597zgStfR0FzmEpS6v03FItkpJVmaHNBwsOkyfmwDbiH/lX14
/0J91XvFVRDfISXjIo+QKAqRJSMtA8VelIpav6aXI3AcsaTkUE5YNOA46ZABswiG
qC1KYtWxcdGi5TRsGv7gjAhLBpgXvkXG9vMsJ9XBmwiHHBh/iLE71LW4YaqowQzw
lFTmZ3xmpYSxPNFI6phR+FcEBBDOh5lulIAxa3LqcabYxiGMQ/1qmKXlnEZmui2G
l9sf9n5WNPux2dn/qJx/e4VBD7leHqqIO3Cq7KMPq11aWPcao7Pxtmn//gWtgC8D
173VGeEtlHK5m1uKi7Cyh+IiQLpewOdiyZuab47VAteWnB5f6QprPP2q8ZVVDdWC
HwdNcqstNEL/dYjoN2R1B5Gco/7g/zIxBy0ZDFFmO41Cop9IpiESBVwz7+1rCd3P
IgX6c5KkxKgCQsjvq5224ZlxZ09pWFGS8QZvZjURfIfNGSIVEdB1Ben5bBpihRkQ
Co3KOqD88utzNec2DqPMe7ML4/3D5zjmmMhj2gzVW6AtfPU2+Z0vxk6YgiLE9DMj
ZWwNAuZ1ybb82jB2vGqBMn4JkzwV54RdgeXRcBZVpObZLEP4MdMLckZ+ZAR5K8Tx
lrr3TkWBw4EZ4atSzTBMXvktWtAsnFGgI0wVM6wTvyNfcNy88Iuh8+xdFpiEprK1
3W8lcgFWssLcQnAUcyYG1ZxBEn74aZFgx2xW8507gF3OBAftHXKQTmFPIhehbWAT
uHGWw5NTI8DOEdO44Q9NqJm23oPdMqUkWfog1SKd5xN69jCi1mK8gEtwNHG+I74c
mirBWMEP2VeUO1yocXhMngb20yqRaqgsitjCZLsjOPggJhuOJqJBO9XnuCK3nmjH
OD/HwBSUozIHOrTpPgRzMP/WF+zBBHTpkj2uw4glG7VzhFnHaaur3QlQDt0j+iIK
YmwR8WvFdTJvHmeTtrs+dockwAHygwmLtgdL1V6fvKhbDQzepE/ZEG3iDTIGC6t/
Y/T2m00hLJvNwtX0z1xco4yKr2n4fJL3eANFgqgpWbg81Yh87AEdyMR+nlDvKf58
1gsqHjhiOZ+pwXubMtQL8dUTgK80R7PZ8JihSUJZV5MGZzWtZAeoUtbzglk1tQLU
1vQsPbwruEiAyqWEfdYJHpfwg/HBi0BV90zffjW3ecFMvFcp6UjKCpDIirNMguRw
dQK9BfdvMa9GGE1HqRYCR0at5MlWhpizSMpQelH+u+MMiJ4ulSdwg03UXEdC5qHh
p11f++J4JOZJ7tqKz0ZSD/e9FAyQ4JaagedwOTHh0ST7/sYI7FHkV52HMTrz+91k
GqBZEwU4to+1CsubTgCLXskb9uWyjTUesCb+tOtgFyMKU4IJpuwAINFSXjwnWSBc
jn5DDk3Ou7fRg75pbbVLWVWswHZgOlJ6+d7N5NLej09dxrt5K38Irc0ymiElq3w3
aHi26z8Ra9YGFpR09bfEf0b6KAz465x7RRIm3Qh8e2Of3mlr0kpxnMtWIaUpY3l0
ZUvFs8KmH24t+Xtjuc6Ye/jXuProYeVytj1slRmgMeA0ziVYOBeAvl3N69vSSZh0
1wc+S2K65chDB382aDno8D5zuTnOSZPsVpbO2qodeWmnif2FE1yz98Cvykz8I7ud
7pofeYvdugqNYclDckjzr2sqBpa4fo1HwenpRcFMq/AwvD2q2xwGyWooihWOEY/g
2uZDTCY8Q5aToUmO9IxRnKZSaMWGI/185u6++j9+UbBOrtkYkkzDtwqMq7RLKetA
dZP2aiHxbm3R46HbEOQelTBzlFWPwL9KoBMZUplaJBQovBAY6m512zrcOWFUB7F9
NFgfZw0ybWWVuYCUHjZC8oSHP4xT2WRpXSSYv2NO0RyIVp3G6y6IONx2CLQFfGcp
ZxRvEltnAE03xfjC7lcfAGYx2jgSmr1QjGjl0otK372E3/TsESkparXJ3sXaishd
l7JqFMcygw2Lm0VW4N2Te2Q1TDcfGUqctfCZAYjLG45dki2e3KmeQWmVlgPdAYCm
YjlMjMLUTSQepOPosAkQPKQheER/aO4Ny3dwRDWp/CTKrNmuO5SJ55PatpP4JCP+
knqODbXkAMyIPXRIQrheVTZyYa5jimrxmrNpBAv1Iqn/7Jzy6vOca5rGAP+tGaAF
MJKTtxFZwgpxdBbKkJWTDZWwmLqPTS5vdBkIPgkF/lnnIiJNP/Uhrz0lVVAvDSVM
Eu6d0DzhOiiovQcV0Pd19GcwTqzwnyp5IwK/L78XuVC/4eTV8FE1kdcqf8setzv3
PvwUzMBCKj1SWL+0Do5Yg9LrZd3yRQD+/KfVu63kFGdqy3tAkYLu49n0CoK8y9uX
0SIuqVIMvH+pp6ickzDZqKppI8eKcmmZkz7KF2Y46BjKLcLZsfuX/9r5xaBFb21U
qd+2se/F0AlayQq63rR3ZSke7GCpMTQS/AztGIdNTpwjOB6xQJ6cPslQC66AQTDk
JoOXbhWSUJFs8vxaud7rwxJNasGVyFObRCCZI9ACMK6ypxEuqkcdyL4vujGBmu3E
3fwUXf3bZEviUvIrhnm/211V9s4QTvHzJ71MZyRhJvvp0qnUfN7AOZYV/1rjZcnB
15t01VOGNZyo3qO0vmrUroCx4Qp1lfT9AlErMsMwXb3YgR/vX7N1r9UmvvG81NLK
/fikY9tdrzEO9cJCzyJPpZVB/gS97g83ccg9smCaOmaHctcl9O2qvnlUam0Eka6R
hdDus36aFSMlVmTQMtfuSCYxxIaX3HQ43YA+gMMDan0NXd4OA8Vd1NrhT+N1/sDk
sIT2pcSCb5UQHlNwOZ8ygrFu1T/NhaStCsBDMcZ7wuCpCDUXNSdkZeb0xxWodC5K
9ijt0Jwb+74GvipjIa7+eJoqIHuyDen98nTDwPI1B52QV+6feKN4oUc+6R7B26vm
ghZJdmIpFyOcIYJ6mYXNVslXYD6GjT6vVrYvUqNFgJUY1clo/GXnowTTXIsAJcD4
wHf2fXMyZrhNlxf/X6HfFKe9/+YPZ751jKoIWh4GYPvtMHNxKT/UykiMVlS8uK9w
uux3thI1UqN3Yg2GfK3EqHfApr0I3fxOw4/6FTosWvBxDsHtJK2LV7OOajXgcyVo
rQvjeXYvIukBjZdSNLU184Xo6/U22u2fQ6BXmfwlMUT9IUr7CX5L7Iiycpj9pWVi
TiXTcx22e6HAwAECBlFBlTS+hcsnQg0S7Mg18oarqCt00iYIbqFMmyhFPz2pzY1E
tFeSXqZ/sudCSUaQSqoYcMt/TbG4KInJsMw0JySQqDu8Q5EzLqJeDGCiI38hpMkU
UrnQseEG0OKoPpg7KflITvUjJiZLG6QiK+6Fh25qAfhhNRP7wgzzg3KhFeIJpieA
n+3uOlfkJsSKcVbfLIMovtRiOgE1nds2zL8XtMImLwA4Eb0GqVXNlgr3/cRm6npR
+PHk9vC9bFV36dKnQSq80tOUyCzlnUZfpwcSpBfEDW36bVZpv32KUpXaHCR4qNMr
QH9nnJVlZJ8+rLGM7l5ANQ56jOi+pvidAhVQfJXwRcNzNOXG67MWpH2u7ucsNzLN
jqNlRWth7o6BNqV+AerZWqMx9KJjA7/wmjx6LlEoDg5toNXT9eXimSVqk4d4Z8sx
/3JcIrieYo8EfgGGblx9cz4goVj324Z7p1eqlm7jdT6VMeMRZbdfBw+hfJAzYS5S
S/1AeFMg0r4BhPxzWRow8ImHSyu4Ly2G2elW/zu4moxEcszFkcqAVxahdU6/Sjlx
3DDIUarEkxvQkDFVRsLf5crZO4LgseCvC8a1I+CobcKeus4F/VrM1LZB2rbU+9m/
rEsKBlSHoXzPKcXFpWeRGcY9kQcgO9KMe+haB1KH2lSsu7Gl9a0ScCWWrt5ycm7W
ewlKtMpjzwPvRsaMV2M9zL1QonloEWthc67ouGeo86rkwk0Btz2ovxQRQi1baBH2
LW7tfw+cj4kQWYxO005UUymz3RpGyx8aTEOv5KKJXoOjxkFH9A8DKBVhhCNecG3r
d8EpQUUSuXBSPtiJaIvgQ3cE69fC4HeJnY1onMe0a7/ydNaFNhojc4X8osQo1Gb6
eLLoMcf8xO1BEnIr4VjSIRwbRiHhfDlv4q7/JER0QA939FiFGJURO7loxRLV9YN6
qkCjs/9jQwLDJyiTI9y6Bgx478oXlGta4FRJ6RIC6TM0WkKO70Un7O9FahfsNrJR
p9XbrJKqxwrBKcWqxh+/eEeQUn3MzN9xaDkBbDHOq+tkD83sSO7BH3+rhU7UgDDY
XZImF5HO3+1TgAs/EbeczJF+ckHoULDEtdehsLBnEXittMe3F3+F2vulutAC0qrK
feE3LmwfatxHWfRyhlDW6MemHCCf/G3/Lq76U+qgOWeU6qFRCwMG3zyp0JNQfjDo
fNHnXO0R7bJ0ZW6BSDL5AQ32Up8UaPBEIpbb2YM1i1295z2KyNAPEJFpr5CVO1Zu
PqvtmlZE7U2LimCJMzyEsBG2niL110w95Hqkv3qqvsvL4U7ltqjtJ3o1ZTazNJ+R
RFj+Cg5H94L7U78iX4e0E7OToqiadyj3hy0ZJ5kYH+Ra4tCW6uJtGyXi0QzZiJKd
RGUzmPZeeWuoorJ6bdxzLaSd59ZraGfcE4MVlGClrcUHQ/C1Ez7/GG0DWu8Y774g
bxFQTZLmeDd4CwkUd/ID6CFB0LMSb6jwDLIqTWBulD1Q5fKFRCmqOt2gnRmI0T0Y
Mf+5HtZIOmU5fUA4scYmIxD2JrA7Z3VtFlRH+15XNiefTFCRbbbV42gBN5UqduaM
V51XepvHCSaop12y9f+iJ3yVtxUZ0Gq/Ta7ROpqOF8e0LxiKPqtO1OnO8lgfbAYT
wkWADdWB9cN9zG9wnQeEvuBpomK8ZTnyqifH6TKO7AIv3NQKD8eqDmkOozK8PeUC
KTcYOm2Upy7gWMA6cIWpDOUBImyrNE0/CE7TrER6kjXUiKITDxp71VhdXUwyUc7c
31FSyewNw8XhhuOyGZber92+NNZrePHZjPNoy6QnaEbLTEo4rHXSZz63Z8HIykuF
clS6TPFge1f+xgrLzMpL2Ulk2/XkXNwAo+iNFuR/7GbxfPXOTbIONIV6SpeWtVdf
kVgCkcRVvTAcZht9y5PmLu8TTRKc88++qQg2ONNdDq0Qx31/Y7iTQAxHfHKCCymr
iCG/0hBATwk/5vKAvsZkKEGIdalFu8Xl0X2Jt/rH/bUnQ31R2oMRfiprZz8nV0lN
N5FZIaLTc61S7EMNqanu1CA4vC+2dGtyH53Aw4Xz871VOEFcOFB2ApAoFM69ZCKK
`pragma protect end_protected

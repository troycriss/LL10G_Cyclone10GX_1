`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
Hb01KgP5kfz6IsSE0fwwQGLaE6A6+hC47kWFj0JVFvZjV/GbisMe+q2O5uFMCoL9
ueyP7UNdaeTTBrCXvPVXhUxZxtMPFZRjMSQyxF6ge7mKc5F1ZaNoRZ/ixBkYVBp1
7HaW003vvZZhfMk8luOeo/EnvZWATUUI7VMUjaZnd18=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 476720), data_block
mnYnJWPPM9UVZoHFc/zqUKMXnk1NLe85vmc9yUz12w804vAt8tyyhvm3rkHbsOkQ
WuEGQJfpydXeMcbGzsePLikenMLCIJdNv2tXTbA8xoRLykyuf/EeDyv8BK472SVW
fY/wTVD69HrSctzQepci/EpaHxe4/a38LId6/nIrUxT9kb/XPgQieiiZfiuHIrRY
+maILwSdiE4OvtxBFdvl4acwJcc6yYY+3rwaTtFrS02XNhn3v9d3J3je7T0zc25t
U0ZqXuhnX8Z6Tuz3ry+hI2IzQ5YwWLWfGBYL0NEBglrTpQOU2D8LGjarBQJfQy5w
8sVhiFPSumS9pJvS1mL28C6csBfUl3rQSbu/rDCzUkBrTplhmrQ5Wk7HgnS2J4dc
IonPbJrONyEKcmAwOO9lg5PZv7/ty21Bpm+karXOx+wQhjhc6o7vpAF5rhun0wzj
8Y/A88Q7vRmG/Gg5OKDTP9P4ux0RPyh41BVuN1IqRK5GlrOUKJFXrAQs6j/PlJDQ
3Vs6qfdsxufw3wuyy9BDYM5gUIYC18ostulvw/XhZOC6kqcGOwoClJzIDP7eB9Oh
/RYz9X4ICjjwS7n6ALatZgFZxjYnfApMELHuNP0FwAJ12HG/PxBu2vMQKqzrAHf0
nBhwu4sgoNzSxol320BrM9LSnZRwOOhksiJl4rprnP/nchDfA6Ehyhy3LDHQzOQv
flmbU4+jNH89qTXcNsn1BuoM5p9dQgnUom50RMaDbAxgVqULuWQs3W1auycepQWT
9ihwIJNAMIo+LymrjNBYLnTEZcF0RB7j+obX4AuhH6H4C5ijCwgbsKTJb6M6X26O
6PjGo7XnC/OyrHnLqIEEmMkFz3YdXSD+V9G4jeFtlRHoGkwyWWfZaUHoD+BEHPt2
LzHlMgxn3LtnPfNIe9e8DBW06L/uhv8veIXT+gznQ43eraaXvh+YRx+kzkojKNvk
PEOA8a1l7AaGBYirU0rdySPbw3tVz3TmB5bzkOI5Bg9MBwj8pC9lDr9p/edadxjK
EU7ULxZW28+aGa1D3Gd9JtrjhQY3npgDKIKEWWxEgwnIV+MrIwekSgt42knLjAkL
zTDY0ydyJ6uQSa7XRQPfyaj/Iwa1Cpi2v1y51xzz+XQGGHbsKSM5HAB2eSbiAmxF
MkVBxcmzDcJrwUeVILs/4lDTc+/hpQJwbjVW5S8/VNCnETj8YgQQWol2VYcJIxz1
8erH8yZ+/lYc7bmpDMEWC81IKEPf8f1a6PxWzBXli8x/qKhomTe4KBrCsIJsvFr7
Fea3DwfiratQIs+sbc4GE15m7WH9sH3NnyLdvSDBPbtoP9FpKqe3tPqRABHQS2vN
y3DyUnb8G0fhM36JGyYbP3CAyIT4bTKdVLTUx0TZErgN9kjoIuUG48DGeEN6HXdn
pvCy6mFN1D6hd8HWZIHtcreQUEmq3OSq1i1BwtKEhU0lFrd8XvjRGu4qDGvroqvq
OtPqLqkC24RZ6n50bW0xTMWVD2kw2JmsruyF83BtTPkSlCur4wdmXYrkmFtQbn+9
uJQrNLuch6ihB4gqYtRkOFKJXlKaBvpDiKrsq1VQotsCZ0zD6Vft+bXBMBAsFS2e
GZYNQnY/33oXZQJcpWt214HWm8Cc7FKMB1cLuTkL9DH1qLfwSXIvKORsElP+ccZq
T+6kyllZkbzlHdK0uoTFv7CAQjCibv9/P2+4kOkTfEcb+cyQmORmhq2dJJxf7/3x
ez5hUmeBAPX1g6LoSHcMgJoES4OeeH3mdWDzhtM8iw6d1g8GVT9nziY4TTJxU4UJ
jipJzJNcA9Kbwhldk3l+1N3fWtlHm/0i4JmsHsZSQVmhbVv4F6CEvhjDjOpQAOQh
pXGhvH5yb8EfaWBfpaIj6RiiR6GvhJoGqZ8M7wZLfUuEav4kbyUOl+vKGJf6AjJm
B+vxLzvHHOAk9POpUqWT0l0VBgz9u2lm5CmM8pfrgKyC7QDP8LrQVCcSzP4kNp1I
kQFolerCy17eIih2p+iOEr9cS45y1Ebv9p/Mj2cagP5Ny1uHX9tX6uGeCejGh2Bw
uNIsDmridSMaobb57brRJXrc1VRvVf+MwWaboxgfcl75EUtCqUTfU9MciYpxVVeY
mTfI5hdAJWezoyjLD3qBHifJEGyH5V4tgGBZ6Dl133AudS1KL6G1b2l+fe7qz5DA
/IC9ahaYxxss6oWQho7hBXQm0/ErzappdOGZsU26M23pax+8FT2koHXZ+VWWHrys
cvJeo46Ln//V+hrXyYWFhX2TBhhW/fiPJnDxvs//fdOe6/jjw4hcP4vnfo0xk8uV
Vu+GTvxQ7awhgKEoTsoymDzX55e6BnJ3Sdk/QD8GEkSncNAWNMJk1G/lpWMlhgxT
dKSQM6ap8kyFTdeU2AbVYoUaAp99qguwjtrYyCQ7Zgd612qO3RRb6ltfTZGHqoQa
lg+HIBeIuMMINK2DWhkqUvPlurQ2Bja7va0K+Cbs921oi3Ezra91+AC1hTMQY3yv
JGel5VCbH2Qz23Dk6nBVpRtVWdU3N6+cQjR04HGcAhVnLySq4g40FUmAaKfSGyZw
7JTsDAe32qckOFeCG/kmguupdrqH7FWDC3KRFn/4l5CMQeb6D/cpg2MJERVpcJbo
sjajxFSVQRCrmqe8k6IT9cJClfWwcka2rIPoLY3zpeDBpyE4AQeXSk0+G0r/iP5k
zFU+EqsDkywWC+81m2vkyCN2V50tlj+R4/oPWJoI/92vZqZik5bInqSaBeIEbYJF
DM4YBECrsrMNfd08l2JA3dnYM/U1VLPiH6vRX4AryYLlgO0UvEl5b5wZhNtqJ+dg
kUjVzf6YzDZanrvaxv6UKp7slx25H4l2lYV3CfkL1SkHi5nKZlGjpCD3hvBqPWPV
4y57a1xRLxadPhnjC/FpnC3VR3jabKPVFBliLJLhCIhNORhv22dObNuWm8EeUg7O
IwZxQG3HjIyVvoHi8O4OQhjUbhuX8mML2PzUvkFfEJfzYcHbAfhA5SmCETzBEGhF
64pqL6/oB95/T7HAZoYMfmvhmg9Fk0q/R9PSyukbLLY+fHHAuRaNaGo/sEerMzcD
rCAumumK65o4IuMDNjiXTSaNxV7Ih+oc5WssAo2hDagFtRwwgNbVJkZHzsOaZP1m
lIjpJlPzXEvvpEvFbTadeZfCnU8c8UCqVmjzeVlCbqiJ9mrVbQioAChWCNmzY7ze
cmyRDk1io4/JGD3G8NTCQP/tuaogYgrs3HJJKJn9vR8RFc+PRMah6HcpdNnKW4yf
5ROKME8cQfOhpV4u/uKjGSwE3GoOZtTARum+IcL3voAcvdlc/nmK2t2d/ej4SyOK
3HTHtMHAQQh7cSSKevDwGdt2LuHRx+x0hzNfM1TyH/u/mFcSIww9LGkJ3zA3iRn9
6pIlVdAQp5d2UX0y5jqfyDS/2B4MR27VpkZUCAzPZtVD1AhPNUs2By4Kk28TXHYt
T4EWPiWrt0eaIkN6XHCfBsChDgBQYA6T64VDZ1HFR7kGkmQkaqcPByIYDzPzyApl
uihARTcLT33/UbRGo7Ju2gJsR8YDY3hDUkfRzUF9SgmmenwSO0h5ssd4bkfCAnPA
TeshZam5BUdjNJ8U4Oo7v9YQuJE/9SOlJyKhr/hiF8rBZul97nTtRzbNjEnpkfvm
i5qRIMclsDyfQlSgzhKHHUxf+RZZutcrHAxt9PmlEllQ0KQjgJeOdYdz4DV4HnJg
O3ccfKWZ5GkAZBx9bCR8PJmYC4dpfV+lDKQy5NIdqlzOGLGmcyD2kQWefWylDoeI
09QyyOwLAcd6EeGFcz3uXikP1fCcnwoxLZoR13iw+eI7Z6mFJMPxeQMsaGdBod2c
AibTzT1ebJvEnof8to5D20nyziDALluLVwW/oDZYhv8kEiWFDc8hKnIDzWOvbpTr
0ZxZ7yrRXm3unea4KSxsls2IW5XH+YF3/1J9vjwOlQhVGhm+r6A0ZbABe5p9J/Mp
iNEgg33wniyB0MZJIT0ONboLiUnxSfWPn8Sz1kwTo2CUt1DLphf32yaqv2Yas0F0
0VqBDolzYsPBQNjaRxP8swEeR/Fzgsd4iArB6APih5eVxO1/AWvAhbLs1qaIpR8k
8wLZmPLMsmOaffqPFz7K4IudMr6CJImlUvWaZ2q0thzAUIkp2ipYGdHRh0I/+BbQ
FqVyR2x/hAClLD14I3GE5ufhXb4ewkzsXNMxCTfX50BiYn8ZUhTl6oOlbAJ+UZzr
sFnOqbxWWjMDjhRybs8McC3I2ken6sBJM3Bnsi0mPmhrX/qCKB2GRkDthPfVDZnR
OlH9aw2qSfdNTwOu8TqYFvZRtgLSDX3UPCbIZOyK2L5I8DxNk/eEJTfdL/WdtjLG
OCRbNoPRNrg7MSSWvq6C6Nzgfcht4oKLnHbazkJHLf2qi5qQ3jD8U8MY3XX1Fm/P
xrqXeeEI3/zQJfKDceE50r+PiJLJq4oWV+1mse5snX6SaJE1hnkwQYoV2O7Z8kUi
CoUxf0zMDVzFGPCFilocBe3DAVrkS0Tlf4F3uwnCn5HBdfTLtQn14KYyBH3SIqYH
i34RltW/gypPV//KpHrPnlPr7jeI4TLxQWqSExc4v0Mzw7Y0YDEiaXod3s0rjVRL
BVzxAulTC97M5tju4qMU1hIFRmVZQ46GKMISMzIPKGWR0+vHRqsZ3Lii08lRrz5e
Zh1FBJEiIEQm+ySnkgx/Y6ExUC40HcfcAellPDHefK4fMz2F6U7EOGvL8SAS2m+x
5ZCBHLn9fj6pXAJumVqPQ+YqXhUCi8leQN8fapfKEVrcuuUGWy43+K0U1H8eLJZv
MD0pyZZEzP2pSfwY7XWx01scgG1ThKV1FU4eZEHdEgw4WAbPOhq0ENSIYXo4tMNE
26uTz0tlgq+dNNwFWEMcQ56QgpKoLnH5nwsv8apoE/4bQF4tfNzDZvmVRV/UdS/8
gmbgRNyfiMPBfS6NsBU+XxI9vvcUA4CQI4a+PrBm7FtVlEGljJXYnkyoFO21EDgU
FnDPAU7IEXPxvvV6+eu7IrkKOAg11hipGbDBjNeOWGSfyJGp3L8thGzb7vTWyaDm
SqzSqazNqOgYtozftP7uhrGb2M5lmN0cMEuUvWB/zCgtfFFQY8fY2x2sAQHjiSPY
1nx57exotaR/yzH8qtz+ZjvagUMfTVgT0gi0tbBsVeWGINFXVjJRpb2xXDmDPQmu
xReB/BPuz3h8DB7g87iJbHBg0aez2yXJXsd1/uLcE5xnHGILObJrJQTfKgh0sinh
/KKwzT2vQ7tsT5dXGZfTGrmuPnqQWka/+O/NAQrXGdxm2JRGjDGu3WaYiUiBxtJ9
rKpJ58JvQyQEoftkbM+hhvuz0AXQWLtbBTXtN190nljPBC/O37LPi3dQzxVYgoTL
ZQbVDYFYhisthujoGgiRYWlmQXCTv42XYlIBAVKCNPwvSERluTF4cW28d1R8U1rc
glFXcSg54h65BSQx365yMdeTym1Ts3YGeI7M2H8GW/7YLzlPsf7uISan8YD/NheP
5u20N9/ryNq+tbPlJCmXJVPRSTmjRE688xhu7BL8I8y+v7MG3Wf3eO0fu52FMjTd
Yr28TXFSZnG/mkplNi2umxZQ8Qk73oAwFhGl59X13hEjLCmiysBSbv/P6zkKkFdH
Qx66/yCcdObXTh8sKc5sMpLz/4mqmC4198fdw3pcr1DOHkwoxFmd5BaJqcInk05s
GEU1+DDfVIusW19e/cfeLsqHeNP+fUfyvFkAelDnYfRYk2Ez3wHeEeyxDO5v01Is
vH7Q6DtHomjiuWfL+hv/6/Lkan5uMdazPmEpYPiqLuPwMcyCcf4gbzeZ9iYlQJjV
lKafS7qhx/JmRKbjIlyzLxilNoej/A2bee6S8YscXqvqpkA8ou++owqjFsIi1VuV
blibNJudFpG7DXac7zQEfS9WBdjta46Tz4HtwW8QpB4X6GVFKbmF9/9keIkTccfB
hDr6fwCStEA7VXphPeVBnwiZHP8ShcG72jAhwzTsn5CYSerjmzmOq9srcEhzC0Bd
BiHwQJHIqNhh5izUfyL9UvFBbzxyMtgMt89RNIuAG79sxifRVpTmrOrx0GpSoqcj
BFmhoes9KXNU0HwyoojVTnXutCBbmsOiNjW1t7FOxAZhjNLaKMSiwcNH4NyMhiip
MfNQSoO16AmQ8dnlPPCji8qQhO4aLIBtQbowaWKvrWnf6797zoCqO1Ci0lWNr7kC
jwiqk0bIY9fnQHKrRNda3JC4oIsOHYenOF/CwqQLZmVYhpg14QJ8LiQA9R+WoQlB
yqVgfbVDFqNrU6Jqk9oCXA1eQtrp4RdP2vWCa/orM1VANuQQsggkxyc8WWW8vuxF
0K4GgDJwtcWsCz6TYSsB0zD0SYhoLSHsiZTzvoGJh1JR6WfPhEcLvlHsTmIbdeM5
gJOHF9/FzrCVGExPjMv3sLFDVS0jqLCdNgkDvvT98PpgRvCUIp1LE8Y3/ooGTnly
REHYDvUHZfRymRoYDctkQ8cO4u3tDdEK/41F+w8txwRfwBlt9JIf4/JAolhbnAsT
/H4lJifsP+n6gJ24sd/5QhvnfJp/8rnF/WQOYcbUIQl5k8HYqYfsegQNFteytgyX
kS5vYbpIAEYRLvQbuTVp1SE1xXXv2LkJlNwKrKFCAwKG2kNBhNJwn3+spmtnlPY7
eOnB4Hg3b6NWBHE0+DxQppgEeJ+lQS6TXtm7kMGjlXKvBHHO+kTyGIPl8Ab95cv/
98pOXyK2Fo0+CY/p0JUafr5Vhs/Jo20zwY1Bjz3bubc1XkkIopyz55OiImMS2262
ymFwNggFg5WpS8tS//mUUvZ39cX6E37MCPltjnem+if5kj0tcxXueqHqgxfUUoMi
XMiDEQKaXp3yXDzRiaZa0QH68o1nQgqeXAAibFs1SZ/p/SKUTsk74aK3HbzwP/NP
TUpY9NVb/Ml/9Lmw39JrxFevud49BSXibtN4yQMPl2UY0qxohuAWZqxUpK4dTEW1
HWD5qKbpHnpcT4IYc+xrHpMWtwZjyjw5rmphXJyUUObCENRqg6ae8JM9gSxSLQzM
FT64jR8zV6B/pTdf4bvqKMEVa16ukkBgjG8OtvW9S8jDZsdnS4/y7DtyJFti/W0r
UaM0+skYlywt7e5aZr6FTOEg39EjyiNPwCUa4O+1h6kSLmUh/HsCdchdFhy59D5g
AoQga3+jSl6KlFZbnnOskZ8y7xrGmW80KpyDK/koGKMAdCTbp+wa+JT2jwnCJZQL
u/MhBcQgtDj2Y9lvioY3melvIQcZdaGQfQuhS1z2oLMC0vAAw55Zu7iVDefRPhqE
ZP42m5rkzTx2kh9Yp4lYOxIeQyZd9aBcTZaMvkQVuBW4e/RUDyb2/HXCtargcNiE
OvEVmMBw2fDp3/Ahy9CqtdfTCbycJEUps0HeC5De7+ZFqyPa+3DfjfaxxnKAXOq8
nuIhQSY1pOMqFQr13KBwB9thZACHkIY7j14J5c1MTbI7aBjsgzJIlVdVl5UunZh9
xgbyU6+QrNo7U2bQB08mB7T3aRQCviycmrSQvr1EdsIrznYL3q2qFPx9QV4WwPZ2
BIN6Q8g+zEL9Pjw2G16GexfWMORE2FmzbFvTmLdz+zGz9sxcSoDcFXOEu3Li1OLm
4KdTsdnEWoB8WT+ZFku+SUj+ldUrxGx8SbJX99WalSiMcIcHURgb8vNlMBmez/3x
pYlhwVdcE1vmvIY4IXDZpZFQOK/01zMpclmbRjn68MNafvefDokk/tkuMHqq3nLN
86TOzc9K7HP4KqlrVctqkDoZfBCnGZx8FHLwwYAZGm8pq91rZqlbuuE40p4MEd7L
ZFy8a9L39NK/mV9lQoOzMEVIyBLB7Z7r6V5uNwrKCWoxso5iPc+a8HmQAWNQA524
WIUmDB3ytmGTVoMoNChXQi/SLMCGvBHDfvoIeiY+Ohg7zIVRhxGfmk3x4/4v5rfz
EpVPoiw9cW1gEdvz0OI+WK9QgBpVKWaZv8P8EyHHTS0b+gCavsa5BnxP3OcXFY3y
L4A5U2eWvnSOJ/B83L9CSfXSWM62Kgd+bz2UfQ6/bcTGWzKDQQoXoYWlpNPzvGbn
7lXvBrGTQD4N56V0SwbLmqXTwUdGFVZZahHiBS6N3VJdDNiGamyjQmqPBwlNTj0F
S2+Hqjckjc/P6cy0A+Ifqx3tua1/0HrA8xEusxZ2nn2kfg4ro/8o/HOsSBR4wMKt
mfRmtLkSemIDh8TJTUwaCYH3ElRZIgFA6i7BIRMQUEQNYdJsEvDrnUag1yB0W/wM
mn0Ot+rHpy+yfkpIzmhCStRfulkVDNmMnoGd8BLVO22fvKw6KVKS1h2wimW4vg+U
S13jzMxpMn6rlJjuHopZkciBYdmmH3bn83lpCbbuDJv2AbefNKQHQHy5Q6vI7dNh
oJCe9HT6dsZ/84KmorMOA/RLbvA0GOLnRyPycmULmOudV1dPH26wQbFPCa6GcnW0
VcvrfUnPFF/e4v7LZ9lTIMmEDTPjPswsPRUC+yhqWXYYFLdTsQJvE5Le/WbTyygA
p+twX2e/OgBGWK1O40L2CM9WowTELhzx5spLTamgLGRITOpxDz3Pm+UqqmUZPPSU
psAd9+5wFFdSyeRWGQV06QM9vlxdJsAuBmLHBpu/sybcRNdPcK204oMB1Pi0rPek
qFnW2xptMYwzL3KDGTMakxv09FWO22WQn8b0wamCjQ9HUBzhrajQETo5zyjV1/S3
/Ue65SVIdnUIaUDat1+mYbXDzqJ+lCIEskIAgzIGPwTRcVv7iQ8ttNyfF5TbuyVq
6wbINYrF90hYWBb4Kl9g0xI9by1vzPDr6wFYv84VKnJ6LcI5rOfG4HE/8z/q3TEs
/x9ono6dBVHVXHh1Kb0H9LYUMG98HZugJs9rTSePGCFJhVAj68ga2a9SEVyJDn1U
PZApvgMxTRt4J8nQB3Hb9CD3e/kj3xfYbDfUrvR8tptS/CbDttNDV66nb04LBsDC
8KEH0Kj0xNDyPlCPVbEdg+mfcqRmIqLUzY3zEdNzbGpMfZZn0WbJw0e+EY4b/xt5
yLOgembzYTuwjCxkc1ICsW8N3iWDmdidFX+as6VIDPGRBZt73UcgKILvMQLohaja
VCNnmZ6xGMNHlc0e9/PdqiVorm0rr+es9e9TkYuMgtIkWzIPjUl6Lcf1CBvdrCJa
EfeL5NqpvB2QUoWVQGMqQEFBUfZkkYqshX5FARzRrvKQstdklYbYdrJeKQg4WD6q
94lKc3TiUAdNNvX7+ia/jHVrgbOjoncFtzCBrkNy3dscL2j8k7QHNRa+Gs1NDEnU
lqoUv/+s/NvUGcaO+qUfmDTWmirmfYEdEgbRKLEe0o8uTCy9PpMwNuErEwzHHG/e
+tOS+GZnynvsp2r8Qx3JcDDk8FYxWsxUAqnVXO6Rbxbd2mml5tnwnGyvxzD/jz09
YEcg5cagMThTk5hVK7nDP6rMGSJLa4dNtdvrdYiOdxL4rFcPkLcTYelr7uukuE5G
Xrrm7n3Y9Zc4vqrBsy2NWS1r4Db+JektCFxiMY55OHSCNCk+Bo/K2K0z3vIU5/b0
FTY4ylyixQgi6cixrDplD7Kk0cuwGCOpwhyGlPfxyQkGsqhlX53IGADqmcgG1LbU
hwsr9LIbteTr7z3cVmxQDCNLyKeucxW0gCvyy9pQYNOvkB+AoQ8k8Umw13uTF5ax
/DRWSJFILoCSJrhAtoh9LA+bXPSdzLUxCPIBhjIWI8xUe28+X5M961ZliCe5KIOi
rPj7GLDXJtCf1IT/uCi/+p2vjthRqEOpP4r1/AKCdMyhqUGfcYZocY++rAC4bh+Z
xmX+O1W5W7gQvlJibRcP7VVaTIro70F0B/QAGAadKwudXB7yzLge56agtMshLgVj
UbPIW9lauMVqD8wALnBsYpmUp8rMzmx6xDp70vB64Qdmj23qh8/rKyKNWAY4+T8t
88RKK0AUb2NDELecn1uOrdkeKBMlgv0GqnPIwcl2wiwsGzUL4rHn4qHPnw+kNcxp
h6Nkc+pnPBNO9T61ygiW4UI4UXu4yCEuJ+nMShIusQTUOaHA8WFCZF1KfUwEKAOK
pZE3zNGF5CIFDA4dXZgke5LmIYQklQMTtjAi8eT5b6KJpkuvmWarThKBrh1UEcoI
lMrgszKkYWVOOX1HwDnwfPuehEbmOjI8XQIC2PmQSWMvuT3UQgHazNinlMywnTT8
ChE+TAQJCbkdGYwpePwawhuHbq21oxrkYEw9jn5PjHm8cJEm0DuGKigREnm39OmP
jRi8iPj7wEd+z7FsR9za6HxuZhZoUSySo5Q4mlQtgtujliJftjGGoU6ZzD4f9/VR
6/VIFsBKSbGQ/vK0tiDsjp/pNamZfQIdiPHjDqUssx3CAHtK0HqMmoa/anzrpXSN
xhXICaRoTu0sYIKI1lKSoyqATvCOb4RrBFrMuj26G3xglywDZk8884njVdUTWk3n
RvNlDxobqObh788QbYKvGGQqq5pQtDjPcVFNOLzg4u+yCjDG6cXsyRE6LY7APlre
OqbMRTtMe8V2jT1r6wwpiMEWJvPFMfwaBD9ga5k2ZSNLPHadFhbYmYqOuym419x3
VtmrWWvMla1nBZM+qapbQe3/WbFLH7l1smZJM6CE7cGE7muWqCVtjUtOqi/2PERI
bgbfaKuOMJZdin5Mwh9/aFwAYznuXj7GjfHPM+hYg/XIFu5kri9+O42xXNHDOvjY
UT8n3UvA0p7eAWWEOHoGMiYA/s063gBb4XxVldv1ER6NwXcRR74Jq9NpBHnfSqmv
aIgj5/FKPvMLufb8WdThaMOknOmWpD4tln1dC3WnjRBnleVYVPPznA305YECgveq
sOj8FNj4mplRHwyxiw8BD3zMGMNoEKLYLXPAkqSkTHVJqrx6ngr1N6ouyATwonVm
snzfKaRVakzVN4t7mQqY3XbHRAILgNF+RklKTeFvKDG2H7HYDKj2gfBRkyd2hEgj
f+NGVGJsJcakVe1EyCmnmfIYo0wdyxEAjXvqxu920UxAUFMdBznuWVX1AbU2GuRK
cF6VpVzVX7yv5WlVwLs48HPt9xZ4BTemuX4XTI4e4pHBTtHWH4B/mUo25Wwv+R6Z
GiTVNyWdLIbHDgu3Jsa93woYAE/9XLW2IbVbkmk7V/pfGf92GXvHevAkTDWKSrPW
vaSW+BJ0Hl0iFmaEg3LHOyfccrIxNML3Zm0ABylIuMlR/Ik1+akusT+DrhGF5XTp
nbl+Y0oyncVzrxTHbGQjRe4dzlB5sZY4qr2+g6j2ToRCvGrAEjsNbsJEHUcHWotk
OC2k6dKxJzLqvNfmoyF3sVY8NicSZsrhPw5dKC4y9K1oQLv+DIAupmRRpCPhBPhq
drlN8jrfzxeXoe9SVhlgJ/VQn7mTuJd2J7EcRStxiqW97huA2fvWfOsksO7ydgIC
5rjkkL743Zxq0k+PIK97uYDUmSj7VgFaZ38ehlLBO3TfrAZhigZKrHltaO1iT31G
SuuPXm1a66E27prt3r+6LwwvTkVjhs6ynlbHpltK59H3HZ75LFDW9olApPMtAzTJ
4VPh1aQLJudZ42CsMKbjOzfTYq1akkwqJ+kHatXYlobjtlz+jVNHnApiFkFCmkWq
xuvkTFiSFNbN+GWAwnDC+U0asDHxW+63op6uMkru6NIX76RCWqJO2Zr5KcYUW7f6
Ju6F99YMZcrhFwgGyP64QjWR8RB6ydSJSLcVMlESImScQXOaReffKNVxZg52O4yn
g6noACEcPkBsbpjrstYmttTRx0iqjmBUDyH3Tr0QyymtwAikSAKjUmdG02yMkSJ+
JJAX1gLrdR/OZjIxnIh+nzYmLjhoQd46e/8SNqcZdNGcBJOXDP6dy9Wuu/OOcmZj
8fUdaAnBAXjOUxPP9HE4PIBmh4Ra7XguosFrEMa9MvrfUljSWwRspLSA9xsJBq+R
LYqkc1WEMvNrolbQu04SMPKGD4Kbg7YxRnMbXPKkqNc71W269p2b+aMQUxIawP/q
gOZY1aY2mgqcyGXV2rQAYzLSoyt1sTNy+lCiwxGM4dbH4P7AoiAGi3PBSQcynk9E
cPNUurjkdu6l9x8WipOhg2y9JbTUJ1teNOuapcCyIMZoWtWRHCkBXDin8pEjhAUf
ylTC+R12WjKyX+Ocv9fX5M/1YGbtP/0r2i0mOPCdNvuylGxqP1fiaNBreksVtPSC
2vFFBz8ldZNAwAUNDCdR9wgTu3DAGpst3WfgVzrltSRx8WYGCP8uQoTNG/Uv/K8R
n8pinKX0MMXfcW+6h3HVZ5r515H8sdgK5+J6VN4gzQoUVvTUfABhBfRPN+J1XmPS
X3nmmLQWgUE9kjiRQH9oHh7RvDAVYDTcMczvqDI7zOh2zHowo/NQG8zwzNL41U3j
EH1ttowVbLT0yjVnz0mF16D3w7b4klC+Hzucs8QQBD4uE2oW41nZRPpSG/CL3DIc
noAjoVhuhXod/3dPNj2P1Oh7RzuM4qnf5iu4MuxpMAe4WoWzCTFVXznW03UA0x/N
0Pult3xULyyIaAJUTwb7fSy9Aul/xqclYlLjGU9oG5jtowzxxgifhbSlAHKyS8NB
lCo44RIIUg/HA5A0X9AtxRzNZAdue0jEUYd1GeNBM7YXiJAqDn0V1hKOrruIXOfN
SooY/xVA7PSC79WNzzXId89/drkpKdKXD6SzgmlZyezBByZg7g4pCH3quSO9TEI6
G12Q17voDdNbryzi7sEG7t0w6CJIF7SEMOOIS+sHVt7ZjYKNdvhy/8rER/oOvElx
VKBHn/EihvSi3KMDAm/9X4YbxPpxlm6k8iN/Wp7gD8yC5ru83pWJOY/a1u+F8Sgr
TEP9Tn0xmAqh7dOBgXC3Ok/12o8HIVrnuUjP9UDxt4YcSCBR4q5Tq71wsmb7+1+u
dJRb39Qxxh6mZJ7oqArjn/VOkvXAmHkXswLfnsw3EvvRVdvKZ+wjFUK7MxHxrFap
JEikEbG3rab1mk9dyYHBlNIoLU39Z/b8f7OLrW7W4Uy7T47u+4lRwaXHMqbQVJrj
P7hNqR/grPt82EXXa1gjmX0wlNlBOuuZKZrCXR2hlVOqHmwK0PAojFx8mVaKwUlI
UNdmtKsywx7K/eKAJB446+J1lrY57m+/OTsNlmj71j8eD9OdFpzNwEaumvbWj7hF
eGHXzRiHZnIvM+BlaymiSqLLVYZqGgJlS6RMrdfEhsIPgihMDBk2R10r4JA+tdRK
So6QIFvPYumQDZz1Nskn5SwCVufhOa0ouFqBTsEyOqhVc3fokIGZ8H/mewU1BeWW
Nv/gIKKcdvgHd9cnnwDkp1ldqpfkAkgmL5nQxq0+s4lyBLJEs6TqWDmgrM9DidVz
G06LaAttg7PRGY6+AkqgstjU5G5uDbEjqHlETYuGfntyj/Uit7VrLZWbtM/9DkWY
eP/wXCQTYXLXr8UembG1jeP9sPvyvKUvNtdGGSqRjjSNGklJ9YZHLIdsgaBseeHI
LHQyxbp22OYrlH80b+mKaRQwpBFxXg1ttqei5muR6j6Raz4NJk7rc+P4KMYkoZ2F
VxGvAdFlzPU+9FYE557ZM67CixWlGM7C1YeHVTcW3AJftY1Gw1SAVKZTLkzw2iXB
YRjBHPBrzQFY6Sq9Cxw8YgUwF3ByYJB8fUPJXrhkPMi2H1inlcyHgBBGAJX+VprE
k29BfAEZqT/YJ6bxt6Nd1jYTw0PUU3QW569pW+JSWJZKHFZNxcUqyqyr+z9ZI/Be
6fXPPZ2ajvssDybCYFTzIzAUyRnunpSp+ll29fvKaW1P3qx0idHhRIrgNcpTuscZ
yAEddEBSsvcZbM9SJZZfbhSoGHxTuDyPg73WJFxC59R2RkVEzRJuahJ6zwofyFja
7MKv9r1kYtrp/4fyliXKm2c33Y9rjsuebGU87A4YTmMj1SZ1lXCtw0+rIEC/AHAh
HwLVZ4MATPlwmyxMmmJQ+g5HiSB2zuir/mrJ5XYGDqOg7I7Knf3B2dCrXZ5x1JXs
FuVQzkKJjwNw9v3PejRTpN6SiK8Us1oaZiYHw4oi+GziHcxBUlBRhQW+KBphBMCJ
abBtNwZJbp0D6htBgjXZEHOO4eLijAcY6jivAANdSenpy567LTwMEpU0UOCplwNj
PzoxI8aXndl+vNgikjtVTaqCVgRgDskZTH24GzBsY74WNrWSFWT8U+X4ZG8raSkk
4AbUgu+dkcTdiruaKB+E/rbIWFqGHwqDVlDKeT+rTSnas06Enrc0jm6PM6pK0Z+p
Z+S1X+r0qS02xG5mgOYIdsdFqr8N8+Ed3NNoi90q4xruuiVHTo8oxfDLu4mPIgAS
UIzgayvJa6ImA58THm58JZiMKw1PDlbthTIjnPjVzDC5GYccLtmvsHkqqULNGE8b
IBZ3ILVPh++87nQ/bU+0deTuMGJ2UDgr8KRXjYD6QOrPIqdPqGIldfcdJ6UWZVYW
I1YIFk+9dS46ct0nOzdGmMe4QdWEqIh3wqVDyTppMA4i0pl2liWVr0Q6eqHF4QnJ
GevE6GiDaEBoGMr9uMu/ghd1i7vTwWXQNRHhN5+kBMNP5YIukxwjPmX82K3ikqc/
/wQCrQIBP6OCIhXf632GSbXLLS5pal208cu/JMia0PvoL9sBn6nwAd7lmOjmasCU
wjdrFLjsePqYuBUO3YgrnBqjQX/QZzOOhUhdT9NaxnI0WWRnBKl5zpWorqMbbH2Y
XTOmVgw0XNey9pEbrRGDXud0WTbboq69+0MYR0/Y86qAZ+DgX1sUquzyDPGgNzmP
M6f6uwwmosZ6ozRSfEF8lJv6GP0ybAkmdV2nTa+0KyPpIgduxfy9JOL8r8q3fQJs
phpUITiC5onViLNw/iLnjCRZRE/vCZwTYd7TZw3AZxZ4T8/R/bfds9urL83qCaiv
of7eEjV0yX9GE6CMbeDjAY9+PmF4asM6hooo+3a2MU5SB4/NzLfSi04ewlKRvfZk
4cra5hQQnu3934baSL88shGH39536cRrykwkQyLouuuWGonNzcXTBcWVsl4lKSwb
eaM0OnhBwGPEh2aTMOllZ3Blt+ksOZhVRtWtwoOT3UxEapgGVdaKnqLOKV+w6h4d
xI5y5L0QSpyu05m99KbafSdUcveYN34sq+qq+NrXvx/YE2uoVRS32jy6sR5zZuvm
USWcRkQgWyqsWm1tnxTn6In77K85tU1lZwPI3Gp0x2N3uAU0llQ127OG4dmcGP2s
iagzKp5PSDIvzD/ogHVEHATBPchGBZfl9u57iErPlSnxDuPP3pfURGcWMPoNxA7R
5Cwa//oLMVZah7llJnaQLJQP+q2cIT/8hTTPfUbAGfKTwKLjr6QYti9ek8wzM+w1
uqJq8x4tCShYGJ38GtGJSBsdhSU6nu+IFqJXc8QTNpFjpSBKKasU29Wbyzao/GTg
rEju6SWMYlxvHh86D352ozxTyXIhzqQoJnk9WAelDTFkCoP2YRn8Gh8TN5hzqm4i
ADQRfQ3mCbVhpZpv/rlmQoyHIVtbTeihvvFDz4/OLAoo5QCzgCb7a9gaJaYK9v+p
UuLw+PfK8CQOj5swVIq28AXqft2VaIxybgqhQB15rmIezLUCunPxAgRxIj0qJklK
zpgDi+c2KgS3wIVpgE8FzMwinb1yblKHB8I+X+w8tQKZhLr3rjV/211LQYN6VfHD
kZCzlzF1TyhKXWQyyKuYcHGYjxmmLXciqthj1OSa33SDxJY21QokBqWyAR9LwyLL
eZrNtheaodBiLj/NJm/gAuCLVXrHJ3HjbUdDCUlFJSDLsr4bT6FgRXJv67cnI4bN
JBkU3wB396p7od7fwIgf0yGwrD8gW9Io8JmlUlLaIGAZi4cI4bdGsWWPT3n0UGnT
JX3sDCbYkhp6KpAPEBnOEW0olrFhiKNK4+JZaNVTMDdbUN08AEermz7t2yLGm44C
HaClLK4c1/OaPbrF7CI5qO2+ce3nnNvXrPvolSsOCof55fzHB6GQXDenhFhqcMNp
xwgAID+r6aqXD/tEmA7STk2XhedaTG+b91oUb/VhcgXA4SNjDKCCRYwdX12m+Lwz
GsbrpB9M+TrGlKsC5ZL2O+JEC3rgnNAPw025w0UVkNBL/6VlrrKX7SHRveO/ZoTV
kup4KOc1m2MzoyT8cnlxoHTRse6gxw9pls4gYarhpOOpSat3PF25GJqMbPA82+uV
cS3MjXQ6c1svbKwRyC0HD88tQ8fLZgOaLl3J0u7sQmQ7c4/znW6Q1MmXGASSnWTO
fefng3n0vsjGBpeV7Ug9hKAdP31U5VOPSLDsn1gA+rOrxJWOHiKm0kjbjd+6Rn9i
JOylMHEnRMadP+BBf0rzk3ytCroNit5C2+0vTuFojol0ghCXQ42+a8i4pV5lHmyx
FCQJmpSZn5yjCHtBJ4Xfg/nCIrNoKFpcdylnM1hr29vdeyWgre4nOT347KCDdYXs
FX+p1U8BmfF3PmSQ6Uke1Z+t2SUmAR0oeBUGnpe7Yr7Iqj2iClu1P1u2krwLtTkC
kEGg+4l6NG7pMz76ha7lbu0F/v9santJxD2KbD1oTHALNpxZR78ZKGNTkV3nMtKy
yw6JHwSffbYiYd3mQoLlXBuRp8ge5FxqdDdnYHluUpd7eHGvTuSLfTx4cTsWNRug
k8/3KsO3IJd64SxNcYaO7epJX4pFZcQ3Z9xA2PvBEcsAT+g9OcWa6K261o3+iM8S
4xfLTmJFAPnKOJtszbJUxDu8pNg7tH7zXukxIgb+7+wmoTqfqV/gd06SVwdZEewN
4KGdOm8Fd4xLqCn1uivhXtfwh5DF3YxXER8RISVWQK68xxzklxaMuBQWGAe0EgVv
bdaDDhDtwOOLlWsJVxHme88mb3VCwfeIdHIeeCoG2IqUcEaHXKkPr4GEwzEz7nsp
IyOTndQLnlyF+BpwNk3f3ni8rDKjLA+MxBrXPGU+ACjveYiDmci1I46IB7Mq+m/T
jWRpKC4aWnYSN5vjNoHJsImcXwfj5MvOPOXGQJBsJ9Jy2lXO1smgxiWYHWczaXZ4
oQuTPZhTtpqlvEd9MbQWuBhkEsN5QU2jG3+Di0tIo4VaM6Xr1nyn2uvTU+qu+OKo
tTzHmSz8FlWI7tz+SmBKK2Ni+4Zbez/g0LtM8ShPqd32fIwcgJpiqh5r+jjQXD4U
EVnv0pyr0P1EHtzh2i/Md7rXdRBAkriY+Vl51c77VtrXjVnT5p+JiNM3CUix4rcW
W6BUQPowBte9+qA2xVuN0Opv2kFSE1wbYuhlpaQ2M0t1PoiY3/5R+QAx7WcAu3Pr
FbLzsHXgN7KnT0JZBmWQxPJyvHV9jF3fdo2FolPtqUiYWEerNciDtFs7/dabhgT2
o/MNkYwI97ARJKlVfkAVmZQE+LhD32Ptz59NRq00yg8dtD1CSzBKwy9W67/41+eV
WoLPyfLGdQWM5RWZA64kWZS8VUxvTF94Wy/fqdOUqfgU8RRqMTrvbSM/NQVvu9Rf
P0nWYXPnyw0Wrq/W36DMQAd3x5dP8xlcSNdpRb4kgCrfo7IJ+2n/s8ExMl1GhfDP
eQvv1+oCR6OIQmX3R5RvEUqCmnVCKCfMati2ezC0waEFySQwhkB6kc2OuPXEpSmH
DvuIeYo2vgy5Bg0QpbvfpD9SPzM6Z+4pqKGI6mc+LyzK+zw0WuRvpgS8jt8XXBTD
4z1HOsKrLhEn8r6Tn7kuGLOa834rpD1DZWEl6MA1WDn0agaFLYF+HR839MVwRL8r
eOdFjvxXf7l3CigPACKVriiT57qJ3xfFrXk1k3EuSL6rqnyDodpXU4CDNQZxAOGm
ODlmhfwgvj7fGbHrbpnbjtTOLVsujWyKks7/KJcr/Lcw3Xpki2gw+U9PAQTuaxZ+
0Ueo6aMw1BAfz+iKaBCjDVc9ZovCHzmQ6hjQKzx2rT/lmD2rZpXCjKRMTgIfzn2E
MZgzM0QLkusX+Y+BrIoQsewWzsSjNsguhCOnLu6fAhFvA5eo8phYuVLUxEJWzOsD
MKZl+7l0lswV/KwhM777OWfdzC/uICdCsMPDbfqae0DrTx063/HnVDMNYNV3RKMX
mMahYb7/mm+xy7rJBtlXZ+jjZiuQ5d9ZRIwfhKUOsRwqc4acPY1cinZEp7aZ4QyI
1PodMVXdRZjocdNnY14S/T/MZ2izaM0Ky6ubJB2P/oB1R1x5Hhtnc3FuNcaCztru
ZHq22hD/M1A8E0LVXMooMWcH7GctUoPvsjmZiwIDHuCWQtOD4+DVgoi2jAQvygXA
W6bkeZYOu05FY5koGkjO3e3j+2bQV1AQ5aZgmLsWPUCCmTlNM1OIEMKamuyyJnQD
IiDDGswqj9vlOBzphbzSPitfdht8APtGrJCxDuYb5IxWKW445SGzJkq3VO4mmN7j
qEUhdrXFEkxYlODt4SvsFB3H5V9DYQE21xswvG9bSavs+ZR7pcbxm78ucW9P8i7j
4CUM/sle5tgXRhvupp0VuZvjTRtoo4aBTNSDMJjEJ9U4ee5pf3QypE4hp+J4/12e
MsLwBEja2aZ8u9nej68RxtJUDzAG4MaLuKm8+gDC5eSQVIwZvVNdNBffqnn3RzNS
9ECm2bSXQ+XpOurKjm8uYD/Et3JA8O93bc1qzJLNd/cHCO1rdS+POP7xD2bRbgdA
OYNJ/WRrVmgFRDwZhD3lapnWmxFv/YiTpr+cltJQBipHVmMJl/gMN16qvqhHsmsy
+PMZbKGYd/c1P60qG6liDAuoLIPfbnXGqdrZW8EX0yOJQy35UT1LhFle0WXEYNE0
qK8fSozsH6AdgjtmzZj/om1z3HFH5wqEhcF9KRma3QUYPddCh79b2BLK0VgEIBLs
WKzCEeHrtxze9AqkIBQ+uz9xwIKYHiwgKTk1KSQET/7QjgWz02YAtxo1xCApVnjc
p1SouBZPDmW8wTVVy3kBC4qq1SmiybjmfJ8vZXFiJbByM3okDUU2X4dtNSMmK/Fl
/1lXteXl9+vEZYg2uB7vWJRE0ZcZU131ZXI5ZElc/yq8JvRNZ81RUlgqV8VbrzC8
PlUSBijWd0s/7v0BgwLUnMoyE1Ta1JnqiVPtlXYmSbPtvpICf+53BPhfiaj8PLdP
oMDrm4hdExSWtmSNtdNBhkRBifSLjf3DtIzsjBgY1uzhMjg9xvuJFed7AQe+bnfa
t4HKrFL/eltMOeri0NnMH83yibhvqvcd7Os2uLhp8k0Pw42Mz4NFgCC22EEQkNpS
UD1Fbs4dGA7StFCMKuDglRcfMYhbyYToPX8ZSW/qDjh4jBZWK9dIt3WE82eZcg56
c7Zu/Rd0tnZ5nwmIwqCVK1Z50QtXksyOQAihORrgUplvb6KZyL4TLmw42kAtX02H
2EQH6ZMeQ0W67QcmJzNhce8mOqv8iAQZXsVQxGYakkYcrEI+C3faYAIrumHBUS/v
OgDLEZfqf04kIcs7LIDSoKKHRrIEBavATBpWfhlwUWd4+3kinboSF+9ULVMb0lbG
CZ1lUWZ/NrvUYufK+scyQNhdthhcuez9Yimvb0BvmlzxRwacC1e61E+NJ3EykIzp
ds+JWRXoSkTXGkTgJOuMCysUmrCzYtCfqU0Slsc5ndfUfxpEWQIzDrwEhYZ8muZ3
Jr25tmZ5GJvMJSaXKTPZQdhtbbevzK9ozPNyjqq9ZukMHz7NR9+kE8Mlry05BwBu
JtuDhgLFUHAG+g67sl9fPnI90rayKfcIloDgMjCvOV1vucoTY1QxYBTgbPQ9cPX8
2FgjuR1IxKRHgkuW0T9X/2uQGcHtXWHIW4Thop6bmOZvsd0PzqT7Ke91mJE/FUhZ
pgTZTSdSnofVgM1W0dzdhMpY/vSy1XgVaPC3cfyq+v09RqT9m8vEPxHdTFx1N+3p
U+Xp+J8qGg5xWtIUXs3Rudz4rBGdoGMjGUP4nQoDSZPt6blbSUllCB99Ls8ASRE7
++7Vgto6rmWyM4jZVeGviuHMyGIuiw/xSQ1f58CO8NlqUA77ifIW/llHS25z42VM
jp5nbcCeInNh0omTY+vZ/wJRJcwOtx/SrBjMVXUHfW6FwlNZyVfnD6zjNVL9K/W3
ElVExHKID7G7dRrAbVmwi26xqvmGAvWRu8mRpbR7F5vEhHR/cPmUXdnmIr0aOP3s
Boph3dfrOQi+BBL5tapGvl8PW0MoOHTSy6uHUPFIZl6QFlqGI7Ivxggi3NbFOgJP
YbqJy3bJy3f2dSonE/S0VjaDi87TFw3nuKAxhQ3Is4P82gAgX7n7cZT5UMcHp2I4
c82H6wxLwqXQ0YWHTT6X3w+S/t0eleAs+93ptjplzDN3gVvnXKlnY+qORIRRY1Tx
W68c8oGTGEOW2tZCvmFrjwpVyQI2FAaug5+M+ecg2ryZuApwNM50A1HrXfIProQC
dZICU5VBy95X3Hf7zder0ygrQsenneGw/zs4FSKv5xqcBHw4P6S/PVEU55idG/hS
Hy9m2oWiDVn/jNQoxXPt7U4YLE6ZlVTNQz3LJYhgupEKjztsvfnEjHYu3sCdaaZ+
NIG1faulmmVgrohlaRosJNG8CgzxAFAtXnCWc3jKVlTab14ysBMnYsmi7mNw0EsI
JkcHKHEh8sUuUrK34X01p189RZYlaM1NdUZkGS6DudbvntXMQXCJVeGcFhiYOWdW
WWUSrg0VkwIittdl/OjOMDMW341Mw9Ih+jaj0SIGnmtPPyVsdaV7U8KKR6/Ogkdt
ZUQsOq/QZsHt5NQNKtVElV+zOyGnZT4lHaWoL0RETvdJ32c+wItEJc80AexP+M+p
fEs8ierZ+eDr9ndi9bKqB3nRKSHMqHBRc/pBjfQnp6LK5pUcwzvRPlo0FDSBhTEp
h9RlRFdBCPCItdZdRflSlW+0+zGfsVcrSZzWxKWk3ClxOWLp36O7dl+qu8qoiutn
RlCr7kt9WrGdbe+tJHIKahIIL5t3O7oe3tuQx3D+xVG06RElKefbGh2o2MnSRRBR
UiT4nIPtY0/x8Secer/jeLdhhgPlnWk3k/meezFbFuL0tyZ/shLIEutVIx7W5o0G
NDlJnMMCmV8Oa6VXmJWdi9CDSpj+DuKjBdX4CJRyqSviTas+E3o7KK/FDNjy+iCu
ZrcDEtPDf56TibXdjyGw/nNPC+pecFNIjAsILonfwJifb+CsX1JJ6t0PqV02agPQ
YN5vY7B0/CjKe7PTQk4S1jVyLdHlAy2qVcKTU94528ny0WzoH3KJqP7thIt683Nf
NdKIIC8z/OSJjnKoOexHYQBpv84JC0FfKa3R6AZ8iig82+2vsIVeJy1wJoayzWnE
8A1vScSUIqX0cT/sc+/tCGAEJjMDZ3StM/kkQ1akJOxewhS4gyECPXAmBIsMX8LZ
qWyHYqQ/AXzLhGuiXFpMqTlIOtYSvOOG8Ii1nS/onlfD2B02tn4/ZD3ZzPn2H5Uy
zH/OXOn7jY+SBsVShLo9kJ0UFNMI/hgkQl0jQb8hQwK6AB7q1WfNVTrm+VeBFI6k
EUSTrz1yErAU0KoCk+Vc6eux1v4mYGU7QHT9S4XI7hg/vZyyg6CpOtiT+3N2cxc8
YJqrtNVGHWNXhzyydHGSRBbbOiWXjfmEGc2/A33nHRcOD/JMY6ugoGt4Vcw9uoYL
I3kGQ4cz7iKxizgWycLvCpTYxaGj4p4FcCO6ed2Euj9V03hauoI9MnN2/PVFgFjx
p1d1pmUZjFAeqpgNUOawtse9sG1fo5MkJB8WqGqHKDnekkcPWPy+iUfOEVkIcJVR
R2HqHUiG7eYeFAwvrXgbcuIULdA46PQ5cYae7961kG4MIMPi8q20WBvumvF3u+La
TN9ylIJ9xVl0RlmvKHVUTjtPWGpJSw3t+Ra5HW5xs1Yumy1U01B4hxaFS5UMGXQY
vGMlhjrAkCrD2milfQzlYySur2lOC5sC5tSXiXgGCPbc+Oo2VsNd1tMQYg6MSTGG
oa1xK+ExJIYLBHA72Ppti3vWSImh+tSoHikGsib+4VOoQFGK7BqA4gqvwtQKBkga
VGAMc+FMtqqfwszohyyqD6K1z2xrFj7uCNUB6wPQUe86Iq4sEy3gDXuHfmsiHrjW
bMUq3dUiCu1O5Ma3gVx49A4l3b4n2+DzNIrZOdLaopLG7cR5ok4g6d9T7lE8APx6
lybO8wvu0qwoYIR0ue97t6T1aXXfoABYNhkKappE24FQ7AI1s6oGFsaZ1WxEDHSt
1KMZ8rUmy5ph4AyOpVnYtB3vMAVSL3grKn4bu5YZtBZvMeX/dF0JcIKzrEe+V5+Y
18zt3hnQPsa9kbKhpoWfvOBFHQmzWCN8TcNhFZhKo+4ja2RujtetgI803CH2H1G+
bSlRRs4rnlLvHPuPeFvybFYa8pI3ApoJNTfMWibOEg7gRKCty1csVJDYEvU75le/
FhVRX7/lqKenUcnGIMZNNTdgV27kT4L685ANc1m8xh2ONHuXA3Hfr4pgTqa1APAZ
oGx0ZDfyYf5VpOT+rcGWjPHIfL0EhZrJmpmQJP6W0KlZXqUBty4BZeAzuXsN0zRe
FaQHLpkzYCZXPZ04FAc5gO96OOff0Hndc/G7gDpOi7jDWykhrxaOZxw1nrEi9T8H
RiRvCRxrC4VcJHFfVglXaJm0MEKzUzyPiq/ou51qG2qUpTXftdUJwv7S7w3FzE2a
LgIyTmWL4952BEjEmaeRtuDyrK9Xi0+UOaBaikqYWTt+XV6NBLDt0fO49ygZ0+/A
81NBxJwEBVy0nIsMBmzXIcaNeZyKVyko/HrKUC1t1d+k3qDr14297C3EqvGXeChm
i07BQRmZ/FaNslCz7PT3SAfRQjvZ3NXRVAwHUp78MfhdUHAviVNjlvk9uHoKLUVJ
pPKtLkD/3QOLDT7NNrc2wxdm2Y8xtAeHTlAvnnl2xHWoxDmQFLtz4AkqrmXCSef/
usClnTlQr7waCbH6kDl56qkO5ldKMQQ2j3vzp4209rG2wL2QiW38B3m91G4dlum5
7nzB2cNG3WVSXiLZMAe+fUsGKdijfKkU4T74TBMuUMtb+MVGCWU4EVMsiy/oVDLn
aZquo30GaCRB7yZ5rdhKAHFYVv/wtHqb/mt62RpXD/AC8O2WZUpbNqj49GU7MikJ
wiO6Goa0k1NqRaldFkM8D0KfoicEz21i4OSlYfRIMcb+t+P/EaA7elvwR1dhTylF
8Inufb3r2mTv8bVs8qr/zL6QLM49t5w40ZVZRrhWcPQBvK9TqV6LX6VB3Cyfqzlz
b9rewcWfxFkn/vox/afSO0VAUIdwuWLn8sZsVzp4K78KNNKmxIBwSY49M13OfP0d
2WNV+6lEO0Nd1ie+IRq4inA25h2waBu1Rz7YBPsIy74EaSJP1qSXXRQsQ/uNXlIG
RcK1chqd2Vp17ojZqaCgNREChBKkRZNkmyUbPP4u90CRrbxvX/hT12puKit4yOJy
697lhxX8OqRExQSEUjAwTOwbJ33mOEuDmDB8Jp6j+pXv6jPIwEhxxGTM/E16eX7Q
Oad1GjoW2WFu3XXvzptXskk4iicjf1J2TxmYQtSlSt6oCBnbjzlHOlDGgJpDz1oQ
8Wq2Eni3EFuORAFhif5zsZGfqc8JEuuSF+xOcjYslAQqzQRLvNYqk6KwmRrZgan1
4hRbE2tJ5hFW3wru8yxnK9tTQttdkiNbTPQO4wOBig11Mqbt/62M2WTenUjfhB0D
02oGuqyM74FIzsh+RC2mzNzGkFNloVuedsjglUO+/AFi+tsqLnIEh8rnkT5kDfap
adFZUks+KdTvL19leWPkcN0f9lLT+TkwCh5ngiiLrMffVTe2UxHiY3OlE9jvAq3A
J+6mzwlC1DSDNNPaNxh051Hx+TBCNnAH88EUMt2WGaiL01Sa/CXvViT4UrWsMg8y
yVpk8QO0cn7WxuETLIy/4fzB7WSa6WLvQmXB70F0GnmXp1XT+wO2RTqnXj+t0o97
zSl9jtrisvpSgbOj5FFpFHZ5nnpNTR6QIZ4Koc2WIIXbPBADcJXPPGzdNRXqXUhb
qtDiwHxtgH6/F8xd7O5smC2y7QsVKUO59XT6Gbob4e8qItQCrCg5qFqft7jfQ/AN
sOq2RN3jQn9nZAjLd+oOr2IsDt7IgJQN4ysAgljItYoH9MXYw9W/YZ1md94fCZVs
SFz51wGeVZx5E2C0vS4GtBNmTSr1qwcZpRbJ6QON5JDAX1zNFw6RnrM0mTqxPsaq
iCM2vwBsmnGYV3TfRGzW9G8iSB5GY5zMQo6LBwRV84XWn0ftgW3JCoAgLe2ppz/z
6YzB5qahRskWQ0iZDR7iTfoZaW6PhZ8LWp6ejQ1bjT/rkGYYLVrZ+Qhrnkajk/TH
qPxpWmmK4/6cCoeXNoDSQ/Xp0NFc7/HRVHTmsAAyDIYC6qzMr1QMLM8kxA8zJCIl
LvVh71dNOCJiYFdcpTZmiQa+0v5q2PCDhCXtEw5XzIDeW9Qh4c27S4vxTV9wGhpJ
zs3lt4Fz4w2Tb73tyqqfiuLTSJg/DHwmynwcN/+lQG4AN6YkN8Ky1bDwZe0tDFLY
dM0RL428CXzOOkGQVH3KFeA21i/H0D0QXzwKBc/rUCaMTCFY7hfbt7jAG7+/hLW/
kmKI6jZPOxR17vOtQJ/uLAX1R+uCAgDcJOzwqAQNS9dKkJwy1hiY+zIc64B5vtQC
rsk5tI5HqCZzO0PtO9a5TScDE0GZo92WB4q7r5NyoHmm4DWaH7tM7ZulVbKomDo0
gEvruGLsSx9GO16majyPGt9fgwsjQuq17Imw7yS1YUUtmWrwC4WYHbU3YsWawNip
zhw/Rxq9Z5t9nDJteP/en3PH3bvvXA9fRZKiP9G6Rmspll/jXVuVj/vudD1Dgd1G
lCnLrwBxIBu4JemsNWvR4qjsTsNqLblj7wqV1knuSS5ctTsRGCROK9iXgdsu/Oe9
h3MVu/xU+KCBMRCT9gkaAKB1H+5EO23WBeVUwfo6YDiu2a8sLkTJRnfEOvoV1mp6
G6QKGumzBgUswP++HYYs78c+ZwBgveaVJHP+NqKYTubC6M7hTnmlBp33kUPNDxfD
tBCvqYH46lcsDEKd8lfei1XaAbc2AQCNUxGAbae2lLnnaTIBIyOhTbtdBAXYTnrl
sRH7jO5o9Vt5WvNNxTm0Y6k4ul5zKYDOs57Eb5W28UxrNQzC/KKU9GqzqMnXwDkJ
BQleisv0Nrdk92wzfdiaemQMbd4NIgrW5ajVlCli6VwzqaCeFZaJOmLE/GItmmws
3nb1NJNyYL9jqYwJnr1xctS2LNmEod4Ph9cF207xVCagIiQdS93vEDFayFY+tdDj
Z6ke+Stp9iWmHA6aSAEDctb8QLmTCfvncEkNoXYchThkgyj0+poDCNLRgzQz6YFe
PsVKdq8jq7QULqFa+HpE/Je14b7YJclF2mfhZB2GuHUPjWXzbN6EoImM2GT1RZHV
RI5AzcIJLjDOMLTrUvKCUZXvaQmcdeRey9b71ZHjOWHGlLpXxvmxymGWhMWov0Jc
V3hQ+5mH80JlsAgY2fmwp5v877lf07KellnFbu/Fz2xy+ISFC/EPEENCW0Dsk0yb
vgMysxutrN1nXRIpmJryh/ssoEYkyY4ptS7+yZfMS0NMYbq0ToFigRBOxF4OdrmC
YfY+pcwuEV5IGAYeZ3Lj1oV53N3JGvR9H2ROAnvXjNop0bn8rFU7rxgYPQG6Xwfi
RL4lM3NGkkc6i23VETF20dDKJIUUcfnyb8ohX6MP27ciK+ejKmb9Ea6iHKseFHR3
kfi7JoSjEasIHJZBP/aVujV1bG3V940xVFA93aYf3f7PfETSw1FW428nAUrErzch
T7dS9efD5HabZ19B3G1+8Gr+9YOYd3nqGcfFBxy8kTZXKYnorj8nFSlYFs0rbl8d
qbInq9x1ElZ1FazHvmPgGSIJtNUdMud/6hR23OjIMECcvx2U4fT1Wd5mHJOHmwPl
Em1myyh33hFpHD3OCqTb7LLmL01SMGHodAjbjtisZgWFB/U1Br8zeCJj9VVwnlg+
fBI+X9d8pOLwXDMJ7cZvKo3t7WK0Y+8VBxjRW4v3W+LlbkriO2hZMw2Jl+A/Auyc
gCa0arD8gi0XKPPqFFYg0J1rXapL/UxNwGhO4ElbCKLdMTap9ChrUHdlWxwlf83D
Wu6dUdFKrr0ZYd3E5gCQM/At+MHAYZ+7znMD1bT3noiV0do3RtDaqr8N8uVjtfJY
XBmd5MWe1Wpnra5sjS28f68vVRocFWVAJfxeCfoqflV6I7zBPU7ehOUWJL1bzIWu
AboEQvPokE/izCxAEbI9rfFj7YsREZ67TofeHkmiWhmJpem7hHAyuk/pCXd6jMUZ
iPyojyg0CiHAQ0blxnVo5TrNsXng2IErXpRwLZEQke6XPR5GBgZpyAVd67aihi98
W/lv82KhVoRc9rlk6KPXPBcYEQUXSzvCRb2aC8j+dJSEm3dstXfSM1kxLlS2iluh
jivPfC1GpLe2+9ZWiLxTWlrVR4d8VKU/8ifPZbOhnIiAmJSiYR1OngEgyTcl0eL0
P4/YrQOrVRwY67QrFL6t+t11EWFGD/31zEo9mPzKJ0HuM58cjR1tmOiPGyq94MAd
6CwL6Jt4PCzPUclz923CpMQYji/ApACbpbEGOdkZVUt+f+9MIWFv8dQktCgmIIBT
k3IcB2TES9SBxxXzbVfSd/ielFCKe8sEa6ZP2NHC3CwaSjJoEWl+mOevr7WoeK5h
FKuGyBFy+etaUNJSuHtC3vpdH6usBI9n2n64oJTaVx5+0KrQr9oo2HYdSRyj218s
HoaPwCS7V6FBlCoUzyIT3ugtHA7zr8AtMDcKhuJ/o7kcGsV459VztSuG7doFKs2D
TIsn9vWwZ9xgFVSVpXn+O2qP76G34IankboHq5d6l22Iwfi3AeVwaHew+CPFenqf
CNMgfc/btStp6Og4uzi59seyoIb9niIZ/adl+Jw8oSn2qYOBSS3nRYYlwZ9EXqBa
TBxoygpCYcc1HIe8E0Zazk5cVOETpx4iRpsV90lnSbRvxdFb4v/YpIApg6YdtKTH
vD1svqmC1yFQVflw2RkSck/dWL5L2DPrKIC+ofWLvl3VEiPU0D0Tgg1vcHqfzOYT
302JzF9qUFiDNxdnjjTs2Ge5REGA9k9U8Z/EfnTQg8YzT07bYNzS1DsF+xI3MG/A
kZEYjNfUI9pyDgNkWwVz4ArxHttNGU+msl1MU8tZ3jpiQoZB+gKSUppQy5TI3Cxb
ts5UtmGMcl6k+hK2He85m2NujhYs4F2+DrY1jvBhxeKT2oWYCbXVVF7W+N/cPgVi
EgVlqRDm+sAbfPzxgHwKnoBW4W9y9FZFhazoiU7hWAuOMQ67WdbYQY/3blbipNXJ
9cysDNPK1qQedgU/9Sgrfmqvf/AE4xJXGrIlZBE0t8HG8Bruyc9Gc117FSBW9Lsy
Aw13XsD2Bb/6DWCYThOl/uXzmJ2PT0bv/VU7Ec7GPzH+hYav5FW12bKMeaONg6Rc
QcuVDUMtx9gmPiuGHnWlmt2ZNsbOh6+VjKOdwRfbBDPJkjtnuwDmi4CCfSEEzW4Y
tvpW+09jEV7L0i8f9/Ea89rFBnFW+mNWjHJsT78hbXzfDw93goZcbYLK4k4IOxM0
6cbOcVDC3mYLmAQPM5o6WWMWh2/aYZn59Ca9CJU7OwPPIS5imtONjxkdgyKX7Gq1
6v6g5j4WdkZYUwuv+XU+PQvZ/glySDn+KJdebJalgnrRybBrXG6efjSGw80NfKnf
8PriNdWXUoxzULLO4aLRCu9H3CN7s1R86onXCf2dFAL1P5EJ0LhpvPxIO3MZkHys
sv2I8jFoVAHiBbaZ1MSBPpD5W39igXcAbeY1iM9S9hJ7zIbE7SlolusJySpEVOoF
8hPkbqSTe44f4hBVNBGPV9vnnjgMcbaMCwTyvUL1aHkZKnDkXJer1eC7Jzx2iuhV
KgGjdNrU30j3ALOMJ398gXqc4E9eogK83pNWnvwdhplSAvnDAutXA7sWOUyZu4zt
Crrg21wyNWaPeM1sD/2jgstJOGuitpjOtBXZQu1XOhblLHtYrRex1N/UL/7x0KSe
uz96cWmTEQaTHhqnTfXI60MuajUqExNBggBISKnT5q8T2fKjrMcklMocT3tYX8K8
xoxaP4dmcNXHtfIxlXrOECDMRkBCyy/ZAvmsdqR5D5rHm5d599fSuQrKDjaUvhV8
VoPhva9YHWWyKCOL9Y7ANGqt9vTaNL5Uxh+rdzuUz/MHwNFnnqPLswhGUU+rHANc
yJVOaXK8IJuc9kx8XexSDVGHKqKzJj8W7Y/7Z3Gx4PqjbLbJooW9Ds2Bq9C5jbJ8
Q5Ryu2jVPRdBMRYb8C7x7XLvakaAr5eoHfXxM+Osoik3ejUYY53qS0i2Z9rhnBTW
kxSp2JUvM1wKEKND92vY9z27igrwo83a8JCKyBhHhSUioeHoiRIWLPU4hjuR81XQ
vGdCa5URVKhcBzt8XhfRRz0FEc0K5YjQlPAtKPMQqAwVml8zlFmf2gEazE0AffXh
hd/fsYRizrM2Pq+KSnlFWHS/RG6asxTGauJSA0iBqvanVgDOn8k341UIAIRYELOd
Qr4WBK+tbFuE+cGwfTpiCTxF5779m5Yx7LRUBbiEX8YT9AI7WjYzwcIXc/GNxCEi
Hby5CMIfQ8p/7a8aLwMUT35JIGYZxdYvLT6fVCnpXHLEQdfcg7YyiUAIo3ErbMzm
HhyWQe0/3vEPK8O0XiKzMjuR3XFdRFxLjv3xsqAVRzukCDae26X4SNmQ8Eyos+Fu
EhW05NJPPnDHrVFiMaCfNae9dNINInEshuj4fr/ELLiBf1I+b08vSx7G7pwGqgIo
Dv7lhQcWXTM/TfdxA4w1mTSWh8iCkPTqHtHm5xC8qqhwN7RsWcIbwVneEK4kpAt/
KUq5bq46j17LspSE9A36oEKw+Wj+sf+H339rKLdpAYx6xOJbrmwg1zBQls2NhuIR
nJh/dcgVBV6LcYAVduw1z6tls7G9FASv4X2md2aOjTOgWFWrA8Ov2ryzbUQ8Vqlf
eOU/H5X2ZekBd2FRjbCi6hYIXtT+ctaOE4p0EKC/KlFf3Nin5BK2rqV0v+XUcMqO
bsq6k44A0NgvCRJ4KP7UvETrFQVvc9kdWxa9NwSmp2uh9MqNnt0p3cSKFHbaNZAT
HWIrNfxA/dGcAcvAkEX55Hp+mdPxTeJTwOx90I04DC3mg0hNPJmSnqRP+uDUytDM
XOh5ol3M3xSZVQjI+bvXsoLwgXGusfa/Gg1YJNCWBIAqbJD7wgaT4eQ+8hkdtDtw
lcyoQJOPnqQpzJyPL6PIaPQXLLdMlUG/wcVMbBCjkDgD67ELsJ9CPem0ADOaElm+
lmu54vSNVR3RGIDEcwJsVKSiY41rwvjKU7vmSlEzHSGdkL345pr+PDZQLB6ux/CE
p6tUr0pDeTasBczbp0VK+lRYapOvqDjnovA2G3jiDDEhUx3qbpGnOGMVAHpqCgek
Dv8y7b1LOOXYQDHNJu1Dml+Tn3BtYYvcDgr7Q1SrzIAVp/NyIM1+woEO0Z+7iSHJ
uDaY24Jk84AyAikFi5rKnM5Ewr9A8AXdztAAJOKBnNwtiBLYsshvCLZ5QOhlrC9w
N+b4B8R4JuBTuG7SVzyTY+iY0HrC4jrgNyRJcUCdvdOoQu/0Ciuhna3m7y8mBhTm
M1AahH3l90AXBfKtH3523u3uXDdT1L6yr4lbMVDbuVVemmRUp+WpHrTP5fEEMYHh
2HE4IIwhlhi9v835Yw4oGrj1TSaTtpV6bxlAFINesqsHj7NDEfiItc8+LG8lwgRJ
ezqJY3+HHstl/ANMAGToebDXpl4u4NFEaahn4Q97bgRANMfx5t9lqZD1fH4oLes3
nia8mjG0qyJen0Pije0/WWeH1V4HoORGbuxeijmQHNu9fpZgKqZXoZw4Xs/dkND1
9+5cvd1j6QTFsOY5y8SYtO/1nCihoFjnQvRDu1vi4HY0r2t7uXh5dXSr3vOoDHgB
2hv8ASYV2pxz1fX++qf7Am63cibfB90W1yaG/d1h73rvFGNNuheP5ccV/yzz0bF+
WdzE+EJ8662e7KJRGm/ilgWf3qvNQITLhqzmNrlknTaBSaS+88TNZUshBeI4/v/R
3KPmVjnEYAidw27JqgGObW9pngqhnabz4cip0k9jte9PmHm5htwgWsyIcIKs0OIT
Al7NdK/5T/+CywGU0kkZAcnTIk+l4pfFHd2x8jAWv4DCZZSqaHwlwvUkXg4/qx9c
8xrqKRd5Nax1AssN70/vPty4rqTTfG6LeyGQy16Y4/eyZa7Cng6Y56/SF5Zb2IV6
DurJLTktArbGp6V2MCf3bDc9o26mOLhjnmk3AxHKG3RqkDmjx06FrOsOSG7XiY7p
QUwkCRFK2RRA4q/BszbdCHANw72XGKDJq/w+DYlnWTC6tuOfnp3rV6rEC4O76aG1
FM+9UysdTQOvWob7UPkdJfy0nX6IF96sntqLnkjvcRWvd0ot1D4TW45LTYeajePA
TXvhCBvy5iLTq68XUp+s+JcVRSHL7frWHTLtLfHJIhIIp7Ecbj6q7oJdaalDnnPv
JuvBpy837WuQ4og+1Y63rx5SfSiJewC3yI7PxYrjXiEYq9N2pU6IPAIm3t2ISg4D
uB72pLNjgxT+uVPadooeyrHa+/T4TNXlq06yoebEIcjxT7JsKyJBEnq/4y8sT9tR
qBC3PwVIur4ZS8KmTpK7Z5V/wHrK2hbRNrUvwq74qZVPNCmVE97NBBqT0JCtV/oc
aIWy/yyxuI3KOc6tYyO4KlsPxPHQ0IPNPV3f3pAkW2oKAPSvnZgGoA1SKascYuNV
d4psSwG7UAi0MUxk4Cb7H0BeU2OjmS+1t+2jBtkMGANktwbNfSlY/iTqlu0sOiyz
fN6BVZyoaWQqa39aH6qg91YRmZ2wK7SYut9zlNSp70xH9PPMgnHCHdWXpWh4lL4F
v9nJ7wvM62XWS7zskAe06yuBrYbahIogFdonXLsN51rWpIU98MhdZlI2aJidtQVj
v/S+k8/kHba6MSPyIdMI0e3BDlC/pDFYsNKDtwMvh1/qvmDmwONRcz3VQBgstL5R
/ioh1lzVNrXjzXh3nSN5iAetEzDQJLNhp9K3HGzJ3TAq6LaxHZgAo9mQLty86YuO
dqBvM7N52LT0chqofUenja1DA4dGIEJu/AHiQao2hTV5MHdPmD4BNE48mTUzcAig
kkTIA/dHIXp5auHbHsW3vx9aQjRFi0Q6i5LqJq4RXlvKxoADuqSAPT3t2PPgEHH2
Fn42f63ifAtPJM+kRduuNOhJ96UInUQTIogD1OLm5KEgNWNNz8PsscemaH3zBePX
CFpNyiqoRCWA/5KOQW16Nf8Qx7TVZmyueeV6IeMRMdubTqU3LmPTlIQ+QEqKQrgp
XIFXxIYNc34mCXQL5WJtu6N9JcLtMjLH86k1HRqTeY/LItHCVObJwMoSMEXt4uk+
EgHmndt/xr2e7Ke+p+iDVrnaRiwglOxYPj/K1no99mXAvbmnl8ntF1ZdlhvcVe31
AJf1y1Op5+Jpq57lC+exW7ffsQgPDVsbUfm9vSfQxhe88mb6CSEQZGfzLRg7OW+N
5gJJypNY4n6687sskJcbgHyFSLBmmguMNOffmoCmJcRfjrjXbi9nWVFj8KxMCD/P
rCDM8gbQVJTCTVmiHdnQBlvU0TH018obm276xw7qQ3ygh+YjxTUo7ZO3quNAcl6t
1WW6mpCMvvVceRpVuyRCa5tqghe6q4ETIslp/BpgLOQvcJATotjKAYmjMSsKt3Pa
fl2mYg5Hu7PyGDphyrS+jlWZv+mBWhR60tb0R6out8ztH7EG9triDc+2eh6zp/iS
FQ5mmK4PH3SRHaSRtmsf8J1aClamcVFADGomygTwRzTQVKfAnJLHerLRYO2rnw5S
WP0JrgEsNY1gDefYzMMXZHLDn4wDDtu1sioBReqQicCQLA/vkFpALScEof0CMpyc
HjJWMeEDJPRGPij+OgsLezIZIllNhCMueSrDd6ECwoC2um+fVeuz4DmGomuGfGPj
xGguWaFLz7ahHr+UjJbZAHe1qZMk0l96zBc6e9ouFaOHJlLJtpxP61DF0lX1sYPv
hUQLW6IEkgZYtSqSksUQ6UWZNw4J+AFeeaMkjTxoy3HRdkWpKq93wYH82yZZV8pa
MxvQ8ujXDWbRfV5RHDb+xKwQrVGug7fY0t0DVcI+Ng5GSsCAqtSSfJ6hqlVhAB0T
FUqp51OQNXrIJBRT6Tw63e3L6e5umkolq8bzGKami3Rw2WRXSLiY3RvnkwOMjqHQ
1sC6HxVr878sL7UbLMuv03kLQbbfMIBSBLD1mJYxAY7/kCDYIGCk8RSWU87OUU3+
ngPrcFtAQV2+u9PQ5LdsNHKy6xYOXP5/6iCGjGjwvecmehEWvjx+cl+CtJF18eRq
j80+68M5CuwAOf2rFaevLoK95D5AMQnRsoqBZRSyg1ICdjYiTQCs0CRptvkCS0oa
Bf2/55S445HcIzZNeyOqYBzh06l4tnhvoYowI74vKiRmKi0aXgZxvRXylRlTSEF1
1jRx5Sgr4U9dXh5NriyrDtv3hPet8mH0qhqKh1zr4XC+ce1qes+LTXTdQ/MBTKVI
7gkjQJSbRM0YVxYumC1hpknUfNdxT0NNVMjQmzm8ZrlpbHpXkDuvErfe+p4UdNo1
gmxrTWfxstltdwUH2wsLqWDg2RTNe4miQtURBpfDWvO/0a/mIT398zVP+3hqqH5K
1zP6r+5yohe8pNoGKG9xXD6wk0MpqbTjYnv6er3dvrN7E+Ej3IixlbsO9QlLXoiX
z+qlshkT431NNgTEJ/Ov0Nq5xAWR9bKVdX6cExcsT8DuAJ3TDaQAx0Y8CRwuW4v8
3fHlpOB/D5qpNi54mx001He+brAE0ZNkBmFEWe5XcijKI2t1+D9SX8AVwyv17uyA
QkGRWJv/yqy/r2y3t712md3Th52nKaSYXABssRtCmNrfAnWbHUF40Zyjr5rYcdyJ
/uXeXQyfVn9k1yYIeRkoSYwvK8TAK4rlwqizeJ17t1OqYJ1v/jHPkJ5ip5UIINZ1
45vz6y2V1FPzfnwb0d2RhoOJs/kMx7mpE8j59vN70ZrvXnDg1mAm4dmucZ20UG8A
Grw53gHgEPLa7L1cQP+piRwzy1XzqE/+sv3ByjIm2kuh5vJ05qgXTGrngTDSZ9n+
+tBBL4H4XyVCb+9Ffi3ZXQ6aNjsEpxkluJ22YaRxirprOVgKoAIoy6tKQmzxa7wb
60tK4McqAHXayuJ3aHRnYttF1EeqGFU8RLkJP9WLRIhJsODURJyHKxP0ykSWiMF0
thzgBYHmFJsRxSNYB1QyfUvYtFXPd1qZTID0CExfj93Mb0/na1pDzPOzAvDxyy/b
aqwtzV9S4sO5mJO8LIORamfJh29PjEXudvFajdUMacIVl5rYpsTGMsC9EfCSFA2W
nK9T5Fsukxi+GEd4UqNz402lvtMbZpI9RTVzvaoUAWCUwWVn/e+h+O2LbakptK/U
OwPmwWql9JI8AIkEl68CbzLzHKzNejf27+qBwn9WVUY/mujLdMZyNB+IbU09fqx3
j02ZIvI+IWockuV6OAcj1snMDpDpUxQBoEKT2jI9NUYwbhswSOeM2G0rlM4uI9j7
uinkyYdOA7PImoCYfnblsWJw18D/cDo9qI9XAB9Hja7FlGO20SnIYkgnLIizs3bP
KgNWiMm8ApQteSuBNXR5HtJJEoZpmYpA3hdbS0as1rptbqGRhNPPfIQnnBVe7d4z
u8UJq8EbfB3TEkSKNKDWbF7em1hYTmTnIooC5JxdX7EFrXsvyKhYVWHeE766WAUY
qYNQ81Za3ckEGS8Ib1Ok1TVHu0tivPwqogKyquKJbvpPsBv1T6nFH53h+FppBOls
tcuW2VjOUjT3P7fS2+O8X2I3ZtFSwQw/fH88coA6S76RlLY2VQgBLWlvIwv4YXRt
lK/dmt/18z5GJCgHX+HfLFQ1yf0dQIWEry7LPwo4oz6/QcvhIZt3cmjmPkPo/k/2
nPY0Z7uqH8aNiS4Og47VnIbl5YtcEUH9nyWd//wgDHr9JPJRWN+Fg0UFtiZctYIo
lACJyjyhjKgTvHTdsAWFoVqGt9CWtb+yPG1MbOT3yvuhFSJ76yXySb/JeH1zk0nz
U3q9+bBSKhkpRxnLVI/eBNR4SqFsmf/xWMFEGy2DZ21We2h6uaEx/ni9TUQquosL
XoGxxENpNYdHdEyJA4L0eS2y43ZCSak0f8MrdwVfhz4vQ+UgiFXC9oIBmWDIVcep
pyMja9kx6MgcXTtKYrN37t8ADUW+FvGHcrSUDTQ3Nd+EITV5yOC/uwS8ju2kaidZ
/USkE0XFiNAhoRLR6ooi/R7WMoauqkJUZlCImjBSy38NlMuqF8uKmgKN14IHwFuH
9tENka1kudXmJBnr552huT6+YBO7ATJgl2xelHgKwVbNhpbRVq8JiWYcO4vd3aMX
+9DbW7GRPnjnsQ0UfSTMt+spxR9Mm4qJUmIFatnOe5OApLTuofndSLmfA0v5Q5fc
pP/EDuGunl0vO/ABdA5qs15tijF2O/ptdet3C6X+eGS0EsiIcewRqfd8Ll6IRE+K
O+jwcaL/TuXLTC5EZuS2DPI7cpSWNwiq76SgG30JeTf2Po1zCoTVWPS+bvN3Yrm7
HTiKe0D0KozVCsEwwnG0vME+8BOzRcZz+nBMBCHv63ds3W/Ed7Qy53iwE7r75F22
4WnZzOAjvl6cAj5lSL5ZFlvTPPo20KX7yJGBDWktcSCAjt3KBvX+/DYJfrY3n3mh
m32k0a6Cu/DmdIYANVlNPFJCOIrGOBhgPnoED20mFZXv0PpUp+dFtjj9OecZz2QI
b3KyLL/fUS0ORXqPw3WOhtwEETStx0suHinzSM0cL/A3k4cKItS1FJSvgTBlPaof
w5R2OsuBw0LjfMJ9znL8Gpq8hNTgiGZH8TTSfEsD/4nWrmW3CuCXo/pOHyiQQA0A
jICG2p+9cI3AWWEC6JQ2pi9qw+e9DWaSOAgtq4sSOxkOhUp7mn9v24IkcUBVetZW
DQ0N5ofcSSg8or+v5aOZV+v7/9hpxpBW3v/weFvfdVAC2geCXnd1ODrvOTLuOB2v
sENviJHG9eNo/uHSZPHcyzwwx+/PT4xzW5qzRTCZAY3TRhDQn5nnUz7RNA/VC2HU
LNsseCnDLXoNO8iSBM9nbpB79hfEhHkYwHo4I/W9j52/xJuC8JuBuIL872mhQpSa
yB+Kc8rqGhIHEXR04ISsq/iXec7AUTTmgGcofkB4EcJo/I0ETLmPCxCmGoiv42pv
o5QENblT2KG1DHLnmBgLP1W0ON+jYOf0kPTb20uMQXzced767uPEvaB2cb4KzfP2
xBcVXEDbCB7lNOJPQcvtuyWWCBP4TrMWnQNFcHzTLcjy6F66pNLbKcrsudWNqx5C
Sa9VM5Pd9DEpaxXesM+FnnuhDo7130cOdG5rJPhNy0zjyGcCFCzdvtMJVYX0wCdn
GhN3RheqNkG4J3/Ph9cvxlVAbao0hQ9G22jf8CLq2forQD0bQRMeEqqD0lGleVTN
8KW8ol/eKgqY8M4kZOzOw3vo8PL1FUJerEuFQG/yp8DfvNZGlqByx8hqcRQsIQ02
OPifrleouWinhKE+d54HkxAWO5/F2mZ663+Uum4Ge5KGwe3p3VPz2TaqBmMjUjyR
D7+SS51J6vjhrSGyNd7afTH6744/u7xNRbWKM7YtbouNB2r8/Fnz9cQcYPd4SR8K
/bmmeuGnztHtIvY1nPhS1UbSYOvWr9G+BbctRDqvCpyuTY4sn4unTx6del46Jem9
U8Y6RcUnkBeM076q2/oZSrHcmtjjOBUNTDuJ8oBI4ettdJsvBnSGADiI1C7kzFru
vw9jKxHR6ri4v1EiiVB4TCemCebfuTcS5h7StP4kwmj87HeZcZvZp4jUUxJ3NMJI
ErRPG+Ou5GfOiaDeh0lXIRywR98AHFuizpOAB7UzU+/IRHqOgMAg77jVoRyoLaeT
k3fV72WL2wgbTOyYtQMKHK/iqTebQRfjvB1J8jHa8Ly0LQBIXMl4bces7FnouXsr
50M7t7anv0PfgVY9xhWd4aAMxtpCzE/6zqsaVAo87eppLYB44KyAQBFZHzOnwS18
z9TZu6eUzbp9Qs/PsW4UZ38Tzi6xOlyFPhP9lJWBMHxSZijFSuv6yBLLXdraapbk
SXemEJFO/88WOtFGkC8TkmtaNcIXWGygkmulhdcu+c0NqaRtsBawPdAEkzP+HeGL
krAUsejdP4/n+rwhL6WmRDK04BT2tDJmjj+UIt9J3byjCIA+tdLXT4WabQ7S1YRx
qbg/Dv0OaVWp8P9NKc4Sq1ZQyyiacYzvXniwq0DBlGhURBxtwDNpBHw1fTxyi7lI
ERlQV9jBq+ZRpu0AzUDIs7xpHuE5Akff2Gtbn6R/CgAgttlXwldhgyaC8MldzTkQ
oGIhll14MnFXhfAdUs+cFKV+JDiXRAJXaIAdYLU9ypMbR5cIWASrTLO6wz7ZrjFH
OiXuUd+xqGvx9wuBzuE0CSGxX60BUSgKba0J25/XRb2jbiwdmZAcmFbnAtv0UGUc
MtrGBDCFYwVxkCDB4BgTT3ZJxlu+1rY+4p1d2QgHQ9Walrzcn5DdTkPWxSn2nY8C
/PTL/ZkJY4YwXPUBt+xzKsqDiIUU5jPAR888zIf/HwTx5ijg9dmzk1B5/FVX0KUK
gNto3E45X1HfU/wJ2FqUPwjlSWb2DDvNt7UMe15bat/BD3LDWaC0/QrH2fCkLrGB
PwAFrYvQkvSVeS7U9HDqjrmimjY7+41BzxtimZCeNIfikJ/UDcKhz91DIg31Cpnh
+0yZSczAKDbujSs7XI1T+7/BFZdCwKvOTR4CX26Oo8Ucdgnx8u//nU4SW3VmVIyL
qqx3ZTZG5TzqMI4EOHBak5yzkWkMEil9zjIx+RQKGNKXYbXQw28JGZ1woxTsUkXk
hq/1sOH27zxbE8pGwAiYZEQfeD0Nlj/pCkDdXeHtN+uxh1IHwL8E/REaKwn2Tzjp
87eN+SRnpNReKDZIEt79EXlVRrNIkGBQ4/jGt15kBbxb2b6nn0bHhm4Vxw54Sce9
HNvQwyKRika8lyWjKsrxOFH6/lIP2oZq6TaTNPcgghW5v7z1ei7oitotJn4ODEkA
DYx8vdOviNRNxcA+SBa8CEkwF1kWFMDr7iCuZYgM5cGnSDdONNFEjAwZbuEEBcWd
j93HA7n8I5xNTkuFeohrtuF6yrR+T/CK8eWqqRs7t5wIhYTxY53kxDJ184gt4KYw
EKAdjZdsa30AyD/Sdf/OGVdp3cox0WBi2sRC6vt0dt+0zR7tEJ36A0gz/uGAckFy
zToUdX7nq6H95KSHfc/GvOwAPLcor4wZytcH77zv0dyApE4y735HzlKmVvGtr0F+
3415H541Fuj6qevF30S7k1RMb10H3xxC0bnCf8ImU2TkuYfv6QeHsX9nLF/8jV4E
XiA5VRwwWVNGfjqZW3AFyDKfSuX4IsjsntMcF0cPhYZMmHjQOlJgnlp/QK6jXG5m
Dub161ZuoXhPdziZIIeSLlnJcLZh5avQa64ekkwClw1wxg6UkVxvfbLggu2EXXwr
gfQJPohYsLNNCdiGkt7Ddn1Wib9co0mEDb/a3fa6poRiGOc/n5oixaCHWgoJxaXb
/zkkWvLCSzdfqnOCTdz8fOiP5bM37kA/wOkpwRq4u1l5w9DJ51eGmp3uf2o+/m5D
zlk3N3J2XWcJfOgl94gTZ6dMONG6syKSLNm9xhqgduuC9CFjglSTxJO11bJneY/l
pbycQ+6Uxmdg775XxCkKjz2gFEMCh2CK1EtAtKNct6L+b9m7cvk4+6VcuLTxpOhR
dFiJ6iCVepzIiCmU5QtyEbiTj4wANF6pIcOCRQeWTPgRyaHEQOl0SEb3OBNfHz6D
LfnIYfc5HoyMyvSctCUHdXRqyHJhaWxuRwznB6puLNaqJ7YJ0e7psKHPuDR97ANV
GyEvj6lrfRlWtWOsmO3jXCwJDQNDZ/7XRSGSHEaE6X/Iw9MAOE6+mfDuvl1LXdf7
RgNRVI8V9bbFagpA2/d6RzgumUHgvQ48uQpOOQZ3qJaqpYxxk6MWCKZc00mI3dSZ
9XQoQ2AOqy7kRlIb/HV8MrAHvPHsidWFmKQwAoAIet3KOv0UeM0htnai/Eq77sZ5
9ijaliheojLsnTRiJRu69BSJ4+rW+SEqcZfMliEQzIK/vD5S5vyCK/wqSy3OOOnY
Ttq4vZm2sNa0Mzx5YzYW0ueD2qMmoMO3xYPAFN3uduBe/GBIyF95ZKstR3Tw8iEq
zGVaA36klKpTCRfidE0KDA7HM/bYpiOxNSTd9k7UK6CRUx8XNMXWGoS7dKyPiz1g
12h1hi8YUtoutlxHpINnsSZ4ySX/3pYg0cKbPt0h7VEtq6bwsz8N8qtOcJtc/7p4
5rHJoEgir50cdb1k+ExdBFUxiBdBE3W+I7H0p0OMHm0s08EGGuj9kh59cDwQghMR
f4QKDR0WY+GFzgrN+OTfW5tMzHkEVixVATyBiRKSTzswcX4k/8MHlCYEQNQC+u1M
5Q63vwSxCvU8+MSP/uksKk1HWKlafqBx2kuO8kgojQ90mR2y5KNgcfSvkyrDihZv
UdszLzn1Q/gKMfLenHUmz/qUj/ycwnemiePRCKvQVp5JV9FsjTgLZZjR34jR/QT3
Q+xynP/EbVxPc/0Ey9RXhuMKi3Cz5jkXEewpJXz76gtPqER7oGwRIYgEezrTODrQ
mIt6U6D0pH59Vmwgl/SrxYIP/oCxLWrgbAZQVxtKusbimCYAzZPGadVphhtkPp+f
Y86NPEUiNh+5iMpdVtmrJUyH60sbJdrZ2NByIgymYVS96RQGS/0WY4KpBmLl7vEU
a2poFjkF9g9Aw3iMThgedZV0VHjYFXZmilDM8b3I5KpFwbJCoToDlgr6/8sEw+1X
4szuHCBlpjYEzJM0PdKPgRxC0rNVOmPuH6onx0LIfnutp/VR6iypCRy241JKAaXT
8/qLXh7JOslK2niH5wQkDcFMVzMbmZ+xGnLG92myhlu3RPjC8554WyHKMq7i6T2d
cpsui8TbAV+0bCSFbgoGzw7lywzXxSoHJX79N1p9aZprUILiZ1XeAk3f0mo26VYP
iZ6uP3pCW26met35J95gIg/Ce1SXymYj47ZUjHdrC4GqNNMaUgis35kG3tZLFurO
7cZrPO6Cd9Kc1sGSWoH2slQfNHbI1rTHCHOlQzkAMbfMCZmInCHIrSWsGst/8j3e
Du+iZ5ReMBAUoelJd7la/Z2LgfRM+0XX/NsYfyaQ2lrhLaZ5RQirAdRO+xJihVJP
PDZ9d1Pd8Ta2q16eVd6Fh5Y6b2PBneacYlsqGrtwESzJOXzJRVuHiLnzhQbDugwj
PAb7ssjJXUb78StB72ugFcG/Ea0REJa7dyeGh2L8u7xQUXax6Ejk78e61HDqKwl2
nFzukLZkyIs+njvsL5D6ZiYIK2txhrla9Gg6DhimXva0+FTiZYHEYkn1J61ns/xl
l1ZOFnYAe808s0CF638J1Q5uGgKiL9aKxH/iKVecmgR1iRogYqQpPzomUd6WaveX
e/z+Ce+1FKcUZPSRCFBKYukMDpWz83ohcYMt68gSx+XrkPlekDwIcnCIhKZYuz+a
KmWY81dI+ksFsFRMysW9ZeH89sBl13JHKTD2Iu1WP0kRygEDq0Novx4ibPvCnFuX
E95hKRhH08ePlRHecTAUxBh82Ypks/JugUmOUd8MXlrSETC5mI5K2i68NKU7tk4y
6rJZfKhVs/VS7yJXtv43qAn4OY0BYbyqq97OxS+GzKsOPHAdAcZAV7YhPMhRDgHU
LaJEsHwsaG+d7FoqhiW04jmdvCuPSp1kK7U0HfxAvbalvaUW0bmxg4OiPTcXMswQ
jSDNYD17pZzn4eYC5XhAD5ELi4pHXO4EfanOmPVcNAPuVYac3i/sAxrieFWfOSu6
pGYZ2FgPya27eXHk4dngaNnbYbFOTMfhGJpGdIaCntx3R5hjBhSMHRUbpopG78WD
c/JiBveaXwI1zmlwdVT/IJDHQ9tTuf9UhobPE/6hcoIwI9oDbnHApaB4k/gYCQY8
JxVzC24nJzmeGCpQrYb0d+cuyirhtB/kWdkgPNZi8wRLhtV18iLHecPsS8vBNtCG
yumNkY+NED/7Td5jppDB+pPAqeUKcSpeMoJt+Ia8IjYtcJfV1L3BRjpYnLAv4IO9
cIjdfGRH3Bs8i0/RFvrTKxIG+JvsrmW7J/JGc1PITDFgoKecT87kGhIStbs9Mk5w
+Qoh3ud2uE9eWAk6E6zA7+Z19KQfAvKCA0yJIs/fSMFx+K0+YdnL85otu3zMuoOA
J1xFdRGOctLrHNbrZLg/EuQSw6/M8yvSlq2VwfvZYQOq3kaWGXq8jGrO31vu+NGP
Bbg12lvZaPCTmavhFrrEREVATMXIhfA64HJhjGzNq81x91gZrC3cXGMCLoy+I++w
F7CcieCKNLk2WctrXSBslXfen2qthkIOgoQZoXFy20SvGWvV5nNrALVNZkvFSYfH
D9ECFHMeM6NMAqEifE3HaczLpC9sdwXFcpK/xu1vaJoGy0rQE6SA6WRc00XgvSPF
9ww5/MN9IXGHqMDfY8nG/u7WFyFCVR5fWYEAuUNnv2lkWdFFA3fdQbzaHWWdLXOB
PdDSDuqS2gJ/iKniV2LfnTx8x7BjW8IGvHwoTxNo1xRzIOjdEkusdbYDH8E5X+Kw
QEFe4FbtlETgbnP1MsFBJrumGL2KNLfzCfYXA35Cl8bpOR0gFHLnx5LZUWoy6iaa
v6I8TCF5zv2/hLhhA7Cghj3Xx1ShRCNVgsM/AwoKJZMNLc+bg4s+qhYBqz749o0v
6IjgVGZTF0dXx+oPzpOqSY6eSOzamn8K1IS1eMo/IIEsNeb+4WAHyqEaq4DGGd5P
EAU6s1L736RXIFJF+BapdHJG4MswU4SjW90p42d8sKl4QxL8urCL+hIoUyD6JEfp
X9gVgRrdIR+/TluhcWPE3XBX818vbWCWLY3s9uNoiZeekhmM8kxSwkT5Uivi9Pj8
IMqyOPqWMSVARucSIXtgTiYVgt40dwDdKGNqvNU+QG1MCR/EMn92xBG6Vd+ronYU
WCbdwv4Ovu8dAJHTC37zCdYNdAHuGE5bVhfql8IemsBZugVlmJZVnOEKNq3Vt8d6
cA0HoYNtlt9vBgZJqH/9Myf4MYo1UkotJNqi9jUBPOudWMWLYQxrErk0hZQuavPy
QDhv59CF3J39Kvm0auuNSnF+UDVBEV513r1mxI38RXNc81LWPq+EDmc1OlFbK8Fc
0VpJZzaYQRONTGUCvCWh5tPHpNVVOlOetq9Dz5/tRHp8P+moaHZe+iGS8d6lQlHm
OfWkrhFZZsPHhSahj1PupaCM5oiwOR6UCGe/Tj5EVw2lq0Le6X6oKS3WyquiFQzy
HGzSYjM6LPW1AhxfxFJ7m51+90n8uO+4zr2zMwH5XUn+2q5IFqE+s5N+QPTDmdM7
TfthlWTwMRRXIL8KkNKBQFHzIRecH5ZrMsJshcU6nMtGCgBtyqPjvJfWD2wfdmt4
tYkBOGmt7fdLUivl9F2AdEYwNV9aJurZqevg2eerY3s26SwosexqeD3OFLN0BQoA
bZbSyN63LbF9lWr6xycSGfKuq7bNQtAPnVeJuwkZljWOTqsR8fne9dV2UmA05rgB
eQ0Eb+LGtKZn5hFAmSOW1naDQ6dDwKcmovrheqlMbbXqZ6zE+l9oRHU7SmZcUFuy
UWPD7CrvjxP2PZKf9Ad9NmdEd5wdm0aqbsrLZhWyB5oWldBoI7265YgRROe5xtSy
hWPSYtgS9Y15EYz68F9voEiJpgjXas+mkLWNW6SO0vj5LYaP0qoB+h6aWnNEmWna
xTH3tNfLetffsL33ICG8o46nso9QcmSiwF85eLTyNbr3BUZlYkODwnkIcSpSFH0Y
8Zw8KUA9Vqz3DBoalia01LtYse16fyK+rUg25GZRlDvUJEfsCO6LYrWVMWtrkhxC
LOjBM9y7KFHF7IaDO3TVZ2mSSzhmkXz3MI6+mLHsx5WKhbrCdUCMr9YKIKNhdhL6
tw62qHLrF7egGo+RHG9q10EYliJQCeUrOwxlu6qeBqkeEhyrwRdm36OdFQngXGBA
ynxbe8fzm+chSvK3A+yyrI7ulG1WuE4HdyP+kwcZwbp8wOceEw75XSTE8f9WM/Bs
8sTQBpvP4nJStJw2RFgiVkaNh+yHWG7ikUqgJBv1RjbRf1qCrD0AJZEh1egT73U1
Fui0AWTym0jZqxaWZ1/UvJ4dUX6p0PNidHKv9aNHeGvpN7dd7tuNBruVOYm4do3F
WcuYvIXUVTm/QMG+qxHeq3YrTxbGK5oUoxUS+gUaJ8VtVkGTK7tD6fq5Q5KUfphj
NIafpuGkS/VzbgJVgBWRzCHtk4A/VTwefusl7IOigKxmTVcVx83whnTi63ommlZZ
npjkRGMNouQvDFjthcqPJERwsEhzIleUKTVtt+3FWqDGd/Sz4vUGDiQd77W09mS8
UUyj/JNElYr4MKWcuip2+9xh/LRI2lmxp0OwiSk49iJkMOfSfj7HBadUIZ6OYAuO
ZKvO1YysZxynTEIEwnKTta+If5NhRbY2/gmhQ4Hao0Sa2bQh5ltlBKTolkd7Gtbm
XHhje4+xbScsh47Y3AmlUVOnB6zLplcjOMlidTRQg0oV0vpspFLA+hpdqmPbeJsP
FCeMu3B3UswvVA0JNFjTxc44OIAl2GlWm4g0++00kdyhcn8kcrZuOsYrXZYeLt0o
h5E97P4fgEEBiglbxt4NsE6Qi6hdeL+P1winTOEEtUqXbvk26nwSUkz0ISCFqO3N
RWXWpGS4DnzZP16Xz3MquE2VK1DuOZHOVAeeen2glZx4eQ1R3u6oYQiVL7u47HeN
TTrb7AyydwWYO6BlHOq1MJCBFFtSKhiI2+sIsgP17s7mDc6ikAPhXDtycHX0bqra
lx9ruzHUVZ+QSAIvzQnWGGSPPsLS44W6c+e6ifBeSG9+VZeeqQKkUe7Gt6rrgyb8
/5OwNqP3VILBUhl08etOhqCQKIyvUhUSPpO7XlIrzxWA501OuwE41d35XKKYeUED
avg/zA5XzprlQMAAjAzgFAA/bJlB9Hx0B5qdyxne60/a2Il07X1dJm3Yb5Du7/h/
Kdlb4jybFMQVvSIm7oXu3ZZFS47W2f4+kkxaY7nPZ1MVr2nqo69B8cggL3Cknjm8
rJqBVZ9CLCEIsM6/L3XT07ki1kJR9XO+s7lhy4MAZG63uB/o/2WxUSzNPDsC3Viw
ilgVhP+hyCRxo3jduTSl4LaMDxD1lcFvWX3uN52QIUXFcDluz7daUH1Og+yDQARK
bRDNe3e95FOctcbDddb2kPjbLFjxQC+ot0Cx+S7vlq1Sjk6xHssMbogL/fE6tRPI
CZYuvgkf9hSDXbLOTBGsmXvNYTqNivT8VSxmknHQYzzLnkZ5QDBVnOKRsaX9qP+n
iKCzaLKyl7Ii44NBnZ5VB+2PKcYxzYIuZCJqv1Xk1fV5QvP84zUEg2R5xPU21BJ9
z89kiJDHbsP0HYsbkhC2+Woj/l8VMVMnmvCjLq2UYGe0xOEkheZgkAJ5Fm/wiMf9
/FwTLLU6ISuOqClkTIY0/e1Olt/F0XzuoiOdHmdXG9PEjNBQTNCqHNY8LQgDzJQv
cIsYVhvCh7532eJgdavhBdqVAP/qlVhWk9kGCINN/LITM/oeV2YVS/Eher1ttih5
by+9M55QuZ9MPShn4Iq1AjVEW2ZGhH36whjDsW0yUgJ/Yyy5sp+vI+3aMRdJT/xT
hlj9D2OT1ZLimgML8qauJpOoFG6RV6MJBSQJ6/+EVykhtVUSVvRffQTdoxNDbxiN
yQQ8i/uvkh1JY5i031TU6KGpTQvXIYKuQGtdS5rdA7vA9IL+NyCs0qB4jYUAwmGE
sGMSlGw6v/v5JkCOQ/1K307K2ao/H1tUNWVKNSxZYcEd2xNQF69jq0/GTpR+dJMq
15iLSpij9QsmJta4jT9mFzxWUq3wKxcGoJ2adiZzu7eZUu3h98gna8qXkRkEPw32
jrJWnsqN9wnBYhIxBCQIcPrpEJshU9Yo/ZDita74t3duqt8LnYw+1gqw0eqDPIUk
dPYfiqui3Ugnb/D3haJUOqfb/QRrsaSH3sbB+LCrPij4e1Cg5Xok32ja6mo43wAn
Vd+umTyRk7NIMUJoYuhqbBQSQ2je3jM+CpdjpuYpFXOsjGyuMCELYfwF067UyGK2
r+gHYiVdPjxqTUzpm974+GbXgqU6073e+YE4pxiq77aEkhz9RhPwsg9xyKs65DEw
Aw4nkV3w8IXGiJv9kpNyEiq2kzYA4aueDrsZAstGszfTpnjccWLwzjW/fbBI7NXx
yk3RGxGSL9F/ANRxlNO9/6rpbr45KyYwuk/jBtqDmILzjLXGezzreUPCqXLYdTau
b8kD1dlQ1qE/sE6mTrjZYtRoSt/ixmFCPER2vu89clQVh2MJ6Ge1K6AXToqIic2t
cyatAn8Growo3PwVeSqniU/4+psCQCFzvc9ygyIkJLlpDcxys9hUmtA2vXxQaOs0
ywLNuTS25YKiOwTCLBFZ/pxYGxwDFp2pNp9LlerJuQedhe8+p9bpeUq6CYLpOrI9
9GEE1zTI2L0xuEuRHAZHRoMygf7L3dhwLpQYSrRBrEdDYFZ03OBlXfvHYczKkav2
FtxG/B59z9eCmOmDjm5n3rgvxQOELry4ise7X9ewptAszQLz/sHpL8+J1F3rgh2O
hG3fZMV6qqbuqM6IWI5uNo2reW1oev/Ig/evYZnMIWfR1dXtoAFkY2Kn5CN2qt18
77pW/4GhGjRIamopCOUJ8R9R6s4mnoRoJGl1i9YYvW2mYY/CMGAcZSi8RGML+1H8
sY4xopfnNkx/1ZotQDRIebnk8W1dPJOTpKOIaq0O1o43ApGGej2iynUiasZSls9a
w5ImAzDVJ02l0+A7TGGZhZQkychW7sv+B6YGRHjfrwuHZFC/3YHTNNdN5EB87/Xu
/0/c+ALspyWq734nz9lYd4kCpvUrpN+Ng2b2sRWhkPqe5jqkPOm5VCRMqpbUpzTc
6wvavw03wV8HQUqDC2R/6nF89cgv9mnQ5n0WIN03yO9ey+2kdflMjPLikr3Se0Hc
VTVmnFUtAErO8EwGVxzj7G0GKdYPNQv2is/XebjzTdQh3FTqTaWXqCj6z9AHQHtg
MQW8A2w6gfZUMXf6g9K6a/NctgQCBB4QKdTVYZ5IzTuhbvG+h3NRIPkyHH9X2sZ+
Ia8G8tByeEVQtVjNG72juPxMbHTPfsKTZT0tCFLn/++oh+A9hhtiiEu67wA7Ax9r
EswQTsDHEMfDXQM/jIweX2DsEC7oNmhzCMPUXc8+CkixNP6InnbvdOJcMXxoFGp0
9UOHoeitG7QFAtdsvc0E7ISHAX4Qczrc/BKGYl3BqMhVYc5i7SJEtcYnuVYV32XV
Fmk8zEEEhlaBQPgtGQRPc+6lZW6YfHk1B3NKujf8gql9XwBr3qEHfquskH7t2b+s
V1UAOIdV5ssqFLbDXonX9N+S4vgw1L5O9a+O7eIkgBCod+w/Ue/nTjH3+aMby84q
z1H7FLNQV+jGAl1J7NXcga2S9uSkDD5QGrJwkWx/Di/y7fbQYAgSZ9U4OLt2AXzX
tmc+uCjvDBtzSjGg6Jwsqa5c87sPBl0Skdq9DDk7Y6pG/M1UiscHejTeDgczSsg1
XIZXaiipaczC59S0vD5izH/HtmVSomrfONHMb5/OWdCtOk7KYqwmFNvvFn08Akgu
ZRqr2dJF5Pykwvukt10aoBlIoUsuJgEEpZMFvmMJiVF39l9w3R6CbFMEoSrZy/Vk
N7goNAGIVM+gorXQoezogdBS/JsuL0f7t0zJCiC50oBkPGyS4upyHc3n/mlbeJyu
CEHiCdA+Hfp4Y3lqDLFVetB2v4HsRWtJmK2K1IsUeeNUJVQ+WsSj+NuPVvnD5rA1
48Xvwi4rOWK+IT+B1HJ255t4cpNZzwLyj8+jcyY2e+hYdoVLWxTVbHjvAFbCxcGS
0Eg4KpuZQlcABVOz0ZoJ64nnnjyCuX3NTpPLjuWC0U+Pxk5NlPUEVbUqYxHxDnMH
+YfLRZtvdXqusg2nMS+AFft+8d5LVNdNWfnv7piDRQTw5c5FPRl0TTAQXpBxRx3V
Qu9caqjBccH6TU7KYV182g+uopdASy0k0hx/iM48WlNP2CE1ypFIZNUKhLbXuR8s
xPrs2PX5pB25rc+cHzb6OBsKsbCDQt1Gcg3Od6BclPmB1RFxZgtImgoBrJQKlEIY
O/K4U9hLXn8J07MIaYFfIAccR7kxpnoHcH0Mz7OkY69LXtJycW2GTG11hiUhSJ+3
c8Wnsl3VEAeYM2ui7nQU0/PKRCPhRDKO48ccAHmAFDgKK/lQHLNAUkuzWcGKJAdh
U2eI9S93QaMEVLNCqG7JUhsWd4t7Qs5j5L4ylfU+vWjvSKONEG13GqQpzY1Ghh2n
dgvNSoxi4LSKmTWyXir5M2UM0wxWPG3TCt8CNL9BuUtKbq8u8hW6pCypy9+/9o/6
6Ws+N24JzTgR65k3eh4m8wNsLHJ+lVWgJ2PTXRRQ1kBrwSPpWv+iKYiFf+2Mfd5D
ozAHKXoTQs4PlCNbPyBK1Ipw5UHBGv+p+N3/F74UVomnwDVn+KvOK3lPnL5Tb5ya
fY4Fez2Pa9nL20CZVeQuWsFYNzbtppGu6fD7tQusVUno0oALI+h4sZC316MvJDyp
CNa4042nsn3ofTEh87IgMAL431SCwBoBOsJE/W5EMFL2j+RHQ6CkcilNqln6dVIE
6HyeVD9QoSdSiApT91jyW7Po7P1HoR3PBUEsKlEdZqinv1PqiUucNrglwj0x/cSa
BMNB79/O7Bw/F5mRS08x0Ni2pDiV4cJumLf+DLq+LlM/Ah7bYQjwOr1dG5lo1klC
pbZRjpM+/rMADSkG/5/WHfrjlqWtj7GuIQo/tUqpIh4d+i8WfcRh0Hrkkxf3rxKb
uWgu5cu992P3+RseLikmCD1oeH0wqE8E5Y41GTKhtqJjfswfoPnvJPUxW7lIbPm9
JPcIMmB41xyMcHLrJjDpB3vbLc23aYUiaG5kH2jJOwG2k4kccKrP2tM6jydNtp4z
0MNeGVnt4Z5+ml3pp40TdW9TLRnsDVxrEg5f6CNHWHCjWqVr8YOYb28/IJM0h7Dx
blUCwMQDvQG4/9PQT23RNAq3vpinG9NzqQy3VagjIXsBL/LBp1HEbQwHMIsKM2GC
uDhzSQ68Lp7XsaGMhT3F/trD9jbeeZZ/m54rC7Guvym3fBoAsA40gOgiTAuXpHvL
7OXAwT1ZA19aoeT51yiUoqh6RRij0sMopS1D/A4dGg8QqrPeId7Imf18MgEhrmNy
teh9486oayXDju8x1+6feiCqottRmnSAS0MjOG8tAOSVq8Gap5vPwofI5DMpPVDz
gSVkRvMrDbIlrkQr9phObePjKpsdLp5wuMAAJtu3vwjkNhzChWUFOsNxN80NbwND
h6FAIO/abQUit53Y/b4ftlzd/ruK9x8UczesuP98ZYDhqNgIGrmSTsFqhTzzlkg4
8bKXBzWW0tiPwGGkBt8O8g/1G5no0DdHk5AqRT2UHMEDXj3iQzfaptqQAznDqL3d
Rc2hGOsgOMmHj84SxPWOjLyxfSL3f4yDqsK/qk6iO2uMYGpzPfUUbhYds6GDLO26
KcOsTEcdhwK9gx5rtxEAb6mLf16Z6Zco+aVrWPWxi9/D1FArXlQrGEYREQxRHFIU
cK4x1zdBEQbYGBPn91BqI1AwOq8Amxzp5d8mwCcOqI4jSPAhnn/YpWfV5YH4JibG
4//3vler4q+0j1zPhP0vRav7jBBKAQgKHt8cwvUdZW5I2eQkldl8n60lFVzoGE03
Dz7QGUlsTVPEb9AR2ksAtWk4J7K2vjVEijwe8YsV8jDdAokXQCU+rOBRxQjpmWbm
RM2jfLE3K9YbPwJjGWRxayJYACkz5oAGds8T5aGFnrftf4uOg95vJYaZqVmr8qI7
Rr/h0e4Q9SeKEIdl2X4Nf2lNW14OxFa03a/qQB36lJIAoTKuPSTlrlFBFrDIGN+v
PT8DDTSCBTwxiRJfkOf3RKNuO8SSPXYSRXV3W7u6BFiNlqDnDbepIfXCE0Eska3e
9piPpVfcXnfswH2ysefR6YpiJfQLZH/Wz+O1PN1krk/jAIchewT4odIy9TIl8O8W
NKZcjYRcdlNKSWjJ26H3HHRU3HtgfgMJRP4pAYVxIoWl8iT6res8xwnhcgtVPo5s
t5KPUaWh0NPZLGDf+cMFXAanaC7QqftDsy6dSL90B8yPIzdP6XZoS6MEISo37k8E
616ab+4cJaFFI1xVvC+QAI1gOG6tNlyg7pN32NByO1Sg+60czZ4X74yJOp4z8Dbw
nZaswaLEiflRvtHwhcEsEoGF6wg6tL5VjRBRiGbdIOcQOK6diCtICHt0C9A4t18r
NhTkRrM+I7BBhyjaJjxhUe7BQ2zuayC7ZYqd1rLHi26pA4k01Xv9XjinkXne2W0m
FMCtsVRZYK3ONdA2jU1awNJ4GCqvoEFg9Q4LfgWQbZJ2NZ6t/gSs4maYrGY0UlEq
Ni/oeC+CKBxSkc9UMYGq82H+js9F7TS5ICqdzbzykMId8fS1Xw+IgG6GUrWdz+G8
W+wIr7buFbMIS9c6yMDA5rrsTPD7kDnv96pUHmMY6g218K4cCiHrVlSba95XGQmD
UQs9ZaWc40/LFDoWV2R0sNkYwnujmaT1ino/1LluIqJjYhhdUN8cMNJGdfNpmmga
v33tP5Zd90lFFx16pY9ueGDrhgG4uO/MqvOElN/OAOf67Yy/M0abd8w8/r+epV9f
OJEaGF7pExxCa2LMHSkIp5tkyOL1dd3b56LldZMSn4Lb/jWYPP5zuQrXAHta0YP5
ePzF0fbTG5phQtFvuPi88hz7i37PYjnaVKKhyXxW7dT+HumoQhSpQbZzWw83lCu8
GJfUQ8BOtZ6dfFSHYNKoOPz7kxVeYQWxnk1txUs0uJBCcU7F1r5/E9goGs7CFnQl
P9vtR1eM7fDf5opdCMEZBaaMGWzoyaELjuHXQHPsCW1Cd745NX8ykloZiKrQlPgu
c3/t1NoHOIYs8POIUH3FjemBumjzL1dQwj9/IGmWBULnduvsUCmOshEbeqp1wC+D
BCMagcxTHi/kqsfiVA7BMDkzwuKwiMAvwGVQmYVIsjK5QqidG4LVnpRpmZn2uiZc
nuXJ07PbIxjfJ11FJ8ecVmDM2TxavlQQZZrYio5l+gcb7y2mdLX2VncuKbJDt1Yr
oC0GnAmK+7GRHpv+QVe5xfAdrvPdlK+JbZKMHUAjYs58A5m704O368juP2Ot/x3M
8wCqAdJ2j/2d3y4tIolppNo4vw7cw+Ue7lmCogZZQGxwTmejG74VRgdzkpWjg75i
gYEvEwIk5FlC6Lf89LqZByWY25UZAKuOb1ObueqhXBSqmC4nxKHTRyzE/ZsEpCvH
vHqUFFa3lcAJhYhGSz7fspkKo0KKfvUHMCRVhbn4tVpKsuMCLzL+dlkOX6WZwbk9
MaiH1/eodyrHEmio+7Y09EEFlV16BEmWWyvqZrmqDS07MwYtEbT9qg9x/9LXdK2X
nzbuInZ1bmJniJgqzmBnvo4mIlOWa8MtN2ky46GGAdnz186iH9E/3i2rBd6gnBCb
gKcd0NOatGfe2R/2Ym5I/trMJghhp8+BpJJoNMJ5ulRpD32BnhTLIcBffBTy/myt
JBADGWm+IBXRydfCuv1clvignqmfB3c0dOukvdwtOg8BrcnGF4cSCuuO4erxpqwJ
xr92tWGRci6NAYOodhpxN8XDHmrI/3Ulfq0EALXcI51hX0xDZfGN2h50PRGPHQHm
KE9r38yd8mJKCxn9QzFRjJi+RBzc2gLUlUam1praQIXYpwSrl0pfjAkogX2j4bCA
LjTWl+2QYfdW0YLyZ5FAYQBobFd3IhmbRDzzjR21CryTiHf5R7k93gZZSgISD48X
Fsbj1mmL9GHO8o4cylD02HdRfh6X0j2RPf+BmegHWozo28Lg8oQSn1hRlPFz3gI1
Fq29aBSWNrpglWyk92n6MmVSGNh+tsltnODdOxsBhTrDsNSHmNa1zQgIT+9mjfc5
LvC5pe1M7RdgcfoC3rTyxfmyf+cFKsSHj8cy+3/JdATHsbgJwB7fv50iIac3dzuA
OQIxlylwCcCoIp9/Ib/XTWhCiMUl659nRys7Yw1tRLDALXm3ZCIoNIWwEcKkSMtB
M1Kdw4JD9hxIbUgZLF9gylMkhGOajvvEVuQ+/yTBPY4vvaAaVmf6gWI58Ey3ZqFK
HMOkqPQAs2i+OMa0Xb4NMtxlpojwgxgzu6Re1OL+52VYJ0XQ3QM2p8cin6PoWNuZ
LQtsOY0gLK8MCmW1XH1XJtFQlfvO3ngYkMx8B2yhEmJ0HM1kfIYS84isJRuivlAE
9mT4hqiniJGlC8IuVTa/eWzkmESXZMALXdFZDsxg4udWWx9o0Y+7HWqPpMHHHSNs
X6JrVWZPIRwyATJtpE8+7Wwrr1IPKwQFllrW5pvJ5j7TguDNRndAkjsQD+SXJI9L
lWmY1zNiKsCSXlXbUmGfGhFSt6i0Pw+4vzUwqXKiyEfMvTKT3/SRNTgc18VKHKjF
GwGlKlu+HEYNhz4pVopWBZoTSmgvKzwTFu5c563gu43KE8fpkaprY6l+fFjN3p4q
fCofNHMHcsQyaqMkrrrIIGdn22X7SDv4ZBHo3e8qp1Cz/2Jmlb2wFC4GRQlWUD0C
M5QFXR06ca88hHasU/k8sn1zIuJ23sinsewITaybfwuEFE/qL/LEXzqsr/uDhNz2
Bl4DvvdxoKK4yQsms2vMmzIIx34ZUksg+LkA017fFZEeRy/yAdhMwQ0oV/1iMMnJ
XzgsIaM3lufytZavATyh7sLyAjfSk1OFqKCDItV06DQC6EsVfmmFFbRB5fxqWZ6n
Xui4oZPZM+corsjrXR5gODQn/kBWN2Hi0EjzVLk+El5WNMiNDlL3CSqwtYnBxpt4
3mSxcLc/2/UMwh8rjrhinCFsKxPdM1GJvU0Dx/lTjibDRvK3CreeRDWtr5qoG1cU
LzLhpdwAwT+8OXqMbjHKb71ctAMtlnpQMXx9//5p8SctL2C+LrWXKl6aJcf3iPM+
ywwm2Re9U3yfowrZvOPvmSGQLEbuW9xX0Qy7QsX1Z7ZcWLKss7TXAq36CkDXKOk6
9DW1z8c7r0js9GVwozei5jmGZp6If3p86Od0negf+bQ0O96IugCSon5UEwAqn1jD
vqQoVEonYarUzxJjiLv5pu+7z2VB2w1BRgU61IfFqVQ0aDOlPe2T+n7trsZ6s5gf
LKAz3xlmuNiUFvLsaYg3AziRf6JKif/A3afu5qT33nkJJPVsyicshskB/pPl3waw
iNDW1nFok29rAOT4G+ahTxOQjM36qD0MiPveUY7ZPsxisfIQq2sj3WHslJ8CG/L6
9knlnp77bY7hRRCyXJ87ogzku/WZLKlxG0ikrVFTfylNivYtxKgHhwAmfs+mIQhg
xDHcb6C0jFHKujBM7235aDECbhPVVgHAzEAE89Kw+Rp9j54Vyir8nuwZde2f+sBN
+QAZPBgchuuhrtDBykNx3hRI9wYm3/ZF7VgipyEjNpVvuCEzxdoS2MrxjhO0kqki
+qjT2F16FtkeffccTgJMe507HPXIJse+iWNHq+9pTZyTNKtV2RVQO/oFswUzbgye
QYCSoLeKL02jdv88qMeJZbEzbONNhqmgj0tHA1anl8AxgYlZrtrYo7UjzbAkmHDr
H3zkifCqMTzvcdRKECZdatPOG49hloFfBnOKyMCT4ygCs1Yz+a19LPbpL5oCkiSO
WG8thOrSTKjQJphsKfXqEiJiIIDQr6oN07jrlKeEvlZxavLb6i+ZXt/AGi2vbQj+
x4fLjDNzesfc8SScADaqNExgp84regkkh1xCJr1F4l3yFDeY7VNtqrPzFWiOX7nU
tvOvR7TB0bW5Q+emzA5Ak//v+V4DQLcreKtJ4YYAOq0VC4BoMv0ZtPt3y+4ub1E3
D/Tq5xLpuaMVt1w6oB/tPVlVielr63e168NSNkPmQiCqjJtvctsfgBq2Eu+RMC9O
wRLnK14vOUvnhRYDrQprpMcBWcYAea5TJ9MtJlkYIVfAnDrpOQqoIvXUDxVjCIxR
bOWMfdyXYwJpvRTNPO/eKF33V+lIBpRCapQfXh3khvHeCNAE0dWvDq45YJpftK2H
A235c3T4/1pZ3yCoXMu0/0iCmduxkfI59zvIwvn+R5b4QWVs+6hKBq+FYo607Mob
4Sr3n+xPnK0qq/bU6fPyAU/OpLlRGfgeWzmfR5vOMBkaflz9mMw6UMgTI4RfmiYs
mzm9gr8CtSkuSX3QJ9LBHEBUFPwEadIxOqwnQKnsezZ8rTVc0RahKo6/WeAfmcud
c7lYXd8o1yqrinJU3j/wdSS9sDb16gmlp+XnW8gsI3F7J1fOgVoIuS64QjdaYDD5
DSg1jF3Q89iEZ+YmabtDZ4TA976zaqFExGHCPfvG3jOEXozjO+y/SujXrXW8gGsz
kRAH41f9+tAKAFoRdpKh3auwNYPlYOAt2scJ+zXAbJVItgq43QMQiHU78KWCbPEu
41J+jg3yVhhq0t+q6XPo7StRMLThfaCNxxOtKy6UhOSakfVVQf2FpKV+etKm0dKs
/GNEQLUjG4ak7vKBSrL2ovjfkXdsJlZ8+9Nck7JDhxWVCOyLb4zgV7N8kEMiU5Xy
IC/Ne3penVYjAeFo/w81cLOIVnVGIR07TXUyU1LI0fYNACLgP9ltYnTbkY3oEZDQ
O/KXt0KTN7YJUf0c6cmpCg0W/wJaFyJ4sELwwOaQZ5CGJGxgTeElp1RwJV7pF35J
9OCgMjOOQW98o9Ljbgguie99oOChj7gKveIOu7xGxzlHC8V/aPQncseq7P84aOPo
SF0SbJb/vkKhNpLvnOb4ux8MjiQhj1jrr0kU+SA4wueCSZQ5y+yYyx1yLNDJX/OU
a48TDGgHqC7HS9gS8ZOPRbEVVps0DRUn7WsQ/fqFUZnDC7sQBVi5SQ1Ck21CkLd8
9UzaBHV5/QBFw676X6DHftRiGuGQTmuaZM0XI6wvElTxmbwN4U2k6cgM12eOfqjD
EJn/zNhP6rh+CzkD/6rdYam1LvrXWiPFOCyVWent6aWK0PEmorY6uyt9un1tMpO/
1xYKcqjogp3wWvDmm7EMADglZ/Xoxhq8r4n4LqYyLtu4M1HBU7qhmBbQSULkk1CP
eM/MA0O+xcDpW/yzhoFFxaVIfVn8CIJoKKMZCduu5NrKjDj3idHMJjWyTtyeLCfT
QPXV3xXmNEr0qjIPSveTEw89bR/UKNDssyWYfAHQ2KAwXBSUPzDNRNo4V8DIiWpa
xh3hl9fVyQycA2L0ollocP9pJU7Avlmrv3ibh3L40ITFOBS7AZHu6eMx8DEZJpxd
8+U+kVXJWIS/LAMv5m4WLPvr8twmc7ZvRJeyWldy5MhIwSH/9AjAcYANFvUPLfE+
ivni32qG/r6qrQ1+SQIFulYoMksOT6RJxNW9kwiE50eJ3OgPUkOIcP+dCcmDHLZw
7oIx1ZgN3VZpDtiehlxTVjOYjpL/Ca53olwyKR/KX5fbnTR/9EbW9oJVRE7Q9MpO
E2OOkKGU6+iTTJxATpfSgwqgYtV0XblrHf99tAx0D3UAhSwDL3m7UcE4K7cDITLD
6WI40DlZNyOo1g4XcrlrzRCsqVbFHibS9p18ud2mzwpMFHbA/m+Okq1kFvt5jEeS
/9vxE2ApnQR9ayopTVVIe5YDbO73EnBY8ugJgXmZHdBd9q2gdnQc40uq5xnWfeh/
miDoe6S6nlOKQ9fiynGqQi9fDnj0F1TkLUX7BLSQIgA4en5HGWWnHc5Fb05gxn/f
jGLxtzllVTBxNV55JLB8mUKqfkaonRk6jqhBq8OW9E1ZIC0RK/+FmcJVa22WGwkU
myow4V5PUg6aWaD+dj/Wf+flqJ4q19mwm+2UJ+DY2ncuSw0g4YuqWb/aRKS75svD
HBsbW1O0WRn4M68Ka14rYEvAp7KrCG7+PWUMtTjvyQpLkMm9NpKFXNHS6CdtIFUI
hqUVHSHalrXmysxmLZOd3YlLzMYoD3NnVwW52ZthE03RYdhAwdpYndZW88ZnH7JF
3PLWU4CqXWhn2UXUXq2TJ0kRr14l0IK/AeGvbXXpSXHZN02bMa7A80skBq+Phqgb
O/1purlpFBLCZUaNxcYxFDzZVnT0DP2OgCM1QXRXjceKKKUtJ5yWRUM0T4XX6bPy
5aWpuSAaxy2EEGkXYbg62bb0hbFduym5BdJCtewc1FSVZLPFXi7XqQmU7gh1rAi3
bhtnq9ynswBrcMwPJt5sc2LnSD9auYXBhMlQYOgSHzs7k4xGJV3/qi30FoG0RU42
bcPubG1j8r5/6/GHG0lsT0PTVZ7AuavcG/RYRo1bZzMSTHQn7lulyTH1UjxosSnA
OVxICiGkm5oVWYei3uHuFPqPIIoX6/AnOmJ/GT+pc+GL+Q4rBDRtqZPwQKKrEAtz
yxYcQ2fCuws690zXvYeT0YL1Mkl1AtiMkBo4pImBrf2DStkIc3arU6Q5RE6vTLRc
FovrL00irBRqh/DYStmavDkx1pWSE6FDeW72gX855Wgr89xqwgkPwcL+8qKwopYL
iT61iN9RZptPpoZDwqAyyZC0Xy7do8kf6gPnT5A3MwD0LFFW+ZGs4VAhqqfV66O7
hsL6ALx8OF7R2rPK8/4i4rhUo8qvcRZh7rjLWFIW2V1vHdubJta2Q3zJ1u5A+AbV
/+cxpkv4+PGDtbH81IU2KqHIOKOb1AixZMGXFzBUu8bRVGY/h7TfRskXkgZV4hgu
wyNECaHK7EJ7TRGUSAeBoWL31fjbsxWzFB5CZIVxmdOX20+m4S3wjq8T1Uv4Bbpl
F86+Eh+o89hcHx/JT9gtv15FsqrjpaCwY/S7JR+wEI4+XwT0yuHjS3nQ2G8Ytk13
RxnfEwisHDtdTKGtpj3h6BjQv57oYNAvzfWf/ir6PQeI/PY++QarO3OBAgl0S+lq
Dl95M8vjTqxBLIP4iF9Gs02GUWeXbSQ7G+esZdBveA606LTUlw5/JSjSq+5rAqqd
5GAYn+m8tX+xn1OR1gPSPXriB6Hyvt/5ZweRG2v6XVz3jS9xlUSZVNj98F/N2uQM
pXW5cHaPYdcAVlx45TX6gJdsVrxHvkYn6w48AXvo1QRNPeFSGXm9nEAK77AFN5VE
UKJQ1Wkso5n3T7wXQMB6xIBnyyVmfir1UNbpuMCwyuRhesgdy7sCUP9dTRXeONXq
95wicMcVbEXfx1FQpa9wpxwyJ+pT/nW4B0hLkqiwG7HeFT5IUmp7b5AaUcIMcw4i
EynQffGXtXRs2r+OVwu/PpoBKGE+prTitTj/krlhNLnD4QOAisQZwdr/GDSyqy61
kcxB8zbfTj+SPO7OF//thg+yd8MLU6I4ucZ/cMTaDzEZCqlXJ0Zjz3nkSJKLeitS
4yarqB08WHYqweGaM1picnIxLgZ+F0cAvLZiLeSyEbMB6DXen5yqt6pXu+C3b6zO
s/UnGdwb0eMTRyrNFo+2322WH9BJmMswabLaeltxidToMFRe+wTmt0y0XHE3U5ry
srH2cGRhnMOH6k4dbTE3PbDdA2B/DuR6tzywE2tbDvnsiprOhDu4rerJYALMtqMz
ApVYuj2pcSNI93X+sjiJGJkPmeW4fsgNYfqCwDx2/Ryv7DFXMCj8zUWuXRoVUwqU
q01sMHIxHHLUCDnJWKgE/owM2+Eu2lJROUp6umIz0R8JbjkyZZEzgnN5XY7j4fxm
kPNjFXjBxzqCYtmHpCn5A6foGadbG6GZTvK7u0BLb5RJTquH9OxT6ebGjkbqW5El
ksBrwa9Um/+wDzSeG8lR2/txN9cLUBgnfSBH2iCOZq4p6it5haOZ/7dntzaDoG9d
5Kv/H5N8nh+mB+Mo7W+/j9pAOZWOn3rqR0D52+TydnIz/iQiWIyJBIRWmMY8sT7S
eZPOmKc4JRoNN6l9X1ZgofZpAT8oL2e1OwkwpdPCRP+1AkWLt0MRhlKkV2ywcwb/
fvaXnIYHDKQm1IxsbsEl+GWZAQ88sFoZg9dCWoHqFbZzB2knosnNbq45dWXES+CX
bFezE76K1ePKvE4oDR/vaXLsm3M/Lxiw2Gc4io1SpjXhcX+Z9//+FBW9JtuE3Jno
l8PzJyq94U7AQWY2MqZq5eqldra5T61e6I4gmU6f/4I8J4OJoMNkpcI8ebJbt/CB
Lap2JKk+f2kvCR/qaC40BaiM+gxc5i+4leT+NL38Fcvc2T56mUbj3rElBW4U0NB/
Mz7SQTgVvpRaPCPiD+xtLUkNMjzVRUaiN32RMLGTi7jz+SkOEcksUw7R6JNi5h5I
NLFNYMvujJSA8mxk2M5Hdsm439bk6GBSSQphRNjOCFJY/jInkgFNbdPrMrVSzFOH
dRE2DcSc19hRSmwwPpwcXFcGqYAGuA4ZNYYH6PVpwuGJvNWFZSPj0V7lesXUNseB
Vwx+VlQsx2e5MfaytqwqdJVKIGDKmWjMK0vrDuZlQDYMzSn/V2c8OIvk33zjqfGH
6Q8NvqROf5zjUPzNNaEfZxISNKfpzQ4H/tipinpVN2F/oA3Id/2lZwjH+95rqEFi
jEByrP+6BFwPy228Foac3KcWPU1uLMIP4rSgTa780YodABQ6iJdc+wjVPBRKx13q
FahDR2fsoLIFKIoag6Qodach43a940s02t+9dZ1SVsQHdT4u5w1cZGskx3gN5RUh
LeJJfEXIGVRIsaFxKOpEcrcr1HbwoOSVmVWdi4FjgztV7LRVHam+0I5ufZ7y4OTQ
EU2ajsVbkkPu22CnkGSjjgoHvCp9+DO/EYZ5Pyf9AbWO+/2PNft0VXNL6Z1AKk4k
cOFOdDu8Db+fTthIrWOoPvptcHZmrymd3nqLSHB2t/ovskrcTb08AP1ihkx5k+qU
zV3uhmhPkGO44vmjpK3cDV+VGyfIIgBNzeE5It7JowZYefN9YrkN4cx8YVdn49lA
anxivKfdM1XBlPOJejwGXOQSzCmAHOUaJu4EFPme+KJwo5N/qla2b6CR1/3tXJMk
iVBIxpdxzhVgKfYSzMvUqMAlpc7cbAnjfjeUDqifma90v86zRNChDkJCMiPN4seN
Fi1BFp7oan50KlY5169Woyq3ijuQtGrr0tlurS4w8rvwlLz9hfD6RJ+V+D676crR
xR8XD8Xtd/3VSI9BcWegCY2mqfYANrYxBK9Sj5EY1dJZShPIWGg24kf8jcN75hkT
F31nETOQRto2JIh9YYKVwDGSoE0u5bO+HL61oinwXVqaSVeWCB5h1tqSuXXQDLhF
1BlV4gdElceaxIFu87+ZpA2oysBeoxuA1jN3uccDD6HA8DTkZOupTE1b8FD1c8Y0
iXaL3KwxaQAQeXjOuSvpgwJs+OYvZIfVXSidTRGjZHWX+E9swFI7QLdjKrpRqeU7
1l8r6VKJCqc5nXWJJDh0ZVU1dF9awLzen+ZicPqpdTULIt9batgSFaoIQP6JDSm+
40YsnpqPQ03n0kHzcpQmbOE5vxohw6cwHF4RHSjWa0CahDZlKDyOIyGcSgVn/nQV
LRqn3LAme23R6Gme66U26LNqmz7nsFstORIZR8EafHi/DYV/uGuJOZQV7ZysD6ZY
+fuposGK4oktMoW4CXNB+sDfEI+yrIgtB8sXxaLjuctcrrBmILveJB/IXF/OAbSG
7wN8xuLqJW3PEb5gQ1Nr0lR7p5ePm70gPhBFwKeDCGXJu+pIPh6c4QluPSbFQhLC
9uvhe4XU5Z9CDd2Lwfj8t/B8KMtB7cd5kGxCIO+dXUIJaJqG6yCfN+nCwTxop3Jp
fNf0GaZH35CxYhCFzOKiSLbTRpikRKSV4nPu4/rMCMdm+q9OMpeeuD8AbTPfy4oC
px8e3oCANlpFib3GXn+heVSTjCr+bJhi7tyx6jG6WJjsPDtejdZ+PnKDca+YdmIT
94P3ssFMMStzQm++VlM+lY4cI7Zh2FVJAzHe+Bwcw/eAVzuh+lftC7O/bTHWSWax
PbNlGyP0umKYdAPWwp5lh8aL6Z2jL5d7QKz/SVBttoZyCkLaexkLPi70ohZwgFb0
E57SL5oxrrqh3Z2E1ocJzvMUp8uJQU5hHcu9uZ89vK6cFXmKHnUbqTlaAnun2qyh
DxHX3qwn/Qkz7tTyD8UliZYSic+nM+P0hvwwFemSbHcTec6Hw/kgKB1CNvpQORKX
uE0vxeCpQxF+BcOP3zE8O8rd+QHJIBCHdJvz6d88OgpyupMFulg/6TQuGxGQLdin
G7C3LW52gvzevipFj4k0qNx1o6EEMh+YwhfbSMxfJ+y/dxajENxp6g1KNb4i8ETH
1XvDiox+CjaWQuzLpUmgkA3xmW1ExjYFA4Ir5cK0T8okkAiTDBT1IO45FTTNh2W9
Ci8NZ/YbwQzFHdmGGwBpcMQSzhOp314Mlep5AVMMCmnyitdL8hOnO9N/SZnxcHkd
2oeKfDJFvCqvgzAJpFfFO64/RKXQfO7LNtSCNmk4CahWNg2h946w6D8f9+EZ79ls
Yo5rr2StyxuJxJ3YxSRCTaX0Zjw8IGPYZ1Vwt244b0kMBogVw8cAqosSpi9/cnxH
oHxSogTjfYmDSHY0k9r3GaoBinIoxlr9DXc74xj16cpu0gGW+ETdXwYZUhJBZ04a
bK3APuogefqMKN92tL5pPUH8kc8e3986gAzDm+etgRNJuZUKH9WoRtFcuRsVIy94
KmUQ9R+xwDfmwQwe8yFqq4BVOnndZ06ZOks1TchomoaRXvxr3mOagv1gqEHsUGZK
MCfnzsO/wTtYDeF0k7DUlQSF3jAgXxYYzQGnNlT41q2OYOV5o9hPmDZe45OZEWsC
UiVezT3hhdz8QPiuMtiM/SiHSFNrlRfM4a1fs7Uk4hrzPFJifvN0/UPH+mDthQ6S
zQ5fK5yAQ2pUkI+KvtjCwcWwKeeFTIU6e8WuHuc7638zr8m1P+Y7PlUwFbsfuPLP
e2s/ZobTdnmwJf5DMl7ZKFzNu8qB8PwWS6k2G2/mHVs33sYNYMLTOgfNQQ7woMn7
L8cEruHYnoB6PQzDOlhO3WwSUi41a4dZx9EmYEcnTP65shHyhTp7VEjcd66G0YX9
RIXPb/xmbGe2rv5YwdsV7yJz5LdVNLTvMzdy5ZPGCmsRaDGHapHNCuxITpNkMka1
iKI7t+MbxFARZtwNGXtedLxQSRrLCrPWZphMDNOEXTT53wiQ9cuosZN2UrIbm4kH
yorlkW00SWK4ARI3OLNGsSbApLbNk8La+nXcEKLDvq8hZnidzgkWNLgIWOEZyAFJ
WRtuCCOk14INonsRoXAYO9TdqAL3mhQqtEVWvhAN5LAWE5FJZ1w0tlSH4a/GEPha
FfWDjAyaGFoBUNduGE+xdvq9vlstmmEKeTqYzjYtTadH+2aEW3kf7JsXoxMIFlyY
X4dnluNusIpw1aQw/rn1f5kruzR50HmMzulE2zPcmv+8MM8mdxkNFfQtYbQgFArl
EDKn6MyXBIl2akMGAas8rKqvL2oFFuOl9gAj1L0h/+kmV+Q/MGPINO580q/DrigA
+E0yfsoIEwzucGwBubfFIYbmEua69KAMSZ2sDFNvmDLHLm8XIcyt3cA4OKYogljt
IN4P3Xq8fSVjk+Ks+LlqtgzT0xRKJFe/W8rm5PhR3g7xoQSO0vQ2gExHCry7BwkJ
6F85CBDETWL8nhoTm5lGpUZAW+zIm+sPlZ0S8OkyH5bm6auL7yusHcxSqaCaMwjE
IdAvxR8IBOTQ3vIqtq08LJdEN6FLJ+9V4Tj9zSKe9wIOGOSkH8oplVqDNoB0M2Bt
XEFSg3g+ZPVmUujFHKAOkUoqQon81q1+cqW5fuREVTPEILKtLTubKo78BMftmhgm
sn+YN/LYDCX57BNQE+EO7Wc3BrF9lSia8jR86l1yxgn6RN4VPcA7Vc3IulyAni6+
TTozevZ26H2zbAW9cfwWHIuOTFIfo5WXZBnHCDe/5Eq3u7JgVVsH2Ki6FGNb8dJ5
MSimWSSbhIFlborB1tdPjyvMn9j8Aub7uqUZE0UE/Q4KJNFuovL++a37pupqMSn2
/DigVZGEUAG6MmTg8P+4PXPxI3uIIPrwpcoOAK2rN4h8fe4VwolzGpu3M9r1p94j
laMOsMdDzlJN6hdIZYED9fJRYFer5S4kYw0NmRKldCaNbQTiYdFllQ3A2OOKOdEc
Xjh8xWWikm1qaRGCMKHU4Ss1w0fDE95tI4VH1zluLlKuBjcjjFS20D6u7xBOVbaf
zCI2tnTow3RETIUQ8ftJzMBulxIPApyz/fqgQNvnKAyKh3rZdyZccw5BFvy6K+4G
mTTTehq9Df3cI1hTqcHaN1RP2SYVgLvzoIhpIc8um7wUjeqx5c5cg9OxrKdNLYEf
DMFkS0aC2bfm/eIiexPdFGR2CHw72R52gwUFnMaY7R8N7+Wl34ucHNPQPuIFvgEH
z5mKBIfD845UWFRzpK0/yyIhlaGWOeVa3NSjSHltoW7Tphg4M3Q4XnZGRzQvzVqs
n9GhksGGV+XJ2KdBdF4mR4FeLAur+rlbfS7kPqmgOHz3LxSgb/ppkP9FER2QaCYM
j+csBfAig43lkl5BHkg3KJFnfC5q4hXIAiDHkC6DAFhc7AajMFqm7Ga2CVD1jhJi
Yx9xeCtRVnZnXfpJgvavu7WXP1Tp7/D4pWNSB3Xp5sA6cy+jtRhpilxr3Y7l6d/Y
3tdQ22BAY4SFGEXlWoK5AuzEkdzqhRx7SXCTQBntsgRzpZh1QoWL9kuyOh+lF+Pt
TzGOxj7ARbkx1FCmdBEWK13vCU7Y29ERsvcsBTT6MEmI5z275zCX4p0GsUhO6Rd5
ZId0kzmVjiMZ7s+1TlBATCBJn+1IcbBnKFzcr1eS/QkpJnrjzgan0cy2VM6ds5ie
Y8YktXYCbijOYDb772hEMErap6tEwjDLhjTFMLbU4jjFharc1dZrQ6EI/3Fb2mhG
FRiYU2pObRbtXv5Lcm4emHc7jxwzWcFvPTfOujb2NPbYo9PDHBz29WTStwQylxcu
LO1jDXoR0jiTPpmwKa9uIOXjJMF2l/BZQQYOtajP+qOlsiMFmd7LrjRzBmxmPkdy
W2OmrHPYZA41pnl3QoaJvFED2vLMR9Roqz+q/jMrQW+JBRGsmYGOVvRe0aQI6HJC
JQ2LDV2TREUcDIrht2Aj5FXmNY5TLWobesKQIqW7sueKFFwZJcS+/BTgxN+fhElX
YhrLhmwhP2tzFOHmMPWgGLJJ9RVPYrN/FgbXuvjbk1w6BqphjOJ3HeLfeSwf/EV2
RzLSv3YusT81wh4l6t9/YwfyMJjdX8mi4o4AkNV7C78+HkX3Y0ivKTTbTSYiVVx1
mZ8DGojWCkOGnE7WRZKpwM8b0rvOXVClBlfLk66J/LMYtMRG8T031Cmype+gZWdc
8B4w4q4EPs+b0spd7b0h4NQE71nlkfUTUmmbJiYC58AynqGERjaFUG6L6NIVeuwQ
dkXKQvIWkVp28meF6ncrIrg8IJ5xzUI59aR6sWt/Gz/bQBMs/Y6ZG2DHQ50kzhLO
MVhMhJ5bmzsama1J1NGuFVVw1IN7LQ9OEQ+EGdXfgErjYksWuqCLv9lbzcQyD5n5
Wop5lltgf6GcI6i7+HFqYt16G3W3W8mGLbVjKoTEfD4LvBXhUwYE+JstknLzEf+o
zL5fe6K4XddA2vltfA5FgCPKcIfXd4EGQQ7fCSkoPEJlpdDd7me2GNndVHG3chRw
ng3koI1QxuH6CLGH37r3O6IjSqPQWYjund1NdWdeQgt3YmEbLBbiGgdKUlZ9+ViD
NAa3uJ9CAQDMl2Er3WQb5VXeE2Psjh/caqryt50Os6w2zxwttwjjrBDjs7vMsyJw
Sjb3cWSVAZYvuXFHF/aongara/sup5KqDKyALM3zhdhXBjMhHnUG0TJ7hFbO1LZy
oCuJ6KeQcrCATmTNYzkoZq42nLSDogd7k/pbdOenEmXRmOBK7uPJFXjNQqmRDN0Y
cbSPKLBqHEBmbfP4/SOJ+oZ/8jI8VkAVFdJ89XCou1vy2L8gQQgjYIu9qVeN84X5
HJhkCksi49uuJllzmk6KDIbEDO2HXG0zkTmMSqGOotgHAF97CZsdvl6JvPl3vItH
hFfthwR78JPKlkshBhiewRuG7+z83MnnhkWbZ+5PF9TUeVL0IfT2jLgFOrzsnnz5
N3augK0LuXs1T5eEmphkQwMavYWmPeNXS0Nm5b4eeqIyE1WfBGNlBN3OF8El5auP
VoYPoQ1+JcOp/sPPA8SxBTdJ1mzQ4wCIvcBR5C8b59ssYfJOeAkaDJI1cu54zSDG
NGBGmFHtYvzigjLY3zsC/WSbhSO1P9UFk57YvW4FvxyNziL/I/Q+KGZx9zRnAFlC
Ptl9dodQn+Yt8fETl/4tcoBoEEtKFe3F6zLX1XvcdSbFF7xrKGXv523nLn/3MR+Y
E7OJQDXYAS9xpUDg4bgRITUQTuTPXDI+xIa8cnOzcTmU/akwUaBYaSnyBWV+NU69
GQmJFx9Z5a8/cLAoAWqfItW/fvXIQSsNpFwzn4biDXJ3gaBVvLeZQ0gchVvZLOEG
Revdy9inzjJfxrFEERn3sN9+uD8mPmwpNSjbg/La6ryI0S2o3TbKLM8F58K21zOh
bvG8us28E1puI+stKOi9kqeQWm+sJ+2FKZyetiebttpBZv4pew4UMIdnGkE9MDLT
uyqCdYiSMhEKh+Vev6qxuC/LJ0XBuqGBOdNf6GH1JZrA0NHkfa23LwmWhZ/jbh7V
PFNL0gUdgN5qAzzZkw+XNAWdVGTOlywwMBABYY7sFw0mzi39K+dvh4HAWYCHHx9X
zVAg/IDto85CmNiUPMe15EKp76D9BsH9vMCpvPYV8aXPFY6if5oVyxESiRpugQQ6
NEv1z0SkehBtcyTu46e++ZjH2Z4laE7/Xn0Uolr5wxIiLO8qjtaaaeqPGQLgJ9r7
oZl8QtJ9prLMdxbyUVvyMktEoZmz4ZBsWMsRCso8qAH1Z6Q/P1nj+6agTQTaesxE
kyDiyaiJEMXmPI62NNfkWSFB/qKbC1Nzuthm0JU0nLlMEQRBnBbAH3CZHh6GnfSj
pQwEBSUrsCrQgbkUUVHJc3mgHiPZwLj3SJBLqc2RHeAv4B2TNCHAjTGP9udjS16V
ZBlgElf311joI9/LeE6cFNJ9ibOsOLlfzPX+ZAz+aYEoJjhy0fyZShl+I8b3VDYt
veIeqFD3Ab9yNAi2qap47UVCLiZB6LNxl20vodVMG33hUb0PgSoGN+k6Q5GlqjKt
6l8tkNpKLqD6dNW5V/eZinDOVizwBaK8EiIhX5o7GUAMTlbXfx/vtCkrsePIDBMD
VS8crKmAVd4+RrY3MzUv9spxm88g/ovgT89+E4WsIJ/xC9FQQdRwuWddGtk3rzG+
1aBA5rCL9/t2o148svWVIMBMc6/h/Mpe0Zv4QQRtyGqRl86/zBd8ZK5EH5FcnJUc
lj9MkomwKaoP1SINQHfsqiDtk5x5SNKsxs5IkdFqTRk+MguQuup0oqhfy+/c27uc
EDtYKJL0eudDpvoMhIyTCr9Mq0HVgKUU4BCoGWuBIA3Zbrwh43VB4uArQ636UJLW
+v72rUWR0vxCzXfHQqYSfX4x7wZ3Cto3sICIXt6Ml0BEoJ47IS3i8T8cxsiO2rNI
ByT36arZhhvu+iq8Y5tmWFCNOrZTpRZ2h2/dfVMXEXHH9trpjvjr7gy2wJRc7RPs
CMpkhhbwIte0qn+YW08v33b7knFOp4w7IK78BUAmsc8XMSlmwRb077bTsNektPY/
hRnMfPWaHKzQC7ekaG23OP4H0LB6JmBuWIOv9kF/Fy+a9KcE8qFXf9OyjXqBcxpd
pmEVgz1/EpzagesRkIrnQTveqk4MuCD3Hl2q9tbJ0CrKh9JdFhYYc8R3Sgs90gk4
JIRIGrpk9NiLIZJ5E841wxckOflwSJQM9QVtq5qSN8U63ziNw0ihxY+PZh0rXAjg
6TbPHWjJQ7dZBcUV+AJ8qn4zZ+LbxGf/2GU4gmK+IFAqUT4wmFYVHwdVm3KgdZLS
6ZmKo+eEDNsjGHCk5ke/6mbfNpclwCcO+WsEDyDrc6qcIg8s/fdXT+LE4iYorwE8
Cxfqx4PlT/qvVo5ZOrgk6oT6zDfhVPYh+qwRvRGUEz/YIfjG1Cy8uuWLSbucr1UH
kBWvQGpPz7a1lXru+HNDatwyKD8/BAxRrT3YS9grHqkhEymgAGdxEv/jz+kClBYA
LjxSdIFTRndrG4lPHH89AVrb9peLGD1qWaW0P+nDdfsJdsKFuzBKoBtxS7QO5JaJ
2lQR5dcdFkGts2e+LGWMgo4M2eXwMUoIb1nQXRv5qqOF+bACAe721TsMPgTBAYWV
eOvcpZwUvDvN37DixTD7cFAX56TUAqpNg6KWQmVIIWeLKCAYI3sAWyBMABdrrEQK
UwrKIawbKNr4XL/87Hj14oYG/NLPfNEdM42kTrp2xkxghVGR9ZAHfIcanE8l7L90
+Y3OcDwlDabg+K7d0F7RgOXkeNxtbGX/qRhVuiyhFz0kPATY7MLvDBJ1HOO7spEq
KYS0sbBIbnyr5YyhCG2DBeEPV6NKpF/bhUFiuz6HNGaPp5JFzaZa7I2hMwxOvUza
l63Nww8rGWsD0xu/WkIxvoO0ACyhiVoJQqoukXdK35vEAiTY+A0Js7swT1Zp7DmD
ezcBX4+P9U53qrz03E6Mi0fYJIbKYmWBVDiQ1YR5MSVC3IzJI+UFa5wymBeMM4Mt
Wz8PfDJxKqM2UeX4pkxejtz+9mq0wwwIXgaTMSOaW8AeYU2LDD1NBkwITer3jDUo
opf/yMcdHGDrdFzn5RbN2u3ZQjhQmS0GhZwXe9zRKO58VLdAVROJ8NbaQIfYC1sR
Of7xhUM8R4D29X/1I9odMiKnTp6fkMF+fdaOgS5cSf3ZxtiHueUd97Vxc/XjBi6n
9F13+784OfczFN/Mlb4yNybmJhGHHi6xjdki9YIKqG/SBuk7/Osl0sOn4Aqmmz8T
+LTK+f98bwAZDyizxeHNKEgpCqQZbv6pmQnO7DQAOjdmq85dOj2pw+fu2OfkpaOt
5JO/cF+xKDx2tiIcBdBPqVV7oO5gJruzmWsiCC9SYTL2TAJpeh6/LF7HARQEEVFz
AOJhVDmsjea5FJsO1GkUkEmwjeaZIANuTBWG4Jel1/7xghWrJ+9VTap73QHo5/cC
5qPtOxh26s4D9r3xHA6ZMpP/tSYh6Tvn1bPog6KyVYukiNh8As3GkqsUOlBoYHkH
qxJ6RqKFOPPyaFu5q7bmTE9b1yZZrQsEZAYsFpjdwVtLKKmQgU6R6S1wncFWvGCX
o6FHYhtOxEmBcT2zdjaY5qozPbGHpnFx8/XLsSTQjnpCAQ1iz5MI/FbnYmw4tM3a
7RGLYUAjtgEtbeTWyd1mm9LnYSGWjIcgByRMt0zpMmDrjWr8zBG34CKpGefh5K0M
0KVpyiJXj4KkT6Rrb1SRs6IAWTiM2ZhuNuIoPcS9QBFak7JdvuZ98v7Hd6jHb807
OLHpj66fXKEDHNK3sLvSEnsUmhK50vSMDJscIOUhXUJcH1Llp25J0sV76q/7a1lh
a46/hFb9cXTObyJVpAKvFpN0GgECjn8wSJpV1zFCoUrPCjlGSCgejD3DX4TFoPC0
Z7Xq5aRsm2i7/qKHQBS7+5SABgdmiX9+hWJouQ5zpPqgR2N69eEeSAkP7l/UaI6D
cg48r20EF5n3nhHOvNskCDf5R0h1XS3JtxT+ajjVAX0D22ZgjXKU5OmzDaRC5Zwn
pBFnosCNSBimigbXADPE/UXbEJYoZX1voeY3AfmUrImf9P87Cz15P7rD8NPJgePn
hpkl1QR2shQt8DqcGeTX+OWaVBx5ExzFPd78KcgOV2gQkAv+jBPYOK6/hYmSbwAZ
1NxO4qid91HIGrFE9+dtXqoUGgbkcaizPXsbUpNisEPjJ/30g7OZZYJ3eAcF79ZK
d5weKki64x4OkW8hVUBg9FXE4sahu+GCDP617TIId3TS3rrmhAN8N7LrNI8baf2L
16T7udtS/kipYKXyv8OxoLSfkgendjCji9RbOOrZM6RCU8MOE6fxqPXAU/WOYr3I
Z/jLwJsn+0rW13pXdtyhIOABIB9wgcBrrGOQHVoISlf1H//ov4RYHSDZI4OLyTlH
r9vvhdjEKuR+ytRqmVpQ84K3Q3RQvXXFSdL2BmmXjlIkL5ei+ppeekNMS4dm/E3t
xHSnCS38jj61VFTsMgY2IPtIK0tQub8QXh7N93JyqEjBi5QnqTmKKzKoss1GpXEs
2/yXUBe5PpTnD1dBEQUGzSgyDDRBIw0JGUNaaYYH23lO2fy3pacIk/uQ0cw1cdWs
sHHgNNNOWwEzvlx2fyV+lTif3BNG+y2wBtGKErz8eVmkrj8fxXezIH7CYRR74zpN
CSrhiZXAHHafYgpXFeZ5dfqxDVExsGogXSMMms6/DhGNUJXm4OxZQnjMaPhrE+lQ
uUxnnms+MA3AUK7qGPUf/SAQ0mCmKik/eCP55r9r/vUUS1ykRWPISG7Ziyp6Ntc+
0WtWMQPdBAFlXH6DUvDvPsccThPLDIrj6nm6j/Cob3vjx5HMAspwSEsrGXjjb4Jc
mLBfmjLIBerhrJURH8NzyOrOP6sf1O9w6UzHcKJ2eS18BAz3YtH/+atvAH8b/Yn4
MpbqBUE0BN7GzLlgnHigU6OdOS9dkY+rXkqzauPMnJRnIcjO32gimjxqy73MsKLF
TVHMFaqHgUB3BW1S/JyEULpquLzvuuxQ6t28KIQvy198jvLcC6hfM1fILsAakF/2
wpN24TPXEiKv/xxjZcsCaF8izaOXXLvm+U6JAWFC6LEY0Rl4PUN7oRbllBRxTc/6
Bf8P5yLPq1ugHNs0Kg0aenKHd5UCdUOxtpgxMxB7gJhw2U6TF7g3ZZ753TYX2x5v
ApinjUTT5CE8Rwjiy5E94nvb4N3hzR5o8Xz/Qb5t0O+35mXN/U4N810zbLT5HEln
ZhFc72/1Q2j9fziHKaxZSWXMIyih/zHhiFtTVAQqerttzK9vtxkZOt3H0c673cXV
B5aWxN9jPRQoBHbnrGNpRr8p+xYl3bNWxLKrdSYGGR/QvpE71FHHokTx5nchA2gR
5EtIEiZs6gL9KgXvTj3OxcGwgZHppWmhUv2LXLhIQ1G9BpTyty7ccdMlq6KLHiai
+Z1GCqR14ZpeDgT4bNcxuC2idZfVAAxcMSibpwOHmSDW1vDfmmTqh38T9TK1iP4C
mg7H19Q9KHH/rdb+5mliKCZOpsOJINa4aSjXUbYZ/Q5gkJqc4VFjfOZqhQOFNLG4
i97H8hMhpyNbE2MKD5VZ1eEs8Gm74kU+jAz2pUJG/YXRR3FLQ1jJh4mL//eEJl87
R6hoh0CvEtZzByJxyItDPW2NrZAb5ucMA3rEg5F3GGaamK0glrPAXF25ScxfZA2t
HapQJFiblBZY54h3YuNasa+6tXtJ0QIb/k4V6LZglmrDvyZr2XpMEHqv4EtGBmgZ
gsH5KdmZxbb4WKNIR2rWRaLpmiQRAgS0W0MNwIRIc0HxwfuJk8cXeVtgR+RoWXcl
M8LWfP1eDmyjMAkCmq718IT34Llgdg3/Cucb/ZV37FzgHjA4tL18jbkI7JIyZWzP
1h4+fGOLZeBXEFKyoZGM7+XKMw4C/Qj6tFZMCGFBfI5nx6Sm2FneLpiETk/4IcQB
zHq5O0+RYYsm9MXOFPfud/aLfEW4RZHCAnaKSgaDmxsME+s3WvKY3rhmFeMFWoEB
M9XAuJ2eM5GXQoxqamWUo2qxeV0i0Iq++5jctqJSIQ4AezE/fxxyW2h6GRR9eKsU
MIsoUW4nT64rEPhxXAlbfhwV/y2mARdfhYG2WjXY46XR6bEbgmW6FKBxj+gcveRK
oU4p0X4mzhpCZfK17sy4eSdngGdGChpHGIyhFy+o87qhmpdjAhlt2MdXuJCaloCX
HxT1j6itRODQ/7Fb6SXJePWurCmZy2l4YiyvDLzaCyc4dAZnlvYfusJxKIp9n2Kn
UqbKAGhZviKMyhgoIdZROcSn/p4cbcUuUBK5TqfiK8ab8iVk5vJrawgPihl+vMj+
ZX99HW86kh6FaDV5MmMNAFVYSNNf/Dy+MzjfGdd+32Zpc9QwydhLAytY6nzju6dF
F9O33dt/VeO0T24FvZak8Ym5Dm85unb1rAsCtKhUCnzQ7Zprw7531O4Omkb5v8iJ
ZkB0KbuMtg+UP5fCWg/FJqAINZb6orYwCK5ILG6JkRgpwmnX6zf/NCKEsNGZbz5s
fZcLzrelSFvKGX7gMHPbmrzswEzaiADr+3zWJXl/ja+WA3fWkCjhqkxar7zZrMT4
LqB+Hw2jYTrkvaJIr1DL/7ZIQiXJo9dxw1VRDzGyZdtj3OpGVWurV2qah8AwDoTX
2Q4Ojl6tF0pT7FAQA0TMD8q0Y1D46UkTKqPNZqAuePBVSoZjyijW/vf5qobmSFiC
JcCso1VLkxGi1JVUhpiokB+/zqY0mTn7cVEsE0o+mbFNMNikVYRylKKYv4VZgYhm
nCT1AiFdxS7ZW2Y/JBBsf3Fwf/m4w2FhBPWrtbsDUupKoi/GoDr+XJhj0lLmKan1
pQggo/cCjParlBvfX087IZpy95LOOCsfu8mQ60GznYz/B79zIEph1SIT7eaakOjH
fOWRwBpTVQYx3BkzQMmyHabZBmzNubW/buPYG+HhMWZuZgxb4ApWjjaLweIN30Ls
0a0j6FBkTsepGRam9Qs3BvaZeBfNI0PthT67y/AmwsRkHMYA9gUwBbqRGzfUh36Q
XXwLnL353uBupEEebqhYHU4mXDUEyMt95ex/Mz7cL+yGxy53YzerEiTn9sxxEaI8
YVDDszIS7Qz4Nfk/7v7iidmDeHEmQPocvJRkerD5ukmj1fz38XE764B0KMg+pkao
lmd+N9qTtzRZAv9AXMk+cgUmrdMoSoZLhh3/DWg3rb5W354PpBVIJcQTXYQuLy92
4kOgoW/SZUdRdP7WXcSx5rdyPFa5G2qcznLKYSzq8/fAq8g9F7AvJGRI/yW7Eron
I6r/+liu+wWtfjXJ4vsuRWrml9ugxJ9o5RT+4Lw9usrRLjKTorZtq0fjcTh5akiH
GYak/O+fVGuscRDdsTpFJu/TgjxUDcZi8DeSHYQx2bCIwKdewAGA5QbU+ef9xvTK
EeUV/AfHusfMSaMUeYNZXOqug3U2kKe4y1F+uzhWs+yeBCU4v4YXS8lkTUnmNpBq
IW9oudFqDaKdBEKUIeoFjIpCSFrcUW/F813lBfEWkIETwKN07NIdbMXBOKvimOmM
vYPP0+EHltu8slE21d3gjC5dhq0DglIed4sTMAIxj8LgHykJtVg73u/R+Hrp47vZ
CIWVlRyF0xltAZe6hE9hEfCFvtmNADCUMPbuYu1vECz/1bqazkWc0aQfKlQY1f0o
ljP6BEyg+L58L7it2rTFF4CAK/N/mF+ta2Ue1fxYMZKQNIu6t7WGd3c9J21s99Ab
hnW1oIHl5ZsJgRzlwji09aj/9ihUP0shqoa03Va5xwXro+6Yt3KO8HkTwgzDqbSv
jG3aREsUXkJmaqu7Nv0Rw+Ccvma1Aaaazp8CscyT7YKElGN8n3UNkyMz7siNeTZy
z0ATN7YNiKdeDWLx39fYjhdInt6RbHNw8bC/5rXsc1RIgXK4pVI14RWb1nkdRMu+
L+T9Hn/lAG2B3msRUeFKupDYtWdUyJSZfaqrrkY4JUWDKmXcgMzGDEqGIA8kZ4SF
EbZBEwi7+N8ibztE95WiRGDR8cQ2lN5XjbQImUDx05BMaAFDLdBB7T8s8s4twu5D
Q+5mab/1TEpEI/B1QFQH4J6fGlCVmXfm8jlJ7Fztp9bPCQjzHIu5/uEHcAI38jcr
eiJn1Twl4QanFKStThsVVkCfdHg1n49k1ktCdKUiOaOlpVTyizE23JN0sMLwttf5
YKtvhnaOFqS9v2BW+EUomfqHNzXg0gKGLOhPWVAenjjDDxSRHAM1N54EKGTTI+LD
OgNdLA/0U7Ahb4RsdA56BBmmI2KqIdK/o2jzyfRGhNuY2rUSsXGb9//O9xSVunQS
tfjYAzufkx0CwF6rdIc4ZJfIeL471Wkyj9GpFnxjMO3T46anZldogf8e/hm5JoFf
MJaePTgPOsyAynhoKOYX7sx5gN0GYa2+IG1qHHZPbAsjFy1spD3JPsHGSSMjKVNm
ZZEan05JM91crFNjLZwSr3zZjQXPyjfYXXHoThNzYb4cLLIh4MXZzpIOwkyLptgM
EvfF1y4GVB7gXaoC43rft1OXqPTjrhv53K48SpAZBcS1H5sxP4daBeVP3LL96gbF
LC4M/PfO5+SnPrAwSa8whoQ8tz3lZoqV28Qzu8WQWCw9POBMb+KUsgHLelsgkF2w
e7k3RBksXuDzBpuMifwk6Dm5T3g+yn6SPHEqrLyaJsfJgeaMjoL137wNppCZidrN
jWRQqOafM7SacbUJN0y/cOHP9pTB3lJGDFWe5g7WK5Fyt4ICuFBwCIAYuH4WUgKq
7z6qWyI80kogXdnrP+rPSmg89y4hPvW1KUYncpqgQJsv9dN3MntKcQkwdJKLnkh8
+k39LAw2qLo8wAN4MZQF/QVb99rvWfxpCSAuQb9Q+ESh3d9jUPeTheke4xi9cguB
YX1xRELL/gjaTiYVEenUYfnSSLiNaVOASRhzRRIrP61JB02JvzWkL/Jd4gcGSzkC
fao2cbMYO4JZaubhOdd9QCUUQaTiSHUD8ZQwxofD2yEFL5zBTSRcO6220zgRuhnC
L5nHNn5s7AGn4ztZzkdD/hh9aGpcCv9Y9l4UFSyAPB9tREUxwwQb2kBGj+hCOB+p
VENRrH36bLjGQnFIS+fbopQt3PmpEm5CIw7g2y3xCfFoflGcHl+px0KGwa/HDesW
lYcmRNgg9W8ZzA8aEDEHNZfKn6DyAj6Ht84R1rWzd59Su74Haq64D7tnBBbT0Lo8
9AWPHm8K4ptwUOzKde65gtzpSmZgAdRCk8r5/bTx3XSp1ojbeHflusTLym5Y5p0u
znrdR0ISh5jLHfn2sxCDqCCVb4vJ0psEkaaYS2Ls4WiRTw895KgjVCV5U9KNo5LU
Ozzgtnca1RR8FppidUgqutZ6ssHIX/NryxCv7QcvCz9A1oR6euyxzh5nooDdXRKj
gN19j6261vt5RVulnVYX+XzA4+9RAGlfju/p2ba5y/Xr/rBK5k31EM0knfHKgdY1
0PeBFRT0JwArBYEkVUr2J1+UQKHu0EjH0ojtGToHsd6JYYtc+E765RapbNdUIHFg
kUaCzjM/ry6IAitAnQUgK3BIMiNAu9bIbqSOXl86/M/5Bn90kw1t62agO0SIKuQg
evOpg5TNIqm5qtH0jcudBUKhFrsSr5Ib/oJVdTs1V1ZgAb5HrUkbECxpFs21OI81
SM+uzDMBN+mg3DlzhoEIMyCrvZdjABRCLioPkUYgwTfkhzFSNvQP7mSlUf7jA278
oZQYk1e44yrwArmJVzZpSiwl5XwkgJ7v3Ny0xB2aEntCAJE3LjtEZRSYTDiI/tr7
RDYMOXMSVmjO+4QyRH5YWXXDoWIwQxbFlWaFJ8hSMnsaYgq1wE2gocjvxrHgUA9L
WCdzVNcv5QS8zhn/trLqncU8REQzrtoAd1ZOfCkrMRkigSquLC4sSN1B41+1a469
XbWsDCVI23aHAyxMk7CHjhy7FTW1TS2GjvLzEztGtms1qkndHU/qINQt8xg6zgJ3
LydiTBF8bNVrv2jY/2nrDYkUxz/hydmaott/I+ATt6JyKDmZ85TCmoMIxCnKHi9s
rVs1+GQ4OOAA0sL0WXFNxDUqgMTwJ6Aujtzn9ANGXUWEK7+JKouU6EO+vTOkAiwi
EEnUYps0CRsW2UTphYl10Gkx7ujJjIl4HoNHOBCIPPkAZndy9Jda+92DB0mNywfE
6nu1gRuaklTMP3FLVDmQYbEA7rCm9+piavyptc21IsXDvNMdBWoHmpEjvioO8IcG
zEtfHKrkssB4jc/s3kPi0cbKsofE7wdULlAlwkvpx4apcPoD1EFIDCprutCUGQIm
KNGoo+fzWNsCRGZ4EfN7mPNgE2U5DJjysHFzgQRKn4kxQ6WRdJAg6yCkxMgvm7g/
6zQq2lLHzXvPlLFfGi3ptjpU7lu80rJiqrQxPJirdBQCpsjFR+yxhGJmsl7is1/n
x1Q/6rZjSRGYQCq3CvX7wkUTgS1GGjvTdzRLiRHa2+IcLRnj2QIDjFVmBuvcegRe
pSdhTJz0L1wdKI88CkeUyY0xmCxdkI/UbGmq2ORJZfIrcNSLfLDHW47ftwRYrzcI
L18ZaOcSxtkZLkbjjknjZPfQTuX440FO2/lMLflNpsW4VT+wvnePk7sbll7MqmGL
AfCBeGDq6b0ZGBlib5XOx0337/WFsjoElqrZRi4QVRpg3COy2dE1VlTRsyjGek3z
LMd7CV/4G1Cg6pUm2iz6rtmEYmLXD35TkQAbJi6tR6YxvnEtrgh8ZNiYYAXE12SJ
WZqFNcSk9kAtM1JLLyb4VNVQite4JMwoUurtbfCxXzzs0n+e+6se1waLd3LB4n42
oFrHjzyY5ao/8ZMnJj6jIDXN01JfHs4seTxxB4qZzf4Qi6t3eQDHGKIQ7gU9PAhm
bkDdwiV34eP+pebrbKDpnbA07e4JlU+sw72E+0sIKbTrVz668jJCxbZFFP9tBUin
rIeQXfItOkHi5cDCcwpGHMsogRFRUTPHpRfgf8y917CPyZUjpiPnGGJNh+UZn97Q
2X8Sl+ALUp6zWFM+GUkQpfxDWXBLOdseBrClTUCpTzLgL71Gd8iW1koD9KG+5OC7
F9LC1Bq1ORjdCzOhk56bpYAZRPaLeVEChR//A82mYnts8pNalYorbI+77fGV6YI7
scT0KWupuhERu/MbfORFSHrGOC+iSP/UBIkmD4GAbbGQMJqmt3/NrczSaQfYIAdg
8LC2cAPgSBraf1e/RhpHAVyPdt1rvOQRHb6KAMU6mibwarSdJbI3njrEdVZV8/Jk
4srJf9f9EqWo/oCThUQCMVaF9BN+sL5dddrPM13G7jShabZs6pUDgWhAFZCvSzP8
iON1h+xfLG9EK/BPzcmpB/OToAiewl1KQDWA744J9eIHm4V4WqlPqq1HZUHUpkkg
exTWG1ppeGhQVqZxPhz8G3VvyH3hrhCAHCnWlwTCJzIN0P/jgHRdDsHsbOIoV0WM
YMtig8wd7tzG8DV+Ye4g1ROB/pDsDf770ZH6y7eqNQYXP8ieoUHXa5iFlTeDuZJl
sPF9dZwP0FBADWybMAlAzVFaO6m8rALbV7nOkPHB1dYvpFUyJBgv/PaseruvjkFs
cOcnUOAtGObqBmL6sQBu6NtxRC22ere78P+4VkBvw4EeWxuXrNhvUX8UKmiw72bM
k4v1XD155zV5yTLoS51fonYCWnl7dQxd7230NNWS/XbBbBlOoJQCERLIs6he0uza
E308caeJFn6w7Mix7WGr0fRZ4ApWawwyQAzAacb2O6y8COuq3mTr+ynHleRUFBoc
Oc+BJ4cUSWU6DlpLTbddhn80VBhsAfBNl4qIwTDA9BQuxXyDTSS6+pC9a87541PR
lb/xK1s4VZShnUXjcsjWtE1g/96vxWnLZLK98P9HzuvDSRC+Va4UUeA217owm3Y/
a1tyhOcYMteZzEWkJNBFCc4HTa/8y0QSNOY/oFjPT9serVATZHcSBYeL7juZJtIE
vr5vj48IieOVblnVq04RsbeYpoQVQPEEnbEeSeAlAbX1Pq1mBxQ48HEtUooXEPvZ
9TYu7ApAbfdXfZvOSvANruzub1MTKFZW0mYbRMvuvBlLFJ2PjsPMbCOx8zaSyxwJ
00deK51kT9uBJwEzsGaRaD/Pri98U0FSnVqM2JgajGYODCL8TS8hrhUOKFxe59O8
C5oFmpt6emOTItYTuLCoEWXhGJuBOfoYwv7NyTOWF+/dCuNFmB6/x5fTUuADUYuV
5XU5asLmS9TAxI2MZ2kVanl7jRSYbNnfGKeZC17BK2ptWohjKhgvrnZx/t5mxL0X
gmBhW1tmEONKwCmpMW74kVBSaDMEQwJiwNog3ERacmf8uekqxCqJPFBVVuwYZXqm
SDKZrlbTZODFtReZebrZcIumC+2RwVbS1jw8UjTx266Qe3Dwn5ie0xgWSdBZA6t0
miteoitbXWP3LK3UCrk2rCkJTZQgKPFxQ9xmBoO30j0PBtt6lEOe4BNrm3vbl9ca
359iKuzvesIrvaHCy86FadJsgzAfE20LITj8FFNGe3IQdVaZakgzkC+TbINDIHPN
GcVf6r8cbjlwAn/E4K8eh3mMum5N2wAADm/gXX74vUbo1YKx8IMmtXBa4WpBAUFG
d5lQDl7O0psOyhY5GMZqTtC5QWbD3LcoTHeQlGGOqpY3KP4v8GwyhZMxINrPn3wV
EKWlv3bTwJUt8CMRpCLf/O5dcJpsLyaW3WP77sXfuxPc7bixJqHdkcHFRLGjXzDr
g9nXEFoG/ysWrHRArFZqp1k1bEtNbBF4bo0lLguyVqwJuTtO6Q28PcfZvbx12nxu
T9sPUK7qJD4OntBakwSKsmdmDuTc+7tjfwi9hF2akJQFVXWnVKgbA/W4Q2f4IfkI
uPzBntNg2CRzjTQ3ELB+QpFArHi58Ci+8+vebAn5PAKkOxSgB6a2RP+RxevIIeoD
BCgUWHLvmU5V0S8Wh05/K/qSXLXuM2ug2Nu0jssIzCWNxoBH1x3GaTuP2D4Jbd/y
iaFrgeEuBF06IcD1vEGEkkXtvheNTj8zPsxl0ho/dQywcgUUJTiOdlrl14RuzT+d
9WEFVdlwObS614+nFvxq1cDxc9SWiOID8MQsL6d5LdIJuyFkmNi8rd9voFvw/JWC
QGKbAcYVTh/uV6Jy4uLbTIOZ4/XWZyXeeQNMFrbldTp8UU4Uhdvy8fYgSH+4TepN
7jbvOpivubNiu5my9swErY8Du9DuBI61NcAmH5EuCYqSmELxUu7Lqjn1wAn0K4xm
EDrb+VvOt6RKc2I9UXqgQy0W++h1cTvOA7SC8iSefvyERCiB3iAZSCr1Ms7kB0BJ
5SZPK6pgPWB77VvEKfZ7o9+EcY8cVFjM/fi1Kv1EgJrFFqtuHMHgcmR1VmPAESF4
Sxe+5p41nnEPJ8zWpsKHPVEXyPvl/CdeHhAbePKmlrx+MlPmoK817bhkPdt4+iay
ZctVH7h5eEmQFcI9PqowCT+kGHFGNffEu9jCuXsBOuYgzvmeOOEoXQsyuwn9AYdh
M9UGF9nQxoJhZEZgd5QjOooaGfVYs58YwLqcp74F1bzpfxsW/jCWlGjxo+arQZGS
TwRrB4FP0MkKTkqO1TGoN3XwsBrYa9ck9bmCNvwyesHK+nzWvvu4yE4y+orbhnpY
EY77oTocul68pTSObOmoKOzAT8KMKfiM6vZKNmkzhbTDKVQ8WVgiEF6H3R9dxRYw
4A1skcHcTYT7nAOi89YUbcPBT94nXHr4cPTgDBlj+ypY8+MqxTyVx14/w2twijOe
obpT5CU3hYrBVVPJ5sXuiEzcIGkG8jwqmW7+VR7Ak8Y+X8at75jcY77hSAxTa9SC
3URaI7zbBoSwzAmXZDH0e/Ye4DP9l5PAI4g/764++m/Gw609OP3xxewvlounKNfr
n4IvJdR+/62dHVUQDtrFPXy/7bV+m8HwMBXFVUm/ykh/SR2a4cXNwUxhvsBDMw1g
robctT3r7z+obhxz1t90n44qRe8vht6Cm/tghQTb/mrsJZpS8B7PMYJu7UCKZbAy
cHzewX8pdHO7cc53NRxxqtNt1EeLG6z7TxtUYsbc2EMZic1ZRQYJQfEdJnJH/eP6
7j2Ce/l2+1E0UfUswPuD10IubXjuJf2r+a1ghZF8r19dW4LOsUbK2x6z/POcXBqX
Z8N58qu4tConnZHC2183bKh68eHLXMCskHd8kTxpuxTgp/DeH0sqsd2H5VBpAZqS
zz6mXf6WF3O75UxtGys/XaAQoIB3B2v0df5yuf5RoCTv5Zj0FC5n0OJdYAt+fwj7
Cxj1pta8kqZP8/UJ9bvTCSLrfXzwGdfex34RkKPocJD3lGL2JYds5JarJGZUep6v
mAotVqsaAn9EHKt5nAerkoZlFH1uYLvguZTdRNFisv8XxlCcDTHx0nyJQb0vQwNi
nF0OEM4ah5yqGokVMgtKxxBb5+iOpX0RBsw22P9eu2U2eglcyQGt+oBAyVmRUCMp
zZxEuPscQMRjBD9Zc+99I55x+rwEO3W8KxRxISAiieAXqttd0cUJ722Hmn/HraqR
90F6veICpNRtUWbsjjfySIS4Bsh2b/CPy134iRJ1ODe5V2B9rpCQvrOKHqMAqKGu
o+TAM0WSRBqVGBFqlNkPKXVHqZrqfzgx4NQE7jmIuAkxlGqc1LlpWah2VCfRDt4d
rYxKwcPdcFEvc5eRL/CpEkzz+3FE//Ah+Bc7B16qNk1wrlj6nk6U9zVnQbm5joXN
ZcwSvyk584dDCTuGEpOydGAaNvRCd57+thqRd62rhfkW2MNv2s33pgWwVEXmUvHK
J7H7qrgLMzKNvIJgDUsgonw9pcE0MIVfAD4hQJIj4X4TJM7f7e4YtTPSkjpTSzF2
XtcgaEVSBjz8LK+8pJFFijiEggZIhLgSg0gT4UHKFY1p9DLAZJvReBv1d0yGdOJr
Ijyme7RRA39SW/g2Bd1TfHuyVsmRNF10fbn2Xl02hBncrkciwSclmSW5sscwPe88
J8aLptOt7XxCQFeHCctBlV8pyVshF9bOr4Vv9CM++IjQuEk0HEly1+SigZRQ19ct
3GWVx1DDyW/+rGwXY5MCmPxzaGShw4aqCZVD1uZy4pS7/aohs0I9RaBG6G7PP/DT
DG7+/sfGOE3q5wRb3yu/rII9Fv9im1MyNkKn1090GEzHD6fRAZpa144HBhysiyDl
TwIZbSGAfKgjoCwZYOJfAJ3JxzV7HprewcHs6uOHmEkqt3x6f+HwIFLJYxMLUwTh
E4uh31kCMohGVZgmqzd9pNhLoLGMLN7xxcGuWKxjhQwZ6vjSVbQNSC4YezbDZCZ5
J3c7IoiPTybrzj4LjQrSeR5gYDIqUOLqLeQTfFUgS46LZ/umwsqPi+MLHnF8PPQL
P4fl40wBXdx6b456f5luguqgdYfABQEaMS9ur9S6ltemJI9lOLOmXgIaZV/cRR9z
9ml22a8VI7FfyW8tDivQQzvUBQtDbPxmejBceXeaUqbTimH7adB8Ss63KRPdJlat
oEpUWpY/Zing9AZe1a6VvSjWfE+sT179ei26H+Q2KslWQjsDFendCuQQzrsVuTXA
5gyQs+WeJJ59yh2Szr+xAlz0r2JCxY8isfubCkhGLnrr2RDMJjwyxNH8jtOTqXTt
mx8HCyIr14Um95OGnzo7WFOofFnN1nAzW8aALnyN9OKskmPRfd0CtMbo96ihkAHn
KoRLqmRVSEnKyxjo1ZmRjAmcP8m8sG1oUnH3xQQ1lCMoASZxhozKxH3GiHkvRtlY
vZDsWtdQyPzgzg2d0emffstcpq0K9pP0KGxmdhLzRYDCY9N/ZBm0XsgpcNT5QUHF
FyBDFEKNuDqw3kUGtNZbXx6SVsC1Wcd1pW+SHE58r/22bGUIbAHKRPoNt13TXFKY
P18/p6rsCsk6ZD0fT9yBdtnrLWgO9WPUC/1QkoTL+XPYcXbpYd4cStZgmAq4aOuN
UBE68Ydabonu05010PZTYTq1f7Qa5br1BgbkAWN1Y9mC0oripcKcFglhsWu6kuN5
sZNfhGrJ/MiF7rm7WgMO+fwz+2YWxg5NWMFGe/pVPB8lInrSNbG9eDmpRbLdpSsK
4KS1sHD1M2xhDWuoWP9wMClNEVQ4Fo+djWMkY24jY2DKNYOs5NHEGu15ywycbrOW
WOPj2iUo3ArIplQKaxHEJkNakxUAgzT/8HE/JZgOgHZDqVHayvNjuPTnuMSaFFEA
iRfU6p3qPCvtJEinJE2BmFAezYVD2mTByjitA3ILz/SMQ9/BJrOs/lD3Uli/QccI
9SPHuoCWoAD6HxjIUEERhLl3tct0TmDrKAsc2Jn/G2XWJZ1ex9fJD+CmYwqa7JVA
M2YZt0dByfd5bLYt7ALvhxB5rl0G78N9q8hTIMLcO8FCCErDfysJuo6n3X9omxEy
1Ha0euMBnE6D6mo5Uoqw3nt2tDjQorEkjymTqwTn+N1HsxjIghv6Pmci7nk/FN93
K0/FITfecPvrRgrD4QEFhiQPqhYRdTG/pKBCNwQjdeBJeiA/gB0IJrpD+v5uaJK6
PYqvRwqKZQA02c+6ENRlPaAW5P4t1MRb/dwOmwy+nZcQE21RpxdNo0s6oyLe5Gzq
DAeXhr6qI+Vf+3mQMfj11OEM7xtYvKiGvwZNRAKBCOlGLB6xrfHbTtjY6x3IsUBB
WzrBzB22dwFGQjKSc3/HyfzsIDOd/DzgETLhiqz4Hu7+GCNwbrtBOiwzzIe1kfDI
iSO1n2lCDgJ1r4wjRqIuufUzqAUzE+v1rUmAo1+U2lbCI7fQyQHz5hgWq0bqsFNO
NDlqdev0Da8iMIJnzOjcuJIzCeE6wW7f4+Rmx6oUYi2HXY/WFhs94aR5ICe32Ym/
BjQjJjFFWcPuN5HA1fTYEcaux6X4yPkwW66Umnh+UTacW8XQHS3Lp2OXiSiUKcQV
bXfpEtbo9PFPQxXzVjrVoyoTl2yNcWPgho/9fMQtuGmYGoVcp2cNQw6qIwMvckVN
17zg23+GnArxbv6K+69lE6rTdfc5JGLAdfiP6UVBmz4NDZAExxHbBkKSHZS3tp7u
keD9uVU6yzk2FjI5+4Es1W1Aw0XYLTXj0/QRtjJ/dhvSOQzwR79shIosQ4qZnYpB
9EjqIHlpAI3Sm0pLUZkJD6DfoBCvUdr8Ym6R9ekCvwc94DtwVc5RJtI7b2Yg7Ym5
rauBneN8zTKSTSc58M1dz/qptLOfbcTXTrbcZ4B6oNzGKTonH/AcmIlPboOmp5/W
aWT4MXXHgTSjQnP9I4afODOJ3MGj3406D3ZzWoXtFJz24GXxhqnU6bTt1GucxcMa
cipt8ydbioNBDx1V+3a6HAlijmd3G7ED6MKlRPbTdNkZgCqBM+iYPh3bX6ffSCxf
7Ixj3nycGHWSifKhtgiyxkl4GL36SVQsPIqf32BXup5NtsP0qye5DdFQgZ35b1Ha
PHjzvWYzjsw7D7W2cQ6RPgIEEfcAWv3pRuxCUvg2G+29THwToSBLqHEQ/kBJIfTo
EMbphg/WRSIkzwYbLyvotcLqaPT/plIAsdbX/NKAziY/rZ30CgZJIXBdSnhb5oNy
GRD/r4SdQdYSTn5j406HtClSRmHh9MeEInPEMa0m5LOZ3bLt9PVLa4JG8JuqtiXZ
H6ZW9hZBqpdtfwagMudj8L1nRtMwd6b0FuKZYMQo5qpK8rxVgFDE+lNyqgYV3hNZ
AtEOZCkzT3djyS+epr3FXgi2yDyzK3dxRBMMX41xisN/3Cjd6hY12mJ32zNRSrA5
rlmVGweIRecFT8sElaiZTzb89zWCnf5G/v1bEOEQzp17/qko08bRGXttCYVSoAhU
TKKorINqe78Xmw/vBpgSPH948+S0WYFEsSFQ/sdbuRiQWB9BiEJVpQWfC9lzcrR7
tFeJsVvfSnqVUbwP8bZcEFtWDbYRbNajHE49q5TbrDIy5pzVvqCZY0NTclbPiH2+
+ZMfWGYlE1b9i6DpFVKi5zHbFGnSeewa2IVm+i3QK/fKnoAc902Oug0wZ+zB7a2l
vsytwaBC8zLbOrI2FaZEoI13FjMymqy3PKVGdjuppqi5ZqHhRLGC/GwBYMgW0gJV
gWmWBunZdpFo0DBTvfYx2aNEK1bCnVkyCfJ5LZTtIwC/4yF1c4h0sBk9Z2q8vQJm
947AMnRQDdJFkPPSBt2H3ReJzQ9d1DCCEgVEnKHjLMFaDJ6VjAaStfsjWkCBBOnn
0YRDBrH6TG4OO/q4B7gs+5q87kgTXFSZotK1tVssljyzVwv4jZQ7CLTtUPyRsGdz
Xh8OiybtSP6ZNXNB9AyUjP2fSBQRwYzizUkpmYXuHZfipBcChsSGvZmFIbBHPMh1
W9cuyXpa9TRGVrxSgiDqkZzTFzidgLL5QDVOE3+ZHL0SqDUpzlBKu+mOpk8/FUUZ
AR8PgqWJYRDJdqZ/OFBoL9shXaYwqSOcgKTPBJA8lGFu2UH43nPuGCacYMmMTksR
vx+NIqP7iEINx8BZ29kNEtUFl0y6ZpC3JP6f2qjvqvogg9gcRF6atPIf+oI/2aa7
Iv58DYhaCP6APZMPWMIis5VYR+Gpxm9kIvO7PqFQFFMzy93PkZUwVu9ZFXHmMRIE
QbNMuRi5QPf+SFXAQkrO7USI1NgyAel2XSWvMZZzIY0ueJc6ZR9/U7uVtiTcErC+
OJ/cpK6uyifJBncvCrgC0MzsCbBKh8WN1IhH4rdV80tV8z2CV0SQjvhqmF5CfLrs
ngjEokj66cI2l0iRMLqtOM/Zmow4rRhMjGSDKDzsN2OUfdAOLZLH51hCI52UMepZ
EwBt9XCHHmwPrWlroHdSdAFA/zIwRCWmWQsDhdyfy786y4ZeAIm228M6XAfD9qly
67ta6iki5UkI0D7j67784Cgj9HtZLYArwEcn9p6eZnPeH4/4OWu1lQB4NbSemiXX
Olr5mfdmItCES2Q9jxHu17hYJl3JoAZ4m+WRLcUz0dQYBaEYc2edAyl92yAm5AIS
+gD2uEvHje/9rwnTmll40qAlN6Fu5bAFCd4giqLvnHqFV0egW3/OlM9WGjuMEZNu
W+jJLRqtWMANjVLibvwv3DhhTX6THEHkHt+J/yPkhC4s94IJD+chN0AddV8lHfUy
RinvcgS9Kd7kYtPJ/tZKGQA343nxa39zwCavYbJ3Ji2cwZ8jdjZ7e24ZRpjhFe7w
KtsXRxK92dDwZTLhOsGWp1SMU66N+mOn6P7Ks9L03EqrsoQI+0f0+Eb579OlSwKU
5OJBkawkzkW/dYiIc0IFI0kvS41vL680OjxbSXFa0mOH6yBC8KHFzKFXdgwx6K8t
MO8N3xSq8zOkE3ABYW4RDVimgXMPB1dttW74YxdKzOr3qF0a5w03dixCviszy9Xf
MCDq7+Ko04GsAtNbkTm3ElINOto5ppmLoaLnbspz0tCWT5LqzkjCUPzWJ6mDnMcO
gQKleJjFLXCI0mdtcQXcbeO590OeyAK7F6NWRoT4cYRI9vZE/AY57HaL67lREEDh
1BNxkMT3NAHtcFXOVcSRcQrjViErDK7s7sVKK1ay7k+4vNm7JINbOhOYbFXOZQBP
dKgo/8jnuC8kkZePfe76tZ4lWWnP7C84SFba+pUeqETxwhZL/pvWfoJ2E3+fMKDC
UZANB4lq218aC0ajbG/WfhEUZssutF3DhEod/fGGZnO6wHAiI5cW0PKW8xvbxBta
4/527DL6Rysl2NQEg1kIX7ETvBpWhu329nZnn414n5skOcbYbO1HGbPZ104ELZ8f
bHYJwcLJK12q8m0hyvxng4xrDc+YO40fvLkIGq84CzPsiqDcmeNjGeL6/GwKfYSN
NPu9L0g2zeBLDCIsBmKCFC3vazXLXO3AxXguJawZceJ+/FS6Hndi/AdP3PT/+OQm
zKyxy5DkZ+3cjksM+HgmwYDx1F9B3DEhEEhs7Qf1drY7DZfwvYI+4AgMnbZKEPv4
PqDzt8SfQZ9TVpqW1sfxi6Mdo7NabXiJ6wsxnPj8IwIlyolUx1Yu3N5Tnd/uid/7
S10NF7TK0QrndoAjvYBp+zM3AI36fst3bimslaucyoGt3Yul/cM8CWse4LLSCm/t
zNz+T6U9mJ4iXiMdl9G3ehGE+pl6Ht2cB3CCJsKVPiZeexE40DfecxDZqnzDERq3
zJeqYbZqvGGkBMgTfW91k4IPbKI59BsMr7q9D1oY2n0zspChrG2eKFjJPOYkceja
sXQm3Jp3479QOKjUyt9Ur7FGJpDaJIRIDaBhymBTn/S7jIcmjS6T2BrDYBpyb4uw
ADaQ1MUFR2MdfMf50wELRJDK3hTHIise2kiJ34tqf3+twfgsfTVUl2IXkPxW63uK
0WAKlYyUdY/rs5+vxftSMFCAyH2KlacdecZfqHrlITumVrXr2Qo6VMfy4sLSIIAp
R2sv/s4aafAvAvux8ZCE/qWCOPLy7ymQ7g7x1tfdweOk14veirvNP9/eItsWXTDO
Y4s7qe1adl6oXTtSrg3o9Umtdp8oh0mgRBv8RraVlToad/XCqQej9X8KKh54jPcR
7aOoARO9ytlc1tT0Bp8BGBssWvKmWvM6mVcHPSbswgyozM7QwUVAilMtfrOGPh8Z
wvv7lbVHNTZSD9kHr5Xp/djNgJ5o9iYQNKl+KDLewGNoJD8/Xyv8p46M8JA+m/yi
CJRFJy5+ZWmZM/kebez+1Olp/bjx+BsyMMl7g9tPmCTwR3cAQTkkOn0O6E86NjnR
mK70eYksKfSvYSynXg8cjiQUGdzZcoT8m72r9Ka1A6PoTMqaAVYuGlIN+K2MkOqm
fhg2Kgub9oeqr52+pkq9aafcPDBqL2oHHOaO0WqCKqUGSSWYOjnIgB6eABGVzTxD
z2F4SUtmz3lfef8rjHb6wKRERtSqxbgh8P6y1+MRYUx9534WdYRlKvD0qBlD+Ny8
JFsCdJ3gBI0tpAjl+M828c7KF/l3thXbwSswJ8v5f+2NxZ6GoJ4bUFmFTMqwR5ff
paTkBWb2Ny35oR6iBrT1aWJMWP2kEtujySGE9JTIgM64Vap3BRA9lZn0nQCIE5vY
g69x6iSW5DzNToRyGpZYOWsq/juf4wcQFrRAVMxAZQLZYmQSq+V2tlYzydRdAhOl
5AD4ZTF414mA9r30eNr/1otkVPmUi4VCM36/aAcf4AUCXllQsAKOWTP5P/WAw1kK
OxwadI7DjUT67yoxLej7BSBMNTHTKBU1h/Kbqbny8Kaa0WuPZyrHZKJXzZVCtf+d
iMzKtHuDqV76lPTK0oQEYIdcYS0hTUkn4nWEpiVfnl7QHQlg0OvrkU6Nj6a0IIHC
b0KzTuK2hlmSje1C+Md0HOMSeizkMhnxJrjLMTUn2TamKAzweQWpMHi2O4dWjtpw
mpV78iaP85huTIPkWyWNZqnVq9aPb1G7JnMSt6hc+9HATCCopw2MSEpNb1HHnHND
RESIBDEgQNa/lNaDNUqWX0+xRBxuOnjAS58UK1Pc9Z5YCArIUKrw/0Iq+xb22Xrh
96zddf1BnjP6N9gcyNWATxTqvG6FKdn/scCXMu4Bcz+aNPa6740eKJndVaa+/gQU
YWtPUoRWp4gSuWJcYOV/ib97asXV7wEt1WAglqMmX/3NKBfjxjh915yd37b8HBGj
SJ2GIoI/MO+DJvdIi0t4GLsTYoDfephA8d4BISn4sAun8CmoNylqhJoiHeyEFAGo
M5ZT2lzCaUhIwJyjk84QS0F/cJFUt/qbiKX5xn20TfG8S/nVl7FMZhrvxmKYV4CK
yveAVSgX0wsn+IVkiTG6mwNg6AqyCsntXDRrRB7uOs6bf801ncPK94T0+zUBDpgq
9QH9QkeoDWp/xRIECeW7PB0R5gRyh8opfxpzoSXAUUl04hmwAIF/ATGmN/Zjvw4N
g/YXC9Lr9ApysphrHocm751SuwwMyFjlNJJMjiQDp6Q+JiedOMHLQrK1+zVC8MPz
oySx2lDgTuQzx69nkNRNDtJgAaoaKSY0Mtv9jIntnzI1qxW1GiUf5uUM7OV59sxH
Z0wY5r0ptQIXDEgic7pwu0rEUJZs6RdIULG6N2TqWayy4Z1ktGqywY2EKeSCQfCb
s/G9UK6I3ZeOmRCFGQF1CXWPbISdYzm+LYDBVwbO6XyrB+28CKjW1sh0ACDUcBDP
EiHn9bmeJ3KFkr8wCqBPQ6uGjllm0yn/f1f4mtQ5npnGJXdzLa4Lb1eP3hgqx+b2
orJXaIi1/FhFaNs6mDFrA6e9FSZFeDJeFUytiarIumQ2c5toxGEA+qTFr6eWl9zQ
U4Gi8UieXJ8CetAjqreZrWHns3c8T8Ogz2I11NFUgmqqJJUrmdW7vYDabU+X3wDa
gUJLRFwezMz51Pm9Z4gqBIHtRQY9zCAz5XZpGKatgQj/+4r6WEVi7BAJ2BXI4Btf
pBO+q0h4GL9GOXeP/WYtvRvSe+GocBNdv7sgxn7H+5v+9sZCbBkvLXN72S25AHI2
uaFyvkxBpY0bwwdMl216YVd0J3Srn0qiVCxxCGT3MVEl/wE4CW/q/xxrqKPweYiu
xA+B5XGUqDtT2czQYLuCwB8paXrbRHit3pDG/G+ofCRi6ZJDqFxJyORXUo+VgRXE
imA3APfHfzqhhEOcgMLhJ8W7HcUZkPm3Cdz9g2h/KpCh3NsvCzFNHV9VJmzxBuq1
wLvoTNonuKX1W6nm1C7Ke+bUYWV2ndF4rF9vHm6fUteglS4yXoaiOczqo42IxXTf
A1r2vaeg7aBvIduqqp1FqkKJz9IMSG+i3LSHQUcNZX01o11FLxR646fj5nke2E1T
a01X+L9D0XfSDf7SJW81GxyM1L2HCcyVYm1itUYSPcx5TjWZiRswZREbD9/Kxum7
OI359qzVNiv8n79iQ3ib7+q/YFAl+kqPl5T2H/FMdv61kjMt7IZMJx0NAGaLqpSS
pGtiA5gP7/HJ3qe/q3qL6nrYgAzO4kYwt00TIXIQrPYgcl6rnfFYo27Y7HmSXueq
gbHAyGzOszBFi3iFW9sv3/Era9x0FCZyyBOAqxfZxQ91cNJhmDzWdAkS/m4FcJCN
9JC0oxJQNkbK/HYZCB4RM9cUAtL0fFnV71EmKwT+a9DiiN5cY9OShh5q+PYfZ86r
9cbgI9a+U30cB1eU1/s2ec2ycBhlpFf/JAGoYDHGkQIIxexq6wQTvwez857mJwYH
WdQgWMVvc/OviuWAw9S8joSLSUrq0Lx1Bq3Jju1cIcYw57j/MpeUINfdwCbvHSAK
E335Y9dDng7Sy9AWd488mM/AJUJLjgkTTvijt0/hekf63EBLjxsBeQc7MCNAO94l
6QlmtC1CLAqZP3r+7WY5NtcHosnxV0+zqekck5byQG5IgGtm962Zl+xkDvwcBAV9
xWxv19RJcFlTGyI5gtOW/7FPkjPrT+39OnjAxI3Zen/Nr9HMx1RIgem1JQJfvso7
rwRG4rW0MET1PIEPM2+/vkJCuFpbvpfABay0EIwW8IZPytUj9Qo13x01nYwB0LrK
NveWVCt4CzNYQsGB3mpblRUqqtEVcwRvLLNQrVvo3g6vc9E1ozj1ww99/jZ0XvBL
6AUz35S8HuKBTHrwlhmZXcbhrsen3tEzElv0Py1RV5eZLF4jIT9XJu09uNcJaHSJ
dpHI/oP4Egft3FkIQ/uDdPuSVVjt6a7kNCik2E5ZUdxr4y5GoTPf15HE6txXAjbD
TTCRAnLgnmtU2wXPPwjqsBZljQVni88xj99GWAadPxvohnp8DAByYv7Q5me3dmRv
XN1ryIXNdwNYMbRzndtPduYoo/4ycWeHOs7Xc+puuojR9Vdkm4upHYC3HXOmrGrV
iLJrIgPHtpMrCh2/QaJMq0ufGkSkYsTwhkQub9pKMJan9EFovEzazK9up6+ccDNN
CA2N2QLYDXC1mchys9GfwWVXlwfD3h4i9oVOMfUskzqHwIs9tuCl1CjgEJDAyMOu
YvOU4NG1zGo0sSG9BuHf6YyLv/fUkm4eSVbSA9Id+/rF4vLqB/YXqPw/yxtNfWQK
/x7kbAHeFolsNpk2zP5JWGTUm5Kala4uNrjSdzizh/LChkrC9BP7T0K4qWYRPrsh
RzocZWA61SqCfnlpqBMW8nfbJOFG0RZgslTpWaBc9PsnJFIToNlJw7qhZhNe3PZ1
MSTHvxwwjuKd3Tdw8oxFn27yztDyI8yK1ReKVALT1Mp/+UIUpGikkYAWQC4NW8iv
zV/atdmmBs18Mtr70mjNJdmLTnaTSpSEZ43GHhLWy/gzJ3It1Bh5JVcxJ1k7GFJf
JRZm+E1EtgOD+82DRAyAQuyd+F+9aHzeZUkxKyaL9IJ7BhrM963QgB0sjeO9+sse
QbE2w0olVrs0SwS2oxrd9wJ1/gjXB1ZzN/bsSbBXeN7eP6RVNq9Hujx9lL859rS+
lLmSGD4PATn9UjZAP6pjDuQc44qo8GApIEc2cioiv5X7x5Bm0CFOAiKw9stbJWGh
NQ4zUXjnBvjLa+kGpF34COyrqqpb5ZQH+ITvfmhrNA8IFYN/BX9MapQLzAv3D0GF
dvrPV3T1ssQ+BAss/K4g1No2MgC8RV9rAP66uvqYwbCwKgkLc5zAnFpqY3OfoEhi
O6RgzdJF7sgBL6Uj4cHxRqUKFRnVQZtaQfnelYjs2IdF1mJSevUDOd2uJ7Whnbis
adb82YnvWwbbUGAzP5Jq4Fp0hXUYnL5o84qyiiRladla3ckKjPdApvXR2z0PY9zX
LqRkU2yZqlg58p7FX0jZfX8oI3y1waSc3QJqzob/1SAr0kYapRSlRqdheJGfwf+S
FYwcfPWpFqDzTNhrHm0F6hS8OHvp4XYa67k42jmuiDqk57yMtd+hVSciYACp7O+h
znpa0JhnY71OjQpbBkwFSOLURPtXQ5O2hohaND8qBCr8eh3wi4t7sBe3OsLxoo78
qgbMVt6w3kXyT7u36zV+EPMSjKJGMvTtfSbxAFAc+Fnb3K5mWVeRU4k1Q1gSC8cn
6e4ypjTdc3oDlm50E+/0nKA64gSLasyGB18BOfFruDpGemCybh8IodqBe6I/dv6t
DdEvzPp2ti+IsFmLhn8DcnSqj3OkSW35g+34N4f3sc524A0OyCjYk4loV26WdJ9r
Vqi8IW85MUUXziNW5DwKRF0iD+gcUGT+i/CRYcnbsSt5TiLsWntjVuE5P2lDXwN0
FktdXheCq5JvRRMcMAOimJPhcRiJz/pqIEJJiFXAYuTfrRxO4+QRVe9HD/JQ9HV1
GVObj8XuUuMgW1GQ3RcvlQtjY9DF96uD1INTc0B1dKbS3c1FyC8aaUCj5XJeiwGg
WFtVqUOXczrlg8GnPloXeNDfs8uSgdz3ZV13PPHKMCpOFwTGK0SzNFs2i442tTU4
vumRuKlrhKv/ntNsSukqc3UEMynS5GkpXtLTpl6Mil1orH4DguHO+1WgqdCTrCEs
KDlOAN2Yyr1zByF35/vYDAUhBAoa9K6Tj1sM+lDTViej7kmKhJUiUOFzxWRFjfbx
KpxkQiXuUIU/kPkltC8m4rEl1G+QQW+XPOdjGWuwqLd5mYKLmysja/6BwVgvazCt
on6UGW9RAdzMPVFYN4ZWXO4uif2eP3eiZcIq2Y9etEbajluggiyce/i4TGvskKlI
UITWMO7nFUbkjHre/xvQM7HetrNPSunbp2tra2+6+/NL8J6L1gJ10eVKYN0E2V0D
JQNCuiqXecRFChpFR9ofPztOmh2SUeRg86TkZumzTrZxs6FT9sQjNUCsuPTm4mR2
tQ9sClsGvRV+AzAMzzuQR1tQTu1CtK+rdjjqrcnpJkxkLf1m/UT2Xw532nAkzgt/
ETSeXJz+SJa3C4JVn4kECKbkFwozNuUK+4sQGurskR+7mTPhGOEEa0360NoAz8p/
+9OCrls7AYkcn+2USJZyjll8L/er/qctXEBiaklbLHuQyYYt1vW9pR5WPOnetVLo
GMP2C144bg7QoP479g0w9RaSjY+a3l6v8Uys4GwbPeffvnV04Mf9mrQ5KApQYQny
uLnDcyYu6zF8radoE+FmYIztuHRBJbavwG4em5ynxTj/R4UE4q/1kl2OuaPaA1c9
wccq0op8Ku2l/9AvTXKSPpoInmIaqU7vyMVt7WWgqLHK7OyfxxyxT1ZncVvC+0dL
Ei33I1dRVAyS8vffLlwUk1NoslRun/X0r6270jTrxCVbQRyFY/7BwwMI4D67Kxs7
i05oCHS5g1+w/0FftsGG0PrbLCGPUFoAiwkh8I8VN00tiDS56G+yC2Q6Fb247k93
BgxWQ1DBaaUHH66aq4CNgzNyimyU4qpfZUBpMCkvWiuzA0fCX/xPTRPjhvnryNIx
aAXpL8mrBpwB3bLNiccWLF2y+djOP3FXITi+o3J0Qx+kNDI/+TiWdpyQ3JrpYBdY
o6bub1/7MCOJ1W/KJKMJ41G1FJWsN4Glmst5Rz2hQfKYQ7GxGwzp/3SFvtoBU5aK
+JgOYCcoZBJGoqqbYB7Bw/tP6FACJ2b5f4vHRm81SFLtJiaiNHvUQT7bh29+CY79
bmkSh7RQ7wnT38V44gDFEWAHyqX9qb5APiVsqntMB3lZreZCckXO60CJRAJFbrJ3
3AqRoi64TT1THjJJqqsbQ+/N5xL382ny4tqWk1+48aCq43marzLRPLm4YD5r+uDV
7xxilU/jj+qF446ChB6SKqJVjsv/TZXvrpI47Z4pTYRVevmLeus/ZNeTH4eDcNOA
GM2sdgwwKBYaxOAMoYyhRedhoCEbSkAtIzjA4rSsZBCV8+eRCY/XdXIULw3K/wOm
CvQWnjeuInJjL0+LBPuTFyXsFRPfUimKcErs3/U/b0kVBPmqRvygkvXgJkPJpn6o
kYpmDsDzax1N/0vFq0FGFidynTics72BPFjoUD7wTFqqEQCKJG+V9FfJYvJmjJLV
XmemOKSx/o4Y1PAP/lsLoklUrRzqxU70qYqQ+EyZffzI9I1FAWbxL4qhnBszeUuI
yu2oQzR3Po6QQn5L4g69L99FUYy+J0L2Guk2+EGt5Ok1zpG1TGs77y/4MLND1y0/
og7z7VUWzfJ1Yl3EZUXZPwYOnMu8/UE41FQjfVdo+ZHeZYiv56xY8PlR0BwMzUg5
jS3F61a4aKGWxn5Lh4lzkmckpFDI6aaGsb4IPoRS94+fd1vEjVzGuVtzU9OKgmnI
oSWRQu47ZisPBta1qvRHWpiH+HfUakai9SFRIYtqrA2f6Ffa2EtZQ/dOnyc/pcua
khsZEUALNUzhyHU/RDjqUCaQamqQlgphQmb1GRKLFvmTpv/bgW1vwsdJ50RD7R3q
/Nj+t+4FddE2a5oz2WDf3ykgS//8H8MYBsBh9o365koS8XZiD/C4dVoOn2EccqGt
z8IHPLA69V0CbOlIF3MFbha4FTmQr85t3AMEl5UtzHKvbH6FVvfCA6gvH9LywKDL
irOeZoXJMArrCsYMOgiU1NL3DLXitEBgql9fqeVb4OFsETZd5FGVRqHQRVbH2JqU
cD5sXr2dnnk0DR74LJ2pxJCsfcsGTBff4jaZ7/eaFkDX7cj3uof9A2i1sgnQTG7T
nx69UDF5qDElLFio/K+TuPTmtvaQyll24Xf+hF2Pk6sZaPkSKVDGKAzsip8xgR+i
NUvqVgLDQboo4Spx3KPeRxdos3Cbl0F2AZu3msLiof+fBWo2l8QEldd15h+/m7ji
kqWBNQ5PC3L330rYs1cljjDCq6Ky9zNRs7CLLvbrfjWJrTEje+deWODv/LItSGb3
fZIEWe8h3AVli7YZHNkaYmwpY0GjqwYtlGvGSYDVJy4fJ6nuheaXN/UrL2SFMVyZ
ytXmvCj2yjMigKJuET/GmO+UryOhbe+q+JVmjZV84kk9jPCpy/jSnMpBZx7KMnfb
aYkYNKwAFZKqLZPANGDhW3JIW9pp0KOIziExB/qlwojUEcv2R3SINoDE5b6T171v
RAdElqihfgw0ImQik4QdRP/4BmXiSurHgcik/sKRuP+LpPIkRvZ+K7ivX512sFPW
6ytwSS9pWfTTEca4oUWUYRGt91iAnDixjV6GE5hUOoz3FP0ChPOINyXp6k9gvkMg
0oFV996YpHHc2ATirMsYZGKJPpSxPEK6+jjOY7T0+1TM1br2SHoPMJI2Uy011uwo
Jqxa7Hb7wEWb9p4wBy1ia0/yJOjq3iIcbcNR95/Ir21EisUKVGEvhVgfmL1tKTJh
pTdZYjtAsep4m2mFve3o7VahTU+z4RGhgdeU7NJBCJ5CQZ0n7k4A5WGD79XJKMMa
NqnZjK+aR9a6YerR9lp3hupHG+qm1mlEFSeAphXxYTKZhbvplNtD7uErkoAjD3NS
hrJ7L4+j9EK+fsbDT1Sa+4tDE0se/lZ0HC6cRfP/q8JZD8ftYmflsnr5w+BuP9Mo
EYxj3/yCYTt0xEAVbbUgWoRL6PExu3kDevSzvCnHmCTlSc1KKENcDesvtasEevRn
zq+ou6x0GhCfyaNo7B4ay3+YeRy7HCobU9UpmILhHH0yswFPvzGIbEvA+cipZzul
vC0pzi2nSbIQQaBBslpAu97F407WU5uXU1Ekh9QK8L9ivLQX624ViadZDQIT2jlN
OGv90dYBQaYpMTvTt+fu5uAVrCYYLSQ6X7CZzfxP3Mn2uQAwnvCoLL2dQ834Hlp+
o3C8flIsxL7rn2+p6ke9uKqNOdAdF0MfJFq8PtfzQwDfJRl3wUP5jh7Fjqiecq/m
sOv7CNZqpRSsbZe6VNbObah5tZ80qyd8XcbTOKlotN2wDZFp7ZCRlsZkYKpsVxmU
stXOlHh8WjDn1/ab9M/2Zy3OOlOH9PNIb/VZ2SlMGysn++23UHcOqgLRW+RwtMnx
941jeZLZq1bJQhTJr3kdKnn5x2GIiKmd911M6dSsBdIhZALxmIQYsgwH+oXV+S6j
Ng5v9uQ53RrtBHziyiGpbnXCXJs/OYLldatuMAEW0lO7h/v9qsdibwiTJyxtuCmD
SbjLjJzkniN54JWbf0JxXn1tpvml1e4qGzMErkApdeI4ReL84KpQqFn2KCj/GfR8
hpJxV5vSw/ZwL/uSSzD53ljUfWqAgtX/co6dsqwf/YrT5hPq+PI+HykBtZhPDGBj
hBTD8ueNFruNyB2wl1xn9jpJUdVpczQlWWqP+Ub/U6g/Uu8MogRLGpdZB/DTQ0ku
K8RxqRe91VMv8iJZrpsqM30DqWqW98DiHXRyxKaMisljmFlMU+K0X/04RIqc7K7c
7w8lNwlJNkDvXYE6f9Jc6HKY+KfVumJzfUX1HLpH6s/LReNoCwHg5sg5QF0Son8i
f5m0kwoV8Hqdqw+/5fWFs0xajFTVw6k2oGc8szOwucXzxzNavPfU0ayGUr7ROEuT
qJfi9gXJJkYtMh5L3b32n+KclAprMVXE/ifLCSeJSmxbxKTeve6XCCs8jVp/k3zs
BQOZvzT+EPz4TP4oHP5XefKxGgD9yBNIFfs/cui0AXYeKaY10A1SIb16OtYloJVz
ZIOEToX0hcIoLTDdDHsZUI2ZTiRELImndyh6cU00iaQbYDntgsLZk6t2ECOKjuhd
xZ+EuwpgeupaPiMuMbi+cQXz+6sGJ9gWXDISrP1gijkXzcPgJK7MUZsZ2NfPtlCo
5lgfF5NOwXobSEl9dH4lK4P3HtJI7k5pvej6LUt3pExgm8/VrzFHY582hjvD13Cc
EizswDbVoX8jzAMYKcYP14J2YJdIF3tGrcXhLs0WOYFZ6PweKjzhEQWmBh88Syfg
I3zxK8Uow/T8MRe1lfn/iWHcm8yyFv/PKV2Zuu/RgLye1EV5v+E69ZARw07VLx9S
Kwb5TFNvhy/XobFcPjqHFvqUPHf3f6BHYGSEYtI4oLi2nhPDdtZDqL5ZI9JyPjQt
KksyaItb8gND0vA/Ujc7bKMDCLoU+KWZhcghGFQUccB7iqaXqGND80WWWA5r3TJL
CBCysi2DZPuu9/Fn1pCk3WBob9zWVBbX6tMywOEXYzGmNa2jHO220V1dYOTGzhyK
qJJuaMllGDUwzGWADLQW5a9EDgs5sHrO+UO444kF3sfueLXtSwTM7pm98SxQUUfj
E2N00ExOkWFYSgygVFChfb6l1fSF14ERYx6jUjVm1J4Q+nkc1alzbGJzTedq+mRp
oDzMSLeyk7ebXfhIF0+Tv/eKpAM+C7+T4COw/9YKChjoJOGGO8A6/08/pt4kQ2zQ
6R4Jzh2GtycGIzjIprM1Jid+Km4T9s+K6VdRlKxwchjxjl1mZ8aXp2cK312ZtS85
Fkt2U+V+QARk4/5aQInolOuUNWTsw1eaUUl85VUAd/nIC4/9RGXq2+eOq4sR53M3
nXREzkpvUFeQ2Z1QkhOafqPkndGgrZduAosLZTxDvnT70s7xrR3195Moaber9gI2
eDuwYLQRAHQoGKDQjypv49v8d3kOpZEk8PMMDrn2UiOaicjvbbu35d4Dq1t/hRPh
muv+WzLXe/Or4bY//MIMuNiH5u/WOg0cM/TYQXlMMTrDD1F/1QxOqSKBBjO9SSQx
Zkbs/ElD1Db/ypr+OZAznOacK/6h2UVd75ypv/PuzOF6dfnnaaPf6FcHGl7WMLaw
44Ubx4z+NarlV5bxZBqgdUs3XioqKc+V/sKcc/iHmxmmfJs9c4azWSrDEwdN/PDN
jUn0FIkJgeHDXhTmcYcAecAUXLFiE9V6Xah0z29aOrJd/+U/Vf2Sa2k+qKYzID9N
DpERuPZGHM+lFs7M0BMcXNO7y9Qd/A5uXovRlRFC/UHBtI/aQrmkQdOy+UfxeWzj
bSkFa9Asc5PD+p0JXfnVq9ewmi/ZovYOuQDP5mOWRAmxkk1FnKwEVP0fw0G+wr+x
tG1wTT4yrumJm7s185aWx1Qf9HHCyfungpwie0l3WYjia20QGBkGXJBh8PUIutFO
H3rIdt800v82okzeUdpjs8c6prHOp1iF+rO9lMOXDr7AfJC99Equ8e8mpsZ0I+lJ
6yLoLhKKk+EcI1gU+tnFSaIqGCKd6+q1iUIEJll7NiPi6JqThXKwP71TVx0OH+qT
ZvDZr5F98AhG7pq02izdSkgfglKLoSR9akCCVCw9paGl82KVFiM7F6cpqzL/j19t
oZ2m9k2OdAjN354US0jmGxc3BcgA4KbNWNNbvo/EZSnNF/TogAzrmA7Ja6JUx4Pk
uXLNkTkV/1sgJTTskG05gOqva/K7Dn0KkbxXrA2k1OmpIwJ6o64AIwJssUHzU3OL
bYb747UkYbS9hkSy9jGM3J2Yt4NBnWBYI+wwq+AtfB5BnFcLlpo06/smGGYhiMio
aVwCa+KmpR1CKabpi8qqVzTQtt48o/fw6r2Iou5RNjYy1/6S62ybRSwmDrhUnpTN
NGGFHZJKMRDjn+s0satMfox6r+BZZwclKyyUhjQtSui7VKMRFS8NSL95cDIHlXjc
XcQFmRhyLpsK6Rxg1v+4rueXHIZ/P6d06zlN0wNTV90G7WahOHDHjSnzFOO9w7y+
asPyKgODd2PXyIe08Iml9aklaLGCb+8VexqyAygADKOC6AAAXpOBUcl4pzKbC0w0
Pi2TneaqObWEtr64XqzbLV1qXZGy2B/5THzcbU72/ZGnYTmeXJXffdDiNuFy5yPq
kVmZsRamFFvUACO8Qvp8zC8CsflS7zrZGVGRaQgT6fhVoguEF6URxoWhIr1jVYoa
QLkVL1cCmGbRMgrTL6DdvSW8mwScqthuji46Rya+jQ514FRF4lRo3gaHbLDPQuvD
KUFYCGI2MZ+qX/3K2zoFqBSdHvDf2U1HGnVy94Y/lr301VzEwKexhd+k+/yGo9aI
yaDG3eRus1Cf/kWFT5CjY8mpRQgBmIt+rMfDmQYvZUOk/lZLUqyrKRS5WO0oIR2i
or24F/qOLuodWLqPYP4bM56fMkg4CxBlgU3ZQeq/Gv1YxYQJnk1Ps8v8jeAoot0G
sy5kBBRoqFogHmw6vgrZ0GeQ4v3kMldCTO4YlaeX6lOiNlAr3FcuCwexjpMxSyEz
vJBmgH9UFwO++/wdSDMxTRBCEY0E7HovBjudExh6kvLV9s3Loujml7N3Mx6ovFDU
vLIjOCLQp+TbNAJ9wUzt8zEdSoG55osDEfiYxz/a5gUS9fILxzqcWbIg70Tv/Db8
Q+wNILTsDbNp15rJYFFLVzxw0kB+hzJCyxyeQtJ040shpQyq4GcuTLzhBD1pddvV
lJRjIX0yFuHGMjmWFhRD0h3B5bkOmLTshhmPw/NSGivVSdb5ECWncZrvjTU1QPTs
ef4K4fSsLN3Z0z10HJyLu8tJH3t4CTROyJXXYPXbylFF+igJHk2NcE8ARUom6axH
bms/XzalAn12Qc2P7aTxW3wBUloTEF4DBMU1tpdemmYj6PT68rgff2mHbcm/PETN
cf8iCggr/ExzNg3LhPNbQ9ckhGQRadcB05lq4KCEJlh86S1lPZGbrMEq6FWH7dxb
VX8C1vCK2x+G7rlEXC9AKnfSF2WKtWyQOy2jf5z8I8qkpvBNTcK3eGbJUz6OqWCF
HQuy2+4Vvb2Dvy0IlPU5N40S2gpne6C0QrIquJoaaVzjZQizIJx97I4aanoZA3kP
gENULWn7QeIbkUM6ZXL3CwoIRhWqNzhsRnlr5qENYvJ2dklyzaCOi3Jw/KQhmVLv
kvCBtumHlo+2RjmKEyV+gKN8yaZ6kSxOVuUOJjCyfsccz5WzVye1Imxxj9Z4fVdA
2FJQnECfC96fAHrXZxk18yAKzslCgFY0piiUK0xSCtJTnwJ8yrpoD+cqeYz/tSrR
GqnebqmVTPMLnE5a9CauoD1EeYB8wfDCQ/UD4mj+asF1TjvKOH9IVF3r0Dkyo2DJ
G0sRBrU2nKXcn4AuFy9gjVQ5epQ2OWwxbI8RjGICEwpSzqWw5aYRwJZu55NJIV3H
mgz9zFM/kL6uF07L+iJPZ5mpJt4BwajddZNLeKmQWBm7AIwydJrL0sDTCWiYa/T2
9wLvvTy03uSMtIH2CYR7R36OLJF/VQnb/sdHDWxZZu+mpHMPBSXP/IYCsd1ElAVR
yr27MU/5w3CgZ6Bl2ZXHjYjMeKtY/HBJavytTKX8WhN81fiacqPGH55NUzZos4oW
FtOwLq93B7tEoO8vgqqv9lqnv7aFWvloKfVEoTDQ9ELR+kfNRyumtYO+2L+s0JzK
2K6M2/ZWTWozoIM9piRZxqeuiOHAHAtRo64qeEbXyHMVonEJnZfzvsJ10bx9RNUc
rcSjwPLOwiTbZXrrv29IVPPh40hBJn4GUz5UGqLAPPclYZhI8AqNetkL/CCMQD3S
r9XGaRavCp81gCf1flJCntpetNUAyg7hoCKMWRKS/9Z6ucaygOfVuTdSzttK4Wgc
VSFtEE7ibn4weFVm+m8w1g9ADIHkzhDOH8bmpIK26ZywpE8IYxqEBabF540U+f/G
jyGb7xOhC1XGplGt2lDuZuzV9+Vy9eFGiDZIodmqd8Vv1Hg5a284QR4qHu/cAwtG
5jgUs1BlaAAYXlRqGGDiYLahZnut5nJZdBQzbKFxYk5fv8+vJCNkoUoZy8vEEBNI
DVfoPqYA2BNu/mCGKLU56WhmMk0L4fE4n4IYZK52ZEyk++5uGWGKpWiy8/hUv3Sm
VrmDIYEPKBQZbTpmG/jRPsBFCljKfUeJXeIFQgnqNdcPCV9DVH3U2pjByS8KciN/
gvEuyl89ydnJObsaMxypCidk4OYJyLwzjndv3gJtoQ+3oqPdr/w/XRgdd683XzbT
2SHhAjCWJlgsvrmvbrZPve7cd1FMtlANSyBJTEKM7jUCP82lFYRutxcdaNP2ILEY
xVtCAKmtNe/STQWwgHaKIzMRCIDXlBl36QQmAdWpvvQIIHYLpRAmA1R03PFboh2t
247SU7urxD9frhoNd153vx4bBivNB4tklWI2i0DTwM/3kG4AgWDyVtjbPhabyMvV
7yDDB2ilNtYbGyLEr5/8O4cUoTi1mZnt0XkUdyKi9KZslKEe5O+KynYs6DkP1u7x
/y/OsSTmP/PhM5sV3IXtLe8q/gavpgnY71apayGqqC+RxmYNU9rMTcic2nCQc69Q
LAG2kuIQGqknVksONF7h66xSk6eK6ZgjV94L3hgvwK0zE4AX77uNFZsI7TUXy7Fl
zztbc3GnjU4HLqShxYs8nL8BnaoXWXaa6gl6CZ9qUEosgCTvPSL5bAjQNo9Pu5Xz
5yRxVYi1rr1TK4ruyVwaK1gih2WEylAUuWqMMu1by5HkK7L6WwSvj69PiajPIr51
iODtEY7/BE9MVBcrjKjrqmdSTpO3sYoVXhnBGXIi0lkJC6k29NCvqMWGndT/xDeE
5ElONfLWIMJoHtuvxnX9oY/O9VXpWR92FpyItKYpmK+9OsYwqxDrhXCB1DAqGs3a
MG4iC6fe0r0kkal0kIegoKJfPLJvxd10M1ItcswssF255PQri2HCUq0sawTYrFy+
VRi+GdqXmfGDySEM6yThjq/qu/hDyqcEnY6MNbLhfq7JLJV82r91f+C8u13mpqH2
DYUPi5Y87DoAm4Gm43pT152EEbvDlT4Cg600SxI0UZIvLh6DsnqRHQfNHMvYf4aW
tTLz2aviEzBf5ALv7kB0p0LE8ZJ8NG+j4d8V2wDIOBJP8pR038hjeVwgDoE05LqE
sfJX06WAgR8XGbdh1nziD9HXiqy65GnEpO7GiRUkFSmmedEyTXgvEaUpnGmyz98F
l/N2yBf60PFD9L6bncMWklcITYWrehKFsHxpkZFpvVdDT2kCv826DQs5qJzRaRsK
18gsvypkmgt1J6oO9/p6kYyLtLWYw08YoHIJlfNQlhJrPafNSF4qC2lNxE3OTal/
amSD8dqe3qKVGus9IES8wZq8vczQUXsyoYCADRFZtAitPs3waWukoCc7hIjY73Sw
oOcyaONvlyele8pTqk3IzqioicLNqeLNoP+n4lNuXCPqIwlqv3QTcAlozHbHa2UC
JppamKTEKKGzz5+nihcV+Ov0QV6Am7BRhqU25YzbLHchbx62kXun7FzMbiBorphG
r5AKidg5Spmkoxhi3VWpDMfoNa6pou/mhUnA28fgLUKKMhMBjNMWpEk5ZLGmdTh7
PRF3mQSDU/8CMBOBk5tg23izYIEXf1OoLYnfYtLXOLfpBAQXLeVtxpHSTHDafR4U
vHpNaWhbsThZgc/sBVoE1v0yMJrDI91Ofa6rw2tcBuKWu8bNGquggq7EOQ9thiGD
uYdoXD8pIVWHJPZtnB5ltIAe95XgvfvSuGH1kMdlX68PY9NWqZMQ/hscgTYNrPKn
s2CdA8wOm1TYnnyWofBbdD8wKFqDCkfkft34sA+h2zFtzAyJLU/YabJmfC1wp4H6
ShGchvEVybUsmYwN6ArXosNVcVMNoo8460b+lxEGkXlKB3a2qu849kH8FWUPuenc
1QPqlzxZ1a4swzPtO1y0VovIFKeET+oAXKhGyEY4mO+RoZbz+9Wz6YMyEYCwQsNv
UY7aPPqS3YAzUy1xigqCETClQKA3a06kI7NQ08kM0NiMUUPNVe9qvOCNH2dosfbe
mpBs1h1sqD3sSa6RXLWDV2+IG387CqOk014+KqqaAtIub6Fq+Uk/5XH7mCrRSHIs
rX+Zj9dvTDQv6XrVkOOmHezZ3B/C91dNcwDVPbZJ/xmM8uSkdn2bv+QPbRhpb+Xb
iblRqsmwHG9hRVdeF0+tdWRA0D2yfzjF/yMjOHYiG8koaBQqgmBqZNyXgO8FTODE
bS5m+3ZjvdEU1wwmp3eTXnRQqid6B1qXarReP1Y8GIp19Kl9ZmfuvmsDRbYV0M9W
VUO/hDuNRwHEKAa1C2D/pn1nONh4uqOGKPVCw4hEHm1/rrcDDcCzt9Nwg1CM0hNR
MGeJvhzgupgWuRN9AD52FzB5gqEB0yvf3QrZwxG+aCqtpxTZNNAxgY2vwYKoNwjn
NQvsb/9iwoolPGejz+2Lurc1jHYtVPItl9WcRuGh70lPWscnkMONhS1DAkowaRto
lSGuDQe/HBiQk4rjfaYz2WYR5N1STDrZkSUFdNgSgw5J2y1w8IrPMI0p8DWH5Q3+
3kg/mWh82n0Z6G9pFs3AI8Nh+4NSZXMo3ms5thC/E817qNqZWKoqxRgEyoGcfTXG
WqvN+pK+mTxSl67OOwk3iEitfubH0rjG1EA1I/9UQITqaP/g0hd7wasUS1+Z/WMg
FsyPP9FAsewo24FWNSFiOE1JxIHHEQu1VxLdVWbZjc6ne3k13dpf2gJbJvqNZIv6
1uR+hYrpTrnRauy4LZdWCoCTyT/RS5E11yuJ5UjVU31cXkyoMxNyvzNoDidQlCt4
Kd2DH8wC3KBjZpHOeBixPx3wln2BTxMMcXjGqnWtSsbkg96PXdaM1rP2uStob2RW
MKxNC0PbSB/3Q8ZCtf10DvIHtbwvZBVyCSZ68JECdWrGKlxQoEsfDer8MGPh0YP3
lTwa9P7pojWyFYujeOjeAwmQZiRNeb2jrDiFiM/pfkOoZSL2v/UNP9krg/onwiOA
auHmNoy4Hf1vIoU8rZuRXfolHSbOXokUbG7BlhfVtpCBYW91y7wheVgmT+/8t8iu
FKDG+v/py2vO4hFYn+hRY3TLe6pEBSourFxGPOgJoKBo2/RQqwV+8mlLGDiOt5wS
iuxV2hAEweahnOMwNWAx1jaOz5UhsuSZxBPRKtIu0Gn3bLv6pwtCis2dGeae4WfQ
5gpiGcbfRjrsesVhclmSOntRUuxblRAuuT4cvXKSWsVIpBIX27+vL1yFFexSrvHU
Ix/DdJs7rAacPbF1pYdvbSunP4SuXNDHHJmkI5aVn6RFg+HDbeYPFse/FUjZEaX3
7wEjSRn4oc/cjanD41NvPp6saOGa6pTbPyZeLVBn3NAr7iASB/SCFdOFj6GA1Xej
52ir+BQzydKaflO0VqgXPARa/ApP42Qm7fNbJxrcTlgofZQ/0DChIavV5PjJYh2s
83zQXAPyF/VqlZFeafp6QDgPvVP/YjfxEPcWiabXn/18Qd72NBzCfBstQiy0VzZK
nHzg1hZVdwPOtii3/GhANE4cIdc6FGMuLJwHEu3cBYTef59TgtAdHTRQtZl70HVH
0/DWQn8lmYcDs4tYXvu/87hXYXLUbcpXHHK+B4cYsL+FkxIRgJKrUF+wSOs57WJ3
L/ioGxu6zV/trfY9U6HVU66m8K0/Kso2oxG4h9jY8Q8EDYvS6UOfMMEummrcKHxM
TM847SMGoKqrIJjyfBzNNExx2xNxbKAcT+f/rXzEnjmBM0sEhVHeGpiTL72c2brv
rsHgrrjPw6bQga6QCXbhAZUIm16gpPeKIWDXbl1zSx07lvFShjkRnTHUQYkYiwou
HUaX0hO9lO67pmk3GNvLtgHjZ/wYSHO+QFA8SzXMUteRO8aGaaPyRKmnBGH69f0e
hAxGDkdoONrXDS9udJTh1SQGR4xaj0+7OJRrHxNDi3rqIimMOK3Qqy+AlvSt0qmH
rzEUwxeDNL9s7apZQqkPxOIqvKzL0UZs+DzJ4WX0D1DejVS3PPb4sXqoOvejv2la
SZD+OIlvAwc8w6DfmRPBhhroO+SxstoKKhDfO+Z5dRICS4ZkUXEK9Wg79bKanR5d
ZI5K4vtaKcRTcGzbvgbFnq/stsUUegoXfBl7H8McYw0KSb6sAyiASOxoXXk+kO5E
3bLne5w3R8ktcsesRVCPvxSvdxYyl8C+A/IMPP5ZAdldZuXfsLhqXmCbltVTUuhz
oqw2P8iePb/b7Vpvvr5OCYCIkjWVrCZrilGCIx+vjAu1xN0Rfe5iG8VnvbbpGIzl
dV64a1wYTAbC8rB28/ma+Y8guOpDeOihJjR5qXeeujnP7iUERSEalBlvZJRLOj2x
YpuUvTVggrRHj6gYtIRpnlaNkT7D4YdG2oNzLMzcgvpQUbZFl0IPY9wV0sFYgFfD
f9A2oTAKm/sqaFSzZB53BI3sA1wVcdp4aQjkvrpUBDjNmj+7Mtzls+DUQfScxaiE
eu2h7Dkf+BqjrStNUBijvoLz9RxuFHWrnmx5Vop5DOSNmXr435Frylbbo3Tsw4Qb
HCkv7VI3aR4t4Rpm3g3qxBKaJaK0PvZMwaghUpZpmAiUzCtQlQEvLipZvtd0Iv6r
aGx8z3ZXIBtbfyPUVhkT0AHs0/eDuqhBDqH2NXDIAQ7arMpPSTOl/iX11uNzf9yB
6WOPGHkVvLzwtfIfjGGzmS03mVKlEdhJGj1LreZOi/t9FgecUf9EcHIgctQGxnxO
GYaTtu3qwbg20+cj1BM9Cyxtp+b1wUWyFXHcJdnmEXPGaftn6Kg5U3/RpLBZfpi4
ByiriNdMvrpuGMEicB1op/1olMmj/ePIJN6EoAvI3njn8gvShePhO+Qh9VT5KhtT
PkMu02i1vzJ3wY76qX+NFPqw2aImWkRzXWvSdotb9qG52G2RP0FUgHJACw4nTpL/
BzmnMrYR2d2jD3GTvAEY+ehxCKiq5vmYCfdy8ZYnH5XDQ0Ons9NsTyPjm3WRcks1
D8YMVylVqyI4OfEgdaqbfk8hMWxEAtqF1ovgnv9CtSzyD1LkMpCFNP/MnaeoRJI7
VzNdP5NuK2o8UFEJObWU1r5CAVxTNJwzxVoYWZaVYvVXN98xbWzDwQwnMqNnyftx
VBAH0kGhnUltdx9iXjFhZQB0DMNJ/3xYYK//VROE9tAAwyugmLRTK+2Q1NEB2evx
TcyPPwUU2FjVpHZp8bcVa7vrOnMHyXlawUd7zBHSqsZpgK66UvplmGLjcoN+bEne
9ajYlxMOlzHh0Vx1ryr5FPBteLiLxRI4ce7EL2qYIdOdIz23u3+h5MMI9bUj/wW/
P4qQoTlsaZgDJH9EySZPHfz4jrU8SGlxpr4olOSYaRzzcOlhzZzwGa7xD0F83u4p
mWvJ6QpSOhkk/ER3350ANuaIffTAUbD5I8P8jjgjyjykOiz2w1+wRzNECEJhimrK
0+9hBdNZPUiHaGpKJGyEFo8UP8HqRwKAnIpbDc36F9WZ0lw5uSqTt1/RAY4+CZEY
bxuSj3FLcjAjt9pXys9YinEHW7RWyCkn2EF2knOie/wiUzmPV8aiNtPWNRPz2jq0
yf3TsJPZZ79n9dY1Cho4nCNqckWKmu4Xu11XW+tk318BkPFvFmF/4XQqIR9kt7Uv
vx7Wwb5ncmvoQSen4lrCaa3XlYxHz6Rz94gKRUk/AwzkZb6fbhH1ryAQfRh3iOiw
o7Qhj731jJwDx3lbXyqr4GE/wBXmMxBJO6az2rgEnQC8yley63L0u1NRPb8rzYLL
8BZqqTjoVhMmDGW80mZIrLpvNcCQQwca2ZpSeghuuSPwefj610cJ5wb6szVvZNSe
nbPSQ1kuVH6Xbk8zMMBRjnjqvTrTo/++A7MXIzw6uJ3N8QP8rgG55nzerpb7YyOi
QvwI4mzqyY92O5KmIrR3hIZSyZLJ5cM33ejLJ8RUuqU7Jt/+bwsk629j2tjOjGwm
Z2kl51yaApY0Qw86T+taaqtPY+3tTtgC7KlzGM+fArqIIgg80RAer43kD8yvo7nK
Bo6/tT716lqom6DLB3+6bfinUz6iUNPNQHNTJu0MZqS2Je1N6zZVj1mzW5mw71/L
k0iRGpV36IEqV196euurDf1/h/163vjGw+W5HM+RyxmgbIqpxhM7ENFKNKDQLXC6
77wRsKKXFKy1wazSk0D6zLGo1scS/RCHIB8IVRDAzFs3PizEk8Tj8XumOb6U97eC
DRrHCbf6FfP6sm15RVUdgbQmoLmKgDCQ5m7bX61Zz9DonszlP3q9NFhnxLNTFoiv
OqguYVy6ZhLkw85QKcErXdyobdI9eEk/LIkMbiCbBbyPAu8dNZe5zIZZBRyawBae
ckKi0ulwvQOGMK25jwELQtq+fB+njN+gA1jkzvFi2VmvTkfZykHvVaInD1vQcbSM
EjsA1dNZv0YSt6WQh1K7wPbWp5v42h/ljfLxcqNweoUqFneiXQrAUqM6AfdlVNZw
4S972JdrJLU2/zBWLDiprRwd1cZ9tRzv0ox6oyMktFZbudpxIdlySn1qWoZ/9KfO
e1xz/YIeB96+t4HIF7wkO1eNIHRBdj8PTFkI5sVqM43ICPQUz3eCTuLEgaEQPu02
RK2oTiqSO4UAMhTTWy7dNpmUhqo7nxM+htMpAwZro/F65d5RuIlreTPSi6CScQhC
voqNjlL6ibMasKRDw2TPv3bhbt4RCSMA+sFdvc0BGtCYdU5cvk3ayou4uGn5RISj
YcsTUalYQMF+VBHeXbJyMYVlVnLuuSCopXvtQ1oFi3cBK/Qyyr6a8mzv+ces7aYy
F+80cXaQsQJvBmoLIs+xlcQZGON7OP42sY1WrF1UN78IhAOUndIaRgdulqRjNTTP
2NecmZgRtvJKf88ZSlhxyiz9lP+b/Hl74V/KtBpurY9SNNxc8DVOdg6LR0xpb23k
YObBBQ7bDIWb45CyAq+QojxnvInVwoR0Kuqyx7n8JCBAr3hk67bQm6OnW3dKLBff
eM+l644ghjaMKvIzfjYp+FSxlD3Kw/wKuvlcIuXYKVpObnMDa3vDKNMJmu/TWaJs
kvZx1VdfU0EsV2XT361l2lLIVkZb/R+BWHSA8nnblgYBle19Trk/OXyxHMZaqa4y
uv2GKPgET4Qyh2X1j7ne8D0KnSJ6QruZ/rX97vepkrsco9LySYPzXBukt9snyeWo
Bt+CSHkeA0QiF3dOzidD835OpkzXXnmlXYFEDaIC/0kNQdKI4sQSXRapMvI7ZWVX
0vvaZrcxQ5OYOLskU1HGJEN2o1ivymS/iIyppvyiZp/ENzs9DSsjmsiysZbF3U0X
sFH2Ta7gZLlH8P/dLkEL/e0JE7RIdBE/KZ7oVGOqvE33WUJKtZJ1mLR95piYwb1m
d3jR/ZoQDlfcvPLO3JXmieIQxzvNhGaS3UugEjC0hC9IrxOiZkdoGhWR1E5rPHab
oL7Np+eOEKMWnIscc3D/B3goqOYHbwIJCROrXiXRAw3q5Chjj6t7FqBBHLpv6Ol/
dRxHxnSN1+eSodeCrvwux0HnqOErqGH70hckI4bLxcjyt9DHoxuXwFVNvHzxc1z+
wiTqfzxnVJYxCj6bZQWZVVaj7VyeCbPd7GmDrFejVTmOTP8mcykwGc619ivbKK/o
A7MfJcGGB4J0IKnaUUCyc+UorWL9NY+/J/ozAy8Jj7tbM+bdQldle3dUk+n5Ikm3
JdZFkIbZKW+lcfdN0Dme/zIvqSN8s+XHP5wF5UVNQHlQMEq387iHh/0yKnQN2yWt
RMLnxk1mm7GjThqfqiglOe5SiNNYJ+aTub4GKMGKmfVff0m9e+Wrvc+rPH1R3lDr
pA7Y/nZYi9Drduq7mkTaz+rAsxcWxHihI/zSqY3H87JCoa186WQ/NrLSAJhPU5Wk
yvJg+p22N4VmrZH0GzM1+iqZjTxckVqZyQtkmXV0G91FxDta9R95Wbps2GwN6h7C
kLGSLVmxbgizOSd+xLi+FtwaW1XyGeZa5FawDW6eeQ5TfVPrXzACaIodwkCJvqAa
Ke3mdxv+3AP0oEm+EkE8uAIanL/19gZXMnD6VOX9ayl2sMQiTc+1WgDyq36gQq+F
OzG7knjZXiv3KQTIfvwMRfvLxvne1b16Na6yaWGdb5R46ilXS0sg6U9CbC9AD6v/
/X9yWyIb8Hc6Db9NnHuaNwrKw5EIm01GOiAq+Q9IhQSrRTlEyu2excp79Qi+e6tz
Uvx5k7XNTs9YVBtMM8s9UOVhyHWbN/bYtCAKZpBqsvRQgs1cFIQ8eZpmwLlUFzwD
IsYgfhqehDbwHB1YRZLe2IVd9sr5DNpRvxN7Utn4TQA0lCnwCSZc2o4kaehaal8X
lM7361Y/yTtP8MtsakPlYXzaEV3gzzeaiP3edA/+N/zsDso5rZh/7XTeeYRLT+OZ
gXHqDcLg7UqnrWp4QLSFQqV0XAEwHQgWEl6W7J/Nk0J2SPClyY4cJkaabwukkl9s
3dlaFM03m/3bLxOCCAyZ/QLVylNYENMBjhq8JR5JHo7MuwGCAehMWiF+HKloqjZ5
m6ArUzbihU6detXwyS1d2odhLTE+Oh4moL52KUbVCRPV3yANSb3rK7JCYY6pc1Tr
gImg5PV4SPztRSUk083BYXHU1mK0k2CBVuOumXl2oLkKzkRCzRCqj88CPKW488W1
Ph0J9RComEUA0zy+wnHZKPi2hRRye/btvCE3hgMlrcQI0/MC7BSyQJYVRvgPpKgD
th3nDsO358yYA8jmHBIOEiIrlFSIJQdQ9jGgMOzuwcEGHeGel/mMfrYxpbSmdlwZ
yzub8uAul+w8kk0gqFvGMQxHkj8arKb4awqpkQeJmVjJQB+FkQ9IySYcda944C07
GcBZJwfm0pw6AvNBPJ4YF1A96MnAZNy4cqFkQi4P3a23QXMxDmxR3Edqd/PhEu/6
J2VuNPDp+2BqulMiRO8x1jpV2e7oEBnw+WLJCMaU67pp/7TacwruK8ly2jPKDxED
mhJisK97yl4fP6AUos+JDhudWIj/qwWrd+QhEKkjhCIgvlmJouEl4tGdvZvj+bMi
5on2LAhYRep+U65tKUkZjg++1qRdDUHhVOpxiE9FeSd7bFPJ4duWw1g57ign6JNY
opudVwY6xX0LRqViymvNqmqHOK7i981x82dJservZS+ASNBac8b0oRAFpa0HiFpf
wSQqE/wpTNZ/VolcCrwbNiMd4AHxQKqINWPBNgn5yOoavcrY0z3qA7fzFz7z7NbK
yllI1b6UvZ+j6EcffYv5caq6l5ITq8eZQM9jiRVJVA+iYhj36XsR/m4YUqW79xns
wSVuVtuQDBBz6tK6frfaP8YP00zAXUKJf7sjprp78ihpmerEOIFkGAm1p/kWssIU
6ut3Y/+2Kx8ynTv5WpADBj/wqKkI4I8ujFr1g7al42vyWPQlgqbsI3St7XxiA513
BFYqoQL10XhIupxLaR0A/4fLgctG38onz3jnYIaYWty3mGKVVA+G1uDjZa5LYA66
bKOR7FZxNlLLV92QFzS+rIVyA9Gh/ixE5InApRMSjuDgyC3CijZlQImvJaTP31d4
FptLzZmh5BadbuAl+Hayl0igUyuUzjnWwAKQ12xMhZOVfDR6RCDaaIDbjeM0B6C6
iuwWIjmQIwZIgzYKAitXGpWiS2ioKl1n/ZHegx+ycatbg0Y0J1F23izdDjBOBtTW
2Nb2KWCsAtK+IuhrZmgwjUNAJLJOF7wOoMwQkFn/6gl1SZBKXXiZz6xVumCjUC8C
8CYrqwNcR4A83ozt/0ud7ZaBg6GK16qyTMI//6EhhhbAdq5ZxHLkzliOhlCacWFs
OEwwzObatTPgwl6LpyVKYrX0GzmYDW5oZIh9BzOeZjJ2k8tMxwLIggUS8SKCEvIv
Bh1M5DkNCppm2QO1SOaEUAjXndLQn0NV6kthw8lXAmXB/E6WGqspfckiRkjUu23F
oc+8IV/cdzQVr0YTCVjS5+xUs7i0f6we+P1xJgPlHkW472SMnaROKcOuoqNPYFYj
Q9nnT7YrjQKMmdX4NPN4h3TtbICjj6/Z9xEyN//KVRZavswgX5K9JAOYVCw/L7jq
YUmqE9RWgZQCJPVJcURfvkqHxtYQzb5sJYtPePYsM0FRDVbao5gQFbf7prtfDCBU
9wqHospBXYNsIB9qn29VtRzuqCfJK/XKBYMzdEtP7gUJkvgR1GhJijdewfwlWxng
/RMf6FQWhwFQ7MrT8c3qE9rHWvwJTPNhALhjB8YCCG0pbQq6C5yAfRQY1/8bcr9l
3UVqNf74Pu1t3imq8XCERhwr96qnRSRIiOV1bj8uFuGvuUK9QKuQHrncrSemALsN
hF6j5Y0zSGHJmwBHIdlW8+VXhPhdCkj+2f6lv4nJJ3U40rmnfsxNqFrnhjiELC1z
Ky82FU9TtEyuafMmtpkY2iZbVcJjngKDvmwVSYIr0nFzHbpkX2nsZnya0e4VbEau
KzF4yGG0br4D1qfggUJoCGPZFPauVUdZfFA6Iv9E0BRecupHSmmPOwcJi4bzQfln
dyY+aDn8TXi6eXdF7c7PTEE7pcnmtQQW1WRwTlsOA9u1jLhIXkptpJRYn8RXVIYH
OditDCSoy7dRIAH1vWQ/AfXAUM5njL7r1N+PmQNbp9VPHHbznYqo68QljXPb6nWd
0ejjSm434ZDH9aHthcMZduCJnav4jfYFGToncaCLT0wCCtBYSZARJK6Pyyg4U1Vb
OZDuhBIpSiTSUradDnKZC8NNbf4biZejXQGEqIi1+BPsAQSuKvYD902J4muCes1B
xTuqWVKgpTQzE3hrKfbDUb1rKWDjIdPfCUroUWgNBxQV+tXLOR6Ue6xvG/n9xBgs
f9JSq7l3B2GMLW6s4RHO/SxohgwVF5fxlxt9twpn+5Zi0U4tXgcOyi9M0epBYO86
rSU8jE3P+EBTlWtI+odyUONEn6CPEsd/to5Pg+GZPaDdvEe0azCvsf7oF9HOMPz4
Fr6SUfeRcyTGjjgfcY9NMaCQjfMXFK31rJImRbBoTzD+6w7oQxk1NhCgBjKBI5r/
gHofyrR5fZO2d+x/aL6/t6zpuGIe2ko6a0x37DAPCV23eF5Op0eQq2SXVqgeZXdl
7ZI41BLDHos7XYnhpBD6Dl1zbZBucEK2jiFLyqGZIVgnOKQm3np2QLrY7a7fTr38
KTH75HnvfpagPtyZVQjLjPhGx54aNEsbCJR/4a7v+HkIAXN/3TqBT1KZHW1YG+2y
MTLyIVEx2gFzU6AxbdH3fgso429vJKkAP9jUIBBpylj6YYK2OJeA+CL8/eGFwt+J
xs2Kb2WOczrrp4p+iN2HLUeM87zrKpoSjh+vIAlKZgh79Qgl5CoIkS7UKunxdEbC
uNJmL5a7W+7fvC4HVItXIpJweUWdoEBbGV8o+r9SnnyA3DEKv99RFcO1kb7Oyi8i
YVCxPHU8T7JsOHc9wxcS9v/KWR5Vf5AMW6jW+fvXe9myTMRE67Zr1iwYu3sCMXDq
O0l8AfdqlMEHZnPQOgqfGLEcAGXJ8uaOPYulVj6U/CFfflB2cJ7AdHTEoRtpRHAE
0D/B2THWspItWSk/RFM6X0Gj65+fxVKK8qYhFmejx0xct0MH9+fRuCjhdBBrghDE
FHkRoxdvKIpwtxnwQ/9wGmw+eVAh995BjhJVE1yhgeEsrIcQTVWNozn1Sxtund4Y
/i+YxW2fGBAfaWQH3jC0ONQz64Xv5QUG6VpK+fo3TLizbq/br1JpJkJYmUDAyWEw
b0NaH7/SMHu2EDCzLOmzPW+mMN2pbkKx25rNBQ+1ZL5wSqqHiBB/3RbsJgdlmHzX
NpWf9oDi8ru43LOU0ZgpQM+WHTNSeFWQKFfukTrNShP0rgKuIjzasNTVjTxGo6tq
5Hb5sThHWux+rtVq4HLpbrrdMX329lDoAC3+cxpj8W91UXVxn1SYwiuRLTNHOMFa
QT3ay8hkbirRz+d9gRFLKWhpMX0M263Eu+1UBOq3J8+Z+jmU/gbBtTiqipJWY3Jh
ilOm/OlrFZhyDXlmWjA9Tw0BTDRG97xjRrv8r2gb4PNzA3U0Y4J1ZjGPe10Fs4rB
gRID7rPxe9xDe6srFYvy6EjSA92PYuuztXIvsL1oUUu2t3+ZN+88dVI2GQud1iYA
KTb9HTjKrJSCo6TEUKW/5y5n+TOoHmFThrH+CHxv1DL1fdXCLhV5GyS0kmI26oTU
5X1YDueAkw1iswXr3z9hmlua7dxzlBwgVMXB+8b20M1TOzvmzZZIQqP7BY+LLRBi
oMr2fM85K7mKI1kUyZ16+iPV+ToUFpYsVifeJ9X1swWE2Gde94eXZJSkrL1u+dOf
j2HPwexHr0DohVVngq6eZowYrOJkbsUSqLG755DmfF+q27zSJ4pogD0pO9trsDav
8+bOq+2gTVewOP+p5I6n1HwJZhx0oeie8kOnJLs/6YTJo4exJrX2vAvtpyNtDgaa
ZBEcrpD/ibM77D19j5Q5JHPB2IwPzstOChKSNDo4cLshxdfIGizY8LSUfaVAeHRA
n4CxbQrI9t2V3d1e7AUkMaGka7Ato1Uo1u60r84ltlgWCB01xzbUKBM+T54WuP5/
r3D21PMUCQRFOljgekQlIdI5gBV+zKqOWM3cMFOqEOKECu6H1DT7uvKUQcFeuIL2
7CmRVpgpKXY1chkUCWjcySgBAw1tmpaM4utLBWdmdenlJwKc9HsnAG0xVC7bgiIm
IFu+sN1eQkTrj9kkXnaEULVh8tkDagz6T55IEZtwzNj6QXweJu4ZYlbz4gMvwKUd
85YhEEJv8fQtojMrSt6ROasBro7+KiTOv5QyRTg6g4QErxIlRc9wC0YVD5YhrOh7
I8KwUkdPa+xzxXFAYATaV5hmY82yPgWmbxgSi17d0uQSu1YWPn8AP+JFbXCPwXs7
Xoj9R+9+9+x99M41tYvTIeNBElxP0AAxUHZlkby6SnX/vrxCW1DLyoocMjJm2OxF
p3dGcTrLzzTv5oD1g1B9/1VcHPUIOXCLLRy1tJRtznvHg4fJusarvnYAN9Lygwoe
SaRsn8HvjvOiLPuZ6ZBGUoVgLAUQa+85Pubur6/SZEY0hGn2YH1K/tsWY/In+ILD
O7FMwBCLGHUvt8nLzHarksyKwniJ/qy3zMH98ykAvQAePd/6RV5c85T+//PetExC
i97uGJrxC817zByYi7wKkjMoYBny/7tX08g6okFZJMUEexceRgT4z/ko2qp0IKfi
5Vs1tXV5O16rgtGVEKnkW8dUO19OUyo+edZRCUj9QkyuTV0yAnH8MxEK9vJZsVQL
2EvfXicg4AWeNcZ0w/Eu+9krU8kTnLy35ylyeIsu0w+U9p6d7Cz8hkIBO6FJyb73
AZf/V+ND1T08ZsQ+U7AlD9dZstZM1gD2ggLh7Cm1U5cXV5fatbpOOcUWQoxlbqkm
8+n49iOCCrCIVbv9nDmnH/WL5ZLus3y4WbZtDji4O7lYMTC7kOyVmBqQjaYQXn4A
FbXRV2zTU3B8L+U+nWv5Z+ayDwyQYF4VcdXF3UCdorCqWPNmjS/z/Ea6ll5BkjFt
9bSKFqQF/YFG2JVx/SxeMH35+fjM27h7/mKm8d8nQM/lVzfs7XRr6oyapUdeCzJW
UjFVGm0E7N7ZwUMSswPUOklYzOWhfSAy2m8nZa9Xlh+QWxGBCY9TDKZHzUReJ74t
Ja6+QGC53MlgukBFRPDncL00jHgaPLcPrvIet6/2jWzpTMTFxWGjELgE/cYCx42B
QKIoTh9ns2yiMcQV+UpWgkL0sxUuO5I7RWL/v0nhmCOYd91NQc/24qe8gv7sfFts
AncRUCIT+XWu0M0JKBKOXNJti0rClPrTaFTs3hEo7wvg862jBqRdDs53O1EhMd1e
Lfhag3vqpSDOsK521iFn1LPkLn87OzTqk1qPogJWLNTwX4/QUaXOpoHLmKwecI6B
ivSNXwX681th8Y5HTsuY3e8G0AXe2KgF5DYis41WSSoASTtiGxfYTrX7/mXMOSuu
Ls4gtLFSfcEjKvBAh5DBojprrC2WwTbZCT4TT3y2oOUVjdeGOuLeH+K6IqfoWe+9
00DN6lSvwhfGLP+deYIt2de2rd+YPCKyrRbsI5QlGocLdcEwsol+r/10OEiqj5kH
yoRHxuXKBBiiYht3PBMwfiT1uJ55GgDZc9SkwlxlFS/7PJ+G2FyNzCD8LLtFVTwB
5DVLWM5pFen3oVktaZrtRSSx9t0JV6Yo3MuhfHMMpFEzwlPQW5NeOmKnIWzPX9AC
1ERMXckTi1nPPAZxI9ZNSuWGQim0dBGzfCzjdQw+RA97CrVgwV0kuKh0X5OlFbWL
lx0oj9kGLW1JLdZGc41vOBbpB+dNIbgXc9B38kQMEV2Agb03soF3RHlOdIOyHumA
swcFFlXsP4X5y/X7vXvhGWo0JSttnaMFlGhR51hvG3xp/Ggc4ehyvejLvJRuq65B
7s70jJpSM5YY9VrG6G2+bifSmpUUV4oOS1b9BWx6or6U+gUh2g6odAcmNWIsfPgL
HSJzeBt/iIjV5mqZrgLlwAV/L7WKGPqfNi4SbRnLj3IFJWmbbbytf7Gkr4BPWaNj
1VNZuDCOF5Xow0O3sMGCDRO0pvDVqfWfdzY+8426WpjhDnkmn/jO955rfEtzaBCa
oPi3QoNL6nM1lFUrVLVFCF1SHQuDs7gZ7sfjamBOz7/hSyk8qlrncgwWmUGszS8p
VkxKATTERSiQpvb4llultWMBceYt8PEgWXd+nKZ1Hc3+idy97IdzINlgQNGO8O5d
sXsegwGvpxmKOnhp1u/+7npEobRiyWZDHSXSGbMnOi4/0uvIFK5LbKjHgPY5yS5I
2f9RdkRPm63mDlvcdHHXHY9zLOZ2kwhYHQIkqEXYgEkKp3qB9761YxaKTkCNkDjB
p0Bp6DmpUCXe7YJQH9kGyu55YkQvwJjVbHzxmYUypn8o3ltQzWOQGmiPcnOOF0xF
sgIa+R/a1dJuIQ6rwAlGMnKzHtz+mlYUmlyZYl0KJLBVmyCUjIYOTQ72aLy+3JlW
lvQ5vIOy1QfUx828L0TQLkk5V4EgYPa3KRYlZt/lkv+SCnjaA/PoFjM1Wd2yMvLy
mH8Q16FEOvs7bRf+h/iw/R/BYGYvyJ0YXDGOByv2JPjtxLKIBQrBOVGnNUKHktHE
e2PYILXsClCq/7XT6NW02PMPQXYyoPHuBDBFSet+CrLDMxGReYf+Ocnut+Iej/xu
sFaLy4Cy75gNhxYC/WQVg11Bk083HBHCqCkKeomj21JogzxGjRaDPlhpCd6eDxsx
Y05/xsXBV7miObwQFXXiCdTbsQQe3IerUfZrsp928q1MbzAyO4uBxUjUVmcEmU6s
70WxCNaGitYVdjtx5sxDkZfL0Isdg5k/t5O4+TkLbKjuTF5zZSE1s0hXb10uJeyM
mpzELMQP1erN6ElZi/0xAOqoQPjN88kWYFxgnjYA1EC5Tn8eqeupYFTe5XbBhzMn
qon+LRUPSpX2qF1xrnbLTE/67HtAUrVDu+l4PmrPAudwkDHMj58SH3as4WI+TKgm
wqc8TjOEJ/friFRjmo1BGSIRJVz5503DorwcBM+f7qNKGlQhN0JLVjbnorfrtPEZ
ZI9IT39Mrh9ho4QMznW/aE1/ndFAiMZoDS7jcRtPjSli47KzOikYXVpwKHDnU2yr
ZrovW68rgakKqqos4oow2Roma5m/XR5+Z+BnMigO/D0GZa4uE+dcAWZjPF7bJ0GP
qf9LfQ4fQNF24fMX3659wAbcVjbVShV+kb8svP3Dq8O3gcZPCUprSdwAYpo7B9WS
pZIvMunp8UnXSXd4xGxllxSIOEsY6INhrH7CKwaEMEaGCDLXqKuQFS0grlbfzshN
0/EA/cJWFg6dB4hwVNJxesZgY3Cpkcak9qnRDCXIEOTgNv0l5ECDyFxrZXKUOv5P
6/bsO5fFTr9ygFgfQf8g4Gksw8J4sZZRDZ3mzDhxlEUsTecpBKtmVkqX9yMmH9m3
grjBB38SvWIDiRs0VbYvDwtiqVOPoPXGDvHTlDaBrkdDz5Soxfk16/Omkjgp0eZC
mDA21laLLpgOgdlE3SjN3EVoQG9dgT1LFmsCuLJEgb5hIw3VoS9bi0Eudk8nsnoG
ygWV8cF8LVkdnvG+NDXDhNEg7DvZ3fYzefrKhuwY3CLUJSfQPaOHe2sg9YlnMMC0
AYRda7XsC14C3m+CkAKrPyEs7ar9IDYZTizvZGX9g2eVZu4xHgdEr5whHil1dAJe
niQf7OM1H/bAwicrK4e1+000u4mtSXJRph8Zh3LE6hyrHAMUL8kQbuXnxPbvp8Jl
0LcPz+Go/Ag2+hdsG3mxZ4sSvFDnEluGBCob/FKjAPlHK7ovdgRi9rUv2T/wnZ7W
YJkul0ASX3C1umdDmOxWUEE8YCgatoWOPc9YiJ5Sm1dq8qqSIN4HY0ujW13se2TL
yjB+YK2ecyKmcsiXfYWELsw4qtdDRJIuHtDC0jc8HZtkl/QytqECnOb6I3Tuj2VD
UJ0SomC55sm81MWGSEM70oUYR8zvmvtRyaVOQkCcFY2pKjykLrHiq8d2Tw5PJCCg
o5EXiVMIkAuxzrl2gGOxT3G7D+MoGxYOI/QjbDT18kDCa8Qn7j8s18YskQzVe2T8
4/sUmbYSamz9tDIUQ3PULDq2D34IJ2re2g+yFueoY7yF3bVzOPUKhqydD3X3BBaF
GtzzID4O4se1x6Emvm7k9cEN1iuDx+fnGKHlNQGi7rn/lTgO2ZhaI7tR0IPNhamT
VcpkLySgAJxxXE3VPwFNkbf2wqSTpiZBTa9Ie3aq7kx/d2GlB8dkpbLw5DSVJHkR
oM+u89HFC+y8+H11ur510al4EcB/SV7p6I8H29TOTmA2cS8Z+L8+jgxdVZ/NoVS1
r/QGVvFW4kWBEHWrd2Q3ceEY+aRvcoPuEGlrlgAvVkk/8Q+xwgGDu3Q/6MQ82tiQ
nBMyj5HLuVHDpORq7nLdpkKuJFtTgf1Tq9F/8zSYnHdMdKY3FwQzGXi7gIVW1uza
fbQBySpqvcNO+RA2x6QlMUX27gG06jpV5oKRHrRPuj02DxcFP6fewAmGjYti8R/u
FoLA65chsEEncnQFxkr2N9zS9oVuuQnJ0dQc3ryINeHSkWdFS+A41pn7xeAifKrj
mB9iekrinBWaiYnno9cvWS52OkwBvc7l2nmtEg8psHVV4d8iyvrMvxXyA90g6JJD
o2B7ptOlxRWOskdd4onDAhlvkHf2XNDqNrFNeuF+4C9aFiQcXRMDf1/37s5miZlc
q9JVkeuw2qAi0+luRkxEl6JVo1yZ2cjKvwX8f2SaLr9brCyJhV68pkmXMeGhbjjl
6nA+FaS2B1l9py1+2N2MmQJINqjcFm9YiPLNtV6Qv1qlwFZDxZ8QEmrFSSXZrEmn
YK8AAx0s0lX7D8Dia5gHLNEemqWA7POQ33dpDXdBmJD+cze4vF1Q2JKwGQdVCatA
rWFN4J5tU9Tvgad0QuggYlJNH7TuZzpllB7StR5Tti4Rv4Ynb2cMr6IR95bVyp/N
LinhzuXjnxeq2WFeOXNY0HTo/9WCm1Lf2GVdrJUgOAzRze3vTFbe7w0SpA626+TM
FbFxaV5LOq/J81XeQnPOsZQ+bxQzrsoTJK2NDC/ZLr+S7+irjT75Us6FjSMMibnj
dp9QzonKFtOh3d3/7qjwpS2SZD+YVXKRwTxAfdmnBI4Cp6VDcTO+Jvzi5t57SPxV
lY17ioAyUFkr0d/nZ9c9x2m0VJOUxefW+zvGW1sfx6OohtiOp8aU/C6uFvaULm9S
E+sW4ph0q8E3HSFycbou43zr462Q1BPCUmY9aCFw/4L3bE3/HR5HGJttblRtjBYf
rZ+UOesNFg7yP0LYpwTQV1ntUZdUoXEmeFO0TwXdROuNPE01yAqc7nUqZh2XAs1c
qgetsQu72qD7862gI4qpK80tdfI/igHeHInl9LGuy3p4LXs/eo0glOV71v5MU93z
NWkPV9RPx2vk4nDarDFBYm/uaTOp/+9igkjq+18jv0vyFRdAs2rhc+S6vR5C6lwh
BYjfdCvbnO32pHb7U7o2TWxHpmItx/yWdzX7pmwt0W5P7kQSigihWUjKeYCzqouY
QK1PF4zV0FgQIRkUkaN9U+LK1Mdh+24dDp/iWo6clQLJ5hmiFRwEYPpXISs41Lf4
W+Kjad8kEaa2L3xM7wlAJgSEoA88GVFzP8p6LjTf+1F70DkxguGineyoUWuuVU9c
otoVjt0rX9kt04800U4jg3RvWZZUdYrM1dLVTw4DGXR1TATjz6kLnP/ydQi6hnNc
t0YTgaKllnf9FHqzUpDnFteCZU88PlcmvxcPrVNB9EKrlhA054wbUxMc3WOHXo05
YfoL+q4jeYAITLp4ZfaqvtwdD1BFBdXdCRKJ12A2P9kh3Plq6gvU2hs/5p6s3t/I
VmIuynIZzxcG5AN6EGtRbayGpUlFYb9rgMacnZkoGy6uH+gt5LuUV7zaimNQzZcW
KlS3haoGf/Hz1Ot1yRcIcct9OikdmPpYicKgUHly3R5qp7xJKQZGsAvXNyWLQk9q
65/o5NsbqyjoCH51SkPQ8xHjG5Jlyojk2bJOd4a/qBX9MOzLiI9e/pO04xGRgjdt
H8JoMSG+5kkvfTI1qcGZuPeYU7YSOjCpS04RQqGzRClv89X45hx+7kZdcPNUju1K
syzC0BT3zEd2/R960kAhsg+YlJ4Bv3VOznD5wYLBr1wng8B0whjJ2WzwIjzH1m73
DbC1z4GyRIttcS/R0O/3Tno52ARo+01xtlTtEvY7NZoHWE20ABxPR6MVSzLvYCZI
vuFNWw69zXrAKA/BsgXN4/NGSKrJtgoXshplAmzKdEb15r6ERihH80B5r4v0TMf0
x3A9+gCE5ur9TW+Elf+ugGkCluSzNhAvjuq58POz9QOITxHQtYfj0HAOFZt7KsnJ
6R8B/QRF8mTslcz7ROab9/Cw0ERO16BYA9Oj1qzigRjQtwiU/DxpCLs2JI5W6it6
nF4tIPox8JBvi+B2+dV+7H/56otT/6dS1RosVHpFffXcupuzE0MXCx68mzSZ6vlp
ugp9FodhvXC3d2YYmq1C5vyLwy/DBxzvM9S+p7GUpXu9e7dEjmOAX9NMfprx4xg1
KQKCZcNUZDkBf/TMh7sJnxyZ/GzLCT+0TU9PkY5HDveJX4/jpVxkFRrQ6iical+f
5HIxOF87cQT3ghzyC+9Baxjjz1Xb15iFKUuIiGDzIaPutbc0cenHhsAD9c753KnK
QtDgdfDBuw3pUg+/LR3b0kZhONFqCWmnlDyXH/ny6A1YdIoahNX8BmtxKIornLPN
snLPHVWOINsJ1LC3R526e6hLCFGM5u8dCYQFftcmo6BPxeek6OPhkKwFMqvfnk9E
SzCBAaPGJ2aIA5nRYRip5U0w5k72nKCvNBoHgnL4M22syJZCzOJ24TlfMcVhvYvE
pkXK+DUlbaIJlpVhEg31IW+VZDeuBc9NLr+D4FsU61y7iCf1G50SmiZRalLufZVu
mImwEcZ4Pop1h32swiW8FQ3+LUXkTKy1VDXCfFVBC+GfcSl5b8OFcndFBgqqg9Gk
/DzK72iP5NU2X/2+7b+U7pXIr6qBTJ/DTw+WK/Wq3/FLMsP8ER1gGGhWTNv9LdNM
rbbr5WBaEKIfjsbOL4EA+JA9N9O4OtWliPSiOSVTjRgoMaejr8ukE1/A0ZvzAlZB
5FBWlv5Fd2uwQFwSNstYdRDot7TiZ5BcstXNyDif1F7z2aL5uuXJiYYaUvnsi7sv
MHOXXtO2dXgSFFAGKImpg8xqe58+w2KAe2UvB4E5ruExxPJEjcpl4XnHpFIvWuV7
NILiy52wuDOcayAKgvYCaKygIa5yh7RcGKLySjZhfiHhdGwZLKFwnvgIw6ASfGsd
Vfh44OkLaz6Aa3ApIPckmSR73USdA9Gj0Wtkw51kRzPywUnKkItBx0Ux+EWQQPC/
nqRiEYaSCmD+KuuHtKmShWIcqBd6Q4mTCLbJ5gVFiLfv0SWxoIHI5S8CBJ+akSNZ
1XxBQgxmROu/GO5WgUQBGT2kmagwoAdXRJAdCyWcLGzFnEyyyWk+JXndtbHeN+/T
9Gfci47IcYaKkXAMCJ+q7CE6BUyiJ937l6fSkCYMSdh9156MAFSzPkm9HaH67kpD
L5woVgBM692CQEYcoX1FMvb9uwvJMEU0lsZU2gRIbQQ4jCI8zc9zeYsCTlELb3/j
n3iFIffZ5HXTD1rG2bWu1oPnyUZJoaW49jf6U6pM2qIw4ifjnjVwJt9ejXL8LBdh
gyh5q2DE0DGfKjuZqcrhi9NLC5L3YR7viQI1Jk+9Gh45UpiqOixNPLz4V7FPqfwN
kdMqdMouROgEgrm6hITc09mXWEIcbTEImEF/nBW7pxWITGrUTyXFbh1BLkFkjMJL
Er4wHnpUjCnVnjjFoqr0Bc5iPm5dvN4CRvoFFJceB6U684uro/IR4ZE52lxjKddd
wdLlEQPLTCaxdphr4SUR3E3HzrJd2TmPh1Gxra2E/9turLrQ94yYbBEYtoEX31ew
fCtYuYsRezu6woKP9dO9WdpzGeIcmQFOd5mUBhgwIqFWxAdEVJUcTBwUUiD2WJRp
ZPSWWoJ3I1i+hG/TAmLvPy0LcwkFjdKRE5vvaaH+yWiA6iJXvQeef9wfBNB3H77C
Sr2KZfCERIsG6fhOdGqtyGe7p8uCh8/R8+L1IU7Wpacj9NgItNO/KZ5uI5w+NEl6
N6F3x7V70mS6ifuzbp4h2lcs2S0aS9PpNX5Uekb/20UD7GVkn6OYg1v3nGCLze2I
yTSahbA+RovrKKr1NYjG7NqZzjtKWLOAjWmQX6st3HzORkcgc4tdroVGCQxFp6wd
jIm/rDqi7erqk/1HH0RIVgnWG3z3ngfIMYBrE2Ou06YkELYN8dFG+02q+lJdbsOc
PEjQ5vnwtLv7dFmjJp9YPLrCqqK8RyQzxBeY5Rmpgjt264Op2hfMrrjIAY4ClHzG
m/O2QyGVp+GWAH9FqliUqK+TXM3imouKhZPuDBACwjiT91rF3rorxwUXvsKpZSXc
h1wkO2sGhvijnj0erpHvFxmoOKfMCU/Dw348i9O6bOR0Ylxb/+6I/6Ww/ca69LbF
IOhxwinRp+WJZwL2L2+cAQZbZemaO0Sj0MV1XNC6FfD2I+WflEr9/ilfZK413vn2
bvs9Vx8rmK6tfo1dGTl8rI49Dyh9y7+oW37kIZC29YmClanSlWh3xgcH0vgerVAN
f1bkNTzSb1ZPz2B6WkTcT2pDhOTeCEyk5/OYunvHZUee4t0nUNcNkHwGV3LafnaR
2ZK9J8t3lZ4LB0G+QfeUkFzPfWsV86QgFJQaGS3f5TTy2fNkdub2wXdXl+cODrrQ
RzV0KDjLySlPyAsTivvZeGU67uKmT8tYkAgfJxY1EqTuBYIN3lsboVSFoenUvh28
78S6GCuO0RIuLggJrV3lgvp/ap+WVXsakR207enjlZiwlwx5nkrL2wBQJSnMnLb4
8EMTbxyRi/+EoP+4zSknT1Cw51Bgt9NkfPVA4p4yX/SoJU7XoavZHt23e+1Q4Qfw
3CxhN0IZpLSrOqe729LXb6BnDUwQBTw/AL1DzXfySULhAuWLz0GG5TNvKoOsKNUO
6wLH/pT6LW+gTM0egSzT+wrBDwJOFXdLeLoX+Mzqn90vG98CBvjvuS3BU8MQFvtu
H4bvrvjXDGrYznMMiIapidna/NCuwEgR+s/GSD2vB+7nDQ8IP25ejAxNa39joCeV
C4UwyMsoS4YTDnBcY8SUVYcScz4SRz1+v7U1bnF8L1wWy2M5ongAtVQ5VoWmWcX1
nsJt/lzWxXBktb+Az1nHtgKUEc//1nm+pEuLrDyK4RG3wG+hY9FGNIxZC2j8Gp81
g18iab4XuU1DAwn3ToQvYAwaxgFsq3oqK/gEfk6eOySlv7BsQ/ZSn7o9NGw60ZEE
grCHiwUofZ6oV5foBEh2BRZk51EvAzpBKjr3E/pfrYdWZ95li+sFe0vxFZaOjg0O
E0rO7ZG56ILSf7KzmGFixY6iCkW1S/6ezYJvsAv733/YU/MNx3pHaYgEfBPPrGCy
KE482TRUUT1a5IAHv5Y8SlYGymYZ+BeNrbk+0npc5t1F6Bmv/qD0DBBL6mwPx7A+
sUUigfisD3AyGSic6TavXmBmzkVdpX76aM0eVi7CVl/+2IIVrgjYEAJzLY4PWnlw
2OYOkI+OayhlI7FQs4Nt4/NunmySOPiUTEN58+bByEcQAVScnkNTNqDUMAwU8UN/
KluB8Epp5AY+IxMery0eOfXEHTm6wkT52EIWWmivm8hhTG2NadbFS2r3ZYFxmYi0
kiBWMUy8j0Av8AztqkTFzxxyMjaJGMNw9QWXWFHloghsjWUJJo/OhS71FnWxGp92
FamRPX4J4z1x4L9GuaKumaTpJwo7XiwI2/rYzyiG4mxf9MUTpQTUmj5IFwX7kEkz
4wDGKPnYNy1LsXICQM9AZEeSdLHEtSNgFz4Rj2dlYKB9FvAXyxDEzTc+yvojGz33
/jiURIyPLHBtn4a+/hmPbBcSL/RWCBAt85GL5JEg+I6/5y15KmWdKhdL+TwpIRG0
oaLrgb5BnlRS6LAn9UyhC9XrXw4KCDnxSBn6H6LjWUZmom8k8nP6F/fShktEbtot
MdLx3ZcbVERQ5NB/FHNRmar/P1lv1s75PU32afwZIrXJyUVENL7VMYn8wZvnBqlF
eaH1EbkXUZrQSE/ELqHMPKvwk0H5s7N7/XplqrpPEM6dXddRsp1hXyDebf9iFCVy
ItozQWfkFDonT8ruPUU305Sfj+Dioom4uTyQiZyeZxsinCTGe0L+art4zY4M/3oK
bbujo42LxqFX+3qIBsRzXafnPOFkg9HUNC55MDE4yPm5kLlcBsGRjeg59OBAjlj/
G21ibZzlp7ec4wbukOc0DwkMoqvl5VjoliF3qmCrnyR89soNe1yshHzqXGwl7+/H
DxRqoUQs9XJ5UdRfJkRMKMmaY10cpL6pRNDOmM6O5EoNmaqV8oppKNaX/q3tb4v7
Zd0Nvwiwf3R3vJEqRD7797T9YLOsTOFJhAsYB4O9wFJ/Qv1w3q820km2AIt+sW70
vpVi9kZ9Yn6kJoLRXqHiQLYvVm62kpXcKyqpnbQCl1Tudep/t+tUsRbxcXHe0UgQ
zuqIH9u2w8wsi1Ut/c8Vvfz6Nd8ZvNsGW+3X4SVwDLX3bHykgaaerP4aJKHZduCu
KoKRwUfeQLQQizwQw5vKMIY+2ihgD/NZiC14u/l1hDDhwbXgwbdnO9KSrbuDPkQN
AYOTCyZedjm8pKRlmIHixyCMNbRCeEkiw10jBr9bRMwyUDLOWIFq7R4gbzsVIChY
RXqCB2Z4C9fNCub/Da5KoN4yRZmtkgguCOFEoidzq1GDLOQctKetLFH1r+pCpeyB
Nt2HG1vKtl3mH0G11ISogEkjprmkZbS2K6Ak4oPSufbAAN8ltaMG29FjAXI8fD4B
zECpIeekpvLNuktcyWS4/zr9Xa7ob6Sas/UBoqv/t58yoMRqvH8uDCjM4cw5+pMe
hD+37FhZSez+Ig8EeBXwHknT82bm7UiYv32/gLNJANGWNxmZ3vf+xEz7hdXaEinR
wmnL2HBYid4QoDXaXED+ledh58sim/OA/5yfyTW9lXf7KjWx25p+WoU3MAt7384u
+lfFLUM6aWlO3MPGPtjMYp+lqsxbeWGOrISc2jlXGGh5k8NOPttNGiq2RQBalcF2
8WaPdHn7O7TLiPfQv01Ci5nXSbIxddwfl3fQiw5TZGI6nW8e4QeMzC+KRzRuZdic
VNHP9G2kCrf2KSTwDYX5vSqdKMd2m814DnR6fjPiM0IQ4qF4NipqKNe8Zdd+IigO
mL9QEC7SgPSDBFrgU+1vXFSmnUzv5I/F8SPs6NK1KFHVZF1L9IjZjLF0tHHoLZSi
+dQ3IB4Lw15Lk5TeOH6KN3Bvuih+erpgI9I//zb1hkS+9wJAUyERZXI26elTQDso
oEdvq7/yPdbLaUJ4Vpv2XhdNp9KCzw9vAB8bW3q/V+LcozAPY4rIiI/tNPw8dic/
ZY5TF74QyCX75PZanMa8O5460Ie6+XnAb1cycJcoMGylLN0GqJAgUG2oxMwy7nc5
S/ZvyrMmWceQnm80RgxjgGLHgfwB517BAUNw9hHwYU9rnA+xy1RxPyHJonGsAbXc
LyFoeVVYEsi/ZPp2xYWorDaTMQBn0NLaOEi+Gppqpy6f0439R6fw/XJZ2mljdAkQ
iLVNa1Aaq9PQ3VIku6fLsfW+nl3/h1B7tcsWcPHHJxrJbw1CP8pl2vxYkUZpgeki
+N9FeNGwkxjrZCZHfZeJg5/x4blB/UOxrwDbxwz3qC3Ft2n3NbhTEqhQTB0NHlLE
cnDOenBfqKYPZNXffXJ0q/RmMXiIuTTD9BM+kk88sEIYXnqTE0GdR5n/dcyJQ9ye
cqTjh/VNciYnBhZj5GG44Uvy5oY4V5+e5JKdHW5Hl2THmA6eKR6WmLv6eqrwN+WI
DF5KRyrnjHO0SBw64afRcU4KlnzXHnapc8vmmhY7xILQxgqaL0/anx7vTCkjMxs7
6yzlw2EWjHdIL3ZOqux1OnWwMcsJej4hPsDZeB+YPilOn5PC7vJdJfF7xdUp4t9Z
Vf16MfnAiMtjlvYmAxaHTCT9eYTwSefA1AqqrHSwQWqiDK3yxiYYHrAdtN7pM3d0
jV8gPsSoTINV8kDEoUqatI38UeJcLx7ITEc/6ADNdhXAmYMoY0BtwXvZdPqsPOhO
etJI4mY3WvooCQEx4Mw+0smh5XL9zMfppoiWiCtrIsCm1GYW4KxPeKIG726+97Ox
wQi78WFVwdUfxi1xWD2T/4+6AlRqa1DU6ur7lt8ivhSrOX37SbiyCNOXKV/prYSh
HWgji+oS9lt/PLqkzi4iZ/Ch+vsxhB1/icJ/VIulq2Ju/nsF0b2cVuf3Wpx1wbVV
u1WW/QP2nIY20fQW+cxhjIFgytkXF5+R2yAqd1rNiJDXBdrQFZ7xqFU8zyH32Hln
TEeWgVoe5FJS+A5LNAckWdFWbc/5Ar6GCJcpxi2093YNxR8M3/4z8FekE4Oevjm4
LacfnLcUNyYpRFK5ahJBSmknzoQBU21MKYCIw22XGbZ2nKcnKFynSJJ4pJfrEKlH
TNWfw/eKWXZLKnyoIJU1iy5pv4pLzWAMq1kwrkzAVsGPdkTo1D0IDhF31JjomVD+
5h9izxxsxDZgIxfoTxVhFwvQxQSmJwQIoFXcfaSbEuzPioa7jUXWBdd/XYpOZT5w
CMez7npKxEAyPfbEM3jsz8S8DnPO7hnbgSSMoFAevvyxWBmyPZcl80FBANpuMrox
UmYkXwhh0Eb5xN+10ZJO73CQws2B1qUpuy01vDHJlKGoMWOJsgtNj/OdHfN304TI
N+pLkEFn+kLjm6i+fvWInh5iPwSQUx5mPQqEXzBtsrvUf0YaJDnmekCf/CLMLg7k
dQorEJVv4SrdGoP7LCPWj0XH+Lhm0tw0VFzkdkY6C4ysb7nIccJHRNlBoJh90iec
+qINeQ6g7wbLOh2OrsWyg74cKqA5Eovqi8qEi0fTEuPxWZea2G9/TWlILebrdz97
HW3pKixmRfGy6alxWz6jE1oKJUfZQfS9e7Y7vqhKdLHRa1BQk6n7C3NC6vYu2/QJ
OjL0XAV4NOHVh3csAr6oCxCx1vXq6ssbeaJJzK+P+uscX17CQBzpU74EVnZSJKeM
5wwq0UiqGmnrfarvUcyq09lwgFNDPPBGPL9ntH078uMvx/6JzBmeqxo+Zpz34oCi
h7l5snMfhVxOZMigKcsbWs1dY3K2X8Fuaeq6pmt7gLxGISAJmzdOLcUmioan+mRD
tA3pbLBVG0HYprdvUg0M0EJQseRzg7ZJeQ9XXswTiiLF+FIdOWga/ORdZyCyib+a
K0o2uTYnvbfWKQjn1TBimJFB6XRqUff2gTyUSSn2mrSLWxhzlXTWARx1Xxkpw9C7
lzWK1CmLmR2twPBnj4i9uPvXNZys44Rm3TF7wgnNGfRLY88Z9LqJgxsQb1W0ZEwb
+vacjEbtsAD/CjXcJUV+sz7D3tSxe63pVlJseM8EQelw3xewCmEQYWtoKIrPNWSy
gYM2PUF+y9iEMZ0ZHaZAj5mfapXwHPFgvB31hOpNMugRUgnSnZqTUfu3S+CslNMj
WfyLbOeYY0P10g5Q8VUtEi7TQuHCEeSghwpHEboVgbVsQMqfFwasT7Na/hx2BbaG
doPyFvNZaXwYCPoUJDLX58yIRq/FTMWowJwGbXjd2M0aJrxAn+kJ5id5tdKmnbF6
ZPQcxdTAkuN3jGbIsZVi6NFUsCyIK3JxYjtHTDaIhMYowy4B4FoeKrDi5vWyPRvO
C86W29xH2JAzcgMU/TwKG8laW3c690apxM+8K+/oELcjJBul7RH1r3Sv/w7DF3bK
3FzIhknlVWV1JcVcT3dqS/vkZz90VgAjDpi8RmRgItG1lub+hUxQ+f0URX8/Dwda
JJCiWcC/1eNOolaKxWdsqxMGeDShbqXWkeo6FxK+/S77ox1L63xaahxmLkbK9lm3
lFbJpe3hPo+9epm800xKb0Dus8nNoONV0Pp8ktyqgXDeakeEfH+foYMWgGGPYYX9
jz856f8FFJPkfvSlkPbiXHX1DRK7OuXbZKojiPRIt0oqz2fHOZZcr+6zHSNNd048
ANM8U7dVkr85W+yE5uy3lMTCCz400FDUhmiQFtfgJ2ZBcuYnuWH2s6svjzlTUTxL
nMEGwh12CRwxjlbXs66Tk6uz64FD4xipG+UOW4ZSkvBOYbcpml081e08hkNW1C6I
wC3gVoQ5OsHbsoFtF06c6wUtCVBSVpdDLjDrUklH3sMCtq9UfOrnZWk7mdSE9jQ7
Z7dClJlBBe8E8L5PxGCOPl2cPIETvPedyNhxpB7qZLkCO8cl6M3wAEJwhYGbGV1h
EkUaKKSCzZqS4byM0Wlyd3rtIQnWcPCburjHKVO4yAqfptaqgU9nh9/cIQzRkgcc
Zhs4nIS9i2FA1Z9HKNmq81FOSbAiQETRKhXv8HlYMh8LYA92b+32PMEbYHs4z23z
/l8hwdh5yhwiCy5Zx4VGQxBjyHdWyCICWFEm3Cf1OVM9MnQhpCrAeQGzlWcI45Nj
F5KrWWfYZJdNMdYe8Coy01U6RaVDK0TUhXowf0+Q7jzGq1RbAsmTF1xHoeiwFhYp
hyvOgWOjZWLEC73gdOpG+3pCKSkQV9VoUOdJX6EmsRRzDr0+0SiMoioJoD1WI96Z
dDo94u7h4Bww34ZvFcCaCP4DFfnoM34CuQK7oTedHEErEUUMZ/GypU+cVz+zUWNl
AgJwtl1zuTIMlqL/WY4N4kebfuKz4vhipd8cVn+9jQvSm/mLSlMi0+MQlHpLfL/p
4ZTGp2+AyzHPvrRyRotFauW8MCg172OgG4C0E70ggdD7uajK8J2z99JNLAPaqUDl
T1Qudobb3bnuF1GRLkWdSUZm2FYLSZDyCXvAovKUsQGxJgAMScEQuAef0g1Dsr3O
duavBBtxR142oZFpTNI1i+33ahbtweq69Rb5uFeqIsJ7Hk81ggVYrUG+BxI0ERCN
FLzaghArm1/4ZZ4pS5Hb8BAVFo9ytJfg5QXNyK843IrBaoiwAc1w1/UN+PSY/ar3
XuxozykmQbgke4hcJ6LeqWJyExuwIpOprGZELHohunFzt/v0GrHAJS+riZpm/HpK
VMr+A4yPwM3BUhzIiGqwBkucQMp7eJ+rX5FJpiLP6H7v/sxSC+vMmXScjgNN5ciR
FDPRK3zQmdmKUnxzZWXyRLd0/IFM1EYv9aFNRHgHuQ6ryi5UNJj2UXbdri1mqz/p
PgnsHkflZxXjAvS4CRXSCKc8fGSao5Sy2lnvAF6uWjJKtFJBEbohGxd0ZJWhNnbM
KcSs4FWULr6fcJZIz2tTmBvRk+x2Ua4o4oeW5BdohVUCpTkmkgzEmrsZjWUdcB0J
9fkx+rwoddMvX5F5tvlcQAaf2BBVH+LKWQmCVmUABqG6VB9K8PyjT0kTtpjlPc9D
xeHZUkqBFwsWnHlPgXraD8dJK5FqKtkHSns3CDD7JUc381InzfsI3YLs1SEdSlde
XFzv0vihE22+i7KK6AkW5nYqoUHh1XZ4h1aJBVdR2W+q4TBIBrqQ9E0V/p7P/Us8
BG1EAOqn22Ok5drvrjVAEyIt2iD45h/AG9xghmyct+QbwaS59uZDlPU1c6fMSEjU
A7mm8kv/IJYtArGTgCpNlP+B3EWJaDwEu/WQ1NGNm1j7RvpHq1YgQhFU0AqeXsVK
YBVT9Wzz5SrQ5YKXVAUjDRL2YfP7jGtttbDQTdRr1s0L/PsiAUBfiHoJrm2905qm
/u++MjJ31Sj45MG9U+JS88GppwU0ft7vOeFqloejc8msYo/zHCXi+aSPO85zI7Db
XOnBtE83ygpF8UoJRtcInXHwO1pszZW4Sk4/XH1DlAz/j5hfvO34MsdI40HnUFX9
AiAXAE0l9tHKNAim19JKVb23HgOTnsfmFk6bcWruyKuAoOogvnj6sk8ULAEViRHi
AOd5C/kDE0XPuLNi1bFbKCAsLQnVkohDX+TngW5Zg0st/Koib2WW2YNLvhTI0B1y
TUkV3T5JOhJ4+Yf1geQ9qKe33wh/Z+Hj2XU8P9YvV3vq9iXsB/3+eOTgWG6kG6Wc
Fk/3AIKLJCm+NMCRS139ujAsn68AbEoWGraIg3h9h4F8BYUBl0K7jxKIAB+AYkR3
gKjxzKMwiTGH4jWKZTFFByYcduccxaKKIFvGutPulQU7GO2L7c6+Siwd/5vMM+Lm
wDpvBlUAq8g08q5zXSKKOEC3uorln3KpvDeDYdjoGVAU+9DSLAvw/3enodU1redw
jbwIonP6Zke5WkWSv65t9sxvEdKPzkCjcvZ5Uz3+Xy36qL2krSEk9gcMADO5Pmll
bJIyzIJ/H82FO/IBBU0WAcmwfBfD1p+qFjyS82sErXBT/8aNsCG0ttQco1f9xW+8
JETqHSJamv1L+WfzAOGJvsVH725blyk0cjNmLpQbFFk0tKgpGTKMx8vxI8PDGU92
rywL22mHOTpVeEpSvLCIqCvQ1WYg5C7YB6MU2GenRZ2N8p6UONSx/fgg1eRI1Ube
ukFIAzEc1rOBBh8IHXWOdYsVqlyfxALJcbFxdO7jEANc4eFDtBBJEt+NuXAbG2aL
gOJh0SLWuZKEQv/JsXCNgKOao0MkWDua4HwKtyAp8Nr4yM7HrNCRTxDota6PIlxp
69oNmUKxYw0xjir1b/c6hsg/f0Tbkfgy0hi8R6F486GcBgTK0vVApgBppiKOmdtT
byyG/Nb9dRnKkKBIPjm9rRJdOF+1HcUqFDF/hEkytrYPljDlDZk3M/HdhF6RzvBQ
gcx4qYGsRqggbXadPjcAkcLDnLx62oUMwmip5deZp+47x6EUYj+Wv/70gnF2Ttfw
9uBOyzb5f2CdXLzfWrk1GB7xBZiu58fRwQqFOuE2z9Nrabaac0gXE8wPG73vxYRj
dZWlCwXWAdBiq4NEpxzfla5CLng9kCg/O716+SfJmfAWi4PWPg//BDEBaycQ2SKl
D2bNs8FbMlPUqCMrk4b/wbWX7bhzLZFahZfLElItXAxi7oroZmxZu4SvqE+YXZSL
rWvOrDV1bh1iqz6rdnxOhkUD+v7RXb1Y1KX0dXU+O3+xoPgYrPGNdmUamsxIgCeB
o6pdhyce6PeFIzaMzgvzb/xlU/m9l0bVEzpIHuiJdTmlFbk6aRjgA9N/84zxS/1L
uOjebjMynRL4Rv2q1mKwZNW5DMiDCJFZyF6G92U6exrN6VB+s3uOLv+MLXCfPpNP
Z6wEv+mtN585wqk3qbMrBGoJ6gKM6YL1NYfdn9XGdMvTT9MY9lH5OpO1ptngiSvw
RTwDw2vivETb85gUMlgaQa4bmSAo6PNA2HGLQGbygyrkxiVIE4fp5KrFqs8J+SZi
f/or9qZkAIRtsvwp8vnoeyGnsLv4BJJAxvZadgjUFZXl9GZWZ/XLt5z/D84X96c/
aRJ9iir1a3jPiJNDTHAM4ia4u07WNG0SqotP1vq+CWK1peeIJsUzTdhGISnsodmv
Jl/yquXF18jvR3ncFOmHXphNyU8d9Ho8R7YKuIP34CgKUyZwEwt26SZRHRYtIjua
mNijdAtiISrt41WI/8X6rgrkuOGe75hZoBBtxEnshnxFJFbZCAzlhvrAYxeJniuc
OxvAbANyBrZQNmzb1t6Rhre8GIH+H3BjJf8gUhZilyUIdtikaLFpAln6UerCkezn
o9uLCVE2m+Su9rijWrJy61huUEssvD/GPhnCyQXqm25OEtX+U2g1T0LBW7FNGfKV
BiIBWs4QtZCml4Me6rRjDczLObkowlFEAiKKnqt0/Xmy93D5lrLcMDPaHo5L2Zwe
cxkkO5QqTeTIDKwzLgtsSX1IEBu8KNIcHdxaYNUdRXiwYTAT/oyt0xNuNZFrnG2F
AVHBS0Z23QncGyVlO+BHZcUHypULvi673GmEr6ih/IkP3RybBvf+7vuDuYBtDGAb
YwjTi2L/Eao6zZTUjz5bd0hgXUU4Bip5qAKp58yFiIQj15BihTKs2JyqKcce2rs4
Xutw4K9DQgdiAIq8b0jexo3XsjkH8R+5yVVkgnPeZetY1JRz4X3Fachmfw/SdqV4
+Qpr+yoGG09DQ4LPv02yPC9BXaxmcxJYe908+NYr20EMVkOJzqQ6BjWxE5C5Ekg5
hSsZfR4nTmQfRMC2zrQryR/yNMoifmGE9UpkUKYAKjZm2oB+PXhnh8Q1kXl2tW+U
cYW3jFsiQBKh2KNedftxzHzoAUQOvZKwga8+G29rM8RUV4qH+PjHBr94YHFp+Crp
DGxYQm98nX5ExjbCLU7ql4BDPzDm/0Z6eL6L41Ou05yN+t5Br4xifSAzUohuQ6r6
VspWK918CRePuJ57/Vvb8G8wnpZJhcHX5ydewGATN7mDtpJ5JguaeCb2fNDjXCuX
+qzHPDNFgXkFgWhBWXvZRL7KfihT8AoX3aQnU+Q1lVi8X3mFQE+Ni07DMh172UAr
TJNTyb+N+AbV54fDYYJQWwNS5zdmY/aYVg7Q5ynoR91oBD7FCzOR6LF0/SWxRCVX
f/TTDP8XNhGlKXm9RbDs1Eww6ffJo5FB9AVNu1XMx8NdGMynxy8zo3NdmnqR+Ez9
VQLNYVf2Zx+09LCTZMzi7rdMMd9kN5pYHgiDEukHtBTNJn37/l0qVBatgVAPerXr
mp/fhbLJRHdhh2+s2aDxIlUQAtmIuL4q4/xuzbsj2b09nPXqVLRNpemYY4AITnm6
GGZAPkdX1tfNcUKCLDjzQG+k7d8/bDafYmHsxIG7goVyt3i5eX7hE8BXFOeUN+li
CUq6+WC7P/dhx0QprJC7yg2Op4MhVV9NHpce0X69Iov7kmbSdEk6QRb/YVgKGlDp
DpwMvBvYVAAOEXmVv56I6W9mPiwuAfZN5/TE1lrMHpZQzuPCkwzvKhOqBwJ458Bb
F1zRfsgNsu2oc2kvitvi17vw/f2r1Dheaq12YImtoOSJQo1BrYbV3669hfevA23f
WSWr1Js+e/bhiADh1EHqA6b/yavlp4i437w7G+uYidvjAoks1tzHDr72SzY4i7ky
WP39erEXlu+L4SjdEqMAX5zia6IyekOix8zMO4l69xZsxrMZkI2l3EKUE0cY7nV/
XRj/59E3igPGBQ9ZQKeA3FrunfWNzDEUkxkEI5TwvaoCw0ml7qeYN/joCtycFlZi
0x7a476z4BpoeFy1bvWa6s1Dojvx1rtON6pwnPMIbrAps6QcejHXzfBUo2yWia8z
99i9N+xb8VZzrX84ccZzkECboMmDOIdnOHu6ya9cvRbglvXWAI1d0ocyhl6THogv
Nkhmdi2cLZ+vrx2rBWybrVEAK/ZtYet70LktRoFfp/CTceaDJXuPOf0Dm4fCcl/O
hRrGM5br1y/kJOGkjVNkj49wRr3gxkv+CwQwc8qvAd+ltN6OM3Wh+3LI4wDil0O3
dkhmwzDkW3Ysm7zwGunVQ9VHqkhshtr8MJMsdjabHOR9keh7UrNBxYN5AXW3e+rU
1ZTmIqgXMHi8Qp+AJI1u9PpBegqXjxI0OFOxsksLJi718Vb+BHfSbpdZ2/r/Z5F3
7QgkR9L2Bjzj8HUDxKzvVCi2RkTuOmlmpf1oP19ZsCTylZbVFeyFpd6e6QDSdIMS
w0Q3sGG2Qe/yb9i/SOO8elJuCXsdFU82rVDSiiQ4c2QIoDuguCqsk+nGpl8p4zFW
/rq//jkd5v3plfhocAAcAjuvRY/5XMTqNvw9Z5D1NCWpVnl6pwEGZ6MwJ1JHk5c5
rr2QHJ7Oa/PaIwaYpy86HSIj/3gJGLKzycn8zGGwDt1ZPyjCxHQ4k/oNvVQexI5I
FTQFRyLkCW/6nSjT9tW6S2cPQIA4rSVRBBXHeE81td/7rAVmt2xMUt0B2jrXabJB
6uz4UF8iVfhPS7SgdtmMnb5UZxictgXOSDkFdvBs3IKyoJEdRiYi2aOgUErO2gUb
X5gz5SNhPNybGZqSMxUGhfUFl1dSFf8ElkyhGNL0RzXvnROePDyY4c5OsI0I6i+d
11X4TGyz+GmLfsU2rnpnYKrFqjG1vZPOfoMaX1Nr5FNzuCL4EvzWsXXdsp0x7uuC
fDQO6BiDbc+5LuiGR3HOsNGXeOB7/UCOT9R5ECaKopcCfwErTE4juBX6U60N1F2V
90nz/tcWOwvKI6cRLDTm9otTjrgoip2JK2d2CXhrF8VvJLzBudKn/0gNSfwwJidw
od+k8XjxihwnlxBl5s8NOcKOxMRXHf0jNDNl4iIoMYnPsM0kf6/lRvtu5sBKDVjv
ocRiQFs1JQBHn7qdDKPSnxKp+lyDXHyNUev+trDR2l7QWQaLVZ+i4PM6yoaVY3na
P9/JxC+vq9Ve8uMN2clRjLjx5xW16nS2jx3Ye3f5rY5x6Z58XKOESHzocT3IqYuB
BnsrNBguWnrO2DZ+nsR9cykb9qCRQgMytyAU46uzalvNLwlRJusS9hYu0KUMP2lU
xUC85A5a6gWLIsmPCBos2On+YR6tu7BVc0ERJC2qZt9BkUyvc/r21L+xjgBAQsgS
VwIGA7ppVuxHsHcmZcmOdlEA21JwEtGDIBSEQgIpiur0eFliw8Fk3P53NkoYGH1a
D4qCOqbWFzvRxAuHLcnt3+wrBmP0L8eii8ksp2e7Zsjqt4rHCkdRazlFQNV/nD1j
AI+vwfHQy7+2a9xlnQo6gZqQ5CCREYs5e8k1CateoXUDUR0XRsVJvWtTw6+uEwLD
eI7lqaIz4ncZuSRIyK1Mf/PSuzamxRqJ5okN2zcJkrRwFB3rTXsmxNazrQHhdJWI
e8G+j8Wbg9H+Hta00lS1bRJJkj0lINb3FID4f2+dFFHxpS71SAp5ywCvHtt77hC7
7HBDCgAAXYAqbZbX5CHxraCWayJ4B9FRlEz6QUajjdTwzXQkjZrUtM6dtIeFfn+D
M8pDeX/C/YCgMLPOx0Je1gxxIYx1hkZFqqbLZnQz5YmBxbnIeRUYvg1icXRNF88q
mX8pb/MmZFqZTaHVFn7JxztFhBWL8DmkP1sc88/yzS+Kf+Ue2M3BJDI0u1x6G5P0
ffqDL16k72YMV79BKBU5tzNsQHOct9mRYfEFKiLv2Hj54NOxJUMdqAZdytbyYiWD
T56f/hBim/GP5FLL91+WwifgyHgzwqVZy8z54xJilGEP/MQzFIYaZdDE7xM/ID4L
1PetnBPmOPCjMBbACBBGuP7vjQFb2Z8/ouPqoBpHJb09PTwPPLmhELW04DHa7Wsu
l42vVAQHhiZU7R7eSVcUuHYo2sTPQ6SsG6k/grCbg7ApeEfq9y7PPMSWwhoI7KvW
JC/+aY8QMGcB75O/SMTj245wMuqoCa469TbdPgGe1YEyu6kIpKY08OdJiWkS6eZ5
YJbj2LDpS9CYiuX5T1fRt1SjT6Wfbt5qGIYyPD+VvAcHIW558n4/MbYxyhMuA/BF
6DuLNrGcsr7X5mY79XGgS9IAt/941kfwfxdVpWQ9qXSaUnzEZfX8fq89TKjOkxCM
S1nBaTpbUF5NoUibbZ7gx7rnxJwg8ce2ipa0K7jlgvJCWvM12jUCOciH+3K9iNzh
v8ZxxyiTLGpu2TZshDYeKwOjlIgiW8L03GkIHpx4hK2cKbUKBaweVh+Zuw1ppS9p
rv+ewOxj/jM9duKOnOWYsChFtzA7s32ofLoFGABeg6AzLwM2b3UujE1geY91drjZ
Chj9jFpN4UQsY/g+t6AQXpGYxGoP6/8sb3mEni9kMisGmCrxXGi4jprnmZNskh9B
egiU/8EkAUweSN5u0JrOLHndtJgbOZDBkMreazFg/5fSM88WcKm1sAwM//ggeU7S
4Gmn3AbwAISCMmawdjuFrr6ju624cIOqWLsYooUKPGWANV34p7uEXDA6VyXWp+v0
wHp1Y0aJPrKPIcLxQI/ukQXbhn0NH2j1kysIY0p2GCOa7MQLh2yNePv5jAoWDpBW
9BLmwkB3TvgsmNbGsHK/eZkWObfq5fTtSjSPDE3uq9fExMqrzVyF6INnYZ0MlMAX
40qxVj7MegXfkmGKPYW9/4aCG9mA50xKyBT9AjcWvGNSQznndli63vL5SaANuKKz
b0A2TTPLLH42BVEkd9TStABy2mAWE8YZpLn2/BZaqrdwEU3mqtXNQ6a8ymhnYjlx
Jv0WON/c7Ftau60AedytFRBJR3GpWZBF3nLEBNXmiUe+tGxiu7x5YVNm2y98DVL9
or1DjGj8NFMuA71dw8zLr2ShtYbPPZvjtfjPvUl9zJEOqS0NhASdL2Tr3jF2a3/9
kC1m1tcL6H0mVLqJVl/xwyMN4UvdtFQ1Z+JW61lP1uUGFpFzQ6Aqhcs7T2Vglkbk
d/BKE3jWckn2SCo2btls5QENmqbXtWKHC83rSsn/u/WFsCgJ08fEtAF4DRUh4MUE
XkTSxh6wM/IYNgwtogFVKOeCp9hv8h4KCKQux8+3EL8AyiwHrllWbzNU5XLXuTsN
UW9vDyqwAX03N7dTHXF2C9qfkOj127vNYLJ3mVwa2KNWHFnF4nw3TwmAoiOoR8vU
dKaVslyZTL9oOHwDO9wTFD3kgFGORyylGTPru1MbrkVOqTOGPqEQpUvZs0HwDC6U
6K1/3QvApfoFT5JACLr46i+GfDBl7M9AseIR0zHL5cMEmgfCZ0M/kggqNfxd8gYr
vDtwM7PYOCAjHqydpabEyLKvSxh9QW2Id+1vR5honhjrwWqz5ixBhiJzh7RXpI09
1KMXaA1lUUXsoZiIRPV0uPvQ4sffE5xlRJNK/U566ZNnazEogqFuICkmly/QFSL9
Rey/ANgiK4ITco+M6iqniuB0KW6wOR8Ma+UUD3HzRvwPGVX9yVpT8NEqGp+l3192
WdwNnkwJ7gQQkPt9UIw8WklGe4mhKHLJqwJU2WfmhXsXVnMzmIevvNPQiSDf+ZYJ
yYm6jIEYM4POLGIw5f0eo4b5VR48lDU9WdHUEB7ok/lbTWqTZDV5akxG/0YT2G/V
uLGVdq8VQ5DAsVkqnVPDPKDocgcA/JmarNbDpasI2fu5n2bxU2N38FBOKzNr6Yyq
TTLkcBW28/79x/tNC5OyBb2UAXFnzGCvuQgSmMllXNDcU65kn1ouq8toZwOVp/Lj
ybANTn7HG4esxE0o1dCpE1utR4uRaCbgNfS+FvpsAy6LMFxczd9QlTSwtWCAV/Ys
27t4uMDDfdQ/JVJphLQwWJ87k1PHSs9m+9CcPxWtOz8pZcWnk9WIOebjHpiCa0Nl
1gTPMpyCll5NT6Iuw+6vPneuomjzyqWrh09vLNrTZIhEuw3YPe9l7j/GvHbqE8Yj
WpPeZpoxL5v2WyxeJPE940fS9fzsO07MTMo9Ws3RM8kgpJrsvhlipkbPa0T8qDQR
pmAmBJIm+CPEKsWix16iGtEO+rV9rE1F1rk8MI++FRHh/XuEkgrhcn0RnDluwbYv
Mh1hghgpo9F8m7q5f3cHxueBuhRTFNfFcZ+nB9Qr9p5goCqcD+YhPGtsrydoV00j
xzApvBcfvO4+rTu6k1w9lEVTwu1qqQwOtbCOcSBFHL6ab6kGT39rI8BNMCU9sxrm
e/M921h1MNJLKUuQ3Ys8R55udtU0NL8kcNj+Oo7bO0oSfpuL2BO5th9315UyZfy1
D5otVhmSCHcood0MGLDB09OskiM0vvOfEiDzF+tU52tgHD09tq6IwfjL1G1MkXub
3iQIzgzX8KtTF2V6/4bS0SPZYh44qsg14PAWU8AqJ9W76dcOmJZzriE5NVKs9U3a
dEJfwAgU6LWOX6J9n3a14bqhxSi7Wh68vHlO4XuiolCTobPNfp9k+j6eSSX7vzC6
hYTH6CDY/Jx1ZgGHOdNxPsc9U6ZcfLrs3NXOpYJVqogryOnpJGNdsEgemlv+LfNc
hAeki5u+pBbJ9MRvbSJy3qXuqLrDeoKif3AY3jKu5NC7k/fPymfB81lJobMZHTbW
v/mkfj7oIevd1b2Dmxbo+q2EVKrGBPXzdFb9TWpyGnYdomHJ0o0DnWBOVc1Kpfwc
C+UfFbpe0uMHTVFRqUmoWM9xIV16HnlyMCfZ2l1aXRJE7/vCLT62F/HbScycOOgG
VpBUg8hPDTXHAG2MFCJY2ZPphWdGikqo+5FtJVvo+nWDMsNoDzJo3hgYHHzdkeBZ
/M10AhD1C4VXjW4HEvLsGF1NAD9KPmBmQqm6ov4vSeFR+v9/pNDpw/WROgNlbHTS
9HozjAO/NRFF/4nBWoZEqMTLWTNUJFmS7jiFelHorf93wc2wE7xsVYzYSIePG2Hm
n0nevfe0iDn1bUH2Z6M0nycI20ujuXtvYvnZSCmq4FRDdV3nlipN6eGOQxCsmCWm
QzZdGD6u2yHA+JHVb/z2Zg/+fKU3AxlPzmJ4gVET0K3K3Z8RSRGWa6A1qwVaTmlY
fsjuqFcGjIzmNTFTSSr1m3ZbnS5i63qqkORfuazh0ZEUJzflOYdV1E1saFpWz/TQ
afuihLS0f1Ax1o5vvb1gp0rbWvzEDEeEZHn6ZeuQBFMyYMAx4J+3BtHCJt1ifug8
zIb+LZZmEC78C5yPNGlggBtNwJdXE5O50EpEBcFrQTPUe/A+/+dwbGHk28Dpx2Wn
pk3rS3OtVuXVe4gOsAFhe1EHB7YHvefJfjfJjRvx3JO0WfqsvPZ/GWBO2IzSS3RT
3Br6f55tNfgIcMOOlaSB3HRltsOmIMi4Eiggf2MibP40kYKtBUIBoS992S+2aTvX
2uc9qyGpLjqz5fBKNgU+si92CzOSGv3DK08C+MV249b3yyH2d1R5WTwp2KiAj8oa
LKaaZqyFhVH9Y5wtmC7I5saOMdfy/G1gqTQZJy0jsWhyQvY19KUjnWiRY5ePn3Ti
MYyx7KOp8wKDr7g7Jw4ocXf3qtyAxGrGyu4MZcg3bcylEig3IRBWRtUzg/hfTAZk
V48+nM9O5ipC72SAa9jPjARfNPiHTbEkfXDKMIUa0S3l/+PGqigYVgN1fwXMSk6k
T+/wXku0b8axLSDKToCo5iBi1w9nrag2nHlUP99S1+wz7sVBqDsESTn+3WDoZwX+
U8K9UIq5bcs1CdNuLOH2FgLAgN4nykb5y60pAfiK3OvAmF0b7v2ctqlSrKou2/ML
XQ0HMmAmOLchreDV6q71dhQqpJECeedviELIj/Zy9xXozM3GLSJp91vBSZ1s3zLW
beutEsD/F71WwRlV0v26fMr+RDOqyupAFRsHUbt88Y7J2UZsqA/dZ3mQb8Et7r87
IFaPi2P3EbTJ19u4R/i1HqK3jlq2ssFRIYYDY5DQ7+loDjq5Ss0kyX6PFMMr1PIm
0nwY/DQ5Aqguy3UIAXN8OhQNZqYmGOVdjcN0JFLq/sRr+I6b1qYM0VjaHfs/GOFz
rG2qoTbFYF6g7Fq1FoaYqvV+7CthN1YdoRzhEQEHHVZ48oTAuivGqw0hu5Z0bndQ
CNquGannzqYkcb8PER/TLekFQIDI+S8DWplNM5NYK904HdQzc9bGq8LzTqTNLcyR
RLhoYE3b/N4dbIpM4HCY6Yatf98xOubGSEYwFu8MuVNKAMnJI8jy5c6+Uc5rqoUR
OBOXcrHopSLXXm5FG1T3vRIrNIpLAUHD0Smc3NES78zOAR90ci90G9I0MBeRkD5T
FQW18yn6XTa4Qw291kKWAY1rjU/Ubtm3hlKquQqFt/VQD2VbUmD+xaH0qcox9bok
Ks7wP6+5jZVHSZEDWn3/oklFj8Rt3nXOE85FBxFc33l9SfTy4CXkeR45IWe8aAR2
8vvbCiKBuyOtoMRTAx/Dx9u9Fi1naFYUjz7cZ2EKTQLnMBv+rcz2vVE9GJ3ZT+eH
Zim2swRmSbmdthoggGO4VJVrdHv8oaNhcR25LRyq2T2cvLpmcIeSHZ0ojvXaoW4m
VBfen8kP++YzCaiNSp1eEhkacVyWS12pOQnR78xEHqFr3fQVlyPm8+FykVBn2TeJ
DBAnbp1JD3tk0LmXpZ5asI5n2NrOCwwPE4coxpRMzLnGFJ/IjfaSj9Hqu+HKfzRP
t2roMpfIUPSL8Hc5GoJmG+y0UdxpLegHZjNO9WoDkdWjvGZagBVnwBhQsQ5qH2oo
GN/CVgaj+GGX9oAJWiw8UfdVvWHUuNjV8QWAcGy2pMd3+fwrwDWAjK5CPCLNetfD
40pNfbZxZr8h4nHwQi53oR6FP5jv/K27PRkvJuVVT/BHYvrkiR7k+C80zmpM/a8b
ToOIkdvupWR9pmU4Lg8+/+27/jpkt8vz4U7wPrqISWhdhzkG/NVq9ja3ZifQXDyz
kDEIxmE6vs894OnCgabvHUHstgjNyqUEYL6It+Nv2S48aMQ9VWlVN3SkgdOSDIgb
f4L8thwqcgss933HxaRTtBknP+WKumFMpVjw51cV9A0uqAOI79mb/nhrD1oS6V+4
J6W1pNRe3ZnkqZIpdZdF1dPsgBQ26Ke4G3J9B+9NRuJNhLImlcbyXi1eqhI6EW78
tY4Qn7C3JRYorexiGO5cm05qSKoIiGqWmquAlLmH3Vzayg+lcO6Ba1vt2oCtm7tp
snEPkZYHnJM2gvzHtR7MefAhr25RI6zr85vtm0YYLu7NOJfzq6r+bKqT3h3hO7OK
jBEgNTKglITStFrXEMVJwiiys1p8ZSIMSmi/Z4ExoMbzeiw4VIa7Y2dfOQqhmQph
rqOLmRYqgi1nfCMIac/6aqYrSrZajVFKcry4rlVSDH3t0fFkM6e3jMahRXLeA56S
pquFFe9Pdn1gdXR9Gb7IzXKpN1qyubpZXz0CmfI9dgYGiRBFeG5T5GaMcdagzB9U
Gm4ilSQVx+VZkkA8UvFJ5Nkg4zf6xWOV1DEBRFpRgdOoAgBb5/1IxLnBJWQwfrLH
jXWj/BUNs4+3/nd6H5N2/53LlvcrR6DMHPl6b5pyO3myTWRMROkAP/DlDsJ9+3tZ
RY0egC04xZ1SuQ5/b0WPGXcprrP38L61aLJe88Kb2c/CSF7LLRPEkT7kM2rU2EL6
Ni+ATZUKCwoSZ5Q14Y3fe3OkzP6sf0hNfUSRNI+t8Vf7CEqbMoH8qx1XJ6LuDo4n
lw+rbdWFclcXhssgIEHA4TfsiqFEdhutet3Q8jYi2yLH5KfvsCGLMP/D3iMFka9v
o76boDlMDg11TM8L6wgl8keXy+h3Sbt2KcnZAh/nRsSQekoR27OTytBisuB3OSgj
ljVEc9FkO2Wpxvpn+pNdcw09wDEsXnLfr+fh+7tvwLeagf3pGPtI0McVC1UM2kNO
v1HoOB38JACiaIlMFvJWWs+uGfLVwFvOU+ZKQdiu0fyoPHiJa37+WbH0ScTTEK7j
GmtSWzzzofCfDjPYXN0AM10Z/EZvQqriEoEfLKQJEDmwwH+hiR9+kmRhEdcZbnj2
DxNLQnwvoTEPp52alM6iQB2ltlbr3j0P3oRTkhCdiMqJVEKbqjntFjGQ2tNonCw1
SP2EMKyNMzmZaL+ak0gXwEZt1/pUKWwRdeDsXNkwNagOfFskeoeh1ePIp0teWzdw
PnrVoxeXcR2765T3cH8LY4DQsMh+1Y7lBtCfiiFBtysOyrou3GUOJrsL96crBG99
ISnbSIENSK5hYM2AnPp6Ax6U3wakyxCPHyX1Fq+wXiU1nEW+mxOkuqO4G4zmv/EQ
9bS86AmmYMIzWlhY7/L+pHdzZ/WEHjKoi4IL+5/FQuBW/79wkU4ivgXetcTcPkfl
jexC71ftbbezu+wzxqGJZ9r0xAwwkHAhgwOOKoKhibtEiQo0PAyMTX9j7NTe6LXq
tUGj3m1O74BhbGLtwPOqgk0bVt32OxXT6iv0m8kcWWdQ/upsXDiAMNhJk09PPPv/
c6xsNOfhxNOS9jvi/gyUeVz89G6L5cq3FjL/7gBGHkBc5bdyskI2gUMjbpVkLktO
Ff1xqLRYBWpZkokPyPxdt5tDZgeNQVgaqxHRQMVehIjTmU/jt4G6fA1nlUrjtVpr
q04+x5eJ93m1MSZ4QRgIPHU6XHMYLRQdn/zBV5pdKH5ZUeMA1F5G+jjZ64clM5bB
FlRBA7FVmi2PrBNd1Zh8+eD4rBYDA7crs+zLcd/UyuW3TBFwi6ebCxqYiTd+w6zF
k+iPY+aYaZDBjciZCScqfqHfyRFTsAaAiB2R66dywYwsWF02eGWTQ39+XzAWnJcZ
aftMeL+Cg32mfaB8XaHXrLMo/2ONc0ArO2VKU6rMMylnf5FKZzrWBpnVwQeNMRha
oGIoJMi33rjyhDLufYxYEWHln3U7QmSM+MPHFF5jsgCDWAwpBjS8ncgbwFhKoBqR
sZJkXewZYppHYs2xCeQQO9hGPEkBUb314adIXXry7AYxZ2y4nODnAO/D/trt3E8q
ipfLEBlZh41fy4ShWmf34E9WIx2EK0XG9hcsoSx1HNVCxMhaA7TbGUf2YvwcTOva
IvCYPbnmJ+cN2a0smJlGcHRZCJc7lRMtEXGEG5nb0e93SzfB4MJ6MaigsV7bQCK9
DiRhoEIixWBCyDiLkaeSR0K6NjhOjHcnJffy54Pg+LfqcVuOmyOLvyiPlSNSMA0e
IE0KanNk4A4UtUGXjJPIj3/Izy6X9go8qWekLAMydCs0nuoOTLDfwc5hoU6BBrws
0iIIrA9+YXXIOG7qT/FX0DTIrkvy8H8rCV4W7WKaOfipuRB4g86yTEzVQeTd3I26
r0Qfi+G9YLlz+FimEs7XrYWA301oifMp9C+8td67blusfXdq0luJDGXNIwpQhK8K
ZAt4QlIlY/Nd4J5yILFZA0d+HfmgeBsX/qwg1D5EN5BzDE5hj/BrF2UkhmGQ9uXU
m/eFP4GebI4pSMjvc79T12Qxdj7BLAm0V28U13CQRi6knj27wyy0Vs8X4NLDlvnS
oPHle5LyN2YBRFvYbVCM4y/ir5aaS+BqVi+jIK0W3FL3CiE6j8mJAhB7xS1Z7s1q
MMs7qQeeF5FzgVIMKsCXipoiuY/EUHU36WZ2udC4tgUrR2Gq6DQHBDPqEF/4x8Lu
JKmhken4KVT4nxbukknYctHO8htCwIrHN2rCWI9Ac847vIChnCaw3iafAKQuyMYM
pFMmvFrTHb7tq2HZ/RFieaYjvhx/HONkMMDYhZQ6Z92DgjCcdDfSxVoEr19gNvXG
5foV2WdRQ8iIuK4DaH7TCYjGUydzrGzJcu8C9+P0+YzZM9p/vNf7NhGZ0zZ8CWaL
b9miLR8TPcc4Fa62l1BVbfbZKrcNOnJQeqbn3tU0H5zRm3oaMBYS9Yv4X3r/aaPd
148dMAp/vy0evYA5lSHv+xW9D287bGEzyVq+rPfnO7Ns0axoKXJDhAILd+wRna1t
coL3yKHJn4sM8U+bt0lth1yMMGHBhVwBLOhiW1lp6mpY1m+5Em3iPC0aAcHkZX+R
vB0X4Qsa4yUpFEZyLMQMTtTNOWxaS+BtsvKida2vLhB1kMpz/ehqDpqxmtMgKWcG
Xxfaksl3CQPcgDfOpdRGyEs6VjOPCqTVFUq2ukZN0KKt8EyRGis+cJNo8S08mEuC
nD/6XhmZ9gBFogAN+cWLdHCOXpGka3uNJFu0k6qyLqRw9sb4gf1OswjGhYTgLebo
j3Gl2ymOTAzcJJfc8c2Sgpusz9RXYGGuyEx7bBKW08k7EAnOsPQTMLJgtqJnZ1/s
Qb3e+JUyU6VncVZ1SfKM+ppKCCRwZ3oirLuk0rIQlZRWQlJDy/4n2MCDoZWgSk+0
P3Vv4spi7HIDhx8PZFY6iW5BIso2kWWkNAjYczEJ77w8XBqU5SRK6mb1eLfKVQZb
OrE7AVBMSZLUQ1o8j789Ey9d5sdvWjVP6nqIC4kldUtRloz05BpzCIOyWFlWTokJ
zBNoLfSNan5r1ISBjaLvaEugqfqc3h8UHJID91CUSB6GMIJyNE9QNQNSmDFhSQ4t
V08Y0lqvA/VqA19Re/GoL9sPYIfzpBvIBfU6hL+8b2wq3OjScAF3bbu48MqFOviz
XxcUuuI1z3zVPzwu9dRezyYoW7aY0BhMR4vfg82CWUtUNfcdzelcksKfRYDjJLAd
IbLkST7S4Go1qf1Te3cmLvIFbI6N2z5HK50ga0M6FphFHfy6hVZ2tlJ+0tANN8ka
WBvaQHwxgvPCkuRkCiJaSSYxWD34WEPbM6CrAqRvyIrf9hn3d9HS5Hwkb2FE3t44
pYUscDcxsjHKXd2bR/FhmRrjRKIQfcEYoc65vHId9+g0QWorWNqKK2/MWxiWwNR9
w8W8i/WcWDOIhsjz2t3E8MftCCTSr7tPbg87bwueBs9fSXbzSkOv4cZ+kHx2A+6q
fbvI96MOAl76LAsP3FGH/6AoX7SG43A9siGbB6Z8aQOhF6KS1jKL7xsMuN6cb+Bz
bhfYEcc8zdrAf0hMXPkhOVt+3wikAHqb6QDYN2x8VEhFUKzh7vuBUCXRwumkqKnu
duzImj6JN5iHRhYWNPLVZwLZV2t7qcv0KbGwZ8UfPC1PDaAdNTr2zV7W48a57OhY
zJrtZPEJZp30+LMchxHd2zLzrbljJWjkQoJOYQI1mIK97ZKRA8/5FEey0uAQ06hp
bqXOTnfD4JkbVC3V4TLpz/TLA+0ku7GwjiQcS/Cveolt2jRXj07fBwFk1V3q63VS
nvrr6H6/wBcNfQMAebncWM6tCY2z6XYUDH2I+wgjIszzSIXF6ghQ0GorBQ7wzPPO
M9gynZty7dWEm1Kq5YPAOn2TuYjFKz31kws81Iv/NtyCvmKU7eRpmgiqmgR0+lwU
Tuy892Si+KnTiQX2Crrjib4DcGxCWnT6dwVJ1eJdjDGmyDaK+DSkzssvO/TtVTSi
2MWzFyY9fFORDmlmXa785H2SPbPW1+oz4SRYxOkbhkDNsXLLxh7n8RrgJOfSqk5H
NkLOnH93kdt2dRpRIqPfE6r2ke8dgZW9Qo+fVRCOUTQ6GocA8w8plh8rartwYjMC
ov48o7POKK9n2IoupndUPF1qGqcDFRCdIAqBrZkUpi12+Uy5MxHJ/+k1TPtl+pQ1
F0gx82HiADIHeVWp513b1bc8SfIJxfQmpZuKLGrGQWD8xefmX3OeOjRWXH7/tGf+
wZWmT/A86s/Lpa38zW5kER5zhmNrkFtkjxsmidnbEzmtqpUvhEwH0j5DNpV59yTQ
+x83VzlZ9WdNErDP2qmaiNuYR7zoG8erN6v7cJsT3nbcHySa2RSCP9okcl5UuALW
BVIfKXJPz67hhGlfbDiqaqccb8WX88/PsVETV35B07oY1icSHu2DEIZHnxltGWiZ
WbhMpKejmoUZkqgxYyifVEqqsXA6Is05ZvFjPYRTqGcmlKO4/D35+SZ+QwBZJ98t
BH7LS7c61q3c3bZFHpjx9zaBYRpcyXI90v6yd3U/i4omIMIO/oNSwryye7LGwHiz
7Q4d8ugGF4kJI7YN9RFVnm9TfVL4q/c55B+pJ0v0rDwtEFkpwngZ+MizSr9Hpbht
LIFo277C/jcIskqTTtxpaCTokqxf/nBh84s+g8U3K0gzqzzyiWVpIY3Iz7T211WM
7dsUksuRzn+eTrYfvt2VzKcAPz/XR57ywLH+Tq+q48+e1Jed3wf8zipn8J36Nsll
zef1uKaNgk9TEmoQuWcIjpEeTDUxxz7OTRKY1Ltpj2Sc4Fcf7E16LTp7WYTa4lsj
XnIDrk+AUKwj37u57GtWzjJiTqbDHfH20erQMI2efOK3eqCxgSeeN20+iaTNwkUL
pTDirgv5MoT0zBfom4u219gXuKp2NDx3aOnCutstgmu9phKXFE4WImQ3zS0zbPLr
a/RBvDbWWHhtaxrv/F/3NqQ3QL05gpXRuPQjJ2yR39+mYXauus6o6WioSgENBTpN
SN7OFufidu+E17bw46JG9HucOR+51XUkCy2Jq/HRgUlIS+DfA1RL0lbN8S96lncv
JkRH7SxGxcB0Tlm647L8/2d+WxOwfEeStlwHreKjyRntRfLzyq7mL9BNPP90wLQT
pZ+y3+7KLrWKGG6OiCshXEPXRZLSAxFBnR+SThykId9PhdRWA7ZJcghX2yH0xbYn
LEtmeuAYN6sGo7+PwOgYOsw8SXmg+ljSZ/dIBNzQXIbz9W8NlabiOREPisid2hhd
C05THU7rBMzvsEAitDso1H8y30JxjJii9MHlnbCPPwJ3WjN8UYU4rPcym3aXwPN1
aw6mKyc0h67GG42/TqBxVzg8ICv0ik6BHfWtA9xPqSFivTXxXzVj5XzkWeHtOnuY
fO80baAPpAixt1YqusQcQpyzwCr/rQ37nqHGEAVhaPpwalov7h6TCrd23KmZBnOh
FTU5UpqqOjOlwYhZ6ssh+L3nPXXKxaBeRTxBLHb2Dvnz0kBsw9o2sk/4ooHX17iv
DSDVPIAINNER4Y+hDYEPoSQZtQqaLAm8UfD6K9lwDQSenIK4dKUKlXO1zyJK/6i4
nya7LNHTkUWIV4p3DEUwLwOGGRYMT+aIVnWOOwvMT1TZy4knbojmAJtaS30DHSPX
J9S7N9FeTb3qxYuRmY+sywMu5GBty+xK9Mei53GJAp4rev/HJuLKTdqOnNiWIwK2
NC2xEc+OTJetAMaJNOLbv/ptNygsqrSXaWj8aiR5b4ggT+XkAg+XeOIhwYaMpEUF
MRhfe1FDUBPQrJOm80vZTGnk1h0oHNH1+8D2vqgTExWh8dW1hYeS7meeuQFwJp7P
EkEXXBD7sEbGkj/xpXD2RVlri9TvtkfgA7OtA9fMOecdc053f1naBnqwTblfVHch
j8vagmvP9Ysb2uo+oZddc0tuNRjYBDSE5tETkGsylb45ynVVVzUmeZqkXR0RE56D
dRDGeKtulfnyxrs5jXbpVW2XsNm51agwofkDqWoWyGd3s5/P45S9MkN++zeOi0zD
9+2YksbPyCfxUBovPBljtQDijrM8HoLZ8DsUD+KsK2hCiANkXcfv9NjH6dDhWP3C
62sgAvZw4fM4tAI1D4Y2CknMkPyt5y4bLx6DlBz9zCaCdqhYy207np3CeD3WFJNU
evbE3E3GfaaiQgcA4zk15K8MC3cptn28fjYeYnTkTlIPJY6w0TUiovo4vJJMeyGY
4WTDQWgyZJOvhBvDi55XDe+9cibnEfybbhXqonU5DLrFM28YRYfKxIbWsxZQvDLg
CcX6am5Pzd0R2+edXQhY7/GOz9JJ78xo8K8DGJdq4qdbJCM9cv/Pg8cMedoypDC7
66+t7YT4gaz0PwlGv+okL4l9kftvo3UujdDAkEj/6qGLYQ7aJJNmooicFui+lwTO
rMZCqsAAOyqnvIijYBtu4s/sbHGgV0XF+Q72TxbYaxueIyaf+szRuXdNwNozYdTq
ou4Ut+tjaU6pMcaIH/+SsIaSYY+GyrYKD/6854apNkhKlJ/XxbHiA9hfI0o4opH7
bh9XRXlJn4I0Wy8dDh+uwjMtUa5zcKMaVMf4pCpgjs3mGSxf9zb/AM3znlkjVgiy
zIRubLjkaCy8HBNhTfWbbSQTZRxi1nZ79Ij1idc05SYYeIqAToW7EnqB8KAIQIEr
pq6NiivGVp4SgdHVIpmDdmxGP6v6a4wVfgorzlkMkgypfTwHorIQwaBTDUUlk4oe
id9lC6RldzwfeN7KXmfd/srsWjGbOZMcGJl5ShQkGxvcf33pBJXRMdcHImmrlTqa
JI1Jig1gxm9F9NxLyC5oU7vpfFIW/rXQEwB0rgfk7CDEx7Vw4BO1v0k/G/r+CJ+L
kwFrl7z+MHdJ70e6YUqdkmFtBuQme5gKNwpZoiQ9zHjopDW8QVCjx0jb3HzE0/Ny
RwcLTuC/0uy+YEELGPZSZ7+ZIb51MlT0k3nvjmyfKLCU9VodvHykc0aoK+whCElM
rdFozhXju9Mo12RNQrsPn6lqO3jFda1Rr3K1oRQfj4C90VlwM5Rgj9kfVNsStM0C
2H0h13pAtiQeuPN8R0LFkJNYADv7axLvRRVjA+4L9bkLCpZx9h1UarvVw+g/MVf/
0weoepseEprea16SycgAMVU2nhZdvhp7qvmPjR7GeEYHXtBoIzBTj0CzJRwK2jC1
sOf/k4aSAkAtqy1l0euTYFH3hsiqSyuKU19fklB86gl3CTaZfjwaYVBouuIY8mUz
AyksFYNI6WNKMPQTEVkxx6M6vJYQO4ItJPmmai/yOUehpo0ZxL4Eh+EBG7XHkdAO
mNdnjfOPlmwC8x/EuOEzPv0f/PV5M+casJJhtiLRzLDpCDGFj7Q4/lbPXovFBv2M
VpMb7s/LLOPVP92TbviHBihnu7Gcvl6KM9qAy1HrLMvI7nX+IwKPSJjvZIIixl3k
Uq5dib5AgF3iMOV2nXJVyCUYccIHWgCmrvDUNaxFUHuRXDuW+09t+r0JNDvO/pAn
qrUm2DWSRTtBTfnlVshJBqLDqCynUN2fjFjKUB1bJ2yYocfd7KVeSBWy2sFLRzdL
Yr32mG0otk/Gs2hx8N/4/BVoL6EeaHqT4oEpgDNlJ/r5J+FuykV7ksR2dSVPWGUE
7bGDtD/o93M/DVBVv9NIrXLaLw7IRzvH6H/9Y0C/kK9uispjSyLaPl/0B2VSe5Mt
JZNsHGtBL/EesiRN+Q0KuRAKw6Rqyd1SMishI1V/H10qY4WLO7nBsu8g4pAu0YOJ
Ly2/b+ZIF2rbw7P3nZfzLhd4GGDwTBcAfJielsUBxxQ/tp9zPeUWMy6AcIKHeZ+Y
BnaXK/eXa2kHQHCb8MBTNAARs2JLtgDELO2RBjxdlwoiouQL/BU5P7mjVrzCl0e1
7fr0gJxv6N90HmFkJOag5sAu0djGeQQuhAG8EtNtXWD1D+34BdBD3MDlnyRNBsXV
Y8ExqW8PaQ9jP/IBBBDQxQ9WMg/u5EPzD1hho/aN2b5G7LVwPknd9la37a3mTAGL
rKlh8DyfGfIxNsUlKAG5DKz+MrHNqPcLqS4NmQt1L5zhDLqTJ++oMZdfufVncD0O
LDqKSk0zFR/8Pm7ELHDmAJi+clvEjm/3ove1fl+sOwVMCzztIItTRNOOY1PpGH04
tNaRervlfgKYKhWqPYOfMtaWH2zmcJeE0NcPCX93giuSLtKhqrTX3an0VhDXPYrM
I5844X/g2NSCwm85KikH5i6xsWEp9Sji/9gbyyODfHFaANCTVJuj7yWfPf5n7CKc
evK1sDyMBybQ7aOH+kV9S7K4aO4BdZ9wya+yIk4dPEy57Y69xbBl4X4WSIogDO1k
FlVnCErO+gYOEbHBiIPvpOWmR4VlfPRjNf5N1rdFmMr23/Y9wVGl1HCD+SXuAkaD
FxZPgmP9b4BrqS8EUbh4ExrvOD9LkpDoAzcchyk5/U/vtSD+rkpI791jcUip9oZo
igNewLff4tL7fzFBq6e+oYI2iadwGsFOCiFabGgZyM0vdYEVVVt8BXR5huyhZNqm
0sYl+5ysPEi4W4TLjbb+nHSNWGyt2boseKgmrxSPntv+Jthn3r/h42oR3SX+hl1W
EGwHPe2VYdhjlwr56K8qzeQZrDuNt1vF1xIEphImQkN+O45YU8clXEUmu4L+J8pd
jFAQARxRS949kNyKT7MXwM/VznNXSRFPhGIudobg/AOQ3YC7J33ApftlPl8Echl9
XYwNYDfrIejGfRCNgqkni6rUKsECFLbWdBPlxbqqfIQ4e73C8Kl+OiufUiQzCgdg
D1mwyUmt3Dj002xODLUaTCbZoYLV7Z4scSzCoapO1iHOt7oSGf3rS7ysdX9fADmB
pkhCRLgtnwcv0ROFuXkUFX0jcGMI6rEij5Yt64IG2UR54jbKFXM2nBVYjCykWlfR
L8Byq9wc+gcSqKBUIB1nj7HJAZYzOqNnCQK8eYI26NGeav7v8UnfZI8xUKiPZ4S7
4Uxgbni0MC+p6caxyC1IDbIhzPa44GeNZFUamE7gXoLaKhjruYzB4bnKmdBKygys
xlOlDxQKbe+5WnVzXyM+1fdYFWDJZFw2vecEgmtgOIXGJ8YkuKxYoWbeg8xpO+4b
n5oNNDO8UBmrVDP4ITiZzdYG8kjKewx3JEImEnECX/1R4gFMa4lCxZrqgdRMPFE/
3lZK/5lC3Wo3ZKARYHTDcQiby8/L6qCC/EiEUZtf74a8+Qqo3t0gYcnT7rOOxiF6
UtDq1DKYx/bh5eKzfTva99kBJ7exj42psc6UwWF2yr5ZkxG3jWw73Zh5/XJARFEz
vBqsm2B5u/N5oDmK4YcsEM8bmIfJ5is2PhXVJFKOpeSkoNxixFFWjyqgdrmpUnIo
Gy9WHTp3UNW/mbRW4gY1rciBMOY6+HKD4U0fsxCuIMwrC+sfhCyotfXRxFdEKD+I
1MvtWNpxUiK77NFdVOHl2Nvydw3wox5z41feHyBf7AsKAymUxK4AKTO19AHEdfjg
fmlt/51Q0Tz8UDIkDA2Id6T3NOOVCPILQtLDu69Tte3vRqyj02UGlimpHsNzOhWw
3rgi8VgHEPqLg97bb28nZCgBp0PXrV7lIYiBOxisma/PzXq2ZxN+HAcTSnQDQnDY
GBZZm1cFHhEB54a++Po/KmRICd2SIBtIFhL1iF5g50ik/QTkvXoSOndd70zy7doe
aCkP57mwasfvXuOyVql43IJBGrmPp2JNokSgZvvZj3IGHctEK3FA5m8mmi483FgT
GhqtEhXjNqA//D5JqFJVsykKDFG55pCeEV8YT6yLq70Qr3LR821BVrOAAPqgbezU
zWlUFk6tzwOs0cchlzE4lODCKC7en3K9Es5WEXlGSSSNnYNdkgu2tQJ+umHWDcsO
csJD5+8WsuzrbkGfB4ReNAopnuRwYaV5IEJrr4YFl5Syb9c7idomm/Jk/Fl2vElv
+TOWAAL+UuqCbmQFEdiBEupB04JwwR/4LnB7gvgwWxuOSNM0nnNipgzdJ9NrrnnO
iOLNXgWPjRxCB8JSqFLx+8bH0R3YrrHdhv/EncibX8I1LoUrccd9ixiW338m1b+c
Yy6hP4eEBOGtWffqGMtqPIOSDWnhUQtFJr94W3JkxGqfCI4Wnbmm/9fwtx0jlEjG
QBpc5ZkGJt9ceMFPiLQHpZkZ4ZMCfepckCkm1CvAmAZBlgEU6ScCuJEWO7U9wnlI
LVrVSDOgJOjAnnI0mxLnGAPB54w6kdqB79hsae7VANLJLVuqnWeLtEZbWneq2JoL
2UcEhwEO6w8yKQTtHJdk1ZNa2VrNRRTddqPXGamSc32UL8gIpNv9VCqhZIdmZGgK
DzGJbYr0AKRz95Qc7gkW7jwPDCZhavhiELrrE5Yo7jG8D706JXuov6t7WKiZReuX
nAdiXw2ettTiqRScPrW02SGJql1xba3JEDGz58nQFdBFkJWcxuOBgYKiHP5IxhJL
MAZ2PncKs7T9iy+95LUwJGQOOj6eIXEue8tbsez1RJtrdK/bzxixYWFglxetQkNN
9bW8+lRshKZwSH7tmZB+A/T3gu0Cye6AE1GqRq+wzJYQCgJEt9hgO1Mu/zCcyWDA
ElnRAHBbEFvMcYA0wfDmjTPKlbl+DfCSnjMfuaQUF0CaekhjMnWXDkvAMXkBGtXW
VrurBtp0DzIFABO9l/qDq8Lf3rnjiClwpI5Wj4Si9E6s6Q2vKzbpeE+tZWHwaW5f
0srEKDfYabwuvgibcXmjLqYo8c9Soxtsgu1/lUUapKlMc36BhW48eIpXHySmIzsI
492U6qxCyWTVCEl1N6asW3hEAPXU7kSbtDQNye+DRvmHyTJXI7HrjJx+TczIi95R
V9gCjT7yigXVNPOyfMYpbsEgIhfwAw17VWapEzdDluSWY2wXV24qEuK7yl8HHuOz
hwUV3pkzvX/Zf0IlRz5Xy5LcU7rTLAmgR4If9SqSMSbfv6JcLDmFd/MhUfSx4dRO
YjzNLiGWxaHY8txysxjZ8Xv3GIQSCa2/9I0M0eEmUCyqrVk8I1nnMRZk41Djt5ij
DA12nFYpcyMSGfzCLXjDFS/FjmtUEkWdsYZtsygjl3nE1rgTXnN58mCrxTkyOrK6
QdEa/fdx3Xm4jPMFFumqII1jcwiqaan4hnNab6DxyKrNQfxoRlTXepB/Ki5V6BEe
QDlD0ZY7iniCmBHB7gMGT90rmLKFS7oKCMBEhc+jqQLnc4xvjA5bASluUtrfw8YM
2WdZQP3pE7JVK0+azzRYTtwfehiEHD+xQ/H9dI8VZJ9e2+0IzBePFiSxgCcaBK70
nwBvgpZi9qDeQHy+m4Qkuwjn/MdW+ARi4+3DbVsooS1XN0Rtl79JFZw4z/aDji8z
Z+jwLgYCA5Z+ghldAqvXLSxE0srrZoDPQYsKXCsrLkcp+o7hClP7wONgYKcde/ty
9ANo+iTXOhnOBjGWySbnRtHl9MBBQtkouvbFOatgkkeNa2XrMFa5ibRysh/THm/N
iysXipnB3VMrOE8MDVGYAtGPAFYsCBDhaS2iu2OqaFsDtzJP5PQ5CwhdDlUCybzW
KoOOS0nu82dvvDiqHgs6mKqsvfqjNlSvWhblTY7b3FANbs5j0owPsXax7RJ+4Qxy
wknqXMrlZaAFTSzpJn+5GIb/MZQS3ACVDVVh3VjVH78AUg3Z4ZoMuF8EFRyx0Pmy
YIyA9JZp6efxqYnsvwJADukX4pL0XIs6ZwNFG5/RjdUXvlGvMELjNs1VGApP3JaO
onCwP45X7QsIc6vVaUFMlvzRZKK+n//q5E8ON0zmzEeL88tu+5ulGuFZ7VeKDYRU
otZzRBBLQhg/ieuM/IJNGPZ0VOiLc6Nzt3pGv/gLM44vhW9fTse916iCnuJPuyCP
CSLBh7C9hii1RYpCKpOA7x2tSuzAov8cNPQC6XDbU2XL49xX8B6v4oV5+GfOjax4
VD6/ZwApsxc0Vae9MRN1K2oKd8vo23077eHaDEdxNuK7v7vmVr3vx+fu/+JqKikK
51aoLibjOVj5xND3Rh9iY6r/p5xEJfTLHR8ve9yHdnvD4KuDD7Ju0ciwva7dZqER
SVKj9J1pge15ilTvGa1c6IQ+KwUF43M6FGD/gq+AZo8Br/MmNzvqk57MxLzdtB9A
wFF0IK7vCGLlluWgbjjmoicZd2yUMG7fC9T4oKorxnQ7+FX7y0BFhlt+n9CsiVyU
hFNALg9f8QZbCrXnRKqKKUmZ6eiPLiu8wLw5iORKM05NFkxoiIZprRtrJ9CQ3HKl
hjI/7S5SlGjLQBv7U+8rzth8PJJAYt+KspGp08p34tyADfxfaGqgi29jZEbSqzeL
+VvMYeOnXNyUlqlPhiFERY4Xj81+n+i5mbo0HYSCHkia5bhapSnSqH0vzSOgMJWe
GBFQd+AcUhUGIpKnVifkq1IhiW1ojUV/nqqUo7egE8nf30IFgJbfSwu1jG/EaBFC
2wVkRF31yUvaPt82JAHOByOTK247olm53UU/icPuKjpQB24zdmsLrVagB8WMYfR+
OtvgCzRwDdKT0o5fd0e/ttJ6xIU6espPtWvinKcWUgTYkfiK8PMz9LuP2WlSfBu3
xYZoyGpjWNR5SygQmD4uXQpaN+M7UtrmFPQ7N1KtJIh/HiEDkcapCaPuQI9IJwBU
NjtuAmLN6LROSTjqRrcHOxQ/HHI1ozzbcbvx5RenxPRhR+qDWBge8v1Ur1UHa9Ph
AzGZZepa2SHNPbtPDjedWpPPdPVfgUzyLus8wCO0nP3E9jgZS9p9LfC8mjmIQhmD
Y+DsOoTJk9vuN0ykhPNVZ6Kf/mWBL1VsTZfKO9LbCfTt9N+IOnWjtcTE8wVWNttb
9txDJbzNQiwk+J/6+AGfUTalyOxdQXNYNbTjfuMURDJRCNHma46YlIOR4hA4e9eP
s69Cb+r3vndo2i8lUQJ/Vm/B4o/ra4SzXw7mr7mmZMYH95Sdu3zSnA/ukSyjTBEw
VMiLH69PqEA29fxRTPfmdEeZEW7a5Fl01lSean3fLlisvgILwuEHUO2svaDyP+qh
tjdQdOWBZ4YXinZTym3ZJJEYSGAAjW+GdU3a1ysaWZY7/a28mRnIiEGmbo1f4RTL
Jl13LWViE7sXjuSflhxLJbwv4Fm4f5MCn5V7OUTz56dQPXoVX05IGjrWUWKZyWI4
eMUytR2Owp0DbaYawoJOxIO3jcViXPs+P6fYPiz36AqF7GpteJncwVjmFUYWN+2F
urOxKtwes3na+RMD2mij/J0SqsTu7xKf5v6R/d0myh3uoqDsFRTc4l/klgHJOvtk
cdLfXFQ7jdjE9rrdwbYd087pGY/gQ1InOxGvaRx+UJM2iHmp4agMOqP35b2yxPdn
5AVEZvbQpZ72Sut04+R1SqHq3VejlKyOIkH3BlebMuzlWhNYpioAVjA2mzI2lZbq
xe+wamvyMj54xBG0Cw42quVL0hVEldBDk/7tRytTbsOXXkH0yuQImbsf5riy8lqR
vkQYP4Qs47Ned3E3Mb9eqhh+j8txHScnsfr4l6n+pGwj1j6XAtKZDwWga+XQK7G9
63TjpZWEoPl1z4ao2BnlLZ9s/Y2faTPrvCrvuCAl4M8+aEBw87N3sOAEBXMpiLxJ
7vxNZ9lGgSsZW0f096POuGn6/jtSx2SL8IvrU/lOwMAPFCUj1ykh8gi7Kfrxcl6w
LQWapIJt4ugwknZGUIk3iNXt5BtPOCYiyf2HxiWP30xkiPwXGnOYwgLhfvhjYFBg
whX082yoRDepyuSgZeHIZcpTipjmbmAOgfWVnDfS9YA4Bm1tqv7nrKabGwgho4W1
/htzgDJssau+BKV4UNrF+X6ZEwlsrhL+I8vwtxduiwrlZoEv47GR8j2abxDftQsm
Ti5WdFmhaZxXTrQrcDXWJKR0O5mgD+htIEQzxpqAgq9Nj85FYJ/SXRanRqkpZB4b
J52rBX7O+VbVEN6LxJcixq9TZAibwQyI//qOeGrXuGBI/ZS0koHM6J8oX78YllXb
fUnoqfSnjrKFhOHg9TzyiCymUGKELF+LvcLASk37Vv0IwS8ShshNGEls4gVHrQc8
6FUChF+isESwyQ+BD4wdso0kuv8S/Ueyi7QCLUiYgmKcfqv99UYiDUoMpWMiTtHH
NWSTtHVIqxt6yi5KsQP54CzMcfP0vy692Yped29bkeH5HdHlzW/Oe0fKhWp1nfK9
PeSX9XORoDu83LbMjeYGQfr1te1n08W1xNKmJbyP3H3xm+86Tk532WQxJDFpuX0X
9wvscRCCZJqyxqzL8cNdrzjZX1RNdvhqkL/4GcE6Lj9qkOs10mqi3goqSeDWwaID
kADv2IFBQQhE5ttEKwxbovIlKsIsFsQOkld0+6TkcD66ctAYj78Zb2KaLT3ZHDrJ
U7M3JIGtUK6C6KLOsvmzYHA5Q2FyCaED9wEZRDTB7rov2+jM0229FuoPKiuw/LVI
+P2f7ckawLZkbAHnLUZylI/dZSwQy3J3MR2TQK7qLqa52RIi6shhRr2KxzLTmJyX
gB/zc5fNgcxtB9+1dLQT9y8Tux1xIvF0eyjs2KOPCwvucqYsGZjXZmQhbWvJIp4U
Z1ioX8CvjJ+sDWm3OhAZPUmfCm9IOEMutKbpS2/yqU1FNaZYfiRsc5kMguW3V4Bm
n17IlaRwiLO8kP9AuvUl3qI7u94vBpEUHehHzm4nwd9csuryr6IzI/jQ/LdPHSAe
EocAXbnxhEIJ6hF6GsKic/8peF00fB9txP9l0a6+QmR2IuDES0DQUYU3sQvnff/D
JqHG3w8p/UQD1X7cAg9H6s7D0tbPyZOAplEcKvUDJA6txPhjGvXoDpTESao6Grgc
Pki7NMDIK19fhj2QQHF/yhgcKCpQ0GPsMnZ8ivJBgxU8FkZZWVnTHRpvo8fobwUC
ybYuQolWnQNPEV+MAy2zHQFZOOwP9/+Hi0XR1iIYlyqoakGhyWL7PwGFL9N5renM
H283X7fKSfS1iFpjBxhGXHrjlKeacCLKRJJBSYn3UbL8hVwN1+iBQ6m60s5CAjXn
11MxDh8omtwWT6QNsMvnUOrFXaeszcO+JPLp8JqfhSK/hUe2lqYCwe5p/yPWwIrk
eKWzV3zQYNDX6IqJOsCMmYQpPSJefgcAhTfyhUikDynZVwi2DMnTjbKGybMXOgIo
WDBtUP7AxA6/Ud3zMLJbMeB8m3vAJRxeqlwdyzJ6HXI5O18q4ZeRPJvCHIqI+inW
B1ywL4iy8+q8ZjOSw7WbvLHQT13CsLhLDg9NxRbH5+Buv43nm0ifHhzj2DyTSzDB
yNXeCbw6fbLHTm/45a3ExMkmXT6wJDioONeD99fg0yMJIJUEXYfMUCAG9loaZMOb
ZnjWStkTmNpk35cRN0jB3ZyZNd3EP3ExnIbrS4zMTq4SlKkRaBa7M8hh7iRFKx4o
PamRZaGdnLOQLCctW/tdMZNaIQVpHiXh8OhDTfMC7c5C02Io8XN0KFC526WarDOc
/lHEjG1J7kpSxfcRqbZcwTIYyFEp5CqGewQzcq++plQO3FF2gAj8nr6UUbtZ4QlA
hUBr9jxlcYTWU8sfL1HOVLk0O2dLgYK8dEDA3bbD6slbGV/1ylHMMXTByAs7PO27
jgL/wprLTUChSPYQNvTIPTDryF4eH5dCskzBTiJR+EG2LooS463oN18A6lU4NhCb
Vff+nI9L/ggciK2zYcIB4p00IU+f/Ph6R06rVb3OEk5sXJuwIYYGPbyFd4vYxNZ9
Q1AeaMCfTQNTFVrrGim6ioD5nZwKklNpfLe51faTcv1fRos72O5ALlFGQgjX2uBR
JEwPLKF80udwiaY6X2yYfR3odkIAqI3LmZITjdtwQ5IuDiXyO0n0PvTTpMQx34Qn
WgB0IHt85z7x8rX5SK8N/EBT712Z1b9K5R2YQRB7XdP60G/Io2DFh8cSuJ15StJh
c2+ngg2fzYeaPWhXDi7Di48NfsNnX3LTbbFa1c5uUhYz++ADkDByvYRT7vNeR1H9
3qITnBXTlRB+M4VOxCniLyEQ7m6KYe4fVrjWmzhp1wOZPc07zJ12rPxAJotdQ/eK
zRbgZKwsQ+2ah3OxtANfJnMWfwgwVG98mYkRq+eEN8P/fB06q4Iu/enEoEnihFP9
CIY/aqjreDi817rAbZpIsftxelBS3UkZtwBrc4lWOPgDLclBXSie5UrVXFZDekY3
V+KziJClUnM2JWZaQ4Y5n2+cd7c/pmHSXexQnfUfgDY8p/IkKm2gShC8lAR4EMh3
8BGpHncMNAz56fEQQ+b3BfeaqlO67nr6pjwo0p9cRRkz0ICswlO++SYwFLVcUl+6
XJK2u3CEZ4hPZ38jvQIYzMz1yBziDdNjEkKhdF/93WmX0JYMfCX7tjx/Rv370ITE
H3zcbGeNsrmqpMvQFy9ixfrAxhvdOluVc1sPI7x9ON257g0zPi2kpcLhmFNgYqDr
yayK+eHYIn35+Dro+0OzubwCIhvU7jh+nI1Q3nzAwxocDQ179xRn2cEyFW8VXmn6
z3nOKNNd/yySvUz/3dTQ60Cf9khZ+1/URefK+rrB4ymP42nwtgwZGHzOyintYAsJ
rfA5bmR5HQf4LY+C+WOgKi/69/6ehP4b1PfiP+L/FwbQ27QrraBmUh4QcQ6DcmZC
SR7E2r3daO8wFoR0078NeLiKca3mofzg5ra4rckBmRfJgR9YjlXG77qqPL7mfmbT
wR0qmuhwpWT+dE3qcUL8fEGjF2SAFYrlvEWWv6tGS0mAbmlGokHsuVZQSGOEqQH0
JnRUMLNtcI1UF0zNaEklxT+DcopKAMlf+nZPsw2u/i6xwGD7hTReZ4czuflbXvyK
f51u7hMcSEmDnuxiYscfWIxXJkig7exAJso363agZCEycXzhEvXJ20yZWpSNvvsQ
9MF2KJoXw0DzjxVERaAiIfj/zcRzl+iBvwDfgOM54C8J6Tp8v/S6ZnkpEgGyeKlr
N+XPbohGGjQx2M6AJHU/PE7NXzRolvL7QHDRInPTSY0Gx9zMuWtFkDtqJg2N3R0B
sXlrRE4W45JOEHLwhg9Z2C4SWdotckmNwWX9Hywd4gRTuwR/sSrGl43GlTj2iP1q
dHRI0zGUEgQ/DrK1s+xndoEiJTA9Fc16UfPUvK50GUnU69ebqCzY0+4MLB5ODYeN
dfEJ3VKYnyogo2M3Lysp84LTGK0h4Y0Y6AVH64FdukqfuitV+DBEM+h+4sloSBly
X58R3ANvwbicqcX8uGU5/lQX1+ojf45zhiRsU8w3YJh0uyHED4qfQ1bSxnFyeaUh
ZWeVj8QJKSYDUU723k36ubscwkDhsQvW4hsEV5rWxB1Ko1MtAPahI22jmsXHcX+4
dTs7ZsLoB/xTjdO4NMn0c46WHqSgM01b1lWs1xlrgeNx4q0dIW6HmCx/OsvBLVB5
MqgfiEtTD+uExC+BKLFTBCj38XVPJKls7V+U1HNE4SRTyKuGo/6ILYzZ1v2ucfkL
2A+91DeCwJctrtVM/rUEoDt/tQb9jqSHA6FXyMUEzXTGljYxbHLdY2PYHVUebNwx
x+LMxNgNy6pbeZ2cK2qWfvvS/IAJ2Y3PI9tQTN9QzyZ/64/hVPvaOKzis9UBsu9Y
QHa44ebTD7eq1sbK8u8PsP8GW50aVkJe1cy/qCisVmFQYQathOUzbMJ8WvovA2aX
HCe3METxqsSOgSTR1yMdfIVXj67IP4ZB7su1yrJJ4m+RY7kwWm+A/m8iKRkbZf/O
LIYV8zXHj2YJDqqodn7ZuAmc4i/FfzjydGukKKF9gxNfiLdew6jyx5lOgUGrpnj8
h0HScwhtxqamUPPjOzJ+QBPz3WsrIo6kJh4z1YGl0qilJ9/PVb5gj710K4qfmkpJ
ADYpA+M935SGoqicVbTJm0NAfMIvupbmEVWkAUa+BORkLC2XogSbfmS45lU4sivZ
M9bg43CxaF/bQUwqpMT5IZrk0zSoutEV7stilRZXsEK1fyITkLTkGLH3ih4WjA6G
Op4bkLNVgQEw2lEVRSeypKPGy7L3/Hp+TZ87A2jLTUy9LACQnFZQu76mLMLCdEwZ
LFAA5ILSQiNcedyxIi0clATRvAAAquXQRKoImbvdoq9p1ICJAm05cNJWHLllWjlI
Xp3o7R58ZhxRdSzfQXcB757OCgqCHC1+HMCbd0d/W9wMPOLSBLbf/QANu+JW1u2y
GuxXEMlKhK/RML7lLQmVcfRNHafuZH0NRC4t2TgTdxE9M/OfZCX/uyehgRaDxpmq
GPE1tGpq26mr9SrCGdrikJ7cGGXG2+rUlao77R27GTaZEhBOHHt00Cx8jN1vBgdg
iVtRnXGYaamRAws/izFmbQ+OCD5ORZlcN/coQwHlrYyKDSWE+togDvzfHb6Gqt/W
kGHnGiOj5XlbIzuzaHpbyWzKUii0IteQeRurwHkJRm0zMrjLtou7EXVKDDmfF4+O
UKBZRxCoicPts4Nz5FfJ/xaqu0aKMiElOEi9TItWRVALvYzJX4F1AUkOuW8wS3ZF
ZBWg6uvFmhMt8LCniVo/nZvqg27osHbkuwIHwHfoLMXyDH6TAAHsS76VpMSMuuw3
jhrpPtqg0U0Mmf2s32oD9OO37WfEEiPE1EYnKlL2fhDIyJP17yey3zRtJG3PnHD4
MbJp8SPrriZxlG0PFhZ3vjqScT0nDAylm+QdcBqhxmz+7Rt8k71jn56Iw4asS3H2
+w8r80Dc3mBovt2H4nmMY/EaTyl60rYp14Fw8z9gi5XlvrMQLUmelyxroPII2xhJ
546dmDr0XFfI4CFw+kxXmTXWEPVFS9mLQQTCz0lcW99KrDyrbVwoKKAyssUadRxc
3EW5taG3Sm6r0tjVsiYWEbfNXgFkEZhT2csLaNyRUrga46ATCuBomG4A6nUafeGc
2lH92fuxjBCd/F219uQJ7HbstP/WK14cDBkerC29itvEQxwTLEoY2xyvl8Ooyrlq
VLyJ29r/nrj8UbHAiZa7g0GNM2aYOjN9X2BgTDry9b0Sh9XsLFZFhB003Z9SIyIR
P53cC2uhun9XDgtgcPXu+X/Pc7+k0hiT9FWQCJK7i7DF2ozS9WyprBr64qguNUcm
YYTLg6L1ejsS8SlUaiq+qc14R+IgcLNIdNBxwTCShKb0c1oU8mkD4RHWBSUkwrug
/qv3jNGdx8gQB3hhOvtvSg/oPCm17NQxiKNqA+/3cNL5anRI90SYNyv0uwup5W+6
y3wJysvYsEEQcheJEGdJ7d5GRwIHyDaArORctI5ZwZPE7UmkZhW3fe1z7mPfoRFO
sC3irh/18fd8TZSP6TOFPWY70PlZSxKTxxCbZ/gH9xFZ29M+uWUJe4Ry5onZEzbV
zaFqHKw1VlQ7r8KAvXcleVBUk7wtvldp/z0bPYIompLap2wdzab6/yhnq6GMhcv3
DGGBqVs8KQXYCknNScXiUDemHb3+FlTE2/huHHN2ZiPw2xSkI88pCiaLBA/Styfr
GJnXqo+Sab9rMdckvsAW02xmmTGBVhMnqiBeJpMehE+LPdlkZ4z2hOitnpieD2ko
nwqqZ59dXeXDAB+4gEVZbkcUoaMxAdVjVNPsXsUWww13MHh9Q913lA5z0KcmtF9+
sgNctJwCF5ukPFk+0AnMkt1IkXt1KDaE++nwEAUVJsRHFKBO6chS8M8IFv4I8WZq
AmG69VdIdqbwLTixJWoXYBVEp8FUhOpF2DQR+ZCwMtJ8kVV/DalR0fCdphu1YwQn
ILszgXhEiV8jQp0WDjWNIbn8khEomh3q7UCzh6r+yxOzxS4DtfRHGkyWrxW4Vi+z
ZqPNqSAUb4QLo12sI46xQtKqBXVZHSPIJ8y4hXlrHmWxvN8m+eaUc1FDlR2+eq2+
PPSwoZNjWPScbsjtu9ZIOYYcIatjBNiKj+uyxN9bYhN7qkm2VoGos0jGeAPVdf2U
nd1O4kTsDsQ241hx2beR1cUjoICNiEnx3S2Kbk8y0byzb9i4N/bV5RkBgmhd7JGP
HjqdGVmEGtazLX+HxpChyhr9yCzWrn+KbaeMwvbL2JFeVGqJM8+BWGfz4Zsijflc
zWgMW89Vo+wN8XR9hXNGGtY0v2Ao/rVpuV4DQ6ogWtaABH/aHZCSW4zWiwug2yoc
p/Gmrj/uCw9gfGRcIwfkg9w1jaMWs/qeV59b0+tP1w/O8Bri8R8yCbUW5SbeQ43K
WZpPDY36KvW9l3S1hxWpCXjqgh+S8Q2euaoiowHDh0dtbE80epKRyFjJp6RjlGNQ
NBdZfwisNtsVFxgaA816O0rmBaRFQMSJC31S4UYcahoBwe53XF41dMd/6dZnHKFh
va5Ji4I2CL1WBFzETvPbtAktlkJYrqTQ8UXovWZ+qUg5vBif+/Q2WRWjjjWz1qAL
BK0DSgTCUeul29DaQ+b6LSAh7A/CKabfBaenlxsqtHAN0OfiZNsGEKffKSb8H7gS
XXS92iBbme5e8xEDP1cMJhmKYWTWLTMjVM9U/lkVFNdR/I+FFGy8RJnmvScUyfq1
Ssz2pvBkO5XXt5j68klPrpy5uX4lJ/DvmiHvxF6Cvt6Ll+Am4fjZviziN6UhPslA
R6192w/hnUH8rmwtycCPS0S/d3N5unVF36UhgiUd1cU+6EkuhkUlCYA9K4ry9cDw
tiJFwEx3bZjRXUNOMQVCW4dYan9D5Au8Vu7UjuLzjiiaWxuwFDBvCnTvCZCKvpsw
LGAIwBaOfbShP3DUZZOjjCKx/+2u8J5U0hpL9NVQyWQFfjSJPFA4qDnGjJxBf4Dd
iYJzCmf+nOt1V1aIZCYzjh4ICrrgcIacWQglqTUIFTt1oMyLXqoCbOB+OHGFKN40
uMqZKy1cb3Ezfg6J2CfMHPt0NZH+H3RURhcyazKG8O4oQ/gJ7nQ3uNciTPWdZDC0
pXNsiieD3TRdP7IA7cTqthqtIFh34tpNLsRS7hOnY1Bb34YdNelSqiNytaq47K8W
Vf5h8qXEGnrbFcgA1S70r9Kf9c4GdlD0DHd+1LoagsE3p9yBefn19FKcqOoGAqyh
2u6Vq7cgR7MmVKzDDx+JLHuWYFcI207P91sLxWo5tWhvu72tOqTQhXgTLVG19noU
f2NTDUVInCB7LABErYR5VKDTlLUPsNpvR4Vw25QR7mCCcfwhCZXkegbeXumPzLrt
0IuzWUMzJxs/YdantdroFg8Rv0+sDLjcxzl9wJmjbo8P+LYo66EiaOuJ3TKh8FuW
rkZ2FcB2nT9Qp/lf8w84UO5kSvHmvr+rsdm74lcRYS3zdmiyml7JReNv6rv14Vd5
5n939I7JYh2aIG5QcCYRHjYCcHcH93/kGIohaoXq6D8TacVUMyWvdJl16WAY6xxy
/0JJ6NZMQZcchGXeSx0PonBY+ZdWAqq/EKJ62bej54qCMg0dh2gLA69M24Rnm4xi
N5kaA22I0oXhU0zcCdFKIH37RDpDyOmzQ+MejTto/Fs1uk5dOLsZd1/qegKsX1yp
1uL3ewybRhORmT9VjxygJW4cflqqq0tQpG/D0Fgb3UnwD0CHlCXz0NzZw0fiKy6K
XRwvBRjITQUoi/O7wVrrRt6KMvoUf3iUSHY4FWnqCmPQ+YEANE9ExrUI/+miE8uv
3CJBBJliFwG23LGkynnhv89+hwIhwV8okIN8BEZTJuiGUi2ayya9go0KJ6waicev
+ZtZWfwdmFouFj4U0A0vpx61koK9J4keLDsyrVNksJNqa0+CvhuRN65udra+LAjK
eUHWoeSM0t5G7hFkxWOJs3ATuL4uyo0o/ma2jevnsurDvZZAOOg9bWaWA4NzIe/O
wYfTYMRkJYwaPsXvI0qs7iVIgyYG3kJPWt4qUQkueEsYXD4H2jr6eKFA5ko95yNx
Pe3IeAJ7LSLpksSMJTTm2Ipe8SsTmKcjx83CgRSF8Aj0LATYR4NF5TFMua4Vma+W
v08gdQZ+DhplG1YTV5GkGd8rqi9zHabSbqC+T2q053mZiZg7kRGaJwedssVpn8Gx
PFEN8lBMW/ZgYEnO8u3ER4TBiLzv4nkCaog94OFKshnxSL9swwgvMfvRT/LE+UAf
WoRI3auWDKOG4A2vKEbfPkPw97b+sA7lPdK2H2rVb1UBSdUf11NNZ3R+wLat8xwj
mMZboVdNuDpMnOL3ClglUV2GpX5wY9nIn+1Zw1fpSVTtH8b1EETyIfuFcmx5Q/Og
kbkF/Lc+NkGbgCcAZyfQ9lvCtNRr5vtNMtJso4gMYYh+mMUPkls3MglrAbxKs06R
NdBPAHhLW3sOq8shK9Utnqg50Jarj6x3y9q10zXRAybV+lSWEHDgh/0HMI+XR4P4
1NoBrA0YSj3Vkh8U/9AU8SflPKu6tfozhIK73u/D3b2MnRDXzJUUJAWNAwIC0C/k
eALt1dAlA7QqpwabOLhotYPdpYUAh0q3X21bVLHJYu5UiE9rMbBpX+XPHZzAzFin
zFAQnkX6QNtZdt5fWS0lh6ObjbG29IFaf8uyV4aE+xBkKEJZnY3/FvM3Ims87sX9
/qK57E1dIRFQ9TDCIdBbOg8MMd56TSItpeG+cep+Pyf+sgvYoOrybVknQUAkI3pf
/mNMhLtm+KfsWj3Ui6YHh4aMOW5tFP4QX9vLQ+2FOELt1fr3IOo52kEN3ylUd/+2
ffOCExflumrYnas179Uw7UL3nbsT/ASt3L3rtJXGVpoTAC0cOxaB0IrpoN3Zyb9C
HUZsKqZdRxJLflq8jjjkxKD3+W+0BKgC1Pd/quvnZOBuyvAMOFP0oRUommbb4EmT
Lst8VoKL6gyhrPnlgy2xtj/FWJrbx2+TqKpLk6bK566NA7JLHQylv9jSGpl2onxd
MceUxiYk41m8eF4eqxoxHmvTSWQqZs1R8iJYgMXn9jJaf6cFHKuELItWrm7PwoX1
Yz4oVbwGV2tc+69pPe80F6Ca8czpijNYHvSRRK7i7o+AS7F9xBKiQWGpIYq9BeT8
WS8L07t6ehi53Wb5QTE5lfZhMtGyJOKlrV25haFCFsyPE6wkVOL+A8qi+RzdkYf8
MAdjAlCHRZhXO87/cRzUiBwUrGONJWw++264jLAWkQwmPbAJkaLH2bmJynMnul8J
uhe4V+KYdeWEK26jl1yQghAA6DQgAv5W9VjhqZUjEYuV/Rb7Z3BUpqGa+BQP1NDR
Zqn2j7h9593ityOFEb9yHOm6PdxD/q32oBBVDXYFugZfyGpjkasWu7Gx5/FRle6j
reF1s99w42CfhZ2NBxMXy82OhILp7jvjs69Jo4HHDob12yW/1KlbZkWjO4CDl4v+
ay5ulleqoCwpzwYcvw4qG/w1oWi0QE5VeQbQY2meU3nU4tH4Bw8+RPV9qtiL6wvZ
a+qflMle7+3S36UsohQRlNdo8oaD19AqZ8KiBc9UUcaINOb2FPtORPtCg4zJ8q1F
Vq1LnINSxYlkd/EEp/qY9sMWymCKjh1EhISMOJHRovknolFbBY9jL+Gbbpca/e2c
bxC9+x3mTZxbR3N9nnrN9mHtYVLkBIcXXG3O8Zsy03c7hbEVlqlbHxpMB05oakAb
4OLwtvNrzmb4AonHhxwtdZy8vpzLXkHpL2wMeVvdJdv08pbnVe8F6kG5sZJzx0qW
hNYB9IYfAXBxHL4gcckeH1kGcU33+UKzkMJnwb9rybG9ps505ijtslSPCPLvtUgK
JF9PZUKdFqRzNDCSFbzbzY1ykJygy0WfWOE7xuYaegYAcRQozEpqNkvvxyuzVFSG
tDKQOq4WyY1kWHsVa6umMCFVH6q5vJCxDTLLVRFytlF5IOEsEFlnaeXSAbM5Kz1s
aj51gZcF5rTs+FQeivj0J10NsdaCRK4NLqeQnSkWB44bRwvSV6oFltZklZmhrznX
jekjjguZD/9Lmrupsk3cKNNAOx2huKG+fuyiM9lWiVqGUKm1KNdXoGf9//wbzwQ8
OZRx2Qfo7UV3oKDM0ixaxC3cSCEmEVnPRfd7RVPRlXS/UkaKV7ODO8cpmzc9077a
eVmcs2fIxBhFlzGGb04baud466t9ly8u0GIgzPfDR77bHkRwMFXFibmf+UlilTZX
BtE1qL6XcsUZPtQenv0yjJZok8qDQuc0Kmgp9lj+/XeqcbI9PeJul493Qinz8SYT
Y4BH72IQxp5XamUiIMUkbfm5B7iv2+jCvArDaLT4x5OS+wZJ6EYa8DP02Kb/tjmA
cxD2xngU7nelisjjPnacGoQJb7jo9eSdExxFWJF2pRNiB6gU0p8VHQekafrB2KkF
WbISVHUONVHteoQ2R1PC9auHpVas+BZ8SGa3WzsHpuzX61UHH7CChRIN1xNk2571
EmMIaMvF0/eIwg3qLfOsGPPJe6fP8V6UiiUVA2EYhnD+MkviAcBc9VPpLSNm0g8Z
Pi43YJo41XiIk1tf6giT+pnN/rdjuXaUfMOo/K/hNXZpcEBIUrjIZ2VTwbvBMADI
ObGEtbBV17H/kPa2YWe4deExQi7pheP571jsVT/yxMTnWHrIwmpII58/JSSvWpGS
aZvPW5Fmf24ECxhi20Ob9oVArUAeaWDBcb3OL+qFs1mKaDO81/AnL/6tjdlFnt+f
CcNk8BPeVbuysddOyxp5VQEhm+DHbsuvUiKns3vMs8zXEP59ex+MqIl39HNT0Ul0
njRXV+1/mAkbqSnYwMHYF2RbnI6RF8t7QjFQvT0UNUwE7WjUo5TzgPTD9nyJrmAJ
r1C4QwxOaoR272wuYE60LpYEbFzNLg27Q36gM69yJiiBWjFR3pBXs4YldhKah2vy
1al/zNYJg2SAanJkQnl51nv/5A28zscX2EmTHhHrMinurI3EDeVD6X2l4ZgtkI/2
GUDblxWXErkApANfHjuwrRR+rH84aKYzMQs6OAtb4zqjBgHHOQg6Tjpewj3/pST4
3b/X1vyAFRqCSlRjzzTA7Tfh/ENnZq65CFrlLig4MhinLRItpMCG/bsdxuuLSUR8
sDMU87FFGdZaYB/54jtsggaaPw3my3tsq4jeBvgAGMK59bRBEjASV88LZ8JO+h8e
vWWfS2AKsKFukYtaFYX0B0Zwa//gHt5lFe5gDXrLBVCpIXQYtWGcIVxfbmAuN8s2
gVqwgb3I6o/reNEq4qy+QzpZ6VqppCoGZwUzeiKt3SJRIeKzYugXuOcxtE3QmnZ+
FnpC+4w9UAEB/56y7lLKzUrMJKTgkzSn2KymZIpL6hTG+fk9D4KDgHC1mtKqlftH
YMywv0RpKMfEgqo7uktvFNS1Hyhy/fZq7PW0ZLL5l7g1JEV4UJ3Z0hxpEzyybXfI
kvIHsU9u2jDqndX49A/RZPW/1g4V9Wyc8ImAmK2NWaitG4B4LjO81b5oYwq7Rs1w
YzcIfpqTSxzFcZrv5Fm6Ib0LKaOfzIwWKGBUVRJ0z/NLR/LrRVfzLrEItkYL6VQB
pEoRiICnZI7WubeEHLllNyXH+4yPeINagyYnZANvqHAfRkVOj68J8+Qpe5oqcKJn
Tf2L7DU1m53reTKwkvTUyqA3PTtkCSg5w06y0NQJHaLRGsxUDn3Tcs5TeNNt5BLx
lSoFbkYMOLhkSBt8eNN2E/3VTGKXyvHTA4TrD2HhyVoT+MUS5du0YFW2Bx5RCG4d
g3mmd6jor3oR75iPioFmW1qwkCuNgXEkbigZ6GC3Jnj4iCBbJP4FkjityiSs0FL+
/LegEZKezp34WIS8MzhzRcHJzvbME/bIla4vuGGY0L5L/ISC1CinyLBGgvf7PTgW
3RJGEfFrXMkDimJR818YgRi+uk1e5IbKFCtU3ht7kvSf1OHV5tXKx1xVIlssgPoK
4Ryb1ecJrg+zy2pLWe5a6xVkzQ3xiiXrH/hgNUzrl3BA6vixLV4bbpb58bT3UngY
F0ZV/jsefbgSQ3zbh0/pJXCuBxM4t7cFVukShz14rPOHHF3IIdvWHOg9UF55drvx
E1ZMiSnCNBB26fF8lKnPL7t5n02mMg29wkvdf8xQD7ztpjiYKW+4CZW3xRskTp+e
O6i3yxIvQLZWhampwciKaLaGkU/lTgWC6zVFr4cdaEtWkJ8tEYp56p7yHtDoTHui
o4bCk2GbTJhOY0R2ktb7AbbZCCCvz3a9LxWPtoVuZ+cj3H5h2pH8ysnJhPraZ2wr
FO2MZ1PF8b6y93EFuEcTD1Cg2WG41y5rDL3yLGjdQbPuS5yQ/8DITn8j8Od26Q+M
uJcbZQss8pb7IVh/wIVIxi4c8+BebcY2EWyJipLzQgjtAqTxdvuYaSv0SIPLNsNk
FW/wIU1cJE/cYN1JlnAxW3OsgIIL7IvH7DWEL56dCElT1xLpehofVQoxpiHCe2Nn
3gO8YJnRWwoJbnWQLxgM2DFwARzLVqop39CXJzgHVfduXcmOzpAgtmThJa5Em7Mn
dqn1zhZasPNITvSQVCM16PtJKgVJvCbblL5slxZ6sQ5hq+cMhGQsRgOV12QuU2qU
8VVNooJbeqiAJb6ugipvdaJmZuA2e655YVdOrv//lWZSmN3jH7TwcP2y7OIISFpH
CxgFWZ5uTWyWQ6+haBH077JKutQzQAiockYpVPQiL52sPUC+TbwbTZv0ZcbuT4M5
lbt7BJd55mC4cPc91yg5RG6A6043EXwmoXWlf4dgBNOdhHGvb/atrGM36m8+r/XB
Jo6inV8bgpruWxcuKawATmPWmU9UinLJ8EGfDdJOflk0Sm4LWUQk4o7xoJbWAtUp
xPaNFxJJmwyhvSj2BdM9YmdzM8aL1nEUOWajjy7wOlbpDqhulubMW5i6aeYqcyOz
DliLz8EXBs6hpcFFPhw7j4bO7Kect5tjOg5pIReNCMpFOnD+njV7GrmbSCJih3/B
4ucOw/TOl1NTpL1TZs0mPmWeXGc7EQ/HIajgmTYvlsWnoYkd1jnHaGXh4D6qiT+G
RU61O2ha+S0gsLU6yP+F7troGDGXfnIgzLdH/ubBB7Uavkav7lJRyohCgpKC+Wps
XuIedCDTq/98vOuJyOdAIEPN2NpgYe3Pw5ncg5WcaltVJfil7REaUoeu0KHT0ZYV
BlKwjodrWu9BMRouNVH6OweyPb9Y42h37sRTjXG8YRgxEhr/IusCLm4j9/JGxk7V
xSBpoEpBTvhIee1UgrGiHfvWApmNyHBNQgX/iRs1VRSyqD2NHUiWg5fRlZHRYlM6
4lBA4wBO15s/D6qgdbX7xU5GvFhtmjWjYeTHhXBav2poHELWwugg1vpQ+QsRc/qX
LFcyAq7qNx0Q/0jxGxqja53liFTLh5yzowuei3DXZf51Yrel/1GrgAa25CysIckE
O2V7qLDhfHkIcVgGI/SmK8FBTM8t3SaP1J/uMswG+XammY8zyc2zp56jif5AXds+
0NGVpSiAMoJJEhzumNcVpK+iRe+WPc0c5Jrgu3lt+TsPluZHOo4QXDr/O1KWL9M8
xdk2MfB51nYMQYN5K+SFsnPn3VkuGrtrP536fJ+iaF6VQpooCxz2j0KyqaEVL+CO
XPcGMMc8BCRS+H1UJspie4vJXyTa4iDjYCgTwxCMVNXtDyJx/TOjkXX2hXfbO7Em
xMdPAaJHE5fShuL/zpCXvCajYntrCZW073mSt/bAwdU9WRFLPE7GjajiLWwD2apP
p0J8XWrVLbWtFuw963kkJ03o9AfptI0fOradzolF9PTWkCVt40hHCgZtfDViuj04
rNvqOBpWyaSuSW5K7/s90fmIRWFD0wwP3f+pzmx1lGRDEbpfQDsWqtedBJ5Tsn0m
tenbFC94b2ydmfBBiQ5Nqtz4WkeGWZ3MRJWeYJNwTY5QiyT9oRK6HpVpGtic3CIL
kgdrBp79sFRuLXdVXc1mUhgkR9Ek9FcrVaJ9+dEmDWttuOmlq6rBO3qeh96Jb4Uh
/buV1nMYwOyolgP8ow2/PP/v8D5XwkvMBzvhwthwVXj53mIcK1BWKFj38w1dIskL
LpUXJBb7h2rWSKPLLJecbt2kOMXIyhKNEDCJmyXun46xevoR7DP5pXhgjHhnRiZ8
y7IujEe8DjRsjH3nDxMfSaAlWTmXoU5b70T8GD8iVc9J2/ubRmmLR+Y/MadfBCo0
Psoy2RhQNjJOy9pGHhc4sGEnCCG+mkJakSpGOxZeB4SRMJQ0fRdU8fyHZOxTXcc4
y665SBdZbaTblbwetckJS0KoE5IZRDvk49opiJAi8Y1r978/t/Vr5D4OCrkXsWXd
7l3hyo+8VZavwJ5CPBzbMx9V6sHfiqpmbZpFES9arWl9epZR9KP5QMhyhQfwWIvL
sPvEwY6W8PvsUXolFVs6NQ53NkydzObPxP6r0vdABNjO1e3dNxUeNDRctQ8lV2nn
fYrnoVpGS23Qh9w0342TUNBC772hpxmKMIiSHN4Iv/h1SLchvnspDXPkEDpAgFno
v1vx6L+y3998GBZ8BFJWjKc+eNiXtQoiQkqK1idEgmlswFGGl2aN0vGyXHyDi68q
vPedo9B1JIyEn3mqUGTR+Pc5HBfzgWw5QFKWwqUE/nfEdCypeTULyCNs9wjYxW1W
Og1eErF3UJ1oD+WPsFgljBOiPKYELSp92ia+QdPmqWe2HosN6frPshYYIDzvsYD0
oVtFVLX5I4BmIRgeG5DscSQIECrvNLMKpPAe/TIT4nYos4dem9LpM/eA9dncBDK/
DAmRZ0IAxwjUvxnxLHqBDRJuTqnsa37lROJTeCWsYFXikpffjuWKUpPfFY792DAH
LITvSXU+CDBOVOmr3svV2KwYTeuXmMf8L+zQaPCOmVykLx5xmchJL3aEgtQMci7i
gmIcIqqThSuK1N7mB7jlMe/hoI02fIOD7tN8kal0F1yD1/hLRZiG07MhIMZD//lN
svgHBrFSAy6h3ZbfKbN5EVxB17hRtjcW9r/eC2AD+wBE15mrEqZ7NSxRMZz+Jc+b
fDqD379mRxOuQWxNQvR95qFit7npYLAc3GKAgdG+YkHwUs2RQDpqLr8CSUB9hiIv
ZZyX8FflZ/mr6Inukh9BVvczYE51r1tjTzuY9Z6wVbTjhpT2678/rSr+bGoUmvV/
iD+Ppsg6WkOWhZHRGQ/rqJG0vSXkwrl9ZeKnfP27mDyRuphhfi005eONfm2KXsZA
bCS82I1hINDPVB8a0w8kyOfztfrRDiKHkFwf7v/DWU+218JvKhuXnvVRL14BwhkX
V4vxyvLz37wKgfGMg9vZRS+7gDzZNsXw5B+H4hY7nQD0BpNEd/Rkwdpo6m2dKTvV
3iaEDv9HYvhXLwafIGSS8sLqxg8uRSk67CYvHHAGdf8B+1KMDRaV05/Drznbm/e+
PG0lOfWpBjSg98LC4yDfFt/Y92qObUq5jo+i2UychfTWHdWwVsBb+LW2o0HjRdfX
kWq9kpPJ7b2IDiWPF8vhVLpUdW2KK9J6bAHcITNd1eI1q0YI8B/tQZ2+7LFQgNE9
K+Rt4H2FZSmcs+viyR0PTa424Ce9nEAPcp2ureEd6tscRjK+1PM+mWzpXUjmOQ6B
HolLWFj15hhaWCUU9k1ZrirorUMePDK4ba7vrVqR7ip58OwIVuUnSTZWAjW7d8eF
aswMR+1U8Mj/QbR3lon4YJOvZ8rl8RCcgwJnDmRhjs6fBEJSTEGGzHlnamPByLS2
xvfKv1g3K1jv2KCdC45vxyY2ctWTld4V1WUd0gdvZ6EIBNdy6BPzO0lwr+0Qxdav
j1lJmSleQBn+MEqGI44HojsDEg8clKd1UZIkUGaVMPMUIFhLbAz6SrVKoA3W36Wc
97dRwEYjSL07L6sGoLpHwMH1F06TM1J4kSVnDlbKmTFq8xrTf/45mt+CqpddcjdQ
btXSlGTAwZWeP3Z3hmpvkOAChOqSV2tj1VYn5pvipEy2y+V49uLLtRcyxkV8B8/9
hJl5dgASuClrlVonaTtALUL+yDBwBp9b2MNIecMnk+4qYprwjrMlBDyz1HZ4MZCR
Kylbm8MYEeEciv4Ugx1peUFtHDVvGLmxXQkSzsOUiOmDpXn6eGIfczBif4Y7VGEW
1eL9uHYcNh2gj4/n5pSCJZbUyyycNntNx6s0cS/7VwIIN36hlVIE1xA+QSzulm0f
Ttg0H0CeYjQL5fFPcGNmPqpVKf5hKWhWo7ZcS7oTUOnLoqGtYivXpjtzwJIXlP2m
hEi/gJsXMwWAaGZSYcXL0XyFuY3CLJpxbHPJsezg4g03rF/zM1c7au2Oex2g8r6w
Mr8xfTQ2XqHBzmyJFRaYLSt3T6E5fk2dzcjWRWF+veqEXqZLatOk69qP+SUkKQi1
lQEjOA8zIhov2c9qXw5O61GpIRPRV0Y0OtDrIgABAL2E5tRO/TtGbB51dqP5/6du
6ZUizSXkWUGIHWm6BZwVU6RKVfDKLnuYR7aDKaNfaypV2Ck1zgI4j87Q3hG4x5tG
bGFnx4qayz0ah0Wc8CfWClDdOh4xFePbAmiThRNIL4dmtRp5QdIihU/8gZvEniPS
5Pjk4x5sZGkX4cU3r8buIqJXlo2DBv/jCu7gc8ExMmrpCMcN2yUKvZDF6bFJ10J9
/xWKw35+3AjL/TKOcOxyJIMqtDavFWCWMp6/pVqc6PkJ02lO8ma1nXMdGZrl2ogi
U1lvmpsoYPRJC5fpqol4tponvoGEWA9cDSXfIkY6YNDAxj+yuWgibaK4DT+MeuaI
uflP7IWcXMKKaPCEEJzOhcZO3Ueb4gkiYFLuJsdcKzz0SbUj+LVG0Zmh/Yn9rsOT
2j+oChiSeGPnsRa8L5rVy6gR9rCrxJvuhSHo4mqidFJIEy0Lfj6G5wsNehBaxyyj
wwPaAwHlGOy2D20EhmOdzhIWJCD3t/ZX/APsrV0T8kzWRvl6QR8bCUHb95RGaNgN
7OTKo6cUqD722M+DCj/Y/KZ/W4TBPAm8QMfyymYEcgkH9XWAZLz0dBqND0/Dj4WN
txXhl6TZB6925JuCE9xOozqxc4u5xESVhpizO6HBXmQkY9kVBagPIaP6VmCfar7z
nlrRusOmnAV753ZtJwgfhblGVOjepYFdJz0OV3EKBdgIQlQYStYzKP/QpvEgdElQ
EZ8n7tCfI9cCcNbtWDHHmkqXPsv85yjsdLDt3ZqU6qoeNM9W8pu+jRgXQ0tEWuTg
b5U4+V0qjnGzy2o4u9HINVDKERjolDMKFCqIuoxRnfykwoUSCaJxnMJMxa4pSr5Y
CMK6OMRZ1O+DZd0yn0eZjX1wPJbw7rUKYQs35dDWkl5dOqpYchvE2B/rZEvbULL7
JqAoCkC5wIvsfmK4+FRH/lqnHV3d98+iNoTpmi1h7vseZRYCgqUkpcfJhfMJgmsD
5oJF8hf/4qN2RFt3Lc4Zf0sf4mgEXiUXme3FEwXjleBFjscXdBKbfVbMVXNDHNAn
AKEut8oAoQFNnaJCUgFatW7MOpzcBu9uag8/7JykfyRJeFDu3lABTd/oAwkLVFK3
nX1/jCrMZhqWV+OoyytEXGHZ7JfRLzCrz9hFtxIGwb++XBfjbulsxNG32/XjbRQX
A0QVg5wD8qa3n1DUZuO23NdMtmh9AW5G67351nLP2WbVeuWdcIx6EAPQg23pspO8
kjW57kPg85JFP+7/nlEJbI1ic58Psz2K1SUrF4V+kMGo3p33MkuuOFynH+IuFHsY
oCIs6Xqw6udLSKXfPhSvjO/WBEuAqnYdphU5IZjusYnCgmRXMDlwN1RyPWpHresg
ClBOdOzgTJmiSJ4QUd0Lr2NQUgSw/vGAQCMg86p6X6mrln/J4pa4cbhEZgjO1CG8
GoExtPXv5x+UFOxWgMIhY5g86RvUUKJpkx9lSGG82WoKtwXkPlHGyMchZu90HP4e
cqtYBkbTjbnX1eLgHPbXiCtMVa2qFxhv7GBVXKuNaEm9rsx/LuBPcRSszovd213N
jOyAd37uyhbrJKbj99k1Bec/lBnibfMV2Dwt+9ftrfKmPsaWpZNTtK31o55sVMeJ
C6Guw3JjYmhIuhvK5dzIU5uifugV44bQoyaw+iSnBXUdd7IoVYuoURD4GZRPRA9g
4yoy+7k06JT7J8L21Q5qMu3m8z3NVQ7aBHjH/zSwh+5sc2e4+xBjzvU6qPjQ6rVv
6Tfi2s6u4Kj2ddJl83EivG5LfgHu01qzz6bPHQ9IU10clDDVcHjBj11oGUIIXJ5X
+LG2PW64eZw5f4ofXIN2Xu98c+A9dEAvlAOKWlHZaObV799H+zR5DCWUUcLtm8sU
J4W8wfVTcyf8omDni59qkJ9G5wRZc1zNwc6W4fAMwLlvQBZWxkVxBhoNlyWiGxLU
2xuNcuT+FjaXn234/XARw6RFiBhWUzJfCDGOumKWnk20Lp1mv/duRbG5y538QBNm
koXQJumxf+V2vyKXBgHjDtDRI1Q5l1bUf3Ez0nYp3XqLIxDutnQPyyk8uEDZ6sry
9NpRfXYeXhaVN3lGsZuyrUqM7Ys7zZxLNm+LOYzntPlRNE1hQvsjviDrCKmMmCcP
/s5LOxt+yEchFR0XEZwUo2Jlx8FV1VJ0azQ9Q0C8A/7OxIwSyclj272SD5wD/l9r
ne6yxdEvQEUWZI4NlOjUFMoJ9ilHnPdmqWaSy+C2c952egsfb4j6EBsPjIO4EBA2
xqIruO9Jr2Z9clMnAtwdEmcWbhK2PxmXpgQr6ewvovo0MTRx9WEV6a678OKRF7Cs
SxAUO0NND3i5uP8W03BAn6ymsyo28jpvwo+gDzYC7Vs771MMKruIDgJJ21+GBgkG
aSl9StNuF+APkQltiPZJ28ooB/0NuinvvFx4QczSV94uLZA8mOxhfhd8Ca91S0kc
ZgkJ03rbH6LYJrdto1zZCIYW1JyhrNxXQ4MXBK+6aI7zRPEaLoJF2iGr78WmmzmV
ZR2/Rv4+d7WgtWJjoiZkaCB+2sx2cqPBUEgNRKkmO43v9yk5kTmYOz42gCRD2fJA
uwpfODqLGuHiPq6GiyWfZHatq+pEkhEcRgtB4okKbkgCjF02s0ndQY1YZ2EAJ2z9
C3tbbDgkJ3l9hWFv5eQGyQlEI+jwuXYTtrO1Vs8BiaTR88f1Vwd+FYteia8hsHqg
wEewdX6qFlAl5GI8i5lvW/cU9W7mDu19tIw/5QyGkGgeYf0OTMCHVxp+cKtSBEMJ
zfqgRloarq9zGDQitQ1zV9ngGGWXv05UcVahqK12CJ+4/G+h9cWzRPwu2DQLqD0X
cyJAoBr6dkOFoR21+Yoo2FxWwylcEeCYUvrNJ1kVYTLFBFFk/EI8h1k9AQjIh5AZ
uWhVcZq7cvSyUf4tX5VgkbYQu+aoM0at0XttcPjSauK7ucoV0wpaSh9ZoXX9Fidr
yPveLq0TEK2aTta4owj1iQ279B88kl50+bUf6I+rWdxjFVblcUSoEhWJ5674zXOq
zYzHD1asglI5TZKynGmxnlXchNPrsGxK5ZlDM0ZSVoorW8JEg3vOsMREnRyXwfXA
rmZDvLfbWs3B7d+Os59BI6gfkN3wcyKE7LV9wv9qYbgVZO5j1DdIG68l2RZ8IbrO
gV0xlWRd7VxvnnWUQbjBn60vgcDogOz2tYU/9lkAGwMRH1yBxoZ/UW5I6XzlDOLz
12TEpAFBb9kZ1vYpBOjfvO7xBIiFwVF6rTWYhml/Ft+vZWbtc7HW5bzTk0u1qh7P
vlz3jVXI6FRqUyzAuKX2XfgxKbgjFy/1VQhAomLeZJwLI9wWlOKVGG482YEC1xi+
KhSG/mE+CcSkwxlAfE9EXkffHCwgicR2QueI/jAM9D2rP/qLnBOzD11PpRg5nd+Y
72gk4Y6Hr/xOvI4feJr5r+iJrVw399/5cHdkWAzmtGCNXWs3G1abWzy+1MS4gB1E
5kE7YEelCFpdlq3XS0Dunl0kUcKpUol2SSgDVh9CzvYbI7PQdr/KJNoIHjK8RRn5
mHUicmoTnO6heIrqmlgYp1ZHrdaLuycfbWySwlfPfvbnlBLeKutjLLBuwVzH2s9u
AK+TfL+K0lV4lOcpK3drwq/oD+kNOGxjLwWrOyVg1kNzsQqoTzEHpLNMEjyOeutu
LePxa0XuFdbhfDLOhmiZhjANKC2GNC9G64JBROQEVYdyjceXu/ggIOU6i/c+QUys
ejYE0pOAiMmDq03Rooy8J66ojTVmp6y5vqQ9rxxRNKyj8QHu1lylQVY3BtAblPYW
qi4MDAiN3YVTfr3ItcNbgS/4ugUUMGKPziVmdBEAA33MIfS5V+PF6yIq9HaP8QR2
dAR91Fpdk077eyNn86cm5prDN2nXwRsnu3C4r0TMsI8cGJBhSDTy7sBDWyUILGYy
Ea1NDhgRvZj9x+fVKfouHNiPAZ3m69gWXhI/ZV6fruHU3uL10TZwJwIBXa8BZwMK
RNEniQKhpDky3GRO/f1cJDTc+5yMAkR8Vq5xLwftIPrMPM57mF1o2Dd4mx/MQ3nT
e/lRPvjS+C4DwP05Ur/2oTeI4YO4J42evTKyKpY7jI0T4/TTP+H9sx4zIWc+I4Vf
hTxiykZ30t2AWHLDFLgScsEdxZNj5gMSyg3xBvcxkCFrhJolQS1wkBAHA89FYk2N
TYVz/fVS0LXG64WeQcNkIebEXTN11j7ZuW3TsUhGRaft4Yg1wgtyq3ydQsnLdQ91
Z9oJmYglAvwHDKaNyfi6HnuVSPSWjMule2zkMeDLvas+QpbAyDqnS4xNe6YZmWHm
qSVLy4xSnzYif1Vmc+Unsov+kovOOjBo87+HVBcBYv+70MIuGSgD9BFRh2QhokzO
Bb7csBknWKHSYGXKlEiLJ6AMe3x6hEMlptpPTQNDB969leXM1rBDhp2JXlRZZiDo
Tx4v9aP0pSwZujKw8c6h76+3QaHgO7f5oaWeqJ2JzDRNkF+EWe5ZUMF6ZGZHU2oV
2/49ab8jDB/k+z2B+fCSU/UaE4iARE7zZUSNFFLTBamruZyszI7HRRFxhWbGvMjS
KvWlDL8BpKD9awF/D2RL+s5eokYw8SyNIApzK7/En1qgGiky8I7E6e+DELk+8cOk
M52GpYDwv3u5vua8OTfCKPnroeaDdARhrgdYyPY770EGCzyeBBWf1sjf012y5gMn
3ngg2XLZ47D9wXrvInck4gWwVvVuIGquS5IO8iMjF6Pxyb1vZ2KOEn46lcWp6f9j
7gNEPosbvYWaHng5AF2G04U5wyH4KoYzopLKwm8AY2JQ5ar2NYGcpoVmyVqxw2ji
G5airdZDxhDUZEbATtKWfLR4xquM2LMRfBe2HV9nff1/8x5nhLfhzdH6MhAmCKYa
v7824/xsvZwSJAnUe+5mZqvLLqh29Yf9zp11WTY0Z50qRiumkNN9xUqdgASGY1wO
ddETX/LdcTn0IieVBxLktr6Rwpc8EYkBa0jLMfDsaDhb6bRzY7Cp5zbP4VA1v+m8
wAOexaJUe1dBlzI8GIz5++cso1pHK+bvXSp8Q6gY/6GwUO0Tcj7UoplcRpp+j0lN
m0bl2slCT4t6TOtLDpiOHmQlgKoCTKqIAHP9EVubiur9uHFFFcZSnVHbb2O92ULU
FQCf2WjssPKZy8D9xJG6V9zo1V/e9RhD92RFDBc9XTwWlTkeQ8LrEwJGouPf3PYf
9XS8l8b27FKfZ9bALp/Paao/gXwthNK+Dr/gQoAQx5BzUdjkh5o9UINl72YfbWG+
qGC0RI+nzXojsdJ+qhDd0cXVzss+XQI1E7sHcF6iRzTvYoeWEaNab3jNJ1mQLDZA
f568mSIKfdblxixMHUsOKYE8nHvecOIKJDtkFvplqAbf/D97URLgIxI87KeBYtT7
yTFsxryTXULIFPGNS0gIczRM51z6928zYvEY3rTDNQ8MezIeVZ43P2JroIdVe9QP
q6xr+/LJGtVld72CKDlaekU3o22rU5OdtHXEs8WBkXKBAHjGsYLJA6Sgq65baCrv
iQ4a+deOkkBgadtonNEdJ4USA3wJifSkXS6LmpIgYHbaBc76xMEZBo0q6LhU9RRP
IsHatIaIMlrWxOHxbDys7fKSEFCiZuAsyH47QaHFo7tdDk9/TNBhiWfR092IYQhN
64nlA5U+oo3gQ/vdWDn7gxZ8uCQYbFuiA/qN4h2MGNRZHdVBBdgERWW7nPrUiIPb
vIWu+ILiOA1oejVSWYSNdUaL56DUwQH8+Kqd4hn+uInz0do6tljjZ/n8Dqg3xFea
ze9+G7HFbkA0bCY+on8ZYngLK5irFC+2HrmrEcyz7dHBAYTAzQ6hjN2xOZs/c/S+
IPPFfkKuhWyS+F+rJYhO6jYPU+KlgESUvixHJrgJSOtXwJn/rddGx/X1wh042N4t
Pmv58RSb/8FDpqbY9R4IzW+gUwJUsMMZJh33YEMSY9kBlPuM3dIvfxRy9TMfh7cb
uA9ZB8i5JkZQI28dP1GclDfQqLsbRH+xLpL1qmBwQG4xVw+RcvRzSf3AxB/Brh0v
l4OdyJdVoXYHy39URlqndLhim3jbU87/zc5UUPep2K6Rfe40rx6II8ZpKuGD//eH
t+Que91iepMkZZ3Lk5b9d3AIpmRaTmBfkpzBqMxV1tbKqshZbB/xU5nE6PTAPi4u
AZ7IAjn/sCrwblGXqIV129q9UNBIIp/SQ5jnbrz2NNkg1smqbPdiezd82KRp1O9x
Wt7KH6sYrZyHbf3LrAt++BWRU4Jaf0PniAXHK4iDklWm3qJlX2tijYj2LAlCMsfI
MpJIMDeKp622n3qouSjEV3fbWB6kE7+iiW60iL0F2169VnN4hRnt8VGMUyp+hypP
W33Zh3K96X06qxza+6GCKZwtcNd+SZ7XaDlvDUDADNe9Ncb9laiYkS1709iMZPZP
i4dBo9YK6NHBmKjyiVCbpGBpZVSr4vJEgAjAiwXlkR3q5XI1/6SCg6w9KQTj7/bR
xJiBtrxi8/lK1hwzln9h5WCVamyObFhubxpEjNcckA6zmSmZbzgV7dQ8si0CPxwa
V2bVDHgNBiEG6EqtJ1/jdXg/ZhQscczbhuau+ytPMBZAlVoWxUPnrwTDr6u0oWzC
iGZv7S9LE48v9OZi140j+stlzXC5zI9fdSgtvscOtORyEZ9osSj3eMJaHQP3p4uc
lig7UNlXjzTWnecs4Gp1hNvSyZZvWmDQs+9L8d2xinYzkfI6+nlaiQhn7V1pzShc
fg7x6KjHMnQOLPEmn+tBAOGprrdxRsdC1e+km9KLYymXQjNH95hxaC8xdQGBmU7U
n7JZHxS4rzhIOYa4JhKwq/nior4NJjkwOzByfweqFW5O2kSke3g1CI6z5nuUXUKR
Y6skK5oxH3RgITrnmbyy/G5GFpk44AsQAOXOvRU9PJyo2qZRHRX+SVsXeVhMUC3V
UYqk3A/DZHZVwBs0AGjYxfVB8CnH6JmpVX3iO0sunb7cTVi2H78MyG8RTjmhDy66
3a2d/nJFniRMNMhdDdEowsKeWQcAKYizAUKpMZKvogzH69qXZcniJv+3cbbtoCFb
kcMQVxKBb1S2S0f4MNBITzZX3CoNMrg0xlIakfWlaqi4rTmniliSfJUBycC9zeFH
duOUXWmVuSOdVq09KH9eBFiWpEK9AGJD11nIqPRayof9tF88zOJyBogF0m041NRS
0Q9zne/qGODmZl2uVv7E+KgwnfAOiJZwr7pXi2MD776U8NIkEH79DtMpZFoJv/Rs
MfKLA+VJ1+CGi45IKKbyQSjSy72EhikbFOu3agvW3YHQZ8xHRgj5JUGgLemc6tOK
0MBO/qLNNbbr9aIe94UJaR0u0Xg0rgYLE6/zxWhjz0dqYpWhqwdb+AzSXaEQIiiB
y1Tc55w9EqiV+tNgbYhgI/T+bhy4TQ5nge30ehu/83DRcl6beNEer8fD1+uwawGg
8crGiNK6tT+Lk8sTjqK+hglACIOuOUQadO4BKdWsJeKDfDWqaENAQuoblmX8av3k
2bUNsmKiXB8mEfVE0jaVb8oeBRY+LOTyDwDAh0MQo93Q5Q9gIB6ahZoVxzJsWRNt
RdxHwaA25trt8umcpR37WiyLH+WwlDqGuUFcmTcHOyeG4vX34qfNojmzFt4eT8G9
WmymjYI5iQCSy8b6gAUlHyqu+SlGo5lZlht6DSZtf7wdihzuas35iV93Uo8JksBj
qJk/HvGYrEuU92WV9r5brFzljLZZWK+a9Nho0xuNprUEBr5TCWyK/33MjiRV+bA9
ygYnOd2Ykcs1vNPCn6Wu7uF9RbcxTeJn4K1mEKQaVf11xhtCyeG3pjqglss5svQS
SX+HRSVBJeHPtc29jZbFkyVPwTHlAClYKWfGdw/oJLA38qp9uyvnwi+sLmzI+Ckd
YeBXzaVxIErYlcQnt2/QP+NTYjaFwU/vb3+jvTAFkmFtsC1cDM5qzXMmDFM9uTDE
CqEAVZgkgTtqZxkXribw0OGr1iDnk3O1vLyz7HWZE+n//x/43oSlZ6d+okJDqxXk
5GxrpoNXrtD3ltsRGW/Fp5kyUy1btwy8w1sD4OQ+YVuG93qEe62Y3i7Bucaq4XEa
+byHdg1L0bCY4+kLzVcGE6hCHxhojOYejaBwXD+mcalUfWp5BiqIIW7MT4v/IP8x
2DqSS3997LflF5QbfIOTGSnjdDfRm/HvqhiWl3OtJ/7e+n1CjGRtcivATbXiJ8DV
ybXz5ej89GH2lNUCys+vOLfRFSmK8c+lFMZIuh5cR912E7NALaeA3W0Yxb52V7o6
ELehNLjD6II7Z45KXeK+1a8IwL4mUGJ2eKORZu5AiILdw76TakexFcLy3lOuG0fy
+ppjPUMO+R7eSB+pfK/8pRCsBYYpcObjgI/CX8E4Jxar8ebgaEfAnzUCYar7F8dw
Lm4cW3y1IpxAY13mIvxcP7enIhBA8p/u73reO7OnMwaqEdTEh0UErnbb6ztwMYrh
Vkm7ByK7yOl5k2QOjrzhEzO32v8k7TSHpa1kfh5X28FgZBP6Qw5cB880xGpImnNS
mUrMk//IZWb7kIzbtIkrhuQuv2eKJwzyiEbBoNB9Fldq7Pz/iYoNv+Ky5AY5X2zl
HTAiK2EYHYIDfKXcYkhLPFVBOlAD3WpqhOLqesvWQryfuqfEQDdnaiUZe191ViuU
HmnMP/dDgoGPxs9lRgFW74MA1v0Ud0epIu7C6Fgq+XoOam6wGcfYCFFd6FNpUp4P
i0XaJaJDsOLLBeMppZ3JgqqnFHwvOstu7uZgMuQVa7uKPG+Z/BMJ83iqcH2/bmfc
EW+uZt+92ogdhThRuZ5ZU7RGgYO0+Ew1O5MR2e+EAVaYS3ELfvYIBxiq36whGjhh
Lg7hek71VWSOAmwgHLKx9bhosV/MDfib90FVf9kX0WDyAMXrVYjZGxUTHB02EbxT
95WExOvlzrCwe3Fn29BiTlgNZbWy0oydZuqMxpqg0neWe/pQnWzJHxWijENfsD6O
1/3Nx0UjT2ZAGCWy7J8kIoZzFh95WlDhSZpPyL1+gmretQtTBGxjQZgIj2Fs+Pfh
7vcOJ+5BETuOaDadpgaVQ2Zib0XnqNzBEppZVjd6l3Zih7so7sTNtxVYki8k3bSl
KXAY8wlYfe0MIfL47ZKiO4DVmdrwXCGS/dMibvofNIJX/lMuqfmqNqKlKdaqnPOq
erR51BDJm3knlq08g3m5yaKxtCWVdy3ZR317OVhTZK7N2FW0iroj3nRb0KWpgDJ6
zVmGE7VR/EstA7e19vfu8bzHGewn9749D699kMrZtX2o/ZS2tHmGjHruH8v4M/U3
UZZDtf+fu9RKqQMZW1tnFiN0gXidMWdegUvD2/ZTAnwi10e/NtGEaEps9TZvx5JS
IckXmAxydnN38hOvM0y+p+EUbaLAQXuosGBUi1+7qVw+B2kawsBpKNBeSX9GIwBy
8cUQFldHJ3hy5wE04CdO8ThW8Hmuwlg8w9cHiwhO0Juejd5QB6vS+gq9K6rDxIHP
QUqYugD2VFzys9hKOLLe5fCBn/9ZSMN+DdI71QbJb4OHsBVYpaHWiTzvIVryEasP
zTk1wd3JKtgECA52kY8N+qPcgdM8mvIPlbKCfTJXjM5FUl873xaH7ax53ku0xePf
Sr5cJNrYhgEzwsbn6e3B8KnWUjcsgEJNUZqMQxkdiLo/x8beBcEEVZhEZBPv0u61
aAIDztX6UizdEiujVHnBYJ4T4h+8H28E1BU1lZEit9Pq/zrRtdRGdrsMWMAteSRN
DmbXbrPXBCJ0tjNJut2SiFNHV4fIMrmK7b39bTWkUv4e2XbynTtRs109T29BX8z3
vgNnjWT/nACNXQrB3RIajKlNILq8AcA0yDm+jJur2g/fp9LV/hMyNgwjrhM2Roxh
BvbUHiNa2ULNKTNOuhr5jynchuxDhwPUgO298ALC6QzDQKFDS++qU6PivyaDA4uk
Ry5ozhEL7bynGQfx1JLOcUpkJmuQEdM15oOea1C/xpnIfo69yiF+VmWY+9vIzRen
CRzyz8qGmQy5Fl4My4ZApjIUUcsikjtJSL5FSvM86ziDG0J1oJbfYBe87O0783Uz
ig2ADQtKAYIbsIv66Cz7qTq8k3URJKRY7aqPL26pafBR27jFrYEfJceceSNm7agr
e/cXe1UzubLZUFdaQ5cbjh5jO88o9QCp7Kb5ySRbr11LWOhZHLpJ3fhuOvpgYWZD
ZLcDlfTXCyTMcuJordGb65FMQvO+ZlFkaupEowov+chor8YheajXxGT+i4lqL/9+
fEAEEJqs2Pce3gMGkiEZUqfgXlirZkxw4SxlfrvCEH54FvBT8WrXeILF8m3ESSgK
ObJVw4OzeooTtDNd+rrGlbp3Oq//C+mPqvLdpTpXLj0R+L9MHVImhW1RqHEV9bbG
YKdWfFkD3agoOrRp83xYVQjBHjApiiOtD9VtUi4tuWpsFcD+qtp/Lh16KJOyZHRu
MW1Q8SD5VJoyunuDOcNVQy/e8hv3UgvoH6iqly+v7AbfCkOmtuJIvoN/JEF9xjwS
gkTyLDQO/P2ODYW4wIxMt28t2ChYcYuihsozBEUfKnPXvRQA5DMuTyBLEPrL/MXG
ISfLxREnskpHiDS6DwRmEkt7jzW8Vr1742yzDnUiLH/GnbKC8JPn4STfdhQUJr1O
WKZI+VUQ2Os3S2OPbYDx6W3K2gP/o9u9nZoag6UfiCMvkbdeXt9XEroiH+0PBAvo
vkrlTbuZVc2sDI/UfuvjI6dKDP4pqJ9TAF0SIzPOzWgXPugMPaiBDzWaYlrDzP1r
QKpkyxDvPV0y57TiDIvXmGOYhHkO9Eg71TZOq3XH5hStJIVhQnqNLeMY7Cv7jOIl
zoJgVXzZXsvzTEU4XCQyufVlmu7E+99ciYXWi2AS2lhK4Opx5By5G/10G/t23EhU
izEBYhUqFUm7SN1oG5+odHuxT5FhlRz1aAn0NFcxyFurtajU3Xt3V1rcS1MFVyda
ff7/ng2ftW6NBIT/VXrH1Du386V+5Lzi7SCUKWSNxbr4muMDVclFy+pcuT11PK7h
zEaRJY252vHm518/Wmlu24f4BMKgy3g9hJZHCJVOz5RTPKW7nKrGsgooDns9RO5c
59VxKm6ORnhFhlMIOVeU448wxT7fvf2j4eCoaoSPRho008aFw4ksbG1RWygwV+mp
iGTR1pZIGniok+GD67fiIZYiGWMiPAkca67qnDjj7SEkB70ikXC0JNB8DmtoFk3E
dbJI7B8vKA23+RdRsLqsv5aSg56iTjdOfaUyVC7LSTUUJq05aWkpoqzglpQtERQo
U0dRCh3E86B2Fs++i81hKB8bsso1TJ1Q+wWfLTCIAEsem2wJJgbEdxwqpOlZwpQz
CdVQwHdoNOiTZ33uXiGVrCNcwgrQtWWol3z8YBBl5ppAQ43yIf76tkix34ofa4XH
Mg5An9JcLCTFJumwg0b1YLoZK4Icycir32FugfAke2k34mLD/jX2gwKp+4/sbnq2
GEgIBx2GpsCW6LefIm4iACBoCeUFOyir6/jlg8FN1622g3f6S3toSzhtwh3eVm6G
OG4ZM7TpuZvoO5q2eszelkZ6jdScd1RbnVgOwip8D4lDu3BPI80X7r63I2UgdrBt
KYUJA/uZM79ONmAZmZJd/LpY2f/rRixmqkGbIoTVon0uoqCT4bVCLYzGtimOk7B9
ImLg5FJ44HvrDI94CCZE7NrDjIkG9WpSzUdnEn/1ZLWHhrWgBauhZKYmt0o1W/+2
SpFkHRyu2sptn3Qb/No1hy967kovTeLw87tAvSLYVIkT0TlgltN82cDvs0XVm2xv
I+CE4UIY8nQFHNydDo5bbKRl25Ymrp+r7oViFeROu1Pct+Hn6oMOI+vG0p61XtAk
uGO58hORwevizz1x4ESFk93wIUpKDifAWttltbftUcAjfJXkUas5u+WTh8i79F42
VQdWfOTTQ6hyI8aVoqXvVRLtFVjf7mhPOaF4KFr4qxqC8biiEXSGWOmMTRT6Pys0
U1JYs64sR50bgAgzJMP+89Z1hVtwSiEn9xYhEq3TywZfdhhB2OWpUemsp60CDxbM
GY/5T2J/PRMw+8UUz3Ab+v+Fr8MAyNAwc3Ic4DTNemmDw5vo+gMm45jAfvcJnp8l
xj5LAznkwPdtgXY9QRfYtefBZXJCjjPQCXAsfAxoFuPJAt2RFx2IgsKKr5dpG/iy
AfACK8Hnai/+H2Dh7KMcZpZO4X+torYpIoxzC9crMo5i8liHm7oKMPMvmYHPraiY
5FqkDmUJ8DtUm6bNMP65ZopDrPiWuWUECmjdLpApM5GAwEmMH4Hsshp7/ceVQOau
vzxheML9Ih2Gsf9VEI2ipMvDSHBr94281dSmtCC1JEAcOa91z/Ru8AxSYnP+KsyJ
TvUoFteFYqX3Sx5DtT8zH26ZSVfYQvgUlpLbxUzmfn0sdOCSOjI5E0w98BCgdwG9
uAV/SDsl3V7ceY9oK+dlqHUL8HiFOLeW8PTcJNh4JtOJAGSLGj03O3AknJkLneni
2+8zmawRuH0RaQUnNSV/sEV8qQSz5mXtooHqwNjK++G+Jfelk7HktGtZMYN7o+Fo
3y1ey76oXR5DVSVK9AtwMjfeG+8LrwAy8zhGzJjK7ABtW3Fp0djB6Ktl4A9Y4sWo
xpOiwlzxqzXhMK/hxU589Rvk/XZEEQ3wHD/xU73tCUCZkiSGZN/QUvFFWdb1PwCB
/C5fSPE/OZNZgQDEQjqVBAX5YmX+RQ5aq2ZIrJGnYcaFnOtmIjlzI2RXE6neD776
BrThhOp/SrsNEq1dAlgC91gMOPGgykny5saGeHB3iBgeEFhk49amN3bcvZ7TxAzW
8ZHTuFmZ6BAH4PRt1EIdk6eJ8nkrOGcc7v0eIKHYx+Qf/xsSPP9bJy1TqdyEd8n3
WytCTcIW9w0sKg6pVEzMxlUoBsC7/tC5VTNLM91xaqNslh9ENqjxdIJE0vafe48m
9mWHXG80CDGGixytA+HZ33Ov3pgjrLHl8s2czHk8qHI5+5aspcaaPr3fKxdAOB+V
lhbcS8BvS1ol3sPgC7HW+i9XAXOsbJ70PGSTMQoFG/3xJJqEEkmXOvoAH/PcXzIM
bfVFFjsxxm5GYsEWH2OYlXdW0mkIgAh5y3/qr2utNo8veI+W6Xttm4EV32HIjplI
2DJ/Sy+FLj284h/akffeoO2RMQrSVNS/8iXPi//BF3Kx9/1GL/JZl7nVZpkG0X7y
0J6HeKv+pxq52klZcBK5BaO+ByVj9Af4x/+VfnNfgsg4v1PIrhAqXG83ZtaKFxqx
znT31VsmE3fXf34LiCqamzRQwY3RFClUhj8lTtSqxtREIaTD0uf66aZeo4dh7nFR
nIDz8oMaezopzSv0VNC4RJRkgwwLSh/xGysPz2o5pRctFbZClqMYOVR0OpvXADpU
5AxTcFc2L/vTPH39S+KbZRjFIOxfS0nHTdasAMhOx88VxtVi6D+0cgB0MxR4ksPw
kmb9KCNajfAMns4jyYfpusejk+46XnYV0tDkE7LDODAp98g2cHAcJlxnpBd+g3Ea
3AoQsLrKxJYFCti/0Xau24QBmN4foo/Nw/Y2gO7x73Y/QJg5OoPOgOLyMu+bAg34
xB7sZScoLcCKPIwoaRM3fqtLIKySrd7/IPz/8XsQbNqXVGv7MOafrhjG7xMaEgVR
eUY1q5gRAecnI5UwIsB2z7cdOt3OsM43B7KfDlw8VGCqTGZBxwDK4ChAj4hGi8KE
5K7j1IyX5KjyhlaN7wWmKJ5SAvZL2RRhZZB5/Qfdnp/NYk3EDsiOQlhFPsREkaks
3rYSjjvHp+KYEH8GIYhvfMm8XmJTHIiotcZX0BvqiRDpE6JjZVHXuNDnKT6XWWjS
KFsIqxNvduVCcCq8XqsJYcuaZyWFVQW+GaI1XPZPu1mbd0wlwS1ZZJ3g/9TBLDnR
R1oByVuCUsI22ds6UmgPmtxU0AJ5S8mZdKeHZMIr0odAbLpRSd6bKnTMKOxvO2Ql
pJqHs6fBax9ICpPPDThmxzJNByV1X+0Ma2TqHug0tRDuXOE+VGZLjc12l6NDlsSx
yVflFetWD94Gmkrq9+2dHubqLXMJNeZBo7N5F2BAuRuEDSXeS4DiivnEFNHeb0PG
uTK1NFM1vI0ZDLUmZr4YceASsppRfy/JfZIQifySoQcM5vxO6HvE3wROaKUBztBe
ZvvIspuA3yAjiDHIQ3ODBFrAeaKjeUOp8vz+D4rAzrhaotvy7/Q+CijQSB/9iUbj
i7In1dg6Ycu2JIFLAhohoOUs4seahrLPhhvPMHOXhKrNmSnzjI5qq4BfIq+IogAE
7t4MR/dy8ruHjcDmVhDWrPZV/Eyu40pHt8c5hKC1Ii+mKicAc9LvpWaO8FoCjRna
xdhDL/WeocjmX/RpJEkMOxjAqgLnAqEayBwYbjvsMltPo2UtkyveEOeVcX95d74X
BEF0hK+LIlyAopIVAltOi15BOJCS89e/0J4sDqDyPBzB7jFFnUw1W77n2ndhP2XX
F3zaP46zlQkVLxPzMTEQTgRqSAGRIlX6T9reRECTWuEppxN5AAnkIem1VAtb5YIg
sAN9iKeJRxGo4B4wbhIaStjuXcL9Zi2TlgYMdrVaLytqUBt5SU0mFyGHREJzToiL
h/iI1cNtZPwKp9Vu3kJyyGlKBnilqKmqTF1jNOHPdS9o7u2Wb6YrgapMNoqUFIYM
zkr6cFQcqz7/5QPBIcznkU7Fmv48nxHl7KN12T2Jh6ss7+CNzA3KJ2NElWJhyb1p
v0DzZugjvECtdW2rHPUrjWFjTXvh7VR5yPy66rWidUu8+pxDU9lGf5zfOzO7KDJP
8USHm4APjnAWEoreKnP6HVNHgGKMskmtobJKaxZJ98jyBvCyW5cLYeLK0xh4fzYP
ZsHNR3KRLja7A05iltd7FhDfHFLJRJYdNNps0x23ek+zGZDwONM2lYEy/UoUhUGe
w7+k7LzuO9u+L1zAJnvx+PAdYQ/XNX3JbVy75uRhLcl68kyU7qquyVcOkl+jpUK1
KBkwgGLNtDumPyR+TGeAJiEYg0YeXWiaEpFVf8g59uV8ZSfcyC9jNWTbymG4Trb+
1CLeWHpDljLhgSjpgYiAbaRpFyUcH3TwnT2J2WTlg9jLGlCq/Ov1KYyKd5SYIR5m
W9bFh4RfSe7fSVdbPwcoNT7s/cPtgHoKzUegr6/oEbuU3zXPgtjc5WhMMmypBu9H
qYVVLRPT7SQGdNjdS0zu6zs6XazJ4dmYP6c9IHP6P7LYKRh/Lri4EmEDrP9kCpe2
2/xLbyOvXWdIzb3OSqOcq/4r30LoL6RqsbZZ+2VoCerBJ8o+7r8G1/i11XJU52SV
Ed4V3aG0MXwjPj35egH9Wv+diYOKxRYSu20+JzH4SFtNjaxpn/zIaIKHbw8WFFhn
xzuAzTlXl4hPPBqiNqTGdmhUknphgPs3Qjg/bKANFyj6vWL35rLH1wdWeK9HYCUs
B70UAKL/lWUR12QGpa8X4bQ2O85Gl6O6nDn+aqgxuEg+tN6mlcxMu5XBWBzeyczk
xKE555EGJnFgeyVmTC+sgKzrst3teYqJctD6OrTWdj5mViqtj58uwukCxJjJEJRl
Ws3TflgZqwrcGwRpapVKlfgINmebh+PPjSS+aW5VO4dQVUw1ewLJTYPxAkBpCxzr
ucT9fyI55Y+cH5865da8Sd7r+6kx4GTqBE3NM0zd4x06qxjHgvZabMI+KJFY+kFf
DzIBup2vnNTGfKuQ+QZxLIFhwejwT9XVmYnrg/5TlG/GuEFFuWJelAHA+oZVlAMp
1NGrrx3d/Q07Pm+ZdVQZ51QoQZqVVrJAVBk3uA/IGvDm9KQeUed9oIMTc8iiwcYS
qbaLkxv897YEMmTk3EuRv5GOM2KkguBgdJd+Hr9GVouoMp9vL/fHs2b9XO/DDIUd
/yJIgUHjIRpb9G0G1CkDhJpSSjb4P2vtTO0Uv7k45MVshhOlL5oCsqKtZCl0GJR1
b8ciuIfVAIWfmfjILQrt6mXvxjr9omOKF7A+HNxBcdMk9DMOKfVHBan98CBsadHO
ntc4t9ACUZEbfh/fuvC3opfRLLibbTLPgEgZ4XPAX8+TUqJrUUsQHRy73QIAKrPm
eliJ+KwC/UtzS8jh/Ga5o4DbBiqFG1PJlEYZyT+7zRwa9ofb1aimf+JtH3VPlRkc
viooMIuaQfI99AW9v70YlpHCdSdzHZ7rieEbN+ad8ly+NpuivqqtfQzLlxZGqGJz
H01+ZAgtGQOWQzcX5yygDb9Y+jIrVaIFpItj2LClEIBFHcG3kr2XIPkF2x2kzSGu
mHiw7oiMjf9VxHHn4iJeWQK/OEzqdk/yxlB74HxPtt4IH+NOMKHxcWfIsCNa/msU
T4O1vHgkAFfyMwCKzIJ+agESLgn8VQQrIZyORPqfF3KqKuMJlpSr/HK53kHbfcVq
j9EDEOY+c1IdT2/JEUlqLL7apQ1sXDAaq5KmBIwRI99/jMRshkKyNG9usH6+YLFp
xMTzWWS2sqgZoZ0YKcPeMWWc2kjR+rjXtWqq8RNQf0MOnbv6HlQFrsWN0eDA0p/P
ES3Y+553bakjfzEjONbo7XIZxRztKYzF+or/kCEoRee4LPpzvmjWR0ZPx1IBXMWa
05kVicPaAnOhF+Mk9UoQ2oUAyazLXzr4Gv7twZUDYmqWoAnMAClgphETT4e98NC+
2xdSn5OGP/mFhpZEaSXIuK4LFHENmMT1Lk6L83e0raKEkCM5IYW9ol8W+DYjVu65
BjKtKYT4KZ433xIpIp5PI7SQH3TcgeP1oP1yPnVSLDcKsm1TCC64oJ3oaTa2V3uY
JoUWy+/hiG/qQ8S5uEXBhubc/HETszBBNbQ9ja7DvScNe/2wFAhjOyuM6n3uhX34
oPqQdnk2gsQ0ui0DPGoBQpHcikVPLkW3Mo/pINLhE8A9zldpbDifx/KnHEMO/Z7Z
tIZtFtb8ImPmZSy5x+whgfW+uH/SGUr4hUlUaNN8NlKYNJPybfw65oZZiYD1aZvR
PfE2y2hNdlCGddzZg9wT/+qCfDIpwb6wnXIFfXSt49hWejJ7eFF8SP1JDyx0/ycG
YIiTRuWE7h2aCOC6ALHWaWxuYyjb7hrawrERO8QjDlmsbFTVw5n7ozwju8rHTSjI
0PGYXtzp7/4PST+/NHXFQYJzi38aWr3qLJ0Y459WzzX64dBcAf5CfrXFcEvmMjrD
32AHg5fo0/wdT1ozprrUTH200dnzRuf4sBb4py+1Oa7BXKihvKU94xIwGEwjUU0W
Kb38Kw6s+wmRVeIxYJhZIsG7RPJqsIy4WV4Wmwc1bKLpvXUHn0Fj8gfZt4tf7l9P
mvCcWLvwng1sH6+NEGDrkpDVweBv/9fccqZJA7JxN7PcR7BNhKPQZ/qZFJd9KxPb
CmHuhCEckvoSlCwMLHD5WMn332x7KBuNfU6kCvunU0P62rpLl7oG+nzUQECSygpj
MeunmHtUG2U5qDXpt/Clz/upAxLtbpVr13LMBKqOmHTSLhEFemPxOwyEkisB4a85
enGz0rRnD8BPjZMKSiRBFpTVicc+EX9KqCWF91P2b3N2Rl3UJyXViXhCaKt/R3E4
GgQ/a4JyKzx0wP0c3eGmNCYt1rsCFEdF8j/Qh/ouqzbaS0ZPdbAqIsLpAATtkGV1
SPUuHCSCHLzEkMulyBH0mUBrmJTGxYb0VNaMVZXbaI35qVgl1q7G9isDLZ5BvY1a
nfsibtCQ2zYKmPKdPmwyStVJWuAM0ZUNLW0ShjmzV+ssDsbyu9Yloqh4a4j1CLmg
xPkdpZ9Ikj45qrCx9dVU7exbicMpWTdlt0insPniqql9immRgu7kXliMMHl8scWi
pgzcCQinvWeNchgnAlgjoYr2Yjl3pZjNGfuH9yntcctWNEDqGJxNrMBLIXuWdU4d
mFT8E1NuGTzWgauXEnXr4qTfkvUBSdP6uidbr4r8hIGrSwc2+ej+a2g07pAE/T5l
p08PTZe549w3OywWV15yfKoIMd9uRlAZOI993K91QOz6yxIRfKsGlz54o2EUO/g9
0xttI1mvX7fKHL1lpLepxEOaP+cocOpiTfezfTjX9zRXC5MexRSssEE9bXUimbFg
at2GNUftO4LbG9USDhRyMueg+rgWWjINHBZ3B64Z1KEJSeeN4Iu6JIF9ydOLQpIn
fvqkXLxK/CMcanvSm78XHzl03jdSzbuBCzzD74ehMYd6m8WSj89aZXA5SN8q3s4T
ECZvR1AcWzCwQjmSj2TKt/yAht72TToZKemF6M50uPKrIiBF0nhOQgY4UG7b/CHz
Aeeo4nUOyiNxM+mMZOrs5KA0D2YJYLWeE8DeFFO8Hy1Lv1b+YloaK9BhQoIYLmYR
c0zz/Vx4Niwn1hwfuNrbyxLoOas1JtMz1yTZDp7Qci0Don9IMbpBPoPejVwys+5k
B2lIOUImY+W+YQ4eCpNmyhDQVp1hk4Yav6++jU+XThv7hEuca8dyxXJOVfSQaUlW
3Hl//MMgWfYIbEXq6laYDzE7R/NaRgfMnHnnjUA3Ojl6GzWLfHtHGG4D8Q9aofcc
/PpF1YdDLvGeejE7Od4QoBIwnDSIo4kKlC1D/cGsLH4T7oRz63E9W6JywP0SiwML
DfEMGO2bgE/CbUP9rcm2GkWcy2oQWSTENiZtlw1SYVCp1an0t77Ngxn9pNqHqk7x
QCUm8JjN6NXLgxJuULW8H4invAWtRxhbJI2tnoDmRPFENth066HSFsZ+Opr4bymC
at2dG/mPx3PukUfTf/KSn/USlofNX+bQNx6PgTPHcurN3u0SvY3OBVqnSUl9wkVM
Jv/f3tyTI5FjKSZx2kvh5grOYDTUIoexKIm4+3qWaV/aNg/GhIwkImwL6P5QI55q
cyiJrGitHcln7W2YTMDpz4Vs3nOS+9IN3ZtQpmXX4BPH5ddpIgvxt8P0u3NsVO8z
RskrGzpH644MBU+zQ4uCJ+aWoG3hPegWNAqdmFbMVQW/2VaIa97uw7KcP+EtPDqk
Q4OnLtnXtKKItrc2oA/5l2Ho8dNdB7p2G28KGLjlFdTTIu5aknXjvnuZLObxZtZe
NkczNnoYhOznttIJwzQQ6mZSjqt52JwBr9lbXDpGNWKaJ+jwGaGRKanacrBvPgT3
CPiNt4+dYXs+B/r8938aoNrGRZsNiabunZuD+DWqbIxMDvu2unNwU4eBKHUacZUR
wAFr475iRBOYP9UaUBoIJBULfdv/rkRdFwLJSnb1vLN+3iY/uDSEUVKN6mdWX+IP
WeE5U3bWWtwv/1Q7+EnVnB3jFbLzpyk0V1BfOYC8W80jzyzJhTZMSCU3f6hD46CX
1aWsoMDuykR8OyYXLS58W4wUfsPNqMV1sxiHWuJso2WLUm7FlcHc/YEZlhNSixtT
dGTDTLP2JMKd6pFnHS/n2COAu54EQ0Ou93ej1GihkUe2g+gVZc5mDmUtC7MaSwq6
VmGkcQK5bIW3Vt91HBpz360yVw/zwvEHqjSWTcDxN9ofiYOlI7weANouN9GJhPNq
xROuTo74B9MTztEUeKo9QVDixD8CkVC6aDd+O1EMgzPJnKH3DvoEqtvRg+ouYgEw
UEJhVvWIrIM4LOBbcEIXZqZewsAQxDK+j+Cv+Q+g7JlkKInI3mXzGfwiwsDm7WQg
QWweDjw4Go2vlVUaGuLZ2qFoNiIuWpgaUgDQNZOz1tA6FtYr+nTWbFMeIak2qexo
g80zyJNM1hwBG1rT/zBDPfrDVD2VLzl2xqfkYPSp9aavDozsV7AR6fi/buNZn5Nn
PLffsnFm2olRCYSQ5idO1uX8cXNTMUNmSdIX+5q/jPy9pQBf2vVxlPCEh8WO8W0D
qQl/RPUD5+fCtsFo0dAS8DRmU1cGt7auzygqqevatziGebVpUqEeElwcCWl9eJms
lPiCpXhZNz+xCHryi19PdiF2YyZhjtEOPeAu4o1dwfmz9vp5Qh4wBa6OVe3z9wOp
yjgiGXFwvjmcOc2f8nAphGmGb9lg0JDXHnTjMwAiAomTPqpn5g+Q3muk3vccM+Ur
g7x15ZUEib8RKKM8UqSbxVVhznbewy4+hIIR+RmTwlh0c3F9gUzmOiae8D+9XLxm
3ph9cL3Wxthdy3GTzUPIwM305gf40KAVOha/KHhlKfwVFQEWbIeQl3fc0v3zvqes
garfrFiCYiX291JN18ZCeME6nzN+1ct2sc9yIpSwlSQF8yekPkNoSeawptfdU3Zt
UIS6suIn17xSUY5mwsFoclZ+9+v6yeZY2zfTrjAdizee9g5wFiFbt3XzWZAns0s2
5qjWvfpaCBa+T6hfvVjBNnvnP2hv/JwIzl6zRK5sJbPe6/lYIfKK/mlr4WhJnreD
Fz/Huu/QH+5kBJw4HN2cdUbqj5q+Ympm9dNBI0EjAeTfK0RL4LloWUD/TFOiPSX6
53CnAzlaHQSsW29eJd6dbily42lGeFBN8aYmTRTSjZQknE6Qe4m3EfhoynneO+Ev
1u5Oh9wjtaqt8QrXGBDj/ytCBfFblOkPFgIoNYl32MYxxujaqN/lnbrW/bRRCeqR
6/MIa61ZWrn9g5OGmIlfY2QyaQkBSp6Jx0OkMcclwmAG6tVLtyuujNPtEjXsF3lM
riGbO+nkomZzAlsNQHYut3EevSfT4r4KM889M5Lyf0AxwwV5LtdfWtr7K+2tXrEK
02slnGLrcxgoN5+u7VrDhuLJuHYfWE1ExQocG0tmntcNV3IqCZ2qxtpL6j46k7Q3
7YR+BHQHUtH/HGAXzdn5iUCVLhCPNi3Tq/klG7UfW9skjDe+9b2I+PQEdRmmMzUo
S7zSuXuUeLyaahrYyuPX9fw0Ujz9vsQWjV+yv6+dXkaDZxyY+gfcRZ0drGs8PzNc
YzLbBGsVI2jJcZe48VRs46kpGSBWcMeuayB47xKw2XxGrlvbphTk2/6XVts3FBXt
Z2A0oZlb/hx0903ag6f366nWAGXzcqaiNenrQ3iMJT0zCYPs4hyctg82rf+uZNUu
pP0cm3qJcWjtplWvkvxn8gIo2pZXN9snrW9HHvgluFItGTJZKUDi6wE8gEsZZewQ
VZlgS8fmpQV5h87pdVJp5Lv+qJX0LeqyJVexH1wQHmyaY3Jvu+M5zqmrSyp33QvI
bm9ybwqnpbWQLlHvPTQhhYmJS5WVbe6ov+DPm7o38L5WYltRLEOVE4KcF/y2mz36
Ddli7w5mgEKxQ9eNSWS+I2yja4pLvEzxp2Mnah03uQaCFrJS35QCein+y8osQlZO
usH88rE90td2SceJhwt2EqgibikF2KUPr/zTA2ECOchCm1DDYGtPqE1KzL0NovYn
NsyMCCa88Jtel5ZHdAj1bNR7XgKe35XcgxHJckMDYnV4eGsdXYVnAz8LB0Q2xknu
DBfbnP04BTprtZgA8DOVIwKmreCEcDgMA+FLlEbXBGk1p73VgcknyiVXKFKPxDi5
QxtVfMzCykRtNOGFD5dwjsfSROqszeumFkovjbSSsch5U1RdMzDacoY1aVJIPUi9
mos0oIHmZ77HtMqP7c7ClPoKAlx2kw7d//jf6K3PzlS62gXPxdZogVx14xZRKRqT
VXEUn4eNnXxJUJh+4eZBuW6+upIzy3zytamVrJJhU4Cn9dIf+Ari4WwDbGtXVcHC
XXJ3yBM3ZNWkjCqclRTuUU4kGyhAYqYBAQZ0XIdo9YdM1Ax17fmMmQQ44WD2aXRN
zliAEW7FRrcGx6AsgHwXk8jC8H18yy4g08In2MGICsh+R78gQxsP7mHZBTw+K3kG
o/ClP1YtwfeEYyGxrqyuOidq5E0K0pPCi47dZ1QJa7kdHYQaHgj5OsfVWQuMMJAf
kKoIb49Pu3QMqN3zQTuUyuBeabQsHYOZGHC6SuaveIhoWweR/qvM6wZy59QhIox7
oUWw0VaXWhGGLXe2Qe0RbhJCPuGei1Y0drVTopBoIAQyqTpweYBtaXBpaKOwts6z
d3GnSWom9E8CZr1xfF4gKt1UfFnby0L4sbGxcl/5AAXWHDfghhsMBgGuJHf3RBp3
DXS0EWM+vcVh2TtESPrGz2feS8yxgcNVqGbR3TeRySCna9wgOoKV9JIxPmtnFGVJ
C96wbJ0YrxITShjfmGuKpvTEORGctU/KD1DeGZhqfssm4ijGVc4vO35T6dMVXesh
/LCJZbQ3BGf8ZeRIKjs7KLtRz7EC9BBtTYG3kdCx10NIga0dp71nDn3bCZgUo/MT
YtOdMALNc5nENNo0b3fkEDanSNcvP4Vi/IpGVnMSfvsjv8FzhDlNmjkyteVTdEoH
dlxteLm+W+4EYGkP8vgWaTHIYX0KHQGQ5OtueVS7E83zsEu2+/eNACTe2JIt1MjH
hGB+gSKEod4xScYMHDvNTNSI3Q18D7ZWuTQE+VvdLuQF2eDSLk1qKQtSMzVIOBaQ
Da6F/oA+zwp21Qr6A/aUCzeaehO75HG1D2KB38PLt//i7n+IPeCRveeREpBjRzEA
OrZ3CsGx7CDmWjn5mqKrfZZwPUjv/vvwgGUlosDT4RpSf/Y3ZcJXI0zh033Zg5pz
v4r0r1nz3Gw6Yq3keXVre8ugwI4ogIvicQOXwxe2UIttSrEAUboUD7MOnX4UW8lO
e6BqSScevtb1THRT0F5i14HhITna07xiT12Xnch7mXbSoY/sjd5ykU5kwr2/JJvE
d9883RNp97Dn1daezBDrWTO9CVdwRsX7tfILk49ja2ee2FQrMdxWVdNnxAX3y71T
qTM23Xt3nng6sOYEH91JM3KEf7nbuyqa/TZQtljFAko7ik2vplKd79DrA/UOdxPC
YEf4ISrdOgyssfYRtIGtFqKBW9a8Ih5syL5GOYDYngprs2VMi7gYYhSOsESLDI7g
DKmqpiT+o4A+7/5G8eO0HPicTazbcZjaPV8BQHGJmCv6bDBkXGbqnSO9oIJ/S2Ax
Ehe6DIsjfUymPno2N58/8YaiVYWHJc4+eHwPfbLprMvlYtrhsXSsJ9dyG27OOgU2
F33MPeIE2hk7q0cARAIEUKtW6HTLbChxWBAszzLDxGnR7mvtdv8ZjwcBM2QAJEpq
/AHxDywRw+KA48CdjrWeN1bqEjbgMT44U8Z659taz/CKSoybkZSYpB5VAqbpwc1n
Lhch5c/nj0Wtu1kJUz0H8jx7zJZ0wOakMgl0yUm8gUCv9YEslK1c9UcWUICuU7lR
OkspTxo2E9XL5XDD/sR/mvEhN86mVidacOweCtoFmEHLRsxF4vnkbknL0FxVS0pl
ryk4WWJYpj8bq0U6n/U8AUScZL+yE7AyAnan8ZJtej5lyim5iFOcBXW6AQ8qLeV6
8j9eUKNbsOE9+iYx50vS1hhabfYGCCHZLV/G8IssfQwoR4SVcsaRw1zsDCrKRfue
2lE2IYiHffIuCbH8ABgYzrsZOaMzdF8mJSeicw+1OU++QcQQX7QOmF+Uz46CmyK1
HUX/IKXI0ZZyP8u3WnTbgGKm1ctREcv1MKHSfwpFh68IQp2/2afr/jxQYalqgcs+
5CVF9ef0OBic+VRP93/6va81aAoKNKjbqmz/AuDvaD5laU0crrdlnguTKPHf1N4N
QSonVP02Bj+VnW+MH0jw1aO/6UonZ2kxLzwbNazY5OnARTK9D5ITNojC9eRGzfxM
zb0NGIvHm85L7X2Nq6auu0EavnZvRGOnjoezceIKoY9eemdy3PtPh0LWl7SlS57R
SXXbvjxbxKZHVMSG86KDdxncUBJJL1QvsLatMklMO3ZYEk00L2baQKw4fnP5OuJK
p7hdz3Mt1DUECQBqbg/enEt5pmtYwpILv58auJNfPN7U9emsbYBauizbc1jKi4Az
/+Z5RGVrA4PS8+KX3UYVThd1WbjcRQEFac3G048Yo2O96XjKgjnt93J47cQL58bB
m0QqtVwyVTkEsVzoZQloBfMEwq8qAkshFSFd+H8eoDELeiFkcyr3k/ru6KD0rvkP
vpG4L/kbsXEjclYpxhXgEEeXbIZG4aITj5LS/eL5L9556dXke/FzfxcCzywCmMej
avsbkvoOXvAZLbaFNSIJgOroqq1wc5QEFC5d6VuRix1C8EHbX8f+46TWT6qk8uq+
cDrBFBPan9tbcy1RyU58fVhlCqLT/+xPewJao6Cwts6731GXvBs3JGw96Cacn9Y3
Nzjy48hYEA9uDGxOMxYZJnKazjbTI1P5WS4HTs9rof85MGVLLz9zTkNn27aM4cV6
JNikbWZ2GGOxxggqVZTuY01NdVAIrObA0NCEfxyq95kfjg0tBDRW7fOA4Yo8tXF9
PzqNSOP6aiVoOEtVqKV19L52n5bn0CRUrMk4VyZ6cStIboHb65v1lMq2YnoCHtkA
+b6zDj8amX8TQnF6/DjDggtAppOKXkZ31z2MbJeHJatSWmWG8B3/dEq1va70na8A
O8G9RTBmJFKlrSBWN+uj8I2XorglQ9gnKInNpSpW0id3sgNzbQ3ejauwDhEU1Oza
nK62rEcg33BN6tCMn994bfHoEutt9qfx7Q+0Tm5tqw/w8pGD5YUwUBHU4npCMODW
55UrPmB07WsVYshR+zupXZgu84zdXU/svj2rhZORJzFWX8fd88K1N0Uq+YChLYw/
P2+GLxCa/vei1ivlR/ZFL6FJqLI3j20IDNBPxpkLTpisAHVNDfK2u3/OYYROA4Ht
41DiNjnTdYlzM3rf+IWFUF3wOWaL08zCTL184gX4GkGW1t2PQj8MUKTaqaQ7e9PL
G0EfL0rxrebk8ZrcZ74sAp6HEyezhgqRIjVOY+vAug0nYVmLFJi0oVfhVEb10NNy
Dyttw/Pm6ak0bPBA09VjEo0lCV+fSnHJoaCP6C2fTRSV4zE75sp+Umj4/Jv7bH6x
HKCxGIGyr102Y5TFbDj9bFsC/x0/FEd7g5omFVh6voqsxc88t5o9tgsgT+K9jnC7
3A/Z+m2h2BflNtrEopYCQdy37DIamPgmYBXEgek9AJaj1nCOcHokW7zkE/Ece9Eq
WXbc8e2xdj/cSjDcOshVkMtnWz/2fn23td59kSVWUvnNT+wineU4HXrDmp7ue/SM
joYFOk8v5hnpvD5xcOUPXieo/iE1oTh9va3N+w2XQ9exoxZyhiNPw5JB4fGvW3mN
ljelUpk4dcjIH42XYXS1ZiDHklQj8TN5R9GKcQuEuBwC4F5/APXaLu0lnOjATKxF
4oG3t3PykIdcbYPTD4fqCni2cxO30Og6ZHygLYPR6MeTtPVAWHBNpzSacLty8PFS
4s0+2dpKqLb8/Li5oRoaRrfheWLp916ZZy05pG5Nc9X+tfjKVIv+0M1jmzsIn6bt
3PTxwEkVmheILQl5DSbciomM1gc1o/3jS7hYMTWH5GYGpCMC4v/1moxIQx55twYe
D3cS9bqcVwTg9oNi4kY1rf6gvksjtNLtbzchNeOM8DgE1fSR4FR46fD35OB669qN
254OkYF44lWpoRFYNgLeTmA2VKR7DroxgOptK2YC1WQ9C6WSnZt2/kAcquiKIo/h
/KavTqgg8OAjOzVAbOAm7nKJ768eauzbnVcBI5tCmipBiRuXUDB6Nh0F+u+3OdfF
nbVgq981u2D/mZmgqWKOehEn0oV5ja9Y3WEzkyu1/yNzXMk40+lFVYYsMTFvcDnE
s7ewtYBlHS4AgJvYIjsjsN95n7NMF+9kwo7JoNnNcujq1MP+DDCcKemMFNDL56nK
UI5F1QJGocPi5xRSp8KrT5d9i+WCoZZ9DwsL65YczUQEgsO4q9o93mJpDdv2MzJN
DY5y3c00tIKLw49XV8n8VW0eIKe1C33BL2udH6U//DofGD2/kgLjxJHCsaJiTR/b
H3Lkk6ooerHOiDev9S/+j9IcZEL2U15tzFTX0KxAhzgkQiBmQrCD5VlFaff7uXe1
m1LmH+4+MA6RCGN81GOYaen/RU0QgFfKbzy9d/cpJwNFgC7W0LMAibVTR1EPTsjr
bxLQg3oHzl8YFSSxxHOvE8zsqNsndLMI9FWLqcZ7ee9mbS3IbohJwvAxuqf608VV
iAL6c9VF1pNNqI2k/b3CozeC0upoRpGpHApOKm2rNc/eh5oPxTK4e4L9YfQ56VI0
6idUob/uk7E2N2M0P80ltFdBiLHnHnzw9fbz7SlFnTKJnj38b5AqCs92RHyXztlK
ZxOvXRxZNV5YdT1AeXWR26TXOZWYrm50SwBvvZma5WLRr6J6Y9kxpMR6rODtaABX
Wn4Mps45DCyBtl7jRSRAmD9ZvyjbVQpI3OGn6mr3mtbZ62isGWNgxjT9LmVTB7mj
Gn4oH8WDx0KnWsEBoyPB7NgAwiYmkRSq5p+8MCpR826OhSIViOzBqgCX7Mda3saA
YzLVA2AMuwrQwId6gkmEsXtPBGFAMrPfYrKxPghMLBbYOsq5gEaggywnRrLMI6Uy
LY1tbUuSNlG35n5MN8S/408z+wHR1+59K5TUEWVUhMUtvukbCbj9Lk7f3mLVO1b2
t67w3UaUam4JngdXpAvVGGl2A74pV2kLzZZhFLXSlgSa7mi5jR3SJPElRTvZoXQA
mKvy+UfqRVkmT8ASOAl+0A6BuA2Frnwz/mtd8DQMe9/xDmaiwu/qYYgT+F3UUhC8
TFF6uPIagv5lvX45kWCXy14Ul1rfL2WjYmdQ1bgd7J9mvcPcf71xYSnqjFy19mga
d39RAKceutO8MVXUlJ+fqO/EX0eQ21dKvUEW3Gnd0pNGAnIokIVX7KQHPU3bnoEm
o8zuiWjJmzsFUgktrK6phJBzX3u00s/DCuOnz68+dJSECe5w6SHoRQ2Hj7PsyI5h
L+MZMUaAIZtXeuFctTVEmk6LUr64HXR7fPw3NerR3SVtOpD4M1Va5c7EMlxocbM/
rxYaB18QW55E9Cr1j8SisxFb2C/aXV+csTp0mSSYbdjCqXrX3m7t36rZMMxQK4oj
3Db0oWtuBqnmSZMrO5sP6S7jVVI0ixZqfT3/pLOKmymKlYfH38bP/xSIM1T53ArZ
F05DD6mrUOqR5/kNcQent0un/XMK9evWVrsgwMiLBoVeH2e5Zom9F88KKa05ZBSo
TUcSUjd4LOmh1LopuXMYlzVkOaZOxC2jYg4NjhqF+TloVozuFOF0byprxjwLimjS
oZrxxd5izheegoND4CtwTtCqFhNQWIWmSCPQVQo0xEgZVymmfeC/nvLdmpWshRyK
5wUit6522RKS6F4wf7TOgbTwlNaHhlfjdfi4VouJ2FRNsF3JzvYKBGxH/qyIXgh0
aUgppZajFc4b/8oYNdQpJCRM2AFs/1Oe8zn9S1W340fkMWbSNYro+95aOUZG5WzX
vkC7bHzd6F6eTzL5rE+XMssVG+eDsxfU4ja+Benn3P87ytXmpdzYx8k3R1V13KO+
AcC0xiqZfzYuiAHYULO4cSepXnyVtHNvfpOiq8xzTPEuUo4HgHTnEfQPXJvhVa4f
LolZtz4IIvebKIkFp+b7GqKfuRyB+RSm4V3CimNeSrYmRxo+Daln/11m1y57Ya8A
KHQ92EDGPPy2YIwt7TuEAY5H3JpRo6dV+6QIdAW4TtBRqXYfIQXJq/UxyeFbbqlA
yd2j9yX8Pz/5pfppq9usMNyANnDeem9A6QSaxc2ZymhxIt2p8Loyef95U4WFbQmZ
JDALwcnabXF8nM8QjDrIMpavGuO03lR3QDn4tc/GF48b3iJuPGgvt4cq5AE0ckaM
71AEVCMu9Z4eFt57CYtUYFG+tiUiU8NOd3KkwUj6Dp1ch7MswWauYIsOrJS3eWHX
Rtrai02mhxWOiKIRl4DJ8uYqi1FN13qQLFM6LwLf3rxelwc7mlaz1CYkYyQfoQZP
9EcUM03GP3Rvm9wgwGY54LiL/jP2sTsVSmGPYsFDjHygf+DaeanESNifba8iQyNn
vypoiWmotzuPCEkaQIYcV6w2MT0jkLpHCZMrtM57NAUqIaloJTviRg1HkfFcPsn0
oYUalGPQ45xYRlcvYX7nCENzhY+yzG5JtIBiStm6M3+4qyE/1qMKdy7GcFFLtymG
2g1WuQlwNjCZ7v1y46u6Rim52EcfEbP4MdoFbbx+r65zZAYW2SiuEz5EkNcZr4/5
kfFU77cv+KEtZCEzF1j5BHh6lRN/wutpEtkPF+35GO66FFpFavqbhuz2C7Q7qqpm
DLk2/UMaaQnjUonJ8u6JVyXsk6VvPaK3FfqaLuRMrt6R9VAGqnelDNiMssHhSSKm
OcCwu9k5STS+8XJlT9VZT242rGmOPfLVvJb8HJm4+XP9nTzbJspJa1ehd2Ii8NzB
0bPRD9rdDlFHfnR2GKDCNhQeKbEk22I0tVqANggAKxrRHrLHgW4se/TZZH9sYopK
io/bxgKlxuPEzqZxDVNyVLlYsrTr1m6hyV8aSHsw3sxk9dqkW6NjTYcMuTYuav6U
o/CB44VjTDKtot3uxy5UBZg9Ig1gSaN3K6qp8bKO9e6N8qlj83AcCbFFkKHz391O
t+yVTnodKuFs10f8TwnOpZY9nkAdOUKrOxHQzzW99GIs3kmHb6pkTAX13rVexY6X
cZhpPVeCJAoxN5SYVPG5Parur6Rg4IGPhhedgegcxlPSTRY8jhsbpjyMpRlMOrf4
sicGD0I/S2O8gzW/+L1wGYwzo38nnjegt7+qM+9pwYbEmdMz66r+YnSS/R53yzqZ
ArB9njI4dc+7g8D4aJYgubiON5E67YtVNH1Ze0LlL/SdAQQ8+FINKS5r6yh92lNB
G5LDfkHXNjlITQFWqyfJvHWvCnvQKDIW2S+xq/kuAKQ5/GgubCFvqd1Q3xSYmBfi
J42yohcMNOCEJSub94C6ucN1LDZMB9u078M9ubJRl8rSs6R8il8QsZLUfmjj/yTC
5P6BSPdSRF+jKXctXKo5Kxd1UTGY+C4s4DBbXsSceeubsiRF0qEaHaar+rww0h3l
WVMBb0b1VVvaxszRx2ZIN7o1vQ2Js2KsgwXfdTLHrJxRUbtF0/Qithr08b9HUBNm
2GUfMNtvmQxsXoq8rStdVnMMne9eeBrrTVFVE4gMZ0GoKIGpNrxH6fr6jjFU628y
LFU3oo6vr+qECler16r0RtCT9aYl4HMuUYgjg5QwF2sYvsCM2ASVoD3HheLATZhh
5atkEz2oIKKezqmjNzwt/nqnRhPmDbcERuKhGavuWbpWFlau4gg2tKe9o3fLGN6O
jljThwiGajNBo1nPu3cFbIVwdblSckh7FxKL6oiZ2eUYTkhabja9mVRdODbkUBsA
+T77VDQcWAoRhMyKYucx+BNLs0klODPRYkKfzlMvbmDB444Ey/sNBAwKWFZTZt/W
bSKaytI1R2fRf8gRtphH47qE2PyDYP7TxocQ9VKCb9AJut3G3APVTYeS3XvFg4Go
CuC/mOSQMym8rqjUbyyy0vEHdJJqMSzwS61pi6ccMXmQLdeoeKuINhtn30mNfFi3
KylPQ789m8jBqzgAMrWw6uAok/+KhVRc7WxET5BW4BUjDgwpmXCtstEUAQ6hpeqC
FsQ2UoUmsHRo3TlE/rL1K1OK4VhASZIKVnsSfWQD6D+E0q5jxncd9swhGUB9aA4k
LJBgUK7bjqBDz+fggMXAcIOuDZPJf8Ozi5umUMQ+OhG+SCXbbAwwKdFX/23tqnq1
aWyIa55bMZ8AKGdTXp2WDobpErqlOapMCcmN4evx8LlhHaNpQSCN8ueThXBUEuqG
sNuxEmuRQcuzsS6JKlUlz2Xhi0MJfvtzshi/i+XpVEbY1RGET4ZAC0IwMMsYuWr9
fbJ1YU+jOlGhvbCKv+n9KjZPVbBmrskxuC4/CnmsrdWHGfSrk98qmP6TBucDNeY+
x3CzNYsMzdJ/9ma7XjMswNhmEw+JRSLmVuea8eX4+atfAAJPFp/myBiy3xA26ciO
N3Qnq5GqZ1nyNc0RIjRKUy4c2sHC/3j+gM5B8J+RqIW5ENjGvN6Qas0ryLuJXJek
6DwPTKOmSAl6PIxG8Vyzviz6+BJtJx7Pdj6sk8eInMpOdTjTtEgq0KxORH1qbJ3g
ePLu49unS5j7XZm4oy/BUxWFMKqPla/Z/q4+fIehszpwStTd5je2rWS9Yp6e6DAe
XSBX7cbjzWwaESDF//mpMaqN/rdf2yTyghtTBvNTaUa2GtZbv7c5YBGBiLBvQSb3
z/Dkjh1/Q/+nm7UWa/6MCQ888gWzS8fJo+eX4umaLBFdjTLaqzIAo6jSHlZm4dCF
AimvoiSBdT40CBiZOWAEM79Ts5RNMEIZapsmlKRdTKse02ZG75sKAwF7N2V8wJCq
O0vsEqO2IgTw0idLLpar+y32n8leQI+EmcxHuY0OSlpEQC1J5EIT1kvpi243K0S0
J6sC7ZmMiLSnMtdBFZX0NJYNtqqzpDYHXYkDMwImxsZtIorJPZuio3m7Wup3qaxF
r47fn+u9/BGPrYbNW3eAvTWtaGXZwP8dIGLDy8L5Mo7u+cNrEqZE4rtzrRaen5KM
JunW1tP+hcIbMDXz6XRW25zP2XmCmuF1xShU3mS5wtUE5MDEZFuF6fay+K2cCQP2
Lnsy7/ZUOs33TAGOw/n8ukAzJUtB1qs1FEAm5SFD/OFQJLyHUeB1oJsQ+8mbHA+d
DGwitTQzh6N/SuVaBL4/V63hDPkHuIZh1bOe0Fj4d+OOUS/iS7Z6Kx6IhnZem6L2
coZy2sfHQnfB6GluYVT52PIcMzBGEanFsO/zmpAc3OiqWVxxifo2DYnkkOQwDjDY
GOMIp+pTY+eZ1W6iCvxWvaXqsx5LHuZLYpeK/CcjbAmcMWM7NxROJyMU7f5RRKfb
W0B/83+yQn+iJDFqSpXZezxoyJ1ugIaRdwmedinuizTLfVB61CpsSv6qdPB63RPY
bJ1nSzD6mn9Ijy8Myyu7xKx4v0Xkk7JjSxh+iFDkMhEPBcI0tJ4RngbmaBRtATGR
6P8St5aS5D+bHCbCSJugUSWzfU9xJ4IKLYF2D+7Dw7m0RIAfzQfCE+rhTWKhTAtM
6P2kT7hx8Qrzi9/9YfMumU/wKoWPvNI7iB4//tL+ZXOvPBpobD5im2w2Xxyk5n4I
y+5us8Mfx/W9zAz9rZyq92xdeM2P8STBpT4u3wCm2o+j4JtjV3wudWjbI9VsYLXl
UdGTFRFIqCpNO/Hea8qzc+kpGJ5i0Bx2DxBHq2D4+lzG9s+pFiPTR2+5naau2tYq
KsmLk6CuWsfkRceqFWmoTCEmGNezfjPLVjGIOxEFkdDIiiY7fWfVYhkSP/p3UWVO
FmcEvhflnyB/QLTpMhfD+EH+mbVLd+FRsydjrubNrhnY6bqCY9iHUCTWCPoUAvby
gT6Yr+c4cnXaHiXLtOofkmQhoJ8lgUrL8PJYWx5yS23Qh/T5UsGh/4QS6vYuKkFQ
X+4xJ8eu66puxDd1MNqO/D8wNSGnAVstBQyTXjzGXgnbxiidre0uikDX5u4oFaDG
UsOuVF0D0Iv4P514pRLTl99cctwJMOpRKdm+EhyiqWAVTemCjMi7uW2/AwUe9B1S
IVnmypArekNUffas/MZRsTmuO/9igmu50B5kFZZsy7bNhRdMW9v7zHtzNv1v25t7
4R45pUOE9HEhLPuft7prGYpPWwZ7nGN+REi/Q9LA6z5mSawjaw4Jo/tL52Up3G5m
GSjqd7P8g37Jv89TXWWWmQVOsTsd/mhGI0i8M2RW6KL7TWXzRTUlCBUrdZZHlM6u
UnjsFKkb9iByc1lxVOuQiy884k2eVjN/+xHcjvyZU3YHWpDGemvcrwVsySDfx9aK
OIohG7Mgb84x+2sIfebrYGPrUkBBGQWHvkACXC91i+/+MoYxrqldyfER9dQCow47
4A8QuxonVb6XnsUDB3Dm9c1IQHJRTKsMAb2vL20iGCqr6uLq+JRqDl5fTjTqmrLp
9XmetnS9GKCkntvvAdy3dNf17RGI8WVM2uWWNwEutbvhj8h/tSDSmKp6ny7dSJDG
tzPtVkm5eJNa43+mQIVkhiJ8JdHmXNJ1bX7jjjzojzGSy/JXvx6sp+eazCMlfN4V
TMYXVBBdSrsitXDYPiycKZ2G8RkuHLKv+sWzdFr0YS0vep2Ru+Jl1BbIKQXhuvzj
RkEGLeZYCFd4m3CtYBmbXdauOf1O8V2PlNzJj15EDEUtP2hRURjy1I3kOYPsMfrD
nFV6Cz57jKV0MVJCWxonUfK56RpwDFXPviW2r+yd2sreIqurf12FKXrWrRq6cZOc
Tdr9JakqAAAO4SLjgFFtufWEZZgPquPuHxBH4ElA/vUNNi6f9QtCXFUC+km+pDrM
ofYOW+bXQu8q2jt8pinkBA/+WSjZIBoHCNGGAi40fLQKllOP4ilXK/zkLrz+sO/8
KfhCAtpqJ+YOaVURvzNdcpO9KZuusDR7xm6Bu2X68NbICY+se9n39AdmXAfp2aEk
NelAKpbbeNHR8awYYViqFxB91wv/W0c1QDSQi0C/wrarh6NOhprjPX1mIFkFnjIA
6j5h1yoEMfjZcBaOtQUnK/24tDvOMM40iacdXjWFiVozVUfgJKUPXK2cgdGplT4w
QeMwV17+vewTWyVP1qCulb+VJRbnvxkv5qIZaPBZpz8O/9PcxvgHWTvXeT8nlXEA
Lp3G8a4kra3bsOycvRO1IDB8abTGTasAP8QX/Lu3P8Q+kU0hnb1n6WJn93MRxHNS
d+tr0+3xAjWFUJ/YXJHC2o8UaHrkKAo9b4KNdw2YqRVW8hRx16wTRVTmeGckJOCe
v6bZTa4TuM6zh5VJ8I1i3J4d9MlaxFFTCa5WT7w+RaCzUiISIsOPD4BTQ7rO/XXa
GFDg72+NICzgVFHG6tChfhq7vlxeG5IX5wRNi5we4tNHF7j8T/d30JI1AoEILP8a
AbFvuS+lxBuAmqcJLEQ/lskQGa3wPqcXfVZ/gfrSEbHs9vJA5jGC7gGuR0XG8YPh
Ah1wiUQ+oSK82hIuHdoXM908PC9iiU6SArgYcR7/jB262nH7uxr+RjNCZPO5nxFi
JU6KIE6Pvn1+DuLC5Vltd0MzEqvCVFLVK7KZyRraneOpEmDzxCjCOI6patDxbb3K
TjoAcdPewI2w4J4EBPguGunGGUImYngihCACyzKS2OiumL68SkDlFe4OZJU+CEP5
bdd6alvXZyUkTgKJhGma4YlDBf5398YGIHULCebvKvnecfL2lcINpR4HES4y9kv0
9r+Rv+L0Uc5k7l1FfmQXepSYoD6za4yfMYYwo6QuIXDJfn6hwg2cjEm2PqlYBLBJ
wv3ZeRDqvvhFONzkYS+E5hCP7dklnK3aZphSv7AeKF65mpbj4/jsLH3EajbxnKkh
FSbdbRFUadi7OrzEUrNFIN0E2x63tk2e0Gc3cy2XckYLfyFhdM0u3oNOJLfuT2Qu
vq9A3HiRl+ueZ/ahP49nYQgK5vZ2fBBFLxbCK459WbTUTRrULpF9tjx7wJCtk92a
ZkvW2VtlWl9j6YCDdzQn8MD5ldXipGyu7MD8UDto0/YpN+B8G7/GPP2wrF9nhPBc
jB8chGwWawF8DMwZg690Ik4CvArj1/ybW14LUZplzPAE53p5Ju6s/xomMlaf4a/J
WZtdqly59CboDfo9ELBfIKbv7perqvXDLIKnx9cpKoLXR+J355iwGoh+tHZBzU2n
fTrlCluwwWOzhm7fbDj7R0TQKE7I1YaDIGMmAKIXiDIahPGyurvzzDmH+wv3kjKv
K45BKCG5OE9HCRc49WcRkZ2np+gVhtpEnp1vuUsuvpcDZF5U2MdyIf1HIo+jElSK
s7Ptt8R4o5fScgIMl0VaebFIt7IT0OYGXa+aYEG8B1ECSyA5rs4iq2Sx85pIolE+
YuvXKQja7N1cjndXWUSraqDhzbsgdyz+djCxGthyO5MNexDVcCHhZbHISq8AQvrf
bq0TNzqPZhjYJq4oCNMW+EB7f3Cg66PsGQ489o1FQXmDK7EQkoKD68rZw+ktXmQc
zITWdEuMbj80df19tylXM2iKA+n3UkMC3BxNhND+Dopbrcon0Z+MGwpqS0cwaCud
YObnNGIfb0DE8XVsgXqrg8nRW0zZHEYrRPepMiQPoqx+IfOhxDIWXRBXRLcwqWh9
aZxgYC+hoXwfq7oGXPaccg30n5rprRVVglVkzLdva+OA0EX15hsrMHme5GZPWo5N
udkmsIL+RxYpJplMjGh1zktphR9ITggbrw2V4g8JsSrKgEQsl5HqQ0STd68KePzJ
wHujIug2RIerCi2oHOkrFjsgMDBrzXz6pxZQFRMa9K2b3wwynr4p+ozoq3cfLBuC
ZLsTJHPO0+SHKQKPY+UjI1jyMDBtHgahfwvt3vVNnOKJU0/0TriuRXYKc0JDtIut
xvuB8uDELSK2SUsN+vrf7r3axYanSgIpL61z8yv3JJeMLqmOj03mjzK69EJNXXvc
YpYk6HA86ZvbkioDeqz0n6sjilFyTKPdyhkhcAFpdiWH+sXji4T5+kLEmX0I2CVS
wIwITytYOpRj4VwFrAPHIuDLOMvstZP+uMiYFvhIWvfdXd4pzKPFRXQdREinIrup
Gryn6x4T9KY6sadPFFyPVgX79HOyBdDVQWhHuJniPQFOIvEB5QIN4MxyofXkaY5p
l0GqHN0y457xKXyW04TZVdiRXYzuddslrERsbsl9fsvxuA1ZK73JYJjB4tDUthaX
G1NO/LqgpR91G2OW00z3RhV29R5E4KVioz2ItPUFEyb8zkAg5VcpySRb9p+b9aX0
F10xQwqlzuf/brmu3+zUqJzcjPVpw6Eztq6+ZY3isUSMWBGeBI3C3npTRivecHHC
WCR1FVLluvFxGzcHn2m2K0Qd+6XD/OIyz8XV69uRtoxPAhvTEPa1Tdw7c2i/MYpr
z2jrKOtIafPpd2sa93O7oIAzKdmwxo5d0MYfHpOj8A95/beRm8lezjF4wLnXaJ33
Y++qDjjroeWgVLp5Dwr2eRXl3X7Q+ySb3uziO7f6zsYCmvVxgvt2ATA5mikQHBJr
gO9qkDoBjKUvlV6ER8X1gsPuoxMpmi8BFu8wQSSKY/zWJ8K8E+cFPbFwoo+09sQe
EqbFV+zyYmM7PYmpTbIByzyPHaZ6ogkCQLvHOkUwWHfawe5TgsBhOuik0MyQrV4O
VVKGbhFIY/2D2v1fZYEjzauXsgNsV9cbrnVoSyRxx0EaCnF9bfL/pwYdEMewyZhb
TZ3CfEXOHW6HEG+8yC6qmFfaZKv+vvY7q++jcBphm/7vjd7zdl+F5+NREquSpapv
qGPdnroWBAxLz5S5EmiTta5sqndBYXD0U8L/8jWXXCHQKi40nG+KhEMUHSqbvedc
UhESqO5szzxM6W6qU4yPpqfwbjnMTNG4vHnpfx1rcIpBFitHr5EjtgAWoChsN0mr
QXQqsDMIZMugl/vyRYpoxeixP5gYR9qOGzx1YfQC5G6B8P5h+Opnkk+E3cwlu4lU
UV7fyUSNcLIgTCJQVzbrUkkbp1rwxhAjSXKPl2fmHatQQ3GsbKqlkgdmLrlS5Pt0
DJ7+MFSQl6JEu2jfCuF6pz/1tDa+XnfN/yT3BXIgCED19gGxzEpUss/iWrMOhrZ6
IO+rZI6I3mF/8tS49z1Iff5TVHbiOGcPfDXdVAhnE9S7j30Q5pmzNfos22R/7p24
Fxb0usCQp6laws/1eETV60cIpFoPaCfTzEMaJ6LpZAM0Qgt8gjWepHTe1J732xjB
wYVbkAfa/coEtTd6bI808d2a718HbgDM3GeVNZwu8UAnZ/m8TGs9Wez7eEtIBHKD
E5xD0UZvM6uXTl2kq3f8Zr/tX/mLdjZYz0g683bsmS9lblVw5TOljtboWCFxDLug
95A1cXM78yM6LNsjC4jIVbBWXP33YUYy2YoQlxC8hgobjtmJIyVI4BxCnYVNK0Al
2Jl24ly9ISfRF1tLcGMQcQU+dTsi+X2OwBEVXrmNh6n3EsjWI4/daqT30x4nh+3/
RZLUA3OUHcOx/V6CjUorYqr8FW8hSEUueFEw6x3jLj/tbCEDiNWOUMONbbjLNamC
rNv9hHemOjsD45QE2KF5yYMnIY/zVYnVQ1lGdrk2qZrjiikM2EYDnnxfuQ0EkplL
tVV80FIKnIsD0EvxTqecHRK5/XjDAyBMUED0BSpts4saM/kdGg5BbNFOgtYN3VFj
Km/P0o8xFznoSdBAGAVQpiaBLm9F25/90Wu8vPLPSU4kuA7sy9K8QYMBmm8aj2hG
tAeD7GqJc1WboL2UvQDZEIMd2YCJO+4sW1+zdLn3Xnp+eYaMHEkfeeqxfMjjUyOt
zMgKXZ1nXdNQS/09p0E2z1Dbi8kzF9YXerrCjhdBfDwpI62QP/IxI/Exqp7+2T6P
j+/3WqPpCitS8VSzCg0Helm+xvwKn8eW+FaKhrfnLPMMEL4+W0S8lN9Jnk/GmZ3t
g0mX64T9g09xdI9X3q/KMPvXAPmYLhnfK0tMJlq//v6ZkOqb6NdWSle7yKLFsk6i
LfNOFK5aOnvKDLKjYn6nOLUY+fDEjABzpVrvA9l1UuGA1odg4Mka8KXPvG4uJtzN
lmMY1QBkvU2Ol2zY3TQ0WyNAiW6H42gATliC2jGt7Fo/SuKjVkhjG/ykWPmlDCQg
1p/0adbpC2zRRKmgWNG2o2065g9UiXbvTercrAZAhImUeP18A4A+vVZZk8TfRYzS
A6vQr2egDnplSpvnxhB4TytbsTVA+WKX8K65qIu3L3ZnofwPFLVddi/FFA+u6O5n
f7Srb3qj5kWerxan5YM+/37aPruR+PVxnwp5IbDggIunBlq1IaPL9bE81+fc5FRz
NSVXrOPVQV31+GUW1Q85QvSFkz28zNdgNJKhqSdk1jt0yYxf9cuIfyBpeKp8rkvv
ZR7xkJEIXzq8StPyjeT8FC3xplvLQaOjZx3/wa628HC0VHq5/AAUVLB0J6m491it
uUd2ybMeEagW/kue/yC6zFcrXh3IIINvuCLL70P2yYsR2Weu1CcRtFSQh7xPggtT
XxglCwnDhFXiC3ijVrOcYjIf74hPIZhUJoLuCQJPEELwK8VeVLr6ja5j1Mumry2m
MbKYlDsucnpqjQIbX20CaMjtAE9Cq5VrvSC3W02Un8r5GNuCjq/Ol7HZ0IMf9VdK
jPd0iKwcvNOMwb3e7O9Ao0oSy38d/lVrTfNcLuUcBIhIpp1WLJwxjld53dnRMjag
hEy3nuE/M54a3E1psst6oUWcxk40p86c+arLaiNV2RnDpC0UIr1UsYbh99xRo27G
qogLGDypKFof77BY3W7PGqsrK1k9pzlOgk+S5j+w8RrKn9gDPZJo2Ibx80sGfYXz
h8NgixSD5Z7AcsJsol9xRDD/jh8W60a/pSu3ZNJr3ANfWsfdW30kOM34SC7jVeM2
FT3dG4SkmlHfGJol5iUIBFbSrCD2Kt2DsxZ5c85xgZX5AQmFPEM9Yuum9xl+z2Sy
wvkHobIjwghcnWviYYzY7Z7hgqguluycSdf5IVoiR2cYD8xE/MU/rNx+7zi+zIcC
kvJ7oPfi6uikYy3q2i3tChtT9EwvvX12u5cMTMkPVMcU+7+9BpyUeWd66nLI2eId
iVbzfTHkzXsCsAVE+HIZ6gmd76beDJRxkVV4raAcbHEPJvRn1poFKDxP/j8rn11a
NO4DR6A6Pz1OlfmTaZ4sO3O+YkCLIzUKIe2yUVMiES/WusM/n7sLFfOSc1XFcn+m
ggRCYqaRLjSfx90K3PcZWvdeot7u61TSWytG1flYcyF5KX1z7EqEsm0KXoQu5MLA
dqHksPTx803h/Q5UKPkqHu23S9p5SaCTCH9ZKuvk27zEND5EzYRM0XczH+UUovQS
hmsnfPCeWmhysZkxPQgPdYa4KB6WrmXlXt3Ch3qQxLMXRwmbO4CElIj06XJRqRg9
Yrm461KZf3LS5+tzj41qqKMH2vWYkOQnUNrj/+vaTo8AwX4wWQVts2UWXv2hvnRd
JjSqQ0jgGphn1OvEx4NSDyVCVdzNZgI/rYcUHFlYkTBr2RGLInrbYC3CQuXfElQh
Up+JM2u3gMUGKstNEKQVSnQu08Vf09346Vg0pkce642NzM17eo418DYTWG6jQi57
I4T28O1RvhdJX2WV27MOt3js2ggniaWid+AC5IuL4MwbTnJ3Zu3r30oGkgE8v7g7
FU570kfuJh8odU8X7swu000MrAS+jzEEJHkuuvNJbaP7MbGI1gfUDNX8sTnsW0i4
g1r31J/4cdCarju4OiTirBVgT4Y0NwZxA8vaeZigiLF/mFtUaAK9zlrGabmOGDtu
p7FVK/CkylMd5fE6nImTn/VUXLr6Cwnj0pyraRmZ4kdhdlFe/gX8STSIzqTJOdG5
4zTB9v+mWPY/QcaCnboN6o6coCowLEEyvqeTtgNLaSBPvOQuzraW/h6DeTDBSeyv
RL4pUZWM5KiZwt6OOEwHqDaSTLX1HkewcCHU7SyBvP+JSceBty4j1uWIIAWhOe4Z
SqBxStWV5aF1GLIzm3ii/l91/b8V1dR7aMSwoEw400bxMK9egCpRUdFIeXdTQUKP
sep+6D5Qu0NesLYtGAH6AbKkZK2e76Y4iMNRy9LcWZLTMtsm1RuBkgUdl3oohn4O
/bzQQY3EZ96JbsM2kkyBwkdzBIDmKl6d7XWlZHeWBsDG0ennamFKr8NMavabca9s
rKxjlZ9uBENerrlqRTPGAhy0q6nYmk8IntZRBd6o2umhOBaeiI9zGlaKbKeN07H9
O5x70XLS2MRta3sS434HQsukJpqi4lH61qRoyBH77NmfpSQE6+T/DEMkWWBVPCmk
N+S1Q22JvTlWM+JqwkVrtgQoGgeTR/dgXpVHiG/jin7xUu01v1XHlaX9+s4QC5hw
B3AIoziIMo5SCVQnmYbUruaTd4sBMfwGeqbIhLQv8O27yuw0OvDBgU/c6YkUE3q3
8stNqHsU4Ph2qYv9oQEmyHT8Etb1SH0/dks1fLX/hs1meyooqaXdK85YSfDbPm7z
AnuK8KZzMjk0Gfh2ltm7dAb45WaMF2oD/VkwSWV16Qb5CClIz8BQn/wKvop5ctfc
DZ15pr2nZfLLaZo+rmKl02/fm2MR1VaihPM3PdQnN5sOCHAwAVZorw7cbr+11ruN
NPz0ilGOO37elxZGtl2DN5FwhEeo4huR/5j+XwYyZf5FuWRO8V63aA2/H2Taif7o
QvX3BopmAn7REBr8VXo6KFE2sxHfy0Az0+lMNEZPofefBqOcpP4V7zH2ZLoFiWIx
KZzIPZv+vg/9WVoBox95H5zcELgvdlKBX0huXm7PnVCOXndudjG3nNcl2DrNoO60
pdacd5iGuv25tcqyHzXurR5qOVkawJmwoads0kfeUkCCUx3P1Q2Lydrjl6qCmbyu
Nfbwc/SEb2LBP0uswT63HbOhBhrmGy+fLOjYWEMLUeLbJolXDZNY9j+iaW7xW+JR
sbUmkDLcaqzp+/B5Es4NQvtITE4DRa0fpUq0X3KlHXY/Y+kylxTjg/5M8K+8SLho
LZup79p5p+/9T75bm1JRbwR4D86DUGpVerp+UC/12QI46w2iXDOYyainTDgk1O4C
rmmjxMJkmXI05YwPrMDYizp1fDdba93pSFc5rVxh8P1K+ESJzodmiMgoRTP1Q/5e
DRjsRSpHueFrVeOQu0/dl6EyQxbvhv+9fvmtx66TnQSPVOdiTauZTiTtaMQ/7AoH
kLYoBusgCrsGE7b07TnOgf3Ph6fwYQ7864BGgb1hKDvGJWTx5yeM9dbrG08K5DNH
uBNzH0Pt2M6fyzsyhn5wNBCo8BbnqavK9kQtRgfz8xPQfS7PsqIKS8IzKbfrr814
7jUNWMSz2bdjsXFMexApoextQglbdkKO6rRMN1i+bQer0OHYswqc0I9cRwR3FFSp
zCBoRgckA6xyCsdVRPj5R6vDmxQYirAMmL78RTBljWUFli71lZ7j4tJv8nFhwJ4A
1XKCEbtFv1PYAcVapUV9ND5SN5aJ+PhjGYrOTNpoGktAiyfmmPj1Sk94qJipd3tF
zLAOlujreLbQox3CBHSimPL5IMZ4JQHX0m40etXzl8coDI3m5wWJuY9hWMpacVEA
nWvMs6z9phOUZ4yQGe5JGTrXysAzbgtnq7M01QJw7WvxAvfVtUIf7VKb1iGipITb
kvVwukTqI4XrD1/c2wLoW9qwROmsVQTGeLNUeReOQsFJIKmQv4yHUOh4GqBmF68F
ZJDrTL71ZfEEZTLI4xx+m7xNjgKTrkRYzEwj8YhsXai9hiyQmFhrm48nI7zaQ8U7
MKhISfgydp0oLtf4dQK7wteNtaUxZml9NGQCYEenZzR7U4M3gBzjJsBYi/PKgX9F
/W/xyTS77J/C4JAkogjy8BUkkVXgea6NtpBy5IVmI7yckveZ8KOrMV6w5ANBO9hj
aPjdw1nDpo7ZRSl7RKV4/aAftHX1WpQRMiBxQRLhAtzNyIHZoCt/omDnznO4Z8t4
3s9LR/eAcnMeqvOwOmq77bzjjFQp1Gygn04bEpiPRFqYQv7aGTJr33hI/7bqZGGY
u1KotEf3IFdQkGvGOsjHkUadOCNzPsTZQ1u5L9np3yMFpUN+RPRwN/sb8yHOAjnD
DCH1PTkW2HtqFh5KekO/aEnaonX2AqfiSHIz3FaeHAahySf9Z+2K/EzoBDekoA+t
TMMRDDPXeOUkONmrUBPw08ofTBph4xKPpfGEr7VvF0sN9RzrQC3ecFhLF9eiDtlt
xcnaPfZpk5BQD+u1CBTEN/R/I5HY4u0YeYYYBHCV3zsF+ZiQKj0VNNhNtzGh2qLI
Gde757F5z170UyNLLtf4zyL9JXu8oIa2I3fxBJg8Eh8IRPiY5X9nAwetyrx19BVX
LKneaL+mikPR0wfmgiWOHfuEh3GbbMygahVuGdjI0Db0LnUR48bOgzjrN8Tlb7NR
9TRcRwPCbyiouJVEdSLQWa2o2SZRCEgZHVR2kk2kPV0FAvCHYH/IhiNvYncnzEp9
eUIH0H03PByZd61Hgy9N5pto/K7NiCpNoqYIXorDLvogjGpofSY6HTpqba2kODof
ItWAJXCgYXz0JUoLr1zQCNWPC7DLf3uN4h50ChfKXcMF203MefX3I+elXyfioGEc
h3xDxqN8kMAIK4JSFoMEV4GHn/CN5TulZL9fOpRHZPbvQA7blwfYBNZGE/B4AFVU
EZhQA8gHr8XB6us/1RPFotTVaZnpsabjckIiVIAj1GcSFCmpUNWbantKfEDGgoGO
QX07J/DUzQiMoOdr3mnKUMrgNwEHKt0CkSIA22wcVSNyLBGgKjLW62U7yC7p/1wF
aY/dyfMtgLSmJ0YrzQbHG1cSeHJzsvRHiXQdZKOm2N+IK7nBD9MVCjucKGwmwKez
xF8RCuTq0pSlft4AG0zeLVJrVn7QdE36Du3v+CYAbI8ybyMHHlCmkWZo48cFl1dM
SdpVMt8IkoxyTZx4GkoqOARrWpK/jSbMcJaW+4eoauEeZyf+uepIT7/KRM/2b/Pc
NgJJKUP4BIknUz/x/KaBb4GdRmCHcQIZHcsGhKrw60gql4acGtSkvLPjgyYsinFA
VdkJuGp6rY/f3rRKwHF0czZxWdIJHYJHN8tm52TEYznf7FcvhytOkPMvb8IjzS+v
SvvsN4kXeASr049F0JxP0LGSb96UfznrkN32uglcTco6AcBsicLIzB3d9ljEf7Qs
7jwqTE5/BC2iYVSnieI5Ru74Jjm6jxp5aDjW4dNxX9Z6ZcdIh0PGwETkVglGieN7
DaMkPz0O8UNs1hYSaNVW7AWAmfhYWEzk9VFiqEIs8dUu6Cr8sPEaAVzRncg7/8nD
NtK2mCrfCotPzepsanUHAFhm4bPmINWOb1o+AWVNScPDj305x/N1UMte6mW1YfuU
6WUzwsoydMak9lV3x57vhvIeW9sgIhTLPcEx3aeNhkm2dYvhlF8mkbuumnqOoD4u
3x2g0Hk7/99ENV+9fvn9tbMm4uLHDkObLPDFBNX2WQ4NZHo0Rd4+Cg4AjcLtYbpY
pU13XOrp9lW/oAyBe+hPnWBVbvPNU1E5cZC/Z8BoRZ8IwDmlg6XbtKQ7g2TshJlk
puvnM0wlXBDy+ebKJe4H2BF/RRZZxXUDIFeG2DDbeDDzCHvRQPO9Skfz4lrqQPDc
pUmb9s4Ix8A0LtPfj8W4ol6rKkW/sRAk0VNA1EUr1fgS9zHYRbWRdBDbSyGmzPBJ
QocgB7tqmt6UfW8ag10xVHJmyowIpwPGM+EsqoPVqj+nQoKnfBt26Bu4TjofQBKB
4/XzaM6ushlyiiIj/H7fjz9XXqS1ChoSR70LAmtJ+7HUcyT+Qcb89xHqNuIoV9Qx
2mMcYH3H2uR+3dRRH6XljTnmjpr9TbXzbxTiaiqP89bYDXFukQsUN6QzND/ZU2eN
I4pGrUTDk4bb2WTzys+I6XzxjHOpoQZqlB65ZarbBs5qhL0QOC8anQVTUscg3YJr
g2vW9dU62K7E0H2K44qh6mNh+uwFCP9fKnLXlPFkE8hwZF94rLr3gpHtVqWifRql
Wi1CpBEDVl+ap/ovY7tx0LtH4W0j+vbsrcdE8nZaPGrUHSwh88HFjcR4YHlV5xCJ
IgiIQsHYaQYjw6bfqQOEr5KXu9Cpnyes7nXSIn3CGik8zRsk745W7SoVxsYBpRqu
Cc0hkSzxfOvPd4t3fk0kU/BsFypWc+kxd+802ek+N8jY47c5pKPfvTVY9mznmyPy
Aah2h71RZIKU88ewp478kXnLBlDGewWXHVri4qgouQvuSn8yqOqHPqQUR193VNxN
Sf+TlAau2rHob+Z8eDsI4hv5zyWXLJSSoj43qkPo2YMulKXehlXtxD2k/JVqxGFa
YLEDlZHpBum6yDt2dJD6fJNXdYH1raN4FlQ0iTHiTqtAKW3aGqbDe9e3Xk5G0ibq
7+xVkTD02SbAD31cTde0pMqIEB1Swd8kJCGhq4/XljE/nbAZAB89v+j/MyVCjKoQ
tYTljO8r4+LBNsSKD/aIyzfUvWIF0z2NUMXO7b/eHpGHy8clS+SlXGFy1aIH9MN1
1E/IRWun1kh0BpOa5H5RJRYRNlUXsMILOF7pZx4foAJydz5XkEsIw4BM/DOufRBB
6DBWeYSb5QChFO8ZmA27IJ2GuxVrKR/dv5UZfwcXDQdCUCJ0OshOeRpeVooFGYV5
8QkoEiQnMJ/uly006ld39hvm5vm2RytPPPy4N0IQRPghtzwPGradBb4HgaGstgN2
7PBoEA6LqYpB+TVFiT8sVPyhyCSa8mVKHNcN7h7tsT2HnCOmrvcC00uX9lK+xvTv
dBiEPmmXkIzPsc9Okx8exOYXoyUMlb5VKeRL0ogHMN3eY5h0BpatNumI8unLKC0R
TqlvRihWgaVe1KBwt+PlVKUCF85Jyn+OK3s+ddJytxoApbW76wJDC9IY6nGcDywf
JFJHUgiD8j5UBoImPOBP3dz/0zcg1aZ7UdHCMOtCIGbPe9joeRBf8ssXz1QSJPEU
kh0nhtOIR+Uh14XxBpuBtcHZ59x7BpY2akqj3wPwKuvD4B+rYKLQn+4/Y8lbQY06
72RXFR8zH4/md13WXePs3xOZAgxazK0knFTIodJXk//oTulh75ESy0ZgbYVFc2Y5
RuU9lnIVjxqkHbgmyT7xczvomTuKh9RkKPfhE5+BwgQfCWZa5ckwviYscCGNP7LW
4yIZqtiN+b8SK6yIb+sDeJO5PSk7GdPBZGE9FrJd4/tAKbU5rcu/Y5XUcLhS3uKw
5oU6srQI85+6TxZ55RyOB7liMi7Got0G6Gzb5WtvwJ7E9CPtQIw3VxgsTMtlKgLw
bGHNiYAt9qTiL/pczPqkNFXHggHrIe26DA8BRv13kc4aCkeZDhnM6qImMnvtp56x
nlo6NFJaM8KPIjHk4wt6qMncs+1pFTKyTZd8RTIzRx0OhG7v09zDhd2Pla8brH/F
TYpNz801egPQ3gNdg8Xj2EYQ36ZlWR0aYlPujYuUOzI0a0orF4aC50nQNEaOMC1+
Pv2jpgQwMq/LOhDKBlZlAEIi9nQUC+9WkBBTx+2xFGMWXaosNNpRLzAzSiMmiUjY
vdf8XbcJ1lQfEkoTEKg56hXWwLADzhcGfcM6jpb5EdE3eFR1YYbWsXTNUhKTQt+d
bVYWRKH+uASMhitRTY+5avw7Kgj6YlQ0b5kFZdsTpfvpwH/LU0SI9D+wf0/AQTyT
FFs+ur1CJ/EZ2D4+aozo108AhKnpOlhLIOV60IbgeGCwjj34vYwlZCy3eUe40M6C
lUgwlKLGP++hKb96lt9yUy4JBlwobsLgRcLQgiwVtP+BwFIHdysB1QYQijaENVyh
ELjBzQKYOtEUtLX+XfvJyqg9gpii8fwQkq0lylKKHzSTSMJ47LrCaR6VYidXNL1E
gPDsC6dVQkDfscni9PQLz3XWrg9hoSlr96ipJzrRNE4Z+mL6kKMaChS1s7ZLWnj/
KyjqR5+wWrtzlg095NUK10sXx55+vtsezMiDyWlUJbuY83W+1oDKtrKOLbA9QnB1
0oKYhcFk6qSAbwcO4hl1swfBl3zutR1AceNrbyqeAJ1Pz6bSg5VJNbo/lAUZI6dT
LN4kj6jPWtblzvlta10V7qcuR4FYpKQWrtXrQJ5y4ziBnRgAV6N5aFmHNprvVCqu
G/WbPyfFGfYG5dcCxtacGgLKlUqY7+snCLQePD5+sVQy6iZDqtBP2+idllnQK9Wp
6CcxiW2yIFUehVgQWyMJJCJWeKJxEl22gmdFy3wBa316ntRx6YfDlssh4Q1XQ048
P7HLWk2LoJRuq/HNWLyJ14ufHHLmyoCt+z6srzxGVgd9dYW57jYHqLL01MT1vx8I
f4r+6vWsu7kxbiZkZ8Vxcq8UwxMINunjZoh4U8j5JpsU6/2PyJ7vfO0+u/0kecMU
FY7IJR2mkAOBIu8JWMADriEBCBxDb3S76CAbM7ryVuyqyJhWbiJbomfr94fg8FuT
+hSdksi2BEYnf07YSe0loXXJyZW7HfeAcMbTdR5i5Be1D52qg0nra07be+n3LKzH
2SXjHaxV2K0D1lZyVMGDpmtrUepTe/AIXE8cK6AIOeqW5yi8dRebjPUPtvKh1M0K
/03+afdsIdIgKp8SzkNzplsZiYdF+YFsWigIalRFPwWBn7BrWM76vYGmxyoey9fA
mmRlBvBjCckipAmjANICqwvipJSQ5ahvTS2N+Z3wGPgNqBp8XvSzfiBd6jSEv12d
Vt1kTN63wwUy6rg6xcxLs3lcoMg9nyFU/xaTgCWVcbn79CFIjc6XDE0pvNTIsudB
pratj8npqxkHbSLrSqnQb8VvX1ilDva9ODH0V1djfR8A/aKdTd0liyNxrgCq91B4
k5qmCso0JWMVJLzpnNRJ0OGPtikDJAnLEIgQ/RCRH8hITTFa+Em7P0/ObyDMK1/N
53dcPOXBBQaAwrUdTBA5F9xlCD3B5fvFYpADwEOad/Lt5xZDUrOE8/zAosTs80D8
BtjtZdN1Ypj0y4Hq8QISRw+r2uv7RoOsTxQ9nJ3EaOQJPaq1/N3hTchfL2p33dLi
O1XD1ZC2U5Dx2YHRZnfaAyMwLjDBkuM6TOKPQQRayk7HNr/zxDumzgbJz37rtHu/
sMHQCf7D3E16+X8Q4+YK71czSRirLgdhml+etDWc+utOrQ7oocrU6lPP9/FLePso
/AMHveAbtovwGIKYqWqb7AaFLLrwFHsztpXtWVtN8gtAJV9nbyKZZbZOdQprNGws
tlDp+e6P9c7F3zDB9dhjka8DhcU/3E/vPY6qZpgVejmiLkb67xWpZixdpcls5yX+
MSAF28fC4qT91wMYMdQZDJLPxs/HpdcT45MNhPLTQ1uiH9s+N+wwYCSM23mRtWsV
H7CXaFlz7yWGZ+TDx5FdGwjvx6AraBIjx1FI1NcUF0dw+scgo+heDEdDb+iWjAXy
ulmAGQrY5VWih0L0/1l15N636cxZj8sjq6O0wo/53gN+ZjBTwf9Ee+h7chxPzAoz
P06hJUhqoubrBSC5k+NcJUi4Lr/Fr9FGWK7PO5vO0TntJ2bPZ6zmSesNBqX4ik+W
Njb65myHaCGXt1LwUOiMCiNvEl1xTOpkyJPO9rDqwD4SIGJVdfwk/pTXR17jcn/s
6uY2ZNwvC2GT0vQdxX93gAbqCOUIL3uqgLSYnk1S+/lf5EpELc4wW7lELiJxqUa+
D7zRCJHA2zP315BYiWB0ohPEogbJWWNug1FIihXX2Lsh2lx5CD3EBS3nyOEX4/0T
J3xJ/Ypy1BGUHm/BRuq6UY+dJ/1E9eu1G0MdcCihujqn/Bi6gaj6GggWqVh7CX0y
pWowEvilFYmxsWtrQVTimlMOs29gPqNPDSm4HXqFoENCwfoR6H7D/g7TfLQxNT+O
p6QJLXnO5s3Qd8kAvYrAxAVrIDlR1fCgfQRZidKumJwd/ZScD6aiJshqlAFv89ZO
zNcfWnjGGV7IUvdcbGc6Tx/aep3f4x10Ew4ypebJuWFWmWQLarxcSvKHCU3NFnji
1lopDdqtckmfmIaVEGdTMr6oWt/Yyvhdbe7ADz1t1UJhrB48Wc7k/c7+FrcdMxTy
YqL1zA8UbW2pPv78/YCdBfWOKwLjFJIM/o4s6KKin2izHZVkoUZUOsGjnS+hV5Ba
/ZeAZiCkZ35hQP0l+acr8ozaBpt92AiBRCGxH+S/MUE3ICg6CuRmLZNqTL1ROr5+
ewttLA7VtjI31awjjuHp/ybg1ft8FFgJZSx98c5ABLq37kFs3rcS5CYjtWO9u07w
cvAYEKdwZ0vNfbntonsMACFrjdf5FglHeZwFGTnAe3QzoGdwG83O0nL+6XPkhunp
1vf749T8b1zhA3CWihTnSFn7O8sXmXKaJAQ84SUHwwZrqsJFJ+5Ugz7ZWTqcX3de
dyokXA695QoqHDvpWUdMeNrc20wwRaii1p6KbFXiq5HoQDl0eILtIpL0q4VvDHLa
k0JKF45wcWplivI2pYsiWEhTtN+mXzyiru+YkV+KoiVFp3OEd7dG8ujnztwcYQyH
Yo1cuCDHx0v1uY6MgeoUhMUE4VDS32sNzDZ2n54ENXqYR8cmxgW3GY/KpHrfb+7Y
Dtwd1swfztfluPZvUuEt7wbLcNY6IlaBUArCVRr05WLmuIhw0hBpDodZobCkFsUM
YTEDDBbssCh4ca5r0rn7PXVgo2BQDYNM2JYCmQbdiyEOkVmzgBPvKMd15NHKLIAq
a7/hxCuM0sJcPm1g5lgA08D+J3+3UsgcrWP5z+OnuQwSLoDJsEftlyEBbVZhk0Cj
5vJuIpczb6CZ2w3D+06ktHT8vTLQs+jHPUIC1Dl4R9uuMKWdlLd0l8RkoXEQpJPG
dBn7mwFK71qM+D8ogEeh9IaggBr+hcYm3mvu2LStfXBIfLyaBLtkBIeN6ZoIW06/
EfUj5IHIl6JoB3ZmTUY3I2LbBYPONYsz+yIABDR2KW/s5tsrnYsgHa/0PHJAgcgE
04c+cxDI3trFSHfg+Yr2bVT3ZGfHPQse1JitHzjpf5i1PEdZbbk6E8SqrAFM/qm7
J9OC1PWDu/OmAhXxtzbBmxr7dNnTuewjZD/GVwYU+EpM46263hV7nGXb20ptXZkM
ykxzo8HUlujJLo94jGCnRrP0dAWU2DcjXR9qCH8Af1Px6/9pnheiEfpMRHeAgNTo
AScZVkfCe7SGYSXMDOep1HxWp90vf3I5HQB4xkucBOOY+9TbBgJNnVMrfsTkNyeH
IrNVwYtdXJxQ2WsIaTKifK3KNhCYhb8Gv0xlfZ9m3iHyk/2pVIvZdV0argDuUnqL
4UFcraaCcCFc9CX0v73glPmOJx7Vt7FF7zBG7oAuR2m3aGwlebAgilyoRTLTLkY3
YsDo+QWv0r1ufnw7VJDQOqVfRpMFOXD3tIzPB6ah/VSOEvP5Yx3l7iv5LRixffqm
BbcXn80aXKMliub5pu/+wJM4Vg4+oW17Dgt1w+mmxG99QHmovFcI2JL9VLZg/Utz
j6z5r3IQAwgE5J7DMKbj0eI4kIouzxlWsrte+usHRfmv36jnbOs07UB4HNvo6B0D
Q6ardvMOcnlE45JR0hTbJU52m6jQwC+8qTkRh5tK5DkOZMsyRJ2qGikMTISMzUm4
WsonsWpHTRR2LKrUIlcisye5+llxWp8+j74JNjNn9L+N63gwF16tluXPveweVgGb
x3nvAkF5HYeLhJOUiJHoEmjVZKNq+LI0ThzRAein7BtyIEiqrg37V7F1o1cr3ECQ
rYxiK/jBPFjDKtLl6U7bGwIPretct6FVpEOU3uNqz7AAqUdP8Tz21DEpJv5ebln9
ZIdAiuTpcbmGqUwbLgxvbG3kCwAv6SW3C3ndo5TCkAFzdsYtv0RvphTG0qG7XkCx
e1PnXMlBEEGQbT+nY/6+KYnzU92UC6hDjnlnGYSGEcRtP+nzjt4FABS0UF11Ze2U
338sZYwQC9R4g+G7B8H5iOHEIYpoXXT5tH7kveJxGjuBlsfcM0xD6vhoc9Puwq2Z
gHy02d30/Mb33q5EtC7xrNHgMpeWEwb1cYt74Y8se9cUouyv3j7OheCdocoZxg8t
ecWW/ek7I9pNpvPRfXl+BDz1hosa3BCPPbg8aV9lD/Q6zQBFxmrtHV/dusg1hPuL
YKj3ODq4udjlbIG9J5hnllJ5ucPXuyorA7JJhoMkDw+kOL+1wVSXgUbTfNFPKsbr
bkPsTN+bRgG/ZfR/J/BK1nu7lNI2uSVdLOI5bpxw9zyVoYLPHIbU/XeNqSZrbbdR
MPwWGRQXSo1vzT0bQdmcrc2kRO3w6oTcTXdkxLXEdksx1JRQ2fk94oqsk9DYd/Y4
F20Rfeu9tDeEFDWr3989PdmeRcwkxmqRJqGar1fFf29jB35tueQGzOHjtvcse1a0
jQqZMjb1KA0r5xxZzcBUVRiwKM+WzOgsSpUP803rP+a+qBKzkLkTzXKFlFsMakqQ
uzTFpe3LL/xiKOln8UvG0+TU13qKIdmD6U1ppI18Dw5qbEnoQ+RPq1ksQ8zx9V2e
1KsezF8kO/OKyLnSu7SSzEctFxd862Vmof9JrQdA/17khthH3HZlg2ieAtXFnm9V
I5c2NfT22usgEyQ6jGlUSYZn3G6ZxPm6DpthiTLi1/W/LipECRs30f4ytB9vj1Aa
xIqEcALz5rPxLsas7YiEaKQ76UOxsyn3m0hCUCXudb6OR/6VO6zQ3o9+PdY9b8oN
6VITCP5aBkivThODxLP5YgHPuOvt8YFrBlFxJWN3qtfaIU0e9F8Ftt3jVdsYj+zr
T4qBQhzXCqym44ljrjTJL9h+Pm9G5DDwu2tC610C/QPR4tigpH7/IGPAKBJRXLhP
rr/0I5+jQB8W/cpdItntYNCets0qPKDJnYG+5xfqL43+LR94Fe+6Mu9jV+WdJbBs
Oiio0SZaX0Qx57SkKzXCskyaozHrCf+eHZxWpSkMldfXAd37Ddg+QIX+iwCYJxPP
GwID1XX3qT+Aem5V+VwSFvD3ahpNd9M2KWk35W30bLs1ExSCvMWrpdMY9h+HWM+L
V7oHqhX4nVAJXTraN03aVQCkchGAXRRVgAhj4AEK2D1AusvitNs7H3CFZ263W3Za
GR2furbs96ApgbS2OjS9cPl4KUb5V37w3hJnrquvNx3DxKDcLOpUZxjSS2hCh2lv
m8LB2qdBRH3o0VW0dbEOMaNLdhHxVXz8j/MvwmeG829YWaJ5dQxTWbLooPy6tMQ+
4a2DYtb3ttOs1577t1W9KP2NKf6GmYnNJIA+JbI9SLdICx3xd/A6/nXSX8ZJXp3X
sIHCP0xuCOSNTDG2BWXUbrxGHw7AVFw5+hcCVaeqtSAYxtfqfgY3KG0HcYsZ2zNV
nMRNP/w/hndP7Lyu8ifKsRmoA+4ZZgI8Sb/NVwranlUP73yJxZkTHeeTU0ttwvLC
/JZtv2oEqSFM33XiTu4uoJFksxASr+qfzQO1lg/zdH8IGbTzElXY3KxDQQhJ4Y39
mmiaObv8mQpCC5bL95Dx6AjjC16SOm0bR57yJyQ86ir1XEfjohRK65IrjaOC5MvD
yflhygyOw8sbGxjdqebiae+gfrdHDwqlfDbfRlwugS0ilBncjKf/ZkOlH9Uh1KhO
iNh6v6T3+qJDggqAW25onzVNgJOovrBCY650LO0vYonxGTQKSaJuBB64WeImWwHa
z+LKwS0fjarI9oPMWlHCD2lh9O5Juv+HwA0yHveqoouUR6vBgLo7cbvPJv7XZOiO
WnsB09oB4twZWwEzUy3IwNJYHVbMVzbbDqFzybO4V2FYD5rXQX4+i39CrY+tT1V/
TIBTZ/aaxbuYmQniUw4TGfJYm22uSp/VHwybCUAxekm3Ezn9ZM2X4Vy/PaPk7AV/
yRtR2vihI+ZxPiZZ+AhrzVAwLRehvMp2fuK8YHVEx4LXZGLSXE2ynPuc/JC3VwUX
YbsUN1zDje/B7Or336N2tqJs1QCdVFxmFEUDaEl3UBwPhE9JOSZQN/AiMZHzyJSC
eVai40LuuAgWOM37LvkQwHpVN+hBfWAZ2JNlcaxWzVoeb4JcAkmnygiitqgCblna
74om9JWit2WTcZGkr0jTIeGyTokHX4eQxw9JesFjx9A5zcpOBKoGIcEvrCgE9Qmp
ifLrXAvEbY3i9Dn0Y9Wv7UuaaWPHtx3unD38B3p3C5hsRqLt5/iqn4s0Vdh5Q7wk
t0OyxXIEW7HOkI6FVi/x3rIp92KS6TGiIJ4SmyZ58iW8yoAT+beJMq8azWiSsB3k
4P9mAX3J9ptEwkYqnJFk483kq40Aq+GniGZFpiqF8qYXUi8ghIOKWmmMtoiYiYcQ
0IrGb4M8nkbVVK964yuQBBrI4MQbQsXEpQeZhae1xqnVVUFXeXPKqinjqCQmYLoo
w4SIRZrNbRAMkAwPw+SAUuWIYT3rgT068DRoXAzsB3EWaEcjgRUR39VBOEf+8qAi
Is2vEuZVRKJDtvhmJUGwMezJtY4fNfccNOurmBeaQjg5M8HOUnQsoYrOf3ttohM4
K/offiiDpefzINixVja00fVIMt5APn4oUwoYjSL5j5BZ3jGoWpwcGiDwUF/2OaRa
jNHldQUVHB5IYlqv9qYKNcU3JyRtZKuVMRyEw5tLJMNwXCVbdv+RZj8L+9tIi913
XAXUUS4K6PrVA9j9b8MuTEjJ0rRS6n4fkwMsBqXpPi6XKF3vfm1z8b3oL3FoBwrA
R7jcUa7Icxz34KyeJVkDWqfxqcbbBBPY1B+KtN6FPHvntJKluq3TRSfn8THuH0mX
8hFNNHfJFreLO0ekDJE4M0AFr6dB452gxOJbT0u/ys2QXz+sKaj1pHKJwGCmJPim
cCHDeqy2WLnE3JLRpT5G2+aGIUuNFT4VL76P7eFUpjw4WjbSyWyBLdwGuWg4Fenm
eTZ6O+CZGGeSAixIrhFgqkSMZ9AoSrSW8P+IZ81yDMqMDpZPxFuL23qo1+OayKfv
VscD/MBiv4OSs6+hxJMffGK9OOnUsyrlMf42/PY+omNsb4SdJubWe0BoAZQP66Fd
OXxOOdakDidZvkgpF1uZPAC+lzAPDgn07+fu4lSQ3jWe+zX0Q7/Q9dJDU4EQXnq/
C2HPoaktodKetzwZigRQg1MmT1n6ASeZdMpni6J6ItlQFSiD7Ffyl9gu19qvmUwI
cuah4Wwh4LJ7jhzrlRsJ6xpCPk9T5dw93CRG06XOgYctbCiE1s1+HDCmZxAbqmqM
bNMR8LZZfstPbF5ta//CdbHLAodd9ej9jrH/5KFMIVi2aPiDj6RKQFEw7MM7a9Hi
xVCdXbQUJ7Gdv5DJGF60pA73FwD/2Lrz75S2YGsEg/jrRLw8wAKK0RZKUocnarb1
j8U2Yh5hhEBWjxy1gKv9l9J72e0tS0g76zK6+tdnwHucsxldnoWOP9T23l+94nnc
tR5MBDJYnghyQWkLgDxUNH/Hf5IF78DF21CzV3H9k2rai7aa2qQrk9f5T5QqCRxv
eqzswRJpItYCjWiZ4ZmWCDMFziE86ksPk2WnCyz13GKSqqa30weTroBONXqnsAP5
UPlWRQUEU4YpJyiwAFI/a3NjgmrKYH4VpUFkWnT+3ufR94XJ00a1GdglBcCKJ5GQ
nCOLXC53ZPj8AAWzRmJYYaMcjBR/sza5IBaUCwmNTQWQDmWAgf7CtAM/XSfQv7Ax
suM48lMsrcHvwXc8pIOcGXERXg6wqmK6cQh3+Af8ltG7Wk6RtGB46J3a9opmQqiE
rnDIssghretYtz/d7akFdxkc5VBwnxJvcNOhJZSwJckGstrzDEDH5CTH6hoYw27X
MR0QR/t5ofF6f3UGhVyrPUBPYERA/w1qaortGJrp57AQ/2Cqn/iBaP/DJjjrpg7j
1ag1YhsrKi8nz/xjcNb3CShH/DoVo552gwEyBKe8OrGHZpVF+H2sycNeBgEmcXZ1
r7nVcoen45HFOLCSWk/P65NMMj7+Rw7rCkF4oyk/50XerM7RhM9+S+yBxlAzTZRv
FCLfPcT18H9ahDjNtr4MI/VahQFMYW8f/IEGLX508Dnwy4fXrYBt0P3f1roRMuvz
RUYyaAa6qcc0qC7k7gnjelTJxi5r5Z9RgBt3DtDBKz7ZgRlQKh21Nn/TSinVw7d5
RZ8PHZzU1kLUuiEIX/peerpL3VC7FXrRvQX6qhkVr9p3hvrffVsrrM11PvCsHpu8
zYjWcUAq4yeb38ACtU9qXTFs4E+6V7hkeWcf/TAE0MyN0xehVOmo/FtduwvxC+Yu
SAkBQE6giUt9SdKrEJJrl45rkYdZGQqDwNvmLLXEhSrp7PGdyxzddnSAIkhOek2Z
TZ726DzXiYBTrQuzManx9+PyGBRVrVnZ7rIn08sY6uGwTkVL43PpBcRkEHczCUf3
+wXCdSVi/ZAiVH0OgXXv+5RE/fziU6R+xq25ljtRMutQaCG2JdM9nGOLJwCbKDtm
5+YndmyC0auqLT3sNZrlCC18VaSMfkvQHJBf47SOS2BzDjeXSaUHTx0GK3UlfbXJ
CboS3RTFFEApq/vT4uV18eB0yN+0cbnbb66MAY8WHZ46RCKfZf7XjknTklYYgjnw
PiLxyC7uslZayW5I5iVr7EB7QbP8VhUGuHxcRqjCBn4OuX255nTEx/BOCGxUSvTr
dcJMSWZzNVAEj6JTtv/KXn0YifbAmsDRvsO4akGVOeQn7iTVRSech/8Yq8wEdZPq
tdAmAseEw8nyMciqsXxxXau2wAL5pANthDvlPVrmQbgR3GU6WQ82xQk7eKsY/J8l
2hfoTEcV8z5PXjsGBWw93E39GuTTUcH2UXKFoC03aP/AJX8SJWJGuk+QVWb/IqBb
TTYPebzf2SYnCrzIzF3T91GV3VpMhnURkuKVo1JSSZUe19InnESpJa+FEqOTRjGp
JeIdDHrukUn9EtYj/tbad1uv/veygx7eep7CT/3awecyO+UzVDva7rjeErUa7QMV
lvjS9axQ3tDVC7+bkWm2JY+RjhSyMpVN9IWlN/zwjCikcPnz1s8ztPRYd9gd2q0P
9qXDj9CrUsU2dW78bCGNl650IGGSGnR5+sCAqEoz5P40sMZVTyzMcS5OK9BQdKx5
XNr9KGhvcGrucJLdfNBt5WY5nFky+ZtlZTbeusQ28vXS8yIvc9/xdhQg0IyjDnkD
wJ3/I+zLRgacQrXqXwfvO3rmGQ2LaTZoY5ZtTqlIsIYWL54H6nyM3xpOzDS7cBrh
hWR8pxGhYB3+H8c9jt1/b/Yh0lir8RFiPrtN/exVV89cGL/Oan1wiSllLc8QqFfv
DedwBK4QAjHjXpEA7Szd4mA9rkYjKb6q+GT5X73QpQ4ngkrt7jXMEcHA4HZo2utc
OZLomUeBGX/D8v7BJ6SAdDfW0GQbWoL+ABz28nzFfCyyzx8lo97wzFB5lBlFOaSo
kAsgVehgCxwBiTCZIDOGWf/32aQUjk+XqHJlAnClR0n1eLlQuSc6RXQpM1WIJdqb
qG/CvsnRMSBH0UKXySpbb2zmv6isYUHSOh9B+NS/dtoA9DGYIvPxLpFBk03JBCAA
WdkhTVUWyjtwohU9hunTXSWtvgbbSCbW1Sb0q8XSnXdAHSLiuNakHRC3uZzsqpTx
ity/hMbrGPjipFexSBsk8QZ4+v7XGCnEOQYBB3cVrYzZqg9fvEtQqJb7lv7mIzTI
mVLwvG37CPzrVgVvQYNe8mNadaPzlU1zHqdAcTe5Qc9wjuZr41c0Jli+6Bewu2q/
GDr0DpWDcRtmUAf2QsV1rosvPvIo1+kXJu1oMHmfbf3RBAGc7tu6xCDZKcY8E5QM
uwDgMM2JWAxbX+FY+nWKlOB2V7lAlFCjh4jwSf2ZqPk5bi1Fe0yDo2Y0vENuK2XJ
gXSwnVK0F3oUYnwwX3KyrX78kfpynUPHzakxMTFQ3vB0TgxnRxb1qJexBbUY7FJi
wZ9+NnPrpJUbh8esV0O5LgMlcQAqFopkbY0h9JKfijBCTMEUQeL0KtyM0+xVy/KQ
MN5Spv70JZedllN7YsRgd2YG/K6yk3UOwUtyqT4p6e0xi8gg5F0pArspLQlrbrNc
HCnxZf1iVy/Xo9taUgp+N0AW/arOOj4uCRETkJV9TuY+XYrJatY/vwoN0JwmwvW/
aLEhElO23rhZ7FcltQQI6RS0/9TIlhffUQb6UMLeYCYVTucuMkg4I2mHJb4zO4KL
h4IYCUgcZMrWXKuWCGoBCKtoHO4kIAecwMadv3i1LeG230EGV2u973juEv6K3Sui
XOmRCn0KbrwIFxt58QRods/yLCxFAGCk06ta5I8ie6eM9VFiPxQZiPHRy8I36CLk
YnRujfN1aWiNTZMwCZg+v0NL8V9pV4fSAgi09M0e+7SDoWlgkF4KghU4QMQnwVIq
D9vNx8eqWFk0yBQLRFEu5Zkfmrc3S6IDlA+s/NyarRrPUIMH08JR1FcJp7HTKh73
RKLbNu/TfJO0u93Vy9f0G+luZJ0X2Ioqzzx503fLT76inFkGYEfvkkZL2AloLgC2
xAJvm5GngXltvKuJLyAQ5cmj0jKhhyDHkiaVMc6Xo0ytwInBwJGdlKiW6qKKpK9W
xiaWg3aj9aexhFqA/bCgaUBQT3Wv2APx87AUeheto8q4J6QJUPbK3JV0LSMiQMgw
/3a6G8dtydZtg/YEH9iqQUQXntlGh2HZgc5mVWLVW3THiKJmJtmdjrOlYo/aY9Ps
pD/8/wixsaY3qSYTa7oD9XWVXKBrnXUCQvA3nVPbzxLq0oekCR+f26G2+r7HWnsQ
tBqqviQ88VCeafYIao1pPTJ6yDl/rpJm3Codl81fKM4F96DyJFCSg+lsCUxBNjO2
yLJQQWwwzD1X947Svxiua9Yl310KLZ/So+zBky9DNN2WiRn6Q8S+kiuAm/KERTNc
/s6qS3x1zgki+JL8ScvO4aXLKh0Gy7MaV+3q4vrWQr1JP6K/dwU8oE4zar8oO4lj
TEmsuWT0T5vcUL17lH8nmORNYHOmq0urNrFsrDx0WDJcz+c5ugFIRrjziaESchfV
WZzqsl8tkdsbDEDCB8RjhBcZgbOELQ3s/3AD6N+ZAj3MFz6rleXlASZz/TPCUPZI
aubBEPF8nqtorVAdCF6GGr6hm4EvSfSDxYll81a00uDVvG43XecboY+HBPu+FPTV
/MZLWe4HJ/i7U56xWOC1Sm/sfHpH23/bEjxU5FzZTi4DeqyjCXB6Z+ZvvrReA7ZN
AFS9g3v8rAxIA0oWZDPovGRw3a3iwT39thTrLCqk0Qs2DsAbzS8KjkmSRnHJgToD
UzHQPd//ckcxVc4QXOXqyTPVXoaw7n2hbNHaEwigSVA1JqWy3mcdEzKAvvLBmqQY
JdI8FppfkTsgxgy4RrIja7p/qxPpAtIB7b3tddjRIxuDCtCzN7BP3JregBbE71es
EKODhxgPe/5H6nkb9dFNVfalarEyqDsHts9HqfTOSHNJQpZLBI/hPlvZD0tvMyKP
dc9eU0JPphn768yRV8rxyi/y0J6zhMUUd0nDcZTizES7D1WBj90mVKSAzPAd5DyJ
VV+mGrSyHAwjzjj/vwtk8r3FXTiOBs/EGzX1XhrzvdeV20M8JlH7p3BsGJnTpdCV
aw8EpQMGH8P0lsdnjwmM9ypn4dX513zjdUgeyagr64r1JsdYbTAjXEvujnuEMhXR
qWOTf5Pi+obWHkjY7EZTtrP508JZrCtAaFQdvKH2FTKStOk9r/pFGcYiHVy5V0jI
1ENUXegY1O3wTCJ1JxkNuryOdjOO3iZU3M1ndxEvmGhfIDi2P74Tx5pfrGTPkvFj
0VSUqsw3oR90jk0x0tCdchjnDkn10eDUzZxki2yqr9cgUTsIcsUScMQNGhBXJuvu
f8i+/UIvqiYhGKWYr/cf47+KANDyk0AVuPtiz0eEro1gkwnv9eb7Kl0u+b4c87uN
SF6Cib1Py8GHUIRheTJKU/oBEI0oMyXXsEWDpBEkX5FNflbH3T/LJ4Kon1oa4vni
U3FXJ4oSj56a9OGw1vSdIkTdjUHFpZ1KfQQcqvrS61W4Y7Zy/DJXJXgwL9XBUj4M
nCVbkDUAsLkMN4x5sNjxdTbIZBRadtOXcPBh3VjS9Q34Spn3n4o9wILWFnDGUTi8
UT362igeqonP1BlY5B3K2YZbOv3ZLGqto7bXBzm7wZsEFQFB795F+5+XkHrLWU5P
qd58G4DrdL560CB06XeDHDnKVHWdfT5Tl5UjFWT39a2PAKVWLu172DEfJKJLm+CR
o1Q+K1cmP5/rUvUIdFpulvi7KW4JsWy8WBYrztXYg+G1k3ONpjMSNuArI2R3F+6S
Aos/CMtZnmDxwuLfeJnRUdlVqznRMa02rdRC5fkU3epTG/W4Om6qWpbW2cbIwHcP
STRumSGL8lgnSYYLB8SKjiNE5MaZhRzT7WxsVYzwRjAK6PCRS9WFRvm2eU/gPkoA
Q77CcGn+7DG95piMhWiqcEs5LkSTybZ4T2Ki/ik0CD1Qb+qxxa9VKgPnAJ10wo0v
dVn+qenwakBf48GVJGhKE7fWt312PmN0YG130MTnuE9Yj3IFib/YzffUzadoC2hk
8pa25NrqsPA69tF1zpRYeCPtSgQhpaJ0+5xOpO/E4sUIUa2Qmo1DPnnacB7e2ZYO
bUD5W5OHjRegfw0owGgUsLU8LkqH94UHL0nATqnrclaiTuz+NU5CygrQgMrbPPcg
yEjVlFKaLy1eagxlhJdZX/o2ZgHwi8wL+sZ+pkS44FuuYZ9CimU3awsu1U1e7aEW
MAZKNx9Cs8JBMeKLh/nedz1+EQMTVTM/xe6UdWUgfi8TlXPLyHK9qlXhVycY4Me9
Arrd1jX34KBS4kQUvWRC/AlsR0lLXJf8S0tAyyhtl52WVvtEQzzqXEckZ4tFvJlN
sJ1GgUqziRnKgZ2tzm89vDwEnps8FkUmlsfoyWy+ZQJAsUpJW31Pq4jp1WNzPCW6
h3lfMlDPr6SInMgLS7Vw24+Ewkt6NpPneALbVKy4XppgV+FQaMasH82FyNLTm8Lw
/vJV/yILw5cUv+baqv7Qs4rVq0zwi3mA36Yem+HFVY9BeB66waUnVKbcgvvWEzVV
egdANEh8LFPZTpOhHupX5UhJpbCxmpfZ4+XwFfHs8CVr+HeKIv32Qdj8jv1V2OnH
sXZxhf9roodu4M79QvQFG2jNLaDcaeN/gtmhg9De3Jh7+R4F7ETqqNzgt2Z7hBmm
C8O0RyfsBahawrFk9soAtOgss3UsEVssWY2AAuKF1h0QVxuuq6IyvMnruHkASHlt
3FLk+uWSe9FwzeMqyBjfQv/tMpArJUzNuxblqoT3JQalp0UNaUhqWnoUCoZMBneY
dRmC2a7hwBTzHE18m6Y2Lv4M7tz5TDAhUr6mqQ/RvxRhmGgy9SaY+l1Mt053hDzG
fI9Q72e29UXO8ImMcYX7/8KjFHDyb6VuVkrwXJVTaTMHmGUYpMs7hCchAB0RIbMz
Y/wtw7G/uaGOz1Ri6npycDZPz8FRLu6lEHkwV/6AMFsTAowPT866OL/fw17OOTz5
W6KZOYECtefrskRYt0m6qujWkPwspJm0jyTOWD8SPPj0ubRRNt5JDaWf0ZCsrXjO
NjmzV00H5mt+paEwkqcz73i/AAZhXkedvZkkpN5JY+RnSC21fhgaTQ9xOwPzX+V6
Y587XYzUzp9cMvxppzvEQd6J54z2g4yOyqaskf6NFlWszOwjyn1bxUV/31447VQo
AsfvZbg58g+8+f+y2V97FRtD6FDMEUBHGVsk8I11AO/n+M1sOBmzaMhTg36o2DnA
87Sv+RDay93bQis2+0NsjizsNDvi8DgyF4cInuaO3AuPOUWuw+yNYGPjIZcyCAVm
anv3zSK49IWYOTPdB8cDDUKC+c/HX5V3LCAQuPLJIHTfGNLp6yNbCOiMUmYorb3L
dJ03B2koZOKXa9bGxLKl9zX2L65/n02N81L+lHUeE5rYWVP+NAqzX+7g/du3Rpm4
Eq8gsn+T3YtSJN5UEfzPMWEX0CJzd2Ex/uNHxg76dGj4BENIcDBP60fD9TkluaSc
j14SPNrwnUwGwgIpcc1tXoMtZLP/B9gkTisNyvnJ8La9LwkNpmKH9NyXyaXgrYRd
V2zd0YAJwH3b8RRC+W7BBfRmM30zqYrVM+u6M7iRg0BU9nB2zgCqygnu2wDU4/15
KD3W0XB1oMkHCvi0LCe7bazDr0zxcmjJZ+643htOGEriwIW+c9RPPHRv/Yz0Hj8x
cUesDh4XB+Kdz6+THR2bPxXluI8C+8DDFhI3HekF8kjmdbKgSpntw7WYyFb6/R7u
nKKSRAPRKWnlfLYy68rL2ITkjL/Uj4+RggWjYo17RbxW0MmkiFS9FGnnVC3tjL1U
zzVUmqlHUAbWnaqQFlsTBDYKD84GYu0/k/DZqy6oAVxT0iUFn4F29IUe4m1Iymh/
z7VDnqM2wMVSzAul/nRtQd1uPMLMYqy7nr+/QuILJpq3zQml/obDlMWpdem5vxqy
moyXtOfdSf6bFtB+BRmhxFvw8XsDM+EdaX+OhD8js6jNmevEYdOpcOBwVB6PLmsk
cY3KeYoQ3FeDJtz3La8mq4xmELzrwDx/47dxWKmJS4qgapJq2tjuax3hYFYaj4kW
kR1EbYF4cT8AdfaYDQfF+TBDLMscVyAkwBoEMpGLrZIbLIUaFuXTcBSOsNj7M8iA
BfFoZj0AZgbTWCtzPnHNindzVMqfczEWasHCz9cSK6fGfMmbCIurEl6biofrQDPe
RuxhSzrgTEseQfmtqzQTqWHqIcXPgU93oksLCMw/aotAu72T9eOVJhmhWr9m6rSA
ymxKUyff/OfuOEepwTTV825HDJlV8OiPZo2F6PtRWoaYptEEL5M3mHh8SiTYK7pc
lQKM+yROysiBHwRZjokJkh4So+yWPgtbqVYszCSIdg1rMeOcD8ZQqDqwB0fpWORQ
9uKdrUMvzTEfY6u8miitNOPR6qN51vSMiAGGRS8f4DqewdURc+p0Npp8GkaA+VhF
nW+jLi4GF/DNtmvmATEVM8A9imt1vy4u/dt59BPDZsxeHRgOra21EOJB+I9cb1PR
pFnIZnfFAm/ckeqYWdA0ZECU54Fl6l5EYgLo5ehWIpKprDo75zHI0a+xfj9P//rA
SbyTu1C9zQFXOjc0e9HafgZmvowEwk1bRg8nXBfLZ+3wfnubJZowoNHgXfVcii6a
wKyLg8aqzFBDBOLeDYGTUWW46ogMHIEL9Glut0A/4d1ZtVQ7ERYPg7OcMNhIKqsk
jhZJlflUgNkcU6jYqj04oDYnWSI9KqBg+05W1L4dnMkMZ/LVDArreW/1HtG+Kwbv
jc1FOAtQ7KJrepjOA/uJ5ZDXZw/s+cYv5WUeM8NFiRYmb3TomNRoYyKV5JeXvbH8
G0PJaSg2hKZqM9+BqWcyruN4St+QDX5k6tnOZU3103zFdZLbcvDpeZ3t2nI/rgKh
plDs8eHoZy2s3bCLRdzZ7nLXu8oI77bAbBwVdxHyPSo6AoeaGUfx1E/r/G/ObcWJ
i5m9qO5Vap+xMIem58NybRcxsRni8aWxM4zGAbBJcexgx7pNgP6OqcJHSclafkvJ
iXWEvRqUQDrHed3FlGzP2jw8nLwVloQyA+2pT3MEM8fLRHdWdzeUC3U0DsrhizZu
ef5TD9hsH1t5OG/UK5z2Ujfqzh35E8xqqHSc+pR09kSGS8r6zSzznK/9ldq8itGj
30GRDKiIrzYKdq2Gy+hKo1ShdtCCbauNwvAwhMBLl1Ely40u1OIlFFNW69uBggIR
NqKCU4zvL964goB1kr/RC9vuznoFYinM268RselZ71kRzEBRIqW6MDon30xCfIis
FnBFpMOIrf+FlZBMwoKpew1lJS/bctzYD/Ge5YTEi/vKt2Y2cZ/hCgB+crCCjCXb
y0Iy5YTrLhMnPnfJkRl/+5xVtEDEqa393NG4CbU1vHSW2UMg6+jg0LmcA623V5xk
wx8Ddpfm7fUemREOETze7dLn/XN+kYT9bHX5JMj3CsfWaXc2sb0Ohae1E+VhJWsM
abmdWpO+BsCQGvdnePvnX9BqNRUG1LWtmO58Lc4zJpksCVaxzha1D4dxdYX79Bgx
2rbtk4UQYuaJ9sYpCVg3BqSUEWwru4uwsuRwv2mU3cTyKjOUEE+ezneITH/l05X0
bDbEgMrhgn13lzqy5rbrKNYUxUhpQPy2WkyC+MdDvdKFWNsgTElVHb+YfrBoS/ym
wkE513aQWRPUQsjt1aCobGgVzUgdp7fKO8EXb4hrRt5CMEI0+tPkQrfW89VQjAh+
jic6efBIRsZjHWQeDXiTEAWJLnMU/ZSpYzb6oOH0DXaqWyEIO6JmD53QR+3pSMs7
LUdX5hX6gzhDPIdWbadpZVG4OONPZMayaDBvQACOS7hBlLR/9L3J/xVOfqHKCpn7
MmTzhK87OCljz2NoiMPztV2jknSHW4HO5n7gtWe6LtXEaCxkbUSWe7qFGCPkCsYp
LbIe80TEQiaQbyqwWRcqJiAypz3NjSArGK5JHpuMq3T6k5M8zMEJINXQLqtXX05T
DSKP78lzeXxETg9YzJ6PKLDMzkDseMpkQOcDbgmz52cmUSVTNrfcUyP7bww4biES
7h4xwe/at+LyDWF83711NcmJFfIKzrctPdHhsEJpOm52Hs0jPmLzQOb6FTCgfO5D
YYtgDJuUu6dvKDYxZ0xJZx3yrorOiGP7C5/92IradszGe0A7F/+EqYRZALIgEGT9
EF1FZTyKL2hYnWQUoajZrXkZ3EBhV79S72fyLtzZbDWuAXxyP6IS4kp6VVmL+HQu
i5IL0ut5WekEkpJDHsiKn71sP4LXReSyWOCIT6aAWSI/n3mTlLJBtCWGbJV5hNN5
a3Nb4pfse73WesyxEl/bsAzNy6rvDStTLYOnKnXrCZInp0Z/RKdK9Yr4cDvXdR5M
AUdj86Ald9WuNDwW+0qP+7HCzBlf4tMfIyVWg5YQsFUlNnLoVGmLRkgpZoHjVX9q
U6+4u3phDe1wzTFykso1pCgwLmagffLTnEog8kkpxnYlvwRfG9bO9ri292w8TGtJ
cKqMufF83FJAGffcTjLqZa1/K079RvzUStlxQAakPjqVJevK99eZMXmvOqB5FIFz
1LcVrfCg5jJPRD8qTfisy/npqvcjcqgDkFZ5+FqVHTAlDyX32WbVReEMIOISEKCK
2WxPqQqCY2nnQqCbMrf+K/Q6eW12v+VX/RPDRaD5I03jJw45MNfrDjWU2r90bejK
DwWoQ8JqlXJh835GTebzf62oCCCsUXz0ifL13UPNl4cGaasutJQga1gELhnytnqG
fSfzwsG/IwDTEZqkRs3n3WUVLQXlpjtfJ4oArHVhnWS88CJWzro92LMoxg8Xk7Vj
AeIyhx2ItN7N+8nH0eXbVG32y8rLw7EhdgeLuNHZ3jtCzY3V3h8jPX6UG+ATkTjy
FjNqwLES4dW7PD1Ns6R0L+3goXVTW60RerDVucEywvcnP/w5sgeenmgdOwPj2LSG
heOnuT03NhysLq8vqlMjOromGgTNsg2Vv0XAsrsjNJC4zvCVJDq2zPV8ha88DaWG
P3NDw5wtwgdhBbO9U/h3ekBDjSOEAihcqQjJnszV2mlHPy2pphGpW72mxSn1tjoY
t2E+0ci7x2ACuwpw8o/+AUHxryXU4HxGur+L2wuUJfPsmHDG6NdMQKpb4f3HrTQg
WP1byxmWN0xk8KMlcUSt8J5aDmb5UjdH/cEpUNq3zFM7tLRmXQLg1HUW7in6Aogo
0cT2AdLvEgr1xwIqqvOCRxyicTSeN5+4vT7TZjDrfA52lWU5IWRNL8ghcRPLUUT4
CY8iPLuBjkme2SEfXT5s0PXEQd2ShCOToCjlzEN1fN3Q+G1doEZwyvYBd+HuDWja
In95/vcRLeQa1F5SuUG5TIFKunU77yz0FvgJRojUAB5KZFGEDC6e0mv+n78kK9xF
tRmxwswYyICriibp8wu4iBNmpWf25QFCXwXIU3UIsAw3t3XBK9bmToE1Om1WPegt
Lxry4ogW6N7qIMAXuwAsQD7rvaplBrnLWZecyuhe2CT4rSa8c+qfZunK36nGEDi+
PAIMmZ9ZIkwkW/bi9wvS7cVeYqDDY+zrU1YS+1EVOn8dAVV4Wiqo2hzJnwXJw2pP
9zL2DrB6oEiW8HG/XodiLfzFTdaSnLapdjue6ooK9VcbzcJLHHC6tXSBD0GiNWNh
c+esfpOafW/IMGC9Ls50LIxDrwQqjA3DDd3kx54A05yd7eUonWcjexJFEsDMh+iJ
0YUIkOFrmBeMYUthWxmuDhKkKRFwJ1uAr2BHEZabFrVsp4b13zkqtYn/oPbH4nlx
lEq6jf88cGhIPpuFKQ/1VwDf/8bwa5OIKrn5/3PJh+WWCfDq+jGDeBvKYgMEYDWc
mCBW2gN2104kSqN67dTUMOWbWm+8zYXuiSdcF0PNMvpRT5y04i3CuaAsiKZcIlKe
wDqMjQz4Ejr+qfjHEh5adA9nwNNyFQ2ZaTh1uo10h7mjhKtzbhmE5ymzhphgjUig
2WC06+BKCRg7w+uOxBl85ekcjVUR9SnoiikJ9JjlPflhaVSkjj3xvOIBca+WQUpS
+JGb4p1nNVacICbUDXWIEYZl8C9Zq5HQNfhWK3qN2QjQ2nSovw9dy6SBQKgLFNkF
78Cn2ZDQBrIkvKP4BPOTQk3lswJlBL5z5UwasGtNo/N4C2RbGYERliPb0e1Q2UyG
23JpdKOKXeaVJsIOl/O9YwNt4SQKbBDEsolslxOnFfdYnYk4dpM8QG9FfTj0TVpK
M3uuzbym3TAViDpmDM2iBAUHqd99Lqjx4AJ8tiP6rmI+hCuU0PbIWAsCBtV/rq+h
aJz/nDu9qKqKiJNm+XJEFQofam2gmkCkw0ErbUu9UsGcKU16FZbq29b+1W0HFVWd
fjCmij/hOgVGSynbOxXtiVKkeYIhA/bBK0aNP9UzH4DLvR6I6d/7LtCHIR5SNhBm
iEjAQf0YuhVhSAtkqYxPjbudNFEW13Wq/iO+y1efJedI9rwbaRxq0vblc5T5NZ9a
6FcLx7PKZc36DUJc+W8ueQIzyUiar2502V6BTctBEWrWh6keAcfUMPuBNQZ3y2HB
EXV9uEIufPd5xtnEYkHPhJXWe1yR4YFX6aN+YITbhSGgncor9elLMnhws2vEr/WP
CPbIrnlAF5k99ho7C2TjC4Ihecpx12uOiuz2xv0J7RL1ZenjCbAAAUBbBbt+HP0k
g4HtR4KxQfJOI9spr3JFVUNJUz7C6eATeJq2yz6wCgxKmlDCvHCJJrQJGQhUKPdf
i3Ub6taZW/jTg9jdO3KZsRuca0xactDzU6WfB9kAAIqGzffk2agAUvWZ/uYFJquH
oK8iP7iBbLehgigGnQlZpRiDBeGMQna39KegvPhNih0J34+Jk9SERe0bRVtSLkIm
UN8ssfIzHv5KDnDPzkkIRaQUF01S1XFu95sixhOs+ymWvJ9TovmWNlDRvrsY4wKA
c/MSqtYcUExVIMhtfQ5H7t8jJcK89vhz6JZXslCXIAwn2j1CSyAZRVXeomtClUjc
lw33LcTQTxGw3RO1b3C1gMaOWD2OWCkiNaLhwpfsutQjCZOwaRBCP3mqTprF+QKp
O6tIDf0q6UcAdBHagROIKJOywezjT4jMERVnVpWQmth097D3pG/dVzJmWNTlH/tY
ohf8wAIjgThgND/kF8L9J8Jjb3b1tSo5PnSMWnI+XM45dthvHJbRvQNtaCVtclm3
G1+dZh+8bAgy4oYgiVsxu6DkFJuNCASzz+CFcUxNn9kAvEoYbFqmBlzPSxHakx7B
lTxzPTtQJ4Jl6p7zUZAKXjI4NwL40jG+4E2xbchqa97HjiWO549qbYn5f9ustZyr
YeWOqwJpuL7EVW94B4nZqm4khuyIzBmuGJp5OIt4TlE6ZIfz86qprKt44IbkPspj
/b3NX2EA54bgJLQpZWm8+OBtwFO275jzEZJeCDyui95a/76tYs9yefiN8CT56kUX
lNxjiIgccxdA9ijxXIV13kvfBV5LImngivsk88LggrPkwFgv/SG4UkDl47jc2z1Z
hXKen5mHbwmcHXnWMzKpZR/DpPbnQPpxBmSMdlMTyk+NlI3Ys6qaOQ2BfRbcFzct
Bhs6QQSNdXZYhpu5RItpsy1LprOVBWhc4sXHJBTweo5G+yoTLnhpGc2oua/9jSRA
iWqZsvD7d81BCjTHbSsP5ayq2VrzCMRWErv1nynAUtlSfPMcNk3eYyIAdxP/Oqwo
LYUtUu2HwkfGrIhJt7faQU/d54tw59FIaT1YfLtyXniWtyMNXdCHiXQ293HON+qJ
JHIevHqTJG5ZrJgQS7SJq7FaTcZlhfaf2LLsAxCZEVPSIef+5ZakoBB64IvvyUgo
LLq6KjDiP5ZmWWINQ7pw23N3wzB6BISEleCiJpm6d9jrdMe5PRps2J4Kt9MF4SY4
JHcIGkSCMWLP9fVbyoCcGqrOk0HIWB/i8uny6f7MACJBXKxCbyfaYHCS3zX2+tz+
Gbv6V3lA8mQVHXBQVNE1N1/S6gknfnb+FD6yxngn7Ig6JF0VGp3dK0VTUxmGpG5q
if81QpLUCdjNZ82mwUhBxZPIHwZOFR21mu0Rcsco52aRrWxqCoyF6A5b1Be+sz2h
E6jLvIyrjvRbk+yMQgmKE7ZSaYlaY0UB2Q5ShVKPIHvRUYvjvov90828Wlx7cCYa
XcddrHRkzuNAxYQDyc+mZHqeU2jjqJwZj7ezFKSEySN62C5JUKRmCN7nJe8di6y2
dEiX/tLxMIcBl5+AdrEJWTUy+ygTEouHyxtRNVEbaOYJDpf6Fw46dLq90NFXeAlw
RV+pgokocn9t+xyQ87ZQXyCmKA+grdmokACFUqdlyKpy27Gg2eHePkBXFnsU8urm
owjI+U5Z7LyUrBOfoSnW+5IFAnADSOYRRD6z2RHTizOX5YSve+b4bgmvhVYOc6EN
GgLcLID/ub16sQayS+S+AogQTmUq2v1IgCPLFECmCfey/6f9A+bFGKG7rEkalRpv
iHNYvEm+AZ4fzlR3GSumJaShJjOj6BudGYaCDWR5WPW0HzyuNRv4lx4blJH3Y5W2
WsSwLeQW8i6X0catlfAKcghj+snYGheuguXXrWis7Z5Yuw9aFfLo05CwpjdCLi4s
ZUar1t1zojhY5O1VInTa2tzaQYbzhNWAHNZ45vcFDt9/K4qXrUXFou2mzuauR8Th
MBRfYJT8jqkbZ8YrCD2up6ZReGfdCjfBdoJ47jxU9qPZUVEJYkbwegsO+YoY9GCQ
olz8RmU2gF9t0JtKvpcd33+Ys4Fqt7o8dc8eesRiPC06aB2cFEbfPrzV7ssv8oRQ
oDP4lYX9C2rFnjPJ7d+d1lLGj6kT2VAzYEmoAMYOIvB38plQw3BTmmXncWPtGvHU
RBbTCSE5mRvK0CS4+Xt1hEMqeYPxcXyRucf05eP00SXlFvHl08ydxrXAuWeZcpOo
0oIpcXz6y2u9kX1ztdrl28okNaJvmGeH3RFwx8FHn7SoKKbySV99jo6SXZv8G5MC
jg5RgFAy5aousWRBvDse12pdeChwTuPkH77czZ1WQBVMwg5GWukZ9puWe5bG8AmB
/6aVd5dZPK0KSMYhyMZHdxQZtUDu14qMiUcO/VOQMiVqBFFyG4MtgG5hnVaTAP2o
QmXMU5c1sYvjHsdEYTCB+4FocHDlFoh4hIpgzcuUJJb+0Y7ML5BGjD3VeF+zTXUB
Mc9eaniVNe6bQJbSNXwLJk6AsDmGIN/eHoLonkWwLB5jwcu7egzrBGq9SHTUeenz
W6/QbaNMwSk9cbFGJD2Iis0KX/34+VjJez8Qq2NAiNJrwcSdpWRLAwx01F+do6KH
rnWjxkLKwTOEVbruWvvEU4sFp3iepi2mNYOSJW20xfVi50sEyp+Nl0gmNbkcy4p2
6s0GnbEeF/RK1b0TbS8wWw6c+Glr0KkY6hc2wgSkmt5TfJdSWIXUhqHs1K2GRLTO
hxQWoDh9z2/5jl+43tu8+d4cECAoAv85eSbKSQZQMBbbw8V4gITgK//puSADONop
fHRI4i3JmLUKRc3yoENl6i3xg8woN4/aJzxKzbP+KLuVGS0QM+8X6eouqqHc8Ilr
uNtkFoW6I81qXFSVIPvxbn5A4xSqTt+ZVdrauP+y3GKpmAvbA3Z6+BohLVOm1402
LvheYD/vj9k6R27lWUqPL1AL4CTuo0Rxs/A72u2nq+TOPhqQglBB4coW1Rub4W3P
Cnfz56Rg1xja4hkRYT1a+pbXuKBwgL2g9SR42X0AGGmfzHMCOX/WXsoU0Au/9vTD
bl3hLeEro0Zj+lv/OWdoHRh5GkkfNYFYsHUKByyh2Yu51U45tOBuZPhE9VTPkY5M
p8b5M2auTo5/dDVN8Z3ia2GvXrVTjwy4FjENkfvcU4Qo2HTxnGBx+iGUxQ/2viIF
aq5GTbZ666xZTtSucQdD0DCAmlRoPasW7W2hGf9JiCA5+jm7r1znp/Mc5Kkvzg6e
ObiAZVwBTytADi95G8WjOMzrU2GV5Jbf2/7i0waR/TZljU4K7ZTTX+uYyDFdaCAY
9PW+kqEMLJt2ZltamWgL0dhDlmsx0FF19Si6BRcl9WZ9Kdk9DOxDy87JRZBEOp7B
ihgczCNy3t81AJqBTyQBRi3cbPMgW8tR6E2jtcU5l3R/OEMO9OEQkz1vfn4jYr8e
FWxO0poaFFIyORwDDi+9rcPHVMZ+dNBl192wh7h8g2p73gFgPybsnvqQp0NszgwT
DAmejIJ7Y4u7c4ZNx2Fk9/QvxtD4z6PGkHrnIX22k8j0aj02l8mbxkfB4ChppGsu
v6szBBwG0qI/XF4W7+vpDyYiwr2Cqok8SyklIsbNAjNuTPilWzOHqMbbokSg6E1N
ZKR77IslsGhI/8Hgmk4wcSO6j00Jieg021F2pJgXEmKkZyHrE+RodB+SYxPTJx0/
mOx/0f6XCL/X4F2Dgw1vFtt8d2RTz7qGAhLwpctNR2f6qrfS2/G99zdVUtUPYO3n
Go+7ZwVokP5k8U9NReeOWXK83Zu+94w/xlvSOBqDghTZs/nnfBspXmAhhlPuwPFm
UW18YsQQGVt8YywvHccAEQotQnAXS96mCHjyBCnav8oV03O77X0HoblXZwspOXn1
eJczrpeh9gVbVNxhuVzFGnAMgyHyE/CPfU2/vRDsd5ryv+w1dwHVhN3q5I0cpydc
vEyOYHnkcRtU05Kmnhcd4IjJmKKX4cp0X0EQVFCiBi2mo6j/er88UFb2Oz8hfihK
6Es/1JI8L7Eo9BkVFPySTCt25ajJMtN9DiTwRY1W9iKr1xRMBstz407Tgcy0VZlC
HAARHtvVERw+9ldlbh8+1DfR8Bh7kS3oBFn/Nbrdk/iiWawoDhQes7cEbUWc490P
L63vG1WD99txw/nJop/GKofBem2kJ2WzyHmqBZF3EKZ8nrcZPXFwxRAtXEvaJvTz
whvlVL/EnZHr0tSoXckfuP8MUfsfkNbP/rwkoUOgXK2K0S4JXZGn/DfSpiq4KI2V
u0VouT1VXNwCaqczERzTG+3DviNIAaOzTYpFsYj7opDKgDdGK+h3X9fCESIHWK7u
GZO6sqc1qNHlxKL24LjBPcr6q0sXS7rkl/VnkIkUG5h2h10FHGW4OAoa9i1k8Es2
evSZ9/M3qH2NeHQGyWrk1nWYvdW8FIYDfGEKEtpHNwRLE7AEFE8/SZDobAfrjVS8
hw8mXX1FCBNZGPzT1Enq1lOLX4XxbvayspYbXTkbL0+WrCSSwQxe0fngS+tZrgNX
LO6iNFtE3UffITA+yDNaLAHJcruN0/jl3KWy9AndENOv5siZX8tItzpuili1pSre
45tb3N6JNA8rV/31gzLeB/A+TJhYlUSv0z+0B88ArUpS9py+2ZBMUbuji1E4rqhL
04LD+6nyCn3ABk/YmreGT4Fm/t2u/yXT3ujo9l45BrIPP/lbTpP67odpFpPmcsns
zROkwp7OOJyZyZbG5GjpTRjmaNp+ZF7pOe50E/h1Ldzoi9fNPe4fdELPIYl3gEPN
pPAqjrmWWzro4mWjXWTFEEIfF2kiugzpHxtUzUPZAsXfXqbD++1bfio8cNsJRs2b
/VbEPdwRkQd3vMGWYnlKwghhGS2he/gOtF7pFv1xQk7YpfAKlB4bUhVHiqzQcOQd
/IiwbWlun16r+YuaC23SqiAoZJ0MZBut+UISy0u2ud0ZcrJ7KHtZLs//keJHacWX
4rUrG6DODvzwmAAn/eXsP8+SorqBNS0WVufRACM+TeNIPEvmjdsoCi6raUO4bsgi
okqcH/lTx36GQBNZrRxkh5RiA8T/fTiJrV9ECf56tvjX0iljz0afBUDWFmJUMMN8
/12Ut7vHDPkteNWejrLj8ve83Yuk52WGU+B1CoaurCVkE5HA9XQ+50zD3MvQNs1H
aOiRTMyTGZs4hJyz2SV+wXWvbJXx66ZL4FG+KYdVqU+TupxV4LGnNGWKti8EIG6s
d+ExP2dsGBFJPw0SD112HCiDLDTgi0L6QxqzParv1U1Khm5mIfJh0DGiwVY+ADnp
jdCAnYghkyjJohtEIR/spzdo5vF78ykewR46INgWI/aUhg5pMI8/k+T3Owt7RVJW
p6JImaAnmZAXYKiJ1WiZy3reNNS/9zpwMhjKmVhdguXU39TJJ82KiPWn9/Gu0M7Y
41i//Ibbuu7yHrzO475sNxYYDyukHwTrksVfMaaZEnCJZsKrrvq8fvT+Jbk+kCs4
g9IV88i0/3ccNBS1b+dwXsRdvpb8nlw7mRVtn+dbaEDK4dwkUhyyRsFfnNAyjGMW
4SEarXEntWFLWnFrUTexzB/FdHMLVqS/H9hyzuI+v8ilrpPmxbe3iH7p4YfEqvd7
5QgaAiItyyHTK7sCD2AqtrFqJcT9NHq+W9q888fk6pdMgxNZSZAhnIBU+Ur6QVYQ
5R+lSFzOzkXnbS4ZML+WzKkb6dLlqNJZIuQEBo1w28EC+avpbgrcR/+1rOu7a5OF
bZg0DghljZlNB88surB7hh+oUbWQhxy5rQ0Mh/ClGeEHLEs0Ja+nvWmq89P1WFWW
hnEhA/8h1CQa/6bHBwII/8LqwclDN735D2Kc68Rvcv0mkpuoGLvvlnX6QLPouyE6
x9frsF1GoQb/6J6/shYODQT1kZ6PpgK++aYAzuH/uDembQfn12+s9mZTp8IYqwtJ
MemD0d0/lFWPwCJ9ZIRLeNIWgSUPEFSb21u6ZuZmx4sLt8Z8LQop1p9LHdc2yAZu
Q7FSf8BZi4exnJNkR9MqSJuO/AA3ozsnPtgAWHCiUNM8f9eOLYwnFsePVFmHLyVr
Zr63y50Mwf6lWueagyV5IM9s5PFCfsNGejrxqc8ChWmUHmGSZEl/kig2DCaZsPmV
FYW63eixHEUjZkGaoeMDCBeJ5DonYJjFZ70Zr4uRzaAS9S33K7mfuNTzHe8qXsW1
xiPtrCWxyDL5Nhis21AFQid3UWj5JZFMfXKkAheIfzHSt5ph2qFlPu5u9rfhq+8j
4wEEcg+l//+NF8kIUaoxOK1y+C0dXcjlIy8eqoLe1kz3eXTa+ji0n6uCwpRIJ0KU
DgkV7dzy7N5evZE02JdFL+hXujjMqTpOC7WJFyks2yKWBfMnJiHFLsXS8T9f94RZ
cZ+Z9j9H3GRL4BxiiBcf8kWHUawOnLv5shJhfWHVNYQJQ/TRGLJicvl36d2Yk0fW
zuM2gP5egKKduk4CePTWGKd5kX85Ew0Ozu+7y+E/5CcRjV9D4tk2JQu9O0tVc4P5
hyz7VK1weKVpaaAScuLYYdqi8SdIRco3CLK6PBxo45sj0scFZp+H/aVzpqqaX694
tdNmOcHZ7UhYhbxEpsXYiwwz6QkDJQFy0xzOf2Fc929XL+kNUqcCpghiI0uHgNDn
dCNKmrsm/r7UB5/F5EpaIVqgYNM1VcpjIG2fjtCl47t5gQ+jZGxSKK0qNJkDd+to
PbK9gz1NONRzdUPcuYGK8AG+9nAuV/ZOZUzQJklw8K6jeZmvnM64AudEnvGxq16J
ZfGL+EHjGSqo8tuQnEoM1A/OAeD71/zB2hIMhm2XHSC2f6uRJEf1hKEt5KYp1vd3
WdRf846PPIH5Pv/Mi3DCKDIU98s9eWGhHNUnS97xexDiXSWdgPdK9kMm9se+Uie9
EkINU62NSpkxQL9DjeI+DCvybgMEUgZeb7+kEyiALb61xmd9FlbR/S+oQvjTG0W5
SRsKOiVnkZDhGjkIoeMSebc368DhNHH+e+AcQrNwt6oXXdb/ys9d9mApe8e80q/u
T8bjsMClsRmMa9DDI1KgwRX8fkw1dDT7Qynnb/rvHgkb+65jHxnl/khMpWlmfBi+
B2Ilwb6RKSEuF91EI6ilHB8y29pWaf8JqShkNglnIYq2tcyc5Lx+0qaSa1+HELkW
9jx8gmb8RqnLmqMjExiR0netPqm0DbcnFjyO+d7BFWycPUqjnno+dar20CpgXDXq
lT30SqzVpv3Ab/Po4xCO1S1+c4QKqes3RwqP0C41bOw5Tl9kgeW0P0WnCGBm9wnc
O4wi2PTRP0IK9a/eAnbgSnrHzZZrehozAN8bLfth/pvBNV9PERGYpU1h0JFNUlXX
ztiHutWYuODn8sXuc2abX6NSAXH8U5sHt2iPcJ75lQqBKV5s0/MMtncVX+26+gVE
uxT4NOaVVHWuayvGDGfez/F2ZrNpruxQ8LN59fmkuXOH1qhJuo2MTNLLJ7NxsG4B
ZCbhj3XTFaxRZ9DsQ+WBrc97rmuNF74/4r8oAEz5Oy78Q1eClw15Cb6306A3SQy7
tKNoCwj9e4QzMsUOoKjVVE+NqRWyGXDaIx4DbDXb+AU9b+nqDENmXFueMUsdCw9r
2C0wpkRLXrCN7SAEodFyNkIAE7oZtP3DnReEUGCtm21kgiuvUurfOWN5XlcCyvnb
C4w42s/VS4O9mgyarK2R4KRk5bXO0Vt0h5OlxeonPw0ohU0tDTalUWROmJBuDIP7
3CFvzfIKgcZKRRaquZfvHzsWAGvXcq5oeEPbmXubwF1ZxdSZCSQCULEJIueeKQ8d
K45/CjNTozt6lVoIDH0A9uTzJlobnlwLKgzTQAA0nl+lXYPI9rC2t/jPeCu/eSAG
0zmruOPtwRxPdr7kIjcmTG35WjmMqFTfGejKjAbeHFubYXAQ9VtulQBdMUnSMcep
rq0cng2JlI0/BBo4QLl1kiFnlTHiUJmJS0EtinBI4AYFrQFqi3jIrj2G3mWK5elA
anaitV8BbXqsxUkdJhMnc55ECvsp5HN928KasQJBko2i2Y+CgPZeDYvrdhIgm19o
6xzJG9K8pg9sUyaJHAe/tIos947nNfxqx4aJ0t5trQzJ9WB1agQbsa12PxlSldTw
yQxfplCiLNUI+DZYhwabu/jsPnYScOUUjAvyhsJiY69VQxvhj7s3rZ5DrUrxuIpk
iP3Iydk8xDIk3CQSEjOEJN3Qp6gRHlAj6UdVzuic9r+R1wsUtdZ2rkPSQUra/TKA
ugL2rutp78O9i9qK+IYQleqKxMPjJKGWvD8CY6Gwzww5wI9RnQjKTTRYvcoW5XFn
Vh+VUpqDz0HARGTf/dZda+8gnrDr5sGWqyOJ0E+BxxGNYCMLoZKfUfPhIdoLC1rL
WEpfdt1lpBMLB5btt+iHime3t2z+psH8KvinCRCP+BdC43QrYfH1Ph5TYp/8qV3B
QDgYLF58XIs8fJDwIdaSGA4scVhg9uRdawRv875/x+EZYePs+BHWSUkktIxaUFHU
PiuzIGfIEh+SADbknrGFWSUUD8UmSEtUWzIlBs5ACabQuSM61ItV3Lvues9fGrVC
16fF7ngEiT3AdjXUwSkYYY54YGd1Ti/RzwgAnaCdE+Q/WpKgvnenyjAEI0nbWWoW
3Dh24pFpsIuDpQxqaFWd735cQeNzDbGOswR3ZSI7wvxiJAGaD57D3YeeauitgpxC
r01LehDTJhd7G0jTU6tQ7vc6sJIHxrUZyT1dZpmlEGTpfZ4GpObKKC+vAubPlyzx
e32dAbqSaplX+gDJ5+jznacI+H4GE2kClNBIgFkCBSxeMz4vRmIVchCHhopvsges
tQPFg9ZfK2gNk8q9C6+xbLsTHcWzHoCBJ6hpkSqF4DaOXl1zgNLMZvfWrOzfGrTi
vTu8wOS8jeNFF58897TCOqSV9rVb6YR7qHzb1qBD+ZxuZG6ZVt8gKgG2YP5Kg42v
DMmCSCK0dYRAvjmZtzrIzLwdBnW4vIILCKWNRW9SYj2aAAI1yvbVk3yfwtBNJT6q
wzaUvPP8rElPIYptuMcbflvM+j59EKrlVUpiIeYyBYBfTA4pv2CP9FXcXh6vnaxA
2Vj1yUN0WtO1QAFD5pHafGxe24SCbQKhebB7BK1aA8LeiH3kSk7kqpQz8/MUQNpp
3gLTM1DRi33qiQ8e4JOwhnYlKijQLecqcV3Zq0k6xdO3KZlJmD7y6X2StW8Tqwz4
i4a+wQIua6+m5xV0lad9XfidsZC91dxkJPBp1MGGdYSSJKBk2sSIizEbpRDzBEGO
7AjPWcaCIc1Ql4xDgyBql7LubRjqw5jWZrksPoztdd/24Pv8U4Nzj2ap4vBdpKNH
SwkWudinl084U2OPJ6NVwapon7UTRQ6A5qkeuEo48x7DB5ssvjwCI+RK5hYiTAF2
WJxFrSIZo8WwTXnQAbijienakDW1I16N0AX88ZlbEqkUS9AC4go5H4zRqpTKxEgd
C137ntnbLvJmYv4Q4kB73znmVF1hX+kHgBxSf852sWXstCNBVw+hymT0VHeRnWlL
Q4Q5y8MXb8zpz98uuRXVPFywhkVd/VB4iBIOyqlGLgIPqADUfDvkKtHh95hIZKXE
F156d65dPRmyFtrUXiQ+keDPJb2jkF8ifHxeRir5pNzQaTIV5X1Ji4+zDRwa2GVh
vvfNUphfLNcl9kXmWI/+YcJoHE1kK9ZR+BLRlb1TzBrwDpmFN5D3jXk1o9QI9D8g
S1cweQ0eeFn/y4/Hk5avDjK55JBxC3gzoX/GE9XAfPkMkRNgX2W1gveDfrKFZhNV
+bC1LMuOUd1yR4uZ4ZvtCY4KPKH/mjpCxYttfjaRqJ0bi8dZJ5Bc+AixV9pvYfGz
OJx/vlBd4DgIADCbTMU8V39pVUjSARA3eB/UC2NKEYlnaLyxcXPl7zQ5Xtq6ZX+C
p5IxZK6eI3wIU4cKNSQ3HoopklRGb0edBq3LJOhB2RBh/pfq3arGbSRFRlcuFldc
Qa2Eg4wVi9jYYaLzqEP1hlQtfSqOPx+Y6NBfEpiP1qePySMJ/1JStlMojGSHAyTW
TdQkfcVFUDiiKwlXwP5Y3bnSM0THecktePVNoxWalp/suuXa3NgV96u7s4JmhoDm
I9f7AkpjeuhlGSi9EW5R1nRNAE1LNe/RNGO12FNmaHVhD9+P8iXiqsroOra0rAkn
8Iv5iuimuWQkekfGcADQsiVMrOnezHBdYz4212jxDp2whvprrhETsuyr/w1gux1w
GvOFPww7iDidz0E9Ax6b/p1tix/ebGes5dIQf98Bs0p8QG7NS8FR0jUBAy0HQ4FK
w3it8kRca9JuwDSyLrgE4mtkAum41OvkJJj+Sdy/q2lTGnuJyAKZNpEDjQ7uKIMU
S72/6HazyTv0tu81ZRzXk8VYTFm8JECcs/LeApzEFDJqIZ8IO/B9Ld/Uh0VI3v5p
0pA7RAnDI5/fiVNGsEFHSmbtW417yGySS7wA/2GyCGC4TbHfFJm3MQxSIY9vRruS
ZPrR6MkfiqBdfiBsAKDwJUTDSN2lIKEAuAFXl9YnNUmO8bkivF2+oN/1e06CZSaN
4YpfiZIOV5mGU1JwQtqHMPDKpYukr/x4g3RVIMYtlBgAzYBrnOcws5gIZUCF1HUU
ruy0RtIv98mCYckd46OXhsw3Ki2KNCzin/EKBDt9X0ttMBKFltaEjhVAdXdqBJJm
wXr84HRltiVgJUjuwgu0U9vNCxiunUzgBzLuFp3/PwOXlm2DDEoMLwZM2bbS2oDd
P3LdX0M/HfoN6ZOMeZOA/omDPqOhfKVd5ycki1UADqyQ92CpXj+K0a7PzsYkt/+3
uGJsqZpY6WHEWrq4cU58zfFx5HmFYD8J/AGH1CvgqaLnE8oOW0+T1QWn/UcR0v9p
4hHaDKraEu3yZxM/3Eepm0en6QvQhFP3Zg6UmwEcuyrbrYf7pZuIW3OFln3Xq0TF
YXq6Yg6oMgfIuCra2IsQLbGREo4qVecDRskJGXa/mV2/tWo628DkaxcLEG3BmE8A
HDLdmZ4LmUaNFs9Qi/NlmfHXmuopBYSq8nS2pPVSBeyxcTKlIgoPc+iN/oaJPu34
Md+ZHJOdY/X/47JMxv69PUMZrab4bDRRhYc5GSpZLBpd9UXsQvOxs3PD3Y/4jI15
9vl4ipKvQhyawdfqcHFJLchlSyP7HReLOj4SY44Dzh84eLNnLLP6ddyMWr8JCFxE
vryIU14/AguupLV1xdMctrnNLD8+DnsEej36BdbCuEh6aTP8XkDkS77kSyNHit2g
ZOoJDwBfuN1tURUWOGD7sE3l6T1AdI/4QODh2w7kpEm4KRiITeV/O+z+wsW+ZDem
ncFqn1bSv7pU/LbYrrBW1gj6nkneo0oNywW5z+QOkGifu0XPMha/tMBQ93cZeo6m
/eyKAqAnXs+MRVxRnGKvpQbsoBJbR4a2EfYQjEZYhj586KpeyJ9NRff1cy4fHvrc
upmpzAIZjZx5LBtwRgMykYdn58/H48BL0SlkMCNsYFza97LbJZM2S9FqkQeXogdm
Dh4lR5IzcsXGejvUyvHgsr3DxCC6lSV9pkKcErDFT0QvDxaKEIJE6sxMnApngUji
arWEfMjHtPgIKGMWro+XJBYXuUTAuR+45iVDetYa7jeAZDfnt/fREPJx0ZL8MxCU
VkWyjcIxuRNT2gA39LAcCmjTF49OMTZvK6rzUOXLrprOCpsyd4xnzc6rlMfizdl8
eLxLHOoiAETKda5KO+DPx5dkIINSe0iQL+dN0X2f4x81djw3PDL0mP4Cq+DsGiC2
nBPPddRhe9YIZomekY8RrPw/d9scWcEm/DFFEdxUztwfLh6b5O6qmfufUw/Ru7Rc
0o4Fr4j0ZBsiZhGGMqU2CNCJ7rFM0HoUTihlGvEludTzM1CmqwoVu1bZFWTqH2v2
6qp5wYIu/Pk6jRTQMIl5qdrNPss9lajUCOMFqvJ1ocT4vnp5ANy65964ECnBChMu
dgp1xePeAf8RWPlle9RQkE54DWvSmg6NPPlNuJNX5PtjWvwiyaLFXN/RwyM+MBHd
7NxZxXd0qXmQKo/A8c+98YxCr45bUcOY9msvvnJHXiYTWQvjaqe/+X3ZYZpm9a2V
+GnhFTzQprpBAoqbj9zyCvoJYBKUmJkjXFAwv/8m077wII6aEKhBsU66A8obKGl0
xWekjn5qkb/F3PSvclHnua50uFFQZdAIdwyySohdobSJEDvNU6nqUz4QD3kXqsqs
tf8794OxhD3WqCuz+GUFDodMGjgcZFeHhX5V848nfXwmbYGmXXo0v9IBmpYiVIRI
qodmdLX5rgvSPrI6nBsO0zTE9HspqXWw1Bh3kzE7m8iCf6ere3q6gutbr3uO7ej7
jSRjLNQUIf+lHHm5xKNFV/KqE+3FLaw2dyOTX1sd1js+CnfQCYD+pj5+/oCfgEz6
UDpgTQWmQoYHXQEZBnrUtGyVOwcIj5TloNklq0kTI/y0icLSm+ln+GLNJAZDnHy7
H04IS4Noq2OwPXkTYsXbhxU9/h2PGG73WhCXjYrR3af4LLQOmzRzCrBVkXbS934V
Ex961AetP/ejRU4xg2j3CkATaXEQoWMqe62/hPSWMH8KTstzhwmssmSkFrywFooW
Wzbk+sg2QWOHDxrK6+OgW72lOU91/CeXfBdaGSXlIJSg5OTX5dMpHHHfqmpba7ID
jYTBkMIiDjZTF3sDb/2gHy1Q7bxaV4wkdG1Hn1iMhv9oC5pCz93OKfsaBVnOLAaK
NeDiFeWX6Uu77ZTagEqEdOAwhptIti0U9z7j+u9tp4v6WkhTvsBhbrplLEkYcrIT
4QKYdbEXadraxzZEYZrGl2PjGvYQeqT3W1izy9QajLu3rixhJWmW6G6bgMFPNrIn
cRTnfgdpMzucm5EJpDG6s9nQN3suhkxzlcV3OSXd/V2EA0DxLqpYRtxHR9dNIFq1
x8XETY2v3Jumw0j7Jt7REpL+h+R/tKA3TpQGRbSuMpXkjkwwiyqqpqtNbMsQcsNa
IJVjIHSJBoIhYi3Tuhch+MoeUaktzxWS043NGus2FjlnOACbhpfn0DdGE4Nt/iDQ
lbY29FNOvVfGdsikccMC4jJ1YrpZbHC+oV/4y8KZQ4/N/45X4bYRrW59ktMRNyS5
yYo/4J5HZd3gnfrdX045JA/3StCfubYub6hY6JqK2Ub3fl9Ozdv0pS84O4k7OONC
Rjs+ylUjHX4XcFREN1cIGU2NrkoLoQmbCRbHMvSd5L7jaon9Ha3I8srXEFpF/BNB
LeW2fKNbw+rrSgM1RMaZ5lr42TplU+axELli0t4NrWreeoZMyQaRsKgB8R6+XOK0
I1xdLj8HwkocFVOhCTsdcbgLaIcyvQmczgvt1FNkgEbHuYfkXI6YnaEvQRRHnz4F
xDdi4rWTFmIqHHqvqfERNJyeeAFXHXikro9N6SFb8ctAcvN1csqxUEGISGFioq1P
cGZ+sAoUgJV8Ism9bev6ohR54c+zeFVjesKiSJirYerRqmbmHjsIgqnXP16G/QIk
JSvhG6oFALM2QcqqoT7wWo7L4y8Ah1ZrWe7NkgVRqKrocIHlHT11czsZRRKHyd+7
yMJVY5bSsrb/S8DcA5oe7Y+U+XlkVoCpJCbqyL9mLGzioIQSfCVYDxhQ45yDWw1X
DGkLtBe6gSaiHfgPYkrAym6V5jUaChSZw4XQbIxDIOvkJoTAT39yoC39CG07BjD5
rA+CupEvLD07yNypMXdsbov+54mzmncltJA2MP6N/8nSWRZyksp9KqhUK8yi/GMD
1xF8FEUNcUYEi9g8x0yjup5KKpcftG57yFvtsBJoAYRxtftDdq+Qh+yxF5H14J9L
l7uzCqHP/bJwIijAB0JZolObzsi65G0RY6HAzzFNOFzQbhcJKOkwXyG21Qup8ZsE
ahpk+borbdJMQAVlL8CyiToExubWcB/DyXMGpOYNa1bJ/KZKmIFMopzSolw8t1GR
9+lLsfre7r9HnUHSmVS+pGAwKrpqwvofiv6rF2+rrI8ntqb16ifWXvBYlSP7IR9a
TXz+DvXOVvycaRdtOvwrSl/tfWBnkp0qhaIVSNFam6pzZ0GFLbOtP80O9NRngTsq
4guklUsr7myXkSzQ1FDXDJhxoIty7/mMGbt4D4nwLLwTZoajUP3D0lGP8Ig2DeX0
Fvv9ns7sgHRiKcowktH3nhUY/eSzihkm2hgll+9yRMW8AKNYyMdIK9T/lHJu8lAu
DFvnH+ooTNvezWzIcJAc4KylN1/oJvvoYC2BMBQ6tm86Qyx56XMp41d99TKi9DRp
fn+AqV1fZQ8hM9C+qcKm+j2f259rpaltZHBxYf21Es8/2d56nrU3ffMd/aTgbQaF
oSUP/jx6y51pKwRizAMrK+VM/LWx3UNZnnOcMFs12F6sIyfjHRyLIi0d6EbAEGXu
OH2cFLR6rNJTNoLrtGEqo2q2t7J4TnEDenQG1Diu5TLxcCp62jjb4l70EfvP0QZ/
iR9Iv/qsSWoFjAe5jiTmSzQFL6l1Y1ondZkqIiHlHbxiFz+f5uPGviQYWto4Mnha
NdLU5+Z6TKmiQejFjfmacT4x2azM+lk/NIPebnt1PgaBHW3MrnfKGSZIdDjMkMmb
ZmO/9S5D6TxChOJKa0BPANehMvmK9FNqnvqJf5uLEgi4a3LwnjGJ5U7BL9qux7/S
C2M3QRJB0s1AKlMGMZ5885vCcBe4wXrhUANNCrOMpeEcMPSiFJ8yeKguFjzXaZrw
cLyqKfv/Md4PFBhIMsyxBxa9gZj7KqAfi7Fd3LioWXfrDKO2X6orZwHlHD2J7/5w
bda7QvRQSGwKQQQ4S70HmGSy3r0XfHjwfZDDEO37WpZ9HivQaPOQGAKsOLOtumYJ
xyJDE7EMzJ7StaCsfTBIOh9kn46MbX3cPdtrVu0qAheEhtbXxk246L8hfJECl8G3
vIG5IJR+qQGC+lGtbanfJC2wzwV6PXWhA3HfJOUgz2wmoHcvKzLjpcu6NGwaZEHh
6o72dhHSkUyi//b998eeLztZFSROupLuPlml88fSI0e7ZatETG2AdKy9X7hAmvf6
/YDXlMuc/X05iaIKEhExvbeG5opjh8RXrbLgn7zy8KSDL/wtutj2boBpO3t4gdIV
zA7I+65v0T9UNjp2e7efg/CszpqvZpcA9QdqSRkr/q6uHCr8VxDW8MV6YYFuSAiW
q6FIJQpIgoH9/jw8acLIXZcLIRtEoHC8zUpwZPmKWo1SDSPvFmo+QpdC3pldv1qq
utfF4opjCrPBK3nt4wHiU+if+eilJ5y5PO8JO4lN2vGG5uAvb4LVPxfPTd5NzErE
4IR3CIB7P3M+zFdwxS1jYSANKaaBXSDZbf6mDjXDzuqOdUsssFAK+ISxWbu9DaIJ
t5S4G52qlEkIub9dZyqHpzGg/rosFSO0MqNhu1zKaknj5AwkVb5W4Imb1/qqok85
pYpxDBqtGOlN1D1wVcBGMH/omi+13ihlQG/HCSwHDURjhoNsVur8vVSImICQaIDl
ezqZhGRVjAvTJLgCqVexSyfqoP0K6KpC3PQ/WGGUHp2QSsc1AmiJxKm04NiDKxOa
+JGZx4oMZdQvSLOx6DBAmx0OIohPuyzPNuguXrBJ/kVZm7BHoN9IcihUfZubAxE5
+HzAyYVb7wHSYXJX0Vp0Xt8Di6HTvKp/EpLU48Lo6EbZ/oSFdg5Np88g083XUfis
xVEZnmE3fRHlf9OJdN8w0fzy5vEMvUzD0aZPzPAWNAYcoy85UAz5KBtcaV/zb7bo
8vxYV3gYGcH8MrQiAtS/H+zJt7vRi3emcTF36vIXY1mgkoKJdKIAeU06DT4hda/P
Fyx+hVfJXwIbww/x0kHe305huMaL+MkbWCpUWgZb+N1Xac+Y5OUYa3ISTLvT+qzw
muoGVENK0sizNqD3oGYC8X+lSHKyeLez/Mec+3UIp5zXwCVoWYk5NXX6GfC+5PRJ
UFA05+4P0XjAy/SVLm+o2vTLHcNiYq+ZcIQBuDOVhZPMxPIE2R8whQslMSmuLBt2
/Fbu5uJAEmLyDgvHHDeHynjtG33/tjMOMVX9QzR9nzs9Eurh8ALBJ0WSsodKzlSz
ttgEh2vYGZCFZM2HzKJdrMuyFFkpc3breSN93IRGtWOdPgc3NUrdX9vTXPKZORA8
Iqdnp0gGl6LVHeQ+bhfUxq4AB+qTn3+HHqlUAjPS885Rt2JKV2j3IxGi1ey6z62j
AUA1XvazZtbVcKVToDBwyybJ4PTAwlMrgIVFTqOyIREZpvWkcmMlW1M/Uk/a+IeS
EPgQkVVdNTN2rgmpPt+jnucpovuqwyqYEUZmHiKJsBNyJ8mBvPk6iuYWdproQu55
KNtA5K4x/kLyuOAByQzTDZi0vOh/CQNMEDl+NpaLBDqBFjChfz6EN1V8nuqIzFVK
vdbZ4EfP7hJt2Sx3g+GODVKrQ7Wh29YynQnvtcaBIYQdNwjbiGuDXtgtq3lLGw+r
gqgF8wb2VRJ7kqNT4oJUmA1SJxKoeqg6I6brp+lby+2lV2h6Vm+Qhlvv4RseFLub
FMJKg93x97/6VKf6NEXoJCcgO9jviWE7Zb9rPq81EWZwdmOS+ZyqZGcxrYDoYssN
o/iGurThKldlsOjGwyzcbasoVExOvN8/GzKzi8wocN5630T/Gs7Ji1nYMHAwkB9p
PGzD5xTt6eAB7OU5FPL07rOKU/8Mq8XPpCnj3Gu6eQYM3if5P0tsAfgPpZDTXqGl
XQOIzx/5E0Yv93+EjON8t//YivOM2RAXFOO/UIZQpjrsTCnsTyLzHkRR9agDHNUT
9HXcI9JRDPyAoFfzgEwulhp2vnhkWES8cQQqWlggYu5r9/j5aneAY98GagVmTgav
olurNik3SnxQpT/b0dCfVGdXtAf2mM9f6VwwXznFDD/30p2M51glD6WYJTapH8j9
8w4KVEmhTSBrWCZ/TD77wLlUB0YjjGp6oSvXu+7iTZE+83UV6KCMuwTJorrExLWq
MqY9CeaMxboMTtCkBWS3tR96Che8LhtA2KpZ0j84/uqhTl0e0G8m5lzbmkx92OS5
K9C21mTfWRplVgLfrg/9bkLuThaI6NYIOjL2GbDdED2W6uuq+pNb8c4R7HhhRrru
AjZxkpEOh6Zrt3pkq+ay69ULe9SPw1d1HAIATTM7Gf5w0V5ja5V1rv16tq9McNMy
yox2rf1mxe3xOqvwmHNWaCufiz+UMMDor2IPponFkT5h3mDwbuWnok4yrhjWH6pu
/awDHR7iBfNe11BVczi8F5M0zh5g4TDRCG4WGB3/MYWoCjFPDa966k9mWR84rF+w
SEHNvuMeaggkiSCEECJTm9pqoclQK/DdZfNO1Zv+Jf6TihBDM3i7QBxa/SupnmNQ
NH0jAv5rVG8uExhDs7CAVo2zupofCO/9LnbuRdOL/Viwb4aW4poVHpZ1Atn1ee0y
Z+o3vujWx3XWwUxqfcqi17nN99x4OeId7jQsfHAWZDMDXM+KbUl0FOorMz94oz3+
YHijVdCQN4Kql9/EWLSYu/QtOddMyitHX+OeBZDCGGOBV1Kof8FrNebrm07VOLye
X4DmOm3pVxM/ubRr/2bpJEJO63HQRdm68BWgnYy6SwAGr3kzr9JxSriVzwzbauv7
SiuBiDJ+ye49EF/LpF3bmkXhKN4pL1hYtYw2UAVBsb5i+0WFbM4jJEP9aJpydnU5
H7FhGVS9XYQEOShJkVD/KGIAP7rAqnmhBY8YlIXe4raljp0r9Ke7Z6c3VhrDyfy3
ZVwA0ciEP4tr/9QFxJplENwjjMvrlu+Cw4mQmRUZ5UPZ1STCLf97cB5P3t3zRavp
egVx0EGgtJNCX4sT1ce3gJUM4+KuXm/XpPCDG7CtfjtdmKzmSrUjfXptubB9CdWV
lnE5SctyveUz4I/T7q2b2cT+44Vf/2UFae1P3HMGUWGbJ9r/6lFHMLoCAHEB2fiW
Trd0XFtVkxkkdzCZpmxpniEvuvXdlHNdpnRLF1bhq17e5DwcI0zcOcuvnXjqJJgF
X95wRSbajYfcCn/cjvaycSeY0gqahZ8DRsg9KtVz1MvuY9xmT4QfIl0yAr4+ljPO
lZje8OSo/390lk4bQZcvFbvoltKGq38cwKN9mF3AH4cYTnUaPaC78kmY5HTce2WO
jvAShdJGChLjq2wJfxwQqd2+H8T3IhoYcAfuBQd88+aUt8IcOq4b9nCjS2AViB9u
pNipY6dVQ91mVYR3R8UM/fZVsxHXnTubyQ5mkpqYgI7XzwFRXghgUlYZ6CJ/VF/M
RURCWd8LArGoEQL7cOOmE8Y6PV29333VwS60wDYL0x8o7OqTY+AelVCLffhy1ar2
07NKRo0BGaSkdGc8L6bL9ZlQQ2iXi6bjhh/HipRR4o8zdMWYPupbNANDa6UV+1kN
LAbVI8/tLgbUPo5G3UaYKiMNlwhXBrZlXZYc131ETdCKggoGx+PPQ2p7wjVXUimK
JBxBoGgwC5nMzdL/asi2DyPg5pjOrAmqNRZ49SnECvQSZqTDeGTZAAcvbW/P2LZ/
spi+5lv9nQSOHPBlf7Km7ZsaL2RcAG9ZHPHrb+ck8kDSfFeMceqQVw8r2JJcSVYc
sktEyeLY7n5eaRNy83o8G4LA/xcK0wgmIJ/XeLs2eVxhy/W0gL+3rbGD2HLOyAjy
Q6IyOZX2WH1oPjt8WwXbo0wzodhfDqEsUqll2fgHEW/PzjeBNqxhjy8MK9Djwvzc
jJMFwYlNb/G/LgSaqGqWshyYaXaY6AizVJwW3yOB6EjvhaOkx4ndQoBxCmMuwHO0
bPyqVC5/spFNXhs1efn4mM6nxOBZvM/sqNUz4hgthrR4T68v+Sf67qCZ87LamFOG
etOkD4Q6yU490IxwtayZhgOZdiuOAEspY6BG0CW67ctqUPZ8ehqm00XCeVMeJ1Rz
xa2ucn+xgh6F5W/rYBEl3RMK3SsXFlJbWgGc9T0qedrdO/qE2wWztC2vHMHOqvsg
I2Q9aYr+8cj7ELICnjk84UqzeIq1i3PvZ1UlmW4NfMUxFrMTCAbT4cMhJ9u9YlKD
/lc37SvwEBUHtcqeSINPcOgNRWlclceLBdOGWqOWVhLkD9pOvNFm79T0TmTJ/LC/
pXo1Mafr7SbclwpzxKlJPcKE+Kv7Vz2x1R3k7+6nKAzYvMQ6dXTDLJMLPkq2cLqh
KVKwWrMlSQfCngHhDUp1hRzw0GsuqR54bxtua8xNqFc8XEf6w6dBhhmvA+mnrvEF
u7kN0ZolHs6K01dhJ4GDAmYFvrsaY7DDlwhDol05omvDT8IniJl1vy1DHFNQfZYI
Kt7zaMy4Nobps/u3Sy/4rW9SeY1k1WmL71EzafOkErFKk5ZMo2nXlQfgX3mnovTb
7XtqGXq2Xxsc/b5wxtuluMI1ji3mxAuDPGOjDZ6xCHrluSrt84Q4p5qYEP9TCKG6
qFFeclzz4XkGUAH16/EwH+XzsgeG4PBrPbi8lrJe1xbVSffcoYF7gH+UhYNjc4g1
v0A2noizhLjKvwJNs1IemEGF2ij/DRGVhFupPC6CMOFcyEIiZnqDwql0rI58f3Xr
Z7C82mslrkPPjGER5ejoiqsTVS7G63au0EIheEjH+y5bBFVgg0paWBbiKNqAPUYd
gSmvI7j+7ZOtCBT9xtxUAWIHfolPR/c35Bwx+Ldd1rWWgKsCUmKs2EjLiyDvxps1
GSXEOPn2xNWTrc1EUYJioJyQtBD0THK4eJzhs2mDlJS+VH7y71QRfwvJaOQfDFfn
vsyaU+kOaKxWA4oMu4fpjQ8HdYA7bptlD8R2nvD9dwaqsnWibJHfI2SDYy+jIzrT
7QguhFO3Jt+nTmRgpj9Zb/xIpRqdKqvItCXoC7Mt2+yJPZb6LaiOnG+1MXhAHgjS
DqBcniiw2Rd41WJnSZpMWMHlILwF1/viCeRpo52S1hTMEHx/7YSvFyQWY7f2k4/8
XvWbSlT3u5w6RFD3hZWmsjEVsjxkE3aKei72PxpmAvapOxInGAQKtIF5nAowfF4b
pisTMfj7EtrbP9As10Hi3LTAueWb+qIaPR2p5pJB80kW8D//4Me2aiQg5DG2pglD
9jS0YVse1ST2x7/MqdnpMhdPIOcW3TD/f/EP4aOPI+Fa4qav3AkjgIbhFdZtemLe
D2RRDccMEkzprIR4pw7XNWlLea1p5EKCh8491BaA67HWAa+A38bzNNOopW4xys8x
WAq3lG4MuVJlpClt/JTMCrCj/BSqfbRZU7+5W+YIyhNoEknN/0HM9wakJwfquqYB
iM/SFpDe5WyLN7znXUIDO+TDGvGgS7H2Uq44YWRj8W0H6bu7qorsrbNlztVVfc7Z
Xdmr5rlq8RSJTI7a48a1iRUKM7ELWnPUZ7jtSCURW8kHbRFNu5y9LmlgQMPV3Bwa
6PNjDDC4GsyQBCmF//+x6xAeB1ewHWpPVUI5EZKTmV58pURcGFAawQQLX4JkSxZr
8jrX9zefCw7pWofFTrs/En8iYDB/7g7hCiY0cX4WlBSYvGYCjvGNBhsANfjV2Eaw
sAqgEYrcryAWRbIEAm3UXMVhX+tFOQdNwOMYI7VgS+5lzYRdqUlmJqIrYo63kJ3R
16/a9g0FyS8dgWS8tkMWCxKS7r7xnC7TDQ6tCN2nqCVj1/fXTC0tnY5PKtvhUoju
M3taaw6mBpNkRy2oW8keap0DfNLRf6LqqNy/NscLA1PlObHzenjmwvAWd1t5Y5xb
ma/zduGfPvJkThrGSZFGRhk1+1JCNGTLeB5eHBGn6AqkmKmsq3k0UrUEc/+DGL7U
wa7QHiuzuCm7B7AmZ3kUhFU8beIaVqgGsr/m5oeurYEDvYjRQEp9OTswNZEeJ2SC
imEyaqhGmDrd8sZyKLG9Om3qWf33IjEbBGo69FwToIHoTARJJt4FSsViBOb4bRkM
leMCZ9/J2Dc1xJ7PZZY3uIpC1fxWSqFlGLn2sFWcNut/BdfwDDiBg6JBffA0xk9j
Yax6vkWI4mSsNhKgKeJiB1qKSrQ4qYLA3L8Af+91UKArDGnKbGWyr5lXyFtufRO4
+G2jSeLGcPXshhGmoRXlMECMmYRBFdc5YPLY2Loi3bUPL+XHpDpECi3hovSCxJpH
bnpltgUA7UGpf5ccm8g3M2goVsArbW39tFpJUHbNyGhOfP3Na7eLcM89ndNpldbz
ZN22wAdcacGOhr1m78FYQUCxeh2sNcF7sLLNb43uvJzh9bXW2aN+mI8vUpgN0CrY
MvE6E2DsE+dlBiZF9gmkyq+kmzHkiDvBY7d6XxdnzaRNCslIqWjq53F/K3bnvxvi
CA3K/2efDDL082yL9rNjZFmjVIY9fuYXQ1y9y9SvGqy8uk3XXm6bflrTuBzmjOmX
TII4BmjAI2wmcueH7TUkPunv4Mf5EowKUJ8cmT6zBAsxvKvEtJFlXeaBVY6021os
k69cqZPu0vS7VXnpL7GlJPQKI2TtM5I9zhUBaBy9uPeYVWZnGgXIZ0x3wMf5pPNq
9C8Oz9RJpne5fu4xl1MkjNwEoExbrMzgJiIWT3HYbDKGnWq0L/yq7zwy/4CIhQJt
DDxILhrrrxbpI075jfJoHGucVni+UnVS2sW3eaS/1c4fDPxGbIVbDseA1QCqEtF7
jBBvYvMnItt4gWda1z1/RxKzdhWM8VtDwmgz2QMnJrAGMMuwcytP6DLaCWkVHvcg
xZAbofWBY2mhRBBD2KSW6W+kasT39uKc+LeIarmA+NV5e5SfskmHtSO6R8WuTDyE
pZBvdt+SU6w5AMQELn7U1nR/gewCB2YR6xAvjYq6zFWlA4rhXPR9Utg4/zCs6JtP
hwPrwVBIdpWS+xQVx7uvPlqr+oJX+DuxsfcrZhr5zQPgCmoiTuIstWGVwOHU4ZIw
WSvds/N8DXxKF1rrqUcvvqe4Wi9+mXZvhEB04x71DJ9ZoQOpUiuNfHfnWQmnPJ7O
1JxlncbqwrGTMdxFaAuMlWAfT6x86ejMYUZAfyTrcno98AgebGBFOj31P4f5pzOZ
MwkcqITZ6gje6jRWeAeAY0J3SbIaOCHCvA8Uiv0y5RnbewVxW11elqhcNqi+LWT0
mftgaweg40uyRthMNSZbPPTiqDzaOuIPY/NccNI/Nb0g6E0CevzJTezjxo6wXJYD
5NRdGR8wGIsBAjsJmpzD5DDjPvTDfPqqitjHWMgLzadaGQCFKldu+PCaDdhxzkwa
V+muWaQpiLe5FyyoOckwoGqDY9iJTk340PeVt797bit7sfxddC1ZjX14SJUpIR2K
Saefa4b5PsElD+v8f+wOImOqc7YxwB/MWOSRYNx/L5/Drf+Nr6J78lnevHkXtc7i
uGkmjD/43nUa2xzm3pfQy8Eb0LwwJtUstqAxPgcjanSyKC58JtfFjMfmQlaJPH8b
R3P3tFmQ5VTJZLEyH3nmw2O9F853j/7Wl2Hk6IHH+8frPomqkTWHzi8jQy2+/wOd
0CiN8qnMS90JKVXHfyslItOkqw7W4ZB5kLP5ganytWoUVCCI0k96tFBZUJIrzW87
kUiaY9WjuelAQ3qU8r2WVJDDhdhOyKqELVuxtIF6uqUwLZceyJt+nDhTDgAW+eCx
rBEBIrD8rqBdqApPzLfEicjp7LD6DfNY1BJ0FFc42JvrJ8K+l67AuTLY/F5BECJh
ZLsnuF2Bbkl04Xip0VEZxjttsA0A8zG202DVFsXaRMRoKFb0pK06Sr/x8nSZSF4i
Shcji5pFr2lIsfMFj2ObOvI8O0e+DP352/gUObKX4UWSg1d16bNUXbBedj4A01WQ
9Dwu5X9s9T11txrGS63aMjjfeAg7ASfNKCG2AKXDlNWQVf5ZgeyGSkJL7CS1WoeE
2hCliAv9Y/Q1J0AlfyIb8AGtuw63QR9HmRQ6J2yLDvf6LAk8YtHJbo567tbKtvJx
PymxbGZWJB5Qcl4Cu5RCsDH+MZk/hcopng+8boQ7GDCsg2t3tFTIB8YfO9NJBPiW
87SfXltvT4303cSbv9xjSEr4FQaEcLWcLEejMOUpv/qa6qugK551afHq8P4IXdFZ
pVVacJhehU3TuIKGRemaWzSaa2Xit4CWEkAjCHdyOK7qyNdNHfctJzLKDHgPPPl3
aWxFhGoqqgiKRdwuGPen4fPh+koUADtBuxqy05P+joJipm+ciwuMmfu8Df1Xz3wJ
4deSOl2+elgtuOe8+hMoOaT+DYeL4eXtWpS3DGCDmLNY8Aqc2KIhO1yxcIZXFXAW
3nlJtEWTM1HEtiIOdtF5dKCnqPo+uqqKCvfaARHg83HyrWHhBz9U2xwP1kRjcVUa
8RfVgDmoZVRB2IyjyG/Ju2qKCHl+g8wubICKk1T/Dglaj/jJ8MhbGe+pmWOCMI6Y
AfLxQeoeIyuk0w3Ex8uvmyCV3LQAT6RMOERbUYQuE5aS9vuMuAMFv7dj5ikc7w4y
7/4FXT/InXPkE4Zp54MOjd7jZgZ/3VWyMDE2T6gGwt6rgSZ7gS2eHc7t9hTEbo9h
X9gII1WriwpQjv4ml62S/rtPc3l4NLVtrUPJOC9QC5SS7S4N68x4YbN7VxdJQja5
Qb5G0DMgiTD7sU/eMMXVS1/K8IgUo68EKIQzaYVvTJo//WE2hF47uHn6uSIs9plE
BKHJVQO69LONPdG99Ss3Fc0eEqIr7HddG/iwFiX0oFOGSYX+ot12ZhC7mD6EgL5+
7Uvio2DYMgUNJ0v60qR0dXaO4l25sA1THN2h/mCjneKHon79Rncu6tr7EfH8uULK
wwTeVCBpMNEz4DhHvCwrZgGyIrDuLHkxWVzQ0dGeYhhRoaHVUIsv3IaepWTHx7Lp
GefG/CBGFNx3ZpCzJIvGQDWjhq8GhkL56XNGEAbknlXp3Uo+EP46uzCUFiN4C7mY
kzxTijr3+xOSLzocclX7xzCXCLpJj+GYJNIKHwmxWyHBB8HIC825VTbOE+q4fy4G
mKyntW8FtNZWrL/iIlKezqMlEATkagbcqL19W7/jbdrWe64fGFMcctW8JtiQTZOx
bJsldTDIoPKfeXDiwgh3/fd2EzICP7zDlHZxV4OjxsSajfivBBMx0ZYwc2Gm5zPR
42MPkBjiI/aYrhwI20UFXYGwQ4ADsm15O5gNVtfJGCuIJO7dxcUpKaJRG/euZIpH
9XVEhJAPDennPdY+3e62Gh8s/pIZRFYEOFaa2ifSSjerhzfcnKeKoQx6axuDlO+q
1stDIRrAm1+KN9VmwpldDb94hyHTQju16QHw2ffwUmPV/U+EmEnnXsKFPb8KXsRO
QZ4AfRG02+099xXkGp5SNeqGMldjozsU8nfoqr75z4qSPjaUXnlYpzg3ECIwaUIE
kYXahyQjo7QHkRMHd3bfXLSK1il5g+Ct4lNMtUfatjUaoGf+iA3/fgUpK4inW51M
VByF6rNx4kbvycrBLjEsFuBN3ZoNbTKJ5q+5P/JqWgxxWtty7RTgMzY6nJpY1bk2
kv/lTRLF60Rhw3F4W+e3kWPP4NNwtTXwhA45Q9yzYXlUmCK2JquZLXhEnVHCKEJV
eZsxwAp4BwdNTibmTE8XcagGc6XNTcihp6mVnt2XPNHLM82CfHvvPlbfH7USCK0g
aCJI6Uwkh05Wbt9edHDcYDe/L6MDUx/Z+xA1I/CBB8KGWoW3DjlrQOYdTV9fD5/l
EF8MYqrOu/BLOFm/eMJHXlqvcbu9K7p/jfJZs+Tk/X1LPU9/D/3u5yecDrHgZ1o2
R2XZ9Ef8RVZdh//bhfvmVEVs238MhefKIUWSMjJZ4Y2S3HDYRlb+sy502Uul7aXz
SJQcfza2gz72xLwqDwh1YLofGZ6c82a12uIF3dGRQSy1///PGeJno7Jt8/A9T/nf
brLF4FQnISMXR7D+JQiqrzf0i2XMWyrabF0GWWFdMkrFxyT1VSWc4WLea9He/gK/
rbpodEAPgjAxX4yTOiNytIwUwdsX5Ths5nLyhSvDMxVpLvfcXrrOyorIP5sBiAWy
ygnMDA4lvlTMnzmABI1vxAnBfPlLfeEFXbieF16huTEBXxb9+zqso7cYmbBRxExQ
/BsfBJwYKwS0cgajrC3jd166jHmgUBYzs4zC5D/61P6Ozbt7f+rZzDfza/QLgse7
XK43Y0Ni320uLZ/O7hnbgIuooqSAetlWJ4ipvrcriy94hmHr8nl56upD80gb2Hul
TmKKLjR/ViF485fCBvSEWLm2hMi8AyevtOtu5QQkNTQkIE3jhaJxbdQPwQHlx5WG
91ll/qtwlnZ0U89sSwWuyLpL59O45J8fecM12ytiX33XiUVzKNPzrcy/KdIPUL9O
3gqB5elC+ySjcSyAb/V/fAun6Cv6e6eyeaAwIp9ZA5uxxLBOeicloBTQkalkkrkp
Kc8MLKfI9wt67TzwlW0kDAgGyC/IthE2QAgNhuDvPZWqJQ2tHK1MTNv4sSMm3fIL
S+D56vAqGsXTtXKImK/D0m7J7mKb6hxRbNa8lAQxgzzEGz6lyD2DVE3618SBoZhR
YkhKzrv8tyqQ5J2aSBjRA0HAFBOPhpTQ9FafB+BbFrhMytAI8ceASS3zj2aRMcAK
UB4LmuEaGxrixHF8loqcUeIFHEYk1MFS/OYWQ1yqisVOSK5ezHejQkEZ++P33w64
TJX2lezVYhmn1NQ7S/YTqQr/PnQujIyht1QNH0nRSHiSel1H+cW8LxLP34g4aVMQ
m/wpMPIoon2yT847n/Vd3zR9tC7+aTTcwkAPjdQvnnXtOQVYIqTXAsGabA7hdobL
jmPkrX8ngkbkHp3wVe4xllIw7mkbIz+90jgpKaNUgZlWcOMIEVKOSCJEoF6m4uuv
Nzfoi6b4WOWzkGxtrqGyHmr/sXz30gfqRzffRj2kounMU6a05QGdXL1+ifdxQZvL
fHrjHYvGr/J7KuqYdTByuVu1SYgHHKvTuxZaqUWcfV7qsMnJ8RwBfFeJ/UpLM66v
1Eps9ufuzhF61Tgu2qgGT6njFWurAtreMIBclXnx73MgxyMRA6J7uJvhL+hUDzo8
nHJiakvGZ6xO3eSDEO6nEXb8EOzbxL3nkCz1OVMcrCu4QoFf5efn98Y+nW26O7+T
8V4CYTs2/oSJs7rlIiQbW8YzdtTPW+lZQPfgIZdmXj+GtfQEq7jS/RO0HoYjzil/
ERFQUaf0qf2cJYVlQpnBm0EEP16r9DHRBZKRvbOxl82bgzl/qiZ2G23Y+bj1i5kr
TkbQAlJDSyIlNLVRLrGyyZwJNheGcOUCQQk9chVXw79bUEVhQl8lnJJj5Z1Ne7bn
Y6crKX7zcSvHaqifjlV9gK+WYU5urMjp80YaYR9XVWQ/rg1vXMT0stbI3vteEQtg
Lg2xI0tnMML1a1bM6DB/jMaNVX9B8wgoaQzmpAw+6BiU1rIZEDM2dkQfccb3euVU
SZH64A/0xlzdLGyAS6Wj7zjn4pwqw7uU6ZE4GOOIjcVNMt+TUUtvStMCN3H9+wME
d8SaZibXbmskXATDcLQnAs2jxJrzfJE6CnYv4byKeM8NOyKGxyZuwGP/hIGQ1+B5
ikngNelVuK8SIASIP+Mn+05w0nd7FNKVBlwsA4zgKiCLYDip/oGg0pN/yNGc7V6j
gt1ZobLoU5sqpX/zl5aa+vsIko1E/X12lGeUQJgvQFlqqW34QCnx58f0IZHfyhQa
/Kz/k1rwgXOHzAOzdmZJjECCg/JoOpDqyEKJRkrm4lrPld6JIQOQJGMZsVCGDxnl
tDcQZiUBHcOqYU3wwBmi3dol6CLwuOcmLevZ+XA13EX9nZksQHPRh8D9C+h13PBd
taDKuzejCZgmqhbHLGUH3jxyrJ9Rd7azoKbqQx4blFEHp+q50NEmwSSvyyx0qT39
WGNPTVttMNYEIvFmSuUxeT2jCgFDk4FPofShlH3O04us6lcUMSCpsgJSno8Qt2/y
t1oaq83fUHD8TkFulwm35DiYDpd263GK6MiG+tRp3VOQ1iBWiREjnVggEtxlgYHQ
iaJTQyT1NAM7rH5gcrzbrDjNxpKwdI/9bBMKEw8korsoQeujuyp+TcfziqJJBhJa
3TbToOIzf5YpYdEI/2lsfW2Yx4BVehDxhtqwJxfpDXb/EeBtp47vsfuhXvq3dyKQ
ToygEU83B2mZd/g3/cJ2oFsNhcX38WnGDZfhR8EM12qUeJZvJFuoj0DYGjO/Y70/
yEiE0zxZNT0q4+ezQ1kzOi5LHPOHRUONRPAIksCtuYp6Ziozdz/Xc5/pClCwyByi
BItwwviIXC/ZQ2brqJuFtITTzo768BDJe91xacDeOe8D7BCcuKLf6tG4RZe8Xj1A
JD6kKuVI3sxT/I9Wx8fr5vRnpNVnzAU/Uva4Uw/Yj6xyTrE8Tl1BPGk5KAE0b5z1
2sOms1zqpPSCqmAfTvVfzObGS71JWnrJ1fymQ1awkI5e4lok88g+JysCs+/95UnN
6VvYdRw9L7524EgHokzj7m8gEeWqt/QDMaKHJfWZ6ln5YsFb86Ft1eyaJrMSSTh6
0t61674SYYcZDdD9sSsgxutwXb3BbKLa8c1haWleq/dKmEoxUt+uGrq3zrBG2m2I
MBkLH/O/uErJFnEHVNxVs3lPdR7rNTstQrn+CedhJSQeMLPO+AGx0ZlGmV7c6FXn
OkyasB43M4jn6LoTHWxWRhv0TnjlxszXGdU/Ner4pMkFqa1bSgagXPTzPB1PP9JZ
mhdO3kSHJYrfDVV2fHSgbUAemupGzCj2rcnSbJQCwccjPvxrYxM3yFqX2Cu/gYPX
evCfZrDKZBIfV4DmQniLh74UVrneu6heEKRxKyFbYkr70fYmNEHdtSBV4Y8QcH3D
RSBiwn39A210k4ajATgtKEbVg7tpNQ3BOara+VFYtmDBpdczZtTm2sZln5xdt03l
LjSNnHjj+sRkhQtKLgY6qkx2VZ5aSFfxiSN+CsepsDn2FIu0iV+ZQLewBO4f6GzG
DTeBbzDeCvtLrJqvhn2x5FNtNUreHruHJcri0eTNAQBg63/LVOM108if8d6fPv29
wxbxaAhNDBTEw9xiNm0FUsOu5417FAhTsHLPKqfgl8URKpMlROJDm7U1dXrGQhx4
VFLr3dPTuem9eA+1EiONpbP2IL4ZN15wTaRMZPlQevzn3wMbIH3QW6agN0TBMHKa
2CcnxHwWgXZsYfxv+mgg66THDIDeH80KTffrz2zMYlurc0H+x/u5QKvoWMShsAQl
nd3k6WlvP9VB+lCmjyTF7T5gXUxTa8j7dQJCNcaULYnOQgSQD+OKIq1BtrYo+q4Y
cc19yiSaFPI48OkbSRdLUeL68Vfegf9AKoIABbpU1lbJbPw4pB0L+G02cYG/Usui
BGdqE/O+DuDnKzffxKdtFKXzwEqReMKkWMLwk2beNe1O+G1A1fREZNYYsCnDCJYl
VoJ+DVr7dB1AYMU+wBwnj9Enl2s7N9gtihWkw9enGyhRzP/9HhukIL72DtzNGqeR
4CGlKnrZCtZ2ueRzz9kN4EMk+yX/X+VzItdYgFP2q1Xhn2ZT6fiAKGFuSDFL3bcZ
sqhHI4F+/RG1D0Dv/FKNIb0vXtZ55O+1GWmEVBwzIKspBb7FJuPiAdlj0i2r97ED
e/cZEcHNwJy0VEFYeFXM80o0VHLlSueWfVgk/T9cCeyXs8283gVeElIdH4nDgXHa
HSlwakd7HAr1fqHbKgqF5uYfHtwedq0Egt5d/dNlxmPeyFJu0UAhXbVZh7vAAbOx
+uOzVYhiHXRSBZFuHw/cKFqyxylJfFpG5dz3mxk2NKxvrDvKMeNm56Kxm01T6hV2
TKNeCnAPUjMpI2hDphPJN+NJ2oqodMJjmg6vbfMyXgcCb37OqfvBcSIlBsWckoR1
/iXtAMCzWxdUoXKkIw+4J95nC4ulAI1psOHqHvpNekj4xp4R9inSMbIFt7u6qWkb
WR6AV5aFeqal41f9L2e9aWCr/ayd7YS1DrK016dIU9s77gHCUl9+oVvkQd2lvtmq
kmerKCb0Hj3L5FyLvD4fkIsfCCL9top7C8ypcrXZJ3vQRPNE1X8t2l6BHvMW3fg/
v5Z+ryZpspiQbnBXzRvapjK8hohKhYZyyop3fnd/ZgseDfzJXdy3rDBKRrHM4Sgm
uTWO1BhFIhfOUULBIQvY7/7CEZult4ix4kSIRvoWPv3ESbzs5+3IsfBna1PlaF/x
DiBUT24cfyrriTDgnAIKjJ/wP42QAgpvVk42u+5AGeX4DcB7l2Mf6KPqqSwsUz6K
Jo5ihJ8mnK3r9gYvX8la0wNjvbawaAaxiH1TlPGeltEfNAkqaqKuHi6bwqHATObP
1jWlanlwuXbspSCHPQRQ6GHXRePQbxxdkGJiL+Dv5tpbdvAqIrWy61QHDsEpO6uT
jg3YFxRT3ZDbhBAcl24xNf5Vz6X9BFOqG/JAy7gncdtmYC/E1Ts/feV2wFg9MFHt
eHOkzHMyOGXP8+LroUm+HEEo2OXLdpqQPgGhI2jEyPJR0NJGq24lLDf5LX1c+Ere
C4YMQYSvWXkUT2bMTokzD9ZZ+oGNdV043QkqqWAqStDcvOxIJH4dRyjR2PvfLceM
e8UTwk0vzyoRQPw8/lfbFol+yeK7wjMEITqGZa/6UDbSc7+6tpbxBtnh9HOya9SC
tCoIwNQhDJwYiNoeK4uzQHSHSfKr+UvqEjDajIc4zRCrSlfbpa1Bztd3bzbvO1d+
jHm+RePopsuHVCdEoUZdGaomKB4gi6EniQ5Zc5seL9E2igk1vNTqCNEhL/69VANM
YS1K1dACMwRlTqH9N93EKYHjrcojx96OmIj0tphq+in7UOCIenUi3pgxvwrZK8o5
m2H/d7z2XE99OTwXFa+jF6SbnfzChmRb9xVrrh6J1ovWr/r9y43dMvZo4yg4WLNQ
EtFBa9m/30/FSnQagFL6HY/TB3skEn6fpx8eiwPMgXEZTH6MrnlR4hJ03Ippti2w
4Y0cC1Ie/lJaeNzt6+uZxr2ge5ZCkWBqvPPKvE9nGbBoCST9IybpjJgTDg+VKkE+
Oy1gC85Aim2ZjZcyKKfc+lcXI1uNq92ZSZ6m4+Ou4oJcd2xr6Olr0ElXXp2+qOgt
/RkFDcL17xyh66goE9I/zFXKyv4jJiv4FMQoi+LwFQPshDajf1XiP2oEF5y7Kedc
Zj0tXxY160nha0iNRfV/Lm2j2WnsHqVKW7zTtziKPy7AUyp1xmoMZKuK3mUr3NrI
a38mDiGeTZQ1Ubz4oE5UU2npFf7tnwNQTbx1pvV0P+6BeSZtOwOIW647JHvHaktX
EtX3bAbgl9RJ20QoPC65usW3PSgsgMRmJLwbP4PsdLQcOa2oo0cuHxew7s9DH4qX
2yzJL2rg+jUmXypUsHyVmpul9tuMdG5DBcS89mr0PKLHlVncfORD5/8DXgdC6cO4
xLOjdoXTZ53u75Eu1LBoWGF4QQyOvBYtQihMJvqmyY8oQ4vsesHanCJ/wLIe0LUg
Im0wZOlBO96Cu8mSDp0rB5B7JGTSwGHR+B8VakVSUxIulgSNUndj27YcrVmKCqTe
mNiDLGteKKh9sQDrHTlXHsuQdlyL+1Lw5hNaJsPNmBWtghRL9d9EIp/c65y+8CUq
Q7OU4Gmzmt3GKhSG/1DaGH9hPOU7Ht/jejqgcj79KuElWAmnmNb7eczkN/6FDWja
WLQ1gOt4q9Dz5a7gBAt7ZvzDuk6nCtSlCpB8pgClqEWDoy1M8y5LvtYUWaQ5Yk8X
kvdR6A4I3fOpCToNkEyRFWEk+UcUD8hAvT5efF6Um9noU0mFp2HzJWTkkuYAeRrv
DS9TJRHoE2NYd3yHZ7mGZakTSHHlhidcxzAovfBmJVmYs+xHPWAlyPEKHfLlwkfz
9H21a66KlPLZaEVFA2IuhZ8VlttIQW1YtCCB2oE3StqKzrod0GdZhV8UuKlGS8h1
1Qkq0dA5hQFxVLlJn2Jriw8GPF4efuefyy8bBwXJ5KfVJoU9cNJt5C1SOl+Pp1X/
gheTS60kMx91qSyFr5qPB3Of+givIO/hmzb2PRqiZOdUwYT63D/sK41Z5AQkev98
jozAnePzwNtESjugyHfyHTyTX2jAKepHYQzjlblzQC93kMHfRsIZ56xOgpDxVyzl
OGlh9XXIE54di7Mbr++EzGgR/SxHb7nz59Fuoy7GLH3Vqz/QQ5MhKQ7eM9Dg2gE9
iwATdaigKezHPOK5HGBGhJtlM8VmOmUYDyX1p9CzmUXzLblWBoquIid+YZqbxKxl
Ht4SVUvdV/U0z0/EEoDB3NaLcUEDrXqHdeE+uscYjAZvOXXGdpuSamMjTG3VoHPb
5ZX9G1jDJ3IPh58h2Y+c2qn4VtCqNUSo47FdOYAt+ZB8EbyCsFOPpYjpOypMhrlq
H1bRtzC434OH2CmKluMa0xUg4hrpYwt0Gy+O8OJqCFdPAIyvTCKlm2VJSqJMqoQb
3YL7vlOzjzpbIXHSzFviDPfJH7T876vVhZCRoFinrL/2XUXUmNRZNMaeYcR/JfS/
cwWPhahQ/Mb0RHyL1z2mfo0Oa/ZyWIJ2eIDu2LCZURqbxRE7Kiv3Vc+6BEjzsoiP
PRHU6e4Az3UKLLF7mzd8qoE9+r8DwjpON8LDZvHC5YeDgnwlFNmr+0ya5kjeboOe
8UYpl12it2d9r0GdfQ8A7qIpmHoCTGymUdVZqsekiKPddc1IKc0f0+ewmQo0lyc7
g0Sf8yoFEk1xECtnJ/zky4/SFwiCJ3Vmdarq1tDsFs1f3PUIsv0kqVdxpxRaz8h7
QEiF5wdWDgADiN4xCCS14EjV955kx0m4HlVGYzQsx/zfYiFpzsCKoKHNZ5odp1As
tHJ3QbirgKoOqQDfXJTh7LzSfqffYfmDZJVITwVeiv6icMK2zqcEAJ8Ul7PwtLOs
QrhGcuTZE6bom34sKw68z5j55giWQJmB4jfq83+h9DfGC/vRkGqaPUPygHgVzqN2
IlEck2qa//YfaHMY3Ze561+x4mWmH1YPzbkjSGGM7WEi2txOwckRv9Ji1OIbXPmr
vOat3mdlGjJPzUd/nhPM0V6UNa3py9LHrizMQhTywlMbMPyhyLDEZCgESGLbUcwQ
NRd0Uqf2XkX7a7YbzL6h1Q/iR7kp/uBKAIp6nQGN7RUZ22lJFrzulCC7X9tJzhRx
17hDjnwPK/RvbRfING3mjiBKbZJm6dshD3l7lV59eetP1WyZmtA3JLjSpaWxzIdd
DQF4QJADchG60UWD5MXP9Y8DaLCf9sHZgeVmCOZ2AkM434pjGYz58n3ZGoTcK326
jOfSFVm/xBIobEJqJFNLeUxy90ysaE1aWawZJbArjKLogT+Hs9f+mxLHKWQPgTRf
ha24PFkZ+Hgz9vdsuW6Ikn/nFcgipene+MmQ3f0W8FJLgzUUX3ekUhciDn0xBtQS
1qA04myPCPzkSu+xXkqsKgHgi4GOtGqm0gQ2kWo5n9j8s0RaZldQmP+UUWLSbQa9
DG0gn6nWPy8k4vfmqX4J/gijRg0Ug5D4O3PLfMCwsPWwh9A3T0F1ol67xfJRule/
5VI2zSas/t5G9NVVtG4jHhTZk1UIaxpBKO0Re//0yNxhR47oqLLKWLmkxNlzHRp+
Zktm+1UwDiBExc719feGsuUTAEPNKtMnGZVlyuKVbNJl4VXIGQvi1yV/tXtCVwET
dkAa0Ozej2g6af3Zvq8qC+6U5iHyVEVTOJmcKDv9nIJvKzYTMobk87jCUA78IIb2
54w5Kq17QMPfi8D7wX1NkTjFVK3dqmw36+dbba6Hkczy849nnHFHT05QfOxD7kZC
+rNLh6vSgesMwOSoBQCsIX5JC9GIQoR5QJr0lf0bvjlCFNpRZJ1xh3BC4k1Zg4oS
aOleWW0I18T46JpQVb47jOMdqaYxmYqS56K5fa9vihIU2m9sq/V6JPNGHCNqGbWR
iqRO7sISEJZpMecS1LsYakpqUEfhOdfCPQGX/DW95kxqyb34CZ07Q9kBietu0Gdz
pXMXWuItpOINf9qeKeesDzKiEbNfsIDZTUygfg8LpvwlOYdyuZ4gSRfgRxg1cgcW
/4/pENyokZc6u/Q6LLt98Hm1IeYqS7IifNabuIAdZG1Sp40USbsC9vHj0iig/x+M
Y04iSkiSb467NaEQoXRXL4GsMw9cFDn66vQcNWTj7RkHH8MsQ6izIkY7+eSBqFv/
w6PRiAgWV6+Hdvc60309k9UHwmVUXhtlLijFTLULxADO8yD1KVYMWVRvYorbZM5t
UrdB17/auAU9AEKsPKi52mWCckC16Cv3i80q/GGUXv1rv553zwhIX1/VMjpNQXiD
L1kO0ZHPDx2gtBSLmtqyoRPbssF9M40Va/x7TQLlJra3P4VW28X+91zZVdDiHVjK
10svsn5e5T+DPNOvjw3opmWIBROn50nN6JppIOPS2EaT3mMAsCvbpNReED3NMQMM
g0yLNzHVR/gz19IOetBCFQ4PSJA2KeyPxgmntridO7gUTijUz/D35SgEW6aubWL+
nV49sP3uck6GZOJ0WtyAhHuP2ViejtMQFKGLOHVQivd2AsypiS5llbCDzcx+7e1K
snBcXARWMPt+mevCdTXdJXkAhYXoGxaP0SSow8MUfpdI3rMNY+ZIM8GQv/bRJXsU
wePdkzKlHNI90/9UgdSBX/xQ2V5/Sbbp3vA91W755tLEipYugp1VGWestBWFRwX2
UA2RExxajolewgjnxwDI/67NHjjY9/vC5hGZ61lrmqPye2UVaA60QTNQwyVjYXFj
3ivYl8btZbSIBaGjQn1CCo2lVVCBB+/NWFYdiPUWuetW49Q8/tuoDOrvsd5jxiZx
vBnpI4gaD+T2cl6gQs8uScnARQgKZnpufbxOeya9LCyHxgf8Z1pwxeRcJdGTk7/j
zDe6mnVnVOPGeVqEfuoXJ32fq8v0dVQgRjolxn+at8/6eYjxg2HADsk80IrH+x/v
TZ8iJ15quZxLpuJ9T9sH5hBsFPJu9jdpP3ntX0WdepidNLIhiTI9XX9vFrHVgXYs
vCI+IpKozDAiglu4klVN8TQZBBmk6nk6foo41A4Ttru7gNG2gB3zZMShKjiY9B9g
HwinFflnzJfFiwr5ar07kQB+OgTpgp0vuIr/XLTNdNO/XbTCtkKiFaf6QPM6iAj2
++RQTBYP042MskqW71VJ+Ye+9pMPyPBmk3m/8y3aPHkfY/WzDavbkpv3HZmuGmo/
QQ/K/pUTgb6yk3OVTUpUdbJCrg2FhOJDmEpf7Blq+S9GxRxgj/4jEmg2JrkCPgcj
RTxDq5yyGlC87HuxEoTTP8rGn0HGz8uVWMDHzIM5t7CgD5g8V3tqtu18RHM8d7ms
js+lLDeYnQG0g54fS6LEkGzut1FKTXAHvvqqkqbQt0UzzrbEEKgsUY3WivZ/C4iP
XLy9/t4ma7XHfCxmoI20elvgrNkuKUibsF4Y7WFfrKCH6cHMADnnujad8mFeknlu
6nFt0Fil8DOE6KES/IBVRb9e5xykDr8xk4mKW07KLVqe0SQ0gErKnlKzwFH28Tdf
VOI3da2MJ2Xvj7chNps1YpI+9biQtFlSgk6MEPSCOurA9JpePQPWEdtXrztk1f2D
sxuOrOVVpUX9bWifEzBM/zRfzS0sxApyZiV4M63BkFmBGj6EYe8wD525qvKmj6GW
mEUE2pajI6mhAWD76iA4Wq1oNNaXhn5jVuYmiQS/kv22JzP5hSB9MAIPFirIZOJx
/OJoDhZcRg3LW6IvNdR7Nc7Hv0ZSItbK3bzYuyEKWxiePAjwx9K+TH4hDtEf8UmT
4+tiksg9C37SpT9kMyW1Jo7SP4DjuYszMYwmpn1gvf3kB1HOqup2UXE69L+R6JIo
hASAWj4RHpygb5/dLdvhQGMv02HBby77QAyZBvrcxkVIJ09CDYnwb0KIv5my5XWn
AIc3/CJpCZzpsI191LnEB5tzmEWloRDbWDU/VgHHy8VRJibjWk3OVT0ig4msn/ao
MH98MCu/5OZXxDNBQDprAZES4Du+eUjpjLZXxMP7QUzF1zmDsTBo+2VfR1bejQlr
F9SrwBEiuYj9xuyOvvAs9v+1mSZuHJCyzYy27+sFs0SqzM0wEPmvjk/acKGXVuFg
atEaIAfI4vZ7FBgv5bBbRrSzynZfuZVedXmwfCi4FsturOjIBAwiNrzlcraWnqm8
t4OVCSN6oHNW1MykrcI8qAgKg9djBt68MXbKEfsRbXSkdEEwrWgWyE8ewXIuDS9p
+AOKJI9/T+4DiS83tPapn5TGBHDGZmk9hmIscrGIYwDciMPVVLpb/AuWBuN6Ek84
d9UoNAS23oUtcXXZe0G/pTsyI1Bf0LT9WpLKGGqAjODb6m6MZvmR41VJgZySvhaQ
cHjd8cqj0Pk1vjTqMqMwz3biH5wOdUpSz6SIy9Nu2hTZYRIW3VCDbxuJKgoEDPZG
A4wHx8d5+gmVnWKsk1JkYjYGaikG5rINcebWfI68G7tQE7fY79ydJTrfryatcVd2
UdKlccfhj1Aa1zDp2tyPAlPMdqLkxbe8w0oP6S742ODBxAiL3UzBg5fiZx8pVrWN
izcawJlRfu90IN8ApBoYekz2/TQudl0WtcRcKVr6GWghkOQN52O8ivsaIIPLK0cp
O5ZJ8MIKrbc9j0rvveKG1QiLqI1DU5htWM96oGHWXgt/xjL0WPR07qh/sGwYhvIz
4wfbSnCNSlo8TOP3nT5tsoAj2556nrjvPJkGvLPTXlLvorKsy6tQD0JXPl3Ytk2O
nqN4ASOHOkBcxuBbo+Xp0CSbMDAAzkyJdXDh/Tu9UiM1we8wBvf5zlwOPXEnktVF
p8vbsiBb0IttBoWC/5+vhgCyRJ5szuh41oJycZUAuOag5LV3cynB5vB4Fr9QocxN
cLgnYNgw0naUifdKgpg1Yv0J2wr5sPsKJTECtZHJ6aTWZwEuxTJ31lZnSrXVIZI2
gF4TKEDJOD/p70lHYne0oGw96dgkmZJsGNDFNCJ+ACly9P5rfsZHcmZiYAiHqhyw
rHXZlW6PY3MAhOQ1cTVH9qtKIJ+PxmXI9HSgq4In2JqBF+l0TFphDVpWzMXH+QZ+
XpagEphj0UA/UksgCi4zxq9dwU5AaYBDPsrDN+JbJectEOBC2PVcV/6QHc9tUiTR
gtG1aRkM55hczhtdKvgmAcSiKCFhiyAPK9pblg6VmiSp9GiN7zBUGN6cxk5IDocH
Va0p9gyyXw40PDVUKSuQnZyN3YacMXxNOZA15/IcscXHjG4fmmVQEuysb9EB2bfY
FUVCPaycoGpF/3HCCkqD0e8n2zZe8Nwuc+y6rkiAQTwr1KUz4ZBvoKEQI6qcA4hC
wKo5iu+3jxJfqhU8aRYOMaXyqP5kFT0TohG/LwiVQZZ0tAkZPhqYokvroSN6cUBb
KsL00mE5gJtlnZYKpasH4xo1LRwgAgnLD7lIVNw0RSjaxVSsqfdt0I0YwR6x0cs9
N/rmd/gyEyvdMv8DEtNIRIYJQV7bOoQO8gTWw9TFopy6QJ+mcvXqlIiLIg9R+0Hv
Di6cnjFoMMXQkUICC085ymBrGGnYuDbAQnkFsx2X7KkkvpGNHbZUZbgGZvZaJhop
qkGh2aHi7uCiya/L6xC7m/67OJNjr7b/4FEz57jQrjWlVNNh8JmSMiyksXpEPlB/
KxKTxNIVNNphG8lsDcp/T661a0J/Tjv20TZtFZ33Eh1dHAPUX869LvIua54l7Y+B
3VzuGcjMl62bv4it+GPpFN4LVCnvS8xX5dgpNlK+iqX2CtKInr4c6nLeC6QuFebh
ZCGPZCREmE0z42JKWe/rstD74Z0HPElkvRV4dYBGkIlfyo42G/svAdoi5n6u5o5r
hTRZ2Onj5lQ5YXhzTQWsoWmu5tJcwge16oME4BV0/Z14esGeJu20GiqWSUsKbuFP
TcVFttrZqn1uycv4dFYF2hKz4rA43q7EOWlWZzAVB4ubH3zBOSPMf6EcrCgBgWgF
7h1JRZ8abKMbhafrxkwHyjasq83ii/SqHFIgKMVJ9druismslPQfMaW1J0q4OSHK
sofZKtbjPpxAmMCl+sokLzPN16TNSFOKCef2jHj2lO0XwVL5B6XRmbobmfj/50dm
JkdIHcZfPfrtZuUYEN98h0t4N3g2tzMb/KtrBjnhpdUOu5zzEQx8viaE7nVjMwVR
oWaGHH68DEndG7G8P1BwyLO+NdtgivtZbKYTiS3GU+I2A67TJAyRzq11l+OxGw6d
BaYtJitkr0h1nkgh01Zy3jMmztYSfrFt1DiBvj+gHruJw43xMzAoBIaTeCxTcWwn
Yf52CQr81gUr77HqNVAR948I+IP+dbEkg9yyNGI2aofKREoMDmiblQfTuG3gNhr0
ybfQtmnV0NsbN/3uPwUnvSUm1sWWpSMRIjCFf7OxEzRLjihpV6RphUKMJcV/VPnd
1n38t31MuWVNVlqR6DGG67Ul6/ilAmxrav3EcTS65v/AkR3A3Lmau0B4MSNzpyu4
3WAl0Nr65wJqOw/OJd3XycAe1lXjeYdLl6nFhiU34cnhsgG3JDLhJ60nKj1yvoa6
R8xnnsvjerXxUc7cNsv0neJFjzk2BLADdL7mAY3ghpUb4AVc/Kuv6Gyb6p3ceO5p
kT8oV2GXQyo627yM68Z3u5KV6oSsVf3O9b4DLjIjJi+JCfLJ9GT+xRr3MnGsEiEo
or6/xoq2sf1HbG1Bkmy7uwJJ1g9oXHrhIfCYSXWp0ysvDiQ0NtiRwHD4NE9Yn53W
Y6IWdg1+IzDgxewO0ytjYmiVrSlhbTsLB+iOHK+togrr/Bm9+xbYIoCQmxPXfecI
XT7r4zvFC8zMP0nrabdjGKU0RVbG6Ju1ssdWAvTz7vW7/hx3EBEa6EHr9rjQeghU
ARKbA82/njBVWqzjcHXkzjCrBKRbrwk/lw6rQWPtQVinFr/JDRaJtvIJr06bJRsR
M2eEBEKQxZTPljQyVZRcVOZ8hi3s+9l5rvaONXq/mwALy7NimHZSQTwu6GXeNBZb
uMP6YhnFdOUTw27W9EH+rn+lxFUWPHZ3i3Uy5DXEAHFMssdYCfkkluORT0jaIUhe
a4zB0tyLoHZCSFzYTghq3sg34aEdXO7aN7OnWiXd/lzCCoSBqWcNEIiacCSurShJ
GFZb8Z/s5tlEBki+NmWIkvRmIKSbi1hTe0naYQ0VfHSI9Qo1bCU9dWrbmNK5D+5o
HDmH222cl2CTKGSThTAzqVV3jVaKAI8mvPZbTh/c+taOKrFH2ydyWoRxvgIsOR/P
Z934C5UdmNmOQO7Ix4Waz/yZhInrZ2rCUIJ7PtCfw/KSA66R/HOhMErNReM4/uZv
9iwIwJcCgrBIDTbvWXbKsapmkrxjG81ORdUKhfaWNLaa6+5ch3YR95eZ6ohQVirW
8Y0KIprWu+ezo8DueqDI7h+dF2ac13gFDy8eOYMXfMEZXTGu8t+OD3bM3o7A6xAL
9u8vwpYSAS8IXU612GLSiJWRfo2RTn9SbujexwOV6EccnQkeZFQH++U4I3AYvGdg
ttlOsIst/jdPnVsYIaY90AuzXyFEi6FFGlRd2HpcJEZQSqxSLqjUkxIcuHN+m9PB
Mv3u2XTz9zVCbr5J4Ft/x5CF6XNtvPNejbmJV2UiESi3P6CPgQqf7t2XMo6BOI7b
KCni/Uf0hrgKJDDPz0nJVOmY3/Q9odUJ257VDKDcgA+nAciKtSxQdJ1mwHZxKvd0
JyA13TkbcUvv5mEfSyq2uNm5WCksRmLkhXqFWNPZvW8Cfz/1HVOilRcC74lDDFec
6BhnbnWkl3ukOtorjkaHMExO3PQGJB8+HTK68stvULDn+EiRx53IrStSWZ9N9F2g
JVqdoXmRHEmxGUfZkDP68jP6Ns55/7vRDZPz9/MzxycYkntrAj29aIBs1nL9FavM
1udWYmqux8yRAf+yI5as9+CJ6PI/IyzBRp5ikI9zbzkaI2R8lOPyGIRuuIkS5z5Q
yO/i1z4TmnKlO1fTJBUuzwe9VM6LMuXVt74ahv9DyOpvGcNKNRtlaxvXrbGQYvnC
kw6NRWqsKvRE4nz/Tb6Bc54hez29Q9hq7fpIjqsMCSy9X8/gKWiEZT56e8Bjg1Nt
Z480+PWgfF5LJ3G59Dow2wypd0C4RlGNf5mbHd1ViXDKRaM6N/N5VaNLRLF0tU7u
aQ7ZijtJzAob6rGz9gqAAJPZf+ZSSHbYsOaUJJgCf0ZsF2T5xMFP0leX2CzVizZF
Sy3saF44KfioBCarW3KRmL6+bHf0kM3FWU1lzCo/ngyK0a5RGnlVw5WZD22FtM5R
HPInnRuDXO97ZtTp/Ygd4q/QMUvq4/96/JEXuGK54krtYyzIGKQswCJyQjW2IQPD
QOx9lF4jYB11AYqSSvsd4fPX7SmsvtoSEx5tfszmqZ8tG5oTgUcO+cW8J1ftN3gL
CoNyoCTwZscAD/alisRfeDtqhbqG1UDGWDN6ux6fnH8eTXoML1gS54zYgG3L/AIo
60TwdxwcMCmHZkw4m4SUh3HwZwjnBrS/K5/sCNqiuY5pCEmRD8yghxGpB8cdC5GA
kh8xjHXiUGc3xqFGrdoqdgLjuecOAlx4x2KeOB7Os+3eHj+iF00jwd3uP/zwiPtE
9r3DcB8GgbT4Oo/cANfIkTIxq5jEg0A70l2jwsJhdfVcVvgLjv4eyjdzMCpJ9DWR
gJmqENR1i8ZT8TnMUUo/2fYUgkhx3iadftAXpxHcK+GQSsFRKGCKVDV0odJpQwDM
LjxHvhgkPbn9nCwoIkm81lLl/Qht5JsiaplnawxzgLsUFGopgWNMWHEGH57WQh7H
KmJPyYwvaFk1gH/u7fopyrF31P49YYxmXpdRTEGZ0g8K0LMFo5nFYujFr3wEEi8v
la/MVdUyXFUmGOq8FPWpO1Q2CX7b2hWkNj4yPllSOlCVSdru3Orq+aMUhEfSTXAH
MRG097AhxBdUcXCz3pveTS/E3nm7wsizyYpaf2jufPPvFFx1E62Wd9IweTT6tu6n
4Q+P5t4TcoiC2y7Yj2xTH14XOPQGjZwY+dbfYq4gNb4z1k5YSmJsCctZm++c5MTU
YVBvjb7PXqk0aHu+f7FcnTE1TJR6YZArVHx3QhHBt+0QHrGKXuGvz7MVg50iZk4v
baWGfW12jvDA0ONW8b3koVQSFl55mbed1UA9ZJvcTkvooHDR732uYy19m+ieTHiF
fgNw4glzt9CueYuwSmsDkZsV2GTdF1L99GuCt5W+PHtLKxMDzO0+zLc4TPbmn0FP
kbTuW878aQuz1cKulD9KniF2iZksPfZxz9QP3eHC7a8RNaFuhm/FYHF3Gq1RrqZG
9Hpf1A7yBfm7LmV8MsrL59fH5VW2n5Qpwco73MoAM4YdNfewdcpcr0ytz/apFhLQ
XI6mJ3p2N2bww5K/dveOZbQkVPTYlAgoArP88gEL/r4xUyUIy/BWAtVP2mxbhTe0
G/Wduj3eSpIqCQnUti/pNe8at73uWwHH6/HYlmBvCZ7UQxTRuex7bRYldoxx0b+y
eAZBlX2vARGerXqagR/nTzVn3/z3iIidYqz2YWZKWtpFGz7brJor2yRafZMTwGCg
0khMfD+DLh9oPal2qYUrte3jFutZHfm4RJ5RG2aDCLDw+Ud0+njeOEEZPO16fQ9Q
HfQf0za2xfpq+1YqSAZ1T/gBqm+0QXrjS7yQOmPnw/WPwtyryYxLpAVO0zrfctlw
y8pk0Ne8LLO99seDtlakABN1UBZjPMV2F2s67lnKq8FLNfbRi4I92nGt+mvRod1I
S1Ak00hop3+eIMKSkVfxKfP5mLy/U1WeUYOVvlC+t8BWaWrj8Zy2X0DIZX921cIy
VbLAOdMM2e8UCL7M9gdEnZbjyEbPEqFO7xOlfggWM0aOSCkz2YpfCIg1+GXodo7m
FkRICITLCqqeKpVBWK9O6IxrPgwkdnNn1SX1AxS0aXp7CTgMm+l/5fRBg1sF/Nvk
z9s6AgOH/5MYsDvspKgqnqbnqOoD69VKGTXHGpV6PkYrf9xHzsTzROdxsYMK5cMA
CQiF5kukjwNQRThlc1k00v2A+jnOhNAUm7CLrQ+X7AGICg/dgamkf8XmDxayF7IT
xBQXqK5eD9p3/e5+C0ey9VpKRq9et9o5GW5hmP7OmnHPloSQQTrr7jzKdn9jhao4
3b8i7priO317nTO0KQik4WReEhcXInpRy1JXxHjs3Am/UveBtdTwws4GyX6HIX/o
PAEDytptC2KAhkhoWAgathhUMA00umXdD7NwZ/kN+ie0aroTZ7o4wuWlgl7K7P6Z
YLhKWDKWiG5b6bYuCFyn5IZB0qC0bEdgpyLzSkOmPOA6mEAyp7n3BgD7HyFCelNv
olg0rSx3EnOKf5nyLB2648xWyGX25Bg624GFE+QUCgUyCJ67jDeI0ddvaz2d+6N2
vCaEEcNSeoXLcaWHIaBwBIV2mmwvLLu8aA2CHOoVYE+M9FI5x/wu3UwrboQRRRIU
XO7hskljaRS7jiQjL+ftdt4/YtmhkBaGTrChcVOUc44PPKWS0ki1KPBaqPzf49vQ
R7WeYuOuPpiLYrjXZBTHsvoQ8fEyZlx71D1DziVbJaSRHRUbhEFOcj5vr3VIYjJc
8W0Sf1MBxhIGuNSPUiV+Fz/HE6lTLQe6rHsXVk6UsFMBDvjkRbSW3T8ABaL7MIoR
xr7yZmyOFucTpX+0OX0h+e+1eVKU+lkzcNn+Zs79MjWlDZVo9EoRRv/jLMLtlpqY
xOpHvGqCdQnfPW/shnIv39QW9+hvEkiP2psLhb4ouikFkQxjtIPRkDvtfTeBnIzw
OF0BsGGPlZOpvb9X9BqPLCB80JO1F1os3W0p8jiprb13ap3jf+Bn0jGZGuycEtpF
50RJk9w4RGli4pc4/U3s8XHer5KVSutiqkklNmDlAKo3sSQ+Xs2yAESN9J6f6HlA
xRTt/6hHVoUZ5masnNfoOn4IQ1j6/OP5jLsRXFvcE1cGqZRrWlPuPqc/1OjCVIPN
wlCfYkKAB0TZj6HZQLooO2WRMopofKG37RRisLM4S5RQ0M9oufm2VfT6JEIpyD+S
f2FTwHcdzBh0Jp+iCzQBsmZ9jaytNNWDPU4vydO2fkxOBBAmEYBEG0mfvTawLZ0b
LGLwWKWROUuljR0c/HT5oyPvhD+G8KRN08dk7k/C7OLLpFTOdBCbvW5lw76DqFm/
iVUXTaG05UWi2rHc5Tw1ZIIXHtY9TXHBDYhnTk7s1DspN8DL6riDZMPpaxyh/9kn
UnWZIUPbua2PdDUtF3hwFOLUdwuwehIsSKnZDE/Arokm3c7c599qnS6ZEnk2snyz
Hbk7EzpKfglO5198IKUgwTtCYsSfBFAp282Qz269TWMiOhAMDSmTowIOCteN327F
Sc041tSG13l2NZYMKdGunTBzez9+4bkWvhsVPaLzfVBZmxz5ZI/5QTBDTwq2gcYy
88ZlFeBN+jHEVdI6gYnQksmIPTRKV0vAq+hNPzEyZ61R2duSTojCntFaCujquy9I
EwgbrCsmq1a4vyaG0mZsdQuuAehLMuB60QHdtyL2oEnWWgj7zQ1Nfjvqy5H2u/LB
msvTB0UvqXhsFNBBAh5+7DmdS4mSakgWH2Z9eKKV+FlLXsew+q7OMTBWJ8Ny3inY
+UcV65W067cv1zRtRjSY0DHlE6EhX1Vw6yKpw5AshCVIBulEsboluStoN31yOURF
dNPAcG7B47gwg6p0/ROZV9J/RQwh3E/ZP2Kp5kfdVM5DjbDF8gJXpDWX2aI4eNtS
v/6OBMDmfwvwCLhXyR3PUYo+jXlYdkndm3LdS+MnQqHP3zJJhsKBVXebfXkmxQdG
bUmc968rSLvz44/ITKXuDrN4ewnIwKdGCRgfFUGVJC2AuvFzQ4g/kwEWRjIAGquV
Ub/NGqg4ffHjWPbWEcdKpy31LxUN4ABfOCF0evWhL3IrmRj5pY83b40Ovq4rQvKC
J33sa1LGlxBtf64C+/n6mJ27Sv4uIsLFyxAcYGo+5dn2YCPynAdXlrC1DYg8DMAz
p3bC+hm8UR4WsNTgN7esb5O4W86aOZUHGhqsX3rdpNwPPgftFb+K8YxFGTdnXNNI
aKC+tAQacbfmGSWPslOLuCxMMYZlMy6IQBmbabrbq5SmWFnpLjfZfTSAUsSepnVK
ybX4yNzeUkPVpuu7WgFdBO/9KauexC03Dz7FYnfB2wLcV2TtC5oNmmvn48kVkgOv
3SzTc9RVAMOQ5FQO1dvQCvqXGCaP9cz7pGPBnFfZQCEc7sVKGye0E+Hn7raZIeQ7
CuwOt4Eh2dXEpnVWWJH8+sfAP0irspZFHVbV8+pHMTvpOm7eHyZi6WiNL0hmZyaE
CCom2teNs2StI4/WoBYs8DDTX4SzLCNwqUjqTsfd/kun9PM9Kar99+T4h2W7ud6S
uEvXntyVgWrRAUzP3bJhflZKzrX7cwT8B9ew5k5a7r0xCPA6IrdZ5QBrubmtcvq8
u2JVd5M2dxk1rgCwnCSsvBXWta0WCveoyZdNo+5o6CYTKx1XOxJA9rwFzQ9wg81/
oVK+g0kBn98mtnL9W2RIWXUv2XR9h7s4IrL8nZRIDjsgZy0Uev62gdQ4/vGA84G6
PqkMw8AXfFSvixKeRoSkXPxOCqLbs4sOrCMuTFOnET01S8fsU5mep/RVoC7gwis1
pSpeqdOduorduQtmvdCz12IBcvP8ZHX1VwhXOoUw17Xoq2TC9+3SnGzJXIUenoRh
7kxbR1f0WHfnLCji22D9tN9ZdwpYVg6fKU7yRSk2j65FHXsCXAKnUZMNP+I7B0gj
PDs6cVYafNgdK0+CYXEozLrvPlVdC9vr6zhGzzUvVG/rzZHYn8XN5EBo9FEBODhu
GYhM2yR6CQJVjSYdDrORkfuO/i3Nzg8gmUegdryq9ymHlUqaBNXX83a0zqiI7Tua
KnLBbUjAKrA/ntTkrGZ0WM475AwinPhnIfYQjo5m8Y+eEPtU7z+y+bnY5xeMby9Y
rOhpYsoWGWdAJJdzN1ir3IZ7eoivwKQDw1zrQ1U7STj1dZS1lDwtzItmXkqFbLiy
CMbz4pGaGNaMbhMOoEMSqzF6oTIyaLrAz5AgrgGkKRplOJ3yPZKh8nxgkOJAGKYy
e9ICJ9uf1sZKzkHZGIU+N0/YUUYBOaOBRtnj2HzAdMDAbChZqCYXq4zgvONToIxK
v6VzmQxsWKZ/VLJgetPAG8LyCNZZematoyIx25ynmrWax6x72C31VG3q7zPnl4Po
CtiH+sQefw3M0lx4v3ugO/7TfsaBibGtPChB5UP0arBHoTjqyIOrSmgnCqd6zAJN
bPJ1ldHZGBGf+uJIRLPFff3toprPCM+K37LNPYqyYEh8o5Y8SATZ97ar9wNURR2t
It7Jv3Efp2TIVkyiCq1TuaQNgFPoA6iBdSvoLwFUwvlPq+r8CY667Mdwc3nUwLWU
h2mfsfmOLHLcVUgN+0Ba6QabPPlQWK/TP5jb+LikjbM1cJ+2thK+25ycezPzYc6Q
kYuGdf+/GzGN7Ga2JuObVhl1TGxvLS6DP/RLfbhxQC9iOmMRn9SvBaxq7PL2VwxJ
q8RCPJ+QI74dGhLav14XEYwVSiXou+ZJs2loymMieQHNFXdHvJM5ZDFoTlEUdnFi
K8SEd1b+Cf1lBCwglKpLQYZ1LZo/No30wOJnZPrWh26+Kxd75zKL1vqW5fLLNSKn
J2zLKQgroqtVTadrYmyj0TFkIG/jNf6NWpeBN9RKVfLNiqLlHTw5ulRIj0sni8Gq
n9rKsu0jQ23UwE3XylbNSy24fvZ1w8+vU7qdcYDeRUJijjAVRnCl6CeIeklMAY0M
gxjRTZ7QdjzGiArPKutxwBPTNyUX94QZbLDGyClW2Ex481hFpLKN1zD9kSmCim7Q
CWlv1TfhhGGST6Ui/KTJUaUUvH1gIp12ew6ALJ8MVHEoUxN2lnMHvojJLIy6uasp
ynqDrJvHKEfL8yjqP9dcF5ZV3dkFG3hvWtUn1tRIwqzK08SiC4O8odQF7K9heyC9
QTYZxZh3Yx9ovNHkVpHZVoO/UgaiDuLoXahBgLcxQ01WS0skys8jz6LeInfcNg7N
VDD4LDMEjoBmihyZkWfAeHOgEVUlX2TSGkrTpeXa+f674gNHa2NI3WaJQYwLGEtP
RchHAi0ggxenxEynKKH8ncZN08OiHwJx4FSO+ZLb40343KvyYaoo5XUr4qsCmyBb
n8wILxZW4tulqbkV2lJYmqwfSfvJKgcLqA1kX6MHm1w0ADetVNS+8eNg3QhahtkR
TADi9rLSKcu9JHA/5wWj//x9CsbKGkFQ2bdF8XvIMRXjdOAhKP3NJ5YI7EKapkt0
yl1V5vr+2iW+ZfGGfD3c/UgyKXmOWqi/EDKI5kqz3DKLHAV8g+pZSiQl1LBE6Ndp
ED5adzkEzT6ixA63OPfcvo0XPL24+URuYn4t35XbAiPCtClNTwOX6GTqhtnm+mZa
jSyV04I5T8pAKZmPA0OnawL0SU7DgWViLxvkDzxUy+rHKSw0o1/ORNJ7uRJVfdP8
mqXhNnkKJxdM0egjEASyjU7PlspILd7C0+P+d4N+0rTdG6w7wDIiflUxlpFAJvkd
KV/BOgVKsciVMtIEXXnriuZyDRf2E/Xq8NKpi4oDYf8KKpyr2X8zLKhMrb39Mx83
ZPDSIi+BvniuUJFWNEzRAKMi2ZZxDR3iO9hSF1hvPGOK/M9iYmzmwSiOox3cTByf
owjjbOezak8ZZkdn3b15j8J6uRMrjAFNLp8F6/qpcsju5EOBNe45JztmAcJUhPcg
FiWlHvA60nR3FlS7NNP8HGMco6p58EZVtQOiD494taLxvyjnfDspr0sbsquM6yrl
JjaXtn7vw/0muJ19cyuIobuZDVqSy+C+6ZxNWnXl5NsHUcf7SIGKufn9+pbHofsk
TcjULE4Tq9KtqGXPsXeTCMBx/BZFQrJw+sYcgI73cZZQNovrrsLmu/Z/Nt48HIA7
zi7Xz1A2NSHLPb2zZEk0rMTGmn671ih3w3CdVq3L0pjYSlIRaJ53if/r4ToaPrhi
IKHWflxaRVjrbWogSt56xAYQVUGAAMU3sL2F1iMJduZG/DB5sYtFDPFEbqLTeKSx
rFctsPe3g3OeuKYO8/VvNCPkPk2WWSgDdPZ5X+iwlJUIJbU8p8j+EXA+vCcqVokK
TwdsF2taj10aPtaxStZ2HwL8fyN8kzbApCQVj2iNqK9XDEo/daLkumSIeDSezKd/
cMYFYL0pJgb2ELUZn3HBsfy61PSgz9D0E1OKMd/1/yGO9iyd3eaFoZBl8YhjnYwc
WviWDbk1iawJWH41jrZqCg++ImvDOs+mJsRt8UxEJE8YNEt5of5DKtDzW38duYkB
+wrzJbCvUXMebDuY/sORYdYY3PTGkYKuTFTllzHNQpxnVo/4W4z0p1HXtO0iU/xx
UbtsuYR19Ac9h2mQM7hBoJnQMDfYvUlu2DVLNTEcPgedKTdT8I2LbaoSyKRralRK
gtxDgzytKIDFXSKt/BtcP58fh9Av7ZlGcuJjSJP95trWHcYdJKxFDBPtv2YnPkzo
jFKkOp7X+/wrxu/Aj3vx9ICz7Voo+l1Z6LiYVhq8gA45ZkoBkskV7PIoFyfGrT1T
fNPDFClVxgJ4YoH+n673KlGana4fNyzedVrvRPaxPkoa9E5itnm+xhk1Ip3vJoZ3
00C0XBlIDLIVBfl6cg0P7ZuBkS+7jfl23LguXxB/Q6c40F3zmZsnK5z3YNGed3FV
s4YESLxl1Bss2cU5jwNnQdVypZCgzIi0l9my4kG9HXKN+86NOlPeL+mvZYRkFV9C
lIEyF9bLszaaVx9HQ8BE4p7sYb6sgYegFRq1jBuHGe225CAjbcOgC2ihbf36DTG2
mjQGBqSlidxFhgYJhHtLkWZgG8naI4cU9AYbX+XCOXYa24OLVVa/U6ZyuuYoFBjo
JhwSgTOEKVaPXSDvKgw8ix+uhRd85YMDd30v5DdyElvRp91L42GdQzr+FIKaYVGK
dheYun7qyGUci6mp0lFIB4pLGvRSwqAvSOLWK+JSgFT54qNIFeurSwz2i5Z8eTyp
rQvq1Opxc8o0XbhDin4gQkhKVXUzt2M1ycVeatJbkd+rll1oyJitpv49TDDu6UX7
UF5OCoBF2/mmgGzau3QzTE7e9HKyUTsHadu7dKNLipcfOVDUvLGog+0p6We8MKqb
yQ/CJq7YMQux310BDctk7OE23t4hlO6ZD/LP8Vr6wzmmiVwfIUfkTQFjvdlQPU/m
qRF6sLDRCeyLLJu1wup2gHrwgrIB6MVf4rD9quperLO4MS985puNN6qS2n4GcbTF
nuvEDIa99HvHF4wLTL3kIKNZUW8WgYn5qNCLoQYiQlw/ILStSIZuTVisqzgfPtUg
ND9vKOyxJG2J4P46rYX1rANhl2cB/K+NezQi6MdPiVXU25ZMjLUSU73dO+/R814M
TMW67Q42EISYs21z0WimF5LiGNM8ash785wZh7kK2wPZ1f5rh1o28emTE0hH7lgi
k1naBmS20WISHqxYYf9c2IgeFUkBM+A5LzIlgF5ih9zA1OzhtLI7SPiKaqnzDAf7
hjMGJWFvnW9SXEbz/9YTnuzxciMMEBiBNowDtsxG36HcZRSeREpux+QXvw/O5jzv
zaAzjmz4I5WOH79164sN4kEQ/Zf0d9mar2P1StJ4mGJ1e/KZ/URD++8p3BvpbfVI
3DkOwvVyttXVJ8tEcvlJk56OvH3OKkGr4H4AfcUS1kMB8Jaf43qzfWYdXcdt3o17
i+jKYxW0lbWaW4lfEzXft/guQwuxN3YJIHxSsZMGUxFFA9dCzPGt1x4swRvQi5l7
VlMW+O1quzSaAH16LsMTB4sK8Z7NHVgbkFL7KDZzlaw1D8xJrx6quHnoMm70eVKL
QYrV4fS0QjzuuXk+R6SgcyVvoBI9W4LxcZwquOuphnVA11uSTJPFuIhZ0w45MpZP
D1EMZiOlq3JHFS28J8BBL8SQDVSHpEr//HGqiT3HJtvBmEctu9xZfPT31Ua/qcqC
smKSu6oTI/Jjj0+/pqimK82vO98zpmOlQZC1XO8L2q7FRe+u/Pa0x3h4knlCjcmb
ZIBjaKB/dwA9bxIYg0d77inVELpkXV3ey0IcYo4b7JYKe0OqyuYcDLfwsWgeTlQe
hsoB/YN0UvvCNggUXZ6RbrIRMHUHOKC0Dxax4rztnpUL2wSgG4OFHnLLzLm0sbCd
B4F/jzBLC9Y1LRqZMUEYVwOqwNEZMDXOvy/7OLXbNAmZR2pCXrzCYO3SEa7VOtHq
B1cJBwdy/50nnaWzM+AVub6/O5chM+7quP2XQJqMKcKqJt/Rd1sFbMOwcP2myYCa
sJs1fwKbtwDnf0jae91TiImAu4b3L/vt2WZOutVUFf+H4ZXbKFWFEMiPmJGwIEpA
LeSH76q2y3psGF2ScaQ3gWsPpq3EFqdqFfdcidfmc7/8/8ftiGlFYjdl7TtxcIwt
sHpTn/f/QZykFKPikIQ94iNXxPXsLTvn5z64agih/yc5wIdQorQhhjoFHXmLtpR1
7r7LF9pEGTiYP9qpInjuVuY/xLlVhA2r+Wu9SIUwqvxIOmTB+m6GTOXjcUF2pqzt
B0p2Rgv6J0aiAOiogLk82qZLguRcNykW1lsf/R1RtbD2e8WpX6ZNFeFpSZwfQJRe
lE5/jh5bVtCVW+xeOZ3Yioq6X84gUhiHL2AImHi1b9ZyWGJgGR/IHt5ySsOZXv1l
3mwM/o/J8ZRRak6c8OV5u+cB9Owwo2kYKMXzL0mlP/ykWCeSFetns+p5tEE+YmE9
AXIJF70+29p6ownuKP6gw8u2d5ZkjwuBKT2+gDpJX91vd9km8fiRkDoOsP/ljmEW
xKEWR50Iv7cfhEszqGOE3bEjvx6CiVpyzamlpspvspc8WNpIYos4ju3b1rlzR16r
fhmjG3D3/3FYa3aIyuVdnuTZgA5pXN98yAdxgu3kWWJ2rQkNot2xDrUrdUHoQSuF
x0jGUQcraBJh5FXPIOaPbuYBGU4GIslZmqUN4jvkWKFEsoWUgrGzicNbKYQPHuBL
0xpVch12LINMTyf3hQU4VdKi+JF11viw3k4F06fyruYJUq7peA3+IhcQaKRS/NxC
emEz9cHiISXiH/fGKYqUVmaubjSEjd1UhkSigVE2WObdjANBnTUJPbMkypknDHZ6
2fu6SvZPYp86cZgj5rolj8OPw1K9BoPNkQSOtJsgljFNFhm0VweJIDZRKG7yP+JN
ow9PMSpQXjBtv8ThwwGCoJ0TUDXteoZp3vgk3IErVCQO/fRygXOa+uK2DrsrcTPV
i7ZtwGEWKdI3JEUioNg0fLyR1moxuAKpRFglS9rjPQmd6yJoq3dUNzCBPSjTvCW1
t+6GCe9uKisihYgg/Foin/ajcysgIXMA/4dncHNQUj9Y7glfT4F20Fccuz88KA3h
C1fvjskFdri/EZCqHTTnXxso5APEolsZqPy1NOJtzwBuURA3m13EgAzm/hs1kJvs
NitMUcVYw6mgM7fOutR1+BtNKJl/Z4muPB6rstixiRR1m/2en1PN3OPzyBXVICgP
8xQb/7s4tw7JOubMCLsOI41VoRJkyOpJAlDl+88DXTtCFgMbxoYPSl/W1FG7wA2K
GWPa/K/VnTJxHeCbKywGM289uIrlT+8yi50SECsz21S2ytu/xrJNvixb0YOq1Z3k
oZhWwp/Tp/QzGNOrMLmg/pFHbENL+RZEHmamYPlJD+dhp/2E2n9OW41g/+rPUmx0
BDVvAtctkEfuyMFEK9W5I5C83KLZS1uj9GW1XFYMfwJjU7W9arqjGXWKZcQ9vMbP
zA621siHaTFODYOPXDGhUIY8Q9IAfxPt1IJVQZBOwzV1KJzQ9G7t/sQzTa+2ayQW
X1j2mlnP4AgUUiqf5Oy2t9rhZmnlZ6KJ8wpkto9FAanedMhE4HGnybdIGklaTIi0
7qpEpYn9toARSoFhYPjIgDjs4AMgDPmRmGHmpVAnWnJRh+g4IjcrjjARLyYmh6DQ
6TXSzmGLJCFrSzwu978bL2APaDefhYheeILPPFOCHFdG9viu8tfsbcZhWmpJdWqp
RuMT3GwFlVrvFPU8U3FFRtV2+z1vHneKcMqZtiPkN2uajlpns7as9sW9FnVMCyEn
j0MsBUURhXvWozoCfJzg6odWIibU4QeRIhm/dojLhr83LOVGAyCb4XVrJLNSP5Oy
TGk1NzZp4FMmqjgu7meNxdloCxGA37XNGPd/hDLZUADJnL9ojQF18cdw5XAaqwsQ
RcAl+/9I7Xhxsj3AobggShLSUCiqzmWv4E/Jp8Zi5A6Kg8xKHNW64dwhg3QvCbfW
/anc+DNhRcBNRi+IR6qPyYK2KDpYIlnxpn3u0ejqmClkNZnekzQa4+UvDoBDP8KC
pgfDtxCe4cdFpqpK8wM1yGnrD2F86+dbHTcUMzCDDZsrJA7Wae6DknMnmtW95pgw
Y+WELbt716eOcNiPGDMmFgQj1sTYvdAGiNN87X/BKgIMRAOd7KdXnqyDlVDViiwV
C+A55VZxkNf+urQeqvPBZySSf6ah44ol1DNhQRWcoE/Ygx8LRLVBGP4cQ9Tk6Qvi
GByqcC9Ku7v6tlv+F7Yk1bHEkdap2ys27L3cYHyWK4c3krWw/wOU9FPY5DnCBQca
+GxEh4H5YGUDYxRxlldADFUGhdN8uBysGbg9v2c4JsiWJppIr80RUawDnlLvm3OZ
OvRGTHRYIo+NVYuIJUN5Hav+tOAxu3DFndiR+m6BJO8LEz9ZsWyy3zBWQKpZrXAB
xp8WikHsjw06uogppSdq3h9aF1cFbwcaDDMx85Ddi0oPR6LUaWZTsdjJH8D4V5HF
Bm28oYLHeYOAXR/KUvs8DwrgvfkcnDf02Pd+sZ5PE8YV8Fqq7vUqHlujYiIbZhWF
VYJw+xCLDm04Aac3Iv7OJLjA/65idqegsAi1lZU66sFOUl2WgSBybkojIoHgUOnS
5L4Ggbnn04FL8Z0p9H3NtqRdRcMKYGkdWHD4cFihDRwEPMm+AKVXy9gyPEx9I3eY
msTIwaEull3HSNiCIDJQ1KsGf/f/Bkh2EisdDzKdV77a4oYvDs+5f812gD55PM1y
v9u44gr2hGXZoKlUb82oflwBh2O+Wohg4mW2p//pMYqHQi2+qCi4yanGkpwioIjV
nr+CG1zozrvGw5xAgsw+inC6UDJNiHu6BNVOWDhQyssonFdA6YyNgM76mCEV5Axs
Ghpf+UJa2bYvj3FbvVE9kz45VDgb0eZbj0+Sd2/zgiFysq6sDU+3jgIZJB1RP4eq
18yD0UfN1mDGA+/JZVDwh3NFEghP0R/hf3ub5QeHhR/BnT0sLfe8LjECSiXJCORt
ScNbwDZ25T37o1r7o4qZocJVXdZ3FeyJZgP7vLkZiBeM+PqFmgK/e19QmUTymf7S
peBKJsDF0XV9B9X4s3rYQZdSJ+o+uha1HAf6M73KCyJjyTAfUAr4vOojzsxSNpLT
vX/V3OWx67gpLxClWibH1a325VagfrplgUGuZuagS4uvQAjoF3r26MnqKXcufQI4
TKxa/Udl+Hptlit1lOL6XroNj4z9HPrMBXGqoPSex4T+zrIHk41nLrcXqNtN3Zx+
fxtrHi4v3R4f+duqdRQhwNtjn1io/Gd6MqMLR8X6qQRXQmntTh+fw4zf4biyMXbK
1zzchwziYqeIf2+OXzEHcli/m82xrHI3H8XrDfLcIY/hegdwxAN8awhkr7ycm1z5
Y/VMBMZsb84rshAZ8M7aJJy2pmdQbBkWq3zhKjrt6jR9t/Lq7af0msn4qGtPcgLR
jiNA40Fo1Wh6bWc3H/YikDhvS5hgi4tNlHpmVp/BJrpevVinuhDE5oqna2zDm2WD
nSdIfNEcGbebgmrbljkw8mhcIvmVtkdDumisn+C9g/6+C9al9vVRXnD/uzrYN4gb
1h4caEvGTMwybMMVXG7hDlR7P+GUuLIFKtwNAJiADNzmQtl7LepNqzUyHtCfJo63
6H1S8DHcJ5JgjterdqmCMlsrLb1Y97Tj4SfnJYrZ/5PyfQqWiRI44BHwH5ME9qDG
10AaTRkmn+ctqM8/M3V/xf50of95OFjCbYr6JcoSw6OS//sc3U9YOCv76mwRncUF
2/+HfPGbZJo+u6hEarxkYMl9rgQSMiCg+jZP0rCBapZRITAb1uSo+xqSWwjmhlan
YHrW/qAXqKKHztwIOlH/M1XfuDpXMbYN6GhpaORNZQZZ2Tj4GujTlzZ2PbAGio8q
dlskD4PLd7I7s49+Ixf0efXnzibObdBZ2kM8qC1yLH0VeRGbJP3LUOhn/mPfn8Pe
FEagxL/g+frV15O4KkxmK3cv0jKbpi0rzymfKJ4QI2hqjGVTX8BIsHCkP+eqyb8J
o7ewAzODdJVEU5neWmhtqQZcM5VdplhMk9Qlg6Sow5U+hZLMcU8wD0Zt57oCnu11
PxU586UWf7vJqQeCD+ZqE2byMi+SKY2p/ten10zhOiJQTTvtbIL2kvWEuhnlsyTQ
XmM7CNPl+N4KXCNp+jomgLwJ5QYjBSqsxFc7QOkThxirF3yDxt474Qp9jgyfJpvR
Itj+TQgdhIfgX6m6mL0TjSVDXvoMTIQy7Qi38rH5jNQiWYUvzYEiwX4A0opw0tdS
0WEMzhwWCCznNrMMyAEDdmzIRtplF3NZoz7zAFUZ1DrVEnd3Ptj3keNunxqHePnv
noph/orne1f8jmHxS7JV3GC9slu5v0QfQphLWZB0jSW13msjUGRlrbyuxZ2Ze/ib
3tYGYPG9X16exiWHXN3zKAfhUrk3lsXhBu0kH5cbLB032/sgWC/Z9g/2lI/cizl0
50p97h8L4VHgo2n2+RcVv2OUd3KUZa5J0wq1BjhCzD6x2Eu0ZvZCMaqB1Ry8Anjl
DrYCR7GC7GvK/xssSLL9qPs4Q1kwmbVwSpdpvArZjvNVzdF7Ti2cZi6+GUPHfUDT
MMI/Apr/2Z+UWdfp1eIbaZ+gowo9/Zc+m9jnBQLSOPeuDOzRyEvxG/1O6c5SJXmv
YkzOzeo7VkID6XFG+jcidg4TtQSBVEQmMXgbGH74aUNsmh21WnOWNfiTMGKaM8OO
liPH1k8aDQFbrDq1P8k5xTyIDohkT8Nz9NSIVreXA5tYuy7vloaSXfF6S9WWJXGp
I9DpyGLDiyxSDjgCHJRlkLCk7xzGSS4pxUl7zJezkr6c5YyWMX7k81ebieScM9Mj
EoJ7JF+schKKYQsa+b42QKQCSyIhIRvJdNecxs0VJ06JV4OdphDZVr96bqMVZe8+
JanvsV7TTJi7RfbMP77Bsy17zENcOcLs1ehB4hxlePMBbR16TLgbvgQoleLn5jIx
1xFmIiouOi4WiFMsIgWvmxMnCPxA9X0C2Q17n3uUGYkVvNwrzJ0fmHXabnAsho9h
oaQa7hFwnC42iZFx4feVZeqy/VrpXQDnzF67gU9D+JM3xerkLJ+lyaGdFFJG4uEw
4HAxcuX+Z8rkmDWv2zHoT+B84tOKFf7LLtq+B3G+KAhOcytf8xynAWRmVaYu8V2Y
+hnGaS/yvfTNqeTlonfRuhqjWWWBk4oreMlVT9OcrNkcXnKw/pPTWRma23/3fvnQ
RD8TjhhZzBQMDJvzRVE9vEn5ZuXz9BXo+k4P8f9ANIMLJmRftajnnFhrUygtjoCK
PwtMyAP6rlwRHm0HmtEiHYipwbqnIRPzogAEaCYcPxTSN6mP+Fv6qNElPiZ+iyae
A75b4pmkmXF7JquO3YeK9P+UL+o7X2J/62FLfg0DEo6zytcdGvKdGFA5/t1I54nG
ZKbGz/ewleL5Q9DfMuEWmaJKMS6szxorbHQ3qno8AFWppgo7UrT/tKlRlOwm0gyG
IVClGLYNsf2ibWkjfuo4YfARnNTG/oZXIkjzEN8M2Utfh+M16Gaf1ode2nWjd5Na
cwf+l/B50/B6n5pOWR79RHJmICYMAuB961twk2HJ85ViBvc8x4AGA7vDPPcILZrc
4wjuCYfSXK+kNNt/ZKmdi3rQQpWuXSjmM9IOewtE7pAZG8J5i4Up/CBt0YfkeFln
vOa94jekh0NuJLmYrtBO74foipZjvIN6MKt4oJEuZoscU7j+c9l98a6wd3nlQdWJ
qJtWiA1PT6mkLIEy/kudpgeuxKy5Q6FRmddMK9oaNvbkNEjAneteSFDpsgkcTsmA
1LpQQSI2hOenGvY7rLDOXfEudngzOuSd+MPOyQaP348yZtscNcmupT5RDlGJGJkJ
r/XSAYEJCGYgLUf26wIorhHJQt9UlbWFzT20em6iGv6D3twfvAKarsemPGnjJ28N
Z4m5QxTMzPR6BSLZBDvY/SmfqmMGvNZkZyjJEp2NKR7QD286RSnuVF/TRwFozGWB
U9AFIg1GwQpZxqx9ohaIe5P3MFPO9OJKP2lyWVQkVnmamRHgzlpVcX8o0i+lrYN4
y2Owvq7r6OTaGvyEBXrdd2eRNdbZL6WHhPhFIu3uotrDVAMVAs+nSixrqbZCUia7
tIWhPRMeuV167sSBbfJ5VfQKih7XBtApowfqgNFA//uOcFBq/SdBsPf4YLg8Dnto
QnOzq/z8BO4cEvuNp+0PW+Z+Y0Dz8u8h8pf8DyxggfIGrIR/14VuxBK8mRQOktjd
nzklnCIt52od1uYOEi3WLie+zm/b0xYYjlgKg1Wmq3G35eknlzI7CIdUXXAM2o3q
9Z979VRMQkikUJLfEMvPTKfCoGONtaPU1HO4wqlKK6hRM66xcqs7O4HaqkM69cGo
HX3v7PYsmt2pCdocv8IWXrjOl80qMw+hM9x2V6koaSFrXL7k/FbT7pCVN8piMZCh
EO+fccGuPQQLYoeH5mzPN2l37eZ/wnspcbfkrFdKK/36sMGib98XyAYFFxmwvt4B
fluncXLAN9TMJzd0gXVKRv5PivbxYgwc1UevPavM4BEX0wkNdr0AGa8NQ39vJ9Jv
0MsasujSjy618APizn/b9BIs+IoEflCbTptnWU4INmwQ2WAh59YTpHWdsi6m1ucV
jlubKZ0GWSAtdBpmp21hzseZYkSeUf/k9OUgoDYAUqR+AL36f4gn5KxYfbzkbu9n
RU1/erHac62c8HfahYY6UPza9vHeq/9K8N7GWIiOr+Azu/T0+lq+1CcsYQpgJSQR
PI4KBeiEdoHgcy54gLl9TL1yssl3TBf76r6JCUJLC4frPBMW1xokfpxWcugKfu5A
dWKQG4K42vFc4dD1e26swQnyMIuvh52cgVYLxrizqJs1MzmJMprbdDQJxA+hGV3D
AI77qleUjaLLwcMm2zGpwS0zdBlQpxlMmZhJ+7RGFKW1/Jk8X7w1mU6eMhUo1Dny
y2eL6H5jldZ+vXG96aJ8rr9FLYjUawqvtZ1/E7UfKaqPgx7UdEBKEx1Kqw8JjwaL
bvCG9zFMleD3JMVgYG0aozBzeVcqCphwbreC1rNhTiw1aLJ8WmUX7VrIhtbwLzDl
khRz8MzUcFDGrLDfED8qbzdAmLXgafDkVyQjfSYMs12kiSiLU9xB2ysJcxrEne5J
F5E9RLVsX4h+daNQESuPKETWL7xjOBUjBNeAXh2Xfvbw3sdZ4uFu+VEnOPAGDdA4
Wfz9W0aZWocJApULeVTqneOz5LQk0JM/10bE0X16HISfUci7iuyLJ+tPUpMFi1Ud
wSvHJCwNi9V+8FF334isfRCqCCmz9yUZZGGuRR3nA0mGYut9tccJ1jvsFhkrsLJ9
vaY3YxtmICI9YJqWAT4Tl9GZ197umfrTwcDUHDJkw+U+bKjM3/YIdVTBv/e3DkGr
O1lqstq+zXeoD8ZwfSSuaRybVTtOQMSybobjlSEr8Fp2co/4pIoAPbSKKOQUhkkZ
9Sv3w+CkS6M7cjVrFrGPvtsRTKOXYLDNqc4872wHqb/2M+OUEBwzAuxOduIi4gXB
QHeXt7aMhl7babEMFM3ghhXcz37rmiZ+0YTmFqE0NmAjOcZEmuQvHIrITE4r2d/P
cP3swT831Aj3V4bj0s3bo7EOWx8rrkdPmnwGozV9wPHU/o7CbVXwcQeo9qkzfhdw
b/xZsssBycn2XyFepTdeMJrgFKGOO6CvvqOn9ZBAbNk26dqWGfmxKAneuD3OIHdY
2Evdm+J0/eZuOZX/zdOxz7h77knSKHEV/cr66lVFggcUAqPYwJcV09mfxal+v+QI
PqPkI2aeY5allNAb8l06HjgZPOZGWYRW41him7w3t2ty/3dcSsbD1k9yRNqST6mJ
nK6AM9aYJOwahEPbpk6UO5GHJSL/Td78u3WCB97xNPYEYE0QiwI3xafUhEomEuhV
fbiuKQRMwoRsDpf4ldcMyW4utgbWvqwPMoAQsotk3R6zKvL20iNrYP8eJCmqHw/Z
yYnt/fg4IaBJb3AN8SZP971heZRyl2FIuIYlaSH1RMihZuuZRaI7tSWefjA0VuHf
LmQG+dOzQRHxHwZDOorn60pPANKZP3W68DFCtd9OJCwx0/y8KkikcbbePnpn2wcv
xddW4Ja5NeTPLkrczCnTu+iJq0QpKm/2cJQGhAqD86LWI0M1RMkTgInVo9/Yhi+L
kKk7ztHBkBOBDplspUrNSG4Ac4qCJQz08m+PyAVj1nSuyzhYJjYa8dwq8FtDLfTL
RygHW9L+4eaWsCc2TwszyKIf/rqYT6gI4ZhGOssHHoTaZcFrPzxw5MpPNc2X9wH5
7T0ZmQh2vHdBiMtobXHlM/P5k0fwwhSCzkyPPx/B1I/+1AhcdXKZSDVhV7AfNTfw
s2+VWNhcOAB1Y+isSaj+XpDK4cB/kFGojvQjYDmWb2+Jduh+TGA134RtlDYNdf0S
Gmgw4D9GjPYxSy3Rrr7pCaOgjMnQXbNrx5cpZ8OJB9leOl0L1z+C49rI3+yXXWA8
yRqxSNtDi0xdiKlRBD6QB5yh1ZoM/D9IWemH8Yul4Dj0PlmFgnHaWJUfqfbQU6jk
2PUsvfiLTkgjK6r48C7r3WTAaovtCve6CE45Imo6J6pGZYvNkKTyiBSKrvjbjmPI
XgOT81+yAgsq91AImTzqPyidZxvXtUHDULrWNxvPf6P9EtFnFehv6doA6zYK+fFg
KaebULJ3fjKyRGqKdtc+a8xIwIAMpurcdcycT6H4XW+Ge+bG4M+AOGO396cVPgt7
x4e84yUiYGIxDyc8u7G8v0JkJbFPRpiLyzTXjmScbEPkg6kHhqOPhCPQtCxE5vlW
XShLVn+dckZUpIxQUjFH1O4BgrZXSGIwdYh73yUrMB/hhpKigzNvM6mCF6vndOeq
uRP5C59wLg1pCpnjp1mWAs2+VUYL0d0qn88jandkP5/xjlhydZDk5Oid8Md1p8Im
GSfjgKRi8SsimWAafBZOjGgAIIes73RAKxu7tHnzp09icIIGZ/GL6dVNRO4Cn6uV
JERrqdrv33hazVnFbWobNpZ/bI98NqIHFeo9KLHjWJIkgdSFl2+yPf55/229t5L2
prwnpIu4Ij39Cw5VWaxw5nudJWVW4IbNOp5JNpdna5nMUJNxttGDQY6kr+LIu3yd
Z4OnXkyS647peBPsP9fAGDo0bRSxRjGR/a84k0RujgnYaa29s/J4BlAUl3cByVSE
MfO+JrKpBOkXyFLGKQ8Ue81H0V0u3ZY5ohnC+JWY6mzNOjhl4FRpKehLlorebBSO
i5MdYrzMZphZMhOcXwg9DTOknLH8h1k/+fQxlUK0iZk7JiqOaDk5mVEwTeBTMUW8
E2ewa5fp8OEJVN/8drcvHPhqgv7wl/kIEirVhFN7A//n5CqgzVssrSO2ObBom8DK
tkk809plEI15d/dpTRY88mGMtHDVYYGo6L3v2sOVYVr8s+LUxN5YZYw1u7sgFD9y
jvluNtmMnivImt+uh0nUVuz+w6umbSBfWWe5yxEM/cJM0o31/xFuLzzVNWijP6SK
FDVrpHXlPtK3vVs1cjdqQ7x0xBiSVHRp7Z1XUkGsF7fI4HLtl4HGPd++QuDrSRKi
0EStgsHzVx0k9/5IY+ttZm/3Y2IEkiLbo6bUsjtpggZV0AQST2mpAzI6V/fgfBtT
Irhrf9RZftnQ42dpjApd+3hgIpbpx9bj6pS3DXyKYUI1Qoq05yNnNVJ63Gkhb2R6
626JfPkexdDX+92aSP+0A9/BrydQBe4OmXKBVfHy7Hy9QdiJjsTgStFo34fnjj2r
R1vEtjCB9HPxHoo7Sh8Rn5B50hErj8dWho9wUKihqLWB2FPjQWR3Rzyyw4uvASg6
ydMLurfh0ZadrVqt463ka2R/6sUeViF6BtNqcFzTyWdAPJjN/qU2OOoGlifDMWlh
ZcVeBYnSACOBTZNZ5Ktg34T1BkaXk+Q201xwIuKS6QTBmu2RTnVazbO05+DKdB9N
QecJDXhofXWLhRqr3BnvC35KKJKq1xrZiLfACStDDXF1WFyhxXoUmEFIrqLLgIFJ
1i1+PgKnxE9htmZFriooU3Wbe7wASnJCgy6sBc29bmc0evoQugc+ybgLaQjuZvwD
YttNb69q0rgbTFN2fSCaaxgVFL/1SvNZzX+WQACajg1ogFXOBvU5nOlKK5+UGKc8
tTE7l2x+zIZzvZLVESAskiqZsj2ys27nf/Fx3frFWoCciebV8r6wUIiPJ4oM1w84
oD1rEvyC3jRWRIIVAqci5jxEnkq37Zp5tDn44PDDh1k6ynn9p6EXjxhV6+Q+LKRF
JiZvx7W2KfzpoF4a00c5SHHseoQ87LaP0QzE5AhCTQP9UuTGlT2U9MdaxHQXojQw
CtK901XJYkAuxjwxJXMq7AEM0a7x7dzcDfx82rTzoQhsNEaGQUJvVWPZqVGUTET6
C3DQt0XXu+t/Wx2xeLkoMM7XcbgqRT0z8m1uHbDVyPRiDQQOoCfRYiIg+wqNfQo1
kKAHz8kdbAjM/6ZQR4hGtKHBWCuRtyYyRr6N060EQ4Oo0dCQxpdg3cVj20yaSHkQ
2npgcsTI6KGCB4fKFhcfUApc/QXarOuVRdgxX4alA28VnSvT0yCrDpFVga8atd1Q
sQAJgx1uE+6+Re0EG4t037HiV6bJCl9YGBj8eh8KS28a6NfE7a8+nswfIuKyCvYZ
6m7cyo9lflv+L8ikKG+82yUc2ejJD8uiUJDUbylJS2qGnRVnzmJbDbFJLhSPrUI7
aUFX41QRyQrqZyexij33Vwu6+t/H274jSgoLfEngeEe9hTLuTgM6nda/7JjG0Elo
uLSuQsVDVr5rM+lEijctaEiWsm9ZrT7QTHpjbQF33IHttK8P6xEhpt6dl7ZcdoyS
DHs4h3CC2+lomvwaoNHsY1O9tEGsf8sKwoSWR6jWDNq+sULSRIRSxedPP8mA22t5
lBvMJvD1S13bzJ4xgLl4CMO7u2lrMN9Czebhfdygt/Rkpo9JjPL3b0ua6y016SUy
YdGUjO9HRR+ZAsJxib69JsQTB9bg9eJ+yBHtYcW+sxZwaj2KEW5wgPlFT3QCS5d+
BboSUwfdb3gkyD6qleWRiAdUy0kd+wwFF5Oae7iZW5mtin0Y9TifJ6P1CB+hER90
tCp8fCM4L3eyzVl6IEFjP4UmwuH+y2l2PeaQ58xOZ+ezm4bwLQPaTAeJzFW1xgq3
njpKZAVdvYcljnbwSP6/qbkEdFo/mVHWqaUWc+ZpwiwUCgHQ4MMuQ3bSiUGDroSA
djXdOxA/NrjyPG20BKbdiStslxfGp4snCZVH3sZONN9TbdwM3JT6grUVmlyNFwGz
jcZLk7Q3LNDttOMosoPURnM1DUnjQ5Za++yGCW+8OvdbVPcNUvibUAOCiI2YGjnK
CCVYi5fcvqi8nF8x97RJdrlfl0mUI3cTwN3xDHeYqBLynNF/PC/nKBhF4hV2CYk1
eOjGqqNKX5BzQIM5ulyoREf7fi+cXkOBCy141PHhxH8/yyMOE57WbR7/o8BKFktl
HB7ZfP0Dh25++fGfg6nsDGImtTjSBwNEWmcdo0dDdT+WGQT71VQVgjmvb4ITubTY
EMRWEDwvVP5I8Fn/LNT31+cMcSRUOgxc7owQSwW/sYiuxkNkz5zCqoom/b4KKapS
9EpjOGUny1wCpTshUrQ+sXn7x6NNlh3a0hqMYvtar6fQ8Ib/6ZJ8dtyXFBTnseRh
u1SNBzHY8BhHuC36zq4IPtvDG2PxtYnmIcdbqMGIpSHBRhEXu5xoM5ofPWzwRW6O
ZNALRpZuHMiJegyWh9VTw6VOsKL5eLEEmjG0AapT4x5ngb/OZt2Z+qdK+0D9tKDS
IRtpat5k4053O9+f7AhSfI82qGPVmytuRLy8dq+IqK2FrTgsrOH2nmHpBAjgmz/x
g3oQ+YLxDMLsrtIGd+kSEFLjrsax++MDZrSgK+1dyyVmIk0BNMZyeKRB2LoT6mAS
pI65mT4OyrS6YNQakNm3gDsVWpozX6emBB/oZnXPE8ONJkTFtrAt7WLPNTIL+84C
TbiQrslzXg16GMwQe+PFKaOymXXQCRl1VDqMZ7uVy/py69aWQo8HWGdogvQ94EMw
KqwL/l1/iyQu3DjC/Vip6JjBWAsMeFoXDbpIlh+LbYp0HdQzURqry/0CCYMcoijg
jS1F1VBdTDozpqUm/pfuSNW9wlRcoMvti7Yn93Lz47ziduQJ2JseOEHG4ZNCdq5W
9ubvsfM8LkjheltNcOh4Qu+KPVfUBWLZ3ukRu0RVv8ro0+zvHyy/32IkuMcU5WFx
X844pir5W1LBRVPkOKPMBusiVR4KimnhYJW+M20FIZuSqr2FbFsHxOiYDEFmeuFI
quHEpPpxE7jo/PI5gxKbHphSKl0A0uoqzVvqLHXzmPrJjeeQxEqa3hHZ89rDR5F6
Uq5NLn8So1QXRyolKkqKMYDClS3bjAH44uA0EPmzesmZpUN0TF5nqeNwZIIclySQ
b2os9CMygeq5IGtrrfQrZvqLY5X8cUyUtWdLRfBK2uzHJSVqFR5y02+PM7ug9gIC
n35gi0b6b2kOJlO4pjjHpLThi7AZz+57TKxpQbON9/R5nQ5GNeXAoA6dVVQuFEXn
M75no/QpEfmjF8LJB3eHsErIS5KZNyxgt+WX04WIiu7pbohcfgbxERXI4r3QtMzG
mvT+MVwC+6qPqBwrJPqSIIfqFchOQLBgVmd08GP/FMg0g83DbxACkDf46zjKIicD
BYwG71gAzqrzrQ2vuKyVX+WwQpZE/gYTAf6IhzAxEAemYEYkP8LOh98rda02Pnzp
9mexP4FchA0eFHkXMxUb7l4Br7ozd/pPHfjoK0KJmSNzVBv5qKO3AxVChbZ1rW82
eKzynTQt3aobJ4MaTej/crbu5WbL2RMXJdllTzluNEwLKkIMIE9NB28VieEyvXGw
U/4HRHmaNJB88OsFue/zNCaz/VTUcPu0vvdIDkMvytTSTOzP3qvj4kKv5rWmN34h
Nbk+dAGaqGae6wX43gx5OkSkv964qN8QU0tWQqbd2BQeXLQ9adTvX1LhZIAT5gYN
kWJx+8seaqj3rqIrELAAiDqVe2WbR10N+dLPqYVoLl27p7QsYfIqjAEONCrgKXjq
muhu9IEjKF76vWIW4B65W0vtstuBBjRyFag00cL4injJF7AiObm+Zu+qGAbUErRY
Q4df/1mqTLYh58IJUFmASyJiMHIEPDNLCoCZ2BqztAMqeAKEb34EIT/1wQ1KOK3q
z0cHXGaEogM1iUygF1chLPSlOk6KGaKG5pk2DwGcPxjlQozV9lwtNObhWmu7Uygp
6Zxex7HcS9a1TCN0+/hSzlI+DMKkutvMnrpHek/mxh/b9BkAnJBVF2sRzOCZNpNs
JRGndT8A1j0vPpVQw6uCdp62kZky8hPWE/JBBPGlVIUroYS7U19t/p3VblXlUjnO
o8QW+7ihqK4a4fTnyeBHneruDjXLJn1uDEq5OAaFQCAU+wy+XFyqBC1vEFnxLGIF
KfVnioYtHRPjlol+w8VAb93dnfoYhTmV0nPTkA1FM6a2PKTwCxpu34/uszfejN9R
DlfytLZ48rq/3H61GvyRWYAzHaznM50Rz9TREGfl80DFh5vL4I78qx87FFbp+Do2
UxUzpuUgPNHqeNiGKHrovVFnbpkyiB8D6+zinTFtlAuGrRXqlt+dMNoKP1rjjeyf
gAdCvSU9tw9JDXOAd5y7L4aJS7zMsllhZUeaSh83HyeXgqRjA98mZeZgL7AWVEsb
VHT/fLbdPHWxDf7MbI10ESBeBl2Lpsl2W32JBToN62CaOJjRJLT3FgZbGMVYsiNl
GssmS6iOWr2oxk2FdNb/enDFRZKP+DZgHPs54CicdTmdwjLKf4W+H3G7RgRNiNX2
/vlkmXsOjCE8f28Ux697EAFDE2TRCMh9B6UyH8dpHKSYW1wiafmhRtlii7Sn+loj
JJ8JZG0Tzv8zHy5KMdSLB926+Oqu64oHwftFDZCHNTQoB9oqQr3qWPxlaYY9tK5y
pVcuBYuo+R6Ab+VtRCRhrILNT87MbyGv8Qtr3PqtdnGXY6+OKG4etUzBVRcP4Gk1
WgX8mivyALfU3d1sEM+mjQJYn7uNDY2S1JMYzrB/HQhzvYDS3jZ0l6kqeCUZWD3h
PfWCT4aIuvJKn7cUUvWqgCkGdNol1kWATwQD3brL4+AGxyZORB8OPH8tPyHeucF5
TE0/1r43cYTgI7lj8ZxBF8itcRu9V3W1xkjA9wZTzoKzH9g1SynZ1oF+V5IGAAPu
CPX8YQPE5P+jIjscbDmBcm8cOWyOL/nn0IYrv0MzQEgBDhFbMGLEaur9Ljm/XX7y
yKt3xnx2tWZDA21lhrd3TZNWBfwqojHNq7YuEbyHXCHHN2rCAekQOMd/OLGujIdk
Q34a0KB+IAi2sbwqVukZ8XgIYl4KQGuSGP1y/X67tKx1++6rW/SqZZmmf1hjqHW3
VeGG4Uwj/E1Ufl67NGE1yTrdt5oriUBknVWowKFGGLJXPSOHiC6a8pzDrJkdvbQN
xcRfZrBGMKK8FB8dWWtDF6ozKpZ5hoUzIZY7Bb0q5ddFjOls7agtF756zg0SCRxN
vTOL8qZOrHbhGj/iMCg0V74E55Ts79gYlQp+0vi4HBjcZ3RWdHalnmYy04b/1r0h
HVajQxlrqU6x6LwcRqtW+3Feb9C/QGMjZgbq8+5mPPs58stANQK3fpWaqRtGU8TP
JO+jWP68XxmXr/rDAZp8BlHgaLNqUYdNgbrZebRtwNAClETzpQdkQ3d6ga2kGPqB
dUokYpCA0ivOCKNpXEPQmauWnYsRIHk/2MQF0AnbS3LEBZe64QWW2L3IsOEU3rs9
zAw7Z8pipYMzQV3mDXCMXQEMz03rORJPGdt4ZqThZSPGZ6qtOCHzM5jhMX9udZWk
e+aS9RuMamg0tymKSx7GjW767v3zJCKBXanKqbnh1cYnMBQo7vwHxfNWFVC2S1Gl
gyDPdhkh9tqxfCT1O2MWhMa+k9w1cOa0KmOUvNlHR/EoWiLrgpmgkfKzsHdp9c+R
7L2zqapfy83rwS6bLwp+Z7BvuAycu+DsSmWcdyCcrDdLwYuGgMaHzvsJwIBJp+io
oBWPOM0JyB1loeGriYlcUPbJu4NRYMc2cxxqLE6qfEUJo+PfLRmn/vWR30uWIfHn
oEocLf3Q1n23HUKmp+DsMg42tqy7lRlCN+jf+E3ONVaS+JEdBj6yxn3KfCUNyrJT
yI1zxYFBKk9tSoggkX8aPgGpTAyu9pnSrC8Skw7j0gkgdvULy+kqZlzdWsAxjClv
0NVNU4HE/MahqtlpRECwPlXoV8WhlMxbEAe3Xq1YZmhYdZADO6yzgGuKL84c4pjj
jVu6mGlB3i3WKSDUrZAqaXP05inhsj/MDr2QJRl9Id/Hn0QTBh4+RJn/fflmzUS9
xTxUrLDNvFSDgyfwyUjYdDEzBzEhpmMvjl/Fr+aESPPPhntoC+yeMHuwszrd8WiZ
bgYi6VcamKyQlI5JKzwzDwiN5Cd3UWPhx7eHO1TyQu6M7xW8si7WO08wYDYPU0xm
65yQqRbUxkUIHYsseWuuqzfz9sPRf7Dqq/cElcV0VXo2zFD6hNIGZ2ZbPVTvWmLC
RfF26m9f+2l6GI+tXS3it6Butl8rUCxyoebgcrhrMbnN0nlhk5B1gTHGQc3OdICj
+nKdpIw9+W7e/iyLeQmExX91QZ1wBNrZ4oby2iB22NHtsM+FWI51UBdb2qPPuRKe
jM5Ev6BIvNJp8FSxvY/rkp1NxVDUpvUmk+WORLLZaNHsHXeo51wPy4vcK24ud6iH
iHykRB+WCUB+xTxn5DEdgWWhRVoxTU0rpBIH2VMu412EsAQWsi0lwJe5HhUwYwze
vyGNViSBim9gocFsWIX+wpMCK9ajouClA8QeBbtlqm2CcAI+uV8ivcMJUbnBsJnt
MJArCyDANmTIAyrVYUIw3JHPnLK5Km8rWgjb6wz9MY3UqA29QMV/Z9Js8sCh+EQQ
YDOBwjzVJ1ux5tc8c39GilJqwJGZ274NwpDMf0lsCsSbdaymgV/ZDHFKF5tOEg4f
Y99k7W8591x6j89BSY6YDq/vs7MC4ONUbhbJ1JMAMGodMaH3tSKI7miEDuhOSyw0
7PCw0PrCXmGqjwKjEjdeqj3P8nXYgeODiZJnNHhNhgGwC2xU2ZMeA1zvhWhE0wgy
vwqfjT+SkNlJEyLj0SN+OwsamflCgv5YDcjH3uuj3tIRSAQRrBJjn7/RFNW9GweV
qmVSnn9rHBRxjCVlm9JAhQFVhnkNy0uf2lBaDqHNBGaOxtOKJEn7A2RZIy5BWBrY
whfbHlMVMpXkC1n5pDbdSmzlKX4CoQNjwFfRLzEj/XhzcXBVU4Lph7qJeaQaqQMg
7ZKd6z67SQVKr8CxT1cxlllDzuI0pbEEgkx49ow65KqIoZ+TMQPoiWprSqLQzbJG
z01WrrRPkrRAkvwA28GttrFSZDgCE2WAoSWM/x3OlmHG4MpxkQj6jRqq8EypEyfH
nYvhjJRRm+B5QZT6+e6lY3yxwyChJFp0ZDeqxCfn6lkhGkc0URAyANDQ4bHEu21O
vBDKdWuBBTCLfpjbJEkJEObGRAzB529i9Fkr7cmiWTB7jV96qQXbwLcvOEgTPPNV
2OzIKJH/lqh10JsjSKzc1VDRp27FsUih1jgBQAtpoTqCTe34kMQCy2qn1F+69WaH
zzzbHzsycrvlemsYqphDcxCejeBzi+PPyvWrj3Ppae3VfM5aWy0nwqqry5RPQZp8
a10BH3dVnflXlQ+T9W5OnYNPueL0py45iQ/QitJ6NC1J7YK7EUAAPwruDlg5cMgK
lBxQDvpkm3rTg6blXISTdiJ0A79PX4r2jkS3fOIhw97F65Kg/Hh8HmJCtCFk0JbV
OGoOQ8aIBWBV/hGrXPdKW6D5Gm3ANPmAUmFswDoHMfleOh27OB6v7exMnB/Pbh9A
8g9U48tfBUajecnv6WfG/g0WoyZfepJGcP3qTrWiFv+Xv2Qr7eGVJhF80u2Wn0ca
UzPNizNyfO+V4+PHNUIkwvaVQHg+7Xiw/J1VNVRgPRAqAeLr/HaqS2IsvAwY1OPm
haN2cligQ5W49OM8gOA00hghHy/7V3C51ZL6eYroPCknP680XFdVJt8tX4Gp7NNA
g0ICnssHeb3UHt0Hr8P+Vazrcr61ezspTd0ZzI/j1xp+aZiPCtg5COeZpJiVoRcA
3TDspNTXvZGEnLSFOUZajuqkCI8CMhZGUPY6Qk/ZEYUb7kIJzf9r+I20vLN9S6Pd
K6766UfvKTcWo9u9mC71sS47JRgeXsQAozVnoMEbnq/EAwfHPL9I+jP694+VtTI4
y72Hf9btZv+hLgxQEEKkjL3FKVJDO7ANaaMqIuOV3bZMf77xGWAmWsAwYcP4ShtM
ht3OvFw7XsJDgd0zfRrN1q04A2EWrg9zyx8IJJLazwVv6QQof5hc4SKpxLe64fLb
eBP0aTqDCujxWqzobL+oEvfrgAPAGAkwQnl2lZlyRNy9Yf5O4H9Q+pDrT3OyQsiH
aJd4UuguEz4B6bXEWY/Q7Tji1uyxYVaqMUy4zu3+fXP+7usorToGMyK4XnLhmx9L
bRZcilaxAAx2P7GPl9nC0N1oyvv/3n2cxtxzxMkhd/9Nw7gHPo/TU0eXCVS7kwcp
7Fq1mDW38D8YmPKaRug+cqhZwjZaUam8TQzrhLs9K0EG5joYMEJzYPTrtSxJl2U8
OoaPdtj5Ql1aVHQ6H/o0MNAmk0NiNg9VqSLF9YBC5KtklxNLEWd1Or7YbMFG6BeE
mBWLUV7fFz/4o/8o/kPfu2AbqIxTSRUqs8AgjELY5nIy3RrytM/Op8CpsBlIpw+w
DI+DtwaWq44aNhV9HJjLP8EyvumswwDWQOyUPYgnKKdjTQLd/NaRdnEr/vj0VgZX
vaYL7QXp8oaAP/mSehlkHEAohVrtKeXVM2w0XMEGrgXObjoQCE0YtFuJakfybJdS
KloJdNeZ+poebEtfg6mqlTMJbkoqebAHjm1/imwTP4o7g/WhjIES1Hz+onM42E+r
ADSzt7INhOQR9roRI7HNHUdlOCt454QaFQX/eN2kUPmyhcJotfv8IObh/msW1vSE
8eXUEicZ2BDVBQna4WHGbcxIVhZxOsE1OIQ++TR2Yeb0SQMUbQGHhqRVN0tN3t5S
jgzr9+2BiD00J0iTUhu3qOAOUv6IK6+s5zvtqlbRmqXczmLr5Cgf/aWmAc0k0Ein
KphxRc0qwChm5YBjNsHhFS4JoGc/w0CG8G+q7a2pkG27uhxwLw7UxK38jeA2r6eN
X8EHLwHW9imcqNXDN21ugi6Zy3qOsHwggJjXmxkezXIp30pq8TmCJNYmUVqDdUw8
mvGiRjsk6KFJcOnvekrm1gmwdmbIC+I4gEcs+sQc+IOiDyvbjD7W7KaCseCZWJfw
RqoBBEbK+rs3CHmO0fagvbDd/Dwyi5G35mrSViqk3n6tTJmEd0JkG1anwzz2WYCY
CTGIWey5uCpEsworqOXVefxpxolnzN5dsvjz8JOT4Hv31kY7ORw+H2CNx8qo4aEF
Erxd/e9n6tOpskKUEcWp3s/d1ujwq/YttfedpIJB4IWAEgvVGA1GBctSn2vlCHHF
z/B0bCBRGMv93LjBP4aeAEq21obZNVzfQw7J3dQlHjdgyuHxH6gGl6KZHAeTPdeX
7bE+/oMPVbZ+UtuoEnn3z8PpMLzWjlyPi/8osHRq03sZIIuPhN151Ky7jpWmS6wv
jqJSW1rEHVAu06Ovv51ILUInJ/+Ig2K2ufBF04zStkTjtGeGmYVtVno+cAqIRlNf
cxx8hOY58Z3PfDE2jGk5mcznLrph0j42Dp+O+u6055plEllE+dwvdmVqPw5A3Aqm
kG9TkAqCM8yne5yex6rk8Xg1ctzRalLzpP0NP5btv0FUMRu4NrbIdxgyY0NuMkbb
r1GdAsd1/bCUO7M0Tzfk49w5j82kfJBLs04r20F6w311rlA72lLkKLyHYhNH/stY
uOs2aFtotJ/FtXQzZ4VUArZ2mBdpQSANf4OSDmrFcZBP1mTwAcLM1rNOWhV+oJl5
OOBlBXU6oQKGSVQ7MxWP5jPwkPfizSOYriuxmUwrPplclXEfv4T1M8+94MFZw8Fc
YgavlSOtURYph+txutaXjFXpBa1oJ3dsm7RyeaD+qjM2PsaLqT7QkZjSKK1L2XOK
6G8Sm/NDAq3JBnVOAgTLT2IaYyY95tv2MP0fg6ZU0X5umJP7X38UB3GUhnfNFfm7
JVuLoVWGFSg7b4WAg7E0jtRA9N+aBMluVzOTvQab7opp6lZL5CkRSVR2EhQ7iluQ
IxGEHDngfethIZZmx9l3yKiGfW95/ZL4T416I8YBqmFqlwkB/pp8t9FYSQToQ8Cd
AzfAMaMTQOu4zltoABQgURir5BwXUjQ4sNIEdoaGZ1tz1peJtvndvrl/zSQ3FRsG
O7DEF4kecXF75TJ18CARAz7U03VFV6EM9oULFXBoR77Vb0fMWCMh3o3ziWK6RUDg
7FKdF6dx4QGduhQi8DTv/PQHZIFJvWFjMbtPzbvV9qqPeRRa9r0SYWOH7xauSOeA
Jn612O/hO8eL+uRlIaLrNOS7npgC9IZ2CVA/CD2MxeEWAoXze0QaR/DCvnmm1dYX
ldRTCVJO+xioHMsRFzzb0KSiAaDgWbXREdkIPYuZnK1AGkUkSg/w1xn0Wlu2i7LV
P1omgHEkOi1eEPuNVLkt3Spyj0htWQ5wPCOTl4cPRD2Fi9kEEod4Pb0GVCx9Z4nx
PfFCWDvmKEsibW93RPHkkwtoGMkiYgdHyRW5OcDFrNXtT0wF2PzuhzPOBIWp8GqH
r+6dj+npwRaEXqnJc2WoEvjJXSV5gGvHVULWOA7j+Fd5ro34HOIx3N0pykbf3EOz
clC42Xu1evvXo9kt0EoDhC64zREynepfeWufyaKKEF/6cvODNtuCd/zouZVlbj8I
5VjpRompR3R81QCrlnclsVlDTSWIzraQIhOaIxBKsThcuIqZmySFT5OAdsHkydJO
u6uY0iU38Bv5M5K0t38/79agJsORQ8j0QbykFlImiNyfMI2kyY73Y2UGki7FZZIc
9AJWjsDapnWybrO5qqriQbzBwAFUdJh7veJk0cWuXYQwfQcCdRF1DwtQ5SoVXxdS
wVekzpK1er54uHgWHjh4mtVFjW1eOkgBaZcPFlvD3FiTN1GW/5f7K6m5Vs2wtuLD
lJoob9rOCHuLehLWlNgUCxojMhQIAEW2bWOIfE2v/T+UAlbQijrV8rgiC5sXqy7R
H/qr+KYjp6okPD6HdRdWi3HAxf6pAyPUKY92JoQ3mSFhaU+cHno/tdwKgxpq2Q5z
PdvWH1xvPviTBUg5yCerGKgD3yPg9NWT/MZ+pa+iW+hU5rQCg9e+Lf0numxuPlVK
JvMhMqJBdQI0nYYYohBmOZ3ryLu17pPYQJ5aK7VQUPVU8lgDJkUBZwgph5RKMXXf
AJeucWIPgQmDjq6und/l4vXHxzX4uooGasbAJDQf+YMHutr+Uuc/RcslGM21RfB4
tP0YCiHF5aK7Z5AJcso3AU20Mi2Q4C5KNpXsBEcrOH+gtjWg3IawYE7jcs9ui/NT
zA5Z54ozL2GJh70mGvdaprQJXxrnk7ztCC91bn0njcVzSnd88Sg0l7UIRsqONsob
Yk6mIy6eKbBm67isqJH7idJybIvI/N8djXT8O8f2YJlb3Bn9aG0+ZVXTh/Va0UpS
VxUmYvTiwLF8olaoJZPOwpL4glOysysGKOwT9XMYEnJRkAotY58KRhWdNR6Fi/j5
epMfJ8TXQmh9+5rq9B0TIsqWQJg0s6iSggz8sWeDWf2zAspwEfrAcqdlyXWhEV2d
6En2KrXXALIy395flJAH6XwQvIVYHkCsxuQyYnpuYlk6YJHqqTze4d0cZR4HLw6C
jDt09bFNOSAu4UV9dMwMu+Vtzo0W5iITyaXhnrk6A37IMZ+aSoqr/esDAahSD8/L
tvo0VkW7dGLqvCEAXIfHJN7aUYhKT3SeEspLjTaNaz+8uxH4zfeIjaRvQOHm3TY1
IQ7W5VSXyUz3F9ucNvjmsrsysUYfv02ge/QMvoTiy2gGW2TVePryrd5vsODMCg/P
0czXitWRpTnLmkSprSiglPiwmeKC05/bEqq4gL8EWJLlwApEfSyIpbLTj+qrck+u
lHUJT99YCyMnB7jN6FD9FeAsM2Y3p4BsTdX9luDyHCV0Nq4uF+wmCfYKmvYkQDI/
Yv9yLh38jkGMy4XQWj4xY6VZ8jpp+I3Sbbzmk1jXrD3wmV4ultpF2T495xB6Eivw
EwbhbCViL8ecZ5kevbYobDlY3kZUY1pCY2zHj6Q2sZdA+ynvhRtMTvZ/dqOdnT5x
EhcUqihzHvPoNRbtJtXI5Aj5BS+POiFVpEkusg56eco++T8ct3PG83Xoky80jkZm
T1DFrBxMfF3PlEwspm3kjxLJ9irkEuTAJemgCNx23VUd1bYDR27L1nVrD+O2S8UQ
44xoMkc6Er25iL6+buvY3Z74QVsZNiV/B1ERTqIIuf0tlRRljnUqz97zHBT1Aelm
xOa3YxEfcvzfkUqHBxA2vr5XymJU9GolC8p49Bp+gmoWjUK6WZeEWJzPosqVNerq
J8p18W+9EBeqWe8c6P7TMfrM6+1/YoYmX+1XO2OUYnXoY2yMbzMMftrBkBexlNZV
6F9FaIVdL5NKQMpo2pDrgdTKKAKwklc2Akl77RYP1R2BtrUweiyP42WouNFxL8BH
TdIymCI6g/mxKoqojoq4ScxDeaFBS4ahiWtAr0XLAKKi95+S28AEfbuUzZ0+tcaI
CtceIHJCedVblhd5ZijSDYOrIjdzFmylgP58KSGJRi2hW8UkRlT8mi+kP9PRd0Gm
ZugB3oZBhnTAO7DCZVqpTq8dIKyvDgnfTKQE0n5UJl9gc0G6LGuDuEouLaD9CEyq
ynbPyrNXdhVqCN4zCrUKmGIuc96usekZXcmWNgvWeCVf7BGNjOgPf2wOdVCQcJTN
1ccNulP6N14EbD4chMxN60eh1rTCFpUDo6GGUHVBXFqP7a4SnxX+16KhX2RN+DLA
3ID5h5fDjBZyj7qRq65/Tjv4r2RYUK9Rwv/QrQNn8ZdHf8zSyrjRbhabUG763nIr
MrzUAE0Ko0ct198KJXVpLCE2cCK58DqObbOWZuNdnXUNb9nlKqKc7YNhelPD+GC4
XuGk4AoMVUFJApKa5JeACrZRUw6WONAkecnQ9/Hay7jgaY5AcqiuINaX20Vkm78K
aEiTMcPzi/5KQAwoAnjyXl+6PktkYsBimHadeo25P6euhtRKFzZxFhgoeSXgWjz4
JlxJ3bo8JclkP8FV+bi7uYovFXfn+pVixxhSyB6rUEPo0XE8SgpSY6A5iXB2XpJf
aoEsFGzYmVnwIoKTgOLKgds7/nD54GR8vsepyCwTs9rCOc6AdiT61eFHjFl6cGPt
GEfSvMBHzhpFCEqPbnbblC84RhweeNoX2zvTApXfAmmB+4KGUiH9HlEgITyCnwS4
nXeM9+MLmU19H8f56Uke4I4Cv5EjprJncYIZpRvHgTrrciRDEwxcDRD6uXvH3aDV
vGJ616eU3q2FL/dPr9+F96DjkQk1lPhcoXy7kojxIqms7TVqnLoN1IGIxb9L8N9Z
qB5FNTRQBgJcdZl1iTFOBPjdt4hC+n3ORaDt5Ju3CZ+3ZGmuseRFMNqFeSXCmAH/
tiKxHjHt8Hq17FaQ6upwUcC/GL1258GBiAfbiky+8tbvjbmAf2/bzY3A4gVzMcU0
E6xv7XxKsBMsxJ4hJas9Nl4VtZ8G7ICsqu6BYd0RarnkHC4h/7dMVh4fKAngmdqe
0VyJtvsYC9NWrp2uqWLjFg9shQpdXGOW6CR46cgqJwzQFyah0Ao8RWhGXaQe8nRd
EklqdtVvWmjEetCPygyiqJDEi3SDR67jpb+Yg/wuIEQt/qVAqtbMANMRJFMKhSha
AuEJm6wnMYN6CYfCfEO0f8iMRsQl1Vc9cMl9uGiLS7xyO9uNKI+qoNoMgCagD1Wl
hYW/vmGBXSg6e5BnwEe8W/3Z73Lcex8aUhAIFZDBYVzD1y6ixU8j8+Tck0iLE0g2
At06Y9FDU7oFXCpwF4qg4PumxlB/aXlbyR3KXjYvnk4Is5VTikkpJ2qd9ajW9yrD
ugznpxVRyeP9DUS4jtjqAGKH8rB66ppQ/002LbnaCBb7boVw+ymSFiKbFNRp2Ivm
M2wNSmewgr4y4KrM+CHKEv+zjR8I9K4kCdeUH5h7rOI5A9AIADLeddPYTwYgrJ3q
pKBns10UqxklxZvC9C2e29iONOkF5U8hoxHyPvwx0iqHQQFqPdpXjPcn+FChrsIu
e05qy0vQ7hnUddtOg/Za06i3fFfXowzwhGoeHBNNo+BZJ1ngUTYDqUm4DLabv875
OnEPSCLwXd95HXFQ3x4Pfq0KgNVFvahOeYK9O2ahmdzGOyKsECZBsGc3GbHgNMAh
QOv1Q2a7f3S2LSg3qyczuYzrsPREQSEi0VMy6lyxWd3VgJ8JPUHKJZ/uqlwpmLLE
eS14udqlEaa3Iffhlxu9thWCRzrgZhue1QNDOxxz4Pe08sh5WG661SoNDPHwjkSl
ioGtoPLrg8qXjrSD7z0d9YjcMfg9OEIHJ/Gpxs3ceD4wHBx8REN7W8sauh0kZmvJ
BKGa3sR9/PJsPfxw4HLPw1Gy5uA9W+x553/tUUabxYdnGJ+PScwInT++IQvU6o8U
0Q5XAp/O2+8/exuQkvd3E5B0OysVg6YmgYiH2ubBWync7SBv8zvM7sJlEq5HzYUW
ngfP2iSyLtd+jR80QicZ4u97N0TKp9RdPv3oxQXbnYW44ASHZ/8ecIYDwQwQLMSt
xu96OjNJhnww8AB5FlCf8oUoEkz0PyWJrf8EtuX52SdFbeVREnpFuQOzHRs85W3y
wZPu9QANKW864thWkbOa3EwZXeH/oKdmZX5LbjSgrCq62PBDcAHQBvnKmV81IJ5E
sHJwa8DcYz5iHiKA4yu9T6fpWZ6rcqouXDMWK5KC7xfARX38pl8u5V5aFsXINmej
l71jGlGTUXmmx++wZpDV7OA7i+Fl10sbcZ2CTGVS3MUBEBDrnusjWuvfPOc0nAYj
Vn4kjt8cTZ3jphTPSMwR7HwZeh/498jXbmQDl1kGnva7q52WDVCfUgfCBHpp+Bbk
ZLfWHSOqSrPcX+T+/TXAFNZtmF6ozvY8EV2VMViWDGQSp5sNYKjmWzYiWRtPG16S
codbYR69nJsfSGizNkNeNR5ClCf/YbzV2S/qTW3kgnK15dzKA5GVIARRCsEzJsXZ
34kYoNK9nFIVxsQCB2QTLZ1paeo5c5uCrKyCHmypoRtVpemrr+C1OkK9sdA42MxR
HR5L1aOUR6qVbiF6lDY4Yx/S6DxtEhqJ/ra4Ox5qIDUm5jeyXod/QWhzPBQiVeUo
EsT64o8ClyyOPEc/ZrpqPwxGMgXonEpEs0TK7jYfXx/OqR9fCjYV8jgOJ7iSWYIO
0Gz2Wx/ihB//y5BoEDmzG8Dal8tTXe2Pza9lOmSwXqU3BjvWB8q4aiQkOAtAaH5y
q4/B3d1nZXG1Eia6Oc3YjSWNst+5KIs/VPwdgZjFyxJf1yi5GBXOOs9T1ZiUg+ws
Fr7Xvq+OkfK0spOzdmoee71S0Sj9JBC30Hfh4lfzarfyAtTph6cbtRXKgbevcV8N
MTm70ZFpCY0HIbhrDNhLMLcHD3qThiZCZDUqYntUOY/ATFngWRBPL356j6QD9yai
nuT9jqxcsUyTxl0wXE2o1Lj4sGZOCEwMAk5qPhJYFQU9LWGanIyz/TDunW7V7cGM
XLGjytRGWd+EmoPNcavejk+MGpLsmj+BKP5xMLnKzAZhm6hrtl4ufTU7zhcvUz9K
Rs/ppm6xrksOlaSJPEGnP9QIMsctW0EENjd3xOc25Mzn7ZqV1AxCkmRb7zxn5KQC
9Q9e1qImGHr+at53AD/3psP+QlIfUmh08eocJFYEFNkFRHptau8sMaIBbVOToPgb
NSqcYtKtf019cFmhYPS9LGkDK/YHhhsE+n6f45jPiQEMTO5ka94F9/VTptKc6ga8
Cxv/I60Y8pk45c8OEgp0pdHeUhzTD001HTZDG5l8zAgUnY/9zCCY34L5l/BByiaf
U4HBkmav+1s65gAleg5gX2r8/8+maMv1vRmDMdILcOMovzkwcYXQAur0sgNbXrAT
i3rVILPKRYqQBuiIbNBDH+oZWLTaXJdgLvAbtDfBkHr/aa5tlyo/l150GiCIdYlC
UIrnVhNbRTtAGFz1FWNQY/QFGHxFqjNP9UFyiTs8J376lpvlSS/jun0itHgYNBsw
0iZfbTsrRbUh2By7qQyVFfzgR/JbyAzRZzf90E7LpFTazpgAuNJVC5QxCFCgHSVn
wCwbEGakTkCRJ93Lx2L6qzD+ui1OztOwSA9PwUdRKve8augyh6XGc/TRrzTUCgvR
+GpbJQfbC1dEn+VaWMHcpzxW2n2gRxnDZq9TEZgXjA3L3sTmzcc/z/+gs3LYjzJK
WTfAohLzM1Mk4CFyJ6rCBrzFAC3xZOU7/IM7n+7OF8qsAMp60LsHM9VvojvDj7DD
kbKexf+3FQkPzxgH8YKAfXyvN43mq5QCiMk0Z0ImwmV2rnAOobGTK3howFl1CRfi
Ht5zo3Mt8sL8otY67RwqAEjxG/uMUL7qxMooGdHxq1VPL8ogf2uu7AnOeqXWi+D8
f0ereSnzZXqjj2xBONoDFquInad5RihjO/P/ROESJDf1nYCFE+QjkOynzM/TyqXQ
MhlKot06b/1STXPmDWNYrydTjy17OJ+BatS2PMVYCG8nsPjCCTH1w8vUvIOgewCK
DLtNfJcaYTYGsFdgKzWvJX58oIOZkPqLQOx4qCVjZsR00EWXliTjAGbYZrMl7gWK
tCSNOK1RD99+c7R8Hj1MrBPrKgZGv8FhjhKK5q5hNLHVC1EoQwiybz6dT9uG/CuC
s3o6gk3hVIFKo1d+HmVdEICIL0U4adgUpCObRSDLsjqPZvdNIb1uSzYR4r4AZGqd
Vxm3Toso5XObxY0Tccjw55//gG9l04uNWCAmRTw41p6tQlvfYybGPf0oAGo4sVGI
Gk7x9wGfVKC85m6oxBuw4OnbjsV2OsNX5L25jySLnmP5BhGz41JhlzPWJxXfHVjI
p0X/UP1w+WhAe4qw8L828S4Rwbn/MVtjTvASRTe8odlkSwFUV/2uJTw8hr2lxt1F
mQQ+c0FmYHGdp2s8Z+tr5Xqgc9ONb0ZP0qRs+ly80RoE4IuVBGwhaGLcbm1KIfIU
xEqSdujdW/6xMZgEgrs1ucHdvhmQ6IioGPoSuRDyq4T2CAE1EvGpgUyHVWeqFyzi
ceteBRpIjQjm3UGDDDX23rDbwNMiknDhl5gXASGytKiqsskO8tZxruwUqgAGrbhb
5bRXFVRoM0gOsPr3n74AV712RiWpJ1RmkrHny7u9LKWynocGlD0XYyvhnc01T4/j
gILas4fw8AGWLUieTCNzOhulE+ZMeHlJXctl2dJxCzj27+//nGzsD0sM21RWmI0p
PSmWccP4XkUdUicEMu8ZeNlIX3sfgXnnghdp9y/ex1OcuHnEgZ4gw/C1P03y5gpd
DrNj6oHGFM/DeaNRBOLQ8Ew3+rpi4yRo+53dHOzmOAzgQwSnOe4uzsWbdj6NSVm5
E7MktaKR9YYf15SSwl8YQl8Nw868Vv9rVh8qOMBX9G4FCVdWsywE0J7vRsydS6se
NP2ahW3uEYFurKk3oXh3n8ctjSswt/6IL+ayNHdfgeRusONzUQYFuQ5Sj90Unnhb
1Ug8XZg1g5Rz4hNDBJtVxIZqFxCFXgYDIVCGXGTovgy56UqC/s41yGOtwnHBQ/ZZ
q3Ye6mhBgCc6uS/FrakIMQ1WepzV4izUSbCD02fFtrVA/9Bw1cs57Rz/umuYgger
s+O0Hl0a732evITG9Hxb/yzaHgu4UnQsE/SV5hlu7SQvzuBlcxyp0DuTxWynTGq3
uxNVIlax7LxaJTYFx2Rb1HfYgU3tIhpBzLiMpPyvkke8arpivt3WYe4fC6IcCwmH
smDGh5uwnP3pLnE6kOo/gMllSGalURoIvw7D3R1BI2QruVCRQu1Z5a+ZXzhmTmNc
DEyT+ZH9yDtbkl/X8ITtlCp8Mj4OvY1wN3c2ra42M8hc+t/Tt9rVloZ8eOKVc7UP
85jb/zPYSrn9Wg+uDVEdRgA285bps+BIW/Slx5wy+pqqb0dBsGtmMCFGJ4SRQnbt
TcdCxgqPhHyc7pYvQ2jDQ5XvLnz8VcQ7iTYR4ToUm9WUPkYGMYLxeOD9eZlyY5zU
AI0tPgXujg5jhizsPMctRkfNbVkNbl4TWgJMW0nm74grCQ5CxWGWTOdnfRLIlR5L
PMuyP7JpBGJXvUE4E2jLyOXjInoC03KmJSibkrYEMdDCF2fye1Q/BSX7zTyhqrx3
f5cZFsWANSCLEk9NH3fCsnXAfDZxLfTk70knx9clWr8TWbh19c/WBgfSiGFa6cfc
92N2SuSgnqyuMTmTkcP9OqJewmWe7W8bGcaxXZ35OsGmLgRvjUWOkmi5FKMU8zuF
6jZZ0Jaqgva0JllG5iKUZJX4VK0MBMAR8yg0yQkCIT/2bN8l6hXEbnuIgNaGHGOl
2G97xqZ25u/GaukfhKWHXIhnWw0DJnU5050+aGkJDoeMx0OD6XrSInJvhut4aYoi
exiuwM0NxsI3LG4ry8iRgJ9jzNSKx1kPtv8RG4aa2BQw8zhzJP8ZjTNBRUfWHDK5
TAlCVeBSlim9EMdxl08CRmTbh36TmcfH6cGq8nDGfwpZ5850yvDMFxnUnY6LwI+2
NfSmnIpY+GW3/puVd8rLkJ5LitqZLtnTenFp7Fx/TaTrDYC6JWmy9R1b9JcBcgA0
yy6MtW01gsCV4NusRbQaQqQ1rmbNUS9X3xQtIIN7R0CUt5h1pHJSuf7FCqnTDifU
XxV5evVhEXl301XVtkUysGrkmMDWv5TmEIG63rx3GiTbUkkNh68mhMtOtd6mEhmH
ElEEwhPtotsoFKxF2oT2P+B70MZNITr/zDEkIO7EQqzgkq3wKyaCOKmVGGboSUPD
SbXv0KLs6I928EEJrZj+qH6RxdCXSle44PrlpIYx5W3KZF8OltBUy95SCC1w2E3n
XNyVi8DHo2iavXEzCCBQ8iCha6vnAPDDWNwMUBfhaG9/5A2eFCHvIF8UBouZRzd/
JMywZ9xnYhZ+LjOlDze5ZLHPwAFdLO5tDdAysvxgHEKNaFwG7Fm6yTm7GbMX/roG
bJhSVuzNTi9FGShrKN67/MEZ1MSG/1Yu/hBDS4XDRHSa0sekFS3ed4PufvC/wF4S
WIxV4cxdWqO09mpocxvXmH1g2pD5YKK8SShVCC/y9zDzk1oCUr6ZQhNXuNGhhiZK
Gb5F7fADr2biqvCrcszXa2heoSN6+Pcdfnj3J/15e4MJj6REowXMqKCS5uKxG+3z
izjENC4K7OXusAsmoHahnitgbgopV94VtWaW5QqTbOCinR1rHAiTTp5+hotTIAjV
O59DSIjn7MXejH5ZyBne4J1/uvxBQ22+Wbn3HsAqai2LtUA13XF6FIZxvhtnCeJB
5HSzqC0sECdEIPhstuuhcWVlJer/LVEiXGnRZUk7fGcuK1nCtXfDrPGjfLPuZfJh
l7EpiX+uAsTeTW7DgFsPRQBfIunbnBwZoMzOf/3E4TmzXwbegTNhSjYudtX3oyaY
ec0DY6y5EhzkiqSfUKumHE9jTOISAgwBk+6I5AhfEdYDsxWqK56+hVUBPZPPbHzh
A97pfMnALljGXFZF/NLAgYSuYKaV55mXYuANzjxelKzp0ZMnY1zB4DJr/GTWVO1Z
wuBYKqozg90TlFXL04lbWk0UQfTD5+2LylJk8MBbT2n1LeSKwj9UazVkb7qnit85
2D4zAZEJE6dsjImfZe+aFqwyl3DWOSamBArNSJkhHwSBQkLSgfQ0flhllmd5oLOL
A1/yx6U7ctYuoC38cNs59t9/Wnlxjqfeae14uMN3W3naa8mXcFqgJ8tWguS8Besl
iKsyf6xndO7WrD+vcDaDA8oZkEWshoOBgMh7utfb7nlh11TyFz3bJdQRSok5ioTi
eP/1k8wKvxbx8rjCuNzUa5EvQ1Ykh55/diz3DjjNIEdeS9v3UcQVLFifsmGa/Vqp
21WRljUuwrx4Mxbwnuxh7xutfwG8u9eofm7NBJg/zCsZap8MFMOMO8fnZ5y1Yrdp
ky1EHOvY31IFEwxq3NlUC/ehtlsqVuQzGflBFMTZ3/OR4+tvnIXyqtLlkQJpfFZ/
34S604BGehyjSIEqgJGNwZXj8TOyTeKPxk4IygZrSkx+3P7R5eUvVuBC5p0Oydop
DpUf8BsGFx7CivIK55J3KSQSjSAV52trUZCnv2cFmVD94A0pfAO5ZLqdEORRGq28
bBA79gyVvTQvbUCeWrs3Aoot6oKTc3HFH94ZZJ4znStqI5GYTf2VRlD1IEojLMBx
qbH5wlqLIoxoJmeb2whEsrEZNvOtyJJk+ezD1EPKBqxnMaTKQbDphLMG+dnrR0n9
qLMB02cvSfovKmN+cJn8kZdwUNZeaVmxExDoUTVp/ouot9BtBUiku6WysrGjPEcK
p3/E8l+xLCpleurPeEwxhH+tZqfr7s+4oxeI7MYz+0PCQqa3sqtvFElwsLjKQrnn
FLlwPBHKRZyIOBrOoeOIaULznc7XyvNPtIATZMTjdM1M+KG1fA4ahEAr93euom+h
lGMGH0ZHvNXQewafU3tCkgISOINPQSLEa/O9lG/O6LvkDr33HfcfKpP9gr12Pmbd
UWK6zHxaVYnnd2xutxWb8S/3IfMwv/UU1IlGz4DX2nMLRVgdBERLBf67JtMJZi1D
dP0D8ws+wr43dFBebIzYnhZx8Y7A6vqjVfBCZwPuVp4D/z0kY5IRtmP0LLmgOVWa
C+w93vv/s9O5Gm+yCSR2WNXLKVIJIDNq+mbjOK3qEyq2u+/2ZlW65C10xopdH5qm
bCWVAu3730lQUupFcOlgaTPhiF1e5I3iTBUSbKxayFnC68udZhuNKfgC5Tv6m2LZ
R4pGk677jnRa14KJ51J3l0ZLITuT+pA911hYr3xPFSRcWdC+K0hAbtIEsTLJ97kg
+GvClqNyC7OuxmC3KUY4VROn8AOzunjBKUakEc5evZlVhgJ/DcIH5qY/hV5YHOwY
yPOR5a5M1eVGiyTe3Kqf3QmJcCQllxFKO3old5NPJ1pOrep8t6zh1IVkq+sGkO6l
5vnu/QRhyJ2fZJEu5vuSifCYeGnOyemD+GUn/LKwL+uHzxvN8xNPnEJbmztKOSW0
2TaJIdkBglVe04+8vTVchkwONzu41gKFRBCNpUu8VV3e+LGPmfA8tvVzoKZFaG6C
yFBEcBwogjDqCrhUHg6oy2dvHg2nosWjn/eUZ2H6If7953zl2nEhqOOzDZXCq6ac
4pHm36AiHD5fr56/pDMhKb5y17Fs8XkE9H6alVQAUCasUOmNECmPMCC0FhcdsYsc
jT2h5JS5mHCWqxhyLaG3o56l/Ae7rm3EjNQCeyG33XnTK7sWA0ewXF/bN3o9MYxs
YnBWdLapi/WTVyWTyS4Gqtz4PW9Op/S22eJDnw0hSZ63jlD86xQcbKICSWlkCHah
pQs9J3GTQW23i7/pbW1gY7X6GOzlE4kMwio5Jcnz9sL+CYSxqnkFSQwfrlRJ+TZ4
tIwhdO47sa+TPrUn87DIF6q5IrIA8OvVX7mN8q8TyzeOQ1GnE5e10F5yk8puA2q+
EzI3fWgPCl3Tz51j7NJXrt70/89QvKUcU9hJOuiYvCSZvxHyeELoeS7CDUMOkB9k
oYTOwBmjKXL7WWojksZG6Ik4jJF5UvsdkaGqNIxjBFbXt3SWZjjeuFvQi9w0Ylde
3j5QzAzT9wkhrbXv3+nvyC7faPOC4owT05KOPb5Em8Hz25TADF69ZjrGp+ns/0oV
UTxUTNiz0SBae3SDD+OxLFiOxElaHpXY7rvKUokumJGK48+2pAZNSHfcI6wdlbg5
op4+3Q3VBRgjB1bDR5vAfc4Lia3FYReyh7YbsrvngocaQSBhVrdr3xg/tF+wg6VB
DMJ/MIsvd7obMhXCxTcGNt56433/6G9mlqOxIlhV+r8qGUvIijDZz7RsNWW2VeGl
lqHFlnrYNh2HnwZ5LaUnIxm1bpaCL4hXQvaNQaa60Pl1Yc1PH9wTlT1qu1hd7BXY
quaKg1LIqNC8QZVlqjnYv87kXVIVbm4+1A35o7jdGc8cvAB+sZ9CrPOnibfnpfNd
/mgyLJVuSNQe+fIJ2xywczGyoMm85EVQpul7K/7lzq9OX4RRdsGdNCLCH1qzNQPT
CB1vShVjGgCuQUtXlF7XhrATB3qcgTEwStbXWoV6nFepgIcea8PGGbYudJakLjyu
POydOWYEx/3d8NeQgn2c16RZ3xjH+zCSBjfpOKZ57JMy/KGzl/fdCl4U6NzCzeIM
JtMCuTUwTYFuNTOS3TjAsJWezNRdl1+8iSFjEVTp5QbckKWAWYQu2nNEdjzVmE+O
CahE++S4Af6IQhHc5f+qi+VIj2Gv1cSboEGlA6TBb8fc6nRKZE6ck/84u/J+LhMV
Bvwt3eij8jkzinoXAT+Slb1fBwI+lpgTC0NhbT/KXXt/bVC85/Li84Zv/w/Hb6jr
op8qI9Eg216wsvPH/z/4xmbLiCeuHij939atk9BUsd9EFrqFCTT2ng2MzjDcSCS5
ALe3QKBK9jk0tjqP8kxc457tVen0hZGtERQ8TSOid7FIquG+Vzju6bBeGbaBODhX
zAOLyYKm21TYo/mZ59a0toNYsJR4192Jgu+6PKHi/SH0y5fjRqNz8GS4RCDPJjeg
F0d+R2utUPyI2MxTH3WFXrGlQg7ZScO5Ic7N3Zh51FzA3XQKP4mqPpgBZjMcSNxU
CvY6lNQ3SJzIahj0+wSpEdc1yUp3R5XCnERaNX4JJ9aDTg8VDb4gASsWmXqDOe05
Yy6BzMnsgw15BGILDrQq9srGw+BGgbdzdEcwxKjYjeS9wl24MOb2HcdCq5d8marz
zZwHeOh0Hwz01CIIBQ0h7HvpGeWUoelmsggVoJBUeai4W2P9QRMLLu2U5yBrUpsy
9Rq/G+oKOPAHpJ0YyEDtpsGvN8lEkWIblVXPlUdztDgYLOc42qjefXuWkJlruyWj
gwXF9bJYdWRIk47kzBifI6KYxsFuofKmSxRoMN9ODawufNl/CvttsOvlHod8Oqlw
w42xv8Weu2PZ5xvYoTaRV5XOFUqUAm1YDKVbLHmK+tv7lZPqKC4nDT3C6ZPeia0F
hI7Q6cTfj0/3+3j5NthJB5uhXmaBwGB2upZdVWopVKM7uR7zTApodiup5G5l1cch
XRMfrSVlGVw8+F8s83AbYAPTuG0tX8KQk/E6z45X0jGQ7Gw0EQDQnjpic57C9yZl
kG8acAapVmiIjEUh0nl+f4DLGNx/Nh6RWO3nR8D0VwzeRTvnmA772wQF++3FmavK
/TCYED2DFASwnyCpSYhCy8rQltMMw6pDcPm8VFQwFwI1MEZz4TR0p7jgyk0IQNUS
7AGhCXDEbuYEOcjQUk+2pUfpdJUH/acfgts9O4IH9W1a2o73WxApQs6R6RKSUn8z
oTPycQOGajPlQsfgO/88/1M5ptFh/WmuIWJWO+tyxW8vtXm5VmNFREr/hSb46iS0
oreXcVdLfsTog/hE65x+7pF4SiYHmCQRGG1a7R9gUvpAdpKy/Tyr7KAu6X3B4GQl
RPKEpdlpD7/eJdn/yRTHbhIMspiez2GZ1ov91jXi0u57BxrXK+4PBsE7pJ+2nmT0
a/bYCyimyO9LBC1picpLtF8xhfnM8C5zMDzaZ5cu6cfCcwrW6ouoNAUaPJn+Lw7Z
ptnRXN1lDYED4M6QPlABfvlURg/WpSNcthdk5wS8y+uOPv/ArH0eK+1PWzQjX3pJ
qGmcvCvS20sxGDP2DTiY4vaRPLtr+LnitvdxPbT7NhzB6LmmxxsYvkXYqs84Q7G+
Q+Io1oH0jwXCGBExoFsE/3gz4kLhMP1CgF1iQmTBLjpjezgRCiDESSAfPa3DdEdD
Ac9JBVnSiM6n03sB2WUDiHCdXy58wjnQTuHNfnlIqTFz6+dlmCD2b0tZQgSfDGkC
cz72LOqEyy3VWqkAPN7mbrgieGC3PFbDnOtXK6BxuqbIOM3ReMFabeTT/4wQ7QRu
+Ex1KB4ZEHa2GDA7b51IoR7ifbcsjSrEkkJ/NHLMk7RvD6VPV3fOie8GD7FeZQW/
mbWmrbx7gE8dgSA6V3T/xtewelWfCvHX9f9Ws5q+9lQHfVnmrEgEa/k/gxx3soNp
rL7qTGHMz/jl6bexq/gU0LikXjguYlvrToikACXWnaAn21RyoalwFIx51obOm8VQ
bgngvCRSYVG2WU22Xec42jhj6k2+l7X4dPzMayFApMGDzKogWXTBnFTUTarACP/m
uNWA9XgnntlX3qSDixOoIfJZFs+vte0S5sXuI3YIlIGxIepDWmeTX3NURdRFgxQi
RiY9aBsGVeUI0viWvq7tH3vZ64jUEr7eThz2lMYthL4AaQoeBkNxCdp1cJ9KNCqP
R3ImQXZyeJGLLcdAycxVuc/6civPsJoHRSnMDFNYWXue7j9U2GA/MJtKXHRxBRt8
jTpACxcjqzMPt4312je0Bgo98MwlFrnYG1tx78gFIlg4UacNAqJ+x164g/xk5Bm/
mwHWIs0V9xXX/1SpQV5OlugCpqY/Wp/T0wUyDMotFbq8oE6N+NBHZU8fS0hKL+uq
WTu/6zm4AooBFQ9ugB0mlZ1fr0vujhEy+KSM+0fM7Z/5TwRaaFbB1EmKIxcybJVR
mwSSaAhDXbjwprxRnlxBHkYNdBSk/Aj3ZOzAirsSmPUV+uqupHGOoDUy2h/k/GhV
lSD6crUieX+yjCC6iKYNf6Vh4XDnW2FO5Il4tpkqVmTRhZgQ9rHy70RLd/r9Zaw0
/HgqgHSAua8TYfP/U+0gfjqNq20SPXEkIbE09IYyvXOfh/dN/GUrpQpUUfbqOUrz
XPnoO2x1h4UYtrar8EihIFZt02Av341ENLVrovq9epHJFsxC6FYcWx8sAp4Q/33O
dr+Pq5L6Dsl50VEshSGIH8u0XRg7+Kb4zaxZ/f2SbmcsyXduhL2ytTx1Vq4EcMfY
g2LZIqpnwKFHvyS6Z6m98tuNESDUzsZDypYRLK83otvefC6AE/AvEPdCHp/iIg7Z
B5tm4UatVvx3XxJL868sBXAyyFAppVzCijDldSQjzlRPrhcsi7W7h4eOoajsuT2J
V/BFkZtozvPcbp43vWKjaWrGr3aV9q9g1bzFxJAc7hROoxQ62lwjLIhOvIy5kxej
JmCAG9y7XmRXUJqmxBj/jz5a/FI8mak8SCFCeCiZNpDJuRCgMdPChLthvnYRSwDD
cZIWvVnVXhF1RaJ66fDjLyGc3xiUjpew6MBBZQrPNPiwi3KL4xCp8RnWiyhqOrHc
gLliZWFZa8TFA79QCTCT+yjBDKESu/kWw5kzSKx5J3l4IRCBHh2kucyfS8LlPDWa
8Ao5rBYxj6Yr8FhZR2qXl89PkQlk1YONS8C7YfMQxebRqijOXNpv0coIIKxSwJqX
WW/1pDwfho+XAooK3EE5jfqw9K4CQthDTL4Cz1psfAtqVBPjyKidiQfWkhc+7iAC
2TBdam5Zc3J5Garmyxedqdlg2VSoUdENW+j53z/w0YBJ/ARrjucQEwY0J4mqpgaJ
t4kljp6DQ4WNSlLJDeRLR0J4nnzvgY43lb0l1Om2bWxW5FVPfiCirJvXwMAR7Pyd
9jGT8U6ykxNaPjXLk9S3Ku4wgo+xeN+DX1fD4jDoYV/+ClzKqa+MrFsGu+N/8Xmf
Cr0udzfNs9UJLRexOJuxWVdkGSyhrIZ+LjDnmVLNszzq6Dg3x2R/LEIbyt/tCtN8
7hfn3pSciyp47gL4y3GKNiHkHmFfcdSArjhuGrQwc65D+Nwb5od3cTkg18GplCZg
EXAyra/OKXAmjF99D/b3yggqEPBr6icutiHz/KPPnqebJlIwuMRHEkRF2/C8u8Se
U5ctec/2xwQhGbZ7Qi8+TZr2Rfv76UrYDTvoHCUHpcfDfCHX3cwdLpb0X88DgVH2
drKrcsumUZcEmxyfjbTpFl9B5DYM9PDY97IvRSqrQH3nwjYYQYcrsfAP/+kZf8Je
QpJC13cd8n68zWoUKrVR+6fzFGegHb9aPp0r+nmpVOOU6onBykknrmwxBuiIkn7i
fcM9vkc49wDX80DzRjMhpVw5QqdAjCPcuvLwZLXXPRSQ5UoSSF6fW3KteVsqCxfY
sTTewfvQ81bXMzUGqdegTFBk/iVwecaiUatZJ99YphMKZOBv1HxIBj38ejYUgPIN
Y8h3ZwrK0HJHcoVtwFMT1P6f/FUuHbD59VE/2caJmlhmhnN3eCt9E7rOPtf4FRwn
rsgaZBUYajjsEdLw7NJaykqg2eMjyqs2E1anwB0UBCZf67NFNtN0UJGPY4RDASLa
tivhmOJK5tsaJaAK9PsEfan+r29kqgzDYRVt6nMrNppTYbLIHR3Jjqe3iyqWDjZF
uPc9Zkm9AFdPIiV/xfdlh71c43b+JFDgR3sbMY6/l0MQdfsJRqdWzKIGLz5RgrYi
Mj4W0d5Wez10V65c2twklXjZgb5tWKFGAkMriD+1Sf0OWnJMJQH+qni/Iz4G/Wqn
fFxWbcjekUGskm911JL9mP48MsxGt4EvLeGkHqf30QBCMnonZeiaars6AFWcnuLE
waBAnkKCs4QoGTjZJlPXdOIPJ+q65MbebNIB4HDrovIk7/T/YWGwU31FdklU2+lk
Sjzx1o/htZ/h8bGMM2LjNC+eRyiXPI4IMkQChWdzy0XPiZRueXJDs8HLyd6ypcSL
2Kuk6C3yRxaRtts/GlcdMOuU6QREaTHm6McgzYNw/YLJIUlNdGnr9YoEO67PvFH6
F2qsbgvAX1OP7Y5iVWGPbagapfJjXEcLfkhuftjvEfYd/PA52SsTY/Do/f2ZI5J+
yKNjZuZ00OGS6LGnZWEMPnYOzmbMwmvCDviK0kWkc36wGUWLgqvKFuTCtOaX4jZi
KC8dDJWiSvNvn12LID/LiebVmRFlvft//YdmLfXdLM4ynDCxTS33ESuyARFZ/ijp
mrrq3QrDcpAisKJ7c6wK22p5yY01O3UE0paEjCeT67MxzcOjgghQe111IeJXa2EH
HlUSPiNNjhuBHuL8CQuTurXYYroMLaXf4phQOB/Ha6I8LI0HfST7ko7JGh1geu/7
fKCVywbfFZ0jcpPBcJGmxBze3iRiQryXSKGRrL0yKBKwuKFzx1WGhtmJvGs4aN+G
pvMJSzgBzCUp7h+mM4gjBToIe3EpSeKh40mB9+B5oAL7r/lD9BMPXq4ijqoT7XWa
nBAY7oLHmZrr70BJddiQjxeMs3VxUJn2eblnWUilXKUjZOT9DymwGKy0qCQ/qnxS
du/PrPMj/RKRDiMLJjyNLQvURJg0DbwjebbmxZl9gWHxpyA9OFsSKsvqyPE8pNft
7mSAde5RC9nWAoXkZk7T30UIOdlYAKiIRHk/Uh5Ej1LpN3WIfE34IEJWVtqhe68R
ASUbfvEK4j9WwEJTvyldhaCtcJp0N44cy+jWJ3wNr6aNh3wOsdBza+TV9RzTpt/h
qj3gOxJITeZ91W5GFJM5pNjbypJr1RcGv5u2A9G6MCosdRUFewmSWt117OvNwTPa
+fgvuHHXBMz0Aj32TgI5cEBpw7qjqkkzvrsJgtIEZBxq5eR5qIw2uER2DP8ab86o
pFdH95jAU1NnH3855j0bIKcXI6gk7EpzNXqm0CusEEZkH0tFzvUUQRgFlPp+kvqK
q+yBW+Sh13SBZrjd+xCsQa9N5EFywnfszNVPadg8Vh0XlP9ajPn7qp9t4vCNCi/p
lH+NItfriLR2Sa8HYIPsKETV6bEKmmxwJJCOC5bRD/u2HrccQ5ZiB/sGPJYn7Jae
YLm1Ze+58bZaWbQvZtkJLwBmy9mLqnyIQFUlV7z6j4+7dcF3aUNwdwJ0Wo+iq2D5
4SaVyKkGLSa7SFrRWpvIOTzZfHDlOVl9kVT10f/9aWWFiJ3wpkXQQnAEaQ0cmDkx
EoAmQJeiFkHBKrXEN/llA417WPny/031zYPutpUPV0Z0L6vcv125CpM1yXQNH+SK
mzGboZAX4VtBbK8hUnNHZEokSsIwSgMsHDqFiKREy53uSa2o1bfT2tQ3q0LMoNa0
88GJ0VfIm8sPdLyrvjqWVVEAnEvcE1wrFm5HN2mTDXhBlgYLvG7Q+DtBMH4Hn3bt
SY1TXiJHk3KxwfYOeW/sQvgH49JQGewnKZq8EOD4rdCIJWTgKa0xFU/fP/fmMFjV
v/DUFvj1BevbbJGnnpWg/j4r4+8R4W1bVxRCzc2IWM3tzpYHOVaxCmHRaBKbG0SV
CVbYUKlJsEV+JOjnqMN3k0nwh3buHyk/Pk2ItDdWVcey+sBp7qimG8JysAGlPT4U
yMUrtJUMjjGCkfCMR7YApxaRaNH/lSuv8znWT9pCfkf/1Ia+0o1RpFrGuyHrt7fJ
ECLJ8MFJtcpX+sINnu5c7mqR+yl/QXIr3SF1chWYNGmL/r7i/ylKNvDaNRNoXe5E
51+rF6JA51dQoZenxrdmOn+ZT2xGx4kKRqpIb0HsIqI9o5GHmwdJWYNNsd/xaJVC
zNr92xYFVzAh956O+JI/LhyzlfUw4PJVfxfe84phWsxfqAIrKS9/CHxp81EmSGoQ
rddusqyiBB3GWHYBPr3carDSF3lvUJERwr7B3aURao8jZ47humwD9+7uOAhgE13H
llLH9qqELoLo68a1TTt8Ev6Q6+lOhY0nsZb65fUoWXGLQ6EU7DzpGHDvzx/QjvkQ
TGvMkIX8UROmgytHrJXiMo01bpoA6av8YheeS624aBs3fEomdzDcaeTfYK+AY0rj
Rvou99XE6IWpw1Rcnvb9f7iXthkRdeaUWKJ//ZPI7Lj4RT1CWXIXurvlnPgWX3Mm
/NxduVtYoO/Fmmw+9KUQdZHFgPQbQ9BEXemLjWK5fSb3isQk3ugbMKrOxskqvRl2
cU/D5Z6EBIwDII3jh1jL8gN96hPzuv3RXSoLLKenlNktWVyrqe/5aGqSrVUjAaC0
exAhGBXRjC1fRAjMjKLi6GWVkO8av3lhkKPY8mly5sAVQwH43ciP1o7PSJBJPqRB
5xV/Smum2JuiSDmc765DyI0l4SlygfcumbHIxC9OkR1UmoDbSB4nHRzz9TsqlCHR
fDkbfaBPY5Ds6fEHMDLWRJYfe2GATPpzNGd8phRAqb9GVuAjliWnsp7mXIsTR2+D
Ym0l6EpN8GNFXmFDjOU9Zpe7u7TDuUn/UtpTqjtHcERglcvCCdXl3shVVHRflzdv
twI/s/QRs0F9IJXjS/fv7oufXQpi9ehczre2jWG4CKC4pF8bNPLjyC3ZYv5+WPYS
ULftr94E5GyHtGREjVEr/HV2IL1V+GSjAwr7HokMKDxGnY+2DnX6d1BxT3oEK2T0
IhDDV+nPZoS89Bf0dP/lXQDex6NoxYEWHZz2rcCNMPpv9eAuwgNxFmpR2rwf8omL
DvicE7V4+WpjAq7PWmWLWcmzNxMaQlMzFRHT+KAlbnThvng3qPp7TY1Tw18HfU67
e+jtrU5ETLc3ei+CNDCP+/bhL3qDgubzg/bTGs/Keokd/8smWwTUmc7Hhew4yIqb
G3Yh+RPaGGWcxyPqtH9FEaky0LVz/XF1HOCdDUQur48IujqXar59McKu4+KISzbw
nJ9eVqjhEnc0G6jMy/2oq87Q+Cj4EMBwsp2LDdE1aVnNQBMYwTtTCaEl4kiCYWZO
b2IFtNBa/mgl28qugKCpHMoUw6Z+xuebICwf4QTEB/8YpceriBLcdMiZCI3Ki7BA
76LIAI/mK7A5g61Ke2PVAw+dY37OzX/tJ0n0R6f1hBsRi6zzXwsE6KIGSmZZa1Vc
YmFa1JocVM5W9C85xM+/EXLLj40udmsp0L3ftcBQVbJZOQSjolRAMndk+XFDaimt
gT50kiM1oYKVR+HNQAU1CjX/nU9HdDeVX15tuXx26k9q0xfjh4wnYbid3NPb6v+j
dDYPFzXujxtsm3AMA3rfn62Iqiu88RAHg0IciuLLh26AjD5CAuJWtoWbqtp4BtQ8
+9PtDQC7wWVyQ/X9asn9TsM/xZm7v7McXC8Yne4NQmhkcieQ4PiGtN0wPpqFprkr
Ah24T9GoIspfjGNkkFHid/Lx4a2+C0bFI/ytlfiiAmipbs523W+RFWUxPqt/0S05
kpj1QfFxXwq55DK1nOATSlcZyggiZc/5I48LzO2ILvzqE9ma1v5UH5bwDs96rvrH
qaSfzeLbjiJmbBLfBdOXHl/6tXS5xY/etTCjKszFJmfmWCJ1lS9tEG4WX3YgOuqq
GcPJ9Psuo0NsoeOtSoQH8Ke4U172cnABjS+8PF/mRPsXqIVUbKmEVRYmvZy2O2XS
U3mfMidN7RZ725sSysb/4Bpz3cFIg87UOjDC3fUhlN6yMf8Hl2cxSF7HrHe74i9A
OeHhULaH3MWDyEeN087+acqyCjSr1f+nhWd1mmQ/3LBlmCkSae3Xt+dtWzuYt08v
rXNXq8n9htNKwtDvae2yqf4YkPF5gkwhgICQvOCcCnzJGj6Sc5fNuCDG3thSfrxe
sswadWqNBIcpHZfzCvoS2EIKGhuCHnkWt8Rvb8PSsXB/fK5bTVobUHPDzjBAH5eY
vQypnJE9ceiQtdeIBn1xSoBedzxygw0BNL/6AmPmamzpgWbf2uMKGGNJd8tyuN+U
VRRK9BcSkYtvr/btRdX8vzBt6hkzEdqJSxJzNQ6yzgtvWKz3Cp+eZpfblP8/O21W
6/dEJwxc8lOnUQIXjVP+mYc64cuPPsqqjOzlye8ZrMDilvvVyO29Nugb5iTTa9dq
46I6O7UeCaaCdDZf7yWDRuttSw+LVTm+PVM+7daZTjD/EoefS8rx4GXfxu81ZNkQ
LR/YpSRAjK93jw0pu2adtsjjcp1V/c8YPmfnXMoHemf/GnRuRSGPhuDYg+IVlRVk
lDZR88MLGp4mgr8mLdhmfeJPJvoB181HawZMaTzHsX7yYroWV8rO8yTEYLbGjf21
ZJt4FRRHY1iuzU/R/k1/fT2RZkXmbZpYuUsqcQI6Q2RJCTCIFlwMb1/KF+4BjATc
al7XfI0DNTNfr7yCkXkeSMTXud3bp5OpA1eHhKI9rl5w0aeLmjKsD/27+BxC8dcn
1l2GOnfxx9xRDEOnfdD2TJ98Qs/eaSReUCc6uvZd8zbPUB4Dbiaw6nZuHJdKbQHT
x6vDt9AqKmj90FKAqH8y1KPNarzP8T7doUl5XDZMc4Uci5Wnmh/F/gb7NSRHeMYC
moKiK6gSiWAPksF3al2zqz8mxCadowWxw9m9SYrKseLWEmHnVi/osodg1ZoPyAq9
xm1GLWvh6BgEmCz+TkzGRg0iJHCiJEjrtsRM4aib9LwqR/PFmxDVACrS6Dd84Nfu
Gd6cSjhM+9JmyirrzfI2vMSaTZ0Ql3CHbgZTJbtWYKWY0WirBRPv6kzw3ep0zkhI
6jWuPu5ZBt58g2z/IzPwSL8YOezp64gd13RnSGRwOTKxasNa1KQhIkC9jr9rxAu1
mqHXmMAtAdaA3q5ovJ4uiebqR0tUUKY2E5uJX7LVfl9Wekum4c8j5CVGmX6dlK1a
agLG871pyWkaMm4AYDvsRIMb2LENOCs4KSjUANxaE2dgVTGQG9BOyWfv0dAayRqN
6t+VePqVqYzyhs8btD1//4BcND5RzDaK2D/qiP72EK4RfK/+888s6z3VHfPVf/9x
poO8OMCX4osGNh8BWEzQOIutHZt7qoqUCGyd5YbKmYYmfUHEYw/xPGui562GIK+R
Ie420gK7eD7rTebVWgM/kX47nTVQergj96GefNpsgcxU3KH5nDnFk9w5F3tz01hT
yyoStHJaJykFBLjNO99NwDjZXImJzewFAgwlxC403bHGCfc5PNTCgwa5+hVfJ6Tf
DDoGsSMCW3Ezx8ztkSPuJtGV52ilHW9Sa5UsbnpH7cgFpY7izp9WDBdS/sLJr++8
xb0QKgJvYHpCuMVBudTQoVB4tmkTNa9P0MMahj35qm33R40XwRvgdR8pt//hVecL
CHfvMSPIt0O1b0JTC6rYCsXB/2au4X6wtw4/OnLri5DNEzKo2y3Hslttr9GdQ5Md
y0jm2F9Nlv4XCgQMTr2771nJ/IyerdZOi06R7VSqGQ3gT09ZuGldp090q6RPN5HG
hCPU/XBpxGnHt+tHtHeO7eC792N4MEVZAg7AoE7X/UxvE22Of/0Wzc+5Q4LpcbAr
McFzU08nRYtI/7pUWu3Ew8zwyVPSZPyLyr6Iy8OJ1Qu3Ed8ci3awFtFqpH8VZg9m
qujHyE4jiK/ZWA6zGyRBXgkL35uvE0L25euWc8hSpuISqZ/oTuK/oHpA3vc3ws8d
TU43ZsCBgLnIeGkSsgA0HF7S0ZKEFK9PB00v6JPM1Rm4RfgLeeEfjez1x9nqLzwb
F1xPaKFgtQnF4jq1w20jiQMhGsp2ooEd38JPUdWle11B+WCPiRCW0awnqyd+hfx5
n3gX4K/Zs+KYrrU7rES0naK24OY4uhblvUC+W7Kp1wZmgDXTE1PoN7KtYrtiUllp
V23pOnvldwNUf1IvmhrcaTLTw7ZvNTrQ0kuOvZK2Gce/MgC8Fep0n7fVi9ILsIh3
y62jrQaKLS2bwdlx6DzQqhyJT0R3y9AXUXMl1WQQ3ph7e00Ncri9KREvmIeIZpWr
G3XFo6ze+IPQEjme1HCsKjUdEEvF8uX/LRd1IMZNAQjJWLFEuiG3ggDm38Gg32df
RxKYIzkcQPFLOV/CKDIqNq7xQM9zB7iQ6UaSnG1/GyQDwst6YGaddfjGoyFuf32b
KI2Bc4NshB22C4oyusYZuk4VqsAgRSQ7SXXmobn6VZMX4XFZv1XsgVH2lb1rNaz0
TF5CoBsnvl6NrosW1yK2+RoGo5QwastOloLAUDc6RrXSTm8SUTD/uwXcLoY6l6mW
/rJvshlFeq25JYwSyKqL3N3mL0+Jp0z+77OvUlu38iPQIZ2oojz98GX+0ibtJLiT
E0lSNsCKq3KXSfUjIta0oEs9gS7yK48646yi2BqxYmotwydgYgtSg/isM61uEN2n
CHC4oGJXlsVfzJGjylyPFX66ZsuKyFbM3lXMj//AocAX/IhA93AzsEzDWohVTJQs
Ge9NEr5IppTQAgUKnOZtaYKK/1vT2whDS8yVpdlRNYhshrtlObFSnlo0mlY2yZ2C
rW0ye/l1K15+yzqs1Qyzq8dWkbE4ESyCHocj1vEWe/wydNh4YYkgLkY87SkTgxjv
Qpf5c624xBBC7GtOc2F0j0U18j19vFgBuYD13RNRBy13ApzBW8kdKik84edjQr3m
z3gY1OZjk44PKTMMEqfHebO4pTeOqpNlQvtLBXzeaMuGSMGeiELuwStmYFVE2YUY
siYqyE8RE8bLnk7bTP4NhWeX1Y2K3CBkbz1lcpGJ1Kzi8xTzUU4VFubS/w+eOxfZ
+h03Ao+tIdXKPH3aex6UwDxGU7jd/o5jWUiQqwLM4jOZ5hi0IKeG+FONArZV5sCd
CkoCFH4XHWlW87gjrEwDkpUwOpEZzlp01OQ0guqeotpHb9Cf/WWtqlma3XmUHx9a
iZ+3ji3Y4D0ORRN7BYxhRXOMECps6IHr2Eb2Jj6vmf/Hqg5snDbpbLXF4XQtbt9U
lNxw2Zr9WKWsl4k4PhBeTCRuRdKxRTq6tW49g9PvBAH47Yymf3TZQnaX7F18ChrB
9LbWblSIJFv5cTkcI5YdFIpzMWb8bu2KU148eRV5mZ8sI1Fr2zln+EW5nCPWQ+b4
Pqc8QTMksKjete8A37MobizO6/ykwY3OaSJi2xfhgrGXrXW+9FKE8pbXQIlbW288
0bHLr2KIbtkZpgO7hVOWTFZX+H4jOVzJbPGCIfokXCpyj95G9zT/vKCR+mROlQ6Z
Hw9vf9caHVs/SzM1RRrtpkMXDmYr3dkl8GneHj5TtUoAHzm52RVIwZHdtuIYFBnQ
UTFAIM8cAApQ+GKeS9wkrI6/OhRUKXEjaT9eEEPZhu4Ta4pnnVXRoh4xes0mAIU5
rLrzSXCXBvhjuWfPMQlx/zAieQQ7qxVJF+HySnFyC/EiWg8+nVU8Fwu4l2ApNM+Z
m6X55QfGiT4mEjwonAsC05ng3IC10Iot57VsNUePzejmjtfZcNdN+2zuQHQaBGJj
mQPPXUoE59Tjd4/LM/+q7UaNEiw8G7CS1x7/VJWVimJlgLU7Np4ffWcWqhPwML73
ywUUxwdZw0xDTEpSroBRcXAY7xNMloFA09y/Ubo8WFy3wahpzrkn+X9cItSkMaL9
cilw8pkVhVjIFSqxfUzfNFn3cOkVw7WifMdYHe25yVCZ9ojE6yjQJZBZolWgYmMN
FfjNOLvcXPiQt5Wtq9nG69hPv9a5Cu2ah2k1VGHnldV0R6vKnw1NeF4uWU/Pm+F0
yAFBCK2cln+ETVTBssi2UA6OdoMNd7KBX/jrTJfrhBxVotTVyJv34LtDf7p6gLoj
DyJEJ/LWCiVK62drzvpDfd1HU22mha5XDaA6jrg9eEL4pG9RbOEqGbRVhHgjyrqU
lTEmVyqeD9Pbk9ognGaJfDTSPruM98HH4SkulGJRtOqFk4qC3bOAkuDGZx+PAWYc
13iBIHfypKJ6aDSzZeeVyBfYSHn/dlcW4vt+BZHicH7Se0ZWAMitRxxhKQydzSCg
tUe4bB3W9hkn5Wk1jKzVkzb2kTImKTVahtC48tgNKYOiO+hYNVk8GydJuTVErj9M
e/HiOoQxVzdIH15Q89p0ll5atDfQaGkw7FE8wlxlGKtknCy27R4LGdSZzfsnIRPg
OH/laxCPlN1fopnrB2BM2ZU/WIl2kUTrZIj1MNgqJTWPPpmEai+54vj0Gk5uhlKv
GiPKDSDy1zH7A0jDrrb9WzV8T53M4Lai5reXXDxn5RSqLPdtB/eqg3VVnMTREH34
3tWCaI/Vlt3bigXTwIJnqeKcB5kzy0NRwOkoPL5caCN7ifApN2+21Zj2RsUR5ELv
g1dU3m4NpYedc/SZHaZevDuasI+WG+EQd2iH//ltgTLzdacfwpHKHJkMnds8S6HQ
4WJIgHYhCK3K8e/rSLFRS1WiYBorK9Tm8AuG9Swpwg4ANYaQzKv43bbiU00aim2L
GK4smRofxVAv+RXpKTCH8/q5P3+UWAeAgrQhLJi2gXIB7PnR8q7eJQGND4Ua4daD
lNmCLxEEFxH5lkc/bIgj2jkLdd7apXOWzA4sVUROpA3UBYv+1ItT1XGRghitqj6/
B8ixFdDwMrAfJoWv2RlX4uSRGYguEjjIU8OzxtIjLdK2SDERwGX3SS8NcJfV5sag
C8NcdB/FtGx9gMGVurzx0y4i3lpGUh8gX4lfzQog7FAyJngKDOU2pTWbdcxmvm9d
5yABmtP1mNoVrH5/r3wqPdFlTaOFmKyBGd6J0DOVKc0WqB8UH4Mok+Ni19Pmp4MP
A2e8l4rKxkYtph0HTGIICAE5c8/feVGHR+//c4Un9b2h98YF3H91LsTs9+kh7Nks
38cGmjGbux8iGmaurSKuccqT1jdWFG1GytjUDDQv2QN6jIdrRF/fBx1S5ujxs5n3
3j6L7XcbOMiEJtZxJTs4PoUP8IjyWBCuYUtPgVdNocdZy2iMmhD9XKyrwHGnLqgG
XJJrsqwvhb3uV+SetrtKARS5Kxwz/2OrsCR3lpjVPNWncqUfmx3Uo64UkCb2L5og
XQw7wr2OFJIDcew5eBtca61ciK6HJTek9jrf6IrqfifLZJr4yeTPMZP/9KxrgKXU
jn95O8+pjLBNZowXP3BBN8g/Dkl1iSzdIOjVJT8T1Hk4vBiPexZLWAvCvichRIoO
r/z83wOv4++IDuxw92QC9jbUahD0FcMnygry0csoutEJNQi/Sous9ksJdRtT4W4X
eq4F0PH6O4EEtXT/NOK3sbtVufAO5Zc6+es4Yf7HSPZFxp9LoHerPAxv8+zIqG6F
nk843U3xlfrrNZm/h+u5GaaziAXVD+7TUTDPhTzYywcN1mdT+lXTl4Tem9t3TU/6
NzsKUcD3iVjYGlxzcRZK6Y2t8I4pQgEHHsRUJg3z9BR4/MTBoyumH0ZR8jvDnIrJ
SR9sLvGlz2LhZYyKzt2tyvw+VrLWcmI89+lYR7FqVVO0E6tLsvp/fVpfoK7wPAvO
ByEB49vxEl2QB0fmvpk17Pmx46JMSJ4vzS7+mantg6yyvvCnp6rW0rcnNOeng/PT
NhmS2gIaPWRLGAQ/qClr8wX/e/GR3WQ/SGd3g5ugtSgJ37lmMN/3H1jtLZeTkqFy
YFncBdRlA+Z+mY1T7OuB6htTMzMAkoaqyd3uknoM+FRPigtDPXYiFIPmxgMXE6nB
t+cPvtxCalwJlIHpV+LmZWRiyeXh07jN4wSrc+Dl5wUpqADzndSsKR2mKM7bdyN1
/RN0f9bH5uPukY8n0r6vrh6krmL3AcbM2McyddkSc39Th35jw/r6tPzyX4EkzJcz
7kWN9manbeyhMDVJsqso8kKhOGJei4nqSRt0YVw48ugYsWcXnUEJg/LVkQ/qR75S
TxUMi74X7Gf3MfrHc01ZE/5htPTqPhgpWSWenOKGJx7hNO+zVzu0KNuqdRz/SIxJ
+oKMUNd1S4rNVxTVjJf+vc2nBDBvZ/ls55WJV3qzIN14BtWE80DgzgyvKy7p8Rsg
1QZrv890uDIjYlG0p44bNVLwVoQZdw8/NOL72cKvA0pAn0E++kQ/Gu92WACzGYjs
26daANbBkp9xXdsvj0yv1LeE//+DDB2sTe/B8AKjsV82aJf9nUhpiZIc5BUCINpl
r8bdvoBk6DYeby17KIc03uHYjpk1JftlIpSUGFlehhUiYsQntQhFE61cMrNUDS+y
rpSqbWUVhVJbgZW4Z7Osm14EFE4DfmnfVVJ6jJkfn8VDC59guhyfKQjK5DqpAZ3f
xX0GIiWoNgg1L1lWH4druP91//GypCafWWywcv1diw02V4oRD5HNC65Mf0/T0w2Y
KhyJ+VQJ3QAIr845af9DOWcATeZFX/4W5vSlwJKXNuypNjkqnKnusTzqM+xfshqg
+X02qwRAPzdCkwuQwwmXgsJB3/l4L29KTp27cMYh5odz4nRNkrb7Qir+jH3PyLmU
9HiIIJim3H1wSC48lmaDMXD74BHkvaeyoaJ0ZaAkcLoJDnH3j9I2YNMMhbBs9GC0
n49V0QzaNULTS325LQRCEHqDGK+9ivolUgBWCiQWqh/yrsgN2G+zSqjKOeR91D3c
unbUfab36I50x4cfzOXyVrJDfZf4CD4V+VlIW+IxMUygUuKUR2LJ8fJGUhPg6TbH
sgtia+OqbXmeuBNaGTb7fqcwFmPdZApvAJppWsaEvWsZtSKQP/m4Jq/0Bx32Kcav
HS3dCFWAMeboUcbZelm855v73e/6SH/w/veNcmoEgQnpAtU/zyjsowDg/DD0dDh+
zHMryiFhzIEBbd8IGUC98sfULX/eO6vFLgpSRmqEzP6cYe7nxfpKbrZD7byj5Thq
VhWt2hZacD9QMRCXNFeh00EuIGyH1nYHSGV/vuoU2+ywRNUWkOxNdkTgK+LQAXKw
wDckkiJDTDqG1u3dAhErqDHVoT+jEn/yCIUZh2oftAG7J6vm89KUBik81Wvfvxn7
YaEfQb7cNIqGne+vIzDboWcDSWGAQUUfb0QbhhqZ6rz29OGnkhRzeRqL0XP4AeO0
unDqt/s9SdtK+K4KpYEnFL8uly8knB2NTWX5MXdBQYhvGLvoupI7tOR5FK3kGvij
UGGxbeogactl1Dzixs1D/WNZkk72/FQ348KyvbIVUn6StyjOJLOeNkpjsN/E6OXh
C75XAzyVj8YQ/8fJj02aU+Rmry+/ES0r/EMFCtnxIDH6jqV6i0npxAvfOtz8kwK4
yp8ZuEVXT2JvpUQTPAi3elz3qaxVd/bTrGvOzN7OtfJzNT3KPhRJY0NwbnPlVkk/
VOarG41/qLp979MtJr1VpjvKd5my7k7urpg1JBAv98M9HkZcx8k0Mv6bO0Y2eQhB
e2zqEHv+QIqTg8dFySDTY/lR7T6g5gf7vo5zPXl2A9f6y1Ly1n7LWvjJWQ1VLF8S
nrZGNOedOmWktTZEsSHMnUDZGIjJvVnUmyFn0RUGov8o6T7ytwI8qXorUD/fr5A/
fa1uT0txa7dnpVctdKgQH75m9r0kqqEOA+wmxZCKFuStXFTUivktmK6B/bYKYPHS
XR0d/3+cHHbgxW6HiDbPF72eljLIcuOAYY993hfZ8ZcnKLHszmxYMq0xloRp0Wps
p6qrTrLOQ/mpB2MHMZr0M7eb9teYU1vvyctzac/CEnnZSBOcUBjvjvKrC2+ZRo8P
bKRSNOlR8XV9M02BBbw80ObJEaHX6/yHrhLXmWtvTTEpLtwA67YyBWNR/9T073b9
1jV+nn3ngp2vuy+k3eKv7cvvC2JkXVA6xvtrXgbarLR0grwX844hoEk4H5ohtG7w
Dx0jMsyR4O5277Nlpw7dmC+pFe88pRrE9mlGY63HjkcVmGyV+sa649H4WkLQxLnm
uZS7s+xrolDtCbmDnHp6bhJU4T0IexieqWKXSdMmrW2H1poE0AdBP4Vdr0eAGohF
ZlffkOcAX50O+LZBEcKpTpgG6hgkWLFsESj5aMavxsOgggR1CAHPaWGqeYYnxSVG
BCeneySPw+yi0pHbK4K2eUvXhN6igx20imHOujFRT2SHok3guuQYL/TNFsoLmu66
OvGJ/uRxWYNbMQBRWyyWyCUHSRoAs2VqhoYHcIXP+h9FrgZoImL+yso03aZUnO/v
cYpZE6ThG4kbPK6f6ygThBXQx4S36/UgYHZGN35FZbokeLtIFlN+YPFpEIGZpwNZ
Tk+gibAbNqXP2Wp0VldIrIXw2rL4lqnSfrMRBRTdA36tA966KpDntB0tod7YcemB
JFpje0D1bRyxvne/TXfUZuLZrdN8VQbR4o9ENpBdnJqddHMawH43qc0KTX8MEjkh
lvKzUf4ArKNkHp/5nHdojLj08KMhuCCeRhCt4EEF63zU/NdnHveLy4gcuMQj7/4l
yn1/9BWF5PujCNhyiWFp31VwQNC7KCRqlw3TfDIgULv2IE9F08VbS885TPdfy3cG
HfPjh3eS0ejye71pEf2c0+jHDUfud2DLGESQHRNFRhQoa5vsmzLrUiv8mBSrSLaT
X+KwsG6BnDou/bnf0nHcWm2TqrMZAyDQVLCMjOBgE8T6GxXeEsEffwLCOWVelkAd
cm7XWUxN+E1Mmw6PXuB81K3myi4axS5rFkCdh1UIxVCWUYbJnaI9r0xijpAZTpIm
gKkOC+eWVz3lzd1gJnI9RzmId929Gr6A3pErG4FChwlBd9LDuWTRgd72eI9PIq7f
puwjXxAk3MNf0vSfHNSwrmgvSTg+2qsexstjXW4Se54SRVKk286+nUtQXXSjzIoc
77bpAtw1j0GSK6uU68FL3xdt9GDuYWpFQqioJHnP3n2HT4K/jlbkE6qoQEG25Gqi
Np2rWI2VPU7Rc/Ggn2o6I5qB+8nm9Y6DiUWD8+XnUsTz+IflbM1LnRD7PJZyCjeh
0/OvFKqOxfQyqLPAdl+zJAMEvMPcsHpDL6hnM8RSQ1cQoN8PI0jluvwtv9WL7X6z
9Eu/RsRBv85u0V3i2TW5C0qS6BNRMpE5bgemX0SndiDRSg+ocCSDcNkXYLh5tS14
GRkW3F4o3dTQOyjV9Mrm0XxSTDORGr6vF8clJGvyVcza38E9wlnkQV6djYNqeLRk
CODN3cBWeZ/4kBTWrFoOM3HkL+qYSJtkbykGn0/8LTOeJRjqXNJ4FdGoBA+Kv1V+
dzmmrSeAImRr/irer1ZO2bBMgEIhd/VhPOLqpJDIRs8g966aENv6gwBXF6qhlTOL
CHkttNhW2UHLNfxN7OLjNS5TUlP302UU++dn2wErEZwTwMopYKRyF8beGekcHVAL
R06nLZPxahFs8uJJWnOZ5YQvq8O+uDvslrrxRFsbUwkbTXwMvigFZD+vYczDuP8w
LiG+PwvITCLCXjGzXFRkxqQG6e4Rj98uu/cAjVmD0N3Fr+ihiv740cyqtOtfdML9
VPNioa+abqm/hJoVhVSCwn17httd3euhIlohNGJpiDxGb2GJf38tZgdtAAau8z/g
cnWreu1+1lppc3Ssla2sFVZqsNwaZh92JRrvDFu9PYhsw1UsN1oTp09DtGCgWR+X
6l8vp8xJncxetGc0fnfFxjYVW04P++yWGdix9MRM3yFO6GcmGQYRAchyoX8zT38A
paKrBJiZd35PtIvpc6e8Jgi+aLhDZm4nr5rAjM4nrUOIIjIm5hUkXMuNL76KAf+L
++waQTqXaHBpHUjaCK5qZy8z7TlA5pWfWo/S3PD/AKdTzKgNp3hDGpGEW/x4vNpI
ujVILs/t5sd+TUBgoKeVWkvNyWxH3qHb9knvR4ifChh5K5FquY3pOEm185o5jxsx
2d76OiA2OA1Xlq7i7vETn0ewLYauphKD598jIGPw1fNd55v4jtRTyZrgi0RxuGxF
9ya2mEmtrWraFtTuekjHBr8QpYeySoK4S21nNP6XsclF7ueg1HBWnFBytIAist5y
z8auxMmbkY6RBAwbAUgDP3nzruLgf2cLUBBTPnYcewWzqwfMrs0q+JEqE+QzWxrH
aKgQPhybntS1zmzFjTIcSyOD7lMU+YRH43J5BCzzFK0m7sPcGv1MhMiNdRNuja2z
weUzeVx4G11yhcqCgSv7cGHHSPwMirm0zy/SxA/X6DNSNzKe4ejMWzZLYw+GFz8k
Xw96w5TggepEifrvGA8xQuRsLL1roFh3Oq8rdx1Hgp5CQiKyKRoslaBvBlgwTGVl
u+p2wntCiSXat5GnR/2QsGUOEgQlu2YkJf9aHHmxQdSJdxN24ttUr6/vyoBcnzZA
eagta5H3867tbARb0elvFsxJOQlreBMpfvmoMmQMKPNTZgG690D6/oCxhxy811yE
fCMCcPSoOm+UroWf4AZA7RlB1BLZW+8BJMkKYuH5rVJ2As4QEPz+Ky0mowMQ+QyG
PSpi04auLSwbyJZ5rSd2oRKhKwxLUq+PA7o+5ggmB5UKhUJq8OSbVaAYbyTi7RV/
qEbe/WMJ5yy6RkK3A8YfDz9zrXJerbdTqxflMZczu7lsuPdQlBo/N7UjS2YutUyu
mLZ2YvpMCukbZ3YW1XCSiWv4Abgs8Ma4v0ciSMAsKRYbF/dlyQ7er9V56BHlQiGV
EBL9uUSBkSum4a+Br/2IMgmukq2ndK6k36e84D9a81UQhU/A5PjllaxF14tnz8pd
prnZTdatlcMsivsVFBt3kMUaFf0oxCGjXJ3B6q6sxpkNasas2GfnK2uD6oFl7ug7
CWpo/9n6pJtAW9OanI94AWGJ0BGl0uuzvqMMm6LJcVbLUANQ5/OtzRbKvAYJjanx
5B2ZjFE21h4tw+C8UukdAr373YOl5mfmVOstQBE1pXY/faN4mOACJVBIcbsP95m0
smYzJ1258ICMV+1nCnjWzVxgK2iGarBjBL84DpPPrKzMcZ3pPvhoqWCgaSPoFTCp
7jO5x7UdKn8MuMy3sqte5qimIW2WKQHKzwyfl5cn48GqN1QfS0Psk3+m0f6lTEa/
1+zOl5SlsvsZWM/aEXDGUi8yBhOSZfHE/aQ0o98AM5UYW7A8ubDYfxMXAibu5ohM
LiHc+IkdBVKbigYMDR5qtqCx0iO3dsNJfzpT+JbLsYUa/LLrTSIM0wkWpfmKS/gz
gPJ1pUINBfUJ2Vk6L0wxMJKbgSskh0herpYqAr0lFWMgtWDXNxjj0oJJEnEPyQal
LLh5msIr7WSJf6tc+VSnuNSvtFqWCBpf+2Ji3LcjtleAZizz3hlWmnCQ9ctAfjzy
s+ADNKrnzSFpWKvyHn8aPHtLL1LLQ7Qd6na7n/DiNUxbUjGsV49nSjf8mzEtMVEs
4vGM/6rB0pnZtGhIgScE9LOTeXBWHZc8chwvyrbv1xTzDe1tWJ+F2RurG3/oot0j
iIv12plvMn1Ck3Pvfa9Up4CrzMM0GQr1ibipdSPm7WUDP017MgicjN4nDDu4sdMM
OsvJmvEks3WDAncFuVc5XulU0QB+b6BKQ7IkbS4EdpbeBTdrq+XdbxpRbMeO+B+H
asiAOL3HCokJyrf4c71kVveWw2c+u5964pPLBxS1/uimeQC87hb34EYzaz9OVbhu
1LJg+NqxYq+z/k7d5yioehQV3KYyIsfuhPiibSLrJ9sgcrFosTDFuCkjpCqL1nRN
2kSIpoIIwiaivCuVQschUcLWTKnW8Ok18bB2P2+mXUjGlWwyFBVeC2uwn+ZuhHwE
ohcOcl+DaHc5b1zNG3OYJZGWeKr5q+JQt6HgmfZgYD0OjhWr1vPzwPrtfZY8hBxZ
eaCez7FdLlRrN2H5GFZ8GCVbcK6M/O7Aw8rs45h8HC1aIIIT8651ga6aupWRxd48
H4cpJMJ4CAXckjYScuoCAe23r47c97kXBJL1xlB5alwibhZi3/jddNDYlGuvKw6c
7N+rIaFLRoOhDbhZM40MbZ7YWtGu85tuMSkmcZ40pNwFiYAQm4EyNOHVYss3ZJ9Y
MPS6vtDomBFGR5DqvUA7vTT2n/+jCWqVzHn+TQe5nv2TIMWPJsEsGPg5uuPxYw/4
V7KzZjA+nBBWQXIe0fQER6ZsyoH89KLlxvOBiDvjYUlwVmwPug1MV+0g6Wu5lqoc
oehAA2cUfQAv3+ffiMef9viVO/hMCWEF3pkTnHyHFuLWcRAzoDL7sh1vwMaX3seP
/NN839c9lSTzOvO4IuX311qP49+QDzv2aau8wvHGJxLeaJyLN0CL71UG/sNJahOn
bKktXCAOlj4CLsEeb9/YNbfjNaaz0myXhcv7PgWFLrk3unYGNvvte+KTL9ujF4VE
9co+K7yFytgTewCGXGvUXfrbXn/P2zgqyihASQX5FvYqIZ6BKLuzk0//AvXYge3R
q/gRAuW1Tf7cNN/BhPqXnRVBVRhC+EjtZa7R5LTx+j3drB9uiSDhMhRsMnHlve/W
JlfOjPF9Sm2Pgp+msAOLffyfOU/Mpht1HBPcUJu4UtqAN1WksjHejgQhVQlqnACV
ez7E7h4be4ftFn/iCzxK+zYLtPvpYQsSjTv6mU+UbqJS3OLHIE1V1UTVW50DhT/Z
3+S+MWQnFgx86ZySgjRMvg2Lr3+JHc2DrL/wXgoU79HSeHUtgcFajSG0EhJVFJVG
Qk/DzSRc5GQK27hLhvbWftaIr7Sr9fXanC0eAyTYD/sPiBBooNICcNN6xHl9H3MJ
G+5rPFoI+6I2mMTvQ60l3ZVSoagyvHeYBzaPNrMdSXhSqmXq6e4n5o270xmXHNIk
9GZcvn+cCUMjvGTOML1tKzOu4C5aeqx7sXKe+2gkCOzG9I+yk3A2wsCWYFtt4zP2
mtRMV+y6cUs1dMB+jB2aPd80xU6uRVEKS10e2gX1oxo/nwi9hQBYjP1CFf5wZeGG
9q2RxnOZf82cq6sf92oAaFBhk9QsstzLYYJ1Cej26ghaUKqlELJW7WhOLRUPLk0U
wMrKBgR+puQyW0gQma7rJKDGdEsHlS1G7QEiLv1Tn8vbap2Cg6uJUwiDM5BQ/PaT
hMdW+NO9l77hUl6LrS6DfCkCKbxSwoHVS5sIFvC6wEBhSI2OitauPQgb2lwSuF2H
6Vz9OnjKI0RVBehaCXFeriKox/67CTn28gEFoCCRkg/fDN6XfV12QBTmj2agdx0Q
y2E8Ai8SK35AzJgmIcPKh+6r5B3Z3Gj8XAkVTFs/0ICl2e3r3ZMgTvb1cVP9Kiem
L3Ri/jbgnCTDuZcp1LSrBnMP0Rg1Kq6R8eG6U/irGKQgmRci09QriiFUOOYE0RYA
Z+Q/hULTXS9eHUsX36NenzqHgWJ29Nd7x2o38eWtfSPIDHa6n/D8fLtXkZip3fMN
+DIB0Y4SPi5U+ARzUPdBzgJFWRURkK2dE0T/R3v1WtXiDpfUOY1cRoQW3EVKMp9H
uUi/tSvECJMmBTCBowF0zL619oiedRLeFZTLaakoqapCJ4XVDRv/bp6B7XN3wbGY
nX40FZ2mB5cpmbjk3NhbpZ72wjfZNuUAqsRrAj6U3M4+8GhLonT6cojXyjuUtXZC
U0Zc7DpGb/BD/h7kRoDZZQh6ZFi4JJ+BOoqRihkQmXiE72j1z89619/RiDhGFb1a
Iuxn0zA0WNEu9v/e3/R7oKPJKRi0GztFD1WVpSS3OcLPFhUKh1it81cIBo7qpLEF
Puywm/uXpkal2bJm3ctno3J99PCksIOpPfBIjmaDim7CoWJY51wuiO4fSbBKmukC
/g9Wg6iPCGsIQ3wAbfXDwd+A2mLUCUOVhL0t41WSAjjUS/wdWoVtzlmTY0oR4KSA
w2dcMTWf+8A34UNYsqJLhnmonC/uRc6BUtqJMLCtrg+G/QGqz1dckIeRFmsGn5Uq
IEz3QsDK1IAKR714Xn8tvA2HGzO0gy8YKhNkJjw9oZ0ohh9zbn+Klzb+LKLRFmz3
JoBcjyQOKGJZvZ4grzU3lTdA9P2c7iwRxbtvecMHV8lyNdLFXNnawVehN1p6Vbz8
oV1zElI1Mnbqm8XXJ5f8nvYn8tJyh17Ik/afeVY3HZQI2xpV06t/cn7hcvcoTqZM
9UO7Sf3e9IihX4mDf3tt8/Fp243Nhr3dDtM/rx/vWUwKq8mNhzAJgbtRn47EWX1A
oDLsKFNeO9EZHlGfR7SaKrW6kwrcXDSGvneOiwyMh1HIEh2Nu4m4m/oQX/R30F/y
F+fWPsVRBkwR1RiPmSG8eMMAKnDyAC9NczLeyknOVKlTBOlJFTeTLdm5fESJOcQi
ppiSzPLS+erBWFO81iQ7eB3WmwSWGZaXATTvY97bAhIk7Aez3Itirw4u58QOOgBm
IaPcX0IRLeuigN0En1vjjGYeaLWf7eqwwB4GpDjKfL3m43MEa9ySeUF/IumrSAWe
bGV88biGbv0ZSqBUuwTgTeyLafuOQsrzYL/mWFix77Vm1Vv2x6IVwnJ7dvThVXyP
ehMqiPrkjT1SzmQ8Xe2ocSgV4EsFTNT8PDRA8Ir8qrJiCQHM2nAWB0inbSvwDbfV
xmKzgKKvh0FY97TqAAz9KrtxfQ6XNM3Ux/rEt7Gjx8EaTNX/rvoOA1XGxMxfW0VK
j3KbrbR8JxmRlD5YACmVhkK+7OG2VNJp3qiHXUSZ/Uo8ed9WF2QQydGBujmEj1gZ
Fp86e4x0NTU16vPunki4AoUquBx/ptPHDql0U86PwojXqwDP2zSiLfYYl7CE8Sx+
6WmpHwHV1i0NRG1OeuY1Yl91UFyIowVOCTz0TSjoM6ZSRXrEZjk2HybyDXF7Cuw4
DF6PDomDi1TLKhYl8+d2Ijz9eVQUgwQTI1znrl73jYJF0+/EuAP7AhyZJSmPKURG
GspI/NGH6bjiCRZSnSyNcQEJFLAWSYDeuCbToKTUfU3TGetbEGKyBltvDvkDAkP7
QlFaYL/g8UzhGANUxLIjtRPyvamqc6ulai3v3upo1MVcSnHIhbwxfLIhQ6MM/2qH
YIX8QUFZr+Y36riHOJEduhjThSbHnwNwWeeSA/Sb/SMhhlrSAPJFGF2SZ1aYYNaI
PzBVvYE7bCD5NGrVpYZRxNS4vSL0JXAs1uYDBGueNddNVFFouXBcGbjNXjYdzsjT
4dMHeSH21RMsB7hQ9sminM8wZ8ICDcT/OGkngFGtO3qCfnYAtzoc5teLud59e6wQ
V0e8mBs2TDizum3cybEUIcJ1Vmy+zLiM2XH+pmiiGN3A1uANiFuumPIpHNmP4IJ/
zPUXvKxgo4Qoo7dF0T+UWIKeLry+oo99VQmhh5lXC+iXaVDIyh00xmLP0KWc9CJo
Lvpu/Cc7rjS2l7LM935pIzQZ09KXeheh7Xm/m9TsJ47lBAeiOlq/QZKdVFhircRC
0xHkDErR9GYs9f6GjV/LTAYmtaKrDgEl2woXZg34R5ztBB3DVO1RY4rfUeGv64+f
6wH7POzthkUHUgRYidABCU3+waVo8ZeHu5XdDpqHFfk+xlzMIeY5yP6eGi6ubDL8
IKRbYCY0FK1C9Dtx+Juk9SAsGVuXINN/4/uP1ybC3FEoZ9nt7wXUFRagLWMp7TQO
Yh1fgnjs4XXeUJkrKejQfHxat/oQwwsfLZ3mI/lowq8PgOkvrn930QEeX4Wc4rOj
9wwAtbLgC14B29VR6fO1wliXlHGxxBy2GHJ+UZFQw4ECfsTZlyqxuCu6nH89WvEj
YFl8JIqEgJxWkAtnBESPbj7u+DOT8dcMC0l/hwAe5dIb88RiTyojinNbiVQt/gAA
xu6Sf+9ClO3x8qD4jwv7IgJ1QXfqsO278tOn1h8GT2QMlsCKIgLSR1JESHm2PjOW
W5BXpp5cFkqr4V7ljzBJseT13UUXN3bX3CQg4XwKolTW+a9pKni+jmciTVFEWKfM
z0HIZOAXlAVNvLzEUv3pNuu5b4+i4VMCMRk7DNTVNxMWWvM2pvjA76qBUqQtNySG
o5X5RTRIA640JKl/EAKJEbgs2jTdzVGa70uUg+17jzt/lseaYcizkYqgdS+fu5AS
iDb76lxIVpWFG81/p2NFaPlvwhctwDatsXfIGziIqEXTP+qBpck30A5sa1z95Srp
hyBdD9pm3R6WBW7IOp1Y/eZoLf14RMURWQNcRvZ/j2IytByzkYe1+Qarn+SDzdrC
QZ+50vxGfMTDIPfHWlDrLBmQHLbgH/TYR4LmA4+xZFSL8P97WOyp7nq7omnWRw5b
uMUr2hL9kaK5e4Y2iFoAgf/P74T1H9wiLHGkjtPGsAhzHDFJ/I0Yk99HUYZftQtc
XAdpdi+Xw/a0MMyM1x5Kx4dv7xKs71ykMZrGKL1rSmO9hEwz0jGXqNZ3oZsTAiJt
k17v32Fogbl96H99LaJOYz7o3KLVHND2D8/VHnaxDzegROkAMBbuzIaMYjhZ46NC
79tTpQ/i3ua5slqVlNt3ET37fBPOs7fFFv8ZC5XUSxZVmV+Shg8NLDZNmf+0hUMz
921OH6wyxAk5+1GuFyE9DG0KlzmU5g76Dd0jUT6lqjU//Vb03ObaIUVblxnOUI19
CISeWZ2GXCyij9G/oXsFqFZRAQp6LT1biH3LzpjC/9ZUjElI0WIzbgL42Vi7fFpY
GGpqjcInBip0A4zliIVwfKBeCQ9qfmnXXKQlhDL0wM8UaezrYGviXVc+TtjjcJxm
IA0xzA0jkk1dvuVW3+fqosy3AIE7cRgVJGDambJnNbu5mMLq5JrAFGOIPDsKjQud
xJym+s9/SknMEpQhdkurNtFtYuPJAL6/GulOrS5QSsK6DcGW1lfAboxAOhsff9vb
HoEGtGzFBmdg4VFKHFY2qfjx3djlnueVc1EF8aKEr1jc56CzfyZmqu3mBnf3VtR4
6lSPpApKL+JNf+n7X68lIHbcTLIb0TSE4VBtME6dMArtV+kEucOiQt/j5JJtJk+A
zeXaturFn8SscwIDKjlsBLcl8Rs7qf3GIHubaXQGHPx/yde+MoVd+llw1T3XXjW4
rOaxxagjaeBvGY69I9SpdU9piIkG3twSvRzwCNqdCmhK8W6VEZB9At+YCbVXQCcM
2DxVVweS11sUhKUN8FjPiUhE3LY7/jwl2PEtOiY7wsPu75c+qorzzabVIAzbu1eO
4+atcgq43SwcmtpENIQ+spBRn1k4XKpDLKzIkhyhyv2Fw7fDuWKB86VgIZkNX38B
w3+8kHZ7PiRJpYObK/190Xl13dIo4uT8YCQ53PjplxcWYHKFAS3aSe28/ypFxzjI
ugyYJKbvkc/S0V1u0kPUVnDZcDci8r95h0K0FJ82And8cm8znFrqGfNXufIyby7b
YwKUErbjybyv/6PIHzD2uSQeuAw4SYKkpoVWy3ZNKykAN4F1E4e+7gME3Dx+ifnd
LqjgDsAA0NuMmY5nbFYkvuA7GeYhEOURMhq0DlDnV17tjaoBGj2AYrQRSo63BtEZ
sZWVxqS/NUXU1NOXlDlzMycwC7SmyWN6UdJPJxeOoovP5BcZjt+ivaIryI7OgeJX
EwDD9bLrtSxeFfDQvrwaeDptup/yZoDhcbMueRM1lWBxXl/uFYS8fcireiIFi7oj
zjI79rMAYiulJ1B4y3aIYJCMODHGlpAA59nAvgvTxU8Qp+9SUYI197z7zCggZ2ik
OzgDoclA7YA+UZeXi5P8k7t+YD6kTCedgsDAQnxLJGpdgBj3Q0nQaCD0Ij2wKQEz
Xm9V6jNbfmauwoFybHJMtuSB4sapJfTzgCw+9Qarr6bOWVsuZbJABeRZmmWNHX9V
nrmzuzBAL0FoXa81yPUIvIvwMw7U9eko4DjLTlsuetN3czWItgMnfvAgKC6wthWQ
6LE7go9F9OlscAQXhJNy+90qLjixpPTXYi5JjqFWCEhWl072Mp80drN5eY6YeKHL
moC9Y8H5PCZpwurdc1kDo+VWVCdO9DH4aVmnnAAAlpEJHxXNJGhIAxFv4+Zvz4eB
Bb9r81I5W7FlH12qGY1ppok1D5ewA55+JwTbxDbGuzXSTr5vG+RawpAKO5ta0uCw
G+Dr8vTmKb9htIXAb1JrqogELgmITXmCuK7fIoUxkurfX0lgsWqwBIu1w4CX9Mvz
iHUWOTnF02Ym0+FLYzJ8cD8ZMDsZly/ijIpO5K3W4cktR4Tkgd86Mf/Uoq+NcHiA
SKNWZJIoDNOHqUWylKVs1qWmWWFqacZQsJqSFlQnckTIbyEL4dDhmCrF23HjWytM
2TFIUyPhHfMfx4OGO0do7+jmOL/Mo3XtvadmJdxlt8cDlbzcqPmSvHvbtSBv6vuT
G2y37NXfTGODQbGodgLunoZu34CC+luNbiTuxDSrStTOgc7eigzJlBse2NzquYJf
fUoCyVrcwU/iKRnz8hl8Q2T6oQJrCpAlOANQErfR5n4Xe6jxqL0eUCfbGARCgNU4
KxeyJLTUfOZIRt+hIYk8uMjY2Vn5jhbQSKyUeeFUKDZmKS1+YrTbolncOX44n7XQ
HqFhhoegD5BCUtmiXD8200qmeH95D+V1BJNc379+vgBG7D8m3uDPZak2EiCMEUCC
fF880as1yEKVd8UIFyucgwmQFRjFMuOaGaSGolMfOGx098t3sOS82pRXbdoKjyL0
16zB+BFipi8D+ICZNWle50RBGxVNv89rxuUsA5TCY9WS9cpPEv7468KgPgr4GQhz
DTLB/cUdyYDUic5ZFPPXWzeaIANzKBNnxWFlQsCUX5sgaTt0gpzA2tpDoiqsBU+4
h/oaVnX6NtK2nTRPQzUvhKg5ywr000XbgVAi0C8d9AeB8ikL0L/aKjQ21ERnv93Z
h5lSDDVZNC3Qr9O8FJZaQnpZDDQNXdCi3Ikp67rqsqLsHinea0lDsUc7xVMyUqd9
ikQgv1cpPSBEw6B+Bv3BnZ2kKvqC54DTsf9DYa+JUnvxVtX8ZxgcW+OQr2X0n7id
4BRYK6EZWYt/rgybO8a8bCg+kwukkI/rOwcgcoyn8ksq/FJAy1eQU6aj/DwJ03Vk
XIRXMk+YbvE9rrgt0OkVc846UdmH2fU5qa2L+nTZkYRlaqXxnV1dylNUKRFx99I5
g8UHT6cCCbsGbHAm5Gl2K9FveFIwRMa/U6Xre12lBZpUO9YqwEKD8ccMhGqiDvyJ
fIsL2+FMvshvsbMeOM37+gLVstgh926oWgO5SfPWJ+x1BO1F0vKIXiAj6DJXfSQw
g9e+z6p0hugZhhgP4+co/a5CrDoRIbLpE8IiGSMxrvcnitjc+JGCj0+Stt2a2Cja
N/0XbDyOJDxQwr94pGfjW5BeshY792ixYxPYGc2N8pePHMG4EeyxDOubVUUP/QVx
YbW7TeqNWKwH8/ZKVkeKsZkseEp+1cOj3JvQTeigFbWfGncnFFuXIXxeDVc3JH5K
VBWovbAqO8hOp+/wm92iwj1jesukKbRmKr3D+jYnW4kmDK2gx2WPp1rot01YfumF
EQndnOX4MNT8lGZ5GorAhgTYQSwJISlG5uYX6LrfTHWUPH1rjfFaZfAE6kOuqa/7
ZiQmoQ7DhHXTieFtvmTqNMg2vjbE8xm7oN08k2XReRQpvDQVMTkfBcrKMFPjEkZB
bD8Lz44S6fbMZtew8+6ZQIhwyDKBle/uGk08dd/TM4Uw0JpY4aHDS6SEsfItD6rf
lS2n2EjkvGmO+DYsZsmTVyMdAUVq82vcYK6AnOIshILcbcS/7NjdRK/wcuP0lv/R
blA5EflXeckpVRMakdQC0GJG+n2QiP+5Jes6ETkqqCayb/dUA1eckC5av5kCne81
+biw/c6RLlpWaavshDsk96ASljUVjsO9bORWugKvXcUamWoHCLtkj5ZGpdW0c/2t
Ka+jdV+KVMkk79USYz5M91+r/giqzQvU+bOzWAaWt5GBtDJsJZFZc+8SkxtyxFA3
LYvYcBjWU44O6fPhLkKVetfk7cFltsb7aUyxvb1RmndTnRKY+Dnrir53/NhH4Lqp
WNuOb6rKWRAPb/AjKjJC3egI9pAxfeLbnN5GDXjm+63O7BelEI/MCoHOIZ3mqW+e
4YZwLqFs2XSZivllD4VjqaCjLDhHm58/UTuxYIi8TaqV8oI7QPTMjc98IU+9od6e
iGlwOEEig1SgDaXZoCCcXan9RpzAR/7tQiDZdeaAt4bA2fiB4Ksc02A/P9Ywd6ZV
Ml0WdIRQpMGu5yODz0Uj7OVgRRZ7tdTonB5k/WpsrxeYIcDsT737vVyfxAkvkBtz
oqpmPwMlZIX0Lf4LFqC3H9dcHFyd+MyjAZvQFh8Or28dnTjAvVSLoJgh6CpyNSVK
so0+FqpOb6rZTN6I0imktmlMyOlJ2ayv4VtIWPhazlrAcghh2jXzzgs/4PlpVg3I
Do3DUIB0x//vv6T0rQL64WETeyLsF3ZSpf82Pvs0NYACm4CWk2SxQjo5yKz/T0LX
CIt2ZvvcSJsh8dIprPEj08NdD+OiTTGhhpZb72LvMTLD/LNNi3P4k2wx8Ta/QjFW
IWYmREcM6qBw8ybmecykdGZd8SrX00A7Mev6oa7ydIo5MrXGrr4zjWOiszMgaTPk
q78aorHir+RXfbeCzMy6eeA/I34vIIxRQhDERYwcow9JLvCoAD0WBxKBy/P3fD+q
aCgeG29nMRjpsOAiO+QIrQwrAjB7ROkJL9+KaGpYg4M/iw6oa3ZgCbFkMFZiuMsB
qh3l619VEOFryk8cmJvsYbl+YEOYysYNTxuKwMaByIog57GyfuEWtIkLqZetvij4
xjSW9wVib0QS+2iTObIn8ERma8fnhYuGhYkdXh8ib1Qgj5b3tFjClEeuv7BaYKHe
Gj44Lav54aOKkNTUNXNW5YJ33B6UqqJVbj2NwiJ2AmFlEDIeT0EBGe1iJxxRn/su
r3dIyV/33X0qqhMcHm2MytsHjNHC6r82DAilYM8XveDaDCdwtoFrMXfkXp5E1MMH
aXaMhmGMCb54R5v/AtCJLEsj9uF5LH+7ur/w+QgCUuVm0a08NcRk7MtwaHOGtwWD
mP6bA+XnuoPNsDJAqfAWCv/HsZuGI1oH9wIbrIJK8xbTpw1mwP3lUQMsEXMAYmSq
UYDikjQSjnvdskVzIa5XK/bbvU5MFJMxQQ6XZ0/6bLHWjV9Gnu91dsjbqJZZtnOM
g5mO77BdKEf4pQm74BsmaQJsQgOvVxxI66bchffGqg8ZkbCBqzPNg154KzYI0W3g
yI98D9sPkRbNHURlIq7lfV5VCMr+9PUH0ibay60OkTleci2/1AdQ2vGe6iRF+ChI
P+o1E5CS6GZoZcpAXm9j6JZB2/tLg1EovRcwvjpzcnDMCa29i7e9HaM7l+fICq2l
7kH7wDP5QuJmy/JFWczSImrSmK8Ar62v+SOsQXa4NFcavbGj7Zwgkrn88NDgZeRK
gasX8VK/qtwS51sMG1UG18llWSOICTEzxfm37Wi/FXHqNCOIEgBvMzG3KJaob110
jqw0Q31BOpK6t7XNVhOGTUH7wdEJ81qyhjMyihn93V/xoP8mTL5Ind+FVu8TIPgq
stmbycxDOi/siO8z8JTCKxwH8dlBSaT5Z+Z+Yw+M8dPEMZOE3T1XaMo4gdIu/VaQ
JYOky885ygR4JoLJGFGrtl79yUBXM0U6qT8FbhBVtbSqxORBgaO+hwD9AsMwF7Sp
9TbKJtDavOxnpUC2zTyMRr7+dSU0AoCCRX8W4FZPDsw33yJZ/5o1UPILw0SewCxj
gxlS4B4K2mDCUwqalEzOF0t+Y9vzxrqqDHgZSKAsX5HN8Pypjol7t20RN5IScwkv
4hrGXcQrQZhOIe5FsrhU6ZRfrb8Oyd1CAQRMVKatUSLMKPepiV5CHncZfQsEqgc1
wg464k2NuIGc3pSkLuJWcV2C5IjMhBFZ8Ks4hSSQaptSvc9sJ2x3wJ5MRHpVAx5k
8J/BlGfm0d8pcKurfBPfo7ukxW2b2moxKGdnSxoyK64sJ9p6C3Q3+rOGn2U6amFR
EFa5e+SFnTYYfGlAS6JMYa93ptfLpA8E/S1IZFjRpawG9RFicZ9gcHH+Q4rSeA85
wyu8fla/yz5k5Ypbg57gD5p8CMJiDfjfOSeCVEb9tuwUKkcRoph6wib4jvIi5SET
KPqNhbRrX9R/w85qpTwzPC9rcWaKEMlPwRa+jC+uCalgYPrhgjY2becJPdF57OxT
K/rO9lXND+6s0RATH7ci30deoseLlpOjmGUlIzK8Xp8gAPj8NdKlKXeZeCD+Z+cX
K3ob5kN02uJdKQnUhJ5r9TcZvfW/uGHfKoFZkWNjmZ2uZBsF5927vD8eHZwsZL7V
h9dCiorF11m9dnA+8vDfK9LGNtO+m36U6K9aa6/a4w2ZxqH9fAy1Z3nlq/dhFIoq
uujpJBd3/YUKp/I6gacy170FBXw22biXxXN8MU0k/CyBsIiuvjNTU03KLwoz8HYj
bngg2yXHMiuZB6bRjIxoO2KQ3VqTAcODgE9eCUfptLIARKrpEfseSopQJe9ejy0g
aDDsgOZKKiB21j0nByCnbvp75y9x4tl7WVbfcbu4xEtGQWIpQnalHznsYWyTr0Kn
S6vae/I3UWM8KCJe5UDMHSqlrtwHjJSAFrIUrSyZBjNY1pifQdYK6gotItuTTIOW
aGSn37QuKDmCoUM6k3klAIaPscPl3TNDlw9EC3EFrudtTH9F1kaawlrMQkBZaxVV
lOPFzj6c+7+aRwVaduxwEx24GnMAZaewGCUrSVaoSngViMRXpALB3HpeAhQXeVYh
4R1X4Ilybjb70cd+kVB/wNJc95U9gxzBF6cOgyJRnB1eopoRwry9tNJPe/1tck42
pMrWs+pUYAGrgYDyzJD7MJbq51ND8ged1fIM1VaDi6J9cDAWwiHIQzLR6W8h2J9p
du8qB4xDKC3ynP/LKquhHxUOvGr5wVENnhienwZBUteU5ip2jJ6Srp51ZFzwcemF
p5mbWa3UPDtHFsOFbMO7VVmywyel8LnI4OOJ0ak+OVEEsF07uWTodOJkLvW+Ygo3
V9WkCpy1fw8CebiVAor4MP43aDCY9F2/I7tu8BT5BQHho2c16/mOF9pn7FRR2dL/
mXGG1GRbqfs4YFKqWrogLiyjwzDLKftyqbh74VJ9fqGcs2DMSDO+7AFFwbqbTrSS
JoVnCHS/fjqtCQz3K4tDeIl20TMFtuvNQc3BzuDX+LXmfYTlLtapWuvQcSHWdJPN
q7LMRxjj1ipfOS4tqv2yl3ypiKLT/juK9Ew7D+CJWlgFsjxmZOTSWwVpCivRk/8e
p/jQDxuh49Vg3YT66fOqxhysZNwhQFQUuAj3T1034m3IUW/v47XbjnzwM2oRvuLn
RbXjHWtAjdZUqZA1jc1N12ztl/cvexTQCLE4GVhZgjheMJ/dcqooqRpXdAPNQjsu
MtD3zIQNVxHaEmu7GhfDHkjh7IGvW+hbL3ThCe9nP+Jp62ByGQyvGPyJnFgGmquc
LdXguEeN83pjG5PAy/zg8v45xYQKX0wmoQVwQto51/h3U1QCOsOsWPtNg01eDEdi
XaPRh6tAaUBEXTluD04opmDc9k1VxUHImETxZs9M3RpPLnGu/gfE3zrEVBStXxkc
sxUj8sZCitPtvjabmsKlIOsX7F8uwWB9brlATcDqRqyLm9NHUncLiHaEM8uvVgOw
nVzdDKyPqE57hPkVUScpMUbFmOVzz0gfyGqWa4kCxuStDa7yoIEA3maERYPJr/KR
4QNlGEYVuMDmAku97x4q1kEJvKdVF4Vd/CcWTCb44awkEfte7/15OO6iYBSJCycD
4wsLHmTc9MmoH/RylmYXckorLN6o9a9r/QEobN7B/IZB00hdqzwGlygAhdvakUSw
FmZF/hehhLD+qxS0/z4ABwoDX06Vou62m8w0v31rV1d+0zvgJ4Bu6jzZABbSbFMr
3xkDMI3HIUiO6pBbakENMEH3kmhsDVNTm/8hQ8vEuzHwn8irpNFHwflyBj4gpDRc
u7EluCir6/lIodYzEdPc3EI37kQ8+DN1XzjvO8rLAErjn7ahr/cr5siiS9w9Np7H
rc+9nNP9qbBq9YMb3RHgmuOdDR7i5yq0H5Pp3KXYtWuyKaBt7GPhgbyfb/ceoPig
tJ13cm7CzZ675ZM+f1o4j7zCNsPqVOkLxeW0rnF/V5gDmz0koyge/7OKsXYMzM0m
rlS1PWW2conj8O/kgzl7E/+O8vJiJdwYGmg0a2cxNjMaqGtEGyAZ5NLEM9CPN9sT
uzr83viVqMK9QICmhVKPdgUhxhbLrtnrYp47pTaOClJjirpkAgXeqYd3xPdNxLrU
GegB3uWhehWrvNPNiw6t5EOXQeNR3hSkGDIhRnG+LXSkcT2JYij8uF4JpOQTCfyF
oeI9DI+/ujhIsTIrUwz//qtIaqvWPBwalg7IIvgidMgOUiE9YOrGasaSoQENKtU7
kB8KxOyT5nidJxbZYPEisD6zM/Ta+BvR4JFSPskKDea1ichUiabBzODcSDYuMMo2
VjFZhZ9KnSo3NX6TsWr3PXidaCiOHc3bImAUTeEpn6s6zX/UxHuu0DD6xjzM8WBg
dSbnSzKpsUMwMEIeqeKKUkoruapQJfQmEQmPI+Z4aZc2p1Ah1103rPPoNRC2G+RU
ZXSiULYVTIHCl9Q7++Odu2lRve5uzOWpablBEeoEdXnZFZLaBtt02pBlJj7hRBST
ciqgtNGl5Bf+q07MiR53CuIuvhKj+YHQALuE/LOWJoPLqKShAVfTVBsouaZ9XaO2
Jt3EHeUjXXpRm0nDSj2sLt20yl05zGIvwaQwpUFrc94OrbOIVcXiTu4WNqZsOq4C
efw3M0G1omceKhuPGIWuc/F31TSTrK8b5kNYtcf/XmDvy8eonvZOu6s/6Nn6ag6p
OkjD3S9QNHUzJag99I/O9TPyaxyEHM4we3KpskLOcuTEYPlCOc3pyWb0F2rmvYR1
6C559tJ7Wjd9GfL7R4LdDQAXuBAWiJ1uwZbRgk9h4IoI0O/WK/Je959mpSrn7qKj
OeFWkN284Z5vfdJb17v0eS81nHoINXtgyIaSj2Oq/MnICDkAv6Ec5UsM3pLLaQcd
WnL9GOK48EHdHcHIUtSntNGeCsmrci9iMCF6bfuRR96+lzp4i6r3h532RLNbWb66
tma1SNb0FMcgu2omR0uF3aRigWFErEz7LNSOg7bTRXmPgX9sWWVAUkHWRj/z/Jdi
ivhValMnbkz7Mt93a+DE52YGVUz60Dhlw8mMh3Rfv82zPcHrTib59Xc3IcrY2m64
zGVyJKiBquHHZulxWLpGb5aCaBWjN4ENjIu3JuLNEDEGGgVMDrJ4R8Fy5p13lA3e
YDwelzprdnZFx47c2c1hbkgh46fgqSCLE/Ol5ymeibB0kvM9YS2NzAGXHic0Qgqs
M3hs38BZrddvhHb83HiSCPIEdEhvtdlrpqWnijlt9YXX5wASuxDLVfXONhmmONR4
niirlesYw7VTNNx8N6v6YAG7tVPAjfEvyZD8bVILshoF2u2dqZxUXq3d9r3uo/lq
JLgoMBhPGpujYNgFS8y1G4KXvHjQgHTF9R5ahBmXnzY7Vkt3LnWHSTHIus/uIVuU
Dm17mdx6AFuNXDLrZOqmF6bQfKJp88ksZefWXtuAStjYW3MXds1zZu5fbx8ih+wU
dwJgo28yJ04oDoW21eup7oL+CI4XsbKgABvZOKFLvBID9ulev/EEUKveEnS7ezL9
F0Vv/SJn6GmEtPvFIcQ0QKsqNtAh6ax3dP7qJFT9Y1h1yY+BJkfr7S7G4hYiLPb9
VLlEcnt4HspA8aL8gcMV7pZcVyv5vLzX5CCiLumWQ9pvi5VT6Cfy4XP4RS9VCctB
4XIgld/DmCf6b9RIIJqEdzdGHutb0xlUTantxCEkIDLmYRkWNIbhSLcnydPUy1Bg
myCKptHeYWpde4oFOIFgLBy865TeyE+15O1Gx6spelSugs1EX/1lZ77XPHchhyPo
/G425588TsDwtK8zIWeQWPf26KleRV/qGGNINZVQKYJ8or77lTzh3Tw0hurAM5LL
ITROF4Ia0dewgMF+U9zqZ/qlibqmH1F9ZapV5t5iNdglVWeBW3LtaaGuGy2aV4CF
Ug4RYSDXzlfpi5esl0T2aJ1BglrjoXGoGtXdz9ckSpZgGr6pxvqiXPbCCRghpfjG
blte7Pcaa8P6KPrLsq51hIwc3GTH5uo81MJzLnl8Ld8CrT0tk+lZXYvjkxhtd/8X
7/C1hu766UIlBqONL7Pzg7NszCHLYlSNhwtyN1lUIlrjKkrt9UoA+Iw62acI39Na
+sjpWNZVZzilt92MJOloY13v+aAOECJZvDJXjwnhfHAPw4bMfy07fO0zol7VAMCr
PLHf/lwIE13xvhFMoY3qGTqjggpABT4KCgnPndgxHOMRFxxsZwetZHURCe6isXx/
LZkaJN4ov9YqZ8N7rYwnmQLehEnF5guxEnNUOIrgPyrJWy8KEFtqC6gUax6Ybu7U
tSqR2fsY3wY/ZvBtGNFFgBIT+13Xgqe0fPmFbbptYv0yCLZklzwnueaNWKyxWt4a
CVi2hs+d8t/5Pj5cgPcMym3ezmxBFEEZ2YXckQR6IQnS8uJ7t1ftVSw7u696dbot
LRNNKUWuHruay466CLWTEsnLeK98binuBTmZrELkqkwMeO0TLXnTNuQwrsrbKMi1
qA1aoTnperr/+YdpLNoxt9DuaMxaXPFBg9MTyFToLG5F/1Vi5H/qDG0NswIhQDeB
/Si83zJQb+0bxDW8GQv36zIKgAMXM7wFG/ZquWK+jUh4axBNyTP4hgBx4HFUrHTC
ojODs6lFIY3cHhEGYqBPj6WU7oNhDJRIdM55m00m2Egy5GPehPzazzJU0hSKS7Hk
RZa78qbHhQt826cKNONvnZBntmPJzIAmcYuIZ/5cDICR8zNm5qjzQoU+7J4SBwFS
1agCaOCo+TJLKIGh9h+vy7/GZlQky6hdxp/C7e821kWiwafYWJd9flmAiAbwydnF
lH8uZzaTzEDpp2cFBuX+xvBrQSPmoPDwEP+0juueKM7dFJYgvCobiVC+AvtXsk5M
rKkoGztgnDgaUQlkrS0sytVt3hHB7ApObSlUzREO5+O+NDrQxaq5RqDqsopog0hl
dMXi1AmQ4Xtk9wCgYMJ146C2PHiqi1deUUI42rDILfCpqS/+MLdRQMQTnmSJbDvn
yRUfqSUmvBU37/oYY+VGB5/QQao4a4a6Mv6LgxdIWBbSuw4E39LogkRUUxP1NTtz
wuc/DU2o1zrVlqrZ4pHB4v8P5B0W6tLd2kzXzjXjIRbUbT/GLXrz7r4dnti/ZeX+
iAsnWWF5Sb+eVm3m9vuLh9fF6h5wRNACS1Z30DUNngA6OFCE0r6NDQggLp6jp3SP
GtaDK+ukpSJFYWi8Os37B6yVcfyyfEDflcBbzEu1Ks13MsT6eKqnkk0FpvBwmR6w
8vHtwHnyFaFOEDc3SEifsCLZ3dU1aNVwLtm9wmbio1dxFjbIkhnmvH5FUzbcd9DF
hDLPYtIn07lnN6IPNISHTHKDzKZA3FGfHRXeS58iAKZa8e8S/6WybjvE+IIkjBKU
6m6ZcOpXlPpU4hFjEPakLOVBxzQHE1nbHZmtD1LBMSRkK9hXGCARIRzDTVnDF5ns
OBAp6E2HuSE8MVWZdusOzlC49QazYWKt98xsTWcO2rr6rH8wnl0mNrH78idJz6Rh
cpEnYK/Q2ip71LaWVqakRUNiIBs7xZUnUv06GplTKc2KzHopKIdItqYWD63v9948
sM64S8/9UmFvlXM8CQXmpJA+TDN54S+qtPxi98nccToOJOrSKC6l6jeycOd29Udl
og6lg+9x9rscAEk+alq2WjHAh6nD6KBYyMKlyTpq6asrFEgGOmPFSH2NBHuIe9Qq
/beNswJwhEFiEKB4D4Vfd9Dl3VM4ATo8bczgVI8U7L46h1Zeqo/BwRN/DYbVPIfN
4doFwu/IDB03FM4c2J321kbmXsh3opjrkyUaxk49DfigZssi7U5CyzxLZoXZuKnh
eIqrYO3axVzDFgdqDOKf8bSkLoq17TMmBi2FS8K3kNmBL75bzdkJ9rxREqUVgIQo
z5ZIZhp2Y6JFMcW4eB1TXVg3/wBSU0zdaaoeXmkv9ByVEkxZHxuzTtA1NA1tO2YV
FIVhZe7oqHXTJdKTU48QRi85hSlRczTsJCM7j2h4okdKvPciUVJAoRB2lZ74DHIl
eq5CykKG4kzp4TIxmTRsc54jBUdV4q5SNg4edTGNVVLcTYvMm0ieLsRm2HKzLCQb
5fDKU0fTdILGfRSmXVoIeMeTliQPgLmwsOROJfofTRspEnYFRtZ5nZcjvPJ2jaSH
ahO2FqfZ5ZQI9pQXaHgWFxFJ319qG3hY/kW9GJ5cT76d9Qo+ugsjpC6F3BHy51Wd
PVJCZ6a3F4eQnJWAOue6RpfXh5+uxZ/53BKKxD9UvwD7Q67K3Dy/R+U/LUART4rs
kWhlvb3rnTVurmwp2TMqO/O1M2g379ksdduUZ/SDQATSR+FGfsKz5RUdSszxGJH8
6q7eyoytXGToVWIInfJz3TQEV4iTBiPrUu9P4w7gJc4bSoOLvlZ4MeeoGdnUld/t
3X3iSOvsHtic1c/snLQI9O46yQwLVLsIrK2mh3748YrLXauZ8o9xK1fvsfpiCQHH
7nWqOrWrhJVH64SHonPGO7vKfjuC8tO1mrngaQTsHFPADM3WkLkGONrALYbVh/bk
Wa7l9ST39+novQUFHeLtUnE3hpuH35HXFkAeRZauhpmceHziZiUgaADMb2SD+6Qq
ibiKxd1uDrfyX+JTw2Cre3PIgfR6hJ56ihtc2PFgoC0z/g8xUcxhtivJPUv/ESkc
Ecvbjgggfmb8pvUiYbhPXUesHYc0aCXjE49ntK6ZxgNrqyvoE444r9Ks3JUFlDMQ
JAayVOh8ZnQ8mihAnaKyoJTNyFPHT7lQwDeiAkPkxvk+y3RQzAWQ/uRpEVea+IX8
zTkhKgwtjRpYXVn+GeTTUAAuABa7AsVYRir+2YwbIDSCuBHsJorQI5yjy7khBYN3
nVR/dscvQNs60klO0HTaeZD3S7kbyo6pQii85pLUxcANeVzubqQf6RIsrpvvNfOr
b/hpBjEeQl8JOfoJKcASZcRIkBCvbCe9MW6FB6f5uHw7Uxrsi7jztnqa9gULs3Ny
hbFH46NGLs0vooBouXzQTjw0oko8oqgiIxWhAQdGgZEP927eQHhRVSiCbvRQRrzw
7HFZuWF3SH/Yad6d3M0t2nCKOIGiUKoxr3lL506GTptlL5sH+HbA2MrjmwoQayuy
YcC/IRJX/atWbSzgwfMC3Inb3ClaMziXSlxo7U1OB5Il04fvqkJ0Nf9RD51w+9BW
b3VDa0i5Ngfkl/xUcE1OngLvntooOyEljPXiE6gHCy/7ENmjgg2XN0rvO3nbjrdf
PW4Ko9zmoWSEdUEGOVU3Qx9zSgAe7ihqJgMqA0lilXMnwpcrqMF8047ZU6Ru//fT
3yGYJvB4X4UMivHKGvY7CyrN8RKsBrbn4+xWI8g+AXwo54lITG5iaUrQDA60kOqx
RLkIqI5BzSJiB/2Tfg2EAIIbDg3f6avdd5PIHZkpx0vymavV4aGGT4lWA7Teq/G/
20nASE8rDD8bv8ZNtH4D+1UcGdimS0lrSUFcgKaH8YCBsFfKEG7edKT/jbG72hdB
hRjCKaUEf/nkS23G5EBHXWXpuWt2Ac+Kk42ujh/6F/i5iCR7WwF+gLHhB1GrLqq9
7wvkLKrYeRvR/V+gYLt0y35lKW+mRJlW39M+P+b5D0773V/wzkFGyuhruo4CPB89
pKU7Fd85TzVNiXMmVJ3uOQj5iQp/h4o8S9gMb49vdtZ8bO/FYDXckld4tCJjUgE4
lJI5DxLKKpNihpgLYN5TTuQLLH50is8rPtIklcTJgcexkYC4n1m8cdjb2ajHvrzp
RXpG5k34bczipldcq5X/ztXt0pzfe01KUhlTY2E3E6sHtevQZFl03e6+2EDjAeAc
djYij4HRhFK7z72TkPocbm5sMUwV29OpiICc60IIruHqFw6ETIvLqfqwClKh95K6
HujkJj2ayzn0G3AnabLSflyL8WK2S5p+xCTcBN0FgPhoW9QRmOlkS73Z5lXzlWbS
RA1VRVAKCEZt6baZ37A0eYEh0E3GZDO4wp10xfjYArnJAN+r2MqLAWNb8Kt5Z5zk
irqogUmfCnnr3reHbIq/HwSdT+YuBeGDcHecvxP70l0gfpvTWsilThOFyD8LnOuI
f8OWXAWoZhS1PAMPm9Do9XRuifJkn2BaZc8z/Qu3OHC97USU4nAQRQ0bm/p/cRg3
9gxy4HMoyMOZJjYSGMFkUSEKV529YWGxdjFMZ4vFc3rCAz9j+Wr0GhqCyasI8NTV
R3QBBACichwaZirWJoz4LOXMK1iRZIlLkba6GruSDbWuL8yxLmze++kNG170PBLI
4OJaKN0qz9LUYeyNQZGEiSbjIkfmSEtZAdqxNCPhZc9AoSLp9CRqhtcKHuK/Ur6w
51FhNmc9fHykifne9Tbs6xAr+b/PLrgkBB/X6t/Aujf5iobDzMVzWEcd/uQEh2hP
OhxIb7kH+eQ+fCzU/wwyiUziArkuneaT3UBfviyMSUCjAvJOK4axTyfsOft740zF
c9NSs32HIbVMGqL0/FECFVvQKt3PDFJ2nBg9Q57PbIDyNTD7g4ITwFugtJ2Oa+gE
PfYHyPQWFnP8JaqHnTCHLcw5QpTT79CXGaU+KoZcTB4iOpRYEPYjO95Dsxr4WIuF
MFn0mhXfjfi2Z/z+D0ULms3h03Pc2X9pNz0zrzvufgtUHsdg+eEg93eiJ0pRds9G
Gm3xSKmQi1Gkew9Dbc9dMyU+aph+Fa/FdKBfXeVVTHWcX1oHuHyJtp/N/7ZMs3ZD
KBXa/Fu79V9oNq7Zt6RXSmGXDsjXUgZ60RfKnP/VLbuzwnJs+KifERXzxLOtmKnX
6FpMZjjr4P+iWqXu2LAy25lnlU4crA6KPLrXlkvVdPtJo4xQUk5y2+19iAoBLkDU
ol7oXQmMbveKSICOzI6zbez+7L+wY1mm7qfPP/lQ8BBdyJzDZb7NkP1p6ePSlccK
FS8hsuEyrkgQSZwrtNGD4Xg7Rr7ODbiBn8pqeTToL5mhVkBq49UvzxUaQvuuSGlb
QsvaVzZ90xB/+K0s6q3OokM/krdH2SANOUvebq5o9acbl4aWSUaDtvCD9m0VjEW1
HT6DT/j0wFSC4Hg+e2L51J+oHtnDLCUpSfbnvTbBg0FZ0Tym2wLfGm8E+FAK/KnE
vAjcN90GHa3n0ssX5vpySTN3TF5RDx1SgcFwWLBeCcFOh+bjJiksc7RZCqfEoGvK
XUCeyEb5s8KwLQC7tbbUJA5w3FdVTu8nqbfgF4k90IKY2YxA/7rTmhDUjjcj2yl+
fqs/j2KJYyW5EO5ph3trjirnGAQl9b3822d+JBbcKuPp1YgE2qWilrPLGbrjDOge
xJ3g/xxOZ34SzvfhnyKYtms04WnGNAZULsM7ZFCHNncp+C7hIXdiHE/+6dYyLu1Y
h5UZPb2HCf/vfBgFiO5u5hhDAZiVl3FhOMxkvFdi3gtC4xTUGyrmtwppK9cuPgtc
Y2OAVLXFAUwYoDDlPUS1yNFLISzHHm8b/bAhfu1ogAhYkRAJyEnsmfUGOfDVLHzv
CQJWQAZIu58W1yj0ozPmPKzKD0hLHFnof+4SelJrW7ulhkGTDNqMga6xaXL568La
slqSWsNIXGRrqFKDVILMy5bKrMLq4iMke6jh/p+i0195VrskIaPF1T9kchtaiQfC
8b7jV9UECMfgjGNH15xtSYWGaDrDrxGqtm9imb/bEczYhZ8K2UeOVA6igKN1MDR4
TmAk/8mytcX8GBw2co/LzyLDb79yD21s/ttmNBAuTZF4YfHfwLOVovtEotG8TT7f
j+e1yWt9GPoAbrDEY+J+gWwWBtqU70UDcznaboLo5frHa+jD/Zw4+J6Xz/chcdig
5ceAb7jfmHFAQPoVtbN7ddCWhO9F3rGGmwa2J503HSXj3bcZbawvdMzpjM4GJhV0
3XO6eOMLAia4oI2lW1g/hkL4JGBvEzL4JlMrCWB+46kIOA/es9uNgmKmB5kBDsuw
MpA6NrDx9Kz+Eq27ig5g9tiY1TjQSP3trCJME/VDMxTHoU0T+z9To0E5mrbxFhb4
EPpODYDnlAe03yNDPi02kh2oGw/iW0MxfvjmeCCS+jp0XzJb7RsIxSiUmPxzb/o6
wC27Ye0hYeo7DQjTsGoO9++0V4ewc66Naped8wZc8lr39nnQcMFmmFDWBPjNBRf3
qq87Jso52TZXw1kzW2niHWlzGto49u6eokR7vLR5lgHfojn8ueM5YRZjMaZ4S01J
hKyi5PrEprxGC5pgLn60Phkthd0V6qUYmJExgnlkhmU/clpqgOD4mwbUbSoNU87P
uYQVY259v/a6xlVUCFhgwd7EzaX6x25YytkKg2N8gYRlrP3mHnan/bAHy8HoZxdZ
U++G7DjW4sz3B5bZnLe2A0SIBox3U/Oo3rIC55QU4RIkrek0bkzvQ9BNnSJm8oxn
hQCL2VUrj2Cn02Sm/2hhMMvLZ2GAA4njuYyurJkZZaJWaFX3Z0IkjqPSbTKMZ4ar
MiS9vf6sN//JtWplri3xNrXhUbfPYe/A29s1W6OSKceqm2A5qQyAOKwFXtmaY2Qk
mfm5lmpEtSZ7p71fg3dIm4vO+wssD55I6HRCXVxiH2fTcYgnYIjFHoad39tjSuvO
yHRTLYBUsPp4GxuCCsYlkkLxNDxBsg4nAB8ZTdzDG5Tt6qH2fI4pwqxlpAQ4ZaZO
PE0baEYnpcC3ZnwW0i+Nab+9hVaAIkBnyO01VzkRGELIYhwVaJS5WqOxwzbNs695
OUQw0lw3kf+JezeOB/OXrBLrnUYUUo/NBLtNJAF/4MG9Z64ctkgY9QI/COkWcOzC
EPFwmBkd8MYAMeZ/6dE08hyt+iWrjG2pYh9I82GMunRGzvsNZY0Ux7zuaMYk6dqA
+oX5g162dECsjVgsSEiDaEFYGjdX48MZGRKu1O51J+fDPx60a00CX0R4B9zfTc0d
IADVjgpwh6SkwWJ9VNEDpUmx+lO668+tLTxx7Qow9CEV/QAygpRnUM0F9htgLsev
akSjquhPkdt0MHAmq3ABsk20efxSrUYCM6VsGusEz50ovU5UeGO98X5IZKpMvkQm
fjV0ClmeNyzW6aS6u++hpOMhsIR68Z1BXwlLM8Pck5zXPuAICDzgkIxads1Cyqsc
Yexj5MuuaYt56CcHIyTBLiB+W4ZiHtsHluC+yZFOjGKwNzcYHfmTfOhFEAbezGBB
GHeSFuxxIvlwJz01NrnONsXZsGXGEJDBzxoaY0NZQ2TPADHnMjNngAzSIR3N+NjH
glA5HDdm9JB02/hU2QgDi8tJzm0uXpwpxFobP2NJxhfOEs72IMTNoUJ6QAaKtc4i
idBeyUamPyski9KcvYn+2lOHwqm2c1YqXRrdyzLmeGQMg0+t0w8XdKHDNFmPyEAh
ryOUqIThIvTOd3nm452sd3uvrVZz/YUQv1HR+Rml+1jfcf+DYgRotlq2Rv2b/JUC
ehujxlABjQr4FYIP6kbsw6hgxDagbjrvdFUHe1CUt8JOXaRQB2i9FHAELdlSv8d7
F36UO8E6iAdzztC2ep3P3kKU7YejclzpuLyBvCnP872J2NwfP8FRc+bBgJv6aH5Z
CiKuzFWi0G6bbVJeeJMxpuQt8j7Mc1muXKRsJADf+ThB8RsRd4ait0stZk1Cn+np
fGrAXwTeMqUClvmGq5bos+Z+4dFg8mwhAoTQSAhZgXbKyorCfrYd5peY06fCrmQc
vocj1eYoEOS3gT455VFVLDomKGHyl/ZoQdZc1KVONCatrynIFkt6QccbdAEZ0rAk
w3m2vQgYdexe8lwD8Y+qmujjbXy26GFYzYa1Jit6BFnQ9OiqFFePOrqYAA6cqooR
NSLwf3efgy0xpqRf/JHpMlQC9Xen9FFag4za6RN68X6Z33izeXOV5wQNOmNlsOBh
34g1Miu1f/YHRxLtITZtlAGGuHnjasOJqrXoiJP7mGoMsY2QOkG9PcW8/Y+ofKm5
dhzEBX6YHVj5Q6HsTvS5upJMtUkh1WoQnzvMZTKOyx7VHDt0VRIoFp1mPj+Ec5q2
cSeg+sxwbWh2n+EOhm+ASBfuWJ9xBzmy6MIOclgPTVoaWAVYSGWS8HZvP4PAQJ4X
Em90Ag3H+an0xgGbuNbLr/cMVawMdjBOGmRiYIrqgv7jEn0Bkcrh6aiz+G0ESR3q
v5tc1xVEUtoAcviqWWVdA44EaS6INrHPfw4ctjlHVPoh1RLxOXhRfc9iyDxELoAd
uSkLre+e60/CPLLufWMBasxaVmMCcmWdRmpkgDqQnxV2VJtOVy8AKSgwJFjqd32z
u+DGBrLBk37xfFld5OfgCUuIdS9ObT0QmjAJxFmfzsse4UZAPsyoiJH17JOac7Ln
4WxxuF5e6pCTZAC7df14MFqMfFb24cCGc2+jEl9jdCj20vwfL/FclcmwEzB/BT3L
JFQG66ESCE09v55sRU6TaB6MfGOUsXMtfJU7lx+kMgf0ZjtdGKE6jHuBiSH1fxoJ
qQT/J9YvG2+pulV/ehTvbkh8FyfDrG7rzfxA6PG2u1HLixYlreArcNd2Dq2j9Etz
e/KnNBQPZSa3YDPzAAO7Yjjl0M5LcUilfeg13bHZm7Dx+UKCCqJc6G/8+33xH6Iv
4kCTa3LOcszCjy4H3tidOy3kgFDShbqgGhmSuLuq7QXXoarPj2BKmG6dKetBlfQD
5tZC51vjk1BPVB5i0dLR1sojeb9halVMrFprfZ1pfSEPe3dwYk8dG5O71U2gozNo
r+UPdoaYn7oQZeavNCJtaGbCocoyOGhRiV0OFqUqK4ykvDE0Srah++o8efggio02
TjkbK19yqPh39tKjYUqouFjGEPtW6BvIHIARODcbftt+UEa+Z7DYT7oiAIjMJBJC
GBDWvy1OyLVToifFzkmdaPN9bSS2rFmqZKHx/ybS+DG524/tijJLkNR5wt5cSAIX
EYkLUQfDSUwibdXKVw8BbtOX4lKj4fIs3vRanZWUehTfd9i3A/2uBA6CMEea4siX
lojYA9ienwt0U4J1K0Di19oZnCzxQhq3FtrZ0WXqFIZ/HP+UZ1phZ17QbY7Cn16V
eS1lmNIRb43vC5nUM54XlJV7CAkC7lVFaiZkzDk5FQUH5N32im+AOynz8r0a/2MN
ZHPnIcWm8FANRS1PZ66vg7SaRTbvnq/pxVid6v9p0gK3YV1kvOpBpJHEYCKXtRHd
Tu8iFGsFrEKXDPFqNCpWy3ag/Z0LVtxWwYCDNLKV7zflE1tSv+zfcwksYvP+x4V7
y56ViwL3Ckj9NYTKuROYpBzWDtZZ3egDA6EYqyqj5NyVVlf24RUuILp2zuCwATxy
lvrCl7vBZmblYNp6BXPuWHDIRm7snX5QRercxB6mk42Bp2heLnPZeaZJjAzIhj5j
gAUmwQl4CNSWkCzLyKDNvMBxpyCRjlEOHbs/q/MXNmCdoJA71nw3/tfZR/SdeOCT
bxPeocTZVbZJu1TxHG7E+4gSISV7Iy9j+/OvGvX4qiVt6oF0FKYlXk2s7yaMmrx5
CaVSjiCk7AxKQgk6vJv0loOiziY3rwTOONw5s4mC+j/hHKZqgwz5OTc9JWsDj6QV
f32fks0BLfXth6xURkfwKWupwlmQUQghKnL2hHEK765G7b8dyX/rbSmv46L9OGWy
Yvq93A5xII1x0dVeCmu0ZY+EpiqptG8vr2SkcVwy8N0ZTjKX9cHDR4pVntv8Q8zH
IJJ7iC37uJDg67Im9DCroRGaCGoNDvnkyRXWp7Iwuya+5FeAuAmjx3T80aMDB26I
HRdKkZJee3c2jg97tGN3+F4l4aYIadUBT/NaunL35YA4w2GecHzN8QYKVosfNWPv
hjh8AEl7ZV7BfK60xC32s/DLGpKMpfGRd5FctYghTnjYT2x99cBcShAw9YFybq4O
7eeU4SHdrXDVTXF1lBKVIJubsOpgYuiwxKRWDDKdPPGVft0ldlNcbTBBvjMwKhWC
Q5uKZpekrCXF4E9UT8lzoa+ZRZRwSTeG8D1/DYmzoiH75MgfCsVQquGhD4nZ6s0M
4VoDogdpd/oQUD7AEq5p4VVPq6R9p/iAjcY2aJsB3gpgTZPZBaSmHba23XPw9y3r
Yw+m774iOYeF1+9ihYVlAnlA02psbqKeDZgr4T6HdCdnxASreAqOlSnCaneVDZ2n
A3bNa/Y/uq4AdusJ5mtCxFylvD62/6p/cut9PWnfRZhblTzx6gGYGY7EXCExOWti
U1prO4Ox113p/oxtY44xtci31mLRR1snx0Iqv5LX+yqfrPpR2m2BJdk71ssTs5jK
23Re0PlmhmYxxAPMO9j8aqBt599xR8mAofi7NcITgYYzktwvky6myPfSeXozjYld
tzeIxV1fHkEI/fKtkI/25naRSdcFhIEZy+JShgFCmYbAAbIWfJMkhYNpvect8FUJ
Yls61j0T7J5d2c9P9w75dIuLqHr2/n9kJ3iNPeyulSYZuChy2xWUMbpLFtMs9Nk3
QNTmFyHGZKVmLGHJiSAAzK8GTzO4BMWUoxpSbfx9hlxmHszKWpBemX7od7+vOIMn
nL4OOyfWYfbOLw53YaVzbEHafcaxyeIq2YRP3SvSrIjE24enbC8T01rLZiopBU0Q
SGc0sfLdPqae5QCzuek34XP1N6PA9cWsPVOlsXLaLLCo8j6P28vGqOWVMOFGvclb
WEDbjAk+3JjSKrI5WDFgOVpJAmkPhLn9NxNw79T4708gvBRHf0wVOA7JtxI9MN8A
s6mni3ElaTtdnwUrh2bKiJyy01k6ojtt4Cs/J37qrxB3jEcqhan31h+8rZvZpdvW
OCDv2G2+8oHxGeHxTEFSg/S1tye/1YlJEOqjknDFw30NDTVWM0eax3qqbhJ43cK4
rAQeW9DsrZ2XVl8YAAv3Tu3XU3ZGda/4ndkFgwnqKdfwSKFI84PQnwM7G+9VXo8g
364CHlZ36AFdpKv1o+P45xeHB7zb/wXQVDMStYGkDGMi3ki9sGdOCpVTWQn6AIwu
/6DSmvvNfMaTvGDABCMN9uVqacOEbUlaBAf46XZ1su/j1pFx8m1yclX4/byBGUPg
9Y7NJx/D6ekhqgfPnfyw+bebuU05acuYTmHmGtPEqypqoCnkWG+O4113ADgYOL4G
r0dhn6LegGijHvjOC/yYMVCyVIY01JJZGqvKaeFUESr+tdqa3PmjLhGZxApE+4B+
ygjptqT/6xiO86EpHdq4wqXE5Tb8ngG0YQus11vqxnczjcZJALX9MItYeMsQoHcH
Uzts/atSpCGMWka08aEIQW+AwkzXtwSdac44RLbqhqK/P/Y4KtCdsI7ubSLA2EgZ
q/o0npkSAFuCz/GmRxDBqKwj1apNBwrWJzv0awxOTpFOJgMXE7PVYuXKOOh0S5zD
/EDlHWn5hTq3KN1WQgxPI8WGDe2DJji+hr8nYbib9rDD3EjrX/42r4H/ahtnRbAP
2b1H+qZFqtV3DtV/orshyhbjOTQou9T7HVs1Ezyz78OTg7+t965XUY6HMwwq4pDr
z6QTSxkXXSoDep+vRGNeZHPLMv9tJP7Z+oT7AfBcQRGGVGMp1Mbx+9zKZS3K3Xqu
94r1rboFtyj9+cZ0XTh0MlgmDyjgJJvSvRQwRrqemJ1hyqYks8IFMVIBMjqUSFSD
6P6TAM/PZOpi2hEkrwStuBGJoTg/obQwzoBXpfOwQgUVh8qccyN7JR2PcmUvqpA1
3Am1Jw8+ZISOcSUSo7g0LXrrALvBnSlyMMdEIeUInp54vjGawfFUtjFjaBN6eHm3
7KFH6NmIBPbxyw9y/FNWpPkssQK0R0Gc+I7nHL5SuRSLokao+8hSGqOX/L3FelBi
/Pc44Y4LXEzCkd46o2iiqQON3OEIpoMknwakj6Mus241D/kcCKkmjpuE8GR2+7rE
k2JkK3wEz2uoUEgCfaO+Elhws4aCh9tM4ts1jOWF4xHWpuYZSANcwRH1dEuXaqXc
3g/KNbajXCL4djkUGQK37kpPWK8R8EU1orI/MJIn0n1aY+t9yqJeasP8nYD1g2P3
Rz+Sy4zesl+30XK+YiEugL/ra6lWhTPheuMyji7LXb7uVvZhDZ7X+4/HzOY7I5KG
0+r5AmVG9KJIZRJsLANebdWekQvHqXAOD+VLtnBUMAbust1CIgegHqYogYNTltmN
a28zCDhbROvgSveZUfy1ESaaRDw/LEwjfwAw4jk7rzQDm5HW3sD9ruZ+gcDUZt3s
TwcIhA+BTIHuNtGYeAycP9W6zukvLBuiC+gO/Er9Pxsd6bTql+agHTLoSzgoW2WO
YdG4qxSz/KYDmG3cei8I7lS8s5c2Zkv35V5BoXb6jPO+6L7doOKe8aPft4hRav5r
rA3UhPb2uvKbnYrM7rGoOR6hVIUMbGNNucjH/EwkubaodFYKMNIQYRG7HQLrofTI
8j4wMVHUT0r6Ria8bG8RMrgUa/WI5pGdWlpfox2D7EXd2v5/fdYn+JyJzaoTnzJV
cGX2vIYp48QsaU/7hjRtAAdsJmySm/9ny4okmVHH8iEHjhLx15joF1rxaScFTqkh
t1l6tHomulDIDLpdYSvwT//1Ayq3oIeHG8YAN8ZMVb5i3/qaell8JfiDU5YRHBwn
v1x339HIHK2wzqWx/AaldWV4gyYzkaIJwGaj//n2gLbHn7L47MT9Zh6w/avuQsPu
LurfbMklD/AnZzwoMO68KP9vmZbBAfdVwjBeav2t4N6PVvIvvp4S4O3XGoBhDHQu
YemCVIIbJCP4DoqIfS+WXYHh9tXZ2G56OJ0oklPOCI0YU5DX/dOeneKSjbI6S/RY
/5vBkYcIIGRA5ao7pCgiJ273d+bBRuXKU/CQ64GkBLObo8eG2hLqBe+PYgVDN7q1
H14EwMuEJGtzzhgSfgW7rBtuBwwp2l157UFpRkZavR3+RI3DZzmIdNpoJLK6WtYk
Ew7wF95CXXHvImd5e4pH5siUnWCdYltY9/7i3DffZ/u4LElGe2Q5BnXEFJOEv5Rd
XBbUCo/yJNdIbBus9RLhjHBTph5ZKOqXPWWmp/Ws7Mf2zMP6ggRoxMU3iy1gxay3
IhhFJN75SQYkgXVHyB8ukPYHXYaQOngTqMuyw6oGXsY9b94Q9O6BteydO94u/4a7
eLherIDZ9AfdX0AsCAaGR8rmroFISRrnK35k5QcLSyfpyIomUjoKnXGRDNzAiwr4
TkVUyAgZCbJ30JUlE2xpAJfm3LZXbm3JoiGXdOV3ZZRB5uo2TkWZ3eBrLtS7Vkj8
Uaw1MgQYD5/VA9HXlQRt9ng16RNCLI/EBJDHcv+bD1FpixaimYQcdy7d+BbENfYr
94nPLNOxLxUWGb+SET+nV2pijpd74TZLkeNFSRhIi2hjiswiVG61qlFQtFmfCoeW
OZUR1hC09IUWebO5zz7p7POSSoIBR9rRCdgdxDzQKSaujx1woYBbhmjZ0i3E2V/I
KvQnAj6HOpq05oQyqHLP8lVgmBKV70SIZQIkeqRLmLn7WAJAaaw3W4tqVwVnrZmw
fgTjpdv1Z4X5KGKu4hUhuCKvPzZa8qbE8skjeZogt+YnsfBPOZm6ojSdWY+tTav8
2dHi/0CDPCXM4HALQkEmYMiA1S5ZkLmC2CYhSntJjFPoQmPVe0EhYqSIhZkch1wR
X2w+5llC0mbrYYgzJ4C2xLJkQpUQ+fyA/Ovt8sd5vyTZi/q6zl8RISi1SPcvuwCV
6KX7uq9e1xhD3RxnCx1hMgziUdvNFZrZN1Zz7ytwgD2JD1TMWdCB5N9MbdcPBx/d
jkC7iBGwwLqCVyvrkhIZv+hHKTp/suGU1qLTQBfCnjRr3+IGJXwXsPPnICt3LaYU
7ww3P/lxRhk+/FCIKvgoTuTvzpDqd/AYwjc+OLD160RIjsomwqF8bV4ivwJ2HMMq
oW3tk3AlS9RrvqqZu8UwKTjjyVnWxftYfGE6aKYt9AvEsTtG4wFP3IGg2tDMWTOK
8VbEOzwBBmO1vhwF90cLih+sZ94snjwTZ8a2D0Hlm5xIPcI89mvU0ntTAXC4faEV
wyoMvo812S9OWdLHydZzD8+z7pbiZdQMHyMc8RpuljRr5nOwY4iTc9Prm5ba0X/V
1LICpjMWQiLGu/8iIupFLhft4NGJmLkWtGw2ydOsyi90Z7ws5rJr6sjG7OEXfJEq
bGSdQ9rq3wX8BH+NbabU5q1+y+QBv//mZp+FdCw2eqmm++rC5MhZCWrAc0SAsNuU
KcIZ8MI+08z0cLR7dnOfT30w2JzLgCS5osIPJP5SgGmGfHCL1HXH8aW9xJJhzubu
xffjJtleJn6+SLtxo5Hv88BPeIywN4ndRA6S0bK0bAGlzwmiN5jV8Y5Ke+b2kj/I
EMp4NLOP5FLtZ2V+eRw3NAIugHIkQVbC5tW4W6vPnv0IQVq3j37XfzUtj/WnKg27
PS9pftSYN532ufUQEMvdFP2FJla+u4l06rNXtC1flX3amQWN1o6eoWTnLoIw8IIV
U6z6k7INmGGvKif3wVSqrDTxKOA6S008Kp2GB4hv0QnjI4wuKlSnyAwaIGQfSN0F
EINr0++NtwGxXUrSusGUCJrfjKwb6F2XbKWiEHaYsPykXRiTIcdn9kbZg0EaJsG+
YIJu+oZHwSt78O2FecQLfCvyMEcIURL7jHvkC6rsrbEvo9+oGGBzz/SKqx3f3uzl
GMHAnF/O1JDJE5GacClYD3HNq3tWDCtaUtBGRlafA6orsEhgXw1pKERc733EM/e+
6gz5LPBZt81JZADl9K2vCy/wVk6ibczrui47kw9o8RUyYVp0jiX5vHcUOS3D5Um3
XhhGmwfVGzVFVrjAFP1QCsZMoo3tVoHlsiUooWlrV5xK/S8vK2FiI8W8MjXDK5kQ
vuyjHBwFrnKEbeLoE2GjKvFqCLPMrK55senMewOYaqU8jolhitMNUjTfPywzlkk4
KCIiF2P9/OVEcLTlmZZrLyokQCC3u16c4ofqoT5z4iRt0gM9Xt2HRfknJ5pf/mdf
8JHIEGJd9r+hDYoUKUiRwF0gIV48AOmWXUATCaXnmIYXBH4K5KVdepWxIUp49s1Q
WAqhCSxmF7SljS2e7Mq7WSlhyVe93DEvtj2eFyitaKkwyHk26DY863ZZ3h6fDDW7
BF9DLmlVLlHewqengSpU8nB3AWoD7c2TqLL0jFhgPW4HPm1Hsix/JAg+Y6W2jB8V
hkydHSHTgQAyTisFRRoKDvzYgSJKCFy7OIoS7nFTDxP6h7AZlequgWSNA08R8hTR
lKCFI0aMQpSPn9bIrIlthAqhyUaTMKd39gae0dMcc5RP4DMK9ovuC5fSQs2Naaiq
J58QGGIp+oA/Dh+vWG4+QHDUBm1wsgn1jX6H6aj5QarQ2uE9TbLmIA0mh9+Kor1t
BNJNFK4kquAzQr+AZ4heER0ojUKUEipo4HYLrNhRzTjsf1gxYKwGhowikTdyDKCM
FVCkfZ3W6zyDcpTn8v8trIpc2bNJWRzmhchpjlIwpjYt54Tnfmo03+j3Q88VAwac
lgv+5LkpmE5C0m3mBWi7aTfquxc452OSJ90Z4RkGvv/2KlsdY3iJylM4QEkvFtxl
UCkqvwOQnY1dkGzbu/eP+oHgZT5nipmrUqtmKDTisO9hxLXYwq1S8EDluvX5BQBf
7fTJcFXH1pOk04L5ftIk69EXHWnc8RZVryCZlfl3AQrIAJ4Wj1TUVRcwfAUaTw50
p0RmJK+3ghN4qjTtKpFzZIBwMjjRMfcQ/7YYy7cZSlnd8Spb6Y4vHspksX0/Zuwv
98JXn0zWc4v6e007LeR8gKLBVArJGb0YQQNbht002EZWoljRkSeuRlL84eQwYXBP
Z8qcRG/05hHB2iy4OYELv/jUNOgj3VpBNOFrPxsZMbC3VR5SfE2QXeQ3ocbTuNyK
djx0AwaNl/m/Mlc2atdXlHV8UTs5Ni6GJuTny0reFCiZOSLd3uvS9EEd0FsEBA3F
+DNiCzd2TrD2I8lLNs6/vr2pYMPjtZrIUPVRPxl3ovB/MrIvyE8FimSsdm/5Vof8
SvpRLRT/dB29rDqtwuN+DLrjdLyV9IXEunBZBG86x938r9bBjldlXfRf7rUclepS
MJ35opHxrEN2dhiB5I4Q+u6F/Yjc/C4lkTlKo2iLkCdN4DPBmnLQKBcgPpR9jm79
83s/y4gzT89PUUPgX5QfMYY3fcBR3F5Gg54u8nAsgXThiO4CCOd3cRudlyIR8nZf
uuYOZcyVSnQgslUB3d771+Xy4T8eKVTTXgdE1I/zAWI31V9CXcdyarJpJrT6AK+z
9b3IvC0nFUKt0/2m3AcMhPTboo6AfvD+CdHVPCXOZGTr1w6/TpiBZiAB+XJd7Ddy
SG6Powe7BmgQttHVryLcXzATjK28LzAdnlP2OnPTaf/aEg8zMPezdcUvi4k9cAr5
kJe1FRNBm1ugAU9ivfjZPP8hzyprGZseGJanLuFkTKm04F/b8CwYf3OJfgv6N5VJ
KF8qyAZXtM5VPl9Ce3fFr/ZZG4H7nXDfDVvgkcaJDk4ZHFXuB8+q9CHBgEbcp/v9
s0nXjMTx8v3GCTCst3KpmGUo+0/BsIHmjF/LYQoXe24f/uOB4czla5xz7UxBCXyX
cVSRcidcenUNX2IAXAfjfldLflHnGhujNUknNzoLQThh+M0hC8Y6rI5vN+v5pkxC
AIA2Cijb83gjc+2Yb95lzMVqik80JZ8m8je9It6WkBofVY/h6tj41sBNDmx290ZD
yb3LEc+XdV8BDQtFBTGrjAydnS2Qurwf4TgXCxhjt3ghBVF5wVwC29UOv5UXa18S
MFZGOIGQMMvGtLk9BvLtSHl4onXeXyzDuG4SJof2pfkYjfvw5B9MFmJVBSsg89tp
B4rN9bOyAb7vJlwkDKyLDOyn4GSk2S/AEVQZ86QP109VKpzLly2HD4crHfrcHHki
wDNbwUBhaMn1fE4fpQNs0Yxpr4mEx4p7C20cugWi1ew1jSXNEFom+mqkWtsfoAqk
HpFGQRZ6RJSjeR2ci1TMnQm1nb9IBuO9D8AQtjzysJkfssANOV4PyDMvUPPcB0wk
ppLsf5irwSfxhDN7PuNFxkXEo34qJMQSPdjRi9R/gJ949P7VLNVS5Dk5JD9MyPLQ
zQqcaIOWlhj1mcbF8IR3KSans0h80VsHQUXPRjcn/TQ5Ei9NBIUsupWST/knTnZJ
3XZU4YjNJJXEJTVsZrmIkw+F9u5+tGjauHrHHYmdYQobEcvLZDUnVWty48cF9XUV
UZMeD4LJod/q2WQnTHAPVSZIkLqDPkBS1lmWoYBUsoMY1tqobv31Dcf0wqlDzJrX
2GsPnobkx7VGWSwUgUu3tgkTDiKFVHgRCiWsi9xRUMTmWaeAW7S1rSkdI86cmTT9
5HW4fMDr8083WAa+7X0H3xmpFLqVgJhSj0YbSNQbaQbID1sEy0bhnhTlC2vHA2HK
xj9pVgEhIevbuEylqWlMXNCj8w48fSt9xlkeHOgKjIKk205xMFw0Sb9vjjYRl6ga
TY9mXUd9Tg0MEbpx8WNkkW2TDWHW4327RFC4re+oWEiNtiUut369ZEheiPAWq4JY
8hxE6za9fJ0j17NLG1IxXD76Icg2n/yp2jinhnGYQo1mvEogNcOt352KnJXf7eTQ
goa6Isvk+SJxS47QfvN2rKWLyakUMJXcbejZdAmk/Ch+Ill1b2F17q3g2RiWEJIs
aS8lB8l5dKtDNhMw7gN79wCanVas0g4fJTGCOYzocoZKXUP9a41YXPTDOlOxtu3c
sOn1Ak+EHDElEgTmySLUONVg8YXRz2iAWXujcd0NCeBg/3leV1sYiHINHZspmbeM
z8nouGeumAk5GuO8+7CfUOoCG+8sL7hIiRR4oknIRRT4Eb30gCC5i9H8VPTF0xU1
5ugG0END0dzRJJMSbsaP4U/qsND/6L5g3+3FvWM+FtlpB9v4qPvjftf0QATVzzEP
efqlri6XzXHhk/eOMJq4nLHWc2MQJ5r4EGWb0w83d9vU5k1r+Ly9tjw01zpbZKyo
GWf4QuizXw/6mVNzym+R6kkM5p0wedPKrw1omffOTDCEfaFiqycDejJ85/K/yeyZ
BarJgU+PIqJFjUJgkDbztIorOvxoiuyNzPZ4ywl6MbpQuRmMHyuIz66MmBZM6M8+
Ppm54z98AOxs2Pdi/lAUGtVWsNEhdCuaH8Yor5CnIG5x+TxB0xN7qdqQPPPEJ3SI
IZ8B+als6vxrkhkiETfVMdHyRNjE73zpQoqcYaSGt2rDgfCJ3EH+M6jQWbB92mmm
SkRiazJPjdv+jklz1hJEDZSwsT0LfSLO4mteRP1VyF8jNY5yjNo43WYwOVM98O7X
l1yr6RPCZkqQ5isu8iyo9Tl04fQk0Zzyj55qQV9i5MWWAs2wAmALYUUpcLlGh+Zh
Rv+8cQE6Oy45o0TC+AkQyanKk+eNtu8R2qJTsN1CPzW4/m3w/7A4MJ6uhj+W5/ab
48ZFUn74ze1MULIDa+lE3AmmnRm8OK+iXMvpAvTVPNf/5AC9HpCd5NX3K/1fMinM
f9hPNSh00o/jI7PrCrHDExvOya3ULJAy7hWLOj9v50GwZllFkv9biZpgDS0oPshB
hpoYKscLL7e5GLJgbt6v1jF6QBmKR+EOv43LuTjh32n5Z6NSN7IBaFgmC9rOyWr+
R7KCyD0Px+NJQzVFMEyym1w1DvlTn1Z9pwPrb+f2vLJ4E7URgYJEafoT6tmAwIOB
mbWa574Tdu2ML2vD6hbGC394UqipZAkSPbFwu5CqE9YjYsKYPPJrhm12I6hyglzc
OsoJ+q49rvzFzfk+LI0oFSfG/AlCUKtin4JYO1cqTKy7SDGp1ktAquzT23k2Gm7g
H8Q5vgQb5Ry+yh5GfOZmhPlGUbDjimGJS/FQYiM2lAzHC/gaDda8QydNxwitKR9m
qm94GnAAeBrjiZkp0+O3txNg9a2n6+b30zobUbVICaCxhyGML9BfaJ3B8HBZ8Jre
e/nOXPBepTXF/h/srxyPYYG8ZS7nLWtMbq1lKpY7T4syzkW6W1gvhQcVIvrQIUEc
28GlMm4mJPpObfEvRuhrgFBV0C0YB8PwWrqZcHgEoKe5kkg+pxPe0JYmB4prwDCQ
gVwVioEcVgSyDMy7apQgi+gJR3FoDO6L56+UkGFw33v6VQ+nYxDWiRu9dI5ySRCf
CjMNKrBNOa+fYntiL7E8C+OBjiJp7mi13SBdSCgMocw9OCDbF2ZIAfIEw15Tp+ff
VLkqFu8EKAR2eZUzZalCiMMptuslsnQ9/+QgtaIOC2A0ebvKkN6uwwj4GgvZ06iH
o2XPk2nQr7cybWcB4zdgnivZ5b6at9zz0h0DrLNkiUbn/hALSbhb6mVg1czSTfQo
EgRx5XCE291wcpZf6qFUPMq2tKbNYUhVMFPQi0Z1+4dOGknhiXj4WQDiiRvw/G/6
uikGqeUAdcTQtUy2MzHoQ+xslmg27i9HeXhyaC6eh1dOpe/9FZNJyczRKEmhHD2d
FKNP95nfplHXA9Iu2DASg0XsjEfPe9im095wqrmQ1ERN05b4BlFODrdCS2jii1M+
qzq/ncg0N6bKf5kMaEute6Zeq21UBelKUrWNq6Os/E/XoUBppLdMwB/DQf6Upz7Q
z742XHRzIlgrwYbd8oJ3hUuX2wqI6wwgMvz/e8ZcMv3ox5/W0XSVM2+Bv7gkl9Ns
HTd6GQ8eBfD/a8D/9sPzfDEsuQO4ZY/Be0ztejqRSKfau4rbL8mUtr7pyuVjc0nI
5hP8qpEzy4pkOTxT2VLzFfCwb/DGxgHASD9tQWxalHokydDXKles1VMP1fHTQ9Xw
fblmgLYRL+R6uj9iJm22iORYrWxpn570V9mV9wzcWZVZKwGzBolXs38X54Ju3HCC
17Yy5zmsdQYZxkaGrFdh8xIXWg1RzRVg5+DOZhNcyaHHTBntvZDiAW9t2rRgVIhT
V6pYF1dc0nkCRWWVGebVV6Sr646J3zdYarZx/rdxTwZcLZeDSCIHAurv8+I4X9VP
YVDECrSOBTRE3HCqeCY1+alIwiBl6/EWm8MsGAhqtqtfuHXlni/TxJZvlE3AbuZq
i98zSuksqGjglHXULXAq16iEt/w0ve9wN1vSL99vceSn6t6h4gWIo60uJ4DCOw8d
sBEScOfgHIc49par0nDDbba4dI8HNlRz6EhXwcPyz3nl8ptt0vsu3lma43gAOQAy
+IVtWv1GKBr4w1YefaznL/PvEplOKKpcYVWqXvOMhj1jbRepzxAg0u1kqMKetChL
wJfl9Bp4mhOSYxHCz/gPWXO+aw5DX/aWZuyshfiRrIiDQPjHnWDKjlNQsrsd3cz4
MARQ05ySaYwvrxssiocWsE7c97187sWoT81i4D0clzMxuh8jOGXL+4lU4eJXtLeY
RUiydCRpauTzcwiAPu2py95kUjaBXbe+Sa8rB0RO726hE4zQHfWZlSqYv3XOl9ln
ySPC/eGMQO3VWEtrY6/guhCTyfGWipsnzBaXJOLo7u4Zh9zhqntwJ8BOINUfyTuI
mBkQnvfLGX7ZRK7LiUiBYMd0rcRisvacRdmJXtw9kkvfdCvlnotwV4Hozxs86v//
AJz5KLVIZ3uye+8jB266llNwp76a72eN3SKS2GFeJ1HH9tzhgpPFcDlFCvTW1gRG
IWUiohMURs6zRqPElCrsG2wniNkiAUqlKLZrPgqfw9D9cGbAAodFxer7uEdKPdTv
ZqUF8OZolEmltoDB6VEBsOf2uHpoDPGxzrhUm4hQbwQ/Y/MmTTmh+QbkgIgQdF8w
sMPaSYJ4Q1uWTzkmVsdrqf39K7Y/eB0G3cWK+UAkHHih6+NEWvovsJVuE3THgwzL
Y01gDZEi1J0xlj4YAOMa0Xi8TMHU+kET2WmUNxdRN0VRZAfwcts2cIFEj01c7Uf1
QYELTo+LnCC2GwdbNbePz4eq5QHrC4bSvO76drcVF+sMlQFmShUdn9tJl1eL1Qwp
rsF75LT4FXrdXDxqq7glGhiGcRCUqc7vFOtVIEevhK6XH1Yf79wqiTEw2Dir1t41
SZmM7eUlRqZ1nt0mQlTTi/8n/Trg37x1aNYfSZNXH2yFN/vDB06VlYWsn4ywJ7Ss
5ziiNCxv4LZSmgmFBJjW4OLE0HA/VceGPjT7h7EWLCwGjgEPKSVC7+EgFYzspERc
BzjWXi1yDpRPjIDSn8kAz9uRbFrFuhS87l6uWTceIq7K7XPaT3xpHejKaul8aVi1
udM/hpWtrVx7VVvy1jHeF5ypuUylAMdow7ENE9/QD+kGmDEbgZBcvfxZjKzPV5dQ
GCsVS9O9Zx7TqwFTmKV81BgFdyZ4rKro8Wygnj4RGpSdfZHpLJHDDnQuQ2c6fngE
o1dWbKJmeii7bInjhGw48a6j+73ZARMYsJk90HWMH1AaYr6JFG3w+KHsUBE/1Nt1
kpGOTEJoNKjl0c9AubZ2VM+5yJbOdPZ7f/rBgJfJdccmkPV8ZUnLbioqdvBnd35s
ADsM9BN7m7EBa/8LrttLBDD6yHOVH6ePfViCsK7S8IYJITWPzZq7Zb6SbvVIyuCY
834XU6dZonRROwZUwi0oKpnBguwwTXInGvsNXYz8Mg8F0cUL3nUji1aeMvgFNuso
Kgx4OeoEXZ/drILvtBf9n92i1HTFUXvxTJG1GcmWRgjt398Iyj119xQ1CjT+h4KY
BtqGFVHV9xMl3eaoWOvidM0VWISU10VaKTLDYrJ/EY93u1YaJraKjxIf/js+BxmZ
3EPLghlqahjC3RhLtMmR9WC2+9Ak41vt83STd8upIXUefYCnYfyZQotxSNvaUKji
Gqbk2E2km5SMcnptpi1n+yBuB8jx2uwHKX127f77YBpHlbVZ1Npy/gW3rQbBMUqg
1YPI184z5enFD1YYlJiErvh8vLblQrAIoQXxzCBaZmZjd3F/ycpT1Jdu+RqP8pLp
mIl66VdCvF1nPvjqsgsnCcmQ4dEbES8inyjxrJfJvOM6niVIOOzmKGGInOWAn/3x
jZm2Piw0QYNLGr34EjKXYo1YAyw5UcK4bQNMK/Ucl5rQLc4KwDar+V+7FUCtEk0r
+oYH0L0cI0H+YLvyxzlrbOOP7KDXPCo9jyfXzFzokAM097CPAuVQCuJMLiIlfyK1
3Jp3Ms4yc0CXXjxOXip87AD8aY1BiNzGmy8mwIKqEFaqPtPHhKMyTrO2Yz2oUeSn
2S/8naX8+8E0LiDcb1aQZsT6vdL8ccSYQDsewmVqIXHfr4cx2rjkY+P2JknSlgr+
G7e2iNTY7WTYNtfkS/ovoIABEiVdjpuqNTzX8q3qb3h98GdDEqkPN5x4GzqooPkU
3YLBahBURdUCTo5FtKyr8dHnqXnS5wKc5E+uthJdw1ORKrhwlZCDyWCYJ1H5AabE
I4U/rOF2DIqtsohFHCWPrqir2XeEpfAumWxccdw9fqCGJgEqazjNkt/UUnyUcWCm
O3DcHw0J4T+SSSkuU4Lj8gvvVyjeokcrfLps1Qd9iTc7KHbnJq2tlTMpVh+7DF7L
UInLLsLTqxzz0I72QrdCve30V2rBvFAfgEY0TrTWRkizzOJ0/q8lGXvHIbY2vYSZ
ejLeQEMNO/e55snC8CFOapG7r+byPEYB3hX6GBsFh/VItmiK5rel5/XzH7vKmH3b
kqGjEwkQIIHvhUYAAFP8OxWeOrDvTSwnEJR399UVSuob8/j98LCbUDRN/L3AGJlS
6D04s9/KiGtuM3u78c1Dwi1dtsklw98M2XHN8eAATYb46W9/RfvhLfafWeWhW2m8
lqOEP+yEXqcYEo/jW0Bv4pBEh1YgkPh5TjzkONKOeTkTTsMBE3y/7QViTpBiZNso
HEMJX2bBTUFn6hBgAjld8QhqkHnVn+fOGHk9B7NRRKTm5zrd/mVTJ/jP6na+tG5F
GqghTODGX5Z8G0s1tJ37NpccArQdkmPMbwFsP9aL5Q4uBRfx+n9cUmQ8ZzhG+1JL
p3aqcLEzoLo57pypWCKWp/4XWgIMyARKmyffQxw/26uhNhVuuxDAx4wqtnqIDpGf
0ARa4FyfoAvBJi6JFVnvXD78rECgfNCx+/kkp/82zxw3hp685Bkdc8DDZHf5xvla
vIgEcbcAwYqj8HF4zxgyc3WtHd7R30WhyWLncOPlw2Q1NtyzzB6cGKMR579DXjYf
/3cDde8UK+xwXuaPb2iZvb0hpex2m5TN0CHjVltleaY0pmJz3dZY0d7I1n0GMFBB
Fnx8xnqv99XhIKusqWvIBv6+bp1ZapprFfgIgI5UnMeScS7sxwDmGrjQFLAPPlP9
wKAcTM/QEeR0LnZ8ummqJsiZ4FViz6+j0ZXhIgCc7+5NlwkIixSL2XcP9I4v/uvU
NMaktzFAoux3XOEn1UeRuiQkK/ucjGST4A1IK7tZX9MM8e9KxeGzOzjY9gZnjhl8
ZX/RDaOfqa96B1jE4SqpfT28UhkOdUzi0pUCijFGsFHt2aMHrUwKUcuvW+vDSVDb
P07n5t+57qEddRAm96q+OPk8Rfn2W9ugFnb+v5IbdXBQbvDMX7VjU8MwIAZfd5w+
UbCUCMX8QkdnLmkfS0a1IKeDSpWN054eBfQlnfVFvXjfgAG6bwMuyjhggStSYYQA
VBMVS354IB0Y0qKVE2rV5DE1hCnyCzqTc9AOWXh4fDFHya9nPaiWpUeJ5Fc/gjdl
09scAC/QXJAfBNpR5hruzk0hWluCk7KVnInx7EKf7iW1MC4GCZwk3YPVzvbQH8KD
EI6tU+IRsEFdFS9nj1ylqYTcqlkZ0QK2xStMRvmAzUvDcpjqs5ET+CvGXr4UklOE
0i3UIgdHGUQxeIBCxobrsGzkb2EprpeFj5vneK4XUj7HA4EYhSeyX6CYbpKoKXEA
a/nxiPSDmxs3utqQPF0mNGg0tOR2H5ChDnL8b3ROTbPXI8c2Cv5Lw51V8Xthd67H
sgSpsjgTTsy3sOox2ZUkrZhcpLA0clMRXpTwzVwD6mxy12pN0oEl6oSa6iJuJCK+
1o4p+g/Aszw7fWbX5YTKGGRqBFVUAxBx1vIAbxdJm8hNU/vP1wnp/X1wdfgDVeUB
i/y+fn/7QTwJEW5hEPgLDAnQwLWCPA4lvV1GlrDydaPGUy7RGRN6KJAMUPiH0A1S
6MFfMaEZxeKfJgBidGt3KB8o9roAAsNPeHss8HNCl4DG+ZJiB0roHjTag42QwbQJ
mc5khKMZUOLjFhWZDV0ge26NnGoc+QIIqZVlmuiPiuIUZgXxFEpBiI5GE4ccVdhX
Znxm0xV3I1Uex9kUCzA77LSguKG9VZNdH2Rm70nvrSpeFgpWXifZqVNyXhr4TZ0X
I+et3YTzifMfi9F7QNyV5f6OvXbI5Q0FKB+/6sy+ySVjtHN11yDlZ8fk77PVHW9/
l9YSUlSwWLLOYz+RypoEHFfhGFQptf6FpYinMAplD4fPKhvVtfu103/DwPAi+Fk8
KQGB82w9hbv0/OLFp7oycs1yjGgr3upRlbhz1vt8CsAtnuDsnK6/SEn0AJ41EVAD
ISgpX4xkY5obIDRco2frMRlxl/RC7wkFBGIlkpXo3tKN2OYrwAxgce50GjyUZ4JL
thHaQ9gQ6n83FqxT2xDKNT+NxOtBav+/Qqc3TqLaP1HfJn4zpDPSyzE0dr+nm4Tk
eDITCc676aBETOYBtqgNN8UKQ7uv0JKwwg7gd5Lo5AF20iLkXQaLXt9ugy67Rvsk
P8hrdR/EaqpPmOcOGM7dlN5Gw5nxfO/uVXPvzFPahLUvdmk6fg8N8lpluUJ3jUDv
RcrW08W067iRIxQcMZSi80jbbDgniawjytbtW5zzes7qpJ1au2fnRv5Kpo2Gs2bK
ZRrroQaMutt8C97Ga597X+AnN/Uf6OQrewe7aRh6mJohNPoNMJ8qMT1C4WDDdrEu
LY7o/ncI/Zbb8PFFJCv7+X8SFruQkVy/8KsGeO3wS5YluyCk9CzsWGgJyv4/PwwT
4/ZjiwlKnebEl10NBjmV/GZVrlY1O7Hqo1Xs0HG028QFtecC4l8fKcDiZUjPnNBA
HKTR2/kGn/+15u5duGu5HEmiXX8bwGWs6INzkWVnZGfuzILKbs35EA/pHC5hw1pV
WeEjYJHKRhD7OBmWxGgrYdjWKlWFjLgjfzziOg7S9R/4JfwnBtAyW/zl3IIbO12a
GRfiUvdxW9NMPHG74xLx6BQmHr0CxQh3vOBKwG+sa+kTBBTOOfkUL1JhCgEqyRlf
PslSfaje/kn4VXqBGkr2eRDTmH3H6euZIZ2RsqeXlNBa5PvX+krY0BQGTqGtHUk4
a2xybpcKbXHZb+SmDojQNckViC5egd/cD5jdtB7Z+JT+ZBfOR/hk4mp7hdDMItF+
TqfSWWuUUdDui+WPt165ffZnjpNUkiIMnDxNPjQow2zoRaxFoE4HitGM0EqeGbtx
QN4CX/4Ge80+fTOsR7HnIE+nn4AcgQDm4rjh6A4f1pmmsvAsftxUqe3b0+H/KgMI
9SVzgqIOezR8w+WvJZHCOdTnOKh45P2EhP727Yunb+I1KWBhYR8pum/eN69TmqDT
yhEvFhTs/kfPqW6zqi1Ihgc4Samj4BJhRDB8loC10PMVF/+dYyQF63qhXNJjmHyu
BHgdLCdbeh1Mq1sgsZqd3V0p26nisqOxg+d4jee30EB5GtzJ3o5cACT4OYrlhiiX
tF+QI40WDecq8QM2iYBsxtLjBe25fwQAhc6zujdor0wQdnpJ1kF4UZhUxKHAYzWZ
YCe2enafkubgYgDHHstKPsSSs/e+GTbl2933ciu/qeNwbgRupkbE9rs+a7MOCaVw
X4r0B7Qtj1B34aZHlB9V+2XM7mQZeb6wODtWntgpJuLRmSQ43ShRlrd+Pz8Csb4Y
pD5jX6VOXHrZoXmXe4HQ84aKsB8p3+YdbVLshUdOZPWc7jC7w/PXtJPEgkR8OaJN
E3PAQYfPSwGoCmNKsWrUMdOFlH5/++xJB6hq34VUj1dVS+Q1yjN1v+6fkoCNal27
pQyZacmymRA1FB7bg0U0lGxbLhtiqeXSHentgO8LDmOV2w3pCx4WCkwcAqE507Or
l2rjMk13DyFdvZc9inZqgZIzhhi1nCD5N3egP+D5nY4lEbil9wL8EFpcWMVNkmBs
UDwIy5mZore5ihBpOsxL5QHHvD5a251gy2mDS+e/6Ra0KwtSZmv0Nra7/sAEFqBZ
P1bpImiyV4mMokCmxdV4mXbcRe4Y4JDwcyxsRoqFhHgUcZlS3SEs8PrBxz4dkkRS
YNeDPgMREym2VyvvWyoZmZ1xrFJG1vfaZ5JQW12yo6h7wke0lL6mbO21UmMb/u+p
cdFShPELaLCra5LToe9AtAjLBodvqWZJ5XJ7TPLbGVFZ/9es/lhFp6FPHWlpgWfH
YdVHQhfUttGBvkaWAW1tpG5uleZMxq05OJBKkOHSc5lZ328AOsZeTlJ1aGlPOMV8
oixMxkysj+nU5UV3AcMff764gas4Whn3CfAPmqGjBeoLlh9majrHIp9UdaSL8aqr
OUazRxcYm6eg7oGFEGVck9EpoufhwA8vrS9oPMP1FAiRkmUDQcWJiwwd+FcCIvt6
VTGAfhAQMOulOFPOFUR8riZo8tJVi4QACk3EfxXi9qPiRm9Lbas/X2oWUs/booVj
CFQGSugjNZ9YZMYGf53jmHwqx6TaHKdWmp81VsLhDU8GWix53HDBeZWNC048IB/T
yAvARZ8pBWju1Eb5Il5s8/vFbj5SAy73pQUUwuR95Km9TN5s9ujr8O7xiYh72iUz
/DxMfc6lb0Fuw4Ub/fSSF1QxuGL5aB4a8PXF2Bl5vqAOgPGxaIYeVPIRZoFVargc
g6/9178+JD1aQVjBM/TQvGqDlFMfisRM0Lk9uRWc08bgGpYxnxlfRP0XngA8B4bs
UwFqLybdSM1PMz++TkXFh4pYDFGXuiM26bJ6ymbUFgtHp6ZDLKW627SQ//3BFT3P
smmgsaHUXxhAsm3ZtAQ3Qd+BAE8iXs6uP5uN6KFdXho5eGL21P7SorVvR+B2P4LN
DCy5NVIvzWQE9SqlwIzMmve/t9mTzt6O3io05nThce3L542tU3fEGuaRpos1hlTS
jXxYvVWS5pw0t8y8AgNhi164ODhN6O0k4+yY9a/lVkIibxz8ra8CMTTF+etdC+Gf
27Ke+fmT37glTNGg7TdKsDMiemhsrVsfYPqZYEjKVR8m1UQpeTUzIMC/YG0nkYQo
YQqfvASBt6+aAcY+MVyAkFNSckkd2CiI7vCDIz+ze/cFBm6PQNDseyyK09Ofc+ib
mntOvtTn6fnNPPYsqxnqYihWOZ87L4d+8n5iKI1dr7H+B7zlYXuB/ECRgJe7w/jv
Xzg33RDKpzjOsx0xtWFr6C5lnOtyjHSILIlByhw33hgBKtrTEcsxKPICvntiv+GQ
3Eizca3PvTwR6VoYO4sJdPHI1StVta1EBFtkKtxHu/ZdcApKHom/gC+RYsjMAUls
3KCPFB/0lcQvq8aMJVrt7o30Be7LLm3FwjTkKi/qXAJHL50LEd0Fj48pd1SBxXg8
MjK4b+HWyYSUkL9kY5JGlr+F24RKWOZx5OqzkDzA/uZ+L3XvnVL3FpdvhyFUcQrg
MT9NqFs3BZv3mZYhHd9AjE3CIV5KlvtCpx7qcLX/da2RxSQdfp20Hn8hSFGql2nS
LOC7b9NdZHumnz2GmTZpFn+EkkrcM73NQNUQ5YUON3G6pb4y5knn+kfnBUpEnxEW
CVUs/aQd2kp4gc4NPlKbAMfyd5nmLq0Zs4MHlcspYgzMoQbHzrRn+G0dgBEwbgeH
xyktWxtZ1Zr1Uqe/21dzPZ8oghl9WdrkOekMLVIxqLUz1yTxVsk9sIPubaH4AKzf
JE0JOnIkY1fjJtRebwzxSemTmgqc0nGODfLPMV9asmZ2HAxSTqEDRwoY4I57ReaN
V11ua7VFmm7yNHq0Bi2rLoHFdjqW6Np9NHi1xe4jEPS2tIVRCFgE7Ve7+di9LDuQ
nQ+KjlV46Dlv2e35IdPeFh/b25nMYlNYVGCaq7zzmwT2cmyv5/8QE2Y+x4RkPvAa
OndD6VotVfIh3WLeCxmDJNsBvb0VRVet8TzPYvCWha1dZq9p9b+tyycB/Vj7+1bk
bjhFookm8wYwZ0XA2Dq6xQPZOLc199MTdMWkChWnF00AW8ijsrHFXlzDjEiixuPh
arQy+TGcpTCf+6JRzqnT8M2RRv+rngztfKew9/AGnHMEWoHtQ+cLyhpepudkYV5E
ytm4YuvIF7H8UXDT1Y0pUgg8mqtzU1e3tA4OzoNtgL0E4O8CWDpwUt4w54TUmXCZ
dutF0iNZQBWE9N34umlFRdkEOOzQKnxBqPQQiQ4M59MfaL7hqpddNWCbPvkt5d80
yCAKUfxiB9g/TIrrOyUQTGb1ZNsWAjwM+tLHzNKkdWfO4IuRYyVi+ELYg0XDMLTd
dAy+c6zzZ8s6VElBbJjo1QqcdgrexE+UqFv4xLj/0/O40aAJaMQkaBS2craQMjM7
MQUHfnoUlReD3SN/ktzSBtKsQp027/d1e+a9osfZlKAceqWwVOf+SalipukMJsRq
0SLwTg/mydSAhfMzIjrUJDmJBAe4hLeWFdJwrzRYiQp1+ara+u81yJQGr264E1V8
3hBdyOBQ/NtJmet/2jyXH1pMrmeu+x61lQ0LTdnYWKgZijhwpy9og989TPDd0jI4
CzXcFuSaclHERQYY1270par4hi+FgrH/iy8TN8iW/XicYrv8KezlM66DjkBY4eD9
CN14C6NK35kl+L0nvqxHsGiHijpPtZyc8mCwdGm/f7mr5NUc3E2LzoButp2MpeoQ
TBVBO8hEU3o0WQ/XNbXdR2i3SAsuglUvx5iVwnkVyG7apBorryk2DsQb64Xc4opx
MlIPs0cR43g1zqLt428ETrawPJlTTzF4eY3rmH51RsqTLKqCL9XcUjCk4KDak6cS
ZqX5NK0sm0n0s12eRO756ZjHv+bQdmP9Qflii+ZqP3ylMUg9MnxpDcfHO9gEQ77M
wL2HBcjiDPA8ROyxYm7qvRhqtnSvIB9Agt1Ex5D5lbgl3uHf0hj5gm/7TJh0Xx5i
kLBoik4Lq9WuhW9qSZ/9I4YP3lFZjXo1mDwM2l0IxsBE4wYzYGtV2m7L8NIJlUtZ
4AjYc7H54FANXWo2lysolATA8EAIZhHIbv97e99vDMv4Go5zHaTADiACmaAoK6iq
3t9UkU96mt4+xw9Lpu8xD7P1QQgcfykA5/m6YjkfTgcB7k5FyxsL8rOa3b6CENjy
ePhDFXBfsT/0To4JZZBe5IWQmUCgwvBGa846vhgrrZabS/uWNTGVDYHuKx1V0QwW
IOfr29K6k0WgA24+W10mxLgmV0ACnQ7SSOtCmL40Vq2k7GLHiFS0L9X5srr53LAs
ya0s/5oBtdWsq882tx8/g6p8zk7LwRQfPyJ7ykl975NZUWNzfLvPLSUdSafVf6no
tgsWiVcP0R3g681UX/SltDb2kJxgxeM59zKtbkksJ/9lchcilAy95viPIQ5ksoao
0IyMdy5Fz/MkyMlFgbgxJ0o6ZhwJ38bryuWLIzHUlFeNGxezvoZUWEO5tlszL1Rr
zKTb/3TBH6G0r0a5BOapYMWm40vkcFE6feb3pUWdBoVDjIMNLgNR+4+2mSzylOk0
uZjc6idSz5uaAI3ifFfJgPGTx1E5IdjJnO+J1JnV+phzH9xf60Xb2/ofiyBiNeQk
vSsk1rpj2HU0SyfaoJ4avgS55w0/fiXlcCWxByBIcaO5pt2OYsw7NuVkqE3uz4cJ
NS+5oqXNuJPVm1pk4olSxL/zII/APa0WqRvqV7zr+e3akgkgO+44OkSNEiTEcbNl
EmVezLW++fV1bfYux9u6bco1wSz8QzCv+fF3Ybquqz7nOQtziZmau3TEDxpcB/Fu
o9JXNhuiWsCC1PhpjEm4EM/WgKAMjXxHwH+/cY7ov2Qb7e0b3h5A14r+0vbxmQM0
T/58jQ+cChj+JJNRMV1EbJ7NQru8utb2oEEI/x2pIKcze6zemNbVgxPBFwcPeIBt
LMClGRzHvUrBxjbTykueA9oGktA3+IpWehHu0CcOToMJGcwvOgbAJOmvOy7RE2lM
CkiLbveoJR4j9haYyFERqYrNikNQVLtjusiEVbFG5vpW2dbZdIT86v5Ku4suLo0Y
meMvMryACtGGr/dZLcQOLuAQoUbLNDAOM4Bs5Em9jq6JzjcRqoC7kVK8p75Ze4fw
IdKp/Hrh9zAjaOXArKiLKqpyQogamNGTZ15UbqI6DTy3CRAfPTIyTyT1fYB/KXP6
UQ8apdZpmsuSXZgCqF+hOHCIhONEZ+ceFjOFH7Cnhxg7dSlVlCTDEwRdXlm1kykj
8gDvTmHJqTAopavTAMRusz5GfY8dVKCslVhKUreMW/XXDQA52TLifkzpuDaI56Yi
SL3agOf19fhYAERCiHMrGZtPe79LODty1URoZ7dNYlTudjajao8L7kyAnjuTeWBa
4LhpA0IuejYWzn5F+LfcDqsHr/ozTInZJ/X9kmVFhdKY/AcZ/rqsi+JZ5BLT2qjr
KH5BjQCYWxbC15ZK9kVPsFlj+CWWenfyuxKm7HNlm/NWLdae5KOq1c8e65eDbBKI
yOhQX5AR1pdN457IbzmMHob962/wmEUfWRVmCtBJpzZ1chjJPaEVOFQgerQeOY1R
Yoa14N1cp6q52pNf8CigJYi6NVp0qqo0vMryEhI56ALA1AjXgTwZhJurNYmRRJhU
zsTXou8hNMU+1anzGM+VZmv+vcV29HlZZiOvxV9Qib72xLetdgUSuIKmD9wMbud7
Nl4JuJ7zr/43DmkkcAoAB51no1trsdZi5pOB6lFuNUe1ztFtqi3djW8J1IYjC8wW
MMy4IjJNMRjEDuXK4BcksVDekLGmv2OQko5bA1xNb9llPSi5lUhby1CY4b7eDU73
XVYhKDWEifqAlm/sKQV+1bDSTucWGsBlupVhrzSo9WUCfRvoR0c49AWPrePi5u+5
uVAvxR4Bf/hjVuEMFVV4W4nsGjOhoPxjPx4LXpFyu1gCgfpf5/ST431JDZ8DssBM
IjmmiX+uTLx6hWhi1NoUKaQhPUPi8kjnEzSwBQRzRWM504+AvKRUCuAqk198cUqa
LC/qS/zWbx+HD5XaPS7/xiV3wOVR/RKTabF/t45mxVfQx5VWLlGj9b3TCYKl7cdQ
hctPcRENU5yMmF3LE8VEgxS6wa77vfaayMDawydKm9w5xDmeET/aJv8hQ/JHvpo5
+Vdc5ydIFSNWqHwks+sd5H6tZKQjd87C3gtuqtniw6sptNh43FMSsota64uxPm67
lYKNpzgB9m+MuEdcoHi9LSnNwyu13xJY1EsivSGNBH5Yg9MyyYp7ct0EKABf+2WN
PLZ7Z837spXYwa30+WnEdpKUE7RjA686aszw1VEG5KLsFOKZ6NiDSxDTO3C7eg/M
h+cYBzlo3/2RA3C6FzzzoVWajyw1lAa5VtH5fZrFhdE+pg2h5wdFi/18lCc7qJxa
wvCmWGXLvmg9FSe//HLiMdcLCzLjrRlKJrExSJ1m7YqwaSqX+PfCUXUZbWpWb0WC
L3CdHbGOIs96xnu88euvKPE9GZ6T97z6yKIAdHUMKZhwwIAhZ2oQfhuNYBrYKCST
qJ1HyWCkMH1w/pKatOriFNlTnJacanV2VEUVvKNw9x3PfZQuTieCg7h+I4XVQTeV
dutjnYzkPsCxkKwAgHU0oSFEfhWnR7mpVSX0TcqA2wqLoz0E/34jY+24KkqNnm/S
CprieV9kxpDc81g7w1giS3g4SmH/Fln/owGJG/141uB/JgHIJNAQWCCLnwl6GPED
JxmTzHw4Vc/Q61o28bda5NWELG6CzTR4E49XAkKSY/9eF5cPsZoy/ZCtTjRlgzMe
pg/weY0CxM5k4TU8EDSKc4OoomSHDRGTebAMe/uHcD6waQUVh78cQzULtlioh5DI
UjumnHRQcc7qiZ73RLBUFmYojyCPCYhBttT1YJsYMGwZbP5cZiVRgA3tCp1G/oki
JQZKFmJFXQEcg37hH5b7i/vYzqEwlA8ooW2cwW3gDlsFW7pvCg9lgq0kzRQkF/ET
+bbXcopKQOyc0f6pi1mPmvmPyU8DHhGmZ+J5rX0BNi3bkYMNoYuZogoyf/1HzdG1
2dQC3YuOdWR2R9ciK2rz5gMCAEQ7233FjrUTjyL8e9CHQeGvXmUl65WRTeI+TDaX
9xlGkahnEaa7AC3xF2nm+obwvnkOWpa85yUWpo6pq8cJRNrXt4qKwXcVT+Somwpa
X4/pdA2c6jUzfpyBwt1aYQeHuBaoPcB9P/nBBBEAiDUSPzctzfwdrNBKTGfYma+J
0ALulv0J/s5JlBjnWU7XQwGESoZt/qaet/QXG59MpO9rP8BxZAg8vzBZdhMZZjcI
5X8ptZR3Sd1S1a0Lr+Jze975OTQq2Lx69ltC40PL7opWVQmDDkTCArI7QmjUQYx3
K23zrByec3TxG02kQEziKltVNWKEMVk8P/Cso20sGNjEkIw5BmWe1FJIGi87Rpqf
KbQN7GOx8JqhjJn5EbbE0tYAtDpM1CEBVUq7dAslW6xsqvcpnkgopmCfevEulZ6N
ru0am2EHMhciWQuwoXyqf1zKROjtPmrNukWDLBJ1BxocEo+/GrFlC1ozu8SI/Wey
Tm4LFP40IQkjXYzvCD7tGXq/mcNeYEgbuiuBRn/5LKH5mNyLYrj8hwVzyPrh5xCZ
oG9DFlRAtIQxRhlCNxD1HjvoqotJw7Qw6gTBeBNJaAPxQDDbKeu8UxfcMGqW3n31
qqRc/pu6RCZVmU5f1OuYLJUfbgBpWEMT+CcLQ2w+nvByXiCx6YOoLb9fZI4cmDAP
mvNtZ7W00YfFEEEaKcrhEd1cFJSbCNgbNAIookoIGjp3X6Qtx8DnzVOT7QVKCSaV
A2aDMv6BuLcoHf9cKg0SQjjwW3dmPgfRaGKT+5iQtaIQs//1+RjTqLH89CBvTx3M
acs/9bM4ZKSka7+V+sQ8yts+B/UiGEJnVE1M2+rOsFaS+a6cOu1Z6mV0SNWlKExj
A6rfwsnoAKyxnLwVu8ESYBfQa01oTfAhBR2Vr/oygtG3a6BGStaj7jf0vQ0ISwbM
csadmzgCoo2vYBiYB/0EONSsRkSZqc6r3/+RZVnfc5XVq/p1mchpzHn6xjhY5YeB
ovrir36P5bNSTeBwgvw0v3yc/1Th+mTadlvjOISDPmXumCiSQNf1XHRqVRtywPWQ
51cYzCqfbFVRlBT6CjWzZ2UpouSbPdf70IGcN3ImRBBITNhoGK+70FOFhfWLKXGm
SVTSPvmHlz1zIDz9UjzxUPmH6oKsfAQvTiwzUzcl1CXoroG8GgG6Zx8Q0gxiC08E
frGJlBMUe4TPuNXAeMb7ojDR+YyxDsvs0La7RkQT/B+9pTt56m/wy+HB9l1aKgsf
Mmm7XJObPMHSrv7Qy0703g+rESM8HKBXL19kCZa06HjLsQ3wwzVObD5rSenJWPUH
i2tLU3QzEN2i+bdBhHrTbKJ2RkhUYCSJABLzZI5rHm2khfsJYlzuIG1/I3p6l7Xi
adSA9vRy5U5pU4CTY7b3mfIqhI1faoryywbyXxg+AhzMW1JreE3DspVGu5FvbgiN
c/+MdhymVrppcZvWIZDu6Lv7lKGO2g4PbPl/24mKYDBAtmZUc2YTQpUwzPAJ6Hiu
027UUfdza3NaExrW8X+P4I8U8wYmapovvCycvwvadn6PJmCjIU6f0T+JeT+bMIia
hQm8UDfbQnP0hQKLl1cytGYmRxN6duecklgGEgtueGBlyNLljz0odE/2A6VbjweI
2iqk0ZDemv6U/EvZJUyxU1HjgvhVqjnIZuZc+fSGcjoVSLTt6/rW+qp69UQ3cPPi
xdZfRjja/IXWG+dgsRvwWkTObbVv47hBaqL4Y7TrL4WFx7+XQ5rC7lp8JdeNvAGB
Y+xgMZwYrlue+ibvhDLYe5HjM/0n+/zfRk217WE1Akh10a8kjeqwHJupRbISNo+0
zlrc60WrsK/bfyn4ir6eDA5Um1eeXSCdRrqR78tCbcvzj3KdfXqtUM140ZS5msLL
oMh0ZsxXoj9v/Hv+khH/2p81J9V37ksqKaOPQlpO4wj4QoqIxwWTtNUws9V4YHIn
+1hWm5Ep6Ib0457i3966D+opERMdxWX2yPu3Kvd0tojuXUfUSEK6KVN6tPjGFW38
sfkXn64ArpYsANB0uh8e1Pqvqa2MZKtWUwKkjqG3HYJNEA3Be3loiHS/FJhrCjbc
WhO4jB+G5I7vyUFTYL6hePidSyq+ut+G1Wk45FAJ/JNodp51aTL7c2jMsFAiQ34i
AicpBYwlC0p9o71H5Kod3jI4O9yW7PWj+jwvZw/4+LVuGDrm4oI97ku6PkuFQ2+s
8qaaITIKTuKc1lKOIIsk5yIHyEjGoev+N7QTzD54RUD1m4y83RiO4nf0cxV/KFtD
VVnZjaPV8g049oBIVlyuBVQQN0s4U6Mj2bj27FzHrDh63kEj1RX5/Xc3QeZ1RPbA
baDDzUIgkcS93qXzsUoByn1QmmZK3/06gAle85MYBdvAz/OzzCek7OpE+1qYswtq
lmC6ji5hNgjbrajB7ksg1TIqpg4M20tUaVB0wKwBADAuxfFtiShhNf+HsAZ15x3N
wJWWfQnV0jyp/ngjnjpvh4cENXt/cLbyqZzTzqYOyj0SIAg3KOXys+k1gLAQNVab
4RLgRWzPhjpdmUzeuxkLMTv/BneLC4aeME1kWU4cKWdnW7R/hAIomMLxZneYN0MM
vSXACws24rcvau/jdd7CQqaIyCj+Pf8L+PcplM6Th1IosovzHyOG9Ap4KHr80ZH/
n8kxfF9UHsej7wrlVt+u3rxerYkNZSNpoWwktiQJeaNEvQaD1FsDeRWcpA+4Ed3L
r6asdGm6Db3B0G4sd68iL51q5Cf2SzPT3JDdLF/Ur6T/SEIxkhK9JOLJa0yiz5/p
b3SGymrsT3xMLopm18M6x8z4qKdIYGV2bt2UtBESLS3bkJDA+vW3yfKj3FjK11ad
Jr+AlsNe8m+UFB5B6VGteANiAtxBNxYeuIsgL7CQIcg44Diu5+/lPvcSvh4uOgKM
+3DomC5plAXpo0vHUMD/Nk+4ylqz+yof5McZtAwyQwTihZR7uIInxyCe/BdlnUHF
SpoF1uH7xP3pHtQqgr4RR4WPw0KkEtunZ0UgQo1lc4S6nQIQbcJpVBRBcj7bx6m2
v+Ppw33aWq2vJQe/NcWcQw76LwH37pgu7PjCQ3tFM8i2Lqwtx+1wSib/gv1A1jb1
n151E5Qe7ExOD1vdHy46vN+BvT+XrYnZbvT/iE5rCgA6uZ3O5AjW2W+pEjhqDBCc
caEVqipFohYYzadrHmhHVCaJWKsjSVdrxVnxbCwBzJVaOG/lsUcBU/TjEtM3CNxp
bCwZE+OPCOs4U0ze86GDaTrDVNOEQ0GnbuWP/ssk+5gtMEPnDPFSV+L3yk3MI7H1
vQ1K6lb0l+0Vy290s+0qmrUiBFqoCOIocfJ+5uLKi5gjTx6/fDC04k3jxo/01auK
bqYpxT436tQ7KNbqELM8w1KfsyDXhtUAInDSI279gemOfLGz1WNIy7+qiQpfHYpV
JJIB7dnW8SGvvCLVy8HtajOW+SSQRd38jrEbp7FFYx1/qgl9CqZBoHXel7fpk7j3
LAqX0eUaT7ojUg2GcUnQ1mr+2DRShFaLSHJZY7HPs80SH4P33gHmUeR25wTN9djH
Z7yAaB9/jhG3KW0IE0ZZGbyNwqoAAN5RgbQsyY3VNMO4CRCid7My5m6uZMPyXrYj
d6qC3oSklr7/u5AYYx79KzxX9fTdHI8Z008QxeKx2NtaToHVPb9JjroBjjtqVS9o
yIlfz3fa5ILSTb630GbJJCWjkIz96alX9UGsaEfl6rexPPId05dNb0cyBU49gBrO
TkLIueda3/EXcZcNxTiA+012te1ruq5EMOm4fzXi9lEU4ks1odg6cmv+0WSInanD
9mV7qgAlhoC3AY57zTHmRNo3NNooIOazzUgs036F/XFH+moKtk6LwqlM0SDKKqsE
X7ZhLt1HbKjiWmuRoG7+648l7zvzblPTCIPIULa3iajYqRY9XbCxqn5pqgyUyPut
k7iXLYIIL7jhQQe/R08OXsR54tI6ZsZlcXXUqj7OyGGqMOzTZ09bZOkDCiZVKkEp
x8WuBvBH//YqZkHddLYIC9PVAi9cu9FsTgv27qPSQ+JtfJGwgNP8gZ4WpZ7T3Cga
8wNUVVr9/tmFcTjsY5hetT8dgUq7oGhwxSZcauDARMK7CCtg6wtenQZ7ef25xj6i
5gcPBL9iz8RC95CZIzljAnWnWb+o1MJYNStOXESH6Gt8Ahjrb4rNwl9HE66T5D2Z
DwRvx/Noj6WVCpl9+g1VDxaodfSCUBlNO70qlvasnCBFWyegt80aSO+1P4fPDKEu
rVdW4nXWH++VpQ/l6JEekH68QivDLEUbwiXEiUdDMdrtTnnrmTvbgG6BauWXWLuh
CgdwSae9rDR8iBi5h1rJFs3VvvZa8bIrZ+19RWWC5aDJkUkdjUFr/RLVAlWI1lWd
Y+75EfhAZsiQmxghc8N0WgJzcArEOs3rSCm63jnFCEBebEffqAW44roKDoEtkF5/
VjT3c5tTOn2LSokuh+Ff6irr1YJpwuF4iu+EcBP6g/qMFa2SxhgCpiNAEGtUJZmj
FJSpQyDU1YCH+Gz/pSF7dBWdiDyzzFh3z4hkxDAzXk57zBAPbkxan4ih9daA11Fq
MS4CyEvqzik1+CUNCiDGk2FMHWv0u4tvVbtVt54nqABZaWD9W/GsYvXl+T0m7lgt
EDl5FNWoZuD4uS3YwGFMQZ5vUzDo9lL6YhaxKWki7f+lbsI7JXtKHefOl+81eeXR
fjBmBjmFGweEZJBHwzszlbAn5D+Ro3PNHz4rwUNBKj1x4eNza6YSsd/zifInTvzg
UaUIWiYxUd9J5t6m+YCPVRRjC8RHC1ULGWZMYRqdNwojjyuT2X5sKKgDUTzQKSIG
7n/ycMFKYYHk8T3c2bFa+y1czBGHxmCWktnnCJhSFzpPO9Hz5/zQEPAeUO5KQbOv
jNT2v1H/aH3E6ITF08J593gvx3m3NfE7oXG5CLX0g4Bl28dN77USCMrW2elmhGLh
XNyQXRCntgYPPBSwFn0lZruX4qtkOL0CfFFVAHosoL7I4gCUl1UmyectcPH9bXfL
eLURDYlID4Vtm+ES7tX271it4XkAUmdSADov9ypa0osUnEnOrFQzdEThzVxC6HF8
LWneDOANcsb+Hl7IkqEAeFWwUKr8gbZC0w1J74PSdTmhzVXaXfoqVoAqKlcW20W4
ya4utCWqrQFSSDuz4NnN9sw6atlltB8lIv2XFPvNw/2H/secfPvCB/WrclzM0gY0
FAL/K3Wh8IO62SG15+Cwg/FPg2XUxflBm9RskAafE54n6qodw1Kvdsf31uhSpaUE
Vrg8jhCVdrAo0HsqR2ovirTGD8j37EkTU/sPl+qXafT1xVFvk1WdS+qu+0jTxsPN
k6kKs+KUpxqVXsaLHffPCcKpjErNG436fdUW7zPRrC0vml3EvDNm7yO3I01eoHD5
sscsYVKYo7czHDwysynV4UC+01xm0p3xCSRWaKhP+WBSn3HqsdiVzAOtAkLW0mII
kqqiGYmnXvXP214FX4CDLT9g+Y2Kr1raAwaeAQHb5reaCfG+2ycs0m7CV6/hmkYO
RCs8QC7mZJv8X4gBbBggbPuyLslMkN3B9xYeq64gUxwBwspCSJLBgah+HOhdQLYz
4Nrwwz3SERydtfEzi9wVv2Alo/xaVMnrFDWuRmeJ1/QkvrOaqi6Y9o5suV41n/hp
G4XBUbFkqzC5YWeURrmrkOCm5uoYqG1sT3Aw6G+Cg10Q+DiCWgVjzZT8QbHkLC0M
dvWOEEby/yZsr+hrKPcB/34aUta60jKUcb8ukU39JVltS3h55ZOlYaWjUSBnRfZq
Om1IEnz7LeNRNbO1cZj0q4l+o+L7sqhr//DFBYy3+US2GBht3ylVQePInaHuqzeo
cotnJKk/L9IbcAhJALdXwVu34ONZZuj6cCLgbhxXnjtf3WV/B4VnM80kxFzaw4xR
lgL8QAFtx4CtAmcohesv16HetawMy2+oJ+I+1TGnIdUN3OQyH9NvC5i/EDh1N2Pg
Q2FnHDB2ANzmsps7vpCdrXlhK3bCfvfcx9NKvskpQYQIsEJa6+60ISp41YvfstwO
zrJx+hy0/VaJIG/URtMpidn6c8ass+VqUcudhTlCfU1YYG7LpbQHt7l6nycRxyr3
iplHfQHfYCtXd63vvGSlHVh4NaezQSoPFzyWxzFO5IsFCAu8ynSb5xXVgd27pg6K
PP4jRD2wrNvRilkPSjtjINDtO89x3AQwfO/ucRpEsAd5O5jp0Hd/XQ/4o95bL/kt
VwM9LKB3WNUbLWMmcoblQBc0btaj5W7+JoZ7pbVw3X4dkKm13LynhGBQtm80YszJ
5RBr3cjTTYBJ0VH9H4AKYBqcXh8EyYvtTCNYuFLM8/k3agDcNt5wE0w3aAibm6PA
yJWLMjegEED8typJB3c2TgbpijGg5trb9gEr3V/T6/JW5l53XMoyCVmelu6gkwij
Xa6fKnERyJUo6EeVT7vOkPC2aHN+1azVpAdLcrWDHi8BVs++QTW9W/vJBRDhfzML
BvuyQQaf4b7ppHI6T38EEm+ur99O9xVpjtAgKT+/LWpqSJRG+jq9HotjSn9+I5X7
lmwcQYaHhT4bSKNecw7zZDXMF9YJCa74d4Mwuw1kkHnFul35lmBgGMuyY7HZPq6/
EtguiNdN290BVsV+YwXSNHOBjdpfVO8JzyB86VIq4Mtj2MEtKDuiSfMUAnrmf4KI
vS6xTCiwyduVGlztUaE+XjpeqFQ1kzckJMct9HU4NqWt5STiZyEFs49qgeF7dO5f
Tq3QOT2zg2QoHqgy40siHeciT9eMKiaEYSfePgp72Fx0+KfLkR+vwwohZxOSOfCy
UEA5TMi8no1FkAu6lal16EXgQHom1eisNyFbytMoQHBs+Uc8byZ4l7aE6xZKxQEV
bgXtQFHwD8uKlyMt8lIcB7RskntQYpYNl96cfxklXNBms8oYiE7nulmNpjr3vXp8
qalaTCc/a0rPQ8NibJYKw3EEU+q80h58B0u2/flxc/x2SDBS21sS+50lcAd2ZkDr
fYfpEVJRDgZlQtdk4QJdcPhjC9GEVqKYI9zPjs0ywV0lzaAcsIS9ebE0/Oryc8lq
9EJVrslaycvYWAUY8W3rX4C/UL1Tz94MqCintRCgG7tTFpDNpCCJOWywQph59PZI
8sKu/Mdu2KpmPlD0hE2riJls1UVEiHpbkHegdbm6Ry2MM+72P/g0gKg71ueAsrnh
n3whigM4QTx1xVO/7fmyvk1SRvz5IITgRHY4MQROTA7/kAbDTp4ozOP0B3Ei6qOm
413Yak9t7hL+IXzd2PUgJVfxL/Bxb7/d5tSvWW/NLqhjljbO7pGPf/E9+bRHLNKM
TrP+I0xBJP11S4ns0v8mx5/ebxM+8nmexsH5+RFivyVXrisKceap21XheV0ok6ga
yscXhmSVdXdyylgK+RW/0oWHuQvDlQxYpkKbWQm/5kjr3SYHmNCuCrRMfOx4rHeR
9+yMvOhjq/4aUd9bmcOKGOKEMA9zBql/Dms2d09XAiQWC6st1UCUY/kbwuiydnpt
WdEx1kKSMBJ/NlTgwUwksliWGRduAbvFz6hJHDHBV6078OZBs13jbahs22HWM2is
Kw0OUlgkjqaION3zIm/JxalaOtsI6u2x4bYsP1OQ4RWgVeaHAKqNb+dje0pvSArD
VleZG9NPNC/oo2VQXlyd7m1rnsFtFKi8inj5uOWxhKr5PIHAW8wd/UoxrxKPse9P
nEA3Rg4aDEJoKpEY1rno/okKI1voq27IGYNDIX5MS3CPvneQBE2oKx12VGQxbr38
JpEWav08eKcbc3ADUzbM+NDY37FczclKsTgEHL0HVuiHdJPmzYuZwiixso7fwH60
GAReRNd53s+pAUTXOBCyqboIjPt0CR4rUomOQEOSjbmz7EmKXbirnjHzm4y4Kwxb
AjMkqKg0uUakadppJ/MiuoCst3ZPnAffCdWDgybU/rcUwMeZg8Pb4RrNZw3ALkdp
2UNB0ZIIxsosH26pF8uPp+JhxdZ+5NCg5rvLuo+Z1J1kyvWBDTXpaaWwyv3+28uH
bdfYWsyGRaUB0OGRmDnXEI2b3czFqLN2iglgwud4ve4tCX0mjd55HzAxWUJjaaBc
oFrAxhfA2SWogeFk7eqxPuyAb+gtZf4wqtEsVonNLh0Thzdu7OUGt4/MgyMsm+1E
ZWB5O5AAgot+Y2yVLSa9onPIg8Ittfz0yWLu4figkut4Y8GkULSLFOcjnp8wxane
ubIkTq9ZfBhovhrZulnoC1BP/ZnTqFgyTW65bziHLxcBbo/rbW/GE1xNleZYVjqL
hzJW8cYHfS9ciT+gdeqxAnJIoRGIeOqXoCOIAEKblX1Qs03oK8Jc7wD4Hcxs2Axs
HP7rn8y7YEKbw/B7DFWrecAFzK+gExD/d8bZP/k2UjzCgo+LrbvY7d6PYTNpNeK/
a9lfig0gZWJvghRv6w+IFUT4AWhcX3lyCAQsVOqg1We/5xOjp4PI2oM1Z9eMMdbt
wcRKltehqySugnBZwFX6V0IdddY3a0C4sYwGXmKJuZL98QnbVnV5+DCC6gh/OWGi
XhI3C4L0eGuqO+dJsExvZoKZyVSl/aS2YmD2y/ZiYbMupGeNT2f93bxesH77dX9V
sD92XJaEwWNRtlC4L/ecEBLY3WoVrrzQQoFES/2dtB1DZLMEGlC9+DRv8PhZ5XEF
/OO62VhdyiNKt1psEBX58THqIMUCbqvNfLqGeG/DxTui4q3w+DHKhb8ZF+lFN67d
FLxkeSBtcWOuTzwcirKrvBLyRzOkXKHaoNL69CagAGOzYfe4fEBwb03g+NSv7kc4
MniRki5vwc4i7Jk3D3792UQnx1KqAfw8upWvRD5F2KtBukXMhwAok0tWx/eCkZIv
pwm41QV+FDbJwuV0b+96TFTnZhGs0SzjTg6xBuXl8MYwSxl81xhF7e5ZVSWou0Sy
SuRqZ2BaGwomyYIbhA+hwLC5PUdrCQSqJOLtAK6oHHwv1bDArvSlmt74ZF6m3nzu
iNS2cZYns3uM1nfxhnYi71HY5Ab9V5nQKs2JG0opP81EOiHQPME9xKoEEl5G1ZNV
qQRZZKKlzr9yQHO8iiaeIS5pJEMkq6y/amHSCmSB8ASiNwUNvoagLA4PzSCdkoQa
cyaOoSV4oilTM977MzS0q7dEuTbLiTy1mD/DX0fdPXNXVDVYy4SOdpk9eL2pJHu8
bSqpbpx5U1JCVUt9f0UTweL2M0KmwkUN31nTyWZPmj8FvxXlk31eG7uaYyuCJzyP
HlatEKh5AxZjYT15JZEpd5zk6qg6ECgqj1ulStzwKm1WXuDZhrESTcmlI7tTSoX5
/WizNKtYGfTfH/SAzfFrqk91HR+NR307p2CD5tpC9H6vnYnOX/HO3XUyoMCWP7GL
D9X5N+ZfJrHMTEc9QJSNRnZitNYknIaN/65SO2oDxyreUoVBlwBhsWkRRAhUbTT/
D5xFIJvegSIfZw6fmJxmLBzbQInsKDehTe6eVcsaDJMHLb2oLWxecBTe4IzEmOu7
5hqYzoref/n8jxQZY+BJp9IBFA2lLxzypESb8s++4Vcjo9y31XcaJopQEoYr2MtL
OGc/FmzhG5kZpN+29Gfaf14XapaIEDj3VJ5iDHatcxFhzuzHS7pgylbET9T63DHk
FDRPpe1g2JIL5NQsgxgxzZv5oT8o3+UhcjkkVQ3U2QEt0YWcA1yGLktdTp83upa9
jyttNZ79uIH26hEWLxGDgTV9pf4+mA/e/fECCGgaEbJIzd+q3vbKaQ0wZVkNZ0+8
1b1I9ebx93Yg7zXEHZFj/hFhH/AUT2h8Hcqp13MaGfhSDlDLHp6lPj5G/tVJGXB/
jDbuv9sVRd3a1xZzuB2OvPjkXjVR2oMFPLcktwlWuiQkU8FMcm1PGCIL9sStp5C5
tfsFabwD1Jos8kqrJ8nH2f4osSEe2ILJM1OrTUN832TOER/dFBS+bf5J+Fdlyurq
iHsyRIQGx/uspvoq8nOpd+sVAgBc1dHm+f8CEI16Y6xVeC1uPobvImndV3NlnwZd
h0RZ+D0zIkBhu5VinFOl6h43VRD/ZVVKoetqvyUu5uCmFMZ4z6smRWVy31L2PPeC
ZmkQkL6vjva1rj8kpKVcKFr01sVLschEWdtLqefAeF7By2SfI7mHN5pz+nGMFG+t
qVbWwDr8QewgihUjq4rtL00Vzp1Ja/M+GPc9/1PlNyJFcm1hY0j/tWKELCTg77iO
eLmwi/1Z8zpdXVUsmAYwNoDdYYkmIarFlThkA1Cqxuv8gKGLWq03TW71b5z7/MwN
/hN6icq6FV1Dg0vpYKcvIaJjvAxoOl3OHuSkEQLWpOhWFvWw7wCFXmhO6s3Zx1Ns
qt9U2pCzCiZkqtH1gDrqvuvsM53dFj00e5+KhpMjYhRTDRsF3Tvfrye18aFhZ2c7
iNtM5Lh71xvjOXMtYrWD2tMBJx3uvZ1fBbxJfADpGtO0qdWlSY5LMyVKY8KMRidG
Vj8BvEu0BooJ6ZNGrHXIYJ2HsnvpR3a9ONWaiKdwPXDANG1eejNcwk9JyH/i1C+k
V/xnRXbsqICQCHe+apinIkAyF7RanHf5ME9JoBPp8wAikf2KDR9T7+TukkoHlb8G
zoDKXVtRncg72jF7IoSgWfvXKsoXtTw5dY3n5lxbS1e3rj991IJX+7p8ymmT5UcB
hOlt9ORHR4Axc7BTGMAnqjpa7zRodYdM/Ms9fzutyHH6F9giAekUPS389Hm3OPCl
9yBKWfDD8bmhYr38ELTipCzKPJsrTbR1o7hJChuHaOhff4RFXwzCEV/okWvRjXaM
K92O73Lztj8R/bjW3PlwQCu4bS2xL/RteQoN+ExodNSQA3SpAMk+FA2tvZzslyGN
MYDH/OByu47hAWCuLjAMsA28QHCS3TO8QXnj5pv/WGhcr0hK9S2K9g2i6ZRocpeo
78uaFoq5L3q+ku2Mo96m3mxuR2j0RrfigEEOGBx/c4t373SNM+mdiOdFogxrEX7W
zNVBAJpcHJau+NPZjdWfRaZoVXDaQSMW8hSh0CJShypJa2CBjfVCDn7QX4pnGc/Q
al43YoTf+PSSOJeTb3QFSAclW58SsLDVgm5LGgeIxOJzo3lG831UZ0ny7wwqGED2
Dlchkz6Y+GspNYafp8ZwuSdnv0g92cEScLz9brWYQP73zRb2JZ61lfGXLe/tVmiM
Ha5cLWDW6OPIDUbtCCQiY1uCEyxSDD42OcvAdXv1RoCHJpfG5l1SIeHItt9nfORD
+kyNER1O5264Z91tkEiY8prWuGRJGzyGpC0wv0Mg+RUWCl0qTtc2ohUz5X/yeGsR
LEeyGNBpmy+gWbP7LnQDqv74PcdYRduvSFjG6cXQaWQ4dfwpCQJ1jPkDIPi4Z79y
YKjaSSgozySl/CB8+pStJJDI58l0ffoGj4Wzx/zNouu1IKvL7TI99/H+D/mleL9G
9K7caV3Kcz1vLNZia9oHr4cX1uroFea5AEq8sdAGWkuo90FAyiTiCBdIsX087dpO
iVrYPDpXN4Xdbz9ISF0DsOPl08bMblcPXH+lzW3wasyRw0PAIN3KeT8ZdvVo/PW1
FFbuJnUFpsteYUOBAIp/Vg5omFpbfGSM68U2TuiJWO/VRWikD8uB/HnngDiDLywx
1mApPVH8lZpLJrLj4kA8SP1XR7mJ9bf1nohZxMgGEqXA/Pi3qrO90MQgj19B6jHn
4Sy8QD+q455Kib4BKwhoZhedYZRwrswMOeuGuknWSkhzb1SoKhDAiMdpZ63PEuLB
cTt+7jg1kHW8GOUf8lxemx0IFqeUhv/LOEfafdLUFHy8GnWZcD/rM54MDrJG5/Q9
Xzujv0RrQ/gT7NnnXWXIdhqZEmD+l/rFrR27XcTVl5US1Lu56tOTaItW0SeYLI0J
RxBtIKwQaywJI8YwnsNssUIjXWzu2OFQ58tP/JUzk2t/iueEofmnLiUFH96S09Jg
W5boc/8Z8X3s4avlTAtJ/jcVvU7YcZYR6lryxil7Piv45np3HvnQYrLtSG7/prW1
rywbJAQYfB9JA22pv65FGOKE+dG9ze4Ou5v+AV+3oEP/HWhePypiLC9FbdJrVKme
GvJeXt+0MIFCcWPogGz+PfT/IOfuCXgnyIFs9C/QJmOdjofZVOMnlB9kZY82fGYc
KGAajkZVFdlEOflspsIa+0vKzzX7gfA60mVFEC9yNXphgHdCieX8kYd2brHQ7uwF
c25I7mIGZb3qXRxe3zRmYBZXuYs4Xe5tj9gumC+hSEohmb2ErWQPIszcMKiLo9q7
0A4+SlWYQzXl0mT+B6t99lRTrQa6KmZOL7+g6ReCuK7k5wQtZIMwM6mN2Y48Ax+Q
iOzZQLD7iTwsgIuo6tgp2/kTjOyX/aq43oPevm/ERv13E9p8nlmqFqevt5JWX6me
hdxERDu/7i4OcbsqNw5z63Ky6wN7vrOdXwLdnBfOGI2codoiNMajw5aMmxqkYEv+
/0PXATJ/+vMXLBrk69sYTLDXd5GNHE1uc2mwDYkfg9ABIAtLxkapRtehxIC5q+ZU
UMd+4THowJZBePehFNPKfkMl0Mc0ZThfCvOuVK1NkJe8oi8dk95TLpZK9KvabDQA
YDENx2zsJjr2qPeHTeowyEc5lIDtg24JA/3SoXOUEoult3wbxc5d5J4U3u2Fu3hO
4kZwBVk+VO4WwDw9roA799ihFQf+eGiznE2et6X6uF7cb3NvaHjIVHazkGG/U5b7
kboTahI8vYUOzrSE8LAtCaCLWSbbyooV4A4g04oz96LD1DbOedCtf9UrdSK+ZgEo
ojoesdRLVY/NBO8zfRf9xS2+pPAs1wBMWCdifilLYN+gNdoMM+SqTYorva+qPnml
H5VoJFHuZORYhZYJG+6i9BG9CxLZUh/uCQ0FS/1PC1xZkhaNwRkazhQGWSfJQ46N
4NM50ZLwYHRNz2JhS9ZNUlfJ0FEJWGyHDm5VZjMdh1FA2lauSbUS5Z4jSSdkEK2N
6Ffj6FK08VHkdBxsu3v3sfyGKYGCUVceqSWAHBonc5ieDrGQh7hrHDF/90Vk1zuQ
xlxwX16Tu1OIg23NST3oImzgw2vOuocTHFkjjlgUxXZLBmQXBgbospbwLDYHLAzN
82whZj4JhYDrJ39ispgU8I6jF0+3c/Qqi6auM1ZeJX6Es95BLqhzquehTbXmtsx/
n7EGy7118nQYvNcP8BdkZIU4GtmTHCX/s+QuFWM5jFBAeGMDjfwQ17xq/Z9q0R03
/+uzyMbjEvFVw3/I4lAJgI/Dx/sX5Ht8IILtAHtEUGQyfTPVdB6GljoZsCXXDqyY
wU9kCAveFvghaLl3ITDdkLmxi2AdrWra+Uf34hArPcAbg2s2NoC0LlKXYcE5dO77
3KnHLFH2TyzY+my+C/G62Kt9qw4H2o38BE538VtH85BesxDdlKJjtGvrI6hnYMzd
r3uzwMhBDO6K/MBQ1/O9Oe1669I0YSUACmBRUL3heFGxROzfFIuDDQ4VtiD+y3tx
ki7pyEnBkQuiTax2I/FXYWLzSaNYgN6OEk1LL/j4tuqVHOdFgsg0Y8AKl6d5Fe74
JpFQSI45iQUhtI4420S3RTy1Zg6AP0v+gtLPar36gqKDoras7CcgE08+NThiSH3G
8LV1B8Vjtq403OnYpQhZvXQNHXudTBp1MBRgsaaCx1MrwqvC69cdGScC9QMuqMcv
1h1dV0Qyd/WYkhBlQ7gfkkafxyTEHdteIWjrQsybbrO1Y9tmY+T3OSEsyNNzg/SA
I067p5M1QRxXlKIAqDt9eKukCMOqHoWTbnLmamuen1Wgo4RNZnQmzCVAO3W8B/XF
Y8DvWeYbFbrbeR4gteIJTH8Q57WeJHQ5epRjzlm89LZkrutH7AyMC738R2+/DUlI
rMMTCQpocfkAnEFm3Bj4UpWSsqO3uHzfR+YemnI9VLC+NO50ZDrSTecNefddnclt
oSnSrenFCA7zxUx5lxJeLURT2Z74NlnE+P6s49P+L61kPjXptRswePoCaNdEV0EE
g9MFg7TY9NN2SBeF1BSnnGRcOj6YVpQ01HT6Td1Wjs5Lz1vBZ47pzsbqcR1eTtJR
LZawPEJ3kIya3VLTKRXELQ5+AomS34BWKqwUuMboOoW4a5ZsIRA3E4QUBdwvRFO5
6yp4Mn4HWuzt3I4oIoCKQNr55V197diXb0Ot+ECTQWHLjmsQmYv+h7oSLmGJn74N
4oEBB7rxewY+UH3PskqnLhg3VOj4PE4+Lx1iVk3fIpMtfUHVwta+f5s1fURXAnYh
0P7zXBZtmbnGJ3iEmYJ1JDTRHF/HAzVoja6RlP0Wp9VgCOGEUjBa84TyhUaglvZA
hFrp4eAiu3uGxEYnyso9XzcFQqHNgtONCiazjZP2n2SxVoKmYJGkLxI9Te4C3VeD
A3O+Lvjm0cD/dbgJypQkyh7mniPJ/AcSygOFo1gawtao8z3QKVLSXdYcTBGgc2eN
0felYWTH1iYi0M2hOiJbyoNC0BfxnJlI7b8GchoxS7AzNcG4wY/kew50Jh2CN8s9
HogLDYv37q960y46MfE7ucudq9eNox+OVyCfYZs2MnwVg96op/4BnPGtn+nk+ryp
qDJe2nujgxHjpv23teQuERPtVsMJTn+8ZWVSzzGXtq4kw6TUVVrBS8uX7SSU8LPB
NVtJAvPVFeIyfI3J3xlve4ZPbt8efwj/BN4rNZhSgPJpmmDzrzT2hgHCbYNzh4os
/EPmInGL3EUo1aETu1sJHagcory5d3js+DRudox78iygQmJG6EcakhgfypygERxj
gItCmEA25b5V8aLTNLaM1+dwDNWW92++czHuuSuhcHHvtfgnqCY7zVcHJ0f7xn9B
5SNCPkiAtBs9dPZONmwT2uFAQOW9Yaae4aY94rwFukCF9TQJoT4g364BnJjCRhTI
7vrQWB0Qd8gY6NP+/qaL3XiluV0eYCFG1VqQLV5llrCAFIk1wWxmSIaD9BENPJmM
vcBZGWsOKXmJ1wlq8Mo5bcSFrRc+qf2/8a5JIb+hQvLnvi7Zfa4FnyraEiGjYej3
a8iChXphsLLSsjhgMCZJ4CJvHUXyMQ2EhL6AQdn1gDODSRiewA8i37nH4gMuhhnN
3q/8w/bBHA55JS3nOkDX12EqD5MRvU4Igecdzhl0rSjdY2FSm+mWX2bN4MIfcEeu
oeseUV8YgcXnxDTjWWlLA6vBHLI1Mkk2ieO1ytNAxsiqRjV1ZJ34Uh0qtF9EST4D
kLXfTu/o4Q/rWzvX4jXLZU7ltMVoH5WyVcStK3GteY7bd2XzKUua+29a4q0n51Ok
4HnM455HDmzobWw1bpCVN1QjW4LcccbkqEkXdrMvcmkxfDlaO86KNld+XoSvPPgz
7eCM3mSSEEwbJ6JRQkPc2TgM0cTVaySQe0sMcWv7nzamhdJkkUN85JjhHnadH2Oe
iSNmDFE8f5oO9J5Z+AO1oKDN5ZpPI7GWcHVpGQaEN/lMMZnW7b1erVwEtildSD+C
1AYUPRE6nU6RrZGPxdavJN3snzcmiMy/LSTJRCzz4OmvtpoNycVb1vp9ohRNFWIF
w0pPszRYvi6FnR/2TseS9dgmFmBmgQv5EGtlTWrWx/OX3Hk/XPdLMfN6KctAeWf/
ZAlBHImXv2Ebq98A4Fg7UiMakNUmQLGBQzESKGKaCy8QDipnXPk5tUBdCwjUP0kB
CFgarhuJ2sPA3BnSB+d8NJMaxIl0WybJEkS6oj2LZv+zPzpRSdfIGPzi7RSnXzD6
k7CYnfuIX/Wq5exe1CJAk9f2Pcbi9W7AjLrtM5vugviyJKNWHpWqwnhZASI4Uac1
TTk51xOiUJGX1mPONPBRQ1RNOr3iqdOU0wPgitkc3rLXsfisypQssTtk8dFedmOs
nAFS7CXJAgHhOB5R751S+DAwxM0EpfWrp3R8eJA1sH+WBD/iVCsLym5cSSnXr2Od
BK5R5YZYC7p69qNGqZ55c2stP4tYf3uNklABXGz80cDqOEmiJLZBoOoVAaEa5RKk
Jv5xfQGqTJzGQ1Tk0pqd6dTDl58JEVao/eOw0hFLWO55XWE62ZdU2GGx/K4AGHqH
19Y5X9h7dVg8NZ5s6YcwrkdvCvJFlc36DR7foebwklOuWyofqplrQ6uimd/eeTGX
ld77ewkH3O783NuGsScAltNTNZqZwsWjHSOtkr9cKUhGFic8JACdRIhnAAkKqlpo
LLoRrAQ/1t6UTQrweaViRmU9LHRyLmKwdHX7Xao9NdEF2++jmkYClMJj+6NUwGAP
4j39d/Sx2OGeozMzMo1RBI6YhtjiBXwfklbgGgt4qebi9MHedzk0g1K7t8j1jtn1
0qoCcThNSQWjdgMzT7x+y4+Vo8npDEfA4OKopRzzBK1smGb9PaUGKjkR82urm6N4
yXsidkwJV9KzJJOaTtLQ/tJDhKIDGY1vZVKKpXkd0wJmR2z1mvYy7vxS2Wx97r+9
hYzlDlx6XWFGztyFHev8F374IGseXfaVGCvemNi/FYTgsDyX4boUHtClu6DX00aB
Zd7Wv7Md0pF93ijflzz+e/238p7ZI7gr1bmUzP03yw6RugLF/VT6Os13zBzI5dpV
vZI3EkQfsbj6P1Qs2z7oXRU24UdGMLNpfWoeZ5WNZDmZg4GH2fCs2ycvpc8ZPwnN
aLP9vayYXflKP3FShxyv2H5cMok9LEXj3pHv8yUX5sG1J0mrguT4IGl4r5awb/Il
7ZnYwRdoYRqF95WXdGo4tEDuvapQVvzUw+EtfiCS44ivmig8kItnuXZmBKzZQDxq
i8gjICNSKBlbF4PefcE50IvpBChfjG6gnk+4hjAU58TwGjCRDM1IUcGwkdClhfN7
vKqMLU/tBgSnhCF2lsl1a1Q/LbN6Xh9JuQFBdbMwI8hrc/GKtUJIoLBBjf+Ww8kF
JMYqAp3ljvoluC3tI25hKyv/JoMjO3jVu2V8mh7JKJWXcTylDRkPWPkKh3/wQWX8
6MHC/4B0D73fm9mQJbAo+NYShCUNFP10dB5naH10PRDHrSDAEOKdZHAqpUguHvSu
nuMSKXrpxMWSm7T/WAoe3DGAtlwT/TOBqO2K87MKUQ0+2RHunPIqlyEkBqBqH4KK
8wNisUC16a9ID5Vqy1RSkQcSb/AIKhDNiGb48H1VcXmWyDT83BWPMqtIABFw98EB
H29g04HIGb2B48+JJRpsHittl7uuaXdzt2nBiLiFXmBes6OJt/fzhuQJ9CUqXVgG
Od+KarG5AnY9/c5VM48/Yy6aTvvt9DRL0V8OOTJYiLWfU2lcmPS/cKwJKjkg3zAp
Q0YSleV2w7TcJoEEEiMOnFVkpDXNOwNmhO9IZJRoqAf7/TnnkJTRYMmcXKhBe6VQ
4kHOzbUjv9n9Nqfh4SyC5X/hcDTsBlobF0gFIO3tA7aCYHTu3A8IxtopbduYmJAi
NV2l3Af9GA+zhPN7HzH0QorRowZK9vlCxOuQr/GKkus5tRvA2MRiRt2AY30zVcR3
DVURmzWmhE2jq3mR0DmjgP6J51yOWMxzIMi4hOoRZdsg5Mx1pc7ns0H4Ma6FO/wZ
OEuVGG5AUn3FSm5M1Tyofkki8EbC8O4cJPaVl9MMOIAUBhVn1uf7w6S+GBxf0iPA
IMqj04F9mH2x+6D/vxfeVpNmhaBfiYsUzJ7nnwFJtu6Tda6PxFMy6qxcl9WO5Yp1
NoJOBDxfRr5koTiYG3TfDmm9G8vyaprhvCl7JXrY4qwlp6TySYpjKdUC93vaBHz7
GqWy2qgV8J/CIcn2z+Z4Q8bin3XSnJ6eq6c/Q/PrMU1nxKuKmSJJ0B7leyzWXzGu
Vdc87gNPPzaDO7x/EmP9d9h+vK0wGxbFlurIbOvvevoahGpJ5jNrGFrZP8KabB9R
O91qBJhyBBPxXDkjDmm3F0EOt7dN5+V7Bgp7Zbq2S+rh4fJe79gpVN7CWt7qJhqj
nNrQq+VdHo8Nn6bdyuoLCNvoWCMBApUbWhHNIBbgZh40OCm+NpSlacDh3VYmrhIE
JUhppqp5obiH6Fozn4ZR39L40dN/19fwzQJSLbmZg9m0gdmEmKzy1ahER9Y49JsS
I0VX2qjVf0seANZfb1V7Ju4fsf9CQL6KzBWXb1ghSOTF/P0DyBF///0ejckyMxEi
HlmHGjaW6qU8o6CNQm2Dc29YZ62tgcnmkdQOPvrfvjtJQNTGrkKiQET3Mt1pVR94
sMtUmKe6A0AH5Z4UyHo83A9eBg+ygVkSwcqFysLMDG3yTjGbShAVX5PXGWhvQ/ef
pfQHVVFqwQs5wd1Mv+glm+mDhM0jlQKZiFUMyij4ypydfbm2Q0KZZc9inoww8aYe
5dwZ6sXk5iArbOE58lOVDIcaZhfsljjnpUP2OvlQRBTMbO4iot0qmj/pFOZiVo3G
glUhBk7XztkIv959jkvObLkR/4mpTWIbSyIgBY6P7O4G1i8whoJh40MZpChaRiN6
G1d1BU2XPXaAfQ1qv0yJDiAGECLUJ70NOz6y6JxsBoTbsBHW3v+u86dLnxDKnw8Q
5oVst8i5AvtoBtLSt7ZzHLCo1hqwLzdNOFbRRKtgzMAhmqx34FviD3VFvTQ4lf1j
NH8fCfilIJjgbyUjf4jiNVXyXv8IlMvG6utv3VbtkKd290mNIGrpPkiBQGC30rjU
Tmw+6Tc4PbFW+6+ySe6bT2llbyN1Uy0pde/i2GNi7MqB8WkKu6WPncNEa7ZS/Lrk
maSMDxTeIjOpmz4aqf3lKlLqrLR66ekVdQJ0CVnYN2AaRJm8kb+SN8dkfZXYPhAg
NARzPaP5SNlw6edYSbIspxTglXzqdSknRUwW1iYss7b8ANHNOEd2XxVKA3wN5m+S
8sRoYMxLUpXaR3OPnYosgfPR8yi2w5AAzyMruAds+LFapVZEPcXIue3UEyNxYK8H
lx57pp80tSYe+aNc86xiGYISzUziiVEslOuCDAlPGRDe4vXLnp1U3ArPKOTaFvU5
6wPISlBn9DgJqsZIMHvoO2B7Ikuqbt0Z7pGFm4d6AuwnWNF+PWQ7fxwByIUGgv1h
KT0HBYpITBwBV5fQ1Vbe/z1CXdGgOLtFAXvOMNjsCVE1QZJcEqh64Y/i1PlztExi
Mug/Pq1S9nzv55GU9s0+yFhGmqDRfE5TQQQFXbl91SUOAJalMrIvrwh1+aqaY4b5
U8XSOf8V4EjYty2JH9eJusXqFrGEdjkdy79mdwMkFQ2Rb3ViZtftQDljai1epndf
BySxvq8MQ0Fq3AIRxp7QBvwC5Trux9DjBc2GXqpqVM33Pp9fV+4+wdYJPu3jvtgu
JqFHDLplz8fjS8B6lRyPsZOamEQcgzUgiuDO4+cRNsg73drQWIx4wS61U0nP1x+s
CzW1NWGbWnXA9d/Xc9rE0wtBheRDKhQLCaq0V9B0jrInDqCvRUOYAR9Mt1ukT+sO
OdwpisfxzICHNm1AlQA49/evm7WtfSO85fssQ2k8DbjqLnnOze40cCHrdzi9b097
cj0g3dMdJZE0wx8T/i8BmvWqvOF3AhumXbDjiSzYpdMTb025anw++0hTHVTzJLzU
L0GUIaAj/Yk9H0zXN1DW6sISf3josRcrtgmbi4bPUxL2Un6N4iKOMyT9FrwnUkSX
oevc56yJjbNhT1chMkdwLxG+vf98kCM4qNCTjyaeg/D8CcfKYiKy+JdHbcHdHV/E
kezODdPh0sZfTSK2cPJnqJ+XIyUQGTIiu51Q9dks3dYmO14T0U7p4ie/I4NWlgNG
Qw/vxZFT8kaytAz+Sd1lpS0EmMeRCvNc3C1mMoog7eg7gA3F/W2Lx6gDta5lC3E4
nXWHuexYk3CUbSI7WkA9gfM55F1rO2+c73EjVbziUAcVWG/57ymBvha5OBe9AwKI
w+QsnHZ5/5FJtfCUZWER9ulCfb5ly5H5vpk0dfSrbOeNlRezgWK73Uu8mreCoRHL
WvX9NRW9DCNbFfXe3EzDYA3xRy27P10uLGnsulRiCNKHjqwmTVw7wFUHWBEe+RXy
ybwI1QsbSqD4cFkGhJpoYdT9/W/CVPDF6yXr0N97Zggk+FwyPr/5CN1wq3QHWfS5
9moVCINY7NAR6M92l4xTKz+OmZ6h74sOH44yl1tRcs/mSit8pFz/eVJvM6ZLperb
l3PDXrpQW+SAd3VWOg1eiK5szCCD/kQLHKExVJytRIUcwwniTR8xS/nZE/L3k8du
3cS15p5bjRpImNW5VvKby8+P1+5zj+uTNESzXod8ITFhPuLJcTRvjYiJZwGLZ8mP
uWMAcONj1DujkYmKwaqegP3Uhzv3bUkxkhyjM9AkWbOVOpiBAvZep2Jzw8nh7q6+
PIEann5ZZrPtMX9ldIJAzD8YcQCUFL9MqAXxiDYG53Evbp3rP9xDC+3zopGmhK7v
blyaAxFxG1NgsJhfMULkwoxSrpyeE6ik+hhynsOvbt+G7hKOPOS5hLtJwwdjdLk6
3SaBkNihY2gqaCQXmrjMhfQW1GEtHEwBeC+MYgy7mBy2m1469FAfSBG2Ee7BeDXx
ppoIU+Hm20esQe0vQ8ydlvnh1gAhKQn84T7YEAiW7qbLHijleDImVMgOwVEw2G69
0MPqMbo1TWFB+sg8uP82YpXLcRA45EJxZTSjRzzlrzjPPz/dgE6ItXTECv95Zt+O
C+UrX2+p4Qa9WmC8rOQs9coYpbzee6bKU8iI6snrGMCul29dFBRP0fcY8UyRFgnK
msswRYBpHeEJG6A9ZldCDcVbNA8HVpcRwN/aN+RAqb/chSi7uhOXuMiSHL2K1OI/
CxTAZEh0RG+CNooaaHiawvLURg4P5xpxb6vaNoDr2FDtFtURm50PH6Hitq8M9Qey
mA6i7Gc7gddhAzmnQScLZRTroHMORDAptkNs1Lx4AnX7ExLo4LPa+ARwuq7bLQSp
QTCtdd418JIwKZ6oTJtnfM5EQE/9tpXlddYXh6lJqvUsEgPYQPR83qppt7JvlUKQ
GnrDmTcp+MNyCcfy7JPyAV7YQJGH/LkGfWR6YfM9CK1ruSJ1JxH0e8f2ObopYD/7
FdhIC+3qFyjhjOiBZHujS8W5ruLPNZnD/qgCRzaNa12LvR7TRAasMfXvHHc1NTyW
9x2iyeDqb72YEBCRARxrs48Bglg4OShJVtHPqK5O6Y93Tq70JsXYnr55+3uySu6V
y6aiirrjXqW6Qat6VSJwbctSgVPygOYzb44/pIfQg7N19n9bjAeiaKZ/PsBrDAEX
bXn0q0/Amnqqz2+vgWRRlD/ySaAkAzH3CjAvwmVQz04sqG5kd90nMWOGgL1FX3uv
UPVgq9vldi6PBI9bz06m5r6ujFQZ+WN+TWDTKHU18VJ1jduNRduv7eUP9tcY6kyF
4n0TYbM3IbZmPazfnaSFb2yW/ouhwpDI1nakSpSg8XEZ7zJcBTrGWsZo1I9LNGKV
7M79ZlCj/xQnbqZyb95Jv5aOqSGzc6Bl6cxOMYdFu4D6hE1hF2yHnOoCnrRs7m+Y
uoCu2Xm4YE5VEiO8Kkwel/2HoR1wQJpbgkQK4eAXRGfJ/YRI5EHeV9s6MK6zpljX
8Lx4tbEel/CwmsO+lCaemmuU3VwniL5HqZRpch5n2FmooqjwxL/OD0CmFxqO9hLi
Fn0hLbo6pjCU3dPvgHM8TV90md2V9zHpWTDx2Wm6Q6mGH2VSUjtzZI8fGOAnV3Xa
wv3HtFAYfsDBiquYoE8YxL8cgRbr9SbcPzKvrFc1Y/TXvKkuB0sgeguhby9pXrhT
TU56e5yLOqwVaDUi87PCK11XBODxWNOoQTq4MfSsLMtWKNCJT3gZUWSYgDBZVSGt
Sw+4v5QWb0llXZYQGIE5xMLYuUWa3wUNEWRVN1Zy+icxtX/SDdAk1GlUgeFGct23
043nKGTXcDqsOjyf9liZfKVyflkjwNSEwvIdYkzEf4omcVLrfcqsPn0EB7buFjY+
1CDb+MMK9+/Xkl3ypKTcGiPCQ9Jslf0DnudGTanlRxiPOVYLQ3PA6FAX17UgX2eR
bQOSlBJv2x6pDZowh8T1TBOJJTIi+tnE2SmuiA50QB6n3XkiL0Z4EysJLztintTA
v4Hueri2yhW43T2X0oGGFp8hFcz7YzWsyRpbxDD/RWHIsZ2+LnJjUTFAX0bY59dD
WRUNNE5yJoJOIlaskTUDRR+qYpy0Cd20z3EFCdR33MQ8mfuZssdkmP4jk/S73blE
nv5kT7XoWceWNIe31biHm8iI5ZmF3lutkIUXItaEHlBdDS4oUFm8h78uexRPC5SF
yxv5C4oaBq2KReZsdaQG3qFNjqH1Dnx78+kfj65nmd/4x3i1dHP3HeOUi508Opyy
lR3oBM6BTuIjD9vLCl5oUlzvHWotgWFQrpGrb+I5pJ5NBBgQnc/29M9PsC/cJQoC
6ONcPPPCokNrK3olt9CFFaqMLUUPGJkbK4ONsRIfaAFXjyWMTnI3KTA5LXALb3T/
MlYv2opwiH4QAqTUE+4sIxHJ9T9hI1Q/L7bXuie0s0e+OOGPKs/K3RPr0bxpWQdX
hvmX8WcipvYn5KGLxr+R4LaiLbdYoxY//g98ZBeizX5M9/XwqlS5QTQ67rQJf8uW
droxwDB2n/U8L1FvNiiGb842Wfc2OthlVf/3moUHrh+mvX36Ay/duJxXO3RfCj9R
QoG7hK+U+AEuhJQnTVUP+SW5OSe0HrvwQkIF+PJpEl3U+VT/HOxusp+GZrlJ8Tbu
87iX2Y2lM3F/1M6FspTqH/BfnksENB0L36hCkM1Ty+SmglhZEyf2+++Tn+O9zzjR
ThiTT1KG2oqIPBjVSc9372j4rJZm2hIFXCKmiObNsRMkSSt3MehhcNAM6kx3/h9J
nOesTujsASQzvaohiHLNWebwsEbbk7MocFjlcxUxktej9ko06YKtm9L41lWv0/zS
A+gOJHO4KwwTlFpPp43ESIfNLj7+NHHwOZH96YUM9k6+SRCEjDr3SdJQoUa5XkEr
5H1fRH9JmbuUJDrATOXBzHSBI0Eah9wIjMVExFCtCtWlZlcm2ZD4NmN8KjCV81wO
5ZE9zpL+CzRF9VenPhXD8FypFCiXDPIbcnGXLSC4WjVokN0yLXqcLSfJRW9cST2O
Us7ubRMOObqKUCSQnWux4AtEJSrCizPNr+XeqO236csBBGa0rqWvVU3q+aFNaKka
JL6xr7t3f4BCBGlgNs7v9AEhk0RUJBxv/4WQMEkwpMhRu+sh05n8X7DrALUQ2BNn
9F2eRZxT8IRZGLNlSkPn/tK70YZxe8H5iiTpsBCg6EGDlqGeBRzn6DIGTLCX8mY1
QqMurG0y9TFmGG14GnTyKA+z5aa1RLgZgwXJpzEx6lcX957MMeVr82L0hbCafc28
UxrqTso9JZ/ET/lKKSzmooSidQbCPU7PP9dpb6VkzariU7+yhwSa5TE1zjoscSJT
qdYDaywAKYPSeIAKwV8/9KkHqUQ/oDHawIF8xfOO4ESZkmJpTVx/2FW0G4/nS3xA
R0Ccg1jW1KzSXZF0cfxoewxROzCAd24eSAXx/hx2O1+keIg4YcPPOz0rPLv8hEXW
sXDe3E4pHEhi/d44Xl8a24yA/LFe9WZD/ZceDjIsnahiTQOYomZo7qC50W4k5OxP
gqBHXgzB+SGPf/Z/PiSaY4tBTXT5O9AhwfgpgulKXUeM6X50yuRpJSWRXOFzVSZ3
tmDOQbtkIE6Kw2NcWoRIxiPK64Sw9AcnSVwY/UdtssSKT2P/vEitv3q8h7+RFg85
nsT9nMqr9O0DYZdaPJDcLyEH9CZrXBa7KKOkJ7/ZnUauEgIhA7zZjWbztSYUwnTg
a/w35+zq8fMOi8nqa0YUnUIz5K4zsWJY3FhBA1de4G2XsVYDXEtsTxlJSjcJhxCz
NphvGfDuckAKK/D9hVl6xMZb56EU18o2NrTzGEMAhwCq0L1oj2fV9xXloCrJLc7r
0cWNhkzamEW4q+eIRORQqEu4Jzi0USElryytWTNH6DqX4O1goLB6zpv2l8wsfqKo
MJp0LAWopFWjMMWTeEWLWs6QqH6TDORnx6KWmgYDCauTSxIXgpflO1t7/0PpVZ7D
bh3LtseJZ7WSdIlQs+KmVn9YO3zqYv2hO5LHr7B7xXkd4R18DjPfi4lI1WrL9O7z
3I5OzMHeK+J1gU8Bfy1S/PfKsSX0Lb93j4yuUapbqs61EddWxyyIeKBGMflpTboX
iimXNDsr8FJr5+hCCV2110oChRH6Bj6PPxlxpOx+0QLMN0y/tA4RQZXUtoAfqZ3C
DwZraZBT2xbrrFiKCAVh6n8TcuWGSoMblXXHemAGc6IhikROn+vNVSFQeTE6aMfj
wdf+jXPRy7JSgy4Vayd4idyk6YPH6Pxv/exmQauU2U4higbX/GfdkBACqSdj8cxO
1mNZ4v9E24fQ3jVupBnobXvZugbmuU6TcaPpoSklgr0nYQxu22Yaf1cQpYm7r0mM
UHZ8K0pybWKVdaxty4H4vf/RVYTVHOQX+kG2Ufg5bPf8C15sfrpUDt6sbULxypiR
i9UjYpjhxVq1Cfzq5gBaTT/BvCsbO4LRVqCtAVxhIJL5A8IhQWRx+FNH6KTTLli7
/Q2N9R/2jTc+CAPrO0chpMBPK0q9IgnCcinrzi3zol1P44igP2fgBo7iTdZEyo9W
5KImes3KZKCDgmvlSObat8VeLMFy7ze+SITXh9gG/YGPBKIe6x8XB5f6ENbx62ry
BQcnJg7Dv15VZKofC8Kr/WNu6q0OkiHHRHQqqlNMutpPW5n1d+XVv5VQBvaQZgpQ
AX2zmAU6qjq7BWbB86jXFk657/SG1vDtK6WorCJr+QxkgVCE/1I9DkBaAiZzcobU
GEhCd7TGc7lAVFg+tsNabor28/RZw7MJvvUAaeFidHFz2L7b1VPPGa4j2HXBwyqr
Juo/iiGRVDXvmWPD0qfFx0JRggsHnOwpQ7HfPy41ylhi8e+vH5T/8jWkBy0NAKCO
PBfzxTENthqRB9TUfoLVOcwZdN+BHMfrv9FVjZUstja58/w2XAHexxI6oPJOHAe4
VFXxbrLCx2dEd67vkxjdNGp2ZaC14rLmCBQaDOfYPnntFUULR/Nsw30d9IcpSNhn
TA/yM71AmQDQv3pg9pboS6QbGjyguPhqKbm2pTth97qhrfeCTUCUzKtS1ia3G9DO
4azdKB3+c/f87Y+PiCePwma5JkBQv6r2fkBN7Q5PJA2R3B5EdWWenI994xSWT07q
6RAayR9ZU9cthQ94VfwX2vMzN/rIJVJdmEnoN2JwN62qj/R+/Ttio9pL+/G3X7PD
CULtDFdZLpdIVjE58Y9QLENGc8joQIk4b/30AGy3I9lW5bmPfVyCDNF8EZVR/cnh
fgIK0BGbHpIcOf87kO9vJTb9WqsOi+mfhVObtUzdXxctvnlZFJPaY1mfPqjprC2l
IZ4fEQ7Bs6rEL/ceA2uCODF0tyLP7utb6k7emR89IZ6hIAV3w6X1kPF8cAjdvz9m
C1IjgaX1vmq6lbFPWE0chAm0Gn1LOib36QWFwtnU1RjV+JTPfIqjXYhvCPAdwGq+
NKqmKuu99R1FO2JKS03SihIBXqtopXnt0wLL2AceiU6pfWDP/dcNf7bZTACPYEP/
mtKQlxw/REWN4MDuQkSfylkpGyKbyJ/3M0+Yj84f3wltokqtKbEvKMk+yQBH1UZb
zBlcfmHJp1auShMwrgmLi/fqWeLgDn1GcmAyM316FOqIYjzfH6MzcHnCbAuLUsBW
Cf5X9+8GXI5LlqH3nItJoCT379q67d4qd0qqwduV9gP7nzaIcQpzOCRA6SZn/rg3
CZkpZIPzfg5j0SJSObDp+fiXdym2vFzhxHnt2yr9ur671x5uWw+Lm5ivRMEGa/Ew
GbnS3oNpRoJ4oKEU7oDSA9bB3Ty1Xz7Xmb9OFr2X4nWcgp2KH3L58Mj5U2sFxuKx
qx9VomHchsQRjxMwbPgxWRRpty8wuu5Hcv9/ChoUR/jY0orA+D0oAInpkj6IQNuh
goh3CUZoT+3/ng4kwqNp7cPoG3grxEs8rCm6EFmr2ZT+Lc8rCPpKtwIdyOj2GQ75
XFSTUCzVFBun+ZH4jynkza6eR5aL7e/pzT44Tnxi++kB2XXXUxZE2t50yGJHvWnq
hyQvegFAxSOaVE0LRc3xIEJeoO9N7LHmPsWZU0qGXHRedwjG7rhlb70G01EUO/2d
te0uVH8ljkdWG8Q//XZF8xoDJY3UAbRSBx+VhXZxecoHSOSt2WhiGXsppJR4lxH3
jDdXSqWhwCPWPyGUUOjbZanKgwMqWAU5yiLZQlbVT10vFULgG4MoF0q5RbD9l2vV
JkEi+NvJCSv9apa3nmqDkE0o+L4D2PmFyOgsSU5IMLymka9ZHmj1ZCvFuij53jQw
Y1rRbJxolAtsk82KzVXUrUIsxfCScwcZpEa8OVCvHK3185DCPfDLsQKpVjGDaq0+
YYol2I1OLGRxyp08d8ZE+egpCvjBsZe63KkaQValvbkEmTt0pcqKG2XjyvKpdCEY
fuENxDzmsAuJEB0ALlGf8JnlVdys0+NtzuItQLtV4L6/fT+3QNpo8S6hggJZmdAz
3/cQnk7pZuG/NcrjyJnfBls1kB/xj5qhkgQQAAHle+uZE6/UyXLaJ/cjgvAG1GGO
xGKPA0w2Bq5cf2BgyxRO8L80dFWzw3m4KOVd1mYRG+/k3Cy98WQCQB0j5O2mPq7O
IY6zfR778aTSFNiY1V3Tuv+lA+WSDIo8NJPCcH8zGaCgYBg/YWhGcYr1vjbI4vpo
gEPS7XE8mRfkM27mr1b3gPPLc12GN8LyjrITHvIZzkjNZHYryFXxLc1rskpLJLBC
4Ehv+ca5gTRyEEMWZi7y623cJ8mRIAieW4Y+Rp0WEN52uE/9R18ewEk7svbD99cf
EmBy8QdF4TioyI0qlj3rGtlbS9+HexRa7ZdE0dFNHNb873iHoeB/JFJL3Aq6vgbs
bN+PKkNGLRRA3t7KI/qxKrQ0VQxFB8z7xH5yTVidAQWO36TfP68Wyx8Vv0UKnpa2
nhA/eB0aTmwb0t82ixGOkecwXtWWgMKSFK/CKSE9i6f+5RzU1IYZyfJj+RBcRb8x
api5mYmbipAGbxsf4aU0hPhVTD90BPyZCoJPaas+DWOEKjkY0pLllci7Vc/ZLTuV
b5m5gBOEkVI9SxuGU06PnknA0LNlaKctSo9vyZA0vLRB57QoFU7Drlwpw/E++ypn
XbKKkL2fckugkZ0MspYCKehEPdQbw3ZUWw/A7o+wYZdUStj0yzhs3DGX2AF+KOUD
3accYff/74ZyIxHDAnyQGJNop2M5ChCh39/1CKUMmwyV1ouOuAn4rBvADqnN/KEX
Yw/n1mBBE86WmT8OXGZ8sOLLQ+M9P8YiEgCkRdycViwJlvDbaaMyFnEovpCnur7f
VyYmhf8cl7Pum3BV6F2XXY9NC0g7rIk9QNxVt70ZcJx1z7U81J2WlAWv4wnqB9JQ
XHsaJZeVavs7cAZj8CglZMB+KeRF93IOp9OcFrjJG9xfYbdK91cM5ZTQIgy8AChA
/AZNliJX0m4LeHZUsYw6/O5Gbn2C2bS6/5Hi+sbd03pCfTaVE21vYqmB8bov3Jtg
9lnD4BxVha3vp0Q2/A4hchk2P01jOBb0pz6JLlRmOly72egQPxSFF8feENpheJkA
CKtHiUzW/A6OUkxlp08AIyJ/svi/uhRMFWoigTfGiKQa9Mo0jMT5PLm4mn8DJRpt
fjif1wXsTKLH0iNahaJoLnxyMelXkfBkTMWarpKgMq+b3AEB0KwYuSCnOsbIXZht
EOECf4ygkTNy4J+QJxpGvTBDE4sWQ3TiM8vSgpkxxcJfzOobQ/EEuIC/jHRPlSmc
t4B3jtFPnt9LeWZ28lhfFR2dPRO1wNntpboY86bVChBlyKmbLal8QXgqoZJhwic8
bFbRLJG4xD/FLF5MPJ50CZ8rljS7bYWB0i0arLYcxFGLI/hy0mYOssEmgVpaTInl
WFo7+FjPG2837U92t1f2+eh67QYeMmY07r3rcZThfJeU7kjqkCYXTNZ0vsF1jeZv
xgGZJwdPXaJXE8ccwFWHh3PtLjHNBjMUrHr5OEL5M6kKIEtrrzmV5UVoK8MnP7rX
eH5mD1/Ggf51+cZcmPzrVfFgL2d1IJOucBmi+4ge5eqX13xh8tbuGDbRmkqvcLS7
MktADjCcfYelBtjyAkD3bfkkxFyN8KSysoTfX09m+R/+gOB6oDjbMysGbLFbFEf3
rNZiIbdooXIfBWKs3YyRjN5dfyOa0kTXEt+oJZs8GlUjUmm4ues85oKen6gCCB0O
rdhKlg5SFX0FtAWxam5mxGFcRO8eAXGTDceYBvaUngSC85GqUH3ZZRP1CDA7rH8m
6+Li3rQ77VfsAZ97eNLceIU0tgs8PFWl2OyzTtybVXAMRY3EEV9qCX2RyHRGslFD
fhiqjITYt0liCa0oOUNrpPaaH0jZPAAh9u2Ufku+u2JHHl2FRbJH0SE11fpGrenx
pCxGte5dWAXUwDYuEa70bIDPTUPH2ZwM+7I1CevlJN0lgAyAGf6HTb82MXFnxvSf
yu1+vFvhHOFVadc/wo03gw7KZ7bkStS7BBwQcwHSnyoGHswKMh9iEpgYr3PlfEdC
o2DrWVGflAUyovTSfbyGGtI9xWOs7xpSkRacHrNxMp7aChHRavu1WB5O45+qzW8A
bePmmvEHy0YS7cMMnNSH/72x5xe058tCJOG6G8X5wx/NwRnvzkokP1O8Rl4xfgcl
l/t5G4x/WGdj7uBjErjHwW9q0j/6nzOMOJwURrtYj3/RyVp55egR/WMXhWFCMOvn
O2bhrWVLFKAA/i1NcwBcUJ/bD+u/rLOMJW4EMmelMqTSRkTVQOtbAlo2UUNRf0Yr
YE9nt2GzMLf0WOzo/XQyOlbsGZErVtIRgFHyUhUxMykCvbHqk3pA926m8XKMlZa0
ZIfz+biU9UNqY2d0LmPU8DVNu5yrt8hSmuDGFzTNikOCDu/SoiI0QmOC1shh6OeC
LEBXuZDeMmYKpD1lD1qT6SitqAB7YM+M5QBQ8IBg4xNnK0/KizsEDHH/cU1yii68
znY/0n+APp0ruV3y8rJ02IudzYM7AHRb8qnARC1WooOTwNfRN19W+C2QfJf5Ev/D
LJqwJQ4g6czVf25x90A305oSUmnfxT1gYiwFwWw24i9dkV1La5DzlhEAatnU3UMQ
f04B1YjphdhYfdqDIW/WEzJawBNxk7MtigQK99sgd9aISQzbbK8nUJSu44Cerx+Z
sxToJkREu42W52BseWV4F7MlqzKXXxcyEhvUzizb/f4k9aTk5CaX/hmTuVZrB9vf
msGk+WvjKLNs7/fLRSsyLdH+OeeW3gCKtGp4g/WSnGG+wAsrwbz1E51aLst/TGXq
0P5hvKcoai+qhGSwK+qNxHrsraW9iKyfwuqvxqpsBOuknOWuST1AqcMzY+gXf77c
/7auIdpjkyWzwdV23NZ6P8bEWlb+RjNY+pQGv8Pmbo0dNlLxCwbLDrxO9K/eEdiu
wviLWKjD4iCDnCE36xiDmCmm6SOkIGwXem1YLQKKcq4eBzN1gOmM3swESKkFUsn7
RDO6M/jsGrmu3dHpBv41b7uCNtUKtcVTN71H2g+up4tVj6clqTmxy7Jf2pizLn+J
DjkLBMmF1IbYb4pw0W0hSO5iq0rf4AKuMEd448ftqroRikVwbxPhd2qDr1NNerIb
khYv+B0z+el8W1nFf85JMpTpQce1xP5Nd45zKV4mYuwm9kaMopifYTbQ8sIsiE3G
D7S88Qch3rV/CBVX+l5ZIiG31Dlx9WTNKJxDMpqUqbt9W8RoHr+TkScE8PuM1Lo8
KSo7/nRwESyqnyM7F9jCCZu+PNu10wrMJfk6a3oNE8MPj6dL5xVET5Z7Wkm6K3Zx
IrY9ENWFXgN222tZwjl+KJNgnh47ai00waJd4BLtqZ5N/hMY9jiT22d9UulQ8pMJ
HBD+O+gZzeEeJZ4WgDSJTukPU6haG6RNA07H+lslVCSxV1CqfvfTV0zijw8swExm
sLu6u45lq602Q2WIQj1tBjiWZXKjxaKwtR8p5xOcOmfVPkwb0Omp0qAVMdjkTvDS
tkfpuOpNXwDInOTbWiwoh4w1TGukygk7B6bkltbTqBrDsM3d+A0zz1bDoNucjZnv
3z+EouW+h0jnAcKN/rXHFk4+I/GTEVjmdXOvsp9tkCKAbS+YHu4VcP9xQgbydsh3
gyMLdkNDs/cYXE8QsfSIOiJHcoZiSswNC8s3ht1cNGaF7J08mDML5knranyHGDQ3
WjoZMgBOlPRFaF1QtP/YT1eSbUpH1Yz5qx5UtM1YOpL66rE7WUthWrvXfJ6n1XPv
7ruAg5nCC4QjEPBbIUrQm9q+r7n7GZCa/ktsYjOF/1TWOfmCdxUMq1/Mf8Ymudar
CndbkpZF1fN2Kce8QtWGGeCBwnntIPZZb2C5hYXq8AZNjGhA0IqV+xFnKpSt1g/+
C6BL89Ey3uQlKTOoTz0uSRkrFDiVOnoP8ssBnf8aB+23Pa82b4xmHAHuobffZV0X
OBf4fRBwcMDxqJ7AKGyFuxxcuZf+svnaqcoCHgTt4HJJDSDhXHFeLyauBOYHm59W
VgebIKRGFKaF4BKlX3Iokp2uVVbM3dmQx5yPNOEJrrRoiXn5AVgIRyXCeROceiOM
sop+nDmXa25hWruNAODeevd0E9VHCjvkxpMAPE+Iz5r701c+vKouFCElsMsZmPyW
TDqmZDc8XdwZh9nZm4Jif/lGJMjBiwk/QQkUhyV/F+UQQm+xoq6e+2fyEY8Ia+lh
1Yp7vynHPbShFGUHBfEF0z9/TUMvuGG6qeT+TSWSR9twE68WLQuImswAs/62Q3eW
Kg4fnJLxEuHCr/SXnRmJAU8kxgk5IofnGj5vL0WPsgBGTcat4vj65qUPTCz37Ecl
F7ylcscMohC7XGhhhdaXNqSNqn85bJw21QIT8vlbbHBI0ATgjklMk8m5I5fMT2u/
A/M9YevR6a08dxZr/1bNYFqfb+7S4PQbIvt6uDsbEp/mFBO1KXjdIa9Fi8TN0qVM
bh30cPdJeS20RGt/2uxTJmUV+2zV/fC9ILj0/5UOJwsRaSf7zsi72bW7+vIXVd8d
HrAcIfaqoAevRa82H4iMtKlmZl6VSCOkc3nJaMd7cJS4DmQ/A8FizUeewkOVB1VL
TmL1MRFcna6gaPnNctwMX9YRze2fSzNknPli+yb1vSqfXpKr8Nkz84tC6OuFFx8m
wVvivjGVzY47uKs6ZwNZs8qZTvmXniUnI8tGvc+V9bBFWKqshzfh5CCvjqSDWO1l
BXW9JqZaxQyZk+/umII1cmMYf/aYRcQ/fleA9Bq+/4u0XKVpFSvcRMG/G5+4a8Vj
1d76QZtyOjV7sd12svZgwRG4jCIzOXSsZ5G7joZpT2dL5KnMkQ4F4WsjDOBg1gJl
j4VvPwiMN3j5DUVqgrG33pXFkIs5XcRkmyNwORKFu5BtFDi6Cxd6jW6S7FYGQLoX
VtiKkGFilgMXQHduvpmA1whH6jfGWQP81/bonqlIQmbb7LyD4gsj65WFq50qhwH+
4lKFC4bCprgbdE7xWaEOoQfcuMIS5w+fnUVUOjQOeqYsco84Xy2WBgttagZuDhmC
XKY0wn7rQ3V7rJIVHBz6/gi2p4r/0NhTKClK0WEj9qvUwToVPsP2UOWrelNRS+I6
gd0KHjNxbwCgj9aBfaiGJGNPel/Lq2+FEwMmu10HQfpoHp+yuRPCS6HU9XqmYuHl
TGNjNiRkHVjLhXDEzbbIECa+I9LSkXupvbXis1Zki4bkWlVd3118hYKA0z0sus3D
4R4LkCrAcCtbJlwZCqB9/k1ROZCd7Q+a8QXU8O73JG2GxD3Fb+O2Xl9BF2z3l69o
fZ7GCDaoad6PW2jONVQGLfZl9z9r7yMYIP3yBKMGO6UP/g/hcSpG9hu5wsafmqLp
xg8u9XxcZiuUEUuiQA5cyplTlvkkS0yQNY+qzdT117EcJWbY6rLsYIYKJvJV8dCY
MSQ2eGUHuprhh1B3NUukedulyUEqjQwAP3o+Fuv2DXNAPcCnICj4djldLIv8xoS1
YYfrSyPiQzKzucfWsBZGjIxSwpisrAcpG4bp8Cx734iZnO6cz4pcLo8SvFoNpDT2
EhjrWhrfqVl5DAapJPyIe5qxBgbZE8XfGEN49BryLK9ts3Rz725SwbSxExEzYPtK
TKi4uU05iJqXY6wH8PjK/AQoy2FIvxr3umylxr0Gg2RC2nHb9d/yG6Q7USauNU3x
QRJG2FSRKBDLBdlD8JfoA/fl936qdpKkn2A1cRHSbcsEWpKYsu9tQJhBDB+POaYn
2Xv7Vi5Cm3WeehA4MrY5fobkyUfb61TNwr48lF8zXnQtVS4mb7EWutWXMnDRD2ZU
+aaHynrU70FgJoDYAAMsemkWhI05WdSccIhNKKBCmcSZYXUdpsw0ogZukM8WVbF2
82At0a4spmkR+/9gkyQXU+NOyihZuBhr9DH1vGUqUcZxSX4pncXc2mgoRVGbfqNp
CR/5J65x9QVr44xNAIFO0dAdofmaqkPZk7NKMyiLGxhwLJVqQLoA1fBpcUDBL3zM
ynBxSkzFDZAN8q/ofUCukkL+Ptxbheutc3SQ42IjXUrz0k4vEPKVOnjF4/IFO0Rx
ukepHeK7rtRvcO/25I4rXGUk5V+8SJEXbG9FXD82s/ISQr8OVx7FYqf2ETMQDv2U
KoEK6R3SM4589O887VKggO/L8/XWmTJ99Ax6G/3dB7i6B5BtdE3UO4vHd+TK12rz
L2TQ8XRhrMQdHDe08yOVQbzRjAnXUOmcUfP0BZS/yASvCfYMVIHHFOintj2YpOew
ww40WmFXp8hRYlTgoJk0YwtHdm7ocRcTi1luSlPh/3XwsDI/Nys/A2v1bFanJoMp
kgofkBHGlEYjI+3wFrs3vLJqC9lCRjcc2gaJBVyTk70DTkzoCeMKz9QnuT1xakez
7gRwKGcKeMidvgaTzKM9IR/8NSiBnfmhl6dDlggTJ8Lgi7FBk4sy2aaSMWaA85To
fJmoRIKr23DfXnoWw8uog1VB8VJ8kn9eUMUsbxXBRIVlY3Ry5abNzAVCijtd/lWo
AmleGfO8nf5iKEBv2txVpSuA8PrZIXitiB4zYaOutTGWtJ0nJ7FrhQsoZP2NB/9J
E2Lv8iFulQJ3GSM2yRP5Of5vHNlmZvnIRHgtw6nF+at7l2MGVK3OvfKWP+004Ajt
S5mY/8xWHmZyunQf8msqmQnsnm2Hr3Jfilj7DBxcS9sIFht5RmPpqFQVYr9BYagx
7SiLvC9nydW+czc5iV2AI1Y6UxL9/mNuH3bzZf9xEEqxVx2vmPAqllgIyq+E6n0h
uGM64m1bumhjd3yGunGpGf3kewRTvkkb+r76aIaUfeMPWzC8MZrHNa8srlvYvg+w
UELoeINtfEjj4YJreDrkoUHXFPXx802cXjoZkVCdBrenwJT9aD9OunKUpEtD2VgO
pxZa9vv/fnca5vRfBt6dp7o7Ve1lRt/rqd7gxxTDahQGdy//2aA2gDKL/6ND+6nm
ogArO5GAM8D54PbVxbkYeTYVlZBf8DOS9oGS3gAX4xqNykdbvZ2nKxBJlt6A+m24
IY7CqeMGqB8ZH72byiVJpCbvGRIDkV8gTkBOQZQH+Z9tm7B8vObTEccAFrZro8bd
LYqe37BucOpVVQdFgHpn3mtr8FAC/xX/qg61gqiPD3B8roZ2EPbCOQPPdq5wLqat
FiHzLBjI/XVnphkEPepXEVlND9f9Z2LeWtI99VU4vJ/ACeK9dD1tXUdT+Drw/1/q
eg4PnrVNHwpcOXdtP7+j4V9YQKHXsXqS2C1K3oh7wiI4WVKpDk9rFu4bcW9FTQpQ
IGiKFT+xECvvBUeeUiDfW7gYxiGfy8YFlvB2gmvuCIEXgb8Uta1sKf7ivcj/gEOC
stk+u51BoEyVkFgv6xS5ou93UIzrcndMG35Wdu6IxKTuU6QkYVXu4LCYPcHFKq/K
kHqz7P7LQdk4UpxrSMV2xeCIVRfpK8yMcnJuvA4TxmpSSfQXWEYbpY/j/yCiJyIQ
lvr1Br6wMRl/Zj2qQ8wjBdpR1ArBJUd4HdqWhU/EnrBwF1MXos79BNiat9rzKT5l
E3vOIj3kQLPSp6Lf9Bfkt7gKnUi0GxVpsgQY6nR3O+R3yjHgdFiF2s6P+ZsMpXQO
SaZgrSNjdKxmx+yx4c5xqoQHIhN1VbLpObwldInteJf+QW9HD4W+plkBrRrvYBRG
VUG1W38awMsOxmS2ynLYp07p77rd7z3Wr0vPAry+6Cq0jNDqi6Y22LeMKjIzauT/
pSXkhf9PXoeEnZAjvyqvLsiuXzTBQLDdFR7BfcAScis2M7vT3g+1HJr4bh/5etWa
WAOum1Cb9zyNz0H/msWl+mwSrsWT4XuMpcS3D3VIZZSEV4vSPOCSGm8p7roQ5IwI
hlnwvnifE/6azq1MBbVLrZL0ekZCC+nJJXtpPYsgLvMoeHHlxOQP8dP/U2g3744R
cxVxEbyillIiOb1Bl+tr2T7wwfGpl4CukbG31TzEHZHjIDLnunORsSVYZJuL7Rpf
6hYBIFlLSjsYE03DmSWGa3oqCtk79T0M2SSKcQ/DWS2C0pn9EfaLQJ/+reJExdC7
qwr0ZGQr3H1TMi/SwzKUJF5HfARrx3QauHXlmaY9cQ+thXy6s0+5yE4M6enwDnqp
SVaru4k0vLwqW/gC8nV/rNXvB8F36EbEon83rcSkFLsRt0AJ7YRM1btR6S4t8Lgu
BE2gjvfkwB4Dx+qCZAW+YKh635my6+ZlaCS1Y9OdyPbBw2slfLun6iOevtBo3AwG
e7C5q2Ebu23MlVH8nt1O8/sdLBF7Tm0jPSL4zyaqcYmJygP45dtxwMnCVaGcV0UV
sBR4EwpmByFqhCKJyo87acJnGtRFUMUZU7Lc6eP1zG3hvUsfi22uHnQz0aXOsPQe
fL5rh3NuYk8tCvUr0pA4QvfNTz4l4TPi1/lvP8BtirKchD0jd8VyKez2CKcB3/GE
5grjp5MSFR1M+wYIaXH0ouyrr83rzcfv4AYxY/QEedHpIYLYYDjpWPj6cYrvZLFP
pM38Z1774rwrI1UJ/7gTbYspwPML4YxI8Q7UxF+3+w7/cXJjPiuYnfv8JdeIlMby
8qAl6JdhpJCkUjNs1ajhNg/iqF/uUtx71jXk26+9rGcPlJHvkbHlBpgx1oJSDqvl
97B4dieYLDa86uqU2fgME95syyjtKOMl+jbMKKqtitiQCn+JJ51/hGmF4tdwNV0W
Yh1rvrUrUx3rTGs9pYUd+ch1xDCBkrN3kLkgpiCTv965EwuUueojMKGa49sQdDti
A0Rd+tHFP2dNy5bRMQ/fJniVBUCHu0XJ7FcPnSd4tS/WPV4MXfCet0/luyzyjZz4
zeadQshHK6Oh/y9C4ld9K+woK9oHLV4DjGg/ZxY/1VYJnlkWmAuNPRg4+Oxc53ta
GhV3mk2qgy5ZaLKSoUgSMZUekbwLrmkL7l6dFauQT7WCPNIOhUFwccgEPTJj/TVW
7VvrlTq+zK1U4gHbM5kEzbvR0YsRySauCKjsjobSwqnHp1xejTc0G7iKtlZnHLKl
BrqXR9csrmukDn4OwF/a3nCMmx2koX6QUz+LffJxeCAco8IgFy+VbIpOE8pLAueH
0dB8WNse1MsfC2vgIPPaFqcfHLdPpAVQk9c0hEoBIydobOGr9pglJj+lDkeigsGB
dX5RgEstI0wFzI27ZwvtQIO8jCrng7iKogR36ZKNx3Wr5sa3C+GS5vQ22BY4IUEe
1+RNqJB5y7oIfZ8BhWhu/FbkdBpcQzbKQ7iJia2Zp1LvOY5YXUhYEakRIgU4vPMF
xahJaaZQDBwC2CHUkxQRLGDlYjayaQ8WovbOxaSjF0bwo5QThqaAFobdrnIRx8c5
+DXGiWxk/6P0/xoKrMIQggS2R93NFkrnsikNg+NvLdBvBHJb181f5NoBrgukxdhr
cMmMOv5ZrLj24ykRI7nhe97LcqpplxJsHh4h1Yqe+umo8RBw5H2fMAQrd8s0Xoh/
MKsH55jUyxCdRkF3dU0yZo4ZBWKYMzSAtWqL1h1pPhfISszueHfF/o3nU386Wban
5+MMuZ1E+XGc2vKXSIkG9Vch8OK9zmk8K+u7F0G2OPn4xHDLyAaaKKqS4sU0sVle
QJmJwArnhVfggr63leZg//0KFSeAXCAt225gT7yzIC/ZkUCOSU3h4bWBRc8l658W
gIdTI4fOKZbOb6VIte/1R68CtYRm6++X9VU3K7NdbxtIo43t2lYUhCWbxLvnqRaC
r2FrreC17QwAaOnDTzTNj0qVcV8KE9drD9jsQNnHm6nf7nAOkYpvTnPdxhrGEr+E
gg5nnaUpZXD0hxCDLEOOx0IPBTCrSgZ5Aa4j0058DERqvq8kLuzPsmZfbiIm40Gt
8GLjZ6DpwVOIm9YoiYi3Efr3y8/TnkixLk99H4hXj55vsgmfzvM36YVSdK6FgF78
5v+VNkMAOGmo51TXzzyb2aD/cSmKD7QuJMZiaS67sEvdaRqN3zWQDcHok2ulsNpa
B+A7Moljzu/vvvp8K0wbEv30EZgqg4n8bDEht2Sc9Hdbu1Lxdgr+Ikk0wfuZ2wlh
vRn5hksf6cyx5LjNtYTJyvpxrufkFNcUUwJ/QMyWx331pVQYDcuRBQtVSUzKdxw+
q/YxTL6ethVh1AVfZWT8KtWuOYYFYxsU0sR/aj/+7VToo1F5cU2oIC78YvMfcIDH
sfU6afz+0yFUauvNau1krvW4Of33r3tbhZP1gB5AWSTEOLKVTvGZf/CXlWQE0yUF
p+v1EDU2SZ3LkmSbZ1DEutFb5R43JHCbPGHYEhM6vZCAy3mWyBiJWIAqEfHmr3lD
bHQxRD0KOE6QcXfCjAeuoWXLZNFQtL7XqAA7I5snf7LfdlNvyy4BV6m+lttjOWAB
fvMegIE4VcDsH0GT0mkvbX1QFMARb+RPV2EXngKJr0Ci3Ov6V4IZ0q+tbWMLVrUn
dgYmTaTSr/I9qfRHVZADfSwAHBWVHOwr/E8/Ize/t+DGrW0SGSPJuFlfMEUFbYBW
X6KnMe8VQAHllAgrzGo/sJ+9g/EZs/T2OW3/1E361n7FynLPqW9cEkqr9wZxZiKe
Z+rLbC8ClyjaLhsR8h3S0mr2iXqbwqVJtdDvRCpIA2KZsyOTFKCVmtUdFE67lxbQ
h2QQUaG+DxqtNcoB0HV+qrgWjZxkoC9JyZxjaeMWebZA7G51cDoMFEFenTEdL8MG
vyHSfhYBxacMn5uD+Un5pLO+YewiE8c9HxAbeexs88dTzgX1MgUR0F4NQ+CLIeSN
TpiODITUocJ2812B5R/wiXp6l2FWjUI8xM+j/pFxgDNKlUC1QIvQSMB9sNWReLrI
ixXFjiN4+ilJR+7WWqctgPC7tOFeUB31BtFnO0/uOqqfVReIbDA8iUB1Q/qza9KV
AQ/wikATmSlUMTQQfi3de7Sy5bWADvEuSQDNFLTM6yCFzWyFoAPc+UhxinD0CfvL
oqQoalmZe4nLFq//v3v1nBDceNMr71lUb5j1GdwUni+sT50W4bvAlmLP68CZfIXB
PrxYRMrpW5SM4EgC8wxx5T9WKOhN1QIn3kQkCWfcgJv+Sd4gLgU+bYVjGokfaNV0
zsKYrtYA0eWU9t0D3gxfjOffhT25i1Yk6MkrPSg045Fwpkp6cowuvDGZFk+x5YMQ
+Jb0rRbRnJ5xSt8Zt0e2wpP5V1mnTSMx89h57G0Zv3rI95uW12AjhkaKq25ERU4k
V5ayZhM2OkueW36JN9shEzj7BvVoepHN3iB/1lpPZwfRbjJ5R8vZPcKd1zTg1F1H
i5qG0EfiMD0EeFCVnIVTzsXi3McJR4xcY26FYOdsRU+j+hTRwSWogdhNOM8/2YCr
sag/o1aSKS3hZuRQufYI86WmcV3D05aDd4KVlyuNmNl3w0P49F6J5PDn94LvYcOJ
a/7p4BLUrN2xhYxKys1XnhGbSkiIcgmjBJ2UkayldiuVFH/x752qFMWJsL0dVqcS
zODnd6KIZbKnSn7Ip/IlhrnBDb1sJAPAC6arOX91Wad31o8uTLYcOGTHtcBE8c4j
7Mr4b+lQQ2tuU+r2jKwyTRU6LGllmceQ4GRKaGfQoq2Bhq62MNoATzFnDTr9AYpV
gKGt7+J3uURtJnf/fn8hsi6YzMghP9tfnApJdT2hN/T0lu/RYXwi8cLd3G0kJP59
O6MfXtSV6z61x/vBTjA5IpBn47Q1KtaZWuyefd1S8MeZ90da0ap4q5V1SF5IwNRC
aJnZXUvXsow0N6zh20h79rBtuUElOjavwm6Cb0RNbg246+Xen92PcG4NdwbubQgv
UTum3qWdNsClWXR8851p3QB6gh/x5K5ZbTz0pqu2iR5HCcloGx6h0FPZ11fe9KeV
qmK3Z55bo8esIzrfKgvW6VZuJJtLDB10Ev+RYyfjQTWNN+Khrc+CqgnodG+EPonb
azMgwLTExpgvk8u2N95qr28/DeDlJCaPg3M7tA3n1Gglvtnk5qVY7NEGdSPAlk9s
csKpiQk2DGXoHR6xQ+Igzo8tWN4dfuCOS5b96I8tHypdvcO4l6qBwGdgpGhEaY1d
Z5pjFkZ4J3nRvJvk3gFoJYPEEeDgY4RzpGb0jYMmn4yVW+IrRVQ7F+pxEPOXjjus
PO9Ub9aflDVowSzm0H+1KUHO77jPOOtcJkSz59JJ0WpFQObV6gCKWK0llLB3MNjI
f4bNvHKGCBkXHzZEm7k70Z3xHwQ2+mnXT8SNvrJffNZG3MQ2JczJLiwQwKZchFEf
g38i8xBeh7sBliXKEHb9cjClp0e3JECJ6vXuF2zGSogBnOju3q4FpCvMXcpI3ewP
aGG/PoQeXOXo5119WaDSWvatS3bLfO2ZnTLrZbPkhxc+HgtxOZxJ4Hnv6UIcBa2W
rAlIZGQBb+2KIbB60rHcMVHkC2ucjWxP8Xhgjq0hQJedPki83/j1kyWipbttPNDR
5CIiUe9QGjQCKtslxOtm9rCeTZ6s9OipTpjHs+z6yXfnTrcEzHUHxBOTc6CLBLdo
WPULYRjOvdwTbWfP+5MyefF2RnAggCRvOl27XpPmem+P6DOJBdCgtD58m0Qaiu1S
AAuvBgFQHqOO/lDdA4OApxZ71m2zOThWDrMoEXy3N6nYYOIk9i9/f3wmBk13glnZ
rwSOYw5DYoiHYWHE+3vHx2wlTTdN4e50DXB7rhxF3Qm6mCloGRL5eICpH2mWHKV/
h3vShpSjcTWuq+sPpFwHC/njocbhKA/BM2x00yO5Lsq+JUUaRhJZkoXk7b6Snk3D
ANDxRd/zEYO635POFO/8krWlzo7F/XXv1FEJXwbeO0hGNbtneLDi2rElSWDVpl5B
0n+tO+gTT+cDGTpgml2bhvBRpZ0VtcPh0vkgczAiYjhFYBSw80ed2LqVENf4ePKE
ds5hK5Q6H5ay8DIrbVfWfTQ1E5qH7CpTBZTORCIzr4qfORsz9Wv9EpMcZ+sW6eP9
rnf5zOZ8gWZ2Jnv74W/Ws1B1uVBNCBVp67u3JXMRxay+i5igo1Oy2XfLNMYly91t
nXi7as9PwvNapo9ruYtvtO+ChUdgjNsXqL1SHqg0jNjSpJjlhEkiuB90+t9tvm/o
UUf09whdWAXpGaq0Jw+BasSWtS++1lHP6HLx5WSQK20dbWdVd6u5q16wqD8QIpFP
DHp9Iy9A3z7YixH59h2yHy3HxwLNblub7Gq2gAFxhdLFRVZ+50+qkQTINlAc20ZC
ry9VkbfharIUUfcfIkAIRq89BhYsKzULjHjpRsNpg5HaRRPWrSlnRsxtYa/TMjUV
VkrW5WKqDKhHLGfP9YIgBav8dAzEZbRhEi4DNk/dixl1CEv9He1AdL7J16kajgb8
LGJPGtDdaHffXV+PompQMuvq/9nQt4dXqTNUcv8W/u2pJLlWkgOuLXvvUNSXg3MH
X1oMh+xmKu0CXLe+BxY19rMziTSlMfkKvb/btmu5xi0tYrtiQjEUAjf7zw/upVjn
VXL8/vbPv/WDgRLkHNWWD29AZCEQfr+NPvC8gkB2SgD2crdyjg7YujIDM11wwBff
BN5zGgzF4/zpqqIMVkzoXz0RvBQBWcSNvfXEUw87xke8pwmWb/sw30Q0vurBTZh1
X+XZRte9+5mXebF3bzz+ajccnXdzuLvmDwQHjszrwB2JHzX8Eh0o+pzE7x+Raj1l
yYpuKuqH1l7ugCcQOst3MKym5AuKTME7q80mMuBo+KDt46QZNgCOZ1AWf2+Lo1W7
MZO/ZT7vl4JqeNUIeMleddUKsIEib3gqLpChF2YB02ydT6cSf0YppCVetM8SGsuP
3Pqz+aea/95Z8xqBgugduw9D4fPRVTxH2lBvIwJyRJntkTrkQ+5DJbnZagylQzf3
O/GB5+mwJog/VT0BzqHDhwf1nOkDK8cumxgm86QUXT9Uhlk2CsrscMJseRVvChyb
RBjMeFzyFwDw9gb28T2OMhCMO1qfW3wVL+DkpN0eELNnxTloVS5loaHiOt1+D/og
BMSuwASXiLk/FywT5QrzIYKAaLCdIgYqK5OJc1abE4CYplRj8u5d554pMGsATH3X
w7UHMqDRW22MxEaiH+EEJJz8nKu8XG+c4yweLqHkhxm92MNp6cS/W2xC4HGi0Aft
F31mRoIAPaXDp3HGcBvelz9Z5L1FL0c0s+X9cNVdgKLxQF/hnqNZl2Sdje47vxXR
Pb0KK6+x4Z6FlGgamJe6XXRVVcasftqcw7sGZ7JWTug89xNO4D7cvm331dRVNJrz
cpPNw+puWNuNrf62zN6vje9BTgsgsbXW83goEkFpYJKlGSA/j+ST4Oa27ZPVfBzx
XleC+sCKQkR9insSZdrr8xM6gA8iFztCtlBfAO5yJ+EuJZFoV91zca0VJc6n5xmw
v/k9WlhHbXGgGaC72I8Pqc//lObopLhkQi6KbW4R32HgMYira4HAHzygygBf4hxg
p7+hB5bxumP1U7akIvUrhbcB2iwKxsHZcnG3aPkitbS9sWSBpNHV5iOSLqxeXnDS
SxJnb3NQYakvj6d+zUlqqaWT061h6BkRdtNlmMyU/oxmZRqpHgoU0tV86XMeN0/I
ksJnWWM+I7KV8ZeXS8lsc5/VbCaONtiqPu9xVBQ9KSccdHPhGE30rrMTZimYhKSU
fHw5eAwmejXq+71VRtnE4stvHmGSr78zcNjn6KPiG3AfbAqqLTePOrgacggKCRoX
KRgEglskY3A+hlKvDYg8KvyryBko+zwuFZCRJh/M6rzROSODRIhljOB2+Ab4PTiU
GfaoLSsv70pX1z11bqHN6QRnedLILDtVvilx7RKh4bJOGkiy/WWtdpXVCUMHYOZm
q7rpv0QakdF1KQurcuTO+mvONY3+3TstJg8AM3jAYeFrMNaw0HXNWFgFzew9Wwua
Aq5Ho3mX/41aDLQ6kUk/pt9q0kuQEP+hxbonzvykHxGtANgoy3kxAFbHacDDLPs/
JriRH241nRwA65E5e/vun/wEH7NYie+G2zX2A4dWAg6kyAIQtwWTy3Mk1ZRWalK2
MiDxUb9i2xzy08BrRbelu6pT2+m91IEsVsT3o291jWnldxgMcJbVEpj0eRyCGZXY
3IYP1eoo21N1ZDa12s45mI1Oqh4M23fNH9zJjmymQhH4lxo3nbqi0j6lghCXYKIC
nZTtSkUD7hLAU3qdsdykTCzErH9+NJvSCTLQikiuLU1KIG+ksQ9NpMj5zLdWNyZl
idwKY/lZznkbg1W19rR4hPoMfdz9/J9w7zkGWJ5Y1qOiZJetHCNnQDm052Biapoj
8ImwuLtLKtw+JVQY5+62u8YsFndgYIlaMxf7w9+eHaXSODJQJp9D807+pZXkd26O
Z8cV9wJXWT9kRX7/mnJbG3UtxTRj64jGK9ZF1bIJsCpgIzE2KyNbVPlpF+e8HHv5
08KuXmeEDz1Y1scoj5JfPTCMS/rBdyt5jXfBf7SynMY5nkV8u8VPuW+lrZ3RSs42
l12Kms16roSWpDMjk+rf5l2SDbMHLsftuVGhAlc0zjhrgOiOQC0ZKVSQbcoqzJw6
g0OYy2mzML0pK1v7oluvub5hgIr/XWbmvxNORf5XlZTfsmFyx80KSoZPf2ntCWj5
RCY8zmWm6yodXU6erjI6qp4o5zT+VM//XLflwgrvFxCxemTUoEyg6XJGEiFUEg2R
a/EO31MEdqqP3tJC8MBWqV99tn6SysRjWm9bzrkaVDUbZUGcvYqMWh4fB1DZKZyO
QYSQVeiiVTeup0bq+D5SPFfJ32xMnwEMPxSJtmyON9ozvaYJheckcqPxwzFMzwRX
fC1FNPcCQDBLWTdQDWjeBLcpGQ5YaUCL8Ih6aginOmTcu+ZpMzg75fT3+V756Tfg
dQo9uhkDOTtoalOlpeiXGx7CA1/K5d0vP31LtKY1bTOz+JLH8DFLqhxAjgm+sCLw
ffapTc55nTWRjyce8fIwwVAcwo05iMwU9CFbDLJpK6qyiOQQH9jYFl78nNrVFXW2
N+9IssnEMkWLUJfu1JlLdrzniauoXHJ9IioFxDWNl2NToO0vNHG4Jp1Q+YFjTQM7
sfmzyUkBlOsVfs9cumtkVDrl+sP0vm8zqFfu1ktUpld5zgyP7XzgTDLsOJvO1B7f
YOrihdazkCNArCnAcnE+OtB7QKQja48LgARiWo537Y51yf17zrmEcUjleRy0BZ06
wPs++/aW9gBWy/mafpNBSzhEKa0c2JUeWR09jnNf16j4pOUdLURTYLiV6Qt0V8ws
dn3XMfPvgHTx9WOgUeFmOeKr2CAngcskb1NuR9919iFxWBSbJa8cBvROfjvKw/gI
hhe627VjQajCr8dkj8L0DIJjq9wsWzFwOUIsvMfZtd8IGRGQZfWFFUVNczlbPkjO
o+kbCFBaJrHw3VkfA59mc9swGSCMTq+MfKESgsxMWwXigR1xNzlQBkwAYEgzf5vA
VXEdcCyAoFQ+4bM9mlsU28m8Bg85EHSEfu1hHeO9u4vu/Z7l7LeGythDR0BwJf/B
HddFvCpt7m+qursVp5X1wCOnoaYqFTKSgVoV0rAcOmB0qLEAy1GAHW0nXEbx9L4W
3pPeuXvH/rr1VjJ+/KA828G+BHqPlFiZ7QwCJG6U0FUYCLrBFib6L5sOogC3ogth
LaA3AAN4qTxilm611H/a6AcAoy91NYKd7hwOBIG7wdWxA2NQqJXPC9a4a/B/CFW8
Di9oMMCFfH1vYx9GHIAxvFnVw5dqI9Dcr7/I54lEIzMZEoOB1z5A81kEoT0ijEQ6
mPOCDlUnQQRKrXsG88sVdBV8Lamb62iiVJ/JZPAhvi3UdaCx7LW2jo5Go6/j10fN
COF4pSYHHSHEMx8o1yHo+vBVZysX2g3gqxxTTd65wpVm8E+r4FM/6YuTTQ/85vba
AKFVapCHIUf9W5C9j9WHdju/TJ0k/ZpSFaZPQnnlGcfBmkfxNHIXu5E4SHyBHmu0
cj4d5vX7fN1yj4zm0p8kLy1cbqDRuTjhwMqtRAMy9Q9srFNf+UrxUQX/y7AKzL0j
0lLI1UMScvWFd6mkZzPjykXqoE8xNju72MTtLDWSYkpgTJTzUfJaTIDbEWNdkKEt
kdRjPt42OGEXOWo0fqdKJ6RIuRxLhvr2W0xXeDxQTRdv1TuCd1/8pVp5yEa99lP6
cwwWfbzyPNB8KjbeoS0kEsEaS/Tm54puk9GdVa7uzahUC0c77oIu9SZxtef4pFO7
SmLdzTxr9KrXB/jc4BZdbcWm/MsJgBCVRJ6I5es2P2nIw48dsb6lYtKfsDOj+2pD
VXAb2yyeEBxmkrr0LqDSD2DlHR+Yr0t4dAyctfEy8XOIw8TVAgBOwV6A9U/6wiQ/
3F0RlmaJx7sK2LX1iNBtMp8K2SGvPLh/RCdvtlDDqerSOpF7LXOl7aUySKv5UJUb
JHkkzu2KxNRRLZ3renUTJL8gfTTpTSEE2TO1FYfU01AcQAkqU1it1nnBDB2ueyTz
DX3iheEJwMbjSuxyq7AoEtDBHFgN5vY63pPop0fd8lMUeLhxiWmJiYNOa3zkY+xD
kwP2u7EKSBsX3HhgFQOPNEgX3FmJieFyYsFSKus1IbJ8Gy7slJVIVbAhDfpAyMYx
7sfU3hFuM4m8LXgfw2mUXHLIoIUGd8xnVZyCsmoQvUl60sr/vqzKwwpa2trJx/H0
NOr7BsIUhgQSNxnAhkcQwqYBjUsUyAlPWrXs3f0jELvgodPDrzwK/t6MYMifw8kP
zX8EpMu4QWpYwUY/HlifavI6BCEhsR8WAKGbE6CmLLBsdFVf1fX1FwaNiqyqtfGv
26jfDrr2CKdkpbn/fLMx44kG4xfC+6Doj6SLWwqtaoBN02P9gtAK20q0xCPM23YE
C8eT7JIcxEvRNVM64iqCnYVIbtQ6iDhOadFIyktF4xau4PcAwE3K3ScB7Q6QPsue
HSixGonShobDCdlze4/2tzh/ju051NmABu6kxpXb3nYd2S4mE4N0ThPNvEr3oMJB
MMSxOtmFDAg4+9Xz3nAghQFuyIMXr9JzVBNphmzGkl6r1KpEgJiICWGJoB768+Xs
F5yVYtht/JcvdZB8JJrrmxFzPsO8yJoLWwtIfWTWwtz18LaE5FPOQz2GsBarCSLp
+lfYhu4gffnei9lg+zcFfQyFbHys6lYKjabYTeHfxoOkuOx5s3eOxc7egBBd3y8F
crrhIaBthtASd+xYTIoGWWosP6bhcRPct3V+mhHKmQO6me2SHg/iL6W4BWKuzBJX
ELx0pM+mPKYokCm3opEWDQPaUZFCO4xmsE4XZyE28UnSUsPuAB+URf0NvCXMBsBm
/x5aXaXLIiqOvXCIonUi3/RrIMwbtOHnb7DmF4TwxtV6uavgLMZALlfUMogAfZwH
wmpR7XnzlJGRKZGeF9rKVXWI39qZSWsqrk7b6x4bcAn2Ipqqv4wWHLiEiDJHjyum
YmmITnoivrsoc1x5uYsuBW5AQQifzOygfoYpJ5J7cWNw5VVwdnoMv4yuKX6B40Sy
rC7BwxBuoKhhVlKVuQZkzLF+pqwcDQg67hT2S+gX+3vZnZQoJc64mjoDqxYbVTuy
1F2PF8BQo+ERs5evWSbRlnnC5Ov5heZX75VMKZcD7t4/vz1r/CmkcaRCHdqsovL+
Sc7rhoxWA2hN0CdOjyQnvR2dtkymwC+Kzxv8ciHS4NK61rtzt9zS422MF14Pbw6n
byPHKz450Kd9rzL1f2fTq/9f1WkYU1O4NI1W8Do8F1JqyBFB09DDsmqRK8uwSsha
yHR1dhiKmdppMDc29nYDYR4uUqIh7kajwUzzwhXcNXViMc1VGHC4p01gD321kpvJ
D+Ztj2IcMM5i8EckNxdUfDzGYbDTYGj9UPobTl4PGMPfQ1brjLMjQ0xIFyINwaSI
AoUfPH7PDhfoDqrwG6/tQQhJD4GgL+E++XbGR0njJJwgiFfzeY7L/pLYU3wQ88/f
Bv3apiqpJFRv4m4LxmEuUkU+SICbl5N6FmclXTBslkqmGzt2hwiFv5dRKkJewgWG
rCA20LbZqYmLdkUC4F4tmcaYmEenyOZ8v1WzkDiN/k6AUeMV+4eNJlHOQb448vam
YncNnjpLdmrUHIh7pvIj2bGKgllRrhbd9MeJBiuVoA77MeJGayolL4nus7RcPPmG
k7RzLWX/9CU4uKtpxqJ0JngiN/bmEwGm4FVdHJpOE2e1l+pGl9Djqf3yjfXnuhlM
XdxbBMEnCAdRGaD7gBeNK9nDSDiu0Q0nWlRn11s36HWoFdh6dbIlQ3kwjMNYM2oY
KLmgj98D1ec/iQLWOeJG9QXBo/e883WBL60rdURVeSM6EqnEkt7NnbKbctv1tSnY
FvYJTmjlppHUcR3de4spfC6kzAiywoQ/Nbl2/fHAL+zcHbHPvVdhtuORxrR7p4r+
W7KXd06bLtqXhFkcV3hROO3M8h73RLRq3s7QdzptJsXMnMn7+3Wbljxdydqx7zqY
E6SNhKYJvhcKyiwYX0yV6LevD2dnduaDI+Y9T8m5ElpvFpGQfZQuP74iDf5DrwZ4
LmDgtf5QzkKr3T7jm/WlOn8kNGYJD2WxO8itM/IDnhCXFY4D/xfEWC9/wzthIE/L
ITDo+xvgtw0R1J716H/P3SM2JIkXmM4S0s0KrTY2IpSCIhItHfmG77ocajGWiF1b
JAFc4WMFxg81e/XCxrp6gxa7R8p+xZuVlOFWdrxcm0a7M8/CxC8ZoQQeZoX1Ktd3
y6B1kO8Sfwk7ohnY/i3RVKOEiuLf59Ok97nQOTRPzEYSzsdOpJYrvaP35w6QMVkI
PxhkuH13kqpjBolGqY8LU/kfUnAnvb4si/D1bcvtwYNMfrTUS2p39UossWlL5W7H
xS1dnqEuEb0aS5ZdCcoJC8bT4qweanMqAeLj3DDeazxnW51BtZ7XMq5ZJAWsXG0F
sChIvr+jRyEYOvmXjPwHDS3xKlY2oAC1W4pEolupPScrXh1DBWmwTYNbkZp23DOJ
xoe8SED3iN5Alb2/PkiNtV1A9Jz1zTN9b7IJniDy/ekJJETKYJI9wYfZgX7Htlaq
Tg8gH5gaIpd0V0ND5fZ+XCfdMWQ3cWLrEXsYHYjH2utsdg2WbXapn7ny57IwJAn0
WPSFjackTx4CBMv9B/nO55yU840TtPWLAW3SM0kLA7O+jW//Z6s7BaaT6Kt0kj41
QCi/RYGK1BFuSIGdiwFzZqMyPdlGuzn8I6kxpE3hkaAJqL/v+9ZHwbNlWUruQBuY
psbmxM+vOgRRfIoEEeQ14IWOft/oZQaHrTl2H2U/yFwtgAzcf0A5E6ejmWPCqtX4
7TaD1kIDDi9mZVNbi9fqg6JVx8NLSecYT+6QCF92DNN1jwqWiYFL+AAAlP8FjWmx
7qaYg9zZZ5YLoghYto1bNcPu/eVIh9Be7kqiaJg9wi0dnzvSogOl/+hhjKGTtewE
nvbzxmqz6jVcu6r5NfhUebJGm/U5jqwUWMJ0ZS5PMfr7w6D7bFPpAPb8J1dkvFS5
iOldFvtRVWxPCuCk/szy9srJupboYrs6xOFzw73gss9BvSIvghIvf/staNJXMlOb
GZ5i0ieZmw1FLUdbNbAOehQjo01Ks58V2JI1LWnUxmRt5h9kLURI4Mh5NZIWKDVd
tcQQ/gSXfh2ecUrylV+XcfnrWBN5JJ+yB00sPlhvsdgcfzOtnhCn6inbw6fJFsiP
sJtBaVl1TJHenE2xdChfkT4z56Sph7CaLTYZljadPADSzWCUd5iHdWDVzf0kYQCG
+VbWNrPcMwHgtnDRMSU0VvIM+Lhu7LGq0kKWcWn1fSWupcmNMVq5JyESLJZmDTxC
LAtpgkL2sWopTFgc74NAH6H+UZs8YoaFtpuPKk/j52sg5/frgU6u8rCrhPdEZIjA
6yWWVML4BNKIeM8HEWxJdEQaW/m9xouYV1GUIuYII2R4Y+A7jX/25+pZVOV6IM/I
tQAFpiM8ScEhQxttjOlA9UNJ5HhAx8MMgZFM7mDY2HPj5jNVKXTpcGHsafIm/4FG
c0x4eCuxiGnB5FGefqDtx/v9XIgadBARcVjFw438zVDKl21IcZ2s0BVLYPMSwcKM
XivJkS/dAKLxPBolQ9H8mP3974rlMQAtwoC6yzBJdPOi5UWl9p4GlfR5mW+0VFo3
i7YTZGTGCe5SG5uCi4Ed9W6hcvpA1zPmIMYY3Xdy/bgtJ/KuJ2IFcIe3TIWDY+bv
TyuR/Yma/tU3LcLeYdFOr8W75236kuNRVDDt+YCGSa+JdYM8DBJCf4X+/i6s7i7o
GIEoPmC/x32ViXJH64oB0ELDkdqtFYc0A47pzGSp6NfSnRNtSnioPZbJ3qAHFOM/
+QGiO4Z6DggrsTMNjnvGjuU8e2tIzcQj84WXDVXPEnefc85S8EMXofuP6Z63jlZ5
juDrrlbNZEZdv89wGaMtZWN6tCCwyAeEdTKBuacDdozb83WTb/ZHdZ7i4kvo9dSc
XJOYIGdnKkuSZwwuGDM0tCcnIH7vTmcm9vtrWdU3QPWGMqwwsDoyMMOscrv3zQVC
ZdvCgnH8+TccUV81PgXbLku48X1TWqX7JmuvXkGxAkAMzZLvG8TlOvAdf9bNUWVS
zm2EMLJYG00oRHpMuaff7FZj0/cXwRVxAFMsdk5Z4uMVzmZrlQxQu5O/F5gquEH+
3NkNbE4JJ2kV4iuohc5/n3MhE6alHpQxCuVv4WngjMRnPX/i0gWurRsfWMjUBJeO
MEgXFXI8qODPET6sjl2E5/MNQyUoMBWv8Uiam6+iyyvoshknXwxN/khrWVfvfors
lNC1Dotl+/dvOyQkLLrvvaGhgivudY3zFGXXR6aoNN4zEIBMnwh2N8/UimLGkFYO
D22i8ehtw1aDq8f+DIX2Y2EIX6OLdKE8r6ccOwvcfQYOBy4i5d86oqMxz0uV+ZTD
4yTk5dhvA4wDkcgdtNKlRYl26tVpLWmmDH32NHIaE8Y458b6Alr/HVSdp77sJdFu
F4VAFc6174aT76NaFAud0dxA4jEbDHs+4nXcavP4LTgHxRjBu0qjvaQEUHZtXabK
aMGNPv+jyW6q5u+t5J5+aaNBnQSRN3VS1++1rqE5ZDDHxnn4P0hsnaqDUgi9w+bu
7A0hV5V+FwRSF+eAafPRSVpFPn8K3FLRrunsGr50phLqaPFNUIICvewJWTdPhrkQ
gfhbz1KHfYVO9ywlar9AAwGcSpB/01yXAbpZgQGBHaF/Mq5hdfRs7pjrTRVD2l03
YTsB8MALuV8nJTjdECiizSgrwveo016jioU+nIEJoY1KpvjpQfJ8HdzTFf7VCjyH
2AB/hxwZN/4RUw3+lj0W1rIiSZmI2DBnQc7SmN4CqU2CdMTIVyaoh9s19ced6Wiv
imP49PgMNa6SdpaUt13R7UQduwq/J+q8w3uABJhmgYNnAwbTsAfbk7TYyuUxjPVI
cWQFZ2KF8wb7qLr8KMsIVn/YFZn2Y2Uw96aWTbnEsIJs1tAk2z3Soe8cj0Dd1HY+
PX2SHZrZZm4F9nfY6dtWcUTTWSWHpIoOHKnmeWmyYEOi232O+3+I8+mbMpKkvGpP
4uTjgRxcCOyj1Z9z7HsMj7FQNlB0/m1Qq/pWBvR8Axuu5vu8r2soE4CB2tOuKMBP
PxMdY8Xm3LkFCW6p+dZfxEjAmzuNPzTyrmDiHP2zPF4bjrgBqQtZZMYr105X97Hw
lFWVollNLB+EJCj6LQcqy+OmpMt53avxxm4T7hQnAI59OSaHkR8YJKop4kHN4Ebm
h3yIU1WFopCIyJptU14ccHymIhUMws9Xr2FPs+PUQFK4c4fOabOH1f4EZqOJk/AE
cTf9IrtfEhYmtI8mqVKc98toMUFyCKJJPfUSO7/V5UF4dgUkG7sAbzHOMPSc3dU+
8GZu+LHo8eUzw1VxXeh1fVYMPUQDm8D9X3X34NS4+Q8kjfWCnVCcAH8tsufN8osh
MKzf7dD3+e7qsITh4nuVxK1JBmrHsbM4udzwHeco7vZX5zWG2FnyVrcUTaq2TBXg
rkKo+6DOw6bX7MiVfyrlR6fkeuGFvDUw44cHeTvRzROGyRZei3Jpd3iL55Yxn5Qp
/15KxjKb8auUPugJ5PgYt7OLAyUECydi9qSagLMLNCNuIR8HMkXDoPRArMcQaSSL
tI1JFkDMOvP2Pe7J7qXAtvFnTHrAGGrzh8ha8cCAu983xpQrefTcTFaoFIlUfiKP
MzaAVDbKRQ3i17XOd7KlT48dAyBQMZrBUQNG765JtfT7CABWwA270GQbnUZ/KDqn
7OHBbtmfD/ySpNWY+bR55jSdb7phz5Vvk2s9VVORo8Iyh+P8oHR8TcAo4pQPatSy
pBZHQ9wT/npzhNVJLWp7zalgGViIuIman01tzIpHd8jsT1b8FeRx0EU2KqOowDfM
q9qL+m/Y3D8SMMjLEc35/yClTvktsdr+aG5hChv+5cX07lITbdrKB1UxUnXNrHnh
wIHtV9A7J+s2mrq4M1jkU9onxbjc/YyOeuMdImFaM5vsQJqrmEAr315G2zcFWoUN
aoad9VREVR5FsqbBz0EkrY/UgfhHmmaIzqBZedNQPLiyVQ/Utyd2KTneRmWziaMi
CXQJgZRur5lwYGW2n+0kOfIMH99IKRLCb1G9oajMzgjaybL6hVlDCMm9qbQOvEaV
ZNhpM1CXtRZ7/+0yc+z+BEPat67qMXXsOWZUh+1GF1YkFZhLBQkM9lXNXhD82WCc
fezAyGdfJGv5ZfSRZNk4DCKaN69Ntx2IuSo25OB1p3v5BlRmEMyW1q1ESRd+DWXU
dJCHVbwCjwJGT+jZcP9rmaIFsjCgXaA4gQook5ZvtTF81S7NNOb/qCbqiwb0s5gj
HXW9lTipvmAE8zjiT8ZrzjjbgJHkrEDWBoO8BeTPqIG7v+t68ykUsTiTxXHJsGoz
nT0dkTq1SLe8dQqeo+1eDjwHoay5d2T4pGZtFznKhQMbBtRDn7l4WdywmP1Lg2gf
6P0W5rWHQS8bMZbZtNHVbHQWYUQ0pjsQfbZjkVe6GlbGAfLcDFQRZDo8NQk1Y0XQ
hibQoCZwmuJo5xpEhXKQAd3VYbVbEQF1w4auw9oAvV+lAIutkBmj4VehSgnwHS4e
Lt17IlAsUPwefJjZHaLMjp3089dvENd/T75lYeqWp0r7UUwA6o+ChhjeEBaGgT/i
omH6I2EmDsYYvOhLFcG54OB7/9+a7TmZMUEihVYJLldHQ7ukfL6xVMBk5Y6cjhpq
5hmKJJOelg/hxPGCBz81gD6qCEsvONTvl47wQCvLcLncXLczJsf9p0ijjf/1bZtq
jKD48mN54rqbInmA/wsjKZkx6YdQzPdvPKSfKylizjkff2R8a2e3Q0hSSsRAbqPD
/3gIjxubBNxS7HmvI5JYOXqgQMx7HLHRTQKNcR2Xv38q0osYnFO19WaLq6lxGirD
rf5A5bnnpLH2WoB0b0F8ssAU28KrY1r9ROzRpgc9FHBbWmEnfbfLCGtDrAJZ+bxI
P0fUbfZDmkH3l94Jpq7BY4z+R3B5mdq/0u7O8Z94fPDHRFLhc8rBiNsQzeP2pRSs
zcXU3eU8t2UOZmUdrWUvyqCRSnw6YL0AdT3P9YSZ3sSNtiv8qyn0Yc+BdLjCr4Um
Gy+WWRxwrqRk4pCbkjpz60w+PrdWL6VTBIt383W5gjWxK6kebDbmYIzgERaXWvl3
gFdOjJJoOOjF7NX9OpYJYy8u4PjYv5Gp5h2rhFUMFH9Dnt9No12nF2oItxnSZsZx
IbeUfwUq9wyAJs72jlWLa8oA9+cpsRJqYkzvY8gN648VDvYh1dhGqYetpmV0f/X5
hR4FGikUsUZbMF15LRy23cmRZw0YmRJodwYppNcPQcNap3Jy5fIIYDIK9CNoVV6O
4INyirRu0UoxyZqVPmj65QyT+hwnsPbjhFp4GyBX8KpxVJaWUn7STFvOOqvEo7Cn
BLl9Wcz3aLUU5xrEEQe42yEJWNwmpshRoW5+VBGFiUg49CrnIAV4G2T77Bwi+JYT
BcVmIySZaIb/RllMyJzCdYQeX5zLyGiB5Lzex9BKoQkR5lWDajAA6nuh0/6YJxCa
oMjr1D//Pr+LuHMRL4NnXCtX1Ee/KHd9qBYVkG5yRV4EJNp4UPBa4+++ogtsEOXq
rfkGQxOwgo/RB2OjW37B0jdLZnPaGv9EDZKD3JWBPHYJg9rhLfY7o0/8kSg3FDi7
3uqGwQB8zZ+4rNcqoYTrTLpPCaS2NUDMPgmcLoZAOX/y3l+nD70hLDNr0PdXwAPb
1ybjV0u5ua0T0gzrnKjDtAg69zbkRR5B5NapkFTQ2Tr94WgVswKm6Oz6BbK7a3yJ
+1n1xvRHKIvMSk8sLVbaPvHjceVRIpllPcDlVcMOK7mDXuWoWEAmgzjvxHzhZHAT
gPhBMEXcU07R7nycMHZLAiLpxrxfnjCoWz1q0Yl7XbLPpsfthh8NAxF0aj94JDxh
zfZfQn/Y0nHeFmlDufQ4QMv+zEismpw3zNzzVVHcjVxdcINajsXYXNjc/1zUvkj7
1On1ohz4m4Nqkr3OxW+Q473gFDCzZKYDE5edD+X5uwSPCOrK7PJ0nmi0ho1Qts8m
7qbdJXQUkplqKCivFYbkwk/naZgaON2e83+2hpFBMnlZrAb2C1+6m7bJ/nyufNTR
UC4FfT4o4UtyohQs9devU7Bp6HpdJ+Ri++nphzpxoSC9awciWEUWMSXawcK90ENz
FDz0Zz0cH3Tbp2FGv5or/2WdeAOZI4Cq3mDr8pHk+xhj81NMUdB5gTd19d4bXH4k
DVDY5Ime7L5renthMFzrr6vhowQncsBJmuU0NO7zs0f/Zo6TI6Eunvz+/1cubndK
dEUHD75oyXMsx0DtMeRNFBlfQBQXJrvX97Cl/JlMJNtzoMhdwGK/r+515+ZCsxxp
wXRJUQ0XDh/DukZegBNgkzzo/OqnLXS2G2aKCHZosE9nFk744kFC1d8lE7/uVybm
lWTYKabZJmmgs2hddD2wO83NHPcYwqf0AkjGQbVArVWcxYULJO4zfWeZTPmsgqMM
rKA+FRedDfjI4oytDzFkPWc9jomQ3hspmLC3tXQF+CQfPzTVw7IqmeWXxvuU8Js4
6gnyeLtgSssZO+z0jXZgVelntpVnYMK6sXpzG9ozo19QoY8aNuAkINFiI/+d4dvE
OvWZloTmc6gNE2qGgB9kgSrv5tJOJW/A5juFWpNI6MxvfexotLl+OYgSzgNCK+NX
k4fwsuUdgWnnIiRtOQ1I9za4X6+csUAxLjxY9leJF9ZZeJX3PGkCa7u58quwtSku
iLbU8tMR1l2jSCYBdrFImno0fBx/K8IAxB88REtMwsLwVK5KBab9PrEf+Uf3rZdD
QzdvRVz+QF8I+CPfqVblZYMK1ylwEk0WmQBgGDPlJojSri7mr0hRZP58uDXoAOu2
Q3FV5a0VXXUnbT0CCA/G89hfAPyn5jY4f5LtXw0V5947Ot6dMR7fuQGrdnmv5VV1
O1OYXgMH7wupjuzS+pbHP+dTavThNvIT4oV7H0zsCT0lb04K4/h1mCgHrJOUjOzb
4nvxvQWl6LdcTQoQr+XbJ9KkI+l7z/RdPfHL1lsdhQr3mbZLreKKFSbY05f491AF
UI0twrcXKzy5o/I1UH64Ef2WdhvbL7hI9+6c/tipvo3N0FCuUm8cw/xs52lDSTER
nL8lEq6X+A0k8zDnAkgMs0ryPRmutmSOg5KkSJUsVn7L22UGxmlAklN5zkMrZQEd
w8eBB8DEr0SfvDkhqQUDzC+7CiiqhI0HSbpShQKEb/alE/FA2b63sB0L/mc41psE
qQmCKZV8T3LwJqknL0z4gPVvdvC+VvwIwTsVizmbXixfwt1vxL7RHCbMxDH5nHNe
FSp+PJI4j5bu+L+mcEWpG3gaZZISDdVKxqPxpJBzN/f8aKUZ+ssiI0yoC56eKMuI
K6DXW+HpYPePJahNvKstgEBTcduTo3VtdqxgW4yjEMFDlRueoKLDqBrvV1vafBjZ
fuKywicegHNpTjiB9/uAKGVQNc5C6TbAwsMSBUy5Sq9lepW4+ZxjTSG275gCZMJ0
D6yYqTwvaPQJTyrqg1Fb7f5faEDn6lOp+FzjAR84CEqUBjBkV/OqBVlAK0STmZU0
bCTLxc/RHsvu+EJqcZGcsh1kpXwUFW4j5PA+46ndj7IPe6sBFCqG73sfF/SY4peC
82uXzYA3hPNkcI/p1RQDgs/MwIqRnn6+Kz7ZZ1LrB1XYAMbGpak5MiKUDfGXlwu1
St5493i468ReN7pP8XcUIAMEDbE48KepRAJ3BsNBp4x27Z75LTkZFFzAi92LFLNU
cdL3rPfK0NwydmsRBH+sXwn9Pu9KHse10PpourETNvRV1FJSoIwMX0Gnygz1w+vv
y+/qbOCKbcxyu/YRzqBjpmCFMKa9czEPs1/kaH6DsvTjBb1u6uk1x+b4wQtt5v0N
IYZlCa5u8nojJnTO10ef3eyep3M0oQkbEDl/Di2zCNq34rpDNvJfTqnWyXGbxMC6
sxCrFFaM+8/nfXhrDHi+5q05ObhNOcutPbjV2b7NffxSLxPxmCe+IrsknkBDfINK
hNYiyrHptOr0/SAu9htpNiO/SvXpR4ejaFY22vjRMaQuay99hqJy3DalbdAca1T1
FmOsFVr6wr8Po7RZVBYsWozvcRxdksbnVGq09L5nx99xwIIeMSxbYNdHrj/8CF39
OWo1K6avXCtf1stxnfUzvQsxv3B2OJtuP81v+VItLVrAi1j0fHgwn3uFw523UCww
glM2woVnmkID3zsGwBc75SuXWyq28EbisiAq2kE0RvRx/9SQ+lZVn34jJh8jbW8m
tH84Z1qassBIQqJ7g1e7QpfcBXtpbIUu3py6Z1LzWYPNLGHkRXbD/mJwxdhSeuMN
ZwHksWbQT9Py2q9Qlj+QRHXyb4A5pLd5B22Uev7nAk4sW1Eyj2HnRsnWZDh44zAt
Hw/MvO8lbbCa2eRYv3X1LHNYVhv3YaevKIKut5AnX6Xa1kKox61uWLQ89hlXKxoc
vgQvjutMrLXQ8qwMPAjVCANvN7YVRkguJh7hrJVvZ5CcH54H7AWw0crJw4OQw5Mm
ucVoIBqi2DxSfFKw81FobZ6Ri4TKsLWPF+5WCvR5KZ/FW/R1WfM5oW/+w4+T1gj8
hI9FPjRlEV9xqOp70knXC7JF3KjgbDtc546aMuFEbdXh/ouCdjgaIHUSOaUhC458
dUF+t02Lbnz4mFZInusje8g7IXjqxp8f0NvKWxNPFEwgFr0O0yBKZ0l1slCvbfDZ
BLnf2TVaaMztLimHG8NohwM4eH+mokJfNNgjJOdwGMIxVbfc/aVuLtxqA8qII4+u
ZWDanH2znMb8rI+Hahkhlsou6hukfywXEn4qgaTD6LIm0JQAPIDJk4jz55MIipmB
OZtG8eDCle/MSfIJsxn7pwENQA0adZk8Y9PGP9lJT3NV6erSvZ03a7nanWl4IVTv
jlnkK5x0gXOu8Bkqgbn7x0Bg1vdDgukkDU/igGdiore2AnIfpI1vC25WpOMXlKKn
Yb89I3I46f1zvvM1/WesOScgAMrrDZIP2xHTz6Ksoe2Z+dzziC9a4vvCjZxQCi2H
YwMOkgoVgugEtqAsPMbKwwCOTHwAfo9Fhl6kBaK3w4AYVsehSz1gN1XTPFqAJHpp
Xi1xKC9cq4zMo/LDXNshF6789msLgcNnF/mvLG9hozInkhS6n4ztJ2OdM+ADsdbO
FdLCrYnxuf4FAF4WCRlc7Qatg43iQGFqmKFikZJbLKrdYKXqci5V2SKzoESd9U/F
p8icIcdkpMr14GXBX29ksVV8Nknm6gcF/DJf/b4FfhFdngAZzBbB+KoiOJCNvPVr
zuhaSdm5q22L8+5GQkqJj6fSUkOD3+9eG0fVIdB8tiVDiKGd8PZQU74gsblidN6x
Jzqw8lTi2EH69oICHPy84CgIn3/Qo94F3Tgimxq1kUaBLg75kmb4eKsGDIh9t422
sDDhWd7LkIXgrDE3IbMxV8DQW10xS3zk7Fe9jisSFawNDNsdP2+wNJWEINUts1f4
sWTAGHZxOjb9zqbYjZCw9tMsszgbGhdCcd35enUYwbgcoUQcrYbi/Suupxv+MubQ
5vmlrWttcWDZs10O2YQAF0WTC6Wk5LawuRQgKL6p+0GyeXFPh9QkpMGRWrnkxczb
pSi78gmHL6D/nE4ss5Yg+yAD4k9LS9d8mRM03wTgbAbTfdywQsBLo++0/oZ0uwLd
41HT+vpTlvowiaIosZ41iMLTftGLr3QVbPUyA1oOu8PeccNVb8UXcWPiBzfgbHKK
uOX4mKXg1w9TZ2Ejuzf/X0G65OxcKkjOFbsMiHh0ZJ61dCMZ3WziWKzx4Z0ivjC4
jiWf1KKJxY8M+/7bw+lhHmQYkwtxl2AO24leHn8VDM7WhZDcsCZ7reFn9piNvdyG
TBbM+IMFcojIb8ev/1DPLLkWdzm2Dk6ADROQQ/eUyEk3nvJyGg/IHXA6E4D3wYKg
SZjWjWnEG82xMLJK6O7I4Wk+FGOWby4wdp6RzY7JVOA5f+ddJ+bwmo9W5Kr4KSg5
cN7usF27CmmddlVhcDQWXilT5ZefY5ZSyuGnlvUrS0XoH5VjfT/t2D65A1usZGRI
4wfecuHD7PaoLT/+II3tFrPBaCxIwKYG4By2p20PNc0f3lxO2BZaWQlzaFPGNdTh
uSUqjwG2+kmwgXs7baK9+ckdFanQwc0n7So6+T3f8Jl4lAlar6T3aF/3dNPSb1yc
YRkIzYda9/IHfxjvYcVCsKjQiWs75RJW96Ldky+Jf9AwHD9DLEJcKUr/rButCS6s
F73RzToJSBokpVCJCcfg17WIALdVEsM4T1+xaRk8qAZGIpNUk5B/bH0ZR4lzypgd
lRvxIrRrXZhOIE+hnptZrdbXU71k8eHmdGlwip4mhvisIrCs8DoeJ0sB7ecp7qEG
qgbdst10mmFDuWq0d0+VfSQ9V/EFyTlVhLd54XUXRrVvfshNrffdbjjyGJMl8B5G
sP/lndWHeeiPfhHcWSCMgmWNFVW3/owAqEcNnT5k14CBakOKMuxI1dJidetGb1dB
Ds+QaFM+3XbfGUOIv3aGoxuCtvlXa4GXg8H40d5R9SwONiWenUqDQAIGwJJv2Igg
uZeA5Emi4DUdyAo7T33qICQGqElDtFKSmHFqdxfvaHIvmrkwVMkaoFBQEZbXonXV
6fuw6pdWBNLvVLVKREnGQ01Pnwotq5HTjxosRPGHJ0bFYqcwlfVMNpsmVIqv4X0I
ivig7PL8shfuGv5qy5aJVTr/k9qWXNmNANHxgdAV0SVvkSMfh9hOG2FqCS4M+rQZ
jvOjQ42YDGVZeH6UW0ous9pTk+Z9OVDyT1EfTtuPStm67WcVzinP8nYHURONfJiy
VY/44wayfy6SAKpg3SvXdFdKkjEwHx2GNUZE8RLI9UNut5vZ06h45mXFWyze4l/s
ISzpZIjmqvA+zSwh9MKF+HfHNOgiANcYX3jETttM19eoXejorcC5kNObdwoxL+1M
PFkDA+ayV0zupRH+R7WWRIeAEfWxylEikZHhxIhD6FarBABeZoGEkjzt6D2tJZzM
byj4LYkifaRDhKVnL++ReZgLmq0TYuYyS8B/m5M7oQJv5RkLurrl81puPKiPJLxf
ihEsogMUkSvjcWp5902HZJVR76q0eoSlB3F+4whFFlccb6K7sUBuS7tnVH6Bx4mg
pHWWO+jHdSx1WflD7BEFW/XPJqHjet9bt7A3Dx0TBerPe+qJsv6PQWzQz4pgQ17B
NXKatwcZd79ilXve2S+sYPTO0UQHbK45W2fUo9tGXME6Yo9S8Jm5KC90K9wsvdDl
o5fVNDmI1HD+GjaLlD4JewDeTVxE/cyuIxaaUocBsabEvuu/i/8YOVwfEdryJM9D
a3xUKzo+PChKTrBWrKSjxiEsf8lS4/D60NjrXoP8R77F3Yrvb50YZ2T2yuVS2pP8
OgdkqRZWdx5a5xnCRJUuhqjyaDQFzizzVBAiogAMOrMNsaPc8YR/d0Nmz3zo33I4
uZg17YRxyOUYcX/R4oyVo/qvrm0UsEnp3uiMtAg9nH92gVQNz02Asy9VzmAKgFys
F1WTsamWCNKE3JYG2l3P+S46efjbPoXwxLX93fINLSNSwf2YkIdh/6LUSBzfVhAH
pOtITTipE++FA0fF8l4GS8i12dx+jnBGeqLsfV/+PAxALpM+tFICz5JYz7Tf336+
CeOclLbUUhJvYWynxugVuU+RMON/q+CDVq9voNMcDHKmpUX3imZR5/Pf2kmFY85k
uRij9wyZah8ouqCTfq74ZZlKE6LHVgGW5b3bVIzSAnC6uEjY+Scc9XRjhXxo2zB2
K6APk61u4VANeH7nXbhnaZ8acDu93wfc1JIURHUWlBwcD09jymI5jYVGH6qNpYN7
+4qEN3o/iktzXQ2NgzTkCvzBRTHOqy7Gc0ESC+iKGtTlbNa3nYryPnBREDJMlcGX
cZDIN4nx+1ijH6Trlz1HD1CxKdzLkQF5ixcUxIa6Tb/x2u2O6YViJRokY87Sa3xz
sDkfvDhUzrImSiFeNoexynnSnZyOzMJVSL6ETWUyyEr5fUUpb1lT/nMbCRHk7I1a
jtxWh4rvLWBmPHYiUBMmUp3AMLqjcU4RLLL5irAhFBw7YKFP6QHmv5dg9PkjR6to
yXk/BiR0XSG24hvdqMeSknP67+8sMRjYJcgVBskEIZuE9nFipBGAZEfDj6qRSQwq
YS4tF6qA3Nonad9D9EC0VPCu1xRuw8MpnTA0wr+0FOnyiVxHv+dqpkT8b7aY6Rf9
koW2vGzQqO26wSN/CVqK0XwOY+0FjR296HGirYVhUP47w6KFp2pYUG/CWEAlG5L7
P7PhaykrtuOF7cZtFv2S9Uu5y5pagABqGaDu8bYq7A5DZreN9d8H+2JN/VZbdPjM
4cQVmslr4lzFv8IWkgxjEBHIGD4vg8Ke0FzpCZb9mjiXONRa5U3/lCiQSo79DRMj
Vs5d3vc3iiH41OmupTCuCPOMeTVBx6y+xt4+wDmZ3IysO+bmbVmWM6hy89e+WODZ
ib6cul5DdJctD88r6xzQ0Dd7ab4W1u4p8o4u6Ix8+yYb3TfxVt3evEUv/l2fojj6
OmTXo9kyhD+Knnz6+QYyRvrF2atcVTqsk58E8i2DvkbUkbDMHqCQYo2RC1zSdK3M
CFBUdDIRrELucz4Ipy9Tr9Noq1lYfVnMAsy6VAGR7PhZSnpw7ZLioxEk346bDJ3J
aQDQaB4pP3lXlsfSPFy8B1b9CY2kviPeOoIpOork/0uAmmSzvZ6KRdYvad9GDAQ2
1gjHzwon0GLCGHYjU9jQeXFW1pHUhjhlvlhrstevXADRB2LpZIHaAwLTMCk+MSMc
+Ai8Pqj1ovW04G51VXtekV35oidj/e9/VpMRsNj4r4rtWF+/ov8ipg5lvaaSzwgr
cz6xR1gxJ97b87nNfuFQR2hMTOv5egU3kyANO3SYKTGE2fg2bvuhFexEtVOwGXgU
iI494LHVMBVo7veFz+mH42WnW/hZyUdFTz3iaCtz9l9yy/LGzDmiFBZdgMtNHNDc
UFU8tiMFO9vfphc7yM0zVE5NxCiXuVcK8Bos5nTahZR0ySihhi6C7KJwUY7R3hE7
ZvfEi96mp0CyyIiasSgjOkdNhpDD2qdYIq+nxl7+GYeLlwin0vjNfBfjnz+eOsy6
Y670VDqBRFBigM1pv2BaHiWKutd33zFb9Wmw9udybvo8pknjrsAqzUT9wGIipTE9
cCM/ivLV5Sgstu4jEd8Sqqgx+76Fzy/ZZFRFg58FQrrOOb8RD2P0AqdZMTcNUrlX
FQcO5xNnOhj6fVr20YVmPDZUulQ7oy/HjNfAw+LvAXYb0n0sOYrtYxNHew83OZWG
3gx2rq1bwPrckhSnToaFBWPFP9/1s3kSrdY3KzOScJKX7J9TonT/kl0SSu2SyvLw
93ZxrYYofVeej5xcfWyCN/97S39834M3qhXZ/RTA8dd8jj08G6SHnwKXjQC0ZsOP
1wdUYwsIV42BOt3qO9hYCAYeNxxM2rV3rRpFMVFlJm6PmnZ2pGzO/M91AlI44SWO
amIO6d9hTq+yusJq2M917RBcfchl9U/7LInEApU4OGBQT3OI77ZJODymb3f8qLcy
taDc2z7tWGg0Ttihi5EHHd4EJXmwgBW+6Qbd2P9WF+d1gjtTxyTChDrfv1VW9QEX
41AUiyVtjH4pTewHa/KIn4AVeJoEB3u51W46CJRyu6glxQdwYSOvYZnBbFEUF6lV
ghMTXmnZee3ZZB3V5LD0pjbqeCyWoP4nroI7EoqlyR5sOKcyYb6rdCqMoFyW8Nvn
H4d0LITVfPiQV0cQtcTzzINyCM6ecLgQ4DqmKZ+JdnR3exCcavbgexkp/ozHMI8I
JaFBVgRedJoH5Wo+WzZ+5pH2aoKvEFQcK1Y2cgU0jU0XC8Mu9rj24UijCqk4F185
rV5P0sMmnA0ZMaJJS2DENj9JJUdY/8S6nWbok/Y/Gg83ZfRi6os9e6OxI0UuHMwE
A8UBZnIaZa8Uaxt3Vk10O6awVLF6EPP2Vc+md9bF6n5YbO1eaItx5HOZjdKtrvVK
l54m0ucqqEwxX96pHP/4/eY6l3TM0DMQFkExc3OHvJuDRFKKLgqt6ujU1tNTaMvD
yaPH+RlvrhD2rdcmHKjp9c9cIBmtDWPERYToY52s512Iyj22V9c+JvvZMgD0nrh9
Z9DpsoscH6NkidtKtDbjG07GQwELDuoaBd/Ae+q8O/8HWrTqWs6ZDhknt2eR/4Ze
R5M4RX9Lsn2rvQzhprUokzbmqPomnN6wLtqJ41Tb9oJP6VJAdAAUxr39iMzwtlEq
wPdt0OVJRm4hVKabG2KqBrKVoY7RA36h6qhWVGNQbFdt4hxq4id7EsRjJXSb8DMf
ZY6iOUgOHLFOrheX4J3jMPrz4JhiefMzHiitqRE3mz3UGWL0Rhfc05Z80ilopwPp
6L6EVjKcmiguabfMhVzwrnxRWSxpsY9Wxr3/uD15WxQi3o7icahy419ULbQhMqi5
xYxfvQ7VliTMGSxVCkYKROP7MYODqqAJsZUj3pZn47bboWYWqqCC+4D8oTmqWO6m
kZjMBKpAA/pn9lPP+ldF2gpRQw7IrpTlEowcbwq0NTeZAhL1wwJHX7Q2+0iiAM3/
nQ1FtOZGszlshnISgCoYiv9RAlE/bdR6N3MnOWSODrmwUqAWCuLpUnI76habN4/7
vJRW0tK05BPz/DPXLCOuoU4LSsw3Oubbiv5tioQsAp6FhL7eCS6JWQSPK/zU+1nr
Iv3Zt16wWEr9x5LoGXmRORV9G3JNAnns1bccwf82w7MgprOt0004CFBQ+KIx7ltd
ZlWytIy52cSZ28SkzZRiynaJDAHS2CCFt5TfCPNdMvMNpxF3Dw6WFOwO0O0MAlpw
RdNBv8vWlIXk4A3GNgy8xSXjYiWXR6eLEMcaYkdcFVPLT05KlfEwxujoSR8xi1ZO
SbFEaKq+c3xpkOKv+47xfMnA1B0hpBoprcIobv+Qi+1NeFXIafMKfk+mKFNOQhSt
cRAVW+cYu0VzgFY8Pm5Xj1KkvgJYxilYZ1fVonT2BXIUtUhS40tVyTgVcTp1HXxz
bbjfQFHpPfVA3qD5MSr84pWzAJV+cRgqvmbGX+7ar7h6QhTI6IZ2x//CQH8sR6Uf
NLy5jPSXbZ2j8b3kgslQpr7QmlsHfOQSSrWnoMgFmJwuPaXIsozz5Vcxqcka+RY8
sKTqpTO9Qn2Y/bKbdhsM6QmFbeMNv3M8PEMdCb1haajQ88Hh791B2nkoH0kdyprQ
7e9cph47/fAaQhyBGc+qgp7qp6ntPF/vhxM/QPDk21tznnOOzsL7qpumSMIQd9Rp
9EKm0R505ZmF6cPVpm+DZoJHiAAOa0V77GSIJyAQq0hmniHtPtGyn6X/h/Bz9K+L
LlLYAMkwe9mYROZHgfrAG7R3PgCwfnVFICjeTbs4N9qscqv5W7cgLeV0Sq9uCsMo
JFwPzVTjFKwNWG1Ht6kTibg5NY0cCjqxiKbTJlJxJNof3bqGu7c9DV7uaVvNdlDU
yksa/X/r4dCzIcctwz+r/2+QiZzCu9WwEm2IFmdUgJBbQ5q9tuTaehA8L5pUswY5
RTiuTLhdpaHzFVF7aISVGTRkivIG8b4JOmn9OcWePgvm6dgOVbCz0qHJVU84QHiI
NtR5Qzrlp34VNZUcHuw3qOeIGUJ3hZgGMqw1F1GcpvU5XoC197+AzR13UVgYidWN
svT/+Z8+0m6OqlBz8YhmS/6bYCmaq6NyJVogJYV+ipImucHkTVMZXBaR8f9o2DfT
jJVI1DUqXb9DidsSIXBCqURgNVzfxDlwH0BzE5qjTMsjRX7zu6UyeE+ljBSIvdO9
6cMz1+UT71JbPWQI8KukawuxT2iPcps6r4OBZSrKmzomtdxtGpppsSP+K3ahvRWt
Mny3WdHS+L1sTefHE/9kDddvC6ld5ToY0Oejj1MEIe9PORPRxq0Ki7NLtyNS48E6
mqpb/4qhIij4BPRoBcvjzgXw/ttG5+pAgVtWehPCnjNNfGo7bPCmhSqbrnS+1TbU
a0jrtOC2rNcba4Cb/ZlHrGBLbxoR/MHzGu8hu61okSMl6l31ZG8CtMpsbCUfiA0h
FFjMjQA+MfSK8KI42bpdigXOb6Ulg3eikAOVShQIbl4ZPzHJDCpMZTEIh01tV8Ny
Q+O0TrSxw0Q7d0G/dx9OvmEwCfjzchhmveC7pGjUhtIhShm6ODfEDJ7E1mePvDyx
yyLvgTRb6Faa/B0nYEDWdwCpgwBHy77qKHSibwLLaVRASzaAObd3hyPgHwUoMvcM
3h6SeftsGgGDcw/adUaitVPXbCt7rlfXm4/jINYOSTu2215PTQmBshn5ZAQ5Mpkz
niIE0b7qxh6EclZnvZ+Batl+axHmGMCVJx6aEQKgJpoSHnGslCDXP1auGmptU7/s
ZhTb77p2qr4efG+v9YOi2Dx8oFAr/4wAHCtEMxQ6ps1EVe8X3QYjr8q23rpywa9p
r342QlhqM/d+pBUT3zWD8+So1J3IWXN3HTtriqiD8NouqX+3nN8IPSiU8o++QF6S
U11eMa5J5GAxHh8+8T75at7DBZI1nUeL0gQMcDSs6Z5xtPmuD8gkEOC4rnqz5HST
1i0vAo/rEaBd02p6cdW4z3axEef+DPnuwcuMbbZKQD2gDAAFx6f5ac+sUffU8DKQ
mXQKY+tjSMSNZ4gbAVw8gV8BYKP/6tF6bW7edfcNwIpf4F4BBYk79XmMyM2nGzrg
WXxpAoOor1qxN2rSbNLV7mA9p2lcdssc4SOOIXdczUy4ASdgWTOXCXkYvD9Ihcuz
M3tPGgHsM+BzcDcP0pY1yGfx/le8mjd+05l6vhlPsasxl6ccXFOk8c2Fj3LdPk9g
0fWVrb0eNEeikFSN0RdEAhOqDI5DeV5tZyfqBpsaY3k5L0TeUgSorPvuryTdOXse
Qb6/TmoOErQf2kC0+dCWmaWk8G2sXldBnnjZRinFHSh+nDnEqtr7q/yLQFXwBNbP
7Y072RRK9sA5GavKyJwTqnLSC4IrMDnVfnuaWOdZZo1AG31RqnD67O+whGR3LAD+
Hqb6uFFf9VhMHz/FExAuMj+3TAEGUP8KGfOfqXad8NH6r/D9TuZ9ptXzUahW7SbN
TzIHZY+M8lWv31LxgdAXmFW2O+BMoL8dwL8eyWSuoSPgixJOnqSh95JS5nkD54d6
Da0dXzl8RcCIXbW0jpxi3WbE8l6iI2V/xT/7J8aYp3A1eMH4YAtVBPyvKNJHu1cf
q9MWvhcdrkVYtr28uz++QLcJDIUf1OJzvKbrXXTXGtM4Q+NwrEcsB/nHc+0MoCpz
+KNZk8vOFTlIJrpb+E593AGprHBMK9GhQjVDLxCN+psWkeVJU7GI1fI22TjKjnP7
tQ9kq6JeuuDH+YpM/VzdF13hjYgOWwt/wVUuaTd3Cv6m6jGL7IUZAUBupb+sYX0N
/a4AY4GTOLs9XrE/sCcSTNOxnN8sBFOJbf4BmzPwO1M8h9PCQPG35TkUWpSYhJrj
IsgEQPdCg2PeN8DQn6SifP6MfsTJ/x37bwURknw+pLXI729rqV+0mIc6XJ0Nj5Xz
76dbEQD6JQLInvkPTHVoFPKZFP7uzeUdeWRRg/v9sShyoTD700hOuPh2JWGNu+Tw
2CryQ+IGHCbqokG+UTyvTeK3dJojdurHoeWjTRnyHzumWAVtOZIuKrUncoXRzcQR
Y6U3ey6EpbPLMaTMeg7L41PljxjKAqBqgqoKelz6n7y/9jjujAW+OSwn0HjQ0sUX
lc6PblZqSndgg6S7lNXTQmwzEO0pRrgJ+jrxo2OIv1iqI0ITrCwUltIepbnrTEVk
XXTQnmBsrckqwJ6GTMNakuBqfAIpxtlc6Z395KaMDv8TVoyfijVcT2PuPZ0UvfBI
65O4NSlAJqN1tsC030U9dq4dcp/Q+X+y8LFKFUNW4H8P4Jdz35NjVFZw2arFS7nb
2u1mVOs8xAJcSM49zq7uUcKA/LS+wKusVYqjMbgFUg3ZXNdL4XVRy740Ng5KBW5m
Eo2A0L/FjRAMLLsfBadLI1/xYOlvcnQJ/8bXCBzydpsf/x4Lee4qiGHrGBeqYjzQ
g1iTo/FYZT4DPU5jYIHAbVHqK291GyuQ4O9t61LxdiLhV9EdrsCz35uFK/6O8pIk
Lrbc+0e0NCe8uoPaBD9x1KvL0fqG81fSSwuLq3HcAFxqallJoOCbzNGDT8O4Zrwz
QlXFgoU5q12BDfDqxuXBXwLKS7S5QBpyqNIIpf78ABQFvCLCktE2OqprzAU+UZaL
BENukV6vDOuBaoqFCSLX4WwStlD/MbKLlw0HB1z5SB+PrZFbfqiPlYKkdaoWMhlf
04P/RrWOOdT9R6msCa4i0acE996SMWSjXo6VJjWe8w4Q+Ft9nPOhOvh+YCj2filV
kbLMkmrYjLyBWjj525C9NVbFbqxIj072IoMLWvKVGr2SlBWep2AtIORrGCU5Q95c
6s/4BWr1o8N+B7/VrVTPVsNqFyX5TkCAFyfXCnZkuJu7ynKC9uVclk4STnfqw3G6
Sz4/uJ8Qm89lUPnPT466QGSFpQA5tgflUjNzJx0PR9SX16MJ7wI02tBQO1C/WmVj
hmxnjzVBizA5a3zCkT2V680Y9wwg2Yre6D5ZOLq7lUBYeNISEAHvbOfYtjmvJ2U6
tq2WiZOQzoRYcrUWdh0qxh3ldcwQX1bOCKEv1njmhM/+FJejb5uNUYGS6hrWOT7i
SekLbN3VHXAFV5cGrQVS872bhkReqmdgN+l7xOCsLXfAR1LmCdfM2gKVZrefWrrA
tnolWZ6L9jcfKfcNYHZ52zP7/geLg9Gw4AHXiUv778g19XlCQuXzHGWcUf74J+yz
lrd13/+dcKk9O/+4cZUAnOV7ayS5Uy9hctDgQQ9n8tQrhy6uwuCemWVtJwkQCIyq
VkU/eNyrvWKCccYGyWxjjzkAubifi6i3QE7dNhTi58eHrlto7tnrryN5WgcSdeEW
CqsF8JydhOZYXuZvoqkeShZQeppHIvFygKN8cK4B6LOlp1H1wDxFWjZ0XD4heWUs
YkcOjA+mviua5u9Aenachv0r+CpHAGzLO63uODaQpdU0ZxkwQBUgQNbX0ursQMFK
bAUCLvhdVIwdOY5ACpwERAO/gQSJxGhDcmlxQA8W+l/O47tnMcyCq8bkGwnagZXa
d+we4cSeVpZrOGgt6RY+P3U/sdl/8PA8wIBLT+S8lBSGMsYQZZOSoDHpKo7k25Lx
iOsf3J8HuWFTHil4fSXwnQSE5c7zo64b2ufaqlmEYzONsMpThsiJ5H48kM9KKzQR
T951YUZLmx9Ie1YCLohrBgnQPTKPUQCazXowwKX+pn1b3w6546gWAYY2Mi2tpfzV
b+pBvwLbWeFak0EoR0YhUFvVy8ZoB9PV01VQLvQQTMtPB6D2BeEjxYQ05CgRMiKx
j1PYmySIbcMwFGjp9KNSdKSndk4gsIvQQkxBo09l1S1ZxA6KduWA6oedHCQ20IQi
JTSxiQjDsi4TH5uTLNz+6v16gzdaXvpPrApX9J9RSeZg5pN+u2YWd/cvrupe/jvq
VhGqpC0y05A0t/0LppGJcYu9+8PuX65phtu1hu9uIjWDr8PVTKIi5x9xIPP1xxST
u1agtANiy6AWIczN7uGQa8EW1I9Y+lbpv3YF0aTm0QcEcjrIhPjb7dgJfarfC7aj
ARuowSo0wB8I7n+GSEq97AJ656/7uwAdPzhc+J3tqNZ7u23qWs3h59HdezWMunMe
bmGUBhnvss4aTYRbD2gikoXlaC3B648WBarmtSxGG+i1WtM6Bi/MGSgWR5nHnQE2
QFxTxCyKSR9sRjuU+7it5ZAFM37oKkdQCjnqYffbSHGl2DWpobmip+F26Ledsa4k
cZoVi/prrb4zbOFdXgNjeHN/2Vy4sdD9b923I8LKGe0ccoyLcfFUR87WzrN1SRph
tkbBllJoPPyBMCrR+2mhgs15x1btKkPFlow0U/mG7yFlaYNr5AuvRn640UyyKdpK
FOYMk0JYcnrGzLeAax98G8lWCUGDa3Q7dsBA4cGcEDk6jf94vvAWGdqB7pnlfrJx
75wECMgzAHkkHvi6RBsbvDnQq4HFbsrA0SLbZ67txxzEYe1pI222u1cyGNi9UxNP
mszhierRDH+L7d4WcvEyUvryDUU6CfDbx63+fGuGWdwHWn8cb4n48nMQDo2XVzf7
lkwO2M5+qsDoqlajpav30QbKHA17oWl+fhjT41hab1u3sUwQISCbj0tDJHIX+LH8
DUrC/hWr+KgElPWieLFIYHCkCYn+EtyVLJ3cnA6sKCWVKizIUwuwVuhalPd8AoeI
aG2dPPYV4upsIsj/VlCIJJOguTq5MwzdZZyLHD8jtf9+QwzudlP7IcWhj/EBkxcO
PpJjNu2SREUOfFENXABhkFVCQ+8rH2tkQ8eAPtX47C2MmkXsnUZQYOGtlgz8hI8S
DG1abxaL5QOiNevwgpbaKKx4zF/boxhdZFD/98glY7UWgXnhKijm4/cVCzjq5Bgm
u75fh6vKCC5ED6Eoc4QDi6DA3dkHtxrhNN8HWOCWK+wVAn3dJDg+TpiWznTHDaNY
ejfGBFWgMGyNO9hj4pzvcPU9ln8liEImoCj5ClFByS55aOzLmCnpyy6mIb5P24HM
KNGW3s8dgjiBoqPKnFaZESwCCmIlga4rkdXVqMYGC4klGJ//KcFRknJEsaX11fVw
i/3zLws/ah/TjMmiVOhpoxnMRjOx9uugIrHo8MHgEfjubQ4TmigNZhMsx78ZMSMO
vSTghPfSce+TlU8VFGB8KMS+nx+yq3/e8P4ZUlZ18JF2cgs6QX6ceapmaUYQd5m0
HMpByNgLaPc2PScNvIqdhUJsVf+M8rS77Ve+BpS+6PCcGycuLZDwUKbSDteE9nuf
2tuKmpIAPf41X26aouC7VxYLoW+ItLvrfutAN5Vn/eoZx4lGsnv39T5/XSu9x3KF
HIn7g22zMDraFNhq1hnQGlFns/m3zBs7LkSAMUxn3w5HJolDLpD55tq7jdkQhVnk
x82egGMACDDxz3+wVB3BskJ1iU3PtKAvXwXcsqe+GID37Yyuwpb7o8dSVj2AzUbh
c2knM+oKytV/snnltzAGWdc6bQRFQ4Shfm7MMgFNCcwyLg3koiF92weFlvVodphT
d2xqX+yQRFoBetIDUIWh1xQyCAjjrWdedfGCYoIuPXYSFxKLeQEi59UQfXcHnOCu
fnflqwbycXMZJJYlUDFskF8O4Zn/BazvesojkQdirM73SyoeIjn55gxOH5v3r2Z9
laEFunPX0C7GaWAEHQ1dC/v6MQBlaa2jLKQKEX+eV0zy7fJVoQY8CQi0cnbudIID
CP+yRjkg/IlIc0od78Yojs5tOKspoPsyY+NkPu+OoMNsQRPToUC608Y+dETNyVoA
DQHTNs5UlUntBOzFc0nQ13pYH1Fs9E0NRGFR5ZV2HCkXr7MFE3C1qBA/FtZ6Vtz+
TRymfcN/tkUqd2VNWDTPrCgq/4XmG49B8T8quefZvKejuxYoV6c6YhHCPBF6IPp6
SeuAXtsDvtJPfygrncCgNa+4mErbesRORpp16QAKxwz88gwmajh+62N1CFnhxsK2
MPx52zHubZqEZkt5cGyQGfrg2WqEBSdupLmq5ZcEXnvySHbWgpEPX5Hx91nlBidf
Z10t3svfaOv04sj0ASSVri0mAYu420CG60IguXViLpzCJ1qyCITSUf2JelhXfveu
VrrSWYEltC3bmfAyBR/zZD0ronmQxkdKCqjqSoFFJmVBgslcn9q6LZUhZzlUIQSM
Bhh6DApOjmfTnexlyMYQ/9bV8L7Dt0kqzUXr6TEoqshqj3KJCwfy+ILrBXxTCN36
QhYnbnrTxOVVAXJprMfturafg/O5B4BwU9O8B3F6bM4GYPp2LHLU7XSOI3PT4jHs
AE4hi0wsyEB3lRB2OBzqLY27hV1iJa8urDFhR46WSSXKBip+mSTVCRrEJft/wXa1
86z93QaWj8Vbn1PQU+zMU1r6HLl422C6cCLFSkUumeXtyJeEw2AGYal+AE7te7mn
hxl5ESRxGtHVhTB5EBXgZh7VmTF6xkSvidvw75KyGL6Eiatt/4ORB1qftVrnbnfo
E5r97usa0mSRNO75WyJDtHv1GfC1lW1hErrAnrbG/WkqZ/2a3OG7GuP08KNUVRpe
bhhQ3q2aLQ5TDAC+UbiKntNOPSIJJLV/x/Zk2qqUZGQ2vgpz8W6CO+hBcgfW/MDk
gX3CqBDLDvT7Z9ORs6rX31KHV7dnPUNYwTagxzy7wKl/BH+6lvlTGTcFTf3ZI4uT
g18AaYFD1M/NIC1XZLkROoDOoVGQ2Tvoo86lMcNPs8nQ2xS4U+vt4QMFWkPJt27e
PnSzjH8jAZmvKt6BqQQHmvzcQGPXsWl1pIa05mdOxeJ6DBVhXL0/zfQzMPdTM4tx
MMlvwQNATCUt+Plb0J9EWBo2NQZviguODJx98aRB5cyG6MdqM9rGk4GzKfHSo+wg
mYwaNrtGk5/xt4L8YqJF5N8Otu3Xlnv1d32/Qsfs3VQCTBm6K7mfDTgiqyWlEz21
/QNdvJZNggFvASY/iXWa2ATbp1YGzKflQsM6V1J4zN6PA9ap3Za5gCKzZaqh231B
RNrxYJj/VBYh362NKJb8VS6XcxI1YnGqoVXjvZoIXflad355dnEmPMozDgTXYyLs
/KfLJJ2uynTY5Cw/IBxiu9w1uda0sKviMqadbXQpvouTdjDUkUCYVDw3c75iE1zh
TPqx3snbr1oPdoSoUuSga0xwQcd7bFNawpM1+GpOmreWa0tHCPG36XeOFiU3/KgP
EdrzHE9TYbLQxiEk+QNKhHaKbqN7O4P2jG2qM3DGVOYCpZbnn37NTRI1MIMm16VC
j/BRq8HaYc/30sWK8uCb8R6q/O1K1XBy5j//Gx192UDn2wq9pgIRt97PBW6JhbTz
HSsxcFdNdE53j8GKLmYn4f8MGPor2e67YGdn3b4B+L71r8jAXuuXWet7z0mdLwwJ
yQfVDHVihzcBzjBRWk++CIBIcfqESbX4KXMD/eRIPL9RmNG9Tok2CzF7sWBKvcwk
bj/rOfa+HNiAk8kAJg+cGfY9nuAEiNsKOrkUiOLHnffSy7C5SmVoSb1E/472qdEt
23OBuGNwE7+UzTYSjMKcl/5vhuqkvYGqtHEGMXIzw+XQOqndDo1S56a2R8XlUmdS
tSO3O6WYSW+QkZe1Gxdtg2SZZfvxUvoc37YEBokTuFTTf3QSUcc8aInq/eUaUH4s
uRgtYgng8n1P9A5c/ltd3SHmMeR7pUxOtT21SwtUgygpQ2FK+Vw1YaEPhESD3QGo
CxfvaQgj0qpytoAzcmgJHG5EzgDIdKai15EQAgvl6+KlzXVR/2J9VpKqgKauMZ2C
WL0IYb4+MbF6werm8A7OB5ItCri6dhDm3giWXudmkQMBMChvMov4JNE4jy9VvXXb
NG3dDq+/kpUBAfpgJhSEDKzMkO6K9hyP/Qh57YYL6q9gBcex/PX3fs6N87U7dtbU
xYdtORAbh4IE1I5gYCTZek12Ak4r2JcqOLw/AJsLgx8OJGs8G9iGtPeqLRUS3rRC
vpXrAFS7HadhcaMCkWUXzpPtECEPl+LgDV7NUnh48g60zRllScmouoLOlnBhjBSa
MuSXWkJ/nevtsZf5+ujw6q6eKLZdfn0usSU4MHo2+o4WoSWwYvUzZRW4HQpKRsBM
Lys+uW//hikzvTU8UbR8fkE6AyLCLV0MLpJJv8YnBxB2tBKhDxGNIFr1Uw38F2Uq
E3m52yCWDuoV73n8sgOZxLSNcVrDzUsEJyG5joPEf1SB585tf64QLPJLcnRNSbKQ
JxaePvfiMUa98/UOxInDiYK7URLyZ9Qy8LqMzzNJPb56uBQin7CpL7jSt7RMnsJv
OGxq+RlWqWB6pxKKIDNuGDFU79NSPWlKCAyH2ohussaTAxZrpdeP6FHGcczJ3dap
c6HPWTLbtMirDa1LPuU65sVFvUFgEFubKh7DpbfnrWwTGncNG4IMEhrAgxmtuvyI
buQToetteehsQGsIbw7fWl6cxOGxp4fprQuijy7oSL5sm8DinHmZHKdtLuuwOtkc
0mU9PbcqpUQSy1iiwc1qasZim8Y2XMmeBN4xmM6ripQBIbRKd2LFtgGEKx1dxr2i
lqT5st8bVU8V2OP/VZ/jfHO/DkFH429nBEp0v8N/GXlufSIpvpa0srSNSyf0Zxif
+4uAOkE54aT2GmLcGpk8VPKbuQv4T0SPyAuTiBk8azyiCQSDWGkAf7l9x7Y6in0p
VOcytUCy3CEgOvLvDPMewq6KgIexAT6x5BxL2Hc6PUW2kCWCnyIXMHUjWejMJj22
1Iorh0o96jH3VavfF7F2SLjuWb81/XoAbAnIuSfH2f2e786+ykVGWihrK0LP2iB9
pUOrn5MOqdRiztlYEF5iCVuWiwhm8mVqBp4Dq/rE4tcPm4Hk711HCld9pCkceRDK
kgaWDZtKmQInDD9Zl0ptv7yefN59TjxocBREkWCMVA1n3GAwC9t9YVU4jj24gF48
NOueE3y6ri24SY9uVEyjwD/1c5X4/UFebAdol4IuBpXf1FwB5mc6+m9EtsbixJqS
RmUBiWIsKzn6flBshUFn2r8lpXJX3Nxz5v1LnSKHdf2ir7YFhowoTmqjrnQ2DcO4
JeJSA857ltPHjxX5x8C5FYYpZCIoEmmVITMV7LJnzVKxRWHnDrxEvU3+CRR4NOgw
TS4ltnKNTxAvKgkMKUn+EKLeGiWmeWy5bo+37CXy1X0aTNKpcZtxt9TckasRMa0c
/EiCFknzFueBYhS9+LHL4um8TSEPzRHTU9T2o7tuGUnQ9cfG6mLkOp/ZJHc0egDf
89O6RVC0wB6m4FGXWsGf2glzjWMHNVO/uzQKzuSvYEhZLlz16ptIRHKmP2llMkVN
6yFO2bs+/NMnRzxbYuL2bbq1gZjOcZ5eneb4gHvzRsfkKViPhahBvVCsZ1JyL4ve
EZosV6BC7rC/EC1WBKWoDAs+Mk+nf/0EmMDfkYR9432gXzXKdQPViugZXwdAMwLe
j1JSP81dlmBiYNXS7Z4qjFyZS4SrIAFkL291mX97MUI4j51Ffdc+71LwoldqyDaU
kgLug+9cDng8ATRKgI/l784J4JF+LfZ3TzgqFpxqXTLFjaaUA+B0PW9at8A1zqed
kv2UNuO0+a74e9Ka27bTTX+GjYUpkEGaa9HTgDnftwOepBAI6QrncZuo3J6VToOe
9qeR8TnfJrSLeSPAJBVJWUmbKr62lXSkCERg97qBoZeNSMc84B8CybS9C9LZ/Q1z
ILpWRp9FLDcKVk2tSNlZ0S5TvUsEGq0G8G4TF1K09KZfDyJcOksNkx3GWp6x07uO
hjUtw3vV6OVtu4xLttKA/EJ/5AjEOulOmLXPh7Nz/jdKMBx/SA3+Kik4sKkWhWQ7
fFvnjXXBeyhdCH1D+HhjTuVdBL8z/H5TiYgKKJXwGu9X8LSc2q0Rm4n/dqOJkttm
OekVUI1VAkenVwf7EWiiMvf0s91Uoj1p7iLrVyB4E4KtSJjyhhFfLsQRHnvbqHI8
U2Lyqe1foeU3veDvGSOUIppw0WA1AYFbTf2jaQynGz1YnGjq3I0T0CvLCA362Woi
aMIJN0ZuHz0Cq5itO5jWoSvfnnUxf1FcpeO4Qdy4gfAgSEBek6Cr4m9V+nRyexJ2
uXAIse3Ib+7m8Ss6zOUtrGzV4DsV///MxqbEOtCznsXJt+vDNbrwO7Q+5m5uXz0k
Ftfo9Oym+4johbRyDG6BeeUlRsnfFxbmDrdX+d/E9M4/bk1FGl0rh7sYLpMG3HLD
kIxCBYgRhUEdXgadWi2wwoR1FSRr+8+oGHwE+jkxKuflK8VES99JHTrohFPpmZaR
mC5TBUOvhXB9h9Ct0d9xnN9xXlKDU2S6nREsUNUuNeo+NqkI0kzj+FiZ5DjYi3Xg
Y+mSKD/jhI+g54OsuFmtzkAURDjBzNMoVZPeov43Ur0gTuA5PKm+ZfqdoB5a2WPA
vGNuGRq19Hr0cyEZaM+3kA7eRw8ZG52pcgXCFh9ufi/Cn5le4rugqCKwXMVZylEu
auUkj4kmji0gYEmqN3wrMvKsYMxlZn3RP+IDPSJ24qbdtn6h97E9TO9C5ujeaeLV
QXJ8qB/T1ph7I6vvCtVG7+x2Ug9hgkZADKkrnM+vDmd0SOUsJJPwutkhqMjBni5P
cBVwjAPGCf/F9XWKJZ9ib0cCAbfR1dI8ns9E5E40TSBO9hYujAlkicFv/1NoS739
i9Nrka95sDYQGC1aAlsx6z375W/EVMq4ygnQXzl74hdlHreBlOM50iApD8gSp97g
HZnoq26yq7Lb5piCpfmtTfn5K+Cuoynn5pfDEQDmr9PWRHHZ49iTw2wtK/9b0Ai3
gj8nNMCld1wbn5Z8ZgWroB1qol4Fkh653E0DBYj0HpKyaXQWMGqNnBiREfgJ1kUU
08pcwHKP8y3cJZUwBxmnTSj2WBdZ6ZEClc4VP6FsCzqaR/hTUTrlVK8DIGmbE00H
QGI+IBAZMHy0E0goIWhFVPevs0m05/tOXeP64wtyv0w7dfoiH+nbqm2anL2HNlrt
MNtdg4suoVdREkNGlhMlNXSmCjG7AlvPv1BGXitKnP52/E5eGj2eSSr6eBTv5yvr
VKGAWiVcWVZIQMBUek+7uVHqpMpXuo6ktNmqakatV/mD38eY6iJmDIpbuFFNhMJJ
JFfl7wKw7sbkjRhOHdqo6OwhcLI5QQ6wRrunukMRuPk+zmzKXfOQoxX4O0hc64PS
z1LIYQ9h68LW5nwA6YLqk9H9hvEfPxYKYOIg8Lh/1yE3jbr3pU8faHXF9ZrYsjOx
sKFoAzWdzw6kgp4Y6U2o80Bk45MUNFEclAsznvLn7+dj8TtVx/V2naU4Y37B2yfs
zk7ac+tqyrZoug0SGjNJGMCccJ34sShpt2xhblALQlUk0sdnTnGNMHrZzwrhDdtJ
6qNG3YINjQfqEqP+zsTywLj3S6rCA0hzEMItuEcm37WOka6LpyZRWW93tjeR29eU
TyhAJq76E4XJ/cp43Nsg9WHTB8BZGKaiG8QT3KEmroiX0gauCudy+J87CDcfZSqF
Zh2SfX3DNE8YUQsijEECnL8sR3EI/Aofm+o+4DkgeqvPqgVaYyNaEO9j6MrGcwDp
5FhefmRUd/4AvM4lQTw729+fWlsnwYEn1OgUOJgdsxrFJc1lWNFXXHUQQeG/GASE
fDDk96n6tvaIm/T21QEdCZs0bOfApG2DefxxyoizZMaoDvngGM/pdhPUpRVcXCL9
uotdY/fPbs+HC9nBkZ7e+DYO/jOGFXwDko+wjBtF7JyxJcy8B5yuWSezdYGgtVA6
0Ho+XgJut/dYRGwvvYw1dZ4WsyqdUipstoeUCoJhA0BbeVoiPF0amYCm/CdqBzX4
GvpmV0XgXhep/kBoQQVKoLF1wjPbv/gNfMEth3tp8ORFCSfjCB+/J9l0ju8FHNHO
aghdg1NTkS9QER8IV29riMPDjkcGZS5Je75fMpeYt+EK1HwKIS8n7nPTkID6tuQk
wdf9+itBcUNJUe4JNoFWTqazvtxU1ukMlBzcPhZmg6M9hYIe4hQxdA9oEME2uEy1
i8WpZQq3zZCUq074heQbvkVnZiJHC1rTwrAVFUImFWR/5eDfEHWEeV2u3XBN76U2
fjrnuiH9mvZhGmL9UITBPQ5p0x3fdUVG09AG6P/SeO4KWqMhZ5HQiz58NuJcb3BJ
rNg8J4AfX5/lk8m7+Y35Q1I24qR8qATbhnHHBRotJ0bsUiwrw8VugD8IgH/xqyAg
3nIqYM128NnzlElIe1rq5f9pbA26RXBO1Y9eh8azhzvFv0FZgxEKQNhRTbI/KUHH
qbxIkthFa98DCdxU4WTA1cphHpTWBkhDMrTGurj5JpJZT9nd4jTV3pI1t+XYjsg6
MKRMJS9WUjKtszM/2gJCgsc96rMBZ2VNfrG2AKCeZaQWBEj26TaRsmtM5mYHarlY
zECGLxovT6e+Yl0rg6/zRvnWMMxoTry2W+/OBOuvCv9+84a8z8N/Ju3UveGhRT0/
L6F8Qp1FdAXzpYGMBO9y7iwB/JAKWjLrtVk2gjerzBeIzmRXCLMKJp8ei2QGROP9
QHruPE50Qu1IYIXSi/5MT7j0N+cdL8STkpHFZk9U4+l1/uQMqiSql4Su52xQV92P
GwWdsqgqlcYee00ORwZPjXuWUMP5+Ze+Fqy8VojSzjNqEvxjhWnAOydOrc6SnUiw
LU7PQo7PmVcMpcKUFE1GkV0yPnnyjhyzbU8GIvH2xAlYvdQpLJrFQtCqaMWtDDYk
Ppkdf2AudAijdkO9Tsr1n0T9hqeU/Eczo28Bk4Y1zfKwp8UU8dEU3n14A3XNWhON
bCiUbQXO97cG60naqRl19QoWlictGkRKlCarlu4vKUB4sadUwjfsmAPgznj68Ob6
vLVJZ8nyPV3umUqc9mu5qgaJrLnNVaolfsJbg1sSZek51tfBo4oUf+MG9Ng3hhq8
fos7JNFc43Pemee9RFJ5gkWkLbShkgO2Tjua2rUyLo0vPQPA3AP04sVms75Mar4g
44Qti/9i6cbK75ZkbvBxVzeFKf7z9ScGzE3QUFdBlK0CLs03ab3f03cfBG1+u4oX
Xfc2YifRx6j52UlvdEQs13FiLP2s6ZaQlcLX3tCuguheYoPqhw7mGSVgr/WUbvIP
DaCvh/SrPZ+XZpiqGoixZGHwio1Ztq5JvORGEfVanl44v9tvzKFL4jyoDle3rFmG
HKqA6TVXLZdkFm7PQpkK4U+YBqi5n01bsA1a2NKkK5queyyEHOTk+y7q+8hOngxh
0vhI43uvt/2IB5se4oED8hkLjCWAteYUm7r9Etx4XKJHwmI/1+7YjOuajIdNuAkO
o218emaGrl/aHhyAo0r0/vw614nmPn2JEN7FTAQ/d/dQa6nljcvK9txJwkdz/lxm
Uuv/U/dH1Epin7/gYQvqIewiEHStt2WF8u9xwNbgTzZmNkl8Vtu+6sKAJJLwgSg5
G8zJP1pW1+xYziGYaexye9/sA3FpZom5HE9M2MtI7abbuUC5eblDGNNxZpXCE7df
zaOXqxQy439qt0oDo28I6v10ytBRUknivQQtAzlUJaSKsobQaPuE5HVGHnQd8S9k
q48zeWvq9QuR1Ay61bddeJxyrDXAjX461xokQIVknitnM0bM4ULZ5cYdpJiuHmj8
uXct/GhYQKRdFjTrViA3QTpWeW8oe/8i3UWtbVKmk7TkHx6JnGSTquMPx+Brpucu
pVptMmiyASJrZRmL6HoERbvfuVGh7iRgfMF+wbd/ecMZcq9UWKfd7mggMUELagcL
TuCDmruYyb+GjDCbeOjyPWMMK9Kg03fKwdpIJ2y8GE0aVqPrmnvJ/5QsFEESSv+4
4m0IQcupke3VUsP5NYlm1xydM/mGo9bVRq4YoymaDdQ5jLhVTTNTSEZwpsPxfYCA
Rah8ZaWERssI1fH8DIWfGQungggoWk/i7PJokg5ZEjdgQUXgoOTfMyRu9z9v9v6+
tk7ogYObYutFFRb+ImnCmWdUZXdKgK5dn3kG24etSkOnBbs2iYrstfRbMBx0nmtV
iGqsqbBDrKniEAep9YnlkhS1+rCpVvTx5neyy3WARiPKq6HPPXBO6dQeDZX2FRyr
prfY7HIPJae6MTNi4tUjlJQYKE4pPa2/h33nGXalH50Uh019BWL3c2g6fiUGYM4s
4XOVXFRBCOw2qp6CnNY3hnCLeQRx/O3lXSHxyq6c1AMc484+j3qR2xyHMVMwRp1Y
4roRgtTU2s7ZaBnhreaY127+C/o16xelETl9UIVZSrDG0awM1HzzFcTuv3SuwlX6
pG5j5h1RXAzrnCjQZttiFf2EgReuxyK9XZNablGnkv1/Io0zq9fR8B74qUMSIL7c
qBW4VsUbqiyFVmLbwyIuQOFEjyh8O9T8wv9yrYh3nPtsUsPO7T07s/UYBLVm/wA3
jLOPdSbZJkFdzEKWAfIhIc+lveRR+YRqBSeMOOar1ezp4h1SNgUn0eWyDX4y48UI
aZ6mWYy/ma+54NjqWIZ23ECyvpIEjbP8W5fq0TlYmXuM7G0GDIWEUD3uEq9T0LTC
xD5v+v3+eHyzPAFYc1u13bfdQ035uz6s80uCHIUI7V298z3AY0djbLv0OwySWapk
ZLWN9bl4b5DU/xbNw0fKlGs3VUhT7Mia1N0VCW6Fe00P+3anjq7AHSSPLemCeFRW
Jj6lTxfkD/A1rXeUcssrs/6dbF3iuXQvJddlHacKKB2zrxaAPXWk4jDnicAr8GYJ
+i6vNHIplMRBY6DpU9AzYisN/hXYQM4T3v+08leA1qOIU4cONQ9z6q0WDq0RCPqK
cx8aHs0Yuy5K+RaxQQ8FFgiU6OLQid7PC8NvoHQFwh1HWT0bOYJwNxXPtEOGdDhg
cSo+FL8jIaUX3+XGE/OWqEoQrXQMR/QaxOEy/XN7FYkftLz/x7MHk+kI97I4d1dd
kD9kuwlyq1nnqreO+YnvuGAueTIGwvhsAc0duq+A4TPQi2cDmYFs/Jz5bm9jUOiM
kwbq7tAtCCaVfFhaFRJGEGANhG2GCueLmGXK2xTQC72EUxLFbyZDW1uARTuFmkch
svX/wiC2oZkv0hfM0mvvfJyTNB4BDfyh3tb+ZyUJJNGix3PEt/fmeplzW3HcSOaZ
Gx/+Iy4zUvunRyieQ68RuGNjIANE2AUTs6sJGFfRf8cshvcHF2HFMia00qJu2TSn
QdbStiGelVNK6RNrLsGqr3yE/A31/YPswXePr/sEupxK5qeda74m/qsyu41A9qM6
S5iAT/F5yueAqzAY95GwfIFLNI1t+Oo1u3oH7KZ1ZOOj3ZA4R5soFedWkbKuhQZD
nedKgDIYCeY3tgJTbM1OowNuJplRbm0HggWZPqe8C1eR+FI20bLPK/h04DnrDCis
jFdEuItIHWy3eyDRK5S37HJo8cXCNX6wEdga1uXlkLNi8reye+7ZllImeic5NGJj
lU72XObK3Dpp8MPIHbzqS6418MLvl+Wq9AYWGz5480YFSJmSzgjaD5m02gwpXNLf
32myBLTGzBpuToH9W1JDCBV+pN3a2UztxLAJImGuhF8XX3rqVsZ1FotCRHGi7xyR
rB0Fx1Gio5RAUNpJWnLu+U4zRT901NOPRUOrh4H9mKS/L3BRXfZ8I1fqdQQiGJ1z
uRK6SNTLj9Are9CSJ0IR9sGXyhT8WZVrSjw2Leb+L2DHF3F7YSf45zlJb+no1I5H
ocO/0d5/2RDk7pjzvliKcIZy+yQoUMG1qbDcWsuCJPvXSblNnle+qnN4BvVZbEQV
gjCyf10gT5udUDQvwmaNzZ+2R/p0UE9w8Inn9N8DTn9iHbwbqMX95FsiHSGVVh45
sLdlLaJAazzTbxt6cu7bnYvbn0p5U0e1lRFqas/KOI7HlkKimR7D0URXy01EA+/o
kgUMSCYuQPJLvu+4W77rNlcB5+4gxckowOZYy8XStUZOvi2bSEoxLel+GdZPic/b
3FEcbONP+x++uGklVzTma/Uqdv9iGtI5AC2AVf3AI68BgNT5iJlIOln0lmHzGGvf
x3mUSvUTQndggHvR2vTpYMXAdur13r17LSVNFQ+COKnhuNOQIE/ufRxaUx6vVq9j
MYu2xLELB15JVuiUieXsIEdK0vlDHsG5i1EX1hWtXpWcfa3RWEmMe4e9/+zbHsfj
Nbe9bxvYH4ZGCcZt7Dvwb0E/qaL2D+TYTYnbQBulQ57v5t71+kL/1ei8+1Vyf7Nm
ihia76ty8UAF/n6zaK/nx2n1HJ/9bX3RiM3P9GiBELY7EOwkI2i36zy25I1LwA8G
fXupMsPd+90HmFtBk2Jwz63jTIxeQuRPL4biqgQ9h1erYtEYpVpSSjrwbJq17lWZ
6P+L/IFXpwKlGRgtaWEWuJIEljoBNeIOQvrTilUgV+STkzepNQjF9FaMW4SN8hpo
pIsNDizyMhxnds4bK/Cmy7Ut1+rJOwHGMfD4bj5GS1M9u3PmWtd6GKB/bpDLmcGF
G7tPBZocRerpQPLn2JcfKwY91fMYhht2uCStPK2T1KPL/Nhwi9z+rA2bawPqJyiu
ueb8JRokGeu2QjJb9qS5uSIEf5TX+GQ5UbGQHo+qv6yfexz9hVXVt+xapxrRskw7
rxMENS0Pk3fvcFRm5zFpGnoa+qndA/pAsyo15CYwbXNWbGtrY0oBKZG99r6a6Xkx
W21bnh9i7YUX7zFLvVKEhRgobgErLi6zm5jSVyIGH5dRocbqd8PDOr8aM1m+gaB+
L40zwn6HGr5QGlKmyL54T0YEiS2z1bQOfhskdfypFb8fRTaNc5gpKUUsr2o5LPqX
7efIvh7WW23sSqMiTp12TnGrmZpNLH14abXmUw+jpPE0CK48syoioGtAKlMZexzG
u6xFnNLlE/cdEF3tcM1n+vifF11+2OKukFvNcS4f88wPwV6tCklbqGGPXnp/AAV9
fc0gOyvp3KYWA/Ur1SbYUScekNhbGeIRAKwaOxUr1fAWi8T994eGBNK8bIPU0Pn/
tk3jSBGp9NI3ZIzQ7d1z/arZLMqc3+Red/mc2/obS/G5aLeLezYeAdlLsozWzjdZ
O0re9QkXwCFHUsWo7chZakx44/SMz17UF8eFN2x9Ba4KlZsxu5OUEl/LhsTLzID+
wU2s4xHKNfWQ0znFSW+GGLIf0Wkcy3QXeGtb0VrY2Z2rLKVM8a8TC/sUApeFWU/W
yDQQTEhCSNw+O0uP4RnTkFe/R+3ZwovZXCcTP7fA5kE5fBjIhyvku4N6tXg3GQmT
qN37k0bLYOSwWbpP3xNTHm9NNYWtdVZEqjmvlyQZ7Kphd/Z2qkeYylPvZ3WgBPks
g9/0FOPnb8PgLkveqfgZSvMh/OqAOnQL4DTWAk6U4XJRjbvEd7/Ib5M/H5nwCVJP
+Ds/1fRLSPXXKKrhbVIGV2yb8DXcSGfwpf077WddSXmocwJyS0QZxkstPAo3UKk2
hxBv+afw5jsKfAoq8ObIVDwqyRNysagZ3hArTDHg37eYtA/m71t+Tjp4j+reK3u9
9qLVcIeEmFmPIpUUn8FraNXjQWyP0vPrTGIpDKrPIwe3sjclVAeUV5lIXIfsGqTy
ltLgpKBJNRZAgI2lWvkOo3nsuyByiJy7dMLZEM/PsNV/LTNi3MYUaXR04nciAPfu
SHaaIkg5flqrpDo7sLOKci9sthpquvCRsPYyP3FpJrJg+Do7Okacr/26SXmuIAhb
hQVABRysXyB4qOn4E09kJALOlsLV/TEYS0ASxFWgjuEryzkrlZQTb8JTCtNURuJd
UEfB53M5QmxRU82jkukXs2if6PD3QbL6McreZ2V43dN7OVFYj2nie2HNceU2seAi
+V0IvK6/oYnas+IJeBAh00mEK642oq4E9UI2mfUGeQwfqYC8njQ0BirIx0fZcWt2
N2JuOzzqeway7hPqFxir+leB/auyMfoFLdeHCP+b6Jr8Dc4n4m/Cda7n6l4vqizk
5/CDmz4sZRckLfBoUhD16o+6Bnefagxw1W74/8mmgVbLl5PHbCVOU+R3w3d4X+9B
zbfvnzPUQIHbu/SiMUtWmEqxYCdMbD4M87THjfTLEzcym+3B3unaFPhj2JmVGcUV
q0g2sRpr4W3+48y+H5rE7TRjbTKYBAe7HhzSIf6hPK9gkKtgf2NEIaZmCJIJ3GWP
2BLZHsPsBD3fijE4lrt51b6U/jeAGReO9xmlkrNumoIP7KYzck7LN8XWg8OC9QTE
tyZaeHKEGZVffXxDk5PW71LI9/4V4f0UiG9Lfaxm8QX6rFUVazpDw314ptv5dbeX
0QwOhb1wj8Xwgu2FXlvdhpIFP+pZ2BFfol7767nvdQu1dmGnVpaofRU+Y1hF/Goa
DpuyXhX0dxRxHJpRNdRVlo6lLr9UmJC//BopQgz3X+EJO3gkriyKYBYpfuI7B6He
orRCoDCHqKLIKMb4gMWGSIgjqQE+kCsJIlOGpE51gDstCiiG++ZyReZoftJv/FEf
iFg9uitCbvvFTj+bMbws85d9qE9GZQ5h0mSTSbqMBHSRLsF6tC4tjCHIf5rNnlNg
W1kHmw4kqcxeObuG0F7dyR2LogUkHJp5084JGviNbgRwnKblcb/xHtUeo1oJ98kK
ha/frB9jCSqeD75QoPErXHaJ5DhFwiJIkSgT1ZVHo+uy2OYsaCI9xPUMrLnFZMSY
iX3Lt4JOMAUc7H2DMRE3p+DFBrhPuFb52Iwbxy1s2Od996sdb/jPheGkaXuIYpzg
t7fV40ZqDOKvc+gN6muzsQn08hu1j68SpfaiXDRrRFJsEC+1CQYwdDDcYfRF81R7
jGbuZXafJlewOuxRnF4ThVZx3Q+0ZpjymGLJx8PsMBT0CB+6IJVAwP0nGcJ1IvSA
beUclkrKCo2ItzZFKCy4GH3aQQ61FYaLRXf10cofK7yDH1fs2jUH+3Z35fecGRe3
/bwcFDKKReKrl+q8uhtLbUZaeEqF3GP8RNAlvKAxoEhm5rG7TK1rRYhYEhpJThOG
NiPowxXYZsBez74d8D+o9A05vQHdoNG38hPUxbRrzZ5gaBTv8K4mTitw2pexlTOC
Z1jK7kLF/8Gs+CMi7jEWImDMFDsvuu4MB0RPz+pEWW/Ci7uDR5dfN4D58FR/tNB5
eWXCSAH5nxIrv92UKAQEMz5cJdYOStJGhDD3O5gXqtMoOilCiVmr/G2Uvi9pQKPN
NCwRpxW2RoEpFznXfMOTU89APkrR+/Kuq0+YdOGLOLj7yiDBKqLby+CSFVegc5v9
fkytYXCSYxZqruyZLQ+yEozT5CYdYopy4X3DAuCvlyeDOADyC6zsUfUP1ATXwN7u
KmOTywu5yPLxiDHXdsF64DAXqpJ0fn/5evNKydYZA330ojk44H+zp5q5oRl6nR6i
jFf4nSTet5bs3mIHVCas+K5WicCSBOXeJfDKBrO2fxRmj/644JFE5dsJbcvMU9sl
2W14Z+ZX5VTduhVpFB56nQ+CB14UkbSLs5mYXEmiaQ9OlhRNYxGGSGgCPpK61t4p
bGQtOw6NjgnUr9oMrtuKDn36R6gYXh2ZE5QXhbqZ++7MEJ8CRuzUuaMLi4HMLJZm
3iJXyfNSxYP7f7d/BAiWtQs76zqv9aTeHYaqN8ngGoKfpmj0L2m21VD6nbOXcXbH
2WKUc34SXATBjGpcALfp8GEM1rRu2T2j2UnOV+H57zWugdhHD/7K/r2c7hNVUrBH
HG0gPc1tEcl0yeU/WkUW4/6EemR9Ctm7x2EIo8EzwxE1QHZBquFBXDlC69IYTTtV
ktEttjtynWUf+CxbhUKKEdHJR4pbqgtGIiVd2/FjZawE1N/sSPhhcMntG5zSD1sd
OjbIUaL0yzlf4c8qnTXYRbqXHWU8mvoDnj7itm/+w8O3Cj3vU/deASUl5M6ms/He
b4jWO2EvKQ0MX8JUBf/feacJ76qjZjqzqsYzrhEUb6Ps3Z5Ms0qOVKe3I2xvZpsP
2oIZLNnJR+oGKB74wlt0WXDaIlBSA29hTrFiORDIT9WWh7C3th0r2XVJxiDfRM1H
9mKHTWHfqtdLTUXdScqXSJhs2axSw2shvS41rPcQYFI/85WyeYkkDS8TE7Nr5zfy
jiz8IHJj5Jb38gRm9GOWZ3jKvf7Co02OZa5+qh+6nqHk6i80tbPt/qjG1h9NU8Lh
hMGszupVN9gWmuh9IwRvJgB1wBxxLQjlds7qI3N58oMb5lwQosN+gJ+86ZHCpsGp
ReuMMvJCBCCI/xwprraXBp5CpdY2ISqOPfMCUviG2lbOl3bIilpFqnB2qV9k/T+d
tKMMVabiH38FmlqeQlVjrEL8jscAEzpMas4+BUo21CS+q1Zf3X5HaI4kBZ+dIp+o
Dpvc0QXkkA5/e5e54yl6dfQ72CdVN/NSEQPpxH/SqtGGILNhp84+sTV77vUFCSho
Lsf2p323PXhWm4eqDnVd9pgpMsV0SQVyefrXMtXNYQuebxCILzgUyGRCTMXF97nI
TA4j4QMAtqDLyBdEj6mYaD53ngHb4xG6Vo8tsV7YGO8qsXU0oMEzBbDPnhDPS/Y3
QKUKCRjG+8Z4tgG7DJo0O2Fwyi5qtonx6wY+SYOKcOiMLZ6nkCezP0nX1UWkcd8f
ZJ5yyXX9PqYuw7VsDNTry0rXzE1of14gtewQJI5xS/iUWMisT6sc14QT0csehd6P
bxhuysGnrK2hjRmkpGIbg6nWQ452PVX/ztxDFF5S9WkMLt7LlBAhRe/eXo83RNwy
b74dWLVAwgcytu59u7YWabSFkWaGxyv2ZxNtdC9skf6ZMGRcS0MXrQ7s0Ki5gAS4
xtJTAU/WQUZBhZ35eowFhGlwot48KDxq1nnckokmWKP3dY9Nwg0ddObia6Du7e5u
fKAfFcK+l7/pApT9E0ZkxIhQ6Pk3BSNYvArjPqTr1BFJMR0VO8u5XzQvvU7BZ48Z
XmrDJoYXm+OJUu2xzsZZ+bxDfrhKVBXaOyctgwUlUF4MpGrmpB4O3sS57j78i5aI
ZqFzEocCFH7LQiWpqCA9YUQPFeP3Sr8obUrFMlKuEJ6OLUA+0s+ghONkMp4+AI+X
H/gmsEZ4gb6i1GhOvnuHdmeat8d6xY01fXC4+RPR3C/Kb+Rm70iciTbu6WoIURBc
ClBN2uZKjqNYwM0CfPBLOMwurDqMsqFl7JSgEtBAx2/Bwame4M1h8pGH0BLXujy9
JH/NQGQZn0appykNyaTY83Tm2MGQdgz3YZ+cjNg87u2zXZUvIE2rnR9hW9/4bbz1
CJ8u2KIJe/uQG4sFHMyfDsKRjF61Q3p1AdLO1wfAjfZ078YBgnuJIAJi4GMm8o4I
TTmP4D42XycBDL7dPlX1EhXe5pd2hKbDyWrVv3NW62AbUZXzlwhATdytupMwbNp+
2VjSuF21UP5suSTalht6nan1QhbMeWQx204qtWKxx/zWI25laWhmpRRiUtp0h0TQ
xjDXfTErkNMKrQ8X5QvjrtUc4HALX8RoKRtusTTswCRODJ+pTTHwGoCtez0SI6KQ
WFbFqhiHPPmtK1g0Amnwj05mBtNVEVKHH3rfoh7c5JHp/2afMxgCIPY36hOKSrfD
JffwetGsnQfZt+xhGcOuZHcKk+lvVqMlY3zU4ZfpELceeorMtO2m0xIZwM0T5fzz
K4k87XLMCGyQ8xC50HbqZXcy5koF2bqHFAGkbFMc/Hdk0Q5GXEM3oxMW4jbI8bEF
4zt2YQyIrosFXRk45vNk98sbQibCYsSsg6K5xGlHkRgaDeuvQIcMqOrtcnJrqwvm
S7ozRIkbdJ/cZds82+ssaurdZzrlH1fN1cLguQdGiZsNDAC3fbT3ep4aYi/a16Wk
FYCH9k9aRhdESYTdeaaPjdtnQ50rmmjDasuyvp+1EniQpa2Tbe3WDLix/UOaaTii
yDom7dkbruyxxrVcSNn7K1JX5g4WtxxmkDu+jvfR5pPfxJiOOq+w3ZoggAhr3zDd
ZdcESFYaIzZmd1UTrse2KnXmFFyqrOpHclGIvOCFxEEzeLu4nNBHSqy5VU8Wdk/7
/2N1bHs3xOQR1PGn42WYWkQ9S8M/l1nhSsDQGeQi/1GaZQxlphor4FjijXnQQb+6
cJ6cRBDx3z/uxMND8vI/TD1DKu6zaIwuOEB3ectpPyvWInn4ytAfS0+19UuwkCq9
A+DnrfLAvnrA9RbchMRuWo1WPzrvPexMq6cQ7MNMDeWtvDcZgKoFFVUJ4ixonk+m
ctreogMOhw6ffOsRUQqteJxljAJs39thayOwT03FoB7zExQIQPx31rHj7cZfx+xt
156FBVb5VwlN5umpbkCjbf7ssXVLKt7gOzKZ5HAs13Z9Njqcn90op79oID0Ys4F4
OIEtWCUs1QFUCUgh/H8pk+a8Ig3GJhLOMArl48r+i++xle+HPDjA75Y76rurRKKl
+Ew71W2QYYAj/HpvZDaIwm0gfy3oKFvDJn7VE3OmnE5RoH1blChIxyb9pgieLm9O
Xs9SALoMbWwJoxin5KGB0QfDsmj4dLpHFiPPfGPbV7eRgOF4q+Qji3148OJ8dPDI
rCEEfT/R0mAwDgAzMN2cFm3O57Ee820MSyjeN5e/3J3p7rqdiGqNWadJUXi3EjtN
g73/KR4FSZv1W5Aj743meEhQEn9qHT0v9XRJuHA8U/Np6UJ0Ql8m4wiP0kOVwPUW
p7m3QTthMForwQWQtP80wY1C/V/YpzFyVLJ9o1e6qzwB7NZnxdA0rytB4VWi34uO
Uhf4xA6V1x24p7XofSxFcpJWsNjQUC+CCVD1Rq9CtNq2hc2u+ayWXBfAN0pv0j/m
TIuJutx+czBWJtlWzWZa3aOQlw8mu490gXm7o75uDDQpJQ/TwMqJu3x7vGsqmCLg
JsCKgLYlI7CUvRgrJLoXXS/vV+8YySXe59myvCoGfGJaIwiXGKO4O/TbMqi7oorM
teCQK4R5oAhmzSgga0lQCWKjuj38vh1KKEQXbiWWb4dlajm+a/5XYslV9vl87R6t
tK04N3PWqvf+aMEPd/nneVeNvgOH4mzWbcf/C0InBMR2Zd1zBeZ5JwP57NCCuoMo
G4cGmICdUv9SZlhHqi3g3D5It/+fLI4trPA6e0BvQ+SEtFkpgbd+0Ih4qbqLwO/g
/n7OsYFkWIKPGNFzoMyeUeeQQ/7kBnD/53DsGPV/3oyL2y3fVkfRRp+tKJRivUNo
jL/6C9lajb1lE0bh7rozmUqchHqACgRDJgbcgAirkneC5L0PWh9O8JP1gAE2Jc5a
D8LX1m0cg6lH9r21YJ5PATokO187E41FdWf2RY8JOGKfJD0uiN1bUv2keaH6C4YD
dvEyV/GpcHU263m9zSylT4Ofemw355bNpB3Jk+DURDE73eSpC+hIr3Syr18mR19n
1Iz9DnLiPSjTXp2erQqduuLoV6KG+j8R4sW6pOr2Yy0pLA3f3l4QujCml3QaGFVU
B/GZfCKGp4I17rK8nloG7Ie87ZWG1ngHsHFo6CDXlQY2/VKI1eiPvCDzbKSBSuFS
nyWdKVYgmxiyv0RunLizvyI8fcs0nhTV+nijAe+ZoloxsuFc8Aud8gJ4JuqXpBan
BYlnH91XjHsz5IuyL1aV2E8XJ8GGCP3z/g0wf1/HeK9/Azrs/PJLeCLHcBnAjspd
y3NOqQZ34kdI3g7E24Cslck1FS/2l6NzIYTTM2Yy4/vg/CE2QpfBlQu5hxZwu0Jg
eagtwDQODEx4xjBSo+fNsI1+TzukYDGOPnfmZpAitUcc1cMplEa/umG/COO8V5fi
zH6EUOEOpKFsyuXwTOf2IKr68iBGEgEASIvtllxE1Me7RoTdEmgilkHIOWumb3zL
WDPMs3FvcQHrD4dOhxN66Jt4tnyTcoC6rHX3RHH87JyZBtPqykInF+q5lin/7e5s
GiVu57RrOvtAvWyzM7cnC8t/NJ88cpWDLMveiOK/upPFoqaGjxuU3EDYVWTCnQBa
zwRz98jfsK4OZJ0DB4tRWYWYTJhNyrhRTLdBAR/GX9jfQost3oCKe5JDJpioBPAG
rPSqCruHuiLGxq2QellRHxaS9nfN1TaIpYeit1nEdLWLEeCGVZl9oTRxYk3holjg
MOC6BERyQnTPok+sFL6GLzB6XkqCPF40nuf3ZhZPT17fAL/yONf+KtChVuKmmn+M
PUTcfAkBkXkz9/wqGQRkUFjGKd8KvuY4mdO4uBVi8WAdAn1NwBoLdyEAWQAo1Ck3
Dc0CSiMFE7DnDPsGRNaMO9GKcD1QoK58qHCMcm77KMqysaBy4/Mm6XaIfrRR19Zr
uUE9qQq+CLM2rK0SiGKqKrp3zZVBH7k+3gsWWsPhGuTtsm3dtBrE+4p4d573ZLri
ItM3Y0NQdhSuI0yDjYmZvkjn2fgGZvqu7J15qmEMUFHJIhTYd2PuxQ3AK/Txvzdu
EhLlS7TNtEhw3UGz2s54MfBTk3xzRJX84sSfgE/ti5dLFVym/4YrZxrm8VQfgVI1
ClKHlIMuRJ7qTsMf6Pb+H9PySIugVJ+KBU/Rhu0A+OkCWH0iuvlCIzmtW2HWwZgG
MuJEH6QgrtDK5Zhz/f0MGDcjIYUj4RsWqc7ew50nGB9A+8ma1RNOjPUA26F8zFZD
UFfl2A1qgxzEEG++yfLrLXa4EGE43NO8tmUm22DKRYjinmNUy6GPHiFqusCr+0X0
01ThqJ6KtdZT7HDuQqDmS+wtFtA5kW+lIreEhC+nXGa/lhOizZr1lSaYcsM0BzJQ
VU9FvrtF3MZ1jT61JTZCYaYIsO5i7yS4ijuoqVGKQgBDsgeW8qfaOUXfwdQSj6dl
59WmUiVI8LAL5oGwG4syN4j2M5Jo76ktcP6HAoH23F6NLcaZRLtmgjqT5F1UODOu
uDwLKf0ABay43wgvdTF4h/NpRvl3e3q/iqn80AXrtI+UEeKzVE6yK2y2Tq1VgN7E
rIA4LsufJYA0F/b5ni2zlio9I4zttb/D4esc3V20fwGqau3RQSgD271PHy0noaiq
DWv6etgpQ5enkXbsF1qRKkZMxVjQfL1xdCKad/7fXMUl5AWVSfrz6t6djC0m+WNf
CEQlTAVEix/WJ3Ka0aP93aSpWXOSQGTiEluYnggjt680ZNsA5F7VJyIFaXB9hAW6
bXQRjLrFQmXWO0d1KBQ1Y1Ka4js9XP5TjQHuyhTrY/1tYBYYZvr/IXxkMJiZ9XoB
wmurgvwWH8FD/GX7iGtdq3MTDnaeJKVgu8N2uluQaEL7Np6qcTr3Bix/xbogjkDG
D2pIjND0Oql05pxmkKi3b20gtD2b5pSUq6YY4E6mCvJq5A9MvdytEaNPa6O+6UZp
ldX0UhBxETSExp0/UG59axL7Gfbit9BWMDtITzePvZJQIHb/ZBzLnVY5pwWbkcqk
8qLFk31mmzA+tEPuIat4CE+swptjEKua/LlA35DoTb1dEZ2ivP7+lKz+bm2VIoS2
teYi+K/5XXaVWy2vHWUHR3oKMjrTdIQR5+atmfhq7DUrK+vsFyg18+9PMbgvi10q
3sEa6H3vq5kxFwwdKIPtdAOPIJ3mEqCEK5J4emWAcOmyvK+CDnkV5A0DyP3srXDP
9aXDsW7t/3geXe9dWm7Q+TDaEzoSBsh8sYoaTNUOul3MHIQnpkGxFDC2CHU5OinK
gQ3ArQDVeJf4w/xJEkKdOsuFA4b/r4f9SnT0rxcELK7eCQL+FuEOFp3B4TSOAKtP
xvN1I5C1j45WNEvP5wV9ASvIHjJVwQaufWr8+GXWB1eBBZ7yHlW/Av2nZmXkJbjx
BwQD9fWBVqxvARZ4c+X0gbKAoGviASyWAWozjMe1Bgvw+OQ3s/mYNs58Ei4i0G/Y
hKKRmzYiVB71i3NSJKxfpZADnuFB9T85NegV+6qOt685Hx9/HLRpwsl20xtpD0Sc
s15mF5MZwzkuFvZ4LhYRIYaFdteMXnmldeEAG5JThtga2En27C2iipm43PTP3G/z
mU5BBwfVcQ1L8TLNIpslrm2vMe68LnPHIXJfVd97iIcZgCjz6cMWvAClGwjE/I3z
21afUpzS4fmlrsHwbUQGgdCDS4EyF9NJbmMff2o/QIAQrcnimiUqMYP/FEpwEzal
qMNO8OH3x9V6lQx43udSqoIpuLGrcHANTQAKBJ5OMbkElZ0+BgfBKBhc6GYPfw8P
FMTsu+1RhDCKXv92EWbv7kwXAEqqrbkgHUs+psUIxV2qsBRY2kOc8xMxJLHvhgul
xAiWPJ/q5AtVbhKB5jaqNJjGDLyJWXaPOeHIYxkyrslom1RYV2FpglX6/FelKSUc
KH5HvIn61c5kMIcrZHSPvHyXi3IXpEcqYi0iEay89R6BIm0zqge8IFFEzF5WhliN
kjeYgwXs5WFNUJ4tn1+vnOfc2HGZ6YyDaR2v6U2vylOXTMtTvkNXf2B3Wkv5IHdv
yrp9r4dnt3EYxTtknjWFdahpUu9Sj/6Ab0L/XYck+oCxOsxqwAI4aggqYZTAgfee
sWH4SY2aheYdOS/hlvWQpvygZDnJIhaGLqQ9iTNWmDECv6N6VuCtvt3Wc7LYeblU
lLjJtOK2B3CscG9fMDZKwvYkt5xR323VhQu/USpwt1Jybs8apuEBjoJQj2tncaPt
tDYOaHRFMvjlL2KGrlTc6djdIcMdJk/xvF/SFuLiEIjBSs/WE6uaXvdDif6/N9B1
kBP0E4G4mehcfhPmlcDrATMIP1HqqjSusjRw9BZyOoiurWquqRzVVQ6e8vpK1MEJ
Hz9TOThKMjJVwLG4abj5n0JxBF+CG4jTwkWjlrIi9VLK3sdZqGZAIZPTV9r2wY/d
pTbJ+lMhakaPbaZJDs0AcDPrNUxfmwRGBDyheYd6msCoLYHFABf2t1UvBFZVskSs
low5YMa38E6PMEFENZXs3eiqAPNEVCmWC0J2OYTzrnS9nOVNJYpjzl/OE6atJhVA
4psgS7kcdLIMPOjK0AigAinuOXwC3cePdnjtH+nNY2493gfcUTTFsl8gTSIfj3x+
VBt0ish8CrlcbhsFcizXsZoGZysty8cKl8cv09s9o4asPs6sn0D18Mw23M/Vk7gb
6IlX4uEt6GFsRviBJmiuAX+dZYBc2oiZjykPJGSUY1MyVmF5qFGJ1r0Uod/14rC3
2MEF16kZ9+KEHPWa9vxqFTUb7+W46ehNd43H/PL7nBcg4TxFoc5B5mNfu40247FD
Sz4NA2Ex+0ZiKUkajU1/pC3EnpDA9J7FbcQeG3/hsi0p1YL9TyUrLjLyMnZGM/yb
h3sbIG8NHFsUHOh0iAoY6fdsA6R1mFGf8G9yJ/bkdQGNQAmMsvUdmeOM5je8z+jO
UfxloF23IY6y8D6CHMUhLgzfOiAlbM9Z+nSf0AzS3m1F0UmrKhyID3ULmrkCW2Du
cGt1GCpV+Eh6/JzelzRCYZS/I8tGIHR/EyPGGgv8xtpNHL0RWupEhKD0dJq89Eq7
TWUVL05QM28ukK72KFVIQjuLwDLi8ZLIle49cwbixjPXU6hP0icCzr9HOttusSjB
fvDeVoIsWXVcpaHr0XL/t73nhsnY0zYAmxdphk7a/frNZZ1P/p9irptDjU3LXJIs
07CTj/1A54HcwMX4zyhPiDzM+0zVF2i0HQeZHVe6k1tXx9aQPdc/kwck1Lr/HkMt
CuWx3Q2aoWoCnqiNVcZ7Fepdxl4LSYr58VJZr+MXqcMwrKNJkOyC4goITOTNLJXw
WjAMYIpCallWR7R0404JCqMK80bR0m10icgbPxpWHNS08byOj7NfXaQvmS9/wrzr
J0aw+YZYYvEj6Sj+Imy/T0kydlQ4XYUp8izid0ai7s63ZMQb+ZPhkcmXhOe9Y4pC
n+y/ejEccCYTNLd7bRtAkA9NarM1pyJTPnpup9Uv5CYV3Nz4ewNdQwE46keaJ+GW
qj+yyVafvQBivZaCO83SiMiuUoRkuRJbk0H2zAGJ693sYM4mzrgUnOb3sJVAxBa+
10LcActv2YEQ1Kv4rnfLJPZvCw2sKig+jvik3fbAlbGP4XVVoZSixAYh3lssYUHx
tF6y2ewB9gzU0WNSuzdR/ShXvyTV2dn7TOIr0a49hitoHLxCh8NeP7PcqIefFHLb
oo45aV2gB2yWrVECFJVu+bM3uAf4BOvB7O9wf0wDLIMPoU8y9PZQSoHg7Tr9V9AX
UbCQjimnLN7Dhgt/qkdOAmClFAvMHth3HnOpaE8PSLHLVkiOQV1yWqUKKoyBcAAh
x3/bxEU1UXZJMK//nDTvsqEZVNBjKHJoaj0ieNhR0yEIYMzWparbV70OMw4KEoLo
9W3hxCa8UYFp5pUsMk96SQTCsXjlr0zudyYPkpEUToZuwCK9JdvccWRtDfAD/UHo
1VFmKifPKnWchdrgYzqYvbbcCyy5/il5/T+XVrwnFTqvDwUAHGXNrX1IkTTfpk6x
zNJV61ctR6zm1wGMcu0rHFI+cI/G44sttVf9CZ0RzheEllywb+PLWm0HzMy436iO
W1gjUnrIvuOUEYqYG85TwEBtQ9eGOOUBEptPTR8OBbguZwJO36/o3lHrpifZ0Gd6
eziIwkBv3VjLzJgtLiRttdZZqGsi5vUSy6441SL7oZ05rOSBY62mBX8f4cZNEZ+A
uYhCd8fezW+cNkPnkilSTjgGoq58J59ZOuNNGaaLifmorDNoCJ5v23IjL7K7bmAl
JE8SeNmHPqiVR22Y9uxperS3mSbrB/FNZSkkGLvPyPvfjG+YsLKWy7rBfb3SbiE/
AB76Zk+AOSevqzxoTr6OU2EGuKvvIL4bFIJP0Kc3kUD55YaTwhOW+TbOvnCRNjRf
F74W9CdokCrlb+Iuc5JGAc5MUNMhPBNurP2HaSgR5cYbahOnygaKZ+Vhy87EnE7S
J8IBRczVBVLR1ca59F0swSBpOEEh0mAnSonldlcQ9U76WTK0dmfHmjJDIMdfGmsz
x8EWE54Cw4fPgnhU5aSzxWF1PsEhC09K3Lmo9j16cQepGrbQwb5AeZlLb9B+sTN+
f0py1xD1R8+ObGnVfS/3FlHuB6PLqovYIKBi5VrNjj7ffCebyUZv9WyLm42f6AlB
AEDUI+U1K2WFT7xf4JqSrVNJeBc6kjor9I4AHk0xyYXFt7EZBO4/V+DgLuyYGd6R
7D+cWDZ0cwgP/kzPc/jtDyIU4GCnkNunmbr3fA4G7ciNkq5okueVo9HaCV65UnGS
KFHxYdZSP2lVmV4sMVuPmNGMaiezGILg87bmZsWzCKCDse4eTZxWm6c8E1Hr4vvb
yEZ9vtok9Q5KnrjRfGEBV4aWuTBS+J84LnWANGKGbds51FrW75UdcnNKLiNif/iW
dqdNAemx+61oT0raTrjE7szV3ZT0PHXpGW2r+v+g3mlAV1dZ6I70BqKBSfPYntGE
GPPNbtVzbgZidmdRw+UhzI9NMjeDS+lUvBwAt5cCSBI9eZghUls5t4zELW0cMKBW
J9PbsoYlbGQWXm3XaPVRe59z+o1L2HeUWciaUNLT6Nt4o8CLa10xiVpf2sHdKBfv
lGCztL2DufxaQZbp+Dc7hDk8drbBw9hQSe/mG31l4WUxHBYHmpe37i8sfRuWFS31
9dB3UsUM/Gz/Tpu6bnlBidLIHcGBsvsWNYgCjAwGJJZHHUH+Q60uZQucHIPMR4vq
ylq66OThSTRV5G2tG+k68BjjbAwxjwKlHw3EbLgNpxY/+XsJjVhCA2P/UHCndMMX
Ksi2+Z5UFijQsaoftHwlndlGdanS2msntiLnnuN8oTkSbyAEErhgEwdhSPloS/0u
nAVg99lYfuafSjs6DUBNBoVrNV02Ao3R8SURiqbfCFz339Zxacib9xXTPio2XlV1
/gAFpPt09sAuo0m1smRyJas0yPnnxzYxW6pDw1Zk+OgarfQAumdYEZfng/3Cfeto
WMfZ52cpVsTE2bqxRdhgJNAy3XISDt2IePCD356kr4yZdqfxaM665uvnAL3V3UI4
4Sd5/X7GyjJ2I8rkrcYVH66md+5iPmpxKue6R2x5lXiSBMDJ8lbfR4Svf0JLWTxV
RrMuTSEcaFsC96h5slLG7XlC7Kxe0KLN9C77+TLZd2k0KR7WlgUAQvSqLK2qnT42
1EIkXtxNFPR5uHxPo2fRBp2iwo1GvchCczd1JtZWwUObKBIYLpdZ6R/HoS/kNBRI
wfal/m9gEwiWMpX+GE9tjclzNHx+C6JmNo5evUuC16CG/bMcN6hqmrP2FUszp+Uu
PvC4UU90bmsLAffLc+RzIcJI1xTsiRthkAQWwYFEHL/UMxUWWNccUGfCg/M4dfKe
yl8EEllhT+l9cZcJD19NPV0IPzCaH2ceYqym2ahJXdHGWWf0VgMKuE92OugGpHmZ
i8SKgsLuZMVQsInBHRelbu7Dhgh9Ew0+5C9d7tLG/4v4EQ3UJuKe2lNEpUHZqeDl
S3DoNhe2BtG/hs5/qkY9ZwPona7ZaXxYe86Y8/7iQUL7h3jQbRA0L8Jg4J8DT98T
ixqZiEji9Vlk5m8JwLEgIoELpftdgtnj7BYfsmf32eP7RNwND5I0u/6+bnkmvU5y
tl6vMm0rc5OoUeZSklv1nUCOyRcDs1WHAnvH9Hwymk+i9dn4uY/VcGR57x69G5mD
0GX/11Yvz9oJLPU8MpByrZfh2ex8c02wREeUz9hc07OwTPdvhKLbn30VaImhvxe6
J9eDe5ymBWVFe9Zmi17BA+uYeVg74UlXtk9XO5EL3+8LFNVrsIFK9APx6FVH7r7F
BQ69+bqwZ1xgBGExsn0+yFqwKukagJkikglcPK6y84+Bbsvx2W8JwgdRT4Seg5AY
ShJ2PVBgcqgtS/F3D4Gho1YJvnETPR8aocU+gw+/B0GbDF9cOYTEoPBNlcN5T7Di
e56b8bca4HZ2ULsYFHtThYPSJQeNALfDShg/GCgBCQMD+PRxjbRT8ihrdFeE6Jsx
NR4VpOIqzRuFjBZwEKCWlZu0kjdfOW99fURxYutBw8wMe2TkSJyJiiLSI6fmzsc5
fqFO/X4Ebd6BFzmEazpiMdJaORfjzQQ+Pa0oBwm0LUqdmsPiwkee8BHxQqkeR1O3
Tfw/FGI1QGBH0t9F38fB5ZgY2QXdr/5Ne+rOBOmlXouG95NJm3d/EuoxnNrPKoMS
OMNjk053BzTaZzfp9mQlljWlsDnz1JctVjIEZIWBqqt/XufsAzUBeNZx7qkfTyaK
2aCvsUXtacx10YNpzigBj0HvctoWe/mlovw+B14Owf/KtJ3jMR/tJZoZtezPHLGi
YPyR68jxos4vIEI9lbsikyyNAOtQUHHnIQ8FpkzKhf66SWniLwxTCyPo1MxhIiJ/
lCvNX2JyQajDJnuRz7lXtX+rQHaT0gGNKVP/CcmLw+xPBg5fQYZHr6+G+fdGtMGp
yiRGaRDLusYs1e3bkF71PlmvTntIXjgDanihzv9WJfMtvNrUfnCzw153pFpCp66n
5PizeNEdIZvcVIzMMGpkGdAz7/xwyO4k8q6eCCGg1ujl+gbh2PAvKZTv3D1+z+Fl
bWVy02GQ0JwN0IBI0ZwLrUSdBF36jnc8Gj4APTnK6vxcHva2RQHTkFuOk40L2MjT
TF2FIGpXh0lRDrSE5iZmuctFAM2MVOhqhpWZulveAwChJR8BACxiRvREgGmZ3bsj
3F+nzqLtLyXS0voEzBpF6owfUjllMcW/r73kXtMpjs+ziEJ4+tcGiyCGTvxZxpm9
vcT4mySk6q5mQAehqsmoHxwLe+Gn0+o+gdQdKqAFkqRzp2Lgugz17NtcgdZRnl51
7JjC6vLVPwPCyu3ukej99B5Dpp8N1TBjt+taGafFVlb8B4+7O3nhBOKSxX1Q+pa6
F3a6Qr0Dhi190nvaOE7ir1klzAl9T7W55jhkmQWanJpqI9T9eYLJjRh9+RVe3j/7
utlFUBf88IWhYTnl1orBk9Kg9pw9QylJgzKy9ZmIeZB/7/ZZcxjQOzkcXHLtv4bc
88DfhSxwgoQTLt9cLoeug47F7DiQ92LnHRHb2hnCLLMMo9a6jssyTwW+lE+0Dtee
umvImAJXxFcxbWZA7vSfqrrxi7f0OW3JCcym+hYrWyaIau5Thed/8bTJD7LemPCp
C87lRlmUx4ktw3I3/ZZiSV0s/t8A1bhVAIkVreOd9QtAiQr0LCOxRYXIIfpydcKX
G+suYzIYLc0z+wiDlLwfI63jH/2XnBqcqTndSW6nu5Y17pbMwQiHgfrY5S0JRDvg
qj1W1pbbtsFlvWoiKA6Su/MQvNzFcYzf7v3FUnKS2d8nFka8l8oqbiMcNOj+1pN0
qE0dp5b2QL5TzDxTrhssuuMpWTxXeWE4BWaEyyn6YEkKvcebIqEfAFWplttvA7jq
QsuajfMleztqxBT/6NZb+c2JNztPXTeH6kgBe3Zg8nnshIITflqwz8fnY1n2YAud
sZmu+qFB76W2ZLpUBEtvbuN0qbQczUr0e+OTnqNiMqs+/U3BwJR6gAAyxtbM4gRO
mSaYcbDpwNo7Po6FWKaQFBgQjoXmRjsgRHEJ41f4a9kVG+uKKYSK4JVGx80ev2Gz
APWR9JcDzqwrQ6YqvBg/Jz3G8TyntgRArFvU2HDG7bkqinZSC0KR6NgBrFKTms2T
ZvSNq1U760fu0nWzxHpfWxTdOTXbIPtfCWIs3iMjzFUG+/kIVVk05faRGuvw6gQq
myeC4d9HPdkt5p2DuuRRSY9Nuq9LaZ5oD22m4thuuu+AOni45MTLB90dZsYd6Mwg
CSeI9wbAypdtpDtdyBYkbCToDCfOc5aitixc0fnIrCxJjbNWQLKB1P4+jFoTT3Jg
G3QsokHxlaEP9no/UPvywD4ISayxrqvt0ffyvwWpXHcRvk7DvocBh9RhHrAO96mf
VXE6mEJVQLZ1UTNQwT27BvQxn6bX/i5xCVQ8S6wU0VKj6BWmbM5vAivINaQ9YzUh
1uNXy/VuAVG6SBDzj+asSKaEkv3+GL+OcwHUfExtUUCoSo6XscuJPhZGv9Nc6HE9
B88ZhxoVSwWSaPYE8azf3EvT6LNas0rFYsyhoDZYhZ5LpO+nh16RQJiUs3cPUEN9
7Mxtuycdv7F5Qee5Ereghny7gGK1eO+2USKxZytt0dm8nZ+CQlUEu+/SFM85vmuC
8LvDf8TApAWtRFJga/7BrXEQ2Ps2EhfU9+3aZZXKAPUikLWN9nax4hu6ZmRbrqYj
G/TKLSF5WkWG1+3+eKXPHAM/ZL2lVg6AqGuT/balN6h1U+ffnNgLiNuG1PpiU1cH
1UjoAThZw90fwigtp0/YKoZixHZ+Cm1lQaScdzir+uDXtBdAczB10MOfxYYQXwtU
zlUPkmXrJdcLDcKQmxKl6/lwyMAQ3f+ibyg+TbrjNa1opE9hRdtltHBVkxp+IAue
R31jRrrw/xvkgqeLTkgE8q5gUyiK8f6TjBEk3iZCp0Jx1d96O7xsPXEv/YE9cM9+
cqrjF9KO5FXsDgh0+7o4tlTi+GPoNd9bBL2Y+wmGhCLKH6ZxWWlDAELwXJ2QDR7U
l4VdGR5HBN7jseBSXbq+O+mnZHB1ALmQ/UMIVms2qyRAw8XUPK2CupPXao/nRw+f
063SO+3TJKE6eLjGWOzJjBh9cRg4XKJqq6UHxTTXiL61ODYC8LEGvxZWooz6e7hG
iHjWEk8+v5rOfdbaPUA6+cOU5kHJl1VgCCaaCIJ+0dcwr7fxGUg7OzYou3KRH2/X
F40slFoSA43iDeq49Vp+dRLarlyByr57Fu0LpnZDzjU6m5CKgR1F1OOSjmdvuBpD
COyQ19YWXlhlV4RIkzX74aPUwipt5fb4GmLQALiPVIcVnhMTwwq2GXzW316rHOUK
uwzOWEP/+0TAfiqUGjpIzq6/DfGAtnbJdrOt8qhUVjTBKyz16rz008W6IOCQeFuj
9ZXqxUPJCrjmc83MdYz8SSqMALNof6RYAGG7joWNgA46cF6woHTxvroamFLo8KyF
hcrKi76EkW6syx8Z3LzQ6PRoPUUDKj7TtOpkW1kOBTAey8wi9pOM7xhDgv1UriA1
BG7Vcv2n08IAb+P+uxKeNWGS8xrcCbRCQNW3qkAU4M3Q72ZjcZ1qJUggY5/Quee1
S/aY4cr9SET9z+smXQftfrhIdWGfOe5p3UMz/3+uI4k6tYPwMZzi/nl5lh065Ec5
+gP2CBeQaJoqzRdgs942zzCV+G4k3rJ54g0ELKCjX7gei463cLfyy1ohBy0xuRTh
ehx8HwaiKDVG+ffkSRUzp9Z/T5imHJhX7yLq+k4xkDTudyQsFV39Ll8ekSOaiQ77
AfQMmFw0fuxdrGj8Xl6qnDTivQc3BMxEE0i3NiHacUElOXmr6vhwrOjI4/Ybe5a2
vKwubiY6SKHDWlnUw0iRwUeQA6e7FSzW35CPpDIp72FYpb9UJFG8lNZst+KIbMaA
9vxp+MY2vXi9P33EXWpl+4cqiSWMdcnHeLyIzGQk2JOqgWWX+uVdsO1jJUfEoblj
LBFXPiynWJy1EQrqqx50FpyTbiRXk5x+Xk7mOgP0OqlgMWNEcRIYWWWS+sZvGFwz
Z7HgJJDtEUrb6WrEE6M5zLLLDckmru8OnQ15J12afG+WMJEAIMfaLzTMpt7hrA9T
aFHFZeP86/hR7fvujRWDMxPSyC+z/KZRIkVMzuPZtvlh8fD8D2kcwVyZfIibBz82
kb7vW3QyTOgo42EnDxGexZFzSJf54cS4s5NSa/GmJLyLW0vkHcyh0ZcF4k297wUW
RoT6/I5en+mYTEHBtajRzEm+doILWKb5a3ANb0NKud56HeiGL+4FFPYah3lpIB27
t9b9HAxeGAkTgKHi+WIwWwOmVAygxpCV8CKY4GSC/LJRYgKxjmHafSskX5domAHI
gTbedH7l4mjVnVoty1h/KWP3YlpA9KkwiQhKk4gd445SE3RMyk1ugFiZjG2ifP7j
qyWqPfWAyF7LJSBwbQjFrT4yNEaqT7dGtv7PoOi3G5QUF7g6q+vDa5WdzquJyNU1
GjLwv2rFrKzqdNn+wXpB+NzlQqMizIreqwKi3B8bkGjcf8msvPIWAKtwvf99jALm
2avfiMyCrB3eYpk8nBrnSbO9k4PxvW5zgRT+AedBWBZWF/9fqsAX32mzwSsYsvs3
ZS6p5zJ15vLgXQ2fgwcp7LkLUohu/zJmjLxtLB2Y0wrmeER44qmuSlibSq6E548V
0jRIN6IreDsMPmMz57Ua9PS3HxjqfmXZf94PsmtET29mmDp848iTCKNWPd1vowax
dnllCHdfC+W45ngul21JRRzgjNn0IFObJYlhhD3jDjlI9D3DFn+v8wg2vIcQyx5/
9RxCXCMhhmLoLqoYyreVvfRgMqklELaHoaMwhfTAeU9Pa+/ABqAmU/YPwcjHivqq
kAiISGbu3W/m2ynKkz+B2uK9okHY35VKxgCR1ewniLQm43z4lu0Z75wentrIQkbN
O2C8egOxiWQd9e04hk6kr8H/Y6o1sQB7libuue7152ALvsmczkCd1D4BKbIHF2fZ
7pUtq9eG71Y3KPV3bZxv34+ItgqGtws8YCXvVrMi8hJUn8UKXL7tWMRWW1TiJy/b
09LDPa1vFUHxjNjSaWTfT9e3RbQ5NLHVVl7q552PuValrt6RGR+HUoUHWhgy8nWM
/mAwhIOkudHAMEhj/Z4kAYpaBHDhzf9JN3o/kyUuFFgZj0gFOIT+scY/RYnGJQJL
VTGhe7PXRKbdGkJ5amuutL5zajy6TEJbIUojNd0iBZegzSOIDjp+KMcWYcnRYZb9
LRkdMWQAFI6yy8ZtcLSm6IiXx6FU/oy8vYcBhmvEe9h94FfBVKO9qtc5PLOhQP1w
j/6SGLPSThCwVmdhvP0816MIy/6q0M365vZhVvjLBL4+dheoP4S1J1QWC8xb8fzL
XujmecCjI7L/lNI/ffiBmdi/KSDyylgVqvITfW4d/RsSw0UHbwlLqouwzJ0qonug
9cTX1wMpttfskmx2n7LpaOg0M7MPxaXhrRPOOLBWKm2LLIVGfB+JaTSEyCMtmvm4
asuLP9fvIlwqOSQfr6o8tcPEBFv5fm36FPuhqY9+TeKuNCJganbsfrQsRwAGj3NM
MsZudRgH2ivjh8clhLTwUrJ84uudneuFRvJ0PlD1bMDA2lhTHyfcddi+WcxlAdFb
IQ38pAQ1ZVK5KM5Fc3/snq59faS7WYfsmg4STtFTPWm0asN8lR/GIp7RqD1uYmSo
CvC2ltKlBtgGJMb9VHBO0cgmDMjEBK5uTjup2b1GhtjrgZtqgvAsSAqu/O0zLB60
A2bz0IrQ7pTW6Y6Q8WEroc6SHipG2WxPSIpbXprs5HcS6DXyOPfrNhcu+OiWu18y
OFDH4ttLGI3oqRMwYaeOUWOiopuUSfZDA/X6uAhJzWAVj6ITaS9WgVbuRHEbgPZB
PAq3gpoEHItZsAS4Io5ILinL71qTCuhxq8FvyKZIq5Ohf0fZOFuOKpbFWPF03/4Z
XJY44uMSDVWev4tMlU8vADkc30yL/YcO/zNvsMm45sPtca1QIF5Tgvumrn51bZ0k
8L/AIQzUX8sZxC1Bn7z23n7h0yOMRv0edAAPxfvaNFdcAyYHP6veYFFvY1Vov5Gn
IijLvuQV74bnaDLzVTJZepjEqHR+3mDnHiOP2GRNHOFeBBLonTxsnoKj+1atEINq
9QgJcwQdOf1vqAAj0YD9h7FQPA/gSUxAI5Y+lyF9CMBOK4rzmm5mN1y/lniG+j0g
SmmyOnJu9yCf+fJgjvaBopcPkwYo0mNOLOHK42oWlOMPEM44eGXZJy1YLrpaF+Qn
YErDJTuIrxqR7Fkrl7J8OVhsU6QiURzqyGPU0tU0KeYjd2kwlwsN2a6iU8uOk/k3
xxLb6Xvkqswzkstt4YxSOQuKUfdEAW+AHtVdybXKMmTDQtXi8pFagsDIpQ1Musip
Tzu0oBxLZlc9pNVYWZb3+fcK8fI+9smos/U7LBE5Ku9G2HOHkZLBnk9ULvQxEHY7
DBvRoi+heu5nEJgk50lVzkXppEWWusrCXp/Bcy+uctWEzdm7RdnsDHIylSpum9F5
d9cJtHfFuhdMn0Nqfqz5nUb84GByV7SdnoZuC/GQBPYLVGu433AKJpkpCrTc7KIM
2JIGfojdSwwY/5SLcIq4Nj/rnnGOM83bySSseSlzBuPDQ1KOnNJdWFe8nlCN7qk0
8tbyD/wYmzWfFi8BzU+Smw+BRothaI3SZwExqOc7Dm6k3XGFyTenQ1cgqL3F7eWk
pPqDeXOXdsetPedQSWnb0TeOXQPwNmGzotx6c9KADTjRVolzjN8oB1hT4cKBcg5x
TmOiU5F6ihNaw+8jlEOtWUv5S2MDeLXY4rH1cZqHbUGokVn6AA1paVQ4aHxWtWXF
bAbC4wG+kCIf/VCZ920t6VnajQE16RQWGf6xzKJBCSrkcQ/ZA75Njg5U29OQ7+uY
RLEa30waoQjpK88lIg802jlLvL/vKzwjd3l91jnzuEC4iArXO5WuA5+b8JhmS9dz
VC1SYbuVrRPjOZtrEGAbNtMlwzrvmU/Fjz0uvvo/CpCPt0ShibBVisBPD3Q8/wHB
hvqy2O2JyBNnDvtSqoPCz+O5t4osyRkB14ILUaXHN0W0IJO/NbqnzX7vGTGBvYU7
tqemoXkl2n1wpKi4hqJBavycixIAt51mQxqOjxCD1kYtWUsi6ewiR1UE36luZqln
Oiuw4+6/WfXqdEZWvHTBlJB81xwxPiCTirFxo8t404qdWXHHNcbH4Q0GBV/nJcHG
N4KG2OtEykI7uXTNep2iFG5hCwCxObsDmJwP/FXvPiH2DPdTM+kA4xwcqDJxNq6Z
T3Gq6RG8ZYq6bjzpgrjue8lUYX12fk2MEqliRWUHNWkB6pAnUy4wNK0j1jNw1RN5
YeJUEt1I9Hz4AibdY4fxFFD109DjDKMu9XqDcki3okqEG/Mr3gx6FV8ANLYx3LSW
3V4RbdOvACsPJVTFUHR2+2UG7bxiVyhmaiSSleez5elkwgDHE+roT8QzIktjdZI2
t2XkLlAMj/RsyKXWla2dgJ6VJtb1bW3SYPNEk6+9er3Mf1ze7uS+y/EIgq9CHGzC
rpR+RX5vyIq6S1ESRThHbUJi/1g6PfvJVHP9NtH+6LybdXREjEDzlUH97bdZSLDB
r6wDPVRZOiCdJ/x0k2OOToUzCy+oQX25w6ti7iTrdVL9wWsLDz58iZU2KHtEd+jE
vFOI60wNG2nCDWVGbK9i1IbVINzX8c9u/Ajl9VRLT2DFWLzx+fnLs5NO5EC0pQ4D
8t8s/mGbmzk5QPuB6CtA/jb4dT9uaUjfc/ygABqLtOn3uSDHMOmUSRZdPS1/GBtW
QcQ1K3lT/H6HEMbfP6Py46ZADlVdRz7yac9/Mx9bXxrV9mlLRGcBofmqg0AvvbJi
B/pat9uRf/K9LCeg3sFMChFbKjBlhWwH4GgNZYAWWW7TlQFatGZYhcG25pQf8CrX
5sb6bu9cOOHW4eHn38siBUWZTaXgSbdaxWD+7Tfn4vOFTwl87syyTCP0oiXLOYBs
BjXSx4IvG5MTboryBCfMZG3Tjo++bylAHrsQMOKUJkkZVIjLi4isVpfCjZprAPFd
SmYujJDPYZO7bQIkoKL+PlJTbAYRTS4IRv6n7sKhnkC8XyWcR/GpbO+UKsarPIZ7
4LzMwSyrNdXGRxq8/iBnqmPJN8Wygy5K1qwN/SsLnTf9ViU58TiELXNkhUuwmKUp
+fC7mJ7QpgA1E2CD6mlXPGuy6TCXFZpruu8ABoL0wcLAdVTEPwCD0CcqBPapY5vs
/U/PKqydGN4xkTKTD8qj6hDbjX7D58B1gGDY5XOihx3ejx0HCBrWVcDFb3M/jueu
uMmtBM2eEt82/SLkvdlIUunbw6cQENNEfFWYe8a5qdfHfu5eeuZXx6CNly6Kp6S6
75PPMhNqVr5ZUvMoZlRcMFcvtv7qHR9L1DcoPvo+LFNoImzolb6KQQn4242m5lfU
Q5klMOoEm3Z8zdf/reNS7AJnbCjwNNHhgVhVUZrEGb09jxd5BYUtmqo99pky1tkh
Pp9l8Syx+sBHvuLp13mvM6Xv2ZGUfVYeUhDxIMwIDft/47YqiHGHZ0UhrpXJLEUW
aLG1+RqGnj5jHFmfGngH9Bf4bq6S5w+2zPdYZF6D1VASIFTadI0WYFY2qow76s3L
xsrIJmni5ulvihZYajvnV0n4ap8PnJ2bgFWuGorPxiwByjmtwKyrnorsO8yzAqNV
PsDtH4If5WSv5bqmgDXKwPyXOrmaHVPIKqVcMN0OzTZTis2ywBoTS8GUX+yKVdMI
baAksjb+1OVSYWEKQjRLBIGb7uhm1F2femWHaBNk3BkKjculo6ZAERs2xzzj2Iem
kOIJJGolUOHsq/lPNyOk49UtTzgHqDRn8A7idP2DC9SdRaRZwisAlPseb429IeSO
KAwZ2YDNSCwX2AS6lAijDmq2kMYK7scIXyGrKN9lCAD53igMAM9qVD2xA4uR/0uR
1iEEXZAL0g4fI48M7vyJjwzZ77nVqrZQ5SJcxaSJbHcpzlCaWS32IAgNiwc7eR3z
QuF9vXN6MbmoWgwJqpUjTkbmFH9uDWA3CYILyodoyE8LdrvFz3+TeKfMBRmUFQg2
n6Vv5MG4teUNphWNqajG39kN803jcLW/EqadCQBx4GBrO6JgyO+vjRgKsCr/hAid
dvsBYV+yd+7KQBXZEaosRZHliW/u5aQ3+JCP4aWvc4Ec9t2VcrFXIrx0ptAMLCLt
1jBtEno6jJTZ6hZY3im1fk1BEsPN6Wy+X4A4RSGh2N5oQb2YFmS6hBAYR1sjHCpS
MzoVctycK/X6Tt1TIQ4ZlSDO72spxj3UnvgXgRuGym4Toc+A+UJuZzuoi75Q3h5l
PL13Dv18HQBJu0HbhTF9OgeuaP4n5lG7wyWkjSpxlvspge9SRpTFMAB4/loGj/z7
QzzQotzttVtODPjc+ckoHMF87veBlzN/HSpl6/XlGmQ7F9JyqjJ/727s1N+HVqvF
i1bJncTSx2S1Ickv2FAFgLoCytjy4iNDrWUInyd0zFfNuHQ0DYnY/Lkg3B+sWpY8
jCl8shbHkcKa1zmAch2G+ja+lwVZ+gCWeoE1sffKF+StArMK8yXU1sI+o5hkXfXm
ydBTeh24mFxcqPFoAJvf9iRKO3NU6FaPzeZSIYAyDsa+hA/VsDSO6iLFPXEpVEAP
Yj/9FqoFTp5rRU0OuPOzZdBy8uAzcjaxai6Le8mUmk4xDnszYis1pmLeyLQRc8pW
XZue35LlqnILtoi2IeIBFsS8jo86qvEeND74lhbZUAZgLQVZopcfLCkbGvyz0jFI
xg9DJLc119WM7qJJX7dfgH0WF4alMPXJ7p0UxO/j+rMLtAOacJNy0rDSU1CSSWZS
BMwXnUU5FKXbGSM4tj1aZkvgalxUj01J5FCEr+ZSHjQq/dwOyDnAeL/LRy+FoqCc
Pxg+1S6svGSslYGH7vzdz399y/EmAtUZvBhj9jbQTITjkZk+KuI6CGuKHKtY8N0H
RrA9heUrehqNXfhGp3D293EfBcQK3PAgNilJamUkIcMz8dS4Nn31ysve0wpQkJyy
fOXzA1OxFNWRDi3/qYn4IJH8fkuAPcSpqw9+ytdoac0TFYW0Boz2ouT4MDrbTxuP
HQeb5Ml4+BlHCe4XnEdnX3i07ClM0ANZM5aORui7Vc7a8kFe87LAqr+jcT50DjRb
dENviqbPspk1P7NtqrK3yKVXCRGdCmeXBeExR1T6AP9ts1f3gssxVXaL9Dvj7kHF
DLcEi5MgFHalEAhtib11c6oNVUuIT2lfnmw6FWyjqUKEoOdwQuhsZGL2+5qr8Y4z
1qjQDX7uUALzhdAS2sKG44LyOdzpL/Cxnf1Uz4P6jPVZm1atZr65UFq69k3B2zMx
rHGQljZ1SJ18WzygAWd/aov/VVXOI6l6l/cDyMBvp1jG7hQQnFnH4zAZiPzWXkYK
/VtrWBtumpq5RDXKROQweBhlrpIz60gAz2K+4PaXZIwxfGoUNhsf6e2U82KZuTBW
T48gYXQDoXtNoLgiz+U/w6WVEyTeOKPcIr5Yl2f/lwaB0ToOMpjYd1laS7TtAUic
vzCZcZYrFdrFVhIhsmpykgSHpU2fvTj3i6zcb3/C+AmmSDmdwYyGrSMPLhMRKyzq
vpK7o/UCycG+jpyTlHwZjK2sLoDgUVC4x0f6EqGTLG0Ota/eN5xYXxxw3pUvwDLM
miOzF7gCR4RD1i0BtJVT5kgIe69cbKrD89thDwAPcUH/FIYjS5iB+U2ZSkw1yvAp
wB85e+A/xSSIZTDUz3cxBcbMgBCV8GUS2DDWqcKpdaYP6iVAzacSghr/VbV0qEkD
SmnuMbj1bKiiwd73e5T4vtHzi/lDhbrMnmDxyK3IDMvD0+P4RJF4k1dQmmOgVz5s
nnFhPrS70k6bCW8BFeyXGOipOVs+dovKL65k1U60fkmAi9K0WnaFhUFKJggyKVLP
C/NcDIPDETWuvg1KijRlL2bDwHpBovu0N+Zz7O6pFP1stB/fhd2SJL7cS2zUJX2D
Ig7XweqObj+yNNJQwmRx37iyjfsfl1tBBfvtBrvR0jAxjdhEV6nBUMfh73jlY8TL
NEdDnIi7t+pYEsuK5scvBCfspOrPtk9SbwhiZ45GJlh216Mhbhaupn7nrLvRxUQz
qfy6lgS1pQxH8eD6FPZrz7BFCO03ckIsDFdHYmZ77sHsSeOZ0vt3WPsFLhNs87z9
qiRiOj4TlZuajcpI3Mvfw/EHwTIbdRURTKQiMmjSV4A5jfdgfnM+ZS35zuLfc9KJ
OtjHeq5xlO5fIF2NEiPwx11mKmKiJqiG2Ow+KjkH3UyX3YlGzNrxDQkIk7EEWFT8
1bTdveIKjUGBgtfqRsrjUF7vAoUNPtdnsMtdFv8QM14oTNI4jiceB4ETo2LXZfiG
Jac5p7qwUEs+XfK+tNYU6uxtxLcV21ZIvMff4NEKnpinYw2dChup0Jh+HyntybvS
OLxKK4OSmsgstaf+RD6oNC9XipQCt5JZPriTqcnj/v4+/YRjCvA349o0Y0+Htc7D
VjM6WAKwNIgNN8nmWJjrCfTywc16IPyqmw1i/eO6k/JZGa4W6I6TG8DAuhaiAwc/
hfgUuN6t6XIgl0eUys7rWt1Txywd3KOiftwXh3yEt3lp8a3bLOPc2w+Ku7wFVIvp
/7Ety8JofZ2GuvQWTIKso6eUI5VGeb+ef0lE0I6I3rQlXP+GkuTVrP2WIHdgaXEm
3u3bZfZfUKwYtA35oXoOd93m7VbZ1jwdL6HKdoqjnqWGu76yZPNtYEP5moWb8vb9
HCjKfaTvyllqh75tj32wfZ/mncwy0WcqBdV4Z40izv4jJATKkHPtcQsBHzMt9xg5
DKqlclfzfTc3U8e/p1O/PALDXwd+3EYQ6XvQQ+1Ieq92Nl7u6KCe5LSoCH3oJmEl
1Ak4zt4ZlCp72M6RLVlemV3pZty6uiDpfYSrvZu4iAuKDlgqol+nDm2Z2PsL7O1H
C25SYTxRk5ymoFPwgPE1JZvSYnKLpiQ0uXt2EkQd9DvwIVYAgk/fb/4lHDK3VIzw
sxtasZcsbPS0IvtTX7qMEkV1it3i2v3xxYSUMdsYLYC2HCjnmxmVzgjAsx9Hr/c+
v2DvMoBJGHHxTH6fdgMclnB7u7hWhFbgsqsFtWH+Z/GBHVvWT2viGXaZM/n4NW2v
XvKMviC/yfANHO50G3vEDBFojm2JOtAEeUAw/7IdYmFiNY9JNW968wZVs0adQC4T
tZ1FKpZQKGw16VEY6NSyx2QuZxgLA8EL19buPGNJhlHd5DBDEezw+Oc7DOd7ezdk
5F6NqRQQSlwCNMiArQJb/qr5F9Z7r52FB8zshwcATkxuuMkgzzCWIa3qqLr0iqq8
nnUsPz80SPHUDKEQWhbp5nrN4LpdbUg7A380hlnHSYpftCkuZ0hjp+k0qJoA7gXs
T1jGuGq6dch/RaO6woitGEIdL3uxjz7Yc3VMWUWj/jmzMNx7SciKu7L4aP8gkBMi
odi461k/UjoHC9bJrsNQ9VgE36tddQkN2SRfmWHPeiLFPrdHt4GnQ/9UBbixedse
T1F7QHasE/x9kQ9zG+dA7DDQmGSSlKrZEOBbUfBJpMa9BAtqEpW/NQy+tjtPz9t2
wKdxmBDbfCFeyuMfkLJphiuU73y5t2LQu5CeLvxbdw+ECk3dqzbCd4ASy8smkxR4
vcUZZE8BoAVvlh83fpyDuIwfIJH72Rzqyl2KO+i9vA3tCNtmC5JL8WaeHKECO5t+
BfWJ7TGWZ/MNVZvfXUwM6iA0wYdDKAUgGPBRUSOIcQl7EdVxjyHOkm6P5vlVftbv
bkL5lsdn8xTBbCu9dCOUB76/npRxXxlBkHJzVn6h5CyMiwCPzuvYdULfEzIPqE6t
o0K9vOWN/6RJiI6uu3YrxcW581/Xvbd9qRu9fcpv+UwpkRu9inTflYky/MfxKhVY
kr9/lj/Du0ZGpauXuVA4ujSn+8q1mqg9mPL4xDDIva84lNjNxpAEPFe9iprKyU/T
0pMFpQabaHN8SMHAVJxZ+NWFHzabZfm6WPVNf4zy1GiM4pG/A1y8lu8IvfVk3xaK
WaAq1HTHfMj8H+ntU04DXMYqAOsnXWQQQwzCNRMHL98sbSBCLfncUWG7FS0ciHGl
wYC3GkxfqIRHaKC4M3l8oTRyl/6eJqnJiRIyhMLLGpZQuc6QPFYgUpKBEQkM/FPp
JrkwnlIxdc8+qVxiupO8IYJkV6sfqDCAztpj1e0UwAHgrTgr+KMxzpZ2iS2CJDju
zZ29q1gsKQkc5mUCLh01Sxc3xsIjQ0xxRFVDnSWfWXdZ8j3k44huh86aNPY1dgZ0
MxO/x9Ic4nbuciz8JXHZPIzkqvw0syfmP+FJtcf7fl8JWrlQ4KqtV8khXL6aHWya
SamgqlP9kFI8FqZTv3Mt2HTVhb+AQCvoSamVkf/It9k/r7BHmdQp23XKDEHgk+Kf
COtxmCH5mzo7OdWcP3HZtZ0D2zaemuyU7ZRkG/dt75O/aLmWqs8wZON26Dsfw3ae
gvrWnnE/EUUM3LEIcBCUyiI0mUzA1WaUN2PECVaq0K7dkrNB9BT6AtoYC7wzWvzy
Q6/CKOEdlluMG0PaJ+y2k66WRxdgio5j9eJpCd6GDo4BlZTywU2ViyHXC4fWBFgP
WHiPMDHSo4AJNKT5CoeNB21+B+qRCMlROsaOp677TjLLOHv3Bq4alLpX+BfJdf+R
P/VXFvcgIMZFfSD8s2L2qRoQtjQuWfa6RpNTYFmfgcDSfF/Oi4ETBrunhtHtxLjH
evzi2K+BhLYgWYsSjb4/3yc0m8TlwDFx0aDkSPz3jIRAPCuqTWkcljT74Us/00do
0eR93/HFUoX/1UT3vkD1vhKaG8iCz1kc4/yOjgE74t/2CE+AmHum3sqkQOCb7hUG
mogp0redp3HAL05fr7p0agXkF9ZHfWJAr6haWMrPuntEQbOvd9W3yaLePH3g1f2R
lE0pjckoY7ZApyUiS5OLHDQWF9Z3zBtaR4wREOwAY4UMZmvDMJw7q9wYpEyYaUtl
5qnVgJcGQ54aeOoHgRcHx8tL1unGDpEWLEx7BpxyatQF8ojYVysFpYGWQU9FkIho
jHbdNxxxVB3bR9N6V79/Xn9FoFoKJGHtVB4hesWU9Hm20Hm1Rk2BXTJ+iymw19o8
PszhIcorgudVUoQnZQ7LVejhgxvKlImKMjElCmZjFMewdLekrADiASctXZIlP92X
HulfEFNijOpBGbSfXjBYlanMKx9z8eBms1jadATa6xePGUu2qjL8kpcsteE6yFHy
TZDV9POk1e3p5m6jce9UIIHEqIX8czSB/W8uKsNm45dKWLnOxH3RMOGRKrDGBlSP
4xs7XWnuNSZ5ko9NTIjj981LEHEYlvrH61M75ZhUXzP8g9uGdVKLDDBJZlauCHb2
8ZdODNPPqtCuaBC6CcBUoh6JmTPOWvhCRJ6bVLgTDjUSXnCxA5bM57BuuUMt/RHL
ptwV/0dikCCCp9bE8ZpOv7yzWt5M/pFFWZRn4lx4M6kuTkHfRa7jw5lhoTcqjdWJ
4JC9cyLRKsoK2wMURBt9IBMBxyYLMOpgoltyVnNTHJhT4AnVixgKphTjWKMudK9i
ALmqwSf6YNIDhFrsc2h6Xxj/L3cwGONWcvBQKZHiX/usNfUX0uZmW/mf0N6FPf3k
R1PedZgdx9en2VLNdzG5htZZgqlgbFsmd5xLgmCR0an9qQ2ti646sU/GVEr6FU6I
TG8dJXEJYL+lfNoj8Oxypo2MSvMv/gLbin2YwD9d3IkGS50Tu8F9VhqsAO22q5XZ
4zJJlTa5hW1bsVnud1wyfr7Ldnx1DA0ONX3RxdZmSvwKSD7tvdX+TbZMkK8RQzt5
xS2JGrNliaxLiM+LuLcgOL54bDcm8vuRsLrh2AKQYmze2OEZSrSEjPd5xMbcBMHH
DCIc3F1DYVrxJ0LyMAcvMEaZH++UeSmqZBB1HhMpNa7xzKmEqIuhIiFlLL43+gym
5JDTpKv9wv15EzzCAI9/qQqV/jrCePQNFXxaFdc5khNzJzPpGUQXkUpUXhhvUZI9
E1lr7sK/8+V37KWBk549aV5z1TLk2ecOU250bFmKPxay4Kh0skgrFGcLTyMx417r
vD31pNO6PJU+U86VReqU57CpH9Qs2lvCG0B6fyYj+HnykVwT0w0eJN5DAXBncNWM
3uUGO1+RbTiqhrokX1GGwNSaufy97df7Qa4Q1jiBHpDNcBf5JmmlhVswrAdKpGXM
wcQm31cYTlM3JOzJboNq/23tqUgXuxvtEhLTzm0SkV3st/EsqXSxNUYtM/aLa6rH
HPBlmAD9dbQSsFIUkLwcfTV24K4QFN4z6AVwubEMG/YlPhizgR1vP63V4lVWyt6C
E7WI69drPCX5nlwVTDv0gseyhlXtObYrNHy9cUkbIVpu0qmDQbGQMrDqw+BFwFfy
1u/tqYJ+aYsID8vZfyxYKvFC443YAkvx/2Mum6/uCysov2iI4K5Of56xVM1ZeloC
LYl0Th4eNJ0zcDvhneOyLH5wD8TOFjNyGQEyuB9GeICbwlQu3bWfQGPjNQ0ygXnU
EFcn7+V92uxyIfvCHxmbgyQo1JBjM5IclHPRPVBaeeU2hw2IbzztXFq1/YOEZ64V
/fGKEjZ+nBvovmuGqqP9M5WQ09x8Wp9+Uvtp3I1PNEbZhDU/fOo0LyS+2KnD8AQt
tYEZiGif1qEEujZixuKK6pj3MCZk/Wl4yHwUOtd/xg2kHcKfgL8c/iplC3+SmGSm
PJzfzJ32Us5hmxHoQNMPPs/hb+xfF9ssNZpLrxKYSGMqN0CVYRkoPjXpR4NClgyp
altGdwQai1UZF3OF6NvTk2bJ2MjWyzImIHmHvRk6OmNoT4Boiap6nNgfK7yjRXVc
7B+JPMQB7atxLI8Umdwwjq1SzRkjhh/WMrE0JXQKiHB705O/ZU5DzRXn+H2xz7DQ
biLmd6LdF3u4f41fAxlThPes4HDIRqt+ZIL3msj832hG9ZGz5D0kThPUkf50YE4r
0Y+VNPQ4Eq2inktfDgrOeK9LFG1N5LMDPNtQCxi+ZZ2jMih2EoZtHaR6kUV+eXQC
omhR0J9ZIp7AiYLl6juDkiZWbJy46OYeVTxYe+J7bWavH8sEcTroT5yalLoiIOaR
GA8kD3fAygjy4BLTyHY2KmNa+WBR0T9iNCxUW/mgM//IxL/dlzJpWSeYlUgA6b5z
TmNSrF7hKJd4JPJIy9E8NJsLx5W5JNSqUCmhQHw+VzysaCQeLz1INy4jqGpr2kDN
WTPxe969y95rMSvMarOgMKtXY5dFXIXUd3Yaq99tqudE2nI72TdheJpjliWjyblc
IMxDOiNT1edq3Y8Gsx8HRMUECEJqu+7sfwmxDZxa8OF8FflQF1HFcq0YWgpjoxXn
JwXplA3EZ0Dt2bOKHs4pe8kUBgZOdKngQXurDUnP4QrXRVM7FEFDlVCihosMkCHt
3kzmT0lnt5lSlZyeea1tMg3tBuMpoHM+MmWnd/rA57PQjOcVGTBZ1E5CYgFw47up
PaqksqYMAppprnnceLwQfX6kqSMydSybzEO9vhIQT+TyXTeWT30hefMiv++bgn36
AL6/iEgyh0K4QPmIl3VWkE6HAVDJekt3xD8K3UloSd8oKb2TjIMM3eNtxMJYQVSh
cO05Hwm9WXnrcMmNprl/+bO6H+2uluvPIPApwWl5qCAGiIvvDw+qP2jnq0Iijiow
IsSX9KEjK5RzddmBp1GdhKwvWEENdI8j9ZKL/xSIJ7vsWVrPVFs7+oqQEEMS8xst
AFsUn/f/o0OyPg8W7tZQH8LGw6UC6yqi0/DVdet0l00b2NNnRwYS6HTKqJOTdPr3
k0m9AhK1z5H92ArCWt8Rejx5cROrhnM25so3tx5pohSlwulqyVJyEJdpgMmhH9ld
OdBTD7AUy6U5z+8TPZWQzFBAnamIGPfUURS/e6ulnFI4BIAs00SeBFYyDSpyigyA
Jg0chq1cAcOctlCsU36GqBAYVU0v174IklfqCK7bEckdKK7yH78PIQxjZNX/omz3
uYyBjpX/YdMaaqpqkD4D7pbSPLHqudWhtou1NcyC9UOHN+rG51EqjHUgmNVRvouu
3iQPoO8QFmadTv06lB8SeB78+YBj4OHHxe3ne+aMl80oHU89AxydklnS7NEqQN0e
PqMGTi/MSSZmbY1Je6Mpn/nxvjULui5zoj2U2tMBNZsT0IZkR5+VFWAfW8/WOxR2
YAtYKJJn8hv+jUS2BBmzRS8XMLaLvsqzI6Z3+DzFU6M76zyd2cGVYnyB74m8LheN
GdAg24R7i8VbpuhfdPihQDX6DwSzH89tV86RhW5eVoCSHGfuMIKiHwbu4tlMM856
evIhA+9IN/eivK1RgY1TyUZsGMmZgcrCH1IbmG433SCZaVDPw9p301nhgcF5JpRF
mp1ZugBEiD6HFctP40W0Kx3XvMjXm2+91JBOTxZa99aJ6+I2bjouHJBKYBD4GHjE
SuEBCBhIqlqU327Aneu2+g1UE5aytNY1OtvzTgnnTip9LeTSjkcXYQ5Ot3Rb+f3k
vVNznrTY2JgpBtMIlSJXYNESzTkg3utww56LC+QdL50r70wY5jTu1HbY1UMflKbY
dN+5gdW8viUKvohmFlKMEDZA8Hp5W1oVfhUUjvUdLOLV/bKhPgwLtqmd+UXF+Zht
idgxf4/ilFJJ22yr54Wbw6PBJpoE0UB50kJt+TNHURlrmZBOTZVhYkHymqcvEIdT
pUJ/1aJj3Aem2Vhul0eDca8uT1Uf+X4Tw4RdEgtEm5rKdNDyQd35WvtheX/pd5HP
SET9nBDAuWapJc82t8se+JtmfchhWMS0t5vGV1wMORkyu6TY3fu5lk4J/NU8gni3
FPRZw8qioO8b1uRFhWl1qXzNFrvr1XTFYRgAQZijCaMhlZduDcVlctPbJgGOCGp5
sZ1uWbIU9b7hFk7IfgC/hGj1A1k8igNErIQ/xKO6oAJNMDoOGmu9E1/gzwYzm3NG
Fs62lQq3jXrEyRpdwMYxpsJggfIOrDWK6zobdkuQxtIb0O/eBSZUwejIijU3ylO+
QyymDTXmxhZGTye7e8YGkUuvNF1DE5bx19g45HFoj30oi5cFJGYM9xYY2RoZoj+U
RLwoEhKIdE/ZDus3sfg1ZN7xIIUFSVy/I6YkYE+QGfpP/q9yU3BI6WAHn5cJfp5p
40/9jo//V2VR3CWn8IygIgBIiILR09cNH57VwoKVflxACTyGD/paMrd3fnkYQtrS
7wWhswu4HhtpVJUmeCqruWF82/tTUHarZHSTR/K0RWKZMXh1oL4wMGIMG1Rvuje7
oeeuCq/1GeSVpeNH9z4TdXmvP5vBFTJiMx2tW+63dRpCkvMftJEL85VwcoUD5wAN
okDDemIxLSZuOOztpDj8Y9f76yqrsV7FatweeVFhXDuTSYNkfmyWzXBUjZVV4gZq
3OtG584SCciKIgEPAb9P7KwTYI7pFzR0D2xnogGgqjytUuwmwvCSVlNhrQrCUFPX
JYEn2JHkdtmecqfGkukPJ+FagSSofmeRP2jC9bOUoKSgMZyDhR902y+XTE/EeU14
rmNaPeYdFWf7L0I518RcmRsB29FXx8cYEq7AeoSkzGR+XmK0tKng6FIVFvQWZbva
dyX8Ki6/f8Qzu6qVfQ0chQPUUEonxAwSN+mQIDLOl0fD3Bk3+TK6bpL6GmxoixxY
V8Atm0zm/jcnWKRxyOqDDH+MM19mJlSDf861xXTK6syaGjo5XYVdnliYFBxlg/0P
fQ7fdX/UzPvQebyNtO9RIziuC0z+kR9ZWSn7WUey6L5wjWlBxUSqj735G4ED3bsn
5a7t4Zmey6H2Vy9dwC5Rb5WjvEnSTuOhYYEVnEq5JtLO4ULA7II1dJv0rb7eeVBw
snCI4sN+n2Gevo6rLDiucDXvx3opNf95wClWsjGc/1Nfgt90yOYE8WlLZrfHS4ua
ILfGGwvN0O5orlx+yRSqj5drS/Bv+/27suIEbkS+25YNoaTnPxB1+ylR/HZlx8mV
E9YHzIDVKFjBEnKIcJHzaeUoG1lCE8EXa7NkkrxMBDrZoUfLKdKG9SRBuFd9emIH
NXyU+1fcAjEo2s3zI0Me+dbo79pYqCMZAXm0q6pdg4Yxafd3DkxtV1Q8lyhK1iJE
oTgkqaDcrPCOiNFE4cUJF27YVlf1HqUfcL3bPcJ0HtSVaO1pX2TZLP9UwmLVnePQ
FAySB4RzauEEDWxuEqZUNP+7hll22uByjJXHQKi27olHmEZQzJPhUl1/tK6xSPjl
dUsI0CLWYM3VFdTQdP5RLEYas9IbEtaRtJosyeNdCXtbP4X+CN1hiwdI4ofVz14L
hAY1b0IEepbcgtPfRkAB7O4oVJ6QGh3FkJs1/UuCLvLrfBMnpX9g/rRDIo0HMLvt
+NbMfqqkjiKAyzdC/pECC/l4rBsw8RBzMWko7xGERAU7ouzCdAuJddvBu6DqiKDu
VY3wCBUqttQh4WjGQ3WTg8d++3K1MpruCQaib9r4ZnOyJ2o1mOBTut1OTPe0MV09
uVLbHpCBkw5xHWbZpexzopsYm4AUoD2wuQOzxtNFKKzixdNrareqpN87GhJmDdOC
yDqxkYsKK3FOmhizLmOz2UQX5lZRUGcM8utrnLpJDp25qb268vAPgnq31gGv2UsB
DmoeqIbKKBY7aMbKfsGsJqx/yB2vfOJC26BEPwHVlhIuOLY8x5dH4SEls+HURMnY
YbXjcgycOb9JfB5yLDRvEYM7ntQ4knhli/oAvdtE8Z3rDqVC0LQ52c36ynM8vtkg
E5+OKqhdJA/PjpxamhA7HU7qixE8suI4i6pdIel3YunWN7AbWbYWusE5PD+nd+47
rjOBRvDP5Q5YTOcWEdPqwvvEcAQg4YQ8Kbxu8ivwSDt2Ilv3kL4s3YYzCoXKj/t1
6Ke2/MdlI9vren6r2QxSobPmW2k6DJ1RTMqt0PmZ64pTEUVevG8fdN9BIfNxUD0+
DVOLxIDCNqj9xiL/W2JrU9UFJv5th1wBvP9m+FQMBPCUuKdf/RPeI4OFrAwICuWX
ZLr+jyWKH9GJwTwObIriikylgYXVI663EJrkCmIf65ug1wYUzdR8GoFT7GUT63er
3szgBHvMeBm3USU0iyV5hRRwrNxQdfVVuHbkgToVvIbWgluFznRQsk666lqDZc91
Spz5ik4jrxrNPDxTTg2+45bUnE1fMPQeezQX9w5Ia2+oX588sAJENXM6hNzhrpDc
Rd/rykpgArHIxZsO7Yur+4fcdtoW6NTOQx7NYmDexdt/3UkSWTvJoaUUL25oy7Ok
Atf9/Ta1/43geNZ/CqPwa0AHzhSiUAMpyFsGMYcpHakDb8s/e1rPSgTr3gBrnXvC
N3/jNnYijOliVbEoGLR6bOgbv9T+Wlj8I8IX23+iDJik8KSSTrQGNfVKXf3pfXcT
hh3q5ugXW6iUzFMYoj6Gtz3LRZBP27GLk9Kb8T9ZYBQfqZEEv58o9fN4kzrFV05M
gMk65pmNUJlp6qO6aLGwFPYQrx+PHR4Fw0aqYJsAwkW2Tdu8ueYJLTlxMTXH70uz
Xkn1HSWZr464pVEbpbzuLETPYVwvNXHOnmtRvuHCszVR4KX9L2B81I5i0FA6sYME
q6j86we5k30Klv3O8nJLobvRYzn4UaIW9Pl1GBRD8gN4jcZ/x/K4wKeDF/quZo2S
wih2iqROHhG1obJze0eo0WEZBzhR2osnHGKlYeCdlXFvY/8X64ILtznAgLVvf4IX
ewCpm0YiT3DNKdvmIpyH84cf6U+renmnLBTcxcuaJfJZwgoZOYkzJh5tAV2Kb669
MDCZ+6Kww3iX5K8odK4H2DEXXFPEzyBf/bczeQXPcRNBpDIWZSuepwYqRs5ynrCX
QSBieNU2mHscl92+3PlkCZFZhDnTdgd/HQT8yts8f+piDFghCcKvNnDfjmdKgIEu
5lFZRsVF64XIlLcNgEEAMLvw4k3FBPbl4VHGSST8osn5pqp9Zs89FsS1pDAytSh5
Nf6hwLjU8KSRsQsHeXrIW9Yxnv/Xn15xo4Swx1edf6uvxMigKRPBK6ew6zsIZaE1
GnMzrnxaf93xZ3ca0EM91EigVXXVwvH8WgwtYXA3Dp/BTlNxQT6zik+FJ1UvmXlG
HfoUuh8C0/+x1pC0zq3Ir1LgE6NF+iRa3ztKnzFPUBQk6WL9Lyw1980FiLtWRsVS
aznmqNMm+OLoP9Ic/+5oKvzYWzNwqphwtuClRaxSSJ2aiPW1JwwvceodGGrZqtHP
INOVFR49WcgfiQIpRFAAbJ7kA8Yjw3rGwtjkfZSc4Y+a6qzBV8wHjqpj/3X2/asJ
6FUmG99eZw301P/ngJNK12EXMjKtwKqdFttW0pqBgdRk1NydPTZfvHzU9wpCrc9A
a2ajVJk9T21Otp6WK8TsAwMp8/DWOr5T8SIy6jkW20R9WhbZObus6JSuT9DQS/j/
wiKtbDzB/CmboAoL1/kB0EnmD2JFMdSfOiUklvupP5v9Kzxs0W6CPlPcy9A44fQ9
P2FvA3wUHp659KesW+m3tjPWdn2BCqRW3QZCifWlURWFz1lMeVoaScbmo7Lv7bLA
+WQpnNa+HkPFaXZZll8yrGF5YHfmio6HdFsc5pp4WRBSdT+ZuM5KUQTpjf15dQ6v
pHu4uztt9rh3LOPvza3LaPwhJ8Jgr4XA3mQvgV8Nhl9z6dVSCNp+z97l6coqrWaq
lwve9n/mzyBoX14m01YBIfwX2MTXQ+e+EOU5R+5XV0nrPZQ5rU/P/x8GS2foqqeF
mLMV7CB1z4/sPzHNFzAHbP0oiBZ18Sp9OoDOFYpcPutIc4CEk7c2JLnwguo8bZN4
rsCCJOwS7Tim5eGg1pZJDAXuLwsLSLqAOfZ0w1Uj4nJLXGh8JU+caZniyBalz7V+
IqW+IHNj0blFNs9PXEu8+CkPh/2GzGU0p0LIHwiIf44039V7TErlYFDQZGvLFzI5
+AUq0CHvhhNXeUS7c+yS6HmxuutMJ/5boftFFBekoV98vOAt7Is2Kq/KVgV57hhr
WoNb8pj2a30ROb4G7pcBFCNhM/O5JHEka9lK2eEzfpTB6+O8/lizf7Zx5osoTWUY
CZ9lMOAqJeaCML645vUXeth8AlxrJoqXcEAEtMbfscnXxk5DpDVKxXwER0fKh5/0
78tyadl+0i/2onjS9f5n0eoc24i+cL7ZIkmrzkLiant74htQ6nZroFS9sXiyUKJc
2cnHcM4AQMzjDItNgImXGusiLIM2jJkt1/NM8b9QwQS+MkgQyFPpA/ZEU63LLm9c
DxwHW+NF9rll5+24Ov7ZCHxOUBnn1zXboVkYRG45gMjpdGnIJw9hxHt/eYAh4jdA
Ufy0HChiNxgwTbh+FCpw96hIc0G2yN7QEYR1JpL7YSDyEKIdmL+0oCTvWTKsb0Oc
VQETBq1xt8rRJXL9lme+xmsK19BW1hxtD9gTjbmyRm0BCmR7e8sRSa7qeZPee6wL
6HIhcEsbOJ81NPXsP7AOHBpkHmZ5i0Y/ZUnyGKO9Wh3l0crAT9MyFL3uM3vRhNb6
ZJ906BrBmg4pcHfe5NwJux/RjACEUcoem3TygLKCZMg6UkRTA14wZPwSL4nn77s7
A9OYeEVWgp3MDf498X+E5umLnyObvRMkgCnOjznSmxacr1PRwmDj/ZvkSmrjdgLL
up/GH4BTv5Rs8rgEAPliIA+nqoJP8phgb7SkL7BJthbVj+gqEW7EqeIN2dyt+Nde
6vZ5gEoAp0YCosD899kalbaLw74A+vv6LUxy4GdawH3X4pJmfC9J2UPkSmlnra/L
eQ1kyE8oFv3Uf64qlvtZUSmY48Bl9gLX6qS46x9Mi7IPq/pl/UYoxX/I8lhYcx2L
awtErfliKGkLGXbwqBR9HiSllPBcW49V+dHze1xXB5FgVNWEqpBTaorv2PvrE+sk
pqdUbnKtwQq6eJe0ayCTxxNuNpvIyjGbiZYYc9hVrOWBTibYz1LeFx1nIjhgv12H
1pgosJ1YWCr35n2uVO0LCzTWvhXa0eEeEWbGzc3k43RC/aLaiiHn4CqOJiYquAtp
HNWjObgtVhUqUQXORVPLkhFJ4qp/QPw4jpBh5LKQ8HKTaBSpe7wegy2I4B+gGHu9
rA5l0MVjHhazMJsncmLNPbEwDsOYDhZQs+jk5SabtyZGlAywjHh6IBufm3tOgyi4
fYRw9FNVx7U3gI1N8BCKM/eOo3WmBj8P1Bcn6QD6Ke//8+ZP/y2mkLqkRiIODVqQ
yai7xe2dod6v8M9tunvdV/Z0VsbLBMmXogysjZUoonpDcfRg8BuX6JWZ5sbL0d7g
0/Oj+cpk5bSquL1aBEVG5iI5BT7CK+/g7QdRF3Jkim/mRQGhfgrGRujSWewZP/Lb
kaJ2XZoNztiiqIWQu0wcGpUr13jwU2dHj1JzD3XpgP/9jTLznrwricDHk0wPbHYv
Gvi0/vy5ZtN33yLQqQ4HEbahzDDp1kHOgfE4n6xDcym4LaD6ihE39iB5tZAaR4DP
u/hW3vY81Ka+qesDJlYSVKddhTWhpw4OTUwZ5Ul0Nz99iCjJarO021MzGNyh+UHE
w2OtakHUWsePiGAh7db+KdQ3Dg+uduVVwq03792Gw78Q7BicoqHLJ85EUvxP+erU
ndlFsEsoTmaoceTjFeFdrYQVrhFpAVFFeoe+taqH54FB1VKOypnCvIauQu9xOI2L
o5BNUFD9lwdAY52adembo8K4k4EaR/O8xeStvBZxMsaslpyI4bSYX+RHMZAOGAdy
OTa/QoyQz7jfCkIJEwKWJxt3g/TqYsTeP/ksgRPvGTMDji2YhkaAGY1aeLyvfTAv
b/6Xuz0pvMvm2DY6flu/PJfOYgcG4/Vk25KJCgKIY+B5wd2SMOabjr0lBFdrw6ow
pEHhjH2Y/LX9ihYnbmbx+6TTIHjli74x8nkRC154N0F+YQqWssXKdLipuQU7e2gX
a2FbY01yVD4ku7SfqwQAB06NR8dNYLoOvSzkKlEU8dT037Tayqr6hr4KDy5CxGVh
BjBh2HIhEf56jI8MWXd7p/foxviFIs5knMr7A3XS9FtpgsjyFtlrZyc+g0Yr/+D3
QZzjBHwQSg3ugCFjRiXGiWDIpQu7tkqPPph/I0p9PhxhsWIJBJ5VPPHkG5xO4BO6
pUXfNLWTdF2cr2IKiUxutdU1AhwSKz/7RuqkFMtNC16HvLdwWwUuSHazZ77Ivm1Z
q/fzQlulZRuTf2/73+8t5dItADVdJDRgsF08czvDh0hZw6Htaimi82Zq/x8YaDJd
MtSrIwfTTgstlQURKkVX0ejT6NldQUaLfC/IC2MP9VNet4rD0fClRo3n4EjblzBH
EZJw2bmJyQQV8pMC22M3fuUDFOw0REmdMH1z0iCm3FE+RGxUviwasQKvqrRJCY/D
BzVp2dvhRcwZnRVp2z/klfiOTWXohith7KXFHsByJFMrt+hXu6BBO4n5MUy+Vp/g
Nmp7fG4XOxoa37zWG864K6AH3yc25tuhy4WoZs+s8uRxg7WDJS7AUhizPVZ4PSH3
O0cFHBHMqQJsOYLZ/+35c2LR88lymo8nFTtzpXXbUt0RKW/Qsztjz8J5LwfgG0Ab
GI1swILvfFpBlnb81KrteeV7Ona1NSA/VnaXpLELDVD0JlIHhWQZ82hN9lFLU9qv
nv5+3PGY5pp1tUUW7QtSvtUss0h/RqtxNKG8eD9SSoQQmRjgCNKLcyisKgLNp54F
ZC/Q0hCTcjytaA3vfc2DgvMswzK48KzwMsqEioO8kkvBqz/EBWbK35vSgz/hLyQu
WiPAFWTmfM9o772j06Y4DRZQkH5qBgLcoQ+7PXjiivRCMFdUBnfp+fNVHcnLFvZv
McBfG4qaVMCaBjd64A10Dgd6mEQqknSJRXUqy7Dmx6NqdRUt8AQ2dibTaIit8X2y
0QgNqRrWy4hLuVuur5fWBORML/m5+Uelo1wR9f6f4Vzf2nb4GNpm1VWMyEL1sl+8
siapcjD4/wt/Sz21oSTIAbluvY9j80EAJBYAzNpQ/dPrMUmaqhSMDzpTNuDbV7RS
aIC7IzuqEgsPhpnuX7jvZeWaE9925jwMJmqZAEZudKSUeLbpL+cwkKiawaVqQGGA
hpL03xY8jMvpstqYeFIt/juhtKjeHczVpPddmGyhwgJKGb1g+pzFuwSN/BrIAW3h
8F5U1mtn9/H4U7XdPULDF+IGFBJvf7jqJXNveaDfFN8U4uM5OvfcNhXTOiUweymL
+aPLJgvKZzkrerDmYlmEAiQTzgjDJyNc+RU1jbdmgZdRb61Okw+q/vy3f4TxSdtQ
+Tl+WUkRkqFPxEoE0ToSb44RsPV+DRr2YGf48bv7qpiW1uxPZdZ0XPtyuDHMsAQB
lwZFS2iQgBYcC4TVhSThF8iPoTAnFb/x+5FkeZXyI2EYHO3XiM9fqljK/oFaVKI6
Q7POdInRzlFIJeaX0QR00NLPgDlH3+h4StrxPowWqP29c/l7ZtxeOAVnMEZ2tYQd
c5aHcXNka+q5w7EyylxFJlZ7OoXoDA6DNEQ2fLi3OyrKbDY4RY67QUFdVPYOUX97
5aBm46SWFBhwWtIW+ktnR/AUVMGOxgMQj0LOM2YIDyb+lgOyPecvheiZrih+X6O4
X8kLzqwBsu4YqGYq99seTPc92kLmd4MdT2Rf0siGZdLmKRPxifOfGHh62BBNjlVd
R9ygM96NgIUPrK6xfbtpo351vaN0Ygrb67LqpmCp/KUBp2VGZ/ZryT77dxHr7a7h
BjwAXgAn5I515SFWnQuIN4Ll6llGIvagfM2GrWNCq+aIhSgWAssrbpCcUQDH8+wS
H8YlimJxuTNPmgG1MuvdjkZk7QvS5vLZWoSLVgUteIVxTMjnoUEdXzu17o28GJD7
KKkAKepbx7NjoZFHtHB+YZs1hYWnarVXRghdk0CjEzOiPYT0AkKGhwxBS0ErFDT+
LukxR4F/zDwhpLlcd8JPQNMJ0yQQmOrxCJavn+NbG12CvKswDN76bYt3e47UZSCM
fqd1KYij/rMN2s50F4BCPJWwqTTYloT9xi1ryXPfweC7ABtCWB/BbkgN7ByWzvOr
h2cPChMKVKXOwDpni6dH/RfmtA2CM6BbB7j8C1NrSYL3i+kc+KbH/wTmReixli+b
P0bRT4DsGgdUZuTT6+Zd8cDP5KGrN8fDzzxSsd6XSd60Ryv7hefUJi1Aar5lCaAt
NKnbfrZp68rLpGDVvDHhTp7AMRZS6NYKW0klQZCXf9sZlRxcuQGUlvTCq9vRHmTE
C2pV/xBkASxQ9f9f7Nf5vft8qLr1RQogfrzpZRpQ6sr9jsd51OMbv1ZVDanbP7LU
TOlfnMJb05hGUBtiGgnWGUd3VKxKGes9Dzvwl6ouP4KQ0BL5Voljvj/NeevxEeC0
ZschY8RA8cWhKEX2p6YQX+aDTWQQkVggzCwpOhIEUS8JqliBpFZYku9RMwV0/f8H
1jj7IPWEeTVrau6zSBJW4/tMxzyjrPWq+c9Xi9cH9qe7eslUqikxBvljGOVJnq6m
quFdce9l/IGEVKYHVVda3/Fevn2MFJ080MKV3RiVJEx/QNTPfx5c3M/ga4zoBWFb
S1J6YJH32TCMyu9eDnr9Lyv2g6RIDgEZcsfZy9Ln3b/flP+dYaMjU4kxDEv2OR5a
wfKRg8n7nUVumSKGoasYGlJxu/az5gR4Bpy2hzL2nP+Jl2lyIl7sckpW6O7G7L03
gxZNLPllMnR6ljWPFv8EV39XcGfQclzPOefnyfiSkHX5yyuhCOZKBtIpRsVCwcCw
MyraShlbhkLR4ejbWLClSAkYzPZ8pM67+W61oUpTybPaAzaz2JUzU0BR1/gsjgH3
Y+597me6mIiEs48t4B2peRmFz+1Uzejms+e34ow9tFMnJmAX6ZFG3MrrzTFp/uXm
w/Dmr8SZkD/NTXpC65UUFMP6cPGeRysLX4onjfa4AKiTlLWyNpJOftE6oD97hsxG
OC4pLdtl69TtDKbNkhHNrCpiivGN+n+xbc5xTDtqcARmW3mCES6tp/alddzTMDXP
JuzoTDCxs/YBcdBb32pY9u6k8gHRp1VE+V+u3HJEgzavv7N7IIGEIio4oYi/FUZx
Z2kDYVNtiZkoyoXoXyIc6qKp4umkOFaqynCx5SXJvaDalAW653pEre6Oj9vO1PA6
Nz1pxc6YlaJIyxHnxXhzD9Ktsp41iEa/pDOaiW7N+vYRV8M6mZH2lQWKNlLX8K5y
QFZ8kHqtBcb5kAAgcQdsTNmpN/o+II8Tr/v/a3FxVYwLXGuzh9VAFO+nLHu41fbo
iDKLKsast4m+5IPF7dJPdHtXBd4btX9t3qMkaEAEuxXwtm2IyyJZOsry0wwk5hEI
Vp8doK2nF3beS7pV7Qly5GjH/K+qy9Luwu8Awo4EpZOp0o49h3JOtWkSSLWz2bhX
Hp6ixSjlz0MWLxhwRILXNeJIy5R6YG/HzL9u5jzMaugfvl8wQqkf/A4zi+D8kzLs
Ldq51gmKcQU6i67THuwlSTDxQGMgOQaE++AeJTSohQ1/aE0djaehNMowGv3icX0/
jG5jEDSTq8GvcCbyuZ4/b6kmuOb7a9xfeVKZAm7pMwCG1tnYDFZ3DhyGEsVXpcpT
mwRdqXUdSZ3Vg5NUXaUr7pd0VVJyrrOVd/zlENse/IPSNWfytEw/VwGQwKL/Y9IA
/kSOcNWS+WhbMGuJZExvIlHnfpOpFXTE6tYDK8C/xfz02shKBl3+kJ8stfTRjRAR
wPhlWOYLMAnrlRGa8EbODVUxbvHDw2XrUJb+cMIrl3BpLj+k5h4QBd69wKApuREd
ZM2GLzZ4m9ZBnFVnL284lPtSb2UYINuxzy7tAj7jD2SLT8QLcYUvuvbL3J56c3n1
yzWA56iDMWkbrl1q93pntnhh235h3Ot2nk/EgwH8Nre+1nic/QdRg9iJFAnbAegP
LjszSHru5014NvhEhNQR7c/+G8bb58pQIsop/I0A1uGb30JtIbgBx/xXODOWNPDA
P41GmtgbEKuleXp5SCXfqIZSfbQqx31RbcN2beEMHjStXqgOWBfJVxITzs3J9Zo+
82nj7a7djcrTknpHFl9WPFtZoejTccYbIJ3usoU6VlASpx3zdT6D3ode1rL3sylN
OyFD0x69rQ1Udw81DbH8NLkxnlsvg7BB9U6b/lrUBTfyR2gmRGiQvfV9OpXVDE08
GKRvH9p0HnDOKAe5Od/E38wt0ZxSsQ1s61DYa7v1VnKhYcXNp1rHR5hTMH4bO9bo
UhQT0+HV+PbWRi3pIxSayQ1YIErWLjO5diEnvfMf9XKbwIbcQzNe4tttWt0LoTNz
zUvGJHpyEwJW2BEPpmdLoHRHbzooLTRjpXnIpouIQH7EOJVJbXdoD9FIC3pEORtM
I+oopI43Gh7rCmjgpv542bcKeetMrUrMdmzA3t76ZiSrK0Bq2gZ4Ktb29TyjCVEj
pMF82Nj16p6JcKK7JY+RfRPU/VWYvzn5aF5Rn2xmhBNsYhkARYCI4HflB/u+1Dz+
+QopB5vvO5PqXR7GBrpxflZwNP5nsd/37ilL8YjycT7fEui+oCSNXEiph6v0qG+I
npetQuLCsEcWdAchy7I3cgsqTlPVli4Jazi2szZR8Dc1+ri+RvClDqOaqhpjPeLH
i3ThBaNNOBKTiA6m3HvVj5jD2OeaphGw1IzTEh5Yw9NtQH5Fs2dVuWR2l5eaghSo
6JPcJHhRM0I9vp/zT6y5MTKxWkEQS+8hebv3K5A2jj/npWlkpm8BJ8tLmiWbUAvL
R+l/f/og3UxFpKQ5nFXXQeZwJGnSHCDxb2K6wUf6k365n5YEDY2/4ncN2PJ7XzT6
zGItN9BHWPPV4T+NFa2CW34lXhFlnhGU+wBbSQX1m+QCodBuMe1zSWKm1Gwt6Y3Z
Y2g+zn2AgQcTb7ZjMxU9bOoLffngy/rGYbB4cMrv8qHeAEIYNgckx8YUHLhULhKA
Ngq6jeSds7voeoRKsxYTebk8jN3C4BeIXATDgrwM8mlnPQaNe7bVHZ2oVy2Ap6yz
1NHmmHTdyeOE0gcqLapNhinUtBGM3iRcW7xVnLT00CgGXNPEs9ID8/naXEvCD/vu
nrzEd6g+Dj/x3Q2fZ9R8ElRS4yhuHD1fn+9CQXrqPqg5zE4BtAoa3c1eOiyyVzlZ
v5a1TuPPQqhLmxgju2Qr8ZGzJcQpfMzL8qV/ZB6kAPgQznFrsV1/TTgXO4N4GQvC
91DjG0nMzre+BWtru45hlhzZC5bekL+yoUwjDa0z/hzS7a7HjQwoOLu6McqQMnsG
Q+TNFbKjy3rFZ/2vMp/VHTzFZTdpJNFiCtuF5LrLr1NqWIV7fLT9dufSohQnZTon
gwl7KCutMtbTrQwj78K5ggGeHjANzWdrsYhcTJPN8i7Qov4Q8bwvW+V9OON6nQtU
zosrMd6girwl6QDsgGDyp75mHW/7hAhrMOLjO3SqqK9ErM8vizQDlFySCq46JRqg
uItEcrZpPOy/V+ZGIooKC385wTOsKDVipFtkQgKloGoQtBit1w75y2KSpSqZdqEc
ar9A7gDmNLrA8MoVMIwNaL5UYmMMQZab33wXtKT7fapo2aBG3q7rPW/CWvqPFh1S
ZbDiErbRjhsY8EpKYW+XS/kipEtE4hMNkrPS+rlnGomF5drBACrEaTYlymAWKJM6
fYBQPYS1H2zDycaPEJqZWhQ1BQRdrxNtaVRM7I1L9J2KNNXIlIu/Z6O8Ykh76AVP
q4RCnJF5nr5erXBc49vAjAUKGn9ToRffhPuPd1JeYalCog0nKdWts7y9litXB5a/
YRi5f1qK1h+y+n1vT97S+G+MHobtb+bYNbFUe3Je05453jlIlAgLBANMCPj5Cbdy
20CcNz/O9zHv7VRe+1X+a8/wwgl832T7mqYmm2SOAhKYhAMAp5mDDoZyZW87k1L7
PJ78qvSpSgNmcT+4ak4/LQUwJTMZs6TirmitV7oGXcu4HcYRc6YYZLrymHGxh8KL
gVHlaRGAxshCfeAz6EWCsLl6eXAc17mPf621GtHmRClOTlnCPCK+JL6ps2ELdXpV
ZuQtcXsJaWQlVQD6qrNI1WM76lvZ+mx4HE1gzO/nYvNPDXL4eVw9l9PSKxSLpjHU
GupGDCMbMiQuTI8eol1RIOE2IP37ijlh5k3QNolzZLgF97amFaEc/9Iq7XrVslTQ
retPydym9AKIonENZ8jrRGnEBbbikBjp5btEe9VAk2oGSHqG7JoaydfGjSWVPL7M
MgzyG/c6dAnhKB2US12Y4E23NRYLm9HotngD0GfMgWi9THh69B8Y6OTuUmtrvCBf
L+h10DBHYbqOwrlFN7tJ4nYX1hNfZqUxZZpO/6a4ovfGi5JoDl1kxKOXyKVGVTnp
9tveRACkIdsIXH3p8Tel6Nb3sLxvBjEnATqLVBYg23BukF5tmVtx4gWoKg+pbalq
8io0HjGKHhZ7GMXvF6bcBIRsIBdjq6Zt64SNsKhPEVrWzLch4QpZoogB5lt3ic7Y
AenBdoPV6Xwbt4evlFfInSLajauQtZmFF5SXRBljVVGuqW00r7TvG+/JJOkH8W69
dQdJXDr0PEFyZMmtXsE2Zczva7kTU7a7aisOR2aUUL1sujUpDnVTkowRpu77GdRT
0M9xC08LP6dyV6vlFvVtyifetJUkFZ2XSE/pFhPLAQdGC+xr8MTHvtjOpWRl9nFI
42vE6imQofzgwUqkG1MURo9wEgCGZ+V1hPq8W994aOyr8eZFog2mlWCSOQntjqS4
LiF/Y2H07s+Z2/F6kfQKbzd452Oe1nRRdclLIABiDl7Pdi4LehAhri38Aqabp4Qj
hCpAyjKySMKp0/nQN128VX9fK4Ue9dPGtjqdms0bNWhJhVySdF16Rzl+lb/ETyk4
CYZJwHwee9t/cFzhsqrF/Wu/+3jMdoPJOY5STXdn/aRHN1DcGB85XRT3+DFyGfHY
ahucsBIlM0WEhOSOBKkrtu4ea+ir5smo5iM04C8DcU0xDgTx/LBLO+GISR8fiC2z
9mrTyHogSOdaGBBZn1BbUX+QUTCvXwDPkImlxUAr6YXvaEeg2ZFrxS2vYkyGN1Yi
Rb53/8QS/c7lHSkYqBhCRV2APZ8+2OSgzGOipXvDYRvAP9w1SG+ZmbS7jBPA5Dck
5fA/Rd2hxk1fe/H0jdmKKq1ZlR5GAhtizjp0ZJfPL8zgJdl34yiLxHCP+f4T0cJy
M5UhM8phe0UcguOOoRGaDOq/Loqdo/BjIo8ozpRVZx5W9dq36u2hYHuaWwIizP9l
SbSvjFsswSWoqc6/IiIklvGml4ENRXeo8bEjqmGfRSRzg3WBrLwbf/Nwk1U4RLAX
AvQyziStjNed13QadnRmgAba0XNeSy/6L51eSBPi3MZDIr6gdFqsjOjIpshuWK6I
+R8KBOBdF4pc1sEP1LBAL6bfTlcZM8Grih7PnSEup3zR2ysV5e32fGcJyyc72BDs
/zmW2r7GImE/hWEMNaGnPW3oOAe08a0ulMeg3oae8ombUZatw1kI3cwpr/LptLEG
oiDBrnMTlFpdjb0jVVIoZUHUhSVoon+kBYIlNXV1i6HvJP6ZOl9umvQd77uDyXqC
xkwpgud+jpbRgNfDi01BKyNiVwqjjwqQHuz2zMrWa3usAxO0IJo8Is+d0Y9a12IA
sLJdWxOL+IJC5TVOmbc6m8I9io+q8WLwMy8UJuc7soGCrWyi3gcpb0pgmw0iOvgb
DkZzmpgV+UfkZ0HbfqFgVP66b2d+F9SSdWEhKBWAOA2vx1rjztWODzy5iF+Z4lbO
LlRtW0jiLCJVFMsL+lKjCSGkpJMJVyiBA4I6upN6joalQmJbPRrmBKOj/uwEL/Ne
Nljt5rWGmJ4/IiaGwXuwGCaJwep1Oy/m0CwdZl2sDFKZEKw+7RIOfAZgGimFJmHB
0PXBUsxiw+HoTPRewe1oCc3x8QcbnzKOszLi1h8aoxnqD41opj7yPRFpVPFQ311s
f7lP2DceO7mjTh9kPRxz7rx78woxREzm9JyCO/AqIs32jeeNNl5sxUQdlSNQ+N02
0nzdi9OjWY/msBbGl7H21rN6twAKpaTeaFk9rmElG0zzDbXAdpD3/QmBjuG+3fKi
ccLYK8yUMPlvtTIMHnz2JSJrylPhv2feHFsP/RrUY1RSspLg61NLZRV3eJS0/ruw
JSu5In5s+rlL4S8OBLQvynutY53jI0T8VZAp/gCbQIQSTWAmy6zZYlsizIpJ2aCG
Nb79YgDRhh54CKWNni+k2yY1s5A39/qZXi0wA37iDXYcgy1f4LVrfDWEodpKMMTa
U3IoEln8FR9M8qlrDQMnFKGbpt3q6DUVDr5uzg99nXdPcQySvmatSKA73RXtsY3V
7DWfgOS4urrMTdHmoZMrHMxWGoxZ9RWq12QFPlXpYDd38eUSSEwgAiSPoGhNw8i2
yDKH7dZDFFGhmM8oKUuQSyUXU6FOAq5H7AqqkUCbhX44MXDpOLUMq3anBoljibjP
p0Z1BcVbn+Kd4OTW1lkyxSxvYPu11DAyGS4rtgJdorPspgjZSaYuQ0pBRzOU+1Vv
x1xRiwtzyNvj+Con6gPZFVE5xQZVGh/k7Z3yzpjbWha1lGPqoBRnm0BUfcenvJvw
s992AFdgFgjDb56ooWu4Dr+WWkabrhLyF+yWTMmgVe1Ok+8Tdxqxz5Zw7AU3Cjfy
8kjUPi4iABek8U3lAS4hxv/1D1ERZOCq3vVOWkM+QWdIGzBHmXeAvMyiRaaLZiUs
1wMOXArc9cdFSsPQttcAphv0BMyZEUP0ZAKTK/JK1EXrocnYc84uS6GVNX9xS5Ur
b1xuePn+PwMZJ8rmciBmf8jgVqFhUQu8PZn9PIKlFGLdKLmzO6LbXf9MXNUwB4zi
d7cZUrN7V34JGYU1UNcljedLlJb8HuQ9DW3P+FFraXeXNaHLKq2blleVM4MiKZjL
CI9tcS5bl4tN7rYSWXndePizqnjTgdCdHQppL43ggsvQeM5Pt3eq3enT0xMdChSy
enRgBijjNRhdAfdwKZpDyd0jt/9JPT621d7zxbQur4d1EAxi07AnhEANr0SGSwh9
L0KzHVERv/1GCLIlLmCjoZUDY/Uu1NlEKTVHUToRh+njVnWmoyjNSoUgJvbVsSZn
oBpwgvDzwtAUND3ZpRppJtxmzDQi/DnJpA3FHmnk0ULZklRFbUI5eF+ADlbrrLCY
wSjzKM+VXC6pkLRCUQMMoigABm0GqeepDSBcpHBlS+CXz8IMeJ5oHZHjSHNy2NK1
RRxTNIba6gj72CEhlCUu43cRKRmf5cHxBGevQPsTpGYjdGEE11sdr4PkbT6VeYfd
D6chaayiJ1CSPWkDkkNcQeAg0Vxqc/8TxDkYBtlb8DnUpB0//cBGa2sTPFxtfCY6
Us4XZH7J1qwLLkibboY8BBcdnq3GCsDqREEuXRAoozJkJQzBMMfsmbMzLR574MLF
kBV+aRS7J0Nrq48+e49cnkAF5OmuGhhavXVkyGV7L9MvZmCW58vrsg52EStK6T+i
nnvEx8r7o4q+XxAMS4jHEPnsB0LQrvpcZs5xvrKG0T1w02zONl4f8+T3fTwJnFnA
yGXa16DB1Sc8Sn1/Tejrk9qI0eiDJ29pVAQiSgAf0loj0+ubkxR0tAKG8NvjA4sK
xuhPy3Sk+xJO2uHwV37nkk2y6x0paLGkzLNTyvZpz/GN0COknaQtBxZYDsVx8vi9
i4ENM1L3twjySC3vBgoZx/ne5yRHFbQD319u2xfjsOib71tRGqSIBt0TV++rQ4Vn
WLqdDlzGyhnA3v7PbPhza+VI+xO5rPJluOJX0wSZjmvbNNL/UK9rVs8EQA5/+4D0
WmrgTC6kdkzcwjcQPFDmw/AXAG+shzVdbJNJormksx7/oqwgWiWKrP3UOeoGoHFE
RPuTpPlf07yx6em0NXrVqn//4rWTFnFYVwfgnacdpbZO/CcYUAF8cNZz7fs6yJDh
QsJIGfL/ciZ8lza+pBSYwwq+cf1eOzfns9czJp7dUPSVLNxYG51ayZsYd7+gLDE3
aoQUKjPLsKTj43ZtQNqIdd8R4sNmCKT/6sciqlvmoeKir9Z94ppIywqayHv5JbWk
8PIYUlGE7uyYUmXgBKNZCPNz0BPjjSzHLas1LI7YuisohutE6WcM2nyezTeZ8Dqz
HoC4E3BFupM8yDcXDpLRj4nXCQjNU1Qox695PtRx/ZHH5p9AK0Xf2pZHbznkkUMr
GcUsZ+MMtivAHEYubilD6m6EqOBbaWl7xOwBTieBefFUcqFPZZqVRMrVUyLQ1rvg
TdMegeyfC8rWEIUVrc/jyVuh8tIoArYkyFZAPgYFFX6UPUDqTznGGzKDQATJkpEH
JsEKFGNn9dd4Va54Vb6PvzD1VPwYciX1Q/Iw69atqsiwb12XTA6zeRbjWtfBueVH
aZhM4eOfJ5hJzzzPjxOMrRMyffIAscF3aDqP/9QciJbPr/aVycvhK9KqCVSUtFhd
UNjQVTTs3X5nYoBa3JmtuRhpAWnPodbvzimQ2LkVp90xs54D/E8+MDAP+loz2Wj6
7KHar0xTTpluyojKVYXeKbOZ4lkNLnK6n7zll3uBFd/CDsn513tpI02jpeeNwtFf
JahAM5SIFEOsdzA96++eU2Un6FPfynYg3OELwNzzgPJu6ODeZWdQRIOlpyZ8qO2M
YQuWDd5xM59gPikYo+bTh7A4sh5aXTTZ0HJtp3BIsWO2AgQZgVWhAf7VKTwdhT1/
0MyokF/eoKvfhLmChW/lYwqZ4EJi1of39rW20ENG1jGy/Ekbx+jrZ7qqBA2gVtes
psnhRN/ab5wZOEuIjZGu6S6vUssWeHjoPGHURlKBtRH8G1k2UCqWXglhaoQFtpxH
jNZO2VAwtgRYJsishf7T+meJjFJnNFz71Kiv/Mld3w3p0z6DvETg8weFtT91qo8D
kzivzzJHAAf8jmoivhtA+qvM+TJbjrqTBkieJB3ZKUpWq8TfH6uY8xkr/tSv/4/t
VSZFW6Js8wD8Q9ypELJybw8nMIu5WiNQ0PL8zvocQdaR7D1n3lc1SQfNxZvZdTq8
oBgfiR1qbpA099wnKdCw1wtkXl5tVKqhn2OZ1sQJ9KwmwB6g6lWUZ+ZkvN5GthKg
Wwky4GiN5bqoBU+RkChM4eKdJg+WNAejVAc9x58KHQTOtelifzgf0++0aRm+FaNK
M58iESpDLIvt3RYSyA/yeaBv/O3p3NwyLSYyZeJfk9zrFOX20IHb4O8ehc2km9dJ
QhLdc+rCXyTEbXeFnsR0b+P1qAxNZUULn9rLGFXD/wN+8pyKskizM23GGIVdQLgf
n/rmxGLGEWghsY3DlfR8wTMjRMcNorNXd9qKkwF24/KE71GrMfL0ArHVEVSVu4/0
UY3OqneVMxknRm3FXTcxhaWSs+H9pSfA4lxoDdfTtKjt2USzeRIPMKq/LvTE4kEY
3n2Vacq+obct4lA/sFhyUzheoK6oPen6NqsOhlzAX70H6HrqFNkF3mgQsF/Q/83f
/fHE1XPyLlf7kEktnC9GBakvOwaqipjFc3rBRFFQmQ4HAOTfBdCsM4dAuTaWbLhH
NV91wlKZiLUeTTQOAiy8YeLrAp94c3aw6Di0vumq5S8D1ti2oFqVFe5dyhLkustJ
xr6xuJmW4frLhjpEGqKWxs1mUl/SXl2gTUIccNq4aEO6A5Ub0VT0Z/YDHZQzPmwp
57bUMAt3jJJzwq905IPEYwTCZpCHGF+ugfDLCVxu2WQRRjytSGvP+X5m70/JW5Q/
uy8Y/sF0mpQZYj09tnbDurRKObHhOnhG0AJ1pgg/vMpuJ8hfAqYehUXDmQA7F/ff
uZB61fV1KqMixdMMpbnIG4w+L0kORNBGSGHiDIqku7C+pFq4kl27KpUmA5GR2eTz
+uJ6E5ZmyTFtNhJvNJ2KtcZMtrUWL/LTdXjvg0PrppAiv5G5FDsp5rVhHouv41d3
RwLytI8+YeXhgkLyYihjxLBpTkQFWDI/TqtymXwUdt0e5VBwi68rE5L98E944Klf
Q2BDG4/Ab3UqcjG3jxdsBOXd58eNQRpjeoKM+IKOZ6HZSU0gfwGpnR1FR6IEgJk1
DgmmRM+7/OjfUNUyDipT2zRaiZKz71ml3dOXqAanuGlvzkhwSKssSX+iIDuOLFbl
FSpSjVIYayr1//H4NBWKNoxwXXy/5vUW0HVskLkgok3gfBBINACEReBjgWfg3xZX
GtOCmr9eEoNfP/WPBfmCPcVPkahhuetWbnDSnP3r6DRQflh13vqNxlWuTnpEC041
bjX6ZpOUCPoyd0Je67U20zLpq8k4rusoKwmy9+i2nO2lMwxGFKrNZCSjmb7EGfFD
/cWwIF+qiGAFp7dJb8MX6q0RyBw0movjnsIW8pq7Y6kO00+5TDLPWBAYduefUB3d
Apaq8/joe9DN9avUapOzORiGrqBkIXpKl1TL+u07PwfkAdslU8MbK7V8azMjidze
4NRMp/P9KG0+n8RPlVFC704lVlIs1tPEGKYIUh2y47PyH+mk+Pxx6ClXvtLGbLGv
oPTDgCqEFoM0/3XOPHwBPJ41i2FzDYzoNk9AnhXnG4BliaSoB70IVOYLNV6oOEIw
3Oe37E8nXXcHMQ7ZIHIK/URiSx7p3L5JiuKPN1iy6NryXTsiPLK6N6d6c9aHBNtK
4jXVXKOOrnuTDNAnfSkYUHood4NA8NSO5Wvf6ZHMtku/eXDo8XkOv/Zu8uxmNL2/
ozAgJqhVUpzpn9FJTp3OrMXZ5NwOOuOB6cFCxhSqvhmcabH1GpyMr8W4qF9zx4+u
Zq/DA0cxAr5yjNUsyW1SUoYLGU5qi2rJHpOdzJe5kvQ24uImC5+s+7PJcu9f44Ry
uBzf1rXDQeEvW6N7hb5Zg5EqfWnkf+atAtLyDQKGcChjrLEyFxVTjvzh3alBTPv5
rs4+4vQfm2vqh6hUKOdClxUmOy5o4kWmn0yJ9InsAUbanbCwxklw07DuZ9DEOEpu
lOcZiybrmQ72pJHY4e5B76/NjHFc4ao5F1enjJ9X2aP8XhUlMatvJn/oHsze1xUI
nj70a5Rfj6loISvXcUyuSGMrt8nIQC0zCg73wgHkdsvmJk8tjuE62TIRW/9y17Ib
z0qdevHGvsIFsYm4xAhuthnWD9LLA1qI6KsKOE4zQCO9KRywTet/jGG3OBwnXWAW
tZRxqFPQiaLuQntvRQx1k/ZhZznhK9j6Hh4m6V7nBoui5sJUoXa6nFEiApOCeD/l
DXPockwm+ljKEmjC1UnNQ9uCVlwJqtl8wJOqDkVFWECzVz3W5XEeNKGzKu1Ck27N
EW0JSQwb8U1z5hDi0YbfJk3dzJj1RfDy+htnaFeFH3KhGwivBGqZw2lUvQzYEaR1
Mlnym9Xby80rNUZKQBS1FoieArXYpf8FbuEZMhcIlGZwR7KOPIJuDvQeLSwrO+ku
aofzK31XnGBZdB7FX/sh7L7JkqYCTXS9MI6BRphQV3o5KB+qULHsiRhTE7Q7Qg9a
CqxufjZcTXSoYUuJPRqLiDSs81SiGmbBosPR9z2oKBw0wYk7hZ+WkVTvlqssUEai
iJZpp2TxCgRPRycWBXuDTSjWgyG1LfcXwu6E0vtaLIqCNvxSimcx7VmCtggm0fdJ
dOhvrKaoPW8cnhQU2LshkDAcj5bcSYAg0zs6Yx/RUszXbszOgECirpC5P+EVJgF6
VlxWKK8/KlZA48hrVZIe/d16qSnnA/1tDQ/1JLiLo0xikhqbVB3QTEm/wnh+RhmN
cNBfkfdeO7NCZHIIoih5AgEskPM34DEuheIVakA6/DBTE4dpz0+oAXadTTUY+9/W
ZqndQqNsB3Tv49qJKJKDf8nS9WbhwDVD1PKvDrufcEHTDno0V7HrZHuYQsxbcNr6
2QjJXle0L6LeoXxhu45yu7k9IgQRZTbl+eAb8KDgL8R6MGy9e0fBfxUjNJ31x6FC
2cU/txmNZG87SSex4XcfSd+EWnDkq0ihA65X5K4wdFHEsSknMKIvy0gdSH32F5pO
/QKtVQBpdnFwwPpvaNYBT/4mPkqOIFeqwsSkjiYE1hcZ709qeY7BkJrSh44YDLQG
ASdUclxijspwvn1NteTyn5jhicdECGbxBHl/0oiwhFHluat7Nkp6+3OdU3rN4g9c
TjWqf4Ed4MUdI0ZvPzUOnW9y0YrK6hLh+YzJfuAX474RvaErLyQWpquDxku+qdiM
OvaeGzHt+4HzXQGcE7aErlXNZK2RsR8vWeC9YBgjUrqPBQrOOtMhG73tP9nZzYJo
YdFBgmTfRzY2fAGRfBkHot3IroJc+jRUajWbI/W53tqblNTuIYDSDmSNzg160JKP
+LulBY3xDKYDiw1WerSEpGwDaUOa89QiVViF6wkyVKlrFGGK5v3keHDybvafmnHo
03WKdkxLJWLIC1mxOBVHRQUNHc6wTx85FKnfCcnRYs7rnGb/d8NV1lEAQ+wxfdjU
zmH5CZ7XHJWgcDk65123fCJhOyvqNvHF3gReMp71wXZ4Pwgtsk9m3P+yoFMgfQQm
2kJtZJtqBmFUwPGnZZC25WRJEgzLByP+J1fS5RTckgxIW9rmxGYiAt+pmIFp/FcY
7zamFiToErxkhVD3aP0M4WUwW7yNRlaObfr7At3Hh1yHKz5QfiniPYfDcEgGeo9x
BPJu+5UQamKRfcvDjBe29FgwbbPoRPMHxr6ZJE/w/A3NT8c9nqRxaYc97nA4I1aa
OltEj7XImz4PyASQGX/8NPyGLsz0tUL2PFn2+KGDWfIK3qS9cXJ4PM0PYQtFA8iR
G0SoVHyyCehe9j8iAWW5HbUIJXfcarOgQrbu9a6yR094VyD/jmJZcCdj8KH0QLSU
hkZ9DNA2Dd0IsnwbSXmeTGga2TrHKKo6FCcWQAbT2hBakwYn0ET78eJQUgkyGVj6
FymYs8aFvosalZAcyXT3EZpduXAB6BFB0gUGzAmttNfSKxlXxSxSlf7dXiKwYWxI
bzL12yEMcn2UP8hAnnyj2DbLGChp+4/wAPhmT7pmixhIl7hTU8Ip2DgJ7us/7cbS
H6s0cWLcJ7hMqVNDlVUjcqa6JXLINysaaOSsA0CknPqQ6Srnz7N3XzxfpB+7ZLOb
6ikouQ6SutctBbNeMx9eAHYLSyv7wQwv9Hh73g0tgYYKKjvQC1fbpHli0tlGyDSZ
a10ExubcXRiy14+hT1Habs1c8JfB0sv4XfV/0V9ascg7eDK1c0ljxCjFdaAwGefb
Tzj2ZaRq0OZ2HwXs10b80u03yQC3G6xsyZQ/o4LjnvS8iBaF7FVeITd8EdnMfUQV
qPtfh2Rs70dkdhcvTTbpja1y0u53Rqtrc/p4128KrJ13DwCfEtRJPOqjBnkV+Q/9
6x0oPdQ2g1HLW+xtNv4VfUhmBLX1neWtDh3AChQ3cUIo5YovvOwWUuC8odHJAsQd
tjRO2ihZQJPc1Eot+p43NHJvpNmUhqdFej3lsE4KJhHrXEyh8dj2PcycU4JORrSl
+KGvR47YKD4UruKuWfwvM/aemW1Puvqp9syNQkH+prOWk/8IeCXa1C+v57Zzu0a7
vVM8753h2tdY0h2Ca5NlWVRnuXtiORVVjEXxdyXUUfAw6bSADpztyEZxLUitzVc7
jzKDX+BlGsKhWPX3CHD97ZlvVsctMQPumAs7UqDWPrhw7vkoNQ98orDxZgWMX/Ae
DsPe0l3EuZSKW5QNP+0vjahouQvHGzSJuZoC6HPTqILc7CKqSeF3nUbq7V1l+1mb
F713GBllBE5C7SZKwZ50Ct56xoi4pdDrRQFJEY+B/NihMU0xQKlYz4M1x9iGurXw
JCb/3YIeCfs6P59yG0NdtcOwBE96a2yll54t6mtU+QA1rksJpmfUg/PE6izrn8qU
IhLdL/uTSnIhBkc1osnQpzewUbAAz/AjETaSBsRPwEcUM6VKnWxQ8yafWOJ971hb
K8Xxjyl4ceNgpiJTEkBBSFeWHrWOOokfoNZOHCEgTODRt9MkGpA7ieS4/0oL7eoR
Zt3IlGYw+B8M7NX34Dxe9PYgUvitzHa0Wn4+P7w8JnrgUJFmN6xN71Hc1X8c/B3I
XeOXvtxd6Az+WYVYdyAXziALqUtxCsZChliIxk8cd8clNYaXCkSka4hvgn4lIDqU
tHWOyz7G7HCshws7HoRMMCX60JLD7hpQEHvu1rXh702YxHjSo6WbfIMifob1FBW8
vQIoQi3sikf2OILmiSqfPzMWV3jP1fBvHvVOxV7sE8+IQ9ppR1UW9BkwihKN79Yf
ED3DPgOTKq3oUmCvElkxk5IIFIVxpVo6pL+DA9A2F4BuFIIApl2fBJQ18nQ4gUOg
QIO+lM8gAdOPD+Ll4kKa82I0sDsNU4ZfovXFVTOZPrB3V+B1+vbdtIiZuNNxYELL
d/VHIMzqPkVtrOmqh/nu0dnbuG6qjR9qXtH/yH9tZuyejWj787zdFegzzQQikiWM
ecuX3eKJBk27gzfq3teRxEed8ND3PQ2G9CLm5lqVNUmL1mel8ydW0sxIjVsjVp9Z
/aQ0N1tyMgNFtwzsFZeHRBNMqlwWqVFhV68LehidYao+oiR0g39HYXMki+UYG5dj
WNhRvIz8ZOvORO/MAMRE4G4YUR2qzRzLbOmxGoYwRQ0hV3wVCyV1mVkUMwUTZTiC
LGoEbSPHynY1xrLCbtmdfmpBruXngyYTqRiPbBwgt3xNKJwXJe9jmczJIOcPnk9c
YfHpeFmbpO0zyqh7SYqlUBwRCZWNV9NvPH6I7L9nUMW20HJkQuMFGjNS7WrDwWup
JVb3YIHkLXdSP2tGf7vZzl7W63NAglBwmq8GDwjiXEue0VcUmG6KZLQGeJJhewH8
KS5gpDHiR34hyxK78YVaWvL3XIJ3fO5SOP4VkgnKgbqZ5lqzO7MpxPC200EYLBsm
+zxr0/WxvraxtBQTGbb2fLAOhOcRcYy89kXbO0CtNu0HVGR7TrbgRfbn5RetiThi
3IPrgdvvxAQdgY9beEKpOD4DdaFVvv9gQyy6pouZSE144rX/NMTdC+uT9nq5KWsc
jz9PqeyAdQ5KOv7Ra8JWXYbFYvA5TcOnDdMvXBgDU7SFFWtlxrmEe3M0F9ZFDOy+
zVW7+8RdwVrk/JJizmbVKPPb/pWDljJHKuKF859u6kNrHANPz/A/TXy3RDhoY0dZ
WTuGCLsSZ8wTl6hd1oLGbGJ60CKH6p0LOeP57PpVxD32Gk1yMyzEOHdVTAwfIS3w
Rnvokbs7OjRXrt6zP/PZxjKyGmw3n5rtMYrAamA+eqXYuaBGzj5fDXGEcG7YwUZ4
Ortp8nz1BRXBwk7W9qVQID12tzBgLLtHn22wUjK+IQ90V8CUBEbjeBrYdoqYNq5a
npeTt7JL+nf6b5Ssc15DBcgUG0UMFESjjL38xVeXHfwIvCvtC1WtDH/ruuzvOToc
TAXuK3gHpMm+VKuIap2SiggqlLTH9axSeHmCZG/rTD0poehMiyySaUXVaTPRAclk
qxiopcLdAniWbb2LNZ2t10Sjtpak7nO+SKY2deiCU/kR9OxPihDfbAtOwmgaY74c
jPHi3NPsEOnUg6xTuWVB4bDIPYtUb2/1IUP5a1v//LsMtgpgFqAJWTH1masAeWSG
oyfl3cSEtwBKxr5KLi11vtQ+rXiCKCrLLiNX09GEWEYAjeVNs/pX/GFh0VAc33/Q
3pH3vS50Azw+DEBjrks5na5F+nvuboUOnDG4/hMUMa9EorBV9zyFJwBBPffG+GtB
2LM1B4psKcb7o89SdXHm6qyb3SKxBT5wEmMtesGO2RifMPvIQKJk4kZr1Nv64Y6o
mBOd/eiJo8DTV7l59uZhFmKOCvQK6yWu8yLLdIEW5hax0dkfIDKLgfpxzbLTFJ7m
oBDDo6xytnNxZTf8pyDtTaG++9b4RBfXKO4GRxx/ZwROZ34LS7GW7k+77DhWzxy4
TmcDrjNowNmqsVBFr9H9hL+dyhnEs1nlLctH5krBit508xSF6Hkw5xlQKyL7nVxP
6fMGOjidAFF7gTMJMnD7e0wqoHyJtdvpLbRyFaZT2BzxE6Q2BQOZQA3VPB1y1Yw6
Ne1nHEtGi+y6dXYcdUp76piL7pzjY6OxMTF4ZhXWGq1gcJ9oYtHnKfdWWajauFmY
yQ45xZ8lKK6UyqP2wDROO+zEnm6YMeImb78Q1A5yiXiqfgf2vG5wh4u862wNmho3
ZAyJT3s85GkjVT+T+sVRlqvQR072l+3zQdnx/9A5Aejw/k6q5u1M6OWru/yx0Jrc
thk3lxGVqfjtOTTq9gsCE6e9Bi8rOIrxz5uDs5IKkDosKQZCoe9k0yJ4nasjNvl2
c2hhHzWLtBjY+uZwB7Vtl97m7qUVoxmS7HG/GYOb1vrXUXBQ4V1SfEHAPNttNgvW
Rdry6VvFI2C3ywhn90E+aa8IlnInwovvtVyzOU5HraFlEh7IGlhNvZr/PJcaeJbQ
xuERWNHf/RlICl6HxG8Y3PN5ZeRTBBNWagiJdQKLMV91rSSADWDOE37AnktKoBzc
lCqGXNOE1+i8gZgnVlBl0GWvT4rOI5wDWLukKLF1yWmg6NZDPKlaMrWLL9Y06boC
7o3fn/UwcjVcIoU/gA1eSwhqz8u7iKZmaKorMCDYloa+emJ5Cb7cD0M3zqzn8SwX
xTU+INqWAp9/g2ig+jA/VFrfo54PzG00xIwSI5mWUoAqEPr+t5z83gy6KhElAhpd
r91kq7ca5ui/LIMvd0Dfw6peoGZjMbNfrm9ccB9xQa1tlJxHj/TRfczR0dtTZ8LD
76EU2MdwjnvOyCh62TUSVnp/iycRxg3l9bf5GMevbMzePBo0B+h25vz+taM2ZvW8
vyDfsT9J2LOnohoKh15wRYVgOpbs6x1HOnceFxytK8qst8E7Tuh4D5mmzwBmJogO
AKgDp69ohOftcHYSjaCEyegq7jxeCYEGSqPyce5HLe7AuO1jQY3u7xOJsiase+Uu
tRXhMHBs1/332abXIyQ3VEz0VuUhOXxF49jwXQe3t7dmK1I2wIb+eaaWjzT0Ev9r
8DWAnRo0PcVknbigTsbsGjST49aKbQxL/CwN7OwPBYJCHpDygC1h2m5FHOVjEfb3
j2gTO1hFP68AZl+xoDEizNyVE3kCBv+gPuQNaF7u7uYkS+46+EIkMht3xnm7UAIy
YJo4GxFgesxlzmkkX5OIHjo5Xo/pWyfOy34HmvzPBZCRJzKnXoQ6H4lquyHdRaAR
4K/E06N1dUquE3xphz9lp3LLRtj6VnmyTrdwkbLu2jiizYh82L/Iaip08FEjJMS0
wDv1X82wHxxBOOP5Dx9Cg8DRn5xOKthfHzsP5TiQthc4h3NDM6ftJDFxsx/3s51+
jue00PqUJKE3Es2/cksdyEEls86m5auir4o6H9N714vkHdvdUubkpUyYcrB6G/Y/
Mvu+1rsQku4M0dIrsKWng34dd+1ewcJALSzTcIcLI/2WUr6CnbnaUldC9LGcvJUV
Op4RR5xFOOyN0c693ARfkeOJQM+rI9+rUULy5J+dfNwGJhWFWo3YBUDr3/EEWAK2
0S8UJSFHwApIy9LpECOSzxFeSCFaWaH5aqWhSdfFHDTuIrcHLuk3BIA8OFFZIJ6N
+4FeU2mmFpE2XYV89N9tDXGq7jguLcMhJNzrxH0Fp7Ft5gBLgpgrIrApNOYjOlEg
kdcfm5+AAApew3aDPIao7weUbKltXWK+DKKNheVfSZH7ZHvE5jb52Xvgdnl3FSNB
vtT8IuFVLY/CAX2fbbp3Rps6UJLm++uxDzdkoWJ1YLh3a2zktJOAlbmUOV76hL3I
vh3KeWUfFeEVFOM/1LwhTcmWktr72l0qcRSyKbmCqa6NQMPHxg2+N0vfWCwCl+bg
mlmb6nlusn4NVtbGzJW2S0SQ5gOTSil65i0iw7DRoQgVWig0cOcKwTrn7wMRApGv
3zzZ0mGfgyxxHUHsG1AQ11atTFqhLMMapUgfe1gqc6Hs3Fz7nmgAKcbnKN9slCAx
uv33i9MBcVHDX1ykSWF91eiBQ3QCd4lwjmtocYHj76Yb65q7wm211E6gTPKfZ2Ib
y13Wv+r/sJBN2uJf/TCzEorxuY8ptyvAb56a4TnmwOmIdDRM0RAWUPge4ZaAdExC
njOYXZoWjNxTX8DKeb9KdO06CSmFi/IAgamUrXFoefoYUs18/g3u6CKE71SOKhIY
vo2p2VOdGCjCLCqHLsyifDOL9c3Tc0ug4emmUEb1coZK2dbCvqLlCnKPKAW8f+s7
eFhsKVUSsHoIBF5A4TxVStKbSjib3Bo1YjtpF3/2OeK/IbFSFmo8PeHrFvebwkCZ
fqWukAhAov2O5KdskAzgpZGWtqtc4z/LZRFrOps2VicUWh9cW+vFIcCm1+wzTrOS
kE/klAAHb/GjLwhIcDtPfbM3cSPvqlY2VHUCEnX93Ys0emeZLR/TRDEdP78Q8dyU
pQORDUk6iYZkgSnY1fj4OLnMOwQavXDQ/7rbc7V9svU3WyMuhh7qQacN802WQfJC
Ue6pdk3RI/5AlmSnuJxSzrF1+Mj12vjZN++nZ76rkF25vud1/Gk962geDt7yRkii
b3bFQO08HkBD9BcYoOlxLP7WBqg/Sg3ONUdhYZg8MXk9mW0ufVAoYZpNsCtpyTBz
d+RL4/1u/DcUTKy52pCUuZefXCAkOJF2t4jaPGRW+my+XdKdlPJ+820OuzjChmnL
WpuCc12f1oOc18D0pNxEl04l0PmVMaUZHOKyIXNH/sPN07cFACO7BBCxh5iZN/A4
cKygBeBSZLzOvVwZDVYgCNLqiw40rRrJ7StKbI8tebrTyPWUCW1hfRDLeqsArxzU
qpzIE4+L/pB1byL6t6E8+RX6PKNvJvSFtSRAA6WepqJHQwx0My4c1yQVdpnC7Eb2
GAjQPjNsJE/eRMv6MhEvopqKxlYMihvG49SxJa5zssO84/ohIzZSvPs/mP+RCJOO
FYfDw6ZYi9F1hjI1OXmPe9kmvBpTXPiWO3RKs79LIB4ewHO+s6zZxzXY0xCQ205U
AA5pZWiIch4YSk9tB+ElioMcmFfjK0t5ELdRWV6DguDLkl+CWptepiPOygYUZXva
4E7w4eT7K9+aH7np6QvOJKdykoljTz/ufOQu2EA3rwjRCN/bowHgF5NhjMTdeG3V
EsoTqVFRla5+0RRBu3vfRvUwviY2FKIHaO7yiHCxf783scpvQsRHVEKC2CKWzSWp
UzZL9tb6rsZ/5ckxuvH4J86k2es7rdGuiees1Qp/dxrl5A1BjTfJ0YMu8SPRKy2/
YJ/g7zivaKiQTzRLzb8Z94pjfusk7E61NN6FMRDgpPKUPwXccdD7P7zdsDaskBuT
OELySJNcIYDC3PRWjYP7WnSggbUzUlIQwsRwBaAXr8+YlOCrzIbGqrKYUyZ+8Y4c
NTNLuyQ0L/o2TJmMVUuQveAeSKFsrrLyR7D7xOuvQnuuvpq1y89jRxuxp0AaT239
k1I4A2bQPO/WKA2mPqKbHdpNtI2uKET+Ro12N2sKFEIxDg2aBf595s4W0uQPBnDA
q1f8MfYn7HwbcnUOMPrpCRHzKn0OwtjSXir2tGJ9mQEj4czRwm9D70B3GQecewWY
eabSKiim1X1eAhUaSSYdtqTbj++3mSG0AA1021vo8W38RG6GPps2GSVwhdAQBjVE
RPZv+pEWn0d34cG4UifWCjzPJjPw3Do2A4E64aNPzUSBcd9hwGd0QW+r7CrdxE7a
E1DPuxp3OY5BPwrZOBL1tGyPhAsIZpE8oGMD3LSzXa2wjAzPm/29DQfvHWi/YXAu
El/5FgySwUohvuW+asRLdivAa6wwSY+vaWzrt/m5VJZwPjX6lDYXfCOgPQpZDLH3
zavveotqIVGPzYRafqygcS3be/E8GoSuIY1fG/Se69eh6Z5tNxoFWnpOsujtaiD5
S+uIQ099vRm5RVP6zS5gX+Ydvu91V6ScQK4kc8xDQNmvllfaUWnnIpbkxFtfmbqu
zoWljD/rvjhNhpO2JTbSWlKoeOOK9NMqwnu4aXK5hbJMFFB2/3wwCkUkzfco99AE
4cEtc6ozhMRSyDDexmn/XZ0KK4z4oCswxejWh4tAYFHmsFfM9ub6sBilbG957QnK
I+5N1iSXznTKU4PncUZxg7M1vR9qak8PN1R+zrTJ2VULArZQ3saTS85awhsjPJOi
wJyBzJDJhRV+gsTzDXwP661AxEIXSq7UTUXeP9kBbXOBaONEW1nn6Y4Ha3yH7uKh
FKhePu++waZLv2imsaHn2S4EVgJn6YNvJ/xiaS5oZvsrp5rfYwPLmYh6mqQdUpD1
N2An+M7QgFvBbYgXXq4B5R7WeTg/PU2AFXLxvjk2HvenrmPGKTN4id7e5/rDtfu5
MV/QfhE2tD3jxuoF6++I6cNxH3A6P+lOuViLR1/SdWKSoi5/Jl1J/8yB3lYZajeK
7WiP/lAGA+D02k8sa34KY4rs6MN7p28G5yWmnGdhNh+yyfcKVo7XtPxI42If9H5x
P98ExkeSUDFqOFgemgh+5Bx2NmjWyT9IRzcdDcNjgManLaK72jXYuutaoGOkA3cK
DMEIAtgG7WSe8NYzGnBEKrEBaPoTemCYOLo1EEyw5vwv6vfEt41FZPD1TcrNxJ+R
6zl+imOahbibNt07Xki6E7HMXK96nV6Gt89aCWKE2GXFqt7o+PD1/Yfpd/8mdVTh
O4VIHzaaHo6HGrzIa+jACqvrRc1XxwhCW0/IjAmhX52rdxS+V/Lp1tAfBt/k4lgd
aYd8eovVDSKGCPva+pJ5HOZzNRZoR1ltqE/bXT5gtj5HU+eYuOpmO/2+3jvXGTth
+jp6oGBMeB2zODMzfSuv8TrWxEW5OS8bJO+j4E7Qc6OI95RqYzIDiV9Y6ADfOSMh
zaSX5Pp+VUUTAlakdRDeQ7Xqasc7inwLwwf5FO7B0t51D7ESQjU/Vj+NNhAW+aY0
uMosG9hNudJempSHZNNq/HU5UMkZavcu5JttuOTgc8kX+NdieatnMEfuKpKjnsrp
Yz4h2tW22NNNDleGaa8iPPSJM4nV99mHIcEl/yUCXtkAxAALLkHa/e3ZiBE3y68J
hbnS/eZEV6cEjww8JJdmSeC6+Bsz9Dkjj7LrVETBylzMoSFcp7KrwDS3K5wS8xQH
wlN+HYaEVHB0ch7/jrBrqSlRsGslOExcTgjUF0X4W9tZkPfEiaBJpq1WBxXCvzh7
Vy+3jlrO2oa7ORbO1mg40oGnLEsEECPLCvGjADPAovKMCDnKJcPtBAZCboJXqA6u
UCL5+EocVJd8IMs0hGCyhCMxyIsA7+wQ3TarrSHbDFf6byJrcqrf3LfBRv4Et9LM
9y9I19dpY+suDaP6xfKtALuGCnTyRAvqalJQWmh4Yi6VBQZKYDiaFf/iTYh15vxF
oCZ/lvx02Ev3wWDJ4ReXEJthNC85woqJ4PRTczjgS5kzqCJ5vo6ieyYORF2lc+ii
U2bSTmmZpPZuvOrOdlZEjVgfOlEmnlYzy+1kK8Z65BAp313VFvwSLWvTb9Iwommi
JAuAH3wi7qXdcT2MLgMuycfkfpz8PvJP0MQZNgilCAN/fQjzrxeGc+mV5mfGwgQ8
Fhem7hCfbu2312tX2lnom2mb6IsXQI5CmBqznD8veLsTntbKWHDILp+HH25LIjGV
8GufO2+5oE3qiuu1gPrSuyvWCYseB5NXwBmzzPr4dKVm5SZUt7/f8F77mXfyOFvI
kktU9krZpgEDV5/Noy2MG1xjyOonzFCBUgRyccQwLxIiJ8IQir4kbTQNtkQu/MQx
DWHQw3LZQShNwe6NS0eV+dY95bvgX/x5fKZNHHzMhNko6EixbiS7gjNuNgbs9zEX
4WhjbLCjWhezwWl7orVNNNaaCPFRW5jm4AJd2wIzFEFdCWoHadEIOIUDaXhU6uIt
NgBdUJQcCPYs9W1Vl6T3idxr2N0AzTjcjF/Dgle9jL5cGy8zbMFfKu3npcEuJUKE
31ys/Hg/PGRUHB2A8Gv3nISGsyBMGcMHCxDaxNEJVILnIipIA1toP44CgaqxRTBV
wGjx9SIdAELDU214xFCRIcJc43Vav5CP79v4xX+5CGNYunF5numkC4OsYBkE6f43
yLnU6fMbid+FncJI+X9W1CCc4T/SR5zhovCyjnVywUwlxhUeVcTh4zhks+VHZxpk
rDJPBTg9SSNh4+geKxcZTVGUr9aUPuxvvOxdKOH9mD0Yupc1hO/D2/iGOd+LAbgS
B6ye+8f6zvWzgDFuKcC8ETxToCCFrSy4w9DzUQ2SFqfwcbHC0EVfNNRUVYLzj9Q8
TR7ZfYZbz6MtnQxKZME0QNPtmICMHKFy+2+HZDICMAavBk0SpDCwW4RUpzWwyzfW
hUi+O+jLRhTql64vxBKZOBG3skCd13AMof5VOE4i1spvFCZijJn3b6qW6R0KDGHW
rGzzPNe6w4aE+4KaQJn9tLJQJjNOGh03gOwe54s6fTDh0G0Ww+FBTayom5fL+eSl
5iniNVr/HfSRRnJ2R7DJokKVLiIFUa4DIxs0JWu77zDVQiBTinTvYh4g+exDKVZQ
iOX4MvbG3mSHRK9O7dFQrRM0SmDV+GUHTJ1n0NtSiHokyndgETfU6wLYkSnPsuP6
LVfJCr7b1QdjC/P/NvSAFm/D1uusZd2g/fP1K7WGVUAfwsy4yNNDQdm34YrqV3VC
V14CBkz1dra01HlGCingHe0LgOhOiK0YQOdptEleeh1nSKduq829fpH0YLOzCVu8
6XDx2az+cUwOzWvoTUjCClYRjM1d+g0qgPUiaUZOjlKyOHZkS1fhILun3kpEcxij
ZNY0qSdQAat5W56Ux2/IftuJwHH5rpNeZ9o2Ok5JGVtNgvRSY1Tz8zu6G+wqEIk/
E0cTtXe4jzuADqEIOuiH+HZXeTIujZnjs/IWWcKERanQJWhKeXiPuoXDW4BXzpMA
Ax+rJx+sEcnDkEG+RWjJPpIBHNWBhLftq35TN9tEPDJNrSlqsGO+wSWNP4k0DI0U
+iUb1IKrkYTKdmPhSIzR5KoGWiyJCinAfaXOSZEbOyxavsGXLTLrYEUGPuUJsgvw
Eebwi65/ZJFzzC9G4ThqPO2uTXOzwYl7uEgrepcycIYf9Lxi7f2FlAQ5m0ggvRUP
vHFrL4ZWJ2ygUIYUe/oFoGnv3nJx0m+33lTiaQDXizLYjdEq0CoeEHCgl717qyTV
6EJUiFPDS8acexDCjK5FjfpckiCGjMNJlYeNjrv0Dvyg+5YC1OCPtjgn5G9Viko9
sc3yVQYIlo/7T9lM+gZ2gXKig/fzcE5Ecy16SzOelHcHRObhF1KkbZ1+KYAsF5f+
hl4bbTVlPUEVdspUuqA+JGDfHOQ56WhWZuV/7UnLA/quXhLvaTHp2DQMb1trffXF
HYPENFhCRhF/Qn6qiKyzOtlvr57QEn7TYjVI9sAnw6kDNGiVH0pT3urxIihgCj6H
5HNytOZlwDmJXkUTlnUkFt7xE9iWB+SN90aY/w1DQNOyWO+KqHx2PDK3H5loYZRL
K12lFNau0f1eTwz7bVMLlXk3w3sWurqENrQR+nr1+KkidKhLZXuhigVbV1ujsXCE
ysGztUeNilhNCjsj62a9DoaYYVo6Te4fqFhdlnDNQumFdr8s/hFWf8NWJwfPrDML
bgeuA2H/00f7hcY+ImPTy09ON3tIMH9SeNg5KFomV5ylWXoY3YM2TlHW4Udo1ufg
bbCxcI3E59ue0g01wre7TpbiKJGjqaFLsvAyaJvwCLaRXM0cFarhwU7xlOiMHZNx
ehYvSKR4tEx7BgwhRq3PAo3WjvtPj+1rZah2K7CkpCnA59x6EblSeKt6YCGrlnxr
0hcgCTHC7EMqWq//RKyzqzCb9yD5rmSABQqgfC9Fbu/9mreXz6PFNEZSYIfj2SzJ
RFy3m0FrRg0sPlB7icGNsbJPBirJjYUZZuKku+tH5eM/f6Q1Dp/fNxBLots6i6AX
1NON3NDugys+NNI3QbA3ntUdBSlPSND7TK6gEze/Uaa+DVGdoJfhLbAphkyCqBk6
ykg3AVqUjmhyaBw9SHN35cgF5hja7mVDOuC7JG816ZEyYxWA7YzUM78NuSObWc+R
8LfUgfBjqJ//2KtvHeG79xwpPL78VSIv4Q9znngXWSzn21eCQ7FwM7Fw88QctHuc
+RUt4toRSvW+if2bpvsyn105vaw12OQ+GUCqlxj5SOucvBl7U2TeqshAH/OjvA0A
IJiN9bEfeZzl25aRDsjLgafN9m1FhjHC8VCukWmUyTtIvTIeJLizOISyWyIEpjmy
KZehiH8eGTvqRQzPkX+qF71yeso35U8rRQzDbFenYpL4iALDjELZQmLj2jK+3SMA
T+W9uIaqeTb04CJzz6N/DQiKcJnccLgxsqs2EqhDLJccCW4UGwhjtQQQbqH7tjf8
Yc88Qig0RTzwTeJsaDCIPJ3SX9Uwhso6KHKFzKXltFfAkiA74W1nSKygtqjEOomC
8rYDtilfGG5/4jKqErwW6smIPF4ZvUvFdOHMBrcaOqx/LHLWhVF0w9l+IZej49KT
mNQq0IdpzhjZp2bDI8eyZr6jUkVqTDDkaKTnO94C2bpRu6vJ57r78YBGkIAfQ1u5
Ce2SoSdf7r5UoeXivBUxShKskxUDT7jrMZrhLruMxfVan6n5yy1FtK+9jCwQOizG
wvsCjKhn2ceoMbSiXtnu+2AUzhNZHOv05OF2mo2jsaeYYPOGzw743A2D6Ht1xwjk
TQBhEBq10sZYfkHIKEv/10vOlVl8R8fGOtVviZuSTKi7VYAKMn+BTHm1t8KGJurR
e4CKmy8JGML4wHMX05NxnNFt5/+XPnoaJNmAPmcd0mszeqWy4emP+hucn2jDOcvH
112MFQ3U2NTRzXezXpbMPRgpzih4z/6Kc5r2CWROs0H7lM5AF0tPLELHvZQETR5O
rcwjMQgJhtoKRBTfCRulApkDhlUnDFywla1hMZGZ0Jqu7e2irUaI0Chv1nXvnQ5a
PhvsXiQowpoyVDU2pQWvWJDdv/p4U2fil+RlQFI2FTtCA54Ryruc+nE0LHo5x0hP
ztiUTNZPI40qxDtXVU+CMTCxUsj0mpxH/IXX+uiPaq5ZtttPj/Q1QNJS316FJ9pI
kEBpHOCMWrWDhZvKDFj2ta6YsIPQtApTARNzUDqx67caa54x8YnMcnk0y06q0oC5
/+KcXd/SDN9LvEB+IPGhcfHIqzDJLmvJPY2eaIGR63Nq8lMf+7uBYVN3bSrMnVJA
sFlrn9B4Ca/68niAcM0FzzvU86/xv1NZWe5Ft4j0HWPvx8iwRqwLsRZSr/YTaQF9
xA/PbwKQkVn8U/2wXoM0ZpKz/aM1oxgcxEtlNcaiP7Pc6JhE1CvXVFLNDP4SFxJF
m9cmFUcfdW8qPXwj7S0o2RF/8MejgcIaNjvirO3Q572wRsFObPWAYYEmNsu5vmIe
vnkmM2fRJlHJdld6dX5oQ6UryxrfM4g62qd+CpXkj4pEzZEWSKdN97xOIctTFhWZ
9KryFrDX45+BKf5Bn097VpCzhtK+haKkHRGMDBeG+uJGt6AY0aDfVCAaK+aVhZNn
efHb/QYRb+IRDc7N5uu6xGd+PhrEUk7bjfUPuZKTcU1SXYX42im3RvoPSSz4vO+H
iVDro2QX5y4RrdJdFYoX6wck0tQkqz4fHlP8vtHcRufOhm2KwiaBHfBd8oU8hhbm
oUCJp4fsw4IyyRTyE/sghP/wUEU4T7xUX0y/8LUiCMFI1XdM61YZSBBisuTJo3ws
k9xbK/yToY7wuuPGPmuSjC6tybf0JCYK5G8hifbWUphAvfIeTc+0dvDxySldaDxg
PUSftOprWpIFCu3V16KiyZ8Lvuc9lBoVQG/Qm9MU+rMyc5jtAJilxxCvI2SorPFm
/lxOWItiMX33yCk//nWwfWssS0H7Y7YNQVnftpJ2hId2CcnG3ex1qR8AAVsLlC1p
ZHNoxNfHggkjxTXiNK6nMPaT7yXYRs5PpUrwx5IgFsMq5pzc6bfsYboZWgN41ifj
H2YIqSbnj5pRMhsZ5OR2kAdqpxtssv9tkcHfn9tOfy+Crtkj2WjMvLrOkM1FZ62t
EHnbguumcJSpo69ykCt+MZK6/H9ea+oP0bTRJwfbiGto35VohF4vObUsU5Vy2WF9
oqbvzyqJKQ44oDPvuarjBBrE9wo2PyhJjYSFDGr8L7/tyD3C61wep/jlAN7zTpRi
ZfrG6Pa05JDdYSVPB0fJdxwvJtPhHkFD3AO7b0Cjgw94b1hu/SQosaYX98nUeX4f
GJtCZDE07TpFMx9Y1tm902rxqWi2hBDLLtbtkr4HbACvWzn4NPBZj/yzHbfUiHfg
lItdwQxlZe+Pu1OQ3Zp/H6hvbfxFmtU2lWWdU90E6GDZ2YDRII+2N0vXqdGhMrwW
26PcVLloqVhCTRHwyoFdN0bYgvPbRFDM7Ot0s3pGZWzgUq37C0WLhCwUNCQFox1t
sJ2OzB84QePNp/0fQiEIMOUPO4P3L7E39/vxjC3TMujovhcx+qSc2O5o9/HzLKnQ
7oWTm88zOE5NRENoO3qV+D2TPe2P42ojUHat6Mapc1KXqlcMSLk7pwPauoFw0Qxm
U2B4qVW7exFnfBNJQYQ4azBZLpsD0L88LQII7N1GHjUdUe7LUQ3KarU6YE4Kyz91
e3iegRuWhiN2xYVcDP6wb4InWeVRQX6KCR2VvEgJRAQ+3bZNYv7gvx5xEHLh8k3K
V+qKFKfBDMCNV+lVmidbDN/nQpOR4dVzR/QdKdVVXq/Uit0yBOTmtGVkvWgrzn2L
1voo66xjxnNpsU3okfUrz1rBWD0EwrVcu9ExGT/3kU/5QILN7/L6w6WVReg262VF
xCxBMMgvlnce0dI0dd7gqVMx657WRLeQlfXMr4LgaFGd2ey/9VMRFocIB6TROFAL
8jrHs0g1c2H1jLTMAzYF8HF/j1DNeVbeSdeWbq+6WDViLGdaHkqViL5FYVNTxHQw
Y0Lnv0XI9yjW3lojVM867E+yH0PlgXIDnkf7+ZDyri8fLlrrdNFY0lbJ4uBJWVY5
oxKi6VN27NEA6BtI1KH7dmSEx6fZPJo7kGh9QEGs85o4I2W/IXD7otRT2FwGVpyn
Eb/07YrEplFusmdGmdJtlOMc+59an2jOPHjnd4LiyBYst4UHFgjWS9C5J9D2bx3f
QHH5zDus4llR3+M+4c/EB6IIBy7pGHDmq/sKMwCBbgU1TlCttrTQa2qyJJxVf8/K
0UbvY0Nc456J/XiO4S/DQHgk5hXkvjui1tWlIP1QsWW1qfpo3x4DGoU3EJY/Z0LJ
pZ7yUHsO9jZrhE73+seqM3c+TD4RKUBwvEzSXKZWS+B/Au1FWb7iqbsJq6gBS2cC
mXCZdYTzr6uRyGwHIucugsvkdT6hfoSQmKqhfTogt6x2AySclWtapvkxhf8zowpt
L6x9xcBb3pRJMmqlzFFSov6yekFrpITt+FrL7CtQMINDtGX7yssbLxgreF3TIyc4
yD3vmCoifsgT5+0F0TdXEMWUJcjrYuDez7A6Vb9RdmRwtQX/Nr1z7voppeTMPqAZ
FflarMMv2fDBTgYeK8jqwPNIsbPRd+tIHh6+vUE9SwTk7twKkTDyL3UcXOxd6GcL
W5WJHu5vvejt72OhXOMV66Jzy40sWbGfLceAuQZksU4s/lbfwEa1T81AdlTuOpxh
hUkc8PWoeq0vDoBZeNnZ/uEoikEEI3rGSIQUcMTb3c2ZqeCHI4bmK2W3pYh6nXm2
lS8uo4PoYqqLkx8xtElVqblQzwBk2CMVESy8CgSGBTRxu+B2OiryI5Y2xgbmnGy/
q0ttbppB9O56nGbp+ipVQ8Pyns2sVkUZupcEX4Uo+1eLOQnTGsh/WdZMF2lU7xg1
aNwENejzgzuFx1qzwjYJfsKwfeQfqgGTPsEDge+cp71MwLvqNlRQUfZGDxnnitT+
ai4cXtOMZTmCo0htQe8yJkNjh+huMEgQoPxZWr5WLjU8wWcC1Fon78dpddY9aPvZ
bo7QC3ESLkUNAkuh4GEcBnlcnWUJpI7NR1IpoBReeayDHzCUY64A5xzVJrE0bIa0
GOCb0Dqx6kJevhscDyYz5lavec5ihAEWUmyKWXFbvE2W0EGn5jGOqmNsixGB59t5
bKbhs9erOKNzaqp3VMFY+IKoXGtzHHTLzzG9uS/xof5FkYyqJwL07ljG411evS7f
niuSkcuHgDbQplHl99pfjcbKDjnnDkgmH9XwYSMHWABR6lnuzFN195x7ptoJblaX
iUanHjZG2ojTCU5BFN9t468MeOEh9/LP9p20HnZ5F6z0V8Jxap3rqoE6jKPFpbvv
594wPWB152YL0Kdr3yAslaDF0uIujUMa5c9iXeCB/v6ciIvchd8bY9wxgPmmrIOA
R2BuPCqVTH44lmqQRX/CI5ZrWMLGLvdD5EcbvePIGJwjRUi9v5V1DoiNHVZrURXO
k/yXseGEA2e9YP6T9qX7PwVdfNbEhepFMsCZOU37ml0MSYT3bXHJXrSxVcGJTjIa
AvkzRyym7+TnhbNaRLDpvFBA1jW/cJrmK5q8GRGDkLZhWC67EXo2IfmGohBlm3bQ
w6UKwEBTJFFhT4tOk2313lO7UX1xRrecU5m5m8bemLuMRmVOG4rtmLTqbN+Nzphj
LI0As95sV3z9EhYAyH1mwMupERwFeMIF1ssxq7vzcFBOcERttNRhRR1KWagXsq94
CkHtOKOsEiul3fh6PhDwRjIgWd5+J5FNCTqTXqfyLeEiV+sn9BTPGqP+A2pujE4t
z1Le23gk8zCXhKVny7ICCFde77nur9RukLbgaguikQC8jrQQiImXuqSnIQYc4DKK
vB5brdNSmLPXRawulX1OFqhnxK8BM0EKjbKbTN/hoT0r9B7/H0e6lNirt4aRVCqB
OlMBCkmUS1/KCkpGJBryU40MxaOd7mYjbFxqAtpq93Kcvxsnk8cJnBWwAbkP5wXz
pcFru3KcBNoNzTVpUBgEA7yEkNWEOJxCjK5qgv/a8tGXxa9cfjhlKmphfqtsLUx+
l4ObY+cgwUAinwJEnSebTBzE/7Tw0owhen9+HwCjWuAxHhFtz0c24ZP5JIPjE7yE
ZuGu9c+6qtgEi0E0WkCcjobPEtCITDZ4Fy4gpLaiue2hF7EcDXwYfQBdzohjB1No
j8saV70oh+yM7NCgqy7uA6bgJzPSrjLCBh5+geYygKrc3PdgLgkTFHbyFkP0dicJ
ba6iqitQIGF0Hse8szvxZsLLGn4NbR+ZoqseBsecCbpx5juUSB8Fl5Cc8bDzUho/
ABIv+TfSudD5UcjBfZSyM6sKo7zBkVu52CQcfNKZBM46rzG+p3e+o+qm2Up20N/2
UcaEkcvHD0sNEHZfUT6PDKuPP30e/I86Gm/w3xJYHJwnl528Dt0HAUBm9/5D87c0
YISy9Vhp7FkzWaMDU+IJVBmG4wG6OrVwjUkOWKgfDmQ8F3zINsllMtuEsrdzC50P
Epe0WGrHWz0Z4EU1abh+j/8EQ6KY4ITgRgKDRAMBGFEm9LwPyzMSyllPzxSjpXuE
rxb1lnDlfgzzMNVc/uvDCm8qtLVaV8gXq03t8I/Ehmb/+Oj+sCHqgajBJVUBRXqC
cbmnAmoM7Kyms3EgW7o0WHcGj32Do30xT0hVRDr892/ouFdbCfIlbbRLhWBG8BAO
6b7cS+6ruT+okfDxJc3Vhvhk0hxebPjTLiRjU/+8DuyAok0nhxGTVyKQKUPiRTqv
1622ethoZDyQXMUJY2roysLuewqNPxNAcR7MeRmK9DzR57Zn0Lb67VFfn0i4RYG1
TXm8quEWTwXYXlYC3v2HGIAapNPSNDa0VXjBIkJaXGmt5XIEL3F4G6F2VkochcRG
u/DI2NP4pAYGVst5AhPUMgR9mr0dUXHf2Yf4uHaiFmQOPymsDL3mhJuclyfmZUdr
oe4yLbRPI9OgEtEYFBNd/hGoOE12MU/pSoPz4kMkT3Ok0mfh1u+5iepj6bDZs02I
08ViDt1SeTZo/72u/BMP3bkrnHIvK6YVWKa52iue9wia+wEQut1pRIqhVeI1ukPr
O4HwmTbYGlg14KN1QsWfNDrvfhrwJy2b3Pe6STXaVCzildNEEuNLYqPLzjfi2T44
3GvT1jcY9OV0N725ZhbLaNNg9oP7T4upLjd4AjB5ItbvUnDT5hY7F1xjLXWZWo8D
vnIZRN+D/xOnlKnZq3qAoONDHqXum13lVjKLDo/JIm3lIuLNk5MHfYsfZxXOaRmr
FxzmGkJjn6Di+zTpghrKwCaQJs/jm6cSZCrHUTOSYC+yp7AU+4mabLFZ9IP5aYrv
4vC5K5Z7xqkDIsZGtaZ6nGOkfVHnqvEsomYZBlGCeXskQIEpMakjNU6eMAs8AR5g
1eri0bvYD2Si4XTTF3CvLSB8v3R7o643NAb2jL2AHCz9MctJzXXXNauSabCuBwli
63DkfRnwdw85qbeCDnxr+Ka+GYTOE+NXLI19bnX1AZWpGSqwX6tqaQWlc96Rzsg1
ohEopE0jAhxkCzdyTcTIgP3htLQdYChgJuIxB2O6eUKyO84r2Vx4CbsvhUw7P0t5
JDTPbbXwu3d8eOdkeVDluP7cKR5hOFm8w70tETcKrjHNILZOw1oiC8v3rt3+PEl+
UNTUHphO/U1mx0nYiQ6yR5VO7NbFRiQaHYwp8G88635CSQgjL8KYHcpQoB0k88QE
FUeaObBuwaBt2WfKjYSunvU9EIXe/2d9vNDHqxwoC7tGbjxjjdnfe/u1kibVuNPI
MbOhj1/mwg4oft5XEImJaBFz/M5B5H1oOGm0jqcMyOQ5vYxIpd1ob33ABULxm0fA
SPrygcla26JLcgXFBF1R9GH6UWIXOZ7xnM9uNAB7+cyjuiDyy3jQwGcUHOKeDI+u
RfvDXMuXRv8A0hqqWFJ5wrG0zdDA4Ej5ivGtsDW3VYICF/77ukPXIytw1S6HBUL1
dqsUcEYIvI5vN20OzvcxeJDZC9zmeYxj4dv/EZvQgqLHXYyBxenwCBYSr747QZeY
ksGpgA4u1EkFxv30A0GJ8bim3ilOuv8hurdOMjftaX8Q113xwXLibBZqEdtfalr0
gTnjCJfmkXNtqao6HiZxoOIOLbWdzPbKUuMSBLznr+fOc0dJw5LaajfHKzpSCOmq
zpvK4E7WgO02NQgIv/wG9sUxQhYj9eRZspKkO5V/HXOmwbJ5hvAtbU+CTqKE0XJI
9zb7zNyDUeCDzCGLgfJvX0htgnod5BuiXew71exT3Vc0gitri9BrfEqzihirA68W
/iF0gTpK+Q8jwNnhgUXgAHSZNZPFCwkWshu11QqjEQjsdPVBWoovWc9Ihoe9rb8p
mYC0Hkw7M040Y4pNuotyXuv5e/feGWUM8T0i+8UNCwlwhZeqkZ2TOCWWFQhAc9bY
APFBaFcVUa3310+74nYKh/lvB2/XNGMIyj7MHpJN07qxBmWqC0xCno25/WtU4my1
nUq3Z87Zn9sXAeRQHOnRr1yrtoC04IbQkyGr+M7C8ObrmeqqhPQBCVUD2bEp8Lgk
poEgn/nLng0LwaWZ2lv0piC0NPsj6TY4Q5pfCHi+l57f6Y3bpJIBXQ5FhJuTbPc7
yga0gjO6Wpywdf5FzT+IwVUpIGzKHvAz8HpjLb+6gPX1gYwdowItz2cvZ+iy6IYa
BTTLMbbE0irCc/U8s1F2zCqDJrFU6rISv4Cwn+NSR3QCSftqJp599+v19JwFiEXD
J/eoj8dFPJji1CFJOQaxyk5mpdzcxFad/pyhtT3ZFuGf5hLK9pFRnoi5OJjPcEIz
7pGIelXhaOOVTJwQwyStAZFoHCvqDilkcfXvY69qG8UDuWxGBu0h0r34vhbK0uJd
pbm8gXwyCO1YtDQffivlofcpAcnCBIZjIh/nmA1Y7/txZUCFT24xUChx7iwEUjIQ
+5dB6X5mlkxAApBDvB8U6rwCLOVtSR62wWEJzxhXG+nsNEohI9F7gwcXxczygUhG
vqAJPMlenO2MRUuXVvp44HdyBeIT0Bj1uwkn7RuJiXziFEpWLjZBRhVacaZnBm17
/wMn926/BGuRS+IjgtyZ7T0jdvr8/j/WZjGHk03pRBcqtF570w+zIkUM2hSbFfmA
LXFSiIj/u/YLKE2QpoVWfOnPlhWPGjxC+7QfDoKvRORQyElm1X5K/FLuHlJi/m0H
kGUC/LKRvWuGtaoxurqXrLxtExReDYJKvMJQTt3ejf+sPLmBdjti2y2NQ59Pcp79
6SAUP6skn1oeahF/+V+QNzbPl1FJtkN6urFuniK0z7SI9fFah/aMyJpgqt7iE9jT
5TGVlBg6olrBn+eCTdiLm2z+ULhq91PDTgWO/L8j2a2yiK+Zk6ucjM0+6Ir/2t7s
sSVDDeBOkmgTEM5vJCEAmuOe+hP47pfPl/IKnq38fbSbHXkXuO0kPyHK0dLWMvnz
NTdYtggEP2+Y62AA9c93e1Yj399zoR6xJLJ1/8iMnhMD4TaVxbXSRjUkp5BEnALg
NTOn+UPJb/rP10FtccuuC8Uo2laKpSfX+abksrkQFX1TCWGbREF1/FpLn4kxNK4k
VZjJ/xoirIse3wHe6PGTRWBXvYqOFYMepaZae1rwkonlZIH2Q8Sag8EXmp0vXMlR
X3Pp0xcQW0Fp2onIsON696vReczV+qpK9BbE2AQlTzHbNpiFWT7NJdUbUIn1DoCi
NZVs/lSMxuXJTKtG28aPkHdeCv6ppaSzlSsGGtr0FfI+xXfLAa+uoj+efCW5E/fX
kjM+fD1+Yn80VWLn7pD03D6oehp82N2a8haEH/zSdAaiMoTO0nhQrqa1V8tLwMd/
SjuDkHp5/nuWPJ0H7shmWCluAg/NDXM12PSbKeUw53/2YkY6EsE1hiC+UyMgVhdG
Yha+aUqqHkm5PnmJ7ilFDOrFvhbiDJCr9C7q1WbtpOmNSlf+WgQcbzAg9wEcyAyP
3NXrUfsyWgyxKy1AnANKV84gssCDMAgO3SOw1vRPvQoHpogCCo2yvpISXjwKtZKX
fuu5pCliRrXvNicYLa4Pzn95Pk4wng/z2nBFhVTv6gi0bxmMeCs0XWxX5BE35ADi
MQ1KLupoC7xWi4S11/rx1nS7cFG/Oe2f1zK4+uyOfBz5VRaOnSfWSN+20ScgkIVh
qUeJblwGwX5UwGdmLTPxcY7MRn2H9HU5T6ulIcvzwZuFfvao7lX/O3t1xmLqz5aZ
sxllgZncItl1fqdzhXrydx2RhPuTIyYYKSYeXDdeybHp1SGs3eJGjr1pbiRmz3SM
ZRsSR0TLQyh4QxXM0zsKGeicQ7kMmFWOOdqhPV9dO+y/YioU/iLupBKqJnPBHjSc
Fc7OOiCzutrqGV6HpEifU8+OTxYxwXOiIgKXGYv+GUQhWqIl+Uh5pn2GuCvUZ3/a
OXDE402ld9pD3t3AtwJ8BwHgSqT25Yv5PZ6Msoha8XV9Dwg0yqCmmylQlB8FtwwO
WCB3XzTs63Eed3k/p+4FIiEXdG7V2YwM3FFMDOSfDYfrS75C3PLvRHgTT2dA8Rt6
dsrdj98K5s9BNlCMxIaN24TIRN6wEFEX6sNaV4cqlnVziSkHGYviuOov3nsDlfks
PjVMjV0emZWhSTZBWkzv5fKi7bAMp8UiQ2pBoRZLPTXKNR8auhXgx/9Y0PQRieS/
CuojzVrFL1JxAeAt9IewNPvtAzMvmjXKAMCU7BtcV+zbzO/N4XVzN70V7R/QoFDq
lZ/iLQbBbU8xP5K7QcGBdFIXFLPdA42AgTvMgzlNqHtZvFqS2jnvtInzCN4ojrHN
oB3//s0dqRw5DWpLNVnJiGU2crQlj0BfUaTL3POaECQc3hk2Y3u5zKCuRT5P3Bjl
eStLc6tcxevjNlKJEaRyMMHTu3chT6Z5PULFrrkDm6gYxQebairuZkuI8+zF+8FK
km92dcbWY2dFQjEVU1V/MmbyMqTYIAGGmwSk3WGope9Mle7thg9wl9NgI0GItiHl
gJ4iagJ+lEb80zNpBgX3sKO/C28px3eOVyYDdrY5RmIV/yJIOrT39K6fW+owim/+
Qa6J9XcjZtaZPqz1vf5AcIMgUGUP07YI+0nihhsRdS9RLRZG/QYT3/79SKwF8Ebj
k4DsAu+Xqy91/MZiVCJMP3d2zH0CHLuYx/L4vWxIt28Gd7p7dIfVmMnpTC/oMa3I
RvHtom+/r/rpOfWIqZSivJXABFsriZXTv2d5mTnsbQ8ET1IcJkoAvpP+FKlWKUz0
9YehuBmLEB5ulER3xGf7R4zXim7HWH2etS4P043fm/V/v9bn9J35YjwjzN2C91QA
us7H6OVVeYpSjbqUjrkqI533+H4yNk+13Utnvuy3goCuTYvKWnryefv/t4S/XBIT
Hu7NP0l2ztkd7AQUEb3AHCG6H3WWxfNYaxQlSlVMlZ6yKO38LuGuDjyTDl8XFuJd
sxfiLYWm5rxsPeqAu16Qr+MvqMF1jmpEYzZsTB0bY2k2lKcyOp5iVti9XvCuu1Lz
lZE6d6ah5797xl/YiiVF7d6Yo1329aFsUSDjCDeQZL8k2t/lnqhE1GdOfX4sO2gE
1Qx5tL2u2PflftQpqDPooK+oF2AydS1HTV94tkCX8plH1u7kPZEdNzaLTl8daNvZ
aB+lwfqq1ovTJlos1Nbd2QiCG3h28KOe1ix1gSx+zqXOSo7AnLxbS6fKCu3SE2IZ
Zs123+GxAqeOvdMJI9EddsmAbTHHyFJzwhNlgg4ptxexe3IJY9Vjo6+fUsTSEPO3
i4n55ASurteiWrSoilsrghXPuQZRTqG/iKkqHIaEmcJm9+y91ys3Dil+HTwR7sIs
clIfRv0qRHNxHzNQDgoynEQEbH8Q36PcDmxS7wBwdbKX3Ews4YDZtbiuR43LcjI5
2jcMDu2tjacqJIp+FWzXSqxUL4CobiIuEDsbOs4z77+QFRzPPWYyewLquJT3dpkJ
6G4gwTlFm21yiQ+wR+w/GFvX+lHCAXUlKfP1h7r0rYL/kOOAWNLnRXE6KAWn/xRP
MFAOmXruPQozTdyB5KQqLdZqttQPeuWD/WqQVy8iYZEossEnCEoRzbRA8ArsyNXP
iltmWgEn7B7+TGnWpVufnGwmINvc+NCGUnsGSmfpFIwOHCjL0r8mqWclnvRMs63l
dzeUR64wdOvN6NPvhrWujygbwbOWxxNDb9OUmD0Acw95Ly7lz1QCixR8RxgI+VIe
qGW2uAGN7jTEEpN4VYc5rjqi6E5B3RBsQvJYT1MH5g5bxICJZqkE1VL+aLhvejn5
mPszOndzciGrWDPYokI1ylGZI/GrMjSNxa6Z0vdkxDYXBbj6qB/ZDcQE1EL3ISkp
HldLRTRWi/q37R55sIGpQpVmYsHeUV3COopG34Q1yXF4KWRg84kuNFJZJT9KEeXo
jk1iA8ZCXkZNLAVuQ4Vy8OyM/Bbu/YdWYTSv7JwTlwE2y64GTWhfN12Kioi+otPM
SUhaW/zDwSpyY23s4TpwXIeapISWAxo5xUMHwuBVhiQj7cdfyneYzLhjHX+hab8a
LT05U1XvD00D7JUdm0TS5dPpf8tgSvd/VgsXCmIN+M539rvjY6NPyPQPTPZkt25v
UYWqGPRefhYoEMvCQDKcRKfwbCb4SkeiMzI3sEZXlNFXKVFzKPUcBNv9ru1zkOiL
vqEuMpu6Ov3q3RhWqtQZe+HuhR6m5TmzZEVrHRhj8Tz/uOo1ye38zUot5zwVvI1x
aCm9r7J9bZ9TcQP4IJ+v2FDdnO0MsuR6ym+cwMu3t85XHA0jxDWzcYTrvDsbQz/b
RNdJCEI1KavU9nVbP+5c0/2D7uQvUYsOI+hCWGe9Fg5REIjnNV8LY33C85eKPb+Q
1/PRfi5ub5F7LyCRTWVrJoCojboBjq3ZxBoEZ4mCMKrEoOKGgawpuduZFn3k2xO3
2NSOs9qJVAdLeELmgkJrBKHkoVJbtYbrQBBnXKYmj5R8BURJdUw79WyjowTO8uvx
2uDf22nNme4Wo7dpHJV6aCVuA+BnBSSFksmLJum4radACMe6AIG5lt05tKC4kKHP
kvI2FureBAoP02szg0LTYIO7YC55xZww2l1j1hpAWJzpTr9c46OFpQ1Olb7w4XJe
RA9lhAJBqBmsRLNQ5C9ZqwRRklgXVtzBWP+Joh9GEJU/0sxt7qGBpvmr9+Q4ZZVZ
/nlY0fCfVamBMIGmYlhFmqGv7HBvW2Q7bfhLu+92kJkqKo05cvuoUs7ujWpXgL4p
zC4fwbe9I8f0DrQIMdPgOR7eIcBi2vlFFcEgtTjkQWPdXp/uQfrRYkU+Ub555QfR
usbPLOi8dKhLCNQ9QqWGGMa2FfHjfnPbvQwESzzXZGVfIWRkwO3udIFPh3SAMUW6
Q6NbKQKXxC4MSPXG3W7XiEbCgemVt1dl1UQi9SOOGK1mBd+/koVoznsRhml3UJrb
2P9BJdwsglN2cF8m4nN8RpXTlHz/2+y3sW3zD963bvX1G5a0If34kNFCfjhNnNJd
DORyp0oA2zJxeciVwNxdWKkHFJevia/tZRlKgHxbd9+mKsC4nWVFCNDVhF7HgDZG
Ooi2WSzL0l3f6iIrdZTj4TD/4SshgYCtX2SCJrok7sEGRebvKxpuSxs9X5w3bPyS
5M5ZMEh612hYlEjaihd+nbS5XSp9JmLHUvTZ3dBk9+Ed0UffmMRT4Vy+Ts5d20IC
5vdCxEJUPaIHWEVjEqZUtJxgR9ntr3xQDBP1nVsWkxz1qJw8/RUpSqznL4DQUUgR
qq9ZUKCRYln2FrI4bBy9Af4vgi2DYR0X/GXGHrLktF0S1s8viAnCL020AH4ynqpY
aUyh8AU5eU3YInjKVOaaDSHH6/dqf4g7AIWYPBKHk0YCger4QnUu+xxK9+e6/Xxf
ypYjzL4cB1LFK8/QNUNv4WastQ5G6Aqyn7UjRlb0qVluJ0YEn5SWlVyKDudK+Sob
Mdzyon4XZ8h5icCwiGy2dRkqSj48lDDvlJnPumYQdS1NUV7CwA/1kp8GF017UVOj
YaGobHoRi19RSWrglx0CgRfblNhl6vZHIPuwPdjpWkm2Gnu06ag0snknIJ8F0CCU
qnc5cRDuEALUCgsK5dqvkqM1EYrc1ar0mFOPJo1MjnWEtpIz3nwDB4Guz6H0lTur
8XeRwOMMlwznSrXG7Dkvi5KMp0oDViv/a4vAQAqlNI6hhqQKND7WUw+VE33oHEq7
sOg0iTqLvHOA9BpWKayldh4wfpX7iji0iDzsX94PhtSNgGyAeCXePqR0HkIktuJH
fx+IRv5kXP84ibSLg4EsMS7YZHBo+r4yUBcoX2GWSE6AtHkIMFrDQDHE2tar0wZH
JTHPqIteocMmrKTNPTeydkv5ceP1MYJWzaKlKRCCjU2d0SH1Ib8w5l2blydVrnk8
A2ZMCW1DRAVuugWB4bcWFmprLgk76s0dJbqtAIDu2dT1UZxVUgbxoIPZTdK1KKpk
ZBU0JNQcxP6RW1w+LYKdOe6dILcvxb7WECc0TGwl+TvbxX2G2B234+lcAw1QrjRx
kmE6fv6syNWl0wk+v2qDJ/P6g+aYvehburFPDMlEYsiHARgOTCYP2i6RoiJVABIH
faDX6c+P3rD1W9MDwI18p+kX8sZYt961zklaVy3pvhjvyS+nHLbuD1gQb+U6t6Hs
jz87YAanEz+yz0p2mdSJYBX/1gjLpzlUh1kvXq3/rcB9gBxCTAtUdsrNRLlX/G6a
iqhzYf0VkjQb9c8WetobMqxjAEV5z4s+qjl7R+U1nzw8wS/JuaORDqTACd6m+nXy
3G0KBJ5ElD++XnZr41x4EI6+5YUTCB2/LJ1SBQp27BZybfEiLubQkWtT6kM1FjAM
H96LzaCmcvH7zXJ3fuMxCUZT0R29cWmB1TuVLE5dPMOQC+dQK7NifwEkLYeejVPH
uS6wUO3KvECxRkr6DgJzTKITGkLr7so8MH+dZUVffyNFjiE93pl6FBbjpF0+IE/A
GlIdDC+FPD07o+EJ8jGRr7zxpxpSb/lsKuvr0FBTJQ+micRItFAI05m7wtaDRK/l
obIybtNbfgtmzOYdZD0EwLPd/t5pzEludOca00Az5hYRcdzfyM6tW1vf4xF95RW6
p+jVZD8WI0YckyDgIIlnl6tMMhHXn7waA2g8jVVUDk4A0pNQdS0FCrGoN+q+ZzP1
MIM8hchmYpUAOcceyNAY9QOiXX6hSky/fp/38RnpmLlYjDPHeZichPy4UrIAsHRn
8JTkDuR8oWfE5zThbHu9Xl52wbLKFh/v8/rvWONQJJol3wOzbcpzzIWeqLBW3Idl
616x8JrnoBOvWCsh9+Djh77Bna3y09gbMnK+HFYgvvoAEZV0D1BtudtttqcFTTrb
E+U/q4/15pv3rAXYiqcwft7Mb2q9VtaSeO9/WqMVMcLCDj84QOxxMwm0Y6jp4Hfj
VC7ArlVuQHUUdjunuvZt6RdqeEGYlyyBRQUoIA9J5b8uxQSqJ3W/M660U44w+aPw
GC2KKU/3IdC+2Muel8Cero3AGY+E7atg2DajOyd8sJxAmNJ9rQGNOCq3Ezc0mQMJ
TuPcTQMC2PCgV6GRTYwQ/TkO43XpPF1TLgM1tY90O1xkbilSHE0BD3X77FPVHF1o
1iuHMmgRh60ZKqY12d1s6Gz1fztF++xpHWwU4ItxmG9bLdqKF6qpEiaxYzd7sRDV
NTBPZmHmVeC51x4B7z9fTd8/dZrgPMDXm+FpycPXOqzT9lpiLNfKoaokLzu4bJMF
6DumkxbEH7+orHb48MpF2FPjxc+8bd4xEAy2k9omzC8G7uuEEztUAGFIqTFSEUof
MdD7atB8LuigxzXdUGr7zRkQz9MVbZVvPD7KdJZN4Co+P7BWQgYYoeWqttX5YNAn
c6C8eKtR8QC6ukaK3/V3auWdkamRd2H5KuX83Q4+SwB/kri0tkbNwoo8u8xU9Okw
rdjgy+k4jvUogoyhH4JPg7SGMUWHI0LxpKZm6SdKTMyFlLo7k1x4Xw6Mkbrb/WXi
5DMNRIQzt9TMt/s5D30YgeZ9Cx1QR0FnhJnSQjtvWZxpp3SLrswo6D5CJyh0+U+I
PpvxQ6/iNmECyGfWjeXdrpbUBkI7XDkic0zVJ/cR8b8UNnovpfMIIS8MBUt5aFKU
W7NubNYT4rLCFdjRUSf/9xdVRmB0oMQKKQZrlihUUuoMuLkt3NUwKxk9sk2PGg9d
UjVvOB1CLPAFXDelsOXdtg64us1dPZuRY+fVqRtQljJSy6UV+UHOYOVuChS+gtOe
u2uWNWoYDt2bTLqXflHP7ld1m11xDpq4/vg0u4s5Aj6kZYx+iU9TdKRYozIf0uEO
cnkDMKgWqU6iqpnaoss/xIjuyjVdKvGZzzkEFOo5x1NFZp3NIRJPYNwVOY4bmGKR
feFPa1x9y/e06rZj7DEVXp7lYz6BMSageh+PV/0rPQbdbNdrQCZiMsTdxJbqJP5N
wq0vuY2333VawhSLIjbBrygZo2zXQB7uZVT8QpU+V8P1knpSXh4AxlzahaiJNj9F
1hLQQ5NCVBS6j7qGEQIEwXr1hN/g5SqZXJe7FVKv7Fg/vJ41/1gfOPeKOAv6kfMF
JyKpg3Fvmpd1dzUuOHmQZCRnPfItbSAD+vqKMGU6nCdfB026a/C6rO6CgAwPvsyr
pez6vPBD4cVBlSSy80PnLpVC6SiY7eEoTtOkrkF015S6IvYy3RBR3PPHurbWnUyv
3pGbfj5SHoblLCsfllU+hPCYOK5/cAQLDf5Djixgwbs+UJe3i1VCxN8fWfeDsk+z
0Bq4OztJLwo8c8yNPmuWmTjMbdRGwuWJXQOkAi49eHgn2T4087au8E7+aCGBWSWs
XwRu2NJnyA2OesQGstbhZDRpJcwFVVQYuGSP3HVSu1wzOFVzQhIUlgnvZrHF6Y+m
Av2MCt1RNY7nj1YggfrkIo+sVvv6Yhget5wDaZm9s27MZNn2wa5vxSxaFTIigsDB
QsB54QRvJAcCccAcIETEuDSW8fAQPd2indcDDfIF0cur9L/px4UxABVo1DU7qmyt
92KJA6CA2IzbgL/ksVMgDDALiK94mpaN2SOyCiUzTDPHvqTHfSQSXLJlgiN0fhRV
f94mCttbEsHi3vhtj8S0irw3qxwM+Jmt2eOhT5Wawm4NuF7NuKN9FlyaSF6i1Bzj
MZGGEErHBtM1ykPNpArxa+eZQZNRKNrFu6UlXwDLOWgu5qA5LX1OOGhhtqStIILT
vr/7S/kkCz1C2rqwSYDkwYocQumpKydjF8B4nGYJRdRLvIDUeXqhUYkNmXEgQeXM
iOQAs17FQwt4ITJ6YaeU4PfjpBBNO90mRQ3VFMASkfRZ4B0kii4Ix0PPICazCajc
9pXelNzWuHz5JCtQjXERjZRRc2koW27IbdkSSx3YvpJHVb90TZmFZnypc4GkTZBX
Y/jqpHHhNWJLA1C8Yqtdh5YCFtTFXep3mIz8C0WSfjVjIRMVbFxCoho5d8US0n5b
OTH7YD2SeRlAZgZVnERrHXq4Nr8RdP4vfkOqIzrOzG+KHaziy5umbPGfrY5G9MC1
/e0kK/wRUQZLad1fj2DSaMsyvgsHDu0E+btZqrUGrmyGvEB+JMtav3m1ptpPr6wE
r35YoZR4ttovt5gWFJUJI9Fa6BgoEDdXabJmC1fgrq791b5yWpXVYXNrQF7IVKc7
YLdkpaw+X+bes7XUoQT8HEuMcISk6eCiYoBuFMTOhI72WAqTd4vp0u4zQfvjX4Qx
JV8V+FBbJ1eCFDz6inEoJFvzXHgZ8N9YLEX3emakHGCaWOwJ8kEos5m30J7hYWxb
8yjABD8IvXcmPLiig0936SLCjVJVFN2TznWcTIJwdAiaOe4Cg4YpuYLetlOtdMGA
MWbP2oBdYebn4TWxrzpEABEP0HiWkVkMuH3OwoCg/gNLufjZ6YpSsairczrF11ln
9bfzLmFHBwdYpWp+J4DVDTjW8QNF6905cLyto3W+rPMB579oCEURFjO9PEh8Ptmu
5TQfxCgHodKZxX03C0RyYuh7XbwJ6JXhLVanXXSDjcKBuITMlJqM5IlspnQrwvFM
iPE6zeqC6FSxh+e8UPyFZRFjvL9wczqyr55z17xr5uU05bnPMQl+PPonQWoxH5Fe
l/zFp6I2HJ+j2wOctlAu/S2fCd98tluwvTTcJenfOM+ur8Vcj/v9vDBNRjcEiS2D
bnth2F1dHdft7wwyv0u4TuE61QFx/ePs740iOeffDLWmoIkkagyONX/gftQVxeEE
caLqfwhREaG2fY9I3DIuDSCIwmY5vd9JinceejYISSxpZUR8xsXJ/nvV2Ra7HtIY
qOnukb/VPlZ02V7E6L7lKrWuRix7ThWSD1WkpEMIdrHYSElmbv82J/rmYIaa/5Pr
JYEhrus3Hgmz8Q7sixbp8jpqqXnK01JUdWGEuVT1ZUa0fjQ4Vv9qadX3Oc6hHRUz
jRW6aBMC8EFXhA6LsytuDWaIpM1IxVbDZX/+ccWM+UsHbfZbHcfpnHD8frOjHxZa
FtIpeUNr7MVaufwlSSn3TrWExbOaeNOG8bnxBxBj+ztXuzflq+As2sZac8Aq4C27
L0GlXRDKthPCjP95C3ze96BwmPYI2xT58YIXYmOncE+nt2R48RhezHnYZ67hR4aT
kom3x78iBJQOM4ILroPqwJfck7f0uyz6iY/yKGDFBa7VQClon1UTXAGYz8cqCYeV
tm1yTm3fi5svwso/WkNHjcQDlUlQ3KUNl4O1ovkqguSPE22gaemLGdiwKe42kl4H
2H8Qsxy5gDNuodBeYg/Qroux1AP3XzuGuTFmgcBvxhBatOrnawJILjrzV2D//1X1
fNjSIuuPEN/vJLqm3Ayr6LehdT6iEkhIKDAaIVdeKiqnZvacbHBY4vorW+oi7MVg
P2H8S1xsG6C+2UlX/8idSsr4Ndirg6VxgboUXzR6U2KEAyRiBh1u6mfyU8ncCP3/
Aubik0s7gczh5bMGIwQc8WCzU+71B+Xhl1lOj4z/rqQcc/lPWQ/hWWVwKvnOQP5i
fgfX6kWGl3vwWh2gc5/Yx1TwUd4gp7+/ufvBCI9EMP0zNR7Piltq4iNF+B9RUMBv
7DiSNXvHBwOAfMwx5MYU0ORBMuN6+k3yUOH3Npd0/melwlTvWLEXKtAIFZSGhnM0
Pi5ojlpc/AkohRhL8PJGoF6sXIan3hRFkhxHKmRvmGscVHiHi29Os5ImWoMZyM6+
Rsrk0IPzkaM14fFCm61gR/+BHVQYWY4MxV/LhY7XNxfe/EU9Q80VeBhBTbDtCAQE
VgQDE+pEPWj5wwjxtT/hz2PRf8r6frsS+NqSj6vLbMGpYeP5zQeTpfhi44RVMggo
LpNkkJ0NYF8l0ku8jp5nkWDnMfpy8HDlYfgwOOqzNmtAyZev7vBwNGCwpS4naAu4
QVh7OAsuxHftTHHGKxzfbxKzxYBpcYXYSD++L6nIGfk7sQt+pIMaIPNZ4rtp+QR4
t5UMxOvgp3DGAAnLNUTn4sSmlnBHd2aWH8Dk0MNE5p4zpfgz2SlJANu2VQ0sY9mp
9TO7gvskVVa0DvYgGt12dop0Z0CMdsLExl8FZ75dfDgZeU048xzGDvxz1Vs9SOnl
wK99F8rJiq8bQUVjdbwSuinMClIAzvrlPQqj0YRZmHq/7oyXg11SqxDkamgUqwu2
VyIQg5XLS2Qgjri7iMayErt9qXpB3QB/9HPctuLbW6hI4I/tOXIk8hfCpC3r0CGV
wyfo9KQt0CI373VjZn/OOZ0aU4Az8lvtqGgcxnqvjyCNMqI+ym+SJd+JkvOqyK/l
eIsR4ClXgZMaik2RHkLTBUev2b3TzVOxleKn+MIG7/YLUtc78tFY9jwE2/PWEOEK
vaU14qHRhbl+DKMA4IX9hCebuEwjREoJtG0VJtlwzy+S/3nw2ZfMOhOi8+OxtY1K
ZHGGkttY4q7l3rj+8IMh0jEli4gXyvsSbfU5m8gNnwU8yfYhaSzzXAqARigT6MXu
rSwiOwOfN/1OSnwAgFjZH+VYlw2IeniThxktQu0Ws+wAQ8EulQNbK1Ehy4rVaP2K
VZlzuRVkVSWMUdSQFHWXqdyBSPhMKQh8tyjAf1LD/dWU78sOHPN4+Ov9ADOIOymB
DOMbcqAgRmCK0r6zRjK+hoP8JFbzkPZqDsqmO1nafg8DvkJTK2dXPzyNfezmU8VC
68x8OI2PwIyj8KqF0BJWsrVA31ZQ3qTnyU7XyuZSLqmvA9DTZsSyMtfQ4l3z8RHl
NfbTt1vMSbDGt/pNo12ryYFPrQWOLQPzZP8BE7jaK1iYvTY3LBpYr8sJIoVJk/uh
3ZlaC9NNzSX34ULfvHFdQyv3HDmnVRQOMLBD2Hx5GXbmNyw1YGab2BUeulCa1A+V
ssLVk1XiFkGOskVSY5FKmswCjVQc9WicsBsPghrjw7JxBZMkww8wCq5jwu3i2o0s
1edmudpRLWG5JAfmc5xPaMP3zaHwA1EY7GNV0aNwA59lOHfwtOb/h/zPKK16qhIP
qlwd3fH+McMLg2DiVB0OtjTD7wVvmNe+xI2W7f6AEHjFhR7ZCG6mNT8kO9gMJvAW
eARvQ2q/XTlVzcyOPGOw2kTlq6qGkeDpNNVDDe9hFFJkPf1yM4/UM1r61Pwtkpu7
GT0qn3UGT58yqha0VwZpzA/SnCRgmNe66DNEbROBvyUwexwObRaTpX4j5gz0My99
H0iy3BApT72x11Cvn0sVfY5IMHc8K9wUtAX2rxXYOV1RVLAiWoBDnBmna4W+G135
RH69VSV+vTuMZ57gWkQEhfM+kT8ePMF6o001j+oZM5/U186T015wtW/fZ/Kqwvre
6x60A0a5l8aR4xXHZnDHAjSLrMKJ85iTifWqTKhO93moE75hElig/K6x6V990i/B
otYL2SuS2auE3nn2HfMfD7t7W9s+AZ4vy/Vsm5mnnI4oXt7eVvBJuUMTowaPJkuR
xZJgBQkVK2b2W+rSHbqFPwxgUBHPNvygW8x5oAHmu6zc75a3Nhr5lyBbrQRI6Uuz
6YyLnGKJWrr1c4ES8nRnSwwwtPUlgknQBgxey3FKsd/BIGQ35TR8sqk1J1W0Gm15
7T9fp4kIZZRFxGQHY4+idHJ6/6qt/Zm9FGxNL1S4fQbO3kEvRjYEdwk8R++2Rq8L
9uZfD7OQ7vL9FAwTaOyxHgcmAlMZbibkdFPeK97hI/bqQHboK2tmM11zjHTbdD1D
3PtamcWAW4nakOrEuvGYH6ysxe4r2JM5TRuUnUZLj9awhPNZqkSjmTCvEODNNteV
iMaSlvcpYs2sHaQAAB7lzUhkO4r2bjZSljhkaLfBxq/CrJlgw4pF7EFqY/XUJfMk
rrO4st2LkVWm7D6o47W1mqvwi5jcDK4DzcLEnKJP5B28mKaC4k5EipTshGD42fBq
kp1ihv46H4OMDo4v6nzpsBqGqbioKwhx6Hnk7hy/rh004EoT0tkLWUaq0A8UZ3Z1
rPRCQTxeVERgNv8d0IqMz0fkp7XFppGqLHUfm9jdP34AEe6dVghw8cdYrirmVJ/j
aCnidl1FtG+CRe6Z8TlX+FyqLJ7UomHaquX/8+SBhua7NCwvFR90UBnEaLbjpqWS
tPf3TmJxfPsdYcLL2CQ1U4N/Q+nGW9oO/3pC90mnjArYoqbm6ByZBYa+X5FuX6R8
RJGg0AcKQtDyyd2H5bvijFIP0Zv8q4c5otDQeOa0tF8IdRff7+Lyv9MJmuiAbjzU
vviCyc4gsSwwHqMLioiyL3731xviu46F7v0v91J0F5JTyrxHDUO52TJtcfnXZB21
hWnpu7f4RMLE63qLfh/n6qwcRylTX6CND2SXJ5HJTTsfogLoHG8c7a+JOcV0nSt7
jFhMKf4sejTsocEASYcFWzFggY954G21a3/b650gVyxPQabib+H2/xaUew2Qavfv
2HS7nm9eQW0m7ZJKX20vFHDKNDhhdKvxpfk9mexGc2JOjRGYV5iW061SCAxGMLiB
f4PugnvB3+Z4K/PXhtrJmJwOLEx0oAqPiVMnzdrCHt8jL/fM0pVb68BVqkDtrQAm
2oqN2ZeGv2+dRHoXkd8ixU7F60bjKjnTWo3taCQRRvs3Izaf3c4BVoc9NnSxPmz3
HCaYo/2s0nOcTBcMwrPhlLUp99JGYl+135yFpGDBzjly4BFQmCmT+9gPwANI6G5i
w1TrAUhZsYpBktOENyIvkD/za1viWoWd0MGPUVVG4ScggPZCzbI2VhBWNahpC3ZV
rPsuDMU5lJmNnK80CobJMxkZR4CirVkOG+eej76xc7FRvWnFweW9fdyOMMoHVZq+
vBjxojrsRt+AxhhccL/shv1o+RK0xMU9ZJt0yKbvMGyozXroWAzFkBykv0BMQeLS
lj2I4AkEN9Oc/PShtdIWRtm02rdSCwNQc/9+U7MJdSGOPSJPsZKfUob+ujgkf15t
3TUSc6Hl8aTQk7dJ5MfAfTsCZIgB2/8qBqjfIBmwsUdfQ0y78w9g2DkpcYSX6NBF
HNURZtB00DRKD2texcYzMZZU2EvoFxst+GEZDDhgaqN4QpGR9Undv72bn/asXs3j
+OxLyKIMqHU2KM2oPbTJ0kg+dTENH5MCz/BVQJm1aUU6HCPleheM2bPcTJSJ4jTd
qTs079pW4hN54hJT4lLPkrEUiXE9LKgmBABLsaCDwBzyI7Kd1pSRVCLEQBN6xCET
z/l9U3h+bj5t6A0yK/hgCCqERVRQYHT/LtGxJakT450r1nLocUZHl0mYjrD23HI6
BdgYKe0oqFKJrLbRSn5A5Yn9uFXA09iMU1xNBTiAl38CaaHYGnjxSHobtCDjGe70
+XVQRrV5To24HbHtIUc0Wia1f4qPkRcy/eqn25Ltr+fGdmaYJ0OE7Z2nGs6DEHo0
5FI1ItHC6G/lQntH0W3cIxXyIhcY3Tx+9GPN6lz2Fc2et0sCVmyLUK+0Kcu9GxSa
xPOJzoFUlOUkXc4b/CsDxmQyCbBU1e7uCrNZulLcD3ZHCsmmGjgpKz/ELOK04yup
hPnGGg4CmvjCfLiq5gOO5pMiBNaDDD57O3vDDw/E+vofCt1CrG4ZCaOLc2KN/amM
II+qiG4xYff21s40MeCQV0XaMEOzr6R4r3G7ltTienotCHpNsM/i5ULP302mb6cd
UjeXz6wi0YmsI+bdodSlEsUKAihOdp72Hj0u1l/JdnyBLf+1ErndK2EYI0cOQ7D4
cY8sEGwP6pRg+/4F8nIcfFecEEDFn7blrmpRko8dH3nKgQ+wlnqZpoQkb9Cvu1NX
AqqxuXX96dEa20XtoXbJ1ab+Ubl4VhaJ/XfAOEvwxAPf4nFyln6+HarY4H+w8wBH
U75cFj/ljxg3bvroavm6+qtmRz1rVk0SlYDo3xO6WfgAwsFJ1LWlpqsGTSwh+aCV
ukQ1n1FzG5Uw6QjYZE05kHuZ+ZAzlknAaaFagBUJd1pb8xtYO71CF30cq2wC3KfK
i6XfbrvTOfDGOELatN0yyfxzI6uKzCFtrCEzEBrY251z/Y8HHPNWQL0MLpzSrOle
THcM+xI0gNPYqbKKSVlIGPV6BTjvZJ3MoPEfH/N8eWprtZ/3QRv+2T1tYTEghQ46
3ELOsDAdCbevx8WaqgfrdF6tRYVJPZ+OxWwIykXFfdTl4cOWluDE6H+ro2AHXNmt
1XXEH0pxcuYULbIcjGic5Exxk6gT2vsraGkaZXszfFD3qk3qm9/ofgBw3d0VuyUe
nGl2W419moPGdbFvi4+R3f0hNSMYd8O0KjQaobWGWhx8hRhHOWBT7qIlHgn1CZob
bLW1bfW8O6KDeOsMoZyZ3HGfDCEmXYv0R5ShOi6MblPpJnJe6bsyRznWuAR2Amle
dLE/QsX7mypEECUPPfEgAkErFTJ15AuPo1ePXPkcSYRM5JHXYP7iWHjaOiPU5pmr
0tW/LEqDMXxgJ58BB52fIKVC21KQx7BkC7yQ3x0v83NzIWasDm4PQ1oE2/xWojoP
8waZ5na/X6WzxhpMb2p8NsmsDt/+/ShkVo+VDj8mJifCdk1PzhVXOsUimST1WzMl
VU/flnk75Ur0c5rdwr5mcozHQVTHgc2BLLOyzulPhlvhXkQeCVoiqa9ZY0DNlNbA
0r7LyoT4qXMzzKtoDqjxni4vDNjmuXzvKHQPfuWpKtOKK32+LphnzYwWAw2QV0eq
2Kg67Wp+gbX2g7NSFADfNeAGEc2qi6kX+yV3HFFQ7lg2ZJQLWmraw2XQYr72VPwm
jt1uXe70GlXq4KaRWgoDxzSxlvMBfTRMSWkC+/Ww9fxU/fK4KkhCxbYYTUQEo/em
df4QoUqQ4jhJbRbOGipnA+c5nYtuD8kq2FrkkUh9aCh4MaW5wHSxuVPKgycSi8UK
eRradwkeXnrOl5Cx9FiGCm1BFzVUH8ArXCUk2CwIQ8W66q60lQ0pgTgRSEKj9UgC
tZ2P2zJCKCxoIhGnQsL/cN0WqEBUZtyGO0m4ewXGPT/9MWMd47lrF3+RCShVZV4T
QSg8TtuGMhLAuvXGxo4RejI7dK66WBPkn1eYjXeuLAKZxBRBzo6U/XCfCJxWc72z
StDUfkmPGnhb5DmszYFciHKxnkgCFlIFgBtj/+P21bvOFa2eltJtsfkd2bXc3SUf
nUmHsVooJ1O4+gpxn+6TWBU7DNKzurrFxQaE3de5pr6sztYX62hBoULd3UT/q839
QKYmM6HnAerEAYXUuYE/0P/azDQ5b98bS/pee1ZWT6GCwGhva595woW/hQr5Ix0u
Rxcp6eHGK0iLH3oFLiZr8KQlhs9By8yYiFlm3pBn2DvZD/5FQdngTavI/z8EFEPK
prioWpcioqAT+OqZji2EOFc0z02M5j7XKCXPeDIRiFIZeccVzv8JbrNru/lgiEWg
0UMGVTpP3DmKgi2zP4X1a4iy9sYvBieU4dY1X2QOdpuuTfZIav4b1YxkHBTe2M9d
fT36VdJjlF8YUPgsz/l7sze/K/9kmlgdgwX/fkEDQCb6o1DmmxAKmx0myI1TPHgR
cuI9FaAwHxVzFlE37+/lNial/KFGs207amNGRvSj3FZl2+k1WHQHVfLJtXXS1oyS
9XILFdwe2YFIJUuvJU52SOkXd32D39+0adkc+uge5Tvd01I6WgmPj2RrE1LaZGa2
diVEabrhvR2VocKYjzLanQQ2axefBEcsKxV0a7yAywFcVpwkunClheyoctmVloqD
mrwKcGis61wCS7733AGNWwDLWdMifwr3zlHSzzYizNTEUTJgv1jNiIFdn5wpikqr
obnStx2IZ7+tH5/qDnN5TdLbfjE/cx/co1m5BQ87ohhUNMKNoUcsW5MK85LafpCy
44Z/cfCNLqAGyx6q1WkAXd3qXNfa5Kc4dLatoLB0MlB5pVOTL26PVBWTgfolGcDD
cuFLGM/nl2UnD4nDXMG31wSe7Q/3+N04JuG3zXn+Z3gKdV6opeHFmB83ihc88bTH
0+hxl9xU/YFFBnU1uW0QSRQDGfy20z7X3lTacJH/ym/4jf7XNyqIoFms8aQ5EQcp
EUBjBqSK1wFkS+GKIf6fwVnpa5OJGzCcIeKbLOCaXF3paWLVRIldwMI7RQaQtTY3
Oi5z1Owiq8JPBzCVIGkvNCtj7TKPtjUW+8dhBmPnMrABgL6y5rz06wRLlMYR6Zo2
WpUW8Ob0Bb2yfA1LP4l6FjRorPMwVf4HqgjRAV9sA/gIJyctkmnRqlYrqu+kJzlt
1fV40F4sANn6m3PCWuYhGy/GzXjR50yJVl6MTsoPuoLAwaVPHNtWt9QKQHezPQE/
kuItPa+ASvxSrmOhRS5Psaw+Kqf3CEbG9kxuyl5dpSLCQqXjH/BolpO5LRUyTDpW
7KT+0ISV9jNz4vilkNEeSfOcYTQqA2icfGXxSA0o6cURUK0YmTQYOxZ/vnqWhbLm
jrhzgUQFRa7S06qKUziQ93q5QN4DDcWhV12SLl2hq41S2S8xug+Fg38UXhbmxGgY
EEfGtvU1H/Eei94kjgFwVUlqsY5btcEE5dkvC6f4as+fEJSjuHFQoEmruACUDM7c
sCh3OW7Kmbab+h+x1P/xXhrpR+caogVru94Yd4d30xMU5A9DBvNDczDzCqJLwWhU
iNg0H20+cVFE2xIt2x5Y4mEkN/lrDnTWpQDfdrAc60yCLFYJnWZihlZY7b5Lk6+X
Qd9YGHmYcEjShoDeXaoLV/vshED+GW8AsIJ4sMSjSMoCydWLFuIhXC5UsKr3GgcM
Li47D25O4r43Wd1I5yrcyN/Lb/1zIxJQM30rfA+pZNmKBanwynBm6V5K7Je2s9YW
x/jAopkoRSerbqRY2n6qWTXl8NDQnCItcuwHIZ/4u6RP0p0AnnBWbCF6jUmVhLNz
94gNqrdNyUqjmkr3TFpVGX6t8U3ZEQmyYgU9S4cNWn6EzbLxGai5/ZsAXCq+IHfV
7WkePXRqMhNbXQcn6zbHgilLr3jkJ68jmzfTZaNGoagD5oHDyWc2DPJucslzyTMC
OpRBvjkO12dOMPqMIWXgkVPHwJ2Sf6/DO87Dofn64uylnDajPTrFcyVDVB3+h1cM
E3Ms467vs35QbIjqGvDf4PEALsEUrQNMs97t02YhXM3V6S1s8FzmmdBS7wsf69kk
DZd2Irro6H3JhnkbfDawlD4wjiInklDX4fBUaGEj7uVJIDs+HIgNY37QrYeRCFlX
326aDX3r7bjO+t8KWSh9gfdXkvm0Hit8ZZ3KbEcvn1eC1DCL76m30+XIlaj+2ojk
zoeW76RxWnx9rncZhesN7lO11Ezdq2wabJoLC7aXOIAmwofd+TaAmgsfe+xiiPj8
r/eobMktIuIgl+xgSpcwuTvh/bvV7EGMh4xCzXIH1IyYAKfsfQnwvUNMigcJYOWK
VKPl94dHiihxfAxaRyLwJA7XRDmNhAz2YlGrCSmdF0NzRPr/N1TwEOBCE+JFPtRG
x4/te+qh9GoAPw6GOPhh/qEnDlvuIi4kXDX/ycz7ELzifwYvxe411dBMmsTCzdUL
J3h5v3M6XLoHLg7JHly8MhMd0EGR/wG35hJbsXQr9wnD8hQgQzIs/BpXuQ90ap6L
POvQLbOI55rFq3XxagauEb3oXcoFq/kARKtYA3hqqyGHovsyAphjfVXXnYojoOJG
0tIR95/6q4x5rpuEvfYoyUW/reoTPIq6r3gab3szaO4ELL8f2BdV6gAMGX08M17v
C9uKJ0YylyVqRXlfUDy414WzFBM20yzI+4R4chDN9A3I7mx98VHpuueNZA+fJX84
GY04ime4yUnXW4RwgYjyPF5v0RU0rqj9acDlCP3i97TrGqieJkfCzR3vKbX4790l
gfXcyaLJU4rNt8ZMO4ktZbyLSsdZwJ0EMG/vrV631lBe/syCDkrhKGAGZEcPCBtG
1oaJxjzpo/y8+73LWCfEbUw/K6tiRvm9re4fvXUPCoREkDuMG/abgTTUqKgiF4Bv
HsKoUwroWEAl2CvHbXZzys6P82MGBxBD/jUn9rvlj6hcO4pUWLfsizgrlX4r6znx
uy2KM4TvVe7qz8jIlfSX0iyN8Ld7YScTIaJeOq4t1hN96QszT5qeD6HusTxtSfGY
dBnxjO7K6lDezfYBTcYYATu5ZOyHxaYXjW8DzszOjnuh1ygZYQXqbJqMg2CzPZt1
ChU5HmRjt7WGANcgeQ94W4JNeqQf0KvV8S5I/vJeTNwFxDMduQRQTexFJ2BkLuM5
oUNcemiSBZrayIvZ5VFGXZ3Ut6JTOxh0Vbe8XhwgspBgrFLTyUY5QJ2/jXIh/WJT
S9GB7qs5ovkCvbPY958RyA7MRFNxap9roxo18Z/8d4K9LfRd2jD+xvQda8PRFW4B
71hOTNy/9I75qWGnWUPcY6L8A0nrChkssjoD0s7B6NzcTaYxHKVKkgeX5y+AXsUI
LKIhBk8ybFXfpqr9Nbai9DRmU0emY10Xtanz9u4hf4oc8Y7FUWX2EeOwbNJRb77h
AEgwkjLfVbkHHYZtv5bfCsVk6TAfDLEgEzKsqM7JTsBnwcSOI4N+BotTT/jqlpeE
RmzO7elolU/LFn0+DN1CtvyuXxgjShGJ5IQyZoFq3HnLge/p+mQ+h1UsRMZpipvi
Z3vM5BvfelLQMSe17EhN3rTpdUTKpD8MXW9q1/SfkVxJoR4tLAH5XmWN7QM6pvvi
bK7qhvXd1PEX96E5aXc9hHGTBBUP0UkeHB+Y///I7DMBOHCH7hULcFIMogjdd7gn
dQvtdwhtW5MM2lhl2CEvLfi1BDWFj/PDCiFMOe76t1cFE5e9+rijq8laDC2OIt2G
ewrp2WDbHihgXUeY5uhvSKHNvDDwVhDZTj5rofvGt9RHiIvcLa+GceYdt6mQiFZE
s4o3aMM0R/Nms3/xMVBbu1FXbUMMAvlrt7efSBmomEn4h8GkZxAsh5zntiyotEVB
+m4JcTu7sDvADknehOWhRcB6ZixYOocEz6vjfWxD37KMSFv/dmF149fJg2KfBZEi
7N+sH2LAB8hcJl8K6cxtwXyt9vY9VNBckOo2LDcIbsB+Qr/5enGbTSPZmbB9+I7g
0OIzE1d1iAvsaAzSJJQweWLycQwhbAld7zNH4rQx6nCXiTuUNutUGnacQZ8G8F+X
S0pOGl8IuvxN4OC5NzryjFnaRbPn1aXf29kUum2tw90tizjpLSnV7rPO/PQ7w8FV
Wdb4nY8GYKI+Bbxj2o/jb9bkQWJLwWArgFx7Fi/14+y8aq1Vuz0WKPq050+QmMde
sNY8j34uF6ifYfKgAbrsyf1ubJHA5a92Diu8HAKMjiAWOb7n6qfuMopd/u3rmII3
kctQ253Pb8dfpIt9cALvHbdOUdFFO7+zbQKh7RPLDLT91RytSDtTm2ONOywqPSOo
hJWoHdx1ZBsApmYSW+UuqOd9wco57vB1RtLlMJhOthe8rpsuh17Pck7hAO/Ggh/s
XnmrMoDk9MOmC+Tb4/zm3bFk26B7mUW0D4z8ADbbQaUInZUAXFDnWqdPbkh/VeyS
qICmIX59HhJ9MO/nGUL4AR+T5a92hxp3dmpcG7aB5LxtKz3v7e9D+IYRqHCQQezn
GCvyRNdlY8H+fAdJ4HqguHlYoHNACYV1l2LYreuBNkfDkvOKmHKSflqn3xitGE26
hXY0Cs0ELvHxSSHKNSMlS6mPHKxO0OI5X6lox+/x0oRzzKVT44dcTLDuBPKtWneY
zI9I0OUgQcPxBJ4/rp22Eyl6AaOCqGxpxgGjRrIC4wQr3Uw6QlDHLBcOC4dtsWYa
alkS2gML+2Pb0/AnasT1mmETWnNnPBYo8t0nOCljWvFrUxYBApr5jUBp7jkjmHO7
1DfU4wQkZBjA/VQjYXCNPyUzpUJs+gf70AMWrq33siktJo8YES6iFYGaropNEOIi
ViqSbrqBMPXAfK+X/OUjOvZZzkWsXnJhdH3VxWs0BYWG5wOrtxl0HDbG/kQhnsR+
Ck51OqhTGVTlfPyz+5G8A3oGSgaagmMx1TivxPulHo63HfdQbAnTEGcaWkadVIwx
x0SjZKnXa5vL/sTw5bpK1ja4pKu9nEVSQu/hkG0mXj2e9g1GLrUdXqlPfCqkU8oO
w/Ijmmm16B8zf/uTdZIDFAhawfBGia9I6K+Z8f8lhrn47c5YOgf34eVblgSwiDou
tpp84j0ZwHipPgWs98jd01liuaJYysD8Us8Ua6UJNmcKL4StmIou/ryZEeLoz1qv
3xIXpehpQaS4xIqkhUzKOsZjDtem84hi8CJebX/73C11sYJ/CNB9KO4bA3L+Pd1X
YRUX4sTFkOGTpGkxZP67A+qffi/p8tqpoyXUxW8zXM+8v18Mx0d0sZweCWGelQc3
zh5uhxYYx1C+fw5PUoMphaJHike5P3+xIEQ1AGfrJ8KaAuPKcmkKP3+LhGQKEng1
MCScuiHOJ1L4kojl9lzXxupP8FwmnsR9GeBGnVogrn1bLMIhaGKe2FVNGkmwXsdg
GFdsCAAInHPFiq7ykyVeADW8T9Q5hCanGv4M29TgQV0xVtUyK7f8Vr9YOFlc2sBV
eVIN0tIkMpo404Bao0V3BYAk84+KYes24OqmNDPTfy/GGFP/FDhiiy19QG+BE2H7
DsjWyHu9uvYqcCQiH3Woqs81nJUGLbfdjy5KzlBPbCbYLvoipJylw6E57+Nmy69h
VVzbo02c0MdmLHRI0eMp83QKHVGNCgwtsPI5Kve9Mn2txML6epjhs54BiL90LBLS
pqnExwXucQJ8jjU7jsjcJLJ15K/q08SoXDKThOIkrT0E6POKdpfOM+Q4+DOImkwK
tR8v3IdExh4FENcIwyTeRJW1WQUkG6AYhzFS5ZtCgJ/ca3/qx8fZ9FcHLmlTLs/D
DVC05pIJU2wWZTsQ45JX4/mbb+/tTmjhVVflY21YUU228quEjwAGPXk0ZV1lAx8d
89hIUg+fLK+FFGGTDbsVA0WX0RExLwb84MtbkUQGi022Ppj7hO5RflhE5zueIXFc
gLZXaebUGZuwl03J0xMP5QKc6bwnHmHM1C0RsxN7XbbLSEnVGZ09R2oqWG/Zv/6B
fyEL8ytDkc5cktmIbeTyc9tcTuEWrC4SyX4JICx9QhYbK4Mzqg1KZTgbiTbMGiqX
oyqvJLlgBvy2Pkh2ls/IoANge4vSUddGBJDR2mpzDM0Dgbr3RyqJHebMg04v0PQ9
opz28zJQMWwMPhnrQ3cRbqK9N4m/zr6kOFG5TQl1FZRfDNhje6uupugzL6utYhcw
Fgyvi6TD0R+9XJgEMXvVd1mvx6eq5SOKo98dsYU26AtssGqc/dZ/wPhkTT2IUhXB
XABMvP0fcUK06Tk2e4FiDzk267QN0alQyCf1g0Z4GwxZFMSzOhey4NtRdH03nea8
g50q4BQ+LnBYGqCZOsGJOTe2TrD4n/dP87lKqC9d5jz7U8fVvjDXLE+PmtFMLdOK
ayUdqeWNT9M2m2oNsuO9GtFHWo4L5MUu2dx1cj2TUxWjkDVNKGW6tBS+xxq+XTfA
/xPfLs86FK6dxpMEkffQykztZWrOt9l8Q+Ot7UWPp2g1RPiB8+9gGM8LSVv5yY+n
5VMqOZCafhlkRLP3z0evnRTBGCctyzLdpjo+EPbQaBvGMq37UKtL19ObDllKW0bG
TxrIQxquAwgEvaAdmI+pXBietJZRZamCTjrkYOaOHe4gaTxiinWj/GM1GpBWzkVd
HjtvZ9Z3/LyWU2VTcB0bd4OPnzXMLZw4/hU5kWnvddjjcl6fFqJ6y8yf5zAcd0Kz
0knmBowqGS7Lt2GPGX74C8KHYapAQvEpFE4V9DZaIHhdOsPv3Fb31f20jc0naDrF
9ddt/4cvj53YdEZf7V0rLNBGMqGXzJwyRhKp0ZYDCqusriq6CyNc2eIMFZmdCQH/
xX9/ih1mRBwETJwvEKSL82QuFV2xP3z6/AtaojGRH6IfCkDlFVZ4iTlWhLgN8c0F
nFXXe0YHWHbryp3LZU7b/UjJ39PtaIosqD2lL/eyleslYQ3CKKfFqxBtQWL0POat
0XiJZomYPJsoZgCARboiGLMhHtHQBQfAnTWE3c1lFx73KfT4i2p9g1WhJgoKtCsh
XMJM7zOIzobY94P28kkdJFMQdQZ1R+uCjvGwa6tI9pp4BHrNiezjl+qeHFDEoUqS
Qe9e+xQDPKYJE757JMgXyM0zqV/KnVHFfcdcRdafShWYDkl49VW5PqgySJYXcdmN
A1YKHY+JaKLb7Q6brdKR3oi+qnh2thgEX4w+HsYEnln2GPFmnpEhEFFO7J7tWYZ+
KIXMOkqPvSBvcBxlxHrZfJGb0D1b48k7b+fgArYjaHf60zCUNuAv9CIUsroQgUVQ
ldqwy34g13+xHrM3uT3kO2IuNlHWJd6s8nBPDiePA2jO2oF88cg7lkgXaH3MIYAG
QaKvoJ8rcUZg+oRG8jvnPSQ1eCzSKIVcSRqsO6jd4qEGHBlnA78Fp4Q0VbqW9ASY
5mKow114hzio5Wvxt75AUL1BLpv7oDiSaoq2vh99UDYW88Zk/IHAk+p8EdxNUUdZ
HZZvRoJAQbCnQ7yLvZ+jfiBTSgb3VSipTFCKVQay0csgDUVHny8VVCe1eZOmRFmN
zpIxLMOv+Vqr60JPGPtvdPa1KygQh/xwhyRbPTVw3DU1ZuF4lI+BdnYd130AaJ8N
Tjxe1l3R7Pp1iQoK5Rh2emc5PY/mSjOaRkZsBLXE04giKTW9gwA9XFpvykMGdywH
yd+SlST600HP8GHZBeLv0RRNJPkQWx0dNoru3oFIhONY60AJAlRbOeq2lwRmLhrj
KJ5/uzDu7G3wRvOonFcGzQLfl21gCnjiKHrVQuGpkvieJfTaNPE4n/I5cA5ZAvuk
b2FmkbK4sYPlJEA+z7bUPJ61eFiDy71QcYVBJH+e7XF0YdXEPTpPATxjJaUROZgx
tHs6Ne2fSjsuP7ETU3Nma8LvDoVdlK0Z5emSqlKDrVRWnUEufbsnUoHlP7930ojy
T8CFh8WGRbLepsfDPIoD0Y2tS7+BN+KV6SaUuTlTYaLjHsfQFGvZcoFiaC6DDluL
YkgOPhPlZ6J8trS9USCzYBcJXGvvF25ivP33bInWlxu7BByf0mplrwlF2GjEU1kD
l/NrKmRdXSrnIhhxUSOY67Tu9vw9+kDq7qLKeOOHfXfpU4CYqbPYzLB8tsPQzdxY
6tH7jsKChvI5BzkYguZOe9Maz6otXTjQbhu9Lna8mSK16IrkuXGUWWYy/Ggxb0yl
KN2Z4IKAy8lreV//mPE+LJNEDkyBP8YBvNepjn7ZNIXEJD+DfHyxPrWrZ4WUZDke
MVpSaTmB+lHvssulhRuqm/FNrHIwBo0oBCJWZp3fMFuGIEWp/IUS9tO10vqMPGkW
jBbhlyf7TlIBO49URHgZ4LKjSCo/k53Xrhc+n04bDt9Tlkp5RVK0Tn2wdHo3/bkF
fSg+uZE68hxk47bSe/VIutkysKzTn0ODQmR86BA1WzV9c66T4VgqdPDGFX59Uz0a
/uXvAIt5WoLO9krD0n8CzA9MXT6rBVjGCUjohMKOfs7NLNHMukxExY2cVWExRhaB
Iy/mo5MXVjHTC5AkqdMO8xzjeYFBxqe2LEFTBF5Y7sYUg+oRfwdLb8d82euQWoya
v7EO5kwUhJkd/hGRMiQJQbpU7TJhrwqwznFwhL/UGXS17rk+2MsZBEjPeMmbuDJl
ZkzZPz5gx6rpeaVrTJNcG9TPNICGIRKlb9QOi8SWM6Qf5bmvUR2Doy6+lcvx7m2M
CGgNC4hn0s8zAlbqclE1dmeJiFj0Rt+fuEqPHq4uzDb8r+5nPQw14jQpGtI1iclC
6gi0ETUJBHGc8K/Sb4SdEbJZQcn0DkAkzfiIJziv/MoaCDGeU0pLlE5biFUqLtTR
hwSF83aN9F4Y/eZ6+RRP+cciZuUxL1E3/6uKctejhRLbF9BMEt1Sl6tBxscUU8Lk
K90/9lYuWSM1xpYbHI8AQJZdoUI9p3LCS5gWBQOBth94ty1Xr1zMyAa+0vv+PdDk
/0KYIkvix2MXRBVymdjSrlHmQNVACI5eMxb/vmvLHVPyE9O7WhXaBFJJYyquD+qF
PaMkx/IVPxzXJdiUMqHFE8RvFw6eIGoDRr6dZf5Ndi07QlYQGMydNyXB8eA3fZVb
+9BPJj7KBTtEg8hsyWJmyAQuotmFi2FHvzsmD39uLUg+ac+A/Sjx1H6MUJBUsQei
2wu04Ae8C6kqslY8XQQq1oQhE65ZGWF6N0+Bwsz/+/UA2h3mhDzMmCW9y1t10R1F
D/RLkwiEKE6R5V30ZeLEh6p4lN7C9pJYQ2YvbLCNt+I8toLk1rbMLKIqNmhO4IFD
j+SUYpFgRn33m1qxckw7MdcAYrwym6fkEZP4V6ymT2YhDEpxcQ2u0zsFEGZj7oUU
XdnTBKkjPtuS2bVQBQgpLO2zI5Eq0eOOFS4iKUq+uEc373zZQs6XxqhgmPu7jPSj
gr0OypbXNPUAqbNMHk5R57hsxfvOUJtHQyWmmoF/1Fv32SfQuRundoLGJz0GwoHK
F9rEKSQJZcbY52wdMywvpKNGMokpSMhW7jF91O1JvSqcRWnI499ZVJgOTL1wfLWX
AInnZsWXIZfZdx0xBcUULfxU6OUlJbqXm6TcYnlEeu95Msz3Ym28+g4s8ji25jZ8
bmYF71gOwqqgToBZwh1SPhXf9lyJfKObGVwbAUl1lYh9X2EfGUu19hH3hy6kEFs7
TYpkYEy1hSsPC+WQcxiTRHWkkhx30CgQSUKFq9YuxeQfQHNVRlRXLHIOtSwG3YL8
adjAkZ5c5+vxDdvuHPf+K6S3FAbmO0ZvlAtHz6lLnqX5ND9+NpV9kwZpPHR4CcTM
/N6vqA4pMiEBn1xVZPQDowAIR/MFOfpAdSLs2B2Cp3B7B8ii4T6LlHnuju7E/3A2
hQ+wcmfBVNS6lIX2NulQzqsmjIPxIxg0KkwYsyPsiBsRsO9HikqirP5rG5EQWBW4
bJAejUQeOs60D0pUEbKsnP1rbaim7kBeUhqyWFToSGW4zA5jc3BDDzESqkwwYqMo
NBJfvWzY88Oh7HSToNNC3n/ihZXdPQLOd8zp+ITWqhAcb2qyp3kSvgxsl1aWNGtx
dcQ4JEPG3vq0j/cogTs6ErwVCnFPSGILYkTzkY8PBTxixykMYa5YqXiDCbgdcAc0
VeXg3chN4hh+cr87XwAzfQhAo36SlQNMIsA+zhMJzwZugVh7GsRePdnPq1LBVpWm
zntPZGQRmtjuKJMPnYZnz2CR1IJAzNZtO1UVi4E+RyqHAnNbvVoV7RohBjAWqNi3
FnrE/vR/g8FOyYf7kqDfriGyg7hr5SJqsRX50vkm++3Hx7jxEUDiOx0mlIbCwuWj
gOnTKbq1Unv4De4YgSKqygMhfx27+DJho/uKjmnajOfXMJv0UrP+rkAVSM1/MBnF
uo8wD3IiGXHy5Vbpo8uDZI23Sq+8FX2VC2WMTaIyV2ZiuGPO+F0VpV+dkG+jme/a
mZ6ZHEOB8wJjAnwF/Enu8kkHOFhRWW89IxbDfYC148fE4frxv78FTK8jKA8hk2yE
+YJoayUrkFz/v4y53hL9FEchzei8SncS2U1RoJtmQzpbTKDhnl/dvfN68CHSxyA/
RnTTH5VQoXmh4XAeii1/impdh3Q4chrRmelbigl4OhHiGGkKqaR7B9uGKRRhfmzg
f1RMxClA3ACVdhmzSwrWgJH3c6XzAbesLDQdZaHTCR2eiwJ+UHuLkSs7SeC6qQtK
i1vpMAakMuEzq3nI2a5sP4PFkBDbauZatikengJKJaLfvo+7QrKVHKjmVTkCRYwB
qRzV9NEhzt9oHkQjhNJB86+GxPhk46Gqc4OSde09Iy1vKVmb3MW2vzOyIvLWIU1E
5tkgAJBLnZJyVvIoJuu/LEpyncUepJcEEWmjteqTEUpzGYeUatuDBtQftLi3prZQ
NjTy087p+o/4ShXbAIHfNKRLelvesH/3DMuzTSwbwI01FgzGZiF6xJFKZRD/F7pD
J19Rxln/DR5+bK1aXLP4K2B64mI3wTqqzRwR0l6pMp61/fGxpnJ/ERmr65cCDiYQ
kcGSbfFihaq//NqXlSks9EqJY5DTa3sSl/XLQymUbfbp7u0gWNSMQDYbdgmEJPzj
P/kODDx2JM5/ZcJe6ltf3GV0eSQFI8YQaZ6fKbV3z/JTB5faEmR3gFz236nQTNac
ZVgpk3uaCkgPZZhsk6rcpbif0AHnZ+ce+WwxkoGBVM+m+/UYWVU1/keaVciJLWRw
wmg38yLTIy7nrx2jJYsFXMfhL9iL4r9wt/U4CCpHRimSRYUBaWtGNOGn4kuOQ6U2
6V1qjd2ZF46y0/L4vPP0MWobQBXCjGK+5/rb4gjGMchN/idqPlcMc/pFBLT2+hcy
FYzde4gLwLXS4a/HXnSMP3zO4yryOUQYBAxlTCHDpMyPnwYkVRKn8qx7ZF9zX/lf
SMJLiwAZI+XCDlvWz3VKNn1RPZ7yKKx/7G1mFjcNKAEFfc2HwbPGY2+CqFhSev/K
sATufEgdCOwReFNYvw3JYl7O6P+R2IvoHOgkF5ucgZWfcnwGqcrNTTIz4w3pZL6I
JvbUYVHbxwL0W+oxcQMDnBq0a5F9C3uuIQT9PIclCE0Tyvzd2iTrkve8IFHNjYlN
HepXQbWov3TOKfXu6hIZ5gdufm6SHSVQL8oT8I95PbUEVOTfVxdDGwIkUltogvW3
LsrpEbc0d3mLYnwvxrKgFeuNT/4bTAI1A4Ip0/sZ7XtXAiob/ZFzNL6ujJQZl2ws
yasgKJEGamnZFpjcuuzAG9yj6Ba65/KKWbRIK6y+4V1UV9n6RfbtU7c/reJIT9Gz
kRlJAmSDQWEkQVNLWA+U/tF9j9W1bEzCQaTOtI7pbOUk3FzDDmAUU9FqZX1s326T
k7CjUJGniCZYIyc6kKKAZ6up+Gczz9b1IOIiQXQ/iLwxBG8ZLbbFIVGvYOcDtWzv
hzpZ3Wcqp3+etB4fnpQJX6dYw7z4uEGXx92Fjg0FkUjDAfEcQm8mibbBCZocqEr0
UdRSyJ8tNZ+mA1XMnmiElx3bh+jXSsXiHszrmOic/8zXqCbpA4rEmiDNYwNpSf+R
h0ORmI6LuJZCM2JRBXwJTbf8zS92yafZE5kZ4KZTXSXDZR3hbxu3E7ITGc1ObMT8
fG5Cy0u/5jJlvEExNUmJaEQOfiEB2gb04deOHCCvu7c19WHW3slMH+01DY/mNDlA
uNzSW5omMqoONhY1HeDWb8z7BzyW4J3WiS4gEyQ/foBORajZPCkAHLnvL3Pw5+40
vKwgXlepay/MiyJcTS4KbHwYnatXIIpsgrFUS9fxbq8zhGCA0gHxkljeUlHb2wvv
awIH2NNMMLYGDOpTVnVysCCc4O9ldevSfys5Jrb6vWJTfaX0haS6tmhOpDHhZY0J
zRpzr/8W+BqgvKT4eQ9IwTaBY9PvQDVubdlf1GEMGKwUdJTmDBwXUtWi5L32/bJw
TJQU1DFbTubXPaEEPVYpxy2AKQuUwFi8QVtJMjHfY0Q6fxeFSUay49L5iuItB++d
IWhiMjnWFWgutRPq9Mpp5JbyjWGXKlSJLM6YU1OS4RzkAevgBiIztWNLcb64UIwN
bE2Hm0z0OWJRl1VV1uruLEQQK/2hdTArlkezN2TGcB7kTJwM8XROOsPKRl04aegz
yL2UowbDIkZfDYoM581IKTa9j6CqA//3WmhJCtEeJonHLzv0CQkaXTBEW+rNZLLa
WcC3FM2B4goCFtPr2ug/bFIVQ5zesmEVbsNSWWuir1jOAlRUlDdKmyg8Wfut7NKe
qhADrEQkyeH2+Ls1zzciEZkGvoHHhC+R6b3dpYHqyabbSnbuucqvI8rq/8HrMLoM
K7WyWCDNGhMp3ow673bbRZnTm2yeoqxlp39W7ozfsWAJLEkqD7vDOA7QjNP3sNCg
JQkNkgLWDpWrSgYY2B9uSHMjYFRzAYRBvk7PT36GIX0amZmWXp8/4rhy/AbP57m4
am/wVJnsG2A8yEz+wUdr8SNn2NFX9pMZXbuhAbOzfTXnp+/RHNDEgOKy3h0Leyya
vw9ilR60K11kH/WbLljSq/kDSDe2IxPyjje8rpIGE2frvWX968RJZLl6Vom8mE7z
l/MYFhi5zqa0Al5VsL+s/g/9sYBI0aBsi8hKidCS01zYWu66A8zk2dPRAAac+R8N
DcCG/2BGU56acq2CSLGUgRS1j0d/Tso9DXqpY5GyhHdIAfjudnTSvKk4EfQODt31
kT3edYSKa6H/59H/BWAQSyn59gqWWzCkEngBrs6gAX/BUAH7nqKMQqqH+HC4ghg2
2i/YfWqpg8NbXpEnGKvS11abN7SdztMnIg/0gkHfRrC7nDy0q53/A1k2vAZjakb6
/iUeQznR63AcJlO4yL53saz6vkc+b7XJnmuMshpqnviZtHo+aSd/8aVsPzX2xfK8
iSJcFXxUvUuii8GURx5j2BjkwuQnxiMeXDBCgiee7EQyIWhC+P4jW4PfQ56LAku2
fN2c39jBRp53LU1/OE9ssAoultgJidXoaWSWAxlqnYi4TjkJX4IaTPtcCzaksm0x
dJg0uqgiYn5nMqfP3+lmxX66V+2vN+oaDl/9s9nin4/L8d4I4vmTGrpVx13C4u5N
5JvOCtq3H2T3ZwRoE2jXvu6ZcsH95TCRG6b7B9LSGD4/+S5Pk32Mm95UPxGJsZ8i
ObeZ0mvoaFajQNZFqXEdX6hbpsbG3WQot4LWyvOP6i5tYpj0olHW8y/S6+UrKtAI
5c3EOKTfC+FENhONXrnzeDyew/S0UeuAdatj2EBgzZHlzgeS9aizkBR97ENORgw/
E65A9ayUDh8TIoGFptYH0r36TuhvXZxijkrx2naUTaWCfL7chxF3ZBGjjKrkKKMc
XkOsirHH5P+H/G86a/GnJQeN8PwoyPWTbtBEq289+GDkdxAH0dMkYr/XK9cp8d+8
VrBtd11zdmus8e2Ki0kW5EV711CaFFmIyQxZiu3op4zZTB+iVuu47PD0xx3iDEd5
MsMmnYerVW1Q/NqrZOLnV5osVDt/diUQ5LWlk1cj9Fmc/qKPGMCfP94N7yiMl14n
LC/mWezcF49FHxirb/xopIdIXeOuVquVd4wSxeR/GXBxQSPQQ270wJ9Lfkvh6uAk
2GflG9xQHDb2i8HTF2bwZil7DLvUBbGwig+7zi3NUNDLxKvHZlK2JraVET1LDQAk
eFS4w5HaoksKn9EqI+LFXyxAtzFGA0P5QPZTEw51mxJJ/So5yaYv8/qEVoz7NL/X
RPSY0DtJ6RKS9J7m9XKmfrptGlKFPsoo6LKjxZASlpwq7LCnk+44WM9tYUHntpyV
2MqRQyQs3iYZcofkQKvmHAFg0FAN2qQ8s+xnP9OjhkK7X7iFiYKZfCz3UZKOEZg9
iNuTxFvglXqPVrG+EEJ10pJWMCsM9mdhkQyv/PL6YENIGBViKOfJVb17MeTc0I9C
oXjI3mI0Qj7ErHfYtKHtpR6V9dvopNXm9OpQNahzSnvzlgE+uU0lHx2gvepI8PlQ
YD/7J3lRuy3rKvHQc5PMugAO0bZhJC2C7WPpWh3kVlufFDUiqadt19hg1DxNyxmx
NHbUpbLzVCgg1By3Snk8JOouro42WwTq+EP7KylzF8wnrk3oT8VRV3aaQzOdpYK5
lLwCniXnQ3I74JuGQ/wMpc0bwYY0/ldQ6bGgE7FgQK+ZiZ7Zre20bohwOYy67p8t
nBSz/Mdg7U9McfQm25/JhBtumr/2kngN7z5/ZRW60Eyxmjtcx23vXu0B3MG9/0BU
HwEzrqszLZhJjIpDHq2yaCiu8dVjMSpmT331hbeeI5OzEzD6ieNnh0kefdYUdAb9
LVdMdQ0CtHjmEB6TP+u8O15xIPze3ymv0dd4+0A6HKoKucZ0X7K1BiML3lHOI7Bd
ekyc6vVb7IdyyZ7k1lMQtH5maLohp62MKsOB4K2eAIBwA6EyEftgNAxEvE8LWDQU
KgTSJRwuDHqd6ob9k0aZqWb/3ZO26mvdwFY7tjZFaqK6Eg1ahwgL4CJt7guPzKlm
ssv5X7CiGeRxrA0JQ70I3WT6FkG4m19OCY3AIkKjpIGDgLSlQbMJ5R5hsh96ovfO
sP3HqUF0+YLdnbkcqY6RTTLm18EYKZ2WOemlwvA+q9g/37ZDoYbQn8szUl55oNFx
qJr1LGKlsdLgdDPBje45M1i0+hx4I4YJkrdgTviw0L4Qmxdd3riBOt7GWl2dGqqQ
a6rWbKC7t1SamMo3mAh05x6sOY8Sy8Aj6NSA/XNAXd6kAPg44eQFhGBT5M+q7xz1
Nq3dZ992yqq1Pr+UuEcOPoXZMJOjadege5cNM7+BgwiPvhNwfT8gXGk7/mUmNqpB
6Up9i/0T3UXm/9cW9UKnA6OROWeoH2jSACuEKMc9IYNI9Xp4jNjxW0iJMGl96IkD
wi9tR71Crs+9R5RyYpxANnoknAmZYrBroO4eOWUhwSjZHtwgH2pVY1h/0IZo4V2P
aH289nDZi+2eSH8+XFPqjOOeUw4P4odNYrUJHfq17ThP5NLvDtOqhDBGjSX0M/Jj
sFurFl9FEAAPg4WCv5JWc2isHTV2asqk0JXJFHoESGDEGCA90aZE6pdJ+WRouF20
IRFDnjSta97UMp6q9Tf5pP3nT9cmGHuT8+WoSuoNluM4ySYJz5/96UYgwjroazvd
4d+XGnwCfqfFj8i0lQiErP4MwRx6n3kG8ZSjwuzDPZrZfqWj5hnS6O7AVGFma9Lb
R5Iut0gqtYaGnnW/NZHi/GMcx3n/YAY79BGW3s9jlC63uswsMgttpmpQjEIb/+eZ
5RwSPhdmoHQLM3mEIRnadI/5CdcfDHuZqZQlw9vEK+e07STspZ2A3XVJjDPtZrut
zvah3sFXcbqVcVJerQ8qn7Ka7Ivpwbg5ePPfn2VzNqyvgGj7o//zbR38SPseujxw
OD8gILXaY0jBc267DkWbJz3g1zvXPhoXZBWyZ1CjfU2qM3sW1k1aTwIiECB0dTk5
/dPCHJbgzCgYZoSEarCiDAWMtkrafXQTROg4Mv/bJM8O9jk8nQBdHD3P6uJSYRiC
gaSpdkDHWctZC2zXl4QAw+0xCETh/MIx+7AmzE5Q0EBwq2mJnCW56yDRdpuqPeKz
O9w0Leu+iGQU9pCIzlfhrcxf6Yl+0Nv6Wq5mzMPC/ls+YxsXfW+9lK9doVvdY9Yb
n7g4vmhGVvqHwObSluhCLZfvN7l756pKDA0bxVs5wDAvtdd6cfs9mnLA+BIiDrcV
vOQj3PLtOMHMLVdtWRKW9l9x5MegVnK4g0wGXFW0CeQpBcgEdlHIGrw6VrPps+Ic
emhRqqDXJjKeFpBPDMMAqQPYkgWlsX0Yx8UAXov6xefpuib5w2Tmv9m5AhIX4U4n
7WnPUvuxzWJ5y0iBwytUN1LgY5xhgr7zbRXkxeE3nlYEnfjxl1D3jJO3GRvslGL/
kAbvY3rul9AS8Gvjp1aX5J9NfntM9ptyKAmTHTIIPTZrnbwYBz6JuoPMmsGnL0mL
W3KsGY2YZzd8iUinnajynqs7fxPSCEHxRzgC09Mql7T1KyVuUvLu+oSZkMZ2xywF
gFPJhnVHTkVhQ4gdTVMWgqatDkj5UCXYVYNTNwbdg7nqyNRCwn/qu9ImCErqNROV
cWMdQ4IkfFTzaFVctsCABJqXQUQh1whR6C9pqDEGgKu2MC5uKHtApyeemhZdjK36
xw9erqwj9jMTjRNOSSyJTI1C4iK7/x1fixZgUI5hn8/5Y5MZXLEbRn/1FLq5aiA9
JZ7Ud0Piz5TKwqRHRUOr2gEftquT+0xeLM2JK3EkbAajwx17Ae36wJmyp4UWUSrf
izODB/Q0ZT0j2V4xCPZM2pLSh0eXR58asu1niEWHcTDZM6sYFyR/6vjkasbunY6p
lt2A9kfhCsOTHPE90Rcp2vxxoCO+8Ntkd6yQ+a7oYmAkfW7NCj5au9kx1avKTDeI
5lCufbJqmfqOOA5M5Sc15OURBg2Mh7ydF6Kei7th0fWBUsJPjvGEb1gCgA6vTrNg
ac0Bbuef/97w1ImsWQYW5M02+yjUaHcok+ibNXM3gjYwy/wvE8uuTM5nLqwHhAh4
+Cq8AI097eyWOQo3bwDicOmmwYxihf9jdMS42s+rOzHou6z+hYGCwtUabIGntx1S
wdJVY5eJ80ULBOvZ4jBnSq7CEh6dAiDwQQ3rJrn+IXxEfPyj2l7a40Ukm40wufmH
9M4+9Q7yQx8t92DYJfbVyp84ke2TQRokJMWaBaWdB22PJW39XDuUKclvUCSJBNvk
Im/svUWmthX70ctLdMSSPmbC1yHpglWHet6f/Ob/vyb7y6i+Bwo8h7j24LSvskQ+
IgR3ZMfgB52CtKX1/c6j9wDU63Gp6egbjAhZ9PH5cPxyMpb7KzjWAv+I+nPDjF/e
dXIws4Q1IzQRf0L2IYYQuI7dkP9whzn4/IfQqJ36PintmmrGxkcK9iDvi/UyRQzp
EpDipKQJsLQF2pOKvr9L0G9DxZBOtxIRJAQ1HwXhDOM3wOkVCNFTvgzs8RtUK8/N
D8wMsBfFuUEYmJDJfcZl8SP9u9WkcyYFwV8gOoqvGTsFOw0ipbrQNsTXuR6gJGrB
iOvSbnc5V3s06qYdn41QzUZweq07F5fdUpAiiKc5PGujg26Y1RIvpqqzqfdUeu8c
Nf6FHFDU/CxXHKrS9TS+NbOLTK7p5grMtIIAsbEnnd/5xWQ5TjRs0Iflu2UXThz3
slKDfV8Mqrqk0aaM7qnYuSYeM1VZ4R08EhB9vjOc2wLBh/cj7BvIbGk402zzYyY+
p2mSdK1UspXT7HQouXE4YZv+ys/w/ffcxxjHhrjcGa/UxnG8EFIn0+zsrNXxqB1+
cGzkL/BZCcF0SBoLAFmsh3u2wDziTHTzW5QkE5RFcO7mFnawMpNUXvpdzwRF7bJv
OlmyjQYAuc8A4pF24vmhGi0t/LPwlCyAV9JUzl7dWEC3q99B0POQdejg333Pb8XB
Gnk1fZfdLujNeappad2tnTHuEJzPz3b5pRGODdTDJ2MJGaY3lqqp9VaQnhjfawdI
8gOWmc4Ley+4dm6zEg8kkDz7QBVnuDWpuHdDMXpQmXhi0HkbNBqFDNkk9MomakgG
8eNbwRGzx/p+Sbm+dbcqEK6n4DpatqwBGpG5fLQrKJYFTjL9DDmDBNqU/rY7jzXK
QGf7bIuKSC4ryRt1u0oNIgX5ZgNI4n51iZzl3suOH342ddRvt/hsQBeieZKRhJ+n
G0nnsn9L5nsq027I4AcSN1PHWCJ9saAwzvj7EOIjPJTmECRKnL3E65JyiPIfm+Kx
OX1McwqP0soNJuSAsewZ/SQBmguvw64imj3s2OqgaukY4COf71UFHM4i1wkyjL6Z
xAFPhct0uNT9pYeeRzCyxgQvs84sQJW4y+89vTujGt3i0jk+VexH9XBMAPaY5CPA
+P/bETnKg8gG5z6YeCpsLegPXgWaMt43M8kGxM90dPLoGn07xEoCsRGXaOrNNh1z
RxApPjQIeCWp2ud+BdDoI/Enjm+yVWZVNVus+t9MpdlfcOQAp6B49ul/SzfqbJeG
skGZxW7Mn7PPH264AN328b1LBR7NpJN3L0kpUhkWLe2haYXnx15MPqCBxL9t+jee
PAsqv1Lx3gnVnkwhh5oo8are7Cc3FhWiAxO97q+/TzkFhih22eML+Nu/okgbx4SQ
aWaHb2NXWm5t62RBbwJ1jZ7UjLMTvdUhNkBxUu5Jt5Nn1S9s+LJvi4rZYXx3cqYG
sQ0P+LaDv5MoGf/UA3Ja1u7FeoFXquBdPxQj2/upKKDlGHjnopRW95F3PJA+MUQS
HoKLd+42oyolCrGVb1N/UnH7I6Rbk9blTZhisBHrJMek6ljQO/vnCBV5V0HKXqRU
1LiwSFQuJQYg3kOW80GmS0ayP3FLys4Ww4UiqPSs2PxSzh94Zr2VKp1Qi8GtOCy5
xZMqkZCNvQMlJLwUxw+v1+s5h2CWnLZT+wvDLtz7Dxb24dsdEOWlqwiaS4xLESDN
hbFbUmHI2mknL1ofSOKjeW9cPHMQfjpdAXvpjzIoQ4fjinQzbfvI7Phg0HAjoZCn
bmu9bkGpLJz3S3C0mejTT1Ir51mCWKiTjPRgF6fLwo0Ei7YWhhCfVzopd0C4EwgL
PF22xxQAoOQj/QiUTf/+2wqTI65NC4YirmM52bOHCe5bVMgD0MYby241wtTg904Z
Gx08SL7qTnX9JVNVJL5VxFFUoJFe/VmDGcEiFTNM2OogBm8bFw3yQuvWSYGKc/Lh
hJJNaRqWmjX5ekt0yb+JfSO0b9CtS3q4ETyhR0Cy2LQ5EtU80PxUUr2JOQmBLxTw
RWRL6au/jNJb8GwqRhcb1K32iwMTh2t0A7rgxqetq4rmoFGw9zxQCv9FpkF1H8c2
U1Sl5t0dqwagX3suuvr9kzrT/cubfpO86HPVthPyO5cFJjwGg4TKlDZVAKkBfaSo
tzNWnbWWF8C6hIdCYebpBNnTcGaL1dXzRkRPT7jNow6FMaa76aBnm23zmwi3WzBF
VY3PKCup8PdQxS0dk3yJXJyy6mnzoMA5pFfNF1MGEg/xqBDbqGY7PiLHSoDZkUng
Pd4bfha3jL33+pSvILNT18vjbAdxWnT9flS71E1qxo6FHjVEGJTKYqqR4nmwPQFw
XHGWa6o0LizJveXyKrvIkvRSqyj81eazEUBYAevXWT4Eio8126j5ngr9ll3O2Xkd
XDMKiIuv2S8c36DiKq+L1e1m6Hl26L69+sqPuYoQbvSw0d+13Mp6hPp7dA+6WfT2
iiUdU1f4vd46v3KfaNMd2wmuSWZY+fpdqaID1BIeL0Ph/SNNWKYEpkzOrApdaFiE
ILplUXl5GymjmRuPlMBHOdioDuis1TeeEbOS6erD49qKvI0cuc+pTDBpPrUcD0Je
x1IIvA7HxVzcB6VpzpjkbdjCudwotb+IAH4VgCkV9DX52VvABgiR9NkPnt7ZoqqC
0tl3LmQmQY3E0o7/UsJiqiRmvJtfyM7H06j2taGmKj2vp6KZXVJ3taBlPhccQKp8
IQLtYHp2Ad2KJgEjhoEnasglDjERfHJHDncVua4hcD11JbCXQj0e74ZQQx/wwzph
Zo+2qJb+ymMd5zTjqdy0MMeB6dISTWVM2V2Zf/Z5ziXi9hi2vY3FQie7Aq2d829k
BEXoDyINnuQEa/MNhPlhbNxW0P4UFAtE+EB6GhqBJMHoA8MqwfjtBKYu+Yyu3Sz3
2k8j6yVXnWF6HAEPrXkMuBBkjkyNj1gCMk8K+y5so42nhyW5nSGdL2jrY5fZgoJW
/kyz6ma4MFTf8W/OIjLdE0zmG8zRqzlJnWKoet2DDpw3ZPLDNxpLoJpiqjAJdd8b
i64DwfRgZxoCdlytPXaI/kqHwMczanPHS4MS/A+UEGa5Yq5oSfayh/RdgwhvUa5g
Gp+/ZCHjDZgwhvbLdWK/315oVGg+SF8clhKjPui5McTGj0fzMA6EUkSMrCLLDjJ9
uYXWY5P0wMuEyKcVCBKDSrgOIrcR/iE6zSi5DUG7RNrms4HW3rhbyK/9Q93Vhk/F
mMY0hTu5YfbhFK+nLlqOsFcogiILWoCcZiUQJiOfcwieRz2RZgGoodQyQIASTw2h
JPrU0dAeGx/CO4wHPXPsCCQ8RCFOev/RRc9f+oDxrfqG3Kb4bXCAhcfvcSTNPZ+r
Jvdx9F0jNGWHOSrXBk2d8wJ+leY89EdTlrWJAkB+u+rFKi0+jV57H98glSzJFZu8
zZ1UjMIbpskr+wDPTa0KUr2k+r7mRyK4nF/lWzKnr98ZSEXICmNAXlYd3AuvMSdj
382KBRM1742sQ8A4StXpnSqk2P2odEQ/XoISxTmV9GADWNBuP+gUveRJ30k8mlGC
zBhykBAUcyjM9ILzN7jBa5ZRZUbZu2+3sdvx5US1tDT7a/PPtlxfj99vVlU/ltjZ
5htcr9Hl35hR9DZ2ARSiksXyekXoSCGInkjr5GkzneZxgzznNIl8O+1UM6a4Nkw0
2hiD4hyzVCuONZeoDYb5KmhIJu4X6El7tpLR9gvMv9oej4TDSskiflN0pe/6RhXC
iTsR+8s5W84Stwa8E43YL9nGQXHTpGEXdSIBHSjEwOW/7IDaTMSbwtxgmJvaLsOj
PTxSkZudrtRFwZJZR+5pWUwh5sKKOllfI0TOJ8YqM4+hdqJRLgdiU3i9dF5pQCxm
ojDR43N9AEev9BoIH46fFp1kadJ6qFdKdMMqDCWcUEqhOAqaAQPbO5am2SUv4X5+
Kphr59Xhas+IqSCpKhtSJCN4oDjr6OBYk1/C0RO3saHKo6oZRi9HW5rzGyVvjqeV
YjFGm4S7zluYu9kORviFzdzrdNPIkNDhv+vIkjU+rNYOoirQptz8xsOZOcOSq7GT
sFHkUr8x1luHx8gjwV4Uo57wAO7qI+vcdnBs9eHuOtO2Won/DOQrKg/Ih208HlnK
6Gs1DsDf8TrAWVgHCpmlWeWxBj50ubjrIgpipGHCwBztCM6MuMqpeMSYjw/vts5e
XNK5BFM/QhJrhzCm2vVNBLs2d+CbvnMSJW+gMs50R9KmAfD+uKmCuRA9xmlVrggM
o956F/TWZjhTcV7oT1XBz2M9fZmxP2+qxzvdiw2Oa+6ppKoE8nSvpPP3mZPGMQcp
xsN7JRDQOY9MjpYp8+mNXm9FL2nNWRXxkwMUxX7s4a0taDktRkCDFtD/1arlEp2i
25FcidOLWvBpvExbFodmivAcmyuPc4jR8+8iLGlPffm7hqpeo5ouEvir2nDiSZ9c
u3CTUt3KjI8fjnUPmQekc5R4AkqVy44QDW67fS2wEaYU8yqkZ/cGcjcejpvLxGc3
zF+BPqJ7tLMxlh9VXnheoPiJiKAICSQ2fwXZgjsK0j+aZer0I9wKf0ZyDR6ug28S
KdYWKOZ4cK3GGeNA+nFLCZo5Tum/1v9nCjO9t5iH8lGXMAJNaZeyRHN4AmpIKUwp
6Gj19OrKgsvMmIlWk/YGs97olNqxoxuDdGX8rdpmUvUarzXai/kydKeIngQfWgnN
mff6210LYgH/vLLBCvbrqt1wvKtIc5zcgYUbr/x0gI4knkII01hN8osFXYwg69Q8
jegMSwfo6R1rbfOdCFWNSxCa425rjVYnupt02gT87FvxTfJxODEp1muES2ObKA6j
zfhu0BC9KMLSeo4X5zLSFUGE7E9RlOGuHk5LhLvkv/mEIhbTgztS+WRLboWRfzMp
yCIXWsXSc7gxL75RwUMFf7Q1YOfbO9cIi7lzRZaOGpyvG1j01uY0V0OW5fU4I7c9
AdgoDIQiFlyK/0tWSxKItOtAHWVFHg6Oh8JcprrJxV/AgCq1anhUiO1i+gmgK8JU
7SgS4cR4DwWNH+sipmWSaANX1v5p3RKM8cx/8ldmUM53yksa5IxIBr8XMrJQvj5p
jLbkjfh3jM6ijJAq9RmdYFLCOkBLRd6DWoAbrPkMOQ+XBIBZ8VJ79FNf5DDXTvBL
5ykM8eWZl7iFQsHk05UK8S3qzpEd7Nh6veG6ypeBHc87s8nVpWGBtYNKjxhjXpRH
7xTHzlChELUfW1XaZOyAVq09evUDcigsP1JOXj/lpkuQsrWRA/CzhJwXlgnCb/qj
xTN0vNUa3+acUfnC3kM5ZAr41KDWvidM4dmBeQbXCWrFzQzWLT/g/F16f1Jaleas
8lSp/aFJem/1zTwrAD/wxLFLXRaOJ6utaYn83VxBAc3zv/XBy27rLh7Wa0cTEphP
nZjxqvE+E2Ba8v8HyvWvCTMRnqe37Bc02dMp4OQi7OLknOH3q7cJ8zlRA4BrK5oB
x/TEVsFtFFh+risLtQHj1+/s3iyX4p91wbkhXnI7emFEBOUHY050e9VgwJEtrvk0
4XK0KXyUNiUOIxa4jJ+Apt6jxk4Vz+5rHHO7GZUxD4tASxK3aNs1x3kWNyoP02VT
Pk4UHF8M0kEQCCFIyjUTL28nXlCHExexp68smpnk+O8cYHnXjfbSxIyJyy+drx5N
aoUMX2+BaDMzGWOO+PxYmx9ZRCrVtpqWQsM6n2yVczx6pLSTIukSRnQI4hmD6coC
0WW9Gjn9T3daLO7lL/C6OQHs3wVjpMIPw1vKdAQfsTH56520q2dAf3RelpgsRKs+
lNzi/SftoLXdW21akbXQ68cwc6bnMQFdOaMPG1luuZl97xV/pO2fZ2rIKuwfMvT0
kda/PmcmLYkgMPXLxg5gYfFQVC8zk6d+hTfJHGnBkPSVIyjnwhky6luGUOjN2x58
tQXn2BSycuXPgfFatXAhh5SL6BJctxUvTVgL8YKiiao5K2Aj+dQO9Rx5X9bdnDjj
291YlLL5xCTYVZ/10W8YeXeip7AoVhIkpvm7w2pJKjUzHVGH0R6gbnViLU/IBkKi
Mf2/7mORe3sxg6o3mqirENAcbqnSiWJQHctpVB+Wq3RWmjkyGVvkNFqYd3ZqeaQl
/Kb7hzneUi4QolDgAqukbSN67t83d8dpDXkXOrHEAa32y+//CE6BLolHngaTUF3V
PKWBtTukegCU5y+H6IaLk2x8af1PidmR23QnZHwrfCvJYWNEflPuXUjT/Eg+emFi
wH7ErWQh/ElEXKcA1jBM978dxQFZbDWW74wmlG6/5o3hfkcMoecNSi8k3Aaj+Cqp
vYOOs3G7I/la9hTjuTnF9ZrkkhEMQfe0Y+wWBBGnXFy5ZWKhYgCxhzJw5GhR96Th
heKGdavrKAM1NQF+aACGMti2tEuWjft+HHJGcnnIpwG1R+M7h2ovqGaJaeujlSvz
bJTX/vJIoCYI2Wm6DlMVGyHblRLLdYgPLiYsBFwZwEHR1b1W9kK5rOwuohD9aOxJ
uvNmNmNQ25kaUNi4gS14ZUHE9alsHQdvJmKNeIJRqh54mEqcg9ka5hLWp8gZ9ZYn
oSuVm1JOqOd3v69zDBlXeUQULfr+QspmGe5d6aW50tvuwXlYPU0Xg642ub7m5JSI
8JBKxTVqzgZqg0cYUAaQ6kFrP7a8+8H49m7rlfGFq3pAYuDG5J8gddlGUflSzpYn
+582nHZgjm8uKrrvJMg1rFIALb3x4Ft5wFZePpt9KGbzf+Neilwys8CDJzCgbHrk
3Cx4pF4t7l87MEeSIcGcrrURbPdpsfoPnNNcDG5jkaGwCrFBx7XjZ0910DybdeZh
xmmC/bTyj1q9ag0+Pz2mcLE+58fs2vE3D27LVZqvxMJeeEUweEYygzpBU/814vIk
Jw5LL8ghjsKCz3Kxj8ZrQ6zEN1ACHGa5MtQZj0JdnI7VPvRWVSBwO/P2cdSmTFU9
EPK4uPmckDDKo34iPEGv6oPdRR8DC6K3nLREKx01uUCMI3aCVKYAmiEAz1SIE1T1
N0eWItWFNys9tf7g9tJCHKjP2WfenWsI4e4o8TGa+5gztAhpYxVX7ddmv+h5TI/e
le+HiNcojpaAioW33Um7NUYxJ2ZdeODFNvKif3tE1L9YWa2nUpczWfIgO67Tv85Z
F3OlDUVbClJuq1Bql38oMP/cEjZSbGNSIQd96vF+WrZ2Hz+SBtQ8DYdMIB34In4A
bki12ob95I9/kPVEnLWvtjZ+u9gKCdBnFiwUQcuIoDydJN3ji11pxtzORO1EBEnS
LC55iMEIZmr5O20Ua7PSG1wFT/v8fQu/q8eTvo1v9IWWnK6jgNQ5DSMQC+8afWnf
oBWCuWATMjbqwxCLQjXZvINybWw6/O6dWlPv46zooOu+TtJ8WKCxncuhQu3QAeVT
D7tQmX2LuiPdy/qlSXwx36036ysnJptCV7K2K8QczaAxTJhGvhpndBTkCiLnwwmr
esueWhWeRyrfBFNcHrEiHjTbzEZJrvO4cnUkQ8i9Fqll13LCtCIdotcU6GuBk4EH
xge8AElrwdOLtoYaVBzymoGbH23dYtuw282LSvHrLGwOidQq1ei16x+feiOpt2TT
2alDFkD/yUySH5R8fSUILivRRQiUEpjfbeTD/DEYzj/M20aB+PInoFcQ1kogZOwg
n74+6nPc+yudDt92tanXd8NrGTHopoDoVaYVDjuI1LSPfnOzMk9lQ5Ua6+rd73Gw
3S7vslbSmPL4mssLP9dyNEav9NXgtih/J77orqRRxjJi3xTB5ojlbRObCgEGHOxv
ucAauQ6fyybcgdDlMPbnneb6SCZkG9I1u29oYyXm2Uv+hG5BCwEhftOxkM5swMCr
jykQpPqJ/XDEI6ZaDWQdnqfP+jgISGuLg4JvIW71wPv5tU0+UdF+BFflePHB5sCO
2HgGCPzQw/k205Yn+pwwCnLxiEpSmT1am02f6E2KUZf/lSEOl0suwhELuPCXa16C
FhnRwbKhHtoyssanUvLK9oPMmS1dcVAVfOdhhaZ6rlSo6h42aID/TH9LrszzRb0a
p4g7eTU5FYWhJstS8MuHZwluYW8CGs6wyZZFJz3lG5x6vXr4CdwtKTUfWA8CT2uO
bkq+2HEblKWcCHJmTEzOcZXWoh+emmZ8Z8zIrTR9sDZq1fw4X8j4ypDGTWhRq3cP
+ljEqkXEw1Kx0H33Htyh88S3RGKc/bWZfs9h3tQSbIwDS41Pbs5UNqOihJz166h6
LMmyUti4aEM54wjCxIvzTbJMruSBCFqvWECCrHituj+7pPbuadfeFIyT/sFxgQ1U
DIM+SdN/iWac+sTntPU37vbPcdPODDiw6XmZiDKpB0NjJ6/S0sXDTkNEiKBG4tx1
a68ltdU3MOykX1pTgutupRjzNR8fflb+d/iOKaCXPjuqQTqjk6ZbHvdigT50t5sm
3V3vmRnoVOHzU/oqDxPuNiOkDatDltuQA2xGTscxo3GOFIuQOtsxA0xiCX9s0evR
Pgc0a6JUrw9ss13izr0SvrzMJfW+y9Wf7813Ifzt7XBEkx8HLiX+PmWDufEAXN/s
Bvm46WgsNGYxYjGm0jM67C3WZzrEpPONSAzFOLXTWu/RVPE8GCcgyp4HjBNAgt48
EZo+HKaFx8KKPDm0yN65JT8aZ0azPVHeZzzWi0oKRwoiGZuHkltrQbM0sNqsYB+4
/bMsUxZPZWu4/b9gT8E+qOoJs9dRRMsC8rkjguNOIrfajve5+IWdp0npx9a6WMVg
lV6RUGIfz5hHesTHB1Toc2SDKcxZqiBcBAeXHPrTDUIBlHnUOhgcUBheBABsR6D0
bq6xG3H0/Or6wtzHW8QKYPupXSeq9Bd3IQXRbL2qatXxlnVT2td83rIH3EiofVz/
U5Z7/6UodXBwjsc56u5Kuz/4n7LVI1ucuNBo3PL1ghB9L8xhAFJ/fxuF0ZueFZz3
PIZ2e4NbZAPknQBG22tDjXD+t2GdtJ4I6EXBrBI4of8x0bF04XHxDcpysv2COKlM
WARKWpDZ2jITk4my1IjIHZDZ+RpCAeegxFox2VhF1ew6EmmDvUd8RL0gWVHxMeke
zb5asM1lSqZJ7IcAhuh19O9zitblPJ49YpjhQl1QrHdbpeqzqYGQ/GiCHJ0RMDve
z9ztHsthbg/c95ZXOc+64IdmPKsUhWvzxRJHLc8U9KGZXdzoC+iEA3pRgS6Z/8Nn
fmnSCx3Usc32tnsFCim9Nne8/oM1GhbFZ7qxOnzz5lvKAnWIrhj82eh3VLl8bL2A
LyZams+e9e1veACENJuIaDtXHX0P/N+Z9HV1OUYjM3cr6yhJP32yn/hZEKjA09LA
Gim0ssrTAInRYptvPJ85UchxqM/YwTf/2l3xYR+SI9u4FyHR3y3R2IWFyFq/C/Wg
/UNzmVr0YYiHjsLUd00cmsWqIYGEE+uXFtiGAj+A0PDiLRW+TQI2QQxf1hlXQVOa
tETcvHmXb0V0wNTwiR3vSCPincQXgwqSw9Aze0pcs9Cc9qqiuPRRdru6oj2gUFgy
K9Y1jWBfsslKDdmdKq4uyyaODmj7zm83z/20+i/oQIAO0uPDGJtVwes5lbzVL3TO
6v/UMstqt6xQw3vuQnghcKjlQBEfmWCm8FkR8JedgZsbk7t+Gmkavs+M2S4Lmowf
Osae6D7qBz2jO/ZdoFlZhfhaHfVX3Tx0rt1RxS3pq5Al83mxxQ0lfBoOb2vDBlUE
OPVcw6hZQ59eBdjrG5WSD9HvdPlBa5hhT87q5drm8isNH5P6H1Vz4EQ8bDThXUZw
M2ldFwvdiNIC/ejszU0Srdywkhn4JMDclYfBz4gUcF7zlr5TkDIBb71jjnfQARqr
JIGA1PENs27hKfjTdYpjxIlRWniQolOjWY5cNbv+cbox3tMllDKg+v7jxVISEMj/
696+trHlpJe1Av7b6P3AEg6KsgUSMivRLTCQ8NURr5D6teEc61xQkMXP+NKnaMaL
ONv7IQQUBJ1nWBBZxkEsi6re0nCtASorycZY71dx4Hyod2r4uJ7LNYWu1ImSqjYI
HBW7KwwEt1BrFOdiorCTjiobEqsWcc/CxVIlDtKmJmHWYBj5pY+LOFULMsfq3qBW
+r9uvcwSBao5PenQW076pXuXqjDyOUfn0WEm+DGbRu1RNtyRqVnot8MawnwLVYvh
Lci+rU0z/qTP4Sf0k8aJTfNFoP34Sma/080u3PRYVDfxcEgN27Sq0tU1ttJ/BPMF
PJ4tWaeg7KZJsIpUPE7SIkumJsoCm60RJcY7rPcy6EpyKX13Y+e1vDRCeoX9Y30N
APC/77lshVultbGURX4NiIc1bKANLQ8Az3JV+g0yFAs9SEuwkygt/DJMztmGuI4t
0k/tsvbdy1ct82gMpvwwqNqBFQYDvEGGNtKW+1/hBi3IzzZCGAfNeeCZfDcFAgZD
iyrEuQ3KTG2aUDcAtSbcnWJn/pAYJ9c+zyK17HtP/43dwidcUdj2wvzPOqykluGt
clTVyWBjXtjLQ2+mZGfaH/4VFkj4ZqsqVayZJBMQDhSDPg0K1H+d37Bm+mEzk/mj
PfvbiAFoVen+0mYTflWzhKA4C+Gd0j7GcZTZ+1beE9Bl8LnWs2iyCtCEkkID4Zmu
/bqJymc/12jHvMPvd4fOun3o2e6+HndZ++vNlr1B1uOVuTKGePNoQOilKm8G4sED
yWn5xNcar1QgwG5jMirGzZecRuJHZitObVTMBwy3UqE6t9/2eFcmpLzrNTXh5Tnc
by6TOTvowc9kNB8pLEgNFM9KZ+L8P4nPuq8s6RyV/eSnjwLGbrAGSDLsVCCuDNuo
8UlaMemyinJSsN9kvPCZGilcVp/CsmItnc6s6/CKHExpIrNWOD9p3fNOIbLQIfdY
ijrH+gAmMT3bcV1DB2rFZSzOliaGkhO68qBGdwUIwoQeouh4aQ8XsVAX/lu+UMUo
DPHFES7z478ipnWaAdoAh01kjltrU3eCTvw+r8twY5P9DayQAQpQxPw4eBY0xJwH
drOQ15yGCnKGktlfyFimefGgU++Bvut526aGss8Xxq8xglit9GJur8+CPMTnRRVT
7wRameQQUbFgj1xwHB+KtGoizIOY6VbkIV94s6TIZ9A3PQDsr3hs2cc9C81mZBRM
vpuf+vgZQ5IG1slPUPHBqJcS221VYBhaebYnjzHUuEjIHPO8P8ytpSqkJNhy4cNm
B/3y5zxxhRsqmWtp77ghQ7Id6vgrbPuq2Q3kSvsG4L1p4H5ztvMwV+6Wc75+pC6B
FletjvW8udl0XjPMOLfDlH/Y/I8uMbIowEF+lPlKa39XllQz/jNF/1844x7jxfsn
GKW29qWB5gjRRh/kdf0lr6et1k4e9X2LYcCSV0Cw4rjRnNmsABvVigQLOaeN2hKA
bzW5JBvO7MAyo9V7wtw2VKEu8GKTXqwfdxJGfiFvHRTkVo60xoXnh2pVFMyMU0lG
yDIzJWOPlRVTBsoKteCsu1Wbpw2IlJoY8hLqy3vK+DL9C3QM89J/N+oNAV7UlHdG
Kg/652fMa8qCbW+c1Fjx4B221slXNlC/KzhbhXmPHpH0J5mIiXpXayYrD1O/dO3/
D9kW9hSgTZHupISg5pqhKm+/cbD0TqPxAAd5QPomsQEp8Ds5gScf7LxtfU0LoDhn
aMcfh46NkDNKj+bqAqw/rn4qHlwQHd0X98Pf3K/npp00g7Afdge0fuZRE9hxR4o+
z52fM/z1mmJJ8iSb6Y25T23TUUhJHho0JKSWgzxoH1d9vVPyX+dKc0rrdZKrvFcH
Voh5f5G4B/sff5EkKDlkWSNAQLecHKGsPMAM2mDe+8r7GzrJFFC7yqugeqX09h0u
/hE/uEXe+vTpTccD/IdL7fNEEQDI1R0GeLOUbEKnYLhRXeXYAFfiNAjQmOFcXa0+
XsFe5C1W4496BPbJL+Whu1HD2+9WGCrbKIdM89JVSe7M9+kpl5IQIfc3mp8Ejmt8
RlOS6pT+cxJKKkwPxH/4cDSikPNn9gX/57MltdmCScTPvcw5fgjetm9bv59dFOCe
hLMcZ/0t8M72/FBxjWhLrWSxULDVjqgoFEH5HKhZofRjzFKWt001BEnIQB0YI0ul
IS8E/9JD1npy728rLo/ftkjiBNL/76vAluqym1PBBp106gBbwyQtZzcdkNdq/Ep5
oCZbIMFmqNBFvUDCv8yrLez+ovPgcpVbBNPup/XvBCAzO1l8mhWXer7IQfVbPBXu
QEMA1T6kFcJmtyStUVsYqImIazOUrJ2v5AJnIjPaOyAFohNXq0zhpMG0BeJNukhH
RrPq8zyaqmo5HIXhqZ0/5eJTICbFQz0Lr374MRhZ65mwtYlW4Zr+1uvs2ZLxlEqU
22IPFZnJTA4GnZ+vPSYRKevIkp0NHBb66TvzVnZkLI/iSZNs9sgDH8UTOu0lSm5q
NAeANhif0nzSXFJkSivfzq0zdf30Owy+eQlpc5brQyq6XW2oVc592J7QYPz9i3FH
JQ2g/f9uBBef6Lux9Ez+BNvMbu/Bt6beKmckbAV7eBt+fDogTh/7NxqTOqoercS4
NUoiFgr0e2CELu6fjj0dDN8r5X7SAk6O+OYG0ZlfBB6h9O98R7bTGbImf8BqhGsL
KaVTaU0l2q5ff+KCyUIO2O3Lqt/sId0oSaDpdhKJEoAHa5bWZIyHWj2u1MxxPnNc
mLR7qj64YaFa1ruFMJOL/6G9zXKKN6hArtfXpghoZf0QBNzDg3klmShHXE9Qkqtb
5U7yovTRIeGR6tL0yYao7X0WAAe5jyHgNryQ/fCUTK3lEYD4Q4OLSbXokWTIyypA
uyJoCPeQ8UOdUrOfsaxbuiQ9v4rp2jWBBBYIgjCYCzcjiEcWGiOBthIQv84s1D6G
ZOy7jHnF+Iqq7Bk3y6plHdc0kztfX6bTNtOdJaiTVNniP2FYtVCg7uanKbx7Wxd8
B0GK5SxagB0731q7/d0OPUevi7FfF5QO2xGeGtcKnE54ymZ2CgkYC8mzSuSYD48T
JLBApoZ8ZKrYTvuXBfgm1vN2sZ1SKOVOVFGf/YpmcTzLBIkSpCibD/NYBoyi3Y2X
LjjPNHWLs1kuqAcWrTjeDNVZYFfjcmU1GnV4zOGTyliLQwHZoHRukXIRilBWu3X5
yy4VvReh5dO0mWXxpXgajIrtphymP5k/jCZKj0dK/rWH3HyV4GXaUJlLfG4nOCsZ
9AOfDII278JmJQRCfF96kdvHuHfZ0ov4cD0IQb+EgKrNcBR++vqmW0A7AJNdqSZz
OW1KN0+AiYY9fU+kL8DisSpJNCGcx2zjAjJwbcHlQqLv2y0w4H2yoSie5L6pLzR3
iZQ3ndoIX+aujRj7oV1KhDBFUNIixtOXvl26R8yQISvqL2PCskslbMjMJ9pFREHl
ZuONvvvwJimUgdMIAD5FWqNq07OODGF/Ma2ZQ/7ms7WYjD5YeJ6e1onDGdJD3+Aj
AEe8D6gibnAN94mXl2yoah7eN8YihaHEloltxWZy1IpBjM+bGgQhsKl5FQ/1GxSw
oNeZBsX9mhLbbwVv5IUd4/+RP+5fcF0/NN8MQxlfvSeOpaGWi0tg1hc2fDxQtBNC
pIgC+ST50Cp3MMfbTCSNciyX+GpbX2kPL87+Vngc3l/AcY51bxu8bbbNII6Lf63U
jk0uzpSPHGzsq5DX5OWOJa/PTRXkUM7MDgmbLolQzOLlGzlNcm7GUscruZjB7mJe
Xod0xTJDDqI83fMDZmfCK4MZhFvxDJvSUsInCtEHNuLrScwy5abO2sl7iXsgaoOj
FOenzXwaIiyROb3LQRP2HXfMm0vENBzl7m3AvkRe4vt0VFQL1/61WgmtuGzZNP7b
3Heu8D1XF9tfxdHhk4tkSN1asfm+u6m/w3pz4c7TcDrU7r60dINJiRabZAXtYi5r
RHa6rUEPrqY+kfNLyJhFaRp6tfriltKDVt0CWkeLu5RbFX3yjwP5fSvm8227fPur
C12DquPfRQTcDDbfzvOFivfJnADW3vhwwDX6Jf+fW2tsyV0clFLA1eWaN60GfbzN
i87oTZpOWSGB7uyWpd9lZbWA4meP+FfSJ2ppgrrOxgAs04BW3VL0LSIdhJ25jTD+
gb+WBxt1WNsbNYbZCYbB1XwBoJfNxgLpEkaQWgqIw7VehwZ4pgjqa2JqhGLuB7iI
kA0iA8ztw3s+fduGmoyfbf4nuTLLT580qR/0L2TNejvSeAwA83QAnNt4wmt53beE
TXrGAkdsIGY4w2H5gaEzmAZPpOwcICWud6Q7PJZCMTndgnHwBZ9BWg+LxJItMOWG
8Q+I4moc9dGVcQpMB1LHwc/7yHES5SNX15UexYjoXS1w6hQFasdpA7SSYmLWZGSl
HRvCPhQ4xKdK3kOSbfcouDG6xsl5+ucVGBHKx4+eKzBL8iV/R6Y7gbGgetXAmgSC
Y6DD8qz0qW2uM5WU0eDJZARdF2B8vZclA3d2iEcwf7lruIjbg7L+ICV2ReM0ObeG
i2puMwqe73JOomAo32okw+mGO4IKoHSwxsMKUkRXAv2yT8r3idFmBMAzuROkxyVB
wZcywEN9UMpceD6HilVJuOxUN3DxXYO1m+HBowen7t6pqzr+AFTzuSiHhdsPtqNZ
LB0uOXWFfz3UuEz7igiKx/GY34NkpTbOwHhqrCZ2azGecyLVtbDn2x+VTNOmn1Qq
EbWQ5IRb0ItyEyofU/gSY4eTOErZzZR4fzhkcM7D0JIs1uCaxtQrp9lGnc+qoYtI
YXa8i+csAjBNAGDlFCAeKVSnYmN8yrRrpDNyF6ZeM6dsnFh7wIPX4HaPb0TRgYdG
5hrnWDM2Iw89Jb0ajWQKZN2heciZ6FOYbFWkXLZ60LnzLvvzfkpiuenizK9biTnt
uqB2PEaiwwwyXOfvLTUC6ABBt8dmRZDd0L7/bPis8ULwst6olgEhGGQlpJ+Ztydo
uu6bdXKEbRQZgDIbak2a0RSFa+bEuNBqiPNKM8dd2J+1eJrFwjHVrx3Mg/vFiq1J
jFrNlvWP3gRFHtZw8J60KKw33aFxN0dIRG4Je4xw2akDgifk/uO08N4Y6EFLcxPu
CpaB/mujkxGItuEwRNBKPPGR/W/n/ipj9J7c7k0iDUEitDxP05h95A/szEVvOI41
qLIM5MFyrcYd6KXlMMvF83H1LuelXan4N/z+VcC9dEEsrPnNdJK6EfD3uDwdw4XY
MldH1mcMDBzOuZsN3Fs8je0R5iimQ2NaPEZDeDE0AEoxanHUvtFWfwoSetMAa93F
pHOWOm2s1uuDRKnkO7gszqlhj9j11yJxvr3JTVdQgF1+ITIvOoo241Z//nr4/Jog
K6SQkuqbxo3Dh0PlCF43gr436142zhDTMl0F2o9LazBPnZvYpZHrsq6joyih4hpa
A3FwFN2ZVY6GVZA4B7p1HevXKQWL51nZM+/dgoZD8mSCXA223sCH1vyQ+ucJV1N4
+7aGDKk3iIYFzLwsK7UpDMUsYcDsYVw/JIw7r9ipiv+eiEHpLxkW0ppdJrbMWybC
AWAD5C/YV0BUARjFANhiduU4vFjexuF5mFKlJqX+a6Wd7RiA5YwH+cQaE6R4+j06
JFxyGGkiyU/TLb9j0ZX2bDXsljEDBZhVsEK9yKJkTlb8ZECMaoBVuqR2LGNIwBHR
DhU1jLDgNYw3ylBIZvNE7JRoB1AIqTOhvcAAQ86OLsT/BzFrHoasAFZzZ1ZEY3Zl
i0krmHFd7VcPTrX+XWJob4ypwgYvFKnt2t4GLMomeBduv/45CThj/c4KEXjmOw2J
AuhKPA/TyE1EXcZ9P7PK56ZfzHS2ivkzEHG9P+dM4EGQbNyI2LpAQkEtM9Mfx404
lwU3+C8FoQH5z9/dtDTniP6ot4PR4ph/M5QjXKSbcwVtbcHq3RCFUqtaBGHUegDq
pP+/8gDhPmCFGOUuYClab1+/DQTyR9ijrPCCH2EVG+AlkcuEphHSXn0Bx2+OOvqd
2tdb6kR/t6mKUceTVxBABBkpkn8p8WqIEXSXhimvWt0Z9c8Bjv68qTA0RINN3EBs
dtuZ52GYL5ZGeRgVrqNBaeIwX0QlhidVT2F1LHryxfl1t2k8NGeG62m5qsP1pDaY
N8Ua+ZfkKsaZ0bjZimnbIfyQosnZosinc0J03dFITKLoyPE08K2wD9uQQB9+jd1I
rnzFaa28rTF1kxT6FudBY3u7lnJEsU3oAu+n+su4QPcQLRSmOuuM+Yo+O+rZzERc
+xiJ6dqYgYlPR1DmZwoJ/EgJwXz5PKVV6ekwObH8UYjcnlTYd9w6vSr4qjCtpNpm
bEtCt5W8noI4YF5y5tknlF1D/0/5CO++F9fmmt0L59z91VwRMMhqFXMMYJviUJRl
bfzZrNMNbOwlm3N1qMF1bExBsf43XKOpnxtISf/LgZBYStiGygN5FqEvnT9gY8sB
xK77kt3ktUPpWPb8TFoPElCP4Y6sKohPVlWGOys7X+GdV5Ou+qAQEgS6bAArIkcE
R9qjgmpbyiv5KUv2nq4N2oqTVhQsD5gCcSlHCqS4SbCVUdZ+eJgQSWXO0MjIjtcG
BoBgnzvbwyf5lsUvg6i+MpJEMa5Xz0c+yYVXuldlJ7FwSXPdues/NO7y0BsurluP
jALiL0euQS5jJHAU06KznpVygOGMhIqgtOwm5AejNGl8NYsAGCKZ06fosj1/xu0i
potV5FOa/LiYlIgG8bPX5BgKtSe4ffkqHxWqZQTqEqPzwAm5MVjKsas61Rzpj5Yc
NFPIYlei/B1EFzBxwq2x1V7Cyr6xnA0681/dFo+mHp/hUyNcBYYcQmw0ryfo5sEu
H8Fd2enGx8HHUw3/B/wzvZPf/4ptvF+VfEI9t4xBMw8AZmxGKhFAQhYasVwnuTo9
2atMYZOc3s4sXUGFhlKNFLnnLqkOGnmAzYKzPkNZ8ZOyUKv/65jvq6CNJqI+UbYK
idCXDtIVYrUIX60qm/V9p60gpxStml9/d234f/Au/b2cAlaqFCGoz/WKil+GRLvA
eeAFfGhCdTtjIU1p1nf6rJTXfMX49qVOvWt/eb0+ItD04opFXWadw4Xk0P/JXyJI
vmhpJYbpwrDY7Lgk4fs8swaCZmmkGC+aqrZI3jjpNLYKHX0rBVG+FOuhU6QrXf+F
Sc/Ch0H5TwQu8Fd6USsccYeRhPWbHXjOToRXQ2OLidRzttZpQ9QbX1kTPqfbJ88M
XybS9t5c/C7c+joTHYSK78rF2dHM13PqQCx8DmyYSZqjZAzvOMkiCQALbAFqFkYZ
PHOqSmXWJKypVMq55g6GHXw50Tmotduy+UPDRe4DfvVciTrRvP4cH/22JwcKG30s
nMdaLvnMRY5Ky+nb4+3fccymXlbjF2+RDn1WaahU+4nvykNinEMl63Jle4b3Zfy6
uAniaHQK2y3FGlJm0ViPdU4Hsma+d8S9VdK8NVxOcFmnlsEWQQ627lgsOnkU+m/5
FcXd+W7S7epLRIyJyT+v3Wi1EeGI6Xtr7iBRKY6txgV/Jfb6vzrH/HyUIlY0i66p
02MFEGrXjhIyO2kA/zHb+FyjY8RWjFMSJQJlr2jM1m7IyihwDmIs4TURVKbZEaWQ
anjlUACGTswnH5PgIP57wdSdVbCBi8o2oRZYuvc1JGgqIH5G/9273xMMAu120CyL
UMdoZnlbDukmd9jhcDlQvGIvD3er8aU4TkQ+9tvBPe4KfU2na2zLK9r8G5ZoBhNm
PJXIv/6/F9wn4DaBe9fHgy2N+nzGMDYeFtmq8s+iMOiTxMwkS00Z0VpBdNDC2WH+
pPw9nXUZ6dRlnGyJRPTpl9GTjmqh88W9wr1zro+XeddRYF2dGq2J3pdFa+9Jr4ai
C+p+SYz+wQY1fjokPNT6U+HyRuCshsPqU6bZmw9DxfClbtj+d7WNhmmVehabjPbH
YyWr/pCIes7zVerXOZIHViSgH+E0PNWZ01X3lqyM760V7i/tlPw3K1kaTK7H4WbH
bwLP2nPMfidAMTgjGhPyN1FqXj2Zq2+KYVGq2IXGBmJe7JWkr3hxlnAmfoJIFTRG
JFnjvh1eKadAOhk+hGHudmKHtsyGpsVPw7Ij4de6jJH8hOPhJC1hSCUwlgq/hmIy
Z5opoLGl1TttEL2VX53J+ts1ItG0RdOgchFIBQVpUNlAsmNJh8fLxvp0Ajp7HguB
Esxr3tzkZqmtFAK0/0bCtko0LvVgSHednuUOPh3qCax28efhLqe1EYGhX5CPXdH6
ZrUVwLiVxQe/48k+TTX6szPyaaG4epO9WvJ89n8Q0svZSDPtqpKP4kkyRuJ8Ti9f
W61B/CS2eA3cGTIc/bA3hEzVlmwvYRTyXqI86jMpsqXfD4TSgblmML8clzzRUXKY
lI/lB1esTcqX4Fm18DNP5Zm8B4LCdt9lNkJSZzSoSwQwIyO5ZRtaobqW+9CoTQo/
hsmvDTnU5KZ6znKPs2vjfda8rUhpg7myEf3IdPgvrTZ+71w1vvjfj7eklrPfcV1H
pnXpfVfQRXFrjt/36L7O8VSWBkf+7Pa2WIgN9SY4HUb8R0Rr99L1ySgv8UfvoQfw
tMcqtVLQVvQ2D3UcSodGMUjfjAW7FFojFGQZ51ovBtRRRc5ovEfwhLvDr45C6iN6
9P3F3sj+f6+qXwXu0G+QK5UDuUsvys/E8TpxDsNJ6ushSACZF61rWOinitZW7TY+
pCsFpTBBijH0Z5Z+R8JmJhH5rwoRnhv8tXRhSyJz5Fk84AM8lWE2+y+/YI178ooJ
WwwH10ZCXqo/96MTkiKBcLaWhjga/S2XhOeCvlB+XNGtbkEgkB/ASb0GZ7I8dr9B
YiT97BomR0GLpIU5cBDGyQ+fjWiuP3nFkqY0vyCVdSH6aP8vRsMzJwzTLtmbUSkp
1iz3NYIqbMwemNdbCAk39z+acQrnpouMFBzDhzjjUr3VGiXnN21o5Yvzthl3RVtL
Q12GNZkupX9FM7tkMY73tbAtWT81YvKsToZJboWV/ek/5MWFR9rnyHZFupsu5Wx7
hx76egt4MoOxgJaB3/2nr6OL2pXBrWbiO2Sw40RdBLeL+JLjQjF7HQrDXdcot9J7
12966NKff5/URwernGtvpH0m6AgC5I0fggWSV74+fwyGbvVv+Y3x63rHaHQ5w/kI
c1L9AIF4ZBGaTd/gFEJ61cVZKTvibHL3ewpRG3LLmfLS3IuqK55CjGfkz2VGP1YH
bHcPZEIgFE8l2eY/+svWvvoCWYKzyx+WlL++dh1kILvsTdjxsPNV9Lw1GWGq7BPI
AMqP3lgOjxtonAP58tSoPFEgIeTEWNbVxuodHEcY28w1kqXHKnk/PACJxZLd0Ktw
Pq972w9xYf3iZyCRDwQ4u/8Vc6PuwA1FtT2GvSnsePOwEL+opGbX9lOJrKMcXvo+
aWfP/D9bxPNfhc5E9c2JXhy8101wxCcu+SDPtEbk+Sy7rRwV4sQ/M8XovNt8kIE4
gz/BiRAvhlhOWnYDbo2y47w925ZwwsfJD5SrYXuYHxo8g4vW6HIsgAhHJaX+86pp
506Izid8dr97jqXZlLd+c9j+QwyOvs9aK+XcdEzZIT3bG+axixlrpc/YoMId7ztt
79HkMMycTGA33f6XeCvWdsKZ+2QyqcRHsD2PeWK1PJujdFg6B+jkH/c7w2AsCG/P
o52NbSWplcNWra0w9hUy6i1qG47EjYeUGlL3PcI36/pavtvDdvAiKJQNrr/ybqye
mXWFBxnc3wycnx6EVLEUD2LrPbThoDXk+YUksFMh6nP2Fm7TTz1KIRXq1+1GJQOJ
Nb6SgcblHpFT74RK+gLVdcRrobTUEKP1a2oNt3NghWmHpLSX94OJGO3pGjTsndFd
Yxf/w/Zl2LR6WITJDCDAtwSIQKBcQ36yYUX+O/mPPmbFYo7olqJNB5/6WBSDtaOp
YpEKCxWbzV4hEfaBq9n5cK+krt6nsgM35I4dtiwbnnyo+OTlQKPNnVKMkY7jCjEP
InZ1CjEyaS7j1DqPmdOx/6CHjp0Ef25n4YBep4U3hiuV2oucGfmBl0j9BAOjgyXK
ieqbEQZT68FGte/FvFwNeiMt0uQHPMsmm6ud/dlxUegslUke5vP3G6eYE70ezWEY
vjILDPeRXedDpejRWCfnR20j2A8Vv5tqSUTzLBG6v0jr9sfkZKF4lUwAQ1clp6yy
c/kB1yQQ9wTeQzox2rGT4hyW8ntQu5vvVrnTlESrX54Jmyk7MkzcZVbCZf29FhTk
is+/NZsWgNCfNVZHmjfunbFYJRZRHBQZCOwsdtmsRKnh1RJtLCA6/EQZWP+tBa6U
t9zMlatf9y4srO13Txe5hz90a/ukIEsPCKcy9JlCNk/k6iQCVjb0689tdq0bGI1w
i5Pv7SXUgW1wVY4qa6DyOdmYPTgrARO1Y5jNWNxHOa8Vossy73TgxsbfALYcbpMo
Uo3wrF2gMqoDXdG+wRVxSNijUVG/BhyfblseRqVsEatKp+I4pT7UY+ltTuTDymsq
xI91hBDls1HgMXQQ+2OgZZqa9+NEud7eJ8MB/4rULr3dlfr9EBKlCeNZQ464EgcA
43/urMkYcQm5JfzAtKJOqIfjfJJaSu2GRMvMxcEJfhEoCivOB0f2z/JGO5VpyyEO
IJKZYRrmzp42n2bnf29Lc5y4ik04NLF/xn4l0r/C2eiCCWe0idb7GTapXWD19faX
gmXRVaZ9eBlnc4uxmoFAv+G/DmSneh77AFvtioy3Iz70C3iU6KJ2hO30bReMxXnd
Clxtnh2iQKUOMQnGLB124lwI+M0+yp4EGfUq4wUvx8WLKHZfSmFT0CDRw/0wMLfD
2bPjgDxnlP1iBCIcJFCebZhxjNdrIMG0/aV1c30+v9BGGxxe/7xNUoabY7QHOMre
j3gYb1KIQN4k8x9nGcR/ssot0iVfbksHZT0D9wAlUNAJFJzKrI/k9qpR1aQB/+wU
UYUHKAJfYzSzdbwqRcQst3YEdPMM/nKlq8GUMDF0Wprk0NC2p+6CJ0UH5+qofR/3
Zw9BG+JaoQg/ftHf4a1FFuXOAWdmrCtDm0NiJ+T+4xxeAJf/3uvHzINlI+KxwywM
FIHnG5QJNf8vhMh9qBZEDFuVVB5xFeWAFE+wcLdERgfOJTpR73++Jgw10W9xjkiJ
m172KjkEG//sYr8R7Pe/hqopOZkoU60TqKLVCCRHAaitG/qr5yGdqEJsyEjwgo0G
LrgnaohdfNqmp9itY12iB9A7lpjZhpLsc32YWtoJDGj/w2aMVHAviGEzrJOpydbx
JSC7gBeeSqqGKFBzD7ItQ1niN1tEQyiBUlVQhMCAFqdLrQ5foye6uo0VdsWTX1PE
WdQw+46Zxun7iHsDq14NZBaKIMe/opzT66BTTW/lOzH26LIaYdosWLfnHFvwRHZW
O6Px9Fp1cI4bOCIURrmIy1fawsG10TIV5ogME6hk/iJsBugEZbJXjUF8dILmr6Pe
iG7gKYycDi15nRa2I9wq+zTyNHmtDmEgdb2TGzmLJhryspU5CJQiKfVtqAWZwz7e
F7+9ZPBe1Afe8A2KvyiMXjf3CYKiJhvrmo+k4vBXCZ1suzfqm0Bgoq7e+UefwU65
yLY7NunZ4rdi3eKX1yDtVNjnxymVNAlLfiR6UfHE8IORlm01Fgb2N/u0xvD4KG4q
36qCLAsExtx13KZx8Nd3Yi1KlQbAfqPfJq6wwDTLYfHlgBc4R+8DvqWhtG+ReFdu
PPQdfJeHXs98VRWs9qpw+j0pcgUybiRTRT6mIESw5ZM21w8MGLNJXhmqezjvIUn5
z0XdMtbuvjhBmOBy1IkLAuKq3RV1RlZiIsYemhGz6T3zlIy0nWenx//zxPR4awS1
5H9/+J0yMdHMZo3gb2sLu78WoNgW7uPHPFWbWBbjudZC1kG6BBuXNFQIrd+RuLzM
d4I7VO/9DR4tu5RCpFMkKYOb72KBZADwtrpzLYK6Id3R+HXb4LGmtlVcqhw97FRL
4E2/iAE8fLu2XHYTg5dp5w2Oo70jVRzKlxIRS2Uk5wv2H+4c99fz5LZ2CLD+058g
ewpofKeCgywIXLkJZMqERGgZ3vhz5y/NbScrKdXS7yJS5yGayrN4xK7kQxGfUsnt
nV4e1HvT2HqCdwsfsMiTPn7A/9755EBPQl6KYTh8NJ/5lLZ7vSmFurFcEAKMQ+6F
Dr/XbaLfS/VNDJR/IM+bSb+b5d2q6qTriCdZm3KgTGapfcIH9GkcMBcUG957tes7
tJsuXrIHMmMh8NvZpk1vRLHbkIU6eSPEnYy0zrQOqF9Q2lkvpnrrxAzJ7BHI+YQ8
dPLybohPnypZRpJzqLQiuAZl9WJgCnKVwKTePsFiYlieu3XjnCeJ9cp2p+MSjxLc
PlUqwdn2W7WYoKUaHnUs1rRmW8XQJ4r45iOqZYVdCFjJpk/j/fzKfpzWaAj9IZrY
p22jF2OYjfghsnuEbWbh2x9l0ChyAzx5SK6Tji18HKVTwISGMELB2tv7hVLsyxxq
rfLVMBnja/e3oo8gdPVBEzIHzX4SQkYTTIgK3LVOlF7dwEWOpbQhMbewj/dHdlRD
WU+wGrX1JH6WYqCP4cBtuFjtqmlz64bq1AbvZoGVCadrQXWhetBx8MwcO2DEvZtL
o07O7fIr5gLIZ/oF9RbvRMewc7zdQ5ZgCzZKhyHuwDdyNUF3XSQGRkW5RDQeiun3
oFrwI12es013BcRE/euUidJ76RKM8eflQ1UD5TK9Mnz6RBgUKAmeF/Sc2V+TzZiu
QHEH74qp4wNrzF9nknx24lh+VSwPv+/NRXHPRvaZm1JS8Ea49obxuoI4Njw4I2Vw
txCGuxgTMc6hHTgjKJajh9KVAtKGNwXdyIpurRHDFYK9xiZf8pJe7cls8OYMO5bq
DYnsCFmsMZrzs4RWV30WcTFz9KjRAQBNoMucboHK5LO/hMcKuDbG6oxOPEmFtgAz
yK0ye94p284nQvBAVlLZYjHb8j0hlDdazgIw4Z5hBB0wt6pICEz0ANKS66eQwqVX
mGEr+Y4g0nM06m+kbA7F7pX3Nub9DNFoscoM1fhPZcK4R9DCB9/ooAoTrw1j952Z
C7Oekxf+pdW9fza07BtoG4Of/BAKMZzkmCoBfsECsYlbecRVdS7//vr+8zv9ezyo
gAqIFTjicxo6z21qHM6b/SIPCkYvQGZuZ0ZNiVNWh6Q6VrNni1L7Xy3J3evrqPi3
fsa/h6M3UKlzDK2dqMCbUNcjDxKSc75tbyowvqECM7s2+tdWiqOzt9Ok7M8xy+/n
ZM5BXrghCB9qOMkjs5pEUACcl64iZ+axVYA2/R0n+ICcRv1Xs5c0vl6g5SQeKmcF
yaseKDdfS9N+j64v5LuL5OdBgyWxWVsmXEWDJnNSxOisLE1kT2ij54TYlwiMs80h
/XNIZV2DfDxyiSc3y6oLRg3S7fzlNrwrW2rrIORml7gWLsRF9+WzeCAOUoxoxl0I
pjd49wb5wDoniJkKufpf5/W5p0bmaMf8MxOtjBYR93CMV+nXseoMFGvgE8PP4KeA
OpQ5Usq15w0q+ZgnrJ5xX75R8Ra7x5Z0F7BOAZ1OF2WxeJurriTg4weMpQlzo/P0
gPbZnpcWzwLJbXxRwQwPLaSIZg2V6f6eEHAzc3EknUPX+8qCVkqnP6XcB2DFF1N7
IW/YU6ZEyWeskUwLgnBuV333wksl4W88CKWck7uK4K29X4WvL7o+1Kg4oMuZVJZG
zsdP03tTK5/gzcDuFhFlEF8IQj3fMF7z/IGvmJKwUyWtsfDgUzuaStDvqWoRzRfs
R8x1hjp8v3DwdQdVXtkwxgUlTOBUwY/KODFFNmNT+ay6mFJ3NG0KVjLCGk2INEM5
JoAdPhBRvia/19Kh6StG3ZniVV003bJH4E6b9Wtb2xXx2umFAxDP0DyZOSrubLAS
sne6VdTwY5rB9HEsWvNQAdV1N3HR8h3jc4e88EUwoKeRTObjfDuRYcImzAUl/FzU
tmEbTFc/bx9a+nVO6Fql4Rp66bdSbSuw6LoxHl5LarY66UMqoGW63+obbCV2nXH6
Ym3Imh3QtvN21Z4d4Ss7KgFgj6OxBGqT8gI9IbjV9H6eM1da7K8Vh6ESeGd2ZinD
FGnKAvSA5LcTaiACXmalQttJ4epES0XM1wP8vuUuH8A2B23gAPOW+im2vwN9elyC
AaGOwYDcXBlFKP2/1v+XBBEv7uyttjvkMxURhO25GFxhmbfS1vjtz3afqpPiYMZd
yZAPhobvyT2bImy1mPWPvc4vcPAnmm+V3zpbcThVjB6diBwJuw7+MdPy/PZkylhe
JxaNfu+LotHssRLhzqID/RLXurYRRpxzXSUotEcjSh0y7WYzUjdH5tTlmzzOEI0R
optN09m3fPu9y/DZiUS5N22oTPJaAnRc0E7HJO6H/c5Q0/bS4Z7OOuJfnuNwJfDW
FtGl796i4lDj3lCTQPEMKvs8zu4ElbfgqWziJgMxzfyvKIxZVt/5rW1mfuGEydrY
yupm6BNP2dLJ+oIcrC4AxPAWZB8LJhIO70pbhd8zYsefiUeXysNZf4cltFFqohBV
9DHtTnjUGOTR/J1qiDcJ/QqRAf1O/AD5MFp/nNlTyUFinmpvXc+MsyOoMx8CYmkP
2HlvGagCIIlujKBChaWR9jZijN3rEJCTfOSgAPHCMkfRjkGiYfLxU6Q22+MVbzh/
GWtALJjr5M55rmi4By8Ap99cFUOy0noAVFYsXLYmyiNe4Rais3aMjRGQjha8kwIz
MRiUpDlSxHaN08EcR31raxMgrkNTe6LehXYmLCRanBOQCw6nHjO0EiZtVPL+G5ru
jV+ZJCF/iEx8MbcxqIShQvi2A4WfVHfkrY8HyL13eA2EPzvQQJfp5SiR1MCzilU6
GhI29RCiQNPyBavHX3ZflvsqIus6l/BWlxO3SYwFJsChHI3wk4853cu8+0X4q8xm
8UETWHYUUR8BpWMNExq9sUHaax5ikK7HNUs3Hx7a6/ideUpayolMefwOjcxie5Fh
kg+XgWzjLeLMoRACIlV/0xTOttvJB7kGmH2faEqN701WYHJF7/hfZiwc44jtPB93
3h7dkGtm8jP3Ui7Wt7gaMnk8jYLseEWFwDkZeYrncaJnEngTXMIIG6rVjaAWUrjT
oTNzypksKQDTluSqNpt3hSQiE68APoIfDoXq5QjkTPK+aSSlERTh3oQHxvNtDeya
7yTqQCOFmZklKfvcfsCyzzwShMgloejrbHRInqnYRMg1gUDrjHv3wB4Hj9IF0iun
e1BAbNa+S0GPxixIenUOKqWwe5RH+h0fkj814HvkEHqyzOw6mpIrE08sJFvlQrqg
2H5fWRQSs4GkUsE3Vbxh2vWN5gokj9d38yuY+kntrq32sJfR5j+nZYzBp1o18rlp
XB+z/ImkWUa7HLtBZlokjcBjVsvPJgXXpMHsQENLBonrGYeU6SRCY+8AGHaCdlOG
1acfaIHNeJfvWIRCJ8KRTgngzXcV7JdcIfz9/UuqoHhmKAURy/v9Iu82e0cWzYaQ
hs/cu3/6ZL4B9V4nYoRx0ibFMtNdtJRtTMLymf50xZU6hsh1Tczn+ynmBnURw1GZ
t0FdnGgRVbp8o7DITwZjsSYtRvN+Ij9tUlPN2jh6vVDjBAcyYGSEFvoffo3f099g
/yjDlyCQXaxAXzUPxfIHUC2BDtzEsoKx2lfS1Ag0pGjPIFSZjOHiVkVw+poBSqZn
6SckEaHdP270eCevHE95yoVdY0M082g5m1LmJ4Cbdv8LjVHKMZVHNC/4KHP6z1od
RB6bKRt2JHS1fDv3jETAhCPhRnqeKQBkkcxKK9kU5hEDHR3fpzQAaHil0tquibf+
9phd3HNlIaSxsWZdQtlcXqShw6bGobbcb+iIxRBmBegbUZh6xNJBOSa9Dc5mDLyc
ziZl/nDq27SOzuPPzJheTbxunBl2gvlc5aoGpledbgzSRNh90guLZvyIYz7tnaJa
L0wEHge6Glc/+Rlk3/mbxQpZA/RHr9saIQFwBntQfjJikCsCpIQAO1GOsONK5HA3
5HMYHV9OjrATw02M/U3R0te4AVlLU4iFmk3JqplQyrMzj6xyTtXImlvENifv4hJC
V6Cie/1V0oG+nd81Skhi3DNjOU3OHS04yZjSHvyUjNF7TCVX5wBgyIbMpcEjcQik
ctzvZAJ9lhDheGFFD5VU2JktxRzN+Rn/pZ3eR+Ag8XgFwHye134hkuEd7CfDknxT
950zvvlfJB7W8r7xzbctOUWSjUrVdLEVd+LmrEMZkyw4wfFVOneCPti3zMRVOo89
3GlrQXkVrIAkdn6DP0cOR9XQ6uw73NUA/CDWSh+//ZWFQyTU2w0l61bh3F09c+iu
huCtEDa5Hv96bh5oe7ltnipSDOUTVPxHvfi+ciC0e5FuZFoESxDJmTn501XOwSFk
aeDTEjuGDmpSS26KJYsUjbiBScZJ8Sq4/xwBqKb6npU62VHCRhDYelaMJEY+IfXN
FGvpUEwaB4eGvHWpEcKZiVizgJI5a/EPs+BBEIrUTZ6P4qWZOQFGI47cgFg2bAgd
v+NrRPh7kvDPklx5qLlaky5dwCTXMvI33VGwGmwAA53jjkesHnYeAtyuksx6t2OM
fDsKFR6N2bM5+xLmbd4memu3FyU73xVd585gjjsr/i5jMF6zPRI5nuexJZrQbpDB
NrKkf2wlsxGGuClIn8OeDFg4cRt5UVFG0AlSt9zM3JLHuC+D3kekT/dt1Npka4Ot
oniC/GZwfR36X/49mSwqQZU0jRJFQqz5631M75/rA5AvAZ7uAF1Gx1AxDjaUvbW5
M50D2k8H0i62YTb/H/ZyBbxGSeQNpedHfyPUq8gvDr0SvwCmior4g0mJ3cgcXMie
CYdMM9VzcU6pR3PTmYU4NtYgpmhTjevTqM+Ap5CF45eJwSEVFmq8TC+O4i+kbPMw
Wu6qBLGD+EHRk+7VUR0rhjuNwHcecpQK/BWfYJi0Iv0xz0spC/QlDVyMog2FiCMp
4DP2HFnmQQKpD5fYdH8UC5uUWSeIHgNBhUYBpQN3g/gQ4hJjzIYuQDz66quk+mkD
hDd8W6xeTCaaaLxrpbNUpuCUDFnF8v+lpMybYuYZFDGXIryg0Q24hA4AZIjgjbSO
x9fgx3L1MQaDyzKTVeB96LAVaJC71GD/QG3voWzdTtqXxBY0QCdCQis8FgNe2BTV
KkyLdxR4qI0YmkHVRbN3v3ailUuzKQQ+nEy0Ly2ALiEeR09lBUqZb2DZd86mFD2E
Akv1+CkTR7CRpxBg+uOO+1I+TydyT3Xr1WnHbufQRWgzkRUmmEpsHhU5TYFTiKbq
14cmoMxh2YTwP7fN4eZL3pQWCcmGBrOuEqBs+ImC6z1SBe4HmkeJO/AihUkueZLn
xQUu13a8Zcd46DDhC02HOYbwi+KlRGgT55wKH2h+LY3m8UoxYulkyLlAxDjosN4O
y2arACyYiGfKGVmv3msNLZxu6XrGRU9uVM7wNn4HsxTXE0NNHoggrhmj38/oVIjr
IpFxKgKsw1he6mf5yBz/Lx7VUfvoTNl16MHeCDdW0wgwZ0RlJN5qwW8EJfUmc4aa
lyPqqDhcmqkkvBMU824JLQg2ZhsyW82vPvQ6HRRIw9MW5mVecB8ae9/AOzb2KVln
m3F+StLFzPZHEOYWGZb6XgXe4W2Pl3OefopwLjCHmou0Fa0tBego7Pi4gzBd25jg
uFoI3UdE2WU9D7xLqJ3ZKdXXYVuGsezRmpaJrpLmxD4Ix++p48oVjI8q+26rv7Fj
CT74I0HC8lIiukLwOlpNyVSwLMG8Mg1aqGd4YWodorBSakzIpY38LtWLZ9nOENFo
b0+F9LBRzav+B23xzT4T87eMQJH2Y9ePAEwVpO6fYq/E7fxA5L0ur3mexRmAQkkp
zKHnbRClbM2S2x+CX99zmEElsXJJDLaF8wHP2RCHOYw88JQabrBFMrHoJCx2fP92
Ty4vaiIOj78rWrdOGMvMRen450TBvcELmUJQpi5LLTwBmG8RZC/SyzidlQK1IebS
IgoAjSDGodlwbszPk/kaLbkVLIq4ro8oD6rGrbTH1o82soW+EawhiskQj3kLVTkw
ljlqfLqzHvhsRrNKccW+xY1jm1FX9x93q5psb912oAk9MeAvwbsF8vOfqyvqpfMN
VXNQ/OC6/1Ohwc67UTl4LUv5dOPL+PkAH/FB29oxvO+92j/KoZsjkHtbUiv1qt2e
gURfG5kM/yPaAKP4dOspJMKSx8eE/svEO7wDv6e0DC7omuYTCg0JIIizlpl+2TCM
AVSHUT7DpZFyWJU7QYCB75ujmuEJCns5EeAuGUe6Up6jm6kNgED4CEIVniNq+cZ9
3GTR66015bnX6klJLA6IBZ6cHX3TyX8i/C2ObqG8/YhMSEPYz+0t7kkk1LxagYvS
fcRupbeLFCNjCaFckaHx/jGt3zi6Dxj3+V1rowlhxvHat7PoL6JjltdoFh2dFxnl
uSpFy9dGdHo6Vzqi2nWL06ZVtUf/X/79bBwXjJxrDhVb0ZdaWHmSh88+86gEIy4s
GQwU4LKJGETnlQW+p0Kv4L7UPKkzB1ZX30nBREaH7YyD9emxmhhhsZLuLfBrPJ6g
bpH5wnUzYnlU07Y82TRYdGfVFXAQFDlz1IQAMVTl6M7qSx1KlOJhzvryMV5sMtRq
yBtM2UlvBj1yROv+cUcGH7NvnPNAQPxiQmUjja9eU3Vni8fMpUBSPLTO+8sttGx+
ou5D5+2ji/VsRjfqLYabMae0j8MtKZloimZCkWuLjxGeTbHH0R4TMCY4ixbR05bq
RICl3bTvi8ymaGNGel28CNZzHLdvdb4O4VeeH6SGQto0qN4PSJR2INlwSAwPbeJp
Z3PZmuliJ2PBvGUOcsofWAf4OL0gSaSnZ1VdpIEXmzU69uPxq9DYqrgZF04in7br
AusdAL1FWiIMj+E4S8xCCFa6BRGF4Qr4jINT1FPBNQ7dAAnM3Xi/Xcmopuz7HbAD
wzdEBa0eu8QTPEyXgrA+9knJMl88XwbPv3ICi462fA26R2qbVZgUeyQ26ZvUodCw
BqVDtCGkyfavLf3CzeCLX+Roeu+2BioeWaieDVtkdX/wMGIddWTKqGFEsnLrikY8
HY0QU+9dWAevSr3s89JR+QjAckG5pd3OAdvzA8JWE5Z+RPss/D7Lu92v5vLa3vyB
rdvNT8BW++Pq71f4IHvE0jaimOCedt2HFCq0dRI1W2zLfhA1XFQZXKslBCzlyo8E
pnJOu2TXEXgPjlLEAOWJP4xUl62ZZNZEY/Z7Ry5n594tVz+ETKlfxHqEjD5j2TBR
6Z8dmI85cQipHXYYQmKgsu5GlG91033Hsr+UVyuFYKqLoPjpUWydG4Bq7w2zWkxy
4cvQbz9aS9ps9eMcxirgrLHi1L4dtjXASadlb0AJCSQ7vApFWAWPGtr6z9Jgv4cy
VUaVp0pTSP93XabIoEUypGlG0EaoFdqYN4CGozIi5mAtNDj5M+CF5XGArAw+kBhN
S3u8eYguht6C4P4pePm3U7uZg/d41bc+Cjh/8GtCEAbvwjeUmSmITwiqjITc3rRx
/JAwCBp7lHkfTNHvG6CFzmRT33iLT1RebaJgc0EQ1R5wU/uGhcSihkmYVyWoZJVU
JpB4Ci4LYoK8WpOma3wZRHNBSINbmBXiKX7P4bBdMN+bEthQSwAImQu2w6zwi/qI
1bhyLlZyMuF96AfXbMTLwkCHUWqbIu9En7oz6QSxC1zxiXTKHjD0wMvgZ4tZC6h2
bvWJbkM4F/XFyMrQBDRLEwm6b38puJJzMbqT7LJM8gfjYG87st0WO+mW1ysiyXSf
1ZFAuj04r5g3BDyKegZuegJ3kGorjvYrC6oKosPwJJ6MPjAsVApCNSauLX2VG4kg
WyH2WV3hAh6nEF0T2uToLGGSXHWIqMRMxVSiEv6YCMKGENl0ihTlJ3jYdVGRTD+Y
p2k15qsqNqnNA4YbnikVVep351O7rcVVeEBXVwPoL2BZzO7lM6C96edfxa09EwHP
yDBw+lni5gt4xaeklklTM3jInYX6XAqPNin0eNTINejlqp1MmumjAI3eV+s7HhW7
ZL2nNf+oqyYD1uFEe6fzQxzlDCXEPNchDB+ZFFS4ePDq2QG7pRWMzMa8wDxo359t
M+ur4/1Ud24921846NVyXm8fd9/unnadAHw1r8VpPkm/dBnm1/NDHxmLT0rPSjed
Pn2c8Suis8meeOgUbGkrgu4jur4sWdmOiD3ttY7TIs4nQ2bLi9zkG2Ga48PewD2Y
Wi1UdCdZiy62AT4uAFZ6Id65z+DHRmNHXl2P/VUyqUKalN6Df8HktamJNyWer6xR
4mR+kv3nUvKPfNMWcyNoI4LoOA0VRMYzqEL7uYLFf+BXB/iSgyiO+yqL5db12+av
VxvrWfXFwXYGoabXIHkR+60ImRlyI6+4+MJ2otlA2ybXLjVg+iE4F236vG/dErJX
qJsilDjZVcGV2qcI4IoCZM09Wz0Nfb615/U16FhQ52qHLlWnCZJ/ngwd/N4Vou1k
g9NYlrnj2HYwrM1LjnDleqjQq6Bzfqp4Qa75f805zaKVGLd0FbM8nu/JJE0Rk2jS
bJ17baitwFQEvxp4p0/canScxrLERqXT1rxJolYh/BH5A68UAzVeE5B7PLAjPApU
QVxW8HddlRkw4sHwqhKrobkrGvweepeXa8/LNzsIPcDkzae/NYYKOcSDfBUh6kLw
ZRu9w2XCpMGMr5VjJJ/Bu94SxY+0uiCLqFSzTVc11xz0gM8Ra4GVpfsrr12XHO7c
5BejksSvv5LX/UePrg76ArZEY3nXaWp2Iii6W7hIHs52j+BxOX4u9V+3Llwyho2T
0xKsa7L1hg2AP4BjVkOmCX2AgJwDIZE8ik4YBN1SP3HcbtJyMKmDmm+y8crTA/3G
8UlmrSwTpbwLJrhSNaTEHIgw9ul35HmCvCdY0NaWvZORGDf3up8L2Mu4TjK0VqBL
b8Qxh7htV/hqsshqBOxkOzN01Z5Ojun2kvCsgVm9yKzhKAUHPQXUsZdARAKD4qD2
CghPNS63K57YhImd+jtFDuoFK+WwypTTx4+XxBfeTA3jpqYnrXMav+cYqwJP1RQ5
glbFjerF6wlNoMQQrzZMkuRWrq1V73jwB/sUxsgZ9DPByHYS+rrxwO3KUlzsW28t
umokNPhHswT2hrNpIA68MGUvEe7Q2hgg8rYOPyfp0HDHCtSniApitrTViHxr2cor
oWIO4Lmi+6j7eIyl3tNzlOf/uGHSa1XHQpRBHGMgqND+nAm/Xe3cZKo8b2bVFZbL
JEcCUAhDDKS+6nfRcTpoY11fkbmB8EyBsue3HFW3ElMOutzY8YahnN+QpZYe3ihK
ehkXunP+3v49Vnheq962ANHfd556dAXmQJwuXMGKd6q1ePJAzpuxy8Y+Ju2vEc/n
FlEmgpvrkJHPP+hnwOnQW4SS6BkfqpGeVJWjgc5nz6KdD+CxPL/NvM3guVirzvXS
dh7J8yjZLrbfx+PwIZ2wa9jC7XwyRmbudf9Qs9Cdh8yxERoeLKs0y53Ze8tBiJ7e
2s1gDEWqtGJDxSdIUxe2uMmW/b/fCTtxDuQpoYCzVea21dMwVPuJK/VU3pVa+Q1a
AIoyiwKleEgbnDAEKfc9zP2FnOaGmEg124nnEOKtwQAxDXSpWFderBrFbpjeCk35
W+1aJBNkDYvlEO7oEAvqAPffQpsyKcwAgmXhTAU11TqG5OJOdj/agKkAfGjjff3O
cEmcmVQ2+l+vMDOQqQ3ScF0F8BgTRcRVI5bzvq/q7zCtLBXqOe3hOzGvwSfaTJUY
PC44LMYHgZNXCFOVb3WgxSyWmyH+AolKDpUhmSURU36R1vkG2nYlfKZ03WkMlvHn
RPmrWJAa03inFHhVEWC6fh13TbBsEB/ok+yd9Ifai7J8H4vxgQKHCR28wU1kOwZ5
zkPpFtwCaP50O71yk5HsDKu5n+PBloo2nYLbVrvUNHQEAJ5+Tsu3IpSLQZ7nS7F+
Ejzj/iJkOit25ZqGqEicxGd0PeDJryteJnyOP2iTyBCpzE4Yb1efCYj8ZOoJul3u
ghW9h6c4DJf8rHGmqh2ORXT6T/LP59qA9xrdjgovpwC3ocqlw0FlqHGCMOiJiKH9
ATIFK6dOdIEL2BZRyNKpT9EIoqCmS9/ulvPtsbKLROi2Cokboecj+1EV29Zi2phC
boqT4a90p1M3EuahCfaYoQLD/79lRJEPLRsTYgCslYlmauR/igVei/VqPOOb2FVL
pWGniWkRNuInI4vh6xzIKt3UYoaYuHTi43GcPIT0lNSapEzfrdtO6oFWborce3C1
dtcHgVbphdhm95LULFv5pfyFIz3eGVf0ncIOfJoFLUq7ydzEL+uYO/AkdrVkMc7C
+Rs/N3ZliCpjZgJns/2AR1Pb0A2HusS4TblnOdZUXSfGO7UGYEMa5ViJBW5kdVTs
Yx6eyEefuGWf8vf/vHCAiqSujEnb6uJQ+YCEuxtfr670OGYpbQJUO7e7+QZFISLk
J7KRYsTELirp1iIhCKSunpJWssxc6qVLwg8n5wKpZ8nuf2Wo5CDOpzfaj/WXVIVq
znhTDATy1jYuoIm8B3bqO/2eM1ONO6xnwXNhxiVt5HZ6UQqMsgvWSgdYll7FIkSj
cj+Tw8md+KQVpFBle2ryGuFcD8MmNTCUc2gnRHUn2uWySbInZa2VeAmRHbN0H0WO
Ki4ju6Xm9mX48NzSEV3mS7mZawtgEr4EFepJAuMJZ0rP1Lfw3/hdbyohUv9PPbFD
B2zR1/NUMV/9V4lL5/pO4eEqIN1Rnl3YXDUc7ap3YWyEmTHVS4AEnBsQPGP0oM4U
ekqj7x/Ff8Xdwzx/UDeIik6kKz1lweVcl5zdqKd8yjAr3Rxjr1QUn9p14PxsfzpD
k+2pz4cnop/4Mv4jBjdeW2f8rHkY4PN/YPlsVyovDaoOxLjNrIG7eoOfHbQEUVMX
j4vm9ICn79FPLp9AsuH5DMI8/QbLEkamyryzpqNG9iE+LANlFINKU6rZNsvPA8yF
ycjxUsk83tHLaKfmrX6jZZv3H+HmvCPeLXkLFHIK17eLegPruVL494DSbEtmWgJ+
euN8mMBkO4gm0CXR3pnABTFV1MdRGdAY/WyWDawUSIDYRIPN7FKw3coY88mk4JMW
RHIMorr1s4x6MXXjlg1jiNaIFRywmGNhHR+9GI2Tvj7iX3IbU6d4L5tBhUfVyeKM
+wIlM4GBPeKTEnUkW9HhAucqvp/2lxmkv2ddILjbD63XLkDotksL3Ienr15vfhqd
Y4u9ehHd+ygcSHbOikSb8WiPtRavPOw7oW04M2Rv0s0uDRx2Rfiaq0PGvOLxcoIj
F1KOJP58ZchYF2/FbJt9CAMHcL+OUCtAp5vsRZnWFdEajLS3/WXObeVYuNOO7J3D
AIpBLFFuGGvLceewn3KyqZffkC6sleBEu/RnpYblkTQtMgMwmoYMEb1tTVf6Amtz
IoHBywUb3nKT6PrFb86CxTUohdKM1wovhB2+hO+UOpdjq3ORbzB4vNUPk/zl81LB
+wUHkhomckd4wZI2z1vp1JgtQnLl2I7Rx8+V75ekW+aQzlcPqeXCRLzQFwpPYGci
ZSZXhKd8GKV0hDPmdRTh7/mF4/G38VpHRM9p5yeqKRdsvuwEYxWFNpPsFXVcW8K5
q+kQ1VFGj6OOP1o3jP8rX13xGWQ2nW1jfe7W1LBF0DS1RL80Z50E4wQmWihMEF6E
qpXAvKUSRSlbUrdc7LJcMxIowGgtbj8GnktSNZvKzAISrz/HUEYY+oWldOpiRkET
9IGQrGCUHFr8EB66GfhytpA5gvy+MjbiCq9mhNeQa72/6mv5AN9l+PmzzayLilSN
ns8jv/p3SMBwcaet9TIYnCfheAoAcfnp/1N5Pr500sgEJDBEAxLVZYmFmhuMfU8L
Y/gUAUzVYvD0l2/lp5OLraLfxRzqTvQhHVanIKSAJY1VIqzuhIwvoybsdlgMR0XC
EnwJDIbH1psl0eCtWTXk/j6n6ssFD4QCPJAwUQPgK1o3flCnUDQ12uCtToJjpRAK
yw/vK1xxdFWwWvHDFlr1+ujSwwXlzU431pGk79K+zOE/MPkV3WwaLlTE2CWoWfLT
M74yxY8bc6dj+43WR/abNlqEBQmpvBlUrbxAe+kF7dQpp9YpgN0D/CPyksacHjn5
mMZweZWA3gOCvzno8+KVjxIEH+Kf5zBQrjsJTZaJrZkoeRKMTCV55ckYjvM4b1hS
SX425go+9Kj/oDRh1oe26B96AkNLFeJeuJ6EjNPb+Jac7bRESqgimpnAQmDydTJ5
Ph1I5HKg+Pcq1GZfo7nnfb4jPlgOx7YPfwlgAARqBduK6iHVLPyBUbha6qPTlXoi
/j8n+QzBFCULi65gSBmRscQZFm0rsdNzyOe3dNX5kGVbvqWM0fbz9hiKqyI76MRN
YIbF3am3EGXYO7t6hvfqedMeWH/z88B/wrf7H2ixHjhklHzkeB0I8U3nB6r8ebru
QTuz3D+WFo383IzNV+F5MjfH+sbOfVIDV9oHMwpuw2vBUGjXXxyCoaX8qUtpW0bt
2juRFKCn72IcfYjorOdmrLRBlE0AYyqpgeqU/9Aor+NCzPAkYZFaUCIiZX4iQvtC
GbJdHwBGEyduILRZ+HNFD6eDq25flvznpD0JIz1nV0ijdIPmJ+sXZtxJnw60O6Fy
zkGOexwc9u0IaABIddwuV/cyjWGrzkU89ewF+5H65qxuohLkY386xxtZl4ebfX1y
97RBxKOLhm2HM0I2J/b6Bb8DBrNFoKjU8MnwxaAux+e+cBFi1byfkSEAuviqkpSt
CSH5hg2gc1xMfO71IUYH9Z3+3VhBNovsqDlDV5hJ12jE43ioP4ZgSnu0BVHmvWz/
4iX5knZJ8PepLV5r4QkKdRIkBc4EMYtGfrqy8wlm+Ytk3fLXpkA/9JaS4Fbl94O0
kDVnVN8TZoa0Kz3E8JGT/XCBJUXYuxrienbsPP25v+tnmr3NnYadB1jykrBa2UBs
H+uvQl4XoZKTfnSEbBpP82haWwamNpwQI0YEB9jkd0LVjIJrQek4oBU/QYAoTamc
1JQrd3xfsihatbYt7AvDyyWiu965Nh3gydqIgoxwL9XaYnXF3rlmBq3QI2750cFa
/+kp8ZTpTKhvQlw4UDwFRyiZpuSfKGx8YBTtDQSGzh521sRPSsn3KBz7js+J3QOa
NssY4yyrRxvLi3yaR4bxTRhLQA9msYjFSrj2n+XBiN6htyC1ga5CSnSkd+eEZFeE
lJOIzk/teoLl41KDCqRp5FjsjkJeF9s+SJ+50y4fW90/UEVFfPDlX/LoyRlq4q+1
OdExtqyudgCGem9+/n23qYsj+uGcuRo4ftNtFNB+eMk3tmZfaTo0yV0gb7wrMl7j
UuI2okqDIImC6FGc54q0LqSJDzs9BuliopRFKIUADJf7RR3+7KH8N8HZzrCyemqk
gOHmgsBv+D8tUlBaqzuR9I5z9Z+ojnuM3Ie6vvDVcX38MOVo8u6cedjy39ktiBFX
8hu1A6MVlfiGW53m3XP7EGxD54jeCi4brp2GFuKWmG0kXbiSnj+fffviA+/7aJW4
8dpcu3FJ7HDxniX4ZlJJIjpaMYGa62T0cKpRHoXKuvIIEFEhb93iSQFPipSRLOSr
BK9lSHQDd1XEKeOxOZflVx4XfeV351WAdV6tytbMhPiyYmR7uKn2B3zGVRX/xfJR
xcEspeUUjo+lWYHaZOBsWEpitU8Bkjmlz/RZw1TvBo95zWAm6q0HO/n75UFjqLgi
yxhFwJrAZqbHHJCVQVvJhY+VixpNVRZbKucTmv4sGKz7/Admo6HtXwNrlaHz3Qke
d0fEu1bPmaZxNbTKrWzs4FJP+NlKC7LEw16TjP/cHups3+ZzahNJevmH39FupN5/
CP3lH78YN+4GEICm3vQLdzSOgxxf+m3g8x6hJKbiDqTVJlI43jo8AGYcht8kXeKe
7OXRzyR63SgJl3x8quQv4ZbOEOmArQbxizbWU4pR9bs8kKCcTM3gjq2p5PkN5ZtJ
hudtkz9ngMkIBn6DooSbi8L8MLIbikH6UOIlJqtWsvuuo6XiAuPDbQnQJbc+oAiQ
lNznrDgCohdU6VmLnyWd9+Il5ae/wwgHSzyXqAftHqC37GaBAaYA/G56DDaX3bcy
dSTjECmWEQKOXwquk3gNK0vldbQirqOdnDCq8y1F98WjLCl/Eg2GiqYlnRfMEL2O
0EzfaxHzcDAgazjE1u35aFjEIxwcBICU9PnNU6SYI2QDfIU6446mxa/9/FVXUjfv
2PtcHt9X1TfJnPiNXG5w/oy27LYTKUlId4KYuJT9N7Kx3kD90q9Ga5OtIAfbUwDZ
64iH8yoMnLByHzS7xZIraGv49t3y9jIz1FiT41RP0vcGamw+rv5upncR3xAFswn2
5/ETuFtVA7iAwFWZoNgVx8HH3bjNHSPh7nfabStJd3ZU0+3V5P6Z8XUBQzPArOV1
48Tqpcr+FgalYi9JyRXAJpnWHSlbsVZNQCo+yxvAMb5iL7zCN8mqAw5k+OL+sjST
tw4pKL7v4/FHIEF8ZmDZcuYWJIa9CB+p4cZ5rbMsrUy27k0uxtJ8b0kuq07mOZX5
kSpsO+Zmo9Fwn6XyD9C95S61xpN1RhFyS0k6bgRhoNXi2/cICXCRdmUG6JOZrjfR
JfJ/lx6r6ZquKUWCfaBw+r5ImMxJUh5o/q0xAfw9OWf46bfrQjzRhMYktNf6QuoN
Jle53iMdmOMfIbo7r4feefYJbexO/b1PAkWO5L4jEvM7BaNe8rai/icVD2rDZ311
ywX5POPUFyd+0n7nkSPC4CdzL1Zh7+OrviI0s53AFUtTdohmGr1XvKMzTAtpudbR
HkpbQ2hsmc/kTagFSi5iAhlHq429fg/l2Qh2/PaDJbrM+sFJ7qi2em2yzU5+Tn3X
F3JglartP4Q0lRbsP+q5vxVrnee3sctdBdMlY0AdCetyR+tEXCWkdJB6YshFVb/G
Fuq1dISZRKpX7uMiYS1k6qg8TnbD5Flg3nyforC06ZJEcfCJdRpttUgHzMUw6I+q
1eL91z18SaUJFmfkFQCaePgZByuE8AL2x7wHILHMVtMEtpg4/wkGeXvq94fqLVVK
yy6mz2Skrwr5pfHn8wyCQTyh+6p43/Mq+Gc34pn7ZTJPgjJr6skdpeXFGDABrSzJ
PB/1nayWeOOuFH+9ZQ4M1txT2hklWF6g9gkc6Ghz/s/UW0laJsc6WLItRdl3oy/o
aHAKP1yGkAIzm8zhnmYTeiRTisvRANVv2F20U4P3sR1l+ewlA/NvgsH1T2O/OyEr
zfv/U5HPOdnjZ3gQrAHWTrNofgFbixLV0mUEDv9BuUWNiIdDrtC86mthdANgtn6o
22/7bG/hykjuxKwxli8L+zVDiWU64qkfmXUT14bZv9lrpK2cKYCaAt3euBKWTAse
9TBVrfcRxVUlPq7FcHR53MuCGNWEOyP2lNRQ8JxT7L32CDALQuOsGfqfp5UORK+L
6yBIehj7BEQtA71jtPhOe9ck/1ErQONRQ0CsGkp5IkRVY/xsQ6a/aLA8iFHkIO9t
/qTWHx3OebQHF6m22N//8kOdYIjmDJCXoNxOMfChO8bv7OkVM0smKo4U7Q7t+Ah2
3P28KUoRnwfVs5Arv9KYKaE4bKPpRby6OFdcVMQnDsKIqcHpDKVjVGTQyqVZ3NlT
WebDkoU+MidEUk9QG+pcOoAvzvCe8yI3PTv7SCPoIbLBUrx6mn1GGRzBgPqEC6qg
S5wQKsvp0Vtl3vhQZJPPyzMp8bcpOjmHKlpkzRCcEYk9EzboXhc4VM+sICGOVLQX
YVIEkE3uE5G2KE4wfgou7yFsKjEEe1Ki9B/DzerlttzV244x/xxrLY7n3/nEybsm
SSTrtsYPpcIy1LQmvjlH9sfk4P6jxGQqYQmbgLJzOUYH4SzVfgH5AV73hrTDF6DO
xjjPSq/Rq/jAmTHZTui3ecQRiZk/j3QNyTKJZ1UEqaEtaCIXUneYUNKC927wNjJC
vY6faUa1SEUNGsicMPRy4SMHwF1kQ/fsYJ8eXlK1ekBeCp2mabInifjrLN4kgYGa
zggIqV7W4li96CSpz6lJl2vKinlxuQlvC6PcvQzjajZRPolFue+uOuSSBKN20GWj
eKb8wvsHd2M+EuYx4MR2zIXCEJQ2LwfikMGgNqaYklivOh5tJWj4OZCQY+iZnUMf
4aUwFTvImpfj/g3VYuMpAy9v2h+XN5/l4AxTtm80yXI6kvyLxudmUBul4lzQ4WhW
bnoqLV2fSmSRjZCRGX6/C9upnddv/xUJtB9cqdLqb8NOf0I0BfMWnKYvi5M3KKWV
yEGA+DxCqmJH0PFFeVpNd+Mmd9SgpBNjSd3jW2SGTLc0U1rTi+FD49odTu5/ZnP9
SlgIQ7uJ6yuD21CoLuY9u4OXS0Y40L5y/mXAKVgR2zbCxUQdMn8KX0PEMMsl2htm
eHTmVJR1hMqdD6Ox9vBuDH9qGkwexAIUmFe44oMnzybHI3bE37KGYz5N4QPFD5g2
MBpEQQ9T6LUAqsV71ZxaXYg1qn1QzKQvy14DH9w9igYZkDWTeh1yLpvN6MGuSWfm
crExuNzBBrpIuFsJTDHd6hROJjQzTVfgdu7y24eof+IM9HWxkTTbUzc/22dipSmw
kWCEwWAHdVNw3Oddr296uGHnhc6offL5ggnCHryuNsB2+Yayn3yxKBP7mkX3RII1
ZO9iNcDs+MKrd3Xmqps9ZFCEaB+gTL5mjplwLixf5ChOKL2g+DOt56YllCuqpTEL
TIGpJ4QslyFzJMC7DJ/H7t4BXkxWs88ArIn9puy7sCItWKzUIwnWz9UezwQsUoOV
x3NDhYLcNPlss/5RxdG9RkS1cwJwQJ092loSodGVw+hYjF6EHZT1XxWHU0K8QncS
W06PkVMgvJnJE4CbbwRazUNJ0c9pMU7rzLDjGcORmVpEFUBD5TM0T1Ed8Vjnjz/2
x3mvLRhivSSxue+jLl8MJZxErUlFWn2Nqiv3wpFBv1ysWReP1UDtqmfye3wHuKRN
PVnMaYIpMVcwCvshHGFBToG3Lhzk7FW1rCBIkbuXV+Gg313fOHa9X0L1CHBySQGV
t655snHGjQD/I0WdYv2uqnmgKPwhCQ6NBVALUQX5DGfksxHfjkY7pTmmuVIfW4oJ
KQVQQyRMsYEbstXCUjzmO7qLEyi/FaSkjYhuToEXG7B0QqUgQQFt7xjK2vsjHAPb
kVo9JahgmhIMNk4Cq86pVfqnlXbb/BMKA5lfl9HkC33K5Ux9K9aMD7D+4MfepGMP
nFmg+anFnRneG3kwVJeRo8yx9aDkTVShKu2ctO9YkAghoEnsXT0zA+vn/hQvNbkj
JokPEUQj9pZ74cc5VB+K6nCf2LHwlSCPoQsD79rEjkHpVhE9MUBHpcZtiULfQ4Ep
VMEErip8tjAF6vPalh84DMqyb6M/LwytZF4OouLoHkXq9KrnEY03krDqiKfKOwhv
ncF2OSUWgn+kWn1rnZlE0BpS1iFfhcARxeTME3Aix4kfxbkbunRAO0Jwku1tgsJo
bGmumXPIUnt8/BKPOu1ZxT5OWMxbW5h/QZIHhZtN6JlK29bwRmMCWQSZkmH8nU8y
C5In4ypxrtRDVMFuBwWMhkphNkDvozMHdq6la5S8JCEUA58gn88ck4WUKOkGvOLX
3rjE02o+is2GCR1BocQYFW6//kJNcoc8BBHNwJtNJriweXCqgJKvM7QK/TlYTBG4
7WuSrJlyyUXXFs5np/UhZYNQWH0HN5dxpZo/7cLLxUYqW7uxbO0y3Ic+NjmMJwA2
XX2O1Ui5r3fsGChHsBRp7y0GCI5yR+XqiJv31bst7gFSpUIdmnxPU0Yn5MXLiUji
2FOej8r19+CbbWWQYrgwbMP63ZP2uABV7cYilAhNZY8pQr/Qm+1++oVGjTjERbk6
JTE+kNYl52A+FeHp6h0vIOpa6Bi97+i8ihscO8EWhJ5C77EBN4kRjj2normJX53s
nEGOVH2ehl7DXNfwMptDpsAYWHD1cOK5Hzxd3zHYpTGGZIfrix6Wyc/lLRTa3ciS
OHpQit69Rzm3ihz5/1ZqCI2nSz51yvuow7Gehx19LjJtxznXvXezRsVHa71bF2J2
ZHMjWv6fZDRAdCuyJmOK5+NUt4MPaltsaLhjYLJO4t0Imapsraqdvx5GzJtPJMJx
H8gJh9vBcL++oWk0pYYLdH6RBXxWUpIuqPqzUN5oyOy6NlO3GQYUyp7Qzg94kncu
xBxU62+tUY5YKNVV+1ECIqQsQyw18iqnHR1ltjdd7W6dsPZfRCGs8oQtoh9gqbsK
Q2kJzAjRopTv1l9gk0aDXvI7hnnrmH+i1VTqPwjq/xY+nJ/UzR1C8dKJQEz2eX4M
cl63yEF3Bl6EqPD+E+ZVQ2ID1xWG9OQVTwo/+kpmN9EkPBJxGwgAXgz1PAFRy/0h
wSUrjbzp7lTahq3Sswp/gXQGOyGhVJydpsQqLtTUd36oNDAg2UVjSfvrAJXF5/zR
FDVfgJdb6HTNZi0owQjWYZeP7FfKwR59J9FMqXiJZof+JS9J8ATVXyN3wR/OriwC
ljUW/e8snF46KeGzHiN68jtNJiI7rwnygAN5zmWo2GAZkd4ZNVJRzNVjwGW+Y8ED
oRCJGC9Ux5pUMPAHC2xlD5hUyitt+a1hnrTVB2as0Y5JfkpyzbLZ6S3NAm6B6HCL
On7FX/dvxz1H4pzbtlI6G7UpEB/oF/H5294DcEzRSo2eCjqtUZ7dkVub2dAw/TLj
OrJGwjTM3tCOv+g3IEAzLY1fZBQJRNomwYGz/Sg0roHcjyrLb4pMBI9YQ69IsqON
9Mys9Yze6tWRvEAK7jDjzr3MI8Mo/5PvdfMiHL6KTJZRRsfXvkJogXcrnEkDRbcK
B7xuS5WIWtIzHKCopspaPVE3rJOQI4RhQXnuFB5NDLh5RqkGwxFeK1k8xPjN7McA
EzyVgQGgODibPXFHxhCBKIAib55FLclx08qDfR2NyxwK5TzCO2CpdeLpklTzSWEO
JaJLgnr/YK8s0irXKudyUeJD642mKorjPa/txKpgX5r0q3X4ACVLgEptck20L2a2
NcQJ0/uDZxx8a7ZY/N0upLZIGTcepqqENOn708eZh3kzC3ahBVfoCIqcShPi3ZZ9
4eZqnOq9TYGEU0IJ9UFuH83REvDFaWeiCag1wH1IG/F2QlsGRToSfhlNzlBaXXqx
bvJO65BpOpgXr3C3z18IH6T37CZY/8e5T38losDSfQwLyVCnM9OPPyKAjrynRaYX
n2Ldeb0ncg5Ua36ZXG4SWvSDHc2DSFHU6RVE4eP2bwf8zbFF9MGonje8ohSdG1mf
1jmw7oDFwzbxrOcLOkhu9y7BgjwjiV7hvjG/SjtRpf4mAYI5PHKDZE/3fTm+YSlP
k9s4JuHF5DO7NM+GJ+QwzvoiXYqFLdICPEa05GX+DidhYfjMXdolmwV+/vlE9X8s
UGKvuPPavvyzLtN0AMlTcAj7bk/sOhKTZnCLv6/nJJL01bdSCLUyD6rELlxhmsUB
qlunQkjwy+k42uxqX4oxBuALmHNAiGD8TZOErOG+ld77rfgQgjAbGrIkTa+W/+Or
8TzXvycm5GwUz8xOB3NVWt/UQTPc847C9ZIjS8bozxRiv62QBwIB8t+SW/JiECZb
BpWFT9QQMVPCjeU3RjXUc3dg5QxPgTN85Kb+J1kevhuWWlo8VDmeak6/0YNQ9XbN
AoRMiTCkuvo6hJPdbEqFBxsnKDLVENi3Tb0kjrQNsmMZhWHhYuEZQC4iPjKVTjps
kpo1+IoJFSwxEipZiVQ09lxUPSxLsBnlJBfZEwijZcfLCmUYXBXS1ez+q/0etkkw
io6lFKRMOWy5BpfpjMGnJ1FCAdv2pV66bZwSSbtknQzeNz17XkDCqhVABiZkPTW1
yIR1I/PU9G4lA7sdETXFtPa7OMqxgaNS0UYgLDb0C3+AQY3/ufDxWbup5Q8DlwZ4
qqdH2nt4kjVRzauDesripYPC+0Need0Mn3Uw4+d/juRyOU+Q+E7eCa9U0AdhRpD+
rsovGHkKE3TqZMnesddt/WnI/QcVZTC2xdHHJMyptqI4HhsUgoCrVwWpCi9P1tRY
MkiaH4dklJnoQgO21blrBOj0flP9QvbJ6aAQ+wtGb3QbnIBEz3r2TPVcnSSkYyeE
lEuz28xiThERqBcRUCjzAQ23irmmAPsGRrCFPmSR3BaHPNlP3VEn5p+NKfEXAuA7
nZxfm2LWLBLenMQSmw5peDpjhgtChSzN7PPMlFdqrtRUhomq6lJwjUmpM11daGJ6
q0EZOW8lRXKUifEZRbE9tlluHv8MZhuvK5UYo4xzVKl3lUe0V+JCErG3mXns6l4j
e70RKZRM3uQhYdOSHz0Bv4JpBn23PbQLB8ytTyVCZrZHeXOuwiPZT8A/8V2NWHLF
QGV4Z//IV02wc8EZZ4CLZ12RBnMOliW/1A8ZGwXqTm/Md6cQhR7ChHX0wSP8vBdE
eifU5ijwxXrCyjjYh2B4FesYc3XgSxk1AYSR+lG/hizxh5uVAnzHl28UOA/GCVaL
+tNopcGDdrxAeyP/mlGMD/WiIPO/7aK49UgQAwT/nIO7PUvBTaBBomYy0MfSfq62
AcKBK3KkEjr2iDh4y3VOiZjVcsqCsZP6EuwQ71qhj9culcpeZFd9GKXL11dXDHdo
km12wgc8iy6BFFjMz/313fEK8XpFWo7iW7qsRKr/3E2tjzXSOkDg711advjhGLyc
nVlNRika54egNiwVGsQnPddHtxspfuPqNAxVAkRfa4zIRYX/25bNuoU9PoJ6TtJ5
cimAfjCk09ctJrpGGDfdnFGsd6YacEuufzgO3A4Bakl/ehJvzykAzNDRbcA0g90I
WN1Uvz+ySXjxfvyoYSJx9KfY078Ah3dE8pun+LgzWEF6tyLDCkQyL09ADSzm53Jf
hmlGv2nxasXvBYrBFedpKgRPs8rd9Pu/ADstPUIhWv/bclh5pBswixenm87ZiEmq
UPcRD6/ZDkOLQJhqgf4rpXDVAEKp5I/2EKkPwSDVHriL95I8znEwa3o1fgLJfxty
FlbFN1u7DY9YT7051Hgdo+rV2eQzYWzvrBhJGHk+hixRbsyfF311Ay1u0Pd679ed
c97//AfgJy9zm9M59Wrx/njRYlUZZISo8CYDVjcZu8zcDzDTrVdpGFoIIwdcZ7Qy
NnioP3Gr9qrHoeu20U1bOPPlP4LdfK0dv+fWNosi4dMqw3xxOOkVU9yLJ9JFzx74
y0bKIMoRt8Fr54xN0KRCbxPD73OlO9/L1fk4A9kRatAD8E3X5prexus+mvf98Bd3
B1DjzPdjyk1ZDmE61mmypqgCJiOWjtgLtuoGoceieoxE263DyHLtB3Z0Pa5vGytq
uKy2y1GEK3oDj3U1VbFfzY4ghVdaovJ2tbYLETZf9J0NwcvjLRYO3HNScEBlvoYd
VJsqLZkOHMejT2NrS0+YiUTZUiI1fF+3N3Y4tlx1jCnLWeCgyGNMeWgZBjVg25+B
Wo7/y8WUAGeOYL2rjynX88HLDlSIZigkQAg3BqVUm2VzV3T93L/xeGhsEB+7wBLe
/ntKOJ6G6Ml3M81hB/lDfVSwtqwpQJpGGqoUXn3zU2w4m061tSektqVED/VdL40T
3wMb+if9nQ7msPWe9uA2aW4rt+fNMFDK/bHXd13Axd2ZNuAu6EkLimP1472NSpZF
/3No9qNlloRxemqHVkw5okpgYjbvwa4UzTsauHZZyIlBgfI1/lA3VSoYvjueqW6X
ptkUWZ+9KI5gU9YM06ZWgSm4JO7QfJfURDDxA9Hj4oZMaZLhaeroQTYIs04SO3xa
wowj3tBfz23e7kRLc+MlFxQsHDYtcte3Cjz9w8ZCSJx5IcHLKlvavRIkLyshCsh4
fIdGIhINQ8iGXMw58M+2WB+34pJWog2gt99vIIjx87BnThgh6AIfQtHpSrtUBr9K
Am68/R3MLHLaK/TXseLwOrGEoGtFNXqhCB5bSUvf6dqXGZ040ZEYcWKb4Qg2Tslk
kPTA1jqk4dyDsgC8GTOKvQz2Ek0+UDDfkMlsKxS6MKyITFT8qh73A1XovyxDjDr1
P8ehJ7doSw+YDFZ/bqaaecK6n1FlWQzV0VBcx4PmBapOacFOOWhi/4VMJ2D8ki/Q
rEP+4FMQkdqjbgvlRwIK8/VbNFJCieqR9UATZboS4fDgdKLnVd43fxrAWJJS6CEQ
Jxbxdc1LVHzTXsR1/KwE60aZVwLbHwePm+a+6gWhl41o/Z8sCD6egCHpCVWJgUL+
6iMHn6SgzezDoAsf/KUS9UZJ1gyqovwb/9Cs9esZg6q+l3/ov5g/W+n/rxNpOoBk
ToBJokGKkEGz9SZZuzWc4qhbCM6DEzWOAamzDJr/yXOlRJo5u99i4sLeZoc/qJuB
iKEUMk7xqbPSHUp6Xjd03JHu/q/XPxVo+2ATKvWhkQN12otGHwJbCPDwacMVNqZg
NEVhxDmrgQSN0RuapRETSkt9U22OzVEo9SV0Yza+FL+V2XZ5oXg6QZLNwjTxjUS/
hcj+kfI7uAb6oa0+8fDRD4no443KpVpelPEac46X5RD2UGS+Q8B5jlCMg2SxO5v6
0r+dEbo/3sd7NtnBAG0wYQXEQyohir9Bm7JefJ0N6M2XHdrBZMtLocbzdxz3fqSS
mEtasDauJEbvM/5yVWZVjAYtF2ZRmYTqnYu3DyO9khYKujpsclrVFvCIcQUOFXrV
Tv4BhMe0U6x6mAs0Ak737awuR6SnzKUcP3/t0YW23edsH/f6Kusf6gIHJ7EH0dJ8
dYn/rGsP6ZYO9l+xaM+tedVV6LnZTT6c+a5berQwW6OyEi1vG/CjdTsCBqGNo0Rl
5sePGDObqIIOgOFpRvolhXMMeT3coX8jTQz0fcsqJN0MkmYMWk9vGMm2EOO7+RsS
xT34OzTcJweLx3s6i+MTvxqUKfvMxx+LHtJbU11yzoJQPMfcQ+g+x5tx9XITfOoZ
S74dIcgzLphDw3V4SSBwsY7+VsApJ5eDZeJJKGgNPB2dhNmRU5XLd6hUeKZYBhRO
jGSe4kZ1JDi+PE3kDj05o11oAqbwPMckr42OGJjuXkiT8HU4LoHQD25JKmWihNCx
rPOPWU/5T5LHJ6rfRS8FXZZL6ksNXXH4/FHa3ljhS9SdBdGUOp8H/E0tjk/trVpF
eZuRI/H5NPYIOqotuQn2AZVpty55sX0vMYDU+kU3RYP/9z+PdtUwcC+D4JZ9dyZQ
bYM72oPRs9CRT3kI0M38DTTcKjyB1nEMNx0PuLx5rkYVNNsjnWG6kfh/K9JIt7vk
BNOa3NVjDYndTspEpbJFIxz9H6NabEqUrau/YlaUyS0tMr60TNxYAU3ymGd1czYc
54Yax8ju9bDbGC7wvwjWDGUHa9VMlTWbh7vyNlpT2utiUYNrM7Zp0I+mpMAGZe8d
r0yVv1hPUjGemFkLuzuMYzeVIPPgYPU50le9UG1UzAwE6Om9jJ8X90yEKS0NQdOE
pF1B92e47oPWXHW2F/+IvMXf3qErGcYcDTDzY54Xq9uRlMcyEvwMinOvJ9OZrhup
eU91CT86/krk9lDErO1s4rFitvtCPN5EGrnLCFmYFToICjhoJnGeLQGzMSATpAoR
PN/pKsIGEQOEt3UJg2/7sLLHliDKM+LXd4NPZbfgz3D22pg0JuKA0CkfciCkRsPG
Fj3p6TuTHKFI/yNW7ErN16yCiOGct6Xu1KZQMbDWyRxhqXKUrS1vVhIb42aroIiw
XijEksyJQTCSox15qYPOHVF90nKjfc53danIjbkY2JyARSwwcpHgL/AJL20fn8vO
A86Qz5rVOV3R1AYNSkWOClNCvw1nFFuWHnm8cc0KvgGkLDiyIYhkB2vJjeqV9YtI
PBye9IXuNwN/WgUef0lJqKE+xcxBeK8uxlES8a+RpXL9HO/uk4rHdX5cbQF9+qrU
9AmmbfHAgQiwwx5RaPBle21EzS6hjcsJVsZj1A/WHVx976c3m0dqvTVEsSVekR34
aiEDQAmsvc4BvLGhFTYNuJ1YmtlHWbotNLLe1kflbxb7+bh9V0RjhXI4MjZEVLE4
hH22RqoEN8ZwIfOUiGl2IDxJVoOQW+vIpg2JY9G0jzNHH8QHVuo91txVYE0CysJi
rZTVTwSRDDGLAUzMeMpj5sROlq1b/1Ha7Ek3CWw8ZNKUfzXTRXuUcO1P5/AOMawf
TrbOYjZnSeLwajNZr5QedDF6Bx8EG97uz3Yjj6Zzo/9rtIwcrDwATAs+fDv+4zDH
QyB9IYd7gh118Q7qZC5RGxqaDd4xxpqpj+bfn76Y+FHF2KP2mZzyGeUFDuhDi8wy
lg+Jq0NFuikFiivBI6ZcpS94x2kkGyiDhadq039Mqnb7pAQrstICiRLPg8L/u5Ej
XTXlESihg72G6LK5QJvpAiflDHXMYIngb9UzJvk8gG3ufb+B/oy3VUR5DwiYHWFP
HA9Xdc1YlnvlnlDcAKStePVbHCzw5Hx8IOttsHqZayRw19NIuyX4uRpdEYtDRvgA
ahH+Uo8wRcZUR6Ns63/jpe11b0ZO8WEuFjQUgfyxvNEmzSTk7kY8sPNJr/k521TB
SzR0xud/HaGCaQXS9SfTbwEo+M8BVE343ZSyvIn5ArqvcbPiNw8Pi9K7TA20gHhX
1MmJuljEBPio8LMqHQjOZ7MAWVEYNoWqo4haX8rji9DBxv0jEcmNHsfYZWQO9hJm
COqsP/TNqWDSrh5PGRdIuEU65G/Tp1Ij5oQmuyo2GJdqFmafAb024cP6D+Nlr46D
hpa5dqQC5Pzypl7NLq4mLMPwbnhq34wTAlEQVAtJ4mucSNSJcwWtV7LINb5i3HHk
EmJKRz7z+dw9QcpfZpUEOiZQcXzdb7aZRhFWh+GAZFQN7fgjzLehFVfW7qdtxAYE
EiQ1pyPOnBwoFunjlBYQHAuKwyCTjH9y8YvbqYno/ULZoINjXOFNgX73ho6dAiGb
6pm6wmo61OI08UNH8b4h3K2fIk76fR+r5Hynu9zchCWemDVenXZ+7NFPIYRZBe2h
8csrXG8eI8GqgZqN0evjnQAY4MX5WTXY5/QLyEnUQ+TJBfAfRR0noT0xloD5lK1v
nG9e7H8Q7tkJLsL/vbkFVccPu67fpcycbBLMLgwpHW1tA8TVbfyrVd63maLNQdJA
TzpPtGQWTnU+fJW/VhY6izJ3bcgXbo/6fwXzqPIONPJi6HKeWWNY+ZOhDcZvz4ZX
UN3OBQh6gF17T6kLX2DwcNXhA7MwRLK8SQFAlNVe3ufptOhaXqeTHjUjCGLb/MIw
iZPC/CqKYnoU5nrK8lqhf0Sm61Pw9MzHNWMiK7Sboa8q0uYU4RT8G1Dq6YVZMdB6
ckhd/OWosJgpKeLC+r7SYBBSHtbKcxWsvm8vNM/NAY3L0W8desQxPo2a85jkcqAt
nGoDVCeo9XjHUK+y59d/g0Xev7TAsxNUTcgtMHG2D6adYBb5YcQgb2HYRTaZSu9F
kfWlRSkT+S8MDx76laqFXIRvDX5iBNvGb38AeQ9AjUT3+LQhjDLhHC+wgTWY45jm
RuPz3ZkyPv3a6aAcR3XLDekdbMRDr71Hr+fiBbstOSiXZbzaI12rc/Mtju3M4TL4
A1LjmoyGA8ddBnYYL6tMFoGR1Mfnp26rAqQWWKfKH3f/UZqb+yzVAU4g9oOIflTQ
8Tr+WWLQX4bDoZ7Ms0KbSz8WlpwHW8SbNphAIS9ZIJ4ExIi134yGrY3xm1HxPvUl
k/8MmzRkynIAkgmRoFWc6wqVKi0zDRn79HvrwiBRpMfMqi+hsSicnDmNGuI3tcA6
h1urmow/NEDJ+oEvmNBgPGQlqkMvAo0ptl+AJIX0SyaxAngHFOI8DAgPPMhu/PZa
baRf8X9Z2ypZ4PrX49FRju8syiMrrB2eSVh5lszC91L2YomW4lc1aoTFi4q8biME
VoEk9R3Ukv0LyQiievlJqjMW1x54CTOdnDt62CAwQvghSVLSCvmZyO0WcfBKu8n2
VAhE8/5RaZBr2KSrCjMqsCAlxLguLoiEopuBmevKohKs/87UAQ0/CpFVToc2PdOQ
QSWlGcJv9o0zxh5p4F1bstLCFZFV+pU1o4jj0e5AAscGingJ03JY+YBJtGWD7xtK
q35wGP9PuGAwpZ0b3ephoxJwozOSUU2sqcjbW8h0icyoNnTYOh3couzVGnOZPvgR
rMP4wosjdZ0jYSCPHuypxn46xbAgym2k8xqc8ev2Qr3eWoIAFg+Y+sLRr6v6egC8
SuAgkj6Vb/ZJHNT7089GadoKaOpYk7ec4wPI5gtOTve+zupyic7kDMh15csWrDL0
R9+0Aw8rGdPoB1sm+i978OnX8NQqbxB3/TCZrx1uUaHEWYVh8aJ1ITbFrm1/YndY
EAHWf03HM8x7L29IjtxGzJSy1QVyuoU4VuFGlc0wXx/G3liGvsPU4X+ew/z0tOFu
nbc64epUUVIZehMQP1KZfOHUzqaEL6Dgq3oxiuWEhx+FxXINgm7CSOLi4J6So0rF
LjNrwPafb6p8kXy7fllH+x4zJEJfEfWg/Lnz3FH/sf8kF+4Wzh4pDXjbiAkQzYUk
6H0Xt1yxwVQ0u1fgw9RsDptluwHmGe4L9j5s8xPGciRxJEayeLYimAYDF/omBnaY
LNcW6DxwcZHx6vpgHTAdawrGipA/OCN3Zw22H/612WFGCPo3WRpZAvglT2I8d3kX
6gGRthxFq7peAvj4FHqE1I0Ne86ZOEfVgybFJfigP2PCsX1DnjsL5r2CP3Eidu2j
Lmq6jXSZKgS67i72ZO0FR6HWMxOKqm7YkzgjfOsBfl4oGcnzeLL+zw8sAxtS375X
BL4aYZ1MbfUl6tbqrLOllsbHE0mDudlnGf9BdB0SQAmvmbHEdLP5fpteCmXdCHVJ
KE0ox3su47DvDhbzPjt7Gfs6h/1wE5znh3r5m7qJgAxqwlPr6krD28k4gXkd/25p
NblZzlvFHRyGoLMP9ALE5dPZOYEFdK9Ck32CgnVw+614qXeKNz4epNtBKXc8rdlx
Sz50Qz9wT9s/H9Ssl2kfH4IWrgpNDNsyeDJVHw5dd5BGHhs/vXxk6y3k3gpA2vUj
5Zp1a/A2KlYj1M3E+DR8M/Bys+OQL/becHQg6Nw5ICn62yWRGmu5hTuxWS3gIOJG
fOiag/WtJ+YMHLay0XGTGqupvmAVMT9+RbvAQZvxYR0o53TtpfNWh3tvCH+13iDX
SD6gOcYx2qSgnndgMx5VJ2GgEm3Y3N91/ZqGo+s83xPyDBTMsya0S5h4X0akTqfz
lzFgwkG8I+aGSWsNFvHw8L1l4FeyZWH6Yoo2pjsilEzP6sgnGIL8U/OOv5ILJ518
dhkCozE8sXYnBqPqCLOmfGVfOFp4wm+sQqqrnNrTKzo5ibOxJ0eSG5oPoLU2ib0L
mtha6Zx8z8E630OeoVRnx/mtkvFE/Xtos32j//4QLhN8HhZ4hYZWz2en6zsGhBxz
uoQx9/+8dIrFTBtyxLku9ZrUGLMNiwLBYs9sJiuhF41iV2gU33+GoJE+AGfrnc5+
kEerVOO4FWRuYEVJ8TwIjRBYvyw/Nl8g2KdyNdbC/WSSIKZd32w1bzyc3KHF7Ea8
E9zXySoq6AFyx83Wk7mUan5vJtHDp8r0LTg35DWWPYpS0DKw6rDJD5hSgcjD/Gxm
b0zhWHeXFPKznHB+xfFEJFCFFGLoyuFy8DGpH4WcHdUoHSUTZSPc8k1lNedY6CGZ
6Z7gBdA6cFn2Lps1EYkYhhQnsbwINpD50rsi+3YukEDwWV0JRDEM2qk8zuuLWBsk
2+Jql4tjtDoDbBvm0jz3cINKdLPDK9OEbkTbFWsf/COPnxzmSd3XYbJS/xqFptO/
LIfnFcp7ieJB1mGHMYEn2OwX3Bw3EGF3rG3QVa9HJMITDZney4WQNvsuMQF/u9Dm
gSZGYsb4SDuaDyGgOCJmBRpe2prBUhTRR2BU1RxjOGaO+1X8mX6cLsNql/U8cIzK
+RlT4NWjytdD1euts527SiFmnXXLM+uunzjgPJSysWg/BsTErCHG7Gwckh3IkjXb
OCSkWQoKwPwYnJ6lfJhQWfuGsvVCDJN6F8IyxG5fq9EkAkN8Giaygd91pEMa4zA/
h+gMmJiGWjMWamp9Ojpljfe18QuwCD+jy6W7hqEOru+S0CH3WXn+Av0Z9fqvjH9z
1e5gHaar8QEt1mbUw5UvA1tEUmF2js4fRJftlbuAMDz0M1OHyJH5K02yeXs1JdMY
YFwxYVrhXmSLSecj+tbhthOMSlj2Nf59ol5s+uSbw7deC5M1lFnZo/+UBDhNDuCK
2Fw/iK6AfM1ZDCHIfo6+dSiuhzLOTZxVK/oc2nclwPmNHUR1s15aowPJ57uaAy3o
0bIEeQRaLOVIgS/6Z0/uB7/zj+lTy0K5WMOCtmsnRCaWyx2TgbM/mPTB4rb+l7gh
8YeKbvKQ6/xD+0lhuVFjYz1yLMKIokZqH5yUDdYNRvXFqRw1ggSVG4d/lgtUC9ob
M4ag6ye5wCIBIm3G3dXQYIRJhGCdv0pHePAbUZGJr62PXyYhCaYqpeS02lsJ8GgD
JRqyb3Ejamu0JgWWwqrLAh5ymXwj+qNZxVi6oAIl8z64N0dFdOFh7vIHRdwKFM15
C7eQeRUek+7UsctTL+lvOTH3yrguHtcZaGAjz1VTnL7xiyyx3jrt6weY1Yg+qcy3
aYdedziMiVtA9LvYm82oJIKOCZ9Z28DPl0sKNax4Q+NlZHGqHNXn3+BYmFCI5/H0
mPfQAiwytn8UuGu2XpNrL26nL+b92SZ2Jr/2JY1L0bb/xxdp+COb+50ncX5qTDmI
YQ4yV8b/u6SxFV1wVcdrncWQfQpsbwBRM/N6t36BVG1rvAaha9P9IZ96P9owsS45
75A3i1aViL/hMgc1VvXb/th9wRwNmYvkRMu1OsDSZa4ehF4014Hcp7C0LBtITEvu
G7xTup6ERV3B+AiBks3hlpZKWz238Cf2olujul8wVCP8ZQC6O2is+E1p9VpzTCIl
rIvkfTKG+3zMM8vz922fQoJ4S5nFt8FC9Qt2EFotic/upx0wTyfuXYbIdDzKGv1y
RkGkrQ3cca50CUARUc/C4w8xzZ3D3ATqBniiuNoKmWyPjEZY+/9Au2sn6jdk7MAj
TiMOp/1olUQqd/n6yEToKbfKPQrKoTBcj2+dIjrjI6a1fjxElEs1q2CNt1m1bsZT
04mnmn+9gdvbXiE2wShjSAPyvz2QdWmqWHR+6WDM6S3/AIXi8RWokWqrY0sL1uja
+5+uz/7WSFFafomt4LOtgOvn+JxXRpHcRM+Uh17SN5ThVBzrmcKxf0bResa+dq60
vkBN+jw4BnJjfmLCLSfovshRYMAGZitJ8V+ybInlxuN8PMvmlumaslL/MJnS45ys
/q6hhgHXX8RuQgf0n3FeasN3Sj2RX6eiy1SL7YknzjOGQuQKvfmWCOG40BB9RBT1
kvZB7zMyshIt+vmy0QBy9lev46T8ck2eZZnod7vnNz+fUkaUVEt86M8mJLfO2mdc
zUtsfbifXlFQxa4h3uehdWjdh0npwG6ODYT29D1pVDPow0ENUZyk59dOdWYCkd1k
3MgiZ0l+ahS7GCKuRJeccQjYGqfztqg2noxR/vmxbpic8IbrtYEuW6pOUF1iwEzs
PLiFzj6WOtLFTzBVbVWjh0VgD7xy4YKNQld5Ura2ABQK1Szb0B9RBRETgeNBelIN
8Io5G0q1PP5u5efwS7R66mDz4rbktmy2C8BHULK+W1R09iTsMVGrUw53ZdMzEnw1
ztgEcEuAf1lemAno6qgtCAISJcY3DB/PkgPa9Ien3m3/RpiYbQr/SxrxrJT2Yjpi
odJOIDIx06WzqtVASN7HT4XS7CnL03QXNJirz7tNDyxJviuwSEV6vIubD7o0A+4K
H0FVsf3yDtU4Gp93T+M9RIxtC9e+KHSx7tnJhQVNeVaSRWr49cY2FrQtibJkQzR8
98NKUaYfkd/ZHbdhsLur6XW9nBGJSZ0RlOBZsZvL7ntSOAO9hLME1wr2n6hcD8Be
PQhBX2Wek+N5/h3hP2mimDuwemNYn8Dy9rv/6i5I7CgMPKlpSwjhaKrpnWHG8Kx7
ZnxHewNsxbhMLjmTNAUNki1Op5+4XpGrrLDDuhDB5NwLcHuoxJA7G0Z4BzNFfiWb
CpXc177TYwJMECwuejL+v6/WeKow8f8Mr+fXzu12s1BUtI2dYfRks3blFDgA3UAI
IjNmW02ZKMwIHuFaf2AHAgTv7FOyAgiO8wxAHSAM95YeuHfWRtub4cYQQY5z7HmY
C5FXxwBeq3MpQr3+Ap4oZQgzgW12Te4/nXdzEYozjk0hwPjDUy0YThBSxOjEUH+I
YVGFt2Z3csziJp4FQYUmNBJIlvxEykGnNJlnxjW4bsSRz09np6le5rI62IqMmZhc
BmPTahkSXF4Gbiw5QKARaamLPL8PQHOM8TsQ5bNQDW4E+TUXw2gkW7dCa5VysW2a
/doBgNOJE5Z4Y4DT09dOlWLnsV/YJjmFm8p2SeS6bPkRJWZF6gAKhf4wE8yC66jv
rRJdiRSSgKh05YOUBwtwE1ctgtfxNMZdNH85w2uwbS9/Wj5SYDFz68Ee1dlCcrb/
Kx2T/TEAWNDFCakfzUfQxvlRR5P/0PEMWU9eDKT3ZoAHwFC14AaMV6JSMbcYQ+aQ
4BFb5Dtwm+Qd78O956SNadv7GHenVmS2lKvPt/0RV/ACmbsqz/XzZoI6kqnWVRwe
yueD3K432y+jPgwHcyimGC7wa3IdZvfiqjZqUdRhTb/+xqvr6NUzealGU8BYduIN
Zxw1H2BUfPr4+s4IYkk0y0LU3ggQBQHxUYfFdmW5Q6wtycivDHEkcwUPYY0UyAL8
jI1+kFTnB8Z+SwGI/SPKw+zHZPfsM1sweq+2dBWVecYbPu+qeV6vVc4V8Ar3meu8
pPMZOX+2Mr5jzwXRS3GZs2jzEHTzDUytv8W2SnMimMA+fTxaNmFnYkxV/LTi6UN3
6KInpTvxC913RwSGyjQbO31CbanQPNzNZkAhE5+us8PHgJXn0u6GL8gaA3V4Girj
/DUz+Kf9oahr+G4G8Qs40n8Ys4YPIaBiCMv4ptl/NRRJIyy6jXnTPn9go87oCCEG
cuRv+CK5/T8N+8S+cjoa1NQf6x5tcFbhnVP2AzOCN3sVEVTU2eUiun2ewxMx2UlF
w/xJd0u0tXAC/XgloT41WGiTvGU4DgW1lc/bQh6UPZNTo/kubmmkSi7QBKRsCoiL
LumWZRiAUTJR//G02MdV/M4hLDIdjV3ot69yK+i/9nsLGb+XIADErolTODVtwbW6
olFPzbFssVN2mUvFla9HZ5XUR9mexVZK/2bSzPPUbJUt2aKMyzRxycPp4uRKJASe
xVtnFqNobklX+2C6T5Hy6sJCeAZZAJT3c17e1+5NquxaHNIssgCeXVhj+50OsP5X
cxmMS+PROj4hsPJOd6/v80seMjDRDGZcm7i6VpCb7fH2lU45AUy1yq72y4zjcPoE
sz+nsBujZGOdAEo5UxHvqQVVZFC8spMFuAPe0Nero2KlWwNbM23gUiAcMdVH5aX7
y/FYLyT5eUj+ILegAbNsPdBA8etD/Ptd2ZwI11gy9VIRwFwLpcLDjuUuCYREH4d9
39srgHRbaDsowgtSYGOBUR9QTpnTUROuX472QMOH4aKlUBeEdDbHuxepdB5x66K+
qf1WkZrI/dwePrKTANeqFaTPgt+4y6HBRSyYghK/ReQ4u37rvKt/tuK2FnBN1NN3
CHdNVDQE1mwB8+MlX/ViP1EEHvdfeqTGauRWmGTvWx52vx9q+iwHn18FcKuNI85k
dStC9JJt50+hqfPLLylBJQlwVCaImABGFQ7+ETcFk3V9xHZxW8tPVU8QxJTNC6m/
XlST2HUIY9SgWZ6sThBF1vbFQ8ZFHWFmA25cqoWcpIQHfcD/7H1wv2KiglhIALiW
O57VPBAGbLcJfMMsc+Jv4fW9PPnfF5f0cYkMpt2gCb+5OEtkxXoHVkNaa8Mme1hm
dVQ7OXotV5ggeDv+XRbFe2jlmAB2Riiog4rSWVLDUhUV4KssjkFWdKKocB0T/GoO
d4AgHBI6HrV/46jjzzNyYF8P1eCiGM3xBZ644KjltCGKWsspA8DRrJ1XhdSME8Pj
eZMyMej35wCBKgFgF9qsop++ZDW9cHKhWizlmPCbhzlPaqwIIv5XCE8q/53tLZ9M
IK9vQs9U8aqK5FKta23yicIFBYhB300SB5bqWNXSCBZqfbAxSukpRuMuw+GVZy3M
3me1H3IJLtFdBR3J0PVA8Vop9GGXRfGZNnSf5HDe7MNJh7EP6uHTa3vityKRQhRL
f48MvV6T1c0Cam0SnJqTUNrJEPhZn+aLoLPZYYQD4zW0RM9I3x3tVZF6FlD0OCvv
XWJgwvBE/lUTrm5e4C2CO1JgaWKcpNQMB9Tw+NcsV9MW8HN8/5Z3Wpnt0gs5ZGmw
XQpmWFqK5iEK5c6mv86q5K1VpYXEduyZi1EW3zXWN7hlRBqH7v7UBOUGylma25mB
kkhNH/O/cvRrlTqiVX5UGvMxymPuRr7r6ul3UdUl0eZUP0RCArHOv0vKLSSknn7n
nXdWYHtoUM9eDs/t/K+cC9BhqlfUSeO7WNqeQpIuq/lJzwOYquOzmfmgbtiRxrIg
l8IRp8U7pAsBQhqyMUNlhecm1qkeIRRAxJvx3gx3HKZv2rqnkU0ZnWIYJKGJp2mE
iz83Jlccbqsa1zeT0m8td3Sd6uryJoRKJOTvvXTklpneoNAbjNzyjp1uWC7zdoov
/QqB1hGI4jXJ48hGsIt+Ccr3B7UW3+qLQpd6b1RpE8eDn8hc73LzJKZv96iu7i1M
SmmFSf3oiXUPyWsYomle0OC0UxKvG46cg+6znK2iwCRJwgZHLqwmEoVjTUrDmqOd
KRkmUD1ALG15Fw4KEoYp1u5p163CM88Id14mBl1ncZkfVLKgUmn8B+5Ff1S3LkbX
r9BqyDuc5EzvF8JF8Z6b//kd5KUg223HOzcnFpRDSPn4zIuFtx3nIqL/WUcdnOhn
YVQOThDWcRMllv5XfiaOTXEDCo2doZGemoaYG7RQzlWtvUTx1AFe8uFJb8W9ZX4d
EaxMary/m7T1M/XoyKXOIHPpf6LqZthCbrASP1EoyY5Nzlr0GSxs8CJT0Npuw5WJ
SL5eFENoYTQOLdoOHLRUlmKM52B8VdcMUMT5t/TlRsFJQ85PQYsjbnabL9/TGAI6
zfXVunfxTFf9GKvghptJjdJT+KZGJUrp1vjuxBJPO2vuyRSpNsPCWE1rylhN58Qp
NpacshH4LcgtTBzyLDyX9ip+j8bioP7Imlz/uYF6JLwbKP1RQiO+QO2PIFWCDEMf
NuUswQmIb/7YwMfhp4hanXpvdn6iFwWbQ8PIUBayd97v2EXhXac8fyVAAvTeLtHV
WUH/eLPOJ+ccH6MgQ9nXAT7Vk0CUtZwpZjpCB4DUfK1xDzST8zRB9Wwp8QEMCggu
Avu4d8J9b/8JV5HxUhTeMdXvrHaRWZ86sNij/CzjAJAPxIccrbp+oHHNIx97IS3o
a/0mna37FI9cR3SHpvivU5q0eJ08e7i1Tp+V7TqWqa1ecb5N9tNxKbN2gJgVf5G9
8lMswkn+0jx/ozJ7RFevrbr+wKCrmoeEA/DP/FX2eIbI5LxHIWwXv+jsn/Ti4wxb
T5OZ6DeBUnAwc7r6y5Hs0L7EBJkM7PPRncUd5abug8kbTfbIjJ4ZUA081VzWg0kj
rEem3FMD2WS/Khi+vT2/3+oBRXm85LK1N/3QlfjiuJJNPD+UAG+fP01/8O5EeNA8
Ar/0055qNKOmEvyay4eTTcfYxcYC0ObpFiNhNi8xYkLdxhCzxwHiQeiBgi+tbmO1
oCziwwQi/+/99XH9XGjz4eSRGDJ8OGgCle/7oGyqa6lYQnsocdaqFuBDtI5PWWp2
3P//CYIOJqIarZFclHhm5xe3XHYdoNYLuLJwEX8uE9FhtFU7sxFFXsXED1kbzPUE
Ei+rh0PvlGsklWlGoIYy7YePiluXfXJ1HLznEe9AsSLO5XLLgdG+obcHD+pMRiR5
BqmCyFA6lmQq1R3f2E/VbNmOY/kYI64h9/51CFl2qieFRA3ImQgLx8CwkGLAO4TR
DNkWeR301WE5KlcbboIvpSmz0aE85OLDC/euGVPJrZ8Q6fQ7UOeVh2r1z+JtRt+I
+OqGVmfrrFxkCxq3fkDhmDtkm4j8r89sOlmQ9v/20MWEM221W6SOLvclYgx4UBcT
dNJweKAbxcySQY8k+vv+yFEPj7Dty/4OswlBIAF3dxcQws0k7JiyI04lcSfOTbQd
vgPZTXs27dmFeFquzF31yckgr/SRaaeujChpcW26mwml3xx6gXocak377faR+x+d
hIbrb31HhMSAal04SaZRXzkaUghwojhcy+UoSKYel1ZuPE6aFR2uBzV2A1OrGJ63
bvSZBcqACjVCc2/AIlIG62hAmNSzR0x4LTML2OpWaV3g75f3F4mayKntlCIqHTgf
k6Ze9vcf2su7HZrWIlDGl8gfADwJ+oMoSVgugrCYH1PLoX1iQ5RE37P0DWBYSJaH
7emsVozPc5uUh+eKZvRwd/igeVJz2hxXRhINRS8Qzsw2JYI4ll2Y/i1jx3KgKfQq
z+JDWUnPEI9fq3hMBX50djkkLPAH2xmQkINvIHBwkYJ4BrT9rXcQu/weDWVzjPYz
rg+YezvNlChoSwZeXJm3fiRWC3aU5UUcLw882veVnQlY7p5i6uR0aKFGjeUZzAE4
o2//13Nu11sUN8dh0Y/9E7n6ECi9kDO3hN/CCf8L5vxPcGJs0rRgbIayI/ha/o8i
49z1gf5nh3cHQ3LpoIQktG9+GK+yAJXZj0ssAvO2Ve7+oQie6dWFQxdUr1kkj14/
XY/ipBwRHTuIyqr9OD10rGJPb/2tVImSBT70OAaDilSYQ4jnxK3doLano0ndys+L
LMoYhjNSfaT3WNeT1Zah3fcVWJPT8gcrdV/wa4ddpI6kxnSMRao5iOfduYpKO6t/
G6Zo9xmv/NGoFFcgQHbmmyFUiN8mu8E2Mtng3JNLv3NRs1ru98xYSUykMeByfunG
eEZWGtTkNxCs+/Mh+fWhSqcNSHqKuMOTpSP7TREUWmYVDSja+GSm6tVwfg4gqbzE
/dB+dPKhLQbdGmSu4egh5NLRIrDQgZMbchIyiop86u5Qo9AjR/U/W3eBOWhPH81i
tyMVJyVFkBdQm8/RXSpcgfOXxugeV5OB4yxtOAN74sas94dEI0NgQiG2QlbejZIn
Z9USKXAO9m/fcS7eK9AFJajb+5A8LdtXcgaqbLOvIggtfPCSDEG4JPFGNTGw/a/t
mkuKzyC0JCXRASSqkAzUozijkDg8rXRjGeChJM5IqxyzI6o5KJqurmYNbsCS5XRX
svjBUQ1fbpwrx5HQP7uWO+jym2iXEdNUDYhDA7yztQlk5vHUcLd+R3NcJHPUoNSk
emhYmA85/amje8WllLbAQ4OjKNuAAGwgKmCQCDcch/A/7Tv06U2tMXU94Z5FJhWs
GvklFJp2N0i6NfVcywKVIRH/kwcopbFZeawCfbKvDuxpOsTnk/3rzTDwSeJYTa1R
f/Xzb4NR31cWMr48U5M1FK/ROeXUuveaBi3J9FoX/jK25Z8CKa54tZHTN4uP+c2b
bEAmPciAFgOO3yASQPO9dwpElQYy+AAf8NI9sMHPhdALNUP6yV4DzwGOpw6BeZBq
Oq72E69hVzrFjqmiHSC3JfUoQHzCHPTgPxOlnZT6SXgjtn/HaKUnYiABzvrkUL48
hBeW658aitW6NvK0yFMhZ0OosyHUX7wRXr08CI6mskRIrQtbPwCv8C+q+Vxv/o4C
qHIS5GHtf8y/s8iNNJmwnLJzaDcORYJLCznCtVmZoU7Bc93iiLHI77DXwTwgJd0n
XrmGzgQfy0pHDpD55MAjdg54cq/POFeUJaLejDZ/OLx9HJE3XhBI7n/yQWir4RlC
D3B+StVxJnsx/BxAgM/Ze2vAzZGLZ+WYXLJbBHFQNOHx2qMqlzJGI75v+dkcXLPs
KonzvSHNTTHJFv3a7xZ/BAj7Ehx+D1odcmS3iJW3WnX9+eP1VWwAqjR3pWF4iEKX
b4Pr5qMHYnX6nt535VpwdlM2nLbOs0P2eopBmkPGLxvDeVjLRfpxlcxG1ttHnKeX
LZhKC/haLk1tMVieZxHDGAHMEKo+35Y6AdXU4KOmPsFjkhh6KYdcyqlLyxEHtZIB
YK0IK/HDHXVDRi3X9absWRXKlT1mNKqV9YvVxky1DHXc7lOpjiJFlLZG3ZJ22fiK
nB6V6TM+ZUlosSgPR4thFOvs2E2tkmw0rKVwSfwNs0EFC5sGs/6lVUkNHXUuKgfQ
ZtX1usGm1rulAA9bK/J5b53eViVRwzfF3Z4ayfGjNuwE8FdDZB6TGIKi929aaJok
IGyzK94b7lQm3JdGeUcnEjQp0mvkWRCMTfCLaoMRZKGZhVodj1PN7nYZ2gpPEBN2
xNSQK6Cm9WRypXhsQBggQMb2OdhBvprVM2rUpp81TVVFqDBYB6VglksdwnKeVlND
97Jt9icZlbvKa9jii3GzDdwM1sSl3pUOgVGAcbjzsOI4hPZ5JP3THx96PMyLlnkt
EgG/yxThwWfFAcqLDBgTe06a9BiTrR8XWKBj4NhFqkg/rY7KU1iUokl76LppnUBz
fFefK8EIQKksW+x+Niljy4eyvLY6mDtPu+tUCZLS7033c/6z/8Iz0wIykHoElu1H
tsj9ezqyyLASwccelKso2Ug67obD6sYxVgolsVcKyGYYFsWt/Dn91x15kaITC9rs
yCOdCeKYuoAQ1NgZPMG2tJQPO/U1WN80lXOd7xNC2UUuk4MDHoFZzdHrq1lKwMQh
rSuxU6IMCOmNJxogXm0NU5zDsFUPs7htPeQ3UZ4oWeE+O305KVNudlF3ugvKVf9d
PI9pRRD32wPQrwgZuNGG0nG3mhKVt1vQlfseQx2xkZd5GliLbPzDXrwXSTw9KAKm
mbaCsyxxSbIZrPWOqI1P3LNQbWE0chKxKIyF9Eiuoy4YHAm2xcR7CvHea6BpxDUn
IGqNZb/r457ENcO+yE+PRwwX2Ii0KNTjCVlIHu3t+mSrBeeyRRsMU+ZpLPt1Obbg
N3jA0pzbtLEISfQKWcGTKj/+St+//eunpNw9ge89+A2adeXyiLLazjoIg9OXRnIW
Agq4842D90c5Vx9fOgI1nVA5Ss/D7Nw/yE7wGVuwt7bvSY8K8poQaZCd/Zk8hJdn
jkmcgwi4gN4IQM76A7sKeBBKQwG9e+njJEvusjc4rq58IOp7q/yqG5qOQueUm4dN
RH0esWz7TDAoUsJXCNIbaZ5K1xYattZwpvWedHZNd5d6SRfdcILgU2mvB1H6BndQ
29THoWZgHx3LbzbgBfs9cKgHGD8d3o1911yQTKj3dGjZjoLH1JT5K0G5FNr14jcK
AVpFshLFvumy9W7C4KLH0F5HkGM/sTi3p/3Q/WF/dxpCu2iurjkhXXK0RvzUU5kh
c0xDiZSlG3o9O9iUCRoF5KqiIP+niI6nAZNKO2xSJg6w2jzWT9ZcBsLEey0TLNIX
KmbsxgK59kBwudZnWREK3QIAhZphZnLjqY7uPR0/2zmlkRn6ZzWupEuL3o20kis1
3uMG2poWHXxM9UTjrMfW6GzigrxpAgKinTNK4Aq5sySoAGvM8bTGZLZBJGHs8dO3
fzsvfag4I+9xyH5BONenycniZtxBQioyCmwerT5Wq0SYgbGSTFvVm0qh0k+ELXr7
WhmS9BTruncchKsxkQhuxsSSHPG5LrlKCLPPS4SWZUdri384OzCikJEirc5qJESE
FL69Ls4MAIbXOGfdYhtBNJuhoT0vXbVoACcSvpuY6BLXYR2sUvJ8ugF09yJV/JPp
noAKr8XrlhxuIxseCRNMYZEChM5Wn8FY3B3kJHthHJgJk3pV9WB+qZfvQAFi3Acq
+wFTvs24VbXmX7LWp4j20hGQtdEE2LJv+tV1SN2FkGHpvx4JV22DAcTeBgE1LpKc
02npwVcw1Bxnh6IKZtRGJf5C9oBdpmBNtFk6HZndCDTPHgsdLe3/Y1EI0/TQi5Ve
JNj7mgo4hMfkTBZxX4yr+eVnxc3ePv2/J55KfyfFF5eAJTn8b+n1dHvj0M64qybL
s/+N4nu/Yc7XiuoxBWnLC4Sk2W6fP8OaQicg4/ZBQLcLVW5RLGCpFjvpGM7D+7RI
UOGbrgIq1W2eqRJdleBtBhSLQb8M424afXEMUXzoQxJl0TGDUOOiizEOCrLiS5GQ
y+D+fvlIYan3XoEMeLagg3wWc8H57tQ3NG5dxSv4/WzzefMt4LuVTn+tidrjBjTn
gOd9sdTfmPOSkq9yfG4DHDcKBkxgFQt7LPmBzf7QtnohANpPMVCIoNaqAekYvIPm
TXnN2XltV95Gq3f229fKsyAiFh+RBMk/7ImAnW0zpA0DmV3evRcscMW870POtGl8
WQ5qaIUHRr2zGtJljdvgz4Xyc6lfKS+UaOQYAqZdCOq3T0WKO3R4YbbnDTAhzbMs
gZerG+HszV11yH64G1cvH4rSTMsKRH6gi4mjc2kIskmZqGtjcAeD3H1tgJol+Dnp
uPiUSCQaBREHTsiNAVnTdKz+yYfcs/BYTVv8JJZbzkPLpLkvkvs574I1McNtSUao
Cb+b0k6blPR9rjhcc/U8b61m0q7ilOl7kZyklevsrJQvsUK6lpGfQ3B/w5FCulDu
lSprz1BYlyxrdxk7WtKG4gZFbyTPoBAdSMsm8O1tMF7iDI8ct8XRan/nRVDBc827
qJIO8s490CLqFfZGBADhOsgF45Wb1mVyM9M2AmUrekl3F5OahsO1UO37sA6ilR5s
w/bKzL6LaXWA1VurLadWDs39ruhloGuF11HPnhR9G2MemtLf1AOkWbM7Vyp8kH+c
25ydb2KAc25039i1M9TX0IeAZTnn0AT9OBYYpU3e8LSZlMX/4ZWVijZUGDmBj0As
jNB52BEi2Gx1oM6UpZt6rGGvV32wYqd/Ne4RujGVgHqhydt9l0a+COxsAeK49Bh+
5iOisIcK+8xPkvzz4y+6++qmsX0ky0d+x8U/Jb2iE5+uKR0Orpyr5m7VVo5A56t8
MFU+6On4r+tzXLEOrFynuSALB2RyYbFcaMoKWkGtQxC1ylL0HP6ryf9v4eSqmt/9
bgwnbEHLJeAgJVUhPae3xNENVPEkn8Oy3MJnaY0+hXK0Ivy3On/UQnCa2Dk1Y+TE
fNCpMTaRIvC8B8ddGq4Eo1UDBssPguf2NygASR6S+uJAemnQVPnih6NrYmj4ATjZ
9HUEk4pIBWDAd6GgqyE8RT+vM0KaEw7HzVYz4n9ohCEZL9tPz8jfyS69mubfJLlv
W6O9xbyyDhcWHmtL3FBLN7/deS0BBsZONlVyKVhEr02+qSwMYwcbGn4y/XnjF8nc
UtEK/SShvFGwwS2thqcIOCeGBbtr0L6+sRHlWo7+xFZ734krCyBFJNYiYZHEc42P
I45ZLlNLdkJTr8LyE5lB82/vgK6P4wjo3jc21PlmF0IobXPr7WrJy37uAs7Etnu/
3sydzaG5lQGke65nBTg6+9yfD0oQe7jhVysHvq/0R98SRJ8jprbuKXuXa8intQTB
RxNKoPHExYRHbke4KjATc59OYeWK8sr5A2Vrr6gp45G5dqFUauvpCY/vJ8ieydd3
E3cEaJdTaJzdiUs1TcC4sywC+xHW796hfT0Cl5/3MSAZeOVmDXSU7AHmHPTxYudT
OyUIRJRCScgyMtYRB6up6IAbTMIePUCM/M/Gxnyz/iDzX35CXcrxfkYeTG64PC0U
MBcLpWoQVuooZr4ANJTvM+V0cctpDDbj+DmA1YcY53MjX+uvyu0CTCYoIdeWSuCC
/OAJe19oldmoq9gJt2erZc2Kiy/xJZTfWHni9fp+8s3FUu+8xfiAYaW/cUJfZKuW
quoF1/pErj+JUAbAupXEKTOyew0Z+93IUYYCDUIesLVihrGhXzo+McxTiPPB9+CD
YIy7nW/2x0cUXEVp4Dnt5Cc7BHDYmvJ6S47o+vgECy3KDZh5T5nVT189kTtyNuYS
gBuwoTGtv89HRZ/Qlq9cFETzceYt2j5qYkoDKY6pSCTLr3iX5P37Qg8lDjRQrhJn
npVoMz/celVtEvG4eLHfNDS1FgQTEALKjYbHdlEor/xf9MpyC+ROSWhgfgFErmGN
vf/XsLEW/+36juhisxDVIEzwzUiLapmW1NnExrKKGWv3mBqE1HnmRnm5sR5lMwEs
8E/dnBNEcvdAmAinqluSTVO29UrZwJONfHkj+6lE0dV5wXuVi3MObgZt7Xuk954h
eGHup9wYafX2xkkRWe0D7W/byfUAlts1aOmkamdkkvhSKHm6zCgtjMFFVMEISIVH
pUSf0uC7l/rFQdt4t43lMDjVevikCKboyZittd+vZzVqGA+ECxcr9xJPGHKpt/fb
oV9f36JWHEncMtSYrcu60czZqjHnuPG+xfBFoMNmtfal2qD5WdBdj1TTl893WfMQ
a7GOTzOnPMMcjOUxDin65tS2SFmmUCrVhnk06jJ54ZeP9mTRmxi05Aeze2Ij9p1j
BRdnJvgMhjOLQfTQf4C+sAYU2P54xRR9kmkn0KMJ8O5XlXu8We/GK+4L8ubccEp2
oRYh12l0Q91cTmMI6h5htlCiLRKTHnovSxWvQJ7Te0wijfkeRzIpRB4OcfW6/ulA
GKXjacgAebUt7npje+Sl12cv/kOHTDUZiV+LEnvwstcyhjj87zp/hOgRVsHukWCr
aaHzyakNBNt34NflYQX+DEI7Ae3CFY6N34EiupaeHF1/OtybzTGJbUKE+kFb7FRC
cWAMzcrIPVPz9uISZNSGE8wjL4EFIf6codlkbn8MlI7yrDmy2zAO0WbuzEbNkTiH
tUzB4Nad5B9vfuuElJ328z9WivwI6lA01dl3UkWiz5evtCF/uxrESRftAoZBdjYv
U6jPU1janwGTpZuwDgRR67GKQkmXJNGGglHLZ+hOKReDSCUIIUHqiqikFPF31fXI
YRs0lvSCMiN1lpfrJV2odo7dvXjoEsvhJBXkfA430ZpzV2pioFbf5Zr72c9MFTh3
HSfqsjoPE8WjV0EogBTi9TVRnoHxpjFtp3AFts6+V2UwVTI+I+vQop7P99N8DUig
IqIS0P625qLtrYkou41NX3NwQAeJ3v6SoY6iHo6YYzaFRVVhNTzjGFB6bNk0Okl6
q3TzODdssxhNTbafu41ig12KUCu2etZl/Qmorh8y3oRhRSfWs+oQTpjtxK7gvg79
574fAyRqO0/WHuf4MsbFFkFPkmBvS6JEXCkLqGpLiYdXFt0Bobz/IUgy+7L5863U
WB4mNPauQGJLun2cJoa3igfhFJpP1lYk19vU8XcN/IWScYTbLyUv8X+5Tf3myiVM
vFCESHsXzAkMTzy3QGMJmRNcy53ZM5mTYdMsNN2IF29yOnxed39gomYWD4g8a/U7
hJ728U1cq01xJAYfeUK7/y6AFS/PfVqEzvmn5mEKxcmtjtbAqAcmWFgfgGPvwdgV
gninRowzQnJgUsikvVao5Ut2AaB0wJe2zfxhxIBehl59g2A2xwtyl/98TdXPiTby
1r0RBaqymU9TPZ+4Y/9qoUmT65D8ANutMbqtXOXBXF0NyANLgwNpM+n44buXbcCt
xlP9wMIqB+H02Glv09KiAnLeu26jZH7kq/G2r+ff9ezW8u312+sRMo4aYlhtbdVp
PEBMGF2FC+saEy58C0g16VH+7Yus+yUiwa92geFxcgMURxlZAM1es3hE2kFLRz3z
KXzBCUSxjGAthnDc59tkAAFXaUA64dqAqlqJ+dVo29OunLS+CqSGDeNFtPTSOVni
3CglGX7J+SRY5fH+H6ls/Ggzv08SIIeu0uVX2D2jgvecu/ypz5v1QGfKudwv1B+Q
NyLGw5n6DOW+Dncal/Lj4yijpOW2lrA8ggQjq2pY35vhhN93YO5VEuEgiHF7HFHl
ZyF/yPL1JQauUyjSqJi/qReFQAy4Dawz36KtoypD70NqOiDNE8p7P4BolWlbMrL/
l5lAN+wWCWabQXz54LMu/GSIDldp0kdI7A9mDYYkfQQOUifBd6uh329+SrvnEf6G
MRTljAL7QwzR9K2i2501lmF40DovtzxtrWi3dMMYyNiJGhPn5+RDs1vNlfWBnDns
yH6SPO9R79RbG3RWztSJUvnWBRnwHeqdI58Cn3zNFVAJMG/mMkHRmqabFR4Un5JC
28dBcWsLgNsHumTeG11WPsacBDeGvq3xdDK/9ugmxZC/Z8IP2D+BUJVKoW5sEagU
PA0L/RgYjGigslqAd6wpJfkpFTpIJbYKN/a5OatBUJlqjn/rAiuTDa4kVv4stvLE
xvMRWID9Wa2WljizCRBPjlEC5U1x7O0FPfwYaH/4P3yspeaWUYcXDNHBbsLEoOLr
Bl9sJSelsLmpoLXMi8B7BNDlSPRcoeNrjEtl/+DD1eEEjIFIaj5iL2qPqhAyL8cp
xhXRJFwcwmNLWOIRXfs2Ode4zO4A43+xVbNYLNAvL5azdFnrA5C+klC26UD9ERU6
boYYsiRTaaiPFyxoqqFUjSy2lduc90jQaBJB8wuY0UsxfRYFsJ/toCOHK4ODbmlI
CRytHerJrGbwFPyznDbNWjGdCkx4BK+9d7pgV2m2h/YKAeDFfAog4CO/EISFbKgV
hA9Z9/0b8UWvwsGypX+7me7PO+Zn9aRVHck1B5nlqRq2ab7Wk8yQycf8qqIOHevX
op68jSDI3kv2EXzI5eRb8QDwe7qfklR9CD9xVfcVZ3BB7ROmP0bIBPzAOxzA33Sj
eJe6O8HRGw5xELL76+PAqoywm+pT4P6UgiiUxaUbGQL18EglQ9DgPuYTcD1Z9Yf/
LlNv6sZIHND0TPT8zZPTFFjm5U+4F7UkVruxgQv7+PmFsn4DzQqm5hjnSKvqePen
TolUWAx1yR+BKt842FghTb5rK+NKCJhnysHBsCLvhNg6Rxz675blpLbpKFVBlLtC
bYsZtvWd1T8xxOASQK09be0JEc9oQlvckKT9f4zABoXm8TmfSL4TVf3WywSg33ox
4UN9ys8jmCF4L822kRyQE35kQvmpxheRJhuCgcnaN9el70ZABnLNbxPlW7OUK7UM
B14ZJIBy84/mIx7xGOkye8vzq9i7mEoXERwli30c/YKRHmXXF1u3qadHfSCakFin
QyQ9wm71oT6mUGHsAJFK5nJVFU/2TG02WZqWV+2/PgLoBMDWs3XoWGD5ro0GgqnK
M35onGW4M7Iyu8ccvNGh/5tN/a4S2XaLPLCqmFdH++q4g/1Pr8NSF0KPIaX+Js3H
7vJqcBGQGc/WRIb6tXnhcHPypV3OWLtgunmpDyMck3q7oc/VpQ0P5+BBTFJ+ogIc
frjz1EogphPx8Kpcb7nyckcvnMd2+4YG0YhUKn0fxXb7S3DqTRH68Kxm/1fxg566
hkc9N1PZZTRjZCfuSPD5OMVxrlPo+31BD4WitVCKocLDhRf3CIbbnQ1qbRUlWWpB
qtpdE5iPNMIysOks6gTeK31qKFMIlVeomf4Uf0OVIUNjq3xJ51l7ds8hAVaqEDA5
no3E7/CTC6JkV0t+RyJuPTB46P4oW7zjXN7dGC2ZJ140MBpI+7P8viaH+EIQ4QPl
b7v5oKszxBnyrrL6vZVTQyeR2bLI7Lzc8LxxvUl0oXDcIuOnWKdcEXqyT4F54Y9Y
r+0dw8WMUg18v0dhJeuSIVlnHGErzYv742YspNYJzBRnET0eFt7kPaRRKFhCXwv0
UXmWcFAFLSlUHKaF5csAxRf94gDKFLCghWkjpFO3fNEbDXUYdoHnhSlF3NTwuMgq
MNj0HZl2+LGrtO/09DYpNoOdUqaPCV8HJh4RbvkVAvgNdcTz7iGDu6LcRq7jPmR1
NDsQc3xxA5Pjgqeiyhqk6XNr6n5dZ/LOFUt0fzpMqwtl2ba7oc1tFZZOWZ5ZFIvk
Wc3U6QSX8Bvc4zzW6xJpVQ/42HajQc67irTmlfhyhXOHxaJdjSUQzk9dKkWKOsMs
Kge6wSbpXk9VQD2wXE2k3J75VNzctxiv9FeM0qdjN8BpKezsfpoQJZvTC3efE7LN
eAW7ysIbkE4OyOWSY5h0XxcYrhsPB9UAmwmfJBcOgrG1v/lj+McPcm+Q8qbH053a
a3j+8mcarzZVFUW7I7c8P8z6zcf1FXxrX7cGd2KNjIMMb15X/nQYqIGK9XvG5ymv
YCOMW8LrsKHlrTU2la95Cl2a5KdjIAD5ZPXHTcvhId9WkUKhQepfhFIufLo4wZcS
s8F+1K4WcO2twoXfibwTYvs3nywkTxHtUB+V80aZDnQF5dWItrmaZSEA2k6Gzvt1
Pu1Pknh8suHQQ/waFdKKo3vYJuNBnyBfwi2L+J6gzXcySpn6j1o1PWoNbSUpLoxC
heMzEJhoAkTiFJdl/OFFT5UZZhjGcnADTZXX4slgG9Maz+dXc8kT5yh/2nZnY+tH
0ip74Y0Vfgtk7mXSGfYWkaRxRWgySx0hSdqz1/fCvLOW3pYpSe+1rNLHZ45UzAYm
Fh5ltm7/SWmegbnXMB6E7TKEav40RvPXMGJtlUfQBUDAJWqYqDkuDKlbGAVsy6NY
BD7jjeJyB8ROdXBz+89x80zxsaW+Bq7Od+r9PQIhLgy/Zji0dMomaYEWaItmd2wr
7rCDU2UlPlrpm/sJa4dcuGk2/2U8TzYRWWgfQ5VvHKUWEmaG9kK0IFav7mpfEaBi
45PTBurE7zRdCiOvz1s+HbR20tq6pgNdTIidgg083HjUQDJpYkNdoSr9KPEGF6sZ
b1aDjPY4g89LW1QliGQq5EjyoaNhTZMYHF971C0p5hgues8IWYPAnEcLPk3a8HLT
xTvR4/dLiksIdpQl/MOcDV8E2CLuMcGHRR0jl8R+ShYsBybdO/+579SKXS2FVTMU
I+GewqJdLf/JWRjzUoY/l3WAia6r004XWnAvlDU0Aye7+LaUTpkDYo0LKxog3C+X
iChZ1Tmh+mb23J53njrN8jiHzPv+ExA9XeS5iEZwZsFe7I4DrRN3t9kPseBpXA1l
/3QlWmYOYDJeKRLn2ecI7UU5Fkt8567nhFy+FjLvs8WlpPiZw4s65J3TidbhaSZj
NL3zl6KZUSRcDL3arSkIg/cSWpL5KcnRIoq4UkJzF63+jc0+EMsGe7eCKY1Vvsb9
5ULjijcGi0CgiCyEf7ri9rzykJ5sVW9XoJAV19WftVgPg86t94ycLOd/LlOdz+Os
O9d/dKdbHu2H0E/90vSK+lLxBZnjJ/m7ZGr+o6iY6kw/eKlRDDq+0NsMhQhi1MmM
CqnZhfN0GPH7XkbCkuzka8KnkS8Qd7a8s1yyg2bDOT1SpJSRnSyZJlqZvBWTUrVF
3FaGiw+RgJHMUEYRIYeF5LxqqF7RLdmegRLCcWiC8tJx5akuSPRY1eMJ96ri1f2h
posOB6zl9gdVkRayf3EwReXxNifDgyNraESEBNzmawQnpVjtQkf2CrOIHEUhrVrL
SvWZLYtbasJZ7lffgO5ajdPBskc7AjXkT4z1LeFQJZEpD+F/rBRuQfBRKtAI88zP
a28o7dzRyRXKM/Di+XrdxtlZ/1fKZGQzCkZthxriq3ht+DbycHxEyzKfjqkaTJDe
a4QMM5DHAySM+VSkX0MrXJ2r4wsSUpfpwR+B62wD7y64IrC7U1GT96+yVPGBK+/Y
4Uq8EXq0CxGmFTG4iY0HzAxoGtRdblFOT3ZRtDu98gHRJoYQJxTQbFlUOLg5Qahd
BAvrnNQwNzxuVem2ANvWgkYR0F4AcAmsQ3I3i3vzy6+bl8d4SosHAVeY4EFoGDHi
uuHMbl5G68ky/rtXGMWik/cNYdfe5n3CLh2zb48SdOZ0OZNLMVwv3kem5n9LtJel
RfqCLEBaQR0vqbnud/jzt+okTob0lNiO+ewnpuFCFFSthp3R31/r5jCoDgl5j+ie
OecjFAtV8a6azUev+guHPN0YKsFV6ybnIfifIGFDqbWJU0oKz7HKcw825eEUiZ9Y
2reApYuAx+zOyAfQkWbPBQVpeTXzMiNbuZ2zhUkdPKrHGj8tq48RIhl0+IRB5tCv
LawX4TdvHhoZJo1YKVaKWKaJ2EmbqAzaSB6K6PFnJo2PxZVCKUsN9cxWLlNF96Od
dOAw2XF0oqOOVGnu2Scb8a7A3Q0g2LPk01bjO7zgTcD92FTocYbZ6p3bOCmYh2As
B2NbtCEnEnvInZOWluI2/FwMzWyldoFnbynOG+UFQh//vuh04aVJNMybZDQYw9jf
LEBgdt5Q/v3ymLW2Y7D2AV3z3ssZyqIRWCQ7NlzInmVH3kqws4JU/IUNSfh/SWVl
kTU+H6b2+SmYpf8m4NMupgL2hlloj8ZGCNJ9wwdAnfvIgBWMGd5gYK2B7VxB+QTR
ImB2UoiIhBgurTKCBO4A9qCOXMrg3nLRCJ7gMJ5GCn2qaFvLv7wGZB1rNJBzmbu6
Ac4tD89cxdt+8si+jcxyZJaC5fcxPFVH1Rm7ldipJ9bZ3a1XbBhww2yC5+3Klf0r
to2859WFoZrzv15+s2XBH12RNsfdsgiscPMTAk4arJBrx8kvn+6INNhX32nquXtS
TzVlc0Uop9sKfB6FiUVEiqSL4IuROa2xxqK/q/yejGia6PTolBrRNs+VM3XImPe3
kPaPDykNn3QZ0xjviGh5sM4KcSjuJx2zN9TaIuWlrN2FfHo4aNUTkYqITHI2XLmU
/sG8cM0aciZYdT0E9mVOdrNhawbhMhHQpnqLU2mXhogGtQX0BW93ZgDWK482oWok
vtRol1/4allTdDoeF2Kd2u6lGrSR1dhOoKtrmaJirZ5uEAX+e3ARRUXq2cCMTCl2
PhvsPs6EXn26g7BuymSbsok8BbqvcwKeksA+qGNd/80dEARaVvoEfHoxWUskvwud
BPCHdefLnw2XHN6zQEzLAn6v/zLTkTxEsxHj2INCRbHPV9//rmWvJoKQI18kSEK2
uad7V+wjMTihy8KgMpQ2PKigM9gzX5O/dEmbdEON5WmMAmhQEtBZBA0bMKotYUo0
FnJbwNSiCgut1ogZ3cXGPGqyhwh11bdT2SeYTL9Aw/Dc0HHwN4NatzZ0l+WjFm4N
tEbRKlxaFidM/UZ2/kFvRlMaeIf/IUP1uIxQik6r60xUhMZJ/vs01sj5vy493Ble
sstdbX3Cf3dUmFpeme3c3yi/dtIo/te394GVerv5GAB+V1k2Va2fMIcmaYEXuvBq
jFLqVnUdsoatzeEKO24Ouv0W8s/ZkRnKldZ04MmVD2zMhcUX0c5WK0Mi9tpnbd1s
UNA6v4Oc728uONPeHn8YnNXFUcIm+Daxcqi1mLSYvxAzfc55Q7MXWBsN6/V6672o
kc5qIg0IkOD4llstloAqWz8J4AvPmRh0hbfM/8JMF+ZiUvKE8Q1FPH3DIftxDom5
6YWcO8pUYMw/qZg9ORUor6Q3lS3a8ypUIHioPFArgLpMtj6vubwHC5h3iUXjfYcp
1z9Kt66Cmj7KtAbkPmQvtKH7ncho402y2rBNu0VtKvH5D1XoniSV7kZdD+VQlgK5
1m0PPL7eJ3M5seK09N8NrMkLjMxKBbfBBilIcCbaj698v66H6vjBW+tVi4d9PxJV
IMoSXyU5dxx7uw3HHQw4x43PmbVG5QPf3v5Xt/kDdv7FpJqWSKym0A4EQKy0DvpX
BuyNc6oUoMoHnVi5cg2aBBwlPI3G0vuH5A+KmrKKgromZTZE/xRD2dvpEbgMMENC
RC+DL32AFLU3iLsOuvQQVmRByDj9ZSgx4DoWd1pfMkxXVv+p06rCuL8vZm8uCj+v
lR8sCJY5NXYPhdA5QmG28K9O7P4rGootbmD9kHLpfjJVV0qOMTeOIpi0itiNrCH7
LCcKgILK9ThQ918raaJRNMQL1utEIhlw7U5pWOO9BNlKLYCEwn/uxFCe3snbwZ7o
f9Xx2Qb+6vpsxVcKFt+LPvVvTq4nrshFrdGFYFoOM058eDCYeyk8lM/eRYB8+GcL
c7uZVOzTbOazalZj5Y3agf5I7hejaGHsM1eCJK+m7cqdGGbfaEpkkfiQoOOFDxgU
WRVBvmtWq0EzlLdJC6dy38/U9qlpeF5baeZczEUCzOpsmv3qJAjCtOhp4UGZ66VS
Cm2g7CIaEq/nsMF85Eej1Iht119nCihoQiwwVPdO3O6qm0U+ZYguO+RulfItwzi9
s6oStCr/Rq00o2/SWXpk2TZMF/Y6VWJmR2Mdkyanppyj6w1jMw67cD1sVPR2BgOp
8Wur8kW9031K+nKAZP3QrXaUd74E00LTZxyLmQKxeHp6AKuJBT2rVGQ0K2U1sTII
I8kFS5Hg6n+7dz8PKH7esMBntD4ogLfCb8QbIKf4y7t4WbNZ6s5Z8/MU1apERAWw
9dH6atVXcKxY1663+JfJpHWjNLJCUTVobEtOI2nhaak50Mt7ICw0OyZFmWqlHqxn
xSbqocMQDaFCoVgVhXoHPICg6Nm/UxIFrTddTL1qgmjR4MZxg2c2ToAQiBXmfrKS
InR6AU/k273N1QWiFk7meFAdljO11Z0DDrAAzp2Yx4xUkTtjbfOcRc5yn14AQ1Mx
IYixwR3bER+MJF5mRubB45CERefpPcpfConFF3wSn44Ob02JWQAJGbOMrrCB5mfo
5DGfsliFHkxr7VVES8cK33k3j7WTajRRLjccToPbJhOxyuRrrauDDXIac4jaKNwa
+lrHGoPZrpRgVp7mMxW5zq0syba/3l0ep/TrONgxsJwtVd9xx3ZEHKBHV7ee0/DM
dVCnx7Atb0vSzSHlq0UL+fAnCkFWzdxg+Z8aAhXrUiZhy0HHj4lELA8Mr8+TESGd
UupsHjiZzpfEvyGfnwVyquT/f2VzHJYbzI0LhDFbEnSamqtWi2knQB9bKTGdjpAl
9cGUih9yPt1j8KdnkXlvnnK77XTaNm1SUwwKR+1BVn+IYqfY2cxTJ91rgBIYmdJ0
UOFyjYGi0BlDKY5WaIQ24tMs/ZWQK2eGrNl2mJOOBZAxHrjoyRSM9WmAIv2LO82B
isS3/iFHUgzGaxG5FXuiLZh1asyDW64oSqeq2ombIja5GNpRBmVGJRCotwsn9B/w
4qf5z47wkF2Fy2N+7OTucbrE4h9EriuSNk2GEMsMVAu9RpOIVX0t92ixjBD5QDP2
8MysDdD2d50TtF4dGsPY/6lxY8KuFBGsAxRCWF3x1pkRU0HxzBV5mxmC5CMUkkmF
a7XgexfrCrFlN8ubPIjdWiWZEnXZrz+h8Ups/h7j8IAH4UpSL0SbPahRYScgRzqZ
Jly6tReDVOyu547tBep43e/ZtPdI5nvbLQNgRbmnl2qich8KmY/eG70qPxDjuWce
Tb3VbraBLHSrD7GfiMQWAgfGsSYJk+k0R+fou7kEa/dG7tmq6Ooj8qJ4KU1EH6b2
nII17a8wxElZXC/fPbPHLgYeqLpdWcuw1Jxm2p7egc6V4xaLMvqpyLC5UYDAYEKk
VpcspSKTrfaFLTPMObncFLuv2Oy/9D8HsFOmlJXSLnqa7v4wF2G17dvnxMFUMjwe
UXbuFnnva/J7OWQwoW986piLoUR3VimjmuM1M9QfVfVcs3YANy8rW7jJEAGZt3ab
4VAMSFAu3/YHoOWA2v46t+L7ZjxZG88OR5vbFUoYULWtA2HP84w7oagQccTYjBDR
Ot+al2SUiQg73ovC3XOpe96DPllhS4xpqwLcumkkD5yY+WURP72xo0a4eA8Z48QS
T9zcbwSnGEdS5CSccqq6P4KvxklvrajkJ3N1rLb0iKgb6Ztb5/ab+Dn4Too1VWYW
/YfbFjWWE4MqDTiriTbFnPPx+J3KS3DBqL6asm/BQjdzXlLEu7kOTlVL7lUm04mC
CsXmnraTftFS+eNVkUgEIIHiy3vcd1pVsMC6iwz4c1bfaAx5X61sV4Y0HV5pFY2N
V97YMkB9oufCwdE47Oj5htZBiaj166PHJyzG5aTaWAHk/biCEDi+ohH5K+pyC0Hc
uglkhYctWYBmfxMGFwzYyNBDTZTIZlnuQF0GSVt2Z+ds7hduBkpFyAHK5Wt1G8Jb
l/QYd7SbB8dLAL8rykNOClNIlfvBPhtZk6T5I+8toWlH6BZf+hyLKJMwS3h3JHai
z0yHarg0yqAEK7LUCxfAWM1FUrO+8khUgIBY3GA/9waKOfaBHBRq8ujkxdoPsafD
61wqUxZ1WJ5ItFGYWA78bLCDOUyS3fc2zFfhLaUpFLw0hPvmpB287Or21HOaCS6K
8bhSJp/+FpUwSDtboQvHwQoGpop7++YZiANKfa/PLCTWt7pzmdi4uk02SA7emVym
VMiR0jSQdxYpqwrUvVyDFS98dUEF3z2mx14R26jW1fDbai/yr+chj7Y2Ji+q7BCE
gqQ6W2kGEDMeLrKrx/vU2I3q0M6GJBDd5gf3HeXxTHHgCpmJEWGC4TNRF9px6GuS
NEKIGE0REUyVAMQuESSjZMxAXqS0ALKkpXBWQZuzyP0US4HRkYSREnoxs9y9fNfk
CiY8Ns0I4qRFpJxpkC3KGPAQgAwCJiGB0Gl8d7XIkwtqGiR+J0iulkQs2eT+oopQ
/PTotMdrv8NfjSW/FMJJieA4FF4UV7R8/0yNW0KMNEx+Cj5SCVk1XW6L2nIrCu1+
YgcP4IX53nx8qg6N+ChN2rt9mkRPtZABsKrbzS9+VKC19zf6TKu4YkGQLbbFTUsl
hO7bXA112g1j9XNIk5Yq/QlRr8ri15yMpQRPC0asN4d9WEHGwEjri7XAd5+Y5Zcg
VJkXAviGh7pIW60IpiPJFb7sIknX7v94wz3U7Y8XynLSCWCdyDI6s3yrtW/H7234
jt6MP7iI0zw76ai9Eb9Jn0kUW7vRUD2+IrLoKUKjCqi/+il/eeSwLNure/62s9se
pLjh4UtK73mSKEUCbFDxn2YnNeIlI1u83+Oxx8eO2K6+CQRyrI/lmXmaHSjmj2V1
6p8I4q2iy24nuby4m9/ehYMm7tlKsi7JgSPTrA345EkGXPWdM8C0dU4PVjbpjzwN
rQxhX7a4rcOLQp7Ojy0WCt2rYE8D2bMOBx/uupF2n/QwYfFpwVaN6yBce7ZhzISt
+PCRf5iLk6Wyqn7wiP74z+uPHGoyKdAh5Sybt6Tvi/PGQI21m+LN1E8MBF334Dmf
3sWZL9pTQs3xP0usjqm4UmVWXK+kd+lTspvHRzJC4D0pJkNA1IUsNxxhwS9UeAhi
IeGKfnIDicZpxi1u3fNSOeB3Xc6T7MVIdqiZzh91eIpeM/M1QBF32SMvBByVK5C3
cvnw3rHIAUkr8YDqi1qLsf1ige7h9hQn5glsdPWN2Ys7hNoMPuGiln8GALR08/0Y
ms7kX9nkleH4uHmDLB8ckjDBM78T4NYuSBCvMW+qe+IvSwG1gN3YYhv/kmuEIMPa
al0tiXYFOWNFn8MeQO92QOuikttkJiVPt7/J4Occ+cfmXKgYpZs9fRztzOsrtz7i
2tx2liBPWTx7/UNKhQzNOWLYUj3JRUiPkFunbAZz737BevEhefw2KXtOc6rHiPKF
698x80J95SfkvmUnr4WuzERfqZp0b8sxyFwqSl3/LcbxxAUmR0fs0oqiYrhgBbL3
gQoJXnOxVUFNqP7T87Wx7ciepMIgrgjdv2lRtsC/erRb8uq51A2yeW9B30hFwm+/
MFLecuJy7TC4CSAGLs1+LzYu+GonkKxzjFeLkTYU/HalVJQ1HS4dP3Eyk5Zvrb6v
6VEZIOCUApi0uBr6W0vuLgfU0fZ2W/RRU06dVAXOCcmj/2NViJIlVjS9SZpNGrs0
GZPmMT/YmCYTg169AcnNDgbVPvmuNmez11b0mNxGDuZCMznGL9oKdotyg4hw2+LO
GCjeOZDqmMlL0aXzBc1DwNGThwva6AuVra7FxllIsey0kLKBirK9VwUOeK7IWpa2
Iu8g5WdQmyUTMj9R0vNTosWiSTi2R9VZ+WaRvCTLqehB5wVnxP+LeRLNVTyKSaYe
Oyb+AgYUGtbH79dUdB56UujIWJoJQbf3tvLqwYeqUIVdbXymbomKyalt21uKA8JP
otM+EkkVNulnHrlZoPoz+xwciMs5abzy5969alUPFvtfVgkwfJ8brBBxsDPxpSNX
OenZeDYbqRY/1UymnwpTGb6huBUKpMSCU9+uvBSjiemvHoADzBmu1lGa48RubIFp
L/4CRxG2orHcDGvKAkIIZcWcAmO6AnzQhnuNNnuAhQo1slMaJESK8w/ldImVptXo
Wcduym26JqPHfBls8bko5MqTRPcTuJKYwc+0cDRnRui2jEScomewD8A1fGrQkxX3
Z+0XBSDNi8h6EhzELxWCbjD0U6SX32W4TdZfD6ujWw7kBbAld71iryF/3oSnzqec
VJ0fF2yHo5xX2hc4CQxazAl2lS7gfXUuWW/TzTKH2UvamW76xTpFEofl5nw6crHr
N9xZ7ohPWD8I4jvlBMfoOEjsOkduyUfiKa+HI2bfQsISrkp6z87oUMvyPUf5FvI3
irNhaMp6MqubSGLk/1x+Qyj/VCoffTwRdNbrq+mfS+GWLyEqu6IDzD9X/2Nh1eVb
WGjiL3OmRglCS9COE+pE4NwZlSubrXeSQPjFK2JWOn9LI12xBvC9O94Xwr1ODQme
pb3BMqoTqxwxR28Y9p98/Up1AdpluNRQli7vpb0UqBuNsUV+bmkLLyrdogkaqsta
aadq8U5lYwaer2IQPg09Rg+N03hdzEtsLuQ8M7LAMijgW0iedSMjtfuFTA6+evc7
33DXtDhQmvO4mqz1gyV0OmqoMESSrwIhmxHTTFHMC77kXls/6Dy5RcVZdRwi1s/v
g17+9BTVe+KW4YBAjHFtY62aQCKZNYGC3o5fJHEQVOO0X0qXeRnjlfuC+oh/7cO9
/HMC4YMEs34uRiC30OXFouNpDQGqJC7UJEE8ZMC0cqDMebRyhVBZkN+0aBkfY3df
uRkoDxqETFpn2/3sEs7O1If6dkmaSbcjjDbcbS3N9S0hEnacxShsAvGPiUO8dL7f
8aQjpGoaaJQz27RJAkbc0h9pxGtxmA1eFdX8Rp/n2yHXojPbSldEEwqc2xW2pddd
ES09w+I7xY7qh6JQ7QpCYEus/vUP/eQ7G1lkG4TOk6IJ2VX5p9xOTRDxNxy6tAUA
2J75xZh5Hv3eJODwcIlloNNS/X5seaXeMzPQ8x7M5meN4h6TTluG+eX4/5g8efzf
7+JBH/BIeNqD1pCLqJkaa6nWTpM1E0xGQApFnNNnpLMlcnv6QKUnrAh9pP6plKja
EUR4VqXrDgJpzsotsDoVeLje3xnEsjTRnRWBbjukaBB8oafu0lG5E51J6i0S67ZR
IdptYcBE4CRwOPIcyUQDEmWVLxQDF10Bvc9SlAnRW3RnzsIG2wbbzlI5BcQQNoQa
Irz6nBjYZmrf5TUoDEEXD31ntIT4v0fscP57WyPlKsL4TgiM/+yRZQy6FZ5NUwXn
opjkBGP783XlYgspCiuFNmlqAUdQYmn1/dtYQZPj+TKg0U21D1KhlXj3jhTRMEL1
tCsrBeEBu49JvK4e5LsLvALBmkzhUtrHXu/hmQPHZq/Kj2t2UXe+UKkvG2VhqrIF
UzNaevOBoyRj/0OoYE+5A+/sgVF0jn2AFf6UmDCUREPxXKigrJ8w7t5Iac3QFAxK
5wXFsAeE2uLWgAxRiZ6M6lk404iBuJfHu9Eygpv8Wb1ri9vpj7Hu2dq2k/TlOphT
NNmC+GTayVR9p1WxZ/g0zuYXQFVRVtgNEStN1/kcBFCIUvHEkTDg0tKxfytcAWMc
kqwBDTPa1b4rHCKVDpt/ZcNXvZQdOIii1ZDAWXV/TT4LSB7dOAP+kMmDxPv06qrx
J2PRB7IWv6w77/apDIR32ZTwMjF1e5JSMGX5TWq8KvRrdrHsYP+de+UN8gYJ5jQr
oHZ7hw4ZEQ4rzlyMzdh7rRPF6reccfQtNrmaKhp1AzSsGP0xytzxr6MTXaMQCMt6
Sy3Hc76MKglRJo7hK9GQ+s8oEDCOEBxGFXHbATk9rRRLTF0lDQ7UOe2Fcvxr8YwJ
3dhWksl/S0j7yHft/R6tsUfH93B1AQNylONNB+lqxcyGCyicw7JrTUKrTO/bseYA
/nYGgFPIM6XZ2wYhdDdYxfUKGbeK67+T9729SD+wTbHAeIyxOYm+v70B/b2d2e10
AguKYT50Gab4P5RyC5t7dxeNasNpi4NRHh58Rreivl31FbTytZhjskkBtKvfx/fk
eFsahN1z8DtKd7X/vF2Vvjgn9bd6Ytwm31kiBrdJKa3pL44D1XX/QJqNJsNTddrQ
Mhp0jPZt79uqO7Zqax33w48QkeKu4Hvcz1lwpsAY3v/sO5Ij4s+ZEm1Vx2E3w7FC
DNaRwVBskiaz5e6r/rai8HGj4c/8HNxo/QIXH2LEjCaYXDRYQUxta7sM9A69xV+x
AnQkGY+5a6+ar5xAdq5EyrYe8795C7i76BpIIyeifxhff3mXNNQiMzxg3WDgHXL9
Wu1AkrzaZAer+ODZknwh8mUzjGAWQet7ZPWOTN03yScYgjYUqYdBgtVyYqfxhiQh
crrF+5EHkAJzmXsvbLuukkpdfkkG3uLUkRt8eOpXoNJamlhOsizpoqixge/hIsjm
bxrZGglK1+gv9cJ1aAJYHGSOFxYvmXLFwr3NBhoiTgvygnqNntS+w+NREoxFfhcU
irAFPTf4iJCyF38M2jUb4GyIQ+rtv/xKEHFtwWEQ2m/xpGeNQUjRTX53B2Q/nJF4
VLYz4+OF04yM8hJlzMN0eFPhgny6Vby8aufsv0CxJIOUP8Zdt7TJszJBltrRRIag
Ouyz4AuVzSNAAMyTWywABXCZ5F2Q1p79sBWyqo/FBL4QYGwM9REQhVDlGTiO71Te
twObvlY8h+ekEG1DP2Vg9QNmqaKfYJ6N+4CzL7DcYrJ1JX2qfZOfKdQ/NQ5zy4vv
0ICIWM+X5rL/CJTfMgLO4AqQUxhpXCaIK7qPC2mqcitxT8Cxfq8SDoAwRPmez8km
OJMZwyPkJifRE2BLUu96K0MNJcq03s8RdY2zILPCjGULyGK9NWKdupfFIqvnqlPe
LZE27Yv9fXTteEeNsdAYFA4R9iqc+u7Rka+pFlo7MKriBiO2FNfqp+aezBNrwrMJ
Uv04ddS8Wps/ibq9gqf79oYidqYOu1Ph3DCDOmbst22JZWmLp8Wvv4/5Y82h5T1q
zOvpAb/0gUhbF34BZbIjSD7zEsqQomdIgvbnQKsc8HlijLVngJGUe3A3+syt4k9Z
8+142xZa9ghA16kr95lLS/PfMT4Axzs362Qhu8wfIQAlMWNuLantrn71C02IGjm/
X4MY2SNhhzXaLhXdGUdQn+KvcQhgp+3rwJSAwpQUaAvUfyDWwf7vHTlo/eVudYmV
rUirDf3QGnYpqi3q7U1mMi7KmpycSEdlA0+YmGRHqnWlDS68k6RnO6zbt74JVB3L
IKdl967DkTvtii+LA/sG7trNABaw3EBiCJR0W5NQj+HRjUctzlfKu1FfMgUQK/WZ
g5Mf0miXygieJLFrNfybfSSnTzXKFDvPfpYO+GBbusXoxiP71tDTae1nS1zoVxwz
povsK2v+GRwUfmKlorlmnMh/jdI60lLYUdPSepY0srBWecRK/CTScM/57rDoVoQr
FEYBvX3QZkxCv21K2UkZ1g1q6ylVLpPVLDScrrirsarkraDHb6bn/kKb9+T7Y8TR
GO0Q9M7ijx9rkqFHkVQGs0K/MNzaf4TU/LFBvAmQIas7/f2bk5dKBSAFyxjr0l72
ykftF9zhy9IVhMlkkPqQqmNcaX5CVKQWQEXmli0b8xl65zaL+1WxU0hsijm6t8XQ
JQ0313IqxvfYqzDv2s8EYGsWK3vpAXiXIhtPs2Xlja2FLDM/LajWqHz4uycqEQ8q
oZaTxgFCbp15n5l32wT99Icpc1OuY4EN1onue3UKgIWqmGQmK9fdUAz4mPn5gaov
X7Fw5abVMc14Mmnu+5lbp8r4ENMrDLyPIcq8H3Mwr4BC4zYw01QEIjZZrGmAdn7Z
RT3CFqsdP41/kENkmmqNzm8S6Hrx6otGgPZz6CrLOMnDrd5PG8h3t7CfjZEngm+Y
LdLWbm+XtAwRUwUL1YlQ+Ro/dwtBLaWrjCkBfK2L1Q0i7ARcoPrJr04CdpyAg82Y
YG4+zs10oNWEpTgTNoKJmRhvTetTH1uX8Sg16/M751mbq81nd0ESBlscZfjPFzXL
mJMP58oaI9Bm6PYyIsKJzWw3y43vIOV/lq6ISZRIjVrc6yaR55gVUfBBbpbfXAdQ
/jHel+4PQQbaI64N2dzzOmBd37g0boWyIyfU2ne63JkKI5vgLesm+4Eo8xy17O1S
SjgRPmgx3yVJPqjd0TV/MhasxsjafjlsVZ7p7fO0uroLIxtkbzA8ypzZ6Sia8ubr
MNL1gukb3oG5eHC2FJkY7Zn18X5XhwsXhlbPwLv1iUEgBV+e46hu/MMQrVjvcAUt
9TUUK/A0mWoEvyyP34SdblA1/iq6N73HfHZDK71mI1j4FYwDC6DPHwFMqfb2COs1
4P8b8LYuXZMgFayC8GiGPEzbCjxakeeMbG2/6jAZv15ti7Je8SIdOOhfN/SWrv7L
9hvi8KSrP6rDIA+DOPmvTBc32N1ABODh4hs0l6xKT1Ow1JWc/mjeSWfefYSeevDW
7sFCn59zHkNZ/yGS2U5evgbSjBW68NTq7xnN94V76AEWXRyWkPRdW7mtXVHnYYjK
sNaZ7cyNEqJOmXHNBwfUunOnTGccjp2cMN7ig8i4PgS5jubxbMVW07QrseC7Gw9f
VrMGzbZ2g3/qQA4vfkPwxT+OjCiueHyD/WHX7sTALuUa8Llw9on23IVUHp9RndIX
75sCNn/ai1HPoQ791QVd9DUni3hrbcyT8r5mHfIOWesfAxTv8W4lMrs604XNk2el
GVyPCIUA5IP+vK2opWDKDdgjuc7iLefQ5wTJcdCCF04R7yQHeA7iel/5JJiwscJG
hKujgRazx6h1YaCTwsvd1N4oEmjaEjhw662UBJeHdFK21p9koqrEJC5+ndop88KS
bER2IMr9Mex/mSaem+cx5mqJUzT6smFtFn/t8203HuFY2CjhKqL6e5jVrs3Zyw1Z
iXsL5iJa1bjlIqUzwov2Hmkoi/EjbOo/WgEpPcnrRH04dmdfcb0OBGUVtLm4COaA
Ifvt+PN2jBOFDm5B3QSe+wLPclZJichCpMgQYfAIkYYPVT2Ql6OIqGVIJvCHgkge
l3W45MKhOh+Pu4Ap2Uc1C6sL9tOO+ZdLbzekQynYsSgkd6E/32Yb36jlcyzYO9fa
8EeqP5IsMM4uW3gyDdUnc2pc5od9p8tTMrUghAQYhpzmjvjzIj0xDQ+XY3mXv6xN
gJ5bwN2TNtqEXQDt8HN/IMTUfnsM5RbYMS8OLMeqYuS0P16ItKoXKFszQ0bENYhF
fCgsrlV4RYlk7DLK9zd79EKh86XCHeB4uC1O4LCmc1TwTS2jwN2T2KTivXEDr2Sl
SMSmSG+UEfNuQuRuf3fAiVNAic3oKE9xtGugBG7PKsm0Y+0b3vJ05nHqGeLqJRz4
8XG2azAOxmB214MbHdXvBU2wWuMx5H4S8FWAyJguhF93v8uaI2O4wKI0YTcrlemV
mgYHV0Qj+Lj/ByI5pOwJiArIarIQoVu5EcYvFDWzW72ApXcmDIzuVQ8ySUsqbMrv
6vZ+SyIurGx+OmbaBNCDKtVqJCvMFF/w89fCH/kdmOY5BVEitX4SaAWhsrgRQzQx
pG3PSq3FN5iw8ihIt6HWg8Msk5z5PB/S9eLSHKSELVJl6uvyIx98msSgN3d91Xqa
nJj3nGDlKg31lHDWvYQMxdtskN5jdLD0MUbLfgc401A=
`pragma protect end_protected

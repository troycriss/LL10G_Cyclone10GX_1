`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
GNKzEqQw1csiEJGDwlBtTqAHvXE23IftE0lZHBqAtSAt2Oe1VIOQxRbQQVD9Se/c
fD/4DlXoy8ou55jdRg28JECsOkD9EeHEoFfcVDP+2UdCxsuRm6rmt3qmrl9Kp42t
Pe9oHXXL58Q5GnTAc9W4rH4j7vwsIqYXafjtqnaXQrw=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 32144), data_block
bA1WuBDoH3UJljbQ3e4e+rA5UI8srj0WLbuquNd2mS2WFnjqZntki8+Jmz/5DRlB
9r2Sy7Wc9zMZTJoSAWY38WLENU9hl+K2Y819rU4WjEt6eFmwaobBJu1GSGTUXtIr
KoNIGEPhVgCEeUynr9Yd7SlLdDz4wtS86feOoXihil7j5AKw4wZyrGgZ6WHjCx2q
Gh18iyXeoIRx9bsifycFFqG+hmiPiz7tzFDP3w5cdnp4b9sfN41dSzLrfpzlo52T
WjQKAXW41+28nzx3cxRLrXGsRmZq4uvKkGma1tDOej9lqqge6YSe+xxvBxwt98gq
Owv1eU1JvZLt2hiF4QNLanf++WVHnMUfsnyhnBum1jvJcq7DdLY8BvYE00uOX5Z3
yYgFkq8Dbjhj/RaV3yIdp4+OWf1cQMPZ7LHYuI0qOay4Qtgypc3OVrpVxZaiJB+V
rLZ1bjf5k2R9WjWHxutcnC2ZYoztSswiVjEryKp++jnpKyz4mvjmWn1i26DngiC0
KUJIdIh/lVr0pKdYJJQfc0Pp9nl4OT8K/sDDY/CtYHxPcUFaRF/5Jus25ssnidLf
hHz16fyJne7ixxlk46w1p6kUz5mS/U8tz6j5c2EIo12+r/4oFUfO0x3XleADo25j
Hpx12sSxbfkuqft4kvt4cO0CubTsEp7wuUnkF4XCnhTU/lXVgZaFuWsRtdEOangF
81xyjyikB5CiXEZuVjXBZHyXBkkr5Bv81bKQZzxYTASxGBg0hm12PU6waHO+dyfV
bcrGCCpa/ggcNYdtgxoEw+C9iKNdvgLRvYZhEUFZKh0U1ORmlC0av8zayoc1ayQS
6ZgDZjp5OXvGKIypPdFKnjsMI9LaZNWs9C72t5mt51SeAsJ5q0+hnkIudJnHinyo
MZIw8Khlx9JL7xZhdc9jgr75fU3g5ZKhEbtg57sB4cxSt3Ti1Rc6OQSc74+m81Le
lfVjhgEiY5ZisEsAutrMvhPFnnzRepEkH6WeINzIjtyzqi0ruSqndtkK9MF+G44b
/apdT22xFUsIjEoYFBJOTTvJrToEGPQAP/eLiNWFiCH5ugO/TD6f0hcGGy4ZFPtN
L5X7aUiNz+uWuwG6QiEPLfEDD0iMLbFEt5A9izwlVKLauxKG4D1kdVwPz7yQVIKz
2ByxzrPh8rdmsmfQ6MsEmc50i+xuIPRow1qCIKq9Dv2ID+6B3ZKRKAoaERVQgAgA
WQgIHzo5q78tlH7jAtgXD/eq8gQwSKJWs7s22mpWpkLgRFb6hxG01rotSwdxKT0Y
HWHaeltJqk15jnU3U6RfbvbLq1xeeoM6og2+NaezlZi/VewUz2OBImgUYFxj09Q3
ZGL2/S8Fu5niKD81hxQGVZi8ILAxHSeSCqD54nJHbj/J6+x6XYD8SQaLG83yepa8
xSyv5H0Y9CCTN0KP0h40mcFQ8bSiaPObCpFmMi36LH3byIsleberVrWrqJBZb89t
Nc5/wFdBVMRY2B4vWlWt+x+5hHW6/dCCVPToLprhVwuZj7n/tTUphrYEN/B3rT5A
wMhOfKJpRa6ynGHYHPwizOydP+VlsuXyKeKX4yCe7MBNdawv2QsXaxyMbH0dybfo
Hjrhf1FLvHa1z8hZvbhHeXIHznVZah8rPmrpuF/XD3nI+OpGBkPZ5pbSSUB11GGU
b1rB9+HUeQX9mMAl0NDLFZ2/Sx9wSzd52+O0rffokNjADTalk4bQhXPzdw32TRN2
7LFEdzgKsQSic5/f0d+evZxmaXLLMqnRRlYjasMu/wmF9iHGBX+mYFt8T50OoBdK
5pW0xsGGqvL4/Kh+n+//NuE6e0oq9BGm1k8aIHNiPhkCFpIBJWxfRvYQUjzJ1TgI
9nuInbeZYB7IvUfNlGcPVZ2rK4CiJDXrGJXwfwD+ykWTxeeMHR6ZnDdPSxnQoYQE
SGFrL/t2nStot69e9wZjAFOfwFXNOkuv5rKN4eDkFXqU0rnSyJBWWD1yN8pLNMZW
hwOdTsJtNMnsFFQCRsRIFPe378J3NrRpflLmGgRwJQU92LKN/u7poehiuGonU/w6
2SHIj+xenM8oF9njpTIGmKt4jaDfdKb5TQ4IjcEixDEZLuH1sFLna0N2kwmBdfkc
CijVzU0VYED+8wnVXYswgtI/F3M+s17BImyL7Fr6bwUlWmSJUv1BGRJbEcH3obVD
OsSnHemOXHfcmyMWrhPGJEHsX0GkAVy1ocdrGhwpOBBFrgXeTv0+oHjj0I7G71q0
CTgUMXWqn55Fq6TatymdTVnxZ3deRuRuGwS2xRk89QhYQidvSy4pAXBuI6wwtsPR
60gMT1Q/qT2DnedOH9rzkbSeqjfeqROddSmhDTiKr3VgqrMQd5FxQh0iBK2P8Qhn
JqwVUZ2bs6mEZ+mFsmwfhd33r6pJPDD2K6k6JL98xGj1pgiNFQV7SagHr0FO6jNA
b7PBcM06I+lF4xqt8PhdSfFPMUQQES0pf4U+DBu4zbbkQrskX+hd34WqSE1+R6j6
bt2nNtDtIQ0zNIDhYS1/qPeyUf63CKzYEiDsLWI0IuA3kWGnylug2+5GyeslNFHN
NqOkeWkAsimqnHoqETDQSyFFhI6wPHthlR0i5PaiXPwLM6r6LmIyRNTTY/RbN+W/
KyJ+zslfDEzDOlH8uGYbab/Yye0s8MvUhvgsVF1W9pWr8T8uuzBYKyYiZp9GS3sU
C3jIZxTCECf4UiniL+GBjLRDqeVdfMcVnebidlhVPizgufiShxXkP++2584wDdLx
pQ+z5H41Y+S0lXw4Pcv6LC51us4ipMxHVWAeiqHqIjNph7wNW8rQH+OpMnbD5z3B
4ibKL2oiSe9lkiaYuSY7/QrATlcUWSlEJIrvDOvh/CLFc+hiCm8dlBjIMmCx0vWV
1oY7S718QVwn20Lh8GdD8GtG5nMUHLFQcDot8uCTHGjHepK7lW9K24URBARIcUQX
Cb9lEjZfHwvy6F8lk5DPjFTglITyUfXrFBt9oKGTA9iFzp5ixUAiMUAgXY/ZmJRj
tChx2VLxPvk7NLs81X9eSwwqCQHNvyQ1wbQ+G/s399/DnI71jKiQJf1oBAzQ7xcB
HLHvS/XYg/AyvBL46CwLJtj0Yk6i7VLH5FCuvaxAHK1BL3yX7tlSi3OXTb47P820
ml85QHXp1/sX8Naofregtgy/qnOWRuVmioDovosNKX0kiyOGk+AWoGnA93Xo0JmF
8WOhAN5m385BOoOSt2A3wXEOt3FWvYwnmMWxN6L/6OkSmzwTUyohhHbqvSNVU5+X
KDoCO52v0Tdb34d+XnbJEyctECkMYhivb1FBTomC0vpFr8F3JWY1CzyP5rvoQmS6
4xiIqX8wS3WXmDnwF3lYzcJXp1mb8rgsBVJ9KffM7CGTlWdNqnIVT3u+LuzlDXI4
YA3Oc+FHjPyJOaxa+A9Yoq/vw6ctDZgbFBEloryWfotjBtr3ET9yjxjUPnPEPt3S
iuVMF1ruLynmAuywva0FcIh6ugZBhSJD+hpu0oo8vycyYVJ60A91Esr+LyKI2Zfj
WR2ykcPFPwwAoW8VIEBHk5HNUiUBv8dJM7COJRS5led8LpX668cFJ6ZOKZlzWf05
8aAR/NQclsPU/22KNKPk/u4kbUz4XPFOrFBcJN1M+lfF4FNDUa1SHORtSPEP5ETg
w2rBtFPaX57Uvfw2WK+CRDJSK44VDYbu8qT2B/qLrRQEIgDBth90M8vEaSUlv2ZK
wa2g0AGHxBOh3y/IpKRJ/ZvVubWQnAkHBzgOuOtCHQsav+Owt8h/eOKd+Zz7HsBW
4QTOVD7RdJnUfOudc/u08Mc/qBLjzvPRwqEPx1QP9dVKdYRzQIXuk4RN9Stpuuot
1TcVumbnBMM5f+w79UdMalzPTPWnjDlugEnE6cZKd08NS+HrE1kXKdkyzx5iVBIX
z8+bWktPtyWyRbhLXEINb/o5Be1ZWj8YVcYLj1jIs6FhIV7vo0xq2cM2YlofQIA3
FJ50h8Oo+q30y5hzWT/ho7q31AptW2ZZogUNsyjZmBhGlYnJ1YURJ4joCuRLK4vl
uHBdtOw9O1IyKDAEoGxKa7rsoYq6jrsv6ioNtq1It8p5+Tz6PL4SmHu35jtaPjOB
jM0phI+jMQZ9bv3Xw8jCP/cbw722yK2P++3DuRc0WAFlG57vKvBbsre8euiw1alS
aqA7allKqq/LV2QkJ3W+SM2WiLx/KhQ6s7nAtomaeuhEEeGXFhgE6iRygW147JMN
lpCRN7HLVoMxSS3Tz0ol7Z7Qv+jShldAKlTbf70f/773mCruPbXof4K1M3Zg/mFw
v9F66s/fhLNUggXXxO9vfURjD5FdLEj/m5DIkgFRl5EjNJjFFp9sVDHXZQ8RSvJg
rJhxWZxYSonUrU/jCSOVEZykco9C2hrzR93B/mAm8GshfkoMwTLAATlAHc3dxSh7
Kx7Mm9BE7xs/fv+9GfW6RE2jXMX+o8SGQhMFupwm9if7iJqJd7B3CIndn5SLjjj/
xb6koZpuH5/dyjacBnfXJtiYNHkrWVJxzSI+OrBosaiLG3t9DLXAK1IqI3dDhaee
1qfd3qTY0opT1sFnxrUaOxwm/qyHdN4+FMYsmyET0bC8omiqqxJXmxB+ag15BChR
hA4+ewv7EHLqO73TZLB5Tyi1AaOb8ckAGKJlyL6+x4P5BoTVECyCcB5BCW83Y81O
BJRCrcquNS9tcsEpuyweTGZ7go4B7YzzQurNJc0Me7fPeARRvMWoFCpXT4V7x43V
fL/pQhK8G10VnnX+Gw+u3Ay7HWWaG3JKTN/BYoEZOoKomkH1kpsJ68buXtKZBhtx
0mTSMVLiZxce2poZ4PVrBqZSfzOUyeYCpRfqd4wRiVIqUaEpTmE7G+dVrT3llMpO
MGpiSAcOSE4Z8wm/cJRuzDhZp2YnPZ1iuLiQahNKqucnQe/1sjPNpAE5Coy9dYFh
UrhjR+FqIWqmP7JVLytEriZElCfWbxgjtc2llkURnDGfURksVpKpYHNf6VJA60vW
8n0x7zAOqJ14XuKR1lda/t5oey0eyH0drVmTHa0t2XgkcqOZUajQEjyXCycGyY2b
Okuav5DXGkME7ztj3yiDEalfGBu5QvJaxHhUtawj+UU1q4/lK8perfNoLNmBEGR7
+4RdrGEFcC7SfUDMFa/Gg48UO1W+d9v3gMLA+2Q5ZX6JDclBFVCSXVw8cD4i/mfb
s+G0Nvo1WxPqmZnrej71x7B2psvHbJZydaVobdOgeUiEFoMoWH3yp+Fb4BqayYGr
KzLYc4On3MoZA6mWlN+UJhjNmvtz0YCJYSWbZcu9CDr3i7LGKuXPSO+jhXNfj3EH
FlbSz5HQIMGJi1DGtivUnlQPfovO7c6GqfRCC4TAnrIbOWdIGwYaIIY0Nyba8FYb
rrQ9dsXsWxslBS+5Tnj9IZ0IpESZEWXBA8w4Zp82AAEgtVqrLM/OIE4R+10N+ECz
fnyZkWPdcBIV8nVu+SR8/LherjYiIK9Xhsqz41J2ress7FFpe5q85pYfaXzEiZuS
TtWtI6yn5BYmJ7urJmRVRKTX+rnpIEYbCJsUAxVVIOQh/rlTioyeTqJyvOo+V5/t
EytTmjnZSQ/Iv5c31dcy3NUrN89lTwHpY0A2horbanpr6gfw4mxsL/ZDHqAwJ4wE
BGZx8zDSMRxSV3uCVXtOEL+AYe5uL8AQ7SbrYwVFFzTrpjZt6QGd63iqU81CbKmX
1EU1UAaSTsXXff8fbEWALf1q5fGV8kse6Qt7dG3L/oDFqZA1GUMDcD4pstNsGU14
vJ/2gPkNVyHE/xRM+tn0fooal83CtB208GmcsdvGZtgPjGv9idgWGRNFK73o14NI
MQnp+Yzp5OgwtImIVlDFaBCAXte1svr/WCg1Nqgu8otx4ioMNZhGtdydQ2aS3uBT
/jYxCuFpew1F10BqJWxK4qIPsuXOmzWm3kUA0BN84B56+9LBnzgIW9EPWa67+eTE
XP+ZnWQUWAozrSxmYR9d1th2ZGCgpQrv2Q/yvgO35CMdyHDwhlx6frgyS7zIXL5R
NGSFPHGl6cwlmNGyAozdSJQ8cVGJcQBCNrQERBsVKK4IeWDPt7kLSSf2vWMJxeT5
5MXOkfXUcsRsAcM263xK7bqQq3jFFCV9WEQB+mEDvZgIkf3MstXgFP4lth4VYYLZ
lcZHI++k02e+gO+UH3GVwEExDQPZAJ5k8vCGBfMfUbVIF5X5VrRwUBAtLryE9Y2Z
PNWa87W8P6VnKIDiOLzp4e8IvugTSqUIi3TyJF5MFQ7ZTmTXcdLaPLLyDGur1i7G
31plt/+fXY9hO/PKo68SjnxQ1iqnpFru/QeVHfHDldS5+bnKrddUF9ojo8vurCxB
ut3a7d3sxrcLjjqxFGe2bswE4R6PcqiuOYht0549aQivT21OwDX+hvuM6mvp4PKe
kybX6UQHXbV9H86NaMcPpVt0gEm99ukGI04WJXt30bw/5O/3nEwH7rAemod9zzCt
zHQ1+VlbJqIk5SYv1uE1YkqEGwTa2dfRKnKmOHFFiyRtqBc/i2XywQeROwMInjE7
zE3yV608O0cCLeW7WycHqUOStjiAFxuGjnzaqcT+Z3ix01U63pnnqQLfTGMOf1ui
/MtT/APMUFUOyAzevoiPLhdnUOZfzP6OmFEs0PhIPHSrpgsxFoQVTgD2QAltX6mZ
ZmhnfI23z49sfW0NaoOMJB8g+FtWkE5eta1jxxiHkH0d0HPqy3GeLwwtBw07sJU0
xoBj+4K+j2tvdoX7Ulh49E0GNeKfoyZkiCVv1YWBHv3xAn6711xJwj++TsJH3pZb
Pu6YmcoM8uP1q2HVAPs8aO8TQcHA7A0EEqr//5MpAZ1jbMLW2xdv7qLt1qC57FTJ
WYn2eWeaqm8uGPcCNeMmVUzO+jCQhdFgFyRXsCqGxSsnadGxUHeNpEdWcHVtrYTb
9lASpnmMQVW63XrHHDP5U3gWwa9afE4XBrq4V9kPLYUTJkqBmiSsg3XkhkEQv76X
ddg3f5WMieUKR3edvL4oKY+IqFODIumYm2n7Taiz7MKtdhPS7XNRpcw+t+zMhPy+
h87aX5iNqhho1v3NdPLsqR5nV0LX2CfeaExvgSBXf003/lwbnmYjxmiSWYwAQoHI
T4nSXuQJakrzAXiE5BcCmP0WIcxS6yQ7tq4NhCJcpqyTpGJOZyOFQwwTS0JyyxMB
ZZ7T/uAzNcebuFY5pxi5BXjt0YBCeBf0ATUFiGwa/Ng/dAp/nQSCLcI88tP7g4gs
Ah+4FOLwFapiOhQyvY6UA8mSB8k04uwrr0NnEHFmISKkjRruN2hLHU+JnIXw1LqJ
xZuJqAvy0qMpWhu+BH6L+M1dw5MqIe5OvoLq2P4cZIt6lsfKu9KR6w/mGkwKPQaz
JbuzVHwy60JaGQF3Zeux66rPLKWOVXKSRPLCSoGncCNkPnftNRftTFCVMwOQpxUX
1mdP7CPrhjfWOTRW5E45o1e02fZmoc6fEDnzAmUQ0/DY1VwApfG4sZ2jO6ikUBc8
IdXgLDa+SGjeak3dQo+FZ4KZcet8d+KygmWi6SVrUAc6ecM+opWZAa3BZECo+Vwm
55DVQQDUhSoEWqEFeZVsKgqILbPn1DGOTLxMRPhM9HN0YV5Lx4JcPssjtBW9PTrI
Zby/etvbPEsEyj1VxH/vIaPhl1usmy1xt7UlKKWBUwg2IdKhbW7BRTccjW4xoYHD
j5dD8Yc32hHQp36s5as3mE0D2ic8PUsPK6BK5cEjEYfD0GCq17tefeh29XX/boXh
FZcv36+OhS60oW+seShWoCl8/5J4V1PAcGyOM1Pg0ti5TJyQiK/iFPz85r6+1FZu
tEqsVCDugeDvpLQJhRpGdNhUe1fi4zInt3pdIyv0YTvHzLc3LzV71vird6vr8Fup
YXPbqde0rWu4aa7N50PC57z7uyvZrCvZ0Y1Ft6YHPtL+f8YAhmifhJy2cbnAPRAK
t3ZWK1pYruh51Srf4cXCHJW46gjtqYRuQKhC5XjxlYiKhqQqW+0+scIZ7N8GLwHt
74pVRFkPCdw4zCBF75vk6hE2jUIS4bPdER+empHmF09/R/YM70t9D7RFuOwEky7M
9ksdoJUpo8dcTtebbpIPjSR1y2/ro4tt2rOHokr9+085SBzaFpC+G7LwTTMHGuV8
S9tBQvP+N/v96H7AYHNHQXEFxw2GKZRSEfFZc1bkqu9e6ebq8VQLwUhVimLlg6db
LbiUtksVGOpo5a8mBwXkzbDdNHTf6Fqroesd9Pp4sVhK6QECbN7eTgOQ4F56PCsl
/LzEONf9R4K/XjXjwxQwej54n/YtK3aXbzLnGjGKrkfDXSARgXjOXXyY+GaRFMh1
Iqh8ScY2iU2KNUYPXoLJA/Ph5v6mla2IUfUPRo4asy2opnLLIM8Qoh0FEmXlGV0O
pSO44a9p5attFVjkeAAc+Ee3K7Vqpg3YlCe0rrfAYIPKdr1OUy7HWQDKHuuhCbtz
oflmnQLgUPBPiJphicdtRpAFBNEDSCu7pGteak52Eex9uWDga6qVRCDZxrjrXOzX
9SN/Q4zKRCESQOlWmVre/RmqUaDrfF2fvpik0zvrmigchh5qtkxJVm/Ik/Ztvok9
1N9/KrPnsjkCTN/eeImHrCSlxkNcS3PHTjuaJ+mZmdU7OVywf5CfySzx49tKAhf8
evw3BvzR32Hlorm7H8/iQm5vHcEdB1N0XIF5kQNKqGD+Ppdb8X+i1b6+5LEXXtNJ
PAVAc536bbRSfBGq/8lgB4jntMTv0kLjJr2h+cmD4x+9frPmsX8AkbmdHNIoqKxJ
6cc/FYQ4KXKA+4B5BzkjkmpTRSjxKxLf2mU1YolER/OdSsBO9fTnCoUtuo74Il/s
RfO7SCdzM8VWnDewvVKCyO11PIf3B84myocstY6aKJKvrP1JQtMktYaw34aqrMIB
wB0NSFBZlup8QCoaX+RY8HDyfeBAHt/UiPmoNAfMCT8IEuGDeKJHSUu4nFi/SbVy
zsY3QSljsqCM6YKOwesqneJMGWi68R3XAtvBcBKYGJ8u2Y0duVHWrtEjwMvPzdZK
HdiIfxa5KiS/v/259aWMk5bxlANd0+Q7ave4BxxjgO3tB0+f/k41FOXVbzbQPEMG
PuDzwrQwR1h5ptdITAt2r4y9AnZBkYZgVBfUbmD3x0Ylzg29bhtwK8RfVQUNDnT0
bQ7dcPpt/iFEYDd0VfRYPOk32pGqsWrYn3v0bMOQHKQYYXMOTGbCZcG29KTs6mjj
nK8tE2wu4YPTOVCWM3irOFE+M1J37XNWSwldz7pXHgLYfEJrucuaNstM8zg2gBuN
nvTaQtwrWH52KPSY1Wnj3v3Of2V+mfDpYsXtUnarjrg9azrmBZfa/x0dtF75R95P
vmqMjt+PBAgUjKP8p7Ml2RTBzov5y2SYEHPBmyfXtWoVEPWrAxSX+dmJSO8rXEwa
6f5rIbxx4xx3l5/3/XYMRaucYH43aSipQhlIUhnH3bY2BfMdXS6Ak7AXhg0OUdkh
6v+a9cEcjxoVDnoIUR2oj8xDpFlRV+7gRyIPzrjL5P8Z+NMMdvfFeqD6XxXtgGGX
s3L+3oGcAtQ53ITp26CYG4txzClJur87u4SKt9xIZ5oY1sApgh/MP+XHT6If/ZCV
XD+DuntJY9GInb2WerC+DBsfjbJat0ujnwqi68ebTp5GyBhIVZMFPTCmW/amIr/E
W2WCzcUwWJm6Y8jD+fydA6+zPJVZfsiL3hvo4mqxowC2AA4jsx9XGEIfFY8cJaZm
OfxIvEENkWoDQ9DgcF/8K2kiVq/sfpVXYszBM2q7Fr8Kg90+i8DT/wyEJEU4ahAV
mAYZz4Bkh0AJe41oVsCFmrUNJkbdgCX9Jog/m5nfRanMTzD1WX7qdSfZWgcsQt65
suO5ggkq20mkaSA448vBIs+Jbv7oWKhmX4OnFAjWTxxP4WXAuZsbVRAlhCMj+ovi
ZridZJw9HRU2K5v/mC2QVVpl8TQPebry3G3A/wyaSPVzkunPtFHluYyj2O3t6q8g
4Dukt71aVuJvfBtfE1KtN7oQilTAGmK+Y0JGMpu2WFQpYIwVyEicIYwrnhTIASiS
DjaUVNEnA7WaMklu3Rk6YRIWaAj3nxr2D9RvENKwLcoK/BAtdb4XdlV6SCo6KCQl
SNth2+bhjKj1P4akXjznAGouMqqjNPW3PhFIHEKa9CVw0bxH2fWbzLO+A079nSWs
UWHb1Bm5s9KIbXbP3Kx8vkBi9ICD6BBXJqrLJgQ1VqB1kEMpA7UvnCg/wShQfRne
RX1RTyFWFrjYhQ6T/E1IrxjbuXbr9tNKdRLRioofX+hO6We/rWW2gtL2REPdcG9A
uhvMv4PPKLAbSY3j9B/0vbJOHExoQMfVMoH+VPwN8RAwK8IRhms1psM3lo7YKK7/
+tlpwxxx/hpy1In9JbdSciGs+EpPiQaGLdUAEg9AXvpoYIWh8xAKv+RpIytjLJOp
DZi6C9e/QpzNodQGOYOZuD80IUE+6VLkUqESpNV490EMLvQK9rsW/V03Sr82yj8S
lnKf2gEDnGm53kAwfze4lzwcYKjmQLsjtYWqkHUCLbSdUYvcO/TuDfhRdU1/huPV
R570FEDpFbZ29CiXSl97Ny/sFLWADGF7KK1s2OcizMkkkiEU3DI1xzvJ8SfKo5D8
jgeoldoGwwbpk+9A2ARX1pf1hCDQhByeEquFiiwnJSADq1rORCIug/XT2EvFwO4s
Z3LCssX9ucr8ijb+hC1FeXN2uSwXQR41QjY1kpQtOeWXjS3LpgieuiN2vqsBbi4K
lQ2TtLf6Gap1VRnVTpzJuMX0kpvx9mfkHnJBdZfwFSBEhOUrj3uDLRRqZ55gZQUh
ACBqOwcgL8hOMNJy0aJ+jT9Pss7bu8/BBlBO949P5E3b0T9VOpY4Hv6s4WLW10su
YQT6Kyb/+cIXojZNYL4qVCquy1U+oy3x54AiDAmZk5cuFJsKGm5zcmAO8N0wdmwg
8RnX/YRf0/+gaAuYkTzu79v+ii7m+1Cadqo/64J6BFq23yhusyO1g9+1fcGUEhwA
UjmVI4cDjoZQ/Nz7PCe4qdBiquqUdycqHVlgAGSDuB8eFXWs5jPp3vwqAPmd4KUI
2htqDV+zHnsMggqvVfQ4kUGgZpNZGUm1Mu6O7SGPemsY1JkUqU+CeB0r39Jeqf9G
LzuO/RGKN5fXWT6Zmb3gCbjRBGtkcFzMMw6JAIGqji266yclqAtsmc7p/hYhEgyi
F9/bW+NvCDPKxxrCWx3J7KUHP8bGK9nwGR5Z6eUySdJcZK0/N3yHLUUG5fREt/HW
4bmqtUrfsV3vRLfzdODafwf0roYTqSq0Z/1a0mk0t1v5bi0ULYamgxykuWwDI0Co
bGSW7ExseT1huc/zfy/xZih39m9YZDDRjZVm/GVrSFyge3ezsgwiQl0Tb+Za+TKh
oDcdTjY7swppaXGcImvAN7GU/gJTjiNyjC5DtvogqsKxASAcXXpI7wlgqUc6dxhp
dYTzYmM4f/voIiBklQX4mDmGNp5+Cl996/a+weFeVnVgfGEoJrx4vdC4saFcLS70
WlS/w/iJsQ7lyCdfIpKeBy7kuilmZ/ED3zBht3+BDs0WMXUFZwrXD/zvNt9i29w8
doFNZZbIKwtMyei95Mhm1eIEqvF/A4uZuV6PJ2iFTFMc8XmR+scHdP8O20tHEbiE
2zIwD3/WYuOe+UNsQyuvDJ53u2EuOyRvQGihJJ3HCrx+yADI9yINMIxsgaDx/eSW
z4fDzTqWI3h7b4S944XDLNubY0HgdkGnuLTFoi9URwF3eDLhwfvT0wFNT8CATLhq
TNjIieIAPOn/UdxiZ3t2bDVC1MX5/L4aEOwG/93pOjci3Dhk1YNcLRwH0oAvtK0l
jtt6gMbfXtnspfbpLjC5r1MBx5gHFRnfoqCU7ZAxjoeD9GF8nFFANoR9XFU5YRlY
gcqtUhTVQlUXOMSJCmMN0Ofc6pqJpAVdkS6UjvG8xxmV2J4Uzitn0haGK5gOeIKU
s5EXd+QTvh2rL2KQP+tpk6j/0T2yViKkcicZOhQzvVt4zZI3Z2oSLwEriVYBW8r1
HECba7oayzFH/IUPWWkVkeTprdTp9XPoXyCuO/7xcd1G42MkkBRgsx/0GtkcuFMt
L2H6o7Dz+BNuDdE0eXU+ATlw50kAMr9FpggQUEctJdOBUdLTZt+ob0No0F+mZlfD
3EG5tqn8m2FiYkmDXXcoH0zklQhPwnFv04u5LYhMRXFrV603Pa+6GexmogHZUmkk
D2XxEcBkIcUyTIQR7OZhg1SNnDiGwX8dbOb9hlIza4gKsQJWFOlZcvaDSH9xDnX6
Igc79/H95uVu+zOlyAOJxvEz1eo4LzXFYYceBpnGJleSFKAhXCqYZfpO0e5GOqMU
6HoPEHkuPNaFJuFzMlI66QRq4Umf3BX/eCpDwD9NwsI5Pg4qS8FlbQBKDtvECgLH
/7X2MDKJznotLWtUvSQNdrsHPDjoCLc5G6zs9rfIv7df0Xx2QS6s5ZAOhfZhU9Q1
vT2zHqqwEPmC3otjEl1uHOt07extJZSNtjVmN+FGg7P8AZua6l4xDKmMQ5V6BvOE
sZBOqsprU26Pte4WyBuxPRyJIhbBn4uI6k4Jxe7YabFBbYGoTryCjDTHVYRCTNgU
491knayVZ6gGZ2tVhTMbgfsqnxPV/uFiBkXhwqKXR59wUPqGe5zw/L/o9jbXuuln
70EaBuAAj49nG60rnWAMTvsraIUyfha+wYieot1Jw+Irrf7KqK1LErIXth8hnlTT
6Yo0ADb5aGbR2uBiFbBuUaKof4zY+RskCzkLIRYi+6Fcjj6hGpx1PM36f30JGUMR
ij2cpNa8SEZ+jABLs5OCiHO4UsWYtLM9CZhto06NLh0i4sE8hI2QYcn9CtMN0nt1
qfAiaKU6aXAwMwKmjNU5R00WfjLjiu0/msRb6F1dRTQr1tUGntlC93F1t3llSHKd
p8hlyPdvfcyF4Ioqw3ctHq9/hqOusx0bKu1Z0VSPALHq28ov/qjnerI8de4BugKx
ZO/2rKVQwW3d5y+zzAmswXv/Ql82n60YUi5PPF8wY4lfnIXx7eOQuOA3t+a+FDjJ
oFYb3/Y2WEt2rfi+6Q49HgPkqGVGr4KSHtSunVOgDwx62pAUndOxv/a1VHOFAupz
Kyu6nnkB++f/89oYRMJJ/eLJsD95i6Rr9VuGMR7jDcImj28N8FxgW+nDHqhMtnWO
gHg6vA6UG0LthfMvMHXbHVkwhGCCsxDHNhHnzaNtjUWOYyFj1WV23ANf5Fr897RM
bHelkbSXqN6R8ejDstvLBLzpVvwL+HzEYeNYhmh28VVO+YfHn4RdFYTuI1vE3RnM
iyOl4P4PURUcGJOxK360yWDvtT/aZqA/vUGLq+/nCP3KALnNYItVNwtiUTNC94y6
mWSsFW0h7kIJvlhRP08ldPaVzSrbWZIgTdvqBclIhTSDgZNODBZdoHEIWsWcXvIx
rKVyW3NSAZokdsvPH7mbXk5fdyhkLBodx72uFUxtgn4uF2JJ62I0XdSSnvSGAcDA
vedyfTRCwDQ/J6RrhbYh86bsi/Cu4ur/Ly4yoWAdCjTi/KJvg3KohYbSN3vpMJWL
O5eLlbWmq6dSRNmqUnyYCTAQt2qBV1x0MqyAkxRDBs0AZOlXK13LPSadFGXjmOLD
k+YFL3mHEHwmL7DIFBxv4j7vuFqVEoZPcjG9RVzhYNzSAyH/whWt2RIwRn7lOIMG
1+Ymz/tZNATBfng/1vBgbbcFdcjvIi8pbszrv9YLBqNgpdE9MEW0UdABUxjPopcQ
Xl4j8RzJ6+nmnWJvbRhnvrAQw5kNiZ/8ifVoi3B1FX205Z9g2/jj5ZPTjM7Madqt
Zbcbshps5Ec9El2nJVRkKDW2aMUgCYTPGSZ5TPY9IDFreJJZzBvZfrKApyxzijD3
Tin6IBGIz39JTT7dReVwKFgzLbMvcZNgnqxzinRSLE+REVPnN2uBNqyh2erZAbSw
M1jJNW4nreWVUcDafAfkR6aez6LOOrxwaVPBjO152aRXhfg6UqbemwuPjcCnk1Jy
jQbFdbjaN0J+mfJDFwMaZF27oxaxkZjUA9nHG3Px02evR9kr51+smdg2+OfrUPWr
7zP9Qoe7wYL5ld2Rk2HdCIt4kcmIW7LJH9oIVHmm7JkOj1eIxMKrR7McupL9WMn6
tXodeMD8L3aPW+5044AYOsEp+aZBbzqnRmNIDU58iS7PJGyRbNhjGixypMSrKQTx
W3wIUTCcIzCvl8aT+/1QNoCLrjz2CVWeB5RHByB2R7vvvhLOqW3ncqApCsyUDwpW
4Pm+yC5zMgKvoBLb8uO9lhFCrFZNJi5eMrl2bHNBynrMIzby9/FDeEVqbjyGFQRC
OLk562zQ6pctWm+QjYMPBYOlY6XqaEayWVYDK1WFJ53TuT/65po3l4VrAzm3R9dI
xh9iIoQuGxnzJidu7mYbvwVvUyOg/tsTAnXl5PhWGmz9aqwoMestrV85d3faqRdf
wQKkioYDVzKm2FlPY9KIoEt5XCLC1pgfQh1q8kasrvgi1MPaYSzhvUEQWXB6tCrg
3479HEbSMQKReMqgXh0Qsg9OEm0Dxx4iYlSUn10CkwvexbgZpx2OJw+0KJvYLlI0
m0DMB8SZmhnz9i5O7hs8/PcSxygCk6WAbd/sydqIvENofCvjUvAoxBZTVGg7p2xG
zaUiQZHv2WYL+iaZFcdK7V49Yv2QYyYCgCTdBbFsM9hgnq0aYT7jyt3UP4E5fClU
6tWpz2y6uJELak5PgXdB56a1YcSVssXxe4AzBlGhEDAD5ivM9OwYnziCstNjt6++
bTo4A7eIrUjUTw8fp6vm0aAOppV4fpu+YNWuckpBQTJjwI2V6tQFtqMRJJo4gEBb
rCFKTtUlQB/FYkeahjyq+8WPPxo13H8FJeNA95shG92Wb7jReQC9hWuL+4aySjOo
bpTKuarsi9BcxmrMWHkD/4roU1VPsQyo05xAD1h/ElszBZsYEo5Kp9kgFea02p/T
w8yvkfknq2X5zEBz3ofLRfH7fnNgBvgIdiYRixjUZLc4cto4LqJU6j8jNLxIVbjf
it5luV5WcOub+Y8FDZOh3N2r5i3o1GKaGk6Ssm3hzUX+ynTsXOGO6M0OBrkPpwRY
jpo2K2Q4VMY2XwbU2U/W9e9NK+Y89e2Wa1ay/cAN47DubZuA7ScRZm/uz2l6TKcj
+xcTkAjdrSsGaaD34uccxadjGfmEeA9rQS6beaEBrhLgCRGrea2hw4csGEx7li6P
pF5uoXoAKSkyTK+4xXGJaGp875y85HrJcl14E/3zeMFTL65W3qGhPIFCRwcj5gMP
vQf88zx6CT+lBTMJG4Rzxzs0lXrj+KgTECw8jckU5kOOHyr+shYNq+3wuK7a9MZH
rWXXr1pOBC1HKqPXX1cwY2OD0+hhhmyrYTCP1fHcLLLMyrQrY26bxN1zjtOGw2jv
JxPVWKcZq/g3L0/oOruA/x26EIjHEQRCTBDOoAjVPYLcjzqrlW059aBHdNUGI7st
lxRpY4ieyK8ypJyDCsXbfVN64rbmX8/AdmUsTNI1T5mcvtoEt56kd4J3AbTsM8Ln
6MlGeTh3roWKKYscHm86qT6XCZXPa+6kOAZasTeRVgGAKLGeCt72SgkJb4NuFoPN
0KcorBq74LME+pGbqmhqfXZznXJ9DjFPDkjaRC2wRAVXV1BXBrc+Xru1F/wRgfu5
NLc9VhoaUJL+MsHL/UEot1s43or+stzMxx7Bp9uAYQCZkj2Qv8YfQdMGQdZtPtEP
SPw+lNFLHry/jgwgcW0LeKVF81abjQKDfI6yHtGgTd7DPJBFFqTdnPIjM07e31Xk
gLdpUJphdHvoTCnIcesKH7oP2VwzFbUUTXaxQvrM8ckixM3bI44vUTUTy5RvjsX6
5ULL/q+P/Et316i6h9FLdkX9WJXZiRvqgeW02Zvx4SRnYWJoGSWMZ9r+7Wz+Asbx
u9I/pwjDwWRwF2d0nQEd0tJPCu6CyYI440zdiNolZHMMwQ48wnZpyk47LbtWKgAf
D0ydTQFor8PvjzlCVfS4cb548TwKV82nmwy8rrszf+u+KPF9XoWK+Uh3K9Wk/32H
rS0aclprAVr25xXenHYjyhhOuIF98GslU4ojgH8D4smTvls5UK0IeJudLmYazELH
TmgkGM7++8pnjiRtMj3DSuDEZVkreGfA6tbV9E94+uYEwzO2u2EgISMkgRKxllkr
qZ/+41u+518ufdRg8P8WN1mjAURdQ5KSMUamT3D0FgwtcYAgIpRnHxH1Nt/OZEbw
nzM3lYDCVGzfZRZR8TeduhxS3AW8Ylr8MPUQBfToYWjfRkMDuvxmpqG4Y3okkqle
p28toIl0JSOORtxYAW1sw4BrFkiJ8MOAIoQr7HUx9Y67fXxCi+T58iQGEHen5w4E
Zx4jTpObCSMH0BmaBrsSdSxLzInaEvFafeSLg+1bLydsY9EwaIaMwANluLjZaeU6
uexvnvH1GfgS5RhcDWQeRWr7O+SAJtRBPkLdQo4dr6m1j3XqbxMNFgOBwDoyZ+3o
gHyv8HOnAFacN40vfg3yXmkIAdt38SdRas0nXe0YuVLUJ8QCXZOr6HjRjfFlqAfS
JMOYJwoPFVyJzhL4K6Kb9OK1Akwi+aORmbncHBbP40l45yGjR4ngiy6DKDJjWy6g
20Nqo3LVzQhK2TzvoSCsBk0TYNL7tDuVPNMdmL641TNSEEhYxRR8cN8E5Rb+uGti
VRvrKcxWQxQh38BiylPuZQTtHHoB5TbStBTAAaHs0CACEWahI7wiNmGrEoOfLY7E
GBZUBqkgKcN04TJo2tZPYMv7glPtWK4eN2KfHpXSICAcCbnQma55NK223e3YZKwM
94JvYazkcUORrFvWfss2NoG8NPdfcwqJTNd+NIJNnrMVxJVxfl/X78pYxzXXWvKM
dgGFvkDd1UciHe7B5TFok4thx4uDGk5sQ3OzGoEQ4iTrFne6vSXaNxrM5TMnSjbA
S+7v1VUbmoGQsMa/2pXmEcW6KAWIFdH+LjRe54cId/Uqly1kX75o/1WdRL53BTR3
kxrbXtNs41+gKIzRX4OWk921xcn+PaMLDA1E6ZPZmjO2i/mKhUhdAAZBnlLLz+CK
/qKvk2xwqLxqOJvgj4wtGKZbIiTUtXYwDiXMt/I5g3tx1J5UVknq6deum9ay90ct
5DI138wt3a5NBN2x9/GX3DqoXnbAvd6Nid3Hsr5gBGw0Ij3k1CSjN9HgRBm1OCLs
bRoxiladY7E8riOAmERb/nHd5f8F81pKluJAH/n38zkmKmISD3zGhM0JvC51NhB8
MCB9qT4+o2FtzENSQbnstiOajrJSTJO5LAnazc3g+/ed3z5H7beNvRI9BJOEbIFk
CxGV5pF0URYHaehHPsHkkrlg4123MR3Z7sKTkpOm+j0zdQsMm3Yujoh+a+PhW/rM
KYoTahjAdnnZLl2iYx1UmqgPpPeetKfAc8DKv4bAwCUS0wkiE2QxaIVoJ7SG01mS
1uYoQ4PXdC0Lj2iudj5GfjDX5uBeVx7QuW0yj5g9z1Qy6j/p1jAg0DwqasAcA6hJ
uxvu+nkcUC9qNG4r3Pg+2akV/psciYijONgesEmdlQOH5LwraSbDOj6+FOmh0CST
Qgiek2jG8LL7jALiB/mrUNDJffjNhtFkIW9oYv/Hxp6PG6w1erz8OXMbQ/e/JLum
TJHxTkd8yB00NJsnRr4YPALTeDebewOD7RFS12CcjH80CLXtSwNk7DylSRAk+8Jb
hmcMOWA4mYI3FJGkpjdgRL2uPWN6Kn1qq0ZO9hxfiKN2V0rlkUxcs1/hjRNE2Vti
eSpKF98+Bd9g+Z/+F5rxV30nDnqjgMX1Oqoh+UdOLQOvu6o3ftVRYsURHLzTG8MX
kNemdtrCNUDqhovOiAR+RgbIRcOTS4BDC8mzjr0SuQJm5G0t7c5usaw41jvEUVVu
GeQj9tqCJ22560iNT3pDc2v0uaQusdbKjH1YMn+Q0Dzya/DfUVEQQqjEUq/QsRlj
4Plpx2HVsfLyNvSHMPmosL4gHg15SMMJt4epcKMWGMr7lG8ILy73Cbz9gTbDtMZt
Jb9oZqlcboyfcKHvA52nxNkfcMLkgjWQ5ZoMtZoUXbGqsJvKUz//Ooe3iSMsZCsu
JaXfH8pgsLxV7wAe1rIJr2ipZKiXN48jGGsS3s+/ESMAvBR/B97AGMVLV8w2wX13
QMZ8O1Defku5YtUkzGBYR+1c0R4k52XyjUqePvJS0tB4FcKwzgqwTa1zvB6QkdWJ
tyCRcLB7Y0ksTV/dOtr1Mb5FVpOj9NwZnvQjsf+nVRhrIpyCq3H3WsDq/zFk4TXa
MMM/TYxGdboVeNPUGSgi6gB1c7EhDWfi70ai1lBOMBkXqOM+pUY++u5gSfBbufmR
BNNt9A+r4TYVqaoLmXkidYapxKccjA4Thqk6/ghPLWwwowfPXl9GyN0Gyls400s/
SqaZuyGi0B+HTF55keHg/z+ypoJPESv70TMgvmtwW41s4LrH1xqv5v04KvutGabH
kDS2HLBobzgtp/h9fEGgZ97+57+pC6suB9GzPoql2WC9m8uAA69IvOmE4PJtuxgW
dGg/Gg/c2zLFK41Bcu2/iQqK7Vsz1aTqnzIiilvMi43GFxwd/UofRasP2RlKFXvb
5RnL7JpUZxn7y5y6ykKRLKGoWhZiviSuqk6ai8gbZq7594P2uc7K+TvDXXtwMKYv
8apmNbNHUitW/wOM9sdWB/uSYjxsTRdGJffr+Tn/KuA9HhGYx3IL7khQg5B6AI+l
8xevszqiZjjOoLfZ66AkeE+O4+k5h9ytww6PqYeQmcJSeobhanRkhQ2a4dwQvwvl
JAXvmV6c+5pAYABTam4aMdHiU8c64q3Yjzg5v1+WMjbxZpewEFONbn8w0dwQGL/r
IIs4L5e5RpZS1a0tBNUqrk9t8k/daumtIdKw+KV9oxq6wxazSKLDw1uRod8I2Zoh
2mTH8uPZavcT5aOA2FEzuZFkG9/9S+d0tp7cSarM6wn9A2eMLQTDojzMZkkKufkq
Ag15GXnTYnt63GZfNDEEc4Vlj6xz/jDbTs6tx1VbscMdN9XIEliuuNTKEuGxWza1
oD56vT3hyzXiB/D2HSPgiYrVMjg9dct0n25KrfftvG2azLWfyA7Qh6jj9GgZ8yZB
lQ1EfuyBz05TWC7EF/GSgrY5iAlh4YZilDViDCYXZDV+UVUDe2uTFe0kUOmTfk4H
oVNS0t6Fri8iWgVjVKiTf0N4JlYarriktXa4anSO6dNcorm/5JvZWLgo6+73sRdB
/qhcOcOtt3uwiMgoxm+wIREPvrjK25XpKqxB+Otz73bzU7II7DroLpvAKoxVZ1sd
RSTKNWNLef5yBEF3qT6FIk5gqDM1wFmSNNdNoan7dZIX7sFMgZhFWvos5wDHHL6a
As3sd9Z2wd+RgDO1eHZgKF4fWxBpPkBH1AFOUUJwbeJmulb82UyndNI5njWNSTUs
zsDc4omy7Ei7rZjXxew/g92S0aJfKViAjrxvTYgZkgjoZXUZ+8M7obkGN86GKdzi
uruiBilGpHTCQTdgkf2+6K+2M5KfhZU+WiY/45dJjhD0VLya/8Gc/u2rU4NafkyI
kA8vXYgO5vEuZKVjQijJ5HUK9QCdXfU4BYAQzgUqWxTdDo8KLwfe489+DwYgzNH0
639m3sv4w7/ShjXu7kv05Qo0Qq92VD8YGfVl9vcdlK36psWiV5o7tC/Y8ZE70s0Y
LV1kkKcE/9LNjpOJAFq1tdqqkmZYWdFaOrj4HBB26JNVswLqmWbb7BpCxezejZLZ
dDSBzc4jVbkhsgUHdOU1p++pAeUaJZCnWAgjxyuvXKpBBBY4/WVGer86Jgfj6awv
8BUkwikYg/S6l+AKH4A7DJN0gH4fCdPr2xZMrS67Fa1QvmqU9DINWZuLqVe57ffY
HrmB8IOARxXmYNZfDIURuLkeuaj4NxCkKgdXweq4MuWkzFulJCQYNEKZSLvbjOck
+gO2+HUWa1QeZCXLjsnSk+5bWYk5S7fu/Xq4y4BI1zqpkuK91Wb6Vt7obbXe1KXV
JqyUlJTDfOfCcnL9KazbUSBwwTMTT+chqnTTgUZwzS8Gu7dpulj8zWxwmLHIhJ+a
HpJP7sZosSjuMAYvBB0BRlesULoRmA4fv1jmxjP/mmpZqUbzd/U9eM2vumA3XaO/
8QbifXvMn+y4N702fkqcX7/s0jWZyU/bFZNR6V4+rnlZNRjVY68dC2gUjiFSEErK
OsBM8n8B2cSsQ69uDlbnzYLKcHqdrhKL93kUyD2YB/6qcVV89Fe3NN3ljBekvojm
RWi4hwrJie3xIIgyr2Z9kxf1y3hi3B6GkzmrODqQ4Ags6g+vjrKmhXaeqHvVbYz6
b6v+MMKV/rGM6OPrWlB4KEvvuUxKLHYMoaPx1j4ZiyN7bkM9k3o/qcWJ+Wm4xbBx
lpeyEdWbgNMV2DvCmIHRHc8KfCxD9V6o4VCmMMVMpiHfCVkWrXcYOnzDyBBI5wrX
ApoHGxw1z/5akExx8mRuY2NjFCoDps3XjZD7JJ2sYnTZcOirdHKF1OrPps6KBTtt
4GvxI3NNjfbmCHyqxNUatqERhimfajlCNtIzdLkLaGgvhIRi6MG06cvbr+5LP8BS
B4WFxLJ4y0qjrJbur16TGWqRxBjxpJzWS8GwfzOZfDvr3mGBdf0JKWttPB0xP7pI
igkuzR0d3C02+BP8MfVX63bLrtWeUWKNJB1FFRe2MKje8cF7XenczvM5JvmI9e7r
KLBy1cneWOI0ocK2RYLgB29L/UQErsY2y5D1wHB1b7485wMhydF6QDFTGlYz2d7P
onlYZH/4lxcHAT0juzO55QY1HgomIozxzL7c2O/6TWFslJOAjnnYMSUPu9ESloal
U27ZP8hZEvPA3mw7Bak6+l4RHB8OsyinzC5hgf9TbHyASVD243J+OEHTHyd6VHaL
GPLnXBHRpUKrj20nMzDCIpvq4UI7sYcVJ4ILjs01Sx0qUX8b2CbhJwZCA/tFQ33A
Fm8mBCSQ2mamEXQgzP0agSt+n0x8hh8fy7hdcXpyNT30cCBtfZEeoUqaRLaE5BXf
CJnNjWkO4cFAUl+buYTEcmHXVuhmugF3diHdawfVnGX1XxejnRg4GQrzOqvgT2l6
fkTD5zQwPPLyg8v6vjRdbMbzbHco33xXGw+ep8yh8Xy3zzIsgC2qhSMsbR9PDCLn
2qYd+ZmAuSUyaah8DHsWElot+0LtgIkTDbIGOzMHc9eIlJK/LfG8vO+RAxq0u3EZ
2aq5fxy3/yPB7dCcVGC5t2zrCpIc10eqg34QiO71v2ARpetQPntuGv+OCU9n5COs
0fBOuxZ5H6yyMDHhyHTM/EgQFpk6Gu4/fVIGMVMWNvaL6jBhfzAgAtS0Cuu+uiB+
qflaQELbCfb7az8Fh6qDIX5tjRSo3G5goU2dWeLzXUmiBKsl2ZPeZiqHXR7Cp1CK
jbVDiCbkZWNTJjIvgWTLDaITmdgL3Dk4J0Ex0XdYFyhXCIza4nHBMNBqwpDgp40R
+cxtJ2CWLkfc5XEwLx68vafuGuOWOqPxbSbsKKJ3cc8UJW0PFRklhFiOcMPKfqKC
exkUQ0NoLLdrhnJbvhGZR+HQgw/gSOrFGSwKVVTzytgslRf47r3wza81MQ7ctmL3
tDchMqTdC0ksehEAg6rbdrdRtZuYxOROw0FNaLryyCvM6E3UDWyv/ZGjjb+ezhdD
2q5BoTpBBobC1/ddVPjo12vNdzYUoJTkAYXLdAut6bP1HbUBnZnt6ieHXEvkArtH
wGBRkuXv9miQvOUH3h84HGyvjXXKsgZJZLqOizwBWN9yoEhx4frsWleFKbe8PsUi
VJxGW70Z0QZjHTSgUmV7K63EKbp5SCuH9njdYjbFuG514GYkccaMikcJas3z61iQ
DD6bAH5ytQbAdosv/jVm1z3j2Vs4GATB4h1OtLnYGvzAWozOUXjwizXlNPhizcij
HQxQItcLfjhA9nxdtLRSbIrBKGuQ5MeYYG+n6O3YAHB9ABFQYWgp6yG0s97RQ4AW
tlFjYYcdvQygblKNZ5nAs8zuNVVcYlr6ML1qZvBS3/fww5iO5aF8c6UzY0eY9RHz
eCb0hx1XA6bzd81dnRYOgxnkhODojAW+HX3R8k4hl0n4KfwrzHml1AQi/rzzMA1l
mNu97elPO880LKPXhR9MQC9rIalYhZ7rNWh7G+Y6jBiwdj3rgjVA8KxrYVHEa/ss
KYppRjXgv+aSvwZfeGYq+/bjTk2RPm7k6pbnWJHUUR/Bfxm8Qkky0/Fp0qEEp8z8
n5RC3H0XHl7asy9IeCmBppW9N5t+HtTEfed1bO9+TKP7CyVxEI/dv3Ayq7R6tuF3
LDg6Qrd5EvsdfivAfhkE8rD6GnVKfimc0VYS1nBxvhxE1C3maGIA5jnA+7Y085sn
Fb+ckUbCW1/qJRljNZDXFjhfyV9JjBJ79pIYMi6LXYXfeThqPGpm3IBsnRye4FdY
+SqtItzI+XaxtfFH+LdG5nRoopL0vR2E3ds7XWp/46MOj+ImMdBs0o0lRuYo/5nK
ja1oB2HZ/Pcx4VpylMxw06ptKlCXOLr5D/H0S/nEZ7N26ErWYXqkrypRdra1QkuO
IR/EgN3kB3wMLXTArzRLx2eRXES5x3TenDqynnMhdrbnpn4xN+jV1swTyc91JXII
Kc3FR1v9WtBeEFFnZyiNcRXW6uoFXKMe3lgbsvrdGyMAih6O4URKbAkEg4SlEqin
+RbZ+s7jzESG3extXBWHiVcvdywrL2G/Mb1r8m3WOuKmWcfT0n8iHf30cGFRhRZv
CccDGylw2WpYew43RskeHA+zWIov14XYYI4ON91Vz0b9T5OFzkbk7AnJBo6ysotX
W9rCx6NoijXsjiTJGxtoeqQOHUdHl13F3V6jen0N8kN/WwrsN37Z7tp4E3q0nDN0
ml34Z1cE3LiiF5o/TVzuoTNeYsxmfoR7yBlVUxe7UBTkAMBlQPQSGu8n/v9yreKq
pnhBfrGYHT/SuzIev4UO7TMrWQx7Tt1U9a06UY9CM0z0n32/JZsEVzRulYRi924L
/G9cAXqOYgIdV47bYDxeHrKvFhcuqusj638Z5oiLLO/gqN3YR/pBMqYdMd+NQBQA
moSpcaLAbCJlhlvPMMssREUqfPd80G55tsnLhcos1ilVEnha5w4qjjjR8Sbas9+R
3FBoSmryCjVt9HnSt3dbvRK2MQ+2+Qj787oh0IRDVM6YQdgB1v5gVVmEFf1qkMNb
JTXbrKpmxX70Ih3QtRDpbqao85cHE1UwvKIha9nePVlEDwfIsrwOj1qhwtKsXgps
rZIK8Z0OWTcXc5W0Ojtx6M0L5g3g7W1qxBLy5N8QLOR2p0Jy++S2z9T7h64WjCDJ
D5rYxDeS/wCfH4vz9fvcjsUgMC/7I5hlh4MgqHbHCOhsECqNRXaOc5DOB3Rf2+ip
Pr1Z+i0JlngO+WiUgtCsv3C27wHxVP6NMXQXC7TbRx7GPei+ZfOTJb2lAuLe5vNy
P1N9WVqCZ2lvblv3P1sEX3g27BXGq7gpIqCTeDfR3oWE3u/Y2jVXUN1VyNwendUc
+KO+6OYOpB0hAbZWwzZ28X6jn/UCqsnGG6/LZXfq/IgxGcKa7A0pxY7O6pxdcxiV
yubD7moTSaI2bJKYlQaVazWT/Fp68fIrcIZrCGLFWu+7fWA2ZZZpNSL9Ck62hRRv
6MdD3+4TaCXcLFwQsZDCPAupNrpM7w1BgbncluOBHWMhTd6XTsWL+t5vBCX88edg
fmeOhP4O+sT6138bUYJY9qLjfXV+IyYf2v/I5xNeDH6gXu3ZxtASIjz1dgdqPM4W
iafhczGrIiqxXNVfU/jmWuKxv5SJHbxnAn/K4wNYgcubqmm1clS/WTgFyuNoD+Cn
lEBlxh+fcFWpaEH2ySOe/AbcFSdDVSjPNGLUtUTlMedrl23pZY3XqWiahGa1a9yG
isZCTFPIBEUKfkFQGVpk8PdOEXge5aQGNZtJjv22K8QpFHh4Wo8HWkjd1F4x7NCJ
COpqDlE0kEhy2NzWSBVmu+ezL6dr5Tv0XreVddYUxU5pklCIC+9fInQfp+R4tBvN
s41OReJFaB69WWCnCvhqXd1OZ8G7MoFnvNjWxQJyEszrwRZ+phcWTLiDeg6ZUdr9
ouucWfQMxNCU/aWRKpUapRM+TmVXYIJzgZ/A0VuFLn2lGamxhl0kSiXqJzPpn36f
4bQ1nAq0bb9tKvI9vk3rFL8Bq+XkKJ1wmICO6xQ8o6mTSVyobGJCmD+Fe4gSL51L
1xx9fCy97G967LAI0SVfP/WfB3HWOCdFafdyLjRlKR2U0iZGy9TxxRzZL3r8TiO9
2k3QZ+JHE6YHQQV8vsbAfLI+ZUbe8ckFVTQwQGCAF6saQtWS2AhyCGVFQ6mge8oe
5TAkCK+bjXgf+Di0aQxXRAbxUSm/Gx6zxYIehoOpbdaGZ4hqRLFmQmr6JVBqDLWk
dnhcmCr4oNrdLO88uZ/mErpjWAiIEwB+RivU2HnFWqz8pD2hYn3hnKyeciaG7uVO
3BTHBs9DvBZ/FvAthdsTDcNvC71EecpJyYIrLQ/vfPFrEk+ZvqOV1wpOBgC74NT4
T985bqHIR7lxUQJpoa8YbAPJN2Ws+2/HQxSVLE4PjPGhO060YSqtw/O/VoMuq3Vz
7SW5ur7GuKVn7Uf3R1XOoPWpgbKWu3pLhnn2JZb7lTnW4gN3QwzCLZLE9DSvZhWb
WUXoqxazdABf+JU//sgsTxrwgdCwjh9hZtE5i7q89HFiS17FmhNs2+g601t4kfoo
+zVMZQY1yozwQHieXBOVE707ozZBLa9c7KcpfEXy/Of5/VxzErpUfzlQvFzW045l
EF++uwvHR7pRPkCLrwJODRnho/pGmj1Rs1VawSRcYPeBTveaF34sAqVBneNr3z8q
/NwkwRHYhBj3ngMqcAmwnOPS4cMzJMqKW8lfP39bqOYt5qWPo8nGdbLhOSGPapez
Hm+TpRyUi0zp6HQ0QacO0N9eI28/VNVClSeN580HkvPWV+Z0IMb544HN0AjQkeeM
W0+znM1e5OoW1Ts27M8TBNzvZR1hFjnEBVHkZL0+0F8w+bHOgmWgLsYFS3U26Nqa
thyN0tXwCs3XzHWvKMrJijx5XuNdmv9bkMXsCAvzvyyN2IZgNsv9KcE2aTXE5RI/
Qu3wJf4te7OBfQDHDTVeIiU1K5izhlPrK3q1jl0YkO2hG+3gG/qgYhVXjdqdEWbo
JENrOGEu9E3ACB8yA2BtrBTdDekHdGfJ1IL48zmFCiGdS5NOPoZpe+QqNryH4+Gr
Wbebf5V6V3d8JiraGmQWeiLWhdG3Xcfo+mBgp4Wceffj4gQCXdB+LOK/mxzFvSbL
qQmXu8n/04NY45haDoJ/JnaORnwJyARXgBfoiyEOSd//VimEEppQ/yuxOwInOriH
gckcYYz1hYoJYJASk493Iq84GWBEBZyL9Dlyc3f0BwGQ8+25y2IchXQJ9lismtHx
fGTLLaqwrPwsWq7+IKh7AL0vjYQJmKPkvjg5NiFDHY1CqF8uacwIn/9egP+U59ee
dHRzgTYgWnX5wJQJ2B/25jhWhoo692LnLH8j79LkQ2Re0+0u0HMlUFAMvJBZ8JsN
6mdP+s6TDnQkBjaDQceKqa6SXWqN19bOmRntsq5vBw6Keau/d4/zWxZ5OU9Ilk1c
abmP+uoc0sLgksI6RpqD9DaV2crvcDaaLQOJBSVBkkCVl1Sfh4U1xVRF5CvQRDKY
cVS/7QcT+45fAdjTsZTs77v2CNGGg8WTYq5aN8OG0LG3zAZBhm/olH7WyEPeWD7/
vN1xHnW6qZ/h9bBstLgRK7Onpe9geJFR/RR4RgecNxXyjSVpZUStBWtcSji/W6Go
qQWXLXiqkuV43mdz95bXt4An8m1Zd4kcXh9GrdYdavBpigSBfxfYiREkT12Wpj1i
qaMKNVvah6C0/4q8YdGgjYkF1DVARpn/nlOgQWqirRc4QzvWT8nM1JoGB+ll+1/Q
wxYtV1d+lFnDddZMMsoItrYFnAUf+SySJd89/Mzw9Ixde2A7pvS2wQXTmQjxZq88
X2t+Xr4fzdt+OtwCPnJiQ9lpifr+3n3H66CaqEM1s6fxxgghSkyl7h8sub5hczb+
9zG11GJaosRvRfi8znwOalnI7pkvZLV8pyxGkULqgNYOQG+1AopAdfavaqFgNAA4
7NB4dgiygMiKas3ALEo5dn+H7YMHARIEPQ5fzigVDXn9chvipVC29VoUHtihoBmA
PbKgdsibZsnEM4a4B8tcUtVg84wcFQxOnUJyCePnU2ZlrlZfJo0tDkmkiFug9ury
vaQopy6RZxGH3S0cqS7uD4GUkM/sy2mAz6iVm3cABd81GDsdsZ+2o+wzz5vibKTq
ne9QGODTQyOU4SdhU4DoWdnMDdtkKN1U+elbcz2utg81mRGLDsEyFDgcY3SZ+0K9
y9MYGP48BRXrOLJYVVyRUzNA+qHSrQTwiYkV6XUkqoRJlcjYiFgjrtHZwsxNTaLQ
f7EDRsjCidLviSU0Dt160bYG8k77SjUD2dgD8JGx2MAx/SXJGWYpDavG4NCLRVo9
B667u5eBlG+Rcqundeq71YOehJGFzB5EkataOOByMXdHmAmLMVsXHiUdvc5iaIB2
egju+olQfyNT0+YTq/9QF1eFcmhnPvDz45kM7pYVvGrK6R/WC3pAYN7LbX2vVyOT
dxTF9QYXvFChlMXvJmOQaYSqVVdf/0PHKy7cImjfaPaMAhfTN3Q86ZOjSjAuvObr
LjObBSVGT9O3uevf8Ybd2/dHwi7cP7UCMGsQ25MHLlgHyVmZ3nnN4b4RKzrSh0AD
s1kcgQouCMHtQEYwgun9PkHdvzftAkfvwudth7BlfPYwBGdQO+92nkKm687+Yenc
0KhZ1N9OJOmr3LqJXHakQHtU30/yrswzUk3L8cLIp+wukTWG9IMCE3PcubFjoi3D
O01Wb490K8lVhYlcpnj4TD5ioVbj1kaAgzS2JIUKBWbVyi9e5dXubsAvZwqOMzwH
xenpoxE/yFIYMlGBmSfZYsymj1UAt2pxMoDGc4vH2u3qSE1C0tc34SIrKtro0Sse
LPfqbAP27wwnPHD+X4ic+ubxlOOS2kSXATzR/dpj7DPMR4l/eNKzHuVi2U5WDQZJ
5ByqtjILmHhsxZkfNkHocTHoCut2GC5ylMOuEqdVdzwvB12UwlL8msw/k4TXiOaw
NjSGAmwQDti3mL7viSaU0GEAQCIoCrCpxmkpGaYdpbT9ZuAMr7Es4BrFnx1M6sTW
+PCLSOTYKxCUjqLEBstrp1uJn/g/nDrnUqJPrIdEzHv1Us2NaDbE54cr3YNpXToM
/b94etLiC992jt8rmES//mJ3tbdfLJAKXY6/VkJQOS766XcmYOuKWdtEpv8RdK/C
sEWaltve8ws2TBVR7vFN49yUZeh32YDs4K0x0LlPfRHW3l7vKDzC8GXs5EZJDWjm
huoQBnXiF8nxzE3zJIHC03tT8Gf1SouEzvpGxT0I2C0eiqXpljj4qPlJSlSrmKnd
NdO9Z06j3XK+aU60lgLrNX/8mSau7rDSg/tR6D/zLvmnUpZSuMeNK7P/VW4wNd7/
HgU39I2KHO8ubmK4MfKavTBtcncYGRyyGXgzJ5AbhMEN6mqSopj86fXTAuXtqM9t
vWpawZ5zgUSIhVfzNdCFy3wEwsBAHMdC9NZzhORknk8neAJd0f0PnMLxLGyNmw6j
t9UgrLyKmLzS3y8L3acQHG8s4TUv2n4q/8NXxiZcklIjIEBgee8s8QOsDHCndb0P
B1FXdjW2MGols1UZt9QgQ9JiRwIOUzyEmztLszcGcNe4usYjBu3IhzF0Is7NT4z/
iz8Ha7nNnhJ4Gnt0HETTK+NOCkfLmhUmXG66zJZulNSwoDjXljB7zLWiDKtwgraF
ePLzfYNdwdLFe9pgMKrIuWkjnkYVGXzh6lvaXbLpBtg5kz6DnTno4v6dpC/v6oLO
4Xi+iK7NTFEqdlnnvAwlArLOGQYGMUK9HzW4X2k0V5VytZfbU6dnKh8WzVcUDznL
f0p6VtZJN8yRPZnP9KYbAuyOfiIM16bApP9MtavfCcp85ONCTQLHG9+ocEjeK+Qv
HfSNGWtdE2Wogfo+fUz4D3+H36nVa49nCXj1DI1zuYOB1uUIeRB8bV8DmWDNso1l
nFJAczR0HlJbE5MUyE3fxaC5bqCJjZs2xHzKJlZT9PAqXIoNdwViHaxcAzmApf8+
TFe/qqWUVXImKdFJtHJrwN5x1bAcc+RzO6/2jo+ZY1g0n8OtvthzEjkHzE2zRfRw
/9yVbHkq8q20q71LYLnOAxmtHU+xqztkfDJcxgdjeV0cXkoCpdyThGiwUKM1jdFk
l/Ri83qqDdNkuyUkO9ybcaAZhVWOqXgBsU26O3x34NnbaXvdjmsmwOu/LFJ9CSxv
X/+AVdaDSHmVewmXAMVMRAFAEdCHlBNx1AoQqP9xAU5J5Gd6OLjy1zubFE5ZRIcl
+DvcKo2hZiN1zaVkAA5+VteT6X7quwBe2lvwPVu7g9+lWADSPmxk5DQdcyN9qvon
byB8B9qvWg4OCciTHVP024MIs+TzGfLpYTVRo5lPtkQ6bZzn2TrHtsaI4YJ5gvTC
lPk/ambxUKKRUVIypDfgEWwJzViGols3G0ATRLJZNUTJYGm6K+FfPFtJSL3id6V9
gcLTCLi3LuypVcrjN9qqt1RAlEe2AYc1QZ/ziFKMaCmQ/xuEqhF54lSJ+9M5yx3w
calePhwwnUOvcCqxb4BGlrMna5FcqiP8lcxRQDq/wilWqKrn6g9nVqcJMSK8iLRx
NXc9qO55kw4uZqlva+jb/Bj7B86gids6UekUwZcUj7IYol14rj0+0tG2A9y/kSX5
9hXruUzTe06jljb3XczsdPNfrdPGvBe25OirNFv+FLqhEu72aRkwOYh1hKBraEsK
gr9jPjwtIy0qmcdRKAJv2gSrfB5uEnD7a07je/KBDL4dTrwQR3JslzAtgQd8oTzN
gfHW0pFOSDjYlnDvuItsZxpAQ/0TRAQIGljeXo1VndPee0DwT38bF30jHVxawuvf
J/umq4BnE77MngHwP1EPpfVnsVRe2ZDeCiUuTVvNYz6RYgxH5qEMCTgivwzDNTC7
QNwq00JQu5sl/csBamSYhjgsQ8IF786AUY1T5QOpxhsj7PCcUcJTvD1udg3Q3hcM
FZesreD7aW256NySnrFO3XZSsgDwU6OnbiWp9IhbQILSR0Xj2yRY1zltgKA25lqP
1WPD9JoAm5X+1yBLW5knQE/n5xaaX8vgv2WGRSKLbn9+7UtdgeUhIezLsTwJqJ3e
dV2q1/6vGpbCKZ+pO+kDwWACsKucR1bhU53GHzTKYM7rZEGFXxtu4VVnQg2A9TaO
xS5Nt6YYC4LcGQXn9orKkh9vcC8h+eIjgiAnFajf2ZhWd0UhWQ5RpnZkMf0lqWOM
ohmftZQUkrwcrD+H0XKJ7pesBgcanhLfFq0e2to30KVuAn8ErYKhZzQ9MzMUPaBP
730BYm02/vmPU3YMAir3L1ptsSVS1vkBHFw+wC0U2ZoJYj/smKdx6pnf8XEM1kyN
ywvBKSggqNr7bSRvBIPaLKhegQ9xttSNKBDX1slVqzaNWi4/fu/+xfWYsJVphIpB
KWB6U+D9xuj1oxrFTWEKwuKAPQ1IvQYC9gw04sk3u27oUfAyzdt9d3raTQyYMy8f
i+Qa87ywR6yPSgyjbg0QfehfsZTl9Tz8z49/4sc/wMxPHKimpCypic0F7ucRDUqW
ntKFlSzGsGqYGHDKjB/cg9zjM8J4Wk2CdCe4lA1m/9NmZgstLcVqnIwgHeYHehcG
OVv494dLi4u0Pkv1T8OtwVZPbkpvGZMlrYOwtIFQD5VOlrztVFwkEp0/sBf6P4Ly
MGAUCo0SK6kdrPmESkwFO2SIWAmM6TjpHDRZ3BngiyP8i+lbwB13XdEvd8vddlhA
bMoxFy84ZXN4Hd/iCFf/+Q6AaHjdlcyy2yrO5xNINUcYm4BVkvQ1nnZS87BjHzja
Aarlw5ywa4baXcwHIU++9WdGNtns2HxDERFNMIchLP86G1Iu179cREiHKeAKVKJu
Ct2dY33BTiA4UEUimhG5ChLT4azFNoss5f6pOD83WuUFGQV2DfRxex+xt7mgWNBD
kg5qLjeR3judVKMtadnO8TP8+BgL9ZwGRLt6LAhbGiHwuz1dl5QpPpVgMwBTs21K
OuN1/+h0Ye5BdAA68SsqKarxzNsJ8w70z4pO0MA6Uw4vd3js5vaBFTAeLfnGtM2a
wuXSAYRzE9g1xt/IyUb44KuxQSjRXNz4avlSo+HFpNcevEAm+Y0bGSQXX8mqTVes
aiv9jn4DsAwBPoox/FoJibS0VnxINq7u39Qo+FZnv7+XUxmqNOGxsorEueS/0dnA
SrR/zQlxNSd7Nx0p/QjkGEq4wuXjjkitGEt/Xfm/U16IappooJrV+VpDDSB2DDjG
oRjiGZKwrriBpZuK+Gp5rqTqXATC0bG6SiBwdeVZAxzO3neiEikXD3oXbry34dPG
+QptA/820ti8iKjvClo5Tbn1QMVWcTC2amL1PQyz06jCcmnn4qPy02HqwzHUXj4i
OZ9rJ11dk7kx/o5P7EAROJyZPF8Gykmwmq1VJnDGZig1sYoxIePEhd8+T2Qd4Ci1
mkDR2S5f1BX1QZCw/6BD9L9fKSYGWQ1aZF6qX6e2L2IJ+1gIXU35XA7lramyaDv8
Uo971sbxgn9xymWTbMU32jWOMKzLkRm7ZdqIyrirwT9PwlxEceP5HWfQlf1rVuTA
WR/EJ/jL0MEjShjzt076HSlVnX3p7EPcN9J3QFS3NkbJCvwdZMqEp5mLKUmAaYw9
k/CrVLSTdvq6P55DUaiigIYszhRsA8YsimHYFdEz3hQz0Er5NVTexIAYoNBB8BDI
zySu4UyfD7wYkheA8O1qYz4SdfKWYyXAY1oWfrpXCnUzfx48pLl88UJOfeanOIn0
ZHHx7bpOz+yt/h4+8IJwpaJipjtNQxgdhBOr7/MJAopZ7MI6OzmmvBqzcEfvcDoi
e7u1AVBOeRDiTDe+KgTAm1Jjrw10uFn02SoF/VU8dWGrlATalcadJLT2DxBRAFiI
FRNNPsHUwhnh2D+39WyQh0QxL4uxUTRTqd+vFtzvaU3xIid7gIAQqReWP3uCyj3d
eF2S5DMaAr+pEUx++2DkGn9ctu/Rw7uOlh8q25EiL5lmYglIZ5VnA+GPjApwvekq
8ByYP1GyXWp033QD+b2x1P2QMfZXTRztc3DjOJAUVlhT/qgi9HTneh7Y6zSg6okv
JTW9f6rTA5Qsc7qm41Ec0PffPqPakV+Lx52ghugh3rJnlym5fZ7C6hKm85aW28lP
sGURFcw/WO6mmeYMI9EQaV4KLJc9Kmsh/fmreaeBVgge+OVed9OHGOY30krWNPGQ
y170WdE/FcZ8ZgMJVKL3wc/vqGTeJR2ReJy0G7PtGjvXRvVX67t7X6KNfnl2KLOF
dgsAG/SwBrojUbZSQQvSYSxctEvMjmbVMCZ8BRzZ0x68dCbBob1I7ydnv1EC/D27
go1vyKWT3yl7IroxdPugQ2G2egMs3SizbbdtJknIh3/w0YAqzfQJO1wZOAVZ0Et2
itvsqYk0IVwfxAB33pNTQa/fH8gNc/k+or91ew2pMv1raPtnr5SFm1NLYZPp/PzE
MwUdgaBmpaaYwl7J5h8mmYWIioHvd7ooNV0FrDrIK/pjhjul/1sIcWFprWwFLcXc
KEZ3rs8qULp8iEs0ZlR1DazrFPjDhDKBj6sX1i6mAhthHw6WedRpKc09smRXyUnN
t/VfIdWQpq/7oVlzqcer5SulXBbf1L7ziqAxuqP5JxJYc7+/oGoXQDKjziVVF59l
FWZUbed3zv5Q+Faq6PdxIb9J++GNDD5zKgznSZTn4MbzlclZ3zEDdUL62wKrZ5yc
HaAlokOEXU6BAZ9bT+E7nBG4q5m+AZWSz5LSsbajNM7mk2uEs5ittl93kmoLktnk
4tv2Ksy9zWECTK5QQSF+WH2gDQzanr6AGAk3ocOB6/ULk7AxVhYqSaXvlHTi88y0
zB5r8cyU5HjiZo7ni6lcFHWIKzwc0tICQusZxv3rtbG9OXreD9Oe8xeRqYaqQqCV
L7J/LGFPeKiws+maLD3Wvog9dRDtgo8ab21A9hDJXnD5jXZjUH3KWDv8r+Q+z6RN
NZD9zxY5zGSHIAlpPyDgUSmnmqMhlL4MqMpd0ouVMjAoJKTcsbY5OosW2Cc7Pl3/
fIGeMvnRz/6RKg1YSZkS/yneOYS6PY6BSTxswMkscNy2iwHnANrMVDVvIiclzx4v
30uZKsz3OQiqoniYANhbSnSF7xt5f1tqxnZpGs1eKLsEFt0FMN3xf+3WK8dBYIy2
tSQPV2E6Ee/QoPtakWElJE2IshhOie3sRaoameIsFrcWWIwJbf/jHqjA+Dx0aJwf
6+FyiKhGK0Obc/NVZhzuvCukksmeRTejNIn9Q1DSfI2Tzy8+gBW20BMHfVBQqpg2
8rzMxM8hcHg0u0iMzLQ2sxNe3ZmgQza4jGQYiutTeT6YIaGf8hjg8PHxdYyY5juJ
324IOzlm79tNBlVI+KsQuikPi/bWmKJ/S/5bk0qnO9yCoAw1bc7CP9sOvxANPDWv
FbtSO9Zi8thnvXrezw1qNzYD0XIAHEqAY9THiMTFHY2aP2O3zzP0LsGaExmLeBqf
JQYnb8FcOvzNCTUBXV/HC0PR8TqFXsR4RaEAaOmRLi8fzqhm4OY3oTo8IplPa18L
wDjEWiQyJI9LBqD7NkdAUaJva686G905YIxVVcD8o1qOj0T0GJnZjXnNKCPpWgZ7
z8qLCnmuXAHLgC9cp7eFrsbFZ8lzhrLqxApScmnxzeAv2JKIvtnuUIWiI+N93vhO
IEJV+WiVgcgh0eOrDnEDN3IWqSTr9aXt2ka5514adCqOrqiFkuVOrsqhl8kdXtdW
rRrEnzBxwPo4YGc/ft5ytECQVWPQ81yu0Mbly0016YTeMOvIvbSEyqz8n7pSFnCr
akrKptW5Vrqbh2Gjefv44rgd6z1QY7S17+NrQ8QheUAnDTuJZQIcpCpJ9YNgA/WU
eeKyCFSYcYhwNBwZuOET0CquXQaatUmdC7lNRIKHsouCbpRxrzjC8quIZead1j7k
U1puax0wivQA1Ex3Wnb41e1X8e7RV5OFvrfvwvNykXPPdIG7Bkm4xbSJF+bz6V/7
8v83mkYCMQFDAN5jMs/RGfM6Lju+Sq1ta2uFvl4nKFYLNqADw1F8ly3jx3vGfcHk
+GQw9LWt5A5vUBVnJQBLY1Oud4Bdc7g+69xliR+NmZkHgyC67Zf6C1eRzO7rBBi4
RzGq1mZ+U7cXYDVqajvWDApFZQkio9ucLy/W5dDiWogKP5Sac8Ahehh2iaGVEeZe
8bYfDjXn0NeVXeWHU+92q99OtaRZk48qSk6uV1FylZNC7xlOtG1V0qtjojdVankQ
+HK2RNV1BFLtsYN2tmHit57p3SnuofceuV3d5tE2l2hfBjMxJWzeRVovZpYrPEo0
wvtbLCAOq3RhaV5Cz3+PppBRQi/KCk/cL8OsZtF9krJ52wDm62xyogIg5FQFfDYu
knJovBNLEW5RF18bGB7xjJcA1+6S9fwa1zf++RuXzDqm10pbE/KEx6GVksEc/RCI
mI2aE5dNYHSDB0EecVc5LqxMPgD+pElQS7qJPfh46Gs++N9CH5ZJdTrDkBPDXhTZ
2agFHLUt248y0L4PPDuRoAeakOQTipJ/FoeXg8jEK9Vaq0iaWbNjh62EbhNTbwqC
dky/lWfzTdan62MhKTiwph+NAy4S67DTnDhONj4gmYEAeT9kagiXQrKARWEiGXxG
c5BABA9QR12yr32r/pGGH5+QdZD85Fk9lc/pW1/7iUDm6JMGmmR2sMVaebl6s4vA
bY2713hy5BagNKXJ3K3CwxOsCXKy6n8JEdUPgRjdSO0DicOwHjp07bx5FDkrnodm
FL6BzIiOMKau2itRllOAKcLMEIZFF6tJ9ADoF2DkMDvA8iBiayAVEIvyX+Qc6QwH
bHTUuVdjidS/Vmy+NYyIRAADyHB2K6MVYNA+PjoRypGsz+WBwJJaK88wzOv4jD5Q
4NEVTyTMjYIoBC12xRxYxCUwziHMWchZBfzLn+Ek+3qrV9dUMh6CA0FkcXLEaNq/
y8VENyySqh7cdWzOHbGAq33sQNXQw9v2iC3ekUMbCOcRyh9iHvcOiMM5sJsmRkQD
N6dQ4OqKkW9+Nm8Nr00otko6XmmZRPhTkfU4ZzwQM4B7CDf8IO69FStop7dnU4Dl
r2agpeSmCMLzXwmbd4owH15fx9+OOj352+N7h/O8JKrc4oUPlXD3l40pP9XfGUfS
BTSf6W4pCIk81KLw28XOGHkqrTyN2pMzYI4B/iorj5JBrd56vsYgpAzdgJ4jnop9
AtAhU9LN0fUywGM54ckOY7pzobTdUCxhLhQGlgWIXLebojcJlRx6+hrlSgYJp7xR
FNrhyizNNLXWaKqR8mn5uGrg/VkzbhlTaPyrJynDBuOXwMwUR3ykz6VVXAy9Dojo
oy612FxZIyYJlYjsu5ZtJk+JhefcRAE6blBu7FtjULWsEgD0Z+/aZfLHQVWULq45
dV8y6vt6DzURFaKS+QinmZx/wVHZlKsQ5OMwL0vvXRG/Roz1YMIQ6CbSu/7R13rB
xOLfM8JBs4WVH0uHen6NtXn4hZRm3cW9004RwbAp7odXkfO5VpLeNaar+6rVEhw/
CaPuss9ro/LDZ1BBlrIoW/AcJ6ZFF7eBc2k4/pwfPE0WAVg3clOqJ0JKgM+JqQtm
X/1dqN2CdQ6b3N3qq+itP/+v+d3tndTGkryjUAjCY8wW021NDW5rQ2VlimG6lYHy
Kx4wARtywMfw25zADmM58S4zq2o+zsV1DuUjud9+wfxgLNwZsFA2em5HZst2pGCK
DhIgbsbg2x7arBBbyWZ4XvmdbUJuw+p/Pcj5PNJt3JC7z7eeNWOekqDCWSRVV8dG
cFnavSth4l2NOD7Khzbi0I/ldOwtHHseb4cRhrtLPq+qnhAKpyDW/pLFinGV7KH/
gNk+LNg29tZvH/w7xstuT3YeMsTnEniPuKmXMNpUPlsM8cXi1SvbHUJeqojXXEl/
14/OoRk0Nw5Nvo7jkkdXB95QOBv0EqYRrMpB+ET7rC/iWmby7SkhP3AcURuOBHZy
vprFoGFa/fNVQmppLeb/Tk1NwZ9HjD68Vu8uq6QK9gir5LIEAl9M1/CAcGlfzosy
3sVn/t7Cf+ESQM90ZSTC6kInKZquOXVtY0Noky3XXbA/3CdMBRulB9UPCtg7J4vY
+zVa/5DIHFWZohmHZaCOh9GoLOTGmClsS7h/6snHN4k04G58yt2/ShV8uXb+Vqcm
jNzWXzFwzpv0k2exokm12EoGy1tbQoomrNeh4JOTeARuZrbh6ZEWmqrY6IbCnNIJ
0hqLIWbCA1V1h4JRctvMKIaNBRYXak10cMtrsMtfGzLAl2zAfAMg9SpK5uYA5T8Y
bD+y3ZxvfCdPcz52yXv9EStkijKJfVZ8xVuz9bZD52jaWRu9u2t8xqj+kCNzgzSZ
2iZAcWJK8mx88K9NDHIo9cwfW0UsoVxqJfjYqZcv30/n99lKNPtaDdWxzBUC7R7G
GXNNpJDISJ8tX6xQV5Pk2HQh4EeQcVu0ynmmD19MXrxwHOrfvgnDmyKYV8tEC8ls
zlzoKA+v0YmJCSM+C5NpFvk4bWjJcVHHywennlhj+hCxBWqo9CQ6icfulIP8tTEC
p9xv6/aqkDEFVUC+31XadbEQ9a8RZIXsPgMRJ6rVWViKpP9r9iFA2bOJZHqOkury
PWFQuRPyuLNhps/ve53PCOO2B+tYsrP7OsjPz7n+bBtrl6yOov8Qbd1e49B01jDy
h6kJYLkwlak5pAocmx14afqI9IDGRHk21kH38q4aj2IcZ0KyQPplMLh86fVltyQR
Y37V3tZd+00I7KRopOXsE3mr/Am927UPFGMd6a/0arvJDTEUCfR57or+WqUeuHeW
NUpaN6uu1KDmSDeD98LAfYjR0uQmapvHGG7EG7jEYPjtTjT6oObID0BR6/xZvv9Q
GeW7hL/UdsLcWwqZDKR/iXJO7NczOS2/3HlxjQTPpybcZmHOaEbndZjFYXFeJnK3
apkBB7xNJ0787Tj2AaXMObcVG/ObwZGV0pkt0SltaIi1V9bs0L5TsVIKL1nai9+j
XONxK0po6VlNu/p1fImk341Y+MNE6qhz30l0KwOSErbQdybxki7nn1lQenOWC3g7
zor6m420I6NsZb4zEbFiaPhxtrCmLbIzLls58IZ2cHiTaGT+m/G++ciDtKrxPOLL
ONVLfglUc+tLRdCqW8wZDIIvb38BgDhXYhClu6h/qmYSXPaMRPlSKPzX9uk7O7I2
nX5goAUJiVhgmpi6QUo2MKXUDXWDX/C/ETkqnjV+QFiTcnmFYKXfhI8iHyweLKrR
f6B/tgO5jfaNtnqBO5XSkwy2p+WSi0VwCZfuSxXo+GvfEcm21OrzmKBqyOSsHp8u
7w0XvgYS9/X18J4GpAgpSzQTZfNfsAVFPtzo3TBC+ONMtba9t7yr6sPJAASNsyL3
O0z2DPKiUt2MEFqReA842LvBKYp/oA37GbiO6QpWix34dMTRaBen3/ULsaUms41h
M1miXxvKenrh5vRhGaOj0jHYynD/uTuk1zjzY0rN4NvUCC2XlCTaBPqaeftTFbfY
yK1pV7n73cptCy0uj0Vei7/9n6ZEuefCKzVz16Dg2INJZh/4b4lK7xPoeJ6sBegt
EuaE8AMCyzcksoYLZczcYc0S2p+Zg1uyOsvkBac3GiDgp3gtV4uHpxWm8hpHZuw/
CyRtWL6UhsIEISmavwQiPvn6OqFvttNlnE64pyhnf0Agf/hZZXWZCGVBk2iah37q
ZIj+02YBky2OqWoYtufOXqSbNbU5+2xExWJ/H9QHAffISwXeKbld+lzoPYau60Sj
Fcgrabuk6uZGCcnHALEk1S3Sfiz7j55HcFrYlnqHrBQznkvIe+RXriFmKTXyWNgU
K1M6YxcNPhBCgcDgl498qU81tkmHOfWOiKPMeB71ER+nthyM04PsmaLIc2u+C5nt
sYm503rgW/RcN74dBu57V55P5XHpMHhEijj/VMRW8iR0hCDup55Dfk3hav4SHdgQ
Xux3c2nv6uDUf9IchTKByShZvubnLlU8zw3xs7Bn3Oegtf4AVMsYih2vmnB1yiS7
8ZG6HHOkyunlgV61NlCHVRo1WLLrk/i+CG9pEX5rVgcKPFZX+y7g6LNKYItk8tZJ
FfwMZc2JiadjQY5qsd6stgko1Z6h5J9CETLNHlQoa+DB1uAjMVHeR561JVU8eriv
1qC7fLacBCIeSv+e5LKg6/Fp3wz2nVxVlY3DMsq3heO2WBWTJCFkIhYSo5rDt9H8
9uGc+vUF5JzFenYqUOhBKnETQGz7NQNSBb9E27BcQyQU7vNZI7tarKHLuvoP4Iwi
N2Wl4z+dc7d42W/K5XuXwh8YbbJmA0qy1qzZBTIzEIjwx+NeHTWnH/Uwwu6UwBhZ
YourqIFki0bZGIt5t81T7tQG6TOFWInOd9wQQIo1YzmweHzEpAD9nsrHyzoVh+Yp
zoFWdLg8hOEbzm2Wgz02+RzZQgOrQfPiWfOfgGaKLiwXQAfnfBKJi2hYgFGXSkrT
5XsNm+JxquLRuLMQghU2F7hMgb/vef1KJEfiAjZFzWr+XgUu7bkvGyy5ZAMSzIl4
CwCBFhgV4tzsqbYgDTL+14ch8UyjueuA5R5/IAJz7C6Y5nvri0QPsEbYjBeRmkci
kdNx7KkDRbvfrT36ruSpyej0L1jYDXrBbCwFOl3oL65Zlwat0CbZSummQPdxKZiG
9mjQlUboIXnxxUfCGt99PYfPbjiVnSJX5Zcsaw9Tr8P7mByH3FVP3MgWGQ1xyB5Z
v9qp/DTKOOppaWRmAGPJ/m6B6o5w0Gy3uDMi4nuDTExuX0Fa5QDVG7V38Jy1oM+j
3wL6u645dIRmLomupHCt7IFC176Q+xIyGC1hB9Y0qNFSl/+kVmyiDpOlpponU9oj
1dVPQdHCREfgcYgCOYObrapx8xmKsEyS/Rdf8yYMZpUtBCquWk+ou01VzGJOt/s9
WeOHkAF8xYcorCTwOqFn/JATariUH72+OpVmm/rfSC5+Q8nLhq3stF7Jlm0xhnHZ
W8XM3LCpC9qXz+iNTWfUZDicnTVcSupAe/GHMTZnddYtkqq15rShvGP6X74ar/oT
pi4/CxuQ4c9Ur9GvyuKF2Hr2ox7cMy3FUnEaQDtqdEfkn4YNo2DWVePitHWZ5fDq
yVl6ESiRioNvDpQTf2drcpzHGwCwZppRyBi0JQGeJrU3JpUq3xQJAQILgWb1x0jY
scktF9KJNPd9FGq4JRtGd93JkVQBUV5NCuB/ecg85iHdSHosOvIbNuOuaKr/SirT
9hhs0IXE7s0Bsowdb+5Z+zXARLZvojUkwJanwj/O4hJ6Jd23TePxYzIKBBOvwxu1
oiOpUEDrKXIiivOYy4FzztY6VERt6A9n8FKxTDEgjm5pq+vqGvn/7q3eBDUFeOgm
mO7yfydV24Ia7WEQSasdgS7jEd0/jfftM5NHXARRsaNiwuiC9Bv/aodgEgUPzG0q
wRsNUKRpSsz429G9S56t8BRHtBQmDnxC+up5CUHHnc1du2HLLWcG/lGk11SuxHMv
HKDWP51L4uDOF05SYia7o+fkah58rff8p0TAlcHH/QbPIO7mdY4itQwr4SW9o+uv
6FYxGr4Gx56iqnuXjs1h9Dmxjl9xWGad/rbAg0/i/YbQOa0QnERjSdsMjhodoYuw
2SwQDulS9oCUo3UoYIX5SPyyRhTSSJSXISzW0u9wJ+Q2sgcwqh4XLQlV+S/W28TU
eWGUX9WJ21BLZu4cnnKFiPoOm35GNibrO47ZNl95q+xRUx6L31bGE6dXXlEKN6LP
8eu83qwKiWs4ovb0FgeUmvYSWNIg0jZ4PLXlE517ofa0bJ7zIAJz/+iJF2TA8OF6
AEPxudKKNMjH/9AorzowzstSKPGf70U0Te+KgCZm0mxAT/lnFrknkwtBfwVI4ODY
CdEm/tca31sY1fpwtlzFtRJbVEzkm5k92C8D9iAwMMU37Lh90rKEX4HWQ8pu8/Qi
Xr3tUq76hr/kEs7P3ITFWSiC2Khun8yliaMt3vvyo9qFAo1r15HgfCgImm7TeNYu
hsW3YRaJbCieLsl/rpL3SoVMX/TB6m0a4f1NW7F8kptpUwTfGvY0kLkgdISiBAfi
gISCAT/w9hLd1jV5isLru9QYfnkw7WfJQxDavDrOyKH+/n4zK5PO7AhWNJQKjbYK
P8PN//59htM3n5/X2VKTcV8FHB0JB+B+ZC3su0JBl+wOplY4Y4M1e6tCznnhYOYH
aaB/vbiB+iQ+mw+AEUkbdFhAmg83r3fA4BvfRgcJYbwlRzLyxIO7AowwyjfW+n07
CijIFtAmihl3bugZMemk0ra13hIctz9W19irkBQFrWSE8IJ1lgIMKG+roKC8H5+d
SLsX3z7CO4XfEralgE6r60M014jhLKxs9EENdyS3p4FLdgIssG4GX6hHTHuvzsri
zvt9ULUoQJ8/bpJIqn/hGyCrOWCd8/cFncTR8ZQRPbIfrdsnMwIFGBz2sNoOBZx9
RddMcFVNpFBCtjK97s0qK/Y3Ldeceu4P1TE51NUqrVyKj0TkAikz8rlwvCP9MFeN
QJZcLNvaCLUiVrP+2aAAwdaflp5lcAvDXlg7ocAjq3yp7GE4suDWIbfxxo+Cj53i
bwKXxJf4KpuU+3oDdwvE4AInc1d3rFCTfcejCdYEaGcP0NCpy4htdqoO4rV+Bq9F
QKsBelCZr7cNNxNTn+IXDZiQSMH8BzY0GemmjE7vVSfbqmaNeiLus5GEqxtQJ1Gg
8XDw3gNiFCZ18CILDkIlqfUchIcodQJD4t5BxuSL4Os3uzFfFItVsG892ZXMBVCq
DHCIjXkMw3oV17U7aFNO0Nev/tP1VNX+2rl0JIolmhlHH7smNWxerQsW3DJrwaBD
mVHbv+/uyC0mwhirvi4w0p2/K15zROzSfJInyCX9n+vFqhUvLC4GUX0VyEswt/OS
nDP2vP5PPCUGceWSarMeIekkKz04IeOKONucXbYRcmkctZW9QOoL3MPH/FzcVbvx
dEJ8rdL4LmvbvxV4fcjPMBnDkpNd09bvr94Q8FH7wpmtc/HKVz+seXFrIl9t4RxM
EdruN2zcALqeVlt0X0Zz6qxykjxUUOF2B2tcIK5e9mG+BDGidAwiIkgJerb0G+0r
6eFGlAcp/MNQ7gUgwHcqaMm7xIfOBL8ej+ofkQLnr9HTomZ51qzrwarb212FqcKs
Uf2PlRwdRV3JOZ98OTJ4qlSpuOufoTvYIDAKovvRq8Sd8zCSlJfTOIVcLlEXxo+G
GOlrVbaQYHMav+5Aarmbb21IQaV33k9zRlTkuBmoZ04MdNaNZn/g1HOq5/TG5hz4
f7qVlCbEDNWBFg9AY4VYIECvjVT7Q3zDGiR2z/4ZLR7eHsyPks5q80bUKWqag0cm
X+GsjvcP8iCb/+j90znaR/4vAQhmzkZFcKBC7NGdmMtbwUPawQgdInoBV/ZEdJSy
e7E9ji0BYLHD4Ki82/jazR/T1gdEPU9vuhGYej2BlHdBBAnrINU6Imh1BCq6t9Dq
+N1EVdDk59+n5/gHEZrswlbncfw8DpjqkNW2Elt2eCMkM2OwaL7+SXz07NCK+V7l
BC3uYrAPObqqONHWDJS6doyiJnW4SNQo8LknGko5SOYZ8OQWbkrNIKq/OVI3zr/D
R3fyNCMtSGPpAg8vfJvrpG+7mDZlveM1QjS23sCBWonW3bHntHLHWUlKpACn0uqb
RnR2z/DzF2B2iJN9O7Q1A+dzt0H4zIgZr1qr/XGHU42FITVrbs9rtU4r1qJ8mNGh
8fjCoo8dc9vLl+pt5rjPsdnTQWYqYRDDpiy3Vf7MdWBEp4ACOb8COqweN/y55xBK
jHI2KD4jBP2U3VXisvb+DRFj1lma6NOR4aZsKeHPb9qK8cTVgg/5DLXkjNTlcNZ/
1CNUtZ98rrFyH294JxJQk9lxwJSpXZhlp1L0Zgaw1qi56lTCqHbwFwPAZ5ynhOx1
2uYolLSawGou+XPh9/c1WGq3TKVV9iglxqUR7u4BqnOkZ+cyLxwOLim2SP4nxxYu
tnIcMZvHYoO/xeTdmYhrYN+56NmIcb9CcXSOGkgCrCUWzAzdHxGjeCP1XL0GG6Dz
8bJKKNpv9ZU/SCRsYa8dloS2GAuGTEHytFAY1bSQaXXXbwxlHlkEFn4yhwhYlLPT
nzMk5EYi9TkA5sE88EEqHaXhM7Wf8tqx4dfCrI1DVDtcPtnRUH8DjVLFnMv0RGb9
Lwtfj6Ge3nLOQKJRn43kDEtZyiqeSUJ79pD+EqElvqhKlA1hZNnDEgK4fcGTxx3g
CqZ1zS6EGVPd9mg1K27kiApl5/6xVPAzEENlXUgOFwTXtTnRc8UJvCZ79KjtPg1z
vSVOnDiaTdjtJy0zsF9BSIYIzfQ/naIjTkRxDwUw5vjnPjoaexWAZDuMwcwMi2c4
Gt8olymhorHA2qK+SXpugrAV6M3edtydLysVfZSrH6/kEpci79hPqURnas5uK4DD
JhTrqZd7sVrnEmL59tPB+zPyefAdAtayEby3leyFRpQ8dX12U0HJKBXwuN85+fi4
wRZa9OmhjIQ+Zq81a50Fo5S0t97+7PlEs29IohKEo60FXo0gsCle/LM0yR3JWmyS
d6T5EHL4PBDWsXLzPjHqUbZwG9M+kTBF/FMJmCyzggL81gbX1hf2aTHK0l0D7DkT
xbe8cOTfVQPn6JYDFvTGapbpu36dhXJWxfgK4z0BfZg4P0slrscJNcbBd+0ScCJp
+KYHUQsbVkKCj0F8Pv91RvP1fKUV6MBPJfjh8jBkeb+d/X1JegBkd/wwzxYUYUPR
5bEFR715oJCKr3kGOMXvc90qaR0OFeDsQBz4th4IZ4pYHjXGs0NnodPOM0AH4X9O
TPG13ArwJj/Ucw0IYQQCvvSV4fOkPYpU7r9ZfKEvtk4kZLrWT/Y1CtcXy21Qi3ve
pii7jNoC1REn2PSQD+jjB03vb/tepNO/cAW2mAhFVl99S3jLDjsolgSZ+vDxUN+S
1mrdLttHWAApaqu2qHJmAI4QZPDrNQLlKsQlNDS5o5xEPpSIVmdD6+TA8AT95xvZ
Os4BmLnYTLwuhO3RzB98FcaVorIAgx+ptwIyqmY69Z3DWlXizFWLrr/Gyfy/VMOy
90oKEyDrS836vR0erZ2CddbQV6mT8uQ8p6QJo0BHN2S7peaKv9QZwIrmlZmql9Oo
LHddWX/CsYTC+mQm9RHgB1HBcuHX/xbzD6qEUdeljNS1/Qvqavao1mfTEAMFkF2a
ybY9h/QGaTV5BgvWu3ylWUFy4RzdkffeF44gqjB0+A/z/O+tY4q2uYQ8dzifB/QR
jeU286SLbeUSBkk4HCZrr+w8u5GaClhlQ4NiUASqlQdgUOWxTGB5LYb9yOdo+m/z
NzXIsegE5JnF5TSVZ17lzewwMCPkgKZiuox9+IZmaWs5dFtmHfJUxlCcKzcXjruU
yupjebcKCXEd2PclFWST6/0HhB1GajcxWVccsReJCAewpbeToGrKdfxoLAqWejmY
smFr2V7Pv1RiSFJqRIIa7eQ+CXPE4wIAsIy6t0bequpJgk8VWSxwppJjdWL97cqw
I5bOfH4+L0gCkZnRRYKtMDdxbjBlpiIkokxBNUa84yK+QqAxxChUhNpr9vWnqBUl
YdqyvavB8hRHVk+Xmdu8RDWcHBlkfaWuAS0yv4Qj34w=
`pragma protect end_protected

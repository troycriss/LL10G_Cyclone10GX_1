// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
Uv5FMoC7q+spXgkwDzav5mKcUJAu9WuD2TJMu1gfb04MUkjU6FfME1kiWahfDxEtBwaWkAmvSFyC
70ey/gMItVq7EZntsSq2t+B6pFnSFIeQgZjpARgQtphYr6idLWDhM0W2kDbpSnVOeb9VPf7+nj9h
bveBCnXpyU6uQmO9ElEOCkGck7SBLjWGlLcn0bgGiDSioEheD/F4oUgnSVePhufmitEbAVqmsBAO
TLYJAt9fXmIhsD9vSCiZi9KYaDqNQcCRiWWq7bN3UEN+ieHNRzmq+VAtmuyMVq8XGlc/OlyoslAK
976k/7Kvaf0s2nWDLVF3wRpMfyvwcEGCBZFe/g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 19232)
bjO1zCI5HuiWUJ6W6xgnNZTDu0w0c128me44L/aEEgLH77M6rp3PhFBYlAPXzZ3Dru+6GhU+iux6
oZjc9dV3FEX46ujqe/5nDJN6pa10MZFyMiniJwvWOuP4mR2bKXE7TAIAOrsfnQ5Je6gbJWpcJqzf
pBy/0gN3sqUwEGMkDLC81TczwrWam59bMGdSEKs97rjYRgBg/werjh9/7h106jrNa2NG370zxOyq
UiNte78lL6APkUpu9KfFSZcb5iMWPVS/VIu/RTeeBkPsTvqfCnNtgAfW4Gli8GCUulvhRHx9T6sU
q1k7h3Cu9hjKArWZOi2RZrp8mdLzJQ8TaDdNotLHO/HkW/8VA0SBoDrCPHzZ9h9wX990subSf6Eb
zTC2hSlvnpl5I8LoldxdboOBE3DI6RgfUqlWTgmsNA8mUzBMvb6+U5OgOEPSh2hz0KJwn08ilGEG
wekAD4SK66CvU8e1b9A4apbvOvAPM/OG0scleZrS0KMp9BJXo1VxtMVBeP8RZbvQtAcjdI1PXQxk
NeG//oVn2/zvDnk3QPKfQG+kFa4QA8j3Q3BbKo6jRFRe5VhfvKFpqE0yeilDx58hTXJ1DpIY88tQ
L+JSHfllWod0YIagYYqXRVYrN+/+lGQoQ0vm0qbZyMWtcg12yChMttd/aqP/qpvFe29ISyxEVl6R
KjVTHoJEX2CDUn6v6lIpEMgSkio6ijpjJoI3J7e0dp5lWsM5HhbAhCKCA+AaU7sbOGG45n1cjQjp
laG6rVbv1a4BUghe8096KArJOiTEprxaSTB5bBPXMG6il1tSt2cNQ9F2PNO5ISqgjdm0nBJJuhs8
ww9q7zHIIG8e5YyQLQdj1Gt0Iu3I79fDliaCPGcUN0aYuhLjM0s0JM3+mw04j1QZVP1BflD5ZaIy
GCXLP1srUGPjNA/uybuJD8fKY3mhqKPIELi20NT8l0As/QR6ntyVhGDGQwj5zlMPq+LRMhnDV97j
Qwx7X2Bu/xFjrix/ICW1NtFcoFUiTwGXOi19F8+DQWGaxjqQNzbPSknVjw5e2RE4FqlvThN72MlV
tbKDUpjFPJMxBrD4S0DSM2pzLFAi5BFf1Rr+ZOocDs3UZYo6wcL035yYDM3qda+0HhoNY2Z9m2Wt
YTs54XqiUdCU3ZrDocSlkF/3WTaKDPjnYhRT7vLEeGA/dU5peMvEhGlFd1XfFSbUc8FNb/++svbI
QRvwlS9NR+swxVUL3/MtIb2ISwtT+RgvTiT34iuKBuNIquck0oo461PtsqLFquBFlvqrQSso7Vwx
h+zap7CfDwtX8MZirDnlO5YTuZSaNxcb8/PUeft6tj6AXGnX1bMAavvzegAdNGHYjT2wJk3qNslA
W17JdgV4yfHMWSTUsSOynNE6nekt7d7pbP+77I4h7N/nKsRYJDqVfUEsNNUNEMMjrIxEax++Vm6M
KrQd7PCzOVZ/SAgbjNyTKpRBN/2PkXSoTwyA0HTrCUeADSheZM5P4Ewy1hn+7svX0HgwmJa45Dk0
Q1ZGUqZIJHX/XvZEYMrbEm3Xc0DkZqT6QlngM4j586Ug+LTrgOU0jRyrF0YKH2j+Ix42e2JRB+qa
MwAlm7VfOUA2nIaC5KMjp8sxY9LOSh1Uzm4rDLRY/BvWB07d4ykajVXC2UKDHKKF1cdq5tughfhQ
SvAgZTN09EJEMbtPsOLzdXj3DLlVDtgkwBTdrff41D1009j5d1vB7r44TeVKED2qqA/9DST8Zwez
nBXRnysX/lCiSx1QPuvcSd349NGxwWtkPZmzq5Ca2gfhN7RXfBfasKFUNB+lvXWR5BBOA4LGQrco
y29bjE+1MMNql8dNRxDyuBwl1JML5v7zxWahr8nmcS/OmBmhTn1c3OwSjOI5HfUp6tCZXYhtTMPi
Z+yPUPhZwi+RZ45mjWyNFE1/KxQUfTR9ojIWtRRoAR7JttaYe4Bu4LwR25LLowFo8xQYDzWuOcFp
2i+esfy1Ez3apENd5oBs6r5TZ6qtdNMyPKYEeBoMo8NZMo/z+62d4/FIi3PjUZYmO7NweVV6Eq1P
w0M5pnb5svsFhv2mhdP597EQq1zCQuv1IRo2GrdvRToBtK3UaItglRMZIxvoOE7Hd4XgUuwxGiR3
Hqmt1jcym6Kwv8KgwrmcDxSCoHcN+Wj7nNzABVgT3180HcvrHrT5AYtLGvuRNDXtxD7tt1YxZqJg
xxs/wPRhm371RjMCWvDZqpU2psKKAdP+qi4Lw2+qsEm03sBoJx29B8+rCLhkKdaiz+5yDLOztu4P
GgDsxTv6oY6Ag1lNY0QY+FVzzMVhYICZ8hHbXr4QKalqWjEU4o2C65o6N7ek/W7vuD8Jg2k01pXN
IVFB5rDl6VE0ypzbGHp+0TjGzU2/V5qoF9utI6hEjRd4Q2W+U9o2Sg0JCypxk8MgsRF7fUhQGLAD
RPnPSXSShyEW3zdiHoLD15+h1NUzQr2q5FOeNQD744LuRvQLna9ny+wQ2oM3veJ07syp1ngl31yy
g1dPNnsHQ8U9OvEqQ5cR04/WxwRdE317dLRfWS3x8U5muUw+RTzDou+53QCZHKuZ+UqZaGb8VBCA
ZyAlSPwcr11oZwDpn/InwNetQk746bPLQI+JjtBax0Csh0CT6m2C3Rep7Iiy8vH+u6c3GehRuLj6
INsbUQVbKKie2UQRuJvPRkW/WFnss+2TsL7t8AactKzN+CxGwfsAC2zG2AhhhPxXaRxV/rDz8zqv
3gpjZz9QlqdkOOK13zNRrk/FjxJ3yvQPg2dSl6WvxRHUzVFY+ltDUEKySPxVaKUKZBenrKFDOOg0
8Lq/mq2SVk/litRhSshH12vytXkMC2+8ISZ3I2lHIx4fUZ74xXc+AMc6wb5kBfhQtGYcZdIaQy6O
U1Mgr/nmPCyhE/IcQqhdi9sK3P3yDYFTNyVY5nn8lYCOA9zRKsfxE7kKd32/W4/AgNByWU+XksnD
dG/BBJaAHTEOniuIfw5DkhtBKrz2NnxPppL32/4omtEyQXpTYMveo4OwWSSCh3g9WNXUF9XGwAJT
lHasP5f3AlWEZTZvKt/IA/Ga1J+jKnfkILzqEx5gZzI9nQKRD34aR6XfwtjPZVjEpnGEkIfijHOE
dXpTqcuLy6/48lAKYLPlj6AWyZIdxS7aQw4T0quIHebivAbq0EL45Q+eSCidPijbcTkb5KWGrovq
ZFWj0bainzU+Ak3e2DAx/A/CVVALAp3lqEaBNFAZ8A8oau/6Po88sCToZGkQzPMgF6uxZdbTM+cY
YWkOXeLT4CQsFeMdjO+5OyDDU2/+Sqe+ZE1deHmUuVnX3X8TS+qFB9jNFmTk/uP9ADrT5IpSI9ZG
KHjOSZaLy2+AuUxIE3JbwDJMdwkRZXwW3FkGwQnOt5sMdX6M5Q9LI4v2QwbEZ4rOaVQIwB8HcCnQ
5lT9Ne49M5gRKR+vKT6uPYHSEbyEkMAZP6pBOB+2KRA1ArbolSYXZ9C8w4iK/vTREJrfvVeqtFnK
AZb468ebe1EVemrihYhqMAga679/1Woc3mZr8fPx05g2l99TBEEsxG5D0YGZ/sHRdtUqlokCbY6c
xJX2W+TESywRuYJp0ks/0MWChg3tH6nNib3TGahplhn4o8NDB8bL7P+m+ngsAILwUazfOF0MtAcS
dUetKMieP26aFflij04NpxJaE1RUxlQpVhhZ/M1VOXG1Pxe0vWPIwkU5DaV5RgO0y3X8oDFxwDwn
HGow2rkBh0ZEVs71mgdWMG09/bLdAAj/6UrCBCIvVIixnLnAJYQYZkYhAilFfrD9Xwu1Rjgc6O5X
1KZxJ9cYgd9D7QfqR923yzinpOu4LzIknFHnSJLG7eU3Vlo2f7gbph+Y2iSKkwj6y1HH1ZkgBXva
MLC7qKirv//5RKks6s+g/UVQUnEfeFLnbNycR8OQSJHHhZD5jsgT1+FwDTLIOH7iFv0DlfCZ/Obe
Mbw6e50+HVeOYHXB23hAEWw8jcqvJ6hV9/bKGL4JtBxRNDNBmacgvnHbxmwN2OkXFZilTcsJvLrb
Y1ti+kffbrcqwFUG9ZDr+2DXlYwhUzZ10wnUxpvV1z7X6iqZvzAjov1iIL/jUA5fb5q9ZVK/zfgn
262g2jwuS9ZiO5kpyevfng9ZWs1dm6BcvpNq5Tkjj4tLpV94dJ5iD1LqjRWpgCcOpmDRpMiQyVxx
uauz1VVM560opBqVwkXFafDVLwFIr1SjQddevPcxuV7q4WKA547+u3qoGZ/Scj0IEXItFgy2ebUD
zxstJh52iBhetrVk3mgwM7+GhHCd7aGvgNGt6NmUXI00NTRFKletsSsZpV63bql25wmsep2QTiCl
PTRboHIpNmYNPyPuE+OWYneAOqnozTjJ33V0lfuykozlulwWvraaHL33z80/ugKZXn5DdrBrkV3t
/BZ//0ajQXFFckloiczlrHXxqR6oqjLGxNT41EfOcABP9mlJvJ+nLcuROl7o2P9cMrcQr4Nnkk7V
RjJRM556//TViwnbSUVzY0l7Z9Adfr5/QJkvbutaVTkeMP9rCEL/yEpfzUlXohBspOISJSSiaadl
SkRS6aBTRi/IQb9DdsDV0UmWwSTbVcbLE0RKvMpurJXqXdBIGP+yZ6nOXikJBU/DQlPkJTjZ+4Jv
la2XuzJPOW5o3uQB5smclPhBqAs++i05NglsBvbpxKkIHWjK23Luunw9to5PelRqcwDpsci4Okbj
gQ7jFYOLb2oBUI+ULYVGkChxH0P1uX8XTgQ1k1qHKXVR7PvpscLvtFJK0jW9AoMkh8uAsyR40idd
qf0PgxyyYpSgPeWAE9Wr8iQOsYLRMGkwlBTxv49B5NKI+dr+YwFhaBg7oxZh8vGVem8KmMPHwBNb
4on4zjy/52OKBxIng9bsG/Y+3/Sc2R2ZfrrkqWRNUA//+BnNYQR3y+v8V1OOQcJq7Rh/cclDeGvt
VN9Jo6Dl9YQq9XPdn+Kd03KeEWL6O/Dn9Fh8N2aKmn2Pw6aXIN2Sges15LuIJZSLKgBlmzxhtZIw
qgdDZl+HFV5++VIf2shU+XCYfsrIfIzTR9pSPDCUSBhkuaDE5vMsz9hvCz0V7EZ7uwig+90anwR3
XXDup5aSPXplLlzalWFsKTb80nx0ZI7tDAuAukTHNTsQuWcCIgGyRd2PXNJg1WBT89PjdtT60URN
JhoQxoYW20sXNT4w+pjgX/NXxu66AcQt/We5sKnpXZDBDkfP2l2zxr9qiiE2yUmmSLN/W9NKuKP1
15ThqI7pJFMk2TFHotu2Hw8kIybI3O3woYnW3bp5JvTRmSJH3M0STETFrPPsDgX9uoErWf8Z5Z1g
4awalNGt0cFZlg3CtVhvgSUhs49UTq7BCNhF6ik2R6nemHXBvbBsU2s+rVcNiPlWWoq9pyb0GOci
+jiQUO1JCo5V7F7vra7H3DTL5MAOmHTM3XEqPPfEZmBezbd3WfSPtzmEDs7BF1+ksdwQ+HjtxgZU
mLS/Tbvs+j/7byaH/mF+HXssrMyfHFkVF4dxJKm1eqyDmXwNaC9Dm7H8WyF1BdrnKgpwOG2h0DgG
JriR1eoGOmMdq7BP5G2IY577Rm2UHriisipnBmOPuftI/6b3000jgNnEgsyl/a2DOs+lI24+gx8r
t4YeNQu6o8oR8C2r88Pd2cZoFl1o2EBfHS+adfAOHFZN9abnO1yuAorgGJEr1uaCUj90n2t/6v/T
RlNeR/eolX3dLPPqKzTLDn9mRywQa9sRl78yxI0i36s6cje6ZS9dJgD9jG7NXUWsezgFaQl8itFD
onMpeAe4/nl3rsJn0cF1Y0ANzTAvYlfJrQDa8YZg+rm1tFWSeHyMOKQ2l4cmFhMnt8gu/76bY3qZ
t8PPsqlz9PXNH0eVb7tz8FkFgHUVudCtOWWhPOQfjjZSQC/VXbwm9mIl9qdkiYwR/EPLZvb558sq
ehyePCT6gcmwg79BUSsDDn7X+58VUJaT4SikRoAa0vh3I9uQC3S2duECKISIJZyaLmpziknem77V
mWEluo7qgVf2xFQlGKEUfVUtn2rGKxoCQ/qyXFIJ9CuKbr39qazK439HAObJmMD05RJgnj1HU/0V
WqJnK8BCAL9V2uPo1FYMNn4sYBP6UoaRCGzSYn4q2vXpnZo22J5GWcjasggvBZgplgWj8WE1kmvw
7U73U+cRDiLvIz1SYC/pgZu4GjFja2dgjWKGHcyqlrLSyLahJ8D7kr8HmLXzPib7F1NHsZNkytts
GX1dxMWY5TVGnYD5v6u20TMuL0r2WzQRfs/CXQWVftS1616j84wwqbNpB969OMuNA4ws0piV3xMa
38oPrl6770z9l2J5buuIWGZiuT+WWI3gruxVTU2VEhFFmrgZ3Ra2TH+PyZTHmmpYzhX5cEqz/e8k
yBfZjjHoY+L9fXrOJkP5XicUG3h7Otb6Cox4EWGNC8qxnWA7bBMFtwadW2EtUiJ6Ww/J6KcmqoDA
EhRFarMHDWmqRNQXFK8WhoFzjysomItq435GWlhg+aEV0pl4vhbGNObHP/OwdEjmttyzNLRWJK+j
HyxORFecuRw+J5YMwOUOUDTJU13+67N7IFG+OI2f4RQKe+8EGWtbDR2UkNxFpqaaJhRDIrjpa3Mz
hN6VgrvMW6sJ6YRXtGMTIck769rpHy881g+WTqbNcw1YASXGyR5j4R+ytmvve30rkflOqMRUdmAe
rb5eSJXsTmYacYEnKPRlP1doJOJ9mE0TKFbaAte5pMx8ZXxXHwQU7kmvUqvOphgEc4YiGIpmWsWj
5WuIdC+6XNcFP0ah3Dy95K+F2oAhdb3d/z4u8xajUXSVDTu4KprvYxb4c2s3Cp1rMtsdGa5PMquC
zYI7U9GX3DeTeWMzdcThlSdeXL8CsFWTIKRA+pzHA9WpLQDyyJVGjvSQqwYX5AJic3E1xcc72IaT
huj1lT42vOxgqHTai4AloIUFt/RoCrUqIkefPzrcA20UksELCgYbg6L3x1saOFDzF7Ln0UvA3uFz
ubk5hgi5YszzRG7OvrwCBB88xCQU7M21Pt3Vv4DeZY/VEA1N+hi/d7Cl5JBZzwtq+c3frauPNdnS
aAVQ9k2OfzFzHoa6pzYCO3WCqJ9p0HKWw/M/DHvKxuLQJoGwJgNJWyIxTSme9rbyBlksK1spcMWx
L2N9q3PpBiWZlyE+R2Qn+WciyVJRjCoCU8Mkog6ave+hr/mHlDeqDVsK6WhiqMKQt/tXZrcelHFh
F+NykGItaKxK+/rYfOHRUQVZFFT7VeEb2CgmDe7lrBMRToZvD9DKncCVk+qQT8n/Ejb85SHjZMae
upgy7nvp4w1IIIO3QPmrlBjtd5SfiOZAkK1KbpTB4xgZsOKYqPFjRNZrBrKfdSQKQHkEJee9GVjC
hZlxpYp8XgDPuyTOBq9AyRJKZvRnd0+egCLw1a9gbQJ2wS1IhhFE0LIm4Yj0wcaLauFkzKfIw5WB
1bTdsq2Uif9Kh9uTethI9Uoe+vgFKAUEUdBaiDIkuORA50scXtUXgeaivNFODU7zsnCI2bqSEv+I
XTPUhQGwQcXOGnvLmzuNJJfi5Ic+vIyg7hmV9CSxhYKPHNQSpr9F7zSJdfH6EtLeHjO46G9QbK8R
b3R2UHeJdffsyfDdl/lY7QXDAqG2G2ED7WXFBasa8eOVeL2r+ge+bxk4VwjSXEAB82T8im6rfeZm
ee1dZ0LZMedQmLSlNE4+nngAq1LJolRuDshcSg7qSPReH9K4qa7MLMF88esmizXp1TjhXKyTGhk2
zgMonQovfXwNXQBdcVxl4rdPCx2KXO54z2NNv/1nWJRlMrBBYszJAe2iCzviMcOzUY0W86xj4nD3
O5odyX2MhJlWDWaTFkhQnDDr5SGLuXRbOMtStGwJw4WSVRy5n9rbhkf/YmKiAkhhLqRIkRIL08KA
ZJUemxO8bX2007x2liGQg/yVSCOSUgbAyYIe/2Yl8dPnlOzMoZ0Km2lkBrtk4WNnea1FQrCzKO9M
ruDjMRKzUmA9HqwrQgU7WkPU8cIKh/5kBeIxFOLzIaoGkDHwnCOZfEMoTJenhhpr/NWqNyzESmaJ
nxS+8ktSrXsvbr/FZxzYGFBkuHp9ALSTUg/EhIkhXUD/GS3Qk6hMOrmJ02DBNtmHeV7uBdjsff4K
AlznnSKF+NdQwYXQ49QW9GnJPi5fYLvPz3L7jyDlb9i/h6pfX1Hz5n3JTM67w+aLrCEHIZMtLT3k
7H6NeIkw+7CpkLgDqrIZpvRC84ZApw5ESt+COFLXjzDqqMeGpYKOFO+0NpTd/ZJ/vbqJH6ejhASV
w+S0wFI/La2lQICuOiStaT46tsg9AUGa0G9qCvLB4G5ejv/q5mVvP1xCE5YGO6gSFvXYqjR6Yh5m
Qfu2ohZPTm/9XhPue5mcwV6foW7RoJgl7XHlPN82bnHp0e2BmREN48qp7tpBCJQY9Ze478cLFIhQ
CTNRm5I3Tb3YhNExcqWmuBiAcaykYl+OTJMBcMp9B/YhvbTQzRziATToJ6l+GKTZqmhzfIzNRymZ
fFQzmBcCpZT+gGvy5LgXtGVnnEkuw/Ao6CjlEDiJXUhwziZ13GJsSv3Ndrr29kym2/wDGbmBQB9c
KyPjOon41+wnNpvIGZ7+p/hEFFn3aD11KlYNC0mckAtLkiyDona+i7YRV4U0eVeOIWra9BE4MsJi
JJ8Pp+gp/JGPZNlPSKmAkq6e9+A3R3QoxqL0doUfTvV6iLVBOss2J1mOfTfQ7zaKAIbfvwh5u5HZ
N8D42BXTFTNo7IbQnuT3hMZFFvEdUkukkOPElFsnSWBDhLOCTHgWBFyCaYdbNVDoYgEOi8ck6wlz
t42AcaJGluz4UiEOHny1ghOvEy8qcvew71QWt8XmonYNrHrpKcxp2fA0tYOuxd6ZTV44savfisER
7HEjwUEwtvzWKJDWxWZAxxKetoMcSsyGkSZtWI5vq6/OyH2YtS7ZAArvd9TlCFyDstLYp6yYYIqL
Sn0IheB2jlLbra6VXSsAcLTK+0XB9STVNKugOWzrq7ihHU3f0K6jjCjHP0g3vm0nB4bUF73F+L8g
pR5DPvYHu0mXUvKUbYy/i8sVm3qxu/8sEVn+X5KJKTbOVQh2rRcNsqlJ/n2OnGF0lwM+SbKbDdJ5
SavCZE1k2VNmDJIVj0zpIOK7Qi12GC705fT3+6WerhWmrHInBcreOUZ1fvmRNY4h23yuC9vbkJvk
bUj2nU+8OpTnr95RSisbZZF+87ourTjXxFnk5wfNBvLQ/4P6goYgDifqpJSAQcJsW7XXTsCtwOQU
WWVn/eIyBb0K0K6MBTn51BzKyHB7Vzy5s9FRcfQvLca+QDdgnxWGJJ8VEMV3nXz3MmoGecMWkqnY
AMJjyyz1fjpyALLZzoVrzIKbhkwhMwRL/e5OeJYYloV3a+128QcIkGdxUTwKk6EZMr4WrZpPYBjo
/b4moYovRPS6Vs/XFC/2aeDr4/vqZV/XXd/rfId1rOefm6zOSWGhjQiJYVImhOt5gwcMdRUkdjgZ
LGplMTIPUJMxqinpN7QE0mpHkLaqj1yIrcVkPdfhXav5lKQ2fgxzQPL3zQpgqTIcgKdjiBIXMUlr
mhhwyKM0AyX198RJEKc5s8D0QMqGi4oSyKTB99btRX/akF9uZ3ITVd7zXkaI0xLeIYGN1ILeCT98
tgV7Ga6YBzH+1Ia8Vq7ci2o+SueqLeIWZgQGrsjDiFjvmlRdCQX595L9/6xlsuLngGPlhoLwszBD
L7vqjUz8c6u1vpukE0R/Cd2AyzxQmgyUgzIq9P9I1gxJJLuIPEOj8uNGJa8quMDR9wD7nUdtWw/N
Pm1nuaut5qSRVyUwJj4hjEc3AKFxvjcwZ4Qj1ULhYtEsPIiFc+HaozU85ypuyUwrNK6rttW+GsZ2
jiBY2eNgi3Qh5Y5DhAZlO8eDfeZHg78IorYHSW8Ir0AN+GFHjhnnSIvgxEs+ayGshFBuHAaglnWw
GSwHf4niEu1rDzBma5Nr18vNDLrBUr+KwAAncfonvLNbVUMxoapevJ9qPgBJ14/syp7nUzrx6dr/
QHlNCWgoth7uYIE3uVGsQBvovnNKm0jgi32IJu8K1AHe9Kk7PVAVS9+rvLi7tysTvjF6cneIb5vD
DndH5Cbvf8oJN8GkbHsE2l9+ZUwSantM/jBZV2LfhW06nkt+rULD4fHbgf1L2GG6RKe9sEc8mXrr
hNYinmx85k3Dq15T0Er9be7ZaT9gn4o6M/CA3CRWzLTUmfzxHniOANu6lFLjrmRA227ZC1Hp2dQ+
xvaIfWF0lVWGcA9q6A4rGyE3hrMkYqPT76R34nhJPQ/8GT2z3C9zPab3MJ1M01tVcGpZ7BgpXOfL
Qg0efIgzHYudhxayab36aVT6Q6fzCyy9UmHqCSKTYh0hOhF34GLcnrWJXnGZdj86A51+CIIHaIuK
s7SmsBVSnVLInjQ70ow0UBMGN0mIDtLcimaSf7Cj7JdI0IXBjjZ2doSnj7UOA9YTr7IllnIidWor
u1y+hHyP/XyCpl1thQiU3LiNCLyj1np1GqfxmDFPyeIIQdki/Du91UYkv2noyO/4Evn6vFkcAO0p
nZ1DbPEFgWmYIkq7ib2iKJt3ItgU8+MtexO5NPCUDncMeT8pHXyuuwcjHSznwjRw4J+vpvE7G3oK
Is65Sv0LSYLsm4cSU1SF7SJbeyQDoGmPtKpD8zUdgVW2hP6GS/zYBs1vzusN+H84p0eYwTt/2rVu
wyz+mHjjR83v+YmMJHizQfJ7zmyBuQ/mL/LYaDhYwDHePMIpv8IoYy5Yocz+gvMECuwVaMR/Exja
Qj/C3NA9gSVDWNRr0KmgjngbVUHFgYCjJYMjkPWKVPY9vA9wcTLfbvnoQz9y3MCtUO+igYZkERD7
YiFy/hrjttP1tBV0HTXdBxodg4dcW+XKG//LRxZ9qUDFK2TZgy7gswKiSyZ5i4oPIu/1Upr8pk6c
2BfcBfi3sJKYGE788G7PHBfowDxUW6fR2AzUB7FZrqD4OQVyU6KUIbJN5S/G9JICVhdSdQC7naZE
IIfzIos9gYfNRmhSuiSwzZFUay2C1k/HuEOM1j1pxD/dO8b98kDh8eg6bBzQMgK+MoJFBGxKDMOS
HN6UzFM0MfmQXwAPyqxmok9WMlgGMKVA9AkbtkNQ0xkO4n/KPZiSs69xpm4G0IYvxcURmpBahPIF
JoX7QKfihQsAKfsx40SNKmavcvxSbTi59HfK4PST5wonaCrns5AjGeSt6OhUB8ehI5c6P30KDOuq
H+LAYCfUpVTRn0Zqm5+w92mUcfKf60MEm1NdlXzxBbqbTSz4ntY+N8q7XwMlHHfd18TK+OwI8xOT
5aZlg9rh4+pOAy/Avv9WTrmek5kSUxDyTh96XiIfl3kjststYJWLWLWwiulFTBd6bx5JRR/ue0Zu
drS0oUBHQI6dt6wqcSuzs8NpfsryNIARE8KnXHjJG4COTpl7eVHN3cHDGHlth2b4Yf0S02bHAJ9I
l87GUrdSqcBxfoHzlYR48Xo9QSCL6RifajvZR5idiIK9A8JGjEc453HUnU2Tqrh0aG3/hFH9n4cB
xXbS3VNKoiqYb8ESeZ+2110DJLGEp4pNmP5s4wBaCs3H3w4Fhmnpczs/1L8yQLecehGU8QYe+mbR
DWw06rPaFkFT4oQlmJTrJUs/hix7g4HYzwqMLpfwX5wUSkr699iRPuUhIDAbJP94PmxsiMLJXkH8
9GfctxdjzVXiVA9vBMG/k2qNsXW6zTvqLF1RP/DDQhKXST67RvcyIsFuDnloPn76H0gJLD5RBWUx
WoFGUE8bqrt6LUCZaZi5pTwF1rPhXJP01YjlDuyn40meIDLnbXR2hINSy6L+4P3AvT+1zi4w9Vaw
Y3JZN4MGdemyoBPF14kViqQgCJpoQ1fIBkdIjhKf+Rwl5tP0lKETjifEF8TxNJ4ffQFaqpLMQwBr
dOeeZ0iy2nYRiOxiY1+XvwnNGC2hiU6W3Np/dZnlyo+g09Tu3oYwjnSjPsAea40qr+0vfALeXWEP
dHY2vhjAVqc9OzvSS3n9OkDrnI7tTdSpzAqP3dn+V6P2Tzo7TjdvzH+MtFyuUH4uXBl2kDRXqh9p
COHv4GmQoTG9bRGvwLjb5OrsGo9OdsHlDcYZvx5BC1Acc0SZXK+phfmv72dnawAOJEqlPyu42CIE
ADqXBQSZJ20G5wRwsfj6buEB0SkdO1HQg8dy5PazMCaZgp8lqTiakJvjOoRpolmW3sHzBh57mvvj
EJ135I9rhT+P4zN5mGYUBZFAhZR1eauc+GCM/zNg/hGcMlO7A6c/Av8tcAQL3X6l4AnH+FqtN+gY
h04/bNnCgYBsRuzM3PeBiMSuDR+CGBDNHbuU3Zh4Bb6QGczj3kCpJPGYpvmY16jfsXzWOTBxZpNv
AUrhB7tAF4i6gC21MafS+VMiOROYFBIox5nBqm/vKFKximkLEw7a/QiFKq9bpkPyZcAwPQqpWuS5
4gBNBOde5jooPy58wvKAoQkBMVWG5fE7lzacCw9bwuJ8SsmesaZh/KcfF+9U51RnlyvvESrlNfpS
EePWh+j/uLP+vPY4g4U5kKr2CgG1n20uzyGSk8+gbFKBbY/rK4ZjtkhcJ0b8yUECi9VaRxK7/HVF
c0KGq1sbxNtKLSPQ7sV9yc386csfGbhli25AJ6wPgsvt8Z9TrOl3K8Cj7PotRSlQRr1JU+6kNDeO
VyI7ynTqf0vko/2GUeL8kdoKXRBtaSDL3904hqC5Q5TArp62mL4hWSvTNZnfoq7gZ3mA61yY2MnN
wKGcY2h51kZ+0rUUpnYQ+vufHu7wZU6eV8om769CfzYuSeND4R71UoYUQtz1KPrGqx+DZNymov+P
29ZuYWS2BQnS51rvchDm5iAS5+BZ4OCs41gB6gjIAlqnjP8v63cd7DLUePyMixyCxEsk16++LWsD
5Gg2Lpxhk9a3aajOR+Yhjz2PEHlVsd17g4nUcUbzi95tXAsHDSIYfPYqK5AHnfraS8lLpzqUjkg1
kBIUiyE+TItTgTqMn6rVk9uPCx5RDvRjQu4phzYcfoIWGt8tlJQ9oEViiowlCw0rEm6o0rmWGLyu
HkREqchZetTrYd7qwpIYHblnA1ZgKWAAtxKycYdLPXMnC9dQYt8o5aQ5vBb4flHZQqupQolzBg9E
2BcRGHDYO5BauzqQ92y3Mx7e6GjJ+INuUVJJPxZcrLTpOFtfvAQkia/Hkch08RsIwLSMxibykvWU
rcn/ihGMKXAPaZfZ4VkB+HNiOBpMVcdT5TfWvc1f7ttV3BOtmw+89ZcO2uI4qACY4q9QcfvZPFvZ
1LygtGTsh5Gi3wHQYaNDz7XY784r03s2HUQaOx9qfWq2y7fopKs4oR8R9FFKf3drUShDplpO6VTe
Phypr0+1NE3X3vffNNU4w8QZWKxC4dv9itqmLIP84KKE4XMFL5Q84slOmOtTHT8YNuYbyGF5CmGg
79+0KtJXc1Hfkr2K1IJ73V9pqnhxfFNzAKB/h3gtSFeLR+xWuBHpIJzK0hepjUKwK0UzpDnL7Fbi
LIrojWSCtpBj/3aoqOHrb5IrOXbxq+Cjr48V8n/RRXI0fv2u5+dllP1dyHibSx5M1g8sy350HRcQ
LuuOzIbkvnBzQEvrsfujnAJzv9xtHkcxw0QHHAgDvdoW+A9O4+ZQeYpB6vPugCYdKsSur16n8c80
cSfDySutOAFtK0BN0gTztz7r9KPJJTiyM/x0mSFQ6V2Vdv7c2klharjXA0cv4golTk9x7x2Nvuvv
YFHRhU2Z2n7aG0J2LO7j5BZbEPVgH8C0ZngGYV+Rjlpzo52+Ul8Vgcp6JuhQpgBji87I3TYrBN4Y
xFnRy18IeZKN8q3nbXmxSTww00a9Boln4Y2E4xiP7fVlLGbUkzUoJrYlrVCQt/LognbjDOoSV/0G
GKyBEvGvp0YpV4FcZPhxOeZe1JwKJGbYElPElHXilHE8K2Drw+Yf80PziMJUl1k+oWbInt+ZuHNj
cFjomo/SXzgIBk1xn0KyD9kZnChyh6/mmtZv7LzHrcxYdjkE72feqQ+uiqoYR67lIaRaqKRdyQhR
o4UKhKrev6tJYcpkn27RKDly4Qk2KGDf7qw9y8bpXuFDwiVjQUqsHIowjeBxuKngMO/0XbsL0e9z
bow+6ezjriE6rQgeBLwjypzwP8jfexI8VCI8JvAhHZoE4OkD/um/nOYoUth56/euCSQbHGWdyAZK
OQsiTCTR4Fj/8UKSxaYLAjZEjRnA+ehdudP2DgymK2iTHFqK1R3RHSvFtjNLFgnN96aXtz9tup/r
lRgVswWuBt0ZZHe9YCSn7vLKwJnkpC963dIQoi6vujD7KFEjw2PjnH+MDcOFlI/G596zs8EElEEX
d69mxLOLHHuJdb4Hv58Zi1ZFcAlu+xipLA3vidcWylTTbynPKlli+sJ1HuI9ILFmQYOKvyPik/7Q
/QS5yvbyJcM8B4WbjfiX7MAtxB5IUM0/KM4IHwRzeSAR54keBx81H7pFkc7XdVjX3mOeXNreP7Yw
dh+ZZ2GKrKwFw2nZ9iSKN+PBXmCXRfbo0Air83G/0xX9sTRtAYKq+DnCotfUyMLFLPLsq9LtC9it
dgHS5p1k8KcJalP38mBOgbxvyIXVHdHZ1viLl5CF5Q/VUMPnsZJ1uVFxfm/+7FRnNMiNPTElzvXC
4rSpdyRbV1JTn3staTDu1h8wTHFUhcyHigmMBnJ5ZdR4RRRYm3/JhHZ0ArJaN1Uv9yT0xBNvqSrw
AvET/T1LZYJbhXaClCnV8UhAdm7eiTvAbf7mZCWNnbUAT+3w7wASABeuVt2YKLe7ghqI8HjOKW8P
n/hNCE4ygQ3r7Jf1TmPuMkFL0N3P3tBczqGLKTdELvMrat7WDpThvVJr5iM0DBnQ6/0TNN23nykH
Ff2SbNkox32GvC3rP8s1RZeNZBbMqqI1Tdb3NLsiOODG9hhe6FFjr80zAA4paHao0KmKRgUN/G9S
s8X6EXCtpkBlRIG71P1o76PEpDwCD/D3UTYqxLZO1FoV1iqggksokV5u93xsOist5cZh02mkm14w
nlq5Cbx2INnQMfkvDqM4y8Vt//3h9eetok5Od8tv83yg3WpVL8M93JdXA1cIdjsw7c2cOoIAijIa
YkhX1KxoR3AA/NLHpRX7Qg6GkXbKSR0r+qYGXzFrdRRcw9bwkkyAXyWoaS5pZI7o50rWXP0R9q3M
y5054rZfiQscsNd5PxMREiQF3zxihT+i/fMX2x8g7TGs/YbhvfclO9QNB6YpTAKlPLmgkDC3nlTr
iz7SK2NqUK+7oijknIQKwNOudo6eL78IO6EPQPSiqn22/+J/GuBU7KI1pXYXViYuIZ0uxyaqvyFU
aUyeRP3/UdpGs5UOmGEVxL9jAr9KAXf+FlnRvtGXfMBZPSubyTvo2RN60EWFleKL7IUTo+fcjXcw
g7naekdS1fEWTr9/vxYKkvYJSQqEvd1mHpeqEUkxXtKj3ZnDY1hFbNLPNLxUnsCOw5tejkLf453d
xv4WIrJ/GQbJsajbGG2fBrUN4OXqKlEVPGGlFqinqK35YkTPTino6VIyNvGSFLxRbfZ8XkpksA7r
5NcC74aLoS1S44bU4WpcxFP1s3NCuU9eRDb/xm5lQqISPpCc/wUHg237dYp/1DBlSujxY9j7y7xa
qPbCF9CysYC+1sWKDcew77j+Glxy1zNIwR1KcPqg+ZqYAo3hcRyhtHtMw15QtGr9ZIFUNHFr19lt
BANd7ruptwjf3fSB9990BgsG1B2K25ykWUR4q3N99Yz4d5kLZQApVfO8gk6K72cpQBQS6pRo80/J
xmyObX2qfsv2SCguYjc1ghTeeTJMA8a69RLorWGmdcVEvcJ3lojUjrFsW+Pi0eVPeLDtk9keYrx1
mjglZ2FUaJL+01bJ9no+xtY12GUcp/xwiEZNoW23mYKgnFnvaTBkET1Nts961XRLrYbjd26VCoSb
JxQZ53SE0wZ3YtnWV5+gDVCt6C/fpUcSQdTbCqP8WTkI6rvAXfho1pen5VLrMqpFd4u+dswk997J
F+pIbCwlzCopjsYiJLTO6ZTgfKlPfTkcy6OOHKWiVlbvdgtPEhWkPVJEMEZS5ip0f3D0q+gqt5kk
cVdIVh0ZVEuw07iZFhaToRdAGIoooNM8uk2xHYqvaB4n2ccutIapY+nngY/qQdCOAk1fuIwLhkUu
OMzb8w4Ptp+dy/jSYZ2Hw3r0AtpKDy5hixvQkMTd3sygd3etqf4Sqo9Ze0QAdRiF2czSufJlHBWL
GEZjnpNbL6wg6NS8EcNmkqK/75wkZ2eb3dNaPRV9e4jWXbWHQMrNgaT7t3EvYCENkrjAxBkOn30w
FK7xue35gWpGivljrBMMTVgwYEBUTfG+/qQxZTSO/5N4eNxfRYRxxxAuAZOs6xyEvUpZtsZEtHKr
ZVDILYncTlEC2UF9r/3gS4M+DPS1pgPpAlsjw45JYA/V15RXzLKB/qargJ+Lb83cibeq+RaQJI2y
oPOsZkgVdR6oJilZBqTmyweJEX6Ir+zXow4kZDTW6CvE7WMvGuxJK8ioedWLK6qwz2MQ4ABljtIZ
L70OFgKuVaGlgbWpqvfVUw+2WelI5QeLBBVsadhUwSTvQKoFkoo6bvB3ZWj+CkbMjB+yjO9Eg31H
rjZdlo9Nt5SnV2AqUndZvz0OEGmBwFTUIMeIdZv3pQBOwBoq6YyTHQgbzoh/EHFAEFYlHk/HTYC9
yf3DlAewg2XbrRgyvRNhwcTd2o8hJ8zTUAY3X6WDsEMpaLcksoVQ2tuOzIj1oJRB1tSxXLPDtP7u
5CEl7dYLECoIuvI2lP+M1NgEmGVCT47UrJ2BQYos9oJp15FKWqGLEsNH/zRAR41q2eYEFJw6cCnq
+TmwIo0acQeykLo9OqD8OY5So/W5wLG5a1fyxBjfUT4nrTj/WXBD00QOuYOfyDFwvVL3ewTNBQRB
k7IjxUXEwqEh5D5SKpi15vuR5vKzac/Fj9QdBmq03h9UrXnRPwNcA3FBC8m0SqP5WrhIk+7xg+nj
O3iyly0WXkEt6ccmJdJ0t6jQNv39loidtkuKby8BKA42AMUrgym5J0EzLHc5sMJ/9EwX4JvXl2t3
P0E6qYPkuQ/5epXpSJtlAWsw+1IedW8C+goAmMIWzDzS6U+PoIJ06FJaC2wPjlw2s0OcW1C73AEe
VfY2rP26kG+mOcXQcBMZf9iEtdmvtC/oZnrlMxtwttomJL+ed7I0PTxRU8vv+P9IoHZF4J0j79Nm
5KnZEGbgopu0PZijK3cApaBWzmpSAPYZLRlksbM69vSfpbWzdZiZuvaBdiqMvcmIkIApGV6NcP/A
WWsm+0Rbu2yMmXsJtE8bv1L2m9EjZlHYIq7iXDbuegt5jz9YZJcph6SJWph9TLtLiChSLauepb0Y
yxVP1Gm4Ajbdputls8ZuKwVOnY/2H/+pnevPhKSi8VBahIBGlT139CAJto9V6Aoo69QkmgN8/UU8
OifxAhD/Ohs9fhCGdYpF8T4zTjPyysx4oot1oC6HemgQpAEsx5Y1MFwqbwD3RmmbtiVVMjkUmH33
6ip8LDO6y+HtKetba/cT+3EBVL+iZbHLUGjJZDPPflqHfP7gOJmhMVLXxUsgxyeiNI/RaEpDn7L8
Oo9Q6sF9pmze1TvvmnP9f+7EhE0YOiA9SH5lbzZXAajiNFGXfL+gJfvoc9cgKRYtMMbpuVv+hGnW
2lw0DhyLroXmBL25AzjrrOxRipIoJntiZk+vdv981gfyUAcs7u9ChmsgHxtWnguitkE8NEjNusoe
Ft+tscSPOQMpFPzX2obG6iesEzsT1kdCiUK0lH36larnjOUFZkCPqvXRSv6igLYxUtgoJ0MG4o5N
P165R94yMxVPK4J1XY5UXUwACEs9zZRxi9AelxL5F6DtpvMycMlFZ85aXtYgomSxahBmPvmKeUwJ
cJBkAYEi6kT/3KfzFXU6rdMA4E4W0+mwLMXmeWgxFRYXtv7iVm5AGnqJnYSigxwTQqi5OtD3Pnjc
bxHzJSyVFEgKekYO8JadiTnvEQhO54Wus6gfrnxMmJVEeAuhe9edBJqnWgHD4MYsHmqL+/jwVK1/
M4a6N0VLp3wRsABhNysP6nhrDRqENIz2LeMfH4BCjcl+N8bLpzTQvYFtrsmuQTvnuFI7YbWbCtGw
XwYmXonKlFTdiPRb3LVshtMUdSuyN8knCMfxe45DDR6gboPA/KwOm1HfbUZqVK02D97WNfURGPgp
axJT+7eYBYC66My2KE5RwO3j4osCky4hRjqTR8xkVkfZ7GqtuME38HA620X0LS6j0rO0TdcQqvAd
GgHZDBC6GWkbeg6v+NIPNrR03HPddBUOgd1cunWNsCdTKuFU8WhoS0tOox8cQMy8nRTHonubHZCn
AVFk+fE1o+NB6G1d4eUjka1DZynVnvHEXzYMLv2/axa9vTq6AIGg7aS5aR7S5xXkrTYbVHQRc9xq
usfs3lChZF2HDCTvUGdLIBHjt9MlMTMkuBVfFIez8w7A+zbyODGDv7S4impggVSpvtl3iw93uBYS
491ugE0cmC3yWN8lxeh2qeAcXq2jHGpJI5k05Jx1kt6p+BZFpf5LLLo7zhPiL3M8LhyUobxynvsy
1ZmXEuEE1GohMnCrZd7ioP3hfiJ/az90BXxOQNoS9ftJZS8ftb4/d0PqD/QHSVFlpphFBKCbpFKw
i2cH0D1AU4gR09bkvQMYQHGWeNNDZ0X2q3oSl8YO3QSjpLuAU2qUrA/53rmOFD2HDXYYJjQMaM5W
OSWhsISGUArrkxRnywZiJTW9Ftnn90Epx83cfD5+K9pZeVmAagpb7MsvhNKzUgkODvxDC0PnBApT
Aje6j9Z/BlKDA1V9Jv7D/oaUrkIBIIhTn3h5nJ/KhVGxFLhFXgXm32fvvDHzBDq6VvfpJ/WmYuZO
WOVGNgi7uK3B+LdzHuJlSfQOdw2OMhldrmWTCMehrNhx/DwhFLvbLG+TswlzQZozTuiMTwMNNrfJ
RVig8Vu2hamUrtXLEKm9RNqWACN2OZP14njbohGyHD13hKnTVKeqoLw00XzUka7Sp7T8w2htGw0v
KLi97UIyHAfxyzppDjsTiNkw10hrgmUspszWrE5hFeFkeL4aHbzGSJrSP8YxM2Aj47VFu4yK7i1S
0xrFpAHICuflDf/ASlOR3vJclbf7mmtzmwDpcHNcWxQIeI77+qj4MGDq6qtixzq8124t655awdjz
8wKGPcuZXkc40R8T0dVmzoPn23Rpgx0KboGacU/maNwRXXpf1nMZgyTw0yZd5stCwOa2+ptviz3y
0SeUbm3O3lRB5vDFkyZpr1ONveQLwaa4HuO66PXQ++OCf/VfJ6HdxJipLDDcXJfEZgRtAT38jhjH
q/QTm8WAZA8XXUxx+U98mhot3AJ43fwLvsWVXTYr316FtsZdZve+l2OrIOyUVjgKb73n6eKKc2WN
Inry4CO5sJnh4fTPYR9xWiH8zzgy0c7gZbl0j3DV+ItAwEsFEYeDuUhlfo1YwRlil0qXs53jFWN7
kMWqWH7lmTSALbwXwk/y0SQOXsfDt/6w3FmocVTInHCDdX5TC8WJ2q0t87eafGe2x4LL31j7nScF
bYyb2sHZK7D+7Q2Yl5yXrEoCpYypKkStSm2HLi9t82YbQTILVvc/za5wS2RWEmDZM7WOKQb88/3R
BY/KLGP+b5RsW6zcWrseoEsRwhkqhgUdfJUq6U5B52iVJxeevnwI8LwAkZw/blBrCA54GSMloqX0
C8wRWWM0+T0nGbZEwm201cjaLicY1Jy3jAZh1NQBUQAm4JTfAhPhpwCXS50qf5iCUhEbgPKnflHc
NhVcXZhzQw9jDl556tb+H97iqSRyVxVdZhWixKdi6Sgt9o+hQL4PuOSV3PiIAmEbo5X36DtfrVTl
lKKT7RYYxY0HiUeqzNf5K6HUSEb0JEeH695j0NdoBRaoDef1wumgU2aF2diGeOwRUzmLZ+z0K4Dd
jyMCwQUhCSLrvfJl0OxALF4Bi59JwiI/gzD6Km75P7YAAt3fWS8y/VRV1PtQ1Xy0FOjcB3VfyJ8K
AS1i4Cm+w8dOpWGEKJtG8d27aobthHDGNGA/v2LGyyLGCBScl6KlE78zb32X56v0lpgHs9a87Y+i
LNftMJTYXum9c+EAH8U5uMTazhYPqK9Wbh1LWF74FWQ3bDhsP2Y6Cw6jxqEx/YmAYByRDJ6tQ1zM
2F9QA8q4zWQZ8wi8lZ+wr5I1gfSIJWvKy5+zTN5LSpPSdlIYz0iSslkNwMN7l2QOPV76sqWOMsB3
cc0/UDeqSY3TfyLUQ+df3n+crr1eXdRIJDyousNSr0A6WPUfmqqA1t7NiCArgRJ2ISSV0kv56XDp
k5QF1PZV2D3+H5kIB/BH3qMAO/b7HgS5jyZofCRcJxlW/9g23/ipZEeM3cZVyMdGhHpH8kegKyPp
/GkhWDGFPGELPd3v2D7ERK0VXNMwilvjHdpxKalKC/63HTOiaMki32TgCR/Kit5LH3d0CztNFvaN
31BOn1G+aLqaQvJFNhenHra2gDbP4i85kav4NWfg/gD8JbCjnLtSlLnQiFFN6Z+prDA0mcDU9fW5
Sh5/9vCr/+in4tZiyz2T0QfAHPNxVpmCN/eDAz86btCQslw/xX8ugW4lCRP1wGTlBbztFxmr1Jzr
hvl/XzZ0MfP6VQEUUv5arLHdY7/hEmIxgJ2o/ZRcJyjExZRlgqXAmqWRwQ95COtKIxqgsOIwW9QA
xuD4Q3uMGC0ZzbGqqB8h9brj0GWVw3xStK2bPEdAhsSoFH65HPqHeyeRDUXZhcKvxguj0FSVa80E
iihRmftctGs/tq1zbHvVXPHkVOD+bpX1Q5QStwF/J4zoEKtJNAJPdP9tSFjqespxxJZ6qDSbBFKk
Xt70HWzWHWu3Kk5ohY4+7LOzuV9+po3P/PUtWmDkvlnnMeGuWS8iAiG3+WyN50fQVV/5kLsysAau
bzsnGJsXpfwsBVR2mUpYQJzVnD+5JMCC7jCP2p4OQKIlyS08GKiM+bXul1wAAW079yA5Ll2Y36b2
YIrhSQ1tpUAg6ZdenwVf/oMHxSIMXeE4CazRUZLEZqWi5lUKh9MpqblQZKZeU+3QlJDuzf28tuuu
7wa4lKNPEBwNa0TThfs5bggk64qZHS5I2QuqjP3uOcZXX+FOnXOJxFGQ+Flj4CGWVtUIeeXCGKat
dwjHnSR2e6LYUE4UxZlX95tVbk+Xsy2GKHK+I4x8gAAthbfCaDolf1vAsVxdBIF1KyE92kYV/Ntz
PwEZUCP0N26kxTZ6cT73uWNcXQs7bwubgny//apFzXiTCc228/cmlYBFovf5u/wsnbJWBeDp6SA2
STYkJSLGI7d6cTEVXh0xkuTx4xWRiIBh723izKL4//pniwqIw5N6KH4jr3ASpbtfEAkkhyKWyuBN
nbWyNgGPCaMRM3g9Wn7PScOqltVjMG0hKyDwDE1fC0AUZ9PpuxfDIgRp4Gy6KbXN/Neuze2Aq2PX
C+eQIsHeZFCCYE/qbVMUs6j4Q73xDT1Ryo3ZpK+XQYon1WKOlnL4pyQX9clah/zi+xskVVNWNcvB
J/xr+R8Z5nLcbCG2vMmAxbH8GZX6VGJnHQmBoucUtpNfxDXXsBJmSx1ost51eRXaJ9NIdMbtohdA
2wkMEW8qE0OxJmOPstHTZpQsZSuxHyBHdmWuZbp3dEAasQKV/sSNQ7buyiu2n6DngrhvECP+GOjp
kuaR7kr5eDaoa92PPwOOZrAtdR7VWNHCDHoD3HOYVsdWx3rkZAX3HkpWZIVwbCWhL7Oe5PFccrnS
SWEQJxMCA2/fy55kOVvkmSSy5AjTeulT71BtIzhzaP6gsl0lfCVlPVJ2IVORXAE3GFFRv6i4UFgn
6MqJgc97p0f4QwMy8tm4ew2keMV0gP4JSRWU5RtJMZjgkw2Nr+5eJr2rFAh3rTLsD5bWZV05irkQ
z3es7B56Gk/XRFhJz0D4/VF2cYx8eQoiIm9sqsSWAmRWB2bjYConHQ6yFr0EFWmX5y2kC6rWXDcE
KsWtI+U2ZU8lw3sZ2Jqud1fQ0AD5PctM/XJqkBqTTJ/toPOQmDA1R08AWI/nHBY8TP2PqxIf7q5k
DWEWTBroE8Rn/EHr/CuYRyeOHWg4QBGtxmVvYjNyWaNGhuLeAATqc44ljOAm6L1JeXbCQwJ549qc
kgt87ZteYDN20mKpXVM/7p9QP0VMwBVMK9n9XQpEUWwlpuZ1w3ZeFAhK/H12Q43rEYM8mgap7z0C
M0qUk7TIR2tC9obF3r2Ha3fN9W1KMRS9R76BENE3Ym+C5H2jrjlFBW1p+ik89ro7K3VIjEtm+OBY
/QXfUNTwlTl4QJu+9BqJDxh6i1i2gE3n0oEBr9xzKnV3hYFZ0pZLqUnh8SCZ43Js8vN/opVrq852
VOQd33U/eL6E9LOnViHx7SkGMQL5gHb5TRVdl6zcom2aczrtgdKUx9c5mVnBHoTeSBExPZJfIMSc
47RsVUeTTnreQw5KEh03swT5O2A6VOvyU2ymNkQozaUGxdyrjh39BGseb2xYZncgCc8oVkTH2X9q
Fg0Yya7AF+txVzmkt2YywVdlIC9TYo5I44UxBgitweAxwLYSqq30trw2NCiqiKzcz02UnVXohBdL
93NqqFUZX5FKPohk31eSrmV8CMo/uTv+/UncpJBhHRIf8hhmOkvb8aMAw6MA3QGYxEExRoILgobS
lDtMQxsx6NO94YseW3GtYFgMtUmYwZ1YqvOmvOhLXVg7dQdvChw+YLz5n1LPrgyS+4kGD0ncoj/9
PUN7cLHYTmDMN8AxI3Nf1pTIZjfS1KWla/BOv6SkQgEtZm91cpwPZ++QSla26xUB1z3ggkH76ysd
JEA7HfTkRhhYsnkh/NcSKhZjlgOGjnESoMnXDVIgEQNwCwKo72yK9R2QjYNGMF79Wt7/+AQx4Ops
MvOhs5ZUR9jwXDKXfGrZnAJyDPdHJDNdS9LWxMMwUktT+GLyoU7Rdbz6ygisgF8LcqIN4xhlDCUb
hTA44T14iwq8+A8kpx1pOXqv8JdU+5fGgtSBqHd8owpdRhnnUBd8RmbPWwhsZDJNPnUP8FKrYViJ
QiSfg393lg48JoKv0f9uOToHY6DQzTAdbVhc9qEOg55OpK0rqt0s8B2PwB4vApVDQYkG5BjcMiju
5nCbV5znpt82yjjLFpLh4e4MB9rK79Pt/3pKFGuiF+vTHUiNH2VERmv83Fner9DnyCHjjRTy2lMG
IfnF5RiO2HhRnr/MREPbZgGDAdmGHocDxoaSUJxfbzIfD/xJk+RL6dbdzCegQ3O0BbLLlicWj497
4GkYr+rI00Q12jPQPSkK1I9y0Sy/4H9MTqxM8yPJ5XZ35pN3eh7db3oy4/xChLRTZMONBfO8bFBF
1xAWAI5FuqJ9M4zGqQ030vTzTS//R0fOcT/39GftAt0E4siBxdPyOjJxJoK08f9/I0s9GtMfhXNu
DnkQxLsSM5XIPtmrbPyTnT8eqhCNpfOnkpKxda0cyRyFe+9sq6sJQgvjt7qq3g0+KypUV3t145Qn
Av+fNLZQRo9QuLGerVtro8WJNRcrhW17Wb9CoCDTECLBiQ5GLvjrvT/hLeCfFv3XTD88d/EzMRw1
uTwDVd7bOvPI+lQ5YrUb/8dzcwwUGWs3kgD2bnQpgD1/LVR66e5gTf9UKv1+o0fvsb/PU95fH95t
s6at154NQ11y/UXaZf1mnTQZ79qe6wBvzsMl19YmddctEstAXLbKZkJcDeq6Sr6z4/VfFdXwiJv3
cFyu9fBhWavZXn/JDRucLgQ6c8JRvMcxuhTZPnsuEJclUT5FuiiQCFIjv34tDzZmR+DbUTLFDje6
1gQTbL+8uR0wgENnC7C4DXwykPTMrkzzvpmIGFeWOVMUbvCYGB7EESC7wRUuUnZdmgVUodGzxsAA
uvbkR8IPjBS3SL04Ces8VXKqtp+va6F/lWiPR5DkoMVKPGQPg2Im2dqaQDKVQ8WqrmwiayiYkeKO
CRzeEXTtNWDAT/sEiBmC7eAXY8SWHN6XRKjdEs3g4DDGdraO3U3nOEG5CFt4Nleten5HG7hAj7zY
CNCK/MZ1734cbDHuULuXI5YpmKA0yl2sqAgA7YJSb16cZ5ugkF7WQxCF3Kz6WfMeVoa8nEHvV8LM
Au8dFxHK4uhdCpRTGLqMJjC5grHSds3Vbtdmb3ymKdXAWYlKcG6hzHAu6PS2mMqNH1FgtkagDPYl
53yiqI/12YwjrejUVcwkOe9AJq3OW4o0zXQ2s2B9bVdmRsFBCFLbk+8E4sjOu3zQgQqnb5+SS9B7
iP8zkkozoP0c8t19zmVD8wnHmPN2uvjNyG0pTHLcBZF/6nSOQ5P4SZAX2AyiJwQ0k/OL2EC7AYa3
nj03m8HSywfWfkj51Ocjofm6EWCzG2VWvfbUOkR3BXPMM8VAzq3yU3x4jnYDc27bLOsJhMdlldjG
2+jzrTmr/ZjBEk5MRJfrF1N4N4Zm6r2WnqjVd5Dwi0+hk1SG8+/bVaY6kpJIo187YalxYrQed7U6
VLcWTYMsRY/bwTZIdcVlMzT697/KZbiQpxOULnsFe+v4K+/YBv+oApMgvCsou2A+PZn7/a5hYDm2
U2RB5ZRZrL9h4071MiZLgNjACeh1veDbx4DpcxpvyNLFJGd8UkwWMooBw2aVSVURmKi7QDGuSLYP
zAFs2uVSzuSVM1UjDdd//Fw/ZBTA5PxYM9be0NGLoYoV9uEGUJaiT9p3tf7LtKqoEXdVnD/Dr/Dl
pVZSJ/tOVFovU1YBv+qyud5+5W46n3hMg5RBzmmlRm7x8qdsiu9bKtLeibcBkvTQrHS+OR0FRM8+
YSRCcgUgFzB79Ue/wYUv7eRDbDpeyGOe6EYaWUpBLujZY4JGSF1Zy/eIkZjUevuJo+f4Q3tqoLcw
71zjbOVLTfuEkdrYV+z+QZis8sJCCF3oASx+YLULDmnO+FZoLgdGrQv8x6kbkcruWyy6Y2ScHgLI
W1PFUEmLDo7zl3Z2JDj0NJhdBwtG04YEysXZNtiOezjboOz2zU+q6F711VE884IMAkzh29sj3yGx
qHWz6g1/KaXyoF/w83BXKZ9f6ht+paldVOmQGgF7Nkp0vwxbKZpe1xSB9KHyKVx6Liq3atSDDuRX
l8uJ7/rpDxpwiIOb6gnOsfDBQECVqcZWVWFtaDGz72OMt1epdilRj610T4/1bCCPnikOOXU0IHE5
xwfvonW5BMp8RG1Jynq32R9001t/tUyn8Qr05m3UGnNmFTMJ+/iSEN98NCQ0Cf4D1gvGXmK6axWJ
0v56P4gZPGhiktwT0IqCug1PVwYd6Rh0s4JhiUsnczPKkYM9j+bX0oWZbcbgY2ta3Rw3NhJVdkQv
ASV4Bo34F/FrNoQwXUWF/2vSc/AXLVhxZcCbO3AWoTsgc5DgTTZMvX4vq2svfThzyQfYLWJK9URD
RfEFktn3xVpCbWdqWXavf/A9a+++VZqusYZkgk+iOBz9XldtCI5VSBwj2OppolIXIgMmdcdnp2If
96LjfLmHGsjX18/mdzyIrCYuAPT8OEhzdXgdkHSqvlUsLx+Eak4GRH9CFdt3Gj3HfGC3lh1+Jq6o
hncgtElO8J9uIa+/2VRSVMWIS6VV0QI=
`pragma protect end_protected

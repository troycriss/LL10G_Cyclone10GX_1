`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
r2oopAxY5qunYQvMZ1f9ume1Cp937C1n+MEY5+JuoH449ExEEv0uTzJ14xGRdhEv
5x5Qcs3xUSwDMOXmBMWrCtOpy6WcFKrsxBProXIas6sn0Jcgi8fGMOSHDPEOhRMY
XloxDNqjuRjxdbVbLEg4hruUy74cd+9+aGFFPc0TcGg=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 91152), data_block
rpfk7eGmD8mp19xmA8xcQdDoFaqbW3xOby6Mpbet1IQ54ZgEhxRH502IdPI+9H7O
qkQvd/chcpJPuK8Okjuzeef0DjjJOFbUfXZohKGIHMxB5XCtDW1yIEVtxZ7RXsqu
P68bnxCO0vfVvxiLZGsHRAGg4/UxB7D5/y30Z2EDvD/nnIx+NzZ89QMpfCPBUmBT
Zvgn8+zyDRMh772luPLpUxHl5Y1/GX3KcLAkhSqdimQPxTWk10hhxxJ6fe5MsZNu
uNJIMbd1tG8VrwuYNy1RDRYiMUFsfs6nji3mcROjzik6ExmUOkEEsBTVf+rQ9bHZ
fi+VnseEuKSDiaGsqHBu1n7K8hMaw7FWNv6e4hE/3pBp8qjxb6wNujUVVbfhCqFw
kSqiM/VWhVF1mc7f6TFAKrgBP7Tn72JY3lj8RT/C7+oa+e1MU41U7xycnhu2OWc3
cwxaoGcP2FHFubRc/Rk41JxShh8J1ORFkwSBonvufFG1l8cfPiPrKINJGzbQcgMd
Xr0Q9vhsEt1sllZ4AOSviLxpaOGXYx/Unhyqvy4zvNk8SiuJZgg/ZG/zbNpvBZTn
DDiOTdIUlYzQ6I31XlVXYU5KWAdvYI4eRm65JqpFYFC51bzsd8vQd9BCgOldFoDk
kEt569MyJgllDt0U7fYUrtkwFLHe6i9A6cB2I122sRkGyOpmU+HjqDr299LdKir8
ad4B44NseJPCUq3x6Z7rDDcDaZqMN3Njg95oFBOKn50XHM/wSIoCNHHCpWFv0EUh
BGg04xrabqWkkxEuqkpchkxa1lYeTuVayrbZ5rN9X9IugP+99cNew2OD8wH8kvMQ
6E99KSTyZFct3WioN+PymoD0XRclcBaKHD/sceY0guGorV3+H0M1V4JC+sDO6OWi
AlvchuCEG3RRL2g4eRgMkVlM+ZXDwObLl4Jl5tlGlEYpBX7W8Hw35iSXyAA7zC/R
irUhNwJ/AekUgM9SjN9R1Ih9GBr7kze1BHQjnPAkMOQs4+sAHgaKSJ7mY9KxOYTc
K3BdAmo/bMjU3FTlpHPkYXr1yMExoZkkhh4ncDUphFijxMlu2p3HEUmkM3qPvQkv
4khaMduUV7Fbp8+iFnvaTM6DfoaUUx7K/LmPs65Vv+ETx0CTuR35SWRhD5+Db2lJ
oZkLT6ZXUOQKIGgv/jS+UmpPB7ZSkp+aVhtNtpG54UIwAZejUGAYy7pL2DineEiT
AHpu4g2PmQk+/EhDGWTW4ikoZ7TrfkiTIhkHAAFJhNaAqLu54ztS/6/6PvL/s2i1
eiJgKdN1xMDRY4UEM0O6ETDmj2kDNzuH3xZN3K/kNNR7rqFvM1aW6Wq/cWpQ72kA
iTUNbIYtmPc60a2B/A4MWp2CFHGDFI7D9LFaXTz54cdaoK1eAq7bUEQ2nv8pL0WA
s+sd8vJwWtv1PdJcMMY8u0sPwu//0tQhpYpMy0SXAQdv5vRH04YJTAKR1x+8jZRq
CtDyolORY0jeQVhiUeH+0ZBgIfArpYHXWg6duIfwGHNF1cqfaAhgXrBcYSOPllPs
3kvnZHUCfGUWA5hstHa335tVfsUiTwEuGmT9/6diWRJNzW2WtXMbY/6UON/KZ+B5
HZpr2gjvYo31cMYNUsi4qAkoyNVNPc8Pzy+DNpPSJnjfBK6vHsqLdZyUyKRLudEZ
qKAsVGb0N6ViD6Syv+AnHC8HAecO7zNpuqjkKYY/88ZJK35UDgLmAKheOhgcyYFt
WxrTjDOi+n0alTWg8s6M8vC8Xon1FeANfxpr5ZoilfC5zmGCwOI0e+5gJTcyHKPp
diqI6EEZAydPx1SG4PufOxa/5ZXpifTKunKMzRulmAB2zS8R7Nq9dyLgUBO43KtE
DXQW4I67wDeE3DAkghEvx401siQU9qB+TVkpcp3R81WN6jTc4F4bQunLwFAcb1Z4
lI14wkuiYcKELP4fAgxcgCI9ORCWmUkjqiVNa8tEQMEP8LRg0BS5KPEYNCo3PT5y
E4W7Bj5wJju1viczGGcuWx8WoZRxSpU3h2BPbqu+hIZz8N2B4tpYiV9hg8kfDtyp
RMVgmNDKwfP5qPV52IDDqb5lqZVrjFnZFej0yrAu+eFx2CzULfCRnwwLsRDgbHBO
HXgb104t2OVluzCGQpn+x0NrP1dtIhAs+XpwnFXgAhj4VTyo0yIKjuUqK5UlNgzb
b+Jpju8G0XpGWYO95PAFx2c09nWsIVseMieXTi73gQoPdTWwwUjEq8WW6VjcogMN
cBwNae8YjFvzcdhYRK2KU64w9A5Idoc7HSZq/bXGLmLQJeRSG+NO/GzoPMiYxWBk
olnys9DBXRxx++ZOjVIMwPdmcuuB5tHRqVqg1Fer7PdPfA74COzNadO5qGUpv3tu
3ywL6qYgwB0xT8lJqn/32Lbd1LiZ5D2pIvei6GKnMTo+8yRoVZiVigTmQ6udQiL6
IiENV40C03VwRVt04rsroc4wHrRk9gax/rFh275+7izFebvo4c9xR2xJNssdfbLX
ePJ/XkeBKAaFIGJ7+1nf9srRxZyK/NDiCXvIDjV1xJDrJD/90PLyK6FoEHx3o3p4
Zu56kPoVrrWk9muuZc4G2PW5/ohMcziA6zspdceyny5n/zT1XVMm19pCvCGpKSgq
nY+pAWaIKm9wryUj/GzzPXp/tB560/MNElJilDfhE4l8n2hPfwN/a67dZIAvY2/3
0kV0kCxjIYg0BP3WSt3BqJlBhVMSSqzaP/ynTMxmmkUmXw+SFwd+lUhyINIsbr1f
AiFavJfvOaD3uTp2+JKJ0Fi22DOdwfm2gNVhPY4XJ2u2/XRalO0F27QuZQZSbelC
Wu2GXufCiJbewHZiYhfAtMg/BNm0UXkJKyLtokZQM3PuFF9HNbLK9BC7k+c8MY1o
0q2eizIscpo6TFDXGLjt++rqM0T7Z9uuxk9C8LVQNt8OArNZ7L+5KXTgNfE2AwRI
6ZHXmr2UwJkIGC20LclaEC6cYgWHpJcwvklZn2X5lRrn33NJXl4CN9A1THLMq6Ox
6g8GwVXoKrXjmnMFXJg10VB5B9yA8laIhzNUJyaeSzWjfnBQ7JCFjgZbvph7yQAS
ppUmhodGKtOWpizVX9lXvMfqpmYO42TmCXpNE3ne5umoObOL36up78L0SNsctX3h
Re6ins++lq/UH5xJbuinb4uJN5g2X0AefbkQfm+DAnDq8ldd0eYCItvMWv4mv+Ue
G9lAtYhTtFYET4BdejcOGEv+ljU1vJNoir98+dls+AYvJQOcQf9GqsgP24kF+dt2
4dGpRMf/yqZlf6hkjZ7XVC14swAWPzA+zBo3HS6esI2fW9Y3qYQBoDKepK1bqGVN
SbOZiZo+6LJVromtPyk7uZuOZ4Q4HFvdG5X+3fC4plMXm2DndpZoEsilacY7ejN7
NSN5CYCi+POvJdXplce2nc40GQs5egFPS+1rHjwkRnwP8gXlvdfnmk2Vh8cd9hJj
xq9orae2msysc3sCOTpMVqjrUkJXlRGugZm7LPCObBCyD3SrYqNMGr5gxKAAysgX
dx/eTl7RuOnS+w610hivEbyISTfAxONo64C0kLlZldj0I5NaT2qxpP9LcrsfDbTU
3dKtrzjP+Nrhdwt5EZ8heBQlbWnlN203vxJX8yCrK4/Wh4n/jG7CXRKxSORO0fnV
6Wg0zYvfVNHa3Q0tJDbhnfj25cmYCGm60sP+x9PpVVFensjlkU63MPj5ksBXdNvb
0CySfMJ+7Qkr64qzxs3376ksBh08DwUZu7/rVk5Xh+HgJnv4jzzZOI99DXLlRc/6
81r34aBLx3TJI+o2StrZCxbP4k+olv7eKzMQCClz+gVDDF2gFFtu9hPIWUSdKxZz
bfig5YVGhpgmqk37ktyXbAsMgH/bX2eCc6ngkLI2UmYPiqvcTc/8UrByvmRloX1G
+FKKo/AjH4ofJMDoSRelV1z3bpTO7In4lO+lUhtr3AulyKZ0E9QQ966rRZU1aXZU
aun2mYfJi9mg8gueU86t1eStNUDmEtxKhIjMEjwSRa3BzxW4zuzGOz9ShacOp9OZ
+tUXtrx0eGjzqBgiIup3zCkqMCUfmwCMWzsfm2Q2wm66PvP2xKuXk7MBb3lwLevS
ksWZSO26lcuScQiCnLG2oZ/zgqEuoMFMoYG0YhMlC9Hc7Q6G3Yqo1VKOcgfbetFy
gWAmcYlT2zzcd3ABKpz81zsgINUPU+yvHP1YP/EKBnFc0s0FOv/lkWLwEsyGH9nD
IWhe4rpELTomkkNIxLld0HAevMuUPbUVwAKYPO7MTEh6O10MGqYby2IT+H2TvH1B
9777U/OGkEPCHHaGdGWWsc+cqjlygiR+7hR41H7nPiwFVgeN4Kwdkn7UcaU+tcvW
OsFiyYbZE3QfoiOgc+RhP2D5GAoo5LUMwUO8R5W5kw9eEMCRyoEpsosmlJRIIAC4
pMD36MhejJmyjLHGLeJc9fpzU4PPWcpoWGWBmc6wJgxDMP5Ai0rTtPTljRRk81ry
W32Sf+k/xEpY6c94ey++0CXOekBiPvdjNRP7n/jEehPLCifISIHgzmiwr0FgrUAx
mce6RKh6glFPmuVB6l4MD3kadeS/lPLQn+KmjGBglVDcXgcWrLBtHMMqav1N8t7Y
uMuLxEveMm/EZfhfbPATmUzw2W8lvGM0etUFRMntMaMcVULMNA8Am6FwThzkRUV7
f9dGynzJBK4XesKtFmI70rIZRDPyIBSYyYDEse/OpZdlj3fIIHghChe8KeY77cLF
w6f4CZRG5HyuNrrbU3+Mx/8IMg4QgMz/LMbU9FU6+7sDWrx6Ln3BwJr4IDcwIaiw
3N8wZGfipS2GTdVqIxDxmuhJz4yIgnX6MjQiUit0F0qn//IgA1G+PSfIWyFsZ3zT
CaqAiLkL8wuLK+UF01hx0Wmp/HDrBVcj1aVUMbuKmlhPimvi6F8IC0B4b6IPl1Nu
VFZ90fgQ1ekcyX8y4Gki2DKRjE3Ta8ooK645RovNfyhpAMTEdJAIKOvCfLSrFHjv
buBLad4pIVeVHfUnYxDCc+140CyjcAq0kWU2e1KujJjZsCxZW7FnDYFpzL6gU2SN
r+nwpPg8EbFjrnkQ4D2rrh/XnWXMvp8vOaIiUbqItoktuOCtPE7sNSoJoIOtAS/t
QqC3GxkouA1dTu8GB9ITzqTAH9dn5Q2Rzy5My0ZuhaNIkf+b1kcsqdKaSQ5NV2W0
TB4PLmvLrwwZk7P8lOQWgc17eYIxzKf+Qfv1H7VefGb5f3Xz+3CTKQqShm8/FyKj
C1mwQwVNmSl1wHbsp5JqGtqaamRQC+YyI0Gu6e8Ga26kpTj3QII6OiWX/l86qcwZ
dsJwZHDNdC+ht1W/R0QIOvQ6pKfQCP35Z33/j2EvEr/g4UeGGrs+oZl0n/cgYeck
6aVFrWzOpap0Fwe368WxjxS6qUkMKYIUK9r/07R8rAGQAohZODIIR6s+vW2ulc3C
1VfHGOCr+HXaf/SCCM4ILdz+DSZzR7pL1Wdllf6CvZLpgDOTTfLIImISKJlN2s4T
1IN4V/9a61JeW+qe1oIt7OvE5CDS2XtpzHnR/g5URqLWblQRtTSvTfuEA5xtegAe
w7Hp75tsPQrMEOnYtNCkhQ2feOWGEQTxX2mMA4QWMwjHzMZttw3lZsO7GhGXZUr+
q27cwm+dNXpNWboCz/NbcrvWRMWpwA4UA/h2j8IJERGKy+rPh47QposMZb6ULym/
tbsK6UbZ0qKZCZvmaz3glggyoSFfVm20Cg4me965LIuieo9YYXAhnDCOwZIk+3Fv
u3ZBu4UgS7Gw4g+PTXLRs/YRiHXtV8SOkLBNK2ElzWLh/hgXhd+ywZMmOae2uGcG
IabKBOhWe0wMsEp5GhAjgg7ZRYG4VmhE51+kS2sDXi2MJzZABOf4htW4R0OfZFr1
beaOdSzr3J9Yowd8EbEPWNy7nY6bSdnCQEWHH/WhFnbX09nSgzIMLKvCf2FuHwz+
s3RHgOgNBHD4D6OrmzCB92+ZBsNCwe7Q7YgPXfJw50LzcHEbjTiZYHs8k/1tBZUK
EummGgucDAQntWt1Kfs0AObAr25hfjLli73mQppmLDbBCKXibucXLLVH/xrI8HgL
pD+71I07nLehuq109C/yulE+56kQfETzQfDmmBed9yJqVS5lHGmwgyoJQzNgFfW8
FkTBZqlTR60S1W8QwXl/xMyEkyZTJxGiKXNrdX3eXU9/unvvEYYJ8v785absJM2X
KtFzAewFE50JUS6ioT8jEWhj7kJ5SgSuGATs3CsX4naEVj+nfwppWkWG7p+KlE5h
aNK0RftFsHkbqn7DVGVzXTfiGcNsDvnALQExh36QZKv+3ZCDo9rFTvvUw1lXmiLE
F0seCHoLbf8v7AzYD+706PSoK9HYbLb6bxqNlU7y+O3qW2SSdmEb6cYHhvOjDapw
yE03qSZT001DpDb56qiiH5EfoaLqH2fUenGmCpsRV9e/VEsuLCuZeiUhNRwsJJmw
OkWofKbbxApiQhXaxz0HYLftkF1mp0QTwAwqvNayL+ItgXqiz0RKM5h5uopPyimY
tZrXjNxZRN0gRpKY/N+sgVl8xc65qSO9OvAzYHA16MocS76muG6lq0IkraYWiqJ5
MLhnXLkn7Lk4N1UhrJ8XLdOW1aMvrBjV+8A5dMupQ925fN0KpKxRrsUzf0ApbyEp
iTXwP6Y5rWqzuwAT+lDjFIZwOeGM5wJeUmdUyR9+AVnsoRFRzAARLmSgGFTrAlNt
P7w47UhpPbOBwIPpvGFBeS1VJu6Tfbh7P32pYH04r7jQjpxAvioBlSKevmWYTUXm
hW/96O8TWPW3NH7mA70zwhz5oGSFeYNzkBy0eFEY/y+B6e9vxmV56id2lDVWdeeV
l2PSzfC7e33/DnKIgs2G+COwEMKHpJHxYCwHW7dfb4LwdV3EQqj9oqqzv0JKwO2y
Xt2Z481wCkEH0YIzU/1intR7cT1/dKwPZ56kRRaUwZNp6Jzvj0lzsdvZz821ERlx
ue8nSfI5t1v3yKZ+Sf3OSkaINedZbyv3eu31KIy08d9pdI7hqy+xQtJ6xrydVAqV
/ttuZsC1zZKQVANDHizFWD+mQ2nRiO149H4+YiqtwFgBQUvUgZ5wZyPtqM6vnud5
38lnlJ1Q7FjdxmeLexpjEPwkvY1LhIusvW4d7qioT0jLsws4z0RdRB7cYSWmqUfR
jy2EeO9xO7afGqS+F1NXLsHXlOKDQa9mD3q3vlNcdciAtOUNcorvPzD7aowK0P8y
PZ2cHelVCGOwe7tKKfpQ+4nNc6KLARxCdbx3pC1cmo4M6iTcJFW0+MKjmTszRLzD
011kuus4OM3nkuQr2YE2bECrmIzXtNA42Zamxh0x0dY84I5I5/5jGUdk0Kjskv4J
B8ndH9n3JN4UeaHj8OGvn08eOWxs7rfcdUda7CGeH/ddK6eBxUSpm+uFj3V7OqMf
0No/d7Th+EAmYpOWn6FQ/IqOzPyhvQ3q4lDpSIL57MPgcNYvZW1VGubvHmjZ3qfJ
n9W55ZFF2HxkDlRwZv9wqBn85Jcfdn8DMx5ebfuI9vdfWoi+hQDBbVXvq7qQrmTD
3ln8ctjtp8erZAG31wY5LoYRVNwnwcaTtQOrPyYLMFfiBJRwDwVN1h8sBnK4jgug
PHuxJkHE372x35HfMdm83ZV+1rFwAi1cDBKPE86Zs3rUwBvzJrLq3Gy7n8Fg3lw4
+X0XtWgPbvOJBTYAzSezA3tSFnYpkVJs281QZ+PN7FqARjunS8oAokEGFHdqQ3dS
rmd0rWnAlZMm0U5u9zB6vH7nSZwngVQfwYqoOLKOZS/CFJ6+Ha5mTA3pvL3ZluRJ
7qMr6PPv0EwpMmGOTzXHfvfuukgevrY5UnXl3YluhmjPWHN9D3xVRF6cdhyPR17W
YdafOmLE3i4LHhOSTaaZjaixSxPqARLkJQGWr599Yr/SfaOdrz+DR11KV9s0gZgX
aDF08GYLl1+u8YUHaO5A1JNA35agRlWPfXLarX0YoNkUIY6jrlYwRPSAJJbe0h5a
2H3A6Ob76BS6H5Jg7Fv/9B/GxhqV7YSEElOly5kjahSVmL5Nsjenh3ZaRCDDREB9
nVLQpfR05lxeDdfaZQqZYmPQ5jmFQaV/kUb+34L9s+5KDBE8HLuY63W4uysz5PxI
bzKx3VX+i8QxbwAtx1rZh98XqGCEv5ukBLkuUEfcUJV8JoRpkkAefHUdMTWaqrva
uBD0ry3b+Xs5NhvI1upzT/numFtAo/Cd/Rn0hblT/NW7Zjw7pGUWvd+Y642wwGxa
dtqoFb6Toj1n3uMPRj5L8tw0JfcEkBg/Mu8vepbMOacwkenSxwCirXifc52zBrBF
BgAqMwD1AitW4GGjhAXRA0OHQem3iras/wrI5bweIWlQeJ83XjyM67TazrJ5tnJL
rM1FrqQ6eOZUbWRK2qIn6LLchfF5N/GUlqPv6R/7ag7aFlGkUoUCJhls2stnPNxd
5NBQzj+7fuZVor8jyrMWI5WUB1M9fPbmRJ9dtlXuKd2ezGPD0lRyfLeAJuBsJByH
ZuA+5PYIvHzoqDQDA1D++q+lxnvFSEL9J7l85e9K+a4WnqaqjMfR3iHTLgspWspD
NS3Iksn3OC2IuhGhqcmGM+485WKW7VfBq/PWXeKChom6ktyHEn8te/0ZRUZsoBBR
pcyBVjK6rraG+xEe+VVK4aXpVnm/Cl17f63pcuqG9SCSdUFnMr0H0SGvYFz+pqtt
acrI+YykALsYuJ+V4Ks9XzgxLQi147UsH3nvHsowDjagtPF47GBbYaEa2TpyFhNO
w/04tNSQMnuJ2Kbf6Di07V3nnQKPhsdrOA/5/Q6lHbAP9pAtTHMatDawG6Ux7F34
7mFGeTeNUfBck4HJebre++WPsnjDbUkQmeODgpe1X643eX/r4urp7UxJoN6JuZeb
NPEvF+lqUePD2n/S3BxJduLjnC0g3fkJgplMfDcl3N85IdA4zShxJhUFvqtdkrgS
TMajvQ4kzkMKTRl2LjQv/bbbdqOeM/blRCQN99M5A8dNo/uxfwdVbgIkTgoBifN8
jPiv5ExJsZKQUp+3nCn5dltWZsWi0vGZr4ZiIrGm2pJEzusCpuoVijDIL6N0r9R2
wsnKR+18iJJINQLemrMkm1dr7RW+KG3A8jQancqPYFJ981lutyl98rDjooPAb1dG
PursPkRm1B+tdW6cf/5ImM0OFuZ06gkRkytsoAaI2JMQbuHzv1F+WsDVVgjNtalN
/zx/DroIRMwNuk1XItvtR0y/uO1TFqr53jX1zJ3+Oud6uMzyjj9WRSBg7jyvJT9a
3Or+o3MXv4ClARZwh44vHPveivZ0CbPki/mw5nooEj1ST3wwQaUh/Fltz6msfC9Z
9pyRMYCqa6V7ppe+vGQyxNfFDFQMdSCqoUk7W2DS2fP4FMIsYLuH5OYkegMHIa9J
cK01AJuuWZvjQYidVOteT4PQAiKd5gKMUN5PvJfBIFtYUWNbe5YD0iPWzOrF3ZXx
U+0OOB1/3+N0ny7uxwRyflAt9aZBtQsse9pbNr8RmUFJMDlsOmNUH6ExWhSg6zW1
6Qxyk+c5QychheMe7zD1b/FNGO7ZmAratO6fUhBOrZweovjeLxyot3oJh7oYUFq+
kKwHW7bZBIssGHfoIVlSGcyzpRfuJWgUnWbufkLgsASe2A7QrlV0XlUzbN23U+Vz
PJqvww20FA1cQd1UhwCtKV9GGaujuioOOPWcTlKH8aPNeliMZYSBF/5Q/uuk/MWV
yFeqURxalbd22F5pU5OaDVig3v8v73jdsiDElJKzBuKhA/B36BCsn+un3ZmJoVD4
+nCZ7/Pm5rBMW+/u9ENSOTzrzbs3bl4xC1oovYymsNPwUvfRBNIf6ArG8eFz5ruz
q6uzMs3CNG+B+AWMmHoCvTI/s+ROM+bMzF5htwHRyGnE6yC6C7il13xU0vUh+Ej6
Wf3BBryDGlXW52AU/wGgQpbje6ns70a+f0c7YFiHLm6EW7hBfv5hgf/m81BAzoOQ
r906OYCQmJZNJZ9xTJY+wqxxujW7I9OhodZUEFHAIupcOt54d64niufkMhjIFCa/
Q26jIqH4amJ2Pj9Van+ru9A/iuqOTEub1CILFpeRKE4N21xjtMTbE8OYGS8NpMO5
tPRU1tQWZ3Hc3j9Ihvr29TK1W4H9O2PsfMBM3k51YC1Nz2jkzUX1CvzKmW8iRhAV
YOrgWjmOgBam9HDnT2QRoABlByjFUvo9wjFSIWf+uzYq5fIKC20VcM1H8MqH1Edg
VERIkfu2cXA+3nBLIJ7Y09klV9WCzSURf6N+cyNCsc3W1TYzMleh0XfuIOmACqLx
yRI15As7SYKNcvGsaKEy/pGGxUiyGwd/UUQeOKTOVARstG36/vR/7+41rz9rW8Nt
xuFseSV4vUSdDIcrq+d+TpIZpdYGVRbXD+zR7kJS8eC/FOWG8+WRCGJSX5YP4Wez
fmE0KHr8GLra6St4oFG4GmZof0aTqSdfkJayU4xPZwmM9kaFQJmSYX3/NVeuBXq4
+Am6ooQL2Abd7NzAHNg25GAtC1CgG8p/j/T4uOsR8sVB7ZTEeXe3hSF/eVUAu/56
f4jb6Agg/5L+kOI47JW+vmrTPExd5wkwUAbDqfdfotGaOH8FYURtu3wQ/2Mxj0mM
hDg1s7xDJuCpKoRwUaRWOWARMOcwFrI7FjFrUxs7Ipl9L4DVss6yLEu3za3yafli
JJkXcWDr6LOcZHurU72FktSxpQMfJDT1gqihTBqeD4CKgu6lwryFFAHW9VkazdBs
znedy96NGZj+RATC2ff1vT/jQhAEFSXtpGXHiXDP8bRGbRbicqijDRW0nam9aU3T
z3Xzt5T/c4vKL2b/W68rsY0eM9nEtWGbBb/g4xbh1/jUcu4ZYloMKCLrMTYX2/TR
jlTKGUsaZTHuKKcWgqemYLcPoYgnKL9zEOcTTpsgMWkELpTD44qJWG0jtL7Fb4Zw
NyhJmrm0ePg188dn0XC3Lgb9KPcr615gOGmvu0QK8gHs5/pi/NyEXaQVjj13ER0R
0gOJC/v+IkmoYfp/1AqYycuprUCyBHgowkatpTHI3Nxs5bwmlEpFqfEhIt86zs9k
umnxOO7Fnjni6Ic7e358jZfpn+RFG3Mb3DhIRWlSpl9Jz55uCBDQLFupS4BZ5Br4
cDbf8/s32a7dQQBHPJY6j7mCpqD0hhofnvzTy9BaI19ONIgrtPkqSca7HN0fkF9E
cPDjLEsF0UxJCr7mPaY3YN4wg24oq8cTGzo7GRlviO8mpHlV74xHyC8HT/VoZ+SB
kBmrnRKLjTpbsoNec0c6Ayj/FnDhUA9XydtcvF6zTzrp6VFuHIxStdfLEhg5Mjyv
Qe6ZP7664rdRQb1ys/yMH9ktN8F5lz+WB0/HJLPHC8qhwMTa0E735HgpauIYPBBX
RBxXxlpxAlErHOxzHBRpZctFUTpKWmECKqensY8nDqerEpwSh5CGOgF7h6W103tr
u1dyJdWeFhCdWnuOnRtVsU699WDPqbsom9NMTvi46xTYgaDS+N7oVGwtmRgywbJ7
I2kTLp4LHPvD0ZNHg1hHP2DKc1AeTgRuozyMfoAYC9Um4ZBC51YxjIBV8hiSZY5P
Fvz1Q2X3/uaaURbufvc2tAqXMBwAxHaGdnjZi9elpBrcLBC2WB+orPpIDqv0pTZf
7i2wjDZvr4Bs07942hz7GSsjHTAMK4qt4p9yRpjZA2x0Nx1jQBiglQkVMrMKtq35
O8af+t0w8JpK602GZSd2zy7AZSGQUp+aaYNBYwEb1kTvTB6Vbhbn5tP9uGUyQsdL
GMstCrby/0604j3uFXIXserpnRHj4A8o785rtBoZ2Dbo+L3guJ83rHXNrKMkT+FH
j/5ZMJGGLYKNmkJpCVWM+Pat0YkBqGJl1sBRuO2rh31HwbBBnElhzNtgL+YwbPtF
U7hS7lcv4qx3WAzHQzLJpvMxqHbypVEd3Djd0+8BrFctROVNnJGS2t2u/X9AGkzB
TyUDYxZrSCWnpz+WL/1zL+MKWj1EJa8VcRKSwwnMZf5+I0t93E4Myd6Z29lLsSYW
HNq8YWC8i1E86H6Lt/jNzg5QFV147EmE/qIpZsCdfhBS/rpGJPfRwWqv4ZhEr+sP
RoJHC4tHswmCihQcmI7G+7jsN0uNTPlBbxp7Ad8zXULm44i3t+u0n/9wcRbM3Pic
jieVZkh5Xo/tvxHtzKYZjtZZaf4Bg3DoL8G+Nnq11Wbjf9/CPwr/USydlm5YueLU
3dYC0U8VZ1H6wH070iu7wyy7KBBMnO84Jp/Wq6/pKDtLi2jb4yUYN42zVXzs8PTh
/uTs/gxoB7c4P09Gh+tzZNHguOqhKRr88OiSlsHqtzgBVtcHe+PKqGDvIb6AFht4
84OzD7toXvYUeAT7fqp0VyCg8aRkqjv8YWBSwxNJRSELIOkdbTPyrKysF+4+Pk40
4XoT5mtntrfGWfttQtUta+9QsitZMdXkkPJ69nQDsGbKB0owCKLmFUd712UCsgW/
AgluyT1S3fJ+FhX+vMCQMrR3g/MRe8jdMArU3mNqUCB1kkVTnfljKkSFyMw5Az+u
0nU0a9oYcCKg5nbSxilT1Uz/b558nQwhKYyYCqbfg8X4fvt3aCkS0RyzxOL32jT1
shbDf07k4fgeIqvVvb5YkPhpFbOTvPMoY6IKnxaEP7ecMKQmwxPBQlM56lxgJ4vf
vO7nuJ+2/IQ5XCKHJJhzj27vdUtXG+ZsAEuzPFa4r9Wj3IdSyykYfSc1fvFe9SUM
tLTQTF/Xm4Md7I5X4lkEnhJcRtKkdECSqC/eWl70+eb3TcQo48yFcuzcAWSis4/R
sRmQeHZTcclPUhStVu6w38vqycRg7PvHr92IYxczxTkrO+YLe1QwxEsePKs4R46F
giZEZD7bceE+9L0hmOXMeHGTcmH6vDnMHg3g0hDBQnSF+PbiGZNA//QuszVc3BoG
Ouj1uHjfQMbo1wMeIivbV8w0fbOvGTwRrKqIIXy2/PxuhmezCeo0iXbGfqM6HZjG
k73K6MnvQQqaEz26ZqUqD45LEEbtVh+uSKFqLWQP7rIHa94ZWhXKu4/UBmaHtJY2
24lPQ55KO9VMlAFU4P7Mz+/VsRIEH94cy8dYgga4qUZPn3M/3ctPr5to1lQ0P4v8
kMU/dYU4mLza7dLeqoIxsBNPb5yI9xZ2kxVvyN/Bf7qMF68TOys5LBbphQbcY/eE
mUphNDgDv9YZOKaxUhkK1JmtCYjJrRna9GEwddVIuB5wFo5t2aEpMyJd3QBKwgtu
PtP2HECsZTO8G23rrb9ckFCyf6IKms6dhg9s93LY8N4urIBkqnJ7i0zrEIVJerWI
XK9eDuDnUbWcOX8CQwLrMBHwsxjD2qmWczpolyZdUi1q5bgmD522OjHyWszkygfk
fYny0qZQhRo1F9A8P8syWajgQZMkumTdtQ1r6Q3SnMacvkKoPa4NjklQl+3POh5F
AGVbamUyYkNQNrffr6J4M0kbCaoTtroz3lqe99tGx+CScofKuckeUmYiS9wrXf92
NdR+uVqFbBpW1y5ybZjIgXuCkkzxTvRBg48QlCFdEkj24GqKnQavNmZsB/mcBIeP
9O35sZMcOnqDexT18vKB8Hl54us7aFj/+O0oBaCZ8wL1gLASZhRhNXXHEnnMaCyf
DuhAAxalN5KAXFqB8cnWfhFLF2T5wQLiHCx/ZGtF7BrXTsoWcac3UBhvDpgiCxZ6
rub22pC0Rt/YpQliH7R3Ezp8/Yv/L5FAGZqEmp3N5UBwJD7M8EXDiyn907qAK3ef
jI32Mgn5kJ/l5P0qYEogSDz4+oUg9GpT8zQmxCX+rTKPUfCR/pOhLRz6S08faE7o
9/ljqtE7toTZwi64k3x/uMbLORhQgJHkGxzMNcALOsuSi25wjskkm8wglVRiDDNY
LG1JL/+h3noEG8ixoDVfPqTB1AUSRemZClGSDldV65WFnA9HFO9AwxOPsX+uWZns
6aCNUxpVTRhqWwdmvZWIeTXmRqjxQbpgjuAEEEI7bAyA49b3a3h2LTYcp8jga5mU
C+xUsM9cHqxjxRSdDD+7gNPxYmw0bdPZPmhj3g94tIYUXUqiFQpG5FfGj/o4wen3
80JpwaQJi52Xj25g11r0NpAdiLSC4hNQYaBH+zvBrzLB8/LJKMkmFqjT2Ljlt6gP
Ph4+XfOPU13Rqwtap0M2URYHCIx4RN+aY1ROClDa+LRTj9Fc4GhAJ5J/jVM5RPDT
K/e4fTzPQ7U7mA8H95i5vOUNPqhMDBIH1jMhDr0jgco6IEynIap5q7KCBUz/C69X
cun8qt1Dgzh3R3AXLluIdZVhGUYKzXYn3LjKy2LftDLW0ujtxcdcXTgrHxMw8n2Z
4IhZmYjgXYlWRfJthLIZ5nBXOAW5i8p8LZNAZzoLLCpCIDCvTbe92wGlfRNUIvzB
2CbeJ5KjlIZApQG0CNdWgPD1fmWzhGVYnlYA0ffXsBU6TDasnsC5DFUmatXDN/PW
ODGF5TDu3LLdAlN0U6q2IBq+p0z0lgTKX9RxNb9PzFZjtiea9MBzOk4XPaILifxK
AjL2SDDqmJye29nkqR5i8O2xfX5tHHEt6+Z1i1egp52q4tx8rldPyccJ+22hX4NP
exv5Tv62sQaPXEKIH6xN14OpQ/6GlWgTf5PBqAW3Clg53oD7835khZNZGXhgUkSN
6yBB3aT9D2xKLMPlCXnYK2lv91dY2QA9TGJvMo2C+PEk2DYgga4JCOCxlGR3YLL5
av9+4qKFHe/08FFdyksG+sW652JcbwuazL/i1+5Snvu9/xTcnol0MdLnYsSuCUCf
78PxTaXQeIo20iPmzw47BgwaC7EXpiveo0D76tiQ8jHTzEmtTPH+cYfouIrq7CZ0
iqTxSl4xLrl3lho6LNRurfKsFphtGfHed5RNbfeLYZ90QrTB/saLiVUS/44E7BoI
cS8TPqwx1jM0CyBf1bqeDTWK1CYNb/4SwN87pAkXz4SmYS9GvCVtgSOZw6eFt1aR
OAwm9CtYT2wOlrauHSKvy5fiBGR5YbhSJkBjkUZ/u/hZFKFUIwQSZMeAIl4ey1Ky
ECGaMpuCCkG9sp1dVdCV8CEappzKjYYmaipKyFaXUhwFZKFoYQqmxdlM+jjd//JY
GL0pbarYH4J547wp+PGwuaKL+LnzYgKFuvYedE+HzULrKQAKKVlQ/65ohvBcMLkW
h49tlfCmiQbdi4HrLJ2Zt8kKdbdO7uYy+K7gb+RTMFUjHCvKhscbRR/XoHtmrTLY
rnEE0NzDICKEdW4VopVFVqbhmhLbwx7/EPKguvlUQt8A2XKshad0qvBC6czuJ5YD
/wWvLTQbKZr5B8t2ijR5AJeNfC43OUOqQQZEJmOXsnhFu5GlVg+XENURik06pLJ3
z7oL6naGI1RbvDvNNiT3FTHn+xTjkEjti4qU8GHC955g21SKfWgBKhhIGo3sy96q
K7uaSjRYQadr4QQTyPPA4xR7V6e9SJc5DE0zX0N/Ffk22/INhQnNWUKeHQaHvIUW
n1HTt7zn7u0kjTVTbI8Dysn1akaCFLas1ZcYh/RHKUhTujMYUf/lP3ADPREYFMf6
Sr4Tizm2J8H2hbNFYqTTS7YWFm6QemkVBCk9f5JvbXWx+7DQvX2Zv7Merj5NvBbM
1kYltr149ZlTiKYMaj+ireRLNwZV5RYzSxpJ0E09wogDtXmU2vPHNQeqbi1ZXAqS
WVY+2XyB1ugz3Y2pwwKxR/ME5KRLulbhneErjrMSO0wt0JH2fUQQnXJGMxPYEO+W
6FzUUeR/4kca6ki0WklzAVegYYXiBjRCuvLh7lRTb43X+pxeIDYuRK2tk7ovNZ0H
f58w6QOQNW2klHaIl5lmauuu1EdvGC+8/n0ZNi/22fdDudSb90cU00QD60Qz9I9M
0Iot5SuiKQP6ADUYQWMgv3e0wnJe8YG7WPL+RssQ8zfJMl4YzctNqRqc8Y9afjoh
9JdpBwxjfihqtCy9YwmZ634v4Ohu+B12B6wJdFBJkvf+dtmh44b5PtUekUnIpq6a
uwUTa0Ax+jnSGBMJZD2diOSbP4DWIGcmz1mvK+7cgWOg0EalHUCHgFQMfoO2p3t8
yH/Jh7f3LZiMguKK9yFtWFjqQw94zL/+/zledR8vHLATj2fs0tWiKQ/DtHEEmH2h
pPrX1lw1KvjNgvGl1U+l9wn1+do+nvmnU4kqaq8olYovQF5msYUOWxNX1eLaBBEx
ho5G/3kAl4iEOeVlpYp9CSsSDosJDIuaqbPVJitgpuwNt38SEcXNr8qySC3mrCTX
6jwOFXDgZkgBHk5iHvzhC+Oem4A3JBmzTSINKZiL+iosojn91BubRsU4WlsqkvBi
RR/R2S1Jv0BRY3JfNKSz0JCY7LLRgZXNK9iRhnj+42wRQKE90IqVWP3Ml6awffoy
XLT/G9P3cWK6pXKzchPSQP9hHGAnGuYKhSXL+ru3XZrX2Z9xuWDKLxhHxVAMxQHP
O9FtUPBzWadSmj4Xdq4x/+Z2eq25DozVHngtzKwjPcTuRdhSlybZA7lPyWT5p9tZ
NZDqoM4ui8BeWSWxckf2VD282iztXih1VsQcXGyDI+Bg4/3BgframAFoCXQhyGnE
sAlaJ3cl6onEQY2WO3kGcFpP6VCJ0nDghlx8ycqEd3nuDI7yvGuobuFAwFx0uY/7
bqQ5P/bha1eRHWbKZPefLQyfc/eMA83CdCFHOAKNW1sY0pVBVUtK++889zDDDyZd
zep/Zk2FQyOfJTUk2qzkFgwPbLX8zFdQKVoOs2tjFlvO2zqud0Pf3j5FSrhPybEf
eSTrtdex93CBm0lWG7emydBBvG05NTiHE94EZA+cRCsYnWq5yF1w5peeGGFSSymK
GRSdoztKTJsYW8ZrNndhrvGBxMedwnWhA/Bg+I7MvgwG0JQOBWRGLtle1iBzSheM
9c+niUHwvjOAuQp/NHYXoxsvKh7SEBSdptP0CanH8v1KuJisEyGg21yhhxiN5EJz
9NHiY09cmFdUfD70RIKmGGed5FbZUUmu/XQggd+F+vgcaRSkujz+hTOSBF9w8MP9
pekZKiyu9aCgajQUCNmCnd1/5ML9T0SbDncDuQB67pFQE8CdjJ2kSLjFaB1tH3xO
LmMcwLy7VgOGtVpcpbR8MzurHQAnbAfEjcc5kzaPadNpgFEGzSgFldKeMNM8kI7Z
0GeOOTJTjnetyv6PPSae2grkO5x6kRh0gjDUstWGqbGWzyz8dncW20nY7krDbavb
uB78pTRXwWTLnU0WNZQ2BFtYKd77hz7AUgFIylit9UCYNrMcyOXwTrPfl8D1VVsj
pdxMenzUgkcIFuKpciyGVUlBmHMU0Fh7LsYRoeg/nwtuu7Z/98Pz4/JCA4R85RVy
zScehsc594GJHA347GqdOBq8h9uU/1vYgoone7+gm54VJyLPpqBUooeqA7zRUPBz
xmt/Qca5RQAODWjwheCTfzSdP+9cDKbGEoTiVpMNHcTDPIOmQmEvb83TbDXm9Sui
tYqehALyAOvBFrgC3Xuz4dkHbuNc8nYG3SfO8RDEUSptKntg7REtuUFCvnTAlVGI
O3FwegAN3vTdygPp3/yebnEbA0wb6nMUEBkr61voc0TZ2CUrwvpOnxE2CytYIoJl
1dL7wHufawcoxpx7OSWKSBJbvJePkAvOPqLuYnWPimm5LDCgy4NaKPUjn6NaKaKs
EiWQWO813oEZwwJJjsTVTX8yikIYCf1wVArXnMw1X34qys1Y3Nr+vKj9NfPNz1AF
OUoajYLFrqwZK+8AX3dpbzZ1wfpL/cFPcktRWW0Q2oCmPlXacIPmF65cleXVBMns
7u8JeXd0r6Wh7fNgvZECpBeJXf5i2MqbDd1OJ5jKD2EbqKwwftsr7FQ6plizoqI6
/dRojaGAiCThililglypnr5eAdg3hAlR5XVpGUQXb7XjrZSZYCA4droanDS0p6R8
twrT49njj4UHrPyT1cjntgcGSLmkzUvMxUaUq4XgTCu3THaTU/wb5O5n3XucEI89
iybk3jxFxBthM70njuRMBCrfSFy3ZaH5MebJcQbLCBXraGw3YF0CwgYcudPfbXzr
KdHX2O+BkTuJYjIgPJCTsUwazh+tjXfw4Ku8H3R0dSYogfOsDmPsz7Pi55BSSL8R
Iol2sW+8ZhmtAuQ3ClXN//+cV34qVapBjfesiofchxYYAW/n9XBQd5vhwkCzxwxA
xTv3s73U4L/YRX8vGx1wdmpvd8iQ9CmB29MtsV21TE8diTiF0Aw0ntQnvfA0KIjA
Z7/Q4xB36p6NtEFFDGX6kEEt+IETTaGHXg2hKYUD/tEB5RZQgVPs8aMulCkeW5gY
eRpvryRC9aVTo9VJmmQ9jVWdx3m9Sp4uZjFN3j/dLfWKDzA/76aQOk4DW6sfUEmw
e7uGAwynU2kbWUlZklZaIZkXVn7L7jE9XKfuaL6RhNnlvm7/mai1Dx6edrl9vMBV
RSbpT1iKc4MIjy2tKYvJIvl/OwSuZFc6Z454hbN3QGl8z3QuyQQaS6wyZj4jQhXr
eNcvTj/MP20RlEZE0eDzYIZU0WBdBeOHrCxv6EACXQmpKBK7j8Im/+MixqVJXxRI
3Ghufr7WcVplJj1wppgx9quqJy4FUByUFskNGiNpqrt5KQWmmK4KV12GbhxD9JYh
3/cimMDXIqOtPnY2ynPXboTvBm5QNGQfurYc0E3k/XmZJmiiD/HziyLFWdxkYIce
rBfRkVdcIiOR4Iz30N4ObVhIS+xZt2pqfHBC4zecCFSLtkwe4dt9CPfy7B/8xhpn
Se8GcZ7TW+bSV2okOiTz1FC3N20B2rmIptz37xFmQzTL7rnXwaOJsujS6lt8kbxP
QR43KvScfU+EYE7LtxGzqM6utwDNdjzqcByCdDNh0Jlp3nYNagKYTN9zqQV/OdHG
D2o7k3MY3UICRGzbF+5TvQjyaOTW0NywIZnGOoQY+pG7DHpTorNUdfWOhWKA7pqy
0F+fIcnt9er/XR/MEH4DBIH2FR+AFXRa2seWfrO7kbyz+Ej4oscQd94qxlgOTuu6
2p/iObz63umcJ7KQ38QaLcvjgR+BRBo8TlvH8PuaOOJmsiGW+XgDa5jcE+djbMLI
i6tCkLg/uDJ8oG5vp4cCTB8Qg9ttPE5RGoBMW73eU2pFzl5wi1YJwys/EqkdqtqC
L+TXlMQJhVtibkfOy1IXNspP8IoU3ZJroB2esRRyrWuTrRq6ccr/eEGn860JJgKT
veCzjOvHcSowRHp6jIwa9Nzrs9qE1q25uXaBikDuRnVin+Yoiu2JpmPcLUt7lCNK
EZH8mfwgklAjOuHXdzj/jybrTBBq/SQk95ImANyNZ9AitLgXrfb0N6v9WRGZMA3a
OVT2irWgTaSy0e7UqlvB5cURwph+1Ehv9g2IXI92CSf7+zzZPoiPBwxN+XEnL+4X
SLGUvJz2gz3GRIQ/F/xPKfnQWISrwn2QPILr67bLyE14LrcKNzc1UwVio4AuLy4J
BK/V0CZ6/2ocW3zrXp+fWIS2rW5XySGfH8E86eoG3W8UZHwkf6L5keOQ953ZVSWv
Zh3bn/49J06rULdzo2s5Vy/yqUY/NpajUXE/wiXgrFiL1d0CRUGAKaI6c8r1SsVa
JU4nxNzL77x1mlTkIYPD5QT24OYCOXYIbr7g6QQkD+2LjxoCzSSnNdOUD7iP0f71
Lq00RpU5hLD1EvVi2Ofi1oHYzCrrXT6ZggtyW67TuSEaqsBMh3bPWRW8Q/+Vpfk+
6IjMP6ry92V3vuiHVK6R3NEzhRfl4RoPu1fkua/tOWozFKlw28IU+TXf9iQK7Sz8
gZ7AytjaOSDmYvMR723kat/mEwy5jjhgBOcVFnHuVjGJAmaX1I4Iehlw3iBrJj6V
pBDVYZ+5sy5TTWcYOy8EJUfTIZ4PWXGJG7HQfW9TcZEFCyqpn28Qh93xMuQ0intc
99fORvXyGAI6IHm7hbCM4jA+Q1WOniApHz7F1YZ2cMfBOXZt36X6st216gmv+AVU
cxb3b1HBus9gpqBMdSdtFt88hO6fwjtvUiHohgFTLNovg8/tPRwD6uYNOf3XyKft
Z+h2EQa3vbhonTFkbgsp5CAyapUybKkdpqFWUeGI2LRQw+lKfdI/R2JtklpYS0VC
XZSWMFranmrqjm7g9SSIaDfJgXYP23s6sLbLTiisKGNoAp712aAdQwKNTJKb2LIS
GiqmLA6e9EHoyrK69OtRUSPB22w0dhzXAjBt1CjMfjvLmxWzSYTr+4hBgAp7ld3b
sHuJOvvbICs/qzp7IcE8giAL4eFNDh6AvHOF/5LtuDJfJA0tx8h2sxjXsIa2a4hN
ogSTnyiUZV3OGMTdaOttfmCSuePxdApyW3tVQNbnsEPxD631bfiU7ypWScK2+PFI
zuR5EdK7UCEQHl8arFayMuVU5Y6vHaQoKoQlmMNR5Gy2XihNOUbhaUKoiMGAcEgS
2xsgBzRCnzUJAOMAKpCNrBJZi2a0ag3BkmqTfo5JY4igQYiMDf6rgaCt6TelgwDM
r5hGyruA/fDwUMwdZgvzsevktMOu09tRXk6wl3J7t+L5kcSFTjc5a8Dc+z5RybhK
4OR10LMZEttztHdr0srfbyaEFlUC8a033jQqhNa+w5MfxTuOq0N1yj4Mg4/BN9r/
Ki1yG1lUmUr+tzjBQ7YPot0R6kyrXDk+MRGNdTwNDFD5w1uvKzBOEl7oIfjkB+kq
XsMkLE2WsvND3w+VCKkOQzoWdFAZmGHusKAcbc5WLmWLkBwk6xF8JjZScqCqgeCf
NyQiuiNoYK6rpfy1//nMgnLU93M6doPf8KJXsne9mh3IND8O7G+6fKn98ym1qD/e
VlqngCxHm8ecgVxE4rLq/byRURv6SqsyfI7pR9azZzo8jNyhX+ejaVWbDV/Bu6S6
pYEUZ4gf10z2ghICq05eEcu9oZQGcAAvXlR+nBYt8jxdY77RE7IKTAyQcqKceG5o
6/0iFJF7PNA6cWjJhXAEtsZ0htD02iCw48HgZhDaSOEQiehSmjkmmkWCVDRaqEHH
Rr+FE9PSbcHnBGpCwJx53VJJPttNyi0xYD4aoDoDOcN1DPXHe3ywyP2HwtHOX7g+
B9qnt1z/WE/tOGigCrCksD5NC7oJ80ZZCha2PVLLbz+wmVDebghiCigNyiIYkPfK
DXgLjYeEhqd7ahctnSeRLtzwWpnGuC/nRwwyIVgrnkodmkbnvXz6TNyOxbLkW+yA
TjeMqfYEFs9CTDuyc0MS7M59JPbpixa0L8oGL31FlTzfCop+yFpABBLNHR110jw2
687UvtavE10IpPSisU1q88dw/5FQXwJWmD2RlBkIQlpMaINUl+otBgBKj3nv58Nb
zXGq3gF20TfJDMGbiwlXynIGTlwzIsd44CEowqNwKNP5vzaKObYAPuPShlIjvkVb
vLaLYdQP3e/nZtz9Ydyha5vcsji2FL+qQttPVRWqgxR2JwYMea4cctayqJfCRpyM
k+m0keo+sp8GZ9oxDXkZBDgJj81+fcHa9O4cuNNmkPaVExn12gtgof2XGjQEBKqf
Bydj5FcIyx/zzVbilbx8erHHLUeZTldnGSvl2BmqnXz0qIcsIFQWbia3rOQZostj
makAb+heVZILr3VaJM3I1cAvWwkNKZ4sZxF3XS3buPuTiDbtwFtE+iG1IhNhFNhr
PS3ynKRooB9wDjykMgm+yiQL3PHoIK2CgRaJt232gAZY+GYkrEVeCCW3iCrXaQaH
C/BtblmAd8M1ideVCSf4ADKW50MK0mmfPDdlH4M4kkIV27qnWQJE73y7tP0n+tZC
y05m/uiDKhggLWPSMMv93Qanb7EG12ok6jW0/2yG3gtDHVjjZHTERNt9jBXeV9tI
juYeVRcc/Ys1CRFrxJCERMoIWa/0/jfrytxts1lNeZhNzs9yJv/1a0i0TLmTWBpP
dekdbypvoxzSriyl68b+5DO+rv3s/mmuO/U/rZ3CYCL5zJJeANIfF4RiRK/bYSci
TsOK/BxgSAUkdvy5pUgRPPS6nRW73deKrH+mWcZCdCIgrA3Apfe+XmmN8X5TTRXd
QaHkzyLfMmsMbzZIRoABu50S089t1J6rfHISEvD+xz6bnZp7ic1YnUlEQmkIXo7/
4B72/ojegjHEGnCWMNAwdAsP3NiA841BQyCceiZLAVxH3LDuY0SBaiNai5Cx7qxB
sKBnstlW4tGtdLcvqxQyn1mpbqmrNGzvVLdMnsKUuA8VNwK6x4dgcCEZEtknV67j
0sQPOv1uUPVtea+4yjOntOWJlUJ+em39swPKNXK3updwr8kswdgszCv7QqcLmNMj
8ht78DUlx0ZA2aDHBxnH/VOQ1jh7+QnFPBjU/kPYgs1stBHVF+A1CMQ7GZbk0KIP
VPEvCdKamKcxl3azGTnNCeTVErCZmFhqroUeHoqCbnBLmwCpywKH4dm+fM9Ac6S6
/ZjIbf12gLpWO4wGHGCJiYZ4Etp4X/v5eabG5ObPhu3mz+smxhd2OVfcwEb3dswS
omcp/NvT36D4Inl1iUOr0YEHouBTzRmPJywFyuv30rY/kBYWeNJNMlhp8km/Ilxj
K4FRw4qYg91hEXWfsQmJPfp9bTXYGfKB/fAN7ot72JVkymtkLIZynOj3gpSCE8u9
YBZYHVfTfec5+ucxz39UosywsaAUUGlMqlZjIGd4DUJbV5n7ui6YC52MPJq8s60k
BdiHRAsVa2ErYsU+zAebG3IHUQvepgLOeuBookr6jo6ssxWOQfVNtDOrqASh+dfp
MiCHai7npp5sieQEaT1awYJ8xc7QH3a0gZ+yXUBPDsKUeKl8ig4Jf6kXv4+keSTU
1nVeWYpaPv1dyIGheEk0brMSNu2WeygvkpPivo213aGtDlm3oIqyQ7KImR443zs5
tB/N5T1zePHFhhekCE9BTUn3R/43r+Jl4HADFCyytoo2OvD75jdUiaggNuVdHj6E
ReGLXH2DdTnNPF2twNYSEbbtZvumml8QcbQvFlrpa38j0kvCdzQlhMhKt6qdFcQr
YEqLyJToA6qlpGDElaMCPllrLRMHTyYN9Bh7o+XFkWAPul3bFYauJ5NW2v0/3agI
ihp0OtABdMb7BOi9BdWvo5dkJLdNzTJ9RyuiS/cOOEzfOkA8ro44rvzyv8VEA2Nu
hfygPfQXMtorn17v1kgVVlD5qFQpdbzIb9GSBYajOrALSU2LjzCZjjsuizKycH3m
QG5T6yGj6DcA1sYn6+OoCbhJ//ciOWLTCsxLOXVYLpaIjlDX9SWdGCiXtMQzYmjU
t252y6ql7+cfpkgtjGLiL+ywdONR0/yLfYrMpz7WxckvHWMr09k1c2nxkiYfxCcj
8736unwvNhk5rVi1mtWV+D0l9H0PY/IlTefwlR8w8pXllqp2oBTIfFhjzy8vgGG/
wj26CEllVdp/UsE8OIxJ5wqs2NsoWyTymQzOniR88sX2FAPH0wl4P5vjS8z/6ZF8
6jotXLeg1D9uBzSHfK06ijDQ81ynPakKBabqYHtofZBVP/MVSkScBQIc/oIYokXq
IMLPAVkvJheJ9vzmwFiWNqkD7xibw4HOFh4mN1hyWc9byo4L/bwO8W6hqenI4RFI
Uv5N4YQo4DPt7jRgU9d3te3hIW8cbLjsUdiLSxkhEY/Cw6rwg18Rw9tbkA19xd93
xen+TsC38axMBBIIfV46LhK5vpXzgeWkBiTwiTWboAnBE7URuYmiz3I/tt+LrLlL
Y0VLAFNHC6EgoM3cxKv6pzihQ+7D8GFguwvZ/x7jCgiLJ6L91xOxUBiktyySDRe6
MUZDUwg7YdGNbfXlKwyKmaSG3SRrw6xjhYohA2O5HLjv12UAw+2Yg361e3cQ8Gdi
nySPvfnJhK9CqGQX1K6kM9e7kYqNDrpq1uSBGkoyotXhJLc6XD3KRXCxDlqwbxUA
aCGpobVBkAsmV3hvsy35Ypj3+DGPVRMhouNNC/9roDMsbQW5KbZKH6mh4sqrsgP2
86saG9Ot7eNsyBV7MGonGuuAdlDhiQWUR5exAE7fU4wQgf179G2MqgV3HRiW8tif
wUSAMBtYVyBNARsny+5huPfhdiICLj+EBpeN7B/DT225WTfXQC/GjF2EDMgotlXw
YNuoWdut8499ivb3260IYc239nZEfoqytGMD+oJrxLAxwLhpP0qkSvJv6jLWl8Co
miv6AuQnP5uUTFftnRdtCVE3zsBaDDBMSi+neiWgRr4BNCmU7/VMlssfZL6wTAST
pTB0C2QCgnjfPvv4+iADxSOfbjfGru9EBP10U/XJc6WR/urmWNOxzieGbB0CUWp/
ry9SzXUNDfPwrAiadAB4irXmrLi9glludaYspy6v7F6ObNRVHNiMk4pQCymbJvU1
2zemVx67NuX9IDRCDn9ZUsvWaTGT5uSlpN2m6RbsdBeD3lv1fWXd03D5klPcRCFu
04Hr+5hI29zApsOqUBxju0f9AW5a3XE3ZKvutBs9sbXQUVFIdV/06bbZztL5ubh5
ERTlC9iErs7kBiVqmNcfj/lYc1HdtJC68vk57vJVkpZr5qWRO3CLKIacBFXm+f5g
wGYlysTTpJ6W9o7A1SdauDJh9b4TQQBj6Z2In5i5BLAFecVnDiqtzVP4xM5XMFuZ
HW66W6EJiTDPHRYDVxsUuR6ni1kyjhkLZx/G35WMRYtrUmrdZLwiMYnkZCswBtaQ
HfW6sbZnap98vxaLPnCsaPNf0GKooZZ62ZnChEi7xWYajVyEkhwVSA6KJFLbsrC2
P9lxWhdTvSRu251nbc7HO/le2DiwT8Ttm6kFoTozq6ltwS/Bz7lOjThG2AKcKWaf
cTnHt0XKOv/Ym4ZQL3dope7HXSJyb4FCoSbRmpXresD/3qJtaUi1//l3jzCyhbzC
NUjoJG+186RoccyovltzfdUeiw4dXwMFI/az28iCYDgxxSKzDrySzuh44sbhlOuU
EdsQyHOqHLFjDI1Fky6ZvGOwL5BKuINvCbo33dFhqNYqXIhEX1KmLbVdmHtLr3KF
G8mt35yo+SFC5i9eFHtZSmdSTd+RiSqG4fMx5MKvZoVaot3sIiCzbZtIh7LWVEXH
A/jRVsmUccoAcVSpLqa+vqnW5xC4OFY2inLGNropB7QjcevPgC58XZgwcp6hRxzc
GDwTrAIr87O+7DUC/8MyD0WtkyvhAUDWZK5y29dV1fIarp7dzDISAwOZ/BFitBkL
E5n6WUQhurz6rYoM4R6rg9xTaLW5NTFErF86KsgTEXjm6UUifclMAbA0XmPVR68z
+qJGZs9iTUcbYI2MSQ+hPh3meSU/V2LRc4NS2dVMr0apSFMl8Nkj9tXFqPz5j5Gx
BIzAkmnakOtdm4Vs/BuqEVVGAQC2cooMeLEJYYSFLLRLzlbzHmhQGaO+q+JwWpjJ
0YHcDEAZtjXFb6rIdiZx7mPmYtkkifRDlHWWfP8ii91hQ+fcoHNPkbG1cC8TKX7n
QKMvXO9b2DA6QhDzIol1eGvMz8kx3wfkALAJNTwYCQpWmgwpuAE4aNrhgFpX2GwM
rBCzXsJ8RtmHvE9ZTXHFQcGh3eFPqIhAUI37WGfQRz37I/dr1fRblTs4AS8xb4qA
2FcnzC211CRf/6t/H8/8D94jOcEqkf2E+rQ2/QUrTEkpUKI0xkmGcJNWkz+AAfVm
rEFRgQ037KD6FZYLFysiWqqW3R2xmtfXuD/q300BREbur1pZpYxIS+hsYYduM/cS
jNAKMAHZ3I5vr4xFI/mRCLJw/JU19hBf6iW7uge5iwhHaw9GPn/2M9ZTB5ul5w4r
URSn4/qk/mI0MLn+0JFyJVC70cGl2xXNBnhQChRSctvzi7rmbnGUcggVukawew2K
jXuqnyiAB4yHCYVcqwD+hII3nUY79izIZPN0xt6ghUfOaA7h3UaEMgrVpNYyjEhG
iPxOt4K3iixJHPEY/bBZHOBsLcHCr2Qq3G0PktFoQGVxIrvhu8vhQ5CDI66Rvg3s
JtjJpZCqGqUc68UtI5Xe4DErn0263oL+7HRLj4uZ2ZY0HPzsHhLwsYCNEdMnXpsn
8LYclRgHY5IQN5JedNXj0uVUn/PCKDV2FEbhNE+X72RCzfab4o+2sQ7GlpzXJvI6
KY5vUjsfxI8rkOKsGmt/L9XqW5z/h3TkdYrgsPNcGUT9Zcb25e9fd90ff96jmsJc
5vdbe3u3TR1BlWyfumdTfFIqcEvzxJqEcOXeYkgtv6TzZZ2LTKQ8qJgdBdoJqpwA
Om3IZq5AUj8Y3Kge8ewNi0NLl9rIkelnYqo92476hndc7sjIv0nQ/NAKi2wZ1fAo
XU9xXeouztBMfS8pMKXMz1qoUQhB7Kxa5u7tZI5x2WgrAzc0PQ9W3qvCGsDBIbTW
fRXv/x6ABHX4AI1btCzDT2NuekWj4QLG6he5TDKD5luDy+WX4r0l3hWvEoQPpkNJ
9cb1bVrsm6+2tkyd7JUJNM3UGPY6GkX2QC/Y9DFSG23O9KC6+VTDbIhXFSm91qh/
yasjkYXa+U6Y9ytyPnkNmad0SjN2dSLSOlYFAA4mkcZsSDPMwMtrCvcSudwLWgez
Bb/cRkgFOVxvRwq/XRA8r3EGL/dCYClCJdYWtGvC1d78bJU76lcSbGncFQhk27jq
nVnevJ5sOpHZF2zSx6pAg/uYFc01vIPSjT+xTfTdLBcyyzAIz9xL2SMaD5sLITHf
tQjaMpOW1EiUZ0tl6M3d0wHRXLmYkPF14YpaP8bPZkz2cN5ZaN8jQYXdW9xVAVfK
s6IvMy42hlF91Km8b6ps07hwi6NT5bgW/+qnVz8T/vYkmzpGurjCmC41KmJDEE6E
g1Jp5UwBaJkiE8Qg4btihhMm3yOsE2g4pIBKmRpTudtpYy91wMO1h2p2GtojA/2F
PeTod8GLDptupTRv/W4VxSauYHFmYUW/KnvWa5Fm76PpWePVIszbvhDG8qIujHi5
mApuyT0b0FhhSXWh/Hi225WQo8ERkuCf+L3rKLiuL+VSicMKqVu5dYOFZIsqYTQ0
Xvk0H0bjvlMIN6cpisKMin8zpdKN0b/GIALJSml4gZvcWn526qlZjQDYEx9bPeFR
4TTdVNov3tpF2XPwm8mEsnp0fnMwQPRYAUKmHfKFRRGr2C7SjMtIvGQpDJ8d/0sB
MITZ0ONfch90Jf6K+0Xa9oBn6pLWt9TzT0E4D8qQFNOxZ/T0pm4Q2u1JGAimXKV5
tVm+9fHKUu9VWAvoA9S4KrB7bUepSjWOu12RwyGba0Edfl12J5YBv7KOgnUHx8bG
qVWebEZ2aGEVQo6vZ9Pd4EaiMzTgKPtLColLeRaVbrZztjIOwFnU/aPLNGosuwZk
Nc8oeImrDwLrQ3Nb0/CLOedr5jmrAtQyoiELfpj7Ie7R9mn5hcYsO2W8gi793l9W
UGKQ1jjaLsFagjXa6BaOi0DXALOXzTMG4oORIKefBX+PUlAfUUAYDe/vaVkDc5Ru
pTm0c+K66p/Jxm9CsJ0SHqoyeU6HN6CsqnJW2l2J/lUqBfy1h8YldrX8APo2NoEm
Rz2kE/TOhxrJTmD+wRIryJHUpBpFV1xhE2uCpjgZI2V9LijESkxAJUJ2QzL++56z
pCvvmzQHIQPqRX+4nN6icFOKdOfTkIv8D+Pn+H+NjRCmNp3trruJqGRP7BTqRIF5
ARxEU5uarVNR4d2wVFBJ3Dyad+EV20XemsbPhaOS2gR3cftXCEKJahG8uLm30GU1
kUOB+UOm+Rzduz+GiHBJUPnmivKvuBSuT6cgLsC0CFwlzk58cUubWXBx78xAbvd4
yjIz8wcumVzsFCXBn3epbsb3zRS/SydGMiMuCDKLYT3wI1hRgJeBeskQTFjad0Cg
gRn8imQZ0AzqvPNygJvOqLoy8Qx3RAlE738BH5Z6FREss+2uxM+pyPtexmfbJo6H
ljFDebXFmUQva53RAIoccrdFtYfUUaBG3IZ+QDhbhAdC51UgHGkzVEMxz0pYpMoW
4BnKoDdSvlkl1RoaDg8NBqOLgxQIqbabMOQeTEyGoSWGCH4A0pWh8wzNTOI4A3LF
I02QkjSmUd4zJ3CUZy2zblMenw5O5KKwQCfm+SfJ5Wd53iFZrk2s3W63kNfcYuHX
cT8niagvWBzl82yQEF2FWyUZf1EACipkklMJcehPIYzE2j2UTKfRvAj+xRusbpOG
dKhg7FzIvpemhQRbQqxZLi7SRVoObT6DCeQPYx+ETu+InFK5PCftKyTWtyTcuPut
qDODxfGlvdfFjrADewq4yngPUDXEKIFWNDFYfu3TolQod/hiNtCi2s0ioeH19Qyk
olOVut/xdGhXp1qWkfd2mj8aSMBsSXW8YvhbzLCtxnzYUuufjccokVj8Hxi9HSUU
axKwDGdHb9tuX6sFsBlJMGtRcQuqOv/G8WE5MEWajIHR3dQNG6qcRgVYHP8IgyG8
rcW0/hzLjl8qH/Ue2G4Fb+WKlCzusyvztUSJfUdZEYuAF0zRpsDKstzq0bnyw6pc
EmoKdR0z+bpWz76Uaks77fd8DXH2ThnsaUXPIr6IgDNyAoxgJUw+yoByG0jmefSF
gbTkVOC6B4ZnECH96BrLzo/gLTK6kTYr8hFtJb3rlwsDAGpcfRqhpoUMPJljMPFV
fn2jTfLYNwIFDJTQ5wKSsSdLocBUsqkTsqbOYHErSiiJ17hv6BXxU9m4xsEl6xvj
LzeECFNY3DQQSHt7m7Mq+B/IJrqp+tRHGGebFn4irrrNgyEuDVrkH7wz874m87Zn
o4m60qJMk1hkwLmALJ28dN59rFUGLAOAti8zvjSnpiZgnWuT0G95AtPCrIY+W02k
+m2UTOwNUKdB4xCyKSAfrKi9ONQ+93xStv4HgKq22Lvs6eTlPCT1h7cvC3OFbD/2
yWIAaInKtwiIXosTPECBHW3EhjBooqwUAdddBQx5/sEcgIV4Srlo0jO0kBAz5uhf
nVyLuLIX84f++TEx61esw/h2qqgEY7rIKlXs0MT6O4SvQOVERHV/GEaJQH/1YbV1
AePA/bnHD0tsC07Ae0yx+/BigpTKuKhOfX7qNeaCpua1p1zJm4UyZ7ruSS/tIy86
2EBKBXEN9dBe/XG3fiD5vh/HQ/rhmz9nr+nEj6DFmjKSq8PF9Se/5t02mwF6rvvH
uzT491N0yVDwOJFK5CDHBARWtpOKTLziQp6kwebK0RGDHsKwnVASrKsbCI1zkTi1
nlOdBBYoxik6GJb59Io9JrHxeFLp+gq9o4XXOc4TUQSOWjSMaoY3PIlDC5Hr4X8+
dXIZwzp50NNmZHhDU0iXoIvM3A5uFHrR3g08DSUHCbNpDxwfst/E4p1U1QEzun+w
ijrc+hDqi/XPTpoJMm18q+Xg5OSPPaByXfGk2mmsn+txEQpkw+CV+O+cPB4EQ1Bn
Qb+3apbF3wx5a81v9NBYrUnSKmaODHyiD1/hhATz2JLvXqRnQjtoM2GrRb9yVTBs
kzCrC4jIqP8eJUZAvrPRBeUChcoYaMiHWTXclLRhNPsNeqM9rltd0OcU4auCZmCR
QF4eDyE9j734fDBDtsUM18OTfbv2vdSZS/DpU7Udlxud1tt21OFWZulViYnsVAfG
aCYMQk0XvHkdSws/mSoBDuxSWM1+dMgAc22uTI/K3bVSjHBvsOR82ErNpO5n5d+0
kUpuKukTcbLR3F3ZXCLU/Ve2Tfbt2yqyQdaC9kFOocIJ8NJgXz9l56Qj/KBs/5H8
98FvxBEeiB7bmmvkgIoyF2jad+MQmnKkGEncJRCI0J0aQIL/DvRR8uaeFKu8NJ0R
bQCTDN1JDKtN7ll2Fq95n3/e2CG++lqgb1ijBolKH/jAEAy9mWCWJPrIkO+mWeVZ
3Qp/C1boPo9T0/V0ERAX3gCIac+kPW95uAi43KKhs4DSf+AL+E+YWjDIQMXDKtxi
OMsSPohkhp3SMUeCFvFbivFjqwLmv5Ao204LKfrpGh7JzMfHNUi3aDNXr3ovQX/3
+jJVV5OVGbeqiwm7NmmXSKW1Ms5uMeE53wxYYOL1cYewrHPyjv172QfnYDgaEUJH
n8z5Sq+bmDG4WrzIXWt6gTI0i6KDVXB7zvGW7J3btO+/1YraDmL1xh78uradMdCO
C+OXvbQny4L89FTsiLJFb62EtjSJtQH7sxz4/rX4ONa2HKG3cM23/6D4GFVDOqHj
GbWILZOtoRrgFhGkYDxR5oaJzH1y3jqA40Qtem/oGkrJXZw+8EUdiGCHOdU4drwl
pf6suLShfkP6ZIpcQuyEGu1LHZjyVhDhgzfy5UvdRvOxKw6F+HgF7PlEeIeE5Vjb
KMC95mT2bZ/W4fZ/k/5BbEeoHeGggOg2Fy1YOkMNiJcUL6QxjgPs3JNaN1OhMB2s
79hxnUHNVc1ZZ+ikv7jYTG9yEKEOEAs+SAt7E69l3DQvmiAHgd+wI2RH5aujLHgY
2WSfozpYvnZpnYiRLcQ71p0wksljBgnKfO/RwNccuCUVEbTmHO2cB8oZGM3KBDAk
eqRlxRSv20NOzftKSzD93YRBfeh7QXTCfXPBv0TRYwnBWOtt5J5B8Xokjyi1lAId
gURhzDLMvTeOevbzbiabguvzHJIhsIyrnhpDnpANuK7lJIgfnjek/+tOxX4MomOH
a3T73stlNo7swDZ1FXDwpIkyPr9gmBYqf6xpcW8ruU+KQwLdrG3YuQYwId4Kmy04
36O5EeW2lT7FpOxEPQ9aaAPfPbudZhrrW3fsIOrbF+tthgntu2sepCGt0yy/PxG+
ARLvAxcItNTOba6cS2Tor/T4Oto6nCQ7abJcqVHz3bJb3a4Yq65BV7tFdKD6IJGf
rJqhzk2cdV4q0/7dpK42mRoabnOe92BoWHrm311/KmbMVGqSUlFliEHcE49Q+T9N
YZFC1M59fRptihD/wnm3/mU9rZYwy1cc1oCdW52hBTXbHYXJw24joEyypKTWtOMd
9Bk+/mO4E4n79aTPlCdrJjK6NvijmxWvrsH37LjVP5l6VE1LGb7OyWIT5FqFMPIX
AVB2Tin0AKwVeSOn2jUgBlkAXbeKhlemapoWCXAdEDJyZksLFNre2tKuMk/uJl3O
z6bgbuUaqEG43CqGVPzoHCNwKo/Qa3cjAHEcVYBSLhDV++EL3S6HPWYya6va/wbV
OfnK33CAIpLD2sfkv0qCRa7/1XF/JFTEOdFq0tZZFncO8d1STJv4FhrZ79Cw1utb
xvLd0IDfEzTdvVNdagw5D38PXRTo6c3Gu9iwUwg+Iy/zJnjkpV1GwgAammpF3Ypu
KTtLxJVRreOKK6OH623QPpvuAubQ9DaH5UFC1uRSKCNwLqwMqrjcwzYti1EXVla7
IcXKcCsYIYc1gb+rcY5oHsnZrBSpkXKoK6ZOXuuWwg35PjjYj4tn3THsMJvkCRgt
6IELMCeDX4OXZNn5LNTf/hoURzndenxIV52Z/iBypclqVVlKtLxwr2XORS09o5eH
gdArMkMll3oavPkeuMdpgj4x3hfGVlKZXRxglywF0tP9JZk7vcKzW3/zFEf+dTrC
cR46NoVZC1EM9kkgG1hh20unSz1QvdC38+pHKfMaLrJEYgG1BJIV4ONyxJ7XrWeB
FhB0Jz2sB1Lt4am8HOZPtOku31tMVoIF28jiVgw3F0/YRAJx6iebsN3vMIWZy9yA
uaJ5rDOuy6RADWactNrZyVI01MiSfTGvrLFvzCMtNE50ILFVzA77vT+kv0NEHt8c
s47dPAbu7vF+huYIrmziISsRHlbLwuUyFVfUB9jRA3cKeKhSJP+bcVgP1YWbpspJ
rVmhimS3RC7t2TM5/E4Jw3Rd9A2ddfHxs+ZBDjLRYCOKmeuiY+ZHwztQZmyuzWEO
qLIeVD98I0e9owKbI6IMEVrSF82TzfyOsZP7PCf4yHdnPL1749CfouZT4tXj/I/y
FctRzaiFFrZ3ESiJqfNqp8iGvsYGC9xfkknOGIWaRHTsR4YavIIMkmjvDC1eO6Nj
SXOqWWT5Djz7H+MlO/OMo7qm6UjJUFJgbcbsuX3L9qjFKIbBHkbAjP45fGzFwvPN
fA7Yuj3WGvjm6g3pPtmXBqnIsKOsi7VVdJRCKz6Vr3qyXcoJQuyC/Vir8USHxIsc
K7vRj8T4LI5n0PTsfZoBoR5GcOTQMz/ghtfFFW61C0tBdTTVgFr9bQL2DXKMSCkX
RaFuwBYqC/fycKFDky/11Is0PENYaPcG/N4VtTcuOfLeDb7EZR2ms2UaIjC13Ese
C4x9pLI/LqT+ePz3UyBPA1NklScaNQC1xbvzWSklCcMU3vqtllMGux7jYD10n4dB
NSxuUHLVA2Qx33ucTcEz4aQJSpxz4L5x2H47c7yRa1mF69qaHncdzocinwIs6xnf
I+rzjHC+98bq2Pea+C84043KbHgvbVQ1czVVPs+7swB4lP2R/fq9PWOuwU6+Zosv
exvD291elGJcOPf3vRP0MkLvW+eCNH/prhPDGvK0T68Oih/OgbSbcO3FylY+dOgg
XqmA18tMwuj4licBZCiKH2TTaCXLfV6Ezr0zfwNitl50aEvcg92puvFaagoPAWHH
qXHFLE1rsJrO4oLGInw5IZGKOUq8I1WXgkU64w1oREr1Z1LShDpEZ8VmioVgCpQd
0QHlQHJGcSHI8BHs08iVivKB9ByHoyObVDTqEBHlYXSOn1fLfrWqJKD/L9EMOC+0
pVEPC76nM0ThzBoUHKj9xHyK0vwR/kEUl84TG7/Wn9EF9QaayaN6nJlrrXauC55U
eX4UeIZ69SC6q+BiUeBiyBYnCo/lIAYHTPDh8gbJr0xZ0p2VugQvSa5M3Ff0fUK4
/jPmzRBAhQA9QuO/vBxLnQ8khI8jfGdxhgqgPzRGID3yJWNVMhiCfY3+sgUhRZnL
OoBTgaV8qHWGYO9dI3UrvCqKEu3+sUebEoNMeEBzq3ydgMeaeYk2t0eZ2YxvTYQj
TpnS+KgKQs2zRdO/sxUECr2UJdiHYdJ1GCZlsuN99utpRnPlBc/fRiSbincAWLn7
xhlMdKjiWF8aQ/5lwpOj6bOfCs8GuhdYG3rlcjkVO3lZnWCgTmootSEwi55nVuuy
Di6drev68p0tC55+TtBUC/wC3C7m7dAZQlGhm98tVAkqTRxmo/V92RLkzJhEqiu9
+XhRkjZzPApndjWLHdnx1z7laD6WSlXdvDWKVQd2KllnEZpVxM4yrzfhTg3wlOTJ
xLxo1O8q3n4ygRPYKxiDxUol0ExcgJEr1T+ZitdWF+Sue+7N1PxcAHZRqeFJA0NU
avcSurZiJ9iWR+oqSxMjgG5VcqLJSSTecVnES3HvkVswyXoEFcUbvAp+q8BH0HHR
iOXFcA2WYhbmLrL7zqgMDkuVHt9/jmeZwqwAX1p8h4uDQ8gVc7HPAR0INkDq5R/C
e0cvafR/Ki2DWmawPiZOUyOEq1zjaxzbeAvAsuc3IBj6dq8OLx3dOsM7d/JwLINX
aRC+L0v8nNsP10f8wbskSpum8DbUVKBz9SjJWaeqd371lY759zf/v3IbpNhfw46I
mTokGhcUXhaXFbOz81+W31pDlMON7IRSwqUZdO5IG2flYl37UxHFkCQHEZ2+V4xr
Al/3PnZX1h/AbglDAc60wDJZVyRQU2OtTvFYSMY5H3wNvl8nLd19oyXA1fSXnAuZ
DztvnNXrcd2T1WmSp9t4oCvpS1Gi+vKH+NT9sRxJ0wG4/G1oubCzDIyB6L7w8N0J
qQXOyTqq3eDIhaxjtsjnVf7HxnJGAsSAwg7v9okDhzCNuQwdDsP1bkqyWvDmjUcI
fUvmM9TGUuhNsgwnhK+Mk9NE4V+wYi0u7x1qVxADCiGXxaWqZPJf3HeDZ9/XPmY5
kQw3EI7hh76evMcFzIUM2hKlvGlo9rJ5A1ZTdIM2wqBluGNRCRnoA2M5gc5EgzOZ
CSVs+IATbaeYSCLj2JRIISMKe4cPx4TooCQwmOtwWkHXeRdUCqHamlPY9UTCl7Aw
pQdE7C1cRB6pl7sxUXuHk2p0ER9PcmTbfv/rEKsR0GkwWsNIC3Z1763irvJVH4Jn
18Wp3de+mk7fFUWt5FfmKpulf3qx2h1u2pYUNotlGpgePgact51k3eu8//EGYmrW
YUHXibFK1JDtISAQ1C7/NpthxCJ1NATm2gzKSDcFi6Myvgle3FtrqKTyr2slsRES
dGmLGkoaQ6rm3VlnoO5fUxGivyDPnigCZw1a+7oLeiM548NZ1rdjUwI1RjyBsLlH
M3dNyup1+RzwlhXYbp1s4qdS6zhfQyukSuTmWE+3QpRfgA5dxYMflt+ue9MQAFMv
ThAauzXKqi2CrTLywu7rmGEmnIMZOd3X3s2cUaVVjFdhhlGHpQF2cKHHOc5gQduO
oxkORyFx/z6cYJEGCKpp8o7bPTfHME622qPv7vxt5kH2s5390iRuG42HhsRp2bI2
XDu13lF64n4kPO1gkf5NmultN3MSMdLjkcY4zlz29FuOlcQwIVC/FjTRUVCjoNEZ
uLwPojK5wLI11xPZSNhVz3AMT4CuaexnSTgjmEfkgjhR75S7L1lxgTB8y8g7gtqw
6MRWd7s8gc+1+Z9+0ejlFp9cDnvhHViJGspCpJPC5nDOPlqG6frzGG8RUmIGOxJL
Kt+4dTm4pfvjpFSvngqL/VECayQ3E6+6EgD/wtajuMnxtu3xfDX2tMG8IwXj/Tpk
RloVeyc2JRCOYdCG6IwB48pYAuubv0inH1a7w9evNGBjBKWfSQh/BuUCIkC8SO7B
xRDmOWVn/0VF1xuY0ES7UPVXI/febQIhgZ1qPqNdogyn/iFoidGZqgIv7f1kBKO9
PMWxYbnKsPHoLYjeKFWnqF1MqWIklcU5PXlw9w+6t6DvT6j1MuHNK7Ol8UkLNq87
nsiGD9f8u7HyT63caj92kt9mkAp5UBnG3u1u4Is5cqxIKuatk/ohFCpwf3YJVae0
m8V+y57SSRUoaHEv5746iA2Fye+0vkIvLvEyRCA+hduemNyqURZI8PfTahUDl4OE
QZsmJqZ7bDw2G6DeueAlmXzBztiFnQSTiCXcw7ipkxbP/48ZAVVjvkjJrI6omxN9
z36t5PQvW1+lphj2SsCtpskhGcqFIekaeK3tm8PhMfI9vFmcymeJbpCXfHjaafsy
e10Tkv32xCWRUWkd1fG3LMnt/BnXSlHcW4zZN1N0Y2iOoTI+KlWbnhM+uO74/zfK
oEW5z7Qs/S2ObrE+wUf3TIENMUeENKEbPAfRLnjn7mg42/PAeXsEmHaj/1IaIzR9
UXaU7NEziIZ6h1CJ61EkdUW2z7TWKsq/KAmUrvlvMzKdZRTKdrW7v9j0KjxrdziG
76nQPjraIup2tfQO3aCp7NVZDv2kARtJJPSfrV+p82haKbKEkdtjmiexrCjieqti
0oWOW1Fx3hJ2ubYcFwLLquR3LmZlZ9IxJQzXtoUB0EygcjsRHNt5cYklMhGR5sxt
+hctxIfu838v2B9hKCikTloGfpiaKV8AH/O1E3iKhrCsJ2XvOSPgoA9NRbFNe7A+
LSJScl06ODHWh7KRt9pDeX/85EivUtK527iSA+gVbqtNnNE4aRHBOyHVZ9Nv/o7C
cMlbNXymlW1uEft15GzroFoXtlkkL4ODn+wbEEgMX0qvfBlTWnas4tAqQuidtACD
c4zz4m6voKGqbCOhpAF14DXkodiQ0UcRzbMXIvDPw98EJ6dkO0Lf50jE12Ky4Oe1
xbrlf7biYA7ANUEYZQBwv46YnK4P5yQ45K6xy91Sg6/Xsq9vPOvHc02TrlCuM3jL
wPzZpv8oHhOnUQGU6iJksSa0CKhbMT0bDaNTKKmMWrf0FqQZ/8wq50zODz3MYCo8
2IoPrWXlcey9EVpKfClSkfVvAFwACW8eg9crZdKkrtQDSkfkeErZ5OzwcL4sunQU
/fKQt2Kd/iIO4i1r9WjV1icKZYJ1NgHSLXPgVCS4hLAoSKiqObtF4S04JMf1BSzh
orComZdtvF84Cr+I/1L3wuTlkOQTFacbg1l4mXhv9aXpalJLKEYHsVXQ6LrBoDP4
feQbIIzKE4D+x4fLQT0cE7Us4H7Cg0eyCr4lwvzN1l2npq3QhcYN6hXtVUqDvUFR
SLOcpThVP9LqRSE1PrRLVkw/36OzcMB5GPCFB761XuRqaOIIKQs7ZuqN92qRMYin
lWMuEQF+zMrZuU9+PiUT3pReSFWVdp7x7yjzjX7bAoDBOelKGX0o0yXdX6vGFoCr
XDWhom5I35rHebqtC/UFpq6ySjEgV8Dqo+EfzDp+JX/Swrc8XtsqeQGV+WolSttx
BOYJ2Y/V0XduUhfiJx75KYSAxSHLld1qi3urVnERKy7zp8uKFkdr+0s3uqM5k0vZ
lGjtsxMoFxP7fNs5EfwXIWPlpVPkiDMDXETxJEOIIJbU6Gur2F5SyjMoaUfoDtBv
WY+3Fpgw5UdELs9XyliWIRPKY76xbrF4939GYSHi8YRpV4beXGfV/3EfyircfEgs
nCNqYRXZYfPR7QOXxudckRAzQl7P6sWec5nBEsry8ljlPq2p+SVr7YES/ao+jKbu
oAwhhPYP3AAFIGXiMulYG8GBR2awpO44EaKjmqLfQGBjzIkPR6U2vSfdHzj4jo6f
/1kGL4IzpqSmEP5c7nziyyiKjEfuJVpirIeUxTJPljdKaHcehM7FVHUccg+qvwDp
5AIydBf+uXz4TJx36TrQ2xPuZTls+6Ys18HSyXilPd7UAY0qGb3gHiz7SsYtE5R0
VHtt7ozNFovtUmoOYsA9fWeqbkMu4ec4srtiufy0/JmoaH2LIqU7YghgL3+vwFIR
tYHltnbyhyCYnRU3QVTj7/V1DX2cmQsLjopLBLmq+HX2+aed8z5sXMmcaxGZUHKj
PtGcmuFOElzoA00qxj6oYwBjM7jfNPp2c+ks8EcHGAdQXCLCBWXXtAwEBK/AbE6x
n17Y/8KpmU4lcgdEwciJ88K2DrB9q0CTwr3G5JCGajACC5T3lCa0GxZeb6yN4SPW
2dlWZqbRLmKS5qgYYnvskDo5u+HNiYu1D3oFPKQJKSBKpmy0dN3FtYLXsmTijvmK
jcFmbj6YvJDSx44GogfGUqTwFG2Iv3aDpCaTmljbWfLaMm4UjCCvqlz/W1C7KvKu
gQwaE/8apWuZBDDTOEJ5iC4yzMEBXOtglz4U4HDQrXYo90+oTjFByX+/8s5W/5v7
JHgAU00z5bBSvGPYgGAin5uAK0Ql6iDClwSrqgadyko5ZJ+2gsyIbfMorXN61aL8
BqVxvIsenifq8TUUxLLWrUpr7xj5IDwSLL95/GLxTgjiyqZeOiHpkLVuAm2hYygA
ePqgtnVhfFBMjB8Ijaj5QtDVdOBW+JGcaETT6ePwGlJHgZubysG3L7+0WX42VExJ
lk6PQfHF26ELRNp3ZpXhKnR9bnTtkrMz7ofZJAGjqiY/aEAOPEkzaW7YDqQ7puq2
u5ax6BJMKporcztqOjQ5Td+NktSCwDpMgzEsv8v0qPL6Yq617phRaR/20LDRc1Nd
qFue+ssvjc9CA7jHLahPM4kuq9zPIjSbG5eCLW6l3dPIru9XrXivuOlogzC4Exqs
Sh/tIa4P8RvYtradKOl14PxOn1GwIiPIYWXq//u/BxnhYpyYepJsezN3tlLY7kTP
DI37V75Zn8wajO72MRSgF7CddHoW1aoLjZ0Hyf+8+vC95OfhjgJjR8+nD2Suxo+v
B3ayIMRYRblz8RdFxCB1wvF2nFSPuhmAtGZ6l39+qC0SdhNt+InjPmFPSHW2+Q1N
np4FQ6kwBlcJJ2GyH4peOb1mQWcUalhi6fdX71n8xTK2Oz/a2iT/HAUerhlwKvql
N713k9sis3DkzYw9NUGbii0A3xN3qW2r6IAoISbqtoIGA06NxULOtkcqxAs0dCzg
xYnBe7vpq8I+DPoJ1HgiugbXLgBFzzs1oYTO7HB50TiFf3jW6vV2amMv/bSl3OCK
irZZO0+U3ZOPnN3aaRp8o7kc7app5dmj5qDcIdVr/JbZVxdrA2/HUoCb+GCZwKJg
B/u7I8RWaj1tRjmBDofNzz97tmcjSSFdWOViP4qbZohxgEvNMQBg7jSiyhK4I9CJ
6hDxPYYUKSCeC+CwvenT1KXOlUvOEY3iA4e7AlLVOEDtIGCgJBmtAb1WJ4jtuWuB
WMzEabclI1rqZ6lzQGhyHOmqhNz2KGTCZO4jCt379vBt91POULb+4MBTM/krqCB+
hPwr3iQWE+KZVYs3xMvRn77SArFRWAi+/K4a8OHggT5BrjA2oPtG3jPX4+zfkAMP
fGBlQluS7O40VzDoa/plGXdxHYOtQ13Jxx5c0RWA3wp4WJzE6JpM6fmtAOmFAmR7
qufWXQMYU3hQXrlvRcc+E3ebrBUefA1FhnnANgfUeaRA60GZ8ks0pF9rXBz1TQ9X
rqNhJQIiBhNHm6DxA+m+86AiUieNmVZQVr9FD/QZIq+kxQWS1QE4VqQnSQUKiIFe
M/dVUgb8csS4t3QRY95vNrBk50G9Z9ZKUbx4faj/B1njj6VL1422iQ+x7W5dmmQS
TI9ZaHwSOxprrgT50mmGiFJjOk1dcoVpH8pJ+PLCBpWpydlUeOolsmhXOQ1Szfjc
Qbt1u79PcxEM8UazCyoRdhbatV2a78me8mjoHPgQFWpEO4HLV6xz3vJygATF7u85
eM+HmN4+TUuRwYLWav4ZedbY8y0DmDONuJKMcmWwc9zT7P8Z7S6GxLNVZtnh2qvc
NW4Ik2S++GfNQOAnqM+vzGWEHYSi+vYFyRwrY36iFOP/xO905ZtxgL4bhqVSUyUq
Cx5mrZhD4ZAOv0+bSO13qH4PpRWpPIXfr3d4d/W/sd03z4LnZBtMxOCVOh/LXosL
xkxaE+MwPQ4Cz2yXR2NgcfogCMk4m9spxuRJKsgQX0dL1VwWCDVu2mXa+aWKLF0m
9R/FGdWvn+oeGL09DIld4mDE4iJIzkfEJB0vRirxMBLnw0zrO6yh0Lg3/NNpSLKE
ap8tZifuuhreK3cGOQfp8a3wl+wJF8XjSzDYhGIzB5FCv2mymTJNbO3Hk0F4ZUZW
z3G4Ud4jwRVSvDgT6ZePOln/gyEDkdA/q+qzPG1iPEy/924C3+/aID764eMHTkFo
pj31sPnbz7gPl2I+Trtk1msug4RvsIkDmAQqPpOjtcELr35uxv21edIS+5+B/LZj
874PDYQsz6Sd8TBIv88UUxzP7VMpByNXk6YdwknDouiYg2schQZPZmf1hDjYXtj4
XBEXppatoqDgdIO5Vb1OPqqFr7xpSuLU6zG82pELnZIdIaFriKqD+N1vm0JUyaFo
ORkCSLIJ3HQR8KOLApKgYkRfppmxk1hsKM0TZyJr92rx5mCJWKBvA2wAY4of7Ics
FXISUZSJ/beiZGM6Fy/cwoFaSHE18Tq1jOI6l6+xLyqCF91XOsXNYai8/OPf2THR
2R+6R/pdyrgFRjjD/GuMP1sG1qg8f6G7DbDZtNJo/kbs0095s2xmg76tyWHPHZxP
P5uUel5E1VwTE+ebQJs/v02O9Huy6shtG7nU8iApVnQtk9roX9JToavBAzOimtTI
ubDh8C8zG0z59YwAkzvPvGA876rfMYEYqcgN/aMEk/nYZ5ekr1vqyvkgCac+JCD5
gN4P+F9LRMNSSgTQEltt6/yuf4BZetheH93ZGAZdLwpFIOq7TDd1b04mJOXoxQGA
HoojT+NB2zoeV6ctraCtUc5c95yHfGjQZc64Odi0NEgFI88tg8m0ptGsdz4bD/uS
cNSMQjqNKM8WxTFKZei++1GkeR6KXQY20eU9NR9JLk+bYmzOsexVTtZ6RxLgjrg8
f1nZnfunmOCBjcI0pDr759DMXLdzAZWwlofLX3xmbnb37CSmk8GOKJ+a83pbpGRi
UziBKBBs9RzvH0DeeAKAH8xLPIQjVT1DopHbUKyYvQq2zWN/NwxPEfSeLpk4wqbX
77ROSgVMClWYOZPV6CAG0ehHB0Z1DF2r3L/wojEbsVsHl1OqxCI7V0kN5jrxhOWl
r2N9DyNOXVonAAOpJd0eFgWyLQiNTjehlkMUTgBBY4xnEPua33vhdUzZBtjg3Lp7
f3scc6VL/RyaLpVck6U5x02pO0HZUMyMuhvyJeOnf7/D76VuQN+PvPlhdEYsrDVx
QfEJVs9V6cfi8qLvZBVd1pCsiELiY2mOlizIsKWEVDnlv8nUm0AEIMuArAQFYRln
ObXeLWCzqqY6r5SQi7SVHZb0TP9t2VJKjmZmL/yGPUawIMnopcFXPPz05DuEUfKl
VY5CgADc5ZdFLzKDLn5lIOZg6l3C3p4bQ9qdaR4LJlGTGfnhxubqfas80fyBd8Cd
I+VJ3V2Qfpa70f/VrkrSDRmrzOuogrrmfd6IIl9JP7Tj7YLmZmfgGn55nrFgIsYU
Gqm/ONe63XZ63IKZ8yEZ6BEIy8dc88BNMl7WogxNb2+Ar8tFfC5EXY0gn+JxkdQ9
UcsFuNRZ6z8mVWArW9mmFRZpMo7no7wLQhpdVb9EaxzT+0foLs+bZKCwoA3bPkiE
uDpsnpQN/JknBOoOPA6Yv9/fAEq8LNtEtozvYd1CKpc3i/fKsnU8ZvKK4/7FUzgr
PAo1CzYz0tRjCUDLVdUsm7+ykwOOHczdhfkFHmRG72r5nFDxrJDRh2GnhnGuZD5a
zIjnhE/e70H2QrTxj9D+8f0eaRxexwq4a67/Div4T/CUYCaP+NOFIRVxulTsTReQ
I10GLFQyrS4qGYS40WBnZiOer0o5RwznPdabCbC2pg8mJDKkC1YsAzRhEVT2He0x
8t8XhKz44e4iaEBnpoj1Lez6R7APtfIT2lRNVmcfWGnjEh1yLiq1t87RLOcdZyJj
E8ELZ6Z0Om683hpEy2l6gYQjsuJOJdXsedrkVy5zIff4er62KfbBmq/5HPRkwDuh
43i2fqiqnR3n5ePVTLJmw1aaEvHX8f0EW2CbrHZCD0xV2w7rk3SBl6bjITWirAo9
aFQE57xItytu4+Eo92PSnECG7rjZH2gWjgE0lCc24jQvFc5X308G3T2K2/fZv82T
HGSLLX9uOiZStdXu0C20+sHMLbb2yzf4FlMkTcSz9LvtHMr4NP4OFOAbzDz3jt3w
sEOYJdAf39CMnQycg2it2YlTteo09cHIiOUcbz6MAmxGas1N01h6WpVZQfBYrX5r
YUS0Bx2aeKScCrmNygwBwANKZG9KoW3ycpt/7yDeHH9n6oM6+sCXqm4eS5IDiL12
P5bkNQfwp3yN2BCJxFz5RRHDpzu1uQBYwpzVwcG4A53d5wvEHyU4+GZUdQeAcIeO
yCPP2uxyQ49YjjZE2zqd/q3RRm6oFImeRZaSEaVMhU+pgG9BkOM4axoPmbAkv8hf
VfNqT0lvW5rQCd0JpqwNDoEsZJegH0+1OngN3alvv2Z9VdSQ+7o0JwddKMTrhPn0
sIm2DXE1qAN94JqEAiXJ0wDwkmgMzOaN9vDnMpcGqygnKa9kM99ADXP1EEQqx7fp
WX3OuMOcTB85Rod2rxkRUzdlwBRVlYINzwJ3w3P+ddWO+hJiboXaQA2ewxZ0zJR5
vd1SoC0s4/jk44rsDm6wxbXXLJAaz9856Y49xNowZWU1wgTtOQ0SnmLZkpVP7qTt
tLBoWUK2KA66SU7Tuu500M6POA4gIDhiozi1QaE7t6CKBxhpudpx+cSGUzlQTYam
OD5rBcwFulmy68v6rQZl1lWVNQCl6gjj94O5kwnEdXnUaeO3t9I/j8nuPsIVsdfM
fhYfrOSja9m8GYFsoQXsxHcoqwxrwWURuyBYkwk26TGbjWtXlSr4fsyn6/U/5Zp7
INDBY4pQlpBIl2WJIBPwxCoMnzA8VJ6ASHGTqHxsSf2UvDgI0oddKiIWp6Fudqqk
e0g8ezi3KsDSJGPCoUYbcG53IlqjbE2HZvOo9xJSJZooRpcv4T3BTMNJXHmrNHVT
N+bCtg35KmkEPXIBmSblW6PBQgG+FQ6GbqTJ2YVNo7xuxf9EeZ0e1yXg8bIprhIs
DbOFdMhjJWsw9l3iKOVJgg7AfmkC2SgB5b6TxVqzbl62+iiEI+MrCNDRtzxove6H
rvBUNHofV1/bp+NNyurK+KL4IWlRPwGtUxwYH44cgFZRjENQaGYgKk/eEfxy/4hP
924kVMWQu7zwUH0h+ati9v+vmvqJSunmAR0I01Er7cCRYKu3kTsrvMt/fyFjRGFX
pEDUJzCLW4w7ojfcWoYfsefQnga924ZQcMYE0BroxLKb5RuiOzNxO4rUZjM+yGla
ziJCc5WGS/oszLhzNxzFXrJZ8Mfj7qr64vFMqoQEXBpxpioxITVoID96U5vbeTCO
VknGN+5zzkOHMgb3mPg+55bQMBcLhK3wpjuaRAOHeuE/uKxqFVcb7s8y4SAYz8TR
CRCWxfCDKYIurhekLe0wq0tueiMyR+fNeE3VT9OR7ruVo88uyC/ZgTKuF2Tfu3S0
oB99sMMeUACK+/7zWoVgnvSetmS8NRczJHX08wKNCMwIqbgvcVEwiKOTYbcK905O
PPyPYW7bYMDHpNBWKr79w9JljjMveqgA0D65pBfmUTEpjhbb83PZJW3xIrGWaVZk
TDC2jhNf5CLpvRm9KNQ6b5vC6alpxS47+ISXcRLUK0rPKUxaiZYVFVBxs/lK3wZt
6pFoKT4PidDpGeiX/tp9h3/1MQximm4f17y6gWKE5zaUdVWYc2gauXn+V6Iya61M
RmW3YbjrSmyCVyvJlAjgI8EnL47qkkwMhL2wjiIUOw+BeYK/nRJozIOtewS16Ngt
m/pTzeCc42xDAcbUqWfQgOF7I7we+bodWgAHZxxmOTmFkSZ5r/QUKBgGlfM7zooL
XpGXJFs8OyBmDob/614PWarA7mJv1F1zwTHucKNS4gh6mItPgX3O9hCWOBoYX0WH
m3J5cSjeM5RJb+g0auUiGD6njw2WnHZSpdqWPQOLrxoZw8lf9Z/sRZ2R8OjSdBv6
ebJJ3YwauINUIOWsPbPZaX0RKTtfMBiZoIm6sNgs/DF22mLyJREdOnIHsQiShs9L
Vo6RPO8A8hjOGcKjnysjQB9LxTfe1ncUk9xGpemYjRXXUKP4lZv3kJLh71IV6e7L
LUd1Fr7AJA4aceL0oYJzh0AVAd7waF4Y6l7PwTBPsu714CprGu3zFPy+tUKQnKwU
tccq4YJxXcunKO8Qt512TI+wTuZAxnXfx3YFFYiaFtZaa7xEVvRG5b15m3GxBSYm
Xx0V9B5P/grKBjx07teWomZN2fz21UkGKskKSYBQi42El+cbZ1Afz56V02VQQ+88
YiJ+cQyoVeZf/HWwu4As/y2pzvZctdh/MOIR7CIbkqMULiEzCWcby5mjAzvuADze
XjY3Mx6Qcy2dWCpVMerJNPj7YaNKw6ikXLczBxjda1AlDzRrIW0ozM6KuPzrWN40
onQ7kXYiXqupWW+IpxDzIlbv3xC9ZFGZkd3hATXaQlI5YD8+dT6n5OH+8wMzay8l
0EsfECPHC+yCViD1exMVXB9WDf3YNOb7oAWqERbeLVAvudifsCjbs3A7juSnhUyw
WvyyaUeV+knST5MUPWyGhsFkQ7nWMGve/nMO/Z4Hny6fTgAl794atQWNGW1OD7gX
MjeIW58CZlgtXvdRkref2z3/nL7wxKOBOd3Qi4MkefXxsu/MKg/i5kI/3BFhrGx7
PPGKaJIySWeukLMv57LZk9v1kLe3hzvUmEUlP21en6vreI6bCspYaP/Neumg7HM1
2h/yHB+NFI52KVXzwxFLTsE44YYjZxvZIXzzyQpCU+l6UBkd6n1IDkDPcysXhg3b
zMk0yq2VhpSFsZlm9XaKIvlu8LKy4ra9lvbxFLfgBwsTrHcHGe6N0kbfTJO5BYbU
d4VVHVrE/jVuZJoCdrbe0ZBYiZ2SXLIqXQbXf7eIBttTeMpDpo3ZtaBHarpBJtSd
aDS/xempqRtTCS5jEN2SqawIN3XbUkh5XvyRHgWG0AQwDJOVHdWCCrCIyH1HWbTP
jl6TZu8Jb3U9uadg/jGSoZMC0CHew2iCeXwYrKrGMAJx8plwSRg/+mvbQ+TM/Mqr
LOdWMBHecGFVPLEZFYflbwHo0HG7kF9KWCwlvXcDzQb9RKrvyWbcpbKZ2gXNXYkE
KjY8HR+hbDi0GPEH6Ip/mHTMmgkr2pUA6jIEqNrQhi0thM4wppkpWj7d6B7HBxRe
LIRcm3HvIoOduexNFw7MWXLabZDSkET02zcxKuje3T/Jt3/5UxAX08can7ZuxmXJ
qx/TXx9zvC8RWeeCs+ub8wonZtwwS5rBcwcx4Qv6Eqlt/l5MYW1agHNq+rA6BzI+
KxHCAUQ1dnlzDw+oGb3f8Qn0dIlmuT9PAMy8WhFfCC9MvNN3PVVd4HWFiKscK8Iw
YD7c3epWxsrl4TDe5dxisd40qRQ2SuAro6udb8qvhvS/Tb0kGZ7gIKflRVq8lqk8
Er2jdEDjyF/F1U8F6oqP6mTXLjuaAde8G9hodfdlgYDhbQAjShScWbzzcJADbJEH
xrhOJv03fmT9m8zm0CU/sb9sXSHduPP1deQTxJylE6C/Ry84Ux2bmn2HGLQpbuP8
WVeDNI0nQusW3wH2lI2jpYziYefuCVDCa9QcG3VEofCzDvfP1nLCzxy/Q26mDlAZ
AtC/dhJEzrAGAmYYZvyVf5kFYz8LuoPugzizHKXKea2fodyn+TLC6sWBOj1FN5zR
wtE6e+1IEzWeHe7HWx4Nw93vqeJYr12IYFfNtLwSGNlGR7vU+Pwmv2TwxG3zmDpg
npv/UD96gSnzXMBqKMGT8mnmHkt8nFQrSercsGFVHvPODT8KPJK7J9d79VfPl6VZ
W6lMj7TwD6Ky51eghQyU6NLzJ+4PqVEgC0DUh/Sst9uq21K1at/jsmfNEUoZwkd/
XMnOMKiHeBxPoL6sCid95DzNOE7ENAYPa0Q7H9mjbRimLXjrbPddFwMHyuSFuVW8
AEDD6V7DvqMwEYKo4UctqSo5/eUgqk95I6YYasHeGNfZXx3fauedVcoAMPLMtn9X
H3LHyKCHqNfucd0wZJaMjnkf9Xwz6Vxpnd3QkyFbhNpOSb13j6OeBcML+vTim4ZQ
UIxtvLWTY88a4Yv9w+y4fxXPAv+jzVmboTUBNwrgqBUDfje4WuQFbQ5ZiUgFf9nl
ypTJdH5Rt+nX5ESBs9O43Y7fmkUKBwo0iiR8AQEG9pLjqsuwNhmBTA+a+fEQ9VuD
Q2HTM21ZWdV6ERqWolEPbvbtTxIHVo9jXEnnA8hl7KxowDzVv9PqSeEvZu+4+ja4
flsFdyeCqUeuV5zYTyly4eDtu0+KqC1TfPE+2SJTvW1URquzwZiev+AuFcnchIO/
0SF4lgZaZxhAjT3/Vx2+OudOo3z/NnQzRbNtvZSZfmEfiZk2fknIF9DQ0HzDlcYb
jHiRBx7D7yUeazl+SXiRtY1lXyA/GwCkppsC4GBW+wJYHjxGooBYZSG2lUrSZ1G4
aLkNsx2m2uAYns5oaWxsFbbrI0KIts5+lIgURI5+2Bjfg92zzqcgtnQ74eoGRTIv
VAtbh+neadTNlrWDNZQXjNC21LJSliQJW/J2Os1UXWUyljSC3YUQLIC5GutAuvqd
ixSe6KeRo677SDUdu4GcvdqxM7B8eCzpP/8gX/oCbZUML+O7CumZOAadh9ix9a/d
sQdjsibJhEBPn0k/jFC49SoiNBJniaQ7riOt2AFbEbz5iLzQZ8KyOe3iKyL18S8L
vhW7zXG11YYpH0veCf7P1zQwBdJ9MMIkys9HIJhkW6xcrThXPxPK93nXGzhpz9Tx
LqiFsLIOprWicxBPSbPXyPfi7RQcijNPyY6R7PrINflOxceQF5rbCy2SvS2A8/k4
pS3ECDgZfxtWp9CaYKA9GVxIVai7Ou0XDn8q1PHbN0HIjLnxTRLFTVzsK/GbEjwO
JxpT3+5J2gEV6rkm4TgjGaQ127QNyfgx1Jtmp/7qeAcIWLkQYQJQjWrTd7lm7/Xz
oz1QHB+FOJgCG9aBCDsryRtc/ju80pftP4hc6rbiWJzeoH8fQpIxeUTuvLajDa2C
syNuOUsgsOh3mX9+XJk8CHeqGpCsdYmQ4OVOglR34C3adMDZ3BKmuSjuLY/rGZGb
HYvS0Z4/GwaT+r/EQpwiwXi4iqLX+wnijDIaLGg5r791ace8ngURVtB/eatQBYRK
cEI2bZo97vke7JBcjLHIsZQHs4aEpnOfnolcOotcPrrkLRbRVVV/vEijz3uK3azK
9F8bbI09pN+wFEISlxFaJNQ5L+XisfpW9eCj31LlqWqUj2xGPaW0k1XIthSyY2ys
XW+eI+065MA0MzqGC7Qv7vgDIVymifpwZG1bJd5/ULMhxA6mrEsr7obtqhJ7z0wP
3N8AQAHKpC10QdRLj276/H9LaEdnrPS+hoG26vFSy5Evd91p10rvjDOVWXAXvx1B
6vqKJovl6pGuhDotNgQkovvSjjdrxx/18S7o/jwu5FmOk60jQ49VX8x99rlNOEbZ
2ZNjZ+93f8QzOuxvsfEskFnpo035SU4LP0VLh5jKplK7f2/Qx3qWthO8TUhLCSmU
FLen4ecQtoceDsSmFXqeWKkvrQw3bu+zs+bZzb40MQDykijS6va5/SofCIh16wAD
jWYKCc6WH4YrNBdCIaob7rfnup+R3/i7/uFmnDRXeQkWJ+0kaGcbA36fUoTQm1xq
9VqpzEiy/wRq/kI1JbQxgEeC8hcaVgKvaGQiRuFGwGSe2HUt4pB6m7vgQVPsOR/R
IkxbprPXkin7hW2/qDf0dsWSbkS3hQwgexnvAS5+r7zSZoc/cy6VK9CneVlyfiKJ
mBmH/wutXU6kFWom4je3KIuTVjAKTt6/xDomnaZgSZC6t3mIuivLPI01s9EUOiVb
ppraZ+OmTrXCw9QQeu89gcvO/lzeIXWZLgWbgf5FoHhb5aq2JfgZ6afc9p7JQSUK
ME4BZp17gtxUHsnc7vInEOwAayi+7FtjQUp7F1e7402Ox56yevHOW8MVFrhHiuWQ
QyD2rR0WcNUnskOTVY+lln40WIgSgb/jLU7R7MBxX2QXTo0EucyGswDNMKJmc0k3
/5JUiBk7yDyekh4UkieDbAsEFqN864/zG6xLu5WH1QhHAlBuzXccP5rYstDxxVdV
XdbEUWZeYGGt+MYQP4D1YFyZNQw+nX9HjDkAlD+YL2cH3gk/jTJbQrXJ52pg6Vgb
aotqBuTF58tB0mIDuM2t16rcpSRimDh3MfyS8QpZoDKxUiYra09P0I9yizzY3OcB
zZxeg2X3/b7nzzeHtqB2AGD/X6IPhYaX62a8/2L+azVP6FrMGAyiZ17TQZwIdBv7
ZG3hBosdcV22MVEG9CjkUPBiHhMq+thvDY6SH/XomHuL51bNi77wgX2MQje9TqBI
fAxUTqbLM4rYXFk0FoSR4W5R0pVhQ9meJTCNoBe7GKGGukPDiK4NIsNd9rNbc0Ks
Z+h65yPoTE+a69JMMghGb8TCh4p5IZ+71gPBM6uWwA1KdnHyBjoEbEOJ0tSnFNaT
7FmmvI7QXKbYA9/YPhIdeS8nRwTqJoAtXogDbGI8mtddfC/LbHvlp6SvhMWBiKai
0SvZ0qHcaqql++GPG9lx9pXFwQcD5X16tFVx2sBG5ncOV5nw8IbmFwhQ1NT6NPGE
x1qUBGHEmitKeF1QyPg58G/4DGTBDvk7bTx1FRdXMxzkF0jy7F2Co7N6ypyyGNzT
Kj3bmez3DGDSF8UQiSBuUwElg/yFF6VIPVYoLRyFsgEqNguJQUD+aLvToZpdmP/J
g9qac3skKqJ9VtEcxix72v+JkL0v8ogO8SVU9X9SRdFL5kQguuE0svHjFa3hiIbx
Twi0697Y1MS5UDxiELSzz2/qvLRC6wb13P6ocqmTJC2Ds4u1UeSpUzjyM3XV8Fub
KzSvm9RWKAerjRP1f59LgTIQU3W1QAL/7gHuZHYvsHL8iG9FqbBy2R5YgfgWjcOj
tIS8Ckd+LvUHxZWKcXWQ7Zhg2808p4WxRVpQlVAaehe64N2NIus4VpOYgJEvniRZ
rK97rPOV7rBs8UqE0zJlxOHhU0MBfZQ5uZod3S/HLR0rFgwZQvPyqNoNWFHbnAlb
IOgU/hZKQq1S488JCu1FrOV285Z/OoASdnpmS7UiR1cX7roema+H1wxgxC6jUID2
rl0RZEJ3EIozY4QEFVgatQJLEyRhDJIHewP4Ji4a3/TeG0G9WQBnH2xkGxfzZG6Q
RdBDj1intJ1OqCaabAeSWEAV9MWZGVXHk/kyqwo58YhdMTajoNYotLqTzTXn6v4E
pInHcUKxSSGJonW1d19AVy4cRLz54WhSJZZrhFVh2hYUjeO5VzuVDA0IKis0T0y/
e+TjmouHikfK0iKaLyVJmvVewQ4X7Ud1LEtFVORXBAqcGVMkKPOcMSx/PFiyeoeH
N7HMuB281u/erk4orW0zyKBQtN8vFD9NBtEI+7XhvrXhd3DFzLzwWjqhzeguzqyy
y03Nc5UqtvkJmP2wis1lN1KuTvAOiIZllF5IMwWgtGoI+kCIRpN0bp7kiYqgVPId
0EB4NKkAvSbkhNyWnqCRzqQCvm5dPDL3YPKDEA6XTHFCY5RCwz5bDy04n4OuoKNE
NcO9dIOLm6q/QNhtyvc1jFvj82EkihDKH3KckHpTny6F8k28Qa+4sZMxYqslJG4i
pm+WnAxyXmC5oVsx9z734BxDv9enVqggS0lbx5DKGQgFDFsnVPMx6ePwNI+XYOja
Nql1HCxnvRFXcXFkVv3rrkz9toWG4g3YD8Yx++FC+CfpBg+G0atJunFR49FFZjSV
KZx50S7s+SeU53FuehCV0eMPTWjcgz2oGRr9/jNNEC0DwcSjJbxs1FkzFS30sdU+
dw1/fQ46ioFPsiu0C9acdb9S0ChhjiKbXuxHNmiL3ZcbxrqPnp5XY0uDbCxKQhAZ
C8xmLIliny3BTirhkX6r3j8pd4pHep9Cp+sYo8sAbShMDVdWLBI+HkE9qT4vDJl/
Qf1vNou5FyEWtYoIeZuVXno+oY2BgZt1DoWyXdd6y9mtoLNFEo+0nHWTsMqjpvZo
z6ZVLos61Jr1s0RRAWmBzy4cvhM+8Zy6ac6lXw4NBA8BBiz6LIlBE+pcXppzkb27
u3RllP6lhsO6xxz2L2sSCnrqahXE0yBlbVccl6CKWf1Kl0oCeo6UOsV0+mDW4H4/
tULXW16bqdxB1NfQCXbGgTGAJEeg/8JHMjGfUedLMj63BCH5r/9HyEemum5CA46o
Um+QrrC/FaiAFHm6Ww3GR8kHfJHKJD5cU0pNiY5ML5tIeB9kBgPIDaiSjZTUxoMh
hPT8F7AeA6RI3IH6vuLR+wSmqSomcVN60wkN4T4BzlMFFC40BGd77FcdLFAFdJSl
WWE04NEXyFr1rfO2QuDKOVNBthpLA+qzHcY4+L8SDfb2xsnB6yUmmDwi43fgiwJ3
ICrKbgHiXzgrDM3HPZBH+OmwihVlqjdpbPXYknumRRFVIlIpWLU82AXZrEtTNI/r
bg/DcTo/LapDsLyUXQJSOxl7h8v+y76zC6jkVMHXLQx3zeqcZ6DpxWlq16EyCHwj
f+ONNEkwycoeIVIGMAOfsVAq92Xm0rMD4mU5V69VVifGNRtN3VQ+ZwXRye3Z2O9Y
moePOGlv2DG6T0fE56BTWyAWK6TsGp8ZWfeK0bZlOq129A+2cZVGshlNdBBgVpg7
Y/1H0T59L6qYZ1fzDc3NSD2+039FjdoKh+4jOQcRW2dLXeggaq6gXad/XXdyL4VZ
YEx8qbMiySYgbdEWwK91oVwjA0hq0uI9yjGSzZzyGcM697U4yGcXI2i0xmXq93QA
WDX9ggeTtWqya7QuF1F217nrjqKxIfZAF2EghVtQBa9vA+jt4zng+3LDNkwRcOdU
ACxJeD0fbauUPnP68fSFGszeG7wBinAFXOajo5iFLdAD2HbvhKrp+7WYPjIBmkEj
HbMc8LIIf6gzg25SOErS4q86NvjnbO8irb7wuqCJ6RMi+u2nL4vSkqfAcDqDs9CS
QThU7czVw4IcpBN9rZtG58NETIWr+9cAIAFXkAOb6TrY3BUWU2+08M25sW/czm0E
t4rGVRne0f/ZeLAZGDvsY+I+cjeVBmsQyEJfWuUcfFTaNFIYg95hnbsPAmr9h+qS
YZKJgHGSh5dkZI3zzHb854FM/Gxze0U2Iy9Xw267r22rjkK4QAfk7l7U2HmBM3qq
q9GT+om1yq8T2bp8DPURpoAhmmyqQT54/zNetoZAfHkPRdyjQ438i/2WZpW1GpEl
yvz0dJXM0ErC0MONcvFfsQY7RiXk2LCf71U1B/h/XBxr4aYcafqtgSA0VFt8pMPr
WgdxWup5MeIc09R4CXkqWbv+idX68Km99kvZfxB0kecMEBRYY42Iid2t5pPCanvE
LthPgKDN5clxKC/y5sB5yICcuTdRnwnahQooZe+QnYJYv+PeKT1AFJtHcEPT2Spx
89+EsoaDF06JH6dLVoFhdL/qYw01sCALq6gGZZtt9ESoOxEDO5F3O+IvKZtqdbzJ
C3VGp5UBomt+oAPBVcUtV2tCQxKB8q++B6Tbj3U+sLI5H6/77orVMSuAhKLBy7v6
56AxCTxkVzbcKFNpw8vA422AC4M/HriEnZp0fM5bjDNcmHuzaJK97WoDnz4zOK8w
0sZqBeDhQStqi25YOx6zXpw20altdy55YQt/oq834UVJq7rd5f45VgDQ2Z8Atsxl
UbYhp5HX9IHp8/O5WKkjyOJ4Sg+ZX7EQUsd4eYjJZ2vfo9wh83/zz3ynzya2+hSm
AumRbz8BZ3A0wFlbaR76HMY2v2Wh/nvnbGpr8rz4YopixhcoUuBFdczE5zNq28KD
eVOR3/u/ScUKLI8wmBK5S4TlcF6LsfJStLg7sjE6LS1Z8sdVlUnSlrvIME993AK3
mNOGnAifYtVNuscoroHcWPzBNcTMaV7STbkqttkX+Y+JTZ22TRupS7pwTvVdZF0W
5i1Sy1PKjpJOpVdmNyWbJbdMNINCazn4tITI2C00NEgwvncsO/Rpwe9C+QBKq7x7
n7tIH3mXB6/ljr3Oxw3OxknXcmd5s4hU2JkOqBzhwCRndjg2fKZcYcK3BzSAvs4T
JfNpbaVbPLksfBUTCBurl4/qhVizH/NlZC6QFyKL5ZEy85qBVtqQbZtnNJHA/pWB
rLqsR645o8Y2pnQum/2dYriIaMNw/5K+DFy13hNPz6S3+MhswdE9mz/auvG/X1a3
493tbOIqa1SVZqJeP8NuqOdjVBtsDVgqCAapT8qkZNpcxMLasOiP79UNmXO35PFN
n//A7/gOHlB/oRMiBv6cS7GWzcpjakXlDfjmhVZsWZGsNNI4hD9CLlCk3LlnZhXe
j6u3fvYgeoaJUVTadVvaERu2EqVxntOBIfCQRcnt7V3xbwkSZAjpebB0tCA7fBPF
9LrDgYmrwtdkXQ3rB/dxckBJeSSYnnck0YXSXpEdgX5vlz+hLj/DGZCkhmi5UQYb
O3UGOTIgOboVNFAqF/IdoIAgv3zxx0qsQal3SF1Acn8VeALL9yhZnpMz3dnk0HaV
fjgPz1Sp6YIJzpPhQHjYfcC9f0YjlHLQ3IdxEohoqwQmeGYD45gR+u0eLrU8bp2q
XtvO6TR/2AVWEj51yWB/fcPjZsdbS2lIYs9VZc87/iUlW8xA0GDWPtETozHCe7O7
jQ5ASkXZXhuC5Gf1DoEtOcq2g+D9FCoJrPIYVgJKoQVFX9K10LSGlNT0hMGydkn4
Mp+c/MBkwhfVvPXeSbhWYRmDkSPRmrh//6biEud1HgwKJCz6+A/Q//omog3sqGCL
eNSlUoP379atKUC8VcUnHPQ36zkE9xt1Y0KcXnlyVd1+2kO2WhEjE8CGlVyneUkn
z5uwbZggkJxsFO4/dQExk5zXRFcmJ6Mn49MxcEcvuH4WlTHxU9gqpNiyR52M6oIA
uuhaMxGiWvgkTZGt/AyMlYK1rq8elONDWbwZUA2L4MfQDVW1oXkNLJvZYNH9UExc
kBtmNLhsIcckip6YcBCWkRgsa/ZAoaLsRkijSw3cyA38pspzhmnMVtjZtm5L27SG
nWm99oq6oixp8ZvTQGtbR2HIDUUvkz2/iasfVoUFpa6HVP8G3iCmD2NKSTVqJJus
4JmRtnBZiC1WSM4LjBCbgz+hCAsb0UKoJ2z9cQztKBUl3zy7hzHkZfaXJ8dO6lTk
MRzpWWDbyPLI8EU1qu2aQAiCYUualWF03WfuGHhm6PRNf4j86Ut8mEfQ4n4Mlro4
PI0b+ThdMxCYt8dc8LpdjfxF+QOxZ+3g6hattWw2iCTXqSTxp3sEq952RWQ9XiA7
12IruLCv8cADyeB5I5iOcXbmyyULNUOd6aHuTzIvw/4nn+MH4Sgp56eStfRYiQyo
Ji21Z7AOxSV2wmoeT1eCNXwL2Vm3y3dH0UFq+9kCtgwHqXS8mRGGsdzoUFbXmRXx
eQYs2WEPjhcjEDGZfumomW1CxPigDta07oLPyYzgRaSibGPgNCBR7JNIiwCGlfAH
qQEOjUxd3IC/a88TobpZWfkFE696XAlOMwp2OLQYcfP4FQFNUts3k75Q9FrRW5tF
BL/f0ZHen6FamLWAiQJR5thVq+IvQgeENk/mwQ2Ilboy20wuLRREMtzPdNkfLW3z
tYKRkvPIQTkLTQKmYm5Q48Hrmp5Ht6W6xrFROc19T/JS3/aGdg7ODm+vX8+2JrZw
OQ7RfZWnGVplvZS2H1FJhy+526ZYsNl4eiAJL8KPf26i0AYe0o+A8FE5c0whkRTF
6ZkFUL477BkJeaHP6HX5pJuDdSb9G7j1sEG56lEZA9AOTsWJbKKpQKDJEzK1hcal
nndkPJ0sdkKwzViQ7BPTQwGF09+eJkG5cYPCYBzzz+XqizyTioIX7Ijr+/1a6KUU
572zLyFrv+eM6E/c9Mu5hOv4fQ/uSXb9iy1CmE1IU96PcSeGfLFwEnmnkFzxvZrL
qf/bbymjfzeHY9YC2yOAbVIvlkTNttTYVIdwGmLFGzOeKU0mb1cV6r4LgmNAEno/
Exabf7SDMOnn2Xlw8o+/yXNpvz9l73mwCM2WFOJew4b/wmq1WT1EEJ8PhC0q6yxY
DLSdncnXsj5LeW9bJrZhNwjaV9fhtK8QcQCydfxAeJo3CXIIHXeHC0l2pG4xvW0k
YqVBShULKqCytYxjyjBOgX4MA3P+u9PfHP6nLaN/u9YUbfoZSUDbZ80mRmZ3dgh5
ggzDx4Dw0jR+DTzKNq+kxKSp8Gw3b/WC2Qk5kAiq2fVn8s+7UXSzStZiNuhyMJT3
6odinS2pR6T2JAlEBMOHV878YF3hPHgpFoO85Qqte9aIKfUvMFRqOS3u8Rs5sL8H
1NDOruxfwVq+G5/By3N2scrG+JK8IzJds/VOu//TeA1IT35KJ1KJF1OXIFW0yIT8
B+ajNazPSraUCqM2L7DN+83Eug0btk3qbdAC7DwFZFtoGUKOP/KYYpbtmQxsDR1J
uj5GUcGoEPyMsA7FIBh5JFZZ/fhR9TgaQP2yusScRurIhu+0v0GrKGhQ3A6K9SUY
MCfdK7X1L7eHfL67IT2Aak1pSb9XtR7tHat5YHD1ToaCujhPd9vVcoghvcC+Ffqd
5YNdPJ/Gx5jeEHkOAPvKRmU8pIEvBjZ5XEpJD8X6nQLXfwxNiXb/lfcG5dePWLUt
ENOy2UU6WiSoM9QHDP/szsdoa9k/4tE1u+AYwkAFHK5wY5HW0t7PgUf/qgJp+D6c
bLBqomz51FaLWOwtDGeMYQ9V/rYiOYHsSTx657Qm0tjMN1Kh4h0s0yTw1UBNHyIT
tgdWiwhQJbFozKlMXc/lSdD202YGL4ODBKyak2kRS0uTBkKwPDcXptN0IQ3KaOnW
jLPhZhjlJObZ6XlBVrc40wBfwfPafNPjXwB6AifdHjAZSW5oCx8WeW5S9n3Iw7GV
K7xJFOLLfg3yPtIbysUxX6mI6ANpW1bko1LLAMRq3KNZnzrMdjQGVSqW4w6n1+AS
MmmBa/6jsocBWwvratu0zo/yp+yakUzZwdbnJx64rg9aTAk7i7tiUKObx1FV1bR4
JP3a6y4v6PMAZH0BoP9Mp6azFx4gPQFLenLNZjYhUiBLGSi443sQ1j+ffmti/Ej9
r8ZGGXQ5QMEErWOkoi2zXwP3EUDxxI0bdOhTG/q6cKH81X9BbtQRmGAnE/MgomFz
nk4PYRMI6x1tQgkjBOA7Uti7dgHrDM15epBsdLNyx+RacPLsezyHzQtu2w67Eq//
Lcql4Ywy25QxlkypWRM62wf8XKPMsvzs/sLQlZFpsHPCOg8UTyefsgZuGan1r1Gi
jJWCMb5Xhn5ocDNRW1OEMlPuws9Ep4WfwBlMM0/OzsC8dD2gFV/bleE/l/2iB4Y2
kNiZZt/ctjf8puTydWHI3YfmCfaGj4EjpqwL53GR3cKLjL53Cge7lDE2ThcBk92m
ncxvr3leNTl/83YWtOmkoMCgkKw3/mAyJrc5lF0m8MbkQ9H5mfKBjOKeMIFXOwjo
hwGh+c8dJjrw7Bl6udo1ZI2PHZk1VrNLbXKtlAIJ0RUyoazAhqCcFO6MyWrp4q9M
51+ONbyKl5OEHCRZdqZvu31Zh/AFvbprJhY/7KSf6VlVRud3N1H5UfEW1keD8aAX
RGN2cHZCwpwI/4AWtgJeaKYefwTgq3yKG7J9LA6Tc4Wzc0DjHWjxQVdNrVkKMyRs
ugiTzBxdavAOxixXUNjbbvF1cjxbn5ts9gRV7TwZjzzpbvdX4674PyetVHGc8yrr
g0hq+cl7qHzsCJk4hFpU+qg2jmcxzd0JC6Y/3VDsn42coMW0I/+26G3Dyr0pg7no
nZGf9+mkS7l7TAY99jcfpDz9I8Pu/j7pW/7fRAy42j6JENSTaGTRKhG4kHv3wP86
UdXpRgmB7vqJnB5ZrAxOMq4Pl1nkQRZpTxMMDHnJYjZcvqEqZtuCZ8WW2Diy+X4v
ep9g60bkIc4iPT0sII1f4fhNOhE9/6V3MC31cpWGxvIOvofE3OWnAPp0mDghGUwv
6C4JCfDlj5BTyymaIiyaWk3YY1P2Y/nzxPuynaDQD4tEpEc6FNPSa0VyL7+2CfKS
ytinp2xO4zQtiTloYv+yTcyI5v4Pko8Rx/nBanxQEXUqXubKHJmYFQs+XAuhyfDt
NCiSJmrIcbyEkw87XL/KTYTbFDtgJHBj/ZSS8c24aPgoQBPByHInfGpf1h0N17eQ
j4bJOaiVIC5NQv7qXFvHQMZvz9iwTQNLgfLTQh0m7ahCtrK7MWh90/ubCBE0T02j
xmp8VqJihRnujZrjC1Or6NTQNYT/ipmtPKyO14BaHETEHm/EP5zO4h0gFq1Ht/pW
5OInquJnefjjHQzchI2fhGJRdU2Q25ELJN0ZoSFp+UeLqYrf8fryracNmdGJNv+G
h3oPLf1OiHq7yWJBZn2tGocj5wvtvxxej5yCkqK8FNvwD+wqOM8LIBALuIzfMEF7
3N4d56ZTmd0O5unXCjQAcv6MZINPxZWkqNWRyNADu6mmbqPCzpn6xXWN5sqP3KMZ
ff40HZW2Ub3ictQI+AOooKo3AQ7cim/OWOMQDpmGVNYKRy93HxWuBGaeuByFT4z0
/3bV9Jx2EYOXihz36PW42Y7DTh4BpM9PXxFb4xtoL5Th+CC2kzk59Bme8iwxbbfE
JEaSJak39xNpBFbySzh4zbihBQmGe539u44x30BO+7XL/Za563oeFJid1khmz1Xx
ZKOjWUSezgMsnE/xrUZyql/UZbL23lF/cP8FijOg7MQrpZQnNTe8TXoynpgqmmhU
ZFqdr6Iq7OB2/SDqBt7bNTKEvW3IjiE4vcJpV17YPuPXwLUfq9BUY1ccCidLnXEy
Pq99sOwTIjpcp/wF38VkfNMKbb71yZknN7dztJQdZKBLDbYAE7X5Vvopvl0AO6PC
mg1GLMNx8wHntSIhzV5gocDeRbJdJOrAB7domVdKEF4PNdU6uM+No+vEVJmI/bTE
DYuTVaTCrX3VVOWg2EKg5d4H4Y9PeCwRsutiMObVQEUW8eD1J1VJpfSMPVRqUbJY
PAeUEiBZZOi4nUepp9IFFwMVZZs6mGWQBKwufwmEN8suQ+XBIM1tnlxxL6cUPNNw
iWNSwb9DQKNdDkUEZFK3+lxvLb2obAwlATBUK5GepQoySnxVkeUekDnCm7oAkfbV
wPwo9N1Exaaul5xfGevq8+NRRadcFv4u9bskDV53G8JFwziBgN0alezSyGJZwxya
CqL36OGtH/dej44X97FcXMTJqcxD+8KRevm+t+un/fXE+sZKAvXQ4MNYTMyOj48Z
sNWDShzJD6GvsNLm8kuZxOQOxTfvtPyBGbVwIesQqQMpwlxc12O3F8u86CeXJ2My
3CeTjIAZeX10ZI5Tzi5UAYLf/fe4j5qSnehYXycWFBHh+pjh3SOgWP7yg7ju8OgO
U8rwm2H0d8FmETHrBI+ZNblMMKPCk5kRo1CMQHJkukSqHqGiu6SFPr0Rdz7MWY/N
+o22EHhLhUpol/IRd8T+JqcuO3Zqcx+g3ZJwE/33kB82kCEvrv6d/vnr2/uXyH0S
ZNKJpWeiY6o96vj1UrpWvbUFAv3fECJaTT8mIN5jGdcsudDtfXteYJ89g17UFR+q
UGKUY7juL4KM77WeAR1IPQmrnEufDNVHosO3mTgYtrv2CivOk9Tu2tgMC2nycWCe
caIIq3BOTyFZkled4CxB3kRYapPj4H5R/E9Ei9EPmVRp6IHvdFIHdRKCm+X8Ep8D
MXWqGCV11PC+xENdSyz+ApkqDCWywestZYUElhAgl/crG9U+WtijVPhqrMQElmvn
39mhNhVOXDZVjBdNbNZSIkZ3EEsWj9T6O8+QcKZoumTlASKgHC0SQuOfCsDOFfLR
nHJfLjcKwjSKWh2RkIeWo/dkK8v+pruCz8NMXl8HhIdD6c+kvDGzA7n7QSEOVZTz
YtTydRMLMVYu1YS4TL9ivdF5IUew53uY1vqUjtD85dw/32BjbUZiyfE5BGoT6n5M
Jm/skENvbntm+PQITxXLm0Jo3Py2nkGKQeKlWT1cNufN4t2cLBi9iLRR2lSoxPTc
5PRYn2l1n/0ckmAuGK/KKhDHBUcZr/5HwIg3Q+4WaleUU/4qNCSNsABykLKDse9A
2LoJ5pBzkj5Ia+iLQu7wxPCG6WGWVd1W070cRaHeCP0v9HoBfhcq7mpuIxv6jqpG
3619oMEnjBPF28FXciUba8d3ZnVG18gL11jo9q4hN640zUcwRHVPeZ9lmVFwYIZv
Z7YJQJLX+KZBHxzL40ubJS/p1Ji+q8CpgOXQ5SjccEhF/O+AeIqLiQMaSLqqy9vH
QKH30I9L7OgQMjQIuyK8BxzGuBxm9179B+KEoMC7BcLLJgVvgZqDsxARWioeRt6C
n+W6Dpb3KNmoYbwr6RKjFsJ1D8152FdTiBHwg6Pr8PgD13hxhz5n7d5Bi2ct3afh
tafop6MvBLe7h9utWMt/RW3r/SwrQrNfhw9eL3r9+kayVJNewqoOfvGVbWvKJ1wa
Td4HcqGm94AGjlsk6d+ovzsQUiBObOsNQxizI2e4HpyLm/MUVcCXZ7y1dMDrbd0K
XiRwBstzyfbkXuWE/uukPhzy5Mz2arOuJfQJRAzLeGGkmyXGvOVBDSSVkTxDkqSi
4iOXj9axdLak3WZnyy6GItJctiwwzH+vspn4NBH7uOX+Iyg1veSl2TSLlBhifSJt
y403mKklGdBgRdPv6nNUcQKHFgH0LvVMK+kk6LYdLVwElI6Bh0HfB75CpSI9Dmdb
XEzijJxl+NT1nZ2Ofx455dXQY3aSxNyqdd3FUQb/ZyYPqeqYzHYvqEyoOzcc9JPa
5H0F+S76PVCtoEWGa9XHsbdwvLKc/3X+pzyWFIEni4Ko8P4EDiSuEO1nrUWBNth6
Et6ZY7VGeN8R49ET3HnQGojbko3RsrLSJqO22UrA7UZG20xwiBJHB4B//lticJn2
w3AdXGvuglXkkmHpyIulo0O8URbYe8iCNL6gQ3IAFrJEyTAVoQTmcgc3QauWakpG
XXtkBIlHu6Nb5He98L4JIee5kcQrUcHX4b1sQW/GpcEoEeJq2HX80iXwNNa0kqz+
y82bdSqkqDsQx6bGsegYM+TnO0rATqXN6x6FOLy0BCbkWqgKthEnom82Wfzku94g
u+lEoB61PMsEKItKYBNuLbsl0tQWIFqktoIb+UWuO3EDwFe4A5PaOakEoSUOOPBV
hQPR7wGDq/JyMRCSAJ+2Aohv2EtymSeu/E5Ct59DJYHGWGv5X5jtLA5ZAJetFDqP
5FkNEuPJoM6gC+YZc91F4AT2zZVFNqoBLAulkexvU8ng/raXhI5NPDwMU8HM91ku
U/yKVBLJxe2m0d1QyCL35K/vGdQeW810H0LsPObLOXtU109OcJ0D8GqAFU45vWpm
zuYc54T38lwWxUXP6WjkBMK/t4te/XX5ojdm3GL5wUHR/0rOOyKOxLZ2spa15CII
YJvljWzIFg6exXBu3q9+O/mYMnSHShwvV8vlPuRQAhq1kwn6ZtH/qLUSuWL71WzJ
M3ymHPD8+7WosbomUgnKgsSi3T/3AbBsKIGxFm+kRuL4g4dw1ALYAJOOG+rD0OfD
NrzHEcfnmUiiNlvIT6Fy2E7MULx6ihSFKoQ2Fpxdtzi/8EpJd8awudIHaQ5wCxr4
YAoGCWePbxYHcrVNiT+RjQRvCGYS0XY1ElSRsL9cqqjAsWEaxBrB/vY+WE5yX44f
cYTcD3ceg3J3c8OfKKJ6129F91wJoMiQ+G0eNW+CZ81yK3XgCFBnzNXLsOoOK/S+
5cRz7S+yE/phbyStd5/cfxeJ86JCPv26Sq8jEfPPvV02atwexim4/KCkwfQkrBnn
RKBCUUOyKcO2xJ5hpknAHZNRZAr4bipeysvSoTIBDrdUWtOL7r7kcxa3K65BacJ+
+G4fPyQUJT9qV1r+w8ruw/Bjr1eTlX/E/8GRt5GZopvSla7KW/cKEeCv3QNJG8ou
MVmR/iRWNcXy4PoWjv8c0BjrYeDrlc+1pkL5sDmn+ZS5DuaYOdJM8uaGD6pQn6C0
2WtJi17OqSYuuQ40LtYJ+/sLH2rKO8P3zl/UG3dyyOMdATbpnHErQOc3z1RKftc+
/3cGIMCFmaWD8kRoYaRomGcObIYKcG6ctkMruZR2TM7JXrMVLkBRi8U2sv8ar66Z
Vc315wL+mVX4lgyrZspF7byYm+6JyO645qBOptU++whb9W8FqUx9TrEOWfgFUqQX
T5yAr5r9lFiWs9aYjWIEqiF4s2B9XVgfZMv0YPho1raoZXS1FQ3HpsSH71lalye2
xnwI8yQPy5NZnKkUzgqNheI1eCdDyZu5CiSGzpPwYC7Wz0x2XNueL/QqarIIa7St
KlxoTJ2Fq5u138ed+oy3463PmDTupR9vgrCPcZwZgklfilxXbC4UhSUzTE9F4sdM
ayhqjXHdsgK+l/1ZDAbJAU74XnXmOr5zM1QDmdQkQe78Lxm/DXrsvDkH8/x1/2sI
H3Ho51uVKhPpDBUICzBtB1v+QU3Thr6H/uTLskfaSeOfOcGt0cQWR8utgxrN5Q/l
0G3aHwBV+57CwIHfwNUu+50R4k4psQoA6GysVumbZR5nEKLljXrm+7Y0Rz8HCrFt
G64xJ9dpearOgs3wBdsfsQyMe5bFX345o2r2xb3A8bZWiPYxv1z+YaaB6vHGcHCj
A+jTlt5L1fVqRyV1mxpCAMy/omcW+0no+UPpT3v/fNEYdQRAK1k5Su7C1xC2XDbK
t+5xpAAP7IKVzMZzmAJvifqF72lMAZUyFMiy3BHDZUy+m61WLhVLuttdUxmfdrlS
ostScsXkTXUFI+UFHl06AXscv4D0lOvOhaOkw3BuIm4zYzPmebApEZVPhens5alX
SxLyqUXdVjXAOObFCHZPFGLySxLHbmzNeDty4jJs7H54RDHODNKLpu7psp9YNe2i
E1Z/BsVMQI2jggUcsZwx0VF88Rm04dcvrI0rLt1iPh183ua9Zj0jR5dSUIvmROKP
48npaVVmZWO5UPAZrl4FGn9y936hF/Iq3U/Zc1Xsjsytw3+bxH4dg8S7DhM99kAz
8rlfnLiBO/aWsv+qVMuDkJAGNnub+aUlOvHIWfsXhBKlSiHeoOhoQHR6zUP6tvLK
4nxMA4XFmY9Os++zbPS23xM6n6lg7ZzhBJI3akfR7gJZx6ak6JtAnS6JJ99cxlp+
LNHL3K4Lpd/OMFgWF9z1wZhh+r+yPUPxQkF+CAwf6GAvi3jybHvaAr98OCfXb6fT
2OdP4PsEhgCsPTULf7BlNO5auMiCCPnekI5IcDXcD86nbU1NS2caITnRXzX4UgNI
topA9yZtd5LQ3bJpCY23nMvm3IZttUdDmf24dyCx+GaQONi/ppd7aqiveOYFK3Cl
r8IarAeBkz55MejtBSrJPihqn128dhZm9tC/GI9ja6bdX1IPUL6hY2gtA0FPP46C
TbGwz9ZqHwvUHn/hFFCEaB9lCJ36zNRIt1Zm/s+g9dBbUylWYME7EZXUbVlnlCen
OlAaMnq40oJNyjQ3CyftIA5qcyqDBfJWaMFFXw/J1YabahHsC51DGR+Qr6vlKosw
phTCCg/xPM927dmO+v3CCJLKzeE9OoDakHoB9f9SiV3bZ+p2GVca7Mm6r17zhxzQ
zDJww6iXcumyhwdjCs7IKb89Z99HSw2m1JIxu3RCVcPWmWmoKY/PYOXXt0UfFDdx
Z+siQjswKmLl3cUKWD/3I/UOxbrMwWDsIDB+R9+pbiULJa6u502fDwrq6wF6tdJA
Jx6Tc9Hx1KUSg9F62yJ0s+m2bqUDhZmtOkB5WB28oMx4k8RZyBtym2SH4AcQezrO
FMxQ7BYdFbT+vVVKp6nKmGYLWIAcwduH8sOx4omdwgj8O+OGO4LrIeTG3VYPsgoP
sUDcdmTni/YAQRLjJTnj5dQd2NVirQc+yQVKPdWnCsp6Ex+twCfJr8tFVkTkJoYx
F9pAw/fJw2nIREtAndKL6Ux/G5E/Fu59PjP7u9PH9SjTXZTSa4d/vHqGxuAYK38q
+54ZsBBAcSo+VB7vYgcLfD8RIE/ZbtU6jqbWKZkUlk2qgBz3waJ0b74nJmMytKM8
Mdb62gSplAws5mfVZ4wgWpjxwWEnQZQ2CyznFBFabuAgLFJEDwxdtuWpRn5/htTq
7pZIKyF8BYibUmefVBa1u5iObwGBBvTIdKv5zbVUQoYNlt6j7I22qcaQpSu9oTEh
yKaI4bBHs3EHhkalDK8XJ+Gq7alnbE/R31bfnHGGf+kstZwnIuWrvZmGM5J8EZ9L
To+liWJ60I+wzebj1154szdRAEkEGAkg9XU0JCxDSvRkyZB8QtQ7DnmWKi36dd8k
x7rEqvb5DOmAA7OUUMd4BRbIukmDUCN0OnjNoY8c3fsTwT9EjDaVybKBR6BMRbJr
0PhJIqDLXAz+s6bmcAZHIcKRQQja90rwY43En2gKFMUVF3Mkb9V271MFgn6jMdPq
+x/rqV04AqYoYcr3gSzwM/2/NQxmDx1ijqRhD5QfJxwtJWpr2y6IRQaUkuaoRHqY
vn1Efd3pYtF5D4YC7KXEA/+IhqfwOI2+IkNh6qOoQT9bv9G7BZrwlZye3PDaOa7K
Vt6QYykeXZFWUfh829hj/lRbmrR2/gTzbfiM4v30aGMgcoINz+YgA66UUpaTykPE
1eGpHjS85AAkUa1j5tba+Tm2cUsprIw3r/pleSYUaxclZyunaj3AsNF6YxfxXkZe
GCxD5LaiefZo+NtJ1JXldlDo8lxAWz9zlEbBdjX3f/Ptlp5fPOLI3Ds2tFAxtWeE
QlngzQK+rj/u5QmBxMuylSkBVD2Vb87yjpx4Oeu4QromVCPhJ69Kdw40cVoR1ecO
7Lo5+iVVOAPJ4bHRc9N5c5ssvqo4K8auKwmOjbkeQgg6UkbJQ0j1QAb5nI43ptdt
26+uZkXdE30wobB+w7MHqbGH27soVVdscku2vBdy26WkwjibWzJQyZQNKjwzBCxm
ikHcJNPt9tdtTlwTPc9iEOgZWoOEef3+3FPB5kUCsBr4Z/ZwzCqNwFaxXVo7mCE5
niv3owNtdDpAafGD0MscJf67vlR8km3C0Vv5Uy0oNb6S4ZZvweeiJDDVD9OeNpGd
UkgmyKX/XPg4jZ5DrzhdoIO09fvpHB5D8WaWSradkgnS7VPX/X/Vb5DpCVQWSH84
2eTHXI0RbUay+rruyOdi2x+atPHxhUrHVouf9Tp8AImoEJ7cltM1sHiArAUc4XxL
qKFZUiKLwYFXqpnKXKQdbFUtPurpznjE6ta0vLx57coqfRIug1S7cALEqIXz6kcQ
vrga16jEB4XI5bKQvIV8Su8sBPluy0eYBX+5f807lEwepowdqf4OV8aSBcLe6iPm
BouONMUQbRQsyn0WzbX25XBZ4MX3Ha8ekjAXOysVb+6eYhhcKpT7+xq4T7EDQd5i
3+ET5GewF7QdotUoKe6gO6+yMGuscm1wNtg9PelUKn14LWubgG40EE02j7wER4aD
phqQSAG/SmmU0Cmmye2Wfzia7O4Y2c4qagDSmKMBS+9lk4ioptPnRKlwbwy6jFII
yP+JkFoKdQ2nD35h+HB4TFoLyC6u/BlnaXeP8T5ipjwaMQWwmkQLOYgInDPBd3WC
/UIKFh1WRPOEHSLXTl/FMLpx6Eeckgez8vCH1VL9Arc0c/e1P5An6D5ZCig+CaGS
NCAXRW5oehYxeS86wbKQnSXiJyM8u+QAl7TzuuMaEiYh9u4EpZoYuZUzWjX8e2WI
KRw15iNWig3z9hNa/eF/swbugRMR5F/NZ0uqZugqKgzpdSh+/a4Od2Up6AYYMEDO
sMowqYJoFPlZgof4vYfoPDtq0DiX3afMutZ48CkyxZmznqZXQGrTk7JMSDiJ+p80
1p5fsx0dvy0/9bdpB+KrYyTpnrmcL6wRol+Y3yaY3Fv//2LyCYVBB/XkSeeIlhSo
u+MEA8NMwlsDXCK/ycrorvRUdPm15mU+6Rp+FaPyfIdiT4BMGbxTL4wq7elwD1dO
pa2BQb/caz21FLJeZ5GhfGd0dPSUCweF9Lv2vYkaCMkXDLZ0mAjrmVAnDu9sBW6m
JHR7UwaR7BmXHGZ/O6H5zXd0gvV64Yh6JQbxxDvXNXbdlLW466DHfZZMCyZ2OUGd
KHBKJVE0ywm7jClRPxasT6AyNTzb+wOkDqN4r51BMY6iLb3e8SR5pdMFPdoiYdg2
0r94nqUB6tNp+L6DK6KPysnOZie1r9v7rn9PVBw263ZY4y76TW+eRUDM7JadiXfR
MTckIdJZUJktu2afaMPWmvBejDgHT51ECCazsYHMXgygAOzX9aRMHpeb/M9YwDw8
yMFc+KQyHR+uPBfynM61JJ3J7E7EZol30NNZrNqyuOxNzINXGGGrF3f4Qtp18f9d
yP+m/Mq1FtXwxJkngLrw2KRHROA2QxrQbgoG+ue38ZpcR2HGYKuWPyxyccYH1WXO
1K0LGT8tTa3gaz6I6bq5hRR6tLpwJWdxnDnKEpKxRvUYoAO15OAxAw8MrqUn4RTh
znFrf6JhmZTtQsxEpqPb6EDHib7zncNqqr/hHG2NAHYFvEvz4/QVYcQVskLoRdPe
7RpOfT4gP0PtlKFKMsAcPOOewITc5FjgtND67WarT4sQuFuCDTtFbX8Cu7a9EBW0
+xCkcStDjyDnYt1tLEe4g/K3ZhMMbg8RtzoCASs2qbfHL1kJ80e/Z2AtNyuXy5rh
dCRAgcgrEXxWjHvcTSNWxRLEGCeXMYL6ttUl8RgAr2ISj8a0XBLXlJ72dAdGSqun
ghL+ZHm83GcYa1Sjq6UdBOUZwukh5RGeWXxyiX6bDHUke1WG2ch/idlMI2DCUzv3
cAxS/YhTIJPu0apbefb9nPsw6ExJVJpqBQr8X+QmusnNZJcs7GAOePcDKavLNzcU
bR96ipXTkVLEDOiO9v8sd3L+O1PVtW9Ps5Wucl+0gweT0uENNU9R4p1A3XiDzN1G
w3v4Sq68vNqSdvJ+ZegXisrSDgdObmyGmcaH6MFwv9uHOeHlO6a6ylazxnpcfm6q
+3x/DReirAs1UEbvybZ9273uj85H42s277vcp9le0gqqQrfATM9D674M+w79DSfy
H/cjGHmHgRMZ5FZXVzNvZ+JHBG++w79I6GdEGFP5bOET2TrhggBVekEdOp6wGn+H
t/6g9ga5nbcGswINA8w1mfd4ybAWKaftPVNVST62V4bAxpJilhU1PVFZZExXyy+2
JfRVraLf44o9wH3bnGjfxoIP2vV4WVoF9X9J/ImwZYYY+lU7m7ODl6CJ1/GfqVZm
AJQuMxzsuxxJsj4aw5fNz2lSuCvdngmHAmA9x7YnhKsAPm/ud/8L7zf6ktCRJvFy
Ps0ViDVDPZBwy0cR/Lax+/zVB+SnBfxXv3bZ7gxEvq+shdeAHXrewc1zMW76l2aF
uEFWy28WG30cNkJmoiELWWk+6C5uzRCqAP2Twt9LQ2xqkbpRqVu15cqjdooD/RnU
Pt5Knfthf+RsCHOUKf8gEVlGmrhhqXlh7Yc/mwH5UvtC597aEht8Z4oUmc9ahM6f
ZxkYQx1L57jpnd3CmNlX5xuk3oDDatU2Bd6G6koV5U7WIySxOgSK+FdVJ6gfBZce
WgG8pTdSYiuYqa21vLd1vzwZh7EaLUJXmo7IXRd8TB0sVfzutt+TKHz0l//JopQL
e3+5Yick1PjbIJAzsRKkT9kNleh1OUkRfJHgBBBVoYkhHU2bOGQjxXRxLlGUwOrJ
gvJdRKl/a63lIeJ0C7j3SaOv6zYgWc/7094ybsYhpt2xAMLxuU5jaaJqzSAx+lNz
ZUT50Mjhzhx5pVfk6GZhI21wAXV3vkKreZdfuqIWS1m46rmGFLKEA7j4BGWA4ieb
c+HzPdLrv7Y+lWV9nUhA2MDCFrHubZYQ6hcGn0vnYkErfSELJrlA5Ez7ZVBAlNp+
h2P5GqEF6AL3pSC4TKg15WBpLf0vnqXEQWaXZ1yYiumqU7rTF2tKLwQ4RBhfCT/n
+SF0DXJI0CTWT1HZYrieiDZNP8YVGs6B+umDJR7g1V+fo97u/6+CDKOJR2/3CyXj
gnto/U1ovNu71j95iwgrAjoLENNQ4aqBNFIN32XFQRNLW+aVt248FfF9PJKf+ZVv
FwLmgQQS7+lPpVJKtXL6UCHyvGj3k511HCAz7D9KRzls8DxBvFOyHZew2QvoM6SY
ssOZnzj0i6Suix6+M0mK/vNpCVlbOvAfIw0PvxjWrXj64+cBvl0Z2D85qoA4IaXv
wQMiDwTqXJs0IYrflYqBZSCUN6Sojf+iT26qnbaKlv0U0GLExE5Osu+b/9dCX6lC
rOsxCFbAmWCW4JQAG45/pZ62kK5Bvsuw2hr/7+/GoH4Q6Nss34LcYAFDBcJGX5oU
p3drfxZZtmPhgexSFppMEEiR/0qmwJrX48cQ3K3YbRYfu18JVPW5CfrMYBMC7PKK
qkYutJemzerimtNG85OsD8DoctF7IqNEnbz7hkMxYBkBjVkvJeeXb5hvqGhgEyHA
d1AxQgU1mMl2YZhYXbssb96KSd3jMgAZ+kdnghRB3zzuGuBK+V3fnA8B9cUYiikO
3vEXxfgIPwgBoQxPGuRBw/JLgZ0a48bLcZBDgLhZ+SvQ9OnwxHoDXGH83EIlE1cf
+q3Hdf46XEVjPC5o5PdFkK0kerfHfFqAlAtp3uG1NTFbF9UDKdZ75VXlITb8R7tp
iOpfsPNUZNG21Qw+IMEr+P9ZFgqU6+IGH5a8eUkbGCk3bt1TPvYdsmpAWkfcdrd3
yGIdrR6nwZWV9edeA+Dv+IpRCHdlPx5D5qtvvBQe+QSIwE20go2qouG+kaBnJnuY
Zmg1+cGu5jT4CJjI7QUD8Un8mXSkNfJaYkbZweTB9rrAmQod5qW8F/OrSTjqBGzm
xICez0jngSNvPe1MEcCaAjZoReIYrc7zvg4rl3uRON1nRJN0xnmCw/J5MRZLpIJt
n8kmXteI/xHBZk9XCZv8blpqRCveJKxWVPj3dfS1g+RqQxuad1t7AX5AbWfw2KiJ
u9CIQFkTztMppyBNBd1V2QFOur3u83yspmq1R6znFkCrfvU6xIuw3kcUckqAW/J8
IPHCQkTyVNq0PZegEwN7xo6qo3ZPleOtlH+f/vr87eQomvazNKZflPys7b3cmMth
yrFgoVDGDiRe7Z7F97CbHwugPDcNQ4avIybiycHxscyq1IYdXMg33s53xkpnz6p2
lxcVBs5fvTVY6ojKU94Y3wfNXAsuWlB5BwzUF5r+jjlJlUlAQPyePL/zkOOxocpd
R1Wlui2Oq4c/YPMNbT6/dq3hVLXOWkiUWqvP0VaNqQ3wC++N8kPOZQ0GxjEcVrv7
NjqCVn9c8bFdghuZ+aFobF1/2DbW0uCNCTQsBsrJ5/cdWjin3Hv2yFnmknkzkrnZ
ph8kbT5KB9vix1JzYrVD4MjJ19WCuSHx7LOmCFVYY+K8EJY3KcloyU4Q8whr2LGs
opQ5oetI+umfPE6K0yNfEgDoHQgDm/DZJpzRENL97Ga1SsEJHzoTWKXITs5gVfHs
3CzVDZdN6uWlLeCtSSC0+VZkVrteVWdT8th1rMn2eF6J0NOF5Cb336T8fs9lSmrD
KkeUp2i3W1pr/TCT+kmxZvupXj3AQ0gZ2zDilf8nmSBJepXIL+rzi/MNtI0meiQ6
8OSTWUqYy8oq2ND6Yd7q30bQD3I9/AX74tx6Dx0ZSanpbLtbvSfXjsx4Fzwragtx
pVHjhiAMYuXXRhFp+TetLXPdrf2jEFYOZ+QvqjwN+szcYU6u4ykpnujt/YyzPy0j
qTwbcHRxUcQEPz/ybWFHySl8BNJdpSYkFQIXA+TLAZPZkI9Fk/cysX8Dap/8dI2Y
Pm0pd/b9Pd8RVWMlxdH5OacYH7tHkQjOpSvS1pRD4nNlMyifEhFKsI8vaT1MV4xd
NbQL1+v/4hQIdlMqpwxbY1Sbar6lEp/FAa0I+X+Ewt2YYWg95MRtOoc7SD4M4vNo
L/gSEl5JhvbtVRn5zEI68bfBBPbqs4/AJOYSg8z81yQ9PyufodJazM2zF/YVuOC1
ZTfTisA6RxQ8/FsXVFWXwsizF2c/60iyZH4XQ5j0o8SZuBO3t73q441o4QaAP+pE
w3fwPqvzR1+kzjbKqeogumQ3AUvgM+jjp8Xaenk4bdtsmbgoUdRWDwGDsh6chwbr
J3s+ajeeMM98DKgDrpu9uY8+rdDBiCZxd6QI5/71RuuEJVm46cvH+lC9DboZSc/v
m0sl9Da5N/cbNsNgB1f65Zi8w6anFekXSLwT/aOyCkEvsmAwD+5Y2/8zOcnz45Pi
ZIh4/dAEg+QUbtla5YbJMEzK5T9v6b8INZ0qHSd+ESEwdW/qQSbYiWVGTDUIVWqQ
hvU4knZV/HS9C841I3L26w3NftwQRjeaevy5nrMKN9QO68h2zU9igV7j6eDYr5ei
vlQ0JjrD7K0/jUs4y4oha6ufg+fL6PKPlm5+QX14QNdTf7m6WIqvYA7YCg4xwnB1
A6GTwlv797bfkzWplYCxO/LZvO67hVAj9P0AC8Ky+h6iAhLvFMjJiu2vptHLddKf
pgOXvJcZtKpx8B85VNhrtDq34EcNVyVrXN2rqLwB0tn9xYsyjpVUYFHgivvXioE7
3E1hhbkh3BboWeXI8FsdPpBJthIvP3yQS0D/9IYAWF1b33q4R22vveX9qKuKG9Sd
Syz2r2KoEXD2+oyiSk6wgxMho9HG+Rhnd2kpQuYp2LydlIb+xs9DoViSRY3ebjTw
790CNX0I3qlC3jGyqPD3KNzzJKFlCQqqVcKPp6hScytKxM0GfKu4uHeHp9MG2cKB
KIJmb7klm+JynFv8ksZvbhR0DHjc/UFeQElCasaFdkBH/FZydejT/dT7TqrUaJ6L
152pZ8TtdnjLUqvzTqBlNvpbknRBp5aHpQ+EgoZ/toXewHVykV+l1qMSkXsn6gry
9ZCdZn8097aCiGvrwAHIaOzwbG+3YzCyhzUmb0R1f8WW/sPgIp5MSaQ+vEZ9jlzD
fikofXK39CNHcOx0Fwn1f8fohXwHnWMS3U56A3h8pn6I8gc+CCr0kQ1OfQgphX04
8/pWQxulhuBd23Zz1KnoHVriKOf4O2LwgTmSYwWf6jsY6oIq+LolSfO9UZeo16Gj
4EggfHtWFfT1fOCwc2GRdVqytMhuXNPILNULHoUE3J6iOfHCthmkv67dWSknA407
ANkbMc/ScQIFdbT5YqjZ5tDCNR01n8Dc5emc6I3bSch/pa9pacD3FunX6RzbFAzL
O/OmJG3R7SuIX+mPsqlzPXEqOVqTFOLrakuCnd2YKdst5FhLAUwI/0Zw0A6BCJhG
OYhwAO22OnaKlzXZzh0YUhoybo6blbIFECbYc7l2RbamO7ssYy1r29AwYTR2qZLu
OtnStglO+Kct6xKdroo7nMATj+uR97CePu569DyFYDxN39cip9Ie6GyifPDN7C82
NGM1meuLBw3bqFvKhtzJdvYGtEWGVWapjh+e6vysd9oeG5wPlzClx3P3l6D1Qyq8
pbY4c4qSKfpQAo39SHSYVY5VsCucdHZe3tA3mlsLHBw4N/Vs7Zm9HmUI0wcf3sUj
BAzbXoA1rjta0HK3eHLyPAbFDQoP1HgYP2wbOXv/DTAO6xHzEAyjvhk3w4Brxca3
ZTQW//4kdktz65+TsMwQxMGRDMbX8wPyvyeso5Op6839yTF+Va9g4blsN3K0Qq8i
TPuHHN2YbrkGPClK8S7DWEnFuZfeVe+6q45+DBo5ab/ezARqzuWbrWyeyayeSn0y
TXB2YVdH3bl0pqfX8vzbbomBu+R9mD0BPwD6e51y7/dGzQv6+flnhbWm15yV/UQN
/SmvbRw9+BsA1MZyeKdQqrYRN8+VHvhFcbAg47zYNxwYdAx4RI9wWyBqoXpwAi1D
Q6FCEpmpk1C+cZrk0zB9gWIgKn5oJgNch0GpKsPA1o8EypDB9ID41F+QblRR+66u
E792h4MbhWY/TibZh2MOizjW44nbqS95jvQ0ywHLcB4x7UcI2q5zoOrD9GacYTvb
iERC66+pai51QUCLTeGEV+mVEBnhkMFyBZ/iR3rUcgKoxT7OXMtG6faaX8sl3x9W
Okerpzoj1vwcenoSRGL8O23YY/qnVsPa/dyeVgqs802zTWrazAHm31kejjj4g5/x
AsvLFLwIkdPBS+8sHDnf16WustUaztKG4EJAYugu/nXqS5jJ/R3mOyX8NEPO4t78
iY9xyUBaaUBbZ0P2unsc++JA9d7MtFXSHbX5YJ86y6/HMyeNST5ZvHON3pxzRN3T
pIW7m57K5cqReL1S/ZQTlHVEXzVx4h513rbnUcIXERJWm0ya0r++pPSfZbiqs+07
gXQEzQoQ8ian+XuzYUVoPr6EsqpeUx+WhP3Y6E+zb1eI0pF2ayzA/ceXcLd+WqGl
E6UByPfsW0GZmSAwMHWSvUYl+J73wEcaNUdYgZ8jO4SaFB8HdC3NSljRutC6M0pl
pCR45HIhGLjUnQ9ysNabgPGo7QpDAAafREx3Ogd37uEnX7TxxxkSI1u/1lGOacSw
MFC1ve5hAjWfcSbN8JDO9yFZmtqCbPT9/rmday92QFUt3oam6b9t9Nothu3exQYz
hatvzVSjdyy4BfrxTOc4bAjdDRtMuKw964BAWqWUZ/UpXQOQfHLirScimigDPtg7
LU+ZIuBTlDusAU9zgDaTqY6wNVc3LzswZBt5q7YLS/z27Kbk0IbVKs/GlR7jC6wX
JLIBcgWUYSks3IXyQGJP7EP00950md2HtUVp6yZlwyNI2v5NEkBsCedfNz7yxRe9
3G+QtiEr/1zUcTwGXXQ9bO8mVskSmR6aOXpL5dEnew41N5zQ4l1IOO7x8b1YjE4r
i88eP4fzsW79BVDNsxN9BdisqZK615deczGgs1JuFUi2A9DdD8if1tC3Ffoy/QpU
oQQmQSVvvCXEvlRQ0uClDBa6COhQ/NgsJf96L+4AAP1+QzJ0G0za/TGcXinwR1xt
Fh4NVktMQ/0IiT/Fj08L0DMBsCYJEXzDnoMLJ8wzgCHmCIihMJEFJW0SGIlOuElT
/P9pKR4gmaNSJZJddBi8RIr7e/tvBmbP4aEk4lajJI8hJSjsvNOlFwZKvUANSGBA
30VP8zfjtKjKXKT+2v8LNRUGOHcpevCgQPs9PmlbL18iqjyDFagMWVNFXZBGmR04
4EAs3Q2Du/rqZcbQ3TVkW45Q+TizCpmHzPsLTSDbmTcBcGzof28X/cUlfaXJMGrV
5UzK8v3UDkMHUPz02kNDE3VDAzQZH5fu+Bf/D7enC5rdjlubznfEg8ArwlDtMZnD
XSExoIsuM0lO86QJwxTUPlmUnrw6mq8690V93rVEXF0ub7A2zsj30rAlGB2+WxKe
001fmtHH/EzxkypF0rFYMMEPm7rPHXrCkzQWQU0uUXzH+Eg3/w1SWCCLc2RNrtWx
eqIsRLyJF52hYD5D+47cRqR9jGNZX98zV7bsu8ElGqbo70SNuB+HjhAVx2h0PvD/
xgL7ppTKWJnXfGIks8jSAbVv36UgumMD9uqaUNU55G2WMpmLe07shIpyVDRvPMsy
QMjtpD2nqQgmy2RabIqoAQb/n4bhkrBfUu4fENPUnKZlnT++Am9wDbPGQ0XPffN5
PuBdeyGUh+vP1aM2p76EXdvn1QWMSoR9vmqn65dZVEt6F1tL6w5ZFVkkwbRSmWim
XOM8sbNAA7dz6jPOPfEgG5CeJ7I+fQWy+9D0/G0vPYa8To9JzPX2BTMJZ1A5Pzvg
bPwhne0LfI002EDAsQNPROlcgMJZqY7t/wNxPxDzP+970OC19XSVRSNYq6mEYflf
NuiQrTTu7hSMhhSNO3A0TmiTHwxaPvuysTPchMcpu5XL305B7hrF8nT7MEeIqFzf
kYIkuXivGJ1IcaQ9egEKLFzPLwjYT40jtzHgFvTcscbj5Pkq59ED1aqBnjkIWRkh
2ZHthqW85wegj8htUTkzvjhqKLqITMiFTcBwWLcFK5Cgp2D3TQOb+deFsjDGBphJ
SblPMhpgORqAFw0k1IrY+F0f+n+r98vZbAYwXg9YZCe8LO6DipD9lV7b5JrY6cD7
+E3huutms+5mY9qPmYpAqH8ErFnNg378/6qDIraCg68jagThjHMuDzLD8U/koVIq
/D0F9zyzerO6qnoifkmh71vVrVSukKX4rFdNjO6LJRFkbuA/xxfbZe8L6VMwwG6N
ZU7UniNJ3DQSNwSL6sp7dEFfkp+P0GLgSMJb2P8GUrTY8dkO79nzGSZ9O6Tag/fu
cpaPTPjSzvtme/wbeGClhuMYrDgAFdEp4nFRyZPV0Zz4KedKS+Eo09hW3/afF0+9
JFcZZuqgas1R5VQP5COWjhuXFCyHdkvO508kS0SRWpAAvYKUldYW8c7HqY6shTA7
9janTmeQlmz4DOPgISs6UcSTUpytONxohLPy937V/G4Gpo8YShd5gS+uDmDS48VS
IcPtu9CmRbZeBGEPdBrwtqBWhXXpD56oW0k0Ofg0gW2veK4AkI2gq54rHAqpDwr2
XgTXCDgUudPsotAECs7wGexfKznorPzP4F852mEnQMwGR3PRyRSZfFkRcPbc0o7E
rLBxeu3jhE6o8YP0QJ9HFBTokVI9MtsmFsqi4GyRqP51kto3uXSIbdfwN5xmoE57
Baz7QoiM96frbkSsT9/aXp7tSpi8H2e7NvTVjQfCQnUHs9WsK4Ie8Rg+eikbyGsQ
X6cH+tCz/saQSoGg+G5CG14rwKX5ZC1DjDwXU5S2pMaiHW1vrgdrp1ScT0udHmK8
evRnsa7Ad9z4Q+hZO+vpqDP2O+H8DzB8+JlRhwRbLBj2QO6kSnH7mN+aqhipZlHn
2m8mFTI5cztD0VgBSc0jVhfFvgumuroNgXz86w4MgscjYltfzHE1HoedAHHy9UTq
6FseL4OYgyCkRCPU9HdzCwiL0UaNnkya6S2IovCvm7JWUnI+LxBUCXAvbsongJNl
2OlKPt5N5FHVyXKxqPGUaWaW0/jNkoKXaE8o0fhJX0LlPyZoFNpJHc5YNZzP4NuR
H8Zbz2AiZlvAUCHpY7ElAfkgcv+WKCw+36hltdmPFSOtolTrudm9mOvcsxyyOoFv
MyyBIzZBfdETXP6QtBouhsWlxKqRWVwTod6mP5e+nBBZM33zGQ1k4/LF2ZLEwKGH
afq+dKyve5Vo8UBxWSP9P0PzMllfKX3GhNNwgis5vM9Ok1I4qgVbokAQKyXB7Xe1
JTyvVVzphSlr4mN75J49mTf9saDRTKEQYWMp4iD+xEyM4byJyciZ30GQ2jRysYFt
bSq2Oein6qPznfDI5op5ZzpQaYFwwsQ34nVgsLB7U4yQtqcIprZ+3ntgVdI3XL3o
LC/9AC1wgauMGvY6Ido8pUDvvjSSS6kt2zSkrqaHSbuIKBNbkLevsL4IblnBBcNJ
nUfWpAg+7IL4yt75lhdV8opk7q3s3XUrrvmQL6l3jGLfW5zuTW1A/lvwjR2DHazs
SAzYSWL7qOcfZiwuCVXTbupXm3ql45MU2AGv7p8eCrLv0DZY1yP5JCkntlObOBs+
sMjJs8CtGOUzjYs8J9KWqBGsLgqlUWCos3K7SpYGW3RDEJigmxJVxhCFT0Lp6W6G
IU3J8rNuTVuXBGcLZX2SWoxJNcnDxbXukxgh103rgVbcgEo212jwDTcyuxAmyiOn
rT7TkFbJWFTruaLv0plv/mKC19nDfOkFKLA/rAbBi4IKN1pfnWu4C8zRMznCy/46
lu7A0jQbMncn92ivvE0kFbG38OlUNaN0kteFTmo3s6jpQ0fICTanWqr18QT1Xi2h
DW/uk9PE7eTt/ydMKzQO4ZYwMSlP5BXcTvxPxL2IKBtQ2pMmjrhkp+cs9viBxj25
mQrbGsTiKdXQ3nGYDMRzVxt0Di1dLVPFF/JhYJYiFWEGUETEwh6nta9Ag5C6I4Dx
6VvEnPmUU1Wzw4SZ4Adu6gNklCP0RCLl7iQfsZ14m5IPKi2aGD4GMWoA2guBEof1
y6ytq2T6I7QT1/BVJHBvvP05LUwZqJ4wvUZFts/JH2vr3hTjwTxwMNay38x6ixvn
vQJIFEeJHKJULn7iJdpUSEE+Ecm8Xz7yHk+uKJmZT3L3X7zXeVhx5cOKT9hBhQ/g
nsNPx3YW8zcg59sVBmgGOt2LFxlN220I97YGNo2alpoGzYbFGH89Be+0prGz+m26
1kOoR07c4Q3Juhha7QBMsMkY0I/4KeVsb1nj6iwFPxUVsIcNIM50xwuY9oPTM8tJ
sXhTzVKmrV5NL1c3o5i5tOYFMIA0tf+Vcf/ZYY5pSQUMno4VWFVt1EUDuhO8uw8g
6TnVV95DGA+hMv2sRG/iI2wcW433m8lXlifU0SkwVTxy/cWPEA/9q+TtF0ha58BK
BVYj7lSxOSKufoyzPE5POf5pzy7Hjv6Owlqjd/EOISgiYH7eppwVqnS3Rst2ujE8
i0xRu1yw5P84VIPvRXtDjrF7QkV8NT1Ma4MDw12n3sISAaUKk9v3sBT2VCi7n+Pw
yyN9G9WCKaEc+daY2ug++uO1sOZC3V/oVQ3BRxSCGOCLAKq3kljfJMxFRL3Frq6G
mmb8hIIAI0Sy5iUXADClcuLoeaLnkTuLnQhW2DmzrblpnLct3iKKYAPt0pHjbD76
WqU5eAEDWNwrLaRvvB28k/FLIA6TtT4w/lny/axBpKuIHhckeI8wS3U3ZxY2l73C
nNhE7DsYtA35+u00Ert1+dVCACthNTZH45hWsW4ddefn23wb7/5Pi3qMEaZMbjBz
+IWcSuRDhmPXUmmGU5QzkV3vsorqNcY1MGtCiO1IwVwCLZNwV2eyXIEPxtXDFVD3
zXx8DZd1e8yotlb8GgIVSgwU34bJFNN2nJHnOjWw7HS8hAze8NuLr9RHKxbj8H85
UKVt19ohlZ9vW4r9ZvNdqf3emw+/nOuP2O9pOadHlPXZF0uVjv/tAvGo/SV6+PCU
U4XqJjqIYxB02K2r6Il/gGBstm+88PfbcGnNEL3x9y38IuJk+ysggJ3JQwS+1QL3
q54m6zJVg95M+zAR5BfrkqMw/1p1SlTFOywr5rIwlTbjmHVBcGdF4a/jk68VzOyT
0bur7ikHxuDlrW5YAqbp6oZWZ8+DjnXT/dpI4dwKGPqRWVCyaoJKGmXOjokRN6Hu
gZJwrqd7ePSGnumhRV8QfuBxqscb9xDjpRlZ1ivJgCEt+GhI6pSJlzPWzyxw2EL/
eo/oUbXpvsO4+YbL7PXG1KwsnVk1VzkWiBMWZcxCfLHBTfQMXagJ5Vm+kSz7XFSw
TiQppaUu+rihN4+PmuXRzmUVYYGgQLVNBOKAYxCg0mhhSBBShmWSW6cyXXfbkIGN
Y7ilr9wLIeNT6c+Zhqgk18VJq8UHnOJMRgsPlbphRvHRgoPKpgIvJep6aem3hrbN
3zQBLik0Qp03GqcLwCByAvz1MGhllUCSuQUtKpbYIbEvZNAYNkByMJ3GWqsCnoKN
trHibizEtFO/KiCs8oLjkwGw2xQ9k2f0qnv8ntwIf2rA3RdkOYVZX4VVrMdgMO92
kRO9q5motFY0wwEPu4OehWpsPI73Bst2+9Y6+NIrb8uJJeyF8A5/Hfzt50yNlSch
EJD8jHJJva2wreFwW1o3o4V5HDrMYNQDvuv29kC07uORz1gsugPgIAKMUD2KXnc1
D5VSLRrVqm1dnx8GzbP7uA6UzzCAiUY8FO8kB6Os2UkOJgfY5puFqLoCngB/PNaI
f99uZbi3Hv7EpT+ZDiceuqA98B7SqcLCNRUNaYngpJi6pJlRN1MoVbdxFuHqJBnI
3xcYKTfUU8/DxvcwV+G3q+Vd5hFAKtRb/8r4+c6o1rkx6Z6vaMllmy6oA2Cx93Ot
DTepOZl5CrxxV1SR6HsTtafeU8r67zh9D8hjt/VDTBr7eWK72gxF+hveMleX2hbD
Zd9gX3dfw7ANL08lRYmHA1nnRL+Aja74+MAPNNqz9pbzhMI3P9JcsJjt82APNhmr
HiXOQVS+67JD7Vl1h8xhA1lyn3gsb6nfs64b+ZpbOGjLyqo5n9+zNMIqduAr2d4x
e7+UM7xopSN4chak+tQhmXCgXAOWfiR14JimSST9yDq7pmJoX63sQIjMp+BIeB2E
q5x73pohFo/x+nH5L9KZ9PsQ9JU9wGOXfAUPGR0hlI1aCyz6SC7JSK9KnWWj4UsC
+TXsY/Rq0OKuzgYwt97cCtJ9UqNvrSpUAcZwY6mJhfyjQwgepsD4MFp2TeZpj7ES
NdW8UX28keXJ69LoIr+TH2+uQBHBL8wtb9ybPqSbnJK7rMoxb/0N0vnkmKCEE6uc
xwbSHBx8oZPYn4KKErZyNaxHLYSJ6QJ85/d3w7bYqwz8nqxIrC7GPH18xQLwoSYH
ItVriAM5lkE2Hyl9uInO242Ldh26ZJnmbI1ijsJl0PQPec1spm7IZhGqL9Ame+38
G/wRWkNaqqxry20c4PO3wBGr395hUPMTtbvPAjBYBUo9aH6BF96wiDfx9A2O/G/B
d4fXbFSkwWtm0NC4H5Nag8Zs9st3n4TJkxLM6WqJkXY+aaT36p29X12QygF6pK6f
Sx5c9kSaDXQyrPF1vlZLdd4dUaaSc7qUpJ3JBbN1nSlfB5FtbsM+vCpvxY5Oeu95
Qsh+aEnhkXd0BIMReiUDLYva2ls57qlXDi19z4zYULmmmiEHWoi3SvjPg6Qic6P8
iyWoSrfGd1Tl04q8Oq+rxoFtkIVaVeHGhP9bY0L4dCHDg5YW88NKsxpbhLpHWoqF
CSe6Io6zgnh8OknUNwD/pJfWnnhMav0Gjmwjzi7tiItkJiR8oQOqxz4g6rjc3UxO
iNjzQ7+IFb0pRyOLYfXiZQ6w0eJ/o3q8c65yFemqtcv6KcYWXYdagWrcOHbYLCov
FzpjpkhC2TAOY7oY6O+CmlXNwHjQC6LxYDUNH81uO0BBGcEmkQoS2B4T4I1KbXVi
UE49x1fF9kbJ7kVBxsj8f5hpIgMWewlZ77Dyb1mcG+Y+k8TLagveCIrHCcRDP00Z
Cba92BalGMVt1BfjtAyhxg+JfUam2ZuYbZcrs2nUfIasYp8CqcAom3tdIXVvxuYS
RHHGX9cyTYWLwS04Hx6yaMXfGm2RE96C6g8UcubcI/mp5nuZIKz06hoymZxbCWeN
E7uCw2Sg7A7+bDBhpWn8kfwJy1C9OQXa92FoVpRfUC+pkWaDqbf+VJCVw/E1wt5P
OSe83yE7E6l2xinIedGl45jWXiJUF/xE4EdGMQrXfi3QOybdCZGkteHFRTPy0ShP
mjQFys9dCYSOQLXzErJy88R3TeYjIiq7/t/eHNUp89NFVjFf5Im06Em26tHNzTR6
SM9BnZwI2NLz3VG9E/YrAFP4XytIPb8bIJlwh/Ou2aPaAGkozyqUcn45Dov54Q6i
7Hb39oLJQtKZL7qLuZrhSc3SbQ+b9FOsB4KydiTlDWafHCoaiKO3cyYKBiLMI0Qm
oW9CiwVIrIfyS/cTKM3cPn5FfFpCstpqCSwg9fs1Lz8Qh7NkQtr9EtPfvQftURe7
013wPFqUrnSr04FG4KhvVGFm7d0R+Z9L26c5W4JVWtCA42+kg4QOM/IQWT6660Gt
CMw7xZYIxe1PlUFDtCG669oooFB0hM3LoJg7mxBAv0N0r5MGitV4j3v01MUiLljA
xZvAE5ZY8sqra+nFc1VAFIPtW+A8IvE66hfD0hF35y8XC50GoARTqU/8TXG28+sj
k7Rdth+uSc/FTeU0oUd1iu24mhbrQkFpilPsE667s9DAK2Gbfm6t51A1oHOMxJ29
sywYto1d0iFhXJk+2la5x/J5xPOfs1PJHZHPAt/IizCfqTAzC55+weKX1V5k3tXe
GYvhYN2TLmFS1ax5iZ0P59rxKvgWredEy0o9rh4ww4SvcbUJhoGjDJvweOvsgjl6
j91DTWA4wpxheDjDw6iREbOfpxB6bGt3XPj9H5AY2N7px45CgX0P/SP5FDt+i/uR
k87K+he5xB7N6F3XfRdyEMfXNm+w2sztkf3tzzFPo+nre2vOK7vaiGWly+c9Fk18
LRskrDFWPeYgwv9PRPEILCbE0aMFgk8o3qqaWglr3/DxMM1NUosgNN3/IoSS74jr
cnaBzkNZ3k2LjfTdr3S4UxhYXjuwu6+RsZ9xwIY0KIKEQ3B7Iob01zXDL16CcsOp
g6UhecmUET3k4BNdW678Ehcm0JGXnyCJGk8/cbhf3DW17OK/kgsRQutmjKsvQsFN
YbeZ3lRSZo6D/GLHfjuqRB0IhSGs3pkdUqz0rf2/UlyQi1AajdLDQhJ9QgojPPFP
oa5lt6mVQv8KSKPQUGJYQOvIIUgo1sDdBkYgelj74lClZzbD0QiHSQ3FBRqIEOCs
BDemkPr4lqKHAmNWWheOJFGQv+qFcvk5lUNTouaOM3/jIZgg/tIkvIhfhP4tTj9r
ki93OwkFmZAlFNcVsPHlQYWHRuuZ4LJEmoHBjDpo8nlzu3Ogjbhw7n9esNbufFxO
wtnCfvGXMyVbsXIfl/uIyJQ1gKyPGX9rN0LPjMcyyOeLSNR4ZhguRNJ4ywDW7IHw
mLTO+MWYo+z6QgFbdQdLOWZ9lnisAkcsO/l9ft/l28JSK25iTjhgNty1n0b53ktj
m+S0HMtVy6Rwgpe71GPx4qXrMOApiBeUPIDdagIaC2U/nQbMK7lwbGcycMYHTBzJ
tlt4Trb+3wLcpyTdGdtE5VV58gmkW5H958nboi3f7kEVtwl45/BZL2rMBiGK3APf
tNTyygFGI61cRucaJkXCDNRNhJQpQy3ySIFlN9MXsCMfgcPk0MII8i/WjE9p3ApE
+nB+LunpnUlSA9PNV9dt3X3PhoVKDFdwpMQqPUoB1JuBN9eLlFUmWdmZH+5TMedn
KAiMHhI7A72DJj+Xu2y2D0gzyFjxslY2sImswKK5edX9ANq9+UiyHo6aBEoSwbFf
accqH+U3IN8GPFSEBVyaQNIwIThb6nrNs/fHScoM0altLKV0SddsdzFU3hvyl6ho
hG+3p+rzHTnBkf8CGkNUoEdfhA1/XbLCoXN/WGrvGfldINDK8C2NiG2BY3JlH3gU
nhg5419JXJ3cdc99WPcPQt/VeLPqqEdjfopLcc4KwADI9+qjpa2IETTFXADeBud2
BJyAjMERdpxA06Q6pKc+9YFJfdt97ewl5CsmWy7gfpsvCCYyLzKOOqedm12Ow3H+
fl6C4qsgx8mpAxWEctdXBAX85MBz+sa9dKaHx4YFavlscepGIEeRLmvyTcCwDHmQ
p+4JN3kXjlklS5oQ5aAjtXSy05EEzaGG+gPakEcQt1Tc11+NatjywjoUrUOV0/N9
6sjhqIiyVvX9aZFXzOZkOhfHV8dkiFi2DVdYyWemaBQJ6tH9z3KEERC7zhdIytOK
WtDPzeVWF8xCC+T5uRvKCHguid2IMbQL1O+JdSNU45cfxRLV54B5umYwu2nTdGzD
r/dgxqAaEPvGOmvjelWC8sXYKD+X1BiCXv5t4WV8OeqJLhlVgN89Ao4q1nu2ZfUa
vKIvPdIbJCyY7KcvKw6FXjRMIWtc4OY6QcTWG8Y9MBI8+OBrTZ0lcfNcyhtOLVnj
732DeqO87YN6ZfHX+6fqS+bgKTf4d9A3q8kF9BCq1d5+yoW9ukc4Jm+AFo/dTnea
YkajJWlmG9AgvNtdxu+IZUFzxAIXYs0yy2WYeIBvhnZDtjq0Ch6QJ4QOBFVezfC9
j402ArTBvy6tyHtN+02N9Ht7Zxv+RpaxpdEcg0QvsDFSY9c/n6V3rNWn6nowi+gh
3bBrOzz7yy/3IOUzfSt/Hk2bCrzNpL3altpW8HWpSjZBKttKL2ac1ltTw+aYAQGx
41szJfQN3Qu+oXkR0UYHAPJHRZvXdUAtJnpn+aVB8QPsNZEM+9FR1BEKP12WfbGZ
9LDNC/+8iU5Jvs97El2wlxk2NM4wdDyMu7Sdt8P/FcXKziQK00nVyfcfaOov5djS
ZjRPzlKrzmO+JURkEhqWKf+/81PgmG3BhSLNVzK8EHkIlsc97yLZ5ceYgZBW1uij
9IA/twmJpD9JIK2uZtjLg3SocTL/nLWMOQ5FdYsx1AJYfhpNArnsGFyOSUO3wwge
1bix0Z7JvDGdXpqm0h0Clap/i3WaciAXk7y/71Iii4folxNebRf+NKoNUBbCLKxc
IsJAkuERopdPvzJiZqsW+xD9HaPumZFMCqJV2wvve/AqOSUFEIMG2U4pd2hg05OH
jUGSRbdLxnS9vFNU2EIQToR2g+PMHXGstVKbuKJA2D8PG88Rv37DElI8x5SNgtCW
XUl+9ZK/UcugqZelHMSro93nHu9sHDYxMbmDUIoPpvvpBIwXck7E1UlGe4zqyJ6w
CnvC5Z1Ew1pa9yyKSoK60NAy5H+ZxsU5PmURrdeCmyxgMZEzfoYb4X5vGTjRQFEg
DwiswQb+srhS+L4lX7c3gZyXsevPBkyUVTjnVudmzKp/8UOqh7UMuf018OPQQSqo
WBlj/V9MWlvw9mgOO/yqmHLOFeOIZ8C5k3uVl94XXxLPKdKHEe6dvkm+R2FVm4Qn
UV83qkGk+dMtYj9teRApz5p3XEHEgs4VX3XXvtHI2I6PTeKM/JtShPNg4dEmSDJV
LCovOke8c4/kJOAQX6Cd5g3ODIjCTh0JRkdnQQVAXvt/Ivi2o9Jtc7s58zDhac9q
SdIMLUrlr6LavOtE2bXrSAFL7Za03+wi0x4ANeCmjriZBhmbJQEWDQ+4yf9G2Bfg
ZSP45mSIGMOBK7IVIZGsPpJierZoPbacxHxPoI/15ru8ScgQzdRIeSWnc3tQb3FR
tk5uNAfkHCohuIzrc3ILKU4vrj2T+mUqPsg7VETXOBAWQaCmKgKmhFnJEEo9K+JW
rl4gwN9OJZ+ieHZFJe9tn60PqLYG6Dw7Ek33z0OW+GUtNwkYQqMkCCukT22b7HAP
Bqumr20YZOQcSSmbZKulMSzHr1cGaTpESjyYCvxJDrnMKd4asllibXD7JcZITuSN
g/ytNN8wK1xvegQMQEJVphDiZlncqh8MtGeNQWmY8pDxtcyM4ZVmcGATOkyDf/6L
S0RDEk6WfSFWduXMjMKZ6xcGMo/GxeFKa/C+vxnR3LvHNd/xR6JnQSSedIVTqHQn
8dFAeeuvetuWIA2gBZYorxYwOmxK3h6oBP+9s0daanzJfULNA7K4oh6BsboTg0gJ
4Imb5P6FwzVUA6e2ECrOigV6ODmpZo7yPW3VMdCHZkLU4LjdSsf471eR8KcIZloY
br/K+9g51HIpWJ9aN8gT/0ZP4tvySgK/AKceiLSaWqv/7etuPwrQ8eLqc0Wpe6sq
9gJBngExqBNdK1z4+mxoLhomOEAQkcsOdgB51rqy+Q4MK+czv7shbVzLqyW5UGO2
a+cbLRIIJwKGgSEQUIMtBBMKUODzaKihhO5YFy0UgqW8+hV2+2Xp73jpLTYYOf24
QpxUqCagy8Ijeau67HFxC+hSgOgssCH+hNgQZ0+LCoM18AdWbtFV4wwlj6edoq69
vf82OfPvDxnsAUlDhju+4KR3dllErCyzMqjod4NqPOZDjuTd53D03BoNWcr9WyjR
ShTnf5fm7G4RQViY6bxBz5rRRxKdw+OmpRN0UoV0HJJC//+itc9Z0i78p9zf34pR
jG004GXCev+7Mzj0hf9gVLLiHci27VUoMua4gxXALAeXsYo+wkdhSUoT2WsTsibl
hb0nm2Mm8QKD3UUYTP6r/HEmDF5+ijttzarLlgD5aUOIBJBLBUlqsxnPDYlFDFUi
7Q2Z83rJUZRdIUT8a7t6K/AkiZgQpwGRyB1ayUay3bC0QAB4QeZrR6WtmXzLe1c1
zsqwiLqlL+zLzxYqJo+x7Yv5XHkpDRxVq3pXhDYx5C29h3OyOT1a7iVDSJ4lKhGT
Tn1APbsFHQhsIgXyR6BC2yZS2jvxzvxVp9NQNPvMbUnJvNkk8WxodABGQjZOjs6o
G2pynl9qhL/pj2ibzGMzwzyp723eSBfMLKliu/OaSUelUMHyU6gLUccnm6eSNnTu
AmzBuU9OBbN/UrciZ0HuzzbTWeQyXXCsVBvpgB3v2PY/JNpzXx5aTq0VyKDGQZcS
QuhB3QP2f9Pvn9Gj5cqRfa8eePy64wPj/PYwG3X4ARBTNFepxoLM30v0kjMDk87S
CnsD/i4QGbdHTJaJM5Dzk9WIW0RcY1sis6w6j0kG6oouNPAPrl0Vfo4FlhNK2Jea
ciOsPCz4FyerUyPFnrPTMDnizbWEKT12o57mZDtbtUeZtJ3ccRjOC1D9zV10/7ff
o9OIQp5n6yeJ3kF2fajDpSnVzw7OWMc38plt8Ms26DK5BvXEwlX2HrePPLE+zL68
kBT7cq33xDsW2/yK37ilOMsyLrkLEtKsIeQaiAxWT06AR99Dp7kywh+pZN/5tY9Y
WUS8kDu951wkY4qP5bYGOpFGSFYYP4AbBks7jY3W9G8u0ixzka6Mruw0HMsMcMfK
p7/nVAkzVCrSUIRP+ZTteFj3c+mm5fpzchXTI6ujEgCkJpGs/gkSvEJNoZVnC+UG
4dSnNkGJ6YbQJUuX3wSp+j0ajHjGggolFYYxxxidMFt9lKJy+itz26CwgOuqwcHl
Di3Y5tPzakgO/Q3+L0FJ0G7mJ0iJEd9UYqIdZoy6a+d1TLktnTJ0AHBnDvsW1m77
EI68i66R9qq0K5xZyohlOh+5nJhgFOVCtyZaGvMTIEgzyAblySmHvQnGab0Oq++1
l4OSvMRKkp8lVJBjpi2GQhlFIe2SIoRgQOwfLxGDCxl2R/bH8glOp1+eprhZEHzP
8jgYwKEcjy7uQPe3O+EoX71yk7VaMChZpHpWmUnJEYY4Al//3f++ErvjRQ6r8gI1
Z24/jqK4XLKcluWR/4TB7mUg713YgzjWHMp/4KtBzXt2DtpcJexTlYf8rgBLf42Y
zrhYHTrt8IokgB12sVX5EF4sandPl0mSMHxLY9abjJr4493q/MQ5fdVvmwUhFGBl
9H/cDGZMgLzcL3mSBKXJqi8LMx2p6t5bqoVgppcbV7fwBFpQwBEQtZRECNjHCv83
8A8lTv9cUhJTRiAHSOIAs7E+nKE2VLPVjDzJ3eGJuZ7jUWrTo+TsyB/EEnWGYZ8x
HeiPXmJLgfHExPpDIhtZgDRBl17QHecD4hozthf3yLGfTSImO6UfQzVI/d3y7vlW
ILSspWrlCRya2MjFfjk66MgI8SUU+ZNDbKkOVZzuRd4XOj7FMOFyX/lTe/ZxtuZ8
DqPdvJ8FAIClZ0B9ldM76Qa8eD9Dsbri4Hv8Yy35y7eO60OIN2Y2ct8bLNmcII2c
MAlcBFN9jscHNwfikPCc4z0Zx330+pRh3qB5cWMyd6N0UNSPLRdxCqq32jRnXkRx
GZ4t7vkhaIcJmgb+mLuCeioDgCU3e/FmHWZYQoyIi7gqDaEpgfdpjLb8feF3uclV
cVewlgqIr324D3tjGapIHehjC/ciG4lyUcEOBfIJ08vu6yWTCtjw/lU/efnvBf1h
I3NF/5cf5ocncibigBhNsLQSPqO8MteZ4+XshcaVq0OZb/JAcLKSts3NpZ9Dd/oR
WfpDyB5b3rV/tjNV41MvgN+TWxztQBHfb18/HEbZgc0hKokO8YXCTxHiyBKAk1VH
7HJzJJ2CB12+mQbxCOCg+fMiqghNPHHyhw+kpVkwInStq14bVZWkgqL8p2j5GAa/
MGJbBO6Uw9sMhypq5FpxlSQetFIZe7lp9A4CD9EzB8LHsZZwC/qwIB6Wb+0ScnNX
iKhyz9eFs9g9RzT7d96whj08T2yqrWErI++LZkENOmXusSsdnWIUfcktqeqw8eCC
yECNBtW9kdGOGAdSbGIQg6nlQ+4N8+iWaIrkteW7HzS/Oi0VKz630w05s5gsoH0O
tvm3lYoj2Yu3E9x0VjpeGXhNclthlVbAqYx08ZzSHctgAKl3C+FGkwmPCnPu28Vm
oo7FKFgQ46IQzibZyPF7IqqqkQ3W5rBOXwE4xUCMA7qApf0KdLBvqLtIq1/NUI+p
PDq45aJrSTOF8SyTqRSygHUesk7hyzdgKbPMxSIjWSqjlezUkdFELHSQtSUXD8mV
gTkYdi20kcYMlmKcw45avY8pajFewFWLkXSwD+n4DTOFsb+jSj/PPQ1Sv3PAfT1N
Oh3JC4zqVRMRbR7SidMaPXcK36V/xm6goaOwHJ3rKHmtMkCaFEhFvhWx0rIC3ORP
zq3iby91MONExXS6FAY+e1YG9c5x8KUOx/W+gDudsdRHiMqEXgFmdYN0HO1LB3p5
wze/hp/Zx/GVElOJ+LehCUE56oN0qjJeV3TX6+l3OVPzN4Nrzg5Lq30aM9dfoe9o
ZQnc/grHEG407hBbMcDI7Glp90t7YDHgDplFG6JAhvk8FGbieVchOpfurSDXEqT0
CW/13/wv4X3yM0OLcgIWaXB+OAoFOYbMGQmVnxMJ6fDbhSPirLGqNbf0P2gKpcBd
lwZDK3E7ozq9HlTS47t7EfrOrGWa5D4jMaa1Z0bFUiOTL6Qd97E3cmAkrbBcjT7f
OOVzTmOF7KMXr4MaOQYU5eWD49KjGyxAB5lbVijo9Atd5/VdR9WKec46eyH+UQW1
n1tPRyDxSkImMJAugE/88gPH101Fc9iSh5oKfDXIgKxgNt4yRMepucChM4VSVSyT
vaL+3+JIFVUsjb+FLs0FLd/XZfErzL0JO6gKwdRmA0487Dng9DHhl+vPdmPv7FnN
xUwpFCrtRXdOozc3DhusH3L8LpswHWRvPWq0sDuveCZWswMlbQb5DgLrj5S1Kj4i
ybe6ppc6P9j09hWL49OgABl0tSO5vQMbTBV02KQzUsg7ixYh3zVpRPBHXazjnbaM
+cjvNHXLK1KpYk7HuZ9+YnMKwygjaP7tNPUYu3TCO/y4l6Owqgu4oV99Yc+IOif+
tJGZqjkMYu/qOWIvxeFfmXAn22aR0EPiM76u5aNF6YJhcIfUnpZVzlSmx014PISh
W2FR7h/Nf3831JegI0pltnQjVrRz4h2oJ+WuP/edVg9Dl9OQCjl+KcIM86LzWC6I
VxaZyu/NqdIcuGOIBlmXdHQxAHCPXQuNjyHSAJ4fP0ifWmfC5FirCXQ9et04Kq/C
BvcHDC/VMLVXIpQ4vZDPGXF/YsJn/hIH1MBgNXhGiMtSDfFExhyttOenMrZEKXJ6
4SWD0kMfXVUbWisQBSsJvfJSr/k3PbIJE5UfH8o3x6s4rfwzNDeJC8xHCgWcWlbp
CWkKCAVlNjHXVhnKhUd0qbSkZSdp7mDhiQHZ4gEmYlW6L/qjXX/3LCrqjQEnGVyk
vMOc/UGEXWXBnqjjtiRsTC7hsqIb31sHc6irK/lsxrtR9afCsDoDNoZOlVOJ1ypr
DCNggsxJI89VNOi6V7fs1l8hPN7pOW9p9jBWXmYS0AULAIjxtss3Qi0odp3C/8BP
IqlJwN82CVoSyqON9ZknCLTIVTxIQxHpMhvzZmMGurb+wQHpEAoEqJqTSBTZ0oOu
bwm8vM20xDz5KO96NkjhSues6LQ3a3ORogQhWCID2t5Yu4mCjtTHh29xS7OBEZR9
aasLzM032Y2BWFd1IbC6NzqveZHBj3FukB7UX66VhLymfm1HLTbJENBuVxetT1oB
uioE/P4p1rXizCHU4Dq5gOnHlvFFJuek66bIz4CJW9iSMT904SrgFOcnq+DSkE0V
eHgAlqVIBcaDMEWK7ODvLdAV7ujFJz0Nd+I0dz9V03tBPPv3UA//jvAUWjx9Ih7c
QJAHdiM2pbG++VlZCvn9O7DuVYZcGxCRk7yqvChAtx5NusoVW07oCUjKgEFRD6c6
kPhIsggn/mQhIDz7eU2zy1h3btW11/VW9zS+qimSB0/NpQw29B+3TPoLUXAw7GQO
tl/kQdhLEf8ApmTksQxFzcaSThnOZaUnSkLColMMZtMTAPI8tMdQLf0bfqvwX8BQ
vscbQY/sHa+3sbmsjEsGEVOZsWzwUXeJjpbn+ot+5YinghcujDCbFBQIqSnSAt8z
5TYLc4VXuPuUu59mGPNf1tSmRrPdEFtLXDApVxZXklZ27kaYI2sm8vk7nc2brL6D
5ulNlH0WZ6+U0cBoiiKyZ0t7yV0XganjhdoV6EzOuLZyhefEOIUC2iMLthJBNoTR
QTyF0OnrQx9ynJ+IM+4s1wWlBsHO+z3U1eKWbcSyUxeXMf6w9lKOMjdguHRh61cZ
uOe+0P2DXuTonDpGwn44JTof8jwrMltVccmE2N1dckieWNlyJAeTCi6hiyUGvY/b
2J3lERF8MKzt4zmJ9KrzO/y/lC3vYZsWmqdMBGKVNzgfhOQgOeDHmpKIKvePY7Sd
7Qjhv5CM0kCHuInH83bsQNl9EfGQrcsLmmabPfEShYIiYx0CWUYz425ctqzovD4R
E5/+nSOAFD/jRYVkOsucMhSVWRlNolkM9nFwiEF+wLXIrChtIMSI8m3EF47Eq0Tg
4t9n9a7tmb5IesjdxgMGmKoaxqjOgsjAnEA7XsFz0LK7kZOYc58suTDId0GwyA0v
MzfUw4CAspheyTC1Jr32qXmbQVruNDWbO/VAL3/KPpe5TiywxOAaiVQv+YEa352n
7tDuD7QJUEfJwm6d9W7RVJSdhPF2HGvotjmG9BFEM06jyEx4krKUWvSBUhOsTti3
Z6mUu/BTR5mRmT/NcTgsAhbXfmOMItjIrx99KuwH876+bGMTS77bI9dMFn7e9Sqj
F3/nWKEQbEBw2dgnk94NF3Pxn7oVGY4NYMIlhI3uGR0j7TsRriIol11rVj6suNhz
BR4z5i9GKrd4x81HJ1+OxNQJWQQkztiGcDx8joa9/cSMieRvO1RBL4BsNVZouiNs
TI0rWarjxj5hSPpQfZEowvV2B7aXyT9UE4BoXu2BRqRqDX1OGq3DsVQwK9hgcso2
L3facDp/mRcY8NBnS0VpKnDIckqP566k6INb4LpX+EVb7+DNEv1M0Oj2GQghsxzN
SAfa7kXTGhYnDwqXlcoSbGIbQE7QcmN/vqytwB442yGD70da+7/ey6rlEmFzUejB
B9eGIy4j4RI51TCgniSjDmvR6dgqDtkjvl/kV7YDgggUEMWPjqX0WfXxL8HOAJFM
y6yeq1iMffslWuWiLje+WwRznqFPhfL1MeXrsCDpUlkERGwDp325APg3EXcPcSBQ
IJPjGP1z1yR+dvlgqAAbeKi3xJhcF2Jhbrv+gvYrYfvrnMYf/j10wccz7oufeoQU
BQCs5XEiFJ/ZhsCoSEFMWChw/eldAfEbS3DZXt1kp3pG9x/qE1KPSHxgVRm1pOfl
YYLtQ+XRQ6TbN3lb2Ur3Uq+PhITo+HFv0VWFyHGIrnLprtk98ZXnksP1HT45Iy/q
fjc69bvnvms6aJAJ8x+H5poaGCuIa1puv7HKov+LjDBg9oYhIBjZYYzH5uFh3EA/
RMAcdlULncI5Vcuq8wqhIPllvoPTd8gItAkeTYdnR76jdJDTCFSmWFWh4OvYcYLT
W1G/ufAynlEJ9h33NYB4AkMK8ckXjWurh9RL048x7QPQYmvZQRLN/Ju3IAfScXHx
6Qfp/HZZezzHYKOI2xzXmyZkscV7buwXwtB/vJcv5HqzgRK7ZQHiAedJJu5cOZ/m
WAVvjpHNfrb+zZUW0eGZpeflUgERE+NgxXSjkBP+E5lb4z1n7C/5UHLknB9A28qK
kBE4UAuMbPO9pQmtsDFIDov7m8Mz5uHwX6LDz1yBTn/pE0xF/gWyhCWLmDUlJYOc
Ho5LvCh1wlEaRZI1R3w/nm21q4s34t4y1Z4mOmkFaKxrpXxI3tj549PED0zM0wG7
heK+TqqXZU4PKzz1YWMvtRsE0P8krqPBw1QE11BKkk+0FONzte1OalyQ5oJjf3lQ
gd0fCm+XfaVq/7psaGbJCme6mnhsOwIhB5CUwJsLviOPtjs/xsjhoek+MtDfbf2z
F4RkTX6YealDkE/MgaabHxONjTEyygd7DQVEeN4Z3rXzgHlyraLT9YrYGiO5KZt8
kpIRIsAYipVJ/3lk4wxHH1C8EY68BOjyRiYKSmAPNty3jv34TuEm4+dRPSQGlTAX
8gLL7KO+m91z3ncPRB4PDPEhph8gOWeSM+jT45nlqfZ89K4r8E2LCEY2PtCGZHeu
uPBXyK7hl9hA68sokBCX9DLcNFSG8OzgxJS1vrgt4EV2KjN+B3xOrkD0ZZ/aRpRx
UTpynwOgZgds/Q98v+YsOvnfhQT4JpqQ97hC26wDDzqATE9oXm8XEbp44lONtDPn
BMgVctpAij9WibXAdWqxesePw/17tpvCcjiaWXg+oDcTNoJe4fupkAMadH1MFOoZ
Mqd7VFiP22bNrC6t/EALMPSgi3kOJvo0NMRHxe1w+OglrnJC7jwf1zgi3pjiWmpz
QVbhpkUKireeGS19k9NB+EcOFZpqu/TRLY7I6VgR42kprRRdZt3r9PGnAAKBcj4T
nw+EDns18pK+PH7k2A8qKEAThwzaC5Gq8dcV8Blja0A67oEPfnhU4/y4LxJnLXBs
kXErYmggGEsx2iHilqcDi9xNGWOlGCSNNhzP4GOHiOZicAiUdjZyZQ9GrLSWaBBs
5nGDaPRIS2DbVKWJtMcWBWSjcX+HunB6YRpAWzTKaDAD/5qiljixF8fS2QJaZ0tL
7blOfIhMXIKkIveEu6ACZjwnNDZGz9VukJHC3bvVVwtb1NZbYNOyfFDQKgcq6Ur5
m1EXDgbjJ6fFsqMNHjXs6nqSnbthrHO3jRTr/QveN32f9E1uNHu3UU21PFOy9GVr
cpH2VTAKOcesdij0x+UnAIyvgGx5Z+jpFvHkNvjZbx3ew4irXtQGAXglCBXyOBNl
MPQthAyU0a2wmLjzeh3Hl756dzdrLoVfEbkg+GBW7WFzqZrf1azw9zMDrglCbj8X
V2ST/XBwKbRharVuawueZyV+HCQzfHVQfXFQtKKZ0QfcRnvDjyU9x81C1QK0GHx5
YXRAzaOqCG64uPMVsqhvsRU0yaA5KDnkOR1vKAxkxqv9Huwofrjy+9Szk2mgz9JO
VB6fqzng56QF5ICBkozIHik7Do9h7dcYgspRg8QET68ulUgUP4VtJJLgOY9j0EYc
liZ6VytIdVJiUav+mxe6zTFGjaMSU8Rufw1M0MsqpFWc1893Rl5dRnuwcQRNfl0Z
e9t52AqxAN6fj6NWqSRvpht+ibFiDbmhXKs5wWOrrzXMbJoTIMe+xFfLsSB48nuS
IuhtO8Z7wj4T3FrtPrVQjfmPDluQcLX52qEjCcyiBrHW1gTvPX7sK6Pfv1AdAbpU
bU2Paiq9RPkCYoPuzX2mXJxu3AAw9yJblhYXN/veHvDcc4Q8Wh0HoCWJUeVFAMnt
BxbFVVgbViTQ17c84BoSI4Nhz/dH7tQfYKjyjoVSq+cBQvxuJgmOYyfmAmyjGt90
xLHiH8bry/oZEBTBUIDOgID4Y06dhkb15ZnAnHmhC6TO3fnxM4iRPXt3kSymDDu3
/YCvPJCuV41gDPk7WE+iyo99Q8qH0SeVqWc4gWCEqOn97lbXct+GWWZ4yW2xw7WW
tQuyRQzc1FGEWC0CjjOx79dTxVgPHHyMsZGH5QWUPobWjmUf/y/mh0bW2SmhQZz9
xxWAjnYJ79D0LvsslwUiDWWEnAQvnZUdr6Bg4b/37HZBTnsMPKkykyZ3PnKn53zW
hX5VrZfTs0EngPOMx4dJl4X322aj6MVJLtz9ChnvXRuaLL9ZyYTXweG3e+YY/hT1
BP/TN91nXozXdNyTuY9c3rUehmV8BsPy7Fz7A1/Q6RMalMViNLlMWP3uEvsnF4nN
wgeqCZcFoVuy2BhvKTLdptMVQ7moOzP4jyPYr1nc3yySS02KBQiJkgkXRuBeEVk6
PtScAyJDCIDnPIHd6Ki5KdwFWh+qc7VA5fWkiFCfOnGgM5ZkY/3DkZ05TB5QHeAR
HyVPvAGFGdOZFe/Y0XRBLcZyng4ZHjuZzR1bN4e9s0i2+ZrbX0xJ5iIGCn4xaoa2
niUZVv/ebBG61lF1R7C2pVQUmBBpJ07PRQs5EEmPC+k9ESh1GQTwHq36e550K6Jn
oCnflPJgpp0lrq0v8146P5lpMqqdpdr799W0g2rMlpqgf75h1oH+57u5e/7VmGOV
h86cIA2rNUyZT/7PW1/GIXs4wXO+lWY8SgXMYG2cNYipjy4h725A88hX+pKYGqYi
NF2KPCE733m7padoIwXU+LzDlCyHuWBEHei8M3+rPh8lSgsH8YcP99EpZuyjxMdY
e8seUGbNE+wj6T09SJdAmjJy4wQfv2980PkzeXt5pa8nSPRkRKEtAqjSRkxOpGNe
lMNyrM1FCZ8yAJyBS1aAzCDc6345clxVULYoQ2ArbMuSaF11ChG2rBmD0VpDo6DO
f1vMqCQ19fQnrqEM2ggyzOxjmf7ONwDsY/9nUMdM5ZDszsG7u8m+oyx/D8mkwpyi
B8DlqRJY6rMJfIsgbeBFdza50PIVoWVuf2PuJ253+H5m7RDQG/JJS6h63zy0itTE
P/8xueuoxStV8cbf+WJBbM9N38soAp2+rkP8fcKe/vhngvICOLUYgJrFgvm262eC
vYLomuJ5QtYN0UIQvu7Fd0m5/e4tNCk6M1pS2AsZh7WyYbXSAwRW+2RMu4XPVf6U
SjD+vHCXGNwjtWzXZ1OqGaQD3IZiG6av3NG/pJ5uJ6r5T1ZwhEbWSjvR9iB//98/
wGXDeJRpsrST6WStveU9+6pt1oGe7uITqabr20lCyCEIZRL97Iyi8f11QCfYvSwK
h+PviiLA3xsWlcCudZyXJga9LE/CAR9NMBrt1yZJuf6FFWGxRuoyl3I6UszWnLvc
JcnNJaivXtYJIiXuhuTnNBm4p4+actXJE2o8mY+mUnqF6O9b6y1QQ9QRRftfLNg0
o9ZoKS79QQ1f8R1J+rFAnU4a7wISMSjMPtmLc2MxtN00+0ucsAhh340zePw5fIH7
Yzq2iP0opN80TgGsDrx8N6xCF/GP71PXEUjO05vfh9VonAKNKieS/VJdBl1E+tDz
xrTcwbhBdjL1+JjkegKip7ikuwr8PkWKDnycKinREs/RGVRmzKVli8JKOm2PYVaU
L/e+/SEft5j6YgM1WFpw56HSaQj4vAV8CYI/Q8jJnrNDTVBbCLdAW5NgPIQhq2ds
BRvKI9r4yx/6taDqd6i/ln0fiaiyDA5OJaT46uJ176WwCGENh6Pto3UuKM6Vi2a+
/0a9LuvKlduSxYKDPHSqwU2b829401RgqAaFo7Lez4V6i2aliP3l+LEvry2YSXIt
vOo6xU2nEA69v2oVT8gVFDej+HumI8TBfYOrdLB9q6ZKgCyWUGc0RYMEryC/bsOR
LtNswDUFNj/dTBx6bIRPuSqhQrn9zV/K8sK84AfdeAs3ykfcLe4yiGXcmX7L26nb
GA2g3PqdgHwwRYLsG94GuHupPhQc92Bp6GcZ54kfS5wLXzIV2oTfD20Hilv2IQxa
bDRNbtpGMvfkOhmJCZHwh9ILkP9omHNG7R/wS30ROcH4B3Di+MB3vmuVAMMCwt/e
vrge2lcVmWuRxRZypiGdIYd8SpdjLCzVheodiS+kuMKJRL6Y7rrcJpYlfh3QLj5Q
hLDz2qB/gguoPdOPvdwuMUhLVHUg+i4VeLW4jFdZ9JS9EZzcKFOjb3BpXQz6jwuJ
EUk1o3FjfOudBscZZtdhSgx/3ucPWgQ+9jlM/xQKOXQyOHWkT/qxAWCR1+zsk9BM
NfKY5ALE+k3JYILmMEhnZuxzPCOMSdCm5mQdfz0z+hPW0Drvyt7weajljscRKLz/
MucA9NI4MTqVkXy5tVO4doFJ3elYEo2mfHPrJD4hqEOGi86k1BrTrXN+/YZry1VQ
p80d5QXhX5dRNwn1D9tyLZBQSr2IKE++R4oQ7agmjh44ca7rAYSW9fmvcg27rhpB
gmcbFvcu41CWqkg7eBUbj54oOEJrGjmLBSgJ8LTlP+3b7xqQgCe4lyOvjqj2KvKR
bzHNcaZlqyC62CbtUWZMmg2l2SQQiFbNEu+2HGd5exZbqBzyZpG/0R9A5qkEtwse
eShqxZ85clZAkFxuVYo95LzD+cRC0Z7V5wbxLlRC/3TyQuhfKopSjHqKUSAWlAXA
8P2fFubpPubvBdLtJuM6FZMUqFlLUPXmTd2JX11au26f74tzpbgyifk/eeRFZj7A
S9etX5qNuKedhlFOe5zH9zjTteiw8D8xMwlaVMNOcOIlG9+W5zz5hm22OGYhX+00
dE84VIGFiBexaat77fMFr3g/ThPWRSFVeEECqmYPZue/EMGPD9Wt2+So0zpVF8tv
gOeSSNYKuejircBYvFlC8sVV+IeZ9VFEaUjVnacxH5NCCUm6DFqHCbxA0RsWLxYI
N1qCigpu2qpWo3BVcew6ZJVZ1isyZ2jJSy+yiqp9592ho9JD2m/sZ4SAJidxzH/q
zspdRQpwIN/jpBHUbBgESyHg/FNdoJSmmqo+9W3LFOSsXdqPPj1JeOZd9QO4fB6d
E+liRmmyYfe/NuAKu0cWCTVzOARxT8SSz3nuBS+Sy2EomQL28pUa21bgvu6yXAZd
aQZ35BRYWsOLRPb7OIWA0Y1vx4wlgeA4UueCeK+ia6yjycEGfoZcKY0pqWnOnxNS
DAbP9fbe9IWykneWpqirKMn5H7ML6RC/vLVPvEoobxbVmfEc1PnpaR+SqZPeEr+0
+qds88ZTlEWSbZh6WNBd5Om6lhILfJEP/nHXbXvF4VokhkW/2a+7V9KZtNYMqN52
R5ga4rWXyzHwMYKqc+NumeyW6KiGz6O64+/4Gxi+J63KgueDr+lbEWqT9AH3qaCx
5kvFCo/KVT/WvSQFIEPhL6iheBjY973fz+T8MraVNW1AhLwRyh9NQbrxXpoK90aO
uJS+px/jcxPyD5lN4bKAfTmwEFb9HRH9NDHeAv6eqtxH71aRIhp9S8jXGOCaJ+TD
vNix5EM8qya+yTVMhzZRRZWS7mrptfnBU4ZNXFzq0oXd/QMDxrEA323gyEJYWfDl
GZ02FM7qTlHAcj1zmWVQsYcMU3vdHQe/pHlaZbCtgdm8Ixx9CD44CnBcI/wZK5Qo
SWKIKLbDEt1FxNkMHUEbfxlQ2LqdvRHIduPvSnFLlZpODvwSIWap5g8NJMhmda+C
nELEuaK0YhvtJrgKteHs7agPHpQkT7LRMHzdkRpBjCRMZ+m/SoOxYOPR86xqX8y1
kEGidqHi2Ts9DiwyntXM5KFJFCTi/LoadWSBs8jRaJoZfxnmpft0pi85/EI4uyeX
see/SdZXatcx+1J0jk0xn6p4kiuWpbFKNMmir+2pu7C9AZr95ECr3NnLOa6rt0d6
wBEdAZouvtdoKBnQHCI1RDkMeK/0RIk58xcKlAEX3wrCfE4g5ZUR3na9Cwab7AnD
ZVC2fxAmBRlqgQ0bYCP7wEeesIMvnCpOso91xDIxqwe16nkn3ZlFxufIpaF7notN
EkYd96tyhrxph7iG+6l3tdSGFNYiF0aCQv7zhrsQ7PgxE6MID+6s7N5UJ9MMj4Gl
yAGhZR0Pfl59EbqDEsY33M/JyZTodv1hwSfS74zXmdrx00ByaNQYM3iLbWLU6/kj
p2+CDZ/DFSYvdjQZPYywuOI8MIy87/Mh2UvKBwOVm/ntR17QkDx3ph8LE/Su0udT
fBGbLy5x4pEbyBhcVKylR2Vs2lsXz/kiD+agXhO9xX9GttKVa6XZIPoBfNEYrpYl
y9/QwaRVNrU1+p4yY0PBEY+L1NOikhLeJyjSc0nUwtgups+QiENWM5rx5/D1irtZ
nVLgFhXxV2Cu3V3QGtp3IU7F1Y/v8+9SqlUHA0pnHesww6h1zycdUXlEFDJQZUkr
Fyu5s/gLy5rMB2vEFTwkZC+yF6l4FDTuUuabG44OrSb8GQLUxSpBqMDKe5vs1uMQ
e8GOidmrSl0H/na+xFKjX81DhxJUYok9cn8rhmE2sUqYWKtJP9Yh0GnSoKvlMT2N
xjuEytyFGj6Hn8wY9r/MxocbM9eEuqUxJ1JjbClpBAcH3Ti6enPxy2ookj28jc+n
wAYaesu3Cswu8MmJwa1w0IJAbfhDESWNHwogJXnbFhcZzqEqHLJxUXp0rGWXwfEC
E42czKLGvx3FRFpsoAJDOXzINoIKZlzXWgPrPz4GN2LO39G34RugtoBDhxyF+tiX
xyQC8Wu/VVu0486Hl3r3RNVCLOv39VAtcoVsEuqSZYuW5TBctWeKLVW44Ns3JQlR
LW1DOJjbkLu7Imixjvbgsaw5AbgAP9YJe/pMEDeLRY0+O9lHgeH9F3GSl10aJO51
LI12gytNiBGfjJ4wcEpda9lTvCWZiRg6E49c/LKyDxwNvOBf7ogWNCHX8NAVLxx2
zMXAM6ww74HOJI2vsXYBYKv2MgfDKTEwCXN/5WqPe9R5fnCgXkuvdXohyLUs6QBX
BHe7JCBAoBRcFr4GUCwMSHr8l3X0lIXcDqN7sKBysvya440fsVxBzHy31oCCjaSt
+z+icFXDETCrxDYg1L4onoqDW6WIXwhhNH69JoLzRAlE8p62676wdxx9E4Smvt2X
OELNm5d8a9lD0lzMXHF/PL5X8K3aCMU3WsZYD+Bn0kqtazxrTfof+q7pAiPdOfab
GPEecObkxT/gvznjmcFCzDs8GCBPPvandizmyGlNUPBhNpvXqh+xmQrahFWjBrHj
gPMYpkRpHdjda0+WXILbSwOyW5Rxg2H2mmkV8qf1osuO2NyfT8B6eL9cNs1W3SQW
D3D/QGJJc1piokr3PDu8pB61jlh0sY1OjxOKNz+WoNtSttlD6+VlEllHXLYdkMQP
qblHAxTLjNNnnlQiTyYq8HUUkrn0jeXiIZzAeO2onlJ7GnsgzxwZPTr1TIlDlGNP
moC4/htweYk68/014p+J9b9Q42v6B9dTVxLtwk6Umc387N+h+A1AdFMzB7+oOVwo
lPkjL5rJjVtRVGNJA4wmE27FyctfT49E+7gmNmuNafsyGPV6RAxFx9LMAz8xCrT8
eM6cXOPQr/nooLaW+xB2osrzCxbowx3BvgXBMzQW0hxTHEb271JCmAxvuZzyq3P+
5v/0lKlmXk9fq4XBdyEjthcuwOCLF7vAG7GKoE4zF4JmbuYo19/EhXczfbpCUdQx
JiUc8VoM2F/M3/nBHMms3pRvG/xYO2IG0AEdlzu1ePjXAbcCYZTo5H0gahu416Bg
a0X4ZNpIzX8Al7q+BbhkfhmtSYSh2kAYALPAOqxCFUXsYCd1wfGt/OKC7mVaMz/r
DrL8ukJ1N6DOyH2lVtwiiQUazhxIYRlBN93Y6n9Lc5Q9Y4G+AMQ6R93dBUHwc9hg
LqdwLlUGBGA/CljxF1CSk3YNzaqrVfuxNWkC3hEF5wX7pDOV9P+TbIGvtkN6tgYL
f56rSBDe4OyHvZRF8IJXtqznils9JJVrQE/pDhvOvVY+YF0MUtTHvnwEXKRkGdHs
aOFrOqkeXty4N5Sx3BCsGQzFdTfFEMDtCGMmvd56mkrDeMXUER53jS5ErWdawOfI
PgZTxWLFnHVnirJpoVIrZTmUQrzka1TpAdQEF9f2UoH78PWJw15VkGjTjAgqua4t
RpvGIPxwclBLqyS4eoCcchDEu9l/5jHRgj4yMV8S6JHMR6sabu1+Drvnjbs1Qose
joUor5sgUJHCmRB+FFUmSqJfhArtP0dDAC81Yq7k2N8CKD0ZfqJyMXSHaltqYNWk
mgAVdDOPxI01EhPVM/3C9klu61zKc5AxTm4RqNt/l1JCLtCNgSAjC1VnfbjDIcLY
gOUV2khNbg2YZG3C1hbfC080qVKMOvg29ysADjGta375KFLdPXwgUylyVoyM3iZm
i+tWP327mcyGXeUrhYGid/BZ/BsX5GU4GBbHBSBzW4j0CxLaOaxqVypJKk/0UdVl
Cua3fuzc1qo9fySJiO3LNBqh0hg68VQgr86hJAGCD5o2fG85NvkjfbDpw0c+hz0v
vmTQs6qLZV2EM4eTyGRmv/u3defgbVPB+KmeVbhvkqpZYCuoYp3mLS2uvdpIpwhZ
+8vqB84v8UbOmak3vIAXR2ylB9TWS7ual81ffhEnpiVNidiGXwOCLj54WEMMBh9l
4hBMIVA2MmDQV0FpgWKPnC7g/ypw5f+KvQt/b95e35w7DJBeOytyEDtO00NColg/
i63jS664iSmvHPP/UO8BdGN98LmKdOb9hkw6lAwwB51Gd5DQrCS424F+SuCzIK77
HjxTZnweDTTMgQZ3uhCHP2cRDpue554RbmFVIf9ZOnal4n/ZGr+1JoJOzzMyd7X/
siLdmSDJO8fNeYgnshikT/U18ihdSfV3UoYGp51x4a1+ile9T+F6CYvdFHwH3SbC
BUQQiBNWA0D9pS+9/MBn2KP6Dn9J6IH6YiD34GirqyMrhZWeAbBPnib/jdgJ48rq
14IFd2Q6d5YFgeRzOwy0hzySef3QNs3tvhDMJ1T6yKy6ryHdfcqSPObYQa+bXORi
BpxB1hOeSvenuWdpy0K7DAfBoXuieVyRkQNB7loe37tyHREdXIkxhS3fhQo1Cm+2
/XeI+bJ02v7XlG+JVgmhXRRgVHaUpeuZWA5s1w/Fnn+njHsrrNa1ccckzcqQwlZQ
L8Ea59K7C9K7r2wT8YpMrcW44etmlUwUmjFTup9GVx8fIXOBzaeRhs394/MXZ639
RJ286Kf2XW1P4jFmU7t0C/uiql2vOffyh6FzWbulO76L8Y9I7Ix2Wv081JCSUbnY
cFqnRg6ErPvS09ZzsFBS18e1aK5DQ04b54lBY8sVMRIbqNC6VkL6Ak2v9912A88U
6iaLazPzHvMTKm9TMkpdWc/QEipaD6/hsyMciTmj5r9nv69J3AD6JmGF14rP/5uI
blJN+dyUTSPh36W1JIcbTUjdb0N/o4Q9nRJuxQmI3pTM/dYdCF8hVOWpsTUWBWX/
XRmuNiYDt2Y2V77zF0cQX/IOOAksXC/5imDtOKzHlmKEglxxvOGWQsiu4gh/Go88
BDmByvi7P29TdfAGPZMoAHpvEDDUvkdQb38I9eHB+u2NJdN7EtYpzy10RhGC3oIx
F5hT5Rd+U8x+ppgVQgVp1HtMdjzEYJJOGQG0yrAEunLqhi4Z0zgxr+s5DoMMsxIy
Bv5BzFqeaCDIQ+/PBCg8k9+6bhZA9KhaQqPXyUcyI0bcnDM6UxvTRzEmHUwU8QTP
LNC1mmEK/1srCxJ2gaP29+OlSrU6OdeLgp7Fhz7TYF7tZR5bDFcObXASvsjtUp8l
PLjvBe8NTO1Uttv9k8AXFEh5fSMqe76RcP9XLEpLS8kfzmwWaNkAqXomgKgoliB5
Pr6y7STFkGuKXbJYCfkQTN6AM8Mrz5unGWpqmob/jIlF0rPUv0fZfwd6l0ExjpjV
5Rqxq+7aGKjDkx+z3U3a1IzavvEgFkooTf1TnfDn6DN+pcd2Cmm5BfNgyad0nxIL
p4OdOlyGkd4Pw9Cae7lbedILULNGAG2cENjAOIOza05GtnbR6EPoSa/vW/ISrQp5
oQW/4NJotRPCbAqOTYYbyxstMi1CH/sWuJihlUEORj4dTjvNn0oOKiB4UhEZNlAc
1mTvb/KlgvHhPRrXESU3ns5lXLhVmKEu9W7qdm33dEjxuaom0G5SUnY2g7v0Nn9F
i+Yt84CVhDsyoOdZx35QDPXgH8rQteJnGW4ZQJ2/dhfgB7PRQFr9uXJqK91pDcut
hJwRfSJQ5QwR3gNzUg819uhw0+vG8Ql3wiE/udOPFZT8UMRd3Vv/e/bVm1ai84wm
AsyaauVumnh6yaxbx9xRVl8TBuRZIKhXKfC3YpWqvneAKyCRqZKwBxCPdjrYMXIz
+Fo63fINbE05ckgDXztI0fkylb2njhO1mJiT7GbxXlkcUoFqK/U5bdRTADyFzkux
PPlboMvPhtCi24s4hAgH8kkNmo/KQ9SQ48rrx5d5dp+txVGNilxWTxL1yFNmLE6H
0s3EGvcZ1XFVxv8bkw5DkKhLK4pag4DFY4NNBUfwKJv8SxUD+KxB3+xtsAc89TRi
DgeEfHEd1//WLc39iuMYKaYQt/y9Idrqy45JhNbDJivfV/6zGMltoc6ibEGbom/v
HP8I1Z3l2B2/9VavgZZTGYrnjD9npo0bfzC/6ocoBDMCbrn53xSZinqwJLzTqhLz
9Tyvj1pcWRL4V+cgC967768zGalLBPhP7ZLH8NVRJBRh3KpG4dy1xgbCvRxYGhUK
C4oGhFHjjjbNWeSy/U0iLxAHpPytF9m1E83Y5lNHOmFA24ds89/uoVxBUXs8FoBZ
O097Trldhrh9xeW7iXFMP/mIcuRELP5cJkKn0wfOQgZeo6oj4P1gV+USoaPJMCs1
yn3Xiqk4zfnpWB/73EPMbmvirIU18Sx3nxufsUI/bWboBYeha7j/LhaIMRkP4Tad
O8zmKtg4QvZKhVX4DgcvkSEwsTJn3sIR3zIi57sZuWLewBC69CnE7/6HahXNgvXu
gpkv3xGLcy7R1XTDz46cUw9o9prSC0vvdhyTx59brwxvPGUKdW7AbExb0Pj3srB0
8joSR7B9vyoAj7JylPsW8saqIuf5b1gPlUNwWuClJNB0azOVo8Tui8IGtHh77EWm
sxQbTcvJ+wm0TBvp0kFY05f5wa+Iizu8vtO3Wu11eLYmlphs2W98hhrIMjhU02Mt
UG/FjnsMrYN1Xkef+FKv9bfPoW0Vdd/iHRhvnNkLjn2WL17wZFKqBrcXgf9vY/+u
KVRcIS++gV/xuyurj+Jz+MxLhko49XvejpbEpzCJi6+NFfk9uI/MMEkBwX5gkSkT
yIpTDYS0FuG//LMWvd+laYT0h3PqJvm7dO7WgAm6KNYBi/qK853PA936kRv3+ePY
H4IBXXpHxE43LlKpSIOQq/E7WEubzXhAaOnqFJ6SKYapkGtexVwGKgspXiiALmRE
TtXm13KMcKqUGBFLPNFhUzlsuZ/wrgrGwOwfM/asEZyVi7wXuDMb+gqecQ2IvKnZ
BWG+ZGiI/Z679WptdckPA/cI83H2l96O/BLh/sNGcldLzBht0pcB61YO/qielZBk
Mdip7VK9efw8azaZN1NTuVdX7/OfiRIA7lizOqNbztq05W1HZve6kLmIR787INdF
weDHpLUMdeICUjbfGTKlwbr/vRPGbUdRNlsTZ05uWZhY8CUbvdp02K3+3qnEHmX2
GXyeWw4v7uifimWRXDZaPU4TXRv8AoUJKc29zUjQvtgiivaXEjE5i4JySKSTEyu4
OimmB0AXVp/Dc8z0q7zwSu+QD2Y2fzRt42yOWzt5hPyJy4/+lHGOIXjPRR3Z1AiS
eSrv/oH9HN5WA1LJfLBIaNYQ200Adgl3NKabWY5C1oTFtorvXmLEM5Qn629SiS3Z
SPqhrqBJhhOVk+13l9o7nwOugWLzmBUhioFKmB3VVIeFnjklYwQbllWW8cOSKQN2
BSZTR3A68grq1BPC3Bwu7GCdti03MWmrPpLBCFMuGuhLJ4NT/oHDR3JsY7myIz1A
lQ9BTIPjT0A0pq68UOZQ33O5uDmWUcBod8/LCs890u/QQA+/+VnoEw7rmwhkzGYF
vQK8jgGKtDzZjJ8fNdUJ+kzPpDaIi+WUWFMGdrpmrm7YsBGG2swdIAVPqDcRqGqL
Ks2LF1ucCU/BHATh4zWRhTHGJ11PFuj8turF/2mp8TfzuDHZq2yW0/Z4km2UyKas
+Fmw0eqUUFK4pJ5lFClf35oSYYk00tFoHJGbSdfi4R08YQnELyl7S28gDdvqFiNk
NA5ycq1i+t/eennM136QzMxGPzvypnNMANd2Jhi+y0/JKMszbwYdXLbBJmCbkz9b
c3WOLDw9cJeVQ9wIvlnJ+YCECAkjEk7+hN+7QBjCTlfUH+qJyoDyW4hO/M1l9QIP
DpDygiITyXov5p2UTSsBhr/OXQeEdjjaJLmMA1CbddDF3ap/HUcooNkm5hSx6FSX
10z98ZlhMorvqXsnPOsTh6KZJxHW64EREkjqXQdFqbjnsayMUxwF5KAktYMXHd5U
xvdQHneZPTgPg6vaTaWKTXMe33uf15xj3WIGPEUIvySXl3Z6Rn+4FFM/8WWL1n+x
PS9xRtQh1A8Z9/g+Pn5WOjSObjTpqy5GIYxkm2RzfCVVjHMsSaFX8kVYhi2O+Jm1
K7t16FclaqV3AfHCyYqTlt0qaAxySK7uRb2hyFxDcua3rBoPAQWhG0ZXkhxaew6N
dmZyYaAk3/72zkbx+igZEa71n7qtrHr71wEaciUT8+aweU6Ag0Y7wqYutxzd5YwR
/3iUIkG0fr+1s31KV97B8nWk2GaY6P50Q++DpHRUzeQVuhH48hCSWo9KUl6Be9bX
IQ+4yDbXjPT3Y3oWforyfKWmjnVWr0ApJSgj5vnZ70jNYYbg4KpDu87ULg0tF4Wd
GOx7W4U1HPHIK+4F7B0giHnwsqYy16pyZUvCgIarAXx7zmFkQFG2lu15XqOuNXTR
vRQAk8ZjDH5tvT08JtHn7/KqyjzUn8UwjxPososEEz/GbVzCWFufyFgYNKu2jm9a
HTRhFotndrdtn8awABWnBQCnnVHa+3pQPiUOmOgOiabFHuHXiehgQqIgH/JGRMw9
gM13qZV+Kxtr8YMtfc/ZgVXV3fvXrj8bu28Q0UjKoDaUXrhiqgmD4C5ztiLS+FuU
q2K7pExxGMBoxzB9Nf8/4ZphRjRFFdAkuRuXkCQ4UjOT7qvK5x0h9P31PD3py5Sw
HTRjtJibMZjCvJM0RJX2DLw1rwzYT1M7ujExmnR6TBaoQfs5nvxQ6dLHQPE1McAa
Id9ZHQrh9HXrP71KloEveGWBraD1IISCEj3ZRuo2lYyrtqZJ8/UB6xPRx9TM4mMh
bxll0wBV3Q8DdZw3WoseB89DCGWYDCrvGlvXqo2tXCCL/i0BzPuthikBbg84CDsy
Gj7miskldg309pc0UugLJwToa3oSc+USQGGRy5FP/Kd5ijB3IwTx7XrURph8VQHa
bqcxZ4epY3CMcU05C5Y2Nwi39GaC1uCSwYVIKeobH8ymtHIdlrFCHzXVPn07ofZA
ub2xuHKK50FW6H4arWkIfBy3ORZphIvlooWmPRYya98kpxkd6aNhQLuaianbljaL
Zy0h96YbKiRArAKZRYY6Wg7yFtK/FFMDVCaoRTq0Oq+HttidY3gdECSExb9k7Bi7
Ik5/xGHK/1POS6dHV1XsOlkqnbga/ZX1nV6r9ea7ZpEphjx6hVCBtety+eDz5ZFO
tEQ/xwDPQJB4ynTFbU9BPJpgGsAvaSqmwXXp5PYEt/sDYp4TDLjEmaUtmOzpEjCN
9uS+BuVBeuTIgb3Eo35pJkKuFXknKkW/KhJydlOUEx3YVDtyb1B/d7mwvPazg+Ew
BgRm8xVxdtshVOQVzEcPx0LM+yRdW4VbqmZM9kLjB8tLGZHtq1Ey3rW1hkLzBzA6
K+uZoQs/ldLZanb6IgtPSENLMsLv4Qx6nHrus94T20Lt30wnzv+sxAd6XNNMrrYD
lL1Dn1XqhMRttqdvZN6ZSYhklO2YLo3oI+nOY0xlP3KWXJptopiBaham6gAJd5+r
nZ6y1pM7qo3CCchgWeaNfLl+mIo6p6mhyJyL2o2bcmKhX0G/IPeLGQuWAH6IKtlC
23P/artaQ0IBEjmr2apqOSYaoB3fI7AsaAu813LDCmTFwbAtuusfhMYW1LYCtf4j
wBd7sUpOE40geurg1sEkQaV+geCGLbUjbMailG8cISU6D8QmNlExDZmNBTFkALEg
ecCnrVyJQSOFReKb/asQc59Qzxo1h6WiPoNKFy1fyuN8LEJbk6IZ/+vztmC3sFNk
5UJ0QpxPv+RPI3ChBlgsffxeEaEpFB9v/765QCP8XplcLWtD3/nlLP5pp84J7uNQ
Xf9no1tvs2i0W/BWzLd7YUoHjtDr2fJEAEtYWFUQe8DqYE+5/pdsxDygXSUio3bE
WStjE86b6I7H43fXfcRII3PES9piaAbvC70rvAKzPGs54DkciEBP16azfY86O56w
K4BUDmahxl/zRzoUFpxEvrXpw8m1aeWu3U4PwXvmnKXi2ajCDTBF7sTzlAlCWJVv
lfRVzfdVkoQcIwDLaZKPkWb+3CcX2IxzAdIVYyaWK3DXJbq2G3RT21Olg8wclS4O
OK14cgkfZqTveYiSGRkxC3UIuTceOZz0FAaUtEt9a32xRedjXYBi2Y3mPJidcRBo
UJkF/IkTAM2FUpkumQtF4cDM40P0RC2gH9mJb8OV5wszLzL4cvGHLdxhkkUCHI/y
YN52Dtviwxkl/T8DTn2YSHXqj8yBTdF+awjTzJcNGFkUo3OMilax/xJTiPLUZMxO
CVGxHwLsFpYEkexa9/76FkAUccnUpOD+Syk/+BVUa7EOXRavQYtYfonLeF99jKga
CscFlNuxGXHhbnkMLAOeWDA0n6iM6YZLsxEUiFF21X/KRhXOX0xNlzRyaFe4Berg
Bxjbcwh8Boospi8rz2Qy169uvoSaa0FB2TYDpE3/Z+EO443AsjGq/6d65SALOEje
rGMWB6048CRuyAhTd6ahD3+j8k50X84H2o9dprknxHRbKdLkubSh5bssMIjXQSwY
gK4CJONYOVh5uTDxkZK6ZTf6Wt5rmvYlPueXgB0MIwQVQ39fj1gBbRtKjJ6jA48w
PwLGD7AnDTov1wvIvMvEOC4S8dXhBzPDpVntpeUacHCjv26sqpC5/xHnrCFHqtus
iZFb6mel2cHo+4x0SMsx7R07aO7Na0i1A5ZKjrMOqjgyjbjhGcHodsCU4UeEWVKE
E/aoJ2dWFoL6B5b68vbGKjpo4if1takVr86wVdLkmJsWGcOU/fZPhMkPFoxYpF3C
Isf4oMsksf7dirFbSVVMyXbkFRriZVWQ7PyG7ydGCmyHstG4Co7ARJUURcUnjsm/
1/crO0ReCmy7+weoiiE7dhG28zL5dsi0I8hgUo6uEBpWZTMDLB7Td9KoxSV3shRi
51Ob8PGIa9sdQtmzIJYUAIg1E4aSh859csEawL33yxlpbdNL4nSVl/78nCi0dbPL
Lo6Vf6Dq51GXBm3LEGVqruaTB03heRv9V+uEGoG++4LEBMbdaZ1PFy+NxuMPT32m
1/aj+s6KdgbM9sifgIQdoF7yRjffsLIo99CYzkmItBAPp2MLv5ATPg1RtL7/jI6N
gzvy3ZK0vJ3UdMPCE3QSVKtbDNOVRKd27zSbB2JqttOb+HKFjsbnLJobQZgnc+NX
Jsf+0T398SVopkee0ENcE7jSaoyxvdpMwGnlh5oMwoeao9acNjfKPf4fX0ymF30U
BStEJ5JXbkaz1s+MilB/iYnUP0tJvn1XwBVAmBUr+04ttATtHnVklCPM0TSBaAuy
ABVB4eOnviCN/feIz03Fr+2f7ACHYXlrmLMBqjVpJzRBzJaOB1ENKEqdU0L3dP5V
etNztgqqrxzLrY1CXKv0Va8BRdaEHwna4jFUw5iCwWkudUmEvhfRDj9das/lQpS+
ohRNxHEn1OMa/74SFa9SP6QgnNUtC1MlgRXgbr3jaWWz3yl5OSSMcq2ZGfRZr81q
daimMnM3QWICxJFtFDFrwoNuBHEoUmYeVfkeBN5O45oxJuaFhEHpuckfLk0UVBNF
ReFUpIOt1vGKzaKroMLsfYwv/wHgR0kA1JuDPo91MziwB2LfZUHfhqfEiudmVoyq
k3q2P1atO+SP31UyOFwlqwyDXDOE5uRNbpVwJWeVKdUjaONAeQjpZxvot8ZyEzq2
v1HOrZfD1Yp9VVXUFebKrNOrxr2QniB65d8q9th8KCVlfY2uqziLscktmfBsiJ93
4Vrt5ebIVeP+5JxSS+l57X1eGSvN/xpEaqS76AOn/vIV6TSSvV9P+c5OYeFYSHJF
0Q1X54t6y4jI6GCvQMaOTsM1S4LM1VxcJ5ubbWmZBrces5W8Ds7KPCSiBMxSjalr
QsLHccaHWlskFHSU6KV3kNw1ELi7cEBuWkUgoJN447+yUGIMUkIOruOCdK7kRw19
JwCYkYFa2NR45niY524S3q1QqE9o0i9Fpm/4pvATnfMjBBh3GCSHvsUiiLlC3TXl
1EeqUh3UCa0XLpVPJGm5kNdHQF4+q3XbpQUWboDAm/7MOyKBzNCvUkbONmgi/kTY
bHMqHFjZs/bsFwEPC2Md668wrG3q/Gf9wL+Vg2a199JjSlJyN7x03U3a5oxAnO8B
S87RXfW3QAkvWGI7jPowzL0LItXeft3IHuRhW7TCMgnqX8vGjwE1Td5Ij31gNipW
qXbjUy1d57NY2Uwtu6RUDl/Rhs7tKNJc+PB0oRwe9k1epE/EQNoy4K/StkKW9OGW
ImN31rMDuQYMZsQrCKH//4/zKj12+N96eJowgselXMnce4H06qkSnyPSWWVfkqKZ
xCkxtvdAeJJpa+uj6vZbFPyxTsWS8yb53hdNM3+wurvNWRdt0oyy8wT1Y23cKRhv
AWrq6XCWwU+wXNpOPj7wBfKzbUPl7ptSIKtcllVXea8v5jAooPxSLO6MNiLHVMJj
5h9crd6QOVVkTrm5sdHcYDn+jujFH9RAPFadAlIw5nP8THllStZ4p/MZpUTARIYV
c4YyYP8456msmp5DQIa95M6R6Zlby0VZNEL6iHFWlu7XxFil93v7NY5QiT/DCeuQ
pnellv71RndwdrXmuvDiuQNwmH2VT9PapCKvv5zICO3w6yee8yle1v7xOMg9obPs
R9Gu+43zOPgR2WRo4TOQNHsz+JFWGDvrY1hQF2fOjmeoBLO4MWdPesz5x6AMNmGi
mRRH5i8EdRcO1iXJSHoA3/roUTvLZWQRvrj8uUGd0tXeU7OuqQidElm+dSw/Pek3
6rk2tyJCYlQn4Sl6WwHLsa0SglW4HoHJxBtqHNJMo041Iyil1w9lOa8HHhT9La0J
av+VDmiiF5l1knda4lge9QMgXurZFZ6dpj9XJfetdbpJm1GuFEXwZyl/G04rm14A
+aYinfZI5EXFQZQK+USEoTtpMoH6yNFqHVN1xgTBIj2SMmYAZRjuCG4IswwRQYYr
UM1Um7jVDOdsEpJfjiqyTPDTpaTxUhSXPRFQdebZUmEK44iSV3eCJaSIH6R9Nojz
IoBaz4kFm6PTrrZBg5yxp7XjWsB4qZQ4F4t8CAsoQiS5EDbDULF6m8l0w/acmzEp
11MPSuzyj3JeD3YxODXh1IHlyJCWjY7DYsNTQSBEuo019KKOoQdN/hidGqg0tiqu
FNdTlG9DADYp/xRS6wjyxYKbT/CfHzHUFH/8A0M9BTrV7I8/8zyVE2AS9JDp5vVS
f2ASWTcs+Gkl9B0aXNYflV85jG3Zrljx7161Hu/J00c+8qhis4jZvL1t2HlhSXnL
6/U5/+6DM2I034SmnP4Su9alWZ/oUTGUGIWziWvSXTC2VEX+wBXYLB3VKB4MoKyA
q6eLvUkUYasq/r0vO5kk9QmNLu9pKTqramhj3IH0OH+4EOsIC9gQ75tm95DigUHJ
9eszMLk8jjlDHCLcO/CYwCcMXWNlrEWd9YvFmNeUZlUaga7V6qCpqd0BiY7Eya6F
Ji51UMZh1ukW7B05DQ3rWqfs7W8INSv6X1ujWkpy/QPZ+J3uJn/Qafa/qfBod8hn
Twz2m/1I8+73jwmcuUQ4/QDlJM8ZUdkrbHD14OT+ctQoyYfjf0Pfh1CzDFXcSbYG
UP7uS1iMZdkb0zZQ42X/PA9FwQ70AO24FtBj/KkShZX1TVD5THyf94Mq/G6LiNsp
lwl+OkZBkhRl2cyJulHpqMUWlQIoiKsa/HnqNfdYqols3aGcnPnUs60/zFILZHOe
xA/lpPhWW9FWcsyimC/drH7f/N2zXqfUWuqZFTeyFzDAhsp711lqq2gmt2A7q1Eu
jWUcyq4hfmB4uyK4ERkxe7fwjbClQySEVK7rrz/ZP9XddHH53TBvogci32D3Gk+m
73B4NpXZhtEjmLIIsVPrg1gOxzLHld9P9BTN15mwr4VQ1zqPiYVOV/S3uuhWkJPo
Mwft5BMDDA9JDKJB5FIfd9ogXxDFZy5sM5xcXh2LIAWUuP6X0UxG8/esMF1CvRoF
BHUV4gL+NV9XAf1dAdbNeSr3WhbE3xUPGlRtg+2wckR1tbB5EE13UQ3HSf2EKcqK
gRWy4OYzBtQMrtewdcROb+pnR/aJXPvWyj0X65HcefhC8DhYnsI1xAJce+5x+8+c
Mi+aH/hsENSk1EYjFAgctwt/NNSLO/vqale/F4fVOsYLeuYTRm4W+0RKKAk835T3
unHRXJiakUWC5y3Y1Ezz2vYA6QD5ghNvSV4aPxwGA+P95a8RBzYMy9x/YY9IOq6w
jNF0zRRE0RUm3ri8y79Rp5NZIoovaSF5JQ8o6YAVGv8cXm4dOA2tlqDikBDxF1Mp
r3agZXiOI05KIuS56QTMcv4Gsy7mE7GnZwClU38ARHP0bYGpVcu1ooPfEhvva21t
/zCo/aGtLsOtcEws5TlC6XlSUlFRZkX2LF31o0jzadGTV0AT7nkV93HXMuXQe7t4
MtjpwuGigKXGkDUa6NQ8d9aIPuFdARsBeTYezLtBV5m9MI0uCwuzflydpkLQjWjQ
y5JPpUy4iCvxqYQukOQ7JrBbnkKnylgnv7/ZnrIHKfqDE/atVkXMsi392199ymuL
Ais3jyhVzzkrlckKCvWN2gV935GhLyO2IqEWJpddhLGD8UTIQEBDb++ANK7zhRYA
1al4dzl5+qvV5rxhsq2/RjcD6J5on2k/h8VOyjHmWT2C57F19ZeMJt7iRKFDYkMf
CTBijmUp3W7/Nib7QUVoBKrk0Y6P3MejuuuAjzinq8XEA3VS6Amykd6U3RumreTA
NwHQA6+35hrfNgMOaBs5jPwOXC3yuE7YqmtfMl++o3ZgDyGMO/yWhr35gQXCaCZZ
kawJyHkYlL1VJLxzsdtEzYyHAbOxKa3UK69paJLmI6+oO4UEdYmyZpb9jwgrwfH/
VbKLmsacOn66+JmBQd+L6IHiX0Rnz7TeJAGZhl8xAwcJD74Rz53kzrlFsPP9iIG5
0326wEjxl2QhNYqRoU6dDBO7RhnHpK0YUVo395EOVVxp1D8kM5BlXsTakTTBx5UI
926q02pGW4mYcT8cqnC9C8Wre49ajhT/QXw5+ka7lPRf9dBO1ywXjjDOk/kALn2b
eDNcfoP0tu1GnD274aXMh7OaKvIB66lBIqqkUsZav/fVppzyiVNo0FeljAv699so
qZKFcO4iKy+KpCqp+TVkOl4uXpPWtA11uAYgr0Q9vWW2/50fq6C7bQgIE6pjjEIk
jfWm01cDGN0ekRt3vU7Rp3NHhcMq5iYjP7LAmsUUliipdaIUV0WrRHlRTz812AFG
odklIfH6I/1tHJaSYqet/p2/v2yHEeAtzKcMT+68ojBDcQmLeiAE7XXjx2PHJiub
2YsVHYJN4gIeLRHk+gBL+2doeTGo4Ts4yzq/mYgD0yi0YGKXKVWvONYtwBHXQdir
IWuZ86HKGI4ybHfzGdKCIbxW/ax3Z0FnV6C75C8uInzlMzQgM4clezgS80kNIdgK
LB/tIx0YKvoHfjxNwC6gjQ7TG+phaP3Gx9qjHpgcZxU6D5DyKiUiOBY1o034/Pra
tDJJnlpYb0XkaTP3Dl80F2T/PWXbvnZDIPpnXsD5wkjuRZ6oEME9R5Ixvd0XEsg9
BP/Mj2CtB5CP206gNDbzvZnPAsRjunZt6RKPfGw6t7nPK/iLT/7mZKjXBQQ8RG29
fkd9jbm2S1dwGOZP0mS6PEv5imoMOLGze7hIGRPPF7NlmQ25VgsR8b6zGKo9zAw7
RuWE2sfPdX1RxqmFF5fIC7c8O5TlS8rR6OTycQw/2ZeXTz3UFHpkbZhL3+rrxKbM
oLb2XSIaoruQwIw13eS6x0XKsKhtjf31wES1JS5Bg1HlkYjO5//J/AseC+Dojw3d
dCc14n6oY2AyVZ4acqAlLi6cKoViewN4ecI0RQb2OWUXIoRh8VWUWa5xTPLXvvSC
+0AqxnlckV45NegSv+XMNMVu99ZZcPonRfRCdlYghAKhYQK36lzLbAqHMnVH2cSz
Ay6ViE4N6dK2M43J/BjpLeYV1Bwdfi3JcktBjsao3sVORKJTcnSPRH5KlDFqWaaD
ginSRBtk/v7RWbaoEu6OtaTlXFQXzldDo1kpgtLtQ03o/Ia+RCCDbQOo7qLTSf4k
/0Ch4+0mHyolXEvPy7S8GIMytpyF6rLbW3UOKbbAj3lFLKmVwxSB63Ub6i+vyHz0
aSOZBjlvTQL5KhKOH2VZ5jgmhQcv+1iiqV5VuRFZmrWHyknWELncdpO/0bXzXQeH
SYARKKXk4UOkoMCwGJtj3XWos5N1fzRlA9ZXRDwI2fW3f5nQSjM7medL3Wvhb8dV
rqMqV8T8N4Zg+gcmXK8Zvhocx8rWEM2wVn81K7xwtPsHrUjOyn2Somc4piQitSdw
goXepP1LZ2PiA+C/eVWvny0mLXWdwqOqguHVeLkMMUBX7G2nEoCXx1UYWOUWOIGP
BIg2+5JNRjcmAqZ41UYof/rscB/hTDoIAkmdyT1ZMT9nIwqSF6AROQgKAHWWoYC0
9ctahLhPZx5sOPvIh/Iv50zzQ/Cu7F0GH/wT8i86llQVQ3JRTpNN708gM7s70JnA
sYWXrMyLntz3Dmekd6quJLnn8ES5/Ph3yC1mIe1/bBeY9RaZAMq+JQ88DUA5ne92
zhvXOSdk5eCvg/0KGHUBqroeV9NdHB8AaBEkLc+88K/fTPSDR5d0CgHpkPupIlwe
tyCWMLDn0481zBzJu3+nBYXkdIe8lfxxA0bUDx4PwZ86/LzihDc44ElmR/DwB0Rb
0TaX1+MiaWP4ASpnA4sZWnwW5cRLujfalaZe9YGOcKmlki8yPV3YyFKjNRKuHuUa
69w+fTA4sMIF0Yc3OG8RtDJDUH006c69hk4AW+T7htPzhsuXglfV9Syw6icyy8ro
dB/hn7yT5SqUK09mg8vRIIRqTL8blbB8bzLT5QWSE11ieGDJDrcE8tM04hDzGx6H
P5mn3CfQxT2SP6oh8CTnyJndCc9Th25OvdCTAf48skTKxlkbWorrI4nxKoTkL9o3
vfcTwMzqX2UVf4ZWIzXAuOvVudVsn2E8qFHxN029ybuYQbG8NE2HndWhWbcMztdO
63xZDetP5toZZwcx98TcsycPJ7WgvHn2leP2TWtDXJtzzhLzim4d/S46qpTG3DCs
5AgwopJKMCUHhqe+INWEdja9LGYRz4obLIFZCyU0fOU7hFyZcmYfpAafm21jTc5Y
J8gp6nPWN2Bt2tRUQayyvA3N4zsz3X1dATjtZBjZzn7aQhW+icQ+c10U+HqDs9Rs
V+wmvJiI715kBP48WfRyFeP6VGvld6MivOPLqO/lwst37/CRN2zPE8oHavl08CBY
ziBnWLaeZGEgL/2g0xa+c6z3C32jvX1rSvsWg6u1IUznJk/B43DQGzPrOdTybYib
e5TJgqJY5JGdp3PBTuoroQk8aSi0fRhlb4WJI4EbFyJ7VRGSiWSQJeqnvNgeZOni
Gl13et0SdWeiAKU8xsKqryl3rGL98QkzzJp9pHuAykZQRqFnBN92Nt727xAnDyYI
IxZ6i1THyVc8cPKuEU+ye7YxEgYhYjhqhppe0VVI4be2de+U5ecXj7FAYL0M5Pl2
6M2S37mr82AJS485HXhX9IhL9NULI3c5eKTNouEIdgeVX3SyTe/yVKzBWzrxAy8A
9qjn1lQ4Gr00iNi0wB4avNU/I8prgfFVAUZxmKEj37yezpw7E2ClprvWyeBB2KYA
SKnTMOXbB9n2lFMR1Hf9sQhEoKH+4bcILOsRplY998o4ZyMiLJbUYr3MZPs2flT+
XvSIIbpk3POxixwRFBrbsR6AOdH2chHaUO66Y9HQ7m5dmfPljFJ9ztw5xz/uMbj7
fLSnbIOpiaCBgAeweJIThOb2uXPcW3tJaxnZOikG/9wz3f1glC31m9cvxLra7uU7
/Dx9yMjKPJoR/SUR2ix73GyiAgcbycx9sEruyW+ZaTt4k0jhoTG7SbuQNRRRkGfZ
3FwmmV6syxu/CUJ4mk+orRlNXFNgQvhkN/7DBkwqiOVkW9jx/iLWs0poGRENmVMS
JT4yHwUggo1Fjw/4cD4Oy+VrMq7jG/i2ylS7y98oZ6DOMP9eqcqJJ4twLIqJG3U6
WsM4wIVo1UAz1PShUct4i9D+XRTFeCtU34Vx8+V86NghVw7V4nw2T0mUu1LuMi30
hZ9xA1ui9gu5Vacgc0C3hte3DubBW2mS4sAnSbB6et5TuxSazMgIlsZPAU8uG2FE
Qlg5sQvLrgoPX37eEnQId6I0Zxs8/SGNhxokBSe0MlbKwcO/xcGwQN4CLC5r9j1y
RrwCswEnLemURLpTK/aL/6zA/LloC+sKIIMstp9nT1HTlEDSHI8sA6wJ3lauTFN3
5tNtiXHYWRaU08R7kf3DtY0jiFpPfH0CMsrFHtJlB8c4vgLLYV5HBg1BvBrvlWDd
HgDl0FT+FOoIbh9QKIIJ1tS1cG8NjWywu+M07pf77kjIe0ErTHFimTa5+bl5QKBc
5PRxiZq7pKKs0TxDLtmZKq+0+jJ2DXYBQOWliHpNkP8Ovg7jk0FEtmhGqDCBIS04
Z8Ds7oLgIMKqlT8sP6CNig9IFZaj1QYVqfZlLkCgaSjVZ/+TV+9QFIe5rup6h88R
T0pe0LtcI9Pc15P3GE4brEFgvZ3JD1m6bsMHvaZ7sN3CPusMYtEjzyAHF4OTZQor
V7FZ9w3NvU+gV97uQ9iInwSNR+97l7zaFOF/NOMh4H0D3T5MrcT7eBefSiopW38i
ABHI0yBUMm1RG0nXL7/81WE92BhyMixbN7tJeV7ZGpxtPQljbqCx5+VE/xvMgVNF
fKVwZg2O6l/1N2uXByigvA11mF5O0BzjG9LYjPoBKGiTE0ORudmF3vED1Wd5dtHc
qHpuNrmm/TOF5e6PhpaymggV8QEPobjO92+h+tWi5OmLI6ZHFk861pjY0o4+jLRM
CvbSRo4TbKDHN9SeRPNZRkv4yn69P0b6aKVphsNqrH6UkqCy7GhESm0mgCNQ43wO
Mc8TaDT/ebNKx0PO3ODBj6vTD3zVe+UR1VePrzXK2vojkAtj22KHJi+L/JP4BL4q
v50ygD9AfsXzmoonMPYh0gtvRkn+v/atzqlyfiH82tV/gx6REOQkXwwO2xyRbdZ8
XHnxOdrbL10tXSXIWsNzpeHdVO/hHGDOzZ3/Uw0Cl8H9fP9j5KxrXGVOsKaxeKeA
3SN+SVhlzPW9lfsJNwcpAxY3FkfH/RW3n1xaqK9RQN70DhTRyHQR6mqHJ7b6rLlG
30nQ+zOczfvavIV9/nSMRvhTtiR6+d5P537A+dfP3GcaLsV6Wl3MaWGiFMF4Z1b/
vX4GcVKjQycrtan9DBjWvOLnG2abT1VrHaIw6N9+QnDbS8elwXozG2GBpE6Wriwq
V9/Q5f5yrNH0QoLJY+ilaKeCrzuFEGN1i5fVa2yckvWBGF17ySZwJnQ3mZwrWCsR
wCYdFdtlAtTr7uBGndD7iDoxrw/cYhIt0SA+Tw0rDamBGScO2rMw9SsItxeJXBGq
5joqosjSXWZJJQNI09BMHB0TwOlxuxt6K2/7bnVRvQFm4uCwTAS/MK+pLCs3Pf4h
KkwQMDORtbr/adOHnCJ700l9gtLeGsteiqOkm+F1/tJKE9FI+aVdurkYowmqb8lK
bpG0cWjIUXpaiWP46Wkp0/8LmkZSZGCdePn2VnULRPlb7u6YN5OAqPM24y9C6KiU
m8q4IIgSnur2DxiRqX9Y8LsxD/DsEplHFVMZncoPZtisFHYo+GKTK7UcS81hjV8t
L1B8CymHAt+baB5KRTuQKT6hugYJBy/qw1KQsi+8XA5lV1BHxLAXYFsjm2az7R7c
xHw+fjFmLIKjRmNtgwGxhO29MwKvQDM++2qqlCgJd4nTliPDFGByO4z1GEAiNgPL
S9XYfhvlijvU/igszEXggE1XtW6UC1dLm3Z8zhKm1HYOwfhl4IvktPuPpQ1nZRix
SOYJcmwPUUilGV11xgjeqfvnIKRNkv7RvCOiNndXhdgJp63WJyMteJ59Jbl6ALDa
E7pjLgkApfKxQMLFIioXfZrIGcG/W+FBXj/lUrbctdlks6FQx1PJiJ1hr2tWdHpv
6sX0wS4n6MZ2xcFpqaFhoDNRVY/Ym6W9OBnlJbid8NEjRDlb2BNAYwxr9P2xFiV/
7WwU2YwVjnnL6WAKN0SkxyivnXrQJYfH0T/juevt8e5jx44ZjAXZLkkGPr/Mqyj9
IJc3EzGzPbS+7txkJezAhsB1v5OMK+IcHZJLAdNNUDXUOMXZjyjIWCpm3+BolyFT
F3tEbTl1UvFi2ZteaJFgeoUAFMPcDAT0vMUzte4Hwu67/CWXoKc8lEocUPckbFJc
i/W9sGvefLzisrHAvWWI5f1dUXvsAwIDsuFTQRs+RPXYDR1UBqCwYGEJ3d8CuVqn
fup0ar98ODW7wpOhqjdOJrKcSgMb9fmAQt7FDkQHcpYXGTWS0jT7lNOZCUyP5GA/
NWxx+OfxItSMPoAvBBcbqA35u4D7iVw3LgplrQkDOvolqeNGXbj4WdchuYsBvmMw
X2uiDOk9VgQZcwzIha8FdphUNsaxEqSKI1QyTuJyhfcmWbZ45fPFdXvAvxgNmP2T
K5fW0XDB5lYYxBIW1+st4rJXGb2LuaOSUj4F09KAcNS3Sf4lcLVkmTqQjOWBFYup
27DWwj6vX+R/+L00HYkKSyzfJNSCjWe1gy0pEkcGTzEpgHzV024LDH0AO8aSILDo
AM81QeWS1QwrdFr3XdZAkKrewRC/7U3EYUSA0td+MYYEVZ05W7ngK5YwxTBcMU2L
8aNJUCyQ++DbGUkJlkrARZPrp78RDP9tuSj1hP+uz81ICuZPkwa2xl8LzxhaJiJt
K5/9+iMdq85+0oOIAVoZ0nV0mNcaS6FTxZfh1MOZA2ve4CsWmspvW7fNl3T7QNFV
luqa/GCRt3EDhs2FSrNelnWO2ZCJZEYhLGrQrdqjOOG/t/MpPU4CQKgxqWiN+ICB
hlutZpo5bx9hI5U2ee99RJq7wJpqoxdWp1/V/lQALKFTq9Jc9wWL75+WfXxl0TFk
u0m0ql5RZ3/riTu7XrAFTPRMyUW1O+baspq3a4BLhawJ4vnBQyO+wuBzKETOYZXc
rBR7T3gClDObmK3Mm1hCt7mOXYzVS7Q1V0mhXLVfUVw1/5WsqbkWuwnmjlLNhk4p
3GPD/q7rzjbCiU39KkhyJUDILn8a2xY1D2OqXNSEv4/BlVZOaRzfFC9r7RmJEKc6
s567lh/uAANL1yP9ruQsMXwdh7NKbEKiv6CFmPFJ1+i76nwSkUkygMNONP73uZ8j
GwQEimd20ZjyK78IZSI+3jFfoWIW0Vr39MUUkBDsAzvwk2B7IMyJFGZOIA5AJjlt
f1TAkmLCIfjMQmjf+0GKX6DHgzs7DD7UCHjpD3H8tgUlbtohE+fTIYEnIDJ/nsah
jZCIM3lkBGTsqu0Wfxkt1ZPD/6vZj1mjMNZTYYVqHHPO4wNJCio4ewWBvrhQcNdS
ve6LBqJ0z19ceJts2FagZ1tXdexrlyqSs4JTe59Pch/52Pvp7hv12t1eXk03hyPO
f8w4dKzTvtfmx1VhAOH25DimouaFOpV5YNbfdQ9kolphQlD1qjmikPcsXJ2K45wm
+j0aP2lB1TcKaAO6T9hHHipLQwGFSeQo/6XSSslOu4bk0hKijyRlD7Cei6bTTMnG
GmvGqY+SImHMnQhs+AdCGLBI4/qn2QIhSllDuKFm5QZGE18RG9OtLhsAy6j6AYoK
ywE/Nh6FP700HqRtFS8P9unv2c0WWJVWWNuxk6WYZMda9eNnN3bI4IwXl7hkaSIw
AaRIPKKajyoCKZE/ceeGFvaE23dX8xERjqr9FAUIsF0vjCjX33rKdgzUXV/PNLdq
qi+fUttFCRg0vUzYL3qUOzwoyX8Y0o//bneWlGPF+NJ0sP4oz2Z35PCkfDJOP+XQ
Pt76Bwl7avrqy4N7kjkbEb9HxTiqH+BlTYakKCd8NJ3Hyk0IxuHuqwIjnrU/Tdnk
Rgm+G/u5xvyr7rN0xHmZ2c01Gc/u1Hs9lbbeaiOZLY6Z4u3y445tXWjn+ytooQip
EsOds78wcwRGwTBZWYGj3rqk3xt/Jpcfhq0PHSilhPkGle35TFqyMgi6p+9yecWD
9HUKrpcVLyzKBw0VtSRf4sXwTL+BWTncHW/I8Pv6Zo0h6sH3d7NOLe7H+20Wwkb5
xVeCckd459RyTROEgxmoz8051Dk5cHC1xyrGul4yUwjZbFN3LAnGG+mRf2di7EFL
e8vVVso0ynn+fKfkbz9SL6bsPv65IzRStgssTyeCu6OQro0w5fAQ1tCo/VED92q/
3QLtmjrM8bMCExuh+eprUcXX3dNZ/50UtTsvwR7wUF9K84HHHROmluIDti/Wp4q5
IzfMFlL0mF4RvsCtdVa0TY3878kgENa6F0LZAIqw/TaZZVhEBSE6a9uEIfW4Dlpv
F13Jm/pdLld7UtZsoOcX9EN0Fmu7UlKjLMkmPt4PQ7zbpIvm1GlmAz2fB3nxvNmG
p6iJvXz64sLHjPjwHcJ/bxEJOLYN9ZPrn0NCAloEizp0TO1wooxYrsrd5jvnZmrH
GNIqwEhSz9YUOYfT7iI3OhHQQYaaZVGg/15Tgsrs9Z2o6X2gciwdueXw/LPA8wXH
cFk7bgM7UV+Acq1u6ImBEy7Ih2oqCNybETssu2mQfp/2Futf1zvpebPtnYFQKLPt
uY51jv2KnYtYD68up/+f0Qa2lhwgVjvGzPVSKA4IiUwyybNzcA4nJJHR2JNx0OQj
BJVD90v5rcAEz3XooPCsB6T98GOMer94fmUbMT1mjMVGvF4nViKpKhAxTug1haNM
ZV8uUuKVA4LhrC2OLNNL2zDKH3eF0W1nyhhLr6v3I4ntujjxFU+pl+y961jMXgA5
8hX9T94rKMLEoCa8N6YwDNoqRtD7I1Ap2vNUhoAShoFxqQfrbfm5PXzeglQmP35i
pkpifSsiePEj6zBac5QaU67LLXfs0krjKWQs6awZEwbKg6au/QtGaMbquSG7/fLK
GjFH3YYFf/6Sj/aM4ra+gaguNaJXNZQrbE0IZQ1/7qjTWIABKtWB7+CUfSgR5QCa
B/HNtgw+pFzBr15cB3gf28C6VTp95/xhIfIXVSc3U3yL5p2EHk2R5nUfR4IlPERa
qQO/fr2X4jzNjXFO4gcxszP2DnI2bmCb76Ckc1SoiRLwyNrI3JfLA62qyWAfTHft
Gl+yUGasOgUp5W0xlbWHAriin6TFOUhUKHwf2RNwNAxkFt59NMdfGFx5AMadj2jK
5vI5ugdHHDzBI6lmgQOiCLfRyradsAc25EP4X31AuHRBGnCdmFrl+HF7rxKLL5tF
RdNSHCkOD/5FwWpen6A5ZBS2rudN2d4IXZYl1ViuTF5dwoHDlPia5k1A6imnhq3B
0Qdhc3Uan9smJkLYxJbvLJKhEPD+Keqy7inHnmPXNp2I7T+1IwexsAaJ9pdOdlEG
MCThxa8D7OlalGnDZ5rBEU2XK++pXBdc09p3z2yuFR2DQw0hK/izWx9QJLZwHzFm
DHehXMGj2Q0EJjTHZzsHEgEauPvGN8R+IkrPnZSXavVvw5+rYnFuaKKnmp4G8xzR
1BUzx7QA/qNbPhguR26VE0e/n0gvAKlMLmXgNMJAjiIzpCrT5SURbqHRA5ywnO6A
vQEEbiJOgE483zMLhTVGhWyHWPOOURPtizPOjZHnZhvRSE/PPH+Qbrg17Q8DynXd
Ze3YnfiGrbS5WQ7LKP8P1k7DopHIWEbdWMIwTE66xyoTvPMGdbtOMHurGNujfydH
CgpACuaDyJSzNofp+JUifCQVGhEGNBBN0mlL1b3fDxQ1XIHY/1+msPvBxr4AQrLJ
3xVubEwV/KKCYY1cSbzAUJfeNjDNMz+k+UT2OA/QdDC5/i7sqAu5Cxt/XrOS0s2C
b9AShaX42tuZF14yUFZWMiS1ukDP18H5Wo+yQUoUVYUGfXN6fPbzxY5+Nh2izGV7
UUFUaW1ImecQ2vtygmQGRKB/1e8/bQVE74emSEs6FaUUNbzTndJ3Gygf2bVBC/EJ
xT13dLLvZ34iHQ7LL0ZnIj53jvVN5fhyiBNGZdE8mOzb8JVfjv1xKD4GOCAqkpZ+
WZShA1xsW2SkngrDvYgNEoJOUoT7TblP1gQbBpgwpr+ap3Nfd7EJ5/FDpNXg/Xe1
252bV5dAhd8PQ9oRjfkAww+/rMBkbA5LAH/ke+XGA+Z8eWk/JPXuXw1ge9NjFSyZ
deXl3TcOMMIKUTPjJXZI55nFYQqfWO1p2L8R/535IZs9Lzmsy5HPWh7Ke7vt6ExR
z2w/2WvkdCylrex+ALAknyyq7qtOXGIMDCIGAoBkgPAOPTgc3ZQ41UXNUL4ZCnAW
SRW9Tcv5PjWW4ZO29kadERL2OpFtMsgC647tehgnZ9IGQ86ipncsko+miPuVOQLq
5gHwtvn05tiQqRqHyjocFC7l5vVLGitOi58MDIMpSrDawPqR2h4PAZvZz6barAZn
KSTT+cPsONstga3pdMTBSm+FKWukqfboqpie+UTn1Lxs73hEdUnJ5vzdu05FwHD5
ulW1N3aB8wEUoGhcoC+M3/OJSlhRJT9dDiY3Ete5CXha7Ayix9r1Xi7AmX+KEVFv
fyaW38fe6vVBZtrgtB03iyTg/oBil6umcs6Y2fzqkAL3U5ImNNzgm1DjRK5ZBNsx
pURpwj588uTMOfehllqtidNG9C5wJYwM0I1mxEmo4swf5oH+4sA5pJN3Dfuz486n
KSmbIF9YjsZ7LuWIecMn+gjMh7PoNNVjDXR30r5dxrJJmyepFdjYLwvbfe7iGMPe
TVPz13iDWiSdXpgGWVZ0bi3TUH3X86irC7nBYNhaceY+PLmi60C6aF5az+8ab6lP
dI0FlVagHY4gSmxOzyUHeB5IRNNYvwkzwfMH14GvglnX0z0iigxeXSc1Il6yKjfy
uAka2/IxYg9kbSH7OTB16TY1y4i6v/9HjvNLK+GGWkBs+HZ2gfGGzkS+J0bh6ccn
IzQQ58zzMgM+yRFQ5RqI9+lCd4J4ZMXL0bfZH00si5DL88Izzeg/UK5cxnvnttKF
egDfywSFR+aiZzpiDGZeLfBVCNLn63C/pN5H3kmihsxvaYyEP/SybJP+Y1B0DbOb
+fKaRMsmkKbEn/NPi1njxbGFhaTkT9GIXj9Wjy3Bf846tijC0mbKkaoktWT+sgbf
OOX89Q9xOJcyp3f/nbwnlsNgzKnYZHJOg9bXdcKbz1eFHOaQfaQ8ZfJ5ijaEVdoH
GcQ8xWguSSIVSzxVu1jOyEtXeW6oQbK2YNPOLRjCdUiOBv2v/BucV8SmAkj4SjM5
YFspbU1qLwz2OVh5KL7Xrlr8M2mx++eIZ3PF35R/5zOBmn9zFRs+37oWG1B10IYY
HS3VS/XuVKxSh+4tANMJUNUCrv6s7mqzcbJ7L+9Rsx9gef+6Ez7r4sq8OA6iXiCy
gHXmnynKYD/dtX8BUDnNRLRzuWSNPNidmkcXVhPqQyqeXl+9DvjSsqot7oEp1HxP
q704LCYzWYmfGOGyv4JcpJH7ivplKO10/D1kvqctlqZr4L65fH6I4sAGfgST3t5E
6bUcLrOgQgJURrjaaNDOPHt1pqvIDiQvHOKWrvKixnIqIp+q0J2IoAFBaUhNp/P3
CzmOD075ZafqaFXE5N6TKibN59AK5bY19rEIhYKmDdNLXAONJoS1J6yjJ4f7Jm0a
djUfHGn2aqzcAFAdk5eEjWK0QTmfN/HXKFf1cRRiUpQfug+tkOUFHbfBC2MQRX24
rWheLFQ0VBzh2wRMIsjMTQEuI/dJ8VdbI//nwn3Q6gCxta7c5mPMAOoOOUpBs+pj
CCwDAj2b1/nQ9cvfcnCjJ9DyntLstNl9aDAdO2QAcyJ+iXx2yuDMYx7XljsRqmrs
K/GLBFazh5hbvbh8hiyiG6POVjRdy9Zf1GHXeD1Rcw4BYntGryQFS4bEq9clGc6x
NT2SYN51c6GsmAbipCh1h2ChdghH4gCGCkn+HFZUCMPGTg2f8fewWJSpWdtA/TP8
fRAxlhWMX+yDzYU4Z2/XYgaiQ8W3L07uc9DR7IjJtx9PkCJy2zNTtNfr272Aj8n3
sTDGGVS4XST+KkmuErBLlMQoa0ON3n1z845lj/ypAgeO3lK3EYMj4Nx1a2PxB8d8
d6Aki0ZYLK904jtvnJWo3VeHq1ZqwLwuRoEPnjCHHsDFSOpBCx4LQ9V5sjhhrJB0
o53hnxLkXU6TawMboV3/Rjid/X1myVg7VP3BzuARiTIIjJviUgLBcv+BDFrb+dB/
PLNH1EXQYLiSvU7nKlBE6k68wvWWjdsH4ZQFGUulA+wTTDhvbbpJjQNrv2cIn0Hi
LNxIlhfd3GgcU2nn4ZXj1U0jsBdvFOEmffpfqlmsz7cZ1rDUoQj5qJCF2FDFg3li
nf38XfXCbwcUOlJe33tneZ/wrywOH8AN9I9Or11kZdPPFEhF3ud7wLO1G5GRzQ5W
0tm5mwaf3frRFLtSJCxdd6MXpCNT9P+FcOeNsVGbVe32rwvUhwwW4H1uNmmvWpR2
QBssudzDkDLG+UOWgITleEgVW4BP41nHJAJEKHFWLhRXbJnW+NGhqu1Z+OgtAl9M
z+EmisVHRnyLuHUMg11KAjSY0Xwc7l1tvFQEW0ocN1YunpTFctff2bYuIBCylKzj
YgBkfBhEqXUzM00ephhaE6djqvehWwVHu7QYPaaT6Bwy4JDrEKVnQCHS6305zydS
5PczZFkWHPiD+En3jV6+Bl5vWo/d9RzheiFtzxPH/LcOqSHSEzwwN62DYGAhJEgr
fTbb8x+O19/VRLQMlP0h3G7sLN6HU3a2Le1uf1UCYSN8omLFx/yD8FSSxGEdxm5N
axh/dBONCUebiA60ZfM+dpC+qB65u6Q0+pxfMmiRsOxSl7B5IAxjhmdbj6NmThMF
DwVQL2MX7OGSlMywOKvpSXPdSOWAd30wwMfjVqWU2eRyxUwaeN1GfJc05n4KDMBl
NuEAGEHx0xQqcI0EEaFdHwr8Z8I+PzIS4OMesDD9km6iXqvJaDK7VO4T0g2JR1nK
hTPqyG+grEqzo1m2kui8Tc2/a5/SZKQQnatRO9PhFek5D7JXv8SNqX8pqodJBF5l
/Lu1EwkYp+2LQQozPWOos+OqWGRHoQb4Tzs070dAolA1uNdOqYI7p0KHh8580Kb9
yprFUXzMf+691VnMoSoeF7QqRIMikWfMQ0gMLQ0f3yPgAQoxM2+9Fapw4DiWo9Yq
CSl6bIZP6TuW51HdXT2NM5Ck2+0bHDJH9KJhJGENhVwMkeZHc2GSMq1Lal8PRXrP
dYK6R3a8mtwx4SxxxWQmQjNtXD1XEjBWJulW0BZ1OIF5cZ1OTP1OqnnYZdbqLN50
Ine9f804G8FcAXBODqwmNhR+gj6y4pcCqfwG3XEJzeukfBhxtELjMrFVbmEcx/k+
EMXzGcqE22R9qnF1Wav+qBKRbBLI4vrJMzzFJhHc6i13piuj+vmIK6G5oaVpsmUC
5jtLmpC1lO/GWWN2LXbvb++pG5h1uy5uVHS0atMgIIFdKvbQNKNTGyJO8DKcUXki
nI4XuSNRi8aNybwvuJUME7eC4sD/P+o+UY+AyHHtBy76ZSMm1KJ99f4VjKgObeMH
P+lam1OiLrGkRNaS4X9q9/MXDiovYva+iLBk5uF7sNDHWk1Lz5uzt/G+6sPEqzny
YAvacKdpPnUW9rOoNEzEGnlSYFb741QN951rfbNVrQmVxwPZFvkfW+cUF+PSW1Dn
YJIAHuNaMVYD/8S9S7DcJs68hEppx2MTOPo9PSdi8a50ZItlgwUJZb9toE4ccXLZ
j4TEl/CnklGly+V7WmA9Vxr1yyWbqhMMxtWiYvrD/Lh3fmNc3vDJ7tRkBJGPEn/Y
iWQiWQ+Qv7ezFzzGIkfCRfQKVy0q0jUDwLWgjVXpep1Q8Zv9RIZW2LkzvKy5c3Zz
iZKnVCEE2Lo4JoIeUv4k5jOY3JoRwg+ISsE58m/c7clIplt3X+a08MADjm2mF+NG
1efMBtyInFkScTCOsOSo9JOz++gIscuEw0licfbE1qNB5yiwrzfu5KMMAB0/cVAl
Faky/GgOu8GfyPiCQvZy1RAnkdC8ZRjSqHrYTAtSRcxuQBcTAXXFb31eBdTtyexN
XNY8g05BVDC6iWAComYFZSbop74d8TiFkZVQYOQwQcEWCC9a4V3JEJxVrzc5t/ZC
674fE1OxXX5zYMy02MCsfxGKT3kOmXNwAuMEp3tMa26igcf80oipDqLMjd831rUC
KOmKMG4ka6P7Wi0SsqeXr0MeYg7SmbyJVgbVfrkdgblnuSuFBu3rw5qB0qe2qk6C
Qc7KVmZnbEnXYbbIEA9VIxtA4YdEx+SGYKpuRt1j3/qxtoqRE5aATWotLwS8BGeN
cfH+6fTyt82ZxMmdlZg92yTMghUbk2eS1WMlJkWt67pdRshqC7m/lfFzgYd/hiRl
GTAyJdBeJSeekAC+o2EvP9WNny9PGc6mb30l8mrreVQKTR4hITmb3gmQO5n2ENoT
q432bzKDbOVSG5rdWg23Z5UJcivXPVl44gq+9/k/mr5Tuf0AbOcf73AMzmG1dbFV
VN0qpby6YEE2enZqQDqIWsWs7YZvaUhHGI6xrxZD9Fu9xDn85ErDZOeIJr8V5g0P
NkdB5cNbbmFb/CuQxVF4WRsXFPPHdEshu6K768cQKPV3AWQJf4K23A5khF7TNXxe
2qd6I0mKgKSAFWcB6+r5pP24A4kW00Q1z8UmDWrorK4An6q7RX22+akIn+cco+nn
tUciPy1sWzme4dAjVw3ic0o2/L86B+MsNM74p5F5QXihGU2zMziYf2bZ7wd3yztv
ckJZLkK35/0O/18BGR35Ja2R4JE/c+MxBVRG/mPOT/0nkxNTG5kYi4CrqOQ3xZEu
I1Ymsm+clmYJXLPfNVk+tNqgQSsV2kKy+JHM06Q9ko5wZIUXJRwqbolw/SkMO4BN
rbMrACyN//zVXplIfzNMVgg6NWL+jqZHgyeA17pR60AA10I+8Hmw/AgpaaCvfxMr
LOw7pn24J+x7+gIcQsU1/4sLuF9tDPJyoZIczs0G427j4zgqusfw9VHt+emtSRvq
DKnZnn8jKAhFmEX4Eiml4IJJO/k+tbZQvRzjolHwClndY2PbFoM0N3FOpY4sLBs/
AE47wERHR1on0UNw80/LDLejzYrbEXknilmaIaUWvUkN9AkM4yYX6IHRYIoA0QOK
DixJpA4UXzO5Cd2mas2pdED7PzSGcuV6/R0kfjHhy8gaUCqOwGtow15kCrmDLwpc
7e9AfPk4AR7laocZpKQ73kTlsy2Wtcteo9AAKaLcyu70A/IVc8+GTzZ7HkcPNOY3
6+Oxp1JnNntwdg73wyzHpKZJv6Ke09SRSAo9UbRlcKn2mzAoqL06tD3EJtBKkPpo
ru2UTLWFxoLucRKk+s6qSUkpGcZoqu0BjCeau3cwsN/OR1ljZdbBXbxBu+g0ruNm
9WnqiqcDGgylQdOBChfr2ZFTkrRMvxsjULanj/65bd1+i3HOs8MlZ/TUUEZkpN/u
JL4PZZ/2ZX3yZ8Wk4S+ISnYx+1hIB2y4nSJlQEeV4c4mJfNzTupTwazX+rnWKPmg
NYqXvIMoN/J5ycyD9/4f3NEwqy/FdwyY4RRNCiV3bwzeVv9l1mYlSXDUb6F4wgyN
ioiQRumwsG6u9qzcLllRTU2pOir2JS/KSMKjH2wXvuEKXAsCDOg1u9VciEJlYFNu
d+rAykoVmo4o/qUI+BU665HDSl6sq3i/tiQ7nJLNRnTl359MEL1syIk3sAmxcw4I
DcJ/JJGuBACx3mY0Pu4+wAsiGfDPERsXusndWZ1BvkmqkDdfKQQsqrYYOYZxhMaV
0Aimhq+LFBZN4ciXhnnErKOFTLswFkW5IX5dTU+RJ6Hj5pzVNeS1m262O1du0HOU
ePVa4R2Iw5dlEL/HajvMH9hLHJ02GnrGLQKHa1K/svvGQ85ms5XLJlALPJzTeTXg
ZJAWgDVryQCQSCUFiK9wqxz3oRb8iSgnDaibVOL6ZfarkTiIpEoHFxRB2qYQQEaM
jQvCHW2D8qqg5m+tVfSVt9wE3CM1QJmCm144AeMrk+n8d5IppYyNekeNuGEU6mll
doRpenDf+0O58uB71Z6hTwhB6pXq3RrUR39hkIo9OT+RqSXnZHbtqe74LcQU/bXv
WZtlegw/OxecgItYp1VqdwmVeXXBhd6ulRntIrtaZP8C9eDMvdGcie35OJEXU0d7
pDCPg4yZ7QDMliRCEG6D4z/+0VyT0m/XWBRMLfsVa76TeEdLSKGXOgCRepJuWSAb
vcfz+zN03rZXuzTiUdZBnCjmQanyp7sZxEw8PFDPqmC3G+VYNyMoSwMLwwJZd9+J
KLP+j8DkkLFlk0F4BeAb8vFN2OccCGesipE/BldM1YDIghjsGIWuZzc2K3Id9YT+
7ItskCskxHnneuXjQDaZ2pP3ZtfgyUkNZ/sGvi6jwP3F4wDeH6wPZkD6asqwu1x6
njywZova9Aqa/d+xaRJCAmZzxzv1MrWWoBHnp5n75a+GfblYrrKzbulMHSlj6/hI
dnKLTB94w/4IkFKCTcEqAP4BIaNm0ep3yz+mFiLT0ILtS1s5Xo6aUuWc5kJe5BeU
zgeM2k2DRLR6aMcwYsJ5nr07Uv+IoXsOW7xgbldaaxuUWH6nuBPglJlTUVNv0DAD
ZfBlf7mCYt0WxiSP5eZF6MPln4fU2XCMO51CvAbCzSM3T2s59HUxBvxATXJrPvZy
`pragma protect end_protected

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
dPM+lcHcz4eXaXhbCCBi9OGRGatSJe9zyupRuRd3VHEcvfCGH9jOWBOLzFuQRwDl
6KCawjwaMz42biGpBUEmsa9gO6RyoNiTXKGSh7uGBw6a+Av7FDm43AVFjow+040R
ud8Db5sii0xlIxXGsj9ms6ws6MjMv0b4GDluN1hljYQ=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 6000), data_block
r9D2Hene2cJHV/vHJWEdwmwout5upvEhs7OF6kq1KXq1Vy55w2T8vfSTyIh+nS3a
zvU785oGcZSXALKafmN9cfhSm2tmayi6BVBhTF0yFWPBv9Avxmt5yjP9lQramzEs
DC2ZjT0xMROYPaPUqx3nV8rtr8ZA1Qp870QC/4P+PZoBRAUSVGuQG3ANpCM12iJj
aXFQRH/6Oclqt4J4p8tuObnekneRHY/Pwl0D6M8qYHtDO9v+lWJLD/pJGtBNeaGX
iSaarXxyOdFStI7e3aru30lupemYxDRjzYQUWE99onQT9s/Y+lQU2s6oDrzdNp03
eFZtZ2ZHsTgFVdzbKTPdcMPE6YZvtLtiscZnRafGVg+SXnaEECQu7I1+Dn1BzV6i
hNMkGnB1cxj97MczKIwRoV3QvJ+rDSPuxUsf84svDXu+aepkBkxf9Era8idu65kq
yLsgv2/czAq5yW2Eyn46Wu5tZ6RKlT5XBt8j+mCxtSjkVnqEnvaw1mnEJ4g8Bb1w
dC44JhHettXnCsIvl0Olmbz1sdnZiEDbKkiONKiFiLlFAJxMKWPSDY1b9vQkTWGX
3Q+4Wh2fIJTy908q5g66aJrSIXdR+BQJzKS50U/k0S5wOwNSivp19LRQD5mlQ46g
Ph9ZIJYbbJz0DKhO4UF0w0kJInEZlGJVrGjFou9q29GBE9BSInFf5p3kFZFgU7qf
hm9lOUOXIqV4hw5lxI3La4tINOLABs84Pm8Hk0nJQcnOxfGf1HOJVnpE3SyHUVvh
mbLrNpa+T5TevKxY3/WBHE70jXO/INywaKcYOwQKMI8ON04lagpPbltEuWYox/+f
bvGePa7Y98/9V7dxjCNnyDFIXWwRjBZBGhGW71TKWIH1ZM0hC6HEhN7PZ5DkK6/c
Lt+UeHimrrpZA/KQYJgFNmLMyvHZ3XxUfkgtER0F1rZ+oRR/KzxHcNN5KB6ncDbQ
Aqm/eRUOkaJ8YJ79o6WjDgKyi2t6i32vGsToA5qjbnfyY5QxKxPH/eVG53LwGdei
Zdx2Elq8kN+RMF1XuBt4C9cAMF0afV84imuNqurk2j0Qh8o4mQsLJGZTa1tjgF3h
ZR/kgoOPrjw9/UI/LzvGrdzit1hSpsxnms25lkj1AX9Riv3blVbUZVFYtxMT7Sy2
XUHMTlSGUYs5Cn1ida3GiQxNiTNXLv9MdUMrmsck6x+0FphuQxA3jXfbochW5ShJ
sbVtjX/vyb3/A5akW1J+47GgPQ15VhyErL62bwEl/zQOMQ5kXJmq/lXxwKz9SkNG
QI4hgYpV3irphN5Rl0yAlguQVC+OYdL7X115BKrV7BDEWvGLnovnK4ezo+WYsii/
84MclPMYWTlFHY/l25QA6fmVhmApBJGWL8spu/qmc6iX0yV+xZYUdcjokTnyZm5B
UVkD8WPwckk8J0D+2SwySz605oS9sYnvGrjCzg7qvoijy0OGdy9hVfjbNehdtcCN
yOzzi49+PrPPF4UA45k5v0DbToEc4tPfjAk9NgHse/T3wnxESmsDaXFRBeEFSSSG
Cn1BIYCP0/3PZnTWMC9AExHZbOrMrbpkXH2iQZ/Cjnp8QCdCcpYRIpVmBv2k48b9
8ej+LBtGfyV+ziz8RT5+j/QugUZndlU+ORAAWwGePU6tDSbmqRv7uu8UFEY5mJcQ
elYWLvWxmSgf9YqkR6cS1t6uMyZsbwOYpEV7FbOtgSJs/3aZ8CQQ8gRzibhNNcq7
CAKFCtff6ujbB+2Yicsbl770rbB0kPYz58PYPuqEjyXD4IxIzreSaKs6rDaeGLQr
jCmsHfU1Wv2eUngMiSeleLTY814ccreLR+P82ff+t+JKAuzUI5RvZzk67jhCI40b
u8RpHJDcvgS5TD9wZgpDfoPB3lo1jLGV0XNPQLOJfMLtbXUw0vU2Tg3GO00RxrwO
pnLxFjwf47Hl9wpMOf4l/nONVQwQ35owoJ+KOxCisJ22jemMZ1DCTS3JT+lJcJIL
5sb0V4Hulb+fb9Jcannj8fS/Iiwb5r+6Le8C2GaSRs63n3++TaryjTtpMSDIiINN
S3WKoL0N4pJT/VOpKyBwJh1ZYEvfdgjpS24FyewjwmIlnGS6L9klugdc2H+8U3YL
FJ9NoNq0k2EZbwyzAKAneV1hYA+MOz7OYtJN6QxWmU1fxDCNJUPo79fIiXxdsYhD
AMNEKJ0cNb/YcJ3xcZeLJPKFiVDt7SLQyDxqLrR1sO8/0JuLsUxxxZOMQfYPvWJf
NtdauiYNr8+dusah/gUFrUyG6saOB2dMZ0vgZkwyWl0yfBte+Avecpg6IX3O+zDa
lWBe31Fb3F9nqMjOSbzg6T2+IVeXz0L/5Z0Bgk4agrGr6PuizdV/kD0jpt3uRGOj
kRtVVkM5CUjG54RQtYV78DdJ5kUpxINFGpylcG7CtA1e+ZctfqKXH0rHmvnPkEh2
4Ow/asj8u6FD7GaZcnSt7XB2lmFbawn1aJ48UB5gm2ioJHfipLQt4nggLLxS1NjG
V53W2YwqdwzniPY8p9ned7VpoYMjejINAc5SwZBak1IbRfMEisK4+er7E4NtrKZZ
9EPraWkgJnmt7pEY0t1Z4097IMhtPhgLKL9LYjS0Gk4ZXES0NJ1Vay8jUxVumU2R
miSgCKNmPUiokuTVZZ/GLtLpkdEaDJ9OMypTisqoIdJQRwrFv6fHpt3RsBm2nOcp
/Nv24BVTryK8jG/OUtIXpKHsLe6r0dkKK+XGU0zhjJfIbXbM7MRgba05NYnkmxyM
y2gu2TarBgFM6LSpkQV4FFGfioLBXTbOP8UBKEOsYLBOOox+ljFBXF+PNvLUGVDm
o+Q9MXyQWd9iEPIFqDiJPOiYGJAfyZ6Yw5cyEaMU4BmhApvAo4qgS6pMB9XPU7lS
qwbEG4khr7voQPeopJVx9WBe2T5hy2w4oQjAUAlBR7FDsniNYYtmXt8QGIzkd+fZ
hxBGr751ILSkuQ6AfPAAI+0Ib0anl04FZ8kpPQf3/JHE+KO5QjTpu6d5Ad/RAqhX
gbwyWFfPv7GXhwEOo8QTcBkxzGJ5vVzIxullFNMXOe+HVyofQKXUqvXsKLi8nZnU
AIa64S4EKxeO9FJ/DfzlLR0PsM+xOnX7RIDCcCp6VPFY1g7z2kXYv4WYNt4C/SnB
SACQCZ+RqTqXxNrfDPcA2hjEJBZOgsEGjGwXU0LLmlV4W474FXpw7nDaW3e3soZf
vyBXYxkOt7EC9PzMB+aNWwK8FkHrndTFpcDSN3hOO6pxDhnS2fFAPNIAoADJO+H5
2K3g6B7CGINZ5mVDhHKENCkq7Tzt5aIjFWHHWOQOcQe/cl0zw+4hFG+pBiIIBpPH
Hhl3p3COIjucChRe71ACJnvKU+mLEZRK4mxR9tH64Bfw0L2tP66TRCDPqPdN+6xb
ftch1w/sGQXJL0WoOyqyhLQ1HKbf3zLfC5DxA5L6LI/ONM2fxE4m9I8qM8BaBcN0
OXV4VDNBtHg8i3QfqdrJe3qF95RYK8BL3Ap3e8BR9vumhfuivcgghKxSgK5q89Xr
Lq6X8fkRwVbAJ8Ku/tuJb2pZ+YswvMgMwaXHEXfvYNLg4nQKlsLV88v4rodGbyBu
FIHtA7r9MLDQ6Unyb28XnWkD2BMkTjduGGnF+lIv859lhUF0X3fTIgV7U5A8VZp0
Nk5EuZsSJ0yxfLUCxrBvrWY70TTYxo7kWP2DUC7u00gs/tHvw6ajxAM3n+nuBINk
GRsiiotUINPsjI3fqR7RDevfQV9K95MJbpygcPQrXxziDFmRDj8ehMxJ4PNd51LC
18mecMEXtX4bvXEftEE48sP/sVFYqMPTa+q/Y+o/CPCMY44MVt9FQxy1ORcFB6t3
GzsyELy9w75p3DxeVom7/jHO2+XS2dfZYV8/uLlmCjU+vl64ATKcjnoQ/hiiIKyp
1DpKD6GvfFXWuKIa3VEh4bGtO6FFerBrPgfmMn6N8FBQyrn3F7qIixVPa2X/tLph
U0wR7GMufIXbVX5T9RhyYnsoL1yioFkjyRJcYsN3VkD+LdajWBciEaPVLMibov+6
4XwtE/VGuYfaqh1+F4Xpsmo9HTBe77QqbLZDSS6PAh7Yg6LwQgv8n7uOF+UimACs
a0XfWRNbwYti9b3TqHuV2j+auNsEo0R5xuzE+Faxuu6BzB1mbYHz62OCMWLkdRyZ
h0mil0cjgYKd3E7Si/wjBsJLAV4joMfB5hvh2Zdnxb0OrPKhfEgvm09L3EIeQmRN
aarD0qnDEJzsZflLR6eJ5TV9hvdqo2OH/OgSfuFjqdv1QalERNQmThVYOUyDB+2m
bI6O4yX5SjY0xZtFct20PE7wpePYrneGwszjUTtrEG4EpVTO+mIfIl+u5jsohVQs
X5PbQPjJci4wkvCAXKTVz5JsSAgUC0UZrkNJawEDlarhG3E0spG8UjmfSlnNokVE
cZwFAYC+ZwhGjAe0gQV6IpTfG6QTrGlMBDptm7dNiXdriHFg3++JKFXrHsMMZhBe
DGXuCWiCgaL9eTjkgH5ji+ndhqa/dTeZ6lIWsl35pciK2v6/omxChCyA2h2LyjLs
ozJ865TBGibiteFK7v363s7j7cJ51NxtEwdmN4fYhUDiakX5FPZb3cHmLgdpyw14
SGKEezd7gsCnTH8BHUY6CuJQ0Fv157IhlCj4ETh78MNhtBhsVGZ9slam5kvcOuJb
0rPoIohELqrG1x5C9IvUMvnPLltMhn7cPYBCARO6H4kdoageQ25/rlMFI3Zt+5K6
MenHlWtgLPyD6aVGwtarmCDj1LdBiiGgFy81M9qAdyr24N50fOw81Xrn1aN+KZc5
9ZTG1jYlUyA6vGfh2QVLrcSIruIIvIMhHuSVXRGlmNr9/DtFOvz3p2IcNqZwraHB
FJtuSg///zrH3ni9XhvazHwCV56YMAQRLmLm4E1hE+2V+ya0ZT/rSU8BPWCD/w85
bOlPZTEb+KzIWj3GcpCC6WWxnIcEi+2mWfDfDmuirCnV0P/E8d6uH4nFKd6B88Li
sJD33zmT57ZliH6d5NhhT52O52cMkZ3uiIroDrnbe/Io5INqx1s+IK+xNa6o+3m3
sViVsyuO5mtb3eAwJbKHpgzSBdc66QqY18kNJ/KfPEzd3hRVo57MPdv6Owv5evKO
GyYoiOKG+nhQbMl6VVV45eM6n7bcSzcNfPv0EgC1QMtHBZ3+NqI/DZ4isFrkH39e
I0jcun6TDKGmm14aiDVe5aG4480cpYyRd0c6LIf2LvJq0Bhr/MLv+FMuONIs2L2A
tXQqiDdGQMFR5qX8dp4dIgXcvaelURzhqJh+s2naSSlNBj3OuXB255Md5bwoCBiK
iTkcgx02BExEX+7N3ft16HYA+w9Eq0w2fg4kC+NRReH3bKM3wJavSotcnAEoSsG0
3M+MlZt+f6JQXykndExydGTjO73DhjDDcxZcg2JD31zI+CBYJ8X43jLLlEyoJ9iO
71NA3S1B6qXe4aIfd6bLNOJQXt7CMaHr3/Ngdi5yirfFpTNyWfUdgoED7JTgrqKl
ry+iLz6p9RC91xP3nONiSqUX1kTjAKY7jsJs7gockl3ZFWCVLWBP6sgdCoU0M7Kl
NfS3HuxEoRq4z31ZJYpLBeAUt9W8j5cht+66hAqJjG/ndq50n47vzS1Wub6GELew
qD35TfVX43AwNirwsgwvEF/3VzTyHTYGSgFgWRAvtoCJCaJ/OLuOlQnZl6HlBbfs
AO8HJEKbaKaR/PbS8fOU7wypjknqUCcsFqE8vflyf9tfXXVWvC770SiQbBdnZ1Ov
iuPkHD7Etyk1xUM8w9Lk5YwEKtaVJE6ZT6NqJK0dRBjd1r5oCqcjxJ0OVzFOrrVR
BoUT5uPJgisaVc7qh15lh8K1SyCpS6SOFMFgJ8FHzsvYpwZ7btMR5fa94adHvh9W
CIwoxwwngcZ+QEbj5DLUJqnp3xelbRtCvg21xXqm5yK6NiXdqKOabF/hdL8tgD0U
OqgzIsQajhv7rytL1UkUZcO3Fjpcdg3WGfCjZE/9zThyDwVya3cO12Qjduse/k7Q
D5KYmqX+gaAdW3iSNoEaFeLFWpKRAkYfyRTGgSwEBVIbLgw29lyaCAtUgFTxmctD
uBM8+BtLWKA5g2Wv8cPpvAYbBOhq2+niVZeD0FLaq0MEJLr23GpV1PNqLfC/M5f1
ek591fG2Kw6WF4RWa1UHaP72fW/nC2+cMqsTchttmoVOJrEHvmN9mHFIokvEdHdy
MB0aPaBPDFudUWEtTM4QCkZM0+J/MPTxo+fUYKM8kXEbrRk9wHgcWS4yA2rtgQ5R
E0NXgnZRdXAXpLpFPnamXBCzVwTLIq0FoqZguG68yXiXT2W4tH2Z1rcd1dcgHYZR
5QRSCw0PE1QYGaW+NFZIfHlbCwoF+RdCCfajvyx/0HaoTJJ/ifbQFTP0/6x+Mo6f
H7Z4Rf/grdRVi2NhGZduNaUa4yMflPaglBfUEP6UhohOV21DhFD6Q6llGqNU/xhQ
JE1zi8nNv8tXOTCWsKgP97kwdf7cECEFbxbwwzRTGwYQuofohmVxMhAV3EptNSID
m39tOOF7JRonfMS5f+m5NGcb9frK/TwvjaC6tbDTqagoilxJ6BMwMdjdqywYBMti
AYSQQtAJCZuomcryqeN0sdpLFxDJ6HqIE1XsH8zl8S1E5OPtZxHl7yKJOc4AnVAV
D6sCBWEZDHa1XUP8OyIUKtxsDeJgl3yoOhRvqvP+fFu4mB6e1DHNoFTGm8yFPiT/
Q4WufpMWcXgWTAWIHqnnp2s9YYlF1unQ1ppBxTCtALNifPDbmcvJj2q5s4WuRqqj
U6bEAFHtJpiaaXPqLdquphwu9hAtugg0VUhM9JBjg+tAgeP+J0zN2HWrmLTBFA0R
WRm74AnFtAzqu0wJKmngxPMTdVyAnKh/bcujxEXu3tMx2vknWqP9hAtB3QLw3g52
IT/A5Fm8N497Gp9aD0QBJoxvqNh1BNjbdI3sfVe+54OXgh0l8wKPIlKjnTEVuw2m
DyhReBP9OGNLkqLqCEXBCR65ItTWn0rOpWzDCYOnmL7AP6OB4Je4YSTJ9qE6jVpH
4P7BuYpyNAgkzKswTFiNK4M3DbJXKkqt+T0gpCAaZ2rdqZGwSJFFqFTjMqBm3+ft
7/I6Md/Ut2i3n2kFid4rQlkxSSH56tcqvsv3EOmi43PLmeLAPKmfOx6mSeAONGzt
YXdwhpo9rRPGXsCCTUtviDI0Q/vKfs2eI2iSAQxGl1q4dj6pB8ntzD1OlZEzszBG
AvhhHVJj+YT23KPS8kdQX1ZiJuopO6aVNNLeeIIUciNVtQNpKZGG6iiYAxS8tTr5
gRJX1FvNm2iIHnHd70u/KSVgWaJI4O8RvxYmEgkZMkfcwsoXcmu4EfpFNWPWHDy+
9+wtICYM7/me0X20vQvBs0RpaY+Pxsa6zog8Hh3/XEnebmFdhaR5QJwXWmhXGexX
n6vBYT4mvLfADQ38QUG84qOzviJga35HflKB+1VB3EX8wKxFmstd8b8A/oXLildu
aA5thsqGpTE0qULPOBodnhdJD8Mqvv5U+z7L63iZG6kRmh09R3gzY66RGJxbm9Sf
IFuOfpxhAAhZ8rP8pdSlEP/PpxPfVN6PxmLTZ1U3xOr79TICPgVJM4CofUb7G+hL
kT0nTIZphUy08vhyAdUSj+pWhz6spGvYfAIxi8pI0nNhQhB5jP2qg/zYczrsOy3c
WXPTG/nHNwKGHjP6eTVR4kpg2l+7x+N1Eo16Y9VRKKZL1+A4Gt/qhjTKY+e21i9Y
PaScVz1rDYDQ4YQysidi1DmlVVy+pZUQg4qmIRw7LCUlLGiOuOrfKWQw1APgTGR0
EuhmkO4ReY0Cps9n/G3Dk7NyHUPMmUoqhIunLXTsb40sqTPkuClT9pmWeuSvKl5+
DvOGkwIc6fl6Mc4UMeX/wraj4ZYcmnAL0haeJ4RNMXTJFVgsvFwovrV0AiGWorv2
WqA4IdwGRe0lOGxb+MvT2yzoY7Ylrr3An1B8H8lWsCXfcJIxoAXhaWj4YQjulsp2
`pragma protect end_protected

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
iNCjmrSIWTN8ZJ3a6Ivt13dexNsHc8MEEQPSg8xcTQAQYgXYGI5/4ppkUhErC4JM
iAs9vYkFNosz7QeNHxlAXOeRpt9/5lqwBe0vZGwmr7nD4/gqBKTEkiK/YtDjz75O
cHpFIZskBHkMx5LIZ21LZNlQBZGqU25xETtIFPJlkcw=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 71888), data_block
EEVwOLtWvcYcvHZc0q6Yx5H8i9hjmWC+a57KJDDwTJ9NXwOM1+hN7uIvTEzWDhnw
LIZeoZqoe14LyZiRMmIhtB+Rs4vKtyp8CDa7eTIMya60lK8yhbYZF18et0cBRC38
wk5y4jsIAkOVgNdvn2b+cROovy8zfdexuFgYeObaAhl1NB0mGbE4sECDV351w+Aw
xtpN3CZR24s6h2L7+PQjRkSUipPvxn1LyBlo1rVvKMkYiNLs1tg6sPHHZW78pkmR
KUVKtbSHC9mPxSVf+3Itwl+R+pIlPlXSPKxFgo1ufw+1hJJzJ/h5yKUnPYLnxRol
3a7gN+F3EKSxgI5HzCMRO+CQ+HbcdeV/EOQfEBZv/6AT63ujMx8TRA2ilGEMAIZ0
e+d6mvKs9O1aXjRuVTc7eeXaEd4V229U0hjtUuuWcC5kBWIu971cG9k/YZlIxVfG
X4QJp0zkGvyZGndGmOYg39OlHqC/LD0el2NYHFh0EHR2aJonibKOCZkjW5f56d3s
zgtHm36I0XSztTvv3OZyGrnf4ytw8eW2SyeD7Nje4EAoj0g5OOGFTQx/Z/5XgNVs
HX8Xt6x4l960eC/fpAm5EhzXiR4OG03bmkZpityQEyGJVDrk3j3AOaLJTArfZvCS
QJm8t/kOKlmbuNlehT/VGqLZK//IC7rmWccEYlYHRQtPZIZabs5WO1Z1rRZObOBM
bEFYQN0kpzgTD2/JmVAYbo/0NCpKqUCJXFyHMqLxTwRY2J6a4r7an0XNYXNUkUOp
Rimlvpzl7YjYYcNmCB6xEQRJ/GvxFmpnpd4x0osFYIZZmuX91aIaFrF/E7HNLnVR
S4g7xUTle+EJkdKrpmW45awTyiVvdrH2rVu4hJs2hGJKuBldIfGdwT6ZBNSV/FbC
QtvUF8JmulU2/xybnBHrkQiapgJivzIb2oIhAG5RQcNtcXHTCJrzW000DpgfTflQ
Q9Xq3aWjuLI517TNRa8JmOLWDZVAlptkcUDl13gbMOCC7UMmLcogSWEyUA7LA68q
uJ/6kjaxN1batN8xp+ePIfvoEcUmmk44INg7A4M99PFOa6muVC7BAGHlDqxD3oqy
2YxSc0Y4TOeVX3Sh5KPMYXWfzESsq/7g6UIyYMqUpigVD0v1YZ8devnKP39UOLWW
8fY4arqT011qwGiaHVA9krMHmz2G5Q95tVMzeLERpG0gJfKiN7GlZ/Ubd+MVyYDB
KgwldqkngeHBiv1h8dXtDZZTT/uiOadB3UszcDkJCOb+0NecvteOzTlzKko3EvLS
IgaI1vZh1fNP0bW5vhk0kFv+HTydse+8UUOD/apYF9JBgxsg+Rhn01Q6AMLzsihW
IVlS7uxHv+OExWe/sqH53p68mY9oNI75TAdF6Bx0XaFsbW54I3kgPN3AYC1zSgLR
dig/g+oMh3ERYIo5Waut1z+o3fTAeDzvcY1HAauzPV8NeaNO45JsSJu9eN3phQ8B
EnXMt4ljvDi2/hTZPmFWznBh9K/93kttdQrUTeglvgzUB+04JVz/NClP11oKOQLu
XIZ3sJmo4oX3jyIRiEp6kntCN1Iw/GINMBzY0AssjpISrvn69pARRew8LgAmXlF+
vP2TopOtXpmixFqh4WNntFuDneebNGIFXkuAAghjLxuKTdFpkPlXSnPb2X5Pm9em
chiPSkyfolcGegD9jcid9oI0lVQvR8AHhDJ3cZFYPAjlLbnvD7Fr779Y2nWni/4H
74mR88uBVRjneimJcfMDjVyJUaSfNdkTq5CC+eT1YcrAx+xlzAx7quyFHIu5Si6x
SCBuGrXbV+JAEUwIwia6iW8Sc1UP1iK47UK54U9yzvDvecKJ66Nrst1+YrXoTQEg
BZFCVD+A8hs1giAi7iHiNCBcrrTYv9lfIZ5nFdy+zvnq9sjvedPhXMZoXGMlIz6B
igiAtnnfiR/jtBnbOgEF4CnfRa3z/cWk489XQd3MKw+f6WX1Wra9ICeQVS9C3sTy
Jy0Ckmd3eVJt+n+5PUSCQv2SvyWi/fGFvokGR2dBpdB21KWepJbpdqUTaYz9QVkD
u5Ks90ARU5SSkUjJEvfddz/DYNNZJYBiMfU0lZZMrmDuVyEFCn1Wkr2H/tTIUr7Y
1dxmpnSs3KSKmjWqgeY/zHWxM83r+LlymYI/c98fNXumNb0TwBifKqkBuPDlbVgI
c3EpuIfzttKP5NNkfUCK6IFz3w1k3n7AXMXPYplxOJxqi8PYffsUdtdauTZbkHPH
c6Lr6ddFjWLVp6jyYBA22OcT9QWMplxGIwS/dQw3nKjiCLFgSh6RlIC20Luxgn5h
0zr7+Ozs/XLqFmyv9krwnK3p1PhPyBQPcpF/Xz/BZSgN9/KyYh6aCoAmq3YMBL/F
tzgXkzWG8W39xruqEBz5eeYmT4c12pNJGPKABNBCuw87OkDzp9XYAgp0yH3vOhY+
hoM2HRSX9Q5nDSX/c/m6/lMbul69BPBFNa26Uy36IlS465fGocnpaNBSjzBqHFbx
E/ncy4LWFfZw30kYPCz6GyHLXUnvO+u3E1VzTgoHVgd1LntFGDUlzOOfeSIY8b0N
7Z4M2K5NLycgxu31JcZVw8YbvWEX3Zs42NcuhtMjdpk0vPa5mM/OI/Rn8yA/ca2d
w24jDkYkQGsWAyhLEIb28g56OXIOIENY54Pq4BdArNWzBgRKNv/PVS+ymsqjahd+
0GcnYHmTOCaz4/fca1Uw8XHZbnXbyYnWMJX7ve+03V2Q2gutMwqHiNTGCqJBMxyh
eXstrbrTH1UY5Q0H7D8Qdow/SV5qTlAi7x5D00FpYKGVC4zUWe/I9tBbv6n9uYml
uSbFWLgEuAr0YKearj1GrF+y9y8ogY3OqzcYAchvFRk1ijau6z0akbCut6FK2jbM
eBohPH4L08T5UxwArDVmgU0fWSO3Xqxpm86P1PD7RZv/oDCBIeQ0mtyRVAgqfA2k
oLPa1F9ImSAawvPhNIGPwN7OwWKrvffXklOL01F2+31bU9tyFpeeB/fXMCZQty6M
AldWy3UxiXSBQNzuuovmRrW0+fMQi7bdmGK51ZHFwtrQZId0LNkOriSvykWDi3n0
JzSJSDQHgdReEphBJjDkfC1AqRpaYPBi1hThRhHj+pluzpev0bOPownExDbfMtym
1NT/o59hi/dGPZxRidMMA++uEVW92hhrklQ91ZSQo47mLIFyGk38GQNppp76QBFN
nwTw+6nciPyMqFqebwV8/t+mzsyxWmrnPUR3UTMcT40Du1H/vLDQQTYDtAc+ohPo
+uVNI7Wdy6e58GZrI9qxMwW8B4sNKbKnQ62mhSmoCUEbo+haZFEMNpjaTQ2HQgH8
fsEi4W8khJy/BvKyRGyEF3iSPu6h/lMwmKmCy3HkEzedfG2covoX3KfmSJyAaKP/
ktgb9FJzoCuzpMQZcq6msP60iF4qIwv5GDhBsQOM2FrBRY61APEng6j8GcK5lrso
54RvyfXTtCoZR1s4N/ZwP0FPPs3otqEpogy0ZaySlDNcXpIeUc1zmXJqPhxMfbTw
s8dHesxnidp0Ii5ElLPYDT4zRZONwudPRk4m2WAGKdwBTXzDIY47VAUDLxYMOVt5
UEzIbdH3//YBziaXt97BpbTWcWeIrU3Qcqk0UA/n8DGcqhF2fmjbmlQb7DtO1up8
QIZSDAoxXTZSAwKPvDCA7oP2rKS2KOfvCrlAgT9R/mmu6Fmc4Dzl5OrgQYmRMTxz
v7CiTObSFDqsBUtRUqmPvReqjHPFykM1n4dxdhf/SSAPKDNHIwn0F/CPGVnj5DG8
l/cWxJJTTO+W+3H+3MmD5gu+RDBbCcn+KY71BbgQ8BiQy727iGKYEmRsf8ww2G+4
Co0A3CK7IARfA/uTtX76n6sp2/bsSNLJs2CLilikbNmHU5gKarGkrR2xxU/oKY6/
9gdXCeB/qVW4vB3pMmG8v6qOiGdf9mSogqhNFWUuHHwY1Hylsnmy3YXwsBPXDLCd
laiDNDYcsFaPdWzopBUiXhUgsb/lkY0kt10hqBuli+w7IWrotJuen3S8X6gMjOc1
ByUgGtc640PEsvq7i6nZ/73560hvmmX+TZviEvWgeZC4TFpuwwLC0wzJHUARmui9
4TMMVeQXgkxD2o01iAPpconnDcibaQg3hUIgrZlIZoW/6SxV4g1KyYxIL9LMgWt3
NqWBvz2c3mY4JrNTj+7hZNwcRiFzNwwjNf1wbld0H3pEEXTHxpZ180x4At5Yirnl
w7aP2lKQyE8VEDBl/7HCLSqSM6Lluq+lnvzf6TqpNeNghVQevDbINLi9x9OlyrKP
HyS7aWpFo/JBHUpSarH46rkJZLT2HQAG9Nf83zRaCQDYZH5c/AgKjDPDq2xiFRzW
9j+/aVbIbHLLMQ8autGjjcxpVIL6jBAUYXnU+isUDYg1GaXJm8ZSOnQge+GISKs4
0vVkDkzJAEcxIkQ0rjtjgMhyou+ZGTsFzjWbSQMQ+dv8OktJ/bycGlbMdPUnsZqJ
u2cMreOv20X7/oiQ7QtwLblJC3UBLxpecCobymqSkWKywuez5ZNP4vIKsAOMDcAj
xAlEi3szZCzrf3NqqIX7GSrb3Ca1L6sBif12JFTZxL1G9CDPUqS7NRYEpbrAbVcC
grqlcmlI0f7Uxu+UH6QhTN24I2NlCkQiWu9MEG1eFSB/oQrK9CTDZkkTsl8RlQqY
bDJQl/3hgabX/y7+nVwfIcXRRIsbvkPfw/Sx2WxVsAol/vBD/riAxxUMfWxYNG4B
O67tqQPHe408PECx3LhAceEbgfcIPTBmc01zM3HRTpChF9/aZBWuJDYgS0FyTx8q
KyUZ9+U+ByuJ8Mu/JAwWlraaATyVIPMxYiw4t9CkKmjW9rpDI0cFMR2fz9aMpgL3
a5Yyrx5hSHTU6uBKClztKdzJeBNkpZLriT0p40g+noB4WisdmeMbmdQ6Z4Z3lW1K
4yFLG1pyN/prxZyakivf6z7KjHf3eBQgW/c0XcipHduZSzHyvZAYLZIUS+NccEF2
HqraSdvWeGdJl2FC5ZGFsk0AXBkKpeoRNmjPbBxftsYh77MkjT5/zVJi7eTTrj22
AZOZ7OAvWqCGnOZF5UrQmeOGXz6YryFbPj1QDD804yV6Nk0siomngS9C6cHgdDmo
jRPvH7LJ6/x6y2EebhvsgkKM3cZhx7ZParahDfaXEZVH6S3VhCiinf/7DIf3DVhm
DalZYMkh2Dn8YfRyoroSpYui7URhb4pzH0Vroo90L8Q6XsX7od0Zzml7Xf8dNZGR
vRxFTZEXPQ+1T7IGUt4R50E/W2uTMstqCcPd7I7b2LdrN9g283UutHC2Nvqkt1Pl
8yQcpMMVz3NYieQGteVjxPR0ojMDdg4BCVh/R5v0NfaKryk1bPs31eSqAcwCiFYf
f16xNWn+oUqkwYjuogU6xMdoPYPLA6dyH5vw+dZuucws3D5xd3ZHa6q/FRbwWMyq
k7ZyCQjqFSIiXn9AwkxKoW/mjEd4oUgtw3vYLGrm2z/44vQtbVha8IuPIftcxKqW
vkUeAC2qRlaQMfs2z72OcyyCP7rqyzlcEXSklJbIiVw/7ZP7l1J+gM1FrYLvhFgr
0HxadEWSkdTGbwkxyObxXvfUbV5T6liJi3iRKvosZ/5BgKZERPLnLPunvjBUo2U9
EQ4PaXYOcYS/EFXyUj07PvEixtNCj3VcTzZc5zbg5okpAiOCK9X18DpWsC0gLjpU
0ZcJ4UtdeW38U7ibj7dgHZAbNWwN7QK+rCtb9w/SEo6WSNddtXuJkQt3YQfV/ifk
L6WkdK6l7L4a3htTiSCw90Oi0iVBW078VIPMIN1M7VNWJ1LwtlTJSJwk9rp8/xkp
BCQ8BUE3Ci/YKx8b4ESMNgNFU26gOVzDcyFnEPsZ01vM/yAzqCp+jIPLtsQdgJBh
T7UT5Ip5nY06OxPXUEy6UVS/FEpvxs2Psqhu0BLMoOW4bODwJLsZkylSYyNXq2tD
t3jhczQpSS+2LNbajx+4ezm+adpBX8wsh6y7cLEDMtMu1IYQSeovWXeq6Fhla+Ge
7CgBhuAVS7EeZmmk9ZSWYJhwUA1DfyOAv0JNp7WtDA5ucvAttyAYQbmT3ZF1+aRH
cF6rJSs+XHTmwOnqN/4aO7lcGN3I5zVg9wnQPboodUSinOBXm5zQoWvPbqTLqgfd
5U+orcEopXGSu5FYex5pMdFXPGC2KCgVfW+xHQF/5zCjeU/rLGZ8eF90YekV7Pi0
rtZqy53+5pYwQDDiLgrDZ+VJ+OBEpLww+GkkFYGnLJOg93YXeX7O4fLZGcE4xANW
AVKd4K0xJuevSUNAGaH/WSX7EcgzlVgCTO8ANJ2jU4WXJXWUVpPw3ZpwmGn/dq6W
3t9KEStqCMa31bgQkny1KlDQo4+7/kYKlXZElBOCEMRrGrIOyUzpGNRSkBtV3YST
12U8dhG+7c4mYBbcGk3YAE8Tdk2jMXzDzncA3K/jH71nLLnw1JOWTDBj8rRy8CUG
9MBfioh3secQjD2w36vHC+ATsx73vhRhiD8svDFstanUZAToDRcjfPNhWZLW/zRN
PDqi5lejGq3eN8A1jij+YfuLf7wgLMIwF4eQxzNZqNtuF0GsoErQZQ/wIKnV6QHa
s8vG3fNzV4K8hBGI7v8p3Yabgiaxg2GPQDKj2rAJssVrvRyHQmDC+LAMC1V+WZCy
Xy3vr8AqciGluv4HsejOBwXT+JAgiuNm+M7z/f8GAkYlSJv7CmJAhphHn1GmMUZi
aebXFj3/KWAS1UtTg59STLmVoJeqt4L92CPCuGXu2Sa5b05d+9P0o9D1dG2377Wo
jqHgmK9AVloI+ewNBPk5oajHpWhvkvk3kUXC/egNu++4u94vOm1MJXFdnKO6Ki7K
B68k0jsH5Cwn4tZO7wHf632Zu33+JebyZJS6NojZmbAfPTK1MQkmqI+Raqwp+teF
ePCKN8txbQ+Ow0Ji1ggc2IR61j1yPtruf/qq874xmeskRprC2A2UbKxOofE8bC56
5h4JxB9Ef0R/rLn3KPHU3PQWIqMYNE2Z1ceIUyI/M05ovOjqTjWvnG3aU5qH3MKG
uij4llu5FSBOlW/519jraek589fJbuV+RRJPxhAPFbUBQhXNhrHWqm9UND+Yes/x
1vWqqJ/ZOxqxGAeamQcwuM/CbGirpnHbvhChZ4/VvURrUzii4zYfJnnqv9jOHdRh
PiAtJLdFmqUimye8I8FQNLZOqEuHwp7tEsgKRHAaiTU00SV5G4JZuz4DQR7vKP7p
/L/WV5w+rlgXmvus6FEqvB71a9Ccz+in9Qp1HvoO4EBAevctonmr4kTlUnIRef8T
mhTEwMLtRnLv7RQgwTiOxiU+yqSg4W+zbYHjsRU8LbfnqrNd1LquTsboe3Cur6s0
tnFhtoQ16gBbn/TJqmO9b9sQ/MmQCNj7uLs0DmYnYSvyqf9FxnqTjA2WZSCvPkDJ
9js/pmT0Bikb3zvGzfaTVaEHSiS+91Vf9neFCUIcWcnG1D20Q8GzdbFGeR71vcR3
0WTmc2EfEaaqVr/nFyE8XI4hno39S0xW3TsOBpTSUqHMouaznhfh+7NVNSbAAlqf
OogX1SN9RShWcL/Gtbp8yBiiQY64orRucLeFINus7n9a0zijcDdppES71fyiNvlo
MgEkQiu9r8Yk67lNYXvLdTbXfVwlcHd+yZc+2unYWynPBhR1meHsrGHdBx/+elSp
RSU2MAmzRC9EQwyNWFDtIy3ijT3+6R9fmI9Tjyknr5PJWgvIwMfum14BkJdyGwna
Q6S5ztIqX71fqTMgwM+RQ5H83V5x/iSuThcu4fD/OmetWsz+OZsKGIZCupvn4tff
z0q+RGyjyPduqV16fhg+DpLJGBLD4oat3kO8w7hgm1wsRnh/Cwb+49vzejD1aVX0
q7gjl5Wj0UNaQq7WgoxF+HV8S3N00Mz0t0Y/cfb2QoBgVBWqeBCXwTAOgUBIQf03
SX49NGgq5fI4KNnOA35xeDajROW6SR6v/E6RgDjKHvx9H4KXOuaHq8rmSpogjOC0
s70aWbdOcJlobVQJC8V19U44Cw178yPc9HFkHhdCKgjsnN5DeQeFj0fe1sZYWpd2
J3kfTUHTzFHNszkdQMy1WJ7CzDaqNgByUaKxkvigM4Pn1CuX4WcPEBZvbs06XCKz
6VGa0jfgeq1e5Fdai6qrGufvn6zgsaNmhaQoYRrlIMlM3NUvNzo7c//DaeAD4rG/
bkWi+7ZwJglxh0qymiDySWS2duiKW/DXOmeEYLp8PA2xu/6f8Y7vgZ2Ser5jgvj0
A9AAA67UFwMj/TWfTb+BINYouwG3hI096HROBBFuyviGBjskeIzfNAwxT/duYQ+1
NCi3iIwA38mRLrgCFbWv5y6YB/8+Vj+0vxUDwB34e9qcQ3jlhsMeuix4GTOgdPSs
oTlL9XflIxMJUNsOVSNUdaw3NhwGFIhmfaAj5tzJOf22+UUwF8RysoaD+LRlZhtZ
ZC5sFGY3hxY9ag/sBQK+tiMC8OiUTsjGYVziihbfFkqhcUDZBwAlg4DKiN9tBBYa
fvDZCDT09vBtNQlY3A1ziIFr7Ju51jaxDIm1BUeCvk+giWVpjWgQA5sgiI9AkM0a
RDPdEgmDvZy4fBcDgJNzRUtPARY0QLYKD1cg2KxXNKrn/BWSx3Zn3iMn1ONOMvPq
Wu3lga9iT4e94LJLfeEwn/l2c3K0t1rnudqSQtEbJj+8obV4KpYLvM+LvHA5qjnM
uK7fhjMJ9yraZgm9fCNk6nYuZCfN3JO3H/lh28QOmrY7kRds7Dn+IB/3J/xEfvt5
OWL39XX5Zmj1IcIq7Mr4u2zkcJYJtfTtYI5NkKErDfCCZsYCmnCBmqxiQoJ7cUUx
ZrwHw6LvQVU3hNUl4hrqYjyBRSQ7+guDMTRX8ePhcW/FCIspK57/+NtwiBCe7oEJ
ZNNPZPHkQQWuP42WOEPZpRyCAykkuSw4QgEHZo8CKUYXaZBAKXZ5VGRiFfOnuDTN
N2YTT95axYLXnRweFs+0O3Y0fYzRNagivk/QxIjrg4HXSDcSXyQOYH7fXc3QM3yH
meQv9Xda+uLFLDX86mpZRn6qtxyUSM+y7oPNIiK99fmZrpycnY4mYQv+amR0XzeF
sjeickNb0jmCY/kGMLDBZkpmwxdxI/fS2whOdSGcnANJPzWp8NrcSeS8yJe7i0oS
Tqe4xd9NWgKRzBN6GHebMHstemIGDCIsWT0uTo+PTcVaRC0F7dXc6M+S6MyEe/+M
JtfF0XOCJORmLrkmUXl0W316FHrVTjU3RrLao8/ZpbLLZdLjOize5gcIqZMu2bxb
nfs8dd2PpECIGfZPl9lpdXGAEI52jtDqhlMM5+Jn0BTPBwsuoeBo5f/H+OR1K9aM
ToRdHG0foATuXA38rTZKFzjhFHl6vrwshPtbFmlmX4eBOebZ3J1hkJBpqL8fl0Rd
cLOOLkGw+JGps2on0Q1I9ES+cwu6Zt8GG7aIx3l2DMloQWbeYuhEfk0puIGmTDNJ
Zeo4sgBWtcsoxyHwV+I1kcGKsv3hrbIIdCFNPdJ12vPoDFslyqf+oKJiKGr+R3yZ
Q1VIPPllgu2YWP8Y/jfkUxAFwpYxFcAy/eMzbYgG3gDXOsHgGWa04qxWBKXaCAlj
wAZ88P4rsJG64PHlYM7UsdB9EqP3jfrXOCOUbOm7cK/6w6xw25r6vQYz9VhjVTO4
p0iJOuSWUXI/xoJDWazQDjoDeYSpP7svM8+mCraDVJE0IY4tqzadSTcS323eZgCb
xv0Nnxd+5QkzQYJnqxBXFunHeGC++AJ6GKbIeLHgCCp/8mOEGbszXub8pGkylOSp
zjHg+MCyPsPE3CWfWHSkpl1Myr6R/nbntCiypmCmn0HRc4eUHx98vrKOObnKo5b9
ZW6weJblD3RJpV+ZSPpZSa2cBwVkBrSF1RpsKE0Wbqq9yWu+Ro82DSSk2CB8R7KM
nE/qKX+8AzCLnSHl11TYrgxs61Vbr6x27YDKMAk/QK9oq4a6qJfd46XwizeCT9G5
Felg71+y7lDFgwGK/k905ev0x7G4mTpqb839blO2CHxVA8O/51fJFbcDmx6rR/Fq
2ZRVPw96EKCCAMDuiKSAj9BmQfKNkU53HPUl61LvbXOwKXXGp193F9xhjuvwc1cH
GRm1rsj/zINDfPn8wWATQMvGN0aWP0qQ3wNxQZTreaaIgYNOoKEGINbvIFU60kL9
bymwo65ci/MpdvTW3p4DP7oubIZznq/ZDhPFQFnJK20yOulqtaJ+QSvVmEOS/ag8
OVV4kiCAjS3dXmlypEvMjJllGeuhi8Wr1vKt39Oziogvkw3bSXIvVRDnqH7T0MTs
KS8edqD3SkSqfi7jltv67zpoqOEEvNOKOe75fcknG4/QPaW/7r7Phe36qn5sQPNG
1faN599CEpb8mLSvuK215qekVESC0jwwrSIOMt6Y2OSjpq4ZNGDW/S3ZwnEHe2ef
4rTxEs8nVlHIsyn0VHiORt7Em2MT2bRFGQQ+qVhNYMFUifxnzBZsIDwE9vbwobch
9fKDNI/lBJEyN/kH03GFVaLxDKhW4dH5Zh6IPACqzGmfuPflqbPSLVvPIGg13EdT
Nvsa3m5zLLBo8RtQAzI4JsfCVVKVH8WoKTBSKcxTrAGXHmECeCiS6YGkcAwSAg3/
QQ/7mN5KUnlbiG01eMcCcesmEspITAB3GUGCdTnj4GSmXUSm07fPXjghI4ORX7i6
EFGOmBjSmJK9vBQ3ZzZHYjrNrLkkvqQGMnRxaDSCLpyDRFEmURaTDjYGugWtRpjQ
W+k8lVi85A9xZaYWSzB8TIXArdGPJcqdkn/rojDQ4q4WeVsnJJBM6gjZet+pp78C
58AkigXKZYNgRlny8otFgakqJwDXQ5Yb8P72mLcXYj0nC6Kc0X9EwDo4h93ojqfo
j3+qCzivSlRGJbEEeLa32qanUG9ICnUfolGJRD4r37LaJ0y7HQEVxn4y2ek8kpdD
ErqOWvIQcMeX2G+f9lbwfmah1dz8EjbXF79cvTdsVq9NDH+ekfmCMKRl41qp8vmA
pHEVliH7Q6qhjuDSVHoEej7kdLucB/NSii2Cqb4dr5HR/D9Zgk4+j9/MShtkE83H
KTeH4Hc861zKTY5r7NomR6CSwjyaUL3NOfZ/e2LZhkqC44r+Iz1spl8KWXAaYtOo
2EfgSoOt/shDi/VQ4bcHpuUr88M7ISKg0h0EabtaANKVPbwQSMDc25HHAFag/Brq
THPk8LOMZSJr+dN6jmnVQ0acD4bh8mD3ybASEsbPIOJnyph3DUNXboMuaBJgz/tQ
lkZcp0WhjJftx/ryOjLjjpBlML6HhClXcHj7wKnzGN0Ww5nojmQQzILu+ISFDNN6
awWkK3FKxn/f9B/FWTCN1xs/SKMBcurdr5cC7iT/UocnPzefGPuWdqB4r+eH3iU5
xmm9sQR74YIIyU5kM0fptG6l/spRno1wv354ANcOFrWOPAY+jNF8iCg4S1eldoXo
780JAI3XEmLDmjRBCb8+RrFcmFy+X3V3y02Upz6ABXrq+1opYu7Sjfi96d5UXyDt
Vy0X/RgessYec411bNfOEaOX/vRjxYMF+D3L3vgWxSF6Y7enYiF+9M6JM/637wPU
buQo7G5hhKFvMttqSXviLnoCPswnSGzt3+pcAI/EFLS/BeGziVCVMGupYr5TV44w
gYAlFq+oZchbOE1WZMI4hj7Sa4mmALcssv/ykJJ/r8VdLdoQGv2ZrEhRUfa/D/Vm
A6U1ZwezJwqia5JWNLRjLmIYTd+i+X3SAjlfmnI7jbNyw2SxBlA/5NWFMECWg6L2
iEZplYYRgD4qCXmcBWmWlzBOYHquLPJBhbuXflI7GK1IRsIdRh7HbNZcGZ907uvk
4y5bMCdpUUHa8Z8NwkVXDlRmn+bV6dz+bTKUhb855Szm+i6Oenn9q3YEk3XbFXsg
jX2MkLlcT0ZumwOUtXTZXeBPSmFGqQ4mqU+O9f6UPKsjxa/uqsJ8UxssHbFtQgyG
Nx+5hqvzcJHGHKouv51HU/oxKBzb3s1YWrAs/irbyagbdfgvz+a4wpzeqkXqPtID
O6QJfpiawDaRjV1hK76IExIU5I1RtBE7nQH0daYtN4ME7PUDUC4g07Xl+v1h8ZAw
LbnVGYozscqBTO3SZS32miZ92eNev8HjXimWh7UqnLJP2CltbRD8Hv0k7QVzdQvB
ouEohv4gYrraAt8dQQw1P+hApdCKoSJSoTmo+QLORuKDnW0DIYZ0kl15fJP4G2EB
nRU0le0uK9XYRx35Rwqsa2MYUv6Gbxpn5Shzrc5AZ+uU84xvTyMLAEe83cI5l8Ax
oYNGc6ft//fs5x/ITc4JANnc2otQPyJ2o48WT0upcSwUv7QUa6hv8kq5SEl8fZbj
qAnnQIC1W2zgGbFGXHne9lDomJpaH4yN+02J25e+duq5gcc2p0V6OxMggch4llhi
tep17G8wOgRvfvdGB+0y4rSju6v9au75sl01Ml8cfrtQdeOwCY26qJYIF7W6pl5P
Bkyegv0Vbso/arCJuVEwgDcb+1jZTUlVYXGhV2IeePzVaxExY+iHR299zDG7V//d
0s+RGulxgymfbt1X5uvnG/ZEQ2qUaQ0oflFYxNkVDVt19tFfY9L3plhraKf8MKEg
QJt7l5DdJnRJymSAsjURHyiCxGANolnEp2VVnXo83Nzt7ZT9z9Jh5n0O5b3VuJqo
BY1V2ymkcoGCsWMUkzLRGG0N4BeJBTHmBc+4ptCrCxYOVv+aRzkW2AYZCpwFsUaw
gSXiw446SruYCXCvLF4rycuR3w0XTYhPFJjMexFyfyvTyvkQB4usxH8ok3HHXUVs
611ZJfHEEoshJgcEIDUr6rxs3MAZ0WLIjZ6eFqjVmmPgs/+PUkoAZPXw++vXnwHe
dZWUoknHGJplDzvzwxETK7ccQTg9lPbabgLy6JVP523nliKevZI8e9i7NVrQdx2b
m0Xszdb1mk9szxN6bztCjDCAV4IxMKRZpYt+klkfQH/k3WL9JrxlE+1axzU6b6k4
KPLLosW5EjqFz42tCRBkauOGtJee34F45dePB6SGGVm/S/mjGeKC6XdaDPd4mDnL
B3y6bDv9+HYX3NuNpBtjGlf+QZdqkzY2E0qnfmH+P/hy0ytbOlfXrBzG3ThGPaOk
clHYqxUg9Ivzl8MP/82Gk8IzPsqydMmnCS7S3FuANHyByq9U5NOViXF1TKOJ4D5z
p5kvzYc0rXOaXJCbIFJ6QWoFz0OOCE0W7PITk2rbdeQD7X/+rvM6AdPwGfZCunmw
kwg/bLnk2OpAPxowRFDcvZssSLSAYbhJlGUCsRlb6d+uxlTg6LkTILKwgaQ6OXtX
7VXfGHYqXHi6zIA8jzAMvqvP4BWME2HDBxXepuVnzvHRK7NWGEJckvmPDmoXvU88
6TeO0OJ1zr3PpI5X6757hTqBvE8wTgFFX/7mNZMt12U4AWBAyRk9EgSvRThtZPWX
pbazNQl94wDpF+XstxyTRLLq67Bp4oZQw8vVkR4QUDSDQgc9YCW+7k4FEuyEs9H7
R0JQ4DUowNLy59maW41BdAebfBHXag1/hh88Yr8CzilJp2ijx9GeVZjkfQwPQVQY
Yj4cT1iKdgwxpqGh+pzicPTux1s3lxUCzMBodo/NoFjy/sC8izr/U58SUQ1uVlUt
T2EwsvQr5Q9sb4Xev1gkFMTnohom/DG9enWuXMWBG4JVks4xoe54snUsOvMqr2ZA
5TZE8QNIg7/e6IYRo78YI+/qXA9pp17j9AhQcNQZiN4f/QjXb37DIqVHpu/1OfZu
/axGBPd+jf9XKtuNudINGUdmTAicXRypUIMywRr4+bg0NUStG9iizIqbDCKdFxYS
8E0FuIh6iZevYhqDJ3SD7zPDqqav/EMLKS+05HFbvowtPUR6tRwrbNlyCvA/4KiA
ygqNnsocNmKab2sE6Xhp8QOXHAV3P2Ln4mZDroeq8VN+5Hsio7n+pElPThU9t74W
UYJkUr7TN80t0cweOlzHaaratlfpEhS0AmCqz0nrNlLG9ioVWPf2Y7+CWoOq6lEP
mwWvy0iwNG3ZDvIBtPlIE8F4MXjxC4JqV7FX43qAeofEpdKQWKDSK5777xumYCUR
HA4AFyl4XC+nYK05QrWywPKg+irsMzU35wRLcbz+PGymiqFuq5jhjT18busOf0Gx
ZACkYPgWY9xJl/Gi5PpY8fodMyUKB/Xq8EQoLZDdBT/NYgxgZkY45aQoFuJGsHt7
8MFuhwv8PDkBDlz8d+43T7WyKb11iWwG+dX0iyrZgBPpIDE+5Dl54ZV8TdOykM6/
8iq0YVP08YShzSyor5kHW6g6bK3jip3zjB8nMEEgnTNbGdxuqhdSlJgqpcP4NghF
8XaAdPyQxA0Dwo02bs7hTTJn1vTuauC8TqwbMOng1dR3axLr3RwjO+RZvze2VjrL
kxFbul3hJNXBKOkVVT9mFstzzJJpQLI5dCNFO3g9Z3QP0twd0sJwzrzw4xgyHGAC
W0eIOzQcIThJ9LdpwwWdpY4OAQ/67hhQHhSYpyOcEl41VTODYGwzAnI6RZMSEr5b
efCXy9WQ200978zNrTBBpQLXPjer7tN055B8rmZThV627kSsqrFWA6Tj02kak1JN
vGpOcFOckjApyEq3xeL+Zgadwu2qZn8ysAFk4LTdw/+BZIJBXUSnyO+TdufzpaP4
5VIcqpXS9Odq2udukqQdrDQ08X5EiG7Tw1ALr435mO+PSN5zRU9MhP5ovjJ92SRl
iNNylf5eR/Pz/EPClxw3PELIostLqtMnbZyxQM2xMSM3KO6EfQ7pPI5rxAStuhqj
1xYYs5AhepyO+OlpVBqJGQGm8zbfRAAaDt4+iedrLxeMRKFlIswee1UTx/50FCSY
SIO/RaPfCL+qDakAMWKtKieGG0dyrY7fnRNSdC8lsr82vQZOtQBX8TTIiAhfqx5b
wgbOtG+FtnJLNY83PZMyTfC9fP5JRhsL0sxigfBzc5ipRKq08NPaPL8XvMJKWKoJ
eC8A42O5/zeNvA+nR0bUe0G7OwwkqNAqG+WFfaty1RfTOmAvsvvCXt1vH9Ya3PJO
IwkdIZvckNHr9fcYbbi9kBusKuVg9gT6p4INrlFEOnplipQstvIeuYsgumQESYRn
9APKbnYk7aUUjFFNDqVrHrYE1Rzvcs+ejKEoTjZkTY5LNVYve4SF00keXchia3d3
hCC9OPtczpRNg6l2idnecN9uACSKs3Su/pdYt5RSpH/0RZw/N77tdXk/xd6BJW1M
/Nlr190VADGjtV3s0ySZbJ989HageflGYMaW7gS5ZFhegIR5r8c7IulwVwDbLQg5
iKD1kQg9qsoL7Aiyr0AD6ywcFgcl1PYQy2giMHAkU4983nPn2gkOYSLAU+5tqlz1
rBRVBdiCO1TMhIWe7ujF3k4LmYmlUWpcVjNLTWz9GlIXuosHyxYBwKiTURN3DmB0
tZab6l9cvqu8YAkhCq6L0wtA5gEKFx+wv0SbyvUU45qtUCwhI+ClBLv1Aqiwueju
clg7mbHhUWFbNlY7dOXS52G8T++3r7U2iY1xmJQjJmoIYxWbrFXrDhdl8J4nxOLl
6rDY8V2k6OXm4z+lVMW1SxkpOs9joOPVbMbEg00NQMk5wJTZH9umI3MJnqCAmGa/
6AaitqG0vNrPrQSES0Yq11FVMdua+u2Csd8HLyq2GwxoLFQuA/4MwSEj0tNSQ6Ju
D2i3CTfipiEPtnS7ChIaYtfgMHMn1LwG0kXapAM1iVmyx8oqSBlNZfPRLQWX03eh
o1oYV2hpzk82WJZrKHvAJM9izEWC7f5hIVa8ReH+Ui/K5tUkgIjDnnV6z+g4snEV
CT6HUe+m44CF4CpGvrLoQrHmfEOcKrkQWtV6XubnVCW9r21oV+NJ4WqFv2hm9Or9
5+u+bDCcfYIRV4cfjxJp9DNjKV6QjA5nKc13LfolFLeDunVCVDq9rjMOuMwOSvSq
lhpa3FxhoLzXTIVE/NS5lN4KYchk314mIxHzP4mv2Mc0ZPiVUx8oBMc6LC5+mFP1
0AgXGUT97AjwZwEKZL48bezrQY2GaBpO1v/+h3QEFiS9zwVMU+yQF9zxc9/bkoBn
Kh+jrDsbXEhGHZy6ei09267VtxK/a+RerLlNIRnR0fbXp+u1MglzNNDwUbJPBhAD
Y+a5mXmUJr/UmOr0AUWruvLnbVs6MGbPtwIy2ebqji4oGMLRvPXXkopem0n3QM4v
xNo5XO8OwU6LxiofrIfGT+2wG63A3/DWDCE5T6GQQf131+qGuwdKqBGvYP+YhKVC
AOqwsaI0y6pwUOjHtvoCACu+QlWJVaD6zKIRm6H1Xh45gYQgk8ET+vDj7LPQicED
eM4gCVQ1mj4B5WfHM2vmD/8Cl8VsX7knc4QPyKX09QwWsT8rbzJRhX5WKv7Dg7ju
Tg0h+nL8IQDSQUMw0LiOW+VnR+FzLrKhRU6QGDxvOEJN4EyA5EE1KIO9fLe0eKg3
+5lu0yO2R5WD4c2aFphAh4849CWboSkpCxodYiPLE7Fg2I0kTPqRtU7LN25IiWMr
DmWngO5X94vhUpRxTmViaSOEuEl26GbCr65+/jUR9lkby7jYjOoeCQwJtfqj628T
tgXueZyxGSHhnWR8ZMYvgSUE6Fv5F2eeeLMwkvIQmcDg6XslzsJGY8re0mWLhVOG
18o6Ug+A/2iaboCefcZTZfrmti0wUZ78EtmJ4WAV1+X5QaT6DqMrOkraz9ulOSEU
zbWFJvoXVWPXSDbrfR1IHKBCgFFi7YYQaB609nfH4a5ArSuY/m6NJa5v4DY2W49K
7nzOnz1trRyRkmIYuKzOoTgY04DlZCnbZArxq/BqlvWiNTAlqW6XDCc9t1d+tFJJ
EWm5MfTPWClZJUw8RzojYyhBP9tJWyh9Wx6TVPHo7yZX6o+M2xb/LLGBl5JJ04VT
wxSHWeeIpNlXbqPpgirWNeGpHRwPe1eDe4K8Ouiy/dbNigIFa8ZsS3Gk+l/k0Lov
luXfJ/bswnrgBExmgelyFjdV5yivfFXj6drHVYfqG1Bd44Iic8ghoTvg+bLpQvG1
9gvR2pFpR0uw/0CHmAyPKwpVd4jvgZb4N84jpwfzbBSSDRGY3sETCpFhK7uVSOWd
2YtXVVm1V5Txrm3shfb5RNhcWBiJ+YUFeBvsjSJ8zGPwu/9FLxhVKAFv7F4NDkhu
FOaeGrGgPne8or90+gP8YS7n+tEnMwtGYSjbXj/EPtvmzWdiBHQwvWCXh8dKnpvZ
bGKGcfKwGkIjt/eZ0+8RPif34V3w1l56xqAgZUA1aAixy7ToQOrKzTBzurbDxEOe
l2XdrUeCSAS2hYurdLpRiO8ZtM64yzrmjqUJdQE8fQzJR3WhLVngkiVvWkd2qpMh
+AXUxNLRrjc5TxTgIr1h8Dfom4LnsWIMo38FA04E3iy1GzJ7gBtAqQhYolQNllVu
mUvpe6sVLHteTQwXfEr5RBlitX3Bz5duTRPQI5sVxMWIZjCAStdlpEmagPPMB3S+
1gDdvKsmotWqeWUjCnfIxGjsD/wz3Iux0RHQmR4fXt98wJQEnIOtcjTXWuq9rxfr
qhwm+tOJ69ZWtlhHRXDuVGVT0Kn4tlcwmPcVDtfo2F/7VAyTeQ0wTRFJL0PQKYJn
ZOinYtxecnAHkaw7/nOM+D8XAqBQJsUFNzk/Fx9T6a8CfXEk8HDQac9sI60/Q+3n
Jh87ft3r9X78yQZF06ffhxGaqPY/SHA443A3E+cz1/zs8lz7eip7HBVGP5tU9kB7
YyUFxbip8zVngwQKEahQkn6iqKwC4uZtml10KdpWqgY8KE0JD0JonytMDeQtQBnr
CgHKrnmFvU5cO2Hmj2Kpe77lkoqB6OmqHQLfqhdFQ3CmxBpPCYa/O1j20+ulYhmT
wHAQdjkQO1JOoZIyZtF9CSHU4tYs2dQwMNJaa/YHBiiUCXWRYt/6F9L+xD6fpvk9
4BYxYTDq+3A94+enloZZ7z1gSYEywJafOMElVmIuzYgp480C035GcUoHEjGZm4cP
3Y6SBmpis+m+Q0PAakDazcJ4rIvUH9c+bT8o249Pjsh0FExicIBN7RCp+bAJCvb2
KEBfiSZ/gatUlEvFlDiplaXQ5WBroPtayBGRxd0JmJMm/SHa2/sQN7RNQoJbcmrn
i5krCLCLYyn4Dunz5mW0qlaVdXscYxH01sJ6U+BTcZnQ5xnBhTxa9+Bl0LYquvgB
mO8AR1JpIBljLYIUHPZ2Wgd25YKQ2I6Qj96kd+B9aLC+20E4vn5re8qvDVXW2rIi
MJn9XUm/Xf9G95JPIabJ6gtaH8Ha0p+yRJ8uyMnI0Iq5h/9bBsdl73amK5pC1ifY
U5qWt8ybaBStH6kckX31lLnBRHeQ9a7vm38+nVYybjp/zVedMMrTEWzkTtplyc+K
uBKdGJmiB18XELIvKHv6JKhkJu/Jo/4lehRWMHjNfKtjTREkh5yo6ueWcp2s/bNx
/eGwTHbL2aaynQ25OKZsb3crF/4jfTH7z0vD6w6BB7dwrG+q6bQlnTal0hXIL99w
zLjWwosnCx/KjKZO96Kus9+NfaGxeWbi6EueYe+9xIv513WgLOjlPs3oQZIQXO5R
EPfzpCuT9/k0+KgedKm7008x/Jwp+ykTk0ICc0xFaCHXUiFjrCgFqEk1GqKUoAsh
+wHCApvTWqQv40r0SNVpu1yESozUmii0Pgm4SucHRz38ga29QidmxcM9mO+8LibV
CHXHqNbhFqW0pYAKb7OO4Gp2kn16WpAtn+H2zGW/KepVihoiTmA70lpGlEef5rMZ
YG7KvXlBgezNzklMALwRKEG7GmGh9Zj/Fq7eZpW/irAOv5620WctmkYr75mtFGpq
/Z1RSpWw9OOaNApDr2N6poFC6BKncTYn6FhrMX4Xu1vF2SBEzqr0T1LOVl77Pjaq
wtEnl+DRwf3XZZ7llEATk7zxzZjPk993earXCC6DExPqad2eMbtGBrlUK7lahVwh
WE+32ZnaeGlq8IwHbCKwvBOiUM7zL7evrBtiuU42Gns8HKrxqCw50AuLvUzg9Jgh
2MCwd9fiTWFs08I0Cef2VN7ALXNsj9z84FIlRgOcNy3Z8u/MU51sLHhYHTlxoar7
vmvIBIXoLBKapccjcc9CJ/Rb/JgMEVFp08blgl6812o9L02DbESqcu6loUPsyskU
ReHNZ8Xm07PCYoiryrt0I7UaGYpZrybwU/JUCerqwM9J1zbqvj5LTVNbSvjRuAMr
9SBl5+x8hmAlHFutphfFVy476fpk+PQFbAiSBN54I8nnAWUEMy8A04kSaOcI8kBE
u+NZO956PKFmi70uvZA9B4EWpD8vrIi3Cn5sO4iLXQtDufEgalJGv1MTw2ccvVjn
GWuZjixnYEMqpwzWabKilAz9s/jzvSPWigrcAB2A6ivKbCeSuIuHZ/U+5FV9ZRHm
Aqs9QAEXtMT+I7YETOP3a4oW28etGINwzuQnS06ZU6gvZYUsx/7LFKbAyXVCNhre
bYhlrTqrMfFewY73wd+7e+1ujGzcQDJRknJyngBllDP9c6Kb93lihVZNS58L8RbS
aryPsxHF2m8pmY9Yl0Avy+rbF8g6Ebpdc5kXzpmjdU5eRodvw4xDRw445f7wl9e2
i5Z/1OqQ2B0kMXQy9l/fruDoBHE0a5X2C/wOtcQ8zlXkZ4Rj0JpoZT2ijiIr2DtB
hRnXiZBq1KmpfZue6zuiLqlSul1XybUGkyhG9wnXHl5zJ4QeyUzxfirN10Iz0jGM
sryBkKtoTCJ/PwycoMMtz27WwLSQydIdncyRqDX8clly0VlmPnc7tiGypY15Jjwk
XshLecNz15Joj4yoDiJP94a8LtznUnH1zaKk43s4d8cb00nKBYwGKiSQZShvs7mJ
N8gVLPlzKQ7IPpB3JDgY7SQn4aW5oDDzI/wV8VbP618i0EjiHVd8Zn/ET+XCw3my
DYb+OAcem0pA/Jxjd3xHrrKVc6SBMl83YprNdT6AVWdPh+32mZ9kNrSkQExvjkaq
OwTUtx//NQiTWPIdBojGX8PEWNEPf/arYNwrj26xeL2VEV38szn2u92QtDTw/+8E
yiypeQRp1HrtBhyT2p2OyHtgZBhWvG88noOI6zwdQeDsnqnQSqOVmw/0w3ZF73X7
H8VmeBEp0MUm4t+9G918mO+86TB/Shis9eHCBw1d/DjMG1ONfV0zI3nEk284d8St
MZDEQkphAN9EmQcE5v9EAJIz/SqM7ZMxoltStdM4Od1FFSg6DdmN+2NWbMZ7lHwJ
guK1txrqOp22vZ2jRyvpkZ5QPmRSBRozmHYNSoosUl95ELVI7KAa5hhZVvk4Ck0T
yRQkEkYm0VmRF4i4wxCPxbzBDN7bXMH7cbbwz7QpoX7w3tNdP4v3yutxKzIIMJCP
pBqH5j6gSWm1mS+1+fBU4MlDV1tlLi4sOlxY9v2yyfUQYj3zA3xLRBG/rKCfXf4R
p0juU/xC5IL0SyrRTvS8CjYm3yZJX+c3g6ZE5xoWT/dW+zc1G0yTNoGQHNanL9Hq
ydzFZnYspSs7x+NqTFr/pWz4071ytmz0fs83k3ddnNPSLDMavxH+i4nR9PylguD3
ehVqIoT0gAjHdawW4KgaZTWA/sKtAq37UEB2ZLr4MtNgFa8CVX8b62uAn7Z0rqzp
QOUx8ftlltSTn5aoRbuSFBm08bSam6B0EOXGvt+8NlVndshW5GHuJvzigqiEGdtT
p1gwMWo03WfDiBKZNqAOuIwtzTPMskxbRL2HHpGTgaJ7jwy+HoziNSWdaUItDETn
rhYTMxpO24TROW6ZMn9YZc2BeiqMh8zAmirHypmWlQ94BLw232E1eLsIZgOouMee
/rZVagAg6QTxZYfIB7HwIegi/Aifu/neZ5K58x6EiSZTVU5BpYuswm92GaOSkpiw
f4211rgXW1b5Kq25b2gbeEde10R+JVz3FnIySpNIrgmDjHY8/nCOqOhXshcQLcoI
zbhqDLKDXN6SbLCExgLtLlkeBf8LBMoszFri6vwc3nCX7F/zOZWCYUVzGrnDLRAx
0OUf04tx/jwoRXPlIwFpMK1KvXAim/OLOGHwvLppOY4kYtMQX8+xN4u4NGmLnEk7
0yVknHw4R98xDYDh2FtbGvYidOdKMKIo4dmU9kMQjE54Low1GDz5NHGYiBEow8YG
h3OBffzfkiCAD4hyCxkIJVRWKZzDPmaapBcteNT4z1F9f4OUf2TLF6K49HeJB06s
T6P9eIWiMsWBNKcSO8CpJTecu/fH/IeybeqzyaIfIKalEdpkMP5rJU26IqZSm0Ux
XVqXkRnaqBwL20ZEZnJBZ6GywFpu00AbDQKhy/L0nIiJHAPrQFs1d8gi68YYNiZB
JXvAav2hpEQjKLENLZ90Jlzixd9FlVSoPggEbRlHNYM3ivwxhlOUS/+8SwpK4b4I
RUqPzJ43GOegKnD2KLh9GjuQ2yNysI1+aM3e5jVk62WUZruAaIWWCt++TK3tf8Sg
iGjDaIRcXi/LpgHTxHxFPWNwVdzLZEq24KKwJykS8v3XJXMDgEHO0/9JzDOHg7T+
/mw8vuvT53VbVmDIZjYnDEwCidXV4n/8FDti204iy6xcj+wNfPfkDVZkbjozOW/y
qa9ZvkNCBBLmariF/PiLaGDH9I/cPow4eLl/R5fVIkGQqsS1R8idddt/Gr0kvAgL
KnJPqXwjiLss/2WQj/uUnv+FY2ZosJHBYwv06R8cW9l44GftfVqsIkxxXSoX+GF/
qakEo6hnbNZrrR3O4tqPjCL3xEHGU5zmjrFZjytDzwRyjP9tydQgnEkY/A8j+C2P
GvTc7R1A/Fcr1wzAvXo0fQRJkJlXY92lvJlI25V95Zr9D/NWu4rF3ZtrzKN0YJmT
1pkpxLdZ+ZqeAN+PhLwDs2LFHBLWK+pkTh9XjrXBOdjzCH4HRSE0PR3XXNTdQQ7g
wCExsTra3X8FdeTycKUGyga5sR9WRro2g+I4lKF43QTPkpavtRAsI1D37lDqy7i5
HxB0ghf4CSqF62GXz2DxLWSh7hScQQbxg6OWltnb4CRsjSH3dNv8HG/xIee/Atus
4IHjSPU0nDm+tHOW64u7JSkpWSC0s1bdDEL8OL2DXHzHjWPRfI8WWxNgbNneVPMR
NAsdVqzjWg0Yrjw6h+CHxoU2aIFFWT3jDZkSyMNaPStUQf5bm/YbZpj3N4qrepRi
469AIs9DZS2yRfxSaqxiM14fuDAhZojBPNDrr/wYg5vs6EEvtV3hii8wg60A9lLz
zZMBa8dsG02j2sGcp94CnvepHq09zirDOrnPko42AL/gId390VU/bdHk7I86UPFr
8T0BPKaRG7QJsYUdaM2yT3FHmgbA5A5suSTpJgjFadKG8BV4s3kpXcKZI4mwJmgi
rKuu6vFDXQdGZRGqQYRIu1Z/6NlrAJu06xqltpJXp+lmrtlj/o6axLzTNmm1C75u
TxFAycSX51QmZOUOUEsWJxF13WuY0ad+7AROtwL+eZqWRknvHi6G5LitumzNTQWl
YCgDRMLbAqa7boNzEmUQN/RQfRLtFPLYcFLd5PBioKYJWIDWN99DlEZHoTabGjeS
abN8w/1uJUv9kNr+FjPpOxqZ+kfnbqbATMTCb++6taeh7d+6Rntdf87/R+a90rnD
5W5z+ZmwttNrg/6XhgzK0U4mIg3yB6Rq5SS1FqewZoTTmXHTwgcEN18SaOkR7c+3
LnwvAnWJ0VZ/GAz6HeLB0hh5tKHsgjiTiwP/iEj3S5MPINKrkeh80wTPAvEFQC6r
6XTJMkAK0JM4O55xRmT7Fvq+X/3KpF3SfYmYlNIw/xjGUTtB3fHMJ9iCrYl6iOr1
KkQ/KSAHuHtVkJN5Np2FFwotwIaDrHzkyQU3rZ+YZ8uySYxMJwwD4qoBwIq9uUqj
1OJNnXnZqwVGui//+YWz1agB3ognodtoetRpgRvNYYzl+wpJa1uREqml/JolDQsu
ZSWWvO9lt+j1hd8iZcoPvOHpomuGxXNzcxpL2Xhpc8R7CBi59hwKrZ3ZwLD+jWx8
BOLE01ytje7wZ6/7gDoRAFhYAcZvR2zHCl0gyFnFkB4r59OACNX1yLTV0Ue1xS4B
Y0xDTL7CegAxeTZAB2DSk3IG8St9cm47jw0X9IHPQmj2rtPLxyx42Tf7JLNtzBJn
L3fpPh7u5lxdFxO3JrzhwEAt8kN2ofuAJZEGQeke7yXUVG5+5BYWrS8j8X2fvGsF
Wsj4PGv5HinQOYuTpkILTzImNRoIXePrJbIu2hcAc5RIAjmyCT5a8O/GO/WFDok2
OgYCxOhXkeafLj4j7bYvbdN7DkNP8q1/wZEdqOwSkTlpoarev2lT2ulr8Zrto/I2
AtdBnAsyWTVy+haaFvxUFxqLU9yHTeNwVJCdY9iZHTOXN10ulz630rmNOt1fQlzk
pYdYacYhde0PeMKtPJfETHYcz1e/BgIhyKhH26lFrH3GdlhHPz30smNpU0tkv5CE
uXhoVlw+IUDcdz/r57fcE0iDRB+ikP1/A6cfVy8flkAVt70M3OX/OVkTalHFZc4d
nXcWMqEd7d1F3qxSPfkO6GNqyXftR2E3QOSrn7JMmF2klWqIYRfRuNFqHQN07eLO
QeK25M/Gzlu0Rqbzu+cqfvZqPOOrasCx3edHN511yxVSeGlbRL1H/VMRa+f9oRZp
2xlQpxZjev5m9kHCN+qSSe+uHcGNOT7vfTz3JFEV1A6vjQA1T47+NNKa+ifNJrU4
xEPmpPEk3LTHHoiSc1gUz349DUhi8ZkoEv8irYQgaIJKIl+a5nuKBE2+JqQ2BZzW
vnbnt93sQMVH18+253XMnA6inROQwgwXVXYEpuSffPeddISNIVp9NarTXfb8WBgk
BqLDEp31wGYtQ0qs31mLnO4TFkpJoJUc8KXwqNPE12U5zGZN+TRyO06CfxQtd1WA
6sJudsvIpu6Xl5t7EAcRkRnGLZZFN/A6zNsF/DxqrcbIBWHfkDPxWTuqfCOP20HC
9mQduptcZsSQ5j9O4h20UQQCp4FeHNIJ195h8qy6NXLlp/MsZ7ScxrgZ8XBJoMIC
jd5YVWQ51Se3rKTnyzsQQxdjB9dOCA1YHYT9/GM2biSWTU6rWy9eXrTa3Spz/+yp
oWTomdOCYi/Rgz7gFWIiRIFAtYtocD0yyj+t2ucczWD43U9lnQnBeBD/SdzodyNv
hC1j87RHL7md7TIhwEj7i3qnIvyD9AI5eHBfPIE7QUXjkW1e3IWWz5a0aMsz2TdA
9UWaPpwLGhYGVj57MogLRqyR6LOV7f4mmMqK5aDznzPpXWwyOgPLHlRW6bt5WbHQ
AgU+VMsvNt6H4fgIKUOcTF6P8XvAcuPpkM2xfsOaQsCpdVCA93iA5k1tkiJY/84V
a2snnWIa4RFhGQgSx/Ln7WVFReFaHrWsYbqpjybsXAlq1KBOaTMjHntcZjN4wlZI
sd5e18RY1pPAtuGjP0AmUGG3S2y0zqkCj/Arn4edV3mZe0s33BBmIJ5rGCPq6R0q
AHbQpOPvusiQJRQccenNJ0BAwYL2JRgnuE22doWPwOLPyiv+gHr2tvW5/mPT/STe
h2j4coM26W+KcS1MMJNeRtysGmyaH66WN5gUcmru+KWim7hV1WDAdp40f0UILF4E
d9LPl6Ik2L3dMDRxdBlQ79Pn5YkBCSYzJPH3dYR7UIIQzzkQfwwCT6zTwyU3mqdk
f3t0gVG3NuOeQhDF+HIBGDfWD9Xnuj7rEgEdKhjXjnHkuhYKgdnNp8UUeIuCqP8Y
/EwsO8heg11Zmvdfd3RseZXO9J+G73kND0V7wiT8c15E+SqXFHNXr1AFxFARVblI
SYqh5GZh0fxuouCdqhvSnmARW3nkJkwwKD44t4C6d8VAVGUtHPbIqXOBGNulT8i+
BiEWbUPwMiyetJHyG97crAoRmbj7AswO+TeNGg9I71r10F1bjOhvWrOH8pQjp1i9
CiZ7lRbE4fMP7LhYsTeHhLNuCM9uroRCHJ839UdLpi4cv0ntU5mEjy/kuOirqQB2
LVAFIRHR9FeI7qiaGPEyoOGTidHTcGEB5WEELYgTHxhmlzc6IvWa7LvUyYcPAW7A
pVxf0XjoCs+jz7f6MWS8KC8Tjnfk+q3ouKny79nXd2cjvVr6LLyjbgl3LGJEGKLE
UWvITkzeITsdBd8HuvNwfsWYEkY+EUvCtvANKvag9tcZzkMwL6bS9Q0ec74Ef/c1
0KxBMVRfrBjZueRMBqer4RxJTEsE3zUK+BbKmmN9u13HDBJib2goxwcffU3rgmHj
BKgCHbJYXVmFbRJqZWEsZ4ehVKFS7cn5FKDtdEb5ysPCw14b9UiW3nn4VWB9QGg1
GMmT8VkIhOxG8gHUU4l/aWEAxcPtlsv9uAoWjDhy6l60GjZeyDn36TOXPhrS2j/C
50sB7vTaeRyUhA1sbWmLIQV71/9Zo6HbfzPRrKker5VQW5xA1pUifkEx+BdN+k3R
/lVYM235HbQa9lsCB6rCe/lsskYTUUDla8SR8jGdnhHl0lo6bXFCm7TpIOQXWCjV
c729B3wZJERTzu3ppcrU3vHN8NuhzRwcXyH/fY2u6NNIWOSEK4M2g5nDXIJj6tjR
ECGPBxg4WAPhUs6sYUyOiL8+/T6Q4PGEMCxMzNkjb0JuKbxIiNVpgFNDiNv3kITc
V43+xs0hTMDi69t9LkpCG4xMjxwCwufKgeh+fD3zaDU1BSZiFBqrxcXE5P1f6QZO
lt/b2OVRQwiHizCPTpz9baFKPSAaPlJ2ldg6D4uCQ0bxb0lqJvyBYY4qEbrZ9+cS
krsbPh/YafCqHjS6TbgAmcvXO+j3Pp4rl8qQcQnZwbhgqydS4NkAUj/UTJmhTfkl
6LE3BMzSvYZPnfhJBkbeuobT4IqBstWI7R5aJByZ6fSLRfijYvMnPHn1jUrxHGK9
OxqWiYeX1nyJ4rwXGysgi7BxLx0jzOlaWFAib3YOim99BhDfLh1WMPVR1MQzdxEB
hE5p5sAjSNOll8kdy39UCm/sWCUTOQZhjTVJUxnyTrgscydnXx7kq0xT3eIN0zC4
qE1Jn1cDB1qEXH/Vw5OzXpvaq+iIFky0tMVmDnURpUYunqsAch/ZDSnsk5sBYara
/eRncM5Q/w5W0jK2z0KboJ4RLIrGIjREbMl8cGwlXsLuTYEyn/BAHPpAmVJYv40k
v5pUFbboAQc/YLeO/1VGy+B9NLw/faQJUoejzSVVSRcUjZibn4TWsTakhTLcnULx
FuF5pYjKlry0NubGuvb7/jK/q+QGGR8MsTCLLnC4HsQD6J+6CUOAo7G/ZcdnaSbb
+fe1+z1LdiSLN5xMXSCh0PnsxYNZvT1f2FRO7qke/Mat+0VBvlSbIINchXo/iGDv
hErHubgJeGTspmuzbm2Vzwl28iccljffc00EPtO9CD55LKVzXgPMkXfTYBuPHIIe
tsDqUAAAWqSSkDmS37W9bJBaDyOt8h6KudI6IpMrjto8qAZSyppvJ89PjOCSvTLT
bsD900bcMvzdYcGA2yEZauHssgijtdGyS1IWXRvI2mNAjWKNDVGw0m3E6qGh43Iy
mgW+PDBc3dGVyFDFUglr0Qx411T2ll5GkxWVC8T0y73hmTmTkW4zv4W2kr3ooeLb
bGo34dW7GMEHULW4ZjA5wtBkrN+aXU9rMAR9Gr3E2upZGhdWbKOM3WzfXKzxcywh
lUUQqekJvzUcKl8N5nIqCu27dsjIP41CE9t3B/fdXkJZ8qlROVM0BXx2hVmIhoEj
Dda5IHP/VcyaKKi6a3noILsmb2sNKEb2w+WAZiB2ZQuUr5W0jbx43BrOOslOdS37
aaa7v3mNSrj0SPblwdWdPH8Op05I1cGr/MdRXq/eFb4rMcCrglqUnqcXouFlSzQr
p1PPzXHinPrGhLjN1pXDzaxXncPGw2jbCuD/c0A3+56c/Mffn7MD94nGs4xF9Jcn
0dM7FaZ/5WjYRliPS3kaehqdMBOwltsZo1lshVO1Ymmy55Nn4ggQc3De2oFN/Sof
5SCay8gfY9+qVRd9tiG0l0ZNWHves73pPRuxWELYVbkofCX5b+u5iiXzAVdt0Myr
KPYSSCguWqK6C26PwVsSbY9fc9hgDgY08x+feeWS/9zyqjrEJMGOxqk+dhQTPV6M
CpuDMnm1o5qmdPkgcTsohLwMKOW5vaa83QIPJFh14ytV6BHs+nkJR+m2DF8ibR/J
WAS7sJnaW8WZFl2bfABp+4vsO2pT9Ugr0KTKMDusUZ6EEHzuBRNtwu6GB/KBf056
dKeA1RgtZt/ULmN+2Ivy3nL0wTtHPBaMaNA/H/RCMwn1acBMOvhavOu9le6cWOem
6qH105tN99U1BamAIIWu4jYR3UJx5ZriLxWFy+XdEIAmQpdNV6UVVRLLeMAZEyO2
O6ClrMxEFcVKu9DuKYD++1S2+Y3Rgp+5KC4WMmKeT8YGuH1LGSU/KKERlKg7sOr2
EcAk2lW+1i6ExoPxGYnFbT7io91HLE+xieBXCq2KXDwaxq4j4E1R6rzxLzzHGqI+
tesIHipz9BIxxF6bLeU4Pa0FlQjCcJRC1GOtJMAH0Sw7YXL4eRhueTS5tJrkROOH
BSCHomGMEk9QsSJ/YH7nKxHwSD4Q2A5Jlv+Vfk6a8lOO1p7hnlcLPXda8CUUFF0J
Yl5Gs9EYOqh3eiQKJacfBvd/ROpaD6l7tURYQKUF87PAy/FU3P4XmozUUjPbK4si
MsIcnHAwMlbvxW5sMdHvK3fqh6htPIJvsYnXRSB9/H9LLWpgOe3G3xe8mKlhUwXr
iMdsqpJ4Y9JCDKiNnhHLkfRVOVKvks09+6FEEFvyUh1GPw9S9md01DbwZBsUPS4d
4Joqk0dXIHbqLUSY69hsAAssG7i2AK4QZF+r9trN911o4QGlnxj8FsQ8n/okjlXP
dC4WmM2NKS3sULLQ/QKEoiL+8IrWHhFxWABnTcKyCz/S2pK5CGRg8QGzzQ3OC3lp
5+vEhEtNyEgrHRbn/2pYysYWu91Wg6JxXFCR5lknRIv5eFMHro8ROlXHP1wpQ7M7
2G4dis3d4Fsj762LPNlcBvWgXZwM2zZZamIlN4/Kb1DfAlNXk3aTAn/PQKfVkQgt
1y53YXlN33iHwWZO0sTz8qbQ3ZhXzvVJL/ffDcAIEQyW0U+ldNXEZISCMWOM5sEx
JnLztr+57jv7knxcUmn4gc0xHsyYjPGcYS9SmIclmd2hHEGkmmb8I0IgOmq/ChJf
YWmkIpDolu6DFo41t73wI1kc+LC9MVSok3a44UmLZJZDNylsFsAZf9aPV0JRJtgk
OQaSEdBwiMjPG2+I7H/+Hkf7e6STHfOyOw+k4Cc4zqUXAw2cioYHj6mpFwG1bx+f
3S+xgxz1CL4YZ1RbbDnJ0Yt+ReaHU9mKzeijnVQtJC8hJSuLfsm1/32QfyN4zunI
bJhL7tCARtT0SAoqCL8K/pF88Ul8CDfxO+sU65tb067a5nSQUb+1vOVXM5H/uk0a
HcSbLCtOC0Tg85C/53o0UUZ0rywCeq/3g+NX79cHZXmYMp+4DANYQAM1IWuq0aJz
eSnKyg6rFq+q8238QVt6ykng8Nb7LTU5G7J3FQIpwFbLcLAgE26R3nL79kCg7Ai6
2RehXwtkIQ8yCLEkrrw8GDw9V6qz+Oyq1TWp3V/7ydXvx4TzJAF6ByjIEqazavGN
7X5YsBFdNJalXJ5PAE/xjr75zMZwiUS8n5pRojuuzp39Lswugac0Ark/0A8lGKpA
X0VEl0fNbD+kIzHQN/NksA+M5y8WQecx38N8pzSGxESczdxHpaH4kbM1MkeeeiFH
CZxt6S5DiOeSSanb706nBm46fOoyVY93BiBRcGAzbx5Y5L85YSrKXUo6LrgLfvuG
gfPGnQ1Mcz3netTsDiHqU5BECAPUGudUodYM4D/HthKiF4xBglyxYcMW1VdE3Sl/
Utj6M0n4mOni108oV0jtS8pUkoDX3ur0dImWiEsvqcAB3rwOHPQPhRJwZLPPq+ZB
X12UVqjSmKqhXtLftIZGe6HNN/k6mqIDnFv1lhKRYq4Z3e6Fj3uPkBpX+WHuguG8
wWWLXu95FWK2k6qHfZSCNLyiq/9D3pjy0++6O0tSBPViV5n3+LmMXfv/qBniR8di
n9vTAjPY2nxTlODJoNiQlBlYz1fUew5KMQcg49ca+bK+qCWJEPR0u834E7+A5Vx8
u1OrReFI521T1UN3tYOCBOGgpfnrXLrbsB1Qkboy0NTATIFFfDeRmPfAGDAdK160
JlQPWx51VaC7/S0dznjopp0T/C+MvnY6W6gw5gxVBMx5SI8MHeMQCu79cKoXbFst
LzvGFzz13OusIsprbg9Wz/1PArB6qw0vmdBDKRZEjsbgqRNUfgUsLnfhPTx1Q7+D
bXBFAMjsUU/Nla1btMNoVGujef9kDt4rdeAAkUI0ReSxjmP2213o/LnaaigzUEoZ
o8LDtfM3NH5NfFW5oY/Il+aJS2GKtJh7DHC7o6/rhzxxXsd25ZgcibSMfQ7o7F87
CxnLj0zTVnbZ+ZLKFAE6PqxA2y3IN08dWUVuT3m4v8VwyoxmWcv+ST3U4K1Trc/K
MHNp+mj6IFXVk+ZN2dfhL+XFq6M8P6/ituzQDaexbu61xzPfCeVnae8t3ILeA91R
/PXKi7/VZfM2vv8Fc91r/+JWt3s7YBSQ86+V+ikiH28bT2a4mv1wtUGbfGvnvu+8
ppKt4Aw/jhMx7lk4KG3mBK9N0tb2+SVkEIfd978WW4bAld/iLn9zdtxYS6LszGyI
xI7K35511iC0/OSf/D1xKjVB1W0ki3WwRBtE2wdC3dcCg+MoJ8wX0eatGuSY0iic
pcWY5SI7pf+qkjwsLOK5MCbTC0EmJs+FNcetxAafq/UFKpM+roeRaf1m2JHvtOpU
2Ab5M9izNAcdaJStriZZfQGzt5+0Ivg/YlnA8hJ5YiJY8qk1GoB2seshmDUM4xpS
CBdVy2jYiogLyLpA0IVKpiX+SzEZ6JKC1cVKmHsVJ31f2cpdZEmiYLmWsjCA1wKe
+INh5VGiYCeiQ2DwbTbIdlfhP6xGJTz6HIOXLjtuVknQYQNoiTFPNRk99/QyDQf0
okR0SCn4hZSM2bb5zWl5Q+qx7wtd0F2KZNjmMN634xyPZaI643TZsu7tfCN2nARs
QH6HJ1eRMQQE4TsU96ZUvunfgyQuOdY8rsqvb4+vkC74nz5YXNTm4pyP6ovAhAuP
loHwNgUv2YJva+pOrc1NowJPLS/HxFH+BTV4TsY2bPv/+n86yDLkrOcq69URElxJ
bMEZtSrbbBXw2jL3dfd34YM7AnypuHY/jItYwCegwb821QaFRO/qiFpcBvP2SIFz
gzpzmSaFmJEqE0tzurNglrn0vG7hJteg2VkMYorO1Jf4f7ojSCoSTch/3N/Qnxmj
rWOEJvfZj6vWNmNZjoRU1tWqFOqDisyG870Mtl82IFCsqgQ38JB0AGSOIIOa9PAS
gbgpSJajZbOs68w/rG65QbNl942BSdKaSemhjBmYRfqL8WK7gr/HiV+2p3XjEneN
/NTyXmhW7F/RYLF8QIdWEEn/BM6E7JkZjkxmqsa4uU2UPq9csUAfL1yAPnrFh5q9
IP5WGP76hyJLq6ACHGI6DYn9lVRg5avEefJIRQqNWDSf3gOXUHdp4e0cZiryDose
Hnxz5dvqUJ+PC1JuvvBuYZ+soEX87KPYSEBa3UfbXXdJfTpSefki3x1yFmiPr2CX
YZyvH/Y8YYpB08YzdWYjwkINQ0FHhnBgCsZ+VyneudLoPPTwnifDXkQUfFvWGI2f
wthB9j6mWtFYKhvmMDC5DI+eYer5fSxxFBzuSX4wcEEbtaa/IgSHyo7cABIygZ/R
5EzV+x/L2c9JxuSio7vB+3jD1c4dqf9as0NB7COV6Iu/Cmb3Bkmq9gOqavBhIT7c
o3QMshDTccc1Tk++K4Mo9K7FYzSjgW93n5MPE1LXDWWLg+4sl+JBH1uMGsP5sBAY
t7i8NAdw3VdKL+fk4oiRS+xc0SAhzK/gop/bsy5nLOz4ojELK3nNcX0voz0fbjXV
aeBdFkbDSjadTycj4bQ++zQJMSG8XNQ3eGmjslH7FR7wOs0NnIGyO/HvXV3Zpdqx
YM3QATbk29UhKHrapxcOoTs8TqrrpTYxHa0ZYo2uD88mbfI1U78n4u3A/1evmFmQ
Lfzv61TOjWsFWMm+fk5g/vgRiKIPk6l3eFqb7qxScz9oM35udm7+1NiwemiS7LUh
5UMJVb05ULZtMph1bciwf+73VYngywzZIBaFh46vUDSfowlnyxiM6C81wStGQQKa
P+R+My782xaEZc/HwvP0kPlB/glCe1VsfN9L0ug7wfPKNrQnd3hQI8wA2r1jxA9I
nWOogBJQR+YsqbWeKcOXgDcw1ROVdYVn+zfzFyH7BzJ62lasGsG6LJiLwU3iuVcz
B2Z2unMNNPvfFQGgpSI4I3cSt/jHoOb/FWGvQxB2+vOjNyvloKJHWeepF4CVMtXV
18SL0y9/202+hUAGPg4lTe6ouU0BPW3y5xU+8PAeLoomNy6MmSHlcEgBfzCC1RI5
6o5uiVxAsf0h6HNDVcBwZLMo9cDvXtGZSgMPjAavws3euiRM5iaFkss0zowx9TyB
Ls97B7WjZCKipPhhFnHJrc5scgiFpSpWsLt7QZZo/XoERShQIq6xbP8R6Fj91eQK
UDP4xmUTsLL5SeoMkhBM7wrYfr2wezgkJ/VbHPLtpe8thgRfQwnGoIeLiYvdQnf5
g+7pise9Ba17W3Xzcha63qhbvy3FBEsV2cjSKNym3COg0RKHfkQpeCOOFVHx2hb8
oNIJaYz615A/EBGNrFvl+JoWN2d1BiQy0XTKOaW0gOUpCIeEtX9YTSSyVQPS6jzJ
lKfDnOFUNQmjSZo8MQGiDwhEn4mnDOKFcCbkCwRIVJtOuOHf4gMCBepyMNlyUpog
vxL6q7sRa4q/hn2LEz0yYAZUIa3+Ont5nuRnV0XfJisd38zIx26NL4nZuPFoCuP9
thHcE5296EuUWOTguI1mSJMgR2C0f66UvD0cdb28beCTPp4+Cwlt1vCPGD0uTpAs
NT09SXidSPOYI7LBWSOftdt7IfdqXpNNDo4BTWcbSH1OvlTbZUYvfTfFeqsbAWIx
7DUj/oF2HIGMo2Y4BJ4yafc0girgU5H8m6e4NQsozpaUdC0Q/zxOUc1bQZT96oZ4
iE1pj+jEraksDREiOdvfH8XLNszsYbkoHfbKkVYVEaaSxrqKJ630Ll9b2rRUWF7C
38EZB5oCoEipX6fvBg+u9fNwoEUFe9D2AbVjU47NKtAPqA1IK8+pxlfeGWejWH+/
0w8AzhiLTIr7zMHFMOj1SjRI8oDmdt8ct6zRNrV0uxbikV0GW6SLMSl+iCvnF7Ma
kAOdG46mW5n8iw7oM/F3FTxPdmu3cyddFEweJ+xi9XT/VJZdJiEdEIWm9dSebsWE
QaMP4ngO69LAZalv1GaZ5PComx0dqnJ71V2q+fNIPyLtvNIK1reeWmimqmWjZTzK
gbXXjGF/1CmYDtJ4p+BG+Lwxm6gz4hnMk8ko5A2maDCpRRmy7flDhh1/UVEr+j4f
usk7NJ8zN/1EJU4TyshSObCp5jZsnbOA/0Gh+PyxPAr5VgyiTe2QrsZCFYpyf34f
4oc24rrD6ixOuX+pNTbj/xAwZ6IW39tORM+hjZhnu9dnstZGrRaSpQlphVGQnTG2
1H3B0CCkU5UXkD9nefVZ6bJeYfaFVldIjBkM7o1xy2zg6PboVagGBMJr2CrYntyg
jmcpMoYtTi06jNv/3f83fFuTXKqG9OeuPnKt1Gspgl89+Z32/XkEHOZQcxwTYyJw
ujB3Y4eDqo9TRve2h5NgqSGzsEe+G10f3hr8lJRPj7FZ0ibK50ZZ/8d9Cm54OH/4
y3y97PpRI4uGJsLCOc2tJR+08Dtv/xIxDx41ekjgWQqU66Cf+Nwj9spipfnSYJNs
/4oZl1Uj8v0lZ6KQ1nj2eJqS7O4aIelPAGrSbdBHjaTmQ7q/cd7WL1eir0JPkWHP
dbNwWUw2IDmD0jNYmHiDhSRBW4LuL2IdbM2GROYM9/ALIaZiq3ajvK9ved44oLS8
ryuWzsd2D/RN6r+5FRJr+cp52/FM4gJKG3ENrEpwuOsUWUKC1PIva43iN6bNJky6
6qmKsfrvdpLGUjmQkhzYd5C6bX0DKVsjQC317+FZXXZWMMyrVEw9ZwhTUxy7efyL
SRy2FWKHTUw3JtH3Dr9meoKyke7/yifPC9RDylNKbeEk33IdI3PHq+U9B1xTxLHv
hd3TwhxdNO+DQLfazZQdv02/n1rq9VWGuFZ1lguD3woDkIItn+6I26EnN9OIlYiD
yeOnHJ0AuXEXrEkfNcZ86rQeHZsyWi5V3VCE//mLJDOB4BdalED1LsT75nDSaq8p
p7p5g5f4FEwHz1a+Y1DRYlo4RV6Cosrdncqgy6Oo7TtoUaUJpWutyQ3+YmWpSrf9
EbtBlERJdkK5i6+T8MeVnTf2lPmWDL7U/uAdGlnk6yqiYOhlsYYT/0nasLfT0Tre
nJVUvDxkOdrlTjhHQg36WdWjA0KRSzBy4pSAJ+VLNlx2lQbvZLO6zdxUaVcdA/nh
qTw3fr9yzIkG2lZDuNp2KrIpFl4a6BRxnClGOBnJkQ9MqiDeKQGFTavg+cxqs6rY
XACHTdsfbfAc9bMeBshEWL5ZGAwExaFY6+H6WTWAseHxUdTFtpPk4Kx80wvp5MCV
0SRJlJemH9FrhXgXnAWhGt/+Dw7OtRq6oc1ksvq/7owpe+DxpeOUucf/0OKKqvtV
nfIPUpvIMs0RcBT7lCzxnthiRJL9+ZWTgoOapDPmBh9Y0/HLcbH487wJVqctol6n
WbCH27yznFb3o8dDZG5a0B0wroQrS0B28H+W7q3T60j5v4nHdEkDnXBwn3IafYW0
uuCr7CpXMXGrTYfHOp1TlZmxI7fXyO6j+smnzUXmwd8V4r1q3okFWOixaYccbXui
7BubHb3SzBU3nqgRpFDirJFwCZnhW4WJDlI2w/e3Q98mI8dcMXmJc/L3IzKk5YJS
0h1hDI/kNNi4S2XsqhAP0U2c7pNqm7XRbfTgU9uzV1p7aEiUIwNz9I2vN0wTE4+6
iY4v673eCeuaTDbihKfgU0GcuoSsLg9FKTMtJeu2G9bjen1PhHEf1viyQvg40Vu+
nKjqN0m+qlm1dVcmUqHZ9U/OxDhsZ3tYzR5/zbogx4BKyRCe3z7ql49HCTFI16C8
e9c/qlYbHyG6oP6fsgibluHoz4dQhFGY1M8TvxxXe7ZD8Myg7+E3NpJAA/H3USc7
0mQQRiJSOBj8u8G4QsKI+dPWQvX5Aquz+8kUaX0b7bcmuGyvGDzrz5rtCmmJRHQa
wtiWlTvI1t9fx0ZuefA269SheJ73ZyE8OWlyOs7wObtjFS8tqJ6WrChMyzOV0PHQ
bimFVtvNbDeFGaaKnGttMWiIDFDeArPOjY+RQUnyii/LvqO7Dh+EBcPaMZyZtYYJ
1nzixSAofU0Gkjvpnly6ARUnltGWzmGxplVod7dwk36CbYezH08lVPl1mTNPFa4S
N+J5AiBTtt8qJ5EHHDk9WiTUQKqmQhon3KiW48Pg2tR0TBAQBJ5kNuwmsZxFjj2+
q1bU0PzVoFPaF00lEY1doNhXV6+X52Jrtm22FMjlm4Iyis/sYPiIKp3hWogdZ/qn
5FydNPT2lZmyyfBlR0VQcKhKJWxYi4VSd/mhY3UkOhvM1DBLRg/FQFrcIB1YbE8b
m+fu48z24C1rJgbZ2nEixyVJS7B7VJcavXFbV7ysopqwqzjeXW+l3ISerWT/ix6h
2RAxoJh4DxtdE/6hCEgYTRi8XDoyJlk0WjhnPUNQ7nChIiWRY0oH9AuZ6ExkQfhc
/koUxpBJa1O8ITYdlVzg93Wu0nfXWtaRITGhm5suo6u29e/M/yoaQfkGwLwqscYF
FA89gcbTdfgYUVQduRUI7dB+jInyVZmyir1I20BM7w8mowCqdDdt6EIzDIiv/ZZr
t6ETd7GiUIcPN+vUFmhCIhUQVFFIPtucL2BxCbWUlFvc7j1hDSjQsSWrGChju1Yv
pd98iYLvfRDKs+grpoAB8s/qDM3OjD5EKebl6eu1etfMqR83AQ0VC5CmowQu+Al9
LDH8FSvzYMPCZt+3UokElKQel/WzGrVbNL6/n2XfjpgHGAH0j4YtmIUB052wsZD1
5baPkvGhQU7PDZd4f0tLIjaXZ92BJ/UZ3/0441c2AU/jqk5VjqBd701P18pZYi/H
KAphU5FrPGB1l4Moo8pm/lxlXiSr9Z/0so1jiWApoCOmS+m0MY9D8yjLz/43CIpQ
iT8+wFmEAA7OM3xrKXeRWAjNm66+K0JO71NRQzvk30qCRrNQsBGzKE3nm13aZymw
tRzm5h7cvEBChVVklElbMJnCEHCFnN2A5nq7+l451dOASrX4nXP72M/HkSUnvjNb
gn8yvDylqJsycXhB6eEsbDbib62eWGvhX2/pUY1+Fz2SEQkRKy+K/1ubKt4i5kQV
22OSii9wMkpUI3nnojByCMhVM5DI2K5YgYGCtRDg9N7TnYTLJfJJcM2lHAohzte0
fHKJG/F1NIOT9RC5Tqm/i1ilxA0ty5ECKJKpV0fgEpYX8QO4dmKDvj+nwcQf4MsR
KG/LE4XGAyY0pNkhBH86tDgBdRvr10z7Ca2YWdyItQuGDLSJGqNys2B9VS2X7A0e
vvE4GWZgaZdFLQ82wqO8pSnioHqMtFozB+tCI9TfwOtANaopjKeULFSnaiRwZ09b
TZnLFthwuOWzRKQjYShyU6xj3g4Fzarg80d24JSEMJPjmgUy/GQhaupo6CbR4ztl
lPXA2xt8a2GUnOapgMCEE/HhYpTpFIcESr2nOto4mX9JM2sSwmihaAdLbJUla3pG
ocEKtuO7gudUK2+ADU+TekuyUyONo8aEUVpygAnsCBWVWtP0tS517neqgrd+ncWR
kTLFuWr+JaJpT8lrX0wEl+bOOkggWxU0g4j6G/rGfGs58l/AD19NLwBSNl9yXC6r
+hYTx2cQdp04BnehLh12TZmR+joZOVCdiPnqJRgkmPol7cuDFtz/VlL8KoLBzsqE
xRZuH4YEjshkNMg8jgB/yNh91/vVfnLrHEhBqJqCGxDMdYWNWDiFk/kk4yLvAPz+
SyyAcRYS5BgZKD1c4/Cs8d9uMtIaCVGNPbhycPAJP4OD1JDpccaOoua1Uu9oLs8u
0AluKE9a7yXrOTzmJER1FTal+lYMzBswws7L81+K6HyVryxMVfWJ/W7vfZuzxKVg
QmH2ael+EFeopwWpTDtuzXSu0yO9Q7q6T/cXjzx2PIjfel8K/SYQ/yAxZm1boyW+
ccCQuARDsHgr1Lait3Fcr38HKXmbgVJ8gTdk/ozf3f8+WKHP1IphEQH/qveT98hS
1nAiIPPtYAPTFI0sA006n2UxXliaYRninvPzJs5NFG7C4XqKsPVyY1f7taPxOxPk
SNFM8XDgruJLfxXQke91j/ijmTuLpgFzYZbaFVou9GT9GtWbI8u9C+jT/NY93xUG
kqs/EZl9c8Z2dfFYKs7aLuMik4RWRgwGIAq27boyys5anvQkW/Qo7ALObkSA1ZPJ
n3756W1iFevFHmCLs4FId6v5JLmzIK7aFvLU12Ai0umW/zxcLC8y5riMvbavDkTP
XZTU6p03ETwDgMHFu8qTfxnyifJjZ7Zx4ZoFtoFaSyKFIYkay1riYqOJyx9uIVxg
G/S44tvXq71t8oCgyiqtCuZfDVXWTmdmHNF5+Jl8KH+7knXValcpmge/JjdQFrmg
VKU4pbkjR51zULzxf1vxqOv0120TiF4m/q/u7zxcpfMq1uqCAWsPR1G3ao3a6kvB
c9R4tDD7Ai5nbu8IKt8ZisKX7nL5FgpchJ+ZiRGwEVAuwM4/yorPTAJBRHbOqba/
U+14uebytl/zKxz+5syNlOFFBrlDRIdec9TNQC6SEUfz+d8IHKXyBWbd2ADrotR3
+lcATcnmP+g5ds3eVNXL7FpY+//ktbFpu9QiuVGcJ6X7FfKcISocz3gMFN6GPkLz
mlkbm9bb0DKBbIp+LBY74RRKzJr77A4WVw+BDuWjUGloQaMEN9FSRENphjhhgu2i
ni3rjf5fPvrf3l/uh38C9+KhVE4lPxQkdAyftlYLY4607Yramqw5lBJv9xnhXqaQ
EG4VbC10DV021lrek/9c/CdUNscK67MCrxdkRny6733q7IZ6vfBKD+1J11bhUe1g
Of/5itDDMBioe+lHVOqEjf3o35D35pX1hLZ7R6TbxmHIvrUFewqpxcpK2iUvt5ck
M8R0XGJp5qxsW93SeRCuJ3I2hax7GSrQBPQ705gFnE1ObBv+/QahjVph7ZtvY35g
DY7HyXNe3B6PMHLTPwS3IPZNTnuNstecBX+sjYDckrVvKAUtdUri7nsWZ9PoX1vh
GU/giTdr1cnVWnlcGqKo7xiU7xUYUn/WPM77moAwl0vuU2fKMaf3p+XpQpQ8jQJA
SSvAkq2tYg4VeDL2CwslW7xOfiFJ0dCWe2Ohl80J6vW/4jjZE+IWTOopdbx0pn0o
vwJxBfJc0hw43TTNgLrGCS8UGGkwmxSY3vOEht/4YUnBYbIy7+DJrTQ/bpoMAU70
Itpmf+MJbws/yOVi+pSykuX6ZdJZtYI6AV+EDXu/Y9+0ef9K7ZwvrGOhcVGn/VNx
GV/aOn0qurIiRZHMuJ4s+0bfibosfdnEluV7zdKeqhaF/GKNviHdCo+e4FQN0HKI
4iTZTbhgLrOUhExq/Sr54tfANFBTxJN/T6I1f1c9NpsveNOXVuC/gFKzPEMku4FD
+BWQuIW11wnfihpa2Dbfm7OWOJEukAX4XRbTQXKkllPmLqZwRBdDwhvdeByxCiIU
E7u53rdXtF3tw14fNZhaGnq/vkV00qfIpr0C2DGVf2XONoJS/Yyx9roaZspVX6yk
Tah2jydCU7amMK9wrfwjWJhCqCDNEUNrwT3aGkU4YGwYErWZcYaCW4yr3BJZvkQQ
SqcxBEh5WAeHibqvRD8qBClxHBdppi97IsWVHmVwe3bHMI+Y5DzZurluZunGKtYm
funbk8zUfD54SwBc2vC5YED9Z5G+tMDNOAELT3A+A3ExFHvNxNJ65JWgfxiQHbI7
uU9PkQLJFFBOS5augOBCdBbfaC4KCXxCnrvnqYvMw2hzsjU6Y2lda6FhsCAAbkfU
9DtihUmlsKjuHxRawMeYxw+vYxEZidMzDXJd+sjqPRdNGl8ffVKtdbPvJhf3LNTW
jKyFZPtxOMin3OtGed+6avfJB7h8vL1mUVEb3VpnjPe+w0EC+p6XjLwSyLuRjqAz
OW6vidWVIkvh/VXqMcIBs0f2XG2aJidAQELjGi6T6BsY1KZTEM/9gluKzp7DX1qv
BCJJvZUKmASFsMdVLwPnTgC3YNb7XaqXNrDXBtqv1nHzAFy1zpt1Nane/0gItf2s
14LvxBCGGzo1oUA4I9kUz9hsQWe6JEarJq0kizSdxGYjVwop2txnYWwFES7e1nOC
SGxTRoUbAgxpOyR4NOIZ2ilTvbRqc0O9pGFoy7lnrUjmERmGr3ZYtRJmnrYBNESe
dPeYe5fkYtBsuzAvkEgbM+IxgzOtTiEEkDRMXNYW6iDnNu4hU66PicijW4E0Z+hf
5z7/xreStPxR+7MW8/Y7Z9BXnK3J2U+15i9TIfCj32MJTvI2ORVQntaC3Q0Pu0A3
3HQ8TQZqswX22iawllymN9k1NP93vEUl/Fcji3yzLQzbAJCUkHGBRJVRgnp3Ny6o
LJeZGP+q4QGQ+OtArBTYCGkFhmutwbsmdDj4cNbI2o+V2BzsZda2QBDVtlbQGc1M
TwkgIkGtl5IevoRZv4pqwMdBy49GiTsQA4flZkL6pUzdb05lJpEpDNQLPvgQWYto
oY5o/GBkb0+hePajcXWAWa7Xpf2GRx3mkhm7wAE7B2aOYeC/aJcmq/K6/E9EASa9
MKLujonZiPkLacVqXxLnTG/Rkr0VLWydCZK+5zfOvKi1v6B+FPZAsKS64ZflSpg5
mYtKIoOqtvi6ZrKEH10W0E58FQLgfdHVyFbDW1AOnf3TyY+eSM+ax3ODieO/wmHz
4cwy/pc07sBExHLYsfFt2EpsOdoesV3/BcNPWkLxvQJOUlqwKpIufYKXd0o2nh+y
ARbgI+SR5bp/qzU+l3w3lgRgQjsO3fTs8soB3f4R/zjc00jXDJg/mYfQvBhjXwQI
E4zh5UYTjVPZkokbQJnsvLh+lIfBdijNAs7gMyB8eYUZQkGJFcVGDK4tN+UqhYjd
v8mDxWauVCpZlzNRl6JBjlIp1hmjwcpooPE7ETJ40oQ1gPcStau0h7lXyxkA09Zj
WzG7Cb72mJe+AVnErEXLrQ6kY23ZZGV5A0Sf5pJj3Bz8mnho82lFqvTKMaCs+QMZ
XwZWMxNVp9CluPxlmi/gdksGymqjjjHLaIL3+LO6MFe9LkjBhUaet+4Wey/QZoHL
6C9zqIx3KKdLdLF5HFutuH03xPzkhyOzenqHc1kSTd1BgZ/H2sIr81mMAh8/JLHV
f1RFjRiU/3GLeuc2oF6ulbb/iZO+VQhfzR48iscRrelFrwvTI39g8kH8u5FdV2d2
IAe19RfcT3PZSJZvaNOsb3AWlgfH3QjQCDhH4rMoQvkm2O/BEjuakmvUH52AsJwm
IX6yoEXXI7hNT+20ozfHCBIy9yY/dWTXGncGvcs+rs7hFfg1qWejFZWxZ+mJpjLZ
ECY+idZa7BGHSM8yn+Gf8r+p9fyZCzKl8tB6Utoqp2Eb/4PzAvzbUVzbr14Th75T
NFJOg8GDTcuzVcRYItCxVbUwOyZRmK5i9+ECPjxybSZFbzw9sULOoH28lwSi0yct
Hbwdy3JjZX36oBoqgXJmJAZ9pCibVj0VxU4ArjoSmzzkCwFEKZ15JKMDoJ0JcjYu
cbG54evl8WLzChb9lwVSNeohuxIHGFyyLR3t4CtF14tJJq2ZyPQJRo4WrKdXIOCF
qJM7evbreICuQpzM/y5ktQkuItY8a1k0iirxBfeUB2gD2VXOT6u0Q27cWCKrbgs7
6ZDZ7yRDQlqdcE9TO5TWkGVq3HyWLZhBEbh9Er7QsmHxnCNPIYETxCFa/RHVYNS5
T/vvxONrFp97yRu0Y7z1LSLUN6kD1QsSZIydvKKLZljYmCKk2MIaghttGYSipygR
hEWzegQ5X6O7D/joKcwY8c1+g/KP5iToWwyD06sO5TwqOuC/kg6p04r0i03+rkLv
Euq9cOFtx6HRYSaA7wb3tORm9LupdjSofignVDyVaVt8HslxThT6FhVi6CWEh7W5
ykSmRfxJaEKHckmwp9ZHnrrPG9tuvEBJxQb49p2eKFYcNdNYV/mX2ptUXbbVD2Sc
E1yKsFVdmav/JXeFGLQJlPEmltX4sMA1f5epGy3VXZ9TIFgCsREj9IuhwI4nk+/6
U1EVEImMlpp8A/IEbCki9zAUjsMkC62+YQGrcAgjH+n6FA8OBL2wBGERiN3sFKGD
ADJ8EiYszP7YywyTCBL+YNnS4VLfnUUJ27rkpV6YEOq1OnEtzuMCKjTuq7h5QpCL
8ym39W2eXIMhVSGLDA1q7QPfAf5OqdEdeTC4c4XD13/3TQPoxkDEXm9LchFawk2Q
Pwm1ZfRcS1eXMCB7EM2Y9QbYP1kyuScvuaUNAFeorB0NSnOSrKHvbARBgUpOGJ2X
ep58t9PZTCBdX+eTfKkrC9qMLf5h/HMmsU1bZfb2NoksYcZcL0DDChlFssZ/gs6w
PTLff9da0WqQSvS9a5DiiJ1O94y8v6BSkkwvOm3/LadS6d29mSEUB5M13K8wcPT2
Mb3SBPcFRWd4nJHsDBL4Op08eqOyz1vLApJ+5+FCCeaRVjFoPxr9FWw1361oWPZO
p8IcfTiOHVS8b78i84T7g8VXktv+XKH8ASuYwSf5dHrhK1nLZvUWHA2p+hLWIdBx
Q/C2HhLxTQzLv3IsxP8hyaPCLsZNfh7gZknsOn8wrLn0BvOSPHLJZDkNuknWu5Sf
hG7wUao4sF6mAGjQ/4vnITX+dBU/dNloeb1J72KCwIB82oHVMtYn+OB4oOX14G3V
Bmms2k7HvSu5JP9y+6UClXZkpOO0v0qDkcFFRxqtebrFuAFOnAtZDJZFeV7+eMrt
rGYwOMye/gJwYTBYxwX9+4xB5EAwqEd5TEH51rYuPJzMx3gn9KGpCg+ZuIMoyqko
qMcZdktrV31VJjUQYWObmtKYUczlYwT8BOMu8sKvwbG3DVrIJoBeSytE6FFPXhpS
4nVysYcqXLiItm962UgRNKNqrU+xBmu9zgGtNsVw7ri7U1pxCmCuP4TpGdxvrF41
ouvXNrJQei/1gFXqLBqjdEi8ISxUCm9B3THgXchHJP+cR7//8HLNjI8s6D3ryyIU
4VwGMaMeNxhih1qDHFmPNfbE2CcZnMS6Ir7SnOyiJ6vpArxjIMP+8SkEJp+e5/V2
NliSAJos/+rbIhYM39j/oGN+Kr6pGplQagX/XZFiNdqH4q15KoXhB4QiheBD6wme
eAi7Vg81V9kqiwyJ4FetzjJ80h3aBdYsVy2r3XDlW0TS55byqKhVC/z0fVSy4xJc
foQyaZJHHVCrn6oVuCCif34ha6OO3900TkwYr1uNNm6He3em4d91qczTPcZ9p/8b
FCSgiqvfIfVv1lVzt1eD18OLOYFhRgUt7iHpPlbjemSwG/7Ib8nTe4SAQsQX7fiE
LScAXKtjqY3NontkOnhscVQq2frbgqzPj79CO0oLAdaqaAYABfCwFRSuaiJvYXAw
J2BYHl1en4wtgOrt6y/fMnnsy0r+eQjhghtad8S692PQ9QHbBrCvZWOPedNuT6ZN
BRQNJ5blQmrABzNQ0yHgXqV7gdd3cJJ6KYMSKHXzmA4xaAuBGyzELo+kLRH2GZ4R
82AxNPtONjdMML4SzDnocCkpbJVa5jPzk44tGwWIG2EWvryGtVL0fYUNnzabQ36E
7VOEXbbGksO5QCiih/Gw4VjVbz93jcT1Zt2bU9MyEkVsbTVXR9O0PahEaEfoaU6Z
p6ia9etaFO0z5AWWINcFso10Czf0fc28tDKBdZsih+yXrsULHDmS5J8z6kDopY8Y
WwWyYYaGMPes+xywk8gsibHrBaOqSp6/dbDbFbbaVvIDo60qMEbS6FHuJ0Xx4Dr5
HmM6q1yGPqI4DXnPAvjQF3ZNhTqoqoeUsUVpCvhWj5gd9Z4FCm3JGxOdu7nAb+pd
BuSc4iaipV0TJkOqFGyx2tdqqKpg40vFlQYSPU1kV05h3NZU5QVW1TfBPG7oC1uO
st1ViFp33ilQZLes2i3bqZAwuaD2gCNH9glA94CfuTj22H9064KLsYHB0EcEwXcf
TYAigNMpFoAnWsBPDOYuIoly64xiVxVl308F8UUjcPhF79Kasm6wYgNOxZ++CUZA
gy+nGyqP8sJJNuieq86xgBSDj+/ofDXMRxhsmXrDwX4oZ7gEuTzQggmC+F/Nb9eF
fl6mlrXxUj1QjU7abqRl2EoXoVXkS8aV3L8Mr57BLh3IVxR/pGU2iW5F2TkjXRc1
rH7eCHz1wqmKLon3vk/tMnKu/4nxWhJhkx9J85/ejOPj1Lfnhvqe8f085AK8RElh
q46+SYz/VZtxSZZnrLG84Sobok4pUbxtC2wZF7oDVWQoZkieMMeXIut9+mwQ7ScA
BPR0Yl1y7DLzTiFyC9mkAwCeLdSt+5xD+4xPCJ9I0CZZKg3SykxT1baF6EVrq/Oh
kuZ+AuBodL1bRxAjn0rJpwdAvIlwq/PZGvebE6tSIEh8HCd6EqhVT/a8cTUM9w3J
zJZbqusu661x86X0SfBYOHB4AZ9Clo/HuOIGjUAf+E76076Z0a4zWmrCU5uHi1jG
LAC/KeEe5UWTJ3QlbxJy9MnRA+qFDlFXKeRnqE1033IbVJkJ2jhQB7py8AHkxHfB
/sCLhgbSUZKUVm02Wj5H3NhD4w8QSxZdAuSXx5r2JvnfFrRLlMcXKwBP2jeNu+hJ
qEFDSMbPiK3fC63gY/aiYj7yL1KEJ/f14/G2BQHRArSWpd2pqFuvBCDaWLgEWq+u
Q1M8ZypLk3exVOSG6SNcm5EwbYQVcABZSfCOgVxocOditWtqy7kZDguZaSytPxes
z91wyHOYU9uQaAWmCZqk7Zf/I2YLWABtYIdm8Z/uF3vrXOupl0WUyXtsi+RlG24p
1Il5cXFSZMXXCElr+TPExwLlGnUJEouv2zrFbSPFAYcLXzn+0leizLndK7kvbgyk
41rNGSV2m3QP+g79phep2oUtoqF7gSaRK1d6FO++x6MknNBo809lHlMk2x47Lgp6
gRi3Tam8Zg9McvItGPqPOQ2UNg1tkkB9TLGEfrFbJ/1cI4guFs5E3YJlbf0NU6+z
MEZDYzRVP/lnR8IKe3HOzpuSEQwUmMxaxzUw84nYey9TK6vnrSK6SxbNHOMexiyi
zej8EoMeN/RtEecGePAgm2oh8V4q+eF6yZ2nF28n+IeGSX6aNbsKzYEndk09JH6o
T0Ca/I5mDj8fqbfNYOMEUgLv4R4yZ1OesUvHvA949Uu40+hbBucSo/YNeNBtuAo7
Xn9x0wCxhVj6NlOfnLamlpgFea15kU4AjwI8uRRA5ur+naNB6Yw4wulIEuxAtXuX
Z/829FI5Rx62GGEou909UDJwCy/6mFpUyn5P2eduQmSF5NNTcVpQSu4XQmWgRaZ1
+FZBfZwUhsdHXkbA6BZj/wbPNph/1K64AOq+ODgfVsJGAvcWIV8lnNuPD6q54jpk
xYKhaUpqss4A536FLAzdk9nCizHMPLGT8fftjhoDEL9ahEQntPwxFaaleMDCt+N0
YaFE5A7okuvlkfhdGXHMoT4Fju7SStqEI0QuMd4VBgXhGRqZEYYThRTqkkbcZ1jU
gzQ42uIgzskoh/wExmnlQjATE+nS06ligRRxLG9dFGwy07C0FdkCdoqJhcM90aA8
Zzup340wNGGTTqjc8B+Gaj6l96u81orD0mTHGLLtEfIcMCYUkwoUwwn1BjjABbVJ
TKswBwDELhSKHI64hB5LDnkJ1n3Nr9z9PTMvYJb7RNKCBMAAxvnFtmQkG34ZkkqB
GH/oJlMIg5oxSXH4j+M8VekAM4oXf/wcZbw0MBC9/jNn93ZqGiorQ2LnCgNJpKH/
Kg5n3hdEoX5vsO78YaDJcLPFe+FAXWOY2ISEFzSHzD4MLr/srlEp9KLgNAJNa5r7
s8dOv0QOUluITuKZ5SXnUSwPLr7GJtpSNiCJb+mSKiPxqSgLEciNMRt0ToRVgOSG
hMQXo0szQHB9eg8QIV9AZ6Z4yrCplMpCPRbYhY5H5U8176msBAe/NKy0VS7uN5g0
UGgMOA0zHIyhyOlSl7+tlLx7VJmMyxBqr5Ch8SJxe558dsLfZ9JLuXx+EqScFQpa
0X2j+VxE+VFpiWOzsKvqx8/1WUMLoaMnjqShlZYJxofJe6+PpBWrHQCsFW/Z50B0
aX+CS1lUP/JpNoO7yuaQzpxs8vC8h8xvRvMhlX+d9M1Jhso0viiKJG4YM7PqWTQK
Oagdxdg1oXKuEW11paE+ZdzgYqJcHmasDkUuvWKplm9DkfqSR81esX961BNMBLDP
vvyvPNv9IfXDX1E5+JjOWxTBjKO9HOQcTNeTYH0ROCueJP+YSgNAnOkTOYeyInQX
vziI5gIqIeqYoaXui+ASDioMwrymKRzDc8WNIy7BeSE5cAyqEKuTFjQuQhGKC2gM
vHGOAO9jXihYosOhJr1w13Tk7ieZpgM0jdBuoKpd2pHo0DS/ySBPQZcadd9A7IDc
uL1NVH7jSBJUCeASfShkc3Uz/EVgGGUVzWvCFni6hHu6Ha4OWzd1BhwiP8jMMdhZ
/LLBcBe4mOEfzIkjgdSdCEpiseei8cIjcFQZKbqu1IyRFcwifMR1Y5gNPdqMHPPk
yKzTsPaRnNwbkDWFr9KxGIQwGpLT25j2PxGnzuZ3aOeSO8mOpug9UGdh35XEh0FO
vmxk6ENllrrGqVY895H/fbz8y1ljDrUt9YcrvSYpdNW9YCw9dXuCX/HpGLz2O92Q
dN+vU41980++m376K2+KxcWZofq5cktCzO0I+DUL4FEJmr23erDcQAi4K7rXLhwE
8jxYMCuqBlOqW/tk0xCK7a9uhJTz/vQqQzzVGKKjDuTWVaoYD32VADQoWHy4E98F
CSbF/Y+f+BAqPpu3w1J7qzOSWtVG2AX95tcNZd/3wONeG4K5ah3WdwywQcc1pVp/
W656Z418cZx0Jq9erFFN53Z8oe6cQy8mDn2BlYxGNXMZsmi1oh44ZuQhJa3BVPm+
jdusRhZ1cnFDh21/d4NLotdy8WUm2549QeP1McQW6jOpHBN4PIPgzlT1aET7VhkN
IpRgYB01RCHnSTVR3vHqapZhJdn4K5i04LcxfXQzdHygx12iwvsrlhyntCnUiKNr
O7GCCZwrJi63p/R0pvcfpRkl5gu5wIeKOtU2qIHGFocvQs/c4AnLupmDXbHu6PEb
eB8y25K6bZqJkzNHZaZYEQxTcH/ZRBjNozyGHizNvzou4jhbpAehwDovHgYeEj4+
Pm8uCgpu61AUTZE6/r07o8IEQOD6CGvqs57+Z20GBHtsTNODgOFQ/kAKXlS7KPr+
7Vc2uDkE4lDkyOJst5tQSRXPEMgoi3c5A3l4q+E86cN4pwc/3peoyu4D6/1HOMAt
+FNC5q5N1+Vh6fGEf9UPnm3as4n8oZ5qqya7ZRrKsY0jbZ3pr9j6VPaV4to124rS
+cyjX5MZ2+dKPxmZX4vnLOCA52zHo2DAwuUHeYpSc18XKrzBlh93pme3TR/+gDf+
Rp+ZBwmzu6Vz+ENltFk2MG9cPMRZjSvCGHN/D9zfzRxT03eYj62Bh93AyYjSbFl2
2Fnsxfy1zy5LzIlrLQu72JAuFFp2n/Vn6EtQeycTnbUrErziYqWksTID19NxeIE9
aWXwowUAUqCT8oesJDS6ORWf9D9QcOerV6S6gVwmAw7EiZtarKpp5NkCRbdxkgj6
JPVDflP8L08DyJwqat7Fqv5AX8JGQkVFPOXOhiObjs+vxrqu6MSAF0bsffJJco5f
xdpbDAEHParKeo3d/y1zJAB75JeLhhg6lmOvcezPEEDus0e1Ew4lkBNt2I5PWl3R
mSRfowBiBuNDnoO8kb3vi2OW/oGrpIijb7PxtFSiw1KvEnEUc1gm6a7HEtpzh3Mx
9tn0CmC0SOkyjqOTF2QZ99d/78Ls3weom9DCV4ISqkHiil0OPvEn+pBTutugZJzH
Bp0nFOMXmQh/+fXSYdBdLYkBCN1XTGeH72hnmoItWAaMgSPF+tV/oQ1RE2qPB+4P
81j0IWh/gw+r38UjUrDe0zJtY51kQnaN/PZaMb9KgfKdJ93exvN5D8eXWVC7HQM6
6Git1W6SNADsUeZFBVQGR+ia7ZRgJ7jsjAtiMy/+e/TKuRWfAaG9y5YURmoU5IjJ
T5xucD9Op200LGgTRHUti5R0mQ3G0WIVh4wM61uIolYgK/4/AgtEHAFZUF4P1jau
a+iuxx9uSFDlqQdaki3XIPI22Xi6zEgiKWmdHOuLLAjypxka9ZSeR+Nyu8RLcg5S
VPwLqeIrO20C3/jKmebDXhMzqaLr9nou09fmYBhhIROgyOAvWpx+ED6pcbDNWkZ9
oMbtFUvnniBoFIny0tteUgzR/Np1xqDmrHKHJ5GfJW1FlOY/S1z5KW00NAK9yfIe
+XKNHzwZrZzGqjRjzfrE+RcAxttpjOgRbkSMxaUxc3o909zb2H/JpECTgFyZ9sa+
rKaolwy1JIQl40fZy+BJazzN4hJ0Tr048ZqyDzA8rX/sALsM5HKFpnLoO9mnbp1L
yTSOVPigG4BWk7MmpOl0KP0B7a/6NmqF4Ov4itvyK6RVhOxhcqd2FBDRZdgN+vvL
Q3H8u+yxvLfbMWmaFPQjvRo5YJ8UJKFPUWpT5E7UZFJuofI/CeH818mYT/btd0Xu
gY6nPtZRptt4qSlb1yn1bUbtTS0Dqe7xowMnfyhNvKDLTGgwc83FuMUQMPcMMgel
LCwzWdM9EFrUanoPnoXc1FyZx8hjBsML5cS3+YHcH4mgaNHQ9Yy24ASE6Zwl90HU
PO9DhikWIxKZ/LvT0/kkK+8mvi/WVKLODBVLbZ9J0HEgwKqbE6kSjsAH9qWcg4pc
VWhb8BAVQtxpNMfYS/1WNyh0uqGnHqsuiHeMmLQq/uxGriLcyJ3DGbGJbZS5TgKM
vpeYv9GQ1qyUn/5yeQFN6kX1QPmS+GaYaQVVN31WdD0qaMiTPMLNZWlxvXwODsVu
ttyezNIC3JuVm3lPTpPEe4Y/nN2KWDP8SE7Ppu3paX/wuUuHhdirEhQn6gBshx/v
puIyEmOxLM/jTqcpzZg8WR94zcYrYHHcvU39ShMqJAxhQaTalsJVe9hwWALkqzCI
7ACuVNH7L2X67ieL5Eid1BAhhSbmgfJcojL6VhxdnlvvNiix04Inr6T1EMaOwkRk
ZQTsKjO6hP3tnmu/4VvuoYOb9YIXKTRw11kYBYc5CZyXcpOlewyaulaXbbTX+eq6
3s0f59LbX0ZNUduW3R1sMOoOQb8jJcHwzbQDMokaf1N3FC/cP8/BDlwAXpuT/BlU
41wSZ++/nfqAHO1rb+C6g8jJcXHGFfXoZ4Y+aCimSxy0A1OulWc2ZyB+PaFU4MV9
QRcqOCKRtPqjBr7cfr154ZmJjQ72OS7Mg9O0ir2MqUES89E2x7smdpPdLs/1J0m6
2HFmtM6NNOgpvvjo7W+O7oR2US/7fXXNoKkloxtlC5HWt6IOHldHjkAZdg8Abzhr
q33/Kt/KQKZMrAzVwV3hh8dhLifVmmiduvtokgspH3uiPC9YCY/NZaGOLoi0X9ns
WjI2yVj5vXawAnq/7d+maYJLa1uj5BF6h4KpZ1yzi+hIiyEZsR0gHGi1azTAm6tN
h/fS70aK6TaoBZMeeUTH0yJllUXYh7nAiH7DQace4iYC5TFYqNPgHgQweXBiIy8L
Mfze9NYDB/J3qHa7QLbyxznt6uZttJift/dKbA9bHqPxNBfgiuCJKHakUB/VMtrI
/LMZ5PS6akdQOl+QrQ3AZ6kPsw6E6f2G0pb6T2bUU1i5jYhWG2riNM7/YUZ0RgtM
QNOS9zH6Ww5s7BVMx//NYBrjoP8xP2YOwPMF0Rcaz7v4POSy+a04Rbene4x8zQC7
Lm9Na4Ws567oUe8HChGWneAq/7M9TOwgLPuCX6kY4dkz558Xg6r1FFAaAe6It+9Q
9DS/62rckQlU0Y7NOsSfQ44Ajq6RNJTITjcBvDolrQkLtJhaBbeRFAA5H2nK+hcV
okkIusNeoUJckA/H/0zDpc/pYPscnjKpUycaiicPXCCl1Dz9JNim9ikQJQzJCbio
4v2FctaEwvenY9UKeHMsU0uSd9ZjYs9qP5KHgZOKG5084xLrJXnTJzNdeAsXRDT+
NAVODSFd3r3kmyK1iK2BGPMhNuyUxDHiHtIIG1951hGGAXWv8Nkj3H0yLjujmRSk
vQ304lMUzqSC9uAC2HFFeX4eY+oVAOnl6hMRrf7lCw3XoJZhKY6CsRN/bkJ3kqXd
/ivjW+QNt0EFXdMYuSYnHDVbr14cyqRxfUgkEU1M8T5faydxvyHvwSjishqpmUTH
vKuwYqhMYKbAi90gSUZRqru7+B7cKaaTAMMZ9cq4ntTUJLxIbFLLyBWndtbvY6sl
CQRb4V09ydfSVrcMkUsbE6hCvG75fA7WFxCW5mJV97LmmRe+S7pemlRU8na1DNHt
H4Szg/H5LqIJlGfSRzgo8sjsZxtUJC6+sYey/hOptbisLj38Fx0aIJVmCza1nDj5
0Twjx+/xhK/vM6fNH4lE7QqyUGgEmiCYsPLNzO9OQcBLB0ZQoB9Vvj1HoX7Bz8Hs
BUxmuLr0IJ5HP9EinoTUhmp4kTGrY1vkzsaGY9v1F8enjFZlaa67UkXG5yfryzLC
SWBmY6sqS4X7q23ESCc9B8TiBwnjwVk8eEdI3JCTkTQkeHuRkVTlzalZpdRtPJIo
VeVKw8hr5mgEzLETx6OkLYA9qXj4j4UBO5RrzvY7SY4lnHpxDq/2tE2876R9mIUu
ck8FIyuPI8h8IBRHUT4cEMwu0lFlp/0r0xipuQ7D+MHowiBBTD/K9pal718/Gkto
3IEv1JoUScoYOhpGchpM3+ZMWZuwipl4NEmt892BbbSsd2OGli1I+fOLGRclme8G
IvR/NVixyHmcntlLjN8+z7RICFVFm+9+lzvSNvCqjUsUFW4/oC2SY41IY2KocSLq
/JDa0K9SRNy4C/FOzuBKWDNM49mO8owz+yX2/vCjdzBJwguPisOXsO8qTtxi+I9+
MB3WsUsqKoEKDySmfX8oWIKbVQhkvZNc7nmwtAFqFpcxGHYh+wF90noM/MOGcy1Z
FsB17OkEwMaP7DmhZZSvnR31e0wGqv2HDdI4bheA5AD5Ded0jbgWW/pj2CqnWGpp
1ihr8EQaeJQMVj+gCOK1wwx3MbpNOw+r/3wZz7bo8NelirPNHLHyIHwC7RTkf1CG
+VAcCsly/v/diD/bvX4tW7ZM2YCbpsoK3syjhkGQv6HrxWOh0cCH765KukxPSVpr
3Y25t47rRX6Nb77khLZo++9yaxqCtqoFGfMt1zlugc+P4RGyeJNmw4ieOVJNHZfc
EhHkK/eLmhEa5T0tQWtkpQpzvP40F5Hv5Iws/JVl1UbLWGR8EGoddacjRLgQGWtj
kXQ8Z7enZOFg+cGPkDEJH2prX9NmBcYWBpTBiB1Awi/UixSxerIKzVhYbmIrgKkF
1TlayEWCwFsEeAQ+dAsgKMyn/ucR+CSmRJMhfB9+loAgOXCd5oLBKOdm5OEY2TRq
B1JvgKUkQKWOpEX49I07SIMNMQyGGEH35s9yBZxaMVf19evJcPaHDOz0Wc0VOaUC
oH1a6Tbx60NdRcVydDQ9V++HqpbG7s3XmT0+SyKUBudIc8UiiVIXKWRqUzIhfsln
njfcU8eSvNy4HVhNkBPBKUidLHGTx9xUr3s161NaWkHvryhSn/WuR+fmaAJKCUd9
EADbfprD1Nqy9DBRenGmTtcEFtrYYtDTatHBRo4n4scQRgE1IRcLtG51OP1moUG0
2UAdor53BBd4yZ2XX5M7035048wj6fECJ2I4M4CEHR7cJc22lfrOZCG5qpzh0Phe
DoQ3DAf+meEKyiXQv4VOXaPDrmU7L6C8BIC2aclaI3V1iO8CdOjdPP2q5kchDENN
uQPn+4E5rUz9UT3G/eVp73G0V7qIDOh5d92GPDLekvm7JFEEKa/7T+6Hx1t6UdWv
VGP6Ze6RHP7aAYIT7Q7Wzu+J80T0La04U2DWcfums69AzK8FxPmZdeFG5j1zPhmd
ErDpDhM7lkBQnUbbGTWa/Lr2Hen3FMYN4MvBuH7UXzf7fw+WpTbSQuPPYr27Co48
zYu0F3YBzsOT8gzGaOIZVZjtzH7WTgbJEEvq8UmLDxT1FQaE0RND/eJa+Ej5w/He
Ph2W7X+tZmT31caOXmnT5ZOddff2OQQ4OBzrLj1R9iBC7qdGtgzL3N5/vHU/vY8d
IP13VNdNKqACGoVXPw+ENKytgAqiYYhpKhKxr12gskmg8Iq6/2Mk4RPrQsHXjV+m
rF8PL9aNNi8dAEpDDTXayhK8wesDHffOmVanWlGsHer0ZQD2D4HjiELaV/3YpSEd
q0hDcdboI+6LDx+LV5QIXA7/+Sp4uzEeXP3ubWT2r0QI1dVCmEH3Ct4t5DwHbCRb
/t7iaIS+02ileOxYLMFiNNjLy4CkPBoUReUZPitrEqg57a+mgWQaE+5sqD2Is6Gq
ZT8cO+ntaGe/mJUpknH8s8AxcOkvp9I/pAeLMQIn1KfUw7VmZNi55+n1xqYBmRv5
zBgkjIh+7W4Nt3qUtZ10u4YpdsVdzny3jwIJggYp++N4qgT4uLtkOZd8mBzxpISf
71BBdkVDz0MPMVA6Q7F8XsRtwrMwTND9g7kA9iW7ZXAU/TMohBK6a06tlY3lBdC2
o4hjxH4cV4/7Urj/MU2ilOR1Wq7j/ThXoIQNfxAjJAhBWGPQ0ZghW6U5Fey+2DJI
4xrloyQBNdRXQG7OyYy7KaKBcAub3RZqwLzIUq9qxlDPV7WonJgKKrT9cNU2VhPk
+XrxWnfI4nl9lFKYrcmMxtHWcX7Qf+TUd6KbdwPgSI4R4NCg+3xgzynyX8mSaIbN
LSrAfI563/VM7olAqfgI1qYbFNJ29veLEZNq9u+FTDV3aqnx/f4sTLzKpJGcUC+r
hhtLd9xijfKG9VCdUfcelTlNsqR3sMBYuPtMyz50tQdQq9juD4WAaKZBU+ENq7i9
ojC64VlUkkw2ZY1XKuAmoBiorIZDegvBcM4l2kF95ibj1JZthYTeF7EEgQQcwTZW
Mr/WbMi+74obOSxzhpzt8VuyL/kaJi8JT3Pv289dppFT2M/Vu0YBKrvnNTpMw7i+
uyKOd+j9SVTC5Q+R4W/Ljv5WuSn75NFisyuSGsDM+2SVHpJc6U7TmglmWZnAqG4E
bAdXcZBfprouxfnd70nRkKz5Zrrtp3Vtbh6OE5Zm5fDV9dr3kujGKo4px6HdIouw
mm9b4gWmC75nfHZ6VAKPa5Mmn+rGNDVtuB/MINgzOP3y8hy2Xb68mkSsYBisfj/A
oapWeVaTaUF8NSfa48Et61VzYwqVp6otuDtL2zDmvMitE0KsJ0uQXxMCDGD3BzBk
LE748aJD3kuvc/d1dY+gT8sD/hIEXqsGyySFuk4YzdgCJyjaDBoYO98HC1PfoxNk
DDheKbp1GgdOF4I6Obm9eWXs6+x/CLK4JJYRCjJKyJxPjynovFwHmF7uBtfQRa9T
MfmhtBHNeJ3Ws8YV308t+IXkUIImky0rujRW9pq0x5heajp4uzXZrKkDu4nMphee
RRnOj+N8rZgPHL/rqs91P247fchXrzid0f0gSqyt7u1BhAHOCRZrB8U1ajI6f6O+
O3PqlgseGL5+mWV+gPR1s+3NzaGlw8ICMA3l6XcZaHO62mZhg2IlmJvSQElAog0o
P5dby2N6BJqLzzwiaDDQjCyzGVWJIjtz8GOovEMlf4My3Vh7JS/iL4O1t9FGR7fF
eAEahN4OUB4YszYFsFx0CXIYDuQ6+XSkb0TWhsAzToIZJcqp2xLshu0puY3rpJAA
Ci6jWSra7vO76m9TQv8dXMiqH0sHHTRrXvRE1II8mCS2Z8ZIk3JjfBAydBOScfQm
WMjkiZJcJswqL6rjQgfvzgXt5qvZ0pYv3GkCTTN11dXN8p9lGBbMrkTV6khKeDBJ
1ctmtcvdPkkohyROIV0TTW0s19sF0k5VT+8EglFLxPKQ4fv+baeAMEhJ8+WmfU5m
x4oMBZ06O/4Stfty0gWNUmKkWO6qTa2HuSB9++ob900fMrPfvi7u+w9urwfz1IvC
x2pP7hRbrom4w8lQL9ScnRkDJ8+tf2E0YdEzI6tdnRIyFRptnsfzUHIUlqquAC56
bvinERKuuC6HFArSXXEqKrWGga9gy6yq6eH2LKPf/r+qCggN2bHjIh1QuZ1sfqGx
zUPHR2RifwZtYAlkHnFwSgfNDRhQk7SA4jz6myBQ0x4a+l2OSlvhiwtF63GViyzR
DggGBEwBcpBD0h5CjUF1Pcev3aiXGJ1Slyl1NvDn5uL8VVt63MLAZml3pypdhuDB
fHVUR0+ZwJPqHP4hOAZV3kVdpbOIhThQTT28P2LCue7vqt5p8nNaRrc1/tgW5eYV
bWPPNIFeotRfd+2WhsAMjEtzY0gOai9wQQOaDmVE0vEIJ6i5Yo2OIrWgSsrp2Inn
vkVebRsarnHhk9dY1mqZmuAjqw9LbKaDHgL4dY4UUrO05wTnQ+QSmnJ8UIHl++V6
BUJ9HSnBM0IejHw602XC0DOkFomxRhKE3+2p/Is6M26Hq8UHv0y6lgy/90A0P0rM
YRg39h5YVp/QVuGFBSbuadDQR1ifAjwFTgoRrs1nR/FNLdKMyka2Q5rKtaT6KXKm
RGgeOQ0RyoejWT4iPpjeAa2hpfb96o7DGobdUZRQ3SFUxgfzs81eOMiBUawckviL
acS/k615+YgP/WNzoYyAIiiX8LweOjzKGwjzKtlX+4M5NGJMKwTW3wum9oNXn/iW
KbwTv527/hMrneHRaxr9uO/uJ+DVeiIjRuJ3PCkKMPDK6mNIq2VoS5NCGINtgsBv
8/N4/UckeADXRadrB1W/H8UdTqgmtfNA3MO/1i9JyDUIAohQr5KQ8DjqNgnGUShv
arFAaAG9ZGjHh/8HgP9mRRKS8RCtR9wsk7t34Ckqvq58j0usIeyDH9cROM34W4MU
Z9CT1dx/aOxnq/kogaM5M/UMjr0rCj70KNEMSmMCU6AEe2BK5o2tgdOu9mWYYTTO
9a1t0j/1CzchHVWAtD6j41sV0H07FEiNgYGfumutM76qZPBapbiyvYBjT2mYAhqV
vudrY4NS9da6V6nyDkil6XGyXjL7ODEKBNrfXTc2vRGufyHehMkQ48tI2BJ2aIAC
440UwBxHhccAusjX+f3E74IU1EU9JMvYcY//iQg+MCaO7Pgg8v78ozVPbSGtnu20
nPoLpWj4S4ykWTd+PTmBxjQH1fd24UOnuOz9UEZfejNF4okfVfYMe41kijxBjLq/
zAZ0GwC0FHQqa8PS6dPznL9nGwhKHUYHTE2cjPoxmu88pqsiSEhQAFlwLHfDozBR
+T7w2339EIbvoq56ex4q5R04DWObpl3pzS/EEUgbU6kavEI+Jzd/63A7FsC16EvM
Ms5zn6imxVTsoh3+nXBqX8/lUDHy8foHbV7DNG6HJJBbvrUEv4LWON5ZJowz0WpQ
pIoACoTqTpBpX6azf120iuv2D8VbcZnclPSKbArQd3gCmfy6Acby7GxBMfO3Ir7t
7rZokYlMs2AR2RengYjGtXswr4ikbyOPR3w7J7zy551V2QcJQ6giq6RKWvFmE46d
bItxdVbr2L2tZrJ5nXbx8bHCD7KNbXSm4tLAv5UhEAG1HSvfwyk0gT6a099LKz7M
gLf/QEoQYuEDpmMaxuFl2gt/m/VoUdKi8g31mOTp2hIaEKLrMlg/JicovCXNNCKD
6yYLu7Q2+K6olGg1Ay0bKeRvv3a353Ch3WS+50+Y6yg3TPpbaobgnSuP+dRd7jGu
JuyFN9BnqeRop2pgroBOQwe3L6s3gjcGM1I8KMYBvYFrD6V7kkzVPU9NKqRibMiD
wGl+LqxRDG60Oe3ZGhJex5Abze+pFDUDERN0C7rCgkHbCzRoiYsDp35H55m+oCHm
tkKICIy1k0OPkPWk1loIT56tGqt4DLXOREWh9BsPcNTw3u1e3s4HWxXxMncGxEmU
287y4X1Mig9Y3GptLQ939qERRoxZBp23SSgv5fMtx56WjEnlgcpzBLmhM5NaUaxb
KSdzj1lWaXYMYhXSOf46IY7JxuAHa+AoeQNImWZfs34m7NK6AUkE3jfxCrX+nAaT
XA5iJzEiMw9WpwGJ5PR9bvERyrh6m8tNbhLj6IPgpPwUcYo8DP5+o9ea0IdiBZ1E
KwUaxr7JXtROp6SYdayS2rtZp+7b0Ic7/m/gASuHnk0PBslJOQt6VxRPC32bHKMJ
9wBMXcC8C80EkqwlWOCCHctfCYksNwuh3xNBnWK62+5OpOhz7FWTy+A5VN77I+bA
/ID9C1RiytQJfdHHIvzjPAFjBKzDWQpG9RiIKzjggbbD0uK0gxl1rVcWCzcyOR65
zgO4nR1QVmoUU5A0mhN1G2iM8T+U7A6eRVskv++N5ByMJNIE8EfCUJ5NDbIAg6+Z
F7xIpGHZkgDVOE4nWh8SJfsCkD2WPsy8hfuF99RDuYfTW6e9qj+SOVdA+IXCzcNI
TCSqbtkIYvRGrOQHfmDXzUdUoFRhgQByVC4oNjv8czkMjyJWa9udEEaexh/NZazE
noS9AOyaebtyrTFIsOpj1RqmlQ5AHRDIXFsM3s0+zmLVo6GQx+5qf/p6nz2xlxQf
qlMBfRtIdvaLGOGbdIv1w6TsR6uORWhAXF9rntMffpiISyYM3pSC9lC4GbBcryTh
jQO5kyfSfRYlLxyTINDJD/OHkMgcJ14WSQHISVvHI25Ne77lIIu3RKwf6CUIXROd
NogvCRKopT2VRlnoGBus1EkKD2Tan6aOBUW9e4Q8r9jaW+ILuOsnXiDs9f4THgVD
GCHUQtOnSdOpE3KbrVw6B6dPMcGMQURtiVkkEuKWejevfMXs186bYTjhBL13c685
TOnGxPvfYuFyIwFxPVE+N75oIkS3FTrg2hZgJf7mR1w5Kw/WLEmRoTxOeB94NdZm
Mk6CqvYxWZBfeuF8i71dyItBm7CC8ykqFShdUGsQGAwlCXuKEN2Oy69WZi5X8SA9
/a43v4SgPq+2cCP0BgywjZH/LsQTXVbOzBzQdOI0C9OOsRQwA/8R9vP0P3HSTplY
A/7vjA2Kbva+AqQ4jKKDmh0TmKl2tTWGt4jW/apCp6kVZi92+moFZfZp2t3wOOGK
DV544ZULgObtxR/B0m7K08lt7S/6UhVPQTqEJGnJqhI7hG2khICAmv3+F8LHhana
D2EeWhhXuNG0A1NADPe2aSv28CHrxNKsUpY/2W06WzNFPpEYxDLfl0FFkOVLXKvv
yBmHsUQMm27juCIqhlvwBMWkJWfZKx8N3Xo1LgA9BLjq32plbVlEzjBQ5Udl5+qS
OlMJvLoEUl6QL/XjqaaZdDj5glJToxOfW/c8TJQsgIuf24qCGBYH8/huk4mGOyBP
y2hZO8hnPD8NnonXbagCttg7w23WKYX2uOZPLew8uBe01RmwLWRObQh/mS3QIliL
MMitu/QQg7D85PpagNe6QZCIHoer20QXUKQ1QNCZvnON+LDiMpkszorEJumzXkIB
oXP2FTmr8nhH8xE5OHCElWW5f4v5D1+kGsTq5t1HyBSP0+9TuhZwFANGK2uAsdfr
3dekG5Olz2K5FIuAYl3f/tDczULFP84UUrIGT4bEJcoxG3OJ4dtNVIBcnhb2LYAw
pMEVTqAquk8h322xefxqWb3rCwqMOAort3muUknEm8sx1dWcRSS9ad8g12rpdfD/
MQdKinC9K4pPui49mcE+/hU0OhHcLMSGPEnj3YeyoUIgox/f3z348C5UBDKYEywP
wbIDGsPwKPTok1rLA5h2DiHDpzob4KhT+hlohzWhZ+pr9yhlUyXZF3/xu6OLkGxh
pH0IYV0HULEJoDR3am9ejeaPnN+kKOwvUNr6N5ucZ0z3eTtrgZMHg7SHpDp9pv0d
3xgQgDL1T0cXzcsCNte9Z2e8/nxA4emsSPhbMsAcDBnobuK4AP81U9dKq41PJqZ5
GgbFlM6uXx/MnM/3hHhSTmzGvPst+TbSnWEK0yL934DZy8PWh/PoqRG5HiTsYnsc
2tB5zy4oQpY7CQhRNMgANnOk8UyG2hCYuWRIRTtH3EVlO7U3R+LC1jR7RxhXHNiF
8sk+4BaajSoy1p3qLjW0Bknz58s1jb77hl+4FVZG3zzU7nPMQJMij2kz8Z0Qo9Re
neh3Wzd5kXbzjk/KnlrSTk4qT0XXHL7y8pZ4eiiOra6vA6DMIClLtd3H3gF2heqw
xWYLp1He5/EUy6dR5VwIvXcGADOI64V1Wh9PrUywrvJMSad+CfYvuD0ZkEjGigoA
PHJ7Zx/9vqrb8b+VTwBUN4AMUqoJu/+3ROl8ZwzbCjfUqlAzrD7llPVNgyjRSAGs
+lCh4t2/EnIMQOle8RWibNmL3oxjFPo4Au/vrR75CvOHJ82g1aen54T8NzrnOLmr
knMv1iLMqSGScEq1xeN9g+WVaRguj2Ry8auH69AEUJpHCpISJ+e+qLOCNzy8LXtW
TTtbjpK725hYTsG2go9WC5Y2WN86AbZ4GTOE1KaoyjfUPPMvxGKX64noLv2SvINw
/4AEYJXqt4sVKPQLEfY+TDYk3UlxqLoIBGD3Bm9tMJ8ZijAffeCcmaqMqYCFLllU
A3ki+WLK93wyjN+O0dvDpgBnI1XFX7xIDzNaq9cfMnCtvTiViiAQTcdsaLgU7Kag
5YVn+6CdboONl3B+2/qrOj1QAWyuMBF5bt1O56jH7gynorIznQCbFkVgFaX4iXZ0
pjzP/lyGpfmdxwbywf/TQWZb7GXQ77EQphwFO2WaM7A+kQ6mvWCss5RiHrYsW69I
5nvTiatKOLsyfUkjzqpjaId81W2tPsE7EZ7UwSONJAoIcMc14nleHJlKNbbdiPNb
EDHXvianqr4EKkRsCElwugUINGermgbyjNNwBE0Aazji6HmXLuK2sxjJ9p4HVJue
TxgkA8pY9Ib/seuxNRHgnHFZXF+uBGbaFl37m+ujNZcYXoUM3TeJ+aEKrd4WX67z
3mQ23T+CnLQvbzBAs1Z9Grvfaqi48eNUlewK4o+YsfSVCUKigxs5G7uPjAOhpl0s
i7EXF49YcO2o/G1a8/T/K23aDqhopqaqLRyTUUNSeKwksbBNMtJCLb1cy8fk86nW
quR2+S8BIp41jGFsnJkgIKqHE8mmzmby3rennUiVxAEg03Qap9pvnFjV9E0v4xV7
bJSnBDy3dfKvDOiL+UbIJM/tcSf4Q6lkQUUuc+20O2csq8xY0AtJFljCURizym2V
+O7w+0LbMoRB9STEtMIVOqQZGEJ+5nvW+ahZSltZpILJ3eNj8RnTBhv0J43JEGsw
1c4Whm3QnDN4yTRzSg2nh+cyw9EN/ENYKzOsR0hvZMN1joX7h72VlXH0Tmg4S87p
zso8lAjUsy5GvmXJilvvwMBQLoTnMOuqIckw7WbICWIm6R0NPt7HAcVcQ/GB8JAI
iZpLoLNV+6JP/6RCG2lteN2RPkczcVrPD2UsGB6MDdmCtVdPCNxVZqU0sZPIXecx
/VPuwEKbxc8AENcKszgGSnHS1bzMcN3kKnCu8VhZ9qBql4noI4Q5ch1ttODhhFA9
ifPayuuDcvs3aSGzxevgZwoEp7z3L4LP6eOMQ5hz7PwRh5GPmfvVA6GuxTZeEtuP
lyTj5EVDuqOJBd5qTRSb40zqA6GRrUAC5eeiwm11ARiBILvqEKm+QSAEmGkA6Vpe
s7rXn5rgPNoRcl2W92u6lL7ZU1vEHS3Llunq0iBQ3IdTeeCJoMVBewqKBlzLh9r1
umVUkVyufAc7dGfZx3HWnzEnXrl3cdXphuHnT0xF91yhBvLv2mbYF0aCRq2E7c3n
1DhXy6euwMPqApVm00/7EWCpe5IBYCBLDbV9GNCNbLud6SXeph2A5k+CU1qQEO+m
Ec536aPzwx04LY7pfTZT5R+TW0BTfMHL0zhEDp2nxfjtpqU7ku5UF7/YVjB4gOQj
1foDz6n82FxdyRkiaotu7A60/gibtrqBsXKNUnwK9zEbe/v1W9xT6ULQ9XtetrR+
VEflgIUt6n5ubbP97yVXR+9eK/YDzOYMce0sjZpftLbl6uu2XyQLRBrUxn7hqSqr
9TfkSyDKoeMEWZIxDoZOn428PdhZ4/bFKlBpsQJkAAjYoXtjMnhOZ92gQYVDc1T0
JdokyG0CJZbotpj76Mv1/FSPt7Dn4QW6ehkILnX9b9Xsl9VT7BT6HabMXS+p++jg
tT07pRom1mkS0WEJ1kC8fO1VVtWO809GihclBjebySgMv9Po6RT7Kwg5phM0QDj5
eMKnK9pHc7NpWlYS7XnKYgPpFecvos4oulcJtmUCSxSCiRxtiiaYCOIkBKDdgENj
BzpXJ8AmsV/a32f0Uv6t2cqg9vYTy+eri0laDhDhnPe5EhUNSB52l4l2BIta9QuQ
5QUPA53pfcsL4WqrhEQ+A1SZ0d/4wEwj2eRb9zCFU6/KTG3r+4F2PAB+O3PK5QIL
ymMoJGQpbY47XKKfZ6V9bSjjBSAZ8j3jCKxBh4N41eenDSQzYRdV3PvwhlixPN5g
lWm6Pm/mmU+OZP1qld/p5VSXB6jAZWP8mfZfF/WJ3v19vdFBHF1LOV8mplA+pxu6
SL3rO7Y02Ai8HsrgRDw4rMG+9ofIy5xhEc8WZEHHg0NhFsCukYs63w8c5tcNRIU1
9KhMjvRq5B3V1VXs11gw9jCxczDFYpbtEuKCbRbR66bphFi7q/kRJtZSmsKzo9f7
rSkQ5kLN//p3Abiy2+l661X7PruTn3GtBfnlmU82gcREBdqlbOUzow0zLGyfRSeC
7KdpMN8JrlIqKzvPpKeRiR4Q9XlwDX2E8FRrzTAQSREyJy6ZZzPmaIDQ1Ukl1s5p
Lj1EvCZflixTV+TArXF5GAMMaGE4fwYH4HGfg4Vhg5tVniLTnxUNv6wW8oBG3cCP
dBZzVbn1tdW79l1NJkYNuzXqRkBY1ch5k1GNFMPe+hG6PF7bO4IrBy0O96PN9+OG
rhMFIPy7umZEpA/NCBldiUUqn63iU6mOsgElvDdI74jt/pLegz4nfKRWnD4BZinW
FRuipFHA6kbYLrhxNhVxmllrbYiwi6A1QYF8+yuB3Ewps3k3eeD/NBBiosz6FP35
OSkf2UgNd/yi9WgX/zc6g7EfmgmS/OiAbf3fF6n24jw62EdMjGPa13oQ421fjpg3
7bRIkIKqGjat5IBOG02PmS1cydJodnVnvlxF1dONXFIFRuuGyL8ltkcVPvywVClb
iRQHTK49Yr4Hh2lBq4WMZq4uSqTxy7QPeK2I5C2FJurwJKcyIK0ox1BRjC7QWU36
/ZnmWVZK7GO5lgHEXyy5Na+/Rbsqq4+6+1yUcgYuI0Z21aeWBhLnPzXzTwdXvF3O
bJ8fJrbQXTpf5plG17caqBVLLnD8Bn5ROtQnP1lY5oLKTXy4ABLNUmWEh8faAtBS
MB0+sN2r/IV1QoA36vb9uEuqsS3BLinu96x79/DA0NtiZEgJBkL34/DQwqMUk4AH
8IUcgvlMcgiPFyxX1qHfLz/F2KZH9ImnYi99tv5/22V7BjKiPE2jfaaBAfxVEFGd
gd1Qo329iwSD3j12xI9QaQ4hd381T3DB6CrzE+2Li3zgMP+zQHQAcmioZcZPQDTG
sWjBKNj4mpLpRVNGLazSln4pTYhM97hVwNEPzXbjBlb/27OW5Uewlz9+6JxlaSEx
8gkOclhv7OkN81h7eF31JMYnOQoFK4ESggO63gETnXI00Ujgqw6w1IEiZQ7VTg4Z
4j7NVY6xcBLT1PMEDoOlNsZTBu2+hmZEoHECI642wwxW/NbHFJ6Zhk2NrA6lmWIU
yKnqZuOgXVIOdsxf2hy/F1P1L9iPqR4m9zjDI1SEFeMYRqpwhu+MmqCkyNnLW4CY
VVNYpq/1MFqOA/61t+VOCwLyfASTOn0whdai9dBj+DdZX14UORpghy3/YmfFjWYS
rY0iL5pdrBlQXN5e7Rcs+vEKfvER7l0vxOjXDKsLRB1YUqzUsMK6g1nbR4r+vF/I
1XGuKXnOQ99DNs5lUwf8X/E+eFC7uUHnRws80HW5QuVgJl/MIhVdhlRpP3OpD9ve
+Qhsa2Z9UQ1GUSSncA1DY/eIBp4cyEP7ck9fCDUr25x3db+rXAq9UiURTTd7Zej2
nUbq5/1UVlWWBkK8wUo1nbpFpkZu0lfw6BbQGdNWMbhqMHzNqeZGjNN91GTM5Hea
bUb7j8jRIeZOnqVsyyqAbKuVYEwupbElAe1WluKQ73BTyTb/pEOoYsuwd9Fx4isP
HnvGiryOML3Dmgv95zuPs/nYS7oDurIiAj4Px12NFis5Alz1kDwa9gOGJcbEXhD3
hvpv93QnytoA13Kuxre8toPPds64pXlTYyF9OIvUWnC6ntYyNpOuAcM3t/5PYZCM
wa7qTwzSoqhPGaMvTisGuA0M7raLy5VZjoQmp7GGcAz3UfR10mban0xPAV4f+1xF
VpdRLXIuusniNroofRCx2J9ydEsc1DzAcMfmaraSXY1r5NS7i9osQWCCLXb8pQkG
ucn7rcNUc+NBjPm37su7SBrsQQbDV3LeAnk/ZxuaaMIOt7zyBGm580mphudludzZ
Ia11xArOuKgKobtRALAs0I7bOQ6CMejwV8X4SDZ3Wns5KosM3djT+8Z8LhLr7EwL
fswsDvzPUXmaFctvOJKWfTGXQy+GIBYu9qziiRshgWu2fwsZ+Y7Acs5tZra52e+3
wFsm36cIr/jWQZx+uWEE1GFK8LAcp8UmXRc4nYMzhxWaEVOpkHsIpHIVcrnVQLqq
VXsl4I6fgJdS54+ZTWFU+lEe3N8XrsMCrXdwhoWpUlfigZzPYSpStPUykcEZ1XmG
zOckr65L1pDxNJ8FTcR30eybLunX+HylU6+TmuNUuy9mj3XDDIRQzcndNTM9/lB0
4naOFE0LFYnHJzI/ECmGajgMKOJaCvj6GqDdR0XGFplkK8oU1DWZTpoct8MaBHjR
1HCgK+h4NY37tFG+k89/IX9i6pDbn5j64CqmoGmhjfP4w/fX04z0yigusXTquUsV
cHHJeCZ4pmoDJ8vbb+R/umTRCufdgMrmDAXIDx7P9RMv7JCbRrCIhbP0HC4cvK1n
ciA12uowVV6DMuPhkOo0ZO/FHGmgBRLADH0nLRcyRkfdL61+FWm0GncSa0BRM2kY
qNkUUM3XxlJiJfyDxAgQ8CH2Pk9oy3/nVeEybD9hUJnCjS7Aod3RjAJc/rSPdXiy
eoQfeqz1ep7ff9YVomKJS9sF1sNZAHwKfU4HXx1TpxFfvfdbDfj0jKFsvHC+1Wmr
H4q12wmCR0Xjw/+XHihu1VMr6AsDBwMz9fAMB0Og7W0nCYtABLsblMNruTCV9aoe
9W9z5DXdmTGenAg0T/e1zFjCcpqT0fqYjgctRB+mm6fj6BFwnSng2w8XIf1cz7Fg
iwC3F/CVFW4181J8CFsUGUFytsYAc88toUh9Re9ri52Ps2sQr5hxb/WGWh6XN4Sg
nZqJTiY7tlBCrxi4FQ0Y1+WAjIpSmc7d4k/HFmX3gFdSbqIKz8MtUBMTPcN04MSY
14j+a75lPEcsafNy4rTBYzPuZcWRS5kZ0RnJiPccdti482CQEVLu+QMnd4XM3EIO
KTx2yM3mnDnJ87K3JtvUiGbAq4n1bkiaNZtTFgyvcMXdbEUqM4MbNYTqGBUZ7vXh
rK59qKrfv0nGZ8SPFjol73SQzsNOry4bL9Hv4ojz9BvbdxnzSJruI8/i+JgudyT/
umShOXkDpVE/VwNfRYuM/S11351SMJkqQrk7S1dhLWwqWrzGl8zXLMewhnmL6dcV
6GLfFzZXQmz+4uoDpBwycj97oImv4pMpici8glY2TH4Oh2j0zmxZKQyzO4nx6NSu
Jm2R4xfHgWbFrD52l1J91R1d0VANYDmJ0K5tLJkkO54oJGV9p+6B6xb9OuZB3JwL
Mx95B+jJNteNht0Yg8tfNWdgHrRLKyJtnlnpcyjRu8HVaoNTCByNq16isUbQ1VtI
iZuFUHn91ETpnvmlW0k9jDfxueQiB+ia4R2/kQhBplApxhTiWWcBOPB88fRmtJS5
celArMC2E6oKia7Forc2bodS09ZJtKWrxlnMDMLBudJ0idaPREggpfoS28wHBH5s
NHgq1vvVZvk0ZRG/QGG7gio0W8/0ZyLAFtW0MHLatVyY2XZcg0eztDT5b9ama68U
VV/+j9wHLHxfkBcODlWAb0Ywo2rjGU0wUWmqjueEtBqHFAukjAzTxVmQ/xBpMQWm
WXB9YbYFISCAokyV0IA4MhfSajO68N75OMoarE3VKS/0c/mSPJYbTvPcRBveorzQ
WqeHH3G008yPzSZIdsYC3kQVlzvUw1KFNmPZ24R4HjyGVqJe2/OjG0C6voi5w3FU
fWdHuTzB7u+rvDW68Zv/Vq3n8oU22Jox848FIsx9ckTbcFDT5gu0q3UYUrxx5ufh
YPwwz1iqhM3keuFVw54X+eYJvPI8+iShEMZo+pZdBGE51GQZyD5z5/75/+QOc6We
IzzXp56UhslRELJp6vxWjcmbYD0xF+8NuUCe16uBajUMaY/YxS8T4KwVz8P25hBX
0gwPHdT+Fcwd2RFevvYTumt0s+KfumUzYYLYR/qXeADrLRl+o3L0LGWzh9D5w6s/
dpLvZ7asJThc+yexeyxgJVpi8g1AvtRrTIxWbk2J73IszYJfNBm4mgd01gBfJHKd
Q3PTE9BLOK+Ao3jeB2VLdtXucdPw8SQ2h57AkWyO1BciK8HXd/M3oasHIbJt92BV
/Nm9yGqVzdmwLD6q1QIqQZSvRNz5P8bL+8bD8bLsKNJ0XcYq+yDMVZOqIssDrZeT
yPwtUKd8O5GTx1CkhpnDDt2Z/TLNS0c+oOc0fRHcLU9y/0UOAiiVLnat1JfSbwCP
UQmbSaQKmECZScdQL5RKpIKoDwgw3aIIES8S7P+/Mk5Jcs8JZhFQFt+HraLOTO8C
0G9CX1kDpkMGhuihq6nec6wK9bpxJpYc4I6KTTmG9dOt0NyOwf5YF5SJ6aeF3IBA
agxQo3cbOA/bv2+SwohpbVMerxTpAZFDjwKmcYPqiqNhWcoypCeITOrYYdcKvUzy
aW7fHtcAda6FRQ38Lj8Di34/avHV80uF06o2jO+NFaVJQKJVVHG/EehvzXrAMpFS
kI8tKeAyOeebQt1F8sK/4M2tvFkUj6K+4L4JpmmCWEVvZD0lh8Sy0+BWk7q26/+M
WMf80JLJocZybQVmWcDd0VWdf7FWgjQK+yA2PqB4cBuBUq+00H9Bkul3xBLi6H1G
autpJaShULYnsm90mM9zXJRgmv0/K31PI0ljQq4I2FtlNuCfDEPZ2wf226D4E7Uu
SqaO/9c9ulc0H2GoQDtM9OpBN2HV/LDLI9fhNzrPj2+O3eeUQ8iScQCKp7Lxywos
zEGKI0VMSRB555AABXqtovKHqp2cuhvRReRK1M2igy3s4losAWY9mgYrPP5VZs7d
UY/0OOZiECuxEWQpaozl9vfLvNVgjPiiRCfaFdYafCZ1ER1g6yjf9uDk3DzE8jwG
+9v9CHfdjdimn1gzd/9+pK83lQ4OnXu283hZEEgJlJiBoauI3tVbgpnWYe3Wtyao
v7sk+iKmH60gvoq/wrlNGg1XUdZteR70L0oVpRACsQASjpAGgBdGX6ali0xWVDxa
2tKLCaf0JSUSW1LtvXtD2D0/Fo7wCC+la1lBwRKZ2Xy3Da7UrQ0UtNo+vs1/0/tz
dBEp49RUia35xREB9dEe65pMfZmNFFItbBqF7t1xvT++/zlVKvew5JJDgFgJhGuK
D4z6ZQLvOPGw7VTXacVJpk2g6AG95xnqG0fid9FMoclMZGoaVIxEC/vJGndIfY5W
ZK1lvJPrCe2909jnJBryTyrwdlEwYUSho0ECt2SRggqKJRGq8lPw2xwHidxAXBN0
ik9aiv6J99ObO1y4MHHXjoXDvMmNzv13+hEvio2l00WHemyJPh01Z2i4msoyLbnM
whW1lRmBJrC4lUpcG1v5EBeVQjgIC/2WE5P17jmOuz4Iakim75poqo/b3zmKSSa3
Foj24Ci46ElVcbvFjZjJ9FFJLQRGKMo2L9DXnZF2Fajs8MaKqz7v8+9F4cmRt6sc
def9gYW3jWKhopE1HM6swygmJGDWvXnMT0fLWSooNpUEWj3dlKFBaQUlL2SMPbzt
AhA/BxNJ3YbmZ/az3V7PyDcDA6Zper1QjuHoPbuOmAPi0HqUxURLeD0ZdytBCiQj
J1/MtXqDUZMXQJ31iI1oSgyU7fR2EYgYHUsBdwTUG/SVMXal6fq+KhZ5IWYw1HZ0
lPxZSd3M7gLs4gBOPHbfA6bz2zKXD7u4KDYAGwEFPFbgShflfsVe9DuFhCe7R+ra
l36j3QpbRYNO6D48opTOSPPyD2fTSjjmjHWj0HXg08Xk3jyrPBNS10nu0gHll8nO
GZTkR6TNON/3zXOr+MNFBgQmjjNylarXNCF+2T/FQkitsTj0xISgcuC01yTO0i+T
i6QcrRizp9HLkk345w8U+Xb/6uLkXled2+QChvZbuZtdtyZ/hRYvGk3+sOGLeRVm
fcw1f87Ceek4uKmPTZvae/bkXhczecmwcnQMi0VyqowuOSYBxqAHdKKrF4Do8Ghe
O4Hw25R2F0y1YorO3IxsEvpnaax/XJPWf/90zVGRsgg5JWfb0aNKd+DPTfOKAA2N
zENyr84OrT9pafZ4yVsx92SbmAMKjDhWwOXiXm2FPzzN/eIn+MWxGHEsoigYHQUX
Q44V/BAoGQyOAXMrbdd7hulBIZWoxbknvbDgOyOHalyrfJ2VwSe4/Dxb0K/zEpgS
o2HoMDh56Lf4R1OFuZnMPki2Y33cpp/HAO1slCrQjwmxsx/gTP/Q2stsyQPtk6F5
w1Fw80j5RluA9vBH4GPUdxYOI1AGSzgzvPN5tBeP7sgDfTHVxwmxhrPZhw11jrQU
HD1vzesaBp1WVkPQwRhDBBuKYjlO2wBbRy+nakDdhz7jR5PvOCSb+gIrxQvjN7Mk
lJXp0M1BdEUxhQpInMJv7QHqaQ5rZqU4eYr7SgnNmWIj9uWzwDKdR5PgQi0uVpcD
/D17ahsIPgPkFx2df6dUzI6xqIHSnln+fd4/qpkKgkoYUeo4IKIEeTnBoO4JIZfm
TnL5wm62l0DH1X5U3tLgtEXPOi7mglxr1mm9lh/OlJx7CZX/idkK5ahe9E02YqXJ
3RM72EpgZvWwUnj0DjU4OpFZifu91CKyikz+oE2HMBrcHNA1GNLKknrFOISRMs+G
+irDRBluMKTMc+bpaiu50GDda6glYw7Cnb29kJH+V2b20z9QnIfUvJUc596Ttw3G
DfftsiiXpOIG+9/2AZOV9N5U5DbgRwGXwW065rcwS+seLKSOuoayaw3s+J83pv9o
HWGSqFFGVJF4HuXtX1WwH5DeOlLPv+PIj9qN1vflN5vXyZF4p2lnk+B/s6Zxbbc4
Gg48+vjOY0oT02U9+EWXHSElsXZa3ZT9kFtQ0D9ZO7xHmMLAbIAzAi8v7M23aupj
zm1kHVEysfPHFE9IVjyIYcAL8OIwkkfiXOV95PO0kKDDFRgOHu3OYx15taEtZ9Ba
v1laC4e562J+TCVcrM6llaXfEVyf7/TTkxllbYRNlpevo5dM6Ptqh63/nw4BvNn7
uVMA10lxtP928h2+awOT0h1GUpKE+Z1Ykq9azOLWPd9l8TEV1ipt6QK2W6+Wts7P
2nqNE9P+aeBCFSiOb/k7DUBbry5yrjVv9Yp1+xVSnK8vDpnBwTjJywjsrnZiSalA
RoA8j8Fdkdkge9h07HkGG5awyA7L8h7PZ/qRC32MxGHhgd2HC4O6zcAkxYEKVTKc
1ofO9s9qICANIVLZB2Fz6xwMdt+qzmW2BhPadtkNYDHIqG+/OBpcKD7KcqglxvJ1
2RJxbqAVmWN7YaYA8JrFIgdIpxWQ0mfdycC2vlZzjzK2gTwUAHGLGlXivJ2JczSE
AItWbY3rarGCtWm65ybCJeXOshU97w3rJ1bxQgLfNn4v1dJ4doAKjshOmHZn59bK
e9dx3cPYM/asrdDYbT97Tg4aWRGESrRigChC54MBbI5Uu2BQVPIol8Y4JUS8Xw4D
jlcff36BdPNMjp4/IzHs+bQqrclaEMe+tvrZJC8i0dZP8Lvd0iOlMhy1v5JVXAzE
+Ooutjia6gjK1KDI13ZRt3AzySQrM+jM8G1GY9hxAbN7t5AQYH5r68EGDXlTiX6x
mX12WlHOVVnrDih0lfpjCAEvvei0ORp5621eGTbLIsd6FiY6vULqlH2HZs7VQjSZ
zAObZkWk3dZr4PJColaVkYCfdNtjse9MUrDfNGBXqbJ+kPzgKiIu+6x8X319c7Wz
YGhaiq7x8eeJ/cpU2/QceDWA5zyOPXWVlYLiqg7NTTXhZXLkO454YZXM+ChXWMie
f+d+mfyayambdJQashKSpXD7DuCHWdE420LjSibRgKgX/Gt3vwGAvJEqaqOa89kx
HnVRk6ynTnSuM0S8MPnx1vjjhynuV7sPaAKsqLxYnlQ+9Av2Sm3UTe8EyjllMAU5
1Y11u1yNlgWJJkBUFXIzq6TmdsKjGRg/sIiFXk8Fx52Ulj/Pp0JhFhQ8lPqhcubH
fgtSKAtu/AxPfJov3luv2682dr4LV4uqoKw0VAxjz8pdhBJEcmTobqsIYS37rIvS
F/00aMF03IHPbv94CvekxyM4bx9wyKKS47eQQ8N/ALF0iJNLON561PZJJ6ttrOXY
4IEb7HcAb0z+RQtfA0xkLBcGFleCpNobvDzHjB0Bu4lHf17VmXRJgdSpqUy0ytTG
XoflCYhgMQUH56kTVLSCgtdExjOSmOO/26nELYcB5TDu8aW9y8lLoCc4hYXxx32Z
EypsRdfbpnTR4ikFEzUP7Ed0OjPUqlpjgoEBU6gaEyKHNGvFdH+zh3URYn8csjch
zJVydQELCM/LgvFlfklcLlbr72dMmq11DBtDwRFeiK5eEEW1os4k9KfPo9M0lAQj
Mnn0J0+2OuBjzMoUKirOOYkq5DQn3+x/Sttc3hJB/sWtJ6aWAPjdEBCFhCF4DCfj
1m6iKHjM5QKTOjFehSpeQO1znoY8llfYjZ1pjNnXNAYqSRS+f2ik/pzM4nPgsztq
v38NCG0jH0qoI3ERJpmFHIeZp8oA32vWvYENwEZ59g0WDAknkC2iFHvi1dZwmS7I
moveFdvmWnvfRUvSIe5asOXXPnjbyEDut7aisWhyAMXRzd4IIGVNaf1d7tbH+TvO
Ze12RmG+QuUlem+KW6Ldosny5dMZv5+Tz5jiCKxYTKY2h3o0bxAJvpSRqiu0+vPn
FpLRPJ9bV0oCVG8gKIIlvic9kk75dOICTbfbGvO3KKBGLGv5tQSYhxUOJSZmQz+g
VHXZSY4yjhYvrlQGdSITJiACc282dnM9+F6JRF18zpXUWMW3Cp0ib6/ly6WIxnHY
zWSo/cp1pxji5JYaCdscU8t58sdE7Xe4ER1Gqs/sawfxFhuz+y2pjR49Rpbna3JV
ez6gavrL1oTFfl0CSm7SjgSlq+KdHxHhePgydQ1nM6CwQC8nNGPDuwKbfGMCDvD3
gLBPVgrN61fRrufY9nsRmJJ6RFQ+PEKW7R2ih1no7wM64wbl/Yx/DX4roLeNtL4Y
N3P9MomRGxsEtB+WPMCkEzDYxGfL38owb58uHtOG7LtKlap1Qy7G7P7BIS+TWrcW
8cnkpMn+G6+8kwCgWIxvl1ij+bYYJ2lQ501aMZGilG2y5rX2pEo6pVcN5Pvq2PHJ
8UWk00for3TMJKYwJOHgj+xM2ng4FNIQJRAhEUwAdBlOZ/ZTDkWBA0Iy4SQ/Mlel
0ll29Se4ezmR51Y/JM8+iFZw7C7eUSWUvvAqk8cDtyxIxKTZ+XnXJ+3pQbgULTGr
BSus6J5fjzkWlSNU0wL5XgjEYfh0CfjmOlQPOnWLmFdPnst9wzJ6dJjM3hqw0LxV
BphYqTEf0m0wP0mfnrRtYppqu1Zp21w5WrIYexv6W71hCgGK1Wl461nJjzFoGIow
tGb3YJbmdeNc+8PreYS4Rg34U+2YwfNIhgziU1pww7caaSnDO7hJANMdnNdWWdiJ
CzXr/kG2TyaGyUrfGyKLbECTwDw2mb3CJW8GLXBAfQnfhc8yeeZVgP8V+TNrndYy
uaU6tGpjT3nNN1ALI9vYdu/m6hOxMpAWV2QSwLmduW8ijePUd1Ac506eFTqnOPET
RT4JPahoXG6Cpiy5xWHBopNPpn+iiSUdXEMAPg2gtREGIqQEk+Dq3eYLEraITpKs
kVutEaTW3nq+OcOC1aNOUeaHvUws7EV63rGHYGwiT20AXcZLMBPv+KQcDbCnyrjE
BOUGOJj1ofcranoDKe+f4G/sVJFpkc8rhm5NHNQNalAfJk1CFvJ57JCU/7iFFFNH
hgimW/YttwRd+T5vY/rFdPvbycrPhKL0ia4UPHhQ/TugvhVaQ5p/GsrQJfzLn8cY
Oa+rKYMl0h3ZvgXkifkvtD5TcLp3Lcr+3t6OTdpAToYJO55YDUWdn0dhbd4AlOLQ
VqVKeWbbVOC1fl/FOhxJUqM4asY5EseZjuPD86RSK8Pfq7RAtRXrMIcql6IZR84+
EmKB/6R+TScdlfnVATiowJ5pJzN5HO2lI5EjooiA8hTWHY9O2XGwPwv4nOSMEcZb
wYGKvzGExx6oAQfFXHmU7LVZYycP82vyVWCLyfy4kFJ3DC/2g9DboLltJoB4N93a
TXozlOBMep7EeeZSNa7TO6AWtxWdoTieJA4Q7rJ3dm/sooBpgX2uMnb7Ox9zBAh5
/C6dqie5rh+wrIHLD7QOW/UoZjzvGxc+c4Ur4Vvm89ftLzrj2n/ghYFpnZIPzUjA
V4db6G4AGnImJVJdQIKhOuSEStVT303zqCW7Djmg3qMpzGCJIHtJ2KOyuI7W4ST7
DR4EJwS9SHLQesaYORoowrOKFzivCu7lYjQtTZnyaqrmqnBv3fCuoK4K0YDb/53Q
DUz62PdT1UwjRHVc/O1nDadZBjMNeRCy8DCV9kiSv/I0htRzKOE4rLEqNfHDYd60
Zv9Z0YaV4ZhletEDu3AFl86lTBQWnZLD1ky4gHUOFiYobbDaxIAZGnGZmSREM7No
4xzWfyvaa7CCWjdgeCxZfe3AsyCr58KSGmlgjZDiNG7p4Krk0tLtLaohgW+8xMXt
WdF9h94jMxDPeUFFyjU7kqAFLi/7HtxiJLa/LlrUscFoIyk0svu7kl6XKmsfoRnc
RO1iMMTuQA7EfHSDZno9tEHJmYaMeHtTAWLiCCvHrWZ5urfHEC7M3p5qnIAkfS1r
WArRhcvXPUfV5yfGivdAhvkR0MpTJiARXMij0WEOJoib0jZVHQc+jW9IWRTPY/e2
4YI5JEGo8pOOWRaLTrfoE9tQD9Ic5KnRuyvNscTMHXlTMS58f2FhULPMHsQsJvvk
a7E23Qw9eoH3cPvXzxoyZL8U58lGnppwC6z0GwMgOoF3mDXc43szKloF4hQ+6jaX
F/qCgjl0d8BhCs91suiUW/Zj2haAUlJARcp2Mbd1rjzptyLjv5HS4pEEX7/Tm7BB
ZWA7FM+QxVcdXC2QvHAC0yXKXrk3QSuqODP4L4e3QGDkFud/snfWdonOOAhl1adu
FM5Y9zWy6tDH9rtleGCqVYl7fvOd24+efikZnCFDPOzGWG9sFsH7qhcWTQnHB/wZ
caZ1qJl1vY8SWFNCHYLrSYMt15gv89sfEX6sR1nZ9gbKuZZvb8XTeo0mmVOqZRoW
VvJIbUt2ftl/TZtFAUDWB/HeKqUblyqOqfDc5FAPGIblaZJJ2JTqQUwUAhkPf4DY
rPBOuH2vbe38SCk3ExFLjDsX36d/gnDC5AfPO3RdkkXAfK2uBZOGJ5tM5b9+YjzR
VgNFmotfgFEfRUxpTE4sAJ8EEModFH0mXeIl5qfW+xRRX+ifN/qVvcuGrgJS5uyG
/tKFmJMjfcWqCu/tGcdBuDpR1FfY8S6AmLiWTVPWC+m491nFU41h7k6FRpxl7KJB
s8UAUImgLRXfsm0f0SYbRT9jZajGPaJvlXgbkRsmfCMTzUEOzXXo4N4qoSIyVZk1
pbceBLCSltnHFMwYuimWd/R0LMxssqmSqP8wtTRzYcRxjReGSOuJiq7ghPCy8Hf/
JiMrksQ4FEtqjfsTdT8R2bkXTZ8vkSMd10K23OIyC5ba595qI+omzC99K6veTtEW
b9e4NvbaltnyF4TN3UN6RT5CZnHWTDkKcGcUVtzF8eL5/9sSDHeLFRaz3wdgKqPZ
RG0lIx4kv866IJ+T4z/tZ/8i8ZPhozOd+njYyB04jvTkU0QIjmDC8kAZfBHAxwMx
QWeopItzxo0uBCdEB/FEteis6tq2whYt82czSpi+wt0e2v9AuWwndk/6lBVlklfc
Ebw14Ob6ixDbskUan5ZFL04JMKfdyZdLK8iGBZ+tinE4NAFeNITKdRiPbIra8PxE
xv5ufZ3Yu3agYxjj/vrgJUfiSupoFtbXcj0sAg1O9JCgZfx3HL/SVV8W2xWoL8mP
TJRzz2AokDfb4GPE21McbTF8uvBL12bDnJrsPrextED5EQ5pHDDosrEvpoFWoVpM
D9xLqzgo9PnS0fmi0i+epIQFk5qIFqkyjD3NVW3aG4YzJAVWCD4BhB92hAX6Xe1m
N6CZUbCA/6Aq/3KuXXmZZNioq0mr+cSVEPURPM+V8B8XoebMrp6PdxHQjBVoYkyd
fOKnG0BwE5pv9+s9UlhnbR7em5TtfCMOBzNyzY6WBvagFoHGRGFvEo5COcEe76fh
FJyGs21gFhh/j7Am+lh6if0Ahv/MgFEB78/FZBCZRZbsAEAa16BWtllg2Kq3tcjB
sAe5pl6N4EdPK22WCNUPxg2ie9pnOSAWBxYdG1Vu+EiYjl3sMr39n6luPSD+J1yM
dAxjs1zT18z1AW0ACqApgB+d+TjJeYM7TukKA1FMc07ZuFuoKnD43jVbc1IA+HoJ
XkjnDxuzViXQXbgTDD3IrBuFXf9VHsiHinpgemmbpfrxYvJAId0XjD1QXgAyqrkh
EO79TeYGaFnyWM/jZGVtun7lb3hMcOEMVmUiSak04g7NtoycrFVLidFPKmcmAG79
ha6IlnZSdumZi7MBtIXiN1sZGPrQ6/PFLE3rUXoALiZRxluTNRlgS9SN8w47yZEl
P8oyvECnOqdRKXB4PXp7XC9kexgCh4I1D/F3yu84W6c1mlt2lsnjED2mV2bOgRbJ
3zC/djCtvkiDpc0UQHmnMZYJBpwAqx961vNgTtxl+f7wt6/JWNiepvE3uhj46DQR
cUZ7ANLsOQSp32ZwHXhYNFo+6ReB5lO958HJhAom+fcnpve+go0rY+Mw6A9WNRz9
dXfjc2EfM6QZmArkyDxQg1qLhTcIWAkBK7wW4FrC0O9VXkwaOV4erHezlEeO1PjC
tWOIWgBJ12vwYodSM5tLBZhePxscwVhLabtzTWPOgEjemDnn6o51/2Wy/4pG6zg3
7ApDcIwl1qD2aV6myTfENuy3fpNYjf9wB5Gz9ijGnw8XKJKMKI5/0uXklj+xYwVL
ewD/lwm3mdsURmKeGPjrwJWrskMl075mjGIe8xqmvskVrykseJSukwcBoHUVZJRC
6WCpoZBnvTt2csSs4DbpO0GtaMYUoH7KUO3Bcs1ZffrUVppPXv0J6k6QU7n3MXqM
s0+chngMwUxM4oBPaKdda0l5+R7GnSXatsE6LaK6wyQzwRGVYWuyx1gvPuzHGYat
73rZkFmnTXffQqomz2jM24QWbEfWtnrjB8L/IAj/YbDaxD0sD4mpReWw+4Fj/Jgk
ahNsbIJmKYgjRnOMaL41429gqRkCowhWhdg44aS+e+ttf+zR+O3D+WpxC/ol4Dg9
gb6NfiW8KZ+cfq5oI8tZ8FQmjPfInc6LKl9vg0D8CfdsFS/ESjl8T9XroZ1THanW
J3XZdklFnlMqL4dLiWKcr+kRTtndShrbFBHncA4GwAUqKNVaPGEXPoyxUSKI81+j
a1yu00DDbSybxp0UvPwz7H4klfyHJgHPw/RxSNMc2vznC7dLQeAhiQNEMpQWfM6K
+V/p/5buA4Is0Hs3+gPg00rQsgrnICiujg3RH26NPhM9iopo4mVVKHLufXiyBPQr
Pm92wxTbtR727Qhh5yyDwewsVd5SNSAAAptwjt/2d+0I9kvu0yQO4Y2TGBSn14Rj
Qr2mXg8d+xqaRApnH31oJvYrv3C588bItYFky6P+D2+eUYH8VwW9JvlEhHFuieXv
VUVQ13y+DwmOiR+U2tXmOWJfhRWfC9q14B7vFY5iZOmtZC9Xh9DsrnUdVF5Hy8S3
XDZDLz+n7yIkRqNTSBNNYQXxgaVk8FRH3zeOUuqgAvej9wSNigwQZQGWjBy/u6NX
D8aHN18cTw8k0gU55qvz+R0VSTpkhWYta5NRiTcBc0oKjjVOAFu4y2HEv7iARE6U
RuLsxj2kXGhRAwM8O1aDNUNAny49LMrUU5EukafWrCGc0IR3rFjlvx5b9VSSsLg0
6umEMGGkgmiKp+uiafmTb2Rm+N/9NLvW+bOp3PD4wafhcRLp5huHu2TH9BDzOKq2
8zK3tvvbr5sRD/P04PxIFTcq1OBc83qVOhfIUajDsGnKSLtCJglZVGhD0bftLacr
YnDM5C9ppPat+Ozp66GoJiPUju84jC/UPHuIZUcVVpIgKY5QcULhg1nEYr9suWal
TSvx98ymZsfsALSfPjg5t6q9s6wVMls98MnTgfaPE7zt4Fj5dMJcbDVkdFTwy+sJ
ywlLCZKRMXel3dZz8XgqANfDqS1U263fN2FaWCs0H92kFLEh7PCIa1ZruvGFtpIL
+t4c7GptIEGq9ql4LEQMrKeSnFmA4r4Lms+yskTzSItdKh0II7wYLWW8l9uipe44
pWs5iuj7+7rvWar42fSKxmr9aDuTtmZXZbC4slrB9XkIkNHRByqR2a8cB/t8Sblm
FddrosTnJpSjhGIcuZ0yoXkLyuMk4QREO3qJ5/SvNxK+Y4c4Np5ZFSlJRT28NIMV
iIfPNEhIOWPi0QiJIMOV0zMBte0XpVSBNZQw35GUilNTC5I69YJHLRi0vFn67sfZ
BxFgqGSZM2RkVX7nK/E2tbYBinSbm1j22NjGXWTJCaV96JFvWsDj3iM4HZqCEJzl
UgtJpwOW/LI5Rbjob69JNsykp+zVx7H5YC7Gl+t8+ZUCmovqBa/B0mkzGcqG27R/
k8/ZYF2Fe8NZPfam3qbEerqLlsj0AvK2MtgxJxjZ3oLqAOWE5iWEfNQlRp08qNii
x6y/JjcifXB99OgCpEFDWMKxZH1OeShhqhc+wyUaX0gsWT47lE+jCg0wnW6zt2n9
g1QTn8IWfcmooUTpIvbI3ZTbE/QG0jGswfa4bSnOp73Oi3wJQc8U8cU2d3DVOJru
/YCbg9z6XLhsQmpMhRGgBoPwKR66cH4zt530SWRrWRHeV+p/t7DVeOWpIKi23bjk
3IN8oYbFNIm3n4MwODTvYtqnxYaum1yvmrkTJrUlbA1M+YFJIfx5xQhlxSQvtzyT
QpJMbF00RjrH45jD959dlxsUsOVhXstCdKHvOmibJQOQsqzHq0Q9vf05leVq3qtD
g9axTudLtvaAkorYrXsmFikghGz7MWVdmcsg/sW2pmcUrv3LN4MKeMMFW2g6xJbn
jfYkgqOrlidvpW/U3RKk+pV/9+vw3r0FfAeH+Iuk3BWfBRZWKyV7eaXNNIQFRuVa
IjdoaVjdG5t/VLHWlZ3D8bP1BITxLtfR1CrJhXA9Oe1+9cAMnlSzMi02mMOa34Z2
2CGd+3hOILBddC+X9pcW/mTfbHZrclkNqlLwzyeW/84NSS/BbQSHfM5T5peVAiF3
K+vAx/Xopolt4eJ1HfJi/XP3fmpfiK61OjqqOWUmsTiygZqET4fzZx7ICG4ST8cZ
i4twDeUFiqKcjXxol99/gJD/1V2C042bQPOof3LnutDhWvZ6cMAnFblIrKigPYud
0hHS3cB4T1RkGLC+jIt+gjFxSS4hA9fPmDjHE63KIQ91gFqfU5AesdkSEaY4OInc
Ivoms062AoIjUv6QmQvg6+dxug7E3B9v9LQP+J13KYWoseX5rg3eB8C2ap2wsLMe
sUyjHQ4ie+cN4gsAB/E+zFmYxhXo8pquLtloFVij9d299zbKnIqVzoeyKu5Y2/4y
srFbhtVPiuskKfyNER9LHTA1g+bQNnpCI9B/72GnthSwvtG41P8dtgUGcgAlu9kn
KRXLWrcQ3x5TNF/GS1MqbRNKbystPIDvcLOzfU5GzX14RU074BcEmhQka7sAZ73B
4kd/l21PHbd2fNFy2IkYpCyPUYe1xkQIlfBMSGU5hA3oFJ3IIN+chsaL3cE3Aj29
FMvekOXhgbH/b5IVMjPgpLeIoRaeGHsxVt2YwJIs4JJCfLOdBjpPBU+6e1TMGANa
CkogtdAZb6jzFVromk1yPYU33yc96QhkzAKTkfT6+odguS9dofQiFu/JuW+MTvo7
7hFhHq0ynKL4uGJArU/tBHHwtphCaeoi4eqotjvJJ9FdorfVTp8wDMMmfAr8lSLK
edIZQxzlm22Z4YNCG/1A3izO7jw1XLAB+3sXPNnzeapp+dEca0INDFrTFRx+9vTP
aLlMstdwJVQuiBwHO/nUBKbySkCP3gy6LP+6QyeEjyLWavrj+LA56SFSCNTlCdK5
s7rosibZilM50PVlf6rvqdbQrkHw9pSFsmLoDj7P78a2LMGPEF+gNSDTgt/uaVdu
6+pTx10NXcc0TLln5/cM+bT7uPajg6FrZNrHAY54h3/rfaLNuUcHZ5AT/1AMS9Y5
nKiUvlzf1avdsIcqYkvsRVQE30UXG2ne549zthExJvUArlVB9RtIoMgcRegudG4c
//txtdAkFZvg5fsp4NBoXBWxa1RruyH1xFxOEefjpYrJlprM7Cr1Hv04pLFTa3L9
4TqULbYiinGNeGAUVVUpLLd4/adiB7QkzPQi0mKCU5f9HL9RT9fWZgn3b6foIBE+
Ub+iOVzc9aShr5B6Q0FqD5DY0Xr0hJJj8IW9fVOu4U82mtLj7PLlt1wa/hEPNu7b
8mDAAwTcgMx253eZtYAQkWN9x91xu85yY4dHRwGHRiBf876z27d8o/PELIpahBNp
FOjBx+dSBYc8XrD/NpjXcja7HVPeqI13dmGONXQv5sArlDkDXr39JEpSC3sPcS0C
S2dlwPZ+ZoRqJLVvsZ/KKFS73v+4VvsLbEd4MJ3D+0MOx8O+WBN6Q1kuX9AOOwmW
6DIw7Hh/ANjeCcTvU+IVR2ftOU3RNAy/l2UfzWUtqHCoM6Iz6d2jm4ELDkUcavcL
5mKvHVshAC0IrbDyQso9SP05K/00odNwftUYl/AhFgqwHOM46AdRYrPdqOVNCJ3k
REs8WP4MziMj2Cs6lIKf6wBFUz73RhxsLQ/3DJW53iT0/YeJgL3ncKReqf6Woi6m
lXXp07VVCxCkH/cIfARXr1vu1UryZ7FVhhrppM1tcS+yUoX9pqGcONX0BDfBB5Oo
oEEcZOOUZ/F5Vx/hI/lji9rq0BoWpZa5nObZ8+2zSv6ri9xz1+6bbdsyEScQoIar
b79CTKRSPfPLq3aazPdpN+bT8sf1MeKfY1RTgVL72tgHPSfR8gZNnIeKCEYFUCDr
moMca4oII7tonpsdwTfB6kA37tLlSFDaYDIzUD3YOaLBMuiOIGnRz2/aFQgUaUTQ
L8EY9QcFZs3Lf7Bnnh3qoYpXIg1dgPG7a/aKaEp9zJeGm4Qcdwb62EQyr2Ug0CSA
8HjkWIVH9o5Z1ndcNs06ag/ZG5Hn3g7yIp+EGEgC8T/lTiHooQYOmMa9N6RM+D4y
8KhR3A4Nqw4uPVtW1MZ0jKiz1TadtkLfyFRDg30U3jueQX4JEUcXqdAoUESyWIGg
IrHdMtMPWKfv9YfmWpmCEDGpwUC1Ndyn2Xo0Pl9nJcm8wDdm0vKHha/L6TT3YCXI
noAMXUMaXPyc2wYDmuf618uq5Cdm7bK4rSoMT4LtjY4/9EMjTdRk8kqrvjg+2iAZ
z3dDIzUy26e/Vw3jhDzzovhHot9gqEpJpuZnwOMsSir8Zrsij39tl9qgmTBTxgdF
rTFchCnTvlV67fHs1haPilU+dHw4ljaB+etE/NuKPF6P1g4t90ntpTLpzZUSSrq6
clIDlBtUKNMUYm/yOtcYKJE4arCEJri0IMVM0JTFOf3faCPE8qSiF/yn5tftQV1s
uO+8wPtVJ1JWNb+wLg3AqS+w3Ixk9yf4AQZrypzQlTCLRRxRwhuSpNYw7N++Ye7b
tvAYE2LfTUrPRuwajpOpL/+DMO80n0iwMxt6wP8QKFZDL59nIbDzGKncP76PTp0v
z4P1kMviZw6X8Yn3QVUBTKQkbZryAtfyyhnVllPzmOaNLN4wP73F0CvvJLk0GMSE
Hc4mgEugbCPMgGS4ibmmJOWJWjlCYAR/9lAT+ZRf1TJlUSPfXohLlat79BHjk0aK
5hKhmyfkd+6q/T6bZRr0FCEVBUL8QPI8ELLh5zT2dnp+4UTEe3aqzY5Rl8ZWHDzU
2soFko/h9SQ4cJfaIxBqylwmDV9Qt+Zs9mWmyoKKQ0hdpxcTXjm0yaTdrLi/fyJU
0M1R9nK1WsL9o2yw/TU58ToxAbRhCFu2qm0DzcXeQ/fE3vWkzn2Syz2LmGVsppP3
uAlalXtO767vqJucpBoSnuziGrzVCoW9bPDiQL6W4MgkesbUlClU6/NG+Nm3IM8I
N0jQt3NOZyz2qUAr6+miXTi5+HM6+qYkkEx4tTZoRl1nwyJC4O8u4EVA/5TyxxtJ
JhIgaCjUMNQlNSMOnBVHjSwPVNDQK5ouM1NpspnHSONfcPn0LrYSGKEtHj6hgKzL
ccbPr7JIotMa3chDGi+5HdHHzIuDvgh8OFvL7ekeB9B0qe7XErKqEGTCzFIcst27
u94InYH6349biltTyArV/j2OdurFEpXJUHBaiRjZIUHo4koYvInyEp10c824/oVf
HWha/NVX7FzdejKHdFSALyHPSXPoCFjLDXG4wV6o0AanRyR/f3jn5wRd6INzrCVo
amFPQThVkIiFRcz+bSiiazlkexqUFpzD6b79kPUyjqo2rvOtHPqL7gF2pmEVijQQ
7aGmQH+nnxsRawYpaRZ/h9gsMQWZI5qwca9wT1fGBUaY+aTT/aSNDeO0Pz4vhmYa
s0WjtiEwoccPurWPlMBcL0zSgMKWrGiZDEpTIejuj4SZdVocx4LUmrxPHE24EKzY
JXjgPvMlJmGLUGHu3VTndjAONe0H5xT2Y4mu8Y6GfAa+SEHGsRo77VsHjyDPo0yz
YAAtdiLrafWwRzP1BGeOM1TPrDPhoW6o4wy3B9vyBjUIGvQEttSsrxZe4FD1PijE
HoasOfCwkof+dzyszbPiA+t5UW1ALM9eaBxAIR2GJNaHgpinFHZlkBV+hDh1QDsv
DqVx7Bze5VoczI5krrlXA2/nxgaj2RHNaBI85rql3wLBFNebyqnCiiWeDcrv7i2P
RjGjJKsMl4itN3jJBTscmjpdHIziQDKh3+nv8RJ77jxw16d52tZHnvsfQ/TUCWIs
Lp3G2xJ/Cpw4cW637yUToesttBF9JNtXuAQfwXOmcp+js1oUc+vxZ48VcYJQonem
8Bl3zXqtJQGIuNFD6y+6bzmV/uYWsLdjGsdWKaZEVYfSmPCE+JNN2pQ007GRYgqP
f1DcO0TKNTfcUW5YBPkFKvyQbsIQPzNd5DYhYgcy/lAehWBUTUDEPKR36P7Da3iO
xwZFB7J5YLwkcMNdBFZ6frFQVLISvI0IhUQrglkRRC9IPOnYn2cyoY8eWSQ3y47S
7G8ugy75AukiYYKQxcXrNXtQvjfDe/cPZA3bLif/X3ScBv3IFHP7LB/+90SGmKHd
Ixpg9YMyA4C4js70p8IPLiT75Xl8RsH2tzvGEzOGhHnMBU9EP0WXATpW6zJ3X52y
AmA/HUEVLtTt3Y1/YSkFuQf3y0xeEjnYTWlyhxUEL5JqugMYRZiGAjDmjffhtmJz
nfHE9VP5Irajcm2WtMKI6lTu3VsUaejbdCiptSoIyAYoyTrh7gSFX+jCJlc4P8Ta
b/uz64iSEANLG3WYdKFoFfW2u4rF5Zm+gemQasWaM83QGMghIFzhtzLYd0V30Ygt
/+8K+YOXK9aaZn99NXad6/UdBvt8IbIyIfucAz8zxg4/YXD/xhHKL67HpzYFMuda
28/EJxFsCLr+FNqxscOedOfwTqNq55FfBMtMT6VlVsR66EMMYwOTcu9B46Tyai+o
TK3/ErFLuqnky7a/tL70eOxVNcwunE57QUWNg5OpzVlxis8Ssx4jDN+Bfo+vLRY6
lx1bZs/FukSb2F1z8YyOBmdCPRb2iSPeEYjoH2UXB9XW1ULihp8lEqatPD90tKGb
KoBatl7K/pCHWkdH0ajW0hC3hRIHiQ4g/wbYAF5lv9SqKMNGXdhdlM/gOLSird/E
u93FXJPTGOwDnHNM+u3rRSnnnLng6HgIU5Wsq1Hx/cab0qO0KKYI4K/woqKuzYku
hLTsFiz+NBWxmvfSFSC2VDVZydxBD4blwiVvZvHw7xvVjoF8T0CA7inVlSLOq89t
AsXSEjp1vHPmS1W5q9d1En3BycPtn1/UsPDEMiGhXGydV3cKVtnfC2+nRy6uLlMn
oevF+qKS2hYxyalINSxu//4eJUX5jy8u5aKBHw7IZh6nlU5Wq1gmBDAK70P9izmW
cDlJgD3FWpmN6jIEtqLq1Afb6ALL1v5yM2h0g7OCJbkbc2D1VUyy24MWEc1xLXaZ
dO4NymelKQ34BhOcU7685fjc+jcjotyzeWxoWwOI7ujsH6/k9+JIc6LfRLMXUc6t
ZKNwGANwRVQlrFE8zHM6+welpOuDR4yLunlnHgg8QtYPC5EB7QRnKFIEE57+GPck
MMlBXgxlRwNVjOIrmAeXawTtC76VMoXNnHY9NkQXGgocvhRtSnvT68ECBHLTAEMt
ePJtoBZtfseKHkvYD8TzhGSvL36xOcKx0HXpM93YOH80ZbwfESMIxGD7as0gjQaZ
3xDZcqB+Y4+HW7S/BlqdVEjsix73i2k6Vwq/eZ+j8bVZaJpFRaRfCFlSCFkP3+AM
6Zzp/Ub/8qBtkqQNbqtAmei2tlSakaHq6abyNg8kk5YM9qCf6kh5WTNMgWUsJelK
NMcUZ7udrL3Dkmpc1FFwufLDLqT8GYuLdNe8vIyB7ed6hBt96BzHQ8nQIckiQDZf
x/yYyhHnaPv7hJ3esdLSHgIKKN/x0mxQF7b9/y+g2qJZwG9zMqNUOlyjHQdiuBsr
B4qysklS/eu6ftvIW6JDulZS8eijqZ4tv53+E/viqNTlY2KVxaQp8JMwkC9wyrs9
05Wcr17loB/bWqWjTERNhDGuP56rXaMl10fYD15F2OnS9pLQnLeiSzIA4JoXdvr1
KRN852uOZ5AJSivKG1f621w0bjeKZsfw52SX/FpMbiz0VRO8qOxEhfajXk5QmIpL
sWnRDIEPk/bF/B47yJCYud+eLpMPCFEbp/LAozKRk2rcQkLOTuLpUSkSNEEIlxih
RI4CsT1S2XgGbSN4Vgtgf0VCYf7cK3Q2omYpEJjqxpIK6dgGsDNk5wq+ZyDgc2z+
22YC3Ih7mTVvCsSTMu8AzO2fW6a1S/tcGV2Kjvz5BjzImSA9/JFCgc2hbX8mam1Q
Biu9UzhJvOhRk1Of0vb2PoAOw+4r7hiVIF+Xzy7pr2TkcihWkgP7EaQLWBCYDFQK
dmRxw4lWb/62gf/wOKutts3iMKHIiIf6ww6mERrNtbg8SHangvj4mceKNe7Q2fQg
v3V8ff14NukItfxTw009JBEUpOwJ7OsS11BqSfOe/6hRz/t+omv9oNxxiyoTrgdu
f8eI3YfBiemqwjxVRQQTTWtXaQgfiBY4s4JogS/v50EQ5uq8qo01zYT5GFMvgCjm
2p3WjplXD6CUTh8DFHjeLvFd2mzzt+BIAK4DQt3aH9bTZSzlRsJNYKOioOHaVFAP
L+0mwsSEBXLi42Q85YcDpQ3MymsUUEtfqkf8IDKoVo2xBBIihDGVa6NpRUf3VBP2
YNsIcnx/oP5ViSFG7HTWf/TqT75qTiTW71InWnGDc5c7P7Y6hfKSOsSt0/U+tFQI
6orp6KvI5jJGY2yv6lCdIWBsfXl8ofbh483c2NzhSp3y+cikYtDXhW7OOlO2d1Nt
DXhPPFeXefT8//xqBFmVrKr5NOZj1n6NSVD4u+WWG7/HUjwW15OASZFlCAaOWEiB
PnDh0CEppP//D+jl9Bcut7AK2K4WaH69HpMDMWarPuKD4YsT3SwUV0YoywyggbUQ
HZvoCMjuRqTS+i0oxxkdFBh1SkCWxgvtsJUVBainn15OCB6YBxeD5vO/deM5jQRI
CzUJcSFg2jGWPkImniyFx6MjjgbKv3ldGZQGzA+d4tt7OwhdmtFC9x3V556gEqEV
oUub1xmGmi/e37QLBgSxcdV86/2RM593uxqvr54GJLUTSzKowJA8/6FZfO7jPk36
GqvyjXy1bQkq7JCWmNLu7plDzf4lchNwAMjylmtA9Es5vAOp6mnKqAPNzFHYKCLv
6RUoU6jgnTvNNdTtPOrOKICoP9ZhDYxLZRDA2izok7JTaW8WWX0Y4FX7pI3m9Vsy
Pd7ABVnkOtTytJ2D7Z4Xute7qSaNOr20xwUYY0wSzngT9F5odOmz7787NGS2CUYi
yKGxzXB31eoKIvvkp5EuEQ4Bs8cDtU+26waETkgdGxBpwnc9NtUvxLV7fl/I2O5G
Cr5zH4cKdb7NDA+b4wNxOu75hcmqWNg5Jgn/XklslprUpzcdgf+aMeipcMX6/wjn
JbqQO+mKpe5TRoCiRCEVmG1kgd3Ex8zXvJ3uptjh5lND1Oz1cQBbeyDwaygiOkNd
vZmL4EGSdE+/B5uU/DNgGMBIy9BLn3Sg7BrNs5taohbqYwWz8iPMPITCpwupAOZb
MdRFzO3KltmrtIvYe4YDsM7v1GFJzSCOOT1PhUUJhfKv5EiFfmnBQ+O3HQu5eloK
auXBkRYnbXam3hrf/eRJT91amTgS+jS0Skm+pO2564kuAGFDZzBO2CSqBOZZzh4X
qo2iMb3yrktDF/QyigLHdXuTPJU9Vvx1eRyt9BcPVcdDbWa9aX6BgcLte9vb5UXk
nqQ8JtnPcKdt2WarESWPIp+qaxqbRJDwfkyJX9RApGfzlIoGWZmMe4z86vahMEIZ
CoN4+HJDEJYqjjXiZsdPngI3aslp3QBBg5gIScbhanLyvgjmd0lbrUZEIl4v5S03
VfWmN27GiycthH19Hvgf3++CEVj62zq9mUmUr9isfvehBjUCS8s6BVOx1+nuUqbE
4dCitK9Wc2Hoh+lpvdGwrEORik52F02V7+gAkZgDxzxVpQR7mILo3cPBF3XSlHPo
dclQWW7YHseEmKU2onB1++XIvGHuX9dU7O0J3gSBaVYiyB+A87iu4m9mDgQhz836
vdwcBhH34BLTqmC79GEBgQkethFN8D/84Uo9HwGKneRSgwdMBIY174AhgUJFR9uj
5nsJl0vgRI6JXck9LhGh+dbqN/SWvkE4o4g1iNFkE5XofUG7lZfgAxupmkP+7mSj
/KhicHjqWrtBWx3dAwK98zlZj6QEhOsRWD6OdDP+DsMt64XnUxUzjMzknQ6T7Uv8
ZJuhGaNitrlf650AjN8Bm8w/u6BA+acsPcM24snrJVcZooQeg4FvlnZtyL8R87BL
ZY72iutYgkRgGJLfPpMsZ98Xvk7n/cT65NoEYdSaC0F4VZRgAiy8Dd65GQMLnEb+
tEbduOmmNOQi1aZhf2/NLULRfR36RCHrL2kkP05CSkeo+GBAuH0WQzZwZRqyF+iE
hfLHriobLWmObRMG1qKp6vAckDUr4sVDyeg28WI5unaf7Dtq00aKDj78h14NFLd5
aV7iKxsOzPfrTYhAs8PamYdUlVBIU1FzpwN7dTZIAef9dCXP5ABUl0ujy0CmqEqi
UXfmFhCFTrhevMvqkPmPNb0xRIcYmU9d1tzcRj9hbYYnQFG1dBqdopj/Z6wPJAKN
s1322+5oDaI5+10FzzpNMmj3RvDZOBnKf7TBBfZZR+tt547rYe/7Suqcd/MifUlr
o0sD/LUbBGt/D2SOLQkXsrtSP8kkkiUaRGcOWp4f03XSsvvCU/M9Ej17oCVTnHXF
NPNa9MgnLAUluxuR/4o8fQOWwXvWXsjDxLHUmPII+1KvPrkdWFB/gx6zERShDHWp
7stxtXnxq/rMMgm8+QhQ737QmFqW0CnNVXWlfz6ohqikfgenB9hrbkffAL/zxyhq
PdPRizLKlmrFtvw8ZICND7SFw/HFpWEwrEfgld5LzZhp31+ZVRqKJYB7isH9HqZG
eac0U3Hx0z/4JHEjqRxI3pGhG4WCa80+MAedu/w9hVeDVYKOybSmCsR7aY84IsKs
KAUY0di000qYoemwqoMCzgKc3w7DiW/Tx746nMaoU9fAgjEXqOj1ZNZ094OPP6+g
xZKF5PV7pJ8m+uksGf2vIWzZOaq0ZcswEB82xWlaW1EWq4E30cJbl/29/4qNgNlM
NkfcBRwa3+f9t3f8mltOSOnZogigp2VEbRWClY30Wi4waIuzCjb7d/oUDaoTVZqf
IV/4Cobeo3O6kxDOLx/M/ABJBBw+wvqgCiHdopfcPTChWi9Az0Kp/zDpdrkpL3gV
Lpsm5ZlcuDsnzBBg1k558/BrvQrJ1V7zYHf/VCCtgapLrQlAaMZo9al5OtiRPPe9
EkTzjaO0lBxYpxpjsDuUV3FNIp8tfODisaoQ3ZbLCT57DJcoW2fHPz9udqjb8syf
25+S6nGm9MIokboEy/IChY+iu4oD+4rrHU1mNCQbZgTKL70WNe8KHOVxB5Qlcg5B
nj9UMaGCoxdN9wS+96270RpbyzPrNSUUII/mFni8MNSNKUHp2RLehlUWb6FOMtk0
bNqDP2vTjgCcDaRLcpdy+Zi2xhOt4oQL/7cL8jMpMj8XYpBXqikMNmuRsgucZa18
IRsnXlLUvDWigyZY/FiQ/XxeGpSeo6U2Rhi/1h3my6F+t0nXpqmdIemY85HcIx2i
+rm7X6V8EOZbm29mUluQC8ZftKwWmul0qGEk1ZTYIq5t3qNJ3qMhHlPGT0qTwZc6
iZewtVN40eIk1Ql9NjcAMIl2OUvBPwORTjKBZwQq4vcuMv2SffFYnDev5gPUizYr
Vvqw9MO/SYus5kpJPsesFF5bkW2sBh2aLv6RD6R9rQRDq3bruKp+tALewwffItMu
ACy8kHmRKwZm2MDMsLKTTag064ctIHLMxjtSaOc0gpfkczhzdU9ShKNV/9jJQ+v+
12ojC8aNyadK4S3WK/NghMViDtt9xSht7gwKGPuwhJR5kkVx0DfU545O7MmsJjMa
EYsJZd0VuytU3lPS0dECmc0dnAGnmSWLKyVzIwTVJ4UufnTQHirNDgYmmRtWQWTn
suIW7xngvbUfIjrGvs73W1pEspG3oPOBAZy3flFpZUT6l94MtyoEDcz7Wk8LQQrh
EIHUy6HhUB/agevSm4/i7JFLfx1pgFDewPvcu7jPCw21ro2E+MypxmufZA48bfXT
IxzkvlBdFtbFybcfZeKoUJluLoeXHAJSYDKF18HpoXoj0uz6E9+lVryyinMmUX+U
tD4PJ2W8xGKZ45Q7hV+3jwu/61ArPrd9X2UXVqZTxhzBqqEGHK3e6qb40mtcku7O
YR2gozO3h0Th8CujUEVCD/0ukCfFA011GhorkA9zavaOnLQlHBSJj4tB71fNp4SG
ta1Bb7fQ3Jj2dRmXaerYiKF9klfnDymLeJca5KkZpYtzhDjyDBoeFAPRq1mpREVL
JmgyGZQLbn/iwHdr5QWWhTOyqI7G/kDs6pZgjIUhVDMHQOqejzk0LYUFFrTEKyqb
JQubX3fBcfH+P+kJbb9CfkP37HHg3Gjc4i2cnpJcuI2NAw0JhZmMCSzYvU4K4c6L
FCF93v4ve4cz1fxvYPEg+pQDBZ7Uc3iLRAG2+xGYi1VRR1NsTqFxJzxNhkJvb89l
xMgoOqJbu9hibr3pibj4a3vZXrilptFa+lYgarc4Eo98HtrpxMfgvUAdSJhAwKuw
pdndqUJXH4Ak2tjiZwfNd+PH958x5fJX0XhE+qAyU5K7rilC1G6Ih/C77k9Fd5dv
3jwUFXy9nag2bG8sQwJht/q5yHhy+H4OkIs6zar9Zz9UtscKJBrI+M5U/mbL7t9R
UR7Oc66tzG1+p2H9C2q71wvfgECYoHibiN5oQauyGYbwdlRtXGGxpVlyyE7Jd3mD
ZVTtctte3ieXhJsls6T9WQOm5s+fo2dbp3BhtE9VEJFGJUNB1rnG9mYW92/AD2ep
Tp2d50O1LHvgd9Y6bl3tPuvGdwLnV6TDLB2lN2UmFCHTxNEpH7BlMM85+IMkMTmh
LIeKcmMtSM7zqCDT68halLkTTSzoSaa2to1B8Giwx0kF0eSpGIeAlOqMaH/ia5Aw
OWY2aWGZZzbDUCoeLPJdQwKhEMIF6amPgADrWViB8z87opkIBvax6nEUvp0+XJXF
UPfqxf0PfB2/NxUnTClH2GdVIjVIZzyuVg5CzFtVb2EL7ynapqXOYpPKD/qP2uYo
w+lTowvUp5rJZZw1BC6t7GOXz20lg091bEgTgofnQG42pGdjmJoRPk9j18GoIJ8Y
0zqwLlv6jFU0vXOV2hvG57lYVFHARA/54DT3+JCsgvwCQRgVJ6bPv/7YIvJiKLIV
FGRYuS6qhD2qTCF1p9fEQbDIkVAzPkCXDWImm9syI88bKYyIzjDTGbOWLKFX6m6I
1Je7CEmkThG+3deh7+AE56q04D1YrQzWPPsesN+7xtgIBVfJxkqqCi+hkszM5Ebh
RJWDaEQIp1Gt5GzrLDHo3LhkGKzhAath51hDswz1Pv63h2FYLv20DEOTjuPfWEuT
lK9I5MSQNs+I9gX1zyARDBK8PGfLXr0ZpOi82cLtp88Knq8iCpqhsZyQPlGLpTDz
clQixefx4l1cJx4Y5A6MuiPu9erjt9ussmvThXkSGgorZCSZ2xtnGmgValE0tq1K
5fBekZi1A1mbGz7mU7lndBMEUvxSOBniGhuoUZXP/MOocvFgSuQctEYqpWi0Ox0B
Yfi+mhnNNgFe6bOYg5SPIs+ThshK/VyAr19UVR8gVYj3wnChh9BLcZGHfMIyTJQF
rDQlv7isY5unMa7FPnvmoorfEDCZoJsZJAcZqvKTNxyIqc5KTXEaRma64EiJouA8
mL3XpQn/lANcpfwsUPcZSkEACCOtwNxrd+vv2hSDoqtme/NRSyzpFlY6abZCYqLg
jGm/fDH6Gv8tUTRr7uNI3DCiVa7NkA+yFZJS7w1a03bLWssKb+0YOKxb5K/vuECI
T0BffpOpphrhXoKrfDmWcFRntWbMONwmtTOSasugAWiEj71tyVy2oWxbZESijXJ3
6CzMiu7Sk7pK7+73zHvAtMFzueoB3O8ZOFclPPvAcTRr/e5vMvKeLkvHjaiuaXxW
Bq2q353Wdwudb16kSMzMFJMQmi62qMyzeAPV1HFI6omCHvR5bhn08RENjcSVaWT6
EhsEwc8I6YfGpT3Zts59Sse5l//imzPs3PEHc1XRW64epmgaDUN171XAiB2xD+0g
zepZgRTFwbTlij6rTNmgYRxn3Y46FPF9bzne9fD60jyGPZmRkiP2ci3GlO1Ol7Xg
OoULK1JuVcgSN3yiaeONzt+X820bfE9Ts3zGhzfW1c8oPKA2zgjqZKdbMS2TO4K3
M+SZoqnIJH2zdJSA5qwCfviD3OsxTtBOvqbujEd8cO9WlTkCJWHr7QA+GiDQ1sv2
4lfllpmmySCUl7/FBGbPaBsCUPkp7/h7Cr8EwLhcR0uPA3YJ9TZvTNQbVL5XYhiv
hctSbhP5z1rWf/Ob58s4Iyj6t7lkDAdkI+7HRDmMHq4XLXWYK/6wF/ixhRKY+HL8
XA1+eS+/m32LUZU7ZSyQVGwFpJb161aBxWNZXlq209VQ++XI1/EbJli1ZwhEx6jk
ndrVAJ0yoKVpExxBYrLBpGuaDmImh5hi5boIijQH7xVvu7cVQeuxULyeWH0nMW1t
J/+yV885uuJ0gtLUWd0Mxyyx0soq4XO+keiL5HqHO0BcRXG5LGGBJcUt1QWrutUj
9DlDxy7aFwWQdmUJCeA9ultEueWB2P0VlZ9rv+CcWf1EsVedpjsSL+svCVzWYrjN
AlRAtJmS+xJHdknm28anXpAaaMKuihTM5iYTFkwZ19FU122XOAIGFqT+R9Gs+JxE
h7Ec6xpZymLP7W8KzSeLjsDphRfLGKKD/9kHSa2Iqp5WtBIVXvhKjz7iK91L/pMY
CxIk4HnLaASvqOrlGJLzPZst+QEm8phdBNDCfSNR68G0wr7kKMThedsD5kbX0Lta
lI2TTFuTVX0X9oahqqj/uytMlRChp+w2+7LVBIdLuOuupJKM8DnEziulKhhcGi5G
6bTeAXXZ7b2rQ/8BvDj88basQlpIiLeSrwocOEiqkS6dTEu1rqLpatOeMuti4Rs+
KiEiVxJI04VnIcc3QLMYrXVt01U7NydLQTUDI8mrNXA/6udvg7/jCb4ula/lHuWV
qXRnZMVw4WWZ4mlJMoTrAWiR/g9E3lWxvxOGHZxjvqD3rqNZ5q7cC6Pg37W7bsrL
x8VOODoZ+vY/ia2vrfVIrPwG9xFUgJkBp7+gZFE7ReOgl01v829CrsyNE2qjjpdr
6VQ+Q+cATNbqf5WZN8mOUFeO1oQCYCI+nFOukP2JV3UKdF3hnczmU9fo81nkCNkP
oVAlFhva9Z3RAKiukMTk+qpkHfc/QtlFzj+SIkur9lMet8mR08NxK/o3Nu3lSv7+
NebM/WVlYKCOOmG7D6eCDJ/ZxWvTwn8dVnzPb82N+0KD3Hb1rb8l2Wnjbs/Lr2BS
oOGssUjaxMMsg1DvGMoeXAeFP8bxd1YsQLNuYa/nq1zgrSX0o4lwsm3RmwQSAQ4V
miE+hyIWTHTF3zFGisEoyyozaMbi68cTG5vvotTj1l5Wot00JfZnzT6a51G5nt7P
sM7U6Ir+DQySJPhWk7v0I7dw8ESA9flCvvni+P7xZbJsNX6LtibQ/l9RRRlNAmI/
2HA44XQAxSc5YKUPVpQDxMVT+VyBADVunWVQGLiPQaIDXALi5ZkihBgZGsapcb2m
iA7tcAoYzVSG1TUEHzul1f7qUWXGU343Lj/ufZVHp/hn/WhpjAsFEo/gTzG9YIve
RFD7H/k8BzAXtaW0++S8kxoqM4fNoeJ4Eu/uoRjnSufbM7CvFPxR3h+IZ8Vu1miZ
jvd+sDGrV70z6kIkhnqSbacBzRVYn66UB+t1mhaV/nasLkosdOQEio/82upLrdVj
1HQvqYn5ag2HnX+gXVzZgedLBCCq8Wk5YybUxQt9HcLuMbfVeCa/pBASg+lH3VGo
6VQTe0pvZo9glqICBboVYVoMnoIyozE3FDE4w9l/oIG/8Q8efofjoHfWHjXlHG+2
CovY58sMY/pzibb6G/eLnI6XTRypXs0s47q/Yg/T2rcO6BqkrwV19FmMphWOfy8x
gHHPBdycA7gLLwUn9/8EI75+eywvRR5yTsCS6xEWdFHI6jbierwFkvUMjJP98wep
7/py6O3SRjdhwqhFVTeKYW3+5Woi4nZNsAvyEH3tRXX4V19YcuyZDtFhP7Gr3LIA
1TRXLjoY45AwfJZboCbRFzCurLRo9x3x8gQdwq7JEFkZwW1683Fc5U0esHTWVA6K
ZMN+nmxT5DDzzZG8iMn31j61SYx2fNvE59VyBRsHBvYnkn/VpQ3TdJhAihvp5OG3
Bj9Khr/+z4M70qnCaK8j0He4ASGWum/aKdZtTBugAo35SLQNvlrbEjgstScFAojd
kXraP5MzrOTNsinoWoTJKji1DUB+gyWXDu9RmTt+gzl5uoTN85kDBUotrrQ2qXMK
p9WNdehqZS4gRzzO/gtdjHlMjQryhX9Vi90WtxrZ5cZzbWqlk9XZQ6mhlUCpgrxj
+C2GxklRRoiXtFgFAYekRto9fi3gJFVEXWVbBDNDZ6MizjtAifOnc/vZnuGxHked
7MmCPrMKoBIx/Cpw2xQQYAGuiDL3J0zfqGEdjNEBOHO7LcEqJVpiYbCRYgWhSyiM
tdqJah42s9ORlmo/Tcj+7uOhDNQFdx+y9cBBSh7SZb2HiXJwoVinx7UQZZ/nfb0c
OiChsnDWtvWhijf8/tP7G9VdeXBndK+gRXNlvEBOURvdZqUPZYJjoduGKOaeUZXd
Xqtxr6V5SieXV7rhrCNdxg+xcKeE7afXV3x5z2UZxmJaiyFE8sYyTr5QGAUG8ywi
WcN2JI5yfTHdc1Iv/TEkhXnj/kKUx/jn8vVH58z+Nq0oFlUo9GIR07oDpMTy/9Ub
iAr1+l4Y8gkk0B7Ch0+b0lUiPkzyQzf3vkXtqyf6D+TrTGkYuGywqD6VQbeRViYG
sWYhXn35lQ8wk0OnL7nKW9uVBrjjZ0txBx/FverkduaQjp2SaUXsNiLFh0i65Vmn
7wYe64X1szWIGUTDotaG6jU250w5GWNOOAcMfdOZ7s620WLXbhX4EUibkllCgRRU
OS1cyS+0UC/gCQY7nQ5WFOpifnVAUfBl2pPI1Bfiv3GocdOfrskZ7Bf3sSZnVbpN
kU6xXwrFyt/9t9PA5wq5ulrYAbGKkd0dMIeyQGBrV8rh3rpcc3wUqYviez0KbzDj
BHfsgWj87GDB7MjOXB7FGVTXiHD3dAFMW7kTAX4zZj1w+9MjByGHdkk0rZPnkfuM
aCVbUlw2da2C1OFuq7fdA7LUxav508hevz5B++7g0+Hnw8agraR9sXQSlPbxwjxQ
8iedxRdviffxPUuKC0DdkS5qeB0sfcwAHwZRZU1fozBbycgueb/o9OWKmKovMspl
RaEm9/NR4VaxHX3YAh6EgyUlFgO/HjD2EtT0CAuzSdMnBPM28zHBvD8u7QQ/39MT
wgAdY50cs1dqI+1dFJlDifFJ1s4syCBirdGW00VIyrpRs/dUbtwRO3IoCTX0xX/x
w3SgOS3+7TKBdfwJ4EOARhfZtrXSpvTsBywzDF8aa9l7uh2sgVpq+QOtSon5PCDr
D7SjTYjv9HPxIxievpTzKRGymobM5zG/V7M4bYfc0VXCrEjgtxK580UP/fd5+Tgu
LRrPH+2u1a++GM07VVV6K+UlnQRgdRBmI+Vz378zQYCGR4pribTd5zdgXzAquSu/
kZ0AOCH3/5+MWtGn/BS/+ju8JKi0J9jvqNRNu51iEP67IXGR3eSusx0YUPpR1B/r
okQnKqrnAoGaGrL14gV/piOTHF37GHOWEwLkT7lneU4o9b737ocmoSZzIOVeOvHH
0o9yhVH8flLxJOSewUkwvF3wPgUSrCgxoLimEjRgR/tFxSTUSJhSj8ttbUmILYbn
C9VdvFlPJP+c3TKMML1kdgBstRtNsJ5t5rM9M+FVc8yKph6uryjTFUsl+1UgeyJ9
HSegR3ZT/tVZBfGxHtAxzI+d48hRv5B6oAdxLoEkButT5j2fB48XeczVZmf72gT8
vHpNBBw/bCq5nkOpo9itM0VFq1LDAQBf/VVk7Ayvt57PHSBEAl8XcLyR2FzQ+CMn
Wn41vffXsTf6gCDqgtVefW4YOkAq8LBApyEWU9KavA+P7I/k49Jcy9gS+BaAW3r/
XGnnJSvxYE3/dIqZw61LoW2wJA15EJSqgQL9JLOf1kSpHdJjBNWIq/saSd0zUEyB
zTLe7Pz3e4lS4Yu41duXxgemPG5/IqwW7XCOFWmLKKyYZpSCR8qbvOlmMjsrFWC/
PxN6cyU06NTYJhaCWQefBgVdU1BoVMX3WZCaj4v7y0oR8i1uR/EYVmqw876KRy4r
AAvcQLJ03U1hN8+GACbR94Jnqr49vd0vQLuwQZg6L5qMbUodbS+EzW6aqL/qa7Jv
KGblpB3QGWzlKAoihdG9OCFLevPQLv7kwTT4ht1oNcotzBwdIynyv93Oy9IyDtlJ
d5cHXjDUh5uvYkZGMet/DsjgWHGEq8Nj794P/dAWzPdS9QfSIRAU5NKEwbItdPwh
vZE7ltpD4XsagrH1uxuQABv1NqmlkV0fABjw0Ov8NfVDjLChWgLmGCN6ITzfFhS9
JnuylEcl/WaadTtLdpYTdK+K4QIvwjQBQb0tgddKXovDenBxeHWPcrIPWw9RwWFl
S7tDHKj3/Q68EQuzKanGLBTP83kCxEV/HIAAXULHhsWb+C8ZufTzczomgRYDXcJ1
P7OldvBb/QtNy+fdpYftPzi59FLmlKDXxYskAOcoFgOAAVGel0JGxLwwuaKzAN2d
nxlv1CFCVZzmRQzxNLJdgqKEXnxiaAIUqlRKlH+OlrjHz5QrI5puhKRsOqyvQ17k
luX9BJ50pQQ3wxzFEL4G6uGSavQ5a/u0o+7wYA0CBz6viZftHE5ZE7YTPB8jWiD+
pvWMF2S6PYRT+lJBecxLW5GsppK0mtKTxy2jPySt+Tf6e4kUsR0FxEyD3rgJpR7K
hJ4F1XCts2vTOj6b4xZEfymVNYtLnabJdMW8A3oFa36q+3Hj/BHoCTO7Beb9NMw+
5bYWbkEYRQ2SM3gyqxChoTXwY5CFMJfAfKTBCOw3TFo4MOtSXs+sFNU/XZTUvxVT
26eOmjfTfWGwzwPNC9ybE/uwHYnqmCtAa3xHTfh4xipYAvTc0WJyghx6MJKXkeKJ
WNLzTHhkOhlASwSbzZpwyW6MsELVnaSVreWaP1vlCYO2No60WdkHUYSjpZh5CdYy
+6wJyZhbJhBdhUZY05SQo3X1fjMXc18ai2BZBMv4IY7XxmDuysI61C6lvs6+df6n
vA3b7BpxhcuptG+DXaaN7pubwMFZsoJmGB1UhHjks1+Bqh0xwXYagrJtlOpWyKcV
D2c4g7+FCGJge3Rmt2X2Gx7bZ8qQwoGURkmETnbEFIeCt326NkgD9bI/CvrotkkX
vf4DfYAtdWvdIGZDDYkmKZ5RKkHwqoS4jB2peEQiNhPItE4GdvOKE2HpJY1Bep0r
rcddvOO97ISOeNdzOBLVEZ72vbKXfvnIl+Ik3fBhy3enNk6j/1r1MtqiiSHEebd8
466BJ3IBARaGbzh7HtB7b1RxGdzJppGkvlDSbBs35ICepF4MQfRzj0i1lEYUfBL5
SPn8sxkvkIWoluIBDr2V5tjKYudvR4toVuQVkTfei5/nRrT5WgpW4rVZkZxNpBfa
iUo/6tadU7THBJcO97IhSsv+NHPzTYeXMyUhOHjNNvG24oTAUh0CEBXyBkrhKj5Q
XpF9W5QPiMfXZSamJ08Ji0ORjH+EL+G3Jy6ZSqTp3U+nqCa2OaOzGBwE5f7pv1jc
vzefkWf5CqZ3HJ8J25rD8FqQcYISBhYD0iXBpT5RzRrWkuSKxzCnVsHuJszX1lsR
CEAzSiM0HfowTIEJTjq1jYaQRMqFrl1zvRxcPeo5e/Oas3R/jXSdmbtnigrsGF8M
QDHBA8rXY2ubC0kybvXM8qc9p0fv3ckq0vBaQbhXHqxwALALp8vVYsUbh+Sgl1xd
UQqKZTgXyCT2jjbyAyTodAmcdtFH5B68tK8BkBNCPUvqY3v8Lp2glasBz8TaIL6N
pl7rF4fEiumiiMrULRQi1C/q6qEdFJeoZCR1rGKqvHUzTBP2gCVI5qUavBv+wiQ8
I+WJwPcKFJ3wPpImFm4SazEwQtyO7ZC8+k1oydxJjq/Fs2nYNA9p7rWi+KvDL//X
QpSKAwnihF0c0vPCrY6uVdcoxoDYnfd6GPmFLgYliOalCAb3rLhex681TC3XQzL/
3IM6gT/EMTLvDIjbdVzGrr2CCUXXq9ZTH7Ueh3M6tZ3S3i1YzbkJgjN0XwIxFjMi
1G/vAGryOzO8WIORzjjXbaPVDqy/CNckoHh4MP7Kt0R8O/jXg5iSTJU6MjiBPVDC
+0B0/JRWy9p8cPUE/y7XrW4hmz0V2wx//X1Aa+qmVQ3nni36H+HbYfCNEHyDlIfR
24iNoZ7e9EjbCJHium8INwvZ/fR9HxYZdT9k0LGKfzJ7JHSqqFvOWz8H7cVCu3jf
hdlVDf0Vrkb7hX/2rs+HdPmCgLVM8WqfJQS8tueJ4S5fE3yZW5Sbk5S/OHDG2/my
im2wri93TFgg4RZ2yzSAfYyGFcfmdv5jUydxkYLG3VLkS8h/2aiWM4/fY/jFFQXm
/6Pz2xVrv/CMfYYpuIbrfdZxpgTLXY+FbR1flcGkU1REQnIuNf6vJoKGlczMmmkK
8K/iiaS0JKZ9sl1t++c4KJex/kiCbwnM0dQCml1J5egL8DxWIx6SmOVTSfypbg+h
Oh48W6iqSAzPYfrBzA49CkZdwabQMLJlKY4CKk10cL/0/zCqQapm1yUkDRbnZvVx
/ZGwYuZaczJW4G0Ze+4N8U4amXdTKnDUyZDdPh8BZ5SDi4L/9D6iq3FioSYIw27g
Jb5c8YR/YRD60vSlLw1Sj9B79Q/vfbo2gJHMB4yj7YNvTSLJkyKJam4RhHMBER4R
MsPafaH8KR4+Mwdr424BPmZJMEm5M3EUdzPG4EKW0ZQUhLp9o7IGaLPY6Y3FnrGt
8caybOGeXKSaTScsLMBwKqUBLX5N88bqijDWJ1xwKfvY0uiTN2mklIyrJR2uee51
EJ5j6mifQezJXb/wMX7miEvQs5FxGGTJcDeUOxYwz78A1yzl6nWaMMKUbYrG2vnM
v3bCbe3SSFmtKwIb/KUc/bH3XsEWAVYBbaYB3j53BYu7iA3s/SD5MnE0X1s570s9
BDhzlM/qGPiXvJxRtAK3TeipqUrA4Ul8IXKB7RO4Zq9T3pwh44jya7tNq8S5WPme
2UzSK0/WASZd3pGfCE4upKK29ujnyk4Yc0KcsCwC+DsjiVzG5oipXaNsyuGsRmum
U/1R6hoM30O9FqxNMAd5jDrQIojdp0+s4C5AvHiW2jpaWQEPB4Xz5hEto/Y/YwRA
HEz8+wPHnAiMhFS6OR1B6ooUyHsF0J5OlQJaWWzI2leKb8M4uA0+VDU7U3V6CxPB
luWyOIN+WAO/uy6SjAyr5QP3mfUyk5cQutBAmBhmsmVy5plACZefDssmcU3Dg6mH
Zi1Bf1IO493k6XYvZJs2p1MCrfcz2CISN4uNQ+GvF+ww73/LGNWDfn6FBO4QFbUo
z1zcVvLXTERHrYqJiNKLBdUvTXKM4JXNC6x/PPqT6YDCZLI6spz4DxyaMHo9js3P
HbHKMnF5QNE0Ktq9EQwExEXwOAncgfi3kIfjUUHQhLVDB0MgTDGRjvWru2KWwAg8
YE3bVilDI+vRP2sGKlq3llk86LrYzD+xMpjt7zhWUmYYnY93koHGR8Q7I/ktAfVS
z0vBWIhis0oR45vHmh3GBeNgPH4zkP6/8nGoDvadOLUnVWthgMewzP9FI1RSw3O0
IY/fmRpPFqq51klkZbdVlzQc78GIt/z/fso+OcpawocTlbS8a72ZzBH+wW80Q898
SYhoRlFBYCLGy5ECnJY/fIY6baNqcI7+E2cW+OEgPAnYiaQ84M0jpOP9hN2OmGrN
xbUy+3VDFBwXuyJhO0MhUCA3GRXZEtODS4vdDiR+loMuOdeir/8JKncJIVU3YIla
rVjKAxEwbQd5FSHfXPHesuam27JHMt6qZtbquTK813yV9ADLirzBgiRqiFA2CSXx
wx4pTCcQR8De0QvZom/j+8vJEiqtNh8KbPclzQOBZDbcpUaZoZYJM6+bgoA63ELN
oAEbqG2x/RG4yk0BGqNgc7g/puvddDK2u3NdUM4QPRD9FVCUpiPj069rShKwWUDa
SgzxNvF8Ry94DPxjLE4HKtJ4SOh+hjeCBj+ZtU5Tj5QUQlp7xM/6ZwKy8TV9whe7
9L2qlASmm+vrLPIZ5WnAWTSwz207LyIGkOwrTKx890bb/YLSuO2XgvuGd8ExlmgV
ElE0+bvIpEGaFTkDJXFIvkrSP4gUxoLGMlPzjWT4fNFkwoZuI8JKeVHMnl9VXDyG
Tj1pJHz1ZbrwIYnanIYVBUdGAuDTf4a2jAJcTi/511bEyAL05NyA2yN9kmx6vlA1
SYL7zNqBVoKvD3+5PA4VrlhyeMTzine18CqT27rSRYmN7BCWRAXoQ45AthncmKMZ
7Xx5pvf9iRd78buUkwEb4MQkSD8m3oBIrcxxNomihU4hcK2mdmGGJY6Dnv1gyGUa
P5c3399pf236M/1qtnpLobYVSIE6kayqg1PfqJ0L2xsu4ERQkgU/uVMe2RBHK7qT
BPr5ByvIT/SGGyqzZ1WqjdY8o8ma31jScnsIUueME+uuaMLjYTasoVYFCDlcRIOM
G0hRb2i3d/dv8MPUtYdZXXhsqEmjb4pk8KmiQV9eNYL77kZpTDqBCIGlpvuE8m7W
Y/SuOwo6MgfjAB2qpBe7DvPkhluK1BPTKgHqyKmaXxFMrT9ZiPyKdH1CbxRWTq2j
mYL+tZz9pcdDgQvbbkOAnmX7cW8gci1W4SKt7hRCQvoGjwmOQFtSYPqiRc80WtWb
QMpM3gFh03Yq4S5I7xCrD3uc3gVOBf3a36zpg3RE0YPw3YqhYdbRC6oiiwVgRykG
juICaKGmkMHLflqq1tpamTO4/wFcad7GEjxlRGEXvPSYESNf+aa4FFkQVR9Dx02u
pCnoSbmvs6jl1N4/okL51K1N90Xj5GGLTnANGOswJ05lSkUD162MWutN4pzELaVG
W0w4P1XBqzjn+ly+p1lfCs6a9RIv+Xu+ECB42nyuMke2Bs2Ern4f3S3vI28ZRFvG
Dj/lS0lWbocceDTiaz+8B0NGgw/Nqldmx11t07SLbuoJLkHehdQzHU+m5PTefzMK
Q1M7LSxqDxqRtm3mQF+iHlcdmlxzMWSAE1Ui58grrBu16Lhlh7cc9i5ycTtJJi/Z
Rn6FTpVaz9D6Qmo9s1pLqDvsIIc+Upt7kXA5EDWRojI9j/lwlVPIq8frl0Q24w9/
5M8NEsZ1AeOwApGwzPOuIzdWOBDvA1dwgNFPqyEQOv/7GMbfiyA7K3sutJ1PKiPb
zIO+IASuI8oXdnLiqHteegWw8pqOUtj8QBdSO6liUefQTDKCT7qRN+gfwk+PWdvU
9jHJLJvPLfXJ5gq3/wJVqbTVbs/XF2PJxMcYBcG6tE9kdH6qLogNEHEmQuUkqAu3
J7oz2GYISgFhCK+vrzAV7v5/CCQPXMhO043pNbSD+ob5GO/dJH+Eq4IGqJepVP2k
xjLDlvU1jkPqjcurDKNf/WdSRjCirvtHrRROXUBw1N8Dh+XN9THVYIkONOIEA4rm
m1IQSw1u5Ua3k0KsUACG1ARJVzDPh5W9KtvgAl6pP+NnQRzLVx0gnhclfvIH1ICK
PIdNz893XJaJc64qNdTTY44j/rdSRv/YXXPg9/PL5AyDDjOwSnS4deIFITWnIU+y
ONOS1s6UTWGLhPIA6EkviRv1FT5L+Zb/mMG5u7v6N9qRaC6C2R9ghn2/yZpLHcRN
q8KokO276U43WAst/wreYBPE4mOHzGVQLkGNnZmZPiLQZ9YJrviKL0yBPgG8P2P4
2ERj/GC1pxgPd8EPtjQhg5lI/aSD7E983N/pEVCdEHDZYhZzO9rROoz1/CBW6UcC
NhlDpYZMtVARcOsakFbPn4s/p2xXIT2dkUoaA7c8GmM=
`pragma protect end_protected

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
bP17pCQajFaid5dhfF9CCwAOYLdLUFuWa3t/wys2X+aieDHTkuHQjPAzpbgrwc58
SvCcL01Jm4nMrUuPEjQ6bbVuDYK08Ovsp+LvWbNQg8sYbdleOQMYHmoRYQXPqRyL
cal/FJynjDM4JSOMByH9XPihoMzuqOVXkZnTdmn37NM=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 2042576), data_block
el+hweEeLWwk84uWnhgzzRfvzOQdmAnxNegMS4og0Ci6Gcubw+GA6IVMeoUkUXCS
F9GTcuA3hVVmoxL/cLdVXIe6sCY1GMQ2vwr6XIozahC68F8mnxEAPSJpUf/AMRd7
us8FDreAwfEyAwHma8O0O90BnyCCyQo+jRAMUqg5ym99GVeV2KG+xuaAEfPBUt6I
8Q+aOcJ1t1s+2esjdpqgAqb1KFusCUBKC13fw/9fhkUkTNJEUSh8nu2HE6wM3b6z
q7DFeGrSo/F9+aMxTOovsISWqwBDsqp7l1HbqXrV25FBsufj1JDQbnJjsJcbM39J
qXw2RGjjgsFjaMNl+IqUGyKXPi5PqVc4ZLZrsFNaCQp+UGwEg/ShqeHc5NtbwNR6
MACYI27CXzuBl9IWmMIZ8cgMakByejxf4oRdDwysFpIFDNTu5g2XTyhtAjYkNMMD
XivK/69G7hXI57kniEVN3YNPt2DrLsGWQehbrusEE0OiEnveXzg9xLEyP+52Exa4
cif3qWdOe4Z/zjxDqxWRECzeFG2jBDoiG0wZ1WHEId/t/v2ayD82DM2aIDI/J4h4
/j2gqOMLfgAkIB3iDCMtz68c3/9Bc+WLl/AFvhivEXtArfEu1Kzda8HP9pnEhG/9
rPplZwFMnKKcScAobPBXT2bMGBf9v46APg2J5WGoOIbVSRZ8I7Usn5c9jRJzd4jx
Dod27Di0YgfIaMel4MH6tysMNv+tDYv1ysftPGji2oKfjl1Zj8lQbpRS3QI1huwH
PaHKjP/Fixg+f9PWGYpvZX7VNBFGwFs+1z4eR0NktKfo5A0ctncw1z4ErHcFS9Bz
DyecA/opff55HvEKCOw2CcnRhdNGN6MXdwDI43rF1z78Z77uELfpwNKSUo5g2kUv
iWCG/EoqHjtVxMA6AKOWTTy8qeSEUXHQ0+TyGAYkiwxnFDMp5pgbRjKI+LY/VWFo
jAk72G835eupvPGUgvu9lG7wu0aUjLbr+zQq0qh1w5+KWXoA4jcdvLrLKoPjG8kU
ifUp4yFg3d0zLB3ICCjSg84vZLe6wOR3+DmCvUbNWCVtUk3vWSwqBHLO50i5yjAS
/MvZzH1yHzUierX8PfXQLo0PUUWuxvh2Zoul44SxkXlG2xuCf7w2FdRqbW/eiwrb
P+Wo3LMqOuollMtbSvgGhVTBJTJjsw+vbcLbafxOOuUw+ooq/AlZT78A+SrMgFKH
BKDkK4VIDVPu7V9fzrLZSQhr9Fh6XahZ8XHzYD+jwkOMT9tc440JAQfdTnNFkq2V
y0OMKSKkSNHkjNqFampx0AmlCBAqda/1GrOM20rZXzBY38JSfkf33QLNkZZkFgz7
26HDcu+/W6cKyonrTXv0YIAHkx88aECKeCDfvjQb3lCs2xZAXCLTr55OjkR3zXEe
IqIL4SDH3/6xd5zS/AYR1OYpO+8qYT3HCaZajJ4+CfbRWsGqcQK6zYIN+AOB5kfL
gati7EVPm911u4aUd21IetgG33B67KuhZ6zRTY68ATEjk3TCGH1M8e1hI66SlFdS
K8DSFUSlAdximZWfNbxVzmTDLFHJbs6lnTKVGhareJEJC8wJkAjPZE4SMI7QvM/R
zhKC5U7FLYvDpPOYsNG5gsdIVqYWaS7D6WbymGYNSHmYDdUrT67H12b6lhfOlc8N
bx+Njrf+GPQQLU49L6wzI6gsiS/BMMJRXvBdOq5cW1VysjmU2Kbzkhue668VS9Wc
iew/mdpm9LSooAkemdnhGYsKs2H5oKGgqHmTYlRXMH64FYmnHz42xLX5TWwb2X+J
MX3ITJACZSJTvWYMERMZHT23pxPPCz5aceJ/KwXRfqbS8D7JNvR1jE0S6v0hAFy/
Fau+EiZYCA4XuGx/ajF7OWnK6ugeqylR5/UJAkHymUP9ukHAT4ookCApQm0sUfNz
WteEbT4IHEXE787fLXIDv2Y/NahOtYNaDFPM7AaS0neEernoXN5bzyLwCFcuqVyO
rMP+Di01PZlLoNVoWjg5H7fN6+jKDyEIoMF0DNr55a3w5iltIggLl7jjPM88H64d
UxtAAvzTYHcpJNl4l30PF/6B9qms85D+U8vr6qBSTjfeC+tWA95Uqv/1G6YA2cuZ
/JcFo0e+gRTk4CQ/MJpcdiRhO1tSr2gGmBXLpSCa9DsuNTJN5/a2Cqy6iQ2tg4oF
C/1VlQugQx3walholTaMwUNHG/k1whhGLWLw0O23Fb6qPyKDENbz3P7ZOr0IJ9BQ
TmQVeyxHDnDjDiEPE8taHZTQZ2Yn9wlQiz3xV8ONe9Inrt4T1KsL0xttj/uWmt+2
To91MERrQcBG6wtgSee+/Q0mPGsIakIZS1BIDhpyfKrDjoHntOvE/dwKXMKmkYG+
js99SNuFQLy+rV+7Iq8zulOEK0Lv96qQTUC7B55XZ+6ESIykfhbyhq7j/vhA/geN
pBv6re/yYdiysrfK9fqxh19zKxNfA4GxJtGeZteiIoqTOl7mAGgpNGBUZ3StFrKS
6hq/KN6RUcyFcecwZbNTnggEydbBjtr0IoPcqt6nz5oxBKVVqBljdYD4rGuSJhJA
/bmU7RQzYclQ6RijFyEMGzMQNW7W11xxQihoOgWKrBOOFxQhzYjQZOn2jLPivOBa
AL4ydrZX+sXJsafJ4FkUD43pAN64rp1dUMD1Njdj4KtyexfxCpZU/KXoyCl3CIHR
8wCneYaYbcsdM53jgXh5vSZge7Yldu7v7/dS5cZua8YgISeNpaY+bOQONsWFxH0x
YaC9lBCB5aCuGaE1te+2h3foN6A/6q3kAAIUyp12vTetPXL1eYB3XduckHpC3MLq
CPxmTs4Lw1ZGI4epOt9TVakPz2EProX4NtFXY3CnOq7SCrxTE3CAAW+mcdM/a91W
kBb/VkdySFUHHLSNpDwi/9TGP3IZRfcwllSy42fqS3/6qkfFnkzjXHYHZDinCEC4
GW8sHTU2PB5FCQJPkKidPecF5LHQh+Tow8J57mbsKU+aZpll8a5oZvwXr/EXW5qV
96+KGZNZmOwthw+grO/rTOqB0FdGX4yX4sqYHlX+Ea1SiTxI2lyMFQig8CrdH6/v
+/Tx3iwtKh0Ly3ilJsAObKx57ztBV+Ds616EQif2Tuopx4vHgFt0NOag109BQraV
Z8jQ9EJ7sAEljsxYv9t2iJ12l1v9xeF/FCBjfJB+5jTvO0aDSI8Jxsjl7maKyytb
7x0NG4Obh8U/bRX2VS227lqn9IliknIo+uHFCxA47LAR0qv1cSsHqoXsf3NhDtlz
95HZpZXYlakNVSfhEAUWzyI0+t9Pw4cWHMDsPX6w5eysg75+wc3yOkr+0E1QBHJd
ipNVcaoUMlY0qCny9FKwfDbxTJ7pBxUAD+bFKm4Q6vM+GMD6PdPCxMKk9V9JxN+k
S0lpINiLxlnvxrPkhzRqikIO5YGEWH7PDYCuUhnya4mJax+o3iljv1oS6GDxB0A2
q5FKajYtBL794aJgDlb2ztljhWoV05Hq88rjZ9uZEsF0fMTouT7H0FthC+5p0UAa
fc2nGA8T3Pkqi3O8MBycfNmTahE7Qi+yk1qIqP2norqrpwh7LpJuYUDFGTMcsoSl
tyimimU5YqKFBFx3YLtDtKk9z5a3kZ0vMWd5aTNgUIhX4l+ltnVa0arA7j3e4Uey
xvHugs8SG4tKnXYPcaV1q7aX860Oh2K135RhCqdzqVPofAGMIFrlFLq9a5BsuWlB
wCRLvaGrFcluE+dnaSy6zcYWrgHnzLYr0GCCLFMdySF+Gp465dBhbPa69Mf+6sFS
o4MRcbaLQvfgfQtoNBLa+kJOddi88OyB0nOqLY+Bcj76aJtmPQtCi0agn7Qdpjsz
Xw4pxBqdfmrhy3w0pgFUeXstCULhH3xZmWITaxY0/YyGczabXcgp8Ezr6HYk+KZ1
/zhmiHIzm1M6uitVJFqndlsOxo+xFl72V+qbUAii9GmkhrDmYi5LPezRMQDaXs2f
OltiJnFbTXqnN7c8oxStajqOxK2CP9IAdEbo8zyvPf/3MIPL/ezKfxobV/fSmgDP
aHBsymmHTP3HbuAmZjwqUuOVYm/jY+1+xfcoHJVTWmWNmHHh53j3fO8GdoQ/nElX
kwze92L/LG0GZgviv71uw/5vHqw+CAkiJPh23pJBO6KFxb89RG8iQFbVU+zXQRAa
7nesHO+OcEaQofkM9gGXu1CndIo8r+4KEjy7XAMNeGdvLVtY26wvil6N0FVnJph0
hJY5L3kQv0hkxQHOWItVof/6+H9VguFIJ97ypJ2MbcjKZy9W/gRVdbgaV40ievxe
iRFd/fSBOyRxHkpxyyWJ3jH8cZyz71S52NFNviAMeWrDNnGo8iUQTfBYigkZEzN8
RvU51aBvzw/wpei6hVrAHUA7xivdIa0aW0Z4qbTWi+b9NtxnMUVuPxYmJl7Xgxb+
1LmjSQBakwS5XhCURDuANNhgvOp+q5toFTdYA2uEeDxj/wo/HN9rxyq+KztCMpNZ
N5zKxCPKFp83QYQnZ/QHZCJkZQIliJz4Pew4pFbTSIwjvvcQU7quw9dkZbgScBbd
7fq7PNJ991tUdaG4rlgwpIDdCfcHgThjJ03EuKhYbybAGAdptX0R7qRJTI9z942H
CG/EKqJq/ZT9pwiDziM4ak/qUqdN8YKJmh1wDkqhwU5O+mNNBD4ZcG6waFYrohd/
6VdDe0KiNAAiXX/CrRbVL42XDXFh5KVlEgFslxAaLUXfYg2mJkLLc9XTzBwuSzBE
focU5L3e5Dq/CORFqmIo9dmh0HHHPYmaVuKI3O7KRQJ3ZIi64mOLS2HAfZ3o12W6
3GrWLBTZBAB6d/xrJ+QpI8qE63cyuodqM1s70T46LWCzCcqXQqRSTWtdEH6fWxjl
9kCbf+gNW0Ptx7vS8XATA8jrTaaks+ulXJqe/OcgXyTMVMzJgQxHetnJSWntmitj
K4/RIVvU6aobSwIzGJQgm9ZXNYVA0eq9ImMLY2tjKN4HwLAemp3gkajzkgYfJiQC
1LrypyOKTTkcAGnO5cg2t41SaGt+joN3RfcQ3y4FZ8RW7ifmYRs21PHCLuxsEVp4
coUHcDQvciXFoQ6KF00wgUPVBARM3S7qZ3qA7aVXIAr3MxFbeZGsb1gTYNEVE31k
Gzap49zmqEwQVzWAXseJjFcYkh8GjDpIZ51IM+2zf8jseZERlizPaQ2wmBoIHF0y
mDH1RVagoXY8JDdStfQuYatehKtyv1bL9jbNvUFRSY8hPPX1+FLDsJv9m7WE5dnI
Rs9sMh28ZLVDzdPLyRinvdJgAFfpt8IEvDIVaCmteFwqC+v0ln5x+oZcWi6fsHDL
6YecrrpFpI5ZEgmCPIKxgD1kXoY24B/yBT+R3z9KiT3ztt0kB2zs0pavdD3OPNzm
J160l2NEJ/b345wKqYP1G3ICgsE+M650HzXNPAwGwt2dyomQmVg2s+wPGAHQ/MSg
1CxgDpt6zFHh957W+Gkzuk3VoYuFvVW8X+nOfi8JZXxvhGxjY1iYC+x25x9KptM+
Rtv5sP/nWZjZ1dvpNMMxV66em03p4VW0wYGbi6ErjIUzhigep0XdA3XZCJxPemed
tN9cnC9jsHR4zvy3Z2JJepsdpV59vU3+hEKEksIHmcyY01Aa6EHLw2Mg70rcObK2
IuuiqRtOw2TYIl2F1i31B2jI40JSQvYisO1HctlN/uKf2Zh/5bDf4FvqlscRCk6q
duRfsLifqnnbkCPxz5Zq5uJNahbXbHoCwj4khXE4bNEtIFze3OUdT4DXNyA3WXbB
BZsNg6IneOz6mhNkRBzCOKTJ2SV7pvF46nUPlNdqkfgz6trGFQozMZLGCHq275/N
tqSILXbGJiIkecJuTmmcuWRh/5bQNnOrXcTtev/YmOn0Jh13O63YpdI4jJ+y036m
Dc/deR574hOZqopBwB+0kV38cwW1RXIfEpYaa/7dwyEyYJ9raWSae1JPbPLG4tgr
jlXYvPpx2+ROdNJTYcsQS4a331Byamqlh5kSyr3Tnev5oh+JJ+dwgBPloGknXgYq
2KYdMYXUr+EWXareBfg+oF+Bx8LA6HZDolB/w1x81zuVu6DP2a6NgyB3D49iiBJb
RKRzhmxDJbC5a+XTjmI/8l2lXx7MlZ2zKRtkazA+lSFmEonCMXycgdLnYI7pP9OC
X9fyxCt5EFsoAjUyKxZS5cINAFPB33ywI8Gaa/+hXZAWOkU5lIDsQXtpRSvo6Hj5
XDTUvmH4lU3PsILyL6c/6ZrEE81OANcoszruYWg2lkGvAOlzX84+rZWNJ3nT90ur
CTqKkqJI35SGWAJ12kdm1nf7sI/GT90U0eoZtP9cQuBVujrd7SCD95BlKE6OCZrd
kyZigq2kZIqKSkLugtwLO52h8D8nibXr6AoL6AicZQBTahTn7Y+3qN3Er2G7z83H
5WeoJzokw1nChliXXWd/PK9IQ2zyLCSDKiGX+8CxG77eNmfw+QQOp9T/xQN/NPTZ
SB7LPHQZ5DyOcD+Ta1u3pWP/a8zshGy4mktrgXmQGSVwNhLaBiwijpMgmyJPxGjH
KqnT/oWgZcU+uckV766Xu4mAdUD64UCZYBbt1J7z2qSOPonhtyll6+0HcInE8/Rr
+SrBvshsewXGyuzFTY0FZb81oB/tUll9MhUc0B6cszflYTmHlSj5Dl/XT7fvM0eg
GEcAajcCsbcST7G1r++0WsKxAyf8gTN44tm3d5be7nBKV1eSZxe9sjTcr2lY1f0I
LFQugPPZ+9pyyVJeVunq6cQMwOCi2M3ZlDOewXJQZXzTgCyQTOUOWmGR6YuGTcSH
k5MdYTE6qCbAZLLYzY6YkXzl+fTEA1kW5iZSstUlo/gbV0RtFcVU9PfxzgSiHXD+
EcSCBNu1VFlMqCiRxyMuDht2ZB/UJ2LPKQhHep8dkAeFHFHcwtpvOqCPeoUtDDAX
PpLEImz+0omC+RJJKWiSxdnSV018iMTo66DaKj/mmBuT0KKdD1OStZjK4XOmonOF
lDJisyAAxRw4Mm1WXJi2O6gg5Q2ZqDRka4FoRyiOGGfNe2yBen9HnhVtGyhSxmqp
Zaw/vInxe/PhAjFdRTv7L86C87uY1vIq0NwYD8UZZYNzEPoTHgiCLqdXYPvZt8Y9
kYzFZsSlmmy7VBKGIzN62mPoyi3IC0+gJ/p3oGf3RDU2PIzJAIEWtQM26rAhy18j
o/GGQYTAZFSSxxDGM0AI6EVlAGhFVkG42Qv/u+wclLHMyRRT6UJELjuHTCGcaIQB
YkhrFqMUuF1FGPUJGkQ9mBqAHim4oM6F6raGWEpgAM+pGw1EZiXrxtNt2R4foJ6z
myqru4VtZtgtjBjGsYnwLrDhnPGvriAIzYhl4larnVLJGZUKsTXI2E1eMrjFIZbr
mceD2j4nNwKicWPNlH1Hq2VBDt5ETWqDtN2DRCcmLU4s6EX3L+W/gyM36Kr5+DQq
6a8tqLx6CIS0Nd4vB1r/pG5QhlAWpNv/LuriOzccqKfcOotv6kvT4LEOgvayfN/V
njuEa3fF+JhLw1el7hBNYuvXDmgWdQ41eOOhh9Ms8HILxf3I1EkPqNSL4CGoOYIz
eR2XDH9+yItboOJ2x+SxgzeUKo39W0fe//6ebRWTZFike8K4JYL5fOq3vDJbjIaK
/Uu4BCIViF6AXx8w0OIelJRx8rGnyDIgRhT3DeJS7zdDQOi/jdcxxg0iRbiC3htb
jkdys8jYH52U/KsGy/InWCtdMp35S9PDWLRq/fJbmDlmgzO5gQRfWPV9D1pA+TWN
6wpbMzczBhEhkVNPxhyheFCsaanTgSg9MY5ELjjE37mpQGw/Hx5iziwLa/jurMoP
2NeXvO6Z+U0jOIoOhiaWO/v8Y09p+c1x1xWQchMjHbHCGk2drfqDG/r6BnCCZQxE
6N1xt4/e+u+l68mdiWhCDM1YxjdD+ZDL8HQSzDDhgNJZr/wF7HyobKVKAXIqLqs0
V2F8wJlYUQREVWFZQg9lqsriUqqjzlZYKHNjvm4vwiVndY4BFT0NgG+QRvxXnSqC
Gu8QuwcNO+k/kdQpxy6UNeUlPAxFevGBXcEjvoYYL03DRQ1B0tKBZFklWmX/sm3I
LHUNgJDdKnYlJGnRZ7D3hGzb1+AHO/fpCbFDf16ueppiow4XorfhHpLZ87BNRBd0
0XFKc05AxiRqgTpPyugefrnCFVpqnTGBBigvOwwQJQykoHwooUxDJUlxtv9DtWCl
p8/5/piFe9BU7ZJCHaolMwi73i3Jz6EvutXS0XY3gOT0Mc8Mr2hrGWEsV4vTT9zn
11qgkQwWNXcdrl+TGeVwO3I1wLC3lHkMp8Y73ymd2k6wiIsDSu31pBgkAAraZqAe
5ExVMlNviGVBTa0L96kJlgc3BTTWLTEVvCb4jWVj4VDpJVjPsqEAfQDGM2IxnGc8
kT6FUgK/aq8FHP53vmst6cB+zXRmFLkyn6EvRCowL1vho5LpYB8dB1tF/tTXTPv+
B4IEnjV2ZZjK5IE2ueWJ+pBT1Dov2XEtwlBXUsD1umLLCAxcLx0eRcuomHzN1c+S
qbLJyVjGfLd4Wx25UcWBJNZXVcRy0darq/OYJmGLahID55ETWama8dsuTv3Lwfa2
Pp1teFuTF6kBVm00o4VHQHA0q+/g1ctE8TWhWKFy4+HIwOQAnWGQv98XBaCHeJ5l
p9DM5x4agUIRXE4kkxp44nvU4H6Ham6/U9rA+HsF4wXLX5Gr3KnKxYTZ6vH7Ncys
Wl8vCvt2LDebCr+JDbCFjtSviRE1FvP61ZCWcnQL4hb/nznT1KxQNaHhXq0mg6YB
LXqAxxnVBwttBLP6hgjTXvNlP3o/IDZoim8tsoEtWsmCWIjnj/ZvOaUCwj/k68uI
gn1cYSyu3WmslQmPBbvsszLLO/TmSGMYL9WQRIVgc3YPSAc4odAgVnJcCVxbTrKS
wCJHsjhqM9i/BCq76Ed4PgWRk50NZt8VPywOVOwt9uPyqIDAG80WvsKzKraL9g9t
u97KauqOovLKLlO06Th7GIktTnU0rzcPbNRu3cFvQt5XBhYOSBA3dGJkpvBsh6fn
UyHKFoosXGW+yWtMzp134BSoi2xmW1b2x+clDLuqlY4k2+Q5sZ+BzELrSznJ2D6M
eEB7v03QVKuNYwDdg9vU9afUa+vy6EnouLOkw2R74AqyhpVqnQeYvu13hzcfykTG
0+ee39j2a/6oGTbUWiWs9a5aHPGWDe03lqeuOjU3B/A7yAP6VqCd+V1J4K4p8YAi
Icm9FaCZOMQju0lW0ObUrgy0TOoLldPCT12RrvB9AoOw/RiVRAZPmPO9vEkc8EDu
KSip9LidnaGKUwcLRZaicad/XNQkEUD/FpkJj3WTQOXdUMQraAYHtV7xiAN6EZhC
dnraYucZX7WeotjKYjp3gxHgmyfFaWU4oOnKrDOqjprESr0eAZJDddEgNOdfIWPO
lZqGX8974EFImLgz+neJchNld9wG3ydSk2tC42mT9QmtreDPAJ2v1tuyqgm5nr5a
mxxn3IuxZIEpjd1AZEfLNAcgsgt3pT2z4w900YPNGSUJA57oGOZZAFzqUbuYv3iA
DpwJct7DTlKaieWbnKkxcIfRwIody6JemnAQLFrsQfIIe0UuFGgj7JK9pWq6D0n/
xTLm9TOQfXmT/8D9v6LQ+LrajRRrJ3ufXLoGbvmliE+uIqd1i7Le/AqY1ES7jnho
0xxgWG9WXYBtfK3aN21nr5vnoF6peLfM5sg4PQD9Yi7Yhzsm4tUT+vB3tsw4gfV5
g3iGMzUBrUfzkVbBJSQgyWZ9mvUL38Vstq0ERtxzUHxZK5g7FOObY30iTEbIxAp0
mTZDTuzigTYY3vR0BGUe5EQdX9xIjVYIaFMYuSfVXiN9fIPpDZjGSUTd6MsOCbBf
MsEpt+SN1V15HbkGFzzQxwUPLDLDSes1gwp2PCqepNsOI4pI+b4dLtW483MfC8Dd
cY+y1fAJ3o+FVGh/1ecj4wnI+LTGmdKHOpXCccXCNvw6wW7zPdlyqm/pIIKoeDwr
MALyexKyL/hSXCDreUgjjDaYInvTf4/Xm0PgobjO0jUN2cbkwCUS53fluGfzCs4v
lJ6HF6B3qfn5D5J77AdW5YT/O34ixLmuW0lr4iErWfPChJP9miOE8K0Oe4VVTAHa
DL2pSXmt6eqwBX6p+jQXc9WRlf+p90HY2Huf1eSR1B+xbWcFhsvbMuu0Y+w2sQDc
O6o9E9N0ni5AvopWNdJgOtOxUer1s6DcAoK004OngYS3PwI3odj2d7I5AYxCmXL2
hPIFjknZQueg+wQxdXUDw0y7gNnqZEyEpWFQLUP6EX1NV+Y1QS+kx66nOl+PbQGr
AGFFdo6+phbcKn7uq8TzyzwqBx/RCjyfWZ4Fyq0wTj8pZ3uftoJe4KfAOoL9ItKF
8Z752BgV2zrVGNrBYRwhc0J6BKHNGRczApZPLGREX1qXn4sqovDn4JZhKWzM2gSo
PMt2s08j0toHT6Gm0A/LhwSiQRKE4IFIpn+SMo3HYwZmTdWuSpSI2YsBU2WJcI5C
vlFhn8Sg21tJaGWRWMxHyq9VYMl/3IUXi5lMv5RgwsOQHbnYkzVhJywMik7jW9ue
fpP7idzTg5MehCtcjoplFL4p6KH6vxW/iW/K1H73EGmUpfUsYsmRWFns2ofZMFhA
7LrIFf5zMcbidWRp5DjkQOyCv10beqchXdSgUoZcpAazCGYuPe2zZRfMHYQmytDG
91+UTj3l60dd8zMsKN0yeQWbRDMJYElN5DLdI+KyoX7Pe2zTMdOCbmKWIlzfRAbq
V2jZXgMeDqXd2cDQgNhIWP3gF36XNvPUHxM7P6MkzXlSNnuLJAU2+iYIy3q6DY5P
5QNm6LGwxBNbJJrEXQP8Kfm/bVh6DAZs4MCemWdJ4ZEqvzSZ6nwaYbIVnIKP5ItI
c0dVYqi7eCUbrEPusixhFiwDipgsrxmkDFfC3CgOCdn5cK2PU9Ybnx9pX7UwsfOx
kRtleVql9K5zIZ0ytx2vVnpllKkFeI+YRei67/NurnHbPQYdy21dmawZ7p3Sy5rY
66J61Ihs7WuxyEgCb7tmWFzbg69f5DjM7wPiEA48DB2/xieucIrln6TtGz0ipHVy
asbXoI+PO8qK3FOPgNirzc8iwzFz1bQ1HVI4HplAa3QeBnikFD9vhwmytqf6htpd
fmondnerC9fMlLi9FR2FbI8QpuIm4UBR/0J4A9PET7tbr0sslplrnviu3N/i/G57
8T9JP77lrasSXVhODI1MaUs7Js4vpFMJTiqAtqMWy0WW44NeOcT9FAiSDlPC+KT4
n/o76jBW8Q9rpRrkP1HKXgYFausXmiRvpR68m2EITxw1ucRMLiy5f/vJ6KxboGNP
bp/BJcqS4GMSC3nI61SYtsmNyniNZBd8lLiMD2cUe6EDdkuY5gAvM9OZBLpWQ6uW
4vAH/osXC5NHmZx+r1Jackzk0PsgLNxa0rLdqFoRMvHrdsBGWEu3Zi1fDr5DwOCK
tqbrJCsCcnv7nzHz8jyHwyYPlNctpCfq699tAXkp2ZjJB9TxiMwA9EG3kpXNk12A
V5nt51wETl9OaA6/hytS2X0AcWGKRJAwRV8Dn1aXObr9N/7TmhkiCW4JCIJL206M
fndL5/v+KjsETRySpbX02dzBR0eKxV0vdcuIE4Yr7gkwgmd2/e4UD28BqbVM0zA1
wodjN2M/HGxyak4xZGRW23gICXLcIGH/GXFMHxqBYhZ/G1dWaEqolJ6/2WCFKwjr
CoLmg/3l8bKwTIdEO83BLV9mePdvaqQF/KlBjPOcb3XhMl/NAlOMeJq4oX/3d5OJ
yKNHXkOLnAHgPruYHoY6AlaFxnA/S6Wx28P/6lc2BwZ4JQazYe0WOPZl1ddJWqAR
lXbS/xSe8DtQ3AkVqfSb76ut2R6kl+qcsLCFxNN+U8GNSlTXRkokI6V7EXbXVZW0
qAculdUiMGxcr8jqgGVKqL713H4yxO7omkDQN8g6vTmqx72ygbN5GUnGERq/l6kY
vFMLRW3YO+0acmAwQWBLGmtkfn8tYevJ05Ww21yHQfD/FSKocFDXp0AR0Hj/OFPu
i3CnP0CYfbNilLJPFqAS/1uETpEa7XcsAAa8uY+XzThsd4ase2nv9TillujOkGgT
/12OU+XVNVIwOUbE2+6zHv+kFqr8jQ6GIDm7OFJI7Sb79AQt9dKGnwY7IObeOeD9
dgFrZ4uJHlHfvcIG4HKBl3mrPH1SOKLbfVlj2yznhsyB3TngjgiUt3kljmfP8WmZ
zLn4TxqEmp0UhaHQRHiL0Tenk8WxPc62vRDHASRXeL9uALLrVbn3KVaFZBeip8Xo
JU1TFxrdnaT4WJ4VKetE/yexG8QB3l69jpxJXTd4cTqlVY4UfLOsH3FX3+p5LW2z
8Xn3msaAX2ICv2sue6PKnFFrCbk3IE2qWYPZUHiUOQE3BybxGOdhMVw/mHq57igP
+AYQSdb6kfyxw6jvwcN+/U0Zvn6nGspbXOzOONZ3E06Ao4UJjG6EmQhyqGYttj+r
pUIVVuysP6UCJG0ylIPwIrKRj9xO1hfXcrUwNdekBcEuhYgDz2WbO8Ly/sYPaf3w
27kHv2Kc0Rio0ZHj098S8Vfa7X3MJ4pZ8aUxHrYxBtQugrl/tiLhfwkvLAYtLeMd
brtWjITc5SuS3zqJFisynqwInCG9TjqkrxRojK3RstrD30wR8S0NNJY/FchwgAkb
9eSHmAMTxMZjZe4mkX3bSvaWazq8Q2IoZ6ycisS1jmHtgQ0zG3bXAXCusMByZZYh
L/6FXj2PcLwjKW8UpcM8MkTNv0KdqL3jGaxhxN0WLHn06tkvxDUxM7uv/g7qgwDX
+2DQVHOkrOKgM5OApmOTHhCJ87N28BmnqRuxAb83657ZcxyziiMffIJYGELa6z7x
3DShYYvoEcj25F5Xq/fihcZU1FUtYIDkJ8TLly/o7lImoRaTBtC/CaZl2+uijhfS
ocXKYvviLKw5afJzXzxbKKlg3ToKai65NLuEsZ4xGTkmFde3P5z8Ghh47Jdl60nO
54t1qa2Yieq/eFX0Djn1cEcs2aqzYjMWYu7VcYbtYahbr2DbgmVjH2xVwG7EEO9b
Ed/lcHepVqsXEl3z5USLRROJTQI1apdBrymfCdDnN6BcvBnaomIENPyZn35BoaDv
ule1WnDmh5bQBomsdlWJY6ATioNEOqcbGxYcoGgSe9lGWMzdrg1y1S2GvfNMH5Hq
n++NIPu+NZT929uY8nFGx9LZuBivmoL8c2QrSl4k5waKHo+hg8zz1AOmksjamIeL
9y1mbyUNbPK5j8QnKv1FieTelnMBgkPj/a28h+fHe32mQ3aHAmerGgfwCif7rQWi
88G5ReEUciM7rewQGKFfyZux6/YEGblfpAJDBfwf91zGSa835BJN9BZXZfsv4kOl
g3v7EEQ5dP1bTEWFf9Z1f05NlC4eXhL60P7kWuCz+LK0zcMLIc4S/LCujqHUiA3B
R0bOm/ExkXZSjpwPbY6btEfRIcKbGUhGjGzOMa1pDjobCaRfqH0zio8IUSdWWZW7
HcsYor9f9uTw9IW249vWWORy5UkrFjDNGB1TCJ+B3ubAMiUSoWZoBvFcFj5Pwx95
eTu5XTXroR/qCpRXOn5mRmdh1nw4o2spXDLXMgSQSZLZunprHSknBjiereHGlGf6
sgwlrVBw7gLhROgtw6OPxXqI3HfvKG7/60n//5MfTpHwHW7KQdogKKvoaT+a53JM
mwJj8+tBnliMytmwkRb/G8Kl9w1kt/laNZYwGt37Kg+BWMgRdyKbomQzp35IeXVG
W9uK4qnOS6f2oT4pBLynLoo1g/NLugWlOUxLbBK0dyHkR8NBglLs06eAtcEWwNIy
fiCPGmI5uw0Vdp2dhfgesFjE1HsLgrQ89Bxt9XptfOJrDexapBHeG3Ne3a969TtH
G1aZqSSqRZg2ILk+NMIZFPp4POzaD5SZosIV+G2I4G7y1EPpidSxT/uFdAvEfb18
rBbybrHfcdlzW324fkwIVEvXLl1uXTiHG56bywp39mmcrSbi6STm/kxXTzaKdvdA
YVKAr4NzEz+wyoInRclucXD66DrfTFei1IDBfDlCdz2yAov7r4dDVCsfBsYo2WP/
bP0gwnuD001O0bPb0F+DjrC3qAoF43lOd8G3CyLljA1J/l/wqTbIoDvyBINmPM2b
0NwpNjrxp3izIYa1dnkU93710tA4SZ4I3ORWaC+sbzFguSHVHCoOKJTG4nz7tefJ
Pd3SeeeeWFsOyTUEOMGrOp4ZHyq6reVwozk13sKD1Yy6uIEzsXkwPWY75ygz3GPx
p70NiwNK2w/itPHE1w3U9Gsae8ek19tbsNlz2AjoStLfuw0mHRZ4UTjI9y9XSNLS
8AIyLLl9l7thdYMfKHOmVQTV2Vp1n5mQZIrAke1U3eE6ct6gySQ8jXxqzuGCN2TX
nApVvbpmVMUeZeSWQ90S79IpOs4ukQ6HmDBR1Qn2jEmWewXqHwGwa2YFjtnZ8xEu
sBDPpMDlCWgR3uLfNSgFPX5KiaPzt+MTVO8+miPud4OfmRsFcNmrXhYfLFtUTI2s
nEru4COWbX4BXoQmgCk1u8o4EILYc2EbxGZH8fDc66s1y9bC/8XRKYqM2pomJafw
SYv9/FAyw854XneWmC+sP1hzNIig9ltOuymDG3rUl1S/BmJXFyhwUy046NxSVRUK
+RoyOP51sK1KH5QVWZJ8UqSTBLgBFFo2bWXAE/DFx9ee9VFOpI4JVQEHNTGyOxHm
Oj3SlaHRUEUF+KBvVbAhkHK3NYKZb/Nsy2G4sZbThkwq6NWBnKYVx0PT9+qpgx0l
A/+n3r+8sQvVIuBHem9q7pSqzUvSOqpxgEeUJUWeP3vgT4QzC+PGC//AW6+FrHeS
/sonZVIoD7uStOoDW4XWNSYW/pDdv/B5BCPoA8hg5Foq9vo3FcLq+KIcuRkMn8CL
XBDdBR7Y2QeUhBQb7rs0JptMJTwe/a6U7u5daTLDKi+6pTR5TqPnhB07XIeZNY7I
vn8nhu9UVL5Cu6xmsVrl9PajfXVdxtJOdpdVrcbqkwEwcsH+RnKaz5wKlcw/AfLr
waQMxOZVB5fXm32AJ54JO4Y9U12PzYNrIKPUNDrqpQfqPBmh23TvwIfe+F3Q8LIz
YT6zM9Jzjh2mUedAc4qxA9Ww/dopkl9Xgm5PZn/QwawBJlILXviQZ+Jk84JHaE6/
LXkSXmge0X3udcJc81nlLceylrx2iIINYq0vaaBiZkQSVYpq9VfhxFZx8zzHy7R1
DzHDOLC/5UbBjo16225/mBeApH1c6yygFBBPx5UQA7Zc40DYiyCzyQ15ltR02GjE
4an50Lce4ocvt+EwvUgv5rZ1wg8TLZWD6NSI86bXkSuS7A0CnKgcwKMw6Dhj3ua8
4M9DJQ7osh6phXAaia8O5XR7wmUGu/LzUoA4Au+lHfzNcjes8YLfwqAEzQ9ZpWhk
5fN2G126yWpqws4/H7aGiXNZDRQqZjhWbu+e2/94IKFEIRZXpK53Lmtyy9/QJJ0U
+fooI0NzfYhEU4C3HTYyTZDiWeeTf5UcM2p8mPHQpDvO/pJyrrCxlXnIdXz9DW6B
7rfwS83CDbRw0Jisql9o9+hkQBz1P2tx+yXQIuViR8uuMdVpIEXdolvX5TuTGRPb
nzylV4SoN0wkB29ptHHcWTkdu54gtunl8+O1XHxEsqKm7jeX+iqlorBZ9KOx6EQB
KKNQOu9d7YyQQswzhKV4/31Mp1pHYzu+/2EE26N8YFatq3NSOc3uQfuOfdzPLWKj
hMDzya2kiimoRCoxdeFV7Wkhkced01enM4q2WYki42g7wM6BEWsVObu87TOCuNj4
zX7CnMx2bhltfIMnLS5fZHLc1WdqRdiwemONU5UC1AYGZZsyIf3I0KyhXSBBgz0J
vPDYNbb+iaRvUnbyI/aKxRuDkyDFRIiVEvHVMlO9UiqAlzVL2o5SeOqdFd0H8aB8
Mw5ZsAyrgvv6C67tZRr1txu4VjdWyCf+rlB2m3CDdb6kkSUH273H7NPgtPN4tCa5
R2D3tmhHxfDS2WR1G6krpHzKwwxAwVbseBdfaXol55wba/nlN1YwRkToA0CNIsct
dRc14lScoPp7j5djetGHFCzM2axlrCYxnxDQrB6NkxKGagDcLobzbZ0g91/Z/c7n
jWVK18FTDTrrBVxeNllIR6hQbija8KnvQv7FvQj32aZE4k5HV3kRcNBwdiCz3bx0
aaRYp48ZVPJtsnB3lz/+/c+BDHj1nPHw9z0Ri7cNrm9i6LLfWsYPL1CK2QtlIGpl
YaWfoV+zoeoPeBZyVmXTpFHMjpr3+NjgN/17Hs/C3ClMOVBVgkaftkglOm+V/L2L
Y1PnsAOaHARuslgORjXmL3xbSu/0Fs/ryGPHK2ISVUqJh3ke+Q0o1lb/pH3eVvVt
yRCnHRzGyx7oY1MeDfjI++Nx+pLROb3bV74iOpg4t2+HPEUrK7P5ol+XQMNkqT09
6ozbzm5UL4+6c8B8/z+ilkhrnyrKlIj5OfPNpUbG0P14pHAtxpR7BmyjI5qCHTpy
i5K1GQCg7JbxIcMOOFVhOuosq7SDMu0S4dVsrzLH8BOyOxgGziEmQ46ptI69NXAq
ItfMuPWja+nHhyklRvO0Av1u0T5gZ+302ki36sj16bv+ydkBpeZiQaS/0cyy7CD8
4HPAs54I5ZtRyrgRMsOE1CmUOzTTkB7ijuar14bWcNxLZJKOKstmXMwaZG41Xfef
fo5MH399xkoGgTcwOrf+oEHuYM/JbAbVjX4hi8HRzAB7aNEdk5VFfRwG+si9smFZ
WsY+5IuP3PZ0Go9yQ51JOntouUq7P1/BTeodjMJrGxumogaRZYa2PfuIiNPAhVJs
DuKO2Ec1n/Mfiz9jCtbi4HG08xItCoaKdFRbVk2lBgMALTbc3vSd8by2bgUgOFIB
rKlzp2ru8ixGb37K0vkW8B/IepDdBtHs1WAEB8CC05QjLbmkSci4tMrl8lMT1qVE
Clb+cQnsNb6uYHsI8pMzPbzGSAI2pwZHpQrvHqbRwcBsZwc4Tw908TMyAqXQO3Ai
jklS8F5KN+ix9SMmB1vFJfOA7gST5NGRKh4O8BU7lW15uXoqbagL3L/cQCfj5UMc
jBFihgd4V7wYynR8GpfmSijx4PAKPyYvfbvsf/b01opMDakPjRiCRLlqwPEI3gND
xLWs8UKbl5Et0lh9UvpInjvkjqGkb9fxlgRQ/k1hmJPOYiJAAYjTjgXTLNAWDyKw
c/pFUf2lvzcZBvPuwIqeywf5qT7kdIThLI8pyA5D4VCnwaah1+vs1P4lKg489QaE
20HMoCywIhkyWqmFxF/xVcNmHGsU9GF9s6WYFgkYMPWjQAjk7SgxexdKMdAHcCku
IX1Cm2FbDh4JE+Wzf0/MHqQuxfAkNT7KeYXZ0OrDXOfpprYM8y2/HBXIGCOH+NE9
kJ61Zyzs9AmoaDNC+EJPDvJZBfGANgziZmV4qoP2TJ/kmDo+RwjYTDTDLbgaCeG9
qfl+KYeeNLMXHxzDHWxbP1w3rLvwusHpGYMo7nfQ+zeGVYyn9r3rDcUVGaOSBPaz
6vd7o/6uBaVsuNujT3tXqceKoR9G+2gnOBTuU7j8wPmuvf9d5xujviDufUhi+5Is
wBAnW0gMz+B7dZhkDkP1NRIYPb6mf1aeGSCOZN7naoKZVfrN6xdcOCkwbPhHSiGV
/TNttpqsXnsA8TR2q1ucSsvmtPW2upFRg4+9KKEJNzlTPiEfTwyJMyVL9lqYY7eT
Pl1ULe8oGzQ4VErytSdIiQZLNBY9v+iixgp1VZ2CSsFtw/v7XjL2nMCVFWpp+re+
x0i4pNlbK98gWTml6WsvrCcplvfCId9RERYPtO70enL6sPb/Gr1hrN7P5VwX4fnN
91fyDrCGVjHud+bLqc3rjGSAu+vfTJI1Yv7Z7ldZNx+rvzfkmN0qu0urO1Ekw7CE
K/EgBdwfIIPh0x1GoqgS5JJeBe7DUxILixeAbyH2LWoREPrXAzXSrWlioXSCDLZZ
2/4C3YmiFW4ASQ2oM8TAJWW2I9/d/pR9RpKP38FmvJDzJGe1GfuzkmUGfhBTU3j1
KeYJmrlXHvqthyddHtrPhu59OMcv8KVaD9zej4Mzz17WZFyg86uNht5Yv4jQ3sSz
HhjM0AyTE8Q+agKY7gs/mwDeFjJSS+/lLuYIQKadeq4jXOUzy+1t/Cx/fOSwdZtZ
bKfMcVWkEE5dCJPs2teTpAsM83mBzbP9IBe6YFtYaPKQahQ4XE160MncaWNhv070
6xM32KH1LMarl3434yxZvs7hRsAs7QhZeWziMtKfbeiHKAUpYudaHb9uJZ6+Ig8j
PH6l25v9OZa7RFbwNE0z+9LJV9VVuVpSLZGT5ZRJB1ySSLYX7qA42pjhJJU7P6iF
k0KgFWfsIiTOD83O6N610VGn/nbmYBsmVTysmMcDwWLE9Sea2zGruTEz8gj9neIS
YlpAsVdAhli2BIL9NjXTYDeLsQ6CB1nQmHsOr6HTCwfawFIr5Ripm4i2CAtMhk+s
BQCcbrvp0V6ZsivsCGx+6MANC7wmROhGt5PCaffzPUCZDA7sDjqVkPtqYgOXn5+C
RpHEckqEVNsG8V03RNwUfppm3n9awdLqmgnpHvv4PcN2fZSVSAn4Q+hoP6cxlnd7
FYHXKZPiyvqSBFhoBDlsRcjy51HTOOj+yQlJjgqcVmK3toucKFXF4BiKwgYNIH29
SH0V8VA6wevYcJ8FRBrGvGSbqZyxjDl7Z17oVNTlh7h29pBBD8Da6uE6YrMqthVi
RkffTlIB2mlYmwe5aU/sFVbjmGq2G7JUHbLoUlgF0GLJw8VlncztFqAXJpLDctWY
QpqDVNNNgDe5DT52XB7OLbwGcXb7E+XkqPUjS/ef/bxTSnZzoDHkeUOv12F89Dpe
UkRyU62gXO+50mZWtTYP9KaapbxgtG56hCG3uNbNdZe5Zio6Nx1/qzvU4GaMWCJK
ByF1YUUk/SiZiydc/8sPOMHAbr4oWNnHnWZKsw1euPP5PiXRy7TKQixGN+LoDYNN
Byo11ec+syNkmXLWJCFG4pAXJ0dA2U3lyo8n8gtuNLDX3/gW4KEdda6tFNJP3nxd
pULGpTV5BNmtPnyBYmC+RNTC6lGiPoNfwsCwTALROG/ZAgtHyenMzqDp5hIvJ/Os
0/1fp2Bb/QFOZI+I0+BPano8971fTTn0H5CPEOPEfHzHitimBt6S+J80jvusQwJl
8/Pe3AIlBSArDcY+zwLfjWP0BnalQN7FItDJoQdkHSuJYpMQWofSQ/RJ8XFrnZyC
5WjjOo11Mn7ZfzHLjUvl4co0NpjLAlp1gjA5V/aCbSNbMY6IzyibjqBeRhNish7u
K1vy3S15/igMJQqcZuwU91opODw4vZX6Oc/Y3VTH5mNrlxzDrJRmY2IWLk62EZAt
Iz+hSokRr1tzIuS4yP3EqL5S/8Y8liYXBqiLDpMT20Bis1h/XVkf0ksORkWLEMGj
zZTHvfJvnDp98j3YkGORMMdLgqbq798pb7g2ApVRS2zWavszGxbYXjYVjl4qSFEa
Mo9eKf+SCidtpFPBxorYuNaLXikVKKDzOoMpgJZ/T6Kb2B+3VddKvVuMILJ7MH7r
c2IU6cNsOUy8qwEejiON5YEbZiKJEU+X/VagGDCjt8MoLvqKIVVI6cSIuLBdwuAS
miUCWLbf8aurVgsjvpp0APFvruV6gntHs92SHqSdC64/u+BmzLwSlgzY54+UB0gy
80gW6aKcXXEp5xeNKoT+0Frh9CaRj36W794y7DGlTA7sNCOquXIeLhVaB/kxIHyZ
WJf7TKorVoAhWNP+ApHNwaU2fYIOZifVokKKQP5uzcp6aeVrJX5XLCIx/jDK3HkY
MhP4ZZx6zAp5SQ4U1pIyv+5CyeOiD5HYEXqJ+7+QVfNCIOtzl5e0jWbeqq0Hhixq
i70SlEpsxQfGcLmLFYIBAJfGsIefWvxjICwT8AQRv6x5LoSSlTy0oYAKedpf06cw
b6Eax2LGdSC6PYgiJZQZZ1lF+dAK/w0916B4tfqeK4q3D2RhMtsQdUt0x1/P9nqG
sg2qtXm8AUvuW0+Lctf3mPB5O2EKFps9KlD23BestM9xMdvr9sA5QIQnMXCWJvJ6
NiiR/CW2RRvBl/qirX3YEl21O1/CSeLZ3jQapJ45a3nzVACPaG+MHoWuEFJwy5n6
DJeYPbN8kgK6bTtC1iLrilidTv2W+yy+c3NPnD0ZUMjiwlZrLOrX315JriFzpXjs
BbVXSesz1M5KB1+3Ycbyp0hFQT2O2G2CZJfwJyl6th2aJKUX6O5pUaH3FDyYeDac
BIXcZCTdXLwSABk5HFJRpf5Ba/IAYPMb/vCeapaGs4+Ecel42imn/FtwhiVcwK9C
fjFgCcRcDeSvaurFd5RL6zSqfvtbx9G09hE1+HOZDkrIYPLJ7v5Z2FdyAFBhrRQd
qWtkLRqAMr7FlZCiYAQn7/OLkWc2emCaSL1bnfMqAO7hCEoD+EnyxM3EDLc6I7b4
1ZYRtS2ALZeB0L1WVBmixX7kALlWq58oQuudWmyNoeuBEgiNIOiAdX6XAgZPWpHo
hQX7c0mu6szlxAb+jgJtQ7xoa/+PcmGCpspCMSpbeJlHW9nJcvzArNXlSFjZL3hX
EUsrIHY+RN9I5XGtAN8uR0Gh12tNjeLaLCHqZKTuJ7oTZTeVO9Q8gpHPi/eiws3N
LtN4Ts/GQ3oTTxqtI3GHLJwmWWpvAdE8M3pitGboAyze35lwSWXNBBzH34+75m5g
07kmf8TOkBlIIDf9fkyHGpeAUJilqFb5ClMRxY/NzTNWNFLSWTvX4lwN/39u0kCc
y10nQoedfs+zXKdNx8BFZofL1dJu4ofV/VBumOSeGwzaJLDWFISkX2Rwn+e9GpJh
0DDWug3aCSQgwRcpI+rIEd/UZMrqlzlnMVdSald5oY5djK4EsMm35gZ69dtfNViR
8bmFBGtiQtsJ+nOn6+bB6Z+bi/oxwzFZmgTlZK8ycJuun5qGdJmctVMzEHRqKOxS
iB7YfddoiIB+88Bpx4gNGDnOXrK0KcxTvrtefYFE3lHfbe8oZsTx9zhLdVXF0nlO
DwhwyHF2HBqJ1568lwZwfdHEZwD+z/h2Hoz/LFul6C66GkumEDpOhyjIJPZSgkDG
PCxmjYcIf81EncSFqdEfiIMiAO75cCkvxRK7DUkuNhxRmLLRVbmwtsHza3t/RW17
yHtRYnf3b4BFQFDAbcyOKV5Ia5tzELxb6mRAjp4XiqTiMPtbOr2qDnlNoGlP5RWF
L1dS78R8Vs9Jzf4YBAk8B4gmOPnMaNyx0SJfj5mFNvHk0aYbhKbYM90GkkvpJ5Oh
cbDWzDxkY6iJvKQRMlQ3sFG29G8b3jdhxSQuPQJy4m4glXD5Y464FLW6BjdCh++D
b3/C0XlFrvF6LVtMMr6CH+0jY7XYu+wEcBIcM3XlNIqVfgvzgKDX0YP/aHckmrfQ
sm1slHKE4uVfI7gcxhw6OrqvUMiqRJ4ppKcSCdBi7OooLMBNFb6571d/KgOXQC9G
P5Y6CsQKmC++tDjBYfHFgwooN7QkQEmaajS6GhxHqLCK7G6Vuz/+zvGc9RnyYFL2
nosD+JFeo26xAW8JR1p9RnC10GDnCceZRSeIvRM04LaSk+EId7WjcKh65BwkzjkN
XG3D7geXOVNdLO6fjRqmFSc+reTIjxxJeIoKNGY7+bJLzMHeZyxs4Gv4179XLWz8
nyOyhDI2j8LwICGsWKTkG6jUz4i5ntrNXFAQt7WB6sKQNaeRVaSZBNRK2NA1bYCg
It8Pxj+I+oAwatofX4mmsYLGppC+SXY1MkxmSaxt1mfYklgo3SfMg2Qrb4k8Dyoh
mhD0Z6AKFEJdyfSxdqp2DUVPIYqwEz4qH+ngTjSkbcjx76+E8ZqZfJipjBQ36CVc
hJ73Qxk3qUHg0kh5+txboHvDIbJCKfqYtahIYHvvrnzGkHyvT087oUbFQWorr4eB
ZMmAsjd1Omw8+g6J+AQyt5QePLDxqJ25Vt+AkzFH5zs2y45p7Ih/Hba7LqzNIGIK
jZ4A7BELdseOhQ7sT0GP+sZXjy0DKutzV4OQz7iUU4pyxOOCdH8Sq2taZ4XDgaRH
uHh/2xZyJ2dTjJ+svoFzlQcJ7dwvGAd3/HyPLhtUSYvHs47JxhIFVVKvQ41YHuOL
/XdeGkWr90W9iPK2epSk+h0zQOpmpnFVVZsigf7u4ZSem55sgvHSPqBhmZnTwQ1N
L5rwdGkd3+0AdOuTlbAR0IML+pMoLFx4z0pairGPZIP0m1mbn/+9nbEHstQl77gP
VsuEpBs2GQuFy3uUsAAkqCKDb7bL3mJPBJfvtftC4OF4XX6s6l+KJFv44pwmemBi
BTlRrtfmo99l1/wOWbc1MXD07e8nhzTvAAItFxbXu4t/hY6tZJLPTtCEgQdIo+Vs
TEOLLRzrQqEnxycesqp+zVvoZT8aPdn3qZpGI9ayRMXjEWaPR4OYQvbmVm/LBNgI
48SoOYBrhLSgSpa8Iavu8ob6QRstKNx5ITOOp4i1UxB8ThQBv8Umv21Vf4NnMDue
UsXziBpCtJmm7OrxDgFHSClrlBW1NBbe4PUn+MMXfbUCOUowP8gmeHRZU/VbsAld
tEKaLUXD67vrzwnDtWofFHRj6sOccxlUSLqrjeTYBGyHzdHBJEaVk/SG3iRc4LWP
QHvfovBoF1ZzVZzZ/lceKDJJjF6lG4K9Opd3ihnG0jxWk0a8Lm4DZ53gTAPF6bVz
eKDqCmbF4TstL7G5Lt/cu5CW9JB8jXNGy5xrsGRoyxW+gxWIWhVQwszg5VWFVS9W
tdMsAxgwX555EELDn5lRjc1ZktGczIwAip/j/XJsaWugi2DJb8xx3Y1T7Hdhdya2
POOGLlsvEUl0KpkzujkqcHsX7SdnWasagGN5i2Qhxpk9a4FD8LQxQX26Omj8OWJD
TaIe/HcsFUPsA2ooZDX3lwZF1//dsX9vp9lI2S35XDKTBuREbfxzOIgmqrFQPh7e
Y/6zXxefefd2Ml274fKKNPvxb6roTpXd0Alic0vU0ArG3ifUbK+fNZvE+3LOXOsV
t2stUDotkZ//MisfHQhjGOaOA3O2xIMHtGErJddxlF93gAk3e+7ELaQHU2zS1KLm
FApD55iF2U1ov9nTF4b53Nzmjga9UJ0WwYUyhoRDmHFkcN0aeZ2Vnl2bFep/W+EK
hC2M3f6Lo/+3S0QdmhC6E9rKaJr9V4+fAXFVgTV3TIEcv/ELIehf07cnu1eg3M4T
J6/t2tGrI3JXao27IpCmKbKEODmcMZ/MNks7YbS7nvzl3aRG+FK4VbioBdYVWF60
rDwK42KH2XW0OsHYzYh1m3YroHolyyEfG4YJbM2PDuvUX7EFYcn0d38g0ryfaS9Q
mqY9FWWv6pF3dXeqHYVxmFyx91z/7JYflFmMCUJuGZruc/2c/0s3SUOMcwWnoE+T
KqpPHEyKY21vsQozvPEkkQU9pbee2fkBCyYmQDK/TILfdDuNBKN4kVzhWK0XVvvh
PpDj1nWP1fc1WDTv6XWZSBhyMJad0NzduLtdqlyD24dQz6tXj9kFttMRSzva2JiM
4qF8CQ8n0p7GD7YrdELMhUoSmXUQo9FCX0kH5/KGsM5BtSdR96JZUXI5V/n3ZbYy
re72wgPXv6hoZfpCgrqvQgiILVx49NVlRR0kHaeia8VTrNOcb7MquxsECsWfnl1c
PML6vKL7FWI6D8Z1Ho6ZIm2qvKWSnK5cl54jekRkYuEoHg/9xg62RQcOACRkB/9A
Zt8nalR/5jr5XIRWoozJDvC8BxGQlDsiFTsHKeGrLzi/V1Wl3j9MpuQbfnc7p0vX
OmvAmGBqzy2hcn9vdjDGhv1ck46LTG3/WIoEg8K7dZgXvOljfG8B/ea7wMp/ewcR
b5uUhlaM/xpvbLYEGHSWvSa2dcmWsORL/s0O50vAeNR4x/o5uHR4UWBL5y1VLMEr
pgwRq96drnt0wZ73r74AYFsRoZ6uWub68zRfz3zDjCx4+opz18Cf9rdyii9CWE44
OA7PDuV6A7brLnfrxn1zeOT5HjoASNgbqvggXzLGbH4SOG87t61yTcDU3hvG8NO3
qA4ZI2H35B4q9CucgrfQEPJbhGh8eUTN3D4J4bENmkP5HnMlz7LSqjJ8XtNWaLsb
0jh80yz6FdAwwIT9UYnHg4Y6JNXBioTPMXVkk2v2jeO+kgF1l2ZfkAD9yt+GZDbP
D0qljSjgIV76lJtGdmp5OeA3SZybHD7su/029+Ovl5lKih1OazyHTO+/wWqyTyTI
Dm+xEVaLD4oo4NIdIjOfK4URKaqP7hihTKA0Qe/IlBolCYEbiQrXKDvAIe2CQur8
hkgn/w5/x1aBA7jaSoEnoGpaGophjAtGt+YCjZSish7dxFJgZV/uqoZ5BpXPvCX1
GeXD5+OYOej47ghF1J659Q7TU/kLI85iTE25RV/DdmIvtTtNAL45Dndy/EZv63Uy
m9gqjZiGMjN5BY7s9g5XTOdOQJELpSIyWmYkeibtxFGBDSJhJyYfMkhIGqTDXL6b
CMsFYoULv2Jb/2N5oXStmUFDkqaT0/a1nEj1LTxYMSLFBhEdrJ6Ia76PZEWgGwSS
I6ZcRFUEdkRsH6fMxC0NNi1EVC8XfD++pPDAfUHFaPPgEYeajWhqiabMWsGFVaSA
1hwKWb+0wEAixBm5aOzTZRQaWj+0cBad79Hz6StTLFKxnJKkEC7qKgy4+6PHVlOk
8bCG11WFP2t7RKCmCtZen0VM4V65J222447+gpV+PXg6zxeuKZ8V9RrU6GGe83qe
0gLi5neIMHxjl5/LjcSchmCMOVXYuSEHPYFrjPPmxv7+Le+MOaUttNXe/cKAqL9k
wgl9jq5x2Ccp4r/N2XUIIqL8jCA7BiNnNzDb4yxu07dD6RzE5QXqbQMA4D/m0a9X
0zUIScY1Tw9snxDiVGN6GfssoAsCRBY6X89IwSl8GKE3VdERaMXdIRziMghyKaO7
y7FCZ1bJDBslk2DCtM26N+d/JIxXyzu9Dk5Ma2Or9v4igoXnJf5rM79rPreuLfPn
xxfYYR8RQ8vudMPN799fkDKhIBFnkqSWt3Tdh9U8BC4DjVN7n8bBicbM5FGiBKD0
gBRGJYeIxLPP8VArbnm0K+Atc3BVQGv/vRs4HEvCKZl1cTVOjKV023CCiCqRCih0
/VP5FxG2mPzjgta9ghgOlhzkMhQVgSORHjRb5fP2Z0t7hOip1e+eOup9T2C0XK/d
j48khYkiGt7+4Eyo8p8kcnJsSX409oMbmnYo8Xtmx/PcXIpfvpoGPT5PEQu5J+T9
0feu/lvBBpq0vdNiKMHM20qZISA7lOrDWqgLF0Bzh0BLdJ/p0/+NW4u8ZcMvJEYH
0LR4EV3XSf0OPHWAkwdqjfrgUuf0f0Ad3wqF8O/5kwdpnYfjh/H+xVrkokgt4GvF
Ae/cHrxSohUMz6JWlLzbx7vVrEGIxhnX0p/dsNvtKtXe5dDcaPhPWsvHMcUoN/+n
MTW4Tn1BpexfXnsVXBv9J8xG3Sz0GsDHGvLUPemXWbdyqMOEOI0Iehv7+dH4K86i
Bv3i7uE/eOCpY2ODbbvc2B8H7dYONMtK8gTTeE1uEJXQvojPLy7D1asWbYR2O0PI
MqBWB9lCJdby3Q66MoclKFE6hmvluu71GQDCzdolEltMQnmQhRU1diQLrvcVi4dh
nSHg9qS1sPe5SBOCHG8uI1fW8r0b4Gomg8/MujzwnQc+dEMXA9738sAM3rOHJLo4
Rq2dvgCt4WTTd8Gg3brx5Zkxzfs4ZTpk6LPLSPRYijPgbpVwTMdy7RxxmA5gtEJP
FBAVuvlykpfPS/c5iBkn+ksX6qAu35EW3BBD9SprcA+w7ats8dj3MsTtOG+kyzXP
RkyrUMdJ0ZvGp9CDDPRSobw26ChUsz1a9hczDiwtNeN2MWIg4sVMsMiXAwMIt3oT
MFBbAGqaYy9nDgffqT0o5glribf3kNbzRkGSGzalAYKDJ67TF63bqQaN9Pfz5QR0
ODLN+FSJawmrw+Ie+OLeNkkOLqlaLEua/S0uvSIe3is+a4VBVPiCku6Z+3gJBDqh
uftAR0GI8ueOUYOYLKzk7rDXPf0WjbaQrBxPRxyC63MqncdZzfFkgpvwY7DGur4+
xoR6YW9ynAQohTmrHQrUmmRFg6U4NzkfPI5Sm5+hRO0n98e9bP+M3NZYZAgTsw6K
GmiVXvL/3CpbLgPaYeuLEQ6EeszAgdRm9FNrwTWIcwxsRdkEIFDtCAoG+mAu19e4
gk4Zi1nG069jWQwuHAfOoScyqhkc9xc7NTVIpMd9tdXKcRgmCN0S5RLx/djbvOiF
Bf7xlCJcCX9QX+Fxb5Z4yVcKzriEabw3vgO2scJ+KzjTcm3LxcIU7av5WvMfBSvW
koYHCEkXOplyvOkU5hOkshHbkvUBfkW0WyRt0LFT5gxumIt5B+VFZKSSwG7dMf2A
ppN/FJUheQOj+PyINrJu3uXk7nahPiW6nge5bwrm/Kn7JkfmCAv4f1CQ8p8aAi5f
f7KzNMPee5Vc5M22oTxy5CPbl4iDzEBL0GTf1sE0FdkvAcsnqN+Bp0/ODyxgLkwt
r0Eb9m5GrmtyBpX6lWHnTQJ2LC2rZCPJ9jXc61K2HNdr031pTruqU+sHCefRrAVB
4Kap6OvqdFv8BrLKZuhyKXcE208lLuLHk2cDORaWJIAS9cJEWHpn/y7egUd0N2TF
hvlYhluR5DwRbyHyMEzDqZgZ+udWEsqxTBH8ogbeAdPfI86/1YD2kNIjQvMAXk+k
cF2O2JKD5im+VCvbbog92/SzrUfcbv3vkLHSFOHRpvrF4aXaI9gEQbDd0LtaWd3p
c9tZUbHRdAZV0mI3X+CoOPQS/oAKTAfJ81qYBDXNa0YF4H2Mb4fuyIuTeb/qnsrG
pSWBj2C6wwrJNRnjodJvmRl64+wcOC3Z9JDDcyZITPZWLpVKNgf/z+3UoQ8I3Qly
jcuBvu7TOv3Wqf8axQoNkoJJ+/VCKRpLA96b4Ht9F1l85gLf9/al67xPHRUneZew
nyKRa3/NTSr/OBN/Y0AyxWEojl2/9zDD7350uIaCqxyMN643ECmeWkHsMwKJ8ar9
lxXznvlmYsObwnVltX9GqrC/bO3vE/bVyCawz1GKlrd+cXGRzlh57CdzCFIaDNdS
cRmzR6DyTkdmTPeycmq1fUUzMvSt9hNX6fUFx80YtlQAsS/W4TGXx7xcSU1zU+7p
tJp5+DtK8iF4L93sitEROcRMXFwTKFM+qZ8lbb4eTS0woLzZvr+Q7eAEQA8l6JeQ
cMLxzilTXHGN6L3chPn+EPNQ+juldSjlT+Lu4RkPu2FxqQciQZ3ClNlwPtXxrLf/
csIVJt66Si2D2Q+nbi8E9qoPIUC31j0go+ojLuuCkaia7Y/b5xeT1+jlFQtWnv6K
yXIymGWk1cjqtife9YsrvHgMtAwNzOFZqiPQPcvT47vd3dLdeU4WFVfYF/ga12lE
Xn/8vLAqFogZqMASDQvrMSG2sxlcnecOCX6MOr2R0XwDt/JMNds6UJfcIwDAKZk9
Z0dz1JPFDhENcjjsHJT7X8SssMTRg29IJ9ZvnL0pb43a4x+4n5vwOG1IMvPVM6SR
65nyeJ33KQEJCW8i0sK4ChG79baNplJmtlDqpibGL0tdS2UheYv4qAHZNs/FqOXS
vgDNynkeeX6vKxcpseeAqxot9r0j0y8G8mTJcBo5fheUU6AUtvFgCatQ/li7Yoie
x4Af4GKowH+8yaVorxNRsz4r2lb8uJfQB3N1OPqBNWey3Nt5AvZvRfUE/s+BT/oo
g6aURZVxKgm6WDR7cq61JeMFtD9rY0I+B3WWKh5R2WLAx0/MD2DfA7aWiHeEEq5x
TBac/vfc3i/UDDWGM1RJdbTV2ni6qG7jqWlGpiNzOQpc7PI5O0gui0DNCWlLr1IP
MRxffiCnoYOBp4EdqSiEWxYWTPWOCU45FwStz/KbO3KIlcu/cHuicuPpQBTXCKps
lw77GRz5ZsKflPQ+jpiVoh3uNebT4Ee4qdRkkVU762tpiVlOtiGksyc7DvIfVlor
9mu1yjAc49z6nlqrdNxhFBifjXapx48GuYWExmhd2swnkb8K1weKPh1C0bCj3BZS
MsdPFxlb+CGEGhV9SSvQyXIqaYVX96tUol855sjKhmxKs7ApzGqQTIAGUhjPZN1V
lHJLEcGFmMnNQRd4OwdedpzUxFuod0azspWnlZhxofbjJbdr0EB7nw6aCT/fFZei
HpTbE8u3sgI95zN3zVJ5qzaiseL5hYkIYt8gr821oRoNFzcv5TI6Hd/RolWR11Os
MegUSs15IikXqXY+EjnLJxQefHR7kfN4N4reGVLzqW2C2+R40QPQ6QMzS0xxbfZF
9USqqbngmD6TfMVb+2WkWtB+SiJcBVohCcsB+sQ8dDRAVbhqtjmKjPq6XcPGBh+r
ND7nVbRlenoLUOHBlgXoxZsWbV5lk+FTnZhMt79cutRfMVw6hdW8TNExqxRWepfi
MutJ6Yujx+Lr9ZqIfMkoWPAsp4TIdNTBm36FQawwFacchgTsl5oLun+A9Vo59jke
hUCU4fN4LOLMAhQI57J52NmR/lYXXd37bhESQBi0Mr9h4x0y+l3hDECj+vnr4DiE
BN4yT1b8/3uUTcjCQh4C+cAMLKOtRkJbva1k/Gf3ell8ZHpahu3A5ZwhIf0PvIua
J0OQvnoDoH5RuwF3gg31eGvFdTZYfPCWUJ6xr0w2FLWwATIvJFK/N/rW5NklPKM7
PLTOLeqQkJ91x8dlxvPiKVgEbxGZZJxLpfZJRqwf367yT9M1ZrAptPI5fTgl5kcY
wqjbV488BN6iLKf7MHshevjz4eNAyvfxuE4eLKoEck6FxSBgHrESh77za7NInlXT
iupa+aarkmh3Dvgmx71VI/8FndsDRTxm8oLikQ9mlhP/ydl3VvggWy6gNPNyjm7P
rRZ27nfz7rpLmYk8/Hx7PpPHh2VkGFbt74skaiiIc9MpS49KhWoxUqZnqlqyVmP+
WjfoQzced1Ti2LjwoonpQPZGH0dScYWH8D62BzHer2tA+qpRUHxLvUwXrD4QHhhe
FRR7BfwT4NbtMSsewzHFHvnX63qEJrL3RW+N+zrt/RJlO+QcP8jgDjvoFg7hHDJd
eo4sR3wj4KrEbal4UptQi8M9S6jLfvB+5U1pRJR+tuIPpRJJ4IDiI6OL4gI8O31D
4O0PRAbODfpe/CMC0rI9wZzqb0jEvVdmBtNqC2W566UulCRWrLyqaQI40lhsLNbj
VmpQCQA6CxPA9gkOAfotIgwGRzTGruNY3BFuL/FE/HU5RVYOEs0uQIqsyZWlojGv
fuBFmWSOPi/1ezZ1PvRK5EokxT8Uk7VaDRVQaPqyVeEHTyVUelwNYKYXxNn+JIOU
2G9qus0adKGOZzPfeWC+S12JYroBJTDHIoaUlITpHwCqtvZsuwElSCaMpuImFjb1
+emsLu41us/161sh6vtNXOiSE95R5K+49bO2kGva5sGju7wYgda7PCeSlgFHrve2
3zD90vGiwjo3G2tH1Zchfszx8WeLMKCvn4EpzOvXeDmOxeF+1CPWefX7xSWIcyCL
NHKozthbxkOE2TUwScV5hnlnRvYm8L4QyM6WoyNyuFagvy3JNhyzSTjDWNc3wWup
yZYGRe76Q3LFjrWDG9tRR9md19KftlCJMfFfzkR+TWiYKHZ89McahMn2NMU2A434
poZhPOIBa+cthmFN5AC2cklcquN9K5M4ECxZlLANdZ9pLjVp106QU+snQW0hphj8
YFkmCkxPNfonT3J2ku+zJdPi1TXouVuwswxSDmLdcE3/xcRSI1RElEo+zSqryAvT
6KoRb9pQGbAzU1wLsAC254jOSz0lqaYRBvkAF/Kcyag7bsEsXWe1t2AcPgRXD5VF
j6f55lvQ5XRZk8svuYo013HjBs3f6FHQCHiL2InTvaz6vrB+pmgFpdYbIVhsCzad
RE2yJwyUQBJOAhLoNf29FWfS0dYYm1f7dRxdJI04EQAQ5761ZpQYcOGL4FIanHG0
XLae9u499N4ipdLOLHTtkaU37qgp1g4aW0xBZ8wbjN9hNOO5WSsIJadpp7/ShXss
pzb2CSvZWvAVwdZJ+sHKs0Ac7CYvj6JJnq9WVqL/4/3NRYjWNoE9lG0cbvGh6eGv
oTmGZ+Le8hlYx6UUv6DFOROMONBvj9PG/gueqXo38CV/jo8JQB+jRTzFycA9iqs9
+CitptNamsFGBl9JMidFnot7Q4YhAPHKNbGcrUoE2qAzhRUiAL5IeSWkopSETeKZ
iQEmryOmnMmFowuAdMORxjWmkJiRib03KGYnXno8e8BaYI1HE0SSTMHKJxhX9LmQ
lPqRr69ongc1JaQCpVjVXZOGew0i4saA//TEvpNAQJ6ibpYDi7EKaL6jB7sBR45I
ZGHs/KoC0BJTvjPxal+HQikHwCA3c45Dgm7NsUZfSPkY6AQhDAcSBHCY9XPKJD7Q
ksLct6I/yIytPafbhT3EeD344AJBQRIxrtsoBOn8x/6hd6o0KXp3maxZjHDBxHzN
xBrIv9nn4yDR0ZgKe1+vpQPLfcBgWMRlPmwCy8eFLbYYDBivm7J/VuguVS06U8RQ
fqd2+BKxqdvEc27GSGPgL7fuL0PfQFqOMrTJzzRrztxrkOkQGlGgUko5nJJKJh2r
ZA5iwF3pptS6V6Fp2GVcjkhmodUsLaudZtnU2hkFqpcZbtH+UM4Dyb3bLd8hYasv
Zi7DKbpPG90820ndD43bo77L2VFCxzORJp7PdBSVz0wWxHiOiztzVh2Kiz2sX0CY
+BxGn7UcOoTDr+5V9kBmoDkC/byKzAWqqIyiLVNz7VnmyCokJ49hBzAdstaoM4KY
9I4yJbmJQsFOa1LBYCqqhbolwWwYYmtJVGBas623XAMF4YoDuuVvsriXNlm9i1Go
LIg7LtcCdPhHEfup8ub+Roi/6uwlZpKLyavBh7vd6kLb2a/+3mRr/s+AOqyGzZJf
ZwR1hHDT+wx72BbLuKgYN36WSaqn/j7tvtSLha8czCWFO4oD2L35o0NiZakZy1Ew
BEvPCDpoROHc1o2m1+EUGcjlUI7kmixaEWGodo7sTIll8GBXTJNpO+Qx1jpEn03b
7CtBgSeV+n2rgzdYXxe1WH97XPWVR0zcdLGLs/B54pdlHcMbri4pkPTC02zeGahM
B/hshOLIRxuLZtTuZTanbac7Ip7qJKJOCq/dcpDO6xPP4PVaDgCRCe+fncm0c1SS
MLJOCQVI0GfzUSZBBH8wHSADJPXQtM3UU6001ja6+J92uRGJSJfI5LII5X1lTaGX
BKdxagBk6XQ/k7CSj33Z6Cf1hyLRAY/ebDo56p254Qj3TeM8cenLqvbqMfcP1XK2
iEPz5XpH0796ZaGYnGNd5q3snA2AjEc47GxrYJ6rRftBOPBrzuk8zU3E5NaI883b
ylX166agbQ0uDUtDbzcql9nRodXLMhFLYaai5W9x/7q3unSYH3BaRNE/REVnt9vh
aO0nN0b3ibcYkFJ2AasTOt4vGD1Ud+m8G4NEWVgNhIMCEAUyncPSaQeMT17Uz4xj
zYdX4VJK1f7/wUIZejWPSswXkFF/g+9b5mwxE7mqUYEDOE4m1ebjcdRCS7Tdh9p5
cGRYerk/6BKgE+LPLTZMGReOggdZ3nmjbTU8rLckdyhtnIegOUrlGZtdT18kXpBi
/dysUNTWolpqVLGkyrlP8cUTRNBh7MWDBPJ71ffBgSlH/bdVCngLb+n/YR+ScSeK
9WJ5N9Xm8czMVyNTt44QXXljXsPRuQXeAZAs9HZaXNGbcNAzlwTTuzd+cyKerUcM
Do4ZRgk2dKvnpOXC42cprldA60vFI8UqVNrbAvn3ipQx/R1UVw3atmCLllx7hBPG
idFWJkcwrMrafG8vLysZ49mVO41nVgTmPQbTCTRXqF9OULQexn8S02ylmKAXuIIn
v6Gfs0v8By0wiS+K3MF+uhaD29omIzmxvAPVGKfyUh1MLOArx0s00YULcomAu9o0
ZxthVgzqQqjiMlrfi7da4T0EIu7qLsfpLGHLemmOBdMpEVGlx8Vgc4wH7TnUoKjl
DOZaSRfFKTa2EEk12aL7iVmNaN77hWBVZyPN3t85Mk+LKBi92++E4sZxFXHKzWm6
c038N2wcSjLihDXW99GKdBfUaCzvagRmPpv/YGh6wJtdGgTnp1NiwTZBaY0mORBO
AAMsoSykaroUa1d/zr4wTvKg9Gpu8MBRo+0+KJ7K7+W46q0LXiCE7+nh4TKCY3+M
70HDj22pD6xH3bWQV8FZCyV554DWMkZW38UMDGjSztWI+Ueg+8FmPZaZkX/Qp8SZ
rKiD65uH8OKUaeUb4ye04Ar7tudogkPiYLO/nW9yYzRM6HdJCP1YfnXUA2wJOXXM
UN6T/jFA0MwjnzBqfJRDo+d/pIoY3yEL05B5vdLDIqiY+1ZKssAk0suqka4c9vfX
8EFJZYIM6S9uGJf/y1oJkNxv92hCLUGH+47oX5WL+zOpg6PujO7Ldsjy6JlvvVZ0
yvvARjTvWrIomc4Jmrutqd8fLOuS60oQzfKN1T3tgaSctsbFlXqGA9CsC9H7qk01
Fy/0Dj/gVI130KcaiwmoympNxUIPKIbzqHPKcoySXx8Z57Voyb9C6cJWa30pU7VD
cFOqxxgUi39C8TInhCxFeBKexJXcB9V/REdWppPSZMqxXd5/vv+SaAZSCtcMN7Vd
1vqdfS5+QN8BxHA/JZr9GjPCXvkkx7ForPGTje2tHAIyxeKQAcbPQsxc1vArYi5y
EVxuPrZZjDJjnecFqUbJGJggD9dBBXkNqpsQGzg4JmDeH4ZeFo33f8N7GJC9XTiJ
FGCHizvQAg2S/FNItco4JBsS9w9d3WHrwYR648Ky2SyhxGYQgVil5cPj/lkb3DjR
NiQqHj/xl57jljP8DBY1cR2Wypb6JLKKykJxP9AOyBHFlZP+sG74/VDkEJsFV8UV
imKWrq/DoI4AIDOnhli9xb50gfXpglBjF+G9r05wyihyn7EDtHCDa4nKUKxnte6C
bbMDcGu28qsNbH23CaNMFBGmx6+izU1qch+5CVKRHunki/lRF5X9xjSxNahW3Rjb
XDAyiFMtPMRPMOOZYnZYtZ6jJKOfsiJywq7OL82Lr48RulPHfcATWlY1+v3jz5P7
7rj/J4B5kd1karRInmSSqlWx4WlzRG6VA356EKCqf32HBYnCoWQE8xHeqrKwn699
bBz+HxoRqmRBPzVCeAuUNukHnz02nIMbJQu5Z2L2CI4zivXz1JBff1NaLmo/DTln
gAh9cTRD6QZatbippcDHebOzcwV427QaRGV6mM3RFM8z8HQVE/yRf/CT/DqN49+U
rWy3o5+QqAOkj29u5vcFymCj5GwojeA2Su2+SQGvnsQvsJkmcmAUiwYxWkmABSdt
AOYh7F0B4ZL5ZEjNqWeUe2dUYzYjzVy97qBroQFXkWdZz2enaHxrqxUyHlS0Ocrw
NRE6GB8I78Q3Uq0DIdYfuwdfmx1avqbH3AQnz8/W1T7XpPkoK01y2lDkz5to3brc
phrDgSoxqsMnosy9S2aX2WfJ1nS5x+AYsN4M356Tl1OU/iaHteyIIOOeXuG01lZE
hPUmGFE6soOS0Xo6G5usv6481/3k4S5whClXoBtvKgjuX77oifIZSNiHjzTpQwSk
r0aa1kd1HUSJwI/56jNVPaSM9Y/dorK2V2xIydGoHgK4MljT/22pyAP2Xcoc82ce
IZlVsLWCDVNPniVrPqJtG1lKkKoysBmhe4wbAtEMhPxzNlqTyuHPUbq09K2LUvj/
lbzPFBdyCVYn3sG0Ku14z97gQl6jCmvU4Yx+7yMMSIBkWDsw3GdbWOjWC8f05agb
mW/Wguo61+zIQq9NlvK8ITzmxsDd9pUIBHgCE3GfoA4iq+ycvaE+ZtziI6oxuORP
vhMUT25xGDs0LkXYqBJngYj1sn0JQvpw6P5KtiD5B1+oRfjlFEPtH4jMCRqrq7m6
+2fKcr4m9YK1vVKqGp/1G26iEtskUwulRAEJF6TdkHm/WOC4IRu+z7rqLzHyfxZ2
fnB3ZIP/g7zlTbx4HpRNfXGWs0pXYd562nNUYx4AO6DWtLT5jwBdPDJdrwG4sHKA
1ViX/bGZqdb1EnqUtvBHyEqbjFzve/gBufQjIy1rURpl5m/SSl3yNiEZ/MVWISpJ
SHONWg8EN+K/h/0HAEH2rLSDQFiGJmatscgVvbUIJNUwUtBObnivngA0FnZoJpGE
tdEoMuaCAsX9DkSIVGnkRvlTpMDm39VE5EZBbnPxheFfFQOGkfUDZGqsoe4XXM/y
5aTeoZa0X2poU1Lck4lnM51n/MXzsW1ceJvU4AY6Or3fKU44fybKEZLli2df++f5
4tzhUz2ZvaYLbnm5Z5RyqKxxF9t+TOZQJoPDHF7lQpla39k4AtjjL7YdlqSfWvF3
mTmM0qAioO2xGsJguDtEMI3IYSVJxZ0JlZq2ABtrvZz9VLDn+dNmFskAQCgGofjL
JdP3p1Art+O1zZinI0aacz5bFkyttzCbSV1JFXFodUYNNAEyfJgJwWkQB9cFo4Qo
asMfkvqqg1vgVRfVrKCSlWJDZQ0SBml7e14cqI6OcmXCYJ54Q0i7FKvC04PfnbZV
dzZ10s8fm0bzxusgrduCDhh4XFulKBL8IIyqUlIsGsAVAxTuv5Emc91f74CTVlnw
vcp1FiVB1t7L86RQcGp9mFsh+p6Aen9jmV7zGrnbRghKd4puHrzlVdFEi6Q++gi1
55H3VvD5ojU8PqTP2MUyXzok3m5kctqdTETJ8z3acNpkO7LUUDTA3FykYa0CZ5xX
b07ioWZWXZVi4iHUXJ5VeAz6SVIOx/eaKyXXYPeJvmvOi5jxzblMsbxK9yzdENjz
bBgKn5qkvXB2sED/70soCdxcBgNrVMpHUDfbstYBucUTZmhaciG/rbTUSM+ICXr8
gWu7v61YbZSy14TaZt/NNpxflfxduz4W+m61AP4GrwDLvNvFazSNx8g2BFrhaJo9
hVY7vUi7622516uhIb4Z51Td+BgN+t7CqtEy8kMCUwcfvhSnJM/99ZRIng2kN1y/
djiTT+jPvqW0iXcDPZZb/dDH2wGB8TVV8zvMGcv9RQ01o6AP0Pwc8zQcEF00kgoL
bryTHUCcPvEyo0iYApXB6kA1VO8rHQ2SzDKxL1IKHisPQq2UJ5WPIrc4H6J+Ks4c
EQmR3O0tJVop8hE/uUhZRj3o+R/Kfd0V+AAP+0PXLTnWfJczRBy13dXIhRSYlEfc
YZ/wl015jj3iDZ2Wep9yD8Wmw4C6PTPiH1N7MwZTo9/+9GKFm1WtBR5XwK8QF4Q6
ehm11taAYuM55Azuj54vxFW8QvXWs73H3BWc3waDne3CDMP1AAopfBW+6B4EOFfI
dwok0agtMgTXG2DuXpPgC2YzSvEpn95g1a25p3vsd5vRB3bGKSotCe+P7+YcO8XZ
A2UkdW2nql5SUGn5GPMD8W7anSM9HqLYXCipuPrZtjubP5jmaoiCXKBrn/AA+8i8
lkDrj2MF3QkYbi/eWml+3KEhaiVei0VlAfMQLgSxAmZyB7YVTUPiB6st/9ETfxyt
ExksA4c91VzkUTgCQe6/eRJNAgjnb4g2Ppa/Tguvw7w8eIbkYamOtVzoLELKhdfd
qT/vJO+YjqIKV+b3dosWI5ZeT5jJV7uyAKbW/wloosaiQ/b92tIQ9amoqsUMsFkt
SMb56J112Rk/eDn6sxcl80ajRVQ8EowByDOOwrvGtPviEj/jr7Ucta+VS0TFWuD5
vTFKC15yWTHqUTwRhgkmYXufyeot6H+RQwx+m62rGXGvJwEfEu+2xsboW3kR7wpV
AFrVP9UpoGMoiXeTQvORMZbaxde5Un8ljF9bD+jac7AonJdnDy3DDpqhlEfcvaUG
ggKUNScdUo9z9004AQChl31qfNV6J9iJikZJ9bRFPi7POFXND6RaAB8R6Wbs32Kz
IRFAkT2bFOjFQc3+sj1t6FlAbVpGiJgPPVZ8svTcuoh1r/uYynckAxi1N9cw66yI
xnSmc65rZGgl56tJUn8GbZTVs2+h64+Dtz8C6I3u1RZ8H+/UuSTxti+f8738Aryf
71o/Hq2B3P59RpaIPqZ0njeOh8j2L0JsduK2s4AI2EDkPY6CD01E9FNVRKQrqvCx
F01EUTGjkyK3bEtfmizTROPM3TJ4Jawy7fltEr4H2W5ByRDlnl3AK69jeCBcSDf9
IKEol4aGFvw0Tyri8KI2Wwu3/BaFQRAotsJzzhjoBixGDMNbHWv0D7/aKQCMR2Gb
PwJlJ46GrQYbCxG8WaaeVmQvwU3GOb+HdckUs8YyE9t5sZSmbCWzGSsz/pyOnKhd
s5rc4O9sTSz9EbhAH2WOapFhOCYirSlogQaUDslmZu3uIJb0KWT6gjW6x3Aa9Rmm
MK4WcB5mJK3GWqvVw/n3qi0EUNnAT/z78mknBciapJA9lSTrRrNhIfUzN7d7lshB
q9dcXqo50ydNdbY2FjKQknE6rodDVwAY0liWE1zo0D2JHwlI1Hd6OTsa1JPr27oe
xo7WipPJ/oF4zu4XlPBPFzeIGvJzoPP/0y5Va2rSw9JUBRZ4rzh7qNsGl04AAOTC
dSsAB4M+anYuy2xDLlp0va2hgbmSc3EVEP0tP+wz+FXL0ZDvBew8jEVWfTW2QqYV
tP1+QfT7DfM6Vy+flUng/X3O5LJ99qgeUlt9kFPflvM/YPrgMRbV51i0jS4zTaTD
gnHDjZpq5DvOPWlXpyqa98q7KX3Mxu/fRXTZ4An2icK2G/PhCoexXI9fH4Wn29Uv
F8jtapWQW38g/wWxm3iyQeX+Mmkblv3fZ797Lga2eoEBh0+hJHBafxDvcV2SiMJY
Ro/H7pYPH9yAtohP96B8kStWbU2ODla5HSkpeD6kZbkCFrkhaxTtylSVJfMHKXnp
KdStQWPLe4gL4nbsMCDZnhTUBo+tiecpIPkBxqntZK+7NhUleduz5qvhDT52dXPp
t54JWM9kZnSV5vGECJ5r+OtlhYPGU8cIlGeYyDyo2rEC1xBfAvngtv2r0Pf4l60L
CtGeRD0VqPhuPHP0tdQLXkbTk8SklwFDF6kq4MBfe0XijPcScXhAuB+iV/qfmusN
nOTl7iLibi+RuOZXRKYxhh4No2KhPBEXA+WujxaICVo2MjLBpX1nhfsZOZ+AGI5U
h98TRUH4M6ki0iSKL9NJuZSlx2M+G665/5dox019eonuzAnaxJheu4ZBrP8fZbM/
KtiakJlotfvuutcj0NINWjOdXUlwDla9EKh+lSgEYogXbhbEH1s5yVQ2n3FoAoob
+nlHnbPiKXL5aKFDfi1tputdipaPzAB7TfmI6kSUssTlwSutF7c56+62/Th9DH09
kMwZROQRHyMpVSssLcJWQsteOD04XNzaeZFR/Nkfw9z9at0CamnwXAnxk542syJT
I4mn5DMwRBwvAoP9+pIHQ8oXujEgKiBWmjVXYHpoxI6NgekqBfNdW4vvmMoZuRiF
fGwl1wUb/YJHaKCeE+lahp1nlaQ0P/obX/TWjcZLecOiSrlAFHpJ2FYtZlF0qh2Q
LXTGHyqi7eDssYYY8yVyUX9PTwVFE+SRRhOetPqbaaNyqntPuv6DCjU5GC/XXM5F
SByMGF+fgERoplD+kIFvt9CGqdCQmRBG0sxxYpETnmCvdB2qvBMIRh+xha6jF8jA
J2L/J3iqVhZBBnHZQQ3Om5hH6AVpKAhlkbMUp6LLGNXGPkp06YQXKfx8n2Xr77n2
LsNt2meCPTvEgEoQhvaRNNE86WiTydVG10IeEDp0mRfO0bnvPGUoPSIj1Y5B2rXT
CcjDT56DTIunNWmmrHqdZN5ppELleY02MudLU0WBIS1qfSfB5k8XKKxDCwndBbRE
1N9aYQn1+QqdQSKcTMik62ys9XSIE39uBvM6Lyc+16TMhTRe6+eDZ3Sh/jUc6mbt
jqLYF2bHM87i/Apulo4yV7YrulqJMe1FaowHBlaJwr5kR8s/e/JSXE1HWnyOaH0X
PlCHuLXSI47qgrWNFjPe7qGO8j9YzOUqHjnsZAcwKCldk3QhNPVIB5clsii1XBRn
Y5ic1Uj7aR8eb2o+SsvE0Kiu2bmpzQl34SGA7eBknxs5uWQt4vA/6h+klcCWxrFZ
39ezuQN0YcI/V7a9OLIVr/JhK4qQ4qnZotsQlrUG5I1ouzf3vIwKk7Ii6JRfqJoq
JQLAikpDs3eNXvIVq4oPrKC8iVATQhztVf8bokUU8KqoNeHrQj14IXdgHYuTdyWe
XFXF0WjeBZgjtOm9yfSb+PyqXR9nWo5+HCuWRT0usUE/U3R7Zk0I6TVblgRLuOnv
QITmX4miNezAA+EbhK3jd1vWtSBtd833D2+HRveOUDfJAgA4I7GvSoHDBYgp9GfE
P3Aw5wNezq2+2FAW+8rhKXdiWF+nJUYXr6eLnwlV3Sm6a8B6ZDU2OEZTPBLB8mKC
kLPWpc9Cimqj+5QaYnSs1bWGpKuMa4oQThJAV5CLGGAKf7oK/lf7iXa2kv96fkzh
YKcF0FKxiGdpVNQgV1rn4kgHLynz/foPQOSg2W33qLYRiLVgAfIAjY+sl9G2AJ3y
DsoMkFdQ5SSCpY8q+YGNoQhT0iJ7Eb0VERsMNLnRciCLel1eoK5qOgJCGbTT4aya
u07dUUzVskNUPhPhYDnHTBI8qv7RIhZchmA2m5s9rlf8rkWCEYvNLZoQkc2jpW9m
0ZRCkN1Icko8zwspazpTmqOKLqGt5vhRZaSsogANao6PKjTrb7vwYoE3tYJlb7P8
GGYO++fFUmg1F/bNP2pNpXhdgddpbTM5z+Y87/0pIoAMVnzm08mqgT0rRgqXkU4S
+00encatmR0vBaQqx3PXMxcklIX/stqZbHKBEYEhmHyjU5meww0IfSLiN+U7eJr1
zjssjsFY8NYptGjZQYhEQQZDQLMU3+2mi8j4NMMOCZvzsmgY266SEwP3wGEn5Ngd
rnu8KycdmAuDe5ICZ6ixPAYrxYqGrasdzNbm/2kDRNh/WuKE4idJvXRl6w9dNCR5
rhwWhXPykcJ7VseKoOVsLyB0hHEXMERE5hj5vIkdm7xoPtLHR7jZWGY2rH3ef1af
0MdfXfT+JyXUVXUcnAgdLVF4ItF2MwiLokripgok5ZVlIfgSQ22ykJ2ZyFeDyS6S
KdJHc9P2eK2532FyHjYP+EpDisggh3TJykvYKSPABp04E+LvfpmmAWz6Q6qfE1Bd
bIpWhhil6XnxPTmPpNreWrmmW91MdXGMSJTFA3EwWS6Z871GVusA49jYlMrjIZBf
UKZVsZs9cwgKJbaOCKG6DqUDGkoJM2i8b22xCyDkNq6SX6Yka40az7aaR00lQXvL
MpONlGPMKY9qY5Q9XQ3+YnEP9peHV2jVv+qpt4fXVCLr7p9/5XFnjPOJofVIzmTg
HX4B/t/K/A83BNLobZwJXr5QTn75Us9uNUG2Xgaj0VsxMxdo2YG4zc8A3Mz+J+KR
d67aVJV2O8IItXifv9LOf1vvaRMByA8jWgGA3mG/eaieN0m1XbSPCgsmx5zHiCLe
YWgMs85i1ETRLewh7GXuqygWdcfSprJCb6pR+yuhs7jd5GoTzGhaxUH8SyUoash8
mjWQ0SwVT4TSyHbAaYWaVBs7V1X20TKUPhJrPiTQ1Mi00cwpCFk1a+P4oqTtzCLd
H9NHazVnbLVBKVHLLPBwtun31q2LXFMOTY0xuBnEl2IzpKokmxkHk0kUEa4VN9o5
Crb3YevfS3QjU1WclpUuZmtztqflf/ZeM8phKUyb6WCs251FWsQS6kPysqVay2+C
jUhRAErDIxR9znmsFrsXV+Gq7NTVosDJFsaRi1Nnflg7IqKXkHIQUm8M4j3yx75n
s/I46/h+hnWRzYrVZa7OphbmzfYjri9Qy5NnHLCj6AgvZJxnzvTfRSJ9HRmIKBvW
btMEBxN33yj+kdYekFkndaB58b1zzLGenoay408FmmWicHBA6zMb87bCpLwAl5ly
XJPuyhCRSxg8BXW2XftKOhdtA5x2wcOQWRJb+pCXeitq5LGe53TSMWU5+fOzlVHV
O+Y24LkFpzwXgBmZUlurljSDw83aS35H7mfVBP7bZyJm8pnJDfUupQEarT3jsfVF
Ll+tEzEqPSzO3bND/oXCovotHBPTUxZN6rWZLUQSR2XQUcO4SVTfeKCJ3yxtGib8
XVy6ZTN3UsOObd0qV5bsagdxGm7dxHhl5t8Im1voMmXRspxYtPn+EMcXMWliVN/K
p/lCiDtPn6djhCAamhb/KHtrMgOrL7BVhV86r5xdtftk0aYtkuskUKC8ERgU0rY2
8P8yPM0L0rYwKsy+9GIwRoCduY3yDNDAVxyfDdteLAq7s86aIx7wygwb9/AFC/7L
xeoXFlfrEYbI2UJAic5l63ofZJ6ml4A59eUqIDBUfc5Qmyj0z437g9gRqx6Mx3mf
nqQPXRzvGSxzowl7KTrXRRlizLebVaaJ6it8L93XedVUn4m468+0YBXnmw6YUKJy
COY/Ul8cSjRkiI78U/oRV6l2FleHhf2Aodn9HQpjOSYZ2e2gjSNgFUZJu4QzpMUv
D/ey038g1IRhXoX3nyv2XJcaBjfL+v2lrS+sf1QFwXo+s85KpTAmiH8lztdRf+Yh
oEq33VWaKLp+xgQ1zg3OpZaj/pk/3S1ChqoeA4Ki0Ufe4TVcerz/oA/UrJUZL9gn
Zav0C5bUfCxtqPoD1HX4Qa0BCDf//npwy2eAeSj0KD8S/msXXo1/P3xBvY915D2W
6dQtaH+YIM4RbTICfSraGI1NjrRY6dOlsiH4r6b/a28B823DMKw/LcDapjCLCcH6
pvec9ihAzQSa7ODLMTSj2zqmpXE9AzNHBe+UdsQae6o/w9TlloK/ZEZB8fuyso2q
dvnudLQ22IpL0bkS2MGiQWFPCXHp5lIyOunB9R9Qw/M7jPTqhgYZ4jGf3d9QV/YU
yLJeL1nDRYbix0gZj6L++/8yWjyfkY1oHtwQwHawfz2LBVAAtBCWG0vIHHEsnayk
bNRjb/khnaL/Mmxp21wy0PLgjAK/Cng/OViKI2beloyOSqm6whYXUSdZjru0xShC
psN/yo1WYKOVfjpdT7L1e6mn7AC8XiiFLIb/mI1J3Y1mQ7hNhSU4wCc0fFzv50Z8
tcz+T4TZrtQ46z2PzDWSubmO8Dwa/vH9QsXzapok/t12yb5u3nlmtYmqQsWPjN/N
b2T9NDM3hHmkx2eVhwefR5fYV+QO3TaQXHIkLNxoMtex42WpyK+SRuKsK3cChZ7H
E3dYEHugkIoAlWj7L+fofTlQjSY/BVHiIWcAUtpgqKkjXZ4NiUC4rOc/MMLawML9
DZKEdRz9xW0Gn8xgJb1rqDaoYFvL7a97X7X6+tTPSrQUwT6LHwu5fuc6z9q6ldFE
QVUBiQxaOjJWPg8eF11W9LGCv2ib8WNsABmJNv61tpK7ON2jh11pAgXDVJoxY4gK
clQ/9cIckVQMaRtjNjh1F6A5ubpO/iAOis4Pa+CaE/p9xfyhOCefEIa1zCX2nZbI
z9R9kLtrEvJwNwRkFfB8MweCCjzm38kwctVJtSo7BWKUNrgmxxRLfpFD5HjeTPgN
Wn4zmtbp+k2pm5IagSdn/eAJBVvNRieQTqYSrQ00sVvRV8fITCQYSMlcI0j5WFcr
2oAQEHLrtf5TjkAaZ5vTLI2wUTlhUNJFP4LPOgBdNlhjAyy+y7wjxq6H6wbDyrQj
H8I0o10/POMl1BPYQ5ryJJzKPdFozOMCqr2p/WxJXT1/LzPFd6S7+6vyV66rkeJQ
5i/BAAOH7JE4TxugDeOKsW1TctXD1s9H05jt9bS1816l9q9lG6domILA7+yfR0xl
wSBj4kDjt9c5WFB3Da9u428ued3NFrpkRhK0QeG2FBQ0NRII5tivHfLEXXhMbz+2
JK1GqpAkAtBpeRop1hUgOgYEok2z9M3HLgPK5jIAzB9/QxyQmgkwhur+H/JRB1h1
qVLjMLAbdvcmIXdfvfa+77NdhXCmHBVNxXkIzB3yiCBQhlOuJVtAG+wRDozEflu1
Ss1faAQiyfdKX9brpCq8cjgLqz/I+wHqLuCM8OIUJlLxKb1SpOb0QmQ1+1PfrxHR
rgCkRHHCXiJrJS5q5DAeuJGHjRSHP10QiZwO8c72W9n1sdkNvCjmwsFwRh0P8N9b
f7fFRwMT9jdOcZNfamru7RF5OyUOXHehki4rNuE6pbP97KAqNb60+AYwXQU/+pg0
nth0J0/Ax8Vi+Nc0BmWrsV6T7Q2yMXAqwsDrsffZLSB+mCViJUUcth/6dOhrsxlI
Fi8pCYbX7edWdE7ZL/JA9xaILWHJuQ73iMfekSYp355M7JJvBFHHY6izkjsHPubK
mLyH5XJag0Jv6exrhTfbVdjE889a4yhmQKVHaqBAKc34mnewoRWQX3WqPU6yUA1Y
5xL4q0RY/6uHOLy5/CpLYzdtTwJIFoOLsb9NgR067yowREcMSTj0KTbvFVU6Jqz3
hdItTPiXZLrpBY9gZAqGJJeahiT8A3UMiUIK6Rd4flKzBxS5zdqwqPEhm2aTicB5
jC2CYc3UGNz7MXxwKyCEBN9XTSE5k7ClDFNCfgQ8OQJEKCipQDACvBMyfBM9910L
iXHqhE8vQMWnOQhOnVRFMlL5eEYfRlE8mNdeTGBcYlou3GrLqZ6oqzJzcfuHxHyD
vAOGmWiFAptFq10mzgQuzcl3jo3KXjeAc/GiiLSyA0ebigUqC8OIn+qEKg+/V2+R
drKpWOpDGYmJJVc4unVskIPScPDTZXhjC6Vh9OwA/Sjj181stnpy3WPevCaJi9eN
SuAmEoTH+qwHb36yiVsOVqR+JGjERPBntLwJ4r8YyqBe7Pc20iHUqBL2TzGx9803
z/bZJvyBp7uO9FqZ/nTI8nIvCPIZMm0KkW0IyoAHOV0lAj9j7/ayO1hXSJB0FX/M
5nLdQ8+vdbVFjpFC2+4e4HqMwAWiyou0q8FZEvB8DB0xq5eVw8aQ1LzQTFyr0QZg
wfh0SzZAffThbrmIYwePRH/4BUC8E0J6+3QpsyklHZPSiYnz4osyWOnVQgjKhTYZ
/7gB58qZ+IvaMk5+mNy4yaQkCkJ/Ls7syFZkquQStS4+e4fMLhLsDlKIX1Ap3HkH
kw32gs48pVIu6uOs/S7L2IuMKXVgd8y/e4bpOZBj2Y37QudpCZCm6tpjRlDasuL6
aUZJFoNnHYZH5P0HXBizIlD9CV/m9yO/M3nMj/FIq5zJ9N8cNZLGX2D7a+tGv2+Z
L2hNT/NWVKY9zcVS6zvTDSbXjq2ayO8Wa7libx0XIdTqBqRZRtzGUk46NJnLfVgl
SOoHfLwDWU2gml3Dz0+bocOPFAq2fqtpoACi1hodm8IdlMUHb5UwKoDx9E/2cDLT
8uOZBrBJSW+zny93vDFlcltkfZJjzFcRxrHWsEcvbE0JBU3EotZCrNx/ewWsHPkO
pss1jxaAILwSKyaMsQArhQomeot43bQf4cP9vhZT03ACSOhJr5lwhP/e8yMmqNgO
YGFi0XeUtrL2iMTl+qHMZblUvbk3hC4q6jhklxHYkFf9ExB2pgUXmSPdD80LLLpF
JfB6X7JcefIjsbXnq+qb/tDGnEEG/rpUErkDc2a0dZSdm8/hZavIJENOzBZaK53/
JKIWlGHjB0JKpdTGz9lOsQCj0w1oYSfkHAXL5bANnTOtTskZfG8zHepTgqXbGAv/
zSWVDDARhYCUkd3v6F3vwm3rIjs7L1xCp3/iADPFMwxu7VBuE+Sh1QEKkXT3bZ9D
/Z/m8PA9pqiAv/Lc+EkdUQgfZ//RgAYsOd2XaIBry54dImqMXpcpzDlVvJJgXqIS
zKzC/W/VvyDxzff2DloSkAG7b2FjNlqUM8hFo20XEtNzCvsDIn6e4/4gLdM3+lSb
bVySJpHMbO73dssevcXUhG/lor9w2CqWrbEEvEaWnPGmsTFqIufFQJZIaICofQNM
jyGXl7+ZcKpgfta0g58bT9rNSdDYnNouS6L4mT1ZDgUzALAflZ9f2b09Nkm5GeLv
RGcAGyyD07jhHgeJGlve2XS3Rfp2UsXq7GTIb31+U01RbnFV08DLd0QBo3gBoUnH
y5hyfZ7vhWeGuzLLKCLco/vkFtOAh8Aj3SGSQ/pCpu0Im/aor8R4HbVelfgC0m0c
O2dyl0LRbz2Kt/lEJKsCfpqbAylPwd/NU/Q13rjWx57mPCf/AjEIvzvLAomy7j2/
wPw1/FRHwY/B3VtTkJUNDNc/hXJefc6BpAE8QKFltMF3qCW4hoE9QXg6I9D5E//I
fR29rF7qQQD88x5E73YzU6AMVVQiCA5nFnF6Bsi07R6Mht8nO2q+33K0vg58UltV
SZhWUBLY4jxHtUC3uM8cqQkJa7zM1x5y9175xyxlj+A3ZQiYb0GmhSBcAEApNDiK
bbfgrPAKjsmI42b530yG5+RcRYI1fcmvcFdUWA5THW66cEXR//oU2ma4yDlmL+g5
mNW78xo41kW8XMl4lJL0BSxaqX8IacF0MtTx7oVG1ofckVH8Gynxzpa4mCZeZAJw
Y7OtdBGw8XAOs5zeDXZw8ikRiq+s8bhCVwSWNd7E6WK9SxcCmKVzDLvfao5rFSG/
xWw/6/Tt3UJBnyEWgl0TCC3UExzRFR6KTMPNXLbyiHO3HPvJTzu6Q9++bUr9/gjV
e+spa31MsVt9tXghk0mPKWGGY6pPWw5SSoLFdqIVgiqwrC2VLgykOFE95PDttRgc
PRIFrmg3Q+uhS5Pun0ewCpeXAPlbtpaNJtwq+dU0tkhIbcttjdmIZbOLnaH0Yhvo
JJtggYBE7mKrobbQf2grCK5S/gkl4bfQM6373cRksNLAzkoiR+tXH79WlmoQVCbi
iXv4oGRjl2ZWngDAfAyVkBOOn8nqzpS+fpEyFkgrx8u/8ZZHN+wNOinMK0yj9wU7
kBwwQC1dJIgg+PXqEa3PJwHzp6cGbag0x5T3dKED9W7GBqXV33mVG2rklH0Iqf0c
dGLBLiDnO2BsO5cOtEzoQK2mGPoR8MbkSOKLhOg/AjHlQyXwqf0UfPtTlkyQMOBR
BV3uiNhveIq72ep88I5DezmcKcajTnU7fsIO+sqZh6P4NTaXHYRnhRhwsZaFTEd+
NwfEp9WtFBRvjsnRGH3zflBjW5R/fLB1VxVLAq8cBD81xXnvjoD8EhNTfFEndAkh
qECdJpncCWBp/b9pCMDwiPxnp1yEKjIpV81LnuqHlyJLoE1VXJt1LO0CsviSxJvE
Mcz/EqnKN5LvV+jCEAlpTZoYiGIxacv6iPg8as5gxExZ8uZA0dUrxT+SSBDveFt+
w/dksSQpzrq1AZZa7z13SfVmKfv9/nZsvbWNbGucicJY/7dJB6G+A5pwNLZrd2UA
iiviUe656ywPRqKAYjnE7WJuuRW366Zm//+BseI8szpIXS4QJHnov2OTY4K9UPkU
XON6O1CyIFDZP7Rv86x00SgO3ONoOIt+Pg3wTbVX7Qk5sD6BCynQ8zyfQzO9KCKr
cIrUd2wmznZPaUClxzUW7oCOxbGh57karRJk4bvTyGMJA+1k9ZAZm09c0XK1sVXI
b2Sr2ANPT1tBMSdaJkDNJNwZ/6S7nWwd/H+n02Er3wnqruIVZCv2ASwlusZHwcOu
SnTSNJ3XkgDGIQtWGXud1B3ttPQST7gJebJ6u9KZofx2ExvrBwK2glm7rZn9cpsU
qY4MQk0V68ZqHsrrUjs5I8Tk5IZ73cX4mLa+E9OxAajDfKnXiq+YgW4vcoBwGKVs
SbMjhI7EI63nzMcfm0BqEJRcdPNvZpg/tGe1I5CIAoSOs97WEPj+USriIqz69Uap
uZNlip3pgBsS06HjLnor9ASCsBE/8IZE7ZjGSy1+CeDyBCAdj2QLPpVFRyDsfsQe
x7Wgbphid5QbzuXQl0iEUVmsE7+MZjMuLPNdQ8prtfy+SBVAaPnuok+Znr4FjIXZ
qmSTyNNB/rMiOXSY4MrRinyR9pNC9Zfp23thEcBrUU8M/8dkJto7CKWYDDD8eKPJ
ZNvr0hUpnb2zENoCfLI+Q6SvcBCsvyGPf/XkCibufHJXhInBJ3ai9/p+ztCi2tOa
VDUM7yI0Mejeo/luFSKD5F+FtHMFSwg+UAgSEMPsg47e2gS7LqLetGBATV+nW9JZ
CR5iU9supdkUO1KuiDSv566XOkGSyoiCNPkPrjAoqfiN0uetEfWN2IVPEpGZ5rwV
ZkhPi8R4wb0y6GQcWFbPAhQResQH1GN1dIBVie1Ste3SpWkZnnhzk0avEppqSWGA
xjbkyseVN/G0RR6UbsBgdCjRExxX7CHkBxmod8CJQkwnt2KiOHagDlLHe3BiENzs
kENWO80b5rMJVaKe+nP4Dr4lHuG5RzJhgqXFPWmL8md8k37j1KpZVBJhBeFuAicK
SlBVyo7xXqwdLd4YY2hWPNIHfMZt3WjMcDSlyJnNZSjaLRqZ8w+G/wfrZzZM/q7x
InVmgkTA1pYZBkQefE7zLHMPdef28II5cWblTyI9P6hSBr4LhmMnf5CSCUJ/81yz
vCMcSBor/YbbswvUjVFsVRyLly8W5aGXlugbdadlmfhnUACd6lRpY0lyG5sBhGUw
93pYDUHc62jUldBa65n4huzm9P+W71ew9VbEflb45f7K0zRq3suAj2MxgZu7J4Mp
8Ec5UI2Bcl+eVaEWH0e+NvZDvPGoDhySjAvV5u8Fve06+E0R3N88butDhFDxB14k
7aLzEZvt6kdHf5FgqboZCrwrXRXiDVVIOsh+jrN13SUUEJSrFe1BN5MBuHwIvOFh
K+7AuRM+KxOipwR/pp2ghVSrE1ibAk0G1OeXBj5MV41HkHqIDaTozty+Zan3cIWu
0qAT7D20oZHDb8ZbvOi4QYcbCIKhVwqxZRweUhhKsZSX6CSvxGOzlxD33g6B8gfj
Z5xiyOYjfqMX7SWy7bQ1fTn+MWfIk79gr6x64DKNNNJ1EbuPQX83z3A9Wc4ddkP7
FTB5j5A+Wy1LErcubypzf81nxvhBDDYdjT+aHL8kdMNJPCrOP36GRGYf9CXKUFbs
sFAKZZMh7uPsGpdNe2FpIvWtDrWHn00hu3kdhPTKItwH5x3qbp08lLc0IgqDvwI2
GPOf2eojv0KeOaWpy5xdL8FGKeCkEaTV/STsaix3r5TQYrKT5uvopGfc0fS4Tb/7
yjz+qH3P0P2sqrX+//Nt/hTfgd3v763CXG4md2UJcbsfeUVNcxWhVA7CpdCIPSUG
y3S5oBc7sgKV8t/WI17Q1Kx/p1OeYHAW3GB/ExNpq0OR5E70VxslPid92CN56uyp
me8r0UCE+M6jvuEXP4KXCPt/vZ0oKQ5sxFl5+itkcv1qgsW/euieopmfmW1f04LU
an8ap0F02p3iUfa7MhAwitPtJU+F8nXkCPEvdp0UBvw4P2BeZequN/NSDgYnfuyc
9tn7PsCXfh1ATG1nCKG8JmCToGCjNZ16rN/djGmOAObt18WefNe2C49ritSfFuyS
QF+RAQnXePCpuAEV9djzviCg9xHHMfYK7WDtj3vnNd9XHH/u4EFhZJZi/Vt8B/20
NPDZPnMxWPEfg+9IfcOQ99XOSqCEclBG9m0Jrrh4V8qwcdrZFlGLgpxrDUIgCyeA
LxRo46fVkNQsB0lUzQW2djsZSaxu1XGGUInaTAp/8geS1qybj0v+jWx0clcPYCa4
7Fby3lmRto6qKFADa3hZWg31XJ/MfS0KyDsXQlI0kk76Uor0xLYr3HUQkpAgnE3B
vEWSPIj+JYAK2HBYlAqOF5faEUH3epc8rLeUXj8j5LOKYFmamO+jHvh314CLZjLr
e60W2Y/md2oXEpW7+h4G7qeVCkzMWaGMLdZ6aRRCmCyrNEwO91kpR/2hmMrl5Nol
qpauk0OYInarnlpmCGPlWkvkbn7qEJEQRpVFGw+zR8HUBT3aAmL54E7uov4B3e4S
UmES8iF8vppF1EnRoncb3xamLtJPdXicHYUD3BtcwxXN+ECaPnD2DMKYfEzCmWTM
TyASWV2qX8GYqa5NvHaUT7aA8ByfHYuArmkOtJJHYP2wN+xlemYuOkpIJu591B5t
arQxzOeUzRWhe8r8xBqiI1b7ztCHFWXE3cSXKMSxX3+c5O+qtZBgiEJ9Yez2BQLJ
2inpfESjkb0D55PwEB3OMsx8ZcT+SdLvcRqAc0876gb+01MjaWbj3D4HpIIbCCn5
rg58wazsMQqImwvMHtKqs10kk80aPFjvjFwwq17mInbUXNWUrhEZC9NddD1p5cxO
+DFvpIC0J+uGVUFldZyReoRiBWorQ9iBGtIf+Oe3YX3RYT5VlTTMCxYotF58Tpgs
KPMR8K4wroeoJsJs8BTCq4Mc6Gfd/BRV7duzaIXPC8EPQImP9JGtYRamRVCJMMHp
TGuMJmMKTHh5soPsA5KdCysRB80+vzloy33vKuqW2Y17Az5O2651q0y29adBio0K
t2daX6Y4uLH0KpDXjNeqT2vbNVo0NXi5eaSW7sAoXe8CeC/6S02jAqS4ll6ZPJjf
CYflncwZISw+7HF9PNrwiU0g0Ha71S2hT/PTiWxRhGab87BZ0w6ykEk9PxoEDk6a
DVc+dt3V6ZiIDY7iEEPYzu/FAUchz2K3xSGpD/OHJm8FN1r2kjuwvfic4IK3mfCy
tfZxF2H2vJLjT7JGr0JIg6LkY92PhZnD6eJkoKA80cm5us4ncr1jqS2lMTxsGIRm
LWUlsrNZHPyFpU7bG4gzZoGIJ2cSIf5ZcF/a78PImvgW1dXlYlWrFFfwaykP24+R
nbBsohCmGuYm5OJwQMlEcL2ZP1gRkyc8bNIewa2mKlZ6n/+S7RFBaSj4WruvXEZm
fQSJhgtqHxabFbWO38oQBH8QCVLUsuCl4kWSFsTqIXIwKQSMzjqD76CBh/9D29+l
A7kz1BQHi86EnkB/o57bLTniZvKUXku7W3Jc918jgDxK6kLWPaxoG82eSmGs+sNG
dkjJTv/jm+AAW90G4SosFuPA1MBpkLcBeONetww0N6t6M7aEy1yxkimOGmXPptNj
O9qYrxVOFGf9d8EpP0baiN0tEiLuV9Yk2nRmLDderNHwxKEf97JN2Z2gDTmGn3eO
+P6/gv/TbgBykPWUfdAF2C2Xpv2pGdV7ySX3LDW2ymVfell0BC4QopbHP/qZC7R4
ahQCvWpKIf6RAGvqjulAvJldkFf73k2Rfdd6tVuucSSTxYEWaISxR1Ab34Nu22jC
OSFrrRKuLJvWGf57Vu5bG2eZCZDG6zR1BlP1uTRJdIN+tN5+0ReH4isqoaz2hvex
5/ytCh8rjd3E9/krbYQtgLGKosWISkughAxxaCQrTn2HWJBtTf9t6nmdPFaDEfT8
GuoayRob1Ekc+yON9nomq8UZb/A1UTtJ0Az03CyUr0Zzn+59wAecw/4vU+/thVy0
XtY6W2zbz2aEUZ2UQPQ1V/A62O7nRYhYdAsNUuvu35kJH/KGwl2QOLmR+V7V+Gh9
fDASCJYgOj8urpGd1+0Hqwz17ouFuTnlpKN9wbL2eSlQBXW1qWvYmPhBk7k/t/1/
C/s9GMdXU7AaxLmOg2JZGWwIMtmbHH62Lwodr0zaAUnan7IHaZ4lg1mwR2fkvHRC
OBeIenG3ITNZxeM0xCBHYr5WjTN7OTo8Gi19w9tgyeCZ6gf9+MFFj7VPWDRN/d7E
P5MthdNBBKTPkCw8u7se+adN4FMBQZSCr490AAcPjGDahXUFi5dJFBKX/C+Warrh
HR+H2ddn74X09oMn2+xONixqY0QDILL3W5ey+QPftnkChYDbxVkpUuJvJQ1CA4Fi
m4AivYNKGIKimEzwG+KKEis6Ak6BaPxQC0vIi3G+XavDdcn8lr9zvJ+P05J9rMAO
L9cPjlnLzFOe79Kv1zcv25yBTN+2QqE8brdYkMnF/YO7Wo4G8kfiMgYb2mntiLwc
xQTfhHctjgFRqBjAD9FHg7OS10ugVg+pNxHE3kEqd1mv8L2LZ80pV6EJ9PAPs2c8
FP+PRWPQIRK9xFLY5E86w2q6O4OVeey04WY0JxmSbpZGjdLIUxa/PMIOdZ8YV945
G8bWWvqLafVSKMNuj2goVcbLbLaL0FkVbtps8WYENpJ7Xrz2khyZaS7+li7I8vTp
HnIF4ThKvU/BdiZvViJqQBXh9QWvkhOBgwjfpBPOVkMIBLxoK2ELhzjolLM8e1Jf
WxyidA3FY6WCz2iK40P/4inFfN5ZdZoS24sYJppso3R8IyFytVeYIcgptzHkzueT
FAtkhdTbyBeVwpXCrVEUbfjWGuI/1YecktP7VdKCR7MMgE/WDZ21sYhI1IW+f3jY
gj4D4lcCT5jYL8OcjO1cwLoZorDZ7PVG2fNF8A2vW7tuQA1fpUYz+tDJCoQ0Y9R4
LhJM36+4ModbwM4xBhLBu6Jw3RCpveUuNcQAe+kmcjeFIMVlb+WQeeYkh3ix6kN+
lyES7vEPUWYHsUcpFojjc5Z5PRy6VdUUNrEiX3dJO/4CASO9zjehjYSQb8fwNnIs
Y9Nqjt77igeVX+0cahRSE77nqZy8+GC5hVrDSNtgw+7BKM1Hx8BHnnzdkYU+T0aB
WxWgFrSXngH5k+YrXzY+VemrcpjoOxgo67d3GWiNIJ96x/7GmWcEAEsHWN4dfZag
vwXjP6tfsNrxcz2XNlYn2EPdY/YCk83qWQik16uNthsjrnA5hilSL7tjCqko7zz9
mUKnX5CBGwBeKDnzVqTCXfXAnYcIactW2SyLg7YDjGBQNklCGddyWQZmF7GoZRg8
yemMgilvLWE+LjIw/aQW5rcOE+sunq5zFIT404hNNmwtXfFh6vW2P/vOPFMsa8Gp
pM90W8KF87IMt57ZTcqgjYAGE2Tzer2pbXo9yOaMMBfZvXGzPmqlLKRF/ooACLKI
1ZcuHIsV+TpAcBXXx5gOcCSdMEHub32QXHxmBtZFLmLpDsK/xAnC1BCqU2nLLj5f
Xo3Q9Bl6iUFZm4QbgIvLu/tdeVPt7gmm51H2z15caCFdo8GR8fwfQZFs7TsVhZIb
yTAtFIB8pTThug5knnjmfI2jtrA4sgMdOIsLjvHrnPNnc2b1Xna90Iotds/2ITAf
HuBfGJHDj+eJhYkFoHW0QrG5atcVSFnn+FTvi2nyw1BOFyGCntiU5+JZzrfLtmYB
Xc7GxypDxciGboEnA3MQLoeMZAO0S9K31RyKDCv3LlocdqE5l8/XykIgMldJuR2Q
zHYiI2afVex472BETwwhqspqM/c0nJuxxeOzZHCbmFJsB48bhIEwA+0MvxGol/co
VxS78kiMbxNNT4l4CX3KEsO8qzn/ydHRBfQFIwI+VONhMMKcBXAknZBqucs1MDI9
ODvJZX6xTV2DRShVs3n35Aa/oCmdkDbYBaZT8nAOCEK4+tmM3NLt1TVr9HSwT3BD
VRrRpYGurQ3nftsngT5oc/JyI8LfbyqYhocebxwJNRARWXs177u+HZ72Xt/HjWpr
sx5qoRff089nROALX+mqq66HZpJC4PndZbuLO1lVUOzLmTPgMXJPYTBXo1ew/+b2
Ld3IbRP7cgiBr7Aro9t2IYsf8PPR5DtUKWN//20+/vWnpF6No2ligH0gdw12uyGC
1NMybfUB52qgmfMkSvURjpAH273k8woznYBG+0riBOPE+28VGxDt7v8Jx6pwq0Ra
ezamzq0HZpDL6oPRa2TVncoMflc4ErPrjrWNNudbyKhEFepxgCAd56gdOPSYNq/f
gJabmHmGlYxGsy2+13zjW/JuYTkGK1OW5nf+o/XrHTYlumBpxnfd/G7yC4GC/Qqj
7kv5knwaV5qUSUtOMP0177JdH00bBF7pLfUXrq5JEVUnaVmNRDbw0bubtMmUh7vf
JeydXHct54hh2+xG8ct0dqN+jE37z9RpMpr6Y+IX4jY1tKjgXLoMts2QxMXf3w5B
vN+eZi8hN2v32/l+E7jG64hxxz6SwZT82Fn1el2cz9nrx7aHc90LeRDFHAJ4OvAA
DCA6Ew91/Jp12eIBoHOf5TLR2GITu+9bWIwL6TgHxNl1dnIhEjqRS2OyVTT9EcMo
x+LYcCoQ5v6i1mF3jEBYAcxUlY7arBa083T0eO8VQymscNjZfeenZ0Nm5DBoxcRd
vCgkPa37EsKt/EXKbUcK4XZkGd8b1HFN6yFAcpICkk7BAP5Pi7OVfDHOLikO1zq4
47sOg5wTeRPhW7JwXLzFUh/O9327rlyl/u8m8CWgMk3ibQdczpjgYlZxBNuYbcab
+h4rDXYSG57C4oUgii6Sb0ogQ8pYlqelOQvBaau4Mz+H7K1svlUQmGTnd3XtmRTh
EdGSPhAInHgyB8D+mQI2CgDBoClfd/Nab6zkAFjdIKzmL9AznxdaW4j7kmatvmKR
nZeQAN5hIxD5mzz7Wql4xscvAig/VK3WRYO3kCoUfcFiYn+BX0YrMLbAyE6vTjCa
nGK5qrhjxDO+e3jo4nfMNGCLVloYYbKoAdqs7VOzcofBCnt0qq0Ey/7lDkX/cOAV
9iAyUr66T+L9uWgzOu8D1q+vMhuQDvMCs7C/Ap1rq11cZ5IieZyvBXz8RGfNEJ77
RN3jpfTnjZNOPeF4ST4+7w7pZMRRgengYc0OU3OH06UHdg4CTPKuIkBSSKMRuZna
4wJb1DY91xnimjXUra9U2NReKWiZBJNZ9mP+TK05FxFPHa9iiaUcgseeqXwx1byI
VI2wMvjDwEVAsJoUNxSIi0Kha29HPefy85WTfiTsVRV2mHwp4cxTGG8FAHNmvGJG
vpCRZ/92sSZ/Q19prF+JqaYSUpcOdpqvQ45OyWsd9Mqv3vH4HPY8ifalcGnlCYj3
VMhjctUZGTlqzmHNLZQ/Ng5VTGUPxleYYbjJ3Tup5jcT/eNaOp8epN4Xq5Ux6k/n
nTse7XvhlnRE2FDX45jCIJv7B6gwVXfLQM+ekqPCKaCs6MS5g3dunSFKn6ILq2MI
Lb98bNq+2ETekLKeP5xDhTrOeAoe/CpvyhfwUC1QfRUV7f4JYb5eZzAUlEOx+BYu
Ja7DfFpmii01oS1SzgeduB1c7uqd7eHZ8LlqdVta+OvHMvudb10YVfcXVMHcLDH9
GzoeXyhnNgFIXMau0l2w4p/4V/CkTL6WhjftJIburEWAYiGoG8sioLA9vNaHKXi0
5AxOWVS9k4srescY/Ijlr5qfZKQz+f2QKzkKW22wANSFd3YdOMwuRNTVr/bzuiEl
gIDwPpCMfiwYb+K9GWUyp9WUIXuZfyd56ZC0/pFOYvaSTYgETybcyC9YKs/EXOC1
010HbKYncpzCJ1FGUoot9efY+TrM2HgjOwi8uuY/yQda2I3UW0cC30gR/UItTMXM
zizxNLPAie63PNft0HVEHMfS6cEb5B/UogJqWj304m/YBBu7KrwLXFltKg0A75RR
mMkxlCtBHLMUNcnL5CedjB8Y8vwoeCf3xx3e7ZwJVEUf+MVvQ4Xx/bf2WVDZH/Kn
bHoBdcxKYp/R3m/f/sMaCmAtDpeNbI5jOV7h921B+p1h3XrBVZSDGl+sVxIMG03K
zoKb2edf8uh+YYmmeWqtpjMWhWRB7fhxqa5l/fiuaKqKmWp+1w/Ax1m2GGr+yFXI
UBO4x816tqkQiBu4pv4fBMILUdvw+5v9A3/rrkcd2kffoBHLnyPCPT8agjvsH579
G9GnDX0nsN43S3ON7RXupzSRHf7CQNKVMTDiFVlokZI2ZmlS58OhZ1RPfVYn2Hgk
cYCmA/3W8UFwUzqML5QVKOtc8PIk5wWbmDS4si2Nn+9z0zAGd6IqJqOPMybHDN/6
Joe6T5+FmjjGw+LWrKI3N2qNJ0a7uayhRKqZMAZ/fKwcJF/IL6IiVaqArWNmymvL
8yPU2K3BT9BFOzCAuybu6t5+zgDuaewpfBx/rhP9+UQLaM9dGIxsp7a9ufEZLrm1
cDcd5ubddHMaW6VvHsYJkuRFuJxoPYpE++UBBuQ3MpU6spdGcf+WYvbUboUQ3Qy6
sIXYlUmzSMhLVNfqE0rqHsZAK2bT6h7sE+5E9e+Zttv+cmuDC2DH9vO1IZi+zbxJ
goCwx6gnm87ifsA33+Sgy0h5QcP00KJDHAxOj3GFKRshRts90rrJ7Ds17P8hPx5P
czmWo+F8hzmIorSG0zrRmgnatW+qTcUbCLcsZjH6cZGDlMEIeIQT74DTnQE0euM0
xypuvLkaAP77Vlbju3/1rNiKVTskWnNxkSnM/dQOV61i5y9qrriHhDAyGZN3rgiP
eUv9OhcUHgdwMpNVVQLtDVS9dxAHsnIYl2Pei2dhyXcUTRqfmkkSJ9/C4wdAn1qr
Yv9fWlxqWadVs0xWJGe7VYDlte0ksOVYL3NTPm1i2DPgOFtd+rf38Liy9yyE6kLf
qOYAEZemi8rBadwcQHkIR46aIbGEJqPB2ZQF8FKi0JerzcL28g5ZDBFqo/AgLYrl
gTp6twdJVTuHp5TXUcCeZOEMLH5/oburfJfjnwy7d8oUO2/aGOOhuTyK0sMWrYTd
6Pj/WRTSTftjS+S/BHUanhwoBAMbo/kH+2yNAvWo/lqTMpNcpuBCXC/BHoXyds+g
ZsUcXEhdw6mndmUbOfCPH5viSs77qx4joj5fy9mpTF84quHy22sBoutiKmcqd5b2
WeHwk1gog1y0+EjUfnKETEaXvsS1xLvHjF4/ktTu+sNcCsMEFuNw5PahAu10HHjd
aZ1THzOq70ae2VOr9YEL6MBoCauKvMSqONSe6I5GY/4V6WuiAFLEpH/hY8ZeMqdH
WAIeCXRAwvGFx9Er69afNPBf+G1xPzyQwpvsOhj7JPJ4D+ZqXGkFmS6B5BgC4ieu
/pU7JtQvTQl0erBbHbXMTI0xfMTfo4Df4+B2QxLUS9B9ZSZjnnAaCWPdUb64ker5
Fsg9+LRfZVVl4ddMpw6SSR9A1yo1yGORujYJeMu7GnWGBmQUczKIpONQUej4lK42
IgPAQ1UTgvic05ReYH9IEVCFdaCrgRGgXtbRMz82+vzmBL7wK3x9vwx+ROHNQqJi
iNKX7vutaXti0lEZlqBMIEpR4R9IuQmFWvO8oQHR3SCfyaABseKBZVkr837UbRTK
dAaWZbfhSTJOn5LuKH846Mbj9dckxb/OC3MeJ7IcpOg6F3ih0uEm1ywHuor6Yt7R
zjaaKl4QwcWId21q/fi/WLOn3FJQ80F1VJx7o8bKIHtkx12NQ/4dstYezH65LOKn
ZehcvoJOk30AupuvKuk6lpony+DRuFP9v2gKN8fjBq4KFNIvuSx1l5YR1mjzpROo
XIrsM3l/azM97jvLzdDEhvUtdIvLtzB5cGZgoqJMqQnN9qpsKtFpxKAmSgIbNoaZ
4FeLpC/cTeq5KfAeUGssSHQNp79JYI/pjHTTHyQeKPtPOYa9kRX2ZjLhmwQQL6E2
i2Mpy0+iOG6S7k5uKidsYmI+5vDhRVbK/WGoS0lQ1+m6FSkbzXL1sJLHTfSkIx3b
O4c5U6yMkbHQqvZQKiz4AYyZUeFVOcjhm/vDu2+4YAqpy4zY29+qLYB4+hDx1Ccc
obb7lQ49PmdWpCXYpjxZHG9mUqObfBYqmNpM3k76T0f+0PdwGuacLTTYS+yZ3B/n
A4m6fu3Ak7FvNb5pWZ836bmh68xCReJS6d3FGNiSJKqhEI1Ut7htwdB0jX49M14L
bqsDKqRCIzksbC3PtCorKYNqL3shsjPuEWYSfQkzqZ5hZFzgGGsVZuWsOiOhbgJu
dKDSWzcR6pUt93ylkFwRgElT9YV3xfafHF5jALejQWH0aGRSZ0NrkwdeTUuWm8vm
pKDkSay8Y5LHMaFLe5xoNEu7H72rCP8bcNpvGtHnLknDJuLM8QQgE3iDFBvPizy3
oCeks6estHUYubDXSNioF11TrnOLHl08p8b6OP20LTMi3EQSD2uoOPUq1UdSstGt
+FZHWtMwvs0DwdoO4nljpXjPCUsAbSIDC4fLK0Ejke7odCI8X0y6lGfVlCrz7r7C
UjVJycjfv7TQWS/ZcuFCJjTbk9077zy3iI7BvdkZei2GSLTM9w8xGTav/VUsCZVw
GqCiQrBz1rVz4M9JXPJhnd+yxyVSyXcfpJ7EI4J+FmVAOGsz2tCDwpTS/Fn2dAxu
pO0z7LPaJzy7FcIvQW+OC70+PcabBQogXbgIqtFZ9SOsq8IEHzZ+c/RlG3jiNr/W
N9XPu3LbfC8GC19wKcrMz/W+PL+ykt7hOoFGYDVi3t6Yhg490UG9xc6Zsb1B28I1
wpXFzHU+rvCyD3pskZg3CE2wNomAsyz/P3zKKhE7qY+kEd9VRzKK1pSqpBVOF3O+
MGaHN1+RZChtr+8nP+x+Qf/aResBdTkyNlGQAhv8CpUCNUoDNfxIsEdgs9rha+ce
7JdATjegqwZZwWRWx7sXzYk8LLANBBG/QKYsgxETd6XbvreUcrZV2lERBvTZki+l
hFP6SJyyv/hKAZOJlwUee4anX5Pde7a5aGetvlK5FaT33WrATUW51/9dTnow0459
H7BjIi+0e/dMUG2uuMAmCppqo8n3SI6r5f8ttAlp4sT6xg62eL6mQitVt4zZ5LB4
dW9ztILr3fdioiHuRWmp7VpS774/O3dZsa5PyHX1lal8v8vMQeissmnVRQLgF5iW
pWQ467Vao2cljlHIapb4Nsh2Js5eyk8VFWYzEJj8pz8K4wM8Xg+8NiAMSqI0sK4y
KZzzcyf68APq56RLsjyeZK3N6sEHAdlP/DrfQX04OFNG1sWxX+jDTmwh6mBcm8Se
XUK3rBmT6kIuBq2USTqXRrZHF7k+rXltIPodmlMxyROv/3zAnyDOz/p87oTobd+P
JZWtjcSsGTVBP7sgrbGvmVVloBwicv3/ZH9MZbCYcsvK8w3RqPyaqKSegvSL0FdS
rZQgwG0MJet3rUlIqjSsfINHsAe+PMxM5nLrqMXs3h+nLkEhkzQKL/Hn51D0BvS8
Yatg4nH28PTc/3HzHLDKIXjuNkLBMUSDBA+sZWl57cmzsZQ9L+B5G/QKwb7U4mIr
7zUg+Q1SKttIYqPlS++rIY694UkQYMMSv2lDhqQRD9x9pZSBLxf9CDlAkt7PMNOD
tajwDhkLx8op+3Pz2fXYSCQaRRL5yxLi7RhmTVbg9ymsbx2EONCbV58VHd32yupD
xtXxsi3SDTepNhHwj68VgqdvbrWMTTyihffh6Jpq5PzbkpIlNI2Rr/Xiibpj5vdX
Q/63vlpnVyyX/p27ke9xbMMldKB0/1PugffTY0pRt8Me+QrPeWhQ5p7QeMs48tSu
dwnq7jcj4aoYSSq8tuQHgs9oiUqkxIoWefw7/TXoU00GCAWTbTI6NuZedaWeV811
eXiLFaHSsrfVr0mt393NGtA9Qug3b2uDcbAw7wdgwf1RgY82PAn/tfrFXG855t2d
7JWBSPreETcvfYkgnE28o+Bz1fWzo/L5N1m60v4ArotGBTeQ5EE5lcem5HJltLw/
iv+A9YNR4Bgxt41+EGEiJ8ENLUlQe0SHnUmmw89fShdyYEwcvnDOhfBwAi1lyAHJ
MwoYHWRv8+b0dPp0rKhRKRHAgby4d4fFcXI1cDUiSN5rm05uYy5iFJR61kdBGC1R
Fp+3L/63C8Ge5vyQCWAhckxcHRhIhRmMY9iWqE4Cklotsx1tqtb6w7fKF36YQErv
6tyGnzpawOgN/ebb8EF1sTeJVdEpc3XWFIjQX9a+OGG6RWDyBpxaFunUJTuCBhES
ywxiklzBjLik7f8P9CR3o0a1KLCAh7fFeWia55BeByRZswVUL0tXuFR0i+EJp0ph
AtmX1I+CxV2droWHR0UvbkO3Kdjp82cPy/o0s2WpshPlIt26lCVL0t6+It0Qm3wS
xVy+FZoF7F1Ejbex1g18mw0uVIPqsE4UYozPtI/pK/T5uSCIREW4zfF6ATiwEbU8
ML6mHvCSzRoX73copolOqnasCGOkF3yySWWicQm/FG9qddFg2DwD6Wv6+MlLtZrA
4vtxCdQ/P1vqrv4CcsfggvLdDyyFIz1eNv/4xv88c/mxyvdEAmMpL5q8SSrflasF
El41Kqu772TuQYUw4IQEYg400+HprooSR8BxooP4cDjJTg5kKjOU8JFnQzame08A
AcVnTjUEptSs4S74Z5i0VzMkN37IL6y//ww9uPXGD7gKqOELZJNphJ8OHOtL9h2E
uk7RrHISf5oE/HuxiihGXgFvDxsVZP0Mb2RjQOkWlY703kbgf60XoNKRokwe1zxQ
mkg1GIRwOg9+jC5XYNP1x6QGeXsXFcLmnT4CTeGIByaPVnPpMHIuRABYXIByQosP
M5b/h3POtU+f2mfHCPZGCMpEruffpdqPM8MS29cmxZ4yBneEyn4CY208OPFgzkTN
eS8tYDDFXvJeALjUSW8dqHwzi1CQ9QqZgNOirOjK5Mh64rgMuyIOKsTFJ7vE9i2E
Pu0Rwyr6JG0UBydPmW+l/xrBoCDf2x8qkKcnFSXpqvlxNvvayHjhEUw4U01a0oWV
cZwK3YYdtIWbrFOth1Km3fNwe5xki3GVluNkjzTNikA+ey7IVma5vn9AiKcnYSix
F6lRehs1sJJRxuz65iqrXxfgs+eIA89MWmPLPzSZccbL/iRwUAQ3CVGTG21Grzw0
+IXnFhkve23va5YpbHLFzHKOpUk994AttTD6014HKwDeVpJIx3Q59HBePjL649uu
mXcKynihdkbQc4wev8wDWndZk6QQRrR6UuRrvZ2M14Pixd55FEmphSMLneoj3PLX
l/d6+j56wDbuQa7JtLp5U9MzKzIC82/vv6puAE7w7SGRDqJKUHYJgveHFSG1MQGL
5OkTBmNckOEChTeZ0blCOTvQlyaPr2HBgzWtLx6zL5n/1VcfeIez1C6W8Icd4FBm
Fua9FRVEwdiv4nLOYVnc+C45gnhija++8Q+ZYiHfhSf5VznS/oijfzBijx7WXOlu
ozCOoNxY6AMfAFTJV/oYKbNs/VAVEBl2PWJrnfefgGbmxEFATum8MY6g59M7T3rF
ny+sfmU+8qJGfx1bGS+H4/LmFA4+HiMFC3fID83vOWgZLoc2OHNWvq8gDKUHuk5q
XZL34EUgMAyKaM1+peQoH7tPQYjnkQwEl1bPHZsImw58oxXBAn+CFb5lBUwWtHLv
AK6jmSTM/1Dy6nYpZKFOKEU+EsmSDc40Qt9/+ZEaA4OqT1L0HN9GATAuvUPBomza
2yjLHSwnkW9Za4TUHfp9nqTFcofWoqTBmmPTlkiGWvo+/6//5bm9D9Lyc7EB0ZA0
1UvrvmrrCokkQlf9OImjWy43Oqvnzhx+Xctz54qhliSUptkfNxO1EDvJY44j+pKw
FRT5f3Q81xdLoZP4aUtcA7Jni+W0BI3tLVoX/XGlZPlj+Fnh7i5CSt4ATXrxs2Wf
FqZA5371q0GeREIVWjlZQTtAa4y9mWzLNOFFTl72qNoCIWX+O2q3vM8YWA4B3phz
yHX0YZZDqlqV6gCc26CuIcLhgxtTUasTmBNF/QTswX8rkcKF6lO62rcIgCim8OCe
NA3CXFm+IE0VevKSNQB2QHggwNlH2T1sW4hPMhaxx0b15jSrzwrK8FJTgFkwTuft
VQPfmfkmFaUq5sc4bXnUUF2cSlQYAo93/e+4o3x/X4TrTLWPj/G4ZklWosnxkVxv
toGk00UdJ2JZgJTH6eb5rn/GS/S2Poq4Li3T1Ik3yZVr0c6zqAJTnx8znaUlE7Qm
i5zrjSEcEg7weUyJ3hnU1R3aN3t10T5fV35JoRW7aJvY0Pwx2WJgzmcCOasHAqYU
ahuPxY3nvjp1qOZoujbZQQlFbCKMtpy7LHVpMdfXq6ApI1Z4k3BJwc6CX2zBqLKH
k4aW9l5fBeKQO+IVxaaoTb7AsiLgDan1P9bnfOlfnmiBfpr6/+Yi7vRr932etgOy
ofwPYFAzJQSS3tHN9wGdUeb6ysIayEazNjCJpFcba/yem98ZZYZtWx6uz2BD5lJ2
q3zqNhFgpPsRBZDMt2PwsK9la6/a6JnFvhb4f6sNnNjZFSZYAhfLbsX1WqT4chwu
CSPQKZWiGVPYScx4bVB+aROuciY7NJ6drP21qX0AzDgQqR11jgr1ra4BRRu06KO5
74i8Qd4rEjMunZpIb/7bYLtU5jceuRfJsVkIo3w8L/bzFGtQ7RcMM2A85zQtLjRW
6kjN8QkZN51qA2sP863XFCMTEZSSjSt584GxjSB1yq+c6E5re1OgfKtDEpTjPqnS
feYp+wXvsWXYEincsKnNOhRVuBxNjupsJqhr2ReTca+o1YEmj99jeHGMBujkb3Af
BYl5kaQDwLeKaIASxY4Np0rPIwgY/P+2GlBSLVL4Zya13XnPn8tHeIDemub8eXjT
5LmXEqNmNzUAyzlnn5nEeefVLZOW8qS/nhMy6c3ec0yvjCSM8uWsczdQOw4YYcLb
OObl3L5Da37jChSFNaQSm3QkaCcu5AzFq9INYQ61flMN3f4ai5hmMYQFhCFHr1j4
Bzdm8MoagBFxlXUljMwd0EV55bsRSQlZKBvlvj6ONTwv2BBBDzrqIQLTtLsMMVmk
4sG96CffYBjszJ727uVYB4Pxjw4tpQMjHWCQ8EnkZQRMRilzjzg5dysxIs17U3xO
eYycAL9jan8UTVXDr9d6HyDwYoftrMS3Jv7V/ZSxpyJk8hc1a4+C5xJ09hSpuN2R
sWBAHhJ3SJ1LolXUKtaCjZmM57zItOWxgtMFiw83C4jZkxcSIk3x+XOPhSQYsmLS
MvHnCosuJks0OeUY7z156UY1ni8TAybOqZNP85maIXvJAyuZ4R7unRcT+OVRYjQj
SIO9tqEuIlNAvd6ceSWRDWlqef4/ABkobOB/6NmYtXtfVDvk8gyBTySCIpvLHw7d
WT+iYDCy7818wBER4a/DpvwCRyAiqgfBC4x2bh5ka2yFdhcWKfXvTIYwNg1gCHbZ
gURa/yBYIpwfcPgdjceFw0TioRqzJoeQ41eUUcfCW25wbDP/mSeeGjeTQhfILKZa
VGd33pjWIWhbS/JcchD3YpF3lyy9PcqzpqjPdXKrECSBVOrrczOQut4Yf+zgBYPI
QWiqPCLlt4PE3Fp+yMhAvDHmfADaioBrZ68Kfw23EPrWpYdgihLxgkVFsW7UBdV4
sHhIf91BTgZpq49snt5p/QsxDXbspEHeM3SkwX8xTpRyHIKt2pXvOe3/2sLiCOFz
1JI2P+7JeeqQi3FkyYFkCDNVisSZKr/ciLxgLkonBcIWajTE/oBBxvgZu5TptATn
2MgBq0NTVPpBo69WedavtKQeU2ewKCKNR/XVfpkGXV8jRn0k50CAg0jMNLAwU5HU
EyFjSaEpilv05dql9taazS8CTGARoj0UqpzsenY4gzZ1sLv+5pG6kSnqXqjUyf1d
5MGZfWq3dssUG7fmiqKOymmEq7da0ua53KouCWEmtCb0R7du10A//kA7BEWBehXD
lGa/321eKlgcLRw7nFld+cNSV3zZV0Dya4KYM52wQxoF2066F83Qa5nBHfpPxMeh
bMwvbolnu48MRwsLk6T8xnRe836J8qnHduRi/PQH55ZDD/JH7MWwRObXBwKUHtNP
5xwZ6OrXZQF8P/T7WQm7ULnpMAAAOX3dIGRpGT8s6wPMc+BC8jf7zYH38cLA9LIX
o/Vr/0P2YnFUlQ0sG0OYSOd0+NSQWzqQRzrF32hTroezgla794InKcIuzCRaQfs/
47GklLwPmMPg22fEwhyUw8KbvtKGCwA6SIdEqU9zFnIvcPzzKvoly4Am6e/X+h3M
wI/ste5neRS/rOXxyhhZhNFee1v/TQZ8bXV2nzIF/PE3J5ZjuY4A8SM2JVgjylL4
hdJWg6Jsrt1ZNStu+uxPGZSg2hHFgWovQeySmTuuCocPtQI0lYo2HTiveMwuCV8E
psuwqy29NTIXT/V8cCnHA376GNVs5e4MHdKfKE0ome3/wVPxM7J9wSKVnGiSqqKL
abbH0mwL8+0mxYoOw6pk4pl/PF2yrY9BiTEeskNvgN47ngAPv6cmDwq0rLj9gJED
oZmWpNkm9+2Qq64JBVIgfBBrf7CSN1wlVu5HBYE9DmSZVEY95a4+qkh6C8Q94Em8
JU4VpKnQ8K2eM9igI2mP2BgoL3N2D94CKISmR4vm55iWJ7qfK8pn7qadOm9vxRct
dc3G3/hSMP2+9y/zc1A6a7fQ7hWOTfLVeXc/fNFpEvlLd9FOo9krfYNJLpHQvIiF
NP51u4hcFkVGQGMhTlYZIZPhsBOUthyv1MfGrxBro7A2q6bGBOMLH22eIbhO6TrR
XOj5yDhEL4w22daCRNRF6WrqPHjXn2GainrLCS2Vt8MQsE2Dxzpl5SrXvN62hKLF
MeP8uj/RM6b4DoD1UUl0/gQeJ6Q6Edv5TaTIpCJNiZUl2CEQV2Unr7ei0/DaiVaT
SWZP1gPRSXNU2eglEVbIRwWffpP6VzuOdN+MI5Gf2jWG+cnl4Ts6Gn/cI+YMAZwM
s34+YDgdlMfCe6aCBe6fN6S6tHtZ0/b8CGx28sWrgCerS8RmxWkrOSE/Gs2uX6eH
cuUGs2LQZXN0zNWqWf5Zv+OHL1SvYDahiFFi7gZHc/i/Y4cQ/YArQiP6jJn3LDBu
gsjXrS0xkzgFAbkkOsKFHREVd5mPd/ikXffRf2xsvQsXrW1WsTkIeubK5WXB8JeO
oM11EeSxhjUB0gtyPgdyVwSTAWQACLw2RJpgvUk0k+jE+LweOLCvmjebMJrQ3epr
svl6KmEaSOC9uDZ+mFNi3e05+8klyt40mQ7EdWJ84w1zsXqqj9NehDKlUE9nDYWn
FHdn6koKzzrTRYP2eeU16hK1VBjTHj6ZCVRIERYGdW4ff8bg7YtC8hykPHDMEbEg
Z/VcA7ms5UJH1aBYw0YFkgChQTNjSF3pG+RS0uHuNVkvgf+SlHCy9gQM4blDobTF
99Cp9Oiq/YIXllVAc8CQ1trYcCF2SOjNdJ9wZVtLPav3U9H5CExjRR/W93eF9iaP
/KlsevDanwxVoB0nG7bjFxCSP0/DTX8aaX6SaB56yRZ6P2Gov4UofwiMlbHJJgVu
PNzXe3ozsaZmkYdXO75SNP+4V3jmblSwDykmIiLdnT68WK9QGB3J0i2+mt7hV1zQ
/J1pNbfMGzVwtvGKA5QNFWhlvbqM4VCui1f5l2oGzP7Oh0BO/uI9v3bqAb3tOWOa
CaeMurwOd1jnGia3vYbKlUqwPJbY88pbjC0gFx4hq6Ar+3aFy2R9WNsWWw0GJYWk
V6uayvVfFHSbrVd+cyTOMc+oRz07DI201Tvrl8hIvL1LhGHKlgBsSyk3tEnYR+sw
kJQsbdWC0SNPVFv0KB7Xxo3d0eLtjwPEvqrxx+BJJ7nwRHhpYIxowec9HBsM090N
bTgclmFKSXE34BTGNU4LKOHtz8xRfg+z2iUHIXnJvFFjar43IfixXY0ITrqawmWX
l3hfW8m4bjYBmJnkokPEeCLaCNR01hw3KawAf4Iqo4LbYMrBSBkfLf9icKYgWJtJ
WAw2jVhFg+W5Wxj9MWkNz9UGcBB+TFYYfw+xKAyEj/pumUxuYKQOjf/Syw1d2KpS
M3BWVVKN83ZRdyPYmTjU9SuxUXt9rJHhZXJdZC7qpgZ1Pjld0sFM3dPbssN4vdBZ
vhslySKA8JNAanryurAoCKe50msffAiQrrcB/HcMBeqh0z3sGAAS71RUbbyZvwwP
eAmz/qR1/kx9aDpZiW8KPqY5FBbQfxp1N00nHjYxBZef7yCcn5F9cR45l0HVHA6N
6/HNok59B3JsEJ98J7IX16xr3OTWHu9TkYFoFFcyN7GUlwZCb2e0Qsflx2GaRIX/
nXjtJbUwuqbgUux0stgM7bx2GGEKAaq9gVG1FX55FHfnAiwioPwGxE3t9AZtWqsf
DmNS1TOTDX0gTNwC8zGSZ+9Ij1Sf14QOyREj8vTlbCugR/sSwOWieNfQOn7cquyd
vWRa+TG9LV5yFVWGlN2RdNA8x24jKWogWCHpnoJ0iWK9zAfm72VJee0Kv8or1axR
4q9i5oJvhbDSAISLAA67qHjqdTcKQa5/nR0YXKTUfEFYotewoS0con24zyE9BPcp
362uMUv0wMo3gzkEWIFN/5BSG81vndnhKV/K0WtbgInd7WtrN2S5D0OhEVtt94TS
i8UynE6BUL58uW79orznT7DPABp8Uud/YIAvS4FsqpInrao9pbHoRqgogfsdePXk
FzQF1xYoeChrQDrU/5AE3Ct1nGj1NJqo+D6sRa7HSLNJGNCt6lOnFOOouZz8iDWn
34JH0IGWBcPO0sRz8Tro9ndmP22iUUc1DUvRqb6owlYSLKGehMHWzzNt03ckXoo3
sXyB3SuxAVkaKhKtu/RK86+yu3G1DK17v/Bgv/CdvtJr/kNOXxICRlo4Cf+9AVb3
3HSjjeu1KaMKEf0wqzsoLBpujTXdveY5RqwoAHdi/rZR7hv/0WmqI/9XXlsRFOPJ
HR8x/V9yWGUav6ouHmCcj+/h07tF+ig9YzDOf2gXmDPuIav8gLC6d2x0nrlsdL0T
18F8NiyRKekKdRHzBlo2hpGnFqUeR1r/XlfN/mftfsvTx+X0h/R8DEcqiVh/0yVt
28nWJmGltBfr28A71D8PqQKaonBU/jjuTkgPek8Tfxv5c4cPZzHClDrCoF3DJbZd
IXaxjSsQiD+iCD20CQkBUmOp3ASH+368514OaLY2txU+4sKZ9Zgj2Gw3gAjwom+U
Wd6VXAId+xwQ1o5c9/gto+NM4CTdYwrKCOUGnqLLub5BRRXPyrT4xloan7Ptxe5x
3HW2AWTfOwY2Oa67ub9kXLnAcVayaoWMbn4rRaII0J2HZS7c+56DJry+Nl/P7ThU
gMRn+epR5W/ikeZQOzjbzcMcdQ1Lsaf/917EzsWT6MVgb6n/SBALvC1y7UwSPxug
g3GZPP64/pewPXFnUyBoXur5K2mbj5Y+bXVENKQ34u80F5SsR1Im66RevMg0mEsw
+e/Ln0+G+BkmasdkVumrcF51x/v5hgokZ4Dlwv5XXuV3XfAsdGtxWlscDQd2wyOR
kw+GqlhHgZH919m3onGAIan8K+ajEAwa8zcC3hdgMikGO2tk6pjGO2wJuyDUOlFV
LB+X0YxrIeGG7ZycNHrSGd14aYxYE0oKS7LWBG88wHq0rtahPbVFSyWdhpQdCF/E
r+/OhJTeQB4M6/Tn36hTKnGkIFGUS1gJE1HpjAm/xzbMttglV6lLL4QO8VSkGglH
mbWwi0wzHFGcXq7o7SboJa7LE1BUoPojJMx+P909Ep2Og2cSatihFsM2t6iR6tjc
PoLE6zH8NNj9Xm98aZmDHvXgTh9H8jTAWE7dv0rgKLXa9mgdI525EfMNGXIi8nB9
VpVu3hwXjZDrOBDSkGegyuqvFm85guoMCGbVYkN7HPTIwSlwWxInrvAaTxQ+TTdr
EJmJ+pDvxsNZlyO8L66smM52SJYzz1PIA5yZ+I2enV3jXqASA3bwzcU+ZSXzLToR
JzFSL6/UOexgHS02Np6n5p5ZU2WPPPOiYvHbrejsBv7SJVwLnvk+dtJH/7l/qW5H
bdfa4ZNmbH0ugn4c+QrlVQVhl4L84TZCySQqbQJxF+NQmSUmqRlAH9yE/crO/PQ7
9qifAvWwAdCJEx2kLVXfVctBj5hZNuxKU8NcuM33Z9zKbeQAkd+NI/vIrJchVn1B
d4Iiw2zKwS/oQAnBK6M4ZOgQnXeRxJpaaDIxUgr/SnkeSSXGlHC71GfENa6czkVf
Wr0PD6Yhoksy7k4mMnZ2Ek+noZbKIgyI4OZiUq42B0ffjb9iVNqTrCUcwlRjzw3h
o/AdeNTmC9y9vu22FggR8TnmSpcgMoiQbInh66LrLx5TRNJS7EM9EWXk+0jkT1nQ
GLNOSaQrxozQlnyWWwrkP/SXlXFQD9i9TMMQXmba72JCv9BxclsZUH4sBM2RLIE9
UxwjhXWIBXQMKY2C4Iwm/JdY6BGkerQ/IEDLejs7yDOeJfB8dXqKRCwnYXyXgexq
8Aoe49jx/e3Cqn7p2pA6BabTC7VbEEVcamASZXRhVNHh0azWDpPZaG8n9wLpMkrp
2Sfj2pbJaQH/xY6VT530oZquKS6SbGfwtmz7L30PwJ+Sb98RXOxUKi3ZFmYCs4IX
qmF81SLAUld3bteNDcoZ0uWK8Ff5L1Mn0yb00IQaKhpLTjwdXcw3oNAMk18Z4wRe
l0hpNS4KUB1IiN5Pob1jTma96R3hVfElWC3NznTTOXMHIdvAH3WYzKeh9nyY1yhZ
Qc0kELJBEOSyj1ZOya63ksQlQK+u78I9l6i0BbgERanHjdwHX9EXAO8inKcSh+pz
grWAOqGsURHDn+lcBx9HeiL7GkvoAVap0IYqcgN8hLl595n0MgbQIDVWYSphbf+2
XtTL0Lv6E6ZmWwhwdcUrcAXpVrnFEN1kJdpp4xOCIusRIa9sIv0WtLI0LSoJkVai
X+rSCTgnmBbGDZOTnafgBvNPEDbQtSBE4Fv4b+VwRxD1Pev1cyhrHdcawXwLD93R
E9s7H/4v6FiHln853WcJ4E+f6JzmyX/x0jiVtSz71g5fEZS3Pj9opfbeqF1+/rfe
NruAioiduFW5fALygosgvXS5ISOBSAmyCReOpdHKWUjtagtDmrDrlHKszEqq9xmq
lv5N12N3IhxAfJbsAHjeLgOIpgFfsLsaRCE3fFmHCyeBmkAlIR7uM/elGtjwWNFf
im7bqiD5Q++7jurDqEUscVvWF3jv4CMceS+G76VxX4EtwlPHIWvhlStaCHRHtww3
tGWf0nmiWrYjzmaIi+8V/Hg3YizyQCspxAXCVEQQyQeRgY3Lwm/hubnUHhZEvhGJ
j8GsEG9a9Pmv3JyTezWOZzfvrUfge8ZrjeAn5ykvdVWF4Z+PRYQa1NNfxoCBNZBz
8E5e9C1V96V6RBshEFzB9637ag/6+2htwUhOH1e+CUppRN10aTQnHdCTb8nGnF2L
diq/yFDzpzPomymaH9R0KJ4oYqIHFfCzGTA7kXBG9UMW5YnssV+EKZZdDqxtuAGW
SM8wcfOIeIKHUQd3atkynSAf99ODVD24XFOnFLYIOM3tf64mlzlbQtheKH1ZQxxh
0tQcnuIYzjwIsC2SAXCC9T92vltkAHtOUwBofhRriROdYPU4hMsVpfwjlvradIUE
c47xGhTNlJ/k4Ne11ZbC4w6oJVNThaAY0DTfyvNXxX+gwQIswoZJpWUcrD2a5qX2
/vfJhihDm4wuexgEoHww87LYww3nHs62hdILn3yGYYYaRKf6LPjUwh0XVcvYZNx1
QsQFWtyiLX1xlMK5bYXNovhPzVq3CNA2lVw1IMGitIPT6TJDQi8II0aJqxt6K17B
N+HBdH4cWfg1se4ZkhMOUUR2/5T0Wf0U3zKYfGZHFG+TSQVUrG+pNAtn5LYRfn0n
9K9K1gWGtpXuwTUdaOsEh51OC7IhvYu9MPDhwTI5aFDO+GoFs4VT2ePVtgQVQSsr
FKvNpVq2KEAKnQff005ZZLzT5JbUcGCKQVq+y2Hf9td7OM52TMQ9LUxXmJJCwPs4
sb7zqFfImbbyWLvEu/hKM3zHhNqeTRyu5TPlv2yz5+IUbx52siZ4jW3QPK8MbSoY
S6y+bd6zKZIurNEDDEp0ilwJam9a9qCaTBbLDR21QtsGx905t/IDfoERzGQRgJ8P
AOehN6T9yTHokaAUsrgYmqKmsb+sL/hhd4wGuuZKyNaHq6aohGuIzsDp4a3GVhyb
+KSK53o2HoUkyiJMEA9boHmYRV2T3BCmmCn7M0xmrM8iq3n6Roi0wUogN4cObdhe
vEfzIBTAuCKaC5nAd3RRmAsqyGIiXRMAio10Aiowo1n1FxZ1VWQ0cOn1MH5Hu4sQ
b6TESuSgAybr7tiKHnI63YZRW7zbsjDMsnVZwzoURl0rmuXyRxwZE2UKCtT1QqzB
40F9IC8lAwyXOBWdvqcjV/LN7lB2t//XboDw3m17CEidzFTeCzFs0XCQlDymnphv
uxRHQZKlqBFZy7T9tLYhHqDUXJNXtU5hPhW/pd3X9J8D9RWln6tTKzhCCtJS2xSl
HO8av5NlaZHdS9h7RjwUSDr4QsasBtIliee29y3MxmHXBbcVXAr8Iz2uF2BTA+1T
fSxL2nRfsZGzJOAmtRdvOMaF4oulwlfLXLEuQxYGRCX+7dbZEsuc/5v/s88oGqWf
uHd0dpZL7HqMP2ylXpWwTT2ZQm5wOiQrpuXIFIRhX/6yk2c+L+UsY4M+WDpjurZT
zhlsIWPcj4yQHnoptFM0dx+1lX3YglnwkszvpEyy+KcBXFwGBoAJmd9hY2yCRYwb
fdfL8DgcfNgBe5Ydo2wMlLHlI6Be64jHuFXQCwLxC41Rl9bZWCnpOn0lahRu0BuO
GT7aur4CJCWkJqyHT6J3vPvU77Lj24+I8Iz8hMhDFZTGtiZa23qLNmt9uVx36TkG
iHeH8e97xwjWe3zoAzkML3blc04mdIkbUK1CXMHVlUIH+7yvPHWNMwmA9buHMnoo
EF7D8x5h8lQ+vWBDQfKaKptk60SKrMfIWdnAUAfMyvOgBtMB/Ei+Is72vuGM1t3p
PVtvD7ZxViSYw5obP4LBKORzllfab9PpaXGpLkw11ipt/wxXRBI7ZAGIOdXjqg2e
O2Z8ihjc0K3Yt++TvahVsMQkuQbCF7EmcC/cQlwOOs5wnq66GvwPMVIwF4hYLjUP
WNYl0IJeNRN/oWeNVkuGhd2loFFTz+/ydzIOOfUj9UNB5kt+fZuub3gDVmOB3WTW
3PrKQ+c/egS8rGUs3n3oFMfnRbSX/ss+07W2brRcBA18L2P8j9W3mwjg4hxfzLX7
z0LLzJbqs8buXzhiE0zCgZZt3VbpBSAyjskBxcaE5YUiH4X8+O4K6aEvdttH/Ask
vM7lAgcUNLhm6r5rddjWR/Vv3i7k5fzCOEtiguhRH97Ts+vx1LaECpuTUQydNowp
PtXGPHRU3O1gunOT0CjRKctn7EcA27W8SqS483zWr3KVMnO7RRdWCYw4bDB6xtN/
XY/edpMD78Kroh9UMAGMzNkOwdxp5RLbbcAzYSeCqC7Y4g9XkAZpSaGQCP16Z/4S
Kk/ZDo1tq9Qi682z9sJK3tH8+dbdfomuc0uyyFpvWJm+/CDPT/nLEAM3+/W5UDPc
5A7XAn5aoghB/wGdbDkcydmYkaTa1ZH6eDHyYSTYrXnhzPjH3gAYI5AFjHmjnhtG
BZifR3McnnHheqtSpsmSxF5liyhuyKnFSRPGE+eB4NcuIMUAoEjc5ozr7Rg4PIBm
Gndaam0Juaee8RfNhEYfmzt5S7VE4kqb+cRAYpYISjbjGJIJRFKSiBuMEnOVYMQB
d9bQfZT4BBH5ValpbPYYbTszsDiEmiQNH0ZFbIu35J/wHMwLArUktJyiw9zigISj
camjKsX28jwqfCH31m3NYH9j99PZvVQB2TPft5ZHyPHMH6MAxkhZYq2szx8cSHz3
tgMWBdBu6NCVlcPpmzyTU/eCIsdRPGgMp/UtoX/+/kHRXSfvbT1YETVWubyc3Akq
1CnDVmKYEGT3iBkjljjGG2sMVyxOuHtxnzeZbo5cl4RTpcCVj2FQ4BsCHUSBnspe
Rg4nK0nHwEVFaMQ8UVLaNc4f5/8zvfpeH4tReJPxmiVLY7uKJFxdP+IKps2R8xL6
Yqw6/HoKR+ySIwrv0Zm6/MAy2AuGLrMe38xVeuRrMbEH7vmqGGZ48nEGNFzxVPp+
Aswt1ssikbhhp7MMhcxJ4MP1P8G+XBez2C0r35OryckuL1PQZvqiev4sEFssvgEs
4PF3iZvAMaMqNDm2JCV7ctaTt0T3w8SOwogUXjS/0B2L4VhGgYeo67Y97ev04cLu
OledaABdxWvpFRGswHqh2mx0X1xJ8/l0sZxPEkNtLjvhwKPakawLLd3ZeXzhmdqL
GjzgmyVv432ml/tLy7+TRSBwuMfR9huaOS/y19LupchQudyCvWFCaPNQGVTH2pvV
3gEK8rFtgednsNCNWuq0r0WOVgxyjK6CoEXKAbkk5a4/bIxz1ygC4GJO/d0i810r
+DOHgNOwyl64DV0oz0sJf9wUTh0j1PscPYv2UQFa2trGV/yhPHbaBBIS4/OTGkqS
seV02wq+Q9AwcPX8ovjK3ggh/t2i8nc+ruZdzg8B+EvIIskmT0yPyOf3Bs5VE6CG
McPSDtcKpHy24QYSJCO4H++e7DOyg0zXzczs/n/pAfn6k/zSyaZuN39kXQxUyHea
F8fXampHpmq95AUYADypJLDLchkA5A/Z9K/iKf1zNDudTCoBDk+wyFuxDlYLA/np
EgcjElSeX61HBlGAQyZxP/WOh1rvG+nxyrT3EmhRC0fnlqj8Y/wSRS2K4tu1wbT1
7OEAlKHaYZNp/aP6x/acR6+HxwzePDOJTcV5in/CpUb25A1kd+tgmlb6U+0VfgoI
gROwYsW/5x4oPafeF16lKJVJYr/m2Mh0R27OctGOfR6F0qOTt6S/wLXMRxHJDjc2
MlARz7S8JsJTbZh64O2FUGbT5s9NRs3MjDkYd2WqSeLCspSaXY6dce4QjNJUHJnw
57qg7YnugS1W97oSqoFKgYS4XY//Oaiu26iNIEYkqm210ebPUyBRFAblsRvn2xJj
XQbqJrrC+yymoNq46wHI1DykO6kcZW3jBth1ZPp5ZSQNODYLqL79s35i1dX7gSFc
YJPkZGv85MsdrgQJzuAkr1yAWNHvxQH5B2RFHpd7V/YXDCkOffO/jee3nETYnxUZ
6xzRgHlyUIB7Xm6vnnsu36dg3GOhGw57wy+tHBB2Zml9/jutlq6YkhHx7+fNioGF
FTFqEzL/mYd743i3HTankNHYgt6VgYA5IYBnWfc7z1fg0vpTDhJRGt994T4uHXlQ
ChROsDpCFB73Klb39EmohjaFeBnOwf4rbgFbAKcXFM2Ur1oM9ihIxFa7eIOP8AdT
GXDc2cJaQjBkIVT06nzvgerapl2rq6mhY+PySNgqOhXASggLWVxWusVKzOXIzgwJ
4QSK+vXoEBtpBuBdgM8D8T3tAAd69taw21Q+kknoLmFOKrW4qBO5+qLLra4j6BZd
TQ0JI+FEb/GEYg/qRXFG8z9GMQxz6scC1LNtkasElsEKglmKAarIvIzx8BM/z6uw
7c+dn5OeD8rpGKBk9nUheUj8DhJcradau8CzSD31e9zjtIUFk64zM5YISL6MaSmi
K6tlm5nL7qFZsVBW72HICvLfzMhqgF64b4dayvo53+YY5vochuaVCSCeBJpUmIRK
tgf+30ehKCA6Bt6VVyL+84KgshDALLMQYF2H4nQxcWIqwD0Yg459QSa8peNEcyBo
/jzLqYtKp//4ij3krtlwiPtjWOv7uwjP8DtmZEVh/fuY217CFOjcvWCS6rzjvObS
vKQ6bFM/n5pbIRkHHsT8no6MA80uR8CEyVF/kMreW3g4jYUHKynRApOE/lDbm7BI
CpCAhf+P7yQgpZ2bih7Hrxi9wSeaXxQQ67oIyKcG1o/SJLF/ysLhiRSrYjmCg8C8
wmG6EN5FvJHn+ZpeD29x9MmkKUJFT/A7pxC4OxVA+8qSgr4lXrqiWv1uSJkiKfIp
x/DUslDxTxcsb5pZp+OJZJEA2gtq3IWuXzqP7/ljsNODnxiPgoL+l7RyOo+1ZOyM
r5fBR7PgDwYIo005UiURM8vvXAOC4Zch8FUmly72TXAqPF1tOUroUlIZcckuzL1M
1XcWQUhgo4kB0SGR8xFQ8aQnOl+h8+BqWC9aa+yttpUDP2l1kqHXFA0ft8q6A9bO
DP8Y6pcDxmIrFnY0mwoIEdM+aadQk+oTEf4vt8+Lp6GAFWpn3hyvdPyt+2VW2grN
7VIMieQ7j7oFMeI1v2W5yr4N7plvrhMCQ8JyindUXU6JHkWt2dlX7jqW5koryIBQ
TsXlbVpxZJbRYyFLqX2PbH2PuCLj5pBsWGC/vXsDMikVpHO/8LkPm1MN2zMqy9Rs
JT2rO/QY5eJd6KW7inchmB5p7J3QpLrf7hQ6QofygFRJmAXjl9VpeUDp+QbX8YoQ
cx2o9kq8TO7wF5/vjoSaTzvtK9y/G22vBWotNepiUj0xUAdk2/uGCw8k7OkRyOuH
dsoiZu0KLEXQr0wUYglstvoVMqiv8zt4pPL31/qd0X2JLc7Y/79LZH15flaYz/UE
GcJUpNplne5lGm8rnKGgRAbLGf7nCKbfOqIT3DurQ8MyAjc6dUfkxBTj3Xp9L6bw
MEbSQHzL7g6BDAUuVfUOtOOqhjtp//qCIQYUAPPl0fb3YosopTbS4TFsO1lsdbzC
K3kzdVwuCMKBIlZ/GD6KYCqh5a4avNo/FQvZ5zYdq1dCG4ctuX2d1gBtWLHb4Dps
qBSEAdvra4oKTvlz3jQzi6ga5/j1yVEv9OA36e3nQjvfChs4iQYSaVe9205JHdkQ
gVGV+EE4OH/0y16c+dHC0AC0C7A2x6HqMGUcCa7aO9m0qZAfXAOjfZgLN8YPBKFT
9OJxixceAkHDB4tmoVJLseQytiKX7SzpCVuy8H1c6DcrsQk3n75tuYeyYL+820/5
OHIDTSim5f5kxo7TmaBTOUEuTpGP1BGneJLYsmAxMO2mDs/HXSQURRlx/1E6HjdM
tL8Jus+Lqbo7XWycVT56cRyy/D2ATH4nV6Xb1SKYfu2cZVVKH0lIrxOFiCUkOhIq
hB8JN2hRN/JDi2cas5T4l48XgdvwK1et/VMU1L8l6yQK8A1Glk2PwTtCtY22W+YG
uZVu0fp3Yw7/su5ozuu85lL6Ug943znJT8K0kez1cT5o1o1W4mOoLbxO5rSCHA6R
kr5QdqWxAydGflQn2wXA5qtFyl/0XRppFZPl2vlqAHW4h+T2QbLmDnSM04tMbsZB
+6j72Bz3DSfUWGSOxs+Ix+yTX8PVws1eEA6suz0j0JFCyHEEKc4dKlHFr1SdoPtn
MiaID4gy5tKWLB+Mc0xcaJf6FdrjTvp5LCT8h9K6kYkXt4E8kDmzIkg03Wm/akMt
bmRA3LCsDCKVOjAoKrm63bM0SEqwvy65NWjRAIPS5YXEyg2Pvi+xYqdSOsZpOlDS
gEZ0GXaiNtwc+7dh2c3RlCM/EoggLHQsqUZOwLz/ebSw+L8KoHbeKic2jR2ct08H
oOVoHLpTZeeUWSOlFuNyjGnnfzCHlKkCPxQ+ls8wQOqouKRRitRg5UUiZEi4wRCX
7CbiC16sKiJwDUqsUd1CPJoOv80vCl/gogkrSHS8S2H+HaKgteQTptWOXe4VbU7N
p0alsr25y5JVjZYKXKY0dX7V0XgKXCFt6qRBZdGbWZpTICtDG+e6ccREvXuOHzIe
uLYli83ZtPHo6yxMVDUVlOglmhi91qOqRFOVK9xeTPkIdb+qkrFmujJEiinVeExT
L0g7s5YVANXlrBL2R+nKnAuqP8RIo4Kf9KSLa8WO46j9lPL4Mt0oICAJEuvVtYFU
8a0LEk6ecllFuD5HMbGCL50yeLa4V4G7LYIr5C9ExajyGmINia2dOD5viT3hFagm
KRDAKu9tAJDmTAfw7VOPlD6lthwQbFOzwnFtf03ephdz7qcrbm5bLSculgtyuy0j
1UeW3par3afQo7hf9NIsFC4HjcUnybAcVgYORCEDwAoDCj9TCC50Qj9GAr33x7N3
zLxZNl5KSghB9HDBgyAPHFvAqED+dySt/9s/kfWju4FzOW7SG4ME/9ocBjeCHrBs
L1Pd/IVJ5Cwmb+BzjgG/Uq2Nc+U2Sc7kwwNfz+pIdEat0dlhymOTnbBBTzvZtFxX
Qp1hpfZzIiIJgZtS/653a2swHXfTK6fHtf4ISSYzyjd5UGfzGmmQdasRL0eMUKY/
nKEwrf79hPndh1cXmhQee2IngaLV0u/imlr35LuQpRd/SHCwGeRR+jsAK+RldhCg
Q43EIicaoGwJVSTgnw1C8DDpI/kcGwi2t+1qaNHO2SgpYMpMHtQ0SqVaMo9p7Ho7
03h0fWqB8nz9UAnb4RSYEkuH/9UGX1sQfIz1Hw7zSw/m/saiaUgfFLCJQfE2PdL6
94+5mHoZoTYV8yyQu0tGUzls218I4InQrV56VTZTD03ogfqqPK8rlhEnyGMCPz3O
Hp0urae+VCug5dvVVPanObJ30+8BAR5Zr7c8jMXP0Wozfcgcv3cZ8bhppLlF3Ect
8yixAIuennRiKz9kWEIl1s+1/Ego+bQIFrJBiFuUKZFgvTxsc9Z5g5TgSmZQWDQy
OuPX63uRfAv3JbPRQnLTi3DcxZKfxz28Zup2B97Qa+46riPDi5rbxZhAr6OF/518
PwPqxkJOUmQuTYr+8yb4XksAs0ACWrAOWOMIwPXIUTdUGi4oUBvfrzkrnqCgyIBq
KDTyPaKqt7mwgsCf32SNjuPFMQJKh72vM6TZf8vfteZ4qDc6ialBcuiPA8y2uofm
T2V1PtzQaLI88OshPLKQMbVAB94uaU7JlXJS910ZCHyC/M2DNF3DSfzzZdg33Luo
A2las1bjk3grm2I7hRQh/qFn+EpzDdOK3gb6mXyV3IMe7wm7+G9U+JibHKWttDHY
NB4OoBVx7xWuvoqPYk7ugiok5Hb9Q4IBRRhjcH1NViCQP9t/zH0oleoolLTRtD8v
QC4EmbOYKya+iRNE6V4gMGcharn6vnA9Gg4QZmXBsPiC0FeNZVcqh70cEd7WTu2S
4KlB122nlmKzPX7LnijAoHg2ao1/KGbQlTupRW4N2OtkqEI+AfVKWgFE7PGU+5O3
zWLRF8o2VTd0W1Jzq0NS+t9bjs/05p7MfXShFCiMEdwpAxiNBULhBA7tgmHAPJ2K
+ZK71681J0xdToMZSjL8kIzBECqM3BCSGrKOi7Likc0NXHZCezyc0DCLuGKjJuTd
u/vQ9FpJjHYHNWsrJm944+LuHQY/fwgClOl5jlCSokdzcRWrSVNfvUr00gBlrDfM
dk/KqPi6gHOUs99zpWPICYtDjP590HwZqluVP7+ez3NYSFrYv09RuUIOopxfJv9I
eeSwG1BgXcBF4Ch4+ILbDDDucStXWzB+I/X/i9Z3dTAwRdLJYQwURvvqwwKx9EUj
TOrjywy4/EHaa+M/Y9+UvGmEa08lmO42fNftF4GErJOTOL57ECNtDbx/SndY5pXM
o+UznQX3mosJNFiAmIICl4RMijskb1COmjiqZEBJC6sqLW+9znjx3po1QqSAfHH5
sW6Csz5plSUaLP+Nxbt2fMwpeuT6R9P12kfloiQg6mF5dbb9R6BK9oCLHqSqfzyt
FE+QOb9HI/vXiDrwnAh6GVr5MnSXCGhgO0MbM8z9HnHc13vQQviYIGjc3l6lRyuy
ZxWOcsopiS4FpZzbgObgw1mOnEm9p8biK3VlJ1B1rcvim/c9GbrjQWXd26W+SMeJ
7GV3c5O88zWGiEOQfAyKJD1qfx8hwNnKJAF4qq+VTkSkHlwSqX3bsdzGjtgLd77g
yIsTVo3/h+BlmQRDCCESrAeep+1XhMYDSUEz9yzH5eSyDi8zyQRIWxbCQh/C0Aou
UlkSUuU/8leZ6bPrnTusgzEP+JV0Pz8XpK/Tf/K/GpPg97lO9dXXGFkgPpnnGFwo
6ScOc8uajfCHdlIxIZVn2AAiGNBgrKZEq0xVRoOXYT1xNAb5xUfUDwsC0Mi5NuaE
Jz+VipDS9rz2qJ/OOwxfPaSVswL0UJP7SHciNEgi2iz8NLMzclu14izSfUHfxWoX
aRn+oerWsp8dmQmmSDE+eRXK6a1ZpBNwow67QDXDNpe83EADS/3S4/ztoeiJw1JR
XZyENm43kIXK6Rye7WXXm8D19kLqOaPEWOlCkFxAbJ5KiFTf79Xm+EsiKVcDDKJa
gMnRcKCGkiK9TRfWMkJxNfQxtTmv05GU5zG5E1xPaaqaiRmCDeFFQ5hvSewnbDM5
HQIRd9iWF4sPciQopqOFyz4IK+sb7MMAikDTmwONkaHp3Hj62uwUKsjlc1QyG72R
OFDhEY53tk4lXin+en3sw+90ca7SAE5u0gidLmC4PLMWz0zTVpN6jQC4LbDxdovo
haTdfvmHPd/+sBc67SS5QpA9F5E3HpCN9KvSflIe3CzgkIPjwUfd2yI6N515QsbO
a3GKsvApkLweEdxNla2jr5e8pIg3yy1ckYuCthTVC485Bn/6Pb8qaiQHKLkmeHKI
w0xp6an5LSa3HN3yCvJSX/0M8lZHJy2kvJ6yJGDsH0ZHAqqFuj7v27087nx4WEU3
day2uCGUISqrfA3MvD2HZos8FsqNMiQu2KSY3CQ29KR9y1CjOTG8Av9eJm8+Atv9
yaB5/3zRqpJAY6hGqU2nbMnfMBUFsbRxYLL2YENPlqWH8cLGSyHeLi6eln1yi8Yr
qoilLtHg3glnzoEewoJUfiTIFNUNk45VskjTJuPNRBd/MlI6ysb4QQeWnfGBCFwr
pQxXAq24gNCVJozCGhvGq/owKDpa3+eLrLHBJoKrZVwBDshtUTR9IBP0c+pFOSqb
fL5+fM7rtrelPyix3eMiZ/j3oYOO1fXG/8NdTbDVFtFkGVZWseOo72K81tK4fSja
2ehVpFxe5nIL3U5WO4dTXVnO4nQL0v5zPuDsymbSlgjyvm91hQu1ydb9D7LDkSn0
9s99ixZCWefWsIQz0z6BNmjjag3V+hJo5IlYH5jf0UiK+ykXehBIsEg3rmnZnodK
OCwdkccIC0K2f/++O4bYtjWQn8r/WmLwih8SWopzxW9YdiSVyZR27xy0Gq9HeU4j
e26JiUDSUAn/9qsqeIxrR7IMZOflV64WN9uNjQ4HD9VPJfWA/zTgRNa+FrnAeqZS
0rjXTSfPqpvhYksi/Q7xlzF4TABpPOvEnczYZwFgeDMO92MeR/k88lMZJCWal7fx
ma+tDDN1P+I1sVV14tWtvqVlhM3ykLdk6c1L4COZatjLRnLgte+l9ThiryTW12Id
n1JRthw9Su90/3Tm3iDkExhvy0/7b5I4f3AeZeYGBro46RqPOMJ1nhcBHa9Ao62x
0N7QoBaqvXlRGezJNkI1IU/Pewsd3qmkJJsFFjSzToBBRF5MqUk27aOWfX/IkeYR
4B5zdcwLzmqFWZIE4W2IyAb6KThnYC+yrfZraxTcaQbtCQLTiglszTWbBcp+FW2H
wJmuwymeT8Sk1BheXHGl7RW/FsBCu5sTLcqydKV3t+4Z8GnszVwvjxHA9miQO07M
hRxNUKaVtx02gb6LEDiSPUe1trtE+Jpq1d3kbCkgkyRpLdi5+caemqEpdKRNzWov
eJ45MTn9ArnEoheZYpv0S5vGPTyKVWPyGmNohVqJoMSmOUpAKJPaUwarr7u8OqhQ
bm+l/oU7mE/mDrUv0CVuZR+D0qucDB/LTTl039J3eJeDt/tmXcenOIWo5Qr8Kdet
cXVLeyBWzzM+GplXuFcMvrsaHDOi6HHVAWMyEk0SbUb5ZONNL1I/dyxn40dAj1hE
gmqRSXRbn0SxQm6yj2hYRl2tOArkyHO0aB49RkGe99P0z9YgU+4oWSqlMNX77oK7
WxDpYg3LL23KL9gSA/sllJ0lhuLe2cZr2vwMuv+VvFItblzWAyEsrSPGimNxeZY2
VmBer7x/0pdQjTLnqaOEQ0i8U/uhJOGfqSyrpugrHUIUIN6AMh0YxWZjF/CEUOQW
h8wrcVB4jOHOc9H1ZS/nHDcbPO3Wbu8Ec6TYBYxbMb9KWlsV537jLTdI/aXMorr/
6EyIO9hVza2mMjKZKFMeTObwotEASpVqwMImeWeJjkUxYXPKLAXeV7LLwuLjtqrJ
MZjl4VxcV4rEbn54ry6yNJwN9Pr8l6n3hIH3265BFxfFkJ+qcHGqLq+sQkgThCW/
AJPOWtWRHhGwGUoujx7Ded8tdzpOWzQcxLVgfksfgqR2UmaXW3S4gyV5niWVT5BB
BfGPQnu7PgeVxlgvfjTc+SjdmV/OzQUj3Zexm14p4zKymI5gitqx4/R8hZcrNMU+
nkAURcqUtRJHgYvXgoz5F1nMKSj6WPAXHMG8OSdTj5wi3OF2O3H4A3SsXgDM8+pk
F/qt5hsGgWiVYcV5cXkmRv3ubRRcuM+m2RELqVJGRimMWgb7vXey8efRJLzME+Y0
uWA1INS+DoZYFleQIjE0jb19y+1Ustqj1RN2b6+EQs169T2Aoa9PSv64yMrPanCK
bp2jAJHhPlxsJ/lOCOZNoRC71ktyO87g6A+OJskBYs7nSaRVPLz7O5X5moBpJoMS
3HgqW0uupZ0/7wAeJN5I2BkzcF5B+qpSuZD9wo+CJS3rfxgtUpfppGjfpoc+bKSz
XTChT/dRiEI14oBv6tVFcY9x73hKR4VdvJEzjh9MFUCBKiUYyCfyHijhsNCmo9WH
99sVw6hBVcb+vWxG+dL817b/s67UkcByPVeKcdSXgEXpZGEIZKgKlrggJlHYp9Kr
JMSgGjyEEN7/R8xHCpH8CAY2RLe0aMy622nOi1hsp9yyq4YlKgersHHndA7f1iKx
EFjo9wTPrT1Ift5q7nJPnxcSVH0+hf76joyBxvs9d3ssDPBHkc+n/Q7oImhZRGsg
NzY5zzmqpH3GnenZlh6lnRjl0vv9nGRYgkwc5TQzufAZWeRnVlCOtAYE20ZWSsLA
ApGq9IPoZ0dRiVSvC8WVr8w0CVRWXdoLCoD8Wz4E/uGdS+nx4Hkzfq9GCBzSZjqt
OY0Qiqn/Dmm8gSvKDbhqijtZQB4TrkStk4iVLXmQW82/KRXruSXQNWiTbZbOSSdJ
SILmPUIqw2Wfa42u5N6MYOx067mzRaG7zES0du8kMpgnOSJl3ehhoWfR32plzOog
AmXH7vX0PHwFcms2W2ETgkQ5uk6UPA6R2pS3qygwEfiDvVDI9dfOO/p4EPlRm1n5
4wakgfnff0eaMTrrzNf5N9dOzvj0/hSjKGRT3kQ3sNwKGDq83kp6SFU19tysX3Vg
cYVmfmEkEzWomDl9z4GDr44wrYFFHb9A/8LrZmkPVBNQX7B5Avg5hDnR2WdsGQ0A
moELSY2G/EJSHOGpBSZ8rJgqAl/ejK3OH6PHAaxzSu1jiWjsU1/cPkFFuUywzO7/
ElUBCz6+IxJCotzY/xW3y/hBCmFnLdeJV75JcG3hbCwNGC/zr1DpysrwCM61FV9K
VwGVnJk+i2gapCr08LZB5jvmXb82Uqj4eqVSNt8KLtjCVigiN6HLWlscjW9kZQau
XcEllGJKyoByqqnhm14eE0UGH8jfjWQ/qOXtFOaxXVJ6qSleVAKzePmzKjvIZYxo
6jwyr1ZF9NYBkSo5hZVH5vmp8QthV5QQ4sqIWq+zEGMKRKsvy+qfTOtXrQwsUdLz
6bK0Uj0QVytRtSReu7jWfvGlKT3IMw9rau9RRcjves0AmiWESraQMJEiRNOEWhIc
aYPg1osgpiW1fCfrkmZoI8bVBOnej2+obMDuDpYJ35DzQD022UpOwlONAgra79Ir
POR56OOihyb5V/jJInFCbSXfV/jpfBEUvQ9tg6+dSxUPv3PzsBYUVdm3Oi5pr/RN
M8k3Hhf8nH5NZWnlW98ph+RTdi1S6d8Y4V4nZxFwIDvd6jzLY4sF01A4sbFVB5gB
K6qhZcJHVNseSpEyEdfCCfCNm86tdi9eL8X9AWNvJP/xo4Pj+eBP21oPqFhDGbZt
6hZpdgKEH0LBcBJs8QcCAvurg4zbmpVCUDyoszxsF19633/OirccsOgEepGKOlIz
gWTfeme68UrmNN6HYz7qbfo2F9yhy5AyUydlkJ/fhZU+Rl2ZSFu15tDPsg1VMuHB
azvz0ttIkf9SRcVnjaSrz46uh4oL24+ByTUVqZ3JYevnKCZ4G0Aa28P2fpm4Qgb1
FQzg6AeR7RMZaNAuaUCWl5itGEWU7KuQuv0l8Rr3Tqu/o5YOan5gFG3oR5AYFaW+
VTa8BpWR1G7OXJpwaIk1tpop7ABXqbwrZ5PhhMdwdFtbPKcZ3znA7V6YQ1MsYMEn
akUuCpUxtNDWWXcoJyKmbaIjgBoGN5LvfuKo8bGmIto6VcW2MquoYOU5EuxNLnss
J/QF+SJm+St1/fJan3qnkj78QgHPRrl0s6gC682fRwv6BzqJxBrkm13UoCaPfceD
C6WIi15eIHZc7LSxWkJ+gjovQQvy0ZZg/zH32admzuZ7N3NX40SC6m9ALaBCN14n
jbLmYvwMWAO54og0HPL5fzq/K2qw/AAnHk6mxoo8FLHdufAHOwzt9kHElRk0GuHA
WNHdTWn2wtYfRWd1VzvY6QdQVhV2onKVnEQsu6GdUy2ub0ZxWKC6SUMlbNknvjni
FUqJ38JF4BqqsTGTx6LziXCM+llSmvDgXuTzSabB2Nq+FPCYdKJbw77M7ha8AJt5
nQjgAtiN2ijJH+HLo3rCXwX0vZnewuvItwDRf9MxFzRtsywvfw4hQxdhQklj1awr
27umSUI/4sLTqDPg3jVuKWqxkkC/CelQ2UH2Lk8nCkQmfC5TRDJ7svqUW/oCZ9Rk
bV8DUSZr+NPyloCVzsfQZ0Qigztu75SUX7ChsptpwrILiz+0hZK+dP++yLTfhOuE
vdI6dcByG2Lc3EjxgWg0ZYD9MyxU/zU489YzPMP0omP+H76TVQQIEIZmzaUAotu7
t+1r6YfmoFlrF2hxbi+idZ0/MVHJReC4g01hyNmKcGIWgVyhSnTPZj+uJlJUACX5
nLein3Dck/3eitHzsC3TAdgEX4+At7ccX23800OTXXaRY58e7iyrYOvVES4dT2XU
ce+CWgoObaqmhLaQOUhMGkJUHTcW8zfpK+A7Tplbvxh3c/+Y3fX4fREXhkGHRTGx
tZ+v7pMNUDWSoNKuDKcI0FE3BgO2XehuKY2ZwO+ffPF0d7tpu5bHAAJGtpIrR1EZ
SQ6K6Q3nMvHJVX6/H2aCxGBQSeGU7SIatU6SanlhtodBRkeXFms1sxXJ+nWgPXI0
rCcDZ04OlpM4sEE4ghITKeI6u+NSwRA4DZAqZ2d4BKjpfAbGcd2TO/gYYrNiQ/da
ckULzj08jvH58aYigfs0+ZpfnJ4rYH/K0dVhIYCjOW7Zuyl3VGtXDUO0nj3ehMDp
MF+jCKUc7odUd1UXMfj+L0Qy+RVHBaR3eLsFxua0mF8vR3Sw5r7fZGv/177FfV1r
hhNoCcpUPkEMrvpDdgdp1qi3kC0+FH0qrMrKTZ7SZAON+R78e46Czv3ccpnIctYi
9ohyVOLYzeiibKsLAwpWK4X+/bX1+z+PPrL8Sy6SyZP5PDyU72zrniXRZgdyCqfq
8f+djCzjkmobPIpnLtFPkfa7l2i8Pkr0DRT6baRBQa/eWUOmCDhcpKLjAt5olaNK
WEX5tFA3MjBmI0sRMSHCld7OehLpxTWdtrX2BvbWww2SB9sqwUE4S2HaQFZHos7k
KplZMGaRsWRGjBehEqZEkrke1Al70zQ9qEPsRQgtABAXW1fHkeUd4vqVzqIrCNo8
ktyzkcQxAMVCBlSGL5+sIk60NMdnBAgPfDCN8qMBnvQLE8mUQW7ZDd4V46MuJm4I
AqvYTwYH8EBuGr6KIEhMJua0yJ1fagooOt1Pgp1WFLyQeZT6Deap9Y3/7VVLC8Yu
ITqbDz20IDlP05ik5T2vQi8Z0Unl14Env08gzf5hyJ7Z1thS2MB4zDamkloaLQ2O
OgkYwiydFgGw4c+iM5YeGKOwiWQZZ8cyh7N2YAPt6Gp9mv4EU7KpmRo5z8AlOVtA
1aROpjhRDqaV78Rjb5aXA6IfAb2ruR6MC7QBJybL2S11+DhbpnfSwmEDzS33Nc70
iK0Xlzv/5OnKKTGsM8x82XP+qu3JWGhoGLXSPkIWXkJN/g05fy44eVJRMNk7Ma6u
o6HVJIqS11keuGHPMaFwN3m2lhrUKBzI1qowwqg1zYlx/vxi8GPpOD+HgSAWdfnN
XU/s6s6XJ+3QtdNc/JBIUZ86y2YheMdRL2qwCWRz3Dx/z5veaQk8A+Dw9AQyNOQ1
XOha9YDrga5y2efo6ZeeP0IBjT7CRPTAvvJ/o9dl1OxLBxpPnmlujbYRh+I46whq
rpyZkbDeNLV/n5ay5yhVfp4jPmvKP7pkD+XrkzoOEXT99KP22g3r9PQQgD8jvENI
spSDg+xSQ6vH5fxIZ6oO16enBXgv9lzlyxBf3GEkMg831r9mxeMM+nj+oDmri+UD
arwqNcOdMHidXjtGXZ7WZr65CIcEGVJxQGmcJmTxHSYVovdYSuoX8GiJPLu47YJt
JKa36hXsqvxg5NBsqm8HNfJ3pdgrtzgRdSUSi/j1AoMw3P3Tw5yfUHqs0EH4QdSR
tyGWHrGowodiyFtZ9mx7svGnEnlO0qavyq23YViv8tx8Nr5YrGXoT/ab1+q2FhvR
WR4NEpjTh9xFQjvjKp8pqrGtSQY3/HwNLqV+ctpWPrjm9KiJ1WpfyPwHhakKNMwu
/DtHofiUapp2JYHvJiTiDkguHfTkY2lFwCAaR3ALtu3mwGvAch6HBXqjOWBC5zxE
RrgV8XgZ2j0w9YR6oxGVG/WzYgHwLqcqvl+VtA6an5rErD4agUIBjxwtJgm3rk2C
+js631J0VzbiPfUZvvkCtHj1yz0kQ0KLkIMlFdxVT9hysKAvNbVAjQDGtKKV2EkY
UAoho2KITcc3VSdpuBJtEz0BtGFY4IRIYFY6aulHkpeypyFpEe1rqSYSBwer6lGh
1ClDyJrUPo80oxbHxHMOaH/CUmmbA/ifPCIonlyKqQe4MTrsPSfA1lmMGjN7LbW9
uCNi2A5VC02/1wdjwau0W1WBPbpjN4ztivhW5U535c3u9pS5ux0wbGs9+h/tlxIm
uqh/wNwbv9T+kENn3y/gnBNTifuiC5TwjpLSQ6rv4RaVbGFiHwlMujHAb4uo26UZ
7JxdsJ0+1ijfNV2kafJSX6cHfe+vea7plfUTq/hlkR6dJymHDRCIYsADLVslCYBG
rJdbB1q8trPJe6ZO0p1cJR9OBSNol4DMDAh25agu7k5Vl0osQX+w8rj3dlZGQGle
4j0PJD2oj8Grxy1SsQ3Jgd9JL3qmdIRsQR+cGMXnd5aH/Cp88BxsWsRU7A3pnwAx
GOydOqifOMFu3vZrXnem4bjFUXInxfvprbBA6I9S+uFC0SOJ+tYTvvz1HVaJsQCE
puuY9nHT3/BogZkpgNlxMQnujErhkPFINN1npR2TBGyuLFPbCw99aK6w7zZRnfqw
mdK3iApUQtxi3KMdEG7INMLVzAzLkmp6R7ssHRx6EBRbHNCAUvEeqm4rcgn88ggI
YddOGSd6h5n2oigZREMQBb8ihAQQsg8dNXMhv6i5bp4xatdGW5B7ieBSvPUlIH3z
VKtsmLqWCh1A7UYVwUVBbkt+TgxqCnjR3sgJPVlzfzBVAqbN4AOGUcYu0UkUuJcQ
pu3LF99yxecod/s3pVWhT3Z+yvIFgistQX/QBRTdB3vP8hTm1zSERxBa413+pXu9
DUkWRkRDOWrPonzJX52eWKLHk1S64SQHQyMA34MGeFhq/pdh4kd+tMrvrV1mccf3
zdDczI7jZJLg+GX7PI+l124nka8KDlLRQo+4Pp1u6tUmaA/khTgbAmZM66wLVqi2
+Y9bAk5tfTtQ6l2r+QXMXgKgsEqDg3ilyPDDVO/lPelhzaqAEjV6hP9P5saMU2wr
mZu1aJGfeQvmj0mQ6vb9DaiYOA+ttcyn/It2ZdnY2sGHvaW0Xbr4g7nUvexPkGQp
Rs8x6UK/+wbNmvgTpu3dESYiXYegdKAq6FyjbIc9nCVzEYABGdfaoR+xoQjjc7sM
3ksfhRp5fJvMP29dT7b5sOa/j67JPvraBcgj0ctkQZDzsQ/nJNPMHmWWKLr7/gYv
lH7Zp86BRCTG3IfIeuZ9RDPJE+L6x3DVBh6XIfOm8K/b5Ka6K8a1nNPGKS2MKjtU
n44LEbbdeKjLHX+tMjNPQ7RY+QQAsjkrDj+tO+yDwdB6TskMEnJkcCBv1pmXG4Mv
cN4XlRhHokKxVE3ABpRKA844Bunnf4SXFJj0kWITVIwWu7EinMoP1vkPjpqFCdYR
pPAEEE/Pb53r9PvxPbeKW+6L24UDLoM+GyK25buEOD2FxWTWc+zgjHOi5Scl09+0
0HHsDGNW5ZVKhNqf2Ucf20t1ccsfFK8A7cJnnhtksFRYVAdRwS/4vJg7jQhXVRwz
8AYK9arkg6sGB1pHJ0rnGbfu6QmbqOZnhNoI0yzCcDIFmMveHWsAWytzimRzg98k
f922/V2t2hN9LewdvjBm4UHqX5bzX3vah3wdFacs7CiCg7vnq7YacPnTz1mWD7Z5
QSbmPTDEX+sKwfOEl+sPnv0lud/i7SPvwjaEogbY9mJFkxxpQNi61EZ80hwBnxjb
kbtSolx1nJnI247hlsKvMBhMxNUFd+uT4wjkUZLOmHO2bwUCj045cM6qNjLzrHww
/7wk4EA0ZNNX/za3E0s/GS6KnaGA1J9ZOxZax1zj5s/Y5mQ9AqnsMTrzSrV1ckFZ
TDUQMVX77r5wXMkTsWwNDEM9YcxIvF6vMWJ4CDu4DVUUpAPiuS4r7MFjQz768+Q9
quqq3kxnNyckzW4zIwmB25a7saDJ8kd4VOrj7LktsLj4BXvaK19zU8qeCxjCHDVi
sL1Vj7jUQHcFz9Y+1j/ABDW4qc7auIdfGEwDqGlShAjmLANF2ru+E1SUYlGby+HE
WPP/QUT5+PjmWMZ2cGHnXeM+XwbIcKtT52GRu37ER9ybK6+dXJBg6gDBCkN39uro
yP7HiQrIP+89Dr+8seJdWoRcyjtvsbHEsLTZ7hCvxzpakhXNTMznyY20FFP1YLCZ
Jxr19riIeYP3ahFQHLfiT0iY3O4ClL/MDVoK1KD+2KwPuYGMRIhO+F0zU/laQ2pc
I2h/GLskCUA1iDlBo8gT9Yk/AbRzoJolbUCWro84Iojhy1wxQUaUmUJQS+DdfYqW
UuaYmnUWOxBy85iOaMntKntuGrUtRDz9hwEMEcNRmF070gNN42c+GBfWwZhPNGSK
OalARweVOqkqBqODkfM/KhqDzEPoawuE+ayheslXOda5UmVa5lC9lfCRn9ZczJWU
3+eF7yf2YEbsSDZnSFMYD4r/FKaJcYIuuOPkYCjVn46WcYCincTqDzTI9I9SOb2a
OQed4RXT2NQKLSECnVC2xUGwkf9/9qeimIiBwniLiW9YP/mFHktx6Km8ydKzjDlZ
B2q66QZGkQeYBbxUcWBfvTWTTu7Dti2R10n5wD2Oc503s39jrTCibHuqLnrZPbu9
+pUwbkt6XVe2rBTgW2hpcBYLS4vMkCrtZ+tQj876HhC003gVEk2YbM8EVGV1eRbG
GoXltYnv/WhCEIPl67nogcCW5lQgpSgdHUjrP4h5JNWxRd12U5OLqTg6tof4LCie
0NfnmeaFD6LdyyH6HcPagaTNmxsy97kO33X3aw6nB/5NCbsTcX0txyqdztBtK6w1
reUCKjagAJ1VY6xYyfWcJL+BsAwwHlkrKi7+9l1lyHqgPV3/QBp0P0F+SCvYr061
tTL7lxQJTRZt4NcazJU6hIsEjv5AtkIXXMwhzBzakvULy6X0oP7Sv/hTjtiru3JB
R3QxXBQRconZZPvwCf0Wavw1ss/xG4dMF8AKZ0MazJVPk/Cl/X1/jKLJQwDe5HxU
alPS4qTJpGVQMJ6DMxrDJapfdLzcwluLGjQlEfkALCryqV/U0e/6+uALcv0wOlRY
zodfxKanN4BFqVfRagjrBX7Uhua+qJPFGdkFeTMlMtTLvF0TXk6DAJs8XJ6RKhIz
eoEI+A9bfU37lfTPBMrksZzZehO4JWxzGvP6WJ4FhUkVfBJa+fpnjSyRWOG24dZl
SLcqjKJmj5YgbJeGilsSHLrmNrRKJFYo0bJW5H/tzMEhcdSk9tSii8eyGEVZ+Tc9
Ocmu60GqmhZjuxlwM6Dj50wGXKBDJYcIpM9W3D263f3isJgkXbdLrz9L5zrErdTm
3iD2Jbho9ozhUNe0MvKjTHzUTnxu4FhHc66SM/PoO+A5hk6C3A2Gh8PUf+sXmE+r
SHfqwM5eG+JOq4HSVuNuTV09NxjlI8H3qofckl2P3KICrQ8F0ICUPp2x1JOta3nR
TwoYubHQ91/xzJuoNudm3Q4CRutXDygrQnMrIfEWoKzaDYaw30MbTM3FluDVRirA
4JtjxNeFP/Nrc+hIY64PwaY5sjoZjV1XylB1qXwr+X5X6WKgXKEPrOiwVVPjeSD+
j8nFRon8+YSUCFTGVd4+TKP3vIyv6uw3Aiw8YD+HJYGzSK5MSp3cxy2swX4AgF8y
bn2CJx8FTt6/YwbtHna8cT78gyeVYNN0Bzr+l26KyNB3KNU05SDckC+e4SUVSA2s
E+fp+kuxqEZqhtBhrTPhnJWkYhhXc1jm33TilQC7UDqKtX3dkZHccr1ZtyTb5E++
QxKfd6Jau3sPE9oK1E047Ctmy/+BT1UXuVAty0e3K+eO9FgFqPxX+VRo5utIvO1J
yjtfuSfTx+WnMw6If6v+Odiwg2pP7Q9mRur4f9HV6EbzoJB/UwrL39cco6PBEA2k
ABs8OJS3GRNS48LIOgwO5XVvpQ5IiaCd24xNqr4Rh+YUwuFd6fvzCQ/f/Gg9fYl/
couwc+MLxlqWdLuBahHrpLskCNMYZBoFpLpbR75pB2IQmQocqMZ6JR3Iu2d/TKZg
7eCnlYqR9Jr0pqv7k3Picl7p+uxRx2p478X32hDan9tUEx/9+o954scJGSXqCvn9
6n9ZGRPTKW5HAURVHtiRDcXFqXfFQMA1ssN2UsCQCeUBAwaRmj7YTe9FLNKLBBJ7
F6G0VBF1t5tPakCQrC8IMs74skoZ8mYNirVMG/88jOUhTjgE2DYoFcaAQYPFZrAS
0WUSh7OvbkeCrYlCI9HP+Ubtoxjm4aO/gpMUWpiNTJpf62RO9iae10F6yuW6NiBL
wAvQEylFkh9ARtljPL2M0ppqup/PgBs5cmj6UD5H/H64TKUixld0ccYgSMtZU5uQ
O6lyKO7jOTDhVXWftyVca/HrgXFlGoGiBxGJZelwZCHmN75KeEMyzRvb0wh6MUdv
2U+Kb3MX5a2WJ5e/Od4LUihfvR35xuOqfwJYhVIw3UO1vzpJJgbXRlD+2o6pHXGn
JFXj+9udVY8lh7Q7gkxG+o9RcPdUlr4CKu5H3nHM9+NxzZAPggDhlNXlPZZg5ym+
gLXrm4VrKd2vjgtzyaF3+6NPe/r9GdU8dqHeV73uSgiJ5Sh9peXPfM/KEQ7ydje/
Pmc7O0OgWkq+/+g/BAnOCkwQlgCMc8JoEXkXqYMNG9LKIjWZuzCzQdh9XumGoUbh
FacxrbHf9N4GL6Z8dpmWdGa9zMWxV/GM/RGA3lSnyVyO3AaNRB3k4zn9h6ENURLs
bzLqhJVI2mWSIhF2qkn+wmwbBXX6FApTsMnKl1zTxx+62Y2cMgK1bEsuUg9/hlfV
amfaeZ0QOzu02l8XQGHBscpcFpOMbOkHQdUxQxnDyqE8bm7bKQFkNS9/m8jd3Njj
juHO9JSHyXogjmUqMPJhu5WiYZNi1xl6RxFYsWuG1AimCGiZx9EE9yR+vdvUsCUb
rnmReCFYPee64+UQANzG/ei3mBy0NK3PxysMco8ZzgAHhGh4S86tM+SpW9LgD1MI
NmmdOXrgLzqHpovCho2qxGRFZrhD7mzV51VmJHKw/butiGtkrwgUcIJzWR2RJ6Dx
QlN6M91orD/1c9vyrvvtf343Z5roIkx1fizFMwCTZrTEhLj5ckT9un2k7AbOMuqG
G+RC2NsCdXfjcITUynJ8+dxk4ivAOoWmmWNtoIshZd+rBDWifIrVMAwehivv2WKe
GxoTBflCXnbqfkyUrytZeGI0bnFuz4JLJxbPB2X+iGpk6XU8fcqjjYBalz/sK8xZ
WJYCA+ysCIZCR+O4IqRGreJ1RF+qdxpLMbmszCAqRxnhVLAlCSHc9MJhQ56J/5fo
CVOUCrKEVHA+yKb4gMG9A1pABCu1j/Vb8taqQDLcThFYaJmyYG3Qdt+05dc5mL4Z
vmwRtMKxuYLa7jbwmM1PSD+Ete8hqY8p3ABRZpxudZpkFSA7lucyVXg1o22WMbOs
y+sM9PJ08Eeww+Q+gFCEbE2k5TL1VdIz2izE49zKA0oIR3F31RIoUD328jvoFy9y
++REHJ39frbHRH0KKdYkgUAprMqpAe9v/FVgMRPuY/xmkvcGjvkmUK7nOHlh19O8
KY7n+G4RhPOXdnjcgB0utj2CGzqhjwydcuZwb5GeCdH5rxQefFPCjry9ohHTS6M7
BmxreE8y1srqH5uiQXhbGQYqYbF5COmBjEIpmDfB9gpgWA7WvUE7+GJoLbN1jt3o
EfJ1RqCmvBLdynjN1BBRa7reKUyZjyEornkm9PAVdaLBybe9+StfmTcDba1tvj/g
jjR3xiK7x6YjD9TfxOe/p3I+PYMvA9nnukd/lEcsQU51ZB/x4WDYPb6NbsZmcnEL
sA0m6JLeWGJ+fGF2a8oCDmQNdxvJctnh0qvoBST1UV0KGMa8lWY1Gbi6B/iHoGcC
Of/xOp7cjuSoT5VzrZroEb2J+iKxhFoTjul4Ds971Xd88AoDjIbuG551SIW8W7ug
dg7h8Ay7wqUQrjaI/TSBYHoTL0MV3PstME7dvdgnSp/BTnPcsyvrclUyl5/GfW7n
+OW119swCSYaQmOtLxJJpe5/rveKwopt/s+osKVoW81WD7iuA9M2wE20mPHn6ql2
0jUx1b47YNtd7i7HQVVFrQKGZwREUNbOo0cSI7/nh5NW7Ok9AXs/0A613D4vdiQ/
wzGYwwmCHbgH4zUEY92bwAXLb9aAAuge8gC8b8vMBQ0bpY70w8DvqQND+AaNpykR
juze3LXHKghVN4rImai3d9AIkQfud2Zuuf5TLNasjT2NipUYIwaIxgMpJnib9XqX
COXqjHw9+vpnjxKb9EumEKccVk/leo226+d7d3hyyJ4ptvuPlwQSD/FbF4jXWbUF
6qLWIlev5LfCrtGfsLPfHTd+1RHdTK4jCzxc3mZlTHgUnxC7P8Mk8s1ZeK7pfGaP
PaGxJOdx5PlcedGhkO+MS2uFd7bo4pNePX4CW8twsv0m4eHtUsoSjvnQMY9CPbxQ
qk/3zrDklqfZXPq4GH4WDydPjbGR/t8LeKBm9qE+rfpPVpbC9pLuIsyrqtTG08yW
6iZlRTIOJeEF5J3PD2Of2vd5sRIeJ0G9hkretsHXBEymbUwAx1dlNhUVT7nykSsO
ktUo0L8rumAQFK9DjUbBqTy0i80cR+ZS+AgaVzNl0DnMTJEDUv9waAqVKmgW7OX3
Gt1TEblVqQ4/GXoDrvHqLAh5CZwgM8vcgPxVQ69bBc9qX+kl3WH31+XI9dk0njxL
nteZvEucPj/5IXCG1ZLmuz5p9xItpLFVETnBOASCkVg05IG0PG1GM0y5QlDfA0DG
2R8CwBeSNI4HdlwMyzWpZTIOh+gnwWRwAynzqlrHegkwm4bcZPeBM0RmfyLAxxNW
P9TK1H2XA64NQT9cYTofKBBdPkO9uP5+O5iYxjb1DJe2n49zsO1C+PjQtD6m+h1m
fm9kQpCO8rcr4gnCXNst1uJoSi3iQIjKZj9PgFmWpzp86nMXgTykdM6jWg3uyH3C
QIMS34lMfcKPTdK1y+uekQ/Uhr2UNO64EQpb8Ygn9C+X6s1gQC801od27CWf41+t
Io3F9LQTPgx2ZQmtakI6tWUkZKZJT3DEt2jZqa27t7zPgU+vDLa2+X84fvRLejud
6iit0mZBdgKhpGaklMbf66eOmc1e2UzhiBGhJ5fhRUHzDxhPWmdnYa/Y4gulJJ/t
t1Ypa9X+pRuds47kcXMxiUnRYqngjga4mZLNQKkNvv8gp7VtU/iNDkM3f8gGGskD
q8sRhigiNIr30pREm9418H7YnLb8q44yCbd7i689M7oxv5g8rPZ8KVMCoWXpnhoW
ru4kDc1/fIVH+4QNXHJ2r33TeqfoPAkL1Mbvng4056qnDd/ionoFb/G3JM+9dbeH
GcV1bjWfubfcRG+tD7lInCJU19ExML9pVAYpJbAyJLjpUvciGZlJDPKQnuBVyeel
NPoTTlpNPjMylscdW8HP2ujgEa1CJyT0l0nrasYY3OSwhFqZtYmJAuvuIbC4ywtZ
QfJCDiurC3yEVxUiQ0SDoE+PeQPwnAkE9iJAJ+3LwmnGHAQYe/53oTBO4+VHRkuJ
K2Xtsc6admNRwm7as7ZDtZer/R47lwUqStzuOGH/bFG8ZbJoIEiSJDbognltTPn9
21/DmDkVXRWb29AmopsRQUY0FL8Mm4YIuzATBJoQoUXnb4PdwcVlI4CqGARUQ/JT
Wi7bK0oqaPK+76s3N6zaJ5uwyNvEkrDN8Qf95NHWJX235n6MaSZ9yE15Lnzb03Dn
baebJoG4OSmQaaDE76NJKLxpc8sheoyv3DUtez2PMTjC6XfvfgCFmXHxF6ULnbS1
y2TYK15iK1DhJrzOH8OlVSk19Oo/hUXm2CA7H5QsdOjJuvdNTr712qgMPvonUU9a
nu3A6v2jG3cNN/1JSAZ/wa6xTpnzbQVjQTfTAjClNyr6fpJCWjT86KBpPANf/vKl
nopG3F9cfJiYbW/Xegpz/i7qYxcZF3JcVRXZXh2W5333wUAUg0/AGx3uUogGJBTL
WXx0T+8LCRyuU06P/10mG73pbuKGzMMLJmklVfbS/OZEWIjxt3DKofq0zevMdzOy
TFZqsVlM7k9IzHccQoI1qtBq4uJBHTEQ2GvUlvxFhCaQHZXq02kTfff5CLBuzmRe
Hl8Z+uVuiT2WMgV8lUysujjUHr1kRZG8R8GM8imMSEVhFeJgwkjLlffemzGJfRkR
bczcMEx0d3ufQtlc0KAnDDCjwVtBmfw1MBmFoKK9NLA6RlgYFenWnO9lIvRQq4vO
DSpjUTzSIxFIHO6EYw/ceAsOie4MlrT+KGdxwLeNGEFTaBNF6LadhYvBJ2diHhxD
ejRqzI+yI0DMmG+IuHdEagl/eROkWicDIYb1vJWBZyJX49licm0C7+qVMv3nNFJU
7UBqW5LkWYn9cXeVr1/noPBRv4ESa8lBJvLVLHySq9gaPl0FdjvJWsmiRibj0GEH
osjNWIEcM0dRl534UwWkSGO8tSJ3CPbNYYhlx9plSljowQMI9c9uo50xcwnMeY0S
zoRvRND5dU0LBUDmS4wniuvyEp6zjFDEOcdcMU72TbJUEsbzL4NFTH9ml1Z2ivd7
GZrL7BNYsD7dB3WNA5s45KNjuBTsoaCEY9OTPynO3go2RFDRIbAHgtYX+Q1WhQB+
F32zzvHWdwIFOrG1Of6YSe+Hjim69TeldNC+iGvMPRDPRMXxuxRCZfaRj0Cel0H/
X5GaJAuc+m5edUrWoDbHdN2+2tBhetm0IPKHWDTS3zuzfFRp9Za7bzGd0XF0XS7T
hJobBVqjJpwtyzKOZWNh09N0qv2qaBnWQJG2rellMbaOVHxilc7g6v5598v0Wzxh
Ny8VJJz5cNRtCn/Yw4d8Ana5+UW4u/uX9nzgmvgY3JUARYclrWal+CNeEEtXrgE/
tzpmcT9NjPeiavPG9F6bEdxzsmYAE2H6AFEkH8iG2BP7lHzJ7sZDSoj8IVQ6vGY2
ZX9G1494FOEl5/tnNdIfkAiVSBTvAphiFhpzUzY7X+06kRbeyRiGxOus9AZEf5zb
yR59UnGKPO4U6r2x6dq6+29uBuFsZfY3oSUbs6rxQmNoQ9ua4tKWRiNe08i2WUTJ
2KwyoWq89RX/zTp5+luotXNefNpoGq1kCKZ4YrY9VUrgmTsmtmDSunaQFhmySbDN
CEtoPdICzfgvTuZgUe/4qW5Ey6pEzJlHLp9ASvZVN7py8uLj1tce3F/6Sbs4aSb8
1dGMWrNU5NWvZZqtrkKI1AXkhUfkSsIzZ4ABBiTPlEBtPG9pz29Vk12hvSnmCW2B
bBblpBmthoRmM0eTZh94uXjRYdtCEtR9SNM+M6sP40jgn7hHGAY9zZVqQ8O1LeSo
GG/wXQ9wvLJa9ubVuD2RvLrylSeys35gVb/5tgGkEjA7tmv/bVJUgIiSA+lb1oTx
oKvSmC44JqFO/+c6Fr8iD1DF4OGxb9IwQj1yT7iqqcuUtGcfZAkMd05wTu0Hgb1t
Yma3tirHrmWNgfqK2t2SHZf5egijvB243Pi523LCv2scookLaa42nVza720+1v62
Z4nZE+DI0yb3XVSKIiHGB24ZTXx5V5/tS5EJ91h5lwrIrqj9iAeD8HuWFZcl/e29
qSrvR5jb+eYodwQNxooP0Ay2qrxZKQT7uckTOz1Prgg+3KkRB1LKrixoTZcr2HGd
7fE+N5MklZNOls/RBbUQ7yyD51KOwOsprmm+NsBaiiwsnnIcN7Qr2Av7vhg2kS5h
4kuBOoCNVraMEPqDed05uyVkdN7BALB3JjGk1HvQDoX7jnXmGnRkeoarHH1NL+Sr
5UDllrIsNhIfKzootYtuNGDTBvegLRieHhvZYjj/Db4kzzHcQzGpkHogd1oY/Y52
OyLfhl0FgZGt+/oia357tZH9IEGsYbOh7rL0KoZUT4nGuPvICLrLVYzSaZIcniCG
ocp58rjbdtbn0ox0y/v6BlcJfNyJ5Al3SQIZQywLEmY2FB4lZlrJcqk4sgM7xnY0
Mks4XYW/qtHS2jbZbJrBH5uqGB0y3r4tGLhHvl5pXgc29g1dv3lLPZK1wAecOHLe
9mx+prnoCW1SlvfmEq5byseHGxQFdsaQzVaCALQ5Yy+cPLFUu3x/eSZQ8CbyWc/D
UsE/HOzMXib9SLtVe8S5pNzra4j3K7Kubc1bQtLKPHH5dO8aUyjLtjIokD4I9kEc
F1TPTI/hzzDZjV4xRKv4DbsRkUwk3AA7voSUsA1mc5SJ9dsZhBMr3UsOxw9CwhTV
OD3mAvYRGDRczgWFK8ad7YcHQKzBXjbEjNWIhkeIYF12fgR1EZPysXUoE+W8HV4T
G9QuRblsWWC+leqO7d0JGJDh2jTZnYQ3bodYE/Gpa9T1zagTX5lfg29Ep9kuDNNq
+JlC1Apl1UpJp+HMKiKuBjR8wAijnqdt+Gtg5joPbVlJwYEo5OjBOlVrHQD0ahSA
Wk9hxmRAPkVm334M4dAd0CXITNodgd+Qzo5W8OJhbwPTCV4SdWI3KcJwp6Bmba6G
ZAuz8r17yMPb//1wjdDbvlGNatSXNTt0Yx/h03PPvRRG6rYk7+WTQlAaJnQyN6Hu
bgrhho11sLbC57ntIjmjSfj28cwpmrU0phm+OmWeQJKiDSk23gOZ9jbkKejo0Kij
mUjsyc3lCekwy7bmMiw+Qxr7Naqo7hyL1yBJJrPzobmIRRZrF9bqgJv4lWDfcmHm
kmYlIbQqt4YB92hbtzuUDu7vegfVwIIeHGVqAIMmbhlLldJnKTaB86Cl42/OZaU9
zLYKN/bOQRDXx/kJ19Z3OjsrJNWF/YrjiAV/3G/lEAmnbKl7p3iQMBZMkCAWXHLO
kW7p57yLvUFT/bhILFhr37EXsa1werdcK6FqV6/WpRmj+MhZRpxTFbfEhDLBaORu
qfvjYzEuyJiGuP0N4MTxYla+xJ4Av7XAzE/79nfOZhSs1tq7rmsaV3nsfFVRgINy
WEbw2P3Fk1vwSptEvzOP5Y2J31uTFxcHgGQAOKxDUj+4/OYrWbNCgr4HSqTGJIXw
NXONbldQrmaFSrfEhjqwFNMKFy5XDRfv/OhX+N7eEHg3DYlcj/WBMXeguRbBlesM
qgKu42rW5h5fAsWB4S1LOnV9VuZAVfWJeaeMevZAMdZegRgV1xlZrDfHM2+pq/RI
7qXmE3D+QKpfwYw+32Dk3gkWZrTn07rdzdbggvsyZS3fOF/19pVDmRXccj55hHPT
7CXuI034BsGx0KwCPjVPdVRhwi6to6OjMaLdG8mkXD4AC0Ij/wg+qjUGgJvh3SqE
MO0DwkxwY7+KxdD0nItMVOZ5ZIbbB5k0Dn9bVHctLBuXw8rugmDpaaPSgLR90/Hb
K+oNgBFdkHMjEULfDl8dI8Rb6AcZlXMg+x0gKFTOjQom55VFFxEwL6UhBl1QnKHx
8ryxlDsKOIccOiQMgO7SyADsVICOdLaHz7wgDZaOKfxU0DtvrmHEzKUsoznzHrCV
KM9ckLEbzxX4A9cpNzTd0uzbXyugyd1zQEhhFcM+bSfXrpNw3cyx/pKCKfMUsqth
wnA0jRWUhXowKoITMwTOvoHCNr2p0c/hyixBdfVG1c0g+e7vw+v4JxBdcPnwKp2Y
JahPKvwsuxZldFkz+UbKYc2HyaOVI+XOvbf+OxarOmVCSZXTRKIB94QHQqGAwJQA
WapWkceJ03XYt4lU5PFXp23+NXRkpeHU28qmRq3V9v/qzbiuMsZHyrJ3NTqfNY63
9rD+JWtkZ11zBU8MauAS1GBROyacGmqAr+Rxcbe/6RY+Pax9u/ht+gpYuOISBwgw
aON3A2fvjeS17qAs8TAES2wWyRZv1fbQ+VGlK06VQu6I/XEQrchx5CCpSXGqc7+h
BxslGJ0s0htCjH5BH2LyYUxKHWkSgLcD5zlKktbxOgpmTwSffqj+U7QmNbb/WL8M
GlVhRhjgd3XTku6ow445EaEmp2qASCG4bmyd8s/r0BvaXdgYzkMdarL6JUc3Riqz
vFF7Uy5euQD7ayPV6tRpF3DWfPO3D4AMQTfnqOGsWnmHEqczSxXM6xMw9e/O2pfZ
tB2VRjG0VBgOKJwkSOSZ+BSYRypt3KUMntI7WzzPbYVX4Ebsr5Ox0ReZe4AI5RTZ
TS5SHB6j2PyVG6o/8dBlDNtprQSkbTUX/5hUjg6IPkx7PP2bvrO2yNh1AL9JXxuC
gEkhNQ4GFmeBces+n6ZC5nKhCihplhj8PHdlp9spwnvYr3VZIPQZRX90CSUOyM0Q
rGHyFdGZ1IaZ/T2C2GrRSFbUoDn3o0ZvIXbDx886wHuAo5XnnYojrMZTIYGZAhdE
/CUJDgJWTllpe9Q16B7aHXgO6Ec7alMvcHvpas92A6zUNHj5rVv0Xo9ZD5748Si4
jmLvxpFtVBV42vNVHu65Tlzi7uu2gty9S88MfIkSS4fUHZZuGnLMeB4KEMQ4EMJg
IJRPrq2zWY8fcK1b5Z/AgdTGHJkdBz2Zrytr0ZOozzzYhOvkNacHph94/ro2alik
VMYB37khbTcCXVG7qjUu99nP2h2qqlDqMO0cuVS7wtW+dyWT9v/W+CWgwvvsaxSL
pOgCx6C2pGqRPUGknjKnFDOyhtwLnFO+P9Ux7DWh53KhnM4upN0v2M9E7lfgxsXG
MWRmbcipDEk15BozdE7ZBQhB6cbj0oal1NQO0O0F40RO6v/12gCwdTfMWBdScIBh
GxDXEmiuZMrugGDV5RLNKhrgfUGe9fGmnb+Br4/vomhP201GjK3xsVdttGcET2u/
NfFzoMKezOAJjJ4dVB/5twWTTH/62lSqnbTEpTlvtmWLtzbf2ZvMdo9+ojcb65MO
6+m3nsbbwEqbm2FAXDS2fdSijMby+EKiNw4tkpHWN+Yolr9YxHWIZ1LvUjPCuxkJ
gpklZXuQdLBj9TLF3/HvjWFO15GJFgPgLNRjmSK+JLmYmNejjMnCkprstjwt/tRM
k3aqzjSxCovtpoxsh3ud7Vw5SfvrGAk+NIYjZCs6eiW2YhrePZUX51RSepKUjqlc
1l5tXQjrlciR84i58L/P204iiFLMCUuPt0L1N2OHIocnBqXsZzxOLJefHImZBZvt
hTjAycb9BkavrC4amkdBaeAR7+Lz2y6hiX4oYtRBMD2HzZbjlMiHzx81GVZRLXqE
c8YhM4fSwcfScEXoBDh5BVrtMqtSMLlDjcVPWof5gRNRvLeHubWrO+mi933vfIkB
B6eQQ64M7cVFrXzA2jr0uq3G5qKWGpopLEHtTJd22HVzRO5e96mEaPVR0hk6Si6o
hzxXz1xz39RalKq2gqlq4veI1yKPAM3j0wWKDQ5TjoyWgSwEkVr9xi6V5AoZE4yj
lK06oFfsw4gpT+Ygk+boTh3yU10yDNTSYf/UqYuppxw3svaCh+w8cMOlAffBQTgE
nj17KdaKtBDkch6Qt7wB3OT3Fq2ise0iK0PbGjs8NksE4CP+1HnhDwu3RIqawUR3
v3jNAqdyBEtMTML/BQN47KWbopj6rdad1OuXlA4ewTIFF4yND7mHr0pweRDh3EwF
vkwjuqdkNcu88aSyZD0E9wZhUMvigO9bBaydhBlT6kLzPupkCSwCdftEh5sd3nDy
lsR0jg9PsKhvi5MIbma4fvyERLvCoobMHW4KQkqImWY4DQsj2ZxfvzoyLEadWIxI
AfiHfBFR4NlhK692el+5dPSPW8XLEuiDPEGt8jVeP2JbsP2WhkWCs/oSAtZBRiWL
1WGgxzEiMOPDRP1PssdD8DngWuvyRHb2Xk8yTvGbuuUAmbflOso/acXjbU8eg5La
C+WSjemFC68l//9QenRnPOhtla/cWgnop3JU45x8CpaTdo45Ro63fmpZQvFnUuiS
wmedEXym4wUlctKWmvRHq562KJjfQPDWrOi36UCg/g6OhepT4/MfkDmdBKAknT9G
J6ZJjKCv/2UHTGHLRhEAD/ljZuSq8PqBcUzbhrRy1MvJea5PBBONdDlSbHLQtdgn
kv0hKlm+rqmOBNz5FWM1YJV4Yy4Js/RZ33Sk/xg8Fq8eBXc6EU3Qs3OeVxxV+bwo
jkwh3sD+krHNo1/6LGr6mEBXQn4VXX+AnRQS0OPs4m1u79ic0dOjyp6iUElJdg3H
YiOw6/lALwuC/EXpepuUrlRC9IXI05jLyjqR4ZhHtB/mbJEpBnwLqLQgUYYDy61z
d9RWazr4PgIf2270Fs9tKqeBFGbMfXVa6vgvZnM3C4nDPpQZbfCdWWeL+viJNlx4
k0jAOMxtZub96iSEmw8+lO6LHetO1N3CP8lx2SWurex3+Sl/FqYC9EHa/5uzU4I8
cZwSQeV8+kJjSpecNr+0BDlXJD2/T4dRrDDSeFJzkTC5rMjpWDO6LQh7DDHwdsPZ
dVickH7WyEUbBbEjvHg+/QIi/q/Mkap342E991EldOukwGTrHXH2bVLGlAs3yCnF
XvU9HTbo29BKh6SjjbvmvIwidxI/vN4z5KzOnLA72P1wh5s6mT7XYg60wD7K68Jm
lBkOrT4b3ahxBwRUm4mAB6z2PtXAsuss0zfhLRmnm0rloSMSKuvtYWoyEv8i6KOh
6GImvH0Of8ofUtF6LevJAyoUgrhVdOA3hARxa5AiU0as8HVmDbye56IhIKOpfK0R
o5JmiFoj70w/tR4QDFO+yvTJCMV7JoYRMy5zFsq95azg3N7HA7gKLE8i/Hax3q7R
zBfL3rvgb9I04G3YqS+r2Lu89Cx5W5cxeAZTQWvjOr8t9avOUZ6Q89LbxjrWoCkM
DCoJtrjQ7FNLAfntWpNg/vh1PjclCDMXVkC2lHKaNM5Egc72xn7rZN87Sj/pqGzq
LgwpisxhOHci9Kuere3un/4LWm+IHg+KsTXTwPPnkIy79do62J+GtHumVa2Id/si
oe0ruQcj9MiHcVuuEzHK6n8UMYdFWRhD9JvnMVpYgVS2Dtl8d7K2IRnxNIME1kmw
7hdX5ew3eH+SePHqjfgJEgLK9oe4joaQPE+LacYxx37cXPdjXorCnaHTJqa07vo+
FiAFouXURcYt9FEon0DZTpnEm+ZiuTbdr++efLTQTcTOdv/KsU9GH7fZDG+65NMu
0Bqx1hUSLZ7U2tGAvGffKVbrU4eSwIWvWx8Z7i9xi4zdFmZb1d2oUq5Mc6buuC/Q
2QeY9V2m0UwZlJ1mqJ0LySAy8xvWHq5dLk1uOPIDMzFnoo+6/kO6WUUI4Kk34Kkz
PdNlcRIArGVU0/CyY3UwJdkE3VstNksdcB4a7ZdvveEXN+lcT8N5+ZXZmIVaoqwb
G655UfD834iWk7xthoGElaYY5TzFn2dq/8DfmoeAWagtbwWL7b9QeizP2TsbU3Pp
gArrLXC6b2mIofuCQYtumd+8lsu45/+iut7BcMBjifYogObJmju1pd6jRfMzgC6R
6j6iwFIUkBHo/OuhXA2/zb1bKOCBPo58VBw6t4qz54L2EiNBE8v8fymakjMj75Wt
luQxUg13pnePIc7PLQgMTlndlF7lnLv95fE6q/AeBcVdtrP+cgfT7sW+hEkDl/DM
UIuVaTB3kjj5zKPvl5PJoJsc2RDlaFQHnyn2FDWmpI8oslIp+oEKiGDXDeoXazv9
vX/G5teATFwOT61+XoxRPTOFTiZn1k3uc7jyP4YTHcgpBcf3tJxgXweTxlFOOPTH
R5QuCHDf2qZUA/r/+a8BZRQL/iunIs+I+TMvzYERHKb8d+TBUUuIneZBK6HqJVGD
oAZpPoqEA5NztRHfS+101z54zO+gQxyh+a74a827+eZIrCPePvMv0keUSGnT24hw
wd1DHdoatBziawFGTxNi0LKZ0SCU51W/nvV4MJvMvFH/XPvnwiFB0WQrRD26P0CY
qtpFDC1RvgfmvtIFS3VCSlrn1I0X61VZID/hVJTkh3QlXuyqCP9errtRTbBpqsex
cepq4xECSbLZq3WMkwlHmlc3yWtyYgtLCCueXHLrUuGf1O0vp6rLJ/fFf6qKxnfx
l1Bz6fFUHPRuWJxBITNEs8+ei8ZKEIL5aOcvyRe+JW+9tr232+HPiWi5cbACS7GP
bIYb7kSHXlCEAwtZ9236vxE3xX85dq3Zuojyu2h3RoZYAHIGT31NcU+AuX6uQFnE
TiveH9s8hmYnX/V0x+XqMkClK8rzautZE8CeVnjsEqZo0TBHz12HnpsUv3VgQVz3
w8vbRWpKXmu5Sp4uWD+VhxUiGGva4N1QkN+OnOJRZvS3izOa1er45AEMJkB/CcLS
VQe2rmyR338D2rgTXyJiI5Grd7/hcVYaMxZysX9A8I0PaHwxGdLZXpID+3RzpSek
/gFU/1DeV9UzLoKyfV2dDL1Q5hsG3gU/By6IHFIMjTnsRkXb5wjFVOR7IGe+MB3U
pCb+09tb1eVwdSBfgQpyvvZ97ByLJ3/pqr5MMvq3Gv2r7RX8Kng/thm4uQLYIJXr
446iOZC4aOKShx9oPvjbPUCF2Z/ncOoTMdZLeY0LTZYmV7J3MQ7r7bdTf0RtA+qm
gLrtgVYxmPewnkMddf/oy9NIR7ScoLMprJLAnvrXV0KTp+yPZlklk1xZIQ9O1PR5
gekcrD7sP5fuxgrY8XXblyoEYKh5StJduRoi/7oAgzVWuvShQ3PufDD55danIqPT
8iUH58whrKvB3inIJa8pt4RojiN5njz5qtI9V8muZ3vfLU5d5AUyZKlxcX961af3
A/rRLxlA0V6Ma5TAEkaAYcUoOWgBOeVdQtfMrF1aQeeOLxE+BqeE6mYVaJ5oF/BA
2sf2oTzE+LX0GpgHOr9lHopPJ9Q+XQJCGF2Iz6BL+4gknEwo3yS7LrQBO5OP1h4U
AXxhcMo9MqexmZtwxjSENFpyBOY126D21EcaTKHu++ZS90qAoyyu51OJn75wzG7x
N4UJvQxL2pm/mqC1EvLSpgfHqIs0ogKulTPdJrx/7a2DU/CRRD1pUk9FMs5vZN4L
Bdaelt76tYIgyOwJw2bjqa8rxzvQGTxzqiynzr7LCvTY0U/OBirInV0PCo6wo1/T
55pa2ybcz/FxVTJE6E9R1MMOiQ4CgAaD52op/E/cO4yvwEo33Jct6ok9HFwi+vWp
k8tEksa1qEJaP/AmArI/xwzqiTScs+/UPNdzjUzas0NAs0modZGc361TMbVVjLkK
DGhreQ7oRhZfcOTFMJD7TPZ02PXUAi2eJJNiLlDJY52cijZWTuWiQ/R2YyHDMrjy
y3PfIKTg8lnKhMG+PW9yzkaB05mOnABjXKINqYy68obZovITvjF5O9dFlILIDYp2
28SioOkj/VVcoN1QhZ6XfdJX2XSNi7gyfSgqmVN3OAKtNcNHTfjFjZF+G1lLcP7S
Dj+dnU9AEzaT4jzSKflwviV/clLm+yR7Y3utsKCzcuePQ+x4fmA2iAIGlIMxT/As
BSEFGSaYaGeCZ2unsJdL3sqm4TfBfcM6Q9rUI78Ehy3XkZLGCgOzobADly277vMX
RS5yPvCvpULI7ggpexpQDII41vh3rksdrAefdF9sf+oUzMeqNpzOSZQO9kIfhco5
VWLP7+tNpCXeAfV5s9DyalKxzcEs4j1I/LaLy1DHsa+7xro5c9ebGLQBHut2jUiq
APBcprlm8F7eTkINvcmerGgIfzpFxuumi1cXT6qN2Z1FxUMcoFIrEzvJK70xloFv
8+Z8zOBc17eAQzedEJyjmiX5NB9WgT7U90PWPLc6UmnOESDiqNbwidZqoUV2zwZq
u2GAstiAN5G9T6aEFEUHDEdPE8nHINLGA+qK/aKAjR+M8rJqfdyH5CBIIF2x1tST
y49clXEF1o0fCqGxlYKnHlnjy6h6anK46C6OA69zunvbOJj9iGr3kd/ju0er9tvY
S50Poaotw4/zwiTgqBNPJGNh0sxnn06JXnVFJduxHXdjyvUHJrQIRTD6uiuFnBAC
oVSLBT+KpDmue4bQnsmTp4clUjyqUXKF204ojVvFIcs3TcrHn/46LqbtF0y1Ndmr
KVN/omYpOf5ZiUMu0j4VAj8kS/cX5/1LK3VzYPsVprYYd4sn7+khjeiSCe6vEk/W
DAZg6xexVtGPj8KsBEvAbLDU6j2KYS1YLIBxLgW4WGjkTiFiZeAjOB60kfci8ocg
uNv+eGdodGTrdm8D1pj8zmh5Cd9dMejHTH8O4di4YFSYCTkSddcwksv9151mNXxC
SLRHb50WXak35t83ZM6Qeh/WKe96NJHU7Rtfh6p4XIXYnvuo/V7A26hl40OvD96N
cHEeo0f64XIc9bqZDkWKDeitUs72c8ptnxCrV3JldBYX3+N3exdGkRMbWsGopvoa
cHdFkHquO1pZSpyFCB5r4ShQ+ui4ryfBXzuGQwjT9EkTM7JNWji+aHAL9yytxZAT
P/CeNHAqrp+TaSXLU8m0SRPWFJA15zqtn1W+45G/behasC0U2Ct4bYGWjsoNXXAD
hYVdfq8+lQQOFTs2q4IEEZFjCC+UvK7/oJQpzdb3NgnBmEaGvSQHeYoIiZBqMo02
8EMhQYJUvkiSePZdW1v/k35aIS1zRop7OR+nJ/znTyfHgNf1Pg3HKIh1iOxnE6IL
YW82AcJmMJ/sUUscZIRYwhFniqrhlZWiHioQ7RRwMuUC8Qqy8WM+er4NlZHuOMJm
q8CRcep1rcl47EyzdLDpv81HgsoihUTEBjg+STtnrtwXbGV8DG2GswGDDrVAP4n6
lmSGzPaciZ5iv1YlJEEvHaimZTxwsIhpTcXQyLEaBJ7gK/4Ac/lycONfX/IbGNHB
UKGleiDxzndigCb2TZ36e014EHeLTED50QXv65K1eVGrzKUZujt6Mkieu75RqXaJ
IVGm/sJLdZ7QUCUFaSWLrQyy4EQgYwY7c+VZsa//q7iYTZj0P6Eo5I6QD4QPI1vH
OdwVYxqY7iImhf/EXESp5TMkThhcU36qfLsWmJemWM3I3+PdDWqJ5kw46Dj1YqGv
Z+gxEXDvXiU0bJlxApU/HVNxqJhmTsOa0Ol/z8//iH6vzu2nfM9m5EtBII69wfqD
siPP8ZuZeTVOGC50/vQKpqYPcE1hDqut6cHoGDHB1EKZDA87zEkApQico1EcsdbJ
eU3BR7d3F1HtJSmp2r8IkU15bh1KhvtkA7YW1u3gNPNpGa4wloIGK735+fsZ3AO8
1f60NU3RPX2XF8Y5JAev48XbsacOFNjNW6tl1D50N0wCzsx3lZf/3/JiRAxV/Vqq
vhka244/ee5tcXpDrs0PEE4qX7BJwXunAGnRAForwN1vs9rUsZx2NaDUgdzzmiil
pXtCRI0IRBXuEp3yNw62GaCWVyI9M9GKS+YeKsos/t79bn2mesU7BsipUOY+EeMG
/e5D5DPdg7F+VAZgUkcvMjpj/4WYnr7uEi+KeT9NMc+kwKFMidpVQpyAJBlBvzB2
WtKl7WAQoCpAr86wLJC0iW5GhC8VrLWHsSz3HGnBWFSoFMNpdpVN3EGc0Q4mhM6O
wjTWaMWiluHoG1+Um+EoauUcE2utd5gjPGr1qaXkhF70XTnNeqYBtaj4xC+8PbHV
gYAVBVDM7U4RiRD3L1H+J9kqRV9YIELhOXUcYKYRabJyepUY5c+TfdgcJ6gIx6FJ
6FUughpRoqPEr2mBe1qd8KjpuisJcCWWQtSuf5Bxb2J3IzxBg4xwo9mj7y7+ockY
CcTnE1lDdWu3Pmy3ZqKIcq/bBvM75skKbyJjvkOc9HecUqqZbJ0UBwDgUYFfqS1A
5tOubyDaGQXjzqQVdK6O9TgHadCtZ5hPfGkvP56gQG1LEa9LlenvuXhvk6dcRDtv
lXi3s3HCZRr69w/MSmrDdgk3Qbp+NAwcoklRdtNuYh7z3P8BWMGhFcgGrlDG+YxJ
lkJjz8jlNLOr9VpOnVcrQDht4qQwX5iGwY3MJi/RNnTQHFIyHhy5561xdniHsTFn
FMaPncG/pyzUzMgHyGSmMeHjLVZsX3mMDcV04V4oI5Y19uNhXYaCnNS/pemuVvkA
V7TZTWrnTQ7RBZ4MhTOyqTrd+mFLxZmPMCHMGuPBVGrOOP4g1/kl0P7BVlo+QNGu
S9NS8cNfDdK6V0Mk9qQmxC7jCDd6qYmSwcJU8cTA9DTogjlGQ9orWFARzodY5JPv
pAwVtvHwV8leM/jnzx2XdHF8wpz8iMH2+b8FmCLOFANDD3K2C5SOQSP0mFnCoZnj
fhxP9rZZ0scRFEeqC/N8/+S3WJRyzEmhDoy65nTY/yE4JToCqvdtGb/uLQw665Na
X+o61VC7+RqtG6IzGE+luhhbtNkb31xIv/CjAuRnuXAP1DbmECkyM+JktpjqSXvV
dAy+BCcu61qzGGPmJ+YRFzxtQTD/s3OVTJkzZuUNzuGj0dbyinnIZHtHetOCrEM9
jRSHOtTHLuP6O6YJqGGenQPYN+pc+l82qw6awP+i5ztuhvN/ulGs2Pi+j1Q9fykg
ZW9MVJRPiTy6YVs3t/V+rRwzqVZ9R57iyzVCIRj/iBnlMS6RTxifjXFzqmSWdeqE
PU3EsXoBJ4MN4MFvD6oHkEz0fdbbmTo8nJIbMsUA1oaicGMV94ldnv5XzjypzZf7
cpjOXlgFgeNT24AQyBf5XL+3BXnGhLhWtw0oFYCxlJ8lU/OVWNop623VSDD8aMJV
TkLQ3mtJw+8PmebfsL48dKl7Qi5hcSJcWQcKLWQSahiUbc7dvTEKUKixzp5TA/GC
G/TE8dzEj/hwPkS6umLg4HLX0Pltl6zFUWaBpXn8q6HFrT80j8Fz/QgGxcZXBDtv
w8eSs0W3cWoBTvPpeEqpzuPOjg311VGi6LbRdHH0o0fjoos4+uyvY0bzDlguKGOi
HwQcCiiDCdKQRxXaAWzL9RAlRp9KIKbpj8R3+gUY4omTmZKIxTMPS+HoK31Qitgl
7NiwsmGrHC9Xfq8LFqLhI7ei4bIs+J+xL1bDx+lRIsy48WxGSnf5xMPWast2bU3Y
BuMRjTh7peSxLWJxk9+cm2A/C97RflCVSdjy77Q5QtdMCCDtU+3YDY327EDdNNcJ
8ppmqNhEIJ3fcO9p6tcpl9pSpen3Yla0uNaG5mjzStgHAP/TScHcbP3Sk+8jeDoH
oEk4MqIfXBOkAx5S56V+zgPBZFcAVdIUz//7bm+F1nV5CcAbN7eZu0XJtuQMSzDT
YAfwQzt+0ogLeCJ+2nob9gNyr1hMeSDEZjSFtBf7QTg/c1bP4kxTgGR4V3EOn+3t
8l7Hi5iNoDngS+F79Ppa+DqQj+xvz0M9UeO0jZNzO6MUjIlQsTLGu/nfnfYhi8dY
h/9jovTGNjw3Enlc4g/thwOpjLd16sYMZb1gxVLTJOcFz2BTeCDdzGqryz9zYdIq
eQGuOB22vsvquQgDX0ANsUmZBPRDQT1y2khfISCYjp2g80yaffmP7aTKjGSAX4/u
vFX4uFgbP7mInsSfmhJ+MkSr53I8b3avIrkTqYXu0CjlL8a/HZGm4vLoZ/s5oOfI
O4+OU6qEcVwSWInsTZSsJLrKilandRTNcnH6IV+loOFt1IOXyLxignzM4KNp+ZOv
ItsGO0qjXqvljCsOL/sRkeXmeVAcUhnH2KTv9jG3ZNCrru5MjwWcfJQMgehFKUZH
L5cHqcHgQyoAPzfjpUwbluHePUALejofSvkbA25OtdmIstzjwQ6UZrUu6n2pzoo1
o2UpB88GAhqlBB5Us1YsIC3UQkpzgbtLCK687a9KtE6zWISUq/wDmcC3GRMEFaQ7
xOKz3Q65za36kfDYRUyptdpCCg7nPMq4KuZ2yVnIbtdpgKK5LSD8eHylKy0dhcvJ
z3bzWRHi857f7sE/h0lGUCCwtBwA3n0o9a6Dk8/3f0ai9F9rQo2gAczHLTmZoTqu
d1by/z3tPrIFUE5Vx7uCY0FXsL/zhUsu4QHLxAYy5olXAOZng4b6Jpkp4VKqNNBO
5CLjdo7hXyxiOChVaOj6RwV8T/kRfGyDJpacN8ma2BQrVnoGgBM43GIcRsdCvHxA
gw5eEc3K50zn//1Y3Fvnq/O7DN6sbumLrFtztjaYwCuxZyfm0h0gmQQfDIUgJLy1
78iC5jq60MSGAxHaBVANyjxtflpd3Ua1j1ykR9lneJTyJ/m6U4vRKZ2FoTU2CLG/
U/saLUpcNVZKOgn6gY4f57FW31iK877UrYzB8QiGlDgixzzBHAzw0cFTOggm3nDt
NecdCXVx7m/B9GgAITg6j/G5zCNBQ6e5+yp57xcQ1uO/3buJs6eGsZNkdVeMRyrF
OEpd16j4oMiwxMe089XNq+Mfb/HHfRyW5CW9e97oratffl7qJXSM0vFbaL5pTYpJ
fYiW+DHoNR8sHRPV9TQdmPHN9FbwYjrdl3KAW7SCwLAJabprPoeu5i5uTLAiadNT
P8wbzMW11DHAH9bDZxCOVT/bpDeTx4gKRkaFq0lLpozZG47SG5xcacOPmkLNkDZX
mt1egWYSlcZm59FQcevbzmoKr+fgZtYXtBLRFp4UbAgt6E7FaxOH/gdx5IDJFwRv
bYy/tRkQtza/dpx7M8t9Mi9GJ5gTZogeldQ3jGcM8auAkRlES68mKLj8gL+itcwI
nixtDyv16FAAHdL5+uMkIYak/XQzKm4z06aO9AJn7pv+7gkJGmPqIBbszN5DVrPs
HmsRoPoWcY8sxd3v0z/RinHhJ83c/QVzN2410g8Zddyf0H9gTlIeZ04T0xcvmNgB
MvnHGL0ii0XUm39ZNTHVgo7mPjNqlfIkr5oegVc6I4NBQvol+L2u1zB6qvXGHPYR
QoXaw4EJX5X5/pk67MFcnf0mXQdxtkATAzs07kxQo3AXr7hOjsouKa4d32GbzaDy
R/eVu3q0nYfdFGkNpNAuM7h9El1LGDU1DqFVp+tNOxshY3u6bBDkB/yMz+eLFRE5
wEa04waSzh1HBuU23ICYqxwoav+bhhYNs5EqJ9B6y30ss6YoyUN1NnVWrRwsXlZE
KZQnWgJTLclCQoNjERreMd96EV8pEH0XykBej0UollTiwvM5E7t7K34Lfq9HNrEK
1srgOd8lWwCtRIw6fn1/JUekyPCQQsxzE+K8qwbYs9krYHc/dj/1piah/KbmVkBt
lZx/wxilPOCLEZqDJu+fulPcX212uzwQumwuzeqdZNcB9jImVBKOHbYhfJSUlKLT
OvGOF43sa/cdJgfyBKUUJGhL1nDr196stZw4A4h6ntPpjSlqtScU72JpntNnzbUg
Q92BDPwjfjWCb0D8TDGVnR8v4ZAsBIDHe39MX/2xC8JwNohx+/+o5RytfIpIPWlh
FjXrX7nZ7HYUG2j6cHZ5C80MBQ5P1g/Lz1rHP+V9wjP1Q1TTPsP4c9cnl4aNqBHh
3tXZMVoLpp/lOlwiP5bfDIfJLYpSP/feNk/jbDrXXKjH/jxATxIwf0JL2D8A2z1h
XXlvCaIE37gkX4VMHwFLhhPFSlO+ILxthSbh36fKbOd12MtQXt1JvPJKwIOv+nvT
guey52X0vvv/uiiUscg/+vQYPLKmyCZO4qnlb7M6FysrjwzxR4t0sXAyldfOUjNl
HJ0iE8Q52NZRvNFpEqZSYu/vtOISIDFRP6VoJ6gEPfMHdcTBCcCPR8E9smN8NUUH
YCMvzO5HD/ZYTEbBsYPXGkSylkXWDs7iReiztylNSXQRxfnc+EvcB8B1KX36x6JN
GiesvHAf53TlxTOW1R/FGg3R8CqPvuxavukj9WhP/T/zYNNIseafPWdnHpH+cK0P
nVFRE3qJXf2f7+yLOKPF1wpj/+gUIta1OICtxhy7b5xfblJRZ1duT7dK9vMcQqP9
XcnasIsdw1FmuL5gW13Ho1tpsfYTq4X5fx03bo7hwGBUB8fpqJ4s/g5gwEYDW/kP
2q13prejim0QgYCJty1NTry+PciVafmi3szMnnWsuHCmh4Dofl1a4Ehwtg6TOUKA
/xctrclZ1sCE5tQVpP4kUrUigrU3ZUyaNeSMvRgTgKk2ga7MZk90fYF0lAk5PFPz
oA962Hlo8bxYIzNRZoMi8GaEGCRic43AnoYEuQGPkMFnppxx27tRjg4UubxaDLsj
GBWL9eFCbx83yu2n/xuZX9psAkfFRVYzvfqegYjOiwCnuP9dSKJ8aXok6UjYDsCL
kEEv0hJhhTOVzRxQ9sXwfLfp7OFSor0Y79K2g+SjSB6/UIkN+P1zjzpl2+1H9rai
mgHLTEH1Ea37XDkEWa21L78QsvP1tsAuD+XdKxX5pkmoe66ZNtKNAw4UWG5Ca0TU
o0LmtMgPzMcND68pJvX7JM6h8F+FOBBNXkFhFYN6BWOFeEmNaln1EE+Wtv5M+lYc
TazqCWHgqHk7XnJzX9c7jacWPQfIhr2mhx8+jc9To71aWGmPk/VP589Tlt5I2mJH
ZGmZhXu1iUKx7m585ymY61UR54i/bFThddDChKPJYK9zxh0LjcDqZoBlVGZr+x5U
WGBBXjYaZWAeDLFGve+4xVFBmK61K9bVWn6zYVumS96gEA3O2LWVGYh5FnTEr9WK
Hm2B3USQb/07clRgGiYwtUNX6dDsQqOxbxp1RzfDgN6MLdT/vBg8vsjJ+Cdb6tsf
0AyAd1boW3/RSYX0s64EzieJDM7O4wIZl4Vd2nWZNX7z/J7NSdSzb0JkCsFy+77S
Ibs40BckbIizFGoBHY07ksycW/6XUOWkA/dBtq6KbMGUo4hlTvFnn0V7mmWvCd8f
JeqAX8VTMhucAZVhIS1dLLkpoVOH2vBxYHl52JjoMbM2FJb1qlUTitUpaQBXf2Xd
RR/uvXcwToxkeg4k6VglPrQx81zzhjUFSkGsEfdzxF/4VFq/NjOlkavP4Bd3ex0w
r/vAdCU3LO8Ql2oTN5Z4B7nqoxX0i+cLWAkR9Z0rjNFAKV7rKoNP7cRRbafO0Xj0
jM3UkivJNbS+6PvLnZR0b6Vqb5eeXWpmaQmjwrqYQWpvynLfosSUGQrSB5DwcN+X
PkuRT2Q2Vy0uJJz1whA8+MRMvH71f2txnqpztJWtbm5XS+Vy8MExgMmt76ER5T9e
PjdIHTaAIxHiEzHkMLSNA8sgfjlHcuHQvQ/xDnifZafGDG/PLDT6xE8ckLlszXPw
qtIhDWcl8tUSWvYYtdMYcLHXdMEtX5rfDESKimtor9nw7sceAEd7YYFvo3igKet2
1jHSBajT48A40odh3Dswp80jWWtDvuiOe63rPP3RfTfu21xDX/8knBE5yLjErhUW
XyHOQwSNyFyUjcCq+D+UBntMNk7QFJVnQmXh3Fr4iwI6BXPOLDA+HgEKhcCs8taM
Kx5nz0rw0yf7JTOoObGaeCRP9+Sqqj9g2Ma+Y8obPMKo0hQnxk7U9FcoDPt3BXPr
KMYxeDlV8xS0/4wMKToDzUFgfkpcgRUWBA0dkynbZNennmt0fsNnZpdY25VsOaIs
1SRSq6v17YbZcII7AOSYrNNCvZ1D1M4wGENvvR8pDdgkRZEaFqfJvaHHc1Ug24lp
R3FLrRZETk21gpufq6kO4dKTZJNyDJp2d1oTAEmLBM80IvprgRYF+czLwn8LDG+6
jww6AFcuSIGuuZH0faqetyfROjUl0kJav2o80jlWTOBnaNNi6oaSTA0kEvPyFF0u
yQFyXNI25pzhzlWGIKzt+2c7txQ/IJmBrjF7XIfnZL7oL9GPrS5zaCE+xTo2mH99
cOHrrSk2HmLTC6CvOaG5nEF9fTREK/wgVaLpGxnyvCrauTe52xO8umzLCyOEy3jE
MzTCs9cigW96HERjEYjhiQetYo9dsI9TDz1DOJbsji/QjO7FItq8NDWTg5vJoIlC
MFzDywau86Mb8tQgw+hh9TAJzsYj0Kl1qB3aR/thwvg+y5T12NsuClbUZw9e76FS
ihiP1qbQ49Nj/XzgKT+Ujm/xpuWzWa49NhbiPD40N8nBr444MoSx0k/YkCzAtW/C
+Ki+2Skgd0ntxegwmy8UY3Eb/ZZDHze2Btw2T4XuLPdtaDcnhsW54GLmHnQtDJfk
58DNqtwf8hEZLMhgxdIodep0lgOf9MxJVCv4vWggTg08FfLoaqFUYxUz8xrX98Nf
+Vm2KoAq7iGv/CqgEYFeLUO/oHMrLT1N7tt7F8LcA8BW7vKLeZhtPmOydHMs1LQ2
/kB9ooz1Fn9YQJ5ykgOER8zkdRVEn+Nmr7lWwYUmCgMg2qGeFoGV7X0/A6e1CPqS
AD5c3aKkI3242IJ4/7I9S/5e03cXRqhl4vYIy6quVn2XFIH/ZUfrtYQjB3hQtlZS
L8tw9rLse7j9uIEddgMBNbxxxonve9HakSZXboztvbKqZYwKt91bLgf2zcUwuHNP
iU4fy0rf5n5PK+46PTP4tRndzX886otejH7QsWY6ktHowyCKlG5FQEbe6FkOozC2
eP30M2Bb4a/qX1TqDbUxtB8G+M2z5XiIkA7R+oRjk3YVep5R7WOos66wesC6QrdO
IjHzPfE49FcCCPYywMBGzNJHOUrUt47GSWcdYWOAn3eY7Ve+sKc5cZIFI+3f+QHF
z9AZ9JcBUFzjhEtJgGdC2AI8JIhEZ54J7tP2aR7NQh7X8GZqhWLQ9RT31VWOpuu6
ADCJDpIzgEJ+fnHBW3ZNYI5yYw3+G6EhfGAflQ+I8fqLe0u2gN0Qk8Q064L2cYeD
/nRttkQjZZ3Lh8Gkgr1J6Zp3ZowRVZvDg+X3jHuIKcDdHDgerOA0ZsK1EyTU1VND
/u7BJ/mAYQRKSRa0K7k4px27FdfKFTHPUmKsaoRBAqg7OdFSb9DiQGH3bVQ6jW3a
HX1jsYxu8dhzbPPTf0Rtw53YnFyIg5bepaTBTnnPfMw6EtSlNQ+zLYiM4dJAIPJv
S4P78qJs32DONfYmGsO1U3EOL/iAR2Y6IljdHeefc1oscxTCooHzl6w2fGtRWOd7
sNqz6P44J4poZoPmvaAOnogLs+/HRiQxzib+OmpKfFhMV8QVgU+BQDJ0f8OBHMTd
R38M84lj/yVQXwky8OOD4YIOZ9KmnKfBKiLVJZ51OYZyeYL4HorLKt5x13Yie4zD
UTz9VD1dyvYM9Gr2hHJv5r85NKuw8x+ApASukPJDKlhmDBmANSADhjvJ0ej45fas
hPk6RFjz3FspEiDaCcd5tmyNNry38fnlmk3vRNcu0Jfmsed00+FXjT4/kJq/a2K0
kU6p0sTK1CX4FHPLXNkSlGMYTLeWjT+zvaOTpZnO/YfE9N5xDJ+kTCIZ2s4GsF+R
DHF4hegdj8npSJPHxkOzXc4LsEpPlREDsljOXEgYFGwc5yPnbB+1x0IqoCkD7p6/
1xYrz0WsTyefBw6sgaC99y8wq28FHGJln1r+60L9fyuAh1lMOR16XCUha5BYaIU6
1ewUscXln4vaKqKgbJHw1m5iqeBGSnfCa+g10KWH3+yjhfnStVMVMachX0sCZk/p
WDcdk4z2mma1mxSJ5TepS+Wj602vC2m7GZIPt45NB5wZVXr19EIOUGXrqCP5KTrB
hIhAgDVzdJ0envLjuhtPOHPmMl1kxkGyvbWB5i9qlMInnU5J8C+VkeKELhCrumfx
3VOQoqkTXxni0TaZm8UYL2lWUS3oUG/ya7cwl41hiFjKNMIL+EVPWJ+KqY23cDbE
QUmcO0pZSdYlbkzrh1pvHoK+0m5hKOczHg0Te7iUe1g/fSWaveMDbLzkypxepsMN
xh7Q75Rw13CcoNtjIiATcU02qRHgiTbaTs1u9X/3WUmBzaUKy4yT+9GiwaYcCI5x
Vi6R0sc8+XfuU35/yFdjAUffJsvrKKQn/vDCmfjc8+kXKl+ZAkgZDOqO9+P3DUHM
g6Gn7xrWkE5CjIeC6pOzMcvmaHwr+cUDLQeyo/2MVbFHSpVOE13nP8pef66gnT3V
kYWvMIozRxGdMroJYBdoKCdGHlgvRGvq8v+Q/LvJzsZw3cqGSl5FAHUNCEEFvNYo
IDHAnKn77TpzOh1x+eHbH5OHt8WiqoWa0prPt4VESu3zXUpPUELwqFwRZDEwXQjf
5yJpm43Os8rTl2Y0CaQFWZqev5El02A0sARh3XXd70J6kHuITzacwrfdrfVpQJEG
YKPmR3h9EKeOmFfVBcVLR/RzjTf0XwGtb+ez9bFoFcAmtxSSGlanyO7yargY5WTS
V/1wzube7l1nVmYh+YrKOEOSEDcgF1gpRlyZ5JXj8rJ9fB6LsnZhOQFqtukz/P+P
LniYTecs+YUKx6LRWuLzN03gmVNcSKFnr2SDAbFjjJTgGu2OPGn2wpuUGmEBgsYy
/h0cMQOUbQjgb3ZwrVMr1IUfW72+1bUL1iXh08MjnrfEyc8OmGKUn8oKtbyqP/wh
cqIu2Ux4NQLyh2w/YZYGrK3oHdm0JtInXyy0TLpiJ/9bBhonZmLndowitC5zHpPW
nfNyCBooJPOFqGid48d2/p8amkOUC19N77uqG7en6jU5q1TJnq7U3IIG+9Wpixnv
8el6qdThhdFwWixlcafjzQmvXxvf5W2oNFK/RKpBzcP54jD66hYEzyZaR068srd9
Q8hyJzQOd2NsjPll/A/By/BmEU79Jc4uo33Ztt4Mdkk1ywCvr0+XEzuAJqdKjRHJ
IcFQYAmIJV4ZqYRXMgWq8ro6HkpLJVX0L2CFvXGW+wj2IAfEziijA6QSLmE5tyWV
Jt6xB0mAlMbGFY5H66dF+kCnrHPJ+8dTdiOmV9s2bKrxZTJmRjBnnBjO0sSXXYXT
b7Q19A49CWs19HU3wZDS+31Wb+pqi2O9yN0/CK0ZPkZ9oG9Q2TMHt3Bg4AMx1Z4I
IbEALsIuW0bQn1/8ZB/32D1ksSmbzsimbUPVe/Ss1k9zRpu8gjH34xQrZh7V7P+N
K83mqsJKD8FM47UWdy/Si2+VPo9s/pMZ0cfaMmuUU2Lo40tdY9RGUQkHAFGqG4zA
vuzN2wt0H1UUbGTuipo74EtBcBnMPFHqSjPOCmpwNTsqFAjpGP/CY7rDWEixCBeO
nzbxkAFiEJP83ix/CzowVtZIm23ECAtwRZaGKazhiTMu4pUHGjLUgz0/JEyHeo7i
BiveE0aSj+K7hXEQ9lsqscwbQ/zHtgexD5vQL9Yq+VxRQjjEec1IG3+Qwr59K2x/
JR3roitIwW16GnUG/WQyNgI/okCodWOrYCvo2EJxWmwaVSodD/C8Axa5M4cJdkIT
5RILk9+ZFFDBCGQVP8XIuK5Ia9SqdddEyq/Jl+5Kq/Rl2ASwqlIKCVIeqC9NLVSy
mqKyZ/qZcLtbwp42hEa9lz4WcRycoB9CSFJdouZlZ0QvJOKsIL2aIyuRG5Pjp9k4
OAKueTXvalE4MbAgM/sNds9Co29OW9STU5in6vMGVEhPkncyXFBmjt2W1IFDCssb
vahAike+OD5GlcjPpJGeDeLHf8J26M9CKfis+dowYI9h2qqg/VOgzKMV7S13h/lm
CIpihNLQ6WBY/uWPmdxnkcvt7fKyx++6ADK4RD+pD7gR4Hcs1AHW/tvgQWEqfsF6
lq663t0E4NhtZA2wV431dMR31m6MiN5eThfN7M7Evqb+5nQuMVCfejX0749fh83Q
wpItDgSLrwJsSU4xPoPeO8cWDtxHgFjz3oNJO5gsE1bxexgdRrummRx3WHZtybdR
KnrSwQVloGBHXOzk0v+pvWwN6i63WoF1s6r/iMwUxw9vAeDOzmiCXix/sT3ZxYL6
boizGi6CWQMgdYJN5XA3tux94/hT4QlMi9wQ9FlhUC5rhzis8Uj/HHXKcVhf/XaO
QHxMrer0L/WQmKBfgPJd87o+R5vtbXrHFG4BOPfD60aYToHC95pHom6ikLA6ooJD
QHyPBGap7Ds+H0wiDUWn2Cc8IAgtbteuloMQXIY4OVbH4EwxEvem7rR1YO+nPO5O
8ueUzLnuOcPHQrVQiELbLNnwMN+pxnseEjhF5wfKvUq8Ehv50NLLcIFIRyFOjuT3
LDtaS1AEyEMfDuM0aaHjxl+g7wmz28n4gnOfrzPcduX6aHrTzpaxnGkKw8YDXl2E
yy7sk7FSXl/PE3MXD2z4f9qGIbiruwqpaWxOQ5yhB758LE0U6z/ZBk1njYA6EJ+b
FyoZQsAX7joAkLfml3NGxHlY2O1jrRh4Jk55IL7VPbx9IR4CRE2N1UtCKlYBEUOn
kKK6qhYTidKXFxlLJrsrvoQ2EWyniakKDhsG+MoEZ+km42Kl9IfV2qGtJwThMO79
dz1UVQbiS164muAyZIW2FCgfEeE0d0K0IIoVI7d5/t8ajd/mzq4xrSJoGWo1lzWe
dv1ab6+dYaHAPjxkhWN3Yn/48py81jOm7KTKtwd+pPJGplkkF7Ul/dQv18BxJDdY
5oJim8txPSHuGkWHnWqDSntslQ8hVaiNiAzM+Z3aVEuIOU5iUV40qU/kErKGjZqh
OZ5aKsD9xF6Prj3GDPZu/vDHavgD7cuBLVqqS6nDpAhm8dpN1So7qPTuz4MMO8X2
QCbhPX0znkvzOF4wPilu0VN5xTbX+gHKBGUKbUJFuwGWGbNohv56HHPQ2i9WNfz1
g0o0gGEd2qr9v89IY/2REx3ajuYQsVeOqwF4P+FFjV1VBZtemejEUCzdunUdpuqZ
0SG+l60WhrFkxAefKAqGUXFhorK9Eht38TzEK3kBTFqjBmwj38d3wPAebLQEvB5J
mXmW3zRhl7vewsHxRZnjiNfV2DbQBj9E0gh1U1BtRqMpQSHvymTtzpoLqQgCX6u0
w3fhOdK4fJIEsf3VsjgRYeODZbqm2pMYoEKMveb8thrvmOakejffrgwgNIfpEKn1
bNyzB/qdvjtSHWvWc0LXXqSOVq04WZuHBE7rciz1zlMLCeIE1JYVZ3OhpSXgEYZx
SiwOtzWso5r5Wc7oxzVuaUMMQv/aGNZpdQO8Ao07jzmvFHob1C7rWToeYYGhPN41
BeRtM4W2XEBx+rw/kky9DrmMDC95BbCEOjubREBrpodpUHOP0+OArUL1zxxuH3nJ
uZ/rOtc3+rGbaPyjn0+oIlf1YN3BrmeVmQZjsx5CX1lpRPm0hMxQdjP9QWTC/W78
K8IHtidSc88g7RcWrgKaHnhU6HighLclTy7tj68WcwqAF2U5ufTk8Wiojpntdid9
dqmfQ/z9x4Vu1Qc5xjijLMlArk0wLX29HhOo7kX3Q6hf/TUR+j0evZc1OnScxddL
0BQ7zzDg4M1CujeOqVAiG3443xF1/LSwL+JIpaVJROl1NuifT8zU/i2C1eu4JXQA
fQkH0vjSGj8C2zq5uL9WiWETqBBvoRbW5sIhs6ZTGoc9KfrLDp3Bpfsm2N3EsmS6
iwx6KJ3hACu+MOumTcu4zBbQQE5JI+G8XR38dB7wx4sQHylIsbbPy9KZwZhwNkpc
meourgWS2tevm7NS1vyoBB92pHEhuosM/QyWrAtIhj1gX5EjANS0HlY2JaG53ElI
PW1VnDekrfLegDh+dvOh5eUyF7xqI4sJtr+fqnYzLXH2FwouWIF0w+KXOPhHxq1i
kkpALKk9qPZmXlIOlpShnjqL9p16PSwCU5XR2E2I+ty6jV/WiaebJUnoWY3tNzAq
KX0jie3HmIELryyCL4axwwZh6ECO1YWBEkvHzNd+09awWhxfPDZbzATB1FSCkXeg
gQDZ8c3skCtVRLTXE89kzvlxL+jVBvUnyeMuyyoORXpoqNu1P8E9CGRqFWAKUdAB
K5WlrxQWmfDeLxc8PLNTeT0OjmgOWxAp5o3hSLJLE3HsHeANLFXxnXxXwhjzY78X
L7mRsblxXq4nU2Zz921A2I+xbZwZ4r1Hpwa+oaGRWNPVHMFG5fWJizvX17UuPs82
gU+vYh/mvnP0bf67U9la+ZW3aRqWAQ9KRq7NR/spBsB4fXrC4P3P4WIsJW3+be8J
/teivqKvZ3uucdkvCduiSn3d3CntuEFrTdYp4ugnrMKbwDfhpN5tSGZNh2K2FOJ5
NL8uMiF+PGLYqdDPBXLktoLPor3Ed9816kDhEKDbPPcddoxFgDY9ztnzzmOoDepD
9yWLew+BCgQzwze5rqHvu/MHtZw9wMplpTzqDMubMaTTOIHoLD9f8tM9XmpGCzge
zb+69JOP9bg2tSM9qE+QEwXm5liSU69HHvu+w7QTHdTipocQ5mbbq3sMeMWPX3aZ
gXX6Vxcya7gkdWSqYXHO7QBTjiloVoZPs2YcLE5MR34VXK5XVud8jWlnyCovX75t
gILk8kO5H56IJ7UwNP8IqhuH4uvQc0Vt+v4T1Qx99QpC7qIn/DbF1h9jAzXnPD1Q
NyqOczi8jRNsxf3Gf0GuYowJqdfEO2GjGAjyS5BEDAx8sMG+caQ90HMsOahu6Tt+
XSvfRs0JF+dSr3lLo47lIXyTkufcn9sLQPqjXLEFJifgUSRwovJFYjVBtejyKjBX
YuSYKw2TezQxGTsMCayRUDBhl7LnrRAqpVsejp5Y48V4CsshFKe0LOt8uezUqBLR
JYsFdY2L6AbE5yxYy1RicfunGDesSYGHE4cIrbU7ekq504xvOQKU9/2oXd2GzZUt
r6EvsVHLsJpca8LkIp/nhBsBuXnS0rpO7jbNuDjYWYH5J4CkG1IV823lmdgAENjI
Z1ASSnr6NE4JKnId7Zc+S4qEojjwU3yGFr5oka2e3/ghJCbBTxIfC60s6crTin41
5ElN9jMzQD16K9HN9AhflLBqpdXRZKmK+IFqGBsoZj0TOLrHhoqdQeSd8EuczGmk
4y6VrvlIdCudUiV4Bg9IYTtgA9giFiit13liJCO0qFaeuHme6mFi34Se9P/QAldE
gpKDJh5oNB0nYyeK8T+AM/FdFsQP/xtfRAeCWfJDjEms3OLCeykSJfhwSc8M4M6q
cTraFYJsQIFCaoIYOfzBz7yfpwhPrnh6jirsX/dIL7aqktp0Af4mDQB7rBKnVHjK
SKNLDEmXKeglTJz8y+mRdz6O+arGdh+5h2VxIgnUYv/AKhwzXRC2PF9fOqSkVHc9
6IFHZ/WlMjMWP8ft0hd2CtSt8M0lvnmrERfzucefKFj9PZMQD/ZdDLPdjCFaxPOU
Bmd/IWTyR8U1rTjBoic/eYONBnEBe5Uk7dqWM+5o4P44gOkhQYbkSRuy377XolTE
zv+Tn2k6sJvXdGvzpGyPWVwjUbZB1k7iUQYDAv1H8aG7SKYTniYxSh9KgCnS9+tg
CvAFK3qyx2QnapUw5OtjFfer7t4mzbMlFhDxqFhsHBf7I1HlQGYo7HbnyIoHixqf
7l1YEUgkwXptbWZTg/2lopRzPW5ZzeSnPBJTJUFZS9vD4u7A2Lr0oT9821Yp25fF
YikXEoBNwxq0xjoEjkr84OQBjsmQlD2WWPEf0aHd3ElApNBRKWYqUqboyDsafgRu
SB6UfKHzOey8FCcCeOs268/pdSNHWsnDjSIdcOMGheqduKdwURnF1mU4YSKzsdl9
9N7lH5Y1AyDJjeJHEbivhp3FAschO0XQEE0oWAtRm0QjKcIfB0B3MAX+1hd0dWYa
t2UyUrrCgaVGz+FGIYtWH6PkfvaBUc30w/iuI3D0dJftkUHpF8LSzLC/i1XUcFwT
UrVkNT4AbiUhff7j4R/AQxvJ4RXqaHXDmzyZlmsN1aDjAP/OVCmOK7LHHXjnIWqw
LzE+PTl3mVLE4744ApBYU/YF/MiKf3xliYEw29heG4MfQBAsAXeWTc5fQAMZUYOy
Cy9PKWmwqVH/0E4DRw/j1uY/EcUNdSVty2Ox5xlMnIAv5GmaZ5ZsetGnUg2XtZ/k
YDNCExHOR5jaEAKiODykvimIHyB+DjQxDpbCBxW5c328ps9x+OvU7VqNzdmYmNeo
RdF+2/Ykzf6z6ZDemUSfmnXRNvx7nHnZpmewOtWAirXk+EUpfrNZCGxPiIxpmJ9l
y40JoXuwGO7WNph747nQ8zoXyhlAaX8m4nx7GQ7cjdp8AxztlkwynaqIlDeXQLUA
bhcRCxU/kb5wDC+FfWIrNEY97YpW5KpzBaKgqHjcI5V4+fEkqWALpBCBO5LJ6ZMM
5VBxTF72hq279HLy29KiA2K7mWJvFRmrHEOAJmGfHcbS13+qmBqMt68NdvhE6ybZ
DVm09gV7EOFToPDCNu5N+7TP6h61NQePJ9WuI0SP4iv5wrUOYi8T+TPbS3kQM27D
RahHzSTYIh86Q3k6ZSfuOPo7TVLDuG9CckrwgjHm+4gHpw18S9Dls/LdiPT05UlA
OAJiKhcA6609ZFRIJEKpu+lmjeN9u9SMEcQZp534e6dJ4jpv2Vl50+WqoAzzREct
43/oOlW5806TfjeXrrnAlVogMUmgzvum2SVOpZrqZsmNhz1GqHWs9g5VnUSVcwSA
GUt3cT8iUcH/ARQIRlbJLCTUd5hchzUK2q5PsWOqs41AsIgUD0o/P9qwQtaPWXyp
Qgizjsgpb1Lqnod1jETTGyHJv4Aiz1hFzOGmWmJeTqeL5IvgPz0Z8EGlAvP8aCiK
pOyfeHYAry3yiWRhUZRacAD8qgXeAQRI8WLs5KZKlFGJVncX1It1ZOLbKeYDKtH/
kldhDQnQn9ZhZgHbKLaNieIoMa3jaNdfPcvEH8u1iIMtAlKKXUjfxRt1PTH76OL1
gyE0fcfUqCtEwPmJ6GCrF+AtndC33srAM3eDra9hFNiJwKlZACrzizb3bksWi9dM
kvJfqQMlHSriZGI6qxS+CL6Q1eDqI7Gz70uaWtQWKiOD3OhzrJjGzoQ1Fh7QT7ZF
vf/hZ+MrEQHtlAQPi8Ahn7K87MBy4zvxV7TjxaOSwlQtRv7OspBxJroZfw3/0IB8
BdNxlJ0IqyQb5QwoezlXxCdohYN9lHmu78ugMTn81lI6JAUsHMfVa6gz/Tt/+Iub
yeUNs8RDnmofedW2diQuIMWPQtxdeCmYFSEsW6+PghTbkUqsAQVxZvY3nSmvAW/6
5blv7mVf6yE4jXIQsZTwmJVuf1fCCCHWmytkCC+IN1lJAqzsRytMT2f3nikbMM4y
HRmksjAtQQP47lAbVqg5Tvi9r6BeO7iG2orXTsnKk1X7irt/Y8cdSOtIETmmzZc+
8OqvWn4azpAhmL8tNm7+nSWt8JcRs7Ja30BJ9pakpG+a8XzZm3djPk7uGJi/3Caq
IzqGA/KQBS+HwSuuguxRnXcGfPJjVt3WYmolsfWWUMpuxe9dYiUZU7ASADkdp3UC
snHAy1p0s+dQtXG+Vd9nG27jwyWmKyVU/5bRnznWDEaNClQn+TRtfgTTCEu6Ntfm
7bW6q0AnPd1GgGoF37CXQuSC8Mb+zFtbc2RnC/E6FJAe0A+X0EvJcNd2sEGUuLQx
Epa22riqGcXu8EAS5P+eMP1e5Akqq4mgj6yObroBP0yVXOlVUOmbXN1+1YyEUdNe
wa36/B088X8H7uyM+wL+xS1hLoftRPbJl08eUqZBw5kAevucBSj17VPGwHz59YvF
4QirtAJvvAdrD+Y0/bQ8KhnK8nss8xj5LlaEnKUYg1SWAWAYqK1+ZEcoe8gNvZd6
+0F+Oha9Ug5vtSgUVfk6KoCkwcJSjnXKYlHlKkKlBJzVGzBeeCunjQyUMHYQcSOh
qaR4uR+TnP6nyoeb4/MK7yAbh8Sckl/AxLsItnKfaUeEjBQqcQCBqWJ/pR5yvHND
rs/ZdCteGeS9Vx6+mSuqERde5IUqMq2O2zz8twywK+qB+VScVb+X+If2iwK4NDgW
1jPVrbK5AC81awSPGhjcCxrFyyAvOkgCtMTFT2tqvNk73nurXADeSpFB9iZiXD6b
rFWiIvhhwzVSSnpq4kQJWnE5BW8ITu/0Sol0omdpDQ1Qxjijqc8zhR807Q62gt93
8/5EC8pJyMD7QkwMye18H384dpQz7Gh+a2f93e/hxrLzvwh22Ms3WDwNTFPJSjTb
D+1j59AVQ4rM2lAt90rtu4jt3Cutat4FvG8vzE2c7YYC5DQ8AjiVNNjHMkJvd9+6
FzksfyjfzEBYIa1Edz9nFntI2FYtKoxKOfxSvaYWo5q8NxIhNYY0fPm67YLvAUwW
GezdEcSmLq2KbilsKuzeB6m934uaK4Wi3zBTz/MCWa6K4oe1Bh0u6cgyhFVH70w4
xQpBur+RzTNcVv8tZLEkzgvpw+VfeuDBBiu9duje0swyiFm1UdTHoJqLw/7O64Kq
sDmsQx+YJ3SrObxcO0EcSOxpyhEewfYxS/xKzQ4+MCn+Siu0vzqxqWKviJwiF7KT
LHuScyR3aFPXamejc6/Y6coP2dR5iyjIgN9+I6YHZtJS6fmrrMFDKAMxoItmP9ZH
QcHX0cIbgARrPiEBIiTrNi6os7j5IXPlNbN286hhAeKHDWH1n/edJMdMYP9rLrnZ
VlCqWNExUXlyP6H/43lJaEj/H7t+ZGbxEtqvvI4MlZ8GftbkBirLpax2qHA1HXM1
pDUPAWg19EpdRL1vya+63y8y3CROmXL/6AQQEjvdAekL4XwurCF5WmV3CM9Izb/9
uBWZtwV5AiR/dQ9/6lwVFRUAjkbloUOrsK2hVaGM/sX0ocIdnPyTqK9AIszV0yM1
GVfHZYsDnIPko3+0BNPslBoB4mv2ApvzYx+iUOpI/g5nVpfWKULdXRqqJ336L93H
kM6y9BRb9zopCXPxD3kuCpyeD9UIaTAS9PgEttT+jJmTtcYYP/Sb0qycJUmC+QQS
Ha+IEklSQosBVzaoXdPWPGNkOvzXFNqqsclxnzeaphEnR25F37cbsoS4wcpQSelD
6c2zh7Rx4WFERxPPr/vRRkcoiA4FpuKjowryycZq/d0ylsCkPsxxz7a85ShDDwED
Ach/N4yke1+4AkLmd0LwsMoihiHQqyW+QupQh9RFyGsscdl04tpMd96js0mdoiW8
9HzleIFymyHtTp+3jM38TfZFHucKdk1Ibev+ts9ElTGHi/lAMmIX2ddMdhHq8aEv
BisYCEDsl3s6TxvNy3ljgAJ9xtTC2HJYSjY6OY0Ex7aLRH0Oytg9aQ5v8v0TwTBr
O7J/El8982kVor8Z0ALLoYlbJTm47CCFgfLt5jHLm11xQHaCNErawPv1bwNL7pWe
qItPcGzMDz4rX6hcd1Io3IK5FdxFOw3Jw9Wy+tx2YELxdgps1svNN1UsIEa43HY1
F/7v7XBstsGywpNJtIEJvbc19ee07jOcEY8PrLwuWS/eGaCOLJ9m+3oDqquYRXF5
EjF0omJcdV6rRhtHrSUo8R1sGzq9CJj1ZKbrSNEljp1YvJsVX9RRygh4MdOnv9rw
R0SKGyaUyOHbFAG8HWuIcHcvWjPQVLKmIM4nppuvUKLx/NPoQieJYpfk9awH+MU3
wxLWPItW0wzlI5w1CgDxZftwuzKncFqMHy4WAB59fFN9jmvvrlTB0ryLuO5k8JnP
FQWW3TB42aSm6rm0kE8FKfP8KOilooHCidfTUtizdOpmyS/hAarDXbyLLpDt9hKl
R/VtWvllwOfEe5TRT3OYSFqxZ96Lcf7tTR0sSq9UZI8A/eaWNk/TbW4L5/jcSBgc
tiaabMLMJs1Y6IqHGG4lTOlZSTTMPrKWNnLkUcDJ+FDwlyDzvMArectE++MMIw8Z
bKVMStyajqf91Nv1enZMaCcM3bi7wBq0dMZFOdJQpdL/T/tcG6Ub66xQkBHbcM37
MM9EJm5gDvyGjVPQKEWBt6PMY11s03sQe9HwlTE6sRtGt3jNHHyi9hEsyikJLwQu
SfXqC+My7ouE2c90T43pseN2Ey8t++2Qvzj3ufrJBaI1a7XMLYLvt57VI6Nok+2h
hIa0MGqMXq2QzAXBy4Yfat6hJvr2xUFQBg9R6H6xUCq7qxYuCMndKi5F+yI4nHo/
rSaIv8A3qeLDQIQwg2TKJE8KHiDXkxolWDXFJjdsahE2zvyvoOCckSrJDlpbQCa2
ASfgPzCFeqbxnnvcfL/a/BWjKJcGyuhJk5amdj8trJ9mSwIROZMTgtHV/yhZN+i8
t89HFVuy+WkSsOGhxQ8iKJ4aHxJKVw0tqn7swOa3oPv8T4Oxc4ZCn34M0/F5GzSx
hoUIvOCXyHCrUofXXUZR0CenvCA5Fl9Lbdy+I4yE9pWqYEUQyLq/sk5BNYlcCsz1
LoTFH34uzgfDSGRpaqQm1h7hkUdj1djLSbD2mXRq2VUHKBH1xOe5IGHnhy7K89CM
TJ5q68q5weyKlmehECLhQDYJVKwZ71mdcnNAsibpUbh1knQAEn4znRoh/dADNck7
GamcR3SAZtenWYTu2MMARERKDmBQYOlsA5roVkG/LSBrwAZ8kcFlL20jzof8r9Ky
Pumo/MsapTOwvDPX1PNV62tzh5jK2mANdzZ7dk+Fajo0TctkrqGOqZuLDTF7Ub9Q
zBH7uT0qw65ddG7vprY+ia/3w9+6sM1Nq9KeI/w+1jAA/KpO+1EoAolxrO7AdzdL
UsRuyaPuypjcGskhxo3QNNOJtPNdlylx+35pW17fD0RE4LyZS0B0i7c1Obu/QXJi
m/XcgUFBU2oXRGWzLu2PK/XnjqZ7mISf67G6AnHBbU6SLIVl+j0ArU+H8cTiSmTT
eXbO94Rl2SUMsO+2fSdP0FHI8pLbW5obSEp8ewSrJTgoBrgZqfrRgeU3V9rOAhIQ
UlJBLIdH1fI/26Bdlb7xXXuC1mv5PFUGc+HMFs68DjRcy7l9AHwlGPV5cKYeMxVa
3E1Vf+1F4A4k3MGZqbSaQm1LYin3mg7QtsRN0thM/j83dHJFpMHzbeP1dvDLeuXn
chTA7JEZtnW+keyk6K7MT6PxxvRAWnqFk4SWDHmPSi3PfDe4mQ3VdpdwfB0NzrIR
ciPljxU5ikCA1JXCtQbrZtjhYhg7kpZ5IWs8Sod8wC0rcUzZEtf1zhJyrYgw/tox
ax5m7AyftSt1z2hxRcmt2LnZ+nZ5grMWrN9t0q2FTyRQIvJbQsFX50WOhafboG/E
OqWe2tVB1oSQ2nY12RqeitWLo3e1VW6h78B7UDsOlRQEPALoJQGm+5Qc0dJvH0ea
KkCeuuMUH/CuGwt55eL6+REFtaG5+JEimFIwfjbgp5b3AiWqbVOyowaSOh/Nzvtz
xs19OSPtiSZj4pO+l+xsEzhe57LV1A0guXWArf7KUWe/B91Bg30cSJ5FN3ENWzhn
PA7d7weMANSuJ2a7g1q7ct24TIYCCjzor38qNIwGnwhjeFsQreDjRw1CAlPauzFv
i4uTSfx0V4GiqreDif46nVRNp+hL+uUCYnxIVk0DEU1zTZvBVogSN5KlQykst9Ci
3N1RUjuMiJiRZ7K2qLdTlewU8d3i6lLIcBlk4/e+hp/WEC9sDn4s8gLcOk4Kr7U7
6itw9J8jfAWBOnG397w7DTuay8Wxr6KtUYjsYxR9EZROf/UJFJ0PU5AAvnekZaEd
evN9XGZb+SRjKVo259VVop0wle4+VAL49UZNSOYKS72yY9r2bi+y8pqyM+/t5zBH
9lPCos4HWt5QrBMJYT2JiCZiOFPbzocXijDQmK8z53Jt9yWcOlXRi5XsuTC08gZM
pHVDOjUgrGhgLsFobp7XwCCUUVlATSA23ERMM9qzQXUtSjzygbFnUwfguzRSnXIA
1uSrloFRDTYSPZGE8G2AFKtkzYzKZuJCdSwWkbJo6uQPUk0UdIpcMbJt+NdadInS
hFDO5LaSRd/Ndnm55S8meLq2FP6x3/zAQI51ivU5N/+rbV94WWife+qZZNgtU12G
9TSUE+SyLBF0G/Dov2QPyVpWTe5t83868S+wPhEFan+ZPA3+7Z5SNDn5FPeFoDHw
p5dItHP5lS8zl547/HWjABJ3yOe0imnFTwUE9K2dF0UWTFb0kqI4k+M2uMq7ZqHy
BPrcoRZb7q58ifkIxDPJs0piiZGP5OaV1bIAMKICTZGYUpH6I8VRBiz7InyDQ8P4
nr43lERUqtvzrZJfPnJPDxRPLDIhn1srACJauc4NyNJuCYmtrCyMoa3ujkA88GZZ
935wmjqLeVU36KjEyTwtodhsX7F9Dg3cOihwg8Bwoy3t6WijV71d2Ie6PS0DneJc
IflYWP47dzBLbGA211k7q4Qw0tS0YzWEv84S2MJpAuCDX/HfQdkjnW5EK9jWnZ02
AtOKtCyMuOG+nTdMY6CaFeKmxDKhyUwnMiMPhNlpipIUwOlgjmGde1r+ID0ctxc0
FSKrozkrgA2yx31z0sK5u/h2sfYvzOlp9r0933BOlqTOtpxbhc0DocNTst7AtOrp
HRr/oFfBcwzqeTF0N0xviZ/2clUjTMvHo3RhYyp41D/yR2c7dhc91bbxcGGlmqYC
OpRgOMGL6GfD195L6RndFrnp1xEMRoizC3C3tymmChn+HKWdNY1ClxI+9G1H+evj
HNNNTZ+GYHPEC8/MsC00VNxB/7JYrQ+XuHEddtzF1khO+uVZQgcWltP/ynkEc7ke
czfuoyG9rOgbtdP2aqFq93YAip/F3R9bWnJw5kMWIgDbj6bRTbL5o2DSjGX2GYcN
Tq0vecVoykp74pq6JychGuXX/jRTDU99dk0CiCaD6GxPnpv/9q5xm9wLEjk7+f7m
9EByGhrGw3ZfUZeCKJ/sTfu/Vl1vXsUxGN63xCeK4lyIexX5Dq0sZjzXw4UCDVzc
Bu8MMgCEnIWr/iL7SCz/g1hwsv5p8bH+KloGHX1B5yyYBTTiNM+bDjkDvFNgqQBx
tpDp9KCrNuIxZpwGfwnbvCayBnxCLFNaZe84pIhwabNPY8hqPQCJiKoKIMKicM++
uWJTeKix03g0Lwfb8qyBryYjcRg6rFZphPjTR0H490Bz4rq+8eYyNRpmsxZdl55u
7k/Q6w9FuWyv8N1hSJKdcLgcrxybIGZuWgt0UBLYj4/W00gpfUWGBJiM/A1oZpJe
xhD58dOxhSrvDFQbMlqhOsx/SRL5PL9XMScElnkpTkjJJQVzA1kM4hoKD7dGQ+63
lAaKK4yabZzGGFCBMrZLUaoUvniCyo+2mikLq2cba9OF0efQPj/masSSHwkucxtR
kql5qrXawhdbL06v9gLuMQ3ChgZitT6Mko0lWpH7Njp+qwfNKei1/fJYjIslOFFI
iCW06CKpfRkft/TPuP0RVVnLnhL+GDeXQp/JvFo7cZEEm20sZgXKHxVyxTrkRw+/
O6QV+cla+XfWsoPJPrrRU/Pp5oIqwrdxp2hIFySL3vxtZMe1gTIOO0Utla/XNiHC
9LRYn6W2cvvbtSzzEDbru6W31PxzDtGivliS12aqdSHkHbq9V8KkfttptfoMab3r
u3HLQkP7L2yWy2JhTdbM8R7euJ2xAcvg5A8xk60RRoVHyNdRrt88m4SfdTWXQ/t6
rtYnm7OnGyOSV1qo3ApqGraHpPvtCQdnLc3NeYFT9kkyyIy1zpCo2vtfXMJ4j6az
9Ydsqo7f66vZI04ZpJGh/oqGQqh8Fuw8nmmTu2ONuxUOrPsdY0d2lzjD8PJ3K/Mb
915mecamYGk34VcF8Dy7DLWcubtG30/rgkjn5pVQNBH78Orx6JXZzfbieW3O9JNJ
iIwMJa5lGiqq3JPU3LXyBm4uXG3AuwjoqfmuZ8T0yVRMCbDrZnzXx13SxWS0dMbV
vxI9OqLglJAvKcsl8ETNlbN2usWpkXHohVQ11NNaCuWbqAYRajIF/v5tmtJ+m7Ic
+ALMPQv1Pca/DgeqF47MhacOcHf5E9Oyltz0CflfY40NlPcTfYm2ttMSatgAJfDA
Jrdmb0yjoklnxbS7lUmCEOUIPLXgj8pvkRtJ6MhYo/ridACy+V+F+kIULUVNl6oX
i+99mS4KLj8IRi7rFZHvc+RkjZBAWaa3KNQI46OVQnIOWuGVfTzczv9hb3FGmope
UVKmlBE/qMtgCVLgdLvcdwNGg0K9YNboanXqNnkSsyaHG/8hK+I8YRxy1mSzoR5H
OgRL+WmV2Zi69qG5PLdka8NeBNixX72mzEckaU6WkK3+bF4ytWMMFUd2YzErDO48
gbcNqb6Q4VDyFv9GEf0gV2QSDEEdD+6/2bLV+Xksse+lkJJnTgHnInOYKLwRA5zu
aIk6YtG2ev6GQDjEHBlFNY0vkYbEe7Diw9YRDFETKdYl0662LGRsBpd9KO3GYoT/
s/09dhmoAyoyZA1CZEArAAu/szuwvZYPhf51Tds6kwjskVQ6BR6TKktq+KUv3svG
Fgz6d2FaL4CiUUblWY+02eW8LpV9PbpPJU3tOdeYYJ0BSB3Tj+5Oi14067vf3/cB
gQpCKT5C24UJoz3dynk+GeJkcrKbcoPePlellA3u9r/q/EJAkKnWHjXyMyK6A6Aj
n93EBwteu5HScf2iEHCpuDpLjnyJEPgES2QFZB1uwIjrvApoHN1jeyTiycOHl5hU
r6U0v/vTko/W+8SkQ1CrVBqVo7lEcZIojAEo1nj9/tInxMGsMFZ5FQOtTKP6yuGn
qpy/T8DY/py1xLPhIrm81fnm3XZBAI07/EKg2Z9ID2qHfpjZ5eGmq7m6D561mX9w
gj4PS7AAHtMGGockAFP0KrCki9PMR5Um+buaj/EpQqnTso/WUyAQCTFdICj519l1
knPN40ZlYgiYHSj+6mUEzacAgc9os11lZGiwgKHnnLn5cNiwyPTeaqXIr7rtVvW+
F7Zy3Qm29GeMaWPfJBHBvr0Y4ABCO6CR6KNukfAP/JLsszUHlq66zFLoC54cLxez
K+QTWGeen6aYQp/eGW5W9GI2TutGepgEOZHpE7WRUu5Pe5g7ps17nkuMkoBWL0XR
KCqJlgHDqGJYb1iYgDKXEZpXEVf/B8W2jdEZGnRATDsZvWgXBGV3EZqFneXk07uo
flm5gHQpRnmHpsyd3rAJU1r0WqBzlPIOTe9GLnPznIMV9A1/6xK4+PCMPfHhz+IG
jAtC/npWptGV5zDNRNaqTHGfozaps2oiSWo/DBZRnnBb1qcC59AoDMC1SQ0cuyAm
EfshbvMeCmwDK1syhxciMA6WTh4YN243MFYqT4NYK3c1hxOPtfq0oNbPfVU/o+zx
bKiG1JKwSh80wyRvJ5mNM9wsButS1tG/m7VPaxocQyKqxbpAqS/6XH7RdEs7roLF
l5WJq4imFK/Fc4sSGRUD5KmZmgYKTcVk5xMtlwXcNblKEEDSstBz/Z08KH21YuVy
RGP9cpEIBaI2WdjAt2afnJO6jSYZMitYWy1AWVzTEmIN7rnRhTxvAcY58rxgfHV4
aFIpayJCCWmOpFRSeNSCQUe2s5LU2YB1wmJjsCIEWex+9ltrbWuDM+VPGMs6w4vm
j3m2rHLua/iBccE1hVlUeNeJBGac9PyDqODZM32MkuR8HHIevqmPnMk1VM1Rax5j
Mnm8vA0Osk1TtIMh0YzP3ZVgQEo30g6iJF10KK4swZKy8264ImCoc+xsIVU/smch
sMmSGVMWwyP9pcxsaIQQAsDkwtBFEf9NDonwqGRDvuZv109eZq/FG83Ri8Cio7NO
dTehCEOg5ONy92XSjejc+PZtWI+6pQ/cf89LnhPSUY0I+no6uLgk3OXmFINkc8KU
6BT2/quhT+n9zhPtlLFMtkmD3TltgAIbWdC63u3VxgLGBxg37qfzZJQR+sImD+GR
YGPised1RWyr5IpAsZ3tiAqzlDsHCEuIG7BjUoEik28JpKDl7YVqtc3zcTAPZ9GP
/JHgHrjkhULdmBWgfFwwq6s0xJ06nsVja98h0cZ7JGUH489Ob8q8Je1VRlp5lbR/
8XLTMISbdGaaNKzyixRhavBTDELyrru4uOmewdD0GRiJq1L8KWHTEM+Td52aHd1m
FghkKS2lSn9Sbase2uXyk7W5Urijz9gZ1qxqNY9rTIViA52nr5EHXLzFqXH2rDZH
8I0ztmqL+vjoqZuMThCmSVCd+O02VfHPNLLvfAGEBFr8VoqMCajDdzo81KNRHrfW
9qTtgTF2h715ns9BGyO3nN/rajExEI5K4NHr+UOAWCKLQZun56dG8wuQEyvjNiHy
6QUnFge/yaqlAZSz4AwH+Bn2ANqxQPCcG6qhAIWn2nySUlxMB3ELjT7edhaC9J3b
QmfiGEFx4rAJxXp9wOAXnSv1+4xI/ooFo15xH1X/lq//oOXpU2BGwk7fqGOHFmGi
HbC8bHhG5vU22zIx/zFlAY1PwrUHL0yMg6X8aw21RlEu++fPjosf0RH6+7z/T7nt
8i23vVZl7QtmulxWr8M6kuoguxXMgVL7yYYP40O236AvIC86RBPP8M+1tLnVsFZI
8D9+QiQPAFrfIZL5ot7zAI23O1q5MJw9UMOl9R9GHM1BocV1SET7BYYY01XQurOP
gF3FPZ8o/eMGB31ZNJvtoNAqrKQ5ihSH9reYP8N3iGudz7PPUOl6xlspNv+pROHx
IFC23BkNDTqmpZKOuR4vMpo6ZdvV2iECz8E8iiP05hNRhXsHN6rYkJwVdbnIbIU/
fl0c9cQcDghM7o9nAdPZLnj4Q0DvIHzvPSAi026pVsl3M2yHEvM9JCydXm7rxXbZ
rEkPkx4QZ6gPE9nBctTBdjYgGvsGdOFMqzskXazbx9EKuLnTlj7aF08BcVzSMU5D
aGY8XQ7tmzBy81iGtqOeNPR14XJq/FgO7BBNmOxgRlbcQZElyQviknntLtb5DcVO
QVQDLGSPumpWxB5BFhNQoAbqdt6N8RCeZZf2VqJLZlOrBnJmUMJ+TNE9/NzJYe3J
0QjSwSQyjnIr8oDCoPA2l5X05hgiD5/JI/ipWkGUxE9gB93en+qmQb56ZMTmUw2z
389Xs7CeFMRGlNyMKiysMSVmDwjxW299L2DR5q75uKPZFTqJewLDu/myckiQBuHD
eYUP7fJmvsl7BdUsap+zMLxIYDiXudxcd5TZsvri6CqW5rLUIKS8Oq1J2xfUFO8h
xCBvl5BhibbZwfw4MySCWMX9sXodmXdelORBgCMXH06NPtmEnJMd2PDbcEaJVCup
4TKWGrTkUpeNU9Mj2fkCVqIGhH60SWR88/MHiDtuBMwzVqkG9BBnqvi1CPXdBI5d
7B+lQ76FO4qfvi8qnjAtu/fH9Vs6xFqQyndYpl2lDPCd6GOACnQG49nfdXsIGtG4
KUzP7DtUhSEStCP8DH/SF1C+yLA/XAv2i0xjkNlcRG79kUqqreUZjqLcsKHGXOP0
rukRP643zOJPhoYmj/Xw43l6ZZxHpaFzQA9bwkub15DTWzfdFEbs2ZBiaRDa1Jc5
YHSH8GeWtlHy+eTwSJike/HncD9mo4Wm/b2Cq5imQ2HDXXDzdlrHNDvfTPQNxnet
2NttfjHUBiK4S6c5eRzilcVzo66c7Tye1YtaeqN4iQ5kbuI3XqP3AhszbpSajM+8
4dsB5f5nh4JkgIvpOjIOn8sO1TXNz4RVyF/EkxhfNcJzmH07CPkqQxQ+O1NcEC9d
hQluJNhHxJ6+A51CyrrYtoVXdfu2RzI8fZp420HmFMArXrMDL6EqVqetmDoXDPn2
ZWHWyL7aY5VLGroHfD2Oc8pccARowzAThWdrcurrFy2HUMJgsyLKS6md8GkFJrlQ
hvVrhg4b5nrNRt6wk+s8ZLsBRrUBbJJRyghg3rJodPPNaZ7tQiR7hc2F5AwZXm8H
3xNcPWSrN7KHihlzh5IsLlSfFYvuzuZWvcILTjjBGvE4Wg5BjyQLuV/IFLD+RoiP
DojYV2TuTAqU2jU32d5v++Q/o7g3FaXQNLdW7+Os0/6Dcuc1SOYPHmh62Zwk+FsK
yWJpzpNCn4qi6CZsojDaNJ2Xm/Nhr/yHdfiC0rXf+qWTpw4z6xSREk9i7qxMs9Ww
ozMK8viUw1Iw+RRr9NZQuIWlSaztGtuiC2wdnaufnEn1gI36MeLKrg5uFSOVwieN
pUk/RS68L0B5DhnJAP+pYFxmFBh/ddEE5Eiz6oX2DfOm5QEYvS0hBMQnsmHmNTbq
iNB2H2VUkge9dCZFk+zgVL5OJDUN4BQYGb37K2ibSk6N8pqec1QySdk/pCMoJ0NX
hJPFuO54OOS+VDpBmqCXDluRYvgReTeEz75ozbAi9ukxUvLYg7PyiTB2xou6C6Vs
o9/raoMffBtmczGoeGAvrd1ws9dD9JI2JsGlKzILxcKDkoVQRh1W6Civk9CoNhxC
p6CW1EwyEWt8vbJmeD/6ACkPuwfi6NhzpjKYpnTCeuLQaOmwKvgmDashZqACREF8
owEDx+6/DDaMNOn1bRSFM0j6iT1fcHEQEM8TERzpSGxX6vKMtPESLHUoyaDPkysL
A82g9RABZ6c8xSPA2fUw8jvZMTEh5QhAFzPJslpoRC9SNWfRk8iJ0xY0fXSlGK8D
NVj13xoJTWJCBad1/JZJgFa4a4EGSUTm7HlHcGOWIONKxKzR5w4k1G3KAYPIqby/
C7y1RxteYPUBxSWYgVu4pAp7z2QfdQJk7WXsbgdJj6eaUQEfjR5hmWzc1+yK0y+i
mmABoV1k6g4wcN8fj72k0tp8ikJBt8V61vw0I3gJLV7U/3+tJzNvHUxG/lKCxFhj
+8+6enrTsyAqrO31W0l027/Fiu69D63s5i/ni2XeSjxBN2KU9Ohah1osvtUfrSqw
7tZEH2aRjtX1pNBQzaBGtwCGREz5b/WHYnXXaJ8L7dSkf5IchdyhmiLATRvUKqe7
49yj2fZMWryvvyw+E3CgrgEUCLk4y7qCR9w3CFDyefLuMPjhyfC5U+/ErwQzJozE
eOYTSCwTtB9xFCcFwcU4FIOPZDIACBPiUVW3IQI7+K7juMDG49VMqE2LufaL99IT
2AA4yZHHavmoiC8axqLJqROQe9MWyuWbPk9Vg2lL9SYZmS3wJG2/ds8HDleP4chN
ZziSFni4g4F3ALMkSMXGZe5oZBPbQA6neLtB99r7eFrRmEIWuQxifoJfWO3cUy+O
/1ZKd//3rFyMKnUWosSeI40RoI1xJOzu4tYWpEGNGkRG4xMx+Ps0H/Nrn6pIDqhs
151DpyMv/PCfOivywZlkrkXHQ0UFoQPg4M8dpRg68r1bTb+Ss6NUTcf+NdaSu/Sd
l6TW3Mx4+MeQs5LwmVeutPqzuoOkEwr8ByScMkz0flDomG3XztBNk1Hdxsl0cJk3
iIuzEDSpnaMu+izdZtHMynLj2tfFZneF8kjMlmxggByJEKSuGdfvxCFuHROZhHIx
NLO8ykn3R9vNZg7N00Owq/BVllMLG165yCfo3Tp6bA6Uls0fBSGos9S5a0yH9SuB
weK5rAsmcIPFCEIYAxTNk/+yjUPpcmZL2odKAxLGNjIdB3lUHrZbmxktN5EanZKp
6tgWcHgRyNXgZ1V30oggmmk2YwAaXi/Xh4jSc+Qks6TDsswu31YuOBPmg3XQAnSl
E5TavSu8yltOdPMhTDLWvsMmc38h+cfAuBCfO0xBLP1NCl3duK6O1jWAddj08POs
YI0tVGFT8K3Of2JPOHXFZsTU4JW3IGY4cuZRKZ5keqqIeyuC2Xw59gTioC60d+XJ
lV3APgfICI1kPVNe8i7cZ90yNhcH6OZNOCW5WiN7HfdTyeFYi4DhHGXc//JXHL5N
ZsNqcfRyrxf2hE5PmUbp8RhI6piMfV2DluC9ZJdFRZG/aQO4H15LrXvnrc2ONgP/
JAuuZjh0eIVYcjtLxwDccVmozSyvXJZ/3dbm3ufrpshTbsius8fUs4Wsvpaykln1
lbA36wQCcw28W2MqB0FdndBw6HVpZ33KmSyDoMlJli0zs9Ve3yRXYxgDgfC8dwpc
VsG/vkTCg/tXeVIdzkm3ZqW4PZ/tzx4oT5mfCDu4tDcMnwbH8vA5qH8QwV/P75o5
BmKTxQp9+r0jg1Krh2KPjXKmZu2WHt6Z/tPZ8GGS1k9NKaBL96dnX+JVAaFr8zyY
4/ApZCDHU3qcGJp2am2o7SHxxW+F0vuXstOqN/UfjTDlEbGUEjlI0kuOCD7wChEv
Rqycm6adCiIAYT5BA0SZkclUr9Cz4xqFgAzmFhPPbq99NsmTmsTT/xsVRvgfkm33
PlR7v19BZUK6Kqg5IQeXXtPCBitl4VN5IebNKTMP1POF5ROKfVEpXpX7Ukg6xjz0
+xdlzYd/fYahFABYmIPS0n/M1J29DHKBbQr+VnBqtOBM+CS5O04U/ZN9l+YPM5cX
k2WXuhEtvvKt3R3rf4nwdN3+KAgvdhop7b7tIE+L8DaM4pu97ToruTCiJNbKLZnf
ct515X5vx4vrrXoJFz/eVS7t0lO1awPbbLfgjVSoBECNZtzFkUULAH3M2laWWYZD
/CKlbSfuCN23IW98xd3D399sEp+4B6p0ifU+zjh1qyWvRJs97g5kYatLw+daPhXp
7KG+st8sWI5rxpL8Vc2IP/P5tDbfPwVM+q1HQJvityqM3AzRz5/9ESHjpk+E7zKo
VfEgrRNPN3NW43WZTpaCmdXhlwE9zY0w4oeO8ul39kmZfKrBsgAUb4PM46EVq/Jk
P03NuRg3gm+KLIFSPqXoYn7UiZ+v714AYUQJEww2RN0Jbfkpe4Fskiduude8EhGs
BKWT7ZZtNvqnzXVt8SQZp1Fkn7A+U94RnJmTPtURLv9qg7EUopUgSADD60Lpz5VF
CNaWqvD64qlBT/S5UCORxZGURYzjl1oq94xe/dFR3VEJfCoNNXHq0ixI3i1Udrs/
ugYg+HPkqfGmI7p55Gg1khX05WO5w2I06616jcMesV19k32300UoGZSt4UA+R+M4
x/I7w3+38CRcEzA0BbwkvKQuqY+ustMTxbv9kDzA9KDlSK1PSunbiz/Iz8msIpEC
Vu5A3smGW6SMogL8wYHNt9RW+ChhXsy1j0k3BzmSDqtT95FStWdVhmtyQEkuCjgQ
KVHMhLdfhFOjPF2qjnF38wp3MwdJ7hLVoYl91sIFFe/rFkfKN1AJKwN8SBS5gF9I
WcRbdfs8rr7cW3ZoUvJxn6vNVShGyo5qcbp7i7cnsbWIHvEajLiJEmrelz77Blu8
JcugfMT7uZLtcwv4xXPeueMPfFMYbRYbK/RQiFfz7Y0VWDNFAK1F4h3j/JfTVl4Z
mTl5PwSROfYETYoV8jjH990Z7HCZgnmvJlPisbAmUw79nsEPhltAD2/JUSwjXwyh
0bepIwdaU7mSRA3yd1zpnCcxVVQzndQfQSsiNqqJsTcXvgKdw2zQXT6zcK3YmSHA
a4LKxKvRbfUXijScw3saye++wUHqs2ArDAuW7VyoCuDunWua0eH90aD97nT8T4MH
3wxjVJrOa1C6ru9lnFIfdihp7P6EDZYuzlpU3bZvfUe5MapNFtog+FD0Q2TyEAND
Or44Zq4Owan57XO5MrkYeAkb87ny5GZS/j5Koe4erYqtZhwXUAOSAh/x1pP2ikne
L+lyf9GE9UGODVv67cVjeHnX/TkwigfChzDh1l7OeGMSZ1WxoTqP/HoiD8X+YDyJ
/fsnxjLoCTnixL7ajuHEMsEvnsrdDdp9BFNlFWurZd7N+nw1H6DNSXzKXsZcZxq5
DKYsMxZ3m104+q6MgOUsgKmPIpjAfbHWTDJCaa9brUPMEGHSsJv+YZmhPSspG2zq
AIaBOGbnnAoba8ojK2GldFDJmzy7770KSBorNrwrXA4rBh4NUPQi1XZTjY0nmii9
jdQc6E/VGAJbyMYjIGL/m8zlTaJbWhbuh90CCucyFBV95PMNASSJcmJR2953D76h
KYNKJ0YzGtfbFPtP2t0gpyg2mmo5If6FkqREfGi6ApAlQijgHvYaY3cDkz4URhM2
Mf1IT6YxSQq/jzoj5+3nY56SByZAheru+/XXcIprbeqhks0BCx9qjUqqCYfpPEyL
8NEXz87Tnwd1ss1lk2zhlsxVZ0P8Vl9Wd/g9pvtkNXsmh3VYv0OHesxBHwfgBxWk
ms5OkmNrX4wNx3yQsOHNNENrfH6d/EobXVLU38YLW2Gc74GCIxpjY4N+hBN712pK
XLtqsXgpfqM//5CfbwxRUWh3J0LY4GWKosKo0INVjAzKVgpECgMn2x1PkrHPvL2A
se3JLH1YKmjmu2Ngz3BwvDIRZ6eSdrlxNrBesK4lIQP3Hyg3wAKP+4yCeb88lRdd
HkqqQtSvfYoXtdYilCtpRJijBYCkCTDgeixSvybKC/Q/RBlkJlECoYm4nLPJh9DV
SxA+36XhqrWqHdCvYhViCeXNm78vKCthCYIDogrid9EDWEZK2VMeZsm/P7iilpCt
BBfZIMCVoI+VF+v+Nukl0ZpK3t8/uKeZm+Yc7v/o0ksjz4OLg+hMbkDQzcXVIQmu
609Q2UWVZMbiR0Wv1K1xSZpGc2idTyxTJ68DKMXKcysAvSQD7CLl12zAKsHtYri9
1XJRG1Oh6ryVIXz+iisoxUFGuPv8TnrRRvY4stbrCm2LfS7F9Ye2ocSBZNqgrXgd
hoQtvYDHK0XLnDNgSUzu34Qoi2x0N/MmHozZeevplQmIN81LFcFcX+kC8TUt/weL
sz/C0x8cCCKDiM7SEMcGQbOQ7oTR2vwPbeHf1YKxkWeA4WTW/oVo7AgQWXLYQ0Mo
pTnuGc8LeHyG1vDcQL0s+l5h2GPqJDw0I/akMFa86ym+uI7ELAZZPSEBOq5Q1Ewq
y8/QDCz/yheNUi4ItdeBuBaLyt+7CuMc5wwGLN6FuegHnucE/xym9CwGMKn7TNoP
VwgetGJMzdTLNbAuxsg02R16DoyX3Rj7hqjUrym8+fjyRgsouCAaTdayhdL5KcfN
f+Pg4Xl6d91hESjIeutKIOwJxe+JWcu9bfAyx1v9eAbZmakr/RFFM9nxRGmdexPR
EoI+ejajXk2r87YLsOAEk+Y2Bd/HUbWRw77QegHmvF6L+rcCLqWv5Ht/6dCqAwPP
TTFzPdGh1E/bRICtYvpa7mUn5ytUcyGr5JaMER3F33B/SrxxqNwlTVi0X+d+fKa8
Rqw3STVMphTxrrpZjWozJ4ZSrZWNdUA034w5ym0UnIWUFVyPh5TuB3WCzOfhqr9+
73cjtnuW475FgdLkILIAKRGop+TvYoO8HTPKvcCHCVHg2mA8Y41wvSYVFhPWEr9B
gySoplwmrNVkTawVP1KaB5u3fU5GkPCdcQ7vsw5aYX98Q1Cveyowta7EgwHRctcI
0vsFqNbTX90iL26wr78vMbXc8Jm6gObvmtHfZ/T8aq+gSyycH/XIeU4JVHOHfHpe
65WCHPKqLHV5lSybxdkBNo3Ou7GGT+YxSo9MGe3Q/4pHo/3txJfhPAFOpDAxd769
WsdBsAcy2q3lADhr3d3KAa8HRTbAs2XPR5yOwUseDRUZOO4Wf0gpGXLWOY5fB8Ry
Ts/m9HgAfRr58077hTwv387FVRS/AF1sVKJz4nTKCSsk2RgQnQsbUqtgMTPx5R/4
c9g2flJ0wqT98xAqOZCCMX7jklcki5qSIFFdxCMoD9cWtEAGkxjeJIT9or0BJ87b
FOTtIVtxoyrLhn5RIilBMKWYiNMVH9W1jsfYdM5i0T2shoPORNU+MBcADf/Ueodt
EJV/rmCPaGWbnRn+9ew4QoRm0XnYEpSaZwBEEsyTzPZ3OPb+jFh8dO4unMxU95j/
jWgUiokSkHBVUIqbbBw3pqjoilCvPZmumxc0Eji1DEbdy8Zv0Qmkeq5iv/N/igIl
nibvBhtbmQg59C3Vvo8q3/5DXQUsqjXRMSV561V3cevm/i/KL5AH62gJM8c2InSI
QEsUHu5+TGMEzNgIhy2ZxtGkmlRYZmwLVHhBsiCV6Jji48Q6nsE97uKi6z/RwgVZ
7MrthJpeX1bj8OkCm41rJeghRtk56lPAu5wGjkaXzzEwMGNJyLJArWKk+MRIc+y+
+bcBCDb8ZqVj4ZB2QItSnVV1U1sLpn0pMOa35SNe24ooDHIdmVthKM7aiNPWoFAu
3efbBbXNFqVt83qiAWgwbvVUNxK0iKH7ZjXQlBKDqD/EonE+XQu+mffS1SDTAC/T
R7NO2s3xnS0lGs5lbomEoSfcFO3MhiSHmx33o4pXb6G2YXeDGpqPqSKas9KZ+d5p
+FqqioGAv/XaUgNHRfH1k8QjO0o4n9ZF3dDaBc7qdGJqJmV+1/LUITv2Hb9hHTtI
2jY5gaGZ8l5EsP6Aw8SJnfP6bE1NqkC4PNNlG1L5bTBrlgoBsEWyKgpJpdQJ9IP3
AMQyZ8h/PczF0o/Pvwe2uJksKIw5ZOjoL9wR6kBPkAZDFR6DMRX7ajvZHvl9C+l5
FZz1kRnHpRNsROGEuUp1WblKskvm8KJ9cw9riivBOA4TvRn3AALfWMTIw3XJsZAR
vaQwK42TlExPV3AcDX1KTJzDwIr4NKpb29wUWM9y6n+3bmw3gkQv+gw0vIlKojsR
wTVKMs4bLAIpg+TGC5AY4r4DvoRJgQhgWyjU/q1sFLVUwgeL4+Y+VEi8eto0Mhts
e95evudbBeZDsGRshMuENtGMDZy6uBSyDBIKuxLufcM08ACjneBP9l3mzjjUkQwX
PafKjpMZoo+ivRy4pREdv27BBmwqaRir9lN8Y6ho505JSr9pnt8/FL2vL6Y1Yeea
BG9b1+k4ZQKyG6ef+POpWSR1RtcwDtc8XhmTU6zScXztTVb12NYpaKxHggoUm6Fr
/H68nMkoreNy+uyEt46ssixwENK46soI5jH2/5uxe+4cW3h281twcPD+1puYYMQR
I23YAQamGVfKmT+dQ+gDO0F4m8aNWZTR3xZ3PX5ubdqxM66DqGWPMjao1I6fDtbK
3GP0d307fttBWzavIcZfBtM//hCNi9uyALuXbO3+hhvWY3Lp5vsJNptS+kA5QwEK
vKNbW3C4k2XBcvIdJ378muc/wv2JoZVjRvMRDTI2DxIgX9g7ryY5Vp3Bklak7Rfq
CvhBl9i1MQBqiTJ+ZI6sfTlXVHxsfJ/YoVunNI3X9VJ1R8luS80WzbY0R8bZ3qsT
A85lsQOMJxJXJoXXiHMjjeMBKUhYqWfqZMlsUGSR+y6U6etnHOuMeJQep/W9PTrI
fte7v13yqG1obiquwEDdXO+ZR2aFhC7nXCm4kCsXOdvSkRAetZ9hmOZcvXMlfmrG
LcoFPtbd0zmdauQZ98s3aJdTFglYxlwEfo2Xg8PCXsgdcd/Pf9vRkbaR5NaQKCny
d2+jRh7zmx+HW/n9cV89dwQB2hy6WHJejMu6KpRuqmAXnjuA8XI2Db19v0OQ7LZY
SNcrpawxb6my2Zhhrg0ofybi6UcbxnL5F8g53AntKvYjJh+Sq2MraO3wW9L0k8LI
aFs9C3FDwapUO2ellYcg20nGZvredVfSs3RhwY7085oV3/mEdCPixL7p65hnvmbL
1Tkd7tOEUv2mrJvQnsfQBbGmPDLj6kNSFd27XbYwu/oQruhBtI2qVbVQy3i73831
tVUo8suQ4A0eIDvjYI0ee8afofGDlOOFceq0cwEtyghOHxg0wJXGadOlFhXYBIqO
2FqxvOwgMKdUDD4E84zUbExEte8jjk/lKAq3TQycsmx43EqNZo83PPTfbWlXyG0u
ZgFRCp7Yd6C/NE2sceZykCcLwRFua7mf9h87WybZ/lvL2kupl45jMmhzoL5Ld5SF
DMtkMo41Lb2IaVv1X2RuWrsk2yNeITxf3n0C2gvlFWsZahpYLEg13mVtIpB0wO/J
CfjBT7HWodJpUGqfTv8//7J/L1OSoj1vnoysdhdHPzD5qUZMVsKF7jVl7MyYu5PP
OYxJn5DYQHJeUghGfFXKN5Sq6NF1tAMJx1wXpfO5GR9Fs8C8BghxAsqdGpOcYY3i
tAp94SZLWWHG6+e4WFrxOETFlQ9p251YEyBxfDyotL2Xkjy1KqtJnm/XfhDh2DYD
iqTPVvoyj/VAdD0KJuYrZhlqDs3+Ix98NlwsWanuH2BYWITw4UzstwcaUSs//W7w
OEQRdul142MUw5TvpjWv1nDa+FH4yZ57mXVQWPHl+iLoEgTWRELUfG7lKRxo4zW4
yJthz8kgEyx/WBDjS9CV/dQjC9Xi+9XJUPBDZ2S8A3WFLGKxp5oSjV6HSJYRrAZX
wYxUZI2NdD8z6Ol/rwzSLd0nK6MxhbhJbPk/+DiUWfQlf+5yGW8hMOyaxpbz/mIj
Sdj698MxtUt42a1fFfpZaOo+dZPbZZl4ZNajVELHUYe6kp3GRmk2AvtCaJgq8P/r
vrvzRBxmjavW7VVIxYFsPQTi3M8SxBDugiIHGwIioDDouAlPK2VD4V3AvRezAZwy
FEsCPS6sN0HVZL69BMbBV+zkOujXXhwh4/WohlwQZqPrINWjYP6U+bpPqKUXQbZn
D/kAnaje2MjXZB6XGYnc77920kqntGcfBwnP2eIBdTT9D2yBwyMfLTU3/ZKLqKlb
Cc+ciXwhHW++C6Cy+PtzLuNKXHmNVAlZfrCnvOQanoacNdhQMgqsO9k4HjPZ5llm
L6okWVP+aAzse/ltCffP37MwiYyHqdBNGDyNyKpgvSZcq6qlHJNOhONNbVsrlaFY
7X2Qj0oXAgBCuX0qRDNDfw3+Rs7tOMdKKw53zKftUwX09Huv+PqzrbOfPqQQJ3gt
PRQulfk6hB/AqVeQsxDEaxoHao6v66OmbwY3kd4K7Ld5TLiGm43cAfHJ6ygmFmnO
TSaics1S7AUxTtsLNh+gs+L3WYPoLhze7Anq47CziZao7iWKEZosb0VTKzFsgE2V
eQA5rA80jm4VOqAQVCFp7W2Qnx2BobEqZuD+yQPFYJCQcJwr/68DbWCDXN2JtU4Y
8DXN2eAWcRuMve93HC+qarbG1/qI/yUQ2ZOgf5Gxs8dR/jZUXz7kcRnp98s7tU9S
6uvoc2n9eAEzoPVCsEGTOn3CDUTg5Bn5QIZD+2b93pUe6QA9i/ZyH3AUE53bukCR
olB5ZIJZX3m7vn4zyKCQ5pw9zEe9Y7RT1xnExk7tR5gF8GL74SSJ+DJVVhxHGYGu
W+iW93E1pW5Bms20+INiX1AF2VjNEGPqbmIOvOZExyvPI93PpHz7J/JZ3waBjo7d
q0aPLqkZvEH+xTXZF0qvgTLrE0eNfan6Hm8H9RNSHqSUkXYV8QhWIRkzEV49X1x3
uzWR0zJOSw/y5Vif/RC4ewxG2UHdNwdDwnQ6p9ECofJccGmwJSBFL8T9v6ALb4di
MzqX30ymg21HreX83/ZbIaSc3IBW/GYDMOnZts0ujiaetvuj6lG9lxJ8EnudPH6E
AXkCPGqse2wR8SnChTFVjceNlwQu4wQ2aMFYuL9detYbkY/Rw+UkR5p6Ws3W/CCS
R7c1h+CmUu9KWGVkCK5SO+6bXNC0DMXrLwyfEO8O6gfHfdVg2aK5Z33e6enkeBwT
RGSxrYPjTNbJzUOMBbppqQGg7ycUnqxgSGtOG5fFgp8g3y7wPz5k9uRYTAWWrXb9
3w6prI5Po/c47q9hLv2VVu9qt77pTrbPLvvvm+6TqDavGs9C2PZANxGG/l/8IYKG
6/vnTDgkksn9xvE+D+eDvxafl+hQQvjQFxa3je6Ml45M4jD6i+wAXqSEKTE6Q0ak
V9BLgD7A9MwwX24DDCVWo3DzB3R6yHD3JI+KTh17Iytm1gQhjFDXDN1Q7yfslN6e
5l8Gr9WDXa1Xe4bTVryItnIhoA26wU1MRDkamUKQI9zd1iaEXCi6M2k1ytvSFrol
5KQ6ZB69ymZaz3rE8ytfFJRuBvl5+zfNnCebJK0P4hJ31zWEbbkBXGrTKH0neLW8
JnUd6FyWuMrNBf2ddGofr3XFsrlv8bIKR3uREChvXyb6HNV1D1WmNoFXYyqCMANb
mQBpMv7/vjOnhxtBU5kcOXRm5Im7wDToO/nBxt/1mRmXoN1kSalLkZey4AfHeqlJ
NXZEUcXL0tsQxvzkwhlEqrMF5eBXriy7TvvU5il5HvmkhcDfh+7dZUd73Uo6gG57
o7i2hTm1W7vkq9V0Ye5CgxpdXNLfXBBVKDD7oUoluh+p9rgsPrCVHGlphnBGqG/J
ew7mKYKkshq69MA1gQrY1xPsmb1SfRqjCM6W4hKw6yPD170Ed0sD/0+rscZW5PNn
ZpiKCFeW+a/QktW/2rmOAmmPA/Yp5FX+jp/EuQ8djBXAS4L1IKl7qoIlu18Go8wD
l/cVndjXRGX3PBKF64rmp4gg8A0qd65tvmu9XrFlo5XESBaVZ0YY/qvKgn07msJ1
sKcfXLdxVP41t98HHOyl8mu4LmeKP6PKMlZaFhhUWeiE4l4fKWa8SPOR9QvFvBAF
Dow/Xlvdsu1AE0O4/PQn6GSB2ngSzdReffTI2TsmnM0JqCVXWBpJK+FP95okY0Xm
yuLVXdfwELwwGFJsTRAg6996rkgAweEh0HJpIZ3BtY1mwyiGokJDJODYFkp4V1+W
b8vLF+Gz5Ty8eMr+Wl05lNj2KGqMYR1XINHxflbjliwz7SP3k3NrQ8ln3uQ/wNzB
D5mfaxRynAuXq75tkfKo4UU/f9NZntohuLO5fb8Xper03NuWa318KV8QLn4WZB9J
vk6OaGxWGINTC69W0/lyMK5B8r3q92+Zbkhjfah3wEVa5HYvRdqVAvZ1I0BbQhSC
gQvpNzjaRHqz+MqT5tWLLpTKCmgl4oPCymv3BEQ5BqUh3CJ3SxMiZgaV3W1ewloK
9Sc4zo38WKyleX8OKmSG2kQTY2mhNs5caQa/PBeLz/K0jzlZRPUGd/rl9kq75ncm
xu9/dhVU6o9dz9jvhrivvNtBJMsC5znAAdDgoZkot0UdUyK9E3b1TC5USqy/cuyK
Ijpe1tPxHm3R6XB3yFVmpfWpk0V7sXHcOz0PRmqxB6QU1IS4z0z1drn+UoyvN5VI
KEXyX9zPSc0MUMhKQwDHDRO8moe0OIHlrL/C5GeLlqIx0og3Z/v2UEs+tfjQ5IKi
ZSCiCeKNwCwOy1k2J4VGH09T1HnDzW/pOSZMbdK593vtwb/4Bft10mMD1XKUPMyn
jF3q52MR3ctzDGTBIYezZU9+NfeIKRpv8wiGwXP1XakZfoOOOLqNSzE/Z8q2RZyn
WjaXnH3S9AwJiCbNiajllx0LW5kn87P+2xTQgAG5lLCMoO9N4U4ttapMpz+n4Ule
T303p+i5LdcRoA/pStPpiIk+os2qfgCgdE0K2fT7mo4Z6RHePzPSngxdgENOMHtz
H5cSyLgbcodq4eXG2hsCapdDL3koNcvUDpHjPwyTBYpd3fik1tRpbFEDdhkZUtgx
tJ2PiQmQBusXru96XRfBSHGH+spukRIBm1jt7kIZK8T7e068YVUwy7GYA3Ro5f2n
Bj+o1QMm3bn12ckwiYjX7FdETQJ8/IYTRGDcVXl23nvDW7MF/rL6UU4plfzrXd7y
y1PN9O2ZFd8LDHGr2oeZ8UeAWlfguMO2XSiMpKZiPYPIkgebyOLfn8bopEwqn3gd
XZz/GG5xqwj7KRMfVUGDxYcCphwnvyM0gin2B51kg/+JoTvbMFHm3dgZs3PqOROZ
+nx0NQlCq6/2LneAT3jWDdpbdBdW606VqrolVgxl39+NgIJS6xYsjgBEeLPuUdOQ
GSFxuuv7gvZMNFuCs7aCjrDu7N/6d+D43RD1GdrhkDjmXPRbE9msG1mZGhHJf4TK
TUaXdBJB9DTC1pVdRhKOe9BFkiZgZBk0GYMq4I6p7mYas1Cvqxf8dvhWs00PCm8J
aYh9jIPHXIpjxv9uenh8CQXGo7SOlGmdASFrjlEFaZx7fekSw6GWOBtDY4z/HS1K
he5lttPCKPHUo4lco02xoEv9OWL+AxRQS2bvFvV7AfMnHl316UWHxvwvnF/n2kvl
9FTRY1lfQnN+OJH7ihCTJlgLDRkp/upbJB81VCY9SMvNWICZpwCT12B82wH49ImJ
tJnJXdEUSCRVjBUDZ2097o9rMYQRT4F0KBcbSwMKDOkCk7i+aoNf0fuUxcL1DFdD
5s5FkQecVi2QnSLrKfhtA53h7HAkMIy25jkJrGh6wEQVXx8cXdke1LBtwXRdj73A
/RPzW2gTQYC250Az2wPTTNw6OaHeeSnl+mOMgZIBPEsofPAfRLYAhIqMHAwKBXsC
TdyMtz2u0gnqPvzVx8MTDyI/wUcojv6X35JstZp2jwjP/0eXrGfjVnthkocbsnIB
aZaK0mNJdu0Skj8TdzqX+vealizXO4w94C/PT/sN8gl+qq05vHMYHyul16aHNzJl
oUmg75sKr9P8oD1Fa63oE6aV0eNeK+KS6enMoHK2WJL/0vWBk5cNPoAespaOAbGC
EoQsVwR1VGdxnc9R6TgItXaUtv2qlxBfsY1MDeAzkikr6ndhmWohTFnX5soc7nCh
IWTKF6PEZD/w6u6QUgxF4YtXkOhSeJhvVuxgv0o6sbMvt+fh2cYzpEAfeLVekhNH
I65Va6gjzzEnamtDocQBXjl3VJZunzwI+VS9ZI+NVWK5e3mvxJZchH9YYXUXGuTA
vrgm0Zws3l76s7/cLP9UpsJqeWz6YiSJUJGZVhEv4LOApB3KEVbYB6dXPcInLJ6Q
YNMbMccNnY+JRwjgwP5JysJ3iCy1mBioyAFfBb5z+v/dg6aG3uYEgojsGzLdiGn9
mGjiy27nkIO9NOhvd8vU4QT6boZsA+L6w2B53RMqX4Gwpkff7YERfPsRjNsTaIYJ
LfFcFamZXDwu0ybEat0++ZhbztcsyE4ggZwfw1vQsDMUuML4d4wHwTwi6faZFzIm
vRLnzIy7cA8MR09AUYycOzniX8EEZDdbnTxXagzJlS1hzCVGZfp03w5t4kpwRE4d
1dOJZwsJzYTksVSA6xafsnueDKW0mI+JH5AGBGBPljjqWIhpcswiA0JB7jbVngkx
ROffxc7dIUEP5g9VXhAz/g254Y20umdZnBJD2SDWyHxaDh7V6/snxr4CZi1l8MTw
8bO2A974/w8d3osVDtvjIRWWnudCcbc3bUX+1xHj5Yi/wWad5WWU3vq8lLlixEkY
Q+ye1N+dRINPGuu7HXgUbbIhKk5dKqb/fu7fS099fg8P8VKlfdee+UqVI7+cJLLW
wwvISOefTvghHtZgcYNSNyd+8kE1N/RrmJlPp7Hk8Gojji4gWWGd+HstxUTaicJ1
YI+25q8aImWQ4ZpLvFfh7tFMByCrnBJI8WQvYJzuSa0sBY740NU564PDqVFfRBzT
EdTK3T7WVlJzY8YOFET0IqQLjGA+jlATrl6jWBzF6Dh4+fpnZk+v0wxXBKGOv12c
Xb+hhzq6b8o+tP8sgtT0l+366vFYjdEmOe+ar9HWBTehCwM3NUNJwW7Mm/Qlv0Tz
tFnq+HOU/IKjuauWlqxaTPWMlDPen5+5+Y6+DatSJ3yX+1Ya3hxG4E2LKhVM8/0M
ztqaF8zDd9I5koU9pSKe7tozOirrEWV3uy8KeGxer7XrhVwJpvsjq2Ub8KpcuE3u
zVavFQM5mi3IPdVkgEE1xF6XAs8ceZ+kUfzZDByEGR0jZoFMejKuiKpJOG/bbbaJ
n61BaKp8e34dEQ/Dacpz5q8RhWVpt4d7LM77XbAQWxLbQDWMiI28wPJptZ3FFWW2
VpQpA3hVpWcRKgNCfMVKOeVSgwul7PwSw0XLVVkfmRiDic6N6SsiTeIAPitcKQbL
wvY/vwT568HJ9yT583Q/7D0GGnV1xl6RzvpVClnzHERPQIE505b2ZRFDJvTjpFQY
sfdBJK3nC7RbUrYX9sL7aES8DKcXpknRkWcO1evNlof68u7uDpg4+n6VR8B34RXS
EHpPJnp2HoK3PIzXED/nR5a32fnuoI/Zv+XzcQnToLbEWN6NNRpnABKHmdN4Q3BW
218F5l9QE/mg5wPf7jFwVg7IIO62Dkx3vM8ecBlN+O4+CFeB3y5kaHMawVgDnPXa
wj4TcIVPhpfuENNu5iPmd1dkOa2PjTnPRQ9vUXH/bwhJvdg6ESGCGCkjgOXCDZh5
XSs+lGJT4U5GMFH49QUiXS7CzN8rTzvszeG/P8EJ4xiTjy2oftS6yK4NaOTOSKsf
D5g+mv/ci5MG+kDXB4qohQ45mJtu0t4bOfcZVE6cc3mtF7UAZ708eRan3sHk7GzJ
KMzhgV1uT6LDn/6ggvtY5fpG5e7bm9Q+/+d9I0cZKGcFT50kBZ7y0jlnu9Krp/8K
Q+b0HTDPV5R0K3jZ8WQNQEY10JCWsQYRFnX1N4s7s//sx71a3Ar0TU4pxTYRtP7p
5Dh7LjLHmvmRADCoI9I+A6LyYPSemEXvMP7b/XiraFRPoIZwjnS5t2nLu0OOxjgn
gfdnvkgbptY+dAF673jAeDtPBnqacq0bn+J1B7GMjWcW9xG3TyX7QDiHLqeFqZ1a
ncFbP+Qmxia27mJWH2aXKnIe9W6F0FoSdGAZ14Ffx4SIlicHIpEpS+bXhS3yWEez
BNd4YPm4u74TVDR5HNovIbvShycWTxypu7lwON80u8hduD7AOOuy8T06R+sU5mWb
uYa8rMPugqi1WVUiJYG1LK+ol9vlNiIsg7l7YR/K7mVajN9F22uzgC/A8ILG/siF
39CQBhu3UyfLd1RfxnS0Rn3aQMEhNFGkJeeMKFt3o8HI3CA/mEq+kY9Z/VuQAI2I
ixFEOduNv87KjuS3Smx99lBfaFIZxbEdQSTubZknEMWEvYg5FCeu3LiEYylGw5oz
7WUiPjsVpKxFavACVu+d38wZGlchAgCJ3IhASS+6fJwLxp59VbfFW2dCV+iAIn5x
0GwUWj+Z05XZhivTIWh5CIOt+e5mRf9eD9a3UHY6PM8UyMvCc+jQmrn92trVVWfI
6nqev8CbCl+O42O1AafNZ6LjcGn866m9cf9W3P/K4ac4VnVvZ2Zmny530g/O+cvs
Si/fQ+wf1ZKUvSjIrc1JE6DhPAISqU976jgqro8OVwf4DT9DFIy7jYgM3H7FVu+z
tSLGglJ9il0MRL1f6kKmMrp0UKvjMR5dsm8/X+I/Py43WWsEKeJLKlVyfovFKNhe
yzt45mS1OexFx4J0HLLIVfUfTpljyhCWOv1OH2ZikES2sAUwz/BU10QNhcwKdR2s
MITLiP7q5kB7ny4KBjgG60n9EF0JdKII8N2kc+UpM/zVSRtiKb6gdWgIN8GvQtLK
Gj3A1Y9UlufRQsQG9xrqF3iIsT7i3LAEwRMc8bcxW9N2Ve31PBx8pBUecAf4KgNk
7jPT++tf++MO42RkJJ3npUMA4KGC6NcmVp0NUfp5YEdPV6ifteqerHklROuSv2p/
F4u5p3N4sGIVtHtOZjuX+trJkUn9PdbRqDMXVQMCbg+eVlpBHUI0zY4EBYDmqEut
c84nQHvninmx8ly7jR2auK6rVM5wKh1D1wsdv/FrJEc15ugXrLLh9nMrOCixu49D
VvNEGhkKJhGyXUsprsSATWladWz5kJ0rLaxpY1T0XpkML8SQFXOtMTs3f/8/tXx3
Cx6THVcttNTpIM8J3YVmeVh292Ni7Ir8Y2WiL+ZPZOpps8mKr7SfwyCCX0jg0h0S
0SLOCFD5T9C4MneBAXbrJ1klJ611Aac4OyYljNChfzZ260rnLOGoJewmkKpJkEBw
h4//QFmgheNQAo9AN5+ZmLuplXL53lGTmn8rl7tpuo41R7OVbZWBgv9Yp/5NYP2l
CVrXb4OKRE7JEHbGh7yiRBZuXpj2jc7iEXl0iPT6teZnYWd0QR8dGHdWbG3D/Ml5
O6ybp3maWtA+orHR/caPSDZTW14fpTKp4vxRJSdVlPIggfvQJ2VWSxKpL0p/uMcP
aEjl1sU27h89tNR2VCOr0rpNqRQZsNgYX2TA55Sok1RZneymTNZ8b4C0OOHZWU56
TAb2fmGcvsBu9jGMMnIoC51aHKy0brNK6DjIyXwXWOKz7pPjyazf22kvlHs2Mvov
CqJPMOuaxQCf6DHz0nGNSfzMuSIpHDoRW8BPPWCqwbkhXIsxbKD9Br56c2ebbkAi
81/7hc5wZo30MAk+h8USLia+TveoyBuVmSMTZBVYbpkwBAO0u0uqb64BXN9r3vli
nBmyfDmRe/kktz9XtB18F8KlVqqKuEMc+A/q4rIoalXiJdLfFhnop9W9UkmPbuUi
Se+0gA4xXbaSldhP0mM5WPlMFhlgAPhHaHer3fDRbbGt8NlNUMzsHzZCJSmcKb+I
6dgbkkkGbYNysoXW02BlUKEMML0VC6njb9jOEAqvT3LPr2k3Jmu8D3mqKrJSAaF/
lPhjVajtCuCoaQdGjBHKTgFXNxR6kZa73rTDSgC+bHQ3Ka0AHshyDAFFHOd27Ecy
LmQub1rlQ4BEhu03HAs2Y9eAIIsGqxciavHSPdotm8fPe3fqDgypIGlGzC4JwPyY
kw4bJmsUx7kAJLwp6B4di5qkjDhs4XlzpSoXA/ZEUy4E1BvHCdJJrIRcb7FAf0E4
hsnuKdTa8gSUGoJVU64zckAYifHcGYL/qqpKO3o0piNg8JtXD+6fv6JpLJMN9Zt4
ACy9aFqyrzgL3wiYqQclHwXVj43CBNIHopv5vIYcbd6Ix0S+pCFBmdvZhdYqZ5wZ
Icb5jvh6+DmRmTklMDATNY6JA7p/QTHT1bnyNa3vvBJnB9Op10kTHvkau/9QDsTE
QGwYM3W+7z776IdCUiwfiptt0YPPUci5UzP1+3wLXyrfsSe+YD9yMXIcJ4mryVDW
opLGrKzB31BvGEUwFtpsbLKsGjz88xHsHEfCO+rhSXWAvBC1Poj+1Oj1jpx5BW4X
1duyJBlv+8iPDCufs+hh26qTishJ1+E7paL/fbDbwZ8BZcNIVHKOe4eMczJBkh6g
/L8YblDW98IFvCfzdaKJNkzVpsm6Iy6ByXcED1BviLPSChruod06jGuCocczDiJ2
zE/On+NK5Cp8nZWC8dyzsT9XwNH/hmNVP1nSDko3AWYfBl4BcERk+wX0qcAS2TB8
t+2AI/yrU4OB2IkZvQQUnF3astaA3oKCFaTRh11jrE9uq3I19DE3WshK/OBCQINz
+Nw6YoauMHoRuuCl3osioALA6y13JRW5+BptOwBx+yTIVkV7MwnXGxCM424NPzZq
RnI+CC/2Q1YsK9cnAXdrb/MqsmKldBKaUbSe5CMpp5L56eM6gAhS8grYwoXml1Uz
YUTlhE1U9RvVr2PvbUEXbCIAs8gJtVu39TiXBdUHZA9CpmzBiEPVjVX59rO/t3Da
QrDTmHuIkV46gB7BkUSGrWLTn/TCerl0T6PNsgBQA9ec5PNjpVZqS9UURy0nApyN
QU+JkNAquTD1hxPNsMXG7F32sw1cuz5N+qHHpufr+UwpfT+9AlaA4+2TW3Q8juDO
F2O9b1I6WxocifTEAFM6z6MofcfE7U5Yd7fMI24qUo8IDcdH92TTuAobR3GkKLio
FHfqEaKyRgd1n5jGcfSByFRP5PhSEQluKkHnazsekGoL9uZD1mNcleYuis1tAt2B
Ye4h+zvyLuydolXuNB1056e1I3pe+j5W810/a7o5EYBh3gboRUPx5e3cpD2Ettdw
GRW0+u7d8maisl2MrpuYyGZSGL3iRtzEsdm1+YjYnk3Q/W2WZKsITHwSOczIm795
HDz3nvVS3UgCuI41sHW0U2yn62pZCno68+aoIecHblBgZWuYX1dARPKv8OnW/i4N
vIo7ujluN9HNQDruxAq7qk5oLM9A+Vs5F/BSG4Nq9rNapGG0LNUes9umKIlC8+Di
97JTWmW93oN1W5XI3r6Vksv3dgvkm06UtV1g0wn53pV5Q2WLlAIFOjt8Lfz62zUS
veSfTEGfxuQnCcXwtkjbjV+03m8S+2NBT6U4Cnzzd1odY+jEKFV94ODcS7nnaLJB
nCTOXYM7K49vVrDxCpZVtqmdJ+tbKITUB81SRrNWT/AW0hCM1wvMT0mZtmzr6LjZ
yA91wtBkeGgcFapsUFW1QPkpR38Esh+fXLWHNglAe6PBC2inAHYUJk7TXMzYCn4L
pRWiZBs550/r8/yzyftN2lbIq5n/SdqvkkPvtN8LFArbdb5BEgi90b3ofHVna0D0
tVJUCYduEDwbn2NOl1h82GxlRGJbJ22sT+L47pvGb0cQQkhfkchp4CfkAUij/uq3
zA7rxIznlxWRyixYwpleTvi6f9JzskJXuYBFH6MX9rWHJKaUJYYMHlpgNWSeTA/O
cVLRGJzM6ATjayXAi2y50mnFe4fDtani+YSab6Cu2C80xAfj/4XiXXCS2NPrPOS8
0eNqMksB30mvR3R9QhkvT1PHXsGGrfhyfVHzKTYn71kbWwo5K7Izw1TmZSTKNpuC
z6ACuPyUd8GKUvgg4RxV1T82qvY1DP5vkOZXc8G/C4lb9cnI/GqVq9YGRIq6vnOV
WeyBJZWQTITQND4jeM+v6hJF8MuVeZdDqdKqPl8KQqkdD0R5wRx5oXK7pAmXdmGE
Wb1UsS1VgLV/COw3w7jBiBFIoZpjWR4acwGiQr4cUayP2JMBsO5RA+nvZcHkvXqC
0l0X5pXwHSQK6NpzdOljoMYqzQqfUzOH2TH8s4iWwdc4/r09RdarPJqsoUeYsN2l
WX8JzY0cdZFRd0b2swGw3c9a1LOavNBhAaUmSsd2awaNZ+3ACPicshV125b4D3fG
1w2PwDPxFHDAbORz8JfjKYTX4XpNqlLEdBa79c6iCoinmOyT/IeuM7RWVbO1zqvq
MI7bSmAFIDpbidjaqlYjpWF1zDO7doDK3fE1MlVVPuvf3E9Z8uaHrfmndVowqcO2
DPI8LpjHO+0RgNqsuH66ztUvbKR4az10mKqCXSy6pkFhc5rSA11Yuw2nOYqvrTKV
BcDNHUWc220chG6UdgCUKKlFt3Yqs+6kgjIXYw/dMla6RrTb76VNA8wu6NIGRO6B
P5mre5ni+JC6M8jQwgnFa7B1naps37LKKsCsADoTSPuHWwvVnbn1n5Rj1xUdCgLx
siwSH41ccTD/VvubXhTUwQIAdKPk+qMRR8WsBA+0x/WCm/t4Gfzd1u+EZT06uKf1
TLKhJufcyvXBQYVZ3DKeMsAjIPS5BLdauEgb0vJKCTK+8ODT33kdf+C9l394Fr5w
B70xJwJmHTrR0SR9OjGp/GoWZ+Mbwg5FNQTv0sPfR+VH3FXWmtjSyA6yOb8GOmq9
IsalSF7XxjMEAgHQQlpfGEAD4PyQCkTc/HQd0YdzSnz8exoSoVYiQ1YSIdeWMDRd
MF9yIxT30JoiOgFqzhWUF1OaodW1CAwCJ7wHrbhR9Fe2XsFtNcac4yd7VZuISeE6
8lUF1waFQjZKklx3FKfji0cRKmUb+7sGZWwOELP9qGoyGqgjJ5eilo8j3TNzv7Pl
d7nVY+ftDdgTvhAGGqz++G1Y5jGRhOrcmZQ8dSaBLqID1fP73qc+H6waafKQlL3W
VuDDMwnBkNcw9U1+vaqnING4X74Q/bP6fiyjNzxAvo+vrWQS0d1gAFyTl7OLqjRK
w4jG+DmTBYcZMQlDVQ7RFG8hkbh3LrSer8uuROnbBglYJy4TlCpwl6k8ORKydx0V
QSSHcCx4sfT5ThqZzIizYJQDzSFIB4H8zaYZZPagtR0stEmR2R2qQ3ZCtylppuD2
KldInegdGwS8TdxuZPWzAwHkNLrnI/Xhj0wqRk9P8/LVpZAC7TwKQov3MqkZZO+r
dG4gX4wkq2sthtv7w9YfYm0ALMd0U7bT/F+c00CiVRO1Bfk4KDXe0GSgu5o4Id3x
xOyoOjWtyLGhT307ilSJuJ0+RbdtRO5gLU/QbgKCcIO1dJjWziHm0PoDAtKOmY/U
ev/sk8ix1nySwCAZLTLoxoI8Z0CIcITq+wQJFfewyxVvpGioo8QMTtoKgfMVqFR6
wDR1MYTRZUF3FcDQ+bXPw8P6aNVIQbVkLIRkuZ23++KvxUbeQtyS502tOUA49IBf
iPl9Nkvqqmy+7RFn8EIPvDYYRaJ2VHqLm6AxRVsjwr1D+bXW0pnbld+xITSc+n41
W29UtJnb15myCbLpDGrvPHdHcroyMncMNuQQNq5Yv8OirG4YnSskjuVaxm1TZEGQ
NE6kIQ7wHsA2mFd+5EZZ5fv4kCDfORE1lOkLY2BVDsVHdmhQpuMj5wTDlWq/RFs2
bAeSIbHx67m68Sl6cqw6dyCEfcNSTA0vxuZ6AB/EX4E9nYWoX0dQPx74I4YtbpOJ
DCW3xf3Q6ObSjks6E3sGIIfg/eCV8DV2n68NtCfRezocjZQa+klJCZ+jUq9qgfCz
SgVG+wbX2kJEGluqw82OgjmI+/L26M3L0CLpT1xmRlB2RfzSeDiCut5M1IVDUPr1
GNd1v1L1CFZdXpB9bvlp5AmSb0rSQKNikL/oBtE0j3w/JE6vHQUEve5MD2DnrIBu
2kJ5kp7xG9Hg4vTKlLArnj7q9sSlNseUZrvmOspzwnxYXdvco9jRKX9865LFPez7
V8UKfhqi16Xe3hr1j/aOngDduegBkV3LZNLHA8bH08b2cprWLQhluI6+i26l/PR5
GaezjTTTDwl7AwTtuowcoDa46ECi50JJ9J4GlObQZ4SUKuIza4TE/6WpmGTuxkq6
jw7LK3pW8tE+pRwDsCrT6JcjnApsk6VQLj+yf9h8LYfp687AEb5Ev0pTETQ4bqNY
MrNPwviYyKgcfK00v52vX29c0e266b52cBvn/GpB/AglHJCuOUD8P8hGh9r5q3/a
ZhlzE+lFfMnu0faEXZ4BXue3p9y8ft7zKn7dD+1jwasm8bPfjru2a8n3WnA4lxok
FkuW+uWRvMmTsl1dINEWonUFO5UGiuRrUUwxr5hoMyFQzteem/1j+/OsUujvgwnb
DJD8+mbKOIcs2dKIITlBZP8m/Om8D+UbNarjqhp3vzzV2ofmAm8W5wRZ8+aIjNZj
myWeyKE8ohUXVTNH/0t00hmGXv8AFFGKQHSJwccMPGHOFwt/Df6lmwjHqt1BQnJM
qh+dQlkcOq/Ki1SY5LNUTVQk90mMmeopkVSls+WKCNa4cJAq3s5uzab8qpvOCkGl
bEQQ+IfVjGQH9qM48VmmOQy0iSJyhJxOQs/zkxt3yYr60+8z9XpWkttHQxI3kzvf
c9W0AlRxzVVjCWTGWBw+ZJod0FhfjUNfKrozDr1oss+n9YALongCfxtc/5I4tdwz
1ZGK37TOQmcVr07W2F1HblDDujBSAb+7PLYtOfzMtLdbhdiCo+C/zATRLcZJinxo
sTxAzYQrg1cFdkh0os883AZhuSpsTv2wXsrZmo+hEUiGgZZccQL9ohUaRhzdCiTj
6SzC/BA8L0BTgIBeZlO95rpWkNFUj5hW77EeF2e/9V1OzKLGVx7kA6dWCamHedrN
vdQskLQmlbBvvG65YI7+tVWtyhzbBXiS311xJf+j4gWXR9QSK1s9Oxv28uyx55gn
TSHYS9yoTAyAnyoNy+Mge7OtgiUL1KGdh+z9J6WvTd8ithT+N1c+LxQ7540JLxDJ
P+4BmrVxBC7vS2GFxV9Jt2xH1YSOS8v6fG0q/akblnvc7/6nqIdsUCX1dMsGRPVX
nb+7QgYwFmOaumKFa7IfF7LkxYmHLIhMQ75JxsBM5LBkVaCUvJmpWQs4qI4wy9uK
xtnBQJNNJLvYAcTQ1TqhHI5GHr2aSrWGZfgYex/yvszT6o9Q3bGX2+zpEcIBLPpl
rX2JlenMgWigeCHjkcdsQv1V3lDYY8Yalke6S8mubIHbPR87gIgiPQgghIWvKINJ
MsEpf8Gz4HBPPGdOQJgGRemMecNK9hdv3dz5PijYPIHSUDT+j9Cx631tpNqNbXRV
ZMVEIN26BEb95krJXACoP2H4LHxYDpQVOa/txImWXeE1hJ+f/EtdctuH2KVz4Qr5
xfVIFykwYD/LaaD5qzSC9NEjejVFp1HH+r4QxbQ2pjRnZSFOTzE7mvxzvHCmEhFX
bNhPJw3k0c1mMyURHsmjwjDnpF3B38KUW0xKgv0CDTMowOGluJ9DdQWqR0rjQc6i
t6ObudchIMwU20vDSP3VHi+8mnsS/1FepXCm8pZVeACWGYhnDk5mPZlG8953Aeq3
E5ca3mDMOi4Zw57j4delS60OcuSrsCHfGUnWP9O2wdE73ledx9FCjYD6kvOGZlwX
iLXh674vU64Vc7UOLVDQgFL/vC8bh5rWYOCtf1UJvcLsYrflc2dTkydBUhO6TSnd
av1Un2mkbyiHOIKTzt/wDQI9maXST3R62E2KGPu6IcLu9yfde9Qv6vIkIwi0FqJ0
/BXTLEC3P233pvj4IllhgKaL5KGGZUK08KeADv1DncqNgGmChxjiIT6Fw++8hA4/
/yrH0vd3QNb5R6oxvwB7rFec3FaMO1yhImqUWmQUWksanfy78/i8i5bv95t8tudi
mSDTsDf6Vya+699CCUYYF7SQ4jXc0EctV6Otozfr7pLa4dGhqujowsL48YZ/A4H/
yqDOUv/TKjYk20RMFG0xnnjt76uJdm8ysqV0WXfU64iR4saJz5XWRQuuBnMHizdX
DVg7gKzTIUOoeCSSPYrD4vMZT+9IRFRax2kh3I2FzVXRWSGJjT8lJ3siPxnJi16m
5ZtFz6x0oVl6skRITG0jHousv2onq2d35Cv1fP6wRV3+4CR+PHaDGUs9ucIQyjOq
6ATD7nHjm3M9Ui4jfFAAvykI2oFxjjoUVPLKv8j69iFQTiJS3OdjJaPIG3K5YHRv
YB8hs6fRoz+uxrwWBxwUkbfp5dZF92+E18d7rDaFumxROmW6Toiat+OLHfpoRMP2
AP+G06F1qBVBF1XIlsUUsJwaHZTVThVK8AnL77vngbnnSn+f0prJESf/O0Rbh008
ksT8ah0uo4ZDsZKqcVnIe1ydOXz5v6f2y1tKr63RwEgyNdzNvP+kIyvaZF7psx38
kcfPCNbfT5N3BQPvckq9BsZoRlYZcul8O94wdEalz7yRrphTvOijRsY1Q7aua4ET
iWgLcjg+t7eTRaimFePib+u5jLVelXU90g3hfJ/w3IFfrpZL9sBrP11rObHHewS3
G6olcDd7VP18E8KuMJkZfHOxSzAIzkg8pTjZXVyc+TTQdyJFJ5la/WFjQOrGVtMk
jneoLjZFFpqYl83sf5rPkZ2vy5duepjPZDBq0BIVgzC23Z+SPERrW7IROdbB9ERo
PJIbfuOQGUB9N1GJutmPPDDp+yivhOVfiNmKGxWhlg9C/Nw5dkHtM05AmWNL8XKB
RNW4U8D8I3wsrEADU1sU3LjgwB/1TMLKt3GeEI3riFZs3L65DD1GnLL0G9fh4Pko
FkG2f79sMQVg5YeS6rlV7sDPewNEgGFWZUTm476kQYhTs+L5H/ydE9qetfprtk04
UXwiVcq4IphcXZ2GIQ90t9FCtGv5YRgIEfx7s3YG/UfNptEEAKaC+Ai+/7k+zy0B
/CkdJjQJAxXrc/y4RFRh8vmcZZ4foxFwzblReCrkOBg7vMe6MIb5w5D4Dfs0Y2em
wV8+fzGWJkjnL5btE4XyxOuFvElnlozpiC+gnpvgP2gsqNlIW0GJJ695AoWR2iu+
aPWHrwzs6nlrOQu27kSrqhI3laqyu0oWFwmEmodS4AvheBEyxydI3//LWmJ1EGef
LcxB1fgwp9oIqqk7TFV5d5BuTT6gZZnsJAV6/ROIGzmMyWO4Y+5kH5jO327oIrj5
HATetHtkQ+8c4K/b4t1xjfaVy4j+JzEnsut0A/vT7Lv9eHtuTF3w9qYCQiRW2vJ4
ULAdGbBpYy5/mQDF4iAllOXmLwjg5xrFAnm21hlVHS6W5qBqw3/UXK0S4edUdLs2
Z38z9xL901ouPtb+CSXYVQ3ebYA+WeqEdgE+MAZkT+IMY8kdMmEQs50WyHTZsEgW
0+kCqQVnic660mHQ0TjKuNBxc8BMI/siK/4ociQBi2ElB4lUN93gCtlI+ZZqnGMm
Xl6nnE0kC2garv7uiqZQNUIc4j8Cw2SN+bzymKWB55UwRfaQY6QATzrYOYINm0Q1
UuSOC22mBSfPXltxCcNm0m9D5QfX5qAcp065DeJJfGJxvAPlR+AJlS5xT0QQcQfy
XFZc5obYweRvNqqoELBug61Z5CrdNwuusblooPZe0dhxkgTmkEqTlNt2tATHjQKH
rbX7b8rn5zOkOthzPNrg8+OQENS413qdM8KMxkjIGiiwShU7xgWnRijBcsdwsKYR
3KKJLIxaofs2Y/JZr5c/NoDqSNs/SYLjnYsvkg+D7gr2v+GqkTAB83XNX2nyQgGf
Y1YAHobNOocXYg029PaWexNovUEqparjBscWxmYHIMQ8vFJUnemOnSEERpy9ID+g
wJWPKhN2ZZCxfsZDSb53tEcfbP3a4Msx82t0jIlTMwXANMp8cjBj61tIDICBjYTh
qPWeRYuDcHM5QxL2gIoqA30Ry+zVe0AzcBpkfFzeazCNVCMoFXbgyh3an1S7feuL
k2jrLBE0XXaCwgIeKZauCM6hI/lCBqhr7VSEltUkFgWfr1PNHv0e7FTWJKIJSblC
w3J/4qO2tyPW4GSaxbwbFb1dBUGZ/YKQimRpOl1w98uMONECmsPn9/ZB4rizlhCI
GUiIZnoMCg21OU7U+mKcLsDQQXI/LhmeKGBma6Rn2/wXS/8qkXiAKSqF5XyCMj6z
ciLOteZjqYj4KJjGPu0FBSD8dOXrDQNu6WdImqNNWLYihhJ9btA7O/KDMNEtTDFN
rFw4AsZZiew5SO7EocODsaSFHp57BBO93DuncbxUTE5z9u5IfdEkHeQb7JlKay8U
F4Ic4c945Vj1ve2fsbsXZ2tnXvxDob7p8AmYgFz/2KylFnDnw82IPERtGLcNyP/R
THYFMJBZVAMD5EqJqA3Nt8E3wbOSCw9GobMECc+JMna3uJKxgS/MHCnHcF2t24gN
Aqz0GqAnPZmyfqhikq6/ugC4gj1OWJOxbZVA+6jr6rYXHeF0H0eFpxeWVwTBB8jO
Iq1XZZVLu7wqtSSiMXV5paSyC2NsFW3sMrCHXEjjdXwI2i4ydb034LgGSCuVFizd
fNWOQ6hz3UfBr0rABcHCNSXo99XEfZCNtzCnzBKi7ciGeYDEA8dNZ99wyn1gMngc
p2sW0sxrxSBQ7znsJVb+4GqE/2NbOyJQ9OhnXPKAhgYV4/NjhuUET8vgMpglg5XI
QTMRQJGQOrXOz/r8/a1c2hWTS3VDO7cvf53B9HxeV0nXBIvAeIsw2hdKpBkhg7AY
+eZ7DuCVOylG2M/bRQZtarzGLQY/bdtfGtB2NHzzbdiGfIVFP5Q64mJnjrKYvVBg
V2nf+Df0dWJuTAiy0iOdDNQ/T4hXcvAzJaNzMcOGqfNQR4ralDKBoCIf19F2644M
EdD78PaH/WxowKktwNydGrUtmUvYpKB9s9+tI4v2KhUwPsMDaZJWsROmnlLUd5Cn
coppuS59EdaijzQ35m+/7qjpPwPTfTf5Y6LNimmJJdGINjIlBKJooLQ7zc2l15W8
fO4oFUbFhZnpqnQ2tAla/RWfeqQZ8m6BHO/QWYI+GSq6fWVm2XAZfohUq9xUpo58
/I96vWy++PBVkm/ezBeJY6lnlgWZ8SeRV7CjuF/8HEEOuCpkjA8I5D86L1bxQ1RU
fQjpJ/mAH0UFAaVW7b0Cf22CfTLlaLs5oYFDdqSnuAvTmOBAoiIDpM/ZCCyQmCRx
biTalvAod9uuGKtQ+JsZs+NKV6qhSzOku3GgdcV2AUWGPcncmrPtniLkTHjfI8ET
lVb4WDe8YW4su7fnJme2R684mRh9unsRrNhss+8cOeD9Tvh42U9PeDLAsHbw4vTM
viaqG5c01nS5Nhp60RBEyMO+2/wPrGZfCnzPl/B09hFNlyjKwN3PmioyyFTPvBNi
HNfbXtYGmqCNgwJx5gL5LyS+TDhrEXuaCwSsdmk1/YG2r8lKeGL7c0vQdbCNtaxQ
M3cK5rxlbJvz+QzI9nlPI7LWWmJ7CCt572tZVKx7g7A889uRs4r5KmKOFSsp9VmP
6OzAlsDyILTJdoFvsoPS+T/TC3+XsNyuL2jlG9GpIDO8VWLo3zkB89yP2gxlLrdY
Nk26pt93iZ5aN2PFkWBF7UYgPYRcBwaBSys/vgk7dwYDinzKaYQsUuyC5U5AfvW1
7mJbWZoE1ndZkLaIJo1yWB4BsKrq8+57vKzeGF2fpK7yyHk9E2Bwyfxd6e2fHDvf
/Q+yEK2TNW1qB8p0u3eZC/2p9RSl6dijC7HSWdN+RCWEB3n4DJYA2varW6wJt7Mz
GMlnK851kceaSqguF3Lz0qMN9AhtqRE1V/27sZOCcdq61E1oT0ylCDGa+hDDf4II
O7BOuZxGws+Fb09PMezQWdSqwszKqdaJ+Kdx/RpbIEdAK13xK0BycI3tIgec+2o5
lgQCAtFR4Ky11hg/ryQbO5X/0SSyXVnvmTavN5f2xdjT00Ki6NV1kzaUZntn+uh0
D3JYKUf69aeujDCR/0QBrtsCXa9rAL1FIfDBSxXaGpPeLUP2+WyYWpmbrR5xGydm
BJ1aefl7UoG/4/QaCf8Oc66qXv0jyjJcfAY1SULEqrZq7Qq5G1D/WJUgCEimEmq0
Vo72mVTgDD97scdwIWCTYPLUSHyAsxQvebFTy4HB5m2TFZ5hdgKbhZ62IYzXeX7g
9ohlbTou1Qzte51y0iInoZOL8BGpTCdDE6c1z2BPPngfx3jVy8QicS+Ay0y31cvY
QRSnk/DeU9hA9UcxxOt75MOVwU7gA5jkkzIJePkPfnAdnjljRPLUjJVo5WcPXv9Y
M+uxN+/7VrFiSazNqtHFPaUOAxyT3MJSbAM4/yO9S/kK4sRRYPllp99v7N4s78/U
lq44u+ylG2lJkcG1/IVGd2QInhhuAP2DLhRToe8slUl8cgMVD5pkSj1UhaUxUteY
yC64QsO5z4CglaU1wo3h3uMcKv1WWUj+I+Ckal+QQekd5lJNdLzLg5nedagxJadW
l1iX2SfgPctxSfHrF51gDYVCoNiutjamHGJhdauWFRR7lUI7FXNgRCB3u9wGDwqr
1b5BwBlnaY/S7F2q22YqFS9/CmnH4hSDmuR391CW8MWWsiPTZ9I8h3lI+pFkyIOA
LG4+BQV9hY8ECAPuMPHGy7aljaXbA4muk3//FPRmdn3UheMh+O1rxdGW3nvetm4p
VI1+zHIr6s1zs1zHLwt5yhfNJ+6EdvKHAwRZ1mAySrfJyAQHmpEf93SrP2CmcPwD
w3nyNcjEb1kNWBxFRcK0GaBuhhrfelekfj9/hCJraNl6PatQA/VGgJEJTVrZQ1o0
MbT41egJte+2JC/C241vQR89ngqLndM/bx1H6B1p5WuAahB3ydmIphFwG6qY0XNx
X8WqES+x7EBnsJMZ+XEv3LijI/xOdDJpyMpmuVT+1FfC30QKf7wWetS3Bf3XIc0G
/C4iHzvlvtXfm3UKkbGEPxMZkUw7Gpy9x0Zrn9HhhOaQCWWKMfTzPcKgJ8bKyBJ5
kn4j3R4Y/raELIOsWk+e0DvKUUUG9zYyjyRdzXLlDddKXpkrtFOzFQ7Lwa9h67jD
wVMTxwiKQSwiUc7WQQ7a1LTfdDLZT4iKfdJ9hWGlZ7mEoiKby11/szU+kxrL2o97
8hR1PZg0jkOdz34+cGByg7cDQaOZZcj/IyGuqKSeLPNArXLGA52LCFlRLdU/Oubv
wUN7fGIgDbjArc3nE+cZRgHj5Hnfk8zxQ0afjb3IH9Zlbyk2QW1W35JVv1oAqWzn
tu8M4IySPkF+Wh2vAyqrynqriIXXpwpfwBcRMRvK1MhpF26BKl0Hj2YmpvfK2dLW
PYQ4R1j3NWVWMPAuxdDOAHH+ktYeWqboxlHRWShujDliHy7yPI0Cy4ZAXzmiRfID
0reHIeyVahPgiE23tO50iBAAEmttGVZAEKIqUpHHdoiCBBm3aWaWKEJdl9zaXakd
Igwc+wF2D46/35SUKW4NJPK9S5/6b5K7OHwvnzLTU7LONWUAzZXjXAkISWuxs9ZS
8CH1LCr3RrSPKY2sbcRKxEf1lloFykBpJXNRus5cytgzQVOmbI61kzCUXAqhqlpJ
uIguNX0+NAgLF+TyKHzNOoM40Y8AZpv0X4e4vdKQXgTIK7pk/LJ44Jx9Olz+tKGV
P9KXOPbJ6O2w7itMDlfNGBcNw27LlN9GC++jY7SPQqqt50RslFD2MQgf+vDlpAsl
ThSeC/kBbUIJcT1u0Tg0fx7X4hxL95XgvINMv7oolCKtW16SEWkPeJMk7lHon5M2
qq04islgbaiGEFROz1Tci8zvfW3Clzm0p2uK6wUp8JtunJCUeKMmsqRkrxZ/62WG
9aaJoNPL1kf/8eIXToSxrHSGaEEyRXJXUdy3LvQieJvZ177Kn4Xa+CLOI9xpYrOk
MXOt8dSmNcQy17VKDD9BeCHxKH5jE0rOdg2H33LaFHv/vZtf6bRbu4H1jBGuW50m
1dZkxxlYgHJqHlZSNtISuop4iL21dplh5Z11cll+AvF9NcnMMgDxnDqQG77r/llp
MVJndqI4vOP79tBywB5X2OPJ64XKmkpfYpwFwIj5DE7TYjKWqJV3zo8rfZSyvOM2
MaZcPlnTY3FjgaPwafBb+Dwrel8/GOaM6TWdAaQDSm50GQwIrBuB5FdQ6crxapBT
+LW3l7mJHpmBcW8WrEeZ2lgiDZdHKdg7JL8JwM8DFEMk0bAB4RZhVxF2wgYszg+r
n4XT2eI98v1HnDrnPtpsaRzCO5tKptQFnEMiUO4JWEmCVyqvLkulyGxkFH/WlrWS
EtD3a6sOtBY62O0HwBlEXxCWEssEs+O+1wx4Ee+5oZ5JeHBs10julbfKYk3IrIEQ
Xm6WxG7dzXseh5KfyuO0KWnoxA3SyJ0A90md1NrO6z4QvhE0LDqrkSLKMTlJ8V67
sOBXOQlXVrjk+qVRD387eZjzLtRZDNSVx35hM7avTXhOTidI4sQ48Y4mj5Z278Tz
IBAFCp7FeGKSHHce1uZfJO1G4OcZ66amf85PTPygwOCcHELGJ2Zow8O5Hp8Vr+5r
9e6cGZTROOeDvbTkTENxV7aBuJJ6TwcSf/hpTyN/TjwkHkOrfULZ/yFXG1kn0UYW
aUq01KGdAngOKSo8TAvDEmzBzGRq9CpK++HUJL1Pr7tEvhV1bcGhW08pl4rP07SZ
m1ix8wYVhk0WbCksUoYMqZpNt4sM+MjUe2Jadmm4owO9KUVYxtGtQdco5rvpXWY4
w3Vx8TYgWzYC31BpisizJScp0sWH4HMB0Hxhi5OYzoAZbvydM8rpN8fiXyYL/wbP
730uwEY/KslM3HJkInbiUVHT+o3nN7qNb5hOw8/SuD69k5DNMl3JSZrlNtsanh9M
5ytr6eO3mXhcymoQnOZgk2tFQYxzM2pVMrM0S9XvYLYnb/roH+LAMwbSu7ocgRdq
4kAi0CN9vYoZGwtwuNRTkREuMX1zyZIhL1y778ioYYaOh5ss0WG1Qpktb6Jotnho
RfIxPjWqYzch/tK01tlNi19YxJ2kL2f2iPjBELN+/vG0WBpXHVwfAp0rSWyVkNik
Xn/KYTqraLP09IqxGhIDoa4lOP6OUdG+REhTjrjFQMxuRnKJ1LY9XoRLMQgNAd08
hw0+sIbrTFkiD+B5nQsLgJ+wswqBUF+fZyvGls9jvK6uPxSdnWiNn+myT2vz48hK
nZavV74iG09sBl5iYfl3CP4yGU7xgfVS5JLTPYEP4976Ue7P+KrW52NrFOwYcUzS
Hiiyi5l2OPnhpuf5xLRCdef9i3DD8How84StwdDNcLA7f1vmsDkQ5oqqo3YFeYgZ
CbpDR9Aojfr8ZWO2rnxeCWVbDXZYyUKl1zRwNJlG+u4b/b1af/oxCuESd2Qas3Dq
k+co9UYVplUdje4ffW5bNNNZcUBjYN6YwbvC0ssg07rwVwh9yuMVlEx8uazTi1mO
aiz1OLcEOCMfi6LokTMfSjiooAZ+aYjYuWLYiF9PhRA/2IlbgS3W2DL/6I+XhFNj
Z4NL93Av+cGwewUK5V6odJ8YQoR6DRocy6tRK5Y9aZCc8J6QZ+KL9xAlII6DFvfU
R3y1SCGpu2wSVet6QZxc+MbjZ4Mc5pwipOKJVSXeUyp4SmfEJXTD0T+0NWTR4Kjf
w2wo+3bS75SieJFgE5cMgjAvzpOQma7OrgpjaiNKfsxQmf+zJ3e3psFu53OcY+e/
T1gb0TLj63ge7JEA5PMw/lLDnrYU/AOo62lpqTD313rdEzm+T7tSD7PntgFJ9mMR
eCsdviH8Y6HNGIh33nF5zVPjUNbId8QTAK3b+RVtSU9p2haFuym0mFGz2p1GktrW
4q6t3lQjIIed5z3lpYCbhjnl+gszy9mqJvkk4bfGecoVp6xDIXqVHViUK0lbdslh
/YK+uPodT0T7MjLzY/dQ9utl8xJQ32jtRciwnx1AJI9x9v0yTEVfvMaTvue7BGH3
xsE/C+MFEql6Gfnq8RSrXntIHrJenP/K3wi98RH4sQMVme0V4dtugJvT3ys0juG+
7yIrIVUpbh0lgrOzo7yUXkzO+p99wQUfo7/v1mJj1zUsk9sAiW3qQkuTFVvNIxA0
gMrHUDwn+1ouXqT5/duTGotjJQss2NBTiwwHIiPxI6W3u6ZA9PLWR9fZTEzYvJGH
0WxIs9NivSxWHVGJt0Z6D/lWxI4PDr4vocqwVWE690xPpLWYn9cSF82mJVlo84FV
xWd53nlmanEaUgyupG373Ht+9POv/k3AbIKwcCdlla6MsFAZNP2BcvYZ7iq1z09X
FFSs9G2d2ZA3qL0mZbzzVZWZbwp4PUUk1jJsyBsEIILnYme+SdAjErwDXCvgNUeb
t5RQBLOQE85EzFTvnZjOwAjrQl7ym1/BQd0Pi2funQiwLcVsnqbBq0bNGmtewdcy
Fd3CLzc0JhciazHCGehoqlNLuwt5Qz0sddcl8+rsUvorU8k7py/4QA+at3EwFXit
tQVaVbTTMtr+gSZyDawAOFcG9f6mBIyYwpEXsq654vL4xmF6LAPWOZkO/Z58QhMd
bl7bctqYNdYrv/rVtrY14UQGNrZHkVPOZ632oG3PMEehGDnLRv9XIzFpE2gVBl/v
reg08vT86axvWpCizji27vL9T2mYt4KW4JHyZ3qQPgPAi/Y+lfMQTtmxcEKU67aJ
kq+aHFE6rSvctykQMHvXMn6EiiS5TJgh2S++Yer2FoagTnPsFUs1vJCVd6OGH0x9
PpFPpawTqgVNa8wjlAEdaTfiEI3jhWNuC2tMfNVvCF9GRoyRJ+ogQBVF8WVAoNuq
/fZSepCKjfznYlHlUIH2bsE9lu7eIyAEGM3d92q5Se8rPxIHlWKhZhLDvku9pag8
SBn/VDu0mPvDJAX3QrcKGrH7GY4PRlea+Z2Y9zKlFwWJnlM/x/s/tT2BdbFi8SBV
gkoLlAkgDZN5tjJ9QwgoYMo+GpVt4GSDeFGqH35UyQ9dfW3t7WyrQloRwEws/ZgI
A5QleRS2Me1Nq1UqpfCxNqKOSkdF6f1urSETjTfC3MRtye0Akvu+LImixIG/zl4z
64bqRcRLqMWosfLG7VM1gclvipEYnmioNHoIvJ6C5FObZJ3e9zKI0QkS6t9tUoV4
bs8Z1G1qFx2zINJZuSdPhOP+4BlErPo5SkYl/XxSuLAwgwUxO0Owu3JT1iNm+FlD
vkLnZU9uXRmznMu5aGGZMaRj9m1D6+I5mQYgQPJCz2CVl/KlFZhUMQyh2n3kSaVX
25QGw0/h7KeRg7jyBiKUAmKPFMRPyG3FRS4deB2TIkOnttUMxwoTEtLgvtTQOUTG
GC9yeQp4fmU1MF3gD4Fa+T4qLo0ZxiYnRxLHPRckbuBCsHtJMjqCo3DSEcVchCqK
I0S6JdcaLr0J4aFzu+MwPW2XOsDrNH+8duaJ+cChaXL4TM5IdcyNil5iDTa/BZiq
jCrPA+rmzmEbijAModMUU86qaK/Vhop7K5kjK0r2aWNhCE1DG2jD6OxjL30eFvwI
nkraMfuoEwWOj7Or1aECRbI7VU/PJSPdsjZp88DDoIEnxhjvh0Xfdl4ZE8kpYEbg
Vq0FwVzB6XghQYteH61S2/+iz9UrZhnSWvKg49XJ7aB01AABl3sC611QsKUVUklX
SotKwH/mQs3ioNbTfa5/ap47Uv4U0zOKHXrUCTNkO45Q31HuSWSD2XF/GUCK8Maa
Jn0h+9Q2GCX1RdKu+HCu/G7+5FT0Sm6cj+/EBg4JdRwA77ybMqNYABd2PEYYw1dL
4nbY8bqBa8XeprJ3HHpVZhtPZuXpNFMCoybniv7aItA9j1Pelkn/pCRalkGM6cTS
Uwd7YgcBmfhSV56CxTPfYBm991nIFUzXX2er8UmpWq2eqIcb0Qp6JLnWwbMs1Ho4
FA4bd+/3Z2AN/w5tw2NY8+pQQoa5z5pT59iWSHMtJjaBc8OfRkxhH3iz2FA5Pnj+
GfG/IDnF4CDNXtMcjD+VECNfWVdc6lykdE/X0ytiCLAVw2nKx2OqDCKNUmfUoamj
GF5Tojp+YKmymKsS1jyVDMUhTdedV1vo+8mSZk/7mxzYXiw61uX7xSxTnzO1ttJ5
g5RIK+hAtC7wPo7ygXzRp3xItnoa2eqSDNHKpNMC9+0ZKmV3jWmlqkCfkn6FYvfz
B4PgcaMMgpEnUatWZlyaNO1zVRDeSeegiVFIgOkiaOoYtAjwJtxi6jPc/Uz3h3rE
DA264hh1Z+80UGOUjTMY+5MlzEj/cZ1vjMzrXab9fWJ36T7DZPLlh5PChUaVRFC7
Dl1BrcGpl8j3T+kve3H1TtbVlBGvpsZt9o0MY1VpQ1Er11uTvCWg0GPFL/9tWL7Q
/AvX9WQ7pETvjBdQ/NlNWRxnV/55HzzKCQKDJRos/upNq47SBx2p1rjD4dF0tksF
N9CdQrrNhvzbvKz75Id3El+JnUQLy5WSNhxuCBftXnaBp+hS9Dj4zulYFQRx093q
MK2YU87zflPbhfXoaTRV1663eObxDXG8IfHhQGBMIq2c8g4z48sj/IxfFZ8TH04f
NL57aWljOWL8N+AWSoapQ+2PuCsemjoWr3BHsXtNpUEaUzPSDB2Rr2bciIZIZfVX
LJVwHK6BxBdnl2sAPYQha+VStDyKgyXR52pdqqEYL4tcF4W1QxaHrQ4fbQFOhj79
2ywrzAYtK0XtrHStv+lsEeUY4Zdom5jAT0+1ANRsC/e7Blba9lCyr4bpdUdvuUk/
MpTLnE8MuMFGZj2Wwy7K48pYh0emcd7YzHNG8Y104pC5YlaTNcIHyUJbGrdkkX3c
T/vePHPnqZI+XumU+dgXfeoc7nPnTN37DVvvTWdVaXWqV9G6FSQxuyO+pL9Dhf06
m+8jLAaAyQjP5x8vmA07PbboCyaPJDPK2wv/kcUCqkL4jMYNAXALaBIChbOlLFiZ
pvBVza8Q1V4i8ZWH8Az7YbIb5NG2WVIDD+aeCmLl6/t//BUyNS5VB0FXEqEKimhb
Jv4tHoKz98ro5ZHTSpfjAL9Cxl0KA3Q5kUYhbMMe3WCjDbFOMlA4Ni9gSjPz9P63
8siRZ7iY7sAGq9L898/Ipnj1ZH2/jqkolOWJD8c7/hd9wD/19QqI/n6A4iYzgeLN
V6NBCJz7SbTSMroyC1RxWYBQxmYEHiI5D7kYqG3HG+oZUeRunYu6auN14Uxvnog6
R1/edeKPeRJerOlK9D2MxeBaNPJkAhd38ZMZ72Chn8ymBbn4cMoeIr8v4Z/wCXaz
qbLuk8bG63jK8wXdJYEMaGVB9oGkp3GzUwRGdnJ+JPwJz3WbUmv8AaIoJ8C0jq9Y
L90kIZ3GDcADb67cYJitPFEVSkwQhydIinSwUH1ldAJpmIhmiyfoPLSBlAEQB7JE
xkkbODDiDvwvDaOVdfC3HSxFnApoRbIlvuOOsyE/vrjTfYDhjBus9A0D4oS+Z1LB
pDLutWQCBHIwq7oYl7JPrVwMkOZMCUcX96cDBp5L0yY3o43CSvxzS/8nJ6Zb6IQ3
/zaNAxUfx9xtmr4JnpZGA2RXQYAK92fW/tYT3C1CqQf5x+wwJMBWUP6x0MRou9nk
WhHgKP4EhtXJ+MQJJBotvvBfeasIRRKcyEbH6bnNAiCycATSJKB97N2OMplU2gFn
a5R9Pwig6bhot4PjBHRmLjjde+nPXc2/qddtOes9N19pB8amlaHiq0+C56J0dLGx
3DsDriOLnNqW/HkBBoWhOixcn7RUL9Sj9ZXKChAfE2UjQq6jNWQdlB8bhB/VP0Sw
BZtX043PDTGL9p9HYmSp3CPK82paqQukn+egjv06N0TYTrKqm1+k1p6Xx9tRiVdp
TGLKU2KeAPNAFFgdB4Ehty/g2n068dIJtmTuJyUb2pE7m7VwNi3jUIzdsMFoOMwi
4wpU9YIVriyzqL+sFs+P4XouZPWPrr69rIJ9lcjoXEBtxjCnKPZzweYNfs5OAr4Y
FeXHgpJW4PUA/DaLzkMuGOi/AERqx5eiGgYkD7K27xZ4cbjWi82itafKuQfjc+ue
HO3T7bYjpgtjmXosz/dGzIu6zmsq0jb6rGlFyJpjC2ty0dlsNU9gUzNUNSC+MH7G
lg3m1zmPcxjWEXdSm2am3xit52KOA890SFOdLoFKnHyV2Jb2Wcamhkw/2y4oZbvB
Gfy/1DzLxdY2LFmX3FDPN4GgWJQ9fstK1fmvMlyO7cNCumYqPrFJmBvuKMSkmyzg
Q1lAUHQw52dIGIgs8kINCC2AKLHgoa73yVo4lE/EccqejPkGN4QJF9aqGsti7LdI
1KfnLi4lIZdIZbKvzxluTZPboZeJZVP4O4QhXp7HkizgO1OQC/bvmdv7H7yXWeYH
//DJeum7wWLLa8CrnaEbQmm1PObHsW8hBkhCJETMnnUnP6dwlZ0HNg2QLmZ9wW9+
ucQfIL9vrQ47kK32l0EDydg9uXn2dtfgrOv16/lwJYTK78MoR3js7ZDF0COezr7A
mr9y5Og8FiI6ez6MrrlPtusgDF9ui2A1a7LL7YzLPAEyS02gj4j13uxpg3lW/i9e
ywWG5VGrldBxEKUK2O2mtBVfNXSiwkwRvcObAq8AmrnnlDPgp2eORHo5oGWZXTbC
A17pNos8UWdPA51reR5kO+2FQHEsxlS7FwXVnG6ZlotzM5Pq3esZB7tpPIGVi9Oc
wCmNzzjPrqv9rh3HhJzIOtk64sX62R299eaKJNHf1GSS7eefj/dAk8SqW2+8C9et
237kmqQDxdGuqleKYKISLimswk1SWkGaZS0wkopXYSbFKwNM+hzUnUFL3mMq+nud
LxGRKA6uIw+d7l3OGFKR+8VoT0yI5LRSDB4MvLj5zkzKhDrieu/rIPsq0//zFIrR
m8j4Tk7+Af7tGZqjzefITI2lIFsX2d34WqaPLnzclsTPeo5WQWPF9aQ9jvNZGhIS
UeN/T0EWJArg8F7AwFeXOlmfpbTpGN1NEWQ5ouXcieeQKQa/WLwd7YgXGRIxb5IU
0uMjWpWhd9RBRMlrr1uR9dpY7kwIV5mny/pAcTYFAJdwuxttRvb7ezGfgSyM8xiY
BOHJ0rn0YJtABTSxoDRSXz2WBwbRiZQR1m7s9tIUYzpiaZcCwDFdx1Wf+xvZkJDF
qxcrhTYh1OsGH7dRur5NTRj/Knd8b1XyvvvQfH+sHw725B07CZgZWgFq5PXD2vp7
k5hg5+mU5dQOjwhiFOiRBnb5e3a3lppdqDtcwSo7c5Xh1TEH84urK3lu180st4bY
VDuy70JzxXUHS0xTc1WFPiuVzBjR1OkYTJbEItZSpXQWcKWi0/4SOSPY63NHYjMT
fahKKGsj2O6igieYR98dv6RJyR7CGSZnD8vdhlGdi98IM8VaCR1Axk/hdWbZdVHX
wlfzM2nkhbXmy0HB14C22dbJ5kMEswNs/UY793mlyObAOhklJmUkCu186fu+B3UO
4ub5+Y2eBpgR70XnfZIKWaFsuqK9xSe+lSPatXKu0jUoTb7w79skaMJiFFt0Euoe
dPf7lr0EyqszOyw1cpxE9klktJrE/V0W1tqDI/1jcVpFOG0cvUF9+rmKtutZUIGx
XsXZ7ywbWuiAJaROypWS1FBqEoLnkdo6euXjlr/219pc4HTUyzUZbDIWht03+hPG
EeoCa4C16Lv2sIw08o7TguHqLSbX5R/wme2v75FPVvIHF9zYV/l/yX3VQpr4gMvI
39n3n7sOIh9KbCvIwH3qAIiGx+rzDSwU7Pzqziz6wuIHylGMH+JwQoWn+9o1vzFs
L2df3qbvqW1NAAC5cjnOxGa8KmOQi1SQ290WukgK+7fF5Ac7gNEva5SNieh2bE1L
zbkb2ESClEam40sprGQmO8GexQyj/9hzM2ZE/L1EuPgLq9UHvqzyYcCoU7OOhYEX
AXXZEJpClU9YvHNgCSfIqCS3S8ITVPIOOJ66TllNVXT37tjQ2PniMBWTeTQy83IJ
AfU4fzX8CB/wqDMhmILbkz86OZLEndJgf5EXnSygpqtzx+wE9CoqE1bPlS1ovRA4
mO6NLPHgKkGaJZo5nW8fxNOEt5aktYgsyOsZ/nXCPBKCf1MFp/2vMCjJHXlsdUUs
EGZT92sQnAoZOGWJ+Cnc3btKD3f3l1yM6hrZwUuUyP5tYkeXDdJg9OX6jZOFC4xX
M2fg0NQLhfu/S2QA432r09WQX0uv4FqsYPP35YzOjB1IxyHy8X2DxdR3h0VIL++o
fFizgIffyPmZg9mmN7+LKfJqXYAuN59QyE0AVvwpHoULxwxf1DToz4QtQhn/MmXU
oZsbBxfG+YySgFMMVhXtOYkkxCnWJg8VJ6BpEYCB31yxA6NC1VPmj4Tc/onFvK1k
LulTskgmhwO6sn2Bq8u907nWP7e/gQ2KpLVvNILLMpvISIUGawuNSxZifIFX13lO
d4dHutyWsYNPSjhr4bmlHePifkTirUcldfdkscRi1TE2tPob1Kf8WsrFq/Vyfp18
a+WjAoi+ga/CbQq1ri4TQL53iHA6BfLHgYxZh0Vj5+s969HdbKDloE2zEGA+ENXd
ZFcQ1C98TXaWmp/ePGFq2scuiNph/cBcu5GhjLyflaUNDjJ+r0KNIz5/el7NG0Wk
LDYXLNYojbh1/cXe5FS2aUzHPf2LcCKDg4/fJSymKl4nCFUleRduYXmSIOql9gRI
4HRYEBgXhpywMuo47j7e93Hl4DRr2yqfv7983kd0jCI5s5/FAXyJ1l7QhYLVvIwr
kqvfeez5mLUH025W2XjtZikjBTTNcr0V8a2BakBwwW1SfYQOS+TURdPxn/xA0fCI
BD00QKyHJPsbdHBYQM9wEU8TZkIb8JT16ZJST9v3FgW6YTjVaAsupvM5ZjiTulJ+
PJg/7FQdmbzpj8q69FJP6XxwsyHMCDVXJyXIS6MTdmP/oXu6Q/ZFwFDEeUFqzBw8
++t+BzI4luEsXGmeTAvEgI/QOLNhUBTVamuxIMog/4kDRgKdOlNh3B4qEadC0OvM
PZnw0QiHXN3oTi31nhCIQsxDwvQh70t6+qEETqJZRDlfze2PN75poGctuC8f4Hg3
4PdVq8PGtXVrMhQqhH/B6Rh1tKuvAZ7wIDlcA1RMldoPe7sJHpqXYUf5ChGuu45/
L5Bh6NI2rqeBZ5oeF8Y+dnyf0d1Qw3zuqB1teR13g5rCuYGnPa2Y33brfwyCa26X
NbW98HMsLf2vAHW0/nl52OMrrg1gzTiJhXIxMbxvjHGvolQ3sHdlXS0FXqHjvtlY
n66XKLjbv1VoheZ8kxMXZkpUXYhDbPmzdlr4QIurtX21n3H5IWzGkY87dEhF+dml
JYGK1h6u4IS5DkLyd98PErXfh865ssZld6AEtbnvgJeb9j6igA19Cnf5zHjn6m8o
B7+sAPc39WiO+o6jG7s8NTYOtqvrVhgkpnYuzigChAgivKQYvMlKhwxyUE+584dF
L8Sxl8DinwMjf8rrCFH8Yl+h3XygRDznTQV4HihXGs3doPUwybTEqpq3rvALQP9x
l6hGV5HaAg6dYTg1NWjgtXaADMYC2MqeyK2Y7w7C4jFkYArJxE1uG80lzViy8n8L
MIVvC2OasgAttA3A4C2VT9sDR4ihKMUcI2du9WN7S5BjVvlKAeW32L47hkw+cr9g
UJnQ7igXiQskcrwSm/Am2WQi2WpMAaVm6ypI1Pv0sq42+WucN3zQRnG4g1adt9Qn
0H7ZVGYhCfgAGKWEqWidHkIE4NDlK5KZ/ETEkNcevk/W0MnB0hbjRMiLyOB+5R2I
YdovjJeP4zHLMypfAlsvdzW7sMd57FsKjhvNNqEnMwRiy9iFX2MZJ90rHgjWGGTQ
Cw8j5HH07K5TQaOgpzgmqbOev7+uHXfqaAG30MP/M1ukaXv0Cc/UzzxmCgznJgSU
RjDW0uhaHKnEXsUQ6sz6FvZJEHZvZrOdJY/CfY/3RD7C7aBvO3ZelT0aTefLZyWG
XeY46UAjAdnVuvCI0xmDTDzevoZqPJy+CaphyMLdOcppbNZ/yfqAUTed83xIFlFI
0tElAOrPIIKAWFBlNY592zxWiW/7z+nkZ3dHSKgDbW0elth5E0C5Agna1XBwuNLM
KN/wn+5qtVJ0jPaxa3dWSsCXy7r0CzHnYbBjoIkWMBTWReSseegMwMNC6pJHayaA
axmYI9GkemTNWswHKbcy6Ms9J8pdWEoMPLSna7vDxsbN5tZJxdklFDo9Pr6NUBM9
a916uN2Iu40Dn+NacJwcxptAYvVz2hzo1151g8Lp/cNO3LqVQcOxwH4uzUrYPr7+
Eg5y0j22kCV7AUAAC+B4eCKuoliYU4o4QgW7ByzkW5n868top22vdkGGzxPjbyDM
p+VXv3qtiu9yBTE6fiErFeHD0MpW0Ce5ZlMZlVP9GM/TBgc6+GpU+suCpHWMN1Mp
zshALq2o35IiUZINd+EkrUtWVy5o6bqZ98P68BdTrQ0fFL7Dz6iWEjnjs0RcG6Q7
IOtGnyE61pgor/o6HJEpw/uXguJ24hQesnw/17CmKTPnoHjpMZVdNGLCFm1Nhzuj
kUag/66gkb0wmn5M4OtKcMoJ6UhPQiYtK57kEIslXoUsTA5L+JetNyoehMai7sl0
wteDyzPwX+uAOwlwM1RlJZpasrEPVqAYwZ6tM6Fo438Q6aP5yNVVDhAXL8uxJOgz
hCAO6La6muc96g4QBCOu23FpyYsl247/0H02ydd+KfxNT6SFP+G9BPhEXkn8qK7V
Wmq/+0W62ibJOlM/pVIW1CLwpY/R1sfoTONqjrKiWEWaVhGCti2oZEeSOykbJsMb
QMawEOec2NSEbCQQlsI7QeilikcGKdbzy+63iA/9hlkjI6DqCNOdVhmDBMxbZJFd
zTW7l28FpaH+E8m85WcvqOBnPvaEq++AVTgJOFH4+1fFXBpc6ytXt+9uIfilYpod
4v/pcKuVRf7PCusbg8vY8aLfGs04n6pbsq5wj2xv0fG4zG/Z1oS4zv2OBEKtP7qn
IMWxghnHSEs1y+XaUMeHaJmMwGqXeujbqU5oGUQ2IhpauS+1ZzA6EBTO31FzVXGX
zrsQDg3qMrTLJ4VZwm6saKXXpBCJBsicJLgs1i+nyguexLsm4wBrqJAjb0GzVx4r
sdPI+G8++KCjoTdOASlF5jDK2+OLa+B2HHJ6LNy0LhIXuwqtC2yqK4UeyMK5Ntez
a1ijotWeVFWzPrq8gaT8Rh4WuW2eIBbwWNbFHVGiu4gKhSW4x6iWtWIZTThXw5ux
M7o98vSlyLKqU6Eamp8MCfx4ibuWwwRq0v8zlaaCiWmmi+tMBS78rA1rIVvnKV26
kH7uGSdOL999HZG1Xn3t3BrUmqGdUCxQbrcXa2mcsPeDPRJ61WSTujE0Kma4z+UG
KorHM+eys0W8bXFqPdFViLQM3Nky2eFN++la3dQlIPBK1fKt+9LzIUV0tytUM63P
/CiLl4M2foDuePkUxUfDz0Nf+/Bc4GnQ4w6QfrPW7+TyuKqGnSHGTQcI1MpETeYF
4kUgS+9LROCe3pce62ssnwGnI5b0u8BE77+x3x2qxKDsZTkIal8iR7FOAb9NpgYx
fwGnQVYOW2z03zwMroqfdJOej6vAwa/qq5IvmR46IQuIaM4mZkRoTD5sSFB98GSo
mflkaql0wlLewC/qmGj0vPhRBYOdbsfPWS2rv7j6KDvI43tUpCx9wojQtNWugdtb
BxQgXydw1wN1hnLdCUEUWmqztPmVAZzwCgG++PeXZre+m5IjiywfbpfAC3DJqATP
wsawIMRUHrd6+i6kmCCxAegUhxKnGClYsX1TmN/aGW8mlcA3h4b7JuOF/OijJO13
s5IwVrHryGrqq63+28KnfaesSrTekT0uIRbI6y1rCHSbFnKWDVK8E4pPSX9eaDQf
rYoiu8ObTveEbjpVxbrUj/PQdWzKpYrp5VjzflIWHYeKI+nyMK4GBsOOfIyIlXMS
VSJ3rCodnOL2tjA85C/pqJiL9Py/YLTBZni1l+7G2f6GZg8QeSfXrlpLbxlIaQAG
CfhWzeluNBPpcJ4wre/9RwuQoKfpSmTd6NwdA1PfvmAqkDeLyk9kSYTMHNUgxUiW
X3upm+KjGTkMiEOsRstY47i/mLvmcWZO6glr5CmC31WMOuU96OAWed6WkdSuPXNM
pg6DPavzSbLtU3Oz6LEBNZzk1SBQTLy2z+KQy4AaOA6+Kz5PClRh3dmyQJa0JQ+V
OWNy7VrbxHLNRA0rKtonUF1hiar7O/37CK5ktZTBaHtX+VsuPcMpqn29x37dvtap
3Xpmi3KxSn8Pl7cn60pHt/9PUPkJmT5Ig/74oIKQdHab4VgClPGJldQahvSmYdAF
u4VNq/BhXlwv5I/GGAWpIUR5vCJhnQPS8axThJwUALjIRUrW2qBQpFCHj/FeH00Z
S0XE1Bjv98BfiSlMeMkzMjDnccBO1TXFBOvHD1nQ/BAY8JaZ5aPiGXadI8tSe4Uz
+I3/yVLVJ5DOCGbBb8Z9PMlMikzN4jqOVaaTVblf8C/FBDSiuhyJG+oUCq2n36eT
I/YTjlRb347IC5dXnIBTQHR6KKu+QLna9EGj/UrElZYLROKz14OFqZTTUHfbZIuF
KA5nG4usvclgeYLBCwfT8C4NGkQdAU72bdIKCDQPIgkUSJMm71tapuLgFCVyW7/3
998GW9KTEUMOGJFhhzgSeTvGByN+UFc2TIjuoIYbDhlEq4DcISKa1ZIsvV1xBs16
Tj7EaHfTtcGxV668ANn/J1p4Hqz3vKappnC8XUZSMIns6+dtJVZBX51CfZD/cT3e
xlPO23BNULdpjsKxvGNqCxsqe48X52UA6nsEGeV7/UEzyNfOSPTIYFw3sngDaSv6
PX+jejQj4XysJBGGGVJd5AqKqyVAsPFlyaVeBtYt64qa0HE1otTJGbmrHBslZk5m
mMCpTGxjhbkSq/wqahA3ElgqTAC352s5q7qL88Yi/sBKqTDjGlCAMvtEYs7fS6VK
lyNFEcG+spe7pHPQniQ1AuYqEfXWqVh5BlEGPWjQ8wPAbDFpbBUH7JnR1rI4ILvO
Ous/jqdt8RzW3kZO6U4XoeidZY6X484Dd1N9TFtRCfwHKOQHc4qO1qzAqExiebzl
TD7MteqSRwQXv1epsKJxEt+aLznlw6UOSu+z3/4viSlNNuUYNqRZzRtNc2Vh1gd+
7FRoKFPT0sDQp1KCtLN1H5WqQu+kJ0MJchfa5Zk3XU82uNM4odo3Le4Szt00j4eJ
JdxGMxB8m8jrA6NLENTwIS3/hDqNdf0L8Wc+GZ0zLD1NTIUmsHy0ERZKpBqQtCkc
bS2l0QExk++zSeWvQS4zcyyeLrswLD3ImdJThST5EZ9MesPc1LZaGR2c32V3jcUC
bRjBBa8EeGJJ9rizgQjllvFRSiNnyzHr57lvB+qtUU34u1jXpqEDXGc4G4FsKOK5
cGiqxKPogQ2bzqyikTTTraCSQyiFtFE3MjPW3r7QA7CvED9gbuCUBL3uDG3JxVVz
L/2XXTpBz4ZpEcSvu2+ni2YLY/fIxRlYyZbd+v2psUB4z8o44fIy9+XxPYiF9xoz
sfw1ZSRyZkU7buzzkO/gqSZMEG7S1S5sbzT095ftdqILLIk/2USeGe2L1IkmQ9zT
RBAUeYijHgILNpMYmQWCLpxHLXFJ9+Uux9yCV3nhW5b0TobVWWmQlg9z3wz4aE6k
dP1OYt0mw1PMOy8PjHKmJVKkcH/oC8oS+pHJxLIcnWblRwrUUdPGgZdjW2xUFP6r
8gRd1QfGTA6gBkIQsT8oV8cCs9ckdDoeD7LYTJQI6crMy4YlSPB1jKau8n2hqDzO
Xi9Zqx4R5pa8KzOjnfrRGkTafpH+n8BYsKQPPzOXATVFtLP0Ekzxz5xv1wtneLTM
nCDAvUd+OIgfAi6JfmPKlaaRS+xjPzA/baQNlS6NqaCPtVp5TzDEB+jFd61iDSBV
18li0Z+7iDCKsEJ7NqipXjPU7c19mqcMoFsc6QBA/Y+sVD8ZKirRMwR2lvClC7TJ
PvPFxc1IhCNPci/TWTddM46EQotg24wODdySQUn+Zd1sp4zOxf+78cI6ZXiKdIs+
fRI8FbXBJokprq1nD8JBgmI//N0rvRkB/EXlCNwhkIdfI86+oU+3TZCdGlQdRtQ8
DbNQskXYHswtLREiCAnbrfiCUWAV1miWJXBVBG0AM/SjXfkgqoHpDJleOAZoU+Ek
5dZRx/rUXBH8rcYZ47LPhGZmST9kPT5luHS/6/nvLNXG7toDtEK1iX166GTtfLAu
Znn52KUIUXKebFjjsMZipCx/Qxp7Z8WqUpOwqnPkGZlgGPfDuG48xHXnEjEXGOM1
ECrcRHeN0VjBZU1Rl60UaLjoOHjBJcp0RCS08SKg6bt7BgWLHsjP1bp5GIyOsnp5
7Q+2hADqpBcql6/mMxzHydFtEtQ9ehEZ6eFQ6LEsJTrqVUdbkjHWNhu72UQrhGDe
fGb1qaAUjoOrUXWq/sudUNfU6pwpFm+KrF3i/Poe/EDa3Mkk1DnwpG8kybyBLw/R
ZXcI7LEfLTKazfiNTgQCDhaq+BrqZe6lYfMucob2OYI2Lhph3mHCwxQewEn2sNDU
1bfggIlJW8vTjtLJTf+4V6Neho71AQKiNSH82jiqOmwhCxvUgM3vtCx/RNdnyubg
6gygdKugyzQQZgzoljfC0uKJhaSCnJIWgXbqYihZn875dn+Ci9VyHvswkwL2VewV
mva6unce/W9NlHyJRMvF+ar2Dw0j0e5i69G0BH99r6OOpRymxrikZlRj7S/Jz/m+
oKDcegOII92KEC4JDFQ/yJvqqXf5HpasJ+cr1tQTSwCUfx3SIW6hSabQ5nryhBzG
7QDTiTOtekFFM7BJBGUA436t9RgI/Fh1J8wYxjtuYU8rgSDzwRdvdFqjVv8nfnQN
xfPBZ0E5OANpBLKRKAg/z5JwmpjkSoG/Inm8m6huNSWuGCjosIFQu5Xmt09veXkn
L9eDHYcZO+i1EkZdhXzIIUJslHYhe5gdX0yMGu2320xOck+966xbrZ9pu3lOBd5K
R4f9JPrr8A6ieP42kYkNBQCk/ZHuzwU8Vl8dg+mjEYMlMS/KkQENj3ZTe7dpWIqA
MJhrzx3kz3iOmc6QUxiEHaVdJ1tSQ4bXI4+ivxeVxNVOnwnk2qaejzFKJptHd53Q
11gm5xgFEES7WknE41R+Jz++UivGF0VWY63uawiNUq/mPqyV5S7DQpcqx0aMopsN
cf4LVkmyjXBMIcDTb0xVpVt1C7pPWPpewcsU+c6nxyiUZGgVsta9/3jPrQlmK3EO
Um0IGHDU+yW9+StM53VeuS0hqb6P8SBA6I1RnzBBXjDGmzdEKdHcuA8gcp3wGUr4
RdgfKry8hVqN8ukzyHdacraP7g9/svnD0mVmG4EgGLv77qhjywbosPa9H7RJi4vh
MwwZr1VOZH5ReWxJE53Z1bF5UcZPRGDsop4Qj+qKC/nIBSqQ/Hrn+Y7jR1Ckd5HB
a9geZ3TK0zK5tArEEY9OgwLBZHt1WtZpWDiGA3mbdOUeSB1l+nX8pEcJQbKg1ymr
jhPcx8HfzARHIoq0jvYBZAuIf4MgjQ9seqgTUG9ZOHzs9agLQXsvSLUpuouYtXsY
5YTKOlrlhKt4goYA7Hkv2iC4PJ109pme/PSL/7VIhT4E1IYL0MaAFieXYw6IHh7S
mJ7Dyfm+Dxq2tjg85seHioGkr5W+JdyGXmYDIWk8PbRHE1LTKWJXyi/LbTbIoP5L
I8/fuuVqRQs6XC52Kghp9zK2c+2ZnV4Ycla4/0kXdgJblr0TDBAVE8OsNEiA0M9k
9jQkWbp5tfnUo8Ave08seZJraRCkTzb8dSNU8wnkTP4Hp3AnFKrgZ5RC77GPbt1y
7yMYsJUGLUaiGknB+7WuT8V4EJS8y12Y4AaSyiqTxGUtu6RGLlZPG3Jq7Y2iuZOv
uwCdjGHDXPxz2VdBuhRObaaT4yaz0OkNx8F/F7yMT37tjYJCFFbbhKDSPzMSTy/q
75kL/bU4cJ4KP/6qse5otOBT28uET1WDJdgeT5QmfhxN+vKo+ckDDSWBZ/taTu2j
gKI8FA8z9A9IuTx1cRz6sh+AIWU1kRrxBOUm/m6YrogJDNVFpRNTQXB4pmpmr6i3
qNpGxEtEVy+BgVFvOGTEQk/UFLFqYGbaoGDvORx0ECd0gbU6XePWEs7gePflkgdj
qHYHCfscQZ1wxuan913pyJD/rea5YJqHzYWj4G0MZuCavjEQ4E4Hd/f17UaEpzyl
gkaD310vIAid+I7YM7JBItv4cqN3Jemflj7I7J3CuNQCr/+zcOuA5EskAuiK3PjC
qvsBR/CexFKNW5S0eHVTTxhJ3Qu+YiVxFyPvZEcd4StLo5N9YD3hNeFQR/sUGC8p
PyL9/Xnt9UH03cWL1PMR40S91c6FChR9x27PtHHKbc2UsqBCtGjG0ZlQrfL738Rh
bcPXUcs/dLYJB2E0esW5o2lFm9dD0+TXkBx4sm/82ULknE96aXDSSpFnNnH4+bUj
NwDsFziP1iQKuY9zgrog6a/O8ftBRIMfQ4y+J84szzwdcVEJaYTcS3U9Z93aWoQS
37OZoUSPN2vUKGKemALFbOjG/yDMLRyKoFmUJTYNTC+1xeKdGkuKbdc/HixS5XZ0
2t1zRvlt14KkaogPqdQnJeH+kUKnQyw5dKEg+h5xqi7TDymyhDXi8OuhoIMMkoLC
s3Aatx/4r8F29NW0LiCpSzj27ZpkT6PliPeX1u5u6rPoy6x9T9sQwAV0rUTgasJZ
crlf6iyLY3w6/9JfYuNyYlEDp5jKcOVnhHBJk5BAs9CV9K9o2oYfaBl0PRNiTLHr
IdQpwTpEA8gsuU5OgZOiOk5gEHlTaUMzWTvK8CceqskYaJoLtEISWBXE0sARZSoz
Vtuu9kjnVHpTWbqBPzOmnON+d56DEooY/+1xmvnG44LaA7MPNzd8FlZVRPdmlBq+
o+0fU7zGcKse7LOHGSev1j6lNLdTXa5ukhe0uM2xJrjBBlVfCPTkpVdAY5LM/P2w
dfw+YORgjEHmrfIdR7JvxwwYNbrvUEo+GqbKVaaf/F8ZTSRgTP8qRAt07yi+vr66
S0AN8c/PzJToXOgeHWTgcodZUBKIcvYwUyDdaIFCQGzZRdZPU+vnbnugnmu4oLHS
xphfdvEnWUDwzQ013lvqc1Dn4Ka9ayLYGnCaWlOz5A8LTGvQeSXcQM3OhhwhBr6I
hy5hRBgglt8hp995UwYL1izakHn1kjuXNXBFrNa1rPyCZGIDk88xgbRg8lKmvO47
wmhgPiiA2oyDnH/SBqQEnmaM2+qzAbswipl5Tbfl2rP3Bkvp43YxNrg0HkAtgNYc
mY96YhBXav4bAEOBbQQ1lOnYLwo8CxCx8FFLus5dS50EP0Io/5ac9vTbejVEttYO
TX58fB2EdWpYxHoqAowaoZVX1K0vajyiX15OJrLw1rhVpmd985umXYnseoO0pMGl
fBz29S8gKACgUV/+vKpd7bNnxTnK/d2GX72MigguONImmwuG4NQe1YTVG9/AjRDC
OVMESRPGtxNcbngcgv8MVOWD16/JiMpE9eJDIwrcaOWEHS0Q+ocvYpAajqbN1A47
1YJLxu0IuL+c7gCBaxzRhV2+K5sNTyr/64qw7BsDLg/6BoTmHlbF78MjjltWVpHC
uk6nCZTOYA9T+X0DNBEeaQpIFHE9azjQ2ZwWAanDaayQqSPF2NL9IhldzyAPCUEp
N1up+GeUbCX7viyMqw6kfrDjQfLhRB00hOBkH/UESu46a53o18+htIFVOP+sZGFM
WxbkFenUhqfatfvM8zp09/BLlahGeq6HgcA7C1ywQ7XlYzJ9ZW/Vn4ZuelWczuQF
gPGK4C41pzdLKUTr2gcBRlVY4cng/LY4BfQhRj+PB66NEUTh4Zor1y9wAPtsbHMH
ClkNZIXmsFESHuWg0KU1qbLqSAurEAOUqZAp6mnJP1+J11bsAPBUrjkt9Pdcpy6W
JFaukmMM5QphGWGkxSIba89+BWnzcTRy3xlDCik5K1yXMnedXQQ1QUWI92CEbmXl
G2EsOj2ywTHkDSRA0NS6ogWujYp3TZVfqfHMP2/PvmoTHBqxvmK5dV7YjKMCJWdh
AXl3skWKAyOLvFzNG2TjoD++6Z10v84fDevq2fTduvrRL/anwmabjgIL4dA6junH
xWNQ5AdrYeiVF9edFAfFfR/CMcXKFlz0RsdJtK872y9ytKKiM265XEo7qULwkVaz
2UpE22XTTs2N2XCgyeuBKQal2EyNDI7Q+6TqGwQVC32BFdIw6Jl5IVWm3Ym3yrPU
hR27iQACz60hSmlCe5IVR1IbLqFtxUMYJsTvpRrgJWjhIElJYbqFKLdPqMjI8QSK
s0zMNweYBp4vvQMQiLT9wKPvu0jOkVrp5/wuqIPboKN4wkR65u85PAC6fCDXRsU+
/cVnjkhFuWP93NcHbC6z6Qf2vSxa//CjXDOI6C80ZzZimSmFG6v/UlY53S23hwcp
q0M2KtYMTmbe1Qog3oZ2LmSaQVMBV+fCjekvXiN90rmiZ8+q1I2CJJFC188AfduM
U8FyaXNpf4n5mU1PSilh6ygIpxxotaZuiQ/SNnbUtcEi6VCHu2z2sJ9RmJWrpmOx
+tCZ6kHP2nO4/fvNCdLa2wtPR5QMGP66grsvhMbNLaim6+yAkt+iFsJgTSGH+wF9
BhWXZUXmiZpoPrTLWq8yzula/z9kmX3rM68mfOh7XSkYEizCYNWuAx7rPDupNcIj
rFQ1nSwzsxSQ7QYPvtYOX2ccV8zLJt6yrqXyLaqbutBm7XKJnfxm43Tk4eCdkGvl
Nyd4RmvS9qjPN895KDTITytLGrEs7AbEiffG8LhpHnE62kHiymYuAP+W8rBMTHvq
0h/wApHrFEuuZVepuxCAmwaEK1dFZleZfqp07cwSxGbaFDHnxmtK0MkScp2CkHSZ
gMiXtCuOxs85xTWPbPNKMk5bY1au7xidRRjZbfUkweRnCJ0CaX6Pk9lmY3Y6zeYD
ptZaGTh2AxR3DNFCmUWqp38dBUPt2JCCVn6l/YKlIdirvn/fanZkjBmk/ChYeV1s
tGPdPBIwvLHg01gtHAkJyo/+EJ805AB7F2N8D3si2jMZ1AehhQvL637XXWt9Iude
ngQyHHcdqM0gCwX9lUz3zAqIKetJQjvNXDfdoonJYi06Gkvuw7SOeZUqmLKU67RY
9d5h3zrs0IQuFNd55rej8FYwFMoqmMO8q9o+OihrUh7LIh//5Ss5oxvEYIUbpy8z
ho2MFdAyVxPOJd9hYHATHh1f9VGCyBSWcIQak/JgehSRm0n0AmMdS4pabJUG6vRt
5LJ1pWaW0xa0BNZFLISeHPp104xLDqJEAm4wV3mBvvYd7sXcJz4mVK0pKZeTwb9R
IENxoqdVQ1lvZvnY7ZIqov69Kcf+OHVtZyTG4pYT6f8FU2tvt5HCa8AaUq+fxBPh
ka5QddHjuiZ6gXc+E3TSc092zItePW6e1/8KX03pPtN39I/keSTYMiP64u76D43O
bxfoXDPPX41UogCzZJ+ea7AXEU2bEzbOYdcm/IGkakz4khVHok3mJMT542oanDkD
F4Oz+GVtiYw7GU+bFGrn2izoY/yeXl/KNNx95jN7dtS7uGrJhRDBW/PhYhIx4FMy
sBSKHYS2A/wp5e9ra0bV+IeAk9u873n+PDBzJ+n19D4Vx9WjFxgnTr3E95E7d/wR
Kx0QqVxkGFuMkIHiJ2uA8uzwv9BBMxIiPWEdIAuYAJ8EksPPrmLXEr+cAgoISfFc
9V8AzZzyHwOvsNXJzcA1eyS9LPXFeDVYETx2l0EED+XfSOQaRk51gsblNHdnBhKq
O5mYf8O1oPc6pok5j0iMVogpTfb+z/q2Mdt1fbcmX+DlCim8rlk0DMXTAhT6UMtR
EKGORnHgQ3DNfKq+O0KV2UP/B2ht4DoYJjZjHxqXHbxgg16CWI48r2vgQy7WNQsn
ekG1G54CNygJDtMStrCfgCAHmLwA7orj+KUgLPLCfXwcCqyf4rMSJfXR/IiNm/vp
pglyMmblsH29xdJ/LLSGyIuQo2u2elL21Xsxu1t6/0R8vcMYJl+E8rZ2BtD5AUcg
FUd3cL++9g0FozUOHu9HnUR9Bk/Z1IKIq0LtuZmHzyqjcsAYihznm7KUl9ZNq45D
rqNqfwSW2TD6nCneVC8+dXCbnuv3UW8OfzojncQPCY/X0y8gXFMoWc7MY1rCKb2F
LhJyY2716eKjpKAOJ1QA8EEdSzREWM93gwlg8gJv4CESyuQ1SiTF7P5mFTnhKJDV
wX7hshnl++zKElZ/tR8AZ7DotREa0xBYhvTXjZz+lPtu49GhH7cT3yWuDwUabuEc
wY44R9wWelRq89pG3YgrDJMB0zfcxUSz4S8f2AyFi17COuEkO86HykkdZkFSAW+M
kRN4wO4TTKjXYjQX14vSKALdeXVNnaSyv5fm1pc7uSxfAO3X/dVnSRfkgo0riPXW
aSM8swkTgWB4A8j+X1Idyed4Z62F51a5DHoUlJkpPaKyhREq8G7Yr25qvMLwQHeX
YOHpV9mEsL57sBcURAYnr4OuNgljgmE2h2M1ZsGlocu5ynxwDck0Z8WKqUxE4KXw
iCu/VJMiLy393FWQ+fvRe2xnAMEh2wrWf4QErTtqDhOGL6KkP6zIwm/Sz18Trv3i
BPiUhmxm/TtlxTaU/kqzm34lMxYV4h6cpvmu78UbhKEUni3auZGT/7KMK9xsotI9
AoYQT28W9odulvWCezJGDf5+YuK41FKWt4Y3OEZrO7Q+GI1cNpsTX9w9kEIJ4K1H
56qKP6RUPw3A/NxvJ/7jPD56pV8T+qYSkG3HF/4D1nQ1wgxhwQGnyW+0og6wnXEt
ywMiV0gj5LNy/IP5rAASijSFewtJtW7CB5htR5Qjagv8Sl5fQFQDXiMJ9mAyP3/l
5uGWvuK7JziN+NATkRsUOCs/3Z44ndv1GBzlbFyGq9ZJGkrtC3hNWfakyE53ncTe
OUbKf2JnEB+lmXN72OK2hOCizxYRxoahk62ixyIVS05+VQRalIuLgoSwPi4AobLt
jcDQHJq/hl9MXlZIl7isKwaD3r/bKKKrMHv/gFWNdTPtzCxqNJX592GMLoL3c1KF
sqolnHRMVfw1zcTub4ThzcPP6M2Co4DB6SpBVNdWRwrt5mEWrpp3uuYvpkvjUIrB
Qaz+ReCP7bVYJSrddrLhPTvErzV+cZcdnmYaIyLJMm54egKYmFBzEPPbrwmitaYr
lXOK6MU1Iqb0vfBlR3XfXJXnVxMGqWMqc9nyNzaDAKVi4RGZ44jXaYPsjuJvXCra
tyQ1W1PwpjOHSZT287MzWmp8ZVJmqHB/3yV3zpBkC1C7r6QpZSpPxwPdvV+k/rp1
W72tSPRSCfQHzqLdt5jDlYhO0jb0lY2Bs5gW7ZUekbMuGRQNK/9AWJYXfFZYNCBy
YD2vBtkZBUEDsS8Cq+cZZUWHUWyT8pYiPnMck2UWRcRVOIh+cj6XB4X2JY3cG3E8
Gz41wNbmEjjAAJnp1WM25PygCg4gtAH285xSsdKFF8rH/vUKlS61KSkrrwRCYhyZ
1NM3AMtcitBMOcSdLy4Vy/OBMfT/cGh2E4PiK0caepa3WbrtOhSIOmEQyysYHVpw
+G7O8vBIsS+FpPB1vVMyewD1DyJ6noM6R93Fmx+8HqSUz27Ze5kKUuHdW8/VFAZC
z15R5JCrhR7DVwCkQHL9b1SNhnT08PZLarDZee9spkBDgNdhyiwppVS9upJ6Dyq6
8rL74bKNoHJgEWNBDlBk8US94Zj5Bd+WeRLfBnTFuqw8Mw67rp7Cuh4aEax8mz8M
sa1wxGpreacMYg/J7UlXNsO9lL98mElGU3aWmz6p1Zgv4qnyFkY0NWfLnNg+sIUN
NctTf+VDuPWJbvTKVFWDPuonnxAGLs6XFAhPZ3VucG+F5r+BwzkA/TnwzyJUC9sw
TfuexzCYzzlFfngQRSAUflFKD2KNvr2htl+kQLiaZzK/MSSozOSldnkW7wCo9S9A
8XdJVSMaBoojMj7rbk9D+8Kk3ORuo5wVTEnVIETVVTfv3zVinxf0x3rIclLjpD9d
Y4MnN3iXjdBqDiiUS8PBjSseftmP7JAWnwZtytBpOw9ppZPklq/eHPccGcaESNxw
aU0Eiae8bQuTf0qWESLU7eizPt9ivB+OzAnO6/GIo8/V5m5prKGtP7XUG3Svomb1
t1KiImmJRLwThgsKMNe55kz8NubaHg+uy8wMvRJ1Eegle0f6hqX0RedXeVIWNO6K
PK28eRRBDsmo6L1l2gwevGfDOM/JxMw27s2DMdvOspV/yKOFTohrr4j4Bl6klf2T
H2YG+LYc+M/mHxPwa32q2avtw16WJinI/sOdeeBQzF763+BSgSsdJNkLPEJPm2gX
PaAuLsWZHTza2GPsAV9LbkJ+N7VoA3U2zr9G4OLaw264FxFVv0fOGNV2SUCJ8CYZ
NR4TY4BeHWld5EkTNZEwbhKK498XHRxajSlG5OjTuP6/XszkKtzLPIHozNvnXla8
wenBauDM+J2kjcAaYivWWKVWduGRkCeJig3cD5Nb1UhK+hXAdcVfJWJ174Xs6cux
ek7vK4HUO25WbQKpEm32qCtNJqmKZdpRODmqj6k4FcC9UNVl/uUEgGmFbG1goB3F
bk7T8EeOODui8XqWYinmhxP+1c/zCC69lwe9XoVklHhVYXsyvVkocrDBwVbFIJqv
eTAMOKbBadzMQ3J/Bt3Tg71I44Qei/pxWseVqZrlZO4U/k7dj7o8w3Yhta5VIeXZ
qiWp2SEz7g0VwIsDRTLL3SvUw+eF3I4uGjEs5053Hv007aMBsiazjfkzKnLkOGnf
1Ootlp81UgsUfjsu0NQi2n767VPqkcqpmsXWisM+0F75sMAUTpGhKueOR2fnLU+B
B+HBOUHPnzhUiVWWF3WpS04LhAYIDWFKl4UaorvZDHbSIEPN4+P8BItw3OWO7kLy
y5F99IJORdwasIGSBIHR0v+kka146wbl9oUfRvslVFJqtEdx6z2KFLZ26JbWKx4P
7puMS7twqeYoI0I/AiV4PtU9rwMvynKLLpNdpV90Usz4XsciKpSZUubYAAMWci9v
rj9dVX4xJA+V5im+HLVh3qBwA/GnWVkAlvMzvoO51QiVCLe0fWgcqcQbGDHuCucZ
bw81KW/xeX7E8bHFjzag1iKd8cMst/iOBfQyYPryviVSXgVnQb3P3mwYPsMm8gYL
GV1nd79AVZaXNYrUxCdZicGp8IiAPXhBZZwMyYaeAPci/A9QX05ehE208RsrYNSc
4MarC9O31xQDtyR6gf8dvd9EJz773FGxIHWuWOktmTubWXDYsF3wvN4PC5ULcw//
Op1tuwkwKi9DLuuh6w+uNExMD4Ptg3cveG0qUYlLRMEpRdTfukg39VNQ1mWtClte
C/HwB4KzoqQ5D8izPM3AP2L3tdi3nC0Z9A7raZO3vwww7m8JDxJ5MlSbJuFGALhQ
omHi1LkWWBjdiRF3Y8KxJlBsmd+dPeACVPc5QW8qbXyIAbaW1kYDmrwJd12abFH0
C0A7SOdqdrtbRLzgs+P8EhQdhRm4fFhN9AHtMMpk2CeV8tGNmobHOLSWCFQ44k0k
eo1TxOpA8Jy2j/IOSenAzGbzxJuNDq3RRH/Kyv9lUvOU4sEY4ywaY1p/f9wd+4Ti
NfaAetSJTW/tYD55r3mNr64+eLLH0NCNUngI8Vgxm0nupWeM/0s8twDT2Ym+oYPb
jp5xpwo/nZOI8ZHVnje3iKs1Ra3UqOMjCe0mm1mYOdabUHRMd/hSjCvvmeZaMudG
hBPeG1jbFCVy3lD5qyiIDQGY33Hhfrx7UcYS5thhC52YCmKekO54G43F0fUq8Yl9
1GjsKBXhuEPuz0GfIZU5MlDaAtr9OfjkZRaZ1Ab/KmbBmf664L67iHSPmn9UiZNY
c+mWUHCKlCLgndlsS7V/Nj0DDVATlxnp+E1lEG+pFwiElMDCexOxCl6Kv7XTW9wF
V+BB2xG0DAOczACOiCxnE1vMqiZBJ+cc3JGn1yv7srbUnwtEdE5jlQ34nBWSIffM
qwXzpaSyQXHnuwRseKfpGtumbLvZQZDLGxLrKDGloMQLS4yFIDsNOaJuMThN2Ka3
ecZKafmMkVQVhoKkfEsA4lG/mdMwM0NOZaN8gENejZW6JMXQxJWeT9tipFm5tVev
EhZ2hk1R/GRvsO44TxRCI1JJEDnU4M2dQggSUE5NPWcSydobXMvHVMeqszjzNUbs
f9q4nwfngvKTR7zLwTldsr0VVERIjjR/HknjYw4v0f0XSaTFYxSjLBWeGBanuO7c
F2HFy+hiutBBdPywlz+GaGvnwtL/u0oPbxaD73hXzugijgNWqfI1QO7SgGsNnrFh
RaF6iZHri5ILoZfEJ7IjBptG8GhiTtLvmZacD0GU2fL6L2Tqi0nmr2/ETq5xOQWb
ne9t5nvHuZquiviI9LQSIWzHKMO3yJ9VFwXwTmmGKtIMgy8NaBhMFJIGgtVW/zhr
yllTZnUSc2KcpqNbnspfWnm0QxoJMUHIHbJ3AlwNye7TGDReZfIlxbmt2mH2S7Zi
xt1ZzabAD7Pris3//ExWhyh87FBpbS1m778b1/TkOv8P7ExwSM0SV2YhJIlwEBnA
28X9ode0+x2sv4244BtKvyXN/W4O7GqAfRwtz6aUzw2rkacOEKLVXA09pZpiL7fM
U8zewStHUCullmHx2CF7arZPaoRgoxSLyrEIfcYhLn6+GP3bdeSFaOurKO3nQjY3
rpiTz2GkSArBCyUQXNFedhxwCRfU8rkjBRSaCh5DcT7wPppTSPuKp0e7+lK4SPhR
4M4l79hQorDRSUwRjheCRkWiaKmR9H3vMnvhvZOlgcvyPYSYTN697MKqG4NOb2Gq
5vQyAoKyS7hAzI+2NDSO+K8FmTvC49lsrOUPf3RFWCyvL6fntsxTwruqPqq4rFUV
yDimp7xriJMxF+c/VRU83kQ6fA5sRV5U1lzAkPQ6ViJu1MbLbWBMYUECy+Hcd0/q
8GVsIjrl88yLORm3TSPs87RaCCc5rpXaNh/Tcbnbs+j134n8prxaTy+qT2pRue5u
aBH91em9FnyVbzZZG7t/H8ckhApyTy2xLWR4fDrq3VVUCq8n3kwhV7qZGjS9BhJe
GV8Bp/vcHSm2B7C2bj/F8sugWUTi/NUlwKbI/LG8UcIRfaSppL0Sc51om3MfQ9GO
0n64Y0KNBtUoD5ynGE57hQBx3KNSuD5fW84pVd53k3fyBRmb3qgsJwFhMSYKtX/G
NrWR1xmiVLYbV94U60HCG2u/ZWJ04M0pqSvYBnOvNT3UFXZ9wJofH3rsZgeBAxtL
R2s2k76x0yPnC77BUy3ns5oCpg7ke0tjnaRkBkuuKEdUSKskO2cPUFe+d0XiSKtr
n9D/nRGBBo++1gnuP6tZmcwB8K/k1igBHINQuzyTQXK2ZlxSDfYXuWc7Xco9okpT
HMNIc6wMNT4WQFkxJNNnXImHHdcgNEfdzUBTdd4gcshFvbDNaduG+4CQ6eAG5dq3
C7zTB5y6WiPOO4El0AcI1N1X2HdKFg8GPBgwb1q9f98Rbl55el4lRIxH4FrtTaus
hxuv7Hk0zkC6n6PBRn1r9+dkK27W9uNg4hp2qtxGtX+UBFJRiiXUME7gl2Pm9uR5
clgkLviBTMmAz0u1Ufh75rjZd3Sc62MbGE8FyURi+pJFIOlbI1fCvp+K8949mxx1
DTFdJ7UVpJnw8M+cD5qhMP610VnH41bNrJ/Tr2bO8IeQUpxbIyZz8jz8ppsPD8SA
8TaWpF7vhv4zapacMWkwLxx/aRyaeV/9UA2n1yye6i+wNtLt/na+SVDb4h0FTO69
7ldsKK8VTcAdnPZEjx3QedQ9K4GNG/6t/GZw8sMLjwaU3cbtqpuUx7a/Atxx/WDQ
uzyw2c6GnhxZUXtq+Z/v42JURhK5eodWt0LcklBh1yjnL02uaPHam7FEuBaTQ46z
Ort6IBq5cXQkKWiXhehbEnVxsDLtiFZpdFVNIdK/QOfotbiNgkLvsAgTyjjH1SUk
x+sIpDpJZ9gKkZ6m2x9LQutm0VDo2fkjmUvLrQDuGLUFdoDZUXr1EzNgcr+Rn+7w
FlPPHGg93Jj0VHYe44D/99HKGmsMzfpavgTjDGq7DMyw8s8FWfqGs2BNoXfW1goA
US3HUvASf9Xd6NbaKkDqcbkRDTK4WOQHw44gxr00bbWfAIjDWnq8TE0LysPwCgG0
vqJb4my8AlxEUUtqlLED3m6YCm84dXQQKIpzf73ojOCwJ3GPVJl4p/OIvEHPSnne
YdxbJTANraS66TK77eqOz0lnrz5hrkEWBO0Fhok1PDfRTZjUfjrVKM/0dppCSEJN
HjvQ+yl/GpUC3T23bNDQGVJ3J3LI9JCpHUkYbnGVI44umJMMRNtz3uq+3j5lJjgS
hVGZwSI3mvfU2xiyvLyn3Onhyx71k84/JBh5gikdHXsEipJYboBiiPKMMGYv7Y8p
Cutq8A+zoIYwQ123gyW48Z8Esmu6TFvGjKpBqBTCcfK/SXi0uZFJVf0iPJcHJcYJ
/ewjPtqd+ms3O8DEyUOCaQ3V+3C6pqSeiU8MOrzskPyNo6kDVclCW/1xBSQ55vxQ
MV8HwKBPn2xoW6sHq4eFQTeIFeSctzKznismyPku7dcnn4VzOW3ocAbxnjucev44
+zbpaDJy52wuPUh/ZI+9AwRrQ/opuCuUx3dEoxctfHRos6jd2JeF3awo84vVPuyn
a4th+XMMCBmnDlO/NWSm3IUykOu5+PE7kIzMlLgztHsKeQMpzhD4CmI4H+YCSscT
OdLpeClr6hpj3hMsz1HW3UhqoE+9NFxFxFcKCs69GCeAEv9iVKB6imMlUx1z3d+D
ZQ1xwTby3oF9E2wJrmM5uHKfZW3ka6179eWFzk/PgyDqiMRJGWmERcI59WNd+17X
jfB4Sl7pFzGt/NWnAm0fCLPlmBKrpc1cGVe5kRTf+w+T0WFKZw+EunKlhlOERZJa
ZraC5s3ghGIjoOzP8W63sZgSjKwfF4h3WkxFIfNSq9xbJ42CLPpSYi5geyTYdi8h
nq+qVxUzzMrbxvVHRgAumv4s/Y705YfJ8HYtmnsQ0ULuy3b2GT0YFl8MOoAnfmDl
FanAC5TWWz8zW4Vtl1mIV+Z/O4xFv6M8DN86FFlJTtL2ksqse8Ov8acGNBsIqRag
eXKMrXImHrEooY2+wo9FeRqzy0MY8untYMV+H3Gmsz3edrtWMnvgE8aNqU+dtz+R
h3NTlwdFfr+CEtgRU/UZtZ3lMiuT4EaMLkZ9FUl5b9zGGPNkgja47G8CzDyGWGnm
YJ8gCFQOPL9xMbt/jRA2+KCwdq8BK2Dq8g0OA6OLDLCPQzfXrQDTciFuoW3biiKj
bRNwPZyp9Bbj1z/ilAfeCI/3BQBwXHfzQPMKSB7yALH9z/i6GDjwieq5Er3MYJop
nwF346ipkVbwICNo4KKqjZfmplD3S6IAHkKcQWuTEvZzckM5lD1hXBo1IG9S8c8I
jwDvFl1m2TzirDKwIGxGJvnEvyKlKdhSQ2AOjukVSFYT0/+uAZRStkQKlG4dBTdH
IdF9S4H7TXqzLHyLw6cQnXOhUy6xu3sy5wwftpzTFrXhCVTGPiLfQV7gw8OCROLt
db0IySHFALgMZn3FvZSDuPj4TX8zp3rlP5tsDlWmMcEuMthFITQy9zEeZbjR5LkP
yW+z/lgAmckYOOkZHNVaXuGWc/4TM5TKgUn6Sr++CyUYRtLKBwjVHXq9clQjtxiD
+/VLVbLNqhL9bm0p/en0n3vrGvFIYt4OnniNzFUqSuNJicPwXLszRTxJ18Xg+svK
0ctdR6Mv3qHLMiD8Piwxn5Wf/LppopsRZzSgU0dkv2wGH6p59BLm4qEbmRkiREqt
4cNpRpJsmgUP5w2XbxaJiPnKmpRiRcbcVt4qiu8Fi7gC+cA4ldASXK8N3YZjJZlN
P5t+59d6GGcbRwsyZPia8eSYA+afqlY0IUamPax7qXBcUEx2GkcXrd6ehnuXewnu
d7wsFME4dPgYuwjmfNQLCVYd+1maLMYoDjIReSnAy5b9/cQpNYlCmCJsdKuAKYow
YpoIdSQARfsjHqXnw96Zq8//syZe6hah//zATn8/wWDfu43ED+v9AEiGDeAPyZPo
N760gKaA4pLCaHKEl6ftpkX2oek+R/6AOiJ7saPMDMZWeCc7ZG8i68w8P7tn+yf/
VFzuBbFJoQzI9nwAyUQElvr6UZ0umAvjwLMZY45l0GQ5MRbf5mrsZk0m1gbEu642
QH5HR/ZTfcOOe7dhvLrHx834EKXAf2F+HDZDwZfdnqbqiou7Kxzq61jjGOEUjQmm
e5i3oeSV5E2DjsEDGGGr/PzHTKV/OtpQvo1331+YWbTmKci+dkgPG2EYllv1pTef
KCAa/eWP1ECbWm5Zh8Zww34X2gYtg200OpbIjVlZTyE/ceqDEmM9YDTVvwCkZTMH
VQovnsYQSHY6C3IzGNR1CwgJ5HeAyg+Kc9GUP2AmjiyRFWccgzjJ+M2pLIOKdngq
gufC7xfr03M4Rdek1BRx41rXELUTBGAiWbCAGUdwj/m8nTzP2CqTB+uXF452g581
QHWMVnEi6Q7oj+P0e8symGfhW675d8FksXdX0cO9ZMQxo6uAtVv+hjXXzh+lzlXB
milSSloQDdk7qSFfdr1HepDm/KkZ2hL6h+bTo0JP9IYACj+P+R3Q782ewnxEYyMZ
J1pKIAANR+u/xowheJq1DDHmcaw+yl1oo2a3yHuZsfrXXhOXFWHUoXRgPKgEFZ1i
R4XFxSew1HfQMC7nIPRaJ9zFzb1zjrTLqv+wx/Y54hqMY1njGw1SJX3GbPEOtr78
dNOHKokCj1fCrdFfa2CXm3IVmLQ982T0XXQsjwA11tdCUsSwy8KH8TAB9kVzg8fP
QZnDHrBBsaQmA733xJSnRA4W0LUWiXYONbpoaoNmMz5GyHhM3Pyv4oJ5EWybvtH2
Gr8Zukz8Uwqk8SOrHLJa2ik4Xv7DStXOQypB8mFik20jwhs9nenp03go54Z8lF9G
UZ4/r8Gz+ydY66wia6BG9a5RL0Y6+DkSIuGB73zteKK4sDaUdl+EnED+iHz02nlp
sP/0bKpmoeGvRkaxjqC2bYelEXA2q17oU9vcsbiGl12HeOS9M8vA/8oSg1+02+vX
miy0w1e8BivfbTQU6xoScAk/774Ed70kHR1bwegyKBUYmA0LR+v3+lOCmGAaonT/
GyylSixnqyOze/D6bxoymG41mYju+w5b+O058X6xlW7IWl9NQsElHF8u8RumztrS
HDN5UCLCFlRPoLvQjZfVGO+hORVNjJJRXSeI847mRe3QRPPwFWGU54Nc7epvMdWd
M+Ev1vQMM2UApif+1G5aZQnpV6aLQ2yp1mvXg9+9Ou+w4jlGD81pao0RqwbezEfv
+eDMyiiVttZBH4FjLET7Cq+xzcTnj71VYsmafda1EjBRk5rwkttwXST71vSXU5u1
5fGcKy1GHHQO8CuOP3FbWDyF5eqVUMc7nX3IGrFAaimHrwyuIMUD9xi5kNP/M/n7
Z9THsghsOUffxJxdXf2sfYF8JEwk/d5bHew2mvtYPO/U834SuGrh/8CjxDWhZcwQ
yEjdAt2rZts2iqEgNP2paoOQ5/IstD3Z874Czgw5LJkZJ6fKkpM+w1keZppsjwhx
pJzpY8KWZtoClv6pAjYFyc5LZ26Ew2SNNPc68srig79OlnsrdpgeUZmkegnJ4uKt
6PO3W5+07kmFTGMOtKU01qeAIFKik3EndjSSIeVSA3Z6KM5SRoa2wf0Jd7uXQ+Xz
GW2LK39g23uGOzO41SFY80imr0Mj2MVUp3/bkwq1IMP+N0pFY16kvLhITBUY27+j
5/F0g3lrHhp8RSLqfQNwd1q4/TzGvIEnlC28b5IJEPHUsoiSdJzZtu+vki1WpkZt
r9vxZH8gLF+0DDyyTlHVeaBUspt3slvDjL7gTDsgTCoxrN0sa8ROfT5HQvN7+5QR
Q1dtB+TkVe1JZU9lbpCsi9AhoFiE0A97y0WJ7YDX36DJrd131YNa7dvpmptv4/Gw
ljWhn0sZBMDPUUVKcX7MIpZC3mN5XBINdb0YnfSQF9/Ow9OwVvhsWPGs45X9/vr8
rCDZDwUwUkoUW3lAxDSgF/Wq9+LEErkb3vAPQ77K4wgLrYXcQku07R16GIHVCNbD
S7LA6q3L25oJT7MBxV7yCxNZl7FKZL3CjFlbY8lfqxNX1emn1wOtOHR9ZQjKvanh
A1As8B6BiaZ8hqXi2n0IllvOjRFK8C3rY2+fHoCSuQezscONeOs77jQExE1R+SPG
x+5ZUj/Ckvqxtzq57ATHr2TvBlmPP5SeDS7Dkt4r0D03V7XqOUBuv9ayjv0nlpMQ
+ZJBJ84oUq3LibVZ+7D6Vljx/poKy0oW/WB2kmL7fQixylPT0IV2EQuJUmcBAOeC
RVWAr+gTPnAl/GmB8zL4yBz946/g1+cCJE+NLoRIbZyos0y3ASAIe3gwhyUlv0qd
XYBwMSUKhDvLb5+yn4WfqCSfhfc6CCtlKHyy+R+Bfe8NxtJ/pFOlKW50RmHZkU8r
/iHXsXMHCKmV3WuCDBDHM3LBC20Xsg/DwKTbLd7E5RziME5JRB+lZmoE0a0jHC6M
sxdwU51xZQ0YLI2tfIUEyQqtGGTW5C3p0vFtu6K86YAFtuthjmCZqf9yc8q1dH4Z
RkVbdwluPOe6Jm0C8G3WfR/Zh9vgPMkqplziy/gdAtUNLfm4mSQY0KWkPDkJzh3k
JEKHXULomX7qWakQqMc1mPHrI72paSpoWkvZNXlaCT1ZBB0/eOTGGdM0jJ15XtKe
pNBlEyruNg++ckEZA1lpiM3kSZCCUAgbtZxgy/nDbNlKFIwaOp5UWQ0j2gAN28yN
APgjpJGZLrcAJYWG1QXNCDly2FTDVIGpxWKr+8xUSe76qWufz3nQknNCr5RLqsnC
ULY9s3fafpJF8ktQu23jysiG+YoA4sMY3AVD40czg+kno7bta7msvBxJSjEy7fEh
TyvwdYmeTmtC5vHn+G3507dhKUBzToq19u2nU4QvRUHBrFkfCA2rvohh1zvROM+J
XIpqsCCq6uknlH6tgze193+yun6SY/PKDLDh/EKLIRutvPyr6e6x47M5XO+/O4Ln
bGsvZOnW+zDTbhdYMSPmgckl9ihvOzH3hok9ZNxgFl+KNHQBbBxgLjqh0//+VmMC
waQAC3M2vGiZ4le4T1n/VhJSAGfUBZLliYLk7WOtEKdifgio8D8Zc2K0nwjwD0Fc
FD0gS/LE9Qx2YSfxnbGEpdG3qKrF/6w1re8v7SI408uHcIzauiFrdCiQohuQEqOw
iiPEypcy5XsjzWy3dsjL5MsVfQ9rFEHm79d45M7FLl+Bz6cvyGP82qjYgwvPNlH0
getvcYju8QiOG57HXknT6Db36v98KoIayjW1ElehPhViedbIgoiK77pkbIqoqBuT
n4J5TKMhDkoslARZOlrNgRdRHylUlr9Nt1IRHpGnYpAdSMwEjR358wBxFbqeseD1
fFDJDoPvIXBszofcMlyMPxGH2/Et3f0A/VTqMD/eogKxZ0uWgfqciCTLcsePn7ho
e3qNtHjtEL8IliA2XfeCPNcRXxIqsJrfXp31KR+CS6DefIJVtdQla2Wql2lswfSP
ESAbi0Of7vxiLNq6qmHWQSdU4C5vWA9z8dHlm7Dt7uhrsPVDW+kiakGlKakHEiCZ
RzugyLBbebY0RpQIh3K6Kk4PwNTgGWj1dYE6hTE1LsfemQ7pDJj36tWhoOo2QzQe
of926uaREewjSjL1LnVtG3miVR9h/THikJW0dbAfj8VqmvLLHKJ8vCwSCpsihUrL
psGv5dktGIDCL595rFwKTkwzZTPRPOcbEoYXO/hSKOSaFaTDuqEVoSnN8QuDuMSh
gYrcIpOiXa56V50PGTyRj2e43mgX+8a83dIhLcMFJwRWIiUZCsjPBVolRWEcqyU9
/jCLVlxisSbgfjNuaWXTduP5rja3TOhEK1rDx5lTrPlkEwhUbNUP9Dh7OZvQW4US
KD8RWUXCgWqEpyyZ0STy3FlgYkDaDr3EG53TUy5eUCkzFduXNnxSiRT/AwnFqprZ
0upsw8SDG/9garVGgLmEqXfGBYLIV7u1+LUOaguEx2GzavddGLkT/Em9YOyc5b+2
eqEr4rKGXHuEUzfFyxFxLQaDgBtSwnoFEcRTTkidVmRZ2zKEzg2qnslx0mY92VP3
lu3re0KNYA0XeHmWEBeDWYRej6K3KErxAGDqxGvRxuT8bWRclMkFEvcH4uglQiOi
769ML6Ed4KaY50lk4aThObJtrY3PMTTJyBZWvIlCQ0BfWbVYvrMxx68kSVoRV5vF
giuYRKvhkL3btTZ0zZKsayWPtk0SXfcWCUiH5JV/X/hj3SUjUVHB3wy1avFnVWvD
2kHPnoxPuZLqQ/xYre/7yVA+mBUBjE5BNzpwKRDae1trn8yFPILVIdwr3vBKrgvE
Brr8vfGOi2+Z83douLJT8iJTjLb20uePryJ1fgx6nGly//iuzsbXSGJgpn/5iT8U
2ZEmhKjtUE+M8d1QkU1wyaZZ+V0haPVKHBcNVd4ea962P/5SixMg/hBbCh6W1u9h
xgL5+EYSOwR8Wl2kOZzNMctb3KO8r3woeUJom1R4cLTR5RHpdZQk/f3a9T+H9cXM
IiGbCSpKQuORexwBsKI97E7FH1fjr4HlFWUDl63he1Kk6HFsdlVjPXAx0QGTy5fQ
Fo1laxrnocZc71pwUDNZ3GaXrcujA4Jxn8ATn4BKkx1x1AJ5sXZFt4sRDTZDvAj4
dtSB/1LXRdlzzJfFVEprg0BOBVA0hGtc0/o+we5v15bLvcgu+4MxaA1IB1xl9fk3
5nLvQhDJ5Of3AQ/ZE2vjdLWA4YCY6ICQw4Pshj3IQ10l4xSbgXcC1Lo6OetbSHCI
gSmGKEnAuWe+RgcOp9EQZ3auy8hn6vcHhMdm7HKQSrSBNq6SruTFNyfBcylFcfLK
MZ51k7nEWugBINFV2EgzMD8wh3o53+q7qC+mV1kuHCLLNmsj37LK5D+VXd9Z2GZp
+hrS8IZS1WR2kQcZdQnKcfspABAp6+GEGCqzWq6m3fJc/oREyZYTVdyv5ItDwlZu
jKlLT40bFd1MtZzVSE+aMr3VbRoVt0s5rof9M/rV8MVh4CTqoXJShFlSqSpyi9WZ
50IztmAhfyjn5xwveGj3r00bxFR5DIUC+oIx9WBHmlJnvzcGU6BT8WYxWpWtOW6P
dag0lrU4VHK6R8Fh3GeDqJz3vqU++EGkjoxobbuphDfb0JTWZ284Ote3+WvlHm/s
onNX3pV/qe+zL7ewRTv5uk+FESHsT59nAWvnjRoV9fuzTKYk+5hQviHJwYbzxQtg
70sh1lfUdbOAb9pofzJ2/3MUs4NfKEUC4gQ0syKV0ITNZdkJwbi77kXLv6RSi7Rp
c6Hn4DRsKVuMMBkD9PyWJcUFnrAYCvWDq7rX4JvH6CBouqMR87jeZd6JsrbzVBuB
zHHf4NF/QgWXl4FJuxshH6X2psS9dsDl4FnlGIgzpTyZm3Uji2KlNo9tpeRp54SX
JreYgDvo/dSGG+OLr1F2geCDqM3J4VyL2DuucKaH+p6/RSrRVBXVh2CoHRVXfUyF
NflA8hXfHG4cjbmG/JILpZndQsSpNuTq18OkBa0xG0Vuf2l7sHsU6ryonuhbM7/0
8wbdY5Wagq7yAXdF/QVQZ9vpRDiqlag9kqXSdQyVXQaqxCM8orJGQiV+x/TUH2I5
Djy36FfUcKPuY+qEy9pP1uiYtMZIVTnqg+i8sKWyYvhL4I+lgTmXcXe2CkSd7idO
xxEhaav1nbY/DKp2mNZeFWHEKHFEcT5PBBcygSu1DlIeOUPgjFyBlvDaXbAfu7Eu
EVa9iIn2k9fdR9ctBAFolXDfNbVapb9E955JxxLFsvHEvbZtKEqEJGT5rX/bTnCf
IqLfqDU+a0VsO4QBuQIPjREjGzcQMrtL+S0Zfag7f5EnfkNoayOM9C5lzzn6qPSl
FoaVyDJ40wGP8FVTX04MpptZcc3LAKf0Kuxu+fDIQZK3L00PpGFUpp7zQpF1MUMd
soEtUTg8xOYtUoC5E1hpl3LlcYpONNUjEGqnJUxqlXiem1dhdojK3V+i5Q9AnNxO
B9Z7DWDOHE2tmSOUqcNsHMTtz0Sr4bTRKdOr0JLuRI2cf4rAByacOcjwK3ikYUQC
xOSSlz5xi70b9ATIhxZfO10LaMJc5NTHcxQySuR0+q6Sv73TVW6pJUrvydT2oXpM
9YndmBAsujJWWA8rX0RmbpjhNIdhComiMyFRMQxUHKK1nH6PEVZQeTmXBpk0STHO
1goNNge9ZCPUTJzvcLyoY1sMiTvpb8c/nWNa5WOB7nijhu1OREy8/KHCl9LvXa85
xNW2vEDO7EqOoFMuZTRAKRrndSWyDDdqMdCmBMtTYmKCY9d3pLh/EPJyxeyKEszu
NxWIn39Zh/35rl5iEIHClmZSv6OSZFdDsMvwbG3aMfiNYnKWM3598E0x0cX6Zv+Z
wS2StkgY/X/yt/H1kAl3yGvhNbfTqwXgpoSH1TDATp4be/zraxwv9Hkn4ffdQnnU
6JyuDJErlQeEanjcGouZi2TF3IcAZawXfzIC4NtS/Wb+KX4WpHIr0/smqi0ivoiw
eonoJ5Zyiuxikx7K+YUEmys61T0O3FRdxHxxpTzW/8AxmtPgBLbNs5ZCItTGD1nX
22WT+PvZuA/Uk4E+9zourFYnB5hJERLSwHhPGY+cnQaE2T5IWFUZXIBqZwVLXqpb
r7BL5XE1F9FgI+eEVYMdB19M6dMOl9EcY5QEqLwME29NFnlIJJOhvsx7TODhf/Iv
MwndL7pe9nBAlYLrInd0ZrsbysGS/o++GfgAsLAF0skPRXDr/YWPkhLvV4hNe7j8
NqjqsBQghzHs4W8mrjimJxuye6FNrHJYJHvF+OHwwrcSJTMSxqRGgdXLB3XkuErK
eHxWsA/OJ3Tn387S9F+H/uSl3DlYjdHqgv7b4ThXI58qslh7oDKIEtD+IBHBfP7C
+ktOfJzESYnl3icZfRwp9YYvcUNf5YY9o9BaMg9TOADO9Udb7SDwg3/kLQot37Jd
GQ50Cyi5Vi2C5yImvdMaCY77tC/6ipfLxGs6B+SyUEy/UjQW/WbaDBzjD28a6dE7
P95wZuc81PlFPsoLobGoXwnjsOwPn+H97LLrCmE+x9ynWa0EkmW6va0BmrsJLVzt
7xiX4DBnFXmH7OKzGE3T1/ottbfxCA0QSJUMe4F3gh/1V1RYSpDuWrjWL9IpQuMA
raUB3u+LjdicdG20dPVufiiLq5Nfo6BZg5J+bj8ocyBYyLuunyIfJ8UXhYU7PHsV
MgH2c32CmYnoQZyxYVjYTh4i3aMpIiS4j9cLvt9QmZRxmDK+xJFTOuojqh6hyDta
ZN58R6JPtKqhHaptZz9SidZruwvMnXIujJ2mpVI0VxBLTb1nviOeWgStB7hF7aE+
0UzRYP2aOAsy9MN+g316ZRhVFkZqMA+Hq63dZyeDD9ybq53SgVtEIu9viVLjMeJM
EYoB58RDSGXly6R4kM5gLi0t/sBNg58AO/rfTqqWKnJxMhs4xxuCYTdWQ+sfVrzn
a+MknT+YwctrN25YTsdhcDFz/dzSRbEZvRZVAQmELxPoMYHqmwQ6Jh/lZMGVXxru
oNkUApe0Jxm5+sBDa754RbpWE6JEtZer74H+vcVre5XjqpRoG1hxbLYT+iQtMO9o
CZvyGYSmkKcK6P4ZTLorLUwCqOH0S7odgZeXtaEmANU1Nnkqg+6w1xwuHPbtPRhk
J738tvdW5PvBC5YJ75uTLD2FETgo6LK3GdsqSS3+M2idDs8tpMMfONBov7wW2ltN
oX3hEK79os3zWrVqjYXo4oOAMj77X9gfJUhjqIYOZ5lPdXumlAk4ZZ5stz+tZ4tp
MOEfoBbXcxvjvBGEM5+8F8g/QMxEnqFiKqMRPOcpn0S62OF8ORJ8/hMeJqeXEwkD
ngnJFOju+ZyjdekrvZIVrty6AJuD4CWOq8E6XWrIssXX3cV43xUfQiMukwvIBKn2
ACz9dT/mUAXgO1yj63SniGMndzGpugIGG5F8ia6YEGaGiFQZl5t4iXLrfETaGIWy
CH0Q32SPEMyqhoF7/xX1C2kDjA4a305RSzJAY4+zrk/hGoSsVH2DHvTlbX7ms5M6
wUQWZfdk9yWvDs03k9G8W7v2FecRQ9umcI5FPFhcJ0mBNd3gU45ILzT6RK/CnmtC
9TETVn23/uw+bdwPL0yidYxnY3jDVJaf0/DOYsaqcHISUY3cK529kQdNvRfFhppV
npFewjr9mX3vefYqWsaOvkhbAzSZma9rFrnc+LlLuaaSDkAp5ceOsOZJpZzucVsk
B2xx+R1iqZ3hrAElU03tDO3x0QS9T4Rzset8IZbAERQHCrLeVooaGVtiyhxa09ry
+g2uhBmP0ULKTRPDzhUI4ytA2ddimoSQL+AorPNSbXf2P5v1T6xAPFwBXMFU1Pzy
c49EC87IE4Ns7957h9etKm8fl+63lxYCAFJMbqs1LOYsiifovb9MWdqxLAMh3H6k
Udj9MBe84QgYjtkCtsn+yWDNjXY05szigGkOca722FuJl2PhK6i5eTA8IEWFy/1o
yozt1WgXfufjbTQsGieCcXIflXCo4s/6x+Wz3v7wWGOnNrOvoqzQErQ/0bxf/+XE
nqeItGhC9mFOUzgc80VHnfq9j4gIV6EDviVFBsH2gWntA8AQfguy0wUlXE55FrEg
psDOvAp/eItCXqNY5PukIyZ/PAVOK7arpA3d5uisJmm/P8tXG4//f203liv6w5Cp
wpXiULkRfFqvPmtKICuBnaU4X88yTvvwo8VFGRjSjXhBgskTF56xvHNFMysLxKUc
/gYwETsnGszCH3FqR88AX4xXq3aNNCfdbZxbBicxzHhmDwdxKNFMcFObvuRTCkZk
qvm5t0oYy32ByU5MclCTCFZ1L8pgZXYS1WiSiWsm2UgCqkqxC+etue2aMnjuaB7H
ezYjLqROBFf4cOtYH6exir0AYbycapqZtXQKvk84PhYiUyfwXmfHrv3oIeJAmB+V
JA/epNmphL9y3/dGa/9YesieerKzpyyC0sT5JXJ/GmAwrfnjdv1LsjJUPTlgaSTj
8saFhKOuN75FPq/aezuHJ939/DaqoJ0jSu2aOJgL8/mgJFOyiNrL3rTS8YlCTGAu
B171fycoQKPJK7Qj7UqWml5lllsmzuWCPAPZLoB3UkD0HNbotIDZo+krisgXzCKa
d/8HxXEkJ4lbnzbVVwlm9CTJRQTHd/PuBz+Gvb4HtMeolaYC+EvkR1hwujZqYW7y
HEHd+neWTJ3dnDkyyr9HgyY8m5Kde2WhPP13RV9gq13qh/iImSZ3Qm/QSn3HVnFl
QB0rbQ1CMMB+e4mnWqDphaBUDCKVBICIY7eivu1LEbkTiMbqDepxtTikj0qWxRRU
PNiwVVu5IajU5RZNDEvy9QunBvYwVP65lTc7HG2BZ8WXpmfj9xmyGBO6eggOmJfz
XSVzG+2Ne9A9z3hOlvHRmWN8owGCbrT+HoIB8eMRYOqhcNe8ctGfCN5fI3YifQX9
wkydC+1w4yyeAHI6igzZyay1JSw5LPb4JvmCpaOcJ4jecHHG9C3R5s7I5Yk2VEmb
xu3ODoCmMSuqMl+dM6TkeEQnNnF+X77msggphPT1r9/vd0vyJkh9RAjvOpuCje9G
vznrTAQ2SrP/gQGyhRSQ3A9oXAcfzSqdW3F1UQMFSQmj0+paXBFAQWcXMUfjZvav
8O9Bv6qWDDbpp86Rdo8Oq2VO+8pROZM08Yo0kw3UgISMvG+DViQ/nPNDB87bRSNR
mISM+EjI308FoNCF03mPJLBK0JPXJ/EiqJvQRAZfngwqTLQnBoCBvNvMbdpJiUlh
dkz4pvX5LwYksBUYBJf39LpGcmdzftOK7CH5XjZNrH+MAJ6ZUTX9nFAnAPRAQsoe
IicaBZNoIjO+yAVqGilakec7omzb5iY2y9wUFDgrjC3nF17SvLNgyTKJhr349l59
rOOtUwilWkPANeNTzj/FrmU7VoRBYAhGbp1FECjxk7d9olZEU7hq9BBiowY859Gh
0IoPsxxEHxvLNx1cnBOUoX88c1XWRSLqRO5AktCSNd5WYyS5BH6SAreZSx9hDgB1
9D175HvrXbFkgFY5kOYXwtPoFCnkCcz+QLSJW6yQSzIs+mlOHA9X+Eft/rrIK3Sb
3tmfOCqQ6HFYaH7iC2yINB3P0p3XMs+YmvvEBqaou+odmKqojMT/qQI46xO0cmIv
mhnCrOzZB0qZLQfknFTZYaNDwdAV+vBwB2kVKiMP1QyseBVXwU0dEJ8U7khfB++d
LhKkiRgjHupq1JRPw2XUzTyzM0jQLKIxjJDUBzmtSvTzZcmu05x6gVJJspy+rBst
ntFchV7Dpq0NY8mImvAAPv+49GxgLC61TO6M7ymbr2GDozJBYhyv19AghtGq1+fA
2zQnNPEFc4hv5y2GI26el4bLGomRxLCvcoJ4XLdfeKHc1hANNri4RcSdVn9PV3su
xGPPEoiLQO2bElAZagg89C1KGIKnFNVn2GDWVjTAsx5yCIPtW8KihGsuI1LuwHXq
AtxYvEdyzUW8z0cmNu6fivWyhsLQ6KJUfplkQWJT+/ZWnvURElGfRg5yqIJtwnoZ
RGqvrSbz9lMdLUmklD6eITqz5XrFvhJ/dS4hKYkYbmAIY/VH9c0/94Q7MBiN0CXh
f9fqiBk8hNwI+cmArHcphpKuA0OB2Hr+r9mt6NAUTGvJeRVUYXPof6eNUZ42YzgE
u9YqECT2GJD8GMi+y+0huH+zMm9g7dBwLdT2rn/D14gObbLutnplXu9bFrAe0ZGn
aKZBtO8oj+YgzUwHTtYQpyunjicDynidkfJaV7cGmCF638TAL7AOMyqd83VWPq8i
MIM/YBFNkcd90mgPmVlaiNMbY2lXEJ6RXcuNB46Rk+CLvhgIi9H40/0wflUYosHp
PCN5GG++11HP8IXPeGrEex/1oA7G5LEaDOBeqhYuxzoxbh3RPp8LyskjgzDGqzkA
UAdBh4rzC5QxLxDbQxgvkbOyMDFl9n0zRHQb/ixq9yt8kAk616LT9wSKv99K+kv4
nkrAVcaTT2Fidm4ZEQ9Zem4uYFjagRnPyfXWJMCNt8OLDJR2+3/IaRKcVuEYUFop
KjD6uWMmvlMzV49f4RbrIkk4cozSbP2M3nqkc/QVJaofRk1/f84U1baH15JyRNGC
jksgyYG1zWwAujxFptUcTVYZ3xc9H5tZ1Zk4/+wRwVe2bHMiDyxGWUToq1CVPAyu
JFNiNHc9q8PMlWy/5PyESVrzkGGt9IEfu+yj43GIwXJasHGhDf02INW/TvLyOYWL
XMhcn5f6drRy/zeRVNyNVML3K4T5S1GyCDXox044BX7sweuvNQYdB64knIPC1PpH
4L9o3LEsRjXPd8j8Pipep8mseAdX0r9ew7WIELfGWSmzMMk17VoEOfqPw41mJ0t+
g6ZaUJCUIWaEJzl8IC71ofe10tZp4Eb83PfZwKRUanVaI0YPH3s4YcpA8CCwzvSw
KiQ4wLX7xPqCgea0sYvI2daAbNvQ8MNJ/nhzyPlfHGm5LWIsVLh9wrdbTU1kuIrw
4GUZYpVfE5lyqpr5ye9COMtjpCoODhAS7AQm/NBjdCA7CMZn+Tzn25f5Ac79dpHI
OP6hNus2VmsK5gDavikp7smoP+5CTiyD8h7JcGNacjAcq9tGX2i2zDtsvvn/m18u
vEdiSSft4eelLVfyv43ghUvxlaDc++W70izPW/78UyCWbV9Y1/QBXzzX59/vEIPn
t/RusUhO69fBo++OmI3mu04J+rnCeFWCekxg80nbjZ0W0fxiBHFEIfIvDOrYEoju
I14J3iTJ+gsUA5TgWVTEjOLHbvpOX6GWCzq/mvzM09og8sYroY8I2PP6n1UQlXq5
/vlu1tnPilAbvfvJnmWOmzUZMk0D8edZkBga5ZmkYrSX71YB9Rm0hM+8NEhocubE
AC41jlxMKBsbxTqeyQsvVMzVjtk37rCgw6sy0n93I1whFK+t16L6lwj6l9he43G5
/IzbGrM9UZL1gtaL6ViumXUaNy6ZwI4o3hSKKKJPTDxiU+IeG1EaKcBxXMSts/q/
YCnc5Vn4zKi/MMHB2Ypi35zbvqs9G+9PxT7m7xsL7sALLTzVyznVm42YnH0zX0+G
UkdmTU34FnkV6z17HSJDK73LZ0cxDupBRt/8A11+43SE4skXrTtiYfGRFFCwLggQ
X1ZF2FGkhlOWDtKZhn/RkueG/ROuOQkZNqopWV0/5UVKe1VZkOt9sBuHVpr8/txx
DQq5RnSjr/FTDu8n7ntBV1upk8rxWlvyQKij6tMEwJ3pH6a2wLf2niEPacvA5KUg
cXK/KwyaX0SMkJmwM163XNtaqhPR6MJQTjwe3q+gTbjD3UrfuhEwjsYS4le6nZAE
oED6HAY5Y1RxWEDoCZjaYO1y3R/qcbia963s0M5jDFcI5lIe3pltJz1NGskq+Ps+
OCKOQUWaOgDVrbi811C66Mb57Mvp6yzx35D/dyJg7X7rTdCIYk+lw4uUdmSmev5W
fLCOCSNAEoxZpbJaeAnEzhzDLX4L4NUVeT2WebHqrk9lENg6IUwZuDiud9XVidr5
YCLte0ioFx3qTRgs/5bdzle+CSlTbvUiIzZ17JyAerJN2ZuQ7RoGVtxUlv9N5/cF
2VX6dNpwiEyziZxQIXD74epEgo4utQ56useHrADbzbunw8tmPScXmceGL/nXdQNt
bUynXw2xgbU9uRqSsqSNfGbv0WB4QIHrsvyBdzaZxqF+/hLm/E17y4tIll3ZsesN
n8ot6pUZboCBSdAyxMu/nZ5Pld1XtLAqxd7YyEUFbDSDvImH+r3dGxo2Eod27c8u
7Q3I8a+6OQZIIMXSUvRbdUmwDO3XaMUCk7/d+Z7byHN5toyuEcs9K9+vl5iMAOdJ
bQHMpwlMYFIicmVi8Z56Bw3OIBshLz3FVSj5MF2gx+d0cTZv3bzCKjYIxBUIlw5O
GO+wOCEiTriChuw/moDY78wTjAGUbIgItUa1jGdRhOrEwoc2LnRFsHsWFcw/KxA7
4DWjS8Y2isB3oFGvRkppEzNN6xSBOgH1c92VBzX9A9Tvpm5psKcvNJCLJWXt7HY9
X5NQTyMfptU+l/KbwKybPlzsYEQ3/a41cpTaqgl+QPfjAd77DMJ/RUhKEwtOg3PL
ho08kRHXWpTothqPXS9M99D3FYAGEYXD6DT5q9c6qCbsB3LX0BpUL4Wlj2CNV3g0
Kehw6VehKtVxwH7kc/TF4KtdnAxTlyqqVFXshVzoJuwNot7pLXdQQFn1YYE9xqvI
sK285YBqkdgRXlmJfCdRR0uue1suHtN6aE/vOkiHuoniKdNi1HcfQPKcgEyQiyX8
KR7ryv3YSUczWwgfj3ZAG7x8E2n3xE91vFucocf1kJQX0kcpkiMlse8Rwt9d/xec
Tn0Lkqji4qhQ6P7wXjyXvwH0ec4B18pkgboWkSakBaH73q6oSuHLp7NKGoM/9cRa
4Ez6+aRvjTSHSiYLttXLwsd2HPKrtosdBa24szNdc++lEs46S09mDC43Ab/GjehJ
Za08Btigl3y9Mejk/W24uu9YR7GF+pR/7FoxgVD0DnrlIicmTnWDOQbzyVi1g4AD
zg/fGQPcKMI/GNW849h58+p2/6UseMFtjtroOYmfHht8PF/0dHXwDw149b/gXvzp
UjbU2VYx1LvNqpGdio4X9z2opirDbLpzFQfx/3gAFwXD28rvhwm35+GBc7BxQ+cg
/M4Q3WIlhXk66AUcpDJR/qx6TIb56m9Sb7u4nWIntPduDnMVyDElU3BMwHECtczx
x/dRv73WVllZJmvHtA0By1KMuSrfk3fzCY/BtgCUmhmuRlAlvdih5nO4pm+5lPVt
IJLSbWbyOLZwFJFGLz+1FZZlk9Ly1275VO7SaUUKO0KEjAsMVRlUUieAK88MRstc
l+aFEaLNteAyTC4o++G3kufekCHMF7uYk8GRtmNMKCuW2a248NbHvIFdEotAr//4
XPwBw2hDJ2jw+4rPo7wsVWwycePDx7OCinUvy68SvQQOS8KVIwRorJe1USZtIabj
J8uKySx/p0lZ8QYydYrqaBnpJ9z6wyjaHBXwDJ4Twnv9PavRy+LQC/EjEoAMBFGX
aRrFJA5wj7sdT74uxjWNfihY95+EjEyWv5/ivuXsL3jpxnylfqyCAPKPmHkeAyMM
J/G7rwo/REFl6L3H/fGTmz4SiW5/dulF/h/dS0fZloTx64qUOomiQ2lvRm6oRAVn
EICyp+5mtBaoHuPJ35isJjmf+yBaK3ORQ7Rd4fB6ryJ6j4y5h9VukuDvOIONSbQD
r3o2pLp5WDiu/tcpQQtQbLp6q3dJHsHUeZtzaJ3gnErNgL03M8nWhV2+bzxV8LCS
1dc5ElfSFYnZY8S+CE9AYsbmK0ew5Bjknf7/hCLja71Gn2pKPEOgaa01Um4rcYgy
EazeI14s9AtnJHXFhLeyGbJUT6KJnYii8IdMC4skichPVp7PvDWnuiMmveZOJhtw
/HwdPikaO178nwAYkAqdoNQV6/3Og0XMMG9OVY8/kizl3ivyDTHiVchSMTxr3cGT
x1ZvOVAlZdDt2yXQdaeQ1prQhoFG63d3mGESWKGI582L5Zw+lCKiJYihO4toj6cG
2gxdJ1a/9LP7qsAHavCjAnd97ExUIfCUEYNbQfTQSvDwlFTZpSDHGbQSYBeUpznK
MGGe0rLeEGsj2uYzaRYWcallbjfzFfUUMc9Qmx3SbLR8ioTI6zK3ayV9/iX7+zL3
5Ewk6150ezPs6R2U5CpWhUCl7v2lomnE7xRWFuTY09I5N3elC0zp2KGLSV2IFQ/l
l9eoU8rS5xLPFOjIk+os/YOMDWxoxfjBC7H6Totnaii+uU8WY0vUV2p+98SNpvAa
rSbi+Ld5+vVE+9JYn+eTfQF0iG5E44nxlaX2/oaX+spv32j7PavNBRuwsc4lv1QV
z04KknZAwfWuXnzspSh+Ls06VWBNPOzHzFogzjGxGNyPdG8d9XAqtdeRFq0RT0jx
POzT0yE+ArjNYe80guI/N0sJ3E1A0EI6OSQhpRDuizgg+49M7SIGKE5FNDAoP52v
qKla5f/cm4FuE+qpLwX7PIlHw35oqA8Qa08dZ+niPobdTrqs9UXOaBm7Qq6/DKwo
Dy8k12yyJx0UNpZWK5j3ofqqtzphoKRDzHhvCZ/BIORGcfgZ3nU+LLUxjLRR6vJW
Uc9q2B1Ca/1hKubnL6eSy0Ivra39x11HubTLVY2wwmzqPw0lggm1+7updRMuDn6e
AnlU/zmlJbjADJqryWmuhJ27wcDmIj5UzptZDh4dTS/qd4LH1G2soEvf3AIloFgI
UmhmZxf78iDcLBqNMuoTRuVmZRcujYNySUNOeWA/RFjRAKpFaUR5e9a6fXkIdamX
qVMYFt7Alhk+jwVN692H482N/K++EN0uV6TisKjw5VjaQToHXOeQoOhk8Jdt45N8
BliwjwHpWixGuvaBRYNlm2+C2wGkVRlwBdHWclhTK9GWu0Mbso7ubaxx9ZGI0VNU
nudZIPahT0qPZtRsEU3yU7kTxCQkaFeO17pZl9WvZn84g+3Rb5nSywm7eu70beq6
gN16eVmryCRlU/RZQwiOLAmkzxcZCqI0gGyiN6jBhM+FeTSL2EEog27+OAjUinHK
vqCVgHfR5lisi3jMlzOVnVU89mb5BuFx6NiMLzj7bEhfc3+jovEP4Q5hkbwWFIHO
DqW5SMx1LPy7hJt8bNaAhcTraCwkKbcPXNDrT3RqtFWkEEdU5XC1/L2S/u+2cSNv
LwsFa0ExCEYMo723eHsLSJEvzaCIaj6lUtmhDghHw+BG1NWSK+cNDiYW1kT99QZO
I0cO4a33vIEROGq7H1hmqHorDWBPtSYkg4LBCU9lJI3ZCJqaqRydr8C66giJ4faT
OtF/oXkTMXnGC2vKtkN/dOmrsDXQQ9Z6LFi3oX6/QEvrlW58APdP1FAYY5GGi7wC
TdMf9mjInxxgYATqjRnHvVCF526p0WQVpe97Hyg89Wh4m9g7Jeauzpql8tA+sBru
Uq8wQWyq7yT8QuBtiumCyEpuXpNMNYUN6iEt9UOVjoKrIR+apYyWLAJp7j32HcEW
7h4/48gwnDRowQeSd+2qd39qk6ax0PPSeKp1WKGcyxO9wzAxbKPWe9GKRfA+o4DM
I6wX5qoTMI94P/Ueq+hSzLk+yrAwECSURDbxMMVQGLX9a/2HeIWi0uo5LTY4Te9l
LtJw56Q0rJJ7yIX3AUWPDKAqqiyuGavGobOlGkhzfv9GLGqiyy7ZSsusyv9Y8Ib7
DshbM63aRkn4ah8ijEdm6Xf/jDNWOIOLKGa2ln1gX0+0WIPv1EEwkMc27JMhf5DR
7czUDEdw8dBYd4O14SpwpTceM0ZIXmhiEGIkxL+6P8VNk9P6Ma1DIw7dyipqrJgF
Xgnn5EjXDYDFkt3CSnFTZalrTdnkbEBHcGSuTokdHXsZ1UUN1moS/EQ1tDSVjYEO
xS6cBmUlqnVuwIrm+nwIT+eOzew37o9M+8zkxFeq+nHuzvQAAasmMK07HAlFqeSD
hKICrY7MiPP4LGVRW91u10Tct2ikZGw9b6ntDIGdH3z7pYV/vMzTdVXRaDxLd119
o2aq1fpIS9102EWntWb9SCL1wbgQE6S0Brb+duvmMQKECw4eneeL9eMp8MZIp1DT
YhkI4MSZw2B2EwplhaH5LvAeFkdKVKf3n72KmfjWX6dxKdS5rf9kFqEcvgW6MEbv
2BO2KaKJ5i0jwh7KyG+mFfK0E3LuPdDmmfK40l4rRq5h1i1knxoQR7QDLKJyHRrt
oimvcdHpqE6seDAYEguUJY60L3nGVYN5gNtP/cayXwz1eSVQ7WRKr426tkrrIl1C
jvwxazs3F7V6tyoBDr3QCfMaFchxGF8PoQiadPDXt39KxqVoId+usrkqE/Zhm1t8
LwNY6kttbgKQWuuyREiF1Q87DJp34ZuDvkA+A7dAvM5DqXlBoiIBziW16cqGuj2d
piGoDi1AyM7qV3KrsiLQvc4WnuXl2rx5UR1SoIHwyt2/PkDd8Ww6lwFZmJnCoTKn
3/crXLuFEZSqGhkbR7DT326qfnJk4y4o/qHO/b6iQKUF7wmObQJ38kyakeeX4OHa
nWJ6XnnRF7b/QVlyaiSUB9sgimfvi+3vC+HS2zlVd/qD2xyzPJEFl6VAXRAXX7dV
yBJnZMQzHZfOS5q1vjk5xGDM0WZ52tU7GgMyoK0rbT2uoXZ/WWjKPQ5lONQVK7Lr
aMXT3Dw4gMAwx2ab7pNwHl1IiZ8y54zqEjKHuwUKVF6n5sk1V/mnDHQR5KoPa9o0
0j6mobElzhC1+7gDXqSdbXPu9DNFNjEh4IdXyjFg5/WL35/VKvTe2fHaPX9+NtsS
5jFVXmorbDnt92UCBo4L3kd7MQRrdV+rLAGrLvq7dnrkPY7MyVsAzgnaWrMW53JM
tJBX2k5W2SjXgO1sDvl86HpmEb79AGvCC9CeZ+jG9RTeAhpVTHD/f/KdXvxvz2/1
E77i/Ab69dWmzAhP8pIx8Sf7RNvYhOO2/ufSjk67wTos2L6i1PTyNtNKKFp6yxVb
EjhRf0gWlzqvtGYJDHTUzH2y6v+1ZFkvhUN+riaO31aLPuicLvT1XsrePXJZsCLN
ef/hk842I+gv/cHCXOuPaYwpb688gMVy/vt/HEMrs0SAIWnGYGOZHBzqfkn2U+Xo
O6E3N6Hqqq7kAxx1IJxQF3Yd3G3mL3DfHUsWbR6x6uUHKBL7G/QE/Sk391NbXeZM
VXwfa1ByXeqS1YLWnR/ocsrVRqzymGLilXVIG2tL/ZC106sYjtQzxpcmlbNUe00q
STIf+9cXi3beLouUVhKdxXf38E3tn/Bv8Tu9RAzO0r3qUFbGnRSoC1/aizW+tppT
DcacLfO2lmDqa4hxdgH0MkdPdnhAZiuMj1gIudiC/g3RBSTqZirfkCFGGFkCHFcc
9mRk3X5RqD+lTcyjXG+8Vp+ylhfdv1RCOI7PavGHGWRJRQjhBOsvvSA8nL+RAlRw
ps5h8ZWwFeOUg93/0lcwe3zw2dJ4naRv6YsqmT67Z5jDPJ939+NQ88jZKDDMRnIb
erbmNCWRJMUmdvPVJXxp+Jeg9rT0xQkfyPo9KB4NyJWSahIkNF0qKzZVKSr+oRNk
B60YeR3yvH9hDXB6VwPYljSPsh1hdsrj3ZcgmKZDNhkVlXrhWYf/fK7FHB17uIPr
fIa1I9lpYYyE5on7D80bAGbJjikqbPP6kjz7AjvBwDbqeLsPticuVk+WXLv0jUKn
0WHvRYe1lbWow/4kEbGjLCV2dlEWaBECyEyQBc0wkGpFT83pGtvmznP/qPoAiFnB
YOK4Mqcnh/mJaX9Z4+QW12e7f3+62TuoNq2twc8QGmEnQpoCZ7v2lFMlXjKhPtAW
TYc+ys3wywvlLoZmppRRM9G7A5uAJ28IRUUm63m7UTkTprs9g6Os0d44sWC6F7dJ
K9UpzFhUHzBTcxTi7oZAOtHpXDGrkwSSnstNoT8Nm0/SpPyy6zzzZvJLG4BadsIt
1+MaqLTFXML6ZHWQ4BBuzq247z0gn3laJmgLTlZJ43czeb9HE6yKVrRHuICfIYln
jtsEPgfliZHaR1MjTX5q5JL0F5XdPN4lwZV73ZEsdLboWnB7kQs7S+xtrUi/zoYz
1dyZ6GVkcbJsOxU9Hc77BQo9sgVlmyheqg93wCnkoN3jvtToEtFd+MuR/bjTszau
hGXvefQoodZ7r6LsBCH+uxclg5j01+O02HDJVl+0BtzcVVE2JRXRjMU47uHpPCUf
mNkpvcT78fvOoU0KrNmW949Pkk1jrHwAqdI5PFb/cRvWvWBs9DDpfO+eIgJdBCfO
czoMq9DBDK6K7GZPkloY5XULVk5uHLUe1rLnJMDOXZmxTxrzHclkhOsRrVWIPZn6
siqDQwmAXdKZ5S2haO4xVtmXegiMmLXJvWnqfgRmD1mNEr0+llpDqHRWGS63dzqm
TPQiU2hHWC6XdS6k2PJC0HCac84ljF7+x5nGVJrr66TwNC4x96B1cG0BltuUYgvF
ocbfs2ghuhvz6YAi58k7+cL9D2NhfhL2oT5/cBDzS6XMcUKCDEkF6hBV9pmPr8WY
h4YcLfWNoiVlnJABU/jxssfZux0cOY+Z/S2xtAgBCXr1riIumcsaQYNDQyt9QKhu
6oLGpy1wA+a80bG0w9P4rg3ro+eqhXN25CAjvN29OdaUjByE0r/nBjVN7HIMQGgO
dBQbSB7KKafyWjAez5NTTX873jtCDtdHENBTrpUQRCqTBVry+SwPRMLi3ow9ZGTJ
Dk9EnmuidAjWJu5kBP9vgL+7VieOHOO4Qm/jegX9T63kBQNpoQ09GG7JS0Fds9DQ
YmWJOCEfCMq+xQhS41qgZSo3p78InZB0u/6JUsLCIk76s+O3rND7S4b3pg2NDG2f
eoAx5/ys9Yn3fHoKuFqeO2sVfwLxA+EemXaYH7S7tYdrBcCSycPDLwdXrDOdI1oM
vlCMrmqX9dUkb9G/IuihHv5IownDYkFdggieEugQQOJvRb9cAGXMVdk0WVnmImmA
iRNAcJN9qpoGrnj70BLxFjp7EtZixsyBwvVj60yVPbRlBjhyytnMv+N7ShuheEOi
7TyR8YaiW1B9c685t+QvnHJOhKfvWc8iL3UxIwy6XPKMt1Gh8+aRgVMnFdFd9fRY
JAuVCHinbb0q2YxEy5JHkJr63/qzUSF41K8lu9jM1l09jhZx9oPMig2SCYvvFsGr
sQR23l29oFTpdE3xprXHKthLuPaOGeoA0ay7RZSQYVdpqAHc2pMaLTiLCoZs6oKv
Z9X4dg5yju/q7C+u0tCAG/cuU1roE7uGE35d3KsbZ0NArSgIozRL33gxhpATp6yg
MNU4x1T0n1B7vtxripkm3Bt32O6CyfDcTWUJC2zlecwrl4SfYX8n8boWHNPYTpOn
TVm3VW0ArBUjhfoRpaNjM9czTiTSkGuJtvSnCZZ6oMURdgOEuJCvBHHQT+DjoOZe
h0vFAMg31g0qkHr3UEkTnxN1+Ca+eg2kjmQWTBhICCk7Uw9B3z+cHWU28QOz3Whx
B8wFcQ8ToHIrVfdLD439M57hrRcSGGnGjUniHmFLCU5tXGIhzcrxHCTLrDrifGy8
98QDgsjA3gcLT30g+Av5UWfrIDPPOM8XYdgbRl2H3zlb5RcjCXFV1CCx8hYeJgCS
UHcXZPqw4BqnpWcHeNkW3iuUuRxwq5afonU6ac8jlHCPgIzO1unmuZRr+C4VuTVL
GMpRhNn/xJKoc77cuS+tZpoEuGEsLgJ5SNBVGUnec5PapS0ctDMioSbKqWSaR6l6
EaEnIvtTiDZ6lkhlYBgX2nxg6AurcH/qF3Flvhw6NcJNOCe8aPqDD6Qz8eAvZvA6
FFiWwCF/GGb6QnbIcKQLuFkozRkqkgZLpB6uc3lrxFnNwivoqbQBjgXeg9odQKFA
2G0/VCmoddj9Scm/S8RJtajXSgojvIOEfTfID1hhWn08xDy8uvIFCcIwCCx0WwMQ
GOYqMlv95h8JsxzXPPxnWDXnebV0e5w5aWRwcG81Q5wEWkoKwaIuzK08RNwdaUGc
bfmYe/cHb0m1RPyXIs8Vkz0LPs/6xcq84/MpD7HhcFWcJRtf7KTBFugeuI6/is3P
RtjF2XRnScsHYjKZInjoiC+TlOrnFz2zqaGMQi8WRWvWEgNhVyqRYJ9sDNhNdQ1T
zT+tdkWqvy5A4H2ep7N8eEYhfDfUlO8RzN9lh7linbgXnBADYS63UBYt4a45h/PY
GEzvXv5tsa0EuumKC9Kb1GuJBWSMdYvFeqiXwvJphNzXnJlW6n7bAyhp03RMpafj
xkZ6S0TmI8+nX+424VTPxgWuwPb/LghgRahnmPzwmbSlWEAAB9fwDUClFnwUekkX
AOIPDVoCyAA8sQb7VminON+uaHT+GtcdhlfRLW1LrnFZpz8PXBRFIUpB41jYX2t/
w3wRIWAOphalFZOCiQUjf5Rbq+OSLuS2vZji2BDDJ6cZSmqtho4NwulkrUpOdk6t
0lx8ndK9Odr0EL7fjkmtxLgSMeKUngB5cskWBoJ6haSbJ8+kYR8iRl4RjEXuSRpb
egHLWpkWI/fx7+NJ1RkpQ/aLF8HZJSs7LZHMZZmDiDicgLJ+Y6exXF+Kbr26d6tI
cNBoHCQhsVOhfAqLH2E7q+RfKUhe65gQQTEBYCa8qEJNToyOazDBiG01gvhkqd6U
5MPKHidvYlAtECAOQNLhX2FJh5L9gU5ursIMQxjAZ08+WPqES8uDpMTZKTdwzA0d
ZmWf433uJeTjBV29vaQC4u/X2XWK27/ITODdJ2EBCNgBW3yPKTijwcb2iqTaoLFM
b1/fsXGWyVnh6dG2NK6e49xZfWYAPr8qxnA0YnOzjHfAcrjpA/t4c3YDRqYBoaqO
X6uiiSQ5OX2p8d8QEdP74OvwFIzF9or3wOS6fspNrGIEl0WpeXcavCO8H5gqNbYc
EbFFAIynR7rtt9E3hFJO4bOUNPrl0F3ivmU1u6nndoC19Cfn2lUMzpc79BYBQObe
xwFZoSuNF6AM/IZs5Dd1vsG6Wh0pxP149W3bfHZX/sCzFapXnzFdMv43DfF/T+QI
jCMmmtNM7hHrpRK58GiOBeshea3RjP3S5V2y/B0P8tHMn+7zoOyPA5mQ0bbHNeFB
72S7Ji/qGpm4AKdlNuFInGB4p8g82EvDrBcd/xtLUZl0Qm/vsNOEJZXtsJuUYDOr
kdtsrTeG/+oT9Kpr52J8gtUbCce8+PHA/bBME7MM8Itf386FaEGZVKyj6IbP9zQr
AU/KRZzTNuddBIaYmp1dhLZ7EIJJKlti2XVRlvsxLEaD8Guxq8N4d20k5BkmVGqP
p2GSnAV2gRpFMoY338OMmKS0dIqdmuH+BwEiLYZAUPmsi5QkpGlXxzjAJwTW4sAZ
RlkQr0sOhp6Elc7BcOy39C/XS5eIFbFNeqMW3tGVnpLwFR+Wk8udttxa9RaKLqKp
cTpCTv7EtCnXXCcavV8wT7gqZP3G3AgQWB0cWOK2+7EtZbHN1Ixibf/XuxhUCES2
AmiwWPvpXlAzUY2sDfIQe1PH4/DZgQyXUngh4LOMHQF8uyDBjLMauSo3HzSnyepq
txgU8oVEW3OIpaW/y/+ia4a+nrrwmGmQj4HhPHb1Rn0+V8Tc8Jzwubn96qPmJ17p
dwbdL0kQ5F2IlIw0tCA45KCK82jaMiWpu86NcTFFTwqQNSRbDZAXEdxLl7kpe7EF
nbfq4N+OZXVCX42RFqUrEYSwuSG1b66VcvfhaFH3nKsgMJPVSAQ+3amCZGdv3bwv
gHVHPiYv7BRIajnk/cG6GuerMbtAjchgP2E2Kz7yrI93r8m8TF6DomDbrsFurwAQ
Jb6MEHu6fw2KtCRp11SZUDnaHmK+vGYJK/qieNFS42U8+4TAtL9wN9E8MpDCYQSJ
aX9W3YKa/pC+y1WjKRq1+VQg95GPqWC6rNvaJfcRU/svVsnO9HO6G6QKYKlWzzLm
TDL7CMmPF2EstubI9DKVCq83WIt51ZGAEFasoBXenStIsuvPTbjdElBMVXEFKptG
fz7FdlO4wuDnZzie8weuvCPrGPvfvajpHShldn23Ug28kJIY4j8hJpPjQ3zTcOux
hcOq+S6xO2nQ9VRKxmbwTwm65Nojbu/kK6GqSbjmcXfjHLB8e1ahAVY/6cDD/1al
HwzH5VFKPFMg26qQe4qMtYxvkUirVk+f17+CdE3bgPz4Wmr4Bg3DwFz8r6YpArmc
/9c/URbXvsHNbusvC+9/oayyVtFC16cWVq8aQJ5mBG4xOzgLK1iJ47MClrRa8FoQ
wHhcCVT1+hK5WiSzOkMnEilXUjwIr9RrSVCoSJGV6sG1nHajIG9mGgR5u4OznR+U
KwMty9K6f3F+dG6ojbbsGjoOAxUZpq8TzPhv4GCXguw3byMfIpJExL1C66Pmod1C
gK81/7vk3W4NVd5pG6au3QxXuupeZZGGzY9mo9X+F59Y3To33kwL6k9QVuU9OkU5
X81dLLkgIK+JUECmlWYOSMG53AdDYtivB6J82ac/C5de+jHOuvWclB4KbNnHiQay
qaONOmwdkIjbEzeoj2/cjhg2LKwpBcMXTT8YYs2/lDcRXx+NY1gb7o7kDmdTwKfk
EP4cMjba0VACSAeGLoGGT/4d6hUXndV2Onm89qFHb2V6DMJRpGEsnXxx/3Q45kNV
avWzLDwCnZbnqnGwImgsMuK3LftuaabwU3u27FkrX7GH7eAJq6fUgYOx+6+xwdSV
60e/BV15gjCvgdXWr/xA4LD0lGuUrGDPMHpIHwchs9pBF5dT5IB/k7usGMxnlqHl
yUheY2+IaqkezTLiuaHzyO4QiFUpaGDrQGLNdp+qFX9I6ZWSoJeYIBZynpKziDRk
57GWQwn1/U7/vOW6p4qE/hIWdQWwYis/9lRtmkwWHN1DPWRG+uk0OiC4BAce8tEZ
zSKBVg48Q/pyvV3Aj+i5zicgmsC9eiKHvxmC9kljpX0KmJcbZBYfoZYithK2rtfc
kg2263nL85Fa7V7P5QUtN8YHr8276v8EbLrSzWa74RImhXXaLNtqGFNSsf6Om900
NaAwmkY+dYh2EpndjvRCUERmIm5MyztUJq3jzQUF9KoCqXq4OdjP2Zl9SQ2Onsjv
U3Qr48fA6abxd1OqHZxewmasgGptrGq/k3ee88FMTqNBsr17m2X3f8MjbinG4LMO
3U6kVfDFAQb2nbqrxssTyQZ5zoeRWlS7kwnkg+70kGsI4D5naDJoJHq3RQqjbSZA
tz7PHwXfrnOuWBCRtJ07MDgad3KoWDBkxZG1vDwmGXJfaA5y8ztliB87vvsuv1my
+TZzsgwr6mMxRiDzpyyLEDh37//U80KM7H8ZHjD4OU7wwxGcbKYwz44QzS9gHewD
rWkkTWfFcJraSxqzkjHgMzcEMnf6WNVegJjN10jVAAW7f4wHvAOZklcj/LXy+Vgv
0vv3v4uyEj4X0CmpORuXWb8foWQwx4JZLgIXcikGHx8iKn4OXOqaZtK8v8jH2to3
HopbS+E5uV8YWSbT2OQU4yHxRoFOfe0+5PkcZH7GUijn06HEvGxc3vh/Pw1ZzrzF
Z28GhDraxcj6+d7fyXepoxj1od3RxKVS6Y3JIdA1mujmcacpreNFnByTpUOtLYaH
F4rrT6OkCm89NgN7tOb9sLUtsI7lQwkH8EHrZPhEDbCHbYG0HvjpgqlC3+zP8Yq8
P0umsDBedabMrZ1L+0b3V+vARn3YHqLNm3+2Gbg1kQ8hFL98WZe9gELXCFv2RQpD
pL3NoiS/2UiNtr6/7lRmPCsrnNCCj46Iko0RJnUsAuW70CGZqisuZFWkVVY8UJUH
jW2gkz/QsXsO0ZZ5eJGF2c4HJY2HH90Y8dbLjaW8fP2fppmOs3oI/AGR5p73sptI
hzk+rxtKA56OvDx42vavQAfyYXdOlA3c9Hnpnlm61M5YQ9Ss4sEc3/lW3Whn9FH6
KAc5XRcqFE5Q3rhTGo1OuNoZcmqkPtCDwzR1cBKliDmpgDcBzD/n48pO/AAfEZ18
CDy613b2c3nmPpZlBoMJIL8iCmbe4Qs2wsMEH73uQjJDcZ4YVm8J/QxrXJsVMphv
mjxI/hRA07G5NhdeXmlXMPewB2gscGWT3DFQEA9T/sGBm/u8widGJ37/hO++lxfJ
7mUs13l7A4+5oWpZ1eU5iITMEVDDUp5HS1WBfOcU7lwHf0uEoANpWtJ50d8R/QWr
DT2O+kSehN2VCECNuxXli67zb9sTwUVW604CF11yW2FOjnN5OhxLtZMHTsdJzhrH
JL57j4PgUIXRV5e2JkwPld/OQvAs0n5nujStcPCl4JlumveL359PTnoTWAFJeDgX
5dCCdWZ/zZZS4m+SX2X48FDX4+n9qglWDtK37ZqkNspZ5q1HCKmlPfGN0hEE31Tj
nm/61KMbUM2+idbpfXMSBcAmpz7nO4zxzPIyXbyJwqw1fUHaNb/vRN8jEzZtfJCB
KSkbBfVtRdPJflg81mdefELog9OnGsRg+jotqypjgmDuc8mvpJpAPi50isIpoYTz
lKd50vd8oh+SK7iNxO4Zf58m6g1VP1DlTX8BBGoBW1o5A9Fnyz289tanFkyDeR78
GhHLQeNL9kJuK4CuGAcnUZykpEZjUIFPraGXSmZTMkjGxRZi89HVjV5jLZ7G2lqQ
PGZNpFG91wfIY2fkOEK/B/AwGoJwWzy7CViPhlKFB02drEDFZ2fWOWt3GFufIwqU
2o2cFw3udURbrTcquUtLb4d1soFQSRuYFrKX62qBhP76gszDprsQjibjQOnMP+wt
vHUIBFfoIbTNO4ZIDtf0hY8Pd9Ioi2oWz+pmsZ99UTYlgmckF92rxZoFq8xfouDa
lV10qgL4Zb8sm27wuWZd4fpvuRDmBxaEb0tdI1GhO0VbVAguPzVxv3ZwOLf8XIAC
tSKrZtJowXLimkpejAKtg2HPitcHdOto/yUVulMeR7hcH0pxo1AOUp6RtJWfAZY5
dK18WTIKB6JEMovG0PPDGr65sydbi1U//XNd60WAOKFC+qv8uBZuIL3aROFoCGm0
28W9Qt1HuozY8xRWZBVM9i6vYSpCRsXIEqfY8kOXIaqX32PWqgBAIp7SM9O6+pCF
tM4ho8QVywDf4c/D2odiu0yBepm/4Mo4frQ00CJvkYq0smBFuFbj/U3bGGpPSvjs
87TtXp6DvL/OCZ9wGcfrnSmkPeVxw18XuiBPzPD96khMuapsKv1lbnNxK/eKOvZW
Ol3HyRHPqQ/RDOse/ozbxZk/A0X+xHgJXYARhyC6zrJ+EgcgoOcBwXZCsubangaQ
NnVdFIgqHLrZShMJDTogD/e0fdBSatR078lipT0dCiWppwBV/mjCuM6g/LVZkOKG
99kw/roE3aIFaixRXpuYzNIojo2KSXmj77k/bTEqTU7yX0QjTeC58TB2z1OvMCpP
5eJEkdTHA115nuJLBcro0E0SD2Lr+ti6HdCTzE7qrn46rLrkx2Vxy69W+PwgWjmW
JV++OmVxU7Fw91QzzpcQU8nqVnpp6bbb05So99PkhmJbzMt8Sv5m38f4ARCKHLlV
mYYn+2J1wYGQ24qMQZGeNlp6N5XFGBSl8ibsGKoLUkIkhUKLlz3vdEIzIDeW3S+O
rwiD2pMGyikEH6PxpGxZx0SoDMBQg0xmB6Rq2oe5iJmLjbQoWp2Hl5N8ewpbf+NJ
/sjHgobf1eta4D3SvbF4eejfyY++LscFyTiwkYo5MrMF4CF9R6+bv90adRiDywgz
PM5cT9byt/1H9OYpFjI5nXhwQM/myX1oIBQofY6f43WkhtIrl3UTNE+N90fM0yc8
zpQaZrepgNYPcZ0h6OOOnKV4jkyrR9EdEKfazCQlAswUE4g8ao37vV+ResDi9xJJ
1wE36IA/VZia6nZGtxlpWNM3aWnHk9TMFGdezHy3Dqhph+iySHSYvsK1l78WyUP9
Gp4nkEPRy1LuegUxOpls7r5mIdiIdMUp1ht4spnEoeGBR5JQ/mXpjDUvJK/d8llW
qUDaSNIZXRrDetG0oMS45dx0Vt4Xh/qj+EjyYRSJrN9c3tR5hTyknifa7VUJag47
/5K2nZkQe4BSBdlNbj2zscIh1V4Ve/rSRLAn7fHBw4u8965RCc+dZbeDXaP77MPK
xzTKD0kc5Mo0RE0w93Zy91YTVVDhSFoE8yM62eO8OFHLFk41NRUMCqbPMnsTlJiu
NOlGhW2ymLfAxN++bNbDZyRxakUrxmFr6AkAiiLYHeTBozFrrfT6Yl/JvdrQ94Pm
z2l7hvUrrAQ7DgUukTnC5e8GAOXzBcS2sWkYSx/AxmXmy7Ks6F7cx8/QIZAxy+j5
Fz5ahAfVBrhCTRu01xPq1IConoepkv7uunHsX41uVe6zH6r+4UW/OjHw5cDRpyox
up0eMmwLAFUrPyzckleVTghkZz9y6VXz9AYOdp2fh1TJsCzx/eDkB5DFIDD9xJcW
l9fs/C51Shv7kjgo36Ta7AL8b9iqsecYKey3F7w5TkOyzZ90hjkcsGgjgXEAVUkk
RjodoB1M2APkrnKCTy3tCGQzfYYLzqD9YDeUKxLTKhkWOBDE8FunsYHMQWTn37zh
zf5tXDWXbtUOXSQo96cJCNKu/LX239cYHF3rUqAtARE7F8DMlKVo/41geXqXpsWL
XIwRgganRwaxDbpRAPYp5p3h4C3NlN45ijRkrAG2yWdMjO3WFxY7GDy9Fzp4rUkH
6tLK8E9H2O9mlX87t9vIrRH7/3Tgfqany3p5Ls2Bp14Y4JF63WCe3ONS+HoUj23M
psT5U1nLg/dDwTbmqAwBHNKi5xVX6xPJ3a693GyQWvF4mq7/9oUHzybmKKAFszBy
lYHt6L7WBYH2paH5Y1d1u9ZYPLwnTkSh+q8s+g8dtZDkY8ENdiTEKuLp674vvxoa
yKRkXs/5DHz0mJaInqYlS627DSIxxnAcfnRo0ZXDHLM2oZD+TAA/7q1fqP0btJxJ
dbIPH2otUGR5j0CFFGyW/pOsD3OGGDgimroZ9fIBT2EK3DbEeIdRhDGdtRzlSGAO
lC52HQECsUvaYfR0sS1T4UbJRT+MzFwqOBK1+WSKU9nUXaOEfPYs3FlYUkbabM2D
XMyVNZLdbubTK8kRiYmFKeVuBBn67zBqZdHNuK9HYOr40lqe+uMWLND2Rbf06d/j
LxX9FD7ea/2TKhPhV7+r2maiwnnOzTV/p2q0YG49VIxqCoyXK4eegJSDihSOuF+N
Q4O0qfNYdv+Qwv87qVKChS1EV/thSL+sZK9UhIga2lNhsNEV5OV9IC8h9RUZr197
4Trv0rXv52h8BG2IIFWNFBkh3IX7n6BBJ+LrrQGLSAOTpZDlOdz0OxrJVXmatIPT
5y3J/wF4ZWhYM8+o+Hgg2It8/SHj6otS/PbSpv6cNrMGxdYKksIfne7fY7HrPjf5
90JnszhZ7aIvf0K+GCTO0pR91psEnh4xxLlF+QAN4Gd7LTnGhTheKu6W0jD9wObY
+3OJ6dD2e9WkUgY4tUDeoVsuvo6MFRfcfeyjTIaXXSZMWmJHQYDyZkoZM7DRNZEF
iTsuYS0qmCCe1eLOOvkEZvRqKuquVo+nUCBD0C9AqMLsYEHIN6y4hLzWq0k0XlMz
Q7cicpRyXWsLuv9zNftlghl2stRkhwXvST6VxvvLJvnPG10lZSnnPEzILl+r1kkE
qR8Xj0JWxzjvQriMyrhdICxwbH8d1V/kzX0Ky/kg6bbEh+tJNXMW0EWpD3oGPp26
pVYivfGqewukIWE+NA0p4HHbct0mLnqXq846QW2KJ9YWpVL8Axb3gEE2WJs/pOMs
hDHh8JRZHK9Ao1F9yRJEPKy7D7LRF0cie/x/0RJDz1S9rEWjKLweCmUtD3WWV2pU
bgN9lrkPTEkGhwNGRKBC1ngqxG/GkszWk0SWeASl6Xh9cOAbEGAQM0GLREU2Ur4V
AkY8wuxLDcMY6NVS8BQWgR+261GBT0fccCZ0hBvU5oFmhWX8spUXXXwWMrBmiYmV
R4YCWvr8NMHN26/ed3IXFVx7CV82kymLlOtzpD52RFWahjqFdJJzRdhGOf0H7tyc
vlmwoOtA6ahOQ2kWQTXS3kRGwhmJET/HntN+6YDjh+r3gzk6g28tHv+Zr7sep3B1
orUyS1LOivGtjKtEKcLwJD/EVfbetgGSX5qczyrnMXVFt5Hl7K1G+O8ZH8j6nv8z
joVc8AVLXzMQ+jc6cGFHSVsLo1miFtS7tX7vHLT9uyRNHEDgVQ33Bg160Fvt606v
3jcBHpb2TyxITrWbEXKLgt8R3txrlgs70cCYlFz0g/VoD0u+IZ2NGLjOqUV9hHUv
sq175XxlyK5F9ClXI2PReVMe3j6d9nj45pjXqA0Yr0CT5d4FmKbmNpdU3Bu0AdAy
001aBrV9YfIeoRdH1dYbEvzXzPI5pxtLOLNNVXr4bMeZX/C/zhgw+aKGSfxkBD5N
xOzqNZBhMitST+9qkrtaJ1OjcuVnw/FRolx1QXzBcMMAc9px4a0e6J7C89l+jCon
Ab9Xz6zBB1sHMMFCEfc/LK48DU0INB1BBj/JgB7ZOUDBR6MPlos+8TK+B8wM5RQg
5iM6IuIfzy88J+zQ9HFp8HuUVQlDQu96LYHfOwVkL/WChGTb6LiYNHxv2fYby01q
Nn3LrC5wG9yw/cuVE46zJWHvX4OvQw+UbWoVo0DBfq6/wb0upBT4dXV9g2ZtBdau
R1utUJkJoMU53jf/72Vz9tSrxE4Tr1kby3lScWuVPUI44ITIgmU/obqb66lVV66h
ug40Ov7aQ51uCLDf5Iw6VLxKZkg17tOd1zXbMzBvqXIcOH+FpNShcoeIwFYkkb4i
aBZV8BBkwvEcWmkh9AFnanX2AUd1PmzEhX5Kq1yg59RtGnywD22ktlU/X53BX3Ku
fWnLqZNp/w5Tx3mhs/76mwgkcu8lUe0/lUZ2KhJZJBnKkfs7Hgng8qapgZO/scxt
v5OSUenzDmIhYrEh3OidQCPWFHmwPbg1kBZ5BaV8U5SMEyE0cssoIBzuFcS7QDKq
OnPXfc8A3c/t4CBbKWJOy48Aboor8P0nyG6Lc0j530BIR6mGb6dJdAe58VzBq6Bu
4zvowuiLTnnKkiYmKBAfN2pEkFDW4b/1VpyeQi2ESdetfzU55s9KU0LMrH9NIoq2
ISfl+rNgDi/cEr07XegOKOCWE9MPyctyJU4E+y44MCnW2QeLRPiSykWN8kN+Cej2
du2/SXLZ4hYiA74tJ+89FUJwSzXLifBT7ZZqPtkqwoq3Qdfx6jpgWDMWlRXP42SL
QNuXKyAwacIr/RKrHZtP3DXw5dJy/sokjMpEOcU820mmuKGyuGvV2gCwVgGM9wJA
f+yS484hgl5ozgmhp7X9JUaOA840SxeSRkx8chtwoHuS8RDw2Zl1tjSO8U9PVdYF
6I3nwCLnKWJ7M2g/YMGME8DZduJ7NP6GUyvoinaMJOWlyxELveGkiKg5EMcH+4ab
HYcjVyn+aQK6CEbQFeePNwATbgIi9HupcHxAyRZB0iG91uC4iECW5re0V2Cu4Mti
4uaKxpMFF3kVZ2njqbXBYOR2RfaY09CucXDbhalhIdUo48L1bgpSXtI/5xChDrP7
/KIp3Z1fDTzC6DyVIqoJP7XfGxAiisnei6KciGOiU8546jlqzT9ONPQeM/alQJws
EgyRHrcXyCqPDv7exmwlOKAYUBpnFDM3YMhbY1sP0pzDWMtbIim9s4CLnPaQJXCo
HsE8MZGAimHPs+gKJlB4RJyWYipkhhNDtzKjnLsk/kqBRRhw4GD1ezvsCC9ghtWd
MV5gARnvv8XGe0rmpjtZzYGStz0rdDds8q0FN8h8ugyecuUW7QXZ6jpR/qhZ/GSR
cYqpSiXNlxNzByVLw+TgSKL71tT55b05d0iB7Da4oi17WgRYCfC3pROvgFGcx4mK
gB/0IaTj9WDsHG5xjOqoOjx7jQC+oK/YgajGnLqux4j5419AfEuzhWI37PVY3Rc3
PVKrEE4xdTXG+iIaGDJIJeBsBuUhVhPnEUqfehrZ60ygMEmZsfhV/9NtiPE6U+GG
bOwC2aVy3ZgHMgLJOz6H0BQQbixbtr4+VQu/hYlM2JfDKfSHGNSwsU4p1SZt22Gl
M0+MBL71bVZqOFg5bXDvESCTxLlu4MmTcNX6uzEpVJwQb9Z0XgfAVLJ+efcqYUfg
kOqo22XIH58v/AZV52ApEH0nY7D5HeQSCqsoXTxZrYBrnJsiNYVDGN+yvDtmHytT
dRJRBVkkSpbtTTd0p9GqJERHgmc02THzpkGjT4U+3xGieV4TT+erDHY8j7ZNznMb
XcovzYg89BcTOnA4oAdLkxWrKv++GG040IwtqqVrMpY0oUgmhKBeqSf3iDeXDIZG
RvNdReQXhmr5UeF6FcNIg+0J0I4qmiWNQBhkdmJax/HMHyG0x55xjAtZ55mpeJ3/
ZLiPfA4BIlFwLU8/UyxiovvQ4Hl62qq3QUj0C8QbPoacksogGCp7is4Q1ivSIAfN
hE7D5iiT+wo5OIAghrkiScCSIpaNn1rlxNYvsUvLG8L4JpaqBqXPYOVnRvDu65tn
0YpZ1OmuxkKuVgBOGSVRmXArW0FjOfDcRBMYpXnNJGQ4AEJf2OEfnekyaUgNTNBC
dWTYYu9Se29c6x9xjXSsOR0Nevn8ffqs8EIBeHErdWAfXJw/6GnIg4w4uSru2sAv
Xa3OnZhNF4LQ5h8ZxBiVt0oRl8Z9dBFt/UlHrfMWMquBs7FsLcvhXB4WPfTx8WGV
1PR80g+NIL8fiCY3Vv4/XLNSOCkvJ1K7BYt50goq4WGyIdqyeRdZHqtNsxJg3vvC
cWP/AG1UflL4KeADRDq0lwkDeex5xQ4ER/7W4LuTIKvqyrvlpOj7W06UO9WmZd2N
Qp8Cl3hL1JYQE9yYZEaMzRZHier3zwJtSGNcZutRjtE9hpmGhm+L5wHvfIxJajuT
ewvypHY/7MVrnfHfiygqVX8kWxaReUVRwfocIi/G/VHzNqBRPx1Zyb+bcsvUQ7ov
JGI/7FKbjUHF392nbMLi/qQtXSGFEnFPcKIvED1AdzyC//Xz4UpitiufdJtOYSn9
8fC3LOxz9gfLR/Xy9ynMDJzc0ePfSY3DZpBgnnfV2yaadzEpN/LI9iBBrgkJpriK
HRPWKlKDjwVqsQcZNjv8rZj5vb8NDMNnvTPWYrZBlHqsVrR0jxxX8BySfdPLTnRW
4ROGAVvz3PkakGME369pTL9xetkHXF4fpVt0qCdMZh3cFv/lOW5Qs6CodZU77LP0
BMfQYJgPRsKelynlvCYPR8gv2a1rhnA0iBUBnNWf+ZEtuOitk+8+phYmuv9dtWB1
5VLHYrhYfcygr6gY+8cOvLySAZc0vgkzifG5YeXSMFSv8OkBj1lbZ70CmiXsei3c
MEsUHR0EUJwv2Z1kU3GW/2NvoJN+E5rA85cS6z0/WUfHD2gVHbYYuaxDVoOxPQ+U
OASf8gsWaaERaiOh8+t1usHwfdrmIVG95De54+QawAmE7DnMPeP07y4S2U4LrewO
1aO4bqiwbmmtcfJNS/nFqBAnOZ3DRi5K4XYEjumfB15u3HAGKWa0LKR1UzODOZ8o
eZIww8wcHF7oDD1qkMm/++ZD9HmIXqZZUx4qbUPtls4YwdjKML0BdSN9s1roqGWA
FLqAgw6lxq6e3vAVPncnG2Ln+TSIHbUESG3QTVRbkCyoGk8T6iAsLJL+4NCvdhck
kwzQX2lvvkNLaF/ECL+VhkTP9cYn9oLzdZGeJZ0WdOwAhnTAzgOqcHeLJNG3AyOq
NjYlKMB+W883+WyhBrhoeE/+LK0XnsCyqYKk9Y4mfJCnNs4KZn+Lc/1FCIa2yVH8
ltd2zvcYk0VKAvZNFf3WDAMPT0srUAB09TAoo4bgCLw2vNQd2+bwyW0E3hWtMwvr
sLT7/Re2FxkkG5g+1Shg9sCKfGv/BGHWV6/XjIwLhiU8TAFsUBJaoFqo58b8zgok
o+B699dEMCS7tTdqh+GeH/ka8zB7ObOsfckRN1qCi0gOUSKiSrQ7pPQTTHzJJ8GN
6rfLC2N0NiRxnKLliLiDOBV7/i2oOBDtomy1juvpBzHFx6CJFtbgIIzGK5bY6YNk
+scgJcSvMERSywRkKxyu/zoFmIP2E2cNn3Oo5uNGyo5iJ6DAIh3Sj0J0prO1ym3k
9EFc6YZ8RVrhXEvfRbmHf5gxhSbFlR7VM6AdmnTmgJ7LYNHEu29pe51QDgbJzISJ
LZcsARkYoLI/YsCkn1Xhb5Y+ZticKYQSvgywTxYfYoB78n9Nupp+mKsGnar0ksKw
biJToHHrz0Q4KijUN4nITKP94oYmNfPvG3/CIkISDebauxcLD+jHdr6EnY59FQgA
PYj5oGrLCeNdrjKmWAwlEMCd+isPfatjcksuC+PWFM0Nzu62D0zUd37v9XfoVAVi
77JpbTjrC5iRwM830LVeKO612O5R3eNP2Jfg+eJS/IO4UpmoG5URbXc9CVspT9d7
W7mvLV/xWOEIuIN/O5r3kAVbkJIHyyMmXpo0lB9UR2mMA2KxIE8UHr/v8dClzFYV
yYaQ2jbbiTqI+jQ1dqPRVbkAuPsdwWfGNuIrIh4ydbdkEk2mbXJhFM5bg3Y3PnXJ
KmTOAxB3sFIUosiLjljtARxUM4p7dD8VTg0zwAbBrSjLuKxLL5HyiKVF9a9KcKCc
2lOQa6gkQOT8sFoXJmz6aUkUXzowWZp6bHzcHOYsgWK1b3Cujyy5SzQO19LbTOMH
qhWOjLulCecfSRpCbCghFZdgbLoARMeBZ1qAdQAaCAqrPuFYofAKmAtXAdgNTNqE
mIbHbCXrO3ljUiqGARIpbxGsqXb0OwIQqAtqCkUO+wlQMXJX3hROgTFAjmNQ14S1
QEldFrvU/CU4rjA5iTqZyLrzhIW+GOK4dS0iXOesIzhIz4IXyBURFPL7oEctNNu8
lSQEUHaNE8QjtOcbueEVV9bn/N8TINre2pmQPlPvAe7016805Qz7BcRXQ0RWpeEL
B8CQeCdClc5cVVigEQ8oSmxDEH33nbe6I1Q9bUCjhUGyqit3Eh6YFJBfTTh9VFNi
YYl4jfhesLMI6yqoNCd0rJFb6iIntMNjz28VPL8K6x28adln7GtRjTqH9ip2YVos
FnC7hb7cK+RSFBCnGiqxCjYyA5vbVma5FSYWM8VZ5vK8WlB0H4MwSLq2b+GUkh5R
Pi4FZuc3Bba8Lc0UyrsMPM105fUWTIy+62WRgRDh+SVCM9Kba6CLM3OabzUaVSsN
Z1xB906G7kraADLi0Yr+115I0DSh5oXECjE9XSV1LuAP5AJuMPiCvfLDeEuNYaOM
2fMzFHjVRD3Kyo7bYVtG993JzCFq6X8pMlekvYHRjDWHDCpmds47CkIr797kJv3M
1nbTY9D3EYcNUh63JtdVpYyPxnv4nQEw24SRBHhUGVeNeRnLzcaIo0SInxaKbSct
moc8kUWQkf13mJMC+Wh7dsy9Tor3J+FmfjxG2FIIZoYXliLlJqekmnxtDwjhfzfE
BE7929FxCSGCDTM68cRyVDxrnH0FR/7hCTomCcV0xTKCvv9wIOrEqJ+RcwZ71slA
BrV8dGJCUXpzWDtBwBUvYuAZEdVr0x0M1dfxEYYL0Gs10Up4hTZGOieMTj5lbZXT
fQ9pBgTSI/oUX/lJdxSBTKusgqCMnYF014yGbh8ESYVjMnqKBSuDJTdtH8889gV8
niSKxpzf5wkhCrjZ5PiZC7cSKo+j8Ai4tg7LhSC4vCz0H+x6eudermZ1JPSbF3Xe
6TjI/Bcwo+FOxD963ZymIztNeWZa8I3J52YYlVTMPZxyNQEyPQe2uJey17Fg2kkG
tIgqFyYx57NNKD13SQK4CyQMuBssTk/EJwHaMwEX3KRf02HoXP2kgowoyUJUkNOv
leWNvlKAdShYjG+8f6ekzl2ZZ1MXtxhyahqoiuz0Dt7dcuDETOXRrH7m26Ay1h8p
XTEr2Sifq7vfvwi8njekND8wHxQKd7VQ7A8z2Tf0ArYlJm/sv9if+CSfp6ScNEoj
pBRnyhihvsY/dOCBBQxW8zJIBePPDj54QccM75pAyGNtJRYeH+su7afqX7zbUo++
U5Jf74qr9s5r9+BxP5agoyihk3SKSCiWZn6kATlZtyi0pKnR8LEY/xIX16PuTiFW
nwhhwSJjH6bZbLdhj4+qenduERf7OlYInx42o09O1SI8i4LaWQNlgpr8gng+rqPQ
DLZpiWq8M0cPujHJITxObKttqAJUVPCbBTwj6BRaKVixrfGmg5hwgmK3bZmoZu/E
IR+wivHF1TTExQkLRRfzZG9XciZEBq96H8iNIPdEID2t2ESTIFaZ4hsyzKOe+uwA
kYnioGEOaNlK0y7If4XTVFH3T8eOm11pmnztKSRQ+5x/gtN/HK2+JuJkRrWt7xeO
aDJoYvfuVdalebkAPVngvCm8rwxbPOjWlAEaqjNCc1kGCG1ICosbP9F8mukQU53r
hFzFsO5xe0RrEq8RRHNKIwiipsIaILjpQxRDQk3kiw5URo6I1TOIyuuYs5RsWptk
oEGtjjOj4Ks7waqtnKkJJBB11TA369Yl8rJSiK19ZVinFGc0PLq+Q0iK42RIt2cA
pMUmIC2Ppr1ykqgJnXdQFB7qzsuo+8I35L4fzVqL5G6bAaTKRpBWhUcfTAuqZxR+
IYcBxGUp6d0auaBdI1IoAULgaNG9y5Qz0XOEPjMywPNFwE5vlvq5MnJN+AJjUSSK
b3YwuenTV361WVgBZmYTThC4XsKVeo/Gw52OjKjQJVyDzQVrn2hrt3Nbcia5FA9T
puZxKtitG0xJi3sPW+ssdbPK/PIxvHtmece265df5nbtIrnuYsMzDURNf78qyoRI
Dt8ZzJ6d0sFuM7p5DuQvPs9Ek08AA4v5nERjqiZ1yh+vb1oJwvW7DX0x1OfClrkO
fcLEhwSHooBY6c6n3hMU7DU9Gu7mJ/5IDw3pp1/60oqZRpa4Mj7gMXYg6JY8c20w
jqC6ClB1hj8eQB2pr1x0YE2NIAmZKmx7e7PLDLXh/zzoo7q2X7jli88k9CiSoO5o
Kp0cLTIRonezQLYZgRE4VPjsd2MVl97Qy4pw21Xpu/GvJOw71oBDncv6LHALntTe
FR7vOj87pmW9nxPoufR5demMdPK863fX5Bor5SRSYl4ThVJWLO+SH//cWXWlFXXJ
6UzALuDA4WpdTg7NMCuY6L8cKscsOCVUgSjc7kWAJCn2V2k8kmqUXL0qXbh+tACw
a9v5a5ZEFTtaLKtnvAzb64pnpIPM44NqXmbGJskawcrmGBew32lknxw5ystE3ukf
HRqs4KRteXZrMhlfX7W5ceFY0grcdHIFrj9ZwEvMTmP2Dl07/990Q2z/k3AiW2P9
rQWuZMTTKgAaddwzRfCp+wOLRDgV5saxgOmwKteGrvyVF8HwPDuzI3KHiSPydXc+
vulLwVOaGISowz+GxvqyIWMO+vikhSKPb2+kolLLzfh61pbdQG94QesWgQzbLXJT
Ooct7LrBsls1ip1WPndFFLTwWuWQqlUzO6Z50XVVdOPt3NmPN9bOBj79f1JRBKil
KJmwZ2zAhUckdW747SM2pPP9nkNuKmDMVrtBp3pMj7jWYv5wmYQKdGEJWcPlA0wg
+P/ErlvH4RxbL5nRp+WVtKQkD4XlJNHgeZPpRuDfiJm1BIIIzriqfMD7R66srqzl
VMp17j255iDC6GmT4IUU2U+pIQnyBRVJywZ7g0B8QrEdx7PGuFw0n4gqoQI8Zvpm
v6F4eS3qlt/NAsuwIBff3dxAkdGsAW+3ZnQOtVlJmsc5voilAA7U9JUWfkc5sB5R
JuCZHD5SPWrYhCDsUGCB3gJ8gxupsa3tafKChL4Q8+YPvoH0d7P+mytk2LYcfZDy
D4NUibPSK8nguNkPyG7/TKSDoNo2P7CzIkNRPwdzaHFkg6AzbUP9UEtsr+a6Lo/X
fWmWp+VrjxtzBhkNw6FqKrjkE9KBzs7Zh3cb+ldsaXk3TBmfcsCT+E6f7QRmuj/B
47t4B2zxBE+UA3+niMf/IyYWjwiV8KoqZtw7Uo463jHe9normnd2in0CJ81B9Vu/
VVs+eDlT44YEfJeWgY+W+iPImwlx5L9LxGVAVbPiY7EK1vAjIJ97todJCUpakXKN
OUaObXWCa6IeQbjz1nzjzanEXgBg3aHB4R8HRBgYrkWT9CFFrFpt7hZMkq62Tn22
xcBC2aPy08bMGpHDlzLkI0x+elyt59/ht+McLwn2xScOFdxy/ya8lwdBUv6t9AIp
XmfHRmnplBrSNDCz1x+rhQfIInHm3oM81qHljPE3R+fp59qamXty8SJEjdyuLJLy
jZ5RfuoLbymTRbFaDiJFDYMEOhlngMceSwekhQuApOQW2kyttJ+BVM06JJ+xMSf4
JPIFbw8m2fPQRfnayQFyq2+B5XffaHwjimXHnRYOrwz+Ng1sBP0bS/cIeZIms0Eg
egyQ6/12vQui0FoBf923TnTooHSGbjL26zW6bk9Je1Nv9yJblhYwLvLmsY/HisPQ
nHelIhYg7+/nHEhvHf95bbRijox9BtQoZiT/8jUelkoxIOreyaxnJ7Pb+PoYMnHM
bdXQ0CcXZzx8dQwprjR1VZEP3R9vI66hsyaIS4Vifro3zCCBj2m0EvQjdanIOf32
p2M4Lk9QBdGPB7AtrKylGfjMeSGP5e9UpfsS9ZB4KfLO+/BhAzhb1dcK5PUEe7An
465RBb68ZmLpqL71G6Fumck1GKXdmgxFwWbOHiDEBFxxQIynyDAjT8myLAmPVD4N
5v0NFQNyAyDYEWEbHUOAoyhXDzQYOHK4F/uxSY/RQbA8Fm/QIc+WnArhIazV8VGk
dcKUZygBU3hiIRVLpmgup2LuyswWL6xh3SdWE4NLGuV0QchKYrBFs9pDI/IsQDpS
CMBwJUhSGfIpVwrHh/j93YIcIOq7GDyx6Eb01VANxz3XZI1J568RfgD0eGRi+Ewf
r9T/Fddt4xeIn3SCf0cHhPQwnFtBq6ruSvcoEuoS3ihiXeTqm+W1Tn497ayU4XfS
uPX+JRXtKvOizifARQNy3l2qCU01gH79eT5gsUW6krazNXm3LLl5dfDEmxlGZQ5E
vqIMbCGypKSrOL+3Ws8lZo2vEGS8ICqjFDIgglLizfRD7jM8zHyu8O/g/VAizCjm
DFjJSW7SvtMf4KWPHQBNEeG49Ulv+dN8YU6VaSd9d787HwySO7yuexCn2YRDkLLw
7g5gjdv8PrBSTlxcttKHGBUpImLr0dmseHp+K9f5McayD9MVDeKnMyWqLnMouYJC
RR9kI8z51TgnP4/2JehR2zMU96x3TlDqNJdyoMKvEacjZU9XXZEsDWyecXr++Wd7
UBv9B/1ETJwZmvo9oIat7QADVPew/B1VCZXcyrDQ5EWev/x2J9Vdm4+6Nmim4yZU
KewCL+lW3I8dKEwiKgS5D9FDZipK8YDyoiHdUEWqXbZKeIwW9zH7bqhAmFznQQzL
O0dFn5ttFOnbMsvnJFT6zPwSLvpyGUWL3mSTr0iM/SYPLKJB82EvH37xzuK3/H62
S35uYV9zhAnwcflzeYflGw8Obqsxe9m8yifbOZPHTFchjm5eavez6Nb0XNUYxuMT
qPa34x/Jk9UDhLzp+6goW7NvXatVqQlkdDxL/cyD8xP2TV1jlTQZa28zHEz8Kko4
wLuSBHgl5y0gXu7gtnYIOcLMH9Ys/49GK9IN4MVTjiJ0JaoaJKl2VEbZ/KkwqUB2
0ocH17M/1c6OnZ3bb+M1aqoT6vakS9dt2MPZ1tx5ZKyRY+nZXSKYoJmgoHJq80kD
DH6ZRF4vIInl1JA2haKO9BxL81bt3M0CWnyEqWjGS1+Azxwl1XonCkRLC/vaBc2V
G71n/bdIMJ5Z1dQVHduffTmUnl5NpJNvludif3z191Tw219RJjHJl5myk/i64iRB
EOXYy0uKhGpRVspvw1KBnEW0t0d7mWN7i37ECC31Q7tJBLgFoKq3l1KcCmRwDaaj
jWo5BRYtXUouIgKO+WFQTwds+JwA2FdbARrJjGFSO08OVcNoEOBgLggDA3RF95GQ
3xXtIX69GS1MCn9dreBaaBKaFeYfksBpxBsy2DxMUFgnl0EO7W++mjqb/TWy6UKQ
HmcKOVKc4tnv2gnuunywSISaaX2+5TOES9NZ8uG4WhpmCBMnOs09IKLdWqfwzvr1
mpmU56G7sKsmPLCMJgP1hKmJEV11/b7S+4gipsv0BvukVPuVSJYJ5gfcGTVrqVo5
emZkjfu7R1fvFYXhfaHTkUVbLugXY/bHOvtUHlYJbNATJ3TELFucxnk3RmP4YxO7
CyvQQejLesmOVDDa/seVGUKITKu2qVMEP9NaVuZ8+SBkV5XkxhEkm53vmSAMG1y0
xJuOaMM5Dsl6vNHhWLFHT2UkTyGLYwKM6ad0Lf4PcNezUXpWZ0rEqVN/E9tnI/Ed
AOufPhX39/mo1xo1khm35T3dtIzje9nLdZvPOaXsDvefugmYlH+E1atOlqZlR7K3
n9WGiRlGBwMRBw34smcjhd7Yhh3FCW7zTvLpzH88j94qrDNvSFIFWpxq6UmIqjQ7
v+m9ks5jtB841tfrY5M9eGs0mGW7OhUAsyaa7CmfHbDcTY/oCaAle4RYFbJH4zrp
BAYu02e8kG6HptEDL5G56B3UPqldf8REPZ5nD+/NF4+u+0IWRnlLljzIil69oOU+
saXvc/ZMziChHH6QvUaMtRhpctR11uwa76/GmziGCNfIVYz2QpdiyrKgBfkLOenS
nFGy8TxZL9UmaQ4RovpLG38/UziSsn2DkUVsqWtLcSt0XNMVPIewF+YJ1rUVFaBR
sUVeXtnBvbRY+TjwnhQiwel6v4tg+6L/DGCYXGBKr0IJmxNXgCETMl3G+Z8M7NG6
ZHvKAzXkV9dNBx27Ul6QgqwyKSEnkcakPgnHZ/0QPLOaviVchDgmR7q5VNyl4x4X
CpXPEGJrwdnzhjtfnNOWDiOeXJZx7qTXOeoNF87PGOlLOYQNDl+0BgaZi8W71A/d
gHi8nZXmFvlPUzfKHIuSgJdX3qSruIEVYpSYwO67nmPMuTse5HCWuPgSdwrtgg/u
V8SnvXX/O3SsCGfbZIut5pWbLOqsiQxMNlkLTScKtLL9tg+zNhUlTcoNruOyltGi
dJMyesJnDuJuSQ6arg93RCfanHxn5l+uvKMrRRJ6j5PCs5E8GlSmAyYhs3dd0SoG
n+xPZsD85zPCfKXpZe3yLR6XwMCd7K5ho2F4b1pkE09aml426YdLgrRW2WnFDSn+
0kLcmjz/Ugj52ZqgM2QSmz0eRfxARrpgeSqVWiRNyJUii+mg7AFeDzlOqVRTO/qI
dkeju9vvm8sJN7v++TnfEpaUL/tqY/qr95wiJYLrtOFD5tu+qVQXQwRGYCkuKGrp
ACMJOaPo1+TFPFSut+Xsn02sRoSdII/VDN7HRpuleqMcM66JyUyGUd2zgjZ6V8Jy
23QXKOxno116iik9GXTY7dla4FPrW2fcZQlWmtMtGNesXmk4EZgXhip4RlIyRZWw
/lKpxc8LAoq6zx9Gpe9D6sCzPuohmj44Gw1ep9utDa0ZcQKawZuP57kAFl3oXMaA
jGxQQ2Zpqpmu+olAlgW+5XVpWbjqHMNvGMhoWAVDFeF+El0sJ2RTrWNISW89YmtN
TfuPYEPZhUbv4FuuOk/hu8wdaxCQeqTNKHwo4jQThGdh7DNQz/wwQ5WhZ+A7vFur
t9Y6QQXOcPxUcy5szSdpbPbMzUvTlwLbiRtZ3KmrCNCpOczL4how2vbIyW6x3A8A
TNaPJNRgv6zWpn7SoSzZYJU6S3bCK4+cAB+o5QBszAEaGzpi+mWPlPNYcgvqtguM
ZKjfwtyouvBChEn5EwuFZb34dMf9r7YbcRKGcEr82J1fHjXJHknqf9+Y/eogti0J
2FXf8U+MTKMEuzB7c7bzlZ/TIl0Fj9LOIup59kIO9VBcKAtza/Co4urnF39gpe8J
mmqqy7Fp2ieJLHfHrr93vEzTZWaTuvxlaA+U0DHb3ImdFFnNONJpgdYuht1sqGTT
sY/1HdTlDG7+3VN/WzROyqrT/sY0fEGDJIWIQACdZePPCDswnKYjPgOwCbCB+DD9
WyI/GQ2bkjBry/f7qrj6EuCahHBtiZwB4dTRPqhL8q7nSiH7ex+inM959Kjz3qC5
I469xbO6nSFl2ZWwJ9SYLg9oxfX9cg7lBo7OWPlqUa+vZgKeJAdSyfqKZY/8SoCh
phDCQ4dLojuk+xCrJ6XxwszCAP6kfJMOtxk8PyQ8FHuJmUoXlfM2kTJU347aX65C
G2bzPR8lkPMJGPIazzAaTtyWbi039vtW2kLIjRhPhqzKHbFUFdYNi1Xnm4OR9L7Y
Tv28yx1wG5lYsSHHNrB4rU3q8Dm3dpnGZk3w11S/Jt5/iG0tIZ52hMBEXcYn95EE
5bUIs7B/wk533aEpG1MaxEM9sd1WH/A166D4D+wAgthdciZPta90yc2Cz2+oW6Ah
PQDzopkAl7qVbpOR/9tsCZ3h2AD5kEg/hvJQ6OAE5RehKgs+R8HlvTfnL99MUbe+
/8tiddTgzKBhhRGqJaE1eZccFcYrJJF0ZQ36ESb21d7tg/buyUxPJzi2qFpcKsal
R7/g0xqNktyn8MTLvpVDY6TUbIJJ0T4tz4j9Z03tdacDbk+m76HLQguSctAo7j5V
8K6TLEUqoKDuCyi1Hrc+nFP3qlbyplLcGfWsnS/jZxmLdmi5yay6Ov71or8fM41N
F7DjF+MA7Tt7nuMpdo3ai3M2Z3hPBAvu+XUyYWp4Fn8QLltiecLrZrvYsILF2Sv/
bg9VgY0wV8nJFHXYL2toWz9sxOLoorYKmrdbjLjdrzzquhaVjgQoOKdKAKVOO367
I05WCqRulVjkR2eCyl26XTB5PukFij3hzcbxIIHzq/Cm4yX8evGSh2geoTe+S4xn
9EntGs3PrGZnhCoowZUWBORXFZDZdYyVzIPCf2Jr2Lb9DZE5HwohB2wP+8KKHlUr
dDXCEyahKqHSmpxqPE5/05fNNtJTSTLLwIr5Rt4h7w98NWjFY7e7NXth6L+IeL1D
fz4x4PYvR9INKrQB2GF7IFRSWQIYCnILVD48Uoq68InTsu5AURTSPlo5o7iweVuq
FFYHT0MwufKbw7kLic64Rvd4GoSnd4bATbr02qxaXZAR4956aHhkuxOKCQL0mrvC
rMMOVEWR6D6WukpLYP+eUixVdFWbRVQS9MSTg6ppBvYTOKlpHiUzeQAMzGYdjAE5
tRx1wIsFgNj3gQvChrAR95eWbJev5Ri+EPNrnqSe+jfMXiQeACvhZHn5dU6yz/I7
V1GSP7alhmRWRp13XKzT7+lGNbHGNLBj3Kud34WLCl+bmU1bdPSlIqdd/e4EsOxu
1VHw4p50PSDKRo/zzMhxofpoHup/hQR6W9c7TxMqPNXX2QT3tAP9pqd5x+JjM2RA
0R8pEYutWYa3PCyliRIm7VspqMp4hSt9VrqR21MxFiaMYIOiDKYDdmSun0Vo93o5
D9S8pLI5ejIQTk/YR5YfS3UX4Xh8sRf4QD/ASKAs2ujfxksahTGiAtOdC9VUikaW
sB1omg4J//l6PC1wupIE96+QsTsxofqslGELHPV3vHKiIOU/i4CLW+e5kOcz+suk
eIHvMgfAvdf0yNItiXve2MyMvTNlQUHt6HEQLaa1UaUJ/oxlcLAOeHSamOGT1gRP
U+NaoQOIVe1l3EwC2Htks2nZ4/M76hJV2nnwAgGTlMDBewA2I6hLzO5HzngaIVmK
OFVHr1qVIanyQlHNut5zO1r1v2NY/gT9vUat52N6LxkytsE1CutR6F6yXKqJTrJY
2z0Krym2RXlg5ilN1k73RbCPFQbnDfNzLmdIDZeogaoNWjim2Jji9eD9uZDOETeM
zKG5eWz6CRKjcin4BkYexnY+8FAifuxTIqwZXY8nF8hswB+yGbxJ4jTw0qqr9B4u
stSmXg2Fg1E9Ggmkc+ZgoNfPHJkGjBLkw6OM26svBguEhIJvAuihfrziAhrOWRNo
2Xr7Ec7chwU6jNKXhemAp2Nszn2wC/JdBcXVpBLDjDc6Ela4sEbmD7OJdvDYUojZ
ooaZ9paWBKjvnKjO0+Gw5dc3aDvg0DvkfRSHaifmUvkHVOTqVUSSHZjJ057PrzwY
J26UUXw2psd8Ah9g8zwMK7KA0oseMR80kf2kQoPJtfUxrA9SDrHjIJ9ZVWiW5bdj
5BgAd4bma9qa43XUTXB9TcP+GktX3TJgv84ey/a4fcLF9zjVtUKj2tC8Iuw+IOka
vFT8VkDASGX1T7BJVy8aaA9aLCC7weoToHBlo3nF6/zJJ9h1CEsmxfkyHjIfJD+8
eZlu52cedKGDeXazQ6QcBS5OMLYCZ3ggUw1jvAypPYMstJKzBQEyzbHsyZqVehwW
si+tY9m6hEBpAxSSKsVMrdw8nJEAimFeGcpEfA7WkYT/3+1+I+AzqaoqzMO3dpxo
fZy9PvU1ZLyK/mOrWKjOSw6P2XbVa2TMe3nNtg29rARR2d4wW0HN20DcsiS3AvLp
Fb2R7oQ5uAn6XD+LEgfiTxLfvZswKMpEUAAsfypIWH3ZdtYOIkjSxjZq8slUpj1n
RYKxvUAHCni4q0xK2zUYJlFwTL1XvG58CA+E0ozCJrSCKo/zm4LhtSZOfyktPV1h
604WtCDea+MdmwaVjb2G/pmpSCgTbq/JvhERVg0LLT5M2OJhGLh78TekqDLRR1rA
IT2QmW8gzojdDsOnYjJzYlCezygCVH20XydpcCubWJQ4NSs3Argj1hZLUdf5qDCl
HNsMoNaK7GFkWwmZjDPtNsc3ZXWaQ0koAAuyGo3ewchlAWcUs11TSrIFTyhycgLn
YrOTSNzhQ0HDM4s5HzVUtPwovthle+IsLyBPeNYMSxptyMFnzwnu1EsgQSScjETM
6yufO/5FiuTr0r7fijK8ObPzhux54r02cPbmgj9zaq1jBx4EVOPTqxomDKIqoA79
PM+fC44c/s2YsOEmt9C62fSOGH1j7xLCSy6e9zDOWjlcgHkkMxlybts0L6KbF312
Kq4rlB/9a9fOy0S5Z8mo1axUT4aRJq444zFG4jMk/CqFahpkCHjr+UFv8exyc8cA
zqlA5eBJQlwL2CKfS78ggaDvjZ/wB9PrsknMJ45n5Tk+2i3PTcO9/3Sk6UtGEMc9
dlcUKVifgB+LjSU8Zh5JIfefUhOcJQms8b5MrQBQpA9NBTvKSjyfwe+sb+Ddmqin
1MvkfIxWIhwE+92o/wsGdtI1FG2cz9IgqNs7I0JxJX9pWQt2FjwSNLEX/rFPYejE
GlzJgYuw0rKXCzybuyU/yu/gM6VIKmUZq+2SNDZKthZ8WNpnIcfyI7HsmEEpeNoz
DtN25130Tr24422AVXqUuNBF5j8WY1ojHOMw/VHV6IxXoicWwrX9qIHtojCZR1CY
ktI1hoWzF52NJQJmkPz3Bt+9IjjQdyiFtDLc4BE6aqjzwgoZSjcNF2Uft1g4EGVU
//xXGUBu1ddPpSfLmUmnbeAUcPqvWiL+X6OBIAiLkXrHRacvqP8wUoMNLSo4kjdI
coGC7K93GRXUVjEcaw6ISl/hU1DgvksEoQIqLA/Gnnld3Bh/G7hRRQ5L4AOu+aCv
KrMRbiqC/k/X8qXANvLc+HQ+02z6QSzIzczs1Qs9y0mFRelihtLZwNNI0O8CZN7+
0n3XM/S9I1cTtMjLQWNYWl4m++Q+uZq8e++O2IXK+E+iE72F+bgS1/iVm9GM/3bg
VF6hb6OzjOASPWG2iWjOsTBwvMItZw3I1a5rhh1uyJdc32gkSvp2ReHuXqG+0loe
9CZu4jLfYwGWZc3x4AWQtN6PeGKF+HSOs8TReurw5L8OwfUy1zO9IEYhYG0N8LOg
30DCo8gaXpAwmLwU0NJaOJAFrhUKtXqmJhP8qQfxmuWypNYcyTj0w4gkGg891XbD
lUA59twmfNRuJFSBvYDBu8Rmk0/e4ILCOqsXGDW5DyLpNTQsbAr0zmjciR1Ttl9s
bEODH83KMjMxoAa9saMlSkHkE4KEaMhcYo5IKiPP7+IVTiDgmAhF1lo/QL8AYX0S
5IIveuzaKIL4FZAiEo7dgal3sxj/TGJHCqTS7ynvGoPu8RuP253mC9KoocFwMwlC
DA/+6zxScNj9nJ8B0T8TgPOLiBSbcteDxntbAz9ObzTuBXARLspiJ7s7iaqitucE
B/Izu0Ny1z7Cg5iCR+qcdNc2HxTjD1P+xa/wwrwPKUWy/3sbWAg5Aru6OJwf/Zuh
uFXsTkyhhiszxWZ+7P+PG+3WAk3o4IolBzVUHb+l16r6lqnZsTr/cc9jtZOKq0yo
JcjDSoq5rRb1FsuEklMDXQmbU63NNzes/660bqu9FVaJpLrzbHYdeQ51JH2ABBc2
j9vPB/L4bB6xRABVZTpirmFHG2XKKBf8x+exaa4RR3wZQ2Y7iGB/G2+GRqgERRd9
rvsGh6lBiBDAhk0jOwzzrOs5TnMEbyRbaVuEe9GQA72Ky8PaQI/zwfe2NO8WWv+k
dGpYoJ4TEYGkmdO6c51f9Me11Ch+r1Jx4A7X2s/aFny6XHZekQAGG4F06ntirEis
Jr0jXXFLwhMg50OFdAZtNdE1nnhQJZ5/EvIaRx17p2SEh5lgMkw6ySTjrUVpK9dX
HxNSWikjB8DvNDywoBTwCVgS58+boEzIuGM6n5cSZLRgohhrsadFGeAwm8LDs8EG
d8zynsKukTBMn6gWJ90ooMhWVWijfibJkLgLo/AqNcnClKEVkwrMuh66y5chyK//
9qvsEIx+l5kgx1W+ykXcfCt/GNmVo9J5qopP8oeaosQNUwiSUs3vSKnf5zOsiNeg
BlkfY9v/mxU9/cKTCjvadpywKBQMV6k55grEg0Tq9+A7ENPl86E80c9p7ds3YoGK
8Dav9qXVuSYSSvJG5XpgSjwImAu5Ow9CC+dYCmdaYKU2Y926ikoT4ALRRxld2utO
fS4u5U7XUKH2JGeCJegQunmc6qWhe5XcbZQ22Vg3JC8vumIEqorEgnGZnHhnspDj
7b6YLan6OxYnYjuxw5gPbeDDrDtFQvhakSX/CP/6RMEzVjIV5jLLCr8nj33B33aD
hs5Jw3CgSl4rPHsCSUWLOMEcGtTNrkjRf3kptmAQm3MsEC8KRHsCqFSdoWiS3snh
yR5DBrb0bD++Xbr33b1VB/CEARN7EEvEhYQ0RojUOKfvBRoxWAOc/JCBXB4lOMRG
8TcXC1cOkJeWfm3aqkG/JLUM7DXAP1Gz7HIOD9N3XSAcb4oSLP4iPhgR9lDA0Y4S
1zmxzeSgoypFceXXvuxh5J5RlyW9YFr2+T6WLHavoKrjEcGr+yHp94am54Jj3Zh3
PZ8KMABaCW+S8vD9OuV+qx019H+UPBOC94oNrbyzO+XOUePbQzkhLfQp9BdSho9/
0gKgw73wlw+DyTFzobb5yzUCW91ExMzQm+jHyMlUIvFv84Ln1zCGSWOj+YMY/fbE
zP4+bXsycm2u5CbYfGLGriy1NhZeTGUw985UZOp5bT27pXh62ixiTXr7gYwFPFDE
mkVnZNJ6y8ue9oEGkoeX4A1myyfBSGNBue/5IJE9XvMqKnSEyN8XpnINFLjNb17W
eZ473+ZdtniomfEODBKCgY+jNd8VGTGKX/HXS8HI1xN3qcObVZ1odrTMIAHOG18+
Eyk5mvvgYfOwvFQWf0zcW3AwL2xDsIWliZC5bdAJZuwxUhd5qfzxkLH/41RWaYRd
Jd2uByvbNLdIMs19dzRE5/gt3qlGz4JDKaX6EhUZhBzLU8ISpui+WV9chhYmIIB2
14CjXkXjRGwRyEyl1tR8XsgvGuP/LXGc4du8kGRp9hGxPnuzYpeQm0LHN7gnh0yy
WbuvYW36XxzeXnmqvH+BEH0XtmtIHP3TJp7BqQS7jdwbkzEZSJ7woUVZgFscQIGv
K1/GDzu9jkUUu30PMgAdzknUukxjaRV3shdYCpkknN5B31eNEobedHL2MQdAfjT2
pt/J7kKYiI6l6sNDjKMzc+CbwGad9c7b4lwOXvEmiQNX+h+pP99w3oI058AFdc26
6I4Y2qlHaLXkxBCNCvC+3HpI2rYQKE8nLZqD2cK6tPdbTVNTWBW7u92saODSOis5
rsaRqKOkuck3vbpdf2Rp56I9KXbo1gV/absTOUsC0vnfqAIlzoXX4AaIEIXH11Kz
cy2nF0V1g4pclnd5l6u0PVHXICFbvUwFGXXa6cpurDG+ww2hoph4ZnLxcWuB5lOI
X8OuVLd2eyx/xjJnB1f/VAUkLYujbM10aA74jpkPsoZ0M7Qty0imQqgtnsTqX1MX
2nYHpkHxmLznKMIklLiSJR44Bm2Ff2tts/LHQI11JncYVOaFl3Gxv/atiKdTC1FX
qSVQ3c+liiI2Dj/bk2RlnN/tAnPHUkJ8mIRlLYGI6N3DOzXMzCq/7Po1l/GcptXX
Jtp8lg5K+7o0J6Y0o+xE6OpQNB5uDFgTZ2sxTkbwUSlm6ov7XnexMhrJ/ZJ47zGp
27OXlgbzddlPwXxPELYZV4bXBMkGuFD/Ftge0sDdkvdbsAOvoJUjEPDCZ5bQ7bMY
UPpcTzMJzq7ICxXFqaH1aJiITBv9ZOZ6KLw4bRHo9YBQgM5xAls8QzdJWRXJwuc/
FmlQStVqEyPvjaQ0icwEfOXdZR+cpw0OYYXBmyBOR1JKDPLHlj/jf5kp2+oMn9Sn
ZSUz7AWt23/l4an+9ejkBrSbkggt94+xbh4n9x0/ueeIrYVsqwnSvQBvlkED8Uqz
ma0lx3ih+e8XYuIpZUt3927wqhiHQSbmCuo6fTZDLM0aMbkHalXxUxpcPFly1klA
PKMsojm2wK1uTyZVToTClGIQa8FlwWot44zaOWwwWajxYDxCSNPmVPR4rqbQlUSh
sk1D6xN3kgJjquSs7R/PYkgRGEY4u1c+EQBPQqN5iu8RwccACqLhcm8HXSi5MHRT
/6aL2k0N4RPjUtkdTniBv8PhbrkBBpTLGkM0ON4z2pduOnK6CpLNgSDSSLYQGOHE
1CuqN6EBlYljr7N4+i03I8q83xe07fbExPj49b+YYFwkuYAkS0VLEeAuCJP7BEf7
IcWZvTAvRlj5g5lGFoVPFyVf3+2kRfBwWQ498+oxbYTSGoqCicrBsknGsNd6kLmp
uCDjawzYncniBKKZVb6+6LQYiYnja1aXB1SAU3MfLdFve21RvebXkQ4yMwzB2GZS
v5sk0fYcO5eusEsmUb9sxhuflpd4om5Hw+0roKefnx1R3phX2g7XJcL5lhpa40fH
j2uWfzZ3MS6cy9TmVvebiKAaMympr37lyA4Wvnp/49OEb4Aj0Vs9lXnrY8Gm7DeD
PxW3jpG8MTIhCJfjAaCVlbmsxrfxMgIEARYeA+Iavw8lL/tKOjTib3X9dRnzFRZW
xAcqByYU5da87vVWUvBIKwD3L79NnTHDggGe2WpUPOPC3IwbhaEEM9ps32hyB9IV
LX3cvqjHN9cJ8k1vDTPuI49flqgqToSBVxqMX3fzlBkkqv6s3Cli5uCWgA1nppv4
RELHgJXfiQqGsQO0dnPiEBWfVekNTgxnN6tosaYs3yUPpDRg+5j4OwK6xayIezrl
D/fBwyULFmeDcDHoHv1DLzjp3QviLYM1EOL0sGe6uAEzG01bKxalXNtcGOKtcFCR
bjYTBL1WRwkiJZ3MGBgtIbw248EHZZFlxHTF2lT+1+y1Fa7oZ31iA7vz9mYMIimv
rJTkuk5yCUavE23SBFa/HC9ld66axkoo9FFm6iXZJw64Xj0SI184XLXxP8i2msI7
s2o3OMGOXLwzWHDI3reRfuR0rLyfJYdQV3PAGOoiWyGLta2WCR8EJdygOZSsvRll
2wxrkXR/p7idZg4zqmUY9x46V3jhrg/GhY6CdwBRIBrh9iyKbstyPhLmIsYToCN9
ST7MLq2wlOPmIIhhpC/kFm4BodnYhwmzI8LVbeHULaHqAIPWgrnr295ffKTJ0jRC
R6YfgRIqdM0U2CkivTk1g6aYndw0hKlIOWzgz0rwE3/5cLWmcErCy5ZSHHM/vf/I
4FW9Ln44UhM7cy8v15pGDxAl0vEnkvN6mBF/+eSFyDpADf2zuiAonypJW2IIVLr3
gksp9yCsU7lduKLgzkTV3W/f2PYlUmZ9S4QvdxWhIi5Wb9/dSg82E185NELIQCyv
zG9vLOYNPnNxSLwdnK1vM7ccGC1mC9KI5fGAh6dntLhKPOBkH6iG/5/HO5iFbXkL
0ubr6AFdI5LrjYgoXvPRNKK1YSP/5t31CWfmGRAVGJYqGyyTXRjCu2OvHYFzLU4n
p6saj2E0Hl8cE+ytg/xp8Xb8d0enA/SVdDLDbbXmV9TK5fGg9rk3LYtqKIJbwDG6
n/0Voy7uWv+ezbY/ZhlfvEsBjDSV8i2bnFblhsYst/dQgoQ4w7Yf18OMhWEWAQe2
TMuw2QVZkt5hYA14GddRpNyS9K8YcGnqBp4hVgVRlVCwdl/CSoY68SvtCVWfNHUs
fWh3/2FtIX6odUkMXfkefgGgdI8bpUGxTM/ZJCD+AujiHHy1W9nBFcVOP1H59Nep
X/6w28Vwb2BDCGe1cgIPJz9TqMQPpHRqkjwbT7n1/rHyMT/YzSXKbYlpf0XSu/X9
L4MXCiR2qDYJRzlmM9MJFgXGndp1PqSmDz09K22clgcqzU/bfpMcsBcsuCTd3+Gm
G3zDISWyY5sUGceJl7e9ME973vsjJfQW7ONmZ0XnQBL9XcAZcdF+607+iUlojvA/
acJgkLM0aNLwVL32p/x4sQE8ZtKsuwZ/HMR/lqlwdWhTQ9vaxuEEMF3SNuJVD7v9
ghK4mpuA+HGVW9JS29cOcSd0aWyDiuhBdBiT9B59Quc2LeDDHhw4NQz79qwT2kfH
Q8sMYBCM6oLmxnGXmF5QCJW4+0f15Kri8SishQ575y7uOpZ8mjqJyBm0bAFLEudx
YPcFQ6+ZJSb20afrznLVcjrXWiXDi1xaNVfORVqtadHnESj5MFbkDiiKYTMcGsZ6
2ulWhARXnrjjhAH8xCk2XX0XW/ur427KjiFgvGhwGoiTzMcXikI3V/aH8joeoI94
wt5qQvh1h7N7qnJND2YwBgOUI5asP1URl0sytwFt762pOzguLsuIxj7KHJnDSqwe
ikD0YBAX6yQq3dckfef8ch074qOgWjxQrq8YuuaW59OU16E1OYtsei6t8Z0o9C7m
sZNe2l5CIZSMB7XakExbjVWfuYGtJX+e6h/JcHVq+G2TiaKe+AfpRs47afwgCnCe
mkq/D6PIVu+DAAFH8iWW1dEARjuQEvRnoSzAzk4aJQgQ6JdI7wp69GvbvEg4Beca
ai/GEVuZ66/GYaR0c09IIco6kKzlFTW49gA8CiX4FVB5mtUQE0hflBd1piYXiE40
3Giazb5NrfJm769CZpJcjLSJmYFWrk3yNpex0NFUmT0J6AkK0M+lo4s3R1RapZza
IyCqX7RmZyEyzgMXiSTM70diwDM2iqq4pqPpoEREewG5hwLLPmFQoHel+4+8kiK5
HQmqDXv8iFdI4nt65dWbVCmwdatLDThlSAuY4q4tmB05RfjgmtU6dwSD72BRTxx8
kgAOtzX9Fz1qVHnIOY11PIGVkuZVS9zaogAV//J/diAtV4wM7eJNHp6IZTebxKwm
UZzdG+QtWshtAvskLxbpEpgBOmgaw6b+3jdENsIsrWdZfhzctSF+F5RA1+GS+NHg
PuIibJqup+BAA4Cc1a1oDY3fjCjmNU1l41v38Lx77ZcAC8OxL5Pk94wIGr+q24Fn
m6sb+ZRsReV+lgC1FNBtP6I1y5eUb2tE6l4iURRoR8THoJ/mB/Jp+tugs+9kWEPC
+p5AOwefnMpJNNIYnv8kMks4cWB6pA6qTsGW1CS6hljOwuJe57omvAJO8Us5EnSo
bpHpLFPK9oY+jKsmUdfjttceIb9wL/OaJfpMdJRoNLrUPEHGfUEnhkxdyB0etV6z
0tF6WK6ze/gspTUV7AITH28b9O4+tnqEpfEkciYujbs2R+p6OhCS/lTnYingpvw6
Qn1k7odeXVVgP+Xy0Xhl/iHpqSUK1KUnPZlBULVuDB7d+X+D7V8xe9cbsRfvPMba
haFiHm0EiyTcqHxW/yAClm/3rWWwm4uDUc7nwLJTLDkW36S/v05dB6zrf0fYqMdi
uTjJvj3T3dydts5VDwX+ok7Wmpc/U2Fz4mMwJBr5+pzVGgPcDdy6eG2jftLxGE5r
LY8SelhvjcHBxmS0T6QZUeqQZQwXwpZI8DV2wj3Yreyd/e0aJFAanBlaGOMLQP6j
ekWBwGPRwsnTKxe4YoD/btIL7R/2NRhcF+kCkW3/yXG80/aytMuGxWUUB8RGFS+2
tO3ffvzllYPFbBN8wh6lQCvybUhVqMJ2g0RIbxIi8mUieH0956Wmys7Ta89yK0jC
Eifxx7ijvk+llFAs51FNJF8MvajZXxlqhBKcAlhJOnLGWUJY1beb3BG5i3wN8zye
rYu1LpUijCq+Rqb9Fn2edd5hkYUMDiIrlT4vag+NcQ1bKn95JY0bqDI04RIjteVw
bi3bTbjTBG1Wr65LUFrRK+BG12yD9YtR2Vbb3XyO24au5DMUzQx2SumT81ASbj22
blvt4eROty4FGDyRuhyUFcUA2IguK6U1GsOcPkbDHCw7ICImS7Z+4AgYX6E0uUPH
XUO5upG0DJxlNv367p5uqsveaJ9OLD+3BxbEzghohH65UXVACJzjNJBRi6opJ1Wp
K4bR0gRlm8cY7oAYQIJj4mdjB1iJxGXRFt078Smj8im9gC/4GBq6lGWpWHKEI/4e
VLPpSpgy5LaK3ImsLypB7MeCPOFPOhJxDQw/0nuaeqs9fq66ibUkkHb5m6wZ32zA
5/MsXE4evjjV9xyZsL6KqWkKEXq2j2e6L9gc/4dxXq3SnsXwHotwo5ymZfhe93c+
BeOTOoBSxvBnv3J8CshZD8ZCOajP+VMK68Y/Pv1zWdvgEHYvQil9C/5LfunPX8JM
EzDgegOj8k6/6GY60XkTDcGDtcR9x2QiGuCA4W8tSpB6PFqzQMcyJYqhu3nv5xEa
klxbjLvyPLQKjDvg9JjoUxVV442dUYc42nP8lqtwtC+nf1dsbBdgDpn9ioESSGpm
pWfK4Y+jgBpFbHWm2o+KrN5y2u5v+L/p91W3grUI3lqlvdm7MzJ5CDudzUa23tVW
/u+I0Um5dyEgFCVN3FlQ2QbC1n6z/yZlj4GX00Oyfru0uxpbZupRxMhWUPVGoZWT
7kk4ra3NXIz/1SfrjJLbOLucw/XQE8i0OykVmEi0h2LpP2wgcVQmPdHoOcx1/TKo
vM3vL3nEsJ2Z/KqIHabZDqWnECd/YjgmerxsMVMymRdQxfzvGtsTbRvZrJKgkgGN
R6W3QOw1QnDncjVW1Rr0lh84+U0IdyJpmx3Lz+KUAqSQ+CiAKMb62gj2PsAUm6Nl
YytyjBzSolGV17+6D6fqLeNRkc7EpswqLyOfVU57q+r5boSWQ17GBtOctAUqgBB1
UBGkWsRZfg9nl4wjEgMtFjoUYeFQubAYE7wNORq+Df8ZqRgWF27qnYvl3Cw75W7u
DUlGUwz4HWMi0/gjGfRnZnjorAx4CbwMdO1WoIAywWnUsqph3p+IGQWIukA0MKpj
W6MbotqEYOeEPMJPPmJ8kbEXYv6PDOad+/URJ+O7Blf1QoV5lLaRRDhe4/GBXvKD
ctREvlIvGiuaIsBtvz1g+OhWNYt5CSdj4EK6SniuDVWYwWg0ZT8T3uYOwoyRUkeK
N0c80BrJ+kFcLDcQGxxEHMdsnt104mh59+IXscmqG/zS5C9UhmVlwXrK5cnXvr5Q
18kpogpKabbED3yWfK5aqUR1NBnxRDv1dNeOTwFMNXu0XrC/WFZ8liucSlg/QSNM
RwYkqWsLYysffIl1/P6Wny+JVWlisrw+oOFyNue+v4umUwKa/A96Q30u5OwjgBAF
R/9ZXKt14VHvzYROfOucDTVtXgwdh2jLlx32raZy8iXYOOeBR6h4q6rphCN9t13b
o4HVUO/JFsvLJ/grU0VhwG3hQ41ByjbeKeW6qQswdjk85DezsxY2GKu1+MggvR0k
RgJ5dJM2DKaz/mbuiGVX0fh0qjv2SPHX3BjvAh1HjaUpfUDRnnYaBi7NZuG2krYL
GPQaKjciwiYWaFWOWVlUYjIhaCGJBe2i3FCtXVrtQYIOIzuNU0XGKAIo/70/PVoJ
TD3jTmQtONM+0xGi4zEyMWi7S+asuuyO+0RnnFTw+jRUzmtYBHtGaQ0I3ol/DCFY
C4JN5AQvnSQLjp2kr675l18FfU5svMokg5mhKmZ5f6Aa2yKQ9AnRsF4J29N1vINg
yHNuEKJeHzbJ0Ngo5PLW3i4hsuL8WZlEeugn6PqcqKzrsvGkWLbZoxYOy85S91zR
qRF3bkloNJg6+ctF1pS7mctBboJnB2TXGOwn2UkTPGkzaFGSVeBujNY6xl4v8wI/
V6vjWLg/M0s8lFeA5hjQmlcj+9T1Ix3ylHEDhenDclvFGsp5UIUzn0NYL1fIZ2/8
OCq8rg2MBom1WTzvQ0TB1A++phxkx6S9iEOhq5FeT/KyWLR4kxGNqlMqirefPNjx
R8L2EQa9mqQanfa9tSAOwfcoh26x3KN9iUnTkQjdCw9/vOK8ufOGPqs6u3DGrZWT
8bvJxWpIWttcEPR7yM+3++PElaVoKbOod4CjwyGzYBwym6IAi3H3uxcjUlwdGdiM
IPiq6sVHW2Iswl0I8KaezBErMWUwmFTtfBpgZidw2EEHSnyF491zSmph/nxWu5+m
BS7hk8Ls41AhiQT8mdAnAZpWSlkgNnrLU/qpHhntxWt+Q+gb7Lq+B3ZuX/zSXmxZ
Kcu/A5mvKA7tLY/4nVzESXXxPW0474hY3K0Wp9ObJMhwPZb1NGNNVXZin/itckFS
Q/QbYA0nVWXCGA1Ri7/CpdQUXAsUk4L/6hBdnhdQshejEjcajbPhQ7jL4nYOjgbf
52f1Kno4AypIn/2TbUo7KvMnNDMPQUYi1+QN4YH7sayDF5feMUYX+9bRPB2OKXwj
06SRkd0qKLioBj171pzKcN43rwCYbfF1FkxnVsfMpDV3Q+y/WuJgnNpUbRJzVmzI
UXwfcfJ5nj0BWFysUJT8l3YMZY32KJaIrxE9HDC15AFUmLRb4cdIcduwG2G1F1T7
xhLh3Lqzc4QpWD/N3DbwZAbP1hxwt2DJw6EL69Pzi5j/KSWZxYK5wlRY01iUeruU
vmXTjS19l8udXNU7aOc5mxcqmcYXXKWctjzLaSrGxdVOR1ql/1mK4s8GGgvjxoqI
QZ4MFjDBsuSpvivWqWw2mpBloiz7SiK6t8IVHUO5dPYwcvIX638tOHJy4vae2p1z
BPquQ0ggNkgyPe54rj79M7LXhdBVToEUOiisVNtsV3OFR7RK8mmGwNumCW4FX7qz
v5/Mzpb+U6HEzTNFBBJNLrWDa3S+iGLfhYCAZSZFtFktpAKCN8LAVsKzGRNIZNqc
VQT+NHTFeB0IYKQJWYfX5E7KAPaDsQoh0EX7ZOO2ciAutBTh7IdG9TdRGucbaium
cMbu6UYdOjIFXfN5kFlvB8/7t4oKFcqslL7ChuW15mnsVhSdwudT8secRk3IySKE
1kgNxEAmeuaj1d0myAaWLdk4UZaf2+xKeW3PEVTNE18dfrKIKyj/gjjpiFmpo39l
lvCEChrmo6kAuX2JIuWx33H0EcLvqjYDyg/rliqBhkpAVf5Gkg5yykm60tavUIAO
EjDY/1YDvpj43OjU7G7ISkR3M0ACvjkA5+dywrSM/XYST8XiVhE8YiD6q2cze43f
t56xMV2Zt4jPUFt/h0Gvxr1hfjHwyC9O+BbeNHQMzpMDmpP8hYIy14wl4xNGayxD
GCa10GErcbahLrUbXq6Wy8gIiiRJPMDh0DShloKknzB05pDuE98SAEwrvbkdCjmc
yhvkxsg5n5myRTEF/cRYtUhudBVH5fLnxClANeS6e6xSGyNQARLZz1qPeeSM6ICw
WCEGg8IJRcxz0eXg7YJAPrpWjBuhzvZg631zHKau6Hk4JtD4UkSaVH0Wu7tq2ezu
2z8lWvnuuAjaIM4xJ21wS2v9h6onrKndxAXafN3utmqGT7LK9v1FO7Q6S4Ic3g85
upmDV1MBAos5xlSiAfiNLJMyKzm719Qf5fKUih/LeJ8eH/2x+1V7/0QNqN+GQqae
vy7sfXnTT+SHaWsk6PUYU+B78+g3+2sgP1tqE1kkBzbL9oozoQRlREQ8mcUIiBUp
wSk+ljL3jgIQHiApI0QGidDsEBTV0Wk+WIw8+7T6rKNjR0hrsTkYHhHNRSRz/moA
42gRDQ/0DmJgJlHSWTPYKFTk8hZHWmP7hlvzRN01mEeKxUDgTm41lwywflaTccu8
Qmydp2CXfU2QhEf6n9B7jnS2KpTddt74TSkEgbS9cxmtSqVOPSkU33XnMvDPy0oa
uGFTbEUuiej7FnH3l8FGKXXl/f8Ha7vPVIVs8PRWHspRK22Rb7CJukmzpVOT8lun
q8AdpMBcEQk+riw8rCxgBd7zoCYvoHFmiHTTLHymkfFWhmB47BvNjtVRWohCFY1V
6twxkmHROyQ59bNxSOubjPKqXeeXa2m+b1GxOErmPjaD9ZcJXV7xMXi68PnRQIDx
kuiyJIolYz0+EDNm7cNsAXD7yt2wkXEzu1rzq/QGz3QarFPRpMAYx9zMLwtS4OrG
zArdACQ7ELyDirWTBM4ntambC/P/Y0JgELdQCfOO9W7cIL5CPAvb1qT6/hp7e/dd
+NhppMtwmmkel/TvLH1g/gC9gJpX+Irc1y+z0LlWD6oTx7oe94OT/lgWMP4vjWqF
ztEheGFfdZXrHDP7NuDE3aP2Dg8b6fXGybw9+ap6XC2A4LmBfjw7GtmrF/E/airG
ZrMadWDkuGK25czAJPcI3QfjgOCrhsYd94xSiPDqL9Pt9BehCDHQdmg10yJM31cP
QN4mNvNZE7VGxRROrvT/ioawViQlsJfPHu0B7z+PUCm9tzd2UKg/XA9iy4+MO+zM
QZ7gVZGYXOTlmxgwa1tGyoJMG48F5Av+oZ7C7tVaVMfhXr2zsQP/9KtDFpZDY4X6
ltExKifEKS+PsH8a3KxdpOtT8FLVMowSm7GFm6mXSGkcCJdQq2nKz7HU/52vUMjt
IMrQDTP/6B3S5LWE2eonJbPi8oTowM9MseRelQfZ18/zQjpmpWIqCVUgSeWGh6Fn
5gXYmMG723LkE/Q63+vqGFVcaud6d+45aWjEzv702yvqbY4VXKTA3SjbWNHJHWWZ
q65UKr5eH10B0O41lMjeuKmWy/jl2jmH3M0Na81CpMLt1042U2M4iKxpSyeVo+1Y
9yH26mVc3zzAmpGHalHGGumYfpY0WOlXm202Vc9HzCr4fPPoxRbS5fvF3fSWwnGp
0xQGHJzlM22srbDFw8wkjArjf9zg4hlXEHN0qfMhU6VhPF8WQoar6yNd+IPMhBNk
5amUMIOtTbfylapwmL18cLHEQMJKsP61Fi+HNRshyZtCUHvZnzxgocBfocshoQrF
Ob7XHRIL1zzGBJVJDvM9mdcsM4vDNo3x5LDscpzJDlUqN2OLcol+R1nm16xOOjdN
XiRQUzLdmXNkyCIYw2ssGgMTKoFDdLcCsdZUEP1y/jBGFThTQZQvZzoJ43ADEvtD
zrGM0f2qxJd6FJ7EwQgjSys4BiOcPSxiWdih5LtAdVW5c7+julQxjy3fIWK0ECTi
kXhaMY5Jx2ShURb39hG3uws+7BoIeBXo1HeOP3fRufQm+X8IGU6NMQNWI0vw88kv
itgBxYpwl0uOmSZi0kwbJaAjMasX7wmqoElzsy8jVMTQnclTjbrrlU8uBP2iDh/f
OpR7NOPIPPn4D6TZjwnOaavCw9joo4fyLb97My4une9bct40nBl27aruUCTfP6nm
+234HyY0zLWqwkRqdA2JHUpOc4Tb/b6cysUIVZEuIfwx+u9erQ1mW1o9SDc3UNbF
fFTm6XnNw4pZNReLJtixuCvQIHjIZ8NV8qXOTKg/XNuzEirBNoHhKL2e9wq5565z
d479MZGyEoKn2N5dtUy4rKlbjpRxurYJTL6z2FIPvMwYk3EC100wHrvbSHpVW77L
2/m5oieQbC3Gy5o2mJkm5osaeQLy0b/NLKUDXU6WW+5QTPF6iVjdYG7ZAIFSBHRc
PhHesiCFP8GqFXAae2QZHL2yXfMx1LJMVVyj1HP8v0gfkeb3mmVOb73qrMC9aqSq
4egfBbYrO6KJcNyEa+5EXyeQB7rL7AicFBHKshxksjFeqZthTkBzvjgc+Y/hw3pU
5r3/yFV39nCDfqf3Jx1zui9iBnQnj5w/yLiJNX8NgEUgBpstz2hGVGGrLgYQatmo
6u+fbXhGdsirJR1kGXI/3sTw0sxJlzM31jEw2HH9eMcAkv24uuqeWBbpd6LN0z+3
+RNOIxJ4sUWQOlL8kx7KZJ6iXSR2dB7YPxGx1fi4ddsNUpl/qn12jAPR+CflerE2
QIk03QgKbzPWj3iXxS5fGNphum+rlyFFrHbto1Ld/dmLGAN7F7xdlXpbSB/sek5I
oqZ+B2u98gdUND+yytnpBVpGUSYMR1UT4odcHrZ0bGJ+shQNpzGyDsBbU36o1+Sf
oqu7/PiOhfqWUDw+n0R+n5WGtz5ZXrOr/jR3bxRgNcDgMFmU7S1awG5226YpQZ94
+2DAu4TXLq9K1AceD55Mn2es/fKG6Y/z65KQA/rnoC+pTzmXwgWgNhPJU0yQb9Cm
YPx8CTWyKo4fm1DjaLt2l/N9ENE3V0LnIXCQIljK4D+uVv4Dz368u6yQlIqwD6Xz
HwgQkbC1WPmCz4t7NCwJVDk6eXxL2g+L+KWeoPo4LIDe8vvvwpCVhZS9PLBwHD+y
GV6qFvh4WzUJtnUTFjERp04n9+iuXnWejwpPMVXZrT/Q4j5ZefCGUN6TIcbSUSUU
wYAr208qZrr5wUUWIosziGpy00M3BmGHq6QNYGsr7QNhz5Lrrq1E/jXhJEYHALG/
tBWZ0CLW5l8FSdTMEweAdMmZxzqrvYxhHGimoXZNpwH5v4ImPA/pOVSQ0DlNmSjR
vjefOaU1lSWsYcualNBX0nk3Qaq7dHZCkYcc8jTGVjSMWe52COvGhx0bBESAYqHb
+Sn0cQ35i5FEhwOxF8qL98t/fspYTfRLcFso4GuH5vp5oFyjK002XtROXcf6nLbN
7EhSkutmNx8ZhFXj/+ExXJc5IRX4RgHWLDKaom1PO4iyt4iHQNSMvgJd1d+VRtIA
cPyF5g5Xg509UlBBpNvZDrr0Po3/cS/iqKicJm5pkua5lOHKNHdUovXEbQP/897S
mb9WbG1u/cEpE+RyD+dKvunEFOMEuI8M/so/XiWSsf9BUA+7NyJiBBUxyMp0D+D/
0J6L6j//vkZxd71eW3u39PpaSE60GmWlztm5W0ihDYHoKfVY3q4zQrIOSEJYitcF
uF/FcXKIaniCEDfGQO/jxBkW7tPdMoTDg9ah57NzuFhFIzFB+rpFkmGLD/t75sMu
BgbFHlZrtZPfQwjNx5NvIO7cqQyPa5plKvaIsTdFK6GgjIr+08qD5Hh1JV49ssbL
dmuoUI6j3xXJ44yIf0akAhZWdnuRRWf3KVOOEUIRCa4OCelK6rzBVmUHnodsXjVz
c7ZX5FkMe5XcFHMsOdgxlDSXqATN4/ycMMuqXHRH1Pmf3UGzl/yEUcYhUZ0syur0
dG2qZbdYGd6s+yf7Vqbm5YBv0a++z8MMWnDDUaNO9AcJHvmZJy3PjHWOJCZkEHyr
dxctagvI68TA/IELxUJ4qgl7YKghEy1vUQBmoVVe31rcKUnajMFq6bHTHuAYx2ed
GeLVQ1+RoOrU1RjQJbTX1cnq7zXxohLOtQGVXd5jJaWQiWloX0SFEJXtlcutx7Ks
7XYJz1buy8FLL5LBJBlKP3cMFNgW26p3fyOoptg5lEqxqwrKwli/Nu/3pH+A57fi
Xwx49syFEUxe61CDpI0y4Z2BMmzw7lLl+AAyaxrx3FQsCMO1Ma/nsKxQ6YuhL+Ld
KGZs5KrduhDJT20GishEnAHw3u+P42nnh3haQ5Lj5V3xfGVmBPFcU4t/d11vHcS4
JEx1wt1grW/mGzwyuUtt2MRN1vUuFvUN9m3nfmYDuU690hFbcsqwxADIjcNzLTQj
s6z09mWSBEBYlaiLvvdEb5dluH4qgOOuDOlw3nKzQKix00rGqLswacgEQ5CvtJA/
w+qgfDAPewDEBzBmU+yfDV7UrfHA8Ei2BNhO2ElmtFpamp86Z81vK92JodcRkOoy
IOSxfAyofvsDpmlO0ZdLKjfUOF+bmQPKO0fSbtArobk5JGeFUMW4HrbqG/QMQq3S
vjnzdCEHNLE7P/PdwVTqJMCKQsrFtEzyfaqaVPim1XWtseF9DGrNM+GjTzWVZ/Rh
oTbHcpwpeWxSryqL/Z/72EgH5aSrUb66vvMyuKhRY3r0UaR45DWpGmnZa6QV0zLX
SaBcopbjTg/X3NV7188rpIxBQNKF/u47HwvvbqR6Y/CBGA0VBlDu0K+a1crHiigq
dZ3JcT/5a/pWp/YvsV8g2F8gEhJMJLfaWsv+nxofUnizfkoxX71lzyRRvj2Xow/j
8YJnUiFXil2G++ttPVIZWn+4hfIyhrjk9WVQpL1P2icpNhn2tPn6FVlZ62M07JJB
y/EkVu9d06bZkcODg/8E/kMA/YVnhE9Rz9z0KzEb2cbEir7q1l3NdtzRj2140xt5
sVIf8j4de+7TbLgI0aAxkVlM69AsVQU4bBy6k9Yxhjjw3/nuQQ6AiyOH2L9zJi7M
I6RyqvOFeeOLnxz5rEl4aFMPkpQvkykrJmEC2RGqrGYQlwO5zb6bI9DtsoO0tIPn
/4qD7SwF8zMuP4DbR0j3vkE5bcxXrfDEPxqrGzLP+nowtZIO/wJDq7fVR1htWJ4o
yedBXfY4ZV2cdHDINyHY/tFPOWKITc2LeO81yLWtWJA3ngSGQV/RITQ1UEV7tYZF
uUvekQydA7SMBvGFYkJjebsAG+nVrZlvBBM7qP3UdrFUm4mYqeeugYtu5vqag2uC
HyOC7Ze5E+HCHIOH2XGN/5ee4ie2EKQAHzRiGxOzxnD0U3iAX+s6iBQVCc6NVtsx
jZBpEDelBjtQwakMZjDToULyQpYqJS0HWBSCZLsBQqpWY4xhmAJoqyO8UwctNU7Z
TgxJmpyDo6xAsnjymdLKKjcpPux/lxZ7h3iivKh7EiEFjYz7AChuJjRWZpEv7qgV
TBfyuHTDDmiiEGrgu4ojE5t0Rzwq6p65o2tLnrgRqO2IzgtK+fzZsYUBKlJNTdsY
+Z3PRR1ltO1Sz3Worf8PbLLJUJLIULf8qME3wjFqf3uqanbhYXcKLOX39W/lzI2c
C1gv5vgNrGK4BbcWh0dyYmodZ2HhaQz0l8cdWzGEnUJRCnMd2lvk5uDCNRD4ojq/
1ARnbo8KnOoXbilQEu6ilMQQt5LYvy0TQyx6CQsze+oVH6/nkXPyIVshzFJRWane
59UcHBJp+R0nNk0D6n7odygnJsPYsvr/rOnCVXtGd+a9ZqeohZIiZQCdQlYlWI7y
LFi/Xdzmv4a/IVfRjmjEk9vhDNkV3RUdWiKBg9p71Gc+xdNa8/HISPh1XrB4O0ZC
ZESJ0q+IJ+t9Oo4bgYPzSTL8XKQ9PfwFycxL3nCros9QKW65KkltCgyQcsG9xUze
7cZek2u893AAMKSHQre/qvj2AQvbLN0iA5xcZiDS0acBupCsocKMVEg88nFqCyHz
hZac9mlxd+opHadhxfVOxLXJ5sllnlYthNgIp9gbe7vLEEQVR7SNUZ2EQOfDcOgI
ctysoxpB4JYu++Un9H/znT/+b5Arz6RISdgFN1a7te5OV7V5cxb2LO4DAXYRHU3W
vkX2zSom5+ClJHfh43Jtu4whX8PfvrmQ7/3Zlz+74RofL+ZWl/wddk9DpoReeUnz
G5zp7Y8+eG6Sl2lWSV11zluvXPcie+n+/FWPmnmmvCTu2VN5abLM2yGLxQHN7mN+
d575Ce0j8TG6gHvR9qSZv/uTF0RN3+HrzuUYPDmTI2ZMFYXmf34Llyk1MRH1ucWj
9mtlqEPPkzGX3ntcWPIk6za7Y9Ehw7Tqlr11SJbHQ5l1En/W+TyZFZj8IDfpzYTi
HlJMPGJyw8CHwIxXyxJTNaNw/LyMTdcAt1kFxOghDkSCKrvGVmnPO2pMT4/0qt7x
R/6pP/32GKyu+Qw+C3w+hiLYysXSCY4V6xUitv638cHahUhCZG8WkY8KpFwA8y+/
r9iMDBJBAW4IM44fhbQXbNFmzJX4C/eYfvhz61WAMH4MHpqDjW/bziXR+jsvLqbx
C+GA/l3tCbz552DK6fTXOsgNRIad7DIUX7PHPyIXL1ZmzlSOtYiQvGfJPLK/FJeD
t3CRtiiyHGYCaWxvWzWrI6vFU0sdPvrfqkvNgbQVjjrsQx4LCuaF7MhfKdLKksRo
hVp9Fu9pzOZkKF4BxU+cDPvKMjAUgHbAPzXSQziBrLuPNELIcv6w27JSqBlTqU6R
8gu7pl/3PsMmVTGbzq1xC9ak+kZXEATkKVSTiQnEbI7DxZSPJrClIH6V+2CpkAhB
B6BN7qSDj2a6PQXeHJJ9CsuPNLbHT62A0mJPQp/Gou3C343iPoaoUPnu0rVm64oi
WYs7AfIvR1Maox1cfLUM4qXtNwL0jwsJQu8L/R94IS0FMof2EKacFaRtHKDZjTUu
DB8DwNRwysBJgHxomelLqvfJ/ksVOWllqElc/k5XzqAq7iCJZGj7L+JAvzRbzTMb
+BHcvueHy5ivLio+KzpiTU7Ita+Y5evZ8xTGwzXg2c/941zf7sjpThSvcaH013WF
7Jyn3XKlYbkdD4MeqLZODyxpDlBrhNjMir9gAsc0dN0lvi0HpDE4OryjFM545bLP
oboulP4TNPTKZcEPoR9L5daMQj4uNXcRuNAdTf2FTVWMT5h0PWyKf9bmvwwpL4nJ
tmGLNtxFcPQv1vYQRFxxxh2wrtgeaGMBehKvG+b8i1Ejobr4acgO7EyM+ow/o+1c
h9TBkoHfCAUeLPnPUkqt4N6n2dwTjH09xC2AalfZqefakVuKYH1MZ38nfPG52i86
H206Ce3pB7aBu9Wf7zHHuJxrVxmjrZ8fOJjGLgIAueMfGWkGMmF3qSxHUsHlfrZ0
d2iS1CZRLx7rdHGE/7o8xuteS8VPvyx8L0jKGwgaY6w9avdE25EEgvncq53f9J3k
FXSmQC1gKOhkHbHjHJUsrg6vmqYjkZoiEuA4M+99YRjaHB/Cd3NsjPv70M/GZ8Hj
PRmyvTqUyG0mg6AM2E7h+4t03sqlV8KUrJDbbq6fc0Udjo+jJyorA2LQ1U9Us55W
ZfV2QmV4bmVZCzBbuiDAvjdIeLc1i/Y1oUgOMvysT3mBwfUPMJQGgu4IG7lDXZrW
/eHzJRcgSK4yhEUStcGPPB2K5hsYf6AFfisFnwDV9DqRotLho28nxfKjqN+XxYfl
y6en+2we3prJhkQQCKG87FGR9jsRI9WndPbl3We5Fld3t17po0fVqmZBJ5VWLT2j
fxYMbNGAzbPtE8qKHp+ZZMLGiSvZlEY0/0bGzCOz8iEsSxL7fuvDMm7QQaxBIotZ
JRhB7wvHUqfyEmgjpieEeNWufY6smpOuayqD4ID+wxm+eZKBIY4fb0eND2kHcdpK
zJUFI412BIt5nPF2Qm3hyMjV3ORlu59UKPhlgWJtElY4YBxDBFRB21xX/V1ymJfU
tJGIw3klWOf2n9Q8TlBFB9xeKC5AT8xNhj0ggMPD31G+aMMis9NWpY7YRQ0LAuwm
1DU3VTHpFBNSXsh00/9n7C3k6VFrPe6Eg4vqz9Zbl3/6RmNEzauS5q89XVj+nWEN
FYJrAMrBcRLhGM+GVACK4iTxdomqyt/wd/4TlmUhfdxZ50XLbYfiE+s2+109fNWh
KghWyYbR7DNZbEVQEVmQIAat9J1X3LF1mmAuz0eWMOMhIE4lUTApoEoYw1SDaTGj
gKFfvLIFRsuydCaWBYS1Fdo30Uk673rv844KMNutdbu7mLA1ybEyVMThJvU3ooyP
B4p4L4ufeoww3rbyD6+3F3lUpF+jSahdfvhXi3NaxPsv8J66PQ1RROfKzXxC1iTS
PgweyI5zEdXAspISJyBzoL9XSBjXC6EUuwsBoxRU9868wUEpKDh4UkSaAbkxCDSz
mw4toinJTiQQgY4UcrjwWqKAXjO78BpQD1LcYyiLYXRItrNZ2ZIopRDucr3LJluo
p2hQAImJcuGSzUbxnDFqSeY5ZWCcHSn34XfajbMmRWHK13SUYXV+IslNQcynrRnS
oMoafAR/ZMtYwMpBltpvjsO5vjJy/wLkvWEdWrMd5rC0lPM5poquYFswc+Cy4sfC
tO1cbg2ZdIV08D/BpHQj4/i9w3bbRtMKTm2BZx+mephgDi0rxFK889aSNLmvJZo2
hkbqq+6Mjzcul8PtqLFII6/zIDGePloybe+uRxSsnv4S3pdhFK45xvJ6L3FRO/WA
w/+vSsOPnHnXFyDO17yTruPxiFM28ydGL241euk7wvVFxstyiyliRgJJnncPY2NN
PhoyNTcrzDnP5QSqjiSqoXYYGIhusBKSbFPpIfmkbuidgnRlnRDA45FZIf9knrXu
eVtAvx/g9HSSpzNxWnSNYKKBoZE1h4z/sYi2y60zZinkbiTgRrXp/GxOVFlJq0fx
rQ532gXdvLuvbOvbf4KkKdxo7TNjEzimGqkRfqJYkQuPA5zs0BUTf0IXv6hNGL/h
YFmDZkhYhFFQc9n6pImHa5Jmrx6WILqC5OJYv8ZrFzTHR50GRddAomek4igmdXim
siJiEsBBKVFuK050gofQr2u/Y/JQBaSPV102zQGakMf6GSouxhruNP64X8wHBzGd
TgxyzD8ExPsh5OcJIz9j9wikImzobyk5HGPsmOgFzFoKzMqJppDgk4op8DaLefWa
2v2NTFJ8Q/SgXXzI1AOxTMbzyLrG3h1+uAkzdJJAn85z9vsqTpBgUbdQCpos/H9L
s7GTYB0Dcvfwx22B03HDABsuAVe6EdXkX8oNG915JdsiCqsmmmLLnmAk7MVbTH0M
wbLNXvJyMSgd05PthncttNXSib7jbWXSZH1tiql9MHNNXadfri3CturR6BccOhZL
LVuH7hCgDlQ0u6/GKAhpbwlthpUPB9VIMHXylmWJ06rte4nEwPZF/V8YG4xG/BTc
9RynG3MdGaheGCbDt0JoYXO8S7MV4kjMScw32mUwhcOAtwF0X/cyAKUqsshcvJP5
b3HlSCcY239tRWvr+0VSwBHP2uzvIm5KWaDFbkWuzvt639jsHBCxOuSClyWfRMeq
944X8PeJCClxkYc8X0i1jXZZHz1xoEnBI8Lq9sRIW6MPgQm1IaMuTMbvcdpu4oW1
7ulDe3ZXuSllVzNabKctRe7CqqxqG5CiHVW64EFhvaEVwZB3QR9t1oNZQUHlFMjo
d0XWFDRiU9M4CHmbV9vhK3M81jMh55mvHqxHuWmEwUacQLcrZjg144+VwHV3cRCH
90McVWX2HpK+81Ji9zTfBywnr/2861LradlT3sBwXcnblaibJdIao8xLR4DQlYk8
fBwShXYEQR0mdw4oOQtlvRSIWDo6a01r+CBLib+jiv7TTcxr+OWT5du5+oyf40N+
pGhIk7buNafQwvcF7Wsauq4rY7XRJQHA8M1lDVC0efx4/vuFMVNvL4hne1mgTrDb
3XHkL99nGhcAKwoH64j+wB8OVC8Cewaq9eweuZsUDlr/dADLAQPenWA9bp0y1aT/
H9JcI8LkbxU65ICLHi4FIfV0QKLKJTWMC1zjzImgp/IOMEuVu3Bq4TOcCQpy4QUG
0+WpTAjILTx/jPgMkTXjNaCjLCnYPrIhB/762z5HVKbQuGbgOarG5Q8ZU9aQtLWj
vIDxGKz6Nx5pIrhscmaP/jOnZfEd8isdhTp2OgiQOHMCYfrcm2/ZTQwjsUfy4kkE
HNmPlhD3bTED9Ra3UvCS0VZDyc9uwubtt0ZyYXzd9I7ZGPIMlLJQ9JrpSDr42M2Q
t+Lb5njSqpFHyzzxljwLQ/liFE5ivHDW3jZLIugpexHHvdXNibuVdPf7iTPSUKha
CwWfFiy1oUb9Rhhr2j1xSIP+hbJNqgprWxAd/MfxUBaZc9lQOThUdPuV6qkIaVon
4QQ7iBHvYod4iu3kMn58nj/TTjPoc7hrVsHG0kQ31M06OIXASxwv8AMXjXtR7HuI
yAjxjsyoX56SKWvglOD4DkaHlxJpxPFMt0Z8asmEsgOz1A7rdGr7T95hSXlPykL4
Yd4szBlRQjoOzERgQyBnE8/BJKXqGaQKI5Op65rIpabz68OTUp6O+mPbR9YTl9cn
hRoCE+KgR/z47U9ctTcTjutkzdbPCYiSYhJqpASxp01+QCt3v7wVT3EYkQh3s4qR
LRlMNtzKzSV1VkDVgiE+pLulop1Ir4UMJa9s2LHs02pLT0Cmfjta7j2Z19C0rQUQ
xXbYMPpmFZeZNOAAYEJTDPci+faCM8LDnwf8VTsvBIPMqV3glr+9eem3WXvT4ZlH
MjCrQt06fjs7uW0qF2aLLskk1tXqs2COMMbLXXTdPOEDY7Iq/DvONiEobi2oKxED
lDBRwaJSbmvTtnQbsZzWOKaC9hL5RKC7id/ApDaBNPyXok32DW2ACwkBceZlPcj0
uNrkvYdOfT5WOyIkKX6QjlXt2/4VEeXeker5PfYatSWFotr2lG6/L2kaHOojh7n0
og3Z3pPNgnUXyqKyIMwbtqVSTjX/WRrExh+oI6fGlCehopHiCL+Pn8fJWgjXIfAT
IN/VtZ56gi9rzRzcrC0SajaJ1j2NQG+LtTjTV5BmVtnYW6zABQwoZtgF/MQp7kwK
5lxZBbMSkhbHONH4xyMFkhO8tF8O1zXwI6zR/29udOs8fxH7Mz1QH9bQcUiSakqQ
GczP9Yl3932smi6AdndBySpdpGzues3EVbLzQMS2t11bXQ8at+RFUPuqNmjPNphg
1y3VBcU+lP+mwwqEs64mKIO1djjuGfh4w9B5tEZbtRvnKx0lHWI1d2Bf/MN5+nJA
Qm+MfMr25RU681h5PaYXw5rvkD+3yJbIb2BiJH17f1wBiDemVPCIPPg5PE/rjfwe
/YMHw28lgBawgOUzxySYpj9aFNAj/+lGiGta66Jlx1wY9xehmo7RoiJ8TnyHncTn
JLw2G8cRpyzFgyCY++5+EiZc6N2JOQcNtsHFH7IXYG6auHU+MDw00qEypqnBB0cI
pU8vnEWgbhvMnEoTXqPYCNZ97RpCtHLnKsW30sXiO6qLeq4ZoMLVbcvyvRp1WRkn
fjU0P4fUJPVmbVp9QMOmhSFS4yjfa7+u6+6SnSxVTzHPJSrYgQHHeWhPSA78zzD9
olN9GZwNjS1lLgTlhARm5f6d/GDrEToxt/qJLjRt+SJLtaMV1IgaeuLpUG6GvqMm
ClxHGiDrDHlvcDBju9BB+IFYFN33w9TY07z5omeHJCCdHVroBY3tC2AH1ZvwYt4k
ej+wGsEKfBRcfRI5UG8NCh3/uEwvEeQ7wO6Yw3PSdUgt9G90Re2YDM0g324K6smT
1b4UIgH/bLOrowt25Fc5pZvYpITVzAnztw4P6rlS+hu8RXWzB8rkjelmYsVMg0JQ
L3ubKYq+LqP+v6jZBdjrmiHaTuSpuxJ0UAgX41ZJuOCZiTuTpgz+4zPhOOWfuwCH
4uk/VSDoCPoG1dkt2kw68shdI9qQIh8ZseM/5H/5K5g5MP5Pe54YZP18N8hYZM5S
f0SBCGAI+99STzEJu0r4aHTgT4XFKfO5E/Gjkr+3Pt44a7pGrHFqvIio/zN1cl9q
sd/2sHcqe/YjIU2fYFlKFAQwIz2VMxDFuKHEQfOYCkrSvt5w4sOUEoK0JDvYow4A
0uiqTCCOlwxOt40hryB7mICxKD5Bor+U5sZmKDCu39qL19XNr+WphsnIv4TGNTUF
BI+nHVSX9CtFbuHlpkH24GTwLT6Rkh3Vs19fdHVFmxCx06cHLztGtcMxhzjePhhv
GH6nuLn2GFRlnRfnYQrxsfshRHKZv+PeJQM7mB0mEFQiUXT2baw3nq6jKlIntH9r
etjjdL682U83HJS+zKYJI27DmXXjoUHL9wiCtz6WMISy+Vejbvm8U4xhd0ocMcAB
fwuMug9dkvf6pq/ssh0LwwNC/9rmV8+fw/cpm20k9ouK/owGC01S/CusfsJXXeq/
xfh+vF66ZNZrUvSrVyJFsFXJzP2yUU96eLUL4Q1V9ZR/0uAzuBQW+LeYySLhRszh
iKPGNTxliKBU2VuiOY1c2MCoCYKCPm5MqC3FSsdHHyQjIdGQcRtlwN+zykw7Zgrs
Ze1K04yE+w8TxgMQBmwg3DokZ7VcsKNNPuFR/vlKOblqRbTDQuA/FbRi6MfCRBXs
WeiiG9oDx2ynTTcXXaLI4bqpj7MPC9YN8kE5xwIC/t7IAn6HUOa5FApImfFKHY/i
hldaxSUdJtyyrbCAXE1uwAjJFt14NqhJE8npJa1Zn6gzu6KY0vDqSx6+l6llENh4
IAg+6Ab54nO8itE9BRQRnn1MEl3KyIMRJsnvAo1FnmpotW576+UZCxSOzPga22vL
o3oRKtLVl1yYL7wzlRHtFbMH7F839ouMzY26S9Z/wYYOfkxtKVDKOPVbH9NxD6IO
Lu2GHrOndN2nMm5Wh9ff6UmfVuM0hot1XxbXz2zB0Y2oSPd1HtbwuUbwdSydnf1F
OJLBNqgO7pmQ66tE9rxtr02HxGAjBrUUSN/UYrUiSdk+/fYmr2qk15Lyo1Y4yhNe
1wxShM9r20el5/oJVgRej0OhUN80CvDNsa03rIWCjr+DO07m7wjWJWO5srx8uALY
tyV9CAnVHtv9ZdATQ2xLNaBV65nm9CHtPofQGS0u2s/PY49M5qC9BfLXrrh8KT0J
C4W41v6tSb9ZWAatmxBdhFQ/L0Gt4uequKPPzDMrquPRSasMw9bZNwYcoSr17wxK
O/tOBbb/1AL4rIycIlfTInSN1AkSVmAYHKhHg8p4XfqEJzCEKfOUbmPGV9VzlG4E
SwwQRvPrSaFgoICmRUC61vt3Ep7MyGYPZI924RmUuIuAnhq4aDrIKy4geX8W42IQ
H6k8U44s9jutDs3boNFv337VlZb3LPsuwWdpwyfXofBXSdJAg44VJ8wJvdR4hcoP
1ga2D1Mx5AgsjefC518Ab51bjN4V2OiR89nggoNfbAM1NPM8mfnf9gd8kZqeU+gN
qnVL8coPQ6yrJh0Sxo9irmy3FDPvExJ+L1vpsj4NFQpCSlOyvw0HE2XUTHz8nu3O
xsxdbMjTfEtYWD1KfiKLT9FU1RJoNEaCoN/QBvcIVHcKsILOrH3I3MYv1FTD62sy
2qNqFxoNn6waIniBZPtEqVb5eRnzmcy73xAGKy3PlIgOAj4BzlJyKvCbaofspg0u
ljnCzm2mK1W5I4543JwK6gkiM/icBfxXy5ORBABdoZewM8mJ+8HaedUUr3UoX9Zd
dUVfeLQcbgTWceD86Sab4wlsJynuc46Quk+7L7e5C/SYkEFai9dLk4zE+1oZfyFP
ZthPLdoXzCoH2Zj1b1P7houRg0B7kSJ+HVeLKInVo/3YxKVYO+kqstm/LP4TsQ9I
TpuUeiRZNtHRm24hwqcIehkaKUVe/eeAcgHfW/y2LOZEGsERe3XikzHBuv/Tjt3E
9qPtmZN3OlQkHqDRjRWWTvds+T3O4bH2EfC4Ok929dgJhAXnrxC2T2zSbTCC6cit
6OTf5elAn/9LldvSdAl5g602+9xDACNqwWloUbuSW8cob7ZXdorVIgGomobyuHOY
eQnm3pNNlPBdqC3GLkrjqTCLq+DKgTEDYFgih5286jsUOnBfadL45udb3VKXzmdH
UTIac6Mn+c6JYkYreLKDRVtjg9QO+5qCUk8XIeUzu1wc6uvo1KbhuQZxqeN3z67Y
lWZfSYTeCcFifmFGUQZTZKBYhlAExvqk+XTY5aO2TD5CVqC11/Tlvc1sCUf55f3b
L4F1uckYSGLsq7M4xehe5bnlCG+IrQtSkxOTQIEGS3Q1kvpGCtv08Z/xR3j4wsTF
k3m8sxLqS3BSe3O1WJ1nw74l02PsXj6cSSqKSI2EtZ/lg/ZOll8iZgi/hOIld11t
XAmoDqL5Ofxph1FSglkmaQRtxkNJI/Xok8w4wcxdii8Bwoa34yrN1UywinqaGsXH
gYTbENH+dMvvKa2FJTW86VAQvZXwVcXYBY+U7E+SjnGkXFpxP6tYDl/UutUNf8NZ
NGCnwH6XSOt2XTsXCoittj41R2zz73OZc4FU2RxTXRxC3Genk4WyFlltSmK3C0VB
uvMQswFDtkN4ZY2RwxXoLAjUK8e9Qvwbje0HjD2RH8fYI5J+xOGGBZWt0M3sRDDX
Y1yqFMxzG0lqiBlGG7Vvf5+NzYwpwErtzYMSl38Po1IKKVSO+Guni2/Mltp6Z3t/
/GHsRkmsCbaAjQ0zL109kLpPCvlcKLynWtJSgTrXpLIXEHM1MVGpsOXPTTARrEys
/LADsZo9yYuKllozV6+V6Gomxys7iWjaBmSrSpCqnCdNTwTqX0BOqPJUAOQ7V9LG
Yp+BOSFnqRQm6aW9SakAN1d0Jh3SQY4Emr6mN1tQzeX0/lwi2hSOVZJc0/DMghCc
deo5Od6p9/SlW5GhRnl1UHN2zi+cq8mcLxCTjri8Rag5n2yAxKsQjY3McK7+DkV7
8c82+7BjnMWkgRtUDuCTcHd6uE27oYSF13fcljPtQy110NV8GRSftmAUGyu0n0ei
J4WezwFPtcuRdBIh3s3ijqD/K4bhJXCfPBfIE5rAEHILpHOLVBCOKfhI0OSwHwYc
w64sg5SrmAjfEr+WB4A8DdApm6YpNaf0xBYlCyCrqDsS6jdxxRCEum6Q7VWYdhOe
/wAcSREMtH3kNguXe3ZtApaQLJZCThpJP2jtGjIVNH1dWlC7OCIo9H0/m/xDgDYz
S7s/CHXE+a6Cb413ssp/AV1b5RLjXcqBg1+rSOVKx7/+z1ZKfzuFOS3brDL//RQK
hLKbqlrpwJQYIBQ+yRuImyFsdLwuhy8XMqmKVkpDwaYnGROXjigZj//k8Pzyr2CO
0yG6Aa3+PwFOw9JaNgyUhTa1iZyeXfkZrBzbQ4A+IjodbIfI2GqAkSmhr1zRKHUy
jB6HG01vYMXkfe0/LXXJxlBO5t0fmBPmyooHsinwD25Lejjk85RK5W3VNT588GAt
dWYs2jm9cb41a7/fMaPRKUngUqjIcp/brnCGvWSW5ix20YAEsaP+9Cv7XO+sBFtc
N3IPPn/i0TzI4jwZ+jowHtrF42QYMYc/keBskJqlFF7cMdRU6q0zG0NL/vBirKmC
j+xr2hNdA7NXDkLVvrbsIcZECkTC0WbTS4NbRyZcJKuITEc07mUSNvE01lFjNpfd
sDlAw0kspn51G+gGGQ8JTCb5ABymfm8U/c8EIZty0kXT26qHnXImM15Q0Dp8O1FU
Jd7rvtjrTxaD2acFkuST7yrIWLIK5v4+Qa893FqWwpoZbHsUNC7FZNqgp1tOue8Y
Ct1twKnDREr2nWORgXOFwdP3pGanOqevnbz3bvsvY8RbjQj6B17bOCbDlRvsBPW1
AYgJeNER1+YzKZk2y89CdJhn1kHKNxts7aAlO9vgtTC+R09XHEbfZsui/eJzQTuu
zPhNBELBS5S3O2pOqXFD4FC5M3oRxzJp5A9e5kKk4EBdXedJ8FnkvD4WR+WswMJP
Fo4/ArNyDSDRMrqedyWXVWV22fSjeCN0cV8w7tJcl9KJ85uNr+nrgs2CwOe2LDAv
+95hOUBhZITjnDK1V7vsOt0Gv1KLWG7AIgLPG/RoDOPYVbr9U92Vz3V8TbbHX7Pz
fZsDu/FW4ee15V4x+F3nWCDtZUltiuxM1F2qL7bTM9D7FGjpfckKGrboLL0qtATq
4KZfopyGry3YQOCCkfzZIKcTHs48sKuM2wfmO1bUG5H3vLxgZlG4ZwbDy+hFG8JD
1vIYWZ5Do3GtK2juP/9qU6NWIBC4+nK+Zr0YB2J01uN72E6QWaUjgLemlVUjE1Cg
+qN0+m/v3Dkj3koPnDKaOIi4+GwE8L+ZloCzRFjVFiGnMJmrybAI1ahhwkWp9i8j
hUCmbl0aTnVeSrq3Jo94fizJ2e+3D/TdADTWg+DfwDsobqtvnwMZwfb6qH3GLeG6
PHLBLezKHrgXKbfqyWxZE5FIguCqMmzGgTPKbLsnCBEIcsux5Vg4XDjlY1iEC8FG
38usEpSUplzRouV2NAaYiKwaHJImD92n57GCEBMxx7PoTsLBOvzHEi6LgZOOBqmE
q9O202C4MVjbMCO0jaPEIJwDzy4dr7nfeJWHR08KXndL0TNNe/1WbUvBYKI2Cqzc
Rqniz/QqRcFNjZn482/PMqJg6/dQHPX36Og6HKUqNdXR3vue9JQG8eoHAhrUdkO9
T4q7SIF4p3hL48akIbAiFcqIvurFtAf/Qmy7GukCSy30Otfc6iFTtcBBEanTUnNC
BwFhIc8ePNOYjdJ8FfZBox43BEAImZvJSsnQnbWRP3EcRlWS3JquFNRWoIGl+nTG
icX5YXKb5wNoOkA35qLAm9b+R4WO4aIiFrtGULghISjj3ILM4LDM5nhUgL0F1HCz
k3V2uHD8THGf03drbh0iZtb9zPyhS3aF7+D0OaflO2piKbhGaAq9ay8EiqmXAtO7
AxX66K0ZunomxPRrtSpWy2DVzQk7gHBtJcgsDfpe6YfdhZPwSK2UK6USxqsfyv3J
r2Jc4Zic1ZpoFmLSeZMJFCsJLXVfEY7ejWxrHhQh+eXz5TCXPDPnVtHrNPdLZip1
eu7zAFKb1n+pvEfgI3y2d7vtMa1hsdB0qXVuxdUKwfixJIh8uEgnpOFBlFCRAWfI
7FyeoJHHlCJSQtoMheUHWJQXcXvA7k9Bd5zgspiAlqfvnI/BVeb34M1muQynug+j
KGGuzVPFqR5mp88qgZM0v4amrbTC8M1ZLMLXCrwkGAUejD2eOjKlCYPzposVThhL
pU3YphRTOqPhfXoNQpoKwyd+256jkJG9JkVqQKcNqJFUl1eeYm45DEYHL/7X732J
7GgJh7L6DWD3bxAmjWFfhjjuaYXWtzhSnv6LxflRL5fyzgN421t20UeViTLVH3AN
CHRHtkP1MIg1emwTH6hlwvGKoXp+8arXICOL9H6bYNrgjzNZIep109ieD+9xNFHA
YDCH93wXyFJ+8+tnfITv3w4dXZFTbeGHSwyIpzLtQsfbM1W75mknvQi/GuOdtB5Y
rJpImc92Zwrubua1LCG9A/PTHiOEIDhN00eS0Cj0qVDFJXugsN6i3tGm8LJizbhZ
MI8NKBaOdmxdhJyFpFGqturLaK0CmnBxu2xx0EmGI/aM5pX40BrVav2s017yD0V/
4erJcEAIQr/9qwjwLQWleVhRSHG52zr4wBS2JAquhUW3aUBZj8i7m1wLUyVQ0Kr0
UbjrFoCzEovKf0RwGeKN4erzXEqjKN/rMfk/VNq0hj4RGqPZ+9vr/BdsssIBO2ZU
thkIDKWSUD4wmk2BXrSgQ4J4WAWWhb0XZPURNwM9fsuHgr1xJMwiBRrvkeKFmLvD
tI2kP9kbnM8NS2tE3kNWeNUyf5pJElKu3OgLNi2dQKLm2qlOuA5Ky0pgmaP/mFrA
FT2NElixcNNr+EQNE6QWvdaZGuYYhSXJDhxKbTBa24GhoH772UE4XRxVbejrJekZ
/+1Y+OmmKnKsdSL6OxyJprUs6hpLqhOQh0BpKO9LrOcwZeW8W0n2K4AODHFJHsc4
0eQUOFcC/mzZHNPiqUey7SVSJ2hZjpU0NNRk33DAxeXIESSo3xHlwkFHJo9NZRJe
82C5z8+ksSrHzvSmyGmcJdbTqbBSTSB6v4mZEKZET2gb6xg5z+V0sIsEC0bM9h+F
t/LNmsWyIYuxoKoEWgCq8ufbqRklBLeJ2SnjUPlkZnEGFQaOX3o9/EDtU3g71O/r
jJlcJEoR5i6t3roQTDU7A71VZbovHCFEnzEV8ZYSsPwfS8k3x+BjXV2ktZs+lruu
hQSzMkmVMpZVcRhqrDifzvmGafUOb6Vx5Dgy29pv/yHtlvP4ECsPOFKHyNX000ox
ZHAQoqeXU5fNknoZAP7WEOCqWeKqbgIGAAxYOYFHqTy3wQj0TIxC6AfEMdRU/LTs
hhLB5OFzW0+OC9III2IJIjLonzIVTjDVMTzWks5cpydYhELnaJgmrwrSZiZNr2bx
DKOFRYeK5sqs4vGF/dafSH03eKKfhvvMvfUGrvDLEjh5A9C8mPEMeZLvHbrBq5s4
CjnaWsvTdckc6TAMXKnImCMH2w5P/ghZT8pB+uP9Wx0e43Uem9d6U3wjY3uJyD4o
eUAzNLsarZ0yEn1eYXq5EpIfNuw7RwqlEJIIoI7Sv+o5N7u5OvMST8JI5mc8Xt9e
kCKPJvHW8yT1fIM9H+PYq8fqbTOIUpzfnxUW92KzKf9RGH5mHLo5ZKl9KMfckmpb
goLJbGMZre0gj9uoyVC6SUKITlMDGg4YhVIrZjuEk4EqVpodL3pKOx86OJyEW0RJ
Q+pDls0O1G6UKGpDWr/hCc4Zr6y6GSu4FPB5wPBIE+gpQ6LAdmeomIxvw/Q2iCb8
uJB3fKmnoBItDygVgyxGYn7U5PWCBcl4oRGaGBcoF2e4M3FAnB1bA40w2+Fw5WWC
513zq/EtZwcwtAGYqXCcgcKxTjnQMS1QiXNF/vRMc/HfWwbcV0gIjQcZlWi0Q37f
/iHhABWai6qoLfEJDTo2vDXDVLoyeS4KVCRabZAjIS+B/x0xi5RdvK3ohVB3fKzo
5vEx57qnNSnjEWBoEiKfAXLgAv6+AWGotxXkE3hgQoBSAlitzfL85RWz6j5rMf0R
NBf4wf0aSCG0sBPQZSiRX0uJzAL1Vfgj2tMxgTt/1kSb0iyUyCk93W2ErkAlDXYH
4smAn/fq7F/DbJ1BulUuOiGKZLyGQ0ZVBjTOzFQtuoy8gJ0/EFN5QffJ5QPIUljh
6RoXzFqvTmVmxoOqokmrUYwNl7g4XsLVdl646DrqQpn27pIRvBHD8fyRuau5ulH9
lSnwrcV//ovrQtn2SWTgU/aHcG9WVGyiRJn9Tx9B52foMOggUXYMjzg08elyxv+J
HpDoBYCicZUmT+itSXv4ddus83O1YKb3VceNhp3c5R2qWNDMDPmBtr9wIKmBAH/S
gX9H10+4OPBpcylq+dgcMios5mvsTJLsZtXkmsU6NwgxcufyW5m6cW/hFRwBnyoN
uoBe4rtFG15QO/MS9OSYgM5PW5unHysRzJfZDKPb/fHg+jMU5Cl7BwPce4TBX6YQ
+w6yfrC6wM/7huiABjaw62zaIXATqdO4OH6njGx+NQ2tzMKX+AfyxyWoqP+devDF
vXWUH4MpKLnx8YKearr1ZT+zoCKmI+dQAHTiX/nNNIU9RXGchSs0SQzdzBzX8LM1
G8LOC6YiMoGS2x6+Chjqr+opDJCnEJSuBF2JhmQaTn8v0ng94wSKaR23ZecYOV7t
57hOFThlKzz/Ex5jBzr6wT7XYzXgQYmZhoeJoP0LXkIcTb8AaWdZAlgut1mh6PZD
Wa1HiId3Pph8XxOB51iZDewhdftJHurcBbxPo3Eh1RX3PJlPLU7pbar5melUQekd
w3u2CzBJH3aN0C7O7tN2gqEGOGd+jZ+PrFwQ3yJoByRVg/no+DyWgqx6tMsosRje
6zuN8DczweNTlNzBK/KqkuU/G9c3OSZrIOqgtOjOqE+Hg/sXbVBkkYLlCnDi+kh0
GnOGNvQMazrR8OP6AKY6fbFrKuA1UDPN3CUAmQoVSxRgMb2lkeKjTXvqvHr45ZB3
4iOLJu7EYlTv1IBkFtin3XaodQ0luFxRd4l7nzHouWWrFImlegiixvZBQucf+RIg
/t5W01R8O2p2hg2ItGbiYmutqS7eaekveUc2FTdwfQarAxjr6WV8pAsVOGlSotSc
5Wsr3UKRnVQpBkQbqLBO+H/C4fzS20nR4TyRX9C2mCHZ+joJ2R+f48jWhH5kJ1p3
K23awdG02Nnd3DbRdny76XG7Dx/ZJ64HxSYcEEjie6hccwZuEniBiWMrwL2FNByV
CywdQ7tM6jr+Of6JrGtPICrmhNzcNdYWr2uIMhZAPAK8lVXM7K728dW8WuV501WC
ZsjoLHwUDYg83ocY9B1BmGX1ivdyEPrLxs2csJ108pAS8NnSqfakzNVFqijS1zRd
g6UdqQqkW8qj8BbvOBUmrRLxUs0cOztZaEYYU12CNt8C04BKHI9bRYain8wMC1go
PdbCuF6H+eDewS2p/ScJ29JEBJtZM2Htl/cUk6P6BZc4CmvcTMsBjAugu2M3Tfp4
hErsVGz18fDMMiNC/29YorW6/Z5esKgDnWnbl3dUSHhYAH3zJl8h+MspSiI40tGc
oxN+YsMYeLlPQm+Jjti16jMiaRzJ2hJvDPZF7VGCm0//KNCYwKKQkmMbHbkh/Xj1
jjRZej6M+Vi6XZswm2iKfFv9sCtWsSaNdzppoQtnZKnxY34neU/igm1waeIdSQOL
8eH0cyBSUByrcM4tP4293rFqjrgNAN/S/F/Bjl0TCbtYX44zUGeenyqRBiquBpjb
Bd6+Vwvyl5LonmhJrDwMjveNW03XyVtV7ZmuHhktkDZpTtBMkIMnsUlEBXuxfSgR
natnxgX1M8ASMHSJuh6PlL4NHAUsguDXihjLpDEM36csZNxVm7U2nwryhx8JQo8v
y/5anp3M/pVKxbPodYEO19gWOx8Sf+ue2e8AelEOxF6HJZ+3AAQ6Pd/wH+dpVTA9
22VmKPHoaGfI1OPUb5IK89ojzoI8wqi3PbNKBoYgECQV7bmMBIxVtqJjAHujWGF0
ztzg9ah7/p8VSRItGf/NpJpFBuMnAuC2D4YrNod7kfbp8mvh0ZZa4YzqV4wvp8Pn
FmAVxpkOgDv/II7bFSx3ugyi+F0bDo9Rt97leioYddzATwuC45C1hXUaQFRjwIwW
E+4+o/RQh7ihm6dDlL1U3mX+huWnTdjD46hFP+nnQTx9AF8ywCCCSasVQbfkiiR/
KOlSA6ovjVvcZF6nMvsjlXAQxPXtmt+DL/IM93vzB5XO7vsjLW+etp1QRFPLs+ex
CkMcd8y7fZ2MArFe2BG3EgOFE5NjAt1HeC4hCq6PniDRo0fkoSM7wwBA0owMdaBZ
Lxeof3B1j5jnBYvB/lvQfq8SxeaCbXeRqj5CMXoJ5GxT2eG8d/Ts/GatHLn/LMSy
C0WzRE2sZbirKr3kk4JhN5ILODZ46Xau4U0okWEfB8F5GLufK6zpD6cywc5otCjY
yzRrPqX9D17l7M5t3vNScEanuMg+BXpgpOTzFa5gmJI/WeIqfmDQjzI8eAPsoPhJ
g03jfRQ2MOgCQ0JRVXf4nd8fi3ySL6QcYwMr6fzpOMdy9RomGmkGo1uUaMOE4SqG
uicmh0LtYlXQFI23ripRrvvbwLQREDtZ8AnzeIRL0y8KRPbcVb9PVbiTMTYH67F+
LhOrX02XTOJO+7TzaMiEtSHJ32H8gLwrdB4GqQPR7KcuDDJHxkyT1rO2QJgcBSVG
x3no0KwVXU3omMNb+KBHKNc12gR94PalEpUeR0NF4srwGcCkeJYZMtWjRVL7fFPM
l4P/n5sbdwmgA9CY/hpAzr3SXa26fk05+i3jNO573ATt/DPUO7OLEIQJxtPcVYzz
tG1l1avhNXqRW15/F/RVUMcGWP42WCybyofiB9vRLcyMMm1RRsvpubDOVsLEm0rV
FPkuTG7iLD84yip7rWqQ39U12tMmNNa+PZXTBtnARwLT3ZFthQWQsyfheeNs4tcY
kh182VInCGhlMlwjOY+MGpdHrGHj3tQD/+YZW2OtXLwUiiQEfkMQOC6h+63IcbDf
WRcbkkIqytfvMTtYcXvf9+NSVpWVHV2WD/j2tb4t2CaBQdaXMyUzfx/bCIeTrCxw
ntTCAtuffgVdnSx+V5HSa+gGcJWoWdlzCiTtTeRLACqj28r/dXBblBGULWYMVyE/
0AGfckvXw+pCiEOhp/3cRwdOO7mowW8/gyXX2IOuB5RtWVobrfRRufPTk0Xz+zxk
1ENn52NY5mlBkuodogRsvjBVQMFX65KmMWCyeBfBGjPbuxcQ7t+LfohgCC3zmptc
WRadbgh0a81Qa9rqGRdHQAjZ7xG0KcUDisXqqzzLlKQv+cv0xNAIjfNvNKjo/qBQ
AywuM+CVvM9jLkg7Ms7/eitXH2pEApNJv4mPPdxSX9aYbo8xE0RQwRo5DOGuoK7f
PpCWvnmOgiABf7AYhn2wuZsSJzKvEQ7h+31SbnLTw33baiM4qq7fbBz2DB+3uDOC
0QhFRkBpQCc4R59zyPWgJpa8PtN0sL92IAESpDbovAmu5JIqui5GfaSRfByX3wNT
jilNKE5Pq+QoQ0NRGNRoKd81TRxV9bY5nhTE+2FY237aUfYX83eh4NIHwZcFLUrZ
Wu8ubIk2LjB39o4IHlB/4rFRTkW6rdRTHhpB+uUQsMd5463dmyp1AGEJhga4L3Ei
XN29QGN1KZ4AzMdOyotfoPWTDRmty4uSOI2b8mhqMXfJccKE0rt6TWDTsu7SX7iq
d1qMcz+wFeqTHTVaxrZtYmJ9Hb/9yp/+2H0EUQ+rpCkTVvu9HLW2rc/BKX6rq5YZ
Y/phca/wKR40xOHvMOVIqexIxI3p2dNJcqEYyiBqxBpVQWuNXM1Y+t3+kG03DE3f
/OJ+ngmXrqntd0i/tfIwuJVAb2XwVQLZ6H/FMndhEmxH+LIdXCRaPN7Q0TbEloIH
+WZdqRLmSHsP9C3G9HBd0sMycB8402jrLllBXHVRexVxJ48vfF3th5CNkcw+PtsL
9O1MPeONvhHw2E+lha/G1f5p4sJykf+G524xApAGFFyqgnrIsAC+SYY32sEIAFqo
9fWsqu5MMYSdXZaO98ZY8H14hEp4/oPu/tvIWgoaAm3iFr7LJq3CPwLLjzmKDPT/
R5aipMHhAvwSwMUzM5BC9MkTaVMDLsESBCOtu7fbiJYNyqI4qFPU1C/yXijTcq4A
8zAJy3dSwU8OoN9KUAwypfUPndg4K4byvsGIJzCV06z/B9xjWTBYzhW+SMMP/lS2
A1blVETTf5GFykZ7nefvz3RSrXAoi1jT3bvqkeEdCfBn+mK0vf5ny6H+w9lEJ0Cc
yr+aqP0u703L1O9PoyBXSi94ndHfPWgnqvTD21+16agkNgHCxahI0b5YqYaZkkx2
4Ut57M034C9uhgjANIbNl01dhcwbsqNWkHYNpmUTQFeIOPSXgZ0D1znPwGftMva8
eUapqkHzC8Lm6n7U4jeBOGMcejaiRJUrK0j02xBeRsiZQuUZhh3nsj6BE7PpgGCY
ebBNGOIcZuzxuPe3Dz9BHcOWK1RL1m39ab7d7ZPbXyGfDpLe5a/lZWmhgZZQjQKx
UChAltmr00EFBHdfqo1Igg4vRF8OJnnCSoor3e8G5Y5xB0/0O9wWdBDVL/6Tm3y5
F7BF1aGQZzTPxD9W6IIHfekQEsEWoOQH9jYOOzIl9mvf4HLj43KkVNi7nxfKBtp2
nnVhWd3QGwpVGXQo+lL7AgWeP4JkuzzfoskJ69tOSfWd9d4MyC7OI7ghCYIdtgIP
rbXgtcXcBMStrFu+K1SLl2T0tOSwPOi0TrpZsN8i1fG3nI6B69rnrmc5/BCpd55l
rnKN4Gkd4maoFAY6sNTghApHXFvZUD0L1F5A/WfUfghvdM9BA0yX7PprdiPAh2US
OxYIue4inOE3KNfYGewPc/Itgl6IjDINJHgLElquarKnDvJO7/ji0QGgGsQaZJlC
tqC6wGXUYhfHgRH97lBCdG7fShosGBAY5fFwnsELJNdeb0r6boYyAKwM7RsSzmGp
Fs00XGMJejz14sGyaV2KngiiaENSl8NBUnUCP06abnbqjqJD4lb+Pp9xMu3ALzLy
O3OKxiMsv63LhB+/BOzdW5h3j4AE9h56nNUzkH53W69IG2oxV0qLjJVftkBvRly8
hamHtkvUXDhvcoYMG7aeuUAzrYqnw2SrzOcF3ShOwaenxU6RkT71IY+iA3mVG/yt
5d+CmCysq5G5pVI2wHOCNNvZgQ/elsr06oV4zMz/t4JdxzcdIehzVf2gEWkE9Q1z
kmLMyk76TwuTZPVF4xh8xUXhROfKkHknYaAF1PHUvCaqQi/+pERHsWaCI7RfqM3T
BrCVw/N7gJcNJf8fz05YeOsZMNZlvfkaTA5rljhAT9dVxPKx+qdLHQ14WTEmWetr
Unk2yuGVnCC8K1iVW8ioPQ0YLyxmAR4/QR34PNC1M2ez/AwHaesazmK/TrcTQjBH
/NF9CyTLst7jc4n02U0+tW7DhLtNxrLrHXUXcPpJXKNYYzjtnR/cyfMAAuzHIg8S
RnCi200LROw7tIqibfEJq6/tcXW6vSc7Ucds337y4Ea6bk57CrGQn6DUbOstItbx
VYXcyQCdMzve7LtSPM2YOAyrt2tJIxhwm1ZsBNtRCOPdohuDwOYXT8yVaiMCPsc4
6uasREA1aY63LeHp1v/aWg8mNXped7nRK5r9g/RHeqVJFuCuZZypy0vGGSVqohpy
qGT1eqNulwl3gX8OAZwII/ydNjcQvBss59wThH4dmtnFk+tds4529LzhSrK8JIaL
ZpV7+ViUL49fNWKNjGlc5YLh6ACe1UCeoTMpYWxybjXoZ2dJ+/eWFuscmaVaRMPA
RaEU3tAVYI0V8uDn21o8vIG/56jF0mXC2sEVrPoNX40Fe2bLJ2MB9/v8mEv7iab7
inXQ1z0HTFIbH9zFF37FksEOpha3lm6lji7HAfE3bj1RSPFw35PbbJ6reP6d/zUd
ls7Shvl+jjo9+d/Gw2yNwN8gKwBbzlxp7F2DhljHE/bbuWdUn052msQJwXOGXaDv
X+7yX9mEDLAI7sx9va+S7diAl0hiuKqcujzoAuP/VIhkmxmcVKLIXt8gyu5+panP
FBZDUci9K70gQT+eF2MZytwNSk2DroAUP5cgAA6LSvIid9IFlgw3+mt0cBtSAK+3
IXI+pCwvTXAN32TBvrQNxXJ7DoHyxzs633xLujKfJZ9SCmYkdCc1uklZuqQT8j0E
Kv/nlECqQOgRbQQE2iwxZeodHoJWkzEHhKrBgiIXiH9B5+mDc75tNRVHEy4Mkge+
6PbTaSJDPhyncFlloe2Q0zliNfTRZxB+mxlxPhP6viwQHeBSwBwNo56nft3mCUt1
0sKpMUpg4NEqxE1qdpYLKLNgLy/Jnkk+4PfD6ld6W52baWYOWNdFN87LKaH7r5LH
qU0b+OYHIxhwyIQ+lsy2UMcOQtGk11ugDTC316NMGL9K9kiU5/33JMUjzv/iEOji
Et9lVQOVsWHp6SgTZC65uEcQ7r483hEFIu1lFSXehJGwZNbijZCJvV5xMWl3YQUx
YAsxVquc3HfIAreTK9AkcswkUILUDiul+Kg6WhUfk4lt07nnsp0tDgCIw5XGQLOo
ZyQKB6uAc+oswmsKQpcicRWsFwyuQuSSGaazG3G3zhJHfrp3Dj8nNrVKKuo6FRAo
XhY3L3sHpLo5k41KhRTLsV3T1EFcUhL+4ewUDmY3NWwVzZTvhMR8HNvf79BNEEp4
R8wBcbNFByNyVQlvkVxmyBtEs9WaE9rFoa832DiKG3pgV1JrslOhoJyql5rD5MK0
6dWbh1MB3AaR4oaHVfPsiydVZ/7LnWDpMLpi/QVgISbIe1KghHUh8kAPpOkng/43
1QK3/0RFk3lZIFvp6UGZaJMRpOVMuv/2LJMrOMzW/qn8xwb/Yw0f5veRousK+OVl
tH6sIQn7Q/hDR91dIR7wSt7XAizDRJcqAOAmfSiFB82rsvHYa/SBxPP4+csYmbm+
2fa+tNo6Yym4LjPsBFCCtP8th99MuAvVTiqPdXK3YjY7WsZECOXYtklD2Tw1H7fc
kGbxFStLBx3oNuEkIv8PJL0qN8GK+UbXyviNeTc1rk5Rdazh2+P3LdaKsrV8Tv5d
YSfhMzISQRbp+JOrmG+6qxRG9t07xGaDr0njpKGNbOZvvHWiUBY2T6mX8yG/xp8Y
39fkbpZ0iNXQzycH4X9qMOxSsocd1L0QJs8Zff62I1RDT51pnh2mQuHeop5GPWlf
uuEdEaokKLQTsZ8SsgYdqx8XISyv8JH7MhvzCWj8QtC4lIEGV5iS5p4q47G5KZLz
V+AjA+BnEB1rw8xAIRq2buhMW9DlyQLJJWtvxsb7JBjLSgC7rhk0qkgIZNLkjEBL
gGYDhn2pO+I3Xv5rpUViqmMxsso1+YYacCLEFx9duSYpCwV+MofZqypHsKkqidpC
JGE3LqUIJ8DKYocMBNouFRvNVFmwzXhIDa94II2MHaGq/Oyca4xwYB+x4+4fpw/N
O865A7puE6hwDuUN7VizS15POv2vX+Mf0ujsWGKioUCN9TdaFXofl4b4QAJgfXJr
4uVdkAI78ATLbZ+vM5gO+ULfo6dkS3FSpKVKOZlGFK8wUQg089AcetmcYZdxGBak
rMwCM9f3myYYWEX1hmeMNNicIKizCzfO0XWHkhHE3Tm1JiKmsMqPZ8o+DmjiKo0I
b03+4jhzype2dwqbc6Rw9xRPFj4XyOqv6mqv7pE0Keau+jKl84J/AVBt3ZAVxEQY
fHz8/MwB1NYlF2KJSWdKoiqDA1GG9SfqLsaPuV/iEtqyoioOFyIMoFqN61U+TC1F
l4LrUkssN2eBd0iJ4qQw43i9SG+Pbs0s9AzbuE82zveMk8hLARPQMTtQjws7S922
TbABuwuhpAcall7r5Dh2DUVA6rcsc+e8Dj7ABCDG0KFlnvr2qdsG7WoIp6QSMUqD
TIXu0vQKjNaEUlPrzyuljqIDvZEvxxBj8oHvKmA3b+UqS9dweAOETG5BmSu4B0Pv
PGQQFviWzP1NZwg16QBLjkpCa1jmG76+PRg0VhD3KYydCcfNkNgQ1aKOkw//ToHP
N2uIEa354SyUOX1aIxyL1J1dEDy37pm+VnB4XbmtUMRMzVnO35h0xwyY9sG4/It4
tId7zDPUicI7iO04GXquBKsGILZm/v31L0G4jPRl0aF7jQb5mw12NDNDcnxQwhEa
ANiqGUs78OlRZ1Wlp3G/HWiczhiAD0KkxDolF7YtyteLO0JfDxvKqxd3F204cm+u
fiW902yY/ZW9cCnNSk2Fg9n5jMMNtqV71orvOFz0R0hnyij6C0tx2JKUzih8o6D6
JiaYABitgUjRgSALwPUXI2Qmdo9KXpXUBtLWmnamss7TrCME30/A5+2Nh9Sb6udq
kxuggON2PJbfE+vmVqObGOq1uiu/bMZY/A95zlyF1C//QivQ7RY22/LqfQA/rHj8
4hIUBBkLHOIbqtsLundYBLNlh1ZryscfMHXs/oSgAQ1xRNpNl2aG6N57m1ewqVwP
f+KKrKqtF0T67NARLH8biLA1wg/93run9K9JLg2TmQL21iEIlOL/Y3f+6ZdUUv6W
kDHctNRRAeAqh/7aKfdt2w5NM3NXzpHt3id0A6RPuvYYvqfWYlEpOQe5uvqW8ofN
s5FKjmZM5aB6AOSMLdkwcln52YHU4viHec4um1S1FEsZAB2TeTbhi19ahB+3UOIs
x8bYR2tj9o6ELNpGRs1QFIRXzSrETITkbfQoOAbN4e8DwLhYuxjNpKopWYrfH2mS
3Nvxhcf1vJNcvNd9EA/VQ/V7AEObZe427hT5auvvKdD4Qq9ylfSbjourJljA+6BL
2u/UBoct//LHSW2wH56RB0yMI5gAj1SY5GVr8AmHtBgjOfokiIEFjmItaZbia+0d
JyQ49cGoOZ8iOYpX4j3Aw02OaE8h8X2A2DN1eDnBodDDOKLxHjXJRSfClxeq26RY
sysQlBwOOn4kJWCQdj5i+OzfGQxHqETpsf6kRTi3x4s7uK6STjUFTUOQ4ksvS/7I
t9pmaHPlPwm3k2OTCoa84p/GfS0a+RWzCUS30vvgouw+YGUXz/sorfmJUNaanExh
j1TziIDtzoh2m7aUUKfkkroFHGEQ8CxqfvrIlmgZmSluOGbjiRj7O3Wb2MePJaLQ
pkMr7yWnk01+XY2ra0vrx2ZNMylFQMdE5O57GlpC0cdUxXcSXO+vOWtLnm8HqWUH
zUxq2EBzxoNeeytesLLcfMVsJX/rdq6F4ATBOYWyVClM8AyoMDqMs6gar5vyFjqs
MVXowq+CkMLpeAzpjKlVQftukXc6paV/oldFXOxsjHP/58szFVp1iFfjTJ9w8yjK
RZpj3+p4eWisQXPMB6YU5ktuQ+DUqoB7cdF4F43gq4CwMd5hY8+CPgsTqWV4XfLL
w0xyREjo5T1S4hY/fFnuOCwmYaMRDmBXDGJcaaFStaAaGctzEz3A0TPS8pgYjCV/
Eyb+uchC+iMUmePxKNNg8yUvB6kmkbIcnaZsW8P/Zr63lY6CxCbTxtlFWSS9m7vt
jLIYDhs16UKahpsnN+LFSxwncdBEorCZ7EKQsGJlXxoZHzHbOrLWNrXkzTnYOymr
ho35tyiKoniB5G+oTtCB5omLdwM0M/NKj6OTDEaFEi2BJ7sNsh6Iiu7BxVlqY4eV
qtjWz8hAW/VsLqVEwviLoJKFLtngjTL0C/8DeEMgno+hm7mdJSDIGcDozLaSfDKp
teUn1OCwJA9Byg4EXvFw3Oz8httGD9XIyo0gMYteWrBHjzq72Ov8bG0b0qIVc51s
+V3zJRLLGvug+v59aV2c00sNoFGjvcfJr1VqgxId5Qa24n9F8pNtdiq/99inYpn6
HhFrt0jWZLxTc+Pd2SYGr8ARo0UXGrIlbpV+kcF252VHPVvROMoTRtvGz0xjL9ow
OEUa/sF4nnXrRkWdMrZbd1fTWMEodq9JeKX/RTOrbEcf8PwbAjusrGghLG4DaU7s
pQ7ht/bUoUPk9vcATWGLKflGNFne0GREDWaMO8URMs5t2avUf0EbgZJPygVpxDom
pWCAC4ShO1BFVUIuWhliaSbKpzaX6mSj9LXzO52C7ibN7Jq2lLC2UC7okb1N2KfE
y23wV7T/+52SJ/NBUhf/rpqGKT9FA4lKPxHNwjRvKGfuGmjO5JXE1s3jVq+yEe3i
J66KB6GVxt9kVTBS2UCq68xDZYr0VeWLf3QzRO3lRhIESNcz2cZ4xK7pDd6De1a3
0K9yCu18bQ8DNx3mExIjvnXcfgaFJK1y72qgMr98cuxJ/rbf4765Z8YOX8LNaPbD
kXH3egJndXvFz5JqVz9NuKSqEfq+PJj4iR3co3iqzTrm8KbhPOg0EWWm9+Tx03VQ
LNKTEwWQrrbrshMLrxY5Ybw9B/dKyJBjeCpgwB3ncrkpavT58IwOflMPWhXEVmNI
oVoHV3j3sMFYg08rrF8PrS7uBVz50LYWHllbSPjlXyQmor+Knhn+0PqzJ4CyK91Q
mI2eiLEK+NKkiZGt/Ux+OTWKWx3n6tjiOzsifeURKNNBurNksRQ/uTqJvkfjwSs5
mjxR0tnDEYB74LdDKiPo+ExzhJx5d2avZqB3h3sxLHgUHIqh/L2KHVj1HOd6nNRQ
9O/2cA/32Ton1wJXlqoeOVpL+0MeKgrPzJZD/qunCEchpt7OlGkdmRlnh7czuIyg
ymjozasC6MC1NoDQD8vAzRkPLqEyW0KL9IsYs/i1WoXJLhPrD5GpqygkFhKYJ718
IvEdCTwurVAiU9L9KcU+t9ltp1rsRLqstfR+1YIhK1Xr+qJBloY7SwazO8w5+GiQ
pAQWEBX69Dl+5LwBBpDUGZ2QYS3UCc9N3F7EE0nlQkNr76n9cgqoffBO+JWwGpee
67cWB8aDzJYUv3KwN48kvrPGq2GggOJq0JUt6vXy/ETdREZHYnlDREDtSCBK7BFs
5djh3PnYGUWJ7U8owJV4uBi4rc8EDiLxxJNNadC7Val7KkOgO6PC5Ml2QmyzVHmm
UYnHNGT5x8wyxiFegTsYEzTSdtd4xJ3cn4cbFuy3HkX2t21iKy0VldxqXWD8yzOy
X+PdC4Cp1GCH6NT3c4BoFafaJd+Vk8BFFivHuMiDoZP6bpobobsdSV3ss645Dc71
DZO2xtLb5032yhafEvudmqnPvXjFmIAj2+2TZUgZS6lS/r3XZRAi02pQDiiSMMhj
Dq6EXNpjpdbGD4vr4wQ0HVfrzlrv8HZFt0Q/V9Vj38IQiIGA01ESSnAYfwpnWCIT
lQWXuSexYEbHffICb7cRTvKqPBFADFsUpmCj3gBzIw0UjOjc0ebXURON6ToiAgfo
SZio024rGWg0M6IGmkH6+UcfryxmyzaL4PcSy143j0vOwnAriRmAnZIJbPVcMUKC
6qfHjUKZIzb3cee4/mwipZMHtcWu8RDaBA+htxZRISD2in24iqNSDuyKCUdv0QPd
TKsKti1A9SRXlnsX/PeCNs0tRAUaR/TPkIo4qIwVjWKzLaDbkITo130SFtq/GG3V
OnqgZNHCLRXx4HqizzeLEz3FTd1S054CKh6Ra7cby3dCYuefYfV1lSQKCUOLZ3rO
5HtmBSFcyXEzfAQpbDJfNN8gB8Flc9byiq1+fStHwRKXTZqLjqr8/6iW7XnuZ9dP
UWXJ/MH+6Rs4jPJGV/vERcFJbXMTuBWC8UJNkOAifsn4Y54HP5DA2IVBgte4JTpx
A1sPnxvOidRkKSyKcBmvG2l65DKPoc3Lw2sA1D9bMY8iGtdw0XoVFiO5Ay7+f56/
spp3S8NeZhDPWHsUnhyQ1tjGjgLJRQ+RDHl6/FuDwVgNPhf95J5bMou2yeDBP215
ovM6GjVTaJidNRy7RJqZQ08wBdaR+YMOvMBaFoBcpi9QlPotHehtdGYLX6wePyHF
B6sV/t/mJGsODC9DxiWTupUoWRk0hVpc491PpEsbjI55JLRqEBvEFGzJJ3H2rklu
ss2HNVwlXlzOvH0vKg9U7rDcN79YwuUcUao4t71A35R8XCfMzAUmj2dfwuB0t4hq
wHryOINwPVe0z+IMW19lpQM3hMjQ5J2lxVWRI3sCkXoK7xNi8ZCYHp9gz2iE1Na2
JNltMEv12yara/FmcAkht0hRId6bYUrB1evIDHRsM6jPi8+5wRWMTqKzacbrN+JM
l6TwTCvHo4lQRI2Z3vtMm/LSKs21Pupsds7+vGNFroyrLawIg4MqYzXN8A4o8lWe
lA5ydRAKMBUzJkhKehbIvNVPRyWqrjPW6WfY6TPBZY7i3rezbg1ilp0VuhkXsazr
vzlwDp8Ef6XnipJwfUdTMRK3iOzVnQyvC3cUROLr6PepkyPerJOPV5HITHNi/+Vr
XRnCrxWxrw/bTE518z59PskW8bpJWi6d1X60uxn9vwidZYtFfodaAyepKF1hs18p
aTYZuDyvyKsKj1kgStCkgLm2eyVy8HsH3zQ9pW4JQSZB1y3U2Bn/VyNpmchAaUxK
OYvm3HXB+/rAcDprCfTRQm5LSBSw5QRkVZ7g0645OO0xqvrMol6bJ6D8CMy5o57W
j+OfvfOn8UwiL89WfkdGNocAvs3m91u2FdaB5qBj8B0/VLVyERYcvkE6KzbmoV5x
G1jBULkZJxjlP6jJ9GfieFYfNbC2lEef3PaL+/t0t1pdeWp3a8RojnbeGiRMbr38
WlxuDzEhLob1O2/EUyd3zZ9e5AB2gVB6FC6ISgEQfCoAG7Jhm26+XukjRrvt1yri
NQwECF76jIu2lgnLUvQPTFgVU59V00Ibx0TLGCQK2IrbUpmIwAChsa9caymg5H78
uCo+o6pnI/IzZrKFErWV/gLJ6fw2cR5j7+eVCZ+YqjsHqWTg2WALgk2Mad7P8VDa
ZOibUVshzb6mOpJX2uZJKZqilTfNdHpkzLCCtpjZELc5B50ZBQUv9ttCAIdULA4c
IRBI0k2blpqSvbwYXBxQA7bTPnxf+ATVBzZMs8qhguGs2rdoYVE1XrHstcpz8C3H
5J3VNr81lmyWh3Z3pnIivtAKBiiZov9iwncEFqGIVUO962lZkClRd5CixyiHN7Cs
YwZJEBqa8vkHvDrYlc4tMyZhr85p00sxg6/ucevuDZPGA9Gpwu8qd2wVc8cuO2GA
1bDQ2OeM+hCMgQfFZjwvT7NolHQJLbfkriUgcWW8gsnopRaCCWB3EdAissX9ZHNc
79DkfeBU1zSvXIV/GJQtO4Ofzaxh1ykt3h9tyjEcF2kQI3F7h/E5D0RmSJaf+XFs
8wFy/KDOf8f+dg2iV/IhIpA7FuwiG608r9jOFJraZC+COPXmTT/kvl787bAvHK0S
fKVj9Ym1NH5n7A9ymVZNMoxwvUiBVxP6hdewfuQidxqMHz9Y/lywauYZm18r5KCg
EZNMp9StyvzvvuFwluMlB0Fg8m63UrHXg/E7tXu9Bgd6DuaUTTCR9FQyar3ztYHC
rLEvPN9J+4tl8lhGybGEEG09KCHlnQObVHLGgCDCupdJky4XXz+qvsb3Lh6diFKH
lw1iWAWRC7R75UAce77GvMaUNkr2QzGyzFt3MSYZyPYWGdb0AfO1CEFEOC2wEl+q
rBGVMvIaPjTKUC0AylGRCdHIo5rru+FYOqhzVLvwmqnzKmIs60CgyaXBbqWVqFF/
v1k3FrhLtliwLUH42s3wJVHKmar8nGrDKqVB1590/TDbJQXkLbHtg0vXx+A3n4nD
gSWBo/GDCO2KUEvd3p+jsup4HPoDed22RBDWTlmtcneKWKXPxzn8sm7wecar486e
nY/iNU+y/H09BleveSh4/4Lo1iCk1noo0nf56QJ1/hQJFStdM6aEh+Hc7EytnTTG
WFi2WuOQM/K4X6RA9NrctfnmwGe2vQitK0GDgyAUGqSh6oQUxJ3z7p55vq9FxuL8
Kec50UxZaxPYt6GiE0URUjuGULvF4KXNdBOA/aglp1bFlxDWc03J5tP2VXAbheCs
/GI/09qNVr3zdkseAPg1Kv7CiY06c+fjX22CGDe2fLYvHYyQZ7b301CL5ZYX2Vum
OmQOhxkxcA61uTZiveQsZfG1Dx3sf0BN/6MK1t/sEXYP0Wf/YRvGhOdQwvDf0DHp
Wow4oYvGQN33IHKbn+4uSo44T64TDVaPceiPXkh3F158Hu2nWDxSSORPB/XZgOJ/
8yJvrMFIsKVul3izpOe2ysleISR38rTG9JrCyWse2nCN03bkHEFoNFRHbgpqvMDK
ectCS/3gJDC8aVOK/AFgqt4843aBBYC4Npmda2iFeiIarrdAKYdryTqVwq+w84Ol
RSOSzy7pzz0ftpeDc0Mt9vkpU0HknSRKhQpfzaJI+/5ImBkNtTxBgcA8UOEOwaS8
T1WI+NMZ8ke8erwz5siJexP91+Ci1f/Y6tOMIU4HzVjaY/jh80lTQA/alGp+OymF
TojvmxEVDy1H9Aobxnh1c98telEe2gRtrMglb30Q8viKT32vwg2srvu4eXLafxP7
3CUWFaSsjUrv+V7PdQhaaTaUMaaPYp3JAbsfzwCB2GYHFkKtorLH864btCXVmzje
NM1r7lWNc/GGo/5vAGUcDGMorOvIUcq/KejNy3HoDnLYUGdDblcVBhbHBm9f70r2
vHJGR326xlmSpmhK3rx1d0UM/zDmvaijUVJL+VU/mk4xbPz+3mGp19HpSY1ogPwH
ImZ2d5SLOV/KUyAxoCgwTITchaw7gMbxp8HiEVIVpKs3wW3SRn7ESebprJEmYHkp
qanRf09ouc0iR5Cly2GWWvIgXG+AfhFXnSuYeYRe7i+ib9wRWbY5kCq94f6DTtEC
7cNfzPzoBTH3scT5GoGahpSbr1Ftf1mYnTl5JprwWEsfejc/6Y1P2QvriEwfMt5P
uE7/soX2Wm79gE4AFzXo2GneayCpZODlYE1S13JIQldGRk9Djm7GFs7CaqAFJM/o
n5i+L8FhM06ZQeFrDJD9rKcOvHJriNByW7NcdKArsxI7I3wuJDTznlr38g6BFbc5
rt+wnrwU/HLSS8o5A5IasJbjqFTZPiUTC9wmZk+fJ+YxmFMwCep3uq9dDEsQidZT
5s3lv/yDDcSRlXIvEt+rsBgBOs03/agOenX8JGzcu57wjYow2Ga8ekZzN9eWEqrx
MTxjnA4DHmODEXmhKd5L3ZIyItu9uCCl1wtn+roP15PZuNZL/seWrOBCd+OwcdEM
LDzye9Np/WDcCGMjTNIuHnGrKn1xW9lkLD6A5aHtF3JLcuxHHa7CeYa8IvR5U24e
7D5Cu8Viee5m66orGp7OIYLF7w0vS8JGBzWL7aKJWqsqpXNg+PH5Ee/g4/eRED2x
FKqQ9RyW73wDUyK0LOkEopKRa/oF4qVK++y0aABows3Vmde2W4y7UwZOsAGbvLw+
Ze999H2enmUYRuwvYYgAEJnjtdJGz9lNoXZJIf4YHBSK9hswZYvkLHpqDODlEWMc
NC3o1mQQlw/BVqmBBf5Ae0kayUsYMxkbksmaDVXAz4uoZdrCQRLwmp5PKw955x7M
9WwvUfodn38LYE/2tAQSLZUn0AB4jjkre8BtMe5H956uLvmgrKYXoUwrxJ2TjAVA
DXAR6b8CVFizcyTViqib22MCTP4qWK4bWX4zpFxegS37hPjzQajPV6do1vzGwNCf
zpf4oqsv23yCKJ4Yw8LB9/rajPSEy5ZT3b+PM+jWZtDoFbAICEwIj34iyM5LH7la
ka8L9N66Ucxb8qn+IcUzEoJ+Fl04RcaqqwD3RtsnbMrc0uF8OlXSgENEP2HoSyjx
H8j3Meh+Mp+9JSnrysrYbeSrcebHMKlBN34LEhnsZHrIA4qzE/AVPKbgZ85Kirjp
VRVW764ZwF2y45qadkybSL2oUQi+hHoS+D9xoLOjQqgK0CVH6674RKGAOK9F8wQo
uT4MmXNDtYvMMgU2TW5r4dvJ8syMkFK/H4UGURVbvTSIbU/DJth5KvZaUWeQ/ZCT
eHc5AQhhmHfOIbuozAmgeaqKthEwR9kcgUVJXlbvJU9yj8Jfj+8kl5J9B47ZYlGQ
HMRnm5wbh5+2besowad43lSfs+WjpfUkHsWKvW6XHPtEQL2f0HfugFpm/UhsG0Tx
UIB/lpBsqUeMkAJwYvMI+ocL9g6uK+wi+xhE3+goGFDA3IUvE9F70Q9vj6WDzv0P
+BG2DzkJX/StqJQ1UXN5B+bPUBi9ix15yf6gev5yy5nf1O963unutn0aSCIdOjvL
tj5sQQ8ny0YUTj8ezisOqTUQ+nyTWwcUrwPOUEujOoL2b9y1H1KF4xYlqq14x/ib
5ITRpy8HcZAOalXG6LZYLAxBYYRG/qU6PAoESOWEGZASdlLxmokXlbd9pT4rZtKi
eKfKDxlWr00c69sJcL3IICVfTJqyGPAkRHHmjsWmq7O5Pfs+F1KkV9y5yifRT4gE
D8OHD8jkWqyyweeBV/zPfLK9FXsZ2H+tgiLbTZoqBSoSbliwBHVy6gbYSWCW8nkb
qw9ceAXOfcD6byGpaYQdd8Ww/cq3LkrD/7htxWVc3sBVjXoRU+oMZjx+GjwEJ+AA
kT5GqFquoGMV4HqN5FjXnrdgG/hlPFIkS8kZiTPgIoQiJw2Dhf/BPeRtXpZ5FGPs
L/CycwWACc+vepR5dPCZ4fPkCDaaRZygGuc8KwNwxVkgumyZm7QqWNQE7nXvTlIe
i6rO3eBGhAKpQ3FXDZPANnWcgLvSGQ7af95OWGfRNLWWbTo/KfxY8+f5qlt4VABd
UL4jogkUQZVX0SsXHIfwpii0A+OJKLxaOIe2V1cWqDw1CthfUHszVyhZMcnlifOu
kWakaZa6PTG3RhLyCqXA8QwgrmcpOdW024xpO7bnbjKksuH8U+qabiHr2QMafkQt
0O4WB1yF4VNRCGpMgrF6xR6a+J1EM+OAQSoOPTblb/gc9ZhwabiZSZX9vS03SGg2
x0NksPaYg4BKB8aLxN4dBQwYrOdwWh7b0hctBeZbNz6vBvf7qqWyUDMfOeSWVL3u
ejwfblzC0Kj2tfqCkA0y8CrtOypcm2Ob9qa+NUi1MFlg8Hfq9rnCmmtjUuxld1CE
hd43YVmzUILXeq6V/NU8vMdxAOTLvhIH0EIt0jV9zvpilzDi7DcOAEJr5P1vvmb9
0DOeO5Z19TSrbHqrfJwFJ7w1RrcSQM2yAroYuYQ2hiJV+DaIopIJ/EE4zwk1NVOX
uMVWNKmMlARszDJXm6rQfml6vVZTO0R/ZXs6NZuKdcOYmrP4V+aOTNbAYGRkMvUB
YMqYINVRfy2ylqDUloJmHbdzq0sQUY14TacryeCbtOBWJ2nKU0GASVNkXzta8hR8
Bo3g/2G7Q6ms5lNHcdtdI4lGr3bNQd1U7N97Ol3vSjYqiuBVCMAzZMGUTtuX3ziF
mhoqWN549YBy0MNUycZDeKu1awbsU1yXEFdyN0FHMNrB3XFBZwitRcc330z/vyd7
CuBcIDBujUgBUvxgbVBKRLhrAO2Xek8AX0gWwmr1tMvKClnyyO2nIuM1Ym3EPvEm
LMLM6T5qDZZ4hLvY4/YazLsa/OK7fD41iBR8w2q4B/2aSakVFkuEq5NdcUgY3X1r
OYsKt2Vv3E455u9FNgU/avPfsZu1DilIU1bqQ2N7ff4CtZA+YVsr2w9sKNwzSTAi
kIvvrVTr3lbqewl5jC/9wcKUv2umbr/zztIJcn5dCazU4vrGa14souzVQ6G8zi/S
baabVHT1viYQ+EBNf9cdQD3UExY7UlOiCPO34Yslw5zTslTiaXrfsiF/QZnNdKki
2Ryhw/Iz1iI8gqxVL2ub54MnZN2Hb4heR+8yf4QoBkubPrtiIcFWVR6Xd+BddMWZ
sVFGSmO3ygPiSCE5WMliKxzLm3LKx1efqrzccr9HEW3H16O1Or2kgDD7lphzx2sy
uysFjkczhsuIV6IAhy4vAL9SDcgWiGsXas7A4lYF/Wuu59UBtN2I6fQNvUIcwxuh
utosr7387dfZbXsBRQY84YAVSsvUv3swKUY+lNnEYQHoCDbouIb0qSH5Lnz7yx+N
CkimubrI/L4o0k1fHaCVA5qvG0m61KblsbLo3I1yt+LHP1rArgJJbtAeeR8R9/fN
eRuK/bq5Uz5UJwOGIFxHqnyeY8j3zutP0PJ/LwJPpKpdCBQLnWqMrScwP/qJECdy
2EBqZ0d62DmEll6GjMrIZ9T9fu9jMay6ycuTiU5Ltm0VIgN/COxKVv5rIZOFRRAN
1xFevVnM1AT8ExCu/o1daE3qNSQWeYtZ07Spj92APkMs/9MVCVjfCd4f4sK+gAXH
LEeqj9mZfrfqz4nwwoGpAqfVw7ahNPvfCdBEr9xCQqiVnQdBpy/g/BXhvV4SF71V
uut21Ls6Ya2f4kPyRkv0/Rp0OC+GRtOv9wWvzJWnrrIBuxyk5Vj8KUoMHH+ZBi5F
DOl7aA78G0oif4x4/vdCrju1VnauFr7dvPJ90LF/Vdg12O62waL0nRtFj2uqjyMY
iFGDNX669oZlYiJHzqOgO41rRguBpfrpkn97FzWI9x+CO2io4rdTIWrFDscA3y/a
dse5+hegQjwyXlYn9xaRwqgwGV6LyDb7c458L3FjPEatGDEMckKZnhwlNC2aPNch
YJ4FjtHOJvXXK6vivBpjRN66ssNoopBU3AEJ+4wPYcpXojnO1w0n0Gey4kNiHLIh
e4frEcnu+9w7KkLmZp2X0MygAQ9zp7KsV4xSY+Xf2sIt4sHeMQEkNlMOtP35DzjD
+5etzBwvJuPC5Jm22+QOzf7LDUVDIieXS9Innxsp1ZEUKgkmx989lcpd7aexRaEV
l0jDa4Ca9UPB8dPpX2IIhBhx/KWcyVgOk1r/KM+BjJqYDQli1UZ/AaDw/4CbueLr
Awag6eX/qEqeYMWZpeTPKPadaqrjsWmv09bmgCFRjk69WFN9S5Ej8RkP+7nmAgUD
q/A+r+fRuKYAR+Edf4jikecebqVovWaWmkXJhDHuKoruMcGxKL5fPH3P144j2/+u
ZxraomGaNog8bwfhzd+Tc+/HdfVSuD/gCJlo3C/+ChYrOSUc5HSQnXiioYfjnOFt
SX5tjwtL29/WIhunT6pNZHwlvSbdos/6bE0O4TazXKoFCdLlxKOc7YQe0SPBS2JY
bkxsoZZYprY+tKYSPf8X9AZxGJypQd0rgOxRFHYo+EmURH80rZFrb2qKgQKUafIF
DIzWowGShpCBAQvZLacwwmovuuG0kDsCccRW0o9DRm45H4JkzlcxRz8uhdxXYFee
wFKv0f7by572g58E6ZVnfI1VphYaNzber6qvqEibJhiBPr+4UppaxP04EuiZDXfs
a6DN+KmX8cWrE1NZ1puwmYgHjuz/kaLQjSsKiYHpFlPAcaBS4u52KXiDalCrMiDG
F0/kelhCE36itL/JjLE4THlMM1tMvxMpfq4EbQ2AC8Pdm8FwgJ8WWi6BZMaIi5E7
Rfk+6WDUTLCevh1j+VJUxRiXm+EB9vYyZxipR/qFRSVNia+/H6w72slqMYvh30ga
1VMUeX2Wmu411aOFjbO+35AesbFeB2/n6tCE+ieKT6MI5iTC8IGRf8fSSkzHcu96
oRd7acRjVn8So4QIOwntsmZn/mzn7EsmGj4u+oGw2ta/3PiadUGW6Qas3gybTjSm
Xul2DzI9LIlzEOuD56hdXgyuvjldHJYUA4PNtdAyZF0o4iVh2l/bhbo3tp011ag5
llY4BIybTTeDTVgaGZN2J0ucEeNpNFqCQ3BOKQwHLFhlerJR0pPge+AScUyVVpjL
qLR69Ks48hyIkpCtrcjfQoNOMhBR0tsUAn4mHgv+guBdX21h1u6l1jvPeduIdyrF
r5DvqYLgweKtQwtNzH6ynoKQOgQAyIqI5vVQ+OcP+pyRS1Xb6wYSmXdkjYNz794y
9veM7LpfDmEvTNVsQ2SOS9P1TG2ukREgUQPSuoPZwPTZ+iZGNiT5eJpGIj/dC/gJ
HFaLFFIsKNwFfjB3evaoQCLAoEE08GXdE10BOVbrshxcKWDqDapaEjU7vQvM7x2d
HoQqkVTY5ffN/ko2SK+sE//M9EmYnW9smJKgwQUYt1aQZGX6C7NTwhbpJQLzCW5x
4yrIpFv8UBW0Fmvb2QvLhEJxUd4fe6SnNpzCcc10Seq6J+ClYXi7yZEgggcK0MoC
yf48BFB4rQUSdXAl8AQGMpvm21rhabWD1p27kpR0VfGjJiW1Hls6TM0cc8inkzLw
+Fi2gJSIUBNcVy+QEcb61YWclv0PWN9KsrxcOjWjZTPV8qua7r28rxXzcpbnXh2h
EMecGgBHjfOFVJBwDmvVqpdO/PdeLQ8fVivY59gTIWQhSkiynCBVYbcTVVLIOoJo
mKi130LPls8SKAbjAhRYfpenoe+XpHlFpqfN5qlc9yM94N3OlXh4b2L+swJyzHJs
GNzxeTsx/IS0MlUe7NKUYhh5ItlGSOKycFLYQy515OoHWfm507sWbC0sFiQRJ/ms
473jRx/kfXh2vVaGE9PuAYlAWXDpt1Q60v9UteGX/StdkLDsdWq0dJg91H89o8rP
++Toys07Rn1zPbn6WIg9UyiPZsSKgTjV+IOraxPnf4ZWW7v/jOfm66jPlHzdZJi5
ajDOwAEaGUifBKy6KB0+rMOx8Z/dpZiMLlX6OoXcBO1bLEaIOlZR2gwCLZ9f0rbB
w3dpdNREHTIFPY++eToFt10hNbpvrLdN3l9w9XrtU9TiVuVx92zKpVo4XTWT8bq+
6lS3SS/jz//OPLzsIgcp04C+r5myEU99yNu+uM6d9bqLXzUHc+7eo8P2dnH3p8R/
Hb20ErksgNKHLwcI/07pBISTqfMFT+VqNuBHL0Xltn5y5GK2OUj4xF58vZTWk8cJ
deoNC+Jtp2ppbisPZ300ga9MygSRVuB7tUkKLAWgJ5lBZPVi4c3xoHWG7OIJad2T
d9EX/vH/nNG/JFu6/H51SSvzzyvBMwHGQGIQvt7WZGKCiX5vtiyyPB4+3MvP72Gb
whcPijSoZ1PxixwV4yVLj/K1QG7Pf5nF7CDNVc3etbsRaCJgtV02KI0bze85wlgl
wZibMnhC7FyD/eFxJL84Zixw+IBJFWXl4EjsaHsot9c6q8UqVPsTAdUY7r/Gf/rs
6LPQZdMhgVvq54pfQjF/UHQ2d5Mcmyogynh7rligLhFL7KCBhRHr2/z5d11ZAcI3
bJ6nZ8SDsfpUARwWCtLwGkCQKO536uvxAR8y4daRNiK9ZPUvCnLNekjNNMOnbTRp
T5MaLY6dlk7zmmTYBY0BCOgEJG2jC12V+dWmwW4KRm/oU1IvaXpnnsiCVe+en7uq
GIp0QnWak4ZIx/sFvZw+F+oyp8UnfGjx/3jwOqF0ulLMu8SFDm9745vnDwVPhZxx
wsrbe+qi2cOw6wdat8G3HfBCyjbLhts5SgMUU3aX3YqZSsYEPDWRayZUTInhgPpp
1HhBUf3M0FasPapbpO+HPdDObUvK4YqnMULOL/byUxHVn3EIZhwJ1LOIwZfTpbE5
TbpxjqEFAGlmMnfmwSzGXQ+FHtPjAKF6qN1UwfRDrFE09ZYkhFecNs3xVfzPUmEV
ZkooYUKozX+WfVziHA+PDIFwhbvuWtaeOHu1EOp/ypXWi48O8IkEPU6B0TA/5H3U
Us+1uv/c1auX+ZPCrNZpfkTsHqlhcHw53TqJozjFW//P8QyJpas4g7hk6NENfaJY
xZKmAXph+zwMO3giwPBaL4z1O1cgqjdTI8oFiRBpHJYZZJ3QooP2qNZFXgUTKRXb
Q+wZHureaAv/6VXDJL52wJ5EbCWm/94/nhVKQO9NGPGl7ewPf7EbEhMSyRQHosoa
n4Ghc63cD3cztlvC/TN8sQzT2Pl6fwEcqZuQz7gvQlZz6CxT2pWCS4iNFFHuEtVN
IqME/FEpm2BDuhnBOktd8vm+4TM74tgTdoNhDOvlzzvsETA7QyozD89dwDAJISR/
jpx2l6lB/QR8Cfs4Z9PbwERF2yBdFGkJOz5gdkcrDilLNNQ/WRxUjDWAvN046A5j
r+KjX9i8JuIAWVOnyft3Uwj5SUL/EBG9NwmVnAh5/ULKVXWk4h9auJpvhkmQbxOA
nIbVs9CEfkaQdArLAnpfNKKepCuCUusLGwuTWJKd7O+dTexHloENTlOgRJoMlpkU
Vl0p/P2epwGsMNxrCqBPPOdzxymSRYMW4uUdMP6+bgKtjHY1ryXS3lsaRABEJzLQ
w9qplEauT0iD4QrOqNFm97Dh/hcP1beKR633qgjvxZJtk+ci9bZH9piZutBgcolX
BpUfb6aynC9/WUzPnqE8uLHgRMftnIKYJlS2Qgsfx3B3TQI7wDv36FnbehnHLQ+9
5lUlQK4+eiTAd766pK+K6ZAFo8G2AyvBV2lg2iw2OKL35lCMh8Y0jH9HbQNvRTsk
x4JtQ5TzexOR/0gA8ITBdHPSt3lOsklTyr0PwK+9FXpQ+qlQ9XTTJdD5zbIaRgME
2FuTbCoBwHf5JQ8/H8ExPzrFT8GBzD5vjk2YpzMSqgLLIYiLFS0g7bjvtu4xf7G9
PXLQvf0uLbfC685yE7mo3fc5VIh8hA1RKWuUESL9GWf5vrjvbnfS3polAJqfTqGC
5LZSdkHMaCpdRtUA8Ad05zGtwcP+Gi6GPELvncTrgDIeoYh8Kx86o9xMJv5CMxVb
MUvJvQOiaDqJ0Z/lMDEL/+72C74vRxx+LU7x22+Am///rWayWQtc4314SK/q6Svb
kN7EYRxkAI3ZNQAZiXrKWrbcO8VzjWJ0HDpZcU1F5xHvnmJtONuwffQiKysbfm/f
43nof33bB95sTCMGjWnBxLDaJ783Jtao/X6Iqq/5U/IY2EY3ZchtqmQ4Ll8Xa26U
Ks95X6WJTBjY16EtOf3sruoX+juTPJU1g9D6dMFzhL0rRSy+xP/HP2/f4heO8Rnz
hO8cc6K9SQCq5BSl+fJxiiVJYTf+J/+OUwFsvdiimPrLRkEHip4yIG2AvHiDMFE6
V/bLKl8tIvvUhoA4rYP7HC8W7mucBUKXbWwZMuSGSftgurmAOChWRSJ3jPQyxlnU
9Y5pBVtnjsSOcPkfwJUkZhLBR62bECyO1H1Hv3gLQpuh+W5pDHLUgTgczgFRVtCd
5c8rIjnubXhIIkeSZbHJDQn5WvlZSVwoN9SwpnZfD6+QQKRjtrxYGEnQUkbhbDNP
i0NyH5hSGugopF1NJHI7drjROQFu3hMSp3NacryosFHUEJUkCRvMd1/2tMQZM41w
iXD6jz+C1mL3G0Z185UP2KnNg8c/U2LUz2g4OL2uLh2XRIiE4xMgAE7k2N6Bz6o7
kK12qcv+VKulv2RiQbk6AqH5YKrUtOJ3gku2lOfsY3UA8l4bopxnDQTw0X+N1X5d
wJaw9+YDLlj2C0qBYeyu9C9ltunaJVWmfHdtJxDrOZltSNoUVj3tccQzpGybUbcz
n7ROuq1dbLp3j3ewDZl7MIicvETeTeDluwfgSd3EwGeyERzC++v/qmidCUrxzta7
WW7pSHpu43XgIWBg6NEfO8DH/IU/GpNyKwxg/tfJq5rNaCUpPreiImOXHXOtB4X7
3MjrF8y64Qkz9wQBZBq2HdzdL6GQDDWlc28A9Un4J//KEJmNuONgLZ8PSLBsm8JE
OK2/ilFz8ae+XIQfK80SS6Mb8/BwnC9HduD9bESOk1Xurcjvnf0fViozgofPLtOm
pAXmsm0ILIcHOkfrnd9N75hWItFfGg1c9HRCnVCK8qjYnX0zWD+WxEhDo8OgGvFx
kzlPJrg4qTSX7Ls6GJRrUDVWIx8TPvjk7qKuANpsiy3Ezek8VpsSvWGOfZ1jd+fM
TcJKc8tiM4oT3iJK8lM5I51CwRRBDn2ooRsIZ22yKsTucvmi+2EiDdMMWEdE9amK
PN54yZkGYmX9JmVqAFc8WLNp1R1RfzcDgiIMq+8M5gbJB9WfGc26y7TMxhKWWvoU
xwLL50r6uoWoYEDA8kP5IQg5KFsj+kQ5noWY0irJ3Cyl6rXRwIP79jsNsJ2g6Wuq
GDjLOEC0qBVLXg665UhNWxIJEfUbxvbSdNso24pJ7TMZ4MiMJpOebcHdTWyBYQzk
5m0dk3r5pgzLPmMwz9tg4pfIG3dsnglX1IZvmBGVkyKGTIUUcitwpx+hu7JdWFbj
BkTp6wUQfZiV448mO8Neod0YTqX7Y2OXukg681FY8va3Y2I3tSBhWAaEFzNISvEo
k57JJxWMl8G/kusRfDbcmV1Ao/qOd7hIea7A+VoIeqAuuBJSFHWioO7yDluFisUO
ShO7mQdZqyjpYdVDpdFC0XrxK5xbW7S51w2qDOGp14h5pq8wSIkBrSxIaAjdUfSK
uD+qpYo925nETGiknK4RrZJmX9IvaezcA3cPzOTH1WBgd4Ozumv2vYecTGH17Wdi
G6B17EPPQvUYksVNWdC2safv9EU5+j4mHVDN++QGCCTa6w/w146pXCOgF/QXxrIj
DK9PnrCAdmwF9f0PCx2Kr4283uzr2ZwYkTXbAnCg7B9nQBs+8BJ+NR428dLNsiPx
U2XWJyBBFYsBXMZuKrDKJ3pZvu6IRb/K+Z6zFR7tqXqPGc5wbJ57J/Qerdjtib5M
iS07oNq9Ty1oeIWr3Nne1s/WmAAUtFlOySgqlaQVYUA6weKAPyH8qi3xl6Cfsk+Q
GpIfAMSSrkjup3oC2ZEDBQ3+inpIzMtAWPjdQEP4UK+fiE1gpH+pzuCRlVpsT97H
qNaJ/XD1A1rs1iVmFXDlQppdoODwo10WNq0b9FNRortxbmR/JaYub8eRGjZIlvWr
bGhgEtH+bW/A5q6VP7LJLtowbpU3M/HBWxEl6yeMWDqoI7hUz5QHhqlEzCFs3NTg
stIi7s303Ks/o5hInklT+kAY+W3y2ZjHbacheheGbxQQbT1PWof8yRhEeE6r1V9P
vVyX+EAukzziqsENNG/i63hrXNu4VOhkhhmLVovauBNVWwxkJQJ9ATTHzYslzeCe
UAEfFQxErAlkSfMFmkIy666XQN2OgebIYJ35t6XxN3eGdaDv2JC9d+598J8wwrrn
u8EfPDlIKhMlXqWl8nDJpQ5mvbLHaUjBYB4ATF+wXJkuxNfLfoYKgd5c4fCEuXDV
utuKzLdRujaIyY8RP9yXCPB3HChfa7ZOLy/0flcq0zzlPQQKx+T4NRAz4GSnDUB5
J5/F7E8JxRRm9iKqS/Y6FAHyNDa4Y9UZB9vmzAT6KBSi3py2dnLA2vYhV2XHGcdl
djxQ+NLGvbI9Q07+w2yfl0KKO5zPdpE8C6DScsDA0L4+vngO4EXfEfdrmAI1j0Oa
veDwnczc2WAVmMBvwtwxhtTf8g3/Z/eICk0WnH04LqvR5PGVTFKhI0hu0A77/Kxv
Nwvx2e1XI4sceFfcJ8UrxACjXWjjS0QB6NaivtCpddJr0LLQU3t/iWsHp49FWdIn
z7O6vFrkfvH5FmnyXbe+AxL7+UZ9bD5EfNajzSWxco8JxZ70p3lN6+x7eOvp4G49
rHkGe01LTF6kfQssSfrUiFyiicrd4mAXfgHd6mS64myLUZ+Efo2pKsg7+wQN7H+r
uqJrUBNKovKtVn5xymUg3JI1iM+c6ku5GsNYKRC483nYdKlOY0GVrkZ17h3DslnZ
YK7NhU71g4La0I5B6hdNIR6tyluNgcW7QQMokHiPOPcnlESqtdMcH583RIFIeSPs
6h8BbR2HPNUlvYbTMlmDydadrfUXb97ZqXUja+y3ECUZl/fi5t2Jp/Ewptwv/QqL
6j1Nwv9lkuNOtG4i4DnybnUot8pswEEbTGLTybiNxP9b4ulXjP9JOHziF971rRsB
UnMP7WJJKulBRgJgfQ2iMIK3sLXHbn+dt5oBOaEiFZSx7+cpXxyTUQ9tCp8ErICK
3DGpjOvMrgVwQAqE3VsRmGVuRNDVt8phgmRQgXjvAgbEwV6GsPh/t+uosiEmedAP
dN+cC7RmKYaYt2pekoR63vy6y91Be9ufOer/nHulu1qT3ywPxu6hQQEiRL4aaLP9
T0THKsTbiaZhQ6qriXvjAF7zxP/SzhlPnY67/fhCuEQMERGEFWLnXVhJJpUQJplw
zHaBLKAN7p0Twcp7riC21eEasdHzxLvOOxhQuxbsTIOLniPwBPQUq+AL0ngwm+fj
Oh62iBDmq1E47z/6DS6qfRnmCfMZJD2BZ4uv+xCywqj7CttOXEoS6wc8Yi0JJsaK
5lDlLSSvRj/g1fIsUGHkub6JvBKxYBfgCv2xbms6UoNx0QYyQG7GHTrECt1r6+fg
Qj0lljlBu8b+8VMTXDLV43HLRDLeXuwXpV1Q90JDda6JlCNg/CSiaLCPxlm7xpk0
06thLYyGQNAzQQbPFr2JcDe7IVF9qe5hVYaW4Z+oNL25NKPo9A7rMSS+qRekaNnJ
RPVhDGvpDek/mbzUkcv8/wVfCF9xxknLk+3XF8ZocqqByDw8YxCDbSOQmmpEbEoz
3c7Eq8qnM/7V6Lfm/0OW6NnsYDkp4oDtLTJbg/jac3PTG9ejdkca5ZwECDWI1pHZ
YEH91LiBt+pTkHMDvwpXNk1F3XP4hhozU1H5ce7TKV8kaUOe4lVNMK2RXSXZvrFE
2rDbu9NXn2zJAaD3KnPZKR2M/sm0E8ul6Z1pfqv/bzmehqz24AcQFtLN5MoR3CAc
ul+Szhy4XsMAw23ZHRsYgh5l1m7aqtroFoPwz7d22o48cEN7GjBCUTjbx1pSNfrE
p7MPqec6PtdZCQqU3OYySMkDqoU2Gj4plI6EknjhiuL537StBtN8Hr0aod+lwca0
bx4FFGSaRfdIazsZMvcHoRzYaLlZEThesV6Gn6jIrV/IHRx7R9d4RH0/4czT6wPm
mei0Lz9fRp1c9AePsHpR6OP6OSI8dF7SLubXoAim3/9/dBD+lVcX8yohb803bMLG
iBbZMCR4GN1IQs9BDjvTrV9uSfUVgGBcNYR6IDsrnQZJJsFYGcpDJOH68FV3tv2s
3HdIYfkoyrKKld5+XVQg16NZb2e+NHActjzG/vH0/gbiIh+5/EeKTPuaSTLLG5+z
h7mFS4FS6BGUAVoytdXanYWSOQhtvuR6UthuuF36xaZeK7fsAsX56SPmpL7eJ6Bl
EfJySC8/mbs9ev0G4QCQ9LEugQvzuis3dwUfls7hONvA2EVa5cgDaK9kKmbFjAEA
EYOOcUSLcl6Ey6yXEJhoQTn9r/W3PPvL8ZjYvwrmTkrJeXbiV9xzeawiT7s2JR4l
gduhopdczljHd6rQnjxuFYzlVV3dxIfkpafdFrbWAz8jz9sba7WbTF0b1fDTWgpD
78pjaYIFqQYTe4gVuY9QhwPpbAWhlkvGdYmK6M3TPpRtsjOXygbULuHgCtUzMCRx
+cU4I3ZCUpa38QWhvIVVBH5Pg7gvAanrWe7S4h2Dxn3AswC+enWXyZuikXKar7gh
2d0tmJIdmsh5z+aBhCgwCS9HipxINzzMyh7mo2SCZGEu/3c8HPYSwWMMDara2CDV
X88Z0ZkIUX6bi20uNAozE+8XdA2+T/edjDucxv1SpdY1YRWgf3Rh7PSuCaW6Q5gT
fPvjyIcXmMY8oacnIiiwk0EyO9upq0KsS6t+/lzzmxZWG7x9YgJtNCHO+IXGvbWt
NhoEzTCwfESB/VncRgtMGFKeFqouDqlOkt0KE9jUqe1dwL2PrGLHvy29AwaTFy8s
IN5+Fo0SojaybTSZDgvU8NX1RM2uF54MCpw/TUTqBiPnWkT51tTbJGVnK6BIgCEA
uvYlVAxLBTkAS7zV+q5ujY3DP8DDnGTH0M/sH/TU9b6fTJU6mLggstlJ1CmdSVf0
Pb8fi7aRqDT++vY9ylwRjtjC8SS1diL+mEUpCPVjBVcXDPl64Gs6W3e7lxYYkeQQ
yaJGZ9jTglXeiTlI+0DqVJs2g35CbUvuK4EO4ZTBCgNOBtlKuNkYBrSFW+Kikm/d
pLyK7qk+2HVNzqtoVa1x3NGBOCXdV7byZMxqZh2pDxgg3bqLxj6Cxct8lrqI59pt
YFuBWUXYYWGwAKqWEGBOOIxnwU6cEHjGThQ0Uz77mvbykhYvx5YRmYM/1z5Rxadf
BggPTcHDrvdo/rzuYzkI3ybCDLUOi8d+ik7rdVSnSBgw917sPnzWHfXxHfc27mDK
/9qS9HAefEC4V82/kiXw0AhPQRCjDVRH+K5Kr6s3ET4+dALtXjyjvuoQZVLcPjsh
ZCVg6pulNmKKIrUaN9kanhg/25mGxmBjz4W1fpPl4yQLaabgDD1d7AAooXn1Ykkl
7F1BT5aotA6kkQ1BfV1fHYcgAiwN+SjDNvuo+7YczO4IaOYUOlCThwDbLvhwA3l/
BmPgTruayfo0d5Qvdk+zyeg3sG6TqIV+ayUHdTvbn4DrqMrH+dHxpS8bWZi+/f0J
8J1KSwGWt7+dxTAJAEyVmWslvuFZGiNfpVuAL4XCVmt/ouP3Jh8Vaiw4KBnqTKxK
c32z3NzL9fvgLB4Ug+R29ZOd7xgBzgu/EbgP5G5ihpxeMms0zPRjEYvQKWERkkSR
4E/5mfJKzGSrADScAxVtl1Wgd7vJy+PpcWBhmYN9oKQD9wuoGhLKpgGW+xAleN7j
nPq+gk4cpcozYmzAi3km3quP2f9ksh5qf00AQHP50eseegP6kqt5r1HJr+5iPjf+
pgtYNkCGB2QlQLIK5pFd0LSy0rWO7PYJu4/r/Qor9NM90qswctDjorBWS/bMlAC3
Yt3fDzTUo9xDiDcKf+gDMJVPgCy05UO8ePzQXP6/ZYsgvisG8yAX8IqA43Rb4L6B
zmzBXsB1P4CcwJ7PkgPSpLJSD8o528lQSulnlfnlkj5EfnCBumI2vbN+eyMpUUAO
KMoq6P1pPj2Y9OWNphptY6iwUeKjtFS1u/tfErzl7Ltf/Xt2VFI4A4gfTJv0RMtc
1gUcbx7O/L+ikqmWpiL3ux0+7ssAyhK4GFKbeoj1jYXrDG8Q48A7x1sSk+7Tyvnu
qDGub9zBxcWdbWblnTVpgWXyRVQB1yb7rRHf4PAWRSnYjonRok54+b81zb6uKYHP
D1MJGSzd+YszL4fGxsGAT9jIAdk2ohnqgEr292m5OSWeJak0fHG2xNeCJN8MN4eM
CZ8MGELIO/B/k2KQltXlQ8X1VyosE1kBdQgXOPr3dTgTqKRB0IIEh/PHhSDRG7ge
hH+Qsz8ISj8mlD7nxy4nq7E+O9TGhmWbIApx6DwPbWq6FqryEawiJNO29KRBbsTi
lV6fXUiXW++miY1S23fyiRIgbwpvXfC6qUYK+CyH6qhxgSdC/tW4JYpR5ncmT273
1H0SrtezEKiy+VHq0YFwwuCaudIf1ea8M6NA4Kfokw9eyTL67zww6siEFbuDyDiT
xxVmdbTVccphKuZgL7gU1GI3OG7gN6jBOaWp+MjAgW6SXw69UV2KclT9tK9yh+E3
RS3r3/t+Xeg/iK6LfMwPzPaxmoBPTT0OAWczQ2qjUfM0lAYlYr7jsC+ELgP0HlnH
orDRLy4eEhmTBD37N5vyoWHWFVGxvzxXifv6aQOihiCybMS0k4fH+DbvMDt69DoU
gnUZBzUdSIxC7Z+cnVQ4ousDseS7jak6AcnWPtBbpKVTgyLE+NoP40h0XHslQsZe
eRzlELFPAQZVpSu/OHtz/CQo5Ijvmj8wGvbitkdgIyY6taqZdrF47xLMzAV4kPkr
GbVjE75E4e0FrIcbB91gO9qzedmN2PnW0KD2XQNF2ak7gy7zRgPMsl4F16UZHpke
W+5D/aDTFOn5CVQ8HXVfCMWEQrNNJtJqbaHVQmcSo2Y2L3CXzWKUnjL6sS5mfS22
dobAehQhwPZ1uAKNZB3AxIuMtz191AAZxlU41HoWySKZsZ/uDDvK6xCsMJDyrXIK
GqRjFHgG/g6uFRyDZphUDtFwQhwRUW4+pdAUpXM3fydAwy03J09NA+1E0EG6i85z
lvAXoM/zikYBRbijADEx6tfQt7le1UooR6kwNbK2fOJ1kAELqznWmLmtY4IDogVK
WXUEWpDhH5ulV9s+oMZPP1TfkMfz7NS2sMoxGdf77fjx/jz/GbFWKeSh6mC79c0N
fw6B+hAYm0nCcxA9AMPFgar3sMCM/jRuOxlZ4QUSQ7p5nj99J66vUCMqKDXkQEOU
ZOAi81OKGmbClzViHSn0ssQFk0jrYCzjTRavI313OwMPwvZ8TUlSkC2Pjz/7Ri40
zmqg9H2fy64epRtWObtSjoty7MVPQo8XQpSCbKxnzBG8rHDdAPCmI2pYnINqQOhT
jF0ZLlMRpauvSvumg98sgXm+TGNkwj9T8C/3JVrEZV1IAS4MkrbQUGeGQJLUD7iM
s6ACd7bYK4ULCNh3dg1PptZ0owONaVbIEcD8LIDbQJ731qnGGR3UfHTuqKleg0eh
UlNL27pOOUaQygU5P1eyZa4Hb6YuePsooMmzHKkUAgONDHNKxGRtsz2w0DdFxbJo
veXnKZ0w+1b39fc0LgYpnhoc1/mJm8GocXA8Hto2jPSBolxl/C1flgnhb3CenFfL
qfL2zCYaVojVFKj2jm9ZhxHnG0YKSi4pldvzVtErjM2rO2DF5SILQmCg9wLO/Fz0
/N+tSPnuHgA2bd4YZlWdefdAfLRQs+y+oXRSnZYZOeh1FoAWNeid5OBeQ1FvVzLb
o6NteU7djiAEEnDe6aFw3SagiRVOe1DXrTlTozC2Ae+LkZWw0/TKdvnFkHwFngnf
dJg63OzrSx/nl/LbJzwzhHrZF/HZlFjFW0fGj3LE/WBlB0L6Nx8h1JOG5L89U9Vs
guulTgEDclTdVa6R4DvAGhuamVhOh85MGKtic3OoBw6Vnu0cdUQRbghfAgd1dcV4
F+TL1ztzbFH5EyzFkdryfT8B5FzQVxkYx2ZQZOXuJkDX9Gs9Tw1fEmNkSlJ9d8Vq
k9FkPSb03G04SxMIoHy7xJegfy5BgzFvIeJeBTl8ad3/O8eys/2QKJtUOfliKEC5
vY5z3AZ4qrSvNDqswzvXDaGBzxTgpIT/Gna4iXbiPHU6QKQB8FIZ0fkCH0pshT6X
CX35rhpgX/kcY7pgP5NBr+opg+SjRRtdK9LWyohFMCkYqSobpmRrntJUzIDvSbMn
ym1/5tQ6VExPMN6PoPqmS8V6x3FQLVRShCMVkdbTeRRraqEl430z3qk1RN2xMzdw
dG9vnjwbtmXMbBVT7r19B0LrcDl5Rd+cmxH8GUb7OLzvClp8QdhDP/SA6/8D0oH0
Hwg9N3BDykEUk9Edq3MaePL9c0Dn6JrFEQV7/IUl3PSEcrPNMTGcb7TZwp7uvnbp
GMcVZ7K+f4evzTGDlypLNq4jDRFihKVuqjy9UXGYCpaZE58dA0K0fNaf0zGzMEGl
sGUG0n6jMg7d4jM1eNnH+vdOaL+tmVZLGZ4eQgheMWT9ISrGfTz3lk0q+LoPfsZe
vh/mp77UMKDXXTadwS0l1JFB76QO01aOZX9kFRfPKGxcRb4XNDfecRBPSRcTDYU/
OJXUJw0tuVUVkpaPGYQpcLr8tGwcXO/mSXzpA0qUDzZfn+4v8XN7Y67x6euSgYeF
kwmEctbB3grvDRoYrAa/H3TxIyYYrbgSc9x9uHq5Q+febG2d6kSvcHLzKrPEW/+O
c1YBsIfRx1Hv/TRX7JWuQm/8CRMhA6lPgfAtwJwlrPmRs8SRXa90vyK1QEfQQQsR
1w2Z+bWfW3LvX3DPf5/pKyTbC9aK+FBJx6MZjgYM/cvmDmspbcO99rtqU7nRDOqJ
1g426snOfIWZS3WhIgXYowCmbDuMxWN0e+0Vd+1pB2ZP0YbyddSBcI6UJSvba7P2
JujuCmSg/If6TaIf+oiqsNZmpKUg6UCAzd9JvUd72E+ralGKvphu/QuGxBwqNBXE
7YPOrhLdHllEZB52EWOflTh6gz4TvxB9xtH+d41Mzca1Wdg0zq3Zh5LZ67mW2KCs
XgUnzP/JJQYH/B7pQau265lGrVlOE8PIG6FHDQJxAnW8AcF4C3Am7ranWYameeAc
6vlbkYeyvMFb/+ovylBHUftRNxeZpkOwvBseAEmOwVUSkXN57GH1qkEtUW+eCcKC
b/DS8pNhD9lG/H12QgYQjjgffjH4cBWMdQbKfP11bxe7KC/0v7TJ/rgCtzUQM0Rc
GOEp0/mME2IHSEOw0T836gD0S1N6q8xgtaiXm88LndXlyzMFcD6DDmr9XxZ+8HF4
4RmzGaBIGSKGaecoSBBXsa6vdHNnuZdbvPTgrKWqj4O17PRPWtsVGeUkAoBsY4Zy
MqBtcUcen015a44eRfi/EJe/7JBwfS0P3q+9ucbHhmOVpMuzrmt6LGapjeDCXwmU
sC2UKOZDwKuRK1Zguh1T5Kz6hmk1jpbjee157qrN/xmOKGYxSaCybx19D3IMTFCN
iHVI8HdKYpwXTSfsFtW+Bth3pIeXEtXEkY2hrCRjjFkOi1HoJXojFe387BiOEkUs
5LWQ1GsBGYTNTA55WnlMn87+NB1IKoiHncsn/3BPJtmth8kTxJyYmS9XT/P+j/BA
KGK8NwnxFSsn4SObMfhp0L4Wldn6rFXyZvr1S09d7V8NGTp8GOsq2BkZXqKUp+Sy
VxOYSD83xn27AmMHBZ+g+1iMhHhExFDS7ohKfeVZfcjFe5k7nMOMBor+p79XtQyE
qnyMlCs3i8Q+yqZWM/2RFbEcNdsC06Ca7nyQZcsOwd32NdWjeLcfBqDp5qA8wBj3
yfsdt+9XrBEx1EepfZ5DqyBxCh2J783lWOE4Sqqtp5Z0ei5OwmWVgtUFsSrjgAXa
QPVw8gL39+X6gDPAcvsfrTL2MaavTk1OSYSsqZzHdG7lBkTWZEyqSoWG0bCnQOcz
XOwAyxdv9JBPiJxWAiWAX+KD29fQOc7gw+49AZgqDSFlkJfD3JWedTvM3Ig1fKqu
amrZUo8e7qAyFYpOCgIKSYsFSwlKEIoFqd6KySz+4QqOu9u8vF/MlaNim1deZVMQ
DickoWvd7xy/uSLM4pvZU/FkZDfJXsizyTyccI3vkRsIwJqqp81ije1jc5bkHn59
V9dG/h1sYrPKnxskbV6Mk++3kkwy1kOsaxeErjINK4ojsE5uCuzuZuvpsOiKoKAN
LMQ7aDs/Z5XHFvjcL8gDROZv91pIKUHo6ebYYoxNaD1A35dUnxNlZAR4BGR96o7B
VhmpKCty5XAPSJnYnrz6SxrD2VpPETUHjF2iFvvU1sRQ/TgcQEe6Uuzrc3441vHV
g5Yw7hrLG/7b70/lKWiFGUaz+QBZ2TDFen2uLQ0ZcXVbWxCS85tPz5w5ITLlWZlO
7uHXIufOf/JSCyITlRnSziEZ23KRQMnJCQ8t3U2lLdfWixet2Kkak9F3Svus4Vm3
VRf8AbpkmN0h6HiyfxE5sGmEVgaTsF2jEXJEPpW3f0GLUki/swCa4Mbzv8mvQxT1
ridCd/esNXFiYOmeP9OAv8JbbqGK36YZ/CQXiEV50DI0PL1TlutrjZrj6c5jpGTH
oLugS4+Lxx2IaZa3IRu+v3QeNcXPOZAbpp7aV/2U9IPNY0SqzMpq831Kz+BFNwji
tTZu2iFw/z79ZAo2stTtDOX/l2MF/kJD5asbxN1DL72G3u7IoQSv8g2maJ3du+kS
TEsOZzTg4u0bnx7fkPK5t3RwvgHxjmOoS7QczLlJJ8F4GL67hvcXFZUARHgb/TbJ
b2lgAFpBKvrzP64yOyuAQWVkKgdEvcldhiXJriDCHk8J5E+F36Oj4E4Ow+YI6wrM
0gutfceY9NScOEh/TkczVRQAZDcKZSesl0yKUZjaaku1UpTOb4hwhyPp1kDJWINJ
uLNfVWukyQ4/N77RARnqfKmpaZbl/a0HpCvpcEhfjEgyJn6+3JVJn0oZk+HN8qaI
dOBS701QwuljoNuWZE3SDz7S8ah2+qvdoNGV7/VJobyotWb3ZW839s+QopszB9nP
NsWUFHBwXE6RGKi4DNxe5Snn5vr9HabQJ9SPPpCM+wbTcUGfHU335fHhl7ea9uMG
EOz2l39ccC6YB/ANGdJN3mXd07ZmcuYkqPdFG71HT/QVk9piuKfbmWt08WQWJ8+z
qyrwDK5sCCKAFaWMsgwRMK6mWKtZf8fnKX2idrzyv/C1DLChRMxkGZ+XpDK+nlgx
W80XvWHu3ewUxvISx+JAcEfNkDXHHjeTRZGcUshpMcZcgpCGZCKWovcm5cBkvMJX
HDdQQ3hEg8eNGfwh/LG9dr3VJvdulLX1nfnSChIvkAsJg8Y823SZEar3emW9caM1
ktWrCET3pzg4JXqYDWz/krhA2orrKCqTROP8lUagVEXItYvfHQ0c/ALUjOU4kplc
17KpblHRzjRz1h4gf6MZYUxDV8aC7xhB8I3zLFYKwMxHEguFiEq0mY4bKfPWfcrf
WEXHDMrzLIREgrJYOP+6QrIUixOCxWdtwxSCP6GnsmAQeNPQiDwMttkSAsC+9kE7
jwZND3iR34Qtu5G3WW8aOstk02vW0/Ww18xpgCjfsQmEBo2woNDjZbWGZziEsrjp
kzwOE9t2sRQZDQ1Fbk8NJ8dSelmUe4OB7BuEniONcQuRjFHl2/kDQkvk4M7RTVkF
0Mo6HafTEOT1MPbm66brpk2iYPnANYyS9JtJdg4bqDvbQYolJlsJw2IzYPERIlt1
kj36NgasGoIjvEQS9uFnd1ovh9x3en7hmOFeufW4g/Zhf5ZDrIbCxTwcyCNmVOII
1pglO+llqg21GYUNiL0AiawZRzevFCY0fkGgPUx0H2Fj39FN1NSos4wMXoBHjiPc
u9ncnI48qfUveVPsuzVglNI9v1Lkp5MvTeQIgvTCSqKtHr1o5oM8ZoSx1eFXHywp
DQ66rb6XPJpoTeLhmy7Qxl9zjy9IKDDf4QufNsvUN6yDdhpoLiUsPG4+5h4rmSoj
pwJuKr/GSxC9O7QGlOXj4sBaG8W9yDMxH4AX4SerKaohXyDQc54f6cG0rqfkeeT8
VfV6AqiBx30IMGkIaQYTFdPvtGHKuJU5JK0USnRbOQNNlc0TXhMdT1NqG+/qHgAc
gBChsj6SzYKDntOJ3x2F1qGBiPUzuzD4sb6ye9DkzS0etzs8ojIFS2JSyH494eJC
GbgsiaLPA+6SI1jQ6s5n3WQtSevJxupo0B+cSWGXi4TVODi/JjRw+euFQOw1Sdkm
jrviIPdm0in+RJ+T7Hi2w5JlyLj2gWyTD44ZIxLh1gLJGE7uDhxcZ6cx00NIquqN
x3LoT+B/ugf4cIODl/J+t5WETQTpCiV1bnPqvPPEemch/40j7AUEeKiiI4YTaefj
NtGTn2AFri8v2Tfw05MtBzmUob2wPTOtuLF81jWEBGebIkjNHozde/HI7e7scgpw
VnrvPQwur5pMtudkq1lKJayGJu0uSqKwm0LAw5Xg27jkm9+DOgBvpPJMa8vTBRiZ
OQjO6KaakGxk7T63wro9WCvze2W6Ree2bJefNmgoVkk5rS33Is2Fb+ddjfSweiM7
WOauiZCn3jWIrOSyDM68rzLYm0mwAyt836YvJEudsW8xSC3a3wkttscn5R2OamAn
MCjz6xXcfjsSplOhOR8ZrlLyIXZPhlGY+DWyb88WV/8M6ztNVU5Q9V+ysreMvWMR
QiOr1fw18pmvz1OkQ8gTFDzxlAk9Sv7xw7J3OQpoT+r4ZVKUdQymj+4zjvCFZ5cA
B6G4w8aXVoXHV3R9hCSQEr5AncQIXGGV1k2IvMrhpHIiRFpUKCdi3DAqDn5G51Pf
lFaHgkomonXtXmcuf8GrA5re9dc73jKcpOoCes/SgTuQE6fZl5uTOisjMPt2caiW
98S2QLr7mhWsLM+Q2ulUIKMyVP0A53rHra0O/vuW/ybl53VVUAjjMF8+pWQ6cHnN
GU01laKFEsH/x0PLdKFixWp6V3mczNh8AdBfsL8k2vXTjL3EZoL65L+qcfH8X8kU
BZtQr6BchqCTdDUkxRcxHh6sdrOmu2dIIT+Yn0LLM5WNJg/NXRObtUxsTqEY74vR
Ve08IvS6svblQZpf/dXPGUu9qniRWd9EkJMO8FA/SKEU2BgJZBjvS6OmTCQmxE6G
5raLU4tsQNI8xe32Tp7VVFAcUWnMz+OOrcRyW51ZFA/DYGBPzJsWhxgHadNGN2RD
utxPMwOtinYR2sSrMlUN4zM6c7juWHqxLln47Upp69mQJ3nfDs3qSmCeGAS+Y4Ef
+wnKTGJVt+ibsgao9F8Hc+oHMDbnmBZ11SNaO1ZRQvw8XP9tdFuhzeWCqOyLOY7L
SzICKLs2kKkQRTe1DfYeu7rLipqUhq7J0bQJ3N8wXxvi7BEsS7vkheukhKqg7lqI
T32faMAiCu4nuOZHAJBYYbsOunVBaGroVEc8GkmHVtP7i7qAVFwAmb0PZhvBnYQV
hfZLMoL+caKVuppPfOTL13k4U8tIt4hJBIaQGoiy8OysBAFWJLHXbFxmGBi17Pr+
n0b8BjO7PChyH+vkyesPMmYNtZWqfu00oIX2Gb5Ht1nxgzAjUI6ilbFYleAMIWuJ
jX3r7w5EplRmKAJcelhNxw/8YDdg8N4v0StcAWV8I03uJJR8cB4uA0JGs7v48xJ3
bODrxjAQ1TfpBx6DIaxhXxws4C9hXaWmqlV12BSXphWZwTIDTA01tCDqiEyumUsF
b3QQzvU+VCV5RGgIEf5aL4Fcxcp4RAL3mPhJAHOKqfjrvhKQLl5g0TB+YnwSyrhi
rxD6ScUN/r3P1scytjoUsGJgB7x2hyIpbyNrSP/OT1rnLAXlKzBaaWAsDZaoqyu5
XqY1hj/0LAqzY2W6j0S0v95egZG8dzbyN53MHq4HVUj6yqkzX6hsf57qi5j+grG1
YyxAP3SGCpaNbcwONqiufFsdE7R/ufAhoxCu4TEtJTpCTowzl21K8Qjeihy+tteX
8ZswmbCtBBV0GHIFXOoaN0Ch7lxBl03QZPi2Cq37eRZ9jDRov+Xl80B77O0YlGZj
aHtjPHJnWVZgkjDC/1e01zbQVxcHxijix811zNA/C0+4kFF5tczml9HGZ+m8Mfvc
jJs60+4VTxxuDU/YIGDZ14dOsmUnoIuGds+8v5YFhkA29FPN1RmxdTQkEG8XMEQd
xecHnB22vjdCr1sb+dCO3XCt+OfNt+hRb8MxbW6g5NWMoDpoOxceLsTtZZ/IuX8A
oQ7smNtd4GxA4Ye3MNGUwdltkuUz4iEYklTpDHGPf5MWPr5RANcPVhW1vU9nX/86
z4tdgdaTm23Gy4yM7ldfbp0pL4iJ31KOL4sk8gt7TuF2TaXSLQxn4SASbl/QblUF
9qsVtNwX+XDL3t0RsUjabXVQFjnbfXudqq2ojoIT3UiiTTdSlG0V3NgQEnfLMJPx
aWp3eSm5GBRg8N3tBdct1dPBiqh51h5fKO5iTnugl/KXj2AW60xhmfNutUl4McQY
avJ760S34kg8VIemwWZYg9iIlmQHXHtc4qKQRHX0UEOvZxVPFp0EkfdclDQH5HQb
cd7Ue8hqr4lpSJaMV14Xx55DEApMZ32ZQjD6E3I8w8eWLs2FV1zx4Wg3NmvQBRfs
cJpQekkjFQ4omQJ7Lga/Qgw88Dpfe82mKgRErawWVEzqUh5sDUwk/jwU+yccWU/7
al3GQawU64HzVw6WIBGRK+F5fEQr9mcFCTqFCdezAujywQLrupUG74Es/htqD355
4kwmN/TaQ4+wugZs+sztFA9/LBsnoGSGwjwTmG/1fMtngq/WTqfmRrbX9BnIayLp
4gzF7lzSJanF0jXEYU000HqWuAAZT1jRSah6FsH+y092/+JsL85cjUlji3UOuh3R
BigzHAH42b0fiUyziCwTD4gvPh38SDlo2KdHMoNX0HEvgTaiSuJK1yrnAUsZtp6k
f+HJ5bmWTcBTD1G3aHr1sX4oDeOy5Qx5QVFptgDj2bhX/vfyr+gmegqSkqsIljKO
BAIYpvc56i/vGhkYJBg5TVtlxTcQNDrhJlMBFbF3P+IFPiDA2yYfqUskvhDjmPUt
HW6adpX25Rd+ca+XJkMPtsnkGOGFbp53e07RmLph1aYaBgo4EOgczCWlOuGDpAjB
JePAzj431bz6ZraUuZ5Gb2kP73IYuKHWQRtXMf5mESgnWFiJt5spNAl2c6BqGZMV
FjgQ5vfLOLDE7Kwi/22mQr9g4gNaxx50lqyNebrMsM8aHKjsP7WfFzWccSsR8Ply
kX30fD/v7OcP6ELR4yyq00mOpv7mhq2PfQWeCBkB8iqbrDGnU9eKjtjsW1nlsN8h
kTGuRlDSnYX/SpEgZWfg2/cvmlPDQD/pRFwdKrq+V1Tund5XhzvLWLobk1AgEJs7
t45HWrpfDNf5+GCH1apFdTRaTtNtoU3oecWQMPP2+OI0C6sSlHQpLMWzGvhSY2eg
spxduKX/aWkiwza1cTCF7tFgWYtAmtELk48FmoksofEET9hWZIucza92sSWaouls
J6e8sryQMehBpnBHhHdQ0jAmZYcSd2cAIgYrZ+vMp8HU7wKL6isxHwefTNxu239z
BadNWmggKMbiQcouWnxw0DX+DO0ff/kFgNck04N+ijYNwzOrV7iIfbH1ydaWdP+C
XQB5vcQpLD07zvI31elb/rGbPOuwZ9qQs1I5JwxJwUFeeLYZWL+dl+u7YouTDxok
bMFtmnJQ+G3ot65Nacw0JyA6g/5xh3MeE0TIk4VK/9bZLUNY/dR1r0Nv6oqDpGoZ
igX0oPVJJvQkK1iGWjXGUGDSQyXwrTtt6gh05ghFS2YBB4KYHfdmDC0ppjWXKk8F
iP8k1uVIoNfPFNjxMX8Ge3U7yg3D5hrQK9ZIwV8kJUyti0JTqzEFCRsTEopyOS59
vlkzRSKaTPLNMUgInBLVRuO9OLbxFX6DF4nm2R6Zrpk7ak3mBAfnvug56seyMaiZ
LmidTI1JgEug8j2AtP35pmC/e6PvgO9wEwOBj4DSn05l8MhnflhP84nlOMqiiHB2
f3KHhPp1BnEz0YueDYGqcLRR9CAJ088NUzaBgKYbXfeT+9LNVPHyOkBPvY7ajL8E
FO6huDL1qgt81cAggZfbsrcUw9shdw+lSTeO319k1VquVpymQmPbEpY9aceWuO9s
8rP4keDRKKLpVSUrFY8/MJmck1RMXgJXgavUhu2u19MqcHGj5LK5tpub1iXHsIy7
YzeS7Z05CRi4YJ+e2arNiGFrf+IClSLYcL3GS0JCJ60d6rf46y8NPP0N50i0YcIy
DiDHn/ncVa9DKQALSf9x7J+Sv5jO3BKijA2fIZ3qieF6a3fL9ZVZhtLd1aQ2iqMO
uz7MWgrK2V7cZ18XNi8LOiNFgfR0BH1P+T7rWn1fXMqaDbThmLiAmS7YiWnm5PsQ
IqV2/AGI7p7zVCW1TDhXmlWZTHIMPtA0m43Hxk4FMc+nUcCmcTwHiiUm16urDVq2
rjs7nLdlf2kp6YX0/jXsE98mMHvpMA0gYHUpVoensvgvTfyzmfYFGPoBU1ZcvZsY
2FO+HMD3Yi/ARQtJYQxZgLU3EIw/WHsNgMFmwGjSK/wE8USUan2YBzK58pNEaOk+
9JeIWsCk6bWWdOXWsfESHDhJqS1+5aVZ8c44xTqqra4rFY817jc4TN2OZBtx45df
Xu6iIZX+UmJhPyKb/KaTwTzap6JH8sk1rLFc8kwjQIyuIdo1kDG+1ud+++4N9d9Y
aNInxBgc2oJjCsKbzi3YQUPU51lVlzo8v11fD9w+QV+ejXuBFkOfrVW9tlKHEi45
LycPld0JsQ0R5LHbpvgU465IzXEY5IjZtzt5FINg3On7f3TRjiY1UYiZZisKst4T
f457AD2IncS93585rUWzKeHnV9F4wDOtVZB5cv+6vtRN+tQF+xjEKK33to29Tx1f
7hXE6vUbNf1APx2vW6A8NC+rUlA4xbs+lvI54mdWvlFGjQOIM7b3rAzkTZ5SRD4R
rOoCJgEEXD+GTiCIyxlDYJ0S0pOiKNguWrZSEYM4yxI0Of40EfA5om+2Hsa2BBXQ
K1tIZ20D8WRBI10arooEKgUKuPRo5gmVvu+LXcQlJvyRsQiHJA9PRxS1WDpPkE6o
f4qbJMBFe3WF/gKWk1vBJ7CkkMYZzJbdIk2cQae9DwdVtaEKB/dg5WPIMpwLRkZq
Vms9OeukSvjl/MPCSfTRqgNS3UWfc5Zqrt6oQZ6NdHF9ncqyUOshRhKuNf4rEThC
Jrq8XPCSspJOPgVw73puIYoY9fMS+EHqyvANS5tpRvAlaW48A6pY6Zt4PtP37ZIP
XStmRuKRPXUZaWkCRXWA+eTe/ttCXiJfMsjTlpYBp15m+PzR8T4SC9ok0GZsY5fy
n2+aX5WyKJlpz7rQkHGAnrQmw7pERktu37hPKw6WVMkK1M0lef8aIdH9o8UWyMd/
JN0o0CswCGzUIVBcE9biPgw4eVGtsdm00xWhYkYQsYggR/r1VqirMVk80Ri8GXpZ
G5AtQtlZ6yGDEmxGuP7zBdhgE/CFCNnDujhxhs9IwWtiVzAzYNdWnAVBPOTj3uDS
uqSuLdEH1PWiH0TsX4mYMu9gSECIeHnm14zK1HTGzqawoV6n7VoFz4uApb2Ht2GO
FzhqzxVydRYrg/gmJeoao1hsA4pG6EYrLNeUEy+fqC3QIQ76g3KploXxUDY7T9/q
ZpEEEo5I+q3I/HuNlFk5uF5KjJbCeL8aQx8ux1x+VjpopWTR85f+38bPHObEsxxr
OBRi7WCVFfqjZP81oDYAh90Qiw8oJFJArZ7xUnm/F5h/mN93b9LztoaIHJYaax8l
jT4Wr5Zewpo6ywM0WvIAcejM3C2zQAV9jCfLuWqp841rC05jRmrZ4CWzKhTtwV4R
bJc4GgDGwHmx+YDB6nfotXOw2S9Q0GUv6dAZK9ZyyDDmHd9+Hlug0V1qFMlSTYyz
2RB4PA9OOFWXI2KrrixFe9HQa46zY0QT8q6d1e4XMqOTd1dl+aVdKvOnQYYp1x53
XQea3k9ZRoWw78b1894MSokf/6l1bYh7pBlqF1W3UWivz/sI4JISMZVUJ9qLinO1
MfsPKjxl7f+bsvZsD/VyK2+4yAhWIYAC5RINI0PE0Ui6ySCV56JbTRc5DfqsKBiI
kWvAsLHXoRx2c9UmcVT3Yy55MiAYAWzlJoiSxmdAi2YW6yI0Utqgz0PyoPot9B3w
FAPGeUcxyHfn1mqmxZcLg+GmtYSTcCzsa4zPNnEcrc/HSD+igWmh3XfQzXOp8pdR
HGk+mpUeYOqUHVKZBSWR8coB5cRpn+x/njDI0vrVrC2dElsMWl9yvIhkijFWIHGv
c3sNdwuji4LrMwXz+OKtzj+bQncOaOB7wUpB0xGuv3flboEwvOdS4QXqq8kTLmj+
HP1IWdop6qjBn3IAwghOzTaVABE1LTTf43bKbkHVF8+jR+XIdeZfAsm3xqSPuY5Q
DTCEAaxemMemJbKr2Pp8npac3NvCpqcuHdvYDnCNp+eZtNuggw+F+T6+Nq6yu8et
rHw4KPQgz3D68l+bqbaK6W09ih24tuKn/pUkgM8lI7UnsPSuVqzmC667OsmCQA3W
GOKsGK6WkKYSg9T4clGISE6td2lhgROxKio/9rxWMgX4ADeNN34Aqw20VMDLQadC
ePt/6xVyd6L9I64QomkPg5Hsquv+3HaQgdXh342btwpjQMSU9WySzSJ25lA3LZU5
6I+8uKnbUUCwTR7X1TPO1vIsDkvUZL/W8SWTA8vYzirxu8ENikcKyRBz7EKyEeK7
IH7+aYVlrQopSGkmF1lL5dmrg44ATIMeCpxlKcD0lpH2BHzhdSg6AURDakCWi13W
J/4QXgXgb8ViOVLavU7K+GA8VUqqBACa9gTKsNacDyCp0dcjayzr3vI6tA5DOOZT
NOaQW7ywNQ7fTgjoZuM0sp8XXS24QaqLh563qJ/9P70fN5lp5A8RHvDAscWWzJOX
b7OwHxtS5jAVsxj8PeI/GYrWuHlWKhMQWden7E9jB0ZOpttrNxrz6idl/xWq7Dmt
pcDXejniB6YPaDj25Ct3j2erMkOPDDuJi2Uj5WP0nhrbF5YpE2pEqG+hv5JFcOTY
oIfdHYtglj6+52lAHScfp2xsQEighVzOI+Ax40EGYkdonmbaKZlKkbqJyTxEo4aw
XDGV+SbG6jiJMOlqRhdV86zhx8g8Orp5Kpw7vpBNetvI1HDNilviiEvXpr+kTxbU
oIvpizSeBUGpxfjoi6xyE9GjODFeASbGVvGevG17wXpqdVLJjY3Wc7DO7T2ODOyU
gfgJtsuwVE9PqS32P4iMYf2jIHcoDgb8+2Br1oCNKGhqEbv2Y8SD+ZJURnY46Eyd
m7JPD1UWWEymdm/3GSExNarPil/fSwADLqXUu77KzFQUXw1qnxCL8wEihd41kOwU
A9BUUigANRiWYeVGnit9DFrWcRV1xL8Ij/paB7uQARkp2UBBuduivVN2Hqj6Daw0
3DT6IU2sOCSGyUK8FQ5D8VyZC8lRuXOtJPGH0wls8EBasIVpr/0nUNXgsaKEO4Ea
NdjOCjbSf5NSte4OD+OT5QTuTpmKzy86XAsZZ0hCLZuQ2QX4Hj40IDVMEbCOGtdo
NcdplNsLxkN6v8EmEVAYkT05Vv1f9k0ZICph4EVKEtY/duV0iqPIzn+W/eO0xTxs
jekmlml1UurURHEIGZ163/4oQs2kjB5b17YpORkscAaWlFOJ/uo2QbnXx8Dn7Oxf
TfO6i9mhJW/7Uz4kwLlZHGPGvJeArq/UTwP2Ve96pSinvpltsmi7SIcHQP0k7TVY
n+CKnAgwVX2FkcCmdj06gPbhHMmoekoL8FQ+6TPFgT0IYZsrSn6j0sY/j9PzRaeX
Om2uGv527e9hIiHEX1G1X8EqfMwrMOzxxZPKg47Mu6AYAM5E/vUKNkijlTktB3/s
C2rlITuekPgme12PRsp673Kn+0L4b2gPDheub0grA9hiVcydQ8cbkrJICly3EAki
YUdfZts5SGOtdu4UuExvBnBhBl8W4dXQPBOTlmnB8tBXfqsfsDfLfFx7JvkUQtf7
vfKWSdmKzxzWGv3e8IwVTxPt/bmiKE4WJr4itP44vqMgN7PNdY+OQWOzh0EP3pPi
GF8zPHSI+JxTj4aAjzxIfTnffOwYqzrLaGUymw92IXpy3tTG4zZMhZkFrYHtnAjL
tMsMw4le5DgVBaux39As2X0G4tMdbziolx3E6ZktdzHVxDQ2Wtt+K2UFWV0xWdtL
JHkTekU47HLOmfGuaB+6BJjSPjWLLqfAGN917hSuPLZaiMJq/jM2PbS+8bLrHa8k
SxCmtywiVV0K4jW7bKZ900yxKIoUizRxQOvrUXfeK9pIPPP1x/44jDZGXK9tveoR
KNKzw2m0hGC4BTqYReiFjYJYWyb7tJzx8t+yPurw0t7A+aUvPphvhMsBgr8qkBtj
DI3tTpDsgSeuG7tJvaEBO2HiZDpMHGL4/z0Th8gwhzsk/JTHgSs1TuOfmjJPkuOX
yxNLjSy/I+RprtcE65mIIQeNFANwA5R/tIBCtT3L/9ANcCPLM0Ql97OnWWjgo5V7
I2GGcuDkMAQADz+7saxZ7ZPs0OIzHykOcxMwFGQzPMqusiLc0/ucc78CDyWO+Dwu
tQKcD89WUk8yOPliA/xCTVa5y+KQMobX14SHdkFk3JntQwfyaafP5yuN/XcH7dbO
YO0V/aLJ6Ke3hTgFplpx3xl3Q7qriffS/vS2/owwUh9eqNCxLsCPthZg+vZ6Qk/I
0SYGuUPYtOiFTrupg4dL0FLXER6oyCIzkj9DKP1q/BUTWLILVkPPWRJQ31CJv5Bf
jHrmUcKQ9AKlE/UrV7Hpogl0Y87MfxQb9c9bH8ZiTbawnJE9rW3KKqT8mYv39obA
k1t6yj7RWgRcLLMFSW9fFClKCvUJppBE1JONM3wUi2oSO/BpbB4KwTlEv0aLmY9U
+TdqD5EQzvnuIe7QvpEGKEA0nJtyPvE+bkIoxQH2VEiE2bmwHMLvXt8b/LYj9lfH
d6SGh896u2BjXcjrpxh/GEWNgy47dRiA0caf8V4okehyKUGl9Qmu5fvRMo2tnBiQ
XNWx1fY0Fl8C4gXYt8fXZ1WN1dLC+fGASk5qsfAjmw+3vf+ZmBDzZS1c9hKiyMeB
ROy+F1hEFMlSNIEviT6U5SlR1WDwCQtCRPuu2VjV9I62vIdsauqGKGfpGKmPboRp
ZxZXLJlW/FKSG9AwUxaM5a4Tw2HJpU0HYJGYwWTyZG4J7TsaSuCk9KGTQoxkJ0aF
esY05OY7HLb4uhtU/ajOQ8h6x35jx5MQf2OoZCuMIDSSzPICIUqFnC1GyxiF/gIP
UhSVOTAxPvVRqz1FcGIQhAuGV8y0XyG2aN2BcUbusUcPLMbPbR5zE/xpqqo47bOo
TrUgNGn59+rLpqwbHrhNmqASdDt4pCiRO01Oh9PeTcPzmHVtbygQpYNflIAPVtwy
WNxxAOO/n3vAeXgZVPdhDTFoM7U6exIIyC+pYUv+XAx8h30kNR3OaowAM4ohNT9u
9GR3eqYRY8yGhOHf5LhOrDPTZ5DKPx+av7mnoeVf1lyyysC5KaCD8zZXxuWZXGbS
Z1dep8aRtgg5xMhpvfjmCwkLA3yF5cUqr4UObjPqN235xUKYw9FCin9+DTfLMOKG
hxzbsbaQl9q6mPws7XOQFCSuZVCuaczccS9Bd+PGaKTr52qZAwQhUbP5C/jNYWsd
7QUJqrPpgmg76brJzwhfYcbYvb5CztwmeUxd+NAUKHXFd/M9oOFc5BzdEN9L2BVe
HJht+O16UnEnbCh8g+Pna5jD7M1FwBZXTdb/5YA6VZR4+ahZGrrScQM11gi98Soi
ObdZ1DC3BSggAWtjzpMmUTHIq3mcJqH0d9F6wQDbHrUwRnhuGcd8UaU0As7T4Rts
4EG1nzSKOq3u5f/1pf95+KY+13Aqky7bBH5qwo8y5v8CaP3K85FxCo9c8S6DKPqz
rYoBx0XA3dXOw0YPjvOWGS6zcsfxxDeUv5JJ8q7LiKlqzwF3I6iZ34zOvAsS3IQg
TpFr8G/eLV4yuSPT7K/g+1SNaeH/Pu4aGkf6meBfEc9QibpztJaDKqMT7j0HoKQ8
RO2cQBfrAN7WI10fgmlRWuVbHCk4iFzuqmnTUjVrwcMi7zL2xnD2Xe4kFAMTttAb
ocUO/xgcpc04V59+MvdgfVdNY4+in6tUNKZijDlOh1Zxs3o8nqivBJAZVvQUnSKu
xcTgT6BxrxtgeX8lh5HlEQxH4X3ROpY/ZGRroTG7mTkjVOeFIGxEjES7A8WWCwfw
v7mXP2fBaoA+/SQVdQ44calQGQ8TK1Nh8HtkoKAbbvc4bYTeJIz4HdFKKZ5aoyum
OaV9Df4fKXI5lA9fC2C0XY7EqRiF9EMUMay21ZFtQDxRvvhlet9naa+6DYwfOSCD
AzCcQncx+Zg8BHZCdDGqRanh4WxpgLjQOoQQjBRqtt3pe1OM3krD/qJ0QQhLBvF2
pC4by7PXIEACUyTiYJyUmgl1h1L1bnLWbP7EhizX0fS7ndGTXtXYcjrUu5VK5FRS
tBn2qJ6qlRUQ7gDx+zvB8TezRgq3sCn42lheaEmVQqfC4fHBdf6TwuawEJfqlhoa
ndALjpqpQfvGH2lC0MqjpMGHjTsXZaTMPARavX1XIYHTis1KTKgIzHkjwPx2gCNg
i/8762sVT1C+LBZATX2w8z1izIDOmOHWFqv73eW5gKGL2fNYN8ywYFL1ZUfl2bJ0
GFFlp5kGxzYgN4lYLLdR8vDN+AggpIcQ5neybZ26Br2aM/fwMPaPiM+rIapGDkcx
VCEFJv7dTeJb7qPoxDziAsjBvqbHdBdvm7lk37IHS6egdH9OQqbSNrPL8Xdbhpda
q6YDXN9R23mUOnOOCRtFHE1VZifYvzKEo77urqqKHEaMcLDHzb7qRGMCPogCnPlN
bXFjRdTZ95Ii5/vlZBmuUJTH94rGAP0ouyeewtCQTFEgXrxKQfX0ezjmk2+Zoeeh
Zfy9Qhtk9fC3ZG7URoFXN/mh+hj/b0FPutGeyxxd1phsDe6IifGAaotCci58XVEq
NxLP6Eg+53OmIlSgr7aA9Ovxg1EhNJKXA1Hc8npdSLWo0LpBhNNE0UMTFtrx8c/r
fCCGSXwo/2ui+qIlOtwTNaqmDRLKPruKxCayrZ6X3E6JgLIwhlMDf+7paMcg/bWy
/edl9R3XRHljMtYO4Yw5Py0oqEOdL42EiJKVMxnpgVBZLKjapf2i6tEJSOns+UKU
QgLOCsuYeFLAIyr8/ZLbZ4wNvlwd0KAKiDXpb5+xYbeUPLZh+r7NEgGdnaDtKp7D
UPmZG2qspp0N+8t1Ipmf51+VbJvf8UF56IYzENMWQr82weABS9HHfNPdZ5V8SWFN
6LSVEH+R421wOIeCeH2XeQM/L684KnYx72//8EJr24RYac+n6B0D6YYartbbKX9z
58x+6alJKOU2Yny24aw45+q9fNiggjLYBTPjlNaXJ7ofDNHTiP+Jhk2BUFd5cdyS
TKq/R582FS+rXPSJMuwV610z8kOwicM6K2Pl6GtBhr+mmf22G7+eg93uixcLs8Lg
+kzc/O7u+PvWM419trY7vDldLH+1tmUg62w/kKc4xC6F49ym2Odl9emktqR26naV
B3ZDgKCRkz4Azym8+471ii3YPUQDmJisaGeCMthRuk/s3FJBjYlPuyNSDA/0+sYR
BXNqp0EVUpp1/NhywKFh4ZG8B9GKQMiw4r6fuSjF5iiAi+kJ+somkFEkfMw83V+T
6/hCmcPY42xVRjH8xXQcP6KH4Ado68E64RwaqpoeeXvU5q/DQ8BROaIkJmFFIuyx
0HC3AZdaSHPKzr7vuLUQB1T6PK8jRtKeG0eONoDjf8ooYev5KBwGXYnFuPzKlGe7
X0ExAO298WxhOqhnfneIFBftnXHkQcf5VLL7x4VNQ2yKSMhiZ/2sfXTE8XFU1cdO
wxHweNCfMb7FOJfVpw3wuxesAFWzhuuvvR6Jmx6jvar6MmOH7czC5CHvEBnIheMi
C2P1U386403IMJbqrAp2i/3uD1r8hkO/y7DpZVKZSMaoDdja4UKS3XIjwxGYV/kR
0PF1tDjovooYn7rC4jW4BJTS0V9AjyrDo498Hi6Xl6Y6ATXm+RUSBFf4m2FVIhsU
OvhhMezt5VKJDknm9TgpX4uWzqNukSsk0oO+V2/PgC43qRM8VL4y8voTVvmk9swm
e5Umbcn/wXNooOADs+9IctYjmLAiQLvxtwszvFyfMvTQKgUHxNcGVhu57Wx6ozCf
YwK1lCFZC6IOFmDdZUTIfvMtwbfwiyGZ5ItCofyWAh/MtdvsMqb9aTdgbS0ade6v
NyBpwJ3XhovcAehhKr6A8ofS0uFhL8YZapTHSz/mlTo2yCTzHGmXZVekuWol1VFo
b+xINIkxe6+Mjmb88gxjYq2sCoJ7dJ3gF5mGmnlJtZfHjFwIC/f0dq9s8gFusYRG
DtjPUinpQAsZ0GQ5Kb/IBQeDJp+AZB9MUYRVZ9xiznDgSRuNNQOdLdhw6LraKCYI
tiD76BlkFzBHdiiJGQAlAjddWCYEK3FVM0V5jkjAOpNtuRzZOaNHmUTHICL7JzL7
WxR2uyQKZ8OfLTBO27Bs7qwIrbBPwx1lE1/5mYxee9blqGxpSAunWaUSyV0hlEwK
VP9JJ/irEMvC6aHEnAMIh8x0T6Ak1IJKkAuidws7xJUJ07Bq4YwWZ4zg+nnkl1EP
ZSrqsFjzW3+7iw8pUfUNDIK38BJtenK4eZ+b5ytNHX/Kgj/c525BnZmLU3PYu6n2
SCjo7qGUrhEoyi7+fhB5Yta3Z5DKj40iax7bxFEV7eLk/hilERql+tJEJofUn66t
4rLc/kw3HR0sOe+ufC2Hbv8cxzc39/VeSHP6vXTUNdUwKHNUR5A9kXOOrmoPetdn
yfce2J+Soh3k6bLHb0pT6URcTe8Z/6k79bUxeoracIS6UjVC5JulN8jPlU6dX6Fj
GTzth006WFyYcwIPg5IgmsaUetwT64wwbNJH0BJtpKGtq3xhsjvk/zr2vTwYryOW
GJ0271ws7JBwPTBzXSCZlH/TJUoqqihxV1wOQvxVutY2ZqK28QydC0UcCHbQX5Ww
wzK6FT/fhfPDqbRF5QJA04w9xCO/h8RszT1MPwwy4TW/kXszTNbCRpatQ5h5nppg
OYlba0I7tueS79uEi3GOK5T7XaaSsnYbEbnFnNr6ctIQzoJjo1eSDtuOES75yAwq
q7ehGiPNRTaBN0hUjYx3DH53b7QK78px07XwcJz1sdOvibupCiww3jbGXKpyC1i/
9M48TmQVnzzcfDw6yTWDqHF8SIyjR4br6tvwlBKV8O2AMIgN62Q6xeghoIw+D0IC
z76FxavlnO2yUmJiwOVkCRcqBiWXBHvEY9/8FA4rPxg4C2HwBSr7ioMtAfGWlHXE
8yej1/bExirPq5/7UYjmQe9yxJv/RGEyHoXkwKtjCVtGjhIfkoNzh2qBzJItB6FL
eGdQGZX+YERQHmR3xSLH5pfDxyJoCIUqsFOJ2c/TXPXv6rx77oOPZgxUpalEsz5+
oS3JJHjTv1SJJecUJuZt/16DwieKcK4hNR8gBQEJwE27t/66J2GYRcRYTqHgSuLW
sL+q3I7NSLfrpEfYRBnLnQTQs4X3hi4wa+uYTjrTHK7whio00lyH+EHUGlqpNZDm
kifZq1iZ4uWPkSAF81DBKjO7uj+jPqlavx7qlcrJfaz2GeN1iLKupg1LbbqBVs5M
HBsTHMFlT0dtOPVyONIcMM3KQpSjdXGt4I2lgWEPiTMMfJE2g59CENIbAFQYv0OA
pg8VYlQYzhxL4HPxP7Y45wPdpXGFzb3pcmRc62xpjU6tSELgjWs3pR0FyQ1hnEXK
TmU9s75f4R+dH2zeXj2Oqg3n0OrgGG9QQyLmTLsQiHdUA0cuH6cvbd96LWw4nUZh
9AtHutwMMxWz/gf1Y4f3QewdBCQ11Boa30IWkvAk9SdcruYppviPKNtHqqQVIfIZ
nsx295Uh+ZhZuiKFYk3VcPmuNmaxljcgjvPctSWHy2Mt4mSbYD16R0rUy0Q3zHuS
0MVupRclzkpL6PB1semxJOdbEa5Q27xG8mNtafYmBnYzUt7hZgXmJ+WaqNcCiQYR
aIfWK510V+Sj3qTe7zwWjyRt7nueop0cvL5DxHiF6Q5nsx/s1TzEFs74Wgvg2HLq
xKEGVWEV1z05bZlSyAcePUZ6DflMcAR74d38gs2rMCIT8yp0iX9niYxnlqIpscC9
HeCqwv8kJUce488hXXP8XtdqDHUYeJhLoCIJG5ZQRuerL7BYItuNvZcvFWqJ+prM
VcGa5Qbv79Lm0A1K3UKQQz4b1plWwdAlCz0OUVGAuAdESCRi9tEgt7wX8e5edpON
33JvArRypwLSAa+qO26x71/aEJ5uxg6U2setJSNF0xgyvnUR5PmcWmxOQWaZaON+
OSmPtI1uySVRuQvmdLhQnmEiw0NKjpAuE0NWNRc1mf3k8Oq7N70fPXCDXc2AB+Xu
NeaQ0YflMFPbLrZX6ESQx3wV+e2RxaddlMgScKS6ln4anK4VzRsn4JoyPFkN3Vjz
yrtpw+ngvsccgX92IDp+vYEKjVj0iWk96dEpyjFCg7Ld2Afq5k3rDKJP08izd1KX
cbIP+pYBKt9p/DJwyCJa0w1LwGaPSK/fycIZp6KFNqv1Nmif9O9wrEjYTVdYD6D7
xla5wgMrlthbWQFgDe7XIeqIFXgk1r9oBhKMqL5UpuUQYjGebygQU2r+ufiIc7ff
AbJvOWWKORkIJjBRI4Z/uIaqlk8aw+FnFDgRa5F7/WsvWNBVUOnUeJHn0PKupyhY
yR51jkC2EB9wIyYQMtHg8wHmh+KDZPgosZaZbmJ1UUz71ASKF8KTYwJBg0iiNCD+
iH3qhcA/W6kJ1jsxzOpOuIkui/AihculuEd5SulbAc6F5L6n1TBuSPjJOxDsAICS
kA5uElAy+JHAPfKzLCsHsO/Qa4vsEj34kvC19gzKVxArcwkNWAEZ+OBD7cWJ/Bmt
qxY/kA8X6h9SdTLdb56rIURpzBY4CUhXnq78V8zeFxaCBQe+NX0ZhbIlxxw5vqdb
ndZlcmgYHhvCCT2Oi+bZpHobrWcOfYjF8jeofuCrr6WU9IIHeUthIFkl9pTZwBXW
MGlsPmwdujKzFMIeduXYyDINKoYwTuFshxYah8ckPzclN7dgwA9ylP611VjpzJjn
fZdjl1aTb1ZRTnKggYt3A2ruxvvBA+LEwLLC5KBfwdlwORM3BK+dN5HnwAKeaXqd
N7lyh8GTW9Z/AuwL6PgMLI6Iw/91A8FTWV58xpqTqapj+4D73lko7S+UA8CcTq8Z
6NisnQid0jBBPreq5Grg2fjsJy3WiKaAZQdgAn4I4+SIEZK35N2DIZiY3TD8YWs/
LDBF9CgaVr4IM9JSsVmRqbsbhalBgBQibHmmR/WSB6Qqab4bYP9qQ5b2or7+4EZW
/jLsohW2EXoP40ygv/1/BHRBSPloH7abyKfU/p3rj2aIpRJwoUe0lGwnrigJAFos
lL0Gc+fT/xa15cM6L4EMecT2v717l3u/LSy6JRP4Tv6kM9FG1gYnj4YUDBCLzPvF
Buae/Avzhumc+K0IFYfOKY1cR6X54UXF+VYoNQ0DNFcXILGzKNmj1/Q6grvQBtBC
Sx0t6UwEMd0241cx4ksZZByHFnxPb29DFvbUtRxr6euRtDsa1O7EhT9Snx4w6PAO
uXb1FrZKWL6LhX0tRQumPXTUFK24Sm4r5/W4npvRaqzbV5VmMUYWFVag0eWBlxeW
71A9Yo5LxgZBRUGSs5qw4m36n0v3rkyhBzWmCruW7pfpFvFgC0ivam2gNRXjD9i5
MaKoO2F1bnLMjZn/lULTYooack9Z5bdyZ0gYALUiafe2F7ZE5ElbHNz/I9GGNMo1
15AbzbzAplD1uV38GouXpcsOBiwRcbKKD5RcGRETv5T4WtBeaHAs8ir/FC8kgnZx
wGxIeQrP0GNBvgZOPq1DZe6qg7Pnngk2PVk+aGK931OeyvdMNAA1bxojoy5qdVEJ
yCE/KfRbm2K0ddaIl7i797Wv5gYxo9Ps6td59oZ0CL0jonqnh16Ivrsa7RbALOYy
FukSpbKvEvt1J3fNlLhozGoQ0iIEE0Q/vHo1slTnSskeS7q5SM6za8NHiD8/5dV+
m2LWigmaXnMP2HCSzngucCkTkuOpYgHNCutW7taDt6u5hyYQ4UD5mr4gyPwsBR2P
OmlVGjskC6dyGZ5PVkaFUY23Vkp8Jm+dJu9DjLdlbyoDg67s6XZlLYP92cAwkbvv
P8azaFiz/7dOspimjYEG8FaHXIF/ltFZqmFfQKZ3csYL3ArJh/HO9HRb56LHuIiS
beGCwccFtva55aMC1tdw9jODaJThM/LMzkjKY4yGZG3xcaqKkE0s2bm0aWiIt+e2
J6HUoABpvMQf4deBBmvUp1Wr4+T2AWGBdyCeqBsgvegWv5+hZvmWHysnT7GRAZAy
W5/nCT5UiDxSQW5tjyleKxxTUDWiBVDLTa8Kc8bXaGE3g5UO2ujjN7K1Vt3OpsAF
kABZUSJsBjsSjF4t2df15abzV7DPJgcicegCB+wgSCmsbQ8uVVtoJza4UTdeNmoQ
pk9YzkpYFLflDbFomug3BBn0BjAZZezycI4qXbi05JYyNMpgey27veGRX3I92Ne3
xyrx5THe49Pj2d943vO6QFkISKLjUMIJs5+LGGe0ncOJ/CqjYx06DY1/0AgTqjml
FJHqgDAU9/1w3sI6ksT283xhJdZaeZyr/+eeC26+qmTchEglUpqM0aui/9D2O0/N
/PX7rGtK74mW21tl4P/gzlcKScqqoF//NXQZ2elBq5vTNPz0m3Nhq1cYX1OPOXVH
NZ30FdVROTDDMb9atSwIUhXk0YIwXEfRB8x8GAbnmNgm1EOP1jySqr4w7Y7oDLud
yrRZGrt1PudfXaZCUUxCFBqs31kCmAU5SFi7RAc/haWhX64knZxxSSCFQS/LnKm4
UIMlk0BBvuxclnoTSNNshq/ep/G8WvjfvVP9Y+COZEYajW8HlSA1cqTIhqP+lzVw
ZtWQzUvhN+jJv5+D8xsZ/8u8/531S8yqVQy+2H7ww/ZhMmvz+xJqFWc21lokHRma
QOA94XgkpaCalRwsIMlFjPfr1oAW0Cd5XPc9v3DOY2guK6+Reoko3bHVhW3ONGZM
GaUGIExrdZXZaDQfoeMvhZ7uAaZ6ZnWZQkDkVu9gpov0wik5yCA2rVZs7BjOtACY
IC83CunwO5C63YbGMoOFFb9Z57Or/x8leWAhdZ7bJahJ91mCvPx5GNtADVYaFiTd
/LcIxg6iATu/RBvtpHohYNVhSHP/XMu/+e4xZK1v6rwIUSWYMReHNcwhvkEJqxY/
iRbyiblNTFSeeoJu4Cr0L4ZQRMx0MBHDMGd9XgHNi2E8CLceBHwfWR2MzNnlF4Ha
jYeIJDdBdXy2hZBHgujanQ1zMskfyk2PYs/l+cca3TDFVbMXKPqi+kk5QiF6kRX4
kL4fG2hBpW2+PKqtNIYPPoBEAT46tU6yt3baLRGjt3BnKoibuzGuE+fm0iU19y/i
Fj4umQeOl9CU5d9cy15StCqAEyfImedD3hZD+NYFs8bz8vqMdFFYdFjyXXZ8tJkH
a+Vyo0ybXbSnd3g0btc7YgwoYKVMg4GfcHky854rzbrKtdBIw0IxsO/kS4cVpn/A
s27DuQsN8Uhkanxr3zlP4ZRaxgfsjnczhN4g+Wcr8FUG0Yhkn4h9CTSNPVWIGwvF
mqA2fK3BxHuXQ5wco3M6aa28i7vjn0DR1HogE/Pw//CMkiwwXpkTVWeE8rnjWoKq
JUPNV/gaSAcKrDyxKFPHPUSaxEvTD4cJOsTnHXWl6/dQ9pem1/waUXYZMGzmqwp2
jqudy+QziPEvFAepxb8Kzx35ejFFlxKn04FO4IBewUvmv28b87iObNn80RNVX9fy
ZwClp2YkAgo464swnOh4C7mpFb2jZ+CKYvNhLRTk9/6/0JlFoiucs1w/AdqBhzpy
XKPXKdREDwUxeCZRIepiWNKOq3k6VXLeL4xCQFk/HjSf3Y3IMfEnLLdp7OGbn5iZ
FzDaCf/Go3o/3l6ZUQFwDLIMes3wUJjELDR4mcp+UApjyyMXV0AISMZ15TMLAD8p
/i/oY7Jw68kfosaZhcRej3fIxQath9awUnGA+NX3nKMDNzAyVTpsnnzXT2CQ5UF5
onzUMT8facJpI7hIn7anr/KQQDrJnGhZTltPfAGzhJaz3Gv0T6O5EnR1bXeeny2Z
5xH7JNM/O0a4B9h9BXUY+GmU7iYQPDjhZQ32X3b1xk/RRFgTWnUKnH8TlA3W2BrY
GHE4IwKxwv//9JNMwUXdHLEswBoe4ReBgGXY5d2s5VcHSIkH4sLZ+kIc39M6Lmn0
o/zpTbdR9Sur4yLmOJAobjqsi3zdr9KXPDscOj1d6uryg/0Az2uFMqdA0XMZ/SbQ
C+zuR1j3mm6WSATuw6r8e3f/M5z9WhudLVK/JoigheqU+fuX5ESQJ25oWbs4TbIF
UpFaJ5Mkcs16N1QCcXy3GWgWv5MaTnLD1vsVqPI1GIUiTxg03m0W8XEgPAyoV5qS
Gb+XX5ZW6D3JtmaZU1ChMbNKtTMdhQDRTwEWUGj5t2P3cRD53ITvlafFy5nAA1b7
nrGIlJ47Wz2uMqIhAo7jmpZ5hoSuIYB0PoFDsMjM84ICP359g3WjKCsBVMXxDaeY
e2RTrKGqJQS+pljDKYPkkatZnn3s0yH6g3Hy6QPG5DABOG8mmG+x8mvmEmWg79uM
WulKgGcMsWIrzHtfPuuEWySMyiyLxwLKzfkz6KJaJnfGhumASbYfGUdPglhezhHS
bBnSmwvr+zV90HLPaa5+o+++06kpJA0LQtq5vrIdgrGTH2pmmsYo66aBtUkgkBNS
0cRqktztoVQxCafWlFOrpqUQpFq93UHgATQNBG1P4sUOtdomp86TaU6XVoUsh4jI
6f9OXERTL4tzPfl6M3eE6m47ECCdKdCmWCxTu/MNYRxtmdKx8ZXm0/20b/i2+Fhq
Lw/3V5CBf6bba9bHha2yT82ENjTFbCdxSw1cvYtoo7muJO9RTkXXIQW4al8aYUFG
1HepzC4nbr470VT80Wqiu85GJDA31ka9ao34GMT/aDf2J6Oqv5yOZnTQnNW7GqtM
NEEra4ZlXOu87MkZWNckPL2LcLTXvrua6VWampLBwIrxeXVvCYWQ7OLvVsvgUjmS
pU9941F7nV5t/yrZp4GNx1pViUtMHxsXQRiPWDcoRKG0HP2NzeiEK9U34DnbGlsg
oZj+Yn41NOJGcMiJoRZoxRbWuQyUTIp8eAp4KelZj4XwmJOYU22MftFnufN0C3y2
hF4BZ6tJ/kxehiNqE9aIgPl8pjwEMT//Vy/y1KEEY/e3fLEpGEYOes+WnSgohTAg
NDLQrey3E5pwlhjuETpLJ5fquiXwcvOOev+mNE0D+RJnTwlNRn8DdbyPLMqBiZmS
qcaLvNrtjchoRAs76M3j72lzL1f8eNXVrDTQfe22MNX86+z3tuoIYYQPHivq3G/h
nPIRdoeuAtM4LdlpQt7L+tWWMoPzgPGtuMDOs7IlCIVRS7fkCdzhtptTOfn1fiQS
zV1AbYRdg5pwoui4/B+RZa6akZIxKV1ki/XV0II9/ZW3C+OU4RZ4VgbRdEVSIYJx
pNxOEASONR111xsl1mOiCtMIazkuBP+gqrNqvF0hIa9ctlcRnQbcREFIOwOvSjRL
N5kMQyQW3ikDUlACG4ZQ06PVvYyZRZCnj6ZxITL3zwJOYXF6nooimyGgpqYFl8B4
AJyHcxFREinB9ypWkrI5UZUrRM1HOqgUSyNgqar/q+glsScBcOU3bmVbwl3lmUML
7AqX89M5CZIA6dz7Lx+lvUEM/LY/XmLkfqQb6vP+MBTzXY9cfwkqxCMYg9wQ1DwC
fKP6hQSBCs+WMLolfMYyYwAor4lDHIYCmbjl2BK3znIh9KWv68/sSPmY95cLTc59
IPHMhlis3sHL19FtELS9MHFqVfcy2LvWXpJ41ssRRtsvrUVWd1gUO2otv9dDG1rV
lWuzMwFVjxDRx0/B8fHdRH7DRUO91yY3iixntTUSDG6KsSnSuzJ0asUSjUJ4TSk0
jIngPgaH/11WVvYVlECbjl456rXyGA59u4VIQfgybLWNLzh8zUQACNF/69lGytnT
XzxNGxNoSQasvuECO0GUHm6Aa3LQjT9sNqdL0CM1YzNCXCE5nrE5HDUNRE6B2UcW
OwkNtkXDVkJpROwopu2JO3D0bxumN/G4C4h7ruK3eT/efFQSwGScILSl5pzev53L
VLzAMZ6mqHUTifSO8NjkHwI6lS345MeesOs0XFxpjwAmDG+QN94hh8E0r4hZZVT/
OLC5Md4QXE8fcwt1Ka3DXYoU20OCOAxkINR/b4ubZO4zTxNdd4U/5VxrEVZCZdci
9m5rPg37sa9a9/gXVfICvpMKHTNTXAJztoIO1eXpddQHsa7JZrfyGkpExA631w8h
6InRe3jEs7AV9C1JrFR5EhNbmIdXTjuKNTnzJrjFl9c18OgSDrskkhSvTxBkK9bD
+BRMdTzA9MVjK9BTbRbyjoCNMlQYwfqMRGBbNptbg1EP54O8aTEC7jHwOtOUgBm7
fkexMbL3r8Evu93ptQ6iWur4DoHBCBb5RsKo2Wvmt1gE+YflIKwwEp9NrTkxzWB0
Fp88iLuXLqeQ10js8wD+64Dstuh60TkGW0BIueqDozxCaYnLsC6M5XzNz3pR3b1j
FNO6wLZAMa/P0+T/hU1M5trpeX7rD3ALQzDCZ0KwDvHE7ApE6Gd2Ikdx4m5UbLan
g2TgLArZVJu7LT27zy3hR9uwF5UxeX8taTIavlzoe+oeSGv2/KRoEp4o/StUJSzF
VYqwRfT7grV8ap2Q4deE8RlCeRIMSSP5sCR5RYVlWwFWb6f66bt06unLri7CcPBW
ePxhE5Z8NishriG+FsrbnlJR7P00m0yX3BzVmB5MWrZjWpQTZhAvXUd/ZK7UJda6
RPaexPCeDKrEhD41/rlC52UrLEhdGvV8qz5wZfYk+YqDkc+C80V9KnpPWXkId/Pt
lfYFgKrNEka1usOyZozZrucqXJzzXRrfUl7iaFIe6RuIBCwyh26c3//D4dP8R67V
ObgThLxWpdcEFOWzsKn4icBcOTz9GA8ytc7n3E5GriGBbLrUg0/P/ksB7Dcwolkq
JIiwkxxiX1mqElG000n9H5BxcQ4L7INJG9S/0qPzapR93in8TXP1Ul+5jbi/mlr3
ErwmP2uKIkRhUT/VwHK5Pyf3n1LhHBVd86jTzpwe3/7p4PPvmRBN9lr8CdkbdRm0
+dYA3UUkxs4IY7QjKN0bTUjdmMB7XtFlYBbLBrIkP9EfUWzURefgrywGp9x9dhWq
8QcvLAAD3K0Zsis+uRNAFZ2FqU7u48v53kIyCqKV6Z6nPMp1Ps4aaxb+IDNx54O+
f5cuH6cUav68QEQogzNpE44/hHX7OrfEp9s+rt/U/WbthxPyEybOaugCxuwzK6pd
r75XJkRlfpVyHhAYtyI0POnEOlHuv1mar5IuM2J0Lnshgm1h7zhVb/u0TXC5ivrs
8oCOnnCYqldQhvlq/B1WyAh0e7c+zHrDVtBjq2C7a85e9yGcG6JzAHvQHspuHd7x
E6juuIuG0EmuqRs84pEFBEPtEzHU4285AvyDriGg8ONiQs31reppAVRpM/2A0v4s
m1Eg7Mp4RmswQK9JUS7OdM2sklgY0sEVRefCiLdXnjBWapjViwj3Y6lET5kBmhdS
YqMQvB1c7aXhnXxjM5tFVFiUlY/s/tmUNXHoin2ZACwsYVKPiFMQoLmZn9sNQvih
xXY7Vj0wdteqaWLNCiC0CoNpbv9TTnZ6BHTdguh8B/PUBE7j2rQP/4tB0ZiddznU
r0n2s63TApsmJ1NBX3DrgeaaWFQSuiLzUAb/XTVlBTofBhdcpUcvWDvlsj/Hv9jd
w7sDv+89z3fe8i0vB7IM4N7mksGpNovIdfSsX8YI9/hlIlnm1jhtylE8Y7BNXDI6
hxeoCoGZ7jo9CmCuVUAs+g85+TgflFa4fBD+ZBPv2A7WRn5Gdw09PLqn1RStXPoU
FIoXQe0A9m2mwYE55Hf8zg7kwrWkgfc11UGz9AjJXsb0a4I6PI0enhFQNiFxT48e
+CpZi6EZuC2sxSs0YINnPJi1zVtz9oSRzGtMS6jML6uOfXixbjMOBHoqamqNlJOA
ZPuUN0bksRa/Nsqe8bMF/atigndrhJ2gqq9FpeVb+HouhFJx0jpCdFi46/A9K6Rq
ywdp6JYm5FyMZh2dXOhpy/fiRZzQWeNEwF9M+e6JoTrq0/YM2Zwf8NwpjEQpFiUs
9LACPBczgoL4vu9gSrmhbovgAe8a8P9/9V4AcdkypogJVbqMc+j4KRI900307nwU
cAIIS/ApHqRm4zAfXUnW+76FWRIwPkd59iBzXy4OK3C3voP02ndQ5jv+17JnuEuR
QVwvE2OJmG62gNC+WLBtfP1/5jMFHRZPYfMzio4CIVsjZ/bkEH2kRnjYu2zzYDqV
5ZC4vj7cbqEOg1sKdq+//fDubnFUiHlB13MVxPBuxuohIpklJT8upHo8hozBJA9j
wU7ESIN5RRq5guM/CgUzc78TK/rQuHPMDXD8A7RQaTJCY9WIbIDmwBMuFGbtIZdQ
ajxJqev4aMv/o3S5avlKlRtdPoMg9ms8mVbvfZ5kwAMbZu8qyZSLFrznkRkSmIuZ
wvtYxpx5ZjY5k1tA6UCkmlbso+cEMsHff7jr2ERYZ4JlbuCihQWjXsfAJJ1UbXqs
lz9VA7jsm5uB9RmWy8w3vrwIiF1W2gtwW+VRlu3Xu1dNkuZbtqAPwptXmbSfHLZ/
nmDn3OOpFND3m7lmCq+EwR6p+xKIPoGrIUdlTcbgE/FPJOtvbiY8fKWslxQdGSYA
lQuizHeyqbWVDreZeptQ/d8Sla8Ob+Tf+p/iBEy29rSenGXOI3a5GHS8sX+Hh+A7
AiRdy42cKOsfUevZJuGjYN56AxGYyzajxNBg1MEHIix60f4mf74GW8KqJdG4U/zf
aS6TJJsWeKMuRCT8jgFH0F+uC3Ky6UAeT2GTzr7WVPf/XUBFdNt0iyBERmkPzVbI
mnTAir4FGSQvyWhs9Dx3wu+O8G+x0Z9cic4yzquZJ3za6en2xIhzyo5u23OAAPuq
GODYAwl65RbsMpfepMu1bgUqQqQSpLQrjG4F1zJWxOwvwC6Z/rb7d+udCLNj/PhB
DHLqJ93ABYH2a+1cjtFViHd3jg4ITwSLtkyfSrpuwvOR0Qye6ow/l1DDzvDR7HF/
/IM89gqQQdTxmufeAtLoFqQkia0PIrFUs07onRKs6lky4lnOr8sK2a4OCz5Xl841
eiYW4R1J+GrKFfHXRDE/rre0TGbnaPYgyY7DJVyM9/Vt64f3AA+QKVYKN2YBMZoB
/NGa1xlvhfoMJ13HfmpprcsPl2KkCVYiI5ouT1FKboAEOWUO/7eP7hgB7Nl6AAl7
u5v7SYbFmnfJLQocPrbls56Fei1t9a8XJ+tjNLzsV3wSPkAIwwSdz1NWI4xc6Eit
S/R6EIlCvq0SQW0/4nfObpVH0GkWOtxU5K6eWDF34ecH6/sBvtcM6hpyNUgZgCxP
bGZdrLtnfmGbbCAiPEuYBWFa7nKxtRR+FS/8DhCT9/nttHJF5ryQU6/cp3rnSiOv
8C4JCgvh2VP66rJSN6pnbtaiBFqLoMIbJGhOTYbbQsRNXTBEWX3XRgNbRoWz1P8C
Dr7j6Zr0UIwCHbEs4pr4MMy/ZtjOxmhQ2+B+caTjVNBgEpKfpuvke80Ha6hfIBqM
RlnPKKefaNcZ5qUfqVUTfAW+/VyXlvQeUys7BxHG9gEflUMiYLn8SM5p1nUuVvLL
sI58jyrUfH4fnUPz9K/wOPGjWbF6keo1BHJymv7GvjPa+scKqboYnucgMHGARWha
e/yulFS6nbMJuwcVp0LIm98teQTPNMMHrY9zkvQWxVlS7pmCKVkegosrz2bDkJ4f
L9OeuGK1S8pdwkWJKrEGN70yJ3xcpfJEsD/wif1LJ+6kcTCtHMo7nXxsIktz2Rha
KyjPZfWrD6Rpcv4XLvIGOx3eGR/fr5MipVrkwKzY6RcNP5FfBHgscdP+KGASOUUS
juHubT2J3ptQkaO9b4XJYDGp/oDnJzinbg0t4TXLUS6lrLETTzFH8XBeJ0xz9SAP
JOW6u6QdJYoLUCOP/Yzx+jGiPSUm7tu04eMMtXUiGH1G5tvayBNMA5isVAIw8Dz/
GFOgLfA8kIekQRAIq9nKgoMw/+g3bNDqbkle7igpqvcaXbQM05EhbSULyhYyh8gG
Od2VkHcQ69JtrMCJu1pQFUpNWz5UYcgomvhXBUgIno/+ixzb92ZKR80OE74irpsE
8sp/77mlJCcXAWVJudApq1pmBbEW9zzX1e7a4c10lYwzD8L61UommY2A/JPK84e3
L+TDlXprK9ZVJzaSGA+D2iThDzDxQKgr2lZYpZ7JAuCXeXmeynrqoLh6/eH7F251
32272ykvLTFeKNbI6Tj3z+iht1hb2i7IOc1bzFHiE3ubh3UzQxdL05f5JppEPKIz
GKv5WwX//xjsoMxUgFXEtzG4AD76TiLpnW/CnLlUAeZyw9HDVQqUSVSPhnk0JVxc
e8UfOwq7ASRPblrq+8TGf+pKV4+wbaNsltSlBhfoM+K+iJM7JUs5vZ/xXUvIK8xd
VTRZbhIahOlJjSelhI+Vis1UeTGKhnkBh6aiYdDMbpAHJaY4FfUkdayJQwZ56pGR
aTPr0OIQslArYus3XBT3Pgai7SAX6j4qU7Je2JqqimmOY7r9KYdd2n7Ww7tRLb/Z
iUnmeKsl/KV3DQq0pVH1s3h5+g28Ze0rpv1LfVGtOHr042NeEoubbJqFgjEliZzU
CVwYihY2WNTu4BSJAS5UDF7i1+0ZfL3pXvjcRAsOuolPHEKC3Fo9Hp7oV0yx7mwC
S2GzC1bQmXsiJnu19UHXFZSIB02fTOjgEstdOARy6kkLaQBzs2on0ECL4TXP6vPY
jo4LRTnAPJqDnEwf+vHnxoQ50OoJwpzeS17piq5/C7xXoMOdPvb9vJf36NT77/xN
jl+59wz0zCtI5vDZjNXPEfwb1jxct0geKr1siCA6cBrcUlbq2p1PGFSx01dBUSet
U74MWYK125/DPXZHfBnC6MtXq0ZOtHDFKZeNaJk1bPmYcuWlgL40CxFkoukH3agP
vFhXSL5gTMDQyPBYtSSuBdHud2LpN3RgFvSQj7V8ynWUNy8Bq/8l/f3aDOrp0Lcn
9JhKFMQxOVryT1BeyVYDfVZps4RyexaffI1TJralG+tlGzBahd9mQxUaVduX23HZ
HKLekmydipUVAh9H6a+YI+A5rTbyofAyMJlbzzfNfhu9e+daMQdo8lec02+f7T2H
zaigpkeVzDT5G91uiktOzM3jiBb08sT06OrBooGG9hVQhsIzAJxZJ69RV2vLcpyZ
IW234T/bAaQWNp16i8TM6qNCrJOJOzCzEvAOD+JPp0RTKLtjb2NXZMmvzNHR+nY2
LsHIlHYKZfxBqssanLsTgnm4QSbAaDaOu8u249ul/REc3LeZdCsMB3nr2rbHcZ+Z
8A9Iw9pWWD9jEey9qFAxToNij66D+izP6hfv44fxRzz2Zu+z5ISeOfJlvlAwZujz
0P8gNpXdEVdVpi93gIxdr0sdtmIegaUHBLSmu0eByWowACj+MPYOStCL31A+f5mZ
R7nvQ1GIsis5FzuLFr7h1W+49v/56hWOXdDp4N+TCu3tWXegRbtEboJC1/nSeecN
Bv/Hb0q00XE8YyVICekzG7y33zDtRIRxWPxM3D5KAiGSy/tLf1aUctmcc8VTqzrg
nRFSSvYyj3wMoZVQxmt1o1S2XJM2usxMWLZQt9WS2MOzMUwMAQA2fnsKf0RYM6jo
GNEFxMTmVElah0OeripFFFXzIVLYwGytY9LrQBGI9/mPLkMbacUlY8592mOLJ8b1
FS2Nfm1yr3EqkdEbJcoearSqUbiJjGca4XOOVUw8XbZAxQu1W1jsQrmpBiNR9SMJ
U2BQdoGeOweCsEkFMnmGO0KmqIPX/ys7ofcScUaQyQH3Gs3UQMt2AgjIrMUm6FS4
FYUvHsSXKj8Q/14ovDfayQhC4ylzBGQSSi/4tcbitpYn/+cuXANpZZzQPIkvZAS+
2AvN96kbooeocsP0edvZvmdrrG/XOJ2X3achY/5wvcElF+75+Yf3h3YKoG7Sz5cz
D4N/TCsF6E1Fl71iQRAcWHM2IpRXgd3zt5dEYl2A699RC8zkALKsqpoL44b6jhkn
AYhUD/CB1P6kytfncT++ETCJjCzfsPolrMPIbjZelNjr+X/0P43w4+Qu3btviLF4
p4LH/Zimi2Mhq3n8HFhFPtOu3W5o/HTTrj/naIuW09QUolVSzzKJEiLzApIsu//D
DscLBKJ9f2htPftyv/hmfQqdmr5W/svI+L++fw5LAlnCKVdvpMUiKUFQiqYiR3O8
Iuq7JBclCExkuLRt/WGDUWiq8BHjbYifT5y3n8/vLxBZIiHxLbHT/UpQkVvWTQLM
IcH7PabEzXBVziWX05Krz3tAwuJN8F7yC66bKLVjDNCwaFJc7QDPB+dkTh3+Ble1
Fih7JZTXlvDNz5Pxcuk/Pg9VhHTAggu+38yVrYL8p+y1NBzHj8fdib5ZLlAaGRdF
z8/Jx9+9XG/CNmUVNeKF6nwczuj5iA9tC4vOVpKWKEeWD166Zu5VlpuFM5Nm0rVj
syI+HOqQBEdJ1py9Mi/HdrqlzZknwhckmrzpb99eFkGDWUHyK5+rv2K8wNlzR3u8
eFR+u/fN6gUTLMBKKK2PrUe0XlY4cQzYzfTp7n7mMNhLqu1pr+glBdOCW3zRhGxu
n5omdVBb+flNNGNBbnbqWo+3bm12kh50LsGTFGcCj81ss7AU4ZAj6hPGxc5Jz7Hp
HMbyOOTRnF20o9Yo7JbZg2iEgo2OB+2HFlGWwGqmf5h9+m+1giBbC77Mgzm0/vYI
Gt5KOGUYKghwobVPvn9V+zUZrm5AQHe4XWbb+TYpPVsY6hVzTM4Z3EcGza+DOOkJ
KQKOTXDNiQh7JG+hSElC+uw6lf4DUVssgrCOjhojiJEI9qbdFhyQwmnhYVTdEFZi
GUIsfYvO3B+uf4u/3CLxyK1512n0v0Bt822Ch0AcD1Yk2/fjc9FX69G4Rv5l3QPE
LGFsCqq1oVa3BtEQTg5ODCiRjNgyyfV+A3aw4FZhOCSZPc9xxZ7vMGClaAB5OaAx
Rs0ayDRXEVQQkIJbSzyCzJuKbNFjIwpSu0HQoDcXTjHLha02E7AYU1sdPAqfvqoP
g+50U+akfzdGhAbPZj/hTAFZ0zoSZzd8t2mgCB51XbbrEIr0WZpDlI4L6djaYfWU
R0rwpIumPS9Qb60t9Og5aPLYRiR3P2PkPZQob4glRW+u7K7tj/SO5WfxesyzhDTx
w0g/7x3GHbLF+MXl3ulStLNWsFqAKE1aETs14eZR8eqHXzrbKjuOregajbKch3iM
IZlflnLeBhXcwVp3Urx8gRUGreTxkkdSPCO6i0Eu8qzJkondYYKBBkAht60ZKuaN
a6tXm2F7r65rLsukbd5m/hdnddWgGYK25aHMbBZadNLYLe72sLpbW6swoG9cBBLY
chYM+LVHvO+9nHeFlW1mQ3dm0fdpGRhYZUo2wb6GLApFWjjrSCYccrgVmFUyvM/C
ilrSW+qj7XkmGiYVw/RoSLXUDSYk9PLOiofb5r9Z6mk+deavv5lbw8HmQgxWkqRl
URrhkDti5q4HZILJyELp2Ms9Mc6GtZdO9PJoCVxGZFqTAA0b6fzz93Qlvsv+RfzJ
Ff2/gG6ZeKiElrt8aMyzEnO92sXtT5bfvj/yYFU/3u4rgYnSblyRqclM4d50rA9M
eoboQuZwnJqcck4YNpPEsL05Sg00epijIjM3rGxs/8oYX0+bHRVUA51Us7aiuxTH
AGE8mk16caYFfA1QDXUJy0u1CWvs8yF0iLtTCbwH0UHrDmw06LuE4Vd76seSuyvd
QVlua/IF0ZgBuSWiSGPfX5rS6kzNQGz9nyWGV3GnG72w2YJXOuL1IQqvzbEaF5oq
yNyddd1wJSv9ndRXEEKNEXe/A1k6L76ZifBw+cc86chM7LqJeZ466JKDXmwP1RtS
+NT5PZ3adCl9FbbwKWqEC2tzv195rJP80svQCnN0ZDLUjjZLMYIQ1YAeAgpeSAyi
GXHiyLDcXLwJtTI0LVA0M6kslkYSydQQw0qSk1bnG99yEiWxQgw2S4WHS0pXGTCO
zp+QEhmYzm6TSLkuwYLP/vaKb21piw2giSTShfhHDZrzDn3d9vRtDqImGF6sicbw
52qMuCuwzO7Km+BBsJ+0ExT596B/89ZWo07eLkvYqvirRv2pO5gDwTytu6ixwo8a
YO48SCj6g8hFEF89MnqG23+DH0kD7mwNhsFH9IjdkoXCfzpONSycn8i7uuEU6GQd
VyaCTREN8bqJorpH26eofNU0oTd9AuIN3mAdewYoFhgI+KHUAnmqDS/OjS+EhKaT
cWbFMTnC2gY8//6flRu+xsQn00jyS6zZqoXW4grMxXT1BECp2htfAiHPsaZZT65k
OVi3LXaHF4J41VqQ7fLlfwd/okYb5Zvn9tbHR+RRPGqetEUzCqjYMw5BTrx7OSch
ooo7R7bD8w0x72XpUTJ3VJYC94qQ8dPpvNlMQLVe78aa55PSBe4V7525XsvdpR4O
nlhv/QBkOfTFtTC2MvKZZFf73bmcel+8fsjQJ6us9rhv3lvJhKkB9PqwObJtwNfA
Zs27xgjZaGYgPnsAegb1QQGFjmUOZ1X1EoXpRJttiZl9Km6HjdjH5J7DeXQ3Y1SZ
Qyy7rPO5ocacViY1eadePLVT9JBKpc7/B5DZy19vD4kqpeNPhEXhsGPX6a6GHxqK
TowrNyvSWtrTpVa/xzX21bEnbHxGbvkj4zXzwyonaxPZ4A8b9trmGoD8hPOSdsqK
rH5ubxsVkocQd5PaTl/1fYi8xjDcY2Bl/r47ogqLtc7kvYaiFdl9crkKrFas3awW
SydUhrAI2Ta2pzln1CvQYLMzrNClZsbYeDBendMbZodpJdwd/pqa2mzIeFbEPy83
i2KyCxPs9HZdhrIUkJPleJAoD4qMW0V7j0MbgdJTatm9qNwNWHat968R/ltPSnV+
9j/yisnha4myCixwCCRZCLSrcR0JKzGdFQBuPAsS5lTRV+AqRSFxc98rw29l4jxY
gFgmUT359LyPiMC6FS82Pz50F7IQ6DB67THqNLWScS4GKkAql1gwijVlXm5gxroC
hwIR7yxQLH5TrbOI5XQAXg33j8jCl8yuzonQ4cFQcaWNMdYRDX4xhuHSUDpUNv5I
PjTexbGXodiyYoUhWx8Zo7DN6kT63rKmdKIEW55D9/Yneb5MgeA2ULH4TGJpATrj
IEMwz4lXlJcO8kb6HIaLriRzWqzAe/C+14qBY2dDcBmWa67OFnjpkpqgvFrYK788
lQ4OckRaG7J1cJreQZp7OcDMpAD1Ttdyg/q7ZhEH6qQsIVK8JYXUQtvrBqyjHvIN
6E8ZDTWC7U9aJ+ITd+NCNHdUHC6CyjPeKST88tWzVLZw0CL/VR2amfEEh5UsWmP9
29vkVifiow/biX50uHarWRk5LrpRiTYzZKdXSpzGUFHBViXMj2NvFTPLkduPwrvn
OMtWVjqNTwRuzFSuagc74KIkbddup0Mta/Z4sN+iNU5bq44xoYNRAta+ERcg3ARz
XXzYnWzYfJYFwY5hMXrUEy5AEhWFMwxdk+D/Ea08ykk7HBUNcm5imhpLAnT/pAdn
mKth6RVtrslvZkfzFPr6gJAddL/6UpUDFW0Kl6r8gbi4gNRwSA53ESrNJcMqr37t
yiQ3GENpkskFhIvNPbeH+vyot067Rl58CWcK9AnRqfYlhG/c5j11m5Gqh6J1Tjeo
daJMb7249V9nx16ohTpJEylfa2mfkBBvVvnIAx+TFvqgascKIN6spyNcUTLnZ2Io
hor6n1EzTJUmDVIqeTi1pWMeCf8A9ndwHwFH5Bz6NJ3oNipg9W8/xlU+8OamG6u2
JwNdetYd1Ol3WPGYSiTGG/0QAmJyNCcHLZ9DhLVhqI9D/zar96WANBNTMYHGVGQO
39ovPBnCGcCOnTmR1Osc8fMih+ErEddF2hlB2vxwA6biZDwjAKrGX6bobZJVQP00
7fuclsx4IzVImFyfgxDpQz6qxcBbWMVHzobYL+VN5F/BVsWBwIM7UBuKPN+cKgLV
lecZE4UehR2K8a7Dhc9X/3aft5lRW45nW8hXPruYal+lXdn0+1BO+GkLk47IzDGC
lsc7HVIz3/+Bk6SrnrhFaAbfvhw8AvsiKfx1mYbONtZFHCUnQioRvRatz+6GnjeX
GiH6nxx9dlqM0dsGvgWCRw5egWy9fLr0UA7N1b3306edzhNqdWpquZ0LcCM30diw
A1AcN7egOewjp9QKjbH9BOm/OVqS1wPfza37GPOJ8E4QLT4EHNnvR/ESgkWp3GYK
9gRHNTfrnotZfWzGy5K7Ej+0U84Np9V1b7TcK8BudKSIGTsAobwtN93zKWa5nYJG
yD12sGf0w3N7I1pV/exJhH5iHHW0OHzcd6AdHJZHjM7xgg3v/KhhCQ0ka8E0sUAA
A0wjxM3neTrqLvPI49q57JCxEaLxKU7QZlv/hfmY9ieClXi8FZyJKro/x1iklV8t
8fELZr/LYUnXOvPbSvuVBSZ8BBxnDWdIN7ToaK7Y3buJonpWd51kpVdn0CSsirwI
QC6H38iNX7yjZgqPzfo+voWxR2DogP3qeOtdeufx85MK3Maq6DA4rD8kuOmw3XWZ
JqENUyrwuZflj7dp6Z7hN9B9hX31iCRiCikTxTotWQ7mZ1MEIpHayTsUB+3UdGo1
HjqoLR+39iwwtSW0RCP6tFlRduJWxaIgAWonmHESorcvRqJp1sWZ0BgcX/0EjoS/
U0bgBhB0bIZaJvSr4Z1TAh0sdzCxEA2vei5llzewPNNo1HIkSGuZNfhQ54LWrP1k
HnuF3NiMZDqZ0KjP7B5X3Zj60Dc8Mztiv9gJkWtyR2Q7Qpp2td3n6QJg8D6g45zh
V3sirEqBreqN69oYSJjwtCUsGNdQlD/zSPrGW4+4qcXn9i1mhrEoFeZLSWVmjvKf
BvUTAMFkS8oYBj+duHm8yHaozWuYe2rbi3L+aM9XmTy9yFeHyPSCqn2ffZzmMFuU
vPAgGnoP4ljuHJ+os7dE+r4WE6JEogGbljvrCtW+10S/yw9Ks6qnq3+i48rAqBbz
HDwhpwwGnWmQ7+yhQuhTwbL0fTTVS4afQXYTmJ7D7yFCFcppaA1Hl5ErqfQ/H+iI
eNM0erZYA4JWwxVILOUOBJU280Q1qLlS/AJQEjkx594VpAQsG+d0BBFyyoH1dODl
BfsRo1c6KoYOyfTOwrtq6aLhwA3PH60/ANeJ8tysF8gZ4RYtpgPamsloZla+4mql
K2GKYEU/pHcpyDBfMfj2KdR8HnbbXwfbqHusvIEkuOvR2SQnIBUb91sXvwRKrA3R
VxYWoQ0FeFy91qv2wqEdec6KMGT91z9/QjA0+YyCW63vmT8vJPSC9Omw9rRL6110
YC7RDVNM/Zi+kwIQpaAmgOTDAOQ61YaGt7IPi4sPwAJfVaK5BXSL2TreYPTPWY4Q
bg5PoEctvcfRsrGQmxO18dhs7sygBlgm7JRM9CiIO21eAh7kddpLAEfr/NxEHLyV
DogJK/6DJaULeoXa0Hy/lJs/88HQXrbhR/QrY3mV3u5oHUMoFEx1w4evozLrcgaY
58PREXcqBEhfNHwSU23F1AQqnjP6b5uwzqSD0E4D15mnxQ4UJJfhy91B+YtSK+qV
PEMZDYOElzo7hM5RaIxHjyfUvV4rSoY99IT1cpzF5wOYg4S1bVTSWJXjPakAx7U8
U/ohxVoXUQrb6U6BZJImRzkcyp2vgdnFrktT5mHkNYh7nry2WJ4vEaBB2a4jnuw0
fJ6t1WRhmh26WS8a1mF4upO9BkQ8T7oRAkgjjRFfu2d6l7j2gWgNrxJZy8c3RtCr
ckRTlXIi6CaBseu4ghfDZcO37ds0AuEa6IKKW9j1+nJkKAoGPuwHRWGb7dp6+GoL
oNF9FhuJo/IsD4ptUCTQUaeX9gfcaI/5Jnt0U8pO5Qc6/E/mjj1HSMkA9ZPyvEUQ
EM4kWXvvczCJXqADCbwpSfdOqeTohuw+08pwgJgPR9D0uUtFqbENvxEHeb2kn3xR
IA1sa+eBhe+17vrILZpApV4Fl4vIlVPqr1YQeQLoI0yk9g+lR3SUfvVHgN+FQB7z
w2sc8/PHmCb19G8NGDPPbnQ74lCYFE3x9fkQ6PQPCEfKIoumucxebXe9ASUVcquy
yQD+xUGFXY/SR9X88GoFTpKTxrnoyhWIkEJBpoh+Q7BdVUfPgCCXjst2epVzwG2E
M1n4f0AmAEmhQKJHqhYLse05zf65QFyDWiq3tzL9yrB947ySVuYrYKnT3eG33mAA
vM7eM3lb/PlO11G+O+0Cg1ishu4Koei7FQnnXKn+vyz9AWXLLgQqWM02Y3N3YDPY
PRx1SsuFa95cKzkUJWbc68DbPlohL3rHqlz5FNqa3ZdN25XNrTGYFWEmpGRqEkey
3C7+OG8g0cwepxU3hj/+3Wl4u0CMkPFuxikVaJ+okME3kmlphIzI7BpPdIm2+sWS
l/wzwPBs1OWXkQdus0IBbCn6DkaqUk2Y4QyV8ytcjm9TgP5YDwc+IcoDgjYkwPNN
L+SvmxhoXHShrh+LobDVfVN7jBMj4mXwgF8CayJUdQtFNtwfckq+mk9X3TKXXALe
vnaBKCBx18fovp2WZ55nyCon0QjoIE/YmLj5Q03M+irO3M/WD/fqxpu41nHTFGh1
Kw7vr0ndaGiqoqOs5uvdcuKqy0QvNqAzwmen1+zo4hItXxD6jfLI4YFDQ3hV/pp3
74wvNToCZBotbdibFi6sZLvkVj8RAE7pi63RnBOSr9sJEaL7Vsms/yXKssL9snR2
gGA1/uaJV8bDoQyjyjP2PBx/odOwH945aoLhsxh0Ug/T679ExjcBEPps9wgi5VAL
fEIrm2Hsy1ok/Q/rKHcjRuYoQo6uy0ohh5vfd2BDMAHhmWzvU4uGZtbVZJcGAl99
MMCZa0HYG//tVFfpYfMAk7OxvoZAU8QQ1MYeg8qUIB28CeKE0Bn3YAgcsTdLbHOP
U4Imy15L9qX2QVaIoxI5h0TyCx4omEBQYDSZbXMcOhesh42srSWlL9Fjz6iykMvE
cX2fYaIjdaJoYeyZUo4k5nopF+Ex+6yKnbfj0eztBMgL2JQWaVWv0hc/CStVlvSW
wDCkbWa7BmDPvNjxIALRtNHM02amp3+lbKOMtPt1ARQZLEONaEzYw55y/WKlVKzh
mhc3dc0OJJbWbs24V5MnQIaQHU7qzXJHDquh58NGRjsvVlq0oczfq6SYhtI15ugD
E+NFOjgJcwAyXYtnwkrdPNKBzPKar1mqfgyZF2YxHSY4snBByWS+md4X8vlpSE7m
2MNqhiAnOvt/1jDe9vhcN94fjAhAn3vS0PGC3LVgOiS5r13m0EGGFqmH/HVsswE0
BNkOYbYWOv2JXdEE+wpdXD+AAGDk2zWPpsZ2AzJ9rkMafKGhaeAYIXlNdpZ7t3JG
mYpWITtNnrvt9YhHeMlZVWL2BgP9VmfOXSfgZFJa08MFBRDezRkLOsmqLg5xhvvQ
hJUGH9LdUdFcGgGVMgQpCcjNYxxT0MrXY92iJB3w0Ym/aQmALved/8x3AUmZqEVe
wx7/uhkpCb+27YlBPGYcGo8vzGCkyeUQvd4tY002vxFwvNnt+vwtcbvbnqHfABfd
8ybL4kxklcdO83CyEvgzbiFVEYBWMHlJFaxchejPs3teWHZJtNugHqA9oBzRjAfP
Os99U6uCylApevB7kJ3XZtcDTVJyN+YycAOJ1q4MVTHqtP4e3qa+cjta0XMSyfQQ
pbX78ympwfadm37Br6UkTz/k3BJ4/A4clNMYyqCHGCJnA9T7W1rHcVHQBfHBsyoW
No11MkUaeoJyIKiNHwFkt78Zrl3N3xuP/wTtWSJQp5AOL83QDDBnoKaQhBip3cYB
CxnQhPPyqenK8bkvUB3+Rs7H/5qjkrUWUU6F3aKSc6N0u0i4tWx2T156YpD+IYq8
GuV4ipS7LjU63nadseDIm9UN9s62yYV81SFemR2WiTaPNjosg8LOgNNmJR5tPqpm
rTvQInpzREjw+X07wqDOzHZ5dlM8a/TQi1zpx8ai1xLwbr/VtM8/5urLZxdQejAD
EQHoX15uqTT8xWd0vlCEZ5haN3Y7Y6E4TMuD7cZcVPN9K/3ZstRE+sp/CaXL3fEZ
B7h2JZuG6UOCMUS2aK8WkiUUJGZ1dC+gqmi5WhnvBGpp5fKbXzlmpZGtX2aMBHf0
vA0Qf8hWzLC8LcwXWPmOHJNLkI4cg2bkNghWI4u+bZqsSedPlKf7bBlvQhSdOI93
ADYMLlDeI/VX505HvgwW/Z97mc/F8/VSnXYIpIPB7rbgAMMgqOCB02hBR+g66PUZ
dht5egGO/lQ1Iumx3tXP5yY357SFxUErmbksASZnY0JlYk94bbkA6g3AX3DNe9nM
VvoUT4HAVwhZTCINZNJ9kxuW8IVa3kZJ7Yz9vl0lZbn5dbR/EBQzm2swXe0ADWOW
sDwdwMaK/e9lZPS9t6JQWG/g+6R5YzZqoXWmhzMEr+TYtWDJbHeQqKoZBmJfFhE1
N0Vbu37ZnzigPLdHdbPYHCGnD1bstKyd84IIYN7w61jmGAEITnnIP2ATM9xiJqRq
+6libcIzSgHUHfE8iWpUNJU8/+o++liKXwiPvI9ViwcLjicISgm8IeL4UeXrzFyV
/OQ8JoHOuZ16umbe9gd2Ux45b3CWXb7qaC4K1kwERRDQ0FS2sfGJrJ/DWhGxeC2h
sDukAEYvwbJ1xGzT6Tue2La5wxDdfOuf8x6BXtcqo4rbcne21S8tykyLPnz7lL9s
3xUA4Mm1he5XdUX+kw6Dyc00opRtUqCtBH1AtqOigqtSGEb5nItDOlqadclvv9Uc
OFZL4se/kqqin9c+4QnEXHUdZcggnkREWEnieU1V0o5DhsM4OW+jit478f5V7fqN
gC4yMINiCigfzPnLKSAZHbwRv6LHyWbB7GKO5XddeeGCWVlkF8TI/oiFFfuvXh8p
FusExur1kvU4+LUYb6XpomVTspd3gNYXS5ri9W9z6UjD+pmt2frrj0I4oQDd6X/I
NR7EcFCLLrISxwE0Un3c3mIcX+w0OWCWpOSN/5enjkkQofhnssRGcNxW2j6woRvv
Rl7cxxiAju7kPZ0G2FKSuvDJgZHAZO1EPGuD1G39DEH68GRNatiH/etmLYsGQDgW
6zh0S8E7uInZTI1ZxRJfPhQU5ZPw/TTTPxA3QzzHrtiysCWmLECN1BLn1nM6gx/+
UefGi2fjSNuRN1NRUOv+K9n9fkhWm6SMc8pUDN7iRIpe0UEusIq4MmjB0WIeeYbE
gGo+7nHyB5xpLf8kEDL+Lx8fxxCjeJRdCesGSGu1V8IklDe48OtV/+9VMVpjofT8
U6xNvI/B04gXnqdjmTsHkqazGbanDzX6TVKN//R19BOFtqs7XgnITzOuUwIsTidp
3Lc5BvbGoZYTmc1gCx97W+m1XtySz/OlqBzZwOgcVMKhc6emyBIbZB4dNkd87Qaf
stPJwYFtTwVH9abAT/cjx305JF5bIzXI/hanKUxSZ+5HrO/zBUrVymX33vOGXX5W
VQ7LRjptvOYeBAMDOvPDx6cVFt7k6mR5Bot1xSNo2v6EfrqxDvKVEoIDSgm7PA7M
aHqtcTtfO9QXZAskoDb7NHe8vzHpLLtnWVtZpf8JfdsIu2W7HxpfpgCgB80b14sU
R8Y8zEmxh0//llDCKco4LrwJLUYkwSxBlLWuI4OZnaO3356YJZAYn2yxbiXIRw+p
YNxxquM6Qd0E8eYhQZxJTYX3Y5rfS/xLYeqpyKvN2zyRcWRxSXcUTVLdiO5IOxup
FGTCujd9ModyAy2sKJWdmP8ITn4kKYX0/VVQOD8gQheoANg+BqYDD7yZPNWYOj6k
TOP25AlmYNGhX6XhmrEO1NBulymqZVQR9M7Dn8u84MtasX9w1hikxs0UY0JlYLOT
9bjf1NP3iq6vQ4o38VRp6GniWtiQbpU7vEozQa9Q7aY0Wpw02SjVAGFCnlp8zoL7
XU9YwyI1ANYXtxD+XhmaVlypMoSQU0peSJ67Omje1MLPHO13DCTQENB3bg/xFjAL
EFy8VB4jUHuOqfBP6EQCMZ0QrSSr656cGGITxUW36jirhxpVK0HsiOEZ7SRJc2q9
uAzmIuONbz2WEibWjkLbfzzYcWptH9xCNjK2hYiy9dYXVjGoGnWHvpYhahhzGmTG
qXtwixMU9cVBybJI2Is62caJ/iXnE8Ytge1HkAmJy2y0diPhJNgPGmWs9D6cC8lz
PQwW6IelXlBcb2CKfIUgWa00y+Au8Q/01bPFBNvJ9jPdQgdhDxvcLSJ5UWfg2bsd
NkPKHk4a51UbVNzFOtLtJX58q4vqglndALONJvX9wOlyKJpQVfYoKNrPAQpqzc23
vFEUl86aXU4bmBdoFXU+208Pp5Qz9Og8ko9SaEzOuzXuTSYSVAuwBlNYMdJtkQ6C
NL9rHBu359fdaElBImL4ClneyYCpWl8Hkg13c53nZPiYmREYAoPrfRL4HyQRoXwk
8A2XHrCZwLFXPauByyg+jVwtUeahDEfj8Tlz+bVgDz304zxuJpjYttjRysvRTmWL
7aZzlkxgf1VQm7VT7KDQ3TZYFKDHjPZ6JgM2FpSZbL1m9mNcjjS+I7hwLGpoqw06
FV7WFI0OKSFQg4bhvx/f70vTgiu1SnQlHylLA0lARNt68S87yL0WfT5Qei3FbEFh
BzjDouo+bEC1jMsQsB8ZZcGTLdDthHezqokuE/0U6FSPI4AYwaoR16wg3AzC0iUd
w/1i+VeNAy2Pl0cc13QNNlSI2cX4vnVMs+VgTQz+7kltfYLNUwPLH0GNPvNjD13Y
OgpoYk042Edv/vrLWOFl4CB0YvuiXR/V8Spn0r77DpH9lPB0CFrpjiL9eJff87Xt
E4eN8T4LAJw8Fq6YTAvwJQZpRvkg6CEdtkrRNLtQ/BgCr2KQHNTz528sFhYTLNEt
cBNsFzwGFpppF2i+tETJjctBd+wdWeZ8qlWYknJJjJHdnkDf3XwQJyjGPz05Qdmz
wWiYh8aZQaDvKbaHo3ch45cNqnU8DJhJJhautBdAsxr2g6ulsmnhbR7Dlg0NhKDp
CSAMsVzXne+dIaJz+Gawz8xn95twmwINzgw4dUChkH/Z/EmGrttLEeNerMifDVcy
H5ZgMM14WBWjfmsVuRB7WVDTstN4yqv7QjnG7QSPVRgPEXECPPog5A3/xn+JnisO
0xP2jjOLLArwhnnfR3bAIMWvKRotD6NadXWHP6NFzv50xtGufghig4RQyKhntjVc
MaIvY5Yw0BfE/vHsLV3zTkV3BAYW2EgwQthrzbYlBZkdHQOVpNwsHnqBcQ08AUL9
6/rOb+SWgdHF6Ri2vpCv02bHHf6pbQ7gG5yBZFq895CTBhnpJY3SMveGr+DLvCWM
/Enm4aSOtp90knMVMqQwla8e/SqBO7mZNsWsPU7hYc6k8/arwhMSYSBlRZtig7SB
tBzeRipH/iaIQTHf4wyBvWwJTg3/c3taCmAc6CdioYDAUBoluASYsL/doib4K9Gw
pybHAZjLoIIEHCtr7gn1Gund5aBA4qch+8J2gewQWyzSdBWczfEjZ7IEaDCGQoNj
PDbjU/pLFbl9C/iTyRlFOVUXV4iNp4hBuoCUuW9I4ZpIV60niovtM5P8E8k9XnZ1
5OfwmqxJzCpCTfJf7bNSV+GmYK2BRZ02+9/9K8U1QEdnnODDCkWV6guWPMYQxn9y
KZ2pNl8P3s5ldFtlaNBF4844aoapchaI7X1QLNCmEd8IW8AG9K5hqjFGpvF5U+A0
EnsKkLLlwL7I4tQ2DPGlfzjDQgfuYWeBLkDs0NUS9G7hkoELCPFViFjSOeGzXqC6
+tPgKwEFbWVT+IWOagRnG6r0BvZX0IGMQhROBgocKutmUXXU3JSyoRdGk/XokdqJ
+uTnDSVT4bUH4pkmJwBY7Apj7heLfpSUftlTez+gNceh72q/LC8NvsceAO/ACBsa
IWHD6u6lHyChSpI33+QDXC5EhARVL0G3WQ4vwvzjGY4wSrU9nJGta00nZI5EE9xf
RDNrMTZmU6Gx6aEhkdzsZ6/K1zVDfyWTKMIJq2Xmf2dSHcXnhHv/YE7vGPayNQVd
viBqyLeXVxw3OxxZV0njhYvqIGgmfWGapi1YMzuttXv3HDY+vtsgMRZRjwTQLv/Y
63cRh9IjwoRlOX6o0dd1p12PbVj85R1fSTck+gCV2nNk1JO6NMAut9j6N78fMxvD
yOaLj4/HkTElpu79zIcv0CqOpYHlMR6GhBEU9zSB16eUABufUKBtdoqGiGe0aXVs
UrbgXRefcjLMkzSecFvi3ATPzro70Xga/dHYlyJFP6d9NPo53oC3TU+m2yV5OU5z
79lWi3qF+N19Yq0Qc88tas9mOALeOqZdY7F0zUHzI1SIwIqpQnEG1bY38CKuG8oY
4KgAtzkX7i7nSfaAhLKI6xZDvF3f3D1B3iTYwGc4Q8hTTqGSs160wUfWj2SHQeWJ
ylYc93j/TuzynOfFtfdnz/eaTZm0eR7Edrxc+N8/wpAzKvjjtzl4Hy3zE+X9x7bj
b+RZgDZmmCK6rgI9Ns3A8wBl/jNwS4WBFPoM2eoR7vhPG6dWS7IbqmPbFIFalASK
V0OfdL4JEnemZLi86tzhdWaeg6XJv4fBj+61PZxFSRiNIluXXUCMT+gV2lsfnWbl
yN2NASvAp2K97FXg5/prSpiYcZrnPgqUn5XUytQxjWtspIGPPiB/yma+JiXvkl+N
azivw2sDzB35agpP9/0xrEl0aPBMfRYV0z95kaaC3JXrbXrUXGPNCfgMZKGt1Lo6
iL40tbg8v6VS8DOwZvvaGxZWG6K2uKir+EmMJjO58L/WL2o2iNRoWB8BGKVapKXF
pQNtBuUJ2Z6DrTBK/vdk9Ia2WcG/6iVa6LTQxOM99gRKQaXb+CbTZw8aKb3Dhvv2
KWJaURfUfTpvXI7wyHjoTG8QaELNf66Qr+XYQy3x7OT0QpbEOI3TUB4GIX5qY+a9
xDpG/ZCinm6NEydar7W1lZM8jUCPXDbKZ0DQ8j4vGPsi3yxDQSi+WUp1O4J1tZDZ
kTml2lm08MvMOEp0scha4BYVdhve6W7ppeeawU7+fK2cxl21lFw7+XGmUhxFv81l
Rib1Wg54fiNchaCEG5/onDhMwHxNy4xWeg7C480Rr9poKNhxxOliwd7ZetkQkTpT
u2XOImZu/FGSrViI84/iOx7F9WWybTBiMtdHVucHTQwdaYbEOsn62nyYLB2SzHGz
hioDLVXQRWo2Zm6WtGstJwco9AOs8vpi1cErIS85sqfSQMbhIUdCaIc5aLytF7hA
jupLAfTdYvZbC7j/4CgYdDyoQ/ufIZLFQP3wsdyBRTBFK9WMC8I4ro+1Lm2856Pn
S/Z6zsnwizMWWQMO52anCXccev6re05ZjF++kN6P8X/3gIsJEd5pIkLUXfccfY+s
Znuq+enKLP6OJDhrE4OHOA41S0Lw14FrII2xt0GPV8MhoSduILZQxt/iQ7asT2xe
DQqD4z0EWCMbyhDah+ZubMwDT/aFbSx10dEfMFzbgjABAU/Lx1P7oCx9qYGi8VQ6
RZE2lEuug4YeNwXOhTojuCXdERmxA2QWW54uEvUZ5cWwTuaXKplhgeiLiwD+CNeu
lb4EgyGwpIsmbwqS7nFx7Vo4RNozdYLaODp9gADhjHUH5CWoqDkcpHl++cmk5dmF
AU37EIuWA2iZm6DUFHNqeO+tCzWClJKh8itaO7bTAtHe4Gw50x1wFF2zludD9PvD
fIWXmvFa2pHNX+VD80KDzHSxj+Nujkh9hL/KLP3kcr/IHr4cwuBT1dnw3x6bKuaY
FI72Ko6RU31G9P+K+AiT+UNbS3agE4h2cXWKtwTevr9R7TFSXuZgiUeitO2kBpyO
UNKBhJaWm6foZqrbN/P+mzxLol1HBt4CH4DIRxB1t4/U7Fav76OxgUszgISTGAB0
Z+Jed8tcdpXH+2s18RaR1gFlastoHUx0dRMFgh6jQCGGAjNEOofA4wILT284CEoW
pUnLgJ+9/urIw0uMioPFtSuFyxtyt02F0Yw4pstdHbplln1o+a1Prtx3ZSO6xczV
tIUuDPdlT878vKeAhqIKWUu7p6GHMYxb4CTEubdLY9YrrTaePdscrV+uJYtxCK0G
f9z3Ln8ZeyWanzDvjKiBe30KUJPvD6Lpuja+YZ5/+/25LRXXAeR7KjFVWGf8EJc0
4+SpZXWraCKAwL/LZhR0bxY8/5f3z5h6qcotBqpaeEkzXZ86fI3mEiXq3yryrZw4
UDTYNYDE30IehTxisnfBkKhSdrCjMPErA81R5XClTgB3TuZDJTzfhcf51x4xEhQB
lhE6Tqz9z/GMEn6HeQd87dwfMniI0NnnRuVUnj3OMhwdbogFxT6B7ntt/C/r1Sdb
aDybvDEjPcE5LqfFNZcLTxrDvyz+z0OCsIr9bb4FvqRMJERM3E7zpS88lZcMY/SI
xqshW8nMtTq6pumKbcPNqQCvXWpkIWRiBBUjT5I6WOvHHwGmNxTwSdvU7leIDUBA
tVsIr2cpQkCIoLTxbKRgsLHQeUH9LhaOg27XFw806oHanWU8QSoS3rbzzvnKhDBE
SSgtDUKMLuWZCiy33YxYNXhL3sPQf20mcHXm01kuQwj1+TsCqx6GQGwdnOg+6YRC
ybth1Z3SmMze7sQ/eCQWsb7bnpwDkCNf6lYFw8VCm2ud/7PbyR4mzkz+GEhj+30O
39JExQ9tNjCIhTT6seo7lfx7t5LBW5VPH82ErCjuArJSMUEcGc4NrZ1gvex5UKIL
r33VtUVJJ9YK8UY9y8LoJX4Xln/t2S7XeolRi/dTHt96kNWebJfAB7dYGyujhSEQ
re+nqeRzVJhguD7xvdha6b6VcaIicjXmH+Iyh9p7dRStKo9dxv3QMKXwi1x0653g
SkBtUDAyis/qcWdApI1Hfgcq6f6gmRLPG/dlciEMXGIpu6lgW8pD75J/uz+lh456
S6o3yZpr2Ew/cDDXp8xpfiuOsnHpDfGDOAwRzNIjH2kzj3G49CFxUyVlMYmoSXFJ
GytpVdpQ6dh3Udna9zAqt3L+qppJO5yuh+06WHsvgGnQVNmLABSzfRG3UuriNEN8
kbBWDhIYHcOEDjieg9XUgW2cXb0rK19OqsPNrkiN4Fe4+WsDbMo0He1wsEmoULyw
jFDJSLHJce1YTSBcs6Y3AfCi6UE5pVAHlJrkYqnsUeNk2DJ4/UyrmvBPwDktck3q
tiL39X+hJDcMwUMM+RcV7/qZUwO9DaIQ6cDkm8MmIBZzaohCqmloeliUJG+1rJTf
w1Zlgxu96XZzpbh/VzymhmSBAuwyctm1v89rBigu1i/JcL1I5GX7W7sRlnbQw4Qo
75/j7CU+iZaPE3rEC8Qw78UiuYQui+BC/g9qOoA2jcUZ4RS6LJfcLvg7ZcZwTAPF
9UmncMprR4puiZgHGVIjW6gTZtnpUjhUZYpg7aHcttWx0Dp7714OcbgqO7c8V1q6
t+O8Be8qirYvFw9/kPAXmhCm1FtPceb0J3Asq6Zt9+aCatFYYkm6ZXqR+xkukHdI
4VZ9IVZ12xSXIyt+X2nMmMoWUF8XVXi3GcJCzvsPF+aqG9XHwJLj83dnjU6sT1RF
frm9dDxjcU3dAEt4Nb61kcbq1WjxDOK37TRdlEkt5pnvnh/Fn675o2gtTPrpLjng
9SpSoXCKNlhureCdggK5Xhf4l8LlpZ/SUEBobS7Pq7VAliwGER0uVM1RS5fR2WNa
giktysqsSq7TvZk6PT/EKIoriPvuyZ/yaKOOXLSy9fn8xRYCZDphzDgjPrHqot35
BTqrgbFvxkDShRnsLtt98X+kLiZlE1FFjcGtMIXAR2CJAjz4/aMp2LW9kfJMI29g
mezJGQmKti3EATcRSMHtDladMqTSO27sG3s1ZhlBbdlHFkqLBSA2lJ65hmb+kjQ3
f1itdwrt+gTPPTH+VrfnrNpI/OxnFVr+Ao/6ChMzw81NBa8f2eXfPAHzWtkydxHF
Ao8B0M5i9SdNi0FJpJJVRUPSEt5DTDwAGQ0yEJmjjHmEh7rYmDmKUAr6IKLpLtSZ
34TH2ycFAl4fczy1Zlru+o2KsQVqtsTbIcOncGBSQaQfZgT/6S5KdLwnKtTCnoHs
f13Y+P40HDaGjryTWbkZcnJ34SeGYWzZp026qCP2pwALkfUHdYkyA/iYRSiZ987r
KrkUwzPrHXWm4Phn0W+/tA+vwekh3NreUxbSAq54KZQMTQj/gmhBANufT6yZ5Ljx
MHtKPeNOj58CjIc0efDdEPPkCFROU0LvHkspRQm+kxomPhr0lMq+bJLqweSfJ9vF
N1toTDfxnNZWNAKHek8XmK/kjHDUh/HwVIYbuD6LwdqkKLA1SfT6s98dfHUc3glG
NGvsWgVXkZgyByAL/cwqhOZUIFL7nazpWBufr4VMGwO1uJ4FpwVZ3I3cx2fQt4qT
f7dHlbXCSB/QAJLwz6tdgrpxW+jpWeQJuuUNJwds8bWQozsJuY3qQ1zOuFCMiGXk
Ns9HzKu3y3SiAcMGv6t1ujZXQmlRNv/YijjV+cu2Y2silvcQQkQcf7VJbLs9iNht
q0hwMX/7+e6TGUDWjgC5cZ3Qe4GyrbKdfBPStUlbP/XErUK+GV8GQRTKJlM9AYZh
KJ3dOvS70sXxp0S5Cmb1kN462MZ2kRosAOSZ8m+eBMiYMu4TQP94KZHUSjEp01An
6vEnUMtcrmf085SkceYxuSWUHymjlUVXBWgO5S3pFsOtBcTSZvI4616meonbMvXl
IXen/RxIrH8wANq+aDmXncCMpCv0c18lJ+d8g3Z9JX0hzgCe7gt0Oh925m4b9CyL
1/+wUA8cRhdbecu3zX0eAD6pLc4tDx7lwNO47JHl3dMUSB1BFmac1PcxLqvBhhf7
2Thle4V0ZYzAlwKMtCXRrv0pGMSzs3okmDO8WmnvX5rnrn3mCHefC4OWZFXYO/2n
+xDHktNKbS5d2D4soiqJShQX5SyTum/w/ztwB7UyBh2XceAhKTuHNWazwjyNY7nr
LMayltyvHyN9Tmvp7mVoIOApvERQgNg+kDAdJfbVJId8ldDQPrh6GlCNxcgQAuMR
GqFk6yfL3scxrTvOSPXdisbdTfpJWHJuEZuhDdRhsubmo9aJjkV5WUNC0SN8SU55
6eiR+Qi1nJfZT7rwC79dRWB1kpDVAQ0VSLZbvgunPcgg02pZOafyzUMhy3VdQMWo
e0nI9n3nchyRsmjobEjDTyVkpfouEcHTvuzBW4akA4y7MCztjxQeDUIKTFuLIuJ2
85dnpRz1s0oJiNZPPo82Xi5/t4kybu6ME/F7U7aueo5slpzZpJaxislTwTqSZkEm
MbxHz5bB+9czA836vTNXsk+06nRQydxqSXu4Sd5ZDkH176vK1FuD1a755URmOeFh
Lk5d4zR2j0ez6sNhpViFgNo5AqohnMD0ss/tMIWPr8Q6KZVFjVH3n8bYbNta0xs1
iA0q3xALv0P76CPkV4Nr5pOHxqw5ql5/9y8tD0x6K1nVBuQd3LPVckt1io//ugnL
OWZ1sblVUFFjvAYDGeH0fiUAlvxW7qksnp7B6s1HBmjwh117Psl2124Q76WTCmea
W8PKPvpTmv+D7AysvvIjxOy3areViMM3g2/weK96yILYAO07jO08pw1fdI1yEsKS
tBIFSndQUX45Q93mq6GJ6u72ddYkJqJws/O8NickfEVZAYDbBu4hHavf44HWx5RG
/TOMXqCpH2fbuCRGg0dKwdYXvQ3lsaOsGoQrBJWBQtvhKQKJzD14XVAtU46nnNf5
4PaeUSxJT6ZmUwSHJw5a83NkuTiLMorhNgzYcgomH7TqMwKQfocSyGl+Umfp77su
BOk5cHOUSvzFWtBRorZS8ZtgGvw2pZZobbK/mjhJjX4z9CJkLtYdL5TzJM+7IoQH
GSWgwz6c7blOnbG3Oe6Wa5ZsGEFo0YkLuk+Xf/x4i/B8FdZcd7Tr2zf0n76uL0BH
TBCDRfXKunpNNII7nwpSsjCjbK+FD6lquEx7nDgIJPgWvB44NBA9GECCj13F2eFP
bKwnwulez1bBwnyzAXLLLL9iluuhyLHHVJHHlLJBKtQoenxPlILC23+7Vhv0U+FA
Vk1NS7QThHx47kugjfdImz5dfBpXnd2v3Ziu/qvfrMF/GjJieQMDLC6lQM6HpmQF
xjEE/pPNyp5nq6W4OHhQ6txCtP4GAc3yH7gi16NNSlHSY0seKIF/heW7Uev2cly8
2CvAeWPDGrrkmBHZ6U6nR44rdylbsQce60vNfyNFINyuuNhxfyWsxsondupiVqDJ
gfXrtVb9Ezf8HyZ/69l4xhlQU6CnwOdQigNykqwqBJvq4H9aUjAro72+f6RZbaBh
KrV0MhS54puGgW0yp9i6FNv57VlznyIeQXIXREC3DgcC3AQysvTaljGW5b+jOQyC
b6kkAxvSxFtFwsTlzskkJ4+sfs9gtr+ewM0NI6f4Jm9Cm1F8ZJ1ltATCtmi9Azo/
yedd8cjVBr4c+dkMvoalC8XldDvvgWOYHTaT7i8xL1PoIHi4qBC5mEydAobBI/zo
H8pKISXBzgkUxv9ct4uR/rvasvhw/8BHy6qoRB0heK1K864kCrhb/4ob9yZSFsgT
0arCqPQqBPPG7KaW+Q9AI64u6j0V9wnFX8HwFkYNlJc1Y4s96d974b2em4DoPq4B
DIDhLzTnRy/RPNENdnMYWI7gK+pxELD6a1B8XwhS7YIZh4ddCn10mG4/LrKqu1mF
1hLDf5aoSj8kam4lpkwNt8TJYv1W6fUDBfNWRXFXV+pGrIQUalwIrQ8Vda/eAssf
qyMlKKCpG/Ws+OYNuN19JgQxvTiFI9bTcjZ/9aJDaxnUJCcE7xONvEriALen9Vlv
DNKCN36FVAqZFHtHLQsXSDxd5BN4A3Ug1bbixIZsJaput84wlqMi4P7vinH7Wjop
Enh3VzWfPztmMSmvIlAqTK/6yodajRxbZhxJqWIAhuzZKI9bIk1l+lw4/O1Dl503
wK23/zdwF+3dxe8WVzxPdKULTJbvLRKH32qXCnrTbmaJvd3lrChpCMx3Nxs2qgOA
8C4DIYlk4r21JiKJ2RAtsrIIGNEzqTrGhnIqc3KdT7/5tf6OBUBMVj7qRR4OUPlh
msLLFwE2DYPM9YL4M8V5BTwM3OMqGj7nvCJAZaYrG4ycyhjNVNTQhcEUBHevMWrC
BOVW4W/tP1x3jouCh8EV39PKAJ3MBOmbHl+X/DRL/PL9cBNVGo+FehJhGCt5Oyrq
W/IYD/TEVQw9MPyv41tlDuHOIAY09vkQ6fiBinRNvvH8q2tiAcI01OVvmzwhzScg
fDbjxj1cN6aP6Aj6sAabFHeLZeJEKCABfjYWjbp1OaJjCVEBnamW2OMuDX5DUYkH
T7pdD4hHVZ5Y5Y8rTqO+2kOVE/ExOXjvRATD5e55i28AMb9P/4ALNu9T+6YTH0zq
0Ixff56SB1NxQJlbAi21AZSMg/W/pR+vZ/F/+lQB8B1MBhagZwML+/rQOdQmh5hV
UrIuDz++HF5rblqNNj6IZwI8X9HpdpNZjW9Z3reqVmSXGL4+bDLiQi10AqVHm7W6
CtcGD/YY0Yfk38KtD3GOddRJ98ynNoxMtBhfNVNPHlHN8QGfpR1xoZi36veVwxKw
sRz8zI+YZvgOY4ZjqujYNKcs9+0DwpkAiKhrgbCvaSjD9m3GWM0EvoTY8rrtq1ch
ZaVtCvfHmJtw/EiDFoTxyx86yXjAUdkAaqIUHFaQCP0zDim8icAFOqau1tBybUvC
UUb7DFYQDUl0asORsl+c/5vEBOEJvqbsloO3bn7YxZGOnuOv/HkwOmvY9qFZ0D05
G7YMug078A9c11M3SvtsXMPD5FL9aFhuofXzn/77P24eL9FyXq/BSAvELYtz6tCT
3Ll5nnx7XsM7etVDJg8Yg1N88My2TR9hDu3vSxNM7hrlBSG40zFltxgiVPglJ0N7
L9YOmnUvK1zZrZMjG4Eh2sO1/c/eNcvhsdBkJQF2enkYhePc0swMhrSYqZnihY5g
H+35oL+/GDgDgPtrRexIhrehHKbFG/ocajoiBSsEoKKOn+whoUe58SEcmj0bs38U
tIYgHRyJ3px02Px0L4jiMJgvE4n9rD8ycAeCdM3daIsdqkLB6ZiBkF0Yu/H/5Zs9
NI3Zscy3sw9ccaLpwqtDNEdU7FMs2oy5VHAVThV2/+ZVSfwOIAgzGl60ISalyBXt
toB5CYNAcXL5HaRscc37s6a1A6LmZYGBS4Dqgyb6Nosd4mq7/UdhXkNtQK5iJQqs
QW1ScKhG0OAmIqRIumWSCNB/SaIyR9xV6miHJFAa+vcmyFDlAqmwZbjiTWNL6vZ0
u56fEiFP040xIWKwKZtSLtmjM7CCNdP2XFvME00g5OXoFWVyyMFLVHjXJKY3xzQ6
EQLl1QWur45VvTLkGJyjRlTWuDjRJmiKFZkq0XFHfC5zVXKwS/nMucunkTOhhPqI
1qHdSUKtVmOzriIsCdfjLwc3rNoYQATpWcxpHSugHT7MzTmh1c5hRRD5PhebFgZV
a30+qoU/we1re13x3IDi4VJxuNfzlPT7SpZVi8QqxMmUOW1tnvVW16atSsBtAkLY
qoAoGkkK/i+wv4r2KUzm3GD5Nhu6CdaDvZqOMTLR7HeGOx7tPNdeL8wGecrENJGw
3Hqein4ALxqWYa0t1ILRECsGY317Odsv0oD1dxiGmeHrCIpvsXsItJxWEUxDVrHg
1rbm289bErvZSEqWwXnwEawbxIDqOBoPeS05K4ROBaOuDg7ziAfvCYVseJcGgv4I
VdmHvPHrPlMxTWmUNYwGU4de4Ljkc6fpZslE01tH8fNFMOWLWgqusSgKeuNXBi3G
4cQl6e2Dl88mFzh8clZOLW/8RT1CeThyE9RAzEkrSjMO3g8ZlvddbunVHzs/WfO+
hw8rwYWLDqTF2d2clU0uAN1N33s0+/sK6pPfQNhCyrNiYcWG5MDIgmwr+0goG1CQ
AyTkPcnaJd6L8NSNyH4A/8CBUqgpGDEZN0fU13Q15eXq7M5sjjrZOBEIt0fMmEan
dKzpmNtm3wKg3qimsnIxCf+3kwL9Za4Dm+D7Q4ThBDqsvVa1GihH3KilZ4kpY7GQ
ZwNZTCRgRNeWQdkI7KuObNTRh3DN/2C2gtQ1VfuTwsnv4Cx8u/FPfAS1mQkl0rwn
GcVuC2+4tLOHR6LDjAeMGvRWPVRXD1VhcTqjs5JTMVmnjmr2CICAIGTzpecbFPrN
aXBpHfgWft0NasFXt1Hf7Wd6B+boDOYvBwsr09xztJUWUdrIh/iueAyfDpWv/zPj
gLRICKuG+Ds86Kd8MPmqu+KQj7BAzF5Qm1ySKpcsViumlqnQQYN1qd58k/dPjHkt
y6/Il3oME9bjoHJwbxWgW3q5AWyraAXWyVT/vzCw0L6Yy8LSH7/upRKP5VCqSOlZ
q6SymUJb9dCNT5FkYOKfukmWEfgbqe13n7vp+wnZdrqbJrzcUp/A3g/liJFKjkVW
6ccmjKrFoL493FGpAV19v92DRS4wIZYq3qIVvH2Fn4GrlYhIx0WDp6c5xxYJqEXi
WkwxK8q2db24Ig1dE+nOeiWmwZ3PEWJpowJuL+JH8T43BXhnHAAmvu0qeJI4Pwcr
YEZ1beANkl3y8VUtWS6RyIq9myNH/P/XW31IWpweBqiHJ4+osL35m/wH897HElN2
Y1Qd9IuF/i0H88Jv7D1NueHPRRlf/+uRoy7EjZnDFsMJERjf2HRfzQyJCJOzXoLA
uNuQySkMYR5Owr3cPZ66tqeCMwpSSvSsKGsJDXSq6PqN2nioDS6ezscSB3UbsyG8
Y6wfKxQZIuInX6n5tSZTvE9Fwtt4B9adMkD9SO3FSqqC6oVyIs0yhjRlvrmksRwu
wZo8jK+G33/O83pnqLvqTH3tuefpF9qey/s75pUKOu5EEGzBNLTYrGhg0gG9j3UB
sBs6bPSdsH7JXtUCdzeePcI+TMpwQuLmGHkUk0oyuuXyZZMelhGADqNe5mZzesnR
QUUA897G3sBXlat/t8P+JWXFH+Vb/nV0BAA0Y4n9LASmbTXlpICftHlt30DAgsB4
PFKbXAGW5aK3MppqfgjdyYApcK1P4Fh2kPCEKsoD7wkpwoAv7BVkCKs245Af6UN3
zPcTeNUQqnbl6ZrMlUU6BYMUf3WGevEYWA7rmKgTgc4zcpSRbsWqj516tmsTS+ZP
K4PQ5PFDDtLouXPt1m61gCb5W2hFxZOrhPc64NNF/aIwex0hWvmWtL3/149QR/CW
qO6KXoFH1PS+zpbshc+Q2if0khVFYr/XyCck5LMB96H+dGXtOqVNG/P8WonTYNqs
jkUAuwUBxGY8fFFGyAsHLbBRLd4KZi2O5eFd2qRhwy/saboaJmor2FFcSqVR/mXJ
Vbo+Kgk6Xa7F1eX51EdU6yf7lCLnxtsGmpAC0dBXGjzxjGAQZAz6zJxJYELsTON7
XXnnnL0DSu/o9vqf75OOj6fjQVKA1OSyh0/Cvr2mcBwhZ10jvzyKxy7BZdTgscK6
6O7e9ZQvZrD19Pv2YaObLwz438f9roSs71mYs186H/XVvX4LAEqxQFIq06xtqdXT
EhUM+g3VklRqK7H6lXXGgjozGaVaE/I5iLGm38O6qqdxKqQVWsR5OIWC/P7jlSUS
NknoMdAtkANZjLCnZAD7joGTnEJzdwvEHn9tWSeLj8GrIZhaqDhahr68KmSwryPZ
XSjWuAfpGetwD3Ppb9vHDP19oNXP6OiU3JxeFMrScm2LCAVMZb06Bxbas8NdFkdz
ZibNoSuwOsWqgW6RYMnc5E9zQNYq03NL5nXlrlQxM0sAGu4JzXqLC7NS+eOTdW2d
6zKUdhftL88A6mdtLHwDAg5FNIL1xEqOiJgb6Xr9Omd2M3hQDBvNjkqIO8c2QI+S
K9+Yn/h9DZNTFbxdRdWD5LfUlOgBN2oS3YZl98U/ZH9z2xKmjQ3JhTgVWqkvV7ha
z60vlKIDtSpLjPWew78oady9Ks4EiTxYZpmzCojWFKYjPAw3UOC2EXrkTxIDDiFx
ZWj/8nFZdMoXl04y7tA8Mde8pTxOOVnvkycp0ghckhducxxz/gojnp/XFY2+yUgL
9ktKlTM4FVVepbWX4CNzK1WVJA2cNfbSO/p9KKjOOK2khgH6OeTvYmfIrJF8gkuB
OSB+yrPfRNCQP/VdQAoP+RuLMUl3ZfbZr0he3EqQWjR89hbo1i+JLf+HmHWlGJGZ
H9GJb5JlpseWeUPe2FgaVLEsO1q2139o8cnnrWLhWuE5gNNm2MrKuBOxTPq6FBzp
o4adc2pzs7D1bu1uAccNFpaEcGk5Zc0HDV+AakXAfQ1lDLESX4+ziH8BD5/TBz58
rofbf3RGZXk9gnPeLjMWUg7xruRzeY1sFAEZ6kvQFtRolw9fzssLymDlt0O/ezFx
6cSsegwefisKgZt5LBne5hnJJCqd/QfIpPEO4hFo6L1DOSe1P2I7OCVO4Vqm0Xz+
sD/5OZsmZG87L/W4AadTuZdL1L0U4RiEzOg/smVjfvo4mnXnr2saWgzLmVd6Gx96
KgZlKfnE0rKlVQSM6JYTxp9RxMrQ8X9uwrV8SpXI67BuCva1Awde3/HTLyrM9U+N
SFZrOTPRFwlHDwZLaeipDMi1xR2c+Iac1Vq/PZWGxtswmd3eY/42LuksruN2e8HR
ZCi85X8+djp3TO8PVFjv+ccUdU50RNe/xPaNo925Ywh9ac/6Q1KKNO7aHD4eEOtd
cRkzus/I1gA+bVBngayFdrNXExzJKSQMkZH6CtMmk4RkL7qeEiSQiUdUn1X3jgD8
3RvK5bj7nI0/dkXRZK/j79tVaqoHa+2efamaYkOj8nkZtYCdIXI/nq2BT/Xlj8f8
4+XVUAWogOSPKHYeaNg7El8GW3axvObTUqmhxbGzsvEWg6JtbkCuaa+AVr8GAUFc
6DS11WZsuDJBZVp07mDsIHfm7T3efHdvlRoYZPXLNQoz3eaAxg0Jc7ozPD/uRrxx
hDmueQ1qwnTCjov/5LONI+JR0O1XjwH11/q/aZVLFTV2ZbWflezCZ2sBgjaH0m5s
ceT9hTCxW0VaFlkADNCVvFD65jVpH0vZL2RQcepHf0oIbz/WMnMO/NsSi3svvhFl
fLkIDfqcSUu67xvGJdFMV2DqThkbuRkbrJBt+hIW81hNSWXtxc+Kmqdm8aPDuWZy
gr24JbY/9/3uHxFkCiyTrd3xBfN7Uio9X9FSNK6qYKqQCggCRA6+2emEfkQsVF9H
yokUa0JXRx82RfzdVMqEjC2lQTcqBBQqyTIp24hcVPSxtjmmgK2D3Yo50FkKdK7K
MINMiPhoaHGgqvDIqjIFRREVJFk4yBqmXn/s9dyK5CWhce4bnujU5fcQ5Ly4lEor
34yKtHS+kXZazBLPkwKZ7/XYOyt6QfXJHhesKoIR1UcTbexaSrKfDX+Csh4X1yzJ
fS3uQv+CJLVEY9MhLrTq6vaES8AQkxyS0WPM00rDyitG97WAtwNycTuQfeVFs+R4
zRd8Q3h3iGGnY0P2wZS8bd18WMbzotymAd3kLk44Ddtsuex1GrSdDC7/y6eKFIey
7Ddw0MnwwISKW7kmHIZgLepunEzPKOSvaUdZhFVSGF+pamGjdkRNdQW9PjomDPEt
j9I5xPbbQOrKpuAdzm1FK3qX71MuzQLOfrRd12IQv7tq1Ck5m+rQVbElQnoa+84F
WHY1lBYB9krv/oIY5fangiYh8peoOXEnh1LyqdyPDw8lUt9UagO2K1teOlEi5NS+
eIqoCQFSX8tWIewbfbVOrnqOCyMtspu/hB2jxhaxx5CPky5tjeV2B1qg9i3hnIMy
e4usyHrM/kUkjGHAgsOnBBulYhSHaIbeqIdVojxCmBi5IRUB57ssEOyoNXuvVz0S
uOGif5LGN+MKHOXZXqiYdykoC7y8asTCdFpefPoBS/Xv5jgH5n8U7YqqTUQ7wM2L
UaQbz6+QKm0qWI2EEUIL+qMg3owz5otINDqtPLTXavNcKi9SX+/K6fT01ioH3CzE
/duRgt4X4HXDOkyU+Hz53dxGICxT8fWrAIFTUt0vVJSmaoseQugDZsdcJoDU8Qx6
4crXjlcDhHiABWMbIfKlUBiXohgc6mEzbVcpqidTWzXZF5Z+pK9XE0LI2LDxxx4H
PDy8nbFAZeOxswbENLqA03ORKYZdHXhgxvrailFeItM3BrNOK8a3/aWD6oNdNz4W
yxJaTHVRNCIKTrlZ9JLFez7SqcKv7MuK96dCrugHtWIYgMk+uTtHXjV/k1uivP+T
ZONy2AxZMhYO77sUJNhFylizwVnrtWC8B7oX1S9BW2BCttCc5ZwPt/zRfRrplX62
gCqrWT+GR2mWvY+mRdB7z4L3ZyJGFl0U64Ob/lolJ1BEbZjRmOUiNqCvoiRFKS9/
zDDZJYEV74lYIAP5JSKfXvLWI2XLkSMkNZC8+LOCWF2xf65J2coqMBMBN7JIX0oy
tgw5OCG1yuCrQgDF10ClgqWVcTKsLiIGofdoVziOi6h87T2E4buls0j2Lc57gglW
4raEVhe+CPBbazNVIWXWbBiN+A2rWtDJmws9+Uh668uMSQK3SUIhZ/3vyxhn+W3c
VDeds9a0+dko1/FneZZmObg0P+acJvF7hX08764xPrKbqycxU6ZizSv6Nt1GK3vF
Sk5XZXUmLGsFMSQyIiMxK13/c+1XajVaRZwC+3f/tTaMFVMWb5jPpE8IUdAWu0ur
qGALad9Qr9NydgXCgjXW+XucGRroEQGQc4r/xmUWEeGeXfJaOljOngNRMzTEZhcI
brGsnM9QPQueaEot6fgNvjKrJZ5qAWlYIOPtHZKPZlV4NjWPRozq6YOBwKXfeRXS
g8rFcEuiYsflfcTTL2Rh/yI37yAo5pTTZkIUb8I4OCV/b8LHsiQy6M3zl26N9VOt
0cfbfG0Augk2FcqYAGKg9TVa4CYb+wd8L1Llhkx8zJo3GiOV78eecDzdYjuPp5C4
14t/B7lhw6h/fKOCw1RoXLLD51tMYCQHnQoUK4aBwRzPBEYbY1NZlOtAr6zExca6
eNtclG8j76VUS1ZWN+nRsFPDy6UhA4KOkG3toviHeXbwdIKopcEm/n5MjKYoJEqp
ohKO/4tRl3hCU3My1+hTSSfiJebgOO6cMARE7BIhGJTPs36+kLoUC/NWfUQcl6p6
okKWuNisw97uZzJbkbY9bmbbYLBmscv22/l90MlpGQH8/x08l2WhuwMPXOaDsFUJ
fTiWil4PbQ9gkvSTMbLFxLaqas9FRBrAd1RDMvQpkobW/qGfOwBpx2/gqsoQo2oK
jM6OA2mchHwvwXmKgMWcXwwCxc9P//TitwqaavNq5DRZfED0/P2BWR7QnJMgJkMh
zMD7J1+/jFoAjt09AtcWqUORKA3GAEnymSeNCLy0wkmLwhFitht6abSZcbTuoygZ
o3t0Mba4xbTRVP7+kH0xGnX0vSZzQCkJPP+AEK6LPbmDyvxRSdi3+0hHpwSWqvbI
Q0987mZCTiH559Poxvnl1926CSq+SmEmVPu9uFEwPo+w7J7basV+fpJsngX25oQM
DJQmOFoRLe17k2TOwGlOmvcjyA7GRAPTKiJW+ugmXtfytAKIii7KX/KZljG/O+jF
AJ3RsWfVNMSwP9uIta7sZOhWYywK3FfgpbVO2h8UtzrZRmmBbgbBVySgwaW8062V
1l8mYj0cLSfGO21s2tCPvca3S5iCqytA42DqkPlT9++zP2rzSy3ODPiTM8KyiEWD
Vkr4ubv9lD4axDFDYRBE6lezfAiwe+RJbMNv3NL86Q7vLOOKcXcM4OA2EB5jZMNW
ZiAj6K40tGYMKWjQsUkLxPv5PmrHziPiwhllfxG+rDw/CeM30XJWv/P4zVKdnAce
xWC0Im0CmDWnX7f/a3oZ/V+dqzFsLrlgkYDj3+iZ6iVGsbbsjs+sDaTvUHRTsruT
oe0UQG3BiTXiChixFkH5yzZnuvKMSGdq2r61R8cesH0BHlRIeAcSeNuNjd7AZTvU
bInT6GjUe0kw1LJ2NM0C12K4fqRdVSZ3Zln1zcuYjjm/N8VRx2l1ZtRFU0AJuyB+
cQBDeLNE0wq6Jld7Ed4LzElRbmi7LQCqOtQBAVIyFeoW8pP3dIxAh9hXHYccM8CM
2KU5EsS01sEZuy+U7HLc+3fe1IuJBbqD/RCPRF370ObJysR+cbUiH2pA4HoVrltT
Dhrtp2uv81rCfMa+NBkS6cHO7HqOcmghe7+yDprdsP2A4zacx4BOd/WJiL0OZxAu
+dBFfPpnSJ6W9CCJjaIjeeFa3U5tEYNTicDeRyOumuDNM6qHD7HKAT+TFVdEiJ5R
CxU0vqVWtY+3qfaaudSZFtTT5YHFbRSdM09yF5LALZzc9513mo26c03DoD2lyydF
2vmJhJ4YRW+2dEncxbMerQlRIhFYYOs4WYtjOCBX4ar3j37i1ebd6rs2WDHWckrp
ogOcWWyjWWEcjmnkqN4sE2/LpvyWs3o9sJir4gVPM7Y+pYD+j7MTT4TNfTrYe8zJ
/cv2HABY56LB0yHzw9zo/ixNvUftQVviKT3XeSx+8+Q++PwmA1F6OtnmnXFcgZfL
XPrn5xGmkbEUoSFylSwm5UraMeaEC0937+lEzUxczIpNIdbrNnRGg8JML3Pv6w0i
xklzbg01tSuaMwib0CU2izUOEkAgCE+wUtl8KtjjAv6at66CcOME4usgMaa02FDA
HYF0bOHF1mDcwocfDZXPnaUubPDVFvbMf/F+yzDmtC72Oy4I+/acjToc5L8yijxh
V3GTAGb7jowFX3P1zmHQsPFSZhJ4OrZuCzJ06W+veNOVEBTmvsC3v5SFgD5FP6D/
AN2wa3PWrbFA+iEC6HZaDjC6JHDH1YX9Q5Zxnbngkm0ZJp5/6QMrBLd3W5cm6elx
uFQuKhOyctjS1I3sW+Ccy2Ukz8V+4Yp/Q+MAIPFguiVcqqm9HI0Uq/jPm/F/hhXq
6SEVQGAk0RzVoKPIDyrQbAYs7oM+IBHX4aefsipxCWiI4o6jXP/CGZxuwKxNjYXS
OiydMuSw5bxEwLpLkqWM7ymGNyYvnSTr/gKPve0Hbra8zJyeh9N2beHvLC6pAKtH
W/fwXIHhwgwQrZwPyxi5zSgfG2uIYLUr/MECoYDMJZks6k/EIrv9UCH/emQiEEPs
Gi0PDrdFcI8Efn4r09YJacvKjHYx8fbHtEYp6RkB9ifliscUwoeJs8xo4oU4vvYv
yOwh0MfK0rrTS7ipygLfO0rHwiJbwQFLwWB/Tue6ETbD9++QHZhzGBUbWQKBJF0g
qyTaeHyEPQOPkdcqCMznWwxHhNUCnGc+T+LkQmg2LVPnRoplMOE6Wk0dTz7LZvT+
k8aBYKzwor2FsiwwCytPgcLzV1jN4whPYAYgFiK31H0oD2qDTM/qnmJFC+5SdqIm
4g4edCi5JngRtZ57hXizidH5tWyNz+RacVgsRWuhz+++5/vhRGd4JQ/D9vbcd5R4
N8pweEJJAa0P8U4FFJhQ1u1oUE2NuxY0hLUDBTDw9U+LGg2DttZdRTVYH7UaEfaP
HnbOmh0/gT+GqqO8plxFKYzAO/ove+fc3kxcqrNoO7rgVEbftAaCAS9mFsCo3ibs
yJJLVcBOCTzS8SXqEAmenFKCk82TGl7ncH9w1x0W2iq7Llirajd1XeCYIA1xdXiK
2J9814i2n6amKp0penq4YPdnX6NTA+SsN7PXxkT1uHV0CIhxk77YU4jYDXSnseJ2
ypy9hT6BXPe7dYoWD9f/CaFSO4Cv2t3eS76WV3bXGeCXARxSlboDdxxCPg71g6xz
2LbdJhmDq7l+ahBJYluWQ5mWYN4AWLKeJO4lcbfh31CR1GcYOhyfZUNbEW40KoIv
Dk4bj9zgxgARhfORf5PvL/rK1T506QXh/v8cBLRbQ9y+k4o0WXTX+Md7qbVcJRiu
2SLnAZiSnFNz4KnV1zkqCqUqKRVABQmlpDANg4I5IH/34BAnWZEhSOdrbKdYLTU3
eMiJO+z+/u7YZ4TD0V/Eui7tLQwomLbbNAtPWv4U2hV0nxEZzdmLRtQCINqkLOzO
67T4pxdNLOkuBRRPpeXS0JxOyggT58pzttGU8iXbYe+OR8s3mbJHG7dGSKwvrJiR
NlNYIUSozpO6t5uCEmLb8ETphki3SL6KcSBnWoH+4FvwvXFovWDA++hI08VQEzed
PCaYfG4C3imFL+y9kVF1SwJq1q+pDzc4Ve0Lg4FaBRrLRwqbuHnaOR38Q6Dmark5
g3cjOWlph9PK58YUzftP572DXdQkf1KfO/ZU30ddyfnc16xALXxxeHtaF6mCbd0S
ClFCf6PEj9vZe8Eaf2hB3zh4fBrSkVSgTfGTNO5CI2OuCqcFk5lY9KGaC7LSJQV5
QK+FGrc67M4vagJvZjSWQ1pbJ0rvR7LD2qkNoqh6R5SzC4OHnBdGWDgXy8yENBtw
aZ7+D6EB4SxW1z6ONfjS5yCtQcs+zyxeU7s7yR4CEyyn0omGjRF7eGTjGzhVaXgX
TSz7pkSKct/w1hciw9p5ZTynjdrU7KWeF+Y4TkHsu752O1NMC9NNBHAYk5IL+dXE
mL6a8LzNTVZTLEgOXWuOvDTfJ9g2LJ0JNa5DUSd24N0IAwxTLGR294BuTX6BB4DZ
tiGGaeMlYErJP501VkTWef946xgxbVlaU3o4Kdz+4xh0t8yZa/4z70qBRrVdAv+M
XsRum+dQrr+CzafI5gFJBwd8TwABEPR4kQIDBrbOOBB/1BTPQWX4JdbJz6k/lwlv
QfysMe1mWi8dcJbPeX51LuoTF8LT97CEymSB0RAJ+M5TFBk4w6afSBWFUHXPqfwG
ZcKlXgsb/ECHcjhX1lZyf9NU7iaP0UbnDL9OxMcvAvsRsAFpXFkHWkO9YJpPLXxs
PqVbM9h9FKJNackmpllh2JjCiPxMdCokAAkNb8OVJKxn4ucX3bZELveejFsaIddI
EYRMIDfpWKZYjxoc7NmAm1rfa0X8DBYV4rQs0Adq8ScOhAibgPopMABxwOW8mXkO
r+nNE9btcUr//7en3Mx4CuJrDdEiGszjgguuzJeQ/javAj7S3d/TBMwIFDfp/0n+
oeosSCAWYWXOXWl1BAK2Az9ON5z9eAhXiYi6Mj3n9VegPU3URsGEN1LoEnlKah9D
4nuKDRjftbKGSzcLKVh8jsr3TbmixWQMZRSuRzjehrb3JBCV/DBfsjX+DzBbEfuf
rHzA+fpc0edhtDcD29LxEtZRZlvJiv4BZsJhJ9WIwtqgOyyfV+TdM4KJtS1XPCvK
uMMRRkT849iJNYwcEunc27aRD/qYnqX4BiTfbJ7tvqJlDUpVUARjfnXcyZXgBi4L
0TtCD5+PC9t0X5kXP+zL0DxalU8N3tMZNj1Ag6YiOZ2nR4x6/qMV6zrjsCHeqS6/
AoDoAm8plbX5r3RAekF8Z3rQ86RcacxV8dnznzC1YUjQDwv7Q9usnII0mvWrH9FK
xetnnTnurI0cf4lCpUPUHh35Q0UAKawR+nb3ufPs/q5kSt7Aa3kKxV+aDamCTfgP
fAfd1z9i/EdGOsgXQf8OjDYbnH0fIEvf64kfiY6S1Fn/mTXeeze/FYpuH/lyVnhu
AYWXxP39Wfz1eBbiVPAYRPQdqU+VMybbd0cUEvYtmXJFP9x59nyPuiLy2EpnuSzM
eAOyAYjKq1Ez84Qum0GH3OmYNEHBpBegulp+fYstN1Z8/UvpdKHorE/0tz7+JqA6
eIJ5XWRCF8zBruRuG/4BWIB5JZ4ubk3pY6VgRcYrSWdaKnyMnUYot4+KYvkUShFY
9oeVPlHgTUG0aRAO9UtHdR0B8ekSGKV9+1WWrLomU2M7RJ6DDIb6JWmdMkxj/T3e
xvi69qj6q6LrpyHpUFyFEm3I8d4e9Co3U1lefqTQAzKjZVg/fhUZw6oHCLAboGLF
b/XuFvlEquryQuZwidlAB38U42zNytz73lvhpOBZ/xIneJsMplJgNCtQkzt8NVwV
jhl3nL5VK9jTas9qCic0jVDG7k0qVhddTx+C1S67A5pduqLP44c2j4XkEqEg0E3D
giXNF+c1qwonxHmtQbNS9CLSPFDf8kJtlClMedVeaeFfUSuC/2SnDKWH+CaLP5B7
Rg/FJ8cuOFVfX2Kz0FNwf4i4wBcHFuSH9WVHPc7VWEiJO8sS9RIr6gOFqrtbbqmN
mxLTGWByFpFKkAu7xvSSopoE5/EDFElJhqtutGsnw4epJms6gV9egKGGt5gRJPt/
rvxHt4tN1wmk0PWa970MguFZwF5rI7rS390C6W7VWJnpHmnKsRqNzaa+zFBMknfa
yqDwZCBPKlxDcEcTkyn7spunhSv0SYaisiRAIuBgjDrjVLqLTJB53xHPfmUWwrMX
T6stJPoI45Ogmf33xqcRZ0FqDsqZk/PfN9pqWRzzGDFgVrNyKhx/zIUaxC2AVU0y
L4aKoqmP/RNKBNwjzgllh1v1E6d2oXLWC6Y1dPC+qhbUngByBHUwflnajmw37DD/
c/CjVt5Brl7KUXcKkQWvN6phsYQwKy3gGrlqgbSXMCtF4aJhfjJaGYrt1e+o/pom
1u08nU9Nqi1emt3W204myPsjVagJXAu4UFZFwaFUSMi/WgI4hkHjBLVcR8Crz8i3
2qstxWaHY7xCEwQI5DnVXV3JTlqDfaLnDHztrO4CGQ55kdmnQNCV4nHg43d2zpQQ
x+LHyVpiffJSev+yOaTSkUh/kMs38Rb/mFEvpGXa3YMmp/3vXBYP1wOpWQ3VxmYq
RABSM3NI3cqrSoTGLg8p6A+e7+QeuqdixW4CcWwCIRLPwvyyjBCjsUJQEd6G06e5
+6yhfK1sabDP+Wom9hndzFc+9zPTx1IO0Zp5ZpZQwaCqmViFz6wuJgrflKEQodvY
ljYFiegWGy6BoFmFni4B2O4vp8vAa4fMvT4DSdFYwKixPl2NdKsROjpWBFnsOiHe
53DSUhuW+8o4Yf+wwp6qkmjRQic81wtgZCJwQXUjwHWZTYaiVxfguihqdeUDLBec
drSseATs+bXol8h+uh9kRhJYbUUWbtavlDcCDriNGe1fAEYSVOyEn1+n51cq0poU
uM/EMwgcYDS6Dc3gDIGwP/5m5dmaozZl40KFsV96jzR3k9WU96ZPO/tUZbmRubao
KRPvND+87sJRDsXQZ6yMwMaDDFQI5QR+PIwHaWh4QAZYSxvydKf3o2GdXWglAaJh
i7mfr/esu2voJCOjyZWhW1psIkl9U1qwRIJ3J8w+TLBVqRFjtmf23K8sBGWA/uk4
if+uJvGOVSL7t+MC8ql1GgzXe3qXkdDg4UApEeIp0rCMvaaIxUD/1u7uXHBabvDW
lm3HWM+gtxn866cPjWOnyX0bUO7u2zXncS6/EJjWHjHEW12j/idIga+YLpK3YlCx
uX2+6kmotHMboJ+00OosDjEZGrzN+DEFkKm6rZqurV6GAHtX69/w7ez7PZX3eW/W
e2tPW8y8kZkOA20E7cjOqCm1H/na6yG5plUvuP9HB4aG34/rupFqBf9ZNYvD2xyH
818nIPVRYQQIbMJRIq5qAZvbo7b2yF56qbsdWENSt+xlpsPBH+lmfu9cCRuPYAfd
xgR6izXook4zqQ9tk356YKzjtoDJ01y2F1ai7TYL76/CrizIrSNZpNTiegFflzs9
YkPcbuno437mk6X6h/7RMauAfDPkNkuN6wVgOyJjSH0vIeCFxhto65j26P8oK2AT
NjvcVgRK7RQz9qHyYYYfzr+oYzAzYEzj5tJ1Z5C9po8XGuu48Zpqj4lxVbAcF8Q/
C6uWp6qw/6rzYPw+YOn1s3V8vrAtAhfkkGhs4J2a31gvr9FXcPSB28BgZFKODZBq
AfsUzAT/fwhuGaWkwjX6y2+RlGHjBuughv8F4zEP2PzdI9fdcgrJyRrIHauiwaAW
hsWL+fA92TNjFre1B4o3YOHMYn3c6E/3VP4wRjCoDeQv16TkelsZeUHF9HqJhOkm
IOvwh8T3WA1BtgFvbpUNgslZGrKhnB9rOVsn+RLD8khrwwP7WBSZOIJExUCgS0KE
UYdfJAebKV6C0obETYwWwm4VQ2P98/ccK+NgaYReSnOnqu6+u2T/sigN5ye0MzlE
TYmZG+kQnvV5fA2SRt7l8jt+mHdM4dZp5drQw8Myvbit/tu7A0fMi7lAdieZB6Si
DXNhCHnnqjb0uk9eOa0A6FCMCP36FR0Lm1+0tZv/i59YGYTieHU50AQC+pfeoxM+
EJSEUBddexHQBtAkRYVnNs6UDJhTwkcD/nt/NvyhObFi1p+Mbf7XzNoPJqzswHAC
J6QqR38LGUeoLVy3+VpJHkngqDzVH6oxbIS5tKUs3yhsaH3gDjE6yLnADXfjBzXe
UATeqDNxbtPnmHOWjrfXRaS/SWbJHa0J92TH8BiE39UfYUHE40K7rKdeu3NT4K+a
9rjUscQ8UldfYaC/+w/pTSttPryCq8KeMJBziw16nMokEHrMHLpOOjY5CN345+Yw
AeE/CezPiEpL/eDCh27CaEL9YQzXL6bmhVGO8ebyRHsGcE9f6uWrYSb18kRibhMJ
HdUpo6IXWM8YnydXTEEPCJXlOBYreSeqkE/mXC5n09WOVdl/e2uN1tW2JnjmjrJO
xXJbud/uW7hcPkDQt2k3y/Zui3WuKOw/xHjacxtMBiFelZSYuL2zNH4aiYBwdy+I
oqRHtjzK7pglCRJFVVa7vIR/r6d0W6YnxhRPZWj7lAibOmStm/PJA10h14TP/tzI
Y92ruQ+xONOIxudTRD9sGg3fxXNspPbEBY68iLGvFmnpBhpULI1gb0MgPTwv6/eY
YtlCh69uXodkvnw35a9x8+H5snK7LAKRpyqBtAtABoat77sOqgCkK/cojaFm6CRh
rMaE7VnyjqtjTh4Q5VYWQuuMEfZzxsEFv+/M6OZzbkdUR2ZliIyB7iAh6ruG54fS
tSJvi+LGTSfaM6928cef8JWsig5sIN6Dy+2oe5nguXoG2e1x4l/G0oXYUBUng9Qs
ihl5Y68wPgnkqoqXJHjwnmduxEgPOXTw6irEroyOcAp9h/vpb6dS5d62QuVPMXWT
KMjoV3Y6SgsSWuVwbdRyQUrRy/UvJojCth6chUfh9Anm5DIm1sMzVVQxlyYv1w//
xNBTeU7jXAEr7vrESrxo1iiRcyje8YwIC/En/ECQ1IreI0O5ENNbAEZ1IJHWMUe8
dhZlmX2EiZvj4BR2uLg1q5f9fPvnhTxR2tgE+s28pzT6uefj6jI9O57R1qzGx8ll
XM1iRlFN8HihuYsmUBFieS4y3Rgqkc1aSVW9pkAyxbtd0vgkslHdpxuBewsYv4SP
XBXEFYB9Vuf7MqBM2Z//2Sj2OqeU1PabJkzpm8oG1sDFH7sQWvRJ6Xbl90XSFCOZ
bj1/f5CJ4tILr+8ZO0IqtwfU3TpuvphiAMXgiDCGD2jPHOmBAvnPcrWnis3gcY5M
HVzZX8tpY77Og/SPdsVzK/DillLW+rQrYlWfFG3IqT9hQXQ8J1pFSIeXQNkBQShr
oQoawY77p9YnmezvF+N/16tHKB8jclt8kokYNhQEs8sW77mwj5iHV9CM7p6tPff1
q/YdmW58jTkXO0P1oGEGvJaU0+s1DsBfoN/NJvlEO9jR3nHrvLHWyAOlG9fc3C82
fQ+MDRu6/WtXclXtQ9bXPms8UyF4WS+hJu0JLYEeOS7ScTvQc36x1UF7+MmHMlTR
F7OYGyAoyHBoSbcp72R5bWUdAhKAl6J3nesg6CUU5dOlQG8e7e5VWjkKtpkpxFcu
TZ4QziYlfuwlV5aP69mlqQvquKj3y/P95siG/rCmY7v08fKhOZD8NHXjxVt3bgrp
MaHkHTm2vU42iO4nEHvtjFBplwM4pHpmloBIMo7qnqEo2qB18Mo7RndyVdhpiO7c
P/SlRjRr49cSih0CnlTfeapGx0MAP+zbY9N179838qqr2Szvox8NXQjisi0/smLW
1eklt1TKH3HfKFJWeDP9aaNzT6P8mEhKsODxUbirJLA2WUCEJZ2d0Cj8yeSqJt5L
6D0NzlRezfLQ+SJLCI6x81yy+ss1zSk5MOcA0RIzFAcg9A0jibfPU6qnTLAY4G0a
ruLZdYBQo/YklpFaYQlpCL9q6eA/TauB9cCqLVI56ZiYV6HXrukd62xlZ+DBumB2
4PuEmT8QkhxEuFPqKhfjfoYDU365ETuaOA81MPk7oG5k0qVViSy+TAPD5QcoLhSZ
8zBUY2X/+xskYFnPsDQqXMvggdHoXQI/nbiT1xTIqJonacSmiTJmIqTY7+UsGDWi
8uCFQLkpBs7g8MBOIxcGmwGckSbX56X8/thEdq/BeOMZl5Mi5hmCPyOdarVPh7fN
DyI6mxKu2+rnWBYNSBh5ykd1PgMwOHIWY4HghZwda2r7Rvi5zblY/i2FazHgl6Yr
OZFH0jOUNdTlHs5r/kBS0qO39uXd+XjYjZAt2xcPWxT9nvKlab7/L/4otIJXyfbD
0knRSLf7+CGYq5sKQiWFazmM8LLb+kCAZJMfYzn6MYaVr+ktakspM7ZXW6zf3wt4
XKrT/A5x8eAPN+LTIz8mMZdl0grJbXgVHIJLTl59FvnUzW32orwP3SsB9Xfkd8Ay
JaIr5z2mwIYH8EGTks8HJI9+ayk04iaVwezzTa17+wrScWYStO7DDuCyNE9wS9tH
cm/Iuezz7+NQCYz7ROG+f65EQz2M3b0zxQQw27P23hog8GEUvS0LwBvysvI3XErW
GuVQE6vOVJgSG94Mw11bMcjIhcwyT1CCzGV/l1McpcHu6c9XqkrILn2NHg7PLWra
htxRXBfU6mAcbowRxWrqC9md8q0etBBK3qwubTiESsjm+xiJLIbHuYC2v7dSKj+Q
VGMGiBMaUBtvsEd6x2nH7/c0TMM/ujky5Uxlr+r1qiPyGXGpQlHSkcrejhFDafuF
JT08mE2Itz6yGRXULI820bWpGcs6VWjsmMKFL2REvZ6yHditP5KkjsuTtS0WB6mz
iO5F2R9BBBYh0ZG8FwixqVTbGZP0wT8lLYfFlKfu08l2wR/tFVof0om1kULNrZHK
8F1Pm9j+yZjS5rD/lIHDNgiAwTgXyAB4x1FD6gd/4Io1E3P6xhsxEzhj4XGIvfTm
B7gHrjT4/2mmKhj2B7ImmnKKUmuyOaBya1Y8G3jeR65T7w2dFsa/B1dikIelgP0S
LIzdRwCzn41l05fwrl6a15lhrHBL1tlBfq4G/gjQnn+75/iNT0dsHUldbFr1j0O9
HeSISMCiRjSzn+Mf79Yiq4kAv25Gg7DqDRf8zJL5rgYJ6mKh9qGTCj6bgNfqTaZU
LDetKLNJjqUSP9W/IwZS1eCZ8iBmumbuj3Kn8gmNyWCRJ6szqN1QBWhNiHU0LXdH
lhHHf3mtiTnFZKeKOWr4g2oYu7sw3zYe84XfLs8J6FH6AEWZ3IOXmI43qqojBSVQ
WOvzhjSUmo19JLQORttbMPWDuL50IucsjN5IWljsjxIHerAjG1A4v4KzBl3BUxDn
aVTJHlSYEl1l8f51DuRIR428PFtj7AGfSFPGqOrndJLuw0JyN6sA1frXrpdNuMif
DE4P30K1F/6nBXsBeXaqIWtQTD5bnd0f6hdl2VwsGr3I9p7ltWfJegIBX3SSVku4
mCraMo7sdDK3wPS4TOi2YvhqD7cfpjThJdqN61IvQ7xU7xTH203QCQifm/awTB1Q
Ygo/ZxghKFXEeHvhIa/SraShAxSCqojP4NWmkyioxk0N44yDY/XA4ZKF2CZgRnuJ
4LN1tLPxv43iweKC4OgINmFlJLIBnjloHEYF/9Nffp/B7FLv0OW7xJ/qvJvOH6I0
GWcgD8NyrsJG4BkmfvMEcOPTfCAYO6azytzG/MUCObhTbkF782I3EJk9qm5Zj5Di
zv9OftC4mdVMAtbFGr+OgtgYAHpYCPDcdjAS558MK/cbXHd5ZfopfWL5BYv3iabK
EO/icdnsH0LaCwpBNyFz1lnKlSF6kJz1z1O78svsdjitgfHUuc9UgAz1y2zs9VYD
/QVPp4b32CWBGvradJtqFVah4Fxy/U5qiWWe5t3YWc48EHx4Un5YMwSD0E5yZtuP
yiDvAxyZ9Yj6O0S5pcEsjZ/KPCmbFeI9IK0KMj8rJ0Q2AJpAcUv67RxtpvCij28G
aALVB5oS7o7Ivzp0FWRq+UVEJPoMp4UTRa2zpS5I6R1x6azlMeGSQYzz9pG3PUA5
LYkG/cAzEoDDYOGXckuEhScbg6evtRJVLV8BQWiEnYQFovWSoaqCoVq7VAIGeuiZ
/CRk1JzHQykpO4NZkK8X1q6XeuoANTe9W1V3mcQqygD8AGUNPLA9CsPZwpiv+zH2
TMWQRCelIi9yh534RMyU3nfUjy7v0IRDkc/On5NhD+hK19MppwXCLnF8nTYfWNfz
aW7dgmPsJfdwgNddzAgATGCOqYvz++4ShF42INdswrPR0ZrmiXeRvol5zB8HQj96
frI5bHFowNWfnUrbWH79QwekCla8Mo1AawUJa1f2cWnLFhRHDwBuNHgeHeWnkgLi
JT3slcvTkdmuNvOhc8S1S8VTqBe73zAjkRcDFJvmHALkHVc9OdQUbdGg1kmh4sdT
+kPYA00lKNSuiHFm3KeMRi5e1ow3eBB9BJDoy+OnfzUgarKGtIXLg/nRWgQtkID2
YRoqW39BTWcfDhgretvX5ImCkn+JnS/dO6JbvM3xzKc8gd0Q4hpav2Nzd4A9KdWS
kkE7DNfogf4cNr9aprXuvOWm0oIWJ2kBdRaOU1PzXi6DEB8UtltlrclT2sA+uLVo
ducjNE5O5ki/ooydlIkPn1gJHxLphzvtLtXAlnnlMx+W25TD2n08IJtkWfTQ2+ov
rGSsscMcmkyXOudSdewRCV4ysb1bKBiKYM6uWqB8llD2QeTLUYvP5ynsiWYCTksh
isqKrZEKSnjat2n7TcV9C6xBe6I5IkpViZmg1QzJWGerG0XN463+xZ5JTuyt+W7o
A/YSXFBOn4H5O9ep2agQTWPx2fkYi+/zOv3azWHqVOpaLw1xgG2hkOc2lXjgN1TN
FN1wY9BR8M39PT+8JYtlZQOP0WdJW5jRdPq+boG69r6a65zbjT3ZVTmSZ2tfJVB5
jXhPooAbU/o+GkQlTQDi/qyUsb5EbKZWNsmY10oWZ7j1JtWKukclJhXo08uhlZum
Ll4SrqlN7ee/dMIrNeSR1pjq8yxP7Pkhx7vPIliDkC7HGXtt3KH4tZxNKemW2kqH
HuH9BIfvpOhQ6PScIzsLlhfRE1NUJIjCmwzjw0SVepUlD/xxD0/Tv/MO9Mk2ebMp
m34+0kRY7MucsdvRjl8LAfzztf0VMJiFnh1hfhu/vwYLc99Qol/UC/i6JGsaA+za
uTu2pTDSlwtVrV91cvhYibG2ahJzG6j0CwtG8/gMcIhgFgzCLFYTVkBgoXWMwGw/
wDPIPt/wK2j1YhstGZC2Ouo18fp3dJhRHsZlnUUkUoL7QzNP1OMdtabHiJzPCBhF
TtjGWkLBiihqnDN0L801CTHd9AIEfu7dkKR3EAwIrp2QyPQLcQNxFie0AWHQdzDN
zU32tVvDi6i4M6RMtLBgqzGmmLKBKoniz4O5D/dyu4DvigBP82QQ2+FXELz6ufBY
u9D6UCwYdI5TIvQzsZ0r3bSFAyezae4ofwz3j61sYYHtWS2Uhjo+u1h+M4ISVjLO
pokrRgsMzpdv5F+u3Nb0FKsniz7jF0mx2SAc+x8hQFbTmuBsRIQM32F7uriGKVUn
HnTJ+fmvKPcaZL7k6ydAk3wqvMYT3XMzlSAiPICrf81y+bYMMV97bgjA8+OsdwdQ
zPEG/3RXlQNfJ3PjPFRtZN+PzqUv08GPJ2G/W5D3cz9QCXYbXxPaDcDWfvPLKBCJ
0OjDKhvzG39RBimwPDQAt2zcYEq7VamxeQ3UMwUjEK4eW8aFNkwPAYbiUkq2QVzu
+7xKT1AFEck9MSGyJvBWHIxRgKARU+Xef8/VADl96QnQh2vFL5d0QjBL4UXmIUIF
e0LNu7n4s379hxOcuERJrKUioY5JPFU5Wso1lhjjR2h/flnk94bYVRGhZmnp5cOC
pXj+RN0xuXRVVU1kKZnlSqe+i0xbxDOWs1CEOnJ4bajS9qw5FmXL9HPWWKlD4om6
cT3YM8RqDadcL5O1HvaB1LgeJAffGCjy2Oayki5sYBdP965qGWEpDN5RYFKuPk6T
eoA13lQO8Rr1y42XTiOJPLE9+LbDZowHilTH3X27rvig83wfko/0HQTX+a9hFkNW
Kb8kLj0RYCS6e5P73V/Pj1qDyj7Wffn8C/AUDSifzqcXNPHhQH9qjk3QyNiOP5bj
n3Sbq326LXyUgG+wzYNX/KuLGjwg/zNnShft/EfnVOtv4KDCWO8CiX0ugTjsjTHM
iUdy+0ek7Vlw/s6wFQgGgZGMiJyUWBmGAMYKcjGrkpCRnDbyNQh1mikN9zcWxNGF
yUoFfxRkW/zcbZINBAloFX8kHhFzhkbwp2fDh+7u+Y0UqJROfyY2WA+B5Xp7Do0N
wDMWGb2d1ie727/SnRHxaivzAQ73UK1ghe6ZvTgla4tt8thMA/vwa6pIkxq+sgPx
Hg/8Y/Ngryc1bEjZ3Lnpg+ilnTcKwuxyri8zJ5IKh6CdQ5mcOWmd0e9dkO61TG1I
j9gbh9wdKXBDKT5u5vfdQ7A8BzamkjitZh0jyrTs6VEezMX5GXnnPjlXjJgY2G0Y
Sal68RVHZYQb7sqlpusFQDTKqkSrr+g1I+Vdh373MiFmS75nfspkHhA57+vH/vx4
GYILN8ZFHjWyt8Kh3XMa5nlYUTRJWpsFOkJsoNQril+TIybZDCFDHxDN/DviQ1kT
PSurD2ygizsEf2P+IoZvFSIgR1VcpUXmjs+IS/cAGegX92KiAPcqY0Pd8w2QUEXI
caP05O+MAYlq7byItU4nevKzAkyGqNJyjLeGiVrapXyB+eRdV+9RpaWObXegrZfu
8l0Z6YrOrAkmOGMURelarsvB46hA+1rbluoCfjNMDpM4zpP6hnL4VlOijHjE82pR
7hFCpR0UR+0abBQoa+rOekFU3gV403mn8cFtswy593kVVwid2Wi0bWfaNycNSWXz
H6e1thnF3cCzVfCom97nq9EfnyfdfNmbRfueP2qMdLCWalJow/INxNVBUVCMGz3p
9m++FDK3bDOkPG9zOaGjJm5HEQnJNyQXJXgaHlTSz1QvJDXAWda+08Oo6ZllNWd2
+yHHH/Jze8R8P2DMkN7s22qZ1McSDQ36ggnXFwPv40bncQ7GTg83Pj3zOXOuwtJg
sHzzxfGeYYBbU1NLNDXyIk6uAGu9D4TzgFIM+R7E4ytIh4e8An2TvpsmG5seOvLM
kDmbh13OKk74qlJ43w2reJJfU1ZS9YmN8JcwKMOVn4rxADSKjsoZCsz7vD1FBhfz
UX6JWYRPPnukObQasRmOtTsdH8v3EBNlD7t+E2Xk5myAr0HWxoOiD08j02PL9u+F
iWKPV7gQvIPlWFwlxS6EYfJQeQWBl1BJhMY6YEvWm0Bd/UINndNr0QkH7MdCrut8
aUVZlCDrZiGPez4h6tufU1hurlgRR9jgk1BsOKufk1Sur+W1aFYKdJjbLFMxuX56
rNGjhTodgUC3JTy4GiuQeasSskJAT5FoefY6A7pwpcFGUC263qtUvqF1nJEgzKdb
XKJcp8ixAxmQ/541xZY28wdM4IaMEXxOcSHcne0AuFsxc1hfkIWaQeMmkLXteoiP
OTqyv+q3C6MsPOBJrMcfFNWcnD+v0w6cwukyyP3ioSTUsgbXznuPXUHKqT56Vueo
y2NCXM4B4zCb+Z8MBEuzLeyD1vb+sOL0qCw00JLIunkY/YXSGydb2Lx+PIvKFwpe
49Nkg6LfIHrdMqYC0kbJSc+Y7zUoBa29rzHC1DX/GxuZEFzMkMG0It8bcGRvuu9e
3eug9owa2vUH4GrdaMfy1UKmOkFVvqoTyWEUwA9n6v7XBClDeSLUMEv6bt/sg4mZ
X2B0SVSLT28TiA5oxC2/NinyCuVNUlrwCSGQmzDCTf1VyaG8M9ZyGw2NIwfblAtS
4Z9aVBGgz+aKOnE0FJxLJOtMjANJEuhOZus/dIabCMsvlTes2dHvqqKKll1JtXjq
ND5MihqRSDloMUyfKSyMUcL5hBBi+jHG5i7/DvqixzP3wDHmimxpiAL9y/dgLT8k
+krWmnUC/NjSTnxBRahYREPmd+B6t8okeTdzcfRexAqoxkJYUzaTTcA2VH++LOt1
qR5ejX2zXCEllMCGsy7Q6USK71gji/rHwwn9YhMg6G4zmCq59QQs0Ckp+1f3BudN
XZabsZAgr8nrDzkVnBcRpLnc3LU1lz5au9iJdZc4DhGnlFyrmyq8OnM/V7txinHk
noWpnOvtPHYbPiRhRXa620eqrVxyiQp9pGCfZ52l4/lPDHD3EfY8u3QoKlhqU5+x
S+aEBFzvE5XkkzpJt9ZiIYCIF2SjUDUaje57uZratWoK7glrHSRIERWXerxnq51V
pIN3ET3fd8R6R+nOLKcDk2uVKfxerjd4omOt2gBe1cZHb1mFf2V9wR7LGKEtlGM3
0bfrcJmpU5V3Ss+DRLVt+UY4BNIpl3gs3OzLDNr7+EwspihWtJtfZtOon4D70jBI
v7hiGc7tE01Cfw430mGc2ov0+3Rb0KxWdGYc48Izm3mzMYtAxDdpavbScQKgUeRu
I/Ofg5SNATBdNZknREW4+Y3ByRJt8+kNjWEGUbPm3TPnzMLEYZCrfiOhDhXY0aJE
4sfLq4XJKT8BcVvw1epm2kns1v+ErTBLu4DYb9aJxwrbCyCQiQDPDZnmU9kvPft8
woxYzlUT3es6EYlEMJSkmoecwQFzoApkhClWzI56Bv+6NtokmJc7oOgsHrY3KpGQ
b6WvOG7H/8nUBKpCI6fYKtlhAJMyKRArJG3TOUb9Hh61760BUeFcwX65b1OcAxIO
hKSsLQUz+MWew3gNg/UZ/bLvIjecQ7oxvPYl1G3RhotAIEkPw/50++PD/sSR9WeA
csTc9QlDK508gVDJbzFbUTeIezoLwsLcdkNIr3HuZe+0+HmlXs2W+IFJZWh3A3Wh
n21MDqkc/Dq7lSHKOf7SikGRrBn7vYuPOxkf0W5rf08Xa5fUNFuBhmvAm+dp9JrI
nzXnApDQdUJSk0lsI+v6nxxeoFwu2D9caMjP+U2eR8XZ8epLPiuw9ldPLMgmE6vN
v2iq9zR7kZrjhk4o6MQEVc1B+POHE3ora8yfrVJUjVEdiGed5+EIe0cyWULYsPDR
rHiuccSqmM8JBadTYWohDC7EKzz/YmAOuzI9cxsCmgawxEfB9VtUCTLj4PTkw4LG
HUCJHJUNULNUMDkh9Z7wgAxiLiUUzy6iaUPgbOVM5KnKSwPmw3Ats+1xka9gUYWy
oqvgZxwzls/OFveFIdQ15StmwJCsO/jHbEkKs0vtt5fDpJFdey9nWqp2vTx4NTCm
2IkVAORGWU7seuJiLeNJHS/AZLSorjaJlRFxkbII3FcZWRSB4wj8X5t77zHdXfhA
sw85NmKZcIlzvzho2dYvStjWXfB3qShylPPt0vTD3kNVtZsUSQcnnwLnVXiy2yn2
vEgcxh6cQSCIljjiHDD22H22cLfJjueQa7iNXSQ97b81haQJpzHQhN/TdVhaEq7R
PQQZEnAN95NZtE5th5jlIVCd8oeiwa52bX+UTnsSD6xHt18sSU1xHuMTTm0ajPFL
SWsmZygGSln7g0I2hgu8FpLfhKon4/abrG/d84R+EzZApJm4DTkcAuvXK+yfM3iW
MXGWAR/VbvucafehX4r9UBdFneeukSNAdI/A447RUDj+tzEplFDucCNzF+1gZo6x
VGHbx2nifuKt5NugrcVvRC+QCQeR6GljJm98oqk1+/Xgi5YqIV5NkEBp+7+3gPyw
3MbIof8ToCyB+W5BLuh1iX4tbfGDl3/nG2pUjMefze9CvVSYJUe9XMAJQv2QF9de
cXjLgjQn8eLgcJOQ2S/xVqHG5lLTC8ypd8gkcN7Px3LPnE+HnB7h7aHzsoan/lEo
5P0PK4Ti8LZy6R5Zb9IbV+JaWgYHQQpJHX3Oqw6iQlAaAQVRwt1S/NiIP8Rwz31v
ce6JkFT2GpL/gY9PDYpXVSua0Cvxs2Vzcet2IRs8XASFuAUb2jGNHUPeJAS5qgoq
kmrQ8z5wVuef0sMw3akdkxIeL4juOhat7dOuxlZusLRWDddBL2g8OUEm3YMUpbon
n/gEJiX1fw9VAVf0DpUNYryABTCJ+xSPUen8/5E3nUaogppgSwy5l7H6/1P2Qv34
GhasjxTuRjz9LwUAR00V4xpbs7QVCDAMa6WxieIhw7b8DjV0ff9huhOT5oVykBiY
/9NLnwVbAPD36fMX+FM6CFHvFcwIXOfkbOoZd3/78clbEDnE56IfNm84qet9gv/E
s9g5MVyPfxW/fdQaWA3WJ9vLQzbdsWsZZfocB+lgwarnfYSdgLD5bJF4OLNwiFON
PBYRondqe1lsTciqkomWZBgrLnAetC+a3PVmrcahYmM+jTCmAyH24tQKD+kGeWf4
JVvE8qybTNcPCZaawyxGf1uER47KJuR8h1b1cRkiyGfRqVbRc36gaYevVAmO1uWV
ya29y32dl/qmZHItDljGm0PXkoGOzbqidtPcJJv+XB82aOcgQaj8GgEcLsEBW3YM
fEbhst5wib40R86SE8IdmASALmBcPB7Bzs5Tuz8bVefUlDDOBmPG9LDH2iA1o5FS
FpzWiX9T67uWO8vqqgq37daACJOS2e5Pphk3ChTjpzykErAhr85zuEdDZL/Mjm6I
tMaYmMAvWBslwxzxx2f/KozpJYTLKJzkbFZoQ6QxrcZPxxK5N/djTytqCzrasjx0
uNzYziMW47dTX8c1u0MkZeufc6zYMdXqrZX3Um/A8ZJuSMMEbrqHtVCRGpMLAWhO
eHIHcaOWNpOxQNzV5B0IO1kXWCcV4DtiP9ndv5RcYDqRrxgETtW7X4OzI4hx3GLM
01Pe+nGOO2V2z8WM6ffAAGQH+stp4WilNgbB3bXRApH7X78Xlv7sDXvfk3F+mwG3
IHZPdBtq12yyb5BaomLHxgiGwKLmO9T9P1XNt0gZJ8vPz2eCshVh5Ep1IOCMNjn4
TZ6bCfYCVryvWd939FAhydqJpQELS30aSEsUZgDQNO1koZFeHN7wuznswavgKI5j
zDl8BoVe3DGAFKJSQsZxJTyguf0DzS6ho9JPF6ZuFou2USgfYNYpCMGsSzyOhIE8
QYJ9viF0RTaNnezj5YXGxEejkPyQAQ0Psy/hWcoE2jOYxhtXDEBMqiKcLe8z6LWh
YIt7zHb1msWyBZ5lSWUopSRsAvtzPeG3cDi6Wi6ZkCfOvjl/PlmdNPzeBo8wJR5m
CfddvECgNwQRDP+7lw6htcEIf6/dC1Nh/inJjFf+nHXgE0wy1tVL9P3cvEoLYUqT
LDHKrEmoBOiQQB/1fsCzXsjluj3ewu2sA92GIWG06NlKhW3kECCP61OLdHEJg2Kh
MzRYuCfq+rblU7gGpw6lxFHrfnBNp7KpEmI7XPjTlZ9v6sStIRdmlAFSzvyHNksy
foiND6AFtGgQMloKonpwH11KXNroxsup0FqRcXIAOh2FXqgvOlFVZHAzX8rtrOCl
Fj0Tq+CcoTUhACjOWBBDGgflNeyA6YOzrg+j8pVoan/2VFih46Lwa4v0TP1p0YS+
u1BJIjyg2TDCYK40WTjC0H0DRV4Yu6gPMJ//tVEJtsl0dq90bL9ICAM6/rVeR4ja
sFK3X0aZgCnuIOYBU4wLKYX0WDnbjE4eRuZMWIxqEtkNgFLu/79swSsOGBpnp3EV
mE/4jmH1Kraup4w1icxZRISdPqMbP7/sBLGtgvRNfLNDeBl8rhhfNCAQGNxz2sEk
j45+lRllkfuHC51XLcw6liAN5o2F+E33f5We4me7jTCyrL6YBi2rYOprZNlDRJrA
hvkuEgHwpYk3Bv841LGGAfugle8/UtnvcEGuowiggQ7LnFVl2mfHZhMMEZr2tLlI
k5AT19ETQub7gE7xAcVT3WkKELej3D48gEJviiQmtNz1FtXFyiVcNNkZg6Jjz0KI
MTBXCaIfC1C1EL9g2sqli8B45vwdOIEjwPYQx8bniW+5plQx4teeM0bbU8whds2j
LnO4q11dZaesgTjgwuFZ5o2As4holjz9UFeSihjMQxTo7T+uAsyUlX7u4/R+N9UC
HggcH87kpiXgrMzVvsQgFHCVi2NyANXFNnMXljuIEKlvU+WvW5t2MFLpx0Cfroxt
1YX/UdDNbcJZD7IJCRIiHV8yZpFKmdaTfXDauTuHQCqjLD0ZprGJogOlv6wVxdK1
xs7+2xtYpYquzf0q2zQQzCDSrUtDgn1DajhAs7e4p5ZIMOUw6mjIJ0s7UUaieWrw
/GRtylY7W7XV5K0Nxqsv7r1XTHaRhEb7u7mhu9/o8WxmxGN4r7f8lsSHr+SIVWXA
DASDiPbPf8HhcB9QA15rV95FWCG6Ee/k/KeHT2MyIUVLFpNMvf8KtxzyCcBJh76o
Ow0zvLm9qqCuao3WjCdtj9ZbPZmANV864FPU9jTLFa388LijtoeJKSeX4zPF4e/6
+4RHi38qibexrfbgVuL7g3FoXDSlQFPxiq+TKmKADNGBSymmZ6U170T9b/EaPD0E
W1stoO8fhmJIsvYzp2hFEKy8W8gHlaIJV6uu9T23DOJkX4l9Kpn3pBsarYrQw3tJ
gwL+osEr5mqgUbbhGFXBOsGz/gQbgDkJC7gW7soCOzmnKAvw9x917Bx1RCr6ZDps
0e8YDKfEg9Xw/rFEqbp/AedSpMK0VVI1eTYpQm9ZJYZJaktT9dZfOPhDqo/YdLgK
nvA3zhDb4M0/7gjjqTmM2eclN1txWblvenHHHTFdib6YZpu4waXSuf+z8PTRp50N
PIk+z+sWZLRxPoL3byEEJ+oGKN+Pfdt5vqZ+mSQOaERsjwOHpst9AH1niRhWo0Bh
PL+DeCKWe2mpB4duDFKI0eJousNHKU7UXH04hiJO8hytKpTMKyIeV4qdDfKfNM2Z
IpxS0KYYw3RfuI+vXmF9Gqw6FjNn6wvaWAXTghqESX+tpHv6ESD/rWryzRlQYB1p
RikHGGot2HAx5Nqjj/80tK5YLo7rpHAVGMbu426zuWHJ0TIukHJsaJ/1GDAHDuA+
Oae/LcnX0Pf7TnB9KavCj/jV+hC8rX3Leb0T/YM6en7yhejlQhlP+M48+xXR3uUJ
QxLtX27OX4ofU350wudY0jbVAPFYTw/FEWsOIdj5DNiG6oQLOAztE1Swl71QKriG
NMybGW6/hlY9zn1IVN/VQ7Td31OlL3Sk88wUXzMK3xVTdYmfYf/TSrSFE59pzUw1
wLf9jkSDCjxjl4O7+5v0wyq5BdCgNFinkmwLmZ6Vn8/80ovaRZkHmh2HvSVa2uV+
6jG4C9LHTKIg8NB4gU+a5sweIaknwG1xuwqyFAaRZPWtxfekZFO48rYMgi18VP3x
/ooqBkSepe1Y8z3QFVdfb/g7dlIFhCAKgZg6ICzwSKSVTkaeMZyj9j2Kbr2D0SSH
r6cIP8HCsmM17RnKge74rUW4QtOG2i9ebYPXrP4feggJmleU8O7NTNbc3v3dlDrM
Fm2dsR2552N+o9i/RF55KaXrsnD8XsxPmFUBxco56PIb95mtjCM1w4UFTZqC/Isl
60wXL8sA3JfSfzyRp5bwhx+MSz3RO8EzokPUdHzfTcvWkuL1Gfdo2gT/FDfNMqZg
+ObEGhiKcWPWPL7J5ysEtivxQ1q1keuSWFJKlOtjao3/cekJIGhOEmBWAp3eK2Nf
5ycJrn/MwXVL6p2MNyQDb3Lc2uzQTSF/vB5useEOG/PXBP/ETBcRth2DkCMTEtjG
kNR2+UVpbGwLJu3zTsyLElrWtSjiaMNT6eawQ0Cw5GuO8KI4SGPSMsJR8dp3Ic5s
r6sgDpFjxo9AxXVd1U9d9w7sEtGZVq20k6xJ0iXnJemT0Qs5PIrAorEwbi1W6P+4
SiW8VNEqfMuW+gYp+1Wp0MskUrUK8kswded85jaZj+xtJr6Q/IXQyK8TCItZY+PA
Ogbijucpa0yAqvXwWAfjb+eQd1/3gVjE8+wwwqBwy/DMDwhZRv4+kO8PfsRU/uSx
Qm31iX1vIIsMBPu6dvjnjnt8IM153t3Cyl6ODQdO+CgbSrM0QUQBza1eDeedINTD
iH8J03/mv1pqlKjmLbfao8xKBqfzt8A43RB7Baft2cnnEO7ucibSk18S0b3YUisf
Aslw7FVy51KjuDJgEvmJD7FdiME27bCtlabd30FIj8gKYkO/pXqK/CDgMFWuIySn
ug1WzIoNNaG88TgrPfN8DkJws8ANcoUnVn+/rb7h4eZ8pq79J0cWEAxCMTMEe+KM
Xb9/qQS1KMXzljZOmVYQwLYctwtkheIHz/D6QiPA6iFbzqlQb1TJflayH9pj9sYD
pOLtNJqoBk6i00oITcqfvjq4k1Ih3jlpH+85cKecxMY2mgb+VNuJ1EA5FiOf1zLV
RyKrAeXaAaQpTR45tqrxRLoyixd/4j5ec9zytE1Ju6T4dx+mUEeYW6SH9fEwN+Hx
lSKG+BMa1zZ1nEtRiO+vx5CspozduI1s0ODyI4WcnKc1JFLX8y2ZHSupV4SNLP9G
FZ2TLEmGmLDD7JrrS52CO88UB/OC3EL3ASttKfFAkIt1Lh4Upo6sxjO9XZbePtgV
hjGXHSp6AssxBX9nXJZ8gUH2aMZwm59HRXUUFgVLXz45p7d7VRcXK+0DY8P/0V4b
kgRGVpEA0sS7txK07De4tLPVY1bC9V+X1V/yehjlQBviq2d6M0VQIsbp/bpMPSi+
jzjzBG8TCjcMJ9eAiJyDp+Syqs887OXCnBfBbHho1vigZJ13SsbR8WlGhs8e2XO4
zs+paghhbpq5N9QwhiMIFmJGyXjB33bMjJcSccDA/9TgiA0BkxWgjN6tW7L1DiK4
z464ooxo8zrKsrRFMc9WXvQE1M8MSSxvBGCdMq3m1sVF6YC4Qgb4X1GXoqBA+7WL
9x33MltvIMVwbPnoGAUlGUBbhZ/ON1zYdnz8Q+HkcU68974XfyUwq12OadiFIymv
vfuYCiU0S2yGYUcNp0szhLqLJYvLyJquYWginTWhUrudJTJDemQwvspftz8emgpR
cfu5Nyvhe6QE6N2bkx+RE5tbZDnezWlV6ohWsGUgc59kaVDJOOg4mE23I1J5og20
xu6UrqDpAq30zyOjz38xSpCfwKTh34xJ/evnzsY7u3bHaeO0MNTst1LWYAST5iUx
KcQdmWJWgmH76Ct6f0UMKc5sLOFb/YtmIK6Bxe4kVEBCdd4RV1hdMU6jziHYduw3
Br5AfIuIYW+SPMOLRNHhFGs8PE/HVkGKLpvuTzim39Vnu2NFW3UVemoGuQM2eG+i
nZAQIXZxRPmPYpWs0FEGT63Onwh5T+J4CHXrN7MyhkmRFh3W8KAqf6507OQwkzAH
C3s+MIe0ue6gQVyUQNvBlVuzoYt4IKRoUg6xkObOz0l4F4SWctsamXb81G7NgCsQ
iY5oH0omQ9aRn1yzPwLEXgSzNlN2Wo3IWnFXfhQVoNDqeSNXEEXy5VhGeTWzTZ9D
pN1xH22bHZ1fbc9s+PQD4mY/t5bO2k3WbCyRYlwic7AmcEmB26pFoY951NmU0pmi
xrCasnCETx+tIkHu+oIbqfzWpc/hjqWY5riPvmMeLaKgg0YgTSl5leX3HWcLMcxb
DDsxZVG/LTjXXbFAM5zJ9abY+WU0Hx6qPiMr+U3OiRJrM0bQ8HFyKQvqyiAIva6x
ZrEVo4jcefo9uMCgw4UWaM407g8aKLMN5oprfmxFyGjsAg8tGuo2mGAHUx0PcF1N
Mzs+jbClb6aQnQDkE2VWUFj35L4QlQXeDjCeyfK0WEw80tSZNrLUvVQ0/murfDec
d+2ccXpqPpCF8via3eXTk8Q7j6v+3K2gkdSAUk/3gHkQRLtaElLFoLBHBZKJoyDB
YbgaSA9CNhuxBGupDLbxCvb2Qss12qi6O1e7O9NxH1MzcxFT1H4T+d3Y9GNJl+TV
LKMOERT/kNaYKANZ7S6+TU+RLno8zDfZfuZtu51C+Ac4kqwAPBILZOleWsLEDB2C
zT3z8sqH9mkd8grxSz4MaMyqxbmUFWjIfXgNKxgnc/p8z8wsK+XYxu7Wg/6aS07Q
Yju0WTgEIbvsGUk8YLWRcmfj1/XpgZDBD4A/HG/9DC+Xg0WuHlvU3WPV9kwufzB/
nvuxX7RpZkpUY/cE7vZjM6BhchBMXKdT7v/d8F0ecsmy8hJRN2yHLS/ieTmb7GWH
xMdM4j3T/0xfF5/O1ro0CD6AERZyAHIH+wN8P3AHsnOli1AwTBALuRptYqmXuEyU
P+2OBvYzHD8IsumF+pK9AVPgNv6pN8Q0k5smY3WeO5NTm0U1Upa9QQG5m4go2Qsj
cfNe7Lm/yKZdyPim5sMLGmodj+/zI5N+WHvqoALsaWgG3U28sWelX5uoFCdwbf6i
W/pBcyj0kz8XTC5mUl4F6Pw2NY8a3tsFmVOtuzTbftFqLKA2Zbvr72RUXM1U+68E
+Vxwkv3gOiqtGC9qAyW9WUR56BC+LAJRRfFBgR4XRe2rNSnadGhzYhAUfED2zDyB
n4g8iZqkXJVn3/0Qgtf9r4ql4z1+xmV2PEbqONbbbJEfGGLP1Sk0qxqVEA9qH6uw
4uhl4Cteb6ow/XbgHRRG7w03OYaBTv+jbmnvujKsUVD8FszmT4LIm8iC3nrmM+CY
q+UsSvtcpr1u/oN+R5rCL+9gIiq5cLX4V01TLORuFStADw6iXBDpsc5Hf8tDDJfS
hTpym7CMy1iM9HuTGweeqFKAPS2nO9FbyRumxfO+3MUKMyL3NYW2+uBkq0zQv1b7
RUrSIMw5sD3SkNHQOkkWcz3WFKNYUhIPeb1SAOxvXUFM/HpFJ8r6CGHuoWjJsQtR
k4LMcgg4k6d+LpGzmGLi7sfqxxCReQpwyn7HYiWjhA/+EoGAVs7XZns90sTbMxzk
PBWuwOpGy4do1gHOquT4uVr//16tVh2H4majhqYq78xdjWU9fKf8bkD4mW3LS9re
isu3iMcfAw6NgJ2w+gwq781Xd6LDQhIeFJYEF3vhMpQGhz3+m6GeFas4JPXLt9iO
oTScci7RsD916qhwwE2u+0LcxVIyh5yg+YyZC2ZcuZnLbksuCzgLw6BKhK7yfJ8C
/mL/9Lj3ovIXkhJX3t9bPcaU5QYGLwzx1vlxI83GFrOP1xBSFU0jlhyGYLhwQGXZ
Rxz89JjINBp8azihKFbl27tE5ZSwT4yEodKx2UWjs244EQ2l9r3iHvVFNj6rncn4
UzBqRkpSr94pVSKlOOQcU+KEvRsfpVbYEB75ibzMQdpkL4eyCvocHINMd3f9zkzz
POijaVfnAltNeR4OBkADA+zxLrmhF0ZPae8l7vTNdBe5x8nYMijs6znpW+SyQ7Wr
nbJoF5mPMZvcnMjCdv27Q0KGdHLQopirBlMYTymRZMKdpFxM2arExE1LS8iliQn3
ODDpO2xCDcYS9xs2iQu34Y72wjbkOhTTGvZcI4ymmUhcOwn2hXFHbyHxf5doCZGW
uuH4wf1kmfXDOEtSLiStP351RI3EF7OWdJNptbyiBtIdqF896vIHxNzhTI+yDQ5U
iQRh8EmRt6KwIoaSAvQ51C1DF3N2Altgo99s5d5nn0Vs9yjZ/QYK+MpLkOdHxHFD
Sr8bM5ZTh/M6mIO2KTkNryQmSgyei0VTFb+7SauySvbiPzr96JnKtuWznez2ETtr
uslFrNHSq50COv1ZKwymqfPmvHlob0s1j0xxThtNmGBWgeqvNcAcdPQ6yU1j14p6
vI2exAofZsbI4dr8fQAZpMV20xICVf7DoqxD5tPiGI22RSHmEs6OJxBMfmPuOUBJ
Q6bgWgBPWhGgn+Kmg5YcaiZSeUGVq9E8nFfbJGWGxgHXgkS2QSVQIdEZn66UBEd7
FdusjC0Vu6ZP2V/xadXWSF7WEYscMKQDejj4OJ7InXRrvQUXrGNxHEWvOh+weBWG
23U/fvfoHkUVHo67j5nt/IvAApYbrAs40KDdPc7/cQMLidLaSLZ6pJLlk9qNk5n3
OEJ8ZSWDGwpUpjH64QmO8bmuxua8ygEIbHIZCxB09k6L0pFPYY39cgTVLOkTljLd
DClbU31Y7AinFb+XY20L+rMRG+eyD31mIwliYN2dIJLVnwAkuWpzT0inxoBVP5PZ
QIPkqX66wT5u44l2WvAAiS2GDzbyHvWCsD7bvzk/WPsWGoq6JrFt0kCbZhI9uixc
0gvgrSIhLVypjk2HRzL2OFeShWal2Z0Gp4I4Pl9yPgeIXTISlh1qMiRw9rCoTVf1
qPA/MB2k58BBxCwmFbWKIMPw4P/LwlckvyG9dpGvljE9vFC4hvzrReD0I1sUm0Oz
n0kI8qqiAMm+u14YRddnvNTH3kCvJ1SJskcMDqhk5g3opsFRvtQ4HjK2FMCQJOsS
FQmMzCDa3FxJJAMmNQVQPpl717BOcez7YapBXRBT0Kj+hiR3LaISyEXokwlV3k8u
JPrfQbCDQ/dEdTxpXTjKcvls1EQh1x+oGGnjROvuOtoQOgD9eZwfG8qMprixDJA+
g+9HeBJ4uZfetiB3ysMo8yt4Ed1BWZDPyyQ5eMcYhqBe88DQ4QEUPG30CuREOWZe
cFWNVoCKX5rSnt0uSr3VUPFw/PM7fylXfMWJiE4zDa7QyBz29U9P649DknLbfklC
Lg/x9JEVnpqHL58BpYzzVT85scQCh7JDT5gSk1Y44dj0hepevMiKJxZORf+hlkty
gh3muYrg4UG4eHfyjI0JarAjrn58kfKgbIBlXgynFxnWELBnQqBVH+Ex1QARiBXB
sCxcIUysXJvpEFBkgXRmtFP87gdMNU8IcaAPeqxCP7Dp7JLr/w28zl/voUaxNT+j
91nftqUnUUuhAQLxhKcz+WdhHzjvdxwjZ27N+urzEhODrwF5TFwiur2PIfWUR49U
oSXGpMzuN2dfKY1L8NtPoK7SZwUBl1CkylJsFTb7azQXuF9s6BlTG2i3krlQW0jP
kH+IpZcOnuq6FY65paVufLqg6RUIFjOdsrV6KxRwsKT/5k7ksMt57d8tvVD/YK/I
LdtN3YGoG57u0NrgS43G9Drq4XgiKeh+yTo3pBmaxuLOMOvJH1UPmAvNCZseHmur
eZcFK3K553aWsGw+5AO0fcbFlZdY6eIEHBeq+C0WOK828JVUbVW1e2XmsSlUDW/Z
p4FTAF42RXdP+xykim0l4z/2tvSaoc8QRI0mXuijq4f3bXQvrSIIIwP9QU2JwYBo
fZSSfQfe1YUETKvb2yjCdd4DmYSCSYoFZuF6OQqRz7JD3e4xTMIxRIjMSYSS+By5
yNqGcu6s2kXt6EhujAVnthrmBwFCinlWecRFbPTONWFj99VXM5YFXivaFH05v+5n
sU4uH8fJwr3YwLeRaYjfptLEaEYX64LCbcOihHQ09LCP29UZQUmLyV5lUkBJZ/xp
960kub/vOhsYWPu29kwYQce3TBOvnuY7dMDOP6/fAniA6TYB6/V65kBPvs/ltOoH
lB9GX8Aru5mb4B2SmAKX6KQDZrzpRpE/7L5WndUF2veK/nF/NEnVw+5yHBnw6pJ3
drqoKCj7ir5deTih5jk+AbP9Y+b9z4xrOhILihaInIeygnfZ1rCfY+fJa5AjMN63
exZzEUX3RUsjMyr1v2fp7wlwRWgNTcXEX07pHOoOb/VA+zG69LnqOwf82LZ2H1RW
fAvV851Q5RslLMk3TTZyqiftbpPAUqk4hRf8FKDvCdIjiuzlwF1bxYfv+IiD6J8y
pVPyEh28y3nbsXOQp4typ+52NnCyAMBmKAZVpbt1fX7wrdtG1oHkPCHebODKdaDp
2EY6XiW3lKWzJYAOgUT7H1sPRu+zCcFoCbutLe3EAkkmEg25rv6bt54hXxCC3QUa
OWnw7771/lbfsoIo1EbqDKFB6NRi7noPngoRPmyVbKmdjTtpKHpmnijdsiSoqRTl
2K5mXnPSNWLFCKO215O9ILAoQlLP5NpQhETzALYe6HHqdPJK2/IPhtngrlPC79l2
dUnTY7YYlTduw+3jwKB9DfOwOcjZ+QuNI8/PrBziSDgW/qjmwBtRt+0dB/xfprs9
nRsbT5ae4WDNRbZVLyRSjy3CdKg1rMSHegKa98TpytOxEe3/ahrpo04y2KLE22dg
VSdAAPOoddD4FZyggjMKYoljVdgCwRroJWgl+no8uJrvsX+Z7OuhmftW7H/1dCAA
JRaegKenweTLl+nAUBKI3TxJ2z71Lvpz6gdJLq1l0ndVo1K6UdwW9nFrFDUvB9Iy
wWZwXHaN3SZ/1J54M5S60sEllOqtzSVH2RfrGsl1eSydqFNhb5JxSCqaXuNVQ5Vj
V0i7A9jPqzH4sbpopCmQ9pf/LOZYf3ZXkkdqeHx6Wq9nPoU07DxZ/bYI1rI8X5Xy
Pgdx5aH6PFwMI3pWve1/6JkLpOjDhPK61vkd/svpK0o/K4ZLonO/DV+auhupCKyn
GuStI8bWMOveh3wF7KZo8LuAxAl3D0Bzy6nn8mx1kOgXsT1lXLVd23jqatYEEBiS
m/gH7V9rKCVYcYGt8lxFvRj+RIS6G4KvfUVZ2FZYs+Gm4abD33w+Hl5C86t2eLZF
tlTNQPS6COjI6cvXWTDW88nODWs6YP2eyRdTSP8fdEhxV6K4368axL80ZjLMKzqo
PFxsPAvKt3ZGX6/zPkRxoRZCunSUM7G37409OJecM/IoOlE7apkcd+6+G/lTtFsf
xYXBr6HfWy05/PG6qrZJ76+BCWGnz8EvSzpDKuy5LgOToChwTfTp5s1OeqjDPGvm
D33gwm96YgfBHmqBY/JiVHdPvCsOsALQ0CCq6KFKbTDkZxkmysHjHLR7/z8zWgrX
IKndDYheEm7KSotKaeOkR88rRxefzxmoi7E/6WQIgERYL2DBVDv+Y+NG0d0bm+Mv
jAAvGRuOprzbVmj3Cp3Ch/tS0Q4QXqglza8fajqIkYQEWcAoj7TI4jpPwEyF83nI
evExQKQ5BdTgWm37rhM4YaIWXmQ+V0hxz9hFSuzJ98RjDY0QSNgboYDi4cu1Y0Bn
GALJgfBfMFi7cNZZ5FrDE0J3uGfUQBbjRmq7CEkAFhoUpUDIzM6q2bUM/f434WUX
esZA+OHjaURg+8U0Mw9y4DvMNH6TBQqgJ8LIT2zcAv5uL7eMhc5B0mYutiJdSSsM
3IeTIEBUaVrBuDauDP0Qs9VGiXXseUBiGae8OjGjQCwdLc4AltCoYJSLqNRy51fM
U3LGMGChK5aWIHggS7BGxGPd5WQ/7dHFLKMiMf5qSnNXKh4OBtuJO+IgHPTITv38
3tVGaoGPhvK1rnJ5INifSBPK2LT4Wnf+ymE7NsZ4ujqDHeEUO+BF/Tuyynl74oxN
Y/vuhnlq0zwHe67mAizq/sZXn4owA1HMcdCnxuVnJrRvTOM/1TNu7BOqF6AkW3pM
KYqjt0pw5K7mSrLZg7hIZVFASEcYWGpkKwP1XJ8oJvjIh159lwC/OVWAd19I7rTU
e6PlarYiBlHGbXUj1xREDLHnCFlVhB24cbuHY8Rn8EkN7wiJeemcMwpZ0yz2iNId
QYVmQTpUd6k/ppsJIalYRqeMUBKvOkb7AzRDCBBAd/jK8eFWNnuLY6CF34gi4KA2
AHvQ6p0+T6wVLHB3hoI33A3I9qVIx7rbyijPoZYD0MNrB0YCEw4qx7Zf2gryrZ2O
/fUwF1LucRaoPtLTeMj1ZHAwLK8D0SBBGBfEytim6IV6JcdC3IZ1+StYGXBWSnO+
/giFvrY/3iAGNUq5qZsjlxF6r773+6nr4LZBCYDdbDYbBzClnhmLwnRbNTzxlHq+
NVHwbCGWxQX+2jNquMnyv3JY6PeUozMhe+7PhxQhhH6IDV/WMKQVHVNH2z1L+S/I
DQi5bKljDoz2thWsMgRqMfkdfIXuZ6yg7yPt0iaG7y2m03GTUQ7ttNmZzwKtWUPW
hncROHU2LN+Pz2DF3w5060EUAWdct+PpF8VqvSyRtOQGPcp0q/QJpYwu2ThoPQuK
Mkie3eySRpn+HEGblgKi5uiFZLhps228UP8icfrEcOxz5AZBe5t4dobfjOj3DBjS
QxjlZJaENrTqFadm5w0ZwuCpSkuJVx68MIkd5PYvZoEQmgrbBzLM5Sg/bepFKq32
hhYVas4P5yNJha29vK2DQXj8NUtmvAUqVc2PW+lv6apJlMG3hmMhynjWmlOTKQSQ
5r+ok+8wfB54VUIFLKrXdBBVy7neVOYQGZ2keySW4c5/bDeVrDjssDxgXRQ+4T+H
9x+VTz12sVTJPewU/wKJSPOTuYg82O/tpn8tUmBaoLU1TCZ8uMXGvfVfdXHOwfQY
Zn39tWP/eXlZQWg1FH+U1fOTVcS0bDrE7UW7XiBBylK1RbwlVUIPLoG0pwcuxfk6
bpOhuaaz7+sSoc/eu3nCYp+GkFyAQxr94eruHh5NCvjM7T/dw/fdTUUiZweBxeL6
+AkOLnJgIPTSG6s1kooaU+tHBcp0O7TWgWfw/skHkJiU/fj8o6hGkbChFxILvp1s
lYZVHbs6hDUVr3iVlcsIFOReLtdyC+buo1oXSc0Ktn3AGPKeNROmhK8LBeWDpc2d
ged+IA86feVN9UiYc4Dp/R0FkFZenNufeS5vHVxTuFM57AvtkEjTBmxRiVfiiNe3
ZptAbXD3qJDofCweTHriSnSh3iZTeKxUwaWVmAk43s1XyIWHKCYrwwnI7jNtV3QY
us6l0BqeLdMZpEMvLCzzATd3H+Ew/ov06Gp8R6PNRmjIcpZjzWwhH9s4GxkO1uLm
PI4sQjqt5Zl5veTNw5OgyxPG3rAKb4NqgBWa76YG0TELt2UHv2FgzBLm2t+AAbVr
F6mLA99p38dpoOnohY4ZXjguKPgzacWoByAPfb82esR/+Q1osmWjpOqhncYGuWzE
2GjogGhKa3QONILRH2NCN/fvnEorFgD+0mJItMU53CjAbV6ERmDrHI5NRbWfDepv
/GzQUSZIrowmBDCUuQFyMKR4f5GWzbPimyeLbABke6bxFJpc5uyzf5vYKwU9VOuM
nZe8PRV0Rr+32/aeaJCJEYey1v+8ziXNm4LIcwHB8mY6DPzBu6FMoW/w5bRk0AF9
MM2t6bRGEO3a9VgR85zErZAZZuOBJ7vIXewq5I/PksnqSnaR18vhfOrVBXESfNlN
XrJVJgOi4QEkpxWd+qzcEc6c4EfoKmBuBxy/fR9tWK+ixGYfFJWZfDKBSAPJ93t9
umFPqdDW7sJ19GfshBUYhdiaXL8wrnQTlfF0dLGNLocwQgszxRqeWvsOSb0Zwsdp
fCuvDfJk9Gh5OPWZF80I513zvTyICbpkdEyf9T5RT4esqdD7dhtBYsRgqkpb0Ssm
Girca0mbaC8u7YjM32K6mcgynvo0VSXroJPEBPC1fcjzT1dcgTkgfyFEGyRphTmb
gCjNT0c5HdBPLwybhjKPp/oDAF172/qKACNHhn5mhVIUkHUlDTz1xKofPsAPMMAh
KrvtJpoALLal0eOtkilBGYG6hoipJC+oSegP6ToRT8X1QsptS/wCafBBfuVMtcNA
d4C2McZ9xxAxBpE0Yy2lt4XQDwiAFV6J7F13yedtUIqjzZrgm5XCAcvJGQVTv1Dd
sYTDBVYJ5P6S/QAtvaIvEhP9Ldv14Z78EulYVy1iqiOol7LTOZqWksWFJYgoIEgj
XVDBp25p5D6AqbOE9nvdlwFN19/QMMy04HTdj+TtnthHgL10Nmn3NYgVIy91gpI3
4jVYBvmGF+uzi/gnNtPRyVIO8c+H+a6k6LWXnI0Sq/1d92gUlD0uepxbqrKz8vA9
xk5P0MPw0SWLNsAlCBM1t/moxWfLiTcmL8LQCQOFdRlIWwtYmBUGlpCczgux5b68
uxexbBpzuC1yAAuhgMNRrsZNnMuUaC2BcwaBuCGsLLFVR5vyHKfTLtN0rirL3ec1
dHe7tN7YVU1aYZQpBlW/ZsMSPVDX6mYtAHQ3wIGMN6o8goxz5qOqZ3BAPlsD6stW
jOV8RvgamNV+cVKnMj90MAxzwLp3/hXFDWNbRQsLxk2i0I8hJ6BCdRr04JoUnaAW
VSLuFfAZBPdzYfjI+4YJTZnAAmUSYA4l2BjmXpDwhY1uzxx0AKtBta6bC30IxbO6
smBkE9Ed2bWopoHOEi/eaZR8tTNuJOrfq9h7xFMsCqDwqjHvPsmNJ7GGtvMI/0Fj
G49Gt3b6FtEgcbAg5IanIu63LwWTdK8xjvmTgs4vlh6RbeWJTdV7JGXIRcN8FpcZ
Wk7Jaq6YuRY99lioOoY3ZRrQqsagaHlvxTR/1wiNgZloAkYszrFRkk8bp67XgUXC
HIQHlVjlUbN8QAyMWJp+3bX8wtS302hovJzacwasdsZTBgzU1Risi0K3f5otyi20
UA2JoWcg1DMGJXhNRbOM3o8DB57Dfr/BjH+yDpDdy11PHOxbVgRilE1z23PdlYhU
4UIw2N+NXgcJdwJ344WIokc4ZlXYLUJb1HO3lWygbBcTbZkq65b9bUzOvdUb69PF
lZOI0LRXtHbo+q7pVJGFbnSHf9xjcaR2trQYd8kb1NSVblf7WYPzb+TWQEmZ/5XW
zjLk7R7pd1v4LelqO2xu07xu867Tmca1KudwozK8Tcwi1H9p9QcoJQY+QqI+vN/G
z/9ou3HqGCRQVHGfsyuLblQrkkXZzFPvhEdxhGg9Q5YYoaXZcdE47pKoysiT7BLp
iuVl6LkXp43f562cDv7f+3ayQrrjhw5PhvX+/FDTZH58OwOXqrmtX4VOZ5VX6Q/0
jk+U1Mx7HOxxNyUI4ZeHx7/+JdtVbDwxjZSQHqT3z9CfWeMiGJUacOhaoiCk7S2T
ek4e3CXuDOi9YcRjD63MtJ7iKURxVzMZabb6AFOjxQAcRZBDKnxjl4vnHEApKt7q
FScGpzYlDFz7+KgC7hSH4okeYXo4X+YgbqWGe2YCQJ/koe9eVAnMhKW6b/iQq6K+
uOMaKHTHBizqFIp3tKGCcHXKU01gaMCsxc+oJ9OfTs4V3bs0SUcpCG4O67AU8aND
GC7UVL/qv/MnP+Bsij/ic4Ic40ZI2LCbTkz7iBqrHtgE58jvnHvvlWF1zku3PYiw
QKU6DZ/Bc6naFt5HaEUhoAkOKJJhEQ9mVGYMf+/HzOejm4dEGvLyPz1SSeO47OKd
MO2qr9mII/sZwh/oJry/9OjdU4dhYgRYawfpZX7iNXi4iJPPphCACd6OkKSvfe4Z
Tj4/zxjuyvnz7ERmjFSTiZzHWDRfHPbRnC1bDuBHr2itRopzyl01AbzOJRNRqoRF
JrNWISHLUQSFl02RYVQQvXjwpb2WJwRg53pIFeb7TjpUNDzv4oQYBS/ovMkLPDJk
7mEVFdiZQCYXEyL8sG/i0McpEtizMlqwyAGSpo3ovlq/kWvA7G1h13w7rtQYyz8z
uqGswfG/CDK01UhUdn9TClih5D53olbfq07a8lnne5BOQq0+fuIidtBaWFLwKml0
0p7/eYhZLdxTycxkYpZOyyLvSJvVTmswk79dBva200BU2E1EA4Ijd2C6I7fyFsu5
79S5VrP9In/kXziQY8BPbqVl/HX4n3wUgDf1OeC7irPoWZ7XsC8euCGEZO0ZufKN
7/imCdMDk4zaj8pcXVB0G+py5234jryIScHNbidsMTXKqmNtQDaBOKPNccxYTEe5
HASrmxFiy9zLrznj1FSTojnOIxXOrcnn4ebkH2IGeS0dEW0+m5nor4ZSpY+iSapE
zzkHQskMr0VeAAo1dMQ67nMchEnJ9X4YGdyRRNdPuxl90Q9IqIAO+t2K0//vu6L5
62eHnKFDxosvsC0efgzGXaL53fdOzF092AuZYB7BXJ7+3pJqiCea6R1DRJUhaxcz
xowm66lWojKkJIeZVk6GVmIZgqlDw9/4PkWUEIk3yElbBT0Yv+vv/dW5ZrobOgtz
Y9Izyr1Y+APMRTrXzatXDp5ka/0gi5i/WHNMnUr9o3PKXE4Ke9Cpzdg7dMgofoSh
wUZ3+Wpt+CHck+KjTMuID0lIAcHO6prQUlDyglaLHQxOXF/ZehjkbLkWHAQkmPDm
w/MTQ2p6LSlD8W7/FiT/Ja3QwdA8XYdybGsHYpBcyQKkUWBGZ5+6dZbVv2qKKPcd
fAZWU3dyItzHmi/iY1FO6Q/wjK27RLnaH/dnEKdGb7a1kirfVE1SPU3uJ/I/kyyJ
groRyqOJcjksMQ72tYGaFFIxGtIhVx/eBODD4Iu09nDt7octXOsmUlxroxi7tgIG
/ZrPKAgHYgttqYwj2IXw+16aDs637P151/b+IsgISUvBIKdHyUgK9qbrCSAMbTKD
RtDt6CH1Pkzf9yjPG0cgXfwQuf+OZ7yG9XW4Pz1WKXT/Cdz0l9fUpZobeGZbI34b
thgsYaV364lCWCGMJwg+NVnid/PufrGM707iRoSwcAXyXPogtN3ef2n2z3zQ2qP6
bHax/3s2CHZotTXj9jR0G4zkxRuQfiP0Y3dxBbGM3c8A4GlZo1oaik9kTjgcPlvH
pfvTK4Dwgv28r34blrbsB2S7/Na0jieNL9NLKeX2jocZBSdfcFk+BFuU8MM6jkDT
QMQAYeTbxtDhxALbOb6vWlmOK44c8ZYBT7KI/yYvZlziBChSa8xcj8QQkELIaFTF
AlDXOqLGToHilRxHAZKdeU/fqwn57aFtzWelR1USWtGCWu8tS1CQqG0UbsUJh4Q5
sPCNIvSueU9tia+NZFcOn+2p1xkfbJGottNoCCkSJVLv7EFLoES1hwudXxYnvkTE
VSFz98QOoZUc9xFYcDqUpqqhhylSV/rl+/E9hnqW0hvNdtTbT+/bDANh015+3i1M
+o8vlrYDjlXYnfSQhz/kR4zO42fxCTZQdb21r2PgTQwhW+P7YbZ4CqgSldy6dBrw
TPPe+QH9ipxxm7yWioEk264LoKsn9M7yrR2P0aL1zZjzKNWfXqQO3lsLUZz+2tJV
KHZpQx03fhldOKj7Zp8GRI/A0Iepsk/J6qTteQAgmIq6HzDyzq9Ai29csZHwfA/q
yHwcH+WetifOx2WDxiM/PKbsrYhafMqu+0/t++/ECApMrQUgsFCzHe83A9dncTI8
VTkzmTEhbgDY8Dinv/i2TJG9ZCP5I15ZlcynufhGe3+1jTgdFBFKX7WskOql+XV+
GBoCBmiUCokM+r0Gx7pu67HFw6fZcbLvl71AG5SxTErF2F5Wba5rqhJBJ9j878/t
SMYCUyjkxjL3hzCQUkAngELCfGu6i9VuQ/V7Yq0FHcWgaUxiKlslkXFMzLQbPTJj
haVWGjo2sOc3/+q+mGMJRvsx6ZnogVwjIt536q+cUEQNGIrGJShxIu5j9mWP9mI1
8cfJBLiIskULMrTO23B9fo+2edVtiQ340WR1zp3ygoyOR0LNhQMwsh543wC4/DKy
ggoUpslpFZAN4TGvvHGppChKutUA0arvFXpDxppqpG4lGQv34TwrklX7JoHnuQrI
MVFh+/ERx76xqksTye880uejgVkUAwri3ABF31Y65W0CR6CE53Y46rDbc7Vozvyf
OtkY/7iGgKh4TcYrwQ3g8m6U6u8xE7KjVkGD3W6b5Zj0OEe3u6baBSGzNMYk1efg
9Kaaw3zOVN8umPFO4NeOwg99HpW4jaDi+VE2p+CK/7NkN/+Y6Yto7OFNGUk2WhNc
Qrrf8ZO0uIGGszPo1xixFlKL0hSuCbsWDB9SE1Vfx8KrPt0DjVedwCt4eRLgVaaD
gGeATKVJ/FdBYYvDVUsh/oPZ/91F7FvZINlVEhV1razNZZDLiyK7RtOTZ7cZ6+FV
uY2b3RH3nq3gYk/iQQBvteatcXguyKy9zNyedzLA7a7kauUab7DilkJv+d7ALO/S
ryQlef5ARmqLdrt7Kyfoul9Utz/7ss+BdbjDFBh3O+XgqWt59D97lxHiCGyL7gOI
hjnvMLcEf6r5pVJyntVnomiTnQjSqjRnZs3n+M3R1KXyDr91LIeVPxNMVNhfHJVA
d8CfLCyLi5tor3J8LNed136SDgRaqUFkpZ2uWpFHuuVFi3I/mNy8BO3uvQ+VYg0e
zYFK0kQ7auwLHaYUfymgYC6lRxPnpsQ2V1inMKWx1i13uYLgsqlOumdj1M+d4iGJ
v+EnP/zfgVAmNR34iY+SQIQa/JvhjLyan/EfxasYrQWbOa50Vwott664rHnwwebh
M2zmtBLD7nIM1gxAOS9s+Kmsi/HXNbdmNSga3bSuXRIbzYsikD9PgmyRPJBfWRUP
/Xf1psonbEd9fXvA+lzcMBX6QZbu0BdjOQBH0QQtbjpcsKv7yD3MLbK9sx3Dpph4
TYC9RiaaaDbRbuijBhtsiVCBoOCKHF20TSHnnEf9xdp9H0qvGHyT6NmfYn/9Mir+
IqA0PfqutA8VN1e+s1AluQtBlKN6w+4qKyA6nixSnMaJg1g7m7otl1ukKTe6n5/I
Y3oRHEFVOo2Cs8X1iHNROadgpbRw3bp4FOTPGdDMPBZHFr9kTydx9MeIPoRCscwE
yeeKcbnM/7rQLUxnqr0Od9djdkbkQ+K+krGz8O19c2Zm5K5kglhQnJffm0wuHx1d
mgorShTE+XHNjVXyoZlezUyz5boYrjxorfcH6OuW7DBeTB2v81FqJryG5/7LH8lV
uA6Jm5oRFv29wzPSuAgo3yZYLcKxGDy9fQVm8hlApB0vKhAjwoBVzhm9qQKB+RrF
4lmakIdKeodyfNaaq8ySqzYFMjeDocjbgxpHXYfuBDez8dUFhdpo/zIw9Vip1G+z
USd61Xm76eOiDmFWXWJLaNhXKNsFeEF6ZfM0sChl6Pq69XXFkawIiC9GDAQj97IN
q/DBkWhjcwK4xd7Y/7p1ID5JGrCUQ5E1P1/K3MM7Vakxr3SdDtb0vFVoWpRMPsaW
5MEYc26DW8307h/I0BWDFoFM+dGW4+HcVt900uZHSo7ClpMix7v4KB13cKggXtQY
MpMLmJ5m+ntWwPXIiTGqmm7S7r6eeQPLrYs+dhf4aDKPMDuEIbfNSU3NCTrxab32
Ga5UOpPCUWkLbTYqo9kD8KyFtZ+ra1dwS0peGKwl3zBtA7/C/3ANRuZ3xJMWJ4aE
GPPzkD+t5bvoFSn/X+oT/3cC4Dq3pXL5sB9h4SKIsuWsBGVnl9p0x0186m4q7WRw
s+OtKCn+RtOQSBkOP0kd+F2gv0RTy6bGM2NNRYYwyhHjNsG/ZgHzInY9WLAoJ/g3
TovgRkpmCDVnw+9wUVBc45IgnObB597cvn8sG884lZHPb/IqvgFGelyPfFp4TEt+
+zVJjsPdpoT0KfmjGTtRvA/IvkNn9r0X7lwATtXPnN3n/wo+aNbupWdU6TR2XqDy
kJVa7DLz6VPv9WduWo0PHrp1Mftiz2cu1SO/XU0x9ctu5W/1bcG8/LEMOlSAMYDJ
FX9NQrk+K3Ml+gGxq/ZwMyz6vlcaJV7WTYvMVqR07EjzBV+gNv89QxzY1LPjwQ1t
N1NhZ9NMqptUqB6AsLGN+UivxHaeUMS9BxEcwT2mWVMvc93r4fIFDXw9tiFf8PvL
B8BOD1c/HrKghp4vg2DoMVlZEbsTVzLrhrNDz6kXcul+WE6AanFUh8kniTjpWtzb
eVXj30pciX6ISHAooE84BD34+QL1GKsBTvjrn0NYdd5Kd6M0w9nc3thjeGcUtduA
RWVrOKdrsOVhT/ft0pFhn0X4XdHF0dcAeQmLoes0WA/qmQZV/V8fPUi+v5guX+b1
SrAjnnFsVVgiiJD/rfdZ6wT9svGvl+KD7j2T7oYFkPb3PhEgck3tTKAr1hR98mDZ
wl0DXDwNim4ttt+w/G49B6FmB2BB0YpvlaqAhCtdnaUk5REFOggW1d6gx2eUwQdB
k22uH92c0KmR9dfw/NaoaHeXWXGZge23oNAbMr58xq6/eEKRDjhjj7JiiD/EZ9W9
bP5xvGiVRlbtVBHmjS5B5ja4JiL/J4jpr8FEXZLVshzQ3tokJqk2psz+yKtoJZBA
2kA2gKuV8lPkFr2ezDLdFbzhyTypBwrdIGfiO6JxhsZe3QJncOtCwu15LAca138L
x0kMSwhvYD4bK0LQJVv7rahe/4O0m/vOaWY/94ei7AnIVdFYAzFIwFr3ZE7iWRRa
AAGMS6isVVws3nRMJ3HUdK/cVY9jLry4Q4/mYW3V1gezyWiLLTNEUJQ6wuw1RDKM
+pdY/k3LX12W+ZrPwiHlyZETHGcbNL0+kFMzTrbEjpJ7M/ZBxVyBe6RGn8hzxaQy
rFijBSpQlWX46W1x85JwYkqjStqTN9Pdof6MSa1f5wnsGnigfWxyTHi9zLKVQdOc
9g5B1g+R6XmY11wugakiZtTgnGQlRvbkL97dO9Cn14KE0qGSnW1qQ33TQ0q28hIQ
EYj5lckb2zG0Uwjgz0rDpEMCmijd7RDnrbLs1A1/Z/EC7xoQSMcCh1Vnk1z09Nak
JCs8n5/oFJtHELbnBUlc5keg9nMcsaVhuPA/+5i+hQMU7cbERV+Dxu4lxafpijip
RuOZnrVmRcIlP6VsC6JU53MqWCq/92RwRhaaQUBlGib2eKIRwMImpDSNz0T9a904
27RQ8MrTOatH0K4OcrG6vXMfQF6rP/G7LZ08Qfm77zw/+lj4HfYQkf+trFkOR7t4
t9K5+PV+ylZghj5EVnP6egiU3uFdsXISinee0OFCQocEmHjUoLZnxvJ7NIoQuT94
aqKUzzMCTVxCGYwCGjkdz/+hAJLa3XG1wzBmMEVt8JtA2j5VtBFYK4cP0mCxOfmQ
VpTVQx4j3/t9rI00SgdDHlDsZbYqEIyuvoYM14UcYUhaGMrLl0rfQtpySy6nS0ho
amo5A1FYHVm330ZPWDUqG5u1dXerlH0mBRhpWoVTugGafROvmHbpl7eNsSkKOCpu
2GnrPdIyrYFNxxPH15eETmnY9x77nxFIanXStivkdrxJFvBVjy5EFL3WKWIlZ1s0
iIiYmFQY+ho4LfILRZLFN2Fai4ntr8oNTk/Js/ekC6Qk6cRBkediUjgIl6tE9qmu
odRocmEPx2It7aKPFQrkBO9nXxyE0YLO5fkqZRKoHsAt7oIX4s3walkdtg4/h9ba
kc/K7+WrxRxK1khfKgkpKTR5AgImJcyd3CVvhmFGaEqipqwuGLhE1BEVcFdts8jh
H+bhBTQZiBjMF4hG9kt9KtTrw7TbewT9ZoQPRahTAthBAolrI7vhGSZpvYP4aazR
Nm/aEOAW60HhVOoiWQesIsmNK8gl2Unl2csTTNZRgkht+PAoONKxdl6jpSHyQFE5
L3FT5BEFmYJwzuwXSftrlu1hOG1Iul5ibUD7F7BH0TT+gO0eiONyYm2ZmqCcf8PX
xNGHFUUjHlqLUMQ6lZvlt95Amcm6eS4dmMHZlbkJdeZW6KPDxXSTD6IsjRRJ+N15
C4+XpW88RlvEChBObUuJNUEhSHw7m10F/Q/NY1jteZXNBBenZLaE5++Ck+TVb1S2
nOd3ZXYQUUqYbZRC5OQ4I+fLIp0GvZdpDONbJuLOolMhoM0YykmCK/ZV/bnYmPFI
EMPfrociA3GhcidTd3Oe5yrO03N7BeHu/9BA6LyuS8w+GbB0yKFeQpdtrqezfoEi
a0W8H71qGj+MLecVLG0GH+2EORKhL7zsQlZfw5RV5Y/gfPVI/PaCqc6JdBb74jwD
dxaLcgkGTtzPo+VvC/xu9uoGvEgzYJPxAIiwmWpc6NC48/RPN1IcrzrKCpUVY+Oh
5K58hPb2qrFutxkh2ZFjl6qyqStbPRCpwHjMfVuHU3lbqUBgayauKuxPwwq0tvou
o+PdUbYJU+Wx/Yc8dHTT9k8EsOvXEW/xzDkr3WhvSvYrx0WkGP4mwHTp91YT9G8c
qTxlR+ivXTSdk6tsrNgb2etHTm2KXevP+3TlIB+O10k04KGmrjs/aYXzro1P1slC
2MwnUdbxXE8T60Z/BSfIat+iZ09eMGDeCFzyom1/xD0f1l7tLHcVlyXd0puMoeHL
eh+i9T3Ghm7xYosN7tLcOm4zHo+fM4exYezH38vv9PoHk2bAMn8hLzePIcedUYwE
wGezdLRA43z2S0rzCKJn0LL4hDP0a01bCDybJFaaRfLZncgDEWj/TO6cQ8dAsgd6
oVr8X8+7BGTnFHvKxe+IkykBIbkr0FNMgl37jKAWKq05+koCptNVvSSrSqnL7xwU
Gs5yg/3asg8AvtehvT5MBjfb7dCOaGv68MoktQX5k/lRYJLmGO/CVBJYT+4b5kga
tOcdPiUMRE+f4zRENnXrzG7ngx+FMsPjYPg+Uv8/9mObl3g2NMsxFovWwVi87DUa
7plcva77WLKFQGbUNJ8hSZYhLbH7LRAxehZXC4bqsLA7iFbYa/yFaPD5jshXNdYO
d8dbZoyEXFaA2EELyhyTkLL2bngopGJ1Ad6PeJ6zhAa3Il2HLLNFRuHxqmTipxuN
9JXSlwh0ZbQX0s5EglA1qTAFseBHQEaeby390bE5UskxfCBMfHxNyoQ6RVBOtH3N
egGAqM+X1ObxT+AIZCFCN9xjDTTceuFJut3TKy10Zru+RgZ9xWyIzAiagSxw4eK+
3DBDlbbOp96Cs3zDxsaHHTUVfWsX6f/dNd4vlbg0b3w09Cux5fPd+5BMWfCPQJZx
qoE1/It2w1pcG7lTQZjwUy7TAttiJlwgxHmnHwqjeTjaAG8I42NDC+2mpIbmnbVO
txYZj7bAXPOfs10QUOxHhFdrsskVnuCYIH81fGG2CkWMr3oQ4kv+uhNIH75C0vSw
D0EB+L41fnRqwLVa5TgpeIe5c+eRVzb1YnaYv+tO8QPn8UNKJEoQ9L2pOiMsGbSb
f8Y3nuPhxRZZplP+p9Kv3k5F2GG+Q90U+YDMwEKFWBO6Pn1Kd9wO/bJ+JMd+2VNs
k1/tR4on2WwDYS28AfdYjfrOQabVOVj6A4YXbUV3kAsNOvLQvIVhke3uTCY6xUFl
Hte0kflCCHUXzEAKyMUYiQlATBSdBYQh+8paF3pPAsUdbdPdyEkKckVWHyNtUpGh
qQgSgYK1eBdwze+Fvl5FAdcJRJaS9Arm/G38EWd9BzW+KON2zpvdO4sBrIN4OeG6
Gqh8IJnfWBlN2MYJnP7P2eIYFRLKbrF8sbHcJvqGaoY9b1UXrrT9kOhFpwq1ekFj
bMQDpCR5jbYyT+kxHPNBWxN9IxEg4ggNqOX/JgLn/i00kRwQia7EAj8dIrcWhnxb
LNkBS1hEPB0Glbcb5WmnowEeiD/Ai36+tgra+v9UuvTUt0/UOjhfgD4Qm99oJ+EZ
HMhh6DpjwrmmbdOX0s6+9DR1RP2awSm9ocP5rbSjinQ0apVVIPt35kzUZIFD10z3
ZI8/r/rGwx7X2kf2/II0s4dzFqpRY2v5Kq2ZYCuV4LsHZ3Dj8YwYc6j4iDTLdDOr
YdXZDtHNwvPN9EsgrWZmhPv3Lk2Bw7wkDYT20cxVF7P57jTX4Sx7zya8TiMRBG7f
rbXnbm+y48cxPgPhKNGe9asZs93U9SYaqEOzjsQ5/S4NX0SKSEch4QfavEBEgZFo
OGdfX+agG8EAGNEZA8v/rJ6eCiYmbi3avZA0bVXQTofO4A9UvkduAyTfancRTcC7
2gmWkRt5E4jgDW8LsHs+Q0iVxdgaewr+iPAfZ9Pg6feMwHB7Jdb8TK7YT2GSekuV
MZCWsf1Wi7Xn3bKGswI+CzE2M7LZSFXMFb6lsp/lGnfDbs6twEAWgUErR2stGVm5
CTXVdGWD8rNHMP7xqx373s5EjhX/9G8Us87X5NjYVgoZ/Q/URu5vULo62l30ODfq
C8JWOxSocDG0tOiEkHB+kM8iZF0a6BDiWXRyFW4YnX6An1nI6V+pZyEMqR2FdIJj
Egukr4MNo5w/wr17mLUN58VeWDfKDtx0Y98wX/yTrgI0OXjMwC9mBZRl++v0FOn8
sQN8/hJZzOAWNfFvNGnrXKqLcIBKQ/2URPT1fZFZd+Kg9AQ6JsWj8Nb3uqgWHaXy
7pZVeN4nQcb9m8X2CGIvOW+NVHQi7Fw6YDjV4V1ji4PYYIw/xzHsyKNp937P3kwX
X6B2u6ixiLvqMcVR47mVg5Iu5d20HQm5XjnEdHJAaigm8QmPDK+Vej1nPrb6VNE8
XMBzr8vYXgYMCABLq8ic4DHS4WKyTn1EFF8/JVXvN0yZY/EhHcuPsL712P6JzAoa
oG2nypyEk6m1q3R+HN8BLrJTmiVoetNpM1+75pnVaP6HKOpPp7keNY9Z6bLGIAEC
Th5mYUtTTShZ8JAM+9r2SUmAXii+ZfrCS2zwDh+iWSuvalbjt7M5YyzI8GsXmCZQ
UckgYt2/fNa3XU+yHSvB4n13POox/WVwJ7lwoO8ClIZtg90uy4hrMO9afDTissXp
ZLUn7w2syh/bNSKD+BvBTE/VVjwbHA2JHXOHKp+R7L7ClyGuKHz7Q4ujEDg2n7WS
+gHVhXDQR/qzvjwx21nKuWvI/gboMVbau2wVgBUNONuYYg5a6w/NRKXCMItu4B4t
d9xFS9eOF7n9ff0llkoxvmAyPB088tlU3333lMdkZ6ENdJ/eOD/aVuYO4HMP0s6P
nhWItmCeK8BaQht0foIgcwwFzY/n3z76Ph44j6VhcpUTzIW+c4Zg3YpIRB+iNBqk
4uFnSv2kqhELOtCYSNwuSHxrdFCXS2qdhlZKjNSC+nQDndy6iscoj32K2rsEQOwf
qPsFH89lEaI224pN6DTP1t84L6+MGfthdKQ1eZOTZseYxs0JXW0lE/urPoNSaYZK
4X1KNG1ppFqSRAun0CpKNSXsQn1PP+xaNZXh5/fiwtl3iYGkI5r1cLl3baJHkrEU
/ckZYGBD/1gYkhv0VxeEFZAPQHMy/Yia++ff0jwPOYFGri214KANZMBGuXD2S3/t
+sjBTCChTbEerrYY28wm0KVASvLYfjQE3TisdnVw+kV9fL/bMXmenlio677UC2tk
286gGrPY+0FG5/Wg36fnr0JjRUoS1fYIcmDZ4RVeTRna0/wTYXfgkB8wrLNp8Ive
4OCmMoDfsTbtd0bHasuGbzEhGrmYnG4MfWVmRt9m/rd08ijZxbucvvxNPEsfCQB9
ViWdKTDlg16zOurVrdXqbo9dN5Oh02/YvkAMLlw+yvrzkoN3d5/x90sz423hn271
9N0AW2/ADbrrprS/zLr5RM7AoThftKIllEW0Pz9uP58ZAuIfUfcJw4jpOb4r8gii
rhPzsjUtGJCBEpeqJovPpuL25AvJsh44jbWIM2SlEB/uMUeYpNoy+4K7/UPGtWh0
WfYwfx6W8tYTTeW2ZTFpKwBz27+ChxuvDPaEDNOx9yExBEGHQuVFfqWuGYmn1ZWP
r2XFcqvtN0G0XDaNoYIul2oOTscQrzFlXBbWtJD/3hZC/9E2++Uy7fc3v8UVdTsm
4cjJLw+EsnikLMyU00N39W6G0NaBaLiw7aJq3GVF//0IKEhfXZS1gExdwcy1RfY/
b8OT+G52RuD9Z06waJ5cGtxOSWoV4QCq0tvAum5Vs1CewwPLsEHbHnyGZjiRbIk8
a5HCUAaWS7Qfd7erts1qeH1qfJEccsLynIXtjxzXUWnEIUKNHKBL6woCEejPpqqR
WPl4Ac6JcFfHN3e3v3NXd60/AveOWcevOUB8ast8zYL7HZw9KtzHFWQPRBAiKNNW
uRnfp3QeAFt1IRXhADHRFPgABbo9rz6Vy/bazqus5URUDCZRAJ0Zvll9uUOcahPQ
d02ifFEMlMt5Vd0n9+9zzhyYIA+WedFMMX8RVUGp9t0of4d20SiPR1dkyGXqN9fc
wKEThNZyS9DCjBzovZIhrYjmhW5vwG8VvATgZk4XFUl5YVMXZR5nMOfEokhE2ZbT
KvPA+8ha78nj/m7LhDa+3V9YkGiJXTrF6MTa6Cx40eycfN6b6ce+8lUOwCNozc06
p2PKXe8XxtsC6Tiz4ejheSBj5EIS4POcHzWJqQOb3idD2QXX4/5yksj6y1OZjjo/
MKxAheLHPWtDtcSZlJi740Gz5jDmw8BvfbVunnuo13oRLzmgyer+a0lhGugvIDlJ
S9tOG5TGMa88utQrryzs16LG7Wb9u+nXFljhQOEiBPLP8GZylyT3b1HS6UHRRObH
l1AIGngSCjLKtn6qeAlXqCXjPnWgnJVHfWVA8jsffIUGWQXK23RhZcjIxNd8MHNk
uja9bNkfwBGeHje5/LuRLE065tHhCB8iSW4KFEXLbxJAf77LoljYYeevl/11Mybx
6VOBCGAmSIx3q39scGm7A+Xemp4oFYSbctNIWtMoGLLXySnfv6emqXNNTdnKs/G8
GZ2pt51X6kRkNwM5/yNYfmYybb5HIRTki3WU4ywqB7ZU66ru/eCgHR6ti8jZRokl
4hVYErNwnvtBuBw84pIxGKpOEPSKAYhpAGsY62w1OIykCrveKhHPS4gfwzo0h0BF
8zka4leq9j4kF9SPyjZm0uGAZNdeNX2Q+2Z+9GNH5PDvlar6b4ZnbxIB0LAO2VSc
+cbuznAenWQSg46Yw0b30VCWkFa7OwBcsRzy7ZW8TnLbCuj3U+TZIYlgnrVilbxB
1xlHjlOLm+cBBxqejP+PNBQO9bp/adSAc681jogU5ve/Gk7FWC/fiHEiAtk45ycw
Twinflm78vTXufjW6UlrDv6DxkG/1e0ewjYgvoaa0tCywozLEHaZOWWD5OPRP1va
c6oNz0JJ3FFeTSvlP0RBRWdmhvIwaTi/CWIHyMJAsynyS2H2oyiAHmCJndCIQy/H
xpMEwCVHUOxFotjxwFR5DdObsAxb4YYCuqv/VaIbIkW9czKzJUgsfBlg+kewTVDK
6gtm7L5IDKVReu7ObToVhTIu1cZ+6P/+yHCD8QF80mS/Hzq6aA9cXNQoUZ2E3Ll8
G01UdL0qtttmxHT9vd0ICcVA/ZO3CjIhAR3knFoVnq8+sHXlANhzlBDyJa8EJrjy
NNShAexAvZAhGC0z44WED3tCmzrnjLVLD7qvrBjLM48I4OVqzMaUgCFx9JdxwH7q
mJGpI2bj95XQeZMX6V7lZHG7sr/fDEWiUDz8AR5xcWoAcexd/v/M3kFx40LeiFWM
7fDnMKw8M546t2K2uS2EgGnDHOm5NVG1DdYiosXkgkpflkL9P03XExDY4k1Lp6Au
+3gGDb/F25IeQ7gAaKriIBigZTC4GX2IurhmDbK3+10CJKmTa4Hg5UBMPk/IS3dE
pclIguodLHGw0EhUZEIYs8lMIFUw2PLGU11Ytwk+8oD5rULOSxlh8DNxzqHXg/2n
XNT6iaSMdM+qKYDK83H+wVY2eJm86BWcPAg0axTxIh+Rx8OpNo2tJZdFWXMJui2q
rfKiQtSvIxnOH4t9KxEvOAPPngcJOIi0B4POAu8cDP5FjRmOxqJ1coNLnjRsZL49
mYkU4eztyIEZnDdXoFOfRNnvg3zURpzKzHb9lQw/y2pP2rzBSt0kePRNHtSY2HVF
rq+bNcnaBFMO+jGA5YVybJAGzR5NZqFzIeSUSybrpoiLc/KYRNBkrxE7JAe8QHir
tvTBmDpuqftbZvU+5+jJlgBi1vNuQKYC+wuRs7ubUUSAd11RlSxZvpoLAC+hnyhe
Y7tA29bQ7l43XTh8pDkx84aRClQ8EobrU0QC9SLkpP05hwJ6J2Vvfc6lQifrxDSF
AsWUhoBD7yNKENISIdtYFdZ5TskDPXAjhNJVPOwpg9Zb8ti7cdO6AwO1BUGOQQwS
XOCO0uxuLcPWrZRQ9YdG4PKhCqI2sejg9jvtW1ZRrdYUovGqTIvN6+nRZj7Zq5wB
Vq0+WSV9BJEGK0E8dNWquy9Sqkx4K5IiRAri/BK9v+AMzd6wWmRJzTKaMsbmIM/n
6Xy3EXU8Gx+SLVbouS0RYvxf9SjXZwn1OWoEfEZ3V83lr68e4narBhGRtKnXAc5H
tATX7q7VqX5H1B+SM5OWl9JUQTcoEgYL6ngPz9x2IW2hwZAvm2kEhl1phn1Cm1hA
87HDslrtfk7gTSvSClp14wVtrhZP4Y710d+NEnm/DSQsZ2qq7xXqYpB67BsPLqix
4CCrRnWEJU4OmwvHSES2zyd+P+n/h/7IdvHa0Uyhjwm60+ba6JkjhL3+P+qLrxC+
CorOSmm1kIKY3VfzByCmnzD/oc/ZNGylrBRtuVGsvGrmLmZAq4EUnDOVnMPjqCfj
KAItm/S9wQOwppjsN64ePM6HVEd6c0+H9ERmp69xS0nLc3kmVXmsjekZWLF6c1Zz
YjfnHPUmL/cWFpgGSMD81eFvxtDg6EU/d0/FT+4LcdNmeFqXlsQNVltuuDZ7WIZn
kJ3M/VZqaI4GJmJKnqmhyTqbluIvqBlmtexfIMbuKwiVg8JySJL3T2ZTmDsCWYgZ
Bs4vpCl/m+tWx48bQNDxnG///yn+t4phihr9hFEKTsvPAcq2gIfcj1IVMlM+4oo0
IR1e8z1pvrV6f9Bp34s6qDV4/Kija2GRXyNGo3IeHcPJEhgDSyUop8j90FP6D29U
Gt/LnSPfJNWBlmJ8GsNBn/dWDAVCui/IevytBGhHism9rED4E7Rah+XAORXJn0xk
H8EWjMjk6CzV47Q25d3Bw02WW3b3n0620uRYi0khC3e7R0VunW1TaB7Fvs/Xqw1C
+8Cw1QJUahIITbWMW3Pi7z1NKrZzl2mCQHbsvI/ezvtE2Uo+WzxnWIgcxt8sXIoB
LQ3QRCTH/yjHjPQMBAVV6Wj+leAgkrUXKmioZWa4+ZZIN4xGVhS80v9FzGr3+gaG
3remeEAzLZpEB/S5uj4/s2qSatOWY5IVXAM+fEmmmswFUGvt1gWSX1S4dcLDWZt8
HOgs7mwC7VgiRaOEESVHpMOUwPbSLW3bu2xpURJmP7xjaIqOwVwA1kzygBJ2LhVf
AOXf5HO/3ACFv//4y4Sj5W4ocvu5msFfHWIYCoH00jqHApa69CerHxo+F7EjBnCo
HMKyFxHPavN558MjyD2/WCEf0NxMQ+3MWiT5S4arq0PuM1VACH4/CkQRGUEa7Mxd
3We9UbS4ysrKF9UvV1gVDkw8Z8hveJsykA7f6f8o17Uwe00OiNxTrlOZ4hV3oStg
MD6qkwBEJYvWVQd0764Ow9pVqv7Yw3uXxShg2aJqPu2kxt6zPYpNr7Kiy288irRD
sa7Ph95JVTgA5N8z905jv7kkRW3QiqVHHILMExm13mgXRke+hUQMk10cqlxVOGEq
zp8I2WmBqSBgVJILY56wuJoZPxwN319qRHRTjl2TP2tM4wr1OmwosTz7qGjVe5/8
Qh7RNV7RrF0bsUYZQOHZfBjrnOkQDRa+ux7FNW9noTkRw5zNMGFuGP6lbGJdmg98
gxUbVnu3n1kbD/B2EQy6ti/Q4gKqcFHug343Y9Xt9UIgOM8EJdmldBwHL7zIVCMq
gr8q38hLLqUIkckHb/Z9Zo3tDR2Cy4FhZuLWyAiVnqK+Xo4i7luDeIqz5gcmO/4m
DO8CW6R/n0Lfc3y7N1cTx9DRAR3DDkzZogYRF09nEqH96CDf5UopLAdSNdVqlq7b
NT7JzKLDZEXoU/iHb95Vehd69A96uXYf+z5LP26+1uQD9P2nkujcaTToHi/wySTU
VafeG4EyXl/sUJkJYrR6WzSM79R3Hi10buVvNoB0+1IK8jUOISBowIH0fDDWlDBz
gcMJJxK+F1X+wIJAuQlYqQ/ydgrC0EUuffEBzqu+7RgEjetfUwTtx8WvrcPvSd4U
ODM6nyoW5gCg6cIjxrR98JTMqDhsDY1cjmWd0V5tUi9Y/+PsjSZjkXKE45wH8xgI
H59UaWbysmP0PmrYL07C72oxmw/dfuiu4gwUpMDZils0zt2ZIxBgJX2w4Xd/jxsL
f/D4uISCBZmFIzmLZizxJOnGs6dPCAHYduJwW0Hf4bcvK3IOJOoIbg1jdfEiMWlT
VLXlyAPDZmU+oMm6ZMSNtJ4DgqYrr4ZbLJ3QaQV2VJo0YDOkI54JdvvofU7G2DnY
yWRd+U/i2LyX0u6KPceCT/PS162aVQzk85mnmYNwVru27bSj96FQMwpveXTpH7Kr
gP6js1QGx6OmpiglJhki5Z/TnRq4cYm3mMuFK3caT8IYRn8cvtEL39zoVddm2XRM
nDPiopPnGFQ1i3958zgS1Go1qfQwZYWozVJvW1oPifswsjBqv7kk9P+Xbna571dr
jqp+6OJxn4TPPaK2cuvw/rH1dzH+wTnwrb3eAHquaYseTvGK+we8mlie6jPo23OK
Dyf+0/KRrHKh0bdSAAbTQvbNkCZUGF+7aNA19IT11DVkgtay1ISu/cTmhDvcNE7a
mXRj12PRQ9VsfVIFNw8V3EtcikJahirL3ypxO3v1buub1/64ecYIMR+2KnE00iol
rO8S1VDBlhqjSrOM2kt7IfWvz9oIzuwXIqU13Rvzk64ukHQDiNOYcOdvjNAQpsML
bBW+IkUwa59Yn3/H/xDMCExlR3ntj9lZq8Dp+loeBOotlazUDyZwTYFTEsub0lXH
fAgHTHRGKnUUX9zhtf8wX31SdAh0xnIx5g62Lxs6q8T3oXjSOm86PCgELu+34hyg
J9pS73J+zwkHupSOX4soQVeBnJW54Scfdq95jM59RM7M3EJfO4Jbm46AcDhMotHm
dpHFa2V9gpQ/QKv8O/U907xJ1qhN1TTi7CRF74ehPcvfTsnOnnMST3Ya/JKFi9z0
+c8xyScXQko0BPlANLKtuosGPZGOHtwSlyKbtRHEeIRnhMmkowkoyzyPsSy+hYcQ
5k27KcJryFmXZDKNLobZ5rMee9b3Hv3I6EF2lZgK4wY44HBtGa7DIOEUBKHRbx83
bpnGOdQvkQvrfBl4mI3M8fjriXRzbikQ8k3S5buZDlDycCkwQLTIFsP1f41dVl7B
bfdJiM/+OrUPafqFBFVOETU24hLzePrkG66K6+sX5WOTK28UH/HhVVZCWoHerhRW
VZpShH1I3hbSy6ySd6ucHxlVtm9vjSmGJEsIQQ4Slbg1eKUKZTd9seijjxEDOiyz
cuvhXsxG1SeuT5rhK/W77TjMzWyzaVI5SCk1t+QVDdO+HatRMDED3eYvyOOhK/if
bat5nAG3xEyR3UzXPYaS20MUAefuHYBZHffrOB2ng3F6s8bErH56pnJy5fIp/nLs
aEqiGoffeMxfrtIzqHKKZF5ckA0rtQk78n/pfVH7b8ijsD+WV4hBkSW9DAP4SS82
g2F9tv8ooiI4aDxhScevxQebRX/JJmACBRsRSKp5MwVuygTk9FXLPxHEF1PRs8pP
RehsS1g7t72BKKJwDNgSFLSlyulDIba1aVJAEyLGZN054Anqk1NpXzx+dBOWUlqg
tgfokCEI6XkeEujLvEW9hhnm63dPsEL/ahVSBbXunqWtlK+p5EEEO5eyrfC1XJrK
arFvpSb7yXQnGwOcdRaMQFeFzj8NK+BHgR8fC6osCdD9I9M8Vm7xfOUOyDrP1B8E
BIXLEpk2sDwBp90yjgZaU5Lx732lJMbIkY2fsiHWQ+iC4LB+mL0KTnazdUpL0k03
muVJVfcFlXhsa/7OczoK9n54rPjSLRvFe92LeprJ8Q+ilKYiJyU/ZuhSuxcU+f6b
vL1+mkbXbDxXfnr1cFGjDGf3ZwFNNJFBtbCJvYV/7r1uTpy6tIpXpxq2LnNYPnlF
T0o8+VQ991yGTxK9MfOZFcTqs8UvAFOL2WNNl09NY0fUt9Owapn+/1BZrmf/oumq
dkmwR9TFO3U4PwQIzKsvXMwtXRmIDlMb4ewrIk0UOxvqcFgYaccvikGqwIFuvkKO
HfaxTuyFM+B4rLZTPQclVfl+I7qQMuewHhpoEmdGnDXDXlqQtRIKwh9ggqYtn+vu
/x2bsaY5asITHAsZOvWfVuMrK8bYCpAemwamZHI6i1KkrB9593Fw2h6sJFReHXBN
QirOFpvVa6yE7iwxWdD4ze6f52GIVdmALcyEjWJ8eXNtZWQbtsV633ia1vqJ6DsU
gqNuIuIap57qhBTZwRI3/77JCpa5pVojcCFjq96QUk4YVnEqkl8MsbHy61T7VBei
kRtkFW+e+VHpHDxAHb4W7acnYCIA/xbsA2sdzHtIuPbHJAWp14uMth4nH4Tm+KLu
Nx0wK7lAnDsJAFc9o0Kfc8MjnG38yir7wnZ134YwvhqDB4Zp40TVKSYmwZ//vBB0
FC8EveLE8HhZ04LbiWTHA+/2cUiaD/e5CLRxBUs2S6OOJWcnhtJv3LSpyq4ZkB2V
aK8bwfxPhBdNGi1XVwUtB+o7gP2fFYkQI79+3AnRTG5MZ41BZb0js0wXHhHo1cOs
Gh4TscEm48aeWZaAehWl8OhqNGZt+xEKsAuLs/lOLITMKi0NYp0ladrCvJZV42nt
6Bi2JkhppzXM8cjPyucPEeH0NzDFO/LdQsDlyS1A0DnP1CZvL2eV3tbvJNZ5vilG
ChpmAKUMDvxaouOH/bGvC4vUAaztaRY1nK7BNSCHEyOxcgOC0m661hl7ZzTKEIWg
a+5BMXot6RQbSZCWyqRALG2CmsWwTrDLsDyp1Qq1m5OcsBMGpgEvjuXVSrj+PmU9
vJeUUThuDeJUi6BRpamk02mpShY2zfjUH8Y/GZyjtZFadEgzWpA4c58GxiGNSY0J
KVnF8vNZwJJAKX2qxDZokvtdljma624mGWVBR4nJVUf3kEOXf+i5ykwkeCNXuMUF
azNUPDDH2mjK6i0XYvxJWJNBhqT6/o7sGk6nV0REXPHGAceAk7Ze/AaOBnikJpGA
QYJc20pLMVSzUlDzpHQlWe7qGxcIyBcf1cA+D/IWJKtgHO+9R/m0mB/ZESTk0CIs
U3LWpkge1GTfroyualvS8An3kySZv5JcOck1YrQq7FwocQik3tfzxNRRfVE+R50R
Ur+aiGS8dt2AoLgFsI8qglAVVJlzluJhsLEqFQntj8WyQ5AP2KHV7+D4e8x/drsI
D0IjbDNXz0hoPW22rXEHc9tXTxdJQM6eC2Xt3vcq35YRB9ofptHFwU3yDIxgmcHA
gVxZGLyZkdNi+VJebY6uQ8962whCg3JHaUj7RsIeWC0pF47Sp+ejmtXuU9Kf+gWk
PaQJxq5QnR14hRu7EY2N+Nq7HuZhOXHgj4o9w8l6HNp53wdkuW+wcz+dqlhp587r
7OemtV0XQ4T7UNggoSDNlGjVXvjC7xksdxtUIKQyob8LOLDGA5Ds2Roq2K8FmnYK
ORJYK/ypov/ALiNJqKUix1NJzfvJ3zexK5DDZ9lvXHTWMHQBd+NYCf+NKrw3YdzK
+riyNS1eU1U07FLXIqDJHsQIk/rAKBXGlZ2RnlIMf3o94fKj8U0/+uSmEo68HPMp
PE6CfPD3oSe8VIOZEm3NcC4/3VZP8+7O0JdIRhAzppF4ZpnEThINL5MYHTmD5pJO
l0Pny4noimHVj/M+sh/PxMkJm0WL1wcGitTWDAr+CEnstwvVCLafby6s3zEngy5m
fWnGLPuRfnHiILkD3VnghQrHDvsIiQ9exUNPanfIQBZB5mFmkO/12nWnbbFkfW+K
LZq0j/gTWPm3uxzHugcriUQ+cbqjb5pEKkQdlHUCoqTaQEj/JP1dpt7HQ/9iAHJK
nl4HmX9XKo8wq+ZQygFIxl6ZZN6zB/I6WYOu2X5F+rdThkpjURqtlubFqYm6Nq2F
drC51CWkEN3mppY0uJokyZLeXcVHEf3oUv4/iThDdIq09dSKk6D2CzdqK2PZZMLb
4AMPSz6ffn5TD6KoNKBkTmIYWjUrLCI2ZjKy3T+AoqLez+9iatla2dKeWih/9Mg2
ANLjLM8gl6BuvmWjnT9FYuNKdIbBf3eDyk8AdmyyBTG26g8XdkwKxiIm6FqxkPcA
QqOGpTRJVWfT7IuRdnSHxMRLdLARa4VnNcgVZPX8330TVrsD2X/9C4wK09VrBxJo
+fLiGHz5zhXgzf1XFNojjfnBFTLe+QaVsLY2SgGvwTeAI1qiG04eoWPdExBZWaC6
xSw2CiJ2bGdC8mfC++9yE2VLWcF59wTe3u1nIAiNa609EOH9dlkoMmDMDb4grh8u
nZFn0Slr9rYnMyxUnlXUT3SqfUpGHvPdaSoJz03Dxvtrs0AZtW2I3xI/JFRvRblM
Vi0TasxtLqvme8QQFr6D24+d8sJk57oZOY7gSAPyX9sxEgaTo0bpgVNyUklPkYno
9+Cam8MRvdxcYjhBLAcrVq48nye+SRAGD0eIZdt3RHuwhuuJJiOBvoElzPz50Bdt
pdHFPr66KBqkJQNMKce5voKYo1gjRR/yBsNUe8SiRHKqznMZKTFcZutcM/Vyxz5Z
nHvsqAgKRol/r3xhUwNypc6gtw8QF/sF45l2/ZrBXxhKd7DBotPvXlkos+jfHRGp
e5tsx7vzUti4cY8Nu6LeDtsS5J483U7GcCfxdtlS/Isx9rfReiftt/QH62IEcWh1
l4fUWjHeZOb+LLtrSvz8dta+KxdzXdG0BG6XVnfJzBJmMz6c3P0ry6Sx0X+p6TON
6n/0a+qYycNg4/YmbAFfETtlluWxA8vfRyafaldE+b6LDJG1m9MOUDlOypeC3MxM
U8JHhE7BuweqE8pxQO+h5nuskLwue27jI5iBXN7saeQxImC6cUG7Vv84j5LA+/L7
6D6A6TuNwMDC3rUf5yEdHprUJOrh7K/zey95sKz6c4lApRgIbnVfIXtPbT+dwwT3
XOWB94EepguYpTXXX3PbIdcgcro7WsPTYDRfR2HKJWvOz5d6sDwC8RhuwnTyZYaH
i2j72c/HeV1zqJzDgU2Ki/Y3bn3wZG+SnE1cEeuaQDrd+Mgiwj1OppLTqujz+KUm
kVxhLZFl/FTMM3QlkXZGqd4PfsSwEtDHhrviqkZF8aZ/b3VJzQSRtjxEdUL5eDpB
j5wRQQWnN80LA+eOIXrreLir9xXevteaiOx8ditbdIdOpJqXODmRC27c6ZGAeDFX
mIxnyNT4pTzzRe0JKe3yCp0b2mfyXfmxz6RvGyNuUJe6wJpU7QBvUjwuSsXWqz9E
JGQjfBASGB+vCIZ4KnzZc6ZNlv6lH0VsLlI4mnibNCmtwCjnk+9piVZk0J5aeED6
xqKAxxuty0TolAAh5OYqR5eUtml4Ni65VvRCmmsPB0gDM9XfNwU0PN0p+chRKbo+
vjatL1pAIaurDTTzMtrCD/a9EFi8bsEk4NG60aPicGnOYRe8jpB/zqzp62/DWrxW
+MKIkWb74nBoj7d5ial6AwuaawIvSoyNJaDy32ZNm5Wxl4jgfW60MfVsh3dkMic6
lgC40UlEVERF2Rj/Uiv037Zrei/zKRe0knDCcleTOwkBDVskJAwJtq47XmYXcECL
Lj0QhoGo3lRK9b6xJ04t26kL+FMQLHaEpb9L4vYOz+ZVJGhuaokX7VB2NMpIni6r
nB7MkG5qBXbjHUOFWGqcuZa5E6qXOuUgSnZD7bR7Rd/Ak/eyeRiw5hwtaUi4dnYn
37gEOyLW9bUxm3H6crb39Kbby+vKZemzirWLk6d+/1V+OtSgMShnmpw+MVKlxeOg
7An6ZnQITMOptE1Pw+uB8wSZ+DTzvWbBHEFZfuRDEv97EVTSSwCNzhTCtxPg2tTv
hrFzyMY4zKzKRAe5qEjSWzYKI/gFCYZXXF9nGyL11I+yBlEt655+1ME6AXpn06WV
LneTfBPU1AgxcB0wHyt2KTMGnipvLpTZa0IDGjmIpoROSX7XMeZIe7z0N//24UtE
yDLtdlG7vVrKXHHdmWhhNDqNZ46RbU9a3KGDY5CWpH0Ml0Ze5rMKene++lLjYSoi
3YyxRHVL3MMyUQVQOxUg/F/r0LBmx85Miex+DAxTpVPbuzCCAcieTC+gZqQYihrL
yWyW0a27cNWx9xGUsdBQy1HGX/YdYBLLvYN0VPZUxlGixyvAGRVTjCms3H9cLzMk
vwIKA8fDKFTw65xNh7a7jO3qThRmVqNe/AjaYFMoYiAEtcWs9ek86BtelP/CyE9r
rsbvgMktNvNmXQWXdetbcTXU+hm5FxLaeyMFYRvtsO59Zhb04MmNOVlCv8YknTG7
ocT7fppLeDWE8SsGLIJZkPvqwT613j6OSUylkyjmzpwYq/Hc8xy5Y5A3KydAqT9m
UO/iBd1owdd6wHzuCcayX8GwOyqdDmy3rbPDTHLHHP9HQtJXsZWZj+IMcVT/7lBH
n1b6MVr/vodOg9cMI1x4HnTA6BVXUyZy5kglnluLafFZXhJVX+xpaoM9C3/3HnaD
mcBKPPFUDKNDHk8A2X8Ir76j20yhJeVfObP7Q6GlWNEHWZEVTlSvsw4FfbGzOqUa
h5cyAjEjEpwzc0JsVIw3akmtuHvrECLDHdFabMtSxyVNqapRvfGpM9XrmFnpwe7t
0Um4Vri7uLKMdoBu8X8PkejDwvI0VEhXrVtYaLl/J/Lbq9l2lFRW8lb9Caq1DYja
U+1+F5mlbYxmR85ZZB2xPZoXvSTNVu9EFM5dTJTFLuHmuYgA2kUf0ro/oRugvCwm
tTTlT4b//C7wFm2f3a5iNoywgXDNbR1Eir2EkrDAjd5dvQlPbqTwPebcH8FRlIor
7Ice34mq3FCKkvUhsOeRGpzp8SqdIPsgHyF6RSnXb6G0yApJl/cjuU8QVDLn8afl
Ks4d5xlDcb2r/5OBe6kdbhRsb3fvs0fHz9B3CueiFVeX7+VC+by3ax4ZbAhzVpek
5pGfoDeM2a30ns9zLAyJIukScazjGTa8Q6hpuLHXP3iEyg4erXZQtedADGJZmFDi
0tBihz8VXHJKaASunNsEtyaNduwRxdbK4CbJCpdMVhjbDAHyatvA0QsV3p3YD4iY
3GlHXag+l/6DdjhdlQcaRvzPp9nZHPfFuirRhSq9Ep/jzhUdtyiwhQpkYN1m09gS
DeVRx2OQ7lRGZzLn7EHUqBbtFTJ9mZ+VeB/+4TNfL9ncLtCZLKsRccQdAHc/hTu6
ff6lPGLLmsLss1ga0+LSIvUENu0xrPQ/0n6m69tyv4DKxSbPIsb2fta1p5VKjOWG
+z9gpWQLSUScGAYTRVgVs5i9QUV5pGMsetlGZAK7wk/BqlEtdL9mNXx2R7MARuiO
AdnaoISeh04VAfF8dLlQFYk5274JCqc3yJgf3I/iut7Q5MvkqHBnKkABrHnpPlGX
ovtSGcQKKNS03NpyR/Otjsj+3INGgW3tVoLOH/kv5Mu/WTdxR8pf7TCP8WDF/xmo
Z1dd3B9J/jdBXQkxMdL1aVMLktJ2kVKS0zmTzrdBGSzqKIWpT/TobAJJ2fuMD3+1
4TrGfNCZZijbHdpYzUe1pdsCw+qEd8szjFn3B5NgEhpEBacokT3QGivZ4csgFPRh
vZ58EjlnalITvK6LpPH0hB+/JkJVzex7/eAZkeqvmtFi4COwKFrXO6VffYCud3wr
O/NWpUfTtMl/gSipoMIMprhcTQ8qfD3whU4tTybyo6YCua5TyQ2lZDD6Bwl5MNzw
ZzwnsYdoU7GF2rii0rgnu+tkWrCpBvLzTweYFXzuNvFK3tnhuh8E7V0fYNMF6SrM
Aakz40WEWBukwb2gRtJRCLdIeLc+z4BN707VRsfIdcc84DIjMxR8JVp99E+EazGV
IkMIwvPquzN18Zbu71lu0X0KjrFK1hhn441aQ9yHafC66nMzMbXKTHOT1tDdadAg
F4D2qIE6+4PwwiultPRvO9RipACsBj7BRKpcy16ZF53nZxlJ5FkbgwFjgflkgQcj
jg7+OajjOLl91VNB5CZfQ/VUn2ChtSkVf0MavQl3ilCo8GAbivMl2wwIfjK3fIZs
djxpTqCz9b2jkxdeBw65GfiCcAy/t4ThPgatFAjlY3lBL5s39hXfa5KAN9CWGYsI
ZwhYQMQTsM7U9DDs68XPGHwsU7Af+SwEbk2j6jC1ZN0Hpojo1ZIAL7lzO99UrpX5
zWQREwgUAB/c1D+uJihIM26ivyYzwjPFG1teEdYKwXIMTdJPs3MB1B6H0PyV0rTQ
IqpuOFnAD5LBibmbXk6tQQfjidZkgLU4sARPZscq1rGFYVcnfJWLRzZ1z2AtZavE
Oe/aEgniaPzh+CCuay9vjYRt3shNDmv/769ni8KDH9i4U5xD3qis5Df5C4ACRkew
/5xtPLoRIUO2lAfNLP7lJJFrp3Glnt/n40l4h8TfotkFEiQxWdsylI20NnpHQ7LX
3hAYNa1r8I70ghheJdR6zAmAlJlwUQbz0tUq/1DECheeaOecf5bRC4wjWHQcV4KT
cAEO5/eRdXGdE9VNK4hYTzTXCd4qecSsMp7J4yiYg1ABNcL1HZo/Sm3gezlBVtpA
o1qYsi+arnevlEGJNeG36G/pVSGjQsf3+WUK9YJc6uRzZWAZlm1151McsZkFU0/F
2aPHHjmInmuYgRKCVtY+5EepdsVk28PNrg9I0k0rue/+Q8S8Gn+CG+NddNXnriEb
Y+9u97igmceAfDza/EYq0WwbYl5xgtWMQbCcuFbrsLtzt4+jRr/nr8nWga1k01Dj
kRTqExIdEyG49AGmRuDv4E5Eitm7W7GvaZvHLtsHTtQHCGDRT0AJvEGxWt/q7x72
imz6bLq8+OF4/Kii8FkRBZ9xyOgScerN81Glk2xq0CgOXbv8qDY0rCH0/HFFwXmI
z+XHsk/gUk4JuakYY/jGZMa5ag19upu4IQoeckioi9w+lDLoIYJ+15/rI2tqt3Ea
pljBkYXGdyeO3pp3lrtwx8IbDsqKtZxo9BvIPJ4jIcdUDiGRheUjVxaIBbcyL7Gx
/EhDaWkQ6M5Q6UMG63dsvgl6l8zDiuveDeTCqW7+ydAGcPcicR3MK2WejivtucIJ
GVGKD0b5773dj/CqcJM1x1yrFK4eyO/a/EiiAsqOWEqBjZmMbhanJgSyKBLUNQP9
rAaoe/mTUpYL5ZxizZlCyse+3XAOk2MQH3UNdfMfCHSHF1/gExEsUCo7cmih/cy4
2zZdplOy5IDiv2TCSIJ/6f89j9Tt9CTbKUn59O6nL7w/5K61yX6LHUaNW4EKbgny
OoaMn+Z3FGcPhYlcZhEEBQsPMFLkW1pccDiz3azcamn/o0bI5FiNnWhReKGXFWjk
t9wDZtlfRn1owxiYmx7X3vT4C26Jkg98UErji1DwFXd+NsdJT11l2oRvP0e+UdPK
5ic3mfsbjduebb2jPNvtlOs88LNzXxHIzirBLwrXd+KnyNcxEM5F4GWc6aZF72jf
Sh+h/16lXuD+Y5o6n2pDQHNirUa7CuqFCLiNFZjE109XE6D/Ml7lotwRPWn+Oa1p
hZp+bCxNJqkp9mLlPVkQS5GSD7a35pAgj0V4hvEg+0KX1STFCE0HhnJKDqPFM++r
izwnw0ByKOL8VYfZOrZkV7lLZtp0FXFwcBBSsI4BFSqaRIdkfEElUezDu3+aeXaG
UPOk6I962G+4gkSJH4MueDuq9k3GCg/MqQAMD3KRhthKQgICEwWyVf7KXda9YR8o
TrjGINi7gpWt/bhbc3XIvaUv/7OWIql+wRxgbfzhZPPoJQBaAt7orEGtfadvHbVd
80BlJWB7c7VNccdBn85B6XXEpAwr9t6S2QiKOCTH1m2cG2ySuykikHSMUIizSVLR
7AEwEGRlXco6ddWHJLEgPYTsuQStic7QAPZW+zNl6DnfpgzKTbd/qQMjXYu921AT
+F29v6026nqmTi+vPFilcNhsh6D2OzD8c7olozRC6UuK+ZIh3BgNxYr7WAWBqLpF
EuZmlca9i/MpiKcNe0W41nKDOvZYdmjbndRx+gYyTJ5BLOIcU7QPDj+U52cy2j0L
igo+IuHZZz1VvooPEO0JZjIdfGH4A4t3azP+fQClIuC8N8igOiN5Ozx63jAMHNqp
r0YJZOjcVzQMHHo2iRNFcfTlQDPFMUrnhtah3kXbmjL3vSX8vFzKoBKTUK4mkou/
71jolfpN+RetM6aki+dIR1oUAuHtto5ZmJTt79KoEcOHfTwsaGgQvx8Qb0v1yZCL
VGVb6REXS1b4TusJcPmnlqwKfpKYmsO6akqRfz2ri03/5u4lzfw84Aji3R/zvfCe
lzbGBKF6IrudWmIy/50+UcMZn/FxfSRWJA7eSEQMKyTramx9E8wbZzTIyPA8FWE6
L1mIVRoaayTGOHlAaICMi48Yw0VTdWkovo0G20RzFk8ZKhNrcrCS+Nv+1zJ7GDO3
8a8aWZCteXXZVSQ7VF8qQV7YMFqu/k5UB0zm/lSK4iJ0T1x1D+tUOOQ8WpHgZQai
0X4IzHwyI4r3lujTwzuGZwH9u6TPPTEuSFG4bIuYOzlpGDLBx9m4/H4aLfNRZZxt
uikrle6V601kke7JAHoMEalRKOX8plc0w+z1KxE3IrfSxRQTJVMOP7cUppIPiINa
/JloIE47dw1YIgt5sq6dMH0IKdL3QmsYoNpJQajdHm2hWU6idbkjOD/GFOYXe89w
QS/EcwPH8TbzahvHaJ0qDaL0FgY1Nv3G0ZPPFSiWqgivM0T0p7eGmQeyjke5fMoN
8Sr3meN9sWPs/fyu10WZYjr8vJzc+Nmbyi7XL029dlUyUHNaO4+mIzFAG06irxjf
jsKXLQfIMqgM46F1o1O7Vluf+XNtzUiFtk8YVzWH5nz5Qlk6nGaItsTrAOCC94ns
TxhGEmBbK3A60kJHbG87osyl9WObnRIBKqrIfZ0S3Utr3xx+tg+xq4f9wE+1Pwmi
ywSzxgdgEjGQsJyYC0jiid5+rH9vT+yghG2u4xs2hDN8NrhXobdQX3iYRUwnfEK7
FBVjs8HYFSysSFyoH01SEC2uJfyO39ciDbpJHlVZVKGEtPueo4vPqFpc12ChYloi
15vGFIWr/TG8UNS8fNTaKAedRZQPR7kzSoVEKz9sN2udgSKDdzJU2HHri4xL8TDE
NqP+pCFWh6UZwxuqpp3fzFNYkF3//qcFYbAzyzsqwQJtBJl2q1ZKLH/w93XUfM2F
YT9sZN4pSC6/ahij522STCUhE+WDx4iL+zWfycJmXqTveJu4M4ELtjyg1Pm0PSS6
ELibw/swCTSUvLCIEr3BCSsFm3Lx6OfU3ARzsbxkiT/dpQar5hYUMfjwLKfg5ZC4
QfD/8jMtfXZffN7G4rr2cxkm6XpMm/76mGOkllq9V8j7+utGQPYP6VHmg9dqCGGL
do8y/E9iSoStAWvwJPbMaxDcrKviapuIKG/XhfJQav9Q99HJas/4rN/Gh++9pVIe
PHIucnqoK3JouFmBvsLq/JdGd18JFEwtGaUhhVUsCL7UJX9f/SfbvHkCXZWbA/8h
sZNjXYRiN97Ll6V21KrEpAyHdLb+FIhnErSeksJ2E0fDQVVbC6WD6o/g4gC6cTCw
ms81//wGES9GxW5GpDb5U4knhcl6Dbz74dyhG/spENMA+dzOnPm0Hybyl8Q5qYIl
lrfRazk4B18f3jnFF7lw6nev+GXM3np57+M6cp4yn42FsDbJ+elXLhFOMtEW3YBV
m9TnQxvuxQySNlNh64Qaz7ACMoFec7zq1onbG2OkhYuyEbCoOqO/hgEIl4Ll/9gp
JDDInyVs2hzyhaV8wfOEmssb3evd8d1S7BOFfoYhMF6EUytfj6YVT1AXh0cXWUbt
jBPj+GAUaYFcIeEn04xMfKNZZkxJqjP4FfBxVyN/WdnXdRfR2NoBUbXLzpMzUL4r
k2yDM843zsePhMdqmY7icNVwP45aGWGOJ+8CO9t8/JXnVmk31y2nCG9aw03gOHAV
KT5pXVv38ShDoYDLCvlxUWQ5ZY6dUvD5r79LZpIhZ40eTKqOjdCrX3sO7yv3tGNS
tuAQWMoZZLu2uEN9ezMvMHqYrYes/hlTDmr5gKE4O1f8WEgDylqV+K44LeAX6bCU
R6FwRbTfZlW3haHCCjOoxyDjraveeE8FQ3glZFG6x381KDptkda6FyhSPD/LvQJD
z/N2Ji5dKCAzXxPW7pRGsfsxLUg82WdpTu7x0abc1B+bsTa/gFuZsO/cdU+Se2d9
y0bL0ptv7YRVdghAfKDwh7XpHTTZAS7m0NZNaKVDuu/i7FCSMEBF32rhPSvoqijF
fDLiCX5zPOCZNTr6Clx0TmZ80NscuJr17T6pLQvrzkZPUHA2DGUF+ZX92vUYsi1/
V/ZOiU/FYQZ0+5nVXL4pMwfV/TblkaXbBPL8jIUw2+qV7MA7yJos/Eku7HeaB9+u
HjyK8Fm1GcLZKjsGBO3xpKcWBrRXV+FMSFU9k+ELrSGXNotuV5EVeUM/kB8Lv9uc
nTmNwzVBQmLdXJfElSPpT2suHYClC+13o/CFnLvLCyFTkcli3rA5V/LQc2duNAsh
/KloyA2r8LlqBvUI9wQdwM6n6ZdtFo0G2GprZUcB8DdPiUpB+jlnQN0GNh196Y+M
OpeYaugK0jaPOP9/p6Dbq8EH0gdwMavO506261D9ECBXE5vInGB2wMLxT4eRtljG
2CAXN59KqkUoIAXrfYsYg4Gc0V8E0QwzBZIHLbAaziV3J693dEWzcZ+zg6XzI5T9
Z2Me+sIpc+UGz0epC0ax+qetOcpTw+vFO10GkonmD3n3Oi9RVVSkf62Y5vGKDvbL
9YSW7Nzmj3nsstGUIjzu0/Ff8V7YgjOUShpartjPAxLuPe6OwgKQ6uWa5tmJHujj
lHQnJUXULTZ8Q/TSmFis7mRvNB2bnn/JRNzpHtooFqRK6FLDRpXTE4ODqOUdOPDH
5zrzQFEdBV3naECVaQtBsWYchqDHAzqOcQunLdIMg0qR/Km9x0iGRGWaj2sYy9DQ
QZe9hgCWuCbDSQ5R1HJJraWfd1itFZLPgsJWVTzKvwBvWMgDDlO6C7nNzzzMpuJD
hF/YCcG759uxDZ3WeFoc6X8zfNljRbzx1aBEHQaVCypAumFjlGbxXrNNuFo5QnBQ
PN16cdx1yy7butodBjILgL3I2LuSFM9hApSrC0FUsTiqpIQcfybvLCsE7OkP7Sxn
j8GQO4amFivw/Z7zoRO5a1xISf4rS3WBYNsBi4s/sujBVZuJzxJmp1nWyNNXYB6M
oN5bOz73yuqwuhiLykys77iUYNDNFnMuu0CQROUli9C0uv4zDU+cOAnplgf7JpL2
b0pIDZs7B5FXFzkazDua5n6U9n47v3UAIbPKDJTPXGlWDoGBA+xav+b1IOz4fAGM
OEOlf2ldvCM3e5kLMsh9kC+yvCAKARvD98p57zSjZR5Yz+gC9k6fDhEDMnhmEw1u
roITCGLPm+qKOaG0LGUXLk4Kdzs3eC6C5+GDe3G8/WMxQJwFzqd4YECwETDuRtLI
nSpeLDzB6r+q3BrbLTjN6xypw8qcpqoJ8d+gXE04Ec7dOhvIrb/62Ernh1fv03OJ
VV5zcOifLyTc16K+PgbAHElVyFkP/5JMXZ8DdY0iKGPO1xO2OkhvGEstrSb8N3xO
asYu1TxFe5G7/yB4qfyjkC/JI+sOMvinMC/e6o8anCttwryyg8IJmQXR9i1uWv6W
qEDn3HFp8v2kUTdhtzdyPVvwEj6Ws8kvQXb2N+jXoquvOEalJWyBlpUgwr4xXvVw
uo8q+Bo7KIqeGThbRNCJmPYceaapXdW0kCxxsaKvdHKneQCsP2eMPmIYcGydN9g8
5zR7C9yVx5Y9KpoVa5z47GZzOYbJlX3sBre2qHXYqAQMLkobjGuSlthdEF2J5Kcv
tAuv7USrXULsh/afH6wiYZ1ng3u4B16FJLgH52ruZdwhQCgGmnu4uwXIPbG418h/
dfRORAH7H/PcoM6RYpYV9lKQnG0zRsUdWFGS8F7JntCsYOtF+hEJW51xeacj9S6h
uO/iZ137o7teYvBjPSWVpY39wzBdq9/CFVL8knNg6wij8QFag6gy6F3BmGq5DSDT
DH2FpqJlk/NuJNEsQ0Wo3eeYyAp1oFQ+l6V4hNOWnp1lMkhku2iNf1dOL9iaYkeL
0jJPjBr/q33ERX8XCyb0yD547AMjp7zyeGvy29AbatG84Fe3nBO4MB97ump4k1w8
6ZyzUPxZ2qIzU33lfW7eDf2um1eEBGhSbeue5yhZJ2UMQ1uQmSO9DUTYUNtkfgw0
ANQluK2gCfv+ZnJZT4eKfJri5HprTFj4RQ/kWdATvFSNPEEr9Np/I0e0l7LSCmU7
xsMCXtRS3nYpL9epHSbWMlD9SvYe9VQ92ulznbt5z6D+xCbR3dH57QDAQI8DEtYR
c3yalcg1F1606M9FrgAG4thdall1LTG1dKU0Kh5awT60jqoaqQqqJ9XkImG78KAA
xlgbcgop1tN3YwrzzOPAMmohitfacnfLkTrZrwp9r7cZjTKzh/4z9wsd0B0yW4zD
Bymd2h2tg4WekG6VH8NupRTOXz4hXAlfGJV/YR7BZCdgopGHGX5LamIkQUHVID4R
HxpHdzSqr8S8rblqeTNoD/xc4oau6uU2P2iWBEfSZiM0+CG68EadfHCRg8KreUn3
Hs4NV32j+5K/D3z3lLnJ0+KfFACZ1M28jYL7mSHyVm4tbrHVVOgjM/UCb2SDmw7M
VoKRGsoNHanBeYdJLaveKpnl0TshO1dT8ixURgnW5o1rsRznDZ5BM1q5EzeLWUlo
UkWiMjEVAE5nOz79WG2rua7etYi5a5H4qwNd9ea0vbsQchlJ/xv8wUbcFAq5Masn
95HNobzISTUZyPdaWeVjW2VqKvQCcSmlJfOU2ab0AvKAQCfSsi8i7344JD3YWXug
00jYRpTVX2ThL/ZrFFg1IYaijGKprowNZNX13+682rSzwwrFtHfLdc95XJWWO8Bj
frVEk3s9vybI6m3jKhRc8CvO5Qugrev1YM8j59V7WfhJYGd2DJ8c3Wc9DpqQZkPA
L51ahNcGXqXCKCTyIPeL6sfsAXFx/Pv30YI80q9QXkhZ5PDrNZR+aZuayKa+84bk
3EauTAgv3VluM7xyBubUyY6OEsZJV9dsHld5DdO9myqfFQ+y84IGezUwNArWeQn+
XLvJs+RDGfn6/rmu6l4UmxinYu7Szo46sixkvPJVjZLnrCkOZQFbNFE3pdDZnGy5
sWFhCw9fiwdKkxTKIcjfOKvd/AnQgv4h9OPeUjE8DtIiXm3TodpAGBgd811j4p36
MoWTI3a9yM8FQDBpw0yIlV7j51yBaEmm1eAohSnr8bBeKafwiZIMx+aDYJOUZDBW
pPT4B+QQbXMGzmBpXvosVLanpVEhoehLpHonX3pjqnbn1vUevcIA1CdSSzc8oYah
UxAhHblDAb0O523FSI6Vllg8wlRnhEuSEt1a8dLasu8Lv6dyRvIdTMn+VBtIcdVJ
czzQVOIKsLN4A23P8quPv2iqMQYM4KNgrTFTHyKYMnSGx97n2+3fcFBnqiCV5bHL
6zLISZG2Z3b8EfkWyK0FrDS0/TkOFiXSG5zDHFRLaFcKCdajFZf6UZoleoMEqN9o
XHRBlMEqpgkFv2pxXhkqwPjwpDfXzXvZamw+d6TP4GaULQC39qhw/ztRYMGpj/LX
S0num4EqKQbjcbPUWvr1Wd2qEbsvCC/4FMAnF4jIiLMZYbNo65BnNWFOAD2SRKYw
TUrRBbxC+CBtxzogMWN/f1DN81pmoDhVrP1Em9rmjqy/hiqPcNei569mXD6d3M04
RASC2PvRV/d/xq5qULhsiJIGCufLqfMzIZPHrVjqTWKNrrS48HmRA+pI/7n4nNH7
LsW4AnOTPFmeE50PBuBKf+GDwHkqOfIMt+Ck/PCW43qZExBsc6qAh/NDRq0aXVqn
9O7AdnLBkQ8dtwbVigtdnFd/wtJf52K07N8SL74m0ByEefIIFmpiK2NZlGFEIRjA
PBFqJ7d3iLyWkCzdeyCveNuPS4AvHREnWrUuMgCNyn4i0A0rvhmYNxBm2WcvAU9D
TRad+REPrS8nj4Mn3l2ZBm31d423/Ax01lpTPgwdv7DaHrblenv0s6w4USKlQtrZ
fWq1dsfmH+kn40QnhS/GmjBnAE2Cv7CgGa0U9eUaUO3RTFvh2kZOTHYZoUTX9WoB
NnawrtoYyU0FWyI+Q1miG3noiBBhn5GH2zMO6f7Tc8JjfXnwgUG4XaDg/n1mgaE+
9tpewCsmYXjgiD3VRdjd5Ddo3uZC4tFqCm0pXje8Zc9turbbwgBrfom4AoTZ1Oh1
jKp4p4dHgXaKokN5LITi9r6uaeHnZalHMTf5fxfHa12VFsh9UIsNek6v9cwMo+Lo
pSJFQFE3nX+xduCNVfkj+j2NTg+tHwD1cvmaFPmczVR3ZBFBZnScywbbDKUIiuN9
1UXLrL59wH2N97SaNGel3G2OnmRFVVBvZIw8g18HGSTGTz0d2FuATVx5YmqX9cmI
sdzZZfFBjyHt0f6YXCpfhVBpjNWK0UU4bNn1uEbN3U4prJcuA51VXee/U+3WYV87
H20YhV7zt6fT8aEI2bvEIESY5QTNB5pfyljk3XCGjc2sLX7qddXekbJ/QMz0t1PQ
GCCNZy9z+ZaZTsuJMrOMNF0ugDYVf+xCZtcaKI/aAb478QqhxTu17h7JS3KVHSJU
pnwpvyyJ3uNu8bQ6WiREeUifSzAYlSI0/6L9RYXxDsqlG9JxKEz3YClEg4LCybkz
KJmZk4ROmK/h+OR9LNfRKTc1EIGnMhn6FdI6LsgTJP44aKJ/j9dY/qUYqTFH6Fwh
YsQLrvSDSYNMC+Tm1b8l5hv/p1G3jMLe2JBrPwZUAo1vYj4+vQhKxQ8W6OjwcweU
3mtaRpmddteDgUncTfWjNvlGAzPslDEv+m3o0xb2mcMoJAuSJmkD2veVc5zsZZz9
fIKHHkRI2f6lsidPK8P7BANd4pVoC+Pm3+AlL0mAtQGFKGHfXb2UF6WAi7WUtoM8
qlM8VHlX/jK+1u8AylxxSyFDZMHxAcuGeoAyIcMgbREOdX6rgcky7fClFYqXTjTy
qkqZz7yG8BaoSnUTx35qZ98hyfgM+/xniEdl415OtmfCU4pHj517TVCXtVlUZ81Q
UcoZPT1Kx9w3H0701/yhwENz/YBjUJKsWr4pvLOYmu47gpGf4PPrIzF3H9v6vVDP
Pb1yRgdgCf5Ag/xHvPPJ85x0nqPtEXKm5DkTkIrvA8ToX+3t2EXm0cd0RoJVbwi4
2D++wlzxMo4lON4y+oumoKPwbIBET7TmpcJhl3mLNHpjVWOdHYe8snJ3RxZiKC5U
hFQ4P2I+ivX1R3Hz/jSCeUtEwrKNA+r/v1//lqQoqving7f4OoFCCVJjyTMWq9dl
xntH5hgRT864laD8E2nP2/PtkCRsgq2/upfJ3EobuHLoPTS4mv6mCG2VoLk7Iw7J
esB9vT+q3movYL0CQoHMQ2Zr5A9iCEHOng/AO3jyKpVNBhmu0G41y+pmP6kQICiT
Kv68ev96xs05LWM5lxiV1A/m72xVTpkoqb7v9ynENd0wlQEnH8NS7zx0IDcZZSYj
hFyvn2JV1uPtUK+X4TkcwTpcRK3mkUSPoYUHgBhMtLSjfENYIqu7uEW2txfwZAdR
HddTEDmY1YbxDnKtlYjKimqzkhA9hQLQ1St7wrV52UMD1ZIBI5jFcYYhM/ygwBxE
6dqUqvqH/BgbikZg2VNjbnaB6GAdhu7TS5Vebinhcxj8CDcliUc9JhZf/W2D+0a9
/4GAAFgSLTb9zffpE03PQmZjZJ9fnVEZSX+er64AScHhPUnW7hgbDellNdwsBRuc
/DcTJIARUDkHvdu9+Bf4TaTmOHo+3qJmmPAHwpUBcFV4WtzYQWXrnk14yi6hTlgL
ZtkiAtbizBVUdEouM2Ta5T9fx8kBPc7Zf2LSLuLmme5DkZKDGBEPKHJ+BaiLDvV/
bRpgwbFU/ll7nnwhJij8gQpblk8Y12Aa+xhaCW2co9HNvtBB3mLoZDmYPjm0pJwq
Xm0NTroiJ1vzfmM3ph7kpy3FdNx6TenebfIybYuSsB/jHjfq7URZrfPpgZrAz49l
wSbS6eD/TXhzqv2DCfY41ieq6MQgfkfiLF8glvwt3nPkJ+GPHXJFhD40hNpzcvVj
jp4Ff3lHF30c22FBrhS8m/s5VHvVIA54G98ww1bfAauODdI4C4Nuc44tW3VrkaEo
YjXW5tkrWOcGqZJBOUh9ug77I+vh7SwKzdft/RhR/0iw/nuMvECwJBFNI9hjoptS
DZg1vCwy/QdrwUF0yo25tj+MqrGnTlW/B3o854+ai+XkLqsVonSCB1TTmSvxLeMx
tAKupF6mLrG2ugN2hjjLcuShqMZ8rTc+5z9e2Dyv2by/SxxM/zJxfFhO+eyd0igo
M1r+1xsVGyi1deUFJiNySy1T7QpKHdH6mEo+p0Hp7q36zWnH0WowH1SGM7Qn3ONj
Z+F2+fbE9But7V/+xDbJtSNH3JfircR6LOonXQd5MTbzu7hvdflEmwQdudNn6Z6c
uJOmTsGB300qhKrTNFTuiQYxwrSG5ZPoOMPdpTkIY9IrSSQvAZ4g4kDG1ay0g5lv
93DxmoAUCh8agOrNMdszACcRLcihlh6u3Si2sM86ylUP9bhk7MBn/NA5hhS18TBt
d9fZieCXal+wqloYLbC21nIFJSVep/iURRbbgWUOvRGiDRaqEC8XP3FWRSpwXFDA
fCaIWHCxpiKWcwpio6vrka1rpuOYNVjvv67mxkGOs5OQdfCFOmeRCnoUiW/0HAVg
to6neBC4NOWJ0JsqyYfWc2V/velW24/Kjwnkk3IS2rKXpQfDeoqoDqHJU/K//Dis
oEf5/bBpIPXEewc/vHhFAuN9QKnODdsF5JmemTCVU+QFAFIorT3qhrtSMqrPojIK
3ViGUnxtV6HYa8Mosy0SOKpKuu4Qf/7wQc41FR2tOQzb6VanaXc5w5MU7FPxJbFa
5e8DBv58irAkRhENpBe95U7oSeD4wTgMbJxF7lt4MUBgSfBwMKHXJNYT+BOTTqRI
lsPiIQ6kevGak28wnv1MEXncFcT2uoL97bkSayTl8LspWDXle7+a4fJOMDv+2wsu
w5/epp0kCMEk1jYSw0pb2sT6VlzHG2s/nw6vX9lErHQaZww4nijUyiuyNwcRFElt
IwnKT76P/utA7uUIdJpkUejPI5BdFi9YwlPiVPzjaggOB8n93VpBI+wzuFh7pzTX
l4XpDezeaGAQW5LHPgd4FFtcg7bnleh++5pY8McfJXlartfmklae3bZZBP3IMhmM
p6foQPIk2vYaQXvO6joly3nJyPpEEiAYAZZ15SRZigILUpD1OZhvHMaw67SPQABM
UkDAaMik13FNwIQcFQqMgz4o30mYIGP4hq4VpIsIYEknJk5EvwkeG6ELOKPdofji
ViJqjecy2awDe6cX5NWT2D0qNQqmp+QQTM4kQfaiHZkFNp6yT4wh1eJoHze+O0JA
xCdWO96Hp9+rfjmbHNp0wV3pcsv9Orur38M9d/6vB38y7jtRQJXfL0aL9UPToHQc
UhpbeBoD+nmOvgM8odZfR0l+Cb9n6RdhbbMse9z/OhxwHZ1rrW+0T8moMix8d57i
QplvO0+B34VoTKkrRabT2FuJR8COHsEjatWr0mXEu9R1kGeXz40Qu4db03rO55dY
KaGHm0RWNTyCPZfj42jKktAXpsJLdl7GO2jbw/gu/XFMRPxEvzur/GcRB4rv4stE
0J9FVecpgJXbS7jynH1Lwpf5sHm7gaNhlI3oRZipIBFLgTP3M5PjMr2vhkwtmmLF
SwC3vsITEaR9NBBeeXXRIJ9IYezCpi3tua+UNRhIrLvvwB3J6p2bXihjOZRygoad
4U+gtmil2kQM4pxJQEhcvY3mdJrSmEqz9JePkDbLiI5wlI5t5PX6yIspw5AJrzx7
keguJKMJV2IZ6YOkHu0CQHFXPn5lFa0XnUEY1uFiennxq4Nlx8gzPEClWmIYlkt9
Tdo2pSGvAfAD9FeXS48nlUPO2J2D5FlverrWnysw3h3VKrOpmC9RqKRYn5vE6DNO
RW2dfU/UYgcHGzUQQ5m/hmOlC112FPfCoXGvotBMzmxEjGvYS/z9XkBdnKmUp0Ew
N5Z71zVo2jWg3pG4WyOysfdLAazFi2RsrGuDLPkkwt3cVjDaRzofo/uiSoTrvpts
B4Q7LZ8yARNHYqbk0XwhnMHQgAKPZgbNys3lLuksGuF8btV4f+kyvCd5y/hj30/D
NKOzUXY5bPxmAd5c1mkQGxzcjS1zLZtznmV6hgU3W88QAy+OmKYAuDL/gWN6Xppd
J8zChhj9aWOu+LO2+Ziwe8OnJU/7ekx+YkXHTOMMdYCwqrYwXwDXHFylsaPpQ1K6
lp4dETXF3myxjVRndUqJKA9/zPmbUR1ICvWpJBSSlSeBx6IXXPvZtmLvM0sNEs5/
rDX4Bc3bFOUXZaqBmqJvghVYsMD577q4l8hJUQU6EyDZf6jbaj/vTM2VZW/LeV/F
uHtcIyiggwe/RAFwPc5ybN2d9qYY95ZeNPriEAYGYSoDueqs5yeZwKPn/kwpNyLN
qm56Rt3BsdWIRH61XlJZJSJ4jS3TiQ5V2ge+DBikd8+zS69uyfyY4w3NgLy6g/4m
MgTMghKqFHiiHQ4ayjYN1ALvPjdUVN1Bpdqf8j9ikiKxRr87ZTZBfFcgtY+igRM4
54pVO1OpnItiUycf9oMBy+4IS5M7KMzlq/RI/1OZnmTFBzc8aCs8mi/AE/3VzEl5
+im+dFVAT+yGbDYunUt4sBJE2I2fciBttPWCiWvSFuA3NMdFlVSih8O+2HS85XeU
/S91a55jpc//VBcKQlIhPlLIh1CvEo5KT+8nNB1m1Pq66xdlGIu5aEaRBOYpg9by
s7oIBMS7QxBFbACHJOnzqIH3OkrsHDrzjOFJqRkhf7AtsZiOdb+RQqLpwwYu1N3x
plp7dIJOfFZ9YetmcpDNwO59ZdtRTvLc7BGpL1d7uaEvlGZMitQf6mY/uQ+WIKeS
8xwevUo6YOCpNtYc0n4JKy73LcXBDbpRZUQEUvIvcpqzsNcZgvR6f7T92/3TEKaa
m7MArZ1xnqfGwcBSTH/KrmR8bSrju/yeQsUy9KgsTOyi6J51WpuSTmmv8iNBycZb
iThnHtUoeDbfGZKJQ5ngZ07wBekDp2UiXqGNS31WCr/SApEzPJv0H0rJ6nlCs0WG
Lez3XK2YtDTFYHjjpiMdANh9+C++AUHtKlzmBSmtp81rL3cz9D3WfK8RFkT6PCjz
DOLe73F4al+RbbP7rxDvhQZhFJBlfMGj4qp0tBgMi44i/YfvVWOxyUxdG4/qD4de
6b8XecMk3jbMLCmpBVILRMzhuNKpMq2YN7F0MqJHkVjDlvqrlBl9YzZXEGGu5ukW
bu3HHL4U8o0HdnxfnQEveb6ZEmu3FPd9+VKgnLvU5FjcFmFRitrdCYv0yEqpFpkb
w5AgnvK1UMmlllws0muBYFzft9m3We75bfEnNAT5fyilQ4BFZrCQxOJ9pgt8YWQr
YhvH/nXr106QLT8TIhibwOPx/O0GLXdt0yjUQSMfOM2qeBQMdckXTic7TExbCC5k
8TMeSm4Ig3jaNN7wdhSVck2qZnZw3IBlduuk/uXjTC6FJKXRCLgS5UX+RqKwrON2
s+L6MBhJYC14RDgqU8xkO/KNqI4BLnBq/OR5WwOYrmRzaVe/+Avg9vGPq7D4y1Vc
H1CIb+SIjMLisSoycPae8NShP9JRq/tSguvGHATrtChU3IqLsUvYfsEuKU8PrUW/
0lcXQyMkDKrSKVV3f2k+jomtPGSuvQkyfxts1mo1J9+mf9FF6BS+5lldl99cy1CG
Rsc/cGxIa7E1MfbH2hUASBUfgWXRefNGSnjh0HHXJzEB2/Z3gb07a5pbrEK7cWN6
A0nSXIFvhhSlsbatMrCQtJR9Lm23kvomLd6tY3Nspb4EsziAqrdyB2eBTWTFw1O4
eeuuQqlgrcJS9OCC1WghOl71Di/NGHX46OOaAyfSOyCzJAgdBeVhjeLU1tuufm9w
cBpIA6peoU5OlGZta/HHl838SCGpXNCzbyYpdUqnt/emO/EsznxE49NDHV70+weC
DK2v1DzmyMDJcsdRfhM2p0sPKDnhcKk1nixM34cwXTkodkX+yu+jtOR+MslL8hFn
j9NkEW70qL/z38MZBQZ3+0H5uaM7i2TksvLVBitVe9VM2+vIs2SKbt/0W44qzgB+
lAY2XzEAVuFHzbGNQiu5nO1bU/CKTyoYn/1YUO2Y+ycnymKsOfPirol3pGrBfESd
1MwxFvwc4iBloLIQfgE2Nu0G1ofEDeVS7pDbxGtRplvUn6AXwLVD9iFXYAFSAFhH
ph4YK23ZNrGCnPRXz2+zOwuS9jJr9H2aMji8VIpnSGl+a69Usrit7EC6kOJY3cdD
h5sjhIFvSFWlmZP7BMHpYTSR/cndb8Zz3RLV27STOKpXoc8u+HxekOZ2V3CNRJ+d
nEXJhfnurz0qGr2mScMHkNealgDxUgi8fu4RLqO64Jcr1iWu94WEGFe7tlaKh/FX
G6a91dru6PBXUBEmUarfvaaFUmyStDW8K66jqssMeYtmduy0elhHOSwPIhtpceSp
lUN1YyA+4ctH9QIvySKrh0PYbNZpBsCYwXrFMSb/lH9Z3dKnCZae7sKfPJLLf3mr
J0Tk7RsBMcYQ1PuEsu2GB96Eu5RKfrn+KMQXYcNIgF9By8NBqs9njt5EaupMsFYx
pod1gb9SYTkea4qT/Q2OcrMDO2m4qYKPJ7/XoGn/t/ZtUjCEqnkAgCb+AjodXw3n
cyn/hxV7sidt8cPEzBJ6BG51kYB+HRx6iCMrq/hOxTznihAhntE8w/PJ2qVcVUpY
cWKKiijI1RyKCoESCU7TvAokNWVzoNVHno1a4L+u9474XqZrLUxGlNkSX3lmcXKd
omBCo0vU8awU/Ks17C8svyFH9FL371WnfvbhYor5Aue0E+nTdXeAVvXSwJlz+vXK
TmChgZVbkw6LIV6MomMVoVXmIRfQt5hFIWy2MRM9QWXB9HXNK26vSrzRYyvLrwwC
+STAR9C0GAavDAiX32Vx7j/eEiLZepzvMsgTSrcQtlaLZhyLVyyvOWjOAubVpKQV
UW3cp3WJJWiW+xS6Gg0a5ydE+2DYYvaGWw0b8WOjXJJZq5cVW2X9ujYepj05LppH
4zSZqbr7J1tfdANhae5SpTAx/MqoHQuUU6Ius9fwRgeIkvRWgroiOhSnZGt4Rf37
873BgJoDJDdOJMUNDGDBB+XJJmYT4l1fo1G3sLrBYEeY+Vux2hmpNa5sIk4YiYUP
O1lzL4W3ca72EHCACNBk/BI+Mal9a2d0mM+jTckCW1IZEShvMx7tSv/qkRk5KOcv
4GgpWyTeGJn48dyuH5i3jpHqeqnsu/pYHCjsMT3MDPZeZN8VSukbD2poGAhDTPJQ
4f7WM2Xe3Rp7sO+ic25UNynYYTWUfRGyePdr1hG5fo5qe9bvfnCKN24NC+lFlNnU
dq1Th3sFnIP5XbMrBOpgH6iKG+hd0O2cr8lkoxhld378C+i2P9cbxmcWUkUdt8ZW
4mw7LIyDtZjYJVe286/isC5PhvOP23ro3k5HBBcwx33/qcY3pH41Tpeb2XEhNsdW
ybjAisQodWdh5HeiXD93W48N4M6krQJv4n4ZkM8YQ5tlu3Vmq4WZ2xDuclH3K/tn
WWYWdpTi16XsO+mKFj6i8cNJezkVXKxTrKG+P4odUXOVEde2PuYQ+vmm0lXnJ3sE
SwmMHx/Xo13vAvS/XrRe3VDaDAnhQefZ7Y4V3BNqOp1PNji8dHyA4Ks65PYlNNLW
orFcH6Qme0LpbZQu10HlE6ATT1SYrFBPgawDD7VzFsRtb8YHURNiF4wxiyI+lkk9
emh4hw59bBzwca5gBRjrtNScPOoHGY6YdDcA+U0lmGtUAuzGVLuQ6IK72gUy7IMu
+stczIJK5vTiyqO65BDYqOVEHAiryP7vMvblwCjuxphWSeDhaNbQX/FDe3XXMU/X
gz5aaFLjbCWgoeWX3vSaAMIxIagLlZRKfEnQPTaDe6TgnB2F81wb1bntURd70N3X
LqV8btxwvXkXjhzY/YU2JqpbGgl5FMfOYSsLeI6NsRX67Pcp+xdRmYIrNTYdEJHz
bGTG+7PVVTjXeCcWQsf2GkGWie0Xvj41LBKUk9Mhh22STXsS7f17zgGB8eBYAss9
f3svWAWBGu1jlD1VcrLa52kxZBonIpzjCs8neYGVXrgF3OksWqpQfywyyBYPRSdY
VBr0IwHyUtd/adR2j09ru85bmBNp3qT7qCgAq0NroIBcUIIjv173JlqlNfv1MX3Y
w4+ukB9iKhn7Bh1yQQV5Lv2Ow2OG9LsXSRavUBkpbp11U1MgCuGUbT9gBCeBJx88
HA9UQpl9dFZ5ky8qZ/tXn6xnWBzYGH7PRHdie72nIVkjT//2A8gdpKLB5hoMhPFG
8cupgTE+Z1QRFG0J8rhFyftkSlEm3RIEpVfOpcrGSkTPlXivDVpoSNM0gdlU2tfD
3+r0VdKfarigz3UB1W4F1MRvzvyzQ/XitjjnlPUeQZGTXuNeeNXt21IRypbMI0Kv
j0W0yg5b96wluQfLcT1MWWxOTtzAWtHhZYVnnW8Jv//Hnn6HJcksk/KKbZNRkWhq
ETfiLZJIWsqGT3UZQr6cytN/rLmRtnvVgA8JbIXRkrMlSd0Sq9tUC/UA2OGQ36fH
yKIBrhx6JhG6WzSm2ltUzjRr74mjoiKd69JWRlfKeuSNQ7/JzxGY9dI7vRAqkzdr
uTvZw6Q+rrqjiXeWazrhW1N5svQ4wfjbrZexw11sbvBTis/XI9isB1p2H6GDzBnF
jEuTmA5uFMdmfgaZ38rvgDGHxbZbQoQH7A/7zvlZyffecaUPoOXgIETZRJIY5VeL
TbI99wOoKEle+z750p699okNnLLsmbWaqXJwepz3RsT+y8TZmVx6PxdPl4fsKLGQ
81fvIqmHwgv8dX4c6nrwRWRV2n6HrNe/6hgqBIWUtcy/j179AVs0RfdPqZre17um
h9DBdxz4lAM70Kks0mhwVcmSnjU/A6/PgycYFEkuX0d7N7/0ABl5hBGlU4stgR9k
i97ZbMB7oiCPfO2Qb7U15FIjiVKlttoBk88SBzzmt8VSn2Tjnxh8o3OyelbkUIbr
5LHeGFvtUUXutQ9IDFM3Ztv4tquLMtDZNzdci2PMZHdGBlNxP47zG8cXdENBCJzI
SSIuyuBGb00Rxdmt1ieEWz03XoT+BBqJhdJeO9fLaNsCPRIeEvDTQz2MFpO9hka8
6djLU+ZINZnS4JBG2AR9VfzhsV9iMke0juOPflb07ScOW52NjC3WBTNmJ0V1XVUH
F92vH9V3kGNsLB4Nb81CbFtRBLJztc5KhyJjMHO7pHrBieiBBydwI80G1VKPpost
bf2d6GP2XbeuE+8oVGjRTB87fsSSDGahQKCwM9UrrUUmfFaqh7VRBIlYa6BEfiQu
LXqsRtSxzfWVKtHb4bVYb6uiygZAQUyODYrYIDPbvm0pYV2C4ePqaxjRCi/N3qVY
uc1W/G0LqthJRliauJOA/5PAHlfZ7m8vKXB2a0xm6Fbb2Vvdhw7j72ChX0UHYmAJ
J8f5Fk7Cnb8mbDgzCy3Z2pT74dtL9KVaEjk/SeaoyOHk+rJe0EEnxyNqTbuaEFzs
iba+ojXInWY39A4OXM8sl1uDLfj7wNInVpOyygbAWtvWIi/Fk2mv8jYa+v5Ldt3e
3Lq6xDx0rTKoww9go4QCys9iJztL6lPyInbLnQU7cahoEmmPL/4QtEkaMbHzLAT6
JweI/xXrVdeGComfZl60IA4euArOXG5MW+cvVjk+C1cpY41yNs0laDdFZ7aBaQzv
uspJWRaE1CXzn6Sc+HNePHtL1XwKjUtz2EmSUnk4oRKlSfzo+EYdwWeSUWHHrSMb
5Lwi2XrVDubiwLftP0r4pauz1RCwUninvDWakjEQJBh8asUgB8+b7/rx9RnU4x+Q
RoZPCqQq3bxAKw0S9uzYY318slTCQY8kcelKu0+hV4gGNaSDiUElBg/YWGbItnyW
ygEZeRIKnhM5QyP9svBUWUh+m+O/PjTpHdwCU2+T+NFKoQa9Nt/VrmpObmvsAkmW
Dm+fOrsci7V04QRAtiVxjGKUsYjZX8op2GdgpQZ4gdSos45Z2g9I3OClZR9svTog
M0T2ofeJUgpsTvGybUw6+3XANqv1HBM9fGabj6glfSiMae9Ca7Mp6Fo2zZrYsLxr
lVilVcwJMq8cPqVAq5PyWsf8WEjfs4P06ijjKaTcnofomcryvegPoChmQArsqHPj
PgMkMxG8txMycV0nanFT07Zw1KB8Z16gyf3O1IbWLh+9MmpSS1wVXnZ6CEJWkymX
y6e+n0QODcsj3d49iT6bqTXpm4skHPhhir/IN9xfgO875PhrgDAkF01nIVnYLw5E
NSQuCc2vkVgOvAWFFvx4wUldwEVI/2jRnU0oL0dibaX4frJdDUH+trvZxCSAELIx
gjheW7iMmxBH8EXdGmQaiGnigTJaagFsDgb6CMWrsHXP6+Qa98dAWyHRFCj6EGld
dPXvSFcE4eD4/ZPkS7i+DCBeyM/wz3JMOb5HpMqV1mypJ8EKwzE2Mi+2+sCVW3zB
dLl9dvfYMXfv0mKdtr4j1m9GDx3NBv5f9Gs5dM9draHK1CNhV2E7HW9P5az9eRRS
mTEatbgePmWPTE3/UAwLbhieUUNuo1b4PL/660Pcqy3tAmoS2f87TII99ueau5XB
Bb8mhQ6w2rW/S6QCnfeyq2LopJ9oQ0NValcQ6QdRqfcBrLPAexyhLn0J3IIHEdNI
9L+hiZXWMesomdA1yupSAJolGrRxr9Bc6bss+O83QjlltcualugX+EWN18exn5UI
nlLOSloBnvY6r6MfVx+Ry0IEUQIUDTARnmlxYQVWEBVQXH/g6iQNQ7OhomI0UjAj
Y3yO9jywwdndIUZwhpXWX1ZNyJKFTIL3SRt+Y+byuc35TNg2SEqa03Dn4fj0i4p9
BdbIV/01H0JxKwu+Z7aMQkw7Fp3dyZjXVozyPya42H9LosYfGlZ5jEb8OQ5qDHeo
Fc+vAo8NSxExg8+wYNQhyejw5MQVkvCGqwgt0MMVjooakZhnQuRpBXkw1QahAOpZ
Nu9LiTCkz1wwBaZQTwVV6RViSdVtP9mBGwBAdnsCb8y45KVdrVosjuM4Zfn1kFxK
33eUBqFPE/jAbKrYB16ABMXZaL4OaKMnb6FzEBY4kr/seAN+ERzYU0y6I4pGKyO2
m5UUulI8kxDygdCi8ioPozAhjUtxz3IAxpBX6L2d3Sz1TGIZkPLuThqeGP8t/APx
QwC2whQWADzduJIzzM8yFLb/dqYaradB/wifmAuvzLxx4TKNQc3Vcc2EYzFbfkjB
SFwW0oc9pcR+n16ezpD3RDLNl3ZUYDzwBOAsWpvs9Ui5PIofzermYh1pVZfihbEp
9mmBcQL7ehC5e8tgD/7STKHOEaJtP4afV47ssWPfvy7k+gLlDA0K+xrNkIyZVslZ
xpUW6CgYyQ/AdtC0GqVS6TDNKbq//Hxlk1LkmScB5VweEJBZ9Z6JAate9JcIQN5v
+DgZxfRfGOQbyHLLekmg5VTMeFNLrS1BEVNhb9Z4xVClqWkBQP0cInn6X8mW3VXd
XlJcLOPLIprjdXJ6wIAXv5Z/CqDm4dZFiEXjpHqs8s6TKEoQjbkzPyVSauSsUjqE
z+VEY01/o41Z6EAgwUm/TeOdz/T75660TA8h4tkjy74mZmkiwvLr0+R9fqsBtrnb
fCEnz9t/PCBu227bjqMqOY0dOGgz3THnWiKR1Y0qG/7+tKx14h9gsbB6ZHyJevRh
tZ6uNQsZ4J1LTcXxn/yvTTdHHOGVZf+cgpjrDD3J2iEm/HHoobRrjmAQtj6/4dm1
RCUruqqlrtcO8ApkCaJpH4EWPifsTU7Dy1QPjt1LSDZt5sPGRNBvjoNjAUoXTNVr
QG1wWNj2Yg8V8xKeXJ4Ghy0FTSh4W9vJXbAIdpjUkn0akGAiE1TIH4nDzoqg4XAa
m2NYtyAuUv0E/UufRvydK2FSo/U0+fAU5/HNooN2t7XXXYM2sBN7V+fQSyqzPfhr
HqOv66oj0HKQId/5oJIIfs09z51AHsFXf4c1Jva8vaXT3W2Yzr6zZuovSzIc1GTg
QmSvGQsbmgVviL2oJMjwxLPHPTY6Ykj+CxpfGaezA5tmSUsozMykwAJ5YrpNUPXc
Ojuk7+NXqDPbGYmZWEtedrZJna+GkDJuu5zh8YfplXUQw8B76dBHdpAv6DO78P3a
3JPOWzUnSMUWwtOuDZmwft59P0BmjdTWFt6HtTAAtJlLs0lwweJd8aFytol15yIX
VXMG9vnQQiISCui3KsPk1e/JqS2rPfY8zm12T93NnsrneZkyduXsKx2OKnsoWdNa
D/z/RH0DDcCK3AGqYP0MwtswvYfqnDgUz1lWyP6NVepweFQzjtyygK67PRLPJV3s
9aWaL3fdpcXpOfNmjep2czCjzGhegcxQVui6go4V43b+C6GVHRKoWQaxJ73Zp5MX
O/9W0Y5SWgDBRuDMDA6IkLpGImPEul3rZnNT0FJXLQwg7mb7066qKGUDcOsBS4Ch
CYnR7/atT+9IAEaIq54e27jgjoWvjb3xT2XOINuIH7a5OirvxWH7boIQqZw5NIR+
cZ7nqpp0L/sKut+Vi5rp+kr/Boi6DQyyS1vg1zF6rrYXxOd8xPkJaJntPLkqmzZE
nt9UgGWp1iSuoKNt+lo9XCCrNyyvuDGm0MAInuj5DZHusb0pKn6EYBEtZzdTZRZn
rHgMdg4QHvVVGjFbg/LlUYWxo4dHKM4GSdaBrq+/DkkbFYEob15tYPenVaEYMi+e
gVGytF5YsuzuO49Vu9/7VJM/pkgnNAoTxkJ79zg/RaSJcphNMET3mEfkF0jIyszC
rcTmgQL5k0orFRqihHzx2rpKHzeS8Yn4tTs0Ej6k/Y3jbXOvur+4U8nyhXc31Fyf
2uM0pJE0nS5h5wojNnaN3oLeWxN7WVQJ4R6nAVFnh6qpOSqXEwf6OMjyNQQFNVWg
N3mYRslA1XtzDt4ULLOeQI8i+pJb0yjbFaMB6y5MpvNpmIdFrx2ffKZSa1mkZtRk
MqhRKEaeSyiMAhPg0K195DfJrEUkS5UR9P0JVzmzIYJXSeJL2M0ErF55ncLtguNP
v8IkveeprU3Z9DCAU/GBqDmgxxBScxutkJ1Z4KW4qTUJ9yCLMudVBZ2W4KeVw9w4
NdXkpyasMXgHxRT3UuNCk2/OiZYvUpNtdMYhwuCoRrngHJIaJYLwp+IjDfVdlbip
9JKuArGiOcsXfl85G+SxN2Ls421GFDzJ+239Ldbr6ukZT6Kwn26k7K0uFBdOsf11
UnLvf4kj34Q9niGgevlVU8ZMFDe8+YHCKyRkhD7UDnxMW2cVHofLN6rYo27KRpkf
ycrsPFEt60uMi4Jtx0fSdh3qCmTaPsbJj+eeQVqijP/wQAVtJ0YemDpIjcGAbRww
CJ9Bxp6YE5mlsYzv7Sj4lS8WkaGQAKl2Duqsw4oeDEGzTCN4gbHRKPqalJikud0q
WWDaNHRMzBARxixndds41gKTGuyvhjiY9Rx3SFAU4+cFizkkKvJ4E3uFXIHWZ24G
mc6//IkwvCSLZlvDxcu9q9Sh9di2uetQvX6xMtUlRVlFeANA9FZbm5mtf4ohX+b2
/shbyEddF5U1aE6e0xJf5mTckz/h9zC3tuNA+boOJ24aYVTAvZckLTvWitDrR3Hx
uSDVo00BTCzB5gxMrklnKCgwlwhkAU9pu3Mwe/9QxRGWFbDLX08vWmSAuxLWfYOd
go6TpWIul7LWtpftVMCPAh/3NUDiKSINldyGIn7MNq8UPC0QoYXa11+DbTOvEmWd
mOv1kXmLSNVRGYfTHO56mkRnAazogSK37ciF2PU36+9AyryZVEtes5wZjzsYBjMd
OC9IE3G0bEJq2N68roFOrK+Ao+plSCT8ZUf2Ys63ATR/qBqbyfEY/BqPCFqHMVNk
R9wmXYMnNrrxYtkqNS4mgWt2l4lJxd8s4jMilLgfiuAnb+gWmp/9CoEH99KTPg/o
q/tYEo4zPLGOm9oAppiGx4TAzoby7MtLVbxIgJj3dK6WIqaCwfb1rfbvpd9oYWea
oUteHvv11tT7rAEWW0IO1z48WWceTDv+AejwJWqm89UJFqRVMchmNRQFU8aCQEhk
yZ5ZAzx8jvX/tKs+TyYFsSYpZ3ItS7wjpRMarCsVoPW7fRBs8M1uKJf1IKPkkOal
ZgUOrJvzM+IkaZcXfXOQMpLMFb6Rss6UB+bICFyNEHjf9nyKsfwogIeZojxvbSVv
OBq/ioN+OMYtgvaCw5Sf96WpA8Cy4MjQ4webdGC2b27tMmccb1wqiiqp/vwM0HJ4
pYWoRRvFq3RsZEvvqBYSnhVoBt0hHUUpeg33tGM4zjkaKCBwXC+Q/SFRz0jUxpgA
zT4DUeyI2s+6UkyeUTUC4UUDJi6+ezW5vxMmlQG4W191Xagu6zUaI9eT95LQuNcu
j/PM4x8qCwaK9LG/rC7yDwsybV5O2y1Eez3GnW8hYxG2qSUvoEEnWvtPTmIOZP0X
3SSZHSpo9Z+cQ6mR6B7KsTgszfw+j5qhRhiVBA4DDZcyM4r1CGvDyAHJaEM67BHs
LSkVI9ZFZoTQhD4/qQuPm0u9TzEvcP04NFhN/Fy9+qAcHXmrizrjGSajCELMXnhT
KZvJ470sA5McVwt6E5KiwNRPPjTjJWhArT6x7fzWc7/Be+p0PpFcnyEeoi6QuSOD
BguBp2Sc1OhptcYbcyexe65v4Yrae6pNUFv68f9A0wWVlDAJRKaoduoYwdYqu4ZU
Qbd7ppADuDczua/TDv6wTG0NPkcvGpEfy1OMkDcegEF22L8nd0P0GAq9Gntabt41
pIiqgzqx3SaIdtmRXgbo7ZlPr5O+GkDiVtqMhRh9V/Dyv/YTg+gmxjasXAXfhxHz
P09vdhOSnvzZXnardlD3odHqU6+1Qk8GglFB/4KBMmnpvxW8Jf1dKIgfUfyb0EoC
8okaLlYe69nf8DZKs9Nv0BllFs69U1RkE6/VFWs4lhupUZRutZrcaKVajy3JPrD7
jagzXTO08Rn8d83jDOa3dH7/i0s2nNxtha1XFLh8y399uEid5K1Cy4bkGyjZ8jLd
Ml6xw4qVepAJClkoBDoWsrWZ4ETr2Gko4eZS0f6MrYBxbepQi0Jsj030NQot/wg2
C0ye6PjoHKd1xRMmYcdoXrQEkXqPIdo3xHIPXOgEuaeWmO38s2eLl4kIQzJ78W1F
vlaqF6MywUR679PZhLkM2tqdamzWdzNKX8groKKgbBHE1vWQTh1rYS7i6bEkORXZ
77rBY97tzcchRPsTgCsXMstvNK/ZitZWBvYD9RNxe5pdtOLiD4l/wi+92ZXGg33k
rhOjs+6PrUCSPdE0PAOkWZY0umXyOoaqhLCjV8tFMao91ITVkp5MeWVuVI3mq1jf
dvdV3lUBl+xDXpXkRYOSA4yUKDxJiWpSsjtIY72RwbHXbWADgXQtanohaf+Pof14
ai7uyvhXcWWVTmtpQ+3YOfk86Do7bD82bJ7yQAX2S9q2KqSGkIMs9vo8RB0he5yM
REniY/g2q3ujbw2oIzwssu97/+Za98hWgXT9n8H11OVBzE7uKvxzDRFXtiQY7qbv
GRjwkrsXrUsLjUXUxLt9ta6darnQqWgnXtUQdY6p9Yv4oqwkbIKVbQnBgFOrKoS6
eYJAjgXUyXNiZEjKrbMko089IezTmeE0NmoxLin/PctjSGxd1ar9HkYPxFbF4llX
6bUThy7n8nhESPqeVgdnqk1YmhDqSWjt+KIsVJ4teLFgUonFljRMM1TvJNUk7MKF
3hhJKkGtAFfxI/BdEs/C6DCFbZ4+S44rtfOlApuml0ocvM/rr8pS9QaqQxcw2E5K
6BQVLxThtiU2O0xxXoUqv1L/Z1VzBWdKvGlzIoZP6BlGRHtbBxNw97CRkPyLRQBU
zVkqtvPqnS5mADIe20BSCbFd/FhdZv7WzwYw8ngoTm8Pz1SHhg+/09q+OQVjWkHx
Wh7BS4u0+KsUppJBvmrxXEjO+K4NHFqJU3LaGkb8lFcXxHxttpNFDsdKcmiZ8ktp
RuhQ87kwaawkdOFIuURA4oeyx04Gooy+qB1PQ1IDaLqiwn9r9kwUwNJ9bPJoufyC
7b3koGCHMQZHBldmUVPP2K+VMOyMOtAXA4QuIKBUdo4bY06KQond/9NhvszNgOys
D/TyXaSpDafw0giK1p+l4xE5wRU9vsk1pX0mwkQCwxvcnASECWovTikaZftmIJeB
3Ujtl2gqQtDt5Q7KUjxpCsoLH8JaWWkAfPny9qmV2+N5IIeHHEdWDSNnUxSVjQQb
lXqRwEWseC3h8P1PLHZLkaVcdh9ikbpecowmJ7g0Oi+IjWlgmBWpxerqosWlhdtS
i9/yF5OY8FfM9KTuylv5uL4cOa5s76xmPP4OL1nvgPBHZm9yps+s1EpRuUOIjbaP
GSLRqKN20ZDM+oN3GezAXxvs8FsbMmeJxgJcpKercETEiucFfJveAdK/MFw/8hxT
Y+l+u1hfaj8a2p4ZewxGnlCgul7mI/F5yIHJFouioON2GlTu/2cyblw8bp3ibJI2
lapYJJleN/QPtXyU50OI+OsxEsNXJ9ujWlkT28cMekAPpax4al8JDN+Hzkhy5SJe
IAeWPAR+I34brCZNyo3p+kh0GTcOU1ioA3DczN/D481i4S18VCWH3UHjP9kulrbx
xG+/cpwOB0xv24l8vRdNBeTveqUf3/rgjVgoLn5yIn9SLxw8RJU6pkBoaQJ4tgua
zeBwh913aX8EWQtVHbVtNiksg29u6M4y6aayTRhCLOhR2yipbtUDq9icxCjyvZSm
HSje0glk6mmbYAkQKbLspIzL7mnfReFM+LoNAMK+WM+VGTwj4WmIvcBAeslVjtOC
7YNAbVI2wVHtPnITPxr6uzcL6pJvyE4dGOUQtNi1BGSAVi6op+JiRunq9EjKU0Z8
yQTsURm2MuVMkl12deHAsQazon7XGBwcMU0HhKQ5MzdLkx/9QdlukayQWS7ChGvf
aMvsTa/GEtGtCzoc+Iz/64PWVZlxsqMu0ie/t7Cid+tsczZ3VWot3pUKXRPXmcwb
AgFLW0Ni31f+9MFCy3wyJ60zSZA/w9whpcHb/BmUh82qraGCDamL12v2Dw4rJG2m
rkwQ7lmDY5V5p5F5zhbemf7eKIHlKTKNwY4kR9wqpPwkRex6raOcluxW33ZWJ/Ve
CcwWpDhYrgNlk1y1Mp3KUbGRMCoLNdmCOt1qa7JK/Mk4WChrGzNvLD8mN5yib9D6
FA2Q2EY5dMhFnt8G466D4NQ/wVDbTeL5ZEFwqEQi+VPqPWUfKlLiJ4nZZSKEv50n
VFiTwRLf9F/NfgqQDuwf+pVPW7pk7z6nf/1G7sz9MDM/0BSpHHG/2MReJwlrUFQ8
M7pf7nLUmqdG5nC1XXOAQepO1ppU3KJAX6CLbqwSWwRbEEzhx7eDRmcCFcKfTir+
V5Yp8Mr+Q/QsjpWTarpJkpjafcVqiFQJvSJP/RvXL23O545T0jjk+vUbmm0O1hWq
1urDvGEXVKRI09pqqaDnV8KV9ZfRwMnnx9ObXtx/jZy4S56/rFwWQyGCURZSqvcV
4jmFCcmpb0H07wJ8AiJzDdPDbJVZ+0PghNvq5AVRqmgM2GFBbGGLz+YlWm0vD+JI
s+cMTJL4bazXk+PJbodQ9S71HM4oj5RjjN02/FDjYylGMCeI977Z0W29/O+feqY7
dB9WQKhduaYLNLu91WH/AZX23KsBlVBU2vqPA1FmFZxVk+KK+VRYn4t1YpN1P+GQ
bm85b/sBO9som8cGzS4AR7tSwC3zUwkfzDTlHCq+pK1yqev0FiAYupopmROelxwc
tPSRuVIaSmIOkAlXvv7+DednoD+jJqv488+OfdnsSXMNnMPTcXVQZ62m65x3qtfW
2z11TUHVFpOHQURtcFpZhLZ2pc1fQh2QKVTz4y5JlUeM3CE7wFCoDJGeLax9X8QF
/JsUbiQwVwTSkUuD5LNKWQJkKqj2cA2nBTg4Z0qd7F7/s96FsQ85GQ2MwmO9wnCt
IeQHaQ6geAuCHYoNdQfQzUqJOk9MH5mKShAuCyRl0UcmMWr3KLBzBXb+IqOH0elA
+GDN1dpRyWw4UhP66Cpmd+qnHDK2EKchRupVaVBBbKgALybCFyEtauDKsVjp2GOb
lx+qUliWIvrrJkp/zFvJVS+ecPhrYSufN1hB3oMMfeWRsWjwzLI8eqo+gfRgmhQr
zX3RTmXvLrXNa1rMxhq6nUgC62t/R13d5zuowQTbmM8x4h3Jq2yQIryFx98FrVt3
yiTeHFq4wQKJcAUcRzA7BmRIVrjndKYASzjty6ImiPNna/Vi6fdaY2XhV4Sv10qP
I0noAflRD+5c8ax1WQIXfAti0aLBoungVAl96hF6LhCgxo0rdqZo4vAhKHM+8cFs
v7OWA/fv4Thj/jhWes4EDsJ5hKa7fLhjfcq2cG5QeMs034rMF5HPJhTV4YxyS+hg
qPRrNlorl1TavIamlB/r48inhbX3kHLiC1ffSzv9FrTsfj4rQCI1Kbi+JHsQx3k2
t33csJwX/dniP3783Ffcvtb/KMxtd99XLF9ofHQ0ly5odO7VPDTc+I0IJLD4rPTs
tNoFyvJP17aqTKvMDfJM6Hy7h/x172FvFbl0m95mhDJY+tVoH9I0+CJ9JzN8klAT
7soHl14mhfLtK7EGTksi1EWscAXUElRZk0ArZxWDwSgF3EpWBPSnO4pdo1GkTYkE
ZE8a5ht5QyJb36uXKDAf2raCqhJeNLwRU71jNwHU9/6NhxbmmJrfoYfMZHXqeXXL
pSogsh2rWYiip+Rja4KxxNbtQA52dYBasPSos8t8vkW9ySZo+bg0QodxAV+YfP6w
zp6UhSZLNS+uC7pV56EqYUFe2hBpMTBvQ6VGLw89oY+/gHQemwzad8bzJyK7o6HJ
a089hxfur7yluy1HlAmHWsUuoAfOJqE19DY9nMDZ37b5LEIMi9n1JUFiXao8mWTV
C0y9QvC/LeNFh7FgX9aNxifHn/EdVQk+nUDWM0ESgQzxYSA2bQZO7RTEpPeicglG
s5VVkH3iZ+xPdeszprtVajdKz+qxQRpoFT6R5xk1DL6cCRgIFrqWiWGja8rMAU6Z
mKD75A4mVvxekRVLK55dKt2nFPmwAflPYbhx7VJLGU3dWGxIRSD/4lb6F9guYFcJ
N4mEV84bxHLEHlj+TnYGyB8H8Ta2WbZwaofrngn/BNNFcUVXDwQ/nVY92a2FVmwZ
yalhp2yXu25iHIfWr+vFhlRYmUTjBUovWmMOvbte07sCX3a6diNFXMrI9gBe5cY7
NkSvUKnEO9piGGejiidVViaWdFtHhqdNzcPxo1+lO9Lm1giNElJyKn7j3LjE47Nk
u3tMcK/BM+QjKd7bQqVbPS6Kf5jVyfVktDUV8F+0M7gb7QEmQ78Gfx0Jd+wzyGn3
SGr+fNOpcsz0HXtVG53o5q2cmE8s+7d/cVLGIkoLb2gB3c3/P9IFTPWylo2nRUnZ
ZGPfoWdn0nowLsk6WNsCqm/HYAbDAYiPGgYLuH1bJWpQpvprhq5UEyq+k+Od0yZr
AvhBJvbvGSxk1J+4E0ipEEQk/o60s/6oMXBccr/6aEQ+UwznTVMVQCoesY/nhgxU
FG6cPWyCQXJWQLbVUhbHXtRf13REYtUDhutlE6Jskr1I0xNDzH2CmzTfTMYM9ggq
cahYORd32NhNFUPvBHCUMGJaSiYRPDkvfCliqUzXbMuIe38DhJmuOKClxQyEcYWS
AE0JzdyIFauNsaAixUslFGkZFaDNwuGqNg/C7/yPJJuvxzCZpOu+OgssQX6dLUF/
c4FJPTb+OVVhe69j8B9GPArI1iuUXeOM3KHyPqDSpGxiDJVz6gcvJZz7fmvTgpaW
cWDNmG/xUwCE8zgZgjq+HdbMnNbD/AH/E38xuLQAMHZHJx7p1l6QOwQrOel1fEsL
78/OOxat+4XyXlQj8nWHxwOGtX9QZg49LrGkQ6Cv2Zynd3L5YhPKv7L5sR+c5fml
2ZlU2QI5BS7C5szzF1ZFieVmAfryDdJPP7hDKd4ZI/t6HH5zKzjCvkLhI/Aq4ElL
VJdTfvlDpB1bbE+ezEXhLwG1AZ7BRpPgNmxHDKXrLN6oa8ORtuUUPqgG7eOp0YeR
meI/Y6nQQlTN9XNTjFpDEsDaiBexDd2iXHnzEmcVOI0gFGfJqjfrjEbNgX4inxYn
ffIO2lPLjgz5Kd5srGGfHLJzPSbdGTeGvLjWV+rdiO7UInXpFD1mhAHwnEl3i/n5
D73OavhmJU13OBO8uQcJZiTQAZQQ9pJs0963q7QwKQx7NCv4mAcct9p4MT7efi3t
WzzPWaRku/Bv9pOZoOHUrE/ZxsaDYo4s/rd5Fi/KO/loivHMkKj2JXH+wTACO6hj
7bTRWua8e+MhS6kyEd512GngZI69XcoERLcaNZEdyZVH0JCO2Qo8lINadRdwc1d5
5jnWfG4YgatF+/w5xF2TCCv8R3ci0WgFwjM29i/XHtIXWQMSaMmsTR6KiWYo2hm0
67JFicS4ObVCbLfxr5my7vcFczIDIoasUdxxYUkIp6RSVuLpJvOmR5MjB6VoXd8D
6WF2IiMHPZTB/hHTkotJzcb/V+87E4p8dPC6A6shGX2VBHOINAYoo5mpujcVp7F2
ByXfm9oUHdTbUTzMxaYvSHP3QNx5WT64PXY87O2JbYXDuLDS3pzcF79WUj1T8yA+
3ALmq5dvG8VJ4iXzw43Wiu9bNdYWPjIC99I6ONvyaE1/pt0ucIsfqlraDKBI0YKN
LgEOS/1JUlcGuEE1FDWJZ6B0zHHJZSOj5Ci82r6/GMd4giz+vccNddZq3O1YhigM
4sOO2WIKAdkTI0oMIP9NUGCp1Qr9aWqSJW7JMvc/rF7rs/TV1vcZLthXPQH80h7N
mGeW069lzdqJIVqa6Z/ki1BAadbgo/NHluQpSrpai4x4PFe9VWYRA7iwUllMh6ni
JUhaC1zA10SAGmicyuIK3/Q+6j0AHBoxaW+kguy3iXAlHApaNIZimY/I0v/s++Wp
nbiz+lnTvCb3o4LJmQ2ZdbQyBuJ6CQH6WQkVjqalmpiw5Rg8HyBzvi9lmkIfhEPl
C8c/V3E1k1QL+LU3dGMKWCFa360lU0NJj8x4AWcI4PQtsLXhd67umZq3sfWvjx2Q
4v0pTh9ihr4LGTmj2bYaTn8zVVFPCv/qH2TiT3bdKmdXU4ohAHVTD3Q+YZR42eE9
7ytkAN7r2ipB3JD7vA9JkcAyxwKBQs3n0uPmADE4WLqmqpqGkcWk3hn6pCgMzoYV
tL3h+6dypMkWMhsq53LiDepStkA3v5Fc6IbFWDlZ2z0GyAD1VTvppM2GJahrKDzv
szPT2ErTMEvNWL+gulkzz24fx0RKX45cpJZuS2iw2s50QnSnNdJO5G9PbWbi2r8g
fipy2ZMimLiFsY93AqbDoOUbM8BRqW8pbMmocTdyrxOvlVtcwEh52BObrN8ytNAI
eyxAvttixBytg0AcDeDsKCYnGLXxupBinAoGMWHplQbFnu6irVMIWKGHA3GZtWhK
zK1RcAbsxSyfzpH2Sn2wLigfXKlhsA2KMY6KVPDHsGSMr+RQqCpKXSFdSLy1n1s7
uJodZYoY9f9GIrvroCHQTmlr21aZg1EJvJnH8hbx0OL3kaPphedDmHY59zRKypQd
JebpVwu+JKahIJi3CZo8P8bNZUXe/F3vtQYfuAnA2CCeBZkFPIoFdx9pl4wxK8kD
s8lThKIeWAIZtC8Y+2BWsmRCW4JRbAn7m/KReVy/KlZJDFhn4GcXvmSCRbb2G8iU
N4bNO2bSb+LxL4qLDa38FmAUtp+xvT+1fhZjuT4niDYq1l7O7pNrqDh/cv9rRgki
/bOXzNitN0XqDW/+E1Ibmo5R7LPrHJxKj2xk5HRiiRBOS16kJ3l/2Ai0zk1N2B5f
pLB++6lTtKzzJVoZg/m8l5T/MLBIDhcrmR096jm16pEc70exFN/o8xfPGYbRSJae
T6INpT+zJBRCzCHqgFzgBoOT8L73wbpuk+pH5u/UULEe/iTZdbiZPJQQ+R8jxw0e
RrE1DtzbgAxgdE92j0BT16py2B4TJl7+QsEDcgHK6LgVmoeDq0bd5ehg5r0hpCXM
BwsVCwS9CibVENCzBoi9oky4w7fdAoCSGErgWa3maETP2oTwvOVhWMZS+7ZyT9wg
9pmTdsLLFZVcXkaGO0NPT9oYzazduoVoaUiGUAEemLBFy1rfDRjzq2WWElfhdtDf
e/3HdB3mc4wCnw+OCvT6IIhcQi/zo/I0TwPO1LwYY8+ALqdGx7wO4MwQZTJm2ANh
ypPzfDsOcTD6D7rYTvg969IItuD/5LcpXAM256HDHv1p+j9OcbQczt/EfYBjnuGB
vfZCJzFCI1Ir40OWbds9NFGJBQ5r090sdeUT7Mjx13EaSZdU89ZonBlPjF/w0zsQ
Ksdm7zr6i1YPRwl3adGxN2ggmq+oB9Y3CCTviBC5Jw8gVbORYsdfrDYZgt7qesau
9YZxCneBCZIx6uvnKGdZnPKqeoRcrVGVPWFGILY863x65oT1Pz0kGuDpNbV5BJZe
M/E8kYHHysbnd8uT4Pj4qAE+LwnoOcO7X0PelvtW9GZrN98oUTvR7lIpeKqwQPZw
2mEwW/8W5aa5JyxNw+LsXqISvGTJFfg9TjI90Js5k2z8mLxpP9OxDEgHZX7F29JC
WpsQUrxAaKzCBd63AA2EWAq2QGly5zXtbQ0GyoNPGhlLrrODu1TVY85aUkIRNppB
2HMGdi3PZVZUASqW/jnQLWApmkCrb1G41YumY34ltitdRx73q+DNx73NAubWaExO
avCm68ie9YcZOp19TXPy3ZuwJXvKa+ggAtWT96o/mYpddTMmzUe44hRamNtKJJn6
8aR45TRkxbS2D+usge/HaW7SQy2Tcrxzm+wXsvXV0CnEgr/kmJDKhDnpGDaXkwYQ
nV70H1f6LinTymBuckc996rw97ZK2f23bMFx/2pcB/gfLwmrxqn8gDXzb1nOtNkH
/KgvtYcGkFwZY8orFqAN4XApd+anONflLIHWbZHToJaFuN1UlQkURKBl3fL3oGQ8
hYWgjQUAYMsprl+spa1YDvv4a7ved0h35V0bjm3uyw2o9y+zPRzCsmOVHs3UOB//
DlsvsCZRztmIn6sBQ2Otv/kEw56ob7TnEdTdBPBkCgC4xJCaF33K9C3birM8lPlN
KVLmGBDlIywvu6I6zLBYuMgl+a3hwR2ZbckQwJ6f7MFSn8kkqFuGMC+3IkJTbrAV
eLClmNKNvVWVG5vyyf2vWq2YHOCXFD3TyL8nE1JWAq4/7YPqFqSw5RCe1QORGlJz
Esv3lZFJ1jJGT3P3OOQMtE3W0/CquuhpFYchs4/JRLhigS4y5oy5VYFNHC04A6Q2
m5gGZEatUhjKvJdfVlENnpDqxbzB4nSVe8A1MlnwhcKDNjEqMFa4ukgu9XjyGH6D
yr+u6NcVG346qi9V1BEJRBzPTYENi3ot4EWMvqvXk92WPNUzPVm5y8qfqT1ZS59p
Ao//gBpXCCg5A1eHRYXIKZjGNqeV6wfCmF1gg1bm3iuynfJt0xYKInSrgMEVsjDZ
2EPOZRb5sIP2Prn2lDglemISlZq7NItld9yjadUqAioC9md8OQU6bakDcisFbboX
3Y7czGwQ52eBIJYTorcSpjt34jeUhmd1Py3LIjed3qJdmy9IscD+MmMOKliYbj+q
y6WKCkThFPo08GNO2j1GCJoNSSOJTzuBu/us+6G11H5k97ZWWzwfSdfQaOIKldur
sY/VzqvlagjsNXv3haQUfp9XJGYfC+c7NUg4V/lDRxX++nUrYaFaqDEhjdZeUQUW
Cir2Ynl/rXEEpGtKf98+wUgXk3DuB15OtULiOO87i8o6ezwPX9CHedvA8P8HiZ23
muBUOQebMCOQFYn7i/yzTy8lzB7Zd8xTYBQrm44fw0NyLFOwiBrBGcbFnSo08iLr
RbryLOeIXqFJnDSX5losS1zMBL8lWKHf6ZdpnxYfrgnPC1fPLHLJcO9E2aoWTGLK
gDzWzgKZyZXkCMMy8mReJqKv3KcarMqoN2GptSKy/rXIg4Zf1Trbjnrr/7KLdSn0
3+NTNU/b4e+hnr9JqGBk38PefYO/rBZKhepNqn6Fm2ikIAPFWb2bqix3CqP2bNCD
fKY18c4KlyNgWLGcYq8vkiNA3vpgtOa0sa7XtGKiU8xjeUN6u75P8WASKHmx4ZVN
hHGe5ko0h4UPX4o+YbFYNTREBXF5Le9H7Qe09xgTo6vfuiRReaRtE83D55G3fZTc
fLUynoiGLFJ0yAtjxZRjX2Y64SsDQQvWv8PUW5jZexumujBcnAoisuRVnfs4Q01/
Fh19f4ovegAhf0tDOh5IBSS8OpueKgizl1FKp7WltFJ1x32ucN3BSoSaf06bmsYT
07UXFaGXP9wJ5XyDNjmDTAfkK6efJ4QFHdcQFkoLWfJf1Me595k9cXSqnoaXlItf
XVACRhEeKmFkOt9ErlslVsbeCOaBicpkR0wJh8aWO7RbVTOpQ7BU6Vxp5cUY7+zH
NCQ5er+YjWLqobWT49ubOZ7HRCUMDdU+ya5XtcOtjicuxQPVRmf6qv04sYRbYjyw
V7NjP8t3rCNs5aNE60BH8QdmwOy76OmpTXg0TrlYDOtd2LgQsNbdT2Z/ze+2JawM
jwmlOFvy5+IlaLU5oWUjgSkJlfiTl942ghgci+IConsCiHERmcu4y3zttFbHy5sQ
KdSBreeLzS6B6Mt1qzAlNvT8/sfQ0gFmaAiy3F6v2YOVjW91FY+vg6G5yrDx4Kuo
t+GJao57OHNdrLYN1nNmQOkjiDM3ttkMOmPkICI4jFK+qqbNZwuJwCK0VSUHAyxH
l/1sqptH7wRoR3CSbOgAasCsadf1pVlOcHG56U8Nbfg6x5UwPedlJH8pEr96/0cj
z33odAZ0bqhtXPvxC7M4gNlaef1r11hbiIV5V8BmuhP+5mZdX+ISItrueb0Ox3Nl
Xmm4iBznTjr8jmhcestroZgiEHBAsMRW6+VNU1OmKZUJU1aMlkSozukb45pxSAHx
IeG0yyWG8KsL25Nie2WNqCTXgZHcHx4USZoIpES/XRnUS7C13TlNs0r7jn/PFMlL
rMbviL66KPZTR0aYMKbiyYiM1ZSmGBTRMZnWxm9S3ozjR+mUtP+P+lXOtgLlPdk/
oaA4u7P5l+TYBBE0hOqDttLsogPjJWA6Xe1apdWMyTE9z/3/8Vlmei5+hzSWYax+
7AbH/NCqxH4tLIcIOeNfhuCXsI8TDcIhd6jHpLWH4x7o345VQN16XNDfm/7QWTdn
nQyT4Fqcvr5o7EMfYSdk/1ZUC6C99R3wC2Izj7/vzaRa9yArZlxgFOSGLrBquVAI
rCux5MXg1KYDCHlq9BGsOVq/QDiM+Vvjpcl6i3OparJHiRSL070cd2TkszfiF7SW
HFB6jMZfSM3IRqtGFu86nedUkAdRxiML7g7/miH2HUofq21C4WzzzgTegqDlv67x
T5ls36GNqYSFFiOwMEpUA+mgYCpfwD1TwOZQWfm5UYflXOWG6VPypy3uCJpLfgs9
uiQQIpgNLMGK8r48cUelooPzZvNAPiw7CZYSGCQPr6XeKiBkm8BTALoR51ZIKW4I
QVFfmo2RvSWCXfD4nwhSBh+hL9FbsuuY1sXz3xi/+kLl2+mniz6m6fRp+FUlEYEw
QlzhkUZoOd6I9l2IoZs93RJL/4WC9Nm/FGqvqRtz8Q5tS2aifmyFS9Ag6+ug3wGZ
oqGPPJOJr6azvjBPKl/Qesegmp9G0xhSVwsUKpuWB4SkhSjxppHAf75rHBlpjS4Q
9h3uv6RsIvQRdUSaVUMK9g2Oi5VEpt70MaPfKuVQ4/OP80pd7NrZUXyICFAihz34
jQxfWYTX0ptg7nbOaobt9/OkRkbHs+5sQIbN7uKmG3TmkRWgWPqPC7NAoBvLe27k
q+5FlDApWdUiIKEfXQ0dfGh70Vv+l6sUJlcxH1ieLBw/gw5JRnjGEFr6/Ofiqt6f
A/ig14dTwI80c8BfV2LdjTvGYRNF1YI0C+wyZ4Ec4M/Agb9Z5ctzhjNPyx6OJZuD
LBuWlCo7UvkZithcOF/tHWp/p8D0f93N7Awxrlonp3TY/NOSR/NeDFE28ah83Eop
ESy+cKAl20cFRGhiFsjwx6NawEA54G2R3vJZz1pxxfCgGgezjIf/DoJ1JmGX/9r2
BWSdpCEBjzyPNeTVEfwXkzDS0JF5mnj6qQ5Hah/xrs12bCnhkhDo5D0zTYKM4hk2
s6UhR2Nj3voTvRGC5g8VGPokfGtue+eVSHIPu2qq9EE03MP1bMkMUyrjtCOggjSg
6HAe1BeD5bqhwaxwYbmQs5wm+QG+pl2Ye952khEFfWyp3JXzlK/dtj/GxXVrWZkD
1s3vBh9PZxCKkN4I8Y57JWyD3VSFt0j0j+4RF0gXRiAOuQjH9RuxAArPJ5rAC/Mj
sHSLx9o1sqSWO5Lu7cxrPNlXKdL8Gp6XFeTSu98LDuF2h+STyUmJZ7smEJrVqBRs
Dbt0+GuRVFXETMfH/l25ucZhUOTA/hJwfHJ4JEqIMJzp1jVEfSvSBAEPuOw9wXb5
QrcyAv29gDqNAQ5LWuToSfhtgRcGc7ucZj2gNIkIHIecgaoIRX/A1VyWUQZMZsi5
taHsV0kYnNVJfiAIDSp9gNL0gFD9MjRkpv8/kj33o9axIkoD+CAl39IS5KBux3zX
uH8dXoWwd/Lg/ICUP95fXQLQRuhLk1dXQ06po/KKMJaf3A/Q1ges150oGudCUCY1
mwcWkIAm+6Ya9do+gkMw3MOkQHS7IZQtTkD8rkPWG1C2BE4L6OcS+5vFkl4/N5+A
VLAwwEvi+OtMdBDumBF+Z7mzRHqunye4X3JipSUrziCJf7dm01vUgdgaysImMp/Z
O3bR8My4eg4/U9XDZ8ZqL6K+MPZlEVMoe71tpwpdJC5uo28cvznpcOD1xfXiGxif
3eC3Womy1kUyc4++dy03EUO44P1OYNqmDaaaf0S4tGDHZy+2Bkae/mBNkK1dPPW6
ByD6Uqnztmu+Vm4vGLSmkixYkw3BOH0ZLmjMqEVBvPhq9MtHrtOA2Y3wJ7HM0uY3
umfnS/25RAGwPbxXtQLx8MziUOs82pz39H7NKxdReUK0RA5F0V2mXJs3wNqIBQAa
LM+JPfChfxD8cVVl/Wk6JTQ1b+HshaMA8iPEx1sukB+vZhUxRHRPYt/OIbkaE0Ue
THqLSrx2482Sc1KAWN87KwjrpGGyjRRWjdaZZhUlStKDQriiGmEVV1HBwIomtm/A
o8819pMIZRcy6FJIcOfq0TuNf6ftWk49Chx8smsL/g7wHs18hPiq9Wipv852UpYJ
iKT3srg2c/SuHXhVDqiwEFNneXIGGdWACzvGFUhMU7wJY2uUgPyR112SjbIYs5VU
q2em+rrhb8DNwgis8P1koWVNkxCzOCW1rXy9TPxjrH3uoloTPyINt2yl+8J6Ld+P
5T5OupCyERWVyfq/tsKdh5Ezu7k/8B1umJRyrnUh5s4c07TxookHdNGq/d5ny8A4
mwuPGxFk8P1g9msXw5IXtKmbTfEkJ59M1qtkXp+aeDEKtiEwGEzUPuCbn+sXgfEj
oBs6mQd+o610Sy/Bz1wHsbBISeCqn8LqlkqiINlZRpGhGIBt7WYXvhsVSgaJc7lt
18QRmEscGQa/cVNQOTrFnPeqFCIKsMsGBZhDD5hdi8GaUiDfmZC2t3jw4snQODsZ
+NvVHX3wOnDE4xUVAzaoaxRpiMPv2H9dMQIBmn0YcoXwWRb6hLTXmhvvRm3JluAe
T59NAVgojKwsj/TITu48KVIAhA/UYFDGlwPZ1xeOMNpJRZhMUkXwfbL6CfGoMpcW
xqvgS2fWSDQR2PkQ4YS32gYvH3v2QalngRXXmAl9axbLd5nY+DdCjw+VicBCwHwS
KUOrSbDFQnesllJ/chvgl2R+GjZBFFyLwePdFgXSpIc59TYscK60xXjM8ytbkSaZ
PkffLayvGh/egS33nGyO6k/Pd+WYoEaCO9rKZfZkQaGTRMXzoUjKHuwXHBJDAysY
ZB7tDePGsOLOxjFdtOEnutfatI+LKBevDJSEJg8+7mkOhyVYUMTb52J/e+IiksEI
KbTCSNA3cUxw23IduYlJBIqWy0OdZ7X1ZAKP4l3P2PTK6HF/4hLw98VS1HRlTQ3A
JmaNuwugCvesPMDat1fbX2gwJZpMU/ZfVz7NGT8GgXRVovshHY/MnfqFv+zGPBw4
wkKqsl8OVc81PKG4qKCBSPqyT+rLoDLwKjdDVY7+1lMWgDFdobRVcVfdW+EXeK/i
GP/hMzgsuz0sfarLcHRtRXz2CCeTDoOKryLurIqZFO5fWSyiMHTi4z255qjWIEc3
eXDyu4rOFBEOY9vY9fTAHqhaBmiu2ydksVKlR3MU6nliXcAVdbuDqVdcE5Xl6QCw
N4V/lz93Bnb4t0LctlbF0L8xWf7wuFh6SpWmDswDrf0hsmKc1ybXtPrXk1eiFMJG
LVdHVxSG+f/72mhlkGHD6QD52jlTyTpQN2hTGkoMxdCOAQ4viDkEKdzLps1moYSh
aw4lzfpw9QbuCRlZNsCqUn3Inbz7ApEg9HccV+ATo7oPbKZqUwkOzRcZuwuR40fY
8aDZuOIc77BgDe2Zts7t5anTnO8oLg3oOcwSXpxxjGp8Zhht1UIgUQtUkeWb15nB
5kkkxOyy1jX5YRuWwG9IAhPi8cvXx8xdgJikWhJ7VFwbXCTQRkyBEzW4wz+bV+bO
GovSCgxSHmZwnmqVQZsL0/drC9z+nTVu5ROvnxMAGJIQ7enCdPAbH6taPUEc62Cu
7vUIbp/G0ielnECwx2GmBnG6u0/Oe8ZcHZclwLJ7PbPngMH3hwzn3zfBgFmhX4w/
3rwzbbvyjkSIDwQvlp6bo25WKo9hGFOzgGVXBafSVOqzTkmdSWsaMD+h6JWUTQtO
Eye3gm48q7EbvFHe6VJG6IuEsJFtFwwHqdKZcXIeMV0aGVPni8Ih7O2S97q62T/j
coMJU4S23c2hdtFpa2RpRSLgNsRfXTMNSa2ZBGd6KA0ZkVp7p9mDjcwwQx2VivPN
6Psb6FfTZqIbyvbBgWLwtOs9ud/N7ozg8LdjeM8pxa86geeLYpaXJ110FG4qMA7Y
CnS7InDOhXx/N28muEAVmdrkFqHryGO5eDDfARRKM1KoiPyqaJv8c38x0igFpSws
lyUr0HibHdaaC+vMhADEAQzgETp3zUgeos3tr9midQLBNEMv4PWtrZ+olxQieay/
GHHyFQqEY4bBLvRVR8bHwbamQ8L8SN75gY6Wraw/shyqH6oYLRui1NNUnwNX9MEC
Sy392BBnm+oCtuY3quVQZZbVyM0yO8aUaPkGSt1dRd6k3yO5lAjMWN6XLGEJSvz1
5yDed6LWCvS9SVwLMwlDcf6VOVq4rQH46mgIiF40f/lQ/b+3mzS8Y8CFPRj0cSoW
Dmw0MCBlev4H310IIyL+3dcM+Rc7TWnWiPZxQz5NGhhrncr2nDflOaoqS+lPydUH
qemJV29kMeGjynqlKp6i52afBqniGhRzqnhgQHl9NrLxMuZLpdo3/3dukLgkVDJx
YDlFmfxbX/1dwNRlPgJ5oa3aTsp4oj9Qb44vZ+42f4i7IKYmA1THYhLGaIfkNQ9e
kBbw8U3Q9emZmoj9HgqvL2xOyQbm21LnXbSCwGtkjqKBeOJZhJ1cDqFVX4iPhrRm
dEM02FR4lS/ak+KRZE/DLuyyFpUt4A/6fQKFe++7MWKGz75OIEpIUynfT3GuSXY9
scrg6W2RefX7rZysOOQr+T2J1+36v6EoQvra125FX6quNBoPsdsVoDAPquf4uXOw
axMwwINM2Uut9FltoAMwT25X7VDYEryhf+qtC/yiKLm+hZTMwA1WR1VDAB+pZcya
fghVdLR0fGzTrfGuZ1cyuTLPFRvU//ysDfJaYZI1CViB3b7jhNy+2WsjZJlzgRDo
lchUbEg2rXAcnUiuwo0Jm6Pp658Kyl4f5V2uccAd0rDTRUyp86yhuELPzB9WPLuO
j9wlp/D750RQ5RYdmxrkd3GpWdLY/+OWDfOJkMcK/QuMAhuc8aIuknPSkVl0n10R
NUDD6mcWpd7Gx+/qBdB3xsWj12hRkx+q01YZswH1D96E6ZVUXz01mRpc8V9ucymU
ey5CfnuUIEdcIHF+ZQBt0MtQC9iaxTON0pEBiy2ixehXGTDiq+EcbjTot/Gw9mGy
3kC6LNmSRYk/Nh7c6u+UiWuDI4eeKtlpbTLoZ2ZNcrShQNRBu7bTOVvo1cD0LH0W
JNQzLMUDlCTSj6iiiu204uNAMkALTTeH6xJiAohCDEMYISRHA1RMvAQlFYMFfp3b
ey/DePvkIsaue45JMycbYtj1OQh8e7PvWFkUrhW4hibneRWiT4qpfQIpceTIm5P8
IQFvBZbXdieS4KtFTLcgCpLkD79GBLjajhHONFjxnzzuYPKFdwuNN0b2adEfs+Ct
GKPLeeEJCyDNCDlJwThHt4xqz1fPEAh8TYTrHFJc6TuJUlLPaULZs+12cSkh/Ep2
QWVtrKOZz+PP82+2a9/8zlerZgO/s6UiSweIE8tqxd73KAfT+SW5RyTDLFKdYiOz
AofGZ1MCYtFuFoTyfReJdEXgrbjF2AMhpBBKKN0TXH26U5AZAb9VuqTBCfeKgFM0
DspVHJis85YbHEDSlohOC9IWfYdZOLbDvh7CRqLJv6BMuor0Jp9z963Sh1F945RA
/qp7AH8NWqLTz34CWMj+gP+OZcw1ITFZFH4YyU66EQmWAnkE2tIIP7a9nUcQIlCH
epz8Ix96EAoRIAe0uhTfr3aUjPQla1PVG195m4ViTZ3SHLBYN/EHYimEhH4jgRuQ
Y+QW22Hv9GHEJpTk8rfEYmaX3UbPpBKA6WgYC2p+TotmgXhG7UCqFfB/XlPEsC2G
AVZg2bDZOnjCEmH1nltamCOGWkSTHjI/a1azGLvIa9dOhEEISAajtL4jMHdLPYrR
DcoQn03IUyxWBGnJJ/kToIjc4rOBP6dFjrMKl4Y9awEusyfwCtor/fqqWyX2rz/0
sjvcPTS1vqF+6MuLsPm6qGvPuWXtrfrzcMJt71KcDJ2Fwu8+QvAVSXhJab5X8E1e
XR6wS20vs1jGKBYUKXZw1drbjTii5b7hO5qVnUc6t7Oz/ZiZTmURGu4hex6K6Nfb
RrKD3BqXKVYMcyZ732SX5oDjSWtg+y1/do721HRmVJnl14v1V0UEa8SNsceIVJlY
ShTyIY+A6h+zUYvHj1bSZrZ946CmHEERVH4aDt+ehzDDq8V1K5OsydsoArHKTciZ
pdTOnsfqOBHdrDmeK/enuWEpbhlaZ0WCXd0ZbxtAUsCrmsPMPVpipJxnW79gTw+g
uaqBqnSODzDhcQTCtnCg+hpB6JYcwNG/A8vBd+TQrRSWZTA1oqoCyaX07lcRfxJx
lq04JiqmoJY5F4eqfIQ844SIw62ogJiUlJfz7UPy0sJG3BQW1ABSBYkF5UmIOkUx
kfkTjIOz9+LbyWjSvkivQQKM+WeGaNA6fzBdm/mnly+oCu5TfhKpCHdQwk5rmUVd
4UIwEd9TCe4LD/rBPdyf5sNd9/XZT93r3ffMIRMKbcbvd8ZfypL4jKL7xbIoirVs
0okRAty3rxQNdgI1r307kr29QJcdJEESsdLmrDNzY5+DLDPiG9QpIElDZzj9im97
QWPvIMVpf2EvrKWosRRUNpV5auSylZa/YI//Q1KFC0jkSNxUz1qvld5VhP6AOpnL
wWJJPxbSYhRYa76sIGScsU7peUF17ChVN3acykl96bfjYYlEE84TpH1CR3/fsA/B
hsJGmr5DvRhv2p65+hiL465X+NTlPc2usy0tT+tx8YNjDQYCvdQYfDCxLOdvs/TW
tsf05aypDrEdDfxEZ893qCnUzyydwqUXevb40fN5OKrEnogIMNh7CwSeL9y4uOjP
8RJVyehZNZO1iX0TOA2ikQdd/oI85iA1AJXNpyRDOsqyaLuwuKCDLr9BnCL4a+AM
YVI4ay0zzGOmq6k8kHsgiXAhM17DgsIG6asW1mc7pk1N5sIqMWFnqpkPORi1CcQR
8yFVXRiUIVVlNoozEs0est/PBT6okBHbmyan+xuDtYqNJ2M4mS5hD0BjayjfdLbI
DLwdQv3/soTSG21MBbzFu9st6ItYNW8vDrBLZA4h16HYcZAljFvIyfb0jmwmRa4f
9TrRvqRyXhcj3zhZ/Y520CBTAmjGsLNlvZOuv6nayUIblkDLNUOP1uvf675oNRRg
2Q9rJlXfixgkt9RYYxjxo8DcovOTvakhD2rxCtXd8DhlISmtZPpWqd2Yfvy3v1e7
dDdYdRVl5kbJ6ZfhI2oxFubDKRtJxnjWPGDGf6BJn+pHyjdXZCeAmPpZ6uKke9Fz
d8iDYFYdZtK9IcD5OD2AOfIwSGTJge5QUesdWc61znjQrLsgQ8vL1SbELNYpH/bE
LJSvAdZVGfQ0aXiIIFXnpcKqgutt+8hMkArjiGh8spdiiuzNTZf8lGXaSbwIyTtC
kyUGPlcqreA/hCYG4CBdorJjrrmuuqCOdNrSKy52QS4Fa+ZJdeKx3+ekV1uXYHLj
jNtb/KSSOaN1AcuztgyjZJ29BYGbQEyaNTLej4BQjM8ylzls8zfxrjeZSemMqa8L
5JVNosdI2jn621znkyE9vB7dE4gwlUjJGf2Si1ko3JKNRLEVIuXgTB8hL8tT/IDP
VCetZcJJ1kvtUmkeItKMyR5DvF4xhMVlUWHdcoSIUzwHfe1/7MQMFQ3+5OVa/yPf
daTLj6PF77cA0zh/O5jZj7nHt80iy3ZpAJ+rz8vwpvZGW9s3Lb4cBnOeP6xyer+N
+JwJdCgrTTWJxr0LhsiZKY8F+5QgKHeK9ys4CU1hd5o/XsIRJrnEepwxvKFxRlg3
y5xOLUXmS3PDJLudVR5cXvxDIQdx2kQXXR9xUbNKjKcdXvrTXX2YqNbu8X1S94+b
eWPnCY1yeOjGvXkymjY2qMpBPZVP8m4lTip/yN5pTFhvqakEuXhDv2Ylnj5GfvxK
9txqrLzhpdTn/1POr0ayrrSYZFVIwwOcVZAK6Q8inG/oWOBc9rIjodkI2nHb2vKt
tFV7ynAkzybunJHs1Vq8TAq1I8mDbc/wDs7VQevAEl9gA45X5lQyXpTklzWD8+pD
xJbBbH0A/1Zhqqxx+QbBWMrW+qrk74pSA1hVp+2mb6qjMFxYkfZdCnp/GwcLaCbS
WzS+aUimss7ehO+BD/hs9pO2HA7lwMlzsPZ7E/JjFJvEx9tFwqSdkfXZftt7LLeQ
mzELCBCKCtm35qyKpXFhQzjEPXPOUHeCSWfuexPMN2xX6TLk7qE1+3LP8cQogEIx
2pSe3B4CIwvMd2rJXV35VC8/cui70Ek7ddDs0yw9LxR9L70miTfxr3MFt+MIU3CX
acO6RWPZznHJG7gRceK2UPVekLaunBqPmWG961py73pEDgCQWSZEaEzPEgWGiAw2
6p4iETWOSN26tsgIaTIF1M0wLKZVa7guy5uryRC2alNa1foSy8TB2rpH8CXW9tvj
FLhfQEVE+uMtAYoXzimtlHaK5aZ8DzMtFc9qleFKhxVWEywPqZj6rQlsAaDq6HGK
tsTB5j+dW0OM/hMreqrnAEuNaJFmDG09kcxX4YDHX0kCGc98O1vd/vubfWV55rI6
csU4IGZTGjx/Xst+D74ID9viUhOjrlC0Fkhfz9m36k3+YbvLmObo0OEooyvImI1F
uiEsb+TLpiU3xPsv/egLq9KZY9Zg1GuVLeUDhSY+YnV+47vFqVsel0F5WmAVlH2X
gNUVTdm137cOFKKWwbUk50CtZCzYOOm7Vsu5lmrzcSpx1AColE7+N2LO4q2ag2tb
n49QCJWs0NnTzLkYhGbreI6WnU+7a1HCMy8skmn5+NccyOacHq1kdIRiMucirokk
jTDzAgjAEOFjZUogsbk84i1gjjvTnZ0TWKGmcjHHDIMI2ajpbFBPC4vGaDwGJNTe
53923xE5OdTMPe3PtKKzq347XGP13KhsADde31M3TyTgybVgjEdriIy0akeEKsls
Qk/Wg/EcDR1iOusR6yBZZSUSYNclYA/D6lDQaonIsYomYEhT5iPje/C15kvru80I
vARNv1KuefssAe7JyRONFdufRtWK8oFTzysR6qlco0WwgKgAFh/BFHE971+gtGvY
X9nv5mept26kHRDvqwXRC4FrUvGLt5bf2h5ALZ/1SulvbMecSA9pQe95kz33h2NV
XLG4sjcKjwa8kCrCcqRavMlW+cPa2+B8hGcMOv0Ob8hRZjd+P55GoGRxK8ICTUfa
QykrbywTAGsj7WqjRpS1MZ6bvrhfUPmLu8NPHwMcVSj4F71UqLwo6Xgo386Vrnrb
M4tHPf5ULMgvXQtELkSiZcUJzP8x9eEAYLEsrWMOOdXde+6DGh6Zzz9boyW1qKuN
tN6zQ+DzpwXeb1Bvni6gXRJ19CtX6mc799Iy2uwUgt3wzBM8MOY+eabgJC/MMTHs
bjd+C6JoYinGLlVUPBgTFgWkLSyBx7QI7dJ77AXV03FC7khIqALpheT7Pm/Iu0Rs
vs34a+zjxdkyJh2ZFUOiWoX5YGDLwtgh7Vqf2K32WcdiNzDBvOwRnmGAcV8MgdHN
ayKt6oo/xUjPeenkWszKytDnSjg/c+25mWvIj/cfWwmyxQEjxEaVgsFtj1U937A+
JOenHG7IgWVqZqp0nIEAbduahcpBk//LUSwwSykJQ5M30dRzLCsfY7FcHoFB0073
q4i4b5DhF6DqVXDahezq5RL0tOAfxSb5i0qA5CZ2Ff96W7fyfLicaPFdfJx1z7wb
FP4lrRdPf9jqrNWjio+XpV06erTznKeGm3i0DPEEXxZxz5LhZ3QFWs8JRJRKmn4F
8ya5X1lD8IFOR3cmXmV/IVVfzhcBvyqRDiG2PxRtxGWADcaUmnHAVUtBFB3t8ajy
RjENu2KJjeNt4iSjHLSoemhmusnQ5hZKVnymAh7Z7E9dA9sSDYnA8tASRz8mixkv
/eoN/1tkN9APKxklKEvIR+BTLptMccavsbGoXTqhaA1IBgHiSL3Ixcuw0JvZiXZP
rk/VdhVovJtjI8Uffwa24SXUwvD4lP2eb1m1wcPQpnp6U173iPmGhG2dAyBr5zn1
a/m3DE6x+2UtnwqOdVTtQuitKrns6f1BepWRgKY/bJRiUvPkL7e3kKBpc6uULHu2
CFr/DuMU0PhIUFyYOb8VNCOmF+QDDcj6dky6lyiQo/QXCTYpMQQGqG7B/q459j/W
wOREh2FkfCioT9DI6ulNouEuSp2VGqihTtAdA5tQ557eo722Y5vylPcWOhvsXtqa
52OIsY05ppwzQmpKRwQArynN0qEmK/tC0mxX6+AW0LRqdqPhzOXWMMCPMS9dzL2y
qVner+6VHONt/JOPemScG9gA+kbbi1A4Ndvl5NNmfHCYT50R25Ec3nmA7ZQL72Z0
RrIALa8QQ1SctG2/lsbGRQxF9R/8a8DQ09z2uQbto9QP+0yItiABHouiZUuNdn3G
wf/ZVYGCWi6AF0F/o15bkxt3XjVN7ed118bBwezD8JySoRtPmtIyTFl56fMh/90p
TapmIdvoHCTJIhQEbheOtpe0gWcfBL0nytaYofYmQroBj8MLWdd05zcT1A02QRo6
yDJbe143OnWxaypAeA8e8ShsOKr3hxcgyay+ttV+gR0hVgw5QQ7agC0wLHLSvG73
sYpI2cN7BPhq/11UkCvhGCXeAjLpccq85FW9x/vUXDyuYKdVG/+6PcV6o5/RenC6
xrlX81ty48mEF8qYyjRFeO5uahBPq0PY6zsnuH2BM+b6nDBBqVZ2yHKH3fSFDU2v
ZhY5lYWYC6VY/iq7KGfSzFg+wlwCV6ti69Ub0gKhsZ9Zo9hUTwZi/2Lorevtrttt
pXyt5UZ9O7plvWSxOb6OmLvMR925UMHuo2Gx95qDJ3xuTFIXk5YJE5nNZzfMLlKT
288XjlrwHh/AB4+pQiCu8kOHhKzPyCO+aGM/6EDZJtezEhXluJAL1aqmrJQK3lIg
LQK3ZnqgtYPRgBnM90YKlFEVADJJSonVjE3Rtz1SYf5lAyG+1caBRlGC/kjdkq0S
xT3KeXQemc5rqddZmnjyaq2WdlkPCbt98HautsqW2/s+WUbje3FWUq7LKy9HaHga
pbZdmqGfQuw2KSfr4GgSYieJte9IR8Zb1pknSOGymITCbFKTIaswtvElk+UEOtvm
+BFyKtOGcUtWK4XvX08EoOzDl9Go/DxR5ilZ65h/Pp9uHEp8jU1wGdyqShMJ5tJo
eqK/rADRR/BE+F2d/qbN28anINYZRoUe7Xn2+uvvSth/vIiQzUr60TqRhCw1Ps5M
dp2knipsB6SqrCJV/17ShluQ3ceFa5wPlahNlWiS2rl0a4SwCKCgeIGYgZvIaI2j
fbOJ5uFBT3f19rNYJKFVTnO2kVwPCNncv//RfMHSoLadxI/O3JBfiC1W5JihkDAm
iKs2xJukyhnDuSaguAFNmzOS/lZ82v6YvLbuRJMNqUa/gmAOq9WBkW9AyA9/+pru
To46lPD2l4VlErct3odQbQhIkjW9kyT7OpqQ29EqJOZhUTJt29reusLbooragLAo
5hz+VOU0B82YL+zOUTA6B0FPUvhCa6A1tPK7Huj45BPORuSfpChgqSNVvqipY7D6
dsSJPn6XpLKyyXUIhVJLwUWr0eI4wNeiEddtMHZEefmG9J3QNhNaQIQ+IIraGHrH
AA0i21yEAwpV/YiSLZyIOgb0urGuMDljZB7g0lIXN33lgCEDwajk/qcDDKC/P8QG
xHEvkyI0v1xZRcg6vz0yoJADudAKO7u7rRidl249m5NgX1s338Rzzrd9AQ6T2ZKM
f8zszXZw2j+7CDm4ukmpMA1eYCQ34bSeE3Vw4ipFsx1mA5cp3psmjHm5yy/+Tvpn
w5RjwLmo1n2HQTozJTOaoYu82/LiHX+sCfIh8qtOcSsF7DTvmHDX4TpsiGb+IcCZ
7b6+OzPeKYchybw1xmZgbXw0//5dmpLRowFSb+So5HTEyZcSgt3SKvoNJ8eNtm2c
FL4GpCCx3otQ8YoMHIErySfHA5KPCtlfglL00SWR4uze52xusTlzBGQ6ZMMEDUB0
uzZgbzjEE14efxXNAuwlaJPDWUNuAicG+UsyPVJ4236hZF0/kLT1UJsV6ihoZHn+
mZ0n70KR1QnmXIXLu56ZmQu7dT56sY9JARIxxKg7aIjVqVkWEWbE2jJhOp8mlfVM
+LxUkDXy8evPtTDHfdfg3U0/p6ymdAU8vHCRUacfGObmcWR8qK5f5oUUEvaP+IDN
uET6njsUKEfS0vLRHAyIIjrLpZ3qevzX15WIiGbWAsaS7OGe/KN3BoxBkwpqtSSW
jupmpNGT+jECZ4WowOuTQiNKNtLRHoQlqzosyJKI3PkhFTfzfW0GauJ1p0t/GDTJ
l11pxIcIvxrn1JDDSCnj5oN7WAx0uN9RG7owfUeLrBNXpIbEzpWNIkPXFGo/wSwm
Rt3JBr29tdqPERN+bxk45WulME91k2gOSVs5gWFZwtpeqgt13V6QXMcF8sjNGCvV
a/MhrRT/fqSRfDnNw0l8yLGKY6O7g9AacvEVKFqN8bJ7ecJvisMmxb9Zq261LX8K
zH9IdLuDtoFXZmrl10zSjaRGKzgGV0LGcnMLHjxRHflznryAh2VXnHtYXhT/335s
2oiwdUCW+MVFd+Sw/V1El5HU1jbFBexDTNEA8OSIvV4vu4f0Uv6fgvfz9aFqRlH8
xkAVx1jldwe0O7Eu7sCc4Ccx5BeF4T3NbrBdaOaqtrs4pdpsAZex9K/aWbQZTGY1
Mywq0yQFMQ93aBIza9FCBwKkGfB2sm1epLssmaCLFWEy0hxCqLuE09XhUqkIOX5b
+Rbpmiwf929AAqeEDP23DNRTyZZdpfepxnbMu123DGZDYAcyMaMJrckoqfntACO+
FRIOX1N8soP6drwrBJ9VWiMRjvEG4AtjR7U2bGl7gj1q8T3kGfzhVeN2q4iniSHN
SgSM5ZLYVX9RNZf95MEdohPBOZCa4F7CULQRDEwm4mlMGox3jO71BMWSF6PllPLa
kTd2VDS0kNdNkncm5SLM8COJMWKPZlyhoYVezM8vdPsyUooEUHoRD35yzTKcR5rO
+1Vq8OJQbeYot72bY6v0xIP4Ngkh1kEhIlc+IkraNTP4iKF5uzbDyid3XO3Uq7An
IuUw3qHMIMYy+HzvdYqZuLO+hh3WXSmn1Ag2fFZN74uKNYSOWUpfKnWiU7f8FoRR
UMSevKlElkCN843g2Bnw8Z8Ghu9A41cXRctjtqLyy7U4LwXLa6L40uMappbEQ6DE
p+5gkkD9gJOdgyZgkxhnOVfb7FyDmt2bqZFhd6Rjnmlnc0G2D9vrLAw1O2zB5EdW
ywMOuwtaE9rPaYm4KbTq9Vu4cf/DOoRuCNdwv4T+aI8tCXcH7fQUbd2DlBpZ05KV
Fsf8bP3SofBzy/vOxjY1sTMC+OYmh6rxBbpOxhWHBOMhDNppW1sMfLRY1rcpgMZs
rbuiOBMt80vUjp0QKLRjLCT/VOzBQhJ193GMNLfZffI0eADB9nKyLnhDy3ZWmH0R
hZqFd4XIPVEQS/22qXZlKKU7LPqKMuYqmNO8OcL6k28I/6fBO4NIdQswQRHO72g9
CQOg3PASNctJlCvr7JQZHtWRnd1ttvZsprloKkv5ThYol3buvYuM96kaWA9VqBOz
xFYvXWwzHStBzKGqBHZx+n0DMxY+ywMR6tRF5CimrpirvA8fzheEVoNVDt4pjTWn
RTHfkubkCDN5/5sBJmSzEoAyAz/VYC9j+9YI+ToexSF2sQ7EK8nqdj6JzFQV9RDQ
g0kL1nYeW0c6csf1GKthbXNPgMekL2izWJEM4unddJAYcNtelV4YahQbHhIOCF5O
oElHCdL1soML3SOoi8qRaeHjr+/0aAJN+dIBA3kBwn4RnMtkYHw6c0iL6X9rL4xW
29OpYoXuWdoLTYEKX9EEdrZasUryIVuLfwnfLL/90kitsM4m4PujAW5jT/0RJrEa
jTPReVlfHfDn1oMBwXzLgQTmg0vXRayWT2bwdJ39qZqvlM2PboYI8Yse55vgRcIm
RQNxt5DTlduS7Mw8OFH321Zi4SZaIBVsvX3a6ob7e5RVv0BDpHwTy7sAgHB3C47u
1H46tKb0b6hl3iRwQAFEy6Criim06XTX5u3qnQn3ZNaEyFsRybBYZ+MtvEBJ0U2B
TO87C5HYMJB19ArTYNAlA5Zrar4KW3EFqx3V9YLpk4//UX6/1g5+vxIgbkhd6IKd
T2WAD1xzTf1jWfxHc0vN1Bb8Evp8WsSpMdADL60tr0a3T+jYWq56u2pbVAQGvGzM
Cw0z022IzW7xtvQ/Eppgimok3I5ARC9PlZmlZWcUxWQrxKImkGYJJNG1YWFEyN7B
HHkHijcRJgDNcOoNl5B8EnaOTzwcweMlJzLrQCJ77Cv560B/EN6yKASUnyjISdon
2KcVga/GhdzxuoYy4fv4siXNFukCbq9hizYI4DvtRmH1lU+wlI8dYAck6z1DKVNU
Rdw3hs4r7EzWeLB+0Q9byZX0z7D1VWwcWAisezQqOkg9A7Pqcua4Y2xjoFq/lAdr
TSnTH7ZFtysFo69AlSus6d6Yo4vMDBo1N+d7V5x8+j2s4MW4HzhSIxXYH914b+R8
TNfVyN5/ZrlQY9OnsHUzb/uwGvMf18kUSXQ2+mX7BerrKgrVYuuPRk3lKZblMnWl
kKyexmB6qTrVFDTpj/EiNPikZLscGrxChIW3Fx7KfzzzcSnGuv4Xyk7cCR08p9nO
KtHIGql6Td00WjxUyhJaUFY4evLEu/ewTQkPhZipX1SncTZqtBft+Iaps2ZPIT2V
nv8QgWqmUvGG9mawQV/EdfjtExFa+DChAgBHdZwFllYRKXQ3SY1nB0hR6a26EjQc
B7y0jf7iQVFqYBvFCWIBCYykF5KKs93gZ4rwihmOo5mTJ51Lzvf3Su7G+ZTJnXEX
AD4mL7yAepiiS6GqZ6kRZVG+W22hQr8DUWXjLzwnH6Gqy7EQP15tbkJKyyUAYq5W
cNbR5+GIo7bVma0K919OmquRxJxjJXs62CDG96D8QBjJBk66sPRzoOdlMX/La28E
zLBLr6f0GbEOmhCzQ4FR0L0R9eJDFQZ8fD30liOUFAwxk/sz1CcuYi5lEpepNZoO
X7B8UMG7QeTtXj0tuuZZ8vXjBnjjvypBE0J/mEudntIHITH2tnGtMQuSMtUhGsMb
QYNf0XGWvm96jNRwmlLRoIfq42kSy3oK/3jIslTjhi83591AVlGNG2t5ckfXv1oF
u/NF35WBxyJBqRUR4wwpe7apJkqiyLGl0znOk+6JBtPltqE5+zkXwlTq03kGt/4U
CKFpUyx5mlWJoIc/BOvI0zLlIK8TLcDvBtOHlMqKKi13YrtEpkGxEr5gYJDFUN2y
CbichHKxnPMpAMgFZKvfZEfUykl1phdtehz2+dOi//tIpCug302f4SHMvcuvRXET
wJU26uWix9RpLU9J+caPTrjXrZ3O73PWSuExJuVURT4+fqZrf1plC1SVK9NeQdS3
8ekU1dv80DCn7wMrgSaJwRO/WPO5XO/Vl5WiEnMZpGkWkhIMe6Nqjf4GG15jMTIr
eZUHxpIiYhWMfvh0FO+XyCxPLNjReusoZYWxCFjLegrIeTQeFkuGUwh63Xwaxch4
rIXA743FH0zK2wtkvBXqCU7esn8PkcoUDqWg72nPRnxg+nm8MZJWpH+7wgImkWyu
rljU4CxCpeHCG3aHh3AYO8YaE2v4LjD5MAN+SY0H2qKsOMPYYLJLyrB9nAbP3FYa
FYZV7UT7n+SoZ4Ue30a0dwrJQdhsZlutaFoUxqzABRMpRYP3iERWxqs/7v3Tuxsk
K0O79p4hsWLSl3gSd+ErGi7FXwOxrZacT3kFU+x6kS2kPdEGvXkUKwt9jhF+AL8o
i0bm/1jcHU7JvTjI+oMU8mEKyLLawd6MYB9DxbE949jx6FU6kNFWT7qJY8KxELdH
VOXVj/0kCH8KcylEw5rNBEbFTR3Y2G4WBYFVAD/cy0tKGJO2JATXKRR5088ba6ym
0qyU+qa78zlZ/vql2+3xjjmawze2QS5FS4o6WTN4Ule17bL7jhCLRlL59RIBhnVD
8aOqyAgsaLhE9fabD19A84tM/LACBFHTm7gKQhFajdDd/RrzaaUPZxuy1b5zu7Lz
ln7piYb/De3HA9oKIT1B6DFVab8mj/Pl+pCfNq7YDULjj7IXMcOikJJv7l/aegkF
ZUqRB6zS0N7gaU53DqCHk1Bw4qKP/Acd/rUS2xFrxg96BnPie3zG3lIZh+t3+9n2
Wh1eaqlIPorjs4+xhXATDstY1L2Oj2D5f3GVX4EqmkxSbuKF2qCgHp7yhkOZE16y
L+vH3JDs9HJr5CvLoQxHtoyQSp010sNeSiumKNGYgsxnNcuu6M7i8rjJtBUpHc21
3bIG1Wstqca06i7Q1EV+gbhEONiSSeMd43Uvuf+LOJnxnx+Ox02pO7w/1Q8/INe/
74OUdwwiFF7Eqp6zg3p1I1h75V2ploR/tkOa6bgUXXVqQs94QFd/U2cCNgzVZBsy
taMMZQJAgNpACmiwfQimU2Y8jT6TRn3/dBJU9hsi5itrM7N/kWFSkDuaqcft/6v7
ryk0P3KR+JFww9lqk6mWCyOfhhJPGu7fKtm1Xk0ms0lxdHMhSEOucz+DI7cQZiRN
oR+QNMhrWcI1tPxF7ixYkZm44xdNyt2L6PZYZ3+mXASGrSMBqQEqD89+UpI3++KZ
ulIvrmY5MI3NmiiEBRVJR1XFC8SwFg/iSlAHntVmtuk7xpIn3zJ4+dLsdakblu8u
zfYWHjT8v1v5R8TwyIsDbC3L2/IiIlunjmeO0ex0qn+mCSv8mmGVpuFPa8pMEshx
PF1F8AyZomJ0SuJnI3Iw+Pyr4d+HXl5DZ+HkNowdxifuDdY1VebAldmE9O3qUt3w
u6M8lYyvgP7dyo9ZX9KjCmz/SRlF/6GUhcLNfy90BZTa3OK3nezo/XwyuPmvdnO9
FvP+sR96H/MUbiYHRUGyeLqSzRSRuUV/W0n6bdMB2Y6bqjAsg9skui5t/xFGOgjt
OoEaFi162O1tyR3YKbVrJb8f32XiWCJg7GMJMYV5Ss0844Ij50JKjGpjPfiJl2XK
zZtFbmZjdqRIgaa93ZawiMsCxwMKl4e8jm/dt0vru1kDYihHReFX8RjL0sOZVXXw
NLKrgKUHUJ5bn58+/4YsAezBE86huyg6xH74bL0ugOW9NDo1bRL0ZdfSYJvdQBz2
Azx8Rhv90VdNGFhDNKOuL5Tdpe7t0nXnTtrmWHzgsaBaURqRqQEUlQ+dBE/HOj7m
uIKKs89Pov6gK2/ABaMO75mjhJEg5VkqUmXONoEV6stw5NZdc4ZNRL8ClRMDsn3B
71WeyAVtHS4DNqvF3IkFkuTbvgZXwOh5vF6rpyffYO/MYsDRdTTHgvOcVnXIFaXP
qbblGV0xWMIgdsSaRa+PrmMHMvqMDAs+KGhgeWWnIyyRf8M80heC2IbHw1fq8Pc1
JO2b6PVV+ftGcdUKad5L76iMFA6p3CKVPr+gBBv60s9g8GBkpOaQw5wX1PJwq+x3
Xfyw0JViR0VqD1KEWAk15dzHNqB9b+V5ii3Ttyn732mmg6vdyXqTeJxCbit+TDRr
gzrKGFxC0a1OWQxoVucNC8pYafVy57Gtn3DW5ZAnS95udMZw755NF2ejJPmGv4iS
mxCqj5NBRRdATjRyYiuR/zADX8wMFamciNbKILmiZRyGgmtzMcCFv6fbcsulsdT5
9zMTZcbUl1Ucbr/17GoNQkS/UkrmCkf7LUuaXkAWPvCvQ1bnxaimG1AAe1SOp/yp
pfRl5jPpU0L/x6Rl2V9rrUskiAvYEsQrH0z/DZ7g5C4R8L15wSukN9fKpmMGK7V3
oCodM/nQIRVdx6JOD3VxBFz+FbFLgTc31SPtfmHfs6/qjDZxvSuouqe21ePTlep/
+BOT26MrS4BzOpA/xmHi3DVKhUTkliClhZBfaiWW80a8Zx+om/Eno25B1hz8IgrI
I+B2wBnnRrbU1vnxXB6+sJcNTMgwxfGEHYEHrNJouglsfoARbzi6i70btozLKb20
AAh4Z8E6FpA0+CCLh4iUCSU1uyIjvOiCqD+PLbOgXV5gsX95hu5KlW3+LVTmDuwn
/ziXS27Pnp9cRfojkOwCzgH3XpkMU/YAMCP2lFA+CpNOJRQ+Zp9tjqsQCVth8dJH
2Ib4zDdzAgEU88NUw7i8BSyJv8Fyd4g4BQ8qQiGlpnf/z9yQD0fDzxNO1m9ZFHND
moTMmarCYDyB2et47wS+tYJZtUVnPcsxpDo258OHP02lpxhCaXLV/iWnENgEQm16
maNJ8rRSfyywh5/aOmJSQxUTmm95mbTFtDJLRApyxMyPYE4Efxc+oC7FelFqpW6+
BMgeHJG0m2QdgL55dscOE3aGBHX6chMqo+AwxJN5AlZPgt9rhNNQ9lD8rpkx0D5w
IY+HQYMWx3k2lxGAwA0WDfk7G9T24jWyxgQHNY0TAK8ttGnCiiXmC9Pb3UOYQiUO
86/C85Ytu48L/hbfSYm4il/hxPM2o8dfQbFAbtxIQMqQQiE9Q5r69l9uoAPgjDfO
kYt49q03uxUJFean/7k9edBU9G1FnLc5TbBaYY3ca1tZHY/vBzZ0acaVe6Qr77uG
87URti83+1zoq7hzX7sZnUcHYdwW3tT1CaSbxgNft9NHtIez7rR5ZnvKDMFctY8s
ITg6wFAL0wqVAUWFsLeAy5dtmLMM+dYR1ADk8eKIFsCzSyzacl3GXlS8dkK/vq1z
qmNRGYlpdxy30ozNy7najUlD/+4CLoGdv9+Oa1/iOdDIAU5/AHNitj8SdffsZ+4Z
jNt4+6lIjCCAjaPeZBZvFbi+mh6CkohAoox3IVhdmcI1nkDTcyhA/ofz6HHWhPS8
+epmUppijrGFlJIBQc9S+foBoTFyaVJlVvxI2ynMyp8Or7n9FwRWTMmx71nPvINH
M6Rpr5t3BtRVt9tm9i7u4yv21JPXnan1ALt8mFK8qlfKXk3r0j74SYnDaTqdv5mx
pmcpv7/tJWLkPud7mDbJ91SAKg55pVqrDbRrX9MWJj+ku9Vc3Y+uSivEVZJuWodo
Wia0BCJy/3erFIoFJpkgOpmbMt/uCxO8NvSuG2gaYdtpoMzanX+HwZfhedUaZLm6
M3cIh1Vcd03/cdwENyKVTIpNoiHmOh57IrTvcQGbH8vdia64haIpbPn2wFmq2f1z
MHc4DFuJJkStuh3IsjeZWUA7IVmBnKZKSpLRELaVITjO2ro1lvtgjApbFfNclPCY
NRLMkOe53cBMWgpI1XQVPDhl/NOtMNX/buidQco6NjnQoNig5Oah2QfUuyFN/GHz
ZaGq15s9arM9E8hfBZ8+Pu62mtd7/AjwLqIWvd9A0F0Fkj1cDAHjqrpm97JgdQ5Y
Gnj/PVVg4E/Y9ud4Z3Cyn/LC/Q+r2KmzOFODtpYgIToNBjqzLqOWgwgez+c5jAHl
jghj0VtfJjqWy3TxaHX0m3tz9LGLO/Ly9ETFTsd+aAf79yIW9z1K4mYNIsVjDhq0
Ld0IBmed2pSchBhf1HWXoKkds4efff3POLIRyTETk+7v6MhV6LPINLV98MPRYKXm
etkUSOj42/FlcYv/yKNirpO+C7LWXwGyKwISldzEgDr4nUooU386VWya6GFEw2L7
+Ur/3EW2M7MxQVn2/Sv3CnP9IgR6ubOb7/buDqX7RH+2kSucsUT2h4Pqj1yBWeTz
6TKsrSD+B+JcXUJxLNWGG9s+94W/BU1111cUjMO7V5WtemoplQA03zQFHet9kBiz
TfdJ06T9hV/yJIYrEldpZ8I73ZlLSQ13G7d2r1BLFD9Pv8Wr6+MZmhlmFeUwf9eH
Xx5NSGtyzpW7X9DlVcGIdHPQd5Pn2TDKvsNiUDH73JtaFR7ea5k7VvF+5ce6q0GO
zQI3ULJgmZimKrXzt0PykQUrH5FaKUdo0dMazpnr437HR6ewN11yOcaoUtdfR+p+
sP5p+WrRjouCEhHDG+JywweH/GemkTeF3wlS0ktNdsCDfG90SHzRtd0lyYpzXMYL
PKkJoehUYLv3kk3rQASkmiO/ULiBYchssoj4JlUJCl2UPOyy2MefA7nRoePQAJf3
Uj+VMvjtT5XkuWG6T+vZEUc9DpViq8TGvqtbSD3CCzv2C4G1RW0LpcL1+P/Yuqzv
n2pvaJKYl6vlFoMTwCVmlluRYNNSSddln9gcHCtjyGUuY0zAno8+jTGourvi9mrc
aV7clE+gEHOg77ToNs4YENP7ySKE2PiM9qL/5RnjueTSMEfgg7hGVvswx1d4vg39
nUys8tyddp4DcNPwzaQhGDQioJu8e9YZigch6Q7GCDgJbobS6wukO4+0XuYEoNKU
ttLgAcU8r2Qn/v4VDn+cd6uNkX5IcKMeBbtXi+S4vq8iw6wytDvaQoO05RKJhGpt
EsWHtMM7221Fmn9+sDaqWvJmsFb4XLeKHZbWgAOJOzLOpVvEgi+Bx9NdhaxuBLUw
FJLMVRppfOcmkmulIUVroDcwZ5vw8YfzlI6QYpTqGFIxjbT18d7VOYwtw/O3rWHL
h9lLrBI+B2qyBtkRimUZORYuB5YnSMOgf2cfXYLF7HZ6vrKx6SGiQPDP4D4we9vd
0c7yAnhLzcMnKgoBsbMt42IhrzhDv8SB/kh7Ln7/LuntTl8gDTTnrJ87Oybay93L
50Zz1IST8MgJ8GPp3liAh6Lgqo4WZOU5YHuzay2A3Ogs6dHR2T0SGk78JrpRrbB+
cCxNQDMdTwMcXUfpDK5glzdTGhwHN8CtWhafYKkJcW2wQyiV6y/TeJh80kFWlLXI
tAqNYDnxG3PSxxCQ9dNh0zC1nt8x8eeXz8S5ThPhq0XmitN1frWwDLyEd0MSbOTn
49DjJHNGwSd92GDqbadHvv4z0N7CIBiI9X1PRC+MNvcJByAEYc1hFYirqokxsQEt
oQzyf1wkl94UEl8yH+UjchClnsQzX1Be/Ynu7zbPnssA4mh+2NKKG+E7pW6vW8NB
Wkh0xHyIUQ7SjvGIMeQcYlgc1Lx3fTzpfiO6XJ6NZB9a6gOfPCJ7EqZDmeS6kAeW
xaVWyl4plLctis0zrgWwwVVfhxDTF4siWOWJ7cbNvIfqS87wBneySY2bZyM5vTwo
NJqsTqY1elEXSD+P2TrPfZSzQCnpTOfz3PqrDa9/FkvkdgXidOorU3JB82i7ybyj
ggIJQEY46fLoXqdjtnMQxlxnO8tFqxGjvTryeESRMavE0NyX/+c533AQYlTq81bU
p3YseIRGwFTSrtk4ttOUCwu6h7YLqTJK4LwH3TxYStuxUbzdFJzLPa08NBAvub7w
IT62zXNZf8yWNM9EuEW0miKI+HTTtsidL4ZTeGLhpSiwDZj4B3uvIzw+bPVI/EVl
aD2JaYcrH230iJVnEwNPCo4LjuxDuKq+kH5rv1YmbGY4m1Nwc0pQYl0n46u4Nt+e
49e3iDgRPvDGKnYIKY+UNZpysVwu/hkjQOm/YvxSS+vOlRCLxAaUqiHdAHzx8Iva
OD6pCYolGgM0lSIm8+7sfFTuAtmMg2fHQUAj/03jud7LmXzS+1Y8q1E9bK+t6mgC
tCr87gIIQzSSwn5rxIYWLujGT1NwniUx1tm+nUzNlboeL8gKtXThFPc4B9tubHpR
m1vtDsXD264+8E7WBhkCHrO3ZAUUe2T5Y7fPKi9P/7gQTmGs4QtO67wYSz6wRY3Y
Wcc/gUZE4HLHEh91qfEVlD8nUYZDnuBmm3caHudS3xtVCMFhtBNeq3dp2wcDKb3f
Jc7j4yFq0myUuacGyMnnPPi23fNuahB7NiPF1/ZguU9EfhLtRHrXlLVhp5gV4vIJ
L9/HQETGcx+7yY0/tB4a+RnbhYcT3GrgRWbJFWhgdm2Yxpn40rGHb/VbGlmATh0b
HlV81vbk7/Qc9DpZ+QO1aSdJUfhtr7nauk4jBhf4pZY5D3u9LzSVhrYYlkPnHvoa
UH6Lc/o7Sbgl3wGk2xY396X0H47VRRHwZzzXEcPOxwO6nmYGv40rEgSBa/3GMDEb
tf5L0bkSW9BON53P6vHejAaPEmB5ZzBQHM3AoN194On6Q5XdssJY/PZEcOihexU6
7OOXmOruIBi12DvwWDJp00srQK5yOhsNCQqklF9BLjOxXCdTTvQGflPedFv4X9B7
6T9h7ntcbVcBaYJQXchA2eBSVGQmjFRaDfNLcVPGy4YJfy6qjAKcDRcArG3w1TNP
I582PUtO8nvzWsq70a//9GxYehuUGLeey6kVPcreKJuaHJOj4mqLUbfpeix7Yd/f
S9g5sBrylE34jiIrGOK68ZuV+DFOdv7+kZ4+YZIwjy8URl+mFHj90w3z48mwHIY+
XIW1o0/ife4YdzLMZulD8GS0SYiA4QaFGpIDf3Sm4JNt8rVrKxggYdGYbKx+CCPv
me0HXKAaqmYa99uayaYEuKIdbxDXeMdgpO+XcKahAcvPDjoLhPF9+CArLtbGCfEV
ScCVNQ4Nc//rrwm27T3TKGGcxM8AA+htX8p3WLL1wsrt2vA3CkBLXRKWEvbwy3kX
JbbUjbZRAGdQ+a9EZbtHSI1R9w8D5pm2I2TjOyil9VrmcD7vHehxjdmQaqZpiOh9
gZwecSaz88dySulBHAEuCzYj6SetsbmVzhP85HopvmxXig6u64W6OzC4zP29ygLq
AnbBqi5npZi9DKvIuRFEU1ZcvakYvzbAysfcq51VmqpS2Wq+gOWy0ric0UdklzNk
1gC37/Np+HdLLnPg5qAGmcEladCR4PNlP598hrG3D/eLfJW6PiKvK5o9qzqIgHda
CZlIIdWBOku1i1Ng8cBAsjFFZZeWZaWnD2UBdQo2kBJrPAbxaxiqjiiMzmepA3z/
AGorYN7eedO7EeltfKmoTcVihecZHQPSgiIUw0Y0MRH21mWrHj9SpvvNy7nKmcPE
QJ4Ev4YVCrmAGxp1n2OcTUTKpjVLPOnguXiYuAI84UnClu3lDxcgbGAz9ICczv2f
wrF8Nsm1p3ovgmQxKjxRMuwaM7Cmoj1x53kqE81IZ25LT3gzZBY4f2jmccJVF7cx
eBmh3V7C6tiNuM+lShMBirqldVD9DBQ4pxPzkgokqzrRFKkNvI+djLBhNJY5zn4Q
JzcjX6DeK86dqjiF2Mbar5VVPMB8867JQ0wwmDUlnyu0C2a5A0A+r7P1c77N4ruH
wYwLvCMsRzD3jFxS+LYIuNucq28zXWpTfeYPt0yu+UDJliRg2++l6OcQstA1ourq
Q613/j4HEScb9dxRsnTh1pj5u7PrrpnKc+xriy3qEvru6Zl2g+yZxHosJq3F7jVw
vg+zcFuA4nICBRMjQyVzkkZWh4uWXk5pKZQPbNt2AfYug8ih+CMiCIy+9QoNAs9M
Qgfo/AkebncUVChDjNath4E+x0zG+UOd7MDh/fBTnNAYp6elHGlUQvvjSC909olI
gfZy0fm82/v5GuWBJdgPTFkYln8EaWS1rsdpJpaJ6yPTVuPkW+Yw4XB747ycd/ZP
JSzPq2gZU6IO6rpjwDxPxTTzaZVffA48uoFizDMXyLAqBEbgHOYjpdZDQYI2J4pl
GUTUBN+AW9noXmpHJfN24iq3XHqsO3NiNRCa0xMSmG98GNZYl/1X8zuioGHOVkdW
pZ72ZrDi6FnAKmWtOtIC0jsEW9U0JcazQVqxZ3iFnhewOy1FfK0Cuecn7JH+BuRd
DfaKAEzEi8103+BwjXEgCH6HKb9OkzlIueSYC1wpFA+6POz4XTngF67WYsp3lomQ
2hJDNEBu5FmGkw/vJ2AUsB96ouUzDLSovD5SuFQzFOMma4CyztH4SqPLmkNNg57S
JN7iA2J0u3Jphw9t2jB8ZqKvhJ1alAoR7GWM7aaNU7mNbLO4K/oZZEOm6iB7XgC+
M5Y5O1Y1M4JAXf+BRXQ14WVyx9qcThYz7763F4xNtQm44tJ6xrXdomJQBbaPzL6P
r8eViViOlZOCjkMNNEp4K2TFd6bR39OQ2kaw2YjlAHXIM9m3/oEI1aMbkOnT3bNN
5nl9W8DPOiM7WETaVEZ3ImU8d45c7leUHhCmz+TwGC0Yd3ryu7mygPuEEiQ+u0/z
02TgJJLYiQubzx/gSF1Ti++9InX63Rz6+ngErxbGZTBsiZvEt6bPZq9Pdlowk+CU
APM80PsfB76rP7XIXGA8PEdoCkYOUIgySEZu85HifXXK/1RhWiWJJEKwMQaDczuf
NU1kFiKZtCUlsT148cwheB17lIbu8svRHtFqCybBlb+Kr4QEZu+ehmrRw8YazEqk
XNLracq5cq5+mOg912U47lSkro67QL23GUIcYPNL+iWds9SdxWNreLPjI5N7B+QX
bmdxD7grxKbP5N65DkNOatoHzvky+yvZvfosDjYiYbRkKVi+eXIwZi+WcSaVBCyB
3kIH5fo2k+zp/gdO37OPcBnN6IZH4v9ZtzZ+ikvbzXalSkeBAiPSuxJ/dNarorTg
qPU0r3Dj1SSYmEbFiXhoXP7k7P8arZ6+gAjWZeuGvh2/l532BtZfp07VlTSnRiip
+ngTJzJ3z1J/E0SMnSjltRJnVRgOImhm34yfm8qTtJcg/oDSklv8dzm90wXJX7dk
zM1Jc+yy7Q8GeFX5C8vG+PwEpm6XAviXU7R+noOANZo4y2wKuVNceCLUPFk2GzDA
PdmcgLJkV49DKyqpalPZ1aJNXER7gaTC4/qyJqsbzmyuA+45i0GPfKSRzQ3+7X4y
LXcCPw3Bw0wAv95eyTGLsb+0s9PFEJnkJFC3okdPwGpfWws7la2oiXbTkLOacsn6
Ge4tGjRKpKiOGL4x3c81H+EOVuK3pVdMaBAxxfYTv4yy8mWJ5NLs8fxjyQfYvrY/
ncasmXjBQ8jHGU2I9ZnRzuhhAd2OnqLHPgS+2T+PIRgLYsnFNwMWG5G751Q+U4xG
2og2N2Suot33E77dIIiHbGJO3SV/8q2EkXU/xBtpzMNhaKnAldAZqW11m5JMuIZD
QHdjjicgps1FTgSv6hQphbsB2TVopVcywcWIYQLxdRmMQu/DntAdMF0l6AswN2Sm
xPC5Sqxx9/IZd7J6vFbmN77uBUQZhOzlkREr4xkWH1d0TAkDpifJbzblQ+6yLLOs
HINokpIBhUXNvzQ16ytId0rAUcuYksuCZFDG6RKr52JCyq68gBBY49Jmfq6So8JJ
+9+AtzUG+wR+MVesfnz7Ozpp2jSlsh2F0OnJsGssaaGncDZf2vl/OjSRcQGt/8bZ
4kYEPRvKEX0ekG3Y3McIO7PBEeMwyF9f4NmvZZ7BO4XjKQb1N/BO4dfnwCkFwfbq
4SAMA9QODCGnaYktfzBU0bQEGEHvIi/hO9g4A7xChEEHpVt6UNQSQQkqJsy5JGB8
gPmxO/kKLkzPJRAIsCqXGeYbdoRahYlPo2H/JEK9thTVSGjCTnNC+SPF8XXTD+MB
Ut+Uh5tlLaeoF4jC8e2hzcRSdDUn3dm6ZOlY/FiMmPlP5NgCmhluMWcX96m6qUW8
RJClF63p+0JDpOlUFeJyVWG6X1Sw2px/U0WFPuUBnuQN5o4FLk3yXxjVTjp6XyZ8
SIsZbe77fQ5ZkAwACm8IV9JwbYCxV4nFvMLK4WYoDO/2yhLtnNakc6nH30UqQhhC
1EzcrNPulC3YxHwjNccwYHm47sKks3n9mamacXLuZKRixMmFMt9h27VfvJmZZ0ET
8brt+ERmbr3ydThXCUgO5kqYdSFjLztlGIfuba2xJIk406JvDqMmEZnkaY+MvCju
6oh9kZMfbMbQz393w3RWGnWII288yFjnawhIz9dl5yE2px1+vnXejTlTVSaGl+VU
JTht0VcsaMQcFAfW6+m0QYFum0kXmu2R13bXQerd/knZFbaUJ4vb5Gmn6FhKuzfD
xJokfEq/W6XOz4GIUETc3ffDYopWC9Zxv+xhk8WuZt8DHngwo66AVYRugcnq76nr
hmvMfSZQG6AzZwqrFEraBKh7l5XAAymWWDcas/R21pA9hlAk68QBziQ2eElCrbsW
1xzIxwfqC/TNPtCD1ggRtI1pLNP+cHuQ47fB3J11tXGHWDvv9jbao2JlClwFp6W2
tBACUIcPt3N2oEdNVNh7vPWRIuDZsOsCivMAiPr2BfzPDfuiLUxuGfz1zA4weNlI
Q5SNvd53TBeSjvf3V+vVFlwOTpiMvuoGCRj5Wh5g8XIvIN0V7BDzp61yDkjIfAM6
pJcKpGt9Tm92ZVvGxbA4Mq23V4nw2DJNRzH7N8fPZ5Pq6T8OtfOFKU6hcYNhRhB9
v+TWJcPYwa+RJSek0IVHN+rT3yYwPky/Kz3tLAlULG15Te3Kkbgxh6U41TFQmR+S
Bd8QlGdJWnh8h7AaZx5b0VRhmQkY67PrxhcD0VYV3svr5CuhN8hBD28cs1chOoNw
sW5A3EdR0Ek76e0EEDWTRx+qdWwx7waMoln+prr4Pol4Rvu6SIndBujHDrQIDBVr
hW6dHZfpwp99mDfPMwaaY1EnnxuzoEFKBHKQBZwf+yh4jbUIwXMnLGBdT1gYONN7
JEGtg1+9FZWXoAD4YFwZ2G2/Fezkl7BVQv/tf7izpR1nblwYWcospQb+j/jxhrpL
NdPSaiOSkDXCRtp1K/Pu3TGhU4hoLCoAwlnutRdW58fd1YtGQFhwo+UVOf5hNMT0
7LTSw5VhwIWKNwBdlXWOBTpRCHqKNIm6cf6f9pf7JeUczFne69qRc60tt62/kh/m
gbUK/hlTAw6kajvdFqC8NgPCmDcRNmZjXrLfUQ6vrqoUfUXcuUZNfBwDoSbViq1i
aAlG6Q+BScceuNxAxTa+x2rJlBqgncNUUxoQwE2f2JiELjKEUdd8TTgoxD7nW7+8
tg4YW43wd/YPkfmETgNGajAdPzpidLfaWbhnRH7xwN/shtNdwkeCdHaMJF0TW8DX
rvEYg0SCtmcDx2IFZbFaGHfXGPhObrSx2QCwiVcU4MQ2WnnOGNU63/cfl+gBeDLs
Nb+1FC2KjRHyO7AwhGQ8/jq76n1NmgOD+O/cG85NGw6sRm6cyK6L4j5vtHs8M0lO
FXjk8+0velSC7b8TkLO0IguVvvYNbNRtKeH537XKHEmoljugTFMf8rdz+FAyORYT
En3yqFVy7GKLFE+oY9C48Tdv2f0ELmrmgDhhOGudo+nrRvvcYEWp4Dea7uUtZRNQ
0yJv5UXj2dKkW7B5mzXX3VcauB9Eyks5B6LDNmNWs6mixmCqszbohr6cyTqXa97l
SdvCwNj8UMgl8pJZ5wc0no1EzB//71tlywJQP6ryjEuNrcI8F1iqhef0bE+0IjAM
hsFevyWRMdR0z2SsRLFYWXiGS3t2dEpYDmyp6ZFjRogJmPfBWWYHQkaYw+oHpfiw
wyad3H2Dz/mV+K742ZDXK99GJRjDCxB1S39gXPdUXUDuKO1KdVEHy/uxBrUp0KmA
JA/LFXbx6XCWDvGTHBq/JhiIWVP3ax3H318S8YH8Gl5K/pxOO3k54WB2KJUNMtOb
afTOlC2EuiigdcxS++mI9twDBn0zDjPiYpt3jLK8LdhlO+rE5dP+bJKw98pryIRx
SE+/A4EdMAKESVlq0ALQP3rNVnyS/mn3ojbe4fV1Db2tfIyAdYcQ5ZMXSyPDbQw/
JnvdTuZXvUUT0pf2LfKPKeIwkHT2vpJHKD5xwxGhT9or0iCclZMCuBcjhAMZKiAx
nbLz93R40/TOC47OmYstTrw4rW2tpf34zOfZrXFzo0gyJOhIaRPaN48GAlqZAu7p
Urj6fwBS4AOnzoSqje5iFxUmyjZAK3FfJHSx17xpPdWsb4Rcmmi/DbKzyPahXTVg
9OBdtlGVeRIwAiSB/kFK8iJ7bSVc9IiNp/gnBkp6PyQ/XIU7TW4VzcNAFOIVKwWq
YDVeP6TVrmBhfEIFaGkKnMR30e8dVE1yJG7puZSjX630lYC+X66QxO9XEELujURD
2yB22C/qcKSMmVye3J/cuxcJMUTuExc2O3o/dtjCgTuYDXYwCqcgevcq15qtFwEq
FkJdtNMi7mVYIEy9IN0hkpXnDgx6oRiRg9MTjb4JsOdX/LTicBbq/XnKAHnhOhyi
hZ97rumKQjAPJ9SGaSl7BO/QxBOUdBzZ9y1b/rK5xIvNnDPopdrezMntFsoITCoP
FvUXwWi9Jf8EW5EcmSrRO60cvdaArZOpDHCL2yWP31XEl3PXYG5jDmwn7X8KnJko
23Qc6+S2qqQrU3OJZqNzn1HmEoH943VDJ1jrw7171/QGdstrHly1Ijuga8UbtBU9
UNYj5F9rn2xoPrdi61vhocrQ6PTXhJmRj44NscrIPD7Qwl7irEjy4v7b+Daid5Xq
/7lNYEeOvthrrTskq0nNy/Nlr2IgLbe7RtPu0Ej1bR5t5t4iAXTbJYIWAoHt4t56
Rsa4s6vD8zGzkl+SXYtRFD0Am7k13S9R7uCDHhMosWcI9AIqR1X4DDGD6nD4mhMs
Df5y45bbd3/o1ndIiaV0JooykBpnZKjRm9YNVjrC7jMo9en9gaacY3JhujfvT3Up
oaDFOen5VN7gR/WBtn5bNEYjcilSLcTebVvI1kQ0UerDqj4hm0xSr1dWhyAfoH1m
Cxcuqw43W3x/WJyMDCNutUKebO/6Kjg/CP6dAxTwLb9hzUTcnB4fvHQF3zkK+Ktr
kqrt0ZM8wbN2HSzrq8LATkb6+AD5pEF31cjQhIzMAe55Sfw9xHVY2P7sIOcUsY79
eb7My5F8KU3buttAdG9P2pEpBW40v8SNnSejozT6tCYk9LbUE+61dRWJ+kfpLnxZ
7Hj3NiMUV1i6LabeTehxtYOT+5nSgJhXqYMPYYO/qJnc3Ubw2EIo3drtJDCHmUZ3
WyekCsHZY8V+EXlSsqrThAC1kF1v0Bp1HlTEUcCUx/xm/x0t4ljZTfEV42srEt2o
pkT6Hz5nGmALIZgMtzhcTmtgLIr9iPlZtuXo2eeOTvuGWK4B7Plb35FkFtGEBnDT
gFP9E0wF2lyIAeGlt2MuTi70i3CNDcVoUQ8Wx26NbImkcOysYoYTUdcAOUjGtZPY
okGxaXbf1DyeCplfZx9mctvAeBD+snrirCH8w9MNfQNEpklBXCDJGP3pCzjqjXbn
G9ABnRCrZ6P0dVQsyQOccKSCkAtLnbpqrqpUYpH4pTD8TtHL0+BoCDnXwdN7xeUT
3a3guJbPfmF5pBt/ndqAaKgTyxJNrocmn2W36acneWmTkFrx6aQj9hW1bcd9koAx
5tNrX+Um7eLyAb/JPnze44qFofDPLjw+l06GK1flwculSDKU1I7pUJXZCLY8+XSh
uGsFP6AM4Mf/nV2/5JyGrPjvLrL/c4TkaBQKqd2Lui1zJkGlAR+vQfl2g700q5Sb
vxAVIWd6DFRnMrCfnfrVNxCaxtpPzWc5YiB0NReHGSY3P9BrYsUIqVOsSzU5sVfM
Y5tS4fV3A7wkYO4Ccpixt7Rf6L2PsyO55QsYLtIrM3xvs6aXITF7aBx39dedNzm/
0pdFNy8NETITi+GvfiZ+/ZMilBg1FnIjuZu0ylXrv3jHmRkt/prkPlXhrSer89H6
pjF2zw9Rb5NN1IFOEwlf7BkBiwR1fbsm4fdxXIWrJdyglBu6Sq4EkEpfL1Wnph5P
slioYh9MFYin3kWb09WTp2QEckuK7C//WytpwPgUBH4nKDFymhGL3mR67BfvkrGb
UxYcK/2Flxa04lvcQPOc07JO/70reNYsrRx/hl6EvtXhUOWRlef8bV1/oF9rSSMH
FWbIHWdTOHfNeNhBQv/Tj21pKxhJ39ln9vUOCJRaoA9zWuLczr9YEk/UD6Q40/4y
8OXaC4TzBmhd96ZsixOKUVHlAPPc4FJZgs26eP1f18lo1SbKFonoFfuUBp8I6PiO
H0tPOw1R1ogAQOYngzfQHKLtgN2g6cGsYuB2PGr96kN0QQY/s3po6z98BBTkhyMI
oBqoNe1l3bU/adi2zgNkOv+FEqnt9dwaS/YH6nNDexTv2Uw+XunUvlTx4AcQ7//D
Z4QMCOoitNaYoAs9bUkdrLnoGsdLbSPfp5vVzBeM0G9PiJPNJW4iV7u51M8KBgMF
u5IIweVYmb+XW7E80nuLODQvhy1psu8Y4TdeCsumAYbXCALAgxJNgRqzdSP3YGYz
l4ZAjhAmsLwrkJMZ+B81EbTFObN/YOFGqDwLiajHay96yr+T4j67bHSy4DkDnGNA
9PvR0OFTRsFtHiWCwJvrmo+t2ssjTSJBO/KiwuEDsMBx1Qk9kRLIlLKn664izyMO
kC5PSzHMGHcrPXNR/FvXU5ejH0J7gtpQKd9rU0HEitOu0AW65AL+EwkZtuW4N/PI
6dXigrBnQrdvvVDG8xwImpQeGAXWpDRaubHkUndpEi7P7fmllihltNuZPAQ90Vdk
p08dSZz92ZadQ1ne+hP2zZuoXuWm9vFcElGuaPvFE43FpHeIYbkrEN0T1+WufbFR
fBfZtLD8FMWztzcxGcGRrmEc9ju7xfJ7vZXcoVfDYAEOeHh2G3md4tldGn05wqnq
R2BNErvaIm5xAz3x9noIt9m2TDUtxLfJlYbstO7YowPJtTHtE2kSd8wGYVjOFTCh
It/xt93g1DemhU8lN2pnBWs8ISd8bfbcPYMGEJ5OZukiEJk3rIDhN48Tw+0PITtQ
hKTN61nI5kksPPJoxIdI1ZartBBzc0xZ/f3b0VMdQW8k7AKJvo9KJr5L8sx9sX1u
mwE17k6Ou8k7sa4PBle5HzCXusFYLuWG6gunwUV0ten3kzz66mRlqkRI5U2T9MOO
+elfHb+AoHR0NJD/DtOXXvWM0yyCmaDHa6XWqgJuWtrNUd1/Fii8iXPPv/eJ4m3x
RkqO+Ul6Od6/+yePM4bmtVj9WTEl5SCrRi1q4+uAYOAMFidGXZ7rqZQMjlT30kUf
vBRN+yojITkImdrm6B6IC8KwEaylZgf1RKfAxQd8w0b4xbvdkqLJygQUkta49PHK
hzHX2qQDucLKnqB1lKOBGEfQr9P7D/VbDMGCTo2ffNmdytiXaJx05mpjF/IOd4UI
dQGKUaiTwWDsl0BhPQIx3/TGo/S23Vif/wrb3ihtkp6TFSGT83SfHoF2B85K/rzD
+OXvsjPcqXsNXAYjKmou3lr359PY+Hj2DUM8B/WS+IZR4s70tVgypJGYbrzRSblZ
tXubGdqL5X0oN6euxj9TXYFQozxe9bSMMoo5J3nuImo9/k+7fYvm+owfa9twXyVX
YM7RmDHZcDtTbvmv0aK8uFezwcnX8V3ijCQN/bMzMal0IlfU2JQnR5B2fR7Ede00
xTPxcY9gnRNc2CcimtPqmbMxO+XgOSUDG0+5RHf7ohcX1SboS/Z6gDM6InOoCtYR
fBGk+S+rMRVND6upLr8dDwGreBUlNXwG9z5dyDrcN9/fkHA6i9leWdWegthISPoO
ftvdenAbjNUbxNvjbvUWj5S/KR10BKSieZn8bss49N6uMJKhlr6m7KWrtPqIJ2Js
AsMM4MY4dKuaGzEwludovQdVe5iH/qCO04Mo2ciPDQxwIPRMB0vqAnQggyNThln4
UyqG5NCBjEeIgERkFlU63ChmogAHAAbkUyDY+2Jg0Z7s0XOLvghYbL3N79DUpAva
dxdWCpZMOhmJ7yfe9wkuew4wCXEyd7UsKnRWtl6CpE5ykgdm6UFZ0q4io3v8pVZi
xPz+/Cdm3TmYPHPfEU7gsKaKPj9B+aEYACOEju8erDWw9aE/sV9VVy7OFc+Ph25S
NmwePskOUs9zJWAjg/oFhOrLr6QeOUxR1IOiq+btxV41TaFomBnUKxVwlZAj/S8j
XH69MfzFGdkgaC0rcicg3lnQksQa+g3JD6vH31jEXV6gDSmzeJ0JfGjYgmZbo0Y9
9M04F09SQ2S4ZdN13wDxC2YFnDdXyyI47Gl1KeRtEHP3s5Z/oiRHE0CxUGAsxo9a
sJspUIT5ql5g8av4CBh5Kb9VMYDF9DdO7f1biIG84MdIzZCmfje33v446bcOXK9Q
qKbuDfaaQnVxKeASzqbdd72tazIL1dHa3q+mZPqNOOjw2AvnT/9esFMyamxeX05N
7Rb1VUwHvBrybKlFi01tt4ZGQGFYie8TkKus8/XXfo8VJK65MQ/zpZv+jHAFr7O9
q0uRrWdSWoeCXS3JDnfmdQ+op1D3bOPtBnWwgh6qM8hY52eaXuxgHS0w0RXK+MTI
/btHLM8GIZ5oP6QbN/4+WEgVfAkutqJ4XvyWdsQi83fGJcAdojKfOWCZ5tLMFnVA
LTlNeKMN8n666co4O6dfPFDFtrzaDlkMtCS2aOZ9Q7BkpnygikRoMJuXaV6NE3hW
HnKk5zYzpmFbBrQz2NUM/hx9L1MABf0IhlXQ3vks181hCFpmaiD2Jk1rHuL6kDP0
G18j19oPZJ94W2wTkmq9T8tD5+TX1V+ixTYK/dLggSQTZa5BDOFmXmCYzemZJvVV
i8dESp+/CCvrf9utQTG4ROL2w+fxM1Zz7GOcwtxrYpisTbNLIlROjgQfTUIGs+wo
s44Qv0PerjsCi5h6lIw/ZFZrmtso5hEcM4bM7wWY0uaurQOMPZK8wVyRvhDKzBwB
PuPOEZUuPqxaLbOH1yqbxINnP6kr3jsJDMZtkKxMWEv7SpkRTsZOQaWb8isZU29W
Y/EVLKBi/2ynUvIvdnfUzIq9rTDlbhWRi8UfMQvFFjX6iViQWbyVd3NzyNAsvRgS
YarTXsnNPJTrRgRXkZrYAlU0KL3aQsS1vYYmrS+gVSDykzY13X7HTfkyXDa1QOx5
Hk8HWOyXEMBOFTC6tFwDqOuLRqM3YlQF0GvSbDSGIW9AnPfO4ZSo5FD7uI+tZ/6A
4QEtRn0n4kOJoPueh/Av9zdNfafokmCwAYnzg6+k5ZCfIZD0OXRI8vPfaezmSZ+G
Hxm4VSYaBDeWP97vwwWjl/wcItEQn+SUN7aDhbNeCbuN5vg2E33qh4c7DFC5uPlH
g8nL/psHBleXEtwYzH6TXH4GVD6nJgiKcZIaY9l5BRSUveHGbxabYWy1fq+29k7S
GuV1EacgdbgN/assynx2KDXxMv1kxvKR4sEK2gpvdFhgAJUrCCkhAWw3VnWqyqAU
6b1iyEiVSj2bmHB6qlXU4rJ9cGytMh3j3plaFJduaCp5eR/VorXQkxRzTfTGSFx8
uPx+Wm4jH1pxvgTWiHio0Wka0RXxttFkToeIFX1YIumyIpwT7t1MT4IfOgTh010i
d7AZ+4SHfgW5cjxDKsF8uAOmFzUkkz9fqDpzVnAFhj+bYIY2wv1ckzZZEk3PeuKO
m7aPBDEhMGOOiJWAjPvXraZN+22GZH86sNs3CvYfFih9KJSMbFk2JCaNGXBI0W9D
9r+XtX4xXc6iiYk1GNLWDLD7vbqfU7QEZYm6nKVeFU3LG2RGObEVP9F6b9ZEBE8m
N8M6uRlJSVlIVFkUVEXQFhStrMjXT+S6Kc6fpkh1SVRJqRnLauq0bnfX5w0axD2H
t54v9xclEJLVQ1ealsYJEnAc1tznvTWtyc72vskpeUIOIniw81RdpUydnA+22vkb
Lh0E21wqDrBg7dKUhQYkJgwPd6zRFKth5GHOUf769KDHhfX/oLnxnZYL1ImzdDIf
ynDHS5wUJm0i5oCWY2ZVaOsQZ6a9ShSwSVI2rU6j4FnQJ8cNbIHUuS1+fOp+fgbY
h6MAN0i7GAnFhKK1JAHnaZuZQcevhLXR7cnZxQp0hpVZZP2eEQT5z5C6OEJGh5LH
d0tz/JT2CkmaIFpdHn6xr6hOtZT6on4NMUCsdZUyEmspWMSNXxYj3h19JcH/JHCy
Txb7j1JTr+X5R7nOgxpCiQEZFlud5AtVWEqPzKMm/Ev6rrmgyXqSDfzEB439n3/U
R6scCL9k/6nyLagVa177JgNmSC1YauPREn1TPd9Vml8oalN36XlZzEEQzJRMVluz
Ogs8uXEG3qMI+/mAbaL+7CSdr+88vKL4e1iFThmz86wOQWA4Ow97URKITIgP3dl2
yzVXLJmMKcgQbual0vKJ60467eG7nQvgBmoGsU4diTE2BENxQ5MEhKYf/S/VLXR+
R9CDvu/dOEii/XC2huSEREkGUUwJKrl/ks7M5V82EQC1RUrjp4xTWQ9SBQp4pxxT
SybAvp0Lqn9cf6PRRHI0uRpQVakSx77dn3uqdE+cecZITXEwwjL3M9zW9tjEoUk+
VEcf5HRl8ZsDrWk5qIUPiqvEZEq5lQDuig9E9KVSOiTMk8gHW0C6Fxpx3jqis5Zw
w0hD0JLnBSDAEBeAs9Qmhacfaa1YdMbWUWap35Xhwc+8jS4ja7XAT0ac+Tfy6OTp
/mXHuONo+EAHNMILe8NDsSRMTp3dKE2/fe2eiOsgS6WphQLM3VM9a0CBl6EF0m5m
iq69JYWcbQ79rBWnZ63IRaJBlLkxCpkW+mZPw3dQD5q9hiGR3XBG6seMTR5YV8nU
0bljYi5S21raB7742FsbRzg3sKg6FzdXJK0jJUssed0O6d5VPpWKBVvW+J5ZCObi
ehPErDqIA6GdxOi6apHTVAAsY+hntIwenZp14OR+jrFmcrvsZ7nWr3ayhCExXSr5
UH7Pw8Pwo0/h1PxpUiOVHzwdb2QSJ1c1Zua19e3ldQWN8DK9CY116SJs/v/oZ99x
r+1JXuv0n+Snf5pJzY5GdavCFuRIwA4IPT1wF4w3wU8SHPseGMVuZiHDZAoP5jx7
kmIHWmOIAVGiWKxBbpSAvLp1iNmenZ8D/Ui2NWuY6GWFaMEx9zsN8+mJWtGVsvYx
1J+oiPV0DdoLehm/aONQGTjOrBMnQTEPNOxlFsQG/4JT0KwY/2M9AM0HGw0wB9IF
8+vGs3Ei9ANVpiUAFIyNxgqaBlNhhmzN8uzbadTjedSyiC3oKofeSkQ+A67QZx2u
eOGzyuMNo1tPdVC4RYlEs3tBEmHjiUoVnlxkdeq70oc8QwjWIYnPTgPH2dxJnHNJ
V/CR8ea9gz6CkaEezfZMg7lhadNd7by5dutjN5n2XY3K5C4SdocSmw4AJsZdmoek
FgzZSOhtCOt3r+tPj0dg1H0TAKXiiO0wqGeNScmg3hctikxT5OqM08JmkvnJKIue
znIbxfqt7MzGuRPPOvGzGND9xyjPx4CMu5SUvctmqYNEQlYThRMA0ki8V5LZ06v4
BXdcuup8KcOaIh70ItNyl+d/74RT1TB1QV2WfWUExUEYrE4J2ez7hDXJLT6U43rS
yphEVmcycY0bCgTgL2sqXWplN4qDks5b89uHjgfZ3aw1TN1z43PZzFZ9Yha80+FO
RswNRv0lLTR190UHX20ur+o/TtJHmGvQFKMYtqMxgDOAAlTzAZAQe7ajTwj4LNgK
q3IEVIyddhUyTUKPpTUnNOhj45IMgs1xcwrNbpNrgtO73Cm/7gYjfJshPgDj2HMi
4dInnLTBl2qxInV3skAqeOxiM00UpPQkY7n5Gxq7XyptYI0R8jof8LwMqfP6wzU3
KUrEnv5XWMxw0fVwbQnyWbK94tIMpe0jbKFbkA5tdWOjEULhJglFBaN/1586RNXt
pYqV0QolMgT8oF22+JIrChV0Fq5/cQGRqCZ7Ms4VpO2cYm+P1Esl29sSLWgpT3qF
T8yCd8GMI/QzA2/J4VHaJVXfFmNTtnX9xqaIWHK2XUf8WWXgMcXIkdtcEPgXAave
IS4ZFV6LkBREE77mQ+FP9ovGsGQlKclz8oqgCyoIjxmz2hN7Gty+q+NcJT6d4kxE
DBOZmBZJHRWBFhACtq857p8RS/hVLlK442UasNYbGeq0A+YGYu4NgFSM74ISl18H
pAhoJOYp5w/Ue4DPgta88myGt7PXdocEjIroKRDdlpLEjLKqHwekz4bU2Cz3Qs9j
RXhGrUaN/lJmsRg9XYbXZboVeSsA51oG6PvHho1Cwz34y4MuLQim8h3IKUb+19S5
ZTVPdc5JF+0VU+w53MeX2CJRptHIaKDDesaYivxqEMpryOTtu0DHcgnW2Goqo2Zv
ORNxDiyyKLXHqtSPn6nFyAgbcR1bz0wdtphoph5Cz0RZWdlUlT2f9gbdqg4NRgB+
zYfWVENIy6dN8JB89LkU89cTsaXWP94I5qWPh+OiML7+ZQCsL2WDkXheZOTnLMz9
S3grc6nmvrygILmiBpmi4ntLg5SCIlr/sYGfMWOIm7ixvzIyFCR6FRVGpmXAY1B5
q2Nv4PXMwo8avDP5z9WQgGrk91WRkvPjupnOH9e49Qj5O2BeaoCqk9hw8jWES+us
sH/VzorhCfKoOlBeVpJz+SJYRxqzOZFctU0uBGoJ8ejD6+KEcsRP4M+3wPcng+pL
5SsCu2SgAdYAIBrq1eW53xak6HyN6QBKYNgoWmMv4GNF1DLeft5rE1+BZREQyGYc
TZQmtWOgxnOWNVkTQ7v07wdRSEC63XDjKJJWSomKfkztRDLFYfcNShS9IyqZJroy
95W/xpqB1v2CPh9UwkFr8PWjbAC5h+axOdAyqToyGyNBs+Cri5Pigf5gAYDsZnfl
yIeKmlATPTmyGiSz724h1pJmccqJfAqnIOa9eWs+LyeMRtdn53o3C4wLKwGdvNEY
O0lU4vIbE2yedFXnMM6OX753h9cGagKFo/cLyqvZUXS5P4LzmycIW3zNgz37SsBY
SiOw0qYQ8GHNewZxFG8JexA/sis2tWEryoX9VZYYLdHStX1L752HxzgKi6xuJexS
KCbZSGXDmbOGkHbscJk2Ju6XCnDMq/OVuCLZ7qKtpPdZc96QV4yHHoyHUuaAAFZD
7cZoTFfTDpUBkDxha6ipYalCxkf9CXzNUaEnZeVEWCXzJy7N7drapANsIGLWYwTT
kwt54qGGYpaKyfegOk48nxlsqO2nOxOM3tLte1H2PpZ7WbYOFs0Mi/tybgjFrcjW
CnZF4H3uOAXIKVibAktTSgs8e1GL1vUN3DJazP8PenPKRrl6MUzPD1BysvOQIGVs
j9b7wZzucOVbYqrUAEpgE7mXnnx5TsNdW1X4C/0ttB+AQXMpMcqM6V8NY42eXCCx
RCfOd1TAv5BBS59P0rHa+6BlDzlmvAjRry7VigdELOljSz5AXTyMLYH63nlWnluu
CPB/Cre7ryCZ2vgdQJaJQGyFwASh1WHh3jv/ImweO5widSnGY0DY/BuY3ewHTHEI
k6i0sISjACPJAWUyEQ7ZvdAYkGXcFrjT1PLhX2GRuVT9yBstQYbF92NZIJlDAoYq
9x8LKhHwF78UZEZhjLpaUFIg0PTYrdqhReJKGr0bu1Gv8PV7npr6tJ5UT3H2IASc
ZL4nihw84ylAd7C6wW+wP9thC+ARTUvJ5c+o1FEXv070r2UuX9zzGynpUSFr8Q+B
FyXIcGuvhTsIWurfPx0p+9wfpuZblf1A6u54Hfvqz6xLeJ3bNETY5GFt4s5IXYo/
dPNqzsb4M/x2gy3bjpBVJrPlqy3YewQL+8reHNu0KQvJuo1lToC/EqCc2kzQ3o+2
369MXQtc3bt2zRH+Q6OVabLW14oJhujkwCmuDjeHdSEQoEJjoDW3AwwlCqjtNYtF
NvUmCP5qJWsEgAFMVNx1bQnP0gb/nANw+3+vmcypl2vE3NkX9EmvC1XCZr1qlAr1
IVyE/ht8NBAX5JU5yJya1kIOHGdXbV268h+X2CSU7wrWOMrSIfFVbiqWmTM9buuc
tcnssEThXYWS3IFBXQz4+BZa3pN3voag8FzoJtWmm3GBa0mU2qG/gb9fyj151yZK
b/NuqLXKopoRe49fP7WtNpZiyu59AJCZtqDCUlxl7sT3HLXL26zkALloNVedFd8P
AWEVh50TI0C48wCboUCd/B+Uc03N0Ez9zLRqlOLE7FbtmT74HHoFOI755qIz0/3w
Tuj1qZXTlGcssKsd8cm8CMaeNsPmtpldMvUJC/QxSjrfmNPAjDDr6iKvxwPqiP0h
C+C0KvSr+AoW54cV4EpBcTx2dUMVZEyJhFWKhLJUosRMf4yW8ZzWrf6dfGvu2Z8/
D30VYgGtD6nXR+TKiKeJnCsxTkjr9HjKPCHFjDO2MJpWbCiP8vTXOFMMEp3JlCxm
SHo8HrOSck0HpUJC0k+6dSos1Tn2ktspQ68YTCUz1sz7lIHXvaGge5zeHCsbEl/y
psHZhXDt75ZhSDO8iA05ra3oc64X1HySmCeiuOoqYo1rqzpOghhThIo3CjbM4d5B
FPAgz3A7jpJZeyxJ0T4+ejaUNGDSAKlVDaymMHZjK5BQaGzgcoe7328mM8S4k4m+
7AfaVshamdxY55eepGABvbnm9hhFCtw0urm4sVmDpWDGyqDv25wGl1yGYWSPHwK3
XW6ezIR8HaERx/221yBNcaGCA1eONa3HyAEn+x809bunknshN4Z0wwIMQ6hnxCoX
fnA4gK5MEwHHwu5bPcWjypdU5GU+m7vxlhMFuuCL37QZbZttMie7ggYKG++DHDEc
bdaU0iAC6cTEqyuqbsfb8uJ5MED1JiSOl/x8zeIeIW9xmsF6djcIHCXrp/UDvZ0Q
kfieCx3zALBXrY8PMEh9/tn9Ar1oqLXj5qTxHH/4HZe9teSGW0JR9ITx3vF6ByUV
tcZrXMX+fqce5q9u5OEJt3B/BhUvWQW75RvFS9A2eXdtR/s6vBKoLa6j8KzO20qL
zD0RpM283NTVKnf8/DM8QYZ/DiLzzMcSFsZiUgAjZxp4euI2IxQn+gy37cGy/oiE
5fM2oLsKL9rcmGGMvGMijRl6skYtK3UlO9xKMrBj2woKNJdaRShDJ16Nst9Kc+jn
xHrAawNU3V0uBDu2P6d3nttYI7Lcep0vpNkGG17SMnJmYAOkjLN5MKVpux14+28H
bvwutC6FtRAznAOD2Sr4vp+xv77VECk7iG4N6TOdgcGjxmpZazkgRLdrHL+gDPaX
KrLFd5+REn/dLVMhJfi1ZxwhgQNICWipYlI6vmL8gtC/8/Z/UCBTg8qjshkRp9T4
aXTTe9eaRkvP1wTko5+PzkGNdWst7bfTdY2M0KFCoh0/1c1jTV2TvssbY+aSMB/j
hESgSzn0tdLAqturTMlYQ/hffbvokzoDNXl7Hm9dG1gHWGDHd858nDcCsG9wsdS6
mmbooFeSovlQ9Lvdo12Ksggfn+/hDANvws+JIMHAjYLbnZ3HQRmijyc4uLnBbprH
7yaEGbtvKmsNesA6AagONTqvb9/RlHqRK5CmEad6ZWFLe0O73l12bNJkviAF43Ir
kJF32zNe5fA2QDIoP/hqI7N4+tdmCQApuQFi58yaKv1ouG9itLMMFm+K5UJan7VW
OWL4bOU8/hBOZOfV4Kgl9vpV2dP5CoVsT2f0w0lk88R1vFVews48t3cZSAHneqOt
sHWjFcSBhxY9fyg2u4og6iPpjV3ASpLKWXEqz70EYB8gQOctKbQbQsbKyI5wakZm
pS9822IJydT5VeGkLwjn+m0DdLz7pqSkWB4mgCJbN5qcZ+hWDuXf/IvsYVdG5tIv
D93VrCTwLxqBE1gRXCeAglk9FYVKjdkOXLdPUZPANyRDIy4sXjXutaCvamx4tYyb
xb96gaC6FfDsa4nz8gqdz4YdoXDYpnCdDF2WuAXPC8R6uQBswWsES4QIWe54Zu2f
V+9WO3dsyfMHBPQYLz1BWamJIxQ8Svs3rA0Er25dAnDCrufPNecsHn70vrGWzQUO
daa8dhiXk0bBuqWb8m+KTpE803YkBi8HQ3I7EK2NS1yVlOI8Vj+L6C1dsU4SyK6V
MITCsrmEXjZJCP2QHLUyEzh9f/D9VS0+0R8b6j8mQQ69a6NvzGoKyAvV9Z/0f3yX
EMPfJ3EATEeq7QGFVMCtneYzRQ5Nf5o5l5O0Uemr2ew4sOT2eJM5NhQp+/MmVYDT
McLEEWaesyW8GWWTZZDJhiSklnGktsKq+3hTQxJO+xPAZUjRpgvO/l737Uy6zim8
v2/Iz7vgkp9JkFXatQcKyLcdJ/G2eZlcyppy1grBVAg91ZLrXSGO+wO+WMoUYaiP
CDw8IS03mH9n+FHuTeX7Oc7H8nDnVi3/tr8Oc34vKMGP96YK9+5ds8hMWVxvD5T8
w5d4oWFt5JmZC7J53xhuDwsg87pHLpUD+yuh9qrYa2x10Xo1Q2knFng4+yFA3Qqf
ElBoivACibFrCm1z1b3oHVNDgP5lq5fz7pHMf4SzZr7ViBtxZWWoBdScUPx8inzr
yDBbQuR7y7yfGGUQS3BCTxqBpkrHi8Juo8+96d3zpkpZxi49S2jMk9U23UMQ0DGP
TFijrRQI3KssbSr2uZQpWIjZs9KJH4qgW51pWsK5gb/qajPfjz6LZuVsMpjZd5Zt
WUWUIlrH6MNDL8ae08RzijO03+/fYrdSq9phKojC/mXrR7kBiP4jhPDcZ5LX7ims
D/0cumGW4f3h6DUcEQKE1fALrGudNw7/Xzt9V6LDPTav/EoY1KXxIyV1lcxEG6sH
R9s332S6xGNSMSaZje8dmKWUYwPimpuHe1ThlFlYx8tuQkpNBG+9lfN3EUOSt1uE
oC2tJzCwnBxaThC2IvrWtV9LlWFIfikEIJH9D3LhIppkVSP87998fjkOlymOnhYX
KMTLP8gEMw/dyONCbzKQCTKD8qrEvpOFanbj8mP+c7SQEwC2mMuGEnVAi0pVhUhQ
bkWAV3b7m250/OedYMzPM2W5xg5Ur/sPiSWZuZfTCgqqNS3kSQ3XCPVXPpkYzkiZ
MrmNV0QU6HT7kI0yTQ8RgW7/26nHXizoUhW4Cy4gxLSXlcODSNBBGeqWm+036Y6a
ZRBEX0QuerG3jXnyrZLRja3VtR3SD71DnNdJ3PGggFufXGLdIcwPFNvOz4fzcOHE
U60s/0i0/RiS2AmCawsCpKyPcNLN5FY85O8Bh0DKxi+yeLlxK0jX6RyyrflmqDic
/bplCxFAed9UqK7Ork4gK+SWJifvHjXkWMaDteQGdNg2HmZxkL4SsQDBttvIRWuv
tZ4qHuOYsKZWD1hXgdtwQF3aWmzDnkeB1Xzriiq03dzWoPN4/vhzN7dW4CzBp5Cs
qgxnSpysRTv02snVAGf62H9zkR0NuNGpJeRQSKMj4IN/I0O6DDgiKRyU/K7wRIeQ
XAV0MLTUE74AjD/HBgvBbxd4TxS1VgoSE91SGUsrEjqcBJN/ANusXikOmdY+Khnu
KwlVYds1VSs213tanh4kAOpL129XeWPSLh3M9e+tflex/o9Xf0rtrDEGr2aNQui1
i/2DLhf8ThnM150RbdcnCBF4yebPp3E44FneIZIXsJuuCHmNXOaFICuhCWeVy6by
epnJtgfwWUIu3L0AWPCPl4w5r9z4U5AFDdzj8tkyZj7eXE0PbT8NyZqpWhKDoLiC
HsmfWTsqrhEBjzSEJZmitJWsA7VYpQRUOsBR9cj8gEUR4JphcNaDmj+rYW7JPUA6
tPDMIdoWKIIir055mj9DfTJUx2YMS1U/dRyccM1j4nNNeeVbUYN31YNKqSl8RLV4
J1zC1e+2FyZewhgyIlTOHEzFQd3d/dzA88XJBSJhVfDnyJCrJq/YSjAdcOGBmzCU
xom+67586bvppcEROk6ckf+ce+syeGUXwkw8iNW0I3/fQYH5mhsThS4hxwW9tz4k
LXWVdRgWPX00KHXVvCn5ZhiGML/vKBu0A3Bd43O9xDgvPUxI+rp/Rjepvn+3ekYl
Djozci7/P+kt9Wb3KRB7ExcBkMhy8S8R5ZD/PTxf1SLENvn+wcJuW+Fr7W4w+PjP
XWWGu/rBtPXHEOHw0UNsEq0gP27szrJ9mzCL0OCFcCe+o1jgR1dR0znXKq3aXr0T
iDqdGrLe2ooj2jLqjzF/4s9l0xGtOoGKssRbWhU8YCHyesqJrcVOwp5fHTUNEZEl
5xkYMANPItemWOOVkNRVPXmXCoiVoL+M3VLUnRXDvB+65amtR0dAxh12EP2U1ItM
7SVsjzk9TagXb+3vpth1+Tr0qisrDZ25/xDElW/hcRLuirD7iw65APqVsLc3AQ0f
jD0MnEdSrB2JLwCFp4qK0i6DQdzhECcLhUBPDaRwCfDQkQU25tFjM95nbcwhgnwB
I0LxJXY40vucCA7kXd7hr9OAVsm134mh2D+kFSFY0oCVhC1stUVVSPOZbZXZeTM6
+x9itIgQrOXRLAEtBhD769A6z4lxxxd54cvYNtClD7Y7Jns7Uw/giMfcW49r3XxB
ibcbWte7Rp9+anQUe3yn3QF4nZnwnTWTuofqsfAGo0jlwNHido69mSDpQhA7IAz+
dHGTej+/6nyCRwu9XP4kUdi6QavNqlLSaMRE0IQ4ebvzNsM4xxTDKkMBGT4FJVzG
A+pubm//jP1kNnwe8/ePalhO9YvgP3pKmGLAnphNINJVqSTvfS+sd2KfovNPn3Gs
rhPtsFsksxy9tX6IxPHSEIxfXBKat81SPPSh1XrDZZLxkjqRwhyo5wg6YDDsSfwI
a1ro167UiSGVFHSS1O69hO++55hrQJkIuDf9u1CxMDJWWlSraA3aKP3jdVexUuYL
x1gXW54ZowYn+kxTCw06GobRZg1VVD5b27RoyD514qfaDhqaxy8F38uWixvIC18c
cCc7ImR61L1PIHMxhfnmVqT79uFseF7QSCPtzrBKhIWUSu/p+awKtKz6+7oIVX0m
c0lNdeDo1jsBC3kVqOqv8brvMaGB7jvm02c1kgjfRy2DpdmaZx8N0hTz7+qr8ofs
rfd3UllDmPY4z4y3nMYy5yRiiT64l6PEWyalUN3jZhhknln/teJrJIBJ/JHEonwC
nkHm4G9OBncXZCoqME44iHUK129KHk420XiimwcVSlX+O8DppGxo9sbLqvEWEo7D
xrsyL9zqagmy0GTsHXo0P1yvnz9R5v4e0Dw1EspoYV5p3QCJ2uzqoRQSCDK51Z8U
VaM3ycg2uxicujAO0zUDEnF8A5IdhwZaZT56qrS1P7RimNj3hCjokDA1ExKbPmIJ
ht/xUxxcWSHQIrXjJGuk7uj8C1bBXznD1hDuN7sD/RFmvhmFxXFc1YHCqhlSqhuu
AgUCjHR528jovxf0DPraMMIDHGrDvNzmMaOaXTxnf7bMJiDIv++PxEa6wtu29X9P
1qgF1mDZFLwwJTNDvT39udZgDNnaygKLjuTZR1DJzJVOL7RZ0pSwf2r+OmBoq4xP
mxGeDHtYdWYGAt0SmBQ0mA0KXi8oPnYJiKj/gQK5fV6FnxWofyKD6lkHqHO29WZl
Plj6KIQlCXQ/bZ506YQ0TKFZwYEqUFCDm7C/nArq15xMX8Wsft7VdpWXu1CjOgxN
dgba+hBApDyy1s9obyM3pZPKu+O2UjQwqjuTq2uG1dMzx3eYb6ShbUxc5hT8/Wbj
ZGk2v4xvnAPpwNoShjdQryIJQWfKP3/i6mWmcHKx8Ug7+iMqKp1DkwVloLQayaV+
AXyFvYDlqxUOwxjS6HbhIu4wTCUta5vc7uwKCcevadVkjR7qa86RxLY2+cBMtsW1
RHaQnX1OSmKvrp0nW5S+FBinTt3IiJwosywmpKXbU8VNS8hN0enzwT6zQEsM3rBk
XIvf1RfV6EK4kicacf2U9HJuAM6hdu07FvktH8D4Kk50vjeDDoWxeVxfrmJIdPtf
GbenLixpTCgoVJ+DZ0BFO90fXAmTtNj20idtwXhQZsWUUUkJ3sXRIGFaeGOP9xtV
Bz3QI0erWuXD1rjeK3VTFqEiM2473BMewM0Cpaj9SKoBc4u2bAkrjwoVLvs6bmsA
n+Uxu7ziX6KpQXYj/t0VcFmeaW+V9MfmM6+n7DTSOKM3Gf26V8iuWCLOaJRBJGKx
FjiXSnAmEgKxZ5kxfxw1mSqqebsBMOCl7qGk5FEGgokKBd1170IV6EUxec5A71B1
q57GwtRbcSAXIIPrvBaf+ZUX+NyEQ+NShte7dHIat0e9vOOlLH7exBcMp424pDpx
x/zH3VR4lPGV8TWHLTZaPeDanJZIPaRvqqkiUPN9tVkzl7IxMRPWFND9yxvSz8Nm
WBd/usqGDd74SF79qVpFlpkb/b115SBbtiP2OX+Z5JJVBmihok3z+QoOczmNW3Gi
T+wFEvBwEI7LJHSWE2bzBj3g5rulx+BI2PXrf+zwnJUlIvh4kudMdqxBxSW2BEde
yK89CJ6bUr2yIqjcXJu5mSKBW89vT6sXi09ASL2BRGaFHsixLy+waEteyFDwZJLn
tP1iXS4NNQLQRegWPxNmbGPJ5mC/reNanaoITBLarxYN1tQfCYUHLYVT2iCEvSAo
geAMXg+H7nnHRFUh8RRBJ9sAVU8VD1Mfe6ynrnPrdcEvsjgo/+vRAKnfw3a3y1mD
lnkml5809S9X4w6u0SV0zVfWBv0QmRdR33Zfb/9rERPUmv0mLVkTW/1HmBAPZ0qt
MRSydN5hLgA5gfLi1Tsbh7VWimoBcutYFJqe5t2NLR0uSq/6g3xWwS8RygV6jwYU
106AKv/cEaPkgHwQE4z7QmNcpbuTOL+kCHjNsFOeetQ1/NoKC420bF7WT53t16OF
hWJ3XXQypb5TqE/MKcwpNkfMSZhrHfasDf7AVE+4XNNCVefh3sEAE+bLBKzG4Jpy
RDgIq3CZIxFCkzaGbkJxalJkxaNGoxqVVFIAWnhKbLiNUq2d0Dpcme+bCpWHeaiz
05KIWTeR/PNQKiI8+aMRHh6edVwEo9Rrp9vwPuqAWnF+E3BUjjtPk1/9CizBBY3J
Wo+GCyEBVE4hWmv5J5Wm0drL7N7euqJL3nnZhqHGko5QaZ0KCY+x1xIXNR2nc5ks
SvbaeYSGZS6xaxGUNlSF20WBVb70qta4vgwmxB2hExf76uJpEED2gbt+QX3Kqg3J
kBTcDbfpWhqTqoFBiNw3HOtv+n00LklUgOpl9Lk3I9PlUU31Rgb+A55RxDW2YwI9
jnWVXTFVWwDPFzx4ZAsxSMSbMlPMI+sfYkgxhEe1ulHXNSgKEAsh0ufUdPeHntGM
BD156gxEodgX6W8Lv8NIt7SppBDrega2mXDAfcfAna6lPEDuFtxC5NIXlokOM5Yw
bJGFOqEu4TdGZqmD4Kk7tmMR13MLvH8tNxzc45+jOd9++HDnt7BwgjjAvSroaa0B
dkbEQgxzAmSJr4+fj0SptR/zCrne6/dTlLnRuj7tIvZc2+irwkkJlEEliezjbxZy
TtUbq9WkUr9BmyTXD5ZOi/sFtgh5RkNRn6si75t7K260kEepPKKJ5N6b5m3o2Ikd
DhdiAwtWbIRXURfXZlYC7psx7+ci6/RJAmS4fI82KZOTa0AvY+/4wGFqsGCwwBQv
RV54oYW47dvPk3ax2e3uBxvsGyDjXFqclXK/qB5uWS+Rb1+7OJEuFCcE3vuQdNER
zzxRK1OkxLGvcfvHgneFKh5C8+1C9RPRUi1GIqVu/wE09i1NbRuijhtOhjAzJNTF
57yNY7wpiSN5sqcjkh9z1DpZjAMOMdqZHOXXfdrZiARDyHCVwmUPugASHM16NdsZ
1f3e0tHBQN9xQyHm9XR0+vJMMQAH++5jPv/NEV0udRxp1Ij2Pms87qhAEhvzVDO0
+wXyXoaWlny9zgtyUFEVDALPAbd0LMBcKBmBtlPtN64tuglSFI+/e4pH5+tQuedx
xJGfRFXyhskUdrKKER4+QrnSqeo73vmpTnJoYpehcEmbxI1romkLnYAAsXw4sbZG
VZkCrhyql9KmGva5WFQvsAC/Yo4CF7NmY5B6kBDUQUdV2pgC2FiUrAABAElPE8Ye
1lNmKzvLsenZ8iXOC3s5xZDl4MvKbRaTt6eP2aSxTBbbZ3KHx3ARgk7ncGA+bRcu
siZWyQqm5jKJEEvQoMeNlIGdVGJ7ywfylcJoy9w0VdOaPkJ5MbWHJR/EYWEFaMrG
+XS2swRKZb/TN+x+HWRXVIjgG40OUodc0PwDcT9RKl4DRQQPEJFF1kQ/yQ6Tm9pX
c2s7bqjAVBJYnPgfnzKlRTdJlme90xIsDDqyDu5UXDxAlGJ2HFGS9uDd8Y5/rpMr
WNWVHBnFSYgRTnPhZ+q3A34FnSAtfKMils290dR+5ZtLnli+/TaB952RLwT+/2VV
8wOubH870kCTfTXFM7Nm37cZ4NoiCfg6Q+AKqHgcjY8A5EIiV47zr1iNOtgn1EnI
YC/MZB3Wvstm1sI0yLgfrJnSrRQfNMRaxhmIWhnCD3J62cnayk/Mb49p8bNuqBOH
UT5KEUG5ysFlj1aJ0M41yPMVIlT2bEHTk8PQ2Zsk2qfc9MtKIqtYTBNJTvyGNTaG
RokJ/ggv/aFm7+193J220KGBQKbtk2+po3SIZ0+j7yfRp/mUwJJDYshdqgA5ZUsK
uUBBuHyrUDRMnfJO6MRWjoG6U+GZJ+0/vrwnLTVOZqZ1HxlPVDhEWE6j2ud9Q4OU
/FmQZqyQgXPtj6qRb1mWFkzeb0M1OpjIf5wN2XpdKLVcFh5vc7hrAlV8Rfh3zDPD
/14iEZQ1gU0MDhjDdFAm1LxJ2ugaGPTVOjdjJM/samp2lMJDEcEfKDcvvo2HX35Z
vDgutYqm6HR9PNYfvF6ZCHLuIld076rCqHMQFJuVFhW0s/OCii8e2ZMO3UYCgsMY
kg/S4TJ660e2ALeFDCbgZW2pTBYYO32D6DvMg/fE7+GUewdY4GLSL4qBNi06UuE9
WpwydFkcpY53Y+D3VGd24pH8TyCg9JI/OJKq3R3uGqvqk6TnWO2tCtqKm1iN8i4C
NvxoxZ+kXcEwygYHONT3MT9cXx4zuoUOihx4W3i1vgJTqSdhh1l/7T/eJzMP9eSX
Pi4Ul6FticHDgdZTuuvb4tBmSe1fK6cNkKqsDn8oq9PU77lDrmK2/3uiZt6jf1Mi
5MQnj2jICti145LFwQGLBnhyFOO75Rn2xfHmB8iGQOA4i0h6vmSSLVWBm+PNWyhN
GfHxDeSKz4TQc7pAxd+eK0qLRIIWM0tqanGsb5e7dQvrWPhYgQzX2NBLFPVHQ0q8
2mwwqzUhUDPO2lT5a2juH9zrX9W2k8uWHoX7qONLtZv5LXEf++NwfPr03pBW0BBN
lSNIQHJjaPNGeXCGZDsunv8YJedUCgpg5ZNF76qCbvn0KWZ1PC2mhtHrNxbdDQza
DY5p6Wsk9AUXtV11Al9XlelL3Q8BW6oII5VL1/IV+Nl8rwNsjX7rQRE76qaFWpBv
CcjgdGD/moOyvegX9ym1ncqmnv0kHoRx3p0GYXHXorFl3GgmH+Z34KQdLZ7E+RmW
AnqyVdNFDyGXYGnOgWLobJXZ5uqG2kFUHEncOt3NUGI+wK0Ilwc1qbF/gnNAfDVi
UJ1uIA6GFCiSpUcGt2i9G5rBe/7WLZ1AV74lvt0bUYLPW4vOQppRi6Ck0mqG6LqI
z3Xb6SbOInYbIr7bR6wMpwlu1r0je/O1XaxxEpiVZz101NmYmzcDaw+Ejdn6HcvV
4em/Ps5Y7lQmt418QWEb1iV6a/70fwbJswciEpCapmrPU/FSUxRcw0Tiyi2I6wr4
f+ZNlMGKmWE3Jghx8P18iW/9JZYDIHEwqgJoMmziN6oZXDeolytq63IULMdUJmyI
7MVFvQ9h3pwva+gh+omSm/ECy2DMKPNEoLwik0PJP7alF4/wYgHbPqkDiRMD0K3s
ygeSUTuMcJXvCxF6ukoe/+w6tTJMEnRU1gjfjXF3cfQcrrr4FI0MP3QgUng6ed9o
59kKA6KrB2w/+3weFUvdcb93Eg5ecNKQnTjbtPGKEWid/tMymw9W2MdSqfd64Ayj
Om9ES8Mbg53l6mH+l1QuHe/g2HiKF3rVyHjIn0vP0IHX9SiGY8n/eszQr6EFXOhw
g9U4IfM18TjdDclNzvb6pDnW3gbNNwpwATZ6jJQ4zoV+6mWHZMtx28/2jYWYQ7Ld
QMB6C50kBsHr61JSYrFGKQjpv2lfKw2fcUthyuCHPj7bvX+55INaW/lMkb6pZ+D6
zn+42/91ZVWS/ampIJ19xF6HBk2FPMaS42fvIt2aRPPV2raDBZ5iqNvKFncnVaHa
rg4YWaXveFbTSprxWk0aWz3C5QOvqpG5VBC50SNScOTMQUOIz2LCj4IdKmGXINN5
k41zBd52bv5HZqorZGNPI8d0AT0GQK2ExoFdcpRHdMqpoDWimP+HntG3Or8oebYe
0LRETbiT9uvkSTrwp5nRBzUWZKjJmjFEMKgacwuVljTKyLgHIrXvs/h1Kwwj0RpI
6OqlBm7nhYVs5mW5lORBGAQIZuI9tqOG0JRs3bfNpTQ6gS/cDIgTRsXeg0i7+prT
eQcgYCJfu+t1P+FLiPD2qJdVL0VbWpyyRUxxvG00PRhERNrMnUCtZBSIg9Ga6E/8
3GehrL0/+NzywK4cDxndoERSz2zDRMg6kpoqgv/fZ5987EQ+Uphqp5I2YXbFLRvR
pqjOPT3TvgSK6p8QfynAl78js/kO+XtyHGloRlreB5UuWoKmjaD2qquhICcieUei
hQze9kj3Oa57/+3oJWrONo0WarXNRmHC1jlS6X8pq8xbH+kQj8HWu073UJaD3n5Q
oDQHDxKS3YXTDaFmZyfNYrUvAoR8gwO7rtU0E2aJFIdsH1PdsbpPlNM2XFDiEXcb
6IANtmvA2F4vDGqPq6XK+Pox839kCOQnGYE+sBFyI4JKyHy8i3S2HT6238gLZcXa
lOH+vWOQoLHOI3jQhai7Mmsugh8+9kQP0yjLv7PMNvS9mdvzQAU8e0K9SmTDG0rb
k1iqLPpAdJmBtDrrVhraXEtWBerI7huqnV0lAgW2Is/iZ6Pz2W4bpHSOkMW2v5fo
hEhDOL1QgsCiYmOu2JeyqfEQ2wfXhDiyFfFw5OzE1SDLbjf7NjsAF1gcAKL3pYK0
gUbw1xD8mSeqTZHBavp9f9oedF09aWzjHz7DLPjxKjcTkpMjLq5FJGqZ/y1TlW2K
+I4XiQuxQJe2qigNGbtX7k4MziUy2GqBtrR7rprIllw9urzwUicTECM8VenLG/b8
Nrw1zD12uwSQjmT+JkO4wJMqNWmfCCxsteQWhDMC6tZqmnUymGUj6jElC31Mrpdo
ujHIXyxsAmaDVyOJcDWuzhHGslR2LPQMPwtVRgGTJeLIWiyqfcODjHozOqAEqkV0
9N0zrewKkjjjBnksKtxtSPT031HLktAM7rnvWODwGmfSqgibcLGRJfbk2TVYCrBc
9E7KJCI3s3k/CDdqZH29Zxest4C4gMtynfmRzao4yQvG/nF1/tCTnqiSBmjQvlKq
2gWoVHcjkJhrvyBgl5UyVTDfQ2z1Rcf4ld4kb6MqsVhm1TxuNh7ya0kFNbdGn8f4
z2xkXHaJluHzXaLVorad+ZT1diwdnJjoBF5qFJ5K5cZKGjRa0W5bxY+3e8/+6v5w
6uVpxS4d5I9P0Y+5Q0nH4jBiwguBVz+RWJysRMWNMpkQDA7y9z8jttJP2m+vUAF+
BWcRDLC8xwE2aGE0UjAUvewTFxjXiT9jreBAOG+yDYWTrjJi1RRSSp0kapOBNw9R
zcO7jWBAx3lpYIG8jurFWZzGL1u2yPZs8wNYPssxdCq8VQg3R4Pw74icPvUNF/cC
pf0B4auFq6+IKz6CHnHDhfT4H0XyNQiXjj2ygLVcHD+/vNt+6Igt5FrPJ1PHSe64
gb7sZIPV881Fs7RBaMTt2+c1C/chqLG3xJqCM/I7z/OGaYGfQYJgsrF2tWMvkmPz
8o2eHq6Wtc6KZTGLn3dXeBdcHj8PXj0vRNqnVjksQGX6peTpe+XJWWnVc+OrwxNf
KHUtvq8Qi9NVkPOzpuuFc3kazL/4gahm1AYlzntXy4w6BKeZi0frOUqEVsrodmKE
wims4JhuLRBLWuvP1uVlDGsVgbRpMXz3TahDdAtZw1R5bt5xca7skGmkKbi6Adw4
X48UMMxcGgJG1+rL0UI+CQYzrsVi+y38+BGYz8OPBP5j6kmcGnlhnsIHx+nFY+5z
EVfi5q3+v67V6h1DwWyOpweIBDmdpDdhKjzPsN1S6jEc1zXD2PdszQH+qKp1DLgq
a4+vnaD2Ydrw1Klp/zPwCl74jHOllgeUPhWLygUaoToZ0+dOlUA6fFrIFFDovOn/
dfVIFJLby/DyXVv0+5tEJKLngXSJz32lySauAQV3aHZNmSjW+0065PLJ1Qh0zgrU
Ox9kb186Wlv4BAet8WcFdPxu306e86SofsCgIThM46+0dz1DOqSbDCCxuymrGs0c
CKyTa3R+z8El/GZm/Kqn0FwM1OhF3if1XxsSKfS6SwnwHc2RChfXnzRn+KBPuZGn
4pqT+lGU/oFWU/L6gLVs5EH3VsFtuBmfX9GwTx/052am1gD46Dvf2m1BOAV4eLL5
vtL1UVisOLitCykfcraWhllMrNfQ9OjkInErk5MgHnUTVz+n6hG08laLtM8fteVW
RiRR0qz94m2c4h+8oPPKFru8FfcBiNgNDnQG5o0hX587NROvOp4+xyH6kY1fc1z5
kUCE6ET0pBQjQCUxxzU3TnDcvrA+HWEg5ziGxei30ZFrlHBNiqoqSPfORxW258Kr
jYDYFv9mh/c6I1B1Ehp4NQHzn2IFc1+so8qxpkBRzgXYV00w9s0SnZ8HPmbmEyVI
HaWN1uORNkm6x3/GIRS23V2aUG6HmIv2T5eq1c6AHeH7SuICtyy0+/HawR0KLloJ
c0t3DOvJPT03bQZ5HlJN5FzdjY4sDcPZ2DYqHED2TELzeVp/3sTVrr5pW+31a2Qf
cbURX4BYhh5U4eqKJxGnGvg7YPYcB7v9O58qCXeOZ9KDhxYXTYv5L0p3atkI2uZN
s8SUSVxH5Zx1B7SggdobwWN2CWvC1GWk3Dz1baPbu3FdBKMBzMvddXVnz8RdihiR
4P90yxcNCq+h1OtSt7vCuFacVq1bMGNjjB/Cl3p5Ld5S8Sb2fXHWaehEOv9BgdAs
ylBtd2YVgN7GJQxKL2F2YTIKiUEsKZDM6sT8wxfrCKETr0gv5DcnaS7kHGJu5FUt
jT/0JEQXaoU4YOdsKqq9/P7VmLIOq/RfP6DflEdwOyPSG09xuk0AbWX5Mxa9BuUW
hbsaW6nzqRoYFMzTUBJQ0RNv+r1DabBsAgvs3aA8ZAnBdrFzPjFyI1yLKW1Ix/qr
3mHmQJcXlpjAxsOd8iZDhQH9el5AUBbeTzqm0MyhWaZtEfApuJb8sDEPg7pli96w
X99+UmdmDZNChoPKuqWGYabuGJJFbiMrmeDgbud4jGb6sYR8tGo/Wc1qUt6WuU9B
hWtPjCwF7Rq1xy2wT+0UvtexYanGdMcdujn7IfutIqlREZMHohPwTzjIdXWVvVjA
5oq0Q655KgjkqJC2qFhW50fSoLfg9fMY/TBlEfau/Q/HZgi1QzKYT8kAF+w0gf/U
NtFD2YDfEEDNig7JHMHOXx4EytOE/drwrkGnc0azk+61BHrIpH81NoLfo6HXWNoO
mQESd2+JdyAF2AHYfCyUL/CkLuzu5vhllqjZRuDuIQiKBrcmwbKFb6bYpTbR+me0
3GV64Nph/BDwXyDVeey5wh3AxZU/N4FMLkBzFo49v7ohmuOYPGYEdlKhrCinydMx
gV+eziGExC5BOpE87e0b1u0Nso5q3KG3myyXynEj1oDhpucDZkVyd+6KcMyL+aM3
29cmtU+pDd59CKxQxyaFfxPxLgryxNU1IN8Rpm5oPSquhufxuYvu1//0Lo3dhCrC
LmG90BfDzDX3E0VriknaeDfqEiKkEeTCsqMvpH4xrPkPxSfXnVEqbz12Z099Grpt
//ZK4xPVOstAqkiSuTFSyemoLGj2coRJyksVlvc+0UyvD46NChwT0EdAVoTl1i8Q
3Yr8VtIP2XxuibIPdQn93w3xz+A8kHI9iarZXYHOCHsKZYFVCG2fiKsysyqjhtz7
RsNBqMyy7s0J1iQTWHgJ4QAErmh6LXJugicu9LiovNsrTqOiBfmwLi8LKFBQntsM
qw8sSx7wNNYbcPK99pWODtU5d7jxI26Qs6EBYgS9dfkUyJA5V4bVIU2bo3IPlXpj
3QyRiDAo1Nhj4SgBtmHfSgavTuSPaC6aA2xjXIvgOk6oF+hCFRuClgh8pJMny9mf
/1g1wPucFAtbaL3aiOhVFfRhaFIHE6UItrukTIneetJogxmOfJgbzFzJnmt1OGlS
r2HzmOA1l5mxCC2xuyMnJW8Yd6gWAlmlMcozduWGqNK6bDPFVQAiFvPbM5lYk955
Og/FOrMfP+NOIyqfUqwqulk574xfeC8WleG1ondcFRgVH4SacwxgmC60C2wC6NNj
G7tRrYzh/fhq7pdT5ua9xaRrNQL++q5Pb2JoLoauvKAOf7G68OCxHMI4J+XGajcz
9rrQpHbiPcgo9j9yJrB+VTHCfrMKq0ZoAAnw8Rsxl8+V+lKNjK6aKejun+uq0Nnq
GK47P1kkNcswKWeNa2/FGQWiAcJLGG/t+cQp+Hw1nGxCC6YvQID/AiZWVS4R6VAP
uYIpxsYk58y6Pkpz3IUOZ071UwO6jRJXXV3YtbM4s9LQohqoiMaweRwAQBtlvO11
kQdCG/6QJj1lRN27GfxKCC0gmH9AVv3ROr89mcUDAj7Y8W0lsIuM7LpatYQTIiWJ
zV3XDl8UibCduCWvX8xDfx8pA6slaNGh7q6RZqJbt/E2zNNsB5lfKGgv2Q+lgK+Y
5Sd0Ax0j7yA2S3NN9EpiumKUqPqLdbg6Hh6Fqz6tErXU02eayJMXbaXfw/L4Eabg
wFCJYHojAjPoNfms8pemy8+PhMoAqXKApopSMX1rYqTi/dQzcOzzimVN7lvkVKy/
xxXH/Daqbrl2eMa1tE1l7vDFe0nkw3HqIN+DfIl0uW3rjw4JhPB1gNPL7JSeXTkB
yDEmFMGdlMJOJNEOEENMQx1Tej485GD8GdEnNXaZwl5WHDObahnWU9nb71eWUp9t
qqliQtWG5WreZNRIEl6/tp925pHxSxtuekE7mseca9adBd63c4XuqmtOkIATSkee
JG8IK1ESxeYk+M8I4/3SBhmDNE9kQRXCbNNaLFVkVMtdBdtfzYwGGVfpGCObLzep
EpocWm1wlIsiddFCpV9a0ILy07xTdf5ZZvMMXBm6H6b/AKmf2xaVsFkDrcY7t3TH
S3y7YMovc1xZQ+xQdOBxtE36in5A3kAQnbtDESHsbQceahtHEFaN1PXlm2Mu8VsG
OT0/2jmfbxGiUVIC7jvYFO5qmb5LLywMifU4zqCoiQg1k7c1O1N8P2zkGrJtbpI1
3lXoTZ0zjPZu/qDmo7gz+9NUz2lIEmujCV9pMGcJXpBVh2aNafJuxa5Mkm3+PV5f
ufGkZPu56+Ncht82LeVHCsGLSEgWgz57fusNFeDPpgGblCVcVgLYOacZpHfhou3H
UT/fCjaBlNdFUT1mT4yoH+b5Nk4CjIsVbFx03HszUidBdWPO3N3R71tsC/HnsmAl
bgbnPvXa4nBpbmnLSRa2gxxcCwFyH504ETnT/DOa2kMbKUUXUmTL9sAjHvthYW7B
CIMc9DoE/UE8Z1IxGhSde3iUD91o+4JjmcpQx2wjB1XHsySsdsA6AqwiGDPapmUY
OED/jJ930xxwqyH7XDoukVixn712n3n5l/iFXH3l27TtRFMlFF+G3JR0DOvisjP/
FdAeSvzc9RdoSC7XD2nM6ZTwQuRnMmmJej2DyB3L2L1Lh/3cWE+Wq8BEtJUcJrCN
2Un8X4uHLkC7pLMUM4JCnWrBpTGrb9wgfMMVp7IAtos5bQK1POMQpn5gS7Q9GCs6
zAvDqTIRvI/OteBt+cwZUjOUmkhCogRUkFR3hV2KB2aHMQP5R8o3FeLugSyjshue
8hSJ/91dpWGzt4PyMCQunjVM4IqmRRKV7tGvp1GjEbnl2JRXn7h4nZSJiOQbhq//
PREBgkKlQdADm7O8RSJj1ZHhgCskMe2t3VUrS8Z4+nQpMLt24s7NccfQxhNT5rjq
ED2RN+1v4w8lhD3KvV5IvTjjGVo0AcAEEMRaEt3UqgV8QFsEV926NTdv+ORkVjJM
pAUoruVHgzlIOLJgUx5R3iYfyB29opPY5ZAYDQ3Ax5TJRaMCh/p1dUerJwRDmPwL
5/WxlGXTDHl5sEA8u5P44mchy2aV3+CNI/aohYCVgP7/9Jk44Bta8b4/cZJiAsw+
cn95gyHNHzsOAvsDwZnk73lEOG7Iv9kasRqCHOu4Xjewbrs8Hr29beykIMT+LxXc
sMltgI8sbpMHxfsi70A5z9NpZiye/Pnsf37cc091kgsxp5fdCDDy8wVlgaXn+EeV
aRDop6EwOZMXT4lx9jn9nwcWeRMrEizFJOGgSEVK/jpVrSIpA8DXDQ73TO6O27+q
xeJ8s2uhXNj9YKNAOXPNBt2zsa2Q4UQh9ZUBCnU2H6oxxtXXdzMun7N4Wy3n3+Xv
mLEoSiBUOtbiAxzd0wxl5eilL5W3L/WgiyKwk9Gdh5gE9hFt7AxsTGSpcQzQYKSi
JcRg37e9oardGi/T6ImHVWV4CdR/iZwb/9YUPLQXNh+ky24m1yKuX1r2WAy7AmWw
lV/GyLLiPhyeK2b4eXWWc+lMckEPOlaR5+rVITIjmRdYbhBHww5Ub/++di65P/DC
RsZFiP7Ak7PXO/XeZc6FE4pO8P3Ba7L2B1mAO8E/jm7qvOlr9j9mSZs08VWiMGAb
hLig2GudLLdCBG6HTmc6EZX0WhFE+c1OVmkFOIzL90L56zmg2nYha32urthrhq+5
qcd9v+Epsx70wZt7uZy8B8CgD70x6d9MLQ8hCuWyPfrH4Lhgc8Le/V8WQd4P2dPK
S7KmSZdx2gARyFPKUtdgS+K/RZ6Ea36fhYqU2eUjXdCIxOyV+Nds45TUCSltWOHd
aY+BRG3dKVb9sFhhAzq9hM05OcKie3ARiqhgEyG2dM5WErc3v/RQxHFzOQw+Dg9z
LQN6B6BtCEOVtbivqg150l9AtGsoTho/PhSBMV8jjcYSId9B/rPI258/ZXPr/6a6
qhTJ72xs220Q6yipmxq8wTF6rQ0drXd9uVVgbaVkZiw2Ld4y1OeBHgv+hMlMLrcy
i36TgqR7RBs0ZSnfwHkWyIseENoMcehp4Bf7chqUzX/yphzSP3LQj5QFkp0xTlUt
qpCs+rfoyk4zfVPejtYuwgl5FSJ2y1hHKrQ3nqF42opcUw9IbCMQ94YeG2YMfRS9
LP2TA+bWAvLYBI7596Mec1IQimora4fYZWE36s2QkTfvI2OevARpWvZCLwiTGISQ
8wlMRUw+bj6Du8jBZ8OrmxLpfrN2umczbSeijxxgVWWB0/Y9bWI1Uvj+zBu8FJRc
hc6N1odFC6K3xEYy4VMItQp9V6iKymBvk4aBEUWw5xxz2QVjZNtvlW1Ntcfv9qOZ
taC7dXYDjc2F3aGNSJHPlLZVIAEFHdbJRBVAXR5XhLfXNLD3LdDoBPqia4DIQ4IM
wDwM/Q+BvJc3XAYItkL90HOKesuCKhwxBZ/PFqU9kEEebem/S8PVrmXNr+E/p684
P8pYjCzwRATS4AVAC/6Z3/fP96ybh6NiTR0PRvzrl9cZbMJM5nDZ4EZGx1FDm/iF
4dHkfwj08kfu/Nl1lu1gd5GEDWJomsrcaN52uUdYHXay08P7dSL1RHYpnXetb8tt
QvkaJgXNRb9c4MwT93dEcvUf2dBCmyZlIGR2QwZgYJ/XZ7HRGwan7oq6EUipYqXY
1i//l4hoNTXW6/XU7uB8NM3Y0dXwFMSqcN3sTTUAcMhu+kTT5s9TW5/8gw8ZF8mB
k2QMyGactNHAcm9PpsNI14Cfyul6QOW7lCP/V5BRvUgiJeWVln/DYh2/Q6ElrJq8
1nQONU7haEEYZh4kjALmtWXw0TxP3yWqOGazteS87py/e6G39ldvKw9Rr2QFHJ3n
6cGVbjQGhcsyM8mJmkiU0hBQg8AiBPUFVXiFiEHxSTSwrotVcXHVgkUZz9AmcG0L
vJ6Uq14BY8rnrwkFPB+8MJjFSGBHOZ55Ew13hEusiE0fI6iVx4jCJLf5/Ah5f95/
8krumGhjlPNUQbNx7PPJGcTovalxDCV7C/3HD/c2Xn+j16xeg0JE5R9xiuqQ273+
qEEfdLv+l9BfnXHV2BSN2wFbfIWLooz4iVg/oWLvwivzLBGWuKJk6b8X2H+ikzJf
/aZ7P3ctTfxoQ76DSlT1SE5z/Iu0aXozgq4bcDE0RfnZUxJiNwgeRbLztHSUjyxr
/f9E2xg/OEzJIoLsFbm3n0ew7GMPJn7eNUqFm1YG+QVnND3F5sFnHvdbjAnx+qax
nnmDUC3WP+UcnFfjlXz36YCae7mlSgEA/QBQ3c0swkYzkB7fspai3+7ilc6Mn7k1
0dzv9VmuLQDfvlVEfNDybHrpzX5nEh4Ft1yeZb/ZNmigNoRa22TYoI1X1a1BUdxP
wLTL+BU6hoUZ3eEqQFFxlgddVXOcSrGTDoTDqERSpsM6ESeVATv/U3nQEKNaS7kQ
U36O472vyPE/voP7Ik0z6Q8P2kc8U7P4WxpSLDj/Fb0MyGNWEKq/EjvRQrWT41Gq
9pDMvo3ta845Uy5aaJKVe5CVzSVrk5c85bDENh2t2ojVIYabYYIwrtKMnpCrYDZo
zGH9QfeGpp8Vs4eMlSBvvIBkmJwY1s3n9PUPvgaeqm39ck+VVdq4Uyf1siTNwzBC
eu3b97i73Ta91KuT0nEgygbvsEZdsDE7yF1cyeB8IxIbtTCuKtwjep7GdAqdfSb1
xFbHqyQkXkC5qM1MATLCjuESQv8+SsyqDiN5sBE+aH+EeJuKTMahLbN+ekiLuuUd
0r26HFbg/AxMLqpuF2Vp9A+XWnTZPVwqVRLAhQGmQHaJ+6S25iLslwVbRarHXrMk
vBWYeq/uE5Tby/GaQoqMwjx/fixyEDActw+tTk2sn5WmKUIPCzwgrPQObBKzFVyI
vRYJzC0UqZTOG4uYdFAfUfdrzjOxJe0Mp2QWsKMJUsFn5sQ98RvvDfjUq8Hzr9MC
nEea//BHRfC1bPg5+V2m6dFQTUANvKiacgwBogdTNO+/zN3A958Uq5VKAZlHGGrh
g2aTeK7VXapsyQQi4zi2MTvKYp4i4sUMOJJEp7vb9B/G/GJZDEYkZf3oxEan+fwx
OjYJ5MtRgogNtHmwvP6+1zNYk0Kf4qKEPvmR7c25JkPdKrS5KIdcNf6Cp0N+Domx
PYlZ3R1WBcFV3NDHUNyGEGP0Fg1MmNgenmO0iA+v0Y6uEApfc6IyX15c4cp2+YBC
LGFqhFlqPZMWQZektiJ1WR0/G2pJJxHKiafkFVenHRxAB6NXVesfAWv7bab5CV7q
4+ocbP8PZsmrAxbuODOCKTlhWDFcKYacS/HZva/h90DqB3GYqPGUkdA251pRa1vi
rEK+KxrIAO0SIXSd5JY8nMACyNX5vs6zf3e9FMWP39cUURh3+ztqNfw6yEh9+f9i
PmlwWNuFHbuft8H8wgD30RPYmj07UTeacMCVE1jwSacrgmv6SMTWc6IGorkTyF0T
reVYfd4Prwg32hqjoaJOVostWB2jWyJxSjVMNoVk90yF8wH6hN+B7gvaISX6jv9U
/eL9qJRC2ZL083JT+1GKgPUinckwU1G5vuUR9GoKksDxe1skNOwM58ICEcy/lCkR
I+TTzda1Moeb0BrWWgbVXxbQQ+UHbs7Tkcjxi3vx5fD65QsHh7tlB5c9rQWgnmba
qLOyoZwqhqHtujVGfldnkXr4Fuu2Y1vA2Ywzihkq/BFYqSV8rWFF0B1OGcSN6eH/
h/4QtwppUlFJ8rpQemRaGzsiwAYQB4R0RAhlX7DRlYB/oOuhuNHkN+BoX4IRwhzj
a5TIH1kTjePMAn52wQCyv5Npte9ImM6U96RMRm9GkWKw+jYAkSRBadX74aTFkOzp
dzzuFEUnGnvHCdfxv+7XO84bb2PAltm5x0UeGIVuT/Is4EQDdF7iF68LQ56SFHXX
QX6G1hWVUIRI8qfZ9CyiV4kXKjenY2qbNkCmbXBSwX2JciV95QsOMKa7e433Cbhz
+AnYfGIbaSFiKRjFp7xPq6DAdzOpTHT1qVdskmNmsV5NpNYyr8Ta2qvmmxUk/tAJ
77+xpZJZdJAr2eTorLP49Ext/3c8Tl9M3SoeiIMpLrp0x24RwSqyAgoDDRJ8DJiI
+BNlIRo+GXadHZnSaRxZw2OJpAnMIizY7xHWbQa539Uxqz6Vip1KR4z4dCEliBrQ
3JDAfpyLCP/YAw128LSpix3ZUM2FP+a4BIjhR5enxYVJDQ171PNfmDlTwQOQ3GEB
Et1Iu4BnXnS50sUHKMLdblJKVYv1emD2dq7mAua5+CFv668htiJDWLZ+sTIKA5pf
vN4WPbiIm/w81HPqhMgDsl/ieRde8md9rhcAWeSrsjwGikWv5Z0lD0djh6AnJRlO
924JR45Vq7UWQ22ksM5zsF0EhVdTWHwCGBzfMNdzadLqVd0baYpaLU7WB48fvja2
+ZXN5V/Q6tnnmeHkTcm7yNvx2rNpbSkEW4M7IBp+yjJeBMwIdVsaURo/i+expjYe
GhoE3gOoBu0HAE9O88+4J03IjvyW7/LHCFYo8HglbG2XFcdM7/bsYMpTwNwMJIQv
dlM5oRI+EXHzhfxvtymGoD4ZIYy81ZHszut0rKLu6lLzy97hrF42ZLjVQC4HehAd
erigQYfG72M+5f3N1++jswW9Mvai6gn9nHXQnqRusVey/AjsiWqAcfDAWSFEUPQd
Fb5wzlVtjF2xxDmTqn+faJpu6MCGpeT/0u0w853AM/B2Ely7qFj955oxduwEfNoO
89bARsxvr6tceft8ordN/zTd3QsnVKleu/Ngripnp3+HvTZD7cA1gPQnAbxCJuiE
eXF2SoaNRyZQNzLxyU7aUqW89sOp8vSa3H0bqLO8KsX9mVw5sDQxy0cx+FE48uWY
PYy0P8N1hq3oB7tP8jZKXduRBR5Qol0/tdLy8IJzI6f7oiA+EcjF6LnwAu73ryo4
vnCNMY7iEKCSZbzW9zjjZF0KjGTf4+3TIifEg0VmM74otNdJS1S5aoH7gR5ZSfyN
reiDO76vnK8N4UJlptNMGrQm+yAQmCmUV42JhzGCyJlafxbmvdFZdUrBPzjeHWyx
41vhHYpi8Os0glXeefR7zbuCTHnflkNMfu7Hd5ubYQ7uNUu2tcHvKK3J18ll4arf
X4cX/WvzxG80MwLNxvXR4NEFCfM3o+XPPcLHbjtn0A1grtqAs/9TcBQ6V1Iv6qbM
TIk5AJ5WSTkRMs5b8xc1LyHy68fu4N5cmFRo1bGosMS67ssxAXp+lg1Av1T1d+lz
tjFHf2U+X68IzULPEff7mMl6tbhPlv58XAkuZo3sz3N7SzLA1EZ0+5cwz8KFXpsT
IIwHuWfnx6CN1Pdjfr+cffaF98Ue/bC0pPODxJMvf0apS+88djzH5jZYQm/SH5Km
GnCNB2RF9OkBeMdpJ2Tx3UQhRXNT+NBIo/7T0st+GwgH1G17s95gUrazHExA52gQ
SOsBG7W0gkciJVQSZ3xqdX/UwiDEpoE5mF0XoLb1FnZDd25wtaQzAtCtwVHNBdl7
WcA0Spac2EBL2576dhTZcKc9qaLO9wpdRD5FTZ4RnXYXhDYUN3ErjUF7yysGe5rK
LwHaZSLkNnAlXjJvr27fuKxTCZbRVG5n4+DNh7veTJx6VjvaT8hLPr/bMjyVu+Db
j2eJkj93DF2tWkX1HsQQLnIL3L9Kdjw0oBnyyVtJi5uNc53wSoRtAEPrRVgS+OcB
Fm7JeaDZQwf+0W0pXzMf19hiZDh68/wVE02orDb+hAwTncJlN2T4Igr6i4pIhEeJ
2oMCK+I+LcjyJ55/J2i1mgeLaR6LypgfrANmqb6JP//0vUAnHb22t1OF6n+8ZS6C
fA7xq5pvpcFiYL/oKMSYL4EFmoFcu/M7LCUVDWyFCNE3umDqf7fglymNuFWaeAm6
TcC6rkfCsr9lVRWkE6aDuEqQNKe2R9LTxdpFPjWAKhyuyizkKO+vTwuhPmZopPaj
Idr+pjQXO5VWAo0Qift7NPkRtY6tR1mGjadJssSMYAr1tk4EUiY8YkSHYa21PE4Q
zvteAD8MbVAjqwWILzoO02hNwiWRipBB0BoD71GdTJsE5S9WyVawRfSoIoB08ovF
yIrI1FKoDDOrRQkeFinpgoqmcaejkyYkKtWQ47jqE98WjfQWI3wmElH1cHOQcCNk
nYD/YY2sxGaqFfdr6IBd2aQQ0u2fpLSM2IJo8mgp0KAZMKagflhT6Gp+OMrdRGT9
kWexvmVST53x+QPVF9aZaI40USpsMdE6nUUh87L6oUxoDWwa+OT59HFW4+9WWls0
PwGRY5l5mCbB8Eu0+GvUWi7iZs1GaByZBmNS/GjYgHPgupQI3etDvb4lbmXp6ZPO
ST/T2jCY8YWd7vAjm3i6K95CblTfC4uNyOsCFRcbSXrUTXwfo+/AdZk4Ld2Zvi3u
2W5g2tKEMpoSSRDiBKA36jeLyc3DTp9DbOuB30ybUtKgBk3TUuCFJmvdb1WaZwQx
20MkoIT+zqa5nOuiBBrAZ0A/VZgH+a08misyMZjHbMwr+P4dE4shdA3NB7foYnqx
lWOYHF4zEuilaEzDL9OVidgm3XaJDLK8V3VBBy2KrE5pqsbPXpXpx0KmcFpxf3Mi
r2ideUonlJSjhkFoDlQGbVQ0Wkm5biZhqrvRC43xFaE1vDppmTAjm1vFEAwYBQ9j
oQ2EgqwJ2gU71wsMi0QuPEYhqEoDA+nKcn8BuhdO5rnWz2Cv4JKh2Rm5boZ8mgVS
/CtFZ2cSJO+V3sgI+Gfc2RTTnZW/NpKVowFj0sQL2vJmXwxQQGVkrKvbcWG4HccF
Bm6DYiDHFj+C5Nj3nBjVl/7NWp93fySufYjygvnGkJ1CmNeSIS0b5qxuyXpc++iA
O1syXKZveDr7c01jk0bcGWtCFYREX4r26yRMcZQsDmlwVE2j5648YfU7mwrPybNY
GsRbpCQqKpOiNAt51sWuS8dcmj7VrMq7RTezpuwctqRkpt7amL/Knq0oj6cVocWb
frjcU8Nbz69Xjxi+mc4q5n7C7/GXa06N5zsjL1SDrvZuYy7iakeU1JEPloMMT7nw
9Jl+IbcPVsAhPxOGXLyRmB/GOWv+qufrCHsomGL9PtrVEQOT0+ree4ZJVJNJitS2
9IL2hTEhX7bB5vKE988u1FvaKxsXMLjAfusF8e7nJsHG1Wi6mBQd1zllU6HPFz1g
mQ4ktT4Pz1/kQQy3hEE9ERbXydmP+Mslnx5slZFoDjp2LoIaNiKnTcPAigpI9dnY
hpbDZdGbCbcbxND+rqMDnaIG7ei1++X3UlUZ6D0rfGxm8lXvGohhxP1tYn2b18PR
Wo6DZrRuyyoO6EM4qX33ke2WNIf5zw54jRiCwtiMGtWMHh4X243Ts7o8ZDLmQF9B
+zd/VWdU8UUoAIXIh7qDxCn//ZxfW1sCnABSLj5PBBGCauNJBtGMvN3HgHeCZHO4
WxnH5x4B2wSaEqfOZDvA5LJUPff0Ga/6EHEcXUUNh3UHdKqrjz4skgv+5OXnjXBe
EKDKVgwBNpd/n23FoJATayOvI3ejbsiRAOhMI/iyJPO/fEzbGbRyh/bimoOIJYJD
QKYgmBHn9SQBhLBhbpqh7xGq2U6smUz1M6dRxpzz71J4wan3DNb582lnjijG4Ant
ikRz42pjMm+HaB55uaZCCYp6NhEjwdHOZQoziNYr2ZLy1egPht2KXu+XNLxItAi5
hcJ/x+nFlJilUEP0CX7URNnVatitGelX74UnnKnlreVRW78qZw22AU4QU7VOECAU
v0Vgqnx6rbuIEA32aJJfRX+N/1GnrdaSQ+QgLySYwsnUNE1JRp7UQGQXBrggMz75
jhOXlHBPoyiqsydKXI8yT819drnmqft3aXYAfwxvhXOrwjgcL8HO8dHRRYsgJQ67
MNp2k9sgYimBpuQYrLVW7d8WiIwbq4bLp+FWRVmwCuasdaBGsYC+spebQbaJMIsy
HSw5kT9pwzKmTlr0Hlg/ObVSVU6ABqMdxo91oiuCWptDomd6s7jmnqL+pwzqMG7V
Oy+VBoZ/5mC1rDLijfRK/kDVQl/NLbY/j6ixB7RRw9GCwxO8+/0wnb1sn8SSenmq
teg7CHpEguYlwLIuJfYwk+UhUznpwG15/nS7+S9TcCrdmyq4xPFHzO9O+Pij1cYr
KYKVPveHxqqyk++7n6B2RGpbePXOjkZloU5NRhdUvbaxCfHSPPfauEVXjiCAYOW1
TT+4jyCxTXzd1uWh7DzfWqaquJlCjceu1nhtvm4v2wsNfco8H40aKLh5y3wvoRJk
0FC4RIm1PdrQ25lrjwAyQt3GCE+S92/4hwJIQmykJMuvrSUez1rlIkawoKyqyurE
Qu/jIbKQtSHOYvmpgL5CjQzKIahu7/BrbpLU6trsHe4pFymEZBXFWcpdmjxn1DGE
5D9u86qF94cAi0hQusHCkTFRoi434zQuB1Ai606G8cDuO6hj2Q1LVr3sQXogDvZ9
0xcUC+j/dBzXDA9c+DNUjqBytSjeUx/BVnFhhwPa9RzmuEwZW71iedU5Bwr+ms3X
QfosD34miw0mcwVWLHmaZ9pjAQnrfyCZoPydax2qIcm6sdCBs0f05sBbvM1qlFIf
mfgi2GsKKOcyvBWnVULQ6KwSikLjrMyLBaTc8tIeoezZWHuWaYg/sH4X3rE26ZP4
tOSAlOWZoV4qGWYgKE8xbQQ2BpMimKHWme+KT5j1Dgq0/yrMmpqvBNsbdU5anzWB
8ScMx2is3zkthEKbLRlcW0hvP5GeWivxmjFcN3mXVNi4hlt/fsRVGXOCJj0+88Hf
3Fo1jQnEqTsqwtuz9Tur3/wHxJSwLV1HNSMg2Dw9XFxoVmfU2441zz0RhrJMVo5o
KYUzUReKb6ef56PqY5/ovJRs/Wn8S37rWrmzRz+jH+uv3q0BPiVxE3pAFPupWCLZ
+rbfKIn7Ob/RqJLwPAdEW4+73TU/eR5UiD+hP6eAVF7EKhTqNNKsmhSMqw9alIF+
kvTLWkR8AMFhCL0SqweZYT/zasC7bbxavcq020Pjx0bK3dWSnQTSh2qwecdG8AMM
S0erbz5mhDkUuy9Vuj5hI3jKRMpeMGjznf4rzVQy6nnClzX/XNrOGDc1uy+sArAi
ea7xX1TGahl8W1Sq+ovAvpA8PWr/rmvKp1S92fUNq7urx0SJCxGZSSTZRAdjvGU9
TydMFgMewrpCafGlRXDbUjriqEcaakFv8xfekF1PZDtSrdRIvxQMtc/wFkPs9j+x
Pdv+YJE/ljb2+MDGlwRmcWdCVZzw9ypgDxTJyo3HG/aBQ1TyNSQ5UdpGApSggCQB
7vs+yP3zSRU0XWlvcUxo1TDOzBWgEfvcepRcEdd3wvdEA/hOeXS+6QBUeOLT62PM
72QA88Ik1FX6Xtl/exXbIInvz34o8vn1gnJ4axsQXdMwZ4qDOOaArHv+VmGlyuqc
1U5khEHPXzyqo2xU4fTRm3aOiElw4zKE7kqPUxliUMbxfgA5nHEqDFeqCRLGRRMe
UJkbqpG71aeE1v3XF9i6D2o4sXG5rJ1KiDWuOT3NxTtXnPCy+wQDOlAoEpmuS4so
TwRZrrxlGHSZ27MG6ioS9F4qDolVexTd6VXHJQf9AsiCSfqw23BgqKBLYNxEdu/h
ocbX5+y998AD9DyUaRj3t+uWG9znmQ689fMMu5ENZu5OojSknbrx+LOBCxR8Fxvy
Imc9QymSLhJ82rXAQsClj6gSmJHhxZ+sji+BY53Sjxadq6swAK2udcGfqVlT+WyN
btdNNA89T+GVuLRB9O+Xfh8sHVMb8/+f3FYYBMKJxZ6vofhpuNApFavcIbhJXzNd
E3N8LjgqXo/2Z3wAle0NdFPISrAh7pSsXqcYHi+smmctN6G2BT+hL4g5AOVcbYzg
wEM1FYMIf8YbDXeQ9ZyDKHUPco04Ery9ZoIn+HJ4SFAFxhX3bA3L+1qvRmqilK3z
PyqhIuX7lJuYZ0h5BxgScOV6Sbj+0FCLx07nMHQwq7yzp1qUcptGEzjAky/+xtHK
wy3dn5NzyKyW11v4eG6ixB85a+h6LETgOiSQTEh+3vuGiqasbNvwQPOZspvBFchP
xeAo1n1U56Gvr2wNKYFThF0A2ANdQYb7dn3GRB+8AVHzhKkWipR9UAE1giPV2Q3N
doVXQuEPAD1bCz0JDaQtGsNInboPahFFjP90IbOYLLET87MJ4mNI+/PPkh03gRII
4JBHy+maIDgzJXMBs1lgzZVFjfF/+xs1i9LDtBij9D4seNDlFwJK7Fjj3e6sDw2u
Mg9pkcvtn9G468joD0ZcMNLmNeJztNZ5v+LGvNHmIkR3EHy/uwMJZWVJk8l/p0vz
SCbCV+2qCeoVNKHyatvbOJsX7rGYU4pmCfPlunbixih+8hGfBUy5PqwtVmi7AXNB
peQXyEF2SxL1z2gikHPjlnNYPKyEhm8ld/+HV24HkIcaPL6C5KutRn0uYCJ7Gxwc
4CuO3KzzrvBUeZCYWUq9SiWP3CzUBbJAA784uwIRXfZU6zn3Q38KHH2+EpJ4AV0N
qWUEh1mUErpWTBcWhK3nyv+4kWwrf+5RNBQdyj/qAemRQXeM0fFPLi33g2C6m6JU
t+Byf8WMjld0Bdxv+eA+gAvtaoVxPDiZlkYkNAOVESatui0C6BB9RwaHlUQLV7UX
bb7irHYWc5j+7zSdCno0ytrgRo0dXz8hM3waO/ZoegJ83KqLYc0Rpzcg8sj7IvEj
VGz7i95dOWRCjLThMYaIFOqz5CUprsHJfBXBc1mTSC/68M/AtYE14LvdMHRmGlBB
T8eU5npCGoAZeQB0FP8YHrarDOhxvm44e2+SyTfarEQgKSgbEQe4hWeN5Wk9+Ozg
FaaUCa8W2bKVUOoA8oK9/+05UBVCq9RGmVFAyM7GikWzGZNQ2NhtIlqIE1YFxiV+
XvyFcyyqbL5JxrZCVRbPPY9IfyZw29PtJKqH8m6pSkZjmOs0pG7hUAoM/tYO/8TY
S5lpheBfZyIGlNi6pq3q4MEUUMbvXVOuOVKSu3KI/kbFwSRMB7RJB5VYljuRfkcU
/OeHYwdq2Qmwqw2yr4ddbWmqpmN633KNVEXyC/yVAU2xbyc0J2A0g5vjHo6JfKuE
lHZ7xB1GcKu4U5Vwq/qqIdUX5iaNW9Obp90wByxBBKs2Ctm6icKESahuFYLB06BN
i8Ujd1ozPAvGcvNGyxe8AD4JOEGeb8RJY6MV+P6Fr+twSsFE9KptLGAvxWbsqKMP
8u2QpttIfsgfwedcTqLdPtlv6DT/J8MQOd3UOTvSS2tSf3c4h5T3dEj/7USe+ULw
H12Qmm/PFAsdQK2+Goy1Fsu7TrXfEcC3t5kLSW9AQxwVY0iCc2NdFlk7mnUy/XAk
cL55huBUEDyTRzN5L/MG4QtUA3as+0OdIkf9c9i+dBZfNPwd6Ob3D7nvzBoflWp9
NG/zjWRmwMqhFXrfWwSgY7Ts2OxKZAYK2Zv0HH1AT2t/qvlVxlnETk+TYIabwMVw
dSOiR2hFMsGhHanCN7oZUz3TH21qO2koDsm8YMd1V8o/0HUj7t3hBKTGWuLW/a6T
w1J0OHZXvKBYwJBqiKmvUeh+jk3Vfc4FOxZCC2U76ZiCDMLS/6YTEtchaVxc4TFk
AD3FtSQaVqgwxghTbb2Cf+bPMp953LGSmHCfSZbVr+3XRJ2gwTcXHFjZZgI9kD86
D2FWg70WwwGng+pe91v26jHq7TD1dUhhX00DY3SCJP06EvCieKA13edi8t1/cF2d
l7oKW3J5gclGMd0SPwnTIGM7E+2ek4ac2xl4dhVw87NNjKWckeAP+u+48MInJbgL
TGzwUaeLPJ2vqybhBlISy3+p9t5W2ibcZwtBP/RxGudJJVqi/jlVe69kAqbgU+QP
GbA7hyGMmT6Jm8D1EGgVT7+2R1Y4NbT9MucMvA6N9JgV8xQzuokFJ3qKs0gRKUHi
M2yYG1VO0fmrs0N9RbGGHoLtntztrc8ZLO33EiBi1iSddHEYR7m3ulycI26K+kh9
aVMlpg65DGIGaCru4d8L7wMIUR6W+PhguXHFnjh+Oc0gzecMeWVPkIOOUDzotv5i
Uzx+QT10yfIpms75xHUzzn/5w2Ry/nwva3f61vVwUVL0nrYH38haLEE5kOsw12a7
6Cqh7Q/OyETbAC6BqYaTSvV3sSpAcbxteIn71+JONTg3lZWZCN1Txtg/T5iLDe8T
PLCWJWL81FuXf2g4iwymJ9B0bWjvWnvlmubYiyGhIN4PpUmMove6IeF4RvllZdXv
QUczV/aymhmzdDdYddpGy//KqqWlYPYjaswjDjipUrFoLxkbi3rIbUgZ18P5l/ng
x+NWYbaSQVAGkAsIxN+XTZQRosPICXHjGxNmYWgATc1TUSumQEDta0q/oE1l8n77
skQJXedxBPzdZaYyv0uR9AohKpYZlIVa4rQ8OGhCOgQLzC9kn5QExyabnXdw/giH
Lrq2t9C7Z0yufFnXjdHhLHbFXTEIU4OCD7BUGLidxLzh0grQd4Ni2xECRVSAXQtD
Yp16D511pP1q2NlDc/JhgQ9He65bqn1T4s8rq/Wjy2CX8CUhPBaD6RBT7J+iVeBk
Y26nVfJPDa+DOQjHe5Tw+T3G/mulKbTTa1vBFXUQ6wLar+JM3MzV93ciHTnvaQN2
tz+IAHGt3crGceGDe89A7v6L1It9WtfMA7xmw/Z4JfzBIf4Ki63ZY833APIrcZpZ
VOphkc2xwRE99XaLq1FYoRwrxlqOBg7xf9PNKlzwtanCGRFL+ktEL57WhRykdlPa
vCBVZFpNiQUM1NoPiXxAJDUAJuGoHl+QOOAPwwx2pxrGYoI8djZl8b9KzeKm2O4t
zxaHOtUkU9G0c+RAJdFUzAqXMDKaVRpLev+ndeE9ThId09DMl9ln0y32vtcB39jP
C3c5F+XHjednoNr6he7neuQgTo/xMbhdSaEmRyUn0IemvsOiN8ImW3mbaJUo91bc
eR+1xY8YbHKVY7EBbssfOoT1oLiwynMMhvkl31sHUo7gg0DmaS6ZSk3njyaG0pwU
YLHPS+8L0i+jX/yrknpWR3A9RwFHlBkx6v3xBE2sb4bXWrgBaoswSMzUWGTDUBnL
ug52g1ovK+4/5pDKGdWuOGLko+HjNmbLgO95abaeERNgSlQduhT71qKhf3KBtSX1
GzRbvGcAngSjHeNH75F0RIAyG1TT7T6rSe09SPGbWCBf1Xlg4S4drX93JlARl47x
iwYZVM1Nmg+XePeVeZOksegH9Gm4KWHoUF4pFfKi8O9+LYL5u9M+iFYeUWXNguLk
wxKcRw2YwlGuXOx7BKCdlu2Ic+BmxNeXLmhnyG8cwPxv17jmWZ0foB1h8uMoFRt0
ls+CqMxBcUyMytpU5wjSNhcYiCKZeS/7W8HgNi+58jJbnOa59PG9HAoz7ZCQB8Fq
9VVlp/lmQTxZSEdQwPQ0Hpd9Gr1uGqqi2564lKMgDBmMoZb59au+/9uta8NqGDhF
ilRWOvzCyiaGyfPhxxPMiOVCIGXHHwpnD9Q7w1/8CiOPrZBOW4tkFSHs5sN+zVdn
mOcpgBfVzHfUwCSKA2UuZPvyxOEWMvDlwUditFpP/JsXJsD2HGiCUskFfs1lq//r
0w768HUNaJtF+1/UrhnAim+oI+Z9YyngLu+w1w7EYQd3ElxO1Dpzp9qIrqTSK60X
zL4+/+anmekPff0y1tByBT1ugEVa01XRoX8ZppOIyyxCZ4Ck691jVy0JQBPT20ka
CW4zU5b0bqosA/3Qtg+oh0gjytOFyZIx11iWU4O5j8QLDVALdFOzunPNvOTZo7Hf
tTGyzV0jF7D1Ptho30b/a48g5V7HlUpzRoCkewrL7dbw59MTL7bdxjgiSL1e3UFW
i6lQHPOWi697G9BrqpsBELR1lflDsWTOXORatnpEey69ZvAqehsvpa8Tz5UQcU63
EIsb3abrOZBwbjmU4KEJ3U/d+jtEXmrS3bFt6BWMx5lMY+Q3bszjOCLnQXqS8ZL6
CGtQnge0X/CUgEd1SGy2HmD+sXq4ugvVLj075w9Lq34ZKoGDkp09G8s6Zo4PKiWh
eVaYedbhnqj47e3gOlNGWJtRsKc85kw6UjxBnDsTUZf+fmE2jWuKcYmHnmwzXd3I
irGdIS6UNLfqckhEePZIaTXFSiF/N+tiKePZJf7AHMSjrCsA4w9nSwbztsUxgPkq
1jLqegC+WDFjkYFjkCztn+k95KBcriMcBXqdbzmt+RA1Vk0TKfonrIXRwiDzumwu
3A5LR53za9VPOexc3+tGE3gerTY7LlQqaPR8t4aXXGGfcLTba/ILc6N8Qz0OG929
34WehLBrOy7tN2oLl2OiYJ8qieBURPxYTuBnIoFicB2+n0JFUxC5tv3XLvmdnhhE
2ozZy1Pi23SMC7LzeiApng/zmhhAUXfbGMSrk2I/pJqBGWShckZPD7ia2Gg2bqfJ
ji/REJFcNLnArsHv47FdmiOm6n1Z3RmHp25jwDgNlJAccNGAPh7G/SNtxXsG4AQ3
sapezxc9BP8LHx5agKKyFe7+VYasB+Dqer20ASgL2IouevSpi3+YxBsi8/8NBDUX
1TaqQkWlQyotd18VTqJCnixeAm2HYel5vQsVbRSbS30SU84RiqhMdggFYNPr3Nj2
I5R/Tx/h3+NQO3W/djuLZMLSsdTgv1hU+2wMLuhsUFMEr4HjXAT8EY3jzYlFmFYK
YwZnQunIZazuB/HEfxxMRxY++k/dr2G3ofeZkpQyPB70oDPL2SQnUotAhvMrxVHv
cq11RH98Jl3n5hhlfAbspJb6V55UwgTSDijHr/cS4MujT3VUkAmVBd7rZ7bJrJlQ
9tPOqaEKeZ03ZJstvD5vsIdBtrF7AduKZfSgrGeiUFHC6SuyeSPLCCxgk0IUBY5g
s4IdHtKB24KywWAY6jqwuJg8XbxRWvDRRNLOq1hEdFrY5GQPCKKI6nroQGuD3Bze
lJ6GQz3i6Ou7K2XrrGmcjs5BSntXu+GfyU/2EGEC57kZQjaZ4yKZxZ1R9R4/+wXG
lkZUkgZQ3/E/zpEoYssUL7NDSyIrfGuq6kTXDKIOuYipzojLUf70wpc+ZBQccY9g
J51z9DJCC0v3QEpZ6+gBO3rkW/7uB7jMZggEB8IqUX6gqTcIR8nDxa7qHhSzfK0e
iHWmbDMnYNrX6Hs50gM5i3D7h9oAoP4gZXufd9+1SJN2TRxHrWYEVfRzJ+/t2mfA
S9hhazG3WGVipb/dABBd0sn5PZJY6jf+afSRgfejsG5op3IzWoqQbRM5U2x2N3bI
CCTh4nDzjjghRFl8FMJr+2eEiIEKgCaIugx6gPpY6oBlbDJOvNd+L7i/suNiesm6
L/IlnN76A6K7DWRYxINEhz6DtE0Hc7GEiQxC+lHO+ZL9qJI4xfBZ2NAwXRwR/3Oz
LdN3Vy598oG0He+TFa6M8hxjxGA5bTn0rljI9WxYDXDF79qH8Uzm5NOQWOi17aae
pzziB7x2Q5qtNyhBIg4Cl/H3OmiV1SSORE/z+biuPjtLaERUIws5Rq9Tybl7lTe8
HFo6H0cY4YVHJp7s4txEkMJ956agXiwCKH1zEw99MrvPqXgv494oagohgJGcaVrk
WN/MBjZczkOaIucoRQjkLqRY/dfYiBfAtyX/CJ5TOLEd8zMz0Gb4RMglbVgxiPKz
SiF3mBl/afBY4qJRzq7YBYd8wROGSEz9QehXZ70i4J1JEnpBXxALEaRjZgpOzSgB
8Yb1Evgwm1i+HspiUhk6Rh/Rp0u1ktK1Uph6rHR02P3E++5g7BwDtu8cBIFWezGB
DJHYCkfDe3C+nKTQeVEFOsM1U4yr7xiemfgpQJ8tDZL0fM6hZo8k8/KBw6R4Pbm3
xULzr0v3KV3ARUDW7qZjWmyxtJAsCJtnyFevh2I3LQ69rU0PrVTp7gN/xhRxalQ6
zOTGN/7YTJsByvmdcYnJj25qjv+mJ5DjrdRgLtX1I+qD4INAUAqJyN+uhTsZpBhA
Msm9ivbA9kmDPi8sc7U9hzLRcJyTQBiyIHWSYMwvn7pFX/6T4v236fnCXWMPzxE2
nZmvMo/DVoL0TcpPqmVtRC7xtERBp9Ym257ih5VY7+QV2KIlcSiZPdYHvYV7efKM
qjJYrNIgLdClID97goWemwUZ137iIQxgy+Bk6OszxGtF+ayHg6Rh3th6Onb3v7pM
pBoCqfGxs52lg2qiX2OSL6nIQeZ080h/mO/WWYAsOT0Hk9wsnOu6YkETVEtdsbEp
t2UP1rZpK0ucaDSF/pOirH5+NHFg173AS+LFjQehj6FCfUighVqd/Ee5iUYc54Bj
wMHISg1uiEiAJOCujufw8QU9JJIJNE2BmJkf/wl60OFHQsMy/Fa6g8ohMBsdM+bg
Q1xB8j9Tz7hBtczdmTKw/1ed3NqlW4pB2V/ukckgMukVnwgmd4+2K06D9YHhhN49
6XMt/PNuyUFOV9SEIhJwY4+o0xoIbfcU6jgC8RClsHb3U2BHju9ZrYr1c+an2tup
CflGqNWtd8UCJ/OAmAax7lgHO6P0PgUmOhvy8EBvXB4q3yG5IFXn3+wwEIee5nNj
LBZBMBt3WZByuSQCyrFwtF1J5W/Y+it5oNTQ3ITeD9nTAUatifxQetylDaSmy0aW
uAI0LDcfPsDnVU+cxgT4AD6YhZRSU3+gE6Mg/ZpzdV47qmUWyBvqTmbfPL0Vk4/u
lnE1rid3cjhIrKBAGV0bOcYX3faj6xa8mwBfbI3TUtv2wpd6qAbPzBYrrX5qNNR3
2+kZZ0XEbdma8LdKXh0R9D1wbgywLP04SamXw671nY9sQwLbU61/lL1eviFrDcqd
VhXC+jrqJVb1Q1Z47pWPFEv8Kluz2gRAI88Ni4v4EizMT9K9eDXK1c4aPY4cC/OM
vn0YpRMi9h/RUfExg91SO4xilCmkvhhfVGNiC2iF+9Hh6papoEGSqrTJQXgbqFY8
NsKdbsYeGYQR1Qnwsr+XSoasuCQRUeNo/of/i3A+DqVzJpB2x/iAwo6D72p12QFL
lflRMm8HrJA+JVIUaXCbKMv2VX4bJ+JF1hBuUEBhoi3kYkbzIRT5d8vkjcykIeBx
d4A8P9/wJnbr2dRPaLcGkmvz5ie34//PPfcUD7+oylMIHZqcSRKu+W6xQAsgU6F7
IoPMic9CPhunvczI9P1WdeAfV8+e/hr5URpOJOsJqIl1vVGqPM5KrRxYfhrxAFPC
JNGCTJLUrthyZnRIPO7f3qlYcBlvQJcSH20kYWv9zOizq91ZZXLv+vbq+8NTRHTs
gZGudo+bgQeiBYRg/WRM5aCYdDcVoqwWPF+DM4109mg7+bbeo2mJuWZJvPyK8ulc
Irg8if3z4LWhI3WrbO6sHWANJxTTkFg885f/Z1mquBrcrooiiiMhKG5HPz7MGsTx
24DtzYIHWWLtlq3G4waWK4/OdNBZtvSKPnIA1S0kGNoCtl3zk9beTqrijqJt1H5g
BF2nCtYOryfExE5uG6IjUND7w8h415XGzC9/DqWPEWESmSv2f2kEFa7hL0ydawAX
ZCF0TWLQeMFkeA6jMVCmIkKH++tTXATkopDiIW1HrgkL94flgmMcJQ0oweaPPqK+
lcVSl1dc2qLOIMOxLzohiZRbMltIcwG0pOI0kNvwcRVT4CKV2hLfUimWvzXT9/AW
8ONfKFYeswMPFQMwjTanFihKLmVWPWG4VDmIymfRgL6OnKf7Nr/P6EPf2aUcu1Q6
0Hf4EYxucOsXstFknuayAw0Oq6hFZtnwEdDjQ218akO6gyJyMg/btw3ITMgQScK/
Y7qSq0b0oDGWRBrw2aqTZ6UZ+W1lzywLICYbeGlHMlhDDFfIeGPq+dh0ogetEkK2
AuqN5ipagpe+Ifcgq54RamjRUl4wx07vHyzVWvYZT7tYxb7vzaMmQ5VLufQ5iUok
89U+yEA2YZ14OCM1UQ3TL22tIHWzSPSDQuFVFXfVTjzQui+gtfJXOOmTOydshklN
cPbgJS01z4cSvLSERczWrNlABXlkxU4x5r8lL59z7V1RNzL13JV/OpsUl1YyGo1p
wbTyolTkCangMyABAFaNzIbFH9n0TDR7WmPRLUsfRfegqdylgSb2s90Qh89BlwGY
anKORhjzWDRW0dtMWdeixf/GLpO2k1glrk0sr1aYPXZZjPlCRGaRvy256C8Ao42k
QMGCR4XiVywSwgRJhPe8L9lJMDldL79mBHXh3ckWuJyk1HgbBbzRjdXEm42g+F4q
fxNMvKgP+PVYyDpTnTt5ujyfczEEaxtulX0grFajZeDMgtA1Dlf/4JYWWAjfqKd7
3HUHGCV2yYaGVR+GEiTfH5Kr05QheRb14nYmmgjiCTyg7oZuy9wUagDlTq1tM0tt
HiFlUP2OJ9ROrd3WJ8wOaWxzn/d3f2rcVUfeackz3zfpNMoW/RMXAsIfR/3ul5tX
n4oHi7YzGigqf0U+ec3p6tFWCy0zn2YkAc4vp/E78DObY/SinQKKR7hCeuRbrUZx
40hGmMVGEf9XxYOSDgGkptu980e4DLQ0T+Z1zdr1xicpGVkeI+3uKHSkVe+pBZdE
87C4vkzzUmqLWA8ZFl4RVwR8NgdCMwap+H4T1UzFA0U0ygK+Mk68XX+dbCzAZ/Ym
DUtKBzawr4AAl7QPvGrlkeZ7dTSVi2T1nkvcZ9hjFHvVIYRWJEE46izlfcp6Xu/v
D0zeSCQ1LXyY9t9d/RoDUHXdVmdum/7ChfTZkWfSmw8Gu24/lh8+plzx63WVChrW
KAgvNDr2wiW5QyMwEaC8Tuy+LpL5WFEcyC+hJUsSpvjM93W7EQy7jxSlz+kc2rcG
vBvURB2F8jetBOFxJMKZBDV3rOyd9tvZL4Fzw6QlXwi2Kq2OJXhEGksMW6C2jM5B
TRJn7Qvoal6qJxpKYZSIRHmvcjFxEVkZLolkHU8JB/zESmuSEFHMN01cOevPDMID
CxS78NN93r/n5OoHb9cdp/Qx9ZOaMsuhLmPuI1p791zWJOgL2eBvI4gN7Ysi2/sb
bGGMnjrgTu/n55vmTXKF0CYfZWQ49vxJwfUI6XOmMR6P+fRkeA7TiRRVDo8bpmuu
aMXLj3cwoHKiXjew1kEeaZPT/d7vnRM4Z+8Us9H17Q0hRTSw+uByrcopLRJjLSg4
yEbpEO2YqBLetsHoUX+Qa+7MZ3/ULkiCiakkT4e7qJlgIAuGk0/qeaCul1YuNOTV
eFNFQC6u3UIqwJhDHaijOi9XcexD8DGeGN2TkhblX1bpCbw6xoabw3lT0jtdE3P8
hnVvOA8nfnASDIcQuCJBovGNbaGcOMgxYC8ByjYMYUEpZeApKk4NjipMgh4oFoc4
QNuLMUbY33KMx0lcOcyiAhFKMqnimdVZL62VhThYJw9nRMozT5Js3kRSPjnKD7kY
coWlM9ZY+FS2yQ6VXDLaA84H1hNGu72MvpOSixyCvf4EFGnUv/z6yXwYAdRSvrtW
1Ks8y4oS2J/NRtrAfXVN33Q6b26jsJJhh1TdQzLq8XR2yyvv4mbvAZb2MtCqPWsR
3OcTk7lhB+i9IFU5tH0NfccknLfE+X/X3ShAkzjtA9S/9sSBfe/IGZ073E5kinzb
CKtRbnYj8dncz7wSiJgTVfW1KZzj14Hs3QY/VLl+CWBQL2hHKPlgETNyzZczyZDq
XS6SyxjQw30CggK354btXINUV9YuBM8VqqUrZdSgqi+YY/I9H9UgSiT+EtE32Ibt
v6At7OhKJODofHuGi3kOFXDz/g97bGb25e3NUkneUkI23lOWRmSr1+yt/i1r9hov
hl4Df/HbJHTtd0Id1bULsvkOLkY9Db9BNcLd/j013Ge3gbjO2BFoTuX3VCCPvcvz
8yj6J/HcIQIJjWANvab8FmZZhu1tvhL/EV2nnko5wfRegAxqGDUek3lJP0DENEyi
2bYduFG7jz8MiiSaV6w2kPMm0J2C0lAuZ5BH/5qXJnzrL/ezMnR5Gzs7zLekBzCe
M4pYctA3Z6d8nWVLDQ+ZufpNkq2xSyAikQrM9m+GCu8pDATzqWjZqqktH1gtWB2G
D26LZB4fOHTmrdpTUFXVFr9SkgoI9FS68DgWY7pvMK7Ks04diou90U/WC0coumsX
y1URkjUX1jXv9DKt7Xx9RV/0PlK5gPLS3zHlE4gCq2wb+K+TxUG6XWxUuUNBJ+Xu
d9r7Es/lcCXlL17lZB/T6ENl+qoXeWUWR4JA+IypDARHHNAa+jEBFl5zeDlNrgmg
B3zwrVaJjP3T49HTuw32caVVNtsx27g/qQkdGPpoA/NBeZzrAdDXjITYlmesJkmy
mDm0JI4OJr3CHo4sAdlMrdL7epodzMR+9IwnYTBVtkCANdTKfkrA80wOqaf+jKYI
64H4oILRGzfs4ZcC8rQ/QTxQRb6hty32AaVV0MSRB2+2tQPMl4qv/F/oU3HjFI1M
GtKgUNGQwG1rwtC1B2do2z5jLq3oG16LElxPVtd8ppXFq57W9AgkRdj2rwu5MLdx
4m1+W6odxCLWMRtq/+aakE0oKJny8WV72rDelh9lPTXWzg2LBOsIPhzd6LWANazR
K1KBQecglyAYxSLzwxFOce/tcUFAd7mSs3UymMjgU1EZFcZJiX71+TwH+b3+Nv1p
vn0hZZ6M1YNVyGq/oArGqueq38IZATmCrqXmTVOBSGTnjaBXYnMNK9YidkPyFLV0
fCeM/rPHlA9QLoMOdke4fh9pxf5akqiXwKIqUJY7XD/UT+q9skESUwJbl4O4Jqsd
opJRP7PFtDmfYpIZ/BmayZqPENxU1jBK24Hp/KcxQBPplxXeoPowx/GLUJw7mpvB
jNVxdau+buICvetSlg3+h9oo3IAfZL6KlNL5APYdvjUEsoRmXNrSDC7L3K3j3nBO
t2JjmHbe6B4fBUpLwctuQCc03gNuoY6qE7BPTOMwxijbjAvV5Upou4YAGIuq/Iax
jMuY0p+7Zr5/625WHQ9IxqLDHhq30vrCLKpCSfFOvOlz6gNkhI0Nd/7ZWRhuxa9K
zH/JxfN6rXLzNZNIbohPnBA81rss7umqTUsC9+325WWwKOqaAxdulFFR3nQpZH7Z
3hxmVtN7pPLxV6LQDofI6Kc2sS3acPVVyLORZDKWAoEYwbM4EdOvy22AU8izDESP
wX7jK+gVRf+tUsszOHpJBSMvjV9ojznuQgIHy0+qRRnOrE4dWFX4BoK6+BtP9207
h1d25xPjDHADwgPdzoPNtenlUq5CkdBAJJq2Cfflf5fb7OxprT96q+f6zuXBZ38Z
yJTtrZ+nnSoSCTwYEh8VWiP7GC0XISbWcjObNtOcviuvpl2V8KzRcobwYa1PNpmo
hEm6RJyEHlqvTVO/ZNDke9JzJ4cU18rZU1F0UaHtLlilOvW5CnjI0SroT5yRKsbF
yYW/tb9Ko2hLZhoZ1OZLzSlSQrbM6DasGcuTT/rpP9WRjKvRRPmUcTRanIPfthUc
CpZhBkhrxB/zP9pOPs/EgmOoTEVxh4wQ/V9lNCFpVYPKrKbwmDbOJMAXYrEg4r/W
XUKq2hjPlBUqYaS/fyKT4Fwfz/mYr92CLbdOmWZEBpPd3WEdhl0rI00kFz3cRUzy
yWNuUDq9jFA++Z2vWpzA6EuD6/RPT2hbSF5fhwlud6A8GwIbw9r/RZc0lHMBbWgS
I07oT7Xuxz3rmaIy52pziXeLigbXPrV/Nltuw4ZA35V4HU9D9Z4hPkb/bejB2pE6
xN1JwGVrOFGvPBsjqVAssLNBe3G5ecwOQqtKhVJg5Ldpfn80eYe92/WH5yqSNn2l
PZdn4ouh2twd7PcFMXcJ907drojELCZT7BBF6ZSoX+AIjKtS6T7/dqXfXQvrUBUE
+5NdyeO0MGXoIDS572hRN8P1+/eOryyIF8z93DF6sia24YRQtc9/DhhGQAKzMZR+
w5lIzd93mRAax7dw66MU7h/yCKHhqcOQWsNF1Cmm/JTdV5P4ul6Uf2VJllUKyNrD
4H5/7WW6IeKb4SBL9F8eWhC76ehc4nSjVBTmOdeiSSqJMYpEBztR/PZCBEqXyMfy
xK6Gd60Lk7IYjmsR/MDq7f0OQY9oTiQg/KBU87hJgvMZi62YM+/f9pnKhHKVqhO1
Bu9hA/xorOi+ROnfcT7kqrAW3Ind6WdHkY/+sQMWsQEETPiGdNGKkB4neSQJCeIg
y/MWGlH2J5IXRX+bqXLmOFsO60x5z7Ys2UvHwetUuiJ9gMKq3DGVQpYzmcsgz1vX
aBG4mvEAAzB/YvTb4x/jaPcNR2Mi7Qnjs9QNzw6ityZXhFlmz5V8nBdd4iasd5lC
G71i/y/9kkZ1sIa9xVc825BPHawIA8msjPRQdR9VVOTnAwfgy4wd43/YS9BTy0gC
r0tj/BQorSS8CBNCHuahb9/rBH8kywgEypl7ZF7VrQEOJiHX+iBuYdKHQ7ahK/ku
BS9qU36v6JCgYxKW7zDJ50BbttUMx4lv7r4pn1rw8J1376Qi+CYZljlksUyA66dU
gNhsR4zV3D5Q/FGl6r9iKWtxXU86zdt+9MtV6Kbpk2ARcXSAXlTrcGACvrs2N1zH
75Z/8per3Wb34yueiwct/DJPbVpOrWSVjKH3FMLUhvRrnEkwYeBAkFyUYIKQY/Ev
PLvUvse04UJKIb6SAiO2ZZkUAw96iuBGrOfVFip8GmYAGcOdnQw86AsCumcelxb+
K8HM9zWfGA2MBJpbtJX+Wc0f94O9vluGKmfAMWidX9p+nLzFiB32XMJ90b823w0H
6EtLSU07NDpAEd9fdtkXJrlGdzHY2ijOzi1lSq8z+BVHUUZdbRG66KxsUGvjGYDQ
2YjCTZUSZpoEJTYeTLLcMe00Ab4uOLdvmZKlkl7+gAtdTboJ9QIerHyDcz34X/ZR
OeXVSyRrXdlLVHN6D0vRIWSJ7Mau/xWNXKX+5m7DHgHhDLkQBxmSiXFkjxkBX63z
a2QDIS/1UUNccKPEzsseA43ZdA0XPRgBkYvD+M7sUn6WGHVUNJy7ZQDGOtJR9yG0
hVgZ8X0m/T/lyryQryGzwCguXY0oxAg4l6rnNkVjcFJohsnFh8jsKlMtyWDMvlf+
1FuFRkuOQL3KiJKnvqe27pWuYhNva4iVqM4POd4EHNeu+cGObvkGN+76VOK1qfjC
DBddYeQH/XBKWV7EoaYrxuXgR8sy2nwG7C3NxE9yXmT4lwJEAN4d6LYlgRAsssJH
lDC69qV0aJ0hGH6r9RpOg6KpY5325uJiax/MuvW35yYm/bm618yEAUGhjWcVCCG6
39NlIqGoG/9OeXZW8wbmsPMx/CpzxCYcKtyuZ8aY6NW9EX5+noAMs46QHwvDVWHG
x4gzOKHQPla+zqkfC7yBF3fpS1087ZC0IAmrD4tpUCKw9h2udIt4Kg2uQy48dxIY
iY9oAG44J6e2SlhFZm4HnrLjAnzySIavdu9gSul7TVVWDGmDOX8TDKO6FWY6JFkR
D4/cZvyq2qTp5CeW/48Q/rm572H8Rr7LEhBpM77d4pb2VzHJ4mNJMyvfTI4c9fQv
h29bqglXauyrg4d9iAgMZ+otreUstOydV17nA+uiAlfwHH+yI0Xyt3tENK9dn4pf
+ocGpb5IX4q/forW9esswf5gO+CcNXcX0pNd5PAK4oH2MsQNV4s/OWVo0ouvp+nk
lYYnxnQPVaoMkZmlX90UG65K0FnBE8r8GCslIRXsRHWK4Eu5p3qgQfDY7lKvwqkr
AtCMrkzz0QhJMzWSXRjLOeRKJYAjrY4IP9JDYBSXkVyUjmIZPZRjumes1SW1dZec
oe+X9U5pHCdIp4i3fDizeRjeFshhe/OTIihfikZVBzJLRTccbb1pJKp6VwMunySp
yXrKrWKlYKgL07zejBRnV9F0bjaUFNcfG/g45EORhr/qXaMUflckRStk5J1kZaF2
tgISGpqsm7PEfcTmHyG5EU1p6swQ08fLu250QIXkKviQaW6qY5XbVoKYexXihe87
ec4kxqumc6fRTdMy4SJNuKqE7nwNXXutdDgtVrMXNTyyoitbepQNsjBRA5YPogX0
2uMMaLqo0mgaz6h7eik8zAi2lBoTKeYD5EGxDa0p28dTGKrQw+kCyxJlLaJsSlDr
zi5bc8uJbn8syayVbJsOHYiw16GbEUuN8/6GlmXLb8xkGfpcxr1hP0jOSRYaALsT
Gll96wdAr2QyfyqEelkVH9TNuR3ybjvSQ7m/Bw+USRFgxnG14mfhxnMU68J7uZAz
mmw3Ao5qw+1xRvC6s4tZMdC/twbJJuaRerpM6akaaaBV5IjIE2Osbm+ee2NT6f8y
k4UTRvH0FjU656ZQUfRY1Xb1mcmXHw4kUJe8uiilKGrVaN4ejUMnKl5YIz9Spuhx
1QTT47u1f2Vf34g6CE49yAikAyrRcG4sI2TMc6tZcyXMOQTfsgupdk6QGq01Ww7K
VXc8QLXId5gPTlVWZ3NhWEfch2oSA3wcvEzmhhe8jzQtLjeh/B2W3P2eEu70ey1X
r6l/qkASwPan9/dQtnsSPFW2nal7guEjAk0sH84Egz8MNAyb1Z4+kCUZm+s+iAX1
AkX/QxyS0iqA69i1jWKt3PfVyejkrbOATeWhqTYgISuK3ksWoDDvqN9RKMIFJJ4m
ceD8z13NWKPaM58qJ86pHRb272Nfe/UB3DWj6I3G5iiVPywMe5WjfHhIoAVIB+S/
A53IeNdVMI2M+HahsQJUp5AIJ58Fw/PwAMkgesrskDLqK6ZTYHgoqt/SmC9g60nB
nu+cdrbToeL7DoCAxU/IS9maiyQCnudVS1nd9AuONSDc8FeCZNFhhZyJlTXwT5E3
ogHvhz/KVai2uio4C0pxb109OeI+igWKr59sJJqq6byyw0R38PG+5DrXHaWGBTzg
fFZttkQnL9zDti2kpGUf13JgnxfhUJHajoLA/CDvLW5LDzfDFaWeb8ZGUxZzqgWr
T5t8qsyKcgQhOkWIdUniIMdQtZQSn6YHVzgYKGfdTvQ6TyqT0qUSyqIY/K5aTV+1
pGpVTE9rxrfq+opgjhYlBhugUrtpnpHQmsCt5L7cMLtQLPbzSj1mBArTwSsOb5c0
oqi8EjYu5AVBO1fLHG/gqyPwcl7mD0yQOf0Is2NtylOGoHt/Oxcil/RByneTG2dY
wezJKzZQ6AkVmcfkv3kqjRsj3P885lEPtiJ9tm6eg+gco2U6IgsEuzgr0wJb636l
xLuGoLOluFepRG3m5xvVrMrhXIFEpouf6sxkdrykxjzG2fOEv+vaHzaKjxNKazr+
rq0Ndr0KQQhzEmWWBaJEkKWHgDpfBeitscbE7qKCw6+f6uTJhvdAZmvpMRMUgXat
w2T6VfTR8PZ2/JCyATdSMkKesfzmi+avWCdMIUx4aezwhKopoxOfjqnBA8xO4D0T
Wdk24q7a9LRK/1SqoDtFX0uCam7LSkcD2nOttiddan9vLl30dpe23tlWybc4iOsQ
MyRZnsUf9r4zeO9NNm0SufKBnL+NFtfJW22+5Bez24hd5gezqyAHCf0ygoeip0/m
nXWS1NZDNebOoDgWcEMo+/zgBdT8iUqwMnIQuivALhIN0EUJxHOrH1S+q9f+/2uK
eeMEgMl7j27YO0AntGM/1Ht1O0EeLCaIZvjqt9/lFCawKk1UUME7SW1pswPL1Cc/
5srRc6yoDW4YZQxWIYxMnwq6mRCXzgv11RSxyNgXX9t3O3eq8rwV6LT+m4PiMz3B
nxS9YXC1QnxUsX/1d+1hR+Q4wpmrOqIaIn1XhcZ+KEE5pJXY94wKEqCESYi+WMKT
g3PkgaQay2DiHk4l8VA1kCBXlWsxSups+oUSc8nXJQ8ehmm9jI/nVYh7WcyWEH0n
pOCavSjgmWE6nIPMZ1PA9ZXgP0lAAfWC4pXYq6LbiRNCswoJ2axPQ4ZpU5c7iwSh
rV6DfGYKLh5QYCS7wDnU5/ZUoR+IiaAGreHVZgdN2YBPb7VbJ5lL6FZ4WLgKElmv
a1cQeh91K2+G9zvNx1bBG65ky/LtaTprzT+5iolmMwfSHv4bdiCMigeozKbUs79P
WlAEhRyzUzzQzIv3dI4E/jK58MpqgMEPFmyPuu0tWqSsiZ8LEhGUIy+3/bSktaak
gWylWOsVCRyw7QfOBFuHdgPLHDljWy/0muBZ4SVL/M41KSEnMXYKCh1iYPJ68M77
wbXxBECZ37winaJsMMNTUoWWzuBXjk47fFtINvc3U8TA7U/winqRS5MTdptr7GSA
ODJC627miy2J3FsFCbiUmY/EF1lI8olsL7qwQzzHFpw2iKmqoWe4L8cdMqSN7qfM
B0lpJnzaoxn9JgFM5pXeMDEkYmYdfNCo+3FmaATkGacwqAbrEhnpDeShIdccWANI
rZrsIb6XiSI2xrZeFarkA2WlszwMUNA5JXNIOstccaIz3wAofnjRKdYNkC8WiWOH
1jnCjqXxyNValF6ftHgwwzWUoyZwXYUx0ITuvzRSunMHu0iHJB/KNW79miBJYwje
kD89B3dANl8Im0UJuTkG70O+siFW05iOxoeuzfYwOjSQcYEz4KV43bHp9Jm8EuVT
uJ6XkJGcGC4LZoA0H5YMT9KVqTpndP8I9cmBKaYYB/juwX9vF71GUHqFc0GhmHP2
VjE0cPZ8trD4BnRI1GxM4d5UAeZK1u+M1KhinUr5cJQtUr8/pC3rC5kk6wBopQYk
vVYCBxixxkjzizCFrfL0TCn4XNhJ6/UKSXh+VKuMLdqJKA4fQHruhE+a0NWp8Pbs
ZXAW9CRssOXYzpMLSY1PYbo/ZtZ+sWPTyHoJdhfweLnU0na/qZDAE4LEdAp8UF8y
dVqMJYMk/XCC3xX+1lH5zlG+jKGDUDw5wYq0n4ab5uY8v7Lo9o1APovV/fzEhi8p
PJhFOR4/mI3RDwXyf+BaFqtxJt9btELgkWhFHN9tB4DHm9YiGDUvHO8bhVLYxi6N
AgdYMZcd7ZryABhcUC2G7n2kctnHmlbxyOzG174N/tbTwrqy4PgyMyJdYc0cnF46
rIAA42Z80aD/XPs8jWp+6mYEEQrqGHqEO9MOyCB0oQVnPurBNl1ZIy5Y00NE8ut+
gu62W0jAQBWWseEeerpPOF/kOyfmjPz53Uq7J5BXP725WjcZytIIfqcaDiLpPjk5
8NW+fIFSd7aaEw5GucNIkDajwT+/cqxNUEnOeHQVdOePUkcRqVMm9VHM6pAY5dyh
4RKgn9CpPJp+KytAP1Uki2uvJ8uu/JXLu/nw4jHPXMBCZKwF+7XqaMvR5RP44ixF
IXJs1JW0qe9tiVEyd5ckHai7e0pPV+eXPGtD/ATg/YwDDUGr0dFUmA2OdUpAG80v
ZKZdrXwTXQIr/o0NzO3kzpEsBLAo/3ljRImInXw1aQ8EvPRAKjk8aIAtXCG47T1Z
iuqk8eF/0EjYX7Wjx3Ak/NcDkn7priIZ9D3ejkw0cHMqQjZBHArJQhXS3JLBBGoE
b8AUGpTHYoLU/tcZgKNJjtBvgk2QIYFNTXokzSt9iUXP0cqVKGbfEo//g/xFal2q
Q2rdy2VizLkyZEE3yTEif2Bk/O63d0g1sG5z//PPCEkuCE/zm/2jXyniRtl0fO5z
YHDbTA4du9yKrR77xDf28mt/jaVrd7iU75Xbx/8r8MC7bF+C5JAgvoBJ1mBL24Lp
Dad6DJ8pu7Wr12DiFPjhz2OoadD9PSgFAoMkJXvm6DW5yQFqhZEhIRV7xRD+6esJ
i51eFq07d5w2v7G49HRhEAb20etHDORqDJu3Aw32ANr8ohJY5wT5jSA0PiubqGwL
dWcQWeZ6gn4nj2JPEN9F22Ummm51yPUDac+hosbq0pjSfg7r2TIsRgq6ODTTPMeV
QSHTQBI09NtcEFn/560TKcabu2oWnlG7yi5LqGQk9wl9zHAE9bb5lqRMsmEKgrVI
ZIrVLRPkkMvenl+bhYMbOkQ3iiaMIft2N2e7IhgCMCYDYXXMcOcl2/Y/8AK6Q1K0
NmSodfh3nFi4Djf3lXivB2+HfurRSCebCEJ2KDlL0vvsQr6BWKi56J/LF5rOyYHu
+Y8BBSD79mxVoJqmTpwls+y4uFT93CwdpbFmuSGDR6zOesBBA8rLvijyukIEL170
jGz1lLLlyBR3lpnUWXtxs3PhUKzvoKGmiFgfT8jzqHS69Xkds3sMKnMHggGPr2iL
me5gwz2Zsfiw4iAwUApDopqLUN8XKfzCYkJoQ9Fojb5KA2qr//THuJwbej8kUSqi
HodtQRhRxdZS4Sl0VTgsLxbbcY+3YI6r7LQKd2TIkb6vn1rgLPM1tKunx0U1nVHB
8NsApjWQkZ5cR4AqzAuts65dDRGpgL63w6qsGYJ2R5PGzb4uTPy3CivtV9vNBZpS
ImM5RFQF10/mFzdaZc/iCS1P5jYOQpXpZmpB9za4hHjyu5b89D4SKH9QwL68+9r9
l5ye2ww4Wm4JQvj/zlETIKQG9pItzbzydOYibxqnxzQrRsJBBpVd+GIBCBc5sBhx
+alkZB2/3k31wavyLx5vA43mjEjUeDt2w6R1PVziyJwzCXNE2UFSYoOXJ69srtTw
yMM7UbVwDht9FWZ7RIxhDa2ACo4F9Cb2XR71+h2voAski/eENz84z9zCJMno3jGs
Mykegtv7OJjPrnEH/OJk6suT/KwnSFvMaT0ZtqZVIn2QWyB6JPpJykEmPGkU7kGG
CTl7/grevVFvBSVe+WwAveRAHwhwPY4zqnDTfsRN9caATMi1rn421UMYdmmZQCRX
EmD2Bq1J3mun+in0U7HA5IF+8IiMxluPnbpjA0g2NgMG1UPYXddhXsY6eFbMtkF3
Pfo6IGwE9IItxs6EhN2CVjtBI7U94jgh1yBlNT2nWD61QNuVpRl3pZGqFTJV/wRY
Y3IQdwjm+/CFXSkwfeMo7f/zsAEP0Nhvf7QuMo3gFHZeJjYmmO4Q95IbUpSIn4xG
OJLlP73JL8IetUFndRJAJ6KCNuysmJyuauBUja/q5F99Zfv2wwAtF9EcYKIy8TW6
trOlhfE9C6FSCoCoEhjSefXdEvcFieQjN8D4BYc8fvlx2V4PlB9qCRAQvK36ruGf
5184/u1zUf5CDNQAColHR4XbyZfYG/Vz0uN4IWi6ariSebIUGIBl5wgB60DEmYAn
cCRdxp5lfoOK9jwqcNlPaYwOuq1TfPU/ua8/2rTeGcDI9Z6rjSFiSfEf9o4hKgGi
71ic7dl55J/LuXkaYhVBf0rnwCTs+AqiIVQpNby0jccLvNKs+iSDhC8Z1sVsQeZk
Os/dbMBfvAmr/73eVONyx0MA1vaUJCufTXn3u0D1mpGvQF889S2ZcF/+UXEp1ZQ7
2awPve7ICOxu8j4MNKwBIuqvDVWhJZnXCer0xRDkQoh8h8lH6fGyaLFu58GFshPS
pGnLYGudnf2ll7NNA/ByVh2ebrqCwUycJZoYuPcFh1netH8562IAnkPEohuLhIl1
YIWwjnkIZoUMTWybvEL9OJ3o+jjtyEPydR24D+b+11Vqfip+VEAtPnYrIpS2Vuyk
if8nVEHHM+FxrsaG/4KDppTASUedggXcmwNsT5QgoWPeiN+8H+KYdwRp2WBW8IG6
1Dy9YYZ4xfdkK3dqDrzcg01TNHT5Igxpt36NKGBfusgaZByYQq9Befhl4TlT15Qm
Iz787wnqt6ntZwly13wdQeZ55agaZt0a9oSDFIvrX/sSxB4GealttG7N9cbGA0tX
A1Q3vACup5Lr4MdUU9l9wMKTiQDvA33DhP1fiizKu8Ax7dbnzAfamjsHerfPMBtu
v4xw2EKUzHsa/yxR7pcvAmGnb5xdNUZ5q7hCgqBZVkcN8mSF+RFlb+uQ4EIyFkFP
HJZZYlMaB4J9HJSKX05AXs8VzBDjy9kO4fxKb8GKm/X3WX4Nuf6UEBJOzq7l6cWh
LJEnH/gZNEB7xO4x9qWyhfwJwaToAG7sE6RvVMWh6NMZuLkA3qi1XhMKI7e7vf/v
AzMrXIRgnP0TntxR+i7BBLek3z7p7DoBC0iK8SGIv+P7r4wc7i/d6MfR09hSWzDW
KXwWQ7RYgZ4aVWOtT6O2+bm8+8dVKcZfKCrLY+cFXNOmaIst5wnCE493ZvHTYsl6
O3z01nvVoP3mhhtvlE+7ZCDwZ0L/E7VvGXTFQDNDR16HUZyoGoJWvj44iJq/fBBb
D/0dm1dQH8OYUw7UOuiFIQrK4lzDtbp5EmU+Oq9xIiF66JnHjdaxsjIP2EJjVPEt
H2sPyHljWYdzlXhQCCvQmiKJro7ShKaFGjs8+61s9MWFJgG6qTbdezvCOL98FdzE
LyYn2xbkIAKhZYKtqPXE/Za76tocfRewRviT/3LlfyYQQzecmI3feGKs2dxQgt/6
kFBA/XlcFmmM+pyf9elFUtfoTP67/2aX5GqiQtIpy56kJT/PRI61l7jJv1mYE3kb
8pJnl7Fe+8uQZ67y+DPLmNBFxwkT4YS62vnrUD1LGOibli9tl5iLd1mYhf7h884V
WJj+d+scberKR/cz55JR/hzcgZq2AV0eHj8nEsmfkJeQs44ajmbSewY4145BXIkn
/qr85w/JpbaM2VlKQZ3W3MNaUxk9twV08bE3ZrABZ3txJCYVfLWH5xcZb8yvbSV2
j3b6t4sMi3FeeuXQ0iGnZoG5mGH2OKUPJ2diMQImJiytglzWpbZx1wRE+yKY2gBJ
mq06dozfntQYbdYUuZERaww1w/Z6pZsTQb1sA51ySpmyRuOji81GqfPi446X1jXF
UP8i1z3pnN+V+JSVhzabeWcc0s5HdXqXBiNURUcIYmWlSM/1xWxGTOMx3XH6IjLV
6ki2B5/Yj0qjeWiRGCP0Xn+0qvNBm/9vIVCYtI12BNWaNa0rd3vlpck940keCdny
djDmsvC7goFH9CFvfL6l0e6ELicCyS+B4UgWJhVjEjOt0WuGsdfv5LsIEXRHA7lm
i6agT9qK9xkvtSsDFKOVrbWSuyCj0BUYyYSaZK3/ES/mBtsw1S2O34uhvTsTpGIn
eAHCZNUfUhjQRRrltxVEhkoxs/6neB+5MlJ92n3J9Y2YnDPGCAKMLAQua/6goQzP
Wk7ji85NbV3mnCZaGiRO1YavNZ7N6Lu9PXQpuKqUKN0TPh/YbUuoapTFtwUk/NsM
ocyKsC1C3HxxqJawNM9slLmjfRu+pw1H9anH1zW+XmA5U4rL08ucMfboJn+YB0/V
JZOiv5KVr2ogsHS0eHPXSteE65+cHHn8EdGKZI7Wv9IwIazKeJ46N8+OJ8V/dnhf
kNBjpP8PwAbs3wN1NsjyMdk58tqGqMLAQqI64EI8ELsmouXTLDAuvZAbUyGng6Ez
uBSXddvTfmK9qi2/QywvBsr3kl+/aVgZRkZJv0SZ+rY+YLQAJwoimKvLVbqVePoK
UO6419PVcaipFOKZWczzjJecQ65bAkdf40ky2re+XhpgJipIXxO74n9uUbL067ef
xdVerlI7RjSoGi3resJevUEmx3DepeeNgX4LVC6JKs57PESzy/Ys9O4oPwD/5G2Y
x+pJQw/nRTDSy8zHpxMcQsyakoMf9JP7N3R04160vmjDzssh9pMXH0gexmoY9wPx
JNyghT5vP954GbZfpJXJCuUrsA3Nrez23tmfIuU/6j0QF5rPxadARYE9OeMIU9EX
3YgUXdGqC4VxSWMiNCiUO7O60USboSV+8O5HHgDYotG3lfLwYcO8r+hHuCKE7Cg2
G2QcxXXmuR4u1Z0DviaA5Cf37kv5nQx8B5R36Y4MpUFffE/tHfWfa8pWyJNl7FhW
KFKLCO+V8T3pICXwuu03FASw5iiDQy5pQd5CeTRouscodjY4xSlFWhIc60ImoQXv
5OafloyB9TyomLzPh+/i6uW8m2zS5ihc92gOw2cDbPQ3/dYlSsABKDgrvVxBBALh
1nxoTmwHgVPrO7X4WTLu54VPB4Bl6v+u7eGwRYsV95Gp+UaPUnATY10hO1QcZJH1
BjWU34IbVZFZ3F+/e1+Ir296gaF0+6ZFBsWGZDt7/w7L5iPiyN0gihhojxsw/vCa
3mI3JOMXaBF2KIh+UVasjKCC6hX+lSF5nRNf9auVF+DMvXOulizdKAYhO6nYGeAi
e48OoqKvKdrM+P9C2XxvXp1Spr2P21AIreGOYXOGd3GfcUNzioiBVz0xldDdg6U+
K1h4o/FdaH6ngYsuq6YXx/RcR4WaVyLQUf3PjgECC7ooc7bK4xUFQszRNLd38534
aCKqC/hYsjDteZrFLIwkR7LWn9YCFcxq16TxAmAhQnVoiQ1j5hAgg0JjHb1awxc5
Q/K0K9KcRUszaIxrwqekvI01YurAU3N2MUnhnjG6chRSFwQ+N8tujuKu/Ap/prsg
zAgh1GadMLTI1KzQ4QT+ujs+xoAchseGNw4b/2+g7agLyjswFXYSog+4hI1LOIc9
YtY3yqSFTxNCpNAo0CuvqhKipaJc/iM7klmZJG0yQBpu8gKEOw71pGkKQcKM4ckV
Ni4QOj4jf8rEFBBucIhMdvlb5WWJz2h0srdF6s7AKtayAuXEECsgfTHKbmPbJZwo
twpr1noqmUKOABuhNsKBJttdetbJD1kFr0bMBCH2J7qmzjD31zOqrc8dTzN2tXL9
1zHgN0paAVyae7QqnNpD1gkNhBHCbVPaCeQ33t4+BvcNKxqfrmFJRCOKEwaCkLLB
ua0cWBQ6/tM9HCUZr6ZmYaI1fOWbsvA07bOwG28ztIrXHC8n02PHyeDTe9w9ePoN
V83KWc04IYCM3eQCFB0ps67xpPa4U9pIYYDvEPVX+TJjl7ebAMfkMO9gl5wVk6pc
HaqXHanr+y3HATiKTg8sIUbqPFDcJ6mCS7adpG19gux0PvqYNtUxnC0U9qQno9Tp
T6FPfD9S374wfX2OYnuzGvTVvGe825SxARy67lO3io+StOWaok1OJOdVtjCytsfn
pQafrDDK6eWpaohpVMH1R3aGskuxhQ5cKG9MEIJ1js/KqMsgjYIssqp8b3fGY2UK
LFQHtETdiwTfz94JN1TyvgGofsT0E8FrgEsaSLf8bpg4iWj2Mgg6ZG42dCY1eSW5
HblrV5oC6MaVChVR3wFK9hilvVO4OxlfBysoBqFi2iZ7xQF4GSokSWR/zCOVLrk2
aq8QQyGEcpGxaRYbz6HVDw/fP6yGL47Vy9m7B7UDLF23zUoLvtr4uJX05d13A9g4
w0L4Dmc/+pSIS7t9oFlyMsNoVGTOHz8ZZH3fdGccFIKeEhQi1oEnXCNiIZAhzdd1
1CPIgfMks+LcLgJCFoiVrdX45AWqNQfUHbIwq1y41KejvuA3L0ZMnTeAhgjiG7co
iA4YrqGQGk90IvnMErgfH7j9YlinJWdPlABp313myY4s9wT4NTS5MNkltJk2p1eC
hgx/fINq/sVpymn2OSUQGYP3IFu5DGTKI9W9yfLWZ7of8yP/tItotwP8C1zI+diF
/Xk0XjD4JttP5c5mCfhZ1a7PKVqL0xebhzO5JYIFAlSaBkXluGpZGmcZG4C2VfCw
LsiuppXO4zZ/bX5v05Wq07YSuoudDKLQj3WcVkEeXKP82q4EoOS+s3BtnLFWqXrO
IG8IboOxr3PGWSp8cUKk7YFeQZUsiX4XakrnqH3weM3Jg2ZEueF4i4Or2RpQqcIw
dmy67dEoEtOjHSkuluVnFMbmCYz1DZG8c6vTAv2k5CVAdu8zZ0VzI0tJj09R9XH5
L/EckuuKUoVB+b/akW6nGpGlQR2vuhHroG+fbyGeUh9Nw1XR6ul309IuPngFMQuP
bMdtZLsW7ReBX56UNQ2Ew6qzdTull1dK/+OShPHUQFvOZmmPYL9PjGhMq084bgCE
9lIQROBFRLdmmcftEar3KsnX3SZZG93pR4ufYH6oZfuQGIxQkSJHSHFMHc2jgWru
EzAbCG0OuVoYZw36kbSe61VZKvVpZovZm4fZ9583lCEs8BroSEo9XeIOG3ZbbONE
NCHGuJxPfhMYREgR20wk0QAhq2KiqSx2AatNufmfOBXiTrQ2E0lCj9cldzZg7Ivk
FSP67fWtvUeqVOUsGr/XP0C4snKDrGkiatiClexEA6URUuleh+tH8aDgz8bqH4Er
pBI3ImhMnti3WUPKHBlUxoBkVtmpFbbvBULczkyhAlAVTSKQlGwhjpFsyr10mPrv
CNHuyes15A2Jk1RVjmImHUm8fJXFZLkyFQ63Ic7sNlgI1lDeYXnKzroSlD8IYkPx
vkUL/NXpzbAFMbXgeRicktVnbEcInbFVGBw5qEgoQuCKxUXi2cXfBXsUYHqys6dR
yBW5seoinxrocQZClvlABTe76+emGDRJ33k1ttRoDxAw+nZgDNBjrtXBDDyi8njA
JPBAJ5lww8UJhH1MBbbfWNBvC1IXeCRKntbLbnwrOXzxytavwCgDafWYACot54d9
65ehDcPo96SkibM9D3qxjU3V2G7hn8TW2QmelPk5NkB2qyqdu0vwZvnXAIgZlgCE
QL/K6/9ErgVepgWPGhnEhn5jCT+zgW8ZPbXsaIswdI7zZ27RZda0V9BrFKBxAVzJ
Tn0Ua2u2ZDp6U+sA40L9qQpjt6lRVGKDZDAR9smHIHbi4XptjQ9LGz6aCGDO1098
QSvtSmooDWJn0bq+hIMNoIeWl0hGKhn0gx0OIdQpzxXIhrH5v4XG2R3zn5mfYyPZ
zZ1v6ilBKXjLNOMPlxMb7c1xPf2GYVlbXM/cJGqPVMC77wWG2Z9niqtTzY3JB9vV
30RSIKKjsLvUahaNun3e7dLT4/1Pe0VNyQKzoaFBtiGztZbR4B04r94zxyIGKkeK
QR5WhSceq9p/igPoZ5oXY/c0WdRQO5///ktxOJoH3d3kR+yPGV2nqR+x/5B6f9d8
ZqMRx+VIW+JShL/kzEiQEcMi4lC6VzFAvf/V2RPQfZ/lQdqrPplMykIKs9XAWNWA
Q58UwSZ59Mz2nG9HwCbEH9682pc04Ln0EfdqVgLgmtI1YtceIDiyFeDr/vH3h37M
89H7EFmJwemUtAQxXJxoXsTgfiFKyb7xz1opNLkuWJTB5oJJTwOVY1whZ+d1JnFV
rKox3dSDn9PSFWRL05MNAla+TLnDtwzcTHExoG38/E/mO/rWoNj7jnaryF34vBmw
F8GzMSzUglmYyCXgwJzKt7IsYlUrZNAGJP0SB43HdfccNdK22Q2oilhvnFwQSVwt
BxPNuFETrxhGcKiNRlNNvUyRcoE+aXp+Wluf4meS92zbVv/m9+LnXheOIV4tWafr
jQrpTjTi5ss368AyXgM4+b2M5tQAdXcLQHkCMQazI/+Voml8R68KZOYNh55msHFq
0FwKvDv20g+ocXGCIP1OhTm2ykk6Q+2HBh0EuDyS5Ft9Nn9KychCzmxQ+ygV0fcP
G0zB4DaFsWOu5mheM1uwNAhKwMvEcVcK04NW0YzBFGEfpUq3Sac/aQuh1MCLfeX9
YewM1MCTIIkHwkqq19Cm59KMVdLdFD3J5tWY6TAL2zekkvy2tF6AzZ9tCW4Es8d4
7ydSa3sOlW7JoVhE+anZT5TlNx/RlqATTlcg0G40A5IMstTCrsoVnxiA0O0ss3aN
BWZTiCOqzCtx5yV30wWNCTdMdhzFB4xDEvyT/DzShxlnllhA5peIHBTBkmkfyTTo
0MlFRgAv0fjtWxNS1o1ApXsvlWwi0nBiba8SGJf0E27xY5GNA8zx4FwmJPlLq3Sh
E4G6GjTxI/ULjPUZrSlSQYQmqxESbbr9euf/l5rSqC80ypd3HFlxuqdns9GXTsR3
2tcEIVpgYbGIQz/M1K6Pl/X7rhZuFhWqFV3wsv7zyFCDx22/pu17j9YIqUO9Wz7I
MmSOrNOE0j4L76PTnuri3O0loD0AvR4P/RfpKgevmJVRLu1z2FECUT3ZOtdG5lOk
JamApyugi3EYW3xYSWpO447ObeelAwe72UitKtc7flfmu9NSnnLq1sMVggrjvVUQ
wYapFflNW+weZkfX+wAVxuuCBf5kII/i8CouEe0NdkoVnzHDH5QK8MPqR9z19o5S
UMbAdt0dh5OxMpbixJWbUeuRj+t2lhEpHluJzDAi5ZIqJ9RShUkY5R4iwxcV1QeR
J8G/1XJpIcrebr896MgLzFGsRKjANdS03ZyfNpFr3RoFCcjrD+57kwsZozr97ffF
16SYLmtfXHSTkekdOmcHNMFZEX8w9K3nr+il4EDZq+c5EmVMw7wqMcs3dEacNe3o
1CR6l1ZphYHd5m2fY6fF1AR52ZlJeqHELt2h0gaXqfFDfcducuXPTjXCC9H2Cuky
j8mBsLekYCEspqfqPsFfYwrzruK9keRBAdFMPMRP8jAcNg2xyOzAuu0EHdMGbnCC
0HkKblTyIDUXwgy9xNQlhr14PSS0o0GblS2QzvW8e85eDwCH/bXSGnJUkk0pRGwr
jrRpSTxGYvMGGLZw9JAX6HaUbAJw/E1dZoXvJ3Cr4ClKpd6WoT7ZoeWX9X8uaM6h
5HAOsBRKpHcpM75jwhIpSQXqoqyleNVZZ3z42P+NVl6uYIzAwVnMMKtEI+oVduG0
vabj3yza5CqtwsVVMSJCX/cNQC1leeW5QpkYUmOwMF76FEQFCU4kvwQtjNiWLLQO
Vcc6XDKspRFI65g/p+Jm2zlVgmTB3qaQldvO5FjvDLGoL4KBP+vydT3F4laYE0OQ
QK1guaVYLvi8acB/74VhjYQEPDSK6vdY5fcmYGC9LLMsIWE/2T6NHUMRR9BEX2mm
wvOJwtZx4xbZN60hAwZXIJPSuR1cCTtcwjF9EDfOLnFyt36VT6Yuz2gnJuRJX3dQ
IEKWUyPRWyX8fgHfOwA269HY7KTnVhWmxQSnBu0rayCYi40eUR4bgC0shOccr2C4
N5cX2N88VrVbPmtnjA6Lx5na2zqM2Ax+OxCbz668o5AU7FdscV3OcG3j8KKBiLy+
/G8NQr58It79MTmeRmtkcOCf6DXtoaTsFxw1XGkw9i1tOLNGTXSPeNgwzic4thvQ
daU+ZGH0WLlB7CRZJf4mGcatkmsQvPgFre6GGLc7DCQWnx+wJQLtJbUQjWMCoVBq
ZGDdhNLHPdmETecLbWuM6JSnO1oaZ2q9NcrOsZZSU0vBjBjuoQsl4pCuHb3qq26S
pPfQnafqsAAaR0nSHyY9y6iYWEGLdIL0G4fUPikTURR6P4Jp6Q+P+j+TfzAhy4eR
xJ0LN261Kxif5hT8p/NsJTk5kkuvDAe+b7ElbglRnIaf0LEdVTOELJBgW69FpFTl
iiIA7M51pxCYVPVxEaRCcTnOKs8r2WnQ2RCgq+NbvDoWZe4x4TBHQtqWdcWX6JfB
O4ZJgSTSgfXiIEDCqk7YVimGXgGpQ1mOjPa7wLRd00GRAmFF2Tq5nj9TQQInslnx
RJ1FhZ2TOphcAwh2nKK6zvfOnVRWpjLC12ST6EK3otK03XBhdqTDiO8LLT3w25zn
SoPLFfVMQeHhz2mWFzScIo5AbNFi7Bym5nNHpUOtIs6jVMIERyX4+G2RUvx2BM3X
oWqLEg+NMjgJvx37aNdEzmiSUCzD0VaU4vTDXaoEO53J3iwtrtRq2lIGBgoBEjw0
XhQAshJGQ1EpYBaXi6Y4cFdG386vHObns3M5GgAPqa9Wm9VfRLXNn3M5+89PvQh3
iehCPbc+UxTny8DqnOwOGdWDugj286j/Xo5ISnEhR+uT4ex1HxF9EqLqvjhlQoSi
vhcr0qVdWF7fYL+ZT4nzgeOd63SFrXDFTFTzhAAQ9TgI+c+2V/LErOWhVPpOAeZc
TeBTdzWCYxUl/Y3ScU2jDpeRGHgLAqBpsDjtgCSlxNQ9C1KoMNBhl46EqpgEAwGT
27tWEaLTAgDXbB04H7F4ZBf+E/xxzeRx26QlO2N5O0w58X7z0SbGA1NLlMzmxs/x
sG9RGqWDHqQqO2CAJ9tG/cbBqyxdApAK2boJCcExTCS63qECzhjR9JdfLhO8NHec
exfgxEVMlFu8zdQpV03WoOQxUxuObOiApW1QFTvJ23f66+MiZSaK/brAW0LRUrlj
2z3CrasNoqq/OTdAp6YxzSiI5Xb8xaDTe3fMhIFhqc1ITgC0EmaIJKwmvxV0sgST
KjHpx/AIm/lY44dR7gA7irrMSjz0sp4IVhWbM6zHdE85sC96rXpEaAbOdipAfO9D
RVFuMUtjpDq7ABJkV/SUrLAazddkKqUY1q5n9ZC4semljeNNvA5TexOXxGxMusDM
VeCTD3ma9czglZJfE6wbymW83erjnwfK+GIaktQ5EAjUovf6FbYaZ3234+afE4em
6v5K+48LTDbrBxQQ+7G82N5+AJY7gL9rHIi/uedPciG7NOL3uuM3oBVhdSMaveiK
gHn3CrXmzCGUdDGrY5KG3yBQNcpfycp8dr6r8Vday9Cq1HI6whCfWQVmaLemGTzn
Ezmr+tSzzplNyNs25EOWguV3OrCGjInb0pkj1YbnI9w+RZEn9Y2mKgFGuXnEP1Jw
WsbQ1Y/obKydxGYR1NA9O+Wi+hCRFZig2vLk8aiKokAapzSLpPE/MtAgjrwd/DXB
meStNUO97ksNkHM4YJ7d1OIU/Qm+oTqvY2hBBcWLVFoSqdggF17McsqkANR1EEJO
F6r4BG5Lwh7J3D+LIXtzBTFWluExsMoxl5aiCAQzaHNQMBeZUUzDisGBfZpEfyaq
E/Q98PSVrGd1jKZODk/iyZ8aUEFq8eVT1uxP6s9ZAwuHkbMq8KJzfuNfS30jD0e4
aQYUuI8e8wBkYCLyUTbwEMyCcrE6r4nNCiOb1nWcpcSl8xb4egxBPUjFBusgeeLt
RtGKb0nE9i0a5j3UgdTahMpf/U2f5ki8aOYkJ34GdkzQnHFn/jZp8rkhuFNiyOer
70cHKmur31ExzLLZmQvKCpOeUvYJM4wa9SM9fNqQgbogdRcuFX9hKZPjYuXiO0NB
SKtrcf9cNotMOiToNktXfDqhPa1VzARBtbdAD7NIX/nP1GFpPFReN7iOgnd4Hjwr
zhkDGRGIPX7/WaGD7LL36y1YytUhzyr4AaBk1kUGXOHEEiv4W6+72QOEupZy6MOB
ghsFocoV8bK0Zd5gk+pRYI38BZcMhSNa4YN2C4khQCwrjTTqOjBjyYOfkfcjWt5A
kS25yoVxzwDV63hXaI7Gnv+udlJP919lSSD8UTZSfU+KDNdezkbvXYxdtnCBgnfj
h5cvQJJcFiusinTiEpf06PVT+IWh/k6pHf3hpgkvWIt6+hxaO47Xj91WQQSlNymh
F4VPUB+a4SJ8CXMf+VYCvW7Bs48IdXTiq4rWXnSIulkFnuMEphCG/Cfw8ckB681k
TCybei7lQ8L/N6j5jSA+E6TkYPUupIucVGdtqPvsPxglzHTqXDPCKB/hbjC0sQZo
W8WiFI2UXTOCKlY/KQy0j2z258hMCTd82hTXh2d3dIVhrrXBWmFO/PuCx9cgmH8o
Zaevaldpvxm0kZhdhSyRS+/s/SpGpEC0/AJ9bzCN2JCxRo6civs4nEQ5a0SwmuRj
pvbDsxZMLHzp5CG7AAiGGbHOrHFHQwf8vyK/3Mo7UCogJ4eklmIhdzN0Vq4bvD4i
0HGktK1XT15f0PNJb9VYZefI0xYMHRhdqUip1Vd5fGzm6BuKdPCTppj3ImIz8xE9
xlVOVM4cQ4B7hreq5rBmLd570x05AcNP1AAfJ9bd7K03RVbvknw5ous1STgNmvDT
o1CdjxYBehacEn4kaIAT7sNfGP+Qqklf6v1CfMJFXxN90ezL9/vnO/QpK7tSdr3E
8bZpAx1Axyt2RzcRBTF0RUGLJvv1LIryu70YtOQ6aUMMCqNUo+SKPl8U7ShvNnF1
RPFfU416vHw5lytomonF/ICfrGOBesBuyeJ1l54lnkBvvX8oCauiCzRruxG9VLod
mtECXSm6TJM7IiRA6JfT8sPB2W0CvGoiVDWUJJkb6j+Z8ck3CDFWEfNls7dxyTs4
7l78ITiNiYa+QHo7KRddKHKa1qClIjbg+9WBTPrf/1a2EdELoOPyTN2t01PCpZzp
oD9wo8Ya85ks7pK45AQbxLKmjtE0tdNqEF86Bh7ot0g2HBnRN0yNuOMXUwLgolSG
lKAIB3T7Ba2OXM8jaUEOMa6D5Qe8lMwIlev7sbFtSvnHnx3qCzqdf5LgilLoiW77
0xaqCWT3Evz6aAn9Cn7MvRscsazJ2eXQ0eU4MFl+3jURIzLNRRB9hAKIQEvpmK80
DNn/ELGwPTPZkRv9kixg6vuwjk8El4JmcNbw7IXrZE0Ht6PyhnB/vdbhBuAJI7Fu
zMHlvKuV2oxZyrEZOUqA+3BxpE2SFhtJ6Ewudgg93U+T0WFB4D6vsFGT9Lo/Iuqe
fj0LjSQp1xLfMeh/y0Mbz89pDqnFqmlkHl3eAH0nUFAvY+cFosew0Zyke7P08jiV
GYQ6FJZYDrJwSMvmhg4V75txGEIfysYiT3UeVUy0ISmNSfP0fPHfF08YwLqzve9r
2jGdy90xom+w6ZVgpMXTrLSE2fPjL2NYCbIJNlhRUOc82gweIjfAHL0wEouQaSjH
cuL7hp/tk4fjqMvE30FdbwtOaS0W1/1EVBww59F9WSAl+JjO22+FskocvrnJpQxB
hII21PZb3ycTUth7tfg77wg3xeF79KA14feLZOmojw7aSMur2tY1dQZqC6PLlFnr
SAVHln3ZL8cfsc79Dxh1Pqfw9vIl9qCoh9tPs6cY5vsq7rkuzkBpTx35ZH3sRetf
2F4KBXblE0y0/Z+p+uNd1PNIPX0DvFNeJ4DvyLSlmiS4IRSwlRZf/1+r30VSO4BI
Yviu35xFbN7sfoLim2T/72cRN9F3d8UOoXFwOqJxapHHtTAHAwBoco+ougYrpzVF
vEhkRcuBHFAUBUANYJccgIbRKx0+gwQwhVjNRxqXggWUh5OqreYlTGVbpXruKBzA
OUGyWA1jgM6pJDsCxtnNtzAJnPEQrbAP31ca1c5YrMAXqrRsKkxgnkNStIQHnjHU
l+MD5tF34RH6nHYMNXUDRitie2NNNU8YXfDlL4mJls7TDFDzEz4guw1Lo/RnM28c
qpf81I2fXJCmHgp53/x267ZKI654OJIMlzrb0YqFnjmBDDyPr22Q3ERSqEqTFYFI
ushHmWB8ndd7lCdkeP5ilDmY+X8Ze8oD01KqW0kG80odnH7RcOq/SUd4qj8WXRRX
G6aMqHb2loaLuXEC1hOuN1/xi/QdbpVzuO2j6CO7P3fl6WTqezyZAM761n0f13/8
kc4Bhg3j4zgCUPU+OGk7eU71VN8LNFBJyHeU1L6HWhKEePjDXirM1UC7MHxF0E6K
o1F8YX2ERcwyQBWhzliiTG3/7kKQeVabtZrIniag74WfnIOb5pIgo573cpG0WqCf
C3+K2XizK4GDnRoFsazblmYZvMrwSmVGS4IDbPYMeTDnVwGHhGjcj5SIa3HOsO0h
BvIu3VyCsyf9aqn2oS9Gw4dhAVELdaDif3uqak1IH1sUUWK3K3jQgYRfAoe0Cwv3
QVYy31BqW0DoCjh6xgyT07kgC6lee77F9CaC3csXohKnM3Ts4OiVRgTygNgdqQCs
HQOCC240jvWLEDE8lmqoBY1uUjRvgMDUK1YtvuWarLSPL5h9wUa8ZRSDEXorfhOV
Qr4ZcfgzzCWpKOempolBtgzcy64Vt1p7Jbhz83NeNuLpcuJRKMzgZ8d5xX56Em7E
BGBdg86IVdhJ1k3Eu8TXqkQeeZHt2jp/ysM76DZIcSSadNYjPbwfEfVqrAacOxbb
TcS79rawiyRtEU1WtyD3wm5BdrvqLhGhnlmXV9CAr6bPaQE6OiMbw15RpLHGhB15
jSkpy6bEzI8kTD0SJwH3kCvBu9hQHTT0aOtuUuGHZu/96o/lZCR1Xln/3GHQkEVo
Rf+/U8fsmc2M38ZD7FljtFAw+LmlGphn2KaSDUkMYmBiL9W9nILFjN9D8vitgCoF
Wvn/yE6mJo3b9uJOfE1odC8eV9VWuut1/BSgzhZCLC7YEPRxsQCDp1loeFbggN1U
uMDQoV+yhzNvpSSRSnc7wQHKepKnLp4hYkLKm0ln97mCHBOxHcMrBQIbevGqtaa1
qHgl+7qftrSZR0A7Ee+GuAPe7Xh7bOHzSo6YSj2Zy7bq6t6f93x5CqVT1q3YnnUH
XDQTunH8q9AiVaY+xRusQOk4GG2THfvD6DcQ+lojTQmcipCW0G5HcJvZGe4zx9be
NANZhrAkD7/i6MqugX7Wb/2qkN+v7JZ38jrjMUVmSBWLgXxcEsmJLO9HT7k6ZiOR
7n9IaWP51+Ro2Wyuw8ZvMC43BP9XNUX37jbYqHcO6jKKuVfrQnsz8rFMELWYKgjR
+qlI/rYrWIBTwvDAcYVK7EHyf7FNLmFvEJ0tqqBqtajlqUg8KFNG+RxWrZTh9oiV
KNpx1atVvbFZgfA2heC2sYMt1AXxjLWilJF9ho4F5kIo5Ac1metXeocWjGRCakOb
ot/7M/i0eeFbESRkS+aoWKyrSKw4J06H+TPTjcxEgJaLQMHo2A19XifOa3ftit+V
gIbI80XXFaPaZpqyW+dSKE8ZAfMCGGPXxfW+BuFrHrv0sYd61kDNAIDxAa367ls+
Ur68hUj3PuyR34pNUko7cFvhxI/vM1ilLbCAaalM+3r1v4hjWLVBvWLSbfRyiV4o
mAvRjqqwqpSJOYYfsSRhkFWrElFmm3+cfsm4wHhYPjeKMuiQkiqwv1rs74AZTdsV
20ru9opyDaHsTUvHtia78tELOtHtV4UHXGrd1xSxnXNL+HqG/G5dUyRe4d3e45TF
qgiRyuAF6wIHx63FcNfg3NUDtZHR/gsPqZUw3SsYEQloJrAUPAa8gjgd8ynYqYYp
QH7RS+pSi/aWDiriBFsovTbTnrgKGxRcOTNUounOOl9v7QBDYlVPa7dsgkjq9Z1t
4B1CzKNxns1vYgBc7hTwBZ2ohq6ZtB8w0jr9csatt4pw9z0ix0bflzWPW9LKueQw
xYxP4nAUdGnCXP8ojRyS9vLa86H3moHkPU8cBoYqRMb03OL1DEhK4OqDUMsW/llZ
sbLm4JZ6WNLLqtS2WfZO3TwSLtItar+pSYOyTiBlHe2SV9HmmX4zX7V/TGr0Jp2/
1vWc1rjuijcbtpZYop4u59A6BMoCX50ON3wHcXHpqBts5Hb7D6AMNTu5k7kQQVXM
KsXwxyJyn7Db6/2sTaYPn2JXF3jxWkB2kzJJ3muUMelOqxgJoCl8sw+Ld5VeXJGx
nqRA2bR3YcT7yhLEhD5u+n/CHAHwTHNxVW52UTQPLA0fWn7ZtjPF+baty7cJQnDf
bpiLqjKXrBiSeukxlQuIcIY5CJAE1fNCJtxM+Eox7c1UjOrWaadCWtYmA/knkbxC
dhCHbY9b4rGUaH/icnA9SGBfBTjggtbQRyV62AK56XrQ7fUG2QepCEKUre7IFFhA
LRL8RzcNREAGmFv31KUt6Uf3Mj2GHvdeshW0nFxEjrX/6aJbPFanrGYYQjWIyM6H
T2NLeUxs8Qlr2VxIsfx6yImIkev+7Gn647IvhaFJQMfZIvl/n+3a2Ug3fCD6SZgD
wbcmcuHGNvmUXkVkiAS1UKSx2XgWz4LNLBPNnvr6z7vI0MrF6WEtgUqBu/THpVEd
218hcxxVGMTr9FPyJJd3aEHA1N/GlENtcxLGz4ESaxxjQekiaU+Cgytd1wJ44ccx
9vNnDaDe6igzVt/Ox37zUUnVIN8fneMr8GWQ74Sg4+mCvpOTyko2wFrFH9MMUWFI
N0LwwhgzCg3koJeH4SRPGxPgq+Ya/PYt/UWV+L0AQd9Pi+zsRJYDRTBZajDI0o3i
qNFO08P1HJKiCvaSESAz6fxSliz/7IJ2EmSEq3Nxmv6YVE2dw3L1jPERfQRF7sw0
ZmW/3gahMWZe+yz/EtTLi3KGiKgwDqih9dJv+F6oIttSXNqIwTOZM3M3HSO028hJ
OYSIdMZfdsFB85oW504ip4GnYn6KxRHkI/0+3H3NRxIPLNnh9GY5vsr+JUf+P2ok
7UNjJAFmpi2bpveJPumVQ31GoCYHwiorV/Ke+X12vEOWfjjsLNOpka6EKgSZReTZ
pAwjK5bAailJRTd21uiRhGA2bR6CWqODl+PrkFBpxGQLmpuUUrFqQMwTwV4Qlvrr
M6Rsw6wZ1zmvps/8QPS/A/EDuEQBLj8Y6z9H01H+ASS45uQFsvUKwzcP+N1TMtHw
nw/iffAw9nz65Ghy7J5zyQlyluIXUsxYvTL87yVM6aLd9uQftUv02hYddH+r4P6n
b/wr5C1VhaQqayDUfXrGEyDazSh7ZIYYCDJC1MAALXsOGLl2bENeXvuNpK6WUlF1
CJVU94Da0dwDkckz+9GS79oQ0i+MBA+Qy2qWUiYMEFtUtq+AuQofAG3N39owpqqt
wrPfZNDT9y9iA3OUrQ/BcNnpxXDgnMoJ/y+XkoX+bt2uhO9uQh8Jky7UfTAylv0+
DcJk2sCIxyeM/kPP1qMJ4/D7E4uN/TvH1f9nvXTYielDm3fJ0mzA1/GPDwbgk488
7GptyQcjFbH3BaQfTlDjLCRD6Qyc5JSG9+1BvmmW6p2ezSEtewF6BQRDa4RFc+NW
sQo3KqSf9JjwauaGYB2kgMgfsORvwVEgoPPCgSo/iKZjpZaXlPb8aCFu8TAoHWeI
zwsTFcLTc1Dv6s8i87bXeI9fcqZPjiOl2Dami8w1YJ1CClZTLQRepAQNncu+gD+Q
HoCVRHyAy+UMqGFpXYUq57XH70EtnYfAAdGKq+HsxiQouhwuckMa87EAP1+JFQvd
ZD/sx7D7cFNm8bfLvcixW+wKxaX/Hu5drYStHbyyuTqjv+a5H3k3ZDFCvNyRMLWm
WLPJiaApBiWrfMjxOQsrAKddr7XbOg0VYU0sdXpOf2o9cngxjmpSrOv/B6uI+Yd3
dU/NukD8iD3PCLiQZsTSTYiB2Tq1dUxcUWc9BPwZkSS0zO1PdR+lPSt54Sdw1A/U
zDXQr4CXmciInFK9miH6uUfqqlkdCYeP71b4oo6oXxwiEmv1fF1UeT+i2A+7gLcr
q+dQ+u8ejGSezXBIghxF5uAiz4gE49P070YDFid+g72cNy+WmOrNdg8tNPk0gOP+
MSnjlzW1sCl2DWhOX/An0afeo621pcyVmJ3nR22nLX7Lzsxbc1HtvO9FFZcLAszu
ITqpbFGep9q8HyLeoS2oXYmQpGD6RrHA5ENwL/330PB8xmis3aGUEy3+hkMMuYcv
q/75osWnV9HNrJTGk7nu4oX9hqgJa7fkuHmHXsBkwA0EQ5HPSD5Hb3n9m70K1LmN
4XLCVvyejEm3I52tGTQE2r7us2xmXIaxrNFIHO8iKaBqN/nqQh8op68EXvl3kBFI
71cfIAa1iN4mv84DGqWoKzay6nyy5KX3iUtle5KUYrwk2hVtt9fVX3kkaW1hBo4S
gP+NuHXaP8gJI/0FRymqB0IemQSCPk3l02CLtP3VtHrQCFkhO69Cal9PycrehnD3
OtQLXy/zZtqwxcNntKAV2DM1d1KYuo8+BmVgWpWI8ERvv/Nngg8c/MI8yjFhu44N
SsLkIEhXWDwJ+71CCq2Ly03in0lWTIFQ84S/iiPapmAWOewUOMNHdjPLJ4SosgQg
bZ4Qjqn5ASeqZ3Nuuubt88hlmntGLLsxCpbap6N4Bu4BRMomqvsC2Tz7cDwdfdZj
9tTI6MkptecIMGc+6vEwunttZfmwwiGuMkomtLD0tnFqj8Y2TMFDZL0Z+v7r6YV3
lIfj7MQlLj7iKhlZ+DLDNTuOnbpeof40X9JFItnKZYB0l/H0efJuPGXx6hW2Eocu
hPx0r5VH+VTydUu2gjeVYM59YLbDWVXEkvIP63jY7wTH/t73qp5j9Z8Rf9O/TXA7
at5Xod84F5xFe/bPJdF8y6AHo+W9bZSY77t34WT/U1X92dRBh3nWTtHs0CRVhegi
qEMzUTN8SbUbsK89HKip69fmFlEsx6y8J7ZfP8jddmJs0FGROzK2mmaXFQqjgGZo
yaE9PzPntB0y8ULSXElnE8RydAhJj1X0j/SLrSgWHwoaALQg7knPk/c+RGr+m1YC
s3/pGE7T99uw2UZ8u3m69tjrGDw9A1DUDtzJJRu2chFzJ9BfXSXUcL1RLLrdIsiZ
RxXnb+ARlt3zr2UWjZiJlvgX54efBemfjQ+bgmSHuobJhzN14LpJOJJPE5kYbJmk
A6gaW/KZzPXjBm42kN1h8LT3Ink0M8YmI++2nQYVdVs9RjteJ/14mYBZxf+ehTwi
Lsc+W06xQeLmIUGovBDrD3d8ck2Sde0lRT9AiEjYGibiRfWO6q2Ce6U3NPnx75BS
75bGI1bnxLUBZ5qkS9lG8dlU0M5P63wf1C8FNqd/FbyyVHd3xSlficqJFHjMBs44
2Hlfc+bnfxlS4Et5W67x5hDjNfpvrOLoKp1/tu1M0KDXBCzII3h1kXwTQMp1Dm5J
EvQFnCGAbbWYYk8CibbEoCruv2ggIpYHC0HOpFZR8jYV8aJ/Xl18rxhwUd2okCxS
jMOeiwvUqQY5O0x7/YjHinrvm/giROYd7Z95uSNv2Dpc9bBT9B9jnx4rbqghT9O6
caR6ja8wKqoscnQX2FUIfD+dk17xKKg4YMhPAEe1JkDMkKpA5IAnLlrbhuz30Os5
5GnPLltk7Z8MTCynDd75uVvlk3slNwgV48IS6a3V3UPPePzYVzzI+yfhH/6QIW3p
FbksCXnQ7Be0717/x2n7zLXPxjP/sYJpmbYu52SkC01Uj3ZqLKN/DmXWAmcQZ2VX
Ho2vcGOb9giYWPlC5+m33vVECaixXBdbDLJm0q4N5DLR1D6gnfmb3vFM5NESwCJ/
297xbTiC+rgCw5IksPAZ3qY7QOd20LbiPQTe14JFolZkKGk4boqIbnpp1eukcBq6
++gm7mrI4uKZAdM6ZV7beY9twBx2YRBZ3spPwwek5TzP4B0RHEaYxsNC9S1x05Cb
75aVdnLH7uf/OVEhjSUS9eWd/YjrMQbSVxyq/CkoPHA/NY2KE3W8ebXLhEFYlZSa
wnejIekiwKjee60cbtxEpH0O2IYPZ7/hMLqXlQPLm3KghjlHMnRUvCjW98LNi9as
VPmCEBvSKeNLOySxrxu2AZ4opDa3N8XXBammGzuOrJ5mETNiFCYgi7ti+SkMPOI9
QNbPF1oTCVOvqK3PkGfUHWi9Sec60HRDgk6La2Tw8Y48pUsyAn6vyKyMG+6FSKo3
xIWIYrkIN2GJDhZIxf2a+K15EVR8ZdxHb4UEMd+mdcb9oiGaAOwDib7lgaV+aEdT
hwXajXJY+yWM4mlzuq/u9a9x4evGdjlUzOYm43/8aiccwx2MFHDyWb8qRUg4ff7v
MnC9FBehQOpKoNrcDx1lNBa8L/wNm+hX4ixYnofLX26MYCneJTyAWgNcsljecd/H
CizyR3fAFu4sUEP/PfbEGPMPxVTnIpsP47ylhTMTEsiEhyyAP1tn3svVw/hbuLnb
loD/SYUAvXZt1Q4xWnajA3HVyptURmqhfctlzLTJ2OfNMY4iCycCAhMjXwPJwrgr
cn9pnoX1XHX1rRXhWzwrONuWSUyCsplM+JoJHIijfu30jSfJ0YMK2h+BF6rBb+gU
c+RiTCZI2mEwexytNaYuqzmEKbXEXLNQZRhQZHrxRNiY3Ga4CrTCfpd2bl3rRXaQ
qbIRPeekot8ZYkLflO7vCdYyDJBIYGxtUUojfVSAmRcnFlxz/11uYq86w5qtCyL7
sJL6oIS38yInLlu7g1tRZjTFb400Akc/i55PYrfaN7YvaB9zKPudUi1sQ8nPLORB
jedNFMgPme+3qrgcytEnFWRGrY96Sa2jo22v2izjmmAAWQLZ2JhQ7YUxR7Yw3/o1
mkoBY67pW10ZV47Ur3oOmUcfchXbMmLJzh3n2X439rOYYRhmwFCrUSuU3VFVw3zR
/S3YT2immiwUxLwTnKEwv8yeoTRNdhWTFfNnlBj6XYYSFOO42bk6zOBTv3s5zaUV
4u2NNbMchtUvWOyYYgYM5Gm+QX7oN7BbtoBmxPZ8ilxeCXxAcdSUVJglHq+VFGz4
p6go8XMLPKrQK2/WYCGZwI6ii63B2Mdkqm79gBQZSiwjmu5IE8NGB2PdIAXVxnjR
8XrqkuyPRpGCSTmTS6dbxg+iWsGwZQ0/gS6AektMP0l92x6VsXNaoFPwNLoVSFAV
CHKEjoUey7PiWuEiGFFNDF43LsI222MTkDML73Za/urIFoHxIkz7Pai5KO0DoDHg
Fde9Vak3XC0GTVEqB5Dlh4e2xBDspsBAVSOcHrsOLv2uazCcxA3sgMZrxxSrc16i
cPrsYCUCUAY8Zg/Cd66v1tEPqEOlPG66TcRegiQ9QnalDwZgf4IgIZ1PzMRT75uX
KMvqeZM4+KKwWiZ2bzvdZ1Pwd1rrvU15oknFWFXOAaORTKOWl2Twq+/14wJU6SCC
okKBbvmsmZqyyal6xvoR1IYiKfVblFN6l+SKVCtO0tV0GZZbINlz/zvnVfsLB8dx
rLFF8CtvNhZmNc41tXZI0BDBlYSRStG4cFX9F9aQV5TOkI6AaRbDkW+5UWJJIpgn
lv910DQAPZwu3xlqr48JYudHRW2g84gDgjDfS5fPmx8OQ0U8eoFdg28Vkjse0gGJ
1B0L64pX45RSv0CaSW7dK+LOSPxK+o6FQeSwzEkyd4/gVlVXYM8q923vBV1PYphS
OtATDRUYqhKW2/xV5ibUBlmAhZtGT8GnvY+owTMawAjSs+oG0OTgMT7ctj3tU5RM
k2Xu8AOf6gugTbceI1wy7kbS2UTyesudVd7P2MUmzOquUWX02M5sYm0pG2cbMtl5
ItpZv3vkMJShqZ3rapLNrRcWBb4ErscYT6KjqIl3MOMpEp0MR61mqb2wm5GTU2IZ
yyaee/1rT1Er9TJbI3ZjG/YONo28ltiP4EDwQVONxrQs/whP53ZcA8AnyK1wpDvK
WrEqYMDQgG0N6SfCddeS5fFkm5wMrva//QjHXdjyCZ5ZjHNqlXkfjtWkyWXXLwM5
StykweuZLk/MLZDqqwiCV3bTuQgRoKI/Nv4CZsK1oVZEl6Tmj9bLPyyk8rT37emP
M8TE4CybH4a/Cb8DTLBvZ3U3v+VT9yB3mkRXcv7gTNL+8S6lSQjhfKPARkzJ3baZ
oUuu7/AajO1CXWFr7ZSgs78oQcdm+1+aIyvJy6LgiS1PEuysUkzgouG/RXka6Non
50qqFw64gV9hUYAVUmE/uWgXnfcdCkBXYHULtzbpThc1SZ1jIhG8yV8Il5/lC2Xa
IDNeIjT4wK+27GszeJPt/63ENNa+UMG57yDhfqBDDBEtUl5dPP/tC7eDPFyTYKgI
LvBo/TGO+DXB6Pbg8NqOmz4VoooMoCLEoILn9CbxGHlTM/ZnKgBRYUELmRt8iR87
vZsBiEePDVYLtbcR3IjecHMw9vW5WBJpdz44FOHsw0Fnv+bENonR5DNKXU+/fprQ
S7c3RcSddCPvJZMRzGuVHhy+GFmUM8HFs16pBfl769fgrKXa4H+H+eus0YVCCgXa
00fBvNiioHAdIDP3Ob1rQo0oXgHe88z/5CDj+pQGVbuX1QQ6HncNnT5AI1UScf4H
ukLDDTeMJO6us2iNGLuPnMivOjbfgpQcfHuFRA35uhLqAE/8fCTxVejWZsX6Jo9p
JZJYw0mPW9YzvdbGvYBV5kXgIpaUXPXvFp72dnhd/hxIS3ts2KwglAID0hZobcm3
K6ajeNMQRpD348JXRXWPi3Cp1dszEZb6dUcGypYrArO5sB57RmQPICROiM2RqLuy
wofnRHON4m9A46qmAd8CkM3R4+hyLz2/arr/HagDCN/ZZ9oFVmXb5/NI5ZEsb8T3
hvlBRDRqKOIfemZ5OaSv5eOeY8N6mn6GUScRZHpSbKlm6+piZ9rPbfdaPRVEr+IO
uH9kxHoe3awDB6G3AvqZsWPY2CRPW0uHrlSaqQ06NP8+hZciduD4QtXkEw1lFaJz
AebUsRMEP3vB6XHcCEF/nxKH5tCevarcSyJ4kpzavkRwckMSKIzVlnTZ7y28Oxsi
HDWutdFL5gW4yMyVjVnowZrsUp2QmRXiG/BZ/9wz6lXyykOZXTSpgfxqWkkRl2J8
EslFs2JFRhbdJLyT8I367USSYIpnaDlb+hdAm6EOGLS8FbIuhJx8PnHPeZs98dXv
fqXpfOjV8nTBAX5DUI1lXHt/hETluFpUiqZ8OTeoN12WwZHg/u3yUsgrrfl8IS88
LltERKlya1eMXOvUwxHH5V2hyDN6YT0tx5MvwEdu4Qos76Xp0j3kZAAf+pAoPTiM
ZdIWbCUqIf5UyE/QYcVwnJwLnm8Snee9FlYioJrgxyNHhCp3FG/MJwTaJXb7k1Gn
tIsnqDJqlceK5gPtGYmkzAPnC8OLsNydNLsD+mFC3RWPL5H0wbZgnu+i2BNhe76o
Dg/l8OtSk2wtnuZWhACNNOtPryf5fROL3sr6G51p4nicsTQWnpXXQQiGSmEAgAd0
brRqKzPScreHiES16YJQBBq0EVoe2EFSUTO5fo3QqGsTX8p06UWaM3H0+03ZdryE
bkrxBQU/PACq9rO+2AgnhDinBmoxVhIihVQc2DNH+nz2bW+3IVAWuGYDTOoXhsxl
tVKFvZeYsCj1tC26XBei4OktaScR5Aa5PaPipS04SwN+YO9+knYKxsTphydwUQUs
lwtGW42UwalLCnLY72dkzDdkPvmHNAo6eyXRLjxAY3REIaBRC72TVdLd9XbxW7aA
CyfRRhkcUvuaVx84tPE50QQ7NdjvKAKtoZzLBHOnA6wMF3NsdJrPZUXVPWOnqek/
Xzm9fCqsEUvdaZm5qiAWv6w55GlrZddlCt8kRSVJALrc3mIDg1uJw1UQKcbsL3SY
PPQV2MvrpW7PstHC5tg1JNVcmCvFQygDzCv3FRsA9iUbfYoa9LSn5hhgWEAIhdyb
z2YSAwKO9xx9+GM9gz7E6GqQ6ejWFiLKjGwkVxHPadKmRvcC83ttxq4VZO9sPCUo
JisohwYQn9/1dDQ4EP3ikpRkhtikzxQ1CcT59eL05RxveomMFl2+Ei5xp0AfIX2u
cppEQnyuv0qW+lwYiq2N1uj7BqTsSP9coSmaSNx1vkMXmsHcWGGbK+7m+YAhV+UF
PA2/m+eTt8wZgmwBTgHKoSD5z9Nc6+RzWV7T5DOI4NmGYEECa81LbuKnB6aSBMu5
zAb9xuAAhw1mFr13eCHGzu1e2eoqwT+XWFBZ/1mHM2PmuekN+jSaIwxo8SjOlU52
ZVzRtSPLaJDdJ/dj6lxBnc0j0GB2W+vg5qUym41HfrNiBNJ97VLgvwO/uxZMQATP
DwcClAq15Grf1dVKDn9oHUzgRbwDFv9eJoWQrweM8KdhywhaSS0a/9odab1z8Rd4
RisOdX6idYwBwpe4lmJ83TB9r5WCt7w6ILVD7kjhnmd1/Wh/Jx7QE1xCEPBRTvAF
cdsoHPytGUAxlVkoTUE1bKiHjrW4V7kPVHvVSGbLW9dFE6yUMf+f3cq/cmF+iMMp
KbQh/3htszT7YGWv9SzhMmnHsWt2eXHAvoCYBAJjlwA9zVUUi/Ux6PAUIWgtngus
0IJP4MZ7CBVzpvuPR5sIOtVYEyb7X8m8qpn0T3upaxLGMEBXi1UzO8M+/Wxwwkuv
R0Igbu26ZaxKOuCTeGrKri5YmIO36NqjT7991wa5g7l+LLWQZmsDkB+xD76recBc
1aOuU39GEXfxkPPLKF4WLDpRCM+W14ZF9aqlhjhBQnZJ/Q9ddoMW/Yus7Dy942wa
1I3yrhug1QuNUuDVzsZZs+NhVTjQQuLnNQmJIcK4TxwrCiMXFJfjaZckKbnkB6hp
owtfRItxoc3/grvGlS0LQ06rAC3nJEQgxeAzPLSle7jPC+uOUdwXONojqKOuU21l
ENjylIusi+n0MDXLyjDDXClahTgE49RtMP76ET6RpuoTRMk16UUnL94zk5vRHyXH
A/z2XFkG5Pd9wK+fp4AKN/E0fjiZckJosNEBxZyRG06C3WxGY1QL8LUpLMQbV3EY
KDldKFabpov/v3xu4ncrh6sNM1M3gOhzSv8vW3glWNvjpOIoQPAX+1trdMQHIMaa
sfTy80UnlIukg5ZU0ezzXzIDjAVhDF8q0psTp7Hhz0GgDJmQhbTPuVwigsE/UxaR
kGvD0/ef+PfoANWPA3jqLp/guw70jax7PdHIgKbwymTvcpgVMa3bAwGg1U9lwlbH
SH2ybl//FtgrjfbENz7Cq1UGYlg0iDjNnwlm9FLdZ8pv20ei3DfHMX50nc6EROP0
i+4BoXKpdn79dXzevARIZ1pPWeg+kWHYI/XwgLHLxdti24m3WABb+qlxrRzY32Dl
OxUVtmDPh0acUpLOtdHU5tP/X0OcrpNCGWoZ2lhCx2P5EmKF+9lT6tFrtQC7Ggqf
rZgg+tSc2xbNDQql52AScRrAHfbMTFbJS8LODc0PU3zmweJGiAgPn9TGgm9e7mSA
WEF6IzXUpR8GW3R9J0TcI7y4rA5vtPGVU62ld5WrpoFdFyleg/LDoOuIHDL2P4Fm
xg1RJG+YuGZrfoB5CxFJgTx1/MZH+X++tcUHGp144ZIcR7Ou/hFDUCSJ1c/hKnFL
F6my/jOtlaaGBgf3H6qdGlqDaAp674OA2NBCHHuzEopgj9vOs0lyGlXOM/kBy1Mz
egrTAzihh5M9yfB/OsTYEWidSwN3rpt9zPLRpCeVx8O/5rGxTOd88D6mbvnDhd9g
YcINiTYLNX5plTbKc0xbB0MQViLeXf4jmgiIxbKGyRZZOxJ11z01zMKES7Pd4hxs
JscdbOJgt7VSWip8KDF9MKKOHjQZfN5raHTgVUgu0ugiMsWZ3qGiH24XWGEF5gkx
LHj/FhfJ2kt+k9+NQI1chaqvv8l1Isf24T1x4QQAtsOco/rjAmcU3G8IDSE+WlKJ
4MVwO6LClpAjUVmcPkLO5jta0XDS2f33HebaGz7HH/fOPDHZIFz03DvfQ2zYzUZn
n+Lckce+n8/6B5NFnWcXXC7+/po9/2wwH3q7JF3gpapkp+QJqcrTScHbhYR9X4jc
YDQwFAhomdnPxqa3vFuu1Ftw+3Yiqi8Fu2SBzWCkOE/s/pxM++QxoUFk6S+6iCiD
wnN+VkLhlRzko7aaLE+zsb6MNt0o8hWxjss4ruqAvCkSd9qf5sKSi4yblNoAVBPu
fF0zsuDHWH+n9eQAIKsMxoQpUTfcNi9PlYqQq+BqgWogb3Jz7hH13VZJqGc3/xe+
6zF+eQ1XZ+aEMjru9Xd/Iwq5nfFwv0Rx++f6dl3wFgg2fLhLzt6GPsARxellsJpg
zAB95jNi23cb6Z5pmuKvp9JaThhXFnkzakJQvBVBMYAt38eENR8nYTlYzITv9ABD
XtxuLXjJ7DYJD5XRLNkqbLdGQyChD4xJSgaBoIuft7zRu0+zeqqCV14bm0KsIP92
Q4mhnVl+4iWwum0a7VHknbGopGRwovxZ9kTCjeXUAB3lyBUzj7wCZ3q9iC260IZ/
yp+LmC4D9L8jauvexyF/azplIYdrL6i0Zl5j9TA39GSjvTNDuixGE9g5t3eqeTcH
v1N3kMnhD8B+HagULtZTsrjveSMMzF9SMkLLxz1ikHrpKyz7a+yCHh6Z7XxNM2F3
N/Qt4Hop5KLjrMvoVNbBi2FajiPGRJHIpuICNzoEmUQknFWUdJbPkfXO4ovJzTyJ
+52yLst3qzZ0Sz+dCOhqsn0sVyTU1Wd67LeaYHaGmgLlcKX7+uUIF+rQJXhl1sxh
S44NHwhQ206SfnnJxSChtorsv3NM72ebckOkw40QGe0sZRv4g+EC83q19CaQlsyF
6759by2Iqfan1dQkLDDkKH1GKEYd4hol3CBJhJywWK81eisGDz6B/HWa/V0mHm8X
mBQTRc/WdAWlZgtfZbFwUcicH5IEBpjSsNggIaUvqN6OPS+RJfiy0LVR7NkqsRJq
g17bv8fuLZcBf2VoAu74WTKo9dIv7BwjPJqv/whV0AnrmHryoZcc90t8poU3TtIg
l+kPbrv87W97MJMK/8GuWNiawZB3BT5yqC0wzNvELGtTHpzJdaUHtFpdc23F2sy6
lAXnJavFR01hGWNiM7ZPfqqNflSUMLLXVJ4HzcIpXcQ19d5wIA+HqbelFmhZOc6f
sU5rl9fFKP34i3RFPNSVIcf/VSlCwLKAyQ5OVRRmSbiTLz2fKuHNj4IPcSoV5Pbu
OTs55hOJpd8NRvYDZHzlU0ZEaUmEoujfELr1pLHBxNGTUPs4ss1yo2WjQXlTFu8N
AeKxjybe/AkPyZieG8FfG3TUtN9aaxCc16NhMGjn5la4nVyRJXrB6jH1i9PZGLvY
WpQPyY+y8PJEP1Mn0t3u8xI7CEmYYb2noeph4r9ZsckzKa7+sQqxYPiI+9ZzCkZ+
pn2OlMpkj3PMRjU1v258Tgt+RvHq0HML48XOeoWY4u1d08eQO2142q21EjRg7OGZ
QbYRkxg2n+zZpVugnBTGoEGUdGUUfgpjLO/hIBv4PjaTAQK8aXHHoXlwoogyMiky
it2NV5PZlnW1e1TM7gtgbDH1WMUj8HvnyDSOVRBpewwIjQqtvkijzzO4TxuAZXU+
LitRdMe8/SxPtSltCJ1olkLI0wUELJOQ3d6zvYTbnkIBH28CDl1jOk36UsvuypRW
RqTXfCP5uLgS2PgUp9AAPeFG8O2KCi9NLV7tWdtzTRam1I4Cw3bPAcXBJINWnPLK
tkQB6ljvGwdQFg5YgMUO9UiD0jR7xRKl0o3k3A0gdHrQpAb3atmNZYJFK0XRi7Oy
eL82CFDTjg8KpYA4amfWsr9u30RW0yXSkN72jPC5vAVdYt9+33rqZT2gB8arcT6S
wIHec97Tvgtx2+7NfXd5pwKFGFHS8YwJCE7tNASI68bhNroVszcai4HndZNadJ51
v32renxydPOv0M1n07aKQNxWcCvbBSQhpI4bFKZnFEWSoeaoFIrAwJzkucQuJipY
Et3vpBq1rliVSESwahJVPxZTPCZmjczQ/1ASu+DzpZHEJ1yv9x+xne9qHKTYn7pH
HmnPw1lBq/pAMIu+l8IKZyLwtxUTtx5C9NzhCDDVkEhEAiSITSbEgGACbfzdqVf0
k1ObV/RS25df5u48jDYV/x6SXGps74VgC9opMlWd0ttwBF7nixt8LCO4TiVrk2A/
6BpDt9aWiTaAcVwZLEUbJmfwBWtasR2c/3VDvrhHYoZ+2JKhVCyBh9joE/RU8TL4
HNcxRRTQgPK68pEZ/ih1mAMt8x2hrzePBu16L8Pf0JP/RdeMeSUlwYrPLMxVfDVe
/hYLZACYL5GMJENGdsB1bzY0GX8SiA1hlezqod2FRgUIVi8mKvta2Y66n6VdUOb0
Q00MRkSd0yv/uBfO6hoLeLka8wfXcpjFWCWYrlE9kJ7yygEbf8OXEv73IPI0zc2m
cLWUQB6IPpNXDp/qjh7Tgj9w6mtUgc5YY7GqZ6DLaTma9nRyw+OcIi3LztorqBPi
CIO4Gwu19MzCdicQUKfv8i50+eaFRChqoKHXwAyrsNPqiMAoDO5D2KpN5vd9gk0T
rx/+w11ceMzabBNh2wxFbFKcMdwsIP71S1NI+8ycVl0Ruwo+WaznxTv7nkYEIkgl
tXojfRqW5CHvUPuss8s0n5CmkHE/VPBi4dQdMKcx+kR/8MPjhxqOAE6egan0BAWr
kKTXFW/IEmHk7gyudkgVUFCXf9qk0xIvqWFUj4Sl14Zw1mTK990pl8UuG5S6qLX/
lFgloKGQTr2bR+4YZZVQLfQlpB7347B5319TNfO7PvOM53d+nPTxUr4CoScRrr0/
zk2aHR/90CmeZLvoTUVG06oEiMQc9dQwPfBeY51ceaUwH/SGVS4vNJIkzm5Psrvi
E4Wo/leArqgQ4SQTynesUz1vYKlV55H0fHWSLQSrutBNKjEp9pikRH+2LTtbrkIH
AcncKYA8njDWIXFNHX9n57wvy35rrkWPbCVCXz/gDkQDX5qmhQ3UDHvYk5mkCmcn
8ZhH7mikvxWhx3qQLUOq/ufRZpqXN8VUjaioLEVnoZTZNN4qWsR2n+JjBlL1t3RZ
UVTR1hP8CtbR6f8ITc/A8Xjd5kLXW74EZm0FagFrdIQIoYtgg/hdOUBg6HEqHiAW
yZYfauVkF4VvIzvBa+RcvRrL+lGkxRR4rLtZ+tu5nnnXo1GAG//zA5KOk0/Nh7uj
H0auVnKg9QGq1JJnnKv9oOWJqd+HZs2SqdjPKaRzM0cMdEflPaRY/xfrUawKu2WW
Gz16hAm1id8CM1ZojHM0vjv+UtRXYNh48O2np1R5zvCbxyGbZUKZI1Nbz5f9zKhC
gtvAD2x/hqvQfaTuspb+MJ58uHcWzzkrQ4sJH17Us0qNUww+wTBhRMifUynr3kCQ
TJcB1uGQ8zrXXMhol0BzY7r3fEd5MHF0WZ4anHZOmUO5PMcSHJORpYfOZREv1BLe
jQ7NLlNGQ9H7ZVaqL340coYxgQx3m2NVq37Zx+SuPGqgfzfXhAru2uHBhDJy/QoW
TLyVTOsZU+3E9AUfAKfRZyLXtw+9sP6PbQb6kHzVVNtuzjF4Ao2L1BUm9JWyRxdw
7WSPTVW5QMWplML1OXXWsu1QIotMf50tu8Za941KaLwvzdfZQDeVFuRLq+24FdVK
asyCI3dJzPQ5Tst24c/2UMxIcQhuTyXhXb+/+oWPgbyPX/bM+GAl8tWlXbmgzLrE
+/6jts1pWKsrLOEpJ24XQH3bCr34KPBoZ/9zj3BaXklrUF/FMqYNvMA0Va0eA9Kt
h0J6YTIXm22QAKSnBl9ZkT6QEQ6DuIatYrXq+y7AhDLcXHa/ASJVvouWkAZvWXOp
7fXCTsq2EFGPuaU1taxXovtJAyv/EUv1Bc8nmlichVyvNHgXD0N5ZztRVWrdRxLh
3NeV52SEvqrXtsNTdpKA3etmqAh6Lw80zKticAaEFPkDadFverb31e156hYSbXlO
Co7ef7hwuBQoDG2DPGdquKe3xfU8Z+AK5C2mN2CYHXwtxQkSBBsSVM6ZKO/9Nh9K
jmGHjXVFGFKl7kaH34T6PCbYnZVwvp6Nz5izg4lIQDz9UzdB6VWTqLl6+n0WIVwj
Ye0DuChe6VlG1ku/gQ/glgHK6YACUTtYlaNKHoNsjVZYFaOT42/k4gKzFHX89Kzs
eLFc5S18J4rhYnGqG0ruXwDW/KOpb7Huit8NmXC9SlfKom88yDS+EqM8SMTNXCRQ
92q3Tf8BJLiOwkbX0tnLsK4xA9ipYPsRZQxS437A9wjj+hL/3VPZPWj2ixv/Gsej
O86mraSLn75Pz38KeKPe/bLSXNJ+1HjwdQWs37ABMIkLnb3HZ55FqZ0NxVuiK6rZ
dM0DRwwpJsBHc4lKIevXmwHHzYJlQH+6vwD/cqEZzktMrBY/61ztmSrXTOHIeYP/
/8BBdnQqaH8wwUhI3oSQQ3KDpz2zgi8O8sx+KMYoigtvjLCy3wx7QjuJz6bEjG72
uX9tbUQSoUsiu7RcPgpCAjYOVXbF7z+Jzpe2BNPsGmX8xqNIAKbgMUhmzryoG6JX
tG6iXQRaH6vY7TmK7KPim7b8ect1zYjZ3jm2regSFDq1/tO/SBXmByD7NZhhpKD9
F25cePPnXcqp390FbNPC3kv6+SVAkZoOevwrLA6I9cFKIuXd/LJV+A1UaNnddBCD
cTvVk4FXkbDeVVI304YkGycmOMvOIEvps+8z3e5AeYXgPTNV0KuwAFaJ7/XyIprK
t+gvSZ+CAbr/NC5tKbvneJpjDpZ/MH2S6d2YGcwA719iTmWay/bmI1e3hOTv7lo7
iRz0ybdM8/SK9ZPm3gHzzdkmwuzcC6zyARJnyCL8OjzlbMO2Vp8HXTRZ8PWzFTRE
UqF4afiOD7DdaAbfW9oGLHI1EFIpF1WQ74OXytO3QoVPK3V0unCPXSQHV9GCUMPk
1J638/0n7SGWW8asDw9YNhRxU/0eStI/ZAK90GhlqcxRD8vQSByKWfZunyYfj56W
zUMLs9s5whn3IHjpiKxqTS9nMO9CmR/J3XLrPOpP7v3gYAuvuTddFT9rwJaEzKeI
9goAqaORSkqlquJBfxyJymTxPwADiP8r21SzsiYuTHJCr6F2DQikTwigzj2iToIs
BEtBwAnkLN7ndB6mljuyi+pSGz5op0oYE4MZS5/d9QuzbKA8t1KVy0lgu0pjvZBd
p5yEIDQhsDd5sIStgKoZiGhDDKFBmyw5qNYq8PvFT7ifGPQuKpq3sQBuYuIeTjX6
5+Lzm0UsFr/hHRiJKYuNxhMjc0SVUv1P3GJBHbjiWgezWwouNE5vdEbb8PcjRiTQ
HLf3k4wTx0ua4Fhs08iN/1TXTTg7D4fxb24IeJUeQNCb0PLPCVariDaktYrXo8q+
Z2gDR/1vGQtHX7RwSGS2ch52v/mWKuWsvT7TWnl/ArHhNWJ3WjaYTbnYmvl0U3Co
ppvVdKAYfyhM1Uhdb1DBpE23bEGBhsdInhGvbWPQ/CrpAfVOff4k/U6wpcm4dO0M
nTYBhO1QM7xXs096VkQBQBypi5xXnBR5dPN9Hok2TIqfFAycH+EfcNARXEyniomm
zLq/ElDIEAQxVpKKET9h/BPbtXdfylHWmsobANv0AcVIIWS2M8AQOzx8dvGSrfNt
r9sYrvx+0pPUzaJmu9uYuqWOyxS01hnDX+VeMzel7Fb3ZB7QCnv1m/83pb35iofA
7IuJ6tj4dW5IiL9MgB7VZk2QS2tVDmxyjU19E55ENKPwLBoxuEOhJIp7jkDl7Hom
UWcyu47DksJVs+tZ0hksAyjexUQjbqqlw5STfndDjphI7YAwMmJwZlc822oPU2/Y
ckMMNJFo+V5utQap7EdktPFpbr73ZmVJo6q3dSBeTmYuU38yDUge7xnECtjRTL8t
X7jkWpwHwcds9RbJd0T57VQFzdsVysczqPuJC+Fhne45iVTVHeFwzE8xWz82H0Ex
ap4qz6UMw4HHC7/rvuurAQ5/QQq+jMGpqPnmdW2WXL+zDCzl3rsx6+nVZd5BckjA
djfCG3ADJlSBL/VcydYR3mU4NdUkt6t9UfTigHBQW9lmH1clzCkWMZ9OMkvVBRtU
rUiQmqNrKWFbtk4Kqa0QspitBQU0UjZElgz53WBcVRK3UD9CVZPM8fM42f5CJ4uk
VyyUER7BHJdhHw+pyCF8rUaZe0c2I+UddyYtTJ90vhdZAGtZ+fZSasou8YaBlj5P
imZUg7JXD2Ez/uhpD5CpdagMNWQTNZyzSpdR+TjoJ3yzLvQt9/lHGo173gSd0wU4
vmLMnf4ASVHf0JLMkIMC/M7dhY8QRAsipYjLd85ibQFHhyIdGBp4IREltNyT8dVo
ENpZw0hqWYH+ek/3btrqC0eVX8x9ZSCmJaZfM9FfGNLxS4dVpENyVuWuVKnuiIB0
+nXVIvE5tiFb1aREh5Q1M1sRwFB4ZKOnRuI7rRQgerA5mV92m0Fm7DqwzRdInwyB
jXvtEFf++iyocqQLOUv4xeANY/BhcwLDaD4hVIROWCCDKwqKFcmrcqfx0iRhga8G
tbakGpjbxWksI0XUooAeqcRcgXrKguNojZOgtZoE7Dd90hQNewZFnC/6+ph5rfik
amnjc5m5sgs4Az3HTQmL+jb9bdnpjNm/keD2LNlBSrpjir8VEquKgv930dPssRyP
d+r8uDq5up7f2kxBJ85RMy2Tt9VQooiEeQ0H5JFEFz+o9vJHpmBW9Q+TAyOXRUzr
TGJispkF+ymq+GpPll+D+Lfp6nO/xzW23BSNhJtilOfLg6aVcH/hj6srtcZjiBBt
9bTW0zC0Wh1FOruiIDU5xebqFWMZarvEdeBOjV6sa94LdS8Is4K4Rq3XwJZukNJg
b5uLSoJBE8lQde6BInZSh1Rb+p0VPBn7FKCnMYKdNzWOTstJDe1dMTrx3Tl5HV5T
tjk73qFbdMiYOmitCcULfAqjfFK5S65cx0wPrT2rGqG0xh5xcVyb2Qh2GTULAj4k
caofPhtyk24sCfPVM/d5Z1wdy5qJHsBXA8wc7Q/iJ7LPC7eegaHqz58yf6Mh1fEx
o57m6cwIS67RaVPyiOo4vjeGoJ1h34E01Fxd+xuDJBm56OVUt9YdMqoSDV9flhsf
SqXBuhyAVY4NcSne9xDIBGklPoH8hDRO2zKQiRw4H8sFUZnPxY5Q0wBProCSCUCh
y6Pijx8/y5WSQSGfW61b8J5Nf7ElRqjsiqkHaV4oyGa3noZdne7udnXUM4EERxDh
5sc5vso485ov9p0MKnnLZFmBEZe54ZqByBdHM4sWrXrGqRhL+ur2VGiuoG9Muigp
mZlCgGahbhIlwdHoy2UjTlk8JFwU19VgEZhWFJCnAmRCg1xCf6XpKeCJiTxzx8Ss
dMu16TgWZTRxTeJ3ro4nkCoYZcmiNX6oGwBGOxQmKeByAfkvvKu8pkYg9jBT5705
bbBW3NbTHruc1CdwN6lPKiZmxJHxaMVZeaOLF4lTk3/SX0qVhZ7j/dlu2Qtfo5QT
ZxsmgYduuvUoRvcsGtAyJBwg2FMwRmQ3L84HC/zIpXVEdJ3by3vdJl8JyK5n8yma
RXmwOmAQJ35y8ntsfbcyEVNQKcDOljhJ6L2EGggZc/P8XQ3A41C3kWBWNFqBbnVT
oxFnlosRc9TRAsGe6Old6pwfypNZHdaKHpyS3+OLRKBMAafjrHTxu+yxYw8imsY1
G96KF4MGQ8+CZrKtDhbUW51JvnDJKKFogIK34X08VP/IUxbay++kAWEQUE525BN6
X5KWvh4eE2exh4lVgYOPs4cDhoX4rPyD4cXluQedMKoilf20jWTrGtdw1xpe0krN
EuTO4ExfiV+zxyJtC0j3M8YnRsk0oxGwn1kz8Zv98HZ34cslDPnkFRosGLYtjj/y
4FSmvle7491fe8NSqpQsAidWgmd+mSC7oV0b8Xytnzpbw71QH8/8kAQBc8Vt2JK7
7srp9+EkJvn3AMQQMCSGw9Ib4ts8ilwDBKK6ZdvwDiAGUjOcIgFcRRMn2bCc+gdO
9kWk0sOwzQ8xeI3zmRBJGhoz2CXBzNtLD7ay+iSx15KSePGdY9W5zqoyy21HDyZr
+fadodG94DahuOG+D2i6TGPhRRlZfL5B2fl7e3iFTvmRMSdGBW6Ye4JKdyo6LMOW
w3gb1pvbiCcpmAU2VBBQkNNIyRPgVAy0TT5qJ8azfXdqu7VdnggtmfTvPbfNLAcl
KO6/1TTSB/QJ+h4uqIbSshKHaNDITV0Fi5UQOTE5mQcuHQM8QZ1ltQz3YGDWsBCN
7oSj0RmjNwts2T3a8rC8roZPntxnz3qjFKZT56Ckrb33aq+W1CmFmSbGaXLXCjsQ
DZOa9W6rLz0pEMSOy2Iu8PRkW6ZQe4K3hGf0Y85ITUvtvOsG+D3+if3L66dik7Um
Rl0qoGmAz0UcNu3ZbFtWdmCarMDX97ukiSRExPxZS0bmKTMBICA9sqipuwkRdBHr
A4yIBSmLJu8QxLEDSg4N9bLrxSosMp3klvmg+uU7G69i3zRoZQ9jm8LkfmlQCGfB
E3zK3vq+WGDqBTlpZ22+MlyWui6ivRna0TtRAikJJM8GUAZzmopi7iIzzCHVrqcC
kTARk3JKR94IqePBz0BTEwdTN7fPaP3wq9Yl7G+4UiAcmgJCSH/iwZ7G/IdAjOvP
yoNVczijjejfddQOAVFPOUV2ABX0PBOGYNcFZ4+Q8ahGO5p9u7nacuEaXDGbF7EL
v4Fo05gWC7GO7ADZ4cj4YB66MkODeryyqOUcXs9aRxrUNuMSYOUeMUF00x6PHFEX
WjZj1PUfmooMiFWU1Bq4eospvBf0ZLQOhet4kxbF8ezsVXvtwuL15J9Gqkcs/oTE
X5AHXoYDA9sf0BoGCgwQbeiJK1YG5g020Agsv5mdscPoeRvqb91PmiV7e11H6cQ6
7SNW023ytK++ujTyiH1xAz91wxLgx76v/6lF1IPLR93PQjcSJVn/zGl3UHFI1w7P
wtmoGuGHZ+gRgoRgy/kQdC4Puo8rT7tq8AZEh81R0lWUTG6PPRI83JQ1u/obsUjO
1JNHTStclZ8z+dfoKqbE2C0ejA2fG0KVeDXgBMIzzY6nkkel1C6wrqPab0ZjlO+x
lxXQsM3NA8XSOePXiljLGf9EelNoY+71F9/07CiPyOKo++qILSbeERXghQkxgvuv
3fQQW0zy11kl9Hy/7WQ+ndrCCATtgip5SbeuBZIfeTaBAfjLMrreWxKLPP5aCNUX
MCC5rO8ttoMiKYDm8Iy0otRyryZdQu8/iT3XHNQSaWTgb0VhVYRXONCpJBows67n
cWHuqspJTWei1YjQ3bFIB2Cwfgn6myInrBjQ0KzIBrZ5jnTHq+63gs/0fzIwqQjA
xxQj4TJBHhLxRO8Rrgi4sBsaP86XmvSMB7zZeWPkE22kjEpd2chdYMXOARH7RW3+
2Cfgy8i0/giUQgwfrwbXh2cQYGMU582dQwz6RKJT2s+1OX8T45fhIsuTS5HJfDlp
ypwLDyry0WpZj9Y8HT+YhuBPQJHBle3MP2LkKGj2nVrIVfOIwrVFHGnHmJoKaDfz
IFux2o3AWd8zEWgzy4vqqIoXysE9OUm/rPmHMVh3rAJYt8gcw8ckjIxxXmzUJh5N
obnC+afyIVhigmNOy17vfKhNqQx0PnDKbBELmVzQI4WX1/teyoTNwuorc4fOpVqq
2kQhIZWLYj7SdDbIPNgv1ZhkTpR4KQTo6gd2kupTGrOdY7+Qr5aWKwhq9+9zhFrG
wBLxFib+yYKmK8RlgqEnY3syNzP3R/rY6LWz0q0aGfiSLFq5gQ20NTEau0euJWzY
YqlYIY1wHKtcb7TV6M6CWg7aZD2Ir9osJ+ObAhIRlrUtlFDGXXtkbuigOQwMBJN1
T0Xy0xgWhY71j8ZbYODZbpI7j7gF2qznQx4aYYEBoDORBZ8j6pWeZgkIRMbnJNEK
NW28R//wYSpZGrishAnk/LFJhkEF9BWt5WwHdm/oAscyEU3GOIOlAWkvK61oGdks
l0MZCPo7ZJNJd+wtZv2Zq1ft6kpz+RwlaSKaJK9zCgAMsJdck9gbWPint7NtZWoE
MfUnj2fiz54VQSS8cf51gCOV1Ylvw5E7zkc3yOqGpphhtjGJQK+gvsGM6bSZULVt
4gZxLwJJu1MElYYHIw71OIhimSGXT0w1REJMRs35nkmsOzTZEtxp/L+mk4ZbOnpw
IS9YofbttWsCUrzck4k8e2OD3mTUjZf8HaKhaTANqhPQ7sNtlDx/cqc8/yatvNxS
vETRnGZSJkPsY5CgKuFhrCa0lCouqKdUHYJgqR8FtXabQao32PrVF45yfJO0O+pE
xWaDQ38y1QL1lY3MrJAcaFUNwCQ1RTulWQOcJmNbaqR4m/ewOm+LI7cvkoAFECe+
uClQ5OhG1dcYeDHP6NyYyoG/B7BhQrs1MFKhF8sklq68k82lxZp/iMhYJ5JbqVRc
lYpdGW8gWvzeQFSw5X6h/B+hCpiii3WKt4z+1cUZQulC9kHxJGyIoeVMdV9Vbd8V
9D2IugUs8iIjIoM726Sj0NFZigPx7O5fMsZTauwhx9wx//Ek+KhGVWjtXAtpcC4Z
zp6e+6UY//+kuaMmQRropvah/2SPGr7GNiN1vl0H6+gh+5twYaXSZMJD6JOYp4xw
rKwJsCW6xrsvWJBVYOS+g48DR7n99dsZ65l7kgtbz9984agUG5f6vz6MNVy7esx2
MxyD7N6Owe4Lsii6toMdcICYyCWtFlhzSVjPyUmF8uXVEwBPvvobBAo11JbslVXQ
oC0rDXUnBQnu2IH2YeJvBhwEvR1KVyi4YJq42OaJIhPEJfw7O/9F7cjDXImam5Hr
e/qoi1/FaFbwjayWOVNZJ1XFKY4GWppcl+cgx3F/QT+jRS9CECup6Q8TZZfP4kLm
jKA+dcsiK+rT7ncSbOSB8Axb46nKs8Fdj4P9c2LoMCQIdrIGo7Bxjb7wz0A1eZso
SkjArtesYY6ODDU/k+lhtYmy2UqQr/m1plww3kcLu2iRHLRMl9xUdgulAZBEZ3AV
QmhbNKW8eRSm5gLV8RUV3ogI65qTAMecxvWofb3Uzq5XpJA8wwJ3fMMC5KiL2YM9
JdBnnpuEVzr+LNDHsJWNjzBJfZZXlb9JdG5ScUNAu8e1CFg36+vGsAUf08tcM5Az
79PhEFsZI0GqQC01reOQFLdcZxOfjGE0aR9iblxL9nDV7WRPW553Rbuvdz9Yfx11
4vdACKQv5XRr12zbIiLs2wMggHV3a01W1gNO0s8rNNv0GeCjDRhamQCZqsNyY6JI
JQGC+aF5PtB6eO6KZozkMSK1rEudGY1hoB0o0bJZ30F0W8ia94gKPD4qKN5aHFcq
tilJaNcPIPSa3wk0F0G5218whW1P9axSmnW6GAndKcUqExdJtE1mO8aDsigVdSJC
AD0W1YgVwMy3JZbsFNdbm0SOo+gk1l6BymjVADFjC3+R56OCpzuF69MHMSLETn0A
qQw0PyV/z1Gd+zHgqDlPiN5Qhc43/z0XFoZYHRaumfOI+uegTmis6RAC2TSeOukd
UL+lTDitcGGQzmfUGurUZpH6lshIJsvSvpBJH3+ABECuhJz0rf4AqK8jmXe3W+2K
OIk6o/+dmkdz4k48gA+O8aCbPf62ACio1TymrjqAbFKuIGSZNk8CPYwccrvMAJ9c
TKZ6H1YvnkYHJiyYZud0276FuSrqEJS53zxN+DFLmOtPyJUwDlh9FOOYmSRPlh+V
29TI7Phf9gT4nlJDkR6K7kKeBsywxTEdPFMVqBNPX3ad4xCkc8lhM6tFJxBQDRUw
YmAfqbAolTZWnx60PmVj7mtsqHSIftu8OmUKyO+dirSe0U/NQPtSE6EoObklGlaX
RSOPcm9/W8Pfe83/0W1KQLUH+IXRdKKCd4OI2/eBelA5SjdOWGmC1YUpV8dLLV/+
rLvhFBvqSaswQ6d/tFN4R4T4Gfl/16BSbY523+ADfK3Kzgv3xojvHmTmFk/9oI8L
zxuwIEztZ6EYNSfjYsC+aa+jCaC4yttbrXG8Oe6Iy9iPK4Ad0Pbbbv/8qjtdclGI
EQwFGx3Qy0k7v14DdeBj30Op3p0kvubSUS6pXlWdEsCbLwU752qe/N59pNlmTG0o
4+3Tp8d8/BlJZFNeeW/VPDLV9WKCdCMbkomKv5LecDMCzgIK8GKduxCgY79pdazO
TSI8ntKl2OWruJF0mV+mkYswdL0LZSYRocqSJ39Tgq0bFxGs9TrbDl6rcex1ls0L
mIo+3gHxQrJtIhqgXibxY0lkqUgsHMzxTHpOPs+CV4osp4rcY5LjLaHRdsiOzGle
HWkjOtfmzhiDpk7x4r7qHxygZbyhX91GoORJPMnS4TWl7EpcAEyPvwBNtRhFvj4a
QIIf6mRB0GaU1X/nJijCPQmagiqu88v3J6zCP7xYX2stcm2XYCIHp5FB3sWXqPpR
aPaBDq0kgQt8Dj408AKdfI8qPADYV/RMNIrSphqNNE+Bh4jpwnNB3GRpTkx+L4kJ
Ve3DigBXqr1b8kRoNpERbdSe05Ve87r4OoMSCn2zpdLzBEkbxLA6EbdI4nJQIHAQ
W+MnO21qxKR2aMtIOaRNHzKdQFCfpY866Zk1gAF/nVAAiyIE0cjrg3+lJlITmrK3
JutZEsUfvQ4ny4GE1ltGm/ZWv21NUgqhMbkz6HTRH4PX3DHHhLNaZhsJsu0hwLIi
VOmA05FrOeMir3mvSfNwMXxBKw4x1L8HtV0b3yl58yXoD+P+EsZMjtVZ7+cUZSU4
SjGCNztq3T9IwVdPJcFTAXJgyRCjJuF0pF5mjf3s0QyEVlQY0RTUMtoCKXQnKexK
HujX44RhRXdKMKbZ19YaQB7Ocz/dBOn1xIzSk3Yva0Z8ZVhCuq9+F2TtGInossbQ
/ajCzKcmPEzcFbtc510hlR3qfida4Dg9CXsVx2LjhZ3WOTU/agelArvMnQeKespb
ilbJ5+WT1WerM5lil/IXftz+FzAEr2k79CsWCGQUHJ17lRBd4y3DRO13hkVk3RiD
beVjMm5/xf9N8JMeZ5T4IeZi1h9cl1Fs7x2HVo0ttZiviNJnRGk7FjmQtz1pm4vG
wgYBNERlKdKsSyhcV3DBVSIeoZ2GcJw7mxgdi2unPXS9xynMMWVSSVwXKzURkpZc
4zfjn9a56ujbYyB5dWOfF7sYY7Pny0E/Ys8b5kcWn+8mfl5JrkFGBFxXaakUyMP4
idIpPTC/ORtDRNbvF8/7/v6KSfLnefFGVTcjy/rXQowMQXBo2ggh8QJK/1hkQS7q
H4RpIrtUEEoj5W6N0hBhwkafEGSiPUGq9MEHYndWGLJrIkIfQZx487NmeK9ex5+n
8CtuLks2TlZ7/k789CqzNqAHhan/cbhbZWs2+wzXxhQKQevemnJdtPT7laAT5IVH
g5D5LPKtlemxhmPPJXuS7qX1L/kmmW58AVsAcVaiEngU2CSQyP03J/vhrTCN/mp3
Sp0xiNDKoE3tf5GADKy44uuWr39rL512QwEguDE9xJx3yGjHkYd9S+foAgKqUa9f
AR42juVPw1oOoWyJvsXj7p0qCa5yPw50tiEl8xY1rSLcjWutXhDgcFtS9FmMsn7q
hP7Wwc6QBg4AiSTehBKF10D7ofj2flVih0cahA4VAkbDdsaYpiMBPHebWkRKxDV1
NjMqy+uVfFN2QBdDJJVqld4YaOvyrF+/7rrtJjZG9Sl52WmQAq0DMZ0wvHYPPvTs
OtUs2IsORAZT8tfqyv09AABf2lGdczMbfaWYro1femYYwGQkZBGTyMFxkuwJKpdJ
d+BfTbiWagHQt2HLFIgTi0a5V+I3pJX2D4g0Ztsth5mx/qZPdql3RJEAIffdgdF+
BfEX7xjqpBKK7YrovYvWodMIr9osd2n0gAujTqeBIqpR4WNPdGybqwPMfR5f6ImP
MjhDzpzQbmSaPNTX8OpKcUkWdLDJF4qh9KPuWRbDeDxOVC0DXlYr5xzp6qRRWG8B
UKEd8iE+3yOGJX7UVEITJ+kLesNu6n7+ZsAKigvDrEUvnRpesNErASqe7cFJwgg5
ecVu7aOGLzd5rEw98g699YhJtdRqASCvtAftfKCcvPiC9YgJJIDuf9zf1iEETK45
k9d+HS+hQTHQhAqHZRUM71D5UxE2XRZUWYN8Iw6AkmVleg+uphErPHuwe8y645uJ
l+KYudLm2txmKfT6ifW8gGtMX1UVOMwiqvx9/u1ZXOVobk9wBUwaJ4+V3EEzje+B
eQfIZrClOEJOM1hfBvl2y7qM6NuX8ZviDTSbr/QtqKjZeqW0z0Q+OC7jaAP2bpCu
L9OAnJ3vpddFOIEYWGe2e6c7RDGeAjgKdn3A65nuM4X4YjknTleiqYnGhgwyhcKk
9HtZEHlzTshODzDnATfL8iV9n18EHao7/FGF7GU2Y7ebP/JVy5/QXf47zQa2KQAV
d4pdUuEJm38MgVL6MxnEnDNfbuhhZt/xJPZgHKQCt/6U5XNJXZwvwsgRtIWr4Rns
8V3lWBaYn/ZLE4UrEwKniWWb2SajwYM8227TgHKF4M+Q86MuPaZ8udYdJjTwUHdI
LaC3V8BNw+2UX6cCJtfZXu6zUWGznYJjtYjISIBNUVDclj/zKLfYm0oke9ugyUHO
xYJCiVLsjQTlWGXdOUR7rvfdKOI6ObBLWJHymCW/Hzl7+opO3CNfF3bUmEVNHJMi
ADMRTD3vPjkFB7nXSmi1n/q/WOODkBeHpk1yAiw9y8qO2l6tKP68lHQT9/BS/Qbc
LwInV9l8dfG7t6qXWkebuU9M0Z32xPgv6xyeDpmw4BlRtZYTzfmBMUkSyi5ecmR6
TKt7V2e9/4ozz59BVN6Hxy9UNW+GL6ytSHmYChi7XQ2Pdvx51PGBRD6wEzeNLN58
g0gGBdHU4hBx2D7r0maNki7UJpQnJ1uaHqEG/TO2DoNXIRZc7BYN/mDK6TTRw/6c
Vj7nFGEz1SEOdpjndRx/mNbn08EuwD8KhAst2si0Z6nHL2ZeR/6jh22fPBhmuG8s
2tBf7Hu72uFx4foL5pZVSZ167+MTE4LYzaNcx7GsWOQ/nZaOrvBIVqc+rFCGktwC
m1Vm9G6aaE7SwSW0RicfSEt8nXTWCslefzrBWcFPXkgOT+cuf6jsKYLFwLN793Y/
yCLCw+UEsmAV6axQlE2M1Dp+jbIUtW0sZBQ2U1bYJs4xmMWqdRqjoL8hLF2uI8og
S8x0gPwWy6FkvtEKqNYLlUAr9Awg/c5VCuoYNYcAkUUvD4HymuTJuxpBxPePwRQg
cwaIn3J/4UCEd3peK62gtayfqoVnvNn5J67z0P9Q8KegMNlkj3o6IWRSZZhfSwib
AqYyTVS6fTZfsUOb06qt8Bo95r9uImQYq58lrks3t/ybfuLCF129rTX9NOPUsi4v
pTZR9K++w5Aogi3fvS3a0ePtFnLVHdIUaF6UCh1zl4//30He+xpcWmy2LhfcQWtB
HU4Nd+1mN8I+juHEy62RBp/FQ5jsBwipaaNXSZh1N/FT1f2gHVA3svfA3lKIe196
PQn972aRwF5+o/x3Z/VgmDdm+3urCEVXvxiIml70qNXPckDKns0+DBiW6D1I7ZrN
UxspSPOEpPEX8YcpS3RKBJbW1hHkj3AME8/CS5Qedo5EnBjpzo8XgLlWI30g5MGi
rNsB1lihRdSvv8Ie5uPqyzzwUPaJ0QgJ4VYaNfWn860Kb69hKn3EnJkgxqYA1eo8
L23AFAW8zvIezP8utg0fjEwUnO76n0kySHKkmQmF56m427ufFpMlBbg4aOM/f0qk
UeyDHbLjtzSopey8cc96qwh1Z66NB9YS+DxElD3ikDy2UF09NTDSY8759e9zQfd0
6GE3aIK81sXIGBQIygq1VMPtEa2Dp5JqacVzCjCzcIaXJmiLhoFAZZeKgedjjuG1
mVvAodoDHKpN6JgUrDSEO1nR++n0p2D7CbiV18hEX390jhKMz4uSkQ71EOkcP9ZZ
xhjg3+TsLJw99P/Opg/qF4jKmhRwUf7GXCQhbNA/Jm70uaWk8yH1oaW9SxlDREFi
UEQ4KmIzAN5cL8db07RwSujCLQwJaM8QMl0D23yjdO3pculBmEwHxRliFsg/VHV1
4+FaaFAnZmwxzDqxWxheR3SWIerpxZHGJjYBeft2ba7cK2JzyaRqy9p+UF4AqO9B
GqYfL6qaLjzNHEcah7plK7jUcFqIXubBfajh+AgXsP57Hg/+iiqrMPEWvX7t8JCd
jLipRQ3Afe9B0hy+5JkIs7+NilTc445UphoYCtrBWSLLV78aji+4aRDcOL+PI53m
UqJg6Ps/kWSV1pGUz8PCjZerOazikHEF8moPQ596kx9vSJUPAcQArbKXE8jv6szH
8/GQahK0jFlaEVua0FRB0pJE7gnKg4D+MSGKL6NshLRr1axhhwxDARDj33SlNv1W
uCvZCD1eiOlUeM8j7Q76kewFtY1uL6aEAnCZywb0b07wiBGND3VTzMjjjiUXEfTc
suCnFNVjN+C8Ph7hYvBEJa4L8NgrSUM0rpuHDpiww3sEYsg9mPExHwaeQYtlKtL1
bSvvyBiJVWbIoh5MFj634Eoc91dXyCJRT/M3Ly18YAhQIFmClKH9PBggyDZYYa/H
H05pzdswc5CCFJDSQW5cibz1KJgN9AGR6wE+zDkj4qZE2DmOjZsOXo1IVcKCXzrt
BLYv5MX3G+jP7CTR0oFiB8e3pBttZUhYOH3QLNpoFmtcKa6SFiHivSJ6CGjhLBjT
wk128cStx0mVowY9j35wFVyP56gGoSsF48BREbSJXcTeJpKddJawQhCogDh9+WTM
qLE7HyUb2KWfDZ5+fk7yCj3MALFrO0OLfarvx5YTYJWf/Ay+j/LU+3Nam1BUQVKD
PfJofaucgbRpbDyjbndQxmAQsFJ0dF8TQzWLEwziNhmEV5a+lDO1iD+gxa8R5mir
vtJEKFLcBAKOCVFvBpSLA/LjH8au/oAeIgoHmL0WKZdqGJExpW6pqAorvcVVDMmd
gRxegKdw1FRe7HJFX5z1WkrwGtrZksdXkRABN+Z0x+RzjCib0kHlzrjecBmYdvMV
Q1BM28gHph4UObrHWLTcg0YC7ePaVDoOuJzqmrSUi/Gf7krpQfDXx2cvNpOXvstn
QJGKRZTvvXEuk4jla6StQJl8TVm4EgM/xhAbnDH1UgjQ9ITUsj/kQsxw1rh4xOUw
YdAiYtCfUo3X6Nf1wypxXicMrOTa6qYzPx9gelnJxpEwwpD4RFrLgfWwMRgNAuk/
4YKd9Zhrt0aU+yfhFjBNxsb2WNzMYxzAmvPXCqViD0pTKI48cUgsz1rb73s4a5cR
1D8Vq1mcRKiyx6aA7aWBBNRnWwpquF4YyW+vpZiKz70bCxgg7p6YWQUbNLEgtM/A
Hfn7n+b1xlHqvE08RpEZK5ZeDbZQMM4bHcGT71eH6V5lcTLq9iliK8LFqnBuMrEG
o2jY68U+5cTDKmYjr72EQRXoq0mh3iMCfE0bxHzyy5CdkmOvO+hey7Y5bPN9mZ4W
9sR/2af6SBUgZa4/pNGt5tJD4GaOfsGso/t07toCPny3VELmn78jyD3HdOTubT+u
tWLyorMYr6YTW8xPi2TWaeReUdy8029zdvoOwOYI/5o+m8mQsLStnmftt1WuvNc1
fbtghckimmpKSIi4VAR6VSyOL+GxlIN5B1JeddczxNRsHVdVNTvV5ie9dsJiBD4P
fzq6ggNGc32SUz55k+bcNwibTNaRfxfBgj0EykuezwGrKnoMraaAC21q1+RgQwh9
I9E/MFtOFnhZI37+6J80BndTLbH6rijsXVdv0KnYtQijsMhnqKBZNP3sWNOlYVFr
eOnzwnN/+RBnoZ3lmLl07wr/RsSD5SwWZCJ5tIjEBgxL4k8Ru8lksGt6UhQBfcVA
fm+OZwsu5TMofaBsScAj+PIdEe3bbvx12J7HYr1bA3MOvE8mxKFB2sfk/pv92r6j
5BmM4ar5+fBZaDm2UyDuSVV+rM9Srz3KsK2HlYQ6yqp/wClQ/eJwY7L4HzspNUvh
otFhjzycYm54S8YS9WzdVpPjPbw6FCuXu7reydHI3lgNtqBjrL9IY4cJW8cwTCeT
IU24QGDYnPRLzqAz6rfMPGr1wlLplTKclTHer5fLJQ5cq08AXcl0899vXKsuqtPa
7fS7+/26UQhNtCfPwZUPvPXL6JnA5PTh0eAuXDRm/LzCOfl7B/sqRf0Q/eYumvL9
4Tq9X536NRyJ42+wt064wdMA5a5SEXVOz0uRGRXTtiqKTfEWGDOJtEcRCRCipDr6
JggkfYcWQ/NGizfr185AnqMudeAyZQetfXrkQLvMIYibvcl7cpsjT7U70YeE4viJ
TqDuP+FLcAoAhPKqlGDIUFLZOUlc+pIbUFCWMfPA8OPR7ogy+wKBr3ua5rFdqjG7
rNR6itPGbsDH7+PSy2VPARBJ+Q/jXD06W15wK+0CtU+gYnKQJG5BfE3jZu3IXkp4
8pz9rGgKGcJy9eSJD1By39JBCUG2ssGYIs8yUuxs3GEb+nznysnoXv7v5yirbKDz
7Ug50+M+NDpYoH/yq6IG7BQrRn4jsyZyw+f6EhZor7/S2zZ4Ufw+G2j78E/EOO83
+23ghGe15fBVckWN2o6Qm3wGJxwlkbZRk7x8VyUndfZRHD5XQu2WzW1nxR/bcpZX
8AvFt0xlBWbFyol/SnhG59B41qXCL5zK6CiyrixbNGuEIuSXhEk+1hLsbBBuQvjM
YRVFJL8Z7xdlDw9t7Gv0UAzun2gh4LWoaEB6WOVi3KUXRTP73jIa4OF6O3d35PHx
slV+Cuf4es4war7vNPRWecJbQxi4yz39LrOCRruSkzNxWyR1Lsd0xcFRtqEu354b
yLy0XLqZnHvxkZswIwM+I4emgTsIGbbCYwRn7VGikno0fWiUVE1XZ6uaNCxlSreT
Xu/1R7MirkN6zpXW6hQlK3jJBHQbVLWp7xve1x9S/vwtjdjICrA0CCHDuIw6k7PC
toKDT5jTxsyWHvY3z0CAN8pYtsxDrYzc1D1ZSZ+U7QZ5eOOr5Q2PTN5ZXRBJrlxj
+UOh4lKkINhYzOvixJ0J3Ya/3x4I6U+Y893BF+URAS9JEyWJCMKq5H5fXi2WBjPN
ItATZM3Pa6C/HiHYgvGxak/GtMXZQrz5U8ZqApZb4qjwCwLLho/31KqZgmcJP+R+
U/qXvo3xwJWFRVQE9X2z/MkNH7VUyXkSEGLwh0gEVc6vMg3/Hm27M/ZNf1iw6h/y
Hjjl/5JGgrXMpmqfz1u6DYz5DySrdZdAnbm868hr3S16s8YHFC+5tp53Bc73d8Y9
F8ylQpcah0YqcAjWaI4wfvN+Hq+x24cIRgSH8YlSdbXGQ/QBYoyer8N5H7bknfR7
ngSyb5krN0E5u46q54ZL/SVF1XTXMvMYyY4tmFViFdKprLEqZ3+VJjj+TznCPYMu
Dq/cbWJMIa+89BBiv71SPiBCGwqOH9pM2P8bv+bl+6Q7VJ6OQjPZrTDXiDBYV1R+
PP4oc9SLp5LjEuTQ4tH3WDkEqa1lVHdsvUzoedVMtooiNVHn1GeeIgMyd68bFWZ5
/fDROCuZ60pI1xMhmcE6ljIstmXbkHTq4ioHld8kb9Ftutb6Eulr3emHgHAJLMxa
MO7IIh4KIjSYQM9KKsUEZgxp2jjkAgcCmfby+qsY9/1nU7Q2yrgE/EuRPr5OZc90
RXhdcP9r85cAYQatiSgl6XN0YsCf1aafx5YfqcYRngPk2g2brtMGSoWBRRudwGK4
cR7ns8hxB45S5lAfJAgXwCNLmrI2tSerexKPdtH1JsRl/ZdcIkHEjiPBJygrYhHX
IWSUHPd1zXmWND79UlE7ArgovdY6IhKP+RG7pIE/EJ2gFe8Cd/QCWidbFALXoJ/y
0c+CzrS27oj4jLQJuoV07XQpM9fsQhKc5GUmDFv6lE/nQkaCw2kO4YmZo95mBNJ0
VO1AGBXgLdu+jiY0OG9IaWWvmMVSfFek3aMI0/pjQHYZloHnrWSD3swfhJ1ppToq
ANrAWdFARLonSmMu5NEtLbNn4UOx1Z/QfcEoc/MNKtQYIrZ3+2ueXJthpM7RFewI
CrL8rw8imp5MYdN3yqEJe167+FKV+CACWw1vjd9aVtGVZryATukZTx7tnSmpI5iz
5w0gBwTyxsUTzUCUt2vUQsOZ2XagFvBmNEL8EOpAWxscPY3qr+wnUiNn+SqUsw+y
Hv7IRpWMi799hvtoxmKhh0GFKU2tx/D9yZ4WtgiefkV+2idNvP7oG41F+Ci9fOMo
5RWg4modlKB8qFXLU1h7dDWciEtczvgoKveyKiV1RXvEOMOPEJxFT2PQm6sxxqAH
MIaAdFE0pIboq8h8Vz8M584yo2ZAmnD/G8sSURdChF+HUBv2fXf6QeOQLhBongFX
F3wJ/eOsuCzNYBacnslb1iK9vkOs8mDXpDICkbU/gDXOgcFauHjQxW3T/jeVHKBN
iFdtt5fIb0ijEx/KWuU15da42FtYtNDN+DvV6MVWHtMwlbQf4woKiv5H3wbxNk0f
zA3C49yoensnq5iNqU50K2M8RQIb2OK8rDFQx4ghINhXL8U60Iw5wlPl+TmYwKQ1
IBrbkFRu+qAj1fV0mcempDZ7qmmtHVqByazZ6utNYclWsCiM+7WTMtbSw1YF2rXe
g1m9zsjKLrJQt19UshSESxSnyO4gPgMhi8lJSgn+A/sUJ45W9oemPl4cq0S5P5Q1
UOxCzuh0K4BDg996IKYvTawztmBQcEVk7tGFeiJC/+MRTlZB5KoDuBYwjRfM36Mq
GEFvr+LGk9uNXz4coS8b9KLqnSsojBkNyholFqtruCPG2tnNJIMleQQGWlYMnC8Z
Us/GjzEfLayFIX7Kh9iXjt348QNkiR8AHo+IJt8DtU3CcGRNDWpzV5p7TUtDYol5
mpLEAOyiOql4URJUFqESiu8QfjjHfHHmuXWhcX+IdlV0GukeIlpu+bcyV4recj77
DrHHm3oH28+uMLkVwf5F7GpkM+wXzbc/pO4X8uFfKrU+yrdFvXoMQuWiyH3ZyBbH
9vluut//G4aeJ9OZlFFgjTZpyKqi5Rk4bRp/6I/UbI5KoNx2wblL4tKmwB4vfTpV
rgHy1BdaxdgyGSVSt2bPrzS+IgPsXxcssfvrVQtHpvPMcsGWej8imo8oBtEehBPF
4IEblrefnoa4h/5zYWmo62MymVr55rPjFMo80WXoBaZrIBvZGz1cVClD6IbBIJFE
F2PjpAqgpK7K18bxjKG6+gkiw6wn7n4AsyVngl6yHvDZ6keYPGF1X5jFeJFYPr4b
9G0l9nAA5q6dgSH1mT746SJrof2HnxXpc2JYkNLF0CGg9GlLDgbQgeEFGaavNMu3
nH9QsrB+PB18vzZnqby5Mcl0xwYel6F7W6DVl3Rx95Aab4C4u5CSQsFSjIRALNbF
fNQjOVtQ0p5/9csji9BjNdXpKO+fgoKI9pTVDu+smx6664aJmksN3N1Uvuzu8Rrw
Za/FM0CDxCpfCbJi90dclZ/MDcDv2+kcQC61BWMrl+paLH3Pr++lcZTWc4N9Q1eD
8WPUcestpK2+br0ZW7QPeCAJEKT8GEFD3ProBk25F5MF75MdrjPlImL2V4wMkeea
BbwXuYHnMca3uX3yLIBxX6FKLwN4aY6YQzusbUamGhD4z/2Ety6IPA6xp1H6UjHS
un5nwr2FOLAn2dIgXVAhJtJnXWvJa77UyD+FS5gTWczY+ttF/dasn+RIudE8vE+9
COucOgWGwg9xck8e9AA3A2Npg4tqhITCq+gy/8hOsUCllKbEcoRlkvKlQvhKAh5k
0H1uYqY3JMtzy4CjUYYRk5IQD8DuCTTl/Lq3wW07q8dXqIVG97EWwoOdZmALd51F
zVHqvMZqWzHugscGdgo2fmLd6bv2Gdzn80eR4oITbr+sfkSNiIcAAfZP0rlxxZnz
fcRwHv1zLGb+F7FfJbbODvIvpSfL6vwd2Ul6TkwWZl6fthS7C3x4hHNWvpZopJZ9
lGyD4yZDvNxMEVFzj7h4czwR8kcOviQvy4V5IxFDCT+HL1kAGKdntZ7as6r+7WOx
P+8GJ5T5K0nGL8HfuXObCSvR/0JG2QDzUaRao85h87sigoYIVIU3dYI1VRngrlQe
wuLkIMAHweD6/ofA/NYGVGTOxQGNV/Z0IFZ63nrQ94jue2KoTLbKEDlXxNV3YFt+
BIXuekEii78cZLLD0BaIbQc4VRgGBnVX38/Tcf5xqDhDjJEwOQ/JDwtmhbIXLEmP
n02mLPt/WGPiTzbQNJ+GeZ8Gr428R1ROO3Xo/x9kFzQqKvm8apEvOlBCxvVCS7pa
94zz6idTJpvGydaIWxpGR/67X7/sqqxTJQyYooBZE+GK7fsFbsJ8zmTZa3jKv0Qw
HVoxMRcrSewH7VWkRpVVuTENcrXKRMc30/YUjBkQKGihgbEs0UDHjwqPxVc2VcH6
3o7WdLDTF2P0/YBm8dvTtXMXpeX68lGP14ICd9jqgdgzhbNP0tSdGhaj7IIeW6h/
x8Y2GNUDH5qqLkx+TpnES4cJAGctjoLHsHZwjNAYZqpme6oUhdobYazKtLDu4D61
rYBa7eo9Fm1Gqg7uPOlefI+uzsgDl3j9Kkkki068A6MATQKHPZgTDrmwaeOKULQW
RDtD2KL+UPnlVdVLgiwZsZlkKGvUpT9VvvRLJ1yU0XZNSXhNORweVcY8XnC/3cFn
DTzbHTVR2FJ5nDj0T7+Tdj9FpZhqAtxJLgdhS8M297BaV7c7k3CIDmolJqx1zH6j
WNswpjTgWk58GIL69Iy5JFUIKCSr8xXVIEdx6C4k1RhX4WekEyzcaty7EoEGUj0E
PMuHsvtWzxVfmJ8Udx/Seu18Qm6EMNLixlWSXxMdmOAwhdOFXD6ZV4cMc1Xbsedf
Dzbx3fvBbVlHj+ZcszlW2cnuG+l0q7RDtC6rQ2xnzp26Mm0HcVRcdctm103ME5UK
hi3RNnK90E8X0kefzlwBYrW1o3a5AOhu+6rdKtUFVvo3+kGbNXSnJ4IFbswhxq3H
jVs5eZz40A4g5gbOCsHGpNAx1nsqxsUysf18Fo0E1Vog0+3/PJpaOP6dQj3O20ax
5HeNxSL4HfND+JqVvotp2nirmzXufGXirLzOjKYbU2uayTEP7jKnJqAf2D0pgIFI
BTuJEQhq1gEfqwaMHHWKUhw05aIgZWATf2V1XyjKL3o+OfXs2uffAUCBsLm0mDXB
IhEeFsR0BgLEgGCllaIYz8fUBNyGsLDtYNPsur16T+lsLhqFa7yqvKlpjGYTOgLb
iEmHmMIvSLjLoe5QLMXC/J7JAMAMMJrRSl788Cyx7pH+c4mU4zT4AK5cGLPX23nr
fVEE0hAiqkU5NXAmL87JZdOGp+OlDLLOTHsEbkNWY+rjpYtrldTtBjZlisKd1TNb
zc+Q5ETqmzL0hHHfkwrst4H60+znI1R87B/tZRMlg+gZwzHuHHQvIRirMjNj+YTD
k6etwLjyQchmI4dIiI+da4+18im7OIpRAPEPLCmF0qlAjODfKan4xbK2xorjogIH
FaU2GtrgGoQpLeik++zdtpJAu2LtCDVu8OpGig71hMigCL+yDEhxDnfNoTBQ34dq
4JQCwkUwadaQ2RLW2c5dMyOmCvpT7VvGDQu8/0rU4zIyp8nacma1kddtotoSa6WS
yMOuEXtmsnHezQ7N+x1udETshaJFArAR73g+/qBV/CaKSDpdKczsW07S3F2kRXQ/
stKQqMZdYveJdorQgzFes9nxwEXjKaSPdYcb6/vO3t2QuRttcStqZBNu7RW8WkoY
Gd87JZx2NYIzxnv6eYp0oPRDqlqJHIQddyvUBlNptqnjnhoK/olsVcm3ME69xohK
1mT5g+F04Ukj7zg1KyXXAxm3AIxxlHIq4NA0PfyIutHz7B7noxmTS/PG1E/KQIhX
WZRfMLvqpl4w7xptv6fbNGVIyGQCmr/501s98dg3G1OZDuzva505aM8TqjfigfEI
hsqy7fOWyrX4qn6qYdG8WMJy6KkGTRcIvqGav15BCOS9GV98hWoDo6jK9PKcFoi4
UJnWX4STHy+cpYnVH3JO6RwtjLT4Uh1i97zlbj6y6jGny70WnH7uaoJ1nxbHb70X
TEBbrWtIGChXa3fZPVExo3DT/Acq3XmF72Lw6PIA169JUv/IneGYLeLLah6+SlOv
7sjkN7yZCoqpwpX3JjACJS4FncDzS5OIvalRD+Yvi+p80266F8mXgWBrSY965qUa
JxdwO4lw+5quPu9nOCHIvyozu+u00s+FrkUeyFehRhK60G+NAB04tvmqhTxK8YMA
IPNHOtAGJS7YyoetwRGfIA2V79HjZ5QmYr/cQs4fh5P1u1lULU2dCBow6dssEUDT
0GKZ2OyNt3qO3sfX9AGV4epAMTNHpbcirqCeHITXeCLN1FfxpyG5lW0SuG3GnGtv
GJIxwiMGnUCTqraBasFtjfBQMN3uQRPU24W5MSh6f1d+5JgNiyLDnfPVYEIi0ACb
Oj+Tf6SDNIrDidhTUQynbbMjb7CiucM11Y+A8sYpZU43S49D4cQd2FvfRdH8/BAO
AXySKgT+xZ+oYyWGqWKWeK1WGUwssL11sIbUwdzuBBl0JQz2v9l9U7XRSV0g8u6B
mLS5KMrB55C9E86zKUV2Z6Oi7Pm/xza8WgMtmAnh54UXRC8Csa4Tfip/Ixhd1BUM
sDXIekhVHGQ/0o32WGOBtpWWg/4/vScRrWhH8AedYlK2uzCasYgDavrYDSUHXRwD
2I+tx9+vTQG0fPf6ESdC9f+5sqhTcYOptv/HjObUe23DtT4KNTgKEzfRF7GFj8Qw
sdJwfFDkN08k8plwTgLESIabi9PHDVg1/C3JFmJv4RktRjHztwkryJiWuoLz4Vm6
WfAgdbU5xBn5GVMkFsCtkoWRwuuLh1qNNg2YbycmimTiUMMyG2vX50Rwq5XhN/WL
oGgLC47yWFDS8qv2jY+G4WuIKhhjIYnPJumcEi//kxNnq0Cfz3/ZujwaRE/JJe6r
h3m4wkbcxtPuoYijbcIfHuFgE5ecXyQTjk/yvcG8V5G6a2VZ4HQzZEOD9ZnRJqw0
LlzFqyQWQuArv4+432qo0Segtl5WdIxr1C393KcDC5FncrdbXgivXpOtkYS+cOKk
Z2jW0jpv6WGkYSFGyy+wZKkUyYIC5+edcH4hC+HL5ZIvcrnRJaoHIhg3x4S3QRyd
7VwFkOSH4NlzHTdJ2cl8Lj0jnvZm1E+jd8fcxtngD++fP5YPJAHFf+3l5Drn54b0
tSFkNVoyY3ul5q8XFnIay28iqGQlSSeqVgHh7HgZQjvM6r8TzOkYbqJ8PfROGtj6
qpxj3DSEASNhffghmrioPWGRCFoyyFqjGtyeCyYr1Cr4US264vZF3NshINAAq4e8
mUTOOWMeALF32g8fELoqQ2CI7q/g6LQcqQZDcXSPl+HS3CTPBCiO4DMGf/AX8noP
pNoVG0ZM1nCsMG6KU24ETpha7WiXHlakHhX8fy7SUmhcNrqA37VIXdNoST+fLcwh
VTniH83Vu56llKKzp7/hX/d8v92Az3xD79CtcR5bZhbCOhPVDXjxmZWqNM9gEqw3
fAAbVYFRqWaUGzZh7YFarwTY7j1Wf+GB4DhwZ28WFWxkMNxpnweifGoSyi08iSJ7
QFN1xcdJiwTKk6WIJuGKxbfKs1jJ5cqCa1jjFqSg7PBX9zH03yov6cZzyrz65YDS
h2tA5W5nZfG+QTdbtYPoxde925LDQXhoiIY8MBWFWMwxcP9nJIkLJjJFeqMAJB0t
futxPMERoiaiRfI7IkVke6ohgdrni/i2l6ytwv0njLEak3xuEK+xn/d0wnek+N24
kXJBEXKOObQKRyUnYTeFl/tJcnsEB07PJgtXywvcsJr6k6iGQrWtDNPaSWCTtnf1
C52/G1RSnHe6l/e9lp1w1sLpPL8cdMxrKU1Ik454gfGqpOuv7bIg+5lWL9fcdazP
UWbVFjDqGbSYeUPWTPXgviNTIoK9Y0heuXule0+wLnKFM8wl3poN6F7RaSZn6IHD
0yXO1u8967UC7zB/uNOrwFddljadrLs2e7WV7r1fmvmtS+lUkGpHryOpVQKkd61u
GlDjrRVTL7U7+pHZlcrady9NyTSk++eoOlLUWsGb6fgyLj6hXkZE4WAcCdk1bjhP
raYHR4zUNgJm0RKAuDUwcak3koSEaqRiLzDZUGAvIOT+ubEX3oEPxvd3qsvzJxNG
kxERF/aXWrsaKTluEYmziOpyK9fXk7es35mMHf0glwsXaAIsdY9lIAAnkW1PiJzg
iZC5n8+9TzJe9+O7TKQd8vfqLOwmX8Fn9neLBzHzK/ictJdfp8UusZrGa3wBksO2
iHaQPGJxihlJ/I75QYSW95U2FUxRD+wOw5Wt1Z5mhIiMGSW3ffN4q/p//dbzbTYR
FkWiX0PUejYvFb3gYJwu7n+wvk27IZxPm3Z/4xmUlhO84Q4v6XS+HBs5AJjeYJvd
fqumw/hdF2Vg1nLpC/gqERoWRXD/b/RxGaTgR0io9fDTsE3ZR0K7KB6mnTU62G01
UbFldqfpcxsIVQmq1iRAMjXTrpC2nu5Mxd+Sn1j5cbq3LYJD3hm25+/uACQCjKYN
Br13zlnTaAyKqHl2IAkLapqn+d3f8+7X7SgQEuXGaCS+Y3QnGpOcUTQAlM4kXC8q
Dg9sA+DFm2x95UI1DEJTJyz3R0BLn/ZTs4DCyw6UbHG//kCZQMG/E0nvLxuCYd04
YRB5+O+j/Q83cPDct9phso46RSfs45q1SB6MpJWLDYswfN2/cBiHSuuSk9VMMQ7e
6AT+0+MgJ/YMhRfntGqjApHgeJPbsbgOztXThO8lea3REvV9B6EizaxF87XUH74/
Cd9kUgZQC5ILhnRUUP8z1u5yy1OrUaXgvhKgSLAPC+Y55HV2q6UtYd8quwccIi7N
WaPTGXP6vB6839/3poF72873qm2lOR8RBThc7TQ5dJtECwL38m4Kv1bo8GOxcGzo
by4BOhkT10JVhn5bNjuiVxDtR1V5bdRAKqs2eStevdde3ojAeuzgfACjj4YVtB0z
gPU2piPAWRDM4ArAWcNYMi5xnOMBd3LG+fjdEmHZHhg3NZw8/dnNW9OZFRl00hFL
PY++/CVXEeDjRU5cfRCBeVSuJY8s+BRmr5IlpK/163SezkSkJ+Fxjyx9Ashcjuv2
QEiW9jl+9+5ss0RL9q0AhLgjVqxILsB4QGCVMRbn2km2w0wNhfEZP8yb2cVldUQ5
SEFDyUte8O/i3ZUnZt78NcMY6XXBz66QT0yDQA5RRE02DXLjKIh/54Iels4RnnDy
BV4++jncnKkfqCReF3yP8hK50cS/IYNrekTcESETNu6P/1X+bs6/Suh7zgQH3/69
XnzeciVTPe650GI1Cx/t+dW6ZQeS2CJWEUlUn24rKMOM/FrWvJ1Uu8yTh4g2/bUc
tKow9g2ancbUzamNV5Zx34tA4M3I9V/YoO4s/j6VI09tg/nPIpyUy7LyoJJ8IApy
Yk+3x24hZ0Xpj7TbCexo9JeWvOXKQ3mvBOurVrcAj34/Lb8Ew/TrZmGE8IMmWM9q
NxR91dGkjjsFVH3I3nIki3opE0w0+g/95mED/pSxOphLDsRtj2VI46jQIroy9ql8
IsPokIym/Ut7Klt9jNGfjlQxGhzCaSOu/k9W+9TApxDBdDk+SwyX17FHmiVqLqIz
WcRSZ9waGxW687b8Y1ooaZhoprGHtnNmoZwYaW+Pe4QN+nCPT047sdVbYV4XM1N7
shFiJKC8tZ2hPU4Un/6ka6ieF0qWG++/Okamh74Eap804Zievar8BmYNuxrFAsOb
XjywLF8geFa2VSAU91S69uIlXhM+oES8ZQOFvmEWCoM6PifyPuULqwr/v4IVUD/L
LckbWrRViakCjX5XVdtHDLne1lMP9ivejQ/QGdykDYb0icO2WEWPHME1vKB2fbg1
qTVj7HBOUpvPfOvBxION+gBhtAVPsccBSNQioGySicgDTtay0qexerWh9/oN+MOd
BNS7cEJCBf4n2dxplKpBFvO2Zc7DfVZMnceWhQL5/7nEHIC0if/sk+bR45BURc/k
GeW2dw9a5ic+d10vMks2wqFBzcRzMbiyV3dZtOLAE+iZYZ1DIHIQZ6KFL8bKUtmv
HFoKdD0VUtfj9F2PELIFGKQoLPrsWuIohTmBSor7yFC68UfjeRLL0L/2OZ5pq+H7
2qfIUv8GEGnwnxH1wUGJjxIaSWLPrmsk1I5LBIDEUwIUjP2P2TIJG6C6YAHGETuy
otM9tu2dB9zJEcaJYo4AK5SDTNsE1HvLf/7wcmfapYz6s2pIE5VLDBB0zc7LlZD9
MUyTGS+fh4FAS9PynCZWt6DXvCBu2AZPWWzR/mT77OlXpC1JVoVpl6gqh0mik/wQ
mIVjckgIly0FtQqWCcvnBsJz33cdUwn7XYzjfHGxeWmypPTQc7x+/HseVl0/MV5j
Z0HDDJpgqBX7gjfU3xl/vXYHurujPyMywp7vcpAKTxX19kH2ABeat2k9yUp9wfSU
qGbzVC6IPtXc5CnvchTTmnvJZbPaav/bnT2gneQiwPWEapFi7PZwWPKaOW2RzaZE
dG8p9Zrxezbm14L0ERv4OSXBD8YVd1/F/KiUKsEa2RUstSZsn3NW1fIdRUnw0JUs
RAy1RoOLhldGXFr/wlsSO5WdywPD2uLAeyfib/cU8u7XlsJ6rmE38EMd6Ukt8MRk
cMUuSqTuNTSiSPZy591srsEnmBlfM9Namak9252Exsya1S1EhNWOF5zvkL8c/Pkk
PZhOJ419tevYDff/Rtb1H4ZGRvQPgGW+YiEPILI9+VWhMESxM7FNu+3BUUVi9Hbo
w3BDNir334f3N2tujK/5PSKM5nB2MBbYeKx3WK4q6V4zEkxTd1QjyXNcJNf2V1uL
aYVUqZlA5A7QIdefLJ1nPJqYuvDpS/6NTWXJ19AU1RDNIN8idqGU4XBt8YraepHA
iM+ixdzr7cn+4mv0iwqEWthjvDzqv8zpveRTJM3I7Ubl8EzTT4cfpRu5eNllGl+I
PbAd5DSyE9ZkJ8Jrt8b13+AdYdc2Q9VewMCGWzcXhDS/cPRdV/a14oeq5OVLQNZ+
PL+1A5hsljCJ/yKdtL6/96Xw9L0EH5COFuaTT8ajg2zRzlfZ4o0acblaSf7VeWOL
WpyifanBX9tenm4y1/nF+3jOyo5CZyCnEAOZmmzNj4HQ3yG3hAjSyTKlhTw1SVRY
spHaEdq3XSCCP9DRPKCCTLaOguWUxhAs/qMfTg2Z2P2u4nn9+S6kcgd14Sj6TY9e
+Bf8I8k6ejRSYxE0Uyu73UGyInjE6u1Z/8KO9xkvydlf3tgDGtrkkhLvIEr2p2Vb
ovJgAFspTQxIXWUjSGGnel0d8jhLPB/y6joIh8LWJkEO3aRYeS17fGXuTwuDd7cT
y/Orul21jIrUMlFWrFHl/Ju7uE5Rqu1NU5PUXPTTevWfVceQsSZF7mWYYkZcfYLL
G9kQBVxlmSd3W6ZaoKv0mZ54RNeibM7QhPGv7uQorj/6vF67MEYHw/3ftagWlg/r
3RTuTaDEYcPfihfU8W8SCfj/hLTJD9cV51q01x/ejBbG9PL3V54A94XXYFZe7hSW
nrwlhGPMLh7Cerq1PTrmaQC/jkEqPZeMtoVAFsxZl1UM21ezqLJKJMU5Noj8KGg7
h5BIqBNMiLvsT27c25NOdu5KrsC4/L8rmE8peGiEEY+g9fYnqb0OGENeMPTOo1s5
jupnAev6lcVq7xCzMYI45fnTYVhtJ1RiZ5juYALVYOeWVJzl63tK7xKCgq74ksCJ
R5+ZhM/tEqG2IMJqY4AN0ylOizxMijmj4QFH/v8+xNeMIGVecSrGfY+FfU+bEcQ6
wvf5FgPv6Z8Fnp60yGgGlZjc14u/QRjj8zaYLvqw9WSM9P1lWlJ9/VsHmCudZH6J
AAL77kVBBW+m64w+wuUTvvsyGHhmuf2I4ZwuoG4CfG7rkbMxgJ5bJlDdTWcDMWv2
AwyCdsNmnLdSl7inpcSGipRjLIgymqNHDj2t5DhtKtsKyBYk1TJ5esg5I3HPsm9y
q3bALNm1OlQ0cPS1glm2ZbRAhwND1M/oVqf238TKhMiQHl56TGkwbo/2kGYdEcNF
QccB9IICJz3/nVBuUah9i4qUNae4qYjapy1ozddoqrozm5aOoz5jrht2MoSLy7Z4
NHfjsH/94NzdXoiR3EU4RTvwcNIuPX9gaicvvxTRKj+FxXSM7RhujZUPJ0wWHkd2
Jhmp/AcZZMZQCm7qfzWsIChuxi8K7mAYUVe4RiRl2W7U3/105O94JS1CPprcI3lR
xzGswkn7uS/WRBs5ILrqZXpWpnq4schU0oCv1HEJMyRGqyCmP4IIp5SyOZzXoYmL
SD/cZ//xqywOQVQliYrKv6I0gPLCneE0xgDCX7wOA6vGvJwG2/lAqWIRRccgE01N
X4G+wZ7bL1TGAd4zl9QIlyY8gF2mn1/1FZKOokNPS68xDHyHsPM4j1HZN1HAr3Nn
PQGNUgeFFNqazS7wyhItOQZxtsOMJzw1BPncmkw0CxMRjsRJTXB8I78ZhMDFqJcf
Ey4R4vOsyS8PgZ2KKa8HIRaDX7sRfEyidY8qOQ1RQsW/5eocY8ZHQ26GB+awaCOE
YQXoofRaIjpD82983JAazupy7yjbzw7K6IvApURzyVXhlyVIK0+xrpzFH7dNg1Lz
RU8V1MgHyHtfqipan86mWDx9nsTVE2okLha1fNWBIvyOjF80qpSTBPCztkeGXknC
sxXMRxKtUDpBjVNCrlBBfrC9MhktisGpOSFSJ+M6LGYm+1NWzzSeo3bDDBxYmsQP
yspH+m9cB5ILuRC0ZwNERlZ/nid9u3dcG4qn68EDgTWrujJVhmmbCgEZqg6aZA2w
duRw/Tgk4+zAzOrBXypEWrXDdZuS3tDn1rCZWAcpMwPyTfklq93m5Wp+cW2/HoLR
SL6pwA6tvRlsNSh8A/MR/8+1OJ3O58ij/HYkKh5zvTRKSMNHmUPxCfr0g5UROKFa
11X9CnhE4sfPRCLNRcMiDavzjGVK4ozIS3Uw/eSQNGtXW95zKhfAI6Xc3JNfAsCA
iWK6fIMAVphfm5b4Uk+z+ipK2VjninihE1Q6CM8YEflX9txbNsx5KFEnq25hXnHG
xcnc0n4setydaXDDqkfiQZdLo1pm61Ux1WAKTyvDMdvoXmChIVxOQwHbKd4qkyI5
omNxJCSTLnOuGMiPoSnJViuOBuoMbICZVGJxJD2yhkPPdB+VEWgmhLIiOhU0JBtA
ZipEngs3zF57O46YSmA8CwfVD3EGhBcl2frtAo4CCJyPr7tOCSK959EHa1OWd4CT
bOqBBpNUdTvYWliNNMzzGM1o6FnjEW2tbxT8Rn+6ck675tAIORLUuoLfxoYwAUsa
M9nlm9ovIFkDrLoLNt2upnIznAFOIzN+CKZPuLS8UmxoEi0CWbLyLXnzNXN5x3hO
ReNNe+e1R6Z1prvEaS8Iphug+7aJwvZmoStK5PSdeOxvuQ3SHyJrIOlG5n3kuvxE
NiUGGT7fzqLCOUgZlctOeSEWchgkDoM8QYD4VFh3YfzFVf13VQy2L4PMr5ALumV2
4zinnN7396GVpnU7y09NrF+65JjjIfiUMnAiif2ik0tfUIie819xmM0tFNubvM8i
XktrWfQwfVV5sexluH4Osem9bdxTiw6TSh0/S7J2f6aDoU3Efgii5ti/ApqA7tFC
Sys8I4+I8b69ktOAOTyF2voYYc0ZPkH3AeOm+G3Sjaa5V57TphnNNqg0NNTKqkd6
VbZ2HpU4oNLG/5Ypb5A5UmmGT9xw9AWFQMGC7aLRwhNfjiyFVVWxczOMXr6w5GTp
lxA70ii2MLZoy+o87kbsUmLtWcvCGU3Yugq7YckgELtNVi4cewBV5+BJAwjEdGlI
xLBT1i8OU+GDGCeEpl/sRbzIMgsS4B3bfStfezwwyr/scbHFkfhxbWih+Lg8zedy
uU2eeKhFfERefab+3JWwZVlrAKgNod5xxRAMJtKAjHEOhhY0l5/aUU3V8toDcTxh
fGpiCQTh0Uk9nvV4FnzzAKKMaK/BIzJaiAi+4P8W7/79BWxZUgSlLnnaI0RN0W41
jzcehAsR/4iZpntGAXX2paHEi2/OKbB0J2+epYVrZx3jAXBOkpR6e+ZL1xqHbPLs
BDokdqV76H6Iy8lRwlJWfVzfl2DDeaD128hCprQG5nUam3NnvaY8oQYdQsOVrcPj
aO1fo84cjL8TL8JdgizYOiNbSwK0/1e0RweILfbe/sFEGfWf0nCOmxFcb1qXcOzH
qhPM/0sgELiAWvgVKCXQzpvi9abltnqAuu9pUYUUG1x3Qk1Zxt9U+let4Dolc9M7
2Y+Snmzc4T5TrVNaCRwua69U2OiBc8zEgFudbFIaxscpCBCTWSNFRBHZXWsua99b
5Zwy10m+iXnoJ2+6BHxZOLZEd48pfuKNRGtaFCT+KJX2T1l3govI9/F/eOJv+N4F
peESmNpfIYbRCc1gJYWB9/hU/10sZ2vzX8SOnopdPbnvxG6FIsA/1RWuDXH2lrRz
y2jC2p7WehbJem9v4S+UnzkGplXwARzPZhAMkVnJvEKFmaCDZI87iOIiowFG6zWb
kZAgquDicIKIHacmeN4wWzHLyqDwCgu9pqQOWpTkeCVcnPMHeJPLjW0dWouB7KmO
hf76+Fof/8MWJp/75xG/qv8FlNLHxj8hfJVM9vNQqm305WsbOO0JD3JUlgYuB3Hj
wjgzuciKamV6SPZrD/E/nAnjzzqX9YDDIlICsBYg1XWbORP7F9642a77eC1iwcn5
2/nrtbWgKtfS6mRHwZSnIa0e7VXbMnHWFqgRGwwJCHGb+HfHU0Tw3/zbaCCUjcsq
HhpyFd6mLWTDjH5MzHZqGroS6j5nGTbOURWs77WPne907voLR0bD13WXIAtF7ANG
GZ0Ep5k3vBtUf2QwgrjXvp0xCPqfLTNZMNxx6dAoxowiELQCsLN6lrzNWni85VUq
gOWkCH/3gW/Rbn1pNSRvLCXn1lls84I+m84PGe5D6+fJQlwTafx3cpoGz6+M8eP1
pi83+B2UKWg8RSZC5SAHWzLQA0a8ZO1/DrjGgsKM3ZPfYNJ9h6bjMJ2P6YIo8Jw/
lk7cZnXggPmJAiBP1QZB8kka0lsL+PuCTCj3XYT4F5fXa1UEzSklUQbhj3DzPCSB
nRUoO1asba1awHbKBJHKoQEuXTOUo2yRildrWS4lPonz+eJZviZV396eNezPGWjP
Gy0l34K1mTil4Etntby/GdcnfahZtsFKrUbu727cgzk5lbukO+n2oyNWcZjGVV2Q
vrGNk8rLDrEsobmMnsmMC9iuGRaeZZa1fo0N4bntzkkxNjmN8oyqKd3jrknXjXdE
CMnKlXm/6iCv97vITlu5Ss1sQzEq6CSb3Nu7zxUSE/ilp0feVa5iAh80Ojz3eMky
JWQw475MnjEKrXfVHRlTq84ZJCsEwOvNLnIce8UGKagOfcqbdAFd9WC6+S8au5PZ
4Wi0yVwaPEX4kPvv5q1KdJAE603i1aylX8e0A1Lorccz92oMCOUb7vzEcE7fqpg9
JNJc9MZO2kPCvJ4aUEzmOFuzQunkbtn8SknqGiCfrjWAz/b4z8oZg0y4baOImUP0
2de7e5DREoF1z01D2V6qM/kNQ99v/B5/P2qOU0MOq5DwM3S2MywWyHiEQey3VpU+
ejfTifXW3RAhDpXYypMxlY9+fjJOTwW5A1u+8v3VqmCVZTy/c6wkD6FVV7GZOzEG
OS8CWVBHwJf8/nHx+qmY1pdk2yiAkBTPZLFOK9Tglj9H0JuL3AFjJXs36Y5nb06A
+9aP3Qi9v94tUtcj8mCdh5jAiKbEwFlueKKWVV0Nq/zL67XJcrCYQfPYNHLbP3zd
lZBN4CYg2te1+qIEAPG1T2ix+7OSkkP0PdbukpbX3w866QXoOtaLS19dyLxJo+Co
7WoWu4QCj/20b6qO1sBqzai5HRWxGdyhgJ1+6jw4v+CrId0VPWVGN63QTj6GBnyC
2skQSmUoAn6AZmPo7SnCCd8HmXvDjQUd61QeZ7Isd1Se/pvcLg+qJohOJWl3q+n2
LqQRX+7CoQMKIlH6MqQrJUHZSjRD5qDwF06V8z0vtllIyGM1s6IUwQrHzVXtPg8S
rH5P3QJfDXHOJ0uWWHypIuj3mWnQDKu74N7KEz+6EOa4YqJn7R+uEoJK9joMSJhU
rFRzGecr5RIf7qEdI5P+M7DeUJy+H+mvFT58GTJhCwqjnAEF9ImIlCaOWYulbrfD
DepttDXCFbVNzHu5iuoUodcmWHgyMRgnK/00HJz++3Ix2l2cg6Mm4vFt6kAXdOqq
T77CRpKibfkLRfGxeFR+5b0B9DoIS4TgL5RukAh8SOtGcTPUEi5nEtN2A7qHZ2WB
i4VgrVpKSOK3XaCz3xXEbD5ijQOI+INUs6JtB7brVWppbh5j8lPsSqAa8RigUKGE
bxothvIDIKuY5tSgKNf6aIImOWxzNAJ0RMd2zC+B3SOrBfEJrSxbgzrs8So5oA62
aJoCyxj+ymAbXLJwh/FyEg4+iwMnjyR1ZtUxVkbHMtOG5hS0xw7p0KGgG4So/rT4
e7KKyGA1PhTtSq2RmfiyxBjuuqffEcNsRjWdLUxilqlBBmhm9ycGA2Gdlz5YzDun
6PPrkJNSOlp3KjEZsuEG5FztxGUqW2Lni7e+e/UQ8Ow+hKYuvE+WlV+vLmkHHYDX
ors+MhDZZBvm87HTouFAxb82s+UkDw8AqO1WDn7xrOJM8kPdOgYXkE7w7YvR0+/f
TxI+/d6gxA8zw0K+Jvs+EaOKtznSLvLWhp2pcrIBtQUF3gq8mPOYYUqHL2e7lp1V
VrpIl++Y+OrG+Ai30bXbpo6RAUK4UqpFboZdqog0vaMkK9D/xjm8mZra7u/AbRuE
o8/Db/rA9iMloXDBAUD08u1pnY4b7I6jSOxoHZZ4Z0gfSGe8P8Y+ZjmOj4kmSgiz
AYbsFlc9zNervvKWHZEYQh4bB71koJb9yNLJ33Ex25kjU7JG6OLkjwzQIeDS476H
pCPhEI/5DhTFg337R3LIRzPyksz4zHVnho4J4QUjxF+ucNEhMt69ewqGwWGw/kgB
fusxSsZSiEZ4/u6S10uM8uDC11fDEgvV2V9rdyV9UdvdC5Slh5xBFGuSlSiC6C7H
XKPmqyaIoT0aRc9ca4uWRMS0hpmyZ54D2US/45H0YFqL2I+xgMgv8Q16vlOV47ko
bCRigsIjZdsjG604uLVr/RnXiKrBleI0AtHldOtsT/FBRLOQIrwAm1G8VwfkkQUh
OOrfIG49A/U4CJfMfBQILW8JWTg6ZBM/rnkHFlA5Plg0NqKiNJKpJ03126LH5RyY
XjZOf24aM6gytSHKls0mOfckXc1wMNAgIITkRq9Z4YV5J88ydW8xU7UdNHncsvEq
FDxGmI2KYWhmuOJFI6UsOlsoJ0F3/5kXDpI/vYBFp8wod6Vh970mBGdEQn8P9rr5
O7bd4reB/yAqrxSfYjQ6XuBiRviHyUt6ufzq2jAa37MbmDty/OhH7zssGFMHHrSL
LrN0ziaIxLu9aiPExgNFB4FWCBNXq7VxmmJbpTKYdL8mDANH6ciaPYoRumhtv8jy
PFdg2YnD4S9JPfowwH0rubYvTIfCD5dqBGyMyw93zaO0Buey3NjMdvMyHwebDjo0
K/QzFVmxk0+lWCQvXIJ5YOPIUiYQn5wd6NMVVn+hrz29wjuOP1lljD9NVNmwQ18/
2zL7j+uEd/qP82Lgg1rrFAzNrly0X28jIzDcomA7xJOdDVwHbzAiejyI/6WjsiYv
pcjWDmRPcbrC5MHuNHWZRMFfywzqI42C8lP8WGiofsrkZ9qHPPPbr2i2TEXDypTG
A0NuatDQJRYTnfaS48m+j4jRxXKrR1WA3oi9UmEWWzf8Em9OB1KUf9kLCdsfa5ZZ
sN92ZNiTzrI9aASuop4A8rlCTzT+aoLq8Q1KKs3Y1NxmgCjBpRPo9sZX7cue5S4A
U8ISUPcnPFnG4KmaSrlJdlLA4hlVqz7St475W5MZuBp8r9I7Od8H8UpktkKLpcv/
uHHQuZIhixIwwZcmf4bNoKPVnc3P//ggxY94CUbFDMBbgUAQry4vko/pa1zTpqYH
EXR7HYVU+mXZxIOaUjwJ2KNZGtDN5onkHOU0AUDRS4sZARvFI4bDmSAbnEoUFLh0
QBuOdkukkreJ2WJ6Xm2u+fdBCNW3lkBZdiYlBWLYnsNtciSw0AeqRnOF4Q2knsN4
zNGHCA62XiBs6xe6Arf4ZYx3fSegUZkB4jHLTK2x/bqAG2rM3UlLhEQMB2GWNeh7
psdS3likYIIQ1W5/wq499nrvFg/NqvwGbJid9FAAZJmsSJ9rWSrOpnA4ILKlCO1x
OCVCMR4z9neLg8iVpCNjOTSmQcbJ7LEULeNpGXHBNO/iN2cttj6QNzvegRPTS/2D
afDXp8VGxoj0L+ZzFMqNci49Nz4s+cx53/togXqN5cHpx5pU7hhl/rvgrbwTbXq3
HOQDa5xg7AtyI/G+Uw6Q9SeaQ4uDvnDnSCA6c8xGrCkqL7Vm5SR5y5q3IWYFjVAs
0E8xPuIDgsk7cjzpgbbDPbg82iUBsr4yJFsJTe9TTsJpcPzA4BssXPGdj2b5tY3T
hyq2cBYuWpQTM8jxBsqf4aPkrVeMdPYQm4hIkyqGCZpDt9dtPfrRf7+yNkqMradu
hfL8TUlk8/lDJ0LLr1sSC0sd1T4Spj6A2rzHhPkrT82Bb1HcQusTtQObEa2adWty
IKR+WCM2bUwRkZKY8IgpbPn63SxIUWF2YbZFY9EaaiPzfXzosMO41IADuE3i3kOA
26ZtXJQvwCtQ/yz0XQAOSx2i7wx3/LHGQxDvvvFkriFCtl0OjA9GuP+Te49Naw7X
cR2fbs3HHR2FAqsXRnrOwp12B//+rsRmufUrT3z4BdGYq3seBw1wjGBWTFy5tnEk
WRDOxAXScWOhBGIXbzRGweQBgjXB1FXmOCPrTQgD5u4QnVG6Jgk+jRmoHeuUw5VC
6aqz8fHNmMJQHpkZLRiOPjQtIQZV/XleOHFH/eUOshOhESybncchMAY2DTHcltSx
lEJ1NcMdBdWaX4Q3/W9NyNkCRo7iEqsCA4XRLyWhRRvPJSRM2DLthg4fylyMghdV
A0aM9cb0a7XFncXCFDW5olxHEToEKvmm/04X/qtDMom0RUk9a4ElFGq4ZK23jv3G
LMDfcwxl7zxrFY74bo6M7p0tiuWmV88bXdnwb5tR/mxkvG3evnyvi34+MsRz/akU
vbHQfEs+/ZA2Zok/Xo0whIHN8xLR7CsTmh2e9USlfbeE4VdMKUok95ykCPNmwgvz
0eWF61dqmWalxBpb9r7Ty3dwJFMUdExE378NL0YxG73PaoTRqCA/tkJvynO02n5p
YFYqumRwBbts4Ug71OPOItF8NFoPhnEKovkRrOddw9kv5a6yBK+olFGZVFTP1beF
Fsx6rFNNDnoBp9z2MhW1gi5Xqyc1R1CmXTGkBKl2gBnhMaP4HOYMcFxe/CF0dnuj
U+M2omIoURw0gwY47auf6LdY6YWXVFsMgB2X5VJtiliLZCPTG47JOh4shaiI6x1F
u1yFGVTqBzHB9TG8n2SDN6xgnaW9qMO11t3AQ2Y5TFdU+87mxHW6qFBKnd3OcnED
WVeyJiK0zKpta5VIGhs2sRBJbrkqKOApylYKZddL6wE/rB6v3iqBCxlFmEUz8S/O
sjQfym4ZDncubeYC6Jcyc22RQlkz4A+9w92+AEDY98i8DMPqTKJC2tMGkInRWK4x
E2htOLOHkyw6Rd+/xdZp9RlFsT3VMWOgoU6kGmE5kBDdG5ukxJp7b1wIMMz13wy0
kGwWBtMVeLLe7wgcywQOhLNjLo4HP80yC2TuH3yfND2y1zESz/gLe5ZSr94Z0GHA
jZv/MarBjHaQXGlLYsECc+BXeFBYuHBqyElsPpWhcqB8K/Mi8nzO1ZTQxjiFIoBk
a3DWyfgDyisqyv/R8+17Ridj9Tvt71JafDHZy6tkDcpOOUs00CGD44RqdR1j1naH
qA0W55517znOI6HylBx0cCYzbrLx9QPhEPppi17MnTFqV0liN1jsU6Kh5PUdVpml
oeVHpMu7AyojblfLxYTGseuXLWxTtsLiCRMZgE6JhbZ7RT2KTa+6MyqWDD0q+g20
YGFIqqF9cIbxtHhVsb6Z3rUm+PiTlr/1NvvPaYaY+GXrm9ne6CN2Vq4liF3a0m3W
PIHnsi3V0FPND4qU8ZQrIb1EDyafiUGF1CONxPxD9xGXsrNvYwAIJsBUToG9rxD9
vMBQSk2j69fXOmaTvz/HF/if38fbDWcitxTiyLB+fGoKU69TeYZOO62eYTZirCQS
oasWb0smW64DDZPYMyamTxvWTJxFNOsCsDGVklk2/1wA5OK79eJwF7iqFUzcGygL
Dhlh60mdCWnWsPoMwWy9kmtYyajACLJ6Bl1Jb1TpBQ+D1i4Y8YDayC5IezBerwA6
F/QmmWP0MD4teo8GV5AONbIEv+8WuDeoxCkRPkNRP+ATHQV0tOs9YiGJaADX8toa
TVBHJ94UKkDCV0k3noNFDdbI0akH7BRl4WdaqxCXRHvGFepwzr4sMpPWdhVlkums
C+4LC7hVS6vJyHeJwUb4c/PgMioCsNKc2vRherVAiRw/OUR69aSMNTMUfhE+Qtcx
8qJiirPXElIYe2yU67SuRS29vTyhy8Dc5xeOUGwh8WOKJBz6Rfz6JQ7+zV+bO3Le
6+Z+Nm+U9lZ1S0vobmBPGBXo/JQkJDkWARYgggXC05EqD6WePKJz9ozntMhW33SE
KpMla1meBncgfqMVfX/geBhxe3A4CWZ1Owsm/G2HGree5X0d4/xR5Am+BvkDjD+K
BA9cNbG/TQv6fMf0RPam8qMYkFgUEYJ3nW4CkHd2wicUhBCPQo+s5x4/tlh84SGR
mIogzyepatZP56jQRURkly/dOE9vDw+h9Y1NvUOIY/+m2aN/vMWoCd4USdNc2JDL
uzFTA/ceGdYAcERAXPrNxyBubcpCfkJNQ6Sn5wiXOek0KoaAh4ntByaJpC0xk8Io
Xh5EjPvtH7mIWqeQcq3aI5BXx9r1Pzbc3LcOnpUiOi/R9iNuTetRKubKH3OyobWU
vkVvZAaDUIvjIA39OSzwpRMTmRdnyPLupM6T4GbXWR8FnVUQNDlSNrMUpRkHbl/3
/o/rogOxn9OdYUWj8g7yjwk9GXSRxpekXgsblPrcOo+V7aArTMnwdkjgsgeYxJa/
QWRLXfK3qjwykgjhuP3emtA5H3ouPN5cqcsbPMl3krL8OpRNC6xiSSKGlqORHGLs
isnKR940Bov8iNpFlSqQI0IWDVGMSaLWLrM4M31sLqbSHUci7/6hKDsr6zjahTKX
rsB9B3cxNb6GnyPmios0XXDrlDAXJsvOESQ8yGW1dCNpt1bezuSouLrjy5J57QLB
RYs+kR6adUrOAk19UhWaJeEPGU08s2owH+bQtvZJEm2bQwgKPm1rTqkfKwlu5Reo
FbkYUdxWEC1DeUILiN2f8fvZAcoCxC0k3DTAEaiy2lcTposCV9YFK9CAQ5chR1Aw
xSjgy8GMXzVdPsN0+LaDlRvwLgEE+VnhTCixpwrzCUCyWC/QuAouIJFmYjZ6o95u
i7HCmi2V99Sw6cHqdj0vw3jtUYW352P5uYPUXj1+Hn0wOaG9tChPaOcNrJNxymd+
KqxvB5wGxZfCw70x3lI0PNaIy0HkPmxfe9yys0Vx8JpuPoZqRb+6/SPDx7+x4zZ7
iiEwnSjTsGe+CEfWKXy3/JTPSXY0zNUTAO4gVKZV2uEoCtmxndLSAIBzwVVAgFxW
A0lIOPMcaXeiw0ReEnaIggmUeIJqsNbo/RlJpv+3CHpWkcpe5GKIU3vs9hPXeQe8
o0EAbUOAWREKfgIOBwP9ZHuqIkKXyIAmdLNLG1pjYl+UN+jRqHqMRlK3J2OwF8Ny
O8wV6WOAgN44brtBx74A1MK2Hsdhe7B2ASri5vsdnNxGrJ5SrgQncN4R6Pjl46yM
PPZ2U62iIot8Dvp+5iW1MHaveRBtVOUakIdXsVqyxeFZ+XTMLH4GC22e9gVOWaPv
EJ3goXWhn22fmmdazGoULmX2nYXtDkOnFv0LnMLwXYRa5GU8j56bv0WWw3xhvC68
6c1dQJ3gerb5ST9jR0GgOmh9D9QtFutPavqwDr/HmMP4raYmCjM34xf/QLs9g9Ua
oHzzE1Y7ND3nB9gzuUdsWa/Bnx3VFhC24S5jnXPVHC0n0S7TEyeWOw8Af8Yg1Jd7
4KdRSFQ0SrmasplqGzGsdPhCmvuC6tTuOYQu0Jo2MEsvgx74/KKxRHMQXKgQmGyl
3UPm1IUggX8Ngyuf5YvFsQ7CjOfTI/Fom6afguHYyXAwLSIPZaxAkkDaPivF7LjX
arc1JuUk9KCm4BkF8LuIykeaO0XwEbshFpF+MqdHV1ukn0l+r7vydY6LDwAAkzDt
MXdIlNPYZa6wg6rTt5eedZ5pPo0guAQp1sjO0pELsrQuwB3aoOk2KmnH0CutbWjO
uDkNuLWFNkbbBL1RHdl10Iu3DCOijb/SEw2BZuYQl8ZOnKC94mJlbfI/fJfST9M/
pyznAOLYpvLLFEEl3Ny6vu5IjCLiIP/P4OVL0xKvYH8wNvQOQlW1SN2eRUsHpuF/
bw39+4/ACIVlFXdCWTdsnd7FkOOXYx9+qZ3fmKlcpg8/kbJkeBdAWjSVzWdeXzwi
30s7y+2AnZRS1DjWdzEDCKGUMtovVcTOcPP5gVTdekhWn59/03vuTHJPVxWd987b
Bl6PwPbIGlG2fl6th9/ATHDHg3DJAYt4Hth0ZAN6PZ4NYK0RpVfsrxutLuFKFc5b
byRiJq98qPNWo22TbE67ucNlly3YQuPn+biofugJJNqsB32Eh/6bEFJz4wp92Fxd
bsdVfNEpjvmzLZvR3C83Z8k/ijvShOu1Yyskimy0QUd1mMGXUS19AsUA6pGHru5L
7kN7oXAm4Pu/LTZiYLZLXcmdOIkMTzExczdV+R1H/f/Sz1RIPPgzHEI3Pbvi+jO8
g+EGBgtIUBLhUEWECPBd6onCZu81F32w9IaEwB3rAYY+rK7J13EhzqRhRzh11A8y
Ilx2erzQhJkY/fx5MUYemRIFzRAd1j0EjivwZDhhSpihaW1VljDBZpNWmumH+6ZE
aW5Lui9o1jwsFq807Qc3Ge9ePA6EJIT56jwHlSdmoj8SN4G5KmY+ZIsi4+Vh/f/F
l8UDstkwjvcUz4FdWd7tQe/3UycDkZkK5GAvPCXGnh7DAWvovsIGpKpHAcLcE/zO
2l/g0R2jl7kpF4wocuLOnF/Hdt8o6uDJKKdpxB3E+6SSDkMNhCF2lK48gpCK+Xzi
SXo62zxBSql+iE/rZ3Eqh3Ichi5LdQ0bZeXMKEtZqETuu1pYzW37Ukq8VmiEsOHl
MhpBUDp0U2CJOvzYnha2scKex4JgH5ngijyb8OO+6JORm9AN4tFa5QgbCwowvrPF
LXc0QuAOVkT3O2IMbZGIJbvlc+KCm4yn4Inyq9yjD6ruGiCa4B+bIbCgoF375Ru3
QyZlvaEI/FaBqlaCkI+weilGWpoHijUizI+5Q4PbEMoCOCZO4koVnuLlUsmgT/0T
7L7zwIOK1jN6MDKBCJYZSIa89n3NIbgerAltVl7zeIr2MTTYGKaGSk6dGRjh6xe9
Y/STE9wkdcQuFGd+kvyZt53pWDAFIoZ/ukZYUL/MeBpbPlQoA8QVtWfzqlskDKGB
AlZ7aB4wABGKkGUuKQW7F/mVYss58PMhlp/zOSTYoMCM59MRBeqFC9Oqzej77K7U
BcUaXOku3LrcxGlxnP1PKgoq7IhzRYW588TtpxwRdrAxB8t36FWXbHOjDurluoCH
S3lBO/trw6c97Tyf6iRQbA1O27xyIfFMYnCBnBMrI1Ak/2DnZKKvtDSkQcTvyz2R
9OlOz0q7RSZjVaECRIJKbe5WwvZ+8AjrBYWedX1Pk1klKDmb2Hu7PoYqSj6K9Hof
+tIT03KYinC1Xtlf659G2+80ucuGinFY8JF24nlTB257cDRltCZ7lHDe2w4qFcUL
cguNvTjm+/5tqKwNSVNmB4Vbdh1iaGA/4haeSeJb+8ocWTj6h0lrFAiC1gendSQG
8yQqMoPTG2MSNFs4hRm91euNlq9YUjrVAiTo96JnWBT88nQ12i6mBiAy19LRllUm
75ZSZliJWmoaVVd0Lp71UNfoirNubN4JbbA/sOSBs/sTBpji72lXA0YQm/OQAcmk
9BmEE5m4wFGm9B4ZAQhWiU6DhAGCScKHnU9ODnnw/AJNXgZh5RVl6LqerVINCWnp
i00KXsQwexTkJjc+HuoEU9FvuHgMXgGIC8xXZMozbGLmHDNQ1J30p+L8Eh+gavDI
BXeSDcalHJJiRysoH+YEz7Z+jMA5KUP7HaxENROgQKXpqBsSCUteHxlEhI0LxjTj
p+X2ZMyGxrXnP5gYKjTiYpirqGmFx/tV9+3o40GXguK04wk8h9IBiDkyHeXJ0hAA
oGWWaVOCuazyaco2MeFLU4wUQY862LzTpiktrBxI9pt4pTkSKjGLRT2ge0JqInPc
E1Q0RBnCGcVKDYf7jGiGp9cuOLrDmfxjAVt43r+th800W9Okex6L/vcexNRqfRiy
eJfNmZaxQl+Mn9xaf4YC4e08ltvtnp340V1ussh9w9yPd8Rid2TmIrg5b6fZeJQQ
Yb7MDBGCSrEdZjd2aVfFBwvzRJxg1n4zV/fyLcIIixmVluxh14lOl2lK12UlAlHb
4z3t62XXCeg2JAItXAP0gC30WjFMZZgYgBImhNqDSXjZlLeRYyELb5ge8Jj07PQ2
XqNl0JF3xcnf5oI52R2475GX0Lapa3jzuToC0KNWIffFTnpR8FNMRrjMYWILk2oC
jYetQY4aYDpuO62kU0KzDc1Y67pHN2+uwwKPYBtfcQ8CqAYn3T15yi4e40w2KbCL
lb//koOA/QDj5mjLhZxVA78gS1BVTwu1hzksUVPbj/2iybJFakPmdN9LliO1/GvH
DYfKLvPlChkGxcFKucekBAScjzN5psg6J5aYEkTIe0jY8JXpQEpTSFLNSFU8Hz1G
QO5zLhp8IDuA8HTKfsx6oO38GOXMDOYGwZvVN1HCd44b9z1W3/01l6r/bFC8UgZB
Rd8K6YRxPXVx8GVNO/YmMPRiLJZ4gGJZ/385tOWm3QwFDLO2esnoY0p8zFNLnlUe
0rVyKpXmv6oo9rfAmKLfVSmpz0EB7sETeS5lxhxkRNP/hAEf6+AdmIE1uHVrVozC
XZK7319ILNmyIhtTqOhb4QIPzjK/xsfG89I6dg4/x2mEJKA41QuLyVBBLKGw5jTq
0WU05eV/V0nbDRKZn2itWjWW5SP3OAWDCQx8Pl6P8gTgbDjeBOUD+e7Pltscmjz6
bPXe3dvGrxNA6k+8CpfID+YjOOArVZOvqtMO6ht+7bxeuDQNVqD+CP4FkMynDXzO
jXQMXrObthMwZr+emuwcEhsbirQmYe5ZQg5yj84gx53PvM1c/4k2oaWAmy6Soa5G
XU33/OWCjkUzc2j6e8qDc/T2NL/6zAsao9dUPlkhTj2bw683cD0FC9mVNtIZmXW0
5J/44sEvCbJe4/Ty82LT0n3JM1ieOVPPiD22hAV24PSSD7krmzPchIlP+PSh0x9e
CI3IwJINzbeqqoyROyHx/YV4RMCMfIE8ZZEkW3c77z73ZQqlbwllFkO7RFfpl2/u
xujV9zYAdILk/u5wFrNiqNuNFg5MjKQaTKeLaAJssnqK3KwuskrwpQIi7IbdDuJB
cAMcIui+q7YXd7ErO+xi8XTZ65o3RfBqf+PB6sRsM3ZqUf34mfFjleiidgvcma4V
jGD9wXSKv4EizWVIeRbQvOKxokqBUdUOZ8paK8HCoJR4J2Nb/9o3L0tSruT6o59i
j03eUW6xsaiTJh9UKmoplJcd4T44GbchukvXGC44h4qPRoUj6c7BXxC55uYPOaiV
AGrbKJC1LMOft0qF6b4yT77UBRUV8msnFCKNoo4HJSdFaA9y7aUTMxR65BhAN6zS
biv60yYvxxFIpcUsFSmnkldQJkNYMGAnZWRAWrLdy0XWEcV+vI6XAQIl7GjZzus9
K8lM0ZwJLqK7ZZclXMtN9WdAWUDNs9I7wSkJQY9W9tEHo+kCNt6Au3Sf+r1nZfdg
/oCvPREKddQ5EQleCXrZb3enptjhnLAGyksMFVROrtDQy0YW0P4k81/x8caF9BUg
iCXsXiX6a1mO821QuvpMdjzxgaXBtLcMauMh2zJ55ANRl41qcY9K5QcFszCBze2g
qinjEVbkABPCezUVxpoYVOuHPRZ6a5SrqPyQ+MxBawM0yDGW/IEbFklaG0Lpgt9y
Im7A35DnsnGKsNChDJ+66oAH7jrZPen1+gnvNBlk+3IqaGwzgtSdgPYpz8LEA7wD
iAgfwuVVwuixFDdaPoruamUBZt8h1XhJ9cNvEhi6v4K6fxLQQoNZclpyD3AR5y+6
1kSlsh6g6/X5NdP4WEGPy43w9pS8LDW9pkL8EA9q/9TEz/WXKlKF2rO6oaa+tviY
z9ACMIWHAI3IqGUwORXS8W+94ex6QNdLx4uB38y91yKaaZYGAIHtBah0jgzRdUBD
gVUkccHSXLeL+mrDZbVtRpwO9BPi9RS0HW7cGE8IeKJdu8bFGPSwdpRCrqcn10ay
nIVFCrd/X1UeIRDi7qnGV35q2u5bqpeoN7WROIcY37it/vFYXAVQwMR6+XESDL4L
KL+/KE/mFPNcFKqY1l4t2ue9heVSd4foZ+EDWBJ68Cfo0FH4sQH+5HFiF1P0KLff
krbFTdbHsJ8Gaa8+ot2dOz6Caky2F5/mdt6hB6wVaB+wAfsFXkjpbRAxdZ4q43Qo
Ke2YloCP7q6eqChGEMdSyyb7HwEKJWUV07dT8qTyrRsQb1HH4vipcFaSQxtpFQZf
8KmQR4ACa0sHFMMlDplbb8bb5QnZ1i1mKrGPvwI4bM8fAFRNwlGoMDlsRRkAu3R/
KbEGnKyKAlONnv8yA9opw74vJasQ7MDqtYcdsRVjqRrJ4gL/10x0YuAhH+Azc/HE
2OhsbH16cTxd+QF3kqhGal3Vic+yFuB9vR++410EEHqRkznOAWNQp4jZlJetbL62
5oh7hHB18nqiu0JDuX+Gpi09bnZASDpWh3V1uIKZhUVWaMjkcERkP7XFnL8thD6a
jED6p/ZJeBVhLpaElW1QNYSd9Hg+3fYxsmojTH5oAwfbKccSTmsE+ASrZjF+Lfr0
RNGD/YsNIyY7IwpIOl+W2MLywLZa0TNf+LV6sEA8JsqQNWXd6/Dvo5dnjY9XHDlL
Y+koPx/V1Os04XX7hCzn8tKSZK2LKNFm+N7XzYgesnqUj2wpE5D2G/qCoiJnoNdL
dVtfV8sdn/JXmu7wOCAWBG2Y9NyeuS93YtMMXLvIT95FmT93hn9uNmUEQ4Ew9MDl
KwvfjmFrHziBxUd7/WeYixVd35ZTmWZfG4ciquGnnB2BXSkxwyka571d91ohZJbA
c1JWnSmPhQWHnvjDdNTHnLlOnuzE3J6OO8y5KB7+gITYYEx5ED6YaTI1aQBx+tWh
4LltexcQ6C4tURigVyELKOn7qDjo/B1o3oLUYWMdQoWZajsOUp7ZDtej/w6Ms6E0
dvwb5L9fqP6bU24IRDGAlL6ZnYNCPM7IAT869YQZmN1LtHsJ2JqsdmEUvctS4G0k
fectrr64PMG2nNHN1NsT2SCVk3tbiMnoB5zL/1KzEJT0yvS9b8blSJlNA7XEHe/S
clpXlbjLGaS7q/5xbfyDbPXLr4x28L6FMGCBPyQYHACL1e9fJP0JOaDU0AgJFUFl
pgqIydZ+rp1MnRvXgQTzcxcWb5sBaq1E8IQJwm+tkPOy/vP93VEw0egpb6bGE3PY
gG3BDlXz7BeFRD+KDdzBN4Ro/7u892hIf29yIIhwM/cm30hzCu01wInP6a4rvvn0
Vr8d+vw1SwurqPEkyiCylvo2dbU8bNS5OWCmzZ/ZhvZZQXO3wK8fJy4R8LBviaOP
+1TpPsNEXCA/Kl5sx7yZSp/Z0vk/SpVuhMTZG4pxGl4dh8XdbgMB2jHhIK/bNvVu
kQLSNOV39JXLuRo97d6La9OmqRDNgMtiSxd9VM2K+t04rElVSGyWTwzridXPawz9
6AbRPjzZ7w43+hy1SQYMFyPoMxCata+KeqPbSWV98d4Su+UkdwQBRN4W7KJOwhtX
MyezSuDaubum1hmc/rorRzK+arabjT9Ep1ZnhMhr9suFxydEz4Aq1qGp57q05YJ3
tvjZG98xwldxUNqbxlnFm1zgFwnU6bJH7kTbrOF0gBtcFnm1eQ6F4l463fE0ry5X
RWNbOFX87vL+FwD8+0DTX1meNoB+hbTZjHlDse8VzOnhV/UdiVZBKKqhzoRhaY/s
W0R4P0M2QdmucLyTMdrVFw+MyxvrfLWfxOCSs+WS1TMiX9wiJ8GsAOhZhpZnmheU
a5c0h2KlcUzA/SDosH8cYytwKiZd8k5Sc3MIiD/JZPtv3boqzBGigkvB8DllutCG
SZ0tQjazoAaK5IKpklTQt04+YoJOyIa1MoqLnc3T7Q5Ca3zX8ZayoIBt3Ef8yqHi
6I8AZZLbOwkMhUnKtKhSmHNxpO5A6AlAune/UEJalN/F1RUS+gLZU6JayYt/8wcw
HEpuiMffRflwrYdFw0KsaOJtcSzfTXaJC/TfDue2aqFYzA0XLHOvspIHSUxd2dvs
17DiOw8x4g3gwHEdUFj32gjeZ0xj31YiCX3GUPCboQypX3F597S1K+6Lzb5o3e47
x6Q9AjygWOqpA/5sGxGhXRvlG48lnkQ8+D9gFDoJ//QV3Sq9UMSkCI6cD/RJXXJn
HjGhoHBLEos9eAf/AgKHBjEDYvpGBkcEY9Svssj3LuUlBIDVVoVlU7KxlchFthRu
OPINCtsR0Eh87L/oc++w7QQlXa6rzynzMpOgbIL62hK8SkxTFEj1z2LqdctMFQ7X
Nqf5goGaJfAUar0EAsDekxV7VAqB7ChsOZ2W0q7JZEdAXRSDkmoapBY97b1zg6tw
eXKC94ycTi26syAQimLY1841GhDi1TBlSsu3DnNQQWO6ZJY59KbTu0eRBxI34L21
JoJsxgSM328CNTR5JR9XFEv+laobnZHR5FZ4DWYD3Z6Na8phHXATNdKoCkI2aITU
TBiDSibP7q9IK+e/3tXjBUd31nFILKPAGFoh4PiwezAfiF4pw9di12l+NdHpeG0v
FX/GR+P+8jyYk3IBqAwsvNy+44iER0IXqEWMdCO5+G0zu6tBjP2IJ5KyeOxh/hI8
pLTxdAh1J5B8w0RaoSCtfh2boi3wkdSqJ8bra5hlU/sbuT6fKVtZaqXA8MUBtkdR
RVjJ1ateCjP8mz89Bdsv3qPC5XRZhMP44KvzUcMoVW2VDZv6aSBuMhhayAryWUuN
+ZCjIfp7R6amDfJIFvOYTXv/aJzviJq55Drt01QGxb5Jx2CGT6Z54HzQ05k8hTP6
CgLz0DZf8X6310uehrsga09DmrDaHS4RVIJNC+pyUB7ScjWBTx1UKlw/4q3uCyxJ
yrGxyYHGbR2Ty3cPCXUbCzcEHe0/5s0ONsSEVqxV89tEk6d4tYbjJH14sHQsVarm
dJE7uWcFf1JTJ4KxNOwT7+gVTjJKyTIOnfDpr+O1JlxxnIf91xWs7kBRLSI0D/cV
iWE2uRDLoGqG7yjHL6GlG8RJqGoikwgPCnUfBtehzZ1UhvH+AaGuDk3muAH6pKvb
pjmS+SthFc45e0pA+pPz9iQ8bhxHR2JwpVV/sN2nk+9sx6bj+gFlRgoNgm0yGEOg
CY+z5H0p74dRzUBQVI/R6jpx8opavJo8msqvKBCfaclNyPVsLKPHL/X3JqOploTN
mOl8N6OA0Mk22I+0rBqHR21hGHLw59TETsT+1m5NmYylYl44dIC0ufTcXujuJf04
D6cbwq4oZ4QVTzVzVkULM0f4ODPWuE5GslIk1D+ih2KrZkfJupbzmTS4L60yo7Tf
es4kMsLRVI1Jb+CzwPEfqQf7Iqk+0sy5uYd0Jm70ZYd9Pi1IYakXm1T7m0DXkUEq
v1UiEJEbYGWw6hcezV3u3txvvS3ZK+5YMH9K7qZ+aBryWpLj2L1D3djLmXg7rMmf
cjm6jeBK0p0mVlysC5vhg5itiUUX0yq6tM7jcKyxcSNKQx9+bkYlH7iyAFn4bTIz
QbTj5PlVVXvfzo9a0To/KNgMRK7/02G/wt0phdIcwiCe0FVgJGqg20btUI+KDlbV
blJMN1PbrNpXCRwB3CO44sHHsghvtjwo4zSBpvB4gYalyRW+pWei7lEYsqddRPEx
FaSr90iRpOozaKCIQ3tk2lOker4l+LDU7ehNUwWhv/s32bIl2g3/w/bQrAbFc791
rtfXiZRP3c2f902gTSu/fIv+p49DxltPTKFXTrkFbToctWD2f34haWPowj/KKRYd
qujltfS9ysxmqQomyyn6K0Xsdebb+IZ4m3gVFc3/QIOXs9v67DfD9zSsbeKDrxDa
3PQKp8+CQrwy+XC99SnKCD9B4vf01QsIyZyi4crr4nAby4FH7QB2wNgd6qFuvsX/
ZDDw0SDDRa8BSkEmPy0ixvfX3P6lx/SvMuT0xgnAyL2hb2RonhQ4L9PFi+2IDHip
/0xpDdd8FLdcQKWgUVcz04037NB5OMImSMu62uwnRlchZH2Ux50tmoEDMADoeZcR
hTtCppsbZTZAk/tTWdczK4tyWaAWfZxXGCMhnTboLHNlGx2q7KZEX+Fg/ZUl7SJ2
8FMWdBxtI+9Ambc6mi7S+PkTEOrFAlgHrDc52xz82K2Vg1XLCaXjhURKb68I/Jpl
JF1aNDpnK/0x/EN+WQqAAdWkYfu/0SXr1wvcttSmWQaKt5ohzJ+tipny3X8Pkp1/
FQ0j+ThFu/h1yjPh7yVNuBCH+g3OKJbzME0ZSVYNtuqvCIrLlUMeEtWCA0UOaXMe
AT6egKgWZwY6Uv4ufr0K3uFiJY2VTx4NTGvInapUkQyZKsdw5QhfPJ7BiN+omhb1
9OkgyBM98FwIRkEOo7nzoAZg8FieARjeyNqjm7iBpw2sQ/d074exJN2L05M8luDx
PBMU+IY830J1S2k8ag9Wnmc54aaIzXDxaU6x0fX9jZGZ8oenXoSx35Z0+xOS5evU
uRA1Ok7YX8Afwv7aVh6itmKoJUxJ9Ee8dsnHjfZQ077HAGWKYHnDhgjWppvvvoMJ
yVydqfAShuYjlB6qlC3HA3fVIHBX4q//7AAjsv8tCSl4qbcNPz4K3bguACL2l9b3
nvpJqbAJBlP+yxS2Ypp/Bd2cdwQcOv806O1SVrbJoGpdYfigsYNjH9t5DBbEh5dU
7z08NGrpdmyYljEZ92vW1q1Hp7bW+ZPuRaVi3tdJTjft7Hth7kUucw6Vw5etxcSK
lcgURkgpvAKAQkbgfYaGCpMAR5nx3XMpmCseAe+86vph/F3adshyEE1lqEeEDyoO
eqEhrjVzuYOL2BH+RYmx1Qh+ZhJnHTxki6i9CAoeJOVVgReUBviUIGMAnv/vhcoZ
P7mU1hQSSDmCm/QwLwJBA9ni0UDOm/cwjJTeQDkmhNu4MsBNTk+hkARB1lvWKRWM
t2FF2cc8I1W7DxXmWCUujjG9tE6eLCXmVzvZulPG81fw6WOLNaKN6dzbfZP9dL2D
xHkjhREb8QcbeFqckjszE3/8R+4sjXBiNy2hMGjRM44C3dpLwXHo9gb78Vy8aBbR
+glgcjX6kSPSZXI3HfcMu8tI3t4HkoQVTUSSytPGlOGyfnCpB0lZsdxhsJbLDdBt
6Yf8hbMG2i9B3CdQMAFfL+mRz/NLANMBdi0PH2vKjzTZjrtWbmO7v2jPXTbOmYA+
9wviX92hP51oNqE9PVhjoXn1qEZmakDVnPZdI3dxH1O2SU7GW1zSI76Jmca+Z2Sw
p7pDuKkzkiukTrkTNQKE/rpsgf1VIHqaPcr/fy+GWHYgtxofdAcja7JRsndEsnAI
kNmi/IKDjDXp/dqF5n+n3nmD2B9l15bFZO38rL4yYIl7zAeeu7MyzsS6e2sb0js+
dI9IaMF2P4R9jv4YY5CifOk1SRHEZguD6vZzazScVkl+S0bwqnpQVUEbNiLGAGfD
AQLK7F5IUMYuRrWjZx2Xs3On7pcgJrcfwS5+kSDO9Q6tyXnxRfnSsXsyfp4xt0SS
cTb6K/WSD4VmiNXMhDn0VPEntVQWkBP7okHaR3HNzg/7w7Ff7Uj6HeJLs3batQ7V
YgA1ULPWp97CWUtuuZ9h4+5XVkSpVZfz359HRw9Nqyv9RPjYynyqPS+x1++tn7Pk
kke3tzP0ixz+fD5hhR3IwUAkmQpGZo2i0YNj/aDFWw46xoLvHSztzKTnrnq3CgCY
brAFRkF6cRtkSTJ2UHMpa90HxCTtwK6linS025ver+upGghynNckKV9Ax76LARC6
jnWsk9sZ+0KI6FxupRKa5/cLtX7zhxMZJ+2Y316itzhDwmqG/tbBeM35e0kT0tue
MYS1wtLZAQvU93AaOWDD9f/Z3aRe74r3/PjYD42jVdK4lRzcwKwEORry3FIQ8ek/
bUNCgPecKyy9S63majagREzFDiKTLHJvyagJX+xa5VFm1MzwVWgjXaZbgFZR5ZCP
t6R5FynuBTbteCjIOFinf+Gl8jr9iNGxHQJjR/oEdIihQdT61U0toVca70tZ5UH2
iMGYMxSLAsQYpQBfwYa/Lqt6JbvHp4T0Q6Zhhk9SBloGYnGf2mj3ohwd5cLNTgSa
fN/Ar4GrpkRe7P233e9ee9nRzEafsE8GxTLOdsfk30uj3QNxudujEsrzE1Qu0KuU
re4EN1fDZcE5C6bO7xMZgSx5s+7TRNIvjGNHbePtCj0X6hiGQoT8tM47FVf30T2Y
qPeznLYpNYuVrrqfANCZhH2l3oZ0bCXFokB1G+e6sT4OP/yGce7mpQcqWX61HWcz
XA5+h+TmI5/zovA1MEmt3+pUdIYbmVdWO/F+bIt4r9hN7uihu9jGui+CR/LSaAeL
0xkaqoZN0iZrMSeElwLB3K+rdnhSVuN1Qg0FirmQ+tU1b7AIPpRGWbBcfpEF2IpQ
O6/i25wejbf6QMj6SbtsgAqwbZumyc4QwsJcHI/fQLRPKDjkMnto/w9Vc1o9UxXU
fIM8w/xlRzESdNfRmN8mGEnXHfGsPdGoib11sJjfeIXQjq2buDqZWXjuhfa8VL2P
Wgd4l4hpOlowMH15buxp3HG4Vd9RJ7kVqXrAxeEUtgAinYrU+qLtATCESvDEgpVP
z4L/MZWiqrxlgeXUiHPyNdOv/ThRGiGWkM7AerOu9OdPtHN8/P16mAAUWQoEl04y
YPuDWEIoaw3BvOTRYk7awZMJrBv5lw0h6YDlZMmXKv3jhvDBsF88tHb3uM+DO+sf
x92HFCT3mP46hGobnjjDnwSdqSeSqZCS97inub1kAngig+NmEd8+pMNA2BWFyGKU
dHVDDs1vM10wEZI1eMMSZXvGCHl8fMdEjwXdZUaJLWFg0xi9YsNh6/lZRKiq2vaW
HpcmBqLaXxrntREEUJtP3e9NSySvFDLkSH8CZTOTXqo3UStoqy8q/ec7DPWagDz8
hxZwX/AwoGGYeBb872siQdxrkZuCFn9mr3A/jVWuFuwAX2Gpuawu7YiWiZgko8Ld
8fpsBT5mK1GbpDCR5XwO+2hmtQoMf0fZGQO7CXXTowS8jLRjX/qgxNmp9tkj0Cw7
n01bGhmj89fmvwOVhpnfi8wtkxvZJrPA6XWeEVhgegLoEakYCV4Y8xpZb2jjXkgb
f5PYNNbk38pZ70s+w9QvubUrI7Yc/13P+yhlvzCcEYTMqNjnlhcHefsZP2yoKMy/
/RCx1H6G1SmQIGDBRt0dyO6zVReK/8Y/oozIZXSNEvoDC0Q0w8hQBWpQYdgTs5Xs
rIm7uN6/eNYpsFb2v3A/dNQBQ2BCUBrhMdaOi7p20dMRdvrnfTkw9OvPaEQ5Hmyl
pBDRV133g2sQ1EDVMzr0TXOEALI4EcCMSCsVxW/N1+Ow2QaC+rSMRWw43x7GqagT
oFUUQD2eDneEbNStLY9HXbJR/ngF1x7f1aI9C7wrTWPbPMUOViDQhg727+U6/bbN
p8UX+nD7iPt2JpfiZmus2h+8+ANrejEIwPdvuoy5DGmNCyJ7Y7BjlD5dEpZE2s0a
POvbLL1hGXnTsc7GxavTYidOmghMZy8a9EBuDO9QeflMY9S4ZHsdIq8f3AR2lnF4
XdAMWCec8t8ZqzI8ZnAadd10omTcPzUTYhgbRhBNJS/iN8grNwZB+53Nv/5CzyFe
im0Ixpk0wQyGf9duxEuSvAG3gkbfq4PROLigE7PyS702PoIZqMI1qI/iWdw+nb/b
g3DgkC++hhsH7YT1v0fWCWwdSAb9a5Z0zhRJvD8b+7NI7mrZYkkHJCwGvjACi1y8
owovp6cHDxzZfZN8X/bxWcdBoeXBrE5D1h9rKOC/C44zJXGvAF34sv8NjHzcSG+7
wpX/4Jy0fctO+bOYwmnHb3mNb5uSHTjm5j3++ylRX6KQWNOqfCBZ7R5nUEyZxNUg
u+xguJ3451OkbcbjH45W8y5smGA/uEdHh/kp/lqSiiPLZaq2k2uGBEmO73wsi4hM
A6RTce2Ry6AroL3G9Y6qz6LjaY7QXvXAsi8LfewsD+p8F6Y6Hck7s+FL+SEmPtCH
QKAF2j+sN8Z+ie0GdQ4msv92fFbwoX+f4zljQ+KWFPX1sCadp55bUBT4rlCh9JXr
OK0V5Z65xQDNFqKtu+OhVRZYoyHoAsgNu5QAlOtahnzcvKwmzAKKZCeNkWmu3Ah/
RhrIWxYinu0DK4q5k9mxAVDkmP7/LB76GlgSr2YEe0xAADAZAF9FfMkRZ63gnHsH
umm3K2p3VhG5F3oul+oKEIAC3D89ereWo3n8uBqZrqAV9yDc8gupXbkkdzjlG76O
lpksT7XD6ICvqOjMXFdK85cQ7CuZTPRqjVLAWLq9/DdLgkV+WqTvwtmOBbOuwnrU
1JjfElOR6GYjamp1TzzTF3cQrxt/hKt3Kc0iHIu7pzeBzn+9H3o+19GDyfbrFyeu
zinEpUiJNHP8pERDXfI8J+0t2V3dc9IdOLg9s15VYIcvu3iJw9Uv3WbES9FpKIX9
pvtEiY+PelXilR4LF2jluvd8nQhlpkYrguc1ZyZsnLzESAJ4TzcvN1ldIDtrS4Fo
gv6KTYXOT0P/dyD4VDAQMjHepOdk1So8lfA/ci68wJ6/u2z4NkgwArxDq7Np5EOn
IKxvPagYWbIl4/xapBbCvNwhAkYYzNyBOtEJ65yBGfYC/X7GhiEqIdZcqxnd8xlY
ra08KTWEw0EGokC9Ow2US6pUPEkrykJHyPvsKdG4TwapcsG7yb4MnLt9MX8Av5uI
U8s9ZxhUakMWU+mcU5MtbNS3SwUb6O0W4UU2dnuWLoLgs8jk1QNvWFzrtacQU9Dv
kCutHx/V5n4Yf0hPWHXe9Bu9GnMo+qOEhnt69gMV6g2Ay9QsgPfuTiKhnCZ61vGs
lbjCOWWLBFmxOdYnR3p5TuZK4T+AoZ2ShELaNeJN92lNf+gLytVypqyfyOVH55iG
bJBsHWKFP39/JbuAk0xIp1/0EBhtzw5LUaH+vOLLbD8/Re2+E6+bArUNLw7CX/bA
Bm35+OLLAhF1q6KK3GxLMMNVPA/uDqyexyGk8NrllubBTDmsjQAIJVkRsy7DqM09
WXa4yRSsGOVaO0zcuJRKj/XZUGK3xTBGZ4Aex2c2Q9Ww/mo74DNsjfLXTLQRSRxh
5gUZet47xYLhGz2tIJLjhJdhx3mf9L0zX0fOgC5EjmyA5SyG0yMWCl+Lz6daGjBI
KrMqjewtJeElzVTsDl3IQWWiCRIOQg2cBAgmSzMoMEYzHlx94HLEEAA0Q/3uCXrj
W9Xss6b50BWFR2SNIE1AdPdFgvt2oY70Au0V/jGkI7tiigBNOL00BwY5wjozbApM
8MESeGayjHvZxlfxyJKwkByECWuae4zOg5Apmd7fl0HxkRvXCipZ7xfogY6CHLV3
QqsrsBo33h+hD0KlrR8J2LJ8P6Vs1ZieKY3KBsc1MmtCQY4ddFrob6YcaUjZt/wP
51M0XdtSrO7w0lNVhNOR9i6XbuSStXLh8Jay0tSisxX4TOdSKUbWcnrQSb8460ki
c0RB27OZSbS6gBo1CN9B+QgNtEXWycrXh712qJ7UnvlsXBMOC6Ke7cP2wdrRSJ45
6UJ4C/9VBB41NoKB2seoAX5daR5OOteTfIwyaR+teAVtXaNn3lCwmL180ewfqKlp
ymPrRoDm/Pd882mf8P2axJMwTtIpEOkDhu+DrtSIgjD5K7734yxLAZKc4imYQ/Zt
OBXpssGrEZCixKPTqGDVaKQBEG+4WArDnyhsTTCOHX2dGdqKUIFHgCK6c5JCYUgC
j7SPtSwrSuQbo+6PB316jvX7wA0h8CZKRcN99ByuZXMg1n7yhn2sXrDL5p5hu1LK
kgjHWhHzbeSm3XdJ3XWQpPtos0wWm0HxVUYyGnNDY1U+pAtb2iPTkeX6nw966DhE
G4RPQJCszBcmv8AU1tuckrtHtBICXeblw9CCW7EU+/irrGUuE/EwC50iMhC+QkSU
5udJEzuO+7fRHCtwY+CXHfg/lrwfarP1Ag5r/kKvqyTSFOLI43Bi6zzMvKxYYdrq
P6F6sJzkdfCgCFJBf8iRFZJ3Y6Ji2hNchpF8Id9aqLW3im5MDasGnjNQiQkzgNHg
kwieBxDNoZjGep+14ZMQ7GHimzB+YBbKOTZmz01DDHTTkR84866/Ge16kDl3Xkaj
gAZoDhHLkEYdyWjXUce0rooW+qUfbEF83Iz3Bqi+xl+IwCWjox11WR/HuMagIi//
vrjn8JUeJApEtBg0wERptgRS7iGGc6r3alDxAgA+d1ldLVSwC9VMGS83CNvwmBbI
+R7MRafkSNeQdUyMXT66NOIZ41FkyNLi9cm0BcSU9yvaHXMitC1AFJRAXHHxsaI4
4zNWreCT8CctZGRj0rSobAqreigWc8iv/U1q4K8RBe/2EN+DTpRX7HnTYT/GKDoW
FdTdaaMTaaR+5B/JeDOUu8Pgyo0knOJKz0HKJru7Mi+4+PvwSqLOJHKoEwo/SDoz
97aem09J49+E/wA7pEE177KKyxRbKSnKS9AF7FR1q0KYRg+fgozAbWvgrFM1Dfhx
RB3cgcwQXWwt5FVCtzXxu1IJXUDVQ/pi6VoNp/t0eoowNzAmFjpnpQJh5BCLaiGA
qIofXWaOJF/zmvKIN3hjs/LME1V1PZ9YqOLk2l7WRuwPEYsbD9nGDzmOiJyIcUn6
hNkRKO01Joi9fR7z6ErYxoMev0x1xuU2jYFH537JzMXTSvNd494jgknF/Q2J8wXr
N7F94QE6Z+zyEHNf/xs8ZeW2jxFAd543AKRfwAWaV479cpk0DOLnCLBOp1Q74ZKa
0Z9pzzTxa2f+Dbf8bMGvsR+T1S+r1kmPN14N/oJlPNR09iGDA0o4J/eW/R/1C6x+
zGCLjmHj5qozDDoZLgJ8F3V9oWfAPinpDSkneDNS3sldb+EiHw9Rtp4e+wQBqhMY
f+/y8n1cXrQJ6YY79DtormIP5PDCLCpYaF1DFzIYrAXFtD4XLPYGd7dV+UCbpxK+
dkGxl3EoHANfRVkJGjVJd1VusoW1NAaBDvSbKFUXGxkNywGmPd/iYmfanSBvXRv0
N7l/y0YObMsZSUOna2ddcnTFoamDaveukhNjsmM9kxlbMoQqU+DJxFsMq6DvDrD6
EBb3E2JdwyDNGu+KIV2bngyoLlaXF/1p9SKvMxNmgJiCYbH5S/A6WjSXBpc7BqjB
vCZyPtkoNVpC/3qP/9pE6TUxzK9Vch1cx5tJiCmjkcFHOSvxYb5cEUC7NopLDqxt
h2U4ZgW6gH8Qywyd/t2J778UKTh9hYfgPeGwIx6JQaSFYO1WCDPjHLkkDrvnXi1Y
c5ZAJ9/+i0jOPsDOw4RPCsYk5WUvdIBlVooGI5G8zK6eeQKhukmTJ5FUutFrjlux
k4mHeyLxCnWGmt+OLBzqzg3YdSSZcZaxa4+rYlyhK0vWoWcWb8sgHNoPDJ2D87sy
C6yTTzsAl2C1e8tLSDSu/97ofwP8/gZuqCpPWLG0s3h58NmMb2LtENs3HH83xeYj
AghQjg2vRdKiUdKPbbGCIVamd4DuD1bIOpSms7MDKhfE9+qizTv2lq8gcPT/HnOC
OUyoRuOq4OrunUVxnLfR9V9rbRf/llkzvL1DL/e9AEJQe+ZpgUEuZN2zgDeZDrF+
sXxGk4UV+p6eSayKmv7iZ6s5naGp8NxWPZaVJqJ+GmkezCjQ4RoOhWhEy1+yCgOE
AxKclXVJ4rGcHY7gyV213B08g+tnVM0wVmzSqJ9o4l8Q0HNB+rO2MQvdZUDYe7F3
vN1JtmzX21u4yIOUO8FoUPQYJMFc46cVie5MYf5in/eGuuZCSyzbVuc78lVW/Nb5
ZMQx1vRqAAV9lcgEd6QE08kp5UfiOjLyUwlf3nNWR3TREI32WuULlOjJb/MtW6ka
5qmy5x6iW0zef+tuX2A+A1f0kAzwZWf3zib7C+cYkhQMfVO/YiieEcdIPpTh+MMZ
U/flpZD7GJvvKzChcfjsl+2uN+y+vjp95L8Qqh5jkBXt6/zEcaK/DVAB8dUT1GbT
nfrf365de5Tbfw4TTl3cIrCNuiIwozD1DUFFvfEY/ykZ+TbakOgsfUnjW6kOvAtj
RtAu16i+CdJ3RoAXzcwLsWlnHlOYqzzU1g8lfdByHRzJROX9TCBB2HPr/LknrYlo
O57r1NCMW46n6osIvxFVFB0unkU6DcUTJqR+Cn6+IuyoVgGKnkg9B54HC7i4aRYj
EU4/PXbgS7GaNP134NAcIZv/HBmkJZPK1EJLjPj0RUmyy8kPVPGPWUx+mtfyM7XO
e3F3KxRrxuwMncachXHwUS54hzP5I2+/mxDAFVjlA1BWSeGvBrzOowkpBI/GymTG
YGma1OjFLTD0N7coEhRRV1RIXi7ObHYWcIUMTIX+P09hu2K50TLFm5kN4fQPPLh6
/+5PD6RAyqmQDfT3gBubb5dowEjHDboQc4agjtSoFxZ8NzpVXP4P4mA7Fpc5WXay
Y0RWCdtKKNdkcogskca7LQx1B/eU5TUu5yqqcSlFIWY9f0nt2EP50rkVHJs4Kztm
ZjesBJ6RLRZ2URpNAK29fc7capi91l/dOUpRVA8uQ05kCPQN8FAaIYi1/yNfVrrY
/eD72oPDTCfUWgxM5TkXpGM+L4mKGcVu/6+TN5Toda750P6gPaUm7gg8IO2kOOjR
+YbjOlnmd0TYzdO6EWIniAT2RcJEN5ULAdYQeBdNtoXZTScyMrSRah7Ms9yV7RFP
yN6Zc+mANPPMPESpEtT8JerYrWLUGLXKlXYpi1DR6qnFIsTcYPTA+ioWWWvL0Zhx
+x8h7xXgH/k+s5UGRLDVTB7LjxUZ7tLvyREltS7xBQ5QUjm3QQ47GugQueEU3eLL
bgX7K9Mg8dPGwsGmoyoZNr/RuH2sjXreH+ZJ7gBFL5CeVE+WWeN8bRDguexJHVlb
CLM3j35gmB6v7niiif0oDbOZ3O77JlPR/akdJSHukrxMGOJLihtykdnGysZ44anq
kpLI+WVaYUatQVu4wZzqrNOJiRWE3wQjpxS4acNs46DoV2/xXiu6Js2k7xOU+eRX
UwFP1dcnNZXv/hY/5MP3q36rUTo4NAY79JoEF7LjeAFd0dGOI/tIya/49Ds44Lnh
LlRcn6JD20Bnaq2QFoTq//d2jHX98ZN0xfLPVb99Di6MHYgu3ocMqpRU65wo/xCq
UG4u1Eqq+vo0qzqbfrC/cMe7GKVlqWX9dgIhNrhl4pJPHAzi9xPuVyOTvJjSDU81
sHI8wRmRhKkZc/X183XB+Cr98U2+8bXozDzvB/LtrZ+8zrxHv9px60XrjiTsiBIL
hnMchvGY1vkmEXhDQcJ6HtP2BqKdc8JpKcao4oVtOPKEk9lbOI4SrIoqVB+kRoGH
o2RbJeNyCfoUIYskQohQDKQCva/3roRnczF40uLMG1aQaPfBzhqnPkNJ+Q93vFCQ
bEfAftVhb2Y4l7ohn8R/EO8xLo+tdJ/ioOQkzJgIM6A0lKyru+rzAezaJBDfI+Bd
B0Tc5VWYxY8XPiYhCENoFSiKeK9yG2P1WLZlSDcblAVI6XRamhrDaJsNCjN4QKLz
ejKX+PCKnji2MKfQe3wBtXBGqcEYeh7reHxx18yJ8m3miewSwjUvG2tEmbU4+nZb
KsW/8o0WECly1YNY72oAaVM35i/y8UYntOk10ZUBCor1GyFHc/wb121oJKZrXBDU
vddQ6SoTSDvy0OpH3rGCA9dXuyB434m9JSWai3cxwPyhu5Nh3ZTKrpBkvrEpUqh4
yBERxG409dvq93dUsTUr5CVeMxVnV0cwnr8bJwedsgiV1e93rxJwXZoD+xu9IzQR
rmydr91tvc9BToa+wadl8YUuRatKbSm15WYQPwVwbJkKnphIATaGBBwRD/FISj/W
j1srW6R6vmLHjZ7dD0n8Q9wW3cos2qdkHv5GRQl4bs44UxDMDLAuseLmfeLjU4z4
QrmULu56Olt1m7k4OWNAAp4BsozewGMSIIEAk17NrwsANHdVdqUnS7LOz5Dg5+6w
5+0vg3khPx7qr1Sarn34Lsd+gJEsACmGLEuqnHyHKxKczf/RXl6SWq22U2DGNoCr
4MOymIDWu9MIvf65yBwwhvcGGixmcZ8tn4E3t17tv6O7djt7KdUPTwwbjffBKlRB
cS9MDONUiTwoqmyOkFl4f5UEvenybD9foSEqHT2Y1bObnulMxza7HCk37POtO/FY
y2rYSyVugmzEK/0AiPp+BaAjaNXGfgXvoJkuBHST9FsQ3eu7xM9wpGjbUa2GYN6J
hZP8gQNdJYqRanJOh6Gamgix2ZDPbOi4bPu6GZkLFr1+fhW1mWOYjtAUn8EenLPw
QIJg3wIlbsMWxCPgT0GROh66ilUnQfI7U2vZ6A3wGkkHmdM7BQJv5Y7NWTanNmOC
710evcKSmv1icIyBwvRdjlQyLrqcBebHb3Ogsu1omFtWFuNR5iujk3QoqrI2lDMG
6hXU2bh3RFh7o3KnVd8gPkakrIRjnrI9WRz2a5Xhm+H2tKvoPtCafxWilnSFTXOP
N8UY5ht3pJKuOqe9eJiPyjNL1KnEwRJzDi11eZpfu+/9N1JiKPyDcyGdst+oukpd
WIlSPnZemVvmbJ99lgj0EzxMQavpOQ9Dqq2nwhJMU3qQs4S41mKEySvG+cJ2nYqs
/vZBnn9iTd7pLxICHDZO+1CrRI6c7jzQTMJjZWWmCOIpMV8RwKs5hp18L45P3rAI
NcLfA6avFrITuSbsMc832pvX1jvvjsQxnHhH9RzGgsoCLWzmLGVWBai8YW7tJLmA
ejPkX0UIOQGaczoNWRQahpUSMzkCX24LSVafUecUgoPATZyFrOQzkubW51w6GaUq
u7+u9b/eHOKPdDd171CsroLZknp7nyQyFUPYCfrxGbzjv/RS1ebODdAVGpeKL8Ca
Yg5pfiYok6GVz2sF3Saex0EEq0vIyhdNEpEjAZgzI00R0IFYZw+wniz0nvWt5LkY
O+8EprSFQRK0mu93Oy/A5EFqNN7rTimQ6qy9qKQXce+nfFbqcHq7D3NU3kMQA/Js
zYjKIwZ6MWksKG30Dcxix4BhCESHuMiTKBQspPQ16N+jtUnqt8w5z8qNS5Nc9DQg
85suMDCtdSF/P1PjtVLutwPr5qug2wX6DEgVjFuLDAcP6oQL0xL/j5ZyLo8/bJfN
ixOftxZw9+JrmR2Mq364PRizMBjboq8CrRnrbPmqhdIp+0hGyRE0grFr++pj93lm
HX5rSyfzF6wTbAD01mzjAK2TRWOexVfJC77I/BBT4SJVvyQXw3hlkD9zzXQj1uxG
YgVn7AXWVxAla9RGQixDeA5Zfv81f+2/vmxIXI0oVmHIisxGCj39jsjwH6pOzsPU
iL2qGq686r86T4IgR/curA/2sfDOsDFkcP7y2Rd87Y964kjwmhlzLSsRMuTvuG1R
XpSjDxSh0hGP75/LudRyideKX18/w1yii+fknSXglEh4s02YcIf3Jbl+XF2bayoU
kprxlmm2uNPoLgm+4yASL+P326+gxEaYh7/GTRSZ/xLjiKF3vontJ+TotMp4LqAC
VP8ct7oO0Zk+WWZyQeG9BlKkcom1qgIP315yDpzfC/3zeWHeQEcTUEhz3rn6svkq
kcq63sB1zBJDuCidLAKgmXYnljYUAnp/Luen8yjoZcTAlxvKEd2fRuBw1XmCN/56
dwwZOaNaGay6UQHeCR/XfvTzU7y3I4fnf/By/yepJbsey1cMDpiMxc39/r+Szz+Q
f2yJChrRTjEErs3Nnf42ZYxjtT5UnSCpRDNtxdGpk2jOiYz/LM+FA4gId1YzFHuw
pSQR+bWq1hLzmZ9BMO3iFBuhC2XykTkDHDSB5KVnWNw/2J2YLi4TZa0KxtQaGrf2
dSMg2gZ9QD34nwwTv6yWXKUQaDjwf5fFTGBn1czlMBvOphqwE1h8fLa5emuV8oHN
Gj4ZkV+Xj842SSlZUO3kBfAcA25K3NXXAv+t2nMKkbwO8oVlZlywFSMCKChBB2vL
3yZIMLAwkfWg1gK8Whfk/H1iQyiDKZVxWtXxmAsBEYY2tjwTXrCJs8QStNJy548g
yuqjE5U9UD7PATcYmhAqpMPzNEFluM4KDs1ifMtKQUFjX0t8UKboFragvOiE4JDL
UbX3KRUodABQCLmo+I9hfGa28HrcTD/4vme39XByqufqgERPIt8MGL+UIZGODr6d
J4MwerE7d99386V0x8bA3GkFAlabgID2kpxqUDOiODCZs6X63kp8x8JMENFZBWBf
6FdLD+XT+jAZvtFwrk70EDtJjGMZLkgCbtfP3wcxXOLCYL2zfziMDmnRf/sIdy46
Dsm0nL0vkV6VDVyH7tMGVlQ5NROqOp16rI1uCEPN+ou1RVUfqM1b2vtoUVDWMorC
0Il8gilLEhQn/532PR+KWK2xr7cayq5oDgt++QO4nmlBPSxyxLb6YEjgI2OOdT9h
QiHfJNzENChpzwh7uSHc2gDkqvEFtkdvguq0ISrujmSGXbceUmeJgG8I0jZ3u2JX
3xvG5bDSDsGrzp2P/UFjmV2xJKVqDAoTCD5+7UPHVTlblR2rjAs0Q9k3zkgW59by
nxjUQoa/Hm97hgEETGxHLlNso3wzYAGno/8jZMNr7/xOt0TUPiGlm4xhqkT4PuOo
t0+IMuK7UEK6O/g3DeLVaTh36FjhlSKs2yr4h/EhxjpVu0GCrIHN6WkLGnX7hdkF
zgivmbe6FXSHoNmD5uk1lQ23humCQLz5Gsv1+5VHUbEEYtpVg2UprvC75XAptRFx
lMHEL7L+Bt0xoSzJ8BfboRrb7L9KuYjiPYIWeAElLTnc7/EziopqyYaFu8FkfVVl
l4gnQqt55FD3QN8zblOUwJQRnlvRQvZ5Sbz0gJWr16ZmkAutq+by27iAifkXaed0
V/M9rU7/3cTTEatSWZMcmbyWJFWq4sMFJuveiacSwQj6uBq+zrV0zcaPQpGKCIuw
PI/P0r+3XlesiOgWUPGrAEcz5KsikOuc1lq2i4QHf8M3p3zcX3I7EUdchkpcFwGj
43eSjXG/PpWFccw5GPfzLiEN432vKDM6MP1xt7zu2QCqzM8D41Nze1Jiz4NpcsD1
xSVCcgnioTXjgcUO6PfFJT39uyJDyGPIZd7U9y0+21VfUCN0E90MLWXP/0ikw9LX
zLhskLBYcrY85XdsotyeElFOcV8/1b4RLG/8RBFqy1uKsSPSFeuTcfdAJPlXSqvR
E119kZ6w6UgyGxTLUA1MKM8mpODeOnGYkcq33dT030Ey86HiF/FPBknjIaxvGX1F
mbhh0gJTafHa8o1lXHs7Hak2kve8CrxwuvYgRFTti4kz1HTxSyNAQOkpnuYE70Y5
RF/6+mdw5WZoQ35uzoSP8Xn5CylohodRTTELb8I/98r6O1TbYcK++PmR2j1D+D6n
wEL6H/otcKKXQ9rOUo33zuuQ1t+XjBGDRsj3SebyBZdMvXVt7BHYIrIQibQ4JtqI
SFJQqD1eHX9GbefRTCy6/cYQ/bi2mJ838htRUyH27i+LX5FuMdRTtEmQgzkqmnQ7
0lBSSnXWKSvfWn7m5VkvjRTRjqHFgCi3uYE/wQqyro5xYSA/W+tooh766maj8O7g
MQD6Aow1ZlJSBtWDKwWZ8LgV58xD8FvnPmniaLAzYBkXYpnoRWODUac4kF+gxN8O
a7fLsLzQcScVAKDX321hXzsDsYv0IH++GnMatqjAPzFiP0OIhwuafpRmJ61Gtd40
oUZbFJM9MbVyFb7A7Tb1PXEPb/GPovhnBF8Z33dvX4NK5iWA1AV3dcdssk0Z+afr
0if+1yKWwh5b6u5aXn4tpE+dH3yXaPTZDvBym5++wETm3XsHSQGViG4y/oxbqRYT
81DtfnjWgkCMeHN43NaXWXxTuM7xbLt52NxZpRiPzKVYZ524PGFcwNrxstKUL4EG
vUsm8RRC0f0CVun0ZnlQRE2TQFm4UDqO8kr0qJ7vzZSOS1p127UJ6GiEi/Py3+7u
9PpbqsEMBLCRbbtYNagpEg5ZbRxiFxDoGgfrUDeG6QdLHcA4BYFtSvasF7qTadR3
LT1mpJtODU7PVyUQFgCTNjn0tWpFjBNh5ZpHwt/OcpcJDDldwVRRhHLnhk5Qw+zt
CQCOpKnHdUyH3xW0RI8dHYAcu4cV+w+umLGPQ5C0y2NScilHXspkZhfWGoP2KeAM
jF7gFYSgAnCfaIDcvpZWn4NxFdsaXYh9093fe3y76lfNGeMFCBoeL+Ra2YEBSm9R
P2oidUQS1aqtRE6CMp+qdDLNn1pMgXuyp2oHpClhZq+72EIPdePXfneLzStl/q0/
ItdPg9lFQ94crb4K/kNKe4nKBPRBF9sow4N7UhzvmWSj314vckjqiJ/LptNRqt79
MI+plRB5Yov29XZgcgl47yqyke54XcC6lIOp7xOrTmINBu4qoy/0/zUIfk7QOxnc
myogbbLpMoh/K3XPfRBlvX7rHaxkU8wTK9C56PAslUs23rINUzCLE5uhRVy+FI/7
/iIeGMjlgJ8m7ravp1A+kL2/1NttVou92JO+D9ECJ5j4wWVwXz+yBDyqbhjwdmwU
c3TY6UBg2B27xulkuI5ZmwECB1PTBwY4lpBY2EygGBGrSpNzPvRhfk5diSH/6izk
HtNxfJWoRkPaR3FJVH7M5QP3kmpzetfjqm2qjmjCXNttLp6k2za1uzeGg2Xk05pg
v388uelr7NU/V9qzfsfferDESi8O1z1Ajjd1qk/Ry7HzBQYwTqgREYQGrkUpRLHN
DGJ2y0hnhL3m1HPXHKzkNyJXuUk2pZ95wclCfn73UInnaJpa0TLU9OuaBP86bNsd
PQl/R2JJwCOaQxt/lkSET+LIibqx3u8eLfuzRmzqVlTMnGM6GoygGXnmCJ0Ct1k6
yW89JlKMlRR4p24EYHNRLHuZh3pG1gBY38RspoEavhncpfr9/frz8i/9KM3ljRwo
ZgxgnPazCvMkk6m5V5VfWPa1J09EGuRJnZX8pqV8V2egM5N/R53pjPfrNLR+fPvb
Jo5DxqeFDcWlzcJ7Ft1Mnwss48GMfHl27Wy82BEOMpliwbTsvZuIaZHfZY3cashB
FgO1x4iqHERCCd4UDwpO86uXpdNlYTNoCTe9Nx90VIUhMHDCMFyNPOPT9jkuCiDu
pSDpsgeksb7aWWYKNZCMq6uTXJr7dbUOBwJPDRAcVuhcccie4tWl0X03mvCwItjH
0Im0coTQ3ljmnfnbJL8lZ0Bw9HNi3vJ6pyARia53Cyad+1oOyzioSQ08yMtxTzq1
oJ31bqoWjGmDAxD459MJiYx9yUVg4kKuBMm3UxJ6a46QonBMcSmb4RN5qdul5lnM
Cq2xxcjlozK/BzgZBkWCPDJc1hc8FTwUBp6OSoU5hN/46LRr2Gc5nWR8252uXJ9Q
/fogO6Qvf4sjE53G18SRaX6d9XMZM5+qjLWRwU/Iw7uOXPOoqm6RsDIrUOBGbqsI
uFU17TkN0cx656V2glShLwcI1M3FV/3Xf9bGHNPs/Qs9SYFj3u6PrHgQDAVGqfwZ
WMreNkYoOymnDuURVpUgPC2Est3NM30gaACHjv6JZ4i975ydG2Q4xl78xG72f4CD
fVFEZbr961K3W/5w3CtBXvLbi8yhg89Gzn3tqbnX14eJOiRkd5PMaP985jqcsEzc
T4ghM8VfVp8Vq9/8JrDSsOcnzv5PE67R5g0Qnc7ZAcohbdkYWvfk4/uPdVO46bYs
zLQ5kv4tUtCWfD3JQnkFubhEfDyF9MA8aCTGTvFEEKwgWxbCesUhq3lZdI/TVcl3
DDpTx4tsbGiaYkSiQWPe+txlU9IwsXkttMkdbqUhCmGaz8cN5KXDJY13GX2S/ALC
olbhBgX/Sigv5jJuZgGa5TFBnMGaoxu+MPkyUIKRDOrY9JFfCC7ZOu5WCa8Wl3fN
pENC2lSSlQQJfow5CRRWO1Z2asS9UylqL1pZ02hPDiqjNZseTjSvGKYm+2hPu4aX
Xyj1x64KcMw55SKcom8wLC/FhhXnM6fx8wbx0QzLtxzpcyBVEGmnaOxtIBxntX9F
90vQlXctGIlTNX6n62kuhFo9WQ4jm/r8eb2TqeewPe1oZEo1xWfZjRZ/pMtK22He
NDuMSOZGRArUtxGOrRHif35lna7KL4/6yCMDhFemq39lLsvmlVwlw1a79wrI0ChD
ZsWcwmLmmVVH8lefkQsIoF/Ti4GjC9B7/mCxxL4Y/KUXD7UuK5PheoCQoZWanju+
uCzuMzb5mCL6SLmqTckNRmOtQOVTdBXklAnPZg1FTzOlL9+cPwGbtDJO7tn0LdKt
Cuf2CkC3JRdZnk98N/B3i9e/vn9fKucaSF/DEfozij3lSooCxsTytY+J50BxglSH
LT937hu0tcxwR1wJeewlrf6OfO1ADa9dmUOBCkPcCr5Wr0fiobbn27RADLbFju/m
YMEf5FNmwWkAjYr/7fpLBX44u+pzAbejgi2KY15ijrqSxB6xDpKJa2lOmJj8KYz/
4trmwowN7OGZmtIvkZ2jNrkhkokD24p9jsKr9fPHDU4RXkXr1z4Fo8fxPPqNgbJA
9ohKSNp/NeftSeySL5aYBaJ6LmRyxkItKBBsa2Vu5uGeIkls9W1aAKL3v1125m13
5bKH/83cCnq0Xjo3c05FPXG67FSvztOWZsP2beoizzoCohgS06Ndc7QQ3lbH9n+o
ETQotoT7QDIrgR9e2x4tA/umWCP50ucvrIHwymM0uN+2jzdB5wHnCod1TomzePle
mpeLP6SV1PoTsJtuxDAb9/fXycvavY8Ua33Xw9V01vY/CGoDENrq9I8zJA0T3sfq
A3ynaMNs4hPwKSgG/+GWrQgWEu66lrVCwGY/qsOHXZYNzNri9CPNXzQhyPyqF9MK
RqWuYIEUEb3LmlYZZS3Zoav+XtvlTExz6ydNIVYLvR/sC8kGdiq19aC3q5/M9aCe
XOZ59i3dSmqFFUyr3X7CF6b0j1pDt0PJzLPVwriZ+2NxVEq2CtDvfYtnsCSGrQAy
WVl3hRBWZmeIoIDNZqOmkwSyNp547hHsxvy9BHk4G0oIlQvC/H8EmhIDmykcn9lj
J33ie0HbQWzK3jSrESQWACQGLyJu7xSD67KeXZExLeGV/JQnIHjLVCcyHZSo0yw3
HHuEgPD3pu3iTnUgE7ZupRevZAmMrhZpEjotNu9rcTQ/RNMz4x8E/aSOOViXwur+
ZWoywpRamiJXEFAoNCYjzVQ4yeBMP4akawLLAZ2/z93gBn5+ekcqudn+CotG8Jhk
br4pQC8Ig+/TrwdAwC0NX1GeFbUk8EDqMqNVNbmmy1sOAw7QzZdpLejh4KF3Kwc2
9vQcROJWnp+sObANoKDJS3wkOaFE2t5mpB8USihHE2pHblk2cX7EfWF+GFqEpy4U
oI5I1SxjqIInA7fBMkY7optraA2GTdR8qZg+xz6j3F/HEboZPRpLHfhzdKxcyezo
8fc2AnDpYQBp8NwinpVChXO9cYMG2r1DKBNuNCSUE0INw7EKTFZSnixJzvqnsWKC
CotiSXaL6rWX+bMBbKLXqtiM5XtkqRhbd1CBeoz7e6okh/1XaMb9qQs1IWRDOnoW
X/1QmM4cgHMsyLX+oF+krYn2KvH+FnBYzfM5Ppx5H4arGr7PLRDlUPL2VP8w8YY+
wH7NbI+x+o63prXTm1EVaUS2ftlk6MjFDxNFcZDlxBQ//EkAkBgg5+a8s4muAGPw
KTYnJ1+MXMM98oYOSWn2aIgZBaalzG32InQYEwX7xPM/Ex/1NkIacu5Zt8u7q+0o
Jb+/ICPlggEDpG+DNcMCpr09KfIZpJiD/G+dttFL/5H1odl9PRpl/iDM5FxtlBO/
dyGvmqHajE+B1Go/R1XRIClll44mu/RRlr7dgeo6joUGHMw+5pBwkuibI4kOG+Gs
DyOSY9Xb6EMZO2nHdtkzB0eDULGhCONHJeb6uSAOe+LGJrdpTN3PZHc0E+fFnyyw
X/jAsSF+4wzxmxaRFOr1Z2nTaxWS8VoARg0rcTN93zgQ57+1hnC4rN7G9VpYoqEs
Au58ZT5EYI87Qu65sHbFJHNgaClLgfmz/OIP7kVFepFg5dktYeDM0Aq4TQpzdgLi
eIby7xE7ISaISQ9tv+UeQKbvog98BB0MefW8ehPkaL9IQ0G7fAp8qtRkrYq5KyBP
mj9/8LrcPHixk6PkgaSuwg+/HBvLlL0fM+T8tqChtloUO4MZULL/JFg3eXB96r8v
uh1bjcRmL44OG7gp4pakpnJHXPmOv7F0fmk6RMN7NmkuFyDXXdHSJrgqzYej2fnB
7q85ZJm2O/Fn7BelttiVSge9b/Zk/4cApbvkVnVqTkKxlFZ3qqUzE90aaq5/WCPy
aRN41bT1Ky/h5WwDF9vgBG5RLrpVP+9GUfz4sspMkEJyNcoldjrhYS5cRN9VhchT
qEVa55ZXr0IaEBsta0Ic+hBEQhFMl3DY5ij+DL0hyUozPmWZaVITl3R4lGtgIcwb
WWICNQ7V9YoDvxMj8MVxNhGxZdrD98CHGSmktENWBwtL88YVUn/NH5MrpVDrt/UW
kbAOJbVS40QE2T4dzm9oF6CfFJXMiwo5M2Y7PdO2f2EKjUkit9/N/aNZfZThCNW3
BrfTqV3nKZfiItpGWEt9Km8Pf6bvvdC8i53NgWjr3zK11yHMqJeC2VvgoEYKW/nP
Iq7k5vutcc0SErqqzzHJm6vGXhuaTek6ILUH3cobx/R5/s5nVzdnUOENR10qNKId
oVpKtBzGtbkoF+nEzbLz3MR2SFl61JnyMvGNiNDnmfJ3FzKtKaqhyLqJYPhRSxb1
XXRIJLhmVVL+Oi8xnrh3KdEpsJWbr9BQlR6dQScsAxO7hVr4DcB1gyWXsttaH9xn
7epE/DG1NXLhjlJ52+FEsfBA+2QFKD45asRhp2zQOqGihyGkOXDmtAZWMoH0BBwN
euPpATJgEKyJAJVKR1DR1NUUATYhtl4p5W+H5NqtSFpniRDrncaOFH/9sMsUw5jH
Gro8Y9yiEbPUMXrTfHLF5+itHcMtkU8hDrrJyGIjOK1R1pvUZE5XRHis/dIgexw6
kqFpLqyoH6V6G5xv7loYIj+6YZ9BIlAQPMc5vbbvz3zpD4n7Gq3cy4MrPxnnltAT
7Ff+kUkLaL4CyyaBX3qrHBdOEVYLyYzGqp18oiadQWfKud9DOAclND3BXI8AVA8u
FG/J+IbSL6BqKC1CUtGlY2r8FaNar7tWZRdbPbH+IoZ75FqjTxhppiAxB+EGjPDR
kW+UI0A0Rpl98h9swe/sdPSZw3GpsyVmpXslGlubrSlNazdLfRZez/U9nknDdQEh
x2CFia35Dv16DWyc3qRlWwnVw0nQyyMDg0xxBax5ZwGCs9Z0xtPaXV1O7XwYeeR3
oAMle/NFhLfZOTY4+WIdXk7VItVdMvPQv+Aez4COpKJJHQMnG/ZVG5S5f16g9Xjh
hsOhrTPDsXQRlufCeN8AQSFIYZ5l/MIA1LL3zYV95rQD75gTQ7TVxXA+axWJfpXt
iMlmAeV2AldspwSVE4vghdPk+s9mxnXYClLqqvGzP4SrsCnMc7FrS31hThtjIiUw
tolDX3lBv7oJcXBVm/1rm/U7teZ2ZWNWYvyv3s8rNZZjwictwHLZOOS3KQOIB7ig
K/q2nLR7rMvVH0A0Nf1zes0RklgSByRw6NjR5Bt5ztTXFCy20BotRmumZoMzZhvK
tIRDAVJGw8kPFUIcSkvWNgQRY3uRls8hvsD5PiuONPm6F/Y7JSsDy/gll/8Lfuyn
gCwRbOZ6TpsE21txuXeyd6rEPSkVIHzQe4NKh3/SvoqT2eeC9yGJwKCA5pS10JoV
2AIJU8U6uRQiCo32JUY291QvlYN5CKmA4+zhNxV8Xd2Zu6xBPueGgXPq/is6lNyP
XLr/j3FeLzAvWC+6wuBGp2cdhaqDN/bQ1oWSpMz5f1bVXp22szeIuV+X9UxrL4j4
tARo5KwBF2PNUwvpiLhiwvO0pI6tdJNo+AMy+dYaBi13OSdDzRVVLT8AidruCcB6
/8biGxbPlgC0fJ7pR3FA6sIM0fTfnak5lnRZFhwtbmg7N5Oh4Kw38Z62DozS8EMh
OWdBpix/zzzcMERPML/S3x4RFu5R646tR04Pp/xO8x/S0iEOitLbumkNEReweqEf
BE4RCfGyY3LoaFksmaq2IrDE406kSed/A1wnOtgxTCGlJ+jIvFzYXRL900KELvv4
F3Af53XJz41FSpwo/EO5NEtLU2nyGXYF7tIxiRumxDV1R7Zfg0S5EUNGI+AwQ69/
KSffNFCH+UVfPgZP0qT3nbEGwUarzqpYc9fnFP0CVsGrBctrNzYzKWlHH4Nli4pu
+CpbhEJteD0KL0fY/QJwO4dnTe+S6UZvDqUt0G+22/2q566eZZPv6yBFZh+DvVcV
GMIJ6ez8XB6w5Z6sxqHbb+szR/JuSCLKUEejl372lvCqD6uYwI/gnc5QNsCsTABb
6NZ9NwJufQXjY7XkN364yGMmb5UEHc2KG7NE/fSHzhn576jbcJNr1detC2XauQQD
9lGeZwoZ62HmVJZcBLSxPoOHxELpdurZTeQm1wojmRA5H8tMPl/rmoWsuoUoPPkG
kX7q0lGJaGLde4AJhfnBv3kT7OON5WpYiBuKVIaRPn5vJRRF++wXJYD063GUSXeK
g2egwhuW3NqG1kxRAZis3hp+nDkgs+yuTjb46mpylKObl4uhurqkvQbl8LaT1rR2
0pYvwbQNv8yJfv4OGpM6Ll51HW8mazW9yX/i8PzMiT1tK3eCwjUgH6V11Q5vICPN
QCRJ+y5Bploz3L40BWnfPj35H5aqLbcsuA3CiYEAyAiYLgKEcm59TjObZckHif3y
2FKC36K/gm5uuC8uQbTAhJssothz6PMVPqmJ/lKykQF96e6rViP3+Wed7TGo4MMA
nQ3nWv7kklx+TxRsglDRlV4Y39GQly0zIIEOJbq2vXuSSlSeuDdAqUxrhkffBCGk
4YDRBB+lR7EuKv34M6xT270aMezPrwxGZMV6OiwTfZeUEFopvTuYA3bMEy0bLS9+
97SkSm+ntX42WU2DsHquwGHIMPSbBSfScz8SaXaMJDaaPKvsSOE8thSqJSGv/lg1
qDDRogs6p9loQh823MO5o+QysevKXSnbxUOW+HPHlzVXc21CF9Kri9OaYMvoUqFs
POHWwKyoHpCPjj5sSd8I4oJ2SS3DoW74fmE22ufTbRTqrTSS4v1P7rYezrASTXgp
gbl3Di8J8Dwnzbct6909HoWp6og1VAUsp05nPXvqhdHRz34v+8H4VUeR95LG/3a/
CLDzgNJAwmwa1hk6Tyh8X2U1snLCNZycoEzCttEtdg/F/rxCFYi2FcokLohi6fL4
ACxnXrVbQ4cY493u2mBf50HVaaQur73HxnFhL+26KU0brGPFDBGOeiJAxHgQMuR0
ydV7JerTK/vpS/1s7DyGJmhMQA6Ps9lbq+3Y0JwLKhv535ZTx24dn6DahjU2PqXX
Yax6mOveejN441u6+fcrArfdrlWYp4sFlYkukUPxk+8lgdHosmFlKlayGoQsXEvV
LWHr36Dz+a0eOd4RqPtnSLMBE9f+Sj0/1tZxCVwwGxkGGhHJqvykXe5pyQftVWHY
dmlUt9zzwKZVQGTqhymKQ10BckPGIziZvqT9x/ElpXG3TimQfcDfqhGB/utnxOuU
jKc5aw/XzAmCef4nrc6RY7X0bHyzJhXYOZWAL4M7/nnHj5dBDfIGlv6TUxoUM2YZ
bzSgiUjcD268X6HVT1JjDR/3Hv+CtzOcQaIgS19nv/6XoCzdrvSuf1NGeWEls2Ir
/y/Bm/VJEm3jcruzKFAkhQIj2ShUTsatbaOU/XagRpLBiaqYDhtIUdHkz/A3K5sb
Noo9d62pLLRn1TQ/ZjVsNg4K+03nZb7DJR4iVqlkNRBxnVVE2CGe52OZtNC+Zhu7
j0qViTSNhFuKDK9/uBIE1hZ9RoyqokRJj2ZwQ2f57FzZ41eNsIDW2QQZHFC/X1l1
ThLJ+AjTr2yCeKvHtQqMctYJTq0wd/1L/wZQHaa/nmOItLtO0laG6bY5rfYfN1Yz
odmUV/jY6HycSDDmJbAHwGPyit0MHrAGoFb/JpeQmGSpQo6AGvWShTy2sOZDrTXQ
lGTdC+jTNVsqBJwTdyvRUf7bGLWY5VKRnR5pvPOLMwDQP0CPJkBD01YG0/DYodZL
kJ4v2foy3v4AEm32w3NSqRNYLadBQLY+dcL8p1GhiVz1OMibXP9TyBBArkrFyrIQ
syv2HKdZNeEWfPGJYhC0fBOGF0mwGm3NK5UO7miOPxAiYdWg2iIEWW+cXTsiaSis
leKfCRbyDDXlCnM2IcI+CfTovl9n9S2uSQC31DnXtny/LD1CUDh38uSU0FZ4pmit
EyiePvOZwhp64dKbuJzSZO936vrewcMyL4QrjH3krHdFrCW6F7I2Obzl7Dyj+H7W
zUNHMoQBk1aXbmb8DLhBjh1R0KYgQcgWCX+2xfXq2NA97q4istxW5W5QNatxHSoR
R0BNtPLeoJSDddWp4FABH+r6v+NBImmDCnDlD+XWBDBnO3GMYpi+/J6qHqRSLWDc
JqT6v5BW1xQue6lzGoMbymWK8+2HpU4BulDlD3rvTQSpqeuclhQXGkA7Q31wccy+
cd3iuaKVix6KamB7ZraWK/D868skP8O7/TKV6AJCBE0HQHZ/ADh+iWZx7uTr7YyL
tldhUXUYORuU1/FAzsxeKMAExxFfWNja3R8ER2ddAQ6+kbVsmmmQ0Jh4sbKAtnva
xR8bb+rDrMCIMOZCl+//zhLUjwLSfDmykMJUpW9D7/EQCzVHyelRfHvxUAj2dw2R
F6yZinUvw4TcVkdk6B5GHeA4vRsiKX5tF1eYqxwAUBZKYB+RAVChogsGAx6FObXP
gxLhwlwkoIbHvGNcdNbddFT/CKjYPTR+ZM1Wg1k304Szc19euW2PVVPirqPxFdUo
RslvF3m5lEMHEv2z0zK6Dmmkx0T3fYjLr80Oi698Z16UC1Sbkf0XLkqE3kbpANf+
h+YP+ZA94ORqIM2chHA6dJSR1lVsx+ouguOerQZvj1VtklVoDN8y2CF3shYcc6ZE
01flNB8AOk6njvOoMF3PAIgAW22RXg9uEVVOMh1eqhGkwNVMatmQUIVbW1HgOUWG
CarEUZGOjhyzu+jJ4/ceNiL10MX7dEqodmV+kvNSWG8yjZDAiyNfQZssknQIHjty
7KPMcwAf4MMMeeJIRmjEtn6y0C4c/sQXdlQ3qtRQVlOi5x1JcHrYZmT8LSmFPnDF
Zc5C/q/1yNOD3Bv2xJvNxk/efIwlkfeyBVXZh+OwhsNyEzOaYVteA1SCwJ8TPzl5
c7yK9WthJ2hbZwTfsJmGk4PxVHNBNoEwfHroPtqUdtQW6dBHRY/ljS/9SfLUvhsy
LtY54m8J2XjuOXJxHQnquKZpugB/OPRu0OpatZYw3r4FaLDM4prXh8NJhtF/znAZ
m9Pv8ObV5Byu+m8/MMratpQKaZ+yNEBThnzKVIxGGsn4KtKPjLm0y52bEnuOnzkD
yKlquK8HKsigHNzE02wFRsebXWNLoDDf4zid11GZ111t537iUfGUjdEGkNMOWgYC
58YLdG/ivnuvD2NL6VfrrlHwPLxK4JS5Nw4qEqv67x/DbF+nANxfCZevBYRe5kQn
mpn29pK9vcHy+zWyPBCi2AWcg2XmlspWPgUIVsVpO2w/ty+LOjDtM2U7i71qU70u
9u5/dmNI6R7opJJUWEO08LRQH+5YxJl1qxHunW9r62eMLhRun8uhf+KKn7/XOewm
QXoOtY6O/7MHeQLYu6g9R9W8nDJro8HcReGwpAV/HU1NSfYZGkxPPHDSPX/K/19h
HJ/6Ws4F7lLK5AjbeuzsIJvfo7FVhdjzbmSAsG35oAuHB5OMG9vXbVrKLygzZ08P
Mo7F4CM3G4HSxx+3ngOCr/MlYcpDyT3jc5OpbK2JfHgi6fWxRhWVCiLrpxLVxxPN
Ez8cHjWQ5Jt+m3qOR+aoa0zBdpGvZkfOaD0ElF6043XjvEJt6dMvdZDRC1XiWKU6
M8gu6M80M6B1iZzeyDQ/PCld+bw4usPHNAsiVNjoRz9Zvx5VO/SAC0iHqyQJGO5r
C8h1zPT/rC3b2c+G5byF2pdUJ/5lXY1a2Wvm/PYv0p/dMZCXkZ9o7tblJVAUqQSi
PPrIz7t7jpb724IIU3g2Z3H+FreeKLtS8AirhVennkttvmOlxIgGxjP+F66zZCUM
k78nVgi1kp9uVMrOmkgk6Ni1TlAUxMJtu2UQZDTHcPc96a79g2aGuwz3dOp+OOyx
h+LrN84DYhGePvcjsIgkfF259uWKS2M9hoZWoRYiGQvfZ+8oFyzd3xo3NossMYTF
evDisJKN3J+H8d6jK+qugbhw0L0u3lxiS96DCe7T1bNkxzGSl+xPHEb+G8jYp1MQ
RDk0d/g6syQzAANJY54+bkgDHNVsC73zofFQteF6A+m1uJ3a6kN5D/ctBBbxEe/t
x6UXt4xXpR/kg6RZXQvch467P6SNdHszadpY4JeR7UHN1aLSS3gfc3SZ6KtmUDl5
RJxdigJqT6edxkIuGiY8NFaLwL8gnLW8xlDfZMs5AOTXOMz3pnfRylUa2/cBIM8g
2/1XzC2k6cU/t3DJyVdhjBIdkSfp7/QssMnaof0451qEIgUrBqCEQ6JAbgZrSOBs
K04a+fJO/Y0l3KH2pFhlc5UHSp7TflB7LALz+mAAru7vAFIEABqtKHpHSlrp0YfM
g+EpFYwdz7R0uIQzR6DiHBpTuJPnWCjgeufFU7O0+hcMPKiMUgA2HSJ4jTSmNeM6
hh3EfA/ya9AXJO7wsa2nhHxNViZpggHWdbOJjRRnrOvLnG7svqNkhx/3WjHeg65F
NoktUyDRM8Ao+5cHnXVyOZfM4/qazz8tJl+wwH1Xj8/+qbi0y0BWwDV9i/zgZpOx
6Q5y98qgpqb/MU45HxJSunanpzRCUERaeuSOtXKM1U3ZvvMh8iYLc4TzM6r1YUcD
6HnjK1L0rTqkP/6Uy2vZ4Q2qQVeXFEYiT0eje7/FwOFApdtBK1EQwwpch+0fPs59
yZSLdl/TNxe9GXUCCYCMFNPhTriyKYYr9e4A0OYmcCEURdLg1AxGU5x2A+sVnGQy
MDQmUEzC40SbcQvc+bHwMCd04gA2d9XDBmr6PA+ufVkVSqKPaW8gX52KQjTYNJY7
nYuQb15M0xmG9c0zAclOn3Bc7MlAz7gliftjF5vLZ2tfEnxmvCIkZLyD82k73IRQ
Cjh4HPIxvlGgm/qwX6jLp/7Dhvhpot9/9HAnG0+SQzZeRIsES+4FGPMy9glwUXfG
3xzavpS1RwmiSRd1pZo4n2d5VYCsqRpvIpTo/WZxKlfjNDmHNJxu7VX5c10mHEGp
/Odzu5Vko7mLM44ib1Qux1udj0w6HxnuXoSt2VDuDKqeCb1RM7vt9HGGMBPY7iV2
ajkp1e22DBLe5fx98Ft2oKSCT90d7UzKp2iLx+GBJrMFAXIPKouH8zebtrs1lWue
0YyPcw9iiY3lQIuS2u1i3BIlpD3l1gYuW9Xzjp1OPmxtAWjhlzZ+Jo6E4fmgJfla
3rEfFqF6J/cgdOtZ0RA0nz769DzRQaROCW6eq7z1lQKDERu1dR7ma+iJsnbLBIEt
f/JhtZK4jOHPKTprZNPdLjl+yyhrr4HGYZ1ifSelboj94MyCj/H4LvbyabaXfvqa
bnUOTkyH3A7pQRnEvuuUhlsOhAzS1RrAQTg8C7jCtcQ7qTF6QwYnF91A7Fe/H/Zl
rVO4Ar2vftf4HxIyWUbBCH9IV6BpJ8F/A3Z9Ts+K5B9ICEHN6s77NihU4H68n8vd
rlsileHCU1c8qfnlcTmMbUDU65IJ2np+iETqZrFbzL2sLck4sI2ermmM3adfC6K8
pJ6POQro3xOJCqDQFbEnSq0PKvKU2/+/YAHSLXAEfvI76fJBRvXRQ4VGd11qbuDk
6qs/VXqYJ8z7cABpWI8kBJx6fISDLtmars3Rdz27bEl/R9KRkZdVas3jQ9vQZEiy
PdtpDzYFyw8HXbNNm0agTEQPGWFKU3xwBc/qO+fNQNSR7b9ReBQyyi/VBWogeY5X
xOeRfjvwUkWvomjJikAeEIhKrmoboEJTBxFZ8vmybsR+bmMUjDXvSMibJVb5xUIs
Ak4WuQJUnZiidPaATRPNSRAmM4aCO9cDhg9rmcZHWWthRQV3RFvSgpork/xIp67q
kZKwGgaW2s11mUMWv4kfnRcvx3PCY4p7wLiXAG5O6B7BIf5cpKZ1LfHRgE5lpmXT
K/r/c+qkZ9XWucd5R/0iR2z05UnKlzoIbhh3FUzMatQC8ZF0775igEFZzL7Xh8zG
OLMbdRupOUd4PlHeylp1A+MKHlBeL/KvPdWkpZQ7qARYnPk5vD5K1w4ZfRL/gB1z
o7dy+xZLuptfjJjHz/biYIx5Gh3U0iC6nhlUkCjn5dNf+DERsn7uuy67XKIMO2x1
T5/wakqxdenjiUmzBy25NXNvtK4ABwjbsx7AqOXWCDvDByLuBEx3QoHS6aH619Cu
Cyjq0ihJyh399KUUftTk9HWzWJOSbiQdcetSfEm7YEb+cqTJWnVlDtBXBCDgn73g
cs5+M7sK9oIcPtlklmDlt+9hQdWHp+eUCOnCuTrsMVfMYCw9GPINStgF44pZNd3w
P7npNRZIxYwdwVFrWiodA+a3UPapuScP6HEBW9EeBjed+03c4RumIVB0jyb2qqM5
YTu92iexp8dSS1uB24aTOmKXvKQNa/Z2YGDYqCwUfKJ+sSt8av+qAylL8KQWAvQj
UOIy70HI5jzwn5AYOBbL9VQNyf91LoNhQQv06wyzywC9Vdd+kZYE0LjHyEnkdvK1
7mD+jCzLLm0KqhRqQlun2hjf1rGEvKmlu38nIXQmPVlFGdCCVsnWNWRVDZ1Rd7ug
LiIxlL/8IYS+dSQzg1+CWbTxiqhaaR/ffguHWaMOa6qkf42Zhu5opX3OnrS8al+J
XEnxCJAPPKWRbWc0go0vwOMb+niA/EMRq3ctbQ9745LGVH6D4DsjAv56WLhIrKkR
EIYAmUme+pBeK8vLbxpwRUgv41iFoZ9ldVmrMpkWkfL221V8X2E9QvADrjTxop5Q
X+90irScUnrCx2Ko65JkhgojpFdDX0miw7TPIiY1zfrcdehRJ7owv7/AfYLhKI1v
IM6QG6/BJM5iVsbsaOD3wuJAJbjUrwkRidJQNQpTfjyDrO0jsFIpKl7ULLL82+2R
q/SrWpoYGCDqaoyamsfE0XdJl559eeK3E7g08uSCsOYQj1INUdRDSoB5zY9VqSbf
pm1UmS1QwSzGolRGMPjw89WakdBgFYsz3epugbBXAdmTMzNEKgmWbGeo3fc8kQnp
PCdui3wVBHStmdo3Xd46fqZ10SZ2eW/ny4Md+uHiuVVyNktAhDkAT931DMFnG9fA
P9OZAwICHjoITpvwRe6wkb4TMj/39H1sxKdW7dNf1b3xSbiMtxI4hDGm1yvtCWAW
1U4dzQkIrIL2I2DfeRzagZYryfB9iCms5e/iZL2Dj8S4axKSPVgacw5ae/k5kWjI
hbnyrARWSVNpeIb6EJ2xiPEOmIBnXd0TBaUXqngRkHW/gzyNlomXv/q95+MMDQmB
1DfA2Y/HDHCf5boJt7y5E3DVLOUz6Jrji21nvCeM1Qbc7AzM5AedZYpNQyivSD64
/0dL43AvWviiUDFwrK3tSLvMcJ/WI9TYIFk3qNGHqUwytbAU1kOmwFc7oDY8pTP8
vreG67LoN3tXzTDdnWru+gCHv3elAeqM0Wa4zJ81nOD/vsV/lqaz3VMc83FJ75RT
Xnn4TBPmeHTkxw8LQiFGtzPY81YWR1j0pp+Th+EFbij0F7c+6JZfyaXTbar1XQdM
LSs8BsmluShBl/ntb9X/b+bhhLwrGeJCvzzQ7GgKB/BfXTJIYuoAvVsKCaGsmS1R
eMiijN+foEjKOEwkSCtVMbJy4yfWZTM5+qS8wbNBU/QsglvDa15gtLc6+gQ7BjcQ
sNdTP5RHsvmoaLx01H3oE5ugNHGVfHhQiHh0a8ROEzQFkmjr11OZ5hyIKpVRkvxb
TkoCpbwpGlrt1AH4ludLUwA6izEJGRSiV/Pd5hpue4JHQoL2kjO3TpndIwuDddBA
tHpqFudcxdfok4Fr1IN+q53rroivVGDtGMdG5n7N1N0rZiyW1PJCcf8y7iwdsQfX
a+E4v9+3vNUtcTLUGvSP95siCVufN3AGhaqIRQPliepLLriPbUX10zhI5Qz7IO/z
BaI/O0PamvktK8QYn0tEDXQ+eDD3d/ejMlpnpcoyiC04GrqHJ9icGrjmCwt5aNTG
sFeHeRCtCZxvQkcCpruapOYUl1Q0AVumNNeadQ2rKTEMS3Ak0isJD6EJZp3F9FA1
LMwgh73GNowf6qlFpnPQuK3rXpy0IgN+ei0S2jsjl3/LKVAI93ZJv5vR3W3WbkZ3
ZDLFs6/aAuw6xTF/YGQSevRK9tjhqJ6jPNoiicET8hZ2gY0Hs8c1m4jyjbiHK5ZH
nwSOuXCnhZcgpfPjfLlQNm4z+/5GAogF0NtQ4QShvY30WCzlMYu1LBsLZnHuHL+C
taDO7378lD1SoEdw8GzkQxswYXSUXT3kbo8Fr7n8z7ZKTjxhnJ1wp45lVxlYCDW5
nfVbth50kh8naJzfQMbez3RgU1p5MHIHA3GucfomCzyCI/2WTEnbhfK44gIGiumW
gyBm0GkzCUnjt3fKFfXodhbtMDzAe/2CooiBOfjP7HvYfj6WE+jJ6JF4cpP9LT3r
IYZmn4aeGsEwavM/OKkvE6/2baIB6s13nxBQsm7L4wBPQeUE3w5EtyXbi1KasdEx
Ywmu56xEiEJbyV6mz3zqzYfGucFTsUcwe+xHFUFgeScIhxoLe24T75C1jNv2RXx4
1deJxioJQLg5S0v3jDmmp0izeRAAm4Y9LVswR/0KCSJUlX3ZVD/ZeiVK+9xOSUsF
qyfpfRMSEdNbEyBdJeb1T4M2CSvzVDw5E1OiNzkNWT5/I5T1dg6E240rnWG/1+ZB
zMP8rFMIkDAZNdJhPkQijtbU2F++u4KP8cvQfRDFlZa2iqklzak3cEfk/R05aJmX
PQKLGQRl25WLp5G71Zes3cr9BI6t7FmC7w7r7Rq+7RIBvQiT7+ocKJZv+/E1P1NP
QiCwkEgGfD8zt65rydlymiGBDFYNqrtfIiTr+PtRrdGNedpH1zGN7ban5nKMH0Yr
NBofhOBGtNC4MH03f18v/rRP/fgX8UlOzCZpr/dLzTiuFAq3TXcFb3fywLbAdvxx
35/2AFmIbdyfLAWutzmlsfEN0Rcp8fwOBkqwzO1656si9m/yTcesX4rIUk3m7cAI
SZyIPE8fPYhcZUmCEajd81TU7IOdF0SuwjjswR20/MXP8aV07N42K6RSuy5YcT8u
ittW3HXCbgN1EGZ8G6kv9Ase/fz9x81g8deYoY/cbG1DQArzTM1w6a3KpRqKHa1Y
O+Tnp8K0X1Bcm8AVH11nB7esQLHZNUab0aP01OUKL6uQkjXIhpyd3OnO8rgve/fA
DNu9r3bU8M03yqW6Xh+jKXTH8A5DgXmGaJYfYU0szgRNDd/519/11m6k5ZiZKhlc
rpjdpehfR5VU1dc9r89gmNH0rkF1ZeB7q3SMq/GkKRMLFIRnJVs84HSKb5JjvyEt
k69rzCBVKayQvG/QHRITeISHu6VcOuK7l6JuKLqjHhMlU1UqmgA8Yd9btY4sRY6N
OUcIVw/DXymsBgqEayAbe7WtIjnlpOzrwfQQkNTJxFZU/qFB8jwnUJoSVQJ9E1pZ
tpDbgbaiE+2YyZpT8YoPL7hpZQfKfISxCbcVtL6T6lVMFDoLEEnXUMdwu7PA3DwA
fJTF1rXHibb1dIo7En1Hb9+vygYv0Kh6S+VBsCuCHjun1zRZ+HLilZtWApBX9iWM
YLKPQYaJqvgfmke08rg22k/dPmvdpfzDbj2q+IznEqzr4ozfCgE+CCklelh3cQLh
ERBwTUBMjlhd9AOG/WYB6noO+ul/2NnSZyJR+R4y22SVSrZebwzkG+20luJD+eEf
SC/Df0wjdPtcsOpdY17Bc2UghEsJyV8UHerC/XkRkPT1Qn12K+247eZq05WhsNio
DEa42fRFpKHmOmloT3ajWNtNNGiJ6+lI81DjEowvEWKWT9IcE2pCIBKKBKg10bQJ
xOFUnPx4r80mlXIZrUlOUSjt5ufBqL6IwVP6KR/LrjHV7b5DaBZBxQdh8XWM4GT1
KYpwqM2LNYV2KMMNndJTtQ+9+s8zJAxYOQwuPE6KPGGjv4YSSX4tpXX/na0RgPw5
dgErS6lUWRbFrIlxCt4kfrVRrzwa9TrjuBugkpp+nggqFVhV9HhF1iLbKPztVZ3q
kzszJdnDQd3mAqgJtaWf2A9092x+WyWWOYRNEWHoqcPXnm7NZq7diSboPc0W7SwE
B+rBHMNqbQxS3vn/ji6UBgHVGiSRl1hNLFUcmiXrSTZt9BUoVnqdvs33w/kDVY/E
sDIEhiLt6rf4HI5HNzgS6150gMZx8mSCt0faE1IloOq+WOLjNGwOLAYEHQfIYfEX
jgKWv7mtLAJxQlkYN7wHtmprti6ClrhjJ757dm1IgI0KDeV8C880nwe4UuSOLuTd
mkpNOJXAa9Qp60wQUGuoU2PqxE7brh7oeiPP/DnybOk3jYsvBJCYFIMDblpV4WVT
otwuDVhIW47e2cjvd1WLreDctENApHgkTK6BZvE8OdALUBT73UmqeosINKrtxfTm
BYb6JmxYAsiip3yBwQ9Dge0aTwzv8cy3f/GR7T5R21HoX5tl3aUNkFFyubpAwqUD
wBFzvPoKRgd83tP9iIz+QGYR1WwYHGBN6jRZ6NDQsKhoDkNk09CrASXgYg5t6Qxm
7dxNNS7RoQhDjFGejcIX7tsxLim6mUuOcfAxga0fT8SAmlPCLdGgZ92tuNrP6BxD
ciy4fuAcJns/ecwKtbMrruxaLuzn17Ris7alaoRJJyCiX5GR7p4V16TzhB6yzkLy
SARkaxbkApyLesqP0gHMlozneFFr6qOqFkHFIfwMkhEyWIlejItz8yk9r/PdXMru
biIxbmUrReDTrIXhj938sqS/Ha/2Eb81BrrN1LEaIl87PznCsDuo4LKyi5DNKQNc
pelQ9gl6nBoeM4/q6fTllpliiSU4kB9etGHfpvr1DwpqkluifCYgQniE2epFyRYd
w+nPzA+dU4h7YFSfOetYasGXW3wFNd4UBT+moyqL3Xo9Up6g2i5xizieQeDB3gUy
DDw1j6mTyQEfksoSemCJpsY9ZFu6PfCB6bQTPkpLhEPZO8T/GgZTCzNzZQxl83N7
+7rzYdAE8+ZEYVYrNY5/NTCpG/3AvmLwGeH0CtEdMkVwCSveh1fAM62aA8KDj21S
K/U8v6lihoedjxRtgdpOH2qvFqHupKvGV3Abhrw3Z7stFWnk7TeHcRqAnMccu+Ra
6cAfuqNHushccIk+KvPUHRVm9mPmPOMXHeqc8TlQLqk14Xuauu2ePN0nJ3GE24Um
AH0gUzPr8oB9CcZ+PgjUwBnG6K5QiOvowHMse9uTFnNR3IpAu10mc//wdQeLlB4S
z9gCiUGxyY9qHgkT+zZXAaOdTkAcQUtt0OacER437UlKK5brbPUX6vW3Y6Jetfk1
Dd8IZpSkRxgf/2ZpO6sM8uZpZevAIjIg6xtnYYFb0U6Bv72aKLzcAiSLMu6asvSk
PHyfVvI7erpMMF9Fr2v3oNcQC5pWDvVQl0ySD1kWuaIi+3kSkUdm1KzLEyfnKjRt
YX9H6o7oABKdg9A2Cmh5E7d6N60BzRy2EYes3i7l6L1fcbgTFojLMBXytMapuVH5
L9/0dchV4B9HFbVihOUmGJ++wZvkQZR0RdxG1wjyZTInPTGqumdZ+opxzusSUR3k
3j6/Ix9On3JDF9OLPEViVFahUb1DxTmNHqjHy1591PT5n0UPIdQlKdo0yHr6Ca7W
DZyV16la6/rurdp4Plv/jUNjT3PQIgJ8fELr9fHQxVEoaJAfJ5mPvsbhCmZ90PK6
HHWTfeW+RPXW7ud/60zyzGN0UmQqs0mEn89KC3QhR1lFKHn9NEvwpgmyOArrimno
HWS8aHzE0WvtuYl+yfbxrtirRtzzyHOaI8GUx/R0u0WJjbB0MkIFLyWj3tnXV+LC
FBVfeyplYNChze2vjRn4RdM6cJp0VqehQTqfk1FGJ98QkBoHXgT2EaQTYyuCye1x
UakFqUe5V2owFDdtaQCUNwk/zrYZbWUVfzRq66G9V62juPTMZ4vepEnBJz3paWrS
XH1DZhkb/yOewcMzPs+kzALI9hR7DlzYKw8YrLdSEDZYTktVis77MmFrOGMabZ27
itmiQknmVmoMGuQTSZR8QSbJ/xiCzU7S8eZOE9ad4gB1t9whkUOLVQ1WjXsqFT8u
XGb3eLnep13xWYkGfNePwaKXcHqjMrfiQdRDAic4elHXm2emHOjHV14mwT9Zcyzx
krLlGa5rMMkI2K1qqLkMKE1ZmK6y3T8Gk0aZ1WdKlJWsfRl5GbZdA3avWKSNmtnK
1JH0sCyhYkjCQfhorFbnDvStHeGUFRP16WcOqW2C8cI+oZEmOiOXqlmbX1z9trEA
bNiTLgU0DbaI5GvZEF7Kh6apL/9Yx8foxzJbAO3evWSXH6FLEHqam9BDgE9n9e4g
+2lQMjBgq56nBBnxcx983A9GrcGGFqY3hRH2mioXB8ydsTzXdrmK7GjaRihis6jB
7kNCEJFNO1fmbQ0X8xt+pUsH3XD99jMEgvAFav7rnQzQXkCaLgNmRhQCr6tTZqT+
jXM0qlNinfjc3yAaNYQZdgPudTuEzhJIA1bhqqXQf5c6oEANSKHCR/ieUoxTbuJE
bCtYzNnmqqaXQL8ugZEn0CpGzEM4fsYfn+fdYQ0QUnH9WQq+tyC+ZDkFLT0Msy11
MVQQq48xwavtUr8t9X4Tw9rwxYUDipbYuOmcQu+6gJWJjFQVTi5nNaI1df6ZwQOk
Q5B5rk+x6dKmjFYIFvCnRJXV/WyDIxqxy0sfMT51/wYISO6bXBKsipyRH6UoKsgT
CkqBj20C+Z0Q/5Sku75NMQsFkv9EWTCPDMp2zVDWMqFyy7uiEgcdeeIHUOrOzLjq
4+X3cmArUMcTMfD7Eln0eYEc4ZR1eDRghQgpCPReUbG2I+XI4so2nC/u5hIVtXGI
XF+0ZdeQHGIzIhAFdSad2/BtQh1xwFBAbpBizP8eNQGR3I/9jpetr3KgVm15tEwA
JC6WfWYLBy5FN0DcJeeFickg8Jem5MruGlf159MCHZMDWvH93gC8dU8boGLy7CKl
+UMEzOw0gaK1OWYmFbB2wRfTJoQrCYUHXryPYFFpirEhVbjeqvq/5VcqlGj9dMLz
U6E5WVObPg8nXAkvEiX1hxxyq7qw450xDSFO5UHrDKr/X3zwQxJ5jaYIwiTTK4Pc
zARCzZYnHu+nkYOrJmpkS7EPe+gwUKCQIi6++InDoJeJOFx7IPGMGgAI0HIdEK3A
He6LrIb36qb94jZJ6lncH0t57GPF5pw0UGCkfwnC36O51xVG4BAVBnuwxKSu9fYP
QlNfwPLgtNWRvFwaDPdOVcIa1PB+4jEas3qegxFGo8gS1f8LWD0wM+paoUDnLN+S
klDHwctJW/ftVMTaDXQ92+ext/0JZ6JwW0uGbUW0IXFPf7cUui/7SrR0JgRlG1ZD
4+j3S1mtBfIskpKN1eoDAVmxQuXwNZg+jEuPnaUx3Wu8Gq8edyNQceRiDYklzwKg
zD1yXyzzwscyBZqJct4bOm6T+ZVY5hL87Um2AxEe/gAQvNZgcZ1NYCh5WlQgR98Q
hQd/6V7nNFjWc1eOmz/X54/Rmqrn9gIrT/xT3zg3PLb0Dz+pW5hJv3M4bqdyoJBW
bqbLuVOX1IceR14yMU+5155BKsE6xjrYjIkqON+qcdpEplgodHus8cRrSygG1DR2
CWbFSqgj5anE8d4WpWZ4FIxYrdt/W5/MBXZPYticZPbbQ+hGwE7abpp9BWRrPvom
T+fn9+9uscmXbXfttRuF+wxORDholl+wkyqV9Ihuxhar8Af1uofYrmYa8tOyMiR0
vWoFM3xxJ2M/0OsF5SMQrjvkom/Riu7jUWziBwbKy/srTTZTCaCCmrQ85fmrazMg
hJESSQvUl5cetw3tjtksl5109sAgbpWylNeAztXPWsstlS5iN0H7uK6Y5c6bFa7S
/AtOh9/3tr813tawVyc7OW3d64RHR8PbYugaSe8pLtVCtNxKlKC39LW2ygUF3ery
/nIQ4gBBi/lh/W6/KFoLrF2kv9HCZKARBj/zsJcjvcCP1QULzJyAvKiOfuZcZyKA
OSy1znFxuqCiVPr5ZMek08HOwmSdMCIf6p7J1cjuZ62mtImnBDh3Vd3lDrKf428C
q+22Oxpc90+5T2PPla0pzU39DXnkBJ8pgb3PKS/xyhrWvbbI3mRzw1IQLKrGoFNL
5/qbc7MBuoTkNxYIsF9XI2tNP5Ux2kOBWVAHymmxzG77NEWRv5j8amNk7PcUd0sG
sUuks/vlO/Lhzfm6dbq53Fk5DPphrNrLKGPwqk9tVDdRkB+Xx3iwJ8wJrFyKL2Jf
4H6q1dr6lGD5GSp78vkfzcydAMebXHSvLk3MMN95Nh4irRkTSDBUbrdHbpv22e9F
ccxFbDfcaewZnhHZKJOg0nHI1Qfasrwkt+QMfeajb5xBgf1snB93YszjibuTLcHz
GomJvFnV+FkVyTVGUFZakyHY3ucaxb3qurGPotUttALTVn7vF9OsYcpdoLOLZmZ2
UnmVedMc1Em7t665ZBVJ8ZpuBn58zLRmHcP7bPfiuJM2Jf1W45TRyFeyskP7O72l
WmyF8EFfLOMGbAgZ0V2xnP+K6HOTgzR3G6Gfo6OW7+B+OsNmWxkPjlssrb86lD37
ktAamg1+1MjViw5zJDTpm1X9MDGgkanJoHvigEfLXFWUWsr5OZzTM5ZPr/EsMQK1
reybsDlD+/fsw4vUK3XxJJ0Ulr/E9aZGryQeGbQFWP7kqY9MqAMgZJq9Q0cHserw
mcyz8chmDwtfvl0bjABwGQhbrIqsIbf7eB1FoLtkiBBObOE+lpxsyA0v62FkQF64
j3UVqN8JxI67WcACAKxE8e554Jo2/AI0SzER25mtBAVhKp1Lb+HDV3zBf6RuZo0b
apc/mpQeF94YIq06LVttfjU6CLPVJYQk3yLCLSTlWNIfhPEdW5rTm0Fht2dn4Emo
eQyfKz58cwnidxWFufHBfm5n/YNvQTkm23ejIgQBjIknPtQcgViPBAmucaSCHC5P
Af64KN7NugvFKV0J63wjI18hd0kSq37SAFS9mkujxMvoFrfmmeIyhITMy2SD+VlI
03th0a6nVxWv+XkX1FBPhCcZtZ7+RwagpOL7np/k0vDFhHnniVU9Tv6d6weQU45Q
/Qr43b02odo6akNQ+A1GKd4MsbasUpf1uYL7pGBzHYZ/+pSvLh1du9J4JQ/c8Nyr
Wh1S3Zd0jXo00BYBRvkEpA4YZTGS4qCv/BF3FxmDiIG6wSOEZKsaM5yIdHscZ0pR
WZglw7yKIhqvrBQ+iKzn5ey+2g7spj9xaQZEdP9U64Tw96Fl6EbftsI0JGQrSg69
8cttXen4UC3bi5YK3yw7cnr1gjpZdpgrdJiQu1xZL7rAyFFkcqgaS/4JbJCDRtsv
jqECLjDFhkgw8BpVYJi8zHAj7yFHRAcHn4IJk++aiJUMVcO31XDv7e+gATtd6L8k
yaIusBMOzKOGtrObeKXMf44Le4a2mW1ZQaPPYTKNmHeD/WQ0ADgK+AbYdj/O0gtu
RXZ05zQyg2VKXGKlf2lmXeeHjDQVPwhCmv5yHMD5i/2CITflUyAPdnIDkwEumzhy
nj9mPXTwRUqIqsp75uk5deChq1CY6dHW75NAs0kApAkG6UXS0lP+GVX/x7nTWDgl
VK51xBYECU48Vk1DmHvVrOEIo2jDKYypvVVhOkc62SUvZIqOCI88hfeVYyohkSDk
mceq4YiBGzpfYBvAtTj9yqD9pttYJYvYdNXVbmTUt5Fg4bBxTsSaAEoL88KHAqxy
eoyM9VMjaGpoYMr0rFbG7j3AsbssgqABjyzotQ+vBuLsTS6kBHyPsgsukEZTpZKs
pxR+EfJlFo4SVnf+hXFGKAdARS0a72R6MGHp/z0wcvLqaRfPcuk58ubEC7kFrHB2
8MrI9pLwSVFIwgTXSS8EOfofHGwb4dwjLkyzZJkSpU0IeRw9tvx3KbUN1yvMxCY8
95d3R9cZ/feRxx5I71ls79iuxhMxI7Fu1xMonX3lQOj/qQlPkiGIAHhDx10fZRjW
pZ+ks1/LLX0/geGlHcVeU9zX6OU8zUgcef54DM2zuXFr5Pqfn8OVRQAa9ElgtWtR
XOWJIcdVN221+FaDRVuzeP0wGxl3/1RUNrCTyE6hnPztswdtzQqix0GUokg4ZFUv
KVElPTMylih2gX5asafFkvOYenuPxUfXwAyFuijs+T39qCwhD5exP4EPv3zjeGUb
Jh0EnsDzs1742eQg4BhLnOpuuxvIPmd/I8M8mxVSMdwetnHuWjLM5z3KiP3HXar/
LCVU5m/cr7FUsIM85dsZjjVBCZq+mk3bXHNB95I2OH5h8rkiXSt/lWG0LKiSn3fL
gNu56nQcbm58hl6Jw87RCcMDA097msQhi6NQ8HLMdrcHQbi5ADKZf3EHJ8IJI1x7
qaZ3XvpfH7ZknBjUIbGBuiy1ALq3AEvSCA+9ki2y5ppOZxBYaGXalUGl5yYCU4Pp
Gfeyym2YaORRrIT+LoBCTi2iNbn65T7Ikaj/2DwcBd9weTklemCRG3SCoolVwExs
tOt+hWpDCgHsDXzZVXkX32ikvYULRE2oMF6bt38V5FvNM1DvvmPou5ow5OiyX9Tj
jBDolnxHPAiv8ita5vr1tuKji4jyBUGhmxlL1f3OQWHdYIy2ZZmxlJUGzXIqAa42
fVxFsnQ+dHHBfJ+G2tKqQFIyGTXD/NZhQMzcviFgiw6GjCdIOX36Nfpq4iOxDeaU
as0qGXR+Zv4R8m1XHgC7eIls3q6vaoh7G7at9w02dJaFvoU5tgCg2xT5OW4hdu/n
2nzT1utijxG3ABfo65ftD4cC63bC8ZAE0gOUGuxX9Guv8fgiz9XBvWU+zG4//+Jk
QNNja5kW3r/WLOR8K5i7QI2CsT0xf4hG4CF0CwqnFO9FNwK57ybYp0J0gag61udx
5s1ahMqq11N1RMGE3P7rid4nmdS2ZfjdNV+Nc5/uSnwPuSwSV2wrKa00G26wL6pk
q83sqYo2b7rpmJei/Znyu/aEiiM36pvC1I2/IhPM4XQl6p+psEpqkajerlkEYIRh
8GwE9R8s8sr9nIJ/vQf/r2YV1PH+KhR30Z2sKs7t3DsNx7rHNYaJGQAca9CDB8gP
jOXxGmtOaeZpqSX3o+zKiEeGgLD4NBCBygzQdBh4TjDnXm7YG7BnWgLE0Zth1SnR
vlmx5Dy/A7aXM4D61ybVj+QAYKigsxcng143uLJd7ELAO4F7Oeq7W8+f/f1C2zK9
Uackf7+sOKvqRfqn45cSqeAh5oAfXVIbdqmKM0tCmHmh7UNoTiQb2ESnknuuwuPn
sA8K9uiK+E2xMpWs7YrFsFvzR/j3Xmf1ZnXvEQxxevlggognWSJlwghzwG2BL+V4
bbXpMxl1afsrR/AT36j59YFMsJTWRTs4vfI0AKSh5JKIHyMnIVBSoVK5ZZvga+xs
5iAXhdwoXjgw15G03IKnPur+apn/6HkTLFByapoGwX77F7xFV7jp6q8MlS4QCQXR
czyDj9X6u7zRVM41nfIOTRUurlvj/jRP6b+S4ukcsQs0ZYT6CYCXxiXIKwe3Q0DK
mCaiVnpUiZZevD5qys1z6gFHXNypQATl+/B+IRzDEAbVHs7VF5D6dFMXKIzY3Sbv
VeCzlh2ExeUBCtJqjRy/h42d3p0HvoHUi1FLEk7lVXweNuphmQuXNkRWLtx+iFDT
ljH5QAiEF1kvbMW1wR+gd5OnVL9Vm2gLSdekgJz4MAX1SP21vamaKI/tO6Y9wznD
XkQ2MQg4Ss0zmtxaNvtRZxCP9ymq3TUNBJ83ZWw8kQpYHfoshsLxhmkqEv9T53CW
ywMUEOZvU/UJ5pHl6nRWdKRLYVrXUUKD9ZYa3UCkd1PIspvKXhQJOzavEehJ5MRs
CFMpVG670h1bg7S/04Ku+s4R7FFBfu/8QT+dVr+Z0SCcrOn660Bx7CSgNyQ6Yd8U
0/FsFMGmwdCNWVbRIl30Yw4p5FKVJMae4/+vczXNlNYetI/eOiXFNKCnJIIdGkiS
A17IUKsz1k28Va0tqEsZCxOcX/Lg9MkxBL3Z6BqTLMOkByB5N4xIcgvsL4dy6l3l
kMR0/t2N5m4f0OI1QnFYRwUkFnmYktdbAJu9pRS9LugEcc2jN/mzs6YD05mcOsjh
4rCcNxPHYb6Labst8i0HV8L6B5vV4gNl364eb+nTsJF3KGSL/g2l3l+kn9juAx08
+upuBXpoaQFFftiO/J+n5FTIgqkH+qkacSB+cXqpTr+d6Cvs3X4Hq/qG2EmLy/xU
KvTMm5b7v7I9Qzckh45Yb97wQS6zXmKsIjd44KlmNKzAafbeSunGPoef1O5pI/Ly
HVwGy9x+cv/eMzXywvQULbvwwGXpESuyRN/tp0sJvFjV+l6KNwVdNXlHsdLrjRoe
T8myRph9Z9DXflLqa8vVs61pUC1nCPlL5fBCTiNn6fdTXbEmzVQI75sGiCkh9Ej7
78uYDz/ona8THeiUW8ITO3ocADg1nT0QXVqXNgJCWUXW/HIC7HARKAjtbzOy60PM
8PmlyOgQjSonMaPwHjTAoSzGsNmn6CVZrzX946zbPgLG+yE7h9SU+vjoxpK6wuj5
8wyr/QeefsjYIDjXtR2vQmMvzN7o+JG2sVYJ57JmYU8cesJ8WB5roHFJqxJJsHtG
moOQAFQ0g3w7ZIs6uwq1wfUp4WkdiL3ndgr/EujhAy1BDqkstkwawuKRBvjlzqxA
LM74gnFd/24nMZ7J3DzSUClCmjfcOhrFCEpVocAIxKGJHUY4FzLMwdDEYf49tMe9
3+ZoSaxExWLqvYCYskTpPsVynpwRp7KgQm/76jJJ4FfcqMuVpa/bYP3lrv6t2xBv
PWcYd8fk0BMZIEFUHNXZbD67iSTi1+vNX5zf8OeR/riQvlCixdlSnyn4iekcAOEH
x5fV8woMjV5arAbhHzxB8qStWpNitUFM6xFzCu/+SQ9oEtRlj0FS4W0VgLGrx8M3
+7HigZ0NHtDYcFVTGmmcmd0bDKnORxw+jPK15GCJctoLtNCdRdZtlCm5GIz46BFM
zF/DQm0Ow8Q3h5Lxj8lm592aW+wPTSztTgJ4hjdJiJr2yrH1m4kKY9EuLPPAuejp
Z9nrvjfaN7Dwdxw65lZyRFZxxQRbjAptvECOrzg0GQhOFuqsQzNwyrJK/g/unmr+
ILsra1diN+zIzmNMIuLpkizc5+rY2IDyU2an0g/+1ijDKapDsWgVfF1AGUTTQX7V
9v94sfIjzXsUgOB9v/ypkDlT2+zbgWRzTMKgjsTbAepU1R8Z2TmpQMgbGbSdOCZH
3CRMXCNF5Uw+2ENLlLE9Uk1Pi5gybYjXvetZEOQwaMw6l5tCKVOIjP/xX3VbmlM+
kgR6qkvilU79yfBXKQ4+hwNq82/C7bRnPh+LKGF+oE0X5fZmI7uy2xG0Atwz0t4z
rY5cDez6hP0dezA9bBBOyEQGPFM1AovpIKtvg25Kseq2Rx+k1uG7gFmNFCLdb3mE
gCjbgMvAr8L6Qxytv+Prr68shpShWtV2+xzSoRQoN8VEd8fdFF138hwbbqWRzzdT
GllSsLY+6CnWmbSeab1lUdfLhM7OmizWh5/3Mj4hI+T1Q8wvD94fAb2HyIUIs1tz
D2MBVexkfnavkQa+3IhgRNv1PX4q7qQSz0vhKfKJZtbqA/LiAuDZL2CGhidZNLHa
YgeDWf5+YSDCDSQm5XTxJuU78/U1OmvPxsHv5RccNn21uj3CFbRwtrepoNXPylcv
NDMA3tF5A6fn2u1OUcq6z4jFpV/kYSBgR3yWfLxzlYoBB9jg+KOJrsvVEf5NITtS
AZGGUxe9LdHk7NMfiUsJALp1tAHOSeHMOrvfCK5Rg1WmTo7CwvjDrBJ9QHvG25/O
T1cktvQSSN1Z4/spKYF+72g3p7vkz/k6Wtp+kiqFeAh85f35xfScaiRVtKpUm5k+
eDjA0UFjG5jaYK2PMzeH/Jj+Osf5iA0IUoAvpNRqQ7ZO1mfvV/SQAiEmqF19l8C/
x1ICMivx+QH2ezZPvoYFUrVGE6DtZ4KabHQA2dWifM0jcC1cP6HkV3Gfa9jZ/ug8
gV4sIb7m+AwaQGNgaqDFu48O2aD/rXa9qSN/X7CQQdo/tOFI7q/IayMi/Ii9yYnJ
9V/ll23UEFbK/zZ08XTwbdDiJtMPwLO017iOG3ftOaz3V76HAr/6dxCpCBxuN5OB
USVJCJT3KIlVJLmzZgV5H/PCOh0j6nsx/EvBY3Jbo/mP0XBavIQtFQirOYfxtM/G
abGnZv9fVdocXAelf7xYkauqLoLaR9fpMI8W0zKi0BCaGc+lM5lB0ZUgGIXdG5Ar
GWP+PAoNbSePhJyYvM69zUlFFL1YB74ec1gYYJiM+zLkXu688ieiPAZil27Kqv3O
Vt1Qjy9BTIHXSX1DC7tmit0o389lYm4e6eo08rjgQIwbVphvU0kTHoWNjQ0tRnbh
YosWw7tXKAmcQLktlKHVbfvv2k8LqPQ00aAp+DiI8mqoRyIQpj5iAMDb+D4g6Br1
8jT85XyU+8FIcoqqtHiopW8+nNjWZL4jVxFl79ZUGohuEvqUkPBCaKVc3o4ee1Cx
Dk6nKDkpSnMXoJ/NE4+EsLLXNQx84K8FYn9j6p+G4Q5FAPcFZH49hTxKxsGDCkfH
A9NyPra96ioZZcVvKdhMD4UjxReOPH1XGh1r0SZlEGSs1Cas2IFUNeP2XV0bmpmc
DV59OvUkUTOQjtZwXxHDpsabrfTQOWUrZek93uvOdJ1KtP8C2QErSEnWeNI5JsYw
zzuXscAMPD27Zv13RAKCOqn+N/nRxnMXy3uOnwogc/Q4cNiPDFuarH9YfWJdFmRe
7xziAvkqaX3hS/Vj+r3BNO+qx1yxxB1cNGAsDGYkfp491EQ5ljuW6mwH2qgbFZMC
VD4nMf9qmGPhyw8LHWBx+u2tMEyA7YAAqoM9shzYLdBrj+L8TU2foof9SWsZyLO6
OpOHde3Jf4r0OaC08j1Kw7QyiOMSvTK9w1z46Xv0bt8WWAiL1tDxcFREyyCwouGt
cG7TkzOYDph+5f/SUNQooxZC3v6CzHoHEqFp79/PKHsyc82zs4RJWMayVG5bZm9X
7T5GvBxWj+4fNCJSkAjxQEYFvbQhpSgMuII6rfbxLbh4PlVMYwI3+g/VpngOJTfo
skrJRqdkhqJy0aZCwxM/Q2PQmwQiXI2ICh6lhsjHHaP9e4TAwlWd8hqHDoi3/aHj
Qn+GIKiCg/7J2DzgttWC9SzUu/IHEJ5B/c5xyxRiJ8S9jAPWqiCoDwhvsGbrNos3
qDYPTkAZakNi81bLE+u2ie0em843q3AAzhjB2oFye+19iFm3gIqu+YQSJHBf7SeI
i/Wbxb7MeczkLTELIgoI3a0fQO7qsFp/cK5oQlpbT+BkfUvEgM54u9Wzqzcj6Gj+
ov3qdUJbMDXM4qH8Y9ndwQKxmNLQZ3kLKSDVFCeIdIGK+jTSUABdcNIDUf0IWeIo
zrjefhAQpOWq3yCXWJHLcM4W21dRNtT9nw8kBaTd+rAWsDyIGEyvycjfH5h5+4W6
Uw9QI87MAVC7SO4FrQMd1+KTG/F5U1zv9kDLWzerfoafjxe6dfq6DAx8exE7Gsvp
RhUVQF7kAzk4IyX8s7PCR6DfNeogXXiJZWd8FefNP35Y4Y5UwJkqhCwdn96pRdl/
Y/D5g0f4vO5ITacQtHOqwQNx3NHNdeht9QDhQjOx4XJ5G9qLvZenkm4zEunakC1M
DnCTNIComp0xD3W2O4DugSGe6FWqQWzvafF/4gkcwL9oTnW/JcR8Q8Ajz079d3MZ
xB7TS1cU5f9oyPNi9m+IEIVN6KzaPehCDYssvhrgruMzgmj3yGYMgCba3OkEOnJ0
Yz0l1u2KyBfw8k7hp9S/mQToB7AQ7CNF7ksEtkT42rQkgfoS2352WAEekAzMN4T+
4H+n7RQ52X1m2uAii2Lbj/r7p3lu0y1dQd6uDZTu77Ah7rc+3dRKN9L9DLoXHb57
z0if9+yuzn8mnGO8Y1+Gw1gXVGdyqhc7FoXzIee/N3379mRrzYvjgfY73JONKCYg
ntPZ1KbgFiw0S84uBm/upRwBUGeqhYMt6mJarm9POdgZxVHQgH07bgL1LO/G/72X
uSKKUtP3aMcQxxr0DQillDNnOXyrC4R0mEcKpH2XN5gP3ym+YatmOZKYzspTUTs+
oR/At8H06Xma7Tyv342B49PdNh0aOx0WBMJA4N/Gh2s5qF8qnPMySmrnV4srk743
dumlmhxgoYr7ZkEmoJsMkKT32GIOeKwwF2IGzAwBqPUQESYOlcbt0QTyWqekALj6
+jIwFdurvBJ6x+VuYv0PMjqOhWjz69fWf01GclBZXcHQPuFBvhFPpaDANWCnYrom
DA+bFYMV09MZ1obS2KC2DXtgDJHac44xLKOYYp1dgDRz7LD0RP5xkfSBnKIiJmcm
9cx6dgkWS0IebGTg7wBZOWbqyCOmaCa+zQFBKWAJqzuvzZPZ5ZE+LBvp7iV4sEdz
it+ZrZUT8bElfoX6UkWA8d0FWc2s7PbAasXW3yPsocFV1FUhDBL2p4Tm68NpqMl6
v4Et5VoSSHmAMw0xN7Nq1hVnOmH8Ecck4cLslAgGnL07uwwWNjhTEbl1g645GpJ4
j7OrgexhdpCRwsEQRdwK/TM4Py7DJUD80gE3d4sdet4jjG2kehZmI1wTiN65dS+2
FMzNvYs7XC4uRdtvaYqq6jNr8mqMBxgZbaSB4cflvxSjCDgpgheDYPa3cyUM2zk3
c0spvLFDPZb9iADe0/iUPTKVOlAU8bpZDagunWdmjeTXs1L7GWFEPdQHP1RqDxIJ
If1oK/EPHJfPGZLqz4Mo0PIRRqD3yWfPQscPmoZoyEX6QJSSCvsJG7qD46Ae9Hja
qj7cNHZf2BBGu/64ue/qpgO2zrYjmAXRRjpRAo+7aqogkgRi7L/cTbEmoJOFwqII
JwxtdDlIXJjxRZyDFR/97ltyFkRB66YFEncK53Ls4ych+a1ecLfC5u45p5rOdUvd
FXi8/5T8y8RH9903RdjVu00R6Kb+kITUkiugxE/AZsT0K2E+MmTHZuijpACSXgwe
VBbRccZ02QsSW52CBiRrXMtBu61QNSd5t4QCQ4Qce3R4oEeHFK+P/+rxEUqjL2Q8
gooZTaAyyeO5ikL62OD7f6UiNJX0UxvEIbLPIK9cweDs7LhymWsSIZjBOi6JLEfK
7CtExR0vPwbogV4dKuo8HHji73X2hdZr5pz8IT4YUIM5O+aUD/zaL+SKQsG19fow
gJVFwF2TWPxnCo6c6JS5cTATpPdDquVNtdkmOnwQpo2kbttGLSb3lBD3ehB3urfe
lvvdA82NHLsnN+qoNv9+IM90Y17km9Zh9l8FqRi+pnvbus9XIApXjsKP3n036jZ8
RtuR3+NotIqgxC90Hk6D+y6nXVhCwqotiHr+eRsSovz26D9sPCbuGBPO/fwM2cBD
hp4UfTR1mQf8UqMQKra+a+zm9HMLRGgodO3D0aAGPlc5qCzaGEAQ973/JHfGUh6r
/vZlISpqOSXmBujgvFIzxu7NVm5w+ubslZqzBKQCa56Yqfn7oovgZAHwNbecVCE7
fxYsgCyqNTmuGj7qNBtv4mGCgYlSnw3Zpf0wM7PSaccVJ5NsBP4hqjO1hqWgH2qH
MZb/ePpqjV+cd0APZ+57S3kzLbeKUCxRyYOM2Kg2oCOiHm80KJd2r3l2sUEayHYY
1SJXDRtTKNx66rs85VLX0/1Egy/dHDu28IHIzDYpUjKXKLt0+AmNN/lGTmr/kKED
JoeDvjwHIzKOTHIeoY+Kw2hYArmWa79L7gYVDSBpobulBxSQsRABRxzo6gyQEM/k
8S7jYB7CnQtGav+nmrydXUD8JUfBB+I+9lozZB2F+cflRaHVtK2k20fSmFZTxPEV
U2s18gaG65InY70HggNN5ou7lVjvkKpcsNQJc9ECdhf4c61h78AaRj3OUWUNwZbV
PZXG2C2g/fXRrvLMDbwLXhAl4i1lrtoR0t0eaKHXH0/bOGFgc4lBFRvhu5yXsvBe
TFF9adc/CeY7sUyTX6q7gitGQwCZhaAaDqB3wV8TP/pgPdq5QXVw6ScvH8JfLbuI
0Tf80+fuqXMlTsU24gR9XrwK9qpJGYcoyzMgveNF+Mi6x0delNKJkX7mKhzU7iXn
kqQum+w4l6uDPptWQbrD+rh8NxZH22TMK2+Oh6KY+TBw6w5/MhNJm3CPZMMHOSof
EXsl8Pg5xyHheSUcHKqMIF6hmbP6ztKYhSs97HNNnaKsek9wjThrxHXo/Swo4W5P
3O9d+pBus7cLPKPnkIOL6f8G2M41WsxbaLDaQVZMvWiWDj9G+LTBMrds+SJTTFB8
uAGn5gUevJsh9am/a4ixJykKctk5gO/YSDEyOJCuRrIdGI03gEZMMtiawGxVOj33
mkpTWcgepSXzq+5uuKHHSQbb9V0BKXWSX1Tk+QxzqWLnhm8H3fVQInkMVMl7QolQ
DIzN6bSEWYglyCQXH0GyP0ALskL1r76j0XYKJMIWy2vXqeqN1SnGDhoXNy1phtpv
1Lm3QEmDmUaXO6czf1NYm1BlBcMCTrUukuezdICxATtCtCBW0c4maasPlXZCPvuO
Hmz/khClVxWTYt+BMLVw+d5oZ0tFXcJG8h2INj9Fdh9UzOqSaECr+EyEhLc8BCZe
at35GRfiQLHCf94Z6DfQ5talyqr3cOV+tbqFXem9pu/sQaLLrsMvg9yt903os8dl
L8Y9Kh8WbliK4dCr+GzJj0xXKgCrgbT0xIK1rWQ/Qfp/tXSUjyVG6t98eUFZNFWb
RYYmoxg9byyQ5NTdlheutjuYUAKKCMOQPB2h16IowDz3b2vkzGtP2PJ8os1pz/g5
OukTQM+7EmE63pNFmAmFO0mDUlVd7MlUCFeOUYxzyis9RIznLAsgNA8FAI8YG9Py
tSpGSVp51YmPogh6TvzyJ3xa0plHes4URld5NPSrYO1Ci3JEOqC5oVw4vo35FWv6
8cyeAE932TG0aS0naI+FX7eoum+ttrjRoatxZxQRckjEKmGXzn0OqU1heVPYTzIH
VBJCsi91+xrktMa3j/8vkX5Z5RDDtGaE8nWklgkTiaWYYbisRGa6uXeiWVbFVHyZ
VnYddnbrYVIKXwcHy7eyff02FD4o81jmz5tdmsMrJiOX7xoDoxB14IC/okG4DN2X
oWYPHNSJRLFdAlRecmm6oyUdLW2oJJ8KekUa/FAYgRK5EHF9ik9aXhTaojbYBMWX
23xqFqqtRcOXN3RlnVUpCx3gwMfMKlgfYoCDTlmuSUEWkucWb/rHXUqvvB+SKrlp
Hb3KBozuE5dbPbeMcAS6FefQnte+lZkTfGcDIF+g6UWbkRc56LOBwlZb0rJvg/o4
06malgyAkcTWc4idjWFL9+5+L8qP+bwT7WMh6w+5UwR7A+Ds8Bla4sjQA9kW+Hhc
DbzuxY5CKarse/5nETLTw+Ida79H75BWfPbaMPXtqEwufzRCsk8cMM9/tmD5l2/x
pv2Qku9eVVWTZfp7LF26pctLUTA6Dbpv25JtRIByNvR1JbMn5TJt7EcJMczA4W6g
2CA0eBfo+C8en3MdZxOFVOnm02aqRKy9axZ7hP6TmQh7VWeeqm+wyclpCuqWsiOS
4tYkAduYkyod7MmP/cx7ueWsZ2pp2JZdzg6VS6fRgh1degg7/tFrS6nX/dfBEV98
sR/RkL7zR7atjlQtafSngnNMx2pJG5DLrb3e2yHZ7XrutYaB4SHt+RxWupCP02QU
jyGzZjAokgq0HotCn8nbt3Jtk8yBHz/0HLHJjea7ZiSJUS+vcBnwiz9bqLYYIbPJ
7eH4yjK02zYdIb0W0AmGwO9kVSzwjtel9TwQagE7PnbqJALOmIWrfEOAHqfSFf3k
roe867Xhap2wKZE6ZX60R7ZKVoUvwyZ60s5TfKKXyUskNfFMhmhoe6NUbjLBC5fb
VHbKA/yjCd/RFmDBbF0uf6rrP2WKVSZW8KX80VItb8zKmLOJbtQhKqqmHG/HK3Iy
2ZU3aciPt6n++ThylhVJSfHT2DdUNy8OUen5crIFY9SYLhioANIZQuy4QqKsjqF2
oTsnjWzfm9+X3zvLUDOYZvrur1Unvn/5zVXU/GO6JfRItpV0X0TBCu/3ewlfWPMD
1JKPW1Mmf3Qe9OlW0zuWlNIgpkUISv525/Bjm06qVuH++cvLUHFkRRQWDUd0GE88
Ucpi2k02yvek0ZMh6v7lWB4gzESF3jFM31EPadUg9MmT+Vyel/rS7WrOLY8fHyWB
r8LGvnmzPZztzF9gTD5gKPEMkLIIDDaK4FjIjSJN9fNoohqKa9Y51uEUXRuUalYg
w+QRx8gN6CoibcMc6yrb2B+zSPMSbsHLDp88WkS3tR42x3hxjIDqH1kiNp7Nptu6
wA08Lz+CUqFcXirMe4zSdQy04Xl3rI902nQm5IbWNRfCQAW9IDonCVzlZOJ1vbKJ
C7kNIbk5pAVuGPMmycaBfXSsdwyajJHrjHSPI6Bl2n+o2bMpehjLEzCtSQvxUcOR
bxQSU8JgJ4DIIX6woeZh0DVwSDGcwwd8EfT9r2NpLiCy8aRydfwSM65KJEGo+Fln
vA8U33cnTJA9gXdhKl/Qqo04SOeqTQYQbrtGcDy+dHM4n8mOWext1JdYUyifuNjL
aHAe3bxAdah+gkLwlUJwczsbFPsgY/S5jfgg3wltpj4lkOc4+/bWaIXyzkkxYAXB
ekcMHBZldgoCqW1UwkktIgeWOteNvsn1CLfAG2vw4TyqJSL9dnl5wGxLD8KiuRoa
Zm8vu2V89c/GTFlAIZiqZTk1LiCq0PC7knVU670bBFqADWwVetI/pBdv2R3aZjy5
G/aRd+BZ/ngkRdvcl+nR9h9faZIVllj6hVlEUJ+C7XOQJ+Ti/tY9lk8qWcV/B5p1
S1MtJVnl8L+3LGbULET4pssIoTQDNp02/hQs8S5ltlfuLmHiuKTxBkBG7LnQe8rW
yhzBXmK5QJSSwfvuZiYlpuFsUvgvdUlw76on7oTzqYZGsNkqUZQoCt/FEnhuLDIW
8uPODGWddrUqW5gcRobyCSrjZpJF++fGvG4F7Y1GyzaVkFMy9BiDmcfZyglWmLqn
sX6fzOp5KQ8EdySxdWUSiRbgfhoZrHVNsGJ29EMCD1wtmN+ANcM9bSvqP6GUL8Pa
BjoQd1Xi08jSkIIM21ZYNZ/DJwPb+iKr1s9xBhBTItGRODVomUHVdRvfm+u8SMAD
Ubve3GHYl5U8V+sZcthmAf0S/IqfhmBsCN6sQPZaxDDIBvnlzUBbzJBRmSIyyN0M
icpIyIEhclAp8Gsf55RDZRGQZwMHUU86+6KhdRGnVCwQtBpNBRkUJYfZs9ELPyWq
84a5dNpwmScNidhx9515mPXJWErJN1Yepwq4yC1KlxtjdkZx7vzCu75blGJrP2qp
0tiLvIL+hzz0FRnjnvMHjFRBVKt4JmjB/CMvDHC3K86npHi0QyjG2iMyDJQXFZPT
7066rF26pY5Z63w5BVOlK4JUFxfhAKuLqed6awUYiiKAQlFp68UD8D1DALWXzdG8
CHTTyaCxrwK5BN84Dkdq2dRzxZjPcdTFzerxiRemAt+i6YJdeStv0sCiLgR2vT30
kFII20vzJ3zGFqksmMaMTgJh2lx6D5B9KdlA57rwnvtsHu53LhO2H+T6VvF0y7dx
0VTDHcNVGFzk4mC6Uv9ZRlT8Yws7cRZ9xuPq700hHsxkIrVuUqzxI0BWrZOx1GVI
sytH3O9o2mo7SaP35F87iYfAz+G37zBXYUj8ikWNfq47ldnrVlZRvdzQnnQS9MYZ
FtqwHHDe1/WCRNuwyTT7OEDRLV/09AE6CGj6JBMabhx7r8s3RdOC+ratFvInxVWK
4vFwU0xb7WZz/HbvQPk+3ede7CVgGHndlZn4dYIWZHS2cvMIUQX9ik/JCOHeRSQ/
stUMlw1g2QvAoxp68QxN8HAWj579zQ2w1rQo+Sgqk7CzB2aiHilH6gR4yd6TQbQI
9YDojaMpWMte+3Hsgj7oCcK37TfnCdho4lcieb91ColHHoFLTn3Q1iiRaYE8TsWq
GeoyIcrKYPd2rdfnqk5b9A2H5Ee/3D5hHviEKqNgTNL8sDBIDGUDPRy1WNPRh9as
xSv55Rh0zaBq6wG8HDQOTWAbiWZpvYhI0/ly6HW2xqUP0nDpWMBFnkSivN8b2EIx
J7m/xrBF/xWSBMgYrWig358YJJ6K/GVcGri4mTDJApHeTxEzFbL5QhOBoI9f5hje
ocXZ0qbetzh54zJ+48NoieRvnRo8lGdwC2y8AztWcR0IaW2lojft9HNiax8ldW5y
VLa/1w36mn/v6kRXvJRfVJfTpiDn8a5AonPhN/nXvF1bCyBj80EQJFFW+gl2bui8
OYE++fCWnBXt5bH910JDrhPXNGWU31N5WLu6G+zAAKHz51ZbcUcraaPE6rpFok92
pdkMXBpLekrZG9gxYQHRjMaPo9KCEOfqB+tCegFhEwhgfXrwSV9G+bEypURgYuiX
SuvByJwgVK3wmjnW2xy0Wkf6Cq+CNg5LEK7miFG3eyM97UDo7ZS6+i0B0D+tTDQj
2A5VZaoyZv09aXQkhmVa7PVi34t31JIiIeK7rG9h3uuAeG3XvroSGxFjjjLqcG1l
dT1PNgv1oIaKTQ6EJ0O5nHLIvAdU8hwI03UyO+Tf0KTvGGuiSLg8+5uorEMvImcS
jAuhttvYGHw9wgNBjjXkO9CRu7zhxQ3R2RO2VW8hfkfe+TWxtkhNzxAWZazBEyBm
r+Io683OoaFQw3Fr5zZPNz7EarscMkVD8pA+Pc6oRmHM4giJGxmXcIgz7i/ieC8M
nMppczMU2/M9dm0nfKL8GnJGW+mF3/ya1LpvmE0zyWLdrzVf/TEyFHi47e5FFonJ
IxcjrY8ZGrc7oAmAmY9tjCDf5mcQGrEUqwMueuJVmJXQB6KZlAkkPqpbwAIfbe2+
z+hyWaZjV7vlQI6i3O//eh9A7rfHlWM+OtA9VUO4qzFp/8d5B0zlgAPrxu4oKScw
XhR+GaXmImNcF/9n58hgy959nE4h1wQmkmSp81oBbD4PPafykUobKjhLBa3tlo2H
enKHXYv/aNodDdX8OxbJwuK6HHYO8tfW056yGkbXiqRJhr3ZltZUVRyKGK+qqwZs
b65JjFM0TlErB20kSDTzLaj62tX5zy3rEcIANKBQ6+XRWb+97SbK30FMlawAnYmU
HGPFHH1vE/YeE5x0f+RlA5zPI0ioVQ4PdlKXcdMHNS1X92NsNXI3CcD1jHAvfq0R
Q/qLB1msH9GIfUZBLfFQssYBBrzQgfG53L1ygD3Eoj2EszNGlYKO5tk1bMBdc1QC
yosv8iAEixpln0Yv/T5KPwgUNjFDzlXPfm+oxfAX3SMTZW6+P7tN62ki2oK/XBcf
XcujTL9rDF1NOc0wIiCSsU+DD6tRf8eE3ANgE2ALP0O9KSMEXaIzm0osahiaEYf0
/5KASoiY9AJU4a+GaJA7fTTLsxN6e3Gua5sa90lBLYwHR9oFo4sUJSqDKfFXwDCb
pfJW6S+lmtlVxOnesNQKrM8H73ish2Dj5HNrNoJPfVDuwPkdIIIoPc+mAxv67Nsv
SienC0c3V7pB0h5qqZDl+tYFixHQe0c/RuFJr2vCbA10HALzrWu25ZfwTnDkcZ3h
AZVcTEe0DPkkUxxvmXjBzAe8K7G0VEPhmvwmiSbHvDxQe78emxv+BOY7KoCPpyNR
x2V5ijlrqDhTO6dSz+V0a+u2qiNkoej1Eoy3hXhbkrF3TgiG0vqJIFxKgNyYqH+y
SRorZJAt06I+dJ0gAbbbR6g22in61vrxIwItD+p49/+gELoxVfLEHZgIdtZ2wWyR
rTCSw42CmU9r3pILKqwPZWNCT6/Gkv9q5stTamUjIfh3cYrm9avZh+xDbIuDTf7w
v5jzG1DOjpdRUPQN1tOaxLHsTOuomdvyCEGnXvA/uN0PjrHt3KgFFpJnOk6tTpgZ
5vxkBNJiRDww5VR3aFrOeiZhGM/7JXAgg+npbSYVxRtPBFN+jvhxxI5Kbs4VzfvX
KiNMuNvr2RFADj3380B0rKQx67SKe96dSIs/Z2qgeunPt+ufl9WPzxAlKT7OSnJ4
gjfCQTtJySnppqwj81QlZ0TMlHK6MSVi54Sp+Bufw8SsC58otWFJI8QUiBGr8X/b
ngYwXw7ZJSlx4XRUbFdU5oCNGGjndoVEspG12Xhhp50iBUrOd4LJE6EZA38Q6XJx
uKrlQW3OSnY/7KjdFV2qwA+A6UO+05WoQuBLo+w2iQqP5zsQwRUOEKn05SxVdUSV
WZMPFWPG8ObjYFrJjJzqGos/lK3cBalOhsHxfkovG6FQT9Nd7nAmu7eGszNItO6X
r4Wa9Y05cIWcaCfWsqYrSyimGRo1pwESAlZIOq248CypI1Y99Kd0cO7FxyHfBCwq
d3FucGc8ILf3FF+GJeqJ+mJBZU3+n+smJGJD5tRNI3/GIX93Uxpx/NZFAOxr80RJ
K/G0xW/yoLanRfOwuwvQw2EuSizhk9GQ54ZnmV/PitR5UfM2sVZAu9QVoPh7Egk1
XbDo7ic4U0EfY+uOMT/PLckzA6lE//jcGyc5xyTvm5wZbxyLE7EJl3e51mqLLdqz
zxd0e0NMe4Ki71OaX7Cqskp6XwX3AsIwHlkHvrjOu5CUcmx3vDCMastFrHeydmXU
Y/LswpVluX5HuXxRoPGoL3HnVLKlnXgvfQLwbWhouCfUSMVrAo4S/TQW/crq0+89
/vvEnvV5m/WNjqlFD2qCB4KVEj1mL6ohaUUPwFpe0qqyQwW7EQDBVXEfufb8WyLN
rIEtJbNU0mCNwhyu8pxjZOowZDbjPpeSnF0++r024a1d+3E0OpJVhrTIkp0d4lm+
oA46k1BQYoe+ExstlkjkcgCkAFti/6xRAH3DN1evVCSeOfV7+HusKjkMRrlsW9sZ
DUFSx7qlTmN8kUsxWzzi7fc5GpsZhlH1GtjLaIByJ2CwWnWJjia0moOjSYVWw4Mv
NpMdZJJrmx30eFd3jHmPLJXzbJivFp+hMcqQ/Yq0PlxmVnuCQEORlaV4xRzezYk9
LyyzcqFrbsnCvO5KoWkeaPoskIH0JhDyILvF1sj+bal3f+vveUB9aK+G/DWmLo4U
Q+QqRDTPutdW69v91sfmn/Fdix4zndNqMgxi+s67HUjN4sX/vb1QbGX7SDTD3/19
6qsRQYYMPDq8WieTWPmUHaLyV8GisRPfQGn3yEaX+z6pTRz77NBD1oQ2g8R4ldXz
UDIrogN0stS/mkZG9iE+vMk3/WxmX3AfhYnGFPTqjm7wJ4kzz2Vrzey5PODyHGLs
BE6nDYIQqbC40XoDYJsh+FRoXe57+C6MwHIsN12REbaVkvz68jyxizzTR6A6Mmtc
zYWSqIdU7y8KW6HKzrUhY1ELTN8c7neql8WMrWXKmb70bNg6cKtQzbmGOWkWpfq4
Y/fmtKP2t7grmUOFZIx/keAedFUlZdWXGCSKEvFSl68+YTdwDN/A5S0DV4PBgWpj
k0WfeddyKpsTjPl/mIGTEJIQt0VAqHudJHcvUbPI1y7QTqJXjz7KS7fz0dhyJj5q
FpmcCg6omUjnq+HgLctXNLoj0sY9d/a9Y6okJrDNJBxy1QYTLJu5K94AYT8RUjS2
kla11TzZr0lXuxVJslXBUGwaUv3ouCssC1wBcFqCUuWCINDv868pNRG4oEu6T2VA
tLA2/omDzsRWXx56bXufs7AIzI5QSfXklvuaSnSR+qY3AwzYBk/RlAb2QKD2VdZF
1rC5E6lB7zQhbmp9z3NaKx6zQHNJWRXasdfDftLb0Qu9tIcRomMm7NNyyeqlp0Ld
w/wn8kNofXYHnwCNVwr+GZLqb3u+28tlcSIwJN5CNt536RuwDQJgIMJ5XJEcL/mv
b3yRztJ3/lO1ZFENS/rCU+k8GBb5njTbhacEtHAxs3M0WIplI7ko7phmQqRCGTrN
BFCgr9EW9ccUBi8pVIpAE0PN9R7dSci7kwW77rUkGfWzYLQCV+1n/6LcNl+/PxRZ
B05QqqiBLjWMeSX/SUhoJLU0ixUziKnLiMnipMnRQcVb+88CKBvPhL/6tJO2lzVG
IXZTNtKnYTTFX9F5L6bBcQvzCBtl8YLVc4cSDbE+ikCi9rXXsHztWuxsLvS6Ce9H
/JUdLqJZQGQf8q8vfrTyC+qZzylNK9GOAVEflRxAwVr2wjWg2PBxr+hL6A6iGwjR
CNVyQHtt/Wog2ZZPS3aFN1wtiM3fDFE1ab0K6pf8R+hHFeKWLO+nRteHgNw2gcP5
Oxn5wDSDlI2Ot0BhuwynDfmZF5/BrjGDW4m+pkcQ3mt8zkwviIPYfTFnEpXsK6H9
fN3zSSNkGOPWcq0uNSuhh4WmaafsJWFqfcfmw/0SKldER5WjGA2fimYiQhUQdPSx
L49xvE1NYWWl6B/ERMvHAps72stlc8/0a/zW2WtYzlepm2AUHrCa6MiYERbrlT4y
43aIElFuxCvYb4wRAV7ynWOPhOKa6VxDyyRtx7LdNHVWlbciBQJo450rEgOtCdf3
Bi8fLA2YyHvo3+pDWocOw/BuqJfdNpqAR/0f/v0XQ2yY/4xi+aiOHJK9ULTBK4Bq
EddcyKiUj2BexC1tD6URG72iLo1haCKkkGFB9TJU8u6Azi+reIjFHIPqi12HL64Q
k38+jsnZSz/ABv0e73iaBWuoyQAou7AimmemlVSTVePvnVrFrJvvHz/TNgY2YlIA
1qaMnwIOqfeD+v0cgEB9nwdexfjdX+0yM3u+tr6Yxznc+Ub+9rABxWdPbijIqxGR
CCLM9fjDyUcm3c6wlsYBK8wuQibsV3rkc20l+or8wrQwKAgGbi6aWNfBT7R5QwVj
q3pu3Ib4ARVJlkfayxO9K16PfdOVB0uWRhjxtiXtiUD7LbYMn4bxLt+Xit0u9Dmj
mu7/IKg2EVLdl/OZKnEuUfIa6bshhwbdQhnZrcOLgLafTVia/YiblDWl4LqkEMO8
qKS/A5hUWlVGPcK5XecC6XzzF2WGA4aY57W1q1rZfrKQO/HzX+9Uj0koMePk4n94
hfuM3krYl+ww2oYZ4NQP5CoQ6ybhD3I//apZ2uTV8PXMctmbqtIbvQs+sBTdkfAW
YdtEgp9ooNpG6+WGmnM7rWApTaMdrU9N6b4XVI4f5OBB7bEtiWOjewWwstdq9hFZ
oXdBokS2LJAiNqh9H+FNDWwWFLjYJ6R1d5T+EwTzR9XOgHedgPYoPoFGwaa1SEXW
q3ojOvaW5AV3zGMnwinV1c3+fs+4msrvwD2kcO8aoX2QcygDoD3qQlZIxKB34AT/
Z/ksDcbT+y6whk+2HI971gw351K/nIfIYcPDttOwvDAszlyXqvpRBl32KE8i0ZEX
ynt5Qstc23HmB+/LV4KLT8G06i/zbKnkACRRoNLViQzB2va190jOW0oKfrJ6AeJA
jvAKrP6NcHeYzUSg3gQQrBpoNOm2nxJ4uekbAEgYBc7EOVZB5xnG7izw+g3ZaZZ7
xLGRE1eXOMCIEobhsmG3PM0aKZQ8RKTqfym89uPx9B6EPGfm36PjUDZtaW5Ayflc
lJm8ALU3Tp50/o+x1FZHvKFBpJaix5nzPBeIBd7ZsfmxSVF0/ZeOAIGa1Y3rXjJu
BV/p1W7YWDHAV1qfNSvhmPtT3I1shZs+zWSdP2KNpdvAHsEOWnVs3QJQ9OErCiml
23CW7j5tf5opKcRVzySohwsdQOZs571CesgTrlqDbr1zGnFktdBZVqKsi/Eo1wBX
g0CdAORydhFblrvrfDRM6vEwrt8yRcs6p7JrMVeukx7KZX0P5CobEH8nx/g3jJk0
vomRwLeJQBTVKaVUMCkkQU8nYqY1HvqTbWH7QdDm0TP8+q/ZCU3NtnNH6N8BBzHr
O2fSN2NXyRsyZ+1+tH20O9TxqCBoMS67x9SC1ZLlOB7DDhU2zwBrcvXKUePhAyJZ
8FhiyemP8SvbC0RIUC6f0zMYs3J1YrCpIbLZyNZqAzVE54mKGBJ05pzKrf1qY1JR
H4sB56eb6wlpsy/40ClvwYAaX5yQ/5zVkIqRLQGq+Ci+g38l4zrXjIke86VyB9mv
HxNSybqfUjFut+BJOg/GE6NtEnhkbDrbDAL6jpnPohL5WaLHxqQPzBIH8IFTlZ6J
BVo9RYpVfpDPCPtpPJdyG02S3srxi5TK+z1PaTwGNcncfIl5Xs4IBVlC/mhCCC5s
oorkduXgPvjXU7njkYgHHQGOkJx5ZtAuydyRRmW5UZaVgStRO0anp+DUwsssFouu
65qlAlAMKgiUCVvr2S7YO1YfjanTbuFd5NW1R9ga0HsIb5LQd8FN+LJAICN11eQF
B6o4Ab98dfQ436KRTIxOY9RWHV3uxJmdrQZ/oyZc/iyK4YVH+DY0AFeTz7/xCqVQ
jN4Fu9EQdaimSYp56EheYiTmnT5t4JxIsO+4E/M7jUnsNhaQ6C+w6BMWGHPwK4OB
w9vUdoGnHdIBOnKOvVZKlrp3GuSnx4DuDy9Fvmf5v9Jy4Fskojb8ctq0NjGtXXeB
WV4NVIvXVRAGHEh7/v67ihewGdYBiJ/4w9vg3dLWK/ktk3WdFeJhiiFzuqdRAulS
nCiFXyweQeYLBcwVk2t4DEx8DofNmhUAf9K0nHmT1suE+Nf9Konzl1yv/WpUp3pG
MrHizAgfmGhy1qlEX2ncu+cYnu6uK04pBHpzcyks8Qgnz7BkJZtsEYrsvELLMLd1
fBByV1E+9JzNjn2bgkxaLDJYJAdFnmjORjjiF7ZhFhxelMJiGDEESI1En60swz+2
xaio4UIDv5EjLul/EsRJ5zr06vGamiRo7vy6Oncig+dZP10h/lo65w8qpyjkRXRo
ewh2EM08p8pvtskTayFHQ9AzgQ6o2Lvcb8aE8mSRtw9BjgCF8UDujhK7TwVy8g+s
X0l4dGx1TDrB5K49ysXCoMoxkzx8tpQLSsqpDmK/JnrotkK4/kzfJyczzUzmBgmm
g7ZTwkDKR0PoK2AVwomx+pMDBphlthCWhrXY+vUWy6aAZSu61X3fZlLnneYe2UHL
pTCNXrA1UAaoXql8xDO4ySkAGPwhO+gzjJJUbymm3OCFY6KQfNDZ9geo6znYjCU9
RfIU9LR7o1dgkOCbmvxIMcdFeo+GSOn4VwtZnZj/as38ZqseHNam4HasTo/+Ugqs
iG9DlIe7jss1RDBys3FSRaxq/3JkVxBR3Hr/AfmZCLASw93J2p676BC8sXclxf/T
Z1QgB0WpQGo/JSKYjwzjUtn5KRlT1fRGQqZ2WNU2NZheNFxdNp1/N4Y14v0qVTc3
AxXT5ON9PMTchWKy9ewA2dpL+3X8UJmTTXup2dFO7VYMuvZaR3xtsWHyE3yqKO3O
wULe3rH27Ehr09ppjz1D2zjL99oijUo7RenXqbCMuR7KEwZKmTPGS0eCJzC59R92
KXLSU57oVu0x5W4+ndcnrVahxgt+YPlgyaL4JuyOSkX1iUrdabwOLoN2Wyx4LlK5
xMCtrwsnk1JULsRHZoLkaE0k2q0ECAoeVI88o2oCNL+2YUXK2WWdE2y2Twqjss6F
8b6UWeuuCIqlhUiFcKLSMSrVfwRNw09yYglCJy7AzhOpc6/7C3sSOoSPgM0rSEF0
gUGhQSa6fry1GMfRk5sCZRLJ4pK0wnrLuGjMmwKJ98OaKz0i8wN9v+U0H2S2oTZ1
3zKDK9Ba3oR4JmBSzHRpt5MJ2PZ9MdmGpq48+14BOXKhaYu6CtMNyisgK40TuLNa
piGWtWUD6/UsCD25KDYQE3Sj59pEfx5bkWkXzptXj+uuh9N11bQbCLgd94oXFe2c
lq+dNKEaFF0zHaa4inqHEqWgy5gafQwhJH9xqD0rCq4Ck9G3k4BpA9sulRwLZzCK
WlErgRXh9tIQAmIXMmg6gqq0zgNiV+n5nLYBs1xxMh0cvFmbQfuvs5OVIbtsQAs0
MlWfc8+l3HW2Skkb8j3CzOhhIXaMrwDAW/4CyG4+IS1Wbc0g1OnVbXQ4+Ul4UMRk
J5dT8BdN3wqCUzokMxIzuRotlZiPPUy56DHFdICVOD1BQNyUT1tlQ4XgJiOMqHy/
qT+8eU7dSlz3G2/SJILH+Cd4IU8pq0gegw/C4BbUr4bz43v0sqPgobwxE78Z4ZYR
oMII+wMY28/TR684kq8KX9vjIni6k5jvXVzejzEkJR1siD0S5PDeNJMWzSuIInkx
bSQZPI9+VcMiiWiKmcMqtr+catRR6kDn+FECSZ/VqjVMu4qGHKbp/U+0xNQpPtp4
jj9itswQ1r5yYXgkNOXXmm4O8wqd+nPZLVs/HarvAKt2g/nK0nCIp8xJVFivY1/c
6cEpMrpxlDYW8Oebk88QZ8G3mQKGsvHI+OJDionQeo39oscpfGzVryPEN3RmnX99
RW4jftzLDT+wxlNzZ0Urg5CFhPRRTKXrdQlcnyOK1429bfShEfJtlss6u8dgM8IB
AjG2igU4+rNY4cX2b6Y/RBt+qswkASQdklk9WV2pgHtvzplq6cjLlNQqJ8440RpM
CIeIYap1HDgc289ng8X5KM43HXgoO+QhkDCyf7+RG5Jbkzk/nnhR9jZd7Q1PjYKs
ScCkudtG/E0w+5/fGeLU/skA42MASRDxhE0RH9AwA+BKIGBVEA9ucQlp+vJghptB
FWVvGRv2K4eyriwOsUL7hdyiTOQB03G6OYr+raQEmm6igDli9lVltoWIuiJ5k/qP
e9pGgmsFRusJCSX37BRmWuZxcVS/0QPcfuleiTzIEkG/aGjYpNgrAR6L8yp9NKLt
ieUgz+FFS1yNb8qZJOBicr35e0qTnIFh5Qt7sZbfvqcv5zpVOtHMfMGKziFscWpS
BvQKE0duHiZa1Y54U3zsKkjCtwtS+Y6uxgJSLc4u6Eb/RPVV9RtCLvYnVWFgQ0n8
o9YWsfJz1nrRqkOb3c3VwGDgiZz/1nkhoAFnZamPZokHIJzAJFVNjPFv2BBb30Fq
lbv5oAYrOOZVxxG9yhFxoxYMJCeU988lo5/20sN08iYWbRPw1n6qaz0CyaNFOZfk
L833g0dBktikJrX8xwiPd6lrGw50lw75qFMxYEIG92onu3cLzGP9rBku4ljT+nvj
IPf8c+K5nsE/XVfZhL6BlAjc7YIFfH1dyCTt8TrP81hi/3SGx4Z2oFIHUwg3A6RH
2RE/w0Cc600PizS7BKOdWwamkIL+PU+07TuVKYhbKd2Dj8/8yiclqQcaRSZF+cCJ
dGltQczn3tanllKJ9MJy7/h0coTR/QkL+Ds9q9CER6/XWvqP1BEqdpvWReLESzU3
s8EXdpI8tG36iTZ/Fim+PmBAgpr5gRKWtlVi8zBJA/yyUlnMvGMhElp1oX6asZeE
Ib4NZtE7BTWVjH2otN0bpLgHFEvCs75ps30/rVEbtK2Jt1eRuOt54isNvgr6FtXk
ydhkBr3A0zplijK75ot2IZI9H/osZ0/P5pLOftO/OzqVCwzWfY9O7Uko3/EN9QM8
HaSI2IQJ5B+1pTYn5wIFVZFOBO6pXs2pXXh0rRhbwUxqfM4fvsZndpy/tIEjNvsN
hivfEVjl9up4uGj3vMAVLUP2ygiNWtUOSmYDDvd3zvHLTfLChUrb4/B29qyg2qLw
hQwoGABjGn51CJcThUBn02pcf4jSKdGS2aGnEZFUKZ7aNqfZDTBzY12BU7N1ILfx
BfrVgD3GkeISr1gJMipgMuMvRP9pTPBl0Fj0Tqlkh7UviYTGedpL6pMDgfiitDcX
K6Rv/7Dayn1fkD4JS6TUAiVxUYOf48dYPNA7MSxRV+mmVr4MOdJmnNyklVQg70mb
9olrogxTBLOmQGfu7kwsUJJRWbD1J0y7IzBU5p2t3YySVllOOuQmyCLxvWaVLmwL
5Rsf/Wzk1706KbIa82rtN/yLU80slPmcDV8OKViCk5Jd79Usqg5EOmaWS7jBRSbD
q90se6Fbr27n4p3JG+jA+49XHnsbEEwSXZj1pADR+la9nPoDXhGSA3/kgUybMn1Y
Hy6UouNfdLjiLG/jkHBxS+xed1K+ICl5thHR39dsnWJb6ewnsVXo4DMvBTBHtKPw
wY0ieumrtDx1en+pjdTgZrfuAVtOZXDNi+LYCzFwZi/tebTy+/lbShpT8AMde25u
nUql6/wzJBU49Szbmg3JzHYn2Sdqi1BmnFw8obTGDcoxMQpXhSYR8ZhePIrZsLrQ
o8eYFC3o2UDQJi6klq1r2OjO5bR1tgzISEOIDHGzhW3IwjUJh1ZgqjbwfEFfS+gE
0WZHOZq+qLWhcI3WW4S7q/iPvKDIOhpmT540An04hWkZOmoILj8A/c58jBxtU+Ho
Yp+A7310pj5iY9l3+rkSWgRbLVUqRAhYDBHlqEL5IFbmClk/RaymDE/55xEYFrCs
1nxnNVtX0jv2nAzIGYa1mGVXEVopEwAWxEI4F5pNrcSW/JHyN4HsO4cQwlufI5J6
cnTofzRbiFMioGu4OxDk4yTESBfRhlU+LsbPk7NtGWEQEmKbzbqntZEQbphWwQQJ
gyQnlq+vadr98v5lgPpbSM+Nkd5eR21A3HYGk3ZzoU7CWLukTLuCz2trpEYmLOfj
WnmYbSwLmu12IRKeOBxKkvcXUwdGD9i+Bdp7o07n13DxBpIk6JW5/wC3htUH4rrF
fmOrdXRQN+kNUrMrBmIHx67LGNNd4M5NcVXHKCnrxcBr/QI4EaqtH6EAJPKTvQDT
zvD8oZgg9J5eNkin14aJI/hQFHJ5FRp+80R+xExJqwb4RyHRPkiwUfIDwRdfEm8W
rxWAH74Qpn8kKVqJ/M2VfCPlK1PeKFweVVKQ8PhbgBJNROogL2VHbhQrRXjPt7++
WtSFGY0L9zWMxnpqUIQErVZY0A5k0o2sucdLzPuybNqumDsdV/XBqR8KMrcpmcbg
Yes3zAPmNrDUFGAZ1zG+ieYIkWcPKUtu6DjkfB/kCUOGEfgKX+MOUFdnK1qGqU4o
y06ONWU+s6PB2vr83MjQtSHqBSPC+e8U+jOStPFuJ4xvkeWeq0kc5X1DQlZA/rgx
Ym26Mv7PsqCtcMRkSDdF+p3kowBzq6Pmej+uDC8eJ5RuRoqRTAyQ994n+bmLLtcx
IuUsA44Z+vTUvE2CxAVnb2wqUi3MAypVusNtxN3T0Xt7y+bk9KsQL52SocF4bT2i
02cIfDMLiB7MAIZ1Zoe2aK0/4tlVdcwBBBU63uurOSyqkviiLKIs5MGXv5QUj/Rk
SjWGCIdSxzG8CR1uOGVKGiXyK8l6wci13z7RHiDBS+ehIj2vr5gFhaSqTe79vwS9
gUfKo0szFJ3HEiGUvS9aEVVduxz6+d04IUEQOmwtyvT2mggkTA82lL/pxgizgbgO
32dI6siI3/c91hY1dKK75BXLbOeZz1Afu6QfM+UoEjRt1oNrcpR7poPqes/eES56
hkCabIpjE0I3T4AtenO5IgO/8/aDRxH3N3HUZyihqUwlA61pPkan0L/EmbFY9uiQ
YJNyZ7aC1nEUI9alGZH60s+unJXjNQo8mxl6QDQin0m1w2iRVMZ9+VoM0tLBAddc
aE0+9qX0x9Ce8gJm0UI6c/Eq1WKOGvgdA4MgL7ENHmb3NxTYZZr3/5LjG12lL5RW
obsgJ9SLaMRLNU5zEdhiwAJ2j1PZqIVabkcwfvMqJpd8RFl3LkAITarzT783jmI2
sw6aLc4+4W7icAzOdPD1UYpMyNBqVyXJCGNlE++n8m5niKdHh16Mf+R54quTeq6E
ANFvVJB/2XyjOKkLqG22KESWPasb8R4VuSTCWp7HcBHfbkvFTvxgl39uRSfTwXeN
ojRT1x/roxW+MTCRlf89K98Y78vrH6azG1s09g/HTOUHy7VD9F7d6uxwfO8IR9Co
/fniXZxsBkMLNm2byhrJdlIKUEKZ+jbJI8smrJH8DIqCU1sG5j/A7b3roLk9l1V4
WhajCtOh6udQ+efqrQNlfig4kHVV10yYdaO0yOWgUWps5w22nhwEvjhMXRe1Fien
/YqzN2FqRMKXhtBilWr0gX5r53/MSiJuww9NJN1xX1BDziToBgg5HvtbPcDbK+vm
6AGatU+3HQE/QMBxapzeKluFX++vRMjBSIIkbY2QFNGPg+eqls7F4u5eK+Y1xTfA
bUHyr6wDgbpsMw+Ry+3GV/COShglK12QM6/tOCBezV9f9/iDMhuF6dXuqyh6XUTV
V9NPmGJfEDUgSaoSkpfd7c8GHdQvWvZmk5ZXbpSreTvgHz8vyFB2qzR+uetSlYtK
gDD0UNro84GlEDg56ouTZD81vrromE5It262nxQT5/uLOznGKO6GjALlxEWfKx8t
u6YWiMIdq7Dp6rYUC7Z4qN8Orv1FlcunnMxsJfuLM/gEz3aTG83DN4Pl/h9StjJM
KVuZ0g3WcCtDlKbO4966cZOc1TNzKR8hBcUcc1rPgUe/tHFKsyoEOA7LKGdSD3PM
ON1uc5cY6S8GrVE6yB2jfY78QdOI9LmBG4f6YDag0cJSRJ/WpEHoKBNe+pZZY67j
N16RkgPMpKxsFvqrEpi1s2kuxa7yyNPdOn3XBV8AeLm4Gxs3fEUjbl9xcKvWVt9m
TiyhDdNm6/+K6tK6CmcqSKTwXRPo7addUFNMrqurbG8nvgGR2gExw27bbl3Id3+E
l73+F0XBQ6pU952m6q6/DV026W7gg3eU+0mjqC3E8Bjj35fHlyo3wfkXsdgpgqLW
oLQHBFNk4gXjt+L0MsTrrLrrTL5GqOrLUC+cHBYbNHWGFMbAhclGHD8/vcLFF/q3
7NGVBkYH8f2RN1Pdh+RvwQT3IkvGRc8T5yneSW1PuhKUOAN+LvhgJ2irsxjfuAWL
vEOrrBygq3dQsgLANamOc5Vw14D+lm5MuTucNfUvPQ4ZZe+m1J4xpvlZO7Jb0qJS
src27pNSB9w1Ipo7FF1Jx0jHHefi4vsS3tM9nPa373mc1WXalOE40bjo3l867Epz
opJphh1ZqwliWATfdQ+Zu4qF9be7l5gHnyM7CG1ONWsJQKKwYt8W8POmiWcM9w42
1DgIUlZ8B8TEoZmIeobPeG8DHny5/bEg/hFcuoIinl84k713yvAqrh7cWxU4Dp/4
M8oko1WS/PzK2lG91vA7D/dXxVBKFz9a9qYpDzluJ5sbAcFzRYv+P5IaDVIsFcxU
Fgh7HqiT6DmnIl0jbxwFD7j0ITulY6K5RloK1j5BDjFgMORK2JGOCJaHvuLVKUYW
CxBnshcVVFnhc1W79LFI7RP+A55e2gkeID5MefVEKWMHGWPyJXLVYScWCTXNr0ti
U1HTRYfG6O9s/Z3xCfy/jp9RIXHV46/0gVxK31V7L7Ql0bFpynq/EPLBmKMYrgTK
c8r3axfn99AWDZ90a7NKbewWInFB6VdSj34rmPK0LEjBHbpuatwzbWQ+Ny4rewa2
JDpoltISdkA5te6K8w1MlNNmweh52U//Gj9yyXb2qbO3f5+nHB4ItvDpsj3d7JvW
ecL7y8V4Cc6GWNKoRxI+izMh5Cuz6b1eMq4/zK7SjW2utj4WwNAew0ZWpOMzz9Wn
0GWJmdkCPUkjm0w3ubkhkTcr8nfoHqL0ZaOk68yIwgxGpwrsGaq7GHhihW3ZJ4H4
HbmBa5ur4vtW4WoUVjcOIBjbZCcdGAJx0R2sY10G5tyHjqENSSMFEXWTAC5IQ4fk
qjlclHcG1ZjKY21gGRgBJuZ/CFu59LzHqlqkFhEznZcldiy2pWdKPePzbR+Ei/K6
FZdDpN2mcqA9qHLF9jR6F8N31NCWQqedzL0bi8qFVNhF3ealv79/Wn/vp1anqGaf
InXHpGRb9pYTCEcSOWJ2GIIuEAkEyxV44kq+t6nwJaT7m2EoCaV3NaPysbxe5xhs
Ok79VpI2YkEZDRYgvfDv/h4z6Lj2J+ikU8+mmg4HXDW/P64dpMSbYwPdqwVN75Ei
FLY65Bz7kLmXuo6ErWVbfR1Qg/Y36SmJ2PZ1krf5Y9ODXhnvUYIDvSaiZUxZ44x0
+ncfofCr0Od6GrjHjD4744iujyjkoIp1zRTKHS3Z46zWYdVRqeKApuq8iAwFoMd+
4CQvLXLXryrDx+iZ4VMZzlDhw8DNycfh4W/d1RrLr3HCWHd2CRIzti4lSLPlmsAl
R6g1dP8bTXuqN2L13A1Ga96Fb1S3D1e6IURKHbryITATbfd0qtgPUIIMp7cFKGpz
aG52mduITtDDOhaj0sbyB6twZZG8VgGM2+IOmxfsnA91po7qlUV/JIuQ9oRyg6x8
JGyL4HlHYk+19cAQXT18GbDg3/w0aZmQvrtYyPuTWlTzAK4fyf3paXxCWyR4MU3z
6jo4TtSYOAErAeyKDMUfOEyd6uAY5xpd2t1iKcJA04R+/e+1mTvJJRQBI6+otnR1
8YLMwYxgN11KHfDQKWf5pae8c200fENfoyRjIlE1fNOMBC7NKGXoKoDz3+v7WnEd
np3VLcOdhc2JcTDvvYq+4ZjjZ1H61frteep4HyDemS1l7ZfrLbi0lNZ5ryj7RuGu
/x5Tk+Qk63E5LRUkmCe5q5j87n6DpvSV3BU/zSUn+JAEPrBMPjY+kFBmtoBQcJWR
1V7CwflIgxX+a/b0MRhKLeWA8Q377S1wM/t/EEHlLfAwckZoPSCCJ5rh8fbbvyfx
sF+7eJW/dZxqR4taPO4KfjYrAoSEIfJqh11FAyzUAnI5kxACRtJvNBUyYjzVZ+LZ
ZbPU91Ijob3OmdGTmoO1btD/Cv1cOT/Fui6vWy5AtpKzbSB/8vFv7LjMzCjnHRzQ
+e8qbDmEh5/yUUFE911UQ3+Xkuqo0SmAiCwvJ9WfIb1hLI14x2MI+VO6rny2lAoW
uWWmq6igBJV0nEAgrNsZyBL7KLzEUqFyQxxcNidgFmtlbRqxkRVm7HbTqhxuAve/
5iUacSV1+j8oKqLO9TW68e2/62sckKyd1jDYQQLlkF8f77chYoUe+fUsiFQSJNgo
cM9nSXJCTVFWeMKsKNx1yg5cW1qQXq2vyqcTokU2ZUYgKrQJahhgGIbmavZWnZ78
tLbp+lzJ7SQ4di6/ILILAg6BNvHyi22pKZ2FomfNn1D6TV2tv7Flv/KhGcc0EMd1
LcO06YT3x6Ao7QqcCPH+Bey2yP56QfhibpiFqQt/A+0RB3JUHdlffGCSi5WNoK0h
0Iay/ymZ1uyWfMeie0bnobM/a7h9VOgDMhiozwfly/4beRhVXot0AZanWHChuXv7
duDlYHVxG7MPDwJDOmbdr/e34OQKPt8uJlYShLRmmxuwPjjlKoXTkcWsx+bQddIc
IxsdgD1JSsuhf4QCrNq6G5Vp45IQDfjNrHGo9uEhJdo4Knqh8j1uJX0DMlC2u6eo
WEBOoF1mDivRDXQButjvWtHgc4C9C+I/9qyph+Z2pbQS+6E5k8BxkY/DeUMqli+L
CbwOx3yhWzOyRuYb0U/U0LksZVkm8m9ASawWIArWpsbMpenqPNpPiB5vMnh5OXQ0
+91pmfjWlhfTpZSgTLsmISwYN35gfOwJJpbz0h1A3tYsI9q76ZQ88gOuM3ccwcIo
tbQMatf+cIEQ5lMs6HP6yZrjXb3bd4pFyFcCobuzSVQU2aIPOvgUfYlv4s/+omZm
JAQi8YcB7ykcJ5s+VS/TeweMq6+GLxHMHe7jwNdvm+l5PZJSxXizisRVTX3fNym2
oBTQJCT3MZN/i6KxVXHI/Yb6vH3XRXuTdmoldsCnmIrkd27TP+tDvOes0rfo0qn3
tt6JNWiRMFSabcnBRVB093YC091AnJRdio6chbg0+7OCDoNvsj8TR3X2EzGovrWz
Y3pnSMmMFt1A0RGFCQfzI+IUpECvO2KysRvcXuvn6MHm7xd1W1RL/ku6vLC33z3B
h1RyX/uOQ3GJYlZGstn4j9B5rGU7OtjasQKsUBMdZnZmBAtGn0AZuouIbmGLR+Qt
iFTmOoIph7XCtzVAqJbsF7M2UR1p4GmZnKPNnTHuurQ0O790KGHQ5J+GupBfs2K9
9b4BQUoB4+oMJtyIo9WbXDGtwbgVfxmuc2qBQu1VyLXWrsbDlkZQHpySlb2T83vW
gwOcoCFydfTZ4tVJOjzbZzrpnQIDIFfUoMjA8xfyeqHgtF+mJ6Ldkrc4HdSe3ZU8
eEQiwSCIngtpKM1laHRKr9lBiQf7YqrRm9eV1kvnACtM+JRXBpobbS1KHLq8JFL+
lU8yPsamLZEM9TI0p8wy6xcKzhjyydwC4nNMRlwnUe5C8MarDT4oFhKP/khPoIPY
886iGZGSC3YMvukWq7ZO5FM3LRygtc1fxoIc+swCpIcp2Ds04gBlmLu6b5T8H/KA
VEvTkQI4HaI0U8MHZ//KgBJZc53mkMdVsVSvMj50CI4sirfeXI3gs01bNjHho1Bb
hXOz1Shc/nk+pwgE690XougH3RoZA8T/gj0e5ESM/m0JYgANM9Nh1NJoYlZQ/EZS
Iz3YTMLa50E7f1b+4MOqAGq/g6+GfxcsEBe03eZryiam3UA6VQmFATbg1QVUUMV9
OJE5OuJAACqC8wDDBP63X01SnmebvJmAhAI6xQ4EdE7etyt06WUhPkSqhmKPEQl8
mfURix9BFFOaTM6JWNFVmHSFCxHpuDkZBQfnNLDZm57Z7Het4hJDlVR7AX+nIJGU
DlBmrqBgeew0zXIRc0RhcB0oEXqqtNYLArmXiJGDxUgK4zfiXudMs5V3lA0628jT
JJTkXq1Rmy7P80Id7FGsGVD4PFyK4q6nSYCPRUspnPnH1xzXbcQcawStVe3iVR1t
uMK9p6AOz/cMA0oAqYXb+b+o3ZuJbyyDGcWcVdIuuKfEbp2/9nslVZGrw9m2hF1r
mdGZB890bq4dds/eb6DVNCVks7AGe6KKS0l9I+i7nW5kIjlyuH7FS+C2k3MZ8tdx
KH+Hd4dClzNQtZ61hPRgtlpauwvubx6cy8ISjA3MLGIcHYqfn8v6cHvrMinNqTIQ
TdBR9q2Vyhx/vMONlG3yWqYzDBc1NyKjr43ZO+Ml+61bJ317wcRSn+WatQMZhr7W
o4sEh0wwARYI8+F5afqry1m6gseTnuvYjhigVeJTDYQG/hwNp0tJ4CQjYPGX88yK
xROP83E58NkiJ2DqX2GLeJzEFCb/Rbocb4a2jxwdSkSG4qUS6HbG5QLpuwYsIBi3
Lo4xKos047E+jD9E8QHdyDXsnX5bDOVhtMfuSl03Emk7O+9MhRVyKidZTTRngtkD
rvivk93VyQ+7O9FCBkzaB9z+HTT4nNlslm743PzFo1MfMAFGTsDxFdLBhZn2QQuN
hi+w5cPP+PT1Amo5oqXjo5ohkAxglTZpkiUrecNW9W1MLp+Mjcodn9gq6l8K3SwL
+d8+5V1QwTWB8oV3F9bF86sDGaJMVUr979PVFHb175pMVJXTdi7zGcaNRFIJ9iIJ
B4Lj86vfT1jn/Z7pWMZp6eJaNGBhXJ0efGj26Gpu03UmM7qyT5HhdGHNqzp6nnA2
CYyDaxq6cCbc0mOVevfCJBKSpQh1FKhyCbIay3kYXESusYnBB7hr77EWG3EORGVb
nNc3ukfkApwcV4OxHn4lce6J/ZFAP5XiF9joZ/Nhl1pqQ67GAUKwGyDm94mf0jk/
5Du2EHUInmE3EdmBJ5a6IrdTQ0S7aC9EPy/r6jbqU+ixLpFLdfjjfZN/+HpA975U
YQWjJC5LsIwf8Xwgq/cDEcMUUjemHBanjQnsJsP4+FwLkbl7RED0wj4nuhLat2eg
f3TdtyMCRbsKCoImrbqaWMD3GXOyxuWVuLkt8lkD809Yl3hsCDvzuUtHYLlL74ke
ZYGVXXZ2ik3QrQiTv5CcxwPobJljiIQqV9y9lJ4ps4V+fOM4L1/kslROOrISjcyB
QJtIn8qvFlHKdJwXJt0eKIlrGR3ZznJOZfenQemT8HKHVkjs8SizAvKTwDy0pDVv
FbSpBUEFyLDHe1tcs22EfZ9OyJ8++Ia7KRw2uBkBrmixr0xnHypTN7uGzkraTakk
zPDfzja3QtZfGrfkPWIta89OzGSVGEJpSbVE7BCjf3SuFcZaBl6hIpfdKyIcgDKJ
IbPj9TE9xSkAb/L1ZGmH1QR/b/3/idT3A+ePsOLVZP4GS509xgJm/ohRgfNfeovD
teMPnOdVu1n6n9VRYANvdsI+uTTZlFUg9ZoD/SQzzkdET4yom6HQQ7tMPX/wtOjJ
7TRXEYH7uw7sIlJe2hNQWqzhhck04/GsF22CdLXShKdU0JmZ+RGGEgxX74++9HwG
LLgxaU4rCsMzUuBM21uVNQeEPig8IoMgFQfqGnJFY7j5pboYHqIGPDz3bLsT3G+d
KrGfnlH4ZXRqJmPLCwXmy+puO6sPIrYY02SJB+QzHaKDGIIvP6RTDrbi2Tg9CAso
0sApHi95/h4BPV0jagaYPh/ABwNkUueYAIhXaoK9AVRikTtJz5Bx/NBem3PfOqNV
Bcl5jzdx2Hvyfgy1f8wBKD3VSqdImbcrMFvDV4QJbD39lcEMuLXv8YLbXbnU+I7c
aULgeJprBWqyHCpf0tb//okdCVIlGVRXxGiltpNtqei0HKGS0gdv1unlGywwaB7A
KcbQB+kwENOh3CofomrTfJ4RgquvX28AE4BMtkh1SQorCeiMglzi4BV6zYS+Zbr+
zSNW3qSBkGZawPuPqAPlYNzPy4bm6CA86bS9Pr9XNqD+NDzP3O7gK9F7eID8C3e0
KtFGfUs/ujqmXTTx2Tn52BnY6YE3NcJZxx4rBrPWfH0SVGhaqyBeQoD0ny80BiIn
ee/uI0rIeMwW4uWGMFIYY9VUl975MarfRETn2piATXkOrtbM/ahiY2kIb7DzQFok
V3GQ0glfeUD3pOkBMHvdLucX6qQPbQybTOL72vJbC0mpzdb2oOQGK+K0gSfR1+E5
LmBmVUF27dwdyDeFxphon5w/m7oL9H4E3G7z6J25vGdtongY++qU7azo+VilM9YH
3bb7CVhMEWvOLw6CgvAJit/3aIWWmb8LdmYew4JZEf9ypgUn1PgDpmWjGCUsZkog
kHRsXZnc8BiVmUWcq6IZc5QCrqgAQMbz2fJjr4WRZSEsI761lvrFhk07oQ/g1UV8
SI/j+gMeScsQJGpMUCVOSGBhnXbwY86/7cXlcp9GLKvj44WnGNGjawspbLgJIj5y
r5GiccFOV/SLhf7TgoeRXXtxoK9wC/hFfFpL66ueWyFHOuQ/BKik8TIWLo4QcNUw
7dwmqT93kGj+jmFvkEomZ4f4QxLF0DuFobk8lASG38Btdo7LkqdlfMYcmUEAkaD1
riZS3ZFZaAypHVSuRoQwx/L4WnsG8gLranBCCV8gJMmLCZRRSAtuhZ+uEgeCaoyz
uJMIsDyZBUqaEm/6XNbZWZa2b6Mjz7WF3oKghsq2gJfDRDnCOWig9EpvULRUo0af
wB5d+yms1Vp+VJW3DOFFs9i5CCGmOMjZJ8e4ql6m29t16b/Cr2WANLH4J1BZOTsh
5ZTY+XjHBNwAw2FiK1bDSyQjDPlcu+kQoE1KAgPXpr/0y6J50/sRV/EM0Zy9Jgno
V9eBuUNYXg3c8Gm8L1ZfwP5Rn/ItEO5pu6+DZf4e0TYIDNjp5DgqaQ/AjYf4Nmfs
niDl/SAZTdcts107xDQvsG4MF5fHA0co9Asb/6/U1x525ALG5ceQrHkR0aZdLGms
ZJctazsY1g+zRsd+q6oFo/OJX0h6Mf+JVAoib4+FmDCZ24kHuClTT/lmQuVfEdMh
rqQZPIuiBkYs2LOFGm9hB0Zapf04Vfk7zAgEw1nbXXv30bzbgc90FeBRM0gtYXsf
8UZAre28uHyfJhttcRynuHICib4j58AxPKDj252DWuPxHhpl/EIwXlaJuUpKshbE
mIbJH3N+Mh43OfqrH05evtWb6gLSUNfgKiDHbACcnOE7CbNpyXCkxD0+upmWNqXU
n+L+TkWE1tqVLWH1gv1j6WtPaAXK24Cb34CB/YI9hrQkdznCKpOdG2mMHQSV/6ym
zCspeFnKLntkliQOJB6jv+EgYHuieq+/W7zzeW5HjZeEY2t1+xCi5rNA8zoxR9xE
ZEWqjXUUvQG8Wy08SZrhNPHd1Fy4INrGZZiz1cQPtlYkujunWecWKalBq0WAn2E5
uUuWmpK9eu4KUqA402AsWUv/CRZABKRifsMC86xIhdeFS+ILuMGfFgobrVRCrBZL
BsbQxADgsuy/We9Fj0MF4FjJ/WHThs72WMMTiMy5FO+jaEKTT66KUBAVHYG6o2iM
3HUwmOQ/FI+/PjcTzU8IghjBJ6bupkoQ5vyrsVkk1r1M+T204IZHonPmmzzNmpRM
9fcnlK1e9VAqh9HIEn4/smDP/bdTCXQJWTHKtFZRArTiVwdakm1zvBE3dPX4ZPOm
ATgmb/xSWHXIKoP189fiEtv4W0JtiVCWQYtf6lAhh5wSWV71TKPokNbZxfeLpLvO
73Hq4m3ye41/f5KWWfmQeCj4JRwqWgqGHoN7JDAvmWa0IShhORtpMM2IY2yqkWFD
Cu2ju4B2ZHce0UQYljhj3veX1Pahljxa1EdC6vu5pVYbGN3Up2jvsJpufc8kUUJm
ZwDLxQwBHGOc2hAEgnckK3EE2A/kd0FklqzbG4AWeErpz/xPueyI/2ZcB0DvTT44
aJrRg+SXGxMxnqeRw8UBo4ZaYh56xgyDB5CFCEDCZ9XBgn5lF3lyAD8/CXjzcELy
tnFBNmG8LDOw3VeKIHaWQitKxw6yMunssS5JvbtIxXDmSOKwrdFYopu+6xlQQmmM
sS8S270ZMM4lkxGvtuHgKJSUHkb9pdFbg1oNU3mRyeLSS3eE9kGgLqrnnX1rjXBh
a7IoPP8VnifXkvMsCTpvCFOAy5d76HdiEN/8o4cZHUJT4b/G0N73qFhyyhQEiRZq
Tu5B0YkNL0E74XA2stEc/EUl5NDn5kQ9gNNPwsRi7nODg324zF2BcMaB6kMTHbhx
yjPftkOXXckpdbt48500AQHuttbVLMWduNFBrt/XFc9wy/ol1IGzN91SKoFDrLur
J6ymEtoO3QweD1ZS76y9J7SZRtAh0DetcnehIar1cb10S3U/6EoeyjZhaK2HqkIv
EyhsK2SIlQydLFyMndzw2QTi3ZCpdFIfcNTbGxLTIKZ7iVhmfUZ012PSFFfXlyt5
fYvC7o6ouNRMW1rWikUtJ8FBLOQCbs0VOsowP23UShCLTE7XN7idJI6dUlrSNGtu
f551fXd7VtzSIrTkXqEBUUjhxBLBSkXFKPRfWPFXVlM4DbW3fhQLlL6Y4cBvC7FE
Hsm88Sts/G53m2vtnBq1R14DYVllUmINUhSPCVRUWdjBHcrNQ+aG77cjrvzBvAWl
yc8rDWQrsLSkpbcvTcklQgCBxxm/2ev4VHnjeMpdFzC33UVr20SljcsRBqJXK72b
Ro0nHL5aIZPwnSrSDFYt1hYOqpkgRHQ9hAWvVihQ/Fmxj9ajZC5JXER6VlYoLip/
nrwXtyyP3/necNeFdaB5yfjYVSQpnaPl0d1tVe/7jGXTClWyl90KBTn0eULHXWfk
vKeEK7Rn1hxQQqiOGoGdmhqlJeWi6JUL+TMFp8LazcrTb8JS/zY8gZqa2r8hnfl3
nN0Ad7YA59gBXVwKBJC7Ykz2CIUNlHwB/P7w9dSnBGR88ufBWGpeTw8TxvBXmDco
OAI3ab39237hpsyG0N4vzfB7IsjLbkertTgJjGkzC/l6EXa3RwhuqjxeGug5UHpy
PRHf3VNPSQrm/fj1262n8e/c3YqsDqZHHnxczaKWzEddcIhifTBZUbmROyVgireY
BvugLH/S5vo6VD9acrkzY5cIkQ65COsIhIZMNCPWwVkBfK1SPYcWiwbhx8d62+eb
nug1xF+S4siZonMu42dll/nqbBjaKeHwGuEhOszr/ZpBxMqe4Sr6MIOKtmE59pHg
VRRV4sKSPIG+vnF5cGvEnNfAbsWdFa77WIIjxSpthXUjOIuvmPuQFTTJEm0S9Kwl
Cg7JyNNYsMNgEbp8nGDgSV9hKJ9hkt7QwMF/asVIaEIkPswu4uAzezp2Blo8Z6xs
MKMebD6nBMzxG/3FmoHG3VXQXl4t0pS5fE6Em8pTASQzlNxk276ybVbFxwBkpeVw
ZofDkHdwQ27AILP31rWFCjO3sk1QIa7oDllaJTiGbCGz8SRYwDTKioUvIn2qtDAp
EZD8RKilxmeI0/39mhajqgc7kWxa55x/Y35VgJajk97mzv7ZHONhb3vNg6Y/EmW7
DvE44qiLHJ2N3nt0I4YVFB/6gwOaDn3W2NgY2rqHZMgf+MSHO6frPRcfCp7CwG5A
lniYvgMjYReNKwDZN6J9Q1EIerDojTxRP/LIXDzKmh4JD/5TZ0woUwCFoWvm3bTr
ClecOycZMQ9u1TfOQv4sh+RXUHDeblRj5lNG+CUqSzKyVjc+B/0PW2z7Ha0YhykG
UZA5uq6htd5Tvn8EW2X5aaD2shZs1aoBA18c2+o46M5cvPo9OLHimRtddJPExr5B
7xsJyTE6YkYPpRFyf7jWjw3svnduQIvuIX+akkp3BmsoOykFwS1LkB6zsB+2NwP1
iUbFlZip4Le+DqGpmSBfoaxrjsNRUsxiv2vZDWGqo97me6RqCrdtb6IJCBX29c/u
EUpRhR0CboNmjabvqADP+F3Y/DScrg4Uo+cV3MlgPD2UslomUEJDbwG87QXI4Fkz
coA6KySPotZ4qW5sD0iXjVTdTjSNTFIjhhwsv6P1ijFWA6PHei4ifm3EenEw2bLs
v17LJxvVAF55NFNxIB4r97pXjh1TCZUJXWeg7IOSE+E6F0jhTw7/enrczDrQuhBJ
MYe8eAZavPltQ3fsb374pDw1FoYwXamLdkWTovDhtpURx8xFJlOW2sOoG8sdo/HR
6B+b5ZZ6Jw3vZpzMhdEQ9I5VHy87dQ1mnkBclQYYqILsbXxcdjdWvUqvSZJwP0EJ
XHniHs6xOVDXWCTQUCsGgMwUShG+OWOClAuETrIAw5GmU4L1hDCkV14OJkJ3B4xx
voSGPN9o027iM3XRvjG2269u2QjSDLU2lsCrQ4QtOtgl4Drg3oF5rbwXagwYLE6T
c6iCRq6gokrZ3Z2qjEsPet1b/qVXWcr0H5uozdAsKY5B0aI6Mzqj67hqxDmzFKTe
1wSZRnWgJ3HFIxfmPFpuZvzC5AFqPTbMNkgimQiRu03rQfqdboj9qqDVYEWa1CYo
y3d5QoaGukB28OUyhG6ytcXuOXyWuK9F7knqt2WGdOjxUCnp5RoiUuz7mAA5BSoL
fLmm+SuAf/PRw9G6cTzT60N/HiALHfxLHyeumUNGNM+496e7iC8GhILJjNnLCdcn
s/w6HeMd463tf/Uj3KjOdaocNFspvEUmnUMrXLkDI6hGCovTNGZyAp/amRd1Cp1g
btLP3HEAur92TEkOeQ1+UtHm7/oC7TyR18HsCtb04ZSQtwAq9Vr4kcktZiOn1vF1
VbS+HaEChBV3BQXrXURIZRVg2v/4E7lsHqbV0lN0RgAW3xMpXs7nAoYJdrxUr371
TCqZOd2O85ePqdaLvCCIUgeICpF+LnsetZp893EbuzlZUhIOliRE/5AWTrJpEiNT
pWGuIGA092bF8lnc8wkxXn6jkz7XgH6qYpi7l9Z+fTlsmteJM0gohhmr8lzCMe9+
r9JvO6JkvBhEIAe5yfyvoVSyn+PbpbiSMvkz0IGzO/6PKqlmMNMbruaEkUEYWrqE
OBGWMRnbY6zWeQYv+LtINkZDERhaInhmRdvrpCSAoA3U4EbPfYmuVRSrUvRlEoS+
EBtHe9ngrtX3s1ul6MmcFKF5g3rrYV5MLoWBYW5W3ECzXqBgjSjyY2JxZhh3yflw
ruvwLnAsomUZht9rFZZlc13na3RDAuW95z8FJ/SHgVPaCI2a+7T4vmF2bsDDUNFW
BwnIvVMx/TBAtMcnv6ykKgdBf/vkA5UJxFi+A1j0LsdFeX/Wt7HOYVC33dXJSv0/
SqZuiujyzT3XVO4ETDFCM0lSmfnhglZ8SsnswtkIUpGSh7lMXd4I3OKhTywGE/Pr
OT2g95EsTBOhkLDI4Helqb8jzRU4ppi3+/YDSB6w3X9In+LGJf+FvqPfT09rV+iF
+pLrHESCukC4W/CxxebgQKbiZ0NJLHW06qaurvS7IX4uMt0vrFT9kNP/gxo/89v/
6rDhzoKRKjVgEWUSg05UhxfoJXBAzxyhI0CtIA8vT4YA64aifQzxSPsxPjnOb6jP
nmeOwOlyFy4FKiU/dNun1XRkfAxl2yqjsbrhMZi/TclpKdsDJhX3SWu/qO9dlJAA
z3eGHI9i/i+SaOnktK8JI/cnXAc85xs4gmIT3uW2oadn/mlYN6u1umW6cvzDDOn5
OJaLdgfK89B9bP0K9sFtqXRtLqwNZhcY1cmYJ1E7En7XrHhtJHYYgTh4G2cN/VaU
m81ebexsjU6ipoG/hmajaH6kDt46MOpXsehAyKjiuvQ0q8bL9rW0j+gYVHq3tJpj
PhS3pYtdA64kNHEa8V0D7xQW9cicWNW/R1XYAMem/UYmxUnTpdqIlswc+hvbZcsg
NlIEFXGI2SgYvLwCENbffjKlIABZNlgYXaw5HD5qzirIdk3jXAvqxN5+kkTsWdU4
nnCIrzrZOtIXH86I1xxBhmo90fF3li42teTcm5U1g47DpwCqrfoozYEI/6tMjD40
q2XrH5BN5AU2HXCPl7/5j3ftLN+0zZEbT2AnfKqc/ZfamWcFnP4bMK609VIWfEhh
PlV7LGumgiS8WACF4/9pDxUDzyxPkfYlL1GpUfc+gGJKv72iuIDZuD1cqMGQ/v+A
4pRSz/mfe8gInDJWSDIqeh9lsiAvI3mJcecHa5peDBs70KZzPNloCJlGVyv00K7P
rR5Iy6AABSPwAHQ7CtBHJB85k893Vb845OMjj5rQMNLYVWyfrOyEzaXtzMowx9oF
xW/ZhNx/mrSvCLedLNYen1kLYJM+m6iSxxN7Lf6dPVAd6W0Y+P7PrGbk7FAifYeY
lJLaqZ2nJavkF3EF0oScLX/2qyMLZNKm8SGIPjBBcewkhTG06GJuuROj0OpRFDxd
ibH1bAzdpz0GKjZDeVVp8OswWpRa6BOKBpG7tn+uaNJnFcZEIkMe83GgFyGoXnKd
JM8xq/v+M2ss+Jr7B6mEFsdmYnLId8bl1H0Wm1bpUs4ZA2+MB9zsi2CSxESf2opj
d9MB5Q5BMSPe8V7fCY1hrGon5209xg1JclNL6k67qsqQBOAyqMMsVcPCCeqwk75K
QOfbHrNHBw50fT+tm/xBRoOBuVIAdoIdbYo6dTXMfYvzCpHX6ges6QVcM9Iri/tA
rHyuOD/4E2OaUb3VTirV/MpM5WrkfYZyBzundSaxJwWhADCroUszcbPUarOjs7ks
wf4Yd8bP5p8zn5GsarbypPMys1GDoInSf79qExShjhOO59YiPgVRv9cxxx9GzuaR
aJZ/Pg+KPLfyfeEce3X1i48VIJfsBB5DpOC6/wNSvvYAw7ifYJ8arVN87dEBqEq/
wRuMKXpBAKzs5DinSqAurnZ+9+wo+lwjlc5ldidEaM6wGrlu3OZr8QVZaWDpSp6a
P3ZCYpzPiY7NSAPKkJQolZmFB6t4lPNK56LbWAFkVgdsYRWTt4BbK1r/PtSgtv8+
e2CKsRfL3S/KNdsXnZ1e1E+KpOo+NjQb312WDXfD26qHOBSCNqmR8bzRkwKyUNxO
Gkh+QdC3OZjIHDncvIIqhnp9edSGOIAdtuzgH/9PlXUgrIfHwI5PjhV3Shc2dTZI
kyop12rLvwxESd0SIhf471M62qfZ21xa2bcvjtMjRtP9vlhwlKFY4KUzFJbAHJxG
unAh/AB0HWe/v5NjOnxfWXTcJ2VC9azA7XdjwZzcCefapWhcZDPQjPMqk6KiFjVB
ErrXaiEsU9s4SMjqATUeaLmGDyNF0ux7bqBCcqZ/taeWNgW7GRgASTrOei/rsKEt
XbRWwOTFl+Qs98RUeOLDQ8ByrQiYljS2ip2vIlyV/BlcbtysUxH7aCxpOqcQsFkf
MujYQ5zQh6dDP7Lfl7J8/EeAiSEEnaLljrNwteXWw0gnyCVQh8wbRkQcprDFA6u9
nz5V6W8h4HfhBU9hTPmaKevM51gjyZg0FEQQpo+DGOYaY/a1udfFrLVGIu3OLYss
PsMxkUvaIwFpMOYmM8b03Rw1FhLMGb9B9ez58kN8CqLXxnDYWEV4WA7No+ArOarU
XE1DFRXr9wDNHY9WxnJAQyQ43C2x0QL+ZkLbfVeb+K5s24QlbWdebf2dwmGwEusx
smxyM5Dl1in37Gs91uc4Ov4k+VwuPsJfjB/g9E73ChzFOnHAdhbxGcMqP3n03/rf
TyCD3xG+PB2OGOpanX2xj4vfQpBJKJCW/1Rac8tcN/+e/5sK6dzu+tmINgB3Lsuk
acvtSb1YPROZ6OxFukqhXVTjzMsStImrIH2KAjgBhsGZBuAKVEaqRxBylONPvLpC
JYWFqz8TzSyu6MTOZDlMKLbuH4c00FHpMonCwCnMSyqHVFdO8TkI9RW/8fc8Vo2E
VeORqeoHxUPMYpH+R9IGQiIapFZA7th1CzwA6SM/A1wLzSECRSpnP0DsPW4a0kT6
0XPOqqIqg3TetNBqh8M/NF3fuOUZ8lpSDa/APWNpFcSLfLFewtznveShEE7RgJlC
tjT4NuxDDJynDw+Zubq1u0PKpu+YrycUm4RAL5S+bb4Ow3SOKN6tIEKPB9cDZBcU
IgJ89Aebw+6A8xcHhcDIKwaRP/kLn5kE+5pFdgcuPiXLAACWAl0pCHjBXxRc1aSA
4/AZWB4T3VFiVdE7y8sH376wjEHN0aJpj0Q7binQ/m1tyjbUZYBwz2EMEpSHYVHH
9CUvjMOMkQg5K2U/cbrpbY3DnQUshuHB2qZlLLOVCyhbhRxCrGE3bEwQcqhgz3i+
q8SG2OYrV3bERvhtRn4f1U3hMV8FuFqf1xJq8BiHPX0sZ0LnSi+WV9lJfXsneAqh
8yOLT14/+G+YrJTflgPes9fV0dZV8y98Essj27kNX5ul+AW5DqIxCUoOuu+LFLtC
4qk5Bo8anZ8LLR1t49y03xH9ytam28hVA4lUeilTum3S7ktpqFLIlvBHlqR5iDpc
stYdaYB3wZo/FeN7sP2dCTcoJlOxpQfZ+b9DRCKsVADedhBNJJgNJTWBcxDyqshA
C/sKQlQakv58MBFC9yE4FDekLFcRuTjytdUnz/ts8JGwBJQVxDYnOCqXI6Vkraju
chMzv2SKKgtx+K8do8B89nikY21VhyNmG8CNvzpfNgcTPE3LfBXY/BalvQgEJEha
jkvKlT/qcKRs3vJ/yUVL29wYJ3J+bbkYBfdZvsD+rJQLQxzpZIUw0jcy9mJknvB/
FMBuyealHFktHSzjSvLMAFXxIprRzCHmccuy5kFJbuqyNZDHYFpAC4JKKRKoVn5n
x1umL3BELPEmfv3eCZuh+CNcZhZKF5pLvsc8w10WOwbl8EM03iLUh8A/z4R8vlWQ
+sqneeDyb2E62p+wOre7/KybjhIJM8X8u/LOHthdydByPjGTYXDBxy2iip+6G109
X0rlU9WLtYSHrtVQRY8BbsYRROxWHChhXK7ZxVasSJ0cSL4fzOQ+KMQIiB7bn7FN
1Ggx26nyXB4OWkhU4PvXCUXgHjUcJOk1mwsAR8V02o5sIKTZh3CcCsknquaQ8EF2
dwMCm1KC02C14RB2H/th5RhSX5vVTlCOSQso9NRxeNKD804P2l1X0aGp4Kp19APc
Wr2wHvLr0GBz5yUrvbRr/O/mQ2gzj3G8Dfk1DuODHVB7C9pHDo8ztdQqBj6HwthW
r4ts5LHf7MKLlE3pDlAeMn/6TPiUZJHW9tHFg7o5L5TgsqBl4jC7hN9Ct9Q7hnI5
xxPL6rYNSURMqA2AMRSvzwRABZa5xKRBbFF3RZHfoB3FxRmhzX6mRubsvESaikhM
6AY4kdSEObjI0RNpx5XxZ9yPYRVxkKgAyniB+TAJ00cBKM2CiwYU5mAoj1a9x5qa
bYiLWU67h73MxRb4bcoVKDDQkrcSiAzKrft9ZxqF0P0ZQ1TXrHOvIFP3V2DQtEfZ
vJRYnRLmaq5/nKsRe4Wm1QGmwd83lbhU/9xtIyDk6dVLYqaRJBekQ1zBxcf+RmNU
f1wYO2F/JCIPrUz8cmFw7ewQfDQAjvR3HElmJ1PiFmknXuNR6YklVN4HCo4MbHsv
017bLMYJVH6qvlxU62bcf7SZkqOhPOHPSFN/pAmwB0aYZAV682h/efoA+05ENyBu
42PFEkiEAny9xgcYZcYgP6UlSfK9svClr6VmFalwZz/2oYUe+oyQusKntwflRNHr
VdD2NI99zmQpAf+aH1Qcz0hM9zfVzYV6FwwWDNVfgzKapNSVTg5RTdj3VcCTseRp
PRrfNm5q7szkbnmA6vCcUjL5lI6/jlqJkI05Mo3zrE9MfJ7krl0ef6xHDQRMyKfu
qNfDfddJvmuBMQGT1XnydrrD6Q7U5blbgD7DE+HRPghNDhNxpBqOHm/h7Dn8eHeP
8cLRUgbPDR3L/Xid2qqkSgfjQgaCA6l697wz5yC9qHJH1kJQviXnxw//9l1P07Up
o7kT3XEeaOch/lZutR9REZTeuDI4Mo47l0hnh7eo7SC3YnPOK/ic3AZo1eiEJbQl
4Mszji/vC0rTfZjKph3hmpRt1Ykm/r1Wu2hfwt0Df46Sawkgpfm+hoP5yjDHDTZe
uPf1Us6JITeU5gBvuEN5SWZ86SVS4ptyYhqh1mbfi17/jE8wmLG0QUszGW+g4TKe
tSEFF+rgSW6BDDmcsUA/JBzBqkKLLtFqKXZhL7MHZLdUNOEHCzwh2+l9fr1RjVGi
dOCw7DRbErYeGdYpFywwe4ant4f7dxvnkMNOnUlKKOYBCuejgc3IXI3SIP7/k5Ma
aFmzjS0Riix9PR8+B6lSUpb/AFL2WuGlVNwoRQ9y579nSga2dOEQ6EUdq2g9UVW1
OUFInCyx4d/U5JR6ao5ustCkuVDf3Y5ExYzKEGJN5g0e2megTUPWtS8hEziFRkm4
J+UZeXOg4C5VK9EbbS64Z8PxiASkogKQQa1k7GpI+mpF9KmJQ8lDKHi+J9UNvsTU
85aJ6Ss6pm3CrTjJANgTdyHfDqKBwuPsQQBVAKD2ddH9zr49UHVpP1nkwmaAaEMc
7Ngl4MES3V5gYiEpKZ7tehe2OnKuNRffqiJhlt8B75OUcIvAqGMKHQNNw2AKcf0A
qHn2/OVX88ND8/SYR4WRQvgOTMgJL34eOhUIEi5HnNIl4JmPFE2lzu8QtA7d892J
c8XKv6yXEShsKj9wyo0Og3Ma4fkLs0DWEQk/Fuo/gr0bKmQW/3gASW34qvLdRUlo
i1jXaM4+7kJDgss71CiI0i7zkrLiEoYFyMr3xJmqUrVsHKE57JSyARuLMYfiZgbb
PPLcDRVT57OPoucLoVKAHN4bBlmAzFF/TqoAmqdFsco99CAmRjjaJlTI2JWWMEMH
KsS6GizlmeYKbK3baMqLJetO+D+dMD/hNqj5LgQ1Z9HOSNBpU6kcRJulo+pQbNxf
jiow0Ch2RCzTQ1UyosEOLYRYgSpp8WuQAGiqR7OrGHgW8ACXtSjr7oaCQOCvGfwq
rWmTTBuPYprziKWzlDGTpypDpzF9V615YvegoKodORg3c6/Z2JI5F5aYvOosQ9YD
IcXBx3J9N6AVr2lWe2sJhbyTN/aHtTqGplZfPuzCRYmgo7qTKPUCQmhLGviSpD/0
2QoBWaBpCWFAhTZCK7SU6qm+0NfWWH77iuLDXrhx63s9x0f3IagiB45+1uBHQAeI
QOe7n5KSmJ/2aiYJALSkr/Yo5TIIvfAo6lr/C3J7u0ByoL/Gj/LjTctsL4mR0x2M
ZYRSvQ5RDNjK28KxNECJ4680LAmh9tpo8L17gUKUpsVXCN2EesJGY0okMXCGLpPD
5qJyKzyca3a7JbcOsYh8HP7+3rZExER9175IBH3MkXSBlhPxeMqSixHDwfv2bDkX
mEM9gGCFS4Ec8M6GJGn+aCcfQymdL/OGHKUSbOIE9R3qmOZnp8/nN0bHD7ONcgFr
BiZGx48t2MGQ+6yLkcnh3Y/+DfAwOK/t3DBuJe5Txj8qfUoV901ddQ3M1UtwLxtC
nvBpD+cftqsMZPcAAdJurV3Dty9SZ1g8HGo7dJWaA+8bILEZ4+0Vx5RTm3FLja5W
ZmVyJ6AHeC6gVKpwkv/KuDrSBPPZUUGes7OBXNuqZpASdYKm5TjvLLMTRO6TuGVD
hYRL198TNvR15opdmiRQK5HjdFdoFAHzgmfuRh1vgVB569sdfkBpLVMZyoBw/Rk1
QFeegNVeXNsVILcSt38gn/N7SLCfdFt0DJ3WewyObPt86waa19m2GUgCKw6WqEb7
F1InHq7AsqdQEwBlZQinOJm1lXGvWmVwedspC0IIn+crLS+GnNAevE8TcINM6gb6
k6dFt9yA+jTBmaqJfSRIOyq6tBW4AmvmJcz+miDQRdUtPL3YDEcidunJwJ/fF9ok
mgYDhTLOfKt+nKc15KSm/PfA5VVRh96wMZTOSmMXe4Dh+9t7Xpk3yGkcl5eS6EQP
CBecgKvWpLuArCaSe9dLst9IF2AY0MdXMANO950w3cSbh+7JVFeWe71QxMShS29M
ulFRUUoepDHsoF5PhGtNVbI1iPzv78BpHZ0aFWxQRDxwNY7Dr6xULGjWkZwWM/hx
PAKCbezFqHGnJyExBEAYbHpGnbBG5xy2EV/YGBw58KtOAF/xzM/eUw28L54vvbhF
CMrjHFDL7Md/ddUhcMpraX60fKLGzzAoepkey72tpVjgkHbD2ZC2VNC6jZf4RJuy
0BIbWqLSoYCrPYmbynM5AII/TFODOYE/aIM7JHAMuwuvpQjyev6iB07mnGm8u4rt
JWvaH5ERRBPUudsBizBIGI/CcDplNYPe3j+M5wLwcRUIdOkczWka24LtT+mDyxm7
HBKGZGbqTfT4Lv+wYE9f0Y/R3d8hFjAM/xFmI1buyCyFKzbu0QqOX7aNdvnsdmhv
+aqPVqiWTAAKQ+l7zlX0NHgdMRmtxpSXc3ai/58UrBZ4h8D9UqlmSelutMWKIqxN
GhwDr5wqpUUR42HNij97R6HVHif42BaM+G+8Ap4T3hd0KP9fc3MkcsAmP02fIE94
B7kei9IPAWkNCnzdGUTSGmRsAK76AI0IzSSzJDRkNdnWCVi3Ullk59gkjzzG4aGa
KkqqlHvQN+rsEsFA7j5eQxKD5iHXUF7FjEcthHG9NgqUQk7SDHKHoGrNkyir4Ae9
+QqiSmysmxjVRDcm5Lm4Ft2DoAURmhFV/hmgSxOIcDn477KXL5ShDRNyG6y3UxPk
vBTF89WRyUqOkvNl+XeiogTJswE1bQUkD0zQPKGAGgEe5bRH7lpuQzo5VyPKgMRM
PdOFSW5B0oKg5+Tk3vNNmc8LO96L5UQtfDzhNAk6vm5YA1FUEeRm70Sir4hNMmTc
3aYUmQv1+XzbqL8u9w3bf8FGt1kHxmTUKJigS8x4NagdV9uANwRxsKlnkTElx1QG
0XbP+64Hs3Yu70Y420B111JXyCNxQuNljITU7/IX8CdXSkWiO0tEiM5I7jolEWcV
iAWaFgdGnPcCfdcBU0M/jzMT7aNp8k1IEQVHHNChv+d4/A/QkfbYCaGQGG4adOau
MQIJWLCofrwsoakCpOZn6L0LBYnZEW1O2ojHC0OLjfnQJQr8yznG6wXyAjg3UNvk
zd9fft36cWQxX98N2x1tG/7NP3S2ufqm8+T+Hj5Qm8peuE8VrQZ9Te2SezYHGWX0
z7FreLZEqFa4WT6ashZjDvmcCItnycQpc5kB8MiMuxE+LuZS252awnFULp/7ZTmt
Mm35CUhf+9RF7KkvMKAHJcWDoluz0V0NRpz3/Z/zLcyGTdPkPDwYkLxdowM/YXTh
+neNdaxuEoOFO3AC6hWqLGB3d0dtEzmhcL+55cVaL3Lxkk4LEE+dXEdiKnOLUv+K
l976rRQSI3F0w3Z8/US84gLS9Jy+XG/TlLv/knzKbFCTMc4+wG/lg47nWZMp5zv8
jkTea8c8H5AEDaXAKNLhc4OzxhUoT7bt7jOPj5aOXRep148/hy/a1B5FPFCzSoUj
GPamDMl1CLxzpnqBB7LR31m67SMVNIEo4HCDzUr03StPPb09zqk0Z14UrxapG/N2
HJu+Js1hwQ0RTcC/H6qYcC2wT0lulwIdB76yVHnLHhfcgFbKRB7ltiPCQjjGJGe3
YKpkRNnQ1hPDrjh4PbL6vukfFRX70Jjkj8XnTxzrSWe8+7TrxGTqI8g6BrYrKwQu
xIFyQfbtha6ieOtg4pcY8o8i/g2Wkdxua5FEFmClYE17ok7mys8IO284ESzvILSL
XjNIeZi7mU7eo8HDMBNN2AAgEsCTW03ix7+Go3mS9gRLaL4VLhh3Ez4hO8FWset+
LvgE+pSZZD/buW5wbBtiPnXIRdTJyfwunnniiAzIO6LIDsn3Yi+Dc+ehiu7MH8YX
DKPyjszEL7cxjQp00BGBReLQQVOfvPw+/2+oT+WkPd2CdcMaz65xQkvuqQ8bPtN3
QqtMr31nPoT9Y/t/b/1/hcT6GiyqWI1pMD3KpWR77FUzTMx1N/A/w7YIZ/qFtlJz
Ju9UjosYPEFXM/by0st+uL8gcoG0Kj4qHtD91onf03asv4QTtL+zGh+ZS0GdiHlF
kn7A3daIG+pfUflEatyBpc0UsfUGEpyom/7EsEu3kEuWDlcfgPwxMlqWl+/cfTu0
t5fClErV3kpYiege1dyocbBMwustmxtsZ2wbknk920Gby+TjvU9elOAizEphnc0v
2HXJMQEUXqzmN+2JcAqv/xP7zQ9hfKcAGvXE2Xku07uq2/nHWzm2xj7cnePvx+I/
hoXELgab8K0cjj9d09RsIXb7MiSfTAlgyq/OklHMMofAKi0TZerFSeExYwYR85Db
BZrWbJ+JUijlz22xHFpCE5QxUKC/GFtU9JFSL4OPHwtAJ436rG5IKMEEfzJYmsTB
j1oL5NFMuha4IupvDGhwgg7ftSAuTqozntVT6UB3+su4vmryn8bTjO5OshVLL5OW
F+D89A/JEEq12gHrNLA99BkoSNE2EhhihZYiOgxddDr2SlCDMW0bMNsEX/JA4680
99mlDAYrySJFZQmvHyFFjRBIjdimrtVmkDep4x27aIN386flQM6eEJDmcnmfTLCD
ixcRl+7rp2XUfnO2EZGPA31CmW5qcQBomBWJNi4pG0wvhPpbiqBXTkTTiVBzw/Zs
+9t2RNuH+eoZcQPG9fgb0aFGjHiRXYQhBufnhsXwV5vKLmbzzO8mPSwPMtlX45Xi
jmslYXnSQgVF7iOiQRMNmY5HRDpLOKD9Xq+XmTwWMx3//nOZPyjdyrtRC3w1B1Ch
0CZ43Gj6wTU426ddh72VzvxQuaM7icIcwgDA76IBpE7JI6299MAiCG1b+h1AFfwh
q006HlLgMDQuPUWaZwnTMW2mN478C/StU6uezqH/ro5e8FzNAiLakiR7041sZRzX
kG6Lad4FrpTwiBb4nIOO2IJNNYw2as/lb3VFbdwRAHv0GbrpJUcrLfeWhORMwDG8
AgHR8fcyxHXhqM+gHfp3xdR4OzlN2EmHjixejDqSPqcMwQpj5O7/X6VeEqpVHdfl
pJerjs0R2nRfy+b7ZSRJ/CLkel8iFo6cCYpd3AyAzBN+Q+cqGlDM8wZL24488kGa
Ra1janEuK49GGMrRXevQpUGlHeE0K4Uk/wkvrunFcxprAV/mtLBw/hbILpzcJG1L
GFXpTHuGksmwgX7DSiXw/T3S88u3Fa6d4imRRoLs16IIqQyjkGIB5oxAq1V+5fs/
4IGmdkM2NH3uVyoHr2+wsWfQcnpaGYL9OwahZjSRZxurPkiNORmPyM2x8rP8czLK
2Lx4Uh95U7uLx46JWzCy2xS0RrYMlSOP3Ip5oFndsdCLkbYDBVlu8rX2i8OahY8+
Lq2bAazRN2bvHVkCT4S8Z0k1EWeDqTOw6P/AIe0YxpqYc6rCJWaHnr8kV6z3Ni+S
96H4M0oc8raH44FX7xhgo/VQw4HCpCIk/td6utP6rUns1WZzy9KICmkGtIoNSZO5
C0k6qGvIRIdCa0/IBjfGo58AtSWwgZ6RaCK9XeqOYcYKTH8OQlfrTNf2cWyPK5uq
R3+LkZX+rOIb6j0dLtkMiC1OcsCRE+gNfTE9swRRtSS9H7eLthjDd5tkCk4SlMjh
PX7ipTnIuQQ+kTwiy6nhTNt9ihYUDqreW3QwwkKNIbO3cuqfwcRjkhoQy8hFSEbQ
0LdIV1PWROgaAvUft0GXS0KS7wtNOfxe7usnNBgXyshY9mN703h7Ks8MqJ6ieRiA
k4O2HrYUAO2TQnflTgzTpBkcw0Fkmg8H2UzaJLrToAt4+ye0Z7E6Jt9a5tf8UUy3
SCImwQdlxRKkPeGv/yUTtM2SYp+dKcs50mcsiiE075nv8UTIjwnr00jEhXB6UI/C
pqW6pVry8tYslDsC/EqdZfhULKvi2IYdlidJr5uB8Ar5UJ+RpAj6Ch54hu7LHvC6
EbTK6pV9RBI1IFVXsIU14wHFf6hYdA++yXP4hyRfcATe7Q+viNve3HPmzuw9Xb5S
q8HAQPoClLAxCAFBD0UNjtv+Yft41jZ5LJGyd6LBsR6RCp9DJAvIGS55oknezUkA
0zevkqYZpAsr/h0Tn+FFKP0r+hoF9+b3X/7R2zLgpbn3KgPVe+VNlUByTq6raxfQ
2AdOjhvCi58/NwiB/zMroflNRS8oNJVnfXJsIZ8+O6pVeWc2jhbv/pNLnFG6yags
Qq1RnYLhm+zFsgipfogZsm8+ZoI0ePE1fVE8GVWQtslANSBwE5GqZ87Ifc0RxgdF
LKiLQa8YNKPWAOWEM+hUoLFccrqD8SfLGoDFKIpUHjI/v2xbTEFKHmnqiJc+sHwk
w8NlvM7irsM7XOxxOtmmR3PneUNZCt7+VOBbdHEye1iKR3daDAGZb9w3n52IPIpe
9B4CvTfs7S62mb4uXznc6jnb/514W7dSqumVdseCTRR1SpsOAH+Cmw86Rmbt9PVZ
7ylcv/CODMoKIK+DcvmQ2DEJVC7xKbxuQv8KWWBx+aqLF32HNr9iR62cGS0NTMuC
lrECeeH/VnSzKuo15Y+kFHgiru8Hct7yo0zwTHQRZ+sqWAIGaoYydoGYCq0itsWG
jqTZEY3JW6MZaUdHH1hB3/cT5LkgyJar2fkX7wMeiPawKRrVO9S3+PpYf+UBxit9
SIg8ApMJLvZn2CJjB26QH4DlK3Zn5FSk7AArJZSiFwxNevcFmU4GLhoxe+iUQQ+K
kGlRKqhwUFYDLEmMtKpnr/SO7g2gDtDKkCPxfVRnpBhj9aHDnbhcGoPfoB0RQt6o
YX+nmTxDp7wR+XhdUf9JywvVfHx0SuRTXKy2nI79fGOtK3cWw5Xmi+pWLkMxN8JV
H7u8hI6O4fnNnXrg1Bd0gp7eM0FGU7rhAn8HPqCmE9cKLImoYnr+l88boGet3wRK
xjidGlZ8a71Fev13BrbWoBN6w5xgRl+SlZcp6/9mFvWdXuswCfsLiH/W05/Jw5xi
4g95fkWwGdYNcBRvXtpQbp/H6RD7dDL+tLuAe5Zi/uN77/QLdDUW06Vhr1WotJGq
5To3AEhO6sssrq5AZIZFxBdC2n5vmeGDCKlKqIeUHTEJym/9GUeN01wzA6ueFdsj
8qRc0aqQRu84IPmnDqwOxNmB+rflB9n+Xe+o6Xe5HzzKfgX+WpqfsgVRnfwy5g0v
oWmkMbZIDx4LJ/2BsITxm8eElgTo4AUS2+WX+QfY4+Jusw/O+mtZo1jiX463ZCi3
aj5P1J6KHYdzTW4uwMHitnPTuezq02dKSS3uy/CG1GgB2rHDPLkTjbT88AA1SPiI
186cR8aFrHlyzSLbIQYZW7Y8pxn308PbK4NsXrCGhtusckAHsNhJcppUUsirEjgb
ZasKRBwo+HoEm5qKtMMdo4g81Q7nCrJP5P9YovI+K4hmWNA5+kSIhY0mYeYpvAOz
5G0V8vB61iyDva9GDoJkDMEmVW8AUrXhon+Z1nyeo5CjvHmU3jrLFxMpKtVS8jcM
ondwTkqjwQyyKepiuukJwQ/R35P27xvCYjWTwmVGb4mw1k+iDPzkW6i4cQnY+QOz
I7UfNWtQVJaltEHTqkfUnXW6QMsd4pOImi5tlyX8v8hxDEFdiCZPFi17VJQrdmyk
M8fOJekg5AeXDxfp1ewA/41Yar+zJkZDRvDzDT7pK1u+Q26AgWR4Lg3vBMsAwkiM
YzFEikG25OgXCXVWy/4R45M0+XdEFj7Yzqqq/CUJJrMwN3GyQsQLTbo8Ru+gJXBn
LJhchbHEy0rNOseFnJQWbeuH+ol15wisOy343lMkqeMvQ8mvsMxm4fUgyciCiDvN
izWMKPJE4zKVimyLgM+EJmxMNKj4WpcJJRtemEMSlGyZtWz8YUWwAMA0P3FKZkRj
tV0NryJiqydgKxN63S609R1Bxv1zCLyBMoFGlwP2uzbJQbBwlD6KDVWoRDSDe083
GYE6ShmrtUIC32iLMfrKtQMj+QtPjlwUnT9pX6OKp36WLUwJGBaFnKvtX9H/o1qy
QXlXbGTOvc46YkW8D1YBa4o6X0kzwsKZhp5zlKOZJI2AAdo+vlsQclr1zm200yy8
6EcHGjTXYfi1haUqRzmgY+GH5mDZtvksBvSx3VcCX/W230pbxr6uWEfVL+6cZdh5
OVeNX0J7Rfs2UzUSLfR9s2oq4Qe3j5iGqL50LjH/VrJsIr/EQYW4ZLTOZa9dbfa+
1AL9wdZnGy5A6BNdkdaXrEDHANcVhc4zsJDsv3Jb/3tmzUAcOpuXHhEahB/ibdvn
vZ1I69YoTvanKmEosf0aWhcweF/wfRmn0w0y9KpV20OM/QbAtMXXxi0A6KnD9llv
f/h1HaHBIYM+C9VGLSshr07MwCU9RX/QmywP0uZJIYc6XtM92alZndFE6DT54VGT
XIHzd9wMGIhLBuxztvghPMW3O1T119Z8zmWoHFO1Vde6npVp4nPpgy1w3FPQ4MXK
muqGSk6Y3Xz+wXrmQuiYg6dmihtjCqF+lwMIsb4RloR4J3iWNFLgrhulgoBBF1KI
VeT7pa9RepZo4SKWDiN94a1d8aO6odIUiCJ3CbCjW6gAQguljsc8j2fFu5hMyFLB
ePA+UL/lLpVeOx9HzKua4frb2ZQtnhKLUBApY6DNSVlfE7NQS8elUfEL9AfO+oVh
5GL+nhMrPq1MCsUiptoKfpHiOnqlkQac8KIOrremP1dgcn2t41YH4yckrzfJzDVl
q+mSCPKqs1VKVdjreyHI/qg2DWl/R8E3Ra7gZm2c8f0Rb+4jNaiZQgbquaFX3oez
NXBvra+oJxu6RKcrdz22q4auIOMC0rZqBwpYcX8MWy3OVBeU7kRp2oWLoogvlwBJ
OfAsWSnbcxHj7v3X0E9TOhpWr5M74rmNYVOEKI0xiWyNHT9vK+zUpr6okcMKX6PB
ANwYo795MBqYk5OP368kfcNoncc0Oc58I7B/g/GsrzvvtcR9cZ+q9kQMWOlwB4sW
/RlH6nmNdlanhbjoSfRBWPnLKUZmB5hx+gFfks+Fu1HF1UFSxhzew/IHnFM4/IaA
Fy0lTNb7mNXTBYR0Covde+GlbyIFyCvcwl0jm4QRdR/Ms2LWWrf/7tYNAdVzhU9X
PdSfIYBaKXTGjKFFIpZ4Hx24acIFxygmX8fv7ae7GXNoSes20pSfaKLEhaWBMSty
9Iw24Ju40iiev2fqT+4OTCjwJndzeKamW7f2EcCVTxvQlgvZLGQN5olPktG8txq3
0r7zZuinwfULwZakHfyAQMsk7fz14EC/kqdYMEHB9yySH+MlRlZ+EuFvcLQBN8s9
Tcgfmfl9fW/VUOZkYwEqc0gCnhzF3/8XIiiYepNQRQgitzYUCLUYXzGY1S9yWRrp
pvKhAjduPJDEm3V5nuYpgSHw9HYzl9JOVC7IxfSPo7Lzv3TOo55K/NGPh5RTegy1
gIHeV2ThJQRfsVtlHH5t074rYR5h2rOHggwXj1v+GZFn40zaJlMn7ZYGxGg4P4vb
9oaTHAVHrIwxN1C6hYiCHvfK+qsS5VLAQCAPai29dKpiw5tUTZv4j1Tsjaro2+4B
rjw5IapkY0F6EBKEy4d5hkt/siNi4bU6FJdYGvoUgQgwjgAVfniBSnYlUOtPqLCn
2ysoHMkgwuUqgBt0V7vsJj9cbkt2hwcbIifithjVaGB0WuBI6mILtDR8cEPDXJC4
Vw0VcUZG5lTsgfrf0PS1+8cx0EQGxHzI4CTTNHjyJHQbOrTvixslYD6b3iSW+PX4
Hzy7Z5i6lPbTknctC/XT2KYW4XK64ZX8voa10WwXBpE2+XA7LRhgZEI8U2lJzmoY
GFVnO7pgVSLcsZgu78mSsnLYEUhn4cmr6Ac0i3zOkdxnUJYH5MA7npRg7QEFb5Xq
9RuBVVAT9mqpFeeQQmAxFZqDop4xCodmHJYRxq4wF20v+xr4Xy6uFE1CLjG9Wg/F
H2oWRhGZOkKTYmEQ2eoUzz97ydr2KbZ2K8UXi5Fa82bgbFFtsAA1A4IFpsDHwRi9
KcQC4Jch1loVQ4CVbEt7dIp4UPTVpP48Av+xd8QnnfPv/jEiZx8qDqFz0cOXklDm
zal365cAaPZKJ5cJ7oaaafd+vKkifXZb0ptFKX11t7JVvLMU5cxOfAF/cKHPrVtB
RZ1G9ZyG+Tcp8/Du+M4fq3Qf6x4IjqGaM3rXhRU1Su3MWFYnNhZFaq7JwpUPi3BF
r1xCV8aanMPKQHTmjCsGwNeglTPaofUxjvNzf34RC0CJcfFOvahYTuLJPo47mlfw
/mzjkTsvlhfwnWC+KeGp9hMa8uS3rcp2Nlakb4QJkuqp//KPuHyPXjiWbtw5U7wP
ttY8ULQmxUFl8v2aCiJTairfijhpIhfe4Zf0tSXCyRnEGw/AOneuJ0LjMbkblDJI
95xaw5e3gyPFna6sp9gqAZLLAMz2AARBe2VtN8/X+hLslkhE71RbqiQbs2fzWrBz
2U6uwWZDUOdAVGd67pM6lqucOkaillWr8k/et66ybnGybNTiqDCbx4Nijzk3n6OD
3yAIjM/717/27uKawb2QEnmratiLU6Kt49zhMjN81/61pQp59Pbwiu3FUPei0Y6I
/6hLr1IvTD1Q8gFkIyJXQOGV/smkK6q5uKx5zWzamXQCo/ROkb9BlDKvnMZMcESE
k2chTVL8Tl6tltJnUCSLNmWw7WYQ5Jo0AJiCyJ1mqlzIY61DkB85F3pZ6yQZ3Bi/
AQmX06ZvKhyM8JUCLX07IfpUkW+2TplroiG8xaVK9Xjk2Mq9J2ZJNU+kvKQwDs4/
lNPw/IX2oiIUQY8idpkxY7rvo3M3c0lbGRcnC7XGYm6VNZWXanlOEyLQSzV2HNxP
WaU+yz/v7gdaFMVq8XG2BXhIKZBMsz+NOUe5FjSR1bMW10sA7an1voB4K1QBu4dW
Oi/X6xjTyx2m9AsdrGMgHlJWB4KmD60PLx2LJ7AJxlTNZG1UAaq5tI/wn/wK8CIE
n4ps5exsGvP/c2N+psQ+F3smfBwUNS/70hTdu+Jf7GdiNnH50EOqo6u+2qqnIC+H
1s0s/yjksqtiQTU/QdqO0WNlCSl5gTxC5ZeeZ2/fFHaft3HYJZ03hju1fbG7bjft
ZXiU7MbHO1e8JZWCwuyeuMoQZnYvfKEIz3TdxoE9TFXexsY/EuPb+B3+jXY5y9PQ
/A6+eFYdI2gpvpq0caKN5/Uzcr2ZmVluxsENT6+xK0RgsxEQG1YwvN7xBYbk2Jqe
WXhmufhDlGF4qyvqHMXt2x03ejZW8WJIZbpG9o7lS5NupB25sdoL3lb4NdEwlBu/
ABdUmUB821FvHcQkbgGgKWk13jHCrpg6vFacECPEzAa56xwTnm0ctV2swlEmFQrh
DKobssp2qGC0K4gE9Z1LRnqovZryFUR/RJeoTf8HZI8V2gw25r13QahvAxCKTr53
45qER4Belv96LsXfEAunEWWmMfeq137vYzrV26uKnZej/PqliV0FUbL0M+nxEer6
4w/iyJk5738uJG22mXCn0NA7Mg9ccnFQXxuDcprY2aBAv1NqUosP3UE9mczy7k0e
TCXhFP6F1PS0XtGYoy//D4jtDsYYKB51BnHIYdvADZCSe6C4cYukStaIgVqJQswE
/iMgAAmFLxnOomau07MnDNrLHVmzuw1RyT4GZ8MATdrLHt0yTVS6o6xuVCbCWeeZ
PBQ/ZW1WcVMoPYqEN7sIqhO8YDahlag89bNEX2/SGbxvto0tHE8gJ4j3v0560CWa
Kc3KElndFfMRN7rHWlbAYY/QYf6nYHU8sv+uORIk1mDOKq5jRV7T6tMUVnOD5rGg
OxSKF7CXWtO6SClK3YW9Tdf4tNnZpTvL0OkP574XTNVTu5PbC7BCWBMAnjGWcRUY
vVQxAOMO0ffafd0mggb0jHRKNqKLAr7iEG9gYd/foPZDAZEtvqxwu6RKkzlobrdR
HV3R8BjjKoSP0seOqw9B3+GkTSWrjYKr06FB6L2IEaJs9Gz2yznvvOrUj7d/sIEc
gIYqaEXhdr9x3PHurecrnoTLJVu+OgDpOsatHbsRXszSvjJ22GE8v7847COVOn4V
wwMH4rus/tkudpAptMklv1YiKoQSKLTGfFCqTigMV8IX8RCEM8KnyyN+wDj6dY69
jtUpDy29xZzYlGWbj2cMIpL/OaQYd5cMRGS+irinnhM2u09/lWLN9bb88VrNFNa+
9uk7L7vCo+RGNuHsMIj62dQiV8DIHxipriGtrvE+xUVOqPerIYpsdRAzqU7kxFkt
aA6/Poeopl4XCDctW+ympAEiwGRgSI+5aDN1gZJWesWClLpvVK6m0tAnXq+VxeB6
RQ0aXxjpfRkG3oxmuRVMhxZDIEf000w97FCn2al5TbzSruEIGdxRqvzSlN0gxlG7
DCcTTat6xIFSExtiF6zEm2ns0MOoC4FDBHG3NVnmlLucjILfYAe9jruMwo+h8PXg
As4lyr7YHKwJkHvCTdQlOk5Ww6M+d/FYkxzzU2i2Drq7kNxmpPKty+P4ZVALh61O
1B0K6gCivbQnzLd5Enm2VsildAl3fKxNsdKfWSWdf2JNsHchqp6PHd9EyTY4gADh
ELSALyaNH/5BNNOcEDbOY0A8FddP4Ayhqq/cxhg7eEYtJJ67c7vajV+CZoCSWcyd
fsp/KFcc49E927HvKJFxpPl0Yz3k7jRIG81n5tN1Ctvz85NtBlbnEVCNBS0FGUzr
mSM3HV0zhI7U/MijoAk25F97yRqNmQtMVeGKX3D8WO3rSK/w8QOeQiaSOm69RDw3
zQD6sCexjXrsccbDWWK/mv7042hhn008jNCjuL0TZTdmT8EaNVHXLIrH0p7OtDFJ
a9y70JQBrjXZvHCxOT8CJbS6Cf6IjceqHU2m691i5J/rsAstq5/gNQAkKkAevmsW
VxIwfh0bPE8GHjXMpRq25kLPlGHNLQDzus7J1xv9iE3K3EszoEMPPa8ecqeTfnZ0
m2Fku4/oargQcMdY0kL+e7aqUekXUHToOeAtpKIjKTjZmv0UpSFcl8hXA8PKjs4B
ddvJHZ066Wc7kOeaVFEW5ZiRYklYrGj/SCxe8/On0wpwKj+EPNuqqcVqi7FOeYY6
qMF6FOHBDqFuq39LEk1t6EwFWaotxbTz1pgdwYeqE4qsT8D7lg6HkO416LROZRdK
xPrB9QECVH3w181qUnlAPNAnoTGWyCNB5XkBUn4B0/LvMmCmhsv2UyjoJMBDKu0/
Lm6grOCCGp7Ip8+p4cvths4SjOaZk0IpSHLpV9mT9ykXCg0HBbkm2gOLysYrLyUD
xFcVtuwmL2n5thRKV8JV4qYz1GPy2EbaDqnSvPo6UYEguTsa+MAuAsM+sbI5Ake/
FevDN5qXTrN6gHn/AsBTNJWg2dGaXWlSAIrIGXd8tt3VagBi1NBE2h45w9X0fF/a
UFmJITKrUyHxf3rBHs6zbEy6Oyrq7j58VKnCLbVRmN0OrHaXdeWDRWFRuMRLIrhw
i1zE5gChFMF/pPdKCBdjePJiyw7UWuBG0BCu1uN2wFMvxioXJ+Ys42eZAuiyElC/
rO+AnpQdNxxiaMl1VeFOK7I1p8zRAtwP9W8rOcG8CEesOCaPimqAbak7IN83zkVq
5qLSzgHpny+G12uff0z33oSZNvCBXpnnY5YVebEOZYzIxDHCMqNmltGti9papom7
64/n7w/kPcn9vi/GxxRWiyb/d8CA3Tm4mAy/Hl7HHpn/IQMzY5QobrkPgw8SOEVv
A9T02UM1TOyRXGs6rz5t99lZPgud/vgsbBYSGJzhAfRn6R998vO2a0eOTIPiIPD6
tY/3uGw30Q81rkdfGt+rBRPmuTgnJkEKi+BeF4Qg5dO+lvRVHkPjNQZvXx3mrkDB
J6bRwSDM7sJaz6rRbw5wU9mMZjG/b2j9nX4fuYN/ERksVon0zv8JYEeFKKFjZBe7
TvY4d3TFGpTk9LipjMnqrQvNV0Y7kj3HIrZ7nUn+nN7iBeuWjQz2S9B1M0BZo6o+
nYuYWsIAjUibxENk5yNqulkob8+qKQuTYbeuKA2v2flrButxv+ssCdPPlrxAYAK5
9WBzPSIBRlgxC6B7dDFRJFM6Y17y06oYMF9iwNOZwsIBwoI+RL9BMaGhBcKdqn35
UGc73omv8pQBzI5glyS7Kiwj+6Z9VPbFJyaVVECRLGagfKc65dM5KB7UP80pkGRw
BQkkNqhOh/ASPGpFX7GTaLf8b+tQsuxFILE4oIYqZ2cFOwoxKY72HerMKlbexSKz
KhhrRSKwyrjUdIwRVwxDY0VyfFHPEnSboW7tvGCfaki4oyCNmVQAdOFygqt5IR65
5vPvPTIgIIT7x9TEbSzRLcRQfwI7yqfUIbElol5BILmwDSz381/KZiOKW+E5tktM
PY6NBhyQyQzG5KPEJjFogqZKAmu9sxR6C2+BOyzECHdkfomgou954eS0u6X9nL/l
s79lMtf/vyduYU78jxTiXZubSQV8a/QvE9lRVUvTCUVBDg/Hdyto7QZjOcPTSXjq
GtnExk+hNPimk7bXqnsuKyHPVwGGfd5BWOAnBhwUBw6tbzZMggnWRVAOVmh8rNXI
s7lDe0nfWzPa6kqLDLhM/x1SD3AFpwulMXH74o8aJRewPOQCyV8+uPkA0yfdru/i
4b5x1ZNmlqM3hg+hsgJ9P7n4QtSFgwjsvYqB5JePu0JwO52b8gKSlapml/V9eQ74
cO5QojRyEewXsDD4hSmPCdM4icvdfBNRJssf9ab7k9vtVddnSCiRgZ4CX9u7fxtO
aBXJJCCvAk4wjua1NfYe5ONwyqes/j1W1f/2HacUahUHB7Xx4tPNPn+qKeJY1aGw
mZy2l/iG5DcqjxpL/sA74oEL3ti1g6Z0dLY1aoWmBKQJoN1GC/No2Y2cunQTY6XR
o8f+1rIkJk9g8DhEui9ixBwftnz2eBop/Kh8EVFKnH6yMNPKi1PSzsw/SfD8gTi2
sU5/CLXKyBtD5njJtHwi093HgwuFBZ+/VVXdaynBs7RRcxHH3mgj/AmTT/XIzyX2
YxIkDIVBVVqm6vIdCiKrKqhCKtKCnvxny3tdQk9nOlWlCEEiRePa2LUtwo9ERp9n
iGJzVq2aI2CLnCn/Z9rKx1s29HTkUmFJW2ShsoFoY8CURn01znktnFNpRFXosFjr
bZQgyfIJ/GQ5M6MrR2sOvP5PR+YfX2ozPvsQMj1oskslgJ4SKCcExMkwNIBSQXmB
HtUtn5mlj8Z4zdFrfkmVSn3be1luJMP99AuEinqPC2LM+gWgz6qLKFQGmT3fTdF0
w3iK1DnSSK80sQm52MLfEusQyCxGA0jIZ32p6Q+3zHUsB6LtxIhfoqxYg5QDAowH
1XAp0FlPTvPHffsUvE/rFgfqwaeeQm74k6oa+TEe/FV7/1DtYQm0oaQbQrVY2xq9
Yt1TYuN+jktUcVoT5ZkB2AKORZzwS+BvW25uFmVHRn7e0oB0uiAK55qVp5f+eCl5
ltmwDLSkb2FS1EvXFXIfNePtvhSGQJKdSUvjHYuu64JXFjSuMgdQCyf3rZunQaDE
0GPjvH1mRomYqvOWFVsdpREcqEBNWFCXfHhgraBEMLI8i3TKgYyS4eYcUZtQn8iR
mOnC1TUpcaATVX0fyeU7FieP/xquO0jwkxdVO7G1WR5VbxdBoBpS0YLAqE848Dgn
3WySkdMt8bP5eEx8Jw6nM5WHNIQXMvRBzj6nO+m4dH+XiE+48344FBKSWmoBW8S6
PcyhcX7Nis0T6pFIvhC5zUkgRCXqd4bKa1HeGb9KESJIOySDNwgPaOUeNgWPmBGX
1FqER2Jl/CnzdntIFKKWmlD325XbQofBD9sR7NVTQYfechcVYXgk+0f1FyEBSQSQ
iKtP2TVGuOKDbMrOEwZ0FSloXvNI9RU5D3mzZEkko0WHEGHDYV03Q7zn+R5KvGsG
ChYBpierkqGdGZY8nuubZEpfJk5hBNBPvXQOy1z/XYnimwhd6zz3QQe4VD8hOLUC
W5rE0bxNTZZkXb8f9zmRmCcKaanSd6l/jPQl2F9xkusoidEXpYesilEKZuCO+2t+
jBbJG9ic8ZYnuRBgez6KwMFxMAuJTdKWTW6R0j1OJODMzURz/ioKBZ+vowOBe5MQ
NHRr5wyCDOSShuVmQLd+fEDJ+J3K83Sa65osUjSlFnpcSlZfhzvGoMTc+ezMXtBJ
QEX2AUQvHP+5+0YJn7exBewaSx/2JeXIHtu2QYohNr8vGo8y9l9OXpU38+wlrAXE
vwnTbUJr2qIt8yTivF0pReE67HikcXMLZtvHmEkYpXvYTDCLifWnAu+d5G1JfqCS
Q6EfBeL6dWudRMv5siv9m6EiU+Y7w0hZ6FxPytxU2F7LhAiNABQoO0fARDlTxZEX
av/1F2f+h6ZH/raBzy8i855mVp4q1aWQ9oQdn/jvGQQlLM6jwIfmrmlw7DQBQ/+3
YYjOQr/t4IqLTgKpAG/IPA/dyV/gw8mhIC5kxva/Lmo4vrNDshkPzozk0OLvbBWe
gqeJYGWcOiKKwoQSGkgLHL8zt4LvtLRiod6020pdJEC+MUH+FGTBYPpy3QHQzjoD
S10ujxxxWwN1Ppql5yPHML6faRUAvl9cZBhlMlBAV0MHLXmPJyLZMI0nQAcj2Oxb
vK3wXgCRw7cI4S34sne1OQj2LBDh6BlsYjvIOQ97R70hnd/mZ9GuiMxo3YL4wYsD
bnQv1vHrN8DvNHOdEM4mSV4yXvfUvyRle1FOZqxVZFsWLq1/L8ezf6L1+HzTseY3
xM+0IMyhCGkbUmcC3RhiFjCw8L1tWA9d9vW7sBs3TYARKoZE8z5Vk78GjTkPiGx4
wKButfwdA6pyBfrN/N7KCMtp/0+pbllmUc53AilkuTEclkkAWUWKR48pfk7cIgv7
RiGLKuvEpDlV9FpsFKQ9oTsw8qeVI6eL1kwcSrh6+FdbHa7zcWxsDq8B7vfiln/s
LcZIXEs5gH0j2CtcSWHuxKxQSAiRH/z0x9gnPZOKRqHr3w1JDcs1w/09VREcnDdc
tqHag5gp0yEXAunl+shSm9+CS14+P2Nf91cg8rSMe2gyOt+BozgbEYdINBo2AoBI
jmZoiRlJOEcArXWTnc50uYrlGqKwf1+RSt95iDczbvfQGxsaYBqGXcpB4kNQPOL2
V5YIfAsY8X/JAHageCjPGV6qLqjkIIVq9vo3lSmvmaLiCHVrhO5LTtBHuJKIz9Fg
hF88nIY1Xs04STdZXEVordjnmsuJySdKAQ+aaDrTo2jDh4bMT/1KsBOv50JrMYV9
2mxJgr1X6teSL3UMrOzYapHdQMxeCz5OQcnS8s2U97kX5JxboYvu+wYhDhiBccM3
yY9KOR00RrP3ldJdU8sT+hyhWeAuLO9BkUFFPqu8cNw+cEM11R/K3jEIDZzKafTV
gwldEfM1yIOoitfV5EfxuhXVe4l7ScvPPZSu3/gLCstbXD++U9xZ2npiY88JXtDA
qnb9shVTINW6aLuOKUV75lDQh+vNNwgkWiaT22mGM5ewvLCpwQgTddNoYitPJtpY
3ZuXlgjIc9Zn/tV3cAKJwITKe2CKUdOTD24b9jegnQ0DPEDyGXcE5zacxCk5+j3F
PPWPtcuu/5Bw++lhTCUMYCjf9GfDqJQE1SQOf0O2jfv5Tw+s7d64sH8xSl5yqGxs
MsTeT4JTaIGUsRRHm9SiaSDUuYnXgBou0owC93hYEhhFtbVgYIT+Vk6aMoEin1pL
j0MKV7RUSKdh/HDWVkw7J7psiSdUwBf2y4lh8LbQVN6JdSSgZGTqeGONuH1U0w9I
WnWO85CeIQ9RsbpcEFAhQZ1+grN5XcrcnpkUpH0Gui+sqOSuJDhKnIrVvfVzA0kc
gl27sGc3xNnfhs+IVFHJ5n4Ddo/7KiOSzPtY7zU05f8u6RSGLbaM+eoIammg8jS/
IeHZM5ob4o3YfS+TBpRdhNBN34WRe+zmMc1pOVD6QMIGUthvtoeCOHbaJRBA2MT/
fNadRKhlXy7FVbhmwldUQU+wnZz72ew1WgPK1DgXIXJ/V3bGBKkGSXFmXYBM9tel
HdzvAW/w7lekQYfsJY+7QHuOq+uMFIYKLOYXnW26Kip4PDi4TupV48mIrtguZHaN
P2hWaJecWwQcfsgXHXCpJjA8QQL4fZUOCvW2r/hV/nPVU7pLZBC6Z3QPSyx1lDBQ
L1vPEUG9QZghGmpvODr6z1nGVGTxyFCFBlpWCYTqymBu+vPhaku31qr4g+zfLFjF
c0jfHNhQm3d2KVdDFPcNEzj71gJlSQGKK9ImVlo9oe+IPPw2XP28PlM/nPpj5rrD
HU5XPWwE7SkUe2imXJFRH2rcmdUCdRk9QCWZelpxrvMa5jI+4ZTc4ruvt7OG2+QZ
3UfErWnn3m/F5MYuagTBZ1rjlhMu5z3dRXRhi0IFdKRbpPLY36u+40nWnMpbVEGQ
0slDe3IyRLFjfh5WqiHfx1YOk6V7pi9hoHF+j2zdJgTuIs8oEgzkLGmIxFjBCVzk
VlAwBiAtC+4A6vm50Y40bfHaBq6Zn2d8Fbqb1Iuo+++/NjuqrfHacpDzab5jS53V
XQd3l1pHchm/4CSMqBY6JXbFMXLwvzZRepRG4lL/GTXP4TX4jDyWXwm4Eg26QBSO
TNLoAj8Il9fQfDMJtOa2YnhhOwWzOoPSCPhD4y43+0ssaOxfu9JhOHBy7B10/e6N
tl1SWV76NcllN8v2VD9c9a0fpJm+JYKY4Gw+wpJQglwQk/Ze+U1OG/gHmSfPOeIi
VtHcbi1gh1k0d7owEVBZs/NnLXL3kjW/TouGMrsqva1CuyGyZ1DyoUNbvUHNL3xN
WkOMsMeV3lN3HW3jep0AMgrw12wh5pTJYiNYHAnOlIoKwvK19WG779CI7AeJ+NK1
2Rt7OhHaOvOSJe3HPMXHdc8adANszFIXhYuvTV/hp01a+sOl5143UDh88O7gyGTM
SjrAsbWHof1TEE2PDPY8BK7owtjEkQ2r1YnyyoR+cxB7/cXdZIfyz8tdBzwv8nMM
be9PsjOZLp8uTU1poAPsTYXTG5na19ZfjB+0Q9KdPDtzstpE6gpyuYHlcq9cKcij
vlmCvCbSxoFDxZ2dcTDHYvCWMW/VjkjBXfzJUZqUUacLrHQXyR2jkDJK4n6V0RGT
sIXDOchEXfhOTM8GNN6/AbQjvxMwhyhTUN9h8HUneNBnbfnFJ3PGKOX1sFyOovL6
6c8xZr0ngifiOjVkR1kbqa9U3461Cj7s4Z28y4RIOD+DZQtk8wQW0sTXM9wqvIJd
CS14n8oXOn4DczsOXp4c1pCBWHGoDv83dOon/MVsB0eVP6hxx6c/T5ayE8h1o9JE
y2iuYKoJCr7TjQ98fPSp5xLzGHK1gwhrHFjabCjL2i/erlUdOT3ygPRb3X6JjoSb
7Qx1ajtOEdAKTCH21b9ni/D2dyNKJLCYgxFfRcOXZRt5TKs6ckf5GcNfDaOUu8aH
57nwFpfcA6zA0XRMb+7aVKB3h+Bvlia1Xc8mrwSDDu+eZ1epfq3w5nVbGwcg2W+H
K3FJGplF9dyPegykOt0zrc9UJh9ElJo3OxXZknXjA788UHVT7QGeW+3IMnd9xO9D
p1O/apnW9lB7DPa6Ra3vI1iOFajgVQJF4E07xukzf20yU8Rq7lJqHdVoPSyAJoLt
TE2EyaYkgpFnBaDh+aKObt56hR3HekSdtHnXrvyNjNvbGG6mhbQj8iFxLOfjqC5/
QSK7mbGWSw1pyrvXQbqlBYJxQ5XXtccQQcdwuhZ6chES+lGbuNVm85k33jCRHPXS
WgOf4yPNvF8M0q8NwP8FbD3myamQHAI8je0q8zm8skSR0ywPBg4/rb3qkfmcLjBW
WltB2qabhkUFReQhCy3yAIsJ+Ur+zT1533wbzORMMEp3OXmS8JZ5XNE3rNkhH5RN
MASuJUtGOxuP1ZVVO8jOoUOKWxctFqK1axDoI4kaqAbwwVb2ZqaDJQqdf6bSMLUr
qtY+r6H5ICWobv20rznNQ12oe++MuAV8NBzIRvhjuki5htyJBKHf0oblrOqqbtWF
dINK248kNfUODrYxKkrFI14SKUtegDn58BOu6nFVjnOknkE7iOp/MKwHe9y69G6T
ezMHkQP9vTWUznAnnc95rLIi+q5zwOSTmKgsLvxExpCtl3B2rNfwL5LilDkc/HvR
DuDtFAD3JpB2/ee9i6GWYHoDHmXk14ju3y11uZbeD4Elr/mU2wChl9TadoePy1b5
Pmnnbpid8ClpuSFd0BDS4tlfcMu5aq1Wo5XidJFES8oJo9THGmtfAXmKAbI3/l64
fy1acgMCBmzv3E8syCyfrK9iBTpdoxoGvyVCnRDOSGTk0Rjz82lOkZFyq4/k2/FG
LZju15V6wu5rlOpCHpDyvwVjfiFAeiLvVZWD+y+rWpbp3No2Acl+HL6WE6g9YdVK
0h/Xs3SGQjC3vMph6f+yv/q5KuGTQiIx4ESTeuijiyC8GUv64Dbt48+gLtgOANLJ
76oAgqDgDH1JnRQZFDxFqCIBJrRLwjGhY7y8TXSrrBTtZeYZbDvWMJKrTFvUUFob
vDr3DMDvvDsW+3UxVBAhtYQ7ozcl5B1zGNxuukpj7t+pf1etIq/U5IIphvgQZBxF
IhAgZDWV2VVMX5oZzVmFmAJ/GyW6Uu7SLDKPgWOVfT/J227NVjpbmddNbhnQOqJM
/m0fsN/eANU3/vCtLszWnKZXWqmkWplyXisf/WOCBKiGbgMAkaPyTgQDN+kBvkVQ
WFscpbQR5tPcvQrFjL1t0Xb8IAh4h5pCpv/U+rJyopTc92IfWvOe7nAuWoABcIMW
4NnCfhifM6JU1MldVvcT0ohLN4t73mVveH5ZxpO7IIAjHi+r529dFK7e3ecarnlu
/UCs0twwVn1/HTHUqcv3h1u/CRKlTbirobuOLin0rMA8BVVbQVtOmP1CJ2aHR4x0
wpBBbBG+gYmPxHU7imMVyGMJCWQXJKN/VBbpfPOuk8K72XmSy/FH0VYWUO1JRV4z
dYuqOfjrL+W611r5tUd7n8U5bXYaQ0B9Me2Dp0muBjFEj1LvHh6rfbvHAEcUlOLi
O9Bov55Gmrmkp72s3q5nagmrNupoddWMXckoB8JxAxPcGtwWRR62L8EDU3YDaWdW
vH5CH03HyWhzv5G09VaGKBSl9DN87IxYYw0KRjeMwYpirHx9c/bc5+LwJFMUYuxX
O5yF5YtMUfCnHKRVgw2azfUQEJET706v+rrNGXF69v9/KwH6sNjtaG8qAcseQjNq
R9Pa5cInHeLF913UDvDeeLm5Wo0tAQSuHMhwOE9nSd3N/AvOwMXZ0fwF0r53+ofA
NFP7i9rN7PZhTR6EkweTQNqSNLXh6u1Gw3w6IOqtJl0Ti6iErvnpCASdkboAK90f
Bacva26B5wJGdM9faNLQxNNWzr6+M5kT1JvoAMH4M8Ros0t0GVRsv3lmqveksXsY
uuEV2BwWDM04g16yiwhSQOfLj0ulWfikW3GZfyT4Ft5gWgt9mPEQqDhpw1P+J0pf
F6+RX11fr2i57UqqGZ6cNi6SAUAp4VjL39Sgs3X6lheKs+afoU7gTZVGz38hbUZ/
WArGZmzl7k88suweC0CmUE1/s0rACA0jkWWkWp8P9fB9+pJnilfMM4R+ieC86Qci
H1/hKhHbt6849peql2Q6nqgV89OE0PG5RBCVDtd/lr/AQarn1FZGiEPXwZJD/wUS
8DaEloTK24jSTNBf6te/njdOJ86ISzi9d1bwQLLKQOqENToCVYbiPivGOYGSB3Lm
UovtT4ad3NbIDvp/lKm6SJo3WrQJClsaiJBfsnoDf8tVQ/eSKE+eOcgwB5o/mb1s
Mn2KPu9U4+WPL6aXwjJwFlkz7y5xzhqvIMGkoHGuaHNBeNZ5COvsgolI6zZvQKYb
3myBfzAANJ+egQdOvZ3+X0xTXpz68+mC7dzUKou8L6oPhXZIZFNrEJqoXK4GEUWX
VlGqH0dOaj9deZPV4Lo7CC+C216VKVu9HbMs+P+I4Wy4ZJBNWdo6EnSkCLjm7Fs7
THsJ8GnkjUL+hEMKhAcWDsojI5fEZCOQECbDh2egV7n7h5kwpeIn9vNl4GtqYvOL
8gWYDC6wJyl6v3NQNIHfcGspDqYlRD9CGxhj/vJkaNr6nJQIZIbVvSCzmRrZ38Ji
onulRbUr4jRk8ZpJOG44Ska/2CuNN0sNCz+H9C9KBCLeiHt8npankGbW5VnFzZ2V
yyVePYgzuCENZamWjEUArKzErFwKn9PvDXHbjk07FnblejQHgEwFMqq15GmoVxcg
xAV+VrqoV9IiE/Zs96AEqud9NfW7D5MsMHmc73H2P6aozDZF2yaL4343t7nLFqki
Op0pLvJ4T3XQqDE8zPQ+4X7SRHFOpaB+BcT4IbTgKrDN4svz1ULKcpBWdD9w6l7w
d6i94pL5ikGSKX3dlWtDYdKu35EJYD0pjPcYM1uMYWOV8rjd1eJ+OP90sxsrCPrA
r/DUcSkGs+B0eZYv9dDANXwxQMfVu0UDT2RApEExEu2qbySou7XubYS5u246VQot
pHZ+7a0pcwUQb3+PSqOIoqyKD9LOUXZFJuT9bJgVZzyaCa81LjyJFl4iAUS40G9i
BdPMtPzxR3sE5Wh478BkQsHqLzZqSoe+9+asfaQdlDYj8wMWmh00L6qivMH1a+pI
ZLzvNKe6u5tV9VyKZRqYcY+fTSUxcoO0w/V01Bq4u8vdOlJz04nVpbSx9tW9ckd4
jRirCV7oYK+L6pByYxQi6V9D7A979XBZIcL2M1NYfM/GsxneBdhSuw0rwj9CWp2p
vLRwxYMqnfD3dGyanXzWAfPh9NBwpaOBxO+SuHsmdk8X6gpv132qIBj5U7GcR4t4
hEF51L3qDuXaansHxMPrtlFfVoj+TBwe13IGJn9LKHPa2eNtnMaSY0KexU64ABuO
U4mLRZLbWbODrpoknd0D1tbjqSVg/1XBurEPqM7yQrvYM8ihEpLVKzroHnJaYzL2
aNadHAQ+f45cKgzwMvDMPF0QWYSU8sITb5bGOIUIOlmaOL8rtFfBIau5mk6yoQ2+
z+jagSptGS6yiPp6UMjbxbnMd7jZeK4vimNz4w9ae2NRrgP1uKgPt9EiIRfH+3MG
hz9RYWBNx1fFsF7/2Ocfs5nDdKyySpQgIS8DQxDmkvvNmltqJHVaWKe9KFE1VKt5
nJAojicFzB4xY4c45/fn4jDkBoGwXeKPBzRS0+2/i2jB2OkB51/GHN/Ba8D8fQmU
gCf/40N8Ch6W5DpbY2IPbHD1w7Pa+1W1hxdrXqTCCRuTf8ay8oinI6VNVplXSv+2
CQ7a22UhTTQwXfg5AEeb2PGDrKa2t6FQqACeHfGF/b0QkiEYER4oX71TKXxBzK6L
gHqvvRlYA77USUCW4bYOj9mIJvK/huR5GE1tQjWMMo/R3stakSWIm8HZZbOydRex
Vpo2I2tTJT37iPuC+E0O36/XjAL12qufn1ZT5w3bSd0aU5pkORdLlS4Wi9hNRr81
LbHvfZw/cUNO0h7UmXjkzJFirzngmDTSlG9MbZpDfFfyQlSw8pYaTYJheSlZy1w6
qgJH/7E7swROoce5VQK4r0zfAg0ep2ffQl5+jWWSvv1Sog2isVUXq7dTeheT/FyL
f1+yEdvznvycQP0DeH8HqoOJ2xjcAl+czhKcjTvVOiRKpWj79IAWvKOBEzdP/st8
j8qfM0ARsvHfm7bnuVjhShjUsvAzIqMDdlmH2DuUYOxynGg6Su5WwD/zTKgiUcED
MMz4O98kHumwLoDWqamtcWgoy+aj8DBwjEyr9OjuPCO5WcKq95mW4WvvqaFXx7rS
JP5GMZSjbYTrJe9JNa59sbsTY95WeEDW2regn+6jhkg7t3vt8czbuVpP5fhE5wK5
W6Bn8rM0yms5i3jB+9/NtWWRqjm7fw1XKUb7xPHVEUhxRclAfAuUD7WAOL5MUMUz
0OIi5t5FiYsNI1ECWZEn86kVhpC6SL0IlrmzFKInCEzFHJ3vi46bG9O/TkfAELWh
SYOaCW+q/k6NkaZhBsFTymhaVeaTdT36P6HejW5T28MRNZhhHxaBPABj95k5zuYu
Z8rHqdxCA7+CaYdbiXmi8L72J27fc3/lBzvpFevMY3ZRA4JmAz/atml4/uOH945q
q7l9P6sB2jWgsNeRD9OSWVNUqaixQayrVdKBnCHNscK0dqrjSWAeKHlqibb/dQm+
G08PB3HkdQqjEe6J2OuSrwx1gBmgkiNuaCzz0XJ3AGI4EaYCyTnYRBIjmL2cYNP0
wqykBxpEhwbRTnxUtvEllVoFByhr0Hab0/olePSQk1kCSvzc37qI7sUbM9tS35Io
yQbZivnm/iq3CHYhMjqhPiRMByGZhL+2qXGYvDvhOFX1pv5rPVAy74V0isJZgQUO
1PStsr6KtosLqbfl97q7/Y9bHLQlYZ1bun8RtccnyJW/sHlHjUFSjbmqujVszQ/4
WorjwlHmeMKQhLb2PR9YK0WKxN+4bkOR+rEzUVaK0gi6csIHcd0ypq6JCp2yOWHG
ZiffGZrwIUHB+fmUBY6fcAFrrnc0nAR6RZFQFvj3ZDfcwrH9nb1E5YlN30G3l1Pz
9Oi1LiitBB2WSAz7lVfH15yUMYVgDQP10/JKpyA+BcCdzmIlJI8sU9VRqJgM4pxN
KWdgEqqJ+UAgHJFF6yvpjFJRJBlDoLeBLQS5Lh0/Bn7lZyj7k8RTlMMpJ5Wo3SrJ
TDACw57Okiy9PneXyBnkz4qS0/UBOd5WQPkWsxMPbUouCQ0edYf84iveUzAsHV8J
krU5dwRoY3oQn5mxPEs7J893ngEAtUcFcl1o78Ql2yq4uk8/iHB9Vk4Vjna47ZfZ
QJiE3Jp98DY38tjIb5IPihRANFFS4qCuYT+mUQaQXPcCMdwDXPWEp6spRnNTtzeL
JhGqp/g6huYoM5+NVpG6tdfM9LGhvYMPtWRcw48Z0aqIcBYihkgcCAc8RwbaF2Gt
t/UnddelmaLTopqC0RunZNy0HX7H5v8+DCRNt+Wa4xs6Cc0uYQ+szcd/6phHEEN5
uBUztwFx+trEu+mAKYUcD2ZRdziFrLPLCILnzfFolm1/8u4aYqqRRlaNh+E+dq8O
hzhCkATq27na5NseEUgWR2QExYIBW2GpvskYe2sH+aC3rTauxv556Pp/nRR/gTuS
qe5xNaiCr00L+tsfk6N8govyfQyZjEv/W7aQDoZ8+stZTGVHKFblNVdtGOHkXu8t
xmxxpabIPLTEbrLoVdkcJN8vItP8XMe2CoHAmo896veOBGhzzo/zBCbMEdEAhQZt
IUL10ajHsgGSmPVyQAFc4Gw5OdDMbFzKTjdWVPBp9o+5/rbkYlYx3RbF8c5ePZz+
BtBAZIjtMx2j9h3pZ/ffexPtfK/UGC/eOsqwK9PBqE+tdZMn+GxxCYlNNHVie/ET
RXcwx05KIhBDqgWievAlIjudjVIk93a9n1xplMYMzZ3W/XBxjaUb21Czjm0Rmaq3
noUoDZ8biq4HkpmyuscYc05KoWOq0VDeAgI1Jr2/iZUFz3Xc1j5KLwH2URlotSgY
NZJL4u2oNImP8XVclq/zm0HgOrx2tUtmKBN6IC2NgR852Ne+Ry6Rfpp1B9aM+AVZ
fFVFJF0W1S1tBIyTbzlJy6WrG40GrmjwMASAbbuZOq7S88rhKggETpPnnASCob5i
PhCJ2WRO4YyUDbXOCRFCG6RiUqRWxrsqHndP1hZ1Jev7saZ64bi/n8swozdgfUTd
PNOMHiGoV7sc7E3skYbVrEmG3ixUxse3jvOnsazbj3Fw1vjbvJsNsWkQJlxvemPx
4QHEGBnfzLZErwgsqV7UK8tOQ6YhDMuf16WpblcdLbJRuWwPayu91tpB0G/rs7nF
mCBlqYqsz4IZVs9UGqr3IzXrAru0/2hGK5KIVAcVH+GC/5ii8HCIzmc8mBlNeXc+
HdJPdKTu1C1qA86nK2etBvBGHyH2cBmtykaMtPFwUQ6d7tE3eqPAmIO4c5NHWmzh
/AZnat3IrEbkQAaU79eXQEj/UgBxJQb+EDD7Mec8zAFC6FL2SH9Q2fYn+Da8t9uM
DjljmZK+oOXkamVx4bdofyg/9/r2q/0l5sSFzriodtOdVB0odvOWIyzb7yFPiT5i
SxAqx6QRlOmTrt1niEs7zGpym0rGRMsJm6xjebckV6izNL7pHOuczVL/WdQ1EKdQ
ySkep23dqQ0EYq6H7qz8qooB8EpC5QBpjaw5THW6zYqExfAWAYFfam5wnzCAg7fQ
O2WMlwusym6CwYQWnwPxOvDhfafw5AbpagaIT0YTxiFUoND52PotJOm7cbhrxWLk
q+u/cnwkqsGxLX9s9c5JT+JsDWzjuI/EtfR3apNYM5rwDF/WnkpUvTTtbOlodJd3
pVimr4QAQMw9Esw881MqZOHdNltlhpRN/EhFqwkIOe8XQ44zHj9u8/hUUpqN4/Iu
I+RVjtsQpxUfY8O3jed30Y7kImGLle8MGF+SDgHvcEKqSvZFB/qiuCTRTmAB2s3C
c/SG7UjF6UJr24mIWyfxyIKobpVBUFQP17zfTBZfSuTdxn5di9Szf3RirZWkDcAJ
2OC7yldwOleU9cs0sLCKnHXuuhkAA/WZ+Le0qBbhliQgflC/dwdusdFC5cM6fJds
yCkRD1UsZhdimfhTWm55jyEKul2E2WoeWBRLDfdYxhPeeyDI1oW9+1kOdA5p8tRm
2emJoAYUdyD8+BSgFJNv7IkmTBhZlMu1D9erYCKWZmpF9+69ISuTSKm+Bs1ahEdI
6gfSaBIm9UZ/QOTMzRnv+X2fde5kELDfiuDVz2YIhMb6nmtve6cywy7njpu2Njkf
NFA3uI1hFtBKvQfb3GTBtUeJEHb5Jnq+p5YbDGJBSRGMG27Hl3lTgWPfliHboCke
+kYuIS7qyQNRq5kQ5RCNSddnlIMaMyVpNIyaGV27sOftkR2+kqgZBCe4Zk/Z+H4+
IKExO7Tm/1uNL5Ln7x/3YPEODJ5sqOARsWtHOcI924AQYWs7FSYg/YXRxeiSBfqw
GX8ND2p6MTKeE5mRBBQd+gL9vQHVovJSSQTIQxfnVy2gxnyOhDMmbGUS9Tuu4m4W
tU8s2G2KLaPU2U42ocGU1xRfQCV1b6ixQo5e8i2oaWPFsdI7XurCh5wyWRAk9oFc
SDPtqOVBT2yVBUZbu+P3GSDg871zQYKas2olPP+nCI/z1UVxgdD2ijVve18Ynz0G
MUHqGfn7tYEmtHZh48/CLjiZ+FDkWOmjqiqgCEA7VECsbpLIkRrioVNYZeJ3oIfg
TfwoeQxi3S2uvVi9WoSpbgS5hHdxqXfUV4dy9h5UwLHde9XUoei2h7coDBZMySn7
ne7uLn428hXxLG7OzBIq8brBsknY/rPLq83I+xeX4FNfKLzH2Kgt+oU7MkCfT5FO
Yxm4ZzGOAY3BuGLKIKSPQ2kuyYLQfdT9v80zMtltsSLvdvGhh44jo9e2CJ9Rfjr7
yCXEt920nzDxp00JxmbZ2tenCQi9KiOBDfp0ZCExGhMBCAJ5s2+uj80SDfpITo1O
LadP7pnwwMTFGyJX/EeneGP8VW2rw7z9Boa0iJmmh83igyUwar0DPqfj1/VtZDkM
G7owDbIMoYws7c2bgEsVgDetzAcomos4K2HzhrycAW77f5X1VX514t1dm0MKoQBa
YahxfvtOV06u2Tgi8SPmLAfC3GeVtNNwFjRkjgNfb2CuIs9JjGimuAFJ+tht35Jy
BoZgkj6a3E7bsFFNpAQE4HLr4+LfLmdDcMKwHfugHg4Y6Xjy3Chqh1X4/zCIgQM7
utvyGOQbkuSqAz/4knq3hDqwnmF89/yde+7dQ1l/ifo/TBEg2nE3t8jQM4BX6NkO
90PXC5O/qMp51tQWFKSXbP9pORW/iQxk8vNLykVSqLMSRDA8QYAvP/g/XSoi5kUH
xDOoYCfwBBVPHWIY2HRAycisJtqxrBoCqYPk7Riok04P/kxiFaFjSWBsklTX8ocn
HRATLWOUP42eOC2TiFdeqmfXWBlHiROaBRwuaG0iaFIG3P8OEQbyVpUKQ6Fp5sH9
9TjJQH6EA39URsUPsK1LvVgyN66+XSTrBN6rlwtb1OMur8+C3Xp02UNE0Obh9E+s
Qg2e7AGxaQtaqPZChkZMLdAx5leX5eK4tA71t99CAk3YL7fOXtTHUb+BWgOVVEWz
VHALXf28dbH8TVMHl1VExI18s2eCrAFm+0iLJkMZVGgDzT42JLO6oipWzNnYwDCK
yxaJ3r4y9wxj6xoWfz6/7fJzi5O7nWkOVfE0T3VWZRuiHtXvhVbjxRCqsbMEb4cb
y1b6RML8Uu8Yr4Aj29LW2rXjyCl8KIr4Jy9PpCBiJdp6f/SeipmB4fmjh1Urdthy
hrDMH1MQsV4CL9AnwujXiTI/b0OyDfIsDJU3KgU6RarOvJX8adj1f3ttW7PvzppV
yKrX+vTlWaJKmfvKkd/Z8iEmY7+si0fZNl7RHtpAI4jaY9tNgnZLM8xYdtWAdTW7
FP4rTUoMHMrso0SjC+4r0hQeo4kzDyrCloGbvYz89OFxO+l5dJKTwQraVmELbxIN
5HCh8FppIZXR1GBM0konuJcASuzphfD56q4sKePD1syU1crGROQJYBam61bOvJ8B
9cqOUStsvcNd/9w5iujQIcUU4h6fuyiH9psmaogG/WEPNb1PhDVn8YaOj5SG9aHK
gu6HIKPdFxDb2pZzPrZVLWnHVA4ZEiKGLobUHMVjX0OvavNIXxBjMD15DTO8zO8/
QSDN1p9T4r9KlzPNxbCdy4LbjnoPGkGzRKh1xPfJEriHzrzeNnRyXC2MCeB8DoKJ
Cuj0c7E9bQdSQQelFGgK71uWzRGXkgX7FgBnjl64uFxVeKfJ0aFjp5bwiLV/gfU6
x86Dab+vDFHDreYUCKwFQu11iJh/CXsv3STQaIHoInvoMEKqN+dKUZSJm4e/ioFB
0xYEu4aCNsYr4gzo48i5c/Z9Cg961k4av6NZ9DHXdc1mhzngFinPViGyy7AEzG1v
OW6p1bOYEwtMjJ8w4PnIB8B+oAA9NdAuDUZuf55I9vHbzi6mqPVHqOhPWhdrjUmO
enFf00xW142jN340a2P7XgqgC2DhsS/bQ+lazru/TFXCfj667IUCyF0em4c1cnyY
SyYm7Up4c+t2Z1NhumxCW2lx5doyc1hF2qKD4RyUhAekhzmY0+LXTsr4WTSKmSTQ
CGDVBVYQfKSxkkCpwjYdq7PiKwrJhN55+q+scjlqzdfPT+up1wacSAp2nYhae3ZW
4IJEyNqacIMdK8iy/PpfIS4XOJXc1vcG96ryyns7lfFW0XcThclxmwrhP5WOFu7C
J7Q1r2uhcVeNXD8UvGyRCQFVjmwto0I02ljhRj7kJEi+D/GhNgBalEku+yv7NlsT
OOxMfA+XgWxFzUwjEcGSQos7JP0cq+PiIwQoOo4VmKUIhl2pAinIOsAYydIVIx8D
+P6lo1ukOAT9YU90KmlIUAScFpv2n6Rux084k3CKbjHkLtTrElEj47slzkEvgHA8
ds7zYiVrL+aaiOWy7RPt6pU2WJP0M0vPVgsLVU6/TJCNjaS/1YtFPpp81+4piY9b
PGCYdVk+O6U8Bg3kFugAkR8yRTFpjuCWynDS/6oDrXH1nRWc63v9AYtzNQBQCgmd
B3BrljyEYfklJwtS6z+ZrXjQu/qiQnWng8DmD649hAp1NCfugIkDdj54dFSxdx0n
z201AwBAoeRXxRj49/gBHtZtpMxZpcigoSf9Pze6MHA+Iv4A+lkqPwxz8leD6wY/
aL/Drb3+vwHfXmBfE6JEocWFdQQC+UbPp4MQu0zwzLz0By+klKa2ROlB5Knp4bW5
08tbis0bJHNozylwQHyDTBzRi2ide+mZp3v3tdtdIEd7irfpWILD6Pg8Ku0x4haN
5Th9SoBst+dmj4M/Kn02UI4e1rnWao6I+U4A3RaEy7Y+yPdGHIK9IrwfCwpE8CEt
I087fmh0UZXtGibIRttoA3zl349/xYcsnItViNHf+LqaUhNQQLi8Ix110sjJTXgt
RaNaKJQXl2mbDjYhVUtDdRhd1xFLkCDl+HY0y6qrh/n24HGypEOzmS/yG/NQDvbK
rgfsEs0HMN6+wIHmMbW8+LD3aqxVXEzsWCX2/ETWeJpb4mi5JeiNVQmBGiLqfPfl
1BoMieUEcWNO989gqaPYJAZ0FaOpnD8+GV7zM7yiA1rrv7RozJ7lsZIDyejzz0xp
Bnxx59Ww9jRq5Zz93lsBP7WTUYVnOyDGmmQHHO9wyfd807vM8debvzGfLxZF+FmE
jaoUl51ufV4jmdcHi99/3oNIUl2lbbTzgcxCJnm2QJ+GLVelEhL/tjynXXbPeDFF
AGd/fDT9jabibRH7O9rt+je3yC5VAuRegyX3JgSOf2wO430zwrkl7o2hrWTCCr8v
IwF8LmiifDamKHr9XUUZMqyqg2j3meZGwR7IPCso41hw6azQRlDL08HTgYWoLV84
ZN4VwBwFGexR2Dw3zIn8ImCR1iC92ULyKRP+z9dcNaEUCKFuPEijq0u4n5kEvP7j
JU3BqPFiuYeCLF9Ed4ybjiznQTCZxRBJ5w00/QJypnq5eWYu3pDfwQ5hDMSmWcZQ
TvcU88zRqAXM/gJg/RAobXm1r1Gjnl6UqXaEa5WlMBgJ385IMUIDq8mRtQU9TirH
4hW3+xoWRfjny9F3rgzBORstkRNKSR36eJ6p3JhlKtrtDrXEUuw/6bLdlJ0p8tl0
L5tDtCNWNj43o/bIZ7k4BPt/ADS3sJ1Ff1irQAoMSxLbJYN7142wZpDG47vnCHwF
i79tNefYdl82hvG1Ys95KP73aEne5Fh/N4Z1CQjlde9ulyI0r8ivoIjEUurW0pVz
DwqLIP5mnfI6Wsd9Ysprn81hDHOcAfI4pWzjY3t3xeLd7iW3AsvVpX0Umdv5LYFL
MRqxAdZckSVfAtQtmXYb/crDrP1Ux0KFGn7T38kl/8Rbi7BeYrQsSD3BbpkORDFg
K5a0fJLzouUGEB8+cxStXoHuiuMXio0zyjRHxZj8r6iPJOxxs+tHt1IbRKcCV39L
eOo4yf3v3GJQup8IxokzTH8XUNdTCIhIoiKW0bR6jTdj24VQYGBS2sjhrdX71dsj
Cnzw+0Uw1O8J786M1G+lQC9gCGaqU5RFFh+X3+hddTwoO2nE0ya7MJy4yUMMf5UL
3iXx/c0a7DuPK203dzVuczT7ENORoNVuof6QRwlOUr3vhjlysbKWFb8MvNO7llar
hx1J2mpwRV6AAKN5pLYWbvxyyO3f4eNGDH16TsO5U/GwTjAv5Ux4uGp9TxmwV/0M
X7+8iC1VQoG28Qaqt0O6VrKo940D5PmiguIorO7m5c4zfi/Jnp7qlDkXMCUFXg3x
Ns3z+sImOiAsLhw0/dY6YCMxxJZXm3mGrEPyiXMoarCtTRMQD9x/MdVuSRDY9sLD
nMWuakvScWwufRnDM6RoqmLtM4RYr/0Fwyjv9RmgmSnRS9lcmUOia6qBGxoaa+0Q
tVWHSLwFU19b++qhL4Gk4/Y3tDgO2TzCPfhn9aaoaDU6vuzSh3jgqGrqttd8z8/g
Xx+AkAWtXkKzyIQRQZCNAYaM4QM53rFIrb/YSykoui4L+eCz4iF/7uEuCV0NV/lM
oUzOxwIBh4/NQDFYv53uAsE2Rq1B/cebphM7pyVqaBAkoHNz8r2SwLQlM8QNNwrP
+NTGsz+cXVVc0TK9j6K0QBODNj+vtLt8j6SLpPuEoxLahlR8yKIPuTeqqP64Ewo7
ePQr1Yv4CwREsJGiGKEQmo07xTRfnvVAdyDmDT7u7Fm2HvQRvdY96sJZ4jWP/wgN
q0VgZoZVIs0DwfqzCrMEt0YzbjDmTiN0MyZygpjZwMaKOZ4qsN7xqeG9EpNFHScv
4hEWPUOzY9BeVBGXv8l89wpLii11txiZOEVeDK0W7NAATVaEOq9ZRVOQqDS+IqzG
ZCETwspnMLKEffcDfTqXcxUfzQDBtRPYPlc5bDIvwdNJ5JWlkR858JHDmbi3KVOo
lKQIzysPVgoxJ2C2K5L04ZJEPzF+mw5aToLHTT4hhiOlxOzd1EwSkr/nxan8WQnu
h8FFnN1YyIp0GlWqoHi2SWH2fgwyd5nWK43/tRn2AsIJJLqfuUXyAlMbkBZ+vW+B
BGuG6Os4kxl7JOVuK3UA1pwhTEW9EzNTeljkQW/5cge+T4TUmkrvExu4gqqyauUb
J085zVZRqgH1ORfscu6cCWmL2T9gNEipvdvhBnloxxEz6FBEoMkKAxjxbcLkSKig
Ncy19xjvsLhpzKG3gUj4bo1S8MYwlmS+IwjfkoAV6CUff7FzEdU9HR68rjazZnDs
ukQ2XnZbAQfTcEI2h6j6yhxsnQRgk6PErVhShit0HEXowPLKwxKdfiuxD9C5uP73
eupGE08HZQQ+sDsRy2GsX0ul9+Q4bhuSW6WhOHodn7X47YFVDQPjMTzC+HO6bF4o
Ggbu5Y8q3wliT6Ui5apn38u9rKEG5aljS9OrKKVMXDFxj+1+2eh/8dLiCM+fzxla
f31+EXit21L4FTODeZT6ARhgqQixLiFvXdrXjiS7uSEj9EVoilRhb1Yy3+F4wwka
thPH8RWDxUbmFJuUQLzzpUyIdfrLgghwMgilVhI5TbfRRGzERxnO2CPUdgp6/Ou6
2KTmPXkGrpVWn5/sNWi1C7mv60T5VsWA2OI0Csud8m9I5xPM5EGnJmMwPGUs6xEI
3JPa1yciR30zuTXSAFbKdXq86gh6ggA5i2wU5/9YjrYOSlfmSjWPYh8RC6R+LBun
o3QBF0KZNPVV6ZiFSbJB+Pbt6rX9lulUWZ31WRpdMIcLU5H6EbWfrMgnS1+jNCST
JEoJTJDiuWoJgZ6EAaWcD0bFFCjZVbQMWs+LVY5INqjaTCzCxnGiQLpBgyJC3J3c
7Yvtabyt5+zn7fEZVdVGLoMfdaKz1n/R1M+HuuicrJzS9pN9B/v1OlRnhcTaovfW
HK81CSuCwr0vuolWy8uKOk/KrQHO9aLV5rcrHGWDGT+Ji98DqlbJkJOniSXRNwR7
UXMrvb7bDjBV60zUXI7YOgmTJVVyGYhH9CCNORTvxhzYFPpmJ6H7iOOGYeh80xDU
M8ZYOITOneShcsBq0ZROM0try3HaelL30A4jtrW8JkMFywzY06a9T2DnnCrXc5HJ
zfaru4R3fBfew2wtGas51tYV4F5wBD4haP9HOBAA4yEp1ZUYRrKTNJFuwTchhPmd
xv38sks+AzosRabOoYZWYd67Gr+gj03N4HYhcASBy4nugK4QQlwEcol/WQjPfhg+
PSdPkChs9tbpbF1bQ1TDXryGlnQ5l23FFJvXi0JNVQxvKEAm/xsuf6DdnhRuaS5w
LorL7WSimY/+E6j+UMlFp8ufCGv1VEj/wBa9WUVtJeibx15yAymezr0TvfJFqqNn
6DoEqLH3JsInmGKQaclXHTrNNmWp0zXxpJomnE5lIiMBt3aYP8SdqmHzi/30H+m9
ck6z2/IBB+QXud3+fgP80NrdxOmhTaXMoSMrqKdfJwANCQMfgakMT3lcY2ju0jNP
/eOcJ6j281Jje52AyxnZiPgZWzJFXxOTqPyj+nLIYmt2gcIb2DcYsN+cihxP3W7Y
n3ByTdxJD0fMJW5Zr8B8XT15pW30Jv9NGuZW7DWfZUrVO/hfG1x/Qcfg3sW6Ag2P
W13UQiM6ySy7+ExlqHxut7w4RM2NoXW8SwL/TJMVGjXc9xYa/4RftPVtk0aKXqjy
l/aIZ3UAsUGO+YcZp7WzQYTgCd7R/TG9YcPF52p6gtP00mky9qKun9ZeX2wmkn30
v9BIy8mU4nGOdBdCmohlyV+eEDj4LpT0YTCByijw/8RCXN9NJySmZVz/LlPAAUfp
33gMXO4sS3I/jou6ZBWlKzt6F6PdiPd6anEZwbmQmui068ggBi7r60ZKnfxHNZ+a
B54EzNCTeHsasr3irDMD+0gEqLdNlaw8LYpx6/ul2/8bNHj4GAWxE+5/4z1O3MMb
FsjtEqo+aM+hGyHoIfaRxOwEWsKUqueiVavr2ohm15QXdm1Jlf7T0+vS69+mn7pr
2AV0/eUGBajkjYwfwKCpkvHBrVMpcnVMa3FyErlcINfRFW5R0gSBQFCC46LWYv5r
L1V5dZjx2lkafSGP3M8jgf2htRwbNaIX7c6S/Nmo/nGayMoCZpDTaFb2/Q4sANYk
3lsw8OcNq2etc32xJTI4iyeRFQx5cebBkrRnVtYiFa5Oxj+D4RCsofb6h1I8Hx16
86eSWIaBoYKykJsWkExK7Lpgoxvn+7iSSoEtyetTl6XNknB+AKkjJA36w5z1Bije
7WaLukDI5h7Lx8MaYFUV8MNdxU2ZmjoKsaeN4m1p9gBuamoVbVvQqhzohNi7D06t
pL6ctyhKmu73Yf4jTB42DgUXRqA8Q1J2OTKI6sIIhnr+eHEu4w6SQLPWeD8EV1iZ
Lma8eOHbGTDUnWBqdOz67qEE9dmjSHPy5uvbfUVXT42g79MjTeKiPGt+IrYGOAHA
UfJPzlLEiTJzsYo7/BBisurVQtBOobFc/gyBD5SinrSKXshPM7/G9i63aSfXod8u
FPVaUl0OSJaw4g1kzLzoEGbMCBGHRCL7gs0xfUgFusNUgTOWNJWMIKSTjzZG1mNw
4fPjTdTk5Waup4Pdp2rNz/V9X+pzspQhQr9ljpir59GtMQQqvyA53jHQxzlhVpaI
GRWx8EJzZA36yr6sCxFdA6TBKTGHMB2IXsMt3wlINGl84l1cJGwj6iTVjHcIzm/G
PWr9cCjw52R/xv6jUJCuyrPY67AOo5iOPmdyjxXeVz4TbGoyMQwfg19DSB5fRyOc
2faU6rtOG7n2jk76xjVos37AYMLH+uy5Lmwks0AYa23irBMsLpiUnJSIGTAPQ5jH
/kJMNlCcWf7SiGPP4KN2uEO8VH2bZ0vavhe0/Fda8gfMOrtgrKJSnVmIWT2FUZRL
Xgq3/tcIYdTO2UmSwOqm6um2oOy+wQXfK8Dk7vvFK4193swcBbBnNjJZLFUXKK/k
zg8v5XvZMzd06+SmLNFPi72OYf7OM/pUAttmNKAXYgrqrJz7FsX+gENCl5rn97gX
YatvUTgS00p783lrpuVL/0upSKjwqKJZaUwGI+JwmePn9/Zu1Ra8dah/Gx82BhGD
QkI48iTmeM+vTKF/s8/rzUnIU1uoHOvbmEsr0/D6DuPfiLPe9nHa00x3QnYvbf+W
/7jodTNAXGb+/yG1C7u5+atskmNfWDwssR8iYilh23m/w0CzTJmdE3IESKECD6ow
hXS0BlI576TUx58KAxXsp6LAwukhZs/6eGhgd1NQ4bxlf5yF+0XXj41+0z7pF0EV
UIasOoYmYqixFrp59eIFRYb1+4I0KcN0S4luU8PjGlQJDFGpdVr18s5+ONyo6OZ+
N5ZIoBgGaTqt7RgOvxDccsZ3cbyu0uU+3Ix+AD6IHfSd6kWF5rYrT9ku+xqT0+fX
NIFANAwpV3tCh+mLmYqPMcC96aGpGKstz2yD/tjo1ksFM2k2ekDm7BzkjUuYHWiZ
DTiXw9a7OYappVXh/r9yqKyIAd36X+E2rglWMEfMqVNgpFdeaXTmY0839x/Q8mjp
SAsP2QZaA3yUMYrZVjuOkqbzOfzS0yRBjAy/9IB1OUIAGaGXOjjjuB8gnAdd3eM/
nmOeDzJEF80LdUr8tL1OWWqTVYEBFsALdLVAlB9D+nq2q30Pp+PL3/SWah7/HCsC
e3E5Qf0SYDtglo1kc4FNIjf2S2wxzTdMUemtF3bc80VM5RKZF94S9fnW3rGjOWKo
mPAGOvtjAzOO3nrvQQJog0tKJ/d286Sx3d+EU/nE739Gn/yjuXZtjqVj5jV9/emG
9Sbt6dy1oliC0yHf2a7QdKa2Cwu399rfzr29MaU1Tx5z2NvBu/O6FINq1BJNR4W1
TE/5LBE6Bz4XdZbqSgnSeTazf0QFsV2+7pslKSh0oT72qBNPJSFlgxLl36JtALCH
DS+0tQfD61nk5q1/7NHwx2A8zAVquPiyVHMeOtuP7HaeRyOK9+N9oKO7cZHz2ru3
KjHpdPIjBHeTC5Fcd3zTInmPj3PRIhYRzz0FOgp6Ssc/i6X/DHJx4/1O78wl9dlJ
eIWHEh1tWbgHwDk8FO1hVhDOFCqCfgZxWqUhEp3eStV7Y6eZRpvV/3BobiDLmjDi
NP7bwNbwfVSbJJT+q/ygXvAV6OpiieAQ3bcaY/eUPjswiNNj9f/SvmuMBba+35Kx
PasGU636Z+beihwp2xddSOuSdECWCO7g12OWO6lBPGgaBBCu6bCWIi/sCLnfrLT8
jpueg3QcMX+THS9mQjXsaCrxp5LaAAmH+zia9uHPWRJSXHURWrEm0Ay1njVobCyq
MTb3vYqkNBZJAuQBN685HYYAFtBNwHF9sSLpFzHMZQ2+SDYKSyVySC5u3fXzHDfJ
j8DQd+iSYb6L/S7G83/xZOUKAml2ggReRW8Jf3YRYD0U/VkE1r2CvOWLW5xmGqBW
eBUYM+7jWRw2sbwmPo368DaByPxMhLQjZDIcsfEfPYlk29J+AJbzNnA28734fLlu
RUWAvUcJiAdOp8LERyxGX5a6uK09wUBl7lZuHAhBb3BfHkND05rkG4e7pt8+1yiJ
s8p2bcXkJdL0fXe8LtMs4GeWZxyqjLX3rNtIXrGTAzkJD2bRvUa8Vke2ZvlKTeGN
uas10PLekY+gLlkcR+WwOKCPKzh9chZcgK2itoOa6h5RBEjyBbjkC7vTR+pmoKGv
USe+zbu/qfXaHdeQFnefOXyufhTu0TkZGG0lQmacMQdOjAATAaoJrodmps5+TJzc
kzk2JMgFockkCqfbKnRnbJnaCNnU4Hh0jRsNOEDEFE9IRlZF8hSzmBJsMs+mkhh5
DF2eEh8ywKY2KA6sFqwtIyT/2Y9P1aJnWHtqTP5WZMMSIm1073QTMZirXgVPLEgS
Odzr1cvtYq0863OAWeEK/7EkLlnfOfRnRdrVBRFTJBCmD+nH0NMNzEP5DYj9JQTE
fWsdr1qWJxbfe/nTtY/Sax7IepuNfMzXwa7qA2reE3Jn/2OgaaXwWtXVpN6CESi+
vueJBc31JIZTQDYEhrje6r/oTyAO/f/G1X+3TXFRAPG3Won0eNE8C9IY+zKHIoLo
9YdtIqcVzsSFsXi0GY8duO8RqTYuObWNH8+VkPvU9dTOniIeuUVS/9pEcUVEuidV
gL1qjOEzGAoRoT73ikNC6HsYHp92W8+Te0lY5hmsIPcZjNLPi2qMvOEl+beYn9pJ
M2m0bK7TOdG6nSjdlwxBlgyZOQ7qIonPNjQ3lfHwJCbwGLvLwgXmm5oGhwYFEFwL
F2b/a3mANqoBRRIXxqUWltaSGu9TFV37eVCfHn6r3vzEYOivXHkq69tGglherBz3
SbReQAslOijVjgHwvwgJ31awBOxNXecQ4uUBYQz5nxRez1atQE6pskEXbBcnR0IZ
JqC8S+gw9jb/LFkyckHzpadRXkOWkD8zQqZwSn3e3jU8OgDOsUFJE3b9buqg6IQy
6JjGmMjAJO3Tg9xDtgoxJt1tueSyrDyA6eXR3kzFuksNImrsdFzbnBJ93hLFPSvi
GsUwniF6SzMIqDx3BBjdwB51ECc888W/40gVa4fcCD20iPa7VkEc3cEAqZgTSKaG
sjmSQkFitWc/WYrT54GBZTn+NbILL/OGl/sPQ+3C2o6DMR2w2o7SU1PUQVN0lRdp
L5idRmtT6LNhOOxJTM2lqXDTmQZIFz3T3EcYQqJ5Ff1+5CjgzOrFrWMdKedEtjNH
veDs8ljqIuEMkBQUgHcfKIDbH1sn6pBInxExIYC3yKcqnJL7kY2ib12CjmMGNOlC
Ful3uADQ/o8l2wfWKrfM9T+TEvQxxQ0pC7oXQQIrMpv3kFbaU1wXcCOcTp/07Hqr
64G7adOTI4+chz4ZLjk+0JrXDSBlzgSNBTWYwFuPSzIUNGyVU/PYYvPT6zlbXE4n
x81PBYVO4y0Yel/9mcQKhtGki8gaJFOVZREH9FzKZQv+8onFvc8ZU/X+Vnn0OS5q
W9cjHAqGgVTUfvfE6CiK+8Yo1YMSZs0k75DHVjECLBLlIHmRz49QmV/0f6cKkUcQ
BlQDvYFoE0mco4s4WaMFcTBz+kMHciSpi2LEMvbuxkc/GwhDhHpuyMj7ikNdN7C2
sOH4jg8jrugfrfFRnKLNJwrj7I8SSZtUI0kqXPQ3oGxtqA5wf1pheWlCEzrQngSH
QEgPfuTRkZnIi6+LsiTBHSh050rnY0zLqU8+3w7kwoX0hwclBAxcRychwr8fG1Dp
A6Y4fSkrWD1XCVfbnVMco1QyPjSpIQ57JumAEDMuk8AbuUtET3jPEAskPty3kNMV
eFlTP+TtkLZWbowBjJHN8ABK1a5wV8TkVLl1kR9TsHIe+rKfkpCZ2yWBIrfI/GQu
PXo0kgHbnjkIo7ZPHwYJ0KfLoE9ELQ+A4mbDywcI74nT6dpmNdpyUjyalyHez+7g
bACKA+BRaR9PgvJxkqN621G+zC/Gzglz0pxJz/ZWKV18QxwCxOdfFpX0JnvjM0nb
VB/Wp2hhXC5JPZcJh5yepwmzyV0byID67QFPtXEfzsVa4rXq+39RVFEiXA2f3UcD
cusjjBN0/L4I429mUmtDO5JTEa5gPR2y+VVtoMz68kXUB2g25kNgesYAOBjC7KEC
3Dilf+ExODfE9DaV+eewoZbifmYAKarAAHY2vamdFCZMcnaTDeFmJQkwpRonORDr
wWdcmTeBnLmmZhAdZrIF9gvjwtIrWXxEvXAw2KBSyNFdQhj5jmrfgFRB8nL6Wmkn
NH9kieutfj6mliT1h4jo46chKiuap/A/McPjXVo9XuHv/MY00zfu3M2d+3/G5uyh
ZuFgeZ9ydwCAjYJz+Id3M4eeR+c1tkYYtZJV85zPFrNgKHxnrtxu64XjOJ+wCuD6
HicPhelLzDuUmOEOjX8L4evA2YfYr3DkruoZoI+hbGVWE36zOpGa2vqhPkrOA0tA
WqLuUN6knZMxcl9kPinsackjJrInvhPaUbDQVC8xBMLR6472SJ51H5Js5v3Agwpr
fWHK3a5mdWxl24UQDXAZdYXkrDIO6vR079XliWsvUxluSgcRWGiECEfoK6i4FazY
HW6Wjfe316N5zN052nceTVVeDecoU6zWV1RgmTZxzyW5cR4PVflAObgTEoh5HmNb
Qzib3y6DUP2506htuND3wmriKqKPTXdTroxYPiL8aG6k/aSUNJ4vFqIvnd09Z2/V
4n11ZfVb93jLTI36aVLtCCSveXosg2xsoUKT29u/QKqjJJfMCoHJ8JmPiZ5Z3euG
ql9hzol+LtwTucIaVw3ia4+UdGcoJC5QRQP3FQsXNIEB3nkZE31H/yq56sZ5ASHB
aUBatEWfyoUUeo46A162XnkleBrgPgsdo+UIX+jv9ye/1/GrBsablT11IM0S2cjM
z+42qteaP/9mPV+VyoCUjH4H7varb4AOxVRMnCoy+n/99OkIyelbCTLLKxOu49xk
lx7GrewQeAJjjj78syYWqMqzu8m41x9NLKcKRC9uH72ZJS/zssWNem+UVOkbKxXb
JUrSdC5Q2UJ6eA5E0KG93rvX488QsG1PwyU68teWNzm5wTVCcINpjg4ARc2yVa7X
4TT4M/YxDObKhYP/0pMqwL3yq79+XaeqcXkcasqtmFnEtALCnse0hNvdS1lQeM6H
/KFV6ELZeqlnoZ2zcMFGZjkmgU309C/vj3UMMRG9rD3vexuy8v0L/87qFgfCNQ32
jeLgBpJydLUhW/UsVWpG/hLAsSz0j4vgbOiA4+9cfOk/2UTNCh1ITZeUqxCRWLYt
GEvbgLXUskRknBHw/Ej48Efd5QB2g/lxSEJuWgNgFjXvqorlkqV6r7L0JRpzXhKE
Pw4BKf6HtsBGh2DwWyzXf7+RLEg+ZqoV4RFgDN2UutdB8z+J8M11k0qd/+TesPPp
YeYFXk5I1h+aWitQTzr6OE6gLzqpPJzGjrbL2RfMm2SnQ4Ee/O+/fUu/alp+AD4e
wKW7beo1UjkG7ESuXpkF0n7aOns8li/lAsewkM9YrxsMa1jyV6jwL1JDFpXbNjWH
sJdLQLT5s+IjAAdJua0KiJQIGrgleFK39L9PQpgGKNhzeXPYOgj+Cd1scTyvTPeO
6KHmyBV9QD89xHdlsCu+DCiYiEL1qd0C/rdY+hNWGhnpkaTHhxWtjUd8/RqlBBwx
Ymie9ZJGmOuUTUNrRWS1HfLky3yOU3r6wmUybGvArp9yGGEkR43jfCVwJ0iZwY9l
5Y/joMXXc5HBW0Yz6tnNyp0ZV13ROsUmsHcypoMntXp3wR1gcmAY6Be3Xp/9Ov7C
PxnELhkakgqWtb8njGWon1StrMGk7v3w3qQl43Y/+Vhd8urEgZFVndZPNbn1LlWd
JDwyvjt/c9LGl5jHhBFQvn7n88R1EwZO4Hp1i/ABWnG1ZmR/ELbNFg0AgRuNmabs
gDgmqeXTDEe8ti9V/WkUIi4qwLPmEoDujEbaR7b3W09u1wPp7sdi7BkmEln3xV3g
hGYA1GLB/WSzrQllI69O4FU7cdeipJa1cCyWeRhbQW4iX98KFEEPUr5RsWAbelNq
6C8FpvvbobqAe75X1YXypQfDKCjcQ0euG/B5bE3cxWeqFGcTNAG2sjIZlegzm1g0
srI40gtem1C1FQjq/Qv55FbjuI8Y8EAyVON0o1md1pcuBNb52jSf6zWU7pO+u43n
rXz3Y6eCyJBwxHN6+rFvBINJhL8gK4LcUmOu2MC2a1ZSOXOI338bQrHcx9mWwLiX
Eqfkqrql87vR4r0yklvbnXoDK7tUvghV31x6wSfGJujEHvoClD86u5MQVc84D1TU
Ba85kO+3iHVUugs2MPj+rroH+ISKbxk3z4yHt0GUTbIjZJL8rcc5y/42JqYctS0K
c7C5pTog4yrMkgh5YmQjhGghXuysQFJ/nFJeStKmJ4gHqEaffgXt6MSUGfWcSkct
iwqgDmfrutttK/Y2abDGnNgQkwJqBFZTyQ+rYfx344o/iYhlPvLFAjUyCE+0jLfJ
iVU3EyqXIz/oqC6wVErlxggimZeXUCf/46uoKH/1kpuI+5PIQOt744Cd7nZ8azIU
4TSqpnFFWnIm6pGPesgZ2OvTuSklBT+4EHfLD4sD9dUPz1sunyuuCEEmeq5WyIIN
ObetZXZPHIRhFbBhaAqfWHPkmD8rkNy71CFsftaoqmWShYOS9B3ME9USBxjIkVEB
OdcmamHHA/pes3QG4qtwa75qjKYDi4ZVMolZAHeC6q/1mGJ759JRiqJIYV9tPSi7
Bv7Fc7TpksppFtSV5bPu96F7YAVSqXBWAk0c0Ka4Fmfimox7QbKoi8ZeKBn/O/B2
5IIc4d+IlRFk673K1cwTu9DaLcnlqlRCAfjpaHgJsLfvmBv90rbe1ZfWx9N4enjd
Ks1hegUjYKS5RR4bs0bz+hcWRj6uDJeprP355hr/6OpgxPHinEsZ1Mf/qziWHpDL
bKLqNtVwRxN5WrMNTyIhQXH27+fGhmYPFQ8qTqQBb97Hdv0xTSHQFmqTbuikcvco
9GhugpieAoJptMxogNX+Y7OeXZfNCE5+nbtopMZ++nxn62Sv/zLBXtAYdcBRQlvh
xs+4gg6R97aMxQWZfA21+Sv6ZL4Rnme2JAQuVzyqf9OvuCzEfb8S/bD7L1jL3lFt
9O4ITlYTjgT4bDuUy0lKVV8idfXHD9r1zucxRt0VZ+PQAHOc5CgCtRU2VrYrrRMi
92Uqn8IaA6oXgrq2KvWLzFv8TwDqeWLbZnHXVyTGcL0E1VQaWi7XU1VW8gasV62Z
yWqxHE7r04pPlhUUbHjAtbWIsFwhprZVSm0SAmCN4R9SL6oeA/cVTsDjFqHMTQN2
jSX7sgDVVJ+gjW08Fpbkfr3i9FQQ8AQ9S7YS/msArH8Cxlp50mRAKJo/Qj0Pecfw
i1XOBvcSUcvTsJhPeeUmGBS0o/sR6b7lZfnBAfsoXgGTKrr+zS1sgLVDs1P/GtqG
Q6qua2osGI1V4e7W3oP/QdA2YjovnjXJ3ANC+3gNVvvK2tKuHcvbPDvIZtEQbi9l
sJkst9eKAPbBVhw1fG3LvQYceYhCc9AhaowyJnF8qsO2jEIMVemTxCgXhwKHJ1qR
CJvCV2VhtJGe9WYGnZDPsEbFgHofpjvwcv4CLh6FZtIqseJ+SVNEASyVr85b/x+C
mkKSRZ2Eo8Da0Hx2OjvuNEbbV6oPxmxrjvSNFF9oHS7oiaXcYy9OBIMfQUbpyjLE
9BPrxwv9lJXPBt7ZqCawY+DZx6tY7gdO94FuDpUMkV3dJk/fCcBBYdINnWFHsEuh
2SfxI7xMwGi87CM1GfiYlAsfSnM3cH24yAwOanBYAcELaKJPw6NmT1ON887XmTnD
q82xC4cjyQtincIXOOA7Ehtmz8flHCWzaS78/P9caEjsdNb+K+pOmB8CN/8HraHr
Cnwe7QQkxkDLbVpkhAuvogTBskAHfpD3LzYbKZzuglq+zrGGrjXHUHWuHwE8z3vx
zLeioAPrDIb1UFaW444EB4ztShuzWwrRsfrZIjI3PiWQEECEuqW9GV8VsiAIxZrf
wwtVJdTx4CJGOOTRt/gzasHVwYI7kByh4aqlV13ES/kl6U7/PvcEBojRI4VFuVZ7
OpYw9YSs7BshLM6gXRvu5/cOjs2UehLo/BML9OC3aU0ksNEkO+tL6r9djvSgfzbp
EUyPXvbFmScQ/4RJeQ7PgNMXNFETcZyL6fHFlbfmuGvmJ+YVu+zL08K/pruCA8w6
BkJzhdvQrh3/4yvQ+G4q6BqF47NR8sW7M4LcDU1WcSF4pumKpzA6pO4oiaba1f0f
qEkQwdcuGzkrnNEaxCPEgELw/nBr3tUJIOXZe0VwJlHwGLbwvhVW4jDtXrcvCQbL
WEBeSDZNfZNMEcjxnTNM/B+TPjfi66ehn0GkcC4HzsIZomaUrd6WXD1mzDaQy0K2
zU+xRuktfc1Im+fBbGncq5uNCitBjFtOsVXpmXhBIhufInOXVj5fTHKs5d6nm9l0
TYnhYi1jJmCQ6YQwAt9uMzMHVRYKhhPYxJSK0LMSkbRNN9xWAL0uIULT5gif20PJ
eQrY7GxPk8VPq+LwdqcHnHeEO7AjMNyKEsECScFvvq3EhSc2tfzvKWmRf1zakCjZ
uQD18DwklEI4FpPqOww34XOavO8js33sn3K3xyMY7K26trCwbAQjlWQ6fyDikzOn
7sfnPX5Pyskwu04BH0hFcWFH2Yyi34xHXofyJ0meECi57qFuD0CQw9A98r9xZbtE
3kMmV8U3IXS0xirr6LAogMBfiRRsVvIePpbrKnQ/8XG2mExUjCVoZ1UERngXA4hJ
SfMIj6R/DEhV7cS8m8+YFTua4ptMICJGIHQRnM1NscQUz0RWBPGKNDpokGA6qvMF
urMF1IioZ1EvVIjg5lsTxGHa/TIH3NMIdjQSj8KYPUY28wGdkKPLxITbMQhXESM6
O+w9FN0nQmhZFCp6KVLAIavmvDiyULxFgx3uaw7cKibmoKgSKRt8KVFyzZ3PE8Je
NtKuiPEWg/ctAxPw9x4IHZHdksDYH5klJ3JkufItj3MkicXeTMVJYgeodhivdH0M
E2UT5UZs6uGvnjy0WceumYtDe79qxpG5stz0E/bbqmlmQ1YDPDeI8U2T9unECUD9
mGgTmCMBQeUh76kk9a+ucpEby2qpdScZPiwTMuly4wNlHciyk03CvpDNMk/77ZIH
lmkKWLTTHYkpf8MnxT6DEXQwsq2q5gq6oAei7Kmv+E6H5NFKwSHUO5wyU8thll/q
TiULA8GyVRtbMrwLl8cI7ZgkNXqhHPY+mPCaLb/N1jmASVA96oI9w4n7pmtIUTaW
zny7VzeRSqxVWXrjUZUJFfSOIiocdiGL50+6PVOCpMiuApFNXjglOC+TRYI0auuo
h2dtY1Cgm1BK+Eqi7mbe85ExLzWiUnJGXjt8c5GZIp13n5tpGUf1YZzjLBBxsuSB
XX+nGxoZIQGoYqEr1il6XTlEODiwm2/qzYLGaMzhIXKQjzlcikR5QXv8OvGSy/0Y
dCBEFSh34vZzk9TmPu0kuRtJfHM3EPlGeT2jpueG9Onn07kN/m6ay9nn1IjUyFT6
07fA+yCB3oQZPnjny/JZn2lWTzTYn9MBp0BIWFMcq22Tvz+owya0vRx7gZFYzEBD
443tPdMgNrqCmaXhkSy8KouajwSqgxKED8g0u8yiF/IWOoGNl4i1jzrYsKc3gRrk
NftF3QyBVOUJK0fLbUM85VQ7yJXtEZfZS7Fdl2u8z+bqQavwxADUzFQEDsM216vs
A4iiGz9gPP4F9AmxhCmScacjkXYbghfGGqk2wytcXrgkbnlnAuK3S739NCIDHg5D
pqcegDxw0nmT3NSSJwUGncDmf+HSEbZao6+9CpuFNOUiSSHTz8RjOZ5MsTQgoJO5
nXN9SZ2bu/B8ULr9UYTVAgRGQE5PVfpiS4d5uX68sAtFia3se29ltumTtgpBO6w4
92IYL7+FHY4vE7Ybxx4bqFw5LI0nHx82I4vFp8pcMUovbbj2g7m2mPFPkvxMU0Jf
Gm0NsOnRfaIFhQLHLWPJzHJ4UPcGKt0S85fueHbWOu1tX/wUi6ePKKPJgYI0WksN
xCzN+fsLU0DS2EbcpnQlq7RwqrRNw1AY9LO9DXWVQZ4xBPr0k85OFuOuIy9wro0X
7TIio3uO6K/EIjdVE894EsTAAsCBTl87hoWDplRGhn/TA0wkj8cOC05smRAV7bjQ
jUcQYFGqgeEbpehkuAzWd4b0L5PifiYLCO7V49WtuXAQcluTqg4nbPjErs6GPZfW
bJI87BFsnRofDm+YHa4iMjwrLc1GXnOCL6PA3oHYgJyzLMrzWberUJaEju8izEyb
lnM2JrqrxD3JU9ytyzTPbNH+jPQCz4IHIkb6YY+bfP3GbmeKxudG5bapY5iSF79c
epYOgtMxMN2ZE1qNNTMicCjtlcQNLDWRiheq1oFK0cHcmgH8jMUa+P/n3NgEe9g3
K4bINCUahXhToqrDZD1B3zkrV1TlpvXhy48hCqKEmV6c1+XismSJ2/dTRX6E75/a
JMluQD9naz9kxrl+NoH9mrSkVOjg0rnV95Ror9+ikKF1bz2nSRTc8HkcYq/L2CIX
/BoE7Ud4RedcHfB7Jw4EhN7RcbALpDIwEm9OLGN4Z9PJA6vFmTXEAprtESvfy8Md
xSVXHc89t8UnJ+6KBH53TKlXUJbf5Chxdbapm0n1jE0euKjyZv2bjTLXZFQvVvcJ
+UHfJT1eC1mkXeQI2gS/Yk7X4Rqey8NGFk2H0ZUmSUlXj+UP1gPjPrQWjvdhjg8P
Kn8IufLCVJaLE6sj0GUbBjz7RXXq56Zl0wmnO1Y6D+YK4ofY8TYS26hZLBHCOe4r
RhzfRX0VG2x/clNKCee9HlUTyx5pOmlmzyEBV9jvz5TWek7azhQgFDpdUL+ishXg
kzuwaamONeOQiePqcvt9nEO3Y0uCihOkaJS9pMb02XergMguit2Lga8yKKb6nsTV
qAa0HJtjmK8rL3EQqaEcXht+Y8KusNGs0HAIMBcuvFW2n+ZO/avUgWk4GUmBpyw6
7pVCHenpprhC0139MYnJ7ZndTqBOR1/HLr6bvPThBd/nZJvHPYZ04wMgrszTgZ4q
ZD7b4tq6cqcnutRCOGaljbuGmIclA+i42CVMQ/n0vMabJJUqrmYotylFKbZKcWsB
XDcJaQLGtXMyqfu/Czxxd0GPTxveXIViv32bFhwkOZklSqWjkgLu3XBV52z1g2Mz
UYmX+VQI/+Iz+pyPrgvg4NyaCWlCbi+WzANnyMhc+xLm2dVHVmQarU5FahbRi9bq
6J16EGYJ6dWT+566i/bD0NSXHtZI7yeFyC/LSzUmZqBK8hjrPBu2IHA7kOxiXrk0
reDKAWs+W4Q6SCDyj7Qkkgdvd7BK6G9p17Wt7ITKSMM3QhmX8IYYzG1xl31QifxH
OUELfD1HkYv/oBYD4fG2o3dMx8eqGWOmOEmwjX88Ru1ErXSqmJA4WYLUMNjgK50X
6gSpE/i0IOdC5fCz0FcKmPO/4TH4GgeEgPzpCfU1GUcYM2iHBCvkzf9242WdZ/6m
XrqcDzWZXId/ZggJBiS3DZmeSvXMNTyvZNHdNBJF8QJodD7UrR1yegyGYfi3xGJd
5/VvtHYKIuz83gTXSVPW5jECnD++4fC3VUqcmD0dTkKYeJ2QHthLdOz/44/pFKp6
Pv39AGVBbPSvD15qTHOlYkeiC1xoSrcbZv8DB9c/U2KZQQL2pP69Bo5Su6ftdDRx
S9+BbFtU4mSUIXWWzBdYb/rsUh5zffv5BxOiAzsF8E/EmtDBLX5/tgkyOokA3okk
oCLuJUJ8WPOjp2s4tVNZwN+Ai2WA5v6I3OBk8OCcDqfA6gNTt19GVTWijFkFpVFL
HBVl7u+gIORV0JXkPtPV7OhX/hCorOBsMmk5itl2xDIJjnyVCotBYhwiXP68n9rz
l22VUEh+u3nnomsZie17Aqa8oa2WCCAaQvUzae1trXMAlB1AFoWzPGFogLuvGlfU
hHPIifFUC9xUC+dk1VXVY9GBt6hMEL+mHok2DMV3hVdEFBmJX6HN3sqs0YPl/unC
DCk3fRJaBLvxDeIcl1zdRixBSlL+37tgdwTpuacbGYZI14GPWRJ2qUvxlOf2Orxa
C10gMAlXrp0dEc2RwHkOGyJIwOztwIapldAVpHtRp9A5CaauitFsYsRuyb2HgCCC
KN1w69N10NUMy6Yot2LcsW2Rk+zbO0RM5Bau/nNFEwPqIxB3dJYu2TG5cyITf8XR
2sU4jIGeYPK4oKtkkpK6pSZvKU3V807BOhZItbdWmwZdd1e22bZa8OxTXUXizrP2
Bn6m6QgUtfhiuWkgxLuGI9nHg7WvfepVjDr8LJV1P+R3Z9L6d1nyqojOjtsGi0w8
HmNUQWh6LmyTE8gR4JOIGRB7gbhWtZ5xyln9Ijn94gPb/4FN1boU1GfaBFzqERxg
4eGFxr7p+NmgTkmq7x7PXIWCPopCspJxZSjJudjHMLgKGiCuyZ6RLJuLtS5UIv7Q
axwdMj4IYz7sm5FAJxkpQKVUkZC5HQoD3MO6g2KQheNQic2OUk+YJYs2lCS3VvXV
JLOyhb4hjlUa0dErLHOxSu3BCG7WDM7yvZRkRsmjFRizKzi2/MEgb1fzgq7VImPJ
/u3yd6sd4nX9oq/OdVn1x1XabvfEbj5eAJCseLJL7nUHyt4DGesoltvm+Md+Kd0o
46FJwtJeyBDYK2PNfmKlZrs7A/a6GihUrDWfBBrOiE5zey9Nf33pjspOLgsUn6eD
5u6SsRUYkOQC/FRgypxw9QFQoOk+lB+6Kxidj5sE27dVpjXzFIVZ0Lm3gQrtSRcr
Ixcuo9eTC6wlVH6tWmwGY0n235PPo6OqZAYefvFZ5n+Ra2efU3dvDunymQp5A2X4
O25QKMKp5gftFNyurvu5rdhvxhuoI6tcoq10YaS5fzxfWX6pV+nNJsFGQeMxDgdb
KgiljshNKTaaPFeEdzLrvszhcgkf19tcjJepbY2jk5htj40Cu6q20PxlQyRCpv2j
wKTbN2PgUIvy30P4DiG8+W37IjJTT7wBY1G2KkEVl3mKkeLO6C1WSey0+42/ZrT5
xHzrd5m/9j4zU70REGdGA/pC3Hud6fLQ8MI7T8I3tEciyohv/DmhW0DwgI0FJreG
EitWAARhBJ6sXd7YibDeXenPc4/aJ7if35FfdxXD+fALsswKc7sd3WyO5iux4PXO
LeRZPC7jMCn3+sAuuyy6ehH7bhYgAaCy2x6PZ947eY4wJCQ7dzLWQT51UNN9B2al
k64L/HmngAw7xOh4S7nd6gufMnwzDDjtJuWBFYIS8HUOIMImtgr92NQJgPRvHuoh
QYX5O9wlLphWA2G7+5mo6aFjhcB26hGgq6TtyumK+9OPnLMWGLQixlOZHNoPg7No
HmRjLPVVyo6f4O9n/QNI+PBuYdJra3reIx4MKLduP0nzs7Cpn4syt4I/Fubt2uiS
WwqdlyzmcuTsaOlsHQooywr1WB8HZBxmUNSKUTMheyGZmBc/ho+83p3q7IQfaoSd
+XFEMopBX7O66aIciY8RPEnjp2Iw2wf6EAHKSe65auFuQ5/G7weaKw/1UNDq8NKu
eSoKzXK6JP4utA8N+Jvq85a45K408fsfRVQSMVEvlG/8Hfc3tJ0VqmeS45jGUgby
ohwmtHqO5qZSd1YQKFAIFnhB/LTuLMcaQa32oalbclyBQBn/atO1muYDGDJincNy
Wjwv1vmeqYaUPjYworgMuQ00VjfSITrQsrvxebNmZGwyj6+6qTW7qVhTYEel4/3v
2x0+VFT25XYko8vHbootLTsz/bZ4O0N3Q/le+01S9rY9g38gb+6okfE06ZoX846f
m3zYwIF8TQmWFJnEklguI/3/MIhWIflyNT5fphGs8ceHiXnr5f6kIyGdch1dpKEH
RmSlfKINuc9GhmkBkLEGfJ84byZAFO3nCnqZEPIM1911t5lNzSx7IY4Cig4dYcYa
5eTjnsUpT8M4WtKuQ8pQCcYYYfBe7dm4bODhWGLpOmGeQJtfGkpFtI4T9LWWegMC
r0aaJo7sYnJ96HMd7qaFxs4eVYPoRslHOokoPeDluH5f8ELFuR90Bg4Gzlh1GqLH
TuHG2sEV3NMmb8paXKjhbzB+bymqAQjdi3zz0onpAWvk9VmcmODzHQT/j8aLmBJx
n3GrkdXNJ8Q7eAb4PRM6xjL1LToxXcSfAZRvG0r0czgVRMH60A88ssHmaosN9v9z
fgfftq74OArlTW2SLXBiaAJzS/sHHc9dzcRD6ngEZnrQ+RYHNDnQg1MFB2bLxkLt
RO+53gO/LiPXk1lVX6vcA+Iw/q6fC/VxF3o0/3ZjFvZIvktL/4fuiiegF0VZWKoJ
VTvAvaQJ0/fmvHwapUjJQN0qX0x+XjVS6uhAxi9i8dIcR/PNSTs4oojFpsWa3u+O
izzKMppHc4jY7dROeZlzXolmsRLlWOT1HL3CT0ToXZkC62z8A7+SwQ5adg8C7YH6
dkZQgsR7klFx/l0Njlm1OrbXEjlvO4bgf9uk9w29cA+xel7MQ4xzUy/LOlAmvuAU
KsIpnY2vrk/BEMYd9r6IcYN/G6cSwP06KsF08kB+Te036+IFeoFhnwbgGtEFZQZC
bq0uXUhciocbIcfhSHebvNBlFnRZTyBOclcayPoJFv3xC40uRJSsOITsTK+lhYCI
8g/4RqnRamSAJ+x1hbCxO2Way9JdZSIYRJc3cMUCYOJeGLkWGIap82Ku9FesncLa
ucksfEAkN8KURdU+jrAk1hkAayti39yDZSrV6pFLIf2ZUFg7Hm/Tvd/M4iHG4dmH
EiJpYbfi9V+wWJ/wIllOPnzzKi6ba/x//dN3y16iNu4qWeUVLAIR8HnL2uCnF9jr
WWsPUBC8Dief45L8HkMjCtt7W0SicRl1o+FKPm/5Wfyr7ajqD8D2Kl6wS8BQ1ehy
03BdLY4SBX4H6JnWlZ9sqZC2dGp0QmsQz1mEMBSKzKhJ0R0nfCcgn7krxroWjs1N
qpYVAB1h8s24JEwgcF40Gfj1R+1OztDAe0OocIsayOl3sC4YDvCClTm9negFu7eE
BVLLlj0btWkgdbx/JqfAkS8oD6oKJVW5nCSTqkuqT/rhwdYfzH09aRZ27cn3gXmt
684tEHUrrVwxKgcKrLjwnV1IYiLD44uf22T5wkpeg2wnQynWSbcQEZFk82zARpAu
8eY66tZcSga6DjXb4RjKXAtJmQS5feqrPzhhLGE4LpLetPVoM6S1en3Uc7GPrX/G
yIO4pEOXBEdvNv3WsmOE9zKClVGlamC4Li1IINMpD8k2oWx1c/S95NP2G6bNqYeM
MsyzCwyl08KWgYMjF82acvelazTXBGkAZjx06aklDWNWLFxbQqFqNrWAiD/Rqh5E
PDPjSLPKSOFpJhQkGlj9uodWhseYDwfO4TXR4botrx8XMCt/QlLvXDClhNWl6cw3
aojQgeQfCFm05geK+hxvRGCbWDjS0QpEmWlDnUUITU6RSyopFKvAeXpf0lDJSfkM
7gSaMBpi0wdlLaMVTMwAK1f+uj8r49tgPj3OUfY9YpAqrpjGPa7bb4MMp5e4rX5e
FS0BrqM2pw6Jwu/+c18BgkoAgsfqU/EKwHYJ662RsLRFdLTZXaR0obLMY3CwLFkE
PRw9YggRcswqg4EyRRDY0SgM+w6CpIF5xgEZNcnVM8+HgDnie4Lyzi4ZMelt651d
aJI5QfO4crt5Z510KT++98VSHC/U2g+MViESCoXNs8/C6SLIv6HnttY3RCOXrbh+
Utv04TnhVf/VDqpqgGlTRj/R3dDXbtP8Qdj6YovOSqk3RRHDMJ/uONualmQ39CAP
4qW+TIy3ciPOothJRHhie5dGopzlpDVCcWQTXUhY7bs77MsBT86LCkbnBy40y5zN
GdRbUbUcQR8VDrNNTuQJCGYq/8iR8GuxJwFdj3EivXGup0yg54qSP3lyxKpxLxbq
RbfjxaIyUn875Qx2c4cm87xsHuUeRZVPI27S0s3CCZPCa2l5WyY79kI54G62JlmL
sKbud0gm0EyB0q4F6eoUHWmN3TSMlZ1UYjj0ntBRIL1mwhAzBg7lHKL2WxHDdLVm
RNz49UYmFiA84uyvPBdIMZUCgh7NNdq0d5CK3vdVFwq+dqSPZ2NaUcfsvZ+L8izD
cl3+0hFlfZ+c7Z0eFiJ2Jx8H1FqueFoX49WfgHWe3YXcyV0O/g7hnwu1YCriyho/
kjJ5nMS1NPKuRFulyPKC3LyJj19vPsvZzpBsVHe5E80UDyJdLNtIYLeaik5Ut81+
/LwtHLLO2GegiVI3ndml91Gh4u2uDs5nWU+iHtbYQu//1M4VhbS4FPccYrM8xccx
P7yTUjedp8yVPNAdj3tceeXjlIGVG3G9iYobZOCtw+SCgBQY+WWz0Sr6kLvucLKG
aoEegrrMIp6UR6bbwag2Jadf/nGBGpatoGpkAoT5p4BB2S0IBeNpZAVVEvMfEzqv
DpbDIQLnAq2skS7ZrqQ7CUSqveTSuDwu7MUvun2aOR/CE6yQ/PAp/XkmwwmbHtH6
Zty8rF/1wFvNiXI9H8Lus5kKgDf1dnOXVtxQqIsDWdavpQn/uCtuePnSfXKxHy+L
yyNh8QeHlyqynDGHOXklN0AX4M6rkJ7X6UQpJy0yb0yUzkMgNt7/vfroxBzh2vG9
UZIUCYmf1gip0Wprt2+7BGE8fFrYFHX/5rKSZyn6ZFY9tOgVMjYTq9wCZ5N2BBcr
mX0oj1YwrD+I9JGq62lllOfJajJifC03Q0zTzHWnlAUGTmJkZNajh5VpNzKIJ++T
SG9USBmENS+lsAsuLEAJz4YxK4wdg1Zt2ibuSKE8+EiCxERVMPz1tdtMQUrQp88X
l46BPSR7UJ7TesJrrDg14tTUByEjsFPfiCRmtbaDcFSvpl3d2YKSCl3dJoq9K8Hg
V4KLnIex/iV5uY1yqyqvBsqF3TmYDYugKaaFuvGjHNd14oIqv9H659Rph2ttBObs
NKCuUfLy3HTDRrIgYigcibpJHO1O3l+IXa4PKNL/hu1CEb99DNvK8xRfEnGK2Sl/
9mPF5T6MhwK9hJgX6aeOyOjYXg2hygpAWr3alTQv6vYpApo66EX0KzY0d/cxiXTx
OeggbHWZU3Mv93mZeH+fPSV0yOgBo9huR5rWvV5Kw3uEQ2XPRn3jHPJptmf/+244
ZRQHHbUczjWCU29qennlkFI4PKcJqdQ9AfJsB0iWOnPGkNs7NvPrmWGCrwASQygP
mq4JviPtqLHZQC5EJR3T+yisvhzJJpTzXz+HaYWFBudHqQey4cgUkWgfxcmOT3s/
WYH7kcFw/hxs4fAW3ES3BiTFLbSI2hE2I2sY9hAjGAOazH0+RRk4b/HYfl7wN8Y4
6Zd7N7vkpkk7khaSbBt43FJMrwDlaqlvFUjXspA+jYzkDkatlCUQL9DWZ87/rgyF
ZGHwBYg97R6Us5L9BHEJ+26zF0LVEN+f/Jzyt1O9wFKVDWiYBIeJZYEwKnx4r7DB
Rwvn/1IV5L0DN7A75lQfsKyObg6dwslviWOIK8fisJHsDqSmZPozbFYcK7hmiQPR
OGvNjicv398jic2qoWlP6MS6jE3e3d7AWff0W+58JhcL3SRUCSSpmH3exYUpYxFX
KI1pYbkU6oh3a53SA2qph5P8G8qoCn55jo41uc9XRX6u+mMFfwXwWBjQwuWGpZov
zikx8Bk9oINEBAgrnnqsHFWd2+xxJSgBe6CupuynLUWD4zYYV8ZQwwRmB8q8qXpr
MQglPR9u3F8Plnq4zg6CjUBV153AQT/Cqj5Bel634MTOlCMpJJiU8KY0z8Sg8w9v
jNk/Vzv9F8NfristukXedtksEGrofiCK5Vsbpe2S+g3ALxMxcRnfkM9akC+wvXaS
LBIGRXKLRIa3piNIA5Usegd+kUxMvS9zQG9Ib90/6v9TRJvrkvbYEGK5ejCtc9DN
P4rMyEkz1TLphKcN8/D0GhBgUIy8GsQF/Y41VA3xZbiK92o3gUNJNQr/aGUO6ALp
1TC9AQOYsOGgLXVUFzNGyeySkeYKd7N7QA/IRTR3EHf9EZIXV119WbYec68UGMfr
c83pvXFcx8Mh2873aD4gS8H6e1pcwek12hK3Xe+dfVX8JNHI8PjFxHfuUu2ExEl/
r1rJXgOJEBvncKdmFT+oQLvWGfKinfOJ7RGzxo3IKgYw4gZAs/c0q2WpVd7GEg1M
4yCnGjU6PMpQ72ld+A36aJgCfCyTu9OSGnwmRFR7NsFf6qeg3psPvTAZzOKrctIe
ReAuYErbmeA9EvOZKevNfCpd94qRmauSEHjT+6Xk65R1Zlo5ch1NmVoh/BqVtxgi
3+l5S9pgza/UprwHilY7tzS6x24Gbk59K9/nCbeJXZl2PNGLkVCcgQ4iD53yMsij
myyWSmxy2CzSBghGFkSDtqPwHAQmjJQ3f4M0NTuBPckeAYko4pTw/8y6Gno3jn+B
gRC2AhCTgGgGzEmlim0R1IZn1do5VHjHF0cK017/WoPt+7Sy5XoJyQ7r4N3Jh+Yi
3WoXtkmS5QZ+us33vDWDb+f+LYHH24rSZYTrXu3cwYalKzVOhNdeANJ9l28XJBuX
l1XENzx5pQtkMxZY67hPYMgYus1wR9HxX4URjGv31Iit6tR2Cozn4Ec/S+ds0WSZ
7KtwyZufaIoOawHdi4rnvCJ0MA7GuoDaRfX2tpALO+MNWf2lJx6X8C+f+xkqa60h
s2aAHRAniKgkFfFYe/PfoNPzd7eVcBcn38dcTEXO3/O5h2eFDc12QbXJjUSd6qmW
YXZoParE1g+kAbvr3FcCAElRl2ed0KiSz3W7fV/J6NWWmMiOtAmESjCYY3Wy8Seh
l3NKOtfglRfDiRV0wU1DeoTvJqpxUG7VXigEi+eIayNoaNoIYl30EMfviLQP2TVM
YEqk4tDyeqJYsOtpooud0hFFWURLUyMCpBnpQ9cCj3zv1Irfr5oSz80VqjPvF4hg
guHFInlwJE/rpI78ZqmmoK9ePULYBJMkIlak/rnXU80JL2ogo0ex6+LX1gDMstcq
gcCNu7D40GZtuyQwWTq9s2zmMyb0R+7diMgrKkkPjpVe07btPQ8OgC25zfzdzIMC
jeoaijCcBwWUbNZkkGyZElT/RjrPWexLVfGuhjv9GEd2yhDQMxUth+g1vXuc7GNk
6wy7Tniba461Vk49LhlTZkBov5KTcLIosty/okS48DiedzP+aJCjAkcEqiB/3Yym
MD3VNKvJcErzLR/6ex9Rlcwd12CGebWRZMMhtJfxKp1UYuB08UC3fdBdkImczq6R
R2mFVT8O2lLTwRXeFvwcveiBi23rRDNOOMnFXjThEdeQchuhnK2vVTEyKiHCBNdN
PWOmwf+kG6Sb+NGf+RINWPK6xKmsMl7+hYZ0L2QRh8SQt7uZwkVRj8VDVUbL3gk+
v6Z7ngRtjpMPOiv5bB+LPtJ2wZ9IHw0M/YoskU3gnO3LPctlcilLrQxIrqfZh4mA
8fFy2n0ka2dYCC+mZY4yi8YjwRhXE51OxZ78h+Vee/4duRlrWZq0+5BQvKmYUSyc
CYtCwAl2een5dcL1wjEm6Lq8C+jX2aW6N3OzkU2dBWbJcPCRY5w+Ze1SgfL1j41X
bKnAJK7heuNul/SRC4fqFr0ZTbApqwVbysgaOXmhYTjFu+qpATyKKJnrGxLBViZr
BQKTYem/z4tUPqhV9vQyMbvmQL6l8VdpOzqwIyl6OR4QO3pXyPOgDLJlNRncdNK6
vv0kwkgakZyS0HVlGbXwPttdokRnJyQ4i8vMF/KxvggtPjWTsHt0TjmmVXP880KR
o5Gt5tpIEFRuOfFb4GyxZfGGrfQl0zXKwIi/suMGabFmQw28ABMnbSgCLKyfQT3j
rsu+FLv69Awahuj5HvpZEgkaE/owryyuVDDOMGdKFqKYeu47VA3qNb/1nzEhM5+U
fRrhGtVM4K/ei+C8XD4Z3K07jRtMjx7+ESmtFDV5Pd0f7eXGsSWA03xG59RJs5Sa
JVZmqyhOboBB2ccdp+SPKL4T4HjzdiRp8gxAf88KWFy/tDRFHa4IXIUwloB7lv6V
1Hv/SuJqnehxgZHmuSYyG4DN8HelXMz6fL6ByO1k0Rot5Ijbx0hP3+Wi5Q/1ddO6
3M99ufKRHyGSKeb6KF/wUkMNPWPRS5moo3u0Lkl2OJdGrzV/UhJesa59roMs3GMR
7H6pyOlm7DW1fwvcGF/gyRPwhfShIirw8802zIdtg/HH6gTSz26fpwlV6qEPcEsp
TdhEZ8M+7nNi4maQOVC6wHMJcXHJGua2497Xl986UX6xeOCuNXQUIEQFa8fs88Zf
EKsHMg5/PKJHVMJP9zBla1eTKY4wIziAfaM1NcxDjTlq8lWWPet2MGsp3D5JpBJM
DyJ2yaL9L38a/YXALhbWgC08M55aGcJ1Ou+ZBrfrX/i+ZSCsYsVQME3X7D8aDCbB
EiKbFdru8A3HRDbxxxUo7MGFEvenvQjwpS1WP8pfc1WDEEbcwbONqgyne1HC0yW4
DkuIJkcXAqrR5VlqclAM9P9Jo0uRmOpNrNwk/LO3X5u6GRr7O63KqxMkZ2FC1On5
RanKwSrFAAzQQrEkXItDNO//q7nMyjrrEqn3WMjkYCjjpHw4sWm+xEwb1dd3S4E+
G465C86YKooFa+gezfNNSwyzwA7xz1ytzFeRd+jYbRTVBnCwS7Fe1gXdpF/zEsFk
iYfVS6vRfgFYruCwzxX+IZxVYYbvHkLldWq4gAwtIciadaJZBZIPMpVc2OkZevbu
KntJzvQoC+AuOtm6sCfu4R32mwZg/r1N+vUwSXmNImuQl2HgR+BHAgzx47U/yvXX
cELQ68dHnH4X/jf96q0Qz7tqJUeYGzH23IkAYgmiHAU9rCUDd/fcvd2kPuk+F/nl
g7dmoQ3q1yQ/w9cFHTi1CHLV7vg7b4XVEOuDPRQh8zy+bR57r6h87AKmDcvp6p78
jUUzbvzr3878eP0iNDnBkC289/6dD3FbnmMlwynpxSDJ9AoyLZsJqKIF7mcMggNK
untuQWFendTYXh9wRFdp1Hl5Tx7VtDng2/AyzB9dV3TxdbLws3TKuSAdYk0rtRO3
AXxo+JI405IpG9ly6ReuWq4KFOPI2nLYEJIwjnFnds/qt+jD66ZbQ32h/lOwx4Xh
TZZotHybYaQeLIfc38CYOJiiAyAjx/HTx3Myy2bld35XFZ8ryYkJ2pr8H8PjsIvi
Y8KIbtVWrFyPMDu19GRp7e8IFDhyiaViNiaOPKXGoPX4+Xh5yk7vv1UfqfxTWio6
ctYWrtkiZWP68We6Z1j3jJ5dCQ0cIc7QdLKhvGQYk3xpeaDulO0NkKILm8Bwp2nR
qswFVDi7idvZWqhAsaVY+UB7460e3IYYeXPrTHikPTI6/FDJuTyrlk6TeH+nL7/C
OqX2dx0z0yQC9Qo6y8jLVT7L1hzDEg3mOv4s7tpMqm+aDQZXihAzkTnzf3UnLM63
ymfrkMwWKQ+JuCwCp1TTrICU6EaK7UtO9DQCVJrX1/XUsKpFQZysL6/YcPuFKJ1Q
Z48IhbuiavnZEFnP7QzXSrNpL8Nu3tpokcpTYuTYS1gN37MbnxQFL1J27Lx8vUpv
iKtokq6Pk7qyGGA1MIfgVVlfSlKa9upu+pFvlaVzrKjCHDEAzn+Fo9Ku7bPLu1RD
5Avv9KRihSXAYMlMUdUJe3VhIRZ6hzvWMtk3l0tHSzpLcdL/HieGpfFfsXTkuRLU
KWJBO2/P0+KibLyvjwU9GYA824zFZs/eQNQ6MX+k4l+Tr5lCRobo6CXfNu2DzFJy
dlv4sYkpoVf++6iaLGQ81NasjiM07USgXVHDnidy7CCDBzBXm6Oqlw+UKJJ+onu5
O4wIh/sDzexVP0eA6QzeY1HZBUDjFUjGTdrcF0XqOjbgf0bm8PqFj6e8PwkSR+lc
OMdTu/pj5e6V/mnvx0EIgCnZTkl1wOeUhpZicqyNoWyRXHqPo3gsWlicMau7xgSk
8n0zJ6gLCkDrCb2wQGTY82I0pkGvFU8w80xY6EzErkNysDzBAaD3fkuoY1n8rFaH
fsTQ4jKO2lAKI+OVAqFWDUGWef7Z6BpMukC/zHDdjzCXGxxtPLq+RrVXKCj5e/hq
Wt2mvjUwnjYLTahI1SQ57+whv00Epd1ja4gxFPhkmaE2ogFgV5qEH1Vmyz0eR8MQ
xdbIYFRMBOjZYOrGqm8cdmppzi5O0y6MLlyNZg8IMyab9jBm2pn7V+N8Yu2MztO2
kcbuX7j4mtMAxMlPEGXbo5PC3D1XSLOnnMzmT40VsBFECgVKQ53lt7YXwFwFsAZl
j6bSbUCJJWU+MDdcVqD6U45CwR+r6D5e3cafi7GTB7OGBxPWG7I/yh+Dc9whN78r
xMEFGfAt4kTEDSqGFk8yM5kY3fBqaWxMgVPajtL0wslUK4hYMiwgg61NVCxdLnGd
2UTPRdY4yips3ZSX8sq6dvpKO3KAVmzTMR8tEAwNUZcjTNE0w95wmEoiCKhd2+C4
+wFo8bwsCL96Jo/vExi8lHZhFw1iiDOtr7jioG3y46lgvmT6bSnCy4xuXWmBJm1h
JRoSk1lBZ2lukUiFLyGguRnIaYpsC+9iARSDhd2j4huNgnwdY8BsXA3JMayde2B/
RejjoeibZkq6rHJWDWmhoSX0eroBgOxtyVD4KVslujhOPp9hINNGCF2bqUN2RJxJ
yLxR6OeITqTZcuPJPuCT1l7MOI2sca67TabZj1jqdQEPoQkcyLLRXEs1AJ1rlUml
aPG2q4Aqo4SZFa8rUZBB08KmqrkRXbQ0bpnsBG9PzItv07q8AQKxDimU6Qo9hQBR
SKDbrdk7Y8Zu6qfON68Yfsnujqd28SKEAfoumnPHCiopmPPfFdo7i3YzIPmaqSAq
pUIAucf9fcG4eIOzFK8GFlUUziq71V+2ywCLyOcfyR2XF2IdHSg/x9SU3tPCt3Hd
Ji7okvFlgzSGC8Vxg8zLsueMncOT1KDVaWGAUDAkaViYLZx5jXQfatbkfK/HhA4b
ALuA4JHWJRg9N7LPyKRFw8ayFN6QVNHSIjNhjly4L4deoyRgHZ72l9KoxzBXwYGq
9tC96kxc/jvn8LxgV8yT085qJ6WS/5Fm6Pdow7qtWnll1yij27xiFkEpAPf5SNU8
oWZdCTIiueunWLoa7P6HP8/vVZHHQGAcwv3GT4lOyhe/ZQGixWKXOtTQTs9lKRvf
fc67AoNY/N+kS5167iqw0FLyucdXwfhulHWQXTW6C7oW673s8cmJlkrculPQDp58
N/PJKw5UM0NDByu+daSFFcVkuup1l6kws/GsweZQndPAAn7cHWU3yxnpCGoPZLD+
+zkDtcXOY0E/64rqkaCKuaKE/0oWacf7rwE72JKtY7F07bKG+EQ2JIiBEKvyH3Id
Lo26pnoQo4rQ76k14FzgRp0euis8YfeWM8SHl5TwsUgR0VyyKH5mNx2O8EMVXTa8
JNme/cMnhc/Sf6IVh1hXND2JxUNtQ10lZFM8xCksYWnvwQssY6+f5VIivBtVUsIf
pddsugkiucf500YqK5oY8dopKjVEFZP2BHRfowAhzphMdZmDHHdD01towVmVPWqv
6PkoIm1vYbVKu+N7tUygS1xxnD3huI7V2pTMjRgmsmy5VIoggiwBbk4tdv748Nqw
HXBsYeZbWFpqo9Uj+esCThMpW24xidJqu12lyxDhMsm2h0GQh9j8RoYHI0O2Fyer
THwMDjRE6s5e88Zk4MTDx9FUztDEhjR2K5U7OAyeHzAdc+VVTHQcoKisrBV0R/0N
gmyxV00V0f4+yGMi/zlUGUxfls8wVL+TnTtsRHr71VtOVopfpJ5a4xPGxhQbGnGh
uAJwVbJNWp52GvkFKy85by+TdYvDXtX6OV0foyLstLG7irSM9wOsobxxwlioXnq5
eDTyJc7Goq0KEohg5cz3DTTQ3edPec5hb74IW2gJXATqn/lcZHyWorpdmwZMiC/i
1Egd0YEfo+OVMWFn+0ncWOZ6U/axYzS6f8Syme/YORYXgrBII+cku7DuL/UrDoiE
A9/b4ULWsbZspqc7x9uCncqneGWnR36edzQn0mMikFXDAMGY2Gks0T7YD2VBM2a0
d3dTBXzXNePQbw1SnwOF2NQIZLPRMUstk2QeLCZAsWMUBwtSEu6WEHMvjzhCP6aa
kWVIPVP/IuNHEWGusmDwGUnGaTV/CmgOHQShEsxWRWmFZVIeHnpHRgxd4eAojmB1
JA7KnwCfJbDq6VLpz8jtF5wEvyaWD1dlhrYn8b/7WDZCPqOA4VROngZCRFnkrmnq
DUFo5RDmZjt70rlsZ5v3OHWRT0LCzjBK3MxV9hCFqRgWWJeY/dvqhubE1sxr+Jii
RUcqAQrSC4J914OEJqDHmQfvLMgXJ2UJQd2kTlSK1yaJec2J9WVasBhJdv4TcDat
k2wYFSZDPiUIerTAzxrWRk0ThFzfFV2p6LLnxh/tP2ZMulBh1v2gT34xI0vvOtAT
83AtiTYxOzVzo1WypnI0MINEOx25nDCpNxuGVClURBwi3EAqj5zRgn3wg/Z8WmYt
Jo2gLzFBx25EgZRM9THzkBu39dMn9FUZSRcvlt2eKppWciW0ivQp2voi117M9bhF
RYaupD61Y3bxINMc2GNR8qT5NMaf05IZNvZxhcBZx8TxeVEvFZSS1rv7q9xSnHzy
4uC2uwDB310YQeR5P1YEnPKR9tMVKib2g5Yxnu3VLtiVNR6swkeX9O7H14Ltb0Qk
B1wMQJy0XDI9mlTwQplgjfQ6/sD6clikUDgoJM0oqhdCjYj2eeX7ohc2j/2sI5bH
rd5UciPolfDJ1I4ir0DNG2CbuRoGqdBanQf+rJSOY6FlZOnT/2q+sIRzFsyfHIwn
yPVr1WOyN7XDf275L/MCU1oVNMi9dB8BSvcbdou8ROZfvcTliqIu7UhcBMs+Xhcj
4iPthuMDefxj9vNb0JxVahx/2pYpbWcQpMzsQlC8kC23NZnNEy0Bcsj0PFcBZhtC
WCkeVsFRIydNeXBti/qxXbgtYrA51j0hEUydeA43uyYAcqLD/T6UncewGFonTPEb
mSX6MjR85GI0ZsJBYIidv1GzrXuMI1wxyE/NUyMtYstr1Y5UMVim1pbXLoNtiLVS
UwaP7ZEzNz1xiycPzyD7CPHhg46WL3x6fEHvDBWmQ3HW2XUriUBjZpmm1xnaQAp1
dhNWBecyUBd1zc4Y+DEaxkMk8pQxVpCqUOY5lL0sip9AwDL9bBK6j+UaG6oY66L7
zLQy5rf5Kn1YRlu9c4I4+uLlfWBztS7lsTcgnTcyt59QE2hJNTQiVeJSha70OXf+
P8oeWnyaR00n4EOad8yzWlZBCypqG6Rki/Nz2ZBank3Hr8xTtKDQ0RTeB/LvOug1
ra5l8lQ2/JD/HsbXvsFGgYJ9PkTRMtzEKjhaDsrXQRhWYCSkAOK3LZyHmsSLJ1/t
e3ZDWzdjD7ZcyPi/yDFCoygmbP7Wzvbg1Gf6zxLmVsQZ7V4rejk0qh0ljOAROSyA
AtBplS/mz+FueqSVxKxfk8/JnBOzV0iMDyyKhQ78HEts94A6hFqBwlCdevd5eQrZ
WUJbtXlSKX3bYL8RnQtbQ6LSsMb8BUhbAmmpm5Z3hBQmpxsMPkOuiDxhMK2ocWia
0+d/Atn/OMNc8QM4qWkP1M1iwEFOO5+5Kp3a1F7nOIXeq4YqKnIegqMqkmLE3jkY
iSCkJIaNIJVHdU3Z5h0GNDzNyE7+QFu4UDWSYChgngGSajlk6t/I28P8Yt1XxbeL
BND3hJW0HrLdwC7xRh2pva3kN//jOJG/DGhG7o5vV7A3ebt7JhsepgZ9NCfaRFYR
h1E2letL371Tbthig642Y7EAzStU00O4Hx2ta1jD8if8pa1/W4HUOye+Rx0MaBVW
HLYXlN88yI4rAPGjr+L/cJrLbdjM4sBRNIexvQ0DB1sany4KmQWdQoMlIQT2ClKD
CSv9Cw++FyP6ZIvGokZtl+g/a8pveD0mcjoRjOvcpI1hsnkh1WHKJKbdRCIV+2nf
01Ff16Z/EcjdJF12pdbqbOVIwxHjYVlYc0iF58TDxGxgiPD1PlVApkwPlhuIMDjV
Vb+UWxNBII9clGZUaWjAsv9nD9ErPiMYUpHfSYPlRWTliTRTzO+Ecp2G0K1AYSE6
m0ZTbvz5r+eTvYqenVsc4zNAiSZejjEDKy5lMaaNgubHncCASlVrGyHtsqPRvo3u
2mXbke8KykXHvnoWheaZJ3MLfd6JyjWdgtnvRKfLli9BNYJAYz9MNBhgAfaRQFlg
ilk5aKoHolQ/Ety2BnAYy+sp3Xlm5IgUXbEzJgNW1LrO9CqcOwTI6A1MBi2YVU34
w9Y7J/mU6QQueytcW9wlG4Xu6RVtgR60p5VoJPwe1qS7Jn1yWtBT9G/SRE40vHsd
jQyD4VT7mgCcGmsJif14VIimIfrX4myJD6GHy4gHeUzxmhcnl/Po9pBRscNQ614H
2icE02wsvkNYPTCSZF2x1Z3ZnGzBEfRxloLOFHwL7ynnmmEEdx8h756K4rWXBsAy
J4IxlX4hRVTkXc4XdLhSXr4hG1+DxPqYKfl9/ylB48cxW1eMVJoCkpdIRPFpEILB
RUE+qlny1AoY2G7F66TBbO/vb2nBecvgHMdXkf9zlqst3/jT0Hwi12z22ZXKogSW
HgCkTS3T82QgVMa43FM447LXU1NCt3o8VTy96guqrZdzOi/OfGV45yQgxLbPTLdM
gzIReZwi8ERWdfWGwDNs8RgusPaX0ZAp83KFT1g6UUJmiyfwuT3ObACTKm4+DukP
lZownNqyDYSvmUz/jL8utxkCgasXm77fqdsWMyIitBVg4x0dIYlkfY1/y7bmvWKt
fRUzKjEUu8VaDFcR4NDh3LXh6PdLRLxf6+1HbuZgpL6ddAqnU/V0IRn1Bx3g7yoE
twS8yYJe7ONfQskV+hNTVXVhkBcy8CL+9IarO4g6N1KGlD4yZE6F04DPKP1P9pH4
1yd623uX7e69Ryz4eCH1A0vCC55CCdlF8XR3EZtV4XwWORVmodCi/RK8wgYolSYO
ME6gAWOTjUCGPf2BnKoa4uDxn32E6glqob7n5GgEKsxytzrXerVSg1AtxrNoKuWO
zSkMhZJ0eH5XFvYWJXqsFF4X8432ymymVV/vt+lIob6Wz36FxPmMooXGMt3mFgt7
16y9WcEINnFByrFZMBzWFeR1W6Dm9QiDwwXNLiyhDXRTZydB2PiHbY1fwaWftdKF
kIxJH3ir9UO/MHiw9U7nqhVPw57bY4QTtwju5Epcj9MNy2C/TiabatMFyiQbddjs
zI94eS8a0xwxvr036HdhWr1k5HTikzjgnNkK4vwpvTcCgAzeNz8WEO8pvk2EAola
1GDlOFMPNZR2VXCpBn/QhjV0g4ehBG02gGUUIPuimWADNn3IUAkkJLmTPKt+9oAf
z5T7Rtpso0YwcHnqBQGTMcQDY1Ona/Nou6DXIsduvM2D2eJ4rksMWRgM4bq3M6Od
9zxWe94WRECAlQEDAQE9kUWAo50wbFM2Olt6fN/V/IqQ2hW2XxBOPH4K8UfkPqfB
MPRQXQycrMKGCI+ouGJQWyx6+qZQHzuCdD/9vHsLhOmGVBBuY6jknU69qgiGn5Wf
QOWonC2SQs/qiPKVqV08cVcLlloed+pfIpLZIg+80yCxzwS9Tws9pSp/ruIrD+cA
IK3r+YF3oizmrRs4TiqvOzwztMSAhTS1a0ExNQzdnBVEWP0bjSlcV46tPGz5FQvX
3KSvE0ID0LO8/EaCMcJZLXkszaCfyU+sWtcjoU6zZsrDT3SUfWvhmrDO2gLJaFje
cggO9NP6XI+7F05C7vi+GH+SRpDnH9pCNSTO31cALnejm0+jX4XAUWtE7HyXVOSb
v1czclMWzLomV4U9pDwDBHoUmTscoK0TyD50DQoyqCjWgRPBAvY8jaW3mdddiQmj
aBqKF6M9NtFraodLAlN8F8P6nHbj+7kWDnxFd2kMTBIaLOujowZ8x7pQT4Bv/ZgO
/Urm8jIby/NnwEyDVKl1rX6iUGVL67dqnRyuslVCQMHCQ7chH1aadHqIvEkNPYcT
fm8Ld7IgquoOGsMHJkZB71gZ+OXtr/Il5UTvKD16I+QE5gDw/x/xj1w1i4m2mc1F
ZnhXOSzJfh1GatgPSHOJL0eFpyUzDDIae7PmareqMTVesfvmFh8h1SBHrQLjvdsn
8zV+RQCcdDp+bZZ8LzJ/n6yb1lNXd7nFGt/iH/AAreO4vmGCpx3cO5AXoU1iOrdB
jq8zjglyHwKmdZ5SZsBZphssFuyGfpWMjSYDc28NVr5HoXppJs3h/C8DWiXLC/eA
hAf1lVPGMrz/Miz+zbyp7qvZSUATxyvbkPvTMFyWPZfRkvfKvwn006GeFxUrzdF6
lpShL/HfU7lIHtjvaF16ggf7IXF+eeU01+ooZpJZ1CXuoAvOcSmVXpvmKPwZ9LqH
yaIu2fSjunH2ggwctVXRInOjyCa3xdMFW3vQn7gxbaxHMuDKOmQ+n4IOEbfkyxO9
aY6DLCydV41NZ2EmOer1Dw6ldResPvAcKSShVP32mtxRQtv5CZ2a1NOZ+0Hq1JrJ
NCk1Y1GRybH2y6IFXpcPUUsPX//s1s6CSct8CjNHs4HCB22whDsPXm4K9D1tQHNp
eUDdCfKda0+aXqtAfH8IEsvnlTSN+rQtW0YOQWz/jEBWfLczcvxKWyNpajZbWy3Q
eMYAy3q7dcr5+AT75cQZoWdbaCy05o1ailPazTRFKbaI3/0DAyeHInXMFdNdkOQ5
xGgCCFtqNDXl8+DLSXt9Wcz7FeF5g8yaTXi2Hg47kfiTOms27MyGq3nNFkNfe9BF
ROGDwcyTaSCmNmRr+/8CZ6pO/qvpjlEcXtP3ulnKOI/BbDL+8v7KNw3KkdFb52ep
fKVgcbOxKFbupxuXNGjR+81cwU4ZouRCVoQ6N3i4UPbpZO4NwC5fb2mPcQYFOhxu
ZjsSfx43y8lWGtZAJxIMOgkcN++1kjmuZruOF5843syk1wJkNYI9TPqsG55Q7u2k
SbSwhZcv5eKvqUsdzrczRV20d/lfp0qmEm7K0u6PZJWdSf6HkdV7V65S3xh442lh
epRks3lrCdhabMl76GKYfyJiqR3/kKpE84XYW2g5y5NvLdpz45e+BaRI17hHJRwI
W1nnkvtR2su3Ny6mUP3VIQQJkeQea0t73vwhDwMB3E8Sbi/+6O2WF7LCEAq7z0rS
jLg5gqZla6HaEvNaVykmNBXwFhXXZaCs+De8p3pnIEAuBWp8a8sOZQgSnc4zCEbV
IWLyLFG/hjFCjwIqNRfTaaBcaN6Evg3Uv9Gfiyegoja/a/raswqXufTx21HBWuSd
PXx4zAzgkISwM7u/ZadStdnEQOd8sJ2DFW7CXZtbZyXLvknuGwto+1/TJMyNfe+h
qv+FAHC/Dt7rOf9Mo4YlXl+zZ5B+OuaMysKy1ZpQeih+uSfBwvo/E3gAtrvSh07Y
mQtEBM6NWZh9SUXAMQ1zUMxO6eQb4+Qp+5dFmZISm7+Bp0gTf8Kzw2X7bwffIdL4
jSZg3Qxekrft+x7HGzgKtyWd+WWooJsX3/H8oPRw7zw3G3gdBxLemLppae3V8ldD
yVcl/qKdmB689VPvBGUOQ1cMUyyLEPcGiRoRlJX3nam3EtWNg8YslpqNugFcYDwE
54ic1fiTWmDHpGIjcJyF6/PzVSFU4bFO+UUlex1WWUps0lKg+xpHzNjbYCTljjRT
0fIzmj1Fa50MkcC0P9DcOBcEzxLiHiLCJxB7FdrTp8+4U1bP53P/R7twypS36B5q
E0w1ACjIOH+E3DGhSdOTjqIaEXHu367llxLmJ5C84Q6DSMWpgDnxikQn9KdNtN4E
g26JZW1I5tSotqidwJaAmSnKf+cSdjOiSrEXSotiP4Q3evb3avNRnk2vmRTFhGfz
mtFWKdNRLd/4727lZFQFIB8WEfzxFgU3j1TrmPP3H4pAeMwUO9U+0tvHN6ccrvfA
iv76/cp79iBSfnzSbvPr5p3LRFCnfwfUoQXLwPLuWiRQoTjh2sCoVe0rUNfwMY1F
MFP756oh8dCr0s2Y2qVS3LYz0SKEo5n4K85N1HKTgPyLqFpPtunlANSAMRaQ84N8
LoXKyPd40w6cRLB9HFliEZG3WEkKTO3kDepVTgNwszsrayWyvlTOoRHUIyRjCsFi
0+IInvjN028uy5rAeSvTMcveMlRBHq7HzXyL0APElbg4RuX2MU+OMi1htYiZDB3b
Qq33mJPENJRJIYhoa5W7xyWWTygjxgVocgu8h0kgXvbNvmA/B+Wu9OI9EAvY+pJ0
U9IE/NkzJPnXCUj48IpZ4Coi2XevIrFW8cY+tzUx385QI7U4QxeU56A2d0i0NqDS
dJ5B5e6X+x42ao/lsmFjd2kbk+wYRcWpgBuZ4oC4B2U3U904Y9g2gQv0I4KGVwye
Ob2j7RDshZ3sgd1cCbjs5P8VknZlO8ei6fVbTRQDe7xcBuIgFAUv41zXeVyKLy1c
CAg/99P4gsPSD+Dj4DMc5PjXQAezzNGfSGGkLYqIkZwx5I7ZN4aYEjxVFAQXGinP
5Nwq9RgdH9PEP7XWnTJWuCTB6SfM3haCZiDbLHlqIfy5H97zr/ZL78ERVuQTCD+A
Q1bmnkls5yxzlDsV+1OgiA+CfhsYweN8THd87vVcla5bGnjnbWIfrQYQWjYUwofj
sxfRN9TTzFTrBORStysTwof1Tvjn7MNlN1wF7gbwDBzSL3S+pswltRJlRBPPJo3F
lLQUOmMgliNX8BmCPszATYIGpd5O2B/qIfdo+IszY2SnZR4sBXu4aIl3z0WwjH7f
obR+twWMFLE00KbqXhMN9ujMXzIuof6ReWcJx4FN2fxx+o47QhjFAvN8+6jcz9Tg
1b340ljOPLOzM9HiNo2d/2gMKrvnbAPEyBiwRfGP+j8pOpk1blGv7qJ46pdlmlfa
OWI76EKh40qKIw8I8ynnDkegDkdNAC6W8lUAQNSVVga7QBVDL9V5gq4X1beJ4Gc7
YyJnoRVlhH/RaZthg7s7GMowsRGwWWmgEj3O8BZk1+MsG469SsPc4bv/hmVTe+DJ
AQL1BYuFrD7m8R3eodiAuMzFx2aFaKaI38fzb8WeQKA3MoDADqkJflqh5e5w87h3
ZvVzUY9KbjRKelfxnOV4pDex0hLHfqi7mO1Vp+Ho1eNrs3nK7NTRroDFNrH/SiFn
dLSfCJ4MRZIGWHDgxT75DO4IScBza3oVtihvQzaNmSCD+fk2B78w9PKtuBc6Ahkw
L9muG9b0TCHFkqj/o+Y1D9u+RM7MjxYKMCC/2RSfmRaqiziOT+lMa4xRDi0ZnyXp
9pEI2EJPE7/o4hyvL0UAf124XF5Sv7zBaSGTUrBhXSbiTUQ2mHgMUksm/hkGmsoi
Ay/EazCH5c7hEM/k4hyqQZoc3aoyWoA+sTy7bRC8/QgTG0gaiPfrRGn3afBrQIjH
gbkmla5WL7cCZuv9b5bl7jWKtO4u0PjnjvRX7MXNj0a3G7dxsgg1D7iqrrChKWH6
CKVlEFTwLvharFIqNPzIofJdbK95LQQUpHp866sD1gXsxA3SUhCE1Zmk1Sa90ceQ
/RQhT46GmsIVDj5+fbzFrZB3WxY4sMXffcvRM80XVHBdTwpWWn/hwIew0VUyYnMg
wpgOyESyFyAsBe1pQjdHdo1U+c6xXWV88+m5acEWzlxrS1JPY7ut9OuJfnh1fttG
gIYCuLwOuNZLqb/CCzy/NuYqbxpYL6AVNFAlr6s0VbbYmJ0T6KIfr7/JFsRVsEVa
1WZ8GEE4VATIlqT3hVg7HHMkBhk/ATTVhMa5lADJeAVqEAVS1sYNcCAX16Fid69P
cr4mgcIKWGl2qkKZVFKxn/hCI+xE9Q6HOt4wWsH44HJoFRJ3UG0Nmo8/wVXT9x38
f0tgE7DRRrK0la+nXsJ4CohJHT+FAscCaPZXDOP9mnzQS9e2fEpWKVWXM7N5gDUS
fwgtNBfCHyGbmYZLSDFN00+QJcp+NasPjPBXQKYYOvdoLCvOJ/0bpxAUjrJpHNub
aQ70lPOuuLD6oqd+60DOZVVDo4oIJo2kQFWpAjv1P1v7w6ZZTHhhCFiLrddj69Qg
zqySBvKPELo83OPohRIi0fnvw+54DJuNwjCink4s976Jd9Jb6zgluKD3xysMf24I
W7NyvFnU7JYlXkqyonbp15+nFD3172t3LnHOMa0TQA6v4aI/t5QaRkJsA9O4GQ7Q
J/6noTcYFuCE5PuSqLD0/n1Fl1vMz9ZQXwlna2F3iRZ0cL9+5+YO/RVmelkpp9jh
j9n0ek7BzJp856M+z+ec6GzjY+KKjFJuJbqHlroV0OCgWk+0Dov+NcsTaw+ZQjNg
ikJYoEI9W5jqxpyCUYZNwYDTbGwggggRPLmmBQaTqDNerzOL1LLNWoeyyrtBCkLf
sC/ag/lpUS7QaP79Yh5KLFYx0CS/GevWlXCoRQg4CUhuTJlzvfRzTShrKv92nhAv
+eeLRRc+d3TFxNI7zepbwx5CMEdnWQEs8UYixHeU+wgZx9JrufHeYBlOwjAqV9uP
4sbNsBO1WfKyCiy26daAo8GT2r7PIZmBrf/oOC726PblSwBLj9jRK/geMU3MpyTN
DVdl2UZxfYvTMXeKN5WLMKgmbTE7j45EPnwRSpo8vvf4QlDl4WbmjoqsQFNfse81
v4jlk7x99iPlWmJGWjGgpUADFras7WeWvf0EGWYPqu02XMuJ0iZ1rmP3/G7S4uDv
W/KyIGtDSajluCc2lLWuOjN4gd6aoIP4FagO/dqDvfv2E5kkpOy9dzmMpUEo7SXd
rR+PM0eFZKeHkp44z+nqLLCjq3stHee9189rGJqASo1vZaGHVGklG1WNrEyHRI7Q
qmDZ23zpRP+Gr3EKjFAt8bf24OvlPmz3zt2M3d9ojbrR/fFsQfwjtdspSZf8rA9s
mr6w68TEpnD15JfE7x0zo0c1exmRxJWu4ckqv/Dpt7UjACEE0eWlkpUpsKosRfZT
FTYukoHYy/q5GuCl6pWRltECRWoIfKtyFXaadUZNLLxIQ/WKnyKabqOpvUeUACut
82O4siwI+ju81QvgSoYVuY17BAlhkeD8B2YXr0Sy6tTGbfH49WFGTX9WBFJNSdBk
fvKJKlT5LAms8utm/g9WjX5ygLRdXfoM2iqZVJIt0/D+hixQDUf544vGNZ1VjuYQ
s4dKDjX67pVyjfbnDfenhXfPRKBwgInOFxFRt+Y7Kh/WnxJ4DBpFNOaE+YMz3y7F
e0fDsP9naSBP7w8odrceBHZLs2EY9fxvk0CzLV+OGGorgXOF73BXxQMH29K0X1Qh
3X7ITurXzJzQYZWPDAC9oNlINWLvqOpr/L3zPYpR+lHIbF2hw2xEFE4AQoY5hPeZ
69jFgB9u82cA5MIyswEkiLVCsYXbjtinnZEsekWKDn7cglxTQhIdpqFqziVn8+E8
EqCGXlYT/W+bxH+ei58zQY+ZwUU/ZXfIRAfNXZ1kMZteuAwEpsWYIKkxN6xKgXS6
FZ2AGSiafdvQXlqircTv4Ttx4iZ42SaR6BdQ3DfuxZGpqOeF4GBPBXEad4WVGua2
CsNx58vraZ/3Dke1BD0ZbCoc/4h1KEjosjv0yKzNHP5nBgmNrTki3IB1f3dABCmB
G3XAHm0H+FTtTDA51dtqytj5j60b/V/IRjfZ7WWPnpNztfDRjCbapvDbuDrFvfiT
O2T1c9DBK0awF1trwEnJygFkwkwzzsOEEDFJrunCVGz+ZWz7zjDR6T71x7TiPw9j
SRIXd/qzLHiwCWOEkgTOZBu3sJjIPTNW0780CaGCfnZk8C8sPVFKSovLsOkG/hUA
E5t1CTZe6rn6+KIdSxm/kJe9gnOVnnIUYVBCln060VDaO+yNXutLgqdaKE6GCK0K
RG+9lxek1JXMXzgRcn97IVpjsvpfYb1y/EfeUn6hV7qRel4F8MEUy3gjrZzihbzV
xpf2rf+dogSEsDODLWgwV/vNjSX8G8gzpB/xWeRvvRQq/QAMCAQH0+/pFCluZ/B8
YxzcT/5ubsuMdueGT/or+qGPwyExiHeAVXklaXrGTKK0mZvnt1oibUjOp0NrehUm
v8qSnZycU04L17BP33W7p5nqhg4RU3DlrTQqCsi+JTzoIifS1r5aSLCGmaXRJmYN
4ogHh+qSn0L7mcJIZ77swOg8x+d36kC924ZFH7vkkVaBXA72+j73URuATDcvuwFb
961HN59vUJppW7l9SlYPpPoTIsKRlFrrqjxHbeTecq571wvMuWfssME2PoqAuJc2
LMmjPDvgcDixxvTnz9vCDAUq4BHI1DWha1q7sxD/s2jtAPe2mX46RjBXAEGkRDX0
C8bHEFGxkMlUnIS147YJ8QOeAlmAwWwd0t9uOH5kreTMwKpPfktteb5NzLR2eIYu
aukui9FsNL+2EJBkfCn2l/WcnTf1Vw/wRp3wN2SdrQ76FHe0qxwirkj8lDOY0jCo
BTTq6QoXmmmpPNyMtltEaMEe6NzkYUxq2it2RnhUh19hdAPW2GLhYAZA8Y6dB0HW
/l9THxYqS2jE3y+X4eqTzAzoXQfkmWpquSC95Zi4c4ngualUHZTqQFkNH36Wafij
cqbLNiyfvKTNmn60rwr45vw9W6oqiXLG2n/PnyWI6yY1HzqkF2llANuIaqQmr7eZ
d4B0ScZ6q6bQAmXATVsM+/mfiBxKgJNqidtBGo2uzEEJhG9XgwHOVvowi6MsKtQ0
FEzyVmlnf40TFse6178HuJD+s8koAO28WSOpTpf3iB2magc84lFYz9J/4eh3Zv92
4j7YtAmMsIZ5RXrbo26J8TeU/BM9zHCa1LUM6uu3EKJilM9Ai2sBN3oNpQWCAufn
ySBPoZIF6UPd7UsbZySGAKCnhKV8gvg9gwiA1hLi4+TAFTeOX3CDPDN5LqEqYsBL
34aOQH8JsHnA/AVZVj10JM5leV9Ry+WJ6wkBnW6NNOp7kB1hEJVcv2LAvaT1x0TC
/3+1dtQHGN4sp1qMrSffk53EwcUvvbVkUP6l5Yj0viqCfPcZm6iWehb8tvWBqYh3
3IRruG9ahTn6gciVUxIDOWXhkQvCh8cEa54iTkyk2j4EdADJTqHFCvJ0FVu/SodA
d9YjjC9MVCCOchGtktcYsejrRP4LMzbVMr7qigbq42r1zzPN2eLyNflhHG2ipIbX
wX7SFleltunqqdzwcOjs2+RXcPrkkgSn3lD/4cixS2zQAyMBGqhsliZh5CTp6rd5
GPdCy9fkGu4Q68xG/+/39MEujcr6OJJNKjYU5HbbAxDSJBK8uuUCEZZmYWJZnstZ
UKn1gmijtHgF60maba2GJadRc00cf4HAqSESftgwQ1zEJVd5Z/FFmC2Dqii5MRxf
jK4GqCRqcWI/T3d7Bce0X3FK/2dfSpN0Rcq1JZHfISn3gsQvoJHaqI2YAZYkH9aF
lkQAM3JVMcdTlY692a6x+0/sRCTt/XJiDCuA6VS3X15aA2WC21L+L30xGty5WNhN
ZqfMpYtt8640K62+9tnyDr4Y0pW66viszLY8BobtkJNxAwIOOEdEFifd9vHI7O01
flgSULgWWSO1vlnQ6JA7SZFQMDtPqCckJ/XeaPMciSBUqQUF9u9yTU5LGa8zpvsR
CqXdW7xHa96ltb4yCDxqDdr8fwInna/0PNDH31Y4I3sxL2HsZDYGdAwI68YXv6sm
tWBgP/TDSBbZ54cj/+fG11nKf1ny5uliBSRvCeXpa9zqU+UbBaHlTsuRuYBrLJZw
WovNd0bfXJfBkcZf3C363nHYBcuVG+Lc5duCqEeUUuFCiRDVg9oVROKfujfjfuG0
sMdA8DGbtncFmV/QLOUmft8cinZ8abUrAAeJwIKq3ayHF01ZaHNgJ5vDP1QIicbG
eNEq8ryoYBkmZv0i3V32ZUfARs3KYwVdQox9UyUSfAgNmmBB+lL7sTma1lmE43nq
rMkqkhsI4MH4XtuPlSRHqJshwX3WaCF1OrUbRAY6KIW/xYAnKeGv9I7iwsRnwHvy
cHXgQ9NdY7XYT/mV6p+JuARwM6xLj5Qo0KPwoebnzTCTQ08JG0v2Gqu7HbUFhOu4
4LsfJrm7lcc029HfhCyM7xtLEy5b4Inau8SyUPx3tSdgOlGPCfqTRs4rjHs9Z+0+
DBindpKM8+kqIVlXert0MFq5TT4/8nYtlbwbWLJsXrrqHB4+pK7s83TG6bLOIyRU
JxL4+JOo/umdybyGriGRhdlIj5yS0vy4z/ifrptq8YToaOszXHJ0XdDf1gfgC9R1
N4lWaozi3miyCRHImlGeAzMJoef1wtT2bv/WATIhPh58oeSTvUbgLAIMdnMJpIqD
HGdFLRY7nCfiijdV9F0c6QJFdz6dtb8ObAIRkI4LRUTn/SsqQMCYnoY5phFw0wIn
vNfBCTdse+7eHWj+/mAeBtcOqrpNx03qLgzlDzaRPzbS7xXfehum+56qfNlqDvk3
I7Q8ha8rC5uj7bhJONz7v3BQ28/jqQjq1KfFrxv9qyD8NHm86eMVB0TehF1Fjf13
B9/EXzL2vz+BLQ3BBoFkGdBVzxQE2fQ4MGnEMEm74EcLo5VWeA6943xuHM6WhZFx
qTYuKrGfoBD27rPtyz7uJzQ4oiuWS5AQXh3wJHIdr0QRLmOxxeo36zGz7Jiz+w69
W42f9RGEo1St7PO9e5bVdvMCfUXVF+OBlU4MKAD+3axvYoURoiwdot62rgU0TIV4
8sLmzivQeLLJIwTuiVesCBeOW7BLVotxsaXqkC7vwsh8TFW4PF4t2WXsMxTEERCF
JMOC9CYV+f1JI0ft3dbKiEVHfpq/ACgoj01cOc2v42XxsgcU6vSCQqfC5Nn67Dy1
rbx6AyHQ13yL/gs4j6Ldf5dyMwNAK/EjhtMOzFnK3rjUlTGL6M8i5nHEUGEctqiy
1ohirc9F7MkDLuw5S5Oh+xpBWSF313JYWVgxnprK6l59AYzhBaYkus8SJW+NHpjg
rGgJQx7BvO11H5RsKCTswcv9jaxvlzHjtVSTdwsk/tR1oWRgF1HOXvvFq0Th8HSS
K1CDehb7IlbWqLIQUcVNoX9z8ESlV2L+247tqDdGun05ZLTbajefijxaQ/thUjac
WhTU5bQ2OIhb7a8Bmd6sgUmgL921qxF9hJpUR1KphENh4sRWsPjkSs5RfMoouSo8
pf3ZbbatX5rcYrajcYCVsForUadXHJWrEZhmrAYg5Dy+Q2EMllrKmdA1ekzD8nR9
6c0O/y4NlK+CttgDBXffQ7C5EMMfJywublWqFbiSk1QVXmaCzBBiSUuHGVF8DCky
/9Is1Y8kKMomLdzwqvRTCLs5KyJ7cJUsvykvtrTw3T9i1XDUCqFWXDqapQ7V54rK
Sc8cVBKiaVUdus2ul115JVPGVbuRdu4mtsEBXFd40i1azSQATeya6v4gg+ZEOkqw
o0E3I2JQrVQB42Ghipx02BwL9R569+RcnPttgyfK3by8RnF9GJ8paL5CBqgRuAoE
8dJDLUjk7k3wd5Kpb4nL9P6QLpDMnnFLkDerJFdpsbuppek2XJFNe+mn7nAVGDO4
dnDt6CfVJU0/kEgWhXhaZa+Ua/Ws5FFViX6jqa6zvaKBIQlSsErP53awUaf/srjK
fWbxnF/sNCuVvYH+N0kgcQZJz/vI77orMKj/m9NyLKbLd1fU1vvVKUxl90CIrTXc
WzqEIRe4S5zM4PYvOLGwKsvlyHQozYoVEbNBdG54zCYiyEj7JTGROBxVcG2SEWO1
Xg8CEUEO3EaPEhSLwXYbcIsGs8OepB8RuNYwp55tAHgotWe2RWHVsmfKcldqX7OQ
rLwJZK19iEQCeyZy+QkJkRTgCJZD0G1yLsWJ98igsF2AcFMlruwGGkgVXSS6iLq1
iWW75UfSnvNYkjYFr/524UOP+wMjE07Kv0tmXdVJ99im5lYurjy+8nF8oQRJBDo4
/UfJEeVfRXQEZtElMkxV94pNZUFzc3buFC6kjgw8L7HTJwToqRnIF4cwO8BM93T8
9S+1+Q+90D5PsCXp0S42qCPZJ9dCCmxmSWOpUY8rNW5XkTInQ9/cVaDtXWEFknL0
kRq7eJl3qaoW6Pd76DU1NyQA5ZeLow5sXreaYLBZZD2wXQklCJhL9PGPNY4XFgff
x/YxPFuEJP4INfuSWVMp/NAtaCtjqFBNVVh0u73Q/3JEIKzuaqF2URC8ctN7srgf
2K+m7GDS2oGKCu7uXXM12A+/m0+nU+vAKXq0vT/zrtFY5bNzxfuL/Lnmm6UZRN60
UMRzK8xzUK0Hyr4WZ7UtDxyBzh19uB+D+N3InFBSkLQhZ82X/ygcfojSpK/z6rGI
PygNxdLon9ZC3LFRYxUSCPMD9pwS/nLTb+f2y3begsBJsjqFdIM78e2gPjXSnnZw
FFjdj9ZIkGt576TrGsdJD9oCJ4Fqxv36PA9/KCIPEqTZPqV417k7lAVk/VGsjxVa
dbAGeQjbi8zMUtvBJ8Q5XsvGioGXvBPfR6ycSEXx7uoHpBUSqWeIJfAkNu/+pyF+
dO0bZYM8IqhEP+sKDufZqBJNlTc5oo4SbwnXmU2FPtIgxuVmNFUFfD3WBPLTc90W
mO+iUdm2PAKZwioZtLw78iGKpAjWKNC6Y8lasd6uR95DBi92pwYUJUHocpi8yr11
LCUcsetNH7zjXUXsOHaJnzI3cD2J3QNAUDyulDWA8J571uN0GGtApGBFQn7u7BHL
Tu5JHkf0sQiXsigaqbvlaC3Cp+3cVKpa8+OWSYXvFFH39EsYPTy5lFlXOZaN2/pc
kwHZ/gL+yt7jKSeoQma0iYRFQ6KyNP+xKlOMGfzgWVTNsUBbnNk9Sl5irFcLanTm
ELiYlQp0UCcJlI4B3Pm3pCrd+FwTK+HF94Su7kHBGKHj2ARtAoC0rY9E63og+Iwx
7jEy3sI/h7JM5dThCxicOH1qK4CN13e+dGJYXWZ2Ve1SaChBcL30/u8i0PumJTOU
2KEtb1Ej3dgdTjSMr88gR2a2ghiGWsse05nMSIhvlWX7e1y1jPBNCFk0l9Xt++Gk
Ock/1KykMeGDgT5hjuFTPMed5xPre//DV5Rd1SGPUXtjNKvB10KRVkwheCdevx1F
1ewCMiwllUkPyACeMj6UMpkG8KAEOS0HlJG5dXqjiiAxLNjpkAGfUyO5pMfMzV/o
RHfkN+fhKBkWvddKgfPcswCvHLZeCw8IBaeE1WYROKb+fW774lCmChhcLW7alJnw
HTCgPCi5iGUlbR5WY7qhax9M6XBRRgCb/p6hA3FOdlvLLAlwLW75X3EvJw3ZcSLN
bN5iRi7YAClL5+VCd7ljrNxVq9WshQyytYV8AVoY5gb38flJhErTOwy/dR74vCv8
+uLC7LFUood6dEi4zTRLMm38/jG2VqbbLOf/k6qzu/UeZSEtOx3lDF/LAqsxzEYT
cd00hYjtZsE/1uuOBxvD57B/oZciaj+Tk0TkZZ9qBNiSUscx2Uj0rZKfQ+vMzXxz
YLCfgcqUU+QZ4Kk6Tv8IDn85yWU4jiDqkAL42OZPYphHUqDCL5yVox9ei28V5tTX
fvsVjU3O/rPwrAEYxFoHTP9z2/JupcFVd8ywFzokuIS0Vedyz89DVSnwQsBE7L6z
5ONuCPq/B4lZxuo6iOBiaTEDPqh+kfruetGoKE1O2Mus07DvIQb9GslCmLPbADBY
0EyvBcs1pFAFe9D9mlaXQcktlpmhEGuyHxXB0efbdYEDMrl96WKF0XA1wReUG/4T
HsedHqqCeh6FDFh5EoX5JUCQ/zjshCnobAHdhg++yC07F5vRHCdHL+Cq4UU4TIKK
Uvzt+/AqMsMYwblltcMXRseCo8c7T6xsjZ2MH9mCQq1ySmdJsduA7HGdpbi6MfE/
N1gDrYkZA674HGX/Il5eDLlT7v/DpXTFrzU0sIWr6CGNqPyMfq44U9twA9XeW3HM
/yEihCAdn/7g5NvPdRhI9ItRdkScHe7qd4lFi4CdgZXv7K20pLDOsUvvMf35GVff
tZsKOxRLBLoo033kVuxt3U58uE0BP5qMwj072575R6IaSbFMkEy0Mcd73AflrsDQ
IvWxmgcLjtaxolZJV5x3HYmhCObTaNLSu7SaI67jqkSN2oOgwFSR8refGIw+op+s
7BN2OXkeVaQN6aM32/xn6f5UsKOv60+xjd0BOpc7LQQ2hrgDWPOkRYt5TB9QMPF4
1JknZ3eU/FQrv294uA0ikw+DwoPEfk9gTdRySYPPElwrlDv02OtG9Wm9FzP2Oqhy
MPK5zh0kHNIoqI7Bd4Mh0Uqou36gt4CmTM/GLPQ6nuIXd7BE0e5w5u8Soj26JMmG
KlWB66tGiUPq9ICOX5DZ14MVxRxgOiw4jJQoe3KSJJWqTDxNdXCX8IYcwGT0OQbD
kUQGb/J9Kqy+8Kf+clmk9H8upXYTKQ1YvubHxA2gnZm7x7qCq0isWJcYKOiHujoD
ZTqjtVSeWxnT0NOcTUxmZ0NjI6pZbMU1QvKymWL6sy0pKEO2yJLhM0ehtDTezBe/
qkxHrtyWSwrnw/9stwi8qGYtkv5FdQcV0B42PrgOqRnG8c5Hw8OihsEGGOZD9zYX
mFkNFhpyurNuZKjkBDeewBmBLrmgCWWZL9w1VPI+s332+ioNLAv2CkIBFk5lxXN2
fI2Ct6Cv7L5iODC2WnUpTdm3A18k43llkQuvNoqWBJeekZzgi/1vCJf1/AEsnYD/
8t0eQniZXsBt3jW+DS6swIXXwyB0ofeHfHZG89o7jvvRAlw6VPAMI8f1rsr2TJ4a
9bt8hJ3ACxOInOhWeXjItZPk8mxHApX3i23zQg8IxqL1Fwxf81jRweBoVPpGMzFs
FQhyRVy5KDOhQtdFbgu/D9F6JvF7Tu9vv1Cs9UPuqD9HPz3oZJviERmDqqiuH0P5
61l4UD6TMmXtYl5ql6FqBSMxcESDQ0zaGwJbyHN4vHti/wRqwYR7PB5YHd5SF5AM
9lMsRP8A4428dv6MVQDGztAEHEGlwkJNfykw/c6c7lh6yDPViQqI23xhqSkO8SxQ
++R1zg+v2al8aflFFFw0MZsECYKskk1uGgi0wcCYHsGVG2OD9z4+LjDYqw/3zQS2
/g0qEWEYBwY4Sngj6EVVfdQnhqI0ZToZ2wfet4AmArXZwDpfm6JiWX3ybm3E19Sk
Jr+7Q4AGUw8qdIWIzTEwbrOocogtwRgm9ZrVtOul9rM8FDKg8mUACp5djZz9IffU
5ppKJ9jrDbGFtS0byTClMTisIQFn6kP3CxkegjQHFARywWZ6Rc9gYmLKJeD+zgWh
TSW0CNOXFV5V2AL6aVx25Yq0eUiXo0O78g0kJ3dUGYSoRv03tOwcaOw04YZVi2/X
uRwHw1WtgDqmNWBhMZ7kN7A5rzIpnuzDvBqltIpAnjFnYFLqtQ3VuUYfi9Zby9dm
ytO+qYp6bTTPHTnUCKsTfKfWuRN9HgNB6Yrx1jup0c8QbVp18OgNli4Br7vwSsFB
jjL/xWUXpqfq5h3WbFESijlu+eL4eZZhIS+OJmO2tncTAs2/5ax4iCpXbs1+5dfP
M2fuHMY0dtf3SqP0Z9eXt1ua9VclwiNBwaZtvVC9Cb/GQvGM2vumqbU9LyklwUzQ
4cZT89lcM9o+WGsDehSMN9Drx+3E+bcZfIwOra4/eOXoMD+LgQ3Wfj8SSVDINzBW
IoneNMNcl5ICsLukVvDWlUWsr9NRkpqRpAeq+N90vi46TYmSGYiUjXZ7SImz1vjp
nKZs/pf86Jxp1tNXrLhw/ASw5A/6JmKa8GlEP3lsx2MMSvs68m6MMsyuVrKpBPUZ
xcjSJJZMLkX5k1rC21HY0Iny12uWZF91cIjgthBdxFb6JR31qVurEoxoyMh/8+sq
vR7bduV1R+JyTG2Q5YYbcO/BLmoLXMdwbUrRAcv5qECcWNz3SbRsmDr7S/dwPpq9
/Jf8j3yu+okpMYLuslFOImqLzQpCvPB6jZ4lDd3n1FZjBkdEK4WCY/EboM/bVwfr
YENp5HSqxOPBjnIQRFmLf4QdWY+uLztuTwen00GI9hrOYsk65tyMeclgUu+QgbLl
QtBoTsffXUlvLr/mizfswwLE0MjjhrukloxEXcKDRGCGrJ7RK/ym+r0OyGbQipbl
Veu0rfOj4pFE0mH8pcND7NMAw8GQDNrGCsvQURGrKX8vUc7JJyuaxt0XjsID0xwI
uXJjlE6m8qEhzpXd6nJMDFxLMkHEefjA/8FUU6Mnk317Bw5ntgkDvBEq2DTJEiSB
Y+cPUdiUQ8pl334Qr2V3DtRex8lbrJIwdfKMnzdxMZJo8PF6/P3W+qBDYCRqqunA
j1K/CaPf8dpoICeN0tl8Jnjwq6u9IXiGxJCKRaOC/TEHHN/JwlVoyUTygzRJ40fw
Wj2NSuinE1vg4kPdWM0iGvxBISeyUlQi7YiVwqIQyd6K+GAvxvaZrHgFM/fvOZi2
A5vvP0uwngbjZyQD5nVoai4N2ZR4bZGlRe20+zzYaC5PxQ1YUbi1K1L+cRvsxpeE
hFBKnGhYO+uwW7NfsHLHeKZsJ9YoMDEjZdZxm9iUU5I9Wo96hfi2b/RUnuaasMvc
ExTQf6jjw0C2ZH886W3Hy9LkBATArb7a8WEOnEIJ7TOAmhyPAuFz5gbTWb97GICn
dMGApPbAJmi4QrD7YV+/Fx4RjuMrWQTd6MgpYOfsNKNG1rrRxeCn3B0OSkGfUTsZ
pAvsgHXInM9WrvEb3S4UmnyxejGgKofd+kcv6p86O0nmlw9X6zlIHmJk3Ui3sivC
xk9tcqJig+QzbWmdYCsZeO7f0ick0KpKA4X0KONvHkZ4mN7yq/VjD9nPMjFF1DA4
nMakjgl63btbfXs16OnRSgRh2bbiVJ3SMY4Tt+BwwV9cYqlkhGVNhMJ/foFquJjH
mK0+EjC0gvMr21QtebTlZQlEywp4zmJM5Krf2QZjV71MmfGPnfFSh/SeL96t4uWT
iMQ8c+7fAhlEaYErlgvTgSlA7rOi0i8T9V6c7Q+F0dBzbLammBeiDX0fDKZrXRxv
am1rJxmlcf0NwithMH2yOgVFnfKEAKTF7oVF1ufoYmPKeXjY2kTqvOiycgKbDLLE
Os9JjCR9RY+gEl36h2VRPSm4IIGh0R6BjbnYYvsmM4ao91tcQYK3jjxPMx053MyU
v/xEkW9KFoXpiafetANL2544KhZpw2xLOdOOc5WhNd5lfd3dSFFrEFfpMr6P65uD
RKjoO5m/jw26u9k4gGHfbgoyg/i2U/QjvETC2GaYkRDRNd76FDb7QDDT9z6/oBhV
MGv0CpQFfyaPqP3Hlc7hQ5Sx04JtpaBXRda5dwGhOTdoLnPxNT8LZxiOliK2nrlp
905ThyZUUUp5Y6nSCvgl7JRotGrx0uiBFDg8OhYV/GfZjYDHjA7wFOkxShCA/m0F
MzjxHQ5mB/Mzg1RUeHRTxFX+LnqX41wjqXoLC7RJmpGeQ+zkutc5TiayGmJm/GHZ
xYKOxhzsONx0ldDy8ioAShQhL4x3ZUWvppph5w+OMWscOr6XPaI0V5UqMfL9h9Ip
LDha3XWgRV2hAx4p9LBpeH/NlauYtIUWm+UNm04uG79PaNiZRW6encEqbHaTnXDa
G3u9r+qczpz57v4/9DbrYsJmUymeuBg+Q0982oaw70yuJRWxdRswxKwE3rD5IW4C
gQbcp31wIQynni1NKOMBDY0LilurvcqVFDKg+ILemLvprRyN/aE4fZ7YyrhBo4Fu
MIHdpHezBU7QZ80Af41Qf7lRm5JsGh6LmiY9QX9WDCJSls11ofq9Pge86KbC1t7b
hEls7p3/zn0CJaWJQyUECwnmMQq1CC8DqdwjfF9iSiJEUP4X9RvxcKkFzCtqCRBz
JeMTIs7yD6Qh9vNiUPdVb/s2xUantnhWXQBLLeDBx/wlv3hn5LOU5TdsuxiqzA3T
jWL6qNMGvRVvidn3X/ukJRxC6tjONLSSDOLXeY44COtkGdNstGRbhPOalHIVrAee
C1lkifO5lXKtvqC3lWN2rZgv8tUTOARFALCcRHxYEFKWkRBuCH18F4ALOQ3ttDkX
CX1WRq5gQro1UvirPAklZG9CbPi2+GeRhYxoeJEi14GEhjaBqWY9HIKurRlN5WVM
/8YT1yCjAdKeFimmODJQmnTW6lfDoQo1IaOOs1bdIpkrRP4OpVGemu2tLxEBuUQ/
iM+Cr5Vuc5aa/aQwv6UlLr7g9aLid7WvkNp9qvXIIE1u5SbuY8YVtq2PfI1VDpK7
CawXGNamvnrvVqok7o2LZTKZzjJSwv2LZ00B+rbbo2U1xZrSMd8833AK5OcClroI
WK81TxLwPjwvzIz3QuCv+7YSknD0eF5rsigxBp242RXElUO3KcCCCyZyOvzlQwS6
csms1kOf5YpBA64x6Wv57dlkzVwquO+IukJaatwsbs7ck1dhsSCG0Km3QfQffVeB
4U/vxKZWhla0Q6AropRjLT3HiVAYoppa2EomJWtyUbhuCwS6DlOEdXElHI7/0tSM
gRryqNU6YatDJEe8dFcxHZjMVOryWIcGaGxW1aNP9HsIb7burzO4nVgUzgJWzw4T
5XxZDAVS4wSdAmGOCvXULiehyNrrvIwY8ZnUtPYv29E6lVRIytzTtcP5MOartRBF
ckkSFHpy92IyJghFJ4ZN07g811GuS0KYDl8hxB12q4+iRuPryeWryNFpzMlVvWGX
cIIv/mz1qIwegEYoMgFdC2kn1HR1Lqqx5Wdn7Nc8GMSYr3Uo/kurRgFEOhrMF+JU
K9a+jpw1KgW88wjSjC50I7cKy2Lj6KKkTYV/Nsz61m62O8o9gncttDmbiuMCCj4s
rAG5YhhEC80IV1Fx5y/lWPVFRtrPGhB09TNNTpKFlbCXjE+Ne6MRlH/FRh1uu1CK
wxm4yJCaUMnK2Kqvm5xWPXmB+wcgZRFhPlQYRHw2KmIBNwxDAsz7Imbu6p24zveD
bxiFc2JhN3n71LgeyUi3ggjHARP1maKBVDaZDGA/B8RwNbQL3xSDlzb2Ndr8EHXN
rv7B9Dribmq7zF36ucsX8u/6dxShdwBAgtfyxkZzoonzmxidY7H9nZWgq+Jpnbjd
PhKgqTsZ1g/Qh76xQtlzQhKpQ4tOoeZfOW9J5EnwSjhhBk6EkjMJF7AooGJDAEuz
xVpgtYBOjYIqCdbtTVygXjnIZJbSTKsC8okuZX8G6IdtBWyZ8utk6iINT1EeV20d
ysKIKGXz1VubrGd8WjJjL70tHz2rOx/IIB20olWlWQx5J2HzbzxoPQBh4KZxQmjj
q0zjocV8Sk+jOyOOQy2wDy685sm1VA/UjTmdl84pGCt64McqEeSyhcK2SRwogeM/
w1LiuugjfHBX3HKAmfQ+xBInFcvQT4IfM/3uv4YKrk7cGH47zV6Oi+h3jYWrH+IM
v6x7LHeF/0Vsn40u/xxcAJFVdv1Fap5H1ksIyBI8lLjFNPB2e/U+wPw8B8QqCxwy
+FEoyEIU3RVMbXxrnQhU0GUfjZkidNyc7HqMgOjKny4JasV7IQ13iQa0XCFDmASl
2vwcscKMTGNtOCY8x9zUKL4ANDLtW9NL2mvri1/LuOSplVSZRh2nQGTCgBxyZC/o
+e6z/oUubTT13DcMpItDfbRBtnmq2hGbcIKBw2S6rAyxXxLlm31WN74qugtI7EBN
YmG61AMxV0RC307d1JAbRLL0Nmw9PKU0PmgpPM0oVuGTT3Mx8i/ZYuuSC1QIp2f2
UxRmKalDpuQsJ9taa4SlP0xCBACCe27QB9jFk3sl6CYDjntcJ/JTh9Q9Aki4mRcW
ueJQJOBMwjspeGhGlsdbCaZzJ64AuR5B9i3ySh6LNwZK0oba4ZuOL9zZUJDxqub8
bbAQJofancy1pc8IFJt3SIUjIkTZsYchgYgOzcn90cU7DeH25lH35wdX7ipAcg3A
mGuJo8Hdz5OS80kG2LhH82pQwFBxfvhC0NAke88CcUn7Nhya3FfpikMGwDGwNf9g
V6BenR4P5rv4VOKA7egSGYKoHCVoQWBvxGNuW5At5urjOlX/8iwl8wMNsw89dFAK
kV7s70C/MyquA6FponrNs9MF5WQewoi0IHPlWgSckWsddRhhSOT26fx2ogvJBwcj
So/ZI3m4leFZQvSdIvPWzNN2QdVzrNWBisuYDYdZlYVct9dGzk7pPIJ+gReeBRHz
QCVDEtL50E61qi1+8e7AxS2qzUNUHmsoa4HQxOAS8WV8bON5d0hI1VBt08N3UlGT
WP/vT6ylxVLMreg+rFGeG4i6fITPiGBH7MEHH9HeLn7UT9h5NGcbMi+pNH7DY0bJ
4p6CH0Oyq2OPMo8FI60AtHK96bMMqe+S0lHRjr9U8ADWVOF5q981BAPWI0WXv+pX
X2DJqZlCQQObYY/jpgCYEt7+HFOUQxb6LVHsV2SzMh63C704YTXpwtYLpDoveslt
MqzhL3eH1bwrclRMpyw085sFMQf8MLNYekyfclGmtfGh/K6UhribcQsVwm6pi6A3
gsBJOS17P2DQsvb4m3168UqNZbLxfal5+lZECQSl00sHMiS0qWTw6SH47hHmZ7af
Ni1xiCJ/x40YU+DCl/cKDeenD82aukbOuYt2VmsOU+PRwJr0j82D4KHwlHDR9NZN
ArVwpqs8q710kKFpPuZAQUa0poNgzNP33ymljrGUdtTCRrwzuvYzkF7e5EA/ApRH
qt0wa7zVIHOmqNkwqUp2pTfMfdcQJJq+362a4uZARkwOGaBOospfNp0dszR1nOJs
pNFhMBVWsZIoBswYplTlZkbyMq7554URitUHds7F8UnVbmKnsZ8dmSy0HtOi4eFx
8UCZ+2ljgMcxisnqXkHAQHhUJYYbzzAyXDL+EPjVA4u5MRUak+GGClM7QXkr+ddD
sCBgXYU4kdIGkpB8Xp44oczgjW2Q7XG4kUQxmfchbtAMDWOJRpvjiihSMejHbcHa
DtempR38irWuRmL52plsQo1uBeVfousjIHuqTxOhtlXmDJTZjqTnQ7pHoT8ijoUq
GeQs5VVOODhW6vq+lKzwy2Tv2F/JXsAUEKHcqskRuaPIy7R8QoL22WTbOh+z3VJb
dEAiAEzieATS9yOSQQedymQyK0pJdGzeOPSYf71KCdPcrE/Ao3bN+TxoByXv91VQ
kGv8GyZOy3sJdjveEzH/PNxUHW13nY3/ltOce/V7TAIEsw1eFWPqsRpW+/nMA4gR
FQuAVqPoCk4ksha3+wIEpxcXvdFXfCBISqgPt0C4cDjNoSeM3T/zHu0BlNsm5nb2
rSHybyYCYO3MCeNYLRxGW9kEJ1Qao5yF7fSqZOyFhRnWsCzwTqAMo4pKtKkRhKX3
9FKU6wYKKYdcdkCg3JHIQDwz8Jy0sXj7Neyv7LEUdFfchvwaeSS85ectA8AvsbT2
OU6fxTw26uC4DzWGPgcO9qbVLVYVUL7HO4atzgdq/0JlXpCfI8QSOL2yOatpn0rc
tBeD87eAsV64Hfo3Wg7ntebTTSAo/L72l0gQ8s/QWM7VZfDTYQ0Fu2FYzpNHYbtQ
uqiysG4SK1ARrIENU0TBhYRNlUxnB2HbAITURohgiveOXol/qdwf+8ERpMRYnumI
uUqhJdi8hLQZo1+sAjU8xGX2/84/6nofz81c5N+peFZJ1IiSqyK+b2cn/frrKGg9
6mIM2vRF6iO0tah7Qi8W04sCBtLJ/7dckKlrDNJQ6yai9CqNSggLS+xt5e5JRAUi
reBJjNgdeXq4hj/Od1zH+OTIH3v7KymA7UMmsbJL3WKCq4fSY+2SHzTvfaUpnl+a
5SIo6Uygf79im+PWtP2d2qWxXiBhvBpNmzDCZg251IcMIK18VjP4s58WCeI5jxpk
gKQ4c/BE0r1gGD2g6CFJGNEFC1xRTBNmk9qvnSj7u0J9GbIaVgQEw5+CeGp20idZ
Ahur/4Uzv0KYn+MCJG1zB+iq4XpzWaMzL1d2rqlfDgFqeYjY/pUNkgjLrqSghZoF
zJvYYIRNrFuEqvprYxkiNKFZluJ1m4YgVlTKWPbh+2cT8T9dVtAtfJgS2KP7C9X2
CpbGnhdxQI4nvINxMMI+vFpjqn1iHoZjk1UisL1ClQAknyH8XZ2P80BH/bcagGYF
VtzyL3IjXbstMs+DVt/su9tGP/ijGgplCEDOVAeJjF2mmeNTj6VpZXU4XTkxt22C
sfYoNgBqVr8Aw41vRzPRLH3pRO28uMAuWSSnEt25OPsaTHVfAy5mMdoXErsuuOmv
B79vIyXcCx49Qf7D5fiL2q5ziwOyRZIh+ReoFg/gxpgrIEcRgufhtlQbFft2Mt5j
sxcmbC1xeTRTIfQyd21hsHK4GHWrB/XJPeSacS2bkkfnZ9qCPj+Jm6u4mPM3G3DS
CKh4zZyA2TeLqUx+y6vSVkZLPHYDu0fHQV5GBhJQvnW9SejhbxcemfqM70xOXGKt
yny8QxxKWYmPJjWJRKTwEQNieZfvOtviqGo2h/jX6+RUEnCrdX0zqLDZZENfdlzd
2uPW4ZUnqo+UBgBq/FvEdHSgTFmPGU3htTZkZ+RG4vgCD2LP/uSg5ZDIIpc2ez03
4WCrwXIr6+yzrOyQzZhuNrGNCIEJge5dXu9ZwFu/cMId9NQ2UNxr50MetzHfj9tH
a6uXOruF7GVOIsHQKyltBWNKUVGYslhQVN2GHGEGi/DupeaWnxPORHphEft2Ugz8
bZZOUxZD7jyrSX/NNbiA5HW27PgS3cwNFhP7rADLeHLuSDRIe505gFVfNFnOv8vk
IDQ7AWx6xU36jlJSVdrvVHdX60spKDQO2meqnxXX2dFrxkI0D9x6XYoSKrvSRKUZ
VtmKJoGLaGKbSL8J6uqpT1U7HSSJP89v9TkRHPMMGmDymEnh4FrLvxJQpvClz48K
tpXc2k0pkAgf5aQgji6cL3+C26S7MNtVZqCK/nVq6x6Pm2imwt75F8fFIt1/NrU6
HPzAjrNvUb0j2GzwqdV/afCJ4MrAtxnd+5KnqvWQW2nbW2Cjk+9p2GkqxyRxU0Xa
8/U3FWsX4Syw+T5gMxhQ21+qh03tp/FNPnT24OYQwP0oztqG+91YjQhXP1Tf3exi
fX+FEKX1qBU8ggOcir3SHFtmXHwi6wKsPwC9yEc83sz9pR7ALznRVY3u6aeanUXB
AjZt2n1yJzOblZVJJPE2SCkkvEFsOka9XJBWSFwbGG6fHuwvDAV4YzKLi7pt1Rk/
mf+5UqYv9uBgxqy4EzMIUCK9HROYJPrhjXri/bY87P73WYkxx0T6oGFdAokzOqH3
4UpXVoKY3ZevyB/9TanZREVfJEYdAS+XcdOkbfWLbXD3/nwKk6kagFd5Qk7ZSZ2T
9eNhYPlA924mRTCnOBxCmEQ7OsTG0ZMFZ4BGFFMX9lVpxvZxIJWipxtVbLVjUEXa
bcI97+aXdMzt1JsO3ZhX33T1h6oHiPvcCeEwAGTmGfGOwRsG2HkMae55CY2zIrJw
zDQMOBTzk5z8XghsJtmlTeyY+xcsBh4tZK5JrpcFrSDO9i2R7Mdae+LoTNbcG0z6
/Xja/S/Hf8jTuejdMETu2PQMCsPWVvfjYS/BHv7GtOa1byFJeZPextsfPmRppgvc
VmTs2YUyEcgp653rXm+H5bhiOl18XWSCgTlEf5ERslZ7mt9GV1KDnvFMQfqLkoLL
49sKJpFnnuuA6imCSZvOSF3h861M7kxXVFQWZLdvGvcrq+A79aFQKmRqli+UYWqk
+RUWfhdr5RCfJN3gXshafEsk2P+Y4PWwGxlWeJN5ibLtJz1H7hGXPLD1gcNLlMmI
9+8/TUCu0kgvYZdrr2i54q00DCmPdZvb53EE5sx20VCgob2jiOww7I6HdnErlNSe
Fs1VTjwPOIADOZYZhEWxVKfyej69DBm8WhnxxrNpPLZOm9UsEnN832Z/sZ+BHqcV
ZBAvR9Um2mfCDIdF/EGLT7DiuKFZw+XhAT3zCNnW+5cNY+Z2yw7Zw9i6dbWU5pW2
dwgm6cGBDCTyTSvoSwpfdjlivFYX1/PuXaERn2F7zbdzU8fyXG8iSumqUJowbVqn
oaUl+2kNBtNrQNuJaVshp03Tor3IZF3x+kNR0hX4MmgLq+yZlaujpxzAPgHuEltR
eTwAj14pABbsM5jkFprkcKq4EXeE/f0+a6Gjf03BVwAwCUznpxX/vV36H1bYkMOI
b4xBXaW9LmnROvu0Zg5455VzCBxck6f7rbqk05sbZHiFQe6yBjk3XiEjSkMWR8WG
Xvw5pa53y1lY2NcO7jd1/UMknAWIjgJ6GY9f1lCQR+eeJAeAKmGVkv/URYbfL/ve
E1/jlqHnlEppko21ZwaQSSrdsOm+gnrv6YE7EkWmEUjPsqyaP1MzzcTrJfaxq5YW
/8ZRuV7wFLFXomwV8QPf4b7tAcEvcaFBJVvAJGc5YpKM8deo+Qaq3m8+dgmAp3mz
iuo7lANgHHUEvg1MV1XOPzTwFhEuwYzGjR/jyIdgWx8/31dns/h0LtIEgKgwi1J0
CwmtjUHOVrNHjivnoC60/aLmN2NkgIKDpp5PmRHt1myS8I3zQv0JfGbRZ9TXulJo
UztLEqBRyPB1ePKvIRAGXObhv+cBogCaAGWoYb6/QRTlOKtvpMqA47ycpqsPXxt+
yNMKC5/1nmCqIhuKq4nGju/2xY1/5DIlMX+G7BVCOlP5YHwEJq6bpFEuvgjtbp71
514gBJJdfdR1b3F24Ee6Keq7iaTSO4qpraZOcU/ncH9ZCBk2V1tx32SgSvq9V3d1
ySsqIXrMM+q3hr5LUQI8INNZXwG7/29iiuzAVk/+qd0Y85cTWQEgMJpcnjPtbKCm
myjmaTHFR+y86RZeZ5eifsZTNKD/mwdc06hez1SCgNpHevS3KoLPjUevveq5+Oqj
N4f39qRtVeowOeBUc5pWcZFAo9XYP9ZCL7b+LUITuFCbWUg/XNxqrnMa0UcsGiFc
WiTb0qmHFniU97ff8v4fFWRh3Rxj1zkK+tguRZEPh8Xk2glt1DiVzBxcmIGJnQEQ
5O03RxLU4sxHnlZMDQyTsu6waNsF0TN31jc/EY5i6rLq/C5SVzA+1JYXWtF/Gcsk
O8EngVSt+zhMxt8s4JSBHrGtiQI3NCjvoUaU0+1MdMvwnV6mqx5ReGezVIJAIBPM
LoMQmlCsT15/4eSdfZOvZtjXh0wd3QdquyIi2tJiyqkq5wDrl9+QL1uiNL5bj1WX
MlLNzH9QmWksHc9J1Cj3xRWE1ZNVgwz5L/X4kwwRbOzPjn62xDzj12eLqcluPpeP
zijzZeJXhdr9hTuiIDufcI6t5Zu/XZ8wFKnOJ08Qp6r+PH7hnzFSTBu7uajROyMm
9w6nNCCYT1N0OND2XmkhQ0ldoMmakNngYoueC4MGe6A2WBbQGQkn//Jl9qaH4lKG
4CYE8p9+HlXlYJC15khHO1YUByohUWoPwonUosPzHLw/wSwBKctxMpKTqQTn7Zri
gU1ksUppPw22CPuqhxxKQQ88+LT10YeVA4HGWS8aeB5XSpwKgUSvPMksXbT1GhRJ
8M5r1Bub7+d5CqwWtStBC9wE55GrcMG8Xm3AEFE/RnDh9Vm5IbsexsdHeIBN5cMY
LNLkQgnu4M9EyXvTJCMXFnRMmrn+lPFlBhsMjlsEtwFlwOU0weNFv1kdCqfN6KQ/
2P7nRyIqylHCfltO3ULfFzsIfDMptmiRHkdFt6fZyckVBgc1dWPhNk4WIzyAWA45
68Kw0QV5yus+hmY0WiaWptrcRRPIqlHO2mst/GerKOU4P2ZKVWWJlhSlrLt7ZIdo
+5ziLJEN5lL2dRELpmikQrbe4WjPfGXaAHDHWnZjsaWjMwuj/jZ/lTteYv/pscgn
a80B/b+UeVHqD2NfHZBIzhpQDzbnbHissZp4v+o5XCF06u/kl86ZrWCOBn+ewePQ
HTRrTrh61RatAklo03FA2suDNzU7CbeBjv0yOTpcwjP9RdxHDuWiGM9b0CnfH5Pt
70brRkywhp9dneAfoKCXSPjx9x1sizDMkjFRVxbZCm//+YYct+7fbhWUvvbijiGn
IXSmJ+dnwnPtAJqrl95GKKChE4AA9XN/fJ+D2kxED1NmzmGoZ/sj+DBhQaNHC3C0
cnTt8CU64OhyvRtFy6QCesrmohwuZ9YdN+rlJeD766zunIh/yF8eG6MCgrq0UO59
0V/z1gFRQ+jEWBXm2tS4t6m59v/IIYO1goB61Y7zaFWmnZoAKXffn53/tRDzpGwj
5ukXBxJKdV7MfUjBoFC5kxnaytV9x0QO72wbLwRKJUAIfgsx6WUx8e+/PtT0pKsd
9ON87uq7J1NeTYz+3kQsd42iU2oXqsU40t+Su+PqlUhAnXZM/tjpMHz48hOCZnSM
6EkA6nC1g9xbXsXxIdIWGQIVhTYdBH6jRqf2QsNx3YzKrtHZEzAzd1TxdrYojyt5
mtXY71UeeYW0dy5JzNz/PCCjJjK9IKxzQGdmcFLunNlHvS4kuCES1IY5qiJ3u2el
Wg3LGa95LscQ5mOrUd40LUSaS+ysEmLdHRpTZQdyqbMUq5IQclLr3f8hcMZL626n
/JVq3n8CVcJUpmOcaMtZyYXUraXMYA/e+Lfetm4TKENfPE87Gy0SoX7rRncW+URQ
YNnunsf2UV0TCHR0jdOt8pFzb9NdOrRXxv05PPb1DPfJuESIXJBnUtOSOQGt5IDp
UblsJcuGpgYnq3Z0+tOkfTThHBUkqqrnPYWRehJPZ47HC+FsUIf5AkbzYWpPMx7P
U7qvxOg363RU9HozUCOTSUSGKLMYy0IZSfG0SdkAV5U5d2pM8VHXdZBi0z5JopPY
qb1kmz4kD+XG+IiXAXcF4bKqwIymkSIGsbEj5xD1ldDPDOFWquRZic7ctLSx1RG9
8H8WRK+R4WyMT1fgRSX9jp/GKEfV1WGWE9/AtQr0C6BRw2BjLKMRM0UvkD2OMBur
to0RFQiXma6FM705NKpomaAPjPan5zsILN0S5DkGTLxgepwXTHnq+sbHIoZ54owL
KVTD2tKI7hFXBErCuzb8/Q9RJ6QrYyDxTbDYCfVeA8IjgVC2oMttAnqR6ZkCs7rv
DIB1+B4I0LENZ/OYjk1uPFOMPQ0at5RBeWLizUCJvVGu6X9XC6meSwUi3I4YH1+f
yks6EpzA5xSzmFBltob2LSI1FS7nX4+tixs4xYrCgfWpFDxQ40qv4DwNqpyqGS4T
8u6U+wBU8pxLxRQO6hAjbToZIoKtno1Sf8M+N2bCNnPAUv2b7lLvy3QR/WLh+E6x
He50Gq0+83/S9FG5oDP8zQFuYpglwot0TC5uopRpuVZz6KvifaJmIondzUVo9j5i
18OwshtT4biQlHbnv0H5Au42vgnJbQKfUKLxdPE72DCAQm/+DOLS/hfZ3a9YwNhN
eoMio2kO76cx+rGUo1FCTf8hcWPGQdb0zXGf02eidPlGniiFJCUecqHO7DU71PPZ
I5AMgNjnw/T5bcdnZTxJbJX7R+5Gu2romYfTLMUbbTuH6+vM/nw8kbmS52j2I044
ket+ifK11u1VOI3sc4C7AHQJatZhLLUlSF8L6I1a46REGaL1k9/P4uljMThRDc8w
vnUElpAy1+lT6a5SPDhTDe/yjK+jpzn1xRYQCxeJ5XjnLP0Y5fx5YzHUaynu9sar
X/LCxD/VYY/5792rcbMGMTvuuW1sAxZ5sh8ZGlZFwc/DMx6nKOlRvdlemeYvUKLE
QP+IYuxw+KeESY8qRd+N1ggybweyzkkGwSCxlV2aYma3Wutfk6EDR9f3I55qHJgg
6k37l/05KzShy7bNdGjuad9jjLAM+jgdnY6yDMgBawa2EP0haimbJ8fKWuHgWv3K
FmWYFiONcnMXWIpoIubtzzSZyxYeB8ZQnyOILTkaGtckDHrxee0pvnqW+KOpEf7x
/DPolURiWJC+73wRZSxW1l2+TstP6eBrDuhRCfL3/2HkNw7snuryfEFyNkGJaO/r
2mChQti4Ra2hJN04F+xGS0AZo1WLDR/1veVjD8hH/1vbe6FIhA+fGYFZmNo+W7uG
WskVNE/e9iLcWAtFhqs//j0ve9co0jIyV3lKNA/rF7w1aoBNtci/MQBuHZuhcajR
mpW/66IU5Q/x99jDhi1x8sF0BcmpmZfBHmDidUoZl9hAbmRfH9Z5eNRt4Iqqrxjo
kM589mSZwfjXXQ3e4g4fUmziNOcHBcNq+OXRcxMtqBePmGUCoOXIBxgiIuOP5nPC
I8Xp/4pQVO3/oR/OQNhnfCdbfwY7vQI9o9B56YG/E391SToGqcRBBVTLbmliv39g
VMsS2sFervWHhQXefPuoFojm1JFEQdLm/zqTKaZ+iFGBTRMsAq81+ZnnJZeZliXX
bvRUrL8dTek2bw9vscSjcN0CGRqQVo+X2L76J+5GgckMHqAvvxOlJctums66Tbpk
wCXa63QqUOVrZEKNOjuuXSlY0Ed5RolO6VsMUuo7Uy1DqByjnjwdbG1mRxwRvrBo
aW74UpPxJx3HlGF0W9PdH6pc5kKwx39gA2sl0iPQKrY2yqcXLahja1NoFTITvg4c
Z8+f2/g6DVNywaimuo5+4qd76ZyI8QgMc3hJSfdeMQPKiQqzRXFFSP8s8CzsbRlj
gNaheXt8oNVP7RyqvA0gbA2ELwBMMgAA81Mty1kRq8+vVzxj9DpLr88A+e1TXZGS
AiHDNNOxLA9kTmskNYPOGx7mddD54z58enJLolTh2VSvyAgHUUJfEIJ4dpA/BwdJ
1usxhMZoZ3cmYqJzla0XbpGxXQLdgr47buiqIBDCQ8E9Rv7US8L5c8pxvdfUoJxe
OTMl5oN+bp1VZfcoSUE2DJ93MCawuxIa48e3zVflCjXpdd9pttoBInvBgS/rVMFU
ZA12v6vCuXo0R/RMgv0yb9wC5QUZNuQvw6/fCLvPt21dYsWwlIc6SIOJd1QvRukL
tOM2bAFInSyVQBdlmzXGEKqpm2nGlRwvXFus2QIvhkFjclYrfh5PK5/LoUsyBLFu
AVupEMf7B9wdAdMjDmbEUD1wofHXr2CBOxxL8hc/je9X7zrUS7xbkgTMPupz+cNb
H/prZmg61TJKD8TfWT0yEMEZ+s1L2FLajoSzb9Ukygbmsdfc2XlB2Y6wYPQTNqrP
3QRoYks9ATlcV+aWEawPCMuYZGI/5+P3PdttTuKOypm4MyZ/M+Yxp5CUNF21E9RH
cT8k+whUoKHbt8jcOzSqZlFk0xDB6xNOZWhFmgkksbJhvsgB3gYU+L3VpJGJlxpV
Un7T72wGmypq3unId+ACdPVOL6Qq/aLw/seuPdM/QEeXIz2Ztq2Xneoyu2v9ECaU
Y8e3sTR3Y2z5tha4DfYDyisaMcsZ0GDBesqKzODa6g+ojNkiFwRgm236i2RjJLpE
u4crqbYKMc3Vuiw7u5K4mCML8f5zAA1kTQJadR/AKunrco8NF3nVsc/+3ufyGm5d
hdx6iwcyQYszi8y2SUxl9X7S7jSIkLevJOKqW+octjsYN82PXLrZb1/di3uYaIfp
XwsPPpUbpHP5zJbCijcdi4/NjURMOWezTVZmNlE4ivYY/f+/rd2wLBM2xn7eGtzr
ZgHEjC1G4ITPyNcy0Z/IoXt3MWB2fOCuqQACB3bgv2OvXSlDUpCiy5EOiNqpFtEI
OZxQOKedH4BVgaMPZvhlFEcGXenhqIGctS/vZS0+lGK6gzo9i2hiccV2IjbYGv7q
i+T8qNyXrrU8Gc7ScS39W27tmS1Uor0xPj2mODyRO6Ssytbn/scXp1MkiWXe0hqi
GBQrSnXteW2MfMt6avWX2C1TqJzgVPn6QdVkkEsFRS6UBdI26/MDHgtNpho5hm+b
68j45cNpCvU4stjCdI3OJGXVxrZ9+mFd2Z0NIMaSBwrrC7glskAvzbfh+inuu3N8
P6LC9qhE62igaQ+puJHYHlZLQPUS356k/zAnz0GQ19b6s+4m9MCOxqYopbJAykF5
/7kkcW4rF85cpWzOPK+JKHbFy4pqERR4J+R6g124syrIlpOYUp0FONaZ50G+s6vj
r4idhQB5cYH+/Ooqz7HmCE4GjV2P5tGPpV2FZvRRlKAHU7tCwL1aq8K5l0G+GSJ2
oHgu6yxcYx9nlk3ZMCiytod12PDHVqqT9sR4JP4yUZt0AK3vRoTlF8bX5Wd4tld7
7WtK2RRx0+VEfKHWHF1ZpT4EbyFqtwXDjDPJWX3kTEuTniO5vkLfgPaO1cA9Hy11
ypT6ULO1FkM4va1R9xPVgiOIDgxgfZ/AMNCpcmTqLaYzNnOjtTlNtr75mlB27c7t
tO+aU1j9kf19XZISzO+jx0Pfv3lw15+QzCEY+j2dBPhxS24RSWsyPKYee3+ij0M3
gCT+ISP2zYPG+T3Aoi92lV3fA0JRnK4iD35VD5eNy6RA4nqfXqucRu1I3BH4SP6G
73HA/AO98D0QbuWyzxysxwSy1p9IuUkZ0Ua7HdG4FHPBSX44bWb7y1bwlA0hvvA6
74yiiU3urNOmKrkQvqNIxoEdTucE9rVWNCsmjOz3QqO5Y1uOZZ694X4SnBG9zhsq
v3gBI0dBzhlEP1MifiNmk6LsRWOaw8SwI0Et9GYUbOIo/saOif/D1VIMIwW2znpM
bK03BzP30NKZTaV8bgzgrMkXMQaYJKXWeC23/ubKKBUJegHdqLSNKPQZLslYeRNM
SL+HnKqUq+8WGWxyK+Or8CNR+HO6JKhCpdGzqE2GsEK/LotAXzGemWc+YOGZAHsT
5dn6kvPmodyZ7vF7KSJAXumgsifVv6pIE7YwmEC9+wZ2DWPVSmIqpmR9s/Tryr/i
MLajKj3q6ID9Z5xzGC+OBXIWDfyWqlWIlqRiJPvli9i3w7y/zLYwzHa2gSkO9dtA
cnBdTAgcWRdQuOSqcIuMXVHs7QYnm0Ll2YGC64j8LmKUaw2jzhHFWXjzmIrQQv89
KlBdadGvVDb3B2hwlf95j23KJFeZJ8lzBR2OySFAOJJyjbQnznlBmoyqgERxqE6e
G2YBfaIXdv+B98uL3GBsfiRmH1x8Pk648sJXu/1Lz2QSg/CiwFubHwHExONjIF+L
6yWd5GtipUm8bvjLN4giGAEo125KjeijbmxHk790z31n5qJ4ETZesj5lFGtv4Zk9
P5e8hOaKqsKuLnpOyF8/l2ZG7s4ZciUdCCM0VXXaJz+IMBEYU4FkX7VhPBrmfsjq
pwe4saZ4WtbJ92RH4XFAUrNsB/HT2GPKOtK++jZndWEUIwve0ZDSmICOiHzZKwWr
y9UBbFo8pl03qGN/sspSuR6N5LX7PMptkgdiLZwRRcUDp3YypW//dbAfPsxLyPt3
SjQigOQbpxI7KBCamBqAz2mjs7CX/d3zLWJr5C3261Y6CwRophp0D1aQJ2N4jNgE
npO6yj/CrinvDljgDZ9UNTG/iv7beZKuSWcMvugvfLR/4LY4eXUn5bDG3PSxY0VS
wz3LiNqKEcNN4Otn+81s5LKkh+DABYmA8rYv2bsUF4ntiYgVJbr1ghFEUiTgTHlG
DAgds0nkXNJlIQrV2a9AUQ1LdM3rwVNZCJTtaqzfJCc0pwGBbJhQrslRJIt9ldnT
bl6OoxKIG8c+kkTWFJ46DqL28RHAwllm8hX4VqYaE0KnB9lWCK7CQG/vDW6c6wnN
IGxqJ6y0MG+hJLCw/2QJuqpJNj16y375pMUYFhqwkFA8iMddRzjc5U9+0G84ezJT
VtWpidyWcBcRgFmOY21CRhxOnPMRYt3YDrQeMJjyaWM+8TNEEssfVuxFDTWGG/9o
LyyNspcPyuzMIhy1Mj1CBgVX0H1LamqTzkvB+b3wicTLPEWDiCH9Xh7mU6e8n3Ar
yy0rICWRm0jvYhOrWKAneuBfq1ViLTpYbrILMNP1n9HKQ12j6D17GXq10eEAugUl
0ZihTIJfAWrVHLselRGXhfUvjb1Ib9Ekq8yiGnte2w9QQ+mbKh3I1P/YHIRJqm3D
rCoT0JsZ/7T0Smq6lYwwsRl61dfMdUKIJEBKLBc9gVo53hzKxOkOInI2DK1bw4m1
2vY/PjIUEFoN2Pb2GSMFqO2Yz7deFb2MvR4RYvrj+XLN43I+loxGcWWJ+Kt9j1dB
mgZBj/YJDh53G7+ykTQuyu+CWZiQsgEdG8so/+N1NgYKlS3A/FOp6ERDGi4op1zd
g+gY/YqfuTZh/aLZVHhlPCyeJW9e+3Oi6Cjn7NQNxaKZfoG72Gv0R3I7/hAeb3Fj
g++rsW5yn9AMw4M7o11NbilBQRcMBqJbq0fBC3hU//8Ln0UMPPAakwalQxbMzdYq
p9tD/0oS8wL38BsNsJFOr4pUZES66IaUcrmo5gdkkaG2medIg2EDAWEGHbo78smB
yPhfrK93RD4nQdvDrxM3Dzt+V77Wknzz2qSlt3fFvi89frMnkcky8UpwNVC15PUh
GwjyldcDso75fXf1DwfgTTHn7TcO2NWcpoOo0jx0QZ+KNg8QH9ZvEyBrPJja94pI
wu+6NmUQ6iR+FDfTLExkQyvm26o8w7CiNQBiZ5o7o2IsVmOlVNcFGDdECRcYI94Z
QcHIHPPwJyrLycMphsy/QjwtfjXL2c4YqhOlu32QIATCEFNe0H8S/O935zc0nZBA
XXRdingvg6bdVyW8SyIX8bPsEiFAZC2TfDUmSO5ra++ugCo7B2fiZH/OxSZ8RURb
XutbJUFvyCYljWTMJYts72Y5R58EFc3e9Ri66mzWuyfs+U8zdvfmLYxpNkHhRMVs
pj39ZgndeMIjihMQnTIDulRSfL/3kevkjrs8EaMQ3jOXjBFwZgiDrdU8gxCLzZBi
1401ohGieCyBj4ZJ0snEAdCH/BraN2PdvZKMPb+kT1cxDsYDRPic6u0WTorGL/oX
aUYssDlNuT8ORQqICtKekQVvzXfPOp1LWqTduGu4UyJu3xau51hUbqoDk0J2Zf8w
crwXwp+qgWNkJLL3Vt5RN2KV55Si/Y50ZokD/rgknzu7OxRK2gmW6b8EcAgNKwhi
E3DMH2/UiGH3qRTNtzLdDl5ocpgzMwAMw0qBb12JxZH4GWczC1yKEWWRCyzH3ppG
bXP8pclLAVHahqU6u9RvSHpKaOrQhlPPn77H9bo72M9D5A/uekX5CNe3TJ/e5IjN
y/jCji678ldcu7wGAXdtvrOZ7sfoxDgNt7IgmNYsO9E1v4Gkj/Xb1ELqO1qhakkJ
ypHcXHT5PVljgDvVF24ysprsz+xxI/Sr0fXj43JSWclfB7lG0GXOJLz9ZTbD1tu8
ZxCUqUr9g6D5FQdqRok5n208c1RR9y7fzqbuo7aBoEZf5adhuffrAbKX3ikxOd4b
xoxuwwCn46LpLm927aYRDQVCJFk3ukp0RVT7oINgvCbxa/F1QtZ6xnjDNBB8q2X0
1K0xN/kM5IfjmH7xJaKIlBnj6VwpnhrpTNXbzSTNjbXGrhxnwSwpJ4RGWHXE8OQq
d5w/OobGvoe1MJIVHKm1qYFgnMGSnDpNRxn46cUbOCXCuLAidMAYC6sphKR1G5Dy
lrhHrlwvSDnr/rrXvaaFfpf5FRQi/7JooOg2gYfYLxZyr1F0PRlrq4aojuDy8NC4
jaCy6/L+DINw9EWb5hLhcG7nVS191k6VVtqVfA9gZA21GZI3+53BlwDuOMxIgNXD
lcIs2MGUiribYRnuvvxYgew61vpsOy3LcS6JNWE42yIyBVR+GhH1n14U0RqpIeZ3
zrheNY1GaL/Pvwwt8hnajdPmCk4ECKD3ZECw6A39VK9TxEvqyPguHWAntoA8KsUc
1/QlJ1Btfn3DhUd2bR0UwgrdCz6anb/xwm0RwfrEwojxs1u43/IBNnxM30SqKolk
2d6VjC1NQXp0iz5r2CzVRL+5aTT/hiMlz/yrVzKYS5rO4dqPTKtjU9XPokyaXv3H
Wj0NO7DAzprzq+RYpTHLd2we8LfgAD2JXTEFJl7A/Us1GEzJT7932voSadnuBTWy
/SWka0fDIeVnbw0pLZ/E2HaFf28LCwYpcCn1vxbNSewJ1tBw8Rm7giOPwW1BgH9K
aH6ELfb0HBvISEZgUzs4HETPeXauLpyx788UJFmWlSU16gl4DolXFGzm71e0e5tL
eXkcfWhAOkaihc3YuDoaO535J7DfziVhxLVcBZOUxtURm/eQc87MTibqEYBEVWbj
icO4P3NcSeXYcqsuAmUVrOoJ7KxGJq9dLryct6h0lpEIX4K02gIFLEu0HlS53ezG
xj0myX49jCHHPu5/oasTOFaEDR5SCdI7jCrd5EJzEDmSfz6AZ75Iy/10HWgW247z
v4L4el9wbMUdAciVOMorGZ5UKFqYMHKw1E3TNOhGgzUJ44pEFaFyWY/Ux9BOl4Vp
ug4M76XMyrur4lQ4sQmQi3deU/hcvgaZcbxNd8MwrRV9oquUrDDizOt1w1XSjjmg
YWMB8ncEsA8qlx01UdMwY4SNqBUBSER5+/RHreIvQIZGa7zTxamJ3Kd6VMq5+nGF
W+K/HVLmQqhE8EIXnDhkoJziB1yyRnoz7RORG/QSKWOtPWU6yGazUPTShMEexo1Q
G+FdB2IhE0xeanaIXvCDjJZ/SaKZC/VnsdJ3dBwIpS8/NcARD4wZN3sZTL/2ZDve
KJbjZ0p/eJvztl+eOW004xthWgoShNgVplRmvn3NfjEJ82dDYAB1We3FpNoeuGaf
ZKE7Zuipoad72mY5GcR56MqTb16//dqJUs/P7dRY5IvBd3GdOf2ozNJ4jGVYmux+
MCs17J7gqn11LVIX4FW46Y8A3TxB7XvONVjLdZ9o7MJboxwi6tihDlnPSF9eHmIp
bkE1zx/RRZ9GiFR0+kgvThgwGJZ4MVRnB8smMTG5iNFjrQa/BodTLYZ/smLL7I6+
fKRnQn1JbNbmgL8ZFUmhTQufkiPvXC7A83pub6tI5t+vkaPeOjlZT0iY2BRDsKSe
ro6bQQFkJ0rC26PjsrALCCJq6UvEn4N+uVm69ij65FEpiTZcVgzNZ1htsbTDs81k
v+vxiPQ+CIey3S8gsKKHpXS/8L2CDZNRXdhX63CicuuSUq0ov7l9kkvDwj4R5YD1
SA2Wg7/6wr1IzvK6KTUCsp/lPByCDzcHFypDIzzovwRAxIKc3cJaoD2Mx4F/T/U2
5dXsk8ZZOVQMrKvi9AGH7FP1dGbXnDQG9EGooewQgR+lfl02ShWxoFD3/da4p/Mt
6jE/K758Q0QIALhYUO3ZvixMyDM4JL1lpRf/Bn48/Cee+qhVUN+IPqR10eIajQIq
VfKcLaN3MdqcEp0cABEPHa04dZPmAC9rKJ//d8T0cpG3pJrERfPM8e52alEA604s
lX4tK+dcMr3K6FiUoLJIOi9GkHSHZbx6Q8EhMzrSiRZSzYr5E4FhFbcK2TGtrZh2
GTXQkG5/2Otg7oBOXj3kf71/xxyRzz5Pp2ESOMV9H/hthcmZyFcRUaToDfW9Go3n
phz+jA8urMqu6nXoCfV03WNDaYtA4VQbGP/9iYLM0jnNaOkg/kC7w/fB5Q9tb4+0
hD/LDeD1AaAhAtUMnxKlkplJETUHY+b/9Uo+J4B7woWZdm/b8Ltwv/Oey0cB49lO
E/7V3Ou6Jr2jxkh1jzhytsmlQIJEB2h1+WQlJEWu4AoHMTkKiLVjxKefgxO8dI3E
SBmiWNhskByLcFj05BGmN3oj+bOBqs3ODpjnbCEewE6RU3z/cspQCfqmqF6aniUl
I66fDrr14s4cJkPtZ+re7akxrkfjaM4xZewxhZnsRb+UP5EakO72lRgwrzOip4V+
KzINdmh2OaXvG9rKD9z4po8RdjxmN4C3vi6UWY6qKT4notWhm5MVJPe7CnzXDbkT
GHi9elEgC3//ejmJkbtdvth5Kmpy1RF65mDJNOUMtvEiD2Inyj26ulkIy+MJ9mmd
tm/kh7snFzUdB8YMWYiUnAmzQ9GawjnwNRRaJv/YTVarzhaTBfE1PO+sPPUnRBpY
ozT1AIUyvCUU+2PRo9iz6wjBBEFEukBBna4LaaOsbvlgBJApvC/FAqPvShxDjeWL
2Y82NhKD264lcElK5szGi7VUIoGSALA7waRUi1VZ/H7I0Bkd8ZzE8OOPplqsU/Xa
gSDKeE+aCvZxCeW9zj5nDIgZa5OBtlRfD9YABUlQMIq+12a7NBE9tYWZ+uQyT8Kl
D4me/OKYKq57A7FyZ9vmiWeCy+Jofy+Z7uCEqPNNwcuOa55SFx6N+vn0IROc1gSH
2urQJXyfW89K4cdR3ZWDGR3Uide8jwbDsGQ+O130JTyKHI/mz7SrQ0xghus+yQBW
nJBPBvJ1j+hoDHrBWccf1VZDRlIZm5vdlVsoMVRZNk8HY4/yGAOelaFSdZc11RSc
ZMlu47Kz+UhD6Zg1zoye0WRMtA7LbbYKq2U/6GAjtb0AureQM/WQxbvhkvqH/a/C
/uqLvcUjkodplt7FczYPSO9U2r2+r4o4t+MFyVwVNPUvo4etL3FDojwdOMQqK35A
GU/qdPcn3/ixxxg+6XfP1VeiJJxklaGOBZGwHpuZQpLbj5Six6XbY4IvFVcYCmcX
dXirssHdDNaltQkb1qSkIbTC3XT8ib0y/8XJOYJ+U7YVSnW7HXjLA3XgEJ6Z8q4y
i9DioXwhZabb3eyrvbyddE0xjIRTCCc7bh6ugEqNZMTpdROTrwQfgft0N/QDs1oi
6QdYQO8SHfkhfC7hIHiCSC7XZZVMhoFxE+8LkdPh2qfheJxwwuxvWY3j9e+pFcbB
KEjk6x69DTxqnS5GgAX0j4KL68Xogdt4w7bOveoSS6yhYbL2wKftZyOeq96Efi4U
vc528De0JqIMDH6MJ6K5IAIuoBjPICQO9i8crSQNOukNFwxF65f61e2DyuKR9KZk
mXHjpLvgtIJUuuEKLGgi8Jk0vgz82Yy4bsrxPbhliK8m/0Q894L9cszH3JzEbMuz
0oejawY+NKYJDLdXiTLSTSG/Z7bziWqYhWU6q8YYpwB4E1gUAzCCnWZrNzBCEn89
55VBgjkCJcd6UCE8m2xVggW9xZMRsdFKa8sGLT0voSGY9HcJEZTcqdar32HCsOMm
nR3ppOiUo2fpqbG6HyXGpZCH96RxAhcIfp8jjC3I76h6Xv0IAdUvWTy9ByMkCbw/
F3GmFpygNxpA9rqhI/u7T35Hk4X36FrtYu2l2cBZAwyxFD+oFiWIhZ83g5KaIqBr
eQA4z1Im6QAu2QqUkEhw5AzphHHCeHCyj7B8xOD8vID5p+8o2likzPoFTwg6ptXe
ZMSCKq7Wv6PNKvH5f/5gtaEgcXKQDvi39bgOwr0w7vdTPyNsj3slz3fynnsQcG3J
WK9phsD22XbjpeqdUo2Q3aXJojLaSHDwXdPUK/voDpgrP84SoUL7jZDNJJqa2xUi
FfHOTQ2Hp0qrZ6Gc/PgarN3qAik3iGEYuNbd2RDIuufy7OXMfYIzs0GFONivc7SZ
MIBhoHd8N3IFK76sYyqMg1xagIzK8WnCqZm4nK8o0FwIjiRoagwS8mA3sVdB6OYP
WkEmDkSUVheIPAqJBUDymEmr93/a8PDRCTUGgYzUDpntk+0d1wl655q4qqfjfIs4
ScdfjVLJd0QLOHy4AhZ8wqK2NVVD/3smgu47Wf/y7nupKaJrm/93vG+/VARW1My6
qEkhJqnzJJGlOh0BFO93fsdLODF2Hpop0IKwmzkewmcGmhKrtsCSFj1nx1TIVjsz
ijWvIvtdwF4hZaAs8ABuncA9LM965VNYcW0wXlTloV+4mTRtinJx99VQ4bkObctg
NTSy8RtiV1W/nghxMkhcTEQilp6OThbEWrLSNYtnpx1YEp0r2ZKSQbJBRYatK+dm
srCCDI5M+LtuNjyO6Mif2q1iw6fUcBHi0zlH9B7gHhYW1giVWDDEZSGyopMEFCpk
q6TWUp6EWeuYIZavB5E4vYwhZogCh/r1ZvQRH52mIy1nRRwC6YGim1rQmWsY27Ii
7OVOLOSbGE1yOPx/7SJEHH0psQLoQDfF2nQ6/pwIQ4LmZ0CJHeWMs3PZsriNVsrc
SAj7dTUE2gkgMTd8LaeWbAO03kSsxlMqbuJqmwZPbpl2zamHtQbxqB7ExgyEKSXG
3QULttBPVrQnRCfEJUnpp+5SeTHu/YkV/ISdHFzCwXFRyM7y7nvQjTSrsnl4f8rQ
H1tMQIK+wvgwLrcyQsO3c+kweE9ZJXKtP+MaJTeBJXXxvhQ+gqM5iJfVtkjfhNWa
M0JZUxEEX7/q/kN6sSgrSetNjvTYYv5mMvtl0l+i0LVmKYCte4I3opPsgSpyOQ7i
J/wPu2Fv0STebyUUkmCSFKEYbZJ4TbUkr405Q5iU457BkZxib9IHppcp7kyf54ov
8mW/p2f8nLpdpEAhIuaE/Z3ap1LpXWNKw9fHQH6PgJGZCo+Ywe3+/HZi8hygq+gm
18wRS0bz80Yurj6tRTRnyIXF0gWnhkZoFtAVqNdvM92lkJHB5Rd5Nh+GlUpZd0QN
qrDoufrSY9Ohp0li+mstZYOcgb5h/93qamyilEjzsCtgfjOKORDyAb7dbRk2wqYx
ZQMSpuN/MdIHoWoHi949hMtpOUVN8S2FHtFmcR/R6NLmp1Va9ALf2dJyQC0mtqQJ
6uosM0vnNR9oa+0fdIWhK7BhavIv0IsfyFi9WgvGmq4zZm2Cmqk9k2vjEU5A3X2K
hBeu9mBcz7cCczs1AFxH2OI2d1zlq93vM6Bmr3AuY7OBU/J1KARuSPKRV8cFkdoA
Va1qt0F17v0UCwlHpdfycGYo7o9cLeUpVMsGfsop9Mk/kIwx1Mg08y8VyaBww06A
2vbziFHM/X4hGLXGcHFI/rATgWFc6cVzn5ZBE1goPZM96FbUmsYq3d9s9WIVr6Ea
v5EsM4He91Psq9s+XTPBzx60RPs7KiZCcaMp7DCH0qWP90WigI0AspN30aTzrztC
d8ZCihpcSo0kAjzFJ0Y/MOIWvPDefWEMR1g68VN4JqBHVVy0BooL9LkwInIi9X9A
MHyUsFIieQN7ckKDs31o9xL1wSM24hkUNja+GxK8Kr9f1qDy6mtuXaJzCDsdOEK7
aDDSaOrupR0QzHeUEaM07ZS0a5jFnehwooRebBm2NpiNCc7peOaelhsA2uZ5DDX9
G8ZKdcXZrADVnSpCWc0zg7qWcsD0VAcli18lwvX0PvnkMcJKj5MLDfUoBUfAlsZb
fqjhHNFkT6jsGnoBK/ns9ymENZYUWVgneCJWhLl326yQaLtC8LiBhk7VfJ4d2RCD
8Qc5Cg2GkficV6b8TcvDuqz4+U0hXMR04es3LxnIepIVKa8jpnfNJJFoCAmMpPk9
tVeCazvYGa0PDOqkb3ZNUYM3oGxUZDYnqNCmTskI02+/HnGMNNVdOp2jrz1ORnAG
ccabKwGdhHnnficAAZc0cwqgUBWohZ70ZQyXGP5/2pnH2qFl3+yf2xAb4JnKFJW7
L2BXce1qU5jbbzLsHWO+ueG8LJXoOO5gbYFzt/fp3nar7sW+qSbhWiCQbVu1wVhR
z4Zzm3NwrAbh86TW8qakpKsLP5hRyZrkP5Wmx6ovAfaZcoo1ZU2xmDa6bhWQe+uV
5Rdx7s7MVSkWoqR9gkYeqiAo5D390LxpvvO6L1koh5Mz0adhYTrvK0/GYEGrU4iZ
vw1hTNWLnT4MaC5uxtJuwwCe5H3WzPRL9qBpcBXmKyo1efat7KlpW94vchKA3fNl
EY6fCbjaYwv8ho628lNuMfM1JTilvgORGS+jkZ4FnHZZGyfikdgem5ugDKZFR+k/
6TW2JZA42ycQ74so+8mE9Qv7Ax46txSKJ0idlx/Y4hGj+IanuI6drFSRJ0Twh2qw
CF7mLvzdrHOVXXHNceUDIKKTX1aCvkIFcRQeYNRUhaNurF0rL5RS412Bdia7qxrX
cvUpDkAI2lV9GaWyaDQ/rQy59vn6RwEBeKK31ycYJYYReG18OO8vbx1P8zN+KwQ6
Ywe/WvR9BWm+pEMK8vii1dLRH8wbnGdWe6oUFaf4WzyaCjClHJ4qzoM6vTt6/4BW
9P25y5238Uy5ThLYJfBo83nT2LwIMPMqgoo5k3lk8aNLRSTkOnsEWD9fktSAeTTw
uCDjzsLzjkUHtPK8lth/Ux4mo0MkEMOvRTPvNDbiKgz91FKhYmIZnPtD0ZwYNJel
LWpScdUiFfi2MklTrnL2k91tj5Hs5t0yq1904UMwT0C4zJlKv0r5lNAnvWGBPqyr
itNqbsnC3S+6If4ChGpyvTo3+QGWaF5jBQ/j0LTkHkLzSWtR6zu8aRBhjZ9zT1EA
Fnv/djA3QP51wRfnbIlPniT5TXVgrRec764jkMAa6DycroRmCgcgPRZCAYruSdId
kCo8GReTCcuzDiPoeWnq2bcl3cdeHNI6LsvdzZ6ijy+qCbnyq8/bE6dFhN+GyYJu
HvzJ9hzwH+gj+DYbqiw+mUAY/WeVOLwomOoShguRWmDzg+oYFX8E/nUmNNl4UabB
+qxxBLMgc61p6EsGKQdyhxvG5wwNG01eDJ4jBV3zhhqvr7JAXpSYE/r7lB2GMrrB
v82W/noU6BSxztrYDbbrHJ0vTPV8SsFNvP35gkl9dPg0doZdVO53zH4bo9qnm8Vz
NPTdkhvC3nE9rRS4SonZJjO0RMPoPcoTkh8EDcBo8Ga6FdQjfWirsWXC11JuLuWi
XXxVLwLWtFfnlyZ2vQAXQvhvk6iSdPnbOjUiO0n0VsOewljme3F8eziGhgVMAcds
0svZafsQf5R4qwVoFhpGGrBmjI9OsTxyaGCVTAM76beRfKXO6MbjgljbqHSsTCuC
Ic23xhmILPN11e8uUAXng43izjSNTPzw0NHIEurbpNVhq3SNGWtpUBpReBgRe5Ic
8tGOknTxMyzBHw4O3D1sv0jI9RK7sAfLR5F/ECU9JdHVpzbAJhgZT9Slv5rcRdm6
0JmJRxUcog3R1hWQrVPpwZbsxCJ/gTqe/c/ZV47WifV0UCkYeznfzYMcWRBOhHxN
cntdR3j4xPXasEHSHS//3vFP1Sf0KblUFp2wbCK8Ac7+4wZ5qjk0anotnIuAgtgh
e1L4fPXck9FR8i+sRSRKYvv84v+VOuCIyZc5nGcFHsOf8/PAdVQIephS9saihan6
joNxR6XvDh9Bi/O3hLdus0J3yR55SdljGfqXw3btMOl5O57vGUuzAfiqDg3VBwY9
LEnrgyaBhHRtedfbhdp08jNgxnlpmoEPu43X6szcri+RgZWsddArIi85J7rwIjEr
Ya0pjRn0o5y8xGKmBQWYDu5dHkwLmVr7ie/6UjB/Epcg6XL4t1LW+YC07gzQKKGx
jVTW/qYVfakP4AyYMSNVknrn43ZtQYANXnbZlsuZLCkaiR6PSXBqevva/h811Brm
HAZ9xK61Hh9Z1/1kmO/4bLIfAbfT/dhGYYnKJ0/yFpP+5TFuk5RGsguNcMYIWA+P
xadXKYlp67ZCPjSMA+pYelLOJLr3X+0Y48p1wPAyws4QRLS5RqprtiHs4FeBYGJ+
gms61/2REpeYswPYmiknokg3TLK1odCcxm5XNblL4WSqKFrzK7mupy0K0JLCmwlM
qhRci7vM+F/B6JoGdJ5JZwKwhuGkeN/3nAr77kNVAdGZhim65Y6jWaL/DPtYAi/u
RLJtO5ZN+HW5zSNoXVW4nSDS/dl+Fa1TI/HGDwZE9KhPcW6pCuVkliRjsWYtm2I3
Z4iZ3oK4qY8lESLEisbQVlvemV52fO7bfn8GMGz0pmnoBWUv1HspA4MNOELzBIHq
tB8rle3mEAERqi5G+Z6J+rDYQAyLQ+xgKp+i5tAvEtHf/9N2RQ0wTNyW6/BAsFLF
HVrQ4+VvkdUM4DGgrZEPDOpknSrsBZZGcey4kO41sSd+6z8p6k5QaOBT8VqEXS4R
4l3WNEiBkA0OaiNYNO40BqQMSDVhhp61AjpkWqixnZhqivyeq+4oMbm/RQgoYj9O
Mrgn4Ot0tYnPdoGOZdKRaecE5aSoC96I1og/L2WV0+iWW+cPSbIV9GoidGKIB1F0
uZvyS6qs9y8jGNaefJPtz8R82Gb2/3ASqdSgI/O1NGNyrxtrALrYXF9Rhbvm2Ury
dKZsEb1/CIuglu+qzaTPr4nYu4ozxvimvxeCBoGSNdPkenDJH8oKhg5b85uVtkZK
sFG3ZUss6eY2fqB0/a4Rs4OxpDRi7YOkLdP3HAZMD0O82s6ZvIWCaZl7tzUB6K6b
77C/OGYCkjCWz3j/EYNkf5C0e/9ykB5xZp3dBnQ/HF+YUjm02sYXhnTSfTHJZZb3
0M8QC7mGnt8BPemrR2IqGr52Hy1x8qSW/nczU6oJJL1IsqmRaGwV1FSdBox2lRzH
lxrp1kvvqokesK7YiZn1pzDmGcj0WYpC72CgXhDLrtSn6zWfh+S4xej2sy0fmnlK
zQcUaYQy4p5vUCQQj3zIs1EUsB4kUNHQVrAvSCQCH5TT/bvYff+0YyD82UtGPp3R
fcvM6VBvIjxgKc53R5etMj2WwHfE+Lepb5qxNVlvNcZsg/xlTL13iaO4CCVGdF6w
04eQQltXxHXheL8gHCMMGeNn86J9O+tFppTnh0dVs2NuPbIVACtquvfHS+Vo2Efi
JRl6WnG977koTBg2TrTOC/7MW2QL9Fzh4uAsqw6zXM3vXtjHV7zcjueEOqgpIHDu
m4YCSO9fzS5sReDkCtIgJRPsdbCAy4kSpc/o5sM7jVcqWTkAsdKqsNk6Md6FDoAj
4hJHH0fKejm7Hejj9Fz6lNB30SRsOAmoP5wccOQo8sn1uvQV0A2AIcsjwkpphqyv
HgOGo37ThUaClCosTxiAheG3MPweOOtrK1RCIHs6SWin/IhodOX5vO1PAf1SYHuM
saPg2TiaoAPpUCdGHUD6CW7u3+SJ72ae7RatSUdTuQFUZOaBGy2MCeTy/1uEpaUZ
8joHmLAdxyQXozIhTOVmsdxlAl2yomUeOhnjXQewFRliwPxtlU+DWTAup+RvxY6Q
7sDO5A6O73EgzYAH1q9j+MZtiu46kOa2t4LpUvQNvhFlVRCAbfJJLVEYMdz+NQfS
KOe8YKSDYKNsQL37EQhEdl4xibB3fj9CruTKZsOeF1/cJDyKlP8HqexdOsZV/jFn
rT8PuqC0G473UMgRSs4QJxAhvpk8ncn08IilhtAxPapyVKEfJdzOjYLesPBAC/kQ
XC6EP34EHS9kV1rAKbig4fIVxIFruH84HwfUMyrYRerTEwGNMEUZrK33dcmd9SXa
/H1GPogQXeNh4r7b4gDHMzdoDGW25HILTO2Up544AyxLenU50vHwThoKeXJg/mNI
KCxtbU5qw2H2YuxTr41Egn/PRg2wbqvXn92OGgCHuFDelQGV/nXnGmF2Vln/moai
vVcfCgunhpAfRx9oyDU0nVI5khU4AMB8/eP0snpqVfaT3ttuzmklO2NQkWC6v3ZF
0WPlxlQjc4EH2Pb5B8wvuvk6QQWdLrQT9Vo1fqfPxmq5Z20fT5J3oPwumgjWGUIi
FpuXFGT2Q8NybG29VxC1avt2uFi0Y6F/jAwznB6D4ybzuXVe9EvBKoxQSP5cTjfd
N7eFqFgqpS2u1A4MJCdXFC3cgD3z6KeVi5jmlOM+rE4uq/D2ecA/TrCGPGE54LEZ
jrMcO5r7VZEfZbvOJ5UHaM5pdYN+oumqJeFmYxomzPT6ig3aqo/3LzekXMjjDl3C
xVoHmn/cJVT+mLgLn+c7DaC1V658Ph6HcoDETPAanOcnBFx/j9ZHzg1rflOTRUcW
dw2CIbFE81m7DCzT7tWN4RDa7MuyKzNE1WhyVUnnmDsoPhW/jGlz/yFT7e+YqH4n
5iKsxJ5Mv41P1O/9RjIP+zewWc2vQltdLq7XQ9PJEb4Gg+FQgYcZXCC1txoVL22x
gXgf1yjV+a5NJOl6UhqRTSzhFBNT4jMltZSX60Zh/BZX9VjwqkBimmBFHcnYuP60
Ee9TqBwlH0zWiIWZffwkKRc6vVAFCJn1DaiuN/ceqkEuUJeCDIS0qBbemUyVypaO
7nQigGAI0RQC8p3zjqgwezMdBjVYpAGE0KLEv7/YaasVeDboGiW/oklfpXRGjveG
pH4dWajUO+WrjOgtUBr5NhnFolcUsfdOtYItrnVfX1yK8lOwvWiU4NPpKeZ/gS/K
9xp3D4JRNkDQs1WEbIArOSx25Cx7uGf5hFOZC/c6/2C8H9RVBOimw/ruVGYhgWFY
xmGeAoRpIiSSRtxY0JH9LcIKFiDJLspbsJAX5hRBYOS4HJrsVxyw4FSFDttRUeML
w02A5Y9IdStMPaUoKSHWShraauRiUgS5I2QiPnwZdH/DCv6A2udlR985RNu/kyJr
q+IHMIhSwMKcJBFIFp/M0rnD+o48Kjk8hooaOVbBeBAVryWxdBA1NNkvi6TILp32
P6sI3IL69faSzhzdBPOcf9BY5CTcRYiX9rP2qKcd8RO0MoxRqRRuZNIeJbAsEg2G
iPr++vmRg2MY/H+cX/kfGzdyk6Ts/aZeM1HKBZ0r1H8RC7smMEnFbfBHuJGLdlcV
+13ZZq+1FpCsAkFvHeEPgWg+fFeQ+0uMTplHLYDmAA5eUxRXMVIxaWH73pZr5wUF
n7cc0Gu4X2lRqYKB1/+X2IkKAcTpwndEoOJdvXW8gLkOLAb4kqNAzOJLdLZaFYMw
m2ddCN5spZiwwqokm2xfquekxYIuu61RyUxAj45Nji9ccR+3Yi346dKmrFNQyo6c
laOoc7khK8/gLKNln5hDl24q7MlqUU3BW4KQyb+GDhayCVKjFvgdxyCkelRxVE+A
6ByMWuVMMWJeJ/gOWEf388wW5jMOWZ6zb9NjmYc4MAmh+yJAE8uF1RSdyqJhJ9IQ
yRD9zDDBK5E3IOMjdUJR8xW8n3dF3CUm5tIHRZQNUDmTBBCkyJxMxDYbj2mQRAUa
pdQpYMFOabbeVhAgIV9fk6EDZbdixrRvCtzyvQSQ1YuVXUqeEWwSVRRjBxbCWUPZ
fMpCW463HOfD1Fg/b+4FKyBI6MEFLFkDcGUpVUMlqpOmVLU6UzjrKkt7oxLmv1N6
xEV/tf8MeZK0sihGNyFWBShOLFggCeBTmLzArTJjFwFxD5uyr1Al57FFjjCQtyXB
mJTbkQkdgjLb+Knb3HkW1vi/ZUvRZHC2pf33XTrZ4d3XFJcG49dy5dzoD0hUj51M
7REZZjGHlubgaD5renROTapoEguvTOQub9AiwFcIYe2BRS89ukvRNT2pump/bLdj
lDTaPyQWhRBEm5sxPhfYqn1LyseRWoJXoQnc4Ij1Iv4sDGL6D8SrF6EBshLtc/Ax
gCoD2GqX5GY4vbA3a2yCRj9ELAgZg2I9tJcH2QnFbTmjXeNOyOU4g18B6WrMOkV+
VuXWFCZdcdZRaLyBATCyPgaBlUTJBJIklSPlra6mZVUZNIDm4JJjfJk6zy2+GRcA
nW90PZLFQQH7meAz/AfehHYrn1+hyBE7bQG51UAqrzhn7so420Dzr3soZRXWE36L
r5c3YVBFX6hNgrIaPYqARbHJhPeKdGtHez7+Gtly3K8UTnL+1LotonurKW7C5gtX
NRMqYpAyfMYdkCt3d5mQvoVwXFdKTB6HFHWd974Oqic2i6tPQWgH1CTRqTB+SdAt
UrEOiQsnpeBhjrU+usRoY1hMiHg6UlnAmHsk8m9w8+1DDVPRY4LK0qesZAa+cfuM
jakNPmJVa5AAf/DvN7gGim7wawZGMYWP/dgJqDKcPxpkVUJ/UE70cFvZukDBx9NY
RQ+3lSLhgRVvr0XlaEaYJ9sscT99obuV+0K2rK/K4qXhqdvNw7lFpps+HuRVjjOA
rDh1V3v8/N/lgqIG5WPqUmN5rquUtlvgxMwuziaYReAsvaC9W6qhJe0VvQcQQSzz
4xbrVco7Oj9xBMBAg88faDx1Rpt1w20LzQEla6c5zcSnFmz/7b1NYeILMXx+cUVF
2PxnEBHdW6ex/SnEIwVeKkOz7bNJ/IyLfrLmfgWkBI1RSWmmGMJou8VZdSn2q21l
P3/Cq91qk6IwbCPBxNYMPMrfdW2iWvB1fHfBZU1Zrd29rBecVBW7PBhZaYiur7Sk
ob6ITuPOZS0zXVAhHfosV07RvG6wkf8NDZaphbAbCLX+dRQ0fiVCy+b1eZ+RSFTK
EVAp/OWFludyETEQ4UeFEey+DNCpo1AwzdoC1g9c7jqi2nUHgo//UToVfvtxdlW1
j9AL51WpAzOfc2YLB4ZDNTPp4FQoWNBVBiHBkVQF5UJeBI2DC4K/FK+1qnn5MONz
Qjxl23qPx5za6+QRStpRxNVoyKHtXqGPOCLc0kYnBiw0X83L4YZVn7Qt0dtr9qdg
crd6WyY8lj3gTVeYbUj7mr16vDfsRlzhtBsb9lZCuYLRFwwju17+1NKAZMYbp5vq
ca9lFGOVxmImc31r8SAnQG762A3YYzlkVknLZl50GLjzgrD0A04+3gqg3h/cdg+F
s04/TtsKSkz2MibkBRzA4205fB3EOSIKrLPCsAsAZZt7vLvjZPZt3sY/xgLteLNg
SaULzIhsJDL1mk4Hlw+y4Xx3qSoAMW5Oh2lJcmdznbIFyEqcM+Pz7tNqVBveAEYd
wma2QEcKEzgin0dJT4IjS9VlDA6fK3kg3rvidzQ1csIEFZFLw/vI4V08VxFVtcZO
g9sM+ZpgGOEasjKiOFoaKWY7WCthHFfMD/g7tW/cISEmNI5Fl82r4p+r/eU5mb9R
jeuontu3l67i1yQfx2CQMsYcJCg8lL2bIz/Dz4hPCVQqmSs9zuMkAFQqD2nlEjfo
EG0dqk+afv1D9n7m3kMm3l+iBsB27OMRhZGYDWrkDYDkC0gJIbxfvxhQCWmm1cg4
DNhF7GgeAg8COaDuOv5OSFSwQZlA+pehSVMwe5fwDevRb4wugt1DEQq5HmFjloGV
1FO2XEpeqhl+ze+ASCwbemBVOsOWhbNIWsX7G8XMISO7sFL1+tqH+k/T5rjCy7R6
re9GlA0RBBMEydqeO6sE1IFxRWxTKtNRpvjSualK3MzM1Hr2A/VdrxT4uiCawu9d
X0u8oMI9OUwct4RdgcwiR5zjJ2mTVPlaa4fB5+LFRxA9g6BIlWhMREPfzTDEEogj
UM4Cm8kaKuqINiwFmgJ84mVFJc2LWwe+i8uecE7octG28sMWpYrpFaKOhDbKvErg
8bih07QRlUag/CrEyqrvZxDuYBMLrg65Aa0fclBGnnodQgJEy4P4VT8ZRNwkHKUY
q+qeIn5kCq8srxUNn1Cj/Vr6MBemCh+p/y4n5eCvQcjAUoHGeVHOvqiALrMBAnrg
xcU4aoZmvFeau0xCBC0shq09EI4Re/Uv2i8CD5wr2noGG9WQU5J5VCcZ1oM8ittN
7lhgA/ZsFFJDJPrUfQQukTWMX5SWaP7/DQS5iRXSUiLtxDKcYEoAFGgXMU1YkrEY
VobERPuIXfgMVR61CfSiau8By7OmUubFSazz0p0n8owxIedLvopIkaGlP8We49UP
/oHbmw9J6BUyuUG2JRVg7F12t5BWUCn0NEwJsDTK+NLejRvro38WPH8+l5tMPesc
CtZypbFA3FQ4BatLvXrrsAFZSbreFLp2l31GYow4J7YxUU7axPk7N3xtw5TNX1F+
n9Dw8aShW80hc137nlB7qkULUr17AJNLwBQgYOL7EobxlMHb7j105KiukdSJvYOf
jMI8S0FNztG4rY6lW4z+RN3BTRoijDdxpZhrcpVf+Vm3gQONlm/3nji+TsxHitA2
1xbqUdh1rIFCi1VauUDomgdmeBncmgUj3J1ZYDy0jTOgudEjKg0sY+o/P7+b0W1p
YQOkRHAyOB2UCGuMlZuUS1g6aBi2SG5aITExY+ApVOjM3xUbUA6dGyAkd6ZkwP68
1+SDxYZZ/Dhsz1DH2XQhVlrsoZYRUq1uGVFpAA6xamVvQI0kFpzwdbpc5P3KgmNO
DoMQF9jieqmG2F64b+YdY7bFtCzJMh1I7ja9I+XVe4j6dI55Cxkj60EJc2NWq5Sy
6vkMkmOqALeXvpPz5WfpjGLaH1rphXkIJ++opusGpHoYJ44K/JZhM9tZfWHqjJPi
C8qw+xE0ENOhMDDJiqf8F7CN86VBIQ3tDmYJjymyHsJGVyVC/MIhesMHCpCCJKqj
bemP2PmSUKZSmLTCoay86yNJBL/8EdAVBz4FlY+lAaLhONCJK4qBT634fbPDhQVl
gFi9Uu270UgLOJqqIURnN08K+CHWKMiwNc8KkuqV5vmJ+QmXZAYYxPfo31olzBqC
XhChJh395Uxn/iYPJXP+wyliC8cK6KQ/IHt5EbsTfwU+UL5ImqBSRzqY+dFn32MT
hMKbBx7RBHfNFaoDcCntN0TnlDxSLPeYRBbjVVxqmx7M0ieVv5CfudnuG2OJ8HmP
YMjvwrkzGtsIwV+dSLUJJTqwSNxiwus9NI/o6nBUknHQyHt4VsXB2SnbhJEcx4R+
JPMiq6T5Q53AJWar7E2WbNhmkXqa3ojKUjDsIoSmGtkigU1rwqUZZzjCmz/0srPK
yz4EvNAslRI8PTSpQdqmeJkxKvQ0RoX4/JIHFSubgjEsGHU9lSSBWHhk9H8WBRIs
Fh7zq+g+qo4J3xAVd9OGZCpfkWaPgkv/0NEo+azsQ8IjoiQPRRhjGXz3ODnrX7W1
igFfc2h/QV8dItnTINWx015N9ppKXQLu4Fthg3+H9Df/grdxvY8xJlgzk3boWSeC
grIq5xEI3H7h+4DZNYsy0438RdXVTtaQ46I2GKpytP9gkYJkrf4fNw0VjHyJGhWW
qqzo5wefKwomi9SEHrVo/7SuclQBpW/CYXqs+OhU0dmZOy8wqnzTO6FmGg/ZqNuh
SxJIVYxg93OCV0BxMOYAyjICBCMdk0LKwZP82Qm+E60Fy6CLfwNf+mT6w/L72CH/
zFb75vF4qRQDYDNlWc138XS6ObLO8j5+Mf44HXZjgX6xBtKQoTSxq36XpT2KVN6c
HHLL104HalktZuf22TifCdqjIAiNvfTjVUixD3F9xwFt3Q5MGPNxnWMJuX90eHQK
ZUXtjCWbjX5tVhhoQqr4eYdtqpI5muT9bIZQY1CM2T3bhbp1VzvdjJgSjvOTGkiU
jCWEIyWXa27g5MTDe+m6lW0QK9EVPzFROOyuZXqISI9ndK7w98kQ7BMsgvDpqwxm
nRAjPP4m4q2uMop2cx4DTGdeRaNrLe1ah4B+gnjKHNhvqMSYlK1zymBvb7Z+qN8a
LWizddq0fwebORUzLzm3t4D9Luac5BYlvq1e3jswPkIWgxhnWj9Y8mebBl4FTBf8
+3sv0XifJg89qgfIdVOXYhsLmr79fwAjTOJVMRZfPwlt1d+Yxs5LKmQEN2wTRac3
MLMBb6OooKxKy+cqM6NZA+xDlmBit1WpaKsvkKnhTAtXF1+GzOr6vdwPPSCQ14fi
X0T0w8xJtb9jM6UjXetcCgeJqrskNEVigcDxAOwg1NUOJsOSgfVrrxTA7rOMBUex
FRQF6rofquBtNLdkkji/Co6jSn21gQKxo+zbQOaXrk7Cr0nWPY6ZU7Lr984x8Xr2
A1DOqlM0gTqal4PLXqmSD+6Kiv7hAJyOL4OoHuY+JSWkg/uC70E92tG5LL9v7tKW
SuWyt5bqX3d79LtZeV3/EMQTbT/HwdY3lPas8nhwNRtdLMOVx4pN0wwJas0Anq3e
l9s5v95ctRc/1STFQFqCXhLb6PgtTiMxx3eVAWsrmyTVVSGhNOkN5RJXxV2ZgZkR
+jLb/kcZyZvQK9/QdiJJgs6Z9duuaUvPQmYNfETYsp5E09iuZwFjjMTVqMXAOh9j
HkP+0OuhyAjBUyjBjFmoueI8W4Xc+SrznTmyOkMWFDvk/hDXOe+WMIzPt787NElk
9ibq6L7M1yYj8oR2Ec+30KCb5b76VOB6Cc4/Ia3rvNbdEZ3BCwN9P7ZTDXYAiQHP
0dJLMa5nncsJUMBMPK7dNaZt4TGz0yy+c9kZhrUpleFk4BOrtoceaavKMvOun53f
tz2SUOTXyQrXEHCfeIPQkBpvLSo+jsnu7m62jkjQqI7hPdIO//SAYSLX+cHC+1SG
Cd+r3UgbZgiC7U1Rniqe9GsduBchJji9ncyzFhY4LW3jVRG1+7CEqlMJHOq9gp4g
qgxDuMTpHF4fZQiVftBSz5y2gBI8e+DlP4WUkrt/hkR0iOvpJ8mS9RxqmVWn1NfB
E7J04uPBuUdHImAGwh23Kz1uYoU4ffQvCjX0aJrhXEcwYmbLQZFYdhrl2E4+NmPN
kRYUoj2FzRV35158Ko2V/OxSMWErYv8ii8Bw66p+hKESI7OKz5+4eqULMGKMukJS
sb67t+aPQO9+dJWqtId5qMfQ97/ygH0PZTkE+vv91Kya/ofXBS2sO/6QmubenyNu
CTFORmBwLK8eGm1N9U7LDGfYgruf6FTqJtiaE4MH+uAm9axjlrqwNjhEctCWx20U
TnGZ2DnZD7T3aO2HAdbz/GOrxm4M8muNDzw87yPVNJOvVNopNcDnEFrWIMrxKrHb
IQ/law7KPJrcYofAxijj3QHWsh0iMhkuVvkzhQexazRjTxPCnx07YbF8oAnDbcOV
7i3QQBdjJAFgLJ0tC1iQZ4WJ+ig4sZ7cqCWrYguuwkk+80fhdu4PXPjTz2cbqSK8
n2TjKuFim+AJrX8RIW+vTRf8PzTCdGACpdYldB/dxX5WxTVvRCPXh2BeIjOaFDUW
SOuaXlwOnqVu6+PI06PDpNRVPILa7m15FGR/JaC72mxg3cRlj2xID5RrgvAlR6DW
rkh4h0oMrG6FdwC1nngGEolLT1PyAOngqcU4z2lH55K6v2coG4HwXEG8gaBY2Zg1
Njm0EYbyHDjk7qU0HvM45krkxyL+M7h401bfWBfw489mWQpWoJqaBeTKvmur1TiG
d0EanoFxdV3kNz1HT5qhcuvDr7XZDfG9TybtgYnlj430d5y2KOxZwrSHm4TxzHiu
17ymUxO2rXCOSFOJ9d8znQGW2FXDypk7TzMQzHUw6XLBXwRDa/PorqW+aSL2t5hf
IzaZiCRK42CBaz2+32Zz0SkZfP426IAEzQX0HYVX74VpezWGZgoyUnHPhgrhyAyD
4QNt07e2mjbgggkk3cN2lvTCnuDH4ngQIFqO+qQwoRGa2efUV5m6GShcuzeb20Cj
6PlXjsPCFN9fV+PeEO1ugPwD/nLuAIt+6+q/rr/JOxEz9v5y+9HSJgHn7RSdvaco
Pc5nr0Q4V8fiKPqlMVPNhMlVQE9FjUfWLZHyOvWW/ite31NZjLhDny420ODIQl1u
CW1MfpS0qvf9l+ulk8hxU+s0IChoJX3BnS09ahHstsIM91jgeubOhA99vUcAD3tu
dbRZof9GCOdhEaDjz9AkOU044pkE/lodI7FvFrl/18dXwXQZI7iHLA03+UsP6+6O
hXcH7rzano9oGzS//68ovgpbRl1yQ77u66zuuxG8RI5+Bdp+jTMXrmmswucgHunJ
H2G8aVFLeCcZyvKTviURNrssCnPonzOsdo8BGEHde9lMo83wgGL6OgtfyCbhQXGT
qMMpV8vMEqYzibU2BsJXxZBhTBQGWtuYtlX9o2a/eblc9KtjXQ9svE7FyLlu3eQe
c39RMfKEvGbT7EzRC5WiMist5+ciwbRBpUV87LlvLkColK6frE+ts+jmPY7k4E8f
5rqXY7L0JEHGtUbhbbCyOrIN+XofsFGrT3jUjd/uhrFtEfYkoaQWabzvreZNqKox
1I6XwCy9CXUPFOmO3SkT5SEzaa99sx8DvZMOmSt5FEWRBM66Mtu+zvbi32I3AZx6
d1+wEDYDeU8h6tEHH8CWvGXebA0/XSNUfuSRfYIZgpYWTNLNg3yv8W3PC7Y5fSvQ
t2PbkOWw8Coh9Ao77pXLRH7xJTPXdQO8Zc6c9tJ72fkTHD5xRD/f7YytlphThoC3
f4fzfWIp6HzCuOLYY/KZ1GR4rQPqRTq8OkZS/ECI409acQFW5DYlM/SIwlKfkern
/3ySHcLU0rA/aJ5aKeVkOOZF9Ca/IGyIwCj7v3HROordcYU1axTXN/w1h/HMKjZF
t3mgFrc/7tLDqta+Kvj1PTJiFTjbSftMzeXPLVSbsPJRbSa4M0ggMey025ipTP5s
ET0DvkVCfBG35vPoKCgMziO025QQ1yXCN1ZwdRrGma0mVPHRdz/AGcoxZHko/AWy
r/8lKsyv1sbloyp/BVPPnl/eUBSBM2rH7TlyFCaJPKcqlICh730hPYxirkzbqnxy
ABUWrBiFhQWAPscktXBNuf0njCr/41ZvOI7PuscmzB48o4VXKJ+KQ9uzP9SvTiqS
UbeW+pSSPCHNDRRYZg4IvPuEeXuDheAOiv2hS7khLwlG2rTFWDA+7UADOe1IrSUx
K8r18uAl0rsBqghkCk9wkNfD2Y4LCyftXBoap1WZf9xeyRVcmoh7hkB/RGCN1h2Q
0+rleLW16chhnMsuNPKgkvGRS6KqDAXfsMQdbSZKAlCgFK8VKxp4n2AYg7UY79Fn
VtFTf+SYR79Y7mOiPbLrhuaMml5Zw/Ju9Z7VUvDMPt5afYWxakDgNXfDMg9zTcQU
4X10BESQxD3M9hhMykWUVJ0ZdRC5LkFRG52b9kh6Q7+TceFvt1oOVdRRKCp63Tle
Nw4q1/B4bMzfHxIqa2gqlywIek/uOweTyjusVARjcadJjy7IHGn9Mmb1rFsSqxiY
IjmKzOhnpN60ojwoF1+37r61BlVZWox16eP5Q+5Gn0C2SB8W7ATRseUqulfLYPwd
kqDNgCjnGWcR6Uk9tck3t3KVqG0IxkyxhO2BgNhqLgSJC0+SPHfgVw6IeUhT8DVd
mfzIwGOhg+ukQ2+fQbRBSR5lvAXADj7R3N1VLV+H2J9Cw+CkqejvfFVcU/L+ibm4
UjxfTduvPADJ2c8NlQsuJ3EHhSHoLq5H9svvR7nqKqrDFBXnDu0JgMknc97BFbYw
syfEFGjqDnMsMwdOjZq7tiyDcn+h26hRn6UG1fZJ85E0+7O0gvISnwhsWq03pgcM
v+gIHQsnfXZZ01eBlt8SPUQF/4diWFTC2HaZa23h53L/ZUKHtJLths6YsZr3L01Z
wDdTl3mNPanj0V0hy1lKSRCHcBsOGgS6cOnf9IjWlOz5g036hIGHmRrISxdI4y82
leoUSKObZbl15lNFA+wpUGkD96wc4iFO0xDVM5Y3sVTHcmD/MN9xZr85zV1ndBL1
EwkczfMIel9RCr4yL0pd7p/JSr8UYqbPwT3GAhF6/Mkatj0LWYGZ9ZOg48aDSBwR
lB5hv+QWUVzxh5uVXjqypSyqcCrdqP8i+O4zJNEfRapSPp+AufdusGFWricRoTmp
ApkPR4vnb6ylIbQPZelVkOY7qi8PxjcTlpIINqk8BhdnINEvV3dfp6E4l3IIj5ro
Qz15HKpCa6fZRybMCRJUMrOQqH14YSOhR6qBZUFlB+k4w35a/RFGqsjtD2f8OVxJ
Xl8NsZdTo4gE4xpTL8ibtBDssFeafbWeR7firkwHZbMBg/JsWoD6Yc8WMpLpIjsP
llj0r2xRhnZphESeYbwhug2zugtDHrjCS4QhZ2TMOpXcbtSwyVK+LE8INzDNaJS7
2TAkdqThdhXbQh3Bl427c9/l6nhdZw8o6WZj+6eh8BaElf6jkGhu6K6wQx0T/pkE
IW5HaLSZ4oX89mTB68kHdiZjXZyqso1NW2Fv/aIoTBLTh0fuJuVdtmTmNQuEfTTf
1ZTwMjKHIJI2WzKX0ES0n7Bq5Zx2tWpDAWAKz5vYwcPqWaxvIQVt32rWimbMi1gs
ARvFUx+wqJRrxvtKr3nOQ5yZLaq0ld5QqKYr0UOIHTIU5x/pKk2uEXaH56VqTwJT
Pq5OCKvNR112ttYzbtOdC6fi2afimpZSGsuriTHeIkwnxKi89Plnx8SxLWlDGfrn
+2gIls3N0QspCCSd4nQeFnExAD9h655XXEqm3r+WCcSH5HbF9LhxFOsfWsRV82e8
+s3nVt7w6096X4B60gr+CY1XQel8A9uI8210PP7UReH61HL/MlOJUTDGvx/TLHZu
qm4UgfDgQgxO9c4CP+js1c3gMmKq0AaFvvourEzDp6ZSvF/1pbNMtIYs4Ydo29Sq
iuUo/BsimzcFnXdihC2Et7k97I5n5atcuG3Czj4nUzuHkWBFidEnr4rB7ul2z0mM
OFsyWOrwQDJsMz80xMmo8N59/TuLRAIOYSpY6lfOQJfLveuDCn76+qFPX/R+l2Cb
Sb0/ps4MPNguzk34cLFj+K1jRTjVNWAy1WIiSQCmxFz44pgG0oBDZ+07vqUBtkoC
eqYrQWaUZbVAgNaFHNBD4ZQLs7BCMiIsUn9SX+t+xxSe0CZDS7T3UvCCaYsGYv5m
jPfYBjIceQsGRWpjfUKdAxd1eMkpHue0Z8isOQSpUg7DJW+dCZH1z3G9IN1KmDkT
hEG2SQMmBeMRhI/T7yIHTExyR3XiVPDlPAAYmNgSi2roJet/h5VaTmOXB79KJ8uy
p5eKlXByNXAnq6kBDve+mqrBe5v/b7tIFtGLovK5LbXfDtMXzW6UmhZymlbRRmHT
IyEgYP1IDMWQifGtM/19xATFZVRw6ZJ9ngCMPnu+Nfnrid5MD1qs/lKuWOfIgWiB
HgUSRA9otaNGR9koAdoIQ/rxHNDZLRQDFx1UP9GNozhvz+MdZhhpD1/fCaQ6D/Cu
JTdM/AmqqOXUmbff2+BT3jWXX4GzI6XS8n73rh/uq4bh3NEQ330JC5g1bIca9So3
J+QAmRg/MNk16n2Aapr+v0gH0PtYwVs8+d0OJb6TE9ipyMn67XgehDxs9rjLG9Hn
qyH1JZHdloeyMUWT9AdAl3QHSA6dL5mdNbkSXpsFZdZEmG3myYCItzFw0eS75OyW
7ZuV91FykrI3yas5/0Ef93EDO60RhKnYrY+9ARdmAMjJbfAPPh7cn2q9QwbL5kah
NQF/nycjQ6WXagfZf/daJJ5SlzNHfOJemyf0EVXcgHcFiQOIgL2gcR5/7TWSiVi6
kK2399aUnN8umNfHXiyes+Tmdj99QQDDd444TBY9Ln+UFdKmLqcTIgES5tYJ2jby
DBfkGatYx1ypn+rLqYVmiRkf/HBkk7GEuydBrtT6AXM+v9aTeuMKAeDi7kpdC1Np
h7m6Z0e0R645teKT8xOCUxcQt5Dnh8TOFYCngtnSPzjXQkxD1/z59TGNZX9a8SSp
e8HEzJlqcug/ZhuEkx2vLwZXX/hUSh2I9vQAefjCIBdaDb6vH1+IXnZjSkU5xLwh
mHn/tP5OMyp4ZA39hw5TjOukdNCY+ij6dRB1anPWx/Kyg2inWg+M5GD3i1WHqpHQ
cTFojhEJbV3vcB+eUDL3VauxAdH8OPWDdNyJvWuEPpQET8zcpF7L8VeMZkpjWdF4
7Wv+kYnSd9JCtPHyqPAr8sLQm8hzRsgoO05BhEAPXisvmM7H7CVwVtPRSd4VcAgk
cV4ZvKj7ORjYgXXZBTr/jPhwt+4z4cEqhwGNZx2BRt50AROfbda/gHj4YrZyF6rs
N26zqxA3FjvIXUMEsk9Yh8/4d87DNijuK7k/zHNHqsxAH/i3FJwc01xz1QebCZFu
foFUc3+hJCa/b0FCaR29MSWRnAe5BD4IqTXXNPkE33yMWlBeUaSUg4oWLVrDD31o
CMl2Z58rB/o9WoBNf7WBfAyFM5xptWeXvKhOrL/+hFMZXUFeXH687G6La+gnRzE0
nSwXCBPnIwt63Q1AC9v3UUs+qr2zr6kAFDNYzfsgIDlOXZEsJX19ba7aTGothXtf
xhqMrzbwx/7kxFk6CHnI1nitJ36SBfctqvhSnp+sVgvp3pllkzcEHIjM4p6YM77h
kHfjiVduXMZS5lzZCbrL/yeDIV+LpcRrIJAo1SoDth4oFNKNLL4r3Osd2qee3wa0
X+Zj2jiH8vixXup6oNNXNTWHoyG9nPbTHrAXmtP1sdVjixjmpXtJOMUix9iUm0JR
ITnXykdBQHfb8xtWGWWnwGlIYxfuQCUtokw2UHj0HTBMlA4/3vWzOv5rz2QN57R9
rtLlOQdp7V/iYIXASvSuPV4DaMjohJq92ZWKG97Xlzaau6VhRXPKgXgKD8GxpT/l
wmDVidlbIQhOcnwNwFE4z9oN2/Sw+MlhokWsSlcBwQqRyheLU+mhr1e9U1Z4IYO0
IDkHSCtTwbfwuSP/g1gj0VH7/+BQMNhZBd0izVFIN0xDGZT60Jv/D9bjuuVrxnEk
7Kc+E0BCZBsKVzd58muPxbOIW6EfnO8OiHlrciSnILfY615GZhWJn+dZW4dv4lKQ
ze2Gt89gEQ7bplCnCoAvxCfx+VrjlekjgvRAyKhas0P3HSatuy9uk3ESjvabXhm+
46FQHExrCcxxvwNSU0Am/LZejnD2BLBCyuTtIuBSY6WEHdeqln/rSQHNAXVBhYt4
Dc7VNCJaWaT2MLzaFVql6Gv75nP6AUmrB9l+9VwjU1hP4mHsv6cDnSxZ0/ocWg6J
xyvC3p5ssa/7hf7hfBBrBuc7zhLJndVJqy+YalhAdGpcLw69K4WBYREf30v8tuFY
5n0jxK12/tAqcMaYmBKDrkUs7SIgpCQom71iYOPZO+oRe3xlTZ4UfcF2az1DIaZw
hT5B1wkWRIv+tL4Pci0kvH0u9kbkcrrmVj75/j4+uKT8rAk5I1OJCs4isT+IrD0o
UxgSlE9QaHMqW2JoUjSPURJ8vGTV9PdFYSPcs1PBWunR1+w0v11oZ8eBsDD3GBCO
1q/xJnLfovYf6cjMbGPtYmyNRYZFw9qsX1+IVTEezEUjdu4OtbohR7TINWeBTEtN
uwGGrE6bCKjynJmz6112Nb7oYwlPYfpYhf9MHgbl4f8/Mb9aM3nYXBmz47uMg4UY
Awk84Dhp2uNMhB8DMlw5ctAOhiH+uVbhXxsgjgYPno4Yx3VpswaGUGjPPEpDjBY8
XkqrGY0HbwVcM/ssbyxhh3v8wrEreCDtJ18Jw9e/e28N5fyPRskzXEshZVmHBTAr
du3y7Y13Pt/b+s5RFeSGu9WoCOenswc8Mg7SJMD67BvTvn7DvinpckklySnt19Bv
DjoJajMCHRdH/b2+76FqxHO2/tiUygS4kP3X3mgBEpDZPFBj8xDKFSmzdhmdh0RS
FqGg4fcDKyuvhSHDfMTJzwCLt2nskWbDi3GoF8jRcHj8YVJlAlcW12+lgWQ5qIKl
L+51QIphXCOxFRbvxhRbLjE5kCHBpwl6WlWL7pbIRGOx9phcdj2e/Udjv4cWcpgI
27WQ50SESt22UYWWg9cdiyvaagkDhNYQA91SSSct1q1BsCK++xjZI+8XT2/10LYJ
5J1Yj442c9CYlXrVqE2+F7fHMisp1FHknJKSzhBto/AUaHqpXSa5kT0Jk9DUezuQ
Ans1f3fd8L7ru/NoQ5N8UEglGEXvSZU3Dx1bGVkcD3F2InTDPh7PnQOfagqiWVjG
niIBOXvIlqkiLHwDil29iubpbD9GGKxnHQVVlaL7BiyiGGFNrkfhkdlrb4tdojok
ZyRqaHBJhXByxFa1hD4OjCzpvbKlLVm9ya01gr+Ibrqc3AmmF8xNXiZrLiLqgV+C
mG4u5BTK8AQ4gSoaTJJDWNAcnohfLQHaKTxg0hhZohxYJbaXl454nUv3ZwfNGyoP
Wv3c1PnIv/mkDYZAH+pnIKf8ksADloCbjFs60l0EKqMg4HEvmt8HpBr7oHuR+k/8
gOOgWp6119RLD62oZ+iipCktV2IHNS327CjkLAtPmBGUA3Du7fI+ouK83XwqwlWp
wG4+8WYSSkZwSByb9PPSUsqdM6tmgc6c0lH/QhVWir6fwqPuhsBCbUHdLZv7y1mB
qMg2/ia7rND4a4F0GhDzk6hW/5FviPVIgHzJiX8/G9/z/xCRUqgcuRPsSW6OQBA0
6qsBKZDzClxApFl4ZVnGJHcEk4vR7ItqLsoCGELPmmxdAEo85OJqOoOa16j+unTJ
rG8T4Jtqhummq/aHvQ2qDW7yj0gqNwWq36JijQmuFffnzuWw/V/Y6S9NUc60mZHh
9xCINlqTv8APjxkJeqfNX9umtcFF5Kgwc9/eYGmqVAbdJOWYl/weMk7P9/ZroXdd
fvGxFA8m8m8lO4OJruY37rEPs5NeBv8KYTE5Jd/ntmy5UPS811UFiRArXgewE3LK
tfwXaV36f9UMWhVnNh1JDTE7fZUaAuyoPc0RQP514LTCY9SEM7DNadFIGuy5LawK
yOlXVOPWLlUcKpj8CXmCxm27uA0ZxUkdqrS1xVT6DOxqEL1h2g98aDQpXW6Uqx2k
6HN4qM5AOf7bbbE8i4smC9KibHD0seaMFFrpWvDKGUqOPC2Zm3yAzBjxM+Q7WzEo
PPFe5+0SsM4U4e0X3AUjwMnA2RKG1oYxNAwTENi4q8jkgY7KtNjQ4fKcD5TduvhU
1Lt6AhS0SNrNO5+06fXEJEmXzm0QTo1nYGe07XdyLGzHRPq2HwTp0oLLueC0/Ppf
LYYr3U2Ktw0YVHV8v/Hb6/SQNAkD85k8BhfzqQ26V5Wj+VT2CYKScC2s2vhZlGGY
tSOHyqWuF8WBA8quJj/3p0k1aSUZVFbvvDDTWEhLNapEuyQXTGUMgaHN2KpkWBxO
kwePcnUVcCXFBAzhw/Us0MCFJNvBopAPLJq8NBchMaU6uGLiYdWvzythLSqRe5tm
ExYbc7fKMUyooUD0D2H9aDX5xVG0bC2jAE1GIQZmyam0/k17YliDQ8k9I9Zx24jt
Y3vU5SuXr9FTgU77QlSUWkZUi0lGKLTSn6SucdN3+8j/KjhadQUIbZldYUKtqt54
koTJ2BEq9AURjW226uj7Ahx2gKhiXt2bi4TmuA+SRhDD8RRq1AFlOV3CSacmaqyL
SZzqGUxWbq3BNTbLN+v558rQlmRHJHt8qzSDg8i4OiW5xcK3iscbkon4XABkhXMH
so2wZykMS5YLpr7jxF62NrWkVPL8zdAS2XNLzBDFalLWDglFMKwxs+/ZHGkCjpTV
nhccihwNH/c8jKHZUOqlas/MQ9s50ry2Qk8Hn2TirtGk0Fwbmf6RAeXpgJ/CW7V4
Z+hYFkPD5/OJzfhUl1+vbjRVP/wL4X1zCVWiuxYkdKAAOY891Hw33qShcjJDH4nT
Q/By4ABonjI8DbcCiUdE39OCEfclp6Xs0aG8scNEHrfw18FN6qEoZIxjyMOnSMDB
AQyn1bOEKNygFfJ13V4HgNAl7BsDR2vw6l0Z5aw2a+Iw1EukWgcVI2ymZxx5fWS5
GsQlqJzGVnlyvR+njcQr4ipH+BAgwTJwlsCi4P2C+guDVshFUJN8C3XzYmo89J+7
UZc3XVclV2ypnnZ9bmu5VGxRyHZYAWUBjPKwJGbH0ZM3tYfjZPJMraFNksEohXpc
LCoyPvnAigEh9TF2g0xjGViJjJhZoMyCQ3w//hx59kZrjd3N7iHnKo6B2GSSGwdI
GHGuwwF+DTZDytWBgL63gk5i4X/DhwDnBg9T01KONeYPxiymRK7IPu+vAo99ojI/
pLLmG2VWxe6jKuFdMNhY6Yi1a+zQOm+V9ce+lI74vc4WtT+wwJRFkiEBY6xRBzRN
/STvarkHKS+5ox7i/8iErz06AXfDcLbTFMmCGBuTOaVvZ9ufnJJ//IK1eugyrVal
qjgLoTfNe6U+7c2fW0CnNRObP1bv7GQEUO7HxgIkXoTuW60hWKxHf44bc51kIzHw
NiZ/X5JYwrnSB8n1AkNJQQpGfuT7JwDGJLoh8rnN4wfz8fCeSg+UiMIlAtNBa08f
JWY+pJav7B8mmnT434KEGhoopwmZ4h4+svxvi3JikRprB+tFiIbYy5rL64A6bMnu
3TukRoH1wnFGp4Mzv5f+84JDvfdlKhd8SjZQPS7goZIyt8liqC9cUF8T1uvqHNuS
xgOMP48vyeKwLGHUP61fNbzHVSp9y+nwa8fkrqyhbc1BO7V7IuKSlUdA2HsEg6WL
zi9XyZ0XJQRc4JnPJJrddjoHgb+WNy+px9D6bq89kle0NTinEy6swmaQXpN04lSs
jG/kK7NG8rOaRrtc8YUbN7o581vdqIKs5cXCxpRHea27eUDV7VFF9/Az/WyLcClR
huzossHCuv8VjWKRrxuP/2Oa99Q/WZoivsGFp/avqE8L5tEQDBlhqoT3/9x7r4Mz
0ivwGWZSmCNG3nz5rVTHuwrHdLJ7Tctj6O2Yhxl57GHRZymhMfPqZ2flHonwGSv5
Qq4XkGvI+4GGZHML6/9Jv2js59vwdJOPP2OqPohV1WnCTJUJv1bAd0TpKlXTiNBl
Hn4d5rm64vbMGc+bt2mlcu4MF+eMbUUpihnilZwDPghqQSpC4x7nYE7UiomDRpUr
u7TCZILxKLQ/PG/3YHkG39stmxrIr8c+M0ZoW2mFUwE44qKnWDkrX5BlI/XJrqdo
OyyjTob5LUiXCQAW5T0ggsufrc8O5AMHKUONLdlwgywsL9ofPMfJgGFqLlnTUIA4
L5pzJ/NWLPtRaYV4cmlALCGPohZrOygXkr2qugy+e2TQ6AhhxeWY4FGIBow7qcHm
pCIP2ZEAqub72jTRXAdDfaqjWkW/SUI/2kqlfGwuyscPhdu6OwVc1+WzUPsdaIgO
YZydpcX8QBKzrLZ7f1EiVNAEMTbnucK/vcF4JLkfWovYfCWyTWNUxi9GV+sT/VrJ
pbj13n2wH6iWrbVH0U16TTXbYdgBkL2FO+jNWgkpZL/DGlgWhU0JqgSrD560dQjL
kpK6E2jT3RgDg4Ct0cLlU0FnKb18guHM5mfiWk4KGM9E9Z7yYTkIHnikAbJAZ69i
kVH4IGWO4FyiQALYiWyf6oknJA40khq6XBHZ466sdLu4U0quLuJYdW067af0HXfD
BZzFMZTywrXCWZ0YSSvlJ3mtFgAcA8f0Cx+qU8IXPWaFhIQG1Ohop5MmHj/5L6Lj
szljknM/lIWCupvZgqOhHKD9xFa0EJ2KG/LfyKjkOfkNWHdLzPQjo/d79sanCz5j
+i0BrB6dTre5RCCGIgMm2JDyKSruvJGYmNHNvWouOo9JAqNvchArPw4BFNQmxY+O
Bo7d7+2FKP5AfVDKdcIU037qm2FWp7zoVrnl14OnwTZFsqiUc/J77f0vkkhlfXgx
/KUtp9Qg9IZj/lDJrfEYG9dPhqhRMjhcFkG7mnBmVn/g+ea4wsjv2/IzJSSGyhLe
6BF8ArT/cLtFTZQHwnRTs5Kf7fYsqnfGvya7WVmWsy3e0jjoiOf4ZVbM4cC6TR9Z
sDWH+1LpXcsjjGs5na+b42shXM+wnXW7wkACB4l2QeuFdbNbMp4PkYTe5Uyyzft+
bKnACnecm15RbxGxRSp9LM4GnRT9uvRPYbILpS8B05Ie/6AR5Iohe/xK1L90IpBr
BxHbH+Ubp/FUni+pNsbUlvM1nmEkxtqZXBboa3UWgVdAcYTG6zFSYesaQHiJijF0
jTCFXoYOvjq3QNyLyK4ZpdsB8pgV3F5jUc0lnKeW/ozJO4Z7B1VmEU5VJYKsfW7G
jyzh57/Z5g+qtEIKQGsbBS/BJ2nBkPRklmtKdMz4H3VcMa7uA3J4/ViS7/egGARa
5LyNBjneC0E2S093DhZQk8zehIl7NwlSe7iHti5/1ejVHhtgCEkM1PEHURJesFK3
302a+I5o9Xeoer07N3Ud7aevrSuLHGe/g4SKuL9ee3ohZekOPPe7vV1iFsKbWeBf
ErkLKtz6U0dwlMimoepLyRjnEjAJZu4cBQshCrE3lpHcxBnpNH9Lv3p+rDCFM7Sk
XYlH5FQS6naYqrQy1ORzlkXzGx3PQHk+5dO0qz3XkJHyQKxqruRGxZp0vk97rrY+
LTUwKLoSySxBh8k/+aBVtgBFU907LwGPr5V7R6QzlJHe/rG/106idHnyBY4OoJmY
hwDTJA6dhSeMMuXxmKlvvr8SnaFKKVCmyhFbjhSv6jJNZq/umIyD0DpbPf9VaWzu
N/yklQED+pyinBBwD3652y/QehCUzbOmND/ToQZlTzYFYCNhEYKZbOuRcP8FaVep
IdX8NmVTtFmSKFCbxJ13nkvdLzKRa2HA9M/VA4gT4GVXgVS1xR/Nh6L1z/R2ma6v
wKInQp866ipdL79NMHMOsPSB9I3gTag7iGx7ZrY8iuwo1Dou4B3pVXr/a9CVbwU+
6k9y0Yqe//jSpm3M2C1edhzdqrwXacy9Qv6sz4/nQVjwxfHcrMHxSkO59hKlwJsf
pBgyezW9+Q08oRo+XAFcehGhzsf7JgJ/s2ryyx0tjDCN/US+gJs+8DifSW9e7yxG
6w5iEF/Ty/lYD+DgHAeZr/9prsnPHo9IGSrF8ONEU3ChjQ52pRVj1+pZiq1Fg+D4
G9FxwyECkQsxk7GLk0CTbIVYt4cbt+DIwr3O+hKg284GVqs61d4TaC1T2+3SQm+o
kMzvZm9GZB7eRMWck3VPvLcliUZ04xJ9VCFGcsncTJh7+OkLxSfokQDDmq/WH4vJ
cDWR3wCT7fS95LYWGCadT1jsnHCvADFODsI2oFZ3jbgD6MSAEZcdSdiGVlzePDfk
voMYz5qThJsRO4R63TvhrDY5Af9Oo37D5JbWabY1yw0ZK//wfskd2tyW1I7wJH31
nh5TvQ2qxtkiSd2nmS4yHzzlAGOlVHBPXDp394ue9cTcLMxWnQqvSZsLYrLIX18C
pUsmQlx4sNMEhqulGppi5ngXRkWiGXfG1F3vpgYyIqn0K5X3L8+k0H/FLAgIb/Qi
qA8X4MwJ0g3bfjTV2Lzxg6TeZT4PWB15AQNWZOrZmuSErr7iSJqbpZQ+urE51E+P
dnZYkOVSg3TUOweTYFYZRLWOrasEZanTB7dDxFjMUe13Pi2gFLRaLmVtvevYziXY
xth+DtRxycT7A4fXleWOGz4hAXEUkKT2ExdsrB7ymkk+hrQWhLa8f73DpITwdIgd
DSo8h+bi/ZDwnXXvMIT48aFwMOmH/itsz3v/fLpiQGEonWHkb3BzSYfIWbwgBMPa
OWzYarkpIFEXGi7/JRBGlO3+6JMvlEcVHfYllGhEzNtLsKNs/qAo78rHcvY3mbjj
Cjmrm21NjljtCb+soKG+a2NoYljfy2rOxDf9Ukccl2fq9KgJAZenvB7T07RwdP7T
PrdCtCeTczvnAtI2uZ7k3bFewEL7il3Y1czVnti/p8VgUSrlcZK9pzwdlG7u1aQA
tFgluexACXmnZKGEnngXAwGAe0U9lyMU0zatBPYTHTBnaOBFlH+YwrFioGReeerU
0PFkd2+JwFUWQhf78GqroyaVWoMDymygzvRDsBCCK9aXRY+W9o3GyosRlir9Hs6I
cn4CGgr5fEaUMprX9Ha2UFvma8/JK7va79HyzMCzSnXlF1o1jq+o4twEQtcHPuJM
9ubzpnZHvYLPHhg6ewt+DAP+g8j98X1h8tA34co8WkzkitFBvuBaSV8sZzyBSA0i
5edaAFygdGHPYgXRZef4t0k8rC2hMgg7jgtEPeXfJH4BUsMgZ70uH8CstzbsPjPA
m4fExcjLHRcBKPhdHRrLwNS7YPHTyeUoiOMg1OW8S6j0S3k9GA/OQN3SzU8SjGOD
TDsnQVN8wSPoVRPJzF4J/tkU+M51OqNRP/aYha1+2ElwwLwq5dzx8bMwSoLXZUI/
77SzT9LjvT4yBX2LS3UW+90qcCkPijGQs2w2Lgd4lk1wpdg/LPtSiTnZNLka83mm
Rc77byDn6cpp8kmwTAw0VQYSkOg6YAJgCCR+gPGmLy59WIDz9wpHSv1YZzswAzD3
w6q0vqyJy2m7ZerJRmPBYbiAnmawwAwp5Np3tzRZEkjXKTpIKYtSl5wIHZFjtfGx
PU/wgU5z0rS9+Iwbv5Pw/YZdYSKCkcPKF/g/Vgk2eRYRMxt3vFd0kXkeWHrF01yX
CwdedvIjSHySHIsNzwwlJ9VJZ9DZRtb3PqhI6gCTzR9luNr+lZdyTMea9Y4r7hL1
viIkgiolueSKaY5fJMBrPBWHTVGNgURfLI+0d6GBQe7Vgja57of24FkjClJGPuZq
kbl/h2GsUzY9AdJnDAJo62egGbpFIIE17kn4gCn7yi510liSaDt05JuRGUjegTO1
QM5TxVySo2qRjzQjodn6bo69SHk9TU6wdmtz5YhpwAGSpdwnGyeOpNqbh55STLMo
eQma3TzexaCZe/xEREx4FSg9rjVBavEk1de0sSHqW6bfoTNIqrvisF9yyo251Ybj
kYSZJbL0y9huEkibCG8nDAGlpvy0cP+0aWkFjxxDCJ2mVh2Gy2s6XRTkn19IrxEs
IhnUTgqxZxrlFPHGG1SttFKV/iIZuWigsCW3MhUtyXLV0W/vDar92VTmwj53H9vJ
3502XWFG2duhrsiyvf8Sdq68m9eLQFvlovwpJXcDItwjNlzhhxp3HsTBEXe0Sqgh
EXOFbrvEA2IMLuf0GG5SCjtgooQ1gyHBJ3YEfnn+kQ4IKbZF4jQhkQkamTeap31P
ECMxb1Ow8TjhavGq/EejwKgfIG8FI2pxpBdomCw9jW7MnRt7HqGcqwP+rW0BskgZ
PLYeA4nYcllZ2ZHV6EPeEPOe1XNJmhBHFoDv7Py3lon5JBU1soOxlPYgG2L3oDIh
L49aLyPG50IF4ozf93IGbgGhpmk3zN04NK4bV3nsb5LsOnB/XJl+mQDdywClg7wc
FM6r0KfYsK3fQoXlZ4QYXT5i0CcTOUmO4UYjtsTM6hVRr1W05JdxWNjBZlzNPPde
EQZR1VxuTtj5N+GvW/WzQ7C8YuivAiW0DyWTXPacwhGOnVvz8K+CcKJBDMDIq6wy
uHNPJtBUxuDaFZdgf4bsIK/1YuBt7DFVDtaWlYBVKpCE+HfpGxzxCPjXWD9fTmpu
lDtPekjSr/92byeQEvRg8rQi31K+hwbsls4syM8isrStH1vtb8tYhGBN7bZ2falo
MG1NB4GCfPfPAO2keX7EVr82MZe79UEvPSnQgACemoaNTJdp+kIn+bSv2gXB25p+
8pIQFoRwsLJu0pyXnGD0Uu9qrl+9T63VAXgj0ZVHwBXwyJQPH39TWCFb4O7dS+F8
4PIlGulHQmIk04jbctOpx/NaK5Urdehl+jB5aB9Y62x66a/pQCtDL4WrOh5l0pHN
30KTqmxyFYk9x6dinuJ6UZjKZ64RLUhATDHuGOMhESv+ImTIsfyqO7P6Mq8MyYPB
9VxipPj+R95HOE4ROS3yfWB2Ctev+gboAF+R+6AisfPQN7Hput8KhtgA533xnZzu
fKqxb5cH2ug/VVn9rK5iDJAxBxdwbUguvbQ+BxhrBuX71xdTUGLKz+PNASmyJaru
UIF/q+6AmWzyo9Eea/A6ANGf+UNVDzBlp40JEiQabwg6UbZb1+IEqddavpAfJ2n/
BIG8LvbeiNugRo4RVCoVsttuYlv2YGAvKP3dbZL2SU04IiDD428cu29f8TQ7oJVp
QPCfrL0T6EeQgtNbLMGSCxw4GLe9pzQk9sFuRUWEGTdIpPnQN6w44CdeklA5lliI
jcpY6cikkW0p2V276G8dS9L3nV6eeCfVvp4Z05ly78LKU66igfj/Ne62ISytvj5I
yEdiYaEiUs8IPEqG6Q8ZHsr2ITsS74lf2VXca2BpaJ7vHdNaYrpDdLi1hQgwQZ/g
eo3xZe2ZI8VmRxJLGHfES38LjHjMsELOPb9Nt6IS04Kn6NHzC4z5TgaLp1wPYnFR
iULJMHAiEyJPiPMTcTOwrQTMrYtuMIMGIm0MQOgPjwD6eti7GTu8FLanxEaz6Dhw
8+zUS272tP6PZ1U1+1udYBzUievnhS+5VTDyXXWyMu/OibGaAPw67gJtYgwROKVH
Q+RyniO/Wx9KJ9R1ddmuYVuBvOLWnK3MVvpxoCGgfk0J7CTnlzou6D9wPO9SlewW
Q0sZbcgrU0SaqqGpnjjGD1uvkP4MWghuYwGBqPpjZ5Q61VpGYB3CaiSVAcKXP/mo
NwiXiKpNT8nKd+wGLf2p9ly+CT6/6PnznCQjESKyRaw3rgRV9qWdm5HHlNb/4IXL
29H117dL2RsXWm0ynl5nd7g5oxKurjPlO0DnQchXGUZM/KVDBw1qDiogF2+n0qv0
SG6HJOVb1oSYHXuN5k73U+7adwvlry00o5oxcjbaDsWpELzY2lIgtInOIlUpWOV9
XIVSAq4r3XG4NkdBUN3E29foUgLxhyNTnFp/9l2HcGPi1LQ4vN9Il0QeXDhKJKKE
zqkq1tKjEPqVzqoLk92py9ihMmNxn+gj+ezmzx7kOHcf/wIwDwXI7OPQIbAisg6H
sxuliBiWU9JG19hl9TiytKEOqbq4b16T+O8eQyVrcZF/TR2KUC6DAkfyD/aAMbqZ
g9pkujVJ+qwHnevumeJP6ApQ6BnHLoFrweZih1Hv02bsT5+m8vqRZVFvUSLhT8z9
zcelirxQuxN4cdvwJKmUxJGqrxSHqNN3qCZ2odvSWLjA0FnXXUYLs1K7sjjSrwv4
iYQe1LMEtpZeR/5thsFg/MPlcziZEbAXviK11U9aGldHmu3nwVnnlQg0nEa4uTPG
PwtI9EF08vJPcycz9QMjsJrJS2iGKzO8+l4JWIJFcF4DQAg49vYVDOFouYsnwlNu
jtG55ydJQNOHbPIJyBgi44t8zdwUmEjPpaM3Xxm6VfuBfbc959gHK5EUBhUoZl1N
Nn5BWUX/VxXRFOu0SBSKUlUDhqLHoIc1vW99Hk3yG2PrHpBSqOloJU4WhU3S2qHV
D5yFwEkITlhAhfoMEVYzXUIIsoC+MwoEvtrHV/VYoixnbM/ZeHiB0kymbAZFurn7
0XgAlAwfrfoqspSiy179nditbnxMoa6gjjhDT/XfUZ+bpeFIwzRLgMeIQzZKbbJ/
YDlnT+6P1ruB9wChqrQtfDQ4BUvVKtnTjO7+mUIjqdW5VDK1XMSH9QBrvL/3GHBs
dU1gYD7E9Nlk5/vBv59UlcRMzWfhS1+vSa68ZJHedPi+T9ihnuSPSZUtsKhL0bJe
0fgiwIB3nLaGdfPOHkvI6DHlpVvkLt4StMSaHMNUwQF2PwtqEWGgnVPzEVWY2hjl
VXLkKoP9gIgcaMo/TbUcti6eu+DF7SVngD1fEP/q4Cc8mnqRtF0+rtrhkh6abcyU
ZVS3drE6BwQbJuVbjzZoRiam/POL9+jis/9VxmVHyiGV2t265ynzHpHtpqJhjtgG
+xyW/ygHjufgHKc+wqQHyxqlC1QzjwoyO1hzZ6kUBZG6tvGBhwc4N1ktcR6ArTm+
8B+8lnzwXJNqvHFl4BzOE3lGte0K20Fp+TmSKwHU65pNlpLMPy0JGgE37xRTYAil
bUp4XM9Ito/UKhVD0fHoB1/VHEVGaUpacTu+X5SK/KeTTbidt4jk7+16g47sH/a8
NBsONaWkwr0pf2jxopvMJ/MDB9GFU8YExajFq9b4NWOa6nRplx4VjkKcEkWdtTi0
wd58kh6GBiz0tSmXwUujeQLJ2byoQ7XMvlkhL1hKXmUyDe4Z+7UnAo8uF6CJ61ly
CL7SCfuSOsNgvSqBUnvOvGoHI8WgSDhkYLDWL+u+GwiQrcJ7s/cIdFdmiAbrXd7e
PBvSaVQND8Yaz8QI2zwuggCtR5Qrx6wkWf26iqRCRA/1K6wCfMDMbF6JUYAFD/l+
Wx18dRmnuGqOiK70k1PUifvRNilhxH34htycW3JSKkPBAmn2M/SEOFXyUdYSBqCF
d6m6f/hxwVIu87T4SwaRALGiGu8f5tX5zOsPRr/Gv0JatIY54Y9+KyWuJ58Vh4KX
y5L37wn7YltB9pR4pkKJUwwLWFIkyu37P08xLGoTKXRjL3QuZyNXYo2MaBP9PEPT
bmVVF9E9vNClcLreYU8+rwZc39CRNNZfqqPPAfhUV6tT+5jh5aDHagy9LNY7JSf7
06PMT3/s8gDLTj973grMAYo/Hr94THFvhcWXyNQFq2CwXebLodw+PvyKyy1now2+
AbzNiQjwhRMVcklcbOlANEtJ2iTAcRLwQo0URzWi80XpF7SuRPhOXNCE+xIqm9D0
n1xmkpZpbyDZDs4o5H5knEAKQo5dzpDjfpl7ln5Bp5VMz/zmros9Ezs1jQuibJl+
/kZoEvW9ICcJ/LIkb5Wv6B09JPI3uuOvBX/xvDsirW06uI0PAegK8G3A38FK1pBN
PU+C/zBOAWHA+Yb9I3Maof7rDlGSoA6bHLAf2ZhiGACzo6GJ5+Sb4+3lrYX5j2+T
cuZDEn3tOHs6BDmkrA8BOSgm3u6MKlglGZPkZxOmWAel6PG7lQqUigvv11AGqKwi
g5ocvbDacyNm9JrAFx/wCrLpPDgT2Njmn8H89155r4zJdH14szx6FJooGrlrXbTY
6GbN998hMXloUcqXvK4+s68WqTVsctCFQohFQK4dAgTA9yWnpcpUVAUNrSpDl9xF
nK2Zmrfy+HGBAtxuLokXWNdbCMiw0E+LG+oEG80MRQ5KDN/2EcBkAtJHoERX0FTa
QbRvUH6hkpq90zLIR6ioCqVzS+Kps757Aybsg7c2jyvDGUTW99a79V9jLbYkrLxe
uSop2oai6/++f3PHUVybod39wd9thTA6j0HlIFaNhzINKHHA7VvgVSOBZJG8H/m3
SEVBFbGzItNyLzq7IKdJin7hnunEbs0gfRuXB0LDuUaKKguzFV4upD2qw1f+joHI
A3YRRFMBr1xdBf1dNqepVWoS28ElQX3iD5N69OWJYkmit/WutenHWJzJrnRJ++iG
l4/QDHReGWc07srrTiPbEfcDYH3w6a/aLzNRdeU6RuF5mZm62TuiYow3KaErMWKw
iV/2Bh2+o7EMD61GWGTEcM6GeNfmFM3FA81fI7USczt4NjbME++R1dfHD/ArUI2K
nZG1F9w9iqKc7u17ZFql00SNCF2NtmFczWq4Fj7pLMthvYNYM+zVYPTXgq9sGbnv
37u7WdCICDG++qCzT4VH1PyuF0lcK70IsguQki7Hmx21BjQ8Brmj3+xYU0e95Jl+
C/iP6NKuJ4a/eJj5XMFYgkb0b9g5pMAwqje08oIx5vh6FXF4g9kiOLlGSIh9Bdwr
3A//D/KWT5848L7fdmudqrPBNYkHmDD3wFhehy/CAdUGdzaHmMQe3/+ydOIECcD9
4ezCTXIqNZdpoK/ipkOTivf75+/ZRZzX0uL/v31FClEMl4S4gCBiMlSgSEPuUw+C
pWZhWAZ4rgi3fr+kX5ZDYmYRe6pEPQFWu4QxiiLtWqiIrSn8ADtn1BvA0aENDhm2
OYoBvBP9Gu8XNdR+P8yS+FDUhlUa8IVeFFtMjr5JIGGzYPqRtLzq3/mK6IyxAJjR
HkDsizaMyjZ8HONptp1zUstXrl3L6lc9ukMgM1FR6+B1eYmZVuTLToM6NCrRtaBY
Ip54t7M7BlHhhTBObFiaoNef+7luklAnm2IIJ/jPjpoz5V7yzObz8FBMneuqIBqd
0Cmf5ilRGIeQ37M5KpqKWRGe+zPiRF1wNsdNvqiCpgjOh8vUYHECu97FwC68As6z
koSHGLI0DQjgaamKfm+HoesZAl54xxaYzIzjJBlT5xEMkAn5fmSAnDuF7gkvdMAb
fjuWsMUxg+ZSVKzgBj+3n3kEHKgQrgU90mq8J1CZ1Nver1G5+cnCodvnNFbWUTQj
hzNszkIdkmAOF81kr1Yh9ah7FllTWsFapGFrmvqPBeROz2sN1n6rYNB1kL2YKAeK
PMlr4SfzP+usMy0oqBKI2Ca392tCCRcP/Yjqe7rsxjkAFuUOXaumpI5CZCunjmhc
iDw0Hih6//KPBgbeJORrciPuPW17lOdocvgDuqcpD6GqNikI+xIh7farHdsi+xz4
xqq5ngth3mbJ3tq693AwfnIS5/3kVjDqF3xz3+U+fHsXdbXpVjtW4whusI6JFJDC
6APTkvCoLdmJRlND10p1yOr3NrzErmwha9d/eU78kjHAPXvA8qNfJzt6OWNH67RV
hsS3GU6nj6TVzjZb6FJ84gkdH4aShAzZRO64CRktly8pfWIeBIlWXUqQehZUCrYB
xkbIJfFk0MqHqh5B0yOI1Si7SNB75CQzZEwLkL18LWWUKsF27shwlUe2V+QW/kXO
U/fuj/xx/CAq4wI074GC7wcOzeIJzGOBeOYcdYl722bPr/W1dryyiPUiVuAU24Fp
UnWNVTdRJGezsnUKc7zGXf5ZjM8x3+rLRBYhNCpZkjhSdJyejItDkQiUFMktp+fG
8O+BtQelqDwZmVDYIZTRRw896xU4Se2rw+m8hI1tGikZhjSlO4STeytTQiAgx7nM
e9k7KYWaGOwxd95cBctAKhfhRtjiyBwoDevlu3gy4M10ndqTw9ACTs3RJK4IkoHz
lQn1SoK1DfW5iHzHi0UgPCW+dXlLdH35m9eG79xdx9/pcP13PnahKs0FTIDgUVtd
//Ju4QlPDu+ZTNm5kk+b/bZuEub1fkVjDKnRg7aI12lOdue02kt3bQKTxcr0r2+3
X4UE9oOr8TTH6BkVlXFl33H04uSs6wtF01Vyhx0HLCY5t96ACo5woFrf5RR0SyEG
6gCx8BVVzx0g48QrmQTkBXySAuz1qJH17RT0/5PjIp/LiXe9zN31TeWJXB3ZlCDg
YGTzL5CGgSfRtloOhDkM9Tbf028/b2sNM0fYn7f1NnCdKDkAkvTcEgymzdaleJyI
My0WKjCvklMgjVZF/niqu4FGmKJfgUhfMfvd5llz+eEjAtQouGPBZILODCgtx0vB
iNon+3iBrjPuQEerS15p6ZOSX+sq01f1udvPrNxD0as3WAtvqgw1BuyNEyxZe96D
VzCxsWIYwgQRxUPK1zcmbPTFbbgVadmimfomX/0WaBsEuWulHcsxK7pIP3lnbh5x
m2noaDzhjkMser46Er38K6gSgBZMorWWS01rbpHKcd6hkDdi/AGD1qWcBoOXl7Hk
JG76WG2Zo2hLbx8xxB60u4TOdw+KkMpkuesbyQgaP/1PaNqW7xzpbYYaqt3KG4pW
14YLWTHnX60AuVH14Bmm+FhEEPRuBICPCVJimc8DHL8bjGeqyS9cY4YGURqkSYRF
vD7csC/eQobQnwcMTt8C1yJgRrI0wU8gi0stWflxBDXFjdxLbJMCNOCPG2aGv7LX
FVcNQzaxydaclQSgRE8WcHYWRpkl55IZ1w8KDuZYsrXG/Dviae+O8qOIg4LgqUr5
tNxgwe5fUqOHgxMXv0PaHxqlyCRqBUeuRJzxDodlrVq8hts6K5Pa9OoaWaV0nhM4
Q4v9VXxfb4KF/QhFq2TvKZ3GokiKS7hsbUTYfcvxxA+oKOJxKIwxkooU0F3hT5Ui
AJrGjrqwiCvDRuksfFejz8F8wFq1l1sqqblotfuHoNVc7QWlqdfAPNTYFqvnO5oa
ilApKJfgZk1KpVRjW3bsAQCgjc3Kyohns5Ju6N356E7hXtLpwZ/mnyh8AnKIDOml
lbgbrwe0Em5+1cpFM/k3GBzzVS7UHfJsescX0duVaUnt7Hmp0AKvVydPPURxZh1Q
uqYgeqRseGe2bXfq4yqbA8J+fc+4i5lXyzdQJjxtzttdR8LQv4T2Imwig2DYiqC5
sZSyNqJJFYea8mvIafqmA+dRyJ4qmyp2A3u/0ffEy+eIlpekGNsJkLY1RwcjV46c
faJV0s/RQHwKZeFTYutM8ng4I1gFpXOo4R2WNmBoUcsQmyDN1pDq8eInkep4js2P
WmiU/TDEAqO/oZvh9EL6IxI5WlGZ+6KeiepZdWFMKgcsm5xemGoB1LmDkcIa33rt
1vQLvof6MSquGLGh3QQMEgHxHJhV4LzPy9VkW9yo2ZLAqrC27EADv9m+GZnVghMc
ophbLjn8i2YGrHoAqXSxjkcxhC+l3/jY5y1KjbXZ42jJRu/2g1HKSP3kIAg/jHbE
Hd/Vfo6AM1lGUh2nUARb41QFvfwf93dSlNI2IFSQOwZ7FD/LOnYFkNXUef8fzgRn
mFYOI4i1OqZIh8rUgIKSQc62HmKUVGtKd888ebKg9us9cij5J9Sf+CP9wA1CobcW
6j0kqJ09ks9q1iJEyLxqd84ZuQKvMD98hzXKjdDc9L4OAFWVMh02jjU8m7wE2Nxu
FY7PhdON58zGR3Rf1/Ln5uVIRQLtmDwKmRDL9df3hMwCZDSZ+rN26ry7INZajWfr
gb/6J0DQUebcEYlL/2PtLelOJ01l+5uQSXoQ/CUDTVev2BM6ZnihJkxXgBaOmCy9
uDiSnuUMfx1L/uiVmfllarBPAi5THkN16CqpenQiYW7mcgYF6K2rItm+xSLjSAn0
8etqMKsVh0G06Bdghaf6Fu6B93loQnkrXB4AZMQ4xtd2TG5AKK/6vPRoVz+TP0iQ
k8neEa+tB/887Z0XWOSgfZ/b9hKOmxfrNrMIlM9+nmvmSu2fz2tXXDNXAKxPpVRD
gPoDofur3fZINl5Ng1C0ZUTqIc5RZhJIUc70AnF8bYsWTqe+9gXbWh54xVFYv2qY
2lIeBaIhcwvZHhYNBRgSDnVFyDEQ06Xz2kfkaOBPmfzA5YkLjLQdlTnkBMpBTJzu
9JLpTr4rzweZge4oqQnijtQvEbxDJN4h7tZHrVYs9W5FUtsnNSQNQGmomjBk58Xp
1sSNqltW9wzILVguvWsRlExSidKucxqOiTkKBdp8a4ObYN3vROvhXjHjE6cdep65
yUeR6II0ToPwFM1TLgxX970T97oly36G+j1NtGSMcBor4wYO8be0GL1ZmhvoGwxt
KTa/LJwfM/I6pdKRyatZTB822fAFWE7jp4mx4mQOVpIsX4G/ZkbzI3gvx6b3QlG0
XspU5HQNYefD4jH6Z3BibRQff0nmx+5G5H5H2xzce8+/ljaafSeCWCrKVh9zYhZy
XdTJkbDX5qzA2C7nR+vVlovOJeLVnoM2i0QsRs+jcoAoqj1F0qsxhI/lMZfjHnRB
n9ozqj/JRM2uyBXhwLZ+/jStQM0a9+80AF8qTs7/gP4iP+oIi/gEak+WbVS1hKCD
hM1U0PNvKzlOznuQRIpUN8wou5Xts/Z8q/Hf2BE0YANI9noRKWssy0zypeDu5M9p
dwZqrq993RmZTbCdVIp77oWndUAb5jJCEnHvhM1eag3Z+NQAc8YAyNHBZ7DeEsrB
lc6r2Kb+AXDiOT7NEoxkkl5IGAKJAb+dw04OV9GOt8sCn5zyyC/xoCLKz+lMxveX
qeaLs6Ef0hazHqvv49Ce/U+sqhQ7tNU112qTsr/ClisPfq58gRg+Om0tNv0J8p+X
KzenJ/cEMSl3Bvc58jmJTDDIk/BqrW8qLwFoiLuYG//L4iFzWJCkuIDM5pyAHtFj
y0z3bqmu/uHat4TsSDggiW51UuN1Ep1fRX+pa0XiGtbpB7Xapsym3iErJEnsOAQk
uGw0AF5NuuJJXYmie5DRXt68W7eTw8Hgkk8b2xzfB/17hnD6+0sid2PXBh/kqhyy
djnSA76R51fH6KoqETOlBf25m2E0A2H5ANANiU4Mazq82j1Q1wL/kq4o+LjzeK12
QmylxgQ21flafUcWCPTuv4QiAZuLOVbT3kWjg/F4gviEfAgbQQjq9RbZc1An0x2M
OzWi2+i2JnHVkkv26DwL6c+95TVSQtj8fCHqgbbpXaFSDD/4jZvCB0rB2xJkvdvf
2jvaE4IlpEsXE2BsvpDXFWVqxRp3kmS5fIx0VCIapuboBGLk67f2GAE56ZdSyQ3i
Mv0GdkGXohjpDiEjOxeFMV3nGg0GK+uIudXI1RN8Y4GSs6nBET6x6ZAAStLvXi0d
L4AYr9RYx1QH9PVhAhN56jRkE7HNOAN3QI5c+2E8g0hWv04dVRJ/twGZqsA6cJP2
w1B5uR7sVNB7F686Ygnmfr1mgXY8uAG5L/yTXG6WNXa4uZyhBkb9HkmG8Yhb14fd
o6iJmauKJBgxmZscuT/4tHswzNHa7t8AmndyR4gFqGWivZmobE1cRypCWNpNZaFe
fazjwMbmimc3cF7ATc4EiFGIHuwutM68nvz40x9qppjPJWgwGWhHp64djZt+absW
3pPaMnyNq6qRhcoT57St7kv8POBFveM18ZRZVTVZG2EQU44RpIMD78DY/N3aDwpF
waBIrWymTvlYyiRmocEKeAwPjAkFlZCrGncTgmMYe7QiYKFSrsmCKwDr5OeobAY6
suMvQhOPwJyovs5eMNbOW0YIRDmjlHWQ5PJD8/rbcH5HSZVtYYWjWp60V6Aq03RE
jotGDpPzv0pR3kGaE4wHgWbyoW5d5BzO52kghJojZVC8/BcjYQrxM6PAH9jcJVSC
2hFbZnAyqugM9/tOMddpO1XDJBs99V/gzya4y1pqUseGlBzDZr2hjr21On9pa3X0
RfR2NVF0ib7Ux4HdnwzaJB0bxNWkHRiuSZ+jW5ifmjJXe0I5KwQn/70DrxQVJDWc
9bYn07t2dp3zpPGqloqKNU4u9hygOvTtXChJlMF/daL0UmgFXjs4ghUUxvgl+jAz
vpoYjwLrDTrveh2s8B3z43ScTgSepd4ZqMNLLCWDJIpAxLfcXCG0BMJlrMGiA7KR
DBC0gImRbin9hqQO99384iPCxvdVG2EyqJwBHtSVIy4krmYzv6XLM3dH9U0fMygQ
mLiZA8+nM2CqjltB7XXyNRcVXvVUGsdnOuwR4O5JLNCyHf3+fhMewaKSa0/MrcxY
zmOoff0U/FLjze5WfZpdV12z9BlMJZcVqTMQJ3yG5DEQChathAFXRuVydlw/1gKQ
+B+zGEkCuA3rybeDdRhzojZsai9mr1PLK0jfRwpG3oX3MensWeAquJdQmJ2VuEFL
MVFfKEunv/l7eeT/ffZjxtzH9iFPh2g0Hmj8ZjWpRkcwPpTNc7UluDHMRVM1OrIJ
dp2rLIem8fbkavTR1Lz2PLumpapefv3f6qX+4dQWAeEPyO579gYx87thaAsY0oSV
9dVhqh2WPPyafmZahGqpDQHRaFytXXFFixr9m7GhaPh7bcCOc7Ir8yhbFGYQtis5
upQLKYcY2mCBU1n+GeRnCDUoyoqH+QOQu8QrarLBTpdyo77R2abEwXnqmQLVj4xi
LgQClVRK3rhBFraiZBr4Hr/oHZkOPG2arXr1677KO7E+6jFq9O3Q7Vb9+Yr55TX5
SrYoclNJkQ/RbRFqRuIGqOq1xI4qToAUqUn1bHXa49helQRjaVmWOClakVCv1PkO
oX9esZ6aLqoIzY+yUrquvQKbb1TZyflABKL719g/eJqvXaEKE63m8s51Uw1yqYFN
fCioWjtFHg5YqoInJp1Ens+ZhpneiGf11ZBNH9s5XcvA0c+lHRxLsjL+bpKQPpe5
pN2l5v/FFIQ7j4UQQwFDgJjG0QpYM+K/hnAFDMGYktbLNDfRC9GQ/3wl3So7FCrS
TUwz76kTuAKQU54xgKf9faUwH5Am9WFHoHD+7d6w5CtV541r6ZWkJLW6ddx4WRbn
oJiOYogozNhSfNnD2jRuOZRe4pDDBNSyJxEQROXImFhmM1xngTT641xyEsHDNQym
iKHEmpHbmriY5yx1VO8TXMsLSS139iTCAsX0bq8rMDgNgyxRZbVUZiCxLSdyY75u
C7beDKMB6/BXE6HvnDR8VMUfIU3EXbWuEpaluId/NQM5dreFet3cbH3LacxuGbUQ
aoSctrbiRFclt2c0hqMA+R/8u+6+zfvFXQz+6KHzfhh0Y0++t4fXKWzQ2HrLV+u5
HbMRwVKOt32ICQMNzTBC3I2AqyuqM+qkbhE1mS/gsPClUpVMqP43aiONTv/fCFYl
DABAziUXVSZk0KjXWb8cEXhi0PRSrT5oaM4Gb2jDeFFE/VfgZ9p2ZqMsSxV3EDBr
NYdU/mt6oG68wap40iXU49MnOu3pMvhuyWzMv7zib24CB6ULB+hdHxK0L2hTrbFE
frnKfcxjCO/0u8hxk8dw3ZoLJ6q0fEWPavYUykZZZJtXjP3tDVY5XAsH1at1jPF1
cU4nbQre6CmRHSGzWIv1ixxKTYcURUAoHajTNuAXR5nauTjdK3AmZrAK19rQ18ac
y129cbmANiC+nEeip72gLzM8DvPoyryy8IOY7wkWmG2jVc3+otMfcxf5JXg85IRt
uu5o7BVktF0PAG57IuM3DROCYJY1ZJu1usyBITK3vFM3iZ6Ch7ecHNpUu5n32brJ
1tfHSlBQPcheFKoUBz+/BmE8iS5EJ7Cux2y9NxAfaOk3d+TqZrXdYLHzTWNkAvNy
WUSYQ51OE7OQpN0M+Ukmg+5/O47vKTza9sJk6mZ2rOqgfFe0VohPhZZjsdyBptaS
FJhC2qqHU3KppGlchGAFeTdFhklhQRyk2vUwPNwoZyBFG2+HxiLgx6bfqufM/VZ4
89fwpc/CXi0l59LivI+sMLsOCm+xf42E2ogcm5Ni45kD/Ge5QpCLKsxVerwxbnGI
/8edgwcgFZEqNEdT4SsXBXzue9EiZXxhOCG5gmyulqT1iWWtZx4cDCE8K3M/H26j
kXmkf1clVejnT6zfbjvNPvX4mYhLrNDVlIK74yFlnTOGXcw+66sUCCJTS77J+m5P
TsuFBTW4GNNOTesY6P6l6B4xHTjll/WzcXTU3LiT8let0AgCShzg67IAJ9AiKT0U
Qj8eWDe+oTb1hFH0alOxZWU8ld2dy2A0hxfc8MWwkQb461IWMugz+MCgXM7efUg5
aWRgC6LoFT+eTyUb7YM94X6JurZ94gmOGFVP5uBDcpL4qRIgSvOq3KcIjerI8wIu
XZyruO2fy8foxZnKVViByaanAY0PbgBzOvzsgshsB+O2pbhM2dM4lo9Xbf1Lrxzr
Yfrf/17hDbF4bhz3SZjgiD+e6ZL1BKKLxN3YUPYV2MPBR2ypAP5FnBXleG2YrzPT
x5l4wu/znxVZMhqvh2uU8bPacFWSzNKswXY26GEG24PZJKNt9Uv/bCtT0gLsv04m
+g0Ay6k4hWuK+95+o+VZ4wrNR4BdjFWtC0oVn+BGU22r+h3nJSbMADoMjKWy5Oa+
WKLDg68JTcfVsrCTyTdS85mBEq6RlrfUqj6evLMK+hVsecqmdxEo8YB1RHgtEuPH
WPBFEynTieA5RW8ozLx9G+ynTsLTk1AIEyAoSzyChYazdvY+w6hwmou0vnhExxH+
/wwMEH6ncgEq/ReRIWhPnrIlPD4iYzd0VSkQPYGrC70a4wRLTI60kPNsRlq4Ub2o
yLIRKx0pxAtXevPnZfi68uSzLz5zQllyawa0CowFfVwbQYKwd3vLor7OqY9OW211
V7zmOH9xG/XblMz2LxiDn0K/4ZyhTeIlczL3SNmiPF/LgrL2XN6CKANfx+i8eoZ5
e069Z/DzEKxZlYF8cehVwW/9244cgY/EFwfskFyaJFb2TDlVR5pwG/8brR1Vgdia
5CJ0cJ3dkyAnZxnHFY6yUcvGNDhEyy4DfgPq2IHBrhvbYmTN/D1FZ1CtAyZH6ONd
kcpl7S806DiKDcdpbxT8t8lH8d0Qe9bjlGZ8Bf2SpslLc+mu53VBbuo6C88HUR2p
yJSBGt1QUsFfp/LeHi2AH6qYCAZ9Frol50hql85upp6XeSPC1ZM2qazVotNMei8P
oLgpIGpMezGnS6StWslG6yXhUZHlS2Lu8ZkGOjJT+SM0NiQsntMh/XeAots0ss+0
rd1+Y7xJPLckTgwFG5Hx1ut4QZFytRkvNnqJVislRSogdfClPNd4rVfrwPoTghz8
TAp4cSFWChgTq8FSspbyZZSyQv48VG7geIP6curVawyLqqXa9mhBresWHniL4frW
gOpCFnUiXU+mc93TTMzY3D+wq25NaX7SfZqvblseYCSnemJ+GO12XlFWlCjznlYx
4D1JCWx0zKQFBDwoPYJGJgHenSbo+g7CSJ+aEEQ24WznAmgXggTUYJLGDjHArnmV
Fv4O95QVMIfg9PI5WXEgJC49AeJPb4f7d+vq5VORk6VeUcHWzaLgwcygXIih+gGi
isIBvxLTT4RKBXxmkeVozg++/0021Jlob38n/3+7IeZgOXzMYFbDukUfbMavDvHF
BYNf3468ETDAcXQWFg9QKkC1e6VYUGAU6/GGBywBvSpXPBJ0HfMvKzP567L5u+9U
CZ38kApooiSjBfK4TnHvwShDHA5SmwHJ5tZtVyxW1s27hvjf+CuM0Y5eIU13XHHW
mTJv7kCZ2v9sfWUG5IwwwaAVX1I3xUWfh/dnVbck10pDyklpc9Hc0X/dv9mJA5Wp
aDjQxdfr+n0IisFCUNSZDZyfEQwYMf7S4LmoOkRmX1wDtoVb4hwbh6vEn20w8ahk
5LOycf17sCKKwdbqmdRHQSIK3IvWPc21MKH+HDieoxDRmeFSPBi67cEHpESSbZZV
x+rK0PRmIgRKNuxyDmsCevzIw9KvAEM11rxOZ6TuTOFOZ01sZ9R89m+lXBOkubl7
FXRTe+EIuJwpjruOYylqrMTDgzbMoy9DA5WvNgyafouFR1eu1UMpXiPT2/EnLsQM
HEpIjs7MUeFT4FRvhoAH8fXAo9pzKhjDUS0ybaX5whhOl82bQaqP+uefc6ROHEKd
dc29szEGdpUgvU3bZ28wM/jJgKZLfOtjtxhwd3wYyN35awLtcmtTxA7q1O+L/fLk
vxgwIUL83wizj2dQI7AQylBtgynvSuv3pgRA6QtGjHaXR7Sny7AJBAITj6My7+4X
IHwYfZ0FXlW/E656F1mUHAP96uSpfkzWmzNafAkrlWVyNh3Z3RXnExJsykHsbR/M
8idjtZNQYpIVr+nW397ftprwtwlx2sD8iO4/7UHU2ftyDFS463qyc9qKFipGMBT5
4o+ZNzQkxeWXlsBZin5w5bS33ShtUIBSqgz3Hhkp7Z0FbFmnWm6WrNho7RQeYaR0
v+egcAIk/e2pKH846Ws/m//aIzSlFiZKlZa8aHJYObuKFNmhqcmt5bbOzp+5on4R
A56uySQPK+l+ZyyiBzmHpxgELZijV2Tytwc8zr3YcGbx8QC7mXMMmevPyGMgWZoH
gdQ1ahQ4bQcHj+Qm2NVWvmjVJPIYdRGP3RoFycxFxSvj+UzfjPQO9JeJ7sEeqAli
KDHPc9a0X0WHSnlIUhrbW/oewdBL90ee2vAKvVtEx0PGKKdvCTqjBemjwJW3Agbs
elNiueGR3Q/c9ud+Zymw67A6S1Bxvt73ouCLJVCdydxg6TbZn6bFcYAIeQPc+qjt
pXeNqP2c9zMY6eBOTDL2rHyxppaxsdS6gafRLTAUAogvy5rDEt6aliWW9monbWRv
PzLRvnhmelT09sGW6OQnTN9F3O019VSYhfI6kcJe+0iJj/i1UMi0mgSw1bnlyYqt
7Xm53SsSA+bpan4Pulr9TO05ZnmEQhIjWCCkqNGJW+aSVsfflfCVT1wqoVENyniT
1UCUQ/TEexks3IWrOG2QIcsJGKBKnJcSSQqYbeDyICGKBc41DZJuLKy5XpK2s7wh
Mxk/k2mRRjHfMo/uRRiLDbFvovpiIWu4JnZXIfsJ+hBmWXCeHVFa/7jU1mlrpmeu
3gE8S8SkrjXZDcKd6fTtJt6yhVJ8lCUsUDYYe0wDR0wXYJiQm/KjgdClmpY3YKsx
xs8FYgQH4v4bogZRzAbHWDOmot+bvbWqiWpQUm46OYFqcx1X+M8YcEWdvqsQM8Rj
xpmrkHqYKwNEZZfjTmm6+WGOAhNG6d84dVZZKXmUIY/nrRgeDdH85+nd6VLLqGCd
aJqfL+WQyXF3Z29yu6zHZ1L/6IXPTfzyqrh7Sh0WFPjdse05GoXNs8qK1pLYGZqc
XZtXultrLYu0UelQvGrREnEzE08iWIskfRLLEVJNPRINbnxRqI2GGYShhUsCaESD
qD4jTcaZ3L5aorfpagy1mzUgxoQmDtKF8KoTb+WhmEDrUicreEDZTAajNPtBGld/
Gcj1SmtjnoSaYuWR2a1d/M7Fne8+/otOLxqItStOyxUIR/nTRFyA7FLT9p6o3MU3
pc99cLkQHPSeIOze0yJ/g0MGbgOZtR/rIrFNtXW2vO9aGGgYGam5qnqxP2pWiKW3
XHRrCGZf2w8RySO155SmtzuISVig1ZYV7Idqfmnt4lkYiiEuKECBuD6CVyy7fxUR
pEdvM8mag4aMjEzu2NugWsl2DIOjBP/xBmsnIAMLZi+BDa0728m5mfNf6YZf/0iY
sJvzJzkgsBQOHUL+m9Dz1izy+KRJJblpZ9pNdfH5KOL7QrZlrgoJ93uoaBm792mR
HwkuWjDjH3EMMl3I0n22fchusvpFUyUE6i6Syx3llc+UoqyoB5Egq/bqWNbhbTCq
Ihj19GB/KkmOIvQu7H4e/qkWcBLQmQjgZtn99aeS3C8GCWnmWN/nPAwayhW0aKDU
FGvM1unkMowlcs7WRFOvLR1g1p6DrSrHmB9XyXN2TkQoTbBj8yyyYxzRQfqKxASs
yh+M7EdjuFny5CCbfOo+gsKDzvhC0yll4ugnP1aRCgOq5x2trYtRi5R5H5S/CNUD
FahBC7qWwxOnKVnOD/frowxoaJV6kmN+BpKGOd37BCIPe0Trhvj4+X0yneJ0w/+F
nCLPUCsDaf7h1ATNKJbOLBadTPILxrm2MASHrFMNCuVifcqFjZs3HsCkExdDFpyE
mO144dR/XNf0nSehEi1yuefMvqCkOFhUHZ/9LSTyXin0YXb6G5XYibtCIax2yeh1
FKRlywTfOocF39wNisQ/jHDjMOo/eyCZ74MpnP3e0D0dA4ZgF5sPfCkHxKuCUxlU
aSylAEQV4eu17TGEJrx2JxxYxEp8xYVA4mJKGf/PU8vfoJonZDLi7QPB316Bt2mP
ArfennsRccaj/KPu2IneZhlOga7TLQPzLREXklY3n1NZfhqB0HRYQXbuRBijFep4
VHbNkq00jHD6Nu5jQUeyf51S4JERAQKbvOV1IAWBMoolzQujpWNPtrfETT57pg5Z
n8G38XB6li8bDfqsqKYcpzkKsMJwoIH1ykM+kh1aOW9yP/tYPOs8MQ6LzJ+C3rap
ZrpC0+6ihEH8IGueXW0qUgIGIJ4z4bwzq87yeRFKkLOXZ4aG3GciSlPu0aaNvX25
8tY6SOOXXKVCcXQEC89/qzMJfDjPg6qfLHo8dy0bpPZJx4vb2mUC99i8YIMd1f3x
6QOKmfU0eO25Izj39O4xKhgSQfOa445l0698M8pcawpksrATUrMy46iPlzt4gACX
4nv7pgLymOESQMkyJU+cUsSA2jR35/tMkZCMdacobo+OdxzvkGb1sa0I/cou4MwX
aKwcbrN8qD29M5bcXggSETj8YX4+bn4MJbHAd/3zbgjfHdq5R79uxW0lt3uA+Ksv
StooKrNxXKk4TRLvKpkAk4sVIgE+xMGqg0UhZJY8rAH/AnznNvN+4jhPXtFb+97w
u/ec7A1dFFkJU1xsX+p7UdiqvKwtAm4QVZRzX8RHYgPWexEJNXFYp5zmYUQXx/7K
z607XUjdbp65Bus/NL1S47S+xgtAiAHC9kZWmJAJhZEZLKsZDvtXi5kLkVCz9AXk
6JuFrbmVPJvj/Ksu7p4+Mn1o4xDVuzpr5nfYxNJWp7UhYBDwFojlQBm3fm86egci
g955vxd7po5XQv3OafmFD1yv8fwpoIB5XzFxauf6m5YgS51sOghvW+oPorqE46+L
xtVTojjT9XaJ8f4RjrXP7zV6eYBtSbFGAVyeHSCfYEPWfljOSYiY1+6PC1dUWHWZ
pUpPUnglapyJaSx+TaSFPF8V2sTaz+Cky84XDq5rVScrJPbMRZxHXQY9Wh2XGlBc
xRH044WOuSmFswJEmIpZ6jr76crrGYIcs86gPENUsAnK2gBvbR7SObVcTTTsv/PR
uuSr67qjgkSN80K40ZCH+Afg97omau5zcUm3B+7ibwho+TxNhAFxo+pBOuI/Vc78
0OwBKRY/PmWmpiKxbbhusPT8wTMwnj6FCHVUFI5zrbRJ84ipAI242H/BmBrQPeJR
SQ7npSW/t9Ks+syBKKHQ/gAePYF+cHTh794ASqlb9+UTSXqMIm12fLcwE4QN10Z2
BqlnFPAAs/MN14LMmjDKpSp+YIlW19qRAQIAJ4VVFZB/BO/pSDvH87oQUgq4nnxQ
nwRFeKjU7aZpIUfgy3ivaP+7PKwuNuxhpuzTk98QA//J9FdAhXf66mSBsqJFDJTD
RJr/WZlhySWI+V1Ox8Xt/2QVM/HdJlpxrvcwktkRq6TJmTyBvE2ePFzhgjMkdtCz
ZLu38A3bRsFm4zLjMR6M37gghzBSJ7BlU8JqhsCF07bF5ZYrC+20/xZ4DfQ0VjXu
Rsp5RxBBV1CnwHNeW3+b/2rwqd8YNkiex6kMdQ5uW9D/e1HF5GTjZAE1CIgCbQlw
7N90E/kcIDbK45/ev9EkYBcSDZkRh3OO/10dhVG1GEkAIOsEqS4y/sWjPG42n2LD
rETgVhy82seV3N6pU86tORP/mcqdiysjeDcKwgVLhhOnx0i212Rr9IL1vJ0OHeCK
4Xb6eyAddd+ODIrBZAZYv6YlWRvG6bNh7EkVvasZ7h/tWND1Dal7BfVNapNwpZ98
EXpgZHo3ye30/mYDivxX4nJtmgGBijCuAc4p4c8Krqgs0lNWkV4P+uXCUMXRd1rr
r6/kctTU/O3BumLabWkfUekubs1AwNQv1Lk2NyKrZtxHRNvlebM8Uq1FBSk5CTdN
nBEhl4eZudnrRiPNJGWuGobOeaSV1FycEK0uxYmrfaPAGbacmI85J4myDxBQcu8J
SNPCjVEmVQsNrS4wGDz9YAFVVZO/bbbgHobzGZQmel0lnnd5J258gHoo3J2Zh0i1
fA7fYm4R7d1ttMJOpv9qQz6rnKEOG+b/eS20FBTwlRR2xEJHQjPQQx+uf8afr+jo
X9Q9myXxajDiZpVKn+NavnZjM3SrhVDWEmLYS2v2qnA3DGxMhCrQP/T2rzQSDMSw
Ak85SyIETBavQlIaGHQ7W5qsEVyYRYAEfUdBNeL8KfHTTY5bpS66GXoSppmTcVjw
WBUFs5LSnKUwaCj8f+kI2RHBhkCApkhnY55u9Bb1o/AM93YXRzotoVhoa+Ou9ZiJ
u+DeJJgfSdgfQ8JWStkih1j9u0rrgidvMhpIXuOOS1G/mOpX8OZjwH8YeAwRewx8
X8dNskdN6ytDbF1tvCpPoFRMh0wsUgHGdsTngLYP4+d26VrR2VgNqhLL7LDcdHz9
LIvYOganyTq885onXHY+Et4sjvdI9i+VyUBnUDfEaY4SvvQ9BMuid1cbHVyuL0O+
f7a/H2GcCYZEsmn7YaF351RE6Tjco/tzjN97HZKv2iKbOIYSE2tBFKeYCJkeT5su
Tsy3vccby971lCo/FgTB07LWLLu6A1FPTWC6XleZMmYN3xK6FNqL/xlugslQ7gTR
ksCgOSCf6YKdodnDuH4VXfyZmbYTIWutVdN4uX+EkmBKROqU4hCQ5dm0o/0Be/Fb
ARiJ1NPq4+a6HqCwFFDSuj29FdIder6eR61FCYsoF26SAkTXMui5y737ACj1yn/K
cL+8g5FPULFhSoTBQnsCYuFWTgIT64o+eGJcm84m6mbsL5V7Gi/hxTCeBnHT06SP
yHSSaG0jxqK0xLV/fwXIhAYjCvoIrufJx+k1/gh6gF/Hgp5wP0pKeoyYgPVsta1D
FGEK2Ct0Kt+T5YjUg5Ux+cH704H80cW4nAUiMaLv8EpugfFXnxqi1QcnOWrC5p2L
IUy9J/Z+07893j76eyxvOLAXT82KADmuXX9So2V69mgmYrukFbRM6RgX9XmGfhab
fa+i8RqGTZ+AQ58ZDymcQ4DZ90gEutHiheF1+h6RoE5z8cNJjEp2pLhbZMKAj8RD
E/2i63qN4BAt4T71YZ/zbe7oBaol36WMuI2TS9oxfUNY6xL5ukKsmGzn8lqsJTJM
KWz0ZGde+BWrI6gAi7GpQBjd+ffRIFoi43JaYxlp9laWEs3brQo+u3ROO8wOLncd
mggEYYckhdIpSSW+YsQbYvNDyUjLx0dmiyxWmH8p6L0yXqBuIdrURwtgHXM7CzsS
kYrUHlVnSwJDKkwNugXeDlaj+fz6XYT2zhs40rHRM/FtA4+DfUDGBR9VL10/cDnB
YbruB42xvPyj4xbdqUMKrHC/Hx57z3KcQd+oloPYKDgWigez/8lAuXQt3uGV6kOW
Vp3hRteUuJqMcj7pxRMY6qPJDlbdRaOl7SbRgFyA6fSjEFYX5KGPCg3HEri3lA79
QxvFz/y1EbRlKAPiNtvJiscnN5M5z1HW/9xei59c+dESXSXblIbfIqsmefVEKtNq
NmP5Fl2wVFdXSEh7iWM7bkBDgV8pTeMfOXvDwfkbPjfRZthx11pxE9VA8Sj8gEDF
Rr9iRuao4KUUyH4DGVGogrU9N/AH+uGphE7DScABfJd5jZJkXG6Fzw9syVWx+Caa
qlTesnlbe7xBxWssibRBUx2jhP2H6lI5OCcEOM8ihRy9JL5TbRLAzDrbSQo8xLOK
eWLu0rfpmh3SA6d9WB+sGpBgXHJd3nvfm0/Cj/Gq/h8tpI4/WEpVNHP+hLAMzIwu
48Xi84DXyL0iy23YK8hCR9+1lWhyb/OLnOTYlkFGphtoLpLoBpA+r6Fs9dNmogN4
d07aq4vIMCVoPiBa8LT1ONejrWIX91HLUhqSs2bM/H+Vx1KLU6gdS1UwwiVK1qJJ
pM4VwwrAdt/dnreKb5+MD0TB+bFURJ31DiK6OXlv9Xxs3bxKe+9yOAVmj2AkogIN
YE2+1LmhWOFTqf7OBkF3hbmAxq40lTlohhqp+i613iakmII2kWdVBujVw/oROplJ
8pEunGW8AZYYqny4XsY/ltSbFwyAxN94twFW0BdbtgDw/xjKjPE2y7PHkn76M51y
GAr/8AmP2NcYewSf/xJh0JwbKD9B7gh9vvG8WSyDtiRaZRLAdClfHJrvYePjnG8w
gNW3gIA/HhGyqiR73xJwdQ5MnupXpF89ja0fRj5zjbVXuDPCO5fVzqnhVC6IQLQ5
KECItAEpOWpsNeLl8PIrxKkhjfD04qZ7Zm5OPOqhWkUssXYntfPkeLwF1kDAoa6+
z4cKFO1Ar6DjvckSp6FGuaafQhnJCAvAx128ojXQ0NnWUkv9bAcv8xhFwFIeahqk
J1oLYbX+N8DG+KWeqOK0V8aCZveq265dYZwjvbNu8n09OoRMx6M2KMRsbKO7Dcvl
fZOL42pF1vUQi8JupN9ZGrQFE3i8z75S6Xy5Mpn3nzSBE/ECsGrkecW7RdIZzhTI
TC9QXCPzMVi65yDi6GHHLGeMs8Ofb0HzRzjWkWzm1Px9NQxNlSbOwQLq7Uo9XtEx
pjHJLyLBXT6E58+Ur+yereD7Lwhs/THVFbClUhidOh62a3mEwn+UKkP3Co0HrgwO
Sh0/4mLJcyDDDNAyb58nxMuvbckhzqOGLnsSIcSo/Tlvp0I0zKNBoaBdwgqJsH1g
4DIW7psCf8AQMXSaknKEu8LFaowsW7Ts2WzSRtqQD0SOkR2wQYnaFCCF3gwONbg7
RlTaeyZPZiOg18KveNM41/D9QHAP2IWMdDbA7iF0AAtHETpbspFjONMJ2+VcrF+K
OzJSp2vTXxAX9GuNdMTPbChAMDyvzvyt5PXFbGwOy5tY0HeTD4Rzr3LI85Dr3RbU
hIOWkZDA1zbgC9/EpQZaLuwVa2vWTMOihNwoUaLxAVFP7A9LYFHuJsoDDKd6jRD5
U2J5Uvd+bXTpunSLxY7lECbepmsMXZ9tv/5Te1YgyiGCWFopsLeHVpGUVQ+1pyvZ
cVF7lLP+eMgNgrHZCxaoqBFvL78ebgI66x4IraQKDe2iNRJSTMG4hDaaGb1s7PXz
6MEmYdInW5mHS83lZ3JGCIVywQsSWjJZRzPyAZfU7k7LV9mmQKezZFLyS58R/c58
0CvOz5iZFA0c5SOGQo8SqgiROd3Ag82b10WUD9NdjMIsm6vx5fxmIJ6K+ResqQde
7NmcNphr6bE6QlJLKi1hg5uxG4FiMa7WxOI3t2jMIj68kRWY66akdR4leiKPIZvO
mmPowWzXB+3WR1NrgO67WGYwuyflLlzd1zicHAk16s6AxZM6wTHVfU0BzKE6xst6
XzxpwpFWGEneMgT89iwetTk19+rNNK0T4wYbgYukeuRkMAD+xfrPSyvgf4qSL5Yt
NJQmNHrgLYaeYY32D76a0KFIW85U87S1enCjeKtRZ4YirCq8VecG/FDoMzWfXAih
QT5mmiE2V6XoZzOJqJHX3wB5MC321e8izcXi3CXgtYo52fpAgaDtKKnZKRK+1C2k
23YFkAotTrqpkH4Csgmi3y9KrPQcHCxNgoRnYIbXYnN5UT+MurQC8J5ifIgi52Do
O+d64pquM1ys6MGJ8jbGT9LqFokD5/5JJXmyfqTqWcmm9W8WMLWQ0vOtLti4rSsl
/4PY++ppQCS1c73iUKVGr/HlzGPF8LUSuvF61WdsOOzWixkF4tCBDfTRtWA82j9J
rxplpitysTdTaNIaYJvzcvBuc2aF+Q+yUkAS5p3ucW0Jt7tahiotGhuIh+1piLTL
Lq/Ixn9/G68symdXh5jq1eyYNQPRhcyg9YFZ2Txkq7+3Fk9iYLteWTmUqS2sTqxc
S3+q+a+LkZPidls68gxDhwdLjwIPJo0gG3v8hSIKbW31ciS1vhBI9YxeJoTrHGpm
pF9sWNcqNKk3+GtB+SJuS5eFi/C+EHODCf4rGYpVYzCRydF4aWnJQYBth1m9/J+Y
FhWI22uxcZAJtegZ3TyzdF112dlqu0VU6lWPAuK8jArZKBF4fwQpMyhsuwLmZPUf
h6rWJu7PYfIqoxvwHZ9r+lTqXwov7Irf/u2kxq5C9SeJFL8ljn0lu6g7N8Nz1qXb
St27uNGjQ+rydIs5a6wE7YerKeQ9aMlcFd8ibYHUZk0Rdm4wkkns2ciFZYPZwuee
1FU2cm0309kLuAMzmd+ZeY5bBw5SZTFD0pCrFHaSkGSkGKxWSZS3roSAUBpmyDR4
KepUahbJl1amtOr5BU4iP9xm6ImEppnH1req9ZquBSLkQ1FXyEZV/hI0DHAqjCfV
uRi9wknR+xyiEij8iezuPD8tYtXvi4JoR4xBZ7+95mdxkvcZcleUkAbwk870SCnF
vk5JNm1R4c3pyiWrLkMONpWpcHuExyTMy57SUS8VHdrWgtr9eWXxhy5om6ph03T4
rTWI+vT9egnP8E7wChWnl3ZgYh8l1MvKkNgPAC42Fpplw1udN3u5En+Dex9xY2YW
evHbIdi3ls6k9XVNkzQFcsUxPj+t1GudUgpfRHEqzMLHiwuuPFycvmbyEPOwIQn/
1fNfmLJJr7hFSjTjKn3QLitaZy9Cahon5AAcHjfRyUYcey6cZ+zG5Grq/uLVKacW
EoKPknFmlZJCsc7EsEbdG00U0xvSlvRx1eg4W+uZbFwwhBwztAgg6uFNrbzN6SNp
sXoW8vVcauXDwAMg04bGCERddihNXuhY8ean0gONxL+8XJXks3Z3ZlrhGEhV1Osj
hBXmoR9hD9ijYg7AOSIsXdSXXXxc5jPQtiWmWJIuvr2qxvAkmNjDFtGD3OONs6ql
fVZEy4X2R7XA0yJrXSUS13OzbeG3RcrNFfhIZ/xJgrnQiZmpZsPi5CjADDqawv1G
f0qGikW59aS4IvI5cNQaiGg4IOhIRtMI0MPBeWx5KqhfPJemeQNnjbkLqu8kqU+a
EqgRu/Bnd0ONB2cvQACcBDMgM7P9f9OoUFwInmaBBXbYh7pnSkPs9v1x6u6ph7dm
9Lr2vCo7Pljo+zCWmNl1vGh0o+dWbGa3FB2+K7N1wtfPzc7xtQNwTg3cKxNksXYK
57EUC6b88REH7+HTXX35RyYdDA4VLvCnq4g2U5Q1l7mtHQngqWlqJDSsAKhdZzGe
DS0yydiy9rQqEE+gp9Lf0o1SAPKDw7BNeOIWO2ZZDopaDmXqc8WdFmtPb35reGMk
t4GzQIFtHTSd6kDwUTGjNNuYSXjC1rOZAxn6c1y9C6LJmYLr9hdjR7Y6jvWsKVbb
CHOw0nrtbuOlk4vebUUhKHj/QRVZRC2QNOMtKWpu2iOBN83H4fUFS38aiJnYLIHy
xpQJvwMuSO18KLjJnJFuT1ekz16jmm2kS8tvd9jxO5XqL6mtH1aObaKgVWPqLs0o
1FgM63AvObGK6Tub/1dklWaPBT0LCtGpnLScxAtcr1CToMAbgNODdhxxp5Y4H094
r4IyrbXQavrEIoy3atXHaI9MJL4R/K0SFttcBItnd4NK4JwuSZWYUZOv22ZZUvH1
fpBRNRPGZwC41KB9A64AaSEhbJDcLArJ37fa4rXJbX+5WvcUKkAlsTJBOxm2b+ku
RHVz4meEYwrbGsGTWKoF7QR3TPWagzRqMUXSjweWTuXvZiQ89Myk1MCDXXB6sJYq
mPpyYPVSvGxTuETXsTCBZitRoffHwq/LZA67X1obpKk4FM18rxxyfvC495eFbssp
0RJ+uiY6sHFl6JrjjS1YAMypu8X+f276ts32IJbqE7zddpWZt4+nY1tzn5/PiczB
28Pdh9qIVHAQbnWPTo8G+mBaj+6wIyKNgiEZZpoegeTMDuWx7+1FmOI09r67LHED
ipM0aal9DgjLDP9d5dAMBJo0Kdo4REqoJ6RsiiSSO++WtTLLcqyYeHMVHmUGyd3O
yBnpDU6r6lmB4fL0qQzTBg/+u79xwNXLZpDMb/8mtJezl0bwcxM9ZHEAh2Oz9wJ2
LA3BseudFlygUnX+bhje/THLHVuctPQOlTb4re/upNaLA9w52qpYzi3ci4mYXcij
SQJF8uwhCWdUfs9gQwlwX8/6jHjgcUkyO8A7ZakUzDXiHsVPFtQie/UTeICjhgvZ
OUzCreu4fdNwywr6FoQPb/aeYJje2NwJqDO3lWqdmEZaH6NspFR+4SIJI61XdtTN
NNO6DbDLic65UrCmFgCLKrWYhsV2C8DFVXqhQ3Abp1ZhzJ3ZYeMZvKHIxwY814D5
GMRPPbuBZ9Pium43UzKY2Dob3eswFlOlf90NqJidpsbr0pXqT/PUNlu/f9quujiY
hrcIfozr9Q5E3FXcgQf23f4Vf9ycYD4w2BLbvb1Ck82ZxnCP414Z0FoswDHmoy1J
xzavuDYLq7+hgY/i3eWJrGKT3CS4NvqEFZR3ejG9ypC3sWiKzxIQRFOknCdMZjO3
8u4oaNTCdylTwrFJ89rmZ/lthO9V3k8vdIon/nQolFUP2v1uj7ZXvJq4Kr4IUl7d
1luXHgNUW8U3sanjQa7lYrL5keNh8tDsnxSFCSSa3zf57xiKmxKaIN/kCo+TEhTW
C2FxjtcMV0IzfyzRtOUxZt0vdbSSk0fAgPk6B0c/1OTcU4mpbfPXokpjT56hZLlq
urKQXZXXHJpp/JigxjPcQnt/0L1H8rVa/8DqnFIKB3vojRpYlUitP3AjpI3/HPBL
9nCyGEzaMi5fxR7aVoVeg2CT7GzLltZWE3dlvBljPuJzvajAmD+5dajtuN6Vfgy6
ucVexZre0PFigerSYUHRRw4u/lTQX83x5BFjVQzr0jPoTz/Tie+25DR3qwpK/9Dd
9+1XNJ22e4voKznTo6Ditre9nolMrB3dr9raPND+MDkAzl9LlnsjAoVwN9fFfb7g
M/2JHXxlcuSMfOxbl+tdS4qEUm4bWJLyFd6mirYEW4w9xcGszTxvdKwlHOGqBKAq
nNBuvKMlL04Zf5+gTi7TXwA7vEDznU02n+XDzW0nBH2AIEK3vsvZfIgLfL+f0a7S
ZJm/R65+UDH6wM3YORp4qP64h0B01Ia9Sj2zWxNkqCzkWP9kEItqSP5dG68ob/0b
Euag2ZwH4qAodWNOfH7R96AErAv3WxED2SwmEajzptaXwEzaUXBoC4o6P3CT9gQy
+zSVOnk2BQ3zfRqq+AL2vVCn0/1SK3aRgG/TXDY1IrpyFL8ieKqychyr9I5Dg3BY
FgUAXBad6ZuPfFaQXxe0LFE52aD1NGB6+h5xL5esObMI9ziEtaIXS0vAQPJloRxz
ELezJhGxsUbUYHvRzA1jpJI0LrjzwhnJEnttDmrJ6obl/M3yTygexpCmv6PLKFiK
JOlVtnVEpR5s1tJDulsNixs4RXrad2xdx4vBf3Q0F1/p56zDjpect5eYDVHe9s2P
Q65pMG0qHsY2wMt9fltGcnX9H2K48qdXvelIYH8sIiEdLmY+CxMULwuS+BqH2Aee
X5rVzmQwbnOW5vzAfuCiW1SDRKJV3K5QhJsYuNc4ArRIxe+1Bbn+xSU9V2oe+3GX
IpNXBjygwjIalvyexIhJUe7DHOsKXzXnPIPx/yoNTGQDvGh7SxC6vYV8kT5R5uxJ
0PEsXSfl/NlVRDFri51ur+zNb9NPeiCwVJIZVLwWdQgJheGQlZDg0ALgszwE0vM7
VTvVNaARVji5EZJSGQfdBnnpk7YlaoTvQ+O6Wk+2114Qn+MKOXmrNmXjLPIxTJvz
NeFMqHeSEXZQIYVR3D++gqSUPCANnPUDBzqNH8b1LhIq7UtUpUbRsibdRwmY2jPK
x8YkV10dIOgFKsUXiwju9R6iGnINXFDtDs0VACQB9xxXOh1HAHGC2rtVuqD5jnsy
EmedsZxyJ6p+TjRkJMxC+LMxH+PwleIFm8xM94ikIIq2nT+Z+f0BPkFVFGvO+8uG
jwatBtW+ynWftaoq2eadjZ+2X1t5H7io58YJICqea7Te4Cgokhv92wcl3K2Oy5yf
urh9EIoJr7uNMnRa8wql9D4I98MFyATEuBso1+Kl/pyi9aAxW3bdZbxsAFu6RYr5
vG5lGDhlnVkSmnr+80C7vVSZ5HcHxs97hqmnBS1E+4e03Jo0vjeUbOI9vRSa4Jo9
jyduumNE+GWpFP+0ZA7U40GSCpZRGiGdAX34u+KOtlXn0HGpRSjn3Ev+G8lFw8ns
2ez8MH2Pup5CCm+2hmhUZyxLbw9m258zIp8WYl6z5+FumV/FQRvMQPwfUOcpp35z
u72BZoB+AtllW1cWbWlkxuab78aB+oJHYz5IEObliNn4oPSBQlV0QIJ3R2PulQ6j
Y2Ny8UUaRGdY4xatZCMVWDHy+NW+589TDCGGG1TzjeuPxgmSHC+f8erBfFN6e8ho
eWEe56dW44yUqEVq5GWPHA5adKUYKTLW5iXMqiTXosMdUN9Ue846x15DwNMbZcX4
+x/ohMs6jhb03MxyHTIrlnQ1188Wby36lMLI7rdo3y2NjSBGw+bdSkhrP3nNku5Y
ZsbXSp3XEXJsgOXtmFaRYp3AKNSKW6cS5e7o1/K/UyHRql0/Ze4UlwJELH6T4FHy
bTEcEBuIh7iW2g2XTaA+OkRbpCDS6OFO0p81YcNrrQHuy6R7V0qVGUPINZjL49m0
D4bhBpCfwx6i1HtQsEYqL2Jeg+rWMa/MN02PKl+UhE8lGupUV13fSZkhGZHYvzG5
5M+zweYp6yy59vsPid5+ceFHKLOfMtxzk7LATpwhJmeviSTEyhGu8Raf6v8vXIck
ZCNSDCN5MzIqu3Cwo+nWIfrTG+1BN+qgSS1kRXmzHlgbTbO+1MkrSjOtvsRoNC3v
1IvtPu0AaTqaKJXiIfWKY21AjxHSJQohx+YecsfKDcxbj0DKAXTd0GEA6Rs/DZR7
vC+JrJx16mSo2e2FlWcVhYNioe5TDnaQC2TZXL/JoY4c3Tp8SXupQ+7MJ6GYnLYR
OpWvinSkcI9qy2Dx7FlD9tASrp43e0sSBXUGTrGeayBlaz4tLmp35IV11Hs63SE1
g5cMW/4sw6sUGGh/0//YLa5XzUmD1D0cWYSejrsbqzNfHM9l2Bq2kdS58mSxhmJR
7JLOzJpiUc1nCd2jhFmJw1m8sS5dAUZyNbpD6Dw3L8yxFoAOIbQ6Uq32PAvH1/kA
Bn5tSz4XmoV88BpmGAYTYwbsgj9dCGi5uIMvs2r/KCTjs56svXcehOHdmW4lMTQW
ZGILibveF7sazy5iUh2FgOBIOuP9Q7RqupbAsfqdkqyuNKe2KUcZA/ZdBBIB2Qrm
atw5H4NC0jc0kQhzyNgaKP6aXuBoRKmHJU7yYj+1goLVCZ2bVzmD8Z5LoPGK8acG
66MF0FL6y1TSQjSnlHUlBtTpEZzeCJI8RF+N6AQYvKxUtu/GpaAIVb1MruoOPCHB
/+ES5zm50Dt6pp7Dmu/4HUk9gAFMIlp+gHGetaKWwMeYJjieIU1etFSBsnSb5pQ0
a2zGM4eYNq94MrdciQrhDHnILzTaCuuwW155mlH7FUe7KFeY1pV5c0sZjyxg3Ht/
RFmXe60AKy3dcPrdNe1qkyMYJ9VVYLmFFftDRjtn/ogXu0513ZzQMCxiaJvw7MtT
V4CJ19/FZm0xXvqMq1nwlO5j8FWl6PqDfwz67VeYYga9ZDPv2ZvAOfTOc9Gc4GIn
3GEX3NWoJwGTbesZJrI82GrNIyxx7/qNNQfLhAic4xZyhFFm0zHiNqpDNPx1eEMd
C90PfyHGrtuWASMiOw0zMKv1eKmnBrXLeWO+lBv/txN2TDLuLIjD1cOgzBjzeGuL
AZrgmYV7j79lwkChFaZjw2JNSMjBF6NvXCrQi6n8aiIlcQikNNkeEroZyfCUFDtV
6OC/LjuKw8ZtUVnZo0DH69d7WHpHkygLOiu/OHrsavmcZ4ofXmXo3jgPsjYHgHer
joJRk9Ond09+CH/1DqH021chR0NnUUYCJtpAK+ayS6t/bZefqFfJ9dSi8SvS/z4n
kODtaypHhbQ6PZXl2HoOa3+PUei6miGQTr4pMveWJzVyqcCYp6TuwfXHLLq/WVxB
HL8jEABYEstRJq/SL/9UEzAUnaMMja7KTPET592y1Nx6hltMv39oMPhwr0zaMeK0
Y740E5KO9AHr/ndF2J8usjLvxemz0YW25/mfxLRxtW0c2AAmq8X2Q61xLuO1pz3t
AFLQCYNpME1mHnq3kZU6eWxgFPipyPBMML3CK64LpDvD70en9Se202/nWFx0PIvg
hP4hkC6DrjvPew40qx2+NQjCfkFygoiZ8X75+Vn7Tv93hRE4yspalVusKa8UE8Yq
C7EftudVUVhXakXb+H3ha+CvUqLq7ib6ZH377yVXMuhXUBZEQW+Izp1VspqYWWIa
xYoKDoKFjkwu8BLWDZp4pc8rSFzNuLQQjZGeqR3vbEAhkbc1gSHHiyWP1dc0L86t
zU2rWMO/geZJzC3UizUZfp5MFgJDSdFWU4o0oDXTWHOrReiVtUvJmWZlU//b5ahJ
PiwIf4Se9bO5Ze6beeyoWtip0niThL4qwjEMycYUi23IwsgAMfGx0jDPIUav3CiK
a4UN8zp62JWpbEEiggEXA+JDoxRQCON0YVuX+Z49a8LgWmToEEmgPsGexJKucM4p
xIbG1H3nRvD1eI8ztN+LuEZINm+VrKraXFNbftIEWba7gun7ShNohncxtfca5+0B
qxbRAPw4hX0lwI/v0EKb2bROlhyjcvFqTcPd4LLcP08/kgwiN3b09LGCoIiJDYIq
XTQkuHQ9jvXO5SJMZqVGsMmc+1ZQ+TQsrrkDEB+AeKdKn4MGSmqbNPopSwJ9oHuD
ZqJsZl9EO3OoFEDgRXKPD1EuQe/FTXVq24+EYMebAlOy6wiXpPj7+4uFMSlT2Np8
ATwZujUhl+Eq97jrJ5MAJVC4a+GVRU3S51kQ9wUDToe2QNoKkEz6t1ejYGFvQzfu
rtqKhGtCkABRnuS6DGnF1XyYhXkO7xWIfYuM0ekMMvyuGL4ux8cKN+PRLizKQWI4
U84SBRP+O/9kpxCcnplD+3yeRU9vAtzjHaW1y5QbgR1MI1/he1nSoghp2qxW+Jav
3BD6C5lc2I8jaHg2/oaXxSIyV9NXtMUTTUk0CBDk4GSGsOrC3ZNTnclqRL866JX9
pCQfoyGeovSKd3/+SFAof5pXhgJdafMGCrpXU6EtZG6g1bAZpjLUxQTWhjPkTpTJ
8kX/sVHldyXTW0mSfvmF3Ho5qF8CdWUalq6CcNYSP6b3BD77fdBztCNWQUifnYi6
7NJsDhlznW6HxAlaWy4JEzrA0cy2Vg9KYnTqG0MJTX2elmxrxActX1+xZKZJGQum
BLmybJvqQ8LPHvggygEQKUPxh+UYD4nzI2QO3YhlXwW0CdlUmNNfOTxUamprh6xP
iO67iwyOSp9lXQLtmNJGZ0YBXWwXJieotNnIT/uY/zkpom00um9t0G2lHBCMkrB8
KMSC04majXd+mk+gm8Tnd4axPvs9MwyIHtO667XcPl4bl3LnYLb4UZoEMelHVJDZ
PQFq3ZJBjSgLxRdUHt8x13tnItDD4qwXZ83LKPwCldg5k48aX3CGrIzdtaqFK0v5
0uYIg8FBbzJbmnJvCe65PeB+eE/zM7JzRSSvltOeHcSkN0BWICKq7TADysjorS5I
XXmJYFkw3W+beHy0z5r84xxNS8OYSQmGWBhtm7RB/XvCmPdXZK6MX2GZzLEQuWbO
D6sqrqzY/nR73IPktb0qeb+9qZhkDIhlsa2gHq05HyYM9nfmblslO/t9FZuWOl1E
djKwUMq4nbBfLlkZIMP4S6clsNBK4tG9PLGNF2uU9GxXzPlIy86vrPzPEFpqAn77
mPhu9XauBndZ5TY3CNl0ERt8GroKFR/0VLfxyFayBSLHeMzJfWxi5QykgWB8JxDp
Cc3AUB5kwEi8suCARZG3oJqTJX78sJGhw3S0l7nPwiXfq9hKZQhxO9dw9to5rqbX
j4VRYgdxMvxQhdexepbPBnv44yDR90zailvh+pGF4ROj2sztkoPFg2AMj5m/u+qJ
ZZ39/TAoiOcnERLadBXIQ6ON+Nj2bbsbA2ZZEZGRBG28+YbWdTefp9ltgvswK/87
0L+norgCBzNEUtZV3D9JNWxFP24fpdElm4riPH636p4ksnC2eYLI8TX7S83PbcCx
EQfv06H06cYGWnaDMeX3+LQZmDdBCcjDDbCGhm/dzaR3p0Ulu+q532yncpBzod2Q
rJGouoNW01IPq3pvknrrcxhCDXmDuw0vGXkDSx5nJu9CepcjJgZXpX6cbTCBVGTE
Rs64oBH9Tdnx+D0jZZhyu0EvebiKWrOZyn17mbhKfSutQw70LUX0Sx1v16vOcWUm
8cUqZ5g2VLXveAW+VIzlHf/17M3g/lVhzgUJBkfg5DY9h9kjG8j4kMxJyMZO+HJ9
tH+rGawskgmFujeGSdRb8YTp9dL2xKa+nnU9laL7mRzOtudib93tcjL9y8KY9jt6
PUhDQbHiRnOFMXwimgouMm8ZAEDwv5SArXyV+EDnRbfUAWrigoY2FD6qJ+M41gZV
bRfNrHVPSCVKoTSiSuoAUpb8O6eiWPop563X2tLdkSbrm4DK/XIhenGwfh6Njd9t
wNw/IGvsVXClsbl7i1jT92nHFUn2o2pC9aAHv1OFquAmwjjvFUKn4N93gc1W7vCd
g0/Aa2yHfOaRHq70605borQubJoG12sS5YR47x09D0n5T0KWSUGxalYHJYsZbXcD
IU97RJB5TMfSFbbho+cCY+I6bwtm+L69tEIxYbIa3Gr1q6F3WBox9dUfH2GEJBQY
RLECDbhoDpMXfYjTbDkLyf367cC/W6Jd1QlAyTNNDhLtahRm4IkyejVefhrjYUTO
G+Z8n3omngbi7jUM6NuUFBWYwUsldy3DccyBj/de7J0n8wVQOj9Eqb1T0JKLf7J7
UmEWARroC2Z94wwAPpr/hjtqQwykSWQWsJbkQH/qRzUVbaKTs9aSB2sUnnOqkDkP
kYmdGviqH8J8mQRmS+HZfUsasu3CB/saA0kVHkLWJP3xt3CKMSdcQw6gxptIrlEi
TxFM5Nn+mLMLMJk8YoS7H5G/FZS9vnUu0T5VSruyn0oxVb7pLG7jDVARUFLsiC3M
/W4P8FMwlbA/CYfuJh3Fun1O7LpaxLI7lM7nkpl9iG3r80FPUfq+/oWyldOTzdSE
NtonOXHJr39e0QLa3lb4KX2DTX/SCcrQB31SIdaxvjtTUhCfr3yyHp5T0tgX3ZFP
3Akxmza29lHbhGhPm+btuhxzrDxAusC+WLmQyrsppO2SdWQk36RP5jF1xdpKl4HD
MZKSb9v6IYOH+ydb3cxbDbFhGFDZfWf9KbQ8pnjp0xSTHjshtBn0XWWZzsAsla4E
vy93qYMXDYy5XYQrLaHpIjtNu2Tbw3IRoBslREZctPlkjqI7gfSrMTjmoQkEBBQD
UH2HfnlkqxlgonZfA83IwYxqRU1s//ztbB2KkD5USdMwEm06erKSxlcv1AvY86bj
YTEPuC+kb09iBOCH6gJx1tomcjPHoGUHgUUf75aJ28VcG/7C8DCnIknUxVD69UHX
4v6xwQpWJkbvX06Lp7wyHsElaPSPHGS/7HusjXVp5BNpK0azSz8JsbLH7DGrqwPl
HnW+2iVaCSb4ieSK0inB5cgvh3jef+z1YLel2EM7Z+1Q7tz2ZAwzf8hIwoaGZcSz
YiDedOfJWV/Qdda8o3uxJSLzlKAdvUWNUU8wuOOzLAgWGuRNlcl1NXbs4+W6wtJt
MymRePdkIJJmQmtw52Gq5dQCpEiE67q3EP1vrTpTqNfv4WnPjHPq6dpp0WZLbKbz
lzCI3A3m2VdfRJXgvCb45ncoOKEXdMbbLc/hOKE0s69bcarNwrTK0lDdrviWKmxE
9+fjvlGhZTJtasvS65UAtHWsigFPraN0iMXhk16boadsXNnPAkQRj+cjzbG43hEu
FWxi6k03IKsKuqtf/oIV0ylCzox9sgK7sChzFHuQJBkokG8vhXv6q/0NMi7+TDW9
JFnsYpmRPnG4jwYRkZw89C0RhNOACMJasa6S3/EPvF/FSeMQMahIOCw/eNGBY3rF
ldfSY8vxyh8iKWMDLW/VOJJ4INew3kiCPpv2BXen2CKJIbypqIkP5n8MZsMHEYs0
k4d1+R1aVhn+MKkNx396VxKefWImTQS66/sASBwIpRotSTLHNCSuXhdtjm/JPjU8
O0zIrPoepEF0Caiw2r3TxL0PhwUtfrAhzTwlVI9DhQCfD1G3X+lWhxslpEZBkrkd
tx3P6GstfTbdaORICuSFAX1Of4s7j/Q0dzNVuClDvSi4Tu3mnTH0UDelwihL+0ON
0949DiFGdr64AOtIfkBHAF2Xj+BUl6Y4cY9Cgh4wDXnIKAq0onSGcVEiJzERIli4
MZcPDriRwosIQgCHb9Ogzd3bs1/VDNdDep7X4KIUnDsO3dKO8vzt0LT3Z70hcRHW
VzfBe81z3yQeLXI/ZPOQ+OfMHwEADy7zE0B/s5mzfcLE/dZQq3W3is2vOqrPxCSh
Y1+Y59CAfsP5vcrRXauNDqZg2f7+YPW+6IVmp61GCJpMsuFLTdfSISeM+NOmMrtR
ocN20tGctcItTUH155mRdRP8k18bMfsssZZFhyCaKUdvfJjZOm3rjz/ZiSYYD3IX
IhCyAMHOz2Y6TIVMi/qm6GgiK4ymu3NwQiRaYYb3EVQyV5srzGQXIxMPrpoGaJ3X
Gs4mnRRxwlSEROIxcwKLiJw0Q1kesfNbsO3YCBRNfTVQQSNuAixVMw4ehEDRWA20
MwZt8Qb+ZItHMM/mHXz8DdTvXR6EzFoGQWKErTTgN79/cyZ0ISP2Pih7DMDVQ30T
QMsS65GRDsQU4yNIjfUBfDgzHbBVXPllLBeCE8IZPDOb4sT4x5y15qgBDuVeO552
ynSBdyU27EVpqeOJaGOOizIHpC7HY8tEh8+8Q+5Q/n9PUvR5Zlue0yWX70czf/yU
+E0FtHmjVPUAJeR3+WRZLow3j31ybQV0GdQxN2YnOyH5FiPue9uMOAOnokoZ/SUn
GkTUU0KoDXOTeqBokSxJQi09yavbq6kks8JOZbo3Gvn4o/AoLNNUdxXx4BZppqRH
gTuIvliQTwudTmDn8Fr8QvPwrGNIK+WOlRLEd6vURGbWP/9NlBvCCxB3BF763sjG
Lsl2ArMeAM+ijA/KugV6IywLaBlP+QM1dGV+8xmn2UfqKneMTBeVYor3wVEu99Q/
BUcVQxO0r7xEOVP2dL4xozA59hUpOKSyM/xFV+OKUF6PmFH9xlWvTZBChRjkHAg3
3uJztzx7PgrBvRf21l8xxeGBeDnoW0rYW/T1A7P6XPhFPqK5vvNMUYgcJeGndO0k
pXXsgCpMIdvSVC14vPbYm3YPP/61+ATpAp/lDC4ELg7n2m8OU4Hs2LDf/CEBTU0u
0CHjCNQBzXmBjgzdgm0ORvULiCUsSGtoqMwzWfBhZTMjC2QdagDeUMAthrZvmawI
mEw+01hw3BGnZx5FUA4JQlKwuW0CGHUe57JF7RmCklNyRrgiXERPPdxxwqr5p45F
Tl+ohZvU5fJmuclVNphKJ4FptmS3A0X/hFZxxnqgVkB3iDW0knDvmbKBS5ExK3Lh
8amgwlO20RFh+YUGSjaU9JCPaH2abxCDj83aRXYCrLHf/wv0RUjWv/cixaojTlPH
YYGDZKiDkkZT8SQsaVWBgaC2v2AJ2TpqxF9x8jmWJndZpGE52iZ7Y7AoKf8q7ump
3PvRxbr6EVj6Y5uo+m5mINizsmxPqw6dpK5bsLYK0y7vr4fDhMvaIBiHk0Ie4XgB
JoQ33SF3gMZ7VR+YquxDNF3oZ+EJ8bq5zCDLwdcSbPN9FSAPqGKDNOAJ36clZYHy
YhP0MET3BYaUx93QuY2P+h+Tzr5YqFECtW9WhLN9xSsLGFG98/hcS6s8asi3W8il
D6A/NPEMBUoHx95RBbV9rppNuhQpVI6KqtpUD0H+CLdNJ5fQzBiaUXbdynEecaih
NIJN/GYhyYoTlwUeFYoBsbMkxMPOKFeWZQ5apwoHRMiouYwciXwyJC0O18DrxjyY
WLu6mJLIMu/YdC2l2AWamkkG8v+mLdK6jB+U3MRNQcVsr4wzSG2iVTrRbaJnRtde
Wz4qGWLVmrFnAThd7y+2/AYJpyHZ5M+WA5avDfNzAcwXMBRr95tBXOWnv1XHpFRP
6h/AbZS5+EhxWLCYoMAd9HcTydObJ0doFRdt9twntatg3s5X8GXR/vyQ4x979ucT
Crds1M9PmdjJhQ41pXKHCXMKZ7EUxdqLdy0gwmK6t5uTDjBdslYBoTBDodZlrC8D
cozxt+YG3KuP0QzQ68hNA9Q2ErE6CUyZSV2w9rYVq/HyZiVCCFq8oi+RsqmYKraU
GpTgDI2Ku2eXOfInF1RboCSZpOxdoOXWqYgaNxWE18/WT0Bm+PAWuH2tj8zdw7nu
11oxszcwutgf6p+AAc/sThyugjlNK/wF2HDubNwMpshk6nI6WoqVKGLt1OG6uhAY
zHA4zqJD4SCBHKRSYRsOv+52/RmvEOj6EsWPnrTdcMGA/bgKQauupsFdD9MRQgCa
JQyi7GJpu/q7QDZJXQeXFQsgtoAyMILgHTkPEkJDPWw5T/oXZI04scdV2MxqpmGK
c/bRgGC48jfDvofKlyc4UcoOAyo2olEn3/AtaV6BYj8sVikEs3s28SHtjq/xyTkg
4SzYPSe+WtcNq83G/PxSj3KzQ2HkDX9nCvvai55nvX496QXIm+NokaLJofDz+AAe
AmMCF8ytZX5Kxqkf4Vq0bOq0PUurgoF0a3zBWHusoI3TpPXK9W9qu8tQd0pifKzW
V236JcfnaAIhFnWoUGFtwqlCjR/+YVcE2vlVF9Csv+hEqUDB6lV5klCLmejnfnEY
u6VjclgUZeC/ms6oLNHQpIhGpYps+I6yq/cDhE7YrAXVAQY+E34NIBRsfxvNvKKK
40GrysuyQT92FnD/y4q5gdKxT5bRF4URGK/BP6XwTq8uI9IGZR2rS6L+p961jqyi
bw5pTtvRLcI3/ZoBI/ESV2cX2m187pJM+6FYNm0Uau7wFjun+vAHYX4APWAOG1tg
ayjdg75fEAra9b9ty6q92UHu7nBBGVpJiijVCT0h/7bJ5ejYya8d8p4cn15TqBo0
NC6R5OKzg+WQ4PEqhFffF5UjzV0GOasVghHcY0vonmixGFkb/Vz/g3GGjjXMm52a
lPL5EvqbWi1/CCUhEGe2EEAc+IPEGdIoXyRWgJuUbRHMV4nytU7AjbpDZnZWxvk/
P+UNvIDAh3oPQBe/OxGoXTk18MTVyggRSKJUaob9Oax3Bn8lB+7a5sKeXYcsLIxC
1qNyi6FnaLqtzBQ3C7mmLX71Doj0jSaQUhZbFNWPsz48yrN2ojDbQU+ZP1xbvNkC
KdoMDhi+ASARrK0/41uJYO0P9pfVgvwrCclm/DSht5G0Luk2SARNGny9VwnTwDGf
VctMHhLS8pPqaj/6PFpH8StUoXOJbSjyrqbYlZ13c/7OAjxqkaDQVBW0si5Kny0l
xRbq2Knu2EqXpiozt2BoWm88CiRk1Ks59OaBVjDXULvc+qnWdRYpNwUJwCm6GY1P
LnP829memwWvefMzzbqycPRJ7MshVqjEDAFATbBmZDzBXMy3xweHxnivKAr7c80d
fqC+9+ydBoFCQyiQZd3m/RGxBac1ho5aW+8U4eA3ey6+cnRBF055SnwDOGuaVygF
oHrFz34AJV3p5zJGUYpz9JfjIr+Q5LZEG/ooDtuDk0g2L8UU0IguaJHaUgTlyaYc
oO/11CixDoZ05VqjfXfsn5LKcBEuBr2N2r7Tf7ePO3lKGDMq2+Eeuuh5hE/9bC35
hat7pGe+Pi2RGXAfjwOMR/gD0Td+91kPosjtBPMS4DB33jmac4dqTHo41r8+nIYD
ZOrzWQ3KiAAiMPzNz9sJJlOHGCuL2WrGO2L25NQ8bLD6u396aEFzixhP5A0cK0bT
wrQpKM5Z6P0m1sp3XgRQJfZB4il67m23q2YzmR7sKGUKYFEKzJJzgO4zIAigKgtK
nhu59EJnwM6RZknZfdwm3T/2gkJwvtVWpSIhdVo8vMIQYGIucV+e6Rh4gVc0ce4N
FY/ZawvE2MhINdLYURG/evbZ10WFwWI1ZHfAxghILs86kIszkV72m+lnHVgXU297
H/Y5jZ++q8NtooUkIyNN7Uwy7qC4Kkau7PMKUTNkOPbEa8C+IYgXlivuCt4Jxpzr
T1Z8xLihAapwC0bKvDiEnYhZFUDmMQzmBxUfHypJUEu4qx+fr0/JzidhEDXrRc2l
o2c4c1W72l87+hM8ZRbrMDeia6z1m8m5KWeq0DYTR7gZ1duzHWcCQF1BuD3wQuVM
s+JZEs9IoRCJhI8fveRyU/3v32zaUDt3eb87LeS83+WgyPgMItirCOjy2G2qbu0R
5klucQgJXySB6oqUBzobYr83iRQVkiynrNCwjm+dFqLxL+bvn2vVBytlo7Lh6swa
XKQheMQ91FxgBfOBThJ+roblY9PIrtpYkGRDxmFgt5cZKdp5tqFjwCbTiSSg9kEx
I/a54aj8CW5sjeLkanKXpTH+P4XQ3uh0lI/AGFJPmbZaOyA17mHx3jmolKXxj8So
8cgcqHp0gFV58frZfg4C6XgBHpSn4kxipB9NgmxGrvSjhZ03c+Y3sGNISQIlavLb
Y6RmJwPjgkDEYcdjBe85wmE6kJGhZPEShL03y749Y1b6ZAXuYqXI0T4A4kTFa0vm
UTvTHlh9CPiRI3jTNanmu77LpAT4PAsRGale7O8VHz7R+LeKNVW1KpAJyHTW1/Xa
ntWFRuU6ldzsRXYeuJTAAuTpiUOI0W0BcPA5PvgISP6FVpM3VBWWDDBZKRPkxe+5
FemIkH7jrUaIeLg6AYSpCcOrC04RAfzKkOVcl12zgehI0ajKAf6sqng75QiUlvHm
Z4GClwskhTMi+Yv5TMNp3VsevCGFlqpPmSo/3DUCGpHOhj7GpPEKYWm/tMhF5cZu
gRo7mk68RibpGHNquBfURsQjUyv5VxBpusU4q8dZZHL5l+fsG3EdqsNHRYYWKhuf
jgpBFfiZ8alFpXWuh3D6RNrAk/r7VyliUbY3FabIblhp0BEXgE8J7/HDqTQsEY9B
+3/mHUrRSUO7U/uf80hsOm/9lZaYJSY03CCMiPRopiRDWWlYbNvB35FJCR6lG/+u
YsY4ZZODJpRS5jvGgxBxTYwcjpiDvC0JohbmafL7Fo7+oLw6gOL8I0iQaiLZ7QJR
czPbLmZak4MMmzmsnKyacMxZiAvxb+cPS9eS/9tX9PGVMG81BNSoVfPGbgyh9jSb
iAhwGJqxVVlF0fiyNe6nOY1hLM4e26aDunuu7eXuLdybM7KFcmVJ+tWjhDlYIqcr
Gu5dGwq9ZrysjjqtYbORD1vFWAXqufUCHQLB581HzjcehTxO27b/8OQ9LgPYN/Wc
fTTIXmDts9Ca2nXyJMtqfod20FGx4SADFcCV2Nd/IZMnM+igfF7ORq1KVPGnpccE
vyHR6sC9jlfcSahplvaMjC+EbD9pywifUMjHS/aS+ifA3yt/n0PiOikm67M+Sa27
GyU6nOGBRMGrXd0a1SUDkyOdtwV4aOG8+1Dy+DEdl2uUpIEFX1VuclYbf/eY17jk
rBbHe1YQErAF979T14qSqK8+tWvGdwve+qhwNNc9OZLNwyzgf4FsYXwTkR1aw1VF
XRbCynGo+x052pyxZhD/21iSU+2rd3lDekCcvwDnOZUB8AhXx0M7w6zhp+Alm5e8
gF6rzdS6SNSZdiUtxPLa+/i4cUMgahOrOSW2H4iDajVNDrWZ/8jGM9JgOFxPbQLi
eB7X2aXUE93SS8Rp8oMGVlx5kq3wjdgOkiDnO0t++inaNyWqiWx/qxbRjnmROAzc
+6y24H4aO1Hj2dKVD7/D9yRcWtXHPvnxkwaWNvnbAJxeoPFjFZxsRheaLySuZKS/
zPLLMajZdZtxTdT1rqj05qIqzVgYg6w2mCnTWR1GDYtpzWE1iOLz4QtU0d3WuVpB
W8aiT9h5ENQnnzksl6UyY0zuwvPwR9CJVNakBT24ib1wFaDVPasldWsetS/nWGAt
pV2dEOTAFBnrYXEVXa3YUA1wlh7b8+dn3mMIn/EBUZwYf6rx4DsGYbTFIis0ZNZT
tmqL8Nrs0I90lthaz2tsE0n/M9M98shBeCId50D6DjH2v68NhFEKiqPFReOSv0MZ
e8YMEmNX4dKk5HzzatltnCr9bEb9sTTRVGtOSw3U76x950eROC2zwO8c7Bh27Axs
Gj3WldOR+46iaS8LhGuJAe6Oly0GDA+ROdu8XSK6IWhnfjG8tmK/Mbr/24zLc0uZ
bSmQq50lIDqiCQ3ymFnXpZwxvcuYKNuH5aBjVSnyzqC3yTM5uzvYrrfSD1l9v6Ct
SzuY5Rx9A8fHpc2iF4UwmxQydHBfvskRBND9w2cxhqzZXooc6k7lIimGtL9vGDu+
C99TbthLnk7ReAXuVkKRAIcwiBSp/Z8aNZDczGeB6hyXOTBRl7uOp3p0U8BQvZeG
zfSHYO8qbq3mnoSOioAcIQru2tvb5FqLtSY35BuhYaBj9nKERd4ErbP5g6uMCNo9
TOpEyKZHmcFtfjpb6sk0sWGRM2h7AFLylwRCsnNS1i6VUc9uOPUUQKXqEdeDjxde
tkIA6tJccPoZp41dsEghRMdXdiX2qiiwkbRbilKn03GJ9tFGmoZbMR2COyO+aapS
6icZhPkXtGQdsPB2pm8B2D7R33bnRuSWefNE7ZINgUxDF/3InyPzx4ubWd5NCzBN
PnSLiqZNolajUtlGTRsEhFqmWSUTAWdKIHziapDvdeCQLpQfL+nPHWCkhpHHLAHM
vYm2d7JSE1j209D+gW42rhZyZf+6e6SZPnEtHBkfDADqXEJrOlQlSGgG4FyRAGb1
fjuU7RHkrbkaMnm1nIZYg/y64eJxKDpD83uPPZzGcX7Y+k4uDrKZrzJw9Ci5f1ui
UYQ24iIjt7fqDjBS1oPiozeERI/ybAuZm77sZM3+aLL0vOk+0RPNJJVDIVnqAuUd
iphcWfJNyIYmTmdpWcJlZzgh2LvGB8Cbk1Me9xVYJBJLHe1m/+rsFR48xd8N/qCh
fRFQjIPek0Jqe/lRvirlhcA76fy3bxMj+MsdbM8ojWxoS7MSMqQ+OcY0MUlmO60A
ICGVb+zdZg+1Tpf7VOTT2VRIplxoP6MgpUbGZtZGBNkC848dPA3wLkmxleTXzVQB
OSkvNdMj4uJnUMQZmUrJN7+yRMMXLWzNS4tejz3ysq3fbM4oUynePrCjK1S5HFS3
832DNrljEyGCF5BeYJ7FYirf6N32WvR1XbRuo75QRFEjCEQYnaJ3CkQve6pPsvAS
PEkbJ61mxsXAptb2z0GscgRvESjoTzBrP0o3VGxJrjl+FEuc+SbshsNJlqWhI5mc
T92EfD19qDRxcF41tYmzafAUKdPL/9APdlGnUnzCz7Y67pN6lsWNAizbGOWvW5re
tA3cmFNKmLAcP7jke3hUxGyQ7mYhaYW0cv6ydVoei0BSX3v5e4BPYOZ6WDE3quUq
A77y+caB5/33VA0NCeYy8kk1qLuU/xzEw5fwhdnVMaqscrOAdemlfg4MFqPO8IBy
f2JavK55BVcP0k3ESBy4KjulVQohUv9CglrxVuZOboaJASJOuzMJHBXzIL5Op77C
lkRb6avk37ZLDC/sskdvWtr1nj8vy3lvRBXHgaD85pGvRLjlMoMccV6/kqNhf7SC
Gr+jGvYptrveoRnbJ0b7IBppSS8tibTXZaLzBVWI0VG6OL+3aqGM5WGSxwEdFLGE
T/hIDVJQihkRSAg1Sj4OtxE4jLrr+YWx/zV2CCdG4rSKA08ZXRIUSJJX28/yCPRm
1qfMLD32k+bIhAXChlV/5YnxUaAeuIb3gR+R2E4YpS6xcOoRGeZsJFHKu1BbpIHT
Kr/DVAhUfBIazHhmRR8RIizfJ6ZclPLlrDMWlulc1ClPLUbuuGmC4pFFhvV0pYTl
YutnOkLC2tV1z3rIQUTcxgAnvCdqxmBxHSqoTD7LoWymx3pFTOFI2CMWJap0ACPL
J+1Nf4YKfG9eKKB04WguWaqO79F7LoLBOCa2dHk1F7ZzDm6dW1RaUrffzNBP5czy
4cPD2Av9eahS1ifVPO/2NkPtOJvhUMBtaAOGYWnGERDeu/wUW5bY77RI8L/yTnP+
hsxsyp2KnfK+O3TmuHObdiJ9/Q6QT8hw7e/Hh0gRA5kefB4UZnwNATPf87HuPiSn
496JUaZOpZeO1G2aWzxrXm0O9C9mS/QEnkHTD5lWtWc1r1XFLt284ayis4ndiXK8
JHdXstjeW8XCgRGjMr65RprK7sOhavy1B6rPyqT90jzdeMbfd9QtGlqDZ8Qzpclb
FYjr8DOQNM4JwVrsaQD4pjL1LtgLkEvpUbRrLUwb+pb4AhghhAp5a3Ckp67RImlX
ERVrZxcB78fH+El5DhHy42XYdw+JTuezlJdZMUBnrN1otSx87YgDCATwSKwdfTKD
fGViP+603fD/1Y1XYvRxz/PtapUjy+UHLUfjmkJY5lwwkxxc+ZnMNZPM1WeuR+BI
PiWgH4oymDAVdnqOTyLzkvyW9e0mwlHES4KDa4dsNpY3CBRZRbRX9ALWJVdkR0Jr
csocI0pGVJorEZKMlBsenKp2qP2eE4CdoJIoH2ajJeEoaM9O7cdXqPfOzS3wzBuI
Y1mZKYx89Qi+tI5FiDt0RglkbgXgaEs5de4UKnHLHe1IUyqHObmkD3wqHR4gpUPi
u/9My1M+FkUjhobMvqng07X5PPUj0hSAML2e5h12pLTWCUkrmYb1HeT+Wbiq8o4a
H6Qg9h3C/EXXDkeef/qaFrqYwEhQ62ab95dJMPBvxfNAdFeVOMSQ1swMGDZGeDnv
ZCaBDZxL5mtdws0z8w5FnTlNqfjOTU5gFpvNH9LWQK8RXco6m/h8NBq3ZAMzxKRo
j1foHVibIsKk5bIXQtyTMBsC/OhdtjkjBor+qV6Vawh51ayWBf+38/rHaPsjfsM4
ICkEb1CsYRy/ptIWhhwzjuU208QRMQBRhPv+VGIjCTPbqhzLFnoVLd5J4mGmCMLb
qsyOUpvVX78GHPAAQz3kgzteGTW8DuRxIKlPMs991zvRB2Hg8a5l7SkHjk/f9evJ
LykUdy1n2+y9jgs9tqy4KMzFoLksfmQr03iJXZaQ5ArxhbHnUNReG3B1qcWX8HKT
8LvpVFTBJlnHElnFLKIOPrfeWa/AL2ABOmZzkQbx0YO6c0pEQiRUTEW/LSyDx4C/
W4YkEGgSIVppjDwYYfCOTdomRlCzcc2RT6BK73gMUIq+v+2AbGxRSAVqjOLqkAVj
3r8ooiqvMl/ldNKouLxa92bQKGDt9eNJiVREY1a1Se7fMBqF0qifkdfm2d31H8KC
JF96cecgX8mXfe0WkDQ8N4XP8rBYbTWXmH3WQihz7y3FGXLGLlFmqSYY800vEI9u
+E6+wgTLBJfNVWaHGyqmXUGjp8IExi872rpJHDlxnFYtcvaRmJ4KDh2ZG/HfHKem
SWNC1TDsRSgSVRIgkmyGGdnqWSA6APvU2efRyEeb11Kv+78lLN4Hvwxy949SfKWJ
k5GlCILhaVboEHK1mecG5fsT3AFcuxyw6hTUfrXisHlrbJ3w4SUKTkgv/Afym42Z
JCs39588zw5I5VH8fqsIqWlI1VZTnvJU8iioUWCgEwqbH8QQGWFmHYUecsppYjyK
wXDFobq4ne63lFcUFVPEASQ40xMX8HZHgVyJ6uWmMO/ze9Gnh8+e2gbsSHfvULSM
RYjmggqKCUZDM6Czx4oYRulxQ53Vyz6k6P1xM6OioVNHkEoPJO1IRGXNUYVzx+5d
IR2T+eZvB1BIWSQZBYkwGLWSAlf+H4drDii1FHftbKoxsx8fprwp2bbKA50Ig083
5rrBaQoBzM3Xl0sbXeugo6ttXS3J2xpYc8kipGoGtiI74i+/fg/Z4N6yus8q+jVo
QCoxKqeTUKVc4a0yi1tf3w1NafQtOoxoOuIL2oUZZAjv+dRyu64WdzyFAGvZ+kxK
f9YpLi1l/PfIjMGxKtS5spL9AxjcE+UvpEeCOhoVuLrH5BTp9AG6HoZvcaeZsnyb
yaSOrx2Uj1ku3NKfZCQsmaT4gPzJHSoJcPXTAaLQnX9/n2bPq8z31PljjpPjo3k3
QXO3gLDBk4+icGwtU6u5ozbR7aHhzRz9ZqoIPybQ5PlpgTUEPu+IBlJilwWfF4/D
y3yMyYRwMcp0UWO8CgDqSoY+pleCCRLuxkASWD4erBIyU8+ovILtCl/6dIo+3oWj
cbCEOIPE28pwPmlnFXjRBqP3wz0z26Mjuc2W76Np6bC5iC+LS+8LIdl6Dpsi8Bfe
UIitomQ2MjgCtTVb48CZL6BXvvac91RVPF4CVLKHE9bN5XJ1jxQalWDXLpVy16Zc
/2ndRO7DoPIq3qIGd8oqsTWNPxmQyWtZzVL57iu8dW4pTILPxW125OThMGR1j5aY
yAGik1khEBSGZqAVUj56gsiNKqtDd3ULjgnHFMoWckDmpx4steQw5wtGU1CTtuGp
mgzvNRE6HsdSbi2trLPlhj4wkIzF1OL5tOQycScW2/WRDgiaCoVQg3liBCwOpJpG
zBYkq+x66N4KEQQRCZLOHneP1kdAbjvc3/xLR8Hl5CQyeYW2UTF3xelJoyppuMDM
1DlbuTdz2dM1f7EO92dKjMy3CIu01GBV6lbHIgLvX11QtdSaSzvjPW0mDVa7wx5n
PZ425+7+OIzlmpJTDD3vH/JNl8sid9X6UwzrMrb4DWH+ou+o2dIGSl2f3njLs2JA
Kz5kqosEbmz662ABNM1mJoW6Yl5eEZT9TuiyFcTjoekH0juJcsvtA1kQJsrcWx6R
idbz3HtDpuoX567xuA0GoUMeM60X9Y4eSYzoQBQhi98USHkIdCPXjJa4I1NvBLPX
I18Wo610/MtBSnv8ldckrKzLvgw5lELhhDEk4BFCh1o0tqtRgk4DetlPhhKsWIGK
dbIdia+cAAw6qkiU628BjXkeRVFIV4A9vUPqF9TqaanMccA8jOOtLT91TQ5H6raP
IObAcpak+BY+/vXvFbsd+RmXaX8H19DEvPzu5ffO8mlTEFA915TItRCCLAhb7rFi
2keMhpfbmSga7o/S5whP1xDIvqttENKnI7iKaRmyxL0dYHh8kJUPISQXYh1ubqIf
ruEVvWuh7ZAPgAihn6N4i2uofS2OAuQdVwJ76rPnD32jqSH8ozyuivFenA3XU9MC
16zBAMQuolGeKApvLGHK0hpLCbAKilvb+yFfu1wmoXpvJ6iop5NNFgyP9l+96HzV
hjImoYjDEZMDrsHrHcdMI5krUpY/nW9S9gaG0nWhDmHQHbJQWxwZPlCjvpi6SeKP
NRcAr7Jx47z2UlAGgbWgC5wMa//ZXe3S6WKjdjLu/t1E/+BU45n7la3VuRl/RRTa
2i35lk2L9BHU4Xsj1jnssr/LqKOBYGnA8cyMxodruKFLltEJPzog22qQTa15Gurj
+jx6w1A+gmHLj0UbcTYrDky70PT+59O1gH4xGYVU2sBI8SulYkWmU0f2jxBpkV8r
Tg8Ejl1URdrnGmrEUcAb7ll2R+P9TAeielak0NYm2WEnEL1kssQTV6w7GONGVDHh
TH9ygiaZYyD2k1UN6Z6Xo86Uy6vB46051QSbLDOFjU54cx3t/oARgog8yn3wg62T
lQZlLF2umkGA94T7krDRJdLGf1avi5zDuOS12IE2ju1cQnP9yDcpGZBs06GrqrJz
9rRVyt9Cx00Fyo6V6Kqyx6XR27fdaN2845YuYzZrMUWeuOShew1he0n/aPYGX7D8
7ETHTLrO5DgnYmkUhhHml4RE44ZOndWnECBLeQZdInALTCtHQVVo48vt2S5AyZwO
kfR4RTw1GEHvotDMLOcA9darJSMMZ56bJS5H/RVL53dEg/oe9zB19meX9m8qvUWQ
ZR93FHVCLKuQxLp9U1fZs8gdRa+zvssT/eDCm/eL/9krp0XMh0vsYUgPbf5t+G0d
IzoEXORXleHvBlrW6ACOKCmDl2ohkROJAIyhPZxjdXBKw4BnYmA9gLjAMGFarLfq
8eG6fClWXYej0F9dh34EHoPRd8LGBBkl+s7bGAyxsVRynCB8mHLzmq5suveyjQs4
5UeK590E4KXvnyF48JqUDvEsaQhgm4S5e/GJj3OJ6x3TM3FjFcUXSAjBbtYyaHYM
ORzizEQ8eRqCiCjkg/UIrE+EC3UH/I9N60xC8/UemMj0+nFqEI8jt5MC6h5lRm7B
mUkMi7vJ+Q5sj9uNvp/kn9vHjRVf9WqWxrvSxRr3joyFJLa1DwFiccJcJcCHv2td
4CtrPoToOuuKGRvUETijDLnCLRBydWsKxF+wCedfR+I3SuoCYGNXJcm6pOnEK0dq
mSsrXfZvXsfPWiCNJtG/IWSw4TvqG8E7NkWdv5J9HovtkKz+a07A3R2AbddiwWCf
pKl4MjnyRksyIo5VSYvhEQOdjwAWTmMvc2eMulW/fMqBSRVdrxRFQ+jwS+g3gC2t
FR9DKyLBbGZH9974ZPN5BYgQlJP8LF5rWGkPmjMFsk8pC6SE/eCvn+x56+ZzO6up
eRRoTJaeNYlV41Pvy276lItWPCFIxyn+H2DAfcKUcifo5ktqmdTbYJOF6FodBrqZ
C7QzFO6x0PIxoCL1wkL5kak2PbzsekrXFBbkIZyokE6CTuo6GNWI95DQcKIDAuOg
lajwH3eWYXnOxXvp67URJ02jlEDVBFgUO7x3pSC5EJZWWGcdOXYxoIKyDXj3Pfbl
bs8+mj5pkspXTf/hp5cT/GEl4Yz/8hzg6rv7O/BUAemCBaXQxdpU8Cfab/P0gF8c
ulj1SVrhNwIT3jw9k3VIXwnuDhkdx0g9jdfKJzpBhIvIx4Vg+2QbFobHeNXOlUUP
9h3rxax01CGLjeoUAAVa+0jiEoVObZX5LuNxAC98067S3C7lkzk0vnBV21OF2cEI
g12MGRu/dWB8kPzWQPR4TXWBjHJieZ2YQI6BL+fNm6YnhZc7GwNxYF4Zv9u4REYI
lkz5OYrS23xYzUL/9ILfJflddTkFaPZwqilyCj1lJp0BrIwoRHexgO6H9RHmGldV
oVd3abjSv4UYnAQbAWi2yKKmSzwGd5v19YQhuQdVFI0l8ChENhrFO8BVfiFMbZvo
T//y54b1YNApMtiPRXlekiiOplsSdsv80MmXPlHGNksdaG+PSzwsclwxugAGNvcS
fJjZzVwnSl+GXCOLXwrAP1qzekf2cPuul5gL5v+CqcPLf9JdBm5aj4ieKsLFb5Gd
DyFdPwEs1Mn7eFkcDcpyJ0YvxOkxRwyejLskoWc9g3ECq9uB9MXBq/Rq43F0Ucgz
2wO/VWHPPDOCdobzp5zaX1RXh6DDoY+WhthfmE4sZHCYEVoMST9Q2uEhnHxQCXAp
rlV4QiWDf7dvjFog0rEsJobyAzVEwdT+cJv0FEdlfWiePOsQzjnPfJtUZ0I6EWyK
fO/VQ5H9uIB3GtKQ+9UjM9siM8krxsC2sgLySIYz74kk1mS3W/TsbluIuJEmLJeM
x3nRIyNSzKyBMdLoJTnh/tZ60yJ4cQIOnC96wkE/eiU/2SYjUVqJOXg3H7YFmhcB
CmmTUmdeUv3Xge9n5SZg3uUn5RpGFz5ZuNE/SbUrYC8S+lUzFBLOawAG0G9066Kf
oY27WApR7KUWQAcKcpnHfkMcuY3cz1Pmb78svnDFlZJIdyrZl1QC0psuL0eYXBrS
c8KEe8xdUH91R2EN7pmP7YE1qG8GTsCfbRpHXQwHa/cEoTIKFFOshhIGaa1BcyiZ
f9P5ThwLDLikAmtvgNCdkP0bKiKEfOGyQQV6KVAtLFyl51wa+mD0C4Wwbe5IB5Ck
DFqWYPw/GTnhS6xte0XJ/JynPRhvKct3/5Bq+9i4wo2ivPcOtO/dLw3XoAdmPtu6
xx35+Ut5HWlHOjD7JUj2K4EC3Vg5es1IvzdrCMvaMBkEi6493UqUx3HAa5U1gaTU
/i2RFlV2VnyBmBz1fmJo9UwgjNSw0HTho7xl+I2w7e7yQuqbrPMxXtmrEP4gP3Db
aXJ/Wq9h6sdae/pc6eZiRiREe0MVPP0OUwfZE0na5kEK0RHCGNNqZl663uKaCmju
tPwmkYYZvWpPRR3YvUEvbrZWw+dRSZDJHG3mOTNN6yFi/xJqM7uhKtDcc9KjddwI
3cCMQbNB2zRHQD/BPTIz4YRnRLR+zCyxjFNUflphGGYgkbc/X0hWb7hWv4kyRefE
EQNEn8QLla1FJCmHkZ/xKcoFSheRRioKEpobpAxqOV5gwZZU34i44LYn0WZrgr7x
Ufkxwwy8MamNQkICjemg1W1XGuYWETvpDwoKBBid+SE1yviZArrGUCKrN+A47YQt
RKbM4Gta0qRcL957DS3Q43VxaBbjYmGYlSjeNoOU5AOUje9bdrbLv95GsJCmkzZc
7khaP0J4KV1uo2jnVVWOYrAopXvKcO+T/PPVYixTRW/wnc3CZRRI9/+EAgMZmobt
yFNeDpfLAF1aVACeZNatLJxtm9bN6dPlOgvHsc9hvCuq1VcPorMHsrr+/f/cWF7t
2SxLYg0q1Fe676SmBhg1Y/ggLe07jrCoYMQUk0qqmeB0YEDwkgiP0qF5zhhdFRLa
fy8wb+AOubWdKfepLHZWKsPZTKPMG9D2yqrDc58mz+noeLDHILJuPlHreON/Exzt
RljYwAO+8rOQdxWpccTj0lHUczPPKWOLISdz2B+ZCV7aNaBmf+tuFg2zokgCjMas
fIZEC+HJfVB88DJMVQJJNAAL+s7FSWpP7eIGqhh2Za7M4ZBb2NBvqzgo0v22fApi
QEbwdu2ukVi+2SEjCtNCae0bt6PEMxa/+52iCpC0fjd2IrdRPMvtCSG2OJ1omu9h
SiOwuF3Lg4fAkq1nc6o4YcQCCmFFOb25XTkNVH/AViJlLkmfxXKRgo1Rc+uOBRfw
ONZxi+EkJjvGnwnTVx4unVQ5phCSk+smSqhRAKWg0hxdaRiwA4vNor1KgnLmbcEm
n0qziCJw6+ita5FLP/st0eRzXcBQiRbFKM3fT99Ojt7isr0w3IPyGqCm1JX2Fo/T
Lo+CATpigascWyo5Uf8J97bfLg2wqUmk7hzaL8fTEETdhtBw0jsPTVTL9mIIrdUS
/K8qO6FQj3Gj1tM/0BAuSEEa/cA66p7dfryBCtXJ17MchO/UtaLcu0JYA+L+SL47
G5jktZ2W8YziNjCzgaOtyQhPw0l09soehxa6nNVnjrwg8TPBrBNUW7arxVTxIYgJ
AEUmP2fTDok69Nt2VpHUszSnFJgG4tbW9YqyjrviEJOoQmaQXF2JfXTGLwEJxaZ7
etseJUqxF3L77YdKX62iuB4zEUhi4prqmmV8mgC56ehyMXM0L/71BIeQN6u80HWk
46r5Wo3LeUay3nPmQbIGVqa6Gr1RSJLpNhd8rEE+jQO61XoxOyVH4ez08LxOACaN
AG56jzmQSzbs3SQLKruTCG0yeNovLoZY00lli3eXWRzgHwW6rrE+uV4Bp7+NsGOt
oBlJrN8UGV1I4UJvyjfQhoWqaudmcofaatWKD3/REKVH/JjaZjQyjpmuXvvSKcwv
wOknUJGAA2AtsWkjC16mmKkKRDyw9g/57w3HMZWofuPsWg5SlFqdyVmyXYDwnLpa
9ToDK9b9VPViVDRfe7Gp9MhexWxxuTcWTV0cAVJzWsoy101V/Peck7pQPhsqyp0T
AtB/vIPQ112ucNim1LTpYNk3Za/6qdVSL6Ay6XGgbwGZnxQzy+AMNIRXHSJo0gW+
+SQfeTvLxfpb+AIjHzxdmyjIm75QcpBz9nz5qxEoGetJt1BIb50fnLMzop2pOvKK
X6oljdCInwQUHoH8PjIwN4elTIjZndRa3XOi64lxQZLG3sDyu1UmQpWV9FoNzNc0
hakSJXsTykAE1RsCTB7sm0PShAlwQvqdUeiENUuAh+bRFxPlqzg/+BCffvnlWsnO
3J3oB6p/02N5GMC3Ee1Y8mFpZ1HDqQLlE+1DBsenjvHN0pK/G/Q4Yi7S3Yv1vO5I
pCK1A+o7OrfI/LQGT92iiY4G/5i4cY37chJSSYUCrJ1IPfj3DtK2RUD+gdoGGHoV
PNYKp6Dzf5r9ERT9n/EHY0cvLe0d4bUddKvjrcyH/Yu9QI3V+tt4lhkI75PDrDOH
k5RhIO2Y6cpWqYQevZf6lU9Qoe4Y30SINPeaMsupxH1kqsi0k86mQ0qa6oRAVOrs
32ZAyFpcutYwZchqOd470TK9GSZIYpQWRFq7gGQBOMN9goY9wnaklEMGgTgeAPR/
Gvw62QGC5o9cenqdye2EbmE/xsMDgmDhxxHrmv3NovZVExHvoDUHJrk2HpZITWxQ
vJIUyHffgZ06cGKJTNJczqMdqmcafxpgo0LcZMQu/0OLM19ljCDkNGxNw6Hs/DPX
YMD9T9chpXSm7mAHGzVSgclM71MyqCRe5kHH3TVgSTSDCYNqME2VCodSyt8DAQCm
EaJWaAATuIK1u1iGT2G5XoxfivQzwcWgtvBJ+mt6R7qDBfzvHfbYrqyOHkGS6p8l
Zs7utt5lqHpAl0x2g1FfVlkIY2vX24Sw2VpDet86N7pI8IwMFOXFWNrUAF6Ci2+v
jOV5WMAICYSOBlPHwN/2//i9QZSwnph8x6dCtIIHrcY7tXkgoyJQZqholO1PhsIA
0LPteMKkSpIcXNpi8kIfvUpD0dIj8VfvKc8GWdA/DzW7Jt7S3Nh5vbh6uXTl9OD7
J8lgsAETFtnUa4w079PavrIhrx/gVnyOa1z5lfeDHy4Le+ibZNngB1iIUSTfZGvP
ngrwyxKtrnfuSRd0XyX9cdYa8Y3RWKE32pdfui7Koq0h4urUB01Jv81TuwOzJ/3b
G3AyuZ1xpRVUUHlPXSNwYO4a65VIV/BF+U5bDpOw+FQVvcMVE1X2c65zyuG9Pysp
crbslkYsMgJJpRw5gj/dNErc1H/Twp7VABzIO1DMoE99pErLCkTIEFLijHFbIyUd
UXNNGVsed9xrEbZ3uvFNkfn/Ce8ORegecIUdiuDICKcJx11jK9L5MgwBGzybk7ve
/zLmtpKfFogh9sXZRn7mh+j419baPYgS0bpz5Xf7JLOvl5yIkzexM6kxrTxkrGDc
bflp0knmB9xAcgnSM4xZCdGnlsPIF2ky8B/0PoTp6B+sY06SQWyCWb8SKrQxCQfL
aTiofbyPv37yYCG+cyjgv2EzVTN23QOVeT9xGognEONMAxXwmSNuiYftQby9NojT
IAbM2ATYcGjyumGfXCtx86OcOfe2q6lm6AQzj+/vIRNAaHE8fLR+qvjbQ6v12mx+
JwQHM0P4EY/EWyKPFVxN7Abh9wTkgmqKoe2GJRyugZRMCFCnMMrJMaW8iaGi9XVF
SyRGMeB8NSOB2xFnfEn/70UmZONmZxWVHlnW5s3grrRT+vQSQlEAgnkMahvsQMDX
ZjNy/TWkO9DBnh/YobRZsSmlgZS/p+fbrWZUbXLrUIw2vEruIwLCcczt9w014Bh7
9RfaQntA+i/3ut5x/Yb1nNQ5Ebh/KKS6M6RNmyw2OrHL6erC4cacxMVwxIKybE7I
DlUOfX5/6zvDdLa+t13EvOPENb1F+wWa8nV5iEMsSx1ylZi2MrjYUiNFL6ioOLWy
6hw+9iIBdKJU19aOq3C/K8Ma/NlszOh59qFd154l3RHpx8OAF7DSPx6gTNKosn5I
MgG0aUfwfbQ598qyFypwNxjRtZHE7tN7mF+g+GwQkF6dm6mNzk6b+qXnqgY8+4AF
WQY2i4H2N2QCHTGtCFwzEQjGn8sxHTjvCvhpg7NCMrDMtJ0++kiRJQ+vZm8EE0Hp
Q0NPLbMHhTZne30878rSLx1ngCJFtQhpxFDA3tha//b/gRui3y5T3FRjA2QK5P/K
PyIum1xSvEeRd1j3bm+o7G1ddLtG4PcSmEvgMXHe489P0LOZfBCXn0yg7a55MIkf
IO/KSzvviTWBbBh+XRZGwu6Y585UQ3cwZbiRqVAqmgQW7vtw8douovxQbeLf15Xv
LitVOpQ0QhLA46unYMUKXald0Bye6Fezel+npb7V0RbUlYBN58wRomxbk/HJOJrD
/AuEqhjOIrfBrbP9Mk703pBa3+iPfuqsne5ip2sKrJxpRJT97ULd5/w2XI38Iu4i
1m2Ae8r5mpSW/XmT0wXK8fF37vUlyIpovNb7uWZ5zI2OHbmm3LydVKf+Qi+nGBfq
FR0SJ/v1tQMYbiv7mbytbx5M3vKwtZyMr7UChSB8yX4EacrrAbsp2nHJbYzsLdzU
Tfu9b3gMBIEaWLICXWB5S7fL+QuUDmQfg4Te6UUewIFfaJ+jW40T2EouJ+Y/9TwG
qfn+7vTNJlOoLXJP21xIg7975G/Fe+W8P0loreVuZkA0xUn6ulPVUrSu0QOBW97x
hDrYihBhDDJ0+L/0uHgfaq/j2XFbYK8pBbuCwvOdeKgH9NCY1xddw71XVVD4kWxo
FRGAM5yrPqqypoa3xCp6nmBbrNwlXeAMYZwSeVkQBkonQ+6bZfbijOW2ZKklRsl5
0yROFy4gyCw66GMWlg4so+T6weakRFEG1wYApIP9p4rvq45zUUt+Kul1eVD7qZv1
Z6mhgTnJ4W7/Dl/AT/JOqvxsbMALyMksPc0C4npD1SVi9Y0JbdLWhvr2CE1AGN6T
DFD3y0SponXR1+zK+OQ7uDJpoq1PZ+VT9TNQkb0kdoZpmRRV8WxgreFOITZxmdlB
j/8qixE8mEtI3yIfhma6jEou4AeFoObV3InnHkIfjBvcZhNAeANnnYeCEKzRRi3w
1w6QiL3Ef7DzZ3rsenbPJ5HBBXkcSoBmATQmzaJh8F25I1BknXoMwDvCLWzxO7fk
UIok77JXyx7xOlCXQpYJtaGOllrnStR4/NCeqGr1mesydin9tnJ9pOQW2F0YAip2
jvxl/2ctqn/1Cx+HsqB1ZRSW3Tora0k68648cL6bfK9JVHRZk9WiCVml7wYsOW+5
T40eohXgQ2zLv7SAqTGqhKA5+wyzVbJvm/pON59+c8v/odlw0NJ1A+hM5ahCQPOG
Q4b6yLjp2qSojBNofnXCK3ES7n0ABpyWIhm+kXC8f729+bB60XwUG4QvVu7G7EHj
wGjFNPwztCkfTAEG20yLZCTzfBCmngi19VpuJvDNZLGocdwvtACl7mQjl/jHn0Dh
TeqGy4Q3JmavzLVQ3VuolJNeP/AqEs3yoGv4Uh6r/WBPr8J0CS/PKNy+NpDdvB9W
Mys7kXeuyJWUVpGsk2/iuOeBSigi/HJB9vluri01NYU1r8SXxikP0pigj+g5Ramv
sxpzsVaETB8Y0t7nM6pPRO/3JpP1fwICM9r6jtby4AbmmZX0H/oXe2a7qnpVhlR+
1P73puTb8q5Mb+lQslIFMfH27kEflKe/471SBuW04gcL1xlpKW81dQYa+pSl2fnV
3uGCnnGc7mxRkA6a/nqsmfkn8d7rLMZZgbBN2PsHmJVAXROrqa0jHJmgeGTfHbi+
AewYzv93G5jzNRf7MlWfa+lU42COb4DjPolp1qhbhWsByLR0evB8RgcFAfjv9fhQ
hZtsSI9vjfqXe2mJ0HVcmO7N5KJ0/FoT7JlyymD1isTvplQoupaFapIWzJp+4Slz
tGyKJRY0rwuiTYW5pS4H5z8fLQZMgOvQCBfSQjvYywQ1nQa2/ky7TDNWe3fn7Cb3
vQdH2fW8OQ1zL5annzMvO6ymb2le50VWB7rLn/qljVohfq0ihKSEx5Sz/gkWcw6v
A2ArEdPiYyOqY3hPuGdpzRaVIIeacCkWCy4cFdgCaEqfyBpVLEFXuOPCVTtcB5x9
waUL5eCL/eCQN+xybrnE1JCbdYb09q/WvUtpjaeLxejniqNDY3HtardPxoTM8E2D
lxefR7Nlg/E97oVcR9Be2DYomFSuUjS93yA5ReD3wJFsXeL6X9VTrqLwIhJOx7jU
QoAhfAW4LWfAQCqpMhTruvRDz/Ww8tlUsvWLoWk52dZLvsEkKom/W83Ol9kHjgLZ
TxHk40SsE0oQuXuX/54XAMZIJbhij2lhSFwNO9n55/ZYgUynjZZoigxuSLcJmtJg
4C2KTWRKXS95sFCF0cPkyzr+piJS3dd9QIaBTYC64C76l5DP3Nd3cgu1DoYB6B/g
F46fwqQ/+C5N5gn6yYIG0srl3ri4h0+a1MCPnnM+AkyWNtapKwREw+btL7iLHpoU
HRqKrxUEwHdj5VXEM+DJkW96S3VSuC8DOlE137gv45jwaJT4w8Dp5neHdeYC9uBF
7a8jESvnfBKiJwMO3qJiRfdSQ7PDzMGVaRKzcl/u8heix9vhPA+131HQgvbNnV0q
xHZdymIR02orcs+MjIq/Q1RSA7phjcnWKcquCc6+ei9wGoMcY3mdZcedASOCdvp3
CKoTNejw1YgFK5iSHTA2DdgJMeB0oWxKQJ8l7Wup9TWn6wul61xLbIif9yAFnKXW
M3sIw0uw5UtTa2XHZ5ykwaqke7YfT/vyomsqxk3OWs2VHDUm9NfLpjP8H0m5uaUH
1tJ7jqPywdSzbfMJiSyFaunuAID/RPRGI5v2ggzQbx2UVrO+rRCk1mG2gQq2bn/2
diqlABmjCagUbpwXmiLArn73XMJnEqq13wECMUDFiaGEDlYCkzSQzesXaJpeMHMb
AdU1xOUuaIFaVEb8F15OtOrrLupkYlHu2mDI2yZkwDXTdQCQZCEK9jdPAQSpwQ8E
xFz+stOyp3C9rn5RyBOXSElWFdwRVhEcpF0q8o8WGaSe26LKvc8B4h4spPhdgwbZ
aOlQyBC+mFnDfH/dsj7jUKa9rsLI0dRcMvsAkHFLcLJfsmdZJ+NLBA3gBXAxscyH
5AYspMxswCfZ2iPVHlXeB/UHGEWnD0K9pEVWCc37do5trg/ndfdSMXpQgssrVadl
ew/hPwTRjTNZCwk1+VEZMcXtsrL3Zh8huBZPoyckI2rX2ZnBl6Lc4aswrXJwJvbc
o8sB+ySLvzffEcxOo/Zu/Njf5TEcbaw3PfBTC4Kl90Ol6ZY0gPhgx//zM+NU1edE
1VSgClb4d/NhVVmRiAFmc5ukCQZfyc+eDAQq+uKwE40i7pyip+QpZNVTiKkgMbq9
A09HTZ/FSgPeFOSPtY5gSKYKtouE0ohDtm/qi0XBj6OYDdrp/CDD9HriqMGOUS/K
+c/hLgvZrcqs7RSDHYy94x/vTJNPFzX94XQYIoi+WITkrYyBH8ky+c2yQW22aGyC
3lOu99dl512Rx1XP2cJRDKKe7qu3OIol/U+ktaMbFbk72P0rmiu4yoXkgJyRRH1x
bvi4N37gYhZ1eH2wL507r/S3Ytker7zhswk66ar+dP3S5Pkd2T+BH8oE9XF69gRx
4z+Hnvy4TyfrmxAlQWgd+HyNKYWWRXI036YPnCywASMjld+KL58c/y7jUewdFOv2
0S8ULKWrl44SmSv6xEkHHL9FQL68ZGVYQztSc5ToYGVEZvidfo/bTkJIL8xsFRfc
NnMucXCoorlS40NBD0GeVMHhwS59ECbj0OIqAagUyg20773Pb9Hr2qPeymWT9cKR
K/CJXlYYe+AnaJWfsrywbkez93iiR/JqoALo0HGYfEhzwZSHQlu2yGobJu/bSiDq
uCsyHcilPnpRR2j7aKvCFO0al9GZzpA4TmN92tcySSYcJvWld0LWP0g01rq4ZLCF
yZsoByihey4Y8huhR07rZdZOu8CGuqu7PINabpMv+LftLcHAfmmYiZQSZwzlvE56
ymoik65Vx7FwBjAh5UhpJsaOxpV2xGKgSGMjlYS0e25EiJieLHcikPsjlrGGo/TI
6NyOE935Xaink/4V2xQHg0jLHEE3PQ79TNl9u+Z1TogvodQWmwE8bcSjVR08/KQN
gjXqdQSutlBRdr3WoER5BRgtMJTDDWM5e3VYzfP2sl6taewiO7okqbfJi0nDsBDs
Vyy3udnN2oBKd/EwP0ppG9/5Emof80hBewlMejaQbgQUuShypfUKjyAzykVDEqmu
cYrPkjl0HZGHqvCGTj7yeCNZA8E+Q4KCjRUzkyyHwvNOcOa8EZi/CF7FNOLC7XE1
CB5lG+9xWDwEi9rPrYGDBI7NtUtZq1tqrFTjdMwl1eR++eI/c5PBunRVZDAAr///
KuXZHgrX40EM+Z8HDLknZcwdMjIiOac6boKqQFHFcqsW/ebwSHyddZk4hulWzJBa
3et59Mc5WiSL/1Urir/CLNFYO0qiFoeVLBkp51ufUorLow7cYztno6Hq+hkHYE8L
lWxXQ2EROpShc6F9OifQRCUM4T7tzmU5FBFoHQM77hKZVX0VHtZvbhvImMFRZySY
2RaQqK22MwtNeiKOUwy8xJtThoQ7XoVGFNtzrc80xCIwEKDhRVjnOTVJKMG7VgQy
sQXokn/dsla9S+uLwpkGQCmg9DSEUVM/muI7HzS00kQG66EigTuQ4QU7GtdsdOKq
U9Q4eb+eqY3V4CLkVFwiDusIAbaxpuW8iycpui5TQitXNd38apGSgTFxb5YCAlDy
aZBDccsnu3zBmGg1AtmsE41//iUjwBTSXqrqCj27LbGSgRsdLn2+4wXAGHlkwiad
7RN1Z1nVS32V0EqD4WymK1Sc5LkgT4f10TgoxFEL6dS0LzXQ/lwvaPjligj4lVGP
Bkd3szX8+SUDagK/4v0oRecFs6nkzu9P9zUIvquzC6LnujhRI/t+pgAcPerFtRbx
UYxWYHkMogtXcgMg4CMujlbJAEzpUH1ktMH5UHAn0Sfh48V+6RFETE6pDbSNHlaD
nyu3j2JoSu1jI+QmEQ/NUqoOdVHMvE5Tz8u7/zrfjiXQ3Qm/DvMzziN0zKpQ3kxL
JjRYIsAr5DTS/8g7QXn9froKGmFFtaC1APp70qK1uzGdWgO2X9/69o68YAwScSVV
GPx1kqYVv5DhdKeUe3dCH5AthJKJpuM0/C5prMDZdwwb1/zlcohhb6dhMwHPVWC9
if+b2xMgRc/w5jwv1UVs+hAdCxpWD++1ru9Q7m+yeKhDvMit1EhqxI+y/cSG9Pp+
tMWHoCmj7TZdoFZcGEsVtCD8AWSK5YZwlpPodD11euvN3BKRNotxGyQbbYtFzQVD
CFHLmOXvVcJEX1yBBp8eh1RYRhVphi/pYODMWV7E3oRVzgn611vMO743OjRFkulv
uSwPAVPQgQrfbLC1lDpW1MyA2xIC1EvJZ2OKI7QIFp4xP8K8vO+62RSj4p8E/wV9
Cv0VbnGlUhRuedpAn3+L6UL49tYnEb0QtMCFvpuH/OubPSVNQkE4OXVnrNdjikB2
aKxt/qtOiWMikQYVsCMRoThFr7Mz8h0dkpUFhx12uxhMjZMV7GZNjcEbG2yhTwby
TbAAAeCjVcF+wy2oFAWkExQYa9rf6i3vI0fpDT8j3/5VHXJhyaoM2wrykzd+HvTl
ttpBbXTnBFpxmxpFUdBTDZkqOeJlnbDfQxVc80AUX3BuZ4eY3wtJKw5dFx8bWYc2
gJ9TNZ1PeqLVHc+oxvvNsEVsDnGnLb3d1BxDu/QJAsYSCJh1JHz1fTUqENFOAHjn
+xvTJWGhIx5wleimG7YK5zSyIvsJA1sCGonTVA9pIbXgQP9eeQ92CJ4j53CV0qnp
JknMowD8svdbefm0jen3gsFhszrbqmJHSiKkqsOhWk1p4utJALg0Ky7/C+9oHI+W
KHbIGsBevFXzxxQYHZwqhVmmdQFUinlkxYg6BbIRupms5UgaBGEwpqTBoMw/qdTm
KHSjCOyiPouLatLpsjxm+DyG36fctMxdLvg1ESQJmxJbokNoAhMT5TaCCCR8IDyo
UJ2dGzQbI0mo+dVSRA4yldiGhGne9JpqWDxL6CUdmu7qTB0xxFZGAZV4QWv9MsAe
DspFny+OeV59J1NFlRILuN+sOanuKLVVEdwuI31BV9O+qHLHRDJ7VTGl4GrCCtOH
aGwnpNGUU8dVD88OmthXlPYcZQI7mrwmxLe0biwBzvXGavnALZR6xmd5CwpbEUau
YIQ7604K7Ac+Q6JL7Fgww3mggdzjQGoRrpa2imNgJNUw372K5ZnmLSCe3bCvFGfN
ETPT0QAZW0u6OlP5sseW0D/lM9zGFlpMeGJOcRDGdoNnNaXe6GWRzxGpc557C/tk
Xb1kH3HOJne3N7mJvC0smk5B3uV/mVthBSZSsheVuw7nXyzfj0yzPnd4i4e8DDlE
5R251XiChy8gXncFcDPGLEQjK5u9nEZz7pC7pEWEYOEXy3U2AryiVrFUEL0By3/u
iC1s5ZqEUM0xttXg+A+B7IRrKefBSeDWtT+tvpMVs5nH2aw0iVxl0UitGvFwiZ7+
nYYFcSgZFsXjONJRWxieXoyoc5txbpcf/+I1HaJ5lqktUgb5cYgt6WpnuEFKwPSO
VSfA0QZHh6S5AZhZTrM19LFCqAUZCJCMfb5UVj0Kapme7zibCvI1sNt/J0Qf9sHB
YOCkui+TJn+Gb3Qmkj4QOelIxTRgUzZ8M73Wggo5Qg2cicHTf8r+nvlbV5h1j6kQ
ZaFKKj7Yr1mtbrNldSl4uHoalA7Na2kumMdRCtI8gh6QD6PvZA6cHTmjesdUM+1u
3GmpNYl4/bVQ6CPcDGRvjByEWxAnp4CQp3z/T5lGylh5VekTCo5U2H5PUVBPEUhj
DGH2kg+ZPW+FPenTWBKxdd7OfgkgK+92JXioAkE4n87Cvt2fJMU7FMPAbwAvJTVC
ZQHm4vNCJTXwMqL7vzOvW8P0Gu/aRvOkFZj5AvxZUewFZkjIyHyiX915t0sdWoeU
8kkLlnUbAxGl6GRIeEWillhSTeweSRsXMM0bdNT5naRbnwoBQgHo91JNC4/XOuV+
DCbpF0tOLP2wIZWA6AuEZ+nEe6XCAQVvdMUPOGPpHgN+YrANFTM5dedtLr1asLvi
kGpx9eZzhOKkT32g5sLsSoJoQLhSk3GgnR9fhN/tpnpymRdCNhXTHunpwh1r0W1i
lvPkM6Y32ihNWTeWme/T+GMGdrIoDSD4GwWe1Ow7/21jr5aTJsAsRg3TNt7faTso
Tbe8XkmPcwYMguwGkbVpesZ27KUTKVhslf87e8G4Do5vzLkS0SwmuI7gztUE6IM8
9JOroaBvG7Oj+wK1Pkp0m/w1BC6CIWz3Ge4eKZcU6tzvjHHgayvzhLqeXZ25imPS
Jz+vvGLN8Y3tgwV6vx9brf8fVt2dThR1jsKNWK5ffInE/6lm2USsfPlFm53CvLj6
LEI1oMiSUm5qffSsYCQbagLs+TdtG8LyDuDerlcvIoFrFfbs4cm9p0E5rjEfi77o
QfXBEWRASNp5rJV/0/G9hGotQmLXZdh0VnjIpcvu10XK6PC9xn44umEAvx8Hm8TX
cACY+6D19SpoZUrjz7Y0I/jYxgUi4q4443mzus1efBiDk5R/jWtciEtC6aYSJILi
sk7ubSj54WaF48EoYYgpuOztindNQDibUDNG7eIQgYQHctGOhqjhK79A0eONFfA7
rY0yxOI3/9zOfj/9i5geUNzeExQUxLDtYV8UVrd5RyLUEE4IfGM0jppFtqEAFIs8
GPDCe+9bYUI2xkrPEfRl5FcWCg7RO/Q313sEAjKd9HhS8YK1XVIsDdyBfO17Ln1V
TCaEFXipn/JIyX/P5CO+u3d129XRwOvErgBuQwtu1FCi5lZqFpOMddEwliKbcEBT
EgiAsEO3AvUSKO0tsz2rW139hbucvYR+U/7iIhyLE+aZZY2dvngUq27fQB8FKXBM
GsqdZPxd5K864h3WqOc/KBr85+gIWV0V4uxefJoQKvSpBHcAafuiYSYdOqVh0683
SxWkU7wPlmfQZ6SedceBulEs9tlcwfxiQLvAoIz31oLisJMj9Kfn8c4DWetnq1dc
hgp9gbiN0GvJT3A3BByLNcsmjqJaw75hMejfPUmoEIOyHfiyE/gLoL/XBNZCPWNH
pVFkMueZbDU70bublwUoGw4bpL/eGnxgvbVHn8oOJMXsZyHEtkLXyCUMvK2Tktbu
9r6kf7/D26Pb0CTQqJpwAMJ5Xz6Dw9h6lCXdfWmSiCXjJSGLcOHZDmMOZ/B0Grz8
CZq/D2rImUng0ol0voCZV2+Nc5q3oFGwBmYJn3m/VFAFrSwe2qPDM8Pv5X+N/h1f
N6Y+A7IGDqRP7yCxfZ11fIYiSE5ElaO2r9NECeFdEQUBZ7zRQKLFhRGwN/USiis8
DEs0Pd8iwCkjpnKlHKMIbvWzGEl69JCx9lW3LvIn+59i6nsZ7sWimem+DZuDdQ1X
NHOmm0yt2b0mnEIIn8KewwlhuHU+JhXzDagAMlq/6aZd9eX5ZjMwGGma3j4j7OiP
nMsmeJQS8eyXMKKUmGvtuUwmfOdTdDC75ABXDQrGIvtr+jcOlKEXdRivIb1Kwpek
tPytlWPC9blz0SsB28ASY4KucxmZdeEjR9IDuXuGb0zt4FoTcPpLaEKXEq9UgGlz
Fl/Viu2fxW7fJN4ar4CNi0WTzKBfLX/IOEsYOmipQTDPgHEVqUryw5AHNpJiKgOj
uYY1b2RYP6DFcZPboI/YEWuPJHla7ryCt26LD0bd/zip6N2RE7Ih3Oh+/6ii2cf+
9h5ghuzg90i4KtzH04gxiFhrw9itoypT8189oZCZXdnjpzErdIcjUubXXfkxCZox
azRu8T/HzSOmSz0dGP9ORZnyfZmSPy3GLtybFMzlSrogXcB//E+m7tludtG7QOLi
4YUFPBdXsAzO4O5huvYuSV6hRQYy3us99TsRIeUlyMeJffnEa/iAETxKFE5B/1vK
qcUD3s79TdxcoHmwGOGavpf05xm22Nur1wxefavVz7tGriUI275Su1Xlael8vxMT
kKaCdFpjwGTl7hH3lSbjSTdBWnbCJjjmrgLCN5Ra4P2wq2f4Abpc1vHWOG2p3k0l
YprgM0NmGSkTf0T/VntXhOzZKegrnF3eR64TFhYqWcxig7A1KOSMcuswFaHHIVHz
pepX6vWzzTezGUJHylTmvIWhXTaM2JT90fd9KtUuMPbwV28HFRwVGqYM8DL8sSGK
kt4NB6WG4/2nK7r3S644hiZ+QjUYS+JzJKMuQXzffQmY7Djj1xJ/Gk51ArwpWGi7
dNVE7KHA5nCk5XehrkbWasqxiKT9KZ1+B2yt7LJphDH/fIgDvDiuMViZjoIUhJ62
ee8/PyTg1SUR53v2Il0nHlsm5jxcfgVMxSSSZUxikB4B0sovxV5GMC+P94bYGovV
zUhyrXPliDQCHyalP8sKwhiS4quFcYgn0dzIeVAvHFdXSdfDIZrnqcyXjvQs72b+
RGp6Bot6V7MvjkwvHsVwlDYZgvfsl9hBz4wO58Wav7czHiFiH/tP2CMbU0CIcWKg
sxTEI4SoGBOC7VAaSNkxZ2ewK9rdIxKzEfivWEX4iSEOQhmOd/IHO7jX0HcrQkmV
XLB0QOQ9tsfvpOB37vEM4C2WBRGsuL4PZn8p0wULBsHGZglEze/frQfM8KfKFIet
UO6XjgV7DnRkLqcvePufreAVoDSJXZcEOTCR3yZUUzbLcaPmY9V3pCuyJzHt4Qg5
4fjY/cRPqZeBR+PTy/3AWn7a5Q4VAsVS4guFdENUI8GDCKeMd9g8Bn+ccuwNNzJ4
ErRKAMsSPs8lXmMNONmQfOu8cpSq/mnoM8SlvRcfuMOknxEbbTt5qW48Z/tp4JLL
g7nruZgmBhb6/Wcl2NCOXsYOtUnuQppd7DHUc6AXE5/TuQe2/j0hNXL3Ln8C65k6
7eaJzR5/46Jl/sO4RRivz78PZgo7RquUH14ZHqwDjJG0HbslZJ/lPXFgvEkBz2EF
80kxbUrIB8mBDiVYhLdf7Eq4s8Cf828p/PjkN6pVLgntlM4EFBVCVVWydMqB2BDJ
fBUe16AC+0yr2Ulpr2hZtk3D+lzYl9LeSwUADh4R8ovfOGXshoz7bvZ2JyIgP7Du
rGGg6YRbfifWcDj6+drZigr0sNrb2Z1qsR1tdEq9YYJFDVVUAvifNlrRLxZrQsI4
FkrLTbZuEOWiqngbBRfbu4q4Afd/szCF6c/cyPHWa81TDjVbKznbqJDOxUdAny6u
s7b/veJzjRSGeKhRq2pY3UC708LKn9q25CkQVxg16pH1vzlKoUu4U4qlEq6O0HsF
I34nlF1uwD/ADpZS9AFsmGckUSvRIhvsJ6eRO9JaCqjTUC3qejpVgpVdnQ/h50iK
U0KmAretwL3iY/80LiAeLnQBoqT34Sg6BIo6+iSLOMEJSOA2rQN1DGxgiFT8CWJ0
79Fmr0/I2Hx/PKh9t3LXRq9uzu586Fm0EfA+B2e2FXM/EoJbsv8GpYE7gVnfaoVX
tUvOw7FEUxiJdnUPLLDHPdSsq/38fzYD5O4L7DtOat3ErIKArjyhzY/I3YNjuss7
nUYH0REZzOUpzFeoEIJ2u2lsRH0EmpvWAVMXjhaZ+LAr8LLvDwLRxIEYpDEaL4TJ
yglnMkUXqoR4t8YZ0ZnodWfVUrsz7kVsUsz6BBl/J0IZalVD6P2FGiBnmRvG4tOI
nacR3CACFSog9g+9buOuD4cQh9mCgttBXnddEvz08Zto4UxK0qQmn3pxiQDg5WGf
HhAxh4AMBUxjPnKBbpsSFZ93XXmkvFPONKOX5EMfQUsZdzUH+zWaLrdGsD6xYDxM
B7hjHb7ekfZRTybvQoiaeDwrw+GOKvT2k6Zu6ZgbA4Q5J1q8Sl/0hmLOMX88ZsRX
8U1cKtV9Ki0qGfzL5DGAWrYjru+Y5K4SOsan9H8Isk0lB+Yk0K2RyCMhFrc+j8KP
g0EWD+QnHpD5TtXuFtrpoUEYjqEKPWAMzehO/vBarlmlPrdQjgT2SLW8Hg3lFW/t
AwnGMzuml4d2dYyMwUvPuKX/SIs6Clk7bBqZAPkb2Mghy5oxC+sfakD2yy0hNjCS
z9Y2eNu/E61u35kufr769MrNobPJQPY0il7iOn0XP50vLMn0kcrsvitZkKxP+ftL
6NTBvXmbzKpCPBcWKwTHz9LnXrjNnPaHZsNZpj4VEucl65NgWLHYKT/PejNRpozj
HYeRwpOeD+cCp10mrypeym39LbT2Kzm0zYXtSBVRZCVssLj3NVl5i9Zs4Kycluwm
I8C2rx6xJe0W9BQaRllWE+epOT9z8eWsNuJZ2/V/PFe+/+sXluBrO3s06UhsxUY8
He7/JqwTEtHkpWmEl2Mh60NZf7AEaj9C6KRgnaEB6MBPKe0ZXPE3gTAqTlz7PBml
3ZZV2JEBbp64f0b4AKlIjzKVabzg+IvL1RhqYd4d0sIeQzuDsgPYt6uRYbF+pigI
9PHZXCOB5glXzqGf8F1RzQk1uloSe+HwXc6gGzh0UgvB5ylU81YYsX8YZJ5TcLZr
V7RVv+JPkjpLHOAK9kxGlmiq7ZkHp1rzfLEngNC3JOyfMr5A3OM31USYsy9vA/ZS
+aBr+eZkvGwb+O1SOW02fpR19k8ajGYXmdU2k4SNM5+p/iHQSFAwtSgArml5y7xB
vGfmEJMeJ6jscfxm2QXPxLEjJHRRPKeFGku6JoTId1KT5/HbLynTlJCSr28vYWcg
jCvqpzy3XorFMFlRh7162ceKuv50BkOFibs2nKAvqL0LwOZrq5xVgRumtqEPN+xO
0+PbTrHHLBFS3JcFRbjxAz7IEapzqa5mYbCSP8Uuf/vQmELAR7C2U2PM8IoH5heN
ZZb5sNk9msl0SS5ZOUq7avyV9NCJV5WijlbDAdZlGzBYRpw/bMIF0MO6FraW82H7
zIQNsEwU7is0NUhDqozRZIN8dfTNsAuTCZBOln3mD03tU4qmfGrE+g+n1H6HKYZV
CLm81Qk2WEMu4WG0JawhM5smRW6NXBmWnR7q24wSdkjFLNmhzNhOrQbQdRqGvYyH
t/lLptDQABYOd1FaMJif9o2SoswpiXbK6QDjxVRR7qxT/0qQqNBa/I5pP2LMSDVI
1w2ab4lVIEDGwEBcY7WPNy7w3nv77nMgB+EqcZ5E3Rxa1EkR666qLpjz3X84t/IW
WECoEpycup06GT9qcZdGZ5T9B8CEpyjsLvqqDio/CiMekx8UiVW+8ih2F1PeHYms
La7WS4p/hi2iGPvI639vlERTIiuARW81m5PXI+JYuAFVbF48eEKytgNlE2tZcuLo
fEbqeZh5lIrN3nQ7mAUSzym4TTi3SoThhpVn5LvGyclo2KzHFzAWcTOwwSw8mGWh
Yss21plx9EUyVA5ZAWQAAAeINmP4EQNL1ou8s2GcMsKnU60uebP+9UxEenehiQrw
36sRGQTr7IUDEJgJK9IFREnO3OwMqCNkMkqX6B3TfhyBKZTRlkQ5ru6MFNo2yo4x
hQC8z8eM0CLzEBrE+TXlSYmK5jUq4ZdNd9WxwuGIUwU4dpy7brwEbIk1O7AryvqT
PXxoYv9ZwwsA09VH1paocxQ8QySiZN8w7kmr0VOx5pfEABFtTZpy3f+suL65tK39
fT3D5LfPeiTN3JTo2cyaZ2gC6HIsb4aDAQj7astKMDzS0RsTNKo1Yif9DL+QdrI4
NkpTWfrzMFGQg0Rk1WSt+l+O721EH4uZqhTFeDR7WAHkFs3aGAX5KdBHJnLBqoZo
NUOGp12IZsT2EYGGe0R31Dy7V8Ux4BXLbNIxQ8VR1ryaaIWDBEZKmg0kzUv3ARbV
sTQFDxUfMHmxtQl1+7H/T4pLWWy/pU1lmFOTMqELA5hC6M/hWdwO5fdYbHyURbh8
durW2nQZp4oCEBcSn10tHLag6jxZgZX1qAWr3lFKnz2uHQYw78ffBzfQUUra6wYs
Cf7XFTbr45S0qUxFXVydKWSP2YW7NrnxltEujf5RYwbgCd9J+KwU8t+YA+u3NRpp
o5fgrqAKViTKehOrZlsXbah0EtoQ66XTYSL5GULHknmzfFO29vzBcjJQaEgXNrgA
4A/UahilOJ1s2NJNy9MLqH1L9NSqGmomleQRPFaIhdkceY5X4I2mwyxTYGBHDxb2
7Wrx/jjhsZg77g4YqhMXW6MMh5/WAoCl0c/h2XEsQik6GyjM5an8bsHm0K9+FIkb
qSicCuo6U8DfVl6rIQCeIXgquLeYKriybkVd/VabXz+z33wfAiOeMCsUlC6la4XN
antCZ1LsbNT5GAGoIgWSE/yj9De/2XRdNBHHKVodNsw3YIklbSW0l2DY9kYmgxMH
iGL5feVJ+yTKLb+gNPRZUB6qYLNtzq6H2x3O0E2TguE61L5fUr0gXECtOS/u8Tqe
HRAjgXgV3EaWfD9s+5NbfkAPtyDasCSS0G4/a3snG34RSzotyNS184A+upPhRgQK
bzeYTLSfkwJKp1HSnleF8y+eL7zdZdIwoKdfL2xTdgdWFRCARgLZnUHRKynwMqPH
A23JmpNaodT2g5ZWDooU1Mj5idHjKm+oNkTXKixnjKlNllNBR//sTVPCjK+b3KSo
uGLJkgrTzhau3TER+CYDgfszVz2gM3bgb8KDDywCDbJ9pvkhZdx2ivXE3AbZnFcA
wo1A21Ae73Dv8+HeLaK6C1D0bcPQpLeONx6YHA7kfHPsDSniq7WShROjk8Qgry8t
4pqyVgK91vBp5TlOy8QflOPQfcZURaEk6vQPnNOUE8eYrMrOCAwEK/CBRhsX0P+9
9LJajASkrNeVqnwT0WutpXd+ztcWZRUQaF+6LXa6QOV0lIczg1M6+CCMTzS2EWmV
BU036RGZddd+5niyfA5yzyjjLO29zyeaMd2sT1hMku8tNaPMtuRdIu0GF6WfThAG
7n/6ixnZ+oMGCgAPCLM5251SWnpDCZcYYQE+zvioQ5bjkv9NLU8pTgnD43TuZ0b5
R7qN+fQ+uvuIhkmz93KvBly2C4oOE7GZ/+aAlAxiUAk72K71ZeSdhd35y6at8ztk
3P7N9exm3AW1neu1mJxbIheyA6J5qeiq0tL0out9tW8eDGWSqaw66DHnqBm2ikwt
YsEJrOZo3kXL84ppQJcIEfqkTCL6jJx11S3ESsxMMfKP+mC6QJcY2jOAw+8ZlU6O
Vsfp0qFPgGpqjKElWq7eTOJFMPIBLbRPBUdd0LtX7YkCeg+v/eFQeg6M1kgu1mI9
uspDXh2pImhGeJRd9TBTjH21796N2sJMUKYD5tjG8em+g96/bGyBLB/Z3Lbn524G
qIV3rmrdAK9IWa/sBJnQTvM61xo0aDQnJdWMM39aiGQFumBem8Epgw0OtHUm0ySx
3OqyLGMlUMd0NduVEpKfAdG5KnxXltk6qpsbi1lVBLRD+nxynfPj6MLoPBSrqj1I
X6cK//W/v/EOxjcBYO+vpWia/7Yma+kPBBAvCuKGEcD4jqKtZxbMSKhHSqpmLAf3
GkVEcBbmbmZJn41cnk5cRSBNppXjw+l0o7+kTVOhP9FbYFTTs9E3lMMghg4UeJPR
k8ma/oDU5dgzsRVvX3XcHE7MMWgT86+GvpVdX+DP1jEv+SP0huEfa7p/VzSp3cHV
9ffbp6OdFJ0olcSVOFCT7j6cS7qv911ciNS24HsMp0uLc+iKeAP9ZgVT6ha5/5b7
u1jqOyMxVMnQ66By8Pm5Y0/HncHyry5i5/M+m6iM/RJHin3varIB+hEeCLmtmI9B
hG4gsEpLBFms5hvqzPkPP2QMkE9fGDIIXHyXInzS7WNoSqtHS0XtOUwGpfyO4cA7
RuDtfl+9yIY4MAmeSORhP5hxDPOkd0BBLPnGEf4N22uMC1QkvUWbd1zQJAwSAJxn
oMn2OysUE9exZCQ2yQzmmjZb+Vz/ErcTbtV3idcA4TQrClIRhxzvd5RuUgvhaiHK
AMZjzWI7QsXhtWp3hZ+/h9C5yLSutvybgs4/pPYF2qnF2W5WE1EpsPMLZYO0rVoj
CDYe72WiEUKHMv3Xkq18Fob6LPy1FJbCr/GShQuDgcSNzGXGYh7Ihgt98b5H2pWB
vDhA6zb15685CPoyD37CZL/x11oTWUOkiH6BQfcJD4LnjZTzUXUGTEnbGKOfW3JX
iXZxN9wRsr3rhje/3Q1gh91j9s8wGV5B0sRhmq1SUKPdkxAxsB9uCRUEZwYufp7y
AYfe5nFpNDdUTJXEYCC198x0ren5HdZbEjeQEvkCQJ0hjX3cymK0Xbjf1ZuZ3n47
WN19uOMB4F27++/jvNkHY7Qg41nOgk1mQc/wKcdHyhcNYR0vht97IxpTaC3uB0RW
8lLvBwjxGyt086NhRS0Fo0+DmIYMm2eCawK9uIjp2BnnUuEIUKv7QPptKm9vYaex
iuxgwllVr0EXmid89vSHpxLyXZIq1fZdK59X6eR7GnYRp4xp4sa7Z75zjOfK0v9Y
1Cioll5vcgoqwOJ3IZUM3+A1Z0+CWlOwsqtA4NU1TNldoH/4WoFtM135/+6dz4qA
CrfTfp6OhGLqUgNSN8orSuqSBgJnY8P0qWM/m8tdJaWAfb0sQrCPPLWAAWp5ZVUt
xGbWaaA9W7xy0f7bzcQ7odwo/iYPBTFvOwSfpt+hg9r926HKDZfdhRW/n8HiTxlm
oyXZ18GQSsKSJDPGys1zMAXZVs+Rr3cZVYV3b4+nzKg880SNvLFolvX+sk4YOEQn
YLGKfxy3hWOwraI0Tjj8Dt9v9lYJmrJ1OwnOYGFJW9Te42suo0opOJRQShX7Nll/
hZRXfZ/yDXGPF06Iu70EzduxPUNWtYnMm+ByQrsF3axS67pN4JWsR+GdOS92wsIF
WlPjbsuETT7WfFJg1vlodAR22oZ1rBJvaroAfrYrDAMfOmURnvx11YO6OrCUu+mH
i91wUfLd70LQOJvSv4Sm8TLU3roP/x/hD7lb5RMA/rO5yAj2UorUg7zuwVhvCPCx
oBuK5Tvz6fFJA4JqZcSpJCSuUxT6MfjnfXhXcKOms6vvWqE7ZKtBzxjRoLzrbcYA
1Umtl/d/Zj5BFPCXP0s5LWUltDDHTDn0hFTM1KEG4C5Skxkar52PFUs/VgvQbY8d
LDPrPWoE3LgDWhs+VCCyzwPsLoT6MlvCeVsDbcXawgu0tPZxOxjmGr7nok3rfeEW
KsIQeocxGffU4vmduFKi/jZW6itnHA7/2lKZ5Gp4oOmbTvT6rVUo1IAClnuHC3yp
ATu0C/OuCPpKvyLYMVlviReriXhrpnBD9CsCv55x2FpBq+QTKmEUioxvUCXVvq/7
uH8X53OMMx9rvFZdU+YlVpPCuR46ryDoDNM8hVBeCDj8Le4AaY5DG8dvNMvtjWoZ
LpPn5CIiyUermU+OXq8gv7bsEfCweEs4HBaveRr8lyVr3XqzZHdHab5jk4Y07hoj
YfPKF0le6oSk+hsFKYJRiOGcGlGCnM1Vvagv5zwr9AGdMz6kWjSAea5ZvX8RWto/
px1jbePA6iWZ6egPSvkhQql3XT4eHej6+GMshfsdEg70WPCwR68gvyP8ZzICLLVH
Yf0tMBORBG8JR39o583Swk1dyDqakh1//Xx6OUEO1K95IsqP5SVjv6qMvZIuJYq1
qbqB59crNCm0PmN5PiA9xfvGfJJNPYE1h+bl8Of6hMazk3iyW+ax9/dmEtY8ikey
+Uzn0zNELujSez99Z6/2LK8EWCq6eiMJeWN1YrudAZO+uoaiDKPUgGlcOcoeTas9
6cDnzRsZdG0sk+VmmSqWwNYghYOCGmbEnfl4WQbZQhJvBuKV9oAmko07w79a1Jau
Q0BW/jMUIYrtYP3VU+F65Bh3o6ntR0p4kV9MoGkna1iiR3SCLqJLI7PuJgF0NUgv
llhaXyqJD1o9oxFiTtfxSqpTdvt8rWFf85vTyJtXKArfkpPiZ22Gdptzoc2Dk8ut
jA++P6dKQ93L8XauK3/6rg4HWzb6TKEjFyA3CHaSZiH6J2ejO0KcpcLnACRuJZz7
Av9wcI1SjDLVrPEOxCtUsBFwmFlij1FkMGL5xsxQRal5+p3zkV8RnJ5a3VKM+k2Q
yceksAnkmXIpwXZH5l7yEeSxL5QmwanEP323quOKh+lMeYKao0NYfiOhMVOJsBVs
1Yq7Ukli/jsKkMiFo6v8E3wpMrvgv5C8+afZeu+kEHXySUfo4xEn1cBtq+23nBzx
/Vsds0KA5nDmOhRrgR1j2T3G9H1V/0JnHD7kRyHS/kGfaePnVapTPdEqs7WQnxCs
vvcNfHfOyJDKsrMnvK7wAZhTB42iFrrdQJCeezC3if8EMCuqPR/nnnL5v8q7RNPu
DwFTEqYMx2j7g5JxDDMFipWhojUAENRdJPM0pmvNwPrGLKa9ruWltBMUGbWdG91o
i7wBcxMyy2YXT5NHy6MrwOxKVlqc4HSonPwjv0D+Fv5628aQgOlxYuVGMp1ZI+mx
m3nZcQOcCeSOiL+fUNaITURaDzfneas061El8lKQgyPDqiTEI+16PiE9hFEkP6V9
XUN++d8PhFaLluo8nOFKC3R3Vy8jZSvaaBA6U3ObJh+VLhED9K3pHfThM2NatbUc
pZK5n9GBplVTh9qzYQF+Ar9odq1o5sd+cAslR9pxM3JKkTt+8196MmcsC6Gf3t4L
DHG7Cv+/IUuLtN/upMomEGjTUEEWEhIU8qa9lYCgUhiRADzCXc3TJ0w8gbilwK1F
5bKO5OexRk2WhNMZbTyVXZ8SezzIYrmSXdvU5xOigWBsYhl0aZhXeFMb5NJj8s5w
l65JBEkvLg0OciW/hPsUd5vZpYQPR6han8W8HHBYl7nfpOVrok4T0GFd4myL4+Hw
2UJ5eZApNQAcEbi5/TIGZYlK/TekyA8QoZv5oJFEgkwSe7VWTaCqSf+BjrEpBgrQ
+FyfPjolKkbCTQAypBlGxuygLR8uVINxNXwZaFaWbz59Drk0ora79h60jyo4MNir
xAY6znRhDtwFzmdXkEB9fYhkMXG7V2HyAhr3tyDVdsrk4Ubv4HcGQH1O18dSYnIQ
lVAVPOkzRjk5HCBfa9rCFDhzIQgcpqLgertibpAnJ8rivczLT/VPmur57zPLZFyO
awQ4n6pZZn0JWMcaDUL9+z7pMyXqH8FXqdXRkfrxbbrTjHGvV1xAQHM2YVU7hSMY
YIwbbFDKlFK+/6g1/KX8K9/rErwyK0uyOjcAdZgFTtqCJlbt2oVi5Xz8GWeaydlW
d+vhbrUFO85/InwbcrM5/IFc+t7ZyVSZkhzZ1CquXicpoEvqdX+AAtfxjq0+Dv+2
UJLVAKbBYtW93QRryW90W8O5kIlSufdwBQEEgTWW8TC99I3nCbl+qsg25Z/+ocq/
Oajtyuw/dOvxrZ92xKzGLcBEjmprfr0OyHM2wmUO0YxdMzwaH7SyOifUNnuTbXnX
TUzEeoCQWDmqXICqxzKm8Fswo/TxfZHJLYhHuHZuHCKkPS3qo1CNMkrfmcQIJxfM
6zUmR1uDnW1dd5xpaYMRSi5Ytw91618c3tmdnQ9ebS5s7nSbKzKIdwk1P5y1pvZU
6FpuatVrBqgySKrCvtztCF6EMlmCHrFvYjJNtVNK1uoKBxWLgooN/kWSGYAWH3NN
eU6H5TeTN/DKgeqoDUzsRt11u10BFwU1wzF5o7nTOeXRpr5c8PZ9J7hvHK6F0nna
04NSncq1PWGru9lnz9VuaYcooOr3OVeJL5JYjGvSAk3DtjXI4uhQ9hjbhrEw+oHg
y9FgH7cvkO7dT0I5UaftwOkoFgzQ2enhogoEzqDYT0QgbFs9sIeRc7XlVE4sS02G
ooHe7QHo6Gwi6XyHQ1tO6V2/KfNqNCfm1UC2BkfCOnfgt737ebOeCduz4um0/bVU
gj3/pB3MMQaavQb5lpocjYNpjecxGosr3kB/T0v6hD5+x5w4XrZVCOd5h7RnUvGg
mE5HI+cVGtYWqKWJJwgZLpf1rfTcPWh+bglE6X9KQg4fpWqtjTpnBMyFDm2VQLY7
KjWupZH838AXFMjJBwIfD0igtUchpr7hWpMQDZcA/M035ObI1OLuKo6wY4YtPZhm
Zs264g2sLB0SPzXQ/1T4KrA/TngJhkFsdq7X0tKKT6pg2+xZNHSxG5Kd5+kG2fkp
7ptTG8wyU49b12LGtiXZKnRFbFa7Ne2Mi+n0OVrN6UuSo+HNc+X964XiSPvpiJDC
8ouvemFpZCOim3poMdJ6+KIFnmCqmLIxigVOosH9Fiz98PatgvZG8TghboRMbGTn
ko1MwnsuuCGlUEf9YXTjU5Yr3J8OxSx85uKdyDq4qMmFWsW5X4DKGway4elcIEJk
Didze3O4OCQ+9xeBsSVLq+a/OPkPPpb0HSRYjZeCiBZZU6RgARc3yv7O+Y4jt11R
LVs6dIkXqBzGOugd2m40sjf01T6V+7JLl0kawdxTAXmH/XyvuVun+ECZcXmx/56O
oC1Wrnd0/IT3oJZfsHuPAcbrBGE2sPY4pYShgXbgSLQ9bfK/3nc4CUgwgsEt963A
p/SCZmVyk2xL/f9FKPv49tQbb12o6sZV+uqrr1YHU3RJkcVrvAKIaPZNYOIXdmqa
QHHjObA8qPGBBe+y55XT9B/EjWNwfZt0UYe6IFEZiopzJtPhRFWosoUDPYS+OfR/
5dPXUPwn/qVBs10C2G+w24kawCkJYwVu3GoSothaCAY0oB6s95k+F9ijzv5ctVoB
q3tCwoyh4OMqgA25wqz+RJ/9MwSC6My2TucZu8TYelYw8BbDzbD4ekqnQUI5NchP
jLqy6THLgd777SCxRA79l6smGBjRcPhAERIKGSrDcOBBomfr0y0QaH1PCx1LgLqs
ZdARz0T48GiWnGkMdjQWipQpum2gKLPOzzsGZt/ssUgdEQMsPfdUxM3D8ghg38aq
jPDYIcZbpbo/3E8QeUleK7HMLwMOKXPXCV9hCLoeDw4svhOBloe32DWaStxADi0Y
PSFyypQAv9Ba0IirXU0aFL0ilPSwpn9qh7n1cJoApRcag7Irg2PPE9szNihsbc6T
JHY6U0DaybGUHppwSLYzgNmkM6bz0c3tKV/rK5ckmCm42aVgCRwlr3Ncy8X8+BE0
6DhM9aFvpLf0RQbU+QCKifHKAzgGa4KLA9oO/iZN+jTcwqcpS5n75n8Vfs1tdfYG
+zpeTzHroIwDH+UExciBNK3l9HjhSikqo2p4DUcY44lz8grajgW3c8e9wMS1rWGU
cZ0QZOihhjTo/vXgDJ2CBsAFG/a1atI30JKDgGVEK7FYA3J0NNMekn5zJXUTXZnX
Kf4gCmqBko0Bt1OJhWqCbtVL7VcVPgnsv8IjmkiJ+kbgU4dL9UxX0f5cGetqwZLo
U7KiGL5S0LoelcePtYqKgbotQTWSl6EwG7we7TvsJKTbgHrTTb5XGFoEwQkH6cFO
Ax5G2rUkjwLigi2hqiiYLgIlM+f8qrjonZ0p1UBdk8edg+Kqpuwvf/npIsQ6mbEJ
jRmuklubuGGARVQmjvIOEBjxO4yb83t42lFq+WH09nnUSaZwDuCDnUkE9c+ksYaG
bUWkB0FakQPPf8OX8H/VrEltc9lZI3mjpE/M45oyDOA3nNRVbl32ZC3tGDyGfSoS
1sb1TOJYW4rqGsplAvdXHixlFA+iCJtYyslVtSOKDEeu0BnTdA1vPhP6P8SWYK6b
rdEHFGzSyLWBJuxDSdxeTxg2Xr5/zahsKXl9mVUdPgrb2MZfBsJMRwRyve4UqBVw
ToJ1Jinm2Anuq74HFbvZbdY49596v63WPp2oi+W6j6Mi43dlZ3UCFlgZ+pDb7olD
0V5thNgDTdzVwbVeIuY2USsjT4JU1sPT+pKCX6SNn8XsJcBUiWo6HfJidiI8WxlB
5ZCEKAZwabcv0ff7uYxmzk61ie/zsUKGjM6qqnivuSh+iM1FeO8YVA+NFpCYZ0LC
8jsilzwBfeD2x5+28ZApY9icIDDyrXg093HtbMGe/YE3fcMr7swwo9I/U3GtDcih
OM3ZAl3Qa68IKOf/dRFSSYUjgJO9phEXWsO9RjZUPqfNmkb00OOvMvNYHObezzLy
DUJCCsmis6sufyoa7L6EPh4riVXAdJoH4mO2JfqIaWtbwF+8p1+QIsD+SBZlOF+Z
7abdWINkf3uzEF15OO40bGTUsWQq8u/BoVyQMCRwSWhlBQ/VKM0gjYoLFDOZbp8v
pDco/Rt3yYDy8NsPx32WFRQ/X4qE8cOq0uWp7VK3XNapWgJTcqxAlslJOokmHOvv
Vm/rbOY7w6M/B0bLB0UxM8H/ZB/qkf6bH5Q2IsmAzFThVbGN9MWK7h2LOa3TAWqS
hoU2vFzUgofSvmyCvoWt+mbTArAkO+B3FlBL+wtDvrrMhVjfP6nbA2RQIGp1X5Yq
CcD87tUFmAUxy8vnucsnYc0HDmWcbpKJe9kYDciqfyLP07D8wFkcLNmljbvtJjX/
KtGwwkIC/eAopb2CKhWNsbYO1tW02o58GnrQCCLYP4w1pizBfN/PC3zRBcn2VSfa
wEp5bMayXgIfkzB+5cph9s6e+jnlxXNocxO4+VtHtepJSR66oD6w3S7L1z4Rdbu7
Yfyl/gPPIypjceYQV5t53qLM1ZabbAkxIdbaa/9Oy13NrzQBtuwIJvqOmeN9wQQx
c2+SqU96SRTkdvaicW6g2LCmLoekhlltuJQpa//mpPvPm5gMwL7u8DrWGWTQtHxw
i19v6Fen+QtdupKFq6kf/lrZPmi/tIGOXv0TsnVvh4Pm9Q9zKZH1EKANUCq+hdIn
sl9KQ8my7NJ8TZL+SMwmPXPqDdrTzb9BfM64pckSXV5l2u+v6NFpBDxVXypffclM
dxwxvuNtKVpQ+mEIjawO3ETjXXu8o6Y7IzJzlRN1kUTf7ecFPxfPx8i6k418v640
/YlF7c9jpo0LJx+SW01L7reV9fiZBZlWeBB8Pl0f9Ga7CJaNNn4zDdfcsYNGiH8X
NRxncHWW0JPl/sXuijd8/RAow27OTt2NM9VJEOk85ZA8VMi7z+qzORdNpnxknWvn
uEz9TEa+0Mruj1/6woM1GywP6hKqQsZXAHhDNQM6XYrNmiK8BrN1s58rNgMJKpcw
QC4EcZk8/JwTXjr556hijk7IgAu8FyizDLBUWm5NbF7vNT+p5n+lxeCfKWqpLrD9
36DrFHn2qFNBtIkCYgabOGsVjoAfenRz9WhznOuH5xrqU08gLDdAVLxmxzxkbZCx
LrPsWF7vUCNsUCPMBZ/E8uc8dtoRR4iYS7dKbJrSA/4yE/q1yZ7sSbBsYVuj7oBp
ZDZ3UMQzb4pE/RJl4lsYDZnpHWLAjfBFcFiRrVPVqjI+LE9r/SBkVY/KuiN6mNdH
FmS/xOK2Kp2KR/+OOf8qEgWo2Xh8auke5WqV5dayQmGL2wuKNgqKhtHIjzVQuB/a
sAo3vA0Tb3vXKz02d0NySNXaAjASg+oH9EVYeAUcc9MfwcDI41C6N3R9MeKF7fn9
JT6RMXKhv0yHt31h630gZMgGyzoTDo6fDCHOjDC0V2d1xDU5m1X2ZlaYP7BktNWd
4XMLxAyRyosRZcD49RV19lYESt99Pt/p1ZeVVBv7SWGSuysDOy6eM23DT6xi5uW+
lSYf4yWgXSzgoNPeKSaBfXi5pj9yVFCEhP7uovmrdZgzGL2PbwPuv+JqACGbJNXX
OVcviCJEz5IB6PpDFXT4t1uyNOd4ADgIGiLCNY7zw2o7CW26qX5jywNfp2I3Jtxp
oBUSUHdAlM+HOAwg2yWYVfFECQfv+vhYJz0AXnQbF37yrhpFsnDshLH+V8ae3CaO
h+EqNDnISEHdQtqCCX2ysT9lKPpXlZby0DsExm+4wuov97OdznqdxMod1f/YIvih
Bn3IbvUbznOa4jAfokX4PKv5xAbFflKJV1aZb5QPVJ+nuCtzo44SGih5nohwL0Nh
LL7wAHrI6K5eoHh8v4cRq0OP80URkTxgMEqIfW4VjhXyiCvAL/2SRVvsHBMuRYHg
ksdeH8jh2Qc8Cgvzc8ORsYfUUxa9OyOcYioBP1wVtx69QtS4pAgnLEGfwy/X+wKb
F6ZwLVrpfIfszCABWPciUYQopLjGYIAkHoT1CBVYXUPuzDrtSsYJMyLPzwmcLGhO
4lZ9zJtU3fQbtGfFQMht0FWG8eTJIHRA7ASsvbEZgR4NMrezyvhGzLk90fFuEFEO
1MM+oDkuQpzxP9D4LEUdWPTuMsxp7/QTpp1UEswiwiLf+thybbJHmJ21fBzDubo6
gPhfzJG5SUsCtlDZHtU4VjEQd9T3xpzUdj4CQsk+OjevWW2gGqFLIb59jly0/0LG
9h7etwHlvJlBYsGbLl4F2pmMNkxhNxA5ZjFVn+DNVcr8IH0FN8B22hZLvZ3VhXYk
UGXU+h6WihcCo8KVcQcvwMhWXic/D6zGZMy5PGueVs45irOabquJWt/d/0XApTvd
hGkeUtapUEAaPdey84wdtTg16H7Uong5/NZU7+x4tFsfYvaF4EU+nqFytnl6MzFE
2jrGRj9y/eoIcjM9x3D2K4xCkUMotchIHvWf7HivHsirSRqOZtFYiA32muC+z1EE
kzvZOazslZF07A5dCN285zMCAgcVDV+/x1gElOSGnYRYSuf47jxjjIF9/L+Ump+J
P0jKIoZ1XDsd9SeM/xjNEmSlwdC8zpIw7DC1270aBiytaO99hWKdnyMeCuCYtKS8
uDmG467GbFvbbba3/oIj2NaVM5kSKuNzUAiFbL+B3Jb0CvL6RMTCceuWcIBDydTy
QBW8ZSwG5MPD08DeTUe5W12N3MzcG09LseOYtz1ZbFhB9Y4kSYdGLajcjAWOGCgK
DtzfqPavSkHu2waG1MeuI35CRZoxNX+RtPAk5eLLQZ2UdGT2XX03FWWVlnR2aG7E
1WN6cPTIw3wSlV95tJ07TYYO+e2uFEsMBB94/BkUrm20vOYJHVerQWL7IbwnUX8r
/Cu6xJ3CqcbR281xmmbSpZk8Qu6pyMYA9RTSsDEhvYiP5D/RyXE+zoVPgPMLkGxo
RHwKPlXg0OPhoLTcOTHWnlawRETbg2dzk0FVh4+D3iYZykvaWmZk/c9OU6epZqvV
DuzxkKNoa2APfhnKRcsUTJVhQ9nwV60kHMVUxohkgGnpDOUPZoWg7WDqKpuflPGp
skw+t/kdp3E6/1+XSP591uur0n2tp+s90FdaCle7j98sTR2RD80BtYnXhBtXex0W
7uaOxe+9hIbZYOV0nWLDjEZL7g0Y4d4i7uRpDlDfqr/EkI89QGGxViFdVtQ6dbIU
Mj3z1S0M93JbDmG4TtT4vDCVslWxjmeGVftF53kMqAK+dhr7rKJUN0LzrfQf9oKB
r8BCFkpaAenBwmJZ7Hz8LoXKT4Dz4afOI02DKfIo2jw/vfzV/rHoZ5adibusIyWD
4V2GAA6SXLUFAP3f+TYcppr7BUMw3q/H5LWkupmQng18PrgTO5hXs9UW4E0X4Fxc
CzFDlMwIf+JbzQbctk5WsAfBaYTY63o3IjpqWwfsiF9Tavk+WmMhGQZgkOJrGQAg
ub3KrdbxRo9cx0gv+Xzs7aKNytVff2DzNyk0PLsH0JOnZn25skAanFwm1MCWdvwR
2HWYl1Q57P9ULtbPLqDgeXDZpHQUCiTThR/4f6Y3JxqdOxw9aSCWLkFVNoYg1g1N
IasihzsX8Iji4xpB6RK/p8YmLYXFzzA9PBDCgsVns8eLpVHYxtmP1mh9JFpplWBt
b/P1dJuDRJ8gAr8dGGJV4J3dqult7+fBoKpMWIpI5EoGDnWu6uSzPPmhtYPdzbPs
m5MM6iF2GROyIXmnQyoVtyhsUrOlk6MeqChjlajPDBJ9/F0gjTfC9Y36vZp9O9qX
00fqOGyib/qeTJF5QSft+fPtHDZ3frdM5w7Iw9XxHOtEKWtDEkg9VfNFe/wVCXya
53H553eEx5Anzsij1wyN9N4wTbK++22rcOEOeHxNJHKLNV2InuYsRMulrZP8ZSFs
KIT5E+/NjHC6GRaA4mFP1qN4s2FQac3QcjjycLJ02Jn6WHQwVgXAXIuUBcf2Uy4U
7wCMk6Wz7h5a4Yuj6AXD1zU/fS3eVHCZiL8BXBXDNvsx0M6zHJGgP8/KkZMUXvju
QtfIl/dnriZVg9gtm0gcOwk8EWiKwm88HkLAZ1UczhOMMb2f848zSgArRwfW/j/e
LFlFNCXi+4ha9yineSadUnsNfvx/j6e7staEVAKJjVuKmub8RY4Js+Pd0cGoiap0
H7JO2wzQnGqnpQNEu1Nhw05Iwwzw6XTwkXicDuPj19J2u4WmMll7p5Mx7aKp6hqx
hf/lzQzGKBBJEluPw7PikEQS4mV19eA4w0ntS3CbxXsvSiHi3j1krR4ypoYU2Q4A
Z/mErx2xdbdC7d7ySxSktc3uYGDA4wJbjr5lN0/jLG/xnqoT4fnEDOP3jDse9slb
Ge+25C9w7pYYuzzMonLSqY2Tn9Qs+Tf6IEG3xPlNAL8zT6r3mMvaqnelbh1j3Jn0
vhVxKOB1CrDM/y7G1L/DuBERAQ3p8HM3cZXhS3nd0mIJl/Ipx/bwVb4MntWFzy3c
buvDclMZe5IW1mpnkmjo2FwqAhn2/Q81WydRsD4S1g3+MWzaaANtpcF6wcSuOE+H
CbAedxaR+jUIqn0+Docyu0SAaLDE+0TExiUA8gPwhp8pRQnEnaMp80NpJ46xG7Hb
BrlC3SxG0oFz/Zz5ejDilciZ6baKoMQqZQY40ld39E9uEdk3j+Ckkkz55IBsWQn8
l6AcHciWVEqbKbfjI6g5C8BpLA2qVZ6On0ziYLAKwlYUougzUsaBZDySE+LETOef
PYRWf2RD3/B4yZ7QBKu4BwpU3Dpger3i1ee0TFSi/j6bTzB6LjB+Kir1PKf5wXyO
ObwiMwgwU+So1C8kTNix+0aJqVNxTDEVa8zqLbzkfIkj+K5Oc8Yg/8Rz9eXHy0sq
AvrnjdzRjRF6owCCPdmCGGiU4tmqz22cwyZ8qRRpAzRhycXbCQUwSiCCjLptIhsB
Jo92njk8V0H7BORIYEePjiVbA8iAaZ7Z288baitCFtv7voDBTSpNkNEoQRAyu0cv
jdogB/DRPWSsPS7GoRFScwq1Ad8CmIsfCJtweO2BdERcHT3R0xrAwuYcqWqeAzjH
SOyqi+RiPhLQZBBhMYAuHd2VmRX3u+vdncqjr1RTJVnYkpQgqSzG6EPQjVibXJcJ
MvyjhuzrlH32nmsP5z0MxEvoiwzHTUN0R5v4Lhk0ODd+1e2QzbkhwSoLsnCXv4ZK
c5DmonOcoi32E1GrOIax8lGQghZYBCWZfwyt16O4795Dqc9pamUvD7DvwFyyaOC6
eoI9qtAGfc191gUjiA4WlatpTk3ufav9YLrsigUZyGKMz+C2eyucRUq5wLlEcvOu
8jWCZIVqmPez58dMM9D+8l5nXWyQRi7GuxWe+msXAFBZRLnAi/jksdINlj3fKPa1
XRWLCwRreR/Q9i3JlerUnSK2Bz8tvo1Jfcm1zw/IPqW0oLpPfN94X0vcUvnkroIN
viLPcdqpAbpfRcI0VT0wAaztukekoeUk5ueOiLFxi++ViIYjxD96muoXIsw64t1c
9mC9HFn4c0A3PpVGSPbUoZBnumeiHgtUcXVpuO3uHhahK+LFP3UcEcHR5H1HoHO1
i0o6+Y6EyJduB16cL68/PvhX5kxsZfLjd3C7OILH8AoumJMXwDiXjJm1cdWDGUxh
S7LJhIhgdbatVLUxVQv+X9leMsvBiA22CmucXsL8/v8yc0TIRwin/1DoPvhIS3UA
dEn2T7qfg7WFzaaMbZBKBUTMSW0PrCz1lNy4nVzyY3alqy9K+q11df5j0Jb/WExo
+d8qKNc1kMK8kyE3EjOwUiOVf9EvHuhfdK3yKG5JVozeLNJLpLbUiF4y9lFT5xNh
8X30ivIao317sy36xHS5E5kYMUH78ee05lKiUxMHrPe0qopuBDVaBHxmOFyJH9KW
NqOGVwpmqpJ+y7i0JmJtWxt41tEGWvmVnVJfzdLKsisOeU4j9U1Eqo+gIEKENGsw
XvHQOf6TNe3/7YMPQ7Vjk42epz9WMqcv9PcJHGE78z5d/dU6BpcSTe1VU69BA/BG
9wE+XfVlZAeGqPweMPsXO0NmChWwf54W0iYzxVRktBFET8HQEP2UC0WdbeGTPwG+
LKTJddgTXiOHb2R2xbAvMx2eQDKZF8bay/E+ly0HQUBWB6EzZB5S+qg3AdYDAmG/
YHxSz6lEPqzsQupZCKuDQ5jeKTAg9QL7a53u35TUJxz57xoPzdCo9cDwB7xMp7Nx
dWQTHCvemkSl48eEbOUVbhM50wUK/hTjGIm7cfX/JMp2uoA2qEH0XUzACyIPazaV
HZ+K8kxxHg9buWBqMujZB4AJIh2XKfuSVm0gJ04g8v1TXu0mMWqDBcs/v3HrjIQ4
MFowqVoqme2inGAbnZSCMhtlUoNCO7ZdFN0Yp/jotYiuCkoECu5R3EHnzDenseBE
EG7ZbVllYzLJ8I1IylDxT1jnA4JExE81EV4c3xLTIrtslCd8Bv1+t4LFv+tBE/kJ
Mftr5A4XDCyLQR3WHLHmmTUzl8KYa9y1ulFR9bkpxtAgo0IP5H7nFBEy8a04f6JQ
ryW2OarS5VmjcQgxl58iUMxSnRIb1NBpsDrV2LlnFg3mP3PUTiS+ZVCuoJtU3+GX
9DgnuFmNFVowh6CXt8FiTVbKGuYak1cFBO3W+8QoIE1wR9ba7L8JZK82yHrYSZdN
x0BsnzKzBJxx/emj9yIeVs4jSHywqt9t8ojW3EWRU0FQLy7XsmZL+/TAOvyzkIPa
OrNf4+vn0ZfyF4BuNAkQW5O8buW6IBOetzSXcxNocFVunxOWX9107JNkVPlDfM7e
xrBwJchr1of0MMrF1kN7bhjiPWzgF8GF27lSU6jQJebOhrfuVsAK54K2E2M/aTXD
H7zGEkqptzP3+vpO15AI13mYizAa8k7O8yUJDMeiq5Zt3rMnlhSeI4CtQfFKhZrh
C044Y+wDateHvhY36fO4GzuhyBoZN7dDLQTEl6+Ae5yPhOhJQwapMyw0xHD86i1j
AhXo2sziG4VOWqswW+V/kBwp6ldJjQAHIU3GbC9k5scECwdPmkBHEHxQRW7HKzL4
5keoJ7f/zey6MVI9BDooyWmypREY658XKA0NDY4n7dj0otAqightDuHO9ztIf0vI
QxiclBtPXvP3VRA5nYuWSRIj6vDTznaxnj6LIZlnXdOohjt20Pix5884Uf7bn2nX
/9BueYIjRgTPyF6UqvMzsG5ANvk2DKAreGoatziHb86RHyJaQhxvz1jyVHbx2vLY
lM7FlDnnhW6f3ithOQkaF5Hj45vt+7QQLt26/dua+mADjRRkScjX8WD5vbri5/9K
lHKYg89SEtU1X6cwwo1hAjaQmdVwfycP59Yt2GIWLw3zlD3tsmEZ+ao3U1wf4GTJ
LGvc7Zo2Zr8LnGra00Cp4Edzk+CrbT8BnO1bYA/Et0kTMYFJ/ISrlV7vz+sAZrLg
DmqQK3XZets/WkMo3+L9UfQKLD+RrEmgsfyjecKS3j7q6H+5Eyw5WxaZbTnTSPFw
6q+fCsPGR0wR0Nr+ltKO4IlgsrWigswngpO7o3ZSThL5KT33EXZFoUjMY1QT7ln9
rr4x73XrmQu4iFTCwFqNQtBWUbBYboaOqYsfOw8YTlGYK3h++G/rd1J6K40pda0D
NIwoZVDHRZRTwE7HSnLpyvHikccmOSt3PTGxgOurp5yb/R/yOikDQZLxE75CHABv
MKeW1C463+K02llwPKpczrihUyzyhGGzwqxSOs1kK/gBGlSG6FbmcWGBDe2Xkdkj
eWlh8oTrmyxYiRPxo9/jPWxnePJo3FR25sL3CXNyt3OPEvDWOXakTKiz3Z4VYpOQ
zk8lmePIlmsAxJtls+GdksLJWIexC2XWRjRoV41fGs1fccNtBdYBhkYqZiIpsJqz
fAik56jQYiX8otRdElzkdzBFUzROqKlntJUI2m3231fML5KAO9rhLsnwIAUbcOmZ
7oNzfABNWAQnD5UjVcoFW1H+XWaWM4g1PVQ2JGnVHXTez9Sjw4ilJDzEZBANoKKm
sePh2rl+ElJYfjC62h6RshvWBnz1u7ByAxufmh6MLFxsXHjqbdezKTXLKnHBYmiD
1Wyot5uFAtsX8HsB57CLp1zeBptm/VUdPodZFIaKNs+HA3ZQcDWT4AIHFGmzWe7i
IajIUE/c+1AavZrDgXr2liesCOXapbJUPxhHN5hqTA8xeuADuRzzyfQV5P3trRM5
dUnvjmvOfnIMf8wJmnSRsFYcXFSYCPsPTtNLBGVtUqXW/8NHBqYpSnJnhKHYAi19
IlgKBTubBsFufiT+mORmNDSLIgErFe9HImNhF5EBmM4v4ZWxo3um+KDlOVpf3ORV
Amfp1vFOrdyE7+3gCmTw/OgmnkCe7DKkgsceKElfNjKttJWT5vr4mk+er0Zt0SC7
/V+nUUfnacjBngBbdjMsvmJPjL/dJc/EXANZh5xD1jdlW78evgirhlAJQxivbRR0
61UTHd3hCTO/UcI06G4DtuoktSaPsKQySBj20jL3PMm0WrFNqSMhB+ipEUBBHWJo
nWZH254zYw1ICGu67ku5vYWoPicsC86dFzFW1sVOVYVRFwcr6adjA+Cc3NUysp5m
l0AGxqQG0aKudUx1DTuUSJbCICGTt2kzua4QGQ6eTqLaHar5oVbtPJkiU4g29DV3
g2/H2Kf1vSBSGCkqpahz/NOpl1zwVnUKmTAi5ezuogMBhfa+K91Ixen2S8vp55hF
RN/JDEjFQ9G/e+8pI5WzRQi8+8sOSSzfGfL6+B8qBtbL0MOK30pRvc3moqveh4qM
rU2F4O3AICh8hSpWTiA2PdLwMLdaYhhfKa+2Wrmd8clTkMQ2V6dNvleO28HoiLg+
H9+RkSsaIs3ufdaJpk20NlXy3CyK1aTPTkeTAY6I3x56U2OSOCvpWZKQCgT+uDvi
lO81yp9Ke3qhY1QmSBl70qhDvnU3deBYm/M39gSpZjdIbdwmkJeOFICTtDVFONU+
P1CpEMpNMvH3hunjMLBx2RCQSqlleR+Trv3tYEkfHWiy4j7orA7XLV6Mo+2Nfo1u
RUkX2mlUm1B5u5r/gV8rrMBwKbD9xJ2Kb9fdrMvdDcHcuva1FwnCMkISbqUKOoxL
KSuaKNVvfMZa1FwCjSoCSazKjAc+XyX2sNCUdY0dxTUkJ97MLDyPZEt/VCaUOi4p
c0aboyjmCLSfdeDYdukc0fH487jnBr0iKJGj/Pvucs7B8WiKSgQEOFVkvvJ5wYBS
Bv43AoP5GjmTxh8ebxzCk/j8MafHNZEAzlV0LNyfs4SkafbpLX8m1kXadjCTuvC9
9Hnj1D23LQEdFZ4iyHBBuVbarqkGg4F9YqTkECce05Jilq//YEhsWvBg11M7sld4
JE7J0vAlstY81WieNSlHyGpLYbqideMtUjRXO9w38C4UNf/bELVQD9EQXv/pV8Y2
rSqAkxcVEIdOz7R28xYCxzlxiP54+tmlJP1oomjlITWzwwuEHWzes9AyBy2QOfHW
rS1CVICuaI6jRFiPzpL/qVwU+nkrXRb8UXgU33s+X75w2crK/zUONvvsFQ8e+pnm
+F2pn8JrtcR/TJJuLMVb7F4h9/tUoXfuXYn9yqve4dsdWqCFKfUB+FKACNT3YFTy
EWoE0Wv+i7LFVfsTx1WqMdwx8O1LqJXyazhtZUG8/huJ6fgCWAb+f6DUMvEP/OPR
b9rBb3IbuZ4V5XJS8gOUdKT+Jw4lWqFFcgRYxMgiLVrGHhPSeRmOXPK9kOT1wbxT
Rlz3/MYPGkfd5774SjE2dB7tqR7VwZ2wh5QrERbTuYpq/dZBMKjgm2xQ5s1Otrid
BL8gkMcVXMa/GO0VesOyPm7RKWGLiL5V9sYgD9/tKvrD311sMCVF/nrI4m8Zs3Rx
SjU5+ZYJXNq3V3+JFi6Dt6vt8wA+bTSQx1SfeFGuovkZk/NCX4GEfS2QiBmHXBKR
trXAZq/nnIqJXRyFo3Se4wtaL4+kziYzwJkKO91vNepqmlRUUM09H4C8Cv06EIzU
lD5JQsYAmhZXv29oeWCOAj/dMWl1Eiy4TVbS75ICUJGeVQjXYAIJyl+7XdCPSzLq
KQikunLPWR2VkCnZARMYRGJ8rBErkBvIEzudbuEpnkyasO/1wTk5g3Ts6cSZgQjB
umZ9/MuOdHRbNqv7hQgkS41YqYhLSqJ28sarktTTPMGcyx/Ka2lQxsdc7zpdL6f3
ffzXoT48d6GisWlnUD+hezr9JM97YOUBOsGEA9Jul1bW551+lPownxRDosZWY5f5
o2gmBXT//Dfy0p4nuArHIhJF8koE88su93zBvHnw9np9yyTPu9xqi25FTCzLobpe
k9gzMP+lNBVU35vuSACAeb+HMG5VsEVPdkqSH8QRjVjHbG9WOWhi5N15y85q8a8R
wnNiF4qYdBIeNCQOnX3wKZCQLhv1Hb9BtaMd1gz3GVFIge0l+XHDCTWNgvPzkCW/
7cEXg0h7i2WE47frXlFpsU+GfzD1w0bDlB/eTOIX3wD7645gMTxqP/5SDScKiJ6+
rQ+qeVR1eN/ZaxOaBCXwSDHwgzaPSgD6EVbjF8uDXY+Z9fTSKDR14jccbVRXiNp+
4lmRij3ojk2cu7YJ+4D4BlRKyVTQjY2fv0L+itxgpLYxXpzayDpXt/bwb8mVECwJ
ivhpd3BcwfGaNavLc4MxAmgJicLD1qBDzzmlsvWTn51ZmhHLzRowsBfDHpFX0DKf
EOluynswZ+rAAI/aW8XlE12FZcAoMA+rYWqwaw/Ty05ZAB6vCuHwaqIXxXCtSuxd
LB1ZLq7HeV0SDCSjzlf7lrL35wxFj+5OTW7nAkNOmEBAYznVGwEnofqfI+TwItc4
3/ZNHTToLeHiCJA7ThP+r2bbuVE3KprY6VSMIAV6MgKh/xnGBr9q1BoTcTcJwK1w
BvOO322evktNRO6afxIJYBoZjvu7j1F8FDwxA5+Cj+2274kasiaj/OuUAkuyJLov
3qcFoyVhH9A/QwIC2yTvoZ1LoX7Tx+X3dZlu02FVGfYCCIGLseVhFWcG3xfLUUP7
zH77K78/RXlBq4HUeSMLcBP/bj+857CrgTmmhVqv6fwy4KW5miogXA/BA+hmdv3t
6O/d5zz5JmzVZDuehrS56R98bY5c5En4NjeJYF4TUUJgZFhBSwMRarXwFd8pqBTu
kX4I2Flb5i0Ddtdzr4rGbLBx3PRMLnfAljP2DunQMW1pNMQRXweaS3kofGG0IFTA
x9ZStp9aj69jmT6sPrVEm5c/vmnCj53aK9WdPAjjK72R0BhvmumVmCBWFhxp8VIe
e1F3ldb0zxb76PFkho9iR+2Vs2Sdv9ET5MRQZThTYrteI8PsxXeQwcKbzYnErM1u
mWfJvfZCzUypQZUA3wc1/XzPTJf787BvrsU7E0XEPd0eIcEqhx5quBa8n0FrF8A0
zr7S+9h7Gi92B10yM/iVN5gAs2hkaYSeRr0ca9BfU/yBX+BpIPdZbwk9nEjm33+B
DFAEFgT9age3dk9OM94BU6/x4mCxOA2XxbS0P2pOawZ6FGqAosY/1DeDmSS8ukqQ
PNlLn4PHN5fBEUAxOAMbNku6zJtTWaG9hYg+5OKqyrluebCa2PV3DUnlI8y5sFnD
VF1fOtJslOEAHmbXxu6kyFNPF+uFjSnXjyGbdmo6BuJeg00Zj4a81/PB5+Q4rcMo
K9RIwOuP7O6T64eWN7yzJzeKR8BFdW5W2k4onhCcwlFs/2YqZd9/DDDk3j72su/z
hDS5BOq3XjDLRsHYgH/OQ10Po56YZtIUeYiKBCOtTEGsO/uL8IfzKmf+09CqBJ9g
g3SG2fJEy5vKVK3YcugKybQTauR6FCXx9GroA3HpZnFvr28G0/K+MbNfJYoiLRre
UYv9HBosmH0DWVkIM7QAq/siNt1SAnF4NoZrPnEOzHuIXgErUnYayKfqdUAC6+KR
kAVT+GvscpW3t0ah3HttiRUOzWpJaAjm/ZfE9mJYV+K0alF29lmFgheTYEJTuJ5y
oJZG2nzkaQzkOS7wdQkwYnocZiP6s2KmrG7wKbYianBvPbOmsByB0DosWXXOioIM
DgPcYLff2/iHz9eIboimyxUR8w2XJAnDuI61tcXc7C231Q9wjtNIfDh9wdFa0SFk
yl45fqDf2YrkxdITP+2JRVOw/lKV/dSMtjqXSHSTta2Wh/q0ZBTegSBOYjDUqHq/
kXBA5pcgUiXgFmAy59O6ul1f8xfiQaSTBbyIv9J5Ijgmo9JglB0kFdkAjQdudj9X
tdXzFDpfAxMXW5B+cFQKVcgXReUwSLw7PKV7Jr2m9Uqmm/bWnmFyopMxEENmYR0u
SH9y8dgqEfQbxW1ICyvvirkv8C5E2Lw3kpIs+Rbzl0iD5Zj5lKRRNR2qgZfIJJJN
muXWXPymZO4xrbYzc4dUp7daaEOsxeb6vRDtCI/nr0/vrF+ivzQ14zLS6UsdDKTO
XxNty1e82CUEIClc2CAh9eKzwOubqj5YJ5YPr5SIH/M7KFsEhoNVintntS1ZNhC9
KE6cTKmxQOMLTevJhytnjvrbVKkJdYtT0PdNn0acIsPyXjXhP7eIyinSt/5BvCLO
E8ZJO6T4F5C0s0gSbn4xkTr87xlkfOKLGDJLcOwQafKFlajvpdCbeObfj2IBOJm6
hGQLxo3Esv/Fys4LcA+truHvtKKIOn/+a63yK6UIHeQsrJU+JxugIcU/LZQiNfIc
g5FImQYN6ufqyEMTb2x0h8nMvwrVoYe2XD7YOm7d37aY4p3Htm25b6oYFaQ7LxKH
0BKeHaNFoDQXUUR3D/dFmAESp93I6KDi70H9geF2DCEwmsh9suAciAkGTWmw2DRq
8D2RjJRHW18bR0EF1Bhc2ZK5wOOl+T+Cyj13levplexNs3P07a0AK/6w3eFVIwtv
enq0p/9hoixp/iNVHF3jcc93v+3I+qvaXsiXdubOSvYR4ycXCDfaEL6jobAurRDA
BHOG0geQm0JinXNAHYGH1XPbw69Vv2+FBShSgOD4Hrae+fFOjq13RO116dKi5Tgr
cFAUZYTwyz/AYD5n3Yfk5mwNaYayqNbA/htlFhiW0CnOsF4r0t1gs+dHgTWs+Ue+
6s7kjamGFTNq3ti7VEnKDg1RUttJo4HXQbi5gQ9/igVJRNAefAuZzsf5uWK27e9D
f5qwLcNiy5nUKVXn06l8hw275WcNY0Dz5uY9yPpieXwGjgNo0gFmHKzCA0WhFMxL
Uaym+oM31/1UFcjKXjWu0LSGsqQTEq/iycHh2OTtcEZeMBE8ibqSG5NJPkCN6Oxl
n5JbJ9akVvZxORjjw0Q/llOSJAmYCEW40tfjUwWGABRBJvWoPZhfB2aaOqTDyHab
WTElERADFSCwlTSM3jNWejFpGxEQVcNBaUz+zeCZG8pP37zM5qKiy3yA7DYEUraA
LFRoe/Cg3z4PR6eeEQbXZyt+Jy3PO5py5IClLtkI6ZDojXNZXwWyOnpKpEnbEIDp
1NW6epCJTOWboTWpW+mgQqP1a+Jl1WMLc7UbrxlFDHkIOQauo2ViZ6i10hvklyaD
ODRx2sGNK/1Ql5gCBfSwCE7nnEyQ1NJnXmNpO1ZsybdGDfFIFnPPQ4A8fA9QeaN3
O/3FUUTvdAShvUqCNu5/PH+OYIpDFbAfWjTUojES3FO7j7w201tIqZqdDd4QGi9d
WwUnbAMkWXxtil/rsUZitoS0UpqPwwDVuBoI54PkzEUHeU+UDx7D9G1A+eHU6Eiv
9rfzDbfTo4szMoFh590SZJ4Dgd1X7hauLU2CV1HwaHLNUNimi7JH0Tfuh75yfevn
qi7lW82eJDIQXdsesbyQjiNDP5G7OmJzRObMJYbIAEgcXanEkVyVqvMVrU4k6WsI
ZjbKG1Lq72MUTsyFbKbMo/gFBOXvgC6c+zkwVofz7k9BlM0UV7+/YeFxvyCZDCeU
qQYsNO79kkyWWiXthk6ivHrRrBBbxzEcPOvdqW6F1qjLlvCJJJe38q+zk7zhs4So
L8mRugRcq7PIVBU8WGN4IiIZKqmNYaBIlJkkx++zFVnzQqP4nhGy+MOMSJbtuF19
9dgtA5qGbPY8Kl4hxbRL+YsseK0Se87eFf2G4vWjvf1TA3VrOh6CzGz3eKyR86XU
V6layMgWEI+1FtCzkeeT82MfaMbqlvrOmQiDY/t4FcVprydYX/JPefNa0xHgpvI/
bv9pl1iIeFaT+05CCVRpKRvJYejA6M1uNtumFiOA2OLcgS89W97FfKR14txWueUw
YWgBdqaXGPv5HF1gOSNF6j52XBJnz0LtJ3sKi+c07xUQmQ0K54z4AJl5UusMx4h6
UV3sELL029XGvKFK8sQ/5m6NZRffyimH5zap9xNh/9UNzaEK+VkpKwWVC3wJJOHe
8TcFJxtpmgCBKV2bPvgvmZI55v1NGyVl9mBxVc2UWX+Hq5RhTd91vlbPSAqpqM2P
LWhuT3rvz1UGxnpgoC+um9a5/7TiGuCOhSR7uc6zut/Ywnt/NjE90KJX43kff/+t
1BPFAFtfW1nGO7k1bba9kl46gpsTXWvFX4vp8OrQUCBjafpwyV0N1VhbrRGso5XY
8RNYHvCgwXVBk4VC9AAkR2QMgVPQqPwaK5cQJHWPPZKBjfVKbGc2sTuGelKrP8i0
WcgIwBdkuULI03x+7+6Se+NROjDfNI0DOR0fEKwBqgCcW4wqNK+2WZhCMh8BfSVT
EEEaWu/FQAC7dBW6gB9OYXXrJXX0ArWh1pInu8q3iU8P+uDVg0/4U6c6lyK6Ghxe
6m/Uv2g2MEB0GWaHb4ei83BRQiWmyI1cw1pU0CYYmTxqcA55waW0YWI+igscV96N
Vh245szJlswgZ4quNKayqwUy3kTRrwKDfV/AIX5wwE2x/gmIC/mKnOJSN27VBGlk
DdICkq4cRO7vbiWZbiEyVvCOeHwmWWvj2Sd1ObHrcFGA5Q5/X8ygY0LTXaygJ8gG
3C6s/64hCubtHEka2lbV2vTBRA+yJJbQ/ww0t3gh43mtJPXj3eCpymBbC0M2h0Qh
2XUodoZiwc0s27O2hKkMvRgNvGhCmJ8nvlPWylkqsuXcEYLuplXuCpjntm6In5Y4
vCfQE9i1250ToIyAYyi3Jf8stLcaOBdPvQ/Q4ikVotp1BDXZT3SlVmK8cis1PCBr
zV5aSuLHHQcUprvm2V2tZlfNesgN9wwYbQ4tiXXJG2o9gL2+xsb18dLOES3xYcwR
ueqIPZmFh5nowMZ7vVmVQYsYGiRs4mhAqxZbV2AvwJ5mNScJuBbIuLta3Nh01+y4
/GIKQpHRt/OKlcLYZP+ijCBOqxfMHLJiVJgsIxrGNkxMm9k0jhaTshF+n8+7+k76
0tkhjndDkKKSGE5zrO2ig+Bvf6LoLAMDZ5ZrqiWA78HVxGSqD4B8yjmzqoex4LpQ
dVxraDQD3gix1cCaIHVrTLbyVHM7fZYCbw7gNO8/MtoF7cPOOwlWzpUXv7IVjvbw
SGgq63Hoq+5AezW+wIOhELxcfwjFHcrf3/cURGgfN6cn2Tagp+G6PWFScPvxgiaW
3WWj3+0pmVQsiBrP6xbDwpEe6zDxO2RRIrJm1Ay08pI6Hg79E6i1IKkG7GkC9klZ
zJbIG+qle0iiSkiiZJQd7C0ctHRNlbY871rNHlKgITdMio50O0k6ZiRaL9499Ipa
LUHVjep6P1boVW023VRLLhw9YXKnOXjh7r47I/blayJ/uOqP5fLUxM0mK1rVom5L
VqD4OWH6Sm6GfSGsMbrEJ8RnRtwUz19Xufa+lso0nyhP4tB7IC/JTAXvdOfEJ/zv
7TtrbalteH0R0mjuKi9IorJ38KmcLRSdNrKrFitRdUAVEq1MPULWpdEW3Dk/RVCI
ZQkMiS7rUQEFU11fs3DUuYOzIDwnSZ9f/Qijoj4J/Q0UHpgrkvGKzh63YBpg7b3E
OFDUwfdK1dxPlJRwevVTNuXGs1q1B8o97ixvll751TqbdEBJgstj6M4VDSyQ4cnr
0lpt1QAqSvIPA+q4lFtTQfz+GJuZaxNKMXV4ABjw3mSwHfsFISfOnz2SE1Y4Dggm
YCM2zW9+l/H3RE3tf1FU9l/K6cMteub9UpqZbl5UoIYrLjGA6tTLhDTsCF6pHR1R
qAVNNpGKx9sUCrd67vUcFdAY55xMPWur88a4Hl3CeamBBfbwiAjI20Rn3EXD00HH
w/gji1eJIW+c2c+OibOnEG3zJnpMK/IBjBVEb0cBs3l05DHqNf2HanPuH8rK4vjQ
LGAbbnvavd8fSNzRJS7V0HjARegrRm0jsxMP6yI2+sjQmFxE35uJ/gEcK5TmMdAh
0GTj9FJWYzWEhG/Yc1WM1YdzkFP+0UtsOvDZHIvXqpNiFMcYkk2GoaOzrTEaY1kg
Ro0Egyqxf5vQT3nLnDwTGVYCWY3COvOQLLWn+qY6CqIeLRYsDOPWGE6QQXmkDhRw
BVeljy6tHCgTb9+06CnloCJXpbardVj7kqIt+Wl2BA7b3MDSiPAE19Vo/HAelAXH
0+xq+L23ykYsGTWlRvURjUR3/tZo4OFKP4hckozx5yHvcJ+DvLrBcbCFV5IGYgLO
HJ1wjQokENYBZhvqihaDmTwQ7+OYG3SnfgSUxrqc80V72yIKx5rmheBRv1x+8ofZ
hoHI20PYcqHyG8PrD3dSY1pkJYvdSGzgORA8YeTiRoim1po4huebf8MTJswWTl/i
YxLEeYky9YKODvMyrpAThgEgqsK+hNrh1URIOr/kHYiaSfR/p1xz37030xhLs+hf
1cFHOil9KFiOZUvYm2Og93mXq0nQtZAydpu3OAhC6JaYjyyHehCKtU1X6vOFVw4y
5+eYlrEvXpGYbejDGW2NQqk3oaJu8Fh8nFV8EHSAZIHGycPMt4bprcu/8fVL6t/n
L5rb9n7gMcALpB/eBcAbEYqERSBDQnB1mGuCkxBG0u5C3Z6UDMCaEv6151NDT9re
osQF5bCoCotJbB0iqZnwh+Qt2k89+OPdb0H3S3s35L2VivWEufnWJOFxDik8idW6
thLaPWJDmLa3hSJffKgkFlTw0AmR+C1duY2/x/So5o9qYMr3ig3fTho4NhB+myFg
BRUGQckTp76GunWaZkBmjc0KssnEGVeNQ0oxBuOJOU/9xGxisRntzUDaDb90iWun
TU/GDN5INcqUF+zgyDjWHw/583VhNFr595x0Tm/OXMeZwEhYifNlRlPq4VZ1oVd5
z/gWkmYpMEvjzjKii5I8puhrSO90V/aap97GcG6AONeQpbRpV7RiVqZAuXM+7Nq4
IH3CI2sMkknkmcHKJiL1wb3BsjLVi0foPxi9nYalKsGlR/nG3C4gBlem94qHfBVl
+OPgRKuErNdbtEBsxmfv2FsDFcWR0vqCrRqF4bgFHo6y4P25zvNrWuf2fcL1HvIN
vwOJQ0uzWyIRRn0NTc6jZkPKSCGApkNDdIpUZzbYZcrVPKTe4XQWPB2Lobo03mhf
7rOLaQOM5R2RwO829LHjrSCpFgccX5Qrins/x2PpSnmszp4WZtxzxHSEm+1I5GIj
S10VmE15pIc0SD6pI3nrNIzOPhXMQISH56iiBSZ/h9ixSNGl9MOKmsifcWzAR3Rc
MuPJzNstSc3MFP2QcKUXJc3NIshGkv2bIAr2DJckX5SdGeEo1sNUY6buHCGD/Dvi
TTpjU3K3enMbgcBdo7OHfsxHxKAkWtI4bSDZXsPRcl997Mffz+/0V+fLGKmWTfPC
okGHOUJGpDSrrIXrbSkjPCKpmKNxs6sZuaP5xeAjz3BNdoo13n0bwNRtBI0kU9+U
SPdWpguC5Ppncpnbg0cLvj0LbccKNIYgQ/q6Yc+H7JU6gf6D9NpHDiMRuhwMFt65
yACSIPeSRvGmfvAJCZn0pyAGApXaAJjjpLEXqX0HQ22zcE/hapi7ShLusxttHQgI
wEjHIi3FeSKfgqlIU31gE4O7rzteaoPDTdacIbiZjxlM1VGP5znHstq6NqgelSNJ
BNJmmCaug8mnqqQL5edLGFP+QJrtph05jzI6BPDzJ2WHgF31lI6Q0tm03H0CkNtD
ZQG8iYdRLw782W9LV5tz6raYm8giq4mQbGW7XhNd9I0LOIadElLioG48381E4/Et
UX7iZ9CmDTR4mK0VbHFqNJddtMAgmnO4akvibaqPyvY1nW3+IwgM8/LqnHOaxjnc
Z2XrW3tM9Ja9k271nNqVZtL3eoVK7uqWN5v5CBeTA5OXtD6Li+LhqrR4sw2mF5Jm
tgUe7nB/NBWgu4wNSxHfzwB28EqsjYY166cdmcCdwBrt3HZuVFTjiM4Vnf640nV+
hmGwgOMxvLnubS4Uxcs6LhphXSj+8jCk5nUQTiC4hLMt3fLCy/cdlVkBXWN8KLNC
Pl0NBdwzMdAQoLjnPvtUZ0wMeyJhpA+AXFF6Io+N11ssWIGxV8/MTIIHsbVSseKZ
6+1ma+FzA8U/UTEbW3KbM825QKInBoyjHZllSV29VYroJI8TEyQfd3q4YKEy1mPq
Cc2aFob5HUnZSR3LUaeq6PN2NKw5RU3lNIrCtXAin9bQz824TTdOt1k+e44Ctb1R
fuBmoF+wv/wl7o+YL3gnyyFmx8MZ/osx+bkeccNsPf+J9AhT5ut7+hsbkC0/oJjD
UxLksqOSw+wURBf8uB9X9SVqghurxfkY3bNRbau/360PIaHon2kRDCwfVSGp3ChC
KF7/MwjDXcUT5WiXBcCh1E+2RMBV77QL9MJ5htBYsO6yZQ567Kjo83ncauxj8fIs
8kj/117DnGt0vvgPYWT3mCVFilAxpDKw0Z2lK04VAcPJVz2zxLUe1QlhY0fkoq2M
jY7j9/fLGTM+BcJwKDs2YZqMziRGymytAUxT4bZfudi5Ji/v7ZwMO5oKi7RWn4sZ
aaTl+zO3P/HUEGI3rhjyj05lGRkry7AEEfM0TMaiDXyRdGmPjJDEUoYjbbxXoPTw
ffVt02l9pd52IGRbNJKwBU9BY+7KMYpThtWwEg7TTNiTqcOcxlGcGWUvA4OtQon2
7B5rKCJhR6T6SSQ7rMxanTpHVY0PoeT7xnLvhZYZHDAg8ciXob/MrKKu8jxkmeZq
tLm06qKfiyivtiHj2ng9/hE7Yt5PuCjwYcKhdqUNfjMv/LL93ANKVIV1D40u6LGH
hasYLmthSnAkPDdNIOINsGFGoxg2V+URAZTOA7bZ2A2WM4IsBVw3kCSDVZQa5SSu
LmefMwDehFWuvIPDIiYbMKRVw6edYn8Aadg5qSaMeMMEs5DEme6lPB138qvXhZ95
IqoNOtJ+g0GQb6vQphu5kHMz5JbIvxj0Kz6k5JzH0GRXFcaR4Bf7IaOmh/o4gTPP
D8vC5xtsZQy6hf+CTAQS4WGqafjrX0U5VFquJOXMd8ZuCtvgPvuFhd6oN5iHT/uO
4Zm6dLd+JknSh3QW+/OvY/lUDrP/wrzFp5r5Xgvvze4t/1dUjMIiDuCPwSiY2tz2
phvEcSCRzULpTymjfdx8uwVm1+Avsk57OvbsyWrBctqrTRYH4DmHbczb/bVcGc5I
x64XaY8MCuK1GepqmoBKXfwVxd6dglNHB37Y/maRULd7uRSyxYG72ewRCZ5JXCiD
9r6nOgIJBum6XZFfiWH034Wm1KSKf1SruL8bQ6VIN+swuY1dWAsOwcIt+5beM8vs
VFtOdORiQyPywb1rQa/TOG/DuXsOc6nU3PnZqllQ6pR6Txl/09f4tVw4WyR4sw7A
3nJVRFWHIgPfFKaoOz3mwAK1omeRZOzV2jKWZPxOrch1jx2fKEfBOzOa4ekGEhwP
5OMfb7TzMjq0DN5Uz/m20lAaSuH5h3xwz15TD+HKEoy9ZsBuWwT0BVOfZ5CLUZxv
tZNGSdy03ojE2ZSEWaL2m9+H/BZ5v35O6/u5ZPtjniOtqfDM32cSL7VSxJrX4PtG
OS4rLyrSC0efKcHwRtzL0W0lDsWXx0M/xVqC+F6rDSAc99RCPAf+3c4u1TlyzCyr
GD7tKid/26HrqDfVtLvFjXBqzmygR7+vdVxt6ezKXfY8iiYAS7vDNXJ+6w0bbyUy
58C4Dbnb+MuSRKfcDXsiZC+POgMuQ7FjxyRckCUXD/Nv0Y9Y/bWju+qkB9wbgayu
HqhKRZyL7GdAl5R962SwCtBqKlvD88q0H1a8AhB+9bp28EJuDDJgeHpBmfGWLI0v
0KorECqcGeKENYGuTHNxMES4pAOVx7n1DRWGiBxAPhuXauL31JYkiVYRcVyIerge
qvN/g3dRd8S6rGouxqUIES8Aa62chfCcEx2N+pzYpQmn8qyufrw8OlSLAYoc2ZDy
VfjnNnZSWFeeXJVsqxC7Gekw11xz+S4hwxsfQ1v8wqRc6Zurka/OHOYlid57k/D0
O6y5LNmrGd+S8++5Z9Dk0qiPfae+0MegtjkZl9FmR9BqFa9aoCV3AzvIKCWWcvj8
O3J8grryhpOX4FCFgDFeXqytwPQB9K1ET21w9dwCoXlRNadUnOwkI5MkPTOEXR9V
Uq/fdrf+IOzu+86cPcYejVnV2ubLk2v7b8YqYT9AhJRnzPbKPk8vJgCSpzGvpraJ
CpdCnlNUIDD+sLurXTZ0bW74w7fBH680IYsihaRnsyYanX79ewiXxeLiR1rMTQAt
cKIleM/lHyGK0fbd9bjGppAqQgNb6Jko4MypfdPn3dBnEeNMoXHAXtFLbNHCEJsD
jp70mbH0AB3lwCn2u5H59mZkzeQ8jkzJta1fZLtGrH/4XNl5pQu2mxZAYe6gG+BV
zDRhFwqxMs/UXfK6Cg6RayBT2gykpLRmbW68og5BeaIk/qtjtzQ7sLfCq5XV1fi7
+NPwrzng9otlhamjGVKRLtlhTjSg20TsFuTiKoRMNJ9M+sJLoIiRSFky1R0WJaa8
I/g28ydnwipSWC3pvlotsSnPcMS4Plch3bOEBlnhtA9lEYnLRgB+bcuOf5IST08u
M1NQ/ear7dMyQto75y0DLU6cmwlcHOVXkJr0amdKXYkcK3TqhU6CJrQ2S7WYAPyd
SwWEt0WSod4Db+HDliTfBYGrkyBdeOO0DD7ejjIuDMcTjDlAsY4ToLoPM4c9Qn9q
aG4HCRNJikfAX8Y2hYbOGthO5rkTScPIDJjy9DYi+AWjQZKSOIs6tvSNi/DTjW4p
ccy69A2w5fkqcz2UXktfjiO/u5mgkfW2aFEmNnJktiBFikXqpNc0dozoKFoZYcMN
4nE+xfIA10eUsUmX9vRRaoWia97Kk+iCBL/lcMiUHJ1XJdxDsrZyd6h1/78ZRZtr
5T5xVvoUVsX+i/2esSp7zuZeycTYe+6mF+1IxAvebYAyDtIiDjJ4Hp/HlfDzuDt8
eivXyht313Nd4jcB6c4RVhETmvhn5JFv072c0f5A8sFwITarnqyPJv/n+VE9tP2Q
QgTqPcpbKKB9HWhFUC1U1mpz7oYE8E5NmUeJ7c76TFCarMbj45wNJrazXtep+FJw
8QbLa45MoOoFMEGTWAfdoW9Td3DDx7+nuWjV1CjcHoTIEN/QLJ91DTFWZFAYPIoZ
vJrsOv7LA+XHUNEysEbNdOpisr7ayj4H2k5fbs4cTWNy/SlbE2UJgx0yH3+gqEP+
exSzh/2QxtKidfs/4lTiBm+eE2BsvetgPQJLsa3/dimXEafAfkhUFWiPUTEnI85l
mry97RSo+9zPOvqf75LvCYYAOsXD0g+8LyjKm01m+FW/8xegubqjsB9n0wZPpqEd
9L9eS4bZwD4VztMq4OUb3s+/QB5StOb7HbWUhAwIOGxcz/9zdA0c3LX0Z/kTqOtM
lHX9ITnVQu41hnCGX/Z+jy2UlLMNRNLonNvFEQiEsccSw7WXsCLUc+2byEQ6RT+L
xMjC7M4dnX4udpuzj+SeGwFOJdxfeU2V3k5xVlItcSFfADTkFVv74ngSTbZh2RjI
p3MMnLwQdxvA05sXhKtDZ/zPRIJ7oh8Oa7J3h1BAWao6ZS8Yia1jz7HSV6d0X6Kr
WHlCZZJTXEcTGbecDJ+6p+zc8rSekvcNmxgCcwOEtntWNuLWdmOyKYt5PqJZAV/7
uYDr3dmXoBe/zLpnPIZIWrNmuFWUJgiK5qglMV+EmXfJZ5ofxv4/3UK3Ibf5L7Bt
D766GqIcZ3LCj/4obG/EamvT4UD9xIn7HRRfNCeo0JnD83LCKBoQYWmFk4vZYKPV
XhdEUmQAfROmLifS3iESOTni0voCwUO6APqWhk3VnqX24Jo/z3t4vwZIFWvoca+G
wB9IOF8WKo/ID27ytMO3MiyO0oNMsq+/jEXkAeEgpGOTbMyLQL+EnXbfyNyMNTQG
xgwr1vfW8biigeMfFzgIIGxyMusq/qrqOQbzZ4k659SwXxK/qZiC+nGZTkcDLyPH
279N3OxrJIC+ssYAy2f9Nyz06l1nrf6aD8bfvtnerAk70Tmbp7y559HALrk7vSb1
SuYH8h0uq5Tj1jrap8nMI52MkeEGBfE+0K0W0lsXWoDrE2hgfwk4Dgo9m0xwd4Lr
92/mKz/+dcew+2BkP48/DGUkTNxqroS9PRozAgczkCDbpuyKo/N6QpYztpGiv1q8
7Y4nbI9gCmwrV9eLF4EysQ03hyUFLiy0nlJYf5YQ6ry/uf6qFVm/MTP5HwWBIb6u
ZQwI6rWChpkIuMuT7LUg6tVQZWmehhGHOHGZzVH8r7Enb6MQ+CPPRkdU6QVQdCyZ
3X+RbTDbIHj9qQHXdrqEEjb/WvgY8x6oCl1lzYuKtcGxHn51WvqAC77awBOFDYBQ
7H7pgvyPF4oQhPQwR/KD2lDs7yRgf9tYlDHasaVrNMhJEj4PNypvSBHfzp1p8ADu
KboG1nAak5S7O+wzCNaPmTd9IPiulx3rKUeqcEP3g91egOgnjVmfEKwdFJAcxv/o
qM1sNHPd1TuaT0ezs6NbdkDR3OyRing7XzrK1pRBj5ag7N/sn44H70gs6OwqKpzu
1L32cDw1i2iLKcL1tIrOLslzXvA07erj/GaH/nTlqLsQI5mUAZNb98Jp1dDTrfaL
1Zk5AzNzpcSd0SOgEW0J4SsSYNTx6OKvcnUU+JnJf/I4ueAkEOwt66ahICINqFVQ
iCrPOBCfTowyQsL9aqZ7lCIdeNnDFMnKg9tw+qL/KDHn17s6XLzjZvEK3Q4DqLAc
DOSOcNCSadGnDUfNR0w00v9wpH0tSW1dWbLEkyYIXUyrpjXZzNLv7SgO8g7sKXz+
p2X5JBHBscH6h3CIHjXwZ9tAYJ2Np/S5+F2RUZdWMb6MUY3qWYUXMr3MsjWq3+Ze
oEpA5jgjDxbpVEMXlaoMXijdkCMM0fdUitq9y58yWvu1G/JALRGtwhOldk4Xu3Is
H5n0yzXMozDldnxnruUy5udZ4TR7Md9u8g66QokZq+Pfrh+nw/HsbZ+ICCAXEupa
L1Tv9vTCMOFuS364KWFypjA2IO4i5ZQ1cfcRCrhe8BQh/WQUHDImH62OsB4trpiZ
lQZZe5G1Vmf5R13DMOhJaZgpxbVGIq8Wfg75iViuObuS+k3lekGla2Pa47eatgM/
0a7jda+TMZtH3OJWu8RvwfAjDq5/33/tOaXmYw5HnakAG69f59qH9xm2GTppnyLk
YIfR37XkzMM+3uZ2BAbD0ZUYudN5WklcBWReJDucq5uVB6muo38kzoESbRZxI+H+
CABQzPoJu5MZo47K0RNwabnQvmTUi4LxD23/6e5c+o85GAcSHuuGsrPAdqiki8wh
o80bvsdx2lO7+WIRvCUsJkEmIFn/966fwXkBD5AdtxPDmHTy2MBK8xWITqTHNNLG
KM5uY6COa21J+0GSyUkW8y2eg/4ixmxlUxd16fSvWOHfVtzD6goC88MvMe4CjXH2
j4agXtDuCYmJeA5xn1yKkX7iILd6tn+4z8nuJl3Lmh9CkKk5FNf8RR8SNujm9ZpF
CdUU4pZSVMRYQwVTcEQJCYpobTGuhWyyRV5pN+mHc5yHo5TUwK2IgdOdnyj7i6Tz
JQslwHUTdEQ9Tvrao/Kym/UXUm8PdkRTMudBWoE3tvPqV9tk5CzMgWDto00VZ1bn
WXKOFONzFR2MFKtTBhVzWoUFj+6O0BTqrCGt++7C5ujhYbFsvV4WNhRjHVrrF2l7
4uiyTAnpKHZuP/aKydEa16CSJL0RDZBrRkW/Yv9pkYfXitOtEVh+KQYdngX+J4Uw
3EnuXbMvPj3a7Ok3/VdnSWvIoEnSTghKOV36v7DE5YepLTbuAzinGfOMXMvEnqCt
3GWuJP3O12Wu+q9Z27fQmC2Jkrj9skJ9gv4fIO1ucy+e2ab+CAoWYiJi1RHqitSS
1NdxDVQieubsjZHRTqnQ+kBJF3s3cToBw4tRPHlNQ+wLOP7a2il80vURBu/UWT0h
vLbBnp9wcfA/O5t8DcHc39ybQ0ftkJAMb7QbuzCddzrs8wQvOla3v6JnO+/wzSvK
SxW5DyV5hg9Nt+WlE3GJaNDAfndsT5E4wFuQLUKiHDzsmvWFJhPCz4o38Br4gswa
UrAIlMCZ0XzgpggRHXagd7dDBkCPDFqiiWLX2AXMHocytKWMvP0CYUQ+6NDB6uPm
F8Ut++2Fbqr2c1kjwSapr69PEiMLTGk5p2exVaPxsGBlJKJWIAb263+UZBMGQ7SE
sH3n7H/07mrbLrGbtNpwoEUD9TtTKay2glRKwH547V6u31Oisvud3UTdecMZLAii
8knnXAoldVu6Zogy2D5IjjRLbA8nV0bu8safY2orgx56hiXYdUjXyG3yVJaZtcTt
QLEAUZ6I9H1CQba2+WXgxrrJgmeaN6E+vyoBTg1+gMd+B4fO4l2zlxXvo03h+mBu
UrERePwZ/Dh25SeS3P1LauqEK1zeeR/L311y7qAQyL5Wy/0k2Bezl7hvhUp/BI3f
gG63GP7Oyn7WngGfaJWuskbCpDmDYzEvQMC/yyK0FAlYH/1/StIBq7p+LcefjdQ0
y3iC6eCExQE7NtTLRxy7Bp+EGpuzzYzC0lIIcL8Fv+TmmzJ4krHKzNAq1IoxLkCz
Lh4AKTCUxD/7X0MH5SO4hhD4+FqvCwhIGDyxWUcxwDA4np4EXaNCttnwp4fn8deY
gOeIBJ/4+w8ONdUDw8nHB/J5JQ2wC57YgkiABNuHOyolSlTdRxXgjYECsx49XoH6
OieSgliZj/sJULMut9WM+Vlq9gerqgXNX61dK5E5Xt60/fVdFm3nCxeOzrnYfoqi
ElYvzsXjCfOBKpUtNxy7eJIbb7EA5igqvGMEwe1wUezIyFUbpvz1o+9hUjQnA5Z7
kx6ZtabVcgJoDHJCOVzb3CDlJlvFbdPXYn0+1uaxZ83pYhfNx9oI3SaXWNXtj7fK
2xQ8MJxJucLdaRcNwoJVG3RcTs8nazXkXaDnwl5R+HV7OmRhRwmLRG63VxWX41ml
yCIU9SNTj7QAh9rRLLHBwG415GI+7R+k2jnYAUkezBxM/OrZLA8d3IG64DKIV7jw
4xnKdKapjJqlxI/+oSNamM5172DSQLVKvz2XbYyFuIN8kzVUpc+KvcU/ITGkOGVC
Z0JsrqK579PZKsAWKJkeAUnm8JwFY3+JRG3SXxEgSfrv1dsb4cITJYqAkV0r4lKr
blHZ/IKQqdjmpOi04jLAzvTOVK+7oaOLIp8oz0Iy8wrp3Nvwl2I5Yq4fJXeLqVbm
aSQOvwkEiTVXxH6SjBECd93BNKsWBAEyoFQLCMLeub405DaBbsjDyjKkawd/hE8V
b7JZ+Unxo2fvBnk7vkJk/vvF6DzBjMF1DlFy2yzBUAK+ojYBbeV7X18RmrtCGyjl
Ak9kaU0M51v0O/4+77DN3HAZWdCcjhEbNp3CBigjXdt6Ihyz/cr/IB07lIKCkk3G
DPMC1gbzcPdxfy42etCFzbXuloBsp+GyOCttLnu1A5G/pb79zmFgWtLO34inM/Tx
akcU0xf4tyyDBs26zNqV2EpkPNUM+GCKTzVrdIv0xQSI8ejNM7j8GvvqaT2/MUH3
aY2OW1vwgfG2kZiRFkfDfcGOB3tTHNbUZrEwr3hp6BWhrQcdqQymM67PHvAPxxzL
ZtBCOBelrgqzeFJBL8eIPzC9Iapb3h4jazOe3WnHElrhjMd5+iOCm2GstXGpodBs
GK8EIn1RJHIde2Z2zkGTFi/ssT1v9iZuC9QnOrK0wrIFbGuKaalSia6KETtOv/Sj
6uNVMLl8FpI6U79IysBObxg8uT/zfRc3RVmMVJhs6plMMJJZmIGCjkGNAU0agvY3
IYUXhNQSgyyONAib75Lr+65wWCdfqSr7+60bFgn+F+sg8VI+0U1iC2qkL/Eexwru
eI9TkxiPqN7P2CS+XDC8TsaUp1FWwtcYLTj72F7sOtRjwLzhCl7uwi7eSAuT/Udh
3LkcqMOqL5luBy2wnmTVtY0QhpZYWpWHbKeTfMZVFJfMQjdCjDiE66abhFe2nkk0
5z9bP4oDkE1mfxVzYr05sU0m5JdHosSTDEZ89u3kxY9VofjL+3r9Hxvl9+KEUpry
fMAZO7aGiOUOw63AQmjVcI3jibQIfAl3J7Da55ag/TefHAfXx+OCiFTaheVgvEf8
0uECA4021t38Qltr0FGK7XkCIZhyF31AmDsdO6POaGj71MwdKdG2wRUCl7ZNQaBy
cP93nWpEqnRkRkQAoy20YC7HYrp51dEfT8a4Q0hdsyjwLnYvvqRL8PHTrSPJhb1M
qVIqdsDjgAL7CMUuGmsj8+K565z2GooMPPrAmSfpFdDVvu5gvgn/bq7/QVoMQPY3
5otjCMDR5lurnZgkFF0VGJJsTO045NWw2167CK7GJ6+jR8tjn2xl0KQHtOBXr2H8
VQARy1R4ZR7TgrSqEkN7mvDct/gMkS74NO/IOAv9yFZ5lf4oyR5QjrLTdyhfh97X
0H8De+K4FbLYwMz5gfD3mai7PSM7fXkxa0nbcSsnbli2GK/ufekxCK1XPhQuZz4c
F5gJVsWBRk9jjLNItDYEDYsv2qCKScWkcL3G1HnXHrwwxcm1Lr2YdJXPw31DWtEO
ecA2HI7SYSPXLHEw9y9IgApfUTDFXB5isOFJAXaTWswEflfzRZ6bsed+T+lEKDgO
NsbW16LQ7TjRoQ67nNLZJvpTplUCuRbpP6KWqbOKLEdjM0nUZAQLyASF/prGeaPX
NQP7YobP4N0dQQpKcB3IrEbsFnWZ/X1NMycSXIx/aBpZkmNQJfORvzp1DwEK+vXU
ojWPmps52Ywm4xjiJf6pRzFhO+3iLx5xik/fOJEXEVx027CfvUdFxV66tYiF2al6
7Wnsq45kkFTkhKk47nwG8wDZ+gYA+A0sXyWz4khTuh7pq3Rj1Hccw23NIzg6SsmO
iJIZ//fbfCT+8PQnHwf3aM4I57/NSacYw57eeZqfYs8xOOQbJdTpeHBAyRBPZASH
sruSOM1M+PZcuRvNzrZfA1iggsfx2dgbPyMlhopET5VpC1j1l0RZsHOUfc4MqpCV
YQNnbYo+gDvflONEFe6Ta4RkwcSX0T6cthb4QYcqYPvG9X2/lHEuf+M8wLyDP8nM
IpEcmj1v4HqMdwc86BhRdz2G6b25lxa1jv1r7dORf1aVZM5ecS7s4I1ZYMMlCsGf
evhDmb0rk6g0XD06SUAv7CBcXGjOvyq90v1Qsoa22eN+Ds7MaRlQsWwniANSn6Ur
QZV/eN9hxyfecYl1UYP/zPrzvPV4RmI1txqHNkSQYaLuJnjeZH5Sb5UfQerJF+NZ
f6zE7qNFCUBN0/IngIX5VNT9IMk8LXHHd6Uy5UNNolCSEnZyjtK6/P4TbIH+QVcy
31lu1DrvYch0s4Fbh5voFlAr2dC3LjK4N9eEYMpGvZpUKoG24yj+r8a4vrJmVWdH
VF4qW2VrKcZulsjrATMAlIFBMuaJjueCMPVnbL/WjLybNGAi4Fc5kGr/UOBSHh27
4aVWzABprAWvURYwojK8APfODZH8Qi53HNNg7HKZ6rSb04BHTMWd2QOQ3FdHpnov
yRGk4Q1ApcXHZz/GVSSoSR6tuNApUPudqTDo3QVRpX5jQskXinRBoO26bGvD1z6A
xFv+8Tb570ZRpmjWWUkaRmt2W07PSblrhdWBnr5oRdqUBbs957ZfPIUxjhNJrfgJ
bpRGiYDqgEB3/o4xzctTry7ocOT+0dEXqS4jvcG7mEE/gNbnBx9srCDCIWxDNy6f
bOJr6M1mCL4+coEZggY5hezhR2faZtoFa2CDLOz09zUiluDxcrwFrKdgSG8f4aYb
/wLjSovhcsSIONeYb9PIMOtLCoeRWZTJyfXVEgzrrRqKxquFJ7Nb5nRP6/9Jtc5X
V2yKEbxZyuFYHcs3RRVbzrE1Yi5wr1GYsKBkx5l0z9a5qlq/PccU7MvdsM87NmtY
OPh0oMS3jG9O67ZZqDFY8xKDjy++eQbiXP6vpDwf2SwXuLvV2uld1i14JsOXj8dA
7Ebrma2/pGZ4X6Rg38/KJzTDUNU5f7gb5TTVzMWSEwd845rna444mn+CaoPWAHgG
kqY/HihsNJeTH5QJi0a0hFPThyynvbxHelRtOuDKVk4ctAmIdKMpZ4/a5uHIU9+M
tzzePZPpKacDaUaPddmB/ipZOaQ6DPc6aueB5CUev6mky/poYljvNbx/lYpJhL9r
h2Et9mkwU9FQdEfQvi7JC33LlfDJ+WLDlpjIgxysN3baYRaWZvdvTCqa4/QwKVkt
mlYwtf2U5uJa+jHJhg61V6rzlDMKLG9cP16vl9wVMqlwS0+rp4CKQES0su5BAv23
DYXNNliRO9h9I7BojUPJeAf150mpwMzjeVlkGIJaGBoGftrmcFj8shUCekPTvPk0
E4QLp4Cszmu6pShUBkpnIV4zRqDxauVLBBFdBi2O0aW7rrPjq4Qwp1+lm64txZR3
qNtTipMHVcymIPa8DR74eZMvkrzml7UVhPwCjXRaL8JF68qPifqU5QMXxWXbguYI
glF4e9cAXERXcpvCDUYFlJCadbRWTBU4Elc2e0Bt7eY/xTY2v3OMvF9wBMphyPKu
B3DmX4f8K4aB89UI9sFJhVoDXVj02ZEAe/v25HKQtBvSWGu4QjxAxxDr52s3PQM5
YUEnpYL4vUReKjMhHETJG1lmINHKHkgXrAnY6pslvee4x6ZYZ7BSUhHM7JyIAI2h
3FVJmP4CnsTv5yJCOKpWwGpx+zlmQmYX/lz1zEn1WJlB1Pm/v7wOREUA7NKhjn/L
gSuh7GiQkM+/+PKh4KGCBOZiuP5UQ/ZwNsWJfAMchq+8+KkarhabdqaVaDw2Nq+x
3krcvGgv/UINoUvg11uFm8PGse8PIVkIczr4sNNFj+Oqa+ULfTp4k4zCEDwZpg5o
OAXmsUAlFcbgRd1GP2hkX5kzXvyS9YKD46qQd+73cZM7uYj5BFUsxNFUjCYnYOFP
GmkNyXKPw2zNc+N9sT0cVAf+o3Oqr6ZEQwNqSqDhghcHev84ap/VaD+iA3Z++WR4
+ZJAF1zEoFm4Ww94/Gf1TGxllojxjTGtzTE8bmkdDEaDnDOBsioguXKBvz6eqfOr
G7w/TRBR23qxM+5VnOO7b720fobbukk5dVgZwJRoFAuH6JlEHRFQHlVGBUaEeFnh
pso3OBfvcOvu3K17K3ai1OHrLm7Tl3g+zsN1GR5Syj3/Ow9iRU6VVFu4VOqrxv8b
YLnc8XVY6+sq4sz9Ahn2cVVzSPdHxmzl1yFZj4SwtyogXKcrVNCvYLGd4UXlGQbt
OL9rAOJH3cFzhqthT/XrSa5anNqXNSSbp84uUI8z21nZvkTI8R8JvgASL/vVsXnh
reOBHrroq8yhAtGKENP2iho5ZSubZ0E95tRWcYmjpsvSYjExUDGx5JfXS6LeArg2
hQ+92zQYBsAZz328pQKMPU2OssO7fwRNvOwbnuR4JBYNrujs2aYWsmoNjeSqK8ss
95om7seB76/+ZDzv6b2i4QEpydhmQU0fD8uIMOWLzNP6fRKySEW7+l7eEvkocyPc
l+fWzkZglUmEtwe93JUTjomnXqfhy0NhI5vy1ceb8XaI7DBwGpDv+8SkJUEKMNuf
icliPdNAuL0JesWCxkTUN1+YXjY1o2DRWMEbQ7LPNN88mUO8iewjjIEn0iYrw4o9
YROwV5RBK9MWv5iGS3TrPV1P/kroHeBsADWRwDWkLwXneuFwpT/JnJJbHpkmfnrB
fJdrjhr17knEOkOyivypX94UryOgZqE0/5iTSqhOvkqMMAHFtG+cLid+sD2UaIgh
V2KsOJx8W2uoRQK8i1/uLmhKu9apbdUgMuprvZk+C5iWhzQvenbHgB0LA9Vmfakt
ADQfN9fQdUbfKffJ4MQ49VhscpwVKwPPTok8WUI/KkafIuxqySOjmUOY2MdJoXNj
RHWBySN69khWe0g7FESC8eZIomknEMYNK1fozXSVHpXFYGfeYOG28H+EwI6Cz5iq
jfWwHpZPqa3iBXB1NMsCuQ/8Yfv9au71HeVv0S+3XX2kEyXsjh6JoioHopzns0ef
w6aZwZ8C6Hwa8zpCAjEC7uCRQFBkR/0vxSRGkwREvzg1z4NKtQo92tL1Gusiz7rZ
fK6foPp2KCWQHgtX/fLxPSHvwSObBXXkWHehp+YziOIX1nbb/wz4mR8e+N4H4qnp
DzAiHCY6KMaNedWYIfBl8xBTEnbioZlceMTAVn7M9cOQ9vqFqMSLJBo93zCVlFmh
mIk0hhztH7PVArzA8nHEiKwAulB3P/IY7JFYxzdHnK4DbZPK0X1le4zZ83HHWU8P
SYwyN3RwuDmclT82oXTDTY83PKBydPttNRL0gF8imRn2oTWorCukS4+IUEODG8yR
eMSLsEc++2cKTPjkEnhMoozwL8ip+VoLMcJmhvdqYxFMCGpxjKsP/1SHoZg+b9lO
+3UldhO4lW2BhCp6bDHlOra6asURamgs2XJoXvPMW6GtOp8Ic/Uvt/BSJpxWMcea
iZi9BoqrTN3lUD/GTJUUZgE9zODZ21CpM6YIvgY8TuFdoPG2EkpZ8VwX2BcL7CGB
0+IoelepvjDf/pmxGzHJVha0go8ZYkNA6im7b22UGuolWWrcx+qAiaQY5BExPSEv
tPjZq/lhaHwczPgHaIT0/pYCzb5RHvaqsqwQVgPIAkSvcz6dbzw28QN29Kei5OPM
xHvw4YGPSJPKVh8EIqOEbHn/fgcpcGnAJ2J83GeTLOPiwXuPcnsExpeCwEm4pFSM
fIyYIm6ezIu9AGu0fyeza+WSXm7ZHieHD/G5Jagz7+M/awiqg31LaWgLzrvZf388
DO1MJjb6O/OwBnonVGdVLHlePlBwcoNBkUCENnCuvqZUQHl/D+LdH5a2pbxlPwMn
YjQLjxm3wwCatR/QjvNIEZAMoVdkkw7rY4Cfx0oZQGfj92JNYMtsIHEOpyQ7vjMY
H8b1FtBsnka5R5fMGlicK6ZE+SNpERshS15woaVM78hKdMVfJFXw7BiLNBSLMyTr
5tlUSAoNrKbuRCueFU4P++TWpgopiiL8rCOKk+kAqsuadkAHbXQbrn6zK/19THk7
7OmeXY7WHfiebeN5p8ogAkgDQMFPmrI/vOahM+6VDKVZXAq28YdGDWeasJ0CeC2v
hRdW++NEkc2wDUbpeSva43ewazdyPECaC9EW0AiufbBX59V2UEgbfQa1hG+ZYM1+
vLWRk15F1hTbMuaWDajJ+uWa5s4ip/LiF92Rwuvm3cEMZcr1Znjh1O+3CrXDgi11
lstyiOXYfn23oqsSPN2RWrcVdgu/c7LjUUslCAQGwAymPtrFGkncHlAspW4h3dKQ
diivitH+8TsOoB1jPTg+8zbPLcoPdnzFGthPsbD2GQQCYIA9pk3vAh4FSuCWVvJq
ylqm1WL4GSJfMZ5gn+PYisR1oiBBQ8xy5HTfu8f0Eek4hYszRg7Sui6/Pp8NmssQ
HMN3QYPMNzWSgwfNxsg1OvMJWouO4ptPkI/qtc8qlAgPzsJR9NY2vGN39zwRXix7
48Wro4wmAdWxoI9yMjHzvnjA7gp/QCTzPRMk1PaTNdKfUoSwIW3fUIkWaDnf5ChF
3dSQU6IDGJxloLeR7MIRmOgmAsnfm2X2xlWLW5sdEGaRqmW2/ZFLlCfvdG5zdXXU
+d/ermZdJcLGSmOe5+GDubLvQfn5sgB6rjcJ+aAgCVp6CT1qEidIhMoM5hwTDPUL
8xDO+n0g7Tn837wN5Ip1gFTXyHeQjAeenH9lNJTxeVRfwjj3PhCiskBGunC89gCM
HU3TJflo52a04A12AZYmtalbdkCWAwbhu7OT7Pd3JZafU08kiIyeBZpnLbv4OMYc
Au8kd0nGKPzy2vQ34axukX6ZMPooOtKIqtpZksUBf/HVVLUalI3q6BuP9WKdrDpO
bV3nCYN3zlABdZh1pT1jAGju713LCB3x80c8BEt9DDdTpIwdilKFkAUGYJUDrt/L
/6kD/CezJFNTQY6RPJiXTpFTGeltH7W8sCfuJVMrJgCahpLzdvzT/6TkPhbhWGCN
OZKEGwe73VkY8xWr8ZWy1N0wgujx+dG7WAl+2SWDA1QViPc49OkrKkK0cUMsfCzV
GYVAhlSIDDGDn5k41DXfZC9zskAQOkNbb0Gt41smdtcG5bOQNabWxKK02fph10lw
fNIzuhj7XZtK/M310Wq4bnwCVvw0NTZ5cVrWgyDOhFSfSKIShTC/NezqBjrSVgVe
UszIA9m8WdapZ4U4DRueOpeJlSHLgCAxxkMYrx0nOw019novzUQCSXV+uGAV+tQs
Py8G7HuOU2f/4nCRK+8ScaAxEes3gDVTCIymCHf9+hBPVGCW18zYV99Ih9Uwe5M1
hdjtAyYSpuUmW0GuY+MKGAHlXIhDl4X9RAfuj/plWxekpXPj69kObs+KzYk5a0SR
iaOJaJDzeP8sIbVscP4uq66YBmmdkFUJ3/+sZI0DBwK1RVxRVgKl2R/QlpHek6q5
i56WD6YsXoRw/kzv75RCBGOoBDprFwGb5apvYaT9E2Oh6KscHLTGcJolZYIuF8vh
PFYZPMry+GEJSCR7yzxxe4gzis0DwgpygozzqrlbJQFwwwtuPzb09ea8yRqojLm0
gd/fXqKwIetGAW6LC4M/VQWoApCuYiulmW/T+Lto8lrVF46m4K8FD3uPIPVDiYbN
B4IgLytQaS3KCDJop4O1SAA3IVtWqJKvHaPr3UVj5wVRozj3XTWZEK1YQKcuOg/y
uUMXXs81PerVLt7D6QfaZOIgbWmkjCSt/RUiBxPSKKMMX94VKsTurXeszV0heLSD
BrSLoJCjkVGHqGwWh1nCQ+6wUhZAzq1m+bIhZPPaEM3Le2+3Xconqs9rJ71JwkTs
w5C8oDn7k33gxHGH4/W7u2hiTjwD5rYQgQ+zHY6N+cewTSMZxpgOd3mo3vlwwY0o
jGzbR7Q//OrH6h32CAhCAh8SGvm9nzWCv/MfxmuF/bsCS+Z3ywsLJDewG6qnovbC
0Zby6JB5YzCO16BnQx5bnUkLwh7Hc6EpTC5zALVvPGvbKYPiFr7t/3/KUP7prluZ
o/cJB+9q9ycNk5Cy4yyppTEJXGHWdlW67wx+JS/S9D5vwa0MRUo8L2FlxX65lB1i
G8KekYsRvbOYQr5Tk0ntIw57Pjjkl/YgMLjEqH9/MzHinSa0BplXq7HrbxJFrDBE
imzdxkBDhSXilSwUNl/VHrjIsZEBnQyEgYT5TrNwpf/7XmP33VAnvBqfe3Bsyg1G
n272mppMlPWbRDWirQJ8A5IX+aI3awsy/DCf9A8Tkn4YoiJ7KEhHTDtOjdWiv3id
Iq9teTaoUNufmWaalZ1G44lRQdH4ejmEbCYEmVTGiIOWVouMicbQwsxoFnZFeq5m
AGEnLjPIafInIFWgRF2xG0J1eXx+15u6lpj7jHFxjPrSMDMnkuERwlUdgnHNy1nA
UoGO9O8oyV1Hcu/HR3P5+dm1roNly9ci88WzuSA+rz6eQCNl7L9NkQ6wvhWd2dSS
WaQhZduRjyyS5LXP68231PqnCunFAFWDH91CbjBIdDr/PTSJTaO+BeE08ZBgc/QQ
svGQYBUQimb2SfehGZswoFkmBPPI1m8rbZQRWtPxsNEpYfzupHkh216ktuv/Oi40
PRC/Emowvpxy2TWl3EqlrIovvxMd6ZG0KRRXjsZE7tjqoucz06Vlt18jPZQhOR8b
GxWSpiW3KOdOVpqJcxaunTyfmyYnTssVjV1kGo5lxbSOWFPrDVFZMWUn/wixd5+Z
HKMGEcWzE6tYpqNZDB9cIrDeaK82fEzHGdp3WAA+UqYGWgEz0ODY+z3nu3CUmIWS
pTYszL4tHIJhmGW2p6U4VF89NWcRpYd4fHF0krOPAtCUeYAJAg+0UGTv00BYY3ne
wq7uEpjpSw38cE2prLO2zUsCOGVuvc9L1JqC2kFECqXCJ7LyQ2/HcMrhqwjRWmCG
puMB4JRNuxawZLhfCsVvOyqnOyt2sk0bcdUT/dUFcwQSMoSislJJOOBne0hB9MGi
4mCnKvlp6s5bWGHC01Xc6qd5m02S86h/B2f1wSdas3SfcnnXTieh6gYVi1eMOaR8
b2K0xU/23r1PHML6qIo6FJSf+1Zip7iCwAE01mJVEYfs8J7CwnxDc5JQmctFoLwa
HK3KdWmqVkFAhzIPQ1VxvCqbEQBPCuWwJ6nPk60EGsMwqZpenmvbG++Q6y04o3Cd
+F3Xf6qM+ctCYp6bcGhRS7YIQN/lyn87CvRnWR5aH6Qu1q2dOkSWiFVnONp0WwL1
1jW/9szi4OAWtJYGvS0yYPq7gz5lf7RYLPUjLP1m1a3hIt+bByES8o95ReJF6Bg2
ZqPsjkCUdxvbaIxQMWUtbtBt6CVZ1bzPuP/tL9hhhv9VPf/YbskuL2L0/wc3t/S9
mUpYKR9Iw5BvcMJPcQna3RtGhX6xuwCFdJAwG4xGrYqhLRrFKe4qHAwFOrE5CDBF
/1ewHiIOkUG3zQSs3tW18WKLsrZ3C92C8NcMrHR3e+8tIaljbxQL7QTgYPaEmkoo
4DEpktgJ3oKeMFU9yTrscLNaCy8nAOw08Rnv2fi3wOtabfTrwxg+l6R0n/YlvN8J
BPwr++OLvDCA48mMvA9whg1pey83OB4n4acXrTrJcZkvZMdWtes6o0pzCYLQKj3l
LZNpc4umQRgKVh83NM1p9BhdjSwy2OtmVBt0cJwrJymimXVVX6Le8O2G3I6/AQvR
zmkFV9W7aM4f0j7jIlMV23lnxjoB9VpvhnIoOu0fEHK1pmwGUh3PVd2jLV99GtYn
mo2tMT5NPYog5CxZZ//Qqt1bwiCOVrNoPhTGclXQIozTNtivbF/ouYkQdTVYkyMF
C/eYJ15GRGh9LHkzWA9e2VKfIlDSX4y/FQhEcWa3z4KXJeqR2Cv/ff1xJcHokUOs
fDCwKcH7rQF5p2tinaXRT3PNHD9tCRJTKGoYhXb2lKu/APr23L38idJ15OL63qiy
A+3QIOyzVsh5tMWlPLgBRZFwNf5l7KXNh4QORJyCwDrgN8npj9CFGi4cXHD+QDac
raKJOK8qcRN/izfzJchbgO6dWXTeImIwfXIouYMdUj1zkpqnFey3uFX3hwHEiBQX
T/NPp1fYx3OF592stl/Q77ScZbHdxe+6tQRmaLjFdfzsv3fFnbHZSGcNY3OfJ/xK
E93GBq43dRTMKHSv7zsg8X+C3vJSCJWsr+IIgls5M09wNn2mhegJSoptq8Wavy/h
8axaWElfGvuz8c7gRjWF7pesHRoi0J+ctwSkPtqzgm26Zki03e7M4ErhIvTZTLDT
hUW8VBS7uGIy9+7sK7cyWPOToAqum0+FTIxDWu7/r4PzaSiyyDP7hGVMRcAPk5DJ
OWONzlmPSYPs9PY6LuRsN6h3vqrAodAWRW9QHa4YOgqtj+rL1n0M3gFAS7wytCmm
zjALWV+1v5e690Y61dM5UMcIHw4L3Ik/HYbugLz1lkaKSCVAp4TwXKGA0cOj/Yly
Of0DFlFeRUdeVZTLDMPsnjVIPCxkPuqABiwEn8rSorl0gol3b3SqoP++NJlkFJwo
LYo/PVCHPfYAywNDI39swqtS1hVR7Cz2s60fOT4b4w3CBk9k1pNdSljjuQNun44i
cHqrAhbvMCAJ3ouWunaNKOQhAUsmhKu6EvS7iYiLNDm48afGMpPvPO/fcec1Tqba
0Wie/s80IllfkXYU7gE2qwzHxGqhUxZIeKNH/T+2F6cUio5mmNVALShv7O41MPMu
GeKUWgVG1jfUPyXS6PDlwxXpq5stSi+KPgZ/5e2oaMLHiCo1ySRtlGbjRymOHO3T
dWjycVIO94JDo7R9jDAH1P0av8UoyLJeowLKKpj0HzV7El9CqzX0x5X09tGB21Ez
0G661NiGjV8puSa9T0zv8Ti9MDCUl+2UvyXkSeDEKA0fnf2wVbfC9wcuqt5iFEPp
hkNbizqs2BasnotuiiJJWRJqG+bo8CwYqkjo87bQzi8vKpsBP5xXFym/020XqXfn
kLtIrnNQMpk1gAhDLU15G4Yx57vK9UQ3Adr076LdBdGB/F9jvKkcOJqUrKmjLlME
Y/5s5MUSNausTQGFmRHUuKGHS/2ewHj4gUyRjlhqGSueP2O4WIPhPmT+GyoVBeSp
bks57OSU7koctetAkvjLNV2BamUz86+e5X9GUjy3ipWdFAFFVkbDuulVXZgSSOyR
TeDzYnu9YpqBxffMQup32yWcQtzAQIalD9F8XUgH02FqiYN9yZ/2F4O4J/6gEV6r
xfZBrxf65uHrV0kunvw2OOehuVOeHbEvOwBrPU6NobKuwq/U9QUk5Of/RmY4KpWS
4GoqSYeokXOnhW87UdQOzrIEvJKUfKa0x8cGxSRrw53wrnhOhHUbYry8E26mxOFP
y+LJZm00M3K2dhV7stYro4QHx/hM0WqLy+2o1Ugt5mJJLLnRHliRfMhN7LKzYb9/
TTKeFDSp7f5jPpyyigSuYo5X9vgRAd94cUOufNpfOMbdz/2MFHuYWhLZLdlllml0
xZbf5daCEzGlGKT3AjudL16n/ZZ4JKgiOWER4DyqSNpcP7ZradTrkdcrZ4FXxrby
ltUJh785KQPhlq7WA/JRLWHLq6fK4P8wES8XL0jh7PA0dEQsnKFzd575F/PZ6dzf
l41t31x+sgVtxA2dGWezr5DW9Yq+y+cFho4txOArGW4ksarwZSKxOX1ywgXWKuTY
5jMCNoC3LNImJJLoX2tEjiMdC3ACuEWjM5sBhrbT48KYi9LLko8iMpRIG/V1SFMz
DgUzaYc1DcvI/fvJrjE0QmCBGJHs9hd/ZGF5SK3vMQiNALmAdp60xUN0M3X19eyr
g4q2YAbehNz1WqVwwuULtGH7Mrmld/VwuEx7S4goXG+6GkuWlGGgThWYzI2Dz+H8
Wy/Q0CGo99QJjkYa/0jnZvCtvD3UEEhwxLZY6Gne5U5iIePNa/qgVYChPxIsDry2
iuk5QNwoK04jL/rkqEGQxTAjTkXL8KbT+9kea2g6GdUJSp+/0a0PmqoS34A8c65k
KGzjXRY5QR8eZNwAtqnKf9WLuSRL4BT3zwPvzEI+qwLPcVWd3MY7Zzd5hfrawhVH
ql6NWYxQ3EIB8lNuLpxujpuGa+UEhJrNGVXR4GkfflC8yDLLDqoIHk0pvSLbeZbd
9lNpyxAXFSI/FplFIygbbNjApdMnskQD+5l04jHZjcomzJ2PxBUD+Lm3bUZ7pyo1
hwQb/I6PTGgU1zBY0q8I2EClaTZFUO2OWCaKk5HXCjBOfFMsBQ27JRrcn+6pmvoL
CVS4d+FJHmUADjXaSZzBMPSFfzmEP6Yp73bDz/866HPe2tKKFHb3RLai0ZCF2/hD
tlYeATeh782K4gJtPp8yz1zyBTI1GHT+mXtueE1qmLXRZKl1Jld8KRVChb/OIuHB
FfUH+e9qJLMIsK1J1OuNARWowu7/N1m1IDEaaqt6qZ/4rZJLcPnhi+TCSEj1w0Zc
Jtc2cfymVYhQ82otgWm+m7JvhaxRUAwbEfTjvZhoM7sR83CMB8r638PSlC00lj7H
Sg6+wPV5rHg+2WMHPrUgA0afvtr9Ohu9h5iDZ5Lj7rQJUHO9lR0USl4VJDZFyRA6
XQTaezDY0wuoo1jL2zLbUAoVZvx4DYrRypibxkQsfzUfJU8FXRfGhTwCilAaTy9n
3UvGXCw703wcn7h0sTkuJy257yTX4Q5gp5YSgZiq8PvtHoKbnHsTeix0w8Dz+AV7
ACO4Xe87tHXuIvtHKR4hHJvT1vEKK77shyyAaNRph1R0HyeKsASotoyYddKnG8+V
P6sQPc8vwsxXyu5UFUo6PhExI2vfpdMuokTt8u3hqYpllzjatv9Kf+TkSsbp0BAy
y3mrMgrfW2+UgIjo8qomw2t3suK1h5MmGCeWlSeIvCsNgo3VERDMbVxW9xkPzL9E
HK0ShELnuuk0EmiRGLsxNxHRkhFj+0yMLy5R+BXCzCZT0WNjqMH1K+DKkK5u9xX+
IKuXgYMbCAuXAz03UmXoK9mLHAj6dtxD2slDhzdoDk9V6/hr/D2c3R0nZzgnHIKS
YXkudcW573S1pHQQ9MjwsWpRQLBfue/Y7UYIoVGMif1Y77VXNzrmUFfWLXm0no+G
U3Xh6Bz45Qy43e4AHKQ0zuGEQ9YJYekutMswNkxOsWcrs5JXyuBoGayDHL/3GrV+
IZQtvQnZ9Teo8eWAGtCDUOOUa4SKNgGm1jmoaMfaRIKfleeq08lOZP9fJHZgnAuC
yeTeJBRxkUI9IYm20rR1lWxbZdfNHQRDtt8Hkfx5xdKzVXJTf1V03/vqM/GDPkF6
jw9N5mYavCXcmASFzfbL8U+JFPCQB/OACxw7TTfgrttt82rL8XtlKM0aLm/Z2BxQ
IjuOYsj2vTdzGR0ToaW1Ll/NaaNnCwEeQDtvXS3DW2+GJkGOmJQYCk6t+27ig9tb
h1r/8xuHnRAhhIud/dCF+9p0tAsG0QKf/bEfIcontOvxpNYK2PChVY9I/2E28M8G
9Vvu+OSYCE8BZI4liTrBDusfONXmgxMDPk++d5grxagbO+xM8BykmMnypeZV2NQV
5uPNM+x/UvF3GJUqj85GJAdKJNtG9ypSnYqgEZ9Tru4q6Up0vkSGx7xxEuS+Eo9W
4SzjCSx7HQmn3ITgER/4g6y0ezIieIkAL6d79z3EnIuNS8YsS+D4xTm6FxXxIxmb
r/YVGYCnJMBI4GRnR0d6JcryDfodE7dYGpUaAnR481Zjo+M1+91DdgS6gqg3oLwJ
3AjapiyUEj7HDNbhdA4bp+IX7Hxm5d6XeRO5kf1Ob5rFryNKjRS59NzqpMU9tinA
n+5cc4tdqMc1tPyVxahrnOa1WIbyaeHHhGMDi8iHzqOsSe66IGAXFHuEQtrMpTIg
mYONidqssRIti//W+OJpVZaScewMRW/9DI2WiT9Majy5A4+VQfSVTM1huuYus/yN
biAitaiJFUU7ezHEA2RvTF6W3dFjA/mi/Pzfuk9ZrUWgHvOfoZ8NK2wNpHe4mIby
GgLW5hpz7p6yi8xxvlEEH8H1IbangjUR9RC6GXi8CXimZGNoZHS3gH4hMBq2EgMA
HeGsS8bZkS4wkctPMRWWlG1/H2YFj7Ilf2ZxYHxvVvWy6e1kKU/VhfsmYXhrpx89
umLjZEKKAdJuqFcGLAbZU0zQ3DO5xhwmWqJNsLUQp6mJyTjT4HEvnTNpo/T/FwsK
IplVr9CXQapYKKBVpWw2Wg+8Vyttj8CW14TYlpAAGoo/EKPj7jWQd+mAx8bmVod0
trM72XeLC48iFJusOCsW4UOfMlpAPOPOO/lQSPRso8+rzQica72gNFWcXmdKQi6b
79dvtH4dACO4fgCkehgOOJnC1nfqgnwUduedcPyrF9Yz2Yr8BUDz9T1BDUvuSOXJ
2ZtN/lp8VNs+AnEFwnCa03e1W5MTYeTpVAGYl6ROpScv5cUU2RHFopRXQFoTZa8V
lOy6Y7akaT+oOS8+7wMeX2b8xLS3aJIqX5pdso8oxw2jluDbJZgLdPaxu4PBWvbA
etRFkDFt2OhxfFWrdGN0jxqSOLKJCY4qbpykZIdBt2/cpSVKkQ3Y/FjjFd1GecH1
pNbWe9jmQRhULcr8IZxSxGfPe4J5jibg1t+ysrS4H1vaIbTjkRQHfwRpt9dDku8H
IB2ZNzPz1hLYfCmWSS/GgnPqyhBEsxBSEEL/CFQ4Ph7jONddaNxq2dmMfjMgJYEB
C88rKo/SsEi1v+vf+OKYS4pK8WJ6FYYNFEcPGpUUFEHu5yxD26h4JVnthR7A3O7e
+RoUIeV3HLux8YAJ0bWk0kjUXYJsiwBHfDeqkPWPMB5PRXo0E0ee2nH0hH1ZKYoA
BxGlNmy2ENINy8SYZrOhrRk+FIxUq6/BHKuQC4kCUbK/j3Ct9FCVRgMiPPhqTy0m
eSD9qDW7JBpEUrMECs6faHDaicVecnFKhBKoimOHHpikVGoawR0u7fwk1w8Isoqh
ku2mgcYi5c0ApqJA518Z+wndND3jQERiyA4xs4CBtfPKqcoRyEPYRZOScQhj3v2A
1nH4h57ni7rlYlc6+WHDO6l+TstCLyrwJfsvl5aK63GJqCAS5YoDwbJBnqs2Gq48
zMyr1XQxk2v03CbutVyl/YRI0baEP5kBcE3HL/EY5K+7KAbeDq9mgUQrUEG8QwBL
kdJBOEeUoWceLTk5Ly+TelJYKaUe9zZEw4KLgeN5VPpZPsuNqXC2v/MRMBWAje7i
BBRjnlfWEpwTPCJS6ywJcMmIbrpxtWRBxN7DqzpcX0nlWfOcf67LkU6uCLtmDTMy
YkW9JqYKOowWjmbUYexUc0CIzskJPLAHmfINsCP3QtzJaCDxL0tpHYLr+UQ1vxDs
9WpzJc8cZXNcRMavsWNTCi9aKiZLQd78Os74rRoaA4veC8aJnQHGHllxwO6NwO/Q
sQk5fJilmELpUpfuQ2FIpDo+BTHHM4+mzcRYqk0BjWowuNB8e/P5mdA5zLG7Ael1
64rMVG18KxGKFR1079/QfpieiSN33pUFxbF7eOnDlNsYflUnqeCavOtV0VqUViYJ
k3gnMRt4AkHYC0oNxDLrkx246YDFPmtUoGFl+IpkDLIFBo9F5edrh7N+KCUXCG17
7d9DirbmRtfO2d4g7kU7AvofL+AKjB+jS6w5blElYZkxPgBaWUQNtIMZ5mLA+OAY
9g62zns+0ymI5rUGUaXkB38rg4iSLyyYUUj6tw5tmk3HTtToi+3Xe2Gs4fC3B5fW
u4ZTqDdICKlmYhYdLvSklpl7VU2wAfEn+t2Ygf1vavc9G1jdQY1VmQCnK4oI9wyJ
C9ZO+pzyvzTJPbBBNivwsbPGY++rYZ9xYTWjL6l62Zk6KvUFuPnYGVQBT9boM2FX
ZOUg1H4ql47L7zXhzkbJroOy+P4d6gc+VhqeImCpZPLtX/EM40E0Fp3BS95doQyR
lY6uGrc5sjyBERI0L39asRHaPYmccdaqz+5W8x1dtPegFsFf+d+bwIGYglj4tJam
F3fB9JXIcB5HLBlUVbJoaj2T5XbQOyxmByTWS0aA5hgJ/CDA3D70GzntA5MqBGXR
maNStcl7YS4BULVkTsQWepOeihRgf/PMTbZJWgJTH+qoPisresliEgHYjXViF5w5
Z7cRKqxO4to/qFx02oGhmTL1/PP1yCfwzbfZZZG0n7szSHrkZdbqM6dU74PPGlr7
OVh9zCqCCGTGoQsi9hZRPPravGcplHE6twag2AsNt4mLne2RSz6Gvu0nVJLLmoS5
hxKQB525NP5YktghB+uDUKqN8EmrCpKhhBJ6Rs/pIZI4UHwedLnNtk2eZgEaZ1tB
9j7a6pdhP67JER83iesvM3osqJclPpSx4uX87WFDeelA2Igy3mrJSaVJoXSoiMGE
QASCn1Ru4nUQOCHYkuc+qvMjemn1wc4/W8zaCsyiNetCO4jX7bKl09Cs41/CvfKY
jcSlrG0Js/e7hoQunLZj6okm/w8/Z/QHTGHl+jA0PzeU8fVa9hCbsluSjzceqVfp
ABjrpRo2aearUV1kfe4VHCSOqYKmeXOKO6WdSbDPw8G4evqEi2Y2MVH2mjxavsat
3jGXT6+1KoURCpG06CjXGNgLGdJMoMye5a7BZr98nskyAaNrbxoqmFEm86Yc+4h+
8pal0YCAHLWTN8jegcQzjCNFZNojW80eJ4s7X++FMYm93vwGBjfB3ml7a/ElqMnC
27AUmhNfpnxA9ypT4x7V9P0xpWz+0LTC4o7iMKwgN32W8yo9em52DUHF8rxJulNO
+8r1AGfEhfc8iOTQ51EQQO96wET+0B/KLoF85uJoxf7tlr1RexuQcHl7Ee6lO5fs
WiP48EZFKY7x98Q8tvoypFgFPf9SpjkXVO1JCOdPmyDa6UPPucRK4qbDU/C4yV8c
nZLcOgibJGvLWql3kQXzSlIoFsG/uDW3AZT+C9d7vlxLRW+Dr+Bo/S33FrRM0Y0g
u+Qdv/Y8k0Vib7xFA+2n2KAdvFcS2qFGH+KVlemvXIhsawcSSGrV1G2kWre5SnT6
S6ogf3UT+IMoG5jFfWsEsc0YfLJfL4WeHWLWdLFFHCQJ/cQ1ul5S9GIHiX4k3Gdn
ZQQANJtR2F7ukqZjaUuOgTmiPjf2pLBkGcWJx2QsV2Fj6DGxqvDMdtDcKcRiLEHk
3PIcVXILFQK5LX9OZUv+rEFFfKvoKVP2cY/p0vPOefAyjL1HtHj6lwSiU0tv2sIh
FRNSPPLqaqrkR778+yV+xtp4hg1cr10wk5ZfItf1cvTn95Zvhud6piM16nUf+Lli
6Qh5WcdP466FqYGnSH524Mu2zybBB1AtBs9nyIpQE8fNaja2SmGcGJGrvFCkcnEs
0mCalF19UP8KxzK2SvvXPofjDjh/zUY/Q3ZlupPvarhljHQobdVosaUarr/8YuFk
5hSAArLdsY+BMadcnpB59pd9eNR/+eFnBo6EycEUW90ZVmJqukztUto8kFMzAfhG
vXStIzm9kW5Q4UVVazoFhwk8s7J7kgSBW8WuzMDsUnYA/FR7SlKsmuOZoMtIBZdO
n9yUDZeDhFwFYUKmDg1UIazYqXv0sl7onj8Ml8P6ENJt2WhndfgiPD2rzIFZhAWt
YpnuyqeUQs0GhkgGZzaY1IwMgxusg6g4t3l1EGM9q5fO2l0oyPgV+SLmLT0dxU+T
FGi3MOWppBMyWEItOZVX9LI181F2/7xRH1B02dkmcCEI1fXxylOYxuZqLuEXeC8F
IwfDTDPmXG1MCMZcZRfDw/TpFtblQF8QkydiqptVegEO/tNyybqWTB0hlejteFAS
YWwrtn4CjcNYZtw8BvPll9OOMjozr1JMsKHZcQedQUwrZZtauehoUqRVq7H8lbI8
OzxaHEXl+4OykmX4k4zsefhsjwA7ck0rZW/GbefKElKDGK9NkgqtkfYVsQNH8ogD
ffsKNHbhr4qbCUv2Z9IGvvg/xVPpjruMrE3V2uOLeHp3azPErMorKAKTFHPPBnzb
R/Y3hjsixAmGYb3NUXiVuuY0cccvURCBrFmwPBEhWINkpFC0D40iHqlDzWoiraCB
NQaSJazzos9OtMHOP3f+zxcrhxSKTCzVC26IQkBvJKVqT+NKWNoBQJPIHbE3hTMj
4Xr/MQFZK3pcaCrzogVwq1ThvNrxexJ8zcYfnI9byzTmUvVbua707y0xHSWjQaPT
vgSGIW947lalQSebYfH9RJifjNhaMocpaWGSCwbN7UpctUGmp9EIfEPzykpurJyz
/GGZfMhXTGiRdF5BHV/VJES5kmzTuNfdS+FshYjY5PllGzXytXQaPpjlMGHQXiVY
Ufrhnla4+Q7CGbyEDVLE7nOJufEo89uQOKQ0CPVqhr+pIPOdYRy3Y1gPNY88+R6h
oYdGwg8ig2iJ6zrUv/4Ntxmxsm09r7YwPp6xWUqDJpF2v6Bbv1RFvKVYbZczTijN
binilzOB313LdXXwk3ZgFEihTB73aEvmQF/yRY+ikVcOkvVAcEq5jryk5Ji7KUoR
AtxDb2QunycmgF8B3AyJFHHSiTAZh0Yt7EW0g8fwO2JEVBngn6VOIQEG2NtqTcKH
Z1mTM0Wz15xduy3qQO1rgbQlf6Ad4wn1/Kw6hUnNavBErEGVXAmkxZKg6x1tEw2Q
haA5nHiagOemDI91p0HtjiocZxqp62P2XN9gzRY+rTh6rFNT284uWX52EWm2r6k1
eM6emKvvhpVclgfL8Zd9Qyo9eM3/Ql7CVuPr/hvVRb8fCg6rLIFLpNytLTRWQuPg
BwNrrM5R2SXmBMDGwObaMK3FEVjNcPv5uk4SPsLdhMVeqm2pcsJm07r9DPS7QKuP
iTmkA5QygMVOmEiWWSGs2Ako1o8hKwsGzOZz3Wu9ufNZ4lLVy83reg+lnYnri/o0
i01OwIAgyIDm30K47qFtnxPRd7xa+onJEt1aQceXX7csnMxOo+d1IHEWC42mRxA7
DJpjwwI0rlWbQ9ny3TWmhOq+e/41hfPU4E+ov/fDHEo8/68lcA1ww437s9+WrDVr
q3r09w+RtykbvxJmX4Z73IbenJuSfEjtTBkL+9aMINuB5JouPSMB+dWXERwIG/G6
3UjZhw1Y9Tnr/zt0Zq9a1SQvpNUbJazg5cEa/d6TQA9CDx3l02yLFMlIQtPqfVPU
rkj+sS1fPPQteLYGsuwMsXPnrfJS6ktn2qXO1N2jvwGoGzTxNGqpBN/OUSe0k1gW
/GQfM0vZkYLd8EniwlUtwNn880odpJVmr+dCcfD1RtrtfGMLdSgNZvAPcUQ/gN2P
ZGE16Ud9zsLiw4althU7QuYk3FzdFfV1+IvZcKkFD0Dh+jI7Rmr+jhQLeSBr6vUX
lZ1sxUyZWNkfXaMPxPCbVzs4iXNCBkjq4DKz+dmDww90vmhLK0Xm9T/qylxl7huh
ftR8R8rdQKJRhr2Zkdkud/iUZc6l/KWkTYpfXMgSjPIRQlNPkH1+PVkPY1OdmC94
cLpr1GPVrlKtVeZAo937YzZ5+dtzcoksXLOQ9NtkKWnzlHpgw4CCE/AcZspo5ASN
evK8V4fXVWf7Dx3cR16PwE6oXSFXl3ual/tTaN1vmZ6JET0/Nqx9VzKE5x2pJN7M
b9LPpjkh5kNFXdH0/nxA/q8tiFjwjpSrVqX06BU3ZTFjVXqM/fe780YMuAbSVc6p
+3HBu70/egDde4LG26+B/pt3p0az3gPpEspPMgnr8hyI9f1HYcpy01skqQSjfIK0
7QAHh5UDrgweMs+Z3az98Mpa4JeAVOYbc7jHhUk32ES4QHYD43xaVFzlR4azdWaS
7yX5Ra+pcpHDnwdzFHe7A0JNmf1mK6b/0YF419di+apD3mOG+/zA6XA2uFhvPAfv
IICx8rwRLgUtfcKtI0/JTlwa8Ms4SMPUCB8uXe8bo6sQRddSDexyili5uk+wM527
s3Yl5daDzXqW+55VqFBXpev/060SNLtbU+hDHfhP359uEjkIo/t1Qe43w/cR6HTq
SndPkDRLqPwzopgBgAXeYKEX2A6aE77LHBVTJ4tc8sFKlWv70O6DRawtADxbw/Rp
1WW+d+qInU9L5nyI33WNh3rBlo4fHg1skKhGHtug7mXNMK9smdpylsfgiaNR6Otx
EHbfry+mZH7SplZoVlJquuI/ENiCXP1LKITqBgSjhE+u+dyh4aE0cE+Nmz19GnA4
qvz8hIKmLlCmLBmdoqnxd8q2pvk4eQc44mZbVkl5IyS/og796g0fVkRxSOXeT0Wt
tMn1etShSaB6MpHbByDvszqrkjSIOS+0icr3wFe2Njl75USnimY3zvIl+CavlBcc
b+6u+HFonU343WQIZQRNz1q8IeFQiow9TZ0SDY2wyazY+sV/EVtRTf4LTJMOdRmP
4QRXlL628dI2Xe1LgdWqlBdsGCTxDtailumxypVgHNV8bQmrmF4aejlM3EtNbhfj
Jw2VXObl64c0bUABjwX6J4sqkR2/RruuI3Jh13sJcaCuDJV3QoJDhJlhhD1kbFQC
0llpEmKwVK9yYZg8J3foq1qfYuKbzr1LEeHG8Lq8PYzyPaElOvFGVlEU3kShv2oX
ANGRQ3heyLH8a7Roz7cQv/j+j+PzEF++qu5YB5vbh9wUnvbafvPOFsn7hjRQzd+U
0mwruav/8eDO9oO/m66qFpO67AQPrQSYqXOiAAr4hsQd0YWg3OqSR5I3G4CPIAF/
cIvaAKQ1GXv7JNgn8TJIHwHIV+f79FN4VjZR5IsZtfev8nGF5gYmP5ZRYBTEhaMd
24C8JGqQMV0G/zzFuyV3C3FHZBoSlV3AY56yjvG7F7JNFiFMBKF/xH8WI6nFooPl
5E4876psIaTnOSgIOxsQHxQUJf1Im/QMyF8UFX9eCpTUF2y6IQ4ArpEHfSGfgDSO
zj9Jf+MBBGSJz+jEYNZL7UIs3YHbpLkxjLQtqlBSJCk/p5ST6tUCiiN6hLt5LXe3
bJvh/1L520d4FBExx0+gC8LKKh1MBZW59HyxcMcMS91Zt5DuDHWEILhozG9uTr19
KDAr79LCk8OJn3V+EewfR/8xgR/93gR1u8fK8Dup4bMFVMXN+HKWxHXMFCgD2dC8
YGBfkj1Fz3E/0aYUNPtF+68CeCNChjOxyyMZT3bEZQ31PsqR7c85IyOtOlBGyjfR
kVDBwXpNcu1ewAlNK7WErHQZ0Xh1EmfKSc8/+lhriWQyhQUeFsxzRw31M5sA/0RH
q5aQBW6RE9xrpbzKVk5dErIK5q3jLihVrPtfIiwf2l/7yCjotAVsJBBwfYAp8YjO
tgjeSW8PbLsJIYxpeYSv/mQAf020EX0dtHI/Sj6oLh/lHqPoziFa8v26TwENQAp5
SmW1DbCZkTEQyorBCWCMhuBD0oebAtrEkW4ZbEZs9Un5OfDSRPDxyDhd3qmkqCeT
BHFEGoPc0o3JUSUZp7MY3ABTE0xEDT33xOe8vC7NtbPiXeb9TtbuHCaASoVOeb1P
Q5CSYgZjq6E6EnrZGufGtipr+T2M9PcJcLjjjKr3SYb63+V8QJH2hyp3NOaWzXww
VZmPnX67GPyTEldGe3cwyAK3duYNYdaIJVWbjkKegvXtUe0CmHFTiPv0bawWevXT
mqzPCzL3b7iZYlCuMjS7s0YkGZC4uH55A+PnU1Jrd/fYZWMvv4TQ3DruEXNOvy5b
hHe+7sWG0PqjmJ/aF8ND5auiNgNJLverjkrdRwE3Z8qQvZfWQAi5A38v0Et7X2Ho
nfB6rjPGJZjanFQXnRzJbmpkB3YUTRxwsbrtZ757JmVHFka9kh9jOsSzf057Itt8
LgbSr0oPO6swgn9MvnZgAvR/DLdsGBHI86lwoS3F1ZJ2N/8Cde1Gtn1WTt5mxWE8
E0kAxUFZkGGzPbFswXu5wWPFs7Uw7CnqqYt1ihTSjXbh73suO4kZC1cFmreLc1Mb
pt9Tyv/SpXNR5FaFNstZeCREpEVQCndnnmlA4lzO9ky9TK69rPU6Ji6Yu0kH/B+L
X1KwOuks7bv6sNRdY444Z+CAB0rw9qNF0SdKK5+t9jAFFHrMit/E5aI4Ktu1n+AZ
Lnw88opfd7DL609YGhieFi02SH2eVy+RkNvtdUrSCc6f7j/hHYQXSWPDeB41rC9s
0T1yL0ewbMnIxx3wmWKRNjd+sfOFlC9mGZimsBSvh4vwRBXL56S0vZ2c6Zuwpgir
HrGxFDwNbXuau2iaf7PQCXOUWP79YnvNH6+lio8rRZkrcl0iYWLo3YRw2WHb3ts9
mQddHFTHbY4Ppr3sq6lfBcFoZoP37EqtvxzbEFaPXxzONp5A+xhT0xD7WIhRkhc3
bfET5rqrbNKsO+5mC+gz3SluZvIcRVuLYbruL/ycO43mQjbOWdEoKMRoIxyAe2z+
+88wX126Vz/I+iUmnjJAvAuicniNVAIvacezp0MHFzsW5P9VOd26V7eJSUpNYxPc
ZLO11BRWwL+RhazF82R4wk2ySdw0ezYDmLIU9zv2gm1IjTFsxj+Q9WHYenRu4Axg
D4UEEuMttpJomJ0ARwwoJrKe4ALH7w3sL98eaGBasktbqHrX0B8x8EkuPaYlVzj/
Rjqy6nEpHipYftMttHivQ9gUUtWhmvWMXgeY7IqrRsLBEhuxWGmOXHRwyttfjiVj
wocfpOrghNkU9e7BXhmpFVRW7zVTdXj5ZOcI5hCKBBa74aT+l5Jm5VscUxMYXLiZ
kzazjkxopPsSIxT8tAItrNb+m7UI9ZMiYMft1QGLNOtxEag+obDWYr5fhebt9mT6
F4kTVyKPDfjEGianP8F0lOp6VeeEj7VKMvx3wXh9hiL34Z5eMirK+E/GScRCd5lP
T24UA6g3B1gY5MKWGl/h0zNpF13Cj5I+7iRXfH9g/+yy2FyKK5mvBpN4WZ88dEM+
Z3yTdpehfINmb6uMTBiiGDNgewU038v/A2/GJ+64gW9DcHh9pGIZ0s9yu5BZoy7O
tTS5HUzHd7jo5Ecm4dUG4PWY7If+b5rrJgkEGnzqy7eL31aYmmswKXGhHmLvrcpE
vvZo8erRuXG2xXwQeiN6wG9IgYopC8T7Q9UNrLYo+S4URa0vG/FUU1/1EUogojkJ
/1hynWSxtgeW1aY/1AKO8Xabq7FO0yZPambgXGZAl1r1NzAlyyFVzVWVHkdRtrIl
eEgPd0uRnlQizwDP+2BJmCTcXVLIsPJ3FHeuvWDUrPr9GpAOYcpPDlJPPPLXsUyj
80y0pg2XC2R8nuUkHx3yAP9fSi9OEujpR2XrTpIdM8w62HSV5JGcVwUudJs1UnWK
jaHYD6NBfOKqYLkhPp82mSEcLCpmb8dkXRVyc9SUBNDfFv2m6XwA/8de+YuRKEmv
VzkMhJGHBZF4RxrO4vOmW43q/wsbb71grxPUIm+pwgC5+kAf7tib2HT42M5i8giw
KV+gVsp5vU4h3i+TLHxd0bJVjlz4HZ7zuEL3k4tjuvtE7g5w828WO1DEWDX4QSCD
2wP/rDMmRz9V4lYTfRVqXsVxHZezjHR8Up8WZulLuRYKQfM7w1LhyxLfnhCi1PZr
aTqxGTafJgCpEj/sZgL+1wO+Xh8oVVSvOHkSNN/jGo5ic3ZUnGPmZDMq5fX5PJy6
CvDlDKcPncfA+HLi/CPuaEJihKSI3xBzqoYyFjWr2ZHumzwjXflS3aXnSRC5QY/1
yuyUtL4axIZvmd+aOjK78dHaH73Uyv+RqzdU32hIejUNPzlZc1f4e7c1Z95c7LCu
AKzkqb2j2QwUlg4R/TmYVgFvtm8WoOP1tjAInmbL0X32fPuACP9vnaJtSHIrJxVX
efE8I6c/9n7VFXF0w14+fk2Xv0U0jy/iQWnBSoRYlebolhLB+kJ/d7gLOZUFszkL
tofaNgj4hwXYuahPA+OnrqRw0/s3pnlrb9KBzOefMb3vSODTDqJIyEwIl/h2Yz11
1Fpb/ku0WFOvqSGrmmjnckVPqg0CYcjKbjH8dvFtN5fEJn2OiyJgLAI5Zwi7zIfK
nwqRDYUDK7StEeDTwP2vnLdoptQU6EjqzTv+tjPB6hhY74ckVcGnrEFjdwkrbXrA
4zD3Ae+1o/9IjBfyXEvOTZx9d307qMbGxYW9wEmMtmxkHGtIWY3QzzQeKVOtHV96
kgwoSWH/RJdkaKKPCW8C1cZo784UGGzA1pXw8WfLia0ugpwO4ZchfwwgbKRNZoMH
514DJVZom3tspqMoI1irKRMUqQ25YyjHHafieW5ayW61WqhGFNmt4nhoeNgjDitl
IMDBZmGLXPy5D9PF7CRldobBoTGt52md8hXc18g9gdhIA4X5JQkUanupkEcKArLR
dR4tF0+EIkdCkHhCfpZnIcn15yY1hOCdBxNm/O2ZlddlFSBUeLJgxesyzYxUSj3D
TQyQHRqTcgbnl/0sRLS4XH01owskjXq3KrNr7j94GQQaTzK4qZvPI7OPCZOarUnk
nsKc2fTJLHgWCmv4FJVt/liqm6i8OArrDnFOFLMMTQdv5xv4+1VB4QjyblykDg39
Z4UfaMtHFzBfEbQo3bRwn16KxiF4ZOxUWwZXxeIIUlvjLqEzoYJF+uecW2I5yCgN
0b7N0jZQV/HcbnIgY2Ra69zKUsmz5Hjf7kkmhOTmyitq5WPX4mLc0l0qH4GEZQeb
EbWPJOaYbK0olmOvrFDLOiz07CiPhaVqaSqpkk6M+FeHgu1Rv2xpKy3Rm4Ts6JOc
QDtumOQkt4iYHvNYf14cuaYaePq4QbGbsRhwfBuMuqlxMpiZILysIll1wBqqNkXM
r90NUUlq5FrIfZxEzhYhaahwFZEhbEnYjySL8OFqMKN/9RBhuRAWCYUZ5GXXRcVF
3a70tIOfomhbflTu0XBwHQMDsfNljEIKJxJvAuH+m7hS89pHK8IGW3PtfgdZUfd7
EczwF+Ej+zw1cKHmCw90Ud7iaiYjm614TlpwNTkuBkx+mIafnevsWvTEYtypgRC4
TrgaOez8Nj4ssx3TAPWjq4sbfrAnmdLyhZv/vwuEUT8c7CUh0cFbW9Gmn68uH8Ym
1k08yQeo789jtK8MD8kuSFsCQ36dlxOPQyxjYoneAeYXE0m269nVYv9d+YHUvNcC
lB43l2nx8RrqR7PekvZjjJ9zu1Zy5o7HFVgZdGcZA7wS0h9CYIS4p5OpaVAbHewo
7ieXMRO/AR4qfaz247zOU7R9zDei9Nq+12HDh590qaLqRhkZiLmM0L0R8A9sMiBf
26CbtbRxk2eLdA6hCTWw2fSkLJRxtQaAk3TMpP5giubsrWN4LWDb9Xds45dHscGa
adK4uDiKJjt57+HVapV2/CeojrpMicFhwqMqp/xM8GPkFsisFg14tFpEg+/2FwDy
S3M8Es3NBPC1kg2/A7gb7Wo6TXObpL/RUaO/GvGN8iORGkRBnXHJ1QK6b+ZlmWf6
gVynPm2PLPkO3VUAVQtZV+9/bd5czqR+ak59x8LiE9HRE/E9YtgpVwW9JRU1veIP
44hEWiK3fryrxsksFNK8WMPrEmc8stdjy9eGAMlkzCTd8HsBDIT5KiuQhOTJkMif
kxYZoBKg2BRan3C1+1RbMFoonP4zUoytRfH7gjcRWNHm05gdkzOS+FRAVz6wGQd1
vcftpj2pZc0avFdtK8PelIAX3wDfNLZHcmW88J1DvVXfLYJP9GdgNtddnpTgik8e
uqqPgJEPKYiVo6xvrRyCiepRU8fFnzMFBzUTSr7ct8C4XWKV26+xO2OSEMe+IT2q
LFI8I/x2TUshieC93rOhBu+miwh0zGZOeUUKM0bHe1KlpCkXNAQIop7H1LCc1wHG
Uj+9o7RTLshy6uiEsVE3iMd+x9mcQHZO7+ESc6vdBvc5tYLdOTlQ8scxR8I2+4TT
LxLkQSh649p8xIPXtTOJCB0jvixcJyuMV3ACOGXFVgx8NpjvymtfzcoqrY3mYwC9
UyhxFZX6DLNWGVyE11TEI0EW094YnZxJ2Dj61teITcSzotsiTRvtyadTVif4ErER
mv+PZcgu/l2Z3W+G9dRRIhE41VAn1sUwQqCcZlzGDPs7WjX9Ic4Wn0iTLMzB8Z7s
Pe89Ky84EJuGZTJ4GzhBoBbJ+8uqqpUfM3QRdbhhdLfk8MAtFmGnbPBdNH7Aw4Tm
BeyLy6zOd7pyUyQ2bTPQeXNlw1XDWaDVIfxYCZ/d+haGXPM00293RzJ6KcFOfXDW
kcYHxHua84f0MLCQdkilxCNh4oCGkfUhUDjJd2nVAppW8usDh0HOhM2CZVzwdFPU
CRX9bD2gMDVjS1tyGcaoDrHkUWlDG+i/SwHiHoTZykP4gSHILaDfVjZwmuJBQOna
KD7azddg6t3GZj0hC+8xwZWt+W2iJLsFLZCoxheIImmq9eyCaAaYDjZ30RLeaatT
OQRFjqPtI6gWplz6VREYtpn6+78t8Ld9Y1D/YQscoLMSt4YbSt0/DLlEsnFKi2xR
TiZwv657xcH7DrQgDBxfzEcrwmWgyZqzsBIHdPZ8u2Vkgl0aG+mkLGkL5iima6ul
xsmBzIq6i/DiM9HD6cwIT36DPU19aCwLnBuxkeOxf3sD+1Z3E1qwOMGTtmTMgv7X
ohpafYH6cUdNe3E+aIaHqnt6Y/YYTls0uToHcOnJxX4PCL7f5ypsZ9HnGlUjyxwZ
3/D1gUwifF3qtv5QuIo+Uixzy/Ma1b+/jjHMIjEiBpzduSAMzpMpXpoGpVgQiFth
qqv/v/l8rBbdVqkhecU731Xn0zFkTmXV0Tq1EExZsbxwTCqG4X5wIqQTiWvPnKb/
bph0bMfUoDAda28MLd+ySIy+TzkC8/HuTzAGCZYs5hCEdfCkOtiHa9Aw56I2uCI3
qB/osL+LL9VaYCF9bOVrS1l2vLD1+Vyo6IpuhkLwB6Pfp5XkFynTpJrDddd5JWfX
0Me2jWxxEJpUyUHqr3tba/5gMC7ldb6fv3i+0mccnq/pYV/L/nUnUZeD9l2UccO6
yDpvao/PaV2B4vltaQX31gorESnALOEBgcQEHl0LjKNtzQvsAL+RwL2ZeAf8fBwx
r8h3D9OApoV9mh/DVcpOyHQja8oPQklwnbwJOPv6c3x7nFS7a7k0pPE7IsEeDT5e
cqVIl6fZr3EMU4W/ilBTQSvDNAkcVeCFpkrJOATJHyvCok7UKnqaYBei72be1UiF
2sCsZlyic9V2Y3eSS5LbRwUpaxv/+YXqwLh283tuxM+wwN8ffjg5fOxIsUv1SajH
dGKMTJ4AlK6zfdneKFMGCe/ArLBj8GQ1aZsSj/jUtyx6uloFgdG9aA4Ap3fWf89Z
8JX+qdfxjC5eMMXExRt2LONziMkBgrNjnLpBbQttOtRJ0F8J62FF8+sd9X2pJAXm
MbUUyDmMk6yZXx0KNYZkGxvXMpJB8xlQ2bGL3H/fC1mnEOJGUSLzH4MEC9I6UvuO
dp9WvbSFnexZQrEIjji8UdoY6GheyIRcH5LtG/8fW+rehuvtElMOyruRZQV4J1cS
a2SMtJij7htas3y3VJEmFr+pH40stF+IimcnYtFxDvoKQbwYbqe5xVILOr7PsK8G
k6iBfxzaChda3QzzadwYtVRXxBJqocK4wQiuKW5JcXDWEmX7JDJjpJ3m0HjOiuPg
Mrdzl6mVRAtLexCsk/4YyfpG+HvhvnFzYjURkg30lLQSvg2lSLPyt2w1K0w6oG/v
yhVCfESKCPwKC2qz1aWud/Lv7xl2dKsQ7w1QDFmAcL2/7Yjoxn6OjYDa02aegBT4
uQyBKrDmtRYZxlVzlX2REbc5KBvqNuBF60y8smNlYAqGVbRd5LH7x5b7fGl7zTC2
eHqvBtrzklrD9WRKGySBaV52OuKdyLCj7L5xOVQKFjvYoES4VihIxiAIOvKyUThk
6Xe0alW/gzD8qNotHR9xgWxgBX4cUdZVljMEKr6fhUyLUfKwRbDBBCS5hT9Tsvc0
y78XvGuzINZlPctKZjy0yT8mdLbZLXN86P1M79BvTTZTzkYF6uL7ZU/nKinJu6MG
9I33p2W8GCyrY6ZZIG+TiuOOvqGqp7qFMJVbsiXUFuxBCni2zpxLw8oYPvnd9SI9
3qxfqAEvU1cB26qEkCJoYijDoRKbW8r7qWnDP2GJT/wE7D7SIRjgswBedIXW+qjC
4GFohuS8HJpdy2nik/yg/yM/eRhTaTilqobsm6Jge9ZY6Ri1P5tTKTBs0C/O2SL8
fG7Tb8iahQ7oUjoSL4NCtJN+ARMzuBUWtdR5V1QAlp2kAaqso5YmlOexRIbvIocY
XI7EUtTzMP6qCeBf8kC1yHq9a8TJknfPYkQ54teSIxkrRP6teCYoFt/PtwjXt6DZ
w8W63MRNfCgcc+AxbB8jRC84flUqt+1tvp7YPImfW7nLMaQU4jHaCIF4Cx/w7gm5
rDUZILeEc5T3K/9fKU2Aqp78np/NFXdqHTM151wzHKHdUFxDiHwkDxPInZliRl8K
BeDV16BsaJ4tS/0DZTkY9MfrjXZE3bgquh2O2z4pEsCBYhHZ1c4F5cdygU9CkgHE
s7x7oFj2eXYWtU+0zt/GaDCrwfaz2xeNPF40tcDuFy9h0UEh3ceOyh3BuXhL/yaP
gYlugEl4YYkfokNMwhPUPSawjY5bI19OXl8HxuKG2uBaf4/UNv89uI2JZFGoBAPo
S796ZUOv1uRX2EwVO6cyfbc9EzbPBQ0Pdo+o2Il/IckfQqX5D61RCSCXLIfLmylp
axFXVoC5nnh7l0RS6f0EbLBrUMOPpTgVIh/0Y/8e3obX56DhkSJPivkK9VJq7JJJ
M4sKOiHMnMY0XXxgmFoGZHzWJRrIi1wuprY9tSA+FrUto/QmbZfdXjMDid/yl9Uz
sYC84iiBEeFehBakCEEn31DFpWt06vQP14TxQPTPft+vRpjazb2KWz2BlyLKJzrX
kn7XOrmvaJC7x9ZCmKx4G1C6bNyqatUCHPF1zWLBDFywUILPMXqm2dh+pbhKkhMy
Mp4MaO7okWQAk8P2qIQr0kc3S5eJBcvoRMQ933nEcr1gS01YdIZokOJQLjJhORFt
nFSc7SY0xmv4CkBo9/tPpngLBlD2zptIyM1ZrW1gDW9PHMIXLRn1RwqW5ep4RD3p
wqwZRXLWTVxICDQUxig49sJ1Sk7AuNKzv1D5Sa+sOxjsjnPggtXEjFEApPcClHuS
0yn9Jp4LGnpmlBwFxQiiWQ6/gpkzPqYujDsk/WJT2vKlMDFHQVYwgPxSS3Qi2qPy
XRfVVY5W/qYAWNLzRB3U6qKsc+kRqWCFPFoXmG+NUCDPTAXusLetzMiD7NmJfqqo
CqRu49trKAdLEcrAT0E+zJT6mmVibNxw/5XJ/6no16E73iwQg+a5xh3Au4zi7FfL
qRg5Omo6WSpEHGf6WeT5X27jCCwSMPgKsjeXWmcKl5YxSlM+8szrc+mw0w8xlFdT
9O6ub4N0a1RdI6z2E2UNnfXoAP6cHOkcD+2gjXkJ+CoT2hQvRT3F+DnyaM09Jtt4
SCU+Ne+JpqwqT+BQpwS6m6TRQ2q8O99tsaDVEvXXgxFMqBWNnpa8iPWhUHjg0msD
mtyLiSWtyjEkT7hjsPpZvovVfHET79kJA1i/kSBsFQHg93i9sVq8I+Y0Nj8vtXMo
o6r072tnGliiEZzOG9SePaotClodPgW3ecndgaHMb86jmewwkeQp9M94skGuyC6V
Denfscc0WakE+GXEViBma0n6KV1/LeSgbGsOQMgF6DhvrkU03fRyr1wkBgAN5XW8
WBBKBOdHXMPNkXEPaLhyJPaDGkCJ7oyqkB2UDtaTvKszidFyoLoyEW4RmV8Oytiz
f60cjQikKv3GCuT8U3o7HniZbrmk3OYD3a7VS3nKKUcRvHH3gmTganvPqLfiUha7
E9ybOmb1Hii159/SWGtknek4JwypNtB2luhLJmoj7+yVTQ99y8bVkEWR3EmAL0mQ
nJbLIaxuOXHqnG3aehfBZ66x1ui5c1MfD5kh4g9bAbcflhateGZAT/xMsDn3WGZW
jeLdS7EC+sM1jdV3rHEYUOhy91Vb/p+cZrz4zbfIOUYRJufhZYpLesuYylxbAutE
nu/J4E9qK7BKSsVbH98M8v9K22ErdJbOlE9FFoTlAXDAS8twDiUP2CIovIPQJzY2
TrpkC+rSdSswQ2J6UfSBG++mtjLRWFyCVUyfkvhQxrggvTjNjbfJyeegG770VzP9
Bky/hqscghX3so5g36HVDUi2qoZNhoXS4dVeYCppl1w0UFroN5xgrf1mVt6oUgH7
v4TTACc2T0rxP+jW6Vt/CJ9ZMPL5VBoG0o3x+zi1BdZRx5wUBRDrwdEay4CAHuPH
RSkoCAQuLtW2Qe0qXrYVEqmR1XMHW8no/15sdyKgVM3ma2k823YzxqkfBXPQ+DgB
oEs8O2lSicy8xNlLzXeZTF8vEAGaHN7LbErdk6uw39EoFixsYfNC6i7UjVTz/xks
QZv7+5uewQwZ8R3OuSI6DwJ0nUc5ufzkuooY709neMcuYAcHVtBiKOJKpnR3qDbh
ONQNLL9NYgsw8xjXSpWufKuOIv1OB8heOSEO3BY00hC3NF/xrNibKiLamWsFWoIs
FaNiW4as9O5pqLhBrYFjWIdsY1Dl3WP8HkweFw+S+GOKYtZGKB5Il91bOMT3M3su
3tXzTKKYDicyTBcVV2Zin1H/EwWylm8PcB0LAcamYWGtgJoWrUXL9AYWKhfqcJZN
Zy91O2hdWXw/MEMtm8Bw+8DEkcuPYD2IWBTbjH+TC2b2Ovh9tZpG8Bw+kUrxmfow
twswa3H+cbi/SMMx/SBQn33K5uFCGwpIyfDXAYkVQ7w57jjyw7ZWbiVi2lnxYfzJ
NuJOAFvXYL3BNs+I+/aVsCTlJDuGrI+kn0U8ZwAIpFCb9aHK1jl8/1Rgl3Z6Gi/H
pDu2yz4U/LkSkUZhX61waLw6zQn33/V/IW2tTARUyIWq1nwvNqEY2h51YHpjkZ15
UUmSnhkXzbsQQqI+554B7FUIMID/jge0ahNGxC1u/zl7Tudt7IDe/5oC2XDhuITq
s0HHo+2dIcAO9qgft3IbHGEpwctbt8++I7yPBF9TRJNHNvlSaZLayi475ufhBif6
jl5Qm5FNVeBhzVrFqEOD9hTfFZ64Tmo6FESvu4Vq9SB5We2sry1iGyoOo8rPe+Xt
ScvNhcl+nLt7aKEFhQRWt7tdVPDvHma8pXjwY9oeYqGF9UL7SMxOf2KVGjtg8rzj
PUH1D4bFGdZ7h46rRxzugHb8MdcvDXbWQ9x2AzKq1rkyORkZH+H17QslMW+rIvjx
bquIBkoepfvOoEpjamkhdIGUqlaiRp3x2hIKgZC+1hLKiLTu82Qp3eNweC59z3KG
muHRKlswGU62nlldvJsHKgo1Ik4NoSLRXbJny+nllKNb80KjgSQ6oeE7zsFFd9b0
oZPeaXHCcEgYgy8h6EtpgAXQ3bsO+4vBZxYZGQGkNLAXOO3mzcomH07Lw0dxctCH
FnwXSSFzfQ7VO2ve66QEuIFhc4MA3w77jvziiJG4XhnyoH9VOzIOswCVuGtknnQp
EWhS/S9ktMFijyh9E6JnfbmWxDelxKvp9jM/AsB8vWl9oAoVd7M4imi2o1F4JpYa
D0tRYsOppDxnDfrbInUzu14g77K06nrDdX1vkjrVGb7M3D2AtWm8dJo1jVw+gDZ2
u+avq91nC79nB3dAL+jjmYfs4WSrYHyex5QYbECdP8Htvgv7X84JIm8OHj6vqAXs
dScEn61u3V+14d4n2GeqIto/0/sutdNSRqxK0RMbBvPOLiVeqctg09f6FECQ9w8x
jZGkqgat64gXru3wf1phwkgDNTr3CEsxTtEuBfuaR6JzVyXc4ExhdN5qhBD20taE
Wphc8vT+EO1SWunujp0pCgeb47qWXyC8VbQ6cRAVO/GbTRhPqYtU/uARp20AxRwh
C7THxy/LUMXvRh23h8ywwNbNQ6e4WldX/e3BKsB198Lw5fMI0VeT9eIJ6UMy1oiV
PAnRQGyKIXe0WuXncz2ZzhbivfQLMyb0jCrcKi53x2yHxCtF3YlQgho2r2Yj38f9
y0ZRi4NRWs3jEwI18FnBZCLaMPpDK+YyQUasNcMPAEq5qlIFmyAe2P+IS9oDnsWU
knxqAoowx79N51tP1oI0xUmrzB8v5952xQ+XtmuUl0gwr5IYrEcuswbtJE8bg80t
K3FIlxjDSCJHsJeKJ2PS+eja7qeE8OK9tParepHNVevWywrQjY2mB6/vZogsPjxR
fMYbdcwiMmRy4Zup2NEya1DxcDoQtlPbDnXoDEEkuOxZUZ7ujsuZq0YTsxpV9I2n
EI8EmpIZnMVtB8h0fNgGnxZ/B5NCLrHCM5o37qqceGJn1ljMX5VDonnRxlb2r/y9
4cuzSGwzjY8FBw7mFcXxtmuYSx8+uhQODku6FbWDNkn3zasvEWt41qVWO65MnOpQ
0W9PCEefbHwk1trATv8R27NOfMtaBI/QR6WQhzmoGWmbloizmHPIGyi4yfOc7655
vTxHLfNhvf45DYUG8wwbt7AcvSrX3+9zvHTv5tOLeDtHoMU7ZrFO125lf0yu5KYA
EgKSaz5xa77er//I+Z52Nyz0ZQYKisOJ5YmMBFwo713sI1hFs7FZnbgykxLZYcTL
BLPRNAa3oBWFET0Jziq0pgaNffIZ/5OMtOyaSlx4DCsHNk+Xc3NmEBXYv2p1dxM0
HSEMc9d8m9hY0acDxMFMywwYZGHrrIo0j0sPhVo4Ea0R69SJ3vC3D4lHs6uEUs2v
vh6zyJ3NT5dim+5TQoUohijf/kKD25RddnoSFW3IjsbD2R2SHMFY7AoXAbmT1On8
XbYuZwA3GH35WlJ2JEFocWGbe3BMc0JyTtIGUV9MgtBFlpmwDY71zMd9X6QBlgyk
gtW+PKInD1fYoLmGSscWJNLq9K43HiGeZOqtdL5+Qr6LMLgXtFEtpQKny9fEKyPd
jIFn4NYNyJ0PMIqVK5crEwNshjY1CzlrmJE+yyGxByJkJOIotBm03pJzMHbZMshj
xS0SzMj4qovyhZSY6kSQGKt+L/ZU02xN3FL15J0jbAPTVReoH84oop774/Ba/e+Y
jjBa6lv6kDaY9bJ4XwJHOY9VmSmQOeL0/vw3lrAZ5Z3DPQMifrWc6k+JG6XvEbnw
Sc58Fl/mUvh8mZmYkIc2KnndtddCjW4+h4IJ5b/GduRZTDBKtALkgfjq2LGZBpMt
Gjlz/gjr5YtGEp6L/OCUhxDTTGFe06AzNQlmrVBA0RUSgvJOfnwUqnHZqGhsLQ7Z
pF4Z5Wzdk5bZUDy5ttKwcD0+tLKxv8QROeYQ/HzLQLTDnKbksgFVd4jZ19+wqpvR
GQwvIUitDoYl2Y4uwKCghAX37wmSTHLQ6H2fvT+xVN/2ZnC9sut7Ctj8DEQR6Ka+
TJPSHrrATzaEogU9qWSoZVOtA0JeBNovxxi5foNnzG6O+LbJaL8AN8WRN7Sv+mvZ
ckrHuIfWs9fv6JG5om+d6zo/ZcbFiiEmwAOG5vWpNvlGrY7gcBqshjLtupPKpAOW
iSOFvEZp0VS9FOtLurlKFuZhNnsRkwU5braxhxs0iV1DQQsJJ7qF6SOHtx5MXFlO
3zWh/EuGx0QmyxWSse4mQbx4YZ8No1roNx34OdedfwYsU4hDzx6msPkii2bU39AC
Bk/Bp3chIcKYfJqCpFDTtDPJ1OJ2gvmLiYNrEQ1T3hRLn2A9VtyzskMTBJ1lPnvd
XDVSiPJ9ea3mt8xjVA7UQA36xUMMZEMJjQPfW7404EdhR313qZ1hXJ5Ui8Q6sddl
mfj+anZtKiivpZmqxH/HaYEbvxImA6hsldZKB8ARYkeok2IhYsYqbEWEKEb4kb6D
6enEzOP+cCiYAt2nmUypfeeyQmKeOZ3DpVopG4k4FruAivsbq5MwTbIhOfb7L1TC
FCgZ3IvZcXtingPPo+kKA892s64f05ee5hCEh2ItP4KV1ZY2volaAJowoMAJS56O
MqjqSAtm/NCSq2anrGkN1E6P8nei6/C7I2QtmFPj6DqrEv9AAkTuK/IARdbIbCmD
jIiFW4FdKWdGM/F/4nCdr78FlqyPi/OiXPov1e2nALh8WVnb8J3BpJpXrabf0YL8
1JwYR2BldhDJR32djP+oQ4D8imhimODOpgV3Q6Wd2x9jCqlRrd97hj3iNCGHR2TM
NZ0YIAb1R8eBn9N9Z2Fuj0toWNtRatVuEOkD1sax5XdEgbB8bREeNVNMWSxUVkwb
WOpYG0MyUpAzAx2Fk8CarNOQucunUgNlsu96J9PuTgCmG3pl4OXQAUqoDGqvNIEt
eUvj0A3wq9kk9aTyJ4y38cnWO3xKQf6D1C/0g8zZ0FZHe+XdlesuP3OBDmqxiW28
NfeGrT5tpqzFT3eQu2SZcfxxzZF/KlMVrDgMXnAlTHomSNEXq5eoUnh9lWKY29LN
hKN06AbOOsaKNxgRq10icbrnChrpN8eH25m0O16H/Uccwd/8J19YCJxXkq9AGXYz
6Te4+CsmfFTdQYO6jCrCx0Kbnz1XlUS9sqC8v6lvB7QaJSpoDVlClS9yIHqip+2Q
44PhPYNr8yI5URaKff+36iPQ7Uo56k3SadzW0QGhmIvsZZvBV6jEivH6wCnvrj95
EctC0oJyGC9Sa5CzOFOaW8HvZAstKJOYWY5sgxZDNr/ZimN5AWDmp12r/pVCdQPA
Vaf83osOPoSJ7kx3sIzoMQOWTcj1bMjWXbYjr9dyHgOinW27avBsOghh3xC/Y2kv
AgMnF/ejqdqHvi3tnfcEGlhukbZlHM8tEAZdlzakJxuXe14RNDrupR0wJqamWJc3
WZbTMpWsY81ioVYoKs1A+0pR5ERvR5TH+Cmr6v0e37iRzzpROsmRkyLa/M7V2q48
LAMU+WM+Jq4pc6xWxTwuytTvHlBsoUF6H4Gp79kcadvlLorP7y2gJ4FzWNF9Oo2b
jkCsse4QoF49avQPOv9JfkqFcclOy9ly76hBWaTmael5TFCg24f9j/RHfD0S7Shj
rQ3fcdwCV/gLC8XI3PCW1YocR9VmVLyQ9PZtxBJ6A7OH8kqZfXy9yIyu/4AMtGMl
1eiFrEaxajCrm+RSxKEJo9rJpvmCf0YDnIKIdVD/72kjRBtUZUh1/F5j7uYjPr5T
zlsOL2TYuFxgwzqz0dU89nl4uDHPemoWzg4UqgYAbM7dhB8T73RNYT77g/RR4q9y
VmVMBklEp7Io1V9ldSttUZBwvYoeXQpZyERH5HVExwUt+wyrVIv1n1ZA7knSwLM0
0lsehAiEx8H9b3MAS4+9NDUkY0PH94ODJtzv58HKvbp7/xAu5p1+4sXVXwKrahbQ
mu7FIC7rDw5b6TJnNYopT5DFSScSx5h4K6uDAWVLVSBYlYL1jLo82TJXLHfO0aJS
4KFojDXANhyN+7W3h+UJpfGqVd2wzrZ+Uqcc5hmcUIQ9P6+pSyot+tbrP5xUUv1q
12hZnBQvIfdjCvdY1XxZliOoGDJvlWiXXjYASdVWikdq2mEIHGYlHaLDApORMFo8
EbxdiEjTUp0UYa5G6E+DAtLoOhvGtVFB5TA7ERuaiZektqjlbZmdkX8rkkQs1/e1
XVmdNjFGXmgYabktYZSNbMtuCacgL7E95jdeXjINo61oRzV7T2Oda2isQTVjg9Ew
YgkgunzVvMamarl2ayHwCKkhiN9fm5myH3tpwlPgrKedIlh6Jhfk7EzN6nMyOlfi
HnqXyNpVpD+yCiKmm+VBtebPV8cfGcPu0xDXZ+WHAQ+pHbJfVHEX4ZY+xY8IUnEX
+cusc1BhGXQSwf8JYJe+bL9XABUmfJVz64OpJky74+Pn8GzCNCWOAkaCEjh3CFWG
QoY2+HtcJYcWvhyU+hkvQT/HJTUr4xeFvAvxbY3cHb/i3jf/Oadz1OhWUP+eHPcK
NEjG+WNQln5TBW+lrWZKF0SJ/OxznhEBQemmNASZ5apkInTugi+24hI4cAwSVa6F
jwvgyw33Ul4yIXNGmnJldEhtD16UcKdbXsvTXrqXjtaomaDgde/S3Qv+ocAXrP4/
1MXuFA1tsiVhhjuNrCFHGtFKajVsVBtlN0NGuyhwd2THyHK7lHGE2zU4+9E6gaZG
+XqXPakaT9X6ctwEL9YXQt00+aFdOzOiWSiWfEU9pjMRGXtAmrty6zgWPwnVflQP
342NOGVeLqn7kMoz3E+gSpTHjGsnAUmqzDwt9BoYNTD0uGtLp0ezktVPpim3Ywoj
zaFXeufRf3vdcNcZsUTbIBHdEWhxFJe8GliQqxYEVdSF9fWRWDgx2RJK3cm7GSK3
pPeyKQsaQH/pEsKyYb5HdUuZe5q4fKkOFC8QEGxzkrqH3S+W6GWukA3dEXWlqswz
XF0yFDrLegTffy6v3jVC56yXTgaqwj8sZyXS2IodMy7ABZETeT5D6h7OofDiRSSs
d2ZU2T8bEriETsnZ9ATgG8UDCVbAzDs6nSi9X198D3ag60gks4I87nrzjYdLoehC
r1HI6jCgHFne1wgiJrwYauwYkAfJ/puoE9mK1MdLF+UbTOxy9XlT16G9ybZRMyG7
DvVSzoTEL7nxXfhZgwthXZlmxVF8o8/f/ndTfXiScPFWjlXEk2mGKI70mOgcedzI
m7QqC2J6XoTRa0Of+Hl7efOf08qUFtCGi4Han+F3L0Mw8pbSJ/nSJYC36JSJ9nEj
eMS18O7bWjMQnWdJipmF7rX6D3P9AwbJ8uXjY8oSSTV1P9UkON+hqPQf37BNwvhM
wcra1utfM7xJNTS46bn5GJkmaRpZkCCi+LgVlYCj9XgeVVzejIzsBg1rKfOAs3b1
9UMkhRcAAe+nUfZ57mY437GTWEtjR10xBIRqbzD4S4if2XR5fYfJjNv2kdpUN9wu
uILINJaWCNPgmsC94v/LsOOgen8AO9oPvjCZDPSulbCHYP2vKCkSkXfteYy/6j2u
d4gEtxhwCUufjdIbN5FvNDNXRapuW731/aaOlbxCBdHIzD9HOrRYEXEtXp75IPrZ
+ssC1RNhq37V77GjFmMwJq0zqnhGVuljJDLn6vBZqgcYRstpN21p0JP3QLQuySuW
gfQ1WAxOm9dc3qW4ETUtJfcUdPdaZQjMq7abSLrNhU0ipkdDff+SZqV0XaEXB1+l
t5rHSLMAvOc0ksaOfGJZuf1WvXQhbdQGSroHuX2KJuYQN1fzaUpNOq9Z6GCGOEJF
hRpqfPHu7Q7Aem7S2zJMAF7PKbt8hEokIg+KOJmT4lYrO6d+WYj5xh7GUqX8t0I6
woD+hpuwL0SK/LLNRcHDOUMNIxZ2gLX26j4Li3ESt6d9cJqUnjbSxzQlngOWNqLQ
Kgb2zfpM7fUt9AEwguKFd8u9bftWYKOpyqZWWHy2pUhgeAczxUQHzRY+h8IErMR/
OhiEh6Ai3BxzVjGDuYyGhaKsSqgbtd0Lk94dX16Gk2qez8+Q+d5GUJGkGP3uyrdZ
Xi3Ufj6fLjLuURDHf+TGbjEfD7N28m9yNBuzeVX5UKMBcnpIJhBx7M723eojNMiw
3F/dC39GWwj1eU5SRz4oqOA+yk/LZ96yDfjNXMMJ1wFGcuetD4PlFNnRCzTHZ8t1
nzflVmzAfD0iDX/E1UVfN2iwdLEK+vTSYf5pJeOz7GxrQJD4seZ4xDktQofXpB2c
T10xrn7GSul2ywHtPghtwKDgj0nREM4yAF2K6b5yciZ0MJD/b0cL1YDbFo//SrmF
mI6EkH+kP1zlaLDkzIeoa4Dm0C5vZbZjG5dKsv39AAX49HbaxUGOowzBORYQG56X
k94iD74kBJ+5WbQwjyzxeo8xLMDtXm4eGnK2p/t2EtvUltrLkFKZVkFyTwXoiVcR
U/dV76cMgJxDrff+PetCne7G1j4yFMHOzEhPKHc4IlEKDxoTQ0ECSM9rS8MxMReB
NgSi8PUB8gBwgixtBe11VicSEp+YmDh7vpFhWLveZbxNktbHH1Nt0SW0Z4upgA+O
K6tKIQhgve8cCRx9ZsDPwHNOorvd1zck0ETf74E/0SWYpfoDptdDhUSnLuUhehvq
dNpkHDLk+IIp3DKnRKahGdj4IlBG7SdP4alKgkaQhVm2cMZ8RhjMp4XEV23s89Bk
TUtVe4mkuQuGWjnGNKq7W6hj9UXfDME+Pb28vnQvOZr8dyKJOrkBPDAGv/U4wACp
YzCBgGS5C8/Ye0cynpBgTwCG5Uccng+p2mtrFvyEgnNC0ZzbilLU5GyVkHlxWicF
U7bWNBasFW6QjKrqqUE0DR5ZMfHSmcOR5vwkSYhEmpejDS7kviCTr+vl9sI/9wmU
G0Y3hdLk9DaNXoaq6uiCOpq15yGtZriEN6ILEqqYIUf09Es9EIzV6eYcinHzN0TC
EdRSkhNNWBG5m0wdVM3oTB5Jd4DEwBITxTiSmqmm0n5pawWRi6GWHzRzynrIVGmU
19IumKEZY3+yD9r9ze5RWoract4bhBtn6VyyhAWC2lMWTp2XvpmleBTuQD3L+/VK
CPF6cbpafzt+vNKsv86Rbai7R+oJFKiL2r4N3zHjbscepRIvrxbA4R6lZxMKOZqD
0GgvJUdwvqaHBNfpMAwDUigxWaeR6B/4FeiAf8nb78q2rWZkwt7LDDMoDxOyB+0y
MZ/8aBTc3oBnu7Px0dIGwIF1qUvT6710Ci6nOnQboc++vNUfhox/v0lNURrOyMXP
8pgfqrZoUcVn8BD7dMHUIqOYW6qIj93z9Y3QelFzymRXKucQNJ/v6CaJbbnO6n6V
xe0du6YdJ9ToADx7S6uSVd5hevQnOx2Ng/GaxvzEaHfmGVMU82Bu1rvALIt+iwLf
jzTPKQnk7va1OisinbJ6mOV+mNluPxyWUGsqEb4aaZQ1QQZWguzGCQfFGZ99zAEt
vtSMkavDHQ5DgSYBkBeCWGhx/ODitsfvkGGGI/HhXYMI826S6RlQn7+PF0qD83aC
aFk8WNPFEk+cwFwn/QFY50N9cZa+YwLQ7psgNyoCObKSiYmlpV7RJD3ha29ky9Vo
OzPZbQYn9/du5yWKskeJPhJJi1eNlWXS9txC8aaiVX4IrhKQSpVHvRJX37PK9W3C
AgZ6GbL2a+YGmUR5JcZOoUqH6xvQmnrGH4Kud0IVND6bqTJxfhvUfw43KhEKYsEO
lqhZTK7z7ksBQmucoFbzjzLVRO1g9zgjMLSxoZpxI69dPlt5Mxf9zmzl2azF2CdE
dpTqFzP97u4fhKhH4J0CE7biLh0Y1uH7CZDO8EOHc+YS3ZmnubOcjtohzTzO7waL
T6+ZRNw2EGSxLr6eC0q8uEaAHRFjEly7BuLtRVAp7Qi3n/Nn0c0s75L7qG+sePf1
wYQUJzLP+wH13vIfyw34BwVSC3oP2LIFa4pDZ9a6y1pPDZ9ccEu7CBRKCPLJ0mQJ
FTCzjvY+hL86CUmd8f7i3ckJWQhJ4Ix/Zy/4g8Y9N1Rs0MK5YHC6U2yno2Vctc/d
V8dni1b2ILt9KWEPDLq3fuk85TLwk7E2PGahj4/gVy6JsKlbLy/S5AVpcd+R4OQq
1cCjaRSuNpAW9vqZxgGxyHbDJVpu8AOoTuNiy7v41VMid56lsgFAk2eYA7ltN7C8
/BhqraeqKopRbfiF1ZhfN2Hoh/xqV/r/DbQJO93zmneP+ywWj6ueahKpb9sHvhYG
Qdmkf6vb/JXtM65PsksxANXRhY1swCOJ1TrWBe0BtGVfXAgpCs2CwyBkWVoPnDjV
DbtD/KYses0kDKgCDZI/fFVCU56qcNzeDy+AVKuSMcdcHTktbenTdzE+kxTDE6/v
Czai7tHblNSlkSKVUsnPcNhYb6pWQU4M51D76g3mZ0Q8fsmjUxniYIv/Bu26lrJ4
gpikM4DB0oqnupLRGsn7UjsQXeVIpPOZgQJoHZt5n99kXpI8IWGnxPjkRAYBGaSI
p7AJ8wykt7QFpq/lkshWMWuEXYkvFLMD9p7BXyRFUB9thPIKXcRJ9lKj8uDuub5Y
z1fMP9UadD3nxUogr7kWMe6Nkd+DbBAvGgsE8RJxyG+GwVJBYwc03C9HYc2zLlf9
bQwHR7NVfG3hdbvhR2Fwd41i0alR7ndCxbIDA/gKetCdoVNiQvZoBsnGIdQV3BLw
SxOu3gVG/zDaGW4/EChwybEHvF8KYYB701e+Uux+/WfSdr3wqnnDeA7dwW53prMP
yQHvkJqXwK0+zN6CE5x2eItqr0JX31d6DOjwjMi7/CBuGBXEyvBwtGh9JaP+T2e6
4totlKIAQIudrC8vZiL8KcKzVV30b+rF3CG5VqkJy1S9xqEvUH9yu+E0DD3P1VKz
cengrjO+Rw3u22uOhypIbj+jemhlSwW5en7REsToMpuyXSh3uDbNPJM/ycgZUSzb
m9oOIY0+7ODwSTxUZ6RPk5hM+z7XtPQx0MckMgTkrY5nLaBSt0DjWXGgQMj5CS4W
yDZEsKrt4wVLyTVUTEFMFwQ0bYR5C9XBLOTK+gtBvObTxbghpWk1ePUFfithcXVt
ia7NekSFfGTlWSjztWFyBtvmhNj2+z3W2QlMUcEA6tHWkuvTkPtrUfkpDzgqRMDc
QrDR3XolUSaJwSVmt84zIlRmnCjyc8qQ3uMyLLPnR1OWUq/lJExRQ4M/drEgGyCe
OA/JPlsllj/2rLkgN65fWptkt7EoZo0T9Y7pYHWI1lE2FgbAlH7sgKSLW1rjUmQh
rzVyExB8fR7vfib2pXuPrXukDmFgDgX2WAsllRN9KIJ/OVd70IQHlbkjpN67aBoD
HdF5n8ENJMHrJFsqU+khCCqb2qV7wrktCn0+2UA6Lr3mVOU9xKo0hz4fLuwBUyeg
7zH0oMwzaS2k3B+KOss5BKjRgd1hcCExfLi4TtMedJiUQWtZWKvumW5dXEqwq9Oj
aSldDicjKDzugSmfTzZ/PTbckx9W1flHVVtxVuJBag/0XiMUjwBeWd+6ad33NXGj
6gAx9apdCWeanIoB4L2/OgCNgIw5L4b7/dcZmI13mnfMyByz7qZ7K8xE6DVI063C
bid2+U7SXFWXxPLQ+Qaegf0Th4eiIq93u6ADje56fFScb2z+Q9iFFGeM9lpum3Ud
QB+Qhti5Q4nT32dIDYehT/QPhg6k0F26zzipMkFquTzMbBlqqA+Cf3Krn04Cz7Wk
++VFzATe00XAkb5VeXZ8fo/usOFozVu0bmegqBKJsZ3sEzOn0AE2WObNLUvbuFds
uOHhHOFozgB2jj2KLZvlcTODYKr4dvtf4pp2xBBl/4DdX6yqBTM33kfRo4y9cVlp
MF7eDVPr2kIKa6DeVQcyc34ioLwWmJ3Lq1yGHbJNXqD+yS/ftReMA3vkI8Fz1xvU
zoBXd/OhABD4t9HqkE4+WJMi9/4VFF3+ph4g07HhhbCq4xKk37A9oKBAv8wnSUmG
FNHYqEfqUul4pFlAwVMS1q7BWDNrvCQI6Mc0uBEqjAsNTFt1T/Q4Si+3YEeSop+N
DjHIAr4FZNkPOloVjLKmwjAT2xlHGBfMlf7RPAqPycTygj4C/At8Tg77619FubzR
F8zOxbBoMYWvng61bcBeC8qJU17hnf27EQgQvElSYQZVo0XFAxsAmtbYdtIgp8FN
hIR5nJ7N7kmM8Ng3sBnZUOj/rsU+iOyW0wbDi6I2jAYZZ84sN6UAx5qbSBvjpCCJ
pFn9rtID3KCvwkyv9HFMwNIu9sx4/6RGXWUp5w2oJCGVhGJq3d5e+QGYV3zuBMIW
JsR4QJJhqs4B/w4SugNn6EcJvMUM6H+OsTaZOji0zhgKhxo70tDMOmbfr0EVembJ
fuxTbK8Q2GPFr2F3DaIU86Lfkt86Ym3SAxSyRAPi1tFW/0TREEA1EruKQ+HID+73
rKU4/bToGKNFCYlaS59erQgyLcAfO1GTT+8vud4SifEhT/6P8gCdG7Dr5Hay0HDh
u4t8SukJqoGvTEtG0YEHi96LjKMPNEjT3p+XFoaZSNXOkzOTzOz70tV7isHJToMy
5jiyewlmVLnjLmrNkeDjSYKBdA9Zx58SrWoR9Qd9KrcUzaJp/PeKUkkc1cUGt36W
CPFr+j8kfrn43WFbtO5Cexu3Iq2yZr8csMkhMdgsCaPjGxMNjzD8a1YQAVD9QdWK
A1o6RqXQJ8drl0ZmrAjF0OwovSBVRoR4aWmOPBKkvM6aSiQwhf1qMTC7PEdqu/H9
Qztal8DMVtltlaSr75S1CAPyDAIKwIelVK+F85Jyy7ED8bSNFrpjwQpatwTIYStu
vZ8Gg7x7Sw0DG/UC4hwGeoTQ4HUTgbNM+0Zm5JpyFg6/3KkVLj2uojIqVYuDoVGP
ghB0OiaZ71duFtxfAmhT0CeACyepQUzN+gq5mTHv2aLIMextmWdvO22t7I0IIsMo
Un4DAMlZIUwdiDSlNAmoVqaJcHuvxlq83B1RlnF9s6BW8NFa87zTDzy3IEWynmnt
/a+iYcurGrxda9FlSbvj6LLzT4FpQERYa98YuJwZuFL+l7l3Bu5O3hAbUwbAJgYO
cFuzegzmuaOEkUBe4d8S7+PdpAL9Yzt53sRejGZklt3ehiPBLSK71fZwKS8D0vcA
mZq0PH+WgyO55+T0z1XLAVtG3GK2FKdpTdBvgFaQJH8Vqnc9RdyC1yQ3BK4qpVOL
D6KGdmRZkkdI4QOvu6Cjyep6i1DVoGLST6zVg1P2O0Z/Gw7B0DIJrQkJQz9u2PMa
5DXEi/xSEN/139Bf1Yrm9b5W4N0xYrMsb1rKzqkZ+l/QONi4HKRi3ZtJZ+hJzCHs
RzCeSEd75MJpuB2DIyVZaE1Bs096Wdlr+Pbtm9SvshimyWLrzFTiNCyLev5TaTu5
wv+EHfa7ZUR8Xt4e+mQUfUN9GHq5HcKopzacAK1rTVHnR4QfDgrjKmHTGpHX02OZ
WuaOw0o9kPblWD1SnutGEEe9RKSOrxp8XDgvyPse/2Un75pf+c7yKGaGauv1X9jD
U5GtejcKeQDfwKab54aY0i/s9g7aJOf4nEalH+mSN2vX4uTsDAKvRLZzmYMtsRQe
DvBUL/eQL4ce1dpeoT1BX7ez0oQiyHQsV8hR2lRXXERnh32wfjjSSURmieewqU1h
MGfvpxgR4eRD0ju7ZJiK0VVaHHVbZEzL7nxfLYYbZaz/si21SWYZfALzLEm3aMyK
WcKYRUSuQUILZ/pmltCfBgMwzZTt7c86ylWlfWyDpt070ij+rbMeKyUDTdxt7mvH
nGvLvGNfFugQhRM3DpCIXTMd2T1mFv2Yt5rAja4msG3+BbskGLY3ERsXbJ+DRDFO
58kKmW0ApfEzMU6PQqtEtEOGMi2B0K/cAiDDW1j+6RZmtmv17xXrlJNeSAd3CFg6
/lOZDz/Z7SoCF/rx5MO5iB1kVmaKNrCZp9fpcu/sU4cgHb4ULAjZHXq9D0F9qrQ1
xgAy5c5NKiillEXy8bYE8wkSL/oDDyao7DLLTlhZq+0w+M9wyn2ckMS1wt+C+Mt0
XjB0cVRdRVFEzGUWT0K1GTOWg/WHv61peOqfYq0H1BLjel9mMhyS38hcHyJjTKyK
XNl+I/RwpJYP6Ne65S5yHYCTPRtO93QAbbnoOW7VS+TWfbVPfPjeuAmZ6Ioej2hl
OiY2PgcMeHKKzdQ3p2KVEm0q5KjtQQDWeEJz1gf0waL2OBjlpz4FoDeI3wg0cR3y
Ko0BNC2NtRT5f1s4JHF89mMsoVuq1H2/O1CvPXgyITz0OvEvXeSZ6FYKP79YPW9T
4IroyHAgWP5zcoT0gf/f+PB6D86flL1rF2X5wwqTOmQ+DpSgfGaCmq+dTzBT6Ck2
fWm5Bg0KO4dMB3klACnU0fvCgFE7cKR3vMtiQ+PTEQRF0kiy3vHOGDPvFrSMio5t
pI+tx4NUBlcJaqPKyunsWwCTJLPUvjiOV23u+NM9+BDdKLs2zJduoaOzfjMVONfS
70zQgeE55aIBtT2x6BOAXGJUHCzf1Debf2hupLFlTZkbEoFzJpC7p9MLKuPn7fHq
XC0TmUXupIzCgja95Hd5y7oj1n2wH2F+oh5rPsD7+z3BtTur3WlVh9NgwQ9lDJ2K
UMA2EOL7sRF36IA5BiMJlyH/n4Hy4wBV9y++hp9yoqDOftmKlp8GJK4x7LlJTAE9
e3LWAFatTa7yu7FYLh6ZcfRXcMNG+xYDz7EC1BglmIHHMzzkOsYFPFuS4wVAD29+
C3bPZ1HQnXJTb2rM9y8CCAgzrZxK3q70kMVyIkpZ4N8bZMOzRKrUR/lZHwvHPzLG
Fpz2dx5sWcUaDdgPeW0THXYKioj3nGMaKqNfinb+WcOTkY30nJLOGBtCXVd37zR+
5EMEu6qyYHDu4hbvtVWc4kDTrgrvgsMfN5iwdhKxjT3nKGXffNy0bajbKD5ddDHx
BSqoTVwPPCywS4iG4MAtNmzDkTG6m+FDjsOh6pKF5PO63qn5V4stITWdMRf1tl+f
dY5+tZNGvlCG/hc2r8PRaTeqJ2gpA0goSayOUftafWT3agM/3OKcGqXTHVhBr1tg
VcYzziEHEhY2h6yZmXjqCpfcI7lWn9UMmsSV1LRA5sofp2f/243uQBDdz5PcLIxM
mIY/hkWYAEiDHxIn/FYN+xYhrKOR+TS+eGVbxHmkU6YdEsZx575akpvR+nRrEycP
yFR2ltUAd5T2dpc7G2oVhTzqGmOFYCWa2W3H7vpIFPEk/otT42JIfrJLuGaCfeFM
cIO1dde29bzkRnWYAx36LhCNYHQk/xUKAc9AuU+Cq1lsPJlcykxKKqvfLEKfQvdn
/Ni5VVv+gx5qpytPVAq5Mfk1BKc1d17KHzfhb5PMMzqkecqgMvcJhj/XphCWcDCZ
C09980oIc9oG8P5FgCqzK2lugG/KqLk4rqswamUKrCYPaP8YBEM70q8k1Qv5bgFa
jY8Kt17bwKmPp1CGYpoZbgm3rTo7xtQM+ADy7ggaRvojfdOWUoV3lIT3Ytmvix/9
V04KvsrfMA2h8gVjLx/Sc56aAq52r8LJOXJOGLZKDmRgvhmxrS/eXLV0Mpjz2dVn
euUDDukOj6G0G9EJhjPC+NbgMPwKjTizR1hujScRm0FqyE3S0ojGK5U4AaXnS1IV
fey1PK8H7ToAVk/2M5Gvt2U35/92BzL8uxEMdUSdkGulwau7K24BbLak1yFz6ftO
F0CQrpXxnIGxK+3yfxlyhteI6dcagQpa48w+UkNJQD6UFloDgQwItZk8qFPH/M+U
btZ8E3+j9Jt80qS5+0gmRXKvC5GgXnNjxBW0ogigQxHwLCMxDdJB19MiXSr8oFNm
Ckm3o2slk2UQpkIpUWDZyMLO2C9181ZXFFmmdJh+8YR+ASsEg3UUZIWlVrh5jXXO
PTEsEidvoU2idwZV7M5YnTAIdHG3+QQirvU+DDyQtbX1yjmMr2jASNAm3ISKz+T2
99BmdkkZ1KxPCrauBDx0E3AQ8iA4YR2j77IYX4THMThNOQ3gHKv3o7j4jNx1Fl9x
mPpDES0I4FEOdleS4J0LGeZmPvhJkfGN/sFatcavjv8JcCqXmaAgefNNU5hGivn8
H5DleUHAWHcf8u4c4WN7P/843f8GUepKC/hQaIglzpCI19vQmAqNhdA0CXN9PmRW
+a0p2LZXKJseBNUF9RFoP6nxRrVpyTGAroLSvsY38EKI+/V4dCgz+iVVcQTYnlKF
jifzQPQRcf5wl2lcLtEKdLbYrQJKbYgyXEdl6Y3cP4akaYQrTpmxMUhsTkBPmauz
JQrzBAVq5fMmEVEhjEMiBSD94VZDVyfXXP2io5aSSIXUOe5TJz7Eu18zQHGhj6yK
wvwiUXqV5jtmMykLMm3xMvgRqAh6t78ZSr8RUCNo3NhylI9jvRBdKNiNDc9GEcWN
ZtIZt//Zin2lNRxXfh49GX6UuKcBxKfzEIh1TUB6vbwvFG6YTQuxj32y5K2UWU+u
6Ipa1u0PBbCtFw+zr3r9JUnsRqqhfSa/+jbApFuOU4Avh90TGse+ZRpxD4jgTPff
6tqOMjBDl+1I+Grs5SKZwRtY4H+QOFBrLS2oy4uy3xY+fnjVEq+oPHanQAr1x1Ej
axp2cJomPtK2K5AgMSX/9EqQMpckR5eyBv9o9GvIBtazFfmxm6sg6xN42eQqRL+u
mnd6CNI0KAxz2C692B5Fm467XYMMHq7qmmUq/Db/soZFZghUSh+eUvIu5FNlya/s
5sfrpkBTlSAs74e9vO0EIOfyDmX7UcGNN8uHwoBFtfdO6w5mO+uPfbipdeUkXnow
S767qa9+AAoIqHlYuacVZYKwZMbQAyoUuPwUsZ7PxTyKbnYpbSCNlXuAJGTtACk3
y/wh5YxRN1HnFlvZal+90R6CgIR3eQJ2WFer4A0WH8cl7QLSGQQfaQo93AtmK6wT
jbXW+nnJtI2jVj8NIMW713hfaORYCVKrW3liVWKwA2xyvl0K0JMlKqB/1RGmFV+2
aSQ/DkpwIov30uC63O4mzaFbxxcasJi4ezAm7jvyU7Tty8uelYCpiUTeI1R/Ht/L
i1HFTBuns6W3l6B5e3D8YK07wDvJzRnW4kIz3RzBT0e2Emo7hcd1mciAhrpqE/3Z
Yvwb3YknxgiEnEP4yz2aVxHdFi6a+diyi4aVbit8hAFpduqYZUXrBBYdeWjLrlUb
sY8+/KDqFOfp/huLBQNxtIWKvXbl2MofgiXZnngPdwCC0aui2nQcdm8pJwpbkHfN
BTNVY6yBEnTM50N168owj/ksxqMoil2Mpxq4bUg62zm58Qub9Y2TSqY8NlzbTCSo
b6LFiRKVhPbndgPTfzy34deJ7wFDSgsvtsHCqykU3nH9tOTu2kr3wkIVE/o1tUUu
vldic4BFUaPfKtnVD0iC/oSMzBaB/Mr42RJAJ4eVRJKVkpy4LKALOwTc8VGW9HaD
7y3cRN1luOVMd2gOXly/hmdCzOICMDawfI4hk05b2VR8JKwm/VSGXPAfnvYntctf
q5p27qZe/Y4ioglLFhfD62WINiXvqU7LJ58B2MxvVJkIQTQ0HvneHA6EFo5WYo3j
fJF/EM07Piur1V7Sr7kMYeZ3DUIxXPDpYR1FKtFLCccn4ZXX+8LDIr5n0R27KBx2
OY5qxQSNz8mNgVw8tMdx90LyJn5DmKiaDjDi5sFrCj30x2W8Yi4ZM2b7+xHCCuEA
6XFXWmJa/lF9ayIso59Lk89ElpQ+zg91YAGUIWbcaxBaN0wufWt5ldq57WcH1FXk
2FZz+JaGJF8Ur3Fttppc0BnnGSdxzEElAL40RDttZQ9tI4vU87rTqzDLRcGZ5KXx
qFr/u4TzAb2v1H8yy3YOGm6dB+RGjnRPjiE2F+zUaFf22pddtLjjkGsF3tOipFt8
Fm0iuN8PVtbmNK72JB1ezKFcAlMyZbcEGqi7+aHiD8W8kfHc6gwy+3DyQ2O3f+sR
nVOgRHU0YF7EAbMkuYboBq/PzqLteW4cyBzW2gt0sNSekCBPH0V9G5c/gEazVcCD
ce51IMq1DO2ihEq2GBZSxNS8IZw9HnAo/TGXwKLk1/aylnaCzgJIZZ2GTFBH1amB
pgx8CdolkKUJsgdQt9XZQsWCjDIiGv3M/ThBI+5C1qAsNIZN3+rSrQKlYKP7L56i
o4GW6NevFey0yVAzCX6OVBrb4afoSd9KDsb3qf3xPdQq4Jh/+YZEFMcqTyA2Qd3y
W2ecSNHSTM505S2dMa3QPrqtZUaH+5eVE5qSKXen/fVpaIS30nHMCp4mRwYIjKRU
9q3yje28TcjXx2JQnxix/M+6jGxRewEPRWO2Lgh9tJk3CEbi5stLxaXhEnQ7x4F4
sMz6pZfo4fzYhtOvoUWAsunBRkEFYSFgi/cXmnF3Tips620Ph0pI9U2ZORtz/KYc
V0nOM36Yk1frS1JRodrBZs/ZYP6jNdmZlnaIsqwNl6qF05UUeAJ0a+sjSAyfsi2m
JHofs2ZikQWKIW3aDhkCzChEtB4EelHJ2NVlZB3jnEI5Y7yUOUuuypL51vFPaVKP
hIX91/VEB6djD+8E/r4uC8tgTl4NY4LYp0ATCg5rIMbbL9rvrjQvstwp7Lp3lB2q
L/FZsyxFHMeoWI4VbyZYt5sB3On19NV9W2nLVgjoUAmO25gf9X7or668cHhg4Nmp
d9Dk2PIp2JV4+21arq1Kl6YXwzLVpdD621hiPBM7rGKDMC4ZjN0sRAjLUrdkJsYI
9TUww3nZB5Siu3V+5YA9eyKVXFbtBKkDOjS2YbFR+HCRHR0XyHoZaY0zHjJRdAKN
BkqGR1vQk2rzPZgW6nH6d6sSjr7JRmzno779wvua8PANcQXrIJVBmaMK/OgAFjQ9
GkO+9Ez+Ff1yc05EyNQqGr3It1RKsqG6xbLlszmsv7IUMngqSOJjG2SLt1Rs2jMa
GHnK08EGP4BAW5yEV6eLbdxnHTEjGZMjZaSZ9ojdLQiW3dGG+aS3G+25bVCscj+x
NDzgnlpapQiLwCkfyq3TQdkDX0ExibINM4TDLGSdg9dZXZjoSZ19GFjNxKL4G9A1
kbGOJkU4nYE4cZFjKy3Qb8UXo5ECeSS/rJx0EzlivAmPBzzkw5/cHTBya3Uu30CX
O24JcZ4uhZmX3uBr47BPqJFAQKMNI40EI3AmrGOOzj9zKS2z6qGINtCQfxfUgJYs
oMV6bjvoFUw6O9u0rd/ci7+Ao/w2fJIUwTmG2HaKOSRis4l/j4zN8f8epSls02WK
Q/QzpGwvKLUZT5k5eT1+weWTMCusNL+5eB5ZlVuYcmRGo5ZS0Me/PTdlZz27sX4I
+BQ4m1t4UyckcOMxm4OLOqyPwqXtuDa6V1q5TP9gwSYuzHNSdl9k/7WQ+FB11aj+
Wztk/E0G69bjtupTDGjv8xGDjS9iUCwYTG8ed+7kYvQSqsPWtNiduazDcblXUaGV
LJy7Bcb8iTl1SUEL14qZ5RhWxBC4rv99Lasg4UzH0BrWfYOsni97h3iwmIhkjU0l
fwR+vbiNgULm09iNvyIsdf6/u+PG3RbbP3J/3MIJ+CRMbLO6rzm4aiFBzU7PCHW9
FvCs5SWzUf87445KZtKZz3m10LD9unAXQltXdYq9IOwJn1NwO47TLyAu98IkErbm
m6tkTQjYni78tSAn/Vwq24nyYPmBWznlJYhhTIVXHkkdA+X3mpQqzh5rJAwQsSc3
7C34WGcKGIS1IduOz7uyiO9t29i9wzgIov/o8aoSBlMVjUd9CsNA3PwiKz7Zn/5J
m8pbzIbCRgzXx3F3NZl/SFkkFZTTpUjaOmZSlqhCEaVz+7hDYBOzFeaYhGbld38X
y3OCB/GTWRG20s4pxewUBXgknklQBlBAkXDIlTYO/Gz7WUWLoKBDFSsia+2BVzc6
DSATSNuPmmK+UptAIypm98LxeIR2/Y2Qqh85/BBnexsprJXWA4aUC8dbI1mZsusq
Ahpm60uLkpvm4FEjTBUIQ1dLVn18WC6jp3mnyCdXSaMsPKYAErWT0X3NP0tyXbpg
7BgDa5aP4vxV7YUTxfcvZcCw8R+vrESapMt0TVXXRPR/c1JoV+GAqz5zBKukTGfY
55T+vPg22p7fxLcshjTn7X2rf8BWO9pf/Q8MpJug6rP8Ef3cp8OWbfzqZ7rsn9sI
sGos9z9Ydu5sJ/q5xOhJyQyWD8gnnXIQjDNocCRvpuPxgpcR8W6zOzp5YkWmiKJ1
H1EUKrp2IocSrZlciy6JLYDer0R86CZ2cChBS1bRaMiLEd2jdXIdCLRvzihcrvds
65T089+GawFOoXCI1rLayKjM9EIPnhvq781iDzHZVbRHipt4Su61GGOmzUGyDGz5
y4dcZ/Kg21RBH0Xypp+Emw4vrKsl1kzfHeHlPTFoJTqhLC8LJOqaPF+bChMTpuJF
hhhb2r8QPHd//DbZ+RUJnHsnHSsThOgAxME/GFBpCBdytVnxAqD5RW3zTKkKuEun
ul0X9DxtSotDfbRXCTd+1fk44V8jNo+3TGKSIL8yrWF4QAhK3sXf5RVtepvDPrgt
q0CpKmwTAXhBoypFg0q/8yFp8MQa8UoHwxlKnjEo/Ls/vT+7G32XTh35/BD3d0+t
M++qOxfqqAscHNlLtMpcsv2VqyfKZ0a8Q+NrPhv34dD8s0rQEhpiCKfKR5yjpm/q
2COk6eN046ufRFtOowPb3UiOFM8rIOC5z9YCuf5qCP/9N5ftB7wMZzQEhBfvh7Tj
PofsG6ZgSm6M6BacKlYXNeXgHaiBx+6uMJJiUYglixkCrc02dJ3/GHjMTKJDBTl1
2Ppi0MD/vhC6Ofj80EzEOpZLDNc+p5GegqXoxRPJTnWAKS1NoX4dWvyaHsjgXpn0
CntPap1oy02duioS+Uy4EZ8FRGkhotkIm0bxHmQn061yE6dnjap878zheh433h/o
3VIi3RjypM8tDWPhlK3WrgsQqm0hFnebpW/t3YlNFmhQmPckHzs9ibPmNQPd/q3x
1WXUBqwTFsUVfi6dPduMpv+SnmjDt1NMJta2c9FQAOpajy7eJFeVKpTIbEJvI5WW
7qozY1P/MF7+zY6ipMVQvHUMaQzs8h7zk9oN/t7y6IBraNNJj/+N7UojUDRggAix
lPsiMSxTPn5z3foMaAw42DbwqsJtgjiy0JGizXnW3BLiJtinclsOliII+YXDnj3e
K8ktuZY8RWFHDgG8Nl/AAcwhGtbZ376/5to79eaQkf2HJYKQIpGEU+vCnlg5ygPh
VBYfglC599b026qiLpUsk1v6jGoiIao1ZLsnjsXc2Kma6LplAFuslbWBtmJFWt/f
RbAeOWxZJEWG33m4voRmBstIxImTKGB9f+d6EHQYpaRNYnOCxhawGZcK0qw465nw
/f2MGaE/y7tYbrna1ilgh2smDBzBJfnBlxzWQPkL66O4lOW/cZmHlPKr/3urNUA+
WtwafieKuCrIknRX8GKVvbzBHbn+x2wKspbJ5wnmu/noWGaMy9Z3vSe8DMaugAN0
G44zNB3E4Ql8g5a1AICO2oE31fNNCP8Xf522TbMq3ifaYPWRAKmY6hEhJe1JYDS+
T3IPHpUFxeCC7MniXB5n0hmmh+vAs99BFve+Ucqh3FZ55+NA0TrK19wmDDAKcHs/
v5CH7h0SBe7T59cTme4vLFb8ihE7OXW2yJp8P95jMq6qTaEN3qbsuJ5YrOBiuhHv
hsb3ou2KiIysCF7f2HAeyCqVNreiEfM5eTyIsy075CjxsuoG1MNasnRb7DyHf9HR
V36KQk762n8PKyinyU0dgvnTEIZGd5BgdE9XUUohGXOZzx56wLL/KtmLoEd/MEcW
SE+7RlsKtLQuL6C8UlcsNMbzAmenSimrDb/0txUJoFlOzvd3XOZPViRmyl3YUpGh
+raA4Zh2f+9SsxrU3JDaygvV6Gy384WKHJxAqy/MZ6rtIUYWPDet6F/rrve9eg1t
ph5lseagjPjhnOsy6u6rVZpSseuXNAcgrmDOv0mUQzb5oIPEGMU6LFlME8jc7OZc
qW5Ey9mC81Acu1vKhqoHDAOxOvJ2MebaqtRvK/6EXkAoZ8/w0Zm3Nu6MTZBm0vpD
KMXVDdzAMPTm92yiG8FQSx4S/m4KZuUHWTjvdBv+zc2z0iiq49JNhJxlxggLt6jF
+9FKYB7fmZ5LCayIwlWsbpLNGZExQcXAfUplUd+yOrrt12JBLMzulhgnaS8/gz7T
RMHWSPc7fgdRJuwlpuW9WaQTttRnXxe01fwBjvbeKmpU233IV0algdaqn6yovIHA
pcyJGUSe2plgQIdxaADlGHoBMsW6EL1IYNH0s4geSiZPhY/l275EELbI8iSOY6GY
71vfy9CXEmbRFFpl90XWeJInIATZcfu57Em7L2sF0ti8N9cCJF2EAHQ4hkuopVeo
RpFRHptLel4j1kAIeMCCFoB9ne3ip/jh++IaT8ojuqkXzHTRBenU5NejvV7TvoHG
weMKd9qs/cNQZo3L/QebhQvT3Parl7iZFLhcK5UJsz0/iC7y/MlRKQTG2KDmqMN2
Ms+1HF1/PuGbVJbbAzozNYnBFePVHNYc9S176P4g5dx1bduMGmJhf9dqmahm6DME
U2mC1+JYmTahvCOpU7nIpRGhgki6KFiQ7XFnNQHwdpyGoppokhihSekw+V1ed51k
NsdPw5p4ZQMm8FQnE+uojS5E0r0WkEQLEGbsSCwUwgmTuYwZR/ckCBFdfDQl0aEN
xiap/u2EwO16/rjkbwn5g8jibhS2jMTTPVBJb749gXwXd87ojh5xPeENhkO+761d
URk3u1h/aBOFLSCmyUtbmVdKw3ndZMBpFc25Wyvm2HyF0O/mSHdJV5scdNJtIph3
9tyaj6L7Y2g9SYcRsv0/3q07mFXbwvz0q6wXwpFXjC+955ONjpkgQLh/F+uM3bWC
hJB4QuMzLtRXNi8p19vo7u0XlMizixsDA2VPSvsReRXeRt+wzblhKL/sYnWnskNm
02kHiYrCP30H/EjQFHEJYZvnQ094aBILwnqmAbzzYs1gEP/7UGM1odtTpxoCC2ZP
hBgsjRoa+ewsQFr3S8tNrgW5YUnwqRi7yWALczHZePTGkenaMEyG6kfuCOYjX7/t
cMMh4TOLNUVmgiumZ9aoEyXS0J+UJF4niOCBDCAno9+TDOpZNOqEBAoUtJRfkpmm
am74G/+Bb66f7KsHdeRJps4B6mUTfMEcLLS0bIBAkOCN/+Sf50tCvcrLtVsyP302
r8/werv1es3VvwmOMi2T7KBTA+kNHaD6DMfq51zEOQchftchtptrYJLDsABIEfJp
z/FfMu5MZsShzOo1feQkLG8em9xgaB2dMqm0PdPIw2xC5nGXPLw5wghLxP7+CLe2
49Yqk3O1/EW5Sl1KCvi2ah+SR17tbXVEXQffH73XntJ3JVUp0Wy/w9Xbni2duu5/
CQD7QVctEvjtKGNuSWacU0DfeGT2bpP+2+ipAgNMGLW4STbqn5oedAn3FS3af9M7
765eJKIoTrZLhINOT+fkw+u6ytq8pZ9rk+1fmm9oH7f6cbtvQkGuACaVHVrDDGUt
jswePCPJG/E+XEH/VQgt/55K8kidav+D8aR9rm9wZtXhfwBW2V+0xHCK9Q/X3+Lr
/R8RMxjlyb4TjygI2cIl8+t/6tCoNG+blo0QMffGWztAauyAMZ+mltArIsPYbQ4O
G/sFqHQZ6YKO5GiAyObzIb+lNckDw56ac8ml9TAJRGwV3lQFIqygNNEjLXyxkqbT
W0YzFynFBubTjP3BjPVTxH8OZkqPMkCuJaE5VeEWMvKoQ9G/feLPVgyZ36+mGjeH
4BW6lDjd+0ac/ZK18RYRep641ooLkyBRQeWF9peygkcH4Tj2dfd67NnIakR7taZD
qeCPdDgCS6dWYSPKzGqFBoxrFsR+Yji/PIe61cahf23gwhL84AY/8I4vEmoHomW9
jMzuA/c0sIrAXwcOGjJEn/8j0v8SqnEe1OF7KI5oRi8xq5Qf/GP5NcD1oFApROot
IrrZtYbdV/8jrmtUqts3xItXZouUMxvtqUVD24XAVbJ2C7LdUS5+noUKgPYVTPha
nVnEWkjKieh+q1kvfqCLOiRFvv36iPdnKUwTuM6vIbyKOOaqA5omQQoHpb3bHtab
m+fkEQTOU+5xdOKJ+njMunzSf0L6X1pafr1P3WTb5b5Q7hHiFbzD1oD3Pjqhg7Tp
tq2gZcoFVk/tjvvnWWi8zo4jpRzqE399b5zH7D0izlwgiyDt3ohAZIVmk3wWLWgp
JCzWKHuQtoPUHUk8MMIpYDkq1YxGeP4wshH3kbHGfKZYXYUdZmTzdSnqN0nEsA8e
gp3BbpP3AKjl4caAWqw8EzZGlVm6/vbE+cMsa6Le2IJINbP9mZHcLyMlFnYnq+li
1swzgxj171TqHNdCyVLUqyHZw1fPtCAedot9r+mhq/dRPxrMcVsI5UosW/uYlyzK
xEvl+MArzH59GUgHeg0Jf0VxYBdwx7BbT2T/dVSKEuaR7b+PggMxx4lMMECVxdly
qXJOHh/iThBIaEFW5hTXsuVMD2y9xUPiDlUZbDIj7I69ajx/tbNjilgK97EJaInQ
3E+JbCdNWnNT518hrfWvTlSIg6N5iU8Kx0PuZIiMWIv+KqbaRi8k3l0ibdMyAm8R
4QSYr4YUSDkSCY4pYKJxGkvv3Zg41NXybtJnwYEowa9D9Y06ORjHPHRwk6AHCCZO
eW79TstDyqb8Vyq4O2NNmPrRaGFwPMXuhuMYp8nPajxCvDMzjuqHJivsMmBoz7EA
CLUSdWKd4/K4sbWoxzizAI4xWamZOhH4kCNNxJkjUkpnD2HLwWO6u7DDMk3NGQQM
z6RMOfuySeNOeM34WuvtkA8mkCniVnr+ZmWvzj+qSwvLG7a4AVf8vYmRB5RSJJvY
6yeLXVEUhAtAc43/hrgZAMsxw80ogMS6LloGBlB/AbLwDMz0xqXoYZPCUF28tynb
fBUtPWkoLoRKFy6rwxhe2YLswotWHZq8/6XTD7c9XfkW881wmPdObfiWmmI/Lu7t
cTpjIzA3iFUe6Q2MSHXjl8A3/UqJByIydb42BOI2OplXi9xis1bccfMI81ecJDUE
OESai7SgGk34dlCd0dgZV8+4LjhUpY4vSfUtuP1E4d33+QvV/3z9Jkr2ytYfM1iX
fOzZiAbW0sze5pd/jVLKitoY/vu7uZYIvDe6XfBaEdkH40GkwHLErhyOLQGZ8HKo
CxnhRdozUAP09FOc6+dPykBhCVAzppx4tMCVWSKlm5hfnC4vCYYNpHDmb3juHEx8
U3Vsj9Mt6u612yeQFZ4fiE61Xk/AA9pM4Ium0HvuPAkrAdUi5UngSg20B6U5cYSw
VXwIubEt24HrgiL9GG9GnvE9WbB+bxG7H569EhEYjh1jpD9DugQwFp4n1c0ajtET
iRpEuhf39u1omgVUOj2R6QvGcp62Yutx801rd1rjVYW/cYcjU/o8XNzcWkwcCGEI
kal5nUrNlvYSaDnQIWeuOulLwFpi8NispYzghllQfMSuICG6oyCDjCotaE0Lz9g5
Z2ZcMIcLELxCKZFImzmmZZJItYCc+76w4rUaxrcrcK+AkOuW8pqhU983GxvjYIXx
WL7W3Cs4gvuvBo9qD9aV/cyp+tKRu4SecE+bJEArLTYckYl1jnm28wZ7Nfs6BuSj
u8y+C6cxIzrSj4CgWld0dA7BfAxql2rUHqYH/yX/U5GQsmcw2G0O6BUZHzQ1x6cN
65MP+ggOUhGKoU9oUPEvPZERya+YJtTxYj0wsMdZJdQsUFsaRbJhzwBn1ixjiQ8/
2x1W+vG4r4zpLoAs+MwkhVyASl643IOYg5CVm+xhgXzdM0/lhxEKyYZSxXK8s2iI
9Pbm1hKKRu0bZPPJ7rnZeaT1TXhKytAW4CS+brNmInuqeBUGVPhVT58FUD2zpt7b
m2nIeOgtq49lgaXGe12CmTEH0wI1ytnMd41PTXQNRkbqcbNVoQ+jLCCyHrjNfUmB
cN9gR5uKbabr7tuGWwqlAcXJqXZwsFckwqDtrnPOoorfsEO/v1oLlUyWhrG7FO2+
Rc7WGK5QEBIIZvABFxBpFVe7/fWjZ8OmGDQ49nfRTHVZrI5ufutitYY/N+GxabCE
yWuGlbaeJgKOSviRGgDIjfg7Dh+oRq13jQcdLsiQ4mybegMu44OYPTJmmwMrcwXP
O1CqX6jOarOsse9V5+8qf9J2dzWC4UzRCuREpDHl3Kva33iOt11E37UUc6kqYOGs
0FIsQdY6SwfPePCsiyFkvZ0h4RtZDduZuqPEtsmU2q1CAA0yn69CzpVjBkBJYTvV
zj0URmq/F17HLyQaomK5nlHdzhctKLWyEmgB4OcYAqUwYz0IOlAq1iZc67ULzrom
1J/45bfclMYBiE1nvuNwWygAZ2FivOp9zi5bYR9+vgu6d0qTVuIyz6uMmoeOOz/7
eM/xqTPVXXORTzU/slqRLgXAylsFSyZ+GY8MZL9Bb7/BMudZtymsaRPMTZIgtvXm
3mccciqkRj3FcSkiBCIDNzmnY8sAfr/xxLdrrbghvkq0za5bwtwxQTT6u25nCgVV
wS3oWKI4QWr88DIH42mafuGihw1I7MPS9dkv+60G+VaDnk6HQlDfOewDq7XdM5wv
khHXL1HrZsUD+JTNbEuO2yuvCRQOQU48Igz/mVSMPQx21HyBpVUsWURjs3fBSw1i
D4S6kdCQQ8ReTxwmpai9aOOkJU5Lqot42TlxyJrgY0WdlpNdAEZXXQ/RESihyy+O
FX1WRnYx+VwT+QdnNt0rX5zS5M/cb52mA79HYFbvAa7T4oeF+jF7FBkHMluXmeNw
jRkwVC3SAdYNoI+9N28SCg9twwO3/Y8I3qP0jJ6cTBv7nG/ZpgEDncNvbFIcb0fl
RV3wgzVubzlE9+ssnV/Sn3N0NckoaUzNNQQ91UdtwSoFn+2toBsJxE4gf+XnDBmH
LFvkyL4ydU8Zm/oDPR/zsSo8UpfCkJGNj7I/0vCfSy1aTPXfTkFjbnQuGxOX3fUZ
aaBaPenQslEkcOAwJ1PQtrwbFKgCFQHOUwAqbLD8QWRCcbcVYl5qtGlMo6CDu2C9
ti06TEZ27+8S1tV3C62id0aOMqunhn1yROgiWrKWlXUVhOnYBY0m7twHOOqKjOA5
7+etHbnAs42frCG/5sXfHjEGQRuCFJ47UUAaARTl+w+rcHiu0lHgo0cccyuQApbW
HmUYP7FOKiH5AOaVsi/h83wpG7sBKbV2xuH9fssH4SmGeAQR9eWvXunqo3iHR0m7
g4GfnfYFwEJFtSLLqZU0/kIbsCvO4Qal5oOsUpcd3BKSWlueg3gaGuOc2qXfSHdH
RfEJ/+AHMIZmP5QlNIBxHtGGaz+h0zOwyJvKZWsc8NlAMRAhZUhDbKm74xPw+bkn
Tbjf0abEW4DTosreDt/wBGUklpO+O+LH58zy91IyEfESG5vVytMOyrtDrAzcxc1c
DbqtoFglPpYRLuhRu6Z2os45Kotk/yf2KVmlaKaQ+lehadc75RlbeUOaBGgtDDNw
Z6T0E1RCRVPicEal08SPw5kdTQFyL2MTrbfk4GNRMk1gbSWKB45v5qsLHL6lQqgt
hRh2xrdDe9AhMap97DolJqW96RFwEVF5br9lSAoJ0mjKJFnL7e4LlvzwE7wSvxUS
lgHLFxVkHVhEEgEmpSWvtoDOS2vfGk/EVNtHAxcA5dfK6i5qfCBPTivT/vjfyqUk
ANiz2mkCo7U0fFlDBpb3rXLjL9TG9Vdfs3Qc/jQ9aQeUsx6fCMa51DoSI5uDJ0o9
+dLNgmhB0Gtofq/yj6NVHfaiJ+vlhjdh4YCsrPrWVxWs+XnYsfdlZGgjVeV0YsBi
jW2uEZ/c2Arlk/qt8ylg2j3YKwoM0Y9hSOHdWV44Z0y79GZM2k1TgV/FDK9SadQv
pHFYgUg+CEuxR+JYm8vgYWIJ7Ug+p9baizICcfaFXpChqAr2Q4DoP9Iul4sfPYwj
E7UgrLGJW+AEJ+lQ8rRxImAk7/SmmWarpagIpQ/p46ywGYbdy62ECDnFoq5YZGVU
6gZ3cqOjXDyuEdYmvDpF57CCzhJiHhPsSJC2EVjq9HftrDIdTveDsLMuhRwbFeRw
EJVnnmjHBglkB5Yx1tPB+9jKs3A82Fpzaba1PNZQ4pCEiRwKlwA01kbqxW7rpNJV
o3Toyh/QMGyZgSNm0NkvIC3mTWqEZG45b7Yn4SYqth1OIHhVY5ouRLCVfp58Kww4
FO4kOShygPxi8WoEY1nTlD0VbcQVkMclRrmLb8oovcJXIT8M3KsR9rCdgVxcxDbs
/F8ZhgsoqBp3Ui627WL/5RS/w6JK2cIQbLANY1MpdWiEA8oRMkSdoypV5ikslbaz
xtwINWtK2l7RkAqw7O4YqjEXyGh4aTOTqdVRsw6kMVWFpThWzNkL3APLobwRFMnK
P/G/wce0ES085i2JMtVakjtGY/ZfyUon+xk8sis9BJ9Fh8PRD3wQnhNH6Ns7DkTD
HgLTDccTSyR20c9hmmgmwml9oeUcF9pCkkWq47DSoyuk3c7iXGgesU9wmCKQXlfO
JqLvJJXc/MY6MlsKCq5QpM524pQ2iaOntQK33qz4F1pbfjI9D3cER10CJlh29LR4
SgwA6ijLtH86YzXt6FbhY5hOkn2axZd5bRqhVNhTuTULtjY8VTyXrFcDmzFUfmkh
AMO6IQDj6i/dzRPoJAHpirp25C00Ub69JDQ23qDegGyjzIyiSMEKCzF6pNo5Aeyu
fZdgoTeEV2dMLdOXNYdmvHTwQhphZVG1yy0L1XubfsG4JK0TJiye66uYewUWskoc
cCQ1l/Y9esshvq9XoXlr+QUJ0Hlpn7nOPr+IdMkskAdaeY25txG6WmZeArPz9S06
UupkzvQ75SbZZs4x9tWeHXBGiNpv0cRHbkf+FFK0oQftokvi0tbq/Ggk28phRcBJ
gvkMsYXJC4y9xcXLeAVGlb1zMJHWbTj3iPAKJc39r1aq+rniWjYmtIynQAfcjfQQ
8O+8eZpeJdRZbVKQIXVHJtF+DZ1btWrwfxQYILKN3VU/mmF9m3XNaE/BkCHblmS9
qTn/Mz62yDUu9pKy3WL/dpGebTQcmrdLLrTC5rnTZc5h7dw7dRMldAIW30ulStOF
WZFArZgOx1UqcpGTZM5gdYgPXRiwJFkpz2DO6jJx3wVA/g91iCco7oXK6V1xMRp0
16mKKGMN5ikGxopEfjlGUIcCLtdLNx0hl7XmQSQmtFCaEnZv7GqwZg/2Zh2f7j3v
hU+Hzj2i/bmlFN+7J26WtGk3VFq+XFD0DcpC3urcA+pI0HKTKVdoWOzIss9Mpyau
AsrJipAkBbaPH2q/IHVEV6pcBdL5q20Ir1qQC80m5Ggy9cT+N0m9kLaqkpqSq2v3
nTOYPLI+rViST5kwW26+h2wHsCY92yfQKBBVmBZoCI5kypljsUCbPN49ThXDxuF2
GpZreL5182x6mtkQ1zr5AHEf6MJyEx9+N7ziCweVoMr+Exkp/1II8GTY9axd68ZS
FsxJ19ukz9sTwJU/jtPWPHS42CP6/Fuv8JZSFEBECJoWQ5MWH/NN1xABH0Tus1yQ
NUV3c2eHmSmjJ78evHoWRWZsskGp1cvNJBAuim1unKTowO0nzbn2UFlzwRaC6LAo
0kSCUBXDE7TNo7HP2KVwCc/QXVnh/4T0bjN5cb/TPk10hQbU9b0pNFE3M0NORgEG
v9BKtNh6S9/63/Tlt1M2cIzEmiFK0uKwaOFd2/IlOImKPn2oozoZatTJ/7/j9MJL
v1VD+okoKQ2u2BjWRgQEJqf7U1C7BUZZYSKmBoPYfuYPuAGvhnSXLDGrEiazx1l7
LEIKp2ZJDnwJurVXKb0+uibZ+7ajj52Zp8gcGE8WDbTVFs/4DLg+Vxs8/hoxqLzx
SOb77tELOCr0wTVIguvuTmWqgJ7X63dAtD8gG0EH2ME0aUDuReBN031fowXvCiQB
Zf6cnas9WrBXM2Qwpbct41YTKA4qpgW19lWD6LWt6ynIhM/bt0Zp5gmMcRqTRnkN
k19MS90ssb6zoHWIY5BbNKUjDJNjiGn8XfT1qSroz1opF0qVhC83qU7BOQhrAH2j
PEVUo5Z26kyU1d/qN642Vil/ZgZM7P0dzYfU5fGPzDpS0x4pTrPJ5wiblCrXLdbr
AckJvlrbOwMpQCvcnZHB56BmtRJpjTVV6x5NrDxtRu2pijprt/WmFRyS/7R5YiXs
ZZ4Zm5gGNnS3gDKn1z1NaM4ARhV1Zq4nbdfkwJGaHvryL6Eil+qcT+16+uybv8HF
fLlGyoR5V6AWXxctU+S5+Kav+znEwYfei7cN2+kA4kvKpAEQIr6YtJixnQaXYqDf
Q7WiKtl2S9/d9nH1HdAp6Cl248LK397qE/ptassaJPVam+TxYVaMHoV5vO7Jr0bs
1BR/h67++0E3ZPCl9nvRnKMiKcAtCNf7fLQFf3G0oxmLUepk8TCk2rQYgOyJHjaL
1AWUI9Orectdnrh4ObBYNl/eZQwSKgPwbheQJhQfqlE8k158XRMHn77XIBAlcK70
mWYnwtFPfiCTpsZoFLRbfUM+2iZFtRdtPi6RW/PU9giANfWAk+6W7d741aGVX1IN
IW/FYITGjkq4jKrXfPmdnukXtIuH8fa6YMDtd8oWxELDWe7PxYM5Z/cli99hsYVK
grOfOw8TOWnG7Wz/t6tPuKChSnRnggp4IekwU3hRl33hV2Wxkv0jLMTHlaVzNPvr
rN2dWcTvn85Rfeai7J7OOyLrAv6lRE3J9lM4Y5I/Wsm/LwHGkAbNld8zRGVrsFMT
s326MOt9GtkAA/9e65nyih/KZ0jZPctitAm5d/bJ8drwr5hqcaId9zRW4/rIsS2Y
eqvqZhf2UoUb37ouP8BHLWd9Vie1OTjRy6fYlm8WpWk+Gyf6dRBMlcdLMjYsIgvj
mVJ2deMg28A+cAZ4cLZ/g2XD2+vaeVcnl4l4sSzC4PTSdwuxhqqorNbF58hHPamo
LL7Ylzc2S/tXbVawJate1/p/lX0Tt2LHzMcKX8oH0/lEPdKjynwryxZL1E46HH9+
Z08/0Thrmgx3gJ1gOq6XTNYQCyP/uxwz+bJoby8A/8N6IpdeV+x7UjoW/86iMalu
b9i3wDykkoBG5tlOkeKA1Tp5yeNUBSLW7DCafHxs+PliTgfvUr/NqFTw6JcOBU0R
FK85kFT+pI48LrRcD85zUm0fdswxpwPVnIiU4axeBe1/yvr/MgQ/88EjsUwCgu6g
KN1DEGeqMVHuKCUZsU738AWKyknMIApSwUYDvRh/Ix2dc4qrHNY3yEAsr35ie/k/
JezRe7S4/1gtvBenTjgegA4zZE/i/YpmphpzMqU7XqRAi4Dq+PGPkMbKWyX15RTd
e4qB06yRzOHDLUkYbaLlDmhs/tI7KnMsy9qfvM+CXwwJoV55M0QPdTRNXDah10Za
Sxl7EdkARoZutL4qT0McHZFlZaKC1F+3Et3rsXMMvUnL72ycq3BVLjiObUGik2bb
t4ut7XLyuaYYXtlY/bBvvRbr9tftNNNDUaUY9ly7wxKdPB3YGw/Hli0HHUuQ7kfK
ADFN5M7b9ng4jlOzF/xwlr1J7c6YQ1rH8Ff0IGtSDugD0GCrWxQyokw7k+xiUIAl
9/y/6ZtPXXHCUzAGqqW6VScB9emeB+D5W0JHLeSg3dBJrAEP9CbzYrs5TTINPKRF
zso00r9DXbiSXMNelqCuLX4PKVs/PBTMN0QZgOz/sX1ZcHpXaNo/P/qVHvZBZov7
JDxC/ejLSAe/u+PgQcexZXwyAB4HOwAfPrRTDb65ZgUKKJDm3S1cMvWKe7MlUueB
dzekePglBoU7naJyAsDpEiXXlmOUf6xOM3k2gWmEEXGD6qCrmnEovpJJ3Xge3o6Q
Ffm9Z6J6ybJTeAXHO8+GCwV94sx1UD/YB5Ao6ltoX7h9JSsNz/8AZNhqkt/Oa1ns
/lFP6egZBt46+B23+VIqqgzc8CS/NmvydbOZXtfOaYgNpG1jdoLuYoAmWuj9weQs
Dpj3bCjfRntm/7UFLbJrAQQ2V60Q66TI21ts/3nVT/oSPv1NcE5apu4szvOdRbCk
+YXcq+h1eok206phDIq8LBJgyn0XN2PvEjAqZnTucPgPU7y4Zpg9kl7Yu4FDTRNM
qhTuWcjm+A4nJOU8KB8SifI1wwTNMk8qpFUSej8mBR82+dnkrYETRGH2wFYOYbKe
ssrXK8xjYGq8GiGiSYRXC0sn++z+PHoUmsVRpf0rN59RTvfrantFs59msSaFpj+v
g1ttNC+Pt1gjYJHcF3whUntuHEQc+sk0v5rDrQHcURiLpiO4T3bj8+H5B5edQh5R
FN5jlm7K4GIizax35zzLAwYRtx+nccQo7D0q4BVFU8gZPHVTq9F4P54cD0/I3RiS
EfiusD8Vez3DFag3lwQJf3X06UaXObyiU7ffCrDS3RT7BaAwEJNyDHzzqYmWQ2QG
RiL3iDAGyQTy+2QgWvK0T44kuscHUT5NoXPaBlml8HmJYNJkQqJDxnaIm4D97kzB
PluVsRUyxzsaKWMRCqw7xKJocFgf50wJU93JdcsjiUviCYPkiRqTKPyjqa2yXhkK
C/WqzC5APQPJCZvooKktgrVeE1dWvHYoVDCqB5HklNawvBvzBJnGioubePnvtV66
nzKlizv94PiVOr46XvIJiRYjuzxj536K3zoSup3RJS2tGOvfUGMKT6hmwdBAZ/E1
qCJmQWBh3e9DmCuIwX3bHlRFU3NLmd4u4VYDwUBzziLWi7dmgsqQo0wyc5ib7z8n
scXXgQJ/PxnzBAKdLL8emCoM046cD+qEqiZGfF5slrcoejJaxLhWpxx3Sezu6sKt
y1VgJIJjC5Mj8z8AOC4MXlQMsyxoBUqTr3lCCw7CcGYb+mUqnV3/LSzCHloEcTph
UD3ZxDlHev9mAnIIxx6xUsjFLbUCeUNfMiJp2T/spgkFAwFtG6NYAX6aPl6lP2R/
mG2i8Laj3q7yrsRwnj+UuA1NWBm5GJQil8PvnoztfJoYwyz5kfzrEZ31RAB2XiTw
jOylI+atZoiSPjlUW1kxhqfctTjCX7bdJIPLLqyS0FacVWg3oAks6izpqfha5vFv
7014NdYBrnOTtqcBCFeXsTKdUcQHhrgVToD2XwR8zbD+ojNVthsp2tGEdvAGBUEJ
XxpZDi2Z0rGF12guxrJkauG1tixAo31JG5YVbJApStXBN0uJD8w8uNaaTIhq0Yah
vPkGM5rjGHx0xBGcnxthdJ4yShNlH4/zs3Z4Yeyb7Ct+U8MFgC+GpRAmFvrbVrv0
a9gExlyIXs6UgFpvk13+7PHbBw2hxIMFiP/+OxzPSqGOzTA/VmT5dJkA2qbh9dGX
enbeUzjYPBoMIcxhLy5LZEHKXNuvjodPRQym/5FekKXRc5lcuPh+pHjIOzwBpJPx
QTgCyUQjUNLkDsNtp9BSBg8kXmvnvmhgmy1swGGbWe0b+gPBhZ8bYyZcpLy8RL+a
rnWd3rLM8726xIRhLaJvPDgH3GIEnSaMbkfNJOGyq98Sr0cPRDJaBIdH1+Z9yo11
3CQET+VpRxqbsPL2dHOpl1o6AEWg4rTSXMuVziVZq+sI9r5Z2yqFjplhKYb8hdd7
gfX1vHStTu2M3oobTZO1LSmAqz8CYQyKtxeInmlf8W5pseUxrqvxeJcvrwEQhGHR
KqRZvr3UK+xBhl0knTsb3YjBhPjX++0HsQt2/RL4gHDibOoTmEWOoveM+nhbme3R
wJu0WAT8loK+fOaQK3eUpazLGtsnGe1TANnVWvo/66Gcfz0RorLTaugh2i/5okOd
0Aeva44vZYsf7GgZfFsuSPoKFniOehluMD/MmyWvZFYDizl4AxoqtUPE7kJijWUw
9grkSkEkPMIoIbnBJQzzHKnn+waSWDct9KF+Gx8C/xsmCkGGm3Ft5OfSXx3slW38
Qz4Kfstx6+Lsb43S2iX3c/3BpPX0KjEEIdPfedrJbsTWGnlZJ5QaueFNHkzZeOuK
btq2+pCXuyzO7bmPFDO/4PxD+yhtVYA9bsXBoCWilBgmCXAiWPhQTfko9JRld1oK
kOrR29cPArYJNrTRARGX5z1fmI+drMb3JbGLKE/YVeSrtxzh5mRzxBgoCaF7/+ly
D7LBaIJVE5CPdwTx1m7zKNMr4WLsIcF9507bz2ZIKEOHNCKboJ5GV9+pxXwrde3a
bQmGjD8HzaHXmP6jC1MkGuxBSvSXVfCfjNM1zAgEP4RxrPDSQpzXR2wBv5JagQFh
aoxensy7CdQ7FP0s3Tjn2D5BDr9ELaPb+nLIa0Wr4shnhd80TRkbK+QHlf8eXTS5
kApg0Jk/g/ya0BgnEPxhTy8YD+1UMrLrDGQRn+XmzLIHm0EThmtFPQk3VOiIPSri
PB9J4IYGAgLIi5+T+eNUHoCrMlyqakJQR10zTkQWY4cw80WHsYKYHxarqUhZdCoz
SOBnWUOYtc90tMN9fehjA0Aw+08LiCLANa4B2bg4ktCKH/IV/LWGDhPu5cNyckb0
9tJp/8rCXhBXs7KJ2p4yDeSNEvUTROuUHionRNFnbgBFoTwPpnwTwQqklKHggI5I
wbwoLvPiyO+2dFJ8SPwLn/ryyzv5Rxvw/DbHM5K737oZkHLmQMel6UBXWcyFDWFN
TiPvZUqU+qhs/GY/c78Ub3EPss1EdHXPDJW6bf67kuLho0QimM0uVuNriAYcnPti
nxnSSl4ZO4lKwR4ZqaCyJ99DkB2UZEIYkNKQJS8BzLQb9geInXIOnVPg+jdA27GU
3q89m0Ea7y8wsu+4Rl+TZXbozUvSpv12z/yAe8CTMCcXeX+rzCzxJuHQ9aXMDvAp
Qv4de1TwH1l65GNbM8MWsGSZU/j/63MyzYK2FO9RosoEQ1fpOUu+OwHUGmpaNOys
RH3GQqTZaCzO0IxGwZIlexqw3sMyu3NBekxFXytNkFFb/gZAj06lcuGpnUER5BAX
52sotlcZGKynEtjuDKN8tV7HXVnkKNGiPmdaZLm00nCskXXEKJrn3HZ71hlZylT1
jjXIDWANpK+/J6wM3zuO2t0NCfnv2jmt73+lX8z7XE+AxaZvlCf/xtDEx9PEnUd5
0JpEKIjNzlUGPXXzqBVpSSmAEAw72cfD6UurOwOOck41yLvK7ReYu2oUrajtisM5
VK1IsWz3e6ksRTlHZpnlVzQy/TewZpGVCPSaqc/TCYb/oqGiBUyyI2/ootsI6Jrs
LkuVFx6X6vbvOyw/NgrjzcxadKNYWWGxFGuKRIDCTLxyJcoauqedwa6qvgtL6Jh/
SKVl+Bo4jIR9vNHVja9Y31lAYhj30iGtnAtMPLUFq3oho+pYhUwb5pzOaOj6f7MU
6KLQln+C/O49B5g7UL8h3DDR4IXnFJOuTaqyXljMB4ztnviulJLZlAN2TGxkB9Rq
acCc/ibGdG4iiZ4SnVeZUTIzawk+4Yz1QqUwFiaKughjgbeaBrYXbVD+iGGACi9i
4T2YU78jGZ8qhmRjL6DpnkTPt/Jec5pRdBsEN7DIYwDSLwhakaub/5V95lBZ/pNd
dfhyHG/KQbXWbb8Ml6WndVzDtiULcHEXU2i3NsPeZ1Fl5f94neW+grKiGV1/cnTC
R83HY66D+wblyZ7g8b15cc/7vfsUUzP9rRTxpV2YB+074VDSjXh9TklLEpbVw2ou
6DpLKtFbmK+EzcXdysnf2Dh31CAZJN69QjFYYYHTvoBdaQggS9gm2NnYWhpgEjdG
YoL2ScorGSOdTSB6xXM05gf7ZYsBtPW+z0AZ9AJzcFfJ62eJl4MaAxpXhz1ZgVzU
nNkHRSfiIeC9PXuMA968xmghSi0jAqZEN/v5toZxUlfzXKrBWjcRd8AjnIyBNHuA
mefwADvDhsJN8vwl9+0ohZKL/n3pDa2rz2IbeZofAjyVsbXLjDIW8Bl25eTJGv/h
mostEYH4DdqhdqXBpLeAztB2kiqTiKOmlEdxMYLI3J43KNg8XC5Eaj1oyX25tCZl
G6HHNakVDIIGvkTDObiwCaQ/Q5BDJgmCkeBOAozttS5bpR1O4MpJm6R7NUq7FMcB
xRK0Aa/viVjF+jv8gLsHm3dtmfvtrqIvpzf8GP86rqbZynds7N06/WomCp+3SQJm
I+ITS0P8oA+UZ9LENe9Aau5XR5w0VvTNXwdpKFrN5X8hu6jo4QuN8L0SYiwliXgA
2+MIlg1oHNpGY1TJWNibKAPLpcfk86MV4fMFppWMoNcSSU8KSQtgLeKR09t+3CO5
Qh3OJRqw/8QsWmReajRR61Xy9ZpfbZTiUvd50fkyHBVqkTBYVJaW3sXQoVH1sx3r
RESOeZWg/OSWNTTBGyxn6LeOKhB6a0O2DeGKN+DVOEQNMnngTYkRFPrpJXo/IXEY
dcoYSTKrW9JOJEI1mylKLWRirTzYX1HQ6SAofiy+rAIql5HQxzLQvVZGwoHJJr/g
eRjoa3Cujev/8SpZ9R4cgckPgOSS3ugVlTFt5h0FJyf6DJ3raVqK9R4QFD1pzEWs
dH2QKUa5hxj0cxPpYKZXYFS5abhdwW13UMQIf91fc28MllIrGEIgJLRoW0LwE7Or
LaAY/LpxMLdNECWnUTtnWfPyTmqB9A1AuD+PZ1u8ZiLgPGy+BbDNGD4S5PRbyCeH
hd0bsehSVxSt49J6EwcOm9qFCRH3sesiUnT1vCPXMpqGKlJm0dEdPfpGmkUOcar0
c3MnEY30NNkZFwRMsQ95XRnE/4EEyiWwaB0BYSBafeFdWjh1rEu5LVEmAO9r3+Y1
VqU8tvy24In0hJw5MgbJA5u89j2crR9LEVXnuRr7UWwNxQR7duw9i6RkA8cHOemC
IPDIf0s6eCl4SGSx+jzvT3xtk5BbRMZzQLMzT9xj+u6LvN4TR3Fm4lWSjDsM6SHe
Ta1wWQaS2pSKR2rJ3WytgYI23RW2vqKZ3HkBbmsSG8Tu0HpVZWMYBprkhoyLAByo
O64WGNRUL/PxchiZzVP96RwUu9Nf4JabNzrf7PLInOg06PMD1y9mbw9Rj1I+EkF4
lw68i/uFr1yw1kCGNVt07syQFSEhYsKinoaddE2L2jWTVIBdpjdgyqk+/TLqzI3Q
y7XGrJx/LKndyh4KhzA2Vk+d24NDCEJOXdDj8ZrlD+AR9gkF7pf5m8Z/wY2SgYdk
8SlgG+SNdwUuj1dmU7oV4tbvyoQUo/H8B3V+hT6wWVi4ofTVZe6B0GruKrHfQvev
wkzgagV5xBbHlf12C78xYqFNTOHG1fiS2ggZAqa0/qOc4umVE7w+Kofj0Z+708f7
5noNppVn3C8ImST6IN7J6VqeNSSRRi8dvoWtT3oOMrpqWqs9syGGEuJEi9Upil46
ljrbkS7nbHDA5b+B4MOlO2Zkmsq0TltAxM06nmiapkgKjLdpfb9xB2HwXgNwAJ6b
xU9g9NMLevYxUZYiycv1xWDFDW1s9hMBl31KCi26Gc46K5mVxPfE3BntVgxV0Y79
gY8a4SINIiHTbUABYNONdvr3CJJuclPv7QcVkqOUSJFL4yu26mYNb56XVczB633j
xPcVk+d3dT4h1/40rWLRha9naZoujK3thdiGQDn6CYiJTdMWPUp4q4I7j0LvWVrk
kYQWH8DCvyQv5Prn86782gZ7MVZeln0F8woLdE9aIJ74ucZ5BpaYJDRjgX9Y7iBZ
B2My6qTHF9QHCQMI6pQJ//u1nXr0W6wAL76ILdQ0XYDpcwgVh44pI6ZW68x8CjyR
8QDS6pc63I3mo1MDL7YDse/3KjsnsuEcwdWnykiPWiV6SDVSdz1ddMwMI7X2LPG1
e23E0IZhgRNrPWCntHvuNQCFIt0YpUxeP5xZBCnVibouKjtHQz7LSUKGTg06VauM
G2JxV45DO3F7BupxQMWZn9hYKemtrH35ok9YlaH+CLDXHj2EEBxXVTR6MZH5ic2X
SQ1ACXKw4nAUv0B0TFgfiIPOAuhlzwRIhdNJqoURQzPxufb12WbrTlHyKqtCGplH
vWdGm1+83A84s58ybsLAVMyAT/m2LCPdc5zCnlgwAnMm1Nm09o0X5+HA9PlEWtB+
iMyyc0wJD+pEOgSjWfEw6SpiDgnpJCPcYPbhHkZGXH7TuW7NrHKL4BLNWSmmJr9X
KrcKGj4bzdR+EN9daoUikjjHuGTm9yXJguQgRN/Qrg7LW4z/P/FF+Yl2kai/09Pt
cYw60zZcjZ/C7y9WzsgmDNgZs+3H8J8uI0KEa3vOego5CCUvcOIfbf4WopGT81M5
nNEny89h3BfVMa+AEPII8BHvUhdyBSK9mVwdi09Cu+he0xvsKcq7o300PHbnfvfG
y7g4vzh0diou/hVMRCp9UY7QVGo0CeqeYPexzWYPhtRJMPPBzuTeKeDzL8MpCb65
kV6Inpbgy/C6mr6Cwkp8eDx10UW4SDFSKOtaNlUe9muniXatwa3HB3srPOsUzR0w
BfjiswUAdQdGwwhih/o1BFgVmYw65dfA4QJjeM6TzGrt/8X2jL52sIOuZBFXHaLS
u7p8WFHw8KfhTDMOxcBniKuhF6MWoCTSamE9PH4B6+EA+/Spci+jat7+rqFt/iUl
j9i5/vDoHZbiVS3tBupqZCe1YMvL6tbfCUtKXGfypFDNo7uKcNP21HCTwUY+yjQt
Q8Y/+EsyZqzwWlLPl3wqb304aysPQ5s6QTZunQhm8dp0K224UhAvg7DJFIymK3QI
+7tO2RQ5CUVPZEvY1AZ0Z+2yGBZ82l/hNE3jn5RWWXhazYWDwhKxJ6kqYZmx9lCl
zJiz9AqpGVBK/XcIpVzuHSCkjG1xToRFpWEQHqwO5rjSpQ/HRDUvYLbJXCqHqOqK
W6EaHNZB4o/tJCIft2+zpud8k6hY3maORFVgvs0PGmu98/CqKWSepyKvLCctmF72
VaN4NoT7HMaBeP0FU5N8KyeQ1sCJG351mLZhBn6OvrUlGQmP5EayEORzU0GIbrro
JU7JJunYNk0IygRtP4cyKV+yo37WcuIdBnBrIzc1CLf3oPwa4NTqgV7pZDEOaWkb
eJVj4VHRqRtfN3axJY6/bC08R1FB/7f84PKSsHRdGdWZ3rE7NwZcxCS2Kxb7STiE
aodq4sg1xpvynuFMKYwwkvF3JO5h5JwIIYE3MHsC3SKq4sjo5JCcKlsRQVaRNMvd
2wO6S9FFm8ANYM8ZEXVjvFwMbm3nx8uF32G67k9RkpbnVDncjTAXoLDSSCXURoGl
ZkncmK+40GEW7Suhh5eiJNvfQ4ke6rDoMbPB6SezmC1AO01BoFMcCOrz691VCWC1
CLCbK0SVpybsZj0lTmdow+heDoBrSYnCXXMtd3sJr3IYtwZ+CpKaMmY3DuiCdodW
Rfm+x2+DmhCt0XFl8vgqI5qrm8fPr7VjFmHyY6HZxg10IeAVHA8QSuDezHYqW9dy
31WTEpLfQY3j1rjg+k8pY9EU301jO1I3gSPkYuVDv03lzaSfT3DU2JRU2bt1HPmz
RFCdnh6msDwAyxOQeH3pY32Psg/MbniHG+PFqZbrK98dWeXhiCEvjaxHdHJigt7L
udnXQdglIzgcAyWbPrUsL/cwVUfv5M52b3M0yB6rLd4vuCKclxFMY4DZVn7pevSY
Q+tDBSsOqYzlG0VyMBTCyltVEfTSspi0UjrtZ4Sjj5L2f4NngsrqW0OXLzWCIGe5
CznWu+4PYfhPxW85IQAIeEvdZsSPBOgPScsnYbwTPqR6Fn6+91G9ONfJZSPCJxBm
wN23Z7d2KWRchSgWFfyRvffmGyx2uh4Pja8uvbcjQqACehLk6q2sf6J0uL0iiRDs
Vk+1BVNhCtTyMLxV55m816A8qUJTtKbp2Vz9tL74wqWvGuAmbTiYH109uX3C+kXZ
/JMRSdesSXtNG2z5lLtadG2j6gswWUJiIqp7uc21stjPuC7ptJy4jHOrutawZi9P
p41z21nZ44oXMFCmG4VI26aYUn95/ZVZo7S3OOMVm/63zXwJebh/AyxfsD0wnYnB
Ej3GiJnN0PPCZP0SiA1Ep/TQQNuYZ6v6M0VKocvrdR/8c5qN6quJ2Xh0yGojlhlH
7yoYrU8skEakm0Bjp7eAtt3eKA956xoxPMppxlzs0kKBJK9XfLyTe6rsQHEVlO1+
tXsw68/39ziyOrBA6B9IbWCuyQHHLTNCSlGcEMi1dyuocqhg2VZ5DvT7rrQLSmhm
oFY8f9nKfeLCXK3wMbcOT1nSg/LDYzkKoAHhJMj5WzU1LUjdQ3hoKmNvohAaOFkG
2HimmakGWr32U0X++QPHVzxnMaBwysRg4vM0dqVPpKqX05JWbV6CY8r3ylQMGnS/
hz6dMn8Ho+o29YOBiNoSUqXuBtK9GSYdy81B5Js/mYwnI10WfEtuohnEVEDAhu7T
wojZtCTODJezdNHAaoSXG1Tp6c4mPILtuHy0ESBySEWWYplj6mZ2TFCW92iYz7eP
HfgwAAgymbN8GHQNg6bxvWc5yAaWwzjBjcfoMGcHTjITR02c+/e+abDfzffil1Nq
gYzb5UL+mfjMN/QrYjHqQHzhjtDl0eUny6xBgbGhJv9ldNJuj781Y67Fk+NeBsQi
kHWnIC1Y/qKHh9jDYml8AdLFJrxu5eKbHyqE+0d0rIKte3gJkwVLs6BOKseV/p11
icXPwJF4fCs1nAoJ4qGUUn3XvIHQEulHnZGgump34uUA6HVHMEnSnE4Inodrz9bp
a3paCFKV9cpJ3gc6AMRC355gPR9ZckEJEMXj9QksL6ZX5X9aJ9hl8EzngY/ypC1m
yzTwIIsYGcwG8Na7yHhQzGndJ6ZQA8mIYOH/wvtOCBKvNiUM7WdsY2tLvxBif2o1
Ds6hyrREMRnd1bJJeypNxJE18y+h72R87LYN/qWmF59KjPeDxgEOCvzyUBPUrz/l
bBvExJR4YEKiFIVruxSB9g33kTVgdsZOTd5YA/Bgxml2tc7334usom/didxXAqF9
H1e0/EGubIMZLwu15fhKX8kHRnYbJGBUt+htfDUgTCyodW3AWhG17UrPJDMEAAKD
5zJdegsmcCq1Vo0niV7lz39k09dDHOnfCY6A/LHv1Db7CZ+kfGqeH0j6anrEUuxD
NVnBWDYwAf/bS8CtFCR3tDlPhXKinlmiuWPwt+FUqgbe8yclNVVhm7D/ILkTLL4J
Uovd+THVQE20/OrGKI56q73B3BY122uw06uhLtE5FPxnQzPTks9vWld1i48dHR/9
NsB0LgWrLOTOjum6AvluL7E3pwDcKZRFdvYuNXKGALWTGr6oH39KsCxjUq+Wt7ZE
Wg3JsfiAIS428XVSxFH1CbR2oszNxwZy9qBoDKrpX/JOe+QiCcr5me8c95jbgUX4
jD8ZFu9gioLuURqQ1KccnhloPPTR6i4N42XFL81GM+fVaPk+NHJaBSaJErYG8soH
JguM3EYMoGv2Nax4p2sVL3oPpTlmML5L19BPUeS+rACJJQTLdlErx+EIVr48vlrO
qHRD3hGNpCu+xneH6fBw0ib138OTi7/cG6/eh2k6Mxu4kh8PafLbsr3Nhq7IiYmW
JIybmK/qGFF9Fi/6Nxwpi6ujxGx+prIPzsV2aMzJHzlu1RXWSjNfiw9zEAba/IK/
q47lf6xpB4BWf0PuYUzUpeh73Ofdwrjw3jjHBMxZUyf+lZKo1vJrpG7i/glOXrPt
1nKOc4A4AWfDLiR+DH8uKNneyXkL8xUo6X9K84kkIPL39h6iylad5rDU9AFwBcyO
TCdRD5CywuWMhtXkoaOCGTI5J00PYAaSPFhoTel+sWWG+1kEyXZbx4GQwG8dyMEa
VziPgDl2K4S09aUXECtZ47IrkzoFAQg0MbvhjIVoI4GeYS4WCLbz30Q37WjDzuxI
wJvHNABbRaSFYhErCMAzjuf1TCs3IXN2Jy/03509lptjl0lgLhP2weDKT0ubvzmc
qV0c2bSrVhaRRadIZBDwwicRY8oe5Bm6hRnOhaRP5VJXvAO7THi7TUjaWXUdGQ3V
aDV7pxy+iA9B4a8W6JbOuFRUgQq1aJBqPngdl3KHe3CBizARcT0dh/G8RRrJgyu8
NvsCrwCB+xwQkbuF+RFj+sWPuKnLImjilpIMQ+1rrnZHfAMVWlZqfseC4/wyREe4
bkQjWLEWdikXF0bMjvTT09KwzmWNn6zjyxuZ+FyAw08tEYDX6JNqQ7kmBV6GvjC1
0me4bFIbD7aTQ9v5uR7XI88YcmXEsSS38axJjMBur6b+HrIUGu1GEa4RT5hIn+M7
PZ7sKLPRzeNMpDOkvFEP1zphxKpwKqMi2hIpbSdJWDiyGc2VdGJaux1MbLCyb5Du
I2h00i+iUjJdyVtpPL5Rv0E+Uryxq8J8rChuEVNIWo76XvHne0p1dYZlCyBBzyRI
EcnsYAfkg5Cq1mYU8jw0kNK62DFHl/LMOJy9sSkNAZWPXf6DYWPPN4B1uCBCpkCD
Po05nMuwCiRQzh4vXzOjoRM6Qeyazt40qEMevwqE+WnWK9UAEtlQm9Dmf8qL529E
g52aotvCS4krNIqTFrSkglNSyTyZVva5IJA9A1rFo6zQzTx+Hlwj2oqVWHmTSQpn
QaDn+TuRpFBbnBw+gDSzDPRri4g4hsZa0Kf5zPMcQBmM9atvPQxl4ipYtb98P9jZ
SKNJalLAxMvBKb6KoM1ZTO2KFVul6jM9RUgAVEpIG1k/CHJRL3d9+8knyRdEzjXC
mLbLNtjAmcBx/H2pEUMIXToBKp3zJ5ugzfmD4KKIpaBA0otPyrhkq58Y2HHaC9r5
dYhq4osFcaNuzhBVuUkVxuCCCPJ94TBMLDCo05hmSCH7W8N8mkpS0DAQcHY+jQlZ
ZApFKRmJKdi9BGqNvTlcdv5qPGanGu7c2eH0imuM7Ox/hxC5nvr5/+0ptSeNhaPl
z790wuAgl9GjLOBCuPLn0x2fFkYFAxvDj4Uwffg1Rz1tySQEBpPYc/CvVfX300d+
6AMPwa9MKqIsUH4WWgA//PqKlFOQz8TS14oPQ/ZWMtyUgmpJ6kuqoxCnBAevK9FX
bUIt4mRWuSteGs8jBjbfM21FTULlUcVTgSl61rGC+iee8DJcXwCUZ53g4UZyqmYs
V/OcgfsD8S5cjKsY5nMeiBsvgHaMO4DTc8GY+ntk+FkOx2sv9pfvUahGIVThTKVk
sgYND7Ob67N85QHWobaCiosZM1Exnerlb4Txh6V0mV2LiDPEbW4bclIPptZSgEVT
n5C5tms8+9ir5yVxs5zYUW9gTdxfSeVm3Qk+rqMj0NXhf0QRQpyqEERVYDFccRmL
iaqF79TKG7NDCXDHv7p2exM0hob097B1bYhm4jcpvpFbxRB2iJJypRVXgx0nmmkd
ZWFXgIOUFZXJRVt7UQdDCHFAlMMAjIEQpLwCGlb6WcuAYwGG/gIPhZ2wb0keOhcl
zZUA1jcsFujtg7gWxUl4jws480G5NUOmOC2Ncr2PNQDRDOBLYw+ACWIRGzohDnY6
LpkhhBnugevYTEpUnjJ1Oz2ooWU/39YVOj0ha6FSiWjj904o9pB81h7nVny8njKd
dVJ2SfaRDgkw5ziP3nubXBSC0SOrT0WKBgCUGR1FoRyst/hKOsj1Cro7FJc7VQzO
cUqtA1MKQZg4TtsOeYncx7Vp6GaOShhl70ds6LupP55TTmql3jYuf4CSldD+KiQK
sCgAafL9XgnXROjMVJcMmWZaO+DSd+xrpqqYQcbpR/16qIupucGHTYwleq3kr1/7
wN046YSBqz3uQUFQLDTn2c90LCtao+NfSpF8cFms8xdvu3GNS/4SG6Q6jeJv0L7h
V2hPmu4hyzohS5JfA6OkGfsbxbcz89ty9kWTUaSHWLHjGt54b3BePRgHKIUyscQJ
b9jh0vxS7bSL/x7uXWfGUgGyGHiWe/qvn4UhmOJD+igHXuNmeYOl7YTZNEZEwFeK
p5hkHZ3U3OqYQjYuM/BKE65MolrYOD52OK6N7Rp3JakUT7/P+jtSg83T5YkCQbU+
MIRzjBgfVmWIkc0y39jE3FxvNCniIBKxhQxlML/kBtt15jDLd9z3XCOhp+1Oe5oi
LkyNrNRkG3/M48ucr2O2yZQC5YNjpjn+VOKbAgsaSCW5sZxBCPBbwLvIeBpZhxXC
f+AE/5aDyK7I+n3yp2+vCb5XDOa1sRnja4zHtwb/AAjNbFGFlsk4Mk8dA7wr1qo6
jGJsmCOHSYEOFAqkSMWerpka1CN9n1vNZEoCRX+1aU97doopLbbNb9KuI+gleQYA
sYPHlrpfkD25AA7jIckZtYQcQdPoXY1iDZNBWVD5zWbzQr5uF0XaFijF3IRwsYnc
QmCV4ZXAAAi2/64m9AgEbXzaNsv4ELnkAzeWz0XbDtKVXzEJVUc2wPIpjYWCnOyc
1KrJO+Z6rIkN7gUd7WLIWUvk0HbHUquHU6Tw8eeT4ZEH9VU6UVuf4SFjkUmSRbrd
+0dBH2/Gj3tAwU49gm5URVn9mBj2fxhw1un/2RgTkTsWthM7lAWUnPTDV+i6x9J3
KBVAAHQ2lnH97UD7hWGj1yAchAcWjlm8zolmpXT+rDKRWBJ2aa45CpGyjokcuF1r
+rK/R+mc5JFOc5NzAPQfM/Jar21pOZaIkYE89A9vNxKgUEiSLd76MPUb2EKM3Icb
uibwDEUcW0SOASlrTWwGBdbt/7JAPSoI+71G8yN2vwSw7RUGwPiCGOc/MyTFLdAO
z+f5d4QDAohrDSLNlEVvscJBBjLKqvVUxJVD9Jslj/ipL8SBN5WbvJHVEeDzGVYt
Oa7q8XmD89O/RRW9ENnw4nXMBoqBjUUehga8VKum2vtaugm1j2t3VTz/lNKsttb/
U9bDhny9N9m6R31BdkXTUpl6VUCtg/0nD/xvq4IeGXTWNXaUN9eqcU9Xn6lqHmgR
HApmdDnHpbxvfMAfUbkSknrdwa5n1DE59rdrZPejRSDDzdmvi9ajO0pDS6rOkVAu
N+8ueUSGZoMihbFsIZvRbNHqfYckU2iANtvuGzgW5ThAlFmhvcQ4/q5P4S8VUbGt
2XfOcVVvV+hXlG5ug6+/SQBABTeRKgsN5lmAB56ckfpJTWtJ36qaDCWMwSRtbh/J
NPYLb3TzX0cc8AiTelC7KWc4fNe2MuBxaB/h0eBCuoNEvXfEXNs7DgbLbyOPpJiK
UxBVpsvBAb7KRetoDkvGUKX2LOQl0DysZc8zjDdWk07JErvJA1/C9ySy6cIlaS0F
oef7vAcTX+bR4qX57GVRwpY0Xxrj+h6xU5NhJaIbctrhMv7qVdmhVClTJfxNP0WW
bbZ9YX6HqSwmOYawsDVDNXIU1AQnIlWDVLQTeOOyGc5YZOOsJpnz1gDJKOtuG9aC
RvEfV+pnrRdxqucDhXhkiHhi8GsT4B0XlJopN9T0IQZB9W4yJo3WdemlwzDgnfvn
RlmtGFDqn+4Gr6XV+gKuyYb6eXMnqnfYQq/+skhqHi9vSMdrpRLC1kD+p3DhGkcw
4NJkzXo2MlKS+Z9JInXEqwYkgBPNsD17ofoIr3HzYhEPsj0Sd9NFkg/hS8dcnYAa
n/lArdLw3Gg3rKy0W+9cVSKzKYpsBlS+RXTGaXjiAVowNbj7MD24EXDJRCyNSqUI
s/vZiJFjnoJU2oH4naAfGtO5KJWeLSSTCe9Q2f5dbZj45p3Ok5G0KJ7VcUVcMz63
+8PKli1eODTLmheeNQJLWK7BdkeAdoNk4jylwW5uS7sZJTyIMRYXW/uUZdsjPHFn
AgDPZ2bHxQ0BRABmreVaosBmrvqmFZKtnSQ+DwskemDBVc+2IQ67o47tTRz4nfUu
EonD76g0K/5H0e4JY4/9yqR+KWfAn3MjjZ3Hvv4nZys46Pe22QNTbUeJV0teRrwN
J6/erIu0EM4JArakLnu11L6BfIWkgpkZS/l+cEsH0N9U1uq/AZbP5YypkMvny+j3
2MNonIl43PjeRRQLnq4EfWP9B+D3HOAjB1WOgEfSvpWR/81+vxuUBnilw4HEVzgK
efDAfE7WlawDxr4CuSsj1qgT/+ADtZ2Mbe8NVcdnARZD9FGF6fHRiSZKUaP/n0t7
5sK64uLCodx9yJXqeRB0rq86zfdkaezIe2pF4R84AWe3lmDiqOQ9Yoa+gUsy8vt7
DSeUzr71cS7Ilk5roeVlRJ4O3WCy1CNQmfWjuqwxPhHwm6MWvTT3DTP0bvSSeLgx
M8oT2bHODCvS/+0Y9rTiBJJ8pwe/HEaZjHhsQv73nCDPfZC0GwnW2aZk8bHYwhTD
SYXM0mNyDmYOemMTa50NV3ntcq9YtY6s+KZLhC6CURsfiqbHjQC0FjbkQsQdGo1w
zKAZn1rP1RTvN5jR1J9CcF3t3C5qAeHtVXeXOCPI+NQzeqz6SD+eaPPnybv3W3CA
jdbizu0O25luKLKugkd0O14RqoXD2dA3o0n4y5B5bDlFrK9aHclBWTTP4mHTiHZP
X9PvUIr73hfTbvVa8geyUE4BKpyLjFF4mHch6rIhrrYuV428H6amHUCJ8qo1RMC3
brK4NpYdGb3kslp5VPemoYOASSM8f6dvllsreP+2GrVTQkl28tqpJiXCKw+1ej74
5RUND5X6GXH02HhVZ8D6RObaeFM26dfEXi/9UPCBmdrLO9aO1BAQPtcUj2eelA72
GBcLfespEkgZaqDv4mDxnBj8NCf52NDvkCuEdELNnkwRyhLHw5JlfIofaqyx9Nxj
isw4eYHJME4SMv8TJ5QS9OisfsqbM35SuJE78omuVMGTzplSvzFbmXVHgo5KPRzs
aI3Ys+y6s2uBx6QRb3+/Oj0velTX6j1IuEOCzIlN63ROZcq/9biyGJY6woLfOAHv
+qijtMgiAFfG7oCpenoJm2rfjcUadJb9C2zQcAHswYYAzbE9HXUx2Y/ua47ZA5x6
28Wzp6HbijQ59OHCOnYP6CeoHwbg55LxHoVzByY9qSe87Xk3wQOarDa625c2j6Wl
D3pecj/GhX8sGNb10zRXtUC/T4rGI3fe/VQHVzlxUp6Y6+aysP6OWmH+9U4xizXm
jaN94cTiUNQnbXlot64vDdfti7zJ1je9/DJx+l+XI67vteEf6dlzrz7PXWXLN6Ge
aygv5J2LUtMsnQlrusJ9Ybi8cuK5InoEsyhMH0E6Lt0dsMJnrITHNb+0WqAUw/zR
W0iAgFROieXhwt2LSso799NtzvK/61kiSIFyuAs02Zi/jFYKb8W7bQOJEH0AmW9T
7rhQeQXzn5k/7vaNqWcyBj4lvDRGem6vTaKskuQ5wr5LMloxebvqxhgsqOtkKjDH
xjvoifm1+TtAFronBCwL4vViEnF8S8KCzmOstcjtn7B1B6hFpYgCLiAruw2kp8Qc
kfGhY6m0m3e4XcxWcsV6Nk+iZuPnkvkLWFIVGwMQFiJwAqYGyJqZkjIahceLYNIz
byXtTp3MHwSwr/p2IW1jDD3ssqdu1kpWv75jGXu+tEmbudR+kr1XHAcg6HZ/wKSJ
LN5h7cNNtVyomfNR4vyVbC83kf/E3LtMblzHlIJM0LcfVQJjbsveZ7GMBFPxf6tu
nke/IhvlLeOk1uQs40ROeC0QJmoeLA4/RMzHfpVglLo+tTkx0uiC0DZTg2qzHKqp
UePGnBc8V34bnrPpboTOZV4uUEw1XLGv2mNescfyUWXWShIaJPFg9M+45u7OlzOc
OKnvkZv4ekI1gnDFnyQmzXR1TS5le6kA0vzAFR9yxHpPPRQ49Fct/s7BKw5Jk+m+
d7gQuPDbcaqhht7eYK9va5n9+PNrySNj0zEBxy0aoAfhRHDfBkYXLnm6k6SxIC2q
ZnM2a+ZGK+AfcIsTlTekm0kXNzN1ztocuRrY/bm6yNbapuEKAfGkmv+iOpJPAHjO
FbxRi0YKZXjY3Yd42oFFcyA86GEE5KVkL91shZmxauBHAL8sUJWBQdqOJqNOm1X4
VLUHLL503BdQCgXjSsMt908syy4tPW/IuATWt8+ytx3PHTNSdQdzXuwNZzE13Dk4
DnHGXvAUaEnLZOAsaK5MPGXVY0/wF0WD+0mH3Gsddu1l3J4RPe5owuzm9P8OLTH3
u+MPXUiwLwzCjVCRl0GYoJg2gVcEhKS9BkHWKzwbYsbY/ODrEPDP2bDtUDA52aey
OBmddeUCrMb9ktyIJ1fd0a/sVtiYkWllk9tm/rTIUde+nqVjYhzzqJbkBzvTUL/z
nK1/IQTCQDTn9+aI5bR95x/6UI52GvQSMmKGB8dOAwYBgVKfvzTJSvLuQF0qnNmM
bTbCHyZlAnm5C0bsiKHhfvRay+9j4sLa9B7Q0pGJJJO8ai/pSXprb6q8JlxP3W/6
HUBFkwNbu9yScgK9/zTKT8r+CEecQMJg92fr3AAA3hE400uV89cG6jc4vAF4j0SR
YKvZYI+xMfB8T9Ybzxpvvnl5MRXCsm72HrZPBZGbqD+rG8PBZj60z4+knr++nfgq
OYF5gHoSu/ecK1R4kDfW1nVG/55/dNlgUXfFP87dqzIsTNRpKRwImlMdj73NBtSm
lL7osD4/AtYYf5+VB7HqvJKZRpaKo3c0xuq3HP3WTT2lOsgRqBD24Jw51lRkoLoU
S0X/YAlOd2IOk+tgUbxCzSMpYBHVg/uulnf7gp1M4yKzf0I35BJdXEScJaRZH/3d
v4hk6BQ1q69lCfbbY4c7RkNnh4t3nLk7AeSLb0x19844SMbn4ZrSE+MrL6n7lHn2
91hGjnWZKIGQnuwafcN/Za1syIi+4BdG+45ObguC8QADqHuhKOHfciN8KsRDpyys
dYO16NTHUeqkDbCpz0jzhVdw3nxvyzUcWnA6nwmSmU9wQwPNuJeF7JXUoM/6FDWT
hfaS7RyFJGYc7JqTep0Bn3fGREP1olbCd6nwo29p5SsJ269b9R7w3hnpuXwUeEZJ
Pszkuxwgtkc3jw3Ha63EW0/ftdhZ00vd9BFckkW0dwlqy1T83NUcrIq2Rd6yxr6Q
2X/9hZ7cI17SEeLMSEXRMX877KHSeQzzGXOUDIAGsOSiqzR3Ugtxa8vcoAP8k4Ez
y9BNfMv4pt4wjDsHwMaOjPJmc6Su8AzDeOLWdEbqACuPOTj3Ryb2Wy2c73hwYdqM
UBMiAMo6/1CFELCHR2n2a9o7yRLVkQDp/kCi5onr5URXBm5QitrTjfEAAnL3Knmb
FO5ZgPyeCFA7kTlrROxzULlbdL+LlEvqY7gp9gP51dKmnaWmy+VkW1gOPtG0stCe
CkzWoGS5AvkOz3rV7/Q6SttDJSt+5cNYoewRTUyb0SgJZudxgkl+ThhG6GdE5KVb
o7OydtoBEF4lPK4pdcB3AcEDjhUE77+Taa0M4mtTaEmYOsvtBbnbx3ZLm7YzY4eX
KHrwFC5nxOnG17RJmtN+itH0Qtrj7s1bvSVE++oh487+DGjvbdn3qR2t/7pOCIqb
C2XFHammGVPBsWkyF2UBrHWXaB7r4xqhd0MBj/xGbFG8wJRjmUulGxHijqrGude3
TsPVJtuUgTiPL7CcpA/jzn9xNKOl6fE24fxEQtXRLOtA3/rYdhcVQvUrd3PZgTWc
n8BTc0HUDeQfUfkVEq6BT6SlQHwJqgLXcjInnncMaX8r6NsOZGsOCA0YirJIjocc
PAWy3ywUxoT1Uc+HzIxUBs/Ne9R16bTJEPOZMFo9wCk2ujzdxsvCz9b77dD0wuHg
mCg2oK8IDPCXfbkTXDvd1Juq1wet3MMjZNpKcmDTyGfY9swpE9PLTfpm9QAwi1TZ
rRgZ7w12kEvnscCaa8MIJxCX7ZtXelIol/9JJqYWPuzyPxXmCnNcGN3D0oBjtIKc
yqkTaDF/xamNrEyrJz5tNw7jHF2msVcNyiiAV7eMgIsYNbj2hT1T/iQzbf6Ue/DD
XjXn8Q151g2IVFBvPmFSi7NZZUS1H54DK/fBmthDsj0+SXY8jXZ4+wwcTIGv902B
ZJdqc9UXCl2c/6sV3yaD0YWp8BOzXV8ab8nBylXctyqAnJZzYjZXfYB4HO+CwWRA
nPnzO6+VbBK/MB+9j9J9JgL7mI9Iy4mZjRYpQEy/WUnsdAA0y03rOq9QHR05BJXh
cgLh/48YArMnD5sxFr++wyn02t1HDXaRzmt0cPEIPamdz/etCqNVSH4aAxujH722
ixeyKvow1DSgEf/DFtUNgpC5kEKG6YllUx17kCR7NbVK24yvUVcY8pppY17fa0ma
fVdbAlUmxmsYrQA+NkHWnPpCPv1j0icv8I1zlD05fnGSv+1WGqj2nnE5QGJ9oqRL
cDmAC0SHA9Yu/SuwQh9CBWkcuuYI+ktlgUF98hlrhvjJ/nV1EayUcm8xFLomu69H
Gu4tNF/p1OHql1/dIxNLzqDV1k0qbIEgiUMcnMgV+RgBt9vKHAt4aAI7hAytnfNs
QeF2TjhQ42kUSrYLKzQ8eFwZkadxJMHh3+qxE1F2fVx0g9g+hAvXFPreJOTTi7Fn
cS6jm9Sqz2zsRKQg2XgqoaBYsUZHebbxWnJbkpZpaVpdPm2bTWYXCU1Ub38CXO1U
/lt5PcgdfVDIrSlzT1GR+mx/EzVijXuIu5p2Ug8kGiBWAK04YirKLI3DRJecBNcT
iiPsgNvxx1hGNxGZWemovhvjOqxWmOwU4ptx/xFvAGuA6AhmIuhFHKW/THC2us0V
Ohmt7YuYHBcoSH7uVwDt+hpM+lLCcXGkU5EspFNhyJf5Jeg+UftSkALc3yjCXjR0
kickjkjgBUXeJBjgSUxU/rTKyRvmSxJcQCYGVGZK/SyexUN0K+YRc8LDPlkRjRqv
pCW/burnsykqvYfh9HVhEvUo0juTlJlc6noht4XMMxnT6ueMDQQjcefpscr5Boao
BQFt0VJDIwxWWBiImGFIoa9xCuwpSEfZA93x0+Ds5shS0j0Lg/w4Bl+wzxs/c0DW
raBrdhDo1wWsMpSC/WqdeFoWeQE9S0A1H8s75YpPMdiQGKH9j8ZFXEdPnlgtdKZL
aZb2hka6JiFtz/xDFEXKyfvOHqtj1rGkDO4ZWk8YUSL7TeL7OTVVYsdG/KECBrED
kXFDoV+tS6q5y3xH/9ltSNDCiwvZZw3/cvJLABeNpasWX4wFdYqfrTvLsehLicao
hEUcnSWP51IlQpywSJ5JPrLitkAqibExWNpr6GYEGmBvVf5Gy+vZSH8ZkD1RFYZr
njHQ1cg1yQWK5G94laZX285RJOfyk3uAfu4kNbg0K2Tpc+FGGFMtkKxj2LaNuSgP
IvI7KV1Eq4Uk/KsfUqEVKrrA/8kmJYfvkHlZcCU0Fv+hSSAXcWim+AgcuyevmTRT
18eqeEMcrst8Qjagu/VQWCCr7PJl0DIPiO6MEV9gAopMUBcijD6tikkUlPospFda
pnxFMyQBWOpUto7kKYTN3cvyBx4oMY7mBy+TPULDJi95wbg0SP88VDCKU8rscNTs
rjKk2OUrGSw6qtjl1OGKBm+osk9zu4hCYTvrtQsDbGszypN/kB6AIvQPc0DAmUUJ
5iFPjdJwilfYLxm685MJKbUtErNENxRIJaiowD4Zzt0eyccYhoS6V9kXxU5uC5pe
ZvjfrWdRqse1kN1ZT+TaWd6GEPzOvBrv4nwF9vagQock1QPo5T0PdvgmlUdnIgjD
G87JFI6MCHBZlMjSIf5dLYeaC7vcqU2BRtt44ueGzq4v1aV3iDwhChZMRYbyZPPb
8//YX8s1A3qQdTR3SIXMkUtVrT707poVhCNmKhVRcy9Fna9PgIXNOIFcDNmAITcW
gkMC8u6BB8OmWmBBSS16eHkAJVVQ0KFncH/wGtyrIZNKYzkfaU9lirnwKKuUx1UY
xzs6KuSJ4DkUElMN6uKIqq4uaYgitF1vdBsSfBy6XWBGKUuFHtrRo5JfKn/a0Xd8
ZZrFClohWj829SstuROMvMdA4PBEfqPznEzhyHgm41SVJ/z7bm9vyq0qtAYEivSS
yuAlckNqEq7ZgTCwX3coQMn22c8LQA6LFJDpXD8rAirujaalb4NbX8Bn7rlooHxQ
wFWubo8jYBvZW3e/KV6iVSwKjyUPiUBEHWtplz+STVQlyv+EFpxDvXR5NgNirSFt
745Qksm53BaIkBfo9Md7pxOVwmwiVgXxukKQPe9IbZHCb5liyqpk95KLa8A2YICK
374meX8uN5bCQwAcvJnWX+0DZJFksQ+gXzXgvt9GbgVrYQz8PwlXZ1wyHYD7cc+K
MjPLWltrkNmW3H6kXmzaTEefNmdNRts9dLoJrEz/EPtrUL3v0VMpEdsaoeeRxQc5
TqRlLQGLZjtGhO7hrnYvPtQ4rhuLEj8m/chQ0hsM3o6/4aolpMH8fOX1C9H6q1X+
tBScGxz4KBP//FaU6DkJiewZEwcJlqz0QOFTOljzd6cNcZwyzE/cXDRSIgvKyqMK
LwtgegFyLqlmmPS/7SIFM9x+bPbFE+ubhFxzyOtuXR7MTgWuxqbpDkGHvkdbH+AO
3J83xQ+L7LQfxMjwOJ9PEXAYWKT2o8FYvd6X7KPIsx++73Zo1T4b7QfJbuetQblU
eP4BfoSi9q7fMOsmvdtm5oNVkj/tuu/bkSHWZHW1XjfAAvHD6JnpsTJC0EnoxacQ
Zu2C22n7JX0UXMy8og+2yhR1bSWmPl2X54RyuodY0v+r2A+z9rIWmr/YmzaX7iMA
0DSsVriqazklVgSRgPov+xJ1bzyEaAgsh7r7krYvX0wlRQcSUVh6+kP4hn7/Yrb8
kNp6gGSWugDmLxeFsQjJT9dGe5JGdMlBh7R3Ics3eraTTbWcEEFYQMEy3YMViFzh
jZQUJGHDCi3osHXCVd9tmv8pVw0kCTUUjuQO+9/xjbOGEVllUQfF5zaIKlpN6ckg
8+w8JrOaA8lg0hwNuS3c52MkFG/bBoYhQMz+BMbGbEUIMQQntsjdSBFpcnxLJ9/h
D4lFFFUhccN5jX0Oou/i4NF9MwgNGQPsmJeES3Kq4luRtEmcwXLcJ4Ad8jSshKic
ex88P/dKQ+Cw2hvsYubJ/Mrxv2iXqBw0v+Gx735nsKK3mBn1NEjARCuA766BxJ+f
NqU0IUN01YTMfDMNQO8YEpllrXwnXbKROAnNq6F6o+1z2rU+/r6rIywFwKN9FqPo
S+hkFYqEYQ2qz5JNq+CKvkenk9vCK7ZhxEMBo5l4KLW99DXliJ4hovm58ZzqqTXX
c7bejou6an1cVat6C3n/7c7RkyAGRHph4sA/MHzFmkaXWkUWLj9X64zNuYKptBfT
Cg+92AaeZGlj5dm63hAHYVeoTtQbRcW74nbF/NSH6DRevqjZpFf/QsY6jPmgMzU2
GDjO9DrCxtvGqDKACC22CQAcWUtcxoGoMItrrFcZNW/RWgnHwo8ba0SeDKQ1iX5K
33PKvHtJ8G6SumIpRUhpg8A9Kl31N5vjf6XjNIvCi7uH2PpDOPh4invE8EYdSGFO
ZO9d23yB7CRBS2j6e/8pxSlE5M0ft2J6T5ND/qyEB9Vb/h88TdRQjoboQHz7jDEH
+9lRXjpmQv6wZpo8Qi7G9qdKB9c/sB5ePHBjBs4AHXgk0O/LjQ00nEjjgyUyox8f
AZkj/hSD4YWRvYHCauY+amFGXh1FUvPxcq1Dml5HDEcHNfgCVHLxn1ScYoIwIJu4
xprHwpIYEAR9uUOw3mzfv/AlXCQ1YzfPwg5v1D6yk2rRAV9SsyUh4QbYsaaHOcab
jrRCLdrYbKdrL09PQWx+FhdkEppYWrocWIYFwQSlB7ITlCdmAt6OqNCCCiDiNtY2
AV/KgrP7oSX+NALyvb11DYOhMCQceNO77cxV8SVAFSgHjPebDGsREY2t40TNvRSx
Cur7elurR8OUysmHURbWOEuG/eAqTthunw/e59ZPzDqltaFzeaTaIQAs5htpnvaC
tufakuxYTsYuUvtS7stNtmy8pOkRn3tyKCwk/mAirSx77wakWDxVMy3/RQWV5MJJ
CMNoF7PetPRcOAubT5AKrlAgY5K1i9Zbf28l22VFMVLK/PV2QCBgQWorY+97lQz7
fNzC/2P/RRO+Z6ul1QVfXJSTEiv4xOSdlxRKvA3+jnL52coOD78gdNPPb2z77oB6
Zu6LhLF0qkBFvIvQBuB9RUuMoXG2fpO1xiGpgwfpDKVJNwusmLxCD5s+lxBco1Lq
cSUIRq5qWzTChFYRu0m3JIgBk687kHn476Pzw3At9WWDLhwi23cJoNBalmWplFxb
YpR2pcCop0ogZCFP/KheIaXmEoy5hFofNemzwWQRyGKdlCrfoPN++bB1ZfFE9KqH
rwrnUg4FyAbTnY1gYTnTksFngc6OsDWFy14UE1Ozu99THlgxMVd+87u7f9WnFOMm
cCxkYNHOROPRHSyp/gZ1hpVPLzQUF3p+6oKP3ljdyjvORpFMMum1DtSA1NklhxYK
3iPLcYZPVDAxH8aWYwhWGZrXlReav+tYSQwcDRBiY6jpz+h4kJvXkpVTu5pI1kM+
2VcVXj5trOGhpkPJW9MB4ArRjWmHWdaWTe7gLywNsCKYAJB2tLSH8QwyNcCtcrLC
iomY8chmigKwQIfQGmnxgToawGd9p+I636vTW72FeMTS69o3ZkPrJ4esqezNPLOU
0X5w71KbeZO9cb3Wu5NCxxQTLyVGq+5V3zlbFuliGhJnLnzV5CwK982DQPFENmcv
6fQ1iMU15+8DTOgmQNg5AH1ZbZjtqsv48aRTRsC6+Vm1RB/CVZ6gTYlUGlT2aMxp
G9h6LnWkwRBB3WHdyE30wRrvezEKPmnC6gZ2VNVWaxD+bqCGea3uw4KnMgYaqTUZ
1WuQciNLU/QoLa2je4+/WnPGPyuDO0s2PjfsC08buZ7yktuIbP8pYVW9DepwJCm0
vemOF6eUJ7rNMRs2QpRBRCef5PmkxSjfsVg/NpduqA4K1wBHexfZjt75WDyAEnXN
d3KShrNUNuLsi1CI1WWKNO9PDH+0e6MM86t9jIDb3C/DVyrNFPE/zPdamjojoJxU
6Sh3Y5rY72RZRWdQSqFu7QOOz9J266xlXPb+HXSzdOUq96kmywlYRiBKr+Mwmrb7
IWLzPDf0GjfUb+8UWpWp1b+6ss6GXGDTlpE8e8yOAguLzNlcYGQnVOiz63NoIcfb
KirwabwS8JT2/AkpXMjPJFSw8iOuF6rfuR4CN5PVgB34KzLpZ8FQffuz6yS406cr
KgNDVVp4V+63HFBDDPUnn7AZ0el/IuBvkUexknVMfHriy0ahBjMG0J7eG1v6zfv9
i4+lYq1Sw8fxdIc7r6DA81EajZ+s+vJKpIyWHNJD1B7+nOlx8M/X+mJradwNoh3T
Jdw2h7nfeSpRwt+KCO18UDKgDzkcLkzXziWmY/zKEoQKagRFivOabHvn32ai/SH7
NFOdr8pczlZqW2uBqtCgeFNK4KFB7PlG6PxMdLJOcONUUKQTHXq7i2eN74wcjzv1
vrlKFw0DN2HKEXkDh34gWL5HJNBkiwFMtqhP5RAxqGyoyeaa2pOhDPLIGbABy2z1
gYawGiP5XmmYLoeecYfU/OX3kQXI157uflwKVFhGs+2Os3chOVFH32qqyDfJqrPW
OPi87uPDKGcdRz917mxsg9QzFqafheq13Zzy5N1tauvqxA9tdamGr8hhMRkfo6nj
VCnHuHcvlQ8Ie4idujEUPymXCQtkrv5h2oB/Y4uPFtzELzPEzIALr0mq9LFEE1eY
4qOhb5MZXkeU0bnv/wEqBN4Sg5+JljfvWUEgJFxD+CEjUZHtNFX364xaHG9ZI1Tx
60S/Fy7PilYY+CGOceRnDqG3KV2h7NMJUpcwuCfipXn3AyJ2987puVyXUargraeR
Kg5x32bpI2lgxpw65xD9mo3aFbClWrOGWdtYIkoKN2wmX4im/C8Cin/aJ7EZHRtf
QQS7GLctMXmChSD5vQoo9jkHpqSpZf2xNjPtsrRT77w9ntMC+JD4LH1kcJYw8zeT
keh94BoxULONWf5R2CnGGH7b9p4RXKnuvN8GFEeoymPs8EbI8nUNcn6pnjv9717o
UKyKjG83s1hoKjqqJ+Jvadx4CTA7kKfusOYInBBbqIH3TieljqIRpdG8z/UeJM8E
yGbUKOWjEZiV6Kak9FQScXTBYf9tLWUa4faIlMAlwmnG4hP5S/x17bYVepS4aot4
fVhCMnjYC3holpwyQSiqghkQksRT4aPQ36c92gAg8gRq3gGu1ZkHb74XHEEm6QXN
UJgM1p4Eg5j0mw24/d39IR1QSCq019aJSdY5VS+fY97KNKq3oF06O/YDtlND1b1d
4TtzWmzNNJo7grEaNRdyE3sTGF+QAC+8O9zEhxM2fF9jBh0NACxBggeNK/UwRx23
GT11TTjFuAAkPN0miPXGTDNCfUdKBDrAjP25sfSbq8tHhuuau/tgCP/olvs2nHv5
4Ka4NJErgO4XZtAv9eUOH4ki1yk+7AWcLZXEI/oznPLGIJ0Jb/7y9xAPEAOWUFOM
VSQoQVm/dZ2nuKG43S6Sx/hFWtQWrbPj5FFLfWA7LVDi0tkhfY4OL0VUBL9q3yaY
FdWigJPjkbGrMXKPMR3B9shYt0MSi8cq9vM6JJ+AnhQ8DeYVrCh8//Ni3KR5vJQW
+SW6mmrp+tr0FIavKqf+eJpCWsz+P0+G4/vYpbZCWnxNoMFYoweIG8JgpDCpTDJ8
SdVlJ2yEcdeLx221mFxzChrVUuGuWs0BRlUVogT6X8iuo+L5lN5ohEj7qGDkbfOj
C8XCY9eH/DyZIlkyksfWESfWI/Y71iZBOOP1JZ9e129x1mtZSsQFeSs/lplj6WF8
9w/OkS2E8R9soDgEl7t6FappyoaXD593HfQ7dvtzhYxz5vEfXv4azXkmX3fFGpXs
4o44AlbCB4tRvjn76DiR7tIhgvZAz1iGGTBLFUl/83zbEnT44YkD/G3GZZY+lZPh
0TVs0A92DFz5JUwpwbGxKuqraIISDQaiXvDD9gXjtl1f2h6XENUKu3qRiURdarla
p5RYXkPMNLB2tqi4raC5DC+UnKoviCmm7AQ9rrC27p+odUcDx5F8roPawH1JmAsv
G0qdsKArixRPUBpH5Mgxv/VophMKX9W/qK+DZC/RNSJ5Ai+9QYOPslyTA8XtESTZ
L+nHl5GaVEZe0jaPFiSY6gRW4OJJmxeI8VhJaLDmGs5iuFa/mQIEXj7aMySxUFIC
RveabwZqweVGpNSHBoW2KXiIuIPUJTfqUJkdIzgqw7RWr0p17QBLBaE09Ea7NNYN
wpXkVnpXRc599b4TZNw8VrhXsuy4VRsYOF7LYkefNlk/IhaXzUSosW5wLLRwLwBr
3ZxK2292CsWOPQkxVvVPGL/LSh/yJSpckzZjWecc57tyxvZIcfVkabLB0zPxlb+m
NDBYIqkIV0Pbxi5bwWb2piOPHILHlm1uCxDAuAGAlfNeysmy0cmICN5cZhgYTBd3
36GCIKhfh1DJ9zbiFavEIpcld5tamXtI6pIwj4kYi+Lownr+dHVDM4Rf0Q4AaClw
RASJsMJYv18IYlaSj9i7L3IfagooskjFhCS8oyQfuaVI4jk14RiNZpl4wUX/dbPn
evW9VBjSiz8Ec2ULgmtBDSATwzqHIqWls+JQUVyGfo6FSy8/x9Nvq1tmoXULE83k
80O3UrqXGPV6xVoFGKsHVyH5t1ZC3qXix8fj6nATEpVCcr65mjHX1PnrL18iRN/X
Bft2nOT9AeH6sYzBIvdKeyBwQT7wMd1OqKgc1QJPTnyVPv8Ad8PyMiLiOMae1wUY
Bmy05B0+8ghSAndYGZe65wDhVBOgtH4V2+PN2T/BgSTNDEAPWUwpCKWSj8kIC0Ny
FRhIRHv/uJ2xNhE5NpO/Fk7onMj8phJVDfVdHpS0zu+cC2Sc2i6NNOsj05UgE7ha
LKRlkPzlhacol7IVH445p6+4fD4uh2o4cNJXtzzIgPqrNyemxXn71m+9DCg8UJSZ
VJBraMvVgvDZv9UoIdMFNA9SzhDW6S+n/QITjW7o6NEArNmxVU+UsANLXhmY0XM3
z90t2hCzXBfm5cQXPixdipyDtoXVpHBFqP5ld6XOzn3JnHm9kk8OZrsoLpvz/PfL
9EZlf+WS5xaSApEuFH469047PC2ClnBil2me7486PpxGqa7D+v1DHyt5nb/E1fRl
XxQKIeiQd5IkKPhbaVz8wP/xz5/sco95jy8SqwYdcr4ho61twIouQmB1uqINmPPd
JAbYUTVHJjH4od1veDJxZKHiUBQk+ISzpQ6SVMk4QUoNc0AB7zWsD/p2pBX4mh3l
EZWacbeaDLI89nqi92K5X2Yn2TcMzbx040Mree6rMHgVBz78hipznPLOZ/eb2UhM
2iWxV3PrH38oq2hxGqKp97w0I5kyMTS3XIYx0olLkSTgJ83phOGnu2pcNuuJsiEj
WQQOsfsG7MWM21zWPRvsiK7XMUOIJNiN8zgM8ziYD+u2W1kFN1In5f0CCTwb6+Tg
x0ZHpB+p6veInnbukKAVLS7atp/D97dlzNRCVr/o4BXHKfesAIdA0GllGwwyM7aG
5hX6iF6m66UTav/2IGzaaHyAFXCRjbJDKybBYEtEYXUjNlk499l+ONQH0wsVSjTV
TNjEnjdkHGkRs6KmyKXKWvJl+1Q6wsXjwZMl6s+6lQmGOx/Ee+rIMxY0+9z98leC
G5N6Am9VKG3V4KWhZ02aBl4nUiExvxjs0UoDCKuyz5QMdDZ4Kn+BeLJdtuBa+Fbt
VPSm6t8S4Znta2egG3sl+wmpxuBt441lwcYSIuJx+Mnlzan3zyQyO+MOuJbBiFRH
zRuy3XTIGYhw4LJ6XLQEGIGAUwRAhTC6ToHr6ixOMjheRlsYAj4eDX69hihUpBfr
Ec+h0XlHfh39PBBuswDqAR+CrFG3IYJozEso4SEz4gXXjaQ8628+fLBR/fu1ttUD
nRMu+0IBEBctfKVKdW1dm1+MVAau8q2bYRFaMaBivPFhxPgIFufro9LSNe+smcmd
RhdPb9qD7ES8ULZAkCXkZoOlJt46akyUSxhkmu/0zDe1MuJjE9WO4Uku8izsCdqc
S9i9iWwoZxqhUcxo0K9r18AVDIZw/iN5cXTIyVBgcbkhkcxyllG2CBJMUT9yJ1Zl
4pcNSKKUj/CAu00kR6VgIqVr/J6iTTyg5zmeBOqT63DD2t8eY1JAhFUCETURax7x
D1oIcyhQJdhhFHq5MieK+Wzx7VjwZymEL7XbB4va8Sl07cX2MBT2RoQx3MxAvtGd
jlWQaa5c9AIJ9chPjFYU5HWpIoEnb7zc4IfRPT4qQJdF5LYvAHjo8stKm5AOpunH
e+PjXu5qaHfwdCGXdGZuE28dUffjMBP73XJLHIjFe/s9zZW7uz+cx3rNDqDgjOeh
OoukxJsCUF3sxYTgKm59HQZy+2vsRyPnt90rECFlkFKIpX/AG/Y5WSKzfJQzyISK
CjtBEt7KZ6DY+ZyIIfmXWil7JWaBCnSLHLr2cKHAVECh+vKRE73aTgqx4RRfJ5fU
lvmKplCm7oV8CCF7aFDwIwEv+SdRPyK9ToE/uNbziTyfDqQ+ssEdcEr65K4y7DGs
DuE9vDhY/bu+YxWJ6ggWQ6YmpqYjwLC4KbLo5xWrbykfsqNC/L6/WQsdot61VqDe
g2i3K1pUkaebuLgNFHpHj/D5txLQ9AO4RbpjY/O5hDVs1gqZJuLgN6IAS4tFbMYC
tArejikzcBmyfIwFn33HXmMstQPuxzuaLRsC7zz1HtkmmqIRjqtZUTfZvNRx6IS7
QP7dJR+z/URhuFnBAgMCwOqXvtkWH82zNM7CjCv/eFMon4riHZTquaJCkE+3h1Kn
4D9cgNmV1DQWEjSxqkgOTqnLJ25aVzjgEUg9QVtGmq/tWViG6jEvcqhKr79fkAQK
HGKl6R8JBO7Gs2BtbcQo5dCKY6OxH5mqvF6oOD39aBxu/nOlNkNIgnnJk8ouU9UL
4N5mMX6YQrYZZAdHCRHbRaisb7i3n4heDhyZj0FbGKWf56rA6hZ3N80S4gekhBxT
Tbxmpd5hAgr4eWVX656NeEzWnlw5LfIIbDystC4KSypbpd2dRl0rf46sby76SJZ2
3A5PBAt6iJvvwXAFel6HOmDn7ZpqPUULBG1dJE05OeUNFsxwslC29h7YSIcRx0+j
Ih43gkGTcCk+2ymBWDIfnovhyCCDtWAHUxFfCMX5ktia6ORMIE77QSPdLeZdQCtt
ZMtAIaHG2yoYx0P7B+roajPLS9WlhSQSsUAN+2+v02IT+QCVPv68J6t4HVyHI4yd
RBOtI0HlHnZOsmnKPENFeyCKOKY+flOQP8nP6r0cObsXngQ4K0euwu8Xdcln76Y8
+x5mq5tsFGkWK2ZfCLglfKKD2VuvjZ0OMh9efDvc73Hs0WX3o10yt9ix9U2WRZ5F
PiFjcsrtSOXlj6HEf6mJF22pCNAtAdx4HYn7sMoveTXu6qPBYLomZRY5drqMwR5n
yYh/c2+/QQto4SKtYeW+yshibpz3hVXDJFIcmXTGhGJtLDieL+RWPT95O/CM+6de
M062sj8c8kMBOKhRlmNxa6l3LLdWqGTVZ4AWgGERpWzh21K0quIgKVttMKa7uv2k
lkRZ/ZWJqBrtFSFaaK7HH3pp0LChSEGaFgeeWCE9xbOtl946+GxtNufKcqKqMNU5
zks/sERlsR79kpVqdqh+wbEu1nUPvX+CcFxLFiMtxxh9jtMx2ru71uTP8HbZa06H
lnFVjLHAhUYIyZxN9PaqR01sMSJ4DsPLkErpG3VNCrQt/JAGdHmejTWgaemenDGG
02Cu/eGFCnKFtrsfN3DafoejKJJDeJcCcYmLwHI9UvZE9xFHf805/fg0xH8/cPeZ
J1BHUBLwZk+xjyHIlxcLgK6GcLfY5jtKQ0CVT5swXQNCHWAPdahGFSbvD9Z0cn+P
/aV95FtNyuCjlILzC1e4xDx63V3r1BMa28qv+dcZdKbXXPO9r3NTTSGIN566+cDi
81Nikm9WFR8vZ1TK8QdfEM/u5AHETLHf7EZMZu9DOn+yEXnm4P2p9UDPnO75mq52
kAHtrtcfDVx+04KAgBxPF92wqgLQqFoVWmWuhIsdieIFnhzZ0xPDxDE8lDNG23kv
qAZx7VWg5pI2dVMGy64Bz/SW2RXA+q5XrCU5c/fYfc7YNw3cw4jHjvIuMfX63rpv
uJpuoPeJJBl53NEvXpLFul6hBpWGhKXUZBvBqQeWDuVQU5iLDH7Yq125UzxXuftX
6W3AGKRFycIuqMk/L1PS40mwPncVlUy0RZ3Qp13zy42TM86NqKtQK59zFnyQofKS
NGXOtFwRhVyv2DbP/hlBeLkLWQkL6r165JX5ZcHEEiOuuwXqpdh7cRQcnU44OrWd
UZhOI9/PXWx2FmBxxYF+cCe5UX8KfA06xDjmh11rhUeiKRQml6v70PPcg2pV+DeN
j+HJslFsnnHIHCPVyHb/f04+iU4/IX43XWV4UPc25aGWTtnIyE/1gSZHEJJRiL60
7yhi1Sd4DyMB/DAD1/dQrnd/q/rRdnOUL8uwDe4DCoZYjnW3cOTyqeim7zxs25m9
Ql+34jHhNeTfbmuwnwyS/1TT11dASoQq0VPy9htUoJPILLWzpnw4uBCK2OgEhGrs
J+Pf+4+Iw8ef5C0pN34U+fjT0FXzY7FEtfm6ooTQtRjGvI2UuiJZKRN+BBmVq8Vt
+hfMi/XKiUILwUm+F1dlqK6zjyheSecnj2o1v8sRKh1RkAk/Mk3dZDRdZwKcgVSf
tCzn/o9vYtCrU9jvlFndcL+a0fG58oqKkebWu6PmCk+7sKTOstDRSvSYD9Q0tHLO
rp/9w2IdUvRfRQYJpw/MZSnZ7ABIGJIq+4ULXrFQKbrx5HVyHMIII751MzEhVnfo
EkBE/PY14g95hvx7s696QchddFJmNAen7uWAbfD7nUyQdaXdMuaNS5wJHQZ28wZs
cXGdV0PGgRkmfsd5wzeH4512kxJBf6UQz7CUtRIu878QG/r4NW40ukp/W+2zIueI
eWvLYgEYYEOoo4Xteq7xAZt870Sd7xKVowq/Er+RoX5DEksN3xzHK+cr1oUvfiC2
/M6G00GwrFyTwYZEr7uQiHn26bnRu8JWNX833FubaSesYhNSiqqIUMnhqAMH17Xc
WoZeQ/TdKDAsdpPhiKH9ut0wTFQ0jZTGhTSfEZa3k8m2cO/TF55+tzF350yVz8ml
WxurAfsjMh+aERyzq1AhGeoRH5rrH7muD7ARzeaWds8b88ArPw2zhVIP0g16yptk
9TWCLkW3WYYp0vq8TqkQi5AOIci397gc6tqZG348aZ3aStdtMsRX6f6R5Akla1LA
gqptBNxIS1VFu85mniURMJigcBX/NUgd0VPgfPFT9a1Jxb/0aaFniPetXdlSKQ5v
uNUFPJfiFgx3LYCkVjRRkGo4qGwoMpd96E8/amyFhQjPOLq4V7ttrG23RHK1o52C
tms7Cuf9GMln+kRtXMu13XUji5WQOxX4aOTbUCOFQvpV+s21tSlR04ndFnqNb/62
HYek6BaHXHbgETfzBmSf5c4Wy4ne+zj1GXqcK05dbBVug9FNrCthRWemYiDMUiPF
BloiB2FQz9l5dm620iMgP7CQ5IMPg3YtOsgy1umeTlp5PwcEjq6SgwwSMR45uvLi
975wh5HeYpikpXOmEobKcETzyBsQ2yAXShxpEFkjpofTNAhzTO1F1hY67G8idmOV
baLjs4mz7szwQ763NATpVic5p1JzInCh9dZarUNQ6rOl6DlqozBLaXZqAf+xVxpj
ZgjC7fr2CnVkoVmFljXgtE2Y1FX4NkxKrP847mAD2Ml8MnZWUDW26VwpO+vRBYR8
laPxo41wEqb7WGr1lUxBLIV8Ka0I1VZvvB4cxIZNSXhY2ALxwI9J88F5fUP8AtXx
CRGvSFa1YbU+9nSrO7JxEqxoDDtu6MfrOtnsK5uShtfb8o4ECpU/R6Z4cKqPXBxs
/D4kOlV02MFK/MoCgl0MQLPIhIf2Feejehfzj3gOzDv+Wso6U0oLe5x+sToXrZoI
rSYIVWub7Ki4OsbOKDbzXMEUurOtc591ZtW1x18xoO/m2+w1W4OqeqrFfat4uiRw
OMNWE4THYUCqDb1iNYEBulFpUXrAjUjXK/VlSdsgLtmTFykvSbTYw/jWhaVzx7ZA
qtQJlkMMaKSGhM8x3kKUYR8lO1UIEEk6C5wxRNkw4tzMhBsotYJBnMeJfbUZM3J7
r+lkdlHqUWH3O/wmZZa1KDfLGlGIUqt1GYK6Gl5LzD4++KBAoYRMnT0aXMVkpsjo
Lg9bzvrK+pgvqoB/ie+j87vLr14L6/EF9G5VByCBPbD1Of2wLW3pAzGHfDR3rWsQ
/Xyq//3rjQiPfRq4tOHZmfMjwtN7KsFFEll13TjBtdS302sUrS7usdFsA30wgoFg
6/igmCLEWZ8JDG8fooEMmfDOICHAJI3YKQO5FmlXRqccSlEEQEzxX8VGbMM1t5j1
bxkJSnBEYyQqtJMu4VwI7t4IoK0FpmACq7ep8wPI9A6wjT+MXHzMaQU6QESV/jmg
ZFNB5W5EzUNDHJLzSEaLjYAmBgpD8XyMvNLBiMcQ0I4/YyzKH6lsiZV/F1ExJ+BJ
wVEMdYo1CLaBFY/LQR7tqT11onmnTZ1QM4oKbWxRheeeZ6PipLlcocAJwneicgRu
1pcwYj1pq9hmc5ejVrL8QiNoTgMJ7UtCKbQpSl9AeR2ZoIhpVodg1Y8fb5Sdpok4
fTD/js5jvXZGIBPItgN7IU+GGoqg2Okmc+dfP7btVrV1KZ/rco/AD8mRbOekmpDE
ehTS3Jbyqjxy8TmvLuY9x6n0k0hHfFUW7k4rOQy7GdTptyDG0kpqu+onj0gfSlFM
OotJh9uscULS3n9Q4uYAxP/s5iL/KL5JLMCXnFADHM8TMrMLOS5IUwNzIfrPoN+r
Grs59vSOGLhjf4WbwnH4FJhzwBFPOMysuxO5I/z4c9mLyxUeh24XLYPcKg7PN52O
TxjYLf1qOJ+OdRnwt4c58kQ+cMzGJdoMGwu1xgE1G9abH/XnxmwZSArcRU5pWNcz
3vSWn6HzxlTmdx2Gp2BW+GLIRSfleHoeuSoEjwtSrPk7FjmO5c2ZTO+byTVmjtI4
xbNEREdydZxwonCWXQU2ZSqtz2/nkQvQIp6r0wlW5Ko/ohS7T88urKEF1eegU0u1
2DYC+TXqpclE9zWqQthA8fVxTxNQQE24I8pMj67GMaY2riYHXwC5OeRj7rP6RHhW
qjexqQd8s7AKAHxPYv88qWwGgwV4MEH5sKZpPfFPQYbcGcalqSsLHUrXrHe33Ppc
ws/oh2Yr7QUdq2vn5bhQxPr0otj6HEeoxaAZ3KCI4qqu7fYz/dy2tMjZuF76k0Df
Sf+7ox7GD7NlDmn7aoBKn1PJ9Ccmqb9bGGn3HzHISBaI/ZtBrv12E0/SXSCci82o
HyswS9Dyct2tQhIu2A6w3i9g7WsZGZ7pUMPAYCE2UjzQQ67p+27YWkH3ZopuV3L1
E1rGZvANL8L8Qagn5gNg1bcm2i1PVFw38Zu7Il+nxgYT9S4D7TZvyX1SOOWNLi/O
B3pZbgWpEM8a+1aiqjyshnbEDPsp3kthRYrJE9z4BYYKXueSI3U87OoofpLybQm4
2OQgGW+jxFZGjtzBinwUoI8GOCL/0D9HmlmaDt+oO+raJJX871Hi2nJmiIy31q8w
53jpV9FHyWCG9LGuXGjNGrePHCrgtXDnuWqU+fS+14so3HMkYpAQw5NEjnDE4to2
BKFHmgPpQcb2T7FOQ0M2Hau3+ic8Djp9sXTpaXBeH+xrJ+mgL+SMBFh4RSnKI9p+
9Pe8zY93iepKQaqOj6AW0KbTmn+2YrShoJznrAwHl4yqhOfUGufPSagl9SEUAm8t
R9cOuvVu49GEY98qtHpRfaOfKUwChiION3rAmPNoSlk9avqB/wlNe8Cy/2+LehMt
vh3y/vmDi9makEP5lqLfyZxa4z8M5ipxqFh9pN80wB4nvPViMVVPVRbhEeAPDrNv
mCkZAgkRW2TwAGTs3vb0GcWKx7C4uVN6mHCjgC33X8yNIz5LriWYeoYgmhv2KQsb
XKGBf1FK5nxPk6FwCW6OeTLWQAtXz6Gm9BTo6oEj//QPnlkwipw6CIkE4qJdFiNT
Ntbl3Eqw/1zZidfkmJAokVTcXVdY1sGQlDyLYn4m8LUbevYsTgIQjz8HkppObBC3
877Nvth3s1fofqQ4yC06ROf3s2wVwCtaeHoq+gCmdbAAxkRLzpLiqBkTiqZuMSQz
Ax6e/pnQrqYFfloi9hDhxjgZ/t9+zF3M0RrW4ReqidxI7eHa+jwR43WxG/OJNVuX
0bMi+4GKyjZWAEU8smV+1H9lFyxnBlXy8dymSka6JZ8/jOxvAHhJg0O7Bt0XMRIH
ETeAX+vwWVZr9zWftiH9944k6P+4NLJarTIxRazAKW0r1V4NG8slryOUXCqBYPpC
5IxxpA1L1HB2rYyLYRTBgYukWXeEbfbcV931TPT5yhMcP2gawls4kR1avWFejXit
FqlX0mVsv90HJV9oG4cX7z/fBg8SiXs53dxRwOSPchk/NR4zUpFFw4baQpkVj3PX
yx9EQ2gd0aBJlpOdXu8KFXVd02TIWMqrMsGhIdJcWgeGeJF68XrIPuEP6bgSMzJ8
3hKtE8Al5qLhl0/e0o+HH3U8T2XFg7FNDB/+23rAsr/SXshsnv9LJSWDllDJtW++
4gX+T2ZZ3BGFNRF/4SSBCRl8SumFlKUQ2XDL0HTDhGY7l/5tSPS4sUy/JWq6mCet
KS5umCXATOXoK7sqpz15sGmBhJDqdpoKdDQZLmepe2HtDaGwXhHgUyYGPhVpASSX
c+PJwpsYP4Sb38tONI534yiXIQI8q9LkMbII+rjPQTNbaEho4RKZrnQL4xyFZAMz
TjkYiDf26yJVyOLxdooTpBhU09D4Gv+2zNPsod6TzUcYp04kzcgZcPKurBQFS+kS
eg/uKIbu2NyWRpnR5RPdX5J3XO1cEMIB6vKKz2VosqDF6x1Qi5RLPdmdgEZ1lSXx
lTCPqBXjP2n5g1UQsa0sq4jBQXc66NdFpSTaRLhV0Um/FQebDC16ZCBdBJFwklz+
J5Dk87QtvwlBuD/VosNCJzFU5Dk/7Os5wFHf+e2DDZpUPRJO2Vc5sMeo35FBpLhw
wchv/BOlso2mLg9ChLRV6TNe3KalLySSbI1/DQ5+MR7l2TWk1Y56nHCPHx0gIB6X
zPdrFR58YGQ8FeB21P4oOGfFYziNMUSJa3dpyA5NWW4M6qtiveqISlAS04hErcYr
t9C7h2kll0VoQ9uM+2WTHOxtyCylpcF8gGKAlqWOdfPxw36jDtXruyb0LIg25mvf
N4rMMvs6zgMSSKH2osGcM614S4ksAwVbjuv8+h6xmUET/TkKLH8IgC1H84y8I/3l
+6cfLxgCKH0evh3LdsPiJmUgb4gzrQG1ggwHPQz9IYcBunPqCTAFMYL78v0jQBV4
+xobDsPqZLyzDz+cOiHM53haEQyQ2HknL1GllDs+0le2j4wsLYwsHrJfGsl75Cb6
tQed6fFqFqLe6194rG2EhYA1yXj1Xlnnj3XCiL8TtR92S2Ranm91N6SJGNsZsfsa
jnT20s3xAE9m28SFl95F3fiwh2JTRf2sSc7FfkeYWFRd/p/0LQGxvPnYbLec2Rq+
wXcb5LheHl0a3KgXoHK9vKfdCS9jlVttZtaE1VnqxmfVUxxtRf18EmGkV6hzSXiE
4SKMNkfPLBPLrC7JXnFG/UQ9U59+CZXanxHa+bSb7tOYAJ0urcLUcbkWE4viUl+1
ccDE0KzM3U8hdUcLlinvhE3SxqlNWBXzkoxb7DQSv72jNf7oCuR61pFhnoVhIYSG
C4VCqPNU0J7OPN1qgc4CyDyIRKIpvSRsxDsA4vvzcwuBJTZrjYG3St6cBwxsxeNc
1Cxy8ZvnFTzSaAGX8yPv+4yrVdwzXQgUfivf8h5+/PnrjFcANp1va/uc0AfZyjRi
yr7h/NPIROgJRacGefhc2snJhJkhvMNdKuKyX5sMneay8RaMHRJLmCZE6q8JSowe
VZHpMQuIIM0ajw++++3NIPKcewi/DwVMK5nr6IAtQbOC5Z0X7Da2B4LIobb+9Q9+
AAgWF+pZ5XKKVwkiFVZAog9LcTpomYahox315xEUI38XjTGkvu8yUm6yU1ElB/jb
a1uuK7lJxovrSc9drXOvd5tk36Xvh5SUQMm4fWiuwV3JALsqYWv8905xRfQSoUP8
RDZqgWfrufo7e3Sjp2U/AXv3YkMTRDEYog7/xVze1FBlzKgXaafA+JnLY6OoXpfe
CUel6tv3+ddLs7FX6/sltHjKXPMbgprkjHLeIAJ+KpA6MZpD9cA/Goz+SjQa42FD
2N3zLj1ewPLRLHPdR0KcDXrqsf0BDt54Hk5SdbkZuIHs73sNws8/SPpcd2fgYSU0
HVOloQSGkchIEWH5S3HfkdzK+Jei+AEiQ6gYQWu0PJpk73+jzgQ60AFZPCISCX9L
dfnzQYk7Uki4AIRd5b45OxuramFqWlPOKzO1l+YC6wA6oEgu4u3ba/aRylRDk+pD
PVfQrbH0TVzNIqX+YxbwmsuOmpgyoPUnrtEMMnJI5hS3PCTpjKIb8MC4qKpTIKoJ
qtk8lGihnWeTDox4omb+tNPpEeeSdJN61M/PKmz8q40rWGRcvUSeCHPWmWBcccYd
L2mEkGX4ifx6VjWIJNZKq2oX6gj1O8QkI/j/fbS4BCvjVBtJot5Za3SesHYPQob1
jQiCncCYyN7NKyPra61gRRKCErJFNudqYNXL0cfgnGc2o63TSXA8gyHHr36TFjOF
KRycxSkMq8S8C3vaxXT4Z+ECZhvcbswMXtq/BrQR3RrJdSl9s5ZQGpN1La7bKnk3
9uu3lG2gZWZdPGl+YAfRReSvZwxIhtibqmYKgmjY3q5rMpn/QHSN5vTq0pTtQZfs
8dJZQXTMmg5uIQTgzyuEQ05SI/hmToDmdViJVxIKFWwSMws5egPVlxqn2yjcljdS
R30x78VKOqbkvDSO59s+hWqov2vplehhVq90L7imWQgF8SaIUqjKBFhs9BMA/mXM
BvP4nPIQpYZkZU2ah/CvNGiiOiUzYf3fWIBL5BpkWfVSH1PYzN8BQhBzqHPusFKb
EWnq7HI2UqMxHPFYfGO8FkOwUnA3jIjKgrO+vBUCr9GjmAoD7pd/A/jAh8xB788z
4VkL37EvEuuPM8M0WUYur0VUw11Gi5c/4vgOlprIGk/7LnLnJoY/kSXk0ntgfeJJ
N128F4euGxPO4e9CTLpHWQkNooD92n0c1lOziiPuHT/NbgYjdFd+tLIK49yChvj2
JrLKjo19cHli7jwTtP0qSJ7WWby5XPP5UBvl+LIJV7HM21tGQXTSX1L5teq1vgo/
+SloznuV30aSbTYE2+cVs7+T9AiVfOhuzbcTIhjkjY+2DdvK8X9gz0JwsuIz6CRq
zCgwRn7U/TLqy54z1wMDATiM/Uj4sOdKZRBsIZZFL7VZwuWDvBtixuDU5NxUn0yg
NjkEDuXRRiDzKcGzuv51tOJK9zzw8XQTQgPgFH/yh7Smwl9xsNBhrVfCtLibVq1i
4OIoKmi2Xox2bVE5IA/Q/ol1keGXnzz52voKLUPHrFZQDA5L43rNj2LTZEWdMTv3
ObnONuhNRfI0hktssFYnUw+XXVnUqX6mB0qdd6bmabi3v2kHsHpCt9STWpBSSZWa
aL5Ez4/EELq0OG80MDXC//I0zvTCSaYYkE9DOzOmZCIlwsmfYkcVlRQrpcsz3DiM
Z5cZ+ceWkwQ88CNLdJdwH3PdLziHyyJ73K27hQDkC0yyd978EQCRxRUyZRKCSwlQ
RsH7FJBwWZaqny9LDAramWCy3bA/IzkxobAleR97ta/lJBm7xwUf38gGIeD9GULM
O6lupKYT/+P//ppttwkN1fcS+bc7MINhn9z5t8JxxBIzkJnDYKIoxNVwSSz4nBKI
l3ZJyUvZ0cOOi2og82rQH64MaZ+xKlF/qvU7SawT0TE5iGWjn8L0hEPEtFhA/t4q
FGAnm048Gr0WsKAzHfuj4z3DJaKGqK/aqkR9iRDRTnDGu+Uy3JYLOajlveDDkKW+
kfmn58d5COy2ihIxrKV1zeu9g9aULRp/pYARCj61jJnwSIUV1gxP7/rtj7Oa7FS1
udzjHwc0B526ke3ii6mFR4AxiKfnhitsJzbZKcuvJotMeISTgXDet4CxhnlVstcP
O9xlcdYP+XxwSHb/w/m0mZ20ix+AIdb96wq1hQKhH8BC2CH+U1Yea2hHjYokpyUP
l2pjWduQv+3d8VoVsxErlYzzrswhx2OeNGKb3B4qYsbR/1tTKo4qjaZWiheqb7sK
YP1X4rBt3dYg+0qnfb87JjkYc7HV8AmXHY0HZlUrpebqq+9Idy62iN+772dzQJj5
dog9FhTBSHkXtrT61F4wRMq42MNDoDNs7pxaThOM/Qa4hvQVRDUVd/+KfybxeF8h
9t9R8Q5gL9yIb84MAIbTmyvM2yva2NPNC6BzQ/vlCszNDSiP9snnBw/jxvXK6hQh
nXHuM4Bl0mQ3leE1Avj2jNTn/hr5yfElBlXDx4WBox9kxSFQvyfsNbGy3gmvgcfX
YuFbO8KOuO5ZcQLK/Zz3DQDbJo0lni1tHoK6bandWoC30nASd5MzM8pem+qR3nWr
SmrurxOiCEOJMFTg/VmbCLOMg7LYS1d+5u8F6eX7FR6l1Iwxaes2Z+kNw/Q0M5Ry
hCk0K+Pd+BN+SWGuW88knBhorMgQxHbbfsEOFA1w9EE2YwDAu3J7Babr/HuDZ3xF
9MZo+6x2NHl5bYbNZN0FgeDdpwh25bwyggt7KWVo+iv3WgkjAvyp3AfOq4CDJJfc
wtiyH0C76GrgNWkzxhP7mdiNBx2k/Nh4IVFHoSNrQqsQoHmOxmBgLPFTi5h1rhhK
FwdKf1zpbMkCFsOQ7Culh93N3e6C25Vvfn6SKREKifMpPGEwDUB987F2fkrGvska
jKQpoVDQ6MhKodVyiSPaN7WSeYRsasr76Eahdr+dz8G3OK2sVcVZR8qz2b6P2olG
yRivC6A9LCsI+2cz/a7/xwdync2y8G8ziFPurD15Rqzlwlvr6bZTaBFNJr2e4Eyh
CeosUAkILbaGjY5TCSWaKZBrssHhLeVndHkg0M7txdC8xjjq1mbDJhv3mTxd/fvj
INf3eM+H1cLFAK78iHq+NtLg4FGVFPh0mOELTYxk6KeV2ih34IgGPvrC6iSsGprU
RKELl4OpWoppXvfV9x6oEPFtTDnrSJHzpOJqmeeWxIq+q0bEY41RGhFbqYgiBkht
f0Jzk2aicdfFD4Mpdg5fw4abmLljb+mibz+YpdSEUj50VW0fy+vmDjvVUKCZd8aR
lGIHaSovBYNNDjiI4xvcV1AjCvnxTHhYeLyoDtDKAkqFjDruOYQybt2Jdxe0KNWe
q5ibprq/2Ef8aYXaI2BqFTpOLKfNSkc+dfObTvIR3bE0vvEqlJwXkdDITfGDrZ28
IfbXChgyLf7EMeB8bx1zUx8VLbsLAMsy8yock2t+S85RD0v/TSjS8M9lkDLjisPf
JhMOL19Uits0ksu50u5hCqmpJUyTcOYyypBEpM5DUtITgsXrsZD/qduou20gLb+D
VOGObY91CG/kW2DW6bT3WYZrPIFYMJwDTh5hslTunJI4rltPhVebCV2XBvRpieXs
wse7S+UQsEZn7aNPAfTvxTKMstzSi555521m+COiUZFHTBZj7sWFWyE6Guxm1rXE
jpZY1v7NM5LwZ/FBXF08K8bdNiU7tJ8qDZvLV+KZ6fJyF1o4Y1oN+w3llcKCoR9M
onM0rt5NOg9g3ryelXWk2GTtbuTZuQBSN1PeROQlxDbjpd3i6+ODKDJHPtfa0YPy
x6wsDuKsfOBSmPqn8vAJPfdl1sAxtsTQbvCFQc/YqxKqjOZ3IE28NvWx2pybBT3F
nvpCyRZvpdMCXjD7uxxdfPkFWD/0u6UfRcWGmMwC2RL6PzcVq2YQlK0jTQOwuI3a
/5B2yn2ncuvbmK4x8fK7w8UDcxu5zC/inYPwACe4m8hAW4tFZQiXqmUK9vTEsy6y
01nM8RYCIIvlgtqDa+bdNDrHH1dMr7y48hP4oiCUyx8vgsikny3EsLEM0CnZpCFs
5IGeqvCHRIZPRVkmEsmYi4wP0PGpnfT6XRJyOuFD/Gw3SYdQrsxz4DKRToTFf2QB
dc3m4zuif4x0ew797cgsp/JSKG3d87GlJgYFYd6lPsGmlxT2G5xlAwNBFicABxSE
7p4Idj0B5LFPQXsI/W72a5jVIEoEZi6bNEHUPF9VQldJPBAwJWXKm8hG41co/PSD
tHL1M5GDhoL4cRbkKjjjbCLNNSmdplq3zoUe9GrMrjwhxSCOSSmWOJMwyP9Zj1vm
LasK78uWVMxrIXtIShzX3EBBSWakUiO2fJ67NyLpIFcNjm9ykb7WTCo9vIx/Wxqs
dAxeO7Ctt+dGILFryGhwFWCItB07rJIxs6m8SzL+IRSVrmY4ZZB7aKAPUnaYmkBm
w6l7WHRQRetvHdt0jdSkio7e/OuHGTPjh89viP2JU6izcdyIofPxBpVL5d6/jRux
c2qYJYPuf357dULWg6GAZ91WMju/9QUgKroZWSMyrjPIeP+3gpC3guMWW+Ga8QyQ
OP565pS6CWBageXq+tRY/wRgQ5hSv5YVl93WhYEGb6ZpbqPdsycLB4itbB3Vk9IC
3szKINzCTWWg5or4gx+jKmBEUkQvpeqEHXAPhHEVtrq5QGM+Phdsv0XSGToEn1HX
gzVllQo6iabTOGQr9u3xwCSD2Gr0C8lWEkY4ImZxgauIisaTYD6NGRr1PEaF9G/G
Tdf8QnvNaWTj8Ld1I3uGLhMg09n76ImuPD4WtYsQOxnn5NIydsCiXQ+QM3bVz2+c
GLZ/1OXTKt3crwzHtxxmADnMgr14K0KmSjIqswXqFRcnrUIBG79n9mMpiE8FPzSu
3SkIdhtbfE61ruYmRkyYrYP+Qy7yBVGTlUSvqn4+Gh4rA+DtJlES+3ZxhF4VCXX0
aVBQc2hmeCVq7Bc5uFFH8kLsu3QyzeTHTu88mltZeINggV6YRzt4lhAlcLRlYNaW
SxxA58TlBvDjqn0uePQiyhDLOU1qPLpUqr37C/C24tGyP+lP0E/dTVw3hJPGFrsQ
cdsDgQZp9HTe61BPbgetG53MRvo8plHw4+Pv98G8ViTo+s9ohrooXU3iMTI2QSoK
iJFZ/mrH8RtHn9ToYLU1DhVZT+rxl4TlAU/NuI0upXqoezShINM/fg6V/n9zRApT
Km9oBEpnilNQgwWtMLwgVWLR2yi+ZiS9fxHVAEIXpIYD4CGlJSIDuiMtyygeMyTC
6a96MtY/5RjCXp/pE/6D10NyE6JbSpaiXojxtcjocHyB5o/e2tPHH/4heQRZwqhk
1958bG1P9hZrs79+LmGWG3ZR86lx/EWzheAXDeqBS2Y4obLLn7mNro63QHHV6KEc
oiDRAU1lykiU8awum70ii3tIS4aGrwTlkHf8SOmdqpa1Vko6BK2gl0SxyhDAeLO5
mZbGmVjbG4WlobXlxUPibvAae7DjAb0A4rq5pbsTtQxKrLM1FyyPOwxj/v+Dn8kn
e1x+GEnHdEZx0NsTqIA0sgGk6s4L0T2xPvy2KlvreNV9PPetcauUCtA6sq+YNYGV
1a8dEfTXP2TTBuroQ3N6Y5XxSObB4GKRdODoc3KL+eUeRffkk41CYZWCXlwc7tOG
EGW4Db3JWA0tzrLoRwBFBuMxs58g3+6qEaskiZ+dPCL1z0B39hgvtytpB+zPeErE
Ia5uJwHtkrGWEXBpnPqAHLx0ewo1p0QPkdvEmYTLWTbBUaAYWCffZc0F9ke9LRYj
kamps1Hkopkgom2cA6ka9AD9h31pDtHnnJateiSstk7odZ1TRvKJAkoPnAM5Ih1n
8VJX8YlO8LMS4vLkkfkm3YlMxY3Va+4r9XtIi1gVN0TiHxYe50AP8H6OdfrQf5SS
GCHn5JAk6X8c5C3Eio3s6H7awWTojLRX0zJn6tZXbcpfAJ+1VkNufXu5R5tG56Lr
SVzQXzpISpD2KQ5bDLnZDLUOdkuVDs8ONEgD+1HQtlYO1g6pmZ3qmMrBcq40mp6K
GtO36ttbGLztiq5hBfPFMRtnGudTCyeNETFduvqUVl37RzJvUHsg9KZwzvRJlIPk
0dj7vs/bac2cN/hgEjEFva85zHHR5kbnL5rnTrywrcpaSa3Azib4TTJkelLIN7MK
WNRIdTxJm3tBIZeFKTX0rceToO8n9ulygxAPvE6OBt2kKk827xCfmeqZq5QJ+eJA
TnR8hlrGZdR8Oo6m4qT4JgZoI619SUkPdbeE+uqjaN/2UgUBDrNmaypNze76m+mm
tuSxdi7OqplDrdByUl65iJhD4i27PTyMNPJNFiUs5mfhC+uvvigcFtkpw/jKQff4
78QYtIjlAGUpC/1aLwccwuWC9dawV8HAkP7jSZJoDnowE/fovfTeb9QaTBHs2449
NjtSFFiwHB6beHo9R9ct4HOrF+afI0EFHVxVK6AxCHixsCi4/kBD0pVy1x8BnsvD
mgest2M8xW7lQ709qAFI6Mlw/wvLFxkDhUYFz3x8cjHHMwqvpMNiSGwH0aTprceE
iS+BNn5Mqbb4+PKO1BUDaU+HLFYjF6+4naZAHFBc5iOE/onRv9CKFTWOFEOoOzo0
839KAWcrG+CfndJ9DhklfxWfs16/JRiXAVM4zhBfbGoyTviBYsL6zhNFJsYr93Nt
zshq7TET+rA48TawrnpfvIa8vULlDEsCAwyhFepCoCYV2zJ3D/Hyp516VNaY4/E1
tL3G91ECeursGTudK8eFKkLqerm4ERf9cf9AFr6cyYfChX8EkcO1SdKQRBQdXUEq
Zznfe1FuGa6XdmcMwQLOd3qpijRJ4eBE4shZVSsRjxgbn6xBpkx1MsES+afbSotM
+cAeW9BiKq0+p2qLJtGNjeYiRjlTF7M/p3cTWeHjV9v7wcifZHxA+jJWOLKWvQuz
iGpRhrRFH/9RdhtXgHNtVeOe8/fB5m+UTBTGUhGsjSrKdqtdDLN1wtny5iCsnVNB
uhLsUZH3gNuxKdaC2hczNy4xsGLvnSzteKmCSWtOEtJD4LeyZJeJL7YROpMe2dVO
sF2qZx8hkwIhMlUz3nXfTiK6c42QnfDVIbDJIL1OYQstupc5TZfMIoacFkNnaNq2
+RsGiNgVx8hb63yFyrOpIlAQAK5+7NslG1C+TWa1Jz/IcXOPz44dYor5GqehX0BM
7P73TKP6vLTIIa+FCNwR2SbKmnYGoGdb7g3lgCAScbkCuCNFY6eB1YIeY8/M7nC+
w2IhTnH8/ux29pKt7V38BbQnHz41AOUiXqGI7a1axJ2iSjFgBFxLwr4YckSrk7ql
yzopklo6292WyX5H4paUshRHrnT5fEzom0ZZx1Z/xetBSXz7wBwsvS9MZeOgKM0g
HWaV0TbOc+RCz5ATSKgl0nrpj90us4SY8dbmgjVHavTgLdLN5rMBnFu4TtCWKHV9
L3+ylvl8h1EXHGdh382LpJ/v+TKm2+NWGHrwgvTW4YxWyPkj8xDHkJWUZSI+MBcA
310w3hsfjuc6uqx7QcsIsSqnIL51ZAaNcezOPZOvh11exWWA9UAkkbCrx2nPUDpC
Bhxm6/++oBLR3j4VXTTwC0Nyk8s1qr/G6Yhez0LqzqPadfMqAw5N+iqjjiWMnpMd
mhVv+VA1znnrmM1hWfMlYfPPJv0SL6adAvGyuV51onJ+03weIMycwJC89qMCL4A0
PQt9+U4G6eO+SGITpGIUVkt+uwWx95Nj+AWCUJCEb1puqINeHWRddaycTfk62rNT
bLIOF2PED6eAqUMlRCFzmnhlSaK3rsQAb/vbHxzh+awyP1y4xFrrasSN++vfJTXu
BsK9NE2Gd7dJq6S+e0KOTvFtm1fco454s17QKj7IkknrYRh51bRbLLi59HN+7WQ/
JzUDCq8OPOCydQXSLKIP2LJAdnt+XInnfsJO8zJ3/a9gWdOp7lLmvTLiWRCvWfbe
zOeJxz8/LVuEYo2L7SvAJmGgbNSxW76kOTn8VqykdBVmyFLzEvqn3MX1UYEhSatv
PEHIrlbe/mUBn6+BfwIXw4w3ldtki5sdmYjRB59G0yNFMwY1VJbO27xOX/7E84K2
J0YqF4uul4OdNnZT9E2u5g6uyFQIs7g3cHaen8QvRKE3oWgK0ieauhD9pbprk6Rp
EmQtk1DG746RhTYoEVsBvwu9fVA1MaNb9QqaU3oe1qnsjMZFKlbnFyPq7UyxuvPY
VtqjW7doDeJ4zKkuSbMw2TqVb1LVo10JAxjG5KVyCKqRdmxXqwMPCDUnr1T7mV/3
yGKV3ywtkJQxB194yPeoP15oRXvD9hjuoRLtyX/TsU44fSVnc8BgZyLe3wR5cudb
2FPU1JV3b7q7rwsKc4hIyso0tIWDIUDxJkP9PXgDQ9SgL+n7cHt1bIcsFOtnWAlR
lZCx3Or3155nYrqH2mYqygWSkmdUttswKhcn2uVGpXTnj/hX5NQd2bd46OmUpHor
vspAXtPTOil/rlam1rhRWIpZp7fQBkJ/9nFSFh8GzhG/Irk/4XJHWl5emY4KeZ84
67WNPPqdavGUfPyfyBqqJRLLghdJ0dJ6A5AUtTSUz45U6UnDTFyeqk3cgk526t2E
s9+m+V+Yg2qZ3RsouA9K9JDOk7eM594SKbsPg8IdAdtTwS3gaVqfG+XfmYzxfTTc
buKdJQPEViUSESsLvhWfnwWvZJZZ4wGw9EZniKyOQAEMjz2JbVDFLyb/Oz/VxZCX
23qAOc7McYnjnSUQ+S+w2vpkaaJGNu2q4eI+MO8gZeVIpRh0yLFeW4T5RSLzHeeV
AerLhcHuWVH2Q/vSZ9eA+hNZbjxzAXDExerWuXsgQaMcjsgZAOIPS2BpyjVhgIBB
PCQ7hVCGF0Ztiorvttzb2lhLYe12w0WvHOJ6VEzrJSNETyw1Mj+z1IcMiu/ZSvKM
B0d8MMDE2RmpwhkDCd0FFvPcQ9usclBrOK3DCazyj30/zC55jO3XPxsoHX29RoJ7
SYtJ3UtcALdNG8Fb0xwNYMJDI9Kan1z3m8q6aO2zxUecwQh2pcslglwlZLiOpzRP
BIhiLQ4v8rNRqpvWatjhVRNlookRd3RwUQvvsMjUf4oaXWkR1jwq1qerhYTNc0vm
vhlKe9KyfmuYSO8+Qm0OaVMqiqer+SzxUwwvKlq3MaoYsRx3iMmYa6lPtB+tB0TJ
jYKj+qnLrpouRSmNikz26XWa2JdT/2B4HcocSumA1gYW156CDjmi/zF0e0SqccXP
4v03AC62sIQUdWYO9VzjZtnhMmt4An/tuUHjE/M2eVLLPbq0d+WHTI5v1pdf2ipC
c524nM5s8I8F62ORGJ5HNbUcRz4jD3fwgNQgKsO83Sd5IwmgQ2PsXa9RbRq4IaXe
aD8iz6SoBA+BZF5dAMyGnbrYIw39jekEUtTfLTr+ExIBTc8dTZCsUFOokHm1OSIS
c64iAMqmxXwk/SDp07MxBojfKyFZC2c/vKO1n+y2SeaZqLjsuuOK0IvYnYzFUrzr
ahzdHAqkSEq4q/rcpfGo/4Y+ZSPEIktpUlSR7kocFiPENGqCb+90BKMWGu32u2ML
7XcLev5pmJWWNSKJx1FXdU1v4f4FiR9Y7fCJZiNVxeVnmeavlNtvj1Bl1i4qR9Zi
dpyxRo1KRXqgVRfhWFz7IVZ1vKfnq9IOXNOpJ5htVrspySwNOvn3UPhNKZtxnv5y
B9q5QR23kh8q+bKOXFjN8lptEAMXXw/cXkbeWpHo0xBmgxi2fqnJiqHiAKJ+o84P
h4Sff+9IP7zp0CBkX98Z8nwaG5nMCoG7jxlRec8LMxlo6Lae10vlGEtOZhybNMOH
Nbrv3/rWJHaqOauwIi3dz1cYfxrv1H9v0/kgU4LLt3MMupkYmLzoCbvnQbTtZRTF
V13elb/FbMb9+RdSjoNO236T4UnnUlE9aFVpxR5+if7C6mDIE5OwuGo7vjOOeGIt
qicpddLz8j/4gI780NJPPOw4/mwRQ/DEZ3FP8slsA4PyZXB5HRsqaYRYVoengZSo
gQLdIW0hrhoAVKDaztPniegfUVevCIkWIMQxfGtMtHxouk7b1ffcM0pj5XAdOybn
DpaZzBlBzbkvSHxlmt+UUKZy8vNVJscFnfaZAm55ZgdfiU9wVg+6vlnJtSJX4uqy
3EyD15R7nQ4FdTtrOayVRcy7DyIytgaqNbi3PqeOHWSrtZp0a+jAWLVVyohO7BTb
Hm/HxpXkAiN7O0g9VQztmhulU6hK4NZmfXtYOJHEkz3C8MpV0hzbvzNexCiEe+U2
vwx0ztm5smdgd9KholcgeNi4dSVy12HAq5lgBq92FmGj7Ok10+1eADumd1L3QH9S
b/C/oaZUB48qMBCClVYITxEetHuZ69BGsWbeQedWfiVAapeBkeLYjqaOmbrjwlD5
kMLTa166BRy/9oz+aHamSBWOMWZBeo1IBoL702EzYkM7RLU71soZYZ/ey8wLYXZ8
dDLVbFIJS+TSjOsRVgUPX80R1K3UEeJr1iJV5UqL2xxF3bX2fx4qLEUhlAn0qu6o
DX//6NV0xxBuV7ltXPALWgP14QNPTrzTbXS96S+tDeCYu5u4ViH2Y2FiRHUPuV2s
mmf5AZYkfQ0Zbga3M7jk11QUGb4EO2/yxSCpBQysrqQAcgN5bGJ0NXdn6zt29szx
svqSo46C39BqECllqbE8KUEiUrq6qNge2b3xAD455EttHP4YGXmgkMZFe7ZjvQVr
phJhHq/Fk61b+VE2Br8SxMkbM06MjuDruclyYgS3Ku2t088m2g+7T1jOeg8lWEfP
1PmXUuGHSYJhlI6ZV8pMKxtzkbTjl6B1rWfe6zwOvx30sPclhCccSJnaCXpqW9jw
hnlvSS2A2PjupndQen7EO9mqimo7LIuswDyx9jr06uN5S8EH+WarMfDkNmwPrO5B
sQPMwYs70K7KRKt19hL3k4R/EDdLfw3IrFqMiyQTTVf0ZVcyDqFD8wTpiL6exoFD
j9Xfx4pkn2QXJf05my1ctntk/SS/rFCw6oTJZF8xRlMBFQcNWxSTk8cUXo8w+GYy
+aUfIx/646ynJJfeReNQETx7silIPJVEs/S7qEDmt55OROSC0vBTIj0ZdXcvj5oM
Hz5y17TYWy9ZSmABTf+s5x1tU2M9YzP+CrHcusktu5keIyEANYrOhV5M6ptT23Jz
c0CWbs5tMTOe79zvhOkd6PRdhCruF2qFVhV6Ifk7lJWq6QgTHNfeMsud0ttED28C
z2KvQpi3VmcKqzt7E6wNR0FhbWU23PGrm5x4P/LSJL1SBWtzNp1NRw8yn957yGiP
/UxxNux4hATA86mGxTbT5MuMyvuO4QVEVcXYCyM+2fE85g1qD6sbnCQkwbnG6T5y
Yrei/f60ck7FT2HGxniu1XJgKBenAI4hqE+rJbtwHzm6KwVQvk1nG0p76EWCvZve
TMpPqN9+gghTi4eGABiB/FVTEd6vH7sGWrgV263lW+66LHUubpnm1l2xyKo3rKdc
Q56LSOg3KhmZpEagMlXqtsFI3un0LB82wEAbiX9Pqsfhg83jbQ97Qw1ZRMtiENE5
5KlSckxSY/V4UO+dRNcuOPVbX4DDI7zMXKE+KBOAB5TyxoFt8injInOlyg1+pWS9
V/0Q2dAPxr0O/oipqEGJWkFSoh4RLTsniTPXw/zUr8WPGo06Msl4keAQ8gwPfp5Y
AWxoOadrfzBAXshM6Ts3dxIBvcMwexKPbCEWayv6/O5NTeKTsPf4Zr/WM4eSBhOg
H72+RDGH1ykmzaskcuVBDptqowymHPSx8qYBES7ZwNOZZKFyw36RWOtED3/wu2Iw
GeNzHdyjKdT7AKr5qQHOHdV/dgoyag84FFlkjEKHJg6PJtIYc+ZQrCGp8+I5/kPK
bAKrsPzmmKXCnN/JY1u2XkUQcAKiRIbrKSA0frk+mEXqSWMw3hEjZUKKcqEiqALc
TIZMsSasaFaXgowL9VebRsSfjcrZvyDvmOlrH9wVsml0Hk8traCN28W0cbwdShq5
oUu6Zooj+bk0FN+f6bWbj8jYzUoaPgczRBOnUgqDCeJtbkd2ykuyT34VdIwW7VUY
Q38StyClXntMiv3NlH+8PQWkP/DZYNgZNjIVZKcxkPt5CbsRzqZswoFowBtAKx7D
rmzlUUp2iszHS3oWnS6i8R7dEWPf1fwDeHAMCicf0jsdPer9SxFABcgNwPZIRhLk
1vstP7CAZSZIvJv8mAGocB2VAZ4TCNafxxAv4bBv2xykEW4uCTd1Ivl0CzCY2RE2
yQz9Cop6AW7rp5yu8mWbsp9e3zz5QFP4a2qNsZy4a07aoBh8CDuCkBmocTKwwQQU
NsQGoV0lNDyHyNMYpQmPS4lVQu2EogFdkbTHxDIcKqMSSeoe2ST/lnpWTo1FN9M8
o36Zb2aTa2VJrnYZRRN/MCaNpjZ9a1Q6cvq77RECYapWTvHyleS5EPoQgi7tV+Qf
YKAuSi45B6Ss+4toHBH5JGSDAgiKT+X+HSTgxZ2hpmWWHmrDzASbfpzq8c7PfROH
ixdoMqep3TOihGMqjL/uWG78lkf/KBS3JLvrippM/wfP2y1b1PUxv7JwvXyjaQLs
h4EzlEPP+SMQU1Q4+8OvJMYUY164tbXDfTuvA9rB0C9cehScEv8kHIM+Ktfbf5Tt
g6n04LpvRbBcDQu7Ggyj1UelTIEmM6zgcuZwO1fTywazOOQSAP3kh5unUfGt5HX9
SkbQxnMdDbkJYfdQ46hq40momD6CFQzC4qKKQ+f4tlBLt9/G471I7d+/6ibwxL4M
R60hAsk2/16iKjMODkW4PvkGrSoaoqv2mto6fBrgX29sTJ2k8XnoL7/5IDQnmAHi
gBePaKX0ivct8Dah2K0k4Vhgq+/72XkJCSph69lnW8zaWiUGb8BzFlJc3Eeiyrmj
aPBJn0paH7NH7p1gLVTk3nlGG64S6RB3gxLRYrLNiiw5lgPBnbv2PqWP0gEppKNm
7piWC7pT+ECBI+T2wlyrWPY+U3zwyQVcrcw9VR2lkbPDCmnCrWeSNjGCDbsQzHWH
wG5qwqdmtHgOtN4AKFC4sRDvJHSPokjzDT3CUFU+clZTj81eaGvOK1D90JVeccBV
4mZQN8P9yDLncWykTnuc7u0MoSEqxT4jXwqdeGNO2y1HQCuxpagMs7DLIJYV+iVM
YE2jtilypP74rbrfpwIQJ2DxEJ3cS04O5MOXWvDx6JIfLXAP14o7fRlyr8EYY+2j
Giv7+5VIKQ5hY65HSZfjQtakQ3MXN7ygJgKrj7xNFMPoxZk9xkAUgJhVhfDPltBS
o3CHR8JdwdM8SWibQtDw5Yspcd7Y9HBngvX5hwaBgsxY9gGZ2kqK09NyktaGsBKm
6DYl9O94eBJ+7UGpKPnY9Xt5ZnyCb+xFFnxC4QjNnkZ/Js9HBi2B/W+Ds612SPVm
vLOXtedjR1aVgCVQ6/Eh/yT6vYP2jbe9i4a14UMmuFg5+VftAjPm0qGI/4L0sPOB
JIyY8LyHgSVKiTifneitlVfEo8veY/s0HG4tvzoBvyXbhw7TCfe8SUbXLI1/j8YX
BhIyUgMJrtKHiUZEM4pv4JsPWH4ZfZkYuzxrkCsvdd9kk9Pm9kEgSdCeyEu39acQ
I+c9WCJjV5WDS+wQCm/07A1nD2GHDdbHF6jiFPA5SfoGirizdgSIxBtIeEYxNc0A
GECQ8KxUO8okRS/Hf9jpLpsa4H0HGZozIfg6zyNYZrg/iz7FqOuu4vzljALR9P3W
zs6e/VfiyLQ0uhdn3FWpWuDdUdfNBhTrALf2HKMQdYASq80Utey6coWiS/uPJ9PW
wDtp1GVtPsdzBzLWxeWyDOzC01NLgHpnG30w5Bdc+YySlA1caWicahVb6AaYtRGx
OrCzCq7ue8bcLZXPd2877UasXN6C2VjSYseKMHqAUS84G/2R+M+bLrCGPbizM+N2
aKrvEQTSMUCmQSES4PK2erERw9AgqTciKAA7JwmlUZfR+NSBSTCmrp2MwWq9Pq8n
aR0LuEQpNqA1vQXNZ+07KDemWy+P73GT2xJPgxmPg+1IUywP19CX0/yQOs0c893a
oZvcOo9M8GYDbRuiIhMkp5k3C7IzFX7qWerRXwhW5WG7ai+DjK9LpMhgXklYLHy+
SWws7GMxoKsQtwEu1c7TcVr6DA2aG7LVgnzMXPLv3cIdbryFLoHgeuhNpAhTDcnh
GUfmXv2G5RC5rNXmN/pTPBjMm6jTS1hLlbiBoJKz+rYH6v7Dc7E1KJEvbXG6IWE9
QCWYxb0FHgEk93MswxMQ5Dpw7kzfg/dNc4o3EHu/WBDYOFbElfFDntuiIe2YTEDo
HBFhN+CPeFBzOSU90pt1IIoSVm7h8Q7Q7d67YJyOB9rmkwuDR1wiIpsHP8EPVwMz
bNhDJdlwp/t10Xh6y7cmpN01ceJgEeXegq+iyPKjpFDc7pihTDRc/KFzKVhRuZKX
l3M9D9yFK73EbMcRsm1Wl5E6xcF56TzpkmMEb8elzaUO4Xqyv+oqO28mWbFD0HEz
tD6xHRlfBP1IWI/9+R9wnA4M3m4zxRRFl0/s6adLONxBspRfJ9i0ip0Zrhidjoo3
cqexRMh09xwnSWTE3Q32vsnGGfnOHYGoej8nrCVBJVisKOrHUJqVBtimcQ8tJ96h
FgIY03qx/MTzZwetLYwyR55jX1X0ds1RokFSwWzJutR1OfOxDxA5EU/j+DUAaR3s
UVVg+KbRlu4lvHNPXdHiG8QwSzMfXdfroSRjDk7hHxU8tMrw+Cj3fMFyqu+GvESJ
hufPyNjIbDlf2v1nyu915beCiy2uC/SO6woytHOQ3HUQYe6t+KxvlSbCnxZNfdxE
UC7JymXJ331QW+4RleDZ7rSALY+VOmdrMf2TbVdtCcmXgjynYgVbyPHC/zy9+Gp5
jjYc1KQOPiHeKCagE/LWlMKiXoXeYFPa4kixI0FaZTbjrBwCMUdwSN0Z9RAFSGLa
JWUvf2sPBP2PeKmeUqny/1U6JgRquJDR83yKSoSbtYozskPpSg9qLb8EF7YEhTuB
Xl94TK8J945Qv17WseR0MhW7lqQ/7V3XR7CTmoUy7997pO1yDFD66v91MsubtE5E
7I+aykAnzSJM/0c2ef4UD0erl/j13NmI6m3wm0v1IJeHWkC6jl9PUgsMuXlYGHOY
5+NrCKLBrj0KNZZqOI/v1KUKjLNrTLD780v7UEY9PKl2x7JvFiL30V2qgw0MK7bt
79CTawTuVN39Pvuhsfh5UHml4yct8zFx8bg5WAcpswszeMM1PLC/LSpXiTA4x86n
bSYy1Dlc4b2BMVbnmHRxYAiB+jgep1mLdzXAe/202Mlx0BolrNT8KrTs0kN5AmoW
UxtdVur6DgPltH2kDo6tWLWUnhSD3x80k7Iq6KVkVyRGNv1TDDSLlYIjZ334mtee
ilwOUdzqMndhVEgFJrzhJWTPi9Zp6gC7Hbz2AeApFMLZOIxGlCf+8zq55Tbg9H9Y
0LVrMtV0pxDAdA4M/nSdpi7QFVCzUaCUzqVu90AWFStsJLYFh8GRcOOKKX0IAisT
Acs00adzgeh0neZpQSPjciZ9L2Nc/r5GarF+CuVyPIqHkQtB8//P499kb0BMIfaW
CZI37f1FyV1zEctIeODGq4i5CDi8u+cnXF1F11/kvp+Ai7ioEx+3T8Q8Ko+M7YTz
pC5LWgyg9IM40Y7Ae7HaEOs0U/u+4rVNLtge48xD9XSkI0TiCRNU6j2/EZP3FV0e
4avoeKhyZbA88y6WO3CFFPw3ODXagfXbD/hfR7JtcahkQyEkGzKOwbyrILg1tBPx
eArVgFg2nV0PA39BuFI6ep1Np5tPeZuE8/xu/fEbkZXdXOjQwRO4r92d6de8X8Nl
ToHNE0xVVLGR0Uo+S8EBT3kPlcrxVG0L4ejwbeRticUEYQVBErVjHyEGFTsy+dBN
I18dopHr0+pDQk1BqaPPB78sbi9nrbetSgz2mMIhuTCOtcYLXASJd/M1xIAg0I0i
AF9/w3WSKZ5D8Mw/atz+vIWr1ZAQuxzfZkwF5VICAqCwo4jZfeKosArkv8XFknae
+tib96GTpIHYQPLz89TlNGziHMJsSvoJgAYR7ODCr7X7IZbawhvrb2pmbPEeyO0/
Bca+UXfL8vE2UZN5tlk2ZSBNZPnqb79FhruAD2JSO81OZ7OTxKoPY6YFOwhrZEP5
11LroxsWy98Buwh04uygNxoe+4uvLYQ4gNpsHXN2gxWILxOKWqx334VgzpWm9bSw
Hh4rfEYK9AITA/v6EZh+zOtEegkrlGX3l++SBlyaqR1/Vkx1XblhfUBj1SzkApyY
ficRWDSNmFypwc6iXFAtdsqWiL+Vx+TT+KZBI7c/XTJ+kCsHcEn7VuBrIxtag07D
ItlCTnTnHn9v3bu2gOozvNnGKiwZJeruh6Z/zVDRggo5QtQa5jeAq+08mVJ14gYB
ewZ8bG19EwC96Fp/BHzKz9a/sAzspdedgoVp5IhkSlEXIfkk9tOupIkHR34pP1sI
v/xGroAux9bxqO8ZELCuX9o6r25LxOkPNcbm9hH3G7YImMbq9GelEyo45LbW6JFC
qbguDUqotA2SqMGYnQB9YxYb5l97VDU0D4knnuzLkccjpNX0zOUPHyi2mizeacrs
eGkRPJTKCr5Y7hBLw/DSyX4YW+Wr8giRVDn/qRI64vX90FvoiegftMTBk1MQw1Hf
iqtHig15a1XzS7jhs2UjkWQ4lOOw45LhYhf7r6vhz25v4/EzcxGeg8CnCZVksJOQ
1U4iWVQpyV/8oU8dk2L6tDi2J540M4RSw6ZZsbNiZa8JnxaUgQCS8Svsj7nVOY8N
0o76A75IR4dSVWd3ss0Y/BqjluiWnPCIvnd4N/GT4ru+QTcj+yxJt5uc4IC/EpDV
HeAjdSf427Vr5r4GUtnYQ6lxER+891JF/GlXRCGfMqepJ4X/mfQsW4IfQM3GXQzZ
e6+47UTdxNSLXAQ+XJdz3AKHxqI12AwTNYDJkGUzKJEKoLlJFCIzMxQr4oib4UVd
go0koUWLhkclYKRkNuOM9s8QgxBNp8W6IBXpjjj3M3UNY63ybD5S9h2CoBaun0oJ
7neI+HbpyM1mmLQrtO+Jflm/p1eVc8QjTovSkLPQDGfq2PsbqzOFxAcMeSVAYEdh
prB8WZ4G19/I70Bap43FaRpBEY+OtjQcib7FjFPmV+64v1GXUIilYKfR35/1rzP1
TRlA96rgTUy8Eqprt59VllW58nCNahri1mAmuS3rEfSBu6y1IKmAAiPlGZQAlHvz
D2MVP+KnEBDtsJIF+kfszaPms5jUPMV7EKgtmAmd4VpWQI7NvTG4+7JQD9uYA9X0
j+RRuDuCXKxGlJfYISOsdCPK43YuwRPMEvg+OPZLMnVq0sv8chdfcUTsm/HY3f01
ZpB3/9ih5hBWtfsRGnSBj4hzGT7Ot57JlZYTGFmdJYcuSWGCMLW4wGsDQ6WyzNDB
VBla3DNbXebViKdOIvaWX7fWczYcVZ34TsAiHl/gjFaFWuAu0YHjVJWfPwO8w/CW
G68AKLjA0SuFXYdI9AVEzYmlC+k37C+aSO6hG4QX9BNXruRy33otMdb9yOcq8OAS
H/IrsC+FQfkVc+K+MQ2r5OdrcLc5pTznMCODVXlG99Erm3BTqeLF/+LJY3bvMYP7
17bq5TBcyEnCNZjyXj17U2EK/hh90WsSMqHUkFMk0dnDshwcG6HkmXZ34v2GDKH2
SgEDmwBJWfJyygv7Iid4QDO8kzGBFljwmQV5VwdZNAvx1yfmwnCQjAKz5NP1e5IL
Ny05r466Thj/jw2ANOlEkvhAOphVcSM/ssvZgRhF0s0MKpyYUmTvTFYLwfGoRpMt
1fiQgXujd3EDNSDyfua+ftl3qjCswJ9W+CVYXI7VluqG3scB0SxJrqL+MX+PsSNf
19A/gWchegKFbwDReFxyb0fdej/9RKJQg5f4D5g59HSJqtBFBd0NMSW3DlSRfzZv
+YoBG/88ylLsHnK96sqZ4DoobuU1qMsCZmmOJqsO8mUfQeUVQPy0KvztJyxXMsz1
OyfL0H4iaROjoc6garO9z3YhL+tlv/pPXx73v7S2pS7Fnu3tT7UZz6YV54YViuRG
YH+9Qfs/Xs6ZyM+twaeMDymalT3C5YagiEf13XDgS00B8kupTEA1jSY9I7aJDCwc
Hpt1iBYiiY15MmU65h870tmOd3KS5+LihD1F6eE6XRxbXC0cUC2YCrptfui3yNmU
1WP1WJ9MzjHtoekDa32/gIG5PScuOypb9aukFFyJ1oX858jL5fwXeHSFOmF7EI/E
D72izLdV/pfhvy0AX8xUnqdOtlpkVHCtFu1L76PlFCz1A1WPCUokQ3/QidhVRqaZ
kzbAZUw4Pzka3jxZl8kBDXYPUIAoMWmFiwfIRcmm6iE3eQ3g3nUtm/NHHVEaa+Us
PHTmPQinpeTnoFvIgeDQoyL9FBknFIS0NAql6n+5UEM/hFZ5Na60xzntBb7vsNsH
fSDZaT07g+LUqw2Ch0mnBElXWuFqF3svgPh4ndcVKrzbhNhQ8JP8cyPNRAcTcPMg
QLqtF58m2jrFdCnQh2sl6kJgQJI0bWf1Tw3axKV2DZE60Ab0ia0nO8Rb7hRgEFg1
Lr08SUqfthQeGoOCiSq/TarfzRUoGto1md+VWCPBZRc0Dh4QqaI++i07p2LIRW4z
I7/wY7w9OPYK5AVw/uzrzokn3VQAxm6IE134RrTFcRqL/QFtStzdfvbMee42o1bh
+USGalXSbQ0HXz/c8JApaWKpGaQK8rolqHgGETeiS6Y+/TXWahCCG7PiG7uqIN/H
1SHCSlSSA4mOzQSDylo9FP0+CTSQCoPpixeXzb5Bf0YRS+sQRcdZXrSw+j1vCH7U
j3atLCT6zjK4piHs66/A9H+2ncSZ0EnFffdYTSKbiC4bTL3EoXiYiNUkry1dsrBf
6GpA7Ch/v5uKPvJ71NqGGdCbtdSUXuUcPPDlN8ajWN5ybYnUv2rTBY0C9M8jE/qI
pMoWy5KzqRPJKA0XALlTuzjLzkhDIuDsztp0EfLMiBNuYmL2Mw8opX5TFpRBKa8Y
b5Tb9YckfTHraJJbb1dJVfiuLrZSArFs6Ll5T28RFwraMUUeLx6mEJ/5ScMskHVF
SHgU9NJzzNQiKFnaL+o3JgmaA6XZNQK9296W2t+FqSwyxI36rAvE3GVwchYY6+Fz
3j5WpjeCJJZHfHe/ZEqea522RUp110YrjpEjBAzA88f16DBcOlWg2OcMyySOvMdu
bXATUsLNxwYHyHKJ0BJSNTr8HFJfMzBHOnp5TLm+kpSwC90py3mpqqo7iUEajjtP
a6vYJCe+xlBoEMW7o7oNJ4dbuz+JFLhHdX1i+lRUyBxewyv9JeOHjuKOY/uEkl8K
UFNC3pv6XAkq+OwpWZIVrXOOySyaoUfuv81JFtaC26m+8D7EFKeYYEZyUvo4XO2J
01Z0nV2iJ/zG0Iemv7kon67fHxcQ8isloaZtE1+jYtH3HxiLe0SEePLXNpa60z1c
tCMqUY2r29ktuPBJV0SxO7FU3p3t+yDvZ6KY8uOWASBXCQpmod2Ply50CtN8qrOY
yFhzZ3fSNrn/c3ZAE0Ny5dyUIvZyELI3Ab2awj/hhnpZPVTIwbGeSykZ1lhekqmM
odS2GJpMcoJ2Ue2SIRmq0lXSqvu2n5JnE+t8iIUDiZK49FXVyUIjRXBhKZZiVbyu
EmGzYcnuW/F9SZ3IzLqtbIG3/I7rA82xv6aHNEckjrmlOkuKH43d1a6nrDZLYVEV
Uuc20kIW82zYCIBUK+HsH4i9ADeNf8WsxippDB7JAeW0rXthOshOotPs62tXfoD9
NWAWQyoamGXRMlXp/0LwQ955VxE1lex+eAGTnVjiTfXukyr44irHBmFM5fGU0hF0
zWt/bjq9HMJoLrqNCGR05O5I0P90WxR1XiWq/z5uMnwE8KI6GIjOoVLsUdzC4h4t
Y+fA3f9MPlghun7IAL6aaF9b4hrbnFoBvC95SiDAOfvpzxHivxuLx9cbqoUismJn
KQ0gEQy18PZTx3RmlZ+4pVq5GbVt8pCpPQ0QReHvvpWejp+etX16zaJw6KQmRJXv
cYrbfbKaVJ5v3/a1vw2Gecg9YTtkIedcWNRI6nft+xUV1LVKknwFXUt3VMwOgwCU
Rn8L1lp+kGUalIMElNtGzgN/v2VPTzUX4nVTjRBmi+FcQv+BgDVJLJmJM3mDUerA
P4ORPPT3Y/Wv6G+V2RjN0d6I8TJSMVEY9uA71b485q4/MH2JkWWTo8gZhNAEDkl6
uWEvTtil3BuqbnpX/giiQdRyUn6h02a1ujMHExxPVb9l5e14pCivzWdVnVpaJ3or
5g8UhEsUvO5WVxXxRGs/sAeCc4ke5sPt5PNpUy/t2cPzLL2x66e7l0T9Kp3lbGKB
MuHbji+sXrp5ssIjJtv7nO5tFOGrZaeGtX9LkMXm+C+nIhXAwU4WuA9G2kWr2Dzh
9n9Ks9zvxCcDaPNPyrsYFyqOXoZwdPebFydvod3VfDApDI7vbVxxzdpfDadmaFIK
/rh7zBYYLJfsd4vAjKT4Mu5cd3AooDGmevjB8ElKFWPO+ud/1lHbge7Mh3ft0w4a
vMlOOqaDo3ZlKxE0SR3zMeC/D9hK8iV2qL9LEtny1tINTuGRGWBWqUl0RVN89uQy
JcCI4hfGO3BwK+ZATeb70OPKEk1Rg4bY5WJ5+8CR7N8nF9ghTTsssNq86YDRtKHt
Ecv3oXz/x7bOPv3VP5cqkphSOtGIwU8fidXPl6s7+m913S58vmL69lIezzWyDe1g
q1m9lw49OqFYgiYMoEoGnVvnhdEfVQlhbfvUauBW8xv5qIptLx734NVuIy50Kn2A
Vswp/YnuBydzZUolbMmv/b9doYcjmNC8u6TtEmPzU6vTMZgyw19IFgNV2dt2lKID
JLxq98ZeYE7thFkdR+PjtMrwKreN2xoSBCsA6eBcgwHbOkh/L2UioniHd9t5MEeC
9IPTubsXvgV2hAWM5SK4zdBLwJQb3mxx5Z9B7iW4PHXExfDaGRl6JHcb3tjgEJf6
nJmbOdhqYRVZcd785uvucWSlvtOKvQQ/LvmQ5v7zMfW/nRAObOZFpp0dlyUoT142
CVQb8JQAwv8kXJ/CUOC8KE6wnLouuqZdaUEDtPy5cIsok14ndwYTigoQCFJmnw63
jWO1dIH5dNfPMEAUFR7sdMXZLQSyQkgK1D89yf8uoVKaSK+75AMV7q6qANFE+fXT
9QTJ3UNXKG3kUoICLgqEKx4iX86L5Gj81UllUQud7ytkBJkpMLyrxBVpL+9Gkwal
oM0LRfqsnMWP4SnyWN+/ErKRxkCGdODL+fSLAopAwCbu6/gvpgQ9RAo5tUr3lBGR
5J+tpzQE7NwZXjo7adzhuScdmdMFOquL1RM9Ugx/hLvQ+BFtU04+JRQl/XlqY+fq
QU2d7p8ZZHovb6+/VIPRJoB/ImzH/lVDhGnaOBjxAYJH0+5MRyb9CZu4Nbx78xB3
/LnHOmDc26Bv3tKpglgTWL+eaHaFWMz32Uj05aQXdGDKFVysoob+fwmfBLWmZp+r
sl79xcn+HtZahdalH1wTa2HmM3VcSLAEe+Ay6biHbz/TjlrXPUdlZGM3qJ3iga90
TGHoNYP2KFnmeviUlpTlgq3gDjuxSvu661vhKA3LVKhgiK3usEla5QaW68nhZUsX
VgNF37FlGEIs+D/+ne/KSb38EsrZyZLaT961GXoRUbHkCMb8crSI9+23dZoyjSio
MOfJZ817wVpRZC+zsYkYmhbOvOfQS71DGaP+430PEjGamBq2Bpq5nkAGzCXqdGFI
f5MqKywBWi9GLc/QngflCCAssLG3EJ7KxKcQ7Z/h7mGqKWcsl/TelWUb4Z2/6p1Q
WoWDjZc96zFxMcOLJb3Ch/DuAu7tZLYuhl8g9zJ1LBij2qlnxW6WFvKQPTapZ/Vq
BLYL4nR7IKeOIRHFCLef1dSIWXy9pIkALoACNQuezDHUtea4dyYa+KR6fyKkUkue
M5Xi6xz9ZRJXEm3ORc2apo9s0kiaXcWtcX9/zHrDa7lxseJuHj87sQFMEYQ8S3xj
GpFy74wsG9CtmkhRrqxC0By2wXZNqhE0iCM1NNJv+FcihzGVSsbwUHg8ALY/O2A1
lT2vv46gvfxpXYkr5tPXAfBgPZmHt80wJhlAOBMpSWGHLFNKguCfePY1UG5kGUtm
cGgnYLngISZM7FtPRblj2+7BahKfZdvTBZDCehPgG4VoPzRQS6x1fgeun6P8yW9G
3Z47UsuBvRwLJ2BXweeviXlILLUKMl5AIbgvyNWNR6kx2DHVJkNjtXCWo20GdQ99
HI4gp+uNyWDUmpsGaKjWMUPdmjQ1wCarBIs56g8rH8r+qhO5knU4YUX5A9sncKkY
/B1VJpriYZTWc9tvASLUzUgbS5/eSL+JoyhsTnLaiYfOIZ7vhWiy3jn0IxTYkR7c
6eDNCRmaQklwzCC05YbTJ9KoA8lVJDuUH/8DWA0VfpVEBGLdnX+QhV2kijsqALrn
ifHvTgqiAVk9jIDDBk25Dns35H1egJrWvuxmjhmvklZ8zsdSiOCWws6fPfG1Dmue
zHoDWsqMxbAS7egTj5GL7Bmk+VOVgW6JASfQP00GK/qMhe0s+8hjkNv42VcSgYtX
cG3lpAelvF9dbx/VPatag235f3Fp90qRYnEnM1BLuNQm64qybCXuTq7edxKVpBQs
FfMinaSakppmGxz2sGtsOlTPV7nf4fiOwqcPOhTsaDzp0p3Cl1EV0lj6SG8YWAim
Zs5tvs4yK8Xc8BaqCx0QcdLawrsuHi0JlpQ5Eir8mfmOT+4cL2gBpDMFeGG9smZW
70/wilhz4c83sm7pdRtOUxVkUSGB50YiAH9UP0eTd9TV2bo+LdHRVpOqAs1j1Rra
SzYPDHcD7Ktt/GFeWsS6qiGQXFQ74y+zQIm3qOgPOa4f6BcnjBeOTS2+h48RKWTp
cB4XWJwxo6G4loVHjvjP5xfCP16mMAp1fg/kcYNsE5sjJnYLDFiRPoO9Z/HHIDzg
Dp9e91OLnZ+eKF32jhbTGnOWEm+Edttcq199yosiz75gt0BMtvJ+GJY0iKQBzZlh
39cvvwAm4MNVic44DR9AwxtOSXfCkENVJK4DCjWia1etdT7/TybORXq+4q7niHWr
i0GwQVzGE1ANm6/eFR5IhSN36esrQx2jFJW2ovQRV30Yu65NJreqsLlSAMmgzpgn
Gp1r+GDVcQRi5MkQii+NS2PfHSpMzdef1T2YPL2rCIEjIFiRt7Em3IRHOeUrgKFM
DBOgw26hmayDD57huyht+wF6/jGMcB1Lyfat9f4EY8RO5jUZP690NNsutjMtkbcO
Hw1yS/wUjDoh5nTrqOazzW6HHGOJsprKb9agpOTUZeOJZmHZ71SEmgrdcopDU1yM
FB69IQZYcDucsCQCZjFY2ZjHzNZikGvc3Z4CrKRXZb8eyJu58d7/HUBppJ5XCPGQ
uJp1h/yWp0lNKz+hJSt7c3dFDQAN1X6byUMzZUDEZN3ZwsbBF4a6BqP5DHfZPicx
oO4l/cww7QThht3b0fXbFFadnkZ52FvEQbBBiamlQmsy/XuFSxZMOJJ7pgfpjEbA
B+cMMQKW1fBWCvIF4zcG/N0VROG8YRJHrZqPmWffOQzgwzP965QHsnALTGmjjMhb
vttlBnJWPYg+wv5/1txnm8GLAXS6/2gyezdHjEyMOZNFhAkk8ris4Y8NdMx7z4eU
TmKFLNpiJtETXR5u1PiujGnb6SM1UD1t45OpRthlVi9lgfJSFPcWPWDQdL9ZDE0q
MYGnK6ATE8EgDtyKj58m+D9JdssJKrcutJaS8NipkWOxkAAyYOWlwt/tqBYD0el2
Yt67rL104cvl+KhGSYt0UhQGFJpqD40HFJK1bY7ikM3Hw7EsBvqGKLzukl+BSFYG
nJmRM/GZ3P9Q5/QX5GD8Jh6ZgGw0k3ttO8KbKntrg/srJ8dC1p46n5qF9z8hp3jV
Ga4RxsWkOPPAKqujXbzW6KZuca3uj07o2ls+ZlvgjnTngo3ku84yCcztiNNacDep
PeNky9pYtpcUXiP5nVbBT+iYoUYHbRjjNFtsPe8wQEeRen5erwW50jvlWyFNJto4
PeByjgL+NS8F9Gk2a09EUWIENnqHBTmSDH2X3PnODmr5JmR/jjdzy6TxIGuc3j0v
FwsiDXFUS7ZFmBw65wDrSifG8bG/25XpAEjcNMhqqqB843h9nR+gaeCLeBlDy8RT
VxtUVSpBzQHgvEGgKPSwbMGdWrvizc/ANXPsX9FsgqG5dMtgwJqRLEQVVcfESbGp
yHCBOjbYLDRc7FhLd0ZyAfRaig4tRHGyR9UsA5fdhLTNwK6VsMVpe/NH0oUw2TuI
FsOkixQiRlayIuZvT/CkyStVYPT+G4SjOnyOXMcHZXAJOasYRqWha2x3ISGi5JJL
uCq4PpKPf3Kzb0whvtRGGLJZw3ujd14Ww/7rVYk9QV8HrFYdc5oEfd4LZausd5Ti
9YA9GdnTaxBKGDwFtSnRL65ZtNelP9/tVggBxBhGUlxDaCNoYzocR0/VE8JtaH3Y
Uhi9jNYiyIpRfFX+SDFgRIvy/46INO2RVq6f+YXiEsAebjvyx9xJ1jlUy2VrS3sb
qWXf3J2DifH5aRXCA+NVKp8BCFPXgV1LsD034i/zVT+Xn+otdpIhF2dSAH2qLwnA
khJ8CM66qbY6nUriA1wWEaRADmbg2I1DdDefSlXVlo0JMV0TWD3Cz6vG5MJ9uvCP
0YWb9PLmKW4P25OeH0ENqKfI4vMuF9682aovHhI+HvOafpKc4S/CjXMJdkvtUwyZ
3LsNjRzoL2lr1SyTCKA60fpE5BoN0bG4hcN0ZxXFIh53oxLFySCcmOf6vhqCV+S4
Rakk6LzY7Qyr0e6I1RLJtfyxpeLrpyJRVbTvyBoL0dNqFQyvjxuYRmvuF6Qkmi7z
mEzuf61h4S8EBuINtWlrEpsBwDQ9obCneZjfgcv3/wM6bFh1eaBMpoIoR+0JrE0B
RHyWj6IgHMRjaT8MLg21cm2ZVP4KzQNMrNVR8SRY3sZ63O57Q2PfUxxLnf38Bm+B
PkNGt8XwVjYpuWNfZ10+HlZLEG3FBc/RaRIFWLaCbSCI2e0qxGPcQV7TNZGVq+yL
kcX4a8K/Hccp5vVO9m1QXSFCs8kNLvqS8W+wJHbESISUR6g5q/uzILaShVTTcvRa
kT0yIaSc+PnHuY2kvq6O/+eS77HTtsdNZP85jESxdww7F7EI7kDaOcZx13I0LFp8
QCu7ji/72gtiq7DU542SAw5uREF8NcbPzNjLUmZ7Pd0K7Haw0zcPrcmBWgpZOKMj
avfbbuaNRXDlHTpwo8sG5aBufPXcu9GgI/Fc7QlU5MPtjbUA4YQfcIVvXs/1dtwO
aIlT7KW8M/iJrmea7qjhDzW9tFsjxTajzpNcimKXSinjpYnjMaQreS1omzwr2VYe
dy2mTxzobNGcA540bx+jCKa3Ywt70vlkJCCg993s6eZfv7xkc2rtuBbeuQi6a1Yr
sDUK6R1GsdOmO2gSei0QyX664qOUcf5ne2ImzcyxJ6UDtQltXRarNOOAzSc/sNfu
sYz2RQvmUglA4BmjnJm0AzWdAPVkBNun7iK7cmKP7XYq7zG5domSxC1qtB94Ihqg
pWTvxl0uVabxWo483ss+ZE4dHFZU0zCQRd7XQYAS9W84kyY1Lxc55wvhWLcdTGat
IB/CnoUkGUr5eiEtG6L/pzme4AKeS/aCo5ZjhiUKM3oYC9Z0jUpUI5JEyJRztvJb
qSID7dqVWsq3fZP2xY88eXcOiXR0e9BOGEtoOuISi36MbGV3l1uJWhN1V3VMEDt7
hR/gKviUw3bd4qJNNM2WUkrB2gNFW3TRPcmOyUSGJoHTwsxGR08ednm9QMwkj5Tj
H4JfRK0yfkSwnM7Gz8xT5i9EPy2AwOUelDf7xyEQXPgmJEFvWDVN3/GEEhCQbpSL
3Fut/unFw4u+EPFHp/Aw+myoIPpESQQZRRRX/pne7C0C9NodwmWI3Oe458SRjWJ7
NaF5dC22JJx7V44WN/xrl9gUKL9ZbC/n96q8gvS3BNmWiFUUek+oCv9nD+FV1vIe
Guc4QLeoMQM83Dbljbb8k7ZFbE2pypYLwIdIm8c/Ls/R+cHVpmK+JSHzUnFCrLya
NRY7hXA8Xl0tJapWDXhsfzlZa0ERqoKkJSPVkhi4aDhsSPjHMsRD0nHgxb/8TEs6
t4zPZLKfeXSEF0Nhq5N3RybgS+wEVU7MJZAE9z5R0PjUyu+TIaE/GjKLqqSkmav9
Y+m4SFCHpxsUfyVWDdmvrFbYwe2lgiArD5B+sX+y8nImRIv/0Ki5+yddfUb9J1l+
h7phRBl2WgJdHhppkj+5stAP8Q+E44tScJmliHNc6AhmezVXBGtFkU0z/N4yskWe
Feo9N19jFfEOa1wC+/JructnwPMXJQUDdDG5Ucr9o9+VGv8y5i6SNPt1E67Yt+lx
rM2f2lqjwdGr8u8HQ9Ovig0q7w97Q/mJmPFSKZMRu2xQY1ivPQRFTMENWIBwM7Fj
82x3vSEWRd3GnBiFNMQ1qrEq/0dvd6nbhxf+YbiXTtmuoRnECG3y+PH/N1WyDSD9
2Z37sx63xmkG7NcGCwwlDX3q/ySPgF2fuNAihziEtqQPO+gSO+PiGNqQOG8u+kZB
Jdo+1ZE1DC/iUh5NCw7nOhWab0dxEkAq11rehVUE0mMm4Pjp/ikQBEXlkunIBLWL
28YpNtE4KycwkEQmETCfU6z9t9dpCUQDfSQZClDpv78MFUaZbQejNSUARmVy50lo
1hrDQEMQa3i7QxwB8/k5TG99i/hlh9Hvb9os+fGgxm+9Ml7gS9U5QyUMLj7t5uJC
cbXuQxZDuD+0bSDaySVweHGdgG00a4tvHdWww7MbHiOUf30oZdq0rc7fYMDx6Jzy
OKFqBb+3PyAIqEK22XsCjQN9FOBqLGFNcsI4d6OEAZF2gH5sMJwpGfHeHnVzYOBt
Fa4z/yBB+qnecsjkO0KWIgmMdtl/ysn2+LcxWYMeJXbbpTtfClXIOuXJsjDp2adG
IqLeh5FyJqitESbwlYW21L/fnTZlUy0NHGA9cr0lGDa5TmE1RnnzKLRWjI29tclw
fnPg0jF+EfKtRH4b/uPxYUGosJ4Ec4et4MoM+hEiJWzzHA49mzLBVCJxcYQjApEq
fX5qSwkan4qUhMUi3ATWC1H7QeKMVoUZMqjG/a2Y3nO8RqA6UT2BTTPzNLtFeueY
t6tsS+27e+KfD5aUPnezBFDDhWo1qFnsFqOR/lbm7BwUtUf2g3mMOr98rm0D30TS
5VkR4+ed6pX+rNr/52wA9KcL4PXRHG8rH8UeHJSh9xNi/Ez/GCxoOSKj1O/4383m
OLHXCrLBY8byxk+C7MdMqCr2vN2oI+je2DVFgxADrY0DeO0ipQQ4tBoxkDstUmnC
ZMUQVcb5cVT54xxmE8SAy7WBv7SEeg/wXRzABGUVK6O1lpYchJs2AF3HbPsSmvM8
wvUq+Le/1CPtgoqA2tOuqoP9G6yEbPgTP/DiJAxFxQueUznugrYG8evsUK5gXMYF
fDhQ68Hn2HfDfLyFN1inXMZXk4PtnYB77wnR8QXMMIKA774Cuk3CtoU/m9Hfz/RO
ar9V3DGLrJo2L9ZbK1BUeQVRoV8ztMzGUqEpCbX14q6vqWEoWLMfJ1clCaqOc6Z3
7stV+zbGPEWRJ2WiZ6wwiyyjHglJFgL3nnbnJHzT8zDA2qTXsM4/LXzvf4tLLdwc
7BjQd00db/tBYZU3JghO0jyOZ6WhYTNM30Dn6Nr6m6G3yBqMB9bd2PuxP0ib7Lri
6g5Rsb36oXoDmSl3IW6ibLmGJSzAB3AfPG53CCxlWREj7liHJ8HT26xaUkW721Hs
mq6+B15NYlzCeGGiBFMzJFnykJu5liRz3toXBq07LBfbWmuGd7SRtCL5cySGrkBa
gBhDXOdXjzHEtHvL1/1jY4lUJwmZnTjq0+OeKOCTj0I7+gGm/gveakO8FST1jbaP
Szi/T7myobJlbPjdHLe///det662nwsOYf5o+Ziy5zEwb9uBaXn0gnZUyk8LAJ0l
TZ2rwcVtY6HaC9rAh8rDxt89DHgklwC0hxkWO5A0q38+uakjNEKyadfyDujggLbV
vgXA6h5WhY1HvjGd61pc2mFotvqNnftOY95fXoJR2Vi4fNXFe2mcgQy8vle3ttKi
d+tNuvSj46T8oAqjC8XTV2sOOtkHkkvKKvydDBcD4YpueQ7EM0Be4mBsIOYKi/L5
72uobgUxWT7I6/GZfDvBAj2E0MUVAS+J6DZzSrrOYU/kiJIVRS3EMpPxwfj8DGJY
2zrEcDAszFPd1G637UhHfo+Z9gOYklTfZzq27S5UKO91WtMFJvEtV2oN38w3ADqu
xI49V7LuIRTzOtXQp9QtOfFGPxF9cE0UWEarImkVyqtEmsbNn6gUb4uHhr8JMJOv
lytPeqM9XMmVxI6wQ0IVImhW7r2Uc2Vw4NzGat8vO2egFeQ81JhyGEqqkLaXvVOw
Hgv5hrjg26vmPR1qM8llORdTg3UuwwuAmvf1WIH4fOsNv1j9qt7v60EeH/tH/Rrd
5dPRMNACgNeXL0uMbGDOmgQL/QCHKg5GiAZ+2tdPZKWkwLmJlb7JkzTW9YHRz4Uz
n98qiGEGw26fRXzp8SYBBzSu2CMZ0vPlk91/JNnibibVcaTkSUgCVoXQzVwSaSpL
3U9fdZIWhnsFQV8jMjV4JWvDHQn32Qc5Bku34gn3z8UGrMxZcD2T2JPuEn+TYDEr
Zac2v7o+MQQmvVeDmMc5BayBdxzsSXgbJphMOO0DmNCGs8iOxy7jIGvdq5OWa6Rd
bRIASRCUXZa+C2mZpTpYZHATpLslodIoKQBrsz4+XBAwYe5mIchnwA1pJfHI0AK1
89jOPoI7lGCLPNYXNUw9Ex3qMvAIDtIMQ6lDj2jdt55PBlAXyTAiEDDxgSP84Utb
ElE9O45EpdnAfqmMNfURd5UxW4LJcfHa+EkZpTl2VE0HLt7FVIwbwhEeP89Ykuc+
RDGWbKqRL0pLCItsYy64fIOWpnjXSqv5mDePSmL72BrVHQAG+V1Fnw5T2HlBE4E+
cng/me5cUEjVjlQxV+C5wArMQZPd0hoHQzx5akrqJzNIJUeYIk6jKa2hBHwYgkoO
MJHbTm+beEFDTfaGIrsu+jU8ggpug792urn32HJIZAtws8+U/WZgm+2dtuFwtHNc
Us+jG3DJOmATSPVeil4z1XSrQiNIsi1Vj2/GltWpXcJsaw/9INPTB8rkmIeebT1e
dJTqblFOZ2H7AJfAiXH4wgAV4lQ+4nc7U8rA8bFa1eIBX/8SiVA3RJdwTCY+P3AH
W6D4Gb2poxYrUcx0tWHjztM9mMt9knFqrMVy8Lswgxv0VbcQSwe3DuVsiZ/+T2EP
0L4+h7xVSXHJ/3tI9CQ0O73DKxPN7ssgP9RfNEtqXD20Q2tSb82NJacByvV66Frw
0us6X7fPFujhDiLdaco4UyPVUP9le2bPapF4nn9amiqNB9UJqAakyQKbh+gR/+Oc
AXC146etaFP1CNocVMDp5k5t3xrXrTwlxM70Zq/6WASWY/bPxZEEhaU1d2vqqLo4
KnlqtGarO6CTDJ51XCZYLQE67Aed7KWQIXaKZzHbdgbWh3Mj0Bf75ZFVCM3Rge1t
Yo+MD4xR707iA2lCGIqq/VM1MoyoayYmoYUCPc2eTwcereiFJodtJcea0FT6y9Uk
H5ZxCdp8aG+TDMh/R1e9bfyZPDdGogRmo1bZTgfrpdBFNywc3G+BY4OHY7sqIRmn
c2Mt4+WMAiL43o1/GakOayE/GH2A8Z97CEguOJwi1fcgLXdskQEazVvrnx3YJCku
fjqdDAF2sbv8SgtGtmOBZTNo8r8AcKo9RcK+Q/qB/P1XFsyefje4O1FIRaDbktJu
bsK6Xla5Mp5sWuldzEZ8tGH3jpKFNq9b1Nt0x4MDPasOeobEJWr/mH2dSM2mXETu
/0zAGP7JEKphC4BX6pf0G6PmU2gbIYzNMMc8WI+U0zqO69p1RP5HcEt5dJhBffl7
s1Ak2SMgCxne8Q71MvjDUivirT44VqWlS4tumxQerxInNVbYrDCrUYOYLyvM9NPS
1yCabyJeTSa+4vCXUlmzvROh5wPmRWmYO71AviCkOtYyXI2LqL3JKdd5AGT2r8iI
gPz5uWuAxXtP6Rr0B+HkmwYvlE18jiTARc/UNo5xgMkRk67q/FJbV6t805j9uZgc
u15YgsXXsow37rIAaxVE1X4MMl0S2XH3BcHVwMpSb7lM8e/ko5w081Jjov2VtAC8
knnhJt90Pi152icPM7HhrxQB0x5+ODjl6RTYFGkUzhZrndwDm8h+cxhRg51GwX2f
u9fGKSS/ZicBYjeWIBoRnGXUl15cobQ9Lh1hDOPZZtIj8NwqaYJHv9Lmm3XANcQH
+AqcSHNkh7NzWrWG6h6UgJg3NpWbcewf7tDeYgAxPVHCxkkVqQhhXZdr5gWkvk0X
T4b/VN0D73G8B59W+syDo0B5Ydk6wVbOgJZ2yIz6ry31DpJV9S4tSBf8YlouP7+w
PUV31Ys6rrAYfr/WpwAt5u2J9AdG4BDd6JSeyK1BTYYT0ND0DEZaxPbMUeCN0HlK
QGAClMMn4TPNL8QfIRqfnB1tlv48ztAtVGD6F271fSR8dTRIGqDAJgLwheIk+GAK
guorwmdUXQKQY8EV+ACHn26A4WK7N3BKq8/9JVT6ZldkX3bNTr56VD4R9aerXbqr
+dRVSsAHBflUW0rqq5LKAx9cFxjpSWDc1kssE1tu8xxFmu1EdKamWXmHoxhAPULc
nPC4A+AS7/TNr9gxDq86nxuS46SNQIeVCyNTGKkbaRDQAZM017a5wzgFMiJaDKlS
qTxNnistOuPZUKqh6cSlVeQaJpG9AxkvHvW6kieo7salXWCXc5HG9HPuhfssDuIZ
K/m/EjR6cCubAkmHj8xktrILQ/axNxHmP4pzVTumv3UyNWWvkQxPP59WsqDxAhfF
gkpgMQAcCrfmCeirSYM4xXo7bqpEnS+ih9/UjGzr+cyhWVfnoTQXDZ7VCnN/uOQ+
f9Hu/5LUxtJlFa+9ej/ZvlNNddwFIzdXcfYnxhJPNGKztkLmvuR+1wN1L+TLIFBm
rjIMsWxovlq6NH1TE7mmr99gFzlmT3kMAxs9m14lU1igZ5cCf/Yz0fC4S/J8ouKc
g4UHUR5MOqqTr6R8yLlBTP1RtnjpGmPTH0jsSygeMYJ4LTJso9prYjqayxIPY9Ha
JM2WS6GV83ghDdqtUdZ0gvPtOv8qZ8HQGtGyAOABT6Nh0qnotEYKdWMtXI7CvDhN
eeccRfkIie8BbeSM44vtL/6dXRQXB64EKzEUCq0KNm9iSbtcva+QCKIOxWu96gON
cwTCZ+hrVc4GIVpysDYeqJP/lddnj3H3ap/B40EM/ftC5YEIOYlUiJvubdMzC5aS
sKmOz/+tNQ+Ub+X0q13NieX3ZjtZ+O9/b7usPG/C1UFtqkypviytb6VOg1HdrBfX
zWV1jTvPQcyzQ2G/UuBjsl6aqac0V8FBLHelRjv1BfvZDRDy56/3v90jY9vLoc1W
Jg7UN37nbSq+Tx4rn4TgvRxeuJbi7deen3pemLSfIxGjJK6AdbhoV0aWvvlYlveF
K7srdm9EAg7ECG83wnPdeAMkFvjPFzRKs6DZURIxHkmuHlHeMAK4HLynvSxdEuNi
l3s8yKlMSeCP6SRZ+4r6g7tqn4fjb6JqxfklrE+Mgqv5i++9jygptjIVphWYnSuA
O0gh/qSw6suQ2Uf5b/nOqyzHwwo1esudxHIxtB1cvlOv2LWjaKumHyD3DgVVl4rG
iqOjyRUSzz+38W1ZkhYPt5GSVPlwwNg24CxpcOB5iBTMMe5eOPEeJlrmDX4dnvIh
E2dEG0zSn68fkxpxLB31KxuMKJQUi6vfbUfo+REM4vv7R9zB7oECzg2Ufnj03GNH
cPkvE8I3w/0SdbqKRek98s51kHD9umP0mHKfv+DsnvaiBmwjsanwarFpx4e/5cLi
f/qe63MoGW5+6dVcFuQpn4iV6wzxz06s08guo1tQH1BxE/dwTYVKsx+nQV9eYkRU
yoV1kj0CXr8zxAuHlzpKTq65vaaE3K0UOKJiHZtvq3LnmXGJ93GI3LY1lawVZarb
RXPJrUzZeMhf15/QqA7DbQX+tiiEF6QQMH41cjcNy3pZxXMuAwgODmTRGE0LLlny
4dlZXjHVl5qhKJ8fXMqOxHzg6rPyl+Bf95HGJk/pVWB+RQCF8bhoMKVTQBByz3B2
DRfrcWbC4m7xrS6916ozVf2MqxaOirJmcuKvoFh7Mw7B3A57kYCCa4B6KVtG6Ndi
EOvZQffjjcT1BKCK01b156O/o7/eat7fommGakCNNX/2ZJ5oRg5BxQguSmpr5ljB
OqvwwcDXIHKyv47A477bkgb2F4X8hYXqsiVPmrV09KHPfxD1ye3gZneefDFztfjW
M1bSs5y+9sRw4NgexS+ARcKtNsKM6anC4gRzW/Ukxw6+kxDZIJp9dQoyBiS+ze6R
6sGWVPn/alKLBulNK2lRNeqMOyf9jx5GtFdLvJuPUwUnsbV2s9UUtQvRqeMaDHso
/63Qwvs+8dM658vlRfQV94JO6iGJf1iENjWmZZz7wEUp0iyYIiNplx7/TcAUOvIo
Onmisws+X7tw7CPjrZPJ/bf+IhXt5eFCQk0wqsIVx86BoSyvZaKitY3OjU4399Lw
3ya+xbm166495Wvd7Z5gQREwd+AejC4UfmloU7i6FePLOZGW2gTJekl+8VBkOZ4f
p6qgAADQmenKeSIsYPx8+D3QxU/bQWb04hcx2rBIYUTeC2JvSq8nBpB5ULf/8anh
NRC7w2xypoop7LEUedxBcOBNzq6T0XesnBgC4XivsgQbsDpVUrL6lDOQ8AmD5Ss2
cx6dZAnDvlo1gKF8onzde+GAVjxvy/w7AFRXaoWf7dNx0jtGU+fidgLOSqWnqaen
iaqKIqFjzneeHEIA5MCJ8fB8uZ36hKVI5584ETZkW9Vp/u4ze42vT8gu99sx8cWO
S8BAedXI6oZ7ctVEVqNxCTa7xWu1cQVUDGWQaVGe8/S1xTUOAIPIH7KkE7QWTHct
Ip6mdml/trFi0ACZlNU+bjccSQ+UJGlShYlZrxxB/5miTnPxmuPmSFkds/HARbTm
5IMktYL0eLtMzx/Kv2Lz7gHaFHFHY5DJhzBJcHC3TNJOyx8TaBtKEOLBheudD2iz
2fsFKoze8JtR9EP6236ohyFkyY6uRQH7XjC43qQ3gUUHwgAIGbZwIcnPmyynMf+r
n2vdmwaFfPVHxeb3aD9OKp1Qt5HYfbPpF11tdIobcfxaF3yp0tKNnOpmQdbpQsr4
YnKSol2hhXpZJoKCUyedMG3xlGedm1O17vaFBErqphhWwqWw0BYGScw4vZTt2xFn
eIXRKr5VvdgdoEdPeXtN9jImWvaVl+a6iMCSr/RWotvhks8Edr46NjvRrZ6G2K71
PQ68pD1nGXsQSAR77SFgVNP4hsr+43nyoXw6zMK/VAOyb9LYIjdMEYWUtlR++zG5
uXyuiALmJTx5yVTzN3fAxN/hL2GLTJlq+kWetLKor9TCrM55RLQZ5eGKRyeqsTIs
ZsYk/swwRIUwZYR/E2UICPoV5s6DwL3U8DUXXAgajjd+ps186nlAr7rV6BlkISi+
dkqsXyOt+jI3ISPeuVH7Ahb0xiAoDk+/qE63JBShcND6qoiDGDM/lS8o4az/QWqj
WMA0LvXvpgMaQNeqWLvbTTiCHfVNbkfiADW5BemDUxFy3q4gJJjpSwPMBeI1bMnp
t8r7SQfiTepOReglmeJ4nLOPls+9XmHfQT3Ka4O0V6wBizXvUJWRjUIeGdCPOacB
y1H57urgmuovnMiZzZxt3UuFaBeKAib+kimWNwrhShDwtlBxKaRmzuEAdthwEkN0
i1U+3XSEQ130fr/oof5DX2FeFpcM9otE/7TRcoyfyRO7UiqvEeOKoHrqkJJr+5WW
2aUhvGA2HmBZiTvvMl9pjLYgLVd8pZM/pr+vnHwuL3ZmS8bCQhnz7tIvElDIK+ED
ThgadJoxPoVIekspskO1UqHVQyG2FoIc4xPPklPg98XkneIWOyuDx0UQgaclfVxe
XnQ+g2JCMjCEfTFoEhf5WS6PhMuiLE1r6s6GhRSkWtBxUrC92LJGnHydb3PoPHKn
CrEuXFJ9vCw8MGxAp1PxkLRcph5WfzT9QZxBlgJbEIa0nKVtGL6gxgPqin26P1BJ
COf4EmDnuo/9JLHBqbU4mgHDb0yZSwcR5rHAmfV6wJTMLED4tlW1YRkbIiVJyzlM
h6zhXykSNjwEXZFfr6e+s0iPAsIEYb75j6nLcZSOIqb93joozqBeIJmFGowrVxyf
1wyKsQm1291u6JpYBWTtFSXKOvMgaCv+0QoKCZG7FOZsV5T8lIm9+DVjFD6kx4eH
0pjxMtQ4TquWbyXQF+cuMo9/tI3iZnYzdfOVcDyi+63WBPFU+pcDM5iw6LKgF5Ev
Lnagt0bl96sKv7cYXxMW+ccp3eqwz+8xqLLA488lOAYElIYELvtpEX+zbQ85RoYu
EqBQwqwlE5GQvjEzgV569mnYFiDqdGzGb9UanV6lI+Zj+QvuUqPVzPnv69YNycd3
PhrKf/+HABYdhFoQeI2NU7HyRnkaRuTcZ3KQRs/q2FES5YJUWNM0rnFKe/DyOIfJ
f7l6AWXGvSQB3jBM2pfbbaD6IZSp7Esz/rUEN5N2BWyew/9x+gptQgYNumnIdZAw
Nf3JMHe99Vpudo7lvlSGv31pEaZElWg/jvYNGhcPGgLW4/L6JZ+w59BJpJulg5o5
38eI4IaB3wlNgESTgh0odJBqODNTa2hn8wBBEy6BeGJiHW6z6gXBOnlmHDQubNw1
4ZmOiaihmIPQ8WakLe924rwRyBAi4h5SvhG5jAyBKZrdnt8/fS5CpQPz0ox1V5P3
YQLQ7mPdgfObDrxgl7fVhVOx99sBfo+MvU5X7/v8deXlGRtt8iIvScI+cQF5TzJ9
8sSDEZk3CpIfYS9p4HPnLqAqfiVNvNQH+M9ll9bQSGMxJfZl6C0zeizjHvsaYY/M
vytk3xzQa9Nc7KpaVfl6y0P4nMFe2dse8hvoPvM4HH6erVIpda5GMhpCsKFS+c0J
/dY3HzoZMyffMpmHkAQ5HGjjDlGi9ZNpsmHAOSy2gdsmVmh/d5AtSHv+Qca3YJ8b
4BFqZCVcA+2nhMFrjEUTZEWrLqF2HPt+fZC/oJwJVFneF7Ox1p/63EzkNA8k0z4d
FPoXGKbvSvZAFPvu2aEGAsFVlvWsE++DNvIblbwHCZGYBoH3SFOMUrivYXP20W3W
t1mIBQxrWfoF+RxnphkXmGjvKNfrGXKNuTZyTeiq/8mHpQS3c3KGRkUwgKnqoxvf
Z6EQPGik1c+seorUzz0gx3EhX5zhzZ+VUy+iKtEMa6yG3kh0MnQx//B8+X8GWlB1
Ak3P7zBOvggflgA0ynfz8nPLrycePhbgXLDvFDGEPOwF0Mj2PK3T4BsP2WYAT6UF
drK60BS/6H4eb+6ZO/7+8ucnmBlPi+2NPlH/zNs27u8NtIoH/jDPwA7wWe9AX7ir
9zAUcoyxcc8F0q3tVqWhjYJ84skAZ31tk75FOjmO/1IkOWYUb2QukmoIfYiN8Qj6
5r4eERArljIhoG+0/65PfG1WIbcnn+tXUTGmGMJdB1TZlzf0CyVpMijnSgbud0gT
YJSlGk/24+zzCdDtMsgWEHVJZ64zF7WlnKX0ECg3iMcmRqOyHhkc37rVQjkxsMLW
yIFtdz+MKg8CWuVEpcwODlaiDAv4xarDjc6whZ+s7SWQ9+7jw2Pe4bmfEZ9W2+kP
4e9WJp0d2Ij2R4oW74YeEx2MaJMdH9rrgFGVzLmU2YTVUUISMG23go+R5KAYiV0G
uur4dgYtrXI+SbBm79SgsVxZIMdBRyxwRS0V4b6V+Ef2dhgf7YNp62HQYccip0mc
tCngHzG8QCayywNO9WGJX5axfDwHoVHJvUNkJQ9EX0nozlXDmYeR4UBCn1x5F8tu
ifZiaEP3/fSRTFISWDvD6txfT/Z3xV1MMZZ6zqufs04KgU8jFqKdY36iowL1IytT
qCzWix2lbbdOZ62MVUhsl6KdfhFXz+5ekCli2RpCri1dJBQhFFvwy19oLncr2SjO
TVxFSM6hIBIiVBczwPUHG+TJMpKzElBrJTHyHf0MIh9K57KODK665aFJ9VRkXLuc
3rwtHPJWi8RuKtfFlePb/f/bzD8AUpOm9ULUN8LSf3tJBQOz8GBFbbn7cr6BbPjw
Pjtm11ZfRP/mAaTqaHrKtpEsJPLvO0d/oyaXBdm4LAgmjpvhUr2Mz7QJ75o0NB4f
19xq6FqrZPA/kCqFhKk7khzs3LVsmxXbA6jqpRYwRi/0MtU+Cn7nSh19vDBSyCN1
yDJ4OFOM1pcPXFbfsVwiCUAzgSJyAM3luN2oN1WujVnfD8DCsfpRANKiZNGLbcli
0xClsC16NfqIGuNN2h1PjkjM2gjrlA8bMWrkwX5J0ZDEdJqx6t4zCaqIsvJ4CX89
yOw0vpY1i0BzZqboUl1rsEtj3/T55s5akdXSt1MVAYXYKKyXQvpL1JbMnSIhkMRS
Mg3ZjBiATy/5T0KB2uJ675q+MofzeSZPOrNMHBFotbZGmWWcz2sceSAcmab+naPD
R1Mu6o0X+F8/8TPD3C/G01xnSrvY6brUQRzzfpnU/Hk1l/i+eDA9+jITvNZoKCU6
0wQL5hzKgWimeTV0Su8Qrz2WvZvtMAkP2wCNTAr+vDecK4JtElKm4MyKzj9CIoDS
Sn/IYUhtsURK+SSop4Kf6qWpeU2PyyzL+iH2siomR07CS8Arje/zd1pkX0A0u2Nq
gWBx5SP7kaWCdt9NWTdD26JKu9d1V2DbVzg6FHiNWtMKrPcH5w4hKBld8J0D1m8t
QqrXrjqzS5gz3zAtTs13Fm7xZrn9cXCO209WXr4hkEbFLW3P3BI5bb0riOAq2v4h
vElMOoCnszGneGZ64TNZAgNAmjUwZV7CVfzCdWXvm4vUlNKZgpCc7LED63lK2m0F
6BvaFFiyDUyELHZHmOAKNz6iE7VzrVEYha7Ji7Xq1pTgX22fwFQ/aKSkxi7Ua5ON
R5/5BYO7vbodhb+taosEae1IQaKZLb5Ey8+eQkrevHADDFbqymt3fEmNnj/mInbR
G3UHGFhO+x9Ut09WZddQvOz4tnWOJNZAVTM0PRbY0qqC5YcimJxxUH2AN52JmVNS
luUZiL0cuFIzt4EuI3+jT5+mcf/2l1NV/BImi3FlDrUp7XNk0g8Fdj8RhEkw29MO
UapMLYbNu3ZuJmqHpBiwEwU7j07AdZgh6U2T3tA4ofy74OfXboEAhlPuVYCGfSto
Lw9BknwpUcrTM9au6CTlOSEwjggrdCO2v/jYlGVphUViTj2CLwI6p8+3IIKA2EFM
U2lCp5YNO5GD6KesvDEux9GonCMY+83BIPcqYyTMgItoCrlmSQndHLZBN9OZbZQU
uvFrJ5T7occHnKwHX9J30wN8PlUgH2pik17AF6GcxzJQyS6EshHeg3rbRYbcJmaU
BHlWiujRF0/AOXPSFoXMPWe9KnHLahvPV4ykjzU497uqMhw6a+ZwmCUAKypkcT4X
2a/sWm6qAWWdB05Nj8/fajy1OI4aJ9T8WS0l4O46KP2gZD3eBTdqvRGjI39EAxJq
htJanujknOMeSrSFGE1POsiUDFSHGqX49TfUd4zVhzCDtjlfQRrc/O/bUJPLZU5w
LYbTfZ6npZcK7rm22NtSeO0tss5jkDtpe9KWi321+KMZv6Op3aYOSw8vKpWxhpZa
YR4U+TRgQ7gMUKweHXYOMQKAH/Ncu5EFUy7kfdvYPh83YiZbypRr8GKAeAzc1npF
B7KN1wrzG9+a3pQhqUHhRyT1fjliUb6TLY0QxhvE5/MXH/88aQljaFgkGb2TQx60
tCvmP6Yd+VDctbSu+iSUDuV51N4wQ+Zpe+dgjdN+VGuErIIdBlDIX7HpEwFpVHEX
XzfKcBl8JEMK7yGVxeHx5rZDBPLDlX4bysuZdgefsoWlDlTdzcm1TQJOsanombQl
WHdFvVjdsOBfjS6SIjymZt8nGOIcJq0UyRvdj5NEvZklv3W4A6OCv/kvOyrcCW+A
MnJSnKTslUWR5rqtJhp00uQ9cXYVsFRh66NWVRtTNVNt6zPaqqALV4Lp5+12Lb37
mob6DVwLhLxVXwI5HpU9a5VpunyzTXbhdQuQL2Xp9rGYno0cH/YwPjrfCzzgURMy
ZAOzLznlybsujut0akrunWMk/xw9Lv+xMXyQrDWcZVnlZOx7RcksT0RpyEAOCM9u
VVbHYAVv2+6lW2zAJHzKKOTgpe3Iwe3+E1MpexK4n9khyhl0793qHHoeWZHxFv2w
vNPA3Ya2TYchLQ4tb+MdX+CX+PyXpoEOUB0zO4p6w+E+1fFeqN870qSRK/3m++11
hqH1vRkQnk7Sr2g5HWpiprdX9Zw1yQxJN2SM2hEOiWCi46RTg9elAenf5WfwFYcq
bLEELL2Ld593ZcqGqlB2Fy3zcpU5Zt+xxmEHxEgUC4kj1MwscmxxTey4YjL9Dbs6
kcfuWYmGNFuGKDYifYmewRsnBheqy6BLkqHyCaiKMitZLnjXDLBetOTqjv1wZqpX
4aJgNejA54Tu3anT5YoXUOjyAa68sYg24difbx/HnnHHWRJkPc71p49xFnduuIqN
EVmasriHshyBgOY5R78Scn2QoXvmFkEt0sdu5kFXcsxJSjD2Muvz7jtzVzossTZP
A1gZ7vcdk+uaR3YP3d833qbRoHQcsjkbXh0Dhfie74kohZbFZZMuSqa31S9dXm9b
nyZtNvypBBMTGf2H+ZYeF7+6mBvopT4dpmOC4rUhG0zHwKeBc1TTzWJQQnqki14j
fvfcZixzSEOSdE2+uzfaU5s6hZhdk9FJAZuw/0zpgdM9CO/McIl1ndmBNS0wqBvI
0lcmODq9b/uLUmi39pM9KY5t5TrvoyrUM1mBzETowFGKLQIid5kfpgYF5iYfzoOA
koZ9d1rBOj9JY/1m2qkRl0KeCpzftF2eZFjpb8iUtloABc76pcjCIbZyjIJVXTCx
8Z6mt2KDvv3C4qFtnStIamVpQVCkUfQ/zjwf5b+edtcWHAp4qusxuzXTqKzwL2tm
pEIl7XlU/raoAQPy3HV2mnUSOU0NpdcRl0WKm+6NjKjrevzQRG812VjX6GPPmZYJ
wq6og2TVsURweOmDp0q36mfkrWudtH417VX0ZrA0oUa5MAdOmquhvoAGc2H9CvQO
pn8gTVNGgSFf286doYuzUkItbDeeuqvaDfdV1oHDg4fyoRWOmsy4/cxU3TUeXT6u
WL50f47GqS+MmdKwB7b5qQrXW2yWDP4ylvdGNBuX64I5L6oufDU5guq/qMg8eNp8
iYSf2pTA9io3g020G/BlKm3RR/Kl2Hhoi7l06p05hALzC6LLG+zJxS/5hdpWzNLF
VLd7IUtf09n9QpFcBlbToCewp+7+Zyz3gDGhuOOviMI7YiC3HHzrwMpqikkc+vv0
qPdvf3Z0RMgsMw5+SmYYJvJw/bo6ukDJpbHSobyjl0E6LSOtCswB93t4XP545Xgf
QepvEceGqRfKCCyTsEpnAlaoAZnzOc5bWW/a279K/E/djRQTX0Dj43Eik5CwTZEt
TO3F35+lun6Ea/LvT1LjE8PF7xVHmsmB94a8Ktf4JlcpaArM4k/EXJ36oHiXM9cf
QKjxCWjoSV2KQJgASXwtEy5WBRl8HT6mIL7AC4gADkt4axz4U+M7RkQdh/IeJhPv
Z9Gg2FR7JDETWcACoW4ahCrBEYFy81xtost6yIg+xA9OMuEi8nQ5XOiLBM90eK5B
zyrx495EQfoK5Xah/GKSbtwTJLRIwX0Zl6K7HVv/XbC+dzybMOqvEljKdEJ4JgiC
adih3hRJM9BYtBV2VXOk1/e8QpGSHlP41tOE+n/VogH8GwsUQZK+AL6N7dWeoPtg
czS/b9ivw1wb/jMgn8ZRo3nZmn8OzTfjPKrrcLz0XTijpN4mgzO4jTTcFTKLzSNu
iDZtRH26185sMhJst2fSu76fxmY2Klo8B7ztldz5Fa+BtGzzlmM6R02E8obm9Vqj
fV+PEOUTMgNQVB9PJrqpN+uKXykKGyeLIqNtqY/ONH1xDZQAJgvfw/y34OmdpBat
kTFolVgfQ451q33G+CLb1Q+wZ/7SWwHudVge3cgQFq9Sq+qYf3l4FUipR3SHSNRI
cEDCHZkA0lu0T9UA9m+lZP5l3f5cwFJbWPmD4sMWSuAeTe10IMmDDCBuXZ0lxpe4
ZIygkAPEfWNoXG15TNawnKZgg+TIKsnGN8DOpIFMlgkt2/u0/UrQPJ2lGL22nxNR
lziDG3KUVVjq5qB2V7RTtQDGLkRRogAoMKkAMODm4URA9OxHyX7tywTQqhmHvjV0
10hbxKuvlKhcENfi5Sae3L33OX/c+VeBKiLIYPLjkBJ8/grUWTe2ZBXCC6/tFDnq
Y4pSk1uu0PlxzbrLPZrC+yQ6yHuWxKtCXt8G9cvEb3JnJQsiakBsQulBx32qlXlU
SJ9kV3VuPYAhTW9nBjHhHTR4upbUt8Yjtak44DH4ezddh4jDJSHlJpdvr+RrhOS1
P8XKNoMBe4Qnl9N22Zmg9PY9e/WlXZpVwQip1rRJBSJ+R2XmnfzKb3EFR7fZ0UQa
8jSfeR4+oAKDxPjV2LvliKhm80k1AJwrFVD8fLrjeERTD6d3dhbVG+18QfQUQtm0
IcsXOiJEoocGxUSKz1Rm5LC9rZmLnXoidPOaDEhcpBu31kmvrYoDu/lTBDAtz3CQ
IAo2LG//qfE5ZhO9EIOwfBzH7+LMaxkH5W7Ayi378iciyXGg14Tzk9AH1mtkLVDm
aoij7H84hgZeEQvoekrMIiYdN8lw7J7cF+Gxo6Q5AAwYYipa3W+5jSnThaHFnwai
YTSghWqahVpKmMz/C0IDiDeGYKl57pcncx0AAmh2+U3fLql/r+V7WuAAA3eCZO7P
x959Zc9DTFcRh/NYY+i2EYW5sI+9cqkUujW7K0WdTL8wYQ4VNXvYeLsS8fwvD9yG
ZjHi+qNLVe52pw7QbvH+s+ZSI0cvCni6JGzTXF69KQijELoxWgJEuBtu+sdbro/H
DPHmeEVgsv49YHlF6BM2t0tDXRHbyQf1pS+bR/Rc3Sp/QZ2oFdYieXxFfTM2xfQ3
pS0LGCMjeeghwFEJdJclU0OYGBoci41Cbyp2qP4XaFxwYUPDcCnELBbG1vSkxIY2
+xAdVzGw/ITSfOdrTv4qHD24c3FKaFIWYkLkfIlLXqtF1GhznhXST1XYAYg1tLGR
ggZZ613Lmvg6/K8QEzYIHXejnmdXeYNwVkbp//CiKBseB+RXYnc0Njdl1OTdO77D
01e5XmcpO4J+TAApNG9JXACKyXr/TS1QYSIiXtnBIFGkT9YkpFxcTE0Tf5iI1c9+
70gdpQnYPLSXKgB0JL5HtAUA5+AU/heWwkUOhpVsLlKADAMJPpLVhS+XICWXWuFS
dp8Jor1A+5ifYzzyjnRUL1zpdYu4bCog1xgKhLb4NWwOsjSXCF7TkLLoQybaz3Vr
jwnKliUrS654qJXhhhSNFLJGG7Srv4KgBCRSxGS7orrrXBcCzH+fFtBYFPUvOZ9g
O3bjHMh5C/4Rk1fgPxCmMSBD8co+03+tTpb5437HhZ7o/yEfw7baPsBaXAeQikgG
XGmN9I7r9aC4E2I1tTezk9SzQhSfeXRMbJ4WYcQK8k+tJj61FtWDpy06u4raYgZW
kMy25OOuwiFCSm3ey51ErrxDqshxjmnpt31F9a2MGTW7Y94Qn+1qHcrKaBhKT6Kc
gseoIqIELM4V/Mjbr2bHkakfg/6rjo8zSNy3CJE9TWOVyps3D2ewfN0ku8XKMsXS
mR1fu2vkJPyClgw2zY0UHDIdal6MQKtL8rERZpdhYnennZItDM49K13l9zdQO5n1
pBxgBT5O5/cltw0a+wfEzhIdWzfI/KvUS9ZzlLCVl0HHMuJb67XdnUVec+cXLV0o
UDN3wTSKqxAzAtucaDA0gdyDBL8zizOIDMsvIfOpy+qec523SNXxBsJtPkToLwqA
pmfrRZhl0TGbDJI8/fe82BOpyJ3bQWQ4TiQdlQN8XZRR4Vzj7U18e2q8uyz7Lu3H
q+ylup+v2BRP/lIxEje1vz68AZ8YzlLs+fYKDF24Qg4hzEjHHShmqHk/YDi8XfiA
1fKlF4Kv47syBZuqnZBUDm0A2p1n0BAGLFwlu02QyVyrZbnWILCLOLLvcoFtPD8F
g8+EAD+ady+JJIXl/PFoufbK/64dwcRESzO1KA5EmrPm6NxblGZr41vpgdILzq0u
wZbACikzvlixcKRvFjrTbtI8tj6JGkKqBKDQKJAoSv2Dl7O43U0Dc9p04t7iVGr6
Ffn4u8hw/zg/Q8/AUL/fSXXL50g6616qCLBlZ+uitpJFc+0rQkqAWFD1YLFJ/QAj
RO8zYuu6GnXye99GWUCWpd94OFU7m12K2mLUu+r8EMHof1x56PdYf1zpiHWiwLnr
3uZmaTiOP0QvkGde01YAmfgNneuepp5ruekDqqujNQnlUpO8JRHM9ZsTMjpumm4v
K1pP76JDtCiZkhw1+DrR/L7L5KuNJoyVVNbI998lIjXJTx39Zm9RStV/IfSaDmZJ
27jXbpm1tTyTOqwqrAr+qEBxxQp0hk2i64ctc8N6m/fb5ORVa4tazuRjgQjQFAnw
7IZWKP3nxZqEehQPDbIBskgKMpjWt7Lk18L9ab36f9q3b+mLeWB71vEK6gTzr3St
OT/p+TW0WOQn1b/EGh1Ern+E4GOAMGvtORghT/WNpuushB+KOkJju5MU7IBBDFkf
JLhRxJoBhL1YpoNYkm9eRdIMWNZDwVXz0sPoha7sRwJI8ejRtwKfk/MaHx42ghyr
MePHvoigmlsZUFBt+u+hBqWHH1QX5+ezWydmLC/Md+41rkCV7IaHnujlP8vs2OtK
IELwsfvbNmCTd2/j1IdcofO0KGlpEpH7oTquJqkoq81hL8PeH8fygIrt4aNfLGX1
d5zSNxLSBls0CfMh5JkyQaQkn+0VbjRgjF48brsFwmoR6+FMR88XsuNDzELaXExW
BUifJczCfkD8E1r3ulwKBGTRvMfapNpXA4W26C8Ona9OxWR2J/yhmQS/he6ZvV+8
ReKBXozInO8BdaoMzP8S59PN+0dXJcOkePh6H0xXtyEfQ+o8tQsjYsFuboSd5dH/
iV4YdNj+5lphAXx8VKUpxxVrGe6civ6tvNJOAYOeolRa39WSC+cxANeb8rDPoDpg
FLdqg0Cap3PhDM59DJI3+ciCaVoDLrEOeDX1vti7Gax7IUjKMrb8/s5+j3qarMm7
9RukE8l/4hDg5fq+MhFePQKYA//WKSPw+/y6x26wBMzBUQvP0LTL4pUZ0RRG8aBx
zBg1jmxmd5+U8AcmuWOaINdeZiz+sayvUB+M8QBOdUgrqJZS6t23zSg26dCBVUtI
yBzPWoBeXfYBXeiDhwa/801Q3voA0edaFRXmyckjlKgTUiXZP1xyUsBxefJ675Tk
OlxZ47pZDtsqEo740XrCaPLGMjHBHyhQQmab5ogd78KkBW4GgAw2vAcrOuFhKBgT
1eV2j2kmJHFfZtnXWJzUJcpIu1ZXZdAYApSsuE3JB5ihk5zeatNiGenIqYIqD3AK
+TIgJpMtiWwMrU13rgCYvlGg3qED8ZNV8cgsDFcrHKZVcxX71YBCB4fO+h5J1Xdo
29EO8x6L5Ob2UOK4hOsPlBINe7lbbEO+Dxle4ADlD0ksqsk8kg1b0FTCSgbop+OX
xTrTTwM14qwQEgMm+VlSrrPdUnpLQJF3ko+nOKu06MxfM2Tg9UNY3HmZLbCvzKYn
12W0C8ps9DanR+JiYqHd6/7+64V5kb4vnVPZES+cqLTgFvut5AOQAO4AIw2JbTAh
+fXGFCL56HqkP7lYUAAczaT3qGvfk4cwxLKU0ovLxEKFrRRWZlda8e4rDxHb/9sx
twvvYQpjvWBuwyqiK6Wh5xDEHF9wrZa4tTa+HzUzMx7crpNbMjj/J90AlQw/0Re9
ZKeGMmBBWSwEBWZzB0K5EFRLEPb9YGSx842g7U7L6LI/w4RIJt1+wZe58qJnep7W
tv2POBgx4yxU/JxRgqeBfGn0lqIt+KgF3fyIPqpA0iiHPh+vcu38vQqg0bW9tbBI
uTSzUoR4nLv26Lw1xLsRbDRHVqPCWLZ2ZUVcgLgyji0mkHKHiBLLlM0ptmVaVvWE
2HpDy6pnWRUQbhnYNiBr93SOlwtkSGGfGI4iijgV4nm1aWYZSxi88NhQha+YR+qz
+snAXe2SOXD5RS39quWykXXjUSzNIO0PaHJS4rT8zsHNViGynWCw9WR2SjwCbZ44
C67XsuNYYEQOf42pLVhs1PsfpCZNWQ6anuRHb0sP1xMO3//EzqcU/4pwEC6VI/qs
OmBleCMdT9ealXKKSK6g+/M3xk46Exh6dEw5J+foVLpcSwzPVV2wI///DuKzclIf
yqM0jTS6dOGPLTkiY/YUDYZB9wdauREPaR/C+aJK45f5EPXow5gPmBDXpYt0YfdM
YuOJu/s1tobF/YDBADPjZVnACUxAhioRJMyadAHXubq7wyjOPy15E3Ieb0UKVChO
fTiTzmcCJIJ5X2XmBpYafDXA5bB3rnnEz2D2NEuM1a4M5kLbt8hCb6KBR5k75I48
Iph16S0FewLZlscQ/XB1HuIC6scuLqGeWrz7Tf3sTFWY8YlGGsF3OKHAnXnXqN/j
A/kl2VIGTJ60jPP3+D5WoOen4+EFq2GomeAEfh62HGW/47LtDMmBQn/lJpljzp1m
Co50Pdyz8gfFkc5C/Z3DIFpkhp5+SwYpEs2VPl1kU39WlKWIkAk6wLGahFFWcQ3T
lIRExnWHeZjAlvIdSfK7aXR9zXZv4+ycqjAMVq4j8SLRMAHJoexb/Fc+57gTkd9H
V3qWKqKCqLhad2lLFn8RifuUobL7EPva6Mtpm/250OI+WEL8/WiG7MSURZvPPABh
z52U5Zie+n+4nDhpm4Qus5bgnMO65vHJ/EJXnRHvF9xxMQRA71of0dzHTyB9/ldN
HjrBzt6EUxkgucFyBLgHhqJYkt0x8MWjmGoutgoHx9UxBjNZ7QHZXsE777vTf5uz
7FijzpR5hoCS88NaAZdR+Xq3Fu0a1R6x4V9RREy20aAR59mEjMIg1yGflLBHmihr
L1z8pFVN2zwUbcoU58lBvPGvEmeR4oSMpueZ3U2dmgyNtjFzEMA+YGrbCms5WXXS
M75S84uky6DCDMHY6yQC2M4lNxMJKEYsfv31DwdFGg2zyVcEfq4dS6S1NvtdNNjI
1/7mU9Yc2pMA5epcGUKl5BmUKSnXK/n9JMXXMXtGujTx+DhIgopKqoFitXtTMfxk
Kx2K1x+IdY15irb/ZcGKV8g2+YYlnGhBXZ/n9srzdrA2nZC4Zd6zkCGnuQID93Db
qaSNhOdnxakF4Pg9ZZ5o8bX8rqE1F3TNo0fUmdE05CaN5RZUgMJmfGeJm4NsCv8c
KuoqSWjrtzNf0sICN7COG7Weoz4ybFE5ZlSF3toxKVLIPLwcPsaq7pxBBBfIxmEJ
XJO3gr9g0ZKgmeRd6NRMUfo2bj6jOJ8x+3NdQ0nvx0rBOZRYSfQi6g+TnqSMDoUt
Ha4Xtu/YDwICmDqI/l0g9Gou6iSOemXV2hHC/W/2a4gP4leCEs0MWiAxxLDwLG1c
VMKjTQNfYkH45k/k3ZGuOWbPdEwloVawQCq0bvxFzql9fSqrdBbSB0pNf2djeGQo
LOtxvT593XaPwUL1Hxqx04UTlijgYGCWzNy6nEJSIkimxpJAB7BYDa6L3nx9kS8/
yIMGfp2bmCjkjptZApmZrJTeVePr+BFWLis9lWU79vOOck65kU2sJQ4l0m4rznyE
byHo5FrH4kCr3uowqphlW9DGbhW4EXmyUZuqgYWPTWvviV2JcGn2pGHbPnk6CSEz
8u/17hEBuRQ5embAYS5bDLBkqqLwq9kRsITmJTtmcvZLwhyJOMN34RRDMtK92DWt
kD6yeNS5y29VP3rZqlyXsieMoH+UQq/eBn7DqCcHq1vonWKkc/uA9T2fQNH1n9eg
j4radAO3UWSMfhQpS8G1i6fiG/VYI0KG+QCf5IWf8JWGV29x1cyFZNA5PTSpYgHy
e5dNfcjeYMbqRvwQiXmBTvzfmExEFWf8ARQasit4DVtie1jwSKtim+hn2gcWT36H
FR3Bx+iHUXelHlhHP/dHYbK5b4rB0+dS6UNTomRb61admrIhpN5lCFtCEiKKBWna
ugX2h0XCJjQJlY86osQygZ607R41ws6NMydSd2A6WSNaNQJVYa0++xdjGjGFG/qz
Q3IGLWIou+sdqxAtBq0zhrUMjtvXViLNx1a2DYaP/vWnnT4IeOdEj8wMJ+hFTfK3
LGRsr/wVrdwNnw+RG/J+Cjh/rqGn3C6+CibAyJf3HxdD2xefHNdatMMf+J0yA+t6
vz2ST7Rt7s8Q3HrgIas8aBY1m+93XPTgEL4BzQbT24bACwR8OuDUMlg/5vUFaa2v
YUY5XFHP7K6LnKEpZqka1PAt+1K2m1VNsEWMmIxVB6QuN6/xT0eaIyRp/uWftXtW
AqxXqsuGM4dm4MrRwLS33ORY9a8sUgvxWJoo4/eCdYv5ogYpgulf8eUKYPSytNwn
qBU16YYkJYcI2BzsAZToRdhPcyE+6+BckgiuQa6A07ZCzthFeqvXUumPoFoQB3qc
EnDDPPeulB7qrrf0k/JrsVEYG94GWk3FG9dR7vJuHR5YHdKodCWQ4zDFNGNk6V9V
EtxrOAXhKuwbSu40WjEt/Ti95n0xgJL6hI8u1hb299JhUsAShgxGHfvnhTHDIKv0
CFMWztHIw42/P6PSnE8bkxcYJMPWOGJhfxalv63XC6Lb5vWsXbTOlFrtZwxb5FoO
BNFwg8hl+jur3Kw9EeYCSFCkaeA4fFJwE8sghZVfjZAJb07OT5+omRVPSkHtzxI5
FLNTbtzfEh/afR/vVi/ZJtqOXoks321/7crdu4nIiapcMwv4G/6AM//ps64P8h2Q
hGUKsJDRuQJCewsUtcdJALNukAD78lN48mnWZhwYJOZAGAj3cZQ4O1xJp50MFGXT
B83VWJf3744vRlkSa35N842VApnx+lMFHn7aSXqjYVT52OBpQ1zGD15RK5Khzd35
cAhrgEBCElP2Ac4D7zvM6E79kVqpk+wF5u0kgr2T1Gz7nWH6eujPrlMhH3m6XPFM
GUld6sSZq3djT/1Tx0PNcD5yO19tqmK62D/ETI304WFu8Et7IJaCDOTssznaKZpb
3WY9qKdz6j42DC6JNDmggF+ntvPLk9q6pXT2igLJApBwR1MG4yA8zaYGX/7R1YNA
g5QqwLM8uBIpoK+PEioj2NumaWgX9UXq/sPJ9eNDPNkz8t+J2pFRs1AWvYW1oHhH
5bBc9nR7gSqLZ03VKiLskjODYu2reUGhaOCLb4+vAqaA7V4hDTTU0Rko3Oy+zNA6
OhoJWlj811G4ONVOAM9i8pUsqFxMk9gowyQfJkYdabd/Hdp8oYUiknqGRk3kJmwf
mcA8Qb5gXNSwDW9PL5V7rvF1lUVSJnsFMzxfXZCHJniyhV7RJvlAcA5ptA5RQdOq
SrCesRFXP4cGqicsn/UQGuxtui4HlnTkrqcCCCT0V63GnBvUblqgCloN9uszDnkc
FMMkVpOXmstKJaJ5W1Y14pldap69IYbp3MtCfC/cfuRrG9fI04p92f7pFksI8Saw
+J2+f0jvELZjhmGMMVEutT3IwjCTKCR4/tWdHOH4yPgv4JMhKzveqq8/cPj6zCSk
I99La8U91gvrX7dHcczqDJsj3DIm9En1SgxhNkTZaFOh8/ZwGAf4Ppq5UPgKVKUJ
6GO07iKiy4jmaMGm1ciVQhm+NGdPWpAp7BcTHTSq4Bb5jOHF5QlKcSdhgxPLI1lA
PwycdCtlJNhpfOK+ZNu9LoX1ocu31SUf0dnOPgxd1gIOqLNY672swfuVdsrLsr6E
DIej/3o6QAWwYvzgsw8oackObmacdvOH13hJCugFhhQIsQqHh8/4vLp0eFc086rk
iJwxfn6BM7VSv9Cyw1mrMWJqFSPyPmQLRpjs7u5E+6DjXqZs1jWE8giBZZ7tuceK
ZnQXGtegDWc2I5JbNOVsxg8/eupNME4ukDikml5Ks+MC0oq62I1a59ydnOE2yl1S
CAU2Jstuhx8woBBXZ9/b1+reYSk6yFlCxbTlT5/Bs9B/ljAEGb53+PAVmzj8zgTq
/uiujJO6NktMT72S3IHLHMg2Ka2EySHiLkaG9GP22QMcFBLWa2/Xq0WIvRSfYWsF
YrEL2a6mdupESQXAPCW3GsjLH/L4gfbDSsUebJeiYlSUvRqxZwHZ2vR3qgD4wKy5
wEsNTf9e1hQzAcuVHgPGfj46PMD0lAT/7krEh2Vqc0HVHEayMi1UtYo7y1gcy1gC
FOrtY1PwAgVlGDk5Z8SNAW33vyBRfNpdt3+MgTnKVcf3+Hto81C81zpVqrqM3sId
zTEEl4ccEoJAqZF48yfVTsFiEPFTephSGCLtvns0Lqfl36J2qvrFgW1QOMzBXk1q
pkkYsbAMjcGKVdYh2+ILUXAxdxyesCZ9POqZ9XMH1T5ToLjjfrNFjRD3/iMpNspi
c1rA9qoW6g/2uMpU+DAky8GO0gHbqyJlDIHX7GMGCMNLo8Qh6pYcic8humMTbHVn
cdwhNbaZAqy9Nn7m+t7KuEkV8q1sif7FnEEcCFNhgfaEB6iuwzhpOls0w5TY80or
UFqlM78S1K+W0Z9V8AEn6Lzpi5XA9Q+lzqSMJDOPG4fhLDlCymnGxVsvDjePgp9p
T+Fi3iVM/Hmck/V+/UYGx3CD4HPJ66ozgHtLT4koTlild9eCBizsQcRTnD/A9oD8
06sVU5QYuE1hteHHQJWhxNxtZvi1uKqWOlSu818NR+q7G5epYC0ebhTLdP7CYpyM
9LoZCxU8H1+fX29NZqWn7pq1Dg9fEsHQDpQg6MZP1IDnkz+dyA1SK4XRetGDcmTC
6k6H98C/FV2zvz6H9o6nw91wb+re1IHV7jlxhj+f91QM4uz6/Ma/e4ECadWIs6V5
Tj2/NpNOPDvYYjukSHSLzlAvU38mTqzkapCVWNpWpy/suV7qCHXe8RRuPBXSOF94
X/01iHZpqoyRvJrlfNLNSMaVnQ6+gkmZdUHXHtgi/VhbCD+gYHQoxFQdCF0zIWur
eyPRyQRULMyxSNYyp3jVNBSg/7n6E0DlJ76o7+3YCKktEZFUx+CUwuamTP6TRV/z
MpLG33mqm08SoBBN49aD7goxig/XtFjvMSa3C++FUvk0VdVdf5/3td8GZkrsPdfo
Ogg326glyy9UhNNYlBQomYQUViZKunHpDmmqKtrf4p6yiF+mXmpvF7P7Bjot3w/n
+nQ4RTT4MOtLzQFLSnhNxN1UQrmqwpyaCqDrAqAI+r4FE/i7yfI74hjzwsRXGQM4
nnOMNKbusrU3JsefQkF/VwYoThgiLOYjYjIXdl8UY1mN/nXCb9eh+Fbre2rQE/HP
4nNXNhZ5weY5B/TV5JPteFRej0l5o4Q+cdYBnXnMuIos9MU9HyhT7XDxMRvvSQ+Z
GolnBQad8pShrnMjEVuEovWhUppaZ3NcRbk+q//PNGYRDH9xFng4bJgxfiWcn/f6
Trg7ylGXbPOn4j6G7nKtFjenLUC/nDCR6bhFM84PUPW4vnSWGDgIbZhxEFVIDMDU
v9NwNYUJRb5H7xP+hTEJjaBoPH6cn0atlkYm1pF9wnNc6dP3Cgs5AUVOCPVbkZvh
z0ydfh1CALnjoYg+C2KdY8hpgWxzFHqNM9SIP2UMXqKm+jXx+a5snCawicUWmXKS
844UcBzMgrXcdkqVGoDF7vEHEd5tyIPi46YtULt0L1P65LDJe/GHK3Vq26yxY+dK
frMSw2PLWm3BYjtRNjXtZUlMLKDv5v7WkJZI+mqjBw1STV49N81AU4xeDLhfbJZ+
PGHjlf+n5aRbKWpzmCYnPoMDXkfooW1qatT1eCBChvTUUkGgIDdwG45gUxTssTgP
/LZYBR2Q0ShbkY0Xtv/EskBmg9jHjIxktaKJ0zfB+GZ0u9IJmXQBmj/ohEmm4ju+
V+AlBjLnyig8VwwbaS/sr/m9cbnkMC9woJmD/P7Qu4ZnVkVlLPT1cgKcL6PXgT0+
H8w7dBBJzOp1YnZTKlmKWVJ1/B84Q3SANBFJlj15MEiOX7WtDZtNhrhe8eKpGtg1
poc7eg9+MJEnEq4eZvJEiDOeKzEB/OJRgZ8S6avFRbwDh0LX/xim0lSjANelzpdN
LkbYzzWlsKYwj+IFPpjcZGTlIddO4xPv1K/y5zG0g5MUgoohTd0ukuzYxEzJkBUT
NVyPunrxIiI17Zt1apgzLzm2EE8lG5VL68jwmIoFEaO8U81QtGk19Zuk76n6B7lC
zR/gMHwnYNs3JFIlrC7Dy8Tz/KTk3NGyelBoQFbKQXYKuL3Xu3HggjuwLiTQ7S74
dJkKQemwJ4fqnO5jir83oho1Rb0DG0EQcM5xNf+RNK5rfNIJ+S8FV+ijEykDMsYN
/aWk9SsO8fJlh/rUkM4mglhhfyQt7Q0c7mIGusGtmD/C9yHXZmZZTUoZXNAvPVST
rtIWsBxvTwK/xHMgIR/BLCCqp5njWidWJd03A2uGkABAUTuH0V7m1CzcnJx4PnSK
nzieu9xD7Y3aaM0ooaNB2lifd4QStKUBwDo2WY/NGAt4kuNPdyDXyQ1SJFBrsUSk
PXst1kCzGZtMToAZB3FJFogL/saAbkJsuzZMkpD32hKZd3fcJif/O5diwsuXkneY
Y03Du+6MRrE8BjnJ0VLvUeBO4ILcvpqS75NQPbWZmCm979yTt0wOnGa0yCMqUqu2
/HNLPYXgl3cKENs/mJZnhpbtA3hUNtIug6QV3tYkC84acjkjgCWnvsm7B8GnWPxF
YRApsL7vVONpr3oRr4aSiC14/5qMFV861LMFuKuk6yBcxFUWnZEkWUXNqtBYq5ZE
BvrcQDLmbhvWSTy3+lyQkvweC7dgKXL35qORO3S4luexJyPFo3A93gZZUFjhqRU4
Yt9o71B8GrjC7IGcmLsLY99j26OYeB9DO9+8ea2NOtqybjuvD0r1VIrmndxN1w9+
Pop7EVcjO+IpyQ1WdQPem1nYt8F90Su30IXz474+mnAKpDrvMcTWbWJwyOhKvSZ7
ghZVEEQQz0W5IsMzZQbOMeV3/H9vkmWusz+DKBPXnTWLJn4Z4u2qb/EjwF3byZLA
DfIjbwIZwRrATVWpXJAdphOG0vKL5LamGkQzAZInsX/A0W6yI3hoGHrAxWsg+7Ol
XU5FAmzeU1XFuQ27mHSewxirFj3LdD2O9Mky4OF9ExGgUAR1kcCpkmbmPDeqJj3v
YlWhPuLDvKKWoyWn35y30VR4WHMQWQFb+18zZ3kG+BJoyMRctcjy4Ew7st1bh+xV
/qZUYT9mKlUj4dlg4A5LUXe9DTzS5pvOxdsEvwbWoVmpXjLTPtqaatLEy9Hii7WP
qvS7z+gG5DJCLIUfcR9ydssRtm9creFZ7unKKSgkRuB2BaouBnb9n0dP3OKRNrKJ
wvHtzGRsIRJZetmFvq3s/tDw5U35I+Hj80kpH4j5/4NTNHSEmKj/imSmwT64bpdW
4gh2SiHUMlj/KyU8/ICn+SYdkePaqvx0RJnC49Apecg/HEricU3g2/3sRv+EpDFY
o6vq4eH3arKqdNUIoFsJZBGDq0tmtMLftOPXXG4nS4cwykLiA+BWX2kzgoTSgUro
5R4J20DFgsOEf9l/XTDsJivdQcXynwBZ7wzkP+OjGwT92lXOA45iFGM5sPw5eiTv
hfNkskIXl9xYwvhJvZbsP9Bhb97ftqQMPwx/G/IhwLg5qac+tU0sS687oZK9RK0M
llA4nx79G71dk1VJFM/DmBp6/J7P0NZ7BHzncaXiwQkzgpTN61twLr+2Vo1TIu5j
OjPOo03ytQRQCdz/zgsXG/5QGXIjgCoFvrV0l2oh/6lg/Xd/v7CyrQtPyrJosFKd
ancJvW71r1/InnO448z6Mr+ic9iCfcv1TFBd0jVV5o8WHRX+tXOQmNgoUJq9zPlx
kdTB3oKOWQ3QZKN6RiSfvtaqsZiYEJY/mFdJXQSzUXJTlFa7Ev2Lch2HUt3q8ahv
Ric/wx+iN59g6PWmZe3cGDbF/AtVHwAD4pG9qwiTWPBPQ8+wcsCCnO3Xa85iZYJY
x8YGFoW0xTymC55hMlc0hiCFTF/PK0RVPOnu7wVxe4BE+DYJxYRGXgDOAx7mskm4
lDytWOD+9PBYzd91IJg9As5KxOQw+ftPNVPGl3N5sQUtKpkHyPhZZ4USQ3k2IcSE
/HPsh7Amjfvms+WNqwTWn+iT7jH7U0IkMZxeq0HDmFWb6SiGcxYQ3TkkREtggJKO
N9FDjuy2g6wj5wn7rbh7LmOpm4+h0qyTYyqRcNVBeaQfm9+foWuT812gVjgTlDU0
WhnFx7jiegWOPQzyiwHOJr/k+o5gWSG79KE18hSZ8Un6EqRAY+7JophAy8MEI6Lj
znJ1KcX7VvCVrv0OsrZRJCewVXyA0hnHbH+vlbRy4Wu3C5/u9ibRbDvs4Qd5QzUl
d3YpLWdhxvgUhWyhrIohBDxrdTxjrDr+siW6dNErmix7F4XKRWjgPb4N5hRkqyF/
WL7DtILpmKntcTY2xlZBNcYqHpUgfVopoSPVFsUqKCKKkSkLg44+9CD4ozIVHmDM
VhapJV8Z64zw/kqk8ccfgvYNW4kwFZ8OEJmfRjR+f5gWgb5Hs2aoCb8e5LwcBzZw
gLSfoIRZoTvYoZLlbSo+nD0K3b//9YUP+4/w0yNkOvLf3X/E3E44ySPoKwKkaqee
qaW5N8XuH+KMhBGAvjmXpO/7nV99ktvQzQuIwEEz04QUHT2Fl8qVfzUEMlKuo43V
SiDkKz+kNX4d6YvHxraDXttTlRDCuTOUoGLwhWvLldOsmpVuThdFZSQTXQyisMZJ
aycfxujiY1K+sndcrp92QvHB0XF0MWjHnwFZbomCxx9KewkXjLCFwDbZF6e9jZBh
7Qq2JM7ZRGtQvotvQbHgF0wMz2fbqPGmil5QvVGKfjx5nhoC8ArP5FksWi6ASpH1
xPBCAjOO36BoPxxsMV1E3d4x8LsRPotQhYu1FoFTkU5CXsu0AlkEZJ4hh1D3aITb
Sx2u7Mc2eY0wcGU5iHa81xlb5IBKuzpGgOXBgmCtNimOa+N8Tg1qokflweUUSaTh
X8tQIctQmpOQUG6iZC4WdImiJz8eA4psWL8nkLtwvsU6c7605U64tBzYtm5eQ6Vv
wOjBTpptI/QvTJQY/nmGzI5wv1kSYld+9O2FeszWBIGQjCgtjny4utbxkPZUIZkm
7wkzixzXmaLesRyCsYs0hlSStqNv2DQyR3/KeUbZxHutyPWNyvL15HSV5vi4iBs3
N3EHZe7q6KlJHw3Ag0KJ3TaFS0zCZmUC4+nX0dbhPFxJmZALKtvMMTJfkSUcM/zf
99XgA0gB62qNbUUlppKw8IQDG3rlV9kUjUgxNDc0K5XX8uqBQ0ZFVSYK3etzLN6q
d3dZ6RznDeINazc2zKHdGK1lxFUTHdo1BL0ahzLKiIDaiICVJ25zW3cPtNQ91kCT
zQDYmMC9KAipGBlhJuhGPbwq7lxa0F3jz/qC7WLxn6WKEd9+ofWromyVLx1WLofR
GC0+WrRj7kubyTfTtCgZ8IgtplkMY6W7c2sWPicXFJXN8JqGH4Qo4DS2qCdjPBSV
ENzpypX8fGcTP9rx7ClJQD6GM/hFFqrWqyVrA2WQ3z62+pwdn5NlV119Y4imilxD
IAUhl78IE4z3piVeTu+4U8TBJ+xUZ+pm6/+g7ickY+6us+vkAZ5brhCM+zZ4gMQ2
UgvSMA1Y4BVchob8JbXI+sB1nXz9xjFlqsrCnrfWibPStypLFWnP5U2Hw4qEFqj5
WnJ2FCO61uNmDZEQKZ6P6BzZ+OgzjZPItmRFA4w+hM1LJQGhBrmL7PQi6hXfQ0hd
X8RXJl13z8orePn1pm1s+Nlp2cO1NE8w4ur7GVUgBPubhNjEvwN/pPGpsNKJNx1P
XcYHaze+74eZYL/VHYHzAb1AdiiYmUqKhkAKY/FRKuXa+sscYyKZadcET9Z6swqx
3DWFGjTJ3m+uGaqWZtkJt3QXefhyYydJZFrAQu27/lveIqm1i7T2ElyS3aW44fK1
USAWuL08YVaGeTKW38o/nVT6M2MggGTV2UqqxAtBKlWtHUXE6u2uTrcAFNvdsaJ5
45uluJmcfqwQLxXm34AiHahIusRmELxqtpYWw2zFsYb4Pr4Lem6qQWl1PCO5rRfQ
BxA5kO1D9RUNfhS7owVQkFZxBfh0QTqCBQu9FRCcO4C8kveXEBPnYPM+WFX6Xwm6
tdhsuIKAkf32iok9uhu/rwGRfVm9VI8qBFCom6Bo2G5mDTjwTwif/WKxPPYggnpN
CVefanIjlcl33lCZs4DNuxUA1HrL1d3dMZqRL2WGikDBXUlalGLfS4UVlBUeSf73
39hI6r05tdADx77/VnGPtcPjSPiChDs478eMDuzyCQ7uCd+XhKzBIxawOWzkoY9I
u7W3dsgB6H4Sz/5rHSOPkjBnvZ67xCpmiflyR0UscCsTLYzSslfZ4KrT1lndSMqc
XV7zX3SwnbJ4CBNKI+HFpIs5bujNPvJj9Ta4yeXChSm8o8T/GJhds6CQHM7PQqh4
NCH9fm12C/1N1zWgvsP+V319A3LFJOdKRIijirfHRbmpBdhNQtlUz8jtB9I9zj3P
TBjlTnBxPxpUF6TTECQAZFQ0NNzGYT3FWadjU//pLFl0UcP9UOR3ZvoTozgTHBzB
kfRoLYnOT/vHfQw/NKptrjmEReSyLdSFbYlcBYX8xA6PMFUjFnzrzeYGEdNCBBRn
qgT1yQZmQrhlZ5DL2uWUB9KoNuW5peRjGKWfCV+eS8ggafyPa8hA7TwX5vfQ/SVP
xRbL1w06SUB+BCQUKuUNsIHwfjT9casPD0QwHShdXKqZjeMoTl4MBFSgbE+R0WwC
i0gS+zPgvIoyWnVnwP2tuEoD8Yx2S9zpBqzXqyCV92enm8KeH0dK3RTO29R50vGN
tYZj/Xub1pOuRIOCn8j4sMzvmGyOzhxgrSl1kmD6c3kMvce1CPvZPgJIHGNkHyiM
o6XpeYhCDIHv4sQtWu2llzY6GXGUmzgkbKnFYeXEKNhn5k6YWjKwcnMEpVuUeTNI
qhr1YvSWIKV6OC0D7g8qOQC/zTL2YNIVVEGqJVNI15UajmYEK9kIAG3ZdkpaJoRx
fCv28DNx/BQWhA6eWFaR2YHTN4ZGE//wa+UeylJ9wEJFFnQkE2ztoKwUvwkTQkoo
ijzgioexzuKaoXxjoT+HJLlV631HAgd1SH3DOyT1WGsP5Jx0rBOVyO19Pno2JhiR
vDhx4GPzFXigfG+5ofK2lPBzTfeUl7YLPIr6R5dAMYDm+xfabpbuR22sWlOQJil3
jCaGS9QXegJ4mAq1hAEvMhPMoamx0HGt6EPVTeavnCMEZ0q2cT+QWgKCtd+8NZHD
ty26ICwARY3fp6/Z88kSDPy8a/3JOU6WotUU9LRZzsP772ECQelsJeKiRWgtGk0y
OmEdYhQePVZJvknNwzFwkvsd8iPqqB0ktAPY2vTDcU1qyzW2l6IMRMv7mC8LSQ9p
FXlAmA5TZIxH8QQCogTfFOyzRt3EeYEKjS82uHYVoLjD/681pumCaqbYcqhfsjsS
iyUFIcbQuwnV1zqNb/YHCirjjEwPoO0RwmHWhtzN1gtJaQ2Mdtgn5HW1xQKk1N+Y
R9DuejyMEiEGkpDjVGwIUxOFPfZCpnfMPX1kKMJ3PAqwOuxogbmR3Ym+Z0B5U6Z7
rQBkx4dfWXD7vCm2OyKc/FckKwqqjgo7VNMpGSnu5V8cW/WoDHOREBvtlCoY98HM
+dH0WwxVjJLrsxTb6B8JJkR3teD2TQ9Wwo9G1zRSJPMWhtWlYNi1FS3SyUG5wgD4
3+SBDkxUSXKema2nadAaaogpPP4HGRJnsImWAxBmlXgDgmDOgBYajnHn7oK/G07h
l/c5jv5xUFXmdDrHx9jM6VVVNO3zHC6wqNFKyzdCfCc0iJWnc2Jr3BA45+TnDPfL
38L+4iCn3bh+kSzl7wUbd25x4T6myMtrweUBdRFZn9CQvpA/UFL/zNR089xOSvea
5tU2gKr+20+7IViU5LTktRaHymUY3DQ6B48BnAFp2eWZ4El8sPimZjpw+nRHiZfI
K4eQBnyPWKGu/RVf2GNBME4IoYMCIk+hG8qfZVz4lfdrGQ30lI7VXv2RSooqLKjI
PuWZC2gVPrnn3m4/GiD87smBtUPP1h9C43YipBx9I0DOPS/AABy0NBQXKSUcrSYJ
HogqF7PaDUQV3wuOSNug50k27auEj2UtBOpZ/n8DI6kNygZsU2jGArHt4HHGWi4c
hSJouIhBKxHWydBwC+PlNKpifs91tSnq0s8VqBL7g/hn448E/JGXT0eA2iycionn
AQS9s6LWUEjzCV0YZ9EepfMS6+MMy0dpa5gW+nvNa9OxoOKkq/XI32SOt7oPFGr4
ajJbKJRzt7Tk4EL4oC3jnFvz9oYGKtRLlLykdKP0vebqA+j7M5TGXqsW2IEpEnxn
vC27LzgYp4kvVGSuLUnHq7RuPr0C+hJnUcvSYA4LA8Gytt1eBgyidS47LPkNJMJp
4KeLy8KyXx1E1aY5BHRaYjJdTCsfhFQuylsnEDb+3uKQi2JhCae3auM2Nky80Ee0
VW8D7jTUGpAJUyw0gOwEqJgVmcLPJDb639X0eyfDeAPWDKqeOIfN2hIvWbEIArRS
w05DMCTcksfZclIsJOlXwsQBRKMXBDhR8JCmpR+piIRT/K4lsYDzslj1edg8DUcx
Lin+m1fQ0klh6X7u/k33/vdjGrKCe8dlkv0/wtWEAfJJsDRrSNa7sp9BdT+Y5L+j
vrnkHHnL+0zAljqWmkQA69XNDwB/I5HxT3sj8UqkzrpuCbLMOxUcGE99WWLfSB7v
lGoX5OpCWY/FzRmFWfq4W/ijgf7EcLEW+K7eAItEW618SHSANmz8LAh0Y8JuVBRD
C2JUoriXVbjyMBhDErSmdQt3VzJ4PoydPAUIN1IIPABm1KCJJv1Z+/Fl0kvlT94k
7t/Hs1oFRwnsZW29n5BsZ++ECUjfu2D/2+yUP1Wlz9n5B9ZMKeFXCN9bwp1VkVxd
0V1hRrjUeUVpBOfuKxb086MyMkXo+Q+dYsng2/Q73DwSmoVtQIvi6Cd+kcVR6Fjs
Xm9cixYvRYBcowpaDZkV4fhAIrBTjc9oSW2D3U17uA+QRkOWENbPQa16IejK32HN
zUsHy8Eg+eQcOmxK74/7+k8jg6ogHeluMBp812Tk3EqUjNM97aqnxwewrLoTgBJy
+7CaAIDVTU7KXySfm5nJmS0EFLDIn1nvKALb4kCKrKqAcvlQfk9Yrg1VWsBNN7dv
muNtVHXezShFRbMwvU7Uwme29rxS6dRvivU8bUIiHdl/sYUf7QzHQLfVY3JOHmU/
jKViS43bvwUtMz7PRyDxGYNlIxY6YM2TeYFUNVotrkZWJqcXSMkju1hNKVOEKAsu
cWlYtCIQ1UKxtpChT7FVrxv/n2HwY1o8U84AC5MKOOYKOuiExHjO8NUy7IHKaUxT
LOIG0W0GLYofL1qFdMjAhGiD6mHrjxqyxpZvunifOsGCHxnwQCeVSSMQek2RCgNf
BLeyPN4peRUmCDUKG2RBnP/rf5tgA7z86RC5At8Ytjzzl9i4z7ukDxRE9Bsa4Hsj
UNrgrlDSJ0q2GZGjPxAytOD6RbnvTNCohCkSYlUWjhuEpGXorfYyOkoqcysrCfhn
S4YIKTf/bW5NZPEY/fucwE3NucwASdDSc8/WSgJY3mGiqdwXKkqOUMlMh4G3uXx0
Ag8T/fIC6Y5dmbAUA5nt9oQITrvPTwIokn62FT/BP4EPBhN80V2EjRwEAOg6HEzY
TRTns6C1/XH4sgpLChkWL8c1PhL9FrDInnd5RLAFT545GbZBCGAZb0FSIkuAp6WV
NlvpRqCgQ/KSgI8gBtBkkZaKySnapAC1T220yk5SNKtyI5Xf7Neo5iljo1d6H8Yu
VWMAxroydv4birFUfyuzKRpdia9SWwcPhmEPiSV9V2Ri3LYCDxDjMwIuAzZuhDAs
pGqX811yWNRpd0ZoKbs6uxHUfD3Do2W/mY/gyfdSUm2VfwGmec96/5GyIPgkYP95
TWV1NFsJNhFZDdjsV179XXyAc+KHYpJwloWAW7U2c8qsoGkoTWjf0+X2D8AuxFv+
QeAEtvUx7SMOFHYgVy+Gg5zE27Hr9cMmofDXuT77gss53p5OewDNX+eBadf/UHJk
DtYMbotfMNzOvRZZrBlB/DpBXH5OYNzrOEBUTJk83HzWxkFus7GymOajTyNaC3Dp
7VzqS90xHRBLR+8I6+JqMFGwOY/nV0oSBgKgowtG21lBGUmDFNXMPXvxZ+hKnFFU
ilU8NbQclSUSEmmK3JMVoy8aFPUcOp7sOn1zqmWJKtYP2ciJlgg3w9bKX2dmQ9Jo
EyKMtTK4H5MoCssyynBDQZ4ZltzqvMAB4kflJuWImLGrqIfAJeYclQ7+f7mkPjOU
B70IuUxb8i22HGrK7FHqwPVT887TO0m4MaiquC3oBnlMt9R56z1YNmpIkbdQPSsT
GXd3u2IREQ1PaHs8VVupflZ04coKicSO7tMJjATculUCJ0SoVRa1F/qWMNOvG7Ih
sykIzgi/JPVHS4bUu3kGalydbbk9xGWVh0nfU2wS2upnim1WIUJIgcvpCY33ym/w
xkrRTsIQgT15RYhis2et0rr9zufGftz4oCOcmbW3Rs0eZsddElm+P/8bKmQDP70n
+HsNdscCpcObV+sQEZHox/Ec+l5A5Mpk2RjQ6REAcvnfFf2A9McUVbcWzqacQK9G
guDOl50Lhu8ZAC8zeulyGPMltmkRW6fPVwKbyLAO3M9Gri5ZNJbxemosc6XmtVQO
3bhhBCFwf5Kd2IffFVPIpb7BUjaG5cG20Go12SgNOzka0smtlkLTQLc+V1piZcK4
Xai+jQQ0oM3SMriE1iLHhvGMgJjTKQL2L/unRlDuZuGBfqU6fzzAcloHHfVAUqIq
c2s1M1PlhDeEijOBG1pxWhannqtDRjGD5D5wZjd++DChtEBWq/zj9IBT7LWpYSbU
g06WeilnqVeS18jyEKwrIbP+W/vb45eljzPwe3ew9CM0XkGLutA6r2Ms5Ftcnsmm
9jgCKg8XQNGd0X0m8gp0/k+Ae2ck3G2pFpv4fVE7voO2/LRaYk0+aOSVTt5fOm08
fcOPiSqa0Wupf/U3ONzJz3i0TzHHFg6qzU6O1XTf7mFF94o6wioVqUq0CuvWKOiJ
hU2CjolQrv0o0D+P3BVkeCaY/7hZlYKV14QfsirurM6GT59govxhIakV9d43Ei9Y
JTbPpIrrSCFJl66NInhgmXNnQJheWizkA3DwAwEdXmtDEYMqdK5/YwAUcbt5vAeH
1rCupy/RTrauBR+K9v/qKPkUVktzE0R13Y+1BmvMCstAv0tyNA/YOAVbfIJew8RI
9KFCJ2HIOCu6a2C/2yxcRx0jAYvyQ+58hDMe1IkFLT/7ITr7RfIqNaSMuqxw/8vO
tf+spZ609E1xMe2cyW5fXy1VP4/Rcyt2LTGwIEW1sGvMrogbSn2pKHd1pF5vM1nK
Md6sv7MY/vnKUAvzDAdwT1HKBbJZG6Rbb8Z5p30E/1ipJTFTnJEN5D7h2DnHymsh
Vi2kVKlD1hjCZoltIjK2zCeTfauj34ocE+86w+7FeVQQqO456ZoKSFZvExrGpPcd
YKba3AT18BqQBJhxrl0MQS9vxEFMY4pbB8fUbZm9qpnnJmcBHAkLgH8PSTqYsj8i
y60VqEeTuLa3q3VCrJjvB0ah6MipTUo2PitdOVtnPNdu63vKzlD+VAakmvXHzH3X
JmYz0b5YMp5Rc1wfRiDQaR0yunUU1WqgrbaLBMVFQpn6TVw9y0c4LEAod2j8FsPG
rO4gUFBE9aDUWKZRPwQuzmYNzHwJimIqLmntFkQwQ0TETcXnWyeg6QMyN/42Ofqv
6D859SyyN5ezuY34mtw8F7dKOL+gAzWQzOHtvainCJjVIA/Xw16woWC7xhydP7CQ
ueg5/9FeXC+tZj/T8sdBedcIvzSBVvFWl5n8T5hIYEkqc52My0ZDH8ehMlpoxhvb
GXLkRv6t/HrwD5qgRAZq2sO56aMaRMkmd6M4DBtdCl4QBZR3A4BlWoTgSdhI7tDe
4clLGgf5Cg19m4vjpbpHlJ2tKdSwEvxHOA3RgU59m1py31LNi/mUaXRSTEiCoynl
VQSkYs4pTV5eLmSLOYeUkO2ChPTvh33a6qFaOiumldgZ2telmf/SH/ENH14hNSwY
TeNW5J3qzfRJqe2i0ojoXSiVdqFsfZWdPJNj8uwnKRGw8istdBgH2t6dDdCIMZ0E
sfnwh7qUdpcpnxu1pNKQqtqL0zIppz0X+VndA0v7mqwVZ3aicOe0uYpPofqO1Jy+
vURL8ecXuaMNLk3AXs+XCGxB1xxzJiu46+D+LvDQKtyWFbIdYL70J/6ijlW94ADX
uXwWQgJ7K4rtuOwc5Y176UbeQo5k9oK2AWFPkD14fsGopeN5Uvfhlu9aIS4TAw4/
tnEMP+t/QWgtvWlkAP4alCcd72I1D7ATynRh+1j+4gFUH3W4sCgeqbhv7XkG0dCD
JAv9WBybSiCLd2OS8h9UGoYhfQuv8KuBuAsUiaVotRZd/fBDfmE7c2br1sKUiK6j
10fhRxN71x3bEK8B1c6NFjY17flYiTwbrmdKyXKU0LtihPEWn0d47NyJ/rrRsDHc
DcRIzsZeHBln1BpRxSbzCCpTx3YCG/mBvNoUbOXD5iU7cbaAATN/ZPGSMmHfSbyE
hijpNJOgH5bOlBraBpOaSeksdarawyJkqPEXQ6RYczqF0QuzlZwJj4dmKc2Iv1MW
LcOMCEEb1QZyUutVzV40HLRo81SMG/ffMqGRQnpCHoWMR2uHhWTi+tV9alGZQzts
hdeV1lwhyGlrqOwEiTJHucHDUSfjFFPwqhx9dfpcS2Jb+g2+HJ0pPvoc6oltePgr
K8KUxdggvgh8qlJSnZtPYti4tKIhsUPt2H2LxgGssgcgkStu//hL627OR/pF/fqf
z1LQhgaTxjA4hySqB2tIHeSw5yNL9F6sHjYbHV3Qs1MBC1HqPoJ5iip9mb12MGwO
A+pA2drCerJWdu4HxYfBeaJH5eUzraNb5rXRNAovOtTI2GuJ1rDih7ABadC+d3zU
w3/LIsdXP8ujo7XCLdXT9f5tC5HS0BZN/KuhoXJ+TjN067PJxhG9zCm2gzBJb2gL
0eGYifFfegf8UR2rByIW/rBD3RWZwNI4gKRO0R9yrRK8bi8BUNyZHWk8M2hnXMu7
D2gn4YpfPgQ7tGvs93Nw2/kNaIbz+oXGQf6OLLfC0hVp5OjXDhfs4yeTJMWTZ9r2
wBDbSWh8NtzxlixkB97Oux+Xb3kDGv8XV9viR4r7VA0pmAtWV7UyxknU/mUcvx4X
FarMUssCeF62H0ZZXXHAqo3+2weLHQlA7QvjFK6iP+BgH6JZH1vR+5V8Y8pRe9rc
ZlemGTlAHfUJ3QS76PUhBSW+AdiE4be3Vc22OR97gD4+PWxv4gYOVjtvkezNmD9R
XbI9rgF8ofkm9eu1zz1BWepxYnT8+vSBaUoOI+7UlwsZgcKwHWMLMOwSowIyjL6N
Oydddr1GzM0+fB0ldeWWLLGCyOwvLTp/GLvUQ/DmVkTk4FdH6imxOZsGZI0o8Dur
9xfKAhx3dwFmw9PATOXf6MdyAlJw86qfnYfSyStgYK0UBk0qJC+UoGoDiTAeqvca
17w3F0FxHkIIpUImPdoUT3afEWAjKu+ag3LkiuQC8jssR9fTmFXab53slxHprIm1
qH62jjpIbtVd/zlQnkgho1xpa+jcELiuvl1qRuuVaVmPwdAOXCMsPKGo+EosJ9zf
bNzvFSSPWrP4YvOI+5ivmkApeUaU8h0elsVJy6G+HUg+89gcyXisodzpQkRtVaJv
ZY7omTv0y/Jad8awJVvCqRK0tZfUDwku2Wgj538pX5upSUBmDvYNqZdz/lVx6WW4
LqO86aDiEL52M4xCIF94WKRzgux2U1D+kWVllj2E2NvsegT+pe5p0wLLK5w3+uMj
iTa8Q1kdG/jcb1QVNRN0lZo00M9cdrW899ySEVlGmIIt/Nur5PWZ20GFq6jsknWt
YGImYTDNiee4GACSHxnCoVsjsNejdu0UrlC59Twi6XKQYygghCYX740RXqOEYpKo
zy4hI+9kA/7CklUg8MQUkoKRSvmX6RYKsoOVqv5elftSKv+OI1zAiRiRpxApK5EJ
DtaGwnrlXXgFZgi/h2313KqFf6ZGDEnPu1PF6Wj9FiktfQxdGguEPkDtzUVVY8sQ
9ZVOwGoC8GnHPe8qGLjYb2g0to3ylE8lfeVOJZ1xR+N98SKhk/MQBVPaxBnvbJTb
yg/Sji3cvy5TIxiVXas793/fjQ9mSDvQZqcLiGS6N03K2y0a+sM1LF7/znnihjjs
Teea5Z+EIQk1w5XB2Lc6iGClOF8WSy2r62oEX3KW8JEpypwa+i6uoUo3cbG+mUUH
I0kGIuexQB0O3Hphdjdm71P8BCodX+6RVq4Vug41fXMnQGLOCUsAcK1aUaoEkpIZ
RlCkR5On8C8W2jUxH/yucTF4xKJwbyak0nQ5/MWJ3RRS92NDblTqf2qETpUsgKeO
2jKdk+uqLuueGzeMg1Z1IKSwL8YQ+G3+tBvAno/ixFYB89QPAINcMK/AXWs6oSla
cSJAszBdEtL5ejTCUJBt5LI689QgJmhi9YsvpD2jzRaf5R8K7ggW/q3Bgb4r9E+A
apwqVElll/UbdvJi5JwD57Pi4qmnhBMFK7GDoK8D8vRxBcq2uy+arU3vgtF6z7B6
4gZRugfV5+QGhDjp0vP1b7mjtZjZA0tOc9B403Iiu7Fn07DlYvgHHcLEV3F/lEZl
OcZ4NuJEUOgbuZ/ngxKrmXeRo1JezvU6Di2HwvFAdQq633gZdLJlLV35U3BajWgm
zpnLEAZgpPO5eEJfWmGBe0aW99eNfKAA3TkZSJTAz8T53q3p9R1sz3gTxoIylsaB
wfGX84oSP78+CAcIgcVLQ8J7Ao9M0v3Fkyz/XdxAsucF0GJVc/4Mn7IcDj4JpxDZ
0LxZ8lrHcJMGHKGprMuY0uLaPL3xu7Vb1th2QrzW1sF9Um+LgL0MbusvEZW8yJUV
SnOBZ3bm89KgXITy185JMlAyRvW1F9LyTjozmepGsH8PD+MJJFbUKtLvAcRhe3jV
QF1W+iA5nWaEPB23J8ccRyJvtVcRA8QOD9hBnV9pBOfcTyAprL9MFDL9B/Wc2oNU
oS0m4jx2gnD+fY7ncaUsBd4AsMAHk40zKsKkHg9qIBf7LzMsF87AwaXuqKuHPucu
vG40BFaUoVF6O2mahLSiNtRpkxsrAk5ooDq1BxVgrWPvkgt7piyHOqZ+m9iPfLSt
4zn8Bq3X85W/F23tv+2zVO+hijofLYFC6xpGcUd6BRESDJlNVAhMG+zvSadBQpPe
Osn1V9s40eqqeVNY+DHSOmWvFv4j7oU4CO57W34nREFydPwoATVRltVEZw4Y6YgM
b1fI+aGIEVylWn4ky8yBXjdsVVWex9eNFtQWCT3ue3GHHkmHd9+fUPX3DH4ya4QJ
uOiuAHgOYhcbUhw88KYzz0qQfnjwKgtruOTdCtaH1QtXz0/PWNrMdbqggL6tAh7k
FdE+FKkQVboOpPDSITqVNfLLFaUc9l7reMrWl2/fUR+Gk4/g12QDCHdvpj9oREbe
D675Edn15ujAi+zeO3I82wkufSVNLaQg75E3Alt1hGvIZu0vY77AOsER2KIrev1w
YlTrSHT45zvcZYLV1aDPL5upXf6DvCadrhRLTjOfhHjto64IdSruq7YCkaxmq84e
5jdSJ5OgHQ0iIsS+yx+ZPpH/IC+fmoJuU37x9JC9tpoaUvScZaRYHlGKUaCHgUgT
AZNYptyrTIxx0eebB00AKHTnYI8gpxVgiePXoNeYWnujfn9REpLwvwQlkgWY/eKB
z8zdco14BIrAllUluXWqVxRNdJyoITP486O869CLpxPLENOxJg8IOL493wwjpVx+
wrhG4rEmIFedKDATNuIesmw1lq9uOVBjBz5mIbiT5nrfaVYd5BIf6MLPcgyTVDSO
IMpn98dehlUhXLatAkKZ94mg6WbGwalRWj+dZnHnWV2wzzpzORLX1IV9pU/9yY25
hWIgoxd9dbQ1nloAcIYcUda8vNhK/rZdxSbINsI+LrCa0LVSIBPdOoY9kA+Mwstg
a/5JEYZ9i5nJQ+/JQVWpnsir3n/M3ezIc/NNOVC61jjWHIyYJvMUcf3nbuDxS46g
8ABgUI6r+ZV6WAiUpZ7r8LlvWdxI7zrRXOFpn0mpQISXcq2oTqvoOYwXKNg2UfX0
BaJ/QJxQjrKeJ/nuHIXeDB86oHtGTU81N2TDeMjFUsJvBEPv6MrV8BaDtM9kt2jE
zNhUa7Xb2v/1v7Z3giG386H7Y1WmTtJZvOK2jXCs8pUHXKvwvBZIcj7E33/Y90Ud
svSYkixz0T7yapG+GO/aCrigOqb8t992SgXlb5VVm1kYpjiwacp7YVtAHva5loxt
zBUDTJ+y6c3tLlppuj4AgxG86rCexHyQeZ8gvWOP82rHC5yV0cf1h+wS0oGnlQ3R
5RH8GX9HS2Tk3efj2DKcfZTA4wCV0g5aqs3Lmm6kHc99+tCnkqCAQyVqa2SSi9Ee
89SWA3HfTGzF0C7OJSAnIVpRM/S5BO1wFqQJWHVgUQZzbkUId3qViBBPthrFj5ZI
HnxHO3vK/a8tvC88V+SWI0Jur0B2iE0XV9IJbQVt+ltXRgq4TN19uCLOUPp9LlRc
U2jmBfC4IxBuIEgmCYNzKI8V5OKT2ZH+mhCnIXM45m002beyl8ZE/UrRxkMZtCmu
Gzy6hVQWXxop/WN5RCrsQwjuhHHkSE27QW8x+SX5OF+21VBrgxtMerE9BEQwOE1B
0G6cR5jSL0UGa9nYFOvu/h16AaY3tn6Vjzk44H7bDB6ma/0N3IdpemhN/E+eLr5W
rIPiZ/Rjo+aI5KvUofiVc+LxZbY4ypcKhKf7gIImshtbEUh7/zgxLi1gwTQu9L5K
qcwqc+DzjRBv4E29vXLatAt4HHm1c4Tb3/4CtWgXknPVnpmdsEOekcpY1+7oHnWg
+4qD2SAwV5q66gfbPRh3Q8TWj8lZtp/blaf+DQlHTc3cBSDVLVvS+PBHmDQMjGnO
IbigzQyjcwlPncMVYMBeKkR9t4tzxrulfCLyzgbwivTI3gDwdV82hnnfrFcxW/uc
2V3LMuTeZYDOXFcTJpueWLJqCfFA4UpQQtpXmOvYH/1K2dpVnZTbqlK6YjjcXYxz
uDBzyMcgfH0W0gM2h5QDx+/QiFzHcODzpPUV7cjo8s9vPOn+/r+3H8HVCMLB6Rrs
J2mEz55b8q7FSubFFuY6gh7/BPik0+hCYvMs4pHkZ6kgK2qkKQlW7SXNGFvDOzZn
jdw10Oclc4CCM6YA/wt5EIi7NPU3U8G4LzOmnmQEr04Kgwzj/Eu3Va+g2dc3BtqT
M9HZ7n6ah0RvWrTFDKB7WRmz2IJG9W7P1M1oHcrRnMHq1B3Jl5fr+3rWr6tQ1e4a
pVaMOF4+NtAirNKH/yvTi7MEwv0Az40V3fpBQZt+Qp/b6xrGkzUjlBSGa4IAV6sK
ilczZWBaqa7NHCq52BYejdvoyFy1n7cjsdtamqOvOC+lKyuA1fSzGyogbwX86fCX
FDDgFHXx1+WxJqcbNNSRt+UA4SRsNK5+Mgo0Ku8uYvj671B16n2Zjg2jepBevdVn
luF8MQazEGGjZd7w+dmp57gFL2ZORTdcfJsGckxsNwxbamIBMV53k+pOPzGZwPy9
20ijlt2Qd4lb4BU2vC5l6J9a4xGLlI2J+4Iz8JbXA8vttAQMInW31XWlsP/Upkfu
bOgGZRxsBGWUEHHLykb4jKD02FizemOqpaueMxjR8G3mw3Q6l+P65KZ/RnSLoyBB
HtVTI3xrkf+THuR6Huh5eVTm+zYbxVbw4aGIW+ToGXTskJk4LXIkNbUHamCxh9K/
zFpKWd6AOOu+qW83O4czh2E+Xb+ovcvxX3Z3UquM4K0NqiGAbpVywriHK5AhtHT9
Hi1izylUTd9L5zE96Pn+qZYhoyWHH72TWNaLDyvmqo4jLZNK3u01pxAwe+PfFKnO
DrXpvx9Qd70i2TsL0SZuVhul5LPwkep8LtQWjFE4iWwzj2VGElu2eRfHlPKcWOvX
tznmYbDEEXgcKJSK9v9LtmoBTJ/1jRnR7808ir32BC7SwGGf+kGUzimScp2VVQW0
Vh+obEwdp6KKp0aS1cLEyqaiKzqLrSLOtX3mdE5PKAF9a2Ipv1GHkJzNdxbVJ2lI
FGB6yKJfbPgvWgO/8ZqcZt5RjDPzw/7FSat74EfSs0N1GeWItLXW6H45wEp9H0uL
wKnXogF5jmM9jBEdA6YIBepogHyLksF3aEShUyVJJ0cIXqMy3APvAvWcUKmwWhrY
8bQU49tamqrp2bIHEYU6iVhruVPjaxlwlrGzfRNn5bEA7FDmwLcZg0nOccIkadgE
QQgveL7ALVuukr1drpnSnKsdcRzq62wtb1LxvsJ7OxAWmjVlvKmWGNjMXDvOZRbu
+T/tiTjBhfrQI/g93WLr/rnffl3aoL+FJXZmBlE3TB2kuVIBguIaVx71/YgskHFz
EjlVFs2fxrUG7Bq24OwiKFTQzeXclC2QJwqlg9jSxqKBniqVRVMEdg5faMTxkcey
MmiK9okW11iBiLTYnWQJM8fxpS1LZjNO9aVc9S94PI5yYySzBDbRFwd7McLxtarv
yuJchb9IR4L+EE00d5x/G4zDtMgkW2zClyj+HHlfQBY3ByIIld6FX+6QEB7azEd1
1jJOpibGsa0pGhE0HbflOjBx15v8axkaGxpOKKGbgOaxOSCY0HKP6frFmttayGqO
H7JblOn6b31rK4t7LtYm6q/NIMVUM2E7mFhuCrYG4iZitMLzG8mZpHjfI8GVg3NR
i0Vt9TTjM2NHc7g5Wnw5YcSNNLiq7ujbFa+KDL/Peszlpaq6hnFtvBmCB5sjMNg3
Lhecj0z4eBsylvdxurFIs49NhwHYFJs4Q3AwPAaQcCLRoCOnZ39j2A4xKFOQzem2
29aTLkPqSNa5OFjPW8XqfQrhNFtqKSMGAXv0cRuynIvER7BR4VRb3+vAXpJhpTxF
+g/1rIPcHJpHv2NIRDhaOCEmHfiMNrOFThdOeFLZYj11giTU9jdBQQInSbPMa+c4
PQmr+I+jvsZIEXjM6oKH9G/IFMHPdx0BSFxiEhg04SKsqGRCLDhxQbHjr2AMqj3r
DAT88O8MxGykaQLSMzNNSS19Norxiwp1Phvj5hNRaWIPEraaivNE6F3KlpjZ0Y1a
f1R9WKz2m2JfH7UUR6ZByPdsfrQsyirMjiJ+/z6i5lUgwSjvLg5ZBC3UpPR5duqN
3T9dAP8fofy8YpGWhGlEeFKkt966vsW/oBYbtBuvDm8S5q+LLwB7fi90gJ9SgIOs
xl13/ydbEu7grWrSwg4P4963Skd/kKXk/6SgIjso4ul1dkFD/Jc2eVKnANhjd+Ge
uMBmpDZvjGf0R6icMkn/YflJ7ESM7Ou3VQMbXErRwhNPJTRepmHVorRF2BXgXiaL
uIu3hXNLFrQImCGY/r6f8Kg7ehBcNOBN3flFiKMBV0/6dQnbCoDk8++ei2ST7kTi
2TI8zkV4Vl1b8VfSHOx9HzDvErjWBKnYSxCWyGidmdrCppVYkhTtB076BjFIE5+5
weg+19HNyoE3THSA/x/Y+aE0Z+oHUfN9zT+WOOqCF0JZYO3OaYHnJdM81SkwSKwY
1jFEhFRAu8G4eEbhF6VYPF6Q8uTnpaKteThV0hKoPT5m6GHZObDmVt3u1Auwj2Q5
aAuoT15DdF5JbHWEHnHkSwJcTT7NVzx2780blRYlnirZNQ+SgKn0JFr9w+m5nGGd
CFAPXq0Ow9B5AQxHKEnjXeNiHpmJKREGSVhqvUg8axGrUl+Pu4lygQdf5Q0apf+9
fiJ8MHIFuxpP+MoHnvw6lnpoFw6LJd6hmVDKYU0Sljy1knvdqsAJHsXc6ZpA9oU4
qSAnNtZDlsgK4vmaDqVKPhWdcaC6jFNsr1sZg9FJ7BugojnbkGf8AxC5tOoFm/UV
Pla+GWQJF7tedb9j+H1MTUSHbASmoamNOkkfXWIQZ6tImjYNm/KXe7rB/v6U3Hkz
+tz7K3En0BUkrqt7yYa3JFzSdC5uX2azXBMfKrWtPAqFyzjH7/17IS8pAtRKvB4n
7mkzPgIVIN5NS72pjF6gqrJArSdOluylZGekLM28UC02E0tDvqLFM7dELK5YVKFY
O8VKD4fIUDFM9GLW5ce7Q0U1E+6RJemTCQR1GmnoBPd2nG6rd874wmfJOIeyUjmy
nLWD7OaTSDxG4fyC6oaONYs9yLzkVi8QvwY23XjEBAhhn2rYkNZsQaq4HpZ8oSua
0YIF+MFnc0+RiAmmDHR+NwnrPI/sj1hGGdWmYopO57K9LpvIUsdU8tyr8xDZV7dP
ePk1VFNlifSZZbiafuN/7iCGZsk4/wuSMAy64FO/LKU0dZtunA4N+Uy+9TczXClJ
JRPoxVWhCfCC9EcdCPQ3ZpjRwt9bq3dT5GaWVi2mLn/A6eEQDzYtWMbQyMk9A+EH
DKrFjd+P5uwuI3ZJKsr/J0cs5MopbnA7myj/5u7tGzm7QnW0kaWB2rS65CbMClzO
Rg/Pg1iCErTF+sTp6RMFD1JphJ973voaDJth3hIsGwGrFY71mOzLd0jhcr2T3f+F
iC4chRYHcYYdv5l3VX3aWUngVUbPTEEniXzjQQZOp3ueNfKtFvUXnAhC4pec1b4f
m6s+NTM1THw3/0nFbm7KNlPlEZDvU3LnCKUq5ySks+RJMofvNQWQNexEP+D5QYYd
7/CPrkgdqv9F2cVLkxnecqRDGEkez7VUp2T4Lkg6nBti33aVm5yPV9s/3aCdUwb4
e7YM53xkG9in+aUE8pm1T3uPjeGBXnUY7kPjDnEDdU88vIhe+SaBp59V9TnZ2hSo
s6ur/ftlpNXm7dcbnRvyu0DLyFmHh6kWmAqAJj+RGTwx9/l/bUg1MDsT1/udCZV8
R1MDSfi9RJH6vpwvF/9/Ws5utDesdC0WcnaZFyg/9IR9vKFtlC/Ooxxm9hLcZW6Q
rHVDG6SiT4+MKZJChbJKwS8f/7W3LiHNk3PbEjeppMYW8qS5Ai/108tuUYOueCWe
ig9F3p00kMCdopmEXxJmrMf68CppnRtbX1esFdne2udEA8kvRqWDEoam1OFi+kn7
9wnxpglLFVwsB8Kdak1sIity0Y7dhWG9/8TRtK5gF7zr3Vgt1mKicChwv8kWqbsL
0006E+YDOXkoAXUFneLyiDZNDP3yrKLFi+g5IMMcTvB7LdKXg0hHzRlWzKaTa+rO
ZJGLQx2DFOCwVapZSfJRY1gGhScw3aIDYzVlw7T9MrJCFkL+A8lkWSfzTjjpqAiw
VY1XXnRxtiF7y5oW+5D5bNp7ZajeQyaAu6rSEo+NAR2Wdl1W6g4srBD6BK1HD0Oy
wKHtyStf61q37yCMUJHXshVoMGf0Kbi8SC5jL5aU3eKyDKJ3fUk7bBj7Fdv5Oxgz
f+5BXnFAjEKFJ+J2UXOWjUYmJw0cSagiRrmZRXowKQhRvlbXoiLOd0cghIWOw60D
1WDPtzCL9GLy1jKCelcF1M2wPgDXd+mNYa6N2wHyQAaLCg6DlRIbCaqqduFeMm8H
YvwEH7jCCkeXDX/8bXi0/7cNqHE9wGrlm79IqtCYRZTzHoNQanO3Ckke2wWEwdMp
WtrtbPhuwvseArqIvGjc1NgjsG85br+EF2Ka+SdMWOF70wWGqTZdSVFPq5Tphdov
ytSAIvxzJy8OPw9qhQNhul4FPrt5PR/ZnTyPQU8IsBlxYofb1AIKBNQ1xCgb+ipv
f++yCIHgDtm9k7pm2OGfyb26tyM9GMkcd/fHtoLUjtNNvmKbjO0pVzzjvuZ/1w67
61Z18IORvDCyAfn3k4fzNispwT23LTygm3cytNjep0DYCGdjcECIsLfB87SorSpW
KsNOHCG8G2t05rzEtUoVGtt7KrCWJyl2YR/ksi5kuRAB5D9hJoBVY/ahYOIY7iPQ
n0Rko4G/+pz1MYMiOXu68lD3c2pfdj9TlZe/2gIeWHRaf2a5b5pLqY0XTYo3hh7I
wJIQ7bTFbMLOshqJ8d+JuY3deecQlCI1xSXijKBlM93GtywepMBY5fMNfMQjQGHC
TXB2+DHGy50uqukrruWzomiGV3aZ8Mc86vnaLSn+6poLTgky6VD2J1sIKNyPI/2J
Ayt1NHri30VJo97G4wk4OSo7kocESrOv3+c12EePiKZYHDQGAaT0Y8xT7o+Dp7Xu
lErBEdcIgIS8WOA7ihAbDocLxcmUw1JjRPJ3vKtJNaEcNx2wyLqTm/4PyDPB7iET
tYsgu6UL8FKVlxOEwveJmspt6b5nUTQy1WjkbmD/rQZjJqXJri4lWr/yJygBRpKB
mR38vAradJt4z7AeqoSTPfApaIlZG1nsvD0cT3o1mYWzGIG3yJku6ZjXFLtBxLlR
zaGbioaQLDa3h6R8XnrAxV117eGrU8vMmxE71G9iO9jhGqKJLs0NvSht8LsesiEI
TmAqxPWzveot6youaKVvfe2ms9j7NT9CFtcZWg0FWYzcfpKypud0bIXW6wQWe++J
4qrVUV7u2EvEDpJ3W66X+nJ/hyLkeHVKmXmOhArPggJRQsAcmblBjlvXbo/4PO7y
dPkS4JbeMooVQwMeMQw9q9GSSajOc1CSAvwSZzSjfAPiu/Mi+pL4DKWpUP9eIvEG
Xf1ifS0Q3dVJuniLVcGJzdyuegHT/mzIr9b0Fjk36sXNoJpIzp1s5hV2KJV2H6G3
XiVcyt8SkhQId9mxisgRsC0EJGIdK1txMedCpBtagxFooil3r3UHDKHv5mJWlw6s
VrpAuU0a85S67DAj5LaQw9sFg1yA0Y2gNA/hZ6Ay+kKIgod6lay2NUiq/9yfCCq3
ir9ynbBXhxHHiRY7eFRkp2mWRPxKZotvaOxnp3lsVWv9XC6wMp2GZhUAFlmxVGSK
ebA6cxsg6cBQd8aMIjVQErzUQq/zwxpEojYux6TtX9rYhCVVH3L2F+a9LBgO4wz0
A0352IEWbR9ksgmr13IP9FBGVXHzoUXIM1QLuJiZNc59WbVxijAx7+F2+UNG9IfL
ZiZwqi0TMuY430p0YxrxzCZU6ji+B2amyWWHOxL899QV8CSV7k67z5/8ULEWqvvw
VkaXf/Cm6iO3hXnxlr+6PfLFmTH5obZ+nExfghU7owAGTSaf5i/sMuhdAbDmQRXi
0EIL6yqpGlLbt8bfxyK6hr7OchU/IPYcO9ZraasWArcYGBfvu57hC+pZQ55XBC1B
R6OUGKKsFmoJF+276NhcJoZg3jvPDyKQ6V3Z2Gl6IjXjOfLcusYUU2hwCc7cwdiv
9S3kj81qYmQnTV7BHIMJx+cbPEv5iM3aGjBM4cFbgBc4bYStNbL0KOpf1BSfUDoe
Z3Hp3R/6mLnRsGS5OZ/yzZlRBG4rSNQ1gGvA+ZaMZ8N6FJ7n09Ty6TsLUwRcN5Fc
0M2Ipy5sjygZYXUdDQuFiK5LchL76/30RpH/etUaYBK9RcsgCzkH9h/lTi+XFEbw
8Mw0jfH6RCpTIhmrHsT1yy6kzrK1kiYVVJYmFWrYyQsQB0ARmRTCkUc5LvE2aSd+
mabRJMiIVEe8+/3rIjfk8kiNoHZhhNI9b29fOdEjUOklGmFapX40rZBWMvxbk3Yf
zTESHnHEuBsUwsZKkmvunINgAz6lEZp4YmO4wrEsOm3Gh2X7FHQgsk58J+jqcMWc
B7XaftzIqaWES15lNm6YkOJoRpNBu9VCE7SttEplFiLF9L2tDkSmzhEKbU5XKk3y
gb6jSoSZDmCuhreNK31iR7yfGCNyrN7VpSwLjCb6g9UF5XEAX/jvIqc/ZEdAsRnv
hDptyGkBC9VSdJVVT9WgSnEsf+lk3JHh/K+cGCMrlyEszFFG4JniwQTDVx/yWZUc
DxftJ/2Nv1/bO5nGpapY99K1x8xtQAwUVblFhOVtzJHDc0H2C5NrG0xR+mxoua0f
+T2X9goKyZTZbJw1nOjt7NhWWGgeHL74JiL5peIq/ARtkQP8bt8ZAxiTO9rEEV6R
QjcBLIBhJw+Qg2adIZ2S5T2Jri5sTIYLN3ezpX7+tZsOooVdYVN34n8jxAyl+jDY
Wq4X26iFLxY4Ai2JPquK2ewrfki6LzAKPMPKY1pI6bXZqcMCvECcivGZUPlzXZIX
PbpHK9hsxuJSHYwhBG67Rp3wzxF7cUxhvHHPFE22n/djQBnViPxkQ4uq4/ZRv/8M
SO6PRws9hhvuUix6ca+L/LIwKp4fYOQPOHGWRNfySOBXZjlg3viCKrKQn9rbwDt6
cTpS7Q0TOfqYgXZjFQkBX3OxFSWHxkLfU/OSGNPQYebF9jUY9om4XeTjfrZfbQaZ
vdna998wfhFihZkmeUW5peFSxSvDmHlxMSLgx0amJNu0nPYTv1FmpIRgKDYfCU7Y
e+dLk9c2v6Gyp21ncVs+vHzZ2pcEwKTKLCg4vgS+7AgngZ7OUDOalZWYw7kA277G
xkrmpjhhpaIk3CRhRCUdc2uqMiWVGKQ2fcfdTb4LKBQ4l+rnhnKSWScWkaLR489i
t4p9keYEFyjaKci9FYwYSSizTfDD4e1Nu1CDbxR6bLPei1eTcGkmXdXYq9GR2JSu
e344VYB/bxUE25cDNsWpLXwlS4MxyxUz1kjc7d4nFogTYHHczxaYG+koLxtWYYnG
SvUJLReA1ILNpa+gODjUj5QatTjHcX37QzRDuoHUIZHYYPauazXj5rtXZe3fYwyR
Dg20jrFiZrI1ZMZ3arStcXYcLC1Viax2AEY917fD1k0n5YQfGkGTSDCOM/vbu/xh
Uv+PCboNqfdqyUK4eCAV2bLmVZcEvGSX5wiLWZmTg8B0BJkj2Q8CUS/dSZf/EK8s
j4KG/I2xl0qworU+qBJIJoj1SW//VZ3jX19InGpu5FtQ7jAOcj8oHAkYsfe8B392
azf/Fd4L6z5MtP7HR9+Rq9FnVS7TDT6gsdUOW3tqer14Y0izOC80IpQ5ZkqBRP7M
rZTCTEpyxLNAjsJ50T0uDl9Mh1KpJeku9DNqwolmQG6gzSZumu7lwMwOJBCJl27E
My0cBLzXojeK17Q4Pv8PC8lZ8LgYnHfxNXj21NhCJcllP0kOGmjPLHZphJwe4hoU
K7EgjBTEG2bq76hKkp0HHzZJ7xYLJg4PuF/ai8ruk47Pj2hqYc7nFtp9ClaM1ocj
TzchdXEMw2l2qPEvWiwm4TbSC86wpNdDHBqx0KtTh01v5Tnf2s9Xn0uRC7eou5yS
jLV7M8+4AkVQJ0LUTm6ALXM//B9zGzdNpXF8R6duIzb1DnFqoqOenTPorBVk/fzi
ICvPx8nuAXZPiQ2jaRxUt2Du3BJNZV/zxm4o2OIOOKSeQGi8b9eYR0NH2wVPXXre
ukLAnxi15GRrwn9LFIHWocObsl0ZNXW3cODJ1mSews8pQdl0q0zdSI18xtAYFSzo
k3hp8+thBKxZK1aUDHo/IYqvUBtlsQjXi3kVOZbtUiBOrpQCouwi2AUPegPxYdOc
8tI2Gf8QTjXShPZUTQJ/95X7j0proswruBtVkFcYzjaRW7xWMbDApcHeqanGW+CA
cA8vaABaan278wys1NZZzdFy/tdd/6x1SMy/9ZtgUSYDEi6rONtN6WM5ILelVlqU
fxHZnxmpFFHyux3QyDT9rNwA8lQY9DLiAu40KMSOyfx1gM0lTz081M4+RN2ApjPX
9MBLh0pPS2VTpFYMzdw+oeVpnplGHuwCMBuLLIjZD2tfEEwnoVsPHbmuuO6B34V+
T88nRsSzl35cb1kZ6RqN+cR3nbtXZzmH7WMhsdLgy+4LhOvkXV8gaWqqxHjAQrwx
BCgPWo0TmzsZce1VoO3MW0C6JkvES1xEGDXYhBMyu87uPx6Qu9SEX+5d51wg2Dn3
tjydDbZqarlaYm3IuSZtPGNDgNGiZRbL1wcHdx3SkLWS3JSjjBNc3GYVCN4LVsXm
uPR4wCSv8KzOoGp9CwussT7VgfQIVnmzDbWHxGXYOuNlxwEoKK5hSN7TkYwjDwwy
G3/mkuWEkSpqmiy+KTmeL2LMmEW7h8hq8f0piT5wOqKImVfwlVJ9agzP5/s1T0kn
aM6iK847Xo845s09A8fHwar/yU5W01z00O3zzA7hRn7E8XkKIH6aH25ynkMeXNv4
05Psn3Uo2bua1QHwqXcrcN0figdvxz17bpk6kH+390fFp/xTSxshDeyjTtnMoQOH
NuWwG+DbInYawOBMGL7bSpjMb/CGaTYzkdzzlLrzj3G0axSbHuP2791xavFsccyd
p5fK+8cjGZhHcSKY6zEc+g26hLA2a3RqZAyYg++Uq+FXvody3gFBUqBDIW5s/2g2
wW1ptuASDy9ICz6W6M0+Im+eX4XIKFdAG1fJOgz/JWT5WYYcaxg+XWeBu3lGicpf
/bf6DvMV2LRXgmaeS8oeH6gL3+oPpFsFUbXuiYsPXNYnnzWNakbbT1Gy257KkiPB
NLgkqFqLWjcozHZlDli/cyghm81GUwuOIXYkvVapUkTIENdDWi6tqE1eFhXoA/Gm
Fy+J6wiFWknMyGP7QFuKMHgBmU4mxfkDxvCkEqIib5XFGCSAY98HEJaWUiTHazPQ
R9jnRoHLVqlgc4eiLmhd8fF8DE2Df1KW3Fs97J7BKiGuHX4UyOfhHPrINBoR6jID
n5mpOoW2ksqKtX1yi2M82V0Q326DYsnYJEhXqX6+0p3E13B0HPWo8JzWHRJtq4hG
wwtb/ESuIIBRicoBIaThokG3nMm82dNf4HayuDtnXfJiqgpUlg54CJZkQZFQBjpR
h7ge1Q5yl/24n95xGuxH2zlYyVZf+heVie6JHm+6H2drzM4AKPDQd52qtVfNExdu
Uw4pv8O+IsCuNO0UAOUkdhHv+J1yc/sMLpZohOUbIyysmUmkIn27scfXG5A3ozBh
yDwBDizNHwqFkmaREfxyBfNtBKTb4r6UrFFz0RyKIOsb22Fwv+DR97wRezQ6Lm1X
MY70AwcedTt3ZAmbJf8KmpWwMCTvSdi6U8vkF0Hj9dJ0abqlaacMy6CTy0XKh7ND
wphCNDP44HOHV1fmJfC3TOOpydVodO/7v2TvnVDhgPewB/Ksfkl09jG5ApX+UMOm
H48a4LOr6zojO6cUcnbnaVsTcZrZXFrmOo9HINgwu8EmrLbhtym9XfAb0I1DT0WM
cjlrvCm0FYzEa63DgaCSzANnqBvhqMEgbIrzay3no6B2T7n4nE7hWQC1gR7sr2pz
q7rc9Zsqr2BFbDb/HHaC66oG8m3kbCRIJKoBrhnkBlKmGqkWzd9DHQV7CQMbObB4
CzZg0vuFPQQAoGo9ojZ6F1M3WRxDJWSD68hsqZuMQkci1GfiRO3thZ3cYI0Pg94E
BqdzmaLofQVKMIPyg9+D1Pl6/CNhqGbJBGq3ESG7lQYMlrix8zXEffRG+GY8BrSh
zPhzFfFzJ7BBNDIkAltx7i+1Kx6cnqrIvubAFNBRLcr3GiB7Irw9TYF6L3IwFwq3
iEUZ+enVXKlgK6mGyrxWHlijUBlfbAIQKvWcv7/bq8N+d1wAJ61qff5Ju8sJWhAk
gnQKUOnCadVdgDo/w4EZ/n4cL//N9DsD1lERZuqhEQM/ETZq60pqJP6gTgrYb3k8
1lMQGQxU2x8Y7NNvN4o2UCHDwUs9FzO3XGTGv1GkKCco2V+g4MIuh5Re/mz8T/Vg
oTuoVVQT/CPbtVzWlid6Uh6wMLJ2VVeEzGYeYC8oF3Qv1fqFomYhSqXLE+CWatqH
F/qu+ITfdkj5JL8a0niM3MWim1v1+kJQNYxGi0oyJEI/+p3ILtSm3CMvkG6gWqHg
YEV4BC1QK2WqP6g/xOocSUsbqQE5hj64wz7OYRDvmi/NHSJ2FpOJRtZ+g+9ogK8p
ekbEXn59GBDm692h4dPbbMKYZJaPUfSIHkmqDoH51NJihJfrxjiH63DKQQegnPRo
QHLXVXarH48oQ5Zf/DCYa9GSsnvoYx4PLyweSTQicYuZAxA3ktWZMnyM1Et+QnHM
wOLuPCEj4muJ3FvlrHxNtl/m8t6Ci0840jtgfkLUQ7z7FdjBljLPWOdpBs0GZO3q
DZbJfdYvf8oktN61lgEk95CywGdWPW7fD+zG1GJBix3DMn/VW7PlUpKSgEFFLTTh
q5ClWcvQHXD9NZpLCYo2EVGjqYLrJfRiWEtkkwrjYOCJ6y96DMq0kkvcKVAB0A/X
Vqh3OShPbjdQyg53KUXeLFgzxBCLLnHMI7Ba6L7zQBSY5/dxrrdWFGWEehe8xcJc
eZamsZZlA3J7g28tfAPxWD0dzviGJdJK73EeM/G/5gJGZEr2rn0fFpNe4Lua8knd
VF/zPu11hL+/F7+cE3SN9b3BlIVNCBi6WgQl6Fh26FriUYKA0w9ag7a0/0rQXw6/
VtNlmQqer8m5sCio8rAJarNogPNB3/e7WcAB8g+kftkqNpWnCQdIXM33iDSN12Gg
7eHgjDPjYTyjKfjujURU368SW+p7apgQ6kmVtaIQZ3LnFzLyrfnl2uzJOBOrWlLn
XbnUbHFne8ZQZ88mhxAuDl03HbfLOAZR9C6Bxj85UTM5XL2QAeVOwLfQhbPxlgap
+zay3DPrZeNExNRKE4iTlXYQYULwKsCbd15STKwc4t+DszyI5sZBL0UWiwUYwmPf
E+EeyoKfyyfr4BojriqzJ9Q7Qm8KErrzQIPRwCC/vcN2fPdiKFp/eD+z6bdkoir5
mUqeaKAO2eOJjPjP5cWsLPQPMazQWOgKLOcL6FpQLUZJ0K3i/BDTD4XqiOgKx8MX
/q2ScsrJNEBi7XtUu3q97ZgtnM36Qua905UdRkI328gGgWueTeY2FAJj9IoJCYUK
a05w+EjBzBNbSW9nzjhwDckwFubUtMahzSfXQPAGXZslXGVwC6pdHMYi5DOl4zIq
voAsxGWQ9q+4u9GBzgukXNFAfYdAxLipN5bnmxgw9YLWoL/35tQXJlPPDXiV8Ex4
y9imV9OU4stMLC3Z3ZLIxesNDqCuEbohI9akI+gAzLjRpG2IiZU/s9lgSKGVbMX9
Pt1qmuwaRQv++n3T/V06xtKYWCEDPvE1VjyTO1JwSe9Puw8Kdw315jD9vR0DYF6o
l6pyS9FDzyyTjwIFlaXfJfun5iOJGVqtFZ8XJBIamRhGEHARULMwLvxloLRXNV+a
6DftH+CT5+/knDBBNdg7LNsczSbwx4DRJzz9iy6yG3fXz1djujrcpmkk1oeHg3eU
cvZycw8xUG7a7i+cXyp8Z0/N60uRngv361xrAlhqb/p8u3PFIqgZpfIjNPCpVsvm
xFp8h8UQgmye+Nsu931d316z9lDAZnyzCNyvGkaHoPfsSVRF5e8RQFmmoiLYKLSY
vCq3/LyXKJUNzATWH+Whl7Pr91a5j7jeyVKZKqIydXCqYVHqYubMeCruZQBp88Ds
I//r73czj5wk9lji3qn7cA1dm47zV4NxIX4FmNchYQiGhq50PoKEBN+hxnzhGG7P
V45US2OeOk+ivf1ZNLE9HD4RNRIzR4WsOhzxVeGt9RyQYEn97bH7v7OrWwX5arnV
APqIyKJXtx0IUCAIyKyIB2L2rDp/SDIknLNFKcMJ5RyWfuIyO5mJlQO++lb+ov08
rQvYYBB5e5b2c+7M17AdNkw/lyP+OUSmSufBPdwcdImhEQ9IqYdPgK2BZRjWal7a
rSJT7QNBd2kp6g1yGU+H7n17i4Qy9812NOkguJfsOtuWTEdFAOPQaMSEYG/4GdUZ
vwF5O0u1fsZ7doyAzRo6efi6QwtuaTlYgP8jF1/m8ljC5Ug6NI2Vsj1uHh6nT0mU
/whTpEsL6BpFep3e9tAoLpjnqpe1vDmm9A1N1BkT/0bO8S/nYkrDJRtG0nPdwKLO
47i4dBy53TG4+zUeI3zCS3zjNX9I9bcbbrn9HDmuCkQ1K+sjRqjOpPXtHf5qDdl/
z8RpfwNiTHknVi3bR4wSfno7Rtu00xYRB5/WD+1PHRuNIiHdKPX3lOgVgBMlDTkE
NgX8H+eVWY5AF2jC7IFuIM35QEMgo62vZEqwVM8/rDhYun9Xolvc5+V2NlNS7fB6
NnG6VG9AjpDN/cug5CCtBAlmZW+qc+L7SfVeGAIdqMDYJdjrY0fwaR6QwU2uS9zt
FYw6ycDLa3dJN9uHveX5p4gV10dOf6nh+N98TtcSvz/EfkMBhSCdt/KDAqxq4z41
tcqNXZmluxWYRqnU9NjnoGmJqYWVa4rEZIFwvUAO8ONV3O9B2GF/u+pUS/LMMipr
HQRR91jIfhSApa9hTwvQYs+apoT6XsD83b6F/jvwZM4742Gxs/9It/UE7lT/u6as
DlCUB5jNEKAuoiXNmxG1nprePQZ8RuJtCsp5hPJKfe0VZ2B7fl2K0uHYjNQOWZvy
ms7GZxG1hyhDNTAxGIaJ2KvOelhXmMmUjFGBWx+r/ZgINjT3QvsQJSIFV19aQEa9
jieoWz6upFP5xkrcdLgOKxRQakfRug3o82LXJclvQRV7vh1HOHFViOKTL/rkdydV
bH1DWmrg50gUFdIZioiu9i8JpkWWq5o1ve0fAjfkNMUP5+1rT+DMVNjTD6i4DCUw
N+HXs2Moon+pL1f2E1AJ+pBc6b0Sf7mnyosLugVEH+loH5xVwM0RXQwPzWLAEyIY
Of2Yx61vNkrvcZoD6v6ccJ9CGBqtUCj3u9cGS+c+lFY0fQ4e27M0GoQPrlmJTElM
81H1AdcEJKmAV7BKlueVThd/kVDWgh6C7+tX5eIjouJxSLYqaVhmS28sMPJvSQ0K
IrcFT9EI+OcB3xEWsWiBeL5+sUawSFQDLM+IC0CUCJj1ZHtm+D85hA64xoF0m/ET
1QhTrloOlbCEWNuSljHaHsU+2WANlO/hh756tPXxu8XvsGgzYUcv4HO+BR3wm4pr
5gMVQvjIe0WaY2eI+TFfnzwwHfL/RqRI76YKI3y7NqeFWsOixqYJaf6bl/avUXPh
ekMlNBjbdNg6mj3KCaM2mWRCkpo+EptRlBk6q6CRcm3nF/6XjuXPxoyzOKCtJs/y
Vcijcen5KMw4vLAAQ4i/VNmltzzqzfB09/RZNk8hXV4ioUCNa/l3cUuRifZ1kTfg
TZzxD1XuZAo8zwJK29n4cTKXxR7SXOY1aGpaCFOS87O8t68bCQhmcDygWe/ZBS9G
u4IKEEmNS6GNX39MhPJMjoPYmHqRI1uwhPMS6gwmcS8ktdD3BdRfpasY65UxYJzg
DMLo9F5dBiEFhhWD+Urz6oYfPFOfMCNX8ET5SLJjPTGjIwjHjhkVhY4p3bO5oi4Z
uNHVLAJ05DW17PlNijK4TW/Hx0k6ef26i0zT5yqE36CPejk84oJJHybyynnZaX8x
4N9mrXNOc+lEHJKmgJHUxf0+zkQEyNtxpe2STCC7reDsupSbCslRMpnagN/gjZC9
FBQqWgs8Y+XcJq7J6cX1YJKZJdgPFcC8fmrNkR281aaMYTxCt+ASvudwpIwg9L3m
oY9fNA410mvxvSoZLuLglT4L+n64K6Xi248TtvJNLS8nqD3H8SXoFZWP5OrXU1Ge
dNIE492TrYPoszYn04oTi4OHoycCRiZ0KOXT1EhhDNsJt4Enu+vu5IBYoVdSV3F9
pPTe4J1Y/FxP1RX0NaKRYkxo2FSy/01RpopbWKDmIo3dXD0S1BzqbHU2rqFYqyl/
Cn02b9RSwjyDcs8dqgsXjLhD/thJNj2v46u++Rz8SI2VHzGFM5alRJzHz5hVpwQZ
AKfP37exJAYS8atav3bEzlmyzhpD8DUNF6QITXfBm3HCAvh96iZBhb96YFt7o/Zq
hma5wxw3AtytwJg/JT8gno7KGw1SCThSjhzh8hi8dPfZeLh9BWZn5nbW/OjadTQn
pU9s9r4WEDxj/Qdln4yp44601tQUD6vCybBbrn4y26+Od8AsknXJdWDxAThxVqkc
Orwb7V6Hdvo6LZYIb1Mj1WTD4PSE9voBTH8Afnu9CLiY8bvvkkb3022STUh1Jpef
Ogo802BvuJk2Y6WoVT7uiK2hB8T+7PXSj+iyXbwlbQ0IVRUFlPt8XpFdfgnZYjIn
L/njRQm5Nr6Wd+1mOyeWAXqJmF4A2xJrICM6Hu2CRwq+KsXarPr1wLYYZ+AemRlE
BpXfiTnnPtZd8uY6WaK7w5cuGkWuP/RBb1NVZh0o1Nj4HsFvX7p/ix/mjwYml8J9
QqzNgzw11xYcEqqR+cGL0U2STu/vKCPXUIX7pYk2eYTUvXQVvZHUXT/XDZtJfJa6
GIUDFBoAlqXFHLCkmWaJQL8dXh9tNAG5GUOSDSnRRq6wQ+FVcL4coRnJ7Gz4iFsl
B1M3WYk7bN23QeYZAYYCQhv75FkyhKYDhzFvcikRXTM90hBLD5Yh9dPNsASSndhq
T3GZqv265KVZgwRNvuRNfWrKN/1Pap+qzsTQ1WLmweqtA3f4R5OPGo5Sk2iGUwf1
IBcXZhwLJbdpkihlFCmN1s/sfIp47j+tA5mhpCc5gtgcFRUKVOQ+apqkXm0WNwFK
CMKm88hZOBrxJmR6fOohmAyMT4IioidXsVjn7fb6E5ZDkgHnwmuMAcaXpgRB2ngg
o6XvC34rzMRnOnaibXTd1JUaut6138Qw+/mwzgzN2XFZ0nYzufn3EV8CFgewr8kc
At3i/4Ry/ajxWVhd9Pr3BKhMdGNBR1hOK60/3gK3eDOsYoubbhFPPPHEC8zCKk37
xpnlHykCZxe1GFc+DRMa7nQSp9z1pJ4zyHbkk39y7v17A78djO7+j+kTNYtri6PO
pDCVNb+5PYTbQs6W9FPcrYvMyft7xdBieI0wVLEEfHLn/21p+VFzk40xl3SXAhQM
0Sfcmlo8+zMqH2g0MFQwRjwbNw7J2YICxRrbIULSd6au4TMOkw65qqtLv+vg2Wg9
+T1bBFM8SsimxZQlNUDvs1mPjxo9hCt3ZLGfcKIhWF1rWHTjG81HJVBDL+BlgBPb
CuC9o+r+xMoHMdPP1ZAawNqbqgmRM2cLHw3RbmmrldTG3X2DN6g86vukp6VEQfsG
VQUbRJCNaPZVPWkpyZFeVmOikcR6aP1eGOFINUCT26BFyN7/obCtLu3l3Ut7Gfzc
CCYurWJo+eid4CL18q9OsJZ1Qk4yQwx2yST6VJJaIhCRtMP91C83NRoEOpbdW55d
G3OluJ/4K0Mh9UYYVUkv3t5sKfTfLG4VTUOxG3g7VlW7Rg/DzLFl6M7taWajDISL
iJ2YM8Q1EtZMG4pR287BChcCvU/XZMnrfl2X5NI+k9vzlwguAZZsaGCFlnvuwe3B
6VOVanh1Ai/rZIiyL2LWXrTDGiQ3lx+ek8Z7AJB9smTyopxo3PmPyjDBFJIYEujF
SkdERtalM6aKxdLx9cmvoHpuGzJqeSein+9qE4IZ2SSYLwIh89c2BAowWhOVNB7e
vI9fji0g+tEc1og9OLmhcccFFTdbZU3evKUfWketdrEHfmPGWNbyPWTeZ80IMnhz
e5Fsq3xF2LL2smvt/7HgZYEyzj1g3ubkV5EJx2gQFDyYPSXmzY85u6eMjOKrk6b1
xKQbOzwAyQhEJlNUGiVOoLoxSiWb2KxftlFr7q3lzZThPqcoX9a8x0Sgsbo1PVil
X0qNMFPbQ7NllP1auAyRwfgW+Kyf8A2FHRlJRK08JjCGq/MEOYbIBDziU9irgIhP
X9wNESjzxBCXkrOnUphXYQon+tntLPJ6k+Ev57P3wBnM9YT0p7IA52CUl8vT8ol0
4NWqQWTGRKIwPyMDUi+VT1XGRS4M7fdywFj7th+bVjYI7WiVDBR5Rd5NMOvLvY4a
S1Uw9X7SejKNo5deZVoNYoVwqBQ3mjdHAKXMdZz1sGNvzSnpb4kpXocu66avHg3L
ge0XulSeWQKX5Mu3E0EDjj0im53Cq9qAMiQb4n+x4U6rKb+KuQGlq8Hrdu8hvYMT
oTvcIbamXjGEvfPQaz8ad0UjWap2yRS95BNGweM28lNqPCmJayq1/2a1smui4Ckw
MSDUPw3csVEV9F85ZiUXC4Zo4xIMhabkpPB/veriCnrExada3qDaUYFDIIOx2EoW
fZlqErVskWI27QzsOxpHIRrjSwrck9KK7Gl0k3fhflPRw3HuwWfhkj5I2ZECfUyU
zYhomOD5sRfNcEi1U3YAxDjEuTbfRetLbLjniQkGg9fgeUSBhsu/ZBTsc50Kyhyr
TkqzVyDB+e3Ab32Fyl0NsF2QzoS5abSllmrc5UD3GpETanViayD6zbMwKDAZrIdh
mCj4XCh4VbydjnHV4Uyximg5SQMz7T6raZ2VktYhNMbhgGzind5QE3JE4O1SWjX9
Crn8JRGSLkFo9uO419m+FN7laB4vkOse5mvHPUTEKjUJ+mn/8thfG07faaKlJBSz
glTW/t3o351GfiefQVSJUJ1M0eUgZhNUn+aPlkGpQVYQqsspktoy9LoKm/f7pLzV
/1ui2l8CIpvg4GTbP6h25/aNNJrtSH3bUwmF63xZlZ27tWRWCjqCLNtcZtBk6c8y
OaaHnvGn9rG2rt2mD8pt66oBNvL6ginZTkQckA8IMkgA4EX4bu1ks4FqUQhXgwcy
scLA7rEx8kCzg08lsWhkW106b8LGhOZzO9/edo2xZM0QvQv1otN2uEqTis3OXCH/
betB6qgk7swma5Spnr4+CS5FdjSPrd9FYGK9IZKGWwpTPVbIHLzYFV8HSHRtV1Nt
pgWhZia5EArrQq032EhwAWsWqDakH5H2kbXDSYIc2ZlqX1E1Wg7xQFh4cjzJYmrA
PbX5EA8wjPBkMpGh3lh03KdKlbYYOaqqyhfR8Zlkm5hEmS0f6KeYsWFre6mWvJvb
FsQCQec9GmhxOsqxCfv8SUAdHRRNmolimm38iKFFQQkTYh94isAlFIX6IoZzPRlq
9aG1am5Q6aMUwmQPJXozrjfP2CmV4jVRBg0yfOGSYsoWyitX2Yd5VjZ5OVrSRmWk
2N3lx1AHh/3hYpYnNgYkZRQcXANHOvF/nYBTowTNu3aBxjsSMRmL4DWMR6OUwroZ
KOnGfBJOIbQLE4fHkBBc3AQ3FzDrPIURKhWg9X7UDOgor0RqAHPFNGNbxygckjw7
gA9O47ylBhzbd5X6v9gTa9YeYXa38HBiGVUxpAR7BWR+KTrdS2SE8R4OfxVCpQSZ
B7MgTbkzIxf06eFY5Dkk1IpWt4oL7kOsb51nq0eRiFWxjJJOR+2JiLWCBQDiyvRF
XdTfbIZpsJfe9LO/WBNn0DOi2qYgQizJ3hS+j2a9z/0jQTXS//7kdixlZqEArTsL
4Njt9ncM0TQbO/8mzMgA3ELDGOARv4li5QWDrjA8fL4NM9DFij+EF6CLixGF8QKX
hQzezHWP74XAwhwFNVveTXnkrl1R95SeKNkNaZgWht91kTwYg60ypJNcMLnfObhH
L2652w9r5t9pce5leXIPn64nf2WVK7Yaz5rV9EAUmWO2D1+MQEmb1WwyCnn03rk9
LOZlGZL5Vw//oePLlqj3QQlRjLeJ/3TvkKdQOUl+CUljHTmOSLWRA6JPQg7MP3Bj
ozU1SYCej+EWmPOBuKaLvMrOnwyJfn5rRjV7697lsB3fD0BLhHX4l4kv1pv7UnHz
be/5IW2Ov7ePvti5eLClPo5+lynoNdvA8AWrxIWwqGgSqQWJxomov20X3HKLsgxR
lXLovfDLge9ujVG5i9ZfsPsMTG28nWosBo/cuW2Y51Oofvf3pfS+lWUYgi+JHjAW
mF1b5QdUqsl2LKZye/D7a0Iev68n4+ZcU5jBHO+J8op2DOwUitJkPKxt6rjVKo7a
OKLUixuF0QPTv56EflmFiWL818P3U31LFcZ1QPR/Ut/sp8PklmivlaPspNIQ/TNw
RGpme2CpVMN9opciziMFlIJteIhit/Ekr58wrsdpTwyiKcIPCWKD2FnRXrCKkiVV
DNAqiJ5ja3psp+swvA8kAQkLOjnXc4yPIG+ttAkTs59dkedFQ1WlrRDdKTOcvBQG
qNsxydpSBMwlUZ2HypSnGSPXwz4r0TQMSNVNnN+xVYnZ8v42EhzgLUwhPeJGwscj
CAOFB+vDmJ8Q/kaTmPdrNVOKi3EC/fjWjGZHkdupEN4qAF5sGY8qBxPzSMYh7ao+
0dHCpwrn8gHT6kZfRUP2evt+SLk57rU9ZRrLFVTl9OPOaKmCwqL85BiAtYE2qozt
m/9mW6rG+VkNaALtFXx1AF/Ow0QAG38j1wRjxush4k/0cuEYXU+HzwuCy4luHRIk
EFrsM2JdQoPNANo47yBI+S+TRdQJjVsx7lgNOgV5FbaNOQlbfIW6MwIIo8uPvfsV
BucnAJIDTUwIR0hHSyVKtfWuTbpEuBEUSH1zzEpEpKV6VJW9jPlyjTIzyqCqsF5N
sLWmayHM66uqhU7jKyfM0eLdRLUlukgMe/nEqeYws5qLt2aqf1kB72/iG1bkXUQ4
L1cQsknapjkNInQ76rEmqT85Nek7Nq1dnfFYa+0fp18WS4ezaljy6hL7WwVY2X2c
gDJkyVCzNBna4zxx4JjOS7H0eSs+e2YNHvxdM6HIeV+4XeUy27Yl0VDotb/17MA+
sD7BRkGMEytPSpNzrcyMqpGMl4UeLzFLlh7NyWSa98Ts+L/KMF+hTro49hT650S2
aKfBZAQSWpccIkg3kvd3MgMSGv8DR7ZfiZ+dBgEk8GmaqN8a3PlS9ZzmwgG5+ubC
OuaTJfvcvTQFma0vxs0rmOV11sqkkhpvgo8LQv8bhHfbPhc6J3xM8CilyahZQKj1
YkH6p5hUz4YviyJ3PYbJiG9z3tsE721+5zdJv/ZjFreonXxZA4wY9FaXHXSq3UYy
wlw/eKWjSdILbS4DvN35UTwj4MqoUwNrZaPopodxdVOrZX6kL307xQ3opxZ6pSg+
qMIkfg6a75mM2b66LblQj6oYfm2zjD1RnsuZzR8IlR4C6xPJvDBpDsLxoktR/NGh
9JT9hy5Zyfu7nNgE5lhM33bpB0ng5fzpdVBNPPC0KkoJLPnGyCc3wg2gtbXV23g0
iGiBDbotALGFi1HUTW6c6Gk+nHDdqd9iPIHA0k9W+mwrFAU/q6fCpc6xA5XjyVvp
6y8aOGI+PeAiV7RhUjxzthsMX2LiYg2kIsBIyS1u+ZOQgignbLLcJp4kWIMG84FZ
pXdIiwYG9dkqXLS/nkDpL1mezrrkAFUbEwiqegM/y+Mgpd8KAv4IosQ0XuWt5eCa
osUrLQwOzlVRMbgru9kulv51neoNWtR+CTlruDmIzKEZYms2l0BT/VSpMs0lPKZG
vIudL640zLm/lUdIqnqHzXJt09W0J1kl3osX4DGhQtz9hUmW651B87k5OgEXqod6
rsD8L9mWucBkSz1/tC2bsCUCFRa+2CN+WntWbiikuFKaxZ6uiPyWMOHtkEpFexjQ
BT5NyYuvVkDux/3Vdexh0IhVsjPGa2SHBNhfTZ/RSQPex9/TDQtNy3U0MWU7M8RE
a76qGkZTx8UIegwrKOTIUH0xkc+d0Q6Mja5t+PL0iVcgRl2pYpnI1XjMYOOMKXFc
jSMS31BFsryA5mxx8ftsBmxPyquyFWQD8NePbxZBhUnteaTDsQmaykAZBMn83W1V
Ic+h8F65XfO2w0b1TdI8dnCFMoMKXmpZa4/Uy1TessYOasPDr3BmraYViyXjoNaQ
va2UQm3JM9bnBOH/S6VSt9pxJ63mdctrm5TiH7XqavK+fnJdnlHR1hcnbsxDWphu
yti1f1u5cEZOyVZxUwCakrFu32WNYMgI2gVfIl0F2JSkSPq0hT4g4YuCWtaVvSWR
yTWjf4sflRboOkXk45K7hje9U7RnPkojD3NSY4cRNCZDi+MNH2xd94qKQiGbr1KA
qlevJHgzqeoKh1uGp/Vmu8/jxZMcwCrnGe/G4qFc4JXT/9MI2W1RB5nuckah35Xd
FvNmMZW3ct+1v0DIXSQEV6K3PXEJ2S+m5vOwyDYl1Ws3AW28icAJVw9EkGFeQnAr
x1/LRbLKJuX0FkcXWTnNcleBasgZr8eX76RJmvhTEu8QT0v9hwnEdXrdPFdNIwhL
ZTOSAzqlxJjKWiPFI4o+W08LOnYLL09vI/05x/Ajj4mWSV0BLx0CYRUXUwtvy1/g
+DHMZoiVTRfaBpVfci0Y6hMM90+Kmm+QuMdB3V1QPqjQFqTWCDCWZvsV+ikmFuFG
oUfA7VOVlIrBB5TiqwsYIRHxYNfVhuClSLu9pkYAWRYhBtE3EuUnmNlY+mNwaLZf
8XunzMvE7E+5Dn/yW7snh9A2vtTHYwbNnpKDVECSFTsL501WHrMVVmNcDgd/CJ1b
BKRlfy/yAqmqtrMKl/gx3s7gWG94UCEhXhxgxwMyM+lkM4+jCRhAlIC2fJf+MjLt
L8cac5UjRqgnYqiOywCA1Ya5orKVf3WBe19HRUaw7t4nzAoGrVj+5f2b+if0eOxu
y0BgogZFGOI0dQSBE4S8D2DfAi0RZheZqtMIvZSmCvuxob/CNPpKTrWe/4ogMTbQ
ZvjVbjIiBx2Wf8W0/Hh5C9QKsjCCSjM7dC/j6f8htBM1EtbPNyKN12tAwIk3DEv+
cFyenSFlLoPaquIVahGk1rYk0wf17nAWcBgMlTb4gdWPvi+ltPBLQhw7jwyRQfFY
tmRPbuHuViXwnoBYECYuGbnMTG077sdHGAzPl6dNS5GStzafDXJ1Wpo31QYG44aV
tqXaLCaM/CLrNtFW29oQAvhUdHFjj0jlgXNl1QQWT0tZANffQbqjoWe7zRKi2TxN
y6qISUQSapMLPYNFsPEx1h7AAlWUK84pCGyqt9w3sdoY3uGNePqC5JVPWmCNz5ar
3S5S9ATSASC9EhJFL1GTaF3hySf0CsPy4jrVtVAzUYbT5O40rZ4rFqdkkzhSJHc5
+qE+lwu41RQf0EArgbf3GHfdrhEyJSBLkBsO+Ye41dnr0D8yrj0vWNOBVs09zbYp
VN30zvTx7EVNo4RSSH4IjyjXrlrlArQ7jV6k41zrCl372XbfmrkBcqC9/uk/A+Pe
RWvY55yd+ouixthBYIHmkwsBS0d+KDPkISYGYmQU16KGf/RaE0UWiri5jXNhTFU2
a8tytuCNUvff2OPicLcy8XneWqFTnT5Xd8tFGauujZ05LiISKDTIZlFBgcICytN7
76VwTQ+rtWexo9rDSjj8/f16ry9W/iB1FLDkE9ov4ujZ0jlzXQMowSg7FuY12TiN
JWixuv7Bh1PrKN+mU6BfTtfHX62Bkrv3r/LSJGTeiaAhapMl762x1wlAT6LCKAOi
UgmXKaA2CpGYFTCrrhSEOB0FpGHvyx0ps2/BekMrGGgdyi4APDHCQE0pBeKxYhFd
HN9H/ER6Z/WTMon/SuljtbovzdC54ouAbkR9CXyk8kdlTIkDBru+SGSXS91JXcsp
DZFxGfpu+nvu4AWhyeI4b11/10jqLooTrxSdFYamLCkZEuWyIy0XX7UiO14V4qSy
5ISm1CdnSu4yaXGiX0wNvZQ7VXP0VNwrblPDrbOqUV0RB44TePIBe/E7I/w1pUdv
gD9azmBjiBPCNCfUxhcyvCTUEqIyO7mQCt2ddq2IBg+aqnS1JxmO4bvNt+/V9ZvD
QteW4hv0ORXd4PsYZ6BvIFqcn6PJaXnBcAMRvnR9UyrQT3kuwyV1Y2jK7DyF4CH3
F7kNkSZk99dwGa+qGjjz3CGSs8Q1rs/v1PLlSLUBV+K/CVL2lZDMlUtbmTDmCqeG
vgr3H5z4ijQMI/iR6TwNA4iqthcpC4HnUdSBUmapeEr2c3jvoQfFrwdXew1/ZVMu
t4mZ7hnS70ZRC4y4Q8B5HfWf3HNj9hvv6wz9RPPSpvZARGoAq6idhfp2akJnghya
sSMQXfCKV1YKn60MIaEr3zHerJgmavLK/TjuK1RVgGArTCp/MOzcCycgYFnHYCOS
dmDNyREGAaaMmZHBzmxAcavz/vaBCPjpv+v3p3Of85QRomFAio2myvRVrBRR7F9h
kRIA2cwhEkYOFotSmOjh8/YpoCrkvCpscNwwEr7yE5uQVkDSlUqFToPGVBR9ewtL
V7YCylz5ilFujcr+tuBToFt39UTGJkdQvxGN0lEoV+j/rUCHivbzKAEvtaoJ7+qr
/O3kdPo7BqhJ14qtpb40zIjpwrcCwjb3M89grcH/uItznRzUlsky2GGIJbJCFoeH
V1iEyUCGTEhwbSILl/e2lcKalIuwAvkzTW4UGnuT/roxe+52tleaqL4uhtuynW0x
17ZgQRbf0l0rSLRfqJlI9E1wchKNJ5jFACwhKU8+HKAk1SMD/O20TcuXLEU8tG4H
jAXxsaSX7P/YSkMuRQFGwkg2Pp1xan0bLNDN8USnGIGkMzcf7W/vWFId+tMQDmR3
c8BJWEvA9VfUbT7fXxu7s1zeraNoWKKRzEfqOGZF6eo+/UpPBxz8TfzvqfGGx3Qz
xD6+lM1G61bJCNAjRKOpTzHC/VdWebsU+H7zU9dbAbIHOcXv7O+7G+mu2Fr37O8w
SajSTUAa9foS+5gUxZKSXD85xxA7Wzw7/iPPAgxOjj1YzVSacu9LmoCRBhTd9EaI
/bdmjLn2LVq3nVoJy9gxjmZ2GqZ6y4BIeP94pz8vsG6drpH4vODqSucywcWcCLyo
Zh2tWzSoC7Kk2VU0OsXJtivTEnWXmSNVq3mYxpedjtRKuvNJC4sz5gWlXm0vNbAL
X9Bm+kQBzHwZQbsPmwOnhB+X+5hBCBjIVWARUMORysoYFsIn4lr4NF99cyGwLcV8
cNQXIIrsMp2aYn+QPQkHiQOrvy9KSNI+0PTSEFBpfq3A1pMB+FA5aj9PdF/149ys
Q1w3uRfWIyzP9Po6Y+m/qJepdLO/8vOtvftWPzYosv6diPvWBdlEN4htWbcU71tX
vgPwgeFVzgj6jJ/hJBbEuS3pcjdijwEv2+mYCBRU/1GWPNuOpu8PWsKKoPf26e1k
dP2P7wuR0M3DPLNJ4IvG1F6yicTTlvv8yzJw00himaJ4yzqHL83WLwYA5Q9a5cvS
mrkDHfugbviUihUYaM2Q92aVFXTX7EMmUT41b3fn3h4LXGqwBsZewEUpqUrwHxRe
5ypwxiQapzCCJHAnPLMdKuQV+m2vrMZg2x6mRndv6WDJcoSgWk8aZEWR66avZJZ8
6ee/MASI6+dTT1ASGAmCAF/aa3RkstwdD9pvvh0ODJX/5dIOnLtY5+TU2qlpoWKV
PNjLlAmUqD6O+j2UMThkIp51IBvB6dHF/th4NUNIFj+iqN2Q/cyXaGVj4xiGDrDz
//clWJxcLCFQvW5dZ2ENGNdKvhnfjvLSjs0u8vLFyYU2zVM8G5C1V3IpNwK9TbZe
rLLA9iAnqv4RxjNXvBfKPi33qCuATz/13cGY4ibzJIzTvTY06Ir9ku0lIHHIj6sR
MwHtEx0SqNTS22Cmp6PQhGiCZooaSzI+LSGzim1rr2rRMdke9jwEokCvspDsrGkE
ziQL3YDXsH5B/11XSczcVoLB7g3BLtBw7yQ7izPfETAnOc4QsRQD6NWP5R21sBbv
4bCQb9HRwoPAT//DgM2S/GSE3TrZhTC6CDD3rx7bHrbaWKD497cFslWK9jU1B4oG
jwW1EC/HZ8+3a3OAzme5pUEC7v8tsHI82UJx12xDqVh+2sOGc5fZDY/uRocgKa8w
NTyerW1ObKLMGx+nnZ/hMZz/khpMoxGxyuTGnfpnc3OBbcSk7PqssbYQ36KYAKof
Yl/IGX7OoTMhxNSqIooZzoHCHLrTpnQlAPK+KYTLIsTm7bGuClC8v0FJcPATeivG
cxCrRgKvJxx/8UR4qz/LCJKcFnmPhoPPxrNQ9zkeIGFZ1VLbf6s5zNigUHXg6B+0
s4IhN3Ezb8BVFAMZ14lyRCVEqXJAKG8bBCtBPWOi8NIHwIoN4z5bNzeKfmYaVicP
tLwF5Fm3Qn3FVBj5VjUlnnAfIuqc/uwim9OqJSPkrTxQx3sIV0jBop9BQuE561Aj
TR4wS0DLlMvqmAy0ZovYbQ4J0bDtj0PjY44RPBJHbFOwYPHDI39mi1HXSzexmMQd
2CtfHrelIQ/sqdlje/g3mGplsWaEIbJRGBBlGSCh4p5B67Y0lXiOYg2k2KFAExDh
cp90EnS5IjHO7ZBZKtziYH3s3L390s7/ARb/twmhSHzBB2G1OIMvpwojPr9zSKdS
ty/vuJ+e6JC9i91Zr0xxHC7rXS6Cykree4Z0tLdi1qQcbA5KVVYLp0T3iX3TMyL5
QJMU7L7fc69cKUpaoxZEg/ZLkHSDLRPTGIpagw0+RNG1pOHqOitaOwJGh85ALE6b
wlsuJ/kaxREnqQHpQvcJRKQ8dq7SIyT5y/yCovXBfVU7+everKtwHynYo5B9wjLf
iXlrfze9pJuPGy1TMqhi2VE4a2FbRIPjIrJ2m4k6curaBY5QzM2gCOakWe3SYBop
Dwla9h3xQ1Kh37xvVeqIcNs0Gy/1J+Kmc/092ZQCWpV8t24yRKzypC9IxekLF5kY
wCjRaX0GDdoXg6fF7vvpK3BPbFWPzi10j7je7wUPtdkf2u4FkOZr3SwawZBT0cBP
JsGfclECJLMgXcm1Um5snsc5ZnSwv7eIMcsr1RDDDAbcMXex8/b5foNZtIaqxMVu
PKl5ySesS6qcvbro8I/pzkumTZ24opLR7oWn52wMVWtMXjwBOMiZdECndZCG8hbJ
tS+zUOClfaSdoGotFZaANPxf46yDtzoN+5+Unu6IdhnRXtK1WYZvMTrB30zkvZ0c
Vyd+5ypIx/IC7RoKgB9bHTRhaxwjMdOtC9kFgp12St7JlH0tqzjIxEVfBC/YBcz6
YHreBnkK/a1EzXAbuASViz5ldDlhAIPkFpnS1qSXtKBpdr6/bb1lZWY8M8qRl/sj
4YNqpZt4cip6Yao/w1KT07QOP1ux1uLlx+Gz/QQLo8y8ZEclzpvudkzwTP/wLnFI
/YLL14bSSIeQY2e0hIHqehfyUZIvVC9BiTzKpoySosn2N4mb5/Ovi+9bAD0CHSo4
SOsxl5PleRer+uaZF9qCZFzQ6g/mNsVXzNZ8CZcZZPBi5bO8sHMSrVRYC7vdnWo6
9hK5ZGliQP0rCthMldDb9dkcUgM4m7cAl1rnd8C6yqDAHLaCPxQKT76mC32oN5ke
48r3m3sfD2ROGKZOw6zQMc7wu1/nMIxneKqO8ZchFTCyIl79WgXX/J31Kod6TRqp
sQZCc/g1VcujMLMBUg7U63HmU1pk/unSOjT+f7B3ZyJw2AG81mOi7INA5sXSFs8v
lDF5dfYYgxzmA/btQSJms4TVy/W33CVNI+2acSF6krADuVfcaW6qcSMGoRi6s8b+
ePZ5fock23KPgPF2Oop2yPOVoss3+FJpP6ibgeOYvgE1YzpqNxeXQ7k7XvpzkaRu
suwK0hc5wbWi6q5ZJZd2l23ep2djMYGHG9tmUMF2eUA//nRx2yPOAeEkRCILH7YB
kLUzZLWThtThR/XH4PfWv1/eILvgem64MN5W0rOF4y273/CXaeRId7MWOBuvnIZn
h4hW8PkACBXaKfRNoBu0egWEzDmVcrCrl97nnBchKr7Es6lSu3DWqY+AsNmrSJuo
HK12Iiom8xo3SrWgY0E235yeUTQizLKuppb7HGCUIZ7yuY3HNb0n4wupVD1JFAuh
RoPlFi0yoOFTMwqSXLd86wWfxvav8GJwT6iiiUODieTVj56eXnGcHJattdfdhUIk
79SzJSFuchHByZlZMY2muP9fGebBXt6V6XkPCnaZsysxQMDssIdj39trBXcxWDL9
AwVratRB2SGE/YWVNRDFCDuTV093ijv4aH7yiYuk1oohdGhdSt3nZgYvbIODzOrR
F5L0oRA3jJwRzjexaFtBPldyDpboQypCt0FHHAwPfIEi066gR6VEjjNGp9TJcSls
jH5wxS0TbIJ5pWr/JU/hM+fEifLhDCkSz1NsseTlQBou2MA1UhtntySMQ4nd7Rm8
I7O1uDliDIdFi8l3drnwE5oIGOjx/vlyK/XraJfqVV6Tkimwd11gKOZATVFNKPXC
UApiccFl4EUWDZ4/ry/gQvtJpqfRk9QV+Pp+ryJ1UZuGnhelbNnyvc1JF+N0E0z9
qLBDPLfuOSPBq2nHd1LOw4NQlZ7J5C0JflriXQT8OFbT+RjPfnDhRUOe1H9vCLqn
kc3aAJtx59aJm/QxHsFLHubztoTXtqcztOTaKWbhTwioexO2K2n3sG58Y7LDGbwh
YCUgxXvfzixSd+a7t8T+uT9DmMCeKZKpcaynVIj0WLk/u4QkqD4zd8EAhpISL4hl
RXQCKNYIvPA/qW0SdHXPmYZHyh8rjD9Po1+voIucMbqG0/5H/3CIHrTmONsB9vnK
ymVkMKobAE85Gry1LBiduQrBCY4IEoCJ9Hsr2aYt+a9cxdFWZbuDODsChDdMkS65
fuNo3eDhkKs37BuXhuBtRxx0TMeF/z6/1jQzO/o7ueCAg608GkmcSS+EdGICT2Uh
JGTPt7caUlxcEa6mP2IHgX4VnOcMv8va1IvOCnCu2JpcZk1/yVUdYymJU6Z/8VDH
HmY9U8/e0migUS5hdBrP72W1YdfaEyHAZzBwGvrSgAEbVW7OXkeAleMwxJ3tztBh
fLuGqTF52uMbSm+/rQP2YuRqjtbmWyrqyd/Rb7N7ji+PUqGr3uWWIXllYBN3Ht25
ekQIBT5kxRfA5bZ7Ps11t5uSjNk/Ml9EL0smD8kVqghWZca+T3eFGdGKHLEheA9i
AKA0BCrHk18JIcVHDK5m6lZeG4FXUtFCt3YBf/OMJsLoa5ORxRoWz7nc+X607qPb
72wbWJPcUeD+C8TyEyE7+fDRXEnffKyR61jGrQ36gJBXF5PxJg1Vghu885chymTh
SaH04TtkgRpmHk661It7/m9F9PfijegYlRWywZ4wbYKkN82eX2PEkE9k15qCF1HA
kLzYjfKYB4A9swMqaWE4L+rl0Kikp510A0YdMLHm96Adm/vItoCZOHqeOuqlENYQ
tuhSJiOrsobmWaVDB0lPERi00hlC51TnoHI8D8rZ7XAnslQ93dxQhHIZhC0dxXOo
l4HQZ4Ap8UX1ubJ2i3xnnf+cpWpBLa0LeWTb019RWK1nTFCGiaVMDCgfC+IXJHX9
Bxg6+0com56p0sXZYFWU2VEOerVqqW44Pp/IzaRFM78DTfMbCh3wUdt3GZGttSRg
Dx1NWBz/tO6iLqLOZhFtY1y3ckwuFua3e3XH9HhwcxTkdbLA18vlf2KPo+2QtUf4
64phgqne1ZQDTRm+kFHbcj3hAx1d9k/BfPHgAii9FMETTh5+MJFBjFVB++GNdVR/
jGMmP7PY9VxzWzAcO89NPn7OAH+fBkgLGoIyiY4xTqiEsPvxBFfHo8J7mwo8O9RD
d7HM3bnTxDmAe6C0sBfaZQkCdRQR4y7MG+vM8YDDi1uVUWwX2LiACWow0UA3jG+9
qlgO0YpVovQNLRf6b6k3jSBNYCWyvdXElHTfT4PmH3wFUdzoqJULpicLhbcIIIPL
buA9Hsb+6umhzgDr/+MNoyACbZUxnpfyouOfUA8+TZ9BsqYBBcKoOKV4il8XTQNP
mAa5UPQbB5cHXrdJIKrn+uhnpw+zRsgJVPVvjQWGot9qp7LYFRanaIbDf4sZirhB
HEKicD46MYERNDlgBxDlstM1w6KMXHdleCCBjIqx5oEwF93stKrdJGP4Lna9udkc
STvKzw5yD0TGUe6gpBPhymFs6vegWdk5kC6Xo9G4dtLWjcetygwiVboWVL0Hsvhs
e8b/647UAR76pKmP2bcaA7c8+p5sUp70Smm6h5NxCg3M0DF/Bf3kFYOXG2OMBqyp
tWFBnFpQvVVdwoANtiZEAfwqhdQQbbkYqCY2XdJ0MGzZwz/mqRJ7Sx6csEeAb9vb
1yIOREjk9Q0WMk9V78mWeElRnhl39owBEAwu/JZ4i8tvJN1Qcqtl75UfmAawwy64
OdOEG653RWuo50ioSmpUuMNhwdGULMzOYHvJ5mUAvUKdEUAmVaWho3+EqWv3OaHI
z9mvAIaSZzblwxG9zXqx64yEEyI1KHkZM4pJL+c1R+5roY365YmEltDaGTFUsdyO
5C7PhWvBuRYN7ZjOS5P6TtvYQux5NciB8Mqp05+aB4LUcCc2TFIeXxfYNuJSnVDf
b6CnoQEaenjr4WYGn69Mw8JMXJp7yIbs7fV6e27QitcCEpfSj+Edv8aEElvSmk1S
qTaXBfAsi8N8HewIeWf9B4BZb8VUhYhu03e+YAUN8RfH1WNdzGXcM5uLg6i87Fhi
b7fjuJPz8pY7N4JQn5Ok0tGHfjmRad9jCa5WEHqOjxpww+1VfbqcAtJpaz0+o4NL
/KcuhmwbWaRW9qbi2dy/K5uyWt4U5mNdiiuGj4yaSy72xxPVF72kZNM4+Qt+JaOO
nuGv8ifFVc6PKe9F0LLkBV/24BvgKV1x+gjHEpVlzIM4ihE4dQaClb85/IBf065d
zF/ndBr3RNE60/aqNR3Fm6wpUIIIeF7vfnE6IhY5e4C7VhU6J6dL9M7a6XVxDxYE
ABYU4OpgAUmExVxBsTVnVdxJicyd30tmZUG9brXS7HEof8AAzBgDr5rRl0H8ja0I
1yFV6+WbebUTOc7J6YNatN/jVbysb58gAEfl3UNGjyI469toHUIoJbVFtw4QTIVu
klpQa04rJ8YLUoeqhsdlb0C8UbVRGwAHVxj2ePUBfh9xX+QM8KHghrgoPpWriRgX
TfOH44spI5+vbbpvD1wDOlNHVXCth34mK7aqL+GkL3LCkvGPP5/m5ZdIwrPwFSHk
k6keaDcF9DJ5QSiVxSo+0V5WybwtgsUz65vntuYtyVZxCzVKz8MxILqNTjZ0UC2O
DGWjvA7ngz0cKFjPgjgrODVDJhcr6vrIXK7lOkpBIwOv9/LCI6dNctvUXnGaBi0p
w/Crknz0PMcPq+P6jiDjmp3wEd10/1VmrYAhQ9vC1ZsNjSruLn/ggQF/vxgKvnXW
Nlym1OH5z0fOj6Bz01kF9+I6X2iTYD5ve8pxjE8Y3OaKsi8Xn3QJNkWQU+J1RlTh
WI6P23ox1SottHMhWwyuVv1e9QsHT0m2gTMAmLzSLWiZK1CSgYkDRO87PMvXtZOm
SKwI7C6FYsD4em0NAPweSF+m3E3FcXWOSFwuGGFuP2I90N6rCmIa2Ck9y/a9qMgI
Ang7hE/1H1rs31G07L+Pn4KBEAPNLs51h+qD40JbgbxdozhpvdmYZoqEcW9wkUL6
3qQRYQqU3v/LqxAMFn5SZ7UFwi4MfovpfNXqNCeBJTls9s2YIW5uskTVuAyznFWD
qqaBFjutPj/U8WktSUFZzq1kETc0xZpQ9lFH+nGXX2o6KwcbAdcb7GEclfm+kNQm
xPM4n1kSLoWAnXpenj8Wp9Zw1sXTnqkma2hpem6s1zOZ9Q2Bw3S4ekWG6MlGJ/6A
C9qISnZ28YV/rF7pS6PHH9ZUHf55+oZIz6HOJlVxuZGKYpuJoQz7lNz/m/Vlql8C
vMva1hhef6Xt7s2O+LB3Dq+1yCUBsm9CV60nkE8o3YUlsuNlVDHZD4z8/rbnKR9a
4KTPUVOP/oLLz4W9imyXmOjAAoUNOEguK113qcQ566mDKTYWwIsEhHSjE6MDnv08
RrBGNFr6lirsPo/clvMpypvf14wl6BX99uC0bpu9SowmpULR9mLOOqEq2teKUavw
MRZiWW12mx6drvUNoYjBldaoDEAgKXckXHccY0kcYB9ShzOBgO073xFVKWQVle7o
3MH3IgH9uPOSR5VWqUXV+PnpHiZO/K/ZY0KEsIO34P5lI9rh/ZI76jl+f5eJMwSt
382Ho2C1FDuqj2oBjs2sT1XEI/Vg8wR4xMMxmyA8v9Y9v7blI29hL7GNKg3cW/Tl
Bu185Pgvb0w1zkJyD2BGZAkiV8ohLGcPLYUI6++SppR29c+lzIlswlYW9c7v1cuS
hjRrdbfIpMqPaNQbdW+eqS+DCCMA9cmhPS47kci1PdKVD6Hg5mFRSwKXk7QyWID7
OslHQAgZMHRSebg79zq2UpZR0GET22wmhHzRVrCbJ5BeZQCFjuiV9pOz5wcMob4l
kfM63cXkBTr9hW3vRp9tXfz9VbVirfjzvsjoBDOhhIr67jp8OeKn5qfo/rtvMEmX
7/qPDkx5ZRL/CVm/sAdYpjwZACbDVGLjERu/qL7W2nWU5RnRr35huw6b3MEcJ0p1
ZqyZysjh6Wz3wwCzFyMhgEUpLDkGfcVlTiDiCuYKpOcjymIjHhYcCiDjpDy6smX1
ApAU6gijVFluizVUS7EvHWs5mRpgV8SRWXD6qBIbjEUJiC+5MYxznTIJmHHYS2xz
ze6UD8M55lRsYSvG1pMHmHi51fEVKM9RoutcVQwLFHAr7oumcblBjuJYtxHdbJLy
baknEtXfZGnMrf4GjngfY+YwVQFvI/jV41QRibZqem5GPPIwbxQOURwbkp+Xr5O6
ogUGOynJ7J3BS6ivJvgdl/sOTmoiAfowQTBaxMhRUrrpb4s6U1csjHLoLjJOxv4R
w86GN798N4JQ13gGhnFgmW5Wjaa9uto+rnCEAl2qY4hl9D++IV/CE+a2+ENlD4Xb
ZFMpqCo+DsJkKZTPWv7BThfBV2XM5y96a7TkAhDiODP0T/mtoAq3vE8FApZylrCG
HOUJYG4TPjzUo5safF7HxOEMIL5vwD79W77XBKz6vHzjf7+6vGF7iRUbFd+em507
SWju9GO7TVqVWZv5MOGOWAteridhbShtdXYUKcow0z7PdxdeZJrmGw6cmMI9XnyM
T8cM9IA7Umb9A0SlXRoKN4K2fE1FRE6KkAn2ikjAcPoyklcHHVs8RwgPQ69LvQX8
DaAJzxzp0yHHTeSYIFBCmaX/T+OLzzwa2ah4PP9EpRZ0/+1DRVxqy0MUMKWrsZuj
fkogL27piuH7oNBafqGmoWgjlZhyJV/pNJyEcCJD77WQTk46nUN9mn7zEJmdW8A6
44Beg1YSaq8LUxJ2fdI7ybDs2ZHZHqzJwWwaZrmypw/AJrHrOpCsZmnkpruK8VT5
v5mInRym38knOxry7DAl2Ojg1saomRzqFcUMJ3pKtI6HAD0EFbGYu5auIGfu6Eqn
8SBCrKzZyNX1xGlOoM1fW0VNK5jSVS9VeDqG3YX4g9sNCfj24v0zTNG0w+LEKBzS
Bg///1MVQoHPk6qolQQG8ZIEyJPy8tv4dgPXgygNAJvi3o2Q4uYD2KYiB5gHLwHb
uvi1VjQOWEl1baNtNJeBd+XOa3IAmv8oB7Kz3zr5BsZqKuz7PjMGL4Tx1JB6JCDy
KFktBifumqEJa1iAuOSBSMFr34sc+z51Q+DaJmIxy45dEPWU40wP3g0LG+2HnBLc
zTlZamn0jteWUQWDVAaqtoheDjaus/3L3TiBZWi+upJto0vJpTbWqYCvwtHK0m/J
DH2k9WHYL9IUwftqwZHar3ELUVuCluN5zpSR0s2p0OXuYVMDE5KkGoLcOpeEwomJ
Du3fQeywMKNA0+nGH2BmQOzZAt7sPllw1kWNcKw2ukA6PJYs+OYf74hxs/swlQ08
LBnT/8IC3+9juTqAQOLzPK26BG3hBdZDQ8IabqUPe2nyDhYyZ1lHLzgISPZLo/p7
kNI7TJKvDR34Ia3eWWwRwBZnW7eMnAL62HOO03Ey5wwZy15cOyXToRxPHOsvasY0
hC6SaIqX5CakXC6TT4hcB0GUkbDtdisXxIlvpq0enk1qyankWvaDIcErw+icJv3x
lNg5xaTsYPivlZssJURviiFv1EAaviY/zxmihYIwc3SWoghQWiD8bgqHOR/Kvcjx
R8kNOpMszMgfpdPb6zEKLIb5yYEK7lJFMr1o5Ttbn4eYT5ItqLmA0tSURNRTtnOr
Cpheu4vJC3iDYsLF0UE3qKtYDd/2uteCtDiKtmt+dkXLrYPD4if56B0+ailUNV25
csNUXyu0WIlzr/G0W5AjD4sTFQpR4RKqTFaGbMui30g7xXSeLw1sSp+ICtPCh+V0
JkXHlXac1E+u+mBtiCiyJP27+FQOCKj4VY+zxZGHYhPmCl+KDFV4FIm++0cyVZjF
FuX5Dh74hIrsAVCIlwuMbxn6npXBqKBENLtbiR+9YD2J4eW8A/AY/KWJOMFL6H6G
8vTxM4WqVh32y/koxj2zzCG+S/HAFhQgUAM4H0w6J4OB4PWPX6E33CVAa7IS71P6
AUoN606dFFg5YFyvl4ig0EvsBK6x9zGVW1r0jM18jeL/0Ptd8Dk/i3px7gF2SLl8
WbOH38qqk2UINGPv1q3eg2NYEhVsslK/ElMmFeDcYLzVMKHjlFm83HD1Z6NavSss
fCgDadObrP4dnIj1L/G23hYnOu73EArvS0RFvCyzTNkUAHsY30SOrcgz8XrRVpxe
6i3qt4GBlQiz4xZ8mEXRZaWMbiQ1SDxJFQ05Z4E56uPuGQ7K+jQ0KqXRG2ZqI+tz
M+KOHB8MZXZN/KHhA+uBY5zinC0CHyjqKNE901V12IoP7//s4bgWGY9EWlUdhmZs
kNq+AT3Ef0Eq+/QnDuFsWMcOZ1Uski8D99oyz9xg6SFpozUeqgL0Sj06y/rjje2y
pJ1aYeKcwrO4eVWbduwlGAt1sDyshJ4KEuPY7y1uY6iVloIWyXbOzRQsooz1hdhC
d0JE7CHmXkXUC+URxHAZ2TxaNoJnHWEX7Oqdj6bESoSo1jHqyGyrKJ5Ok7YmNmRC
ikurIfkQVYNnRFVVMhZH7fRF6zN+ldSdBhe7I0hlGq+QeQdOq4ZGxAa973Uxa1eW
3dr6OcCfSBCPI318+gAJl+2m2fQ2cTI+PHWr4dO4TCN7R/vyv+hL8hwADfnWdOnt
COk1SKzfRD1YwfDcDihdHLBePBo+9C7FH/p1XFkd54Y9qcfxgiovHq98HZMdXRVO
CUfUMHTzRVFYvkmnRP+enZ29FN+e1C6OTRPmbp4ttR6xIIs8u6qEUm5BH1zNv3Kr
t+m2vWysP3OY50oushPlCuPWAWAxIyOZfOfFz9NHLhPWxzhyCZA5bu7dKGDScr4Z
VwqXIpNByB90eOz/GdQoarPWzuQq51yKlh2rfCdtbaqf9ufDlF8L5+Y5IqI1y3g4
Khuj29ZUqFsTNk9OEw52ivc8RcLlwr+qr4/VLmtSM8bVLwChWEtwoB2s8bhKSAWB
S3FB0Arsoa6eufJ/SJy3lyev8osCyoos3VCsokIeM1jx3bVlnyUAxWENAq9oAFpt
iqTcttkIuGpwa9IY/CY9roXIKJ/M7KTgbqIxXUD01osCwrehAnKBO93JJ3M2VkWV
oaKOhxoj7lHbelK15AAUVD24SdNlAIklGzFBNDlKeM32lKSVZtMUKvgXxcssdT3+
RS1C8nvXoKvC7OV5obivMCHV13S1I7UNiSRvHjVDMXDZiC07anHJsdsBQFpdPt2B
vstMW/WM3dsz/5EQdDs8Vo/TBMPaE3H+kNxJzBotAib1L+5+2qKk9rwdSVTVpfwd
GUqA7Vx22tfXVDHMIZ4t9OANzFyM5LD6sS5nrUT6d+O+FA+JL+y1lwT/wdfR9vRy
WG3CakCSUfEvWVarlbBLL5a+3s8Vj3aHAmkqKdCuolLol+eWQ/iEzsFGOEuynVdH
oLc2CczXAvniAzbOYoa9f6Rjl+WaS5aYaAUBhOsTmsiGqOmMX4ty/+srD68jFKS7
w1JTMxc+TmKkfA8CZEjVhBWRgDQns2XJKRRo3BHdR440cL1NeG3s26S1XhcRJ0M9
aNKt2k5cgh4UE9peGdvDyXk0Vye/5s5bgL/KV0RqT1PLldfh5BAVPxmtQzoC/If6
KgpjXJOBPqvc4htTw7P2r3Srl6vkfsGPowOiXrQgJL06zWFdEPK2S38gDzOv11ll
hDWhSxz4IwzyMxeEIKDUM7VUWvwNkM2OHpytkDF85OuwIlrWLuHWyPXYI6OOKhnw
Jc/5fxeim1e/m/vwZdOUOBCutnaDAJVkQ3znz+I2UqxL5vtECWrgO6TIt/CKjAir
eD+ly5UmlOateRTm0lZcHpiLzJZlEDf5xMkmSX9Z4Egt0bE0qHVOHmBM25+0zoCJ
MfX/LlBlMkYVdF2eoYNSBoFZegjOuyBYhU2h1abTyyq/ZbtXB/OogMpfFMQuaron
AoljYmTLDhoUlJNg7gDsWRCUinSWj5/YxGh8mkVgS28FDGdLYbvbtMIN8qNOkZjO
LE7uW4f2JnEramXRqlcKlaIT2tutW4BOeuwWK2DDZvoEGqDLR4FYhFq3mf/tIwfa
HAr4nrp70x0syXjNEnq3cKYo1Q6LWL3Pnr/VcD8vl03QuKiFd3sDMWBZKEjln8cJ
aImyLBbzWCdiYdhYBH+8PDZkmFqhNkiTsk4qUn/nNQTkXKyZsbmgy9mlW5P5clbp
aEbEpBkTnR8/Cb1vN/slN/TnmCauK4zaNK3XNvJqPo66rM9AzYtPdsyxXKkyNS0P
PXoOemBRDa/U4rjffX110WPZuBcuIBdAdn6fcNvH1nhTbVul9dgF7wve1oDSLyeo
VcN053bbOhbJJ7BeHL94B3pQCB0QdHPxJJpmHAMPCsIpYwx+B1FYkcxYPvYyk3bs
c1UApCD0c3fpZLic6NYDP6EGDXinSJaCbgRUPuyUtSqjcbP9BjO73XsQelBkaxLK
T6fbx7/hc7FFNniaOGfnU1F5YtGWy/kWLmVaEhfRzev+SqZ2RuKklAyP9j+Nhzr1
6q1ZRscOVXm2b+EI8EeNkg9LnOOYBVuqqyHKuJQAARAlnURN71q0fC5dx2oxc7Mp
EhvNtD2Jn35ZlC2WAfa7LwhW4CrFwBHrywnjBfpULqP5SJ4Gtl0KDIz7qkuT1JEr
QKTLC52nrrIKZTYBVY4RvXPIDBLlRuaiarsAd+QFlEj1gdCHpEn25D5XLYOc/EHV
Bujd+M9swX+K3RGx5ONtSp7+N0kdEAG7GJPX3KI6/8fOsw+TFThYP7bF61doMgtO
RIsx96OM58dgJSXYcYKMAlBX+VrWDyWC2GJEB3iwxLHaGXQbWNJX8+MT3e2jcUEo
Yt+wGNppADb1o/Ya0to+2/aNNQz3Mjg4KiuZapqhj9YZxEffqqzmlLPAL/75WhHl
tjRAOHnEteXUzVZYarVsZXAec3gLOcFfyFbTRuMDrDRH6JuBzxa2hkqqJLRuOZ/i
42hQTLHLl8aAZ+ikLB9jFEo9AuvTAj1Zowk6dU7Mz2qYJ8pO4aS7HIurF3URXHMT
bABHXMtlBU+arB4Ax9aq5wCeujE+J8f7Urz0oofWqZySYJ4VSW1JuQofDWc6Mj3G
bhnkuvJNiPW4sXwsHSCGTeChKUbzSIid9HXkum66mhAJbK5As598DmunPtYzEvZ+
vfsivTjQo75926eF2a63LIO/YP2zECY6GyPcrrLzn75m+61FgeobcGJgtSzrgCk8
mmUY+VB74Jg5kFl4g1DLL6NQv41Z1RTlOLRd2NQuDrjynkkS0wP0CbY3/ENhNGGS
s02QlX7Cfip6y5C2lUDfL5JawESbzDTs9CYjurJbN9avhzuf4yKpC45/DYy1liE6
IKUmi0dv7D9MdO5PXml+crKPkyneT/mSlecIndp6kNyuFWFLYDcTky25+v/kJiMp
9T2GgCrkMF/iMZqsNzhZVktV3fAgxvkPVkg9sSkI0W+FYIYPBAtD7lUezrruXygJ
ZhidSP1QOhZoIZCvVpvxJR97vCh97OWiWz4uzNFr7+ltM2aRz+SuIf9wW1GXfal7
aJvGmRtbJS3BbDq6PdpF4L9Jn4aDM1MwWXQOnZpcSzRJK7B7MJFh9Bd/z4OTva5X
1dycN/PYkKidw0h7/KKacaCl+XUlCL31Au15hPcHvUPAaVNOV8bFeV2tG2ffVju0
y5cjZILEMtcE5sSTnUtHbg+18VdLXwxml63ZWN6BJlypcjq2cFCAKZ9KaahFUljO
V5GyXK3YmjY+vy4Z42iyjbJK6CJOVK4LojlrBAWOqhIO4a452l05idRNzNwIpR6J
TftxPMd74zSL5nbodFfiw5gBqXWkEBvCvuYrS5tUrGIQV36Z9rd4BR/DGAJVqB95
JwuYuhSNIS70MDgKHXlDoQcgrOP47HE5ufZU5bP8XXjbUahf4ZafYvopwgVRpnvl
V4Bj++Rhyky3Lhpn3CrlBzrE3f3N/CuIBLMcavVt6hiC+adjG8S/VtUbyQ1NJ4Lh
C07MkUyCO6JO5nss/0WJBudUYxn/bfvnb15N5JLZu9anHUMV8YBdN0n/zQNaL3Yj
pqGolfP8uwesFWiYLDrcum0zINYKZurd4knbAi7RkqoIKAIRMPKgs3YCfDWwlQie
NgH6Ih0zRov7Vvg3olnppN2VvcYDZJKGxvlS3wSb9iHb8JmLFXpyRUFbcKvWYj1v
pFPflVh2ZX+Yb0UFVXUJi3/RCCHHT+UqHgBO82W5N3iRebqs2m18zozqf5IkJh87
C+7/7EiqoeQXAhKSrO7bveOucEx3r99gbXP4B/CD4hRFfVMgV/9CGBvIo4Df1+q9
25234/fkqK+8LxLChL6Ty9FmDHes0bSLo0V0t3S1FTwSo+UmY/bB6EUOck9amDH6
qGggGDrkEi2WHvk7+cPVcBpUEFSrh4ZegyhY4HDUf9LA4FFwWXX+LYjAGDkcNfk6
ZHDklQ71zsSOPUwPBtF8qz4yU+T1qyr5EnXlWyJZ3I2P2es6d/KKz8d949Fvjcij
Xc8QdP5IGG6d4NrOWuZhwnTK/m6tULA2hvMz21x8MyceeN8695UvGWpotXYlvDye
f3MmdM82kRvaMpfBpo+meWxmx+P13eyeFxMA5mEDdbpGcKfrtD6Wzqp6X0BLXaEf
T4HO+gJNFdPnSzGqkv9EToFaxpqheypihN0vEDxtw//EIy4Kajvi2/RqSwSqk1mY
z8rqxncXzNGlIQdYHBWURK9Z9T2P2DVmdAcPzbksPDF8St/MwpvbAnzXip5sq25D
VkEvOtB4Sq0gtx92zxFs5ohpXDRR3fK+VbEVCxpGDVird6+3JGAF+MswmVTdsMVj
4o4RuHHMy5gm5Z4N+hNv/ntuFvImW1hkjdjtjdn6DsVz5UDVJHDsAdiqWlYQlqKZ
dNPaCqwkutiUjTkPROk1wHyVQUmGBM4TU0EqNHavGZsLIJeGsEB6I7i+zPWQzXti
6eW6lnic7o5rpC9TcsSArLq/r29ioXUQt+FGjdQ5SLXGDvjgQWHpzWozurSmOBLD
6Mwf4BrxbXOib78/r8CpkB53mO4AN/R6GAHVSYFusMzI/wCNX9L+f8i9XsDDFQYk
uTVNT1IfGuqL9QLdtdRn7wYYbJXXfNegi0oasTwIWsK5BbkQYxP7kQSc+GOKDfFJ
Y94Lo4rjCvbBUImnmlRVKsCe6HUflWcvibh0uNbEB6nBuMABtyTZpyl5is5ehTIb
Ha2D0DCvDtFLs9pr2Wxf+30gz70qF9udq9/kv/oqhyROoVYD53u7rid2Vt2XEQi5
6J1NKdO+oIluSzkGRO9BcewWNAyTe3odiRRLSrHd25E2cnBHH3Yp7GEE1BFRv4Dy
0Qi7h9Mhkc+NqXepFdyBt0+hexXYPUvjay/nrt7O0deZJzJuO7d88bpSCWnTBXKk
faH+d+9T1R/cDKpoBtKY6EhRUEBai6qZgFN4956b44TVhX6Z++FXQvtq0ULQxBXO
kZNlgk7OZHTwAL03+DPHIsUJDQEjBTdJ3MFvsn8UJ9eQCHgCbY9AugVuZcJc6OnE
MAjVqquLH6f9zlNqpdqO/Wi8H1WMR0n9BB/8aU36FpRoJzVSKiL8l+IDYj5ROQyn
g4OOyR2V4i7KreT1ihk0s6WZFKt7dZYLytEkjjcsZrSl2HHao4YENQxsBt/MoEvF
qHfXZHW8TKG4lr/d9aOHJb4YIfbLGu6jQk43bVYEId7AuV8PjQocZWE3QrsE4vdi
BVUPYnoy8F1Mt+B78fM6SKGMCrdBktjlcEIbwNyaX3qpYl8quS9JfvPdhGaSLECQ
lEfLj4GdFIRKyPFYic4ruZqILsbpYt7gq3N4EkQXym/KrYYsBddB7UNX2zGJozw0
Mz9iFwFohd9d+T7TeUYUGF+AucnMcw1rPm1xfIuC9CRjUW2QAXCkRf8fUTr+cVHp
RRb7ov2VdfiW9v90rXaTgqUE//CYCgOUtt4wECorA+/yPk0ykr6q8+S6PzzsHzZD
Sr3YIqUtDSMjfdiJmBwil4Sz13C9mYKfD3GRa8hgNOuv9HXpMluVVcnBT+IiSVUf
DZjzhhYha11IAaOiABmrEMYLS+jlDwUyIjXVNWjJolKDv02+vZY7NJecWpWMI0Jb
bTVVKkFxzIzpk6FiHwa8rm+Tio39HuaPRRrh0Mg6IDo4Strf7m5CvsK1psyAvFRN
FgwWDRdsXevNrL61r//I97/NmG7vzWhXEyBtquoeXcv9vvb06T9K4PHg7WLP+Gyi
0CXZLFa17p1QNiEC5CCe7cAM+v8kQSIQ1RwrS7UrnQMvoYS9ZnrS2LUd00benZU6
JJBso/7NfOUaCPePk/v6G7YBB/cuxnVjB0Pnfoty8BDdkg5DALv94EMm7V02STA8
WsBUq51ldjPPsa40zGCL9S+guLPtDzUBTl0NZc8DeLdxoATZ+RMZaT5UF6WSYJ2t
sRj6FnQ0MyKMyeezxSUdxXHp6rj4v1t7wzc5KPad9iZTpOZZOJc5L5QFB8Bi4jMW
cC2PXxOw+ntxL+e1ml4hgQlUKoEOvh4uKoM3f8Sf9nNyDeLzOq6MluiWuLcToQ7s
7rRWX9zPQz9GRcm5VTqt+O+l0cJKZBSQSirzb6rhX5gWUfIpZMfCYmpnDBtJriaW
t1kq3KWcDEHjio9Rb3/SCPiA++ym/l75M+b5Woms82At0A6olvm+0/44smi7Up8P
8B+GPjvT6fwEAFgDiMagpNbtvkVL4PwCPOv1Loq3fqwsdRg3zOdwCPzIs6etzqNb
lujSEm/4ZakF8Ze17y0P9yWXhe4RILzyeOTfnk1Y6q+L4ECrYo1SMNvI1vMgCRU1
yAf8tK2UZeeLsvkmszIuc8zOqBbSEepTtNfqQADdqBx779qFUAtpIc5yH0wh9zqQ
dGoX1beCs9hXnzq0AdpWCAmWZJjZ/Kw3r9xXT+qwi6KEBlszTuV5XmlVYMXApqcJ
39bp0d5cib0syFQZUtkmNrpXAMGzdCFE7VRm0d+xcAILegcCtJvNhLL/TQc/wBxH
rsBUHp47dSnYbbUzp1VIxJDsoG4nNI58h5OLvBImVRBT9PcunaWqM7wnoCZj2wsY
m51qHDI7PqI0OiAt81kGYRq2ZsMLKyhwvhUILNxdojwntaB984F329AnOle6VPyK
gidHjmrJ9ZR++snAvSFgwEuZl1+dqhF9CXlDA8HtmnOAOBfNn6mMXpLtv2R55bYM
lt5z62Ch/7fgWfXs1qT3ox3LxB+/YY4d3EX5irXoIfdBqyQbKxGOQNSdoMIomdBr
Bp6IgcGJY18d3JdJlafSN5LiqTyDDLcs/dHblzj3h22r9d3UCCoeDygXaNl1IZnA
pqHhVquOVfWuCPrmhf7YgQO5Tp+krBPpvtAM85DH1LrWo5R0ZLj2bm/OfWPvmPpv
7qCIHuG7rxgH5HuiWRutJ2GtgKsW/YqDYeZFz6BrfHkYfPp1frkWDEBKtYTUOv2N
4X1y1SITz58pZyxe+sNS6AEiAao9K34imbKEXGnO32ghuaQ9G6vPg50rQBPgpR4k
M7xnXNItwCLdXMQQcz7zZGERuPRRqIB5yG/BBaSBy22nTxdwbOa9XPfzgStZr4TM
o/UWirSWk0URLDMabT/LUVXxvOgRSGd+vUlSm50XtuwGp5dcnM9Lji2If8p9JWxj
mJzf3HDLjYXNw4+jQzMRVsV+uMonSPKUPYz7Ls1H5qaK0nW6T+UZRXLRpZGL1WBy
9LxnZ1L1RAiVKogFhJV5aO064zP6EItK6wJGBFiPWcLKQDBotlcSQr1pEUpp+Qn+
hL4XBW9+7cNSTXwi9YyKPbzydhCAp6DN2YwnAekbrSTHlhJ8ul840AR2Mm+dhCkx
MnjFJyJGUzgI61peaIZjLbJroabXzbkA8Q8bzDoUio7u7tTQtjNSoR8+egYC2g3f
+/1Ii1JeVsaQil3rJ+hzEkYvbkM6vzABdqePOPsHyuYU5mfJHWi06/RKlc4J2Zoi
tqHToLMSDHzuVa3MC4gmmnCbNqoJ3tDUUTqFv63ntk3OB93eOKUelqSnAdR1yoZr
yTkZXASv7GQROEpkGdwlmluNvVOq75jC7TdFM60N8L15B7AwpaewyWuhWAOVp1+h
zZcHgU27XOLNhv6LOyoiFg/r+L92q7z5E/CagndBeYFJTXSfxybbHVOp+Fy0zRPJ
oiVfc6ecy94dMw5pirH8lRIpsd6EgiF6RKhYRA3rBnd9QjZaOkJAmlbPtOwWmfZ8
13GQx+jC1eZ/fzHfWfuAk4Wh9OXB8DKRG+oYl41nhsO3OH1ua6xfQb9uAKQVLG/Z
g/2qoAh9MylG8OJjX4Xhy401OhwDxLhWEzySd4SoUpdQPFxjLt50ODOxEDx/V0of
MgxyGaIM1LAqIxIpJGEaNQySc/g4Y2FdbY9nGKbs+Gd0bd7LahkdmLpDSE25bOe0
ybnW/hG+uFfWis1sf8d2tZvhtEBiIEZAQoXPM99S0n9M9uHRpkZ13AGd13NPwX0j
Za3X0trgpcZ0Fg5kDT3RfiUzQE6tDhy5lFQejTauJ65U0VcOjubydjrAHZuKXFmS
9byCeC5mkaoFqueRqayhoRb1t5KnWPgigjJqOo4Bkg93497wuZBHefiLzvA1LGLw
v5oyTiNtJssAWDa8zvbI7xTnxhAVmvdpDOK4LHxTjr4Drm7ummEKmYX4dsYIZ/yr
4oeEx9SfC4yiY0w7J+2sIoNd18E/0vx0E+i4l93rrSppuJsjEwz7g4WzrhLS4o8P
XiOtJgYU8vpdt9ZoWRHBeY56maj1ZwEC1S15J5z9tVEtUhU9cRV9G6APGDY7myTI
Z11bDFndZmpYSyroroALGIihvAc35MGGYVWNpPbS/R9G57/gARboJYLuzLcH4fPT
hltkeuELL5O1U2JjKRkKM+ob0R+HXNC5IQmbq1p1wMONvaj0+PAxLblMyb52mKXB
wNCH3Gk5+cdCW6vu3C20SQF7KYB2JUdnix++h2IfYDapbmip8wn9HoZ0tjiCMCaZ
Q0baaMYmZH7DL1e0Dd0CTPuJQMKvkWuqZ+O2AJPilbGuQZzWnspodcQcALtAGnNa
vtpIKiDjw2+50EFCa/6WtJIOi1eK7cUJf8QbMJi/OYSbLOlbDxx8Ys6EzBdyHJJm
QNIz3yj4vNbDwCAdVLGlcIekv/kjifkcr98m7x5AcwwfBZwtcIXp3UT5cCG7yL74
IbesAWp0mZagNEdklqce5u9HfEIRFcg1loctlkG2yjgoriAySz1BdtrPeiAwb5yk
0F8HOMnRXpQVCbFfQq/sAxzsHRzP5O2WPXhQ1+/XgKh2hVTQmktUCGMimrme3NZz
XMU6y6d0zzSwK0z/zs+0R9ZPD4IMRQru5Ar0mJsIKLiPJFpW9+HU4pbu1O+Tn2rs
k5OJeRQABwnO2Rxp01Pys3cmpph1cSM4bEDmRfrnuODuZ2phvNpr+RSD8inSROhF
MHTtiY2wre+Y83sSYoRe8ecNzARCDJK26bpkpt6LzWuaSQ8ln9RyY3gQylgYt2bW
4a/IuiJmXbI2Bh8rbHpHchcYd6W2EYweINUOo4IBgAIN18weYf2e65rWavLQm66a
5+r+AXF0t95mtIzvJSKlj9gYCQXhu+dml/uD99+t1AGXk5nfdf8dq8vUyKAkpDMD
WQyqKNe6mVknGDJlHsyWxH6MTrGQSKQDSmK1p/vxb8HOYAOcXdkdtlQ659Q01qh2
NZ4tW0ZcBP/Pkja8v5nVYsiARWUxtR+UFGZZ1BPhuswS/OsH3sIbumH0tcQ2FAmb
3502ZwVU9RcbN4abgEq2H4uCbC4YVhBH5WnRZhGitZ1ZNOswN3OF7E65RCh+SqL8
3zRy+EhTtRMfXGPG/WG2OuOjI9z1+i70UeyYdrEPZgtjwvmdLwqT+vW8678VXQQP
br5uyU+9Usqw/evDU1cv/d6yn57k5dhVJP5AdZDE3wAGsI7PknCbggaFuddohn7A
9Q+EfPP+KejuLutZC3HXre3N/BYpaH59clBJ9MEDYLLeM4YYrLANCLdAgGOZDnzW
I3x/+7FZF7wGrKRje28GzGP5ENvhNBY4WjRN3mIm1R9/uU+PdnwhPg8s+z7mUOvI
wV6WJ4adc5k4TbCxdyDZJU6fE5Xq5PVqqMotA27fUdemLiCoaxmT39TEUmuLD5/K
0n+UOAgp+kA9OOCia8GUE5kAXujGOwOmAdDotvsWH6BhX6q3hxWrcDhbdAU0fDhR
4U4XfQDV797scLhjPA/McgcY/ihhyVV+ebDMP9xptu8JSFHZEwfPoZnxh9dMh4wR
w6k+i01QCKE70VaNuJZqon62479KHlzyQBO/n6EOa7tEIHZXDdUHBgrQJAWuGsDU
vaNt7WHivshrkWedLEgCHVXN4+XnK80Gkw03ekKD4bgXs6dLki6xSgCppDfTk1Ws
GTOH2fwe6KwkUJZ0SewGykp3tLpyo5oFicfWuWmzLqmmpcywOBBt+W31coyeHXlT
3UV0XNCpW3vmsZsDPs+zvvJrY2gnSH5WhZG2O43PSu1Wq12bMR+S1aTiq0Viw+/x
5uMM/yhPgOswagnoXHpTnkvuf0Qjy3U6LAtKl8BEmrTN/sdsYjzSgEvrXxlPyTnv
I/K30rv8++jN0dtqG7Laa+7z2K0kcUbFltpJkfLxHSmRRkW3PyU7o2cixGASAnjp
4mXVKHIJQoc8X7Ik79e6PwlQYm5riJunFZegsUqIlIATn9uELGMaCyjJPoQQDK7j
HfO8Zaa8NcMV/n3Wfil/oYSY+G2DqqOC/ycD5Kr+KHsU/j1KYEXOzru0PoscIERl
x2p9cvfuuS2gAkoXYvZexgtNdDWT6lcbRgwLHZPxscg2g3C7tayIp4ZB0HHqG12v
NqKDwTRUF4/XvjWfDHOrc1kux49riZP2x5A0Cw5LzsTMHcmrDObxG3YR1ut2N36M
rBWKIckX+O71o+mC+Dw1ToAvenqJuaqqfXoYLREDsesbgtA4MujkAaplBJA22wBS
3v1hAuYgXPMDGYAamZs2SizmvOHg38tI5XZrdc6hryBp6erNc9q66OWOwfDvsowC
6P3cMg0LbNkeZE1yeFvdQLLee0K4rE/STTaSnhuWSqvqm0LZdtlfug1lXNYKqeji
wQunJyngx/xAuOEBnClynw6aoXR8Sz5lbwQt6glF35Q3ZNpmhelrLXaISYEMOa8W
+lEDV6OFBFID15DVvmLmOxR9bqnG2TOXvQw0S+3sZctq5Hc8KvtWxmSlQ1DoQrGf
FtnParFzWo9MABMXxbRGnwf7jFTgilNtb3pHDju1ZusgwGRpIK10hra0D1NWPfXI
7t9AuFzyku8e5JmW38VYqlHggQz4ugNNBmA9WAcLFDcQRFlxg2az0F7i/KsAvMBs
lRGXIIvldssNcU+Bw485MI2S3Q4Sg3LW0wcAilFXLAuixgGJs1/3v5/3htx7wrOl
oKkxzLWWUDvuqaxibbo7v1aNS6lZE1/v6E4qnp3/LM1zLWGz60gH3Yt1RawZtGUG
x/+LA9FC/OVmtAER9q3dXFBBnseEk7be4UPi4WMUC0lw14aBTPuYjZxge7OMYPyN
AU6UENNu6gPshRArT9hfJBys0BTKHUMA7xyYmCfxqwxJ4WHNgIzmjiE0JhLStCjC
ClxQEnKi8kQkXhtWsT0GaROce3pwQ4QM0PMsvSYYlx8LTOBx11EIUdRgUqu95+pD
qWFB0f9CEioy+J15sKRe3op0jPE5GMpaTK+zPPKrF6S4+FsneJ/1uaZEhHZcl+KL
UgL0wtmqBmzV8ouKMJZG59Q8UbwNmB+8tL4d+aFIfaNNMboQrKM1FC7aeC0iINx/
62XtsN3t4UF2Cj/3jO0kL20O3L5iN4SsZbQ35b1ePxJuWVnK64VIxboFCG3aDnhT
clfnsu3vpRa5UGzXyFwGSx5y/VFdmbRDUr0AuXPNe683svvXveK9ylL5b8Hc4FKd
ZV0YwxT5AKsUmBeOx0RYzaX6jmdg6azWPUmks69cnVKsAVua9siP/Ay5pTClBTxF
gahU2CbJoc4OE2GJI7LGG5kTMdmRMCYxgd0+rht4C9876U3e/svt+E0SbkdPXcZy
poyMCmnR6MMO7FNryww7YkyQbYxtSN8yNIHklxwj4n2j8K6RegKiHZyu5N5bb7IR
VYqI3EljoPrR7LJSMF1BnmNYg5nJdLWU0fXDJNdn+5NFQsOnMZIOR1mf8Lg9HCJa
ttuVOJ13tq+lOfpeqQAE9JDRiMsBFoiBU5CmIFziYLY0Q/gxXA+9h2H8rZJAvPCt
ozq3VKh0E5KaKK8ZKdTTAvkpUr0W/2ZYy5AsWDf+XGCo/IU0hIJQiiHHaqvF13Jv
l5lRkL7wJAhVnCf74ytacSELMA0e43tWmfrTWCthdYJwg+r6WQ5lxJCPNQhza525
SdRxbcaF4QaCVByOjVFKdN/X12+8IIcOfZIwurqMXojf7uam/Nvwpo3nNONc6PQ0
c8RBqrEiSPXQnrER0FZa8+emtmJ4w/+pQZqwIFxGajmH7voyeTOhTpbnp4VCv3/o
PKYtmJUpXwxogNWK4DX1e6Pqy6PcOko15cmk60OrOTqUbG0raBcJW/+jwUP/P/lZ
JTBBZvjzsB3JRtfO5b5SV6ZAP/4KJXV/YPTHA78d0JM7uIvYayKc9GQM1GynF+0T
GuDCDUf3KugxbkcKzaD/TSfOOzno1rM7mlUrmWm5azfJffTW0CCh02SjI+VWcBQA
Du6d1zVNmfLhbW94rQHeRXn/f5NjYKUWjL9E6ccy1wXEaAY0QZZ3Zh1HRC4Rpevp
E/TNDxCWUIHSy8u7FKAWzSszRxMdmkpq21+2yzaTBXsdXOgMJTJ65PK23ZOtu8WK
kP8YXARPzb94FxhDUwO8Tpv6FSjPbDVGcRXwVxUwhQEecXBhe3o2XMOMLRdry/Qi
saTVHlx3IfZ1kJizXW1a7OH+rjjmAmU7vYKa8NNSOmX8YZyDpsOoWkumNyTGpcYC
sCn0AP4JIOFnbRUmrEpteVtcfcyoLGiGJ1pejbX15VnmKT0ZPATxXHmhmqjJgcYE
O0NOeM4UVzO36jW8zmtFxnLYU1vHK6ieR4acy018hqPZJV0MhD1Cv0JciY1xwVX8
6SPlhZqPSUggeAvjJGsBvUJO7t+BNa0lxueYr1ts/cZhpqDS5emSX2QMUeEUPIht
EFIW+flAQ81sTOX05ngqSZOTsMs06Nnt22cepxE06XrGINh5ifoFEQsrvnTdzpQm
7to/zbyI14cgaBvsEjvSVR6iTAbuxRpWI0geDOEOV6MmzFr3JrmLpyu3VGnmgILY
dbAzSEiOjthYfuDMemxbUn+ZzlBNRmddfdTRiAPECOOFul4Bs3A4JlfxyqOiJkfn
OJQxBLaM2uhXf4Ub7bSvJDjJdIBKKLyvd9ChDK1PQAhc3Nw5JBNTEVL4xeNN4eSk
H++ryOv71ERIUypeahg/NYrg2a8npt5IBfe6lgvwOjxK4k8QHQs9tM4HbTcjZb0+
X1gGNF8zxhJb9CkqaqZ8D+S87DeEYQWXy7D9DvgcbQEdPhLexnsK1uFqFSES5sIA
hP/TQGmIU2wiakmls1h5CnAa0Yby5I0Iy30V1raGre7e5r794c0QR6WwsZKHX8Ve
IlC2nk84B6ibFyeOWF8t4S+AVRHtL7XWL4HCIP4Xl+YijJOVX1SUHCji2Eqy/ZDF
+mNPiiWuV4aPalretToGUy4ZALXuKkSnT5onHVsXKclE/bUeC0ZJV6W30me2tPOB
tsFVuq38zm+RHA6153gDnLGwxv58VwYYPLszFoJkSLkkwBCl2UHMeto0jdpK9Idi
NszyhjxMAPCES07ROmYx3DZOgoCDAI2TspztMAU2VdWpYHRKbNwFdx3RMFrk9OJ6
vXiw40yARlovYgern0v/jzTbhLPkAcsEfdJqZEqTN7IGZX9tbq51u9r3j3pzNpMG
FBGuWh3nE1f6rmTaMA1bnhTgvL7nfWtc3a8Ed2EIR+x2hQNf5YBNf7oIVwMZrABO
Hy9rGXJe66wtoXZ54YFaVyAYlN10h678D1TrnVrFCoeZabt2WijeZIuGx0snGOnL
DukrQEM/O5yaqBkUUY1W9UM3LXGqOx5ZQXwjSMa7fI3WjHN4rALNvC5uqkzaEvUT
l5eTH/8VSmaXmEqSwS+i3UQmNhY8OrjNxX3nltTl6X3Cbadhdpqmv0gfu9FF5Nmz
r+8V8mqgRtWqzTef4uTg7EEC2JF5Rllb+x7PQBWpK0G4JlGtlNryPma/JJTrkHsi
/bEy6iyaX6RyR0SG62ocv7cHiPrEX9cIhh2nvzgla57MnJ5Jj9YjkhWtCNOKqx4L
Z4W5bG9F8JcW5N9rssQmbFtbyLupHETdG4Ch4fU5QvwFD9NZuvs5owIEGpN7xYas
Pf16hrbiHAZ5BYwjNtdOrBnnjbEzVIsH4WSpcdsieaCzXKQr9s5SKTbeNTLB2e8D
1ofKTv2wpcQRK7QLJTUfD6gm+lWbFm/1cAHuRU4jUH/tAUgYTQftAbNO4X61DMi+
kYlkUCQXpgmLbUDahA2OORulbSl9p1PqJCBvOHxo8Xnk4gJIYizQNXEQOSy/CJZu
tKNJGvJl7dAWUigCCg/8mBqHS8ck9s1vbwcg9dfNdHTmkWBZWAcqBwl1rxeLePwJ
sS9OMhucgTFOZ2km7BiBGYko9i53ntFpe/5uPU0oCv0kLHV2l7e3YaHUdUruQsTP
4qNpIS69sEYopi+9AM+zk15b98r1sx1sPdyuaaQOM1dFhsl0qGCmam0icMDM4xqt
u8ljyU6mw/y/8CjxYBwsAka1FLSvSgHOOHQoMqq/JehXjo4vzqw4Eo3zxnkgi6Yh
AFCoCRTmfe89K/Upp9EcOHX5A3/Jkesxjd125GJ/ev5ELCUdooXKbrp7uBqygosn
VxeJjvMHRYx3mCDS60ks39CNrYczLF9+W7DmMk3Gelf316MAgBlthuw5VTP2DiC6
qx6WXrn2MmbDZ2BBjDPBNsQieSsC8S5INzhpiUR6DYgpBQtpxwdAklSTrla8/TLF
13FLp9vE39kicRydHv2zkfyXKNQC53fLOUufDxLhj+PWLLgEnpxsXJWYlZe3SGbl
Wzaqh0INH8Fcf3QKuKZfy7fZtdSJ1tcvVsjI6fjwRiZP9/aGDk3uFUoIZ4XW9h7t
ETXhAy89VyuT+X2BMyvfox4fS0eF/tMjHQUr6IA+UJF2rm/TDZCbfFLoA+HwN0mu
b2/OAKp1Q0NMqdK0fitc2zwd4zD8qjtGvXHWEX5fTpTdzPw1kS1ZIfcUIO3nZmn1
dxpu8TIYPOA++gmVSkZjQe1TQDV4vjqOs6bIvrE9OX3xMcEDl8hAifG7NVSwkBRd
g+as8HYyTc5fteoheyNFk/SclRdIHizAgdRNuQcm/UPCvv3ErHz1Uzgqrbigsbci
/vGaFw9EFih0zl3/uPzgdCC6jKL9a30OUg9aRfmFUpKhmvalLVgp9pUtTRarwYiR
wbHfII6/rSO22U70/XBZcXor2UKc2kptVuT9jZ8J0q8PVwB68uhDI4XAHkVEOJ1/
EF/F4Ht6f/f2UcYh1/WFomukaPPJM3cDEn/cwiubEeenb0OJk2UHXyT4zr4qZ3yd
7zMAV/UwLKJahITIHkTSviGPCZf/n7P/LbUy0Gt4uE+U6mBX8liBxQujPDwlJn/1
UTUbfOq872Bqe97WBi3HUik4sVjdAjlf0ouXd71snXlSK685vF/hChYY62gafppb
DzbEamXBnK+GM7M2lvnUDpCjC/RzXrQPqqY0PBQoMQ53//gDVLsiiRb0o6Xx5K8n
zmQmMuBrAVan0r7Ca/EDu4Gi/Ksq7g9OdHJVkwAoLRzudWT0uu3T6SxfGgMcJZQn
sbMrpZJtowfoD2i3mPwH4Mq/4CecGCg/apoMYoKjnZh9DyUKY5EdIPb+XA1eHC6b
PipR4O6dYQH+IteBOPIrym0eVN2kRdEtERiPiWjK1p/gPqAfEb9Khxtek/jGHnbU
Hv7KydXLtv8r1rSn0gspz8c0M4LKHyxXt2hIEgtsXLmGpnXWX2cJ1ALXLLY7ePCb
6lI3i+lxQAshgoX8LAOfb9V2jB/sKE+wtjUb/MkJDTQWn7+XeAy5wbthnjh7eIOy
8c6P9FXYciaMcHMNOGRyrp3eCIfgXHCT23fVBIv/KPSrzE5UVYAUTP57jLaGT/7p
iX3Ufyb+GcqQ8yy7/LNdd0xhHV7Kz8VL+WYYi9qNyWoIUxgQV1EfFYstLlUvZBQ/
dKIUDYiewE1+ylAoyK1hgMxat/6cV9nvgViwf5gXyHpjkueptLeE8Io0XjT9w+07
3xRpp5J6NdXkEVxahu8maatW8V2FZT5OK6nvRGVs/kFu4iBw7WofTm+InwZ3DwV2
yhSzUeJq4yUBSf9Hh4YU7pkTVVTzFXdWsjGPdN/2fpgd/yZvf1YHxkoUTdW6bi6v
iX8EZ8qIMNECm2cxCDNhZSrXdg7Al08bMChP46Pmm1InArEHjuVP8VfA6WzM3Quw
NeLqDvp+KD5QrKUe4ymSCz1LClKaCXhQteVHLBtODpR/y6cd7Zy23vPTe4zn5xnh
t4xzfEod2e7Ci8Zv1qaiFgaXxAiobNc2l4BZ2GIp1wcbrKOMYrDF4zsVXtFfT2aN
Dj/OghRxDJcTnqfGCP5kiPLrlhoIwOXMSd7mTOJWKd3jNCLWXSmE7hIt/eILS+nh
JRytlTA7kHWu1ha1+vN3em2u0LC9ZZCmx8RW7iVrJUnGIsGLcCFtHIlk+4ub66JP
A0Yd6PY29l1gZM48EnW3h/oWoRbSPSsycYSW+AcV/dvlfOM80S0sWBq7ag5u18gE
kcPeG7MWOFthLgLuE7YsGr5UFI/43zvtjX8jf2lxFTacz+hxRa1+GOpQSqHJCWND
wZorQnGD4jCIawPtrvsT4QyOcwfhU4FFdehxzg99Xs8FtOd07zQKlibUCo5Uy/os
Aeh+9KDNWG75ERlGC8gzIWwaTeGFjXlws4xJAZ/NAxpbtpAeoaSLETAt4Wt5+bcF
kJtrGeTsi1clqfZRyMABu78G46kWTB7Fcj6dG6Kv09iw+l0nmJ+tT4zsvavdDC2z
pnjKzsV3wmdM8iuGGNIaaxeN6TiBqqSYFeC/oh8obWpLl8awq4WL3oKQnFZF9/kK
HYTN7R0D+RoTsZtUuutdo9EpFfcFAkSJDeyiR28SSxxkBXvzFp87uucZnEU0NWzz
CWvzNgeNHvOvI3fU7oc1nHeispuCxWNcc+Rn7dcptfV5rXNAiRJTWEx24g7bSyO6
ucJNCMwIE9sGwwAeMKDXn0J1pKEamAe5mZbK6PSKfC6nfRlC4Z8ykrWZHo7vliCP
otQvMaZzr5RPfR8YmTAhFDVizfaiSjwsIOaU1gk7bTj0PNyZIqa6X4UR5Gf7esQA
/XU4ZrjtXcolvnQUM6ZtlLSzcKq2NSMEh433GebiILOoWECawVjewRKmXyz9VaSS
fd474rK7lZn+BOvC8N9yoSQU1tPKChnUaF+gAxw+GKT1f/o2HbLtTXQaUvVBGnhF
8oYWGCeR3QCdrHZYfNryAXawyCxIOyN+0d82rY4PKve4rT5+kAqmb56FIGuZVPJV
pccVkXxvBJEZKvCmhYYgOSQK/9jLT01l/o5VyAzMdkyNRJu4ljSFNA0NAPzxhB/b
wwtWWTJaV1Y2RQwXWbh5zCMNCNYsmAfwMXLKGfsKXQZFZZYBsUe9EWoMRCez4AlE
2LavhOKGa20vGYhmuk9791zhudG5bABuzvJ/4vUl2OWqUnYSZDyHXbiynEdXy8V1
+ao7PumlXEL6hpBVx2z9gjS8w8nz3RSeZA3GBaOJBZRWl601tHW0izqfFKB7Nd9C
cEOGk3vMCp6dEckVow5Ly3VbGM52uWRLM4XDoUKdXx/AohVMRpXdGQ5U3zvn8NlH
DerwaSNFBGfgJjF8o8cYYgCutGvml3CVUPKv/YcwFlHxlF4TaMtOTu78GtgCv2GQ
TQYR8cIxzCl3GMBZ0aLWBgsM4ByTT7f5OarkwxgeuodvjDL+i3uWjQAontujyzRC
Um+K/E8mW4RAYgMIxuHJdwcxEptyi4iR9rSbnrXftBrGWSFdUETPwaNR5icLYyO/
vsgJEZF6i8YTp0v0dAucgOfvIire7jsiMaPtS+T0YldU4E/SPVygKw4vZ+IiVVZW
Yz9aKIucjsLLk5LdWkYB2GE1fe82YrjgTFriK/zorKZDq6q9KayUIprX04knuPWP
KedXrBx/dHm1NFKN53MOdjuxzG6Morjb5gLjS6mQAOCL8+TyuIq40UDqeALtRn0v
pPk/yz6Kbi3zfkemOQYVA/f/60HoeUOovAcKHziCnfsg2mltSTqFwoSBemynCcXE
NDsb/DRZcJifJD/DZv0YkKGkOT+w73kNNzSIY3viR+sJZVHAwZmw7p2W+Olyb45r
gqDyR41iykMSVKBwrmLdOGsGE17kyv8x/3Ec8yM1pbo48ackEWsbqQwt7BsNZ6gz
Sx60Qbq0qtlAYQ3GBPj/jeXCD/FDvLeIIgtJypvomZoQxy9QwZjy6Y+PpnnYFCiF
/n67Hl0pwuV/3zrTUbYahm0kG7tsAaYEPxqKBK57aHdpImt5NOsDeidoR621A4Je
fDEZBRnn5d3vu5q8EWUILMd/KLekGFVN3Z5Q51BwHBC81rRXOk6kmsAcgD/ZipUU
upfJ/0Mej71rf9UmAu70igNa0tVvXlS6xUYTJSLYe+cda3rMNq5R1BsKPfcl7qI2
W293dTGVAj3/E59zFuHl6T5E8YbHH3h4STLxjakpnVmHIpnzERx2BWW9vapaOspw
uMKXBciQcKoUVfhgaOKa3D1GL0kwMTbRlySs10q0BWZMXOvOFseQQP5bMx0Nu9KL
ao87qJVfwCviliCW923IHQaL3pOaS4hXFZB1noltsr6VHi0cDE1tBu+we5Pge9q1
FJCO3K4kyRhqrd8Oe/uSeGmjUIafh5neEarMaMHYtDcF3gnu7ReQCRSwKdA8bRCn
ZI2n/sSpCY7gHc3K2c4nvw/dy9Dv8viapOp3w6lwvJXA9IkrTNAm4iyX3BF1VZAa
SAFf+WTvDQ+D3y5d+KrqC69ecg51UUyTBjOheqttmv+mcd+Wcnuc43ih/KV4cjMx
ULiNB2uweluyQsdZIcRzokQBJeRLmF0EEgs9wJFR7ijmSdidRW+VjvJSTheyXQvj
Sw6KEDLI9JeOZVfMg2t9emENondHjOv5Qgxu7FtG76R6NEfqNQ9SFCdPJo/euL7q
wC7alZBtQRkEiDnfeRidWt1z1dhkjhCpZKt3/j1F1aZOTfLI90+HlojuCkTEUFib
wuHKycegyaGqaQFOzTIMV70s7YimzsaqlLyTdXacO4Yfrge/KQ0No1l+JKZvq6vW
H4+QvFM+M+R+Psl+/Q9qA84Wel4kAvu7S/J9xPtkJfVzbxoIx74xl7Vg2VVl04Rr
34BaVlgrCTeFWRtxUDuifQ65vuP0ioKebnKdg4hYQMN92z0zGR/Nl5oDJLB2wyq4
tBtx6g5mYWUPWczdaquz/2LaCNHNhgjqPtmwYxAiEpgBsoiZtQ92IkaCFoaQsEs8
jXGadP/Fq5a2J478OfGpZWcvfauOhdcsDwaLUCVWCDYSojA3ze5OBuqI13N1saPG
U1sYPg70kTyB25Yhh66Ynmf/WY5DIOecYz1GtDiH+jQv7OduydyPNLchs4ryKWlh
USh2kkz9gIXkyf31VrGlQKqxp66asc9cKs7Lg+qnVVvUdb3KOhjSe/ECOfXlBY9D
AGcV/QopIcBNnmpO5x513aot71pPHKOw4c9htzKza/5i3SSZs6/WR1stWtcrtfUw
1RKsk3UJWWKpLRW7ZCOPY+0OFZYjyoDJPNGQ1XKe+GOKjr9p7x8n4b7RxV9lVUUg
Qb2R7ldEuMJJIJNVGx8pGnY1pVuMRytJzxDcMLodY2YLR+4ATs7njQ74gUjsjl8O
fPzZz7eHrYMhvzjJu0mIZCpG4qR6rZDwHB/KOodwQX+tGbnJDbr13LqgcPQM0Yh/
p5qjLw7lIB3GGZuEXWTxHGiAsXwvdVY6i1KEAft4xRLBbLiUHTCjNwUPUXpc7LEf
/N4FLKnw8pJ86+c5qFQCbP1wNxraBXyPEq0BlDNeykbrlmNmMqjqX3joaXUV9ULB
DDTRHKuQIqgcCK0d9v5VlCtAQI15u7qe/mpvRyAJOIGnIQiAy+pqFNwedad98JpQ
hUQxxUvMKj5LhGo6YXzS5WhRYZ1Ru9zisEpiqgbFvANZH9nkGcc/Gdb3xtb0U3hb
ePOVLjzIazar8jP5BBmBZrgS6ELK/N68nrH9LcQNsHPml3MIpyAi+U1FAez2XjKc
Eopb3DEn+MkqNTgwKuSUuCd+wKV0URAwECgNB98A5ti9CWlyG/K5JXUNjDM3n+RB
3/Yp31f9YR6D8g9VEU36+mPSdg7gKfEPKX/supZRe4Dtb2zdSf+hqyPWgrnO0kzQ
58g/YNwxG6x7XciMupGU9yfK1CLnxPzJThHrLw4FEzymLXXIeaYVc2ypB62TFAjz
cYo4XEP0CM2XQ7+zD5+VkhzXtcujOSNY2WjosvRwUVg8ks0IU8biB/No6l5jwyXp
Dr4NiVbR6a7EdKflmYteb+/iTQwFiWIFEH/GDm2+/8u41U9WB+YK0ADQNrRfLK+0
/WXhIxAOkCkZj4iQ6yXnagFkumjygThX73NO4DTsUcrr8rjzbHC9yo2xTlnbOvG2
CXJuLjmK9QSDj7ZCjmH48XcEDQlsmJ+xeEjkQvUqgBd5FCZfSkzq4gW8utfDZjSg
6PWUyk9TxRYcV46KBuxDjYtljL8vrO0MLo/gesHSZRWBC2dKeOy1iEvzOBRVKsTZ
SUJXngJAi6lJ0e8k+NHAtOYNJdC3UhExUweG13/Wt80daphhCh8+zZOHQl4OXe7D
xQ3JI/ZWVGfN53yPqRC9H15KkwMXkW3zWEBnQozD6TLDDwqvbqUmKQLtN14cGWPA
KhwjbcjXFAUKN21dSStdtveoxGFhLauYvp8tn4YKOkVtcvlbfrUkMinO3+PzSzr3
w9Kp7Y9D9VLXsvuTmY/z2eLXmkifQO0HQvsK0tBTG97qSo9HwDOHcyjVtIHZ16eI
XKahnu46rot7vewCIh0+W1jDHE4KMIoE4QzhAtR27RTCNcxozjYCkve/2AYbdsc4
Tr4DxcNYhvgQWcKSprdsahiGhUEpmLcrv39ra/B64nEkqWFfSqwii/1T+m2yspsB
AnfJeUgOZI9+ChcS4q/khTc69kS14NKn8wgAdZLY6YEl8NnNqr3r02WHY39Sl/eQ
TwyBygw22/DsEDVgGNO18MKwnazfYmVM1c2akUl2e2WSs1vqPW65txl3UsnAor7W
dXn8CpNXCgopBfBrRdDIdmCz87cPM1Yve3eB6QnofEoHHiVAAcB18XHYVnM5LVMn
y1bqiSJEoKvvKhdgMzzcTAXy1CfTrj+cvqJX8NkJ19jtvBxrU3LvPNfn9KEgGfQy
auY6ECjNPoR8KkNIYbhRKMprEXtpxPo2bZShbnZ0vg9IRTBCIC0H+M3qnK2Wyhix
fzlg18B/uHFjEd6vtUrq9os0uVXf1eoEi1hPVLSoGwn1b+osOJcTqNNhJ2ZaWF8r
lIuNz/R7PMs5hjbAd41tWDjP//krJuYDdVgzWiHAlGtHY7GrqIFB+0dE/gRTOtUS
Cd+o1KrpBd6wBoNuZ7MPzRNtNuMKQ9XwM+vKThXpxQ+TKZv1T2zVtPYw4cX3do3y
E6JSabscSTwRIeLahta4LeiOSZfXmUctJn7Lw/huoskPnEK91Wgb1MezlMcT0WV1
ClH6iuZJt/+663+0aRflnpG55PxLGvKRsHVhxG67tdgW5FFtjyly4OW/Iw6lWvrp
hZ2vEUDsbraRvya8HzRMsQuTc1yBJdXbffQykef1BoyzXfcJo6FTb5F9rCXKJtuM
iODuiNeEbniThMCybcNK2C05Tup6KvuuoV2U135QtlDCGSRkmspINuD7kIi/9qSL
rge+JJ5aJnEnLZvLp8jksKhNm10CM7nwGAWoFyOCZUpfVc1XN4u8awssQyK9QCVh
QvSxf/rGmFveG1EykLbJEROM/XwYu+4lqWb3Qn1zHDEXNiSGKFLt+uGTVT/CtMla
trXiRqYyqRHWv6DMqxnDcjBkfZqLpNyTO675SMm7a4ckeQ1yNyemlMvOV2+oeRtp
Ub8ZFMDcSdaVpu+neOenLJ1ROaGPx2eBStGroULuKslbs3d7csYW52jbnaAusvPy
8CLsfGGi8f5W8yKoca26BIQVmIDNSO37zYonLPdHi1vrxmD0BidGEBvW9avu6hZQ
MNIlNSpSAaFOsRA9i13G9hZMQj0Qzv8IqxFxbFKfKymzgu+UOV0yqfglEwl5pJ5x
OeKIxopa7SDnjSu9whRMvlms5I+Z3QOPR2pxNkaEpcrH+G+LiDRgNO0Cw19KwyE0
ueBoCdH8rthrcy4DojTf8j5cScbiEpGt1yIGoumltGTDOhAiPr97Vx1wGwudiSuf
fOTTcSNtA7HG+4d2GdlsO1UYrY5P+bI66ZerGmajc4Q3/7jMyS4cLCDI+JV8oxHm
79b2/vtVa/E0QzlUn9ZPqvE3hzhSARi9JSYMY6vc37UjjSkgwety3Vs6g9yreWXm
+UeN38iBRXIQq/InhBUFAH7/j7OXsIan6ZGwEffzhDUqjvO0jYfGf7uBSOtmj53z
leqi/pfDsimoSsFLwXdSjcT5br33Wra/1ieXsJs9jvlyxjtHmJQjmwGuKAjmdF+9
dhpG21eCoCRBHcRpiicOfQerhncrDkt057jPquS8zWeV8uhoiAlEmQcjVTYpy/8v
qk4q446PxV4lwX8dqwos0+n8anrThEU5I51GHz1o7q4CDGYFvCkcqSNsMkRzK+6E
gXDGCixYMD3mTOc9b2IcjCLKbukJxrukT9qF7QZptvaXKuegwGkiwwE2iqTSIFbZ
xZlRTAMbZzmx/9umoru9f5SnIEg0PQPcq2mjrvFEKwR4DExZFfKCkk60llvi1jn/
nLCNdnjs4SDePe/Kj7PSiBhl5YvolaFSu75//MQT7jf97n7nyoE7Pm+6Co3uibws
zx22qzbdtDWPiCtOVYrB0h+6TICzvIoPuwAp6ymXRLyKzN6Gqc8C60JDSzUL7VQo
4BMHT7UaVSgGfj5LiiePvuHJvbtCd7DWcflQODUjlIx/ZoSnYRk/gFJ9RfuEyA4Q
wR39VyUvKWIXFEKgIBJZmVDJHlYWozAJJMT/mgsyNZDohaH4/idzLwVXoE8pQ+eq
wtpCkJ5TbrKMYr1oLNUgHiHLFfuVSZKCkxGOS9BHWsrDrOwtNkGyDlU2Fix4ZoWB
8PRsc6fhwExnq9eGi2uSSvml/ERCjpqh7zOkdrW4EkPUa3X4EfOF7XG/bbLEuTDD
Qz3bl1tuFe7pLZywqUOMkaPs520Ohu+VfHiSUwKEcMyzAFc/Kz+6j/Y6cgAWvS8U
iJlwUczZ7zYlCIhQeqSh1ebvunyk0xBUTrJd5++P/e5oS7MFWhd3oMxauB3c8LJ1
cVj/4CHPHY1ArF/OzAhjodKGJ2Bc0f/YQSZniw+B6SF0fpPQ1SUZn32PD840U7Oo
jxZRqFtqMdyk1+kHdlIEUNkorp6QqiNodJAug7osWQwADRVCBEL07Xbdcd8+8tFh
4PEPvX30lpWup/aHPQ5g8wKdjYKZdpRrwGujRkFRBcLVxzhVIg2P7v/iwDb023eM
EEp06AH3Fm19qc4x6ol0NNcBrhV6xazucAJtees3QUQP9mWqK35sFn5X5tfp9Eog
fpvcAG6fWq+jUUZl2E/Nw3KWOwMuJ2BZMExUfwUWpE0BjMdLPwHKjcwt0gW96BSN
ew2RMvqP51IKsMB1T78wZCu37pWyVSg+seuAt0bYW1+hrTrOpXs4CaKO4CuGjsgI
2iF6SIJkFBxmNoJVE7rjvi1Zc4pcXJ3scOpKneSRib7hYKrBKVP893xdT0kWmY8H
C1t0Uheae5YIwN/Db7Xh2+AaEzkfO4zvWWsXFo+n7GH3W31Clmizz7GU3RN92ibF
J5xru5SBAxUFL4YPmnkSDM5KuYQQOOaPuqSCEkEC9t+1n+DWUPKgOTCxg5wr8yrV
fRwR4F2kVeCwm6FC2FmOb5fs9jyC1soJlF3qIPcs4pxpMC422q8PfyDtIf/Cgtrp
7kHzzw14T/PacHd6LOU47CS/sDil/kV7m/GnPZa+mKPvV3HAxF1r3HpuevEG8T2F
R5Myn9KnQIDYpl1/vW2CX0+J6xm4BjY3DY32Y05X6xOsV5pcb3iKo46KyupNRrXw
hGNNEfarnKCKRqJrIoSLcDblDs3NpDArAmWc61oO8qnYmfVHSbMj/XyWnY661P6T
VadaUNixpcUgQvV6keMf7EBTgnc/8E82q8kymHapP5Ug+3mcKBNgpOV7WkpPrCi2
X2vUF6KI2ONRwq7Z2LsEEhpXskmkZ+CNccH5uGV6EAeNaxmQzXKl5zd0o9gZzdka
NCLwO1T6pMDOqyps+CGlZzNGn9bIiJqrWqZOw05YIxO5FUkdTpuPDO+Z+HAeFmFB
drFfUZjqKYWc62bMVsVCLGDc4PkIyFpXJ9mDi1FVAYtX7CanKFv4X4js1NXhXgVr
ImUGeGUPSAEjBH8A+x2gS6ymauImmksOPFlFd8O0i8dFVErj0XJpaOnnTqYOYYGX
AmJCOlqRi4PfFPQ2wLm/OxtAy5aaAmCo9YeOf3wovnehkjTq89xTQzWQ+qArwrH1
Xb00/litwl38n+MWUIfIc5sqs8Su157Ap2P8hWC3yGQ6me8sDAVhiuqb8qfpM7H5
eRCEydME3IXAxHY5xRnp3gpxSpnZkcYeuUILFuekIqnWdxg/ETpubis5zZ5p67eg
/GKkdi1o1zDHZZbyMkYKKnBmXwW8MhtPDubm32YXj4JFQwqph6DXvYaGJSK1dmc3
6ylbIHupVp094ZwFmdWFSYeDbKuvZ1cIjVIUNs18MDp6QdkIs9lWWY6O+JeFM8/F
jN9PKrijFbRL5DtXm91yD3EScRndoZXeiheguV2IvugSgzr0odVf5X1oM/u+AN31
duIamyGLyWxUT7C+lAYGQSh4QaMWgq+uKku2KyBK/gpCj1L9NgLkWb72Z/KzWmbA
37ZXk2FARnIsqQyu3n3+Csj4a0uGbWTeoTzmClIxujLexJdN/i+L4hYj/xN5oH+4
fxm0FM8MImsh0opcxikdgoZucuoDgsM+9KRkSavCO3JIr83iq2HzbYu1ZQ9qfI2y
4p7fTO/pwah+axhRfm9i1rN45FLsTU0fdwUv41+VdXg7myjjtGlS707zko6smsin
A4wHoCTCYeOsiRqpHIdyTv+c4J56Mc/CuU9vehVbWW4CLsmCGOqAYdbdJJmROxuW
8Q8lG9lYluVzg4hgRNWTgOhjFxzRbRXcQ4U3dnYy47GmjS+WAn5gdUNjXBmWU0l7
mE7GXXDCElTD+ZMG/J7T7lhV/5MhEFHubSN3f7ya/6SNCNiUwxONQviE1XV1dFIZ
joZRrFnTpurMw5k6JPXgdFE/IA/VyFDq4IdL4NTMMl6FpztzzWGOmnfWVr3co1J5
7eGkI0qTgTHN93P13bzGRY6PqNUPqSEy+rGZcSwfkzUmcKEsPmbMvgpoL+YAK6i2
atf6WcK3L/9iTKELcu0xYHvPJaEYj1RCBlC7Gj2TYB7f4lcPhGVX70scKZI4KA+Z
Km9AhCZA4EPREcfeaSrrwWOdlaDkzZLWX8aKoC9Mf0TpVeHNTYdhtz7rH0OKGpfU
my7AUdHy+m+OCuw4DcXC9bDyNsp69klx+NB9xjAV5GoeCUNfDOoq6jnpDYQ/ddWX
htAavHWfPB7W3kbHEvuWnncQArAH/zLNGYz5+StL+VXb+9M0iqUa2sET4nRs7CX6
UaYhs1Hj4ShSFnAFCm+uWn07yerDvuhDffcVH5zbw8UrCsrxxnB5ic82lpYckHJe
MZ2oSVihneT6b/P4m+uWrInUdS7sSLKYw+6KT1pltNYG5xFaxyWMuktWljI2LJo6
uv2jAO0SeCBuEdhYVxiapCOhdtSAaSrViPTRWRthR/ZHsNNI0A8n9QOsFLPLFrY3
kWl6uxQhOy0e+WfSj6HyEphlWqeaiJKBCL1RtplXNJM0iy3sAJzINMYwqSgT5AxS
NOZmFnFxPbZH+PBfs9EwAT7RgQWS8CHCy8k6Dt/n/pcz/yB5E2QYy5NMXoLQ4as+
dXISPQiUjR0MkDhRmsFl0IMEVQ7hKmPoLTUkMLQ2eOFPIUIGCaL8d2fXkOEVmTbT
/IyNDK7SiVVtCntraV3sDYgkddmBdflTBqRoS6oFJUYj1/pAe+oLL6jYu+x8/ICq
WgCwux7wFhFLIeDro0bB9U8hi0l5cli5S7SXkWzlOAgQuoh7T5Ib9OaNfayjFcIg
/AGC14OpReuhA7c+qERerJhmChVQdL0TfSEa+9I5ZkZM663gUk9ztHGaboUJYNex
SfBSkD8WKqBkyjZfm40joXRtJK7sfghuq1rjvdB6Z5xMrQLRIbEgxEagaOSRnhRI
MEk/Fa4134FY3f0XQKIaYdOCSzAoxV7mNJ853lcWausDLaXtFMORHqqZkxwV42+0
VkM4y+nEwfq29hyMGvolV7pAWXJGEf0oKmaD9SgknbhSP+wqu4wZYwBI8JMZsHlM
qhS+EFg+W4Y2OvJf+LvqeaIlbVQpqGkBlyheM6V10lUOF5wWmsZw6gwQqgoAVIWD
TW2evpB1Ex9oDRarHjNBcBdCZJXqUANoltbixxfv/X4sZNIPOFpB0xzBIa0dcvoR
W3jZg6SaRqn3CpCNLcGDOcnLEUCML5o74NEZYk/6OaEJoYn7ArAll2sd3rxMHVx8
/rGmU1wMgwxVMjel1T3rAVwtBFlSZFPMbYTlCwQQStdkRGZtMVraTeMZICYQv8W9
6bQv+DsRkzZ6avMAHFKwBs1uTS2U7WimoJoa5Uns3jVwGxDvYTC0M8hvFGuJXTyE
ImWIHvtClNjeUBg5iFj7mrJuPVmueNyJMmhEXwUphJgI1XoKV+X6Ep4hWeQqwZYo
3wZwyQn6I80Jg8PZ5uO2gkbK0VgEM4QeD3zdn8qnB/9aIb0Tg1VNtJeEGR1WQ3Rg
Ybd4w080P1+Jk59Zn1c5q8K20Kg4Kc1oPmTPRBjHp8pnFFm2zOe0SN9mQ0v006+u
s5gbQfwkYootmAhlE/kUqU/3LdJs+YzaJh3u+YNMbz3/PZ5b7zGV1WkJS6BBYHt1
cg7THDXilh1hcD4r/C8KWn5J/LSjRk0AfnqMZ0w5eB7cSGL1rs93lW1sttcTThmJ
DNqBpiSjI2z5I2Gh5m5uJQnjQ49y9xM3hlSOOt338nC6HKaPtslnDv2sZ8XyPA0O
wngDAg6HbPhHz7OPkREFHXacDBbmeSZ8elhNYdz5Q0WtC/rm0nRSwX3f0Gd7pmqy
U60ugxv6Gm5Ha6OLMZ+wk4clliMUefoF6z6K1vWozE9JZNrprUnMbK9CIah54ffY
XmbLlse6R+tqLgBsyUv3DBPYxr4B3odQXNVcgNtEGWsaT58Y7+w+CvxVzcMnqIjd
JUP5eRl4/C3330R/1vTFvLD7lnSJgcP8thL44TnvOFRFtnlNDO/18ZAiZD1tRVNe
1RgasyqOXh27oS3Dt7Jp1nNGWjATpyBBAGDbPW/mdglUHPBPg09Jm9vTOt5/SpKh
5qOwx8oAVWXzv91QTq4cbN+XSUxQALLIZm/wRyAHsVzlQQiS+l9OmxGeteQiO5ye
iiMZ/N3701e5e5KrvLDPq0nTwj9NajKEi+KD2a3UZMRcEFO9154iv+y+4/s8qsKL
Szd+Y2yug5EWb5ohNg59Zm0ceicekwX3UTPaQR/L6s0Ob+zuMzYn1DtN6e6vXwlD
5WJadgbPpBKl0t5m98XOrCV2JDC+oPKvdlV2msamuwrXg4emegiwM/3kftO3x4MN
BM7fW4N5rjZkSTMARs+QkRtmiS01wpfIM0M1sRFBrjoUSCsMXVbzQOVB4prxiex9
y6mt6rzwtsJ9X/jqjN7y7/LI4vsvi0Nux41Wo+sWwXlU+8/BVstNRr/AQ3R+uNE+
uheMbJxmy5fjNWTAyoESEPErUZ6Vx83aPwzJdteCtFn4uHyCRbQ42H0YR8CHA5Fo
oJsVwwObQKy44tzH5wZpyBWBdbjmsOeAMZ8hhVaGp4RMWH+sg+qAHoe8ya+PYDDG
YFFar7gmw2KehITrXnZp/DjrSfrMriXK2z52vNFKZ0QL0qsHNCmfwD8vjecdpwQ4
vU6DnFP2r65xSXWae3KZIMX1t6dT2yvbEed51QzIjaxbGMLDalis/8sJipMoZ7n9
OffwqbdvEVHYaaDjyu1r02rQrtc7papR5c9DKiEnfL8Z4RaelwEkO40B0I9s6X6m
97uDdMYz8JLdyds1XF8Br/W5KRu57CuzYtD+OGmN4EbcFFB175EWwG0SPEu/wV53
bUL9PYDrNwigINDM576lcZYPDttlwats1+Hv/C2fadjsWFF6yFg+gOGb48SE6Yyw
zhfm0eGlpXA9ZGvXPsBfwYV81sjhp5vDlODxdhmRnPpgwjKqwmNyxk0vjdlHZJ+x
CDjLBYEaBoUjR2oq/VI5+MyIcBWnTLdGvg7uyUU/TuH7nVVizmSYZsYlsxizWLBY
9HPuu+j2cE1PApBnhAYpcvqnZQfD8IT7lWPLStwQlqCCmZLxYrqZuzh73LiQtBCi
zAfbjjH/uSTRM4N1BUD3KHNnv2JP6rncahbk8G5tZpIecCOR+j/MuOzUt/686cya
rzz9ja5777iDpmdwedpEtOzU7IOgweM3a1aexLounMS9T5RF0+9HkgbvapoZ2+vt
4XDo/CwpaaFwTLKb6k6i5YOi8GdFrrSPIBl+pcrlASDeuvxY7WNSt1BEq4dE9w9L
L5GaCZYwXZ9e29g9KYsEuBDc6PuR95IgduokFnsOc8IHZbVFJKnHfwUlPDBaq24v
7Cw72fUOiza7INsosy1Mf142fOP0goNtYYvHzG3DMYX8jE1Gv4Ajh9CQtbm/JAqT
BVaQEujIV8QjkCBzaJ3yjMYtnurQcuS3ujvJIT/xaqNb+GU58XlL401kuVKmrijv
5EI5G45b2VK78tKJQGpyRtzkvcnhfsfg0+aU/fJ7qBH1kGeHAtP1wwSOkWL8fBCD
/1rCPPMT5jOYpOBFbpFjQCExRpkRG5jGLi4avkx/DxJo0kTthKjMVDBx9YpaaV2/
LvifMm/ZwEY19ZG1hrG+Os7lpnzDL3SJDilnM4Hw8NlCpG08CH5iVchg4XkpdO0K
4Slf1chFU6wNjkZqw8W89PjOVvT8m90geitJ191YsUPe2ED/u9N7CAkIS+S2k/Mb
P0v9YXQfzQzSTRX8I/PPqk+z+6wv3DY+pxQEqE4M3TUT8KhsL+E6iO5AV1FzpZYU
pk9GQ+sXallYhuUOUV1V2VDRHunOmES/aY7oHm/m2gKsS9zIHMWqhAkl2Z7KEs9W
L4mqsga2fUz8YSflooL2E/+x+ev3rB96rDmhtBcBXIqXswUkn84wjKnu0LaxeRw2
aRch8IhD0tXgHWsrK/hl+nEY50+WMRxcrqk4/EAi/8jYczF1prRen61YkudhEVhI
eGkogmhQsPKBURQymn6ACMwV0rExOGoWSqjf9rM8TJtouFQwv3xrE1+Z+5usWwAL
H2vZ8r3dPf4zFs1L34NfHOOTbVt3WEVY/8w6txOThmpRpVPta6/WS5TqP02om8j0
cIoH3hqgmMdMKSkVwEOo082YzyZXoS7IAMet2VqmGUnYJi57njMR1hTu+duJ9Zht
e3OgzMZ4vESrK1scJPYz6j/IjSHDu/ke4PbsP7lzH8xBKEX6oXnSxDHwKI4NDv80
0vD4QCWSmgBbPb/zw0opc6FJNk3RaOhANZvtZHDQd6TjBxyjoVWwp2m+xPyo9ueA
vIYzIJvR0/DANewVjR/Jv8T+NkFO4fSXZimNPisMOAiLEJxMSSsKKLlj0K61u2F4
2IvbY0F0GnIrWUoQJzZ3ZwOWjUSfvoiCZ1z/oiT9pduIswHyqw2nrH3C0Ar5dQre
8WV8S0TUOWnP8SOW4jDt0NZL7A+FMXN8dDDnSL0+0tRIgANlv1Cl5F3j2Ogxcom3
Z/pEceudEUVOu5ZZNA0PV9OgkJd/md3QHWkxAGvcjnjNVRCsDM2tp0yZD1qSEftt
q3KcVVeIau3ju7jQ52aFEy0g47u4iMq8xar8idW5c1H0MtgPZ5zME717DUt4xa5O
zH7Pp/YCvgCKaIMGd9Byzc2t9FDieCPQ8UDu+THBq7uur1003x1BrAJMF8tb1pU8
wfFUv2JkfNOTQ5rWOPnyaeCzbDBD4Zu83Z1UrfxpkvJrh5IQnMIWMCd5Q8KZy0kE
lfS3mbSiGATrxVy2y+pEcieJsYHELUVOqMEJ8H+0bcXDGjZHMVIdkdlw82fbPpjd
L1qaiKR+Af+/knx2xDiND7rhlndRIV09Xw0Rks/3ETdGYWP/gbdAslIfwkj6usSD
svOWeKgqM2+ikWFXLwtWCUVrR7BfBoEkzOVlNweIwka0S9Z1r3BbOjTPouH8ZmUx
hrHuQRlU6eOmEEOI6io6vaqzCXjPjc2vQJ39sh/R0iT9hDqH0Pcqm1taiSk6gtCT
QUN57a3zW4sKQ+UK50tQ0jR/3gDE8sPzpg1fdTCyJ8tp0zM8Xn0dLagc3gFj5tIv
DGH6H4GPRHgtDKfor0azuKeO5zOudOaW8B8FucGrdA+8Q+1CUAfGMhxd+BVW1/9k
1ccs00fEYvRwnhEGGKh0nqa3C5exlOoRCv0oNKTcYWUSkKDxpNjDuEF8XDKu5XTi
Itfk/JNz56akyXRcUmTkdlTT4+owvNNMTk9d6Zs1rXc7YsDYXm23ykP9nWILbP4T
UTkKd4sDn1DZKlwFFql0Q6wMwRqpOaasK1+7/wruSPUBuMgE7mt4CujFTyWuzXJ0
oUIt+yui9cgmAuQg9ptfWHLhWeGn+OQM9V1NJbyN4yxD2CNQ85JVIKr43Mlvo5vd
/o/WOpiIm+yv/gbaCK69lDHOaSaeQHDKIlynSQmE+0CPHAXroXGpJy0qY/QkzySX
04u8e3SURaoeQuaQILwDAHClsLzwG+ELXjvMtkCY7Ho+dJY6DuQ9RmBfyEl5Xrdg
Zj+P4ti/RjRAGSc7mPg1ZRnzAWDnxZH9hlUo9mIka/LOmGe8OYHGO043r/9SIaFP
T9zGQNlpCM+3yfoPdMM1BifwuY4YoW91ZBK6qDd6U2Q6gUnP2awPk6AeBa1r3bsv
UC9bjmc/sJqPi8NpmrehXMJp1PMjCq+iUN3/si+rObf5DC+BHPKXlS9MKyZngTjh
8kMZUT2F2ZcbufTa7gjnKY2DI+mN4EObz2/b42pvG6J2M7g+BY8rEPl2fJ1QRolz
uUOTGd7CiFAcglRmiLCx6NqXLTlheH6pa12niRd0SYNoCBYOaLumggt9CuYo5OYk
HfxkF67jNRwazS8OB8DS4qw/ghG9/xXhGAotQkrNWOdahosuAGvFToWzto0rJvCu
I34DaaK5EgU/YDPXOaTVWISdrann9Ea5gGWKUmzmPMrNFucDB8FrPsbXJEcijf0e
yvJTHta6qKA3JinaDsKBquD1qvanes1OGu7oO3j3sFi0J2R6/Icb7R7XhIuqL6zC
qjwRLaCrTQEYvvbXzdq6zCGp9/qezNfVpAI+mFP3tJPngoenKii87q0+W6EQVWB2
RoU8APEfNbixvLgJtHqdEz/8m6YaZ1fW9vRv/SK/JbQJilKCeerJDhxyUyI9+58Z
IIwQsEtr9SLAslOw1rsl+N0632d08xiPB2tZDO0c7qRsVRPaI4K1Lz8jICSNVZ9P
8nVrnnJ4r331Lw+wSkcgJ7gKxhu5tlP7Fa20KdiL8IUy4C1nI8ex5N4hrD422ioB
tXOcome+rf9ASgUB1OgefBBR7PQvnNOt3U20dFC7WVRxiuR5Is/TlSGjgLi/VwN9
39RNU+MZP0F0WM4hab0OYYDIhK2KYtuq9Pj4GSJa72CLfpiWOrwKQdkd9JdQvkjI
gsfxkDrJ090jvEkYQMEvLKNg1JNVblJ6NhsWXdZkqwuteGK0USySlnq9UkQoCbFW
rxe9dqtJnSKbF1Ra8YgyRNrjdfLsULtGxS4o2g/FcEw5uk4vEOdEtDVt+aIxZaNb
Vb78nbyLg+POi9VWaXvCeQdj7EY11yZom+Z1InzsN4EzfaS8Uscp6YNCKTmmtpKj
erCB8xLp1QD5aOVqMfIdIzic9QKd2SFSyCt0nMvhXT4ugV/mY0vBBXYiS2cF9TVF
xiPaVdI5YjxldbHZhy4QwgdobELIkcHuJTAcLjlNooS8u+OmOvFdkGJ738/qFDxR
VM2VaimEhKr0oDAdroYsh2rNQ/b2WcJvZxeLejUutnqdaMbW1P4GwVf8pHKNsfRW
4iS9rWkDbjwzLu9zR5PDfGky/ttQJd6FRfqSfm4/Iu3nyJk4bYDHLDs88IOiZPW+
vxx7VnU7YcV1admV0Gr5QyxVeBgzuIrlUU4VKg82VJTwMJbatKThRGzhZAdDBvsG
3wezA3Eywk52C0/zgIgWQB0kPk0vodSc8FbNmvAEVsSioVuyb6rBr0HUEowdz/cv
kmxj6BhAg0oTE2wIh5mHHzYkBrXRmINnHa3imQuzGxQ6RhHbTqYBa3c9y7g2HOHx
gzc7p0qtPYnsmbfyxnO7bD1zV7wdD/s5580DECGy8t98+Pml48iC7ZoxGRmPfcTe
lE7Z3DAvwRID5UqBeFEgv+oXQr4cWvrEwrbkSiD9mlW35ki/xINNUAjxHfWjFNxV
0YhMikmPGsVWpJaKYJIt/0R7qmecPMx988M9eBs1QlFIkAKSvJKz1G2XOTkURbCq
0kcLW0cKpIf03TIzl32bN+TmhqE4YpukVGpqdsT2vh3dG/XUhpiQLS2UEu1ot+OP
vgMjT6K+/6zlX2BcTWTMoJ7Ce5uqG6jtzmWhZWJzdhmTvxOVPPgVGFZT6dOfN4qW
qbsYR9T6igcqwm/sMISkiE293ozcqlSu5+yfdC+t18F1GqUPLOU7uYyg7RbQhfSP
r9bskA9G2I/TLlfI9YPp/HrSM2vg0nYhAulSudBspWrQ3ig689BhLdI7xDhKuSXV
TYkcZiOrHPfb1nGcSG+I7ZJm+fpBSqKLdtcj/FSJfXjhcth3o+X2LG3J6bsOA/s+
W/frHuWxm5lzqLr+meKqv0UCMLPXn3i2BALEfQGKThuXLg2so/Sy4nUoqOrki95W
W8hjwJDK3C/5+VTDC6nFxQLt1ChMlnZajQ0dEkr3rwJ0Rl1NxN+A3LNnnRf1jbVL
W9qjXO8bvJ3fWVqsBgT05chvFDECtokmAwiZH7bhdwavncyueOehwkErWIoqmwbm
yI9iDomv8zZd33LqgzRrPe44Z/sM/o9SGaPCSckCo/OBBMPmcF146ofMgNfIIcch
GCgIS/qAO/uCuRktrn4SLHtSuLeFHvMmQqxz9VSqOFIHWquYcNE8/K6p7QQOY0Tu
vkr5VHPS/l7r6B6G8539pafxblEaCxmwuzPI99CztAGEJBEoHkaIit6scEx6QK6J
VD3NHCwb8ZuxYVYmgerXbR1CgUixvrC2rT17SDTE56Xh1PCQMFXMmayDKGUF9BcA
iSw/dkqi2WVfigztIOuCmmncsdYU6zlKBcOG3QSxRLqRJeD4Vukc7JONR4YoE8GS
2YHjvrf/jy0+T8Vb27V/M5h0t1vOD6jBXbkAM7Nmm8J05L6DC93HD1LWgddWjqSw
nBBTsd5ePXb1xHc660gwwvbKc+ubMq7rjgKXt/RzROgxEEZy9Cv/ekBSQ8CXrSV2
ye0jaSvHMXDzL1YvbDG0iRVHkdPs0+0nx2WFBLJEeCdfD6t6AGs1FiEMvUTkLHj4
ObcTvvtST9/ysxZ+iO8UkIVbs8uG223zSvp+igLccAfID4Iv+K/tMt7+SSt5TCOY
Ug9DBvl4kpNA7tMiensUCWJXOj4qQvhbkPfb6JD+0F6XrQ3EqUJg/wrOS5CHzp0b
R23DR9Rrja1t8kW9Z5hn5+9rtB5l6NxK8lZwZN6sBOfE4OUQnyNbxzoLOdGZQj0Z
ySb1Fp3S2RCRqrMlIyrZ4buB6pQ0T9iEd7Nz+XRt3ZVEiXrckI21FkyyEMyb96a8
ru4v0CH3c5WEoteJaKoqBfUqtkBy6QlQ1Ra7EUg4Q6GO6LxEyOzL1s70FOY177+D
ZeuBU8DzPphf/r2ac6e8ezbapxXUkbfVqHf6BVIUlbJ67fJYvv6zUAqIRgyX1iS8
z4es2wa7+4Vjc4Fsxmmkdw3qWzq5mRbghDM95HZWO292gyj0gxlH00RkqrC697UK
lhxjkYgCP6ngexeIh83Y9iSxfjbvORLVgW4VMwX1Dgb9eOvw/nK/GLGJaanygIsB
+IohbewnTlaV/ZrTvF7IVgjSXtZMZjaLjAAri+kk/auUCgGbNx+kaQHn2quTeJ7d
xpJQwHLzRAEWYeld51p7mEwohqYIUw2AVHY44/IBUMRjD/ZHVZq61MgccSUsGJL0
o4F0nqBjkuVeZ28QVuq9SJ+YyNuip9F1tUXO6jcgW+W0m2l5GZvsR7nPlVIV1HPQ
TZzuwQOspWIfvEczN5A5+RevawIY6C9NGq+1BmPk5adnIEscriCiO2vvHF+9FAP8
Ie5DYGOfIMa26wSI4XgNlaM6DhtkWmNcWy6a9LfZT7VH3UPeAFLfHc6fB1uLhcAG
b8fhG6HSsRF3SRNJ1/6Pa4vxUuwaZLixB1bR2b+PRCg6PJLYlMC9kg17CwphSXVZ
64pVi/fEAfdT3zfyF8NP/tBjMJBf6P29fp5RnnasofsqLDRoJizJAaCdPLVsh+rq
XokWe+aORe8Pp+bbEDrRFwJSGwIyh9nVYFZtUYyqTd5l1ZZ9KDWL5+WAa/IwVyJG
7AGm+v4I8mkbxAmH4cbmdd77JpX/KtJVtt6vktXTx0nPePIrtgovtpEPh4dppkG1
pTakcqIhHv+Vskd5DEc9yuQrylVaMvlJWbfU6NVXnKaIf+ZahEcF6S+IM+/g7qFf
2QediFiUKLI09essn44/Oeclsvzs0mg2Z9KSeGPXjNOcd7HAKZ3wE6HAb7nWoSZ4
Ualwxa9Yg91JpmJ6U1AYEfnQsT0grkgt/ySM8McZCrV7ge1WZx+1voGa7EMW2rJp
NvCTmTY1DmoV4FUyNIgF/OYwTHJMp4uKjTsClLNVBeRAmtZW4iNOsQvEnyGMKE6H
8oCAx2TELqWZLNe0ewPysvZz9ittZ407uWpZKdxvWTXHHWTyQ5eR++VUalENJqbS
ZtkAlJux6lI1r3wyKWgpe3AsYx0YMtRnu5O3LxqtiW1VmUOdNjSruQofhWEPknGq
PrwfLbQIl+c77qCT2aGaf8WC71fCfYcXBXSkxv9F04aI/PbJuZK0g4NRF2nr57mK
h6H/dMimj9CwAq7DGmykPHhwh65P/FHZFXdu2OfX6VQQ34WyKlfnjSTKH66BCQwr
meX4WHSpoJm5E2frY33l+YahI0xwisdnGw1t+iOz8Dy7ueDm016MoNr0y03DrRE9
1bXro17Opba2/fIrSsU7icUR/6psJfJDH5cT8ZowzefvY6GV6L4TsuVEGOAWH4K3
7zXdEqlRNWbHDfWmedFOouGi6o2dndAd8kDLSM1N97XjlqL3lyCw5HbMIpFRzj2N
m+bUNz2rDz8gfSUfe7nU+805WSfDghyTHm1JyDzpidav2eiVZ8huMo8+QjL8qSI9
EG8q8imYWQdBV2h7HJoPWUFi6L5APmwr+KwEod766o+3eR1ERVdKxibfTG42RgJM
+8vTBCxM/3C+WQynSFZOWG+XwAz+pp48J9pgQLKykItOUNzQU6pT1VZREnWXPBEX
g9LV6EkUXrmjPMKSkA95V5oga73ZksHTAQcoMZCH0nFrz5cqHJEdfXXEa0nPSPBt
pOjrQrD0rfqvnSKZ7glf7wI06Wb6w0ysLD/5oxjCKH39huF1XJy5QjglCZL7eTZ5
XnXJ7GWTrGNxPrxiiA2ur0OfZhBwiDdqvRqoQ+DyICc2wZanNfBudJic2DFAK+fx
/oQaaP+yjupBg+b2Eb9ySZcZa9ktAcAMXf5TmdJMTOrdk50AELndyd5YanGOM50t
jbwXePazMeZe2X4De4Jx77s0Qrb2Uk4hpNzYF2uzsqz1A2mFTvx9JRLAwWR+KND4
DNBC1MEW3MnkmHmpAeQ3+lhbqCZjvfWahXe7KSR9GOTIgxM+CP0hO885P8sAOjsZ
Q+9ZlDdRDQAT49KlmHZsA7ohvHwHiJKE9sfBYNv9HpekX1DbgNpriwLetOuUGmao
2paNXQpVEQtHAcoh9X+HZMfuJATLHkS1o0MDTrVrkNd63RRX09mcnvFTLW7/FyFc
74/X5OoFjC6zeRbb/w1J38MTTr3JunAowdAFgBU9HAPhlQKcB7R80nmay+GLNZ2j
ttporLoqDnX+IQSY4uRvC8ShEIyYgXAXVX69zY5ztBR7qoMPdXiyZp1sOdnExx/s
gE1TEyfM7aSvGg6yH/h27sIz+rKPRryYFJKN9XR8pSBpdQlI6lv2gyq4QV56s0QL
PJCY3rroteAlqbM0Q5Pryiv6ePx6AGeznpNA3eEoH4/b04Ol8mawITj7BJ3SrILA
t7/2I//A5iFj0GamBV0R0BXeRgshPkc8YC7VkYuerbAXsdV19bnoZ5RfPrg+RKqi
5gUR+ziAAcbivDfq9w4r1XRhDn9MeHWrW3lMK2gqgs1qX0crN3bizOj6BhWSlmOP
tptQmxfzU2sv4+QeZe4fF4f2UmAuUL/edzqdGEj2pVEP9AdbZeb+Qlv7htjzeXck
wQU64YCMvIG/qqttDT9wRRAYHftWPEd0dcEwE4zcU+HDlLs4lZoo3bPdqWxcfTiY
5UPg6eZjiF8YEsj1GAk+GVCfEI9wZuJsH0uLehHBLAfPAL0pgMEww78T1P1hBGx3
HgPBzZygqVDqwujTGf2toMAYmjAXTmWp2xZcJbHjv++TUDOTBxNE7GaeaqRBbbHd
Y1UGm7jxPyQ1stGh55dcpTL/dP3bO8x6IK8zBJjjoFkoc+DWLdFjsQBTubAN9vdH
Zaw0pyoQq5UD3CMhfrTx4AXoym+6YzDKt/wSZnudPM1Gq8uZqP3rr3VKDw0sv6Rv
+LSRw5R6ONfvOirm4OQwQDUs8806TAqC9u8OU8PBB7opWTnBX+E2ZAhbNgzR/4wJ
hyydxWFmOg8mA6dmX3XgCTV4EsG7zhyceMV53ur0bP2Von4mAQhXAV6PdPvi516U
QbgAQq0qq+RkO/6i5TBlrdl4xFN+zrNdkM+ehJ8rIyNtd35bMiFJzTSOTaeICTIE
stW6bPdBVzNxv8C6LcR+LSrFvhqcAylYxBY13s+5yYrLzSGqPVONzPURgVxrVtDv
yi9Wg0GqEoVRFzRXuFI334jiEdqtAFw4MrX13GCiOyjXtijFsItc6XX9Djc9Qf3k
idzrykG83FDla2kLCKpEDwN9fXKeyxcMj0BscLxcyjNSOoM7KIww5/DXmGU900kx
uWvwKjbBbT4oNwW3yh5gJ2ee0OeGkm7SBs//7lA1xdyjtXjufy2ybDdiHDOMruN/
uG6FGSqjRXQLInALpv1p8xoW3iHJykM0rEf4IsDMlJ7bGmxBK0ABb3r/zdOVG+Rx
ak2tYmkxFVfeiXz4mf0lmmAQMqGmKtYJl9VVLtypKBR5xPmELaEeuhlIfVsXoiMP
ilp8wMBx8zXAjg3emKe0WGtnV9bv69IAWRggxB+pGfUekcLfMYBKtw8O4H5fMj0b
hv45HWZVckuLJzfDxbiwa21W2ULRQRJblPAPtqz75Fa1ABpX+feyplSE/wrjAiHX
su6+wPJuZqk3IKDhcGIsejyvjeqwKujclFzmFq4aw0AWyDRbrTsru5lmW/4JGBvD
+0OlZAfAlnJLYnxWalrZYH2Q2PFgqa1rlOZTte10JysUwrPUulSylj110Eu09g2h
RV6ntLJqMEpYONSs/N7lh53XTs1gGAkODjrspbr0VLY/ouX4wiGpxHSxvOvV5u1b
eZyaYLkPgVtCA8UW/1p8Hpx3XfX5AnFo2otCdw82+hi07HJfiStLdiXcJcHE54ut
H4TrwJifoIdozrD+vHZ0d0IB+0Mzt8ach3/+95fPiBIPxzQ2DkvgHWBjEtVXXcLh
0U0oxX8tRJRA6gV5vYHV5ybLCEgeAPZrtYMuMtia9x+3ydUM4vEv5CXEzv0bsf+k
kY9xY5Xzp5GRqGE4jJLn4NN5bl6x5qAvVqZK+tq62V8tbLTht75h74KncHhFQWlX
YjYToRih67FvckhNT20nAmIsqawgSzikoc/Pd05vjHr3fL265F+Dqs2GgcruJxgV
Ll/rcxS1ycVlc5T7JrP3NSVOQC7Wbuz0mrCfChwfHwn1bXf8kI0wmNcR7oGpk0QN
rKVEG1DgMsInrq988g3bkb6x6NaMyhaPpT/kh6E3N+DpMy+G/XteO7++nV6FIV0V
eh3cbUmrkWDFSl51sEUpnJgPIp8NGHrpa19HoY5OKfERXs0qx5Jn4ePpDDuSYsxe
iQrPgmZ2vWz5vyKGJJKlEZyAOaLbUaEY/n0wPhRPvIDZT6y3YJtRr2MmLXNTa/xo
17KV+cda4grlYCYHOw5TCu7yJ6rk2XyUn1CXk7Sln04FzeXYmRX6v8cDa01LAziM
obB9vyBxqLMagmBCprU+QcbCDI0WYiyz8PYOELXcRq7yOuBXqkAEIgmljQIizK/q
knidlKfzYOsovBwCfhxuTp8dYyzLLW8l5HlUgKylhrtrOElLdcXIkC0uU5IE23KN
T5uuHqVfIpyzX+RWZRqx2gt2P60LdA8F5AkkKCFfWMU3v7pq33StppAk9VOwHgHc
U6z7sXn4aytc1anshbJWQ4EKzZ95lb8OKrbxYfC7va4gyMnC0aIr9+jIIimK3sbm
pjvADZfiRwMkPjfhlYrAVUQ5B8Z5dhZ0xKtxIne+nZmW6y+RII7pqEweXPHY3bnV
62u/ZBiW3c7M7SBWoocwzutSNwyOrVCdAIdRZiJXFPj/ypooyLKlFcMgR6C9Zfdr
1JaojkUbEXKE15mV6FOQ2iG5LCbwHxjKZhZvHUZOO144GIeoND0M1fWF3Y2++RvC
F+B2Ru7yUHq3PSpVXHChd0Vgh1Zi5XqMtjXdAvcHIrOvL0/v6YNdRcYhucled7bk
FOoWsnyokpS6RY0gdWVCzSVmZIiWJn4tWrzD3hWsED+5b+TRRY07zlo2+wAW9VQu
B2n+IxNOmiwbYpL6IykS94s3tcFrim1oYIP6ABE/VX7FoKKt7WKP/abss3GmVoF5
xVJmbZHvN4zDqwAR+NkLcaaQu9YcdiCb5v+Z7Dq80Q1qEF4JnZJlpzOHeaX9A/Cn
1XdjszGxr0yAhgN+ljN2eDU8ZboAmyoo5IeuklaLhLDCs3UJtUp0+9gHXViSoooM
/biiMBj2JX0pXzgoDXCe1gimYDMn0FqZavRAyBBIrZaIkn3DShZuU0zJEH5pRQB+
/TcA9ZPG+KAAYvzsSdrKwQ77UNhPVlKPDgryngUs+CMfUb/HFTN3vvgXa4e6tXBN
INy5ow1KGSECqtwWQ5llf0M6yVvLbi7hS7UlGNYqxBDPFdx9vx4o7Bzb9jSzpQIp
WRqEw39qWJFKu3hAKpMb2Hrq5BWmTQKAFq2d8PuKwTMKlBVe80dnnUYkkKqmheaZ
sKvtBqUwE2Z8cH+/zEObzZH/SPgazSAX4gkdAHhmqQpqcW3wfr7/JZeAlDU7TRfN
gUvV3eHwTzNbhhW+xZW3NcpA+0Sf1UpB3OHklSTXjsiWVVMyid9s4UjzYfyvQHWp
tUeY+pgdgVi2w2FZgyxDiKguWRnaN8rqCFVMQqiY4X5FkMR4Z+edmf0rAyp6f/Hi
PVWCQBKxPK17KrLz5WLROZwnXaRWGR3JIlcGXyGebX5nX5JAL4NJVAGDldCkXMJz
AKyq7jzNZPZnSDbgcRpJfRsPWb7lGRXGkTwkgmO5BtnO8wdx9tjt5WBpntbOeMhy
/cJwu84SGKWyvCp5/rtwkCPeSb+En5qv+L0WFg58tFX1QSX7CmfPzHx/2PWqO1FM
+q99+eizxcdm3sQR9v8jFAd65F0Gs/1b5uIebUqtu+NcpBZGLrm/RXz91gFcoxWE
ERMnlsNaTgWOJ9CuYAVdc8YZtUBUmAYQa1zJtg103Lptss+EPgAQX4kTIBHamTgF
lQe+U2lB3KO9DKGoUeUEXPK1K7wWnvX//q+AwGctfJb3ZFUgEzLBWe5GuVBJFfLf
7kZ6CsI8bVbs+ycah+e2tj3pfNK8p63H0arxdhLWaNXznXdHnt1EEP2M5L+NYipg
hGfNaRevUhMFj6k1DGaJgD2El53kW4K9PIYQD1pMdnhV4E2CaK5DP+P3V8OYRxsy
ohK/FsfFuFp82d/oMbHm4V4c5UzPl0o9EB3WctkJKKf/3RqCQhkp6JuBQ3EBIhsn
f8dQC/o9+AcClW8Q45wRpPWSFbaF/IVFV5Lp4SuNkFIUqMoI8Kz468kcjei+aZrZ
xm1t5s87j/GCdbc+GFfHgExVDtvAt1ykMC7+jqVHUQHf6nuIp0v02NdFRKsq/iEN
qlHNvQxs9QIi1Vh4WSxaHWlDnCVjrxykCVjL9FjiKUK/1jYPWVPvYCzyC9IJgC0t
x+K5xuB3VsnCwGhcc/NIVG38l7FLfv6A6BKR6MVYfg8DIfDVQpTViR9yu4ui2IIk
xaJN9oT9KAGvB4MM5K+LOKQLYizhowIrbe8tyhY2OY26llEPyEpcrkaSjZnihS/x
Q27HXUfSSAcEXQrbRCMFp/tH5koMZ3st67RivblyzPdKDVvbFEVGlJ+YBq49IWwJ
khOKu520DDKBzlU8VTjanyKYoNn7TWGW5sc+yOf2e0hDG1/AEyHwfWd1AenUxSfi
+bXNtwNSQelFaswoLKwkJvpt+Rn3EyMKJimts9V/zX9pmFW46mO3UqKjNelt+UlZ
TkVqbZnaRqZtjT+W5o8rZWX/jSsa9snDkoVkFxdql/xVMVgCZsf3Ad3VUIadnrXM
KIGC/fSdRI1Ed7ZJqetpiP36K6SngipvkQA3cZ4XO4v/ZugxXmOjWRlzje5qOymp
12hFVRfjlG/SMqA8gXl7kJUN5GCfrwqueTFwfE2nvGCT84LSWuKcFzAZVeG/B1aB
ig3igy8xaKzTCb997LQsrhZ4lBXRONk+WYHk7gvjjOGbkXFzOR4hbuiW5xRjjmcL
AVB87u3UwePj+9OKZ+lSfkfdPsPCArAXx4KoGlJnUKoe/elaVaXzOCbuQtg4Eem8
QiQxryi3Rocowd8PwmBfC2FOA/gYMlO+PR43npjsPC4nAAaq56ZGsEDq+Cyi64qA
QKyobZVtuQ5V7WVD425Xw+ttns09uD7pNCGYtHEq/sogTM1Wb3I3zBrD2i1HaIa0
xO1Pk0n53rlc0LSA26tOEY5vuRo9wF0kx+yzRryk0Z+xCNx6PVl4KiO8ZQ7tacTR
FfyScDQv3f62vJgOYHmITLrPiUraD/4FVoxUDeZz3UVD/0UyBslYWM84RUYGtxOX
QFJUMuOYVoH0xUxiHH6HZhXWBaTI66vDIFLH5brViytqI/v/SaR3SOxtoAExes9v
GWznSsofM6riNi1rqhr0nkSp5faCpuFSrfxtlyKbyWHq5KEHEfIQy3ws80Vb2PTS
/6w28ibyhGz6KaHKcLUzjUflwTAxtFBjXIZs9L3o5cbvgJcFvLap0RYSnW/RqKw5
jAasOXDwe+45AAYQ0qMZtp7iim5nU30KLCp1ae67GOC1KHOREDJ+sWeLKDsKNvoz
t5Ux37urBUY2R9R0q0mElWS3xbdjz1O5UppMqlKqVXlUuixPUsWWDf4p7l7F8baR
yEI9jkwicOkkLT2zmBLOkLnvX0f77t/vxi7F28xHGEK9oGK74kb6hqT6p6G7VPVk
xH+21twRbWU0AhpU+f0k9yzUy4P8quqJx8D2z7/xfrPwfBO/2xRGgLKfQea4hK3P
5zlUQ39WDQU1IFUhEFld1bZpO1O4rznDkWuiQqFq/lvef6t9pMJ07aV2Doi93DJ0
FJolGCKMCQpS5IBzEumMQkPTOxmRVXGNe9bWfn4wIk6xJ5cvXZVuGdAHrejPzT2F
cbkIiq4+bqL5WaDAW6EmXRl/mB2tpzfBDF2ihRXQZ7L/4Y74li4jze16443W4Ahp
u3m3ePV36YZiIfCbLGJLTZmVQ/Z9E3RGHhfLUNOv0e93EEvKzi97bJiKG4YDLXe8
q/6MKic5t0Xekn5QbQwChgjuhaY5kG/jl60otQBH4Udg1nCe46dG0ZDpYSgPvYMd
f8GE1vm28LO2zLub6wC/yJPMHeih9TjMjTxo4jpAAeSC5la6yiIMK8+KRhPZ7Hek
JAR39PTAINRkcI06Ap1np3aiSiHmIhlzLYx/Kv8ZkFLVylSRrvtx2Q8gAMfeXPra
GVk+MiiaBlsqtK+/AIk67KQZZBOKq32ZcltrybtMJ34QDIIqaBMXcuvx3SENLyzv
PRWdk8NAsy2x1hsk87W6t/4Od/ghgo2xFL1Zqzb1LsOTrxG4saDmMjj13Zp2VrAl
dDtvnvURVeWYc28wgI8eCXqvOALfP2yFHsIiPUqjphzkfBsfvMDYuGRQSXX0OLJ6
GGYPnRRxQh7rjtsRk8vCU/RRD0lbo2KmseZWih6wDjp1PgRnlG50hC+pf51cK0Jg
lWdnXJvu7wVFXakCapkZdXXgVy39IffY1L/VkafEmeaZymWtV39ROpQjnBH5S/aJ
nB6u3w3h+SZajatdZU8xMz56u+Msu86kQeY49pepUm3FQQDsmJiL75WF0bbJ2tvh
Sn11mRum0tXDUdgOlPGHaqN33SVGXwx4T7neOsp3qnm9Pdbtp8dQXjmJNbhF8jPv
FkdlDfrzDjVSMmYL9Dc5NKt1lwPYrK6EZICBb2DnWRamzkaDkp9isTY/EN3K9JgN
hbP79Nifd4RJr4Vd8vj/Yl0vkzWWR4u589FZAJhDg0bG8AF0SolVseD/gC1OlRog
pL/KUYWGl9F9Vv6Tz8WgwO7BZHtlrF5Vgm2CH+wYE1k1cTikxylYUqhfq/fDv6L1
KT5rQmbFoymBHeqJnbF0A/BCbWZjFX9HRQkKMhCsS0WfB7J/2KbnCLsUQvlGDFmV
Fk7kEBqw53BrDs01TWaoJFnkI+yHSaW0jOxkXIMLbkc1INcXZsiLkCDeJaSmQM+X
m4TvE1artmMQkBrDK0Owd137bod+uvxPLDoGiv0ovaDMGvCnx/NOVhAMdRS7Cunv
Wz/YNPAIGCn3Qkfr8FlfnDqLpd6iavjWdH63wGQFkLANJuw4PI2pzbQImzVzHd4u
QtXLjB5jg5qLtTtMBBRsqdGFF+WPW10obr1oRbuStXozI8YS+ksKqQ2oxC1vs3kJ
kWGNdviE/BoaHH2N2W7cXCb6IX1sXVc8PvHwfht5iIdqKIvD30DfuLUPXlH19n3b
Cd5rVxtPEfUDsNM76+64FTfs2ZrebiXXm+T0w60hfvAOo1QsXB4wl3FLIRDvu2MO
tbVVoKfHFObgQdhbEu49NIIKRvB9mgCqkKwNplMp9VZGC2NGbah0FBLUE8w/qRjB
LVD51T2NCphhyzanHd5CBW9YNMtKZkahAIz7wbkvnQJ7swlh5jJ9Zl2G8tOLc6aK
It9+AxtqjhwT/uClgYRgGgK7ZqJq49tSEawcwAMkqtwTg1vCBLT7Jn5vtL8HeR2i
ls1oLVFwrfLzE/tBkwNmmFG84DX0Q67nP6/pqTGzlZXXKJJ0Nr5ClAY4qTHJQ2mT
Fe5ESPfHkCRyV8WKI7Cp2VokSsJQPcpNjWpv/AxHrUPgWVfnuaX6jX8+/GPSNYxm
y+Ngiy69OLmTSqfO/Hs/+TMS/wfm69zx4iEpNw2cooCL/7OnUOJcUPtYA+/2CtC9
FgfZD+WWk0qDnVRqAM1A/9hxQHYI+7W7/k6Fsq96/EtyL/c4Nd4GoKaAQJhLBKlW
PIzuaWb3yZUsL6IFttj695HuDT4ap0pI/Jt91T75QLdbR0geZo4B1C1jarlcSLIY
FJ9CCOtDXpsNVeahJzmolDuMDIdI2pf4BvTi5RuRFzuFDbdGQP/F3f6gNKIZKeh3
rj4oN5whdUq/FcA/iXg+kaYj5cM9y+cdvi5mJRlMXYdohxLKL3TrOW71NKmXWDcP
EkzDqnOsPD0FIb7Zo9ns8SpgCXos51ghZqfAydwHNRUBJAhtvrWBUGLfD34xc/WV
SCvx7jIqJzVHi30ukXr3WDivFH6sJMa2WEZYWMgmQ4gomsRAMxn1juu4d384ZCoV
3j2lAVcTYkWk/5d9bZvtyAoeIKAOLsSAH15sIbwZWwjeKYfAUrADk5nOk1a8zWEP
dFfa4LUtsnuxaodPlMx9/eRen+xOqk5NssslSNvww3iNhr/NcGWbmnYX1hx3IU0G
3OD1EyhtLC9yUH0/1NUr70sgUI1IDOvIFxDbPoZIeKGbzxxtfz5VMrQXO+ssDpwl
/Nio70BzAaayn+9xzBfVtm3LS+mPp8nlowKSZKX96nR9o63e/x5EGjYovPYzuJeq
9Ad49fRNrI4YWdmzWAyerzYGIY80xEnOOuphusfHWf/CAWkxHdSZNHCY6xD3IJw8
+QPxlI8E8H5AS75VOIvBLE/G1ujfiAV3AJXlsGGrhh0YyO4BD7cmlpcuybhIfpLi
ufqJVFnUs3VpTkepagbMWkirjCHA5zp2wooMS1Kdg/DM5gKd3aWytuzoa7DsCIee
/JWfGJ/DMlccnjv8gNgah75j+Ek45YqoPbdT/c/faw/+KpITEdfEVLd6SfWZpNg4
IPad+gbZQ2xUihB6CvbP46+jlgd8bJptO3XjtVJBcKnrPex9+jox2q+NBSKUqYoS
2fxd+Hxj3ETr9tJSU2S2ol10BSh0Rm31CTtJSLE97rewAbrzlcdD9VZr6VWrJIc1
tdZcnhLx7nWvaa9QzUH/m5nkjxy3NPS0G7QtqDdUW3YFX5ExG/KDiZaRvoH08//p
iNfPIbWoubNzRmCvNZEpSwaJDZe/GtaFEZYo8uNlgmrCN4Qbx257UZQpMoi8rfu7
uJVd44N81/W/SfR6Aqi5e1UCWnWt6VimKAgqgyntS+5a9zdvLPl3w08iXna5rTTA
1xcXTfZD8T/aSfU3J0UaNpzCH8YsnVGBw6C42I+8PXRZAhumRhTnbh95nw/lhTCj
fvrC+P+yJzpvmzMKcadyI1q9wurDtkKCS4BrAcJApAgOXs2/3WdVJrt02MzXngiq
Ofo3AkwNTRPQ57glXNinuul8OFf51b20Ez6MysFk0Hl8UFEU0PeMnKXZAl/TpYBd
RBlGDek5r72PD2dJ4h4TE8SipkmsxJN8JwqNbr5WfjtSw4PcNLYn1GjnZ0G2gfYh
TbqwGzwXCccDAE7MQH2HeAxvl/J6nEMMw4vK7by8clsLNPJidz8NmAtzKL3+9l7R
iA/ewVpc2C0VLQOdxVlkQQEZ+T7PzsS5mJVEkhouB6aOe+ZVXrxtx7idbTNzpjpg
0GoMOjGav7SuVZGhKbXV/IJAOIjas3yJHEnEihCPOPlkplIqn8V5OvaaAEBWrTAd
REbu6aujoYyBx15bmJwD3zRaxVEjEjwYehr08qTdIJlEC/lvlinYJYY4h3SnFaMR
FzCG3UPpa5tLtP8izzAaCH4w8klbnDj9dLZWVlhs3PmrSMMWK0DYj5/IJPDd9/nl
BvgU6JAv7JOhDfGqBU0/Uuivj6r7/ljz6UMracankWyvvEPvuTNoySGSzh6yv1E8
Ay/XPKvTupOK+8nuvgt49vmRT9O9DUtdQGkaWbBsWuSJ58OKmyzyOa7bElmBAnUC
vXE3jzdXZi8VEH8/1j9HYx3gpnSRtOYxQBCw2nwYE3gsWnv2GBb3U4qykBEmjsHp
IhgvdxNiKwzCLJ1IH7wC8DUYUMgJa2K56dQGxrwIumuJV5TSbuPduiE0xRsu7bUC
4p1SQW31Hw0JDUfK94FHmjFgi3zS87cA3QBZ/dvqRnD8KphzZGixHKnvJP4LZeWK
HFfbBrW69hThbrlG6fPfD3ZX+qhgv4Nw/V7MwZA5Mozc9wxnaOwzLqYvrfKy8ZNM
soA3Qv4/ieOcsjvH6uoaAcbtrhlqUfm/GYbIecpsMdCnB+2sd2ttGWQoLCZyYr2i
8SimyMh8sl/tZVfDZ5nF4LE6mlGd8QH/qXLlj7DVxb/fzRiCnsOGQaepJPUJZNyo
W4zHrDCIpLrKpNcSbA/z2SyRlLGXsEDWVdvvy8ijUC1hPXVUepECEkng0MNvlcG7
wgmRhd3Cac2dkS0w/A5Br/3SqeQGiK4L52D7uucTKRdI71Gs9eWd9jUQe4sFxyRI
yWmnWg/d19cSoKtsREpFXkIqDsfPp7cCew4H4Hcw4YIyD5eZUXMde+FScdhJuKSc
89AtdRoF1xwHvUhuJDINh/vcVJayOtVq782+lTlMYFMsgIUZ9OXxnXGg2zm+AORU
/sBQSQAWkFoSEuluYV1KLo2KC3xfxAQv22eDje1MxzMy8pmkCC01WLttiNEW5hjd
P26dO+oVVdB0UXd65F2EdjDO7/1BCviN4EVT7xUeCROTb1p7bAO9Tv3AGRcHT/3P
D/P5jj6wb/RGvgna04TWYTsTuc0fDp2LyNezBVv4f6bgsGykwg9FhFslTZpYKhiA
pqBCywP6R7vNGhkr5Wam8lytCXfkBv6kbCLOmDgFd75SmkfhZeqBrl/SpO2p5TSs
VjUAms1RlXgumbtIkHd5qMenOaWC0Xr6atrL3fBaMdjenwIho0XnCOv9wnsGzbJ+
xMSWFArSiU0prJiXYMh7gI4XpBXwq/JAoGIz2HGBwD5tiP26Mn6fND42OIFb1WVU
7AmqMfpc6s8JV3tk7pRZdfI+N0GCFQG1MNfOGHtcdG5RU/j4/aV/ZkIrL5Avik4u
DDQFedsFeLOD8LrS2h3TfB7pK4U+Lz+U65trU/j/lwyPVC6RhPDK7DtCINBuQHdn
c/jGc8+olyyR5igwzBfe81/fWXYDUVNMBN4c9UuCpMgJ6EldgrcGceD+PyZURTiL
GJCvs1pTXZHhsfP4lHJ0Oy08hF2J3VbUYUo3buLov4q/TP4patLveDZNtvTrqj1l
8TknYDyIeTeC3ExE6rVMhcicPTPcgmx/4W/XRmY2ZCZLIX/TTxVJYd/8UM17pji8
HfErZmbPmvNRKukjObhtk1qHUd3kJwslXvEiHy4GgYg/YIL0H0J9qZsId+y09G+Y
JCg/3SVdkmHFs8n1zrYHBhuB8Ou6wlzz+FhKh+QwF9dfFGyNQOhuEnW2a6Wl0cvA
FYdbAr6Eo9heqlrat+MGzYJpwPGpFn9IjR4/o/mez/9ze86QjE57Mg3OPxaXrDUe
MiRbEG2zfm/KvKX85nu26queFLGN/qn7s4vkrv6sdC4CRP4oosxQkFIgUv4VJfrc
OAht5T3Z5MsLkCYicV6T4A+cCnDkesSpxQHsPsw4DL9V7SpCe+03btNjLGjNaI8v
Lj2u2m9mNf34jY9BVzGaoNYI7N3rF3ZUmSnRRuhtI8gmAAELmr4xl+2+zlaJRipL
bGRVpZ7XXcmuTrJb3HGMO14zIkpBSdM6ewRueM1+hZQa6nyaYel8QED7evoQyJd6
73tD6AnyQfyCRlK7y2Lf+w5dSH9lCGbjnZ05JaTQ1NHyt86yWjWLTEXfyqYOVDeJ
bhuchsVHEYIkflh+DXvsSNrzjwrNOsQxc3CpCg66N7MQyZFJGIEVg50qKYpSbF0A
K2i3NOvqjY/5g116wBaGjDD5Pw22gp+Kf9x6Tp60H5R7g/DjaMFvwflncjiEAN8Q
IY9YwkO78oQWgK+FijyWSZLRxpm20HU6WTqqHsQasbU7A0aOAu9rvCLjMM1lMj34
OMERQZddujRgaCnWOHxjF1xu6R4DDBRI8Mt6jAphwIxL3kvJ3VyiDuSds8VXQr7h
nB485DlKpg6ejT8S+XhHi9xWQp32aTOT8lWdF+FZu3VicJeZV4giHYyTIDrzoq8U
U4x4g2YLidSf8ODCthHe6spDpHjVvC9INcae8VVQFSbVe4cCVQZhBUvWnKPRA6KN
Huooz/0ZMMl7O/HO09FdOBeyK9WsmzUp9LEHDGQORS4kEof7Z5O4d7daKQ1UfYlQ
Hz6zIR+BHYI7XxNh1giMfB4brIDwBU+UlZuAmvktLBNqqrm7fzoIJWS6wXJpn3+M
1/Ne6RT0mm9mx75O7dfgqQOKlM9YYMUHTFw0HzR9frFsZFFuwh/Szv69N3N0GdMD
wOW33HoJPQN2P6vHqBSmZaPTs9h5SCKvW3+AKAsBCo79c1GfT7ZeIkEKKzwip+aD
B3y9+Uzol41n1zWApvbAvjSNCQdpqliE2iLOEjlSSZY5iUmQmwCDAprnBYobV27j
D8S66XrxRWF7UDx8q9CASKS0eWUoFugv0iDbaCnO6YaclvhirEpHTKlHU/WcZhrv
DYcw+Y+fP2NjrSFM3IEb08/kwG2YILgwrO10PCtLbKF3DRqk20h0GiPJ2/LFMV3c
y4HUw2Pf3XlCfPKCZITW9rbwwmwa49zYu1JajfX6Q4z3IgIVHMtTTkAkMmasIr+o
HQBJKrXmptj80LI9KaImVcr8eJU4MRllIzGBlelcq9nkKEFZrXriBR+Bp5xIB0KG
ihYadBMnFjgbeY4K+lXMIc2dq1jy8udXK50VsYwXUkyc+3chrPxKIbzP6DicK8dL
nsBJ17Vp62LZVEqXwA/UWiwnJWbLPTLwe++ZJ2VYtBdupVKKexxoektr7J6Nqm7L
zmE0IBtHycMBkn/DKIR2Q6GXpbU/lFdKuR8X+C12PN6lk1UE2L+B/A211T0ah9fg
K5ust5TbyNrZL0nOFZRwi4pvWobX4EOwxi5WYqBnStUFRIrHhEQcGJYK8XSZBj/m
GHoa7V1zGaOraSqUovZG+Pk8J4aakPh9riNHs3+SC8k84i4G21jidF6WSh2i443N
6Z6XmyKVTnLJIebTkGJLr64XJ5RW08oyQZH2smeJ5tDTq2dBrEqzsacbc4Z4U6/b
Ii0ww9OG5Bvg8fOmQ3ugKICvXWPSp1gwqeBTiyDuDoE56sZS5aq27STfmMvk2het
WSFvKakxIIOIF3VXb3w3eb1NDW56impgwXX8jZRt4gUVqrVBXaPdMW6EeVS65ff+
7G3VoKEshaIdAreSpeAQTSIkEwIwHFYbFxnrYrhv5kDPKwiXP4x+1Jr/TKh6psNY
73Wb0vZtZCkuhPYtDcfseEeGC+9dco3TYNJ6186toWMz0WqktJQBTyJJf5h8eOjV
aWyMuqZvLLB+K+DllheUMe3lUSMpg0jc0X8zwqSMCFe2P5BZED4wLEIRZTJD/yZ3
EMmElygXoRoucpGcd9ccY8rjSUwWlsMzEPhZj3esniqHRthIzMvePJX+T3CkqLTz
/rWDWYppH8SSC0grCO24V/xfQ4vQB5PNlFQ9shoOUcgk2KLv96urdaBMLxHlldzk
wztfxjtDZFQRJl+74Yf5iS7Yxg2dRbCmVCLtJ6dcarxdcRpKk3qs7m+D2qJDDVuz
kw6KkHPVWeX9oUTe6NrQKvR9RPL6IdyZUHnvdqV+OslXk2HcyMX0yQPfnztT1JnG
PswzVaIJ4xWSUWbr1iLn9pR/NKwrbW+Ms3hp4CSDpl2R7VJSEaJhiMXKV9NuwF9Q
5po/YsxeB2HjMVMSmFmTYvj+oy1nCC4t8w9xoByuvBMb39PlKsv79TZsBbT7CNnS
mSE6kCOX7U9n6Pi86UQyb8MxTfVM6rL0Sh29YNaHCTcwmcs3CH7Mrgyxlkg7143N
Xl5qWT7HQoiEKM0kPmQPv3dzZLMHM8uRv82bVWVIG9W0aJ3JGFxPa0e/cLAhzQnr
NM8JPIitqGZWZMr4vHeXWm/QkpQBdJcfoXIX6QY9NjHtOeZN/xanUBUDbzlb/VaI
S0xkMxDkQ5eXsqTc+tI6gQbXDIhjfULZfpEqty8PMC3oHw+V5BYoExXCFe/Yb1Uw
8qzgb3Vp3j+Cs5fyvzW8KbfVs+XlYVfuHs6Azmj35RxtM8bwiNGQY2NcYxLUwd+p
Oo3Qna4dcRXpvFL4I/oy9gHzaLQ3TICU5+nwU0oRqY/iBy7o7t7DFOgRYeUjNmZO
+hMr7gcaBGmCbDOy1V/rz30r9cO4A2uzc6lI/Yujdabx5zFPgZSCR5QBxWDs46Nj
U4hQDx1uthUloK+gWTv1XGkUsRUc8FgH2RY0Ri2yfNfr19xFHuBnnE8xz09H1ABU
Ldy4qR9yeEeHg8ibtlHqAKcpCpxq+JRRlYthXS2/HhQ0vNi+P3Qf2QgCxoeit/3Q
5M/8NBzzrAOXoRQGOsvAu/YenyMe4o9/TtajbUQwucqSnXeDqCCfEdheVuXoM8zf
sXlFXWozMR9Af/FSznG1V5dwx9Bo7WazUbB5LB2St2PtCQHTQHtwT7Hx8obyvqCP
T3fgjj63s0QdlB0sjG9mQ02dhybWFt3Lf0XcmPKnlnPxzX4F+x+gRRbpTruu4b/Z
N8SCD4xqBRCmmTgy2iO1mZrrqGNAgQkGxGQNjsqNlm0WQahZ4pFDck0hxOnixFuH
CnB5baZlDR1Di1/tp73jinzbTSvKTVE1DuUbynpJ6fnAWsiv9mX1Jtt2xRR65PKM
Aq308FBD5fgePuZMneezT0zP4R35bCMW+77tYwvkWWCOZ0mX0rtDkDO/MAoD8pQ7
PehCuc84hJziQ9SxMfvEoO1Qe8Wdf6fiFVGXok2IEZ2QKhwujh2DlCKPAuN8CS+W
24ijw9EORgnJlCC3nOYpame1r8xlVfz9o3pLc2goLjUfBbZDsTsx+WmUUidm5k61
PsSf3O2qMmHU//c6tkJk5r8NggENOw2yW9G0TxXflTwzAUS0f9uF5YDtfXozdiUR
FyJc89eOwTEk/8M1v3h1QcfrRM/5RGke+tiyevazeVSlX6q0X3nvvtPZjeGSsBb7
mtR6nAn0smpZANv2zcAyDRQd69wVOFxZhLXcgsSqgZ1wdhl0fXRaHKMZSakxjQiU
v1MWJzEiGAGmIXxoOIHUJXTB/RgU5hkUUE8XMyfGl2YunwAbe6/ZvOuIfWo42iir
9pxEAtzp/XBBU1l4+61XmG7KDQFRQwnr/0/Bz/Z0BKYT1cU22iwVkbWNUtbdR+4C
/cfx+fwDp4s6hfSoJNi09SKAgOrklIKzziN2tlHrGWLbzWP8zujpCDV1tIvGMCKE
C6gSR7dMnBPhNKEFm6iAQUN1r5M0xuEdcqA+WQJIU/lf/lRz/GyoVWCU1mO842F5
MKiVbWL642Pe/eoh92ue2QfE7fm27cSHC76ZeNQx26Wn01ejqoiUCFR8FhA0yPys
RAr2Tcj1lCUNV6ld2J3PH7jGwTEnK4mBDLfS4XLmq/MnIHSKUiTxssgucmIO96Ys
4vV46mVJzjdjm+1Ya66jVgRAdi446/Uxnr6hrT7jHyKKp1psGq6ebZcafByA+9rI
d5OvDlZtJ4m2AjpaNFNxz0VxHo2d6k1qfMrJUMKgACrWTYFV1cs7fYWoDsbOOHr+
r6JkFVe1E+BvqnG9JYd6kDtzBh/uZg+Z7YNOgBmgB7MtWR99cMKuLdviAbgoE2c5
9IbhKp0uSO/nX0SXSZvnSlnzafCuru1bhUbuXdbbJAen1kcu9fDz6xxJzMNkt/CV
3hcSbGTbp7w7fRkRJVr9q2ozLtalxtpT/FOkM3+eoLHFt3kMh+X1kkjZ8DhGeERC
+PjIfX5hoR4YfBT1Fp4HMoNHiMZgmBdkg1w3nbWksTHEv7L+v/al40iNGW8uwTYo
M8lG5WV6Fk9zKaoVIasz2P5503zUaLxA52RP4NHiC/JxefH+QASQGGp/M7igMQU5
fuuPQx0KX+XoGZTqvPxUvstKNCiqD8TG5BCJOsQdj9HnxI4SShrh7dyxVMwJR72F
0PtRmM7ln1UKx2arfvuw4J/grQ7hSaxLgqJo5c6Wiynqlpn74joqM24dAkFKGFaV
1ZzlA4St8Dc2zDwN0mzgOBLRxT2XJdKKPx+WNGW1ZkrDzs6vnbu7TudTadGjgxIe
fn5Z02TWH0Ka8ACXjJLSL5zcC1Ro9m3LcB2DipyTGidtSo5i6XhsN484SSF8dJa2
oH23yY6afh31LuP/a01H52xf5imXraygEYVh7oFc648gpydVvxsd/58Eq+Os0+hx
aEGfXRyYFMQHX8GDpyLsKInkL+JHGSefw/jYUx5HMBIckFWO9Gbv+eQGk6VyVjiT
q4XtkERF6X4gSK4IlA26wPR9Q5QweiCEE45AY0dYnPB/al4SU6k2Ns6+ZXzoAPuh
5pJQzzUnoIRL0ASlbP2CUHtDgZKfVD/igAkkvhgDzaFMHx6zy0qDMY4EeKwueTqp
UUOYZJhiOIIs93vbTeDdu3gK3J9amT5w8vzLw3lXCkG5l1WCnRBtH7zcjojXCCTW
17U2gcE6lwZWYIv1JYidRYiSKduQ5Spk6s+W7lw4wN46G3USabl1ATEpTr4DqgJR
f74ZHjogRBPTWip5ZlSwExys6fbr6v1ZebfINANHxrM4Xdwi5IEyc04TBscAPOg1
2XCv6lJT2W9LhJ3Y5k5SYIsMdlSDJTJ3ZZU9L+7DIkw7S9YECj1aFh2T28/t370y
OwcIBOXZkqq1rgeHPMXRs+MvveTkfyC9RM/UcBeccny9N8sAfFI6sa/MZaDGUfZV
UthFQ+yNXsr3Li7/bK7bhMyPE9HHoKWf93WRecuWClB90k6ZTHM7UgA7wr+HmSyY
ig8L+Gl7R2sJs75r5JvEUGwiY7vbCqkeVJih6pQj7vwzzWwS4eGY/lWk+77kleVI
+uT9Gj8Z2ob69T3CrrI0lKVzHsDXe0dvYDsCf07/fODpjEjXJm9Z1NMBZUeLASdt
iP6Dswr7NUZno6VZ7id4fZeu47WASnxVN46aR6IB+7WqnIkumvJm/g82/6QIt51s
cForus2vroDuU0RgK3itCvIt6fIeMS85sKcuV2DSHOazAFqRrwj3lFElvS1R14pE
ZUEHezoLXEOO2MDVqq/jkuc4o96myfToo/S0J38Wmom/yJrmNHejG4HGJxDxYicZ
C0q2xMXJ+Hs/uZtNDgK3mDv+NLqBWbrM5Jc8/tO/rxH0+OpORA8ft2ab+TXHybNz
L3+YUAsveSq4xXAviuKhA4FBOHKCyOdlzukqBJyw2/1QAFYPj6t7Di1GLDt6Om+5
Fo961gTekK/wwzufKSKvCIvkc/COX7sh3/9K8orXfqehlTgstUp9hog4etl2QX17
5omYMJtINx+ctSuwpIoW0QRpFjcCRWuo8H3/zJmE19RViI6DcS8nPYRuAcIglnxE
ZfFmVUnKU5GNGLINtLjXooHL9MBEMQu8VaWF0K4554UyKnZ2e7OkyU0H6+H16jRG
1jkTMw8hfKjJfaV1Q15olm4TVLBga/ND5uwvGpvoyt1r/gGq/qbcZfjQqShEweqw
n4oq9a++dzCjNtYOMxAxkqnJvVq13lVDz4FTJbnAWf4m48sNuZeFzxKvqtE41Ns9
NeJBIYbINLavYIvNDoQIu/g72S02N8USS4irMszn65C+n7N0otjoWUnTM16GCQf9
nG/CGNBcnNOBzieVgGevebb/ij6m174b6Nv2SKYKg/igaK7NcTiJ+1KHdLCMHFmg
IGSjv9sbhqf0KZEPfo2SyRNfuq7itITxRyCzFnQR9MSe5N8mJMUzNZnzLJ2QmASN
/hmtpKYgG57D8uJqi8e5Kh6L0i93xdUaI6nOl1F0e1ojQi7s3lRa6Cg4ryBeJ/xL
SgwrhkyZrZ+Y4NPkzxT0BP64vSP8b9Fmr3lqC1MnP2KjwqoVu/xLAWX1ILjAHVjR
MwQeId7A64sR+HVIiFKu3VxKfvuo4NliRqhx0iZ+Z4YJV9JzyZ7Rou20R2smx50P
4z4PPSj4KubF+mvCBbN4w4RBvaHTfE5RCnMJuaBAZ3dhf+pT1zjOArjKt1JXIRyp
v8n55yYfnK++mD8tnOqnzIxyd8kOIXZpAWjcIgrBCzV4hiX1LQxuIL64Bjk0gBkb
nJbdszXz0nz5OtoAAap4nGZjbmrZidv5Q3O9S9WI6dnT0rkBYWrqZ9BDAacRP5Gb
f7969pvqO0DFsLfgbHFgcjURpcJ51XlWc42L8VD1NrpTX2w/fAQ4ce0bbIhvM/aM
6XElf+UqQFPZaGNd1Jp3vxmDtz004fH2OO9PAs6+8nfFMHVzCcuuUDQVkBzXytqd
DEUn39DOOru+F59eTvZ4MKRtXJo6sTBtpiVI+2zOXvWONvvGkogKvyAEd55neY4k
3Pif+yGYmtWb+1tHKbe/ne/RgeMPHjtyMKuREB5pcjP6dqJQYl2z+EN+7FDBJSbX
1V4ubQMCMRaZlBVcXMkkGryNFA8z3UHPKBUPzqHoBLaCRWpIHoBLeUY0jjiXiIFN
UR/P7Us4rXgpln0N0X/JOQNX03s6LlHmgMeGaSNZN1kMa+j45kKfErDrq3J4EhK7
TCVWwnTfNLXPgWy4ZHprD/q5px/GKV1xI7cKHx0Vl5OIuuoxqp9esWBtEoWESy87
8OJsDB6M8U+M+1kbDP1h+aXRffOBmYmuckVt646XM1bHpQiFDM+6PQi59JVRqV+7
2hNo9VWL2VdfvX2beYlAISsnXr0ifYa2XHEF7BD4gqFF5A0DEh0aq3d7aAwOhXLw
2vtb1A5TdD8IaT0YbrsXam5B4QGcu4o6lhvnSb5ud8wi6d8c2R8cPYZGfNwos0dT
1tEDNm+73EH+Uudg2+0lbSASg3o1/R24ZiyER9Qv0AJj3LgIodj9FPZQiDOkU+z9
w4vpxs4afS1zOMDJhnLaWM7MOAYjFSB2TbqBXIr91TmFxmfk8wLnEw1fhAKRKSbo
c27Ql6LVeGxlZ49Z6GGelbdeaD4zsXu1wHNXqsM1o1Rr1Ngx6718WamkV190qUWB
z/7OWRU5wpG+mlV9iDQTmWjPQ4v7crqUQq++T5Jb4DftjjsDDTfIaLPJbS+FwmAT
uMDrMaoysw4AlenQRNSv/p50+nIgMrXG993Oj4LZwzm7a+MVPeqeoppdh9s1BFPV
DwD/EYqQveULCZY8PW2e1Q62ixKjFNATcekH0/1YEUd4A12HItGfPDy6cFsolHsw
HNjBZrVsTDM95lOpNmVKhg4cSL+l55VTY5CPBKMciWF+W/NhDNMRMn5uHCKgxY77
ivjANRKoAq+ymlalcfIMcicU2MhZe05TbhpV/Pa25dQT++cMgi5qzTAGDD4ySpcN
fRPSVdnKPpbv7MUkg2Gmma5NLmGt51OV+GgeSxXaprGs0H4BVTkKzsu8MxBAqAOo
9oiotbcMCuIw+3Ofhn47pCUBpAayRzjVY3e2HBJp6xjjs3QyILHnP29Zm6pbqK7u
YyHelxCGCw+w7iV4sjoC+xRLsuA1BHi4mcZkMDFOoyY349rP3XZsXybe18FyH6qJ
ZUELgG+lBjlCEjg5PAzBZE2+w7Vc6svb7WOfOX/EXDOIqW4k+OSlNY1OYrQPNiEe
KUKjUd3yot56mnKq2sH3f+n/vKWmGoDET4kHV6WDdZpAbh2XliIhuchJ1yJIBB44
1sIY34Tnjw2uqFA//oUoofbacqoRQVtTX4gRiWhRTXLhsdqYvxTIrVtvpLka9koX
d1EBNW1VZGz5znZx9q//ox0fwAMGkf6b8y7mqTpKJLoINc5Klaq+UlpcG47lp5dc
3rc+jFybpycGG/EfPYQSQA/BW28D3+qb+18hbPPHLocCaxFYWV2UYRz3Y2Modcmd
HltNFV4tgNDV11AfOWgwAVGumhEK2Vr5jLr0EC45fyZ8+sdCU5pWfZwk0T+UPqXl
Sf58tm/MOUcplbNpwBPD+xi5dqZ0FSohgRa/dEbOkbaQZJyw04RYOogrfGfERJRn
y3okynR0ArKCGChbZR+SrrrWgnyThIL83Wz2QTcurRRyDYfiev57kxaKiTy6zyPi
CAcEE6Xg624/SBmQabWyUo3qmkRBXGneG29ss9fxyFUIf09UeMZl3j6RG0jS7vVg
cnsSn4zpSPBoqXvz1C3QcTZeWTuycl0dKeeYVQjG7e1lrlX2L5oXjvkIJERJrnmf
T0ypsX7NcrXd3t4PPums9RsXRR+NuIary9tXiNCyf8Ih+M/Gh0HbmrhwVF3vRXtv
6PQe2c8aXyROB/cdxQbsU9FLMDwvoHdZvlqVAfDaM76B3pUTGaQUuB3UhVGpcjtG
PVaOS9yE33KOPUMt7Avuh1PVZgFUFySZvqz6Q1vOCiwf3PBP2MmJaIeB1B6jc2xt
zf2e/7hRHaxJM1LaiMkgtWZX6B/YanfUPAj5F2oKmHKZjSr8csJ2l68ndo8NJ5tu
xhr35PWnGsEF7c2AArvC6BX9XfJ4b4iJAHQJhYWRs6qySabhgh0Q+V43fOSq0v1m
cDyxwEciNnRlzQZC+/sGYGUlXjcmlBQZxajj7ksnWXS2rQsBPEzc8IVtLsIEFNhg
aT0hHSn3s+eeDolax3lJnJh8PBZBC9xLSAsxlhDTMyi1BwXXgKURv/BbsAmFAzzx
5ig36u2Ov3rAZXr9SE/zz2u1rP8i+o8lhDQkQ3hCyurpQHKoYarcQsOpbNRyTq3/
tCK/9D0rVWCpjW7d/bVtiArJKR5/TLSeWcny56rCnSFTbMU23Y4KdzEPdptasEX9
oUqTnbSqNldQ52hobJgp/eB2R2ZwfLzy3DYXUcFr0U7ykszA2RU8ujlyf2fv6pqO
0fKkxKzTqPCdAm3Mblp6yi+G15ALD7uVVWm7K8AsyOuMomUP8FBW9H4qIsze57nW
1Y8FspT4T46VBu3DDcsAOETKoH5nltkToS/27EL8thzyc44rxM0HdDufZksqt5Mk
ab3d1Mf2ddvWte6cj13XM7JdWs94nf8wUNgu5PMN7pL8iOnPXHr08yS8eTUz5Zea
tW68b6Cy/Tofyn8qC6hE/lagFSwHWUNDaAx7wiNuduZ255EbgunJqsbEPMJZc5+l
x9oiYEqSOC2tKlbGfrzRm1McI66D8g9aBdV7Gi9R3rczsNVUdn4Bq50utZHiH0qs
/CJ3AoqPbZULI+VaUP9gHmeesY/Pk8xTbYjrmymWKg4Q3RlglwHCmyi6d2jui1S/
BkHGITQoWxMkAG4LdaoHd47l1N/30zlKoRO6ViYubeGFal1ZORPzhe1iQybDLICZ
oQiXFUr8XfPPwqYL1pwhcbQm+mYZvtSqGbptMczawN2h9wt04NCcbPZqoHZg2ggq
ETJ4Edulgpo9PEhVHCxqvvMQGsuw2CKbQIwq5XtLtaiQ91l19eiXeyhT2dMuu+LY
rdEvpmYkEUZ0+lI+V9eOLG1OHhkof8fHX1vU9zhaOLop++flsrodHnldW5GQJgOw
vIzpzDbtq4zx+tPk7I12CN/C8xGBW2dAliKZErGXxcjPLumtB1OMybnMakv0dny/
BoYfRDjUDYw5bwKpQRMinu0wrTlzFOQVtTu7RoLRnvxalJNEsNUAySBFYuoqkkGY
bjiLWcks3TjagH2RCvFI/sjbJw9WWfz+s7gGY6XXjtBNkyDZ8dgWJEvehmt7MVXf
botuKEx1mBPYxxc92bhQ+FUP6WXihaHLRMeQnnrsqsTEwCGgIFQcqQhfwrqqNc5K
vmxSJImYf44ZRce+dGUZ7nA/LO8Jsvz48DrdRk9QsEKG4eCPdqjV+P5kIJuOXxh/
Acurm6u/mqEnnH2KvqT+lUqAD7Ucp6OftLYjHUKHdIvNZycdc57Upt7/xhYwfO/G
8/Mjzc1k00+NtGCWgq7tlF6wqC8lFkTQFDEWzlkgHFJtXSvd7yTGaLVRsngbGlSp
bMB18kbB7MMimBygj3iwztAkBrfW7PkvXhwFPvaRsnDvpMow2HtsCV7piAXWZiZY
LOI1PevNPm+abnnyl3VyO6UeH6p91eK8x2vg2gh2bQ+2Y1F/X2lAly0h9NEUxoyx
WPtEZDCbUoXagNqUwPTzAR4e2fRPnWM9dFqjQ+4k9neSbgDNR+JrgtUuulUiqiqO
nAFGF1FCEqYSW4yU8I24z2G4UGdULuJv1fSf8Q19QHhWxvrqfiApIF6Q4OE6y/fw
9nNKtL6klx6XGGg7ceiMwX5WDWs22CED4gItrn6iLTD8aTUfsEwzK9ns6C47yoJT
Ko/g4MLFOTKZSTcIuVzKXeg1bIDrjtzQme+41AYiASDLNOX4W6d+Bz5BF4G4vs8x
9jX1yfsc12EBqHWM1PblHUKj6u+obIFEXsKoDFdKDdhEtdDVJ38He8rkMADpPXGm
LpLiVyqh0wLKs6AGSX5XLtsq8Mi/yRft2AtcLQ5Sb9zcX21JXPtnUJQb8L1hjIiO
f0gNGLLojwxR6/AYTLWAwfC1S3PHzmoA5gFYQls/l9v14N21jSlkfjAd4Ic76bw+
tTQrBbBR524cpJwSgqA7cuNDIdD1piJaIFh4iIhX/iycpCTehBtR8Msg1yN7Sbkm
UNAsgIGq8qP8rSwJkiM4vR6Y/BmbLJM+crA1r2psDSO7x8Dpm76OC9hPA+S9Bk2q
o4zDz1p7+UiGB3hMHZ9kb1Gjc/ulnGOlRXnxya+eOZdiyjl62QlCV8eTeDk+eOrc
o/6q2JieG29NeD/hlY6GndOSuMaTcJgTZX1AvYUlntBUlcXpJjmqtTil1ezvIyja
ltllDTKTeUZgvLyV2A6ebxUHfMLOpfPMn2ZpVLv4eEXNeQ6fbbYvB36yRLjICXP1
XCPbiMi83YBGHqkJWhg2p/yhxc8gV9YwTDMcLLRtKD3H6SibA3Ak+4CUWLhuR3cd
3QkytXYsAznr6OeLWWIi9vBLu/eSObTC0oazCLEpOJfzNBTJhVyAFU98UZ2FVBGz
x20TGql7LUlYoi3F+AHH0hybClzjbB10XIvU4eUUHGS5VS9OsBskijaYPJnRPMzq
nLQ6AQLr3wW3KfP94m97gIDv8acRJpr18JBuVxmAxg7oFRYu7gO59CHNF0VyAxZs
FW0YP68lfTDbwcOIZUVeY2vmXYGnq9IrE2EypkNBqMQ0AtZvrQgofd6HLu0kHNC3
PoNsUJ0xt3BPA3yNK5WMajP21REe31C1ATdrzSf4uqZw80Lk4MZAdQKiT2NPf43y
FJb+q6mfsBoHzLWBXrQ2klk9YdY+eijvzlpWIL/8xaxe1ci9OQoYxm3fCjZcM/d8
KYek8/eLQTFB2b2hodi4Igcv3ttH1SpQ4C4oq8QXDUEc6V78yaqsZkFCxW2Bz1PQ
CN7BGdIxn/Fl55oBSgX0WfzhfHYIwKlIVhDM0TeSGiF2XPTEc4AkHW3H/3g5PGpG
8xiRN59o28vIpMyGDWAdnLRWIjbq22oBdyAf/xfT+t7S0iUZXECYI+MxVDNaEckB
sLmZ+7wZkyiTRSwT/wUq5hcxl4kqpSoV34m6LQjcLd/0miz24sfTKlxUvdhJlvNZ
hx7EkJXwjU0QeV66oI8DaQs9/NwmZMjoiRiEuUbXpH4/+xp0/U1CCwCi0Ac+DjGt
PQ66+ajxWmlz7YTVwesgRHPZO2vrE8MfppQhPRtMdGNNdnBOEqUpZRZb92h2sUAX
rJ4aRRDlQl+AaSfW6hrqeR5fT1GKO8CnFQECX8VLwrqNc1t/XAIdOvN5SwyzLRb9
ayFIRfttOKnljhP3RRNI3Ml7Ypgb88UKkeDR+BpT1+Z5cy0Dbkl1ZWDLAte69Gnu
+ENRWTU38MiJ9Pd8RUTgnapb1G4z/8EQR3AD3KNb0Xm4Y9sOubOKqHFe66pxSpFH
aVP/tHiYXzn9fT8BPCkXfGY2bFGcnEtx+oBjfRDh9gXEl3SwaYXgC/BBjRsIR1vh
3Dz6O6YPqL/2h0e9WZRAIgb5q//H9bPdOfFBBvivlWMjkKRAQ+jqEFbEoEz0GX/R
pmKeSxQkMXQ9sB92H/LG4xig7c1pP6iQ8HecUriEI5lkZq2DkNU+26lnaZ/r443S
dQEstlR3UATiEFBVVMquYeIkKk0e2COIQQcy2r56kyxEHrX3E0XwfzFwivDVz0Kt
7Ic2jPiTDs5eagn2TyBoHbBXlncwMINPSfiKdF671wfXlSCTsJHfk+w+WlL08JfN
Sc9N5voeahbGdrJ/Bqh3BmjGX4pltw82jol+2jOD14sR+i8qQnSgelCJsLjI+G62
FsFrMpupGp3oyaukPHdwrkl92ZxqAucsg+r01+VYimblQI2YHX88Ewf+ooB5Ri9r
oRpcqXRPL8HgqoKDDz3Jbg562jzs+z9A1aCVd7L6s3zNtmteFOBwL/mgRPzvIWXK
cclv8HxFd6jy30nypvnsRrhFXFFb3OFP0ekizJRzZv5/Kv4JbABbLll+7YfwH1tf
Hg0pM6Qz12iv9tXU8uf2rkMdOgYJoiBf6VCxVD8tpG3DDIOMti1MErKsJVMYr+sh
M1Ho1OPOTq05dyrxTcHmd8sjVW8CdKICzY54wbu7Y5vhbn19Uvcl/oywwhjKbOLX
8G3vc8b5mVxG3iZZPYGnkjbM5fmLTyd1+Wfn4VFpnaViaJ3egxpTxG6t3o4CFQwB
09yLyRdiAUidNWhDQdrbh4fqVLTLGC6lkunmGNDJDrsiqy8jdRUsOznciXIG8lLS
KO7ZsUxaqM4xL+cnTET39mM1Q343jeO5q8Viifub/eHSs9YGPY88HgYJi+NQZIlW
Wxcd20AdpzyQ5Di7czagApxkcjuItDRA6XI70s0P1StUMMwQSv18EEOGBnuzESQD
+1YqdAco1sB3tvn7Bair9hbZI90MgJAaiXS6ANNHLfPbHgo0/BfLVa07h9vnPrGn
u68xesnAHYoqBVra84UwEHcosVLQ04Qkv2yPSBXcMz/iAFiuYi8llbR9NAXXDENv
wWoC5PVlNeAzdr5r4/xS4ERGdDRHLNrOIuCoAY5U/INfgDbizKyj2hjpfPYgZ60A
uXxmQAEzFgWFFyRrRi6ifeaZyXxs6IV6PutFVWZL4OcOc/nd2ktCzefGZmJKWo+1
Bb41m6LP4iV15HO6dJyVpKPwoyXU2uvd2S6rF5TfKh+TopBsttCaf+4vYnRDbCSX
f/rqbbMAwWCytKXbcqz2PAt6m/s9nc7+QkMP/jIj6YbWVOq7H13bGbbZsb1WVBlG
RIPuFXHxoYCRIeeo4uEsuWI8uMDhQFhPBzVEB8+Zuk0qc8SP0rQCe589J1t8o8wz
cRRfgiQf1DvBLpqgmPD0OomRmaB16ufUA+erlZ0iQvClJhvAVuqgcrm6gjbNBJei
CGBcn4ogkQBgm2UwppGAGt2G6rNaBxmaHVI5qJ2NV4+PP6Pi9XDIfi40pf+wFwtL
AlOnbo6KusT2kqHXOsBEJOof78MEY/XNNkru+v60E8C0AqZfXNSprv53AxuCkRAo
Y2lC8hS0/Fc6xFAvWxF8mupm4zTGo+IpNEuqwPRZ4jEhONmWRrFlhvetpkQZalgl
1yApBGFLFg8aPU4gxqp0ecZFU7QZo1giAdLtHdvG6NGIlIJKDsOiEVt4fMQ8ETgn
pnWgXGI2phSZFp5pDF3FzMuUWkKxWU4+Ht68CO8xO4NXNSExPODGTG5YW1IXeg9r
0KpUMYgXTZ27gLV+trVBfatNNPWRckQUnxio9UWG9n45rzjPR4aP0jxRh2zVptrL
tzgPKgip+SfIR/4UPieyJGiI4EXRNZ3KBzZOmBTvX3FptFEM7FcNQwevJFSI9igR
Mgk9/+s0sjt2Ik+8PvJXEI3BaKL5Vyb4we24eaYZgLupSvQ6eQypotm3kfLMltb3
y4FCpxZnBqqgKQ2YTHnql3wXPV1uvvZOKhKFS312opn+n4WPeLBfPNL8NUhVcvGW
UXIsNNRv5/QW0ZSDmEBRwPj2UyjRAfjZP1E97AvltFt/Ph9URLec3vQA956mCBDc
JHWDHFdlU9W1qmBcHSdO9Ed9Zo2eI+BdzVTKYZ+CHvDfgIwuBwi3j5IcOCqDatnZ
Tj+5kLrUFb9brbgjyBR38yOv8BXB7K9jFmsXSX8qJcSTWd1uAQlXOzutmEWbDaks
x45rpS6x3XfiKzTI3LwiE88L+nSXVdL1ifj8EQ08eDtbyJtAYvMrl8Jx+FYBeJ3v
H3Ycmk7qY22mdu7T6SiSV87TreHKU0l7MoaYt6qnoWSV5dSIzs+F4MlIOs25s2e+
E/RAKxYO+F9ggBpRGSBpjE0FZ126zqmz0P4V32wO2cvfEwf216/moGPSlXMpgefe
jDZ6ebYAp6nHHkEvEsXJaUOLrbZxZs+JQzro+4kYwqmbcOYzbjyH3cvtEFImKQhZ
kkuDxUOf8+jqjkyHlBLF/oZb5g+ZJhYA62YHvw4x4Boz1RYZ9qnEZvAxe811HTI7
VxmsMfcaC0ig6mN6D4uoIB2ZL5VpsfNxdMYqk4KSHMniWD6bd/xhp98kZxSqihn4
/gKIvVN6JLdoKxpIJ8bjM1W/DCiEbPWxrdB9rToE3gPc3qz3EQAX7THm4BLpKz/5
Pmi3+aVMvShVvtatkdgccOSfw0BKn5ewX6sOfulr1vE41do7ivFgviOvHk+R4ka8
ai0CmIjsznnOaV8g7SRURWl4+cY85Vuu38jiHrj/2qeZAhvhJ16/iCOOS4WY9NyT
/B+SnUtRsSeQl4CcxdHIo2CAeDIjayawsyEB3bmYtZ5p9SB9ZL/+TOw1RruKqPol
XVk64RbXWdXg8ZqVO4Dgo/4LNboa51Eyb5qzHPcV7a0zSNPhz1dRCKsjdpU3tOSN
aAm1BPzz5yxZUwxgRbVYI6MG6DpPDVyoqY6CFLCOjV+ER9th0d/rIfGZ5T2DGpUS
/Eor2Kd+bfNJUVkJ/AIZwC8Ct6knbNH83t1I5Jl1t/JDFHexPtSiUZQDdQWqnppC
T0sa43CnJXyGAbeGE9ZEyNao044nePCJrk00YE2Q6IhSGFk54DoMJHFRwMvc9HLI
rIqBuhY2qkQeMTiMPJ7BKyCVm4m65MaZC3uihMYpx3xEtgcL/v/8At02snGPCTwM
i39iEGsow2xYymF9HB/pSW46DvvpTtB4lyr79CD6570ezjjdyNVuDHIPqKjuMGJF
CmujeDMULKYUPnX4cGvSuGHnJhejNi+TA1fXv+AFf8i4dGUtagaYp/vj563Hx23/
+EcPM8LspA3nUwm2cLDdex7YthCJAT3RSyYCC29jL588PnxuzIisA+siE5/s3gu/
k1pJtYTE/W7aorJKIKwcR5hFBhsfi+26QuJ/AnWaRJe+sP4nDGGBMGtkLA+osjBu
wFinhMNAaIfiL78anWqUn4suppY6DmTpmBS1Ocw5lkylkRBW6iCBHuMYhcGDtk8l
GVOnSjqbuSB1LptsHKWS6SKItGMCa6Dm9a03/cVmHKZa7quNLK4V6LoHtJ2dO9LR
TRF8ct+oS5gGcU6Qr/vYYyYK12XjAmsoBz0rFY+eUsHYe/X6+k1KkwvMZyWMtj7I
Xo7pC8SAcFLA+kbGVj7Xgspm3YJVj96mBiUM3sqW+Rxwivz+BXJwvqU4WKbpFYdY
neFPvvoWxgBwSmXVlQc+8jFf8/SlPqtAe/8lqnIA8ufex4XkxlSjFEzljp56n2BY
X/M/cr0t1t7G0cpwWC5aAl/Gluj5QttAB+G6HFzXNFewD3t6IqSqPcgjrJyqxPvk
xgVfvFfdI5tvRqDmVpjxWQr7Joz7e8mvSIxT+pSLftMRvsU9pBQCLfTLFjKVniP+
wMzKFe3KNuhKb1GEq9dIk3f8vny/PY4sekbslhpJ6tQ1rqx4I+OcbQ77jCPuIrqI
bB4xrsa6YMLVLxApMUmM33xUXJZkNEt8P6Lhtd0Js8RWybnWzwGYG47QsUHX3FHE
/yN2wZcBIhRzpv9RWqnrliUzkAMP8e3c1xFp6BX+8aqFg4kPlCbsDy7EFa4/8nJc
8iuW1gsyBJmBXhZ7NnjBi4N3ZriFGpbALITt7d0hux57Cn5Da/i53LnehNqNgOQf
pxyetMOIHH5sX4MhHg8dZwWv8ujD6dxEXU9JuvX8S06fRZe/5lB5MANT6qqI96t5
mHregIBhXICqO6Xj3zwd1UYKA5ibbau+5Svmyp5J6iM6mh7qTYsVVYivxN6Fq9nM
T9jevPWHVw7btsJqpGlr47uTNl6VNg+MKleSsnVkTu/6gyN1pczkQ3JPNRqWINjX
CYT0s6/DS95Q/JVQgR66Kkl4A0uXh0NM7dn5cHvkH/kgqpDHrJ/5uZW/hCIUZxmz
f5+Yv4GbZWbq1MQ39WBusoLRIyzFN4bzc3D83IM6ySsg5CmR4PwF+l2AIA10GS3P
ZUQDNj0H3TM4cCADNvYsHJ8Txa1DShOgQzNxf9zCTaooyuikkjp/pBDJPLnfzEWz
MuimPYhsqriHK0ik+wlPUkGjjlJw1oNxuTFFvFFeH3mC9n9WuB7VfMM1LdfzoHVg
0NHJRYf5piPANzRFP3Vt/DEFxIO61b1zbxWNFFuIapqsw5G1U8feshjCbu5R5ZuP
T3UUwMnqq5J59lBoGJg+90jmd8qtjOYDGFkArYf1VnarVwYoPM5DO24v2e9FyPKb
fOXC8AGMgH3HVnyX+mcQe6ca728L0mFkb2VCWp9YORNxOX4vz45o5fQlbRGq1y3V
95ZaH7mwxRAnHCbj/DBcs8tOw0XWR5AYLWnh/VCIkN5g0kMih+ULJkGEkky5uXXO
6s6/MG8WjWMk8/X5d4e/DO7Bwwh2xSrkkLlM4dHDJ4u9zC6ZOSvVsbLVJ42RtbTp
QqyJ41l+nE0Eaw5UVC6unCmkVFeiiMp96spXZc82FCFgKVF04iqq9POdByv2ndJV
hix1hdXLOUrmx3Y336yDnnzt8X+qWkrWCL1hVeMPL8UVp/oNbbp6bECaUCceZVzu
3dvf9Is+jZD6Cs3hLuk0JbKYigNjK9Ni0Xq6skD1lYVsEc2YizoVpuP9/jxYrynb
3l9tyJSX/uQCCRytcFbaHzxeDkKzJplhLZGC3PLnx0RlisGqFRwuXKz/i1p7y/uu
2WgHxiGm/jDQo5MCDqbztIZF9cyMXHHPJMaJ8vKVrI3WPYlPJ6wAln72eiz0JVAo
i/zM0QdUhl9JQutuNWqJ1FO1HBGTRJToVqwf1X6ILkZIjc9+TZH3Y2UCrOI/N2HS
Grt/UPTfUqNvpmcMNzPGygx5z1iLUT0SwHjaf4kWyHxYL9V8FhdNhfSE47mSeIry
GK4509k31de9yrJaxFGXU1SL7F7qruqjRTRgIhf4/mGJ1z5YFiTCwmVLd+Z2nGjs
d/HEQlKlORhNo/18P/RWrEoqKa6INv8TieGs9uFh2yb9OhowPHEzrsogMANo44ZL
R2DuKbJLR49aYS6t50KB3gNMdXwtd2HrvwCWWDhGn5yu5LxwXCYwbn1fItZN2Sc6
WQKXhJBuHzHG3y8xvs/iLLt+kv5oDXnNMIapIblnMF4C/82VBJ6EdNQHkY+fgd7K
a8VNML+8o1cjqYox+6kfHXvfESVPHfyzxXVCyV3qoydrT8Uaj7mn76xU5VMSSxg6
1oiU5VOAl2QgCfv8ffjGNHKjqD4uNfWOhdZCoWp3gjGC36BUKEHDSit5zzl4sCg/
Ebd/e+bx0t4NVFKV4NgNgR7+Q/yWF7Q5GnXT3aV/pO8Nc2EzOSmkJhEtEbvtPV7H
xRsDPp6sAb2FqLL6ykhwYLkmQ1c/VNHI7A7MiIpNvfc9YstqQjPjsS0nJHzSNvKh
k9IoCEfK4zOa83wKUeZkUQwH0OwT8JsWFzCzf6HppfMp6yqWV7SOZaINsfGKVxXu
PIbMCnQOKii1dxKBNCagiowuZxcTyl+AzGfB2lJso5pbSgaYh9R5QpXOp8Hl7DVS
yUOxqMw/41Btb2lrNz8BBrXn9cFBB7i1I+9DLbtvaaGW9Ned2qZ7CBTWdV2oj38I
1+Nzz/qO8HIdy0B3mA8ZI0CEY08CQOxBuXjcXHsQhf4FQYgyK71Eghb9b8KSXfR5
iUf8iwrOPdIWFn7O2YrAqsUPyyQzlz4U7TXzDQSbzJesxYQgoV7HRT5x1l7E9jyK
/SypzMiXBYcv86i7zNQMZVXeLroXJiV/2T0hAohe8zfsjXRJQIwass6tl/n36H0b
ZaVM6wxb8NfHE+zsVMzVpF8iat6WDkTRWtvW5Qlw74JZkvydOtEuwMjex+5RsFIY
k1H48UCElyOooxMIYqh/qrf6jOsg9FaKW0SJEfVvVO/tW8G22VVoSaz+y/OZ+2vX
dX2BQob2zh/CEBPQr8BgJPBNYpgj/nZOdtRToLpCha6YsfH8LHJctrqPJTtX1K0N
RPO+ovY+pVgY+AHyciusUiBRUN5cqjp7+KCERxP2Fea8TiM+R59Z+80paTOt8P4h
PsF/WlGhBaPSNXu9Zp8/uywKkBKY3+T26NhHkhfb8I3K02ycIFZEORhY3ku24bX2
SleTRMQh7vVir6mFTquyESGsKUoOshfQCE0WjVy3iaJ8d/KtwmxCUgwksq/qN7fx
YbY+KhIb2TsLHmzAjVBGpqVWIyNO5l5yLkO9zBjB0tl1b5W/YsGx4gK+jQEJMcC7
tp677HpA20F68B1WMLwv8JAUa6q0lU+fX0jF3d63W/WlE1bbTrjcjfEwH3NrxG1A
HlPhQuLSirvG+MtAtuH6bE1gVIEybKj301GsPYUWbLAveQFnZ9oDguSYQ3Pdb7Uo
+2PT9Vc3veqqOWrr6LKcIOI1Gs3l2/RCbXq60A9I+vPOc+Mo/ws5mcekrjCZc3n3
jaHyMtBOwml6wTm3HOuohoUjZALF8oKDd2KgjZK7vM89DvzYXz2vrD5qR1YG+IZs
bJPBWmEm4+w9A/6d27UcH1cFyp2PNYmWYVv11Rdw32GdlW0zqD3vbR7mTF5hZ+re
at87D5xyo0C31aAJd+O2v31Kgo7unU+pwGzYjFKoXEpn+tiZtnMje2eueUmXZdbv
Z/nq33/u9JUDCZXBktAcBYsG7QpDruDHJJxsVH8OF0HlRreKWkipfqobSTaCiw6B
vz0UIG7cxZVu/YD98as3jYFj4+inyMT1AO/QcGaSs2nqViRZFTjPXrX0G0YRRGKr
BuOIoOxyH8mhf94CVf3fEFtKNbBSsBEyPGpoRlMsUGiCZbdfgVa5QVP6NOVLx6lG
LBlvxn998TkNbHObMtMlbo6TZPJ8L0P9Kns392vU4bWnFSjxyw74DdO7HtdMRUAx
+VFhp7D6rmXsh8371r0Y9XavCud5m/BMRCAb5iSU+UMidao+csp0n4EsWDgcPf3g
5Qvu38ApteBfdoQlh42+SRbR2AXdSEZWxpAGOuNwEudQGa358t2uzfCgufMJ4VZz
gsV+AYDE2WvAt26l4w1dRUQvmHnSpu345daD1xoIrTkZs7J4qWrhuUgm6bw2TLmL
T/1mEKW5nJjc3YXkq2b2cF4AFcCEbBapcqalUghmchfJOm0pCM6Ymj7p+K3RMDNe
R+lG4cp9QHEm61LPbBaWTnKeqVeGnCRoeHQV4yHGAP0cIdLgbJNYwRuk6G7EAXBY
VwtP+OFZ9T5o+8kOOOokt8qZvlqbd0heSaAqKt/M9F+fWh5MlMZ1dZqfuFXvFY5f
izib6Uf8wfcnF24rlH1nJVv0S0doubz4MtEGXNN+d6mXe/flgMVxCTnXnX+6VN1c
4DcqXu5/d4NKAYr0LyVyR3rJtvvyZJ3SQApzujqCgHrAti20aSXCL1FB19nfXLWg
BAa8MWxlxpcSELkqdwjBptYZnYXNUXY+upqHDbqT/bIZUNjpYUAyPkd+g6TF3Uhj
fZNg1bfxw++J6MrwECSrmMMib1Utm9c+3mtFtVn7DozQOzZ1FVplcg7q+ddw8LpE
jSPtqSZ1gjW5IEb0P5+JAcnUDC66RpPYfepInSoCA0wcFr8MPtmNWJw5KX3AYRPz
CZ/6VBBJ0+Yi8ekNNHkWWqW3F/Wlid9o9HM2xyXEXQL54g6lwpIi4r01pO9DtKDz
qhh72z/NtFJk3hQO0qBtpLmBpVdO8Kv3B5PHrbeG6SBKnE95rrWXZ4MrSsG//QdE
9EK45tNjOGUYckIbBSFE/Ip6GyJgOvZ5squ0dkXyvq6zC+U7I10Iqiu/VGcgWAKj
altHmX021Uu5a2sSwusa7oe2ljlkzeh8KSYaaHqxPefnPOAbPRsIF6sclwQ2J3JK
QfNXMcC05LJsd2OW0nJ6QiwzHbyzC2E4TwJPsHVSzkirOX2FtNmcpopxe76D8fbX
LzoI4YN1mq5lYYln5GoC3eJTxfmAJFMjuK/GB5ychXKgjR32IANOcX2T+F+A4bhA
3ym9Y5NSKdT5EUgNsa4fBOvtq1jYfGjfzjY2hYZImMSF0hSaHZHpFqvZwb9GBYtg
i+Zph6wWN5Hudrdkpt89x/6D9auFXEeWNj50r0ZncupcwZwncnXHgbaxNFmFhsTy
faIcNKQkT3h5DZYlW/SlYyVCNokcNoiyzhzwoq3y0KsbR1F+MnF7cBUV7NyWFCNe
lNSTMH5sV7EZHhBzp0fV48QC5LW42J/qZjVlVQ6TVScLYxmc1aqexmvkXEXl/KUe
/Uh8NnQoDI0GPq9liqkfdnq7ELuvSdaDyMSnZvyaSf041bQuyj5yOtOK/ZBZpiJs
rNCsha5M/mZ2lrcym6EyHUMOyt8sBly4Tjyf1KYf4Dj6xwV/JNe6xWAqxV2W/4k9
qcH+yNP2axpgjNsU1CHvxj3UusOEHT3bvyfJr6rMLT553XDWH4OgY1SdGlNpnsNc
nzqMIsQNLthqMiimzV/akMX6NzItN/jTa2TH5/yvWh9XKAYuuDKGuyxsvAlLlS9o
xeUff77V0ppzir8B08zXqOYQUr6IA7dqJHIa51YUqT00+vF6goJ8nJ8uwtqKSrj6
2op0UrlwOYIokAE9NadshECvwgLuTnJ5Hmc8dS6V5kHE70pZjbx1VGdjUO4Avh43
bQPupTaO0r6SrsQeziESPThbcPBr8coTbrqxUmlT2H+utSYcMgJ6oM7wUxzldaFe
UHTiJnXQrRn8pSNcmJMMy6sxmC62DNNlSkcxqvtd4MMu8kSgggSCRkJ3wYRjnCuf
MOhRCoVeISbuaysvai/OX6C/yhr8UlmdpcnhEop4cHqutuppuOzGWIIAn79z9qUG
c8jlTxFs+UZkQEvNiyoPdTz/o0aKvgHOhR4v8j27Co9hpeoWqlqvmvrl2276UAtd
6GUnN+DTsEI1s/oqRuxgGCC2my0Ir4i/JQPr7izexKq1wWOEKbLsuIMzlALN2N7C
/RJ+FNdt4rHf6o+EO3xp+yn/wYDtpg1oMyElkqvXMLUCTuCncpyR5J6WV3pyvfC5
dFaaPNQpyY+Z3W3pPHBD1EH64Hzrlng7d6OHCxOc0OTlx5JDCU+aH7GdIcRcUFpF
2LIwmLAKNqZOrMiCn5GMQ4YtYnFwpXXWMwAsYNw46JUr1RV8OvBFouhCK48580q8
+puHQWneojaAAOcRvhGewT2RXDgP+izOk/Fc+2uj0vL2IJGWSkaDQ+iGhpHEmfxs
NNQFoldjF7Iy9Fo4HqUyQbtu/g5esOvIAVvO0NGxQHv4X46Z3K1yWXSc4gvYtiPs
jjvxc6UmvVC9pYbBxigSwx7qr2/ZeYTv7ItwpniSLF8wOYBN6ufFWcYzBpVL6vpn
yaB0xo09yce2AvtBAXA1KfSgzNOMgUvV50LnMg8Bmu0ryZhitCC9P6yFLJxuBs+2
dNh7+gAgOXC8smr759IH2AEEcN+vudcwlKziVvgCPWqx4jAqyfZ6E6beTkeae/Kz
URnciwI1qT7mhBtsFqIpzUCq5n4lhealBaOI39w7V1rmlJAVKo0YQoqHTJSEfkRM
ybvOAT+PMxzZQPivlj6TF8CGcUE9zYUWfZfccXdDOUO2FuHNAtS/YtdZpWlzfFHo
QfJUeo/rIcB5E6RrKgr8j1XZ7O+RjqafYy0QNqIY8m/Aoxk34CxuunTxxyTb3eGg
ea54yVZP8b9Ha58ucufQHXgTCqE7XXWAD4C2dvST/HVTAO9aAjT9nUw/h0hSVrnE
8g3ZflAM/5trMuD/l7IM19wkdZm+CWkzM9PXrG2lROq0VWQj+lfwg/wullHuFXfk
qsnJ/F+P9WGpduUyORhAZC5OXTcma1VIoly5cDhCl014KXqsT30KyeRVumISTF/E
povzziAaLvpuFk6xloF+7cUN6MtbJpl3G7hSnW1ZjaIvGnE6L8z+M50gkcUEOzvI
ZcLb4JiAX5QPKbtH/jsvtlR8FXX34h8uDPxUbhy7aCtoP1YCrfaqRD8O07+/2Jfk
jTx9g2XMtTbrEmFew4XKpinSnSMhNWES9b954H5dHMsT+2B/BcQR9yElzgMSwbDW
1CoSKPYLKQvJbuozmS9Kaw5VYxrgYD6DfRC+BXbzlEm+j24QKuPC61YEqil//2Ih
wyGyOy7kjVw4A782jNKTnObNYoNojqpd26DtazTlwUHU0ydGHa66loR/LS17dNps
AttVBRET6GyRK8zAOl8AfEmHnY8HZ4cnV4zAzJqghYXRqTACzdJLGTiGVRnyeaxS
yE0BwMyZrqMNXwmcDvo5pRX1C3UaEhs5lJrlzZK4ZnjDaBNRYGA82T+wHLMJHcUr
oICRaDJGaIpudQMG7NYiQcaFobreoN6wgefOqjJhx+H3aBWfh00d82L0nJLr0aoz
gJub/osIU1EVAnlob28/eoV+4VZHRkwWuV6OWTz+Q0fXA2V3Ug6u4xE+F7ph4k+7
Q1XqGnx57O6HkE/wfkkd4Ofw/4RjBIq6wB5v7bKVIktaBVdrq2gfnKrzO+M2Jsov
bWbBpN5ZVusqpYeACbE5OGmqrB/l525tYBTiQkjmsnlffjhKgmSWAEgtsSwjtS8r
E/MuWPHdXv0QDAqaTyIOJKpOBKRYj/HtcFRbqoNZB1l4AetBTUNP0mWaups9eYCh
4tnp66rg4gl2qNqHhxZKWUBLjjyJEyzl0OocqFhSNj+W/g9eZhElqy0/DcvBfPqG
IWvKkZWNDQHFMLD6/WgQeT4ia+zMJgf97f1U+x5cnt+QmU0UqoM8TOCh9zExou5j
SPOJwvU7cOJsMCZVLTVyn3cXT9DNBxFLqccQ/RvvdgNo8i753/9kw2Vc40Q0ZzCg
/QvrQ53gFf7etCcZM6VUzLjcJ5TeYeStTPfP6stWUIrIgRRKBB9GmjD3twxk7Nyk
o5pm57xfBiKqhdfYhtfJ1v0DWtu1BJRaSSBywvSxV3ldB3M9pB1TrOCk6/CCNmIs
fVs35BFO31bmpzdi7vDdfi11Zzkyuppnf8EoQ2B6k4TxKBdk2KFMbTpIiH2zAeqX
vbdAkTsCdYECNfed5xcajLE8DAiZ+d4zbGrUVkbbouZgfDK8YZ/KbX/fuatf6U2V
5Kt9r9EqvgDcbI/hyZpX+Ji7UsRlYHSxlYfn+c5vXP3TVxe85a48h18CumheCtgm
5BvvNqRu8qmVb4e2pfFVn1/sJjMwa+QQ/QB/4zbjxRLT2UkyowBXK/C7IZaMsatf
ANbr17OVLg7CGFaJ2NBVgvLGiUsjvrFXPr9fSSAolW/HWyEOiQAym2A0GOrXctqg
Yg5SH6MsFtpf7AP55dzM1w8eFp4gAQqvHlvoCGasezFV9H9FoKMNaeKlb0DVhnOP
ynAcGhhZbcu9UUCjCKRKBmyhEXMaofhqripTr641BenWXaLlczIUqmavF9ncqQPa
iBiYjKnlIK/R0X84X9gNQ3olmYKenCki2/3jvy8kw88F8js9WtmiaKalx0A7ykxe
IVSdUCrhh/nPMMY9wZEtDxOpvGiJuz2cQX5Qhyn1t9lwnP3ek2hL1/2G5fcSLAG4
Bwm6xg/D2atNsxoHfL7wGhStJaoXmgqAle2nFmPcPq5FgWOkw9+lXbIoI5jml9ye
7s1dW/tHszHUU3FUybK1lAblBeEYqHvSJLpNn8zU2zSC+tYVBdPQYgkME7tyOQ7H
ZlLE9/aXFjVFYLjSkRyvmTfMWsxELOO9av/KtjeBAPwrXCRNinVDWEWj2Vh8sIWf
gi2u8Ne5ckiot2KWnPA0YJcjf1Iw+UrnKH6pqz12KS4Z9fDEjZiKzwrIkTGkefvB
5+AYQUDK8wuTUV5OcUkXdB7HZrvzhwf5Rfn4GPXtfQhRL5WZJ7CL5LH78gK1+nSx
m+/TdDLCa+Ta3GzWH9yCYM1QrgIzvAG4bNbfwjV6bPaemDfcg23ItTqkUFcp/ySw
8diYoW3aZqi2iGO6X2fwQMYC1WY6UoQCtFcTh5MSlbudy3eSjA5Aqc9s2uzxU17g
6Gha+bk9XAx3ejxL4dEjseWhruhzBoFC7obrn+Zn/fH7KTzuHBSR8MsQZTHSupZm
YI2q0K1IMba5sU/lL8JsfI083tnvSnfINrZE6zaX5WcmVEqTVg373OK8IztNqAwp
LZLEkX9iVWPzTKnp5b1eH9WrKFZXIE4KbcLkOjsGGZDB1wvNoIDOopM5JDf9uY91
vwtQyosyvuvHDVic7LqVb5AbQskkYerO1CbN1q8hdwCYIi34l/UJYWlvxJvJAFiM
/lm/PjqEpnGv2is+8i7EyAPEM//+vvo/D0my6bf82lxFMxckjZy6Pp7ZhXR8ytWT
w1ScwKhzfkwgwQzFG1H479DKfjqxEcmNgWuO2mB2bHQDdug+TalmsMF23146m4fD
H0bv9/dACZ6zr5vORm0FgtPGoP48SCDkFDBr4+33yhEBp9ID2ZUm21lQqXju4m8p
g9TNS84LbjzsGEWFlMyPZ35LneV2NARoh58QUy8a/Vj4dPL32KjFcz+JxdUaG3pb
D4Rfxo2xoqYLUvHauIDMPUfHKcp7VFgzlW57xSWhKGGGB0BCRqidSOGQQK5zour4
uXldPANNOM5wl8NNBLeZ/emChsnfke8R+aAJgscVXr/KDZh6K6i4xte0M20SrFy8
WX7KUuUASvA0MBEnl/MUDjXlRiAbXk9WKS2lhHUqtgQilUFJW82BiVXc0UJNr+y2
OZoGqIdlZ/ozVM/yEmFFY4yYnjt6uoPODCZ4cgBYuZ4+hIl/eRjDsyfj/PhZ1X8c
ZEMgiDaer7+Q+0nkP+5iVXiL9W7OB9Q8WEw9HQccssZVsW35xmOnGtxiRZwxRAYv
ZXtHaQBo0FRINejm9+d9fbmK4B7EcNHR8yQHWvXLhWLy5LK3fb95wCsZGoX+YO5k
pbaORQsXv0DtoAnLbrFsMkiaU5FkbejC7UTfAl1PudlbCp5NW2XL6yrx9sUVEp7t
90qe4F7sTHzCxIAP7gcxDMXOz9RxEaeG4W3Xgm94JofNkRhEFzNZZArSZpAvb9x2
IJ8kJkQ/wngmU/eHXQCXF+kxMY/V+D9r2h57Z7P9YOODdylFap1J++Wvf+YM2YDx
AtvlG80W2Zpm0ts3PCkQEsxdjG4gmDpbgR49zAfQK2C9qBWAso/OezY14AqWKsrx
guwGO30UCXDhAAbRzCo/3LRZZpZjPYur9FqCqlcGQpEyQMdUh/10/gBS1Tlwhwi2
478GsY7sdB8okhXCTCXlPuOiUrKjlvfaFYQXGzkNENY2WdiWB6GIoi4lR62IzBqV
B0kaqdPtG86YXJIdQQOqVAxDWeqWR9YEUNm0qQKtUI3xgg+VeiJtX8nWd7ey15lb
vRqO91/VLtY3rkPyxp1ykPDxfeyUFLb1ZmfGXthMKyfNCyjItvRRRQYdNVRmKe1C
EM0eh7UpIYNDJSOnXUNCpmWCO/uZ9LMXbhtCslUyAgqPEazjFek2uILb2az1idAf
sh3JDzBEa3c8ItfAMaLaVkf7np+P+mtG3ZY8SC7dfsOwBOzKFt+unu6jCDQApgLA
udEOq6BzPAVHiiaE9av6Ahv5JEJCfk/woRkNOuZjsezW+HApQX7XefMVMCA1NIXv
yx0FHJppiPNdGRKq0K0eMvbqeOSOsTioGLMrN1Q8PZkvcYN/aRNN0aJISPdEMvfJ
yf6ZXX8Xn9wCWwMl1bDnXvmwAb2MOE0EFzaPJG+Gs0Sj9VZdazODzO4gMtDVJkyt
yWgo1Qld2hJ7Rm5sGUy/RKRiL7UgBD6mKG8HyYTUiCUvKtAI4b70vOZKSWnL4xX+
S9fp6CWJ7MjPMkJaGuBfSAz1FeaeorQZqOj0Lg53+nQ+HFKr7xAK2YBlKok+Sf61
0j3L+5+gCIyQIYXATY+zpUAMmdXS9q4zbUM2NimnNRzGsT7p+lypJyayfe7XZ27F
GlgxAw9JqlLP34im/v0AyRdefH8FExDO91UadJ36t8H1m9kRxxOwDeJnk56n0KS3
9KOFuuB8nVmkkGwYu6YqnHqzbfhJZW0NX3wUzI79TNZnbXjD6jmUIBPxjfLBy25Z
IzDcwLvX6qyPzROkoLMH8Yqrwe6Oz4vXuQvG5esvCDgrtOWH++JFoC3ZEG1gS0fz
dZDqNMgshlLjDGSW1j6I21PQuvn4LrqP3yGcO4uheozhj911QSXSS+F70Wckrz9S
Y5sy+4/L715bTHKIfQtSV6VqMEILG0b6rJ5MGbJr2hIafgh6LwQ+8trRR3FOr/Fr
x6ySih2l17YvI83UgHYxj0uYkZ3NyKAXU/N/khjg2JwoSPz5r4G9HXd1XmWuBSzR
o+l5ekzfYcQwggE5tsujmshPUWR5LpTR6+5RxuvgZCdjYDGwzl+pmpA0rQsDV3sC
dwUCKYAdUmMyQXJzICng1pyJm9JUR9Ixtn3lgJ5vsnzQNsbTMMA7BzdMYG+suVif
lhZ52UkcTLd7hEnIpBvSC7rJ6rlS5iw0TUI13hCJ6BSw+L2u7PlBuCT/ZmK3zKYM
uldLFj0xiFYij7090wIGfPPkyYsC+6L16uX1jEaKokE+j+yI9OgkYWDOOyXpe9p1
eAiwObo3/5HTc1vIZQnQKnM4vgDcQzPDkjKZ9SOcMRvzR8ZEuYA4mA83WRuQZjFs
aQ7h5WFcZh467OgORHrnWw2/PAcoKK1alsYrwLHXj5iTAfhlhRCl3rh29IHGCttb
NZu8t8YTpU7cUvT8JR1f9c3bwiPn8AqOTTDz3F+pHGqS9yBcjPa+x5EMvxbzGbNN
22OYC8JSTDMhN1jaEd10oc44/eCM5i5eau4EUJCwPmym2n/eGlrMf9ygOeeYeJcA
Uz3M4mRYQESxJdsHyPNsdGQNdGboFmLoXqgPnMdq7ADzAG58qJr8LYwwJJrns95I
Bo/B/qT3mWVZPIFoDfXzMI3GqQa40sHh3buVFkp/Ly2fsCyhRsd0oo1at9pAHiIo
ZozH1RP/HYQd48WDDHY2UTnuPXjUclxcgxdeF/d5Txv3c8RlyFJuy7DL6ihV2tqJ
alLdXPCMnw/GlxlgPrgn5NEkszPrtmwQRylMeJwwlxx6GktL6Kbid1JXG2whqZdY
AOjttWmjrLegZ/b7ZvB7xtaH9oGp85CwQtkR9SOOUTytly4J2W1yU68iosfTwEFr
QlLwpSheRsDHA8W8D67y6Zm10VYQsyxQ0pSJRb3pYJNOQ6noUN5zaFdClGmORvU9
QbH2Thhj81PedeKa7+2xU/RVZAJTv3RQfoLh6QrTCAD7tc9QrhOQ8Qopd0bM2tRx
FFGrX9bZ563pPzspGxUlCJrwmT36FJ0whpE9XmIG1KvG1WQb3vDbG6IK79fZRsLL
tDwy4hUpZxb4E1V5q4a7LaPTfogOg5if9iiBd/ybvtb81GhtVvSChswTtxtz/Ape
2q9THOVxBrHFWLe60KdC2gDdxc7cnH0v+X/0g+dOP+J/utfPch5QXSXv/G16Xap1
SuyLcypOWAnxwax5Du1gRNcOQvV8XMSEgc9bjr2NC1VNAx5B2LANrr1M2Bpwp4Pw
1qw9KIRwk4/f4+fh1ru0v8NWSGw6fMaFl+/TwTZ6DipWkF6akP1SWjBSYFhUGAfm
UtbGhJ/M+6Kmc1EuNuQjd0SypXQ3tIscrqEtcjFxn0BdL4LTYC94KbU36nQG7Z1S
Wsr8OeEhejeJhnbvJOKZLE69lNIQo+shqSbPMk3Ttryu9TfyS2UdeOGN5RNCKLYw
22PKqtgjfdkLVkAlw9av/Br6YwR40KOV+fhOvHnueJBiRQ40sXVGVcTTnDK9SmEH
6UNsUC7rFtBWIjOa7bbSMc38rQ5szTeYic79WW6GgMLZ6M3JkFbJ0BsMdppU7QDM
EnnUUMmqTWZIIdLCO/ltSpS/xpIhG6xq1MC2dU2LpSBkqftPHTrpAeLeB7Eg3c90
tPTb4fJYDudDD1r4h+6JVWW1EdwBUnzvF58z1SR+o1J7ld3h7GJR0L+eqx0axSKl
GELwX5cfxPTSQdqQg6h25qvW0CwWeVBFeIFJjogeAS/Zpz0U0vuZtciYc+MXCseJ
RP55egvBLjlvP/CUm2j8qAP4EaFrXgeNGqhguIX7bUzQBy/lJyMxTDJFObSyOFbJ
tHmbUQcjA+H3BKkRnkS/91PclfWlUvHHMOATpEzJlponJnShjh4GQiGViPU2+FZ6
PpnGXswFx/Gz+jgB5QM7Ofl5+P4z2E7U/TMQcmBaFct/hYYpYF3R3qlnSY5nmVtA
N//wACMsYqqwjwJGrXEnY2MX1zI2TqEDGqr5qyIVz3+3HL5g+hvidaSjH2j4znRB
l6K5ivfsZoIr2KlkZw8O93rC+lGYijRv0m+qPXjyYWFAQNzL2UHZOQVIYzBCbUGO
DfZJKyVYZ9PXE5vrc17WJiLuJxFJvWIIo4sjRPuaQxfNbVayx1L+GttvUJrwBQJz
rNqZlk0A80QqIZ0kwcYjTksoKjNCX0l/YQc3rDE83+DNK2OYYgmRVyq2oPdVeDHj
wXykCd6lWazK6duPKbvTgVeb9nMl5xnhw+lniEE29g2KQnW4FDM8eSIknHHhP9O+
U28mdjru1TejzHx30anZAxNoQNZtRqbNjvChgzmcxCGJmZ1ouKjHVjFJPIKpAaVV
O5LYA6LKMsszMl7hI9rAkcC0xy+zkbnzd2+IFLcAJO5R8TKMDW6eCjUI9//4J/KZ
Z9nUtCJC7uIBImSrmmyI4Lueb7V8+mapfugwmRouEGECiM7tIY35yWtpnScYJ4/6
ec4oLkyu+iazAAmIEQI18L0TBO6wq0B8M6FoTbXqZsY2SghDOdwD9Be6TU0Cbvyq
vA3b8L/NUkedZ+U4cw7tZ0orsYaOaqMkumdnK1iPrL140+5LWRAxL4sPtmLmHKPC
NmeWEuSnTLJzET8uVTzAID7/axp3Uk+C3wWx+tkt4US79RMrT2iuxNImpiF+1k6X
3iaYNDsugPuBeFHAedrQbfqRpEif9eu59AehIOqmYYAky1BAasVifusDzMm6z16R
yTyJDGoR0TeKmo3p+9NKhLAOubbUIZ7pr/uaX5Mhy+spq5sJaAr3fRub7AFOIy6X
lGfKvvAxmdaSz22hZzFXX8kSYiCmhfweEPnO/fDYEGtq1XibSdVzM3AAJO6o8rSj
nUlgp99vtw7tL99efEiMiTq+BEFnZHcZ5bGiLBgvstA8X9LSmByvyWuaYF5Rwken
vhfFFvXfGeGepVXczUwo+tgot1ZC8a+QuuvyZd5tKPnmD/0XXxM861V62qAOifeB
3BuLo2uVOPYWV4G4AIXDEkoSG1vdXURgZGCQF/sPPJae/kBOtGssWKJayIwXQS1y
V3HFyqurtib2JSzHeSixqoeleq2qwbX/6EyjgIFzd9kq/bH4se4RDT5nfelz5fLl
hv6l/95NMV+SiGyPZMU3yYRv9+ydX2SJ5Vy8oP+CowYRyZZWXgIf830d4gwUNz7w
c8bTVQJDKp5meHKNJteWuqsR3WvlWVU7+17hu1EEkU5mToxIbMS4i6okNm/sJL1O
ehyulbVIa6yq5FMUwH/gF5LceDyyJ2Zo92g5kHZDHXj8+vjbcuMzaHSCw6XBhgHf
Zswv+0YlXTtEOJCfDXfKlgIYUBS8gYyv14oGfD5Wuui2WBmOjd+FdD/8GZ2+jE/U
aS8W8pLXS1uDSQgviAkqArVNGl911CtOVHEzjEtVTYNM04yCGv2DVLqvHyZJQz4q
QvQxW+7VcC8ymnQLyk0qhvEt+TWe26p0lN0oXlW6awdCbhKSB3UeJ3FNu3pO5z/b
irvusYkN5TWqW5ItP5yZKFNSfg4RNYrq2bKr5B9z9Gg1CB/YnXmCmwyr1KlEgXT3
Du1oscF8QRsR/RgOhc5SgZv75MCx+82SzAhUToIziAthlOepwl49APfoQdcG70PK
mnRq/YDjRBpR8dlyuuTV3pnl9pVdk9gyUOtuCNsVF+NAh1xpOa9P053cwRI0tnAw
brwEAvXkfw+XYn8npi2qYPNsWyMnM6nPELPf+ZVTJyqWouFFS4UNc37QhqDTv20O
Gk1Ux40sO2cRsE7KGBU8bFrSfF6x4H8MpVpDh34SWUijFAMZf2nM0eRX9eWrIQgO
qKmPEgeWeO/Av5l1/v8jb3FGVztcn+XESh4nG8CiqkO9qWJKrkVOYCxd6fTa1o7w
DZYX8tfkZvxOh6kU/UlT3go+eZ/pWaCciqtfa8T8Au/syclwddGJdGDTP3c4INGI
nZmwO+7p/YMIp1PtAzsdDFq7KjHSwKWb1VNZQeYCSiarS+xiJAChFk8dUnK4l4BX
tdt3OITvQReRdsZDf7ywoXcZUkYPi37ntFxTxoG/qA/nkuvQ6nMeXT3TV3C9y4i0
9TPNAUBhR/3RR0koGmeuCCfvszM44FtsLfNb/KYyIdclDp4caPcYes5GQaejqRcG
SAwlAv0JLgrzFI1jV6pzowtV0Rbdda+0ri7R1dOkHkrAXqwmQQS6ZVrrkZsqaKnK
77BNI+nF9DsWW4ltiueTv0eWlsvQuBHYvwxhk0S8ay8Wdf3JvLTquR23XZokhILA
OOUHEl99ULMBamh8exFiVznh2xHK3s7A3N6BZFNsdQrHpolrqWbA2AGjafAW2gmQ
nkLLAEm1mU/WgLVNAoxSq3alITPqZGQM7AOX2JEv9hXP/Abd73Ow0eRw3waClEKz
QK2iN1O3HBamtynMf6LV6ZsSzZDIkz4Zg/zvgy6IUxzmRz+S6PJK1EPdkkFw0RpV
3hRMyLrGhWhZhFl9txn4zFtis4M+AUKbcU7nyaNSq2Xc3b7SaXGiD9NT83KpdIBn
rsDDaxiWW5IKygNUSbhYh/rCGyfO1kA4VvbZKCmJrLngyeMpkcXdelqXk8JujVxO
qQHJy4gEaUUfantIEJD+laA1tWhslVkfNgqrmIiLeGyGtDZJIovzltG7G+bhyWcR
RtWrFraIsvLeb0vcbHcN0JYRumeXDcafvjwgfVvUTO7A1l2VJkyZbWJ50PxvIXQb
Qp0HHC6o8NT3yKxfQB6Sfq1cHPpqy/nIOKluk3N0cbATr8n/vkB1PUjDP8TqO5qC
gO5uX+DP2rrniSg5unWM68RkN1q8+iEvhb/mavJjZKgCfQk1gBOMrQ2uy7SLcz5I
6UxjwIbdeIXGiN5VH8o0ctIjY1gbr4JGCRtZP4wRQSs4Mh2U+EszbGL5RuokRf2u
F842tdRQa1ztcP+7/01UvNHDU3ucrAcVHr6ow2xNTwq4FtUJJ/pY3UN31xAGUDIi
Vd3ctE1h0IZcAmsBBdJPfHNe7l7Q6UAI3GkyPmWoqYpM+MYpSIfpW9bW9wJHX134
Y4PFKpxUyo0mUYhM/zyVNoBd9odsCSVoQ+TwRl7/Sau9OL1wwdbVQPbB88YqnZWb
Kj2h7wdJajPs1o5gYZDA2PxtLMURv32Fc4DX4eJKRvWChFOpLBQLk7iVTxIswmHB
gqsF/SENhDXA1vEUyktO7s20cwLNQKtavrMjJ1odZKYRS7euv3Sv1oLDnHpnTq4L
kEf3zqK8vEeiVs6C3nCvfAnL2FNiBVALMXSx4bGAIfxoqg7mWIdQMbWwUvtT64p0
0EaP4ZD/JlDd2Ht+VPBAvVxuTiMnt4fgtDoHx/PH7EcQ9LhBtY9czFMOP/3pXafd
WGs7Hwqwu5Bg2okCZrlxIAEP/+nnfvqbfWtoaQQcMCDSKHEcwzBRYkWHmOWPFicX
96lgCr2nAftyCM4mxQncJCM9Y/f5oLiuc7Y42UX7Mih/KoVjOYttvlRRZaMfHi0I
KoNeMeI3KyUQ5LjqKn6onS9wHPVdFJF27uC2tDHFcLEhz0HvWE9HxBsRSbkTNaXs
YF3EJ6iuuyYb6CW/JlLFhuZGtuKGA/Pbtmav+gsODiGgeyNA4mEXM5xeXHm6g47z
ztzYuCwa3osCT88zNRy9ChlM2IPUtFPGqiIQZvnnebmR6lgK8SJxapioCbVO+5UV
the99ZAxVrNWg2iLsoGCgrw6sSiKDE1Isz1AcWxNQmQzEndJgd2Xxt+NyM9N1jGY
2WrpkvvjNW0TsElD3xKopXwVj5BRSGvYWHM7hAbRfOurAefwsaqxs6lFJRc4I7Yw
ZbdQbA3C+K+kPEAcBh8mxtvu2ei99ORcGZXS+pgE8p9b0R7QblTplCBNuTgXETnD
RDU4u3geKr29RarE4dAO9ICos+aWf3SH6MHX+kmuaWEXMOrtx/dxXorQukrkNl50
A6xVToAO1G5XWYF1DIPZ2L9PAm8oG3LqiyHVGYO0oQFR18WCu6r56Sfo2xwqjfgZ
TjMzmEOHyEPR6GW0z83QsCixND/gEHwO59uHQTQDSi+u/SsdVsayWxM08OG+Mx9c
xcBPgaLbGLSryeR37PLb5YAi62nTbmizDnz4ZGbqbSgO6N/g4Q25vnfMOZejDdd/
VUUKEkDGmbrW4hH5f5Lvg8GRg271NkWulh5f4sEZx6zspXL/CwZAll/1NC0lEbiL
57mWhO6O7ukVrIGQU8Aq77B+gtD60TZJenhmVvE+aSbjb/O5fsTdhm8JBVSZFZdQ
DHc7wQCVcbLKeD3s6/ZYDQXJc+YAIGZ0pNU4n/5FM4cEVaoVoQlx6q+kHMM499py
yQM+fITVF8sNeu1kVeNP5jFO8zUAc2zyi+cmeic0Kbbgq55mwkRVvC6+T/VIBV5E
hidmWpQNbuBjzb7bzQUQTtKmD4tMTz79OaY1pwSC16/HyPdYiqUtPKmNnJnim2af
FVfmb2KXkGtbAPmXmGqkc20U+x2u84lw7uk3RXry5aVWXw0BpXpWil3jRIcu40FD
pZ5ZdWqcZ7zCGygV42WCBeN2lW6epb+uKeVJ3sgO+6ahD4/Pr6k/A5rBQUZQfEsg
HbOawS58l51+xVgE0As5aV5iYm9zRwypyH7H/4KYMiQMpnWixPD1OWaRkOdmRDfw
yOtfm1mio2lvPU4IEM4N1guh3/YTaBHt//FB459PT2KkqU465xQJTU7VHgc3P1Un
DSmqNOyWAkmKf4dVrZ5e2hi4uHTFbqd1lwgvnnzgauSehvi8f18Ku6Q/ZukENkdY
uRh9KFmQta98TgN/dtRpyY6QYiRAJ6mj9UJ0tIUnM34LSBqhIc1omj9pGZrjk594
0qAq/TOFt95lf+Q62y9/YQvhaLharnBpuVr35w1A+Ghl6InvCjdQCeutGhaMdPNm
wiU22Z8/4Q2vxn6HSlo4BboPNJSXRKzz0eWmiFHFEw3OWd1tAWebGt2HJL6XjD8J
iEKxswqP2g4DP6s9DjTQQ1Zxvt24/nuz3Ta+p4P4LX12Yh5RGDKUTqo7W3r1EPC+
pyk7hoCorBiW1np64/WtM4z3g/BfpkGO7IzjZRjKMapW5k+oPWuqBCMBVOPqxiVR
2/GO4DJGB8q5oo6OEnVawL8xeIOVxQ71njAjOKLPawYmOhTftP+siNTubsmzFSmL
7B2HAgj9XCVO9dNQ0oveO941YZl2jAB724Nu0KEd3HLUizbFgmtAkItIkN4fUTLF
9ZWG/EkCvjckm+7uadDpTSv7XWh5K/FZ+33X+itswJFf88HChAwlJf1M5BTsCiqJ
8v+NtJZKRzaRLsnSa0iCj2QOIjy0CsAve5biGv97PqCirsk41WV38g2BxRaxQY11
f2ky1jnDMcjo5EDegOvOsSl01Y7sXP3bNjiPqnlDQiLYI2PdR+vlSaSmkmiie/L6
61yU9w+LgAd3wnYqOZh4z8JpmzYI1fwdrpz1CD8YUQuWTI7Igm8PgBQvSjduwLho
dNRVtWh05KTpHCIuRuv9XuRG/crXAf0WuXSq4GXxUu/r02Kl/64WbIMo6Ja++W0/
pmD+xgGpFKKq5x9jPp7lpQ0Pwhbl6TDGdekUa2b55chZsDlKFbOK0J2O6P9cELwt
m4q9yXvv1h4GnrTwAIPeyUkLwX7PlKaANqjUwN90M5EiuiJd0xl5dg242Uuoa9BK
TCn5c38XJ0QtC1GOCUlEL7LXwMfp68Nm8n6AvjPpVQNyWJMyb3w4+y2vk2WBPHVy
B/noMQOqrsEWvJubk8G/FR2dJGD+yoNZTANZdkjdRAz6D/CZppC6q7XdzAzFPLTR
VDdEdoA/DNWuHajF9gR5/cex1xH+0Lo11ALJN39IToNSExTyqNj6UUyIa7D9j571
sL4lICyWKsg0O7uQf8UE3evoUOfSpD/uOgBp2Rw0YV0VLn3yRyCg/qTJk/yArgcB
r3bxuUx31Itb6Va9avrUrle92wj0FvhswxoPceSOJu3YjmHGsHNmK6d2ijKVofE9
vFsq2zq8c8IP/7khVAk+2IGKM1t8tWnpc5x7Huo0aGs2oJ2UZTruKMufMJ2nzJmJ
+epqUBi4BkkgQFUIFy5Amc5l2cz3GvxqtK3z/MZMqUw2afxUQroeodXHVQgrF1ei
WOdcbgNP7QXfjEUw3IOZEWxsjPgnT8DQidddwGjRmmUzaLn4oRFOKcKuuh1ZINgc
COVlD1gNuxdVBv6EPKOeNUWTa+1OpJU1TZmPaXGvwYL16NrIegBzt9HlID8RSxec
bI26Xqf+eJgeTon+7S2Mw/BO/ZQrRcxroW4Mh8HHLll0db8UPHfpFn2t6dx6/kRi
G4Ikj1PCYpd68dAWthC3yFckERjr2tmPFcK+S9/lMhsRx7h3I2+CLooB2KuGVufy
hffoD40757p3QiMUzV+F1LLnPBOVSddcbLQ6HSDIYkkndUDkztOwuA95VshC98gO
nYZUVuqLzErYKi8YLAVq4mUy4zjZdzlm7p6trUrE/7BK9o9akeTq9QtrlXi1TQRy
UnUHkZdzcf67dIJFAIy8S8/B1x1dfvgBBZSrpw3wAFyUnrFzYp1R56YDTxU1Buja
CttLm0B99au5YIJrslhR3Rjky0Qkmcu1OYDQW0aFL3BSfzWgFFVPwif7uVg9o8Au
p2j8DlLuz+PW585FZt6M8P1otOZM4cbazW3DUD0VcPG4ivTPG/8WeMI0ZJ2C2Zw2
OcvUq1MPVJ3NWU9jwOQvTWA5ufJEUvlAToODgUD0neqZ8gTDlsCGsFrcRaYs43+l
EA2GisE1amdNJ4F5L4kh91YUrcIimIyD1qfJEGQPCELPaNTT8rRLn/R9GuEXvEkq
jAq8iCFrGqUq5zq7ZBWNHfD+weL+QFAjuwwIZO11429u6U+zKWy7EG8kKTx9mCla
K5HOWNAta86UBTWHhx41mN1Uv67srqKFvm5hjjfuU5r6rTifnBLoAasmC7EJQQ8t
+frnYV3dsonf+f58yW/oV6fKInlKoAyP76A2Y9PSZ3AwiCOIJ1UpmZ0pi7I+mhio
kGnwthfCoWSA88O4lVgwRVzXY145NT/OkmoT/ti4fllLTO+W9lOZ6POpbLrrxnTd
rEwzfiw2FzqsjaXM4fmR8V6oA/oFbu6I63WZtoGYqYseyKoPglcES8fngIh9+oE4
S5tWfhApvQJuLTWX68c1S/Eu8aiIwoXYIsUKGDDasguXttmJdpsxX9uGYn8wqknk
2coLtEg4IU9IAopRtlogVpVWyoUMnwUd9BFc7nxvg0EeyT/Rl0ug1GeVnztcYe7i
l6snr+guG5DguQ9lBghOToJ7ZHY3NFFcroyQOESkLUBSepuPEcqSAeklhvb57MMz
Nr6L3ICkticA3l8hNcdGBLYy/x8yXJtXpJSuUdlRkP9HhcT5LxjzcyRgheQYVDqT
mHGysW0gqna0yRMTOoGjU41O4iZuHEFUyRWNN2XUxQ74E6LXfX0vU7o3PFBBQ/5I
2prBh+E3AhM3m+dlxed4VgURFeiNtlV1AneK7VJcY3vrxoPWNYbu6W0i+HxBfaHN
NclDpsVGFHH+a953GFa2CR+5p9/33tg4in/2Wgge+VTFMS+lWN8nbXmleHmPrza1
3WXyaZIb6n7F6ORwcY3mkMx3TUZrGzDSPP2vDbb0zB4HZoaL2+7E4PMVFz5H1oqt
e6jHrR24vYjuPgPqBWmGqS1bMAe9EcuRUObE+qZQcy2EuYg8Upiy+gnZm59DIFqy
4ewl+6ANQBq5MkTBTI6vcKNblRE0qMLw5domIr6KVjhSprMWqVaBOHTHzyDU6U8W
Qwfdd+xJ6SFFiPnaGqQnFMwrXuAsD0hWn4PeS8hJnLUNFStPNQlmqXLNaFaAAQEw
AY7mpHdWji844F0NTz6nHkobk0XfLE/Gzgnd2YVRn5S7KcWZ99/S8ZJwJ/BGdhVR
b9a3NLA7oSoP2VGno1d4+28eWC9ljK9YSoTvx7+sl+LXw9dwCh+FBjoM/shlr3kH
D8GxE63Hb9Ck1UM0O8RWwAuUjnTaLLrmbKJ9dg7KTu2z8KdLzhNHLKdHGtnn4I6q
Eb4caN46s+tfm6GiLco7tRzHOfOpO2HL/rsZNgfxsfo7Po3Xa0hgwdl/9Gi2i0Ww
GQVnwLfjDxRLGE883GizpANCkIsJL7Ud88DUMQekBICxHhBoXyPgzGGdka6AGuQ5
EXLYYdLmpWLR0pBw0mWmBlWzPclq7IR0L3GmR2vr7RdzLQ7OIX1LPklzj+u87bIp
B5TNOwUh9bfIjZ+CMsYUQwYQUDQ+VEPzRE8XTf3a37YbXBuYjZMDYkAXaLu+TZey
CvFQqoyeEFew+Xb12aUIiG757KOoQq4NRJp7tLtuSy3+VEVO0a26oUfgf5/lxe/X
Fu78GqwdbhiKPzeLdT00JtqWpfS9KYrNRhRgWczcWnYFJvw+kqPu2srIo8tsKkG2
vrUL0FxEx8Ok69Hc3z99FOrNvVH01n+N4j93cwvEJvtbPRBcswNjDyRH0UGRwZNf
EptoGIwbh2llAW6q8vOy+Erl/u0HjF0Oh2W8rWdg8h2chzj2ng2t1LZpaAceDihv
uAAtaun1qIwslZkmO8ZhedFvZv3ib74B+6Sr516XEk59LjGsYkmus2gC0RwA4sWI
Bpp/bsoJxJ2X92pqNDY6NqcwOqDmsYjGfAZpUOCTmbB/tRtLCWtt1NjHFFVTeNGq
hmxfQlDRxGoHUiUY8dz2lMv8Exh3moqQYdXcbTrF2xpRavVXDcA6dramjm1M1L7e
8fR8iw6ELGiY4rHMi/vhV9qRY1CVG9cTu5+vAAG6g2e6ejWqlXLjfzSf/iI6FxTG
ziwZT4BLJy9QwFdDTZ+mm3eBG77Gz3yRw1aNk83WlZYjNCXYdIDMyClTjQzr6lyT
J/3W7aDClq4jjhvSM1cN94558I5Z2u1tG+LAdKZ5Rv0r0MWk2yYo9IHgcdpP730b
xin/Q+P7emUN8BiU0WJipn7RM5ADrkwB5lAmSI9575wzUnq3p4G9tsETLpanBFtI
X9NhSKuhaPeutiVtqvh5b1ptxImrtWWrjA3lSWpyl6kiCCQ7bVcON2r5TYWRGSOo
meCiaYK6ZTKH61hWIesMXHvgmLgJffBjnXnhJiGfQVx98Hlg5CPzxAPPwg9Owc+y
pA4uikzG3pYGJYsSXRkg/2Vb4M11070rNiNxH15l78e8DEEyDi27QP5ht2O9VwM0
hZtmhPtGBtAXSD2HAUPEVy5UwgOLhhNz+sMLoRNUKA5cJLvBGuQffdDTzXVeMqQM
ziAlJvmzHIL97UzemZlUd4pOdymFbGmuQWX5XHGirpGq/OF4fuA7wDTAfEel2Whi
NqfyN0CTiWQPt2I6GxmC0B5M01gyAHHFX1fQfzrkbwMbGQ/GKL9qkCd/3vMbMAVI
xKnrFJHf0hMKxORyE7aCJXkA55X46ZtQ9dQpVu7pKF46OFSuNLQye1p1vxuRp2iz
Q6FNgKnM1P5x+f4gsmFXkL/HcntIp8pkG+/gMQIcrrRC23J7l6eq1zcTigbEGwt+
+xbGZC5A3tEgXT7+NRfCIWQ2Cd1CPsM+W2XZw6osJyggzDa0dGC6p8tmuS7Z5mqe
C50XalssSX70lPtAFxtLg2tBsQY0k0/4fa9vzcKgOReKfOTgaW+ViFlcJ3+ddUO3
3K5pG+Me2X/i8t4Kz/pEVIy9xMlSIfuAf5wRaRk35JgQRCz+PUch3+lbzQNRT9+f
AN4sSBqxsnAqRtKqBzemhO5R7CfZm5DJL9bHmuZAZLM6wa+69DBI68usuywC/bYY
BnODjPYn6GIwb4FxmtTJevX+DIPNmIQtrPYbJN0TbX3vzuu79LbcO9ruzie2zWwG
PW/JhZRIbXa1lOB2z4ofzkFzuW1lbmTrq+UJ37WaGorvtrC0u7AzLdNRdpt7Uiaa
EDdkJ/J2KRJ85vJgQfLEt3aMzV3V8XE8cB/efkFcxtvp4pIahjBWaUOupmFfwEAn
nlNGd15hhDYeSgX0oxtxLhBRVw0lBdZpNrJmwVVj+LX8KZ19aY0+EgXLwireysX/
btGaWYUbKlK5lo+ixjfeA27Hu9iamiO6QVXwVK6Y0YCNS20asuwqRhC+zPPKKMB4
p+5SFmfFfZ2t/kwQT8jR+wztj9oCakjxaIDXkyY/OWj87y1hsdXDDVLnubP336JK
C4MRdKm0F0jjnavVMHmJanqGdS8Z58rJR/MA2EqizFOdnAAcjM1N3RysC4vcOD7/
4zQg0hlRY3pHMbSEd4QmoYD+H77dxqyVEEfgHySn4bUn2VBI/KIyQ1y6QLnYk3p7
zXM6HOe/2NN7pWsfk2DukvfndaC3LyT8WCTx3aTqTm+2vFYDb+BoofManm8ydoIB
ga81kwYLiHYOgufINOlwT9SnNNLxGpz9HYPh0wKcLLG0KKHM8YH7Xv38GLmJmbn1
coL1uh+XCYFykxJ3xkZgtdG5XibatChNRe5j/kdNtaBPjotRZkPihf+6+68l0+ui
E6P/C+J4mX8a4ihqWwd8wHOeBVBiffDMHQUK5hf74eLeDpmTUDKYWyeT3VQ1eJRx
+V7LOM07zPcoXxsh3oJ8ir8g1AdmBkvhCgcOMhU1EnI1F8m7vRTaMqnZyV5YKcE8
BG+TG9DJ9OhQH6s38yG4szEbMlzE8386+7k+uzGcB6AbYjtyJj43UgWGu4jkJIht
aizVvFkiCKRNuYUNyQlfOBxkrhy3P+2SLHmCWA+We/ZYRCOsJHdf4NNAMLe/MEpI
2aUwfJLwoTFoHkv0tF7LWWMwytVKf30+aA1hsyrTgBto8yScSuv5+3pjWOJf78VK
dwFN/QDvWYVPyLWmciJrUxObX4sWOmgJ5Of+XJA9UZAHv5BeLttwwqmmHFoFcRpM
IC81IWugOwZf6IQKDCWQ37f97VLBsBDEvCt8m+9czNI6ShsH2XPJAPf7y1P8oAL6
YJ3fGYo0d1eYJND3BNEqx34ksFW+CNdF3LiNzpHXv0yDryRVxf/87dsR7sBtFE+g
aVxm6Rf8MbUYA52SSmWRm/Yw4MUc+mRDMXLt9Lfo9hkHgWGHaFw9Lj2dRdZvSlpT
LfKsd8aqeF2lAGV/DHHmXIfz71sBWNC3wmo7RyDYdAyppjPXS+fK131kAcVGQ1C/
4TZ7dtJpN7+/hclfwmUmSJkgon4DLg98hdTElbTnqxgqgMVu4UXsdZ6RaOIlpyDk
+dZSLLrmm0Wb6xqaNoWayOXdopHOHlL9bbiB//Eu5FxRXqomtdApvJaZp+jgiWOe
I19RqJc9AoFlIRBC9aRAP9/MaGJB2XStbwFcibuZsiveHXeFsNSLnogos7jD4N8Q
c5uw9DKAnfKRuKyvcwrEwb20ydEVsEzSgYMPuCyhehmWoSNTBzPWabXcM4KYV5Hd
LP1o845PcQqIVTe3AaKZOgXXKR3z9MIV1t4RJrg575XhJfJ6QqPI2gkrSFjuxm1J
S+KV8pBsfdAUQEY5x7bmw5bUxx9ms6XGGhVaNEgC+lioA/xzUKJ81/HvSBBc88RT
T7wGsIT02SBxMIJfQeAEwv0WL1rk4iDiBiv+H8HyUPRNVMFy7vXMNI7RHvnMQTGK
jVcK6CEn8y3/Fuan44UB49dRcKheC38W6OzicSn6zkKByuj6v9ErV8jdafKXTYLQ
3eCR6E5ppkATyNXNTiRxbzCSb2laaxYH3P3JJ6Xx4IuajDAPXEDNmSjdwiwizkuK
2fneAPcz3iYjK0hM3MexT7cgfNVMYeTB+RSVr0C9eAzHysg1MjOGWz3v5TNCOK+U
+gw85k7PIZ8uesP9fxaUZZvLr0X/Ln+kOzz5qkYk2lwwt4Qlor62a4MRodcLB8g1
ztEVpRryfkUyqN5UZQwVNQ3khfyjQVECiMuC72QZe50LZAS7JP1ZmG8tEAB8GueC
nacP6eJiUA3YjqaUOTjxFHSEIREzLsoo+/WvJQCuJlSVxRvtBxklhUsqr3Rq3a41
sV9wxPv/ctE7RrGirTY5HZxg9vzsirqsDXVZ7/B9v7hI/bOhU4KW7ocsDrSVHP6T
WADx3UIRQUEkMN9KV1qlOy5/CrKWU3ySTssBtt5tSZJqlGp9J/5mWr+g3iX0IA+N
KszJldLaXXzGtihVwaNSmf6KZzl5BuszExiSRu98mGctf4m+w+0bTI3TnD5D4gvt
Bmn2eIJd/A/C3+aJy+QYH31T8DJc6Xdihh1oBgy3OqolrCMgQkJ9xSMGQvPDFYy8
CzyJzhjoh8XyujpKjUQZgpcaZb5MdFV20bEl267cWsvkIg6zQioCuVyD4zwh+3ga
D3JHwpDugEPxvtGLjXbm/jvZdO2obmkwdGv9giuaILB+ImLU5Zu7St4Y2eqUQUAu
DLp1Z5THpIJzMon+7jAMqQ7TMvGvLbXdTSg8vjv6TRzBY74aaBfUzGosGtGAXGqy
VedJ6LZ3mFocGoDjRXVyjGjc/JBjOMlT6ffY91q6V1nx4xGDFAaIRyZn65UB7lG8
depz6anmaLJf+FL455hvx3CHuvsDNtvclzOwd+7r/1o8wvOGV6m1f6XnaaYF04W4
UX3wP6kj7w9sQhwN+01CgjvX0DqZ1wbpE5qppUgpUvS3ZBUwO0ccQYn6pZT0IsIE
E18HJR9yvNi5mTe76vp7DqSzEqAcTx5/z6rZmYlXtLcgKEBDCT4gXf6zd1+BPG7g
senqRK2hbcIy/SqHDqvxJDIFNH9zlldaky6TAjMOz4TeqjmVb5A1ZBcTmcQIBZYb
wsOTKtCx9UKjKxvqgso2BDV6sKSM8+Jqb3/yHcULzfDH7eQ6xAOZn/HrH9kQLCAf
1ovr91jhLdOPTSV2YsgNZCq9VithP9q70ch4A+pOTP9yzVsu4sSCy86EIGvF43zs
twd9mA82XJ6sOQYacZpO4Gah+BlESC8v5I7g5AHHVCkUqhrNYfPchfVKZzOfCDLS
kiQK3AsFIoEJ6L9jDisJp6wH1Elapcyr5HlhVuy/w4CbvG0ZCHPAKDLw2NkbHV8P
14nEZPc8qomHFVAxODwXgyEYuFrwjpVIq54mAoE92wNGCEZCbYkKcQmTIT2zPLFW
ncsTlqUYeRE6Z7qDNRiYeaDnqAxNNjqURlC9ssK+koDcjfVMM3hHGYl2IoSNqQHT
dsnlQwSo1A8gVHpLmwijmYcnNmfxDBn26F0o0ATc98Z8ov7myIbzQAiHG6ns2yEO
q7i3iCjlEQRx1X5MMRA3eTnds6HJfrZDRaFUiC6/LDVl8XgRbPCCQmo518Z7KM/u
Zn986pyWfqMpPyXXseykxRdeLfzA1owUuX0DqC++AMfgE2C94iBRmNM+FxRMiMfN
epccjq8k4ORft6uNB713R9Jzr8shVE5O9kD1B6icKbVZBzH57r/h+HB5eEzDRk3p
8SBmDi+7Qt/nXA5tRfWzhVroLE3goIyO4dQ4qNtdK3qkVCZvufF6VPm7qK4NJ8pL
SFTfg5tGgdE7jFaB49xIF/GYeGfD8SJBuq7upb0mBRf7SMl4RKzGypeaLzMoHiFE
UVIuLFflDcJ+1Klu7hhzVbgWXMMc4lRMtsv9StyAu7135DHrc6EsUtt5eGAyYdZB
vGW3hI6S7Yqlr/FztehWZ+cUf576N7AL6oRqLjx/vit/0P7hTEVytfQzqzazWiph
m8eoHrFaOmvA2xLjLW8LT+KKqXKsDd6dB1XaXpoNmDyyR8q2c4AJrme0mDwLIzP0
4Mid4RELtW5aokxCJ/wvayRp3z+oH7B8XOy4C+xY/EDt1Tnnd3DOmZIUYOUH7DeZ
RNzSNXjRPsVfpLvCQuoNDPWTa7bmgRQhVIBfveuro+LXrErvCVWPkMiK/+UiMKpC
xwHx4Ri7Q+XlvKbhqOgm5+2r5c6rO8WONqkxo7nCQeOdZtt7C1ZHvHYVJ6DNVR6z
Brx5xexp1D6Umn2YuSPRlrAm3aWkcXM5vtq3AWYIjsVBILK7+UCViBUGa6bKFxgA
4z02dsSxTLeYURvPZKJE0ENV/JvJP1/41qzS8x3vkyXh9EoTbe9/G0lpmLmxJcsn
A8dpW4+vUO5mSkeZscRldpSyViyNIfKfD2QPin5YoIht7d+t5P6cNOYhIYczD0Pp
e3B1x07qHJlFKOt5kG8kxhgZQPVtNKpmUMWa57F1k5TXnwzxfMJ+D1jTzsk0gkqn
eb3A0Pm3+J2j9As24sHyegGRRQmEF/AMwXDvtNERwBA5o3iHcivFpXTTCcDKX3Rj
oXHmfyP/N2jwg3PG+6ehfVZw+VbZv6Sx3WBycSBpvEkvt8uWcD75svTNtx8eL7W+
i+ch3UC6hk89uIvxw958/znL31iQGqCdgMxDx8Ac7R1EpJoG5GTVIx9zf0JLT8X4
BfCii2G/nEsS/YYch/BmaBDEpGCFSHApsXbjvGFtrgf+fYRmjtiioRuXzgac3P0b
9ewkC7v09Tx/EqebG6OfvcoSIRosWoVUDcd2Ips7+GUYHXAGC2Y3nqntCGWyKK+D
wyCzC7l671SwWr8Dj9OQTUFqZGwuypVC2i/fLsOclLZ4bSIyRmShz/9i/ndG0nv8
DTnl25HJBpiqmxV68GbUK742Svrc/tkkvXI8aMDoCgeqfCF/AY4Ijf3YVlPUCaGg
/lZ9OctK/r11KSGyR8MEMdjDWTKpf1jXJnKL/yC7Aabe5HtUUI5id+N1uw6Miv9t
gY7teLGRgOgGvvrw6X3sapgnBp5UdwRNsFZ6/Vhx+H2k6p+fRBmg0o9XS0SHwuW4
GHFTADFgaUCwNlATMs2kaiaBCyygERapeqBEm/qgFb7dw3hEDEgi+O4mvsrns4a0
KNRwivbFySNxEMg2g9yTpdSFeUryiy54mPrIKM38zHPoIRb3rwJ83t1XaiPo0Uf8
w+nObSrGX29aeLPSN5nTm7HdoO40w+qVEQ3o9BM61qW+YgXw1EUm5bH65Kptsf+I
rGHvq4MRoi+fejGmhTiNKvswNhR5DGg5JCf2Ub3VDqJbu+jK8IRzDs3rNI/4JeOb
JUt/F0Wn9QsmWEo/Sm/3mE4dGEezcafJ7Cq1ObMs1jUaHWbHPybrenf+oAKE1f0e
oomCVqP4kAvApVC3cpM91wNI5qNE3F71l+U5xZvmy41h4C95WmRojwyEn95SOjLV
eQZLqz0hJ2HdGrHxORbQ+Fn5zVw2tGkrRpE+0UJhaRicSAskE1WUvACyTDLi2dij
R4hZQ82+7WCVp0C1sCHuio7VQKPPs6pfNJYKOzmGhURXbYI1N408veUKtxQpbXd/
vUAxTTnnzCe5aDFRfM1uE7OMRrdnjXRubK7fZuMF3M6yTX3oRtjobPrI/2qw314c
X1KOS7oNi/pMVULtS6+pVNO13UlW7asxpnE7xs1fdNxhmWGo4vq76fGx9mfFD2Cp
VkilqDgF9C/fS255nrCQeHnE+Ccz2jhYsGBw6KcysNGuEmY7zAZqOxy51fMxLogc
x8okJyWMtEHqbgtyEJLTou52NqqEexT5HHzoXEaW422oZiTShfTPmz6X4rUu6sWf
6DEVAZICQ3Lk3DuFDeZHCOVybX4joQM7kvuKC7nOKpYdnUrchmE87xoaJcQ5EW1u
lq9mM03UK69A2kmhlXLpQnTsVS2b6W3EiSg47JLE/O6KPhxTM49SfSoaHkGtK5Pm
JAiKrxCmg1krGzNPRxnny3j04dHihnVkUPOQ+XxONnX2khQQFgO/pMds0hTnCvj7
q5TuJdf3GLyB2Z3ZgnIun6yoW044Ja0MTUbePvZJnvfNxIijk+fa6eO6l279r3TB
ccCrQQeEMzOZgwZknQsjf2sy4tcUWR3sO0fhYelENO2YYa5VQTzHjStHZcUAtkT0
ohQRd7emZr14MyS5jae+ubnDD8Xu14a94br4BeasqtXwhVwjN6AiVTpc2BUe934J
/ly32226eJQ6hote2QxLN8qs/7nCMZTkbnhBsS1LRjxvMAY6Zdlm0SkEO9o+WvNe
WZdMhRbQWLtsgwdfkrOoE6E1RYDjhqCRjMtVHvpxVzhjaXJL+NpKjDTlD59hqWN1
CT2uYkVHscJtlHmnuLgEyaduH97UmEzA+p9JbKTet+h2CoQH3mm46/MQWHudFVsa
NS+/x8rfr80Oc7PBVm4ghWMYCVYBzAh6t+lv4y0Y55hS2sdwIMCU8BcmUvIDgBCf
BHfoHDU7oXPerxCAiNp2IUTETl32hcO63HEaCRkPQqtVXiWkUfbexyb/Wcou3GXB
TEB/kOQUeV7fMhTguzStml0FFJcdNNxdKENQKpd2hfSG28Rt2VEM8XxQPk1xqULl
AMsRVkqouKyqNU/gyunMk9LZnnjs9h5F5NZwTZM+t0jTba+U8Mjc8QubO+tzZpE1
SrnX4KVP6DKZ/vzuPjwgWDPfZ46MyEBy33HWWZEDLEGoqCrQRwiZIat46BxtDajE
9ZLfRakUZbfzwOSunzPEXFeIHONPrKgA+mgIRYDZBxLW9MtwtKmFlc36yxk4rgAR
gSUNmJTCixPxqHCq67d1Q0/xML2r3qj1nlxIRr+Pou5TMoDj/TMM0zqk3pIGQtVj
2/0HRB8VlFxQFQ/DiufbLRMqiKwoRF4cugWfu8b+N6BlwuK1JIErCOAv4VUWEtGd
x3nq2PbatGky5ChsPcda1WuHnWPEpQuwPHFl+rMzzg7Hw0HBdku9+XzFs/N2VjUQ
9UdpcMAbE/Fu0FJWmPA9ip8HwDWJ2/2JTXt4y+SHB0GcvbUoXB0Z5BgxGibNpzAp
il3J59wlWFi3HhfOhpYBNAI+K07qX7Lz4uyryDoVixv6RTA8bl2w7vrL1HpmbR1l
N84ssf5FUd9OZAQ3tbBhgf/BCG/jLTozDMlFYFmGgCJ5kuz64SZk5/0pW9YTGJCx
5UuRvE1TzlrxLJ7/gzBJwP/hvw9zH0xOARnw/dPlUWrRhUI9O43tj9AzjQuY/+4F
5wf4WTNO2qBBJr1kts0qwHn80RxtxiAVqScMMFKjRstIi22m3DxCN0AVX/C8PDHf
8D/E2HUd3oLj4S/Ug7k+A6LEYcMGy+WnaVFdpnjlwWuh4glUPZ4xKnr523/YBL2W
lGArxP94zMywRz7Q3WEuI58IqT7wjICdYOk7tJEVJH7/l6RrwUH4v6zS1EzJOuJY
Ax9sJZZX8BobPJztIRO3U2L8b+FYxa3bzuPpcVUga+il55dgxGWGEONfST1JfR7J
wWzsIDQ3V8qgVhiTavoXZJMt9Wl3ZVrciEJMVXC6T36XviMPk3c9CMy+o/sR8KNk
GWvRHPjz4vXWdzcOGJXtmJDmQhpRwn6lySeOXZnYDxDNmbkt0xi/Zgb2IlZM40Hm
DMiqqUymkqPMDqUwpDJYE7bTR2TuaRWRbnJlyxSGeD4t/9FQkY+x7Km4CksMF0/R
Qm8t1NDe/FE+Z1mmwWo9hybSE/i4Q/xUzu/zRchzPD2U/RoHlv1N3CCUHJI6jUnl
8YOgJIWrdzdAjzi6olbhqevoVpa9gY5HqEbABS2cwJCrtVkbbxKhCkm4ylH4aBvI
okT8AJkwQLfE2QuFS3oOt+1XVsbnGPxtQFTMg4Pe38Fdj+VVREoRkA5MD66QS8Tu
0/8bHm8wtALV+E664jY2Ipciq20woifRQYEV/w3Wj/xm5OIPqdjpohlg5gFk9B1T
42vo5bbJIh4VxBRNsRz+URmVMFNHDWd5iwbH2HUnVuCDkUjHCKFiMvxY1KBkvY54
jXwMRZdbx4Y6AtkXlQgc7GB/BDNTWdcMbEALIhirO2yfVp12PfPoggpkqJcFEihw
tiSF0cRCQ09XQFaJH/K9TZ2QeKadC24ST7/83CbBTSlXhObfw18AYug/a7lL6kcq
fe6PESj/G9ELjBTpPMRGeE0MbqobeIoU9D8SdhrBBR+yWDuXBWoZjFjWDrRHU1YJ
faeSJbOeC4WEc/GFL4VC8KesvPGrcX0T3jeb5QuhijkTTFfbhGYdcFh+jf/GAlsY
NalUw4lyUJtO6ChtyHq/R436WL1Of3UbJk5oPmQKypi3wZHyEgoKnhLytpKvKOI4
uP6Y+MgH+lN4AaIKL0GYPLkJuxBJDgrxgYnLo3REb9PfCRuCE/F6QRds7cs9yWNC
Zobh/rbXwpiU+gfMsFSwvy3R7VMIRGZSwTqkEyGBKivYWy+9a/3dNMQk4xY6fGtX
modyybOSEp+YsoiPSly/4rEXa3xgydC6xCsE3HETz97b1G8GKhUx7Ye0vxs94/81
5VfWGsltpCh0sKKn1Pn9B6kh6LohdsAxTAu34g2SHtY4Jgl+AEw5s4m89elUnmwf
NWeIgoxNIx5RSeppiG1LLTD2T1x2wk96EEQWYa2mQPTsIYaNXwFSUIinezGVY/if
d8tiscP4bIEt0QLakg6TbrahdVdbC1qNCUbvQx33cJ99QhI3AohO9CJ+1QJ6ObVe
xcLe4pDvArOBp3Z++5m4OvUqVqVCtJCY8OJiBdfG2izIvgiSRmhVdXZTIIsLNA34
/BBvYDd8IAOqG9I3Dq8BBr0gabsOPkgCJt9Xuryk3gkOnHw8QM12unzBBw3QjFQ3
enbSzhI6OxIH1WdzTzfzto7Glg4jq8xtP/if8k3eMVRxY0RPL8kofrCd3xYEOb+s
bFTEGpW7pQHXAZimWxeJxMukBtpS/stYDuxwK3S2x0enKXXq1JFLcECsSc385sNT
8BendLsTpYdRyRY+TFkiG54q/p0+v6lNOgbX6hPvhKhG8jEVp9vk/nttleCTTLWR
wD13Rl8k69YqbRcBOwuBoxdfC4sSNQvTHNyWWYK7TFEv2bKg1E1q2jodiwkrNbbo
qJF+NsVM976a9y+TJZ4/+4K1D+yIIXBNAh0BaC9P5BNsiluPHGG+lA4M1uGNokVj
c8TPSX42ehciG6H/pEUxhWN8SPS/yUvFdWq0pZdBdTlRYgGjSA5bV7NFmja6DoTX
DUPkSMMBSTya+D3PlR9hQWKBB9rzP4vUP8r325w2enjXdv/0/yc/UvsU4a1jNNZx
e8LZODbmVyRdZGgkwGEwRRXqFCVwA3ehc7hUkerVFxmrSZbwxFmYZ4IQYn36WW+e
wT3RFQg8J7mpgah8Mjyf04pCK4fckjEnI160AtIwAyKfXpNTZ7+Bya32yjaqg48a
xHMR6Tblzlkz13Ky/tQBrAq7YSzhznQjgYqPqDbm1CN7jqlhX6fO5lI80uZKdbyE
r/60Gp12HJtSj+YLEvheYW331ZItAlD69GNzGF6z/SqYtJzO3dL42sffYTLBv9sb
DzQ1v//34a8ux6rwvpyCjmQ4Aq3b50zN+ae1sMtEARXgHOX2IezwlAOg6oeRHsrI
v8/ZhWN/EXNoDQ7yZ5mAp7iNw2FYigMGtkk6hOhTPeCvPAfL7gH0VLo14QYA8FLu
6jbpUprNUJmFKHBGBOTOTugk3GLUQo7eq+vzhF2fjJQ9uwTLVk5Ar2CCVQkl3Sdc
0QcnxAr/8VsOwnoKykZGKAwFQ80Kdl4vqL7eDEFWEEoOf/TwK5+jxN+yDqx8WKvE
5WiGhStjntkAn73aIWZXN8PwyCCo8wPgkSqlkXPRYV0/SYYf795cirZSIxfzvySD
aCIFKrIgOkBrjjdmIBGPrVTyPDoO4SXrJilh9pB6EH/W+MT0RBsYzjvLIU+1aOOr
6Da3Oxdzy7dh2QJRyh6c9DyGZDaZF6AUbQtitbVpfekAvAZ2lprk88IkEe8KkkSX
XBc2M6PByXL/vl9M7vm1RNia4pB9cDpLubpNGOVY5ytOaOVtGq5dhPOctEX4QemT
U53u71pVx1ZCzkbC81WTqZYNNFGi1VN21zLSPIroNWDtmmargazOWDZQSKYU1atG
bKoZ3EM7mfxpz4beYEoy3Wl7islhwyvoWfUBd72lEwhLL1T1JlytP+z2BiF+Vooz
Pl1skCwpF70z2O+zEaf5LsvaAyDA4TWFsH+CtRHdvKSjDpZervB77DNoswxRgUIo
1SfK3MojmKXn548CDb0RJcHKP6niwy09ugbZTfEGecI17qMY7C0Rf4CCrjAIiDne
dFpjxEyVhxS84KXMKZhqXSdXtg+IIZqEsWYOGRdajFbc9Q0+PXL8dOAd/AmRC2YI
MBGvY3fEPiA9QRFU19aJyBeMJUzHv9M4i5a+/qw0S6Vs5NYhKh1NQu75gs0b5YjO
2kYtuismO7b13dX3PouKtGmXLjBtpB3oEbtHh5ow2KvTjMuVw7NEGKNj1Hc4xPqC
DAV/TLppJzwgYfssMNQO8FPFbl2j5vUp0TIJwW3J680y5Pu5ePdNcsKjflinY6CN
K5zim30MD+++DjlO1GER9vntlyZhQHRa86h8Qno36U4x+/YYTGuA+Az6nTegzv2a
9tveuyn8ZCHgRDFh71Gk1KQce+5DsC8s0lAtosB3Dq1H+LRjpTJaqTSAcppuS4DA
te9HsCcxdMHOnkeRc6xNyCilbFqJ/E1vj9GcHjPupVGJ9mOmF4HkdMQ5MtlaBYLq
2csCkBFk2MMCQ0obZ+gFGGT0D+JmU7QJvdaPe4AUWmrIxTKCzk6foeXsVaQcFPCD
EuKAU3q8aDoLbKRj8MESQIAXiooa5zSnAVHocRjcmUw7C1RMTV8kWzZqNG7IlvBX
npXCKXofCR9WRp09EhAhIg9wBQNVcxMnsj5n9d9wnRvubvzGeFtFh+b9A3BNPadV
nHZpHtz0p/tHVz4Ct00QfzqHULeLxkI3D4hSxwfeWfyxJAONgtvinIUPIMI+/9JF
EIkTN2bccmpEo1SNoWyvyP14h2Fq7lRqhcnb1Ljp840hrrnt2dD4fDrGLn0ulc9/
t2qbawfviC2llZcOlMfFq7greb+LyVX+uNnvyZoLmQv6g2Zfi59UlVhBsan3d/ko
vEASkzU42w6RO0uUS1GG/cRoOvoFuEst+xXcQQOB2kDm7Oq6un16My/tcHfVznnf
g1LjabLb2waPvtVs+stoJuoO4Co59beKs98syu9oi+RG3KyUKHihoulZRq3jP6Pw
qJcWKAZ+RsMGoApOh7jkDUvnwamzOxEEDFHMGEMYXbAWZJMC8wEtlmwUGNBGKcQR
Saho0fo7Bi+J2azEEFkzyVmxuySa15rmrJ7NsveSuSwYEIWLJ+YGs0ByKCHLOxJM
/wKsVFws8UyLBxDevtUkTsOq9VUfT/xqoj8dim5WWqHEAfNZcvf6l8HilICaJniA
5Houk818/bmcSf1OLKf1P9+hzEB3P8B+Oh7HUX01uH37fBzUTqytiwa/SoyVeVij
dnHuG24R0FX+wrqxmw0IgQ/pnTnXk/PK3YIXnNeTBzOpdYolnSXbwYgf3Zpe229P
tlOsuTd28ayJSvaQJdmS9yFIYZ6Q928RsPdwHU1H57KXyMOCA1Hdruo/6HZedL5p
qnfisoPOqoj1kU0xd+iDYDQYnjzEg6NNVarVDx80Q8zb0aOfyvfljdslyN3/UbSJ
JrSiUJQLuB1AsQ9eZQkSGeAwBlmF79E0xLUQaoVZknp36C4myIDrHLPB6vn2DsoY
/IMZXCVvg++BvT6bpWIiTT/WT2G290oOuE7fJa7OxbN/ivnDg/Qt7C6DET7JY+24
uEe8iX4PGB8zJ+w4Hr0Rv+xca7UCQzNeM/VM9EG0X+dzWHr2FESgQcPrIb5995u6
7mfZ+56nxaPN2Hz6TXHvGAGkzNH2wIbz+YEDNnUz3Qwhx/0OJLrR3gMqT57/ZzW5
8Yt0jf6QpAjbcRUFMdJLMCqqEG61xN34td8Gl7ASXx1mN+tHx4mOBfwtAABFPgpb
pnKAmdD6VW2OsAzAvt7pdDDWUGGrPi75jM/2A6FFcn/vRAcfn6yvkvC+EVUPaaWN
nAoPSfS1QKbvo9Y73ioDAdkbAl0TerYxSLmNPgNLB7Oj1G1u0UiAYSqPCz5LHU2U
3hMQAZz+hEyLVPwARx6vgc7IyIh88Vg8SmIp44YHAhZKJFSMZhK1ux5duYCYb3rR
LS3PA3HbjwprVJ8SdiQMnWBvK0+PhReNiM+TsVFRQLWlOV15JsVv6oNcbda06Kf9
+8803rg2HXtylOtR0GVHh0krvdjCa+JqlGYI+gJ5WlvbYILP/X6I175TPsZPSpmM
au6qsi3Dk4s12EmcOzzEZujD3WnIE3nWuJA64x6/VhOHdVWhc8Htt2RDxwT58XJ8
x9EN5SF6GNnJ6+u2I7mbKGXQadPqTmK57ofXBsnjvb3kGMm6jtpNQNYf5DgP0nIm
MeSD6Sl007wTk8dlnG+vgP+JXgxSUoibjPzAlWdP9J1wApwJn8TtF3D3WdJi4ptK
xX/5jGqgbmcDSQjBJbs+2j1XGyQX0WlYoqomPnMFB/WKFhs9zfQJsv+vXHeiN4ql
1h+uE4YJLe22vk3Es0YF4znntzDkx1IqTl2M56ulkk0jHO9zTNTWAQFju0cl0t3b
3pSVGxDcqkmP27PyYBwkKh5/mfv95D0nA+Srnib1ADh9tPXfSrUyjP2yDZqRCBBf
QB7o8B0dxdjaXsjxBWcWROeXCibk9YoOs63itiVrEd74YgAsjeF+u+Bd9UbNEh09
hkBcq1va/AkHJ1JbzH7lnbhUWIvVlhbOOA3Wjg4mWnWlCBZEV17XGreroEXBtud3
zD0kJhY83nyE9gYYrTh9baOX5ldRq54KcTSKwGY5WOZjtWl+4WPtpOGr3dl35BBC
EWvRpZqxJamcTc+0JGfU1sBNp+gygYMSNMT5jhO0dLFqPvCa2gaT0Kzd9RI0I+a5
tsMbBcQiw08TQIDxlGN8rgYDLAMaQfVdXXMrRqdHnbtibXEdxjoaWItDTN2IFuKt
bvQvhSAQcxmCzgynRMmT1xEa4RpGkcoML4sN7frsXgi2VUfpQZ86R0c63chr0RY7
hSUSX6pFjgcF5N/ruBPlGx/fHCi36rDBLsN7X2PzKnhYpEC+9YYdk5wruohLzonV
UktknBv1S8XKRfbMVxlMozheNssDYtytlFDwNcmJkRWMFOGAqRZuGAdBUrOif9ME
Nu0MGbEdNOER1fxgt8ArbadmzxgYydIX3MpylbaogPd6Pm6DP5aD5WegmXL0UJo7
gQdFhVsBfm8BAlPUtSc0B8MESd9EmD/9Pe3xKn69mYd849/wzd732VfiPY1OBRDv
c6coWC74fKPRvWXZ7mFprUiKwWmQacY7fztefvStx3MwypFOGyUixB6xVNhQlclO
I3sEUB8NU5DGmjVtGrAWtgNw2mTwz0uUqcXP9mYSiVg50knpz/lO2GtXzcd6UjDE
s0zA+xY03URl50pe1RenBlaY3oH0ho0Zu7KPEpT1Tm3qeWsGS6TUiy11GUNEDtHk
qp7/4iC7Qifo7DZHTgAifrAHE6BdVaTrqElpfb5I5veQc50sO5veWgdWj0TfNIq/
K7vcktAJskxhPSk7+GYksqv/lIMIj5BnNtmdkOHS6tQPF66k2x0nGc5iM0uxbzhc
w85vFmAO2d9BBEAGWVnwIg5PdOw6X53cJqyv2xr9jgn1HxGMi9EgJuQ6rQElTAnX
/rXe9aNGTYJUm65mfifsSwyq//dAd1NdL7eOceDx/w/E87LJDCNrgPcfxvixl1BE
sNpz69zWc6I2e6ZgNrUI3kyWWhdEuiSo3q50O020BrxkhKtq2JxfEcNwiUxzne74
EOjqXe2HuPVvLRUi64NHPjByRs4hkF3IMuI79YjBsVMGzlsVj3J/4Bwi8muuFXSH
ID9pQWi4R9bd6P6I57iPWldjDKSWTwSjXz/ibNNEd7yVSHlY+yHEiXdZgIRBfDYI
q7hR32n4SuAnldUIfYxgTEBa8PcxyKZOQtCwHZaItpo7xUrH27Weu5dPm+6tWOrY
bZEZ/3ecZxWmDmL3UC5VgEmNxCmJnPZJvblDkpYfwiaztvkwBkDAAOjlW/wfh5Fu
ucocWFA9xN04dVex5bwfoMtQsviDIfqlI3a+ZUqrUHIaGFh5eKASIqzJlKhoGJbq
yNsewoLQWneUPN1ZLlBUYsxcsgtT9qFLK3+k/XgTI0mYh5oaRmvxOJ4YAb7hbwh+
K7/3FfTeN1BxMcmjpD/odkpZsEz9biXCc5PWqWNX7/qt22Wg49TRCtdnR8mzmPYm
djmtQLeEvRwOzFUkNthzsGVxFtURZ380DK2hM7MPljEdsUgq7E0XQLKvPxyseBs9
LHw/nCtrepooav6tBaovtrkQlAvAMk0ExMKnHxpj4QKYgXRnTyfLQgLfB10OukD5
Ps9NafMQh25Dhfs8fLZc2jwAITHDyRBTYVjWjh20uF7mNQ9SD1t0E2Y/j08H3Ulx
B6EWmE+t5cuc+3Ps0AACFKjV0O6Txt8a3zYNjHAXju2FVsfVVD89R+fsaZT5WEgp
rMXPTD2arv7ZPNBt2dqG4VxUVCcukFUE2tvIbPkmyVHlWtBbkAgnjWnXVKXMbZVN
qEvD/4PwwBC89vjsCWtpVjwRbLEO7KcQIl11U698lhgmvMwHHS6zgISI9aKaho9m
xEf0fhg6bHNDUeBxjZJb1d4eYFb++WCUrHJILDPbjm+8EucfNuzM3FQvHVSFZMYz
EcVak45RKp8MdaZHwqeaA26iZ+FoTWMD/PEilp7r7MacD25G9SCdu2PZ1OZtLx1r
gCyj94imIafrPbKiF5DjwtviEqUwmkfG+UuPtipEfDGYM8nzVz/u1g0P5VL5fYHh
t55LrkgEZAc89uQJjVPOv11zwMmB6p08fLdjPS1+JIvnVaPS+jM4tRYe7yibrn8L
pI7U0bQaIT/pY95fOvzRm4Cyg7UsU/wZyJizj7aFFAiAsXHcNI/qRY4LWuBfP5eX
xpgmb/P+OVPTKWOm6OUP8aFvN/1RGP1WgKVPC9p1yn5KDD4BSulh+T0Piat2wExU
D3iy0rHPynd+Bj3C2nV9OoiyJG6x0LX8jU2RpEtSGMnEwmJkaFtRx6nKpz12dAt6
vXuGBZLddW+1nRQDkmEb3I6fRDExLCkuG8UqO7fhWSyKZ9DCelsaLjcXNlRoS6XE
6x0cIxvG4jrTb2wrcpy9Qv9s7A1/mw21Fym6W5gePGh/pWBmqK1bk2vfCrQ6szAa
ZWRUUyJYOIXoEJ2JJbyo1kOzF8k2HaRwmi9vnrfkl45OlV44bPpKhikwwpeKhzrM
jHU6OkrExePSD8kxaFttFQ0DEgxshmERpTShIcDOwJrQsVmtf4unXdRnIXsmBAY7
M1evayfONajSYB8T5Xwozs1kUN6SqOwzIB1PoW2H3pb2Fy8ji9+Bm5/a5NddQuFY
0YbKN86NrElcuI92ZlJ0KmLEx/aISGvxEJkGqDcdzmOpx/Y9ZeSliASq3ICZKi5Q
ZMn6Hvpe7DBxmbCLUv0s4gn5HBjP/NUm9k5o9Wo1nb3O4y4vQZHpPvapn8e872Gy
kCcs3v6jULcJM9JjOZEIho1Ot0++xi1PH3JqFQbEnWq95hK0QIFLgSbm9jxiJKSM
lrFQqig59w3jc7EDbw3HdLy1yHJ+qpGEwfOPZG2wnir2h/YU6MhnZ35Jy2VIuHyf
3qGWNazJGlORNb47GUsWdMymRGJ3FjiTZ56Xt/ZmOt3ganPvcc7WQIRiEc2+sZb+
YejbDbnHxSa70ARlbP5tp7eQPLwrvD/xgY1CR67APxEUQoGNYsBTSMkwH3VJHb1S
m1QM7WngjcDki+Z5i3wYrQckrchNBJi5BLDIXnKas/KU3WbPo0ges6o28DxgMUCY
qCvI48n0BSiLdpOXxWZT9JFRUoT8shM7yBI1ItSBCxGq7gqmsi14HZDvTvOvtq+1
U0YJWRNda+ZLXPmEETg+7foCFO1LiPiDgBGSLxbcuLtNmTeoDpS/WFTY+B+99Kjt
YT4/S0jiPzG+ePIiJzdnINDOoTAVsykbfulJZigHZSL8jfd040Mb7Fgfet6R9vVD
m1Y0AIyxileCkJ6lWIXk8Hj+PbT88w5It5TolkdrujzVz45kPtjiEctTcoPOvx+u
a8NHn56/FCnBRZ8Rr1e6tTYeyNzJvazcPNJQ84eZfal7EOyUCnR6HARxJipr7v+W
8/mQZqa3C+9gS34p+/EaTipwSR7HNa8IqeX4QiQBHn9L3pSBklEXdqUpD0J9JW7O
VkijArCY3Xjyzc4j4d6d9iOZD5I+D2+fvuYmMp1TSIj5sh1Ag57Fk1dT502aVdRJ
bX4Pr0uMotp/bIwDjwoSRiZgob25le78UBscr08HbEMz4mqugiQzMAruzcWWp7N3
eNOXbIWMof/XI0w5R8LDhgHFHsmXp0v2AY2ibDe+Mmou2JaH5aoVUhvLJ1uN+vJ4
YQDQxhGyPV67ZwbUNEHjS544sbwGKP5j4Pn44Vt9Q52+Uv7ZC6BgbQGBOXLGNVIA
o6a8USWrwjf6tGd6BhFtq/N41C5VrktybH1VpXu0pZE7vUvlLfQyer67uU9WMh5i
BifcH+0/jGDU4cHJzq2VztKbEAaiXP7yDL8dwhOhCPI+7hC7jACVjBd2Le1+187n
yAhdk09GHpV91kLMqFD5hHWTA4E6vJozf05LT196ZRJfiNrWzMyIFxF6XwhSyxCG
K3ZXt94KwHV7XWiXH/+SLFTaKQrx3MK1GY2SJLBdfV/oMlBR894NP5xwKu8yOP12
1nsQ8c/zIeY2uTRiA8QnJLzpCIFg/udh+fGTXSlcDu/Sb5D1I2dH2+5Qeuxy7NqC
8CwFLCahDHOkZR8fWuM1D3bMLfL1PbvgXaeZM5/lG7iFMRofijNRqm8e0PQWZ/zF
gMMHU23KFuf9ad9W0Tm0tIP0gnTiJgs+vuPWYUPlmg3haFkch2DcRi5zNLhQuooc
ETfsc68FjCG3wfGp0pvc7KKLockSIpvS854hYnyu/ALf7W0pZvEjoKh7ab6VNsnx
IxxWGKcqp+J9pOCMtY3vcDZKu4GAQNhR9AxJrR9BRO6whYDDCKtkeJwE+YImC5cx
h13RMMwzXnTTZHLtCnMVJA4l6C5DIRdRLu2jjNHlcCOYCzq3ID3wqknr+6xZ68AM
OHk+K4QslyxH3uhIhSeBex7C1JbgM51UqUVE95PmRQcA1JGsMHO/RTR8/6iI5hK4
MrC720sUAL27a2ZrEOswnepQWdx1DsX23GRAZLM+6JJixH4baEKuBsgx9hN9Q7of
dxjOZzFqYDYL24c6/+ON74qWy0+0ys+sAIRW2ecAXJujjtrcDp0VP/x26Ey3S6gn
sHf1UGYs0OYAVQB0jiAE8BFD+05LAFnOKtoDHB+nbNj6qeQYm5hBE7ZnZNFR7Tj5
8eSlrDPMD2J4Dw/7qGAgno2+bf0cO45cW9V9QBRe+qsChPiJ3o+rvcx5vh9gExJ2
rJv9fxNegaIdoO/wA37nq7avdFaG+kQ5G81CW7gC2SqgQcWETFRIPt4h/It8wH+9
pI4lFayrR+Kj7UFNYEuHtfjVVzqgRKq20haVCx8iuM8W4N4bfcwhXUMCLmYCaYoL
NEPG+1n1VqxAZbRNwXaI5RfpJyrdEGu/9g1B5upGf5oEaAcw3V581oFH5JQnzMeu
BPmTKVu+OopV8rosv6P6QTT3ouElx3DC/gt36Z2Y8WIT/er15Wpr4Q4wZu51Nu0q
xSsnn/bmNfjHkaIKCndEQxgHiA006DQTx32jtxhXaTAZAiL6g3vWdGIqd/D0s1w9
ETVrWJV3eZLREkrDYZFxPy5X8NYm2qd9iLVYAqJQjk9hWpTKlGKZtpZ1g5jUk4xy
e9G1OyAxOXR3yyRv3Dil6XyLmnLLf4rah+xwikeO2FbG6uASJ/9VSPSZcs9mg+UM
o6wvHhhz8uVxGWmz9SHL7ShCAVlmgmkSVUhVztHGP6h3w6Vm6uwHgpmylZ74VvH3
BMH/sbjahDCFXHnRoUsRRLsDN79+tBeJfHqIHfWceK3Bm7MJlBuOe/WHIEam6Scl
0hUiw6vMZl9cb2Lh3I/5lH/rAPOaNBvHbVj75TiyChEH78WxdMkioLcPa0c8iYTR
9dxqPszJohJi8NXZv0XXVBd6utrRf5DISQB+tJpbUmiSngtOKhkdF19ljcKFdIk4
ZKpb5Oq+WDEpwyDO2XBCWySeV8cB2qTmIphpnjXugBl1AwJuLj2hItfSfOGDZbf0
0hyU531e9B02u3Bbs2WvzAN4vvVERSc+0+Vhil2S5bg0Oy942I+oaqm3LLUcSVG8
0+X3eikCebIpICe9flxfUgBa1PFOrbjvFQhOtF3ebNv3B7+23/UFyFGTblQSyRT4
dMtphzoEyC6nGWctzPueSuR7nJIuh7c8xRdh5DNK+SfQKHbYOT+odCJJUm9cqG1N
/pxKxnIvMokMYbYuzcQXd/XVe0MIYE0PSYrfjhcTAwvRt5L2JgEhLWadTZCr0/yI
tf0bcDXcEv9+zAYgxHRs0CpZChENZ7RV6FQwLxRAmDEyN1Oi2DoLllr4XpUm+xPD
ULR4RkkFw10VnO9q7e5Wbl+4yp4HR0p7xbL2Z8KdSiKRyY4G8r0oqFD3XKVh5/EY
BrpDRNmldHYky7dcVkwOZmGpIjOy+FeUWGk1+0jE6qG3Kk9tJ9zqtAFbDsUzJZLg
LdVx1X8GuxJdpmxBvQSCMhwJzgoWLVgPgslhJkrLfZxt2ZpkANi3vuWdfslX6yBY
XhSKbAGwARhLmPPv4ACdyl8JSSppabn8PcicrLa/TAIcVCyN9jJqzeHi72ckRj/h
BvHvD+uRXJPKxoJEQTWJZfvFXh2H8xNK8ZEBX+kOsIZ8C2yqUOj3GiMXiWB2Clzm
wJqBOcdGwO8+tw1H86r7uLN8DTSRhoRiYwuAZ6zXNy4ZM6oDqi9EnP/oAq2DAPpv
OvBJ9VO98jh8kAcxzU0BWkodn0h2DiWziwkYnpygxr4JGu6WlfIxnWLxWMfIq207
fuqqja9TEcZDE4XJolkoBSAoCpPkYgoZmvpY088Sb7fmb6op3JWgmYPrYZI+AAMc
rS6HtAMU45p/HdZMO2d+Yz1to5Db/VWoGfDZn9CeqtZimmyzRlruXrc3Bwhjh0vR
RgvQuwFKLyEddYE3UUaG277cdA6B61OC9F0VFDu9FvlEWrCmQvAj8Hz3xTQYkLmc
LRdcteztVS7CLvk2gqwl3SnDWQXB5Nde90+huQD4Vzz9YCfx6fhhzEkd3CTryPK3
VMGgWUQ5kj6WvkBTGogDSCsTjq8v2hh3OZBJ4S0Y5FU22poOJ4bJo/kfOyRQpxEh
PgndMMG8E72kVWS0VWUUR63tSiz9NlV+pNVQfpoM3g0FzXO1zXdspBaZC+9+LS9v
/6MTZ28S5cm6aRgTKS9z3iwKaiMGxTCGSgtT5y8sQMSz+dGjniyCwNwRC10JylKN
O45WDiVfVAs2wowpnAKCAPgKpE/W5LPAGdfpz1/izIX1jpyl4cdvLyJMaT3Rs3jn
Ye197VEF4BsDnnbOFUTWOrPT1guWuRuE7wnyXvbgSPWFLWlM42zreJnly9Nh49fc
tpS5rJih/ur0DrLU6GH5kkOU3OUGzzLi0eB1hCQsAKAbcAXidX1xbX3LxgS7pJYe
tMRxQhqDrPohsWOWudAcHuQcuEGnymTxGx7/uNCexhVjXECOenimmmNnH2EXcNM8
BSeF10tYnN1urNXtr5oW55eW0znhKw0nqsmvvDjue8HhEwbCx0jcyA6X5fDgEd+z
ORMcYAAGzyCWNBeeOGW9SPo0m9id1MDq2n0jfiWF/uP6HkONqzlVnvLpkSk9gNsU
P8PaFa7F3Lc6XbznB6nDukjMxQu5tnxi2l/G8yNiIPtrm+zlgXvVr0r1MCAgCStR
NJGWfd66sxWrnGg3wnCStlgpXoscvN1OV0IJFj4SG7BNnKv1yoqbnmuOCQpVfDMr
loPToEPiHhZ1Xv+1JYmftOF2t0JTELmuh3v+0H/Plyw5dYTzqmKEtkvL140E9HEP
/ArCyqT8ryY55v18X2EPUHrLNatj/Avg8eNO23PrsYaqnWkRR55DapHIasikC3h7
j+4xiveqb5avfnocBEoxJVKehmj2qYclCBnIlURgpI9TH1sLqYLv1x+s1BGVmERO
+J2heCGFBj9DTgtAAMIKFwN4RGab27dMPvaYEGWmxXz77Xrza8xPGTq15FYLfLup
b13jG3ssqn5a5r4uXQrHMi1BYKOusSwk1YT5mW6JRLuYvTUrlUqqyrOMVG44h7N6
sdmqRQXdXeiia+DNB8XcR7qmnZRTJH37xVCRINCJE8Vh/6JOlAAZeBfhjtUDqPF7
BxpLCSl2nxhlONTrx4ss1OUfMX2BoCXQjW9KgusOp4Cz702MeOfurfwOY3yv5wmX
48jNXMLZnSP+QGCyac6RY2IBqvRo8ontgWV6N4pMEqPHShh/bg+qT6ABRxu2HxRj
MtqzOb9zp1Xhky03cscs7XEuDYVVurFlvLu2dkuzWBRARn+Re1d6MHKEYDc4ajzC
AW/Ji5IZ2dnks+AeW1HIzoN0HVfqRogX+VISdzkA83SW3y5flbqdnUBO77+QB+qE
ZCYYFRu3G/mmGURjc7vYjB7LMdhOK61EaM0cK1TeZb1sP8y87tK+SBB4uh/uPldZ
XXb4sU1XCltXEC+rxpucSqMocMll6Mey9OlejbFk33KDHcqFhlzP0zvBMDa6PWfM
bdK0mbehIOmYVliEBhotqC2BVOLlx+J5hcF+1xsqIeEoCgZcGTqRSnshPO0H0SHS
v42+yyTOkaRHU8TrGVeA785YOgl/gv8Iw4RjCyZDVpHV3WusI80i8yeocJnjM0Ik
9z08GDA47CPoXuI5A6VG3TmeRFObZ9lyj1d+uyTiHSDzQK3WLm5Qo3VWPU6qmoQC
0bnrOOKk55uXJqYj2qi/qY25l3xQvrf6eAPMuaMDDabnH4JNIJgxrevKXmeyBiSY
uv1vkMB7n5h6Nwb36qZNeHRHiwOh2JwKucz8ypYDKsSlMA/a3pEmIMniLPY9VG14
9CZLIu2KZg5w67S5nei166p8krSdXAxp7nBh9DF5FT9WkI3FXS+iZPosX/KvKMQp
EWbu8Qqu5zrCNcq/AQ9QPEsdzff+rNk7DMoD71a829TNYXptFnqj5cAjhFKEEF8L
1GvyryBf7uLQ6OoOQTZJTlwKL1GQmTEsfACUEr8aNT6LZucrVLnPOxANCt8HTQPm
6Gu3BYwpoJHjRp3QV3DwpC+EtdtWCTxrLPEg5AP5oPZWtB1fZ198lAWJUVO3Dmjk
Vf8XS3dM+dFbkVjKYcIhmXsUUMVGqP1TBKkd9pVHjM4UwRfTBs4arWHYHHOYIBzk
rCf1cAXyWflQULCYVpyga6ouDjSo6370lzPJC/4H3Bq8o8DGHGffBGzot8KqRXJh
7RdUok0KGm4p0otefCIFAEwVgBMIJZchdP5fah/aJLNEuwbghzjzqlEtwsOcrAtl
mCuXsu88kpHbp7E1+4tZdLeILam2d78QQtKxrNyCuJhkFfvYr1Brc0ui2myV0AgK
7Re/bdGppAGoUUuQESh40bdWRwFAWwdu+deyVCqWyciWOHXzDP9Hr+a3eOzkPBSn
8CrHB8vE2II7SsxUhEGNNKpZhJhiLSlDxPliExIt6kYh/4xuEvtOXRopGiAJ+Hca
do2Gvk0WUyjIA5FEYu+di7WLJShqJ76bSm58wO2q26+E4F2rgOjI16IRBnKhbWkM
eMQa/56lcLQERQxBbS1rQnLbWTDTeN8zDuUmGP8KMubPQgrFhOPsjY8cCp9Vg7XZ
hlO1j+65TYqeHIwVjpxkQnG8YTPHEe2e2qnlIZk+MWrqtO3BHhJvSmxjuvRZEN1+
ebhWRn3UV8knsTGPOsRwy/suAloZFSezjGvDdbue28PRfY02DkRPgkQ40RVV2cwd
vUPRntC58D0odU1ecCGKbfNKgHv8Qnp3i+B42jwPUVBbp8jbJx5uIYO1Gng1RNa6
eLcHirdbjR5ip9AG57codrMXi+SOgzXsjZVn4OMr9NKRnJo+p+2QGzoJzAMz5/SV
tsRvqJxG+tWhoMY749vFYervRcflFLSyw2ardUNTyU8LtixBrNQyCK2u35xkrWOX
2ETxAS/ZBIgSMyGW+GThwXhFjpbw0ArW5H5CPHNnqQlNtNybf+IpzzLZvJN4Uhde
lYDltWYiTw0zNT0eExfFdbPgZdSIjeuy1sMbTfEIhCmErHd2FJyISp9eGagqeLvf
9hz//BhSolbh6MDnX9qBqMWsZKQhf4t0tyafvN1Ih7iP/ugGrQ0jeWMPGtHSVxWG
B1RoG4/cOlnElPR8T4w32G8jkfhfEeeLtVjY4OpnJCCExyOTKT+Q/yokGCljL8vR
5LXX+bBr5NhAeTKXd4D0gjv+C1e3Y9zIlh9i3j6erq+ZDoIpHPDF5zotwCQzHWgS
z59jLwv44ku5ITCBqCHCgo9S2kbiKvPegLcMCEwNnOAeJWv3sf+loFaOtGgQKe1K
GhQTC2FrZu07LWnwPaZId24nC6Yh9W4gPnaWzWELVKNTSN8mMVFGD5QaB+OWny+4
ddBJT7+gzpS5oG3rxBGiD3f2CmGRdmOhZUK1TXYdoPRTBwXu4yK8DDwqIZyeC9oh
gIkfEtcdsxpyMPD7DdS6fkO0tkH89knCNWofs0EEFCJtvC5ywtyP8QMGVIr23SwF
Zr2i5g9BXNf4R4mbh1GtLOG+nBr2OOFsdcxhV7kUIc6yOIsjwXyFVW1Kcz2hHIDe
vrU7lkUcjc2V2kSLGNuHgv+Rm8FakcTPkbSjhoVPtORaImFUwRH5DFRjkofgwrU5
hcDlOpCp15l6Iy6lUcmRzLnTmstGED/LmiU8Z1PL+/I4pKcQok84UoXabG46M82U
PNELA2aOeQo6wkpZAaFpvvNbmshx0YlT96xXFwozXBvhbom+MwjcegnI6KJWvpCD
XJy/gj4g79tCnzlw1lbnKGNTHzdxJtGkQrccxSrkwjHUMKHM6GWqtRQgsFdMbLcJ
MOL/lsbPApYt4OsvC8YNAnRteLmXYH+jSs/x6dqxdemnLcZ02ftMf9K0hkcW0ef5
USKMOJDwomTJmy1aNo0bLQle+TmwQcjNEhJWmb9HdzvqlEvfjUJ7JntBt8oWheKe
JtUcNoPgWx6EWFjWflWKl2xDRtTM4/pmSzfgU7u4rOwOS27BXLPttrao4OzZxELq
xPzHNp9iVLHm0NM9T0QI+BWAZbqSCUrTAmw2D3ePaVw5WWL92Y1zOuYYAIoM9KFP
qfc5qWB7kTK7gkwQVGMwEs0oSxKdi+FX0F21yDovqQgLNVoiJEFZu3bF06odnps5
dxwH2c05djmEpoUqU2jRqiQ4OVaDcbZaau+gaBmXqZnloY/PUMTz6d15wiITOA7K
L5qju/d+mJmBO6wxk8SLKs+UI8u5/JmiewBrqKCZQqEzHAoSJKjmOE/YGZHtO7kB
fVQbZb82jOLFWI+Oa6RUhp1SVx+MzPO/GAMQyAj8Z6101k4b2b3IVgA9z+RIxZjp
fXzEV+v3vQbOKrDL794kMiv5K6xCQIEzrTRb+Dqmm+0XD/3lUGsLNEjcVjfHqB3P
Lg4XoTajKagvT3cmtQH6tim3GXMYRRsv7CUvaRw+skNewOprstmkMxYlQhAdsoZO
jOTrtvMvPQSgd5mGEIltCWK/6KMC81J6gv/vYmR05fgLpqU5v0hQqyOzQw9SibS/
4FjtRW8hPuYt27GAY9sCYdSf5vtwCxinOr5yiGcQy+uOOPOIWV7gJBA3cDmzIVby
l/01NmkSzp6+e/6SHh2QLHk6qR7TDVKQUodTloI0Vc7nSas5MkvJvhi+/PViGFUU
cQmnRLZSdsNMJI/XCl4i9mJNnMaIR4ocZaRaDZwE6r6U7JVK4HIAYKDUUYZPRNAR
DPUWew3JYXLu9/rD4YiQNDQgcVacrNHoOdzLbNxZ+z0FJsMhr0DAqyJ0CnP+CUUJ
hyr4aXcAWr/pLYVuDc4JSDfTr9OxYIOj8zAmM1hunDePkz9mxbnVYj0/eVEpUU3Y
6Ip5JGBHa0+p4CPeNcEMXXUpuiTki9saJVkyV9bwzn2Jw7xW/FmmcFhW0LtKideZ
It8znTIu8xaxBVfgV5t8uAazBdMXjt1FMAyzZbHd4n0WGWf2/lFnArEOyfmFj/ER
o6qV2vSGDUXKCjVEjID3vefkftc62wl984Rvi8ydF3QU3s81zCJumHgImQ0OSIlS
y8LXyl+SBsViczg+Vrfh8lv+4al5q1mJj2mKn+w4/duLoJx80N9pN4eReuFaH4Uo
NhIXkxs0EVIFKRcaXcpXccYqziyVCGcyiEkUVWgHER9K000jtFxRw7p/UL9I41qT
+OqYCeu6RGS09VZDc3vwY7UeVG7ynp7uP0GtfQBzhreZb6DDlZZkLUYP++qM8Dbo
LEqaZfKV1PitotZFxmcAeJ6NDzh3SS/go7K6PnUIsDpRGP18QQJHF5+rKXkwe51H
WpFN+6cTy63p4ej77CTGMIb4Bmsgz3ANlkQ21v6C/1Dgt4kgo2dlqMbzs64eOgzY
3PZNxI1dAyS8UbtA7g/45o7int0nPnbumGc9Xj8wCAmaiJzDuP8mWGQL5+06VVf5
gXUdjc/NKiJFFuklNiGaXkOhZZfJB/fw3Gim8l81E2C7rVqSgeRKX7v6Os5kmGPt
lxaESY+U8INPmPzmPffLscNq5KHZmrUXCiO1N4UE79dEy91uhyzbVuGKhIQc47PF
g+aYc+GH6etYJW2ntGTlm+U5XZRq6k2dbM/hcFVUTg04YCThcGa7xJyg00HdFTNl
v0ygiuLLPnkICXGUeKRg9jNQzriHmD16FL21jeHOHmuxo0pJf5QpPNHsDC6YxJ0h
F8P7yE5vGpnCYsEboVE3xW+//RXtIJTsumQuT2I6IoX80fYRtQOsJrm/9z0rkLPL
5XG8VLwonMgIbuNptNS9WvUcmRCIdV5XXWKenMUlB2MoCakOqx/Pl/2AWfuludK6
/ZaNenMWja7VbkJQ8DB4eTWMmpPDG/7RK5JdBay6Wu3JukJ2qVKWSArmx6ebVTpJ
aKyoRZQH7xZJb2QTDSltHdTmazxnePM60QmXU7tI+8nAz3mjvrq4TQLVvN5Y3+Ag
8xeK2VQWbXdwzUKaWCfW9EYsiQ/a7F35tPU7C/AcjtmV1nWI6BJ6YL58lCA3h82a
G/u2yPJYGiltNo4QEKZEOpXdSQuZyb8cZbHT4jgssgMSSbmXH2wncM0eLA7iC2QL
PybCW2oZAy6D4/AmPvAkWFD2w31X45ML0Vqkpf2IE8Vd1fvnbUD0MgxVmPyCpcms
FGQCLgLLAtJIIDTQqn7ovGZSiSjZTiaK+lUVFWkVuYEDrAnmKMYGwFoZxGGilbtu
gQ+VdM2A3U8LB5mFYrkgycDwrtzoR62/PeqEwo8/7uZHh3UqoGvK0tCkOaPf3dOB
LHo3WUJM1iCdg1jEyqcXFkks+2mKHb8FmT5rFCZCx+zLnzXa/BVzPYr1UuWg+Tiu
dSGDMNhyxL4t0D0XDkBQnrwf23q6kOya4stuJ7SG9xoLI990CzeBdHbBDyRJkcAa
NswFilbLiXaWQ05vNtd8auVgn+5GDoRtyqMLs6Oc4o9RYYVCA6ZI0HZ/9HAyOPQ5
bD1TmnVZmNykZnu5sB0yWaLuAhiMuKoXcgiQX78dSNm+FIQPu5ELP+uVUR7ZQi70
Hz5CtQ4sazbyQ029+q1OaKXiryr/CTKHHUEuzXBvSMEWJsChe4D1ljNSF1M1CEcb
Zb1EgggXr790YbWwMpodAyANEBA5zLOilALbW2cfFsbnlGGZ2B4uzbo7vl0Jo3/e
P1KBjJiLmk1wIiQA4m6lOrC06wWTlLiSC5rFn1lYoSJ0u9SK4vytKRxbeaU/G4R2
NAcFxyLNQYcDl+eHUXNaoiyewxuUJUrJhfkWa2tr/56aIKK/yTjHbmvNwpuH243Y
XQ1gqgsgwsQOCsDkayMRRzm3l+63gg9z1ptw4bcFYXvNwGH2NP1EvF2Cp2+44G7M
HV4fzEYID8E30ntjVvjouE5T1l6sjSOYg7ZBMJ7X8Z+syMWSmUn5xNASn5NVAOpA
YIbhDjkkNdITHLmm1V974oezVq1okrDdIrag7yvkTYxPSsrU51wyDybNm71De+nJ
qfOU0KO/3OJWzhNsTxw3+3bcVOzNzTaQXcIVDvjQFZyD/Lqss9YHX1j/hy770vrw
Ymbx88WKvdTS3TMF8vZ+MgEpv+U7Be+sd07tSasEOsZZsMXgb94tMGHDhXDVKvP5
6dHOGv9dPPBpyZwV2cXh3Sl6qkQiiMb347jC4W1CG+MGxbB9TtJ1dCB6fP57Ll/L
LaHOQ+jukqty5bF8g8aQQ1CqXWiefyqa43zslDRSLN6sUliG1+G26C8RxQ8giOit
pgr0BMjPaJ6r/s5SPMVCyYz2V2KtcgRKZUce7WlZ/str6yE+i9LHVofCh8FJ4pE3
FVaI1RxkCg4Rt2g2eXrxfKoxU/Jjc8t29f4bcTWtnS+pLFJWvFNES5Nrkj/6qlzH
1FCFhJWftbfNRqOSovDZNX1bV6SgscZxQkpW/XidzH4m9A3KBjN5vfXsMu8SKX2j
cmgCLcaVR4q66xYFVI4y+Y0yRmtyA8VUTK8nNo9/t0qI7n4qJ2Na0A7Fr+4iKY5T
94EBMAqsr/WJRkGeTDn75TGNXxTbccDc+aFii0sRyZc6ZsV1vx3gCZSBaMC1IHiW
BmkjN5DzNvmTZIvWzx/vXTOYwA+8RotZ8ha912P5/0HoyIXlE55GZn8lN9ddsMIh
V8KaGN+BuWPUpMXe8u/YnoAZ2aLIaAxDwAWrW3E9w4sSu5O9WT1Xu/FI6XSX3OYz
X31h7LP5JjDFI3q83fbcxrZG0Ru0E9UIATTH487hqPxa58mamnbZ+8BssMJFBJr+
gMkZxf0Ol0d+VDxTpio9INNbPurCvVhZWT5p7T+0U5gX9r7iCa3R7Lv7jKJSCIyV
f19Sup3Mhbtr67pUWAqVe9DPech4XbozusFAQITZQ/OrNd7BfnYlCWUxwad7Ah1C
QjfY82L4x7SLbCGvSRD3JGHRT4EKPR6pSOKk2LYstEyPGCdmEPxvJ1DVXSq4gArf
OLfpplI7izzyXf8851NxmplUZW4FHV6klHDCCKdAlOh7qp0v7pQgosLfM6ahyghc
DCHJRwx0JIsTAdbdTdZeyO9ZUIw5go85pG6LvdXSXOIcay9EDDGvuuz+d/+f1pB1
Vwd9+DglI2JdSWyOlsSYPauLFfrggHLUBCmJFiFptpAB1gy0EheGLCatMHAl3XXe
OKi70jWxi1IcfMzTVRxAXuVSU27ljdEEWz4xFtZx36DQLwPRJkJLTFDx6xHIy2bf
+kdGMjgoxHjizbeYCxKXb3XnZI30+J+gJhmO/nqQtqoimrIn+xvKrnLmHP4lBryV
HlV+U4JwC3B4dSFGewQAbKX10G9ulWTIOdhs+X7NTarKgwwqqtHWPty+4/Y316Q0
mzVSi/1evRdrHT5MeLb9HTC3QdB1E3xy527oWJ3vCUSfRTdp44toFRM5FatP5rGd
YJS0DIqrHQjH02nMFDj42ZxMK18Pog8VKOgbN45w8bCPd+hyJyHCjvyOdUw4ueQT
QPjHGUChGvYvX/Fpuo4Jn+D4PX6XJLz+iOHcyQdr2MS/JAHRGIE3xZN+VJUkbenl
eyubpu0garSIUYS9RtYOfmz+DU9bVNfrh8LIEJQg3/qheOL6e+3tDYdApsEkcU4X
mw3+vPeGl8XIE73gUNypS8avpLSCUaS5Y2/T7qev08BCaKdYXBTQDUz5D2OrPg0J
4prdgkPok03ZRaPP0ocP3ga5WiIxKDLpvKpBqDirOCxn0KvLtQE6Dez7YIPaI/o/
mpra9LOgvrtonmskQk0FDLxEzkg3yAcx/+he+owtwdVRatgcK3DdbzXy/0ZpIuR7
DZLQJ9DTLtMP3j0nmnPFm/6cQonuX5sOIUCUFsfkiTv+GbfhK0XfxKAZ6CowJruJ
xYyLQB+/P0C+XtQa7/IaYNf7Ms6b5/bEdopBileEEDJWi3gPi/qgk7TWaOeTHPym
lxEjYyDXyTd54ct8rMeZVADdh+3TRMF79cb0IgO25id4VefRiR/9q90lhFV0pt2k
Uk+EQZyewH146toaplcMiqsALbuFad51RvI7l+8Kyd2Ncv6Z89Qz+FHT36tQlMz8
6d3OxhIXunxHDV+xCga7f1T50Vb+fDWwGFp7rvIClc/OeJCHtZTJ2fT2aGJVw0WK
EUIjGOomLWHvnpNgIs13DLZFJF2UUDDk87k1yfIsfhxP8GPrvfP+0v45TWLamqzo
D3AwRsnj9d7vSWeupMVCMwBV8SB9AiM1m6eDvZv9tCQeXCt5dqlwQ6OBqTek8v7O
0B5yKqgUZI2obx+kU8P3ighfeoMk+bXs0OZ5q7BNfksF73YlvDr5mvY6ch4DUHol
HQuy0RGzzXhNdaeNN3fauDgtSwKAbJbzVyvnNXdBbkV7cSB4WAHWy3ahhGjD/R4g
ATAn+JQOLc8w6Piai0VnDW0kpft3rgqVDmBC2dW40wSM+Sl2TrzhRPQG6ZK3nN2G
96TF6WBNSK2y1Nzk+orNDbXV6wkM6YjaeujmEwduFLvMSWZk2gy/aviD/cFsmQEC
6JR7+vfK0e8T1BEG4YkQfiOmzkm4LDLewvGATsl57YUM7yqbDjDAs3Wz3yLGa7/2
K8SQHGMilhE2hm8WTmsJfHHbeskHnri2WWKWXUcCpicyS8Yu1xu67mW4RKYJdQfL
CeklTBt/rSdTlpOAKY6IqFchVLr6Ju7iqFkICXjJyPH7KLVHeY512cuHtrKaH+Cw
/ijMV1+JE3j8Iehcql/CG8lAOl75pzJrV+M1/C/4zBpWLqH+ogg331fdfcz3Ch/F
MdJSzHZk8IbCLmLwuE/BPUtpeMH8J9rjPI3aUrnsqHC6gRh/lo87Pb7O+mgrYLfC
hgAW9WRKxQERXlAKTNKULKtVrQo4UMU5x25UHtSnB8uDe9hxH7+5q/Rj3X+pr6+T
RMQS84uNfTX60x770ZGx+Yy18h0FKAnFOSS1vopqAbyedTHONE7CU0vR0kU5oAH4
fgDyTVOpiFTHADAAFHxbITMvyyWCU/uRqrgWdckVuMLU075hd+cFWOOFaxoUeX2W
wOsQYlvCnsrWMO2BoyzIcUXdnkSdphKLlann1M/NM1nUp//M7hYORHSmPDX599ou
fhDlaZT7YrHpd82i+rQogEarH2rWewatRw+2D+d8zrmzQA/nTm9Tdn6Vmbhof1PQ
2e1BYNnAhkJeafprNHCvtNwFjoqgGYNEEWHZSF7BskvCyGtP03mMk+8tJwupmwlg
ztmUgua/7s6trXB4DcyIzNbTOgVKfYfC5ae5CHi5bCnKauWgQinKDzWmDyD8F6MZ
Du+qHPGJoSj+IYjJ3FlCzq24HLkPLIpAQIc7fykJc3d8o+SlDwan3T5ZFqc15gIo
tUItJ6zEhs3s8WQm90BZW+rBL8LNzIJYQHYQ+q4SV5KIju65esFwBsiaCgcpiIw5
fV4wAJPbqRoguxp0c+VGDZcxtkVRbpxjBj7zeIuNJPAwFd+dn8o0BakUbtgyvBZF
FQecXlAb7OrnWuokA7jzXFGePjyxp0e6qkjMZ5+i5BtZpo68RMvd3yxwo67/2zzS
F+kJNrLewCxXNI/SFxQ0Nvv8InMlW0wn6/MPMcqhU0ENqW0g9OOGz1gIe5sUYD9w
KO5oKW2YURReixMF7m5XwXikbx1MsFIhcJfeib5Ypq24Ch9QRg+SK4As4vNAtw7k
/jxRMlaJWw8NHirKoHVFFfCnOzizpZGVhh3qFeQjoASVAJ8CddXY3cmUFoKdLjjI
nG2TgbuPwMyOBgLM3qJ2ejFUjkRsMMJFeFPbLvRF+scjLqmytht+Ua/EOSwtUZro
uBPcQ9ZVTnizo1FhhHMpzNREAEtbK7CVXbOxfKkTP8S+Qw9Q25SFmwgLcCpt3SgV
la2owbwcC84GGlTs83Hl8bDLJjRHJeC0L17OQiRzKWF9gesU3pfr5xmFHi2yAAxU
ep+FoX3E/QmJh+cuSi7HWjTBFMumpvjmhzE3NjMRiV5EtEfGO1VnaPn9fWJ5Iui7
QqxexXZNIwK6rrCUNh+jjYiDC7EM2nLyii7rHfW0G5B06yEqpLzIg0n0DskWtFSb
Nq935AA57+m0EJopT9wXb5Dis91bw+wvnDLkiYKfr64w0XeVJsz19aYYH08E9sI+
uMZMELiDLJx+aeO3VHzK+K3yqsPWtUIbs9Tq//rxc6RbxaxTtVo8IOdOVrP6xZtu
HF4dLetSL4TJXsvqi/WnFd0WDxSN4ZerUksXYFl3YXeEU/UKlMXIslhxHt29iUaP
Si3OMHE7L3JBonb03Wg1yUX8era6QC1HapE31RB76u1QgGW3HZ9N9h4H7N5jWP/W
EnFfxbrfnr7goNrtjDadZj6m7M6zk294NrEiHN9+2V+nLVAzcsnQDEaOMZHY5byg
yzHKO621t3jhtDvzKgJ8PeKUwj8PrnLTpDt/WANGijyJzkhrfMgnEb0lxj2bkVYR
++6ElGTuAe1qjB23DY/nyano4krzQyBX9UEYcoKPQHpZC3kEzCRkk1l6wHtbsyj+
/i+0c5sOlN1C25LwKcP0iyBx4Ty5ulxhZVbjMewZoLkAXb5LVnqOjyHVkUKNxvWY
bRag8TODXYgsQ4QpcewAk/s+2EN/EdggORLW1guh5kjYUskW8RZZOYCoQf+0VBfx
4cC3ucsn9ixJ6GnCEN6UvaZ1PjsM6GOHKykrSHMrfan1qCr3uQJ9hGZQxknOiwg4
KQWqxxZHA1SV4Vu5B8QNKHxpc+6r/p5pg3kB3bOpZPpGQG7IXpwSAJ0VMZV5Xhf4
FAufxaeFxyrXL5iIp9TVcv79DwfauAO6zvjaXE7Ybnbij7Z/bvUsAVLcb87j+Ngq
JqUsJSaxn5HVrSKhoXvqk8IXa08P82VDBJ4GP79La5RiZYwXBwjFhlOQBDkl2yO8
78t5sMkfYBcsr3PkRh5Nw8pEbfvLSI/AA61ahOsgfnWzD2qq0xfKMjGrxuDiDG4T
gA/iNuSWk9AgE/oprzf//pTh4DrnlaI/DpHsFCtd8Yd5uZ5pdmbXPkX3ea+3EOE/
9YsAidr3ZzI76PMX7+ft9c11USjDgh2GYdi2SQvTh9eDOv5jlZ4j19pEabRM+pC1
Gmo2i7/c4T8b14ihNWhJ2vI0P3+QgC1HLdYnjPhFP0paEqq1BNTyYE6xvM953WxS
COHtoSpWe7pXu2nphhgqIwCZDD3XebpDdeTSTH7H5vLP8HITv1ZrRROfATcFfqQC
e+fQ+f2yE6kBYQrocLBsE+4PH9979DqNtJhD1yRQR0CIZwLJ/73oLvDp8acZoL9X
jBAavbYbMfWevDj5O2Ax24/vTxOdcn5F5uOzifZwhFatzUP1QIxtXfbkOkKN4uWH
9XEhzV56Af6Phr1q4Adak5s8I4wIk8pRs+adL+H9cN+RtShdze0MrvJOgF5mdZ7Z
1gcpRwJagSOEk0jhH7AnDpa2yx9zqB0jd0ESvk+1baNiKc/COdfPHc/SfQ+tK+0X
QqyHJBWJrXovkrEq6GD4JMjhR4YPthvrsyOczov3e3KONXSk627Tlvry2cGf4JN/
sxEBUtGMgFwG9FE/euuoAGP51UPFzRJRyBwLFXC3w584zUakkYa4IkXqKk6xIW3e
0QCbtudNG9vw9g75J20I6XvVEHibIU6t1IIpXN4BgZJQQHCWN7RUkYvkH8nrKu8q
qWRMcAwgM6eE4v5dU29mo8PuBTkmtHzx58chCtKcLDcQt18qVT5GAatBgqCYnzN3
clme2rMmZx0sxx9q53wWb1oIdUg65gJNx2X3bcE0IZlb/8ngd+gOAOkJi18Rw+nc
S9WC90LOZ1b9z5s7qEWEsFSBIisZ7Qp+VXU6uw8kvu80mPBRJw0LQyIj2MUtPwXu
AVa5AhUzL3CdQWaIGDKrYZIf1HxNJ3MQk/GMR4pYPrpa3msyCtqHk41p1P7dSCbV
qsiwDQNxdO5KDAILS0DEMvPOn9pBoXZw6pwWyctdO4FKiY4MVNnNZURAY0iYSf/7
q/7hw18pr6goCra5h73pfn8IzQbwoEUbiJhimju6hsYmeDJOiNgveSCLIShfGqcs
i7+pYLNMKEPptOrwph51biBHhmxbzYZKPg6yDQzbAUZ4bHZw780URNWkNye753g3
YUwMdnvfk7IXWdoBzkEAIKSoI2ZDfVHgamabCw8osTEJBOVoVXRLqqy3lmbMswaP
M84YyzHaWb3STGdIdcvaIVHBcF6BvDSNlsBhnQtqw9V1AmD/GbwRV5sExKRBkicw
HNV8ObDVu1JcEWzgxJHsFRYUsxuasnL6Jce+VkM6f3tVBIj6fD5/rv0rlorFs3sD
r1AvntaRt9DVW+jpjnEddu5o7SPdEE/Z0Sqm8k4ipFc61oNnLAtZmB59vHlRe23t
6iz3cxVasIHtZKyBP+Y0ggLjPvk3ZrvJQcuTMy+LYBctKTkgWnygv8I1zqPj9WW9
IWSW1F1ZK2ycXjRpjXPITyx0XDmUeSr0LOTb4z/fgEGCgr6pn9b5G2cH2Zh4G3iF
q68Izf9EpDNdhg4nmBkBwK9pFE9u2HNKp/NNJg8QQHEakOP1Iu8TdjZTb8Uu1uDQ
/T6oM5GRz07VJ5OwSxOFY51pEfQz8oH+ZqErXyW4djdDaV/LZEIySKG+CAU+BoAp
NwHyuJIW1ynbK5LiNjvMampiVqLPm7Qe1+zTEGq3b0fLXhI9JKohsNrxGQh8J/5i
gLYo5c9nMBb65k8wFisAdk+9Anp7ybzER1o8H3pIBdcYw1QQI7CpWQ+rfDqp72Xo
pPphKSYWnX9pFIdoDfWKcW6IGdRaG0NHULUgA38CAVn/HAlFZnRkDREq2u6xJMwy
344HORpDwZvXvfF/9T3WXI3NnSa9VlPOy55ZDb/b4gUAtJYNwk+7qCFYtTf2hGDW
14TImZzPjPhLEpzpqpzJ9jyLS1RidP6hHgPzfQ2tAZ7xDNh8se+v/QX4BTOk0RRw
Uk9cNBJMS6hlQCzPlqq5Omqg20NJXxPAdErhZiooZxiKbf5dbZRv/IdLXwNSKRdk
KKNapabdQE3QChPVI83UrvY3TlOqTL0niGfR3LHfwztuKdHytKiBUCD7XZwA7yhW
Ouz/OzP/pVtha1bjwpbmxdxfW3+Vuo7a97OaBro0gi3XUE57HaJ1aCbCuve8KxIQ
ksGUjuRekiL9U126xcB84uwS4626aY3pJKKjWNWNkZ0IdoUSMUnN7nSGAs0Fjd9S
dTrRxuaaLJwGGMDBjPZ0BEVaFBLcwQhDRGT33OL1cIRZI0pjU9N/X+dm+cPQsmJH
Ygy6TEN2trPNX4IbjBZF5sf0bqB7c+kbZ5DLHZ8v3oVLLEAtCqU8TSx4GUY1v+Wd
RTr2gC6dJFz+YrPMMRpBMz1HQZ/L1wwaSn9zjR8p/pJGCs1dCm+5BItqS/36uJGf
XbK3u8YYxjEmaHevQP6kbY365kdm8+HsygoXaIgkpc9C8VALCOqRkuJqkO3bqpTs
a3MW5jQe+gDkVpU2ZyfNyu4XJZ90DsY3vuyGsApNNUeJE7d3fM1Q4L5iaeCeMCcN
eh3c2rFp4V4O4xoyEyg+oCKo5YjiJcExDRKFoBexC9JgFT3OKhN/9oLccr449HTp
FB9T8TRtPy5Nov9chPDmjIpF28F+oYUD6YudBb8ccqalZvHA+35CxIJ9ObIQb6Kn
rAPWes+pVxCDUt40Cvzhj3VUB8M4yG7ObaaybzfcjM1oXUIvqk4hW0lUwjv37+0p
ZhpZpRwulIHekAez8FqMC4lBrCMUu4zpYh+zjZNpZvCvJSR0KL8EIey/Md/8M33N
6s/vL1NouwvB9fzSPBYkhJHYCbuOkhFagKJmhn6NM5ZZtbpkG2WxNulN4E1tJcIA
0PK2Yu+z/Blie7HwlofcxVKzBfGCGou9okmN7djEWC4lhKr9AWY+FePK6S6gxMDr
DUbiDJXr7KZew1bCKvSfulm6BtANmrylryGEPZrIeryGmNbLoIQr6dj8RrChZwM9
kGHadLKAeFUw2THDl0ShgtqQESyPGb9Juk34M003+hiPJnD9V15BnHiRtASgHrzG
zZhrikUt3Rf+lBxndGLLQbutqsetjPsPU7s55cEDAp3ulXXb3TUsEBbptWfzewPU
x9K9BNjiFJCBkYsMoEAMl1HNKHTWaNhHvUTq18zJhLePnNZp15txQ6IsAZN2I0x7
40fNKGV9bWk4RW4usR/NV510w5RBhKOeEe9sN6k3cHjriX2RlkAKqetvpQjKfedA
XFCYkLm3TuFZ+Zadjse8PHYlT1GDMgzJKixTRiiVvhE5QC9zeJZek7Vv7QFWyqGd
emC7FW0sNajGdkN8a3zocdUaxT+bF9ncshou+EsXGyXiEiSyrkZWTccZDqV3+ysQ
/qer9DStRJT7tEBbFHi++IgSRKoJ26kGmfsDLzOzK/sTDOc0DpYRaR76AiymDx4w
dkzvjVTAPkOZSA1kZ1WJqCElRuTq3AQFDkwmzFrYI2mRfMhzxYCyrG1Z4KLxL4P4
fdEaxcRNHSC4gfxiqErfWjtOOICpCtP7jrJvAj/lTkmiLJ6NU4cwfvT3v0yJd5+l
5prGrI2qV85O+hi1T3E7KC8JthqyZGQRvgOrrztN5CwBjDpGKooCyMtmPQpOFBjq
88c3R4crsaW6fAuPOQ4SPYIGKzjIkF7HlapqpNywERGaKh1twR7B8iN82SHTaXGP
nec/u8olPS9lySQnElxGUuFyuoYr3nbIw5SY+0JiAnaWzZiPEZQHlxIp6IYL7/BW
CY0Q8i8wJwfgd/Qa7M6ih+iIIO5EBzg6ZUk37yECguWS2ktYK+Vty2qp7ezENhtw
Xtf6Q+yJWvpeX0bFcGC7UuoIHlYlKh7Ki2KkJ/STThhce+V+8p21+BNhHyqNf2vl
l5GLmtVxrcL1Xc3dGeNcNXIwzEM4NCesfGtQHzr4TEG+2xdB75e2kQrh6Cs92zQ3
jr1Nv+5qMHx4p4lpUD57tWhLFHHZxbdJ3/EunoXQVtWfKtaCsezq0Lbr6+83YAPi
ziMqPoWtPaH5oxNqLdIJHtOs9uyzAx7INtaAZh0EkTBSWkzsPUAq8n4WegR2bRQK
jO9Z2i6TZLRSbAMW9lGvjonzaE6biWjgP4DyQ5osrBkw1gwsAITX97UQ3Il8wCjf
4Glpn0fzqaBzancxnu7uOIDqD7WuSyJerDYcLFepyTUkqUgSnBGzR+WZ1PRjQCNE
En7jj68ZlCPuX7D/m03h3YiGVxaRiBFxE9D0PojvWMGvqXrr8y8WdW0UMo9yEIT3
nXGGvosl6CGMFw79fkyxzewDNBnUG5f9zw8J5l+eSCAZevSMICIdcj7xQlzgOE3O
dEnNanG/Zm2xY2QdNRbFNQy+H4ywdWVwKPZz2L9W0AACcN5ndnpGA9aEtuHv3geM
EKqsQDG4u2cc5YC8Zq76kPaWwFOmDxe1nQ5JFEcpt81lKYV6wKjnPyNJL+Gw1E5d
p2F8VYuUhv4Kuc6qB2kyq3Ki4+biKJuLrwrZZiA5LZu7LM24S/2Rti015+15grMn
BKrP1phEBzc4g33vawKH47m6kgoRtXlK3JVYlnL6ZQSgGjtf9DsxiY8JY3oTxJzt
56z6tjKsvYtosst6AcbQJTraflQqdR6T4S2wNYUS7vv/eHtkdo/JjHVBCnT+mQp/
J2+1GhBWeyWXkwUUbkCCqy61BNUduCEp5FooMFu6BHBxn0F6185DfSwvAz8igjOm
Fyd7TiiJSGaco32YZ+Ec2uYkLXgQx16ZRemGFYabKxwUBy8FBHoQT1Hf1DxJvTr2
XZBrB+7UMrNgK8B/Jhg8BM1iQdEC9NefFGIxoFdpSCThltMXTQn+q9jShM6N0RcK
peJlJ6dCLLnaxMXXKhIyTTlabI/f82AW9koLndpHgsqHSXj5QwSAMjyLst8yRrmz
HEVTv7iMFfi0uTZpoUlNT6TiFl1Tct2b5uGt3gzcNa4KeFDJedBiy8BPOlVCkXH+
cIpKMyb3pUMMiCmzRCQm+bPkoKkK6QV78CK6nZaIKb7deZb7Ud4AAsb/53Yf/BXP
GYOrAHBCymhVYCbYhmJvpCzhFb++CtLymZsjyNH4KL146Fbuh9qbBYXwCFaqCjfF
ylw8LChRoNaNl7VQNhWcezuEP9trw7sSFHD9QVtW9NtmnJH2A+kQ2LXtdkXJF+V5
J38AOIWIh2Wb0zY9gDuci9Nly5mCe0jF3bNM7s4uQMgpn8drql3qdITdo9JayE07
8g0iFQN8gGwM6vnvKm9+8Gx5y5EJ+ju8LMIYsDIU4sw7liOuXW0kS6V4DT4rp4Q8
IhOmNfs0FGBE8hMXUna9kRG/Xa+zmVUnLByYGiSeLw0a9VAkPpy/f+HH7MhwSqoK
WlkrKUBhv6tLH9c2mGjZLLHvBs4boVVHylP4Rg4UrLwV0c5jGx8iPUSbpkeQTMvT
dKcvlJPn80oijegwFkeBN6dfc/WMSTs2qCovlnmkU+bmK6DaDpdotqgavQsWE795
+2C4F4rGadkuYVkZV1JbEL+bC338OthPgji3X+2gN3VSzERH7LAwia5QxzFmfRTl
KVkMhKttv+CGRIFIpjtBEfV5FJ+R4RjLoDepprppXfcJibRjJZccGX9wBKf3VUw2
zRgql7ZTsRqc/gcXyAFuiXcxO9WRs5B6PDeU48dejyvU+NtzK5atx5YT27A7VBgs
OTr0s4Hys/Q6F4S529qenqLlb+H/hW0hViV09whyqZRJqzXuX3aWJKiRdSIZoudH
7GiwyR3QJP9sAA08pTaZ86oV2Yk8Jxl8+LUvoS/Cfh7XAnLNIs1yMsIBtQLjRDLG
qJHgh9+do1JXCMGbrdU6Y74qYEY431KgsbNRJe8D8yBkalPfNfOVm7qVOgQwng29
RpT8m/QjkEdt84Fk8N5k80iHLvARbBUdfnGVoOXqdBMYJLjKl451GCn1T8lODIhV
+wKu3mqN4ugNfW0orZ4oN+TIHOB6DtUSrcFvLs4wWwjfIt+1XqKVGuGCPWQ5TLhY
7MLhUjJo0vOCbuwn+Dj+pRONAhIX3dkol2EgHUKpW+IAt4987KBfRaZB9kQiT0tn
b8xmVswDlOjl6NVQSWiClAO+yNCXoKUcraGoZ3PuaJhPeZe+B5cNGuLszDvDeFRF
wtiidWr/M5qXdU69TzssKfhUuLU+gSE5mMzBfOatFxiNBcPM7nOpt2uoCPUcVleT
BQUZuMb0XxySmOYOoyq3B1ta+mQKkLKe+GBDg+QdiSIL9ZnCdpx9+5JjoM+ilUoZ
TnW18/A98eATtbMPdS1kA9sJXckSHYXQX+JWneBlo+smkH3hIXBjZiiJFYbefQr9
Ve7QznJLac9v338+ShMPg7Jkt5IIR+TVOdPUOyhJyyytr7H563r33b9EZVHnyW7g
3IgHzIJ7Ct2d3DTaEPjCMBBgqoqBHRH4wSQoVXuPoHM/egZCxhIv3vqsYnwF+9nC
dWfh8hadDlzuR3illj5WNnvw+dbdg646eoD2Kgs1hCqieIbmZ1ccK6fhMVdMfXSj
2kGR3OSGy2sUu6SwW10lXldTFbH9WD90T+tGtqkUlz3XGm+KRQ4K2wz3yzOFD6Og
L6yKcwTXCMQkvlu5OpYV5mWflkdm1nIjJEI1GsdS3ZPi07sFqiB2UrXsbGN+XLgW
g4QOrRPtek6nyN6aNVdc0XJ/NY+otriLm/yxbim5y2d5LZYFVS94q6Zuu1E//Lzo
SB4UX229hf9sPpdQOvSpOMTkh7CkGMyIFs0Dr6ZUivz84INxJRVQPSywqeTt0vAs
D1xdc4WHf5K7eJXeJCNn5l/ysBujYp5eSIOhmDLkx/ADHBzkBUtJBj9BR6CsP8Od
9K9dRGkqFrGZV2MOupzGtQj8jA/qixT1P06NLG/3bUnEqMNeV40xM6itigDWBbvt
8KMoYD3fo3ziVIMWkDoxIi34h7ws0D8phHg8SfjHHiGks2DsfKxqx7E3AYcr0o+m
dTXQLaCEO79S5RsKQwwMzBhkKmRQSRuBbAFa4zGIzSLncUfUbOaMMn6/LJc1R2TY
2SyaU52s0iMx68z2c1HLeYXJ0q1nGPxWEYue6tJ50LdpC76U3DcbYY3ZZLgtFVk2
g4qMYoRObBJtZMGpqd717uY2uoJH0+eiV7NoeciD7ovIgGwzLZXCEU2XoS0hRcBn
LOay/XJFEo8fN4lFmfX6N0oKUwAyul+BCBNIpAAtuXN8ea0u8sER3zx0jLpkBh/I
WnIvY2Jj7dfzGcsTalYDgdUrN+x/nrji1HB3CoG+5Oafwd8QjQ8cOIVU+WKF1PCn
Aadbit4P1WMEFfgBUb4RiMJxklM7KuBTAyhnvyI+ZnFVJXkWz78g5BoKSE6HpaKt
LfdRDBxkyKahuG+mxZuHcIk94Ws5JDH7UeMTbpy35xga/LN45FdJhqaxaOSWCYEh
EvENjgXqpGwjvrP2Jl+aFOmp9gQTTrMfvAV4axvXwVYIzSP/d2/h0ppJxmqTHm8c
LcT2Ulnnszb8SK9bSJT/Xvgvf1vPBmhp9AsvVCOlbOTYhDqo/XS28t590iuOSyob
7aSbB404ZDleAeMS46hpPoNhcdYcZq7BzJIFnRKVj7ytR7c4QBPwnLa91uit/5Ca
kfr9GurZ7c7IwC9xHYh8/uJatJbOqxlgLWmWOttx7ZUGhk68jBW48si0DEYLjEX9
Ijkpx2AzVPncC2UltYzrYnIN2uE9TYIJzefc+8EFCsyU22snvAcPhSf/9NbxsiP+
3hT3/AQSEfyGFrTqoCkGKwLxV1+LSB2RrawBAcevy6CcU+a2XIiO97oybtIR6VNp
q672u8KlNKCs11uFIRFa1Jop/P4+OxEHx9xxHjWdyGUXrEnUiDlZ1xlXr9jkslMa
F+5cwqZWvfy+8Bn3OW0Dum2MTky10X977J17pDd7fbNtuiNovTQzpA0mmtHikBHV
SqzF4j3Ak/wybXzTi5J9mTtxWmjF098Pfu8gDJBmmKw/xE2dLuVxNPpYUrBuWygV
4czK/WgRfhd5WyW3HpENnnJqKplMfLyPTAHKr5ZPO1lFTkSoLRKYgPwK58rWj66k
kJ+gLJFrzw11dvJB5bGl54IrwiejNPJC+ophwN8XNfp083Cjbpl7UHtKSTd2H9vh
Nqcb8FEHBvJvJaD9vJLJkwtvBcRVYKOY7WkPQ0dLhoy92Av84CmnVLVu4K9rG00m
7oHVR8nPmZEWdSioYsq1J0UxZDBFLnb5cwlL2R9gpaBbJ7E6h3JB1LCKiisRj5eK
5HRs1HjYMh1EVXxLzAGfQtntbz4SN+gb7hZfx0tbqJXEeSuz6af+aod4IQkrq31y
5PrlKh9b8RnIWd7OgLyE70LnhtfjTwF3gV+Bp7vUsxfTceHqqBAzqP5BsPtS7tpm
Edo575iyKBTf4/HFyt3BEzaIZKSF4HaQRNRh6h9Lwmd/jTpYEEGy9f2hdgQUDsgc
53Jluc+FEgCQ6c5hzM3FlRjZglWhF5zzzK38Pr24pbwuzuTPPGokb47AAM/nwmVp
WyZTvn7xxb2oJApXXWyxVd+kh2EQdKyOO9PFaSMyL5msvfdINInFRm7hW+CA+dqZ
0WfJiLCs4SNeUZL6S8kNjUv+o96lWqAZhhIAg668XbeRSuqFAZyIx/lj1WfSpl8w
Yln/KHrL71zzwgMXxqHhsWaSUGd88gWAP3YsdFCxboK2Q4D5F4tWUr2sdLeOEuIc
WZnCiiKWphZUjAj+HbS82dyhN2qNbT9sCOHKMTnpoXl78qLOM9uGZh8N3VZAec6K
yzKf4sjNbniLkvu2LmSnOIEgWJQahnp7Jir6Babx33oewTfz+LEYehRCNnqI2MjW
FUHLf0aHfJiYs3BLcUwxLWwYaN00rb5sT2iZWP7Ximx/e8WQ05CdwdaaZC2+bMgz
TOCoKfGBA7xruqKoChPYACN45zIdfI0XWEIDLUsYwc1IVj9CylK6C8tDmIjAbw8q
1DRRP0OvqpstSbwxQbxPnUSqd3LoX7WX0dzPzTzMdejjYoJ5OTWrYpSWP5kQLTnU
59JxP4YNl3d0kMx0yxJX6Gu46rkB60NDG2w1Vn+sZd4n/CvLflHlBp7DoSiTzEDg
+tv4Br99kme9aZDzokaad6p0PqBY0OGHea3+FeIM5IQXJi1x/tiy25bGGAsQgPva
NwFRbwkAlqAKH9XJ50MhXZfgiGN39QrCksL+GDZym8GIWdP/tR1XaOHb3clCL4aj
ophdJV62uFOg1C+w43t+ieUrCs/+xS8Qi7YA5fEst687qTTJjGj88S5+adz3h5wi
41yP5U8yPQekJSdIO+oDHDczw3R2V20vb5zWnafh1ihMR+vi9HB2ewIGF6Xq79mD
7+BVQ7eJ2EVyuzRDOqio0uCCYjl8kbyibOE0QCB02tQ2ELBwjGbCUAIE061X2m02
7XctH5NkzO5trpz9IxOA5cbwCw/2/hn+LiWel2LR2owv/fY+OOPB6CrZVaayzdtx
ptrl6TTR9Px1oGTcUxcuZgfrzK7x2RqxnfD5luPQyvMCCEne8BVpc9TFJEhnbT1C
FmxYHDfSxrPHQnxRzPVxpOedP9KW5iOBBHMXIze2reYj8eC5u2rv50rrKoFLfnjD
gP3bBrTO0E68WeDUy+Enu0QVk71BkdmIG4C/wLsR8YkT2tnWJFpxgSuyDTNh8fyv
p5Nt/IZlUklvZzBNg6PlgNpG5LYN/+TZxdbBTn6CwAOxGCMMLbW57dl5Eh7sednD
KM+q2/qFeqy5eUWUhyelZkAb2+TIjL+hz2WfwzhhHynnr3CBjxDoWZKxWcS3MdX/
ffTFrm2r4I9cBoiuWbhialriEps35mjlQ1WpeJXKcmKe0l8AqD8A6DkwAtI+vMyK
QNrheH5Oe1Ku0v3WQ9AK+TJ6e8hhgESh+nOVikbamSP5r2sfHJYjfSunYcHZibep
3KGZeM2fwX0uXd8iZSAzZN0KsRIRn5VscpEjS5N1a2JxaqnltXYXBCtAbrocscdC
UU4QPPRPKHJx/RgzcS394F+LU050vHSGbOJ0aEFhn2PzIl9sCO+oabkW+jwHt4V2
w+9Au3L9Kz7eVKc5gM16K0e2KRwLOCiJ1zbdJSMPbMSiR/M8tzlliKJADv3ALFrV
PkXptKSeAz1Ed4PIkRl44toUIu3QXR1TYpr/6W7Jvv5Qls7MIVDlw6j3Xe+ONfEo
ZLIBhYt40AnE34e7EIKUOWz+6+fPQSD+MBlJeU9uGuXm59C89WOQRJKfMM1G53jP
sIYCkSm8fFGDQruUtQ6NEQyvlDv9pK4jXRoKf98DNLlUdC4Xpuf5Qv2f00Q8QhC3
mu1hawShv1ScR75y55KFB5/gEDJ6ENUCgId7etR+32JGeLBofeExbywCqbatzSPG
mXKk0Wd15pXTHD5Dsirp5RWxD9soM1yxmmdnKHpqrcKx2oJgCUy3eKMzQVM9fsu4
wu2pkO0KwXl2Zaeip7rtQI15PQaGCtwhQV0j6L2u9Yxz/ps8DjW3v4varBn96uDK
ATgiDcZaS0pDg4vuc3zxhjV/oS+QZ0X8vgiWVaZ7J0XT7JUEdiMxKTE10w3Rwu2d
eUIvJL2qtIYG/p6cJ8cCOh+T/04dOqtAiNpPG8iVTNH29nboeG33aAsihd/wWn3Q
/ELtdLUrWO1daMSUBgzq+jz/e6YCvGMCNNxSugv6aip03gaytix/63bpuhK1m/n0
+27sotQMdjDp3fDz6l+X7yybNH7Q40EzBTZi2yWhuHl/KNjkzBB2ORN5CRf5bI2K
pJkxKyMUC0Z3ezPshmlnckIre4/ARO0QPph69VwS0WcJ0VaN5lKQcmvaLAJR7hUn
RfMU0CGOSGf+glY+3m4rOx2bwFGN8i9WtFGSuGdTahqagm+6xUlPa4roAk08G6P0
e/0xK7nLI+ll+4eUihtFb8A1hQufa2m084HmWHqXYU775j+DW1afxe+4l9JX0ZAL
E0Im4FiZ9iOMQBnq1MSZnGxzOisb51SzBreIjTzDdv0KrGj0vnuhyd+0ZjzWrZCz
c0tQHIoMCBx1dppgg3zT4o0cHkPzqebD9OVptivKIwZ678SGR6zDYpG2cyAJkBD/
VfPL4CAl4vRNI/ctFtbEkfhAZ5uZq79ObeMRWnompy1oE2FvCrteyFdbdO7lzyiO
vb+UYd+mtQbrk6I+YXuN1vw7XBvUU/7XXE0xdPsCztb0HJ/ZbKNnyTwn7xtkTHRp
y6pZA1jWY4+FfjO4lOIB/nOV/yni5osUIzTJoldF4ic7XBIrgK8gujOSG95qGWcq
TA/X7wlvtxmlU9KZf5q8vc96E1EsoJ0/JeGBDopNpKsqPcAu8KHAoRfx/DPUi0gT
YRYcs6r1WJw2kc2GmANdV+h3OBztDinZOB/uestyZhBiN65/lpeuE3+oWgY6KgZe
nrGT//ImzQOjk/VpS7ORMe1dczivMeI+G0qVrbCilmiGmPytUR8CxQCc20q/KDIK
UQB7+XOKClaK05vl1isBcAhs0phjuoTzkzC6+WNIPM9rRPpMC6uSRrb+c8uAfDIz
VcJoFyx1yarUZOpOwIV6I1O2JA15KjjeH7SfB+Ae+H7b6a42sIY5eccGMa7MUL7I
FKSRG9xc89MsH2uPvS8L1NfaaNeaLxkmKUgT8wojSckaLOlCEysoVgGK585v5Jm+
DFNAwRWyZjcBcExilF1oLbiyYP+9toUuZjQ4toqT9tKmVUXvn5FXNu1/egNTb2zT
fK6ncLMZ6bKjdOTZujjEsBz5UFlNVeZOfr2WYnXqYFxgmkhBRyNqxVBCYpzPEjIX
OAKo+dtvniBP1zIgJ1TSUHksTSNhkdho92q7VnTD9Zxs5u8MXy9B/XTRTfKpJ1jO
NaOcXGtmx/3PLpMA3rsM5E20QMCtHR857qb4ifPNeH36/4WsQARY9zAcm6bkMTO7
Rk19kozq1XNNiBmPH11MZ32iR5nY9UoLKB7yBvakVXMuQ5urZI1iWE5UBFT6MEDp
WMPYSJoq3AiTWnTxMDVCNOOpt50K7mQlPE9wx54YRQlT3w6K5IXCqE9TfoVOxe84
prYtzE+mKHkT7vjapeHa1+j0cMSS7jnW0t0qgSikMyd6a/VtBchhAlv+mV76nn9K
dKXYYa5KeERkBKg5hwh+qAZc4UCMTI50m2fTNGXdc0cpcprySUsZ4rlMMhFOIqqY
RSFqiEweNvWox46mV3wisWE5H45wrZn7LtFNjkpljUqNlcAtzmyel/4lCbgV0NUb
JV2CYOOPlfWLJpS/6d7oRffPtvxTPudR1NS8cYt8rLqNzsXJ5PLYLiAhWVaD2Lke
aAiNMkHclydi7G/ZWsNYikfImj4GOGVaSty4XDem3F1N3SUavjTGeT4zCQQTjTJT
QoXKKkFG1MBN9IirM454GEBUCdMPGXumQzqS5ggO4lvEmt4rh2nN0GVWjZCo/BjE
isppoSFTUiwuVT3MXhHEcSbJ/DJEi56GyKeXWsAtYQ5DAe31IAT6oh67UgSo9UIj
7J8hlLqt4k/hZEZl0pRH6jXvQyYFKuab1cPBWD/TSiRMVn2ZNpidIgB+Ge9/05Lv
12VWjom/b1syEVzmxbFsng7I6GWYcgwynAk70dELWFrBOVElZk1aq01Mje7Qiyxb
DS0q/G1UYM5Ky4vq7zKMOlnyMP/M+WyMfjCnZNZXW+lVLvtccQ6Zk6lXsUMUqig4
NRrhZYmQT+XyIYMIZqI9F4cV6FNBSDKKjl3F3gC1RQmyeTXo/67b5TCb/vizbLIL
cfoXOrkok0sWQ4WNboFy/sxbnnRUoHeXu95xqvKRJkolV2E2Mk47mNr6WQ1+2ITm
i0+dck7yrrihAKMTp1U52Yx4H1P0GO48IoWyn0TTLKZbi+ug0DUQUubcPzL8cdNZ
KDT+7ibJFhWZayfVDg/nXAyHZTgAg45CJHs430jxXW+cOJtT8Km8dtB5jAPKTaCo
gXFDnEgzRZuWLKEg6pemayHArHl9YtT/4OiBHk1/iMNs1pay2XGq4jYvd4p+6ylD
lTLSSI+vJYWuc+wwjYl3mx9mX0VS0J1idXCnWKDSntU2qWcWDXVtQeQBk5437ntS
wJdPlreQld2aoYeRqJHQEWc2AGtOJm34SnlcrNIOmFakItN5RX+3kavCoWC59WPe
qlXaVA5moGqCfgLOVxQueJAbBKXoVzAgl+paFpnTivpWMpXqWgRhxvBG/tCDLAER
9Mu1fc23EYOjZssRUxZ8cXKszTzI7oUvtmDFBO+1RE+hkZqJpauFnXjEob+0tEo7
WLfeqoAKKocHlnyzB8o6qgtXXK8z3PkzhiW2W8Te67uTP9yXPtYFH+0y5yCXI03l
POdDle20WGyhjWoZFv9T+1ZN6i//at0Fuhb4PCbO+v6sl1EMufImaVIDcnKzevSO
Gj45lP61I1Lk0FOj2TT+qz7zap0mVpYlqHJdUrJjxRVXKvZUy8XQxN9bL5AQeVCi
F1nJDt/i2GDmQ1kOOoQ4AjDG+V2BSq4JZJyb1jmIUmRbbZiG17OtX4RqxCKrS9vy
d2h/wGf3Kf9m70VRYFxv55wlAh1LixvULY0FiOMOJ2tDaJSgDlBR5BW2bDqzPBYF
n1w3sX5c+7KHb2A/efeDzasKDspjoK1/r75sM0f5PZQMhLJe0S0pHDivdNHT0u1e
k0LGTTYU6TISAMYCpHnoil5Fo3UfmU8+zVFZi5r25jwcT7VRvnuskCkw526DPJpg
0ZAb57WOi2jIdk2PJ7enGLztOza36i3dE6DmM7W0CPTyhqw/ALChQAiAhpopUyfY
I8qGtd1B9CFhMl6hevh7MkAzZdMBKKSiDmZAmC0cv5TawuSLYcGsw8VaL5sVPagf
qqxTcg5jGQcVzon2MXzCuAuGeT8K+N/q3mNi9XIYGupoPHw1VOBGHdX7O3wE3afT
mu07vignjE4+C1w3gOvhFEVm4+IZtIbF8oIcI5NqatdTi6Mw03aZ+JMcYOJKeYe3
KR9LyV2RJv5anqBguw6TnSoszR40u6MO1tdP+eKMREfJZ9nG6FDEYsURmiU6RZP+
QhRNCjxpfGkTZyodhXRmSk9m/SEqnZkPH5i4UtR9PBHKMce7f8AejksrHwMbHgvo
T9UGaLFeUXUVuBcLaB/1TwAKresdGsyeMIagA048d/pXsUFmBto44ckN2qvCt2u0
/ISfomFX4S/ORlsuYfIe47XrQaU0/KcvHZHjX6XX1j1ApluW6H1LUZEMcvX0SYpu
1eyklFrb6aYaqUQVNLoOyXHOqpknvymXCB3xpB5MZGzNrp4R+qlkTAj0CgrMTxIH
Ih1TONawrz6JWSDFaVlJNhqkfl1L6H99Z2EbxvBjxMYi36KaRG5ZMeJeBfIF5geq
wVJ7paehQ/3Ku4y7trTy3atPQBJlxeHynRs4/Cu0+xu1UBXEYbTkZ6yPp049+2hi
K1KP61cruwsrpMXgXSGa6H1MX+NTQDiSCp77KjZODjzLzOh7F18EYPstgAheWjxZ
WS8gjHX7TNqT23hfEi3GMNgoYwGt4GIuVSLk7qT6wlfW/bn0djXmqMOkdBu6S4ZW
L04pUmM3/IBXiX6gh+f5c1CTdyA3Dnpgynz9xBdbTObyX1bqQzbcJP2iJEuF+24H
IvTKtP1RUeQBSDDcq6INhhHBpQuIxhpph/WfMq2iaTD6/GPD5F90Y+Y53xOiKjRt
F9T8gDuhB9vrEKKJHKO1CXLLa4LpZQTCSjzJPFEB9W2/IsDA+L5Sfn2Sf8UK7GL3
huMtX9u7XmNAbBJL37RgU7U2eyRkOJwWZYigbH2MAjcKgP5KbaHpqEJhFwvplznA
5ghvJkO1+Jg0NNXaL5eQHGlVcrrDHfjRttMrVLx/UtFbJwjpFABziVuXO49qPi7f
kmnwLMNnE7CEZmodwSRZwYMPK2rWz29oSIlCEkd+4itrmS1uKJHBTeyMtx0PFD5A
JSOteJL68YGfvpwdR0B4D9gpZwSglflqOWM1foeoSHaOLDY/wq45uhXhd8eLi10i
yvO/2LK+Kgvd4ZiuzJRER70jE08r40xCuhIfV+4EPLXdC2Bz5fXsGsjrGCKeKcVo
y/60e1Ph6/j8KDWOn88EKxal6xtjeccG6OVOQqEFd8/AFDtkv/a3jz0GxAjOIHKc
eLzSx8hFUhXXvKMiXWmgiKW1pfEDcjNV6OI8BU1UwuGOr1x9BrvAXrkXXq0ZJjN2
qTcJa3TfV8GZFTpQg6hxIkBBR1bIg8JYdE5iyvB0A1bBClUoyG8ltC/5LV5JK4r5
WEV2js2c74qqgqEKKJ0xFMZp/LG69Y0eKj2eTD/+pS25v+9COYiMXdFmVMdeHX5z
PF3K7TqrruiXbwwD56QMZ5NW4cDUmS7IMQsYfBDPVmj8ZP2LYGapFNUFWFql7+PB
JIBYYaHSsMq+BRws7+7VC9Gk/quWcoGjpqWffPmHfDljZ5h/EwpTwzXRhLdzZgNX
ghXl1IqeJwAGt/gf8uAUnbJUjX6HmM3M2WEkkSJRkH0LsUowsOwtxJLR4JwlgUcW
8tm2ucbYAgNznbNX03+T7Bm0ykyFhnmJSQH5FSY43GVyDiHjs37gjwxPWCiy5i6I
hBUH5oTVJK2qy92YMJ0qzXdIk3Ezm7MDwDZfJfuTWGWFY70y9WiYHiQtoLvExJMc
hlGZbU/AzcdCohTBXv6Fqel7Se8WHnWzj2ia7u7F3B1F9fjh/mME6yrQNl9qT7MI
LM/M+bKmP8HmAtWTAgtwMNdI5LyBHCepKK+YO9F88cW+lgb6os+bVx5G8ZKpleHa
ymORAhS9m4Q+xY7Mu96/bmXjBkwBwtO5GJnM1QtfR5sVEp9tnDNAYySh+k/7gDdE
DrP9QUTvBhsSFIDS7wTrmlXuz5QqlKot6yTdlW+QOze351rVfMdh2HTjlDFVZuQ4
jFuwXmg89dFO9y5oNe+jp+8YHLdP/q/f0xFZsLS/5hA3OSz+742AFADdiqCNAC7i
aHCm9FU1CCmPk7eWW09/nJPdeg67ffGARthtpGgwTxhXfw6RUCN/vy+GZM07DDBh
O5SOLnhcuCj4RHf+9zxVNeoOYZODC1HNvSHE9eQSmgJQfEhUhrZqMRS9y4D4BhIq
lJvdDZx/hnuH94S9jeUMP2vtgYDMQfHYsrLx3fYTvIHbPqX0WXzeoTVPsz7pHp6b
BZcNxPgFAyBN31FINuIV97OaOHbJvinRiXo9NKwvChhvYflSYQXYevReLms8hbYK
ROqKKLJ/6ZKlkPAQhiI3xSyl7ddjoELGFtb1J9lwtsRBslok+vBgo6lg/kezy6Lr
zyzHYfMeUcz1GaXxyx3TL9VmBmI5elx13glQ2PsdCPVnKatIBulUSON4u6PAKuOp
yLTKK+hD2MtPD8CpWe8KkSLBhh+2xnItq/pJ0dMJ8LY+aLNw1zURMn9/oTp5NQDK
/wCkk+LbPa9vB6PEZ0VAsyvYdXxiArC0oQ9G7s42+107L5DI2IjbnN/opmbRHVqJ
enGVBFwBrMzUomXF2Ck2KpmSB1vjOsgTqODluUbvpAa/gWvyZt0Maey31Vynbocp
USa+h25wNOn9MyXcMx/NcvS/zQrj96mDq5fJuoTyuRbj68VWKUnC/H76eJZG8DEW
IHko/bUIvvNUAX2HeXDao67VtVc+7bEZsFfI6Ugz9EuzUr5a03Zt148M0UWzBBxl
pJggbdP3u6oCjjxlAyh4HxmjbR7sZy0ZA24ZgpCuEK3RWahAOTrPwU5ZwNY68X23
4LmnUy4kvtbiubIItRA5Ex16oWfL8VVEzvLHq0sz0lWweksDqIizo5vtsezCGB2p
yD3EkbahNWynK3Tp6VPk2M1zfoxwY5pOh5uXMmdJgdIbP4tuJUhOlEbNeRSz8BUt
idFWOkAaoYfhbPUjQTxBUYz4vZsEcmry8m8j9/JYAsGISScrgLcJpeo19ixU6vKS
gTvZeDMB5Qh4WG3HPUzJ/Px9Ov2gM2eydlG3C/xsB4xdHLJV0HbfZIzgkP22KbO3
AeQchwTa+YC0DPM0RBHTz/RvEUIeLfuWPuBDRLjOpoeVfcGdm3x2FPsqneluMfSF
ZD+rLmU5weQG+W6E1RP+FuTkb4Zc1TiiLfBaG/mrOKOsZs4iYUHmQZlQye5qiVsO
KLhyJ285AL3LzRztAEt+gJNeuRCI7pLfHZ8w+YAYR7RtbubJQrbLgrGQPUR/fQVo
LJYlopm+DzISddVAZbu4EWD7VUHDwODEo0JC/qm9pq2bqOo/89IYlV0wUsZ34pEP
ZbEug9dvrkzkstPpKqxFWzNkYywJLfxp4N0wD3iIfFyyA5ZYnnY03CNvXq8LBOtK
2ihs1nG4DIl5hLtMCFYeeZ/rdkoGjM7ZZsvRSIXMUy7sEBPigkLw8EwM5KaujK44
0ccVKDcEDumx3hq9DgsfYsW/VbPlrZAtHuSec7+8JpTRavpNfvD4v7767xKDe4QZ
XRDvE7I0u7/JzAnTVAy+OYyX2HaSbriXn44n/k7oRNOAdZmtiRvRiE+7FvdYdEIk
fnHigZfkxp78VNH07PsmsbcmLi+dKNpSeoKl0xuRw6MU07LttZeLuYNPthuftcov
6qqUbOSl9tQ3xS7zh00Id/i9aiEI+4ooJGkKgNdLAa3DcAsPWuW5iWsze/d/KNSK
qqYk9FfTAgXWo2pf/Jm5eRDYowgQONLQsXwRs3E+RynSvV9lt8CNNQhaquQKxBn2
PURBA3o4ioDSBCgVwscImI1/Tsa0JcXO6X4CmkN1ZyJprTVnMCGynwGM4ndBf/vw
32YI5vmJI3OWjePYNsG2kwDafY2xRuvOPp/j74OSrmS12xT/MKJ5MiA3C/wyXAe6
mIO88BcuNYG3WakFwSuhsry/HaTy6dOApzNLZnlaUOBLkKvWwlmY/rWbLxPATdcm
ptcskwBkBwdAjRl9Y2p5J4FCRU81+Bw5bJhWG6HXU/r/DUpUrbtHL3wr7cO/8off
yJAaLC3ddLroYB3YIL7neUpJ6h710nHj8YfLgD0ROLUy5ThqyGiPRoQXqmz/i+1S
angsBcPGuz6BiW3Ijk24WMrhHMGiBqsAyyc+sUjfkA3dsfi+WCoaa1AFhRa3JFMS
7dZDBex9z86sLs9dpU2HFw9/EK1rGdqxV+4q5ul8i+lb1hFQ14yeHpLcFWFhAnbv
KIzLs8IZPJ+V24rIufmj6qSUn8XMmyfxSUz3MkDUT5HdQ7WZQ9R7f53bdaVaZceQ
Kkxg7CD+urMOquaScyjs3XI6WS27xee1RUDV/xDf3wgJ5ahhIZ5zKkDDYcBf4rK3
zCCyReyh0LpG5h7mdZ7sbFozpwgJxvvnobrDb90rxmdCkcDCfuVfTD4bbEwOMKsY
whfn/YO5vqQC8O7XqhnPYhW0PT8yPC4NsTdbHcyHweUr5bZpwJflmnDe+sEurT5o
or9kVnbXiJL/QU46hBo5diKpaACnRgVzF/lcH6cmD/l1UNC/QHDIwQnbFgjKdFU9
5TXZH2ac2DEY1PappAuJ8/nd7txczlZ+6A31JMTE9geqdQ7VOFSdqpinhLaR7ew6
r9z4cUUGBpHaUeeTyJ0ft5WB2Lf41g+AlVNt2gBZMd3j57g/8Kwkt/H2dvM1EV08
u5urulBVW7cxsv1mL1/c6TOZ2l7yaBbIvsqYGDTg53gVCg32ZqDNOXG9WOkVlOeq
1J0FWZmpgW6FMvsthGZyNTJhBuf/bGG5o3plNVIG4Qc0D79M6DE/cEbpRafW08s1
XyZInPtKUF3klv4Ayl8Ehzynhi2sPNXMSeqhbgwQkmxweZ4DCYLiy+f9QmF+DYBi
sK/m0kxd7pmkLulGul3UIUTjMK6V/WCrZuBAB9YHr9FKiL8Orkost32Fh0gT+Fyy
y/WiBWIqRPskQWe49CY50k8Dp9/EF4bwxnG/5JFm80LwwX7C5HOC0U5KCtFkSnBG
NxBX8vAIa+Svxo/BA+mRdSRN4A6BSd4vthlDdgBVvn/NIBBo5g2dggZU7nZHqeaX
IBbQCPx579d9PWPX2PIPCoNA2fmfLTQWqIrISzx69WVq6vE8TUnIPBuWBeI+Vxcx
DMTimE/s6Oi+2vqePmkFDzQmKUAzwumD7IfhbwDHj3ygN8sw9JvtDVx7hfX1tBN3
idAFbkX6SbZ3mm5AakbTDHO/GuuND8chbqSxG7W+WRJZwYV+WOuLjgPm+NwSDmQe
Qo6Be05/h72V/hwi89+6Ld9GCIIyHC7L+re6ITGdcz6S7xjQQ0VKkFJG65jV/H9W
gy5E0mnEbyqQQTCW2lLVU4zmvZwjleSNIXjU7oScNtCVRj7iScOm6wcWQ47lZC0N
xmytUwtGlj90GbwcXlAARbfsUd6UwTHR2yELYfOfAQZfe85RL10QpB5DvwmxCyYi
adwtlH+6GxsrrAVsVBpb3TjnZXbWIb3V1X8Jg4i7OvkTF6OrKF2ZwUHVnQBDkKlD
t8kNZaizbKcRqkjVDBH13RifsfGdsgaEu/iuUrWxpB0u+eP0fajEuCWYFfIZ0pge
uFx+ne8ZWv4138o5ipgvlAPXrql97BOEofWynnyAc9ZBzabS6a0tXulEsJ7fu5/F
aZlW3vss71BI+ezk+38o5l/4wFObPUx+zeRwD+gpgbUSENYhRXhfgw+9RmmtoHm5
p2Qv2PtchaIGc3LMW2IUesCxgHu1QxNyUmuKs5IIvExlc9JkWNTqz/6ddFTBZnEk
7LHZEBN2nwxThVAGcfK3zaMQtWUcMtfYDz3ZiPk+8gCp2qIXwd3M2j89CcYhGIJ0
1tyCETG82T1Ag2R+URPdpiF8YccM6IlImTeiSSAiPuf3dPanB4nZCgrZz4p17Qks
V1bhc5sWNwooHE8ukleGvyXox6wRmx3OH0q8M9VRcnw3lClcC7xo1Qo1lk5YwN0C
ZglAP8BJPn2SaxaZuBdboORmKt6r9W1RHZqUu7pHflXVvkRVgxQryWdBrd+18BPh
W/H1X9sdDHbgGoxCA/unhjvU3ArtWyFv9DPXTLAUiGkYAlerHsbYh7TC6gvt5vHu
Q0OklR4Qdp4z9271OOO028f6vYRbGR9lQB4R0jAa6Yek9kWPbYLgw4amvSM76Bzf
ynxW8OJWHVdLGUfVOLyTQJiRx4k+vrw0D6qewitSUECPNvKQNBQcLivNAvjUp4IR
P/BUQmLia459Tu3P8kzp5oHEJ/ncjRv7ck0sktJMbK9Qk1fl2P6rJ7FQ25kiOQS2
9AO9jU6IEMQamhLE1BZGOqc4OBAQSYttlgQqvteeuz/sTjtaoW6qRli+blJZewIR
DPWyXxB/pBD8da7gRq/cSSPsTdIOCsAyvhdlFwkO9lHTeWBfgZbIW0J0SA3NOUjZ
96bV7lpn0w/D9igHddlsv5x7hSE1Jv2eGXoehxtPsHgdjYSVZTLIHbrey/R7mcjr
pYeL6V6apTw6NkP3be8FSihHb8NevyeaxJE1CWacOfdwUabQ1b+rFIrZGsxXFJbU
tohqCHJoZocvp/eOrPhs4/hKBe5hqZtbQxNFjItWBzJWDnO+OE/j832RY/18yFqx
RlGEx1Yem0NsD/JheDYwoGPIkFsh23bNVl0k19e5v1l+DMLnONW/k4XzqM/rPq7d
pEvq21uajiMF3d8hlNP+kuKJ1FPUWncql6AkS8x+2rb+K4VF1JmuZQLsc4FvmxO5
CiKRqEUCD9uuaO0dxPL5KmB0cWJ6NfOASmAwo+MqkI9Nx7XeylYWp/yMJ+0CPcQ5
j5+ODA9YIpu360x2JSbHdu3kxBjeSv9R+qNI9hT657nMWNHtqUr/gq5T3O2FMpk6
mmxh5vUF5OQx7PioViw4CJbl6dK5cMrobHRZMPET1Gu4rmsYvoHTmElSctM/D+nw
QO5cGP6MxQXGJ3NXToGHs9E1MFGOsrfxhGSH/OgQDfVJ/D8B+2Q13jQOkynxdop/
Svc3lp1XzflIf0yU9FnE49jIJfd+pxxrWqAXW2wex0geVlgr19m880kdlrem/sJu
3gbqrg9SoEJ34iIDh9NCrtKDmrG+H/MND+16+Z6EH+iSnK8rLqDLK1wm8F/WmAc5
NNG0F01lWBYnGncHx/pXozIngC1xkMBB0mNL0fhPeRleOy/H8nfj4VMG5if2+wdb
VQouqnAECoKwiqJg370+eaAkNUUrYoQ1eR6TQPYHAFkCGjIxQMh3QIUIcK4BeU3Y
4zIYDAhmm/LIy6h+InP8a+q53UlUgwYRNcrkzASaTxPInNJLo1Sj5zwEQFp41vrp
Z3Hnj6+wxyfeOJMHOk3LSMqG0E3DMKhKHx3Pfnfm9qLnaZTrRv0w6MJMv8BE9zI5
QyjOLSY4Nmol3KDcE94kiEYlAHlTPz4hcDU1aNc+JpWIkFU7CP/hG2kPqkhEzah+
kB67poaWB/myVnw9nhxuBCRRWTTVkph5/nouZwJ0C8F/rjY2uec5X+7d72KhtXNr
/YbPj/Ep6ppfHBLguaa0EDlwFQt1CC9eUvzzwsGQlnfbPZvhEuRb0gR9oq1ReMin
PljnebWFrGIOG6TA/hOvS9N5UibBwYEcYBOX8I9OIkGyhZo7RXseeH345f7AIRxQ
IJPO57gb7M2HEU2WXAzujwAOzFTXwHBNYY0dwdT0knPTJMDQszcVa7AyF3SOBj4I
GXxjYzKNyvKLoIOoR9V7NJi47lnNIdpYGUU9C+zzj1DgFNFprTqnaD7TeeBG7yuw
ergSBnauocklrnFXVoFDl8+PLk0izik89K3DzGiutaLRbr6hjX8QUQr38e9bTVWO
ExjW6ayT5NVs5awstVfu0brUA4JF9iJPQGoBBDzPlvtUMDVS76TZ4dGTiPirbLV/
6IQqN/25Lfnbi1Nqjp7z9ahE3udHlY9oyZxyJY8N9SOz6wDfXH7lwhCfJEXOJjYA
K1P6tRhZscSy7dNVYS9s+o1s9KWLUD/dAZ7sBXsxAa82HCoFCxLY3O6iBX4HVvrw
qYSVZNiKqGpSa4aWLzaJowvmMl/Pe7mmfdnBgDRcbhW3AQIGHWuP8i1EPBP8L/OT
5CFWUnqHtkpME0ciFzfR9hZY7CKaiPh4LeNzoDk852KAYPh+GblYGk+7ROjfQ5V+
+V3B+cYS1w3p6VSINRM+64K1XG8Q4lz0hdqsdQOCR6X2h6RPgWkeKSPlXfy1BceU
COGEjILcsyuYS1th1No8sVRVgvjrn2pJn4e9NLmsK1Vw1lV1Hv9n4pdaH/kakD9W
b8C6QgdnQ7a0+FXnKWadlb92V5Z2NY/rS+dBZerwpC83DQue9yaUD6DJFNmEsPa/
HOnp9Vpg52RAKkQ0PtKddo3usXrtoGZX4V21Qzex+jCL5k60ktE1dG4OQOBKBpHx
hC/x78Tt+szulXRTrnnY7sK5MMj74y1JhnIaghXNY7adKkU9LctnJ1tO+58xZEWw
/mt7UjR5WsUXg86aV3zEn/jGAgfZpm4AP0qNkYCuE2O0fg6B7YEVD1hW5ArW+5kC
NciOAHROMYkQSwaJhYfDJtQILlNA+kdPeR0a5KswS8f4CC43DTkElhAnhDbK8omc
FXrC9gTIa7zgjmHhI45wLwDBAahnM+/jJxvlYF14nvZLUwXZ3v0gGQs0WvQMvBmt
Y5wplKi1DolAOFzkJr/OtYqQImZV4aAYqjAGoRnwr+NoV6ki4gyH2dhD5DbEnpIv
LoapLFKYybnnFY15n3hB6MLt5WjT2E+MwQIdT3sanlueQR1nrDsXSRsdKgthl+P9
6oPPQYJSZMtIRhBaq2d8iyX01ivMQlt9CggZlxFh7G+sX10XgZ1LRw8dSex5lLh4
rT3gFaJsySuBCko+t0DmhJcF5qt7JRm21Nb79r5pM4c7Qt+zjyUPGPwd3NVw8gld
BSdaYr/H1QSuliE7K6g1UelWpkoz1rP6RtcW16CRIMsuWDHEdrG8qxnfRmelbVOT
Aq6xyN4aFpXQjWhTmPVipXl45JIkZNOgkHPoZXdbWHNFKwYRRPffL1i0oXl3B6Mv
vBk1mavsY0dE34bCw13fH2dRekm0u2g3CTP0qMvpzNmL97gCgigTrY3g+GuVifw+
aE7GlUrJpqxL/lYcu+KMj+nhNPshnaqtX2CRlKQrza6ORymgWasrAs8mKHeg0t8G
bOpeQIDcrLl2SW6BAv5ZvxUlEthqbbntN+ru/KbbGdQyBbazeYIUt8IwVuiFv7UB
3Ahojd0OAUNmIh4wpARLgOkBU2afgy+gb17syCdAQnd5H9f85QcNsuVGD58Ueme3
/nfhwKgTmhlyuR9oDAihnl+KwmCM2MNaJ/JeXb1lGl55MBtf+NfdcZIe7XNNJMtv
COv3hatmzZhGU0ofzLdP+xMs7ogcu6LvKaTiuS2Jm314fH3srHeE0LlkJBrW1fh1
/wXnXaxkqxfRDuZLSsnfwcvTURnlgRcPrCgdPMRjWP1VUwt0iS9BAte9OMdZLB6o
5zZE6law/Rw3yFc/aS5CfxtTuR/poz9JL57fBwHfwK6n2Krq/7sJ8YxS1ZRA55tW
lxt4Vu8jVeoalfGB2Oot175lg+BFlpK6lAt1eQ8v6/cX/hpR/9XHb2iE/ise0w47
AJmHOWagr/9+PSY3w1MH0TN7Kp892hDdbeGyzE/59BM+S4Lbt1Ezh+T9heP7/b9f
DmMSKa7c20wYpNV963txt5fUIcpURMO8tJSDJopztJfo8YMCgBeQ84uTteHUql3u
tGxttGZHjKXHj4nW3qLVplieHOfUbdQtOXqYGal0JgATwW2x3svYEObYmH7HFSmK
5xYmwdsuH80xrVWZWEv08VXkWUJYLahHBBHUhOzc+QCcXeO73edhx36cXtz/nJZu
1GcPv4Ibl9C/LLLhwseu0qphGGQtYJ8HSVGbKYGajffGobnY7ad4czU45lLy1rL8
y3XJfINBXLYx/wxZKq+qUp4iHZWKaubpc8T4z+Xjn5JVMV8EX0PUhcDx/NDQ4RX+
1eDyNdPs4HmvIeT+LiQniw5kv7iE+KtTshtno4o6QYYgV8nHXFzfNdJHvAuwnO5z
+Nh/h+VhjRSq6gz0ie8t6vovFCQ/dZAPw5OJRwSlfn5W1V2CcLP2wzsTB2WRCsyN
emEYym1Hj/NnTurcHTmPeJoW1vNb5FPJ/5KSn8iOFHPAfj/MVcy4b/S4ergteqzH
orYG79ad5zLLcAWXqwWq/6yyyndcxz/TqgbzQEI/SRZxpdqh1aRAFs1JZFsHUdFL
t6XauBY5CiglHyQSxf7a4gYZcKG/0J27ogZqF0gLc95EMHAKH1FoHJBzIlAfEBec
kzAfrLN7CQkwVs8148BWmeKC/l36ijve4e2XuLPoxh4FRjksexB+UU6mnw6ceJCQ
zoB1whr9ovMhaDCbZSd8EX0NhS40uSjQy8zqDbe7BtknKUAz9XS0KqDc5I9WjYuK
O1lLnFkrirjxes2palNiKj8kU+7VxV8VUQPWM9hqRjxao4V3KabEfx2a1TGxiuhj
UZzxeJYI+0atuMnhuM07je9Eg974Yccsh/ChqOSUn5OUtKHbEhDRi+gHYCtpBibM
N3wGiBjKSHZ0IPQOY8GDNtY0oSc6v2MS3WIUGUHaPNKOHxzlOz9hIVEBkm0Ex033
Mf8sqFAdwLuFWvQtSth/J8dU/LyCt3eyUvgMoAeZ/MEnNzK19lT/DwKIYnQvQKsj
j0GUhKVf+dANOgNx+DQ/ZmhCjc+Aei08xqYONM2TyfYVpFJ1s1v4heCQbOoj1aWy
3/pPws7lymfn9rgeIUDYzyilIt+x24UOQ5amV3MijGt+Lkgyj5CYPTrseywpH6tu
SVbc7Wdm5HfUtfJx6Lon+Vko8d7UZtOruic9/mEsFy3j3UbfNvQ/t4fvKjMPTjjw
rhp79G9FAuy1gnssK6RnDn7AEJKRkScUCuaudwxrE+PVyMbRpy0xgBkgZFGIgnog
Q3jfI29DjzUSsabq96zU+e/hex0CTKCuW+yLh4Z1zhAThRFdRbUvF+7Ej76WLy/v
0Ne+mJBOrm81rhNjnr1yjUw2t/b6SmMYV7Z5TnvE5xC1cuSVl1zcCrB+rZyZRycL
H/t4FiNES3ctSGMThSkRZGtE9QfxNui/s7noubhlT10V6y+uVEXvJbciH5FszYz2
CUxn8DeIrbrrk9pBMSArLLVyWQ6ksSTB4IqLe6BHdXZPC/xzyU1PDnb2yRWweBdA
t8nAPXW9ud4aAd4ET6/Do1D9Vbihi35rzDkgQO2V8WTBw9uNh3srt0GHRxGat2Aq
Xi1MbZX/mxu2dTdpr8n41J9TLOqG0fNCXnB5nuKkkI/gz0lgNqLoAtnQp0i219wu
OTLUjov8vTNQYe3T/VYieUC4Jo5KaBQB8eZYm1oHVZD4O3ko8PnUBaAMw8KONv39
KBn8Sp2aUFpbdzAu9wo7HflSWRaHiJGtrWPzNJBl90laudOUVHpQXK7oT7vuahIl
VXZRGkO/l2KJWh20Cqch0Xyc1o2UTJdQDmWJf49WCFBsudZex0ZN7OYYRaDknSkl
lKjmNH92eFJCY2XYnBKgv5ltar+Q3sSSj7eJx0dGekQolNVUcm/yx9VLM9+dF642
8ai028kpEs8rD10PoxIHPIwnvvAf1RYj8tttBixky3lTzx2S39LElP3yGFrCSiaG
GFe4BQ4vvoTW66ZyuzhIoQ8XU5mgXSsQj/va5rSJT+t5QnJ66FvRSWeqgsFCsmBM
uvAG2gWyQxzeq6/OxwK5k1uW6KafHi++97pqnPR0YiAjsT3HETWFtH6bqaRUSzr9
e+gxFfQQG4rmNb7WMNRCSZbaeswmRtAaFdqpKX9w1+zcPp8xkC9cX7Csoz4UBCtb
CG1ff969ja9DZRf9BSywzn7ZsZLsm/eFiFuZJXIhylfgwgTOG8U1Qd2Vc660lEWa
Dso91LINN/FiUNH+iqldBBDUMYTKNs+9z7SCyGxwzW5YE8U8mcoQiPuroIlILEzj
l70exc7d/5encROPJ1iQz8DEL78S8H3XBmGqI7FWwZ9KkoKE+iskzQN0j2uS1tV5
vsj11G2kTnJ7sM2QHv4HNlxOQzVovuKHjCYIWiZfZ9gZaZfE/wkxQsdc/gFhhmBb
7IfQOjIGEqTcr2XbbjQvxl1yOB7iuCtmghGpgJdGLbs5GkJVnRuL7N5jjclqgrRO
/Xz1MnCPScIb/txfefrjBDkKexK2VqOQT0zap2A9SHpnkAMc6uVpCuiButVnQG2s
FxsNI+etnzlhVmRtZ/49tmS88WjKrAQTk8irf29yuvsDoDOvuCRtUHrpp5w8b8kO
8cpiX2cqYbirbv2+OGFllj/stbEMAxTzwCVExmNQLAX6LfiuLEs5jLlfzjZTfR4V
oP9b9j0nzTuFIA9u0/6bSN1lfFjozstLuZBIXJ/1+5kdFaknIl1CklyKKK0y+8Ri
Sr/edzX4C1TjXpJu/WIZv8eVMyZ8LKN3gvLfyZIH171smDnje7K459dZ53nYU1Bp
2yhEk9bDzBvV18g5VU5Hn/8o47KfSmIGA2t6Gw8i9GguTok8QQwnoSyUoz4Z4Gav
sJePOEM7zpSdw19P9BwtInM+kkwTHl/zG/Qz/OqQRkvIDbamSUJ+pemDn0rs0g6f
7l1yNoaNqvpXIDrwYpKss8AcnNoyHHOuFvTVix521Vc3fzhyULyxGifP/mKOGXTl
JMtdySbP3WLbPSrmJJwJjO7N8qzpfyW60sDBmp+TUpPkUrBAqZAzmSrgWfWHLZ2i
zABAz9+D37YzuylRLZ4s+EhbeE8/gBIBTebdngdrcThUdZ/TtJR00bE4pmrYuN8F
AXxx0W9IuZQyTlcgYhAdhHNMFsz0oxMU/rmFBjATFtRUvUYCpWksmTaTAbelnpDw
jGRSK2qB80uAAcGABX8xRgoxD1StZ7/2uSGisp5iI/lEBRxE31y3IqEYE/NpgvUO
Dts/8OYqrZFksjfP6KPFnxHSdDk5ZRhWN79EXI0ZMaaRR1QVpGTuSNHC76698D/j
N86yPgs41khPmJT7jLGzOInwl9YSvMljk9L1LQLx0wpl62V++MwnEQUocP5kBxWv
QZ5GoYKWJEF9onMpWYU97odD01WsMaD4tgaMje8ucBC2ugX0VlfvP1dmQi5ZCk+Q
XOPy8LqEqv8NTmKi2Vpn0+UXQo1TC75/D4bdyu0vXq5ZV6HtpTJzUhZK66nzk2GE
u9Z70B5kzJiwzr8cBMAeG3azIvxkwHLX3SgkKCDvNSvcoit3TBHhc4hiwRCI/3Mz
T+GEZ/17gWc1wXQs+b9X21A1VQZTwK3myrkkvH75x4QUiWf8cWDklYjfcigBlCJa
7zPuBY2cZmQ5clvom7OFBmZOzr9ofRE3n9oZqy3OyXRIX7GQcLztyZjILJ7iAgia
UoqnkXNUiToe8aUg5u4gszLZUpmjtFCKCTthKRaj64rIDWiJq18wRAFm/HlMwuBr
YbYS+wfH7UX96tVsBs1lQ9T9NY2tjGgw39KyMujv609g61cp3cBmgxbZ2FlPlfBl
/u4h0D/KBJog8PpcbBuytBasD5x+jNMhJJluqAPaaryPYs/ueBPCEG1MwuowhtHd
TQOyG3rKKC6OJY6dqJCyWXXXVWrJGccCBKybRYLoh389uPoQ4ADXPXqKYR90Icqh
8HP9DqjrWbjlS15lJcceaYwzOCUcvvg0IB1H0+e6TgFIACukbZE9OnzvDtKWsQeh
3upBJTKtoMuLVaK5GA3TrGpiJIElFUnjgyhIwH3HXDd6wSQ14y/85tANwZAlLoA7
WqB5g+VYSw7jVIqhAquNdjv+L0WSWxjpOVu3ptHJkBt5rGUzcMAo9c4r15JEVD6s
r8k/g1v+EY9OBQiie1SPOpn+/PZuB5Sd/h/frMGdRsZoKtz7p45pw1L2j7Ytsilo
6P6zOJZqc5LT5CTYuWPBECVLNUlXRfY8gZC7w+SrUcjM7yn4nrBb2I1RJz78Hqun
t4PoLrrdk9/tBU4ma2NlVa6rYeBTP4r3sadLOmU063/GzKpB7WRzJ7/TPBz+C3FR
ZEAp1gqVlWJv9uaIadhhwjNzjD39ztdpvHfgNDnd90HwLhlAjfytNgL+SRealzV/
RwVvhn57/16RRk87jwxzlnkANTa/MQAPOPMFIu1ueeweYl2MbnHVr5m8eCKvQzgh
IvMdlM9SHcr9XUI8ISAqHwIMjiTyvmZIBrXiGHWL1r6yicC7owWIyrwslNKfQ6la
3u4OI5AE+IdNYI4LctOji35zhfJYI1dVER34Rj9MOQuTlP/umXSIb0+dz2Om0wSK
R6kOtfN8+DfvUfSZ+iL3hsrhHgpFsCWWiG7nV7voJsh1pJQD5o7Hb2J9S+a+GtGB
T5t8UPV3v/+SReHp59AUW3tmH1hItEQni0JPBYPRtlGUpsPpzdRqIzeBmue8TK62
z4SGdXn41ODqxZOsYtcMbM+t2gq2Wq+/DmnX67o7mdfuPNWkoAAuLhTP3fDIWhzQ
oidZ8JzHOAniPcP6T33TZC5od8cgOvZzwPNHcICl7PmweM1EllxBjy+amjCzrewF
tzRwL7TlK8af2Z80oP06R6tsm91fwgGMyjAHaENxNDfz3nIkrzuWP/1I+BTBERjv
kZ85GNuhPCCtQfbrXMvBENGBY4omNbcu5G+9OwpgABQY/oLbblUElxoo97sZ8m9b
G5wi2s/CmtFfl6TL5AchzbIRlPM+LeS+hK5xX80XntqIiXRJAEaVzN0qZyfhirXd
CyZjkDxJJxNR/o8MrbSckYQaiy4/trYHjrmk/i8LB6VofGHJX5LeRGRGh5heKnTg
U2+jKWHVXUi7f7vcfWGEam8AXUSPz++WacvJEGXR+nusEQZsRn8kDS0rxKvx3ygt
Rx5yiXwvNdVYnps9BTt+rCUUu6CmERLVObBUhbLLsoV+XBIgO8O+qM+jw4dHVCX7
R5qe+sNFGM6XVfhmazDwpvukBLkHUJpiYzt4ldaR1xp1n2gJQLmmf1JhqU6vA2iH
HmXvmqRawQwV8shB6UNy6UvW6nk/nYCK+ZDXe4K/48EKKaQG4gaLG+mYGg6XC9NG
m5maR90ejFPFnxXPMq2ksOapCxulruUDb++boNuQHZApTK4Yqj64GrQggiSH7F0H
Ojfp9YvpMRNZ3UvVBpUl/oJ32KTawZ5YB2p72NlyrbSaREuZ9vcls6+i1vs83nTb
ePoMl4serArn4yn/JvtQ6W/1zhInX2dew/M/4LvdNJsNRO+INkt0Z8kaLCz6APA1
4SLDezcXgtAxOqnf+rFPaoePizfslDUo6WO3MKnXTY9a0naOdksFsBxAyiUnLeBd
kpIGdp31Mi0LOjZ7cBGpeSEIPERYPSo/hI0+vDOfhsVQ674LB01hrqdp29s29K0N
Fccn1aw+yDnvvb1yfeWIQgm+Y7T26ckRjVjJqx83ujlNPSIy51EgLHdn2lmv80YR
BWAvYdG4aXdHCDvmwkZcCSoQLPNsq24ZrsEHEcsvSdYAtKG6VnP0KjwOJ4Ekv3mq
Vuqv2ETCuoGahdbmV6okWBCCXPu69Bj1aO2bJe6MyMbMZQ12xzLc3vlterzr+5Tj
e5Z7qvvU8u2ziR/qm4jROm5JUqhk+uJS47Vjux628RQV+O1aTGJxmhMVWR8EFUQZ
XqWxuLednjP7O0XUdJ7nsJOAi0nDZXN6RZG3S/XlQsRET221IrODW7VE0b8RrLTs
ONuGK4JDX9gBTYYrn+FlgvByFdCuZm59ssnt1rMjSdCzkH+daD+0IsiLpUVtSgBq
tJAonDXTY8cXVMelDMVLgEYBEvzaL8I9J4VMqKBOjMJd0SGbIjl/YNAUNF7L7ihS
ftASvc1b190JJheTOvuLMXQcMa7ET+wLPjIaIdSgY/r6xU8Am0eOwFXrt2/RY7G4
U7NF31Pa35tyv2oLPu0ZJIodjyeKiepkAntSuxOL3xHmhPJQUZrlI6aMMxV7XJSr
RP314v7YUu+4VtAJa8qxh2r+psDZcq4TiPTKGmikN+FJq7xb7ooXa62L7utVqKet
yjmfP+Dmc5U2LNFA/YzIRY+cySF+p/DdQo+a1ymZlVg4JOBI1b2sOL2hd1J2iKp+
/YNTsw5BX8gT0mVktadMtMQaeUAs2QSkGgJt92VuGcKL12U1tV7OLLnhM19FunUh
uJIwRDpgLnPhoRb3HIrDsDUlSsOb5apitIRxTtfHgyKjIIB9Ex566eX/MdFi93AX
UM64v8bQp0hBoVK84NwQ2iyHgtDd0Mh0GcgE6vfbZPjEQuv81sj2AZdP5BJe9n1S
NLxMoujR5T+NTKpHa4pKSff08mcGnyTlSbPhaBXIbj97hZOp8clhmtVpv5jqptiK
uWh/m757GC3DDA4sxPVUqqtDRTXobz1+batTyCE6Dwa+qRVHBfXu4LtEcJMfNiz1
CIIh3hBhhCazQ3PRhtVtTIT3V76Zp1sEBUUUFKNlD7sa46CAZtu55TeceeZg+0YN
9gcRfBLBiEW3zoNFWUxgevhWB9qRmIjj6yzfd+JFAnPvk7hhPd9kIPuSPvHkcCJF
X4Oy2nx5qL5qaVgMszubZ/GWOVvIPSC8EE47Pd3WqKJkE2ItWuJoOr5tt+fB7Fu2
rfh23lmEFanUcHYG47aY/Qksd3U8Qv44caTpxTqmX84TfVAvOIWkhUKDz/NMrwUn
REXabKNvHAFxzP9zU2EI9RAV9xn0Uj6N1nqkj1XcWfVJruEY/Aps7R7S+IC7ZqVI
JdFYPV1RErIKO7P+8xGVngeaibbPSsT/ivt6oNhHvtzTFTob8unkJGlXuS1YlqcQ
MuSQPGVziXBWumUho/a0i4ZaGHjB88r8/EpcSVECTkoraFsOwyo67diLLtGCDb3p
Ls5MBEpEVuiZpHhLfozMH47RCE90Rz+MLmWmMgO7o1ISeL9EeQP8K6hP0tIutuSe
XC76oJqldPEMD64i1g1S8FY4O68vxlgwpaBBCxGQr8L4xsw9Yb6XnXK2SjpSmji9
0MgmWTQ0kEoM30FNpOySsCdi0qN9tgivqwF+TrrFEPr3lGjJla6PoJpxz+PjJ+3R
u+oTST7z9E3KWNb+ApF/VJEd4v4/8NXm2NvpSqsQX/Rs+0XDS+5kr5YpJ3JCQvog
kPP2MZ6LKKM5z7o/hSJFwlfQIgMyklTsC6Vp8Ji18le0C9WWJPqBLiOYnZMm1MZB
T48mgJxJd88qvrhsVta/nCt8FmHj2RUUSHkJto9A4quXBi9zXOOSlDVF2gGMW26g
yAw5kosypEdu2VQOuAqD546IKA4Clmkz+hnmxMreL+hQxOe4Nwwu65jwJfV/IP8t
6ewAWfg5Z182iXyPMLBh99K8nmV6hHaXsFHUmagYKioxQhXtAirm5N/hao8EYZ8I
udJ3iFNuUOPwJQDIRRVDdgpl0S3UWS8TW6+s95jtWXt9NZjwO1ncEpGy8OXB761P
vfI8sK00Bdd9BlY8yKAYnpCCV3Z64oThI9POrTqzroSNdrFTQwn8SLKHvSQouEeY
LFqddK1IBvRs7v6o7Na5Yf7Nmm9T/nUyTvIR6PvzB11OlDpAutWgRZrN0gD1WRmi
MamRrB3iRp/hUnkPM3rYl+tlRZKk+2JEa+DKsCRjOdXp8Hzz+1voVXhHT4GFTt2o
3vyYrpC3oCXX2YMcm8bDjIaWhfzz+DjYUTTBy66DTlOxIonrpnIhxuWcYiAsGNur
2AkHiPnvVxelvXj0//myIVkChOeQZ5ON+u5+GboOAuDfsZXwQC/pue8SePBdR7Ir
VBXl46R6f+zgtsmJi0pG3ekl72Pe95dH2vFvpuiRP6CbvRAY9Jv9e79dJ4zOgG92
Le9AAjkIBHkmaHCcXJGwotME/yvJfWycwTdpbIX8lbT4GV2VuV4u1e4SlkIjwGu5
PX+uJu4zC8uaG7DfW+YjWX8hEjprEEJsqUspHzUe2KaYI2ECA2sWPTijc6a/QGn1
Jmp0BqS8fVnXgZ9fsuQmvXOYm89M3WNURFqFkUJnpwVDrm7o62mclTnJZ5nGG5ek
Cb/ZqxJMOefe8zhrnk/yQed30uLQQ0LD1iZwNfwjdL/OTxySZo6VoBsHdctB/eqa
sd2nSzPDoqTZrC/vK7my+f/PHxhBou1IMEFgDGHEoqUKrJnwwSqOpagqvMyTWD8Y
0Hku8QIskeC7y9BcU2qffx0wgHWdTYsfnRERnfSW4UHCU5SRP/TuWY9UYJy+5pyq
JUFmI+TLpqplPeeBvwa0klcHJjkh4h4B9f/+8lppN4SKkeBan1QA6koteM1V+JJZ
C5djOChPnpuaQJy4SSGUiw8sRw0pkQzmVjfxGB+1aYRwSHyZneGu/y4y8mRziUjJ
J3SaXntB1UMIIFN322uWHrgngHmr4uIeGIGfMfUHxHVOiwrbqiHqLT14YPkLLQyP
Og0txl30flurllGmpJ6dUC2l9fYyMmwl4uOqhCpExSDtTY66MMZH26/pRfnfD3Fs
dYwnHpDgohRp2G1hscDYuGjehmQ36rjOATYmVfwP1Q+n0fAjvRSNaMatkuxFnEEm
zf5VA+XZYLtSnq55hdoW23JlSkKFMksFeHUUrR32DAyfvM87V01ydDcu8JMTtr+T
umk73AHu/IC1RetPDnqkBFuGXia8V+EfXtm5gnNox3BMUKUaAVyDQNkaTQeaKMij
AzbaJsFwI2meMM0Pyc9sX8e91Djhf0RWAjVqAzVH17wSz6jI0FYCE+86ZwZs4CQx
AvYlkvWdxo0DtFIN0vR772ZKX8dmXxjEPDre7ekX23qfgr8JLmBf0qpxZQx/QsLL
EUVlKs0JQpjiR81i/kKwyN1R+nV8UH5cfYUQWqlN8NLpswVNCPCMFSYbHhLlU+l9
Z1JIEv9/rI/LrhnrCmZhtKB3pJ6+tkC5SQZoJx8jamz+zVLD/+of1MK2roTjbsdq
VM4IoXzKEf2WYQmMJS6pN4r37C22wHx3PUFxCdil1ZZLje+veX7rrBGIJn/nBjlV
R3p3l0VVqwxoi29aIa7397aS6fzC/lwSkCsUh9Ul2IULWMho4FBsy5Q1WuCVSSeN
aaaa6aF7da1tF28rnTiMeAi40c9zqHKIvc+lspXXAcE+099+aFBttkkdmEkXg5Aa
76SdIyoCELfNtsY/JmyLrhcLZzaibrcRWvjk5iwwwnM8ILQTugrC4SIqcik2Tzzy
U4CYsZwYSiHsztfw2OS9GkaVZ1suep4YUlCXWRP+Fo22bRT0wxkZyG4x6yMmSK2r
VLplzag3OFQEBrfd9QnsPUl2b9NrY/qGFd3rRacreGMnvoSWUg9uoplt9E1quyc5
s+xVpAQHWaYXOD2mxrjO5EO+UUT1qrdlVzlET/a+psgCNVMQFielsiOIhpiHqV3q
CuWXp2iijefgcHpejO3bzvnZg2E7dDjx9qd6x714EbkoELkTlKPSGtHna1jI8SUj
XSZYqYAqKhFMmm0EqIB7e7BuQiAHo3k5AH2SdSTLROrtD8hn3xHiNKPS1aNWVfxD
/Vh7ke2DtdNBufbrEndr8Wy0Mc5SD32oMC9IbGi1nbrHVl0caEj8HBBTnVQH+/SM
7vp1ro0r380i539vUZrlc+POlSaSl886BWYBk41NDL21VW3lE91c+8eIPj5O6G67
Gk3henZJvWiD3aAaiSv2Yaw4W2GTcQbito8Em2m6RFK492UWpIXlMMfJE89yugtA
B3ORlAojwBZu+jwRkJnw6L+PlzybdKwZRI9//SfUqir8GjkXhKe/ETVLNhYrFR9t
eBU7CpQRd31TiHHogqzEIoI2wFSHPzcqnFMRYIi5UH+FZwcsJerwCZLzY2XDDJDP
fOUCNmhjwKK4I60DFtZuEx6tMQ5xe/RPYqJzu/mdRgOL9VKrIqf4P8XJ4N32p3Uh
QE9BnGfRx9rOLTTfbsKEU03G9q0aBYQem+PSrkR9twaF6xxKqt9wzeLGZQ/wq0mp
JXBrXGWcanRlo5iWNFTdG2LBe2Iz901nqwyFUzWIJ/B79AUEGqZ7LXqr5jRzjLOa
2v+dqILu+KuQETkz0mkBZHrM4Y8z4CCh1BKatnHi4JZdUHKEn95bGgcfEwexrgtr
TRNPhoo7XiXAwoTaQIfuUsQe04lFWO9fKXkbhSN5TYFswq/xQpwqBhmweGsr3Kud
D6vW7csRBB6RvhOCpVXX9CwkBmbRThAmu8EDeNG/3Gyx0XzwTgMfX/T7HgLsbsBF
Czs74pnVjOUxgTYaK+Hdw2jeFTby38jWY++94it3txfCKpuUVfq+p54auc97TjF5
WkpU2fVp2148UmMMMIS3DGkGQXXRk4NipzhFjF9ES4TSbH3A7pxRLKDyNVLwRtaZ
7VOjL2IKTU2yfLtPa/wTMGcAHJ7hKyr+0WIfV/6j/mrawvIvwqLzIXkcE19Q1cQ6
H5Ub/DePjeqRCX7SnPE5BfyUuv6Yu9beNYsaxrES2dpxv0MNEH+o5QWC/le34a10
dYod4i5yuakyVGBQAgKQ1V65GGVrTUgkxxeE2Fy+/cSr7EreAbcYSimWAN2TLdKI
G0hz9xr8JkWvhfhyQhqR6pIteX1dKwpXOl3e/Z2hI4nYbxCzSKfU3cEY8wXOojoO
y0T3JgR+ELx5fzeIW1CambSqfhF4VrBIYKFU6ds3nHgeBy8kpp/VEYHXq3mX3omt
c5jXMIbeL8/pFQ0chIssah8BVaiiLlFoVvS8SLkjJKmt4eax12h9gfjdwteH2eYx
YEudl4FkDlN5ehMuzO2Blo1RUbJ4B//cQAbWRl1CEhnYuk8skVlCpJmnSg0xsnYO
x+eodncn7e5LLRQlhUytkSZokoTNyPkEhR3OLrWEoo7wWdmS88/MVIbeDFJjbBfm
pECfyMz17JW7m+sPyCIojIfxJvxIt5XKt3MeUgAFMorJqK36FwD/FSN4I4wvkwQS
jCDCy27O5C3MoyDQsiK8He5NwenF8z1xFjTgCB8gGE/87x+5f0d1hiyg/kxKn1fM
RLb0fo7wBLNeydiVfzhsTLLDZ6yMMUHecO/byxwUQSEzYLqbo7OaWQic27X5nhXa
/adwQapui3x6zwzfvng+afYJtpVSY8B4UVbLmuV3nPKjzzyBvwOms2/5eRGxf3Ka
nYeMS26ARddnwXpOiPGjJ7Pvl+vOxifF2YalAUu6m3s4l33bXtIdp08oTmTmobiB
aSxim0nD+XLXZv+pF3m4mUeQI/zlZX9S7s59wWYZRAloOYQcl2Z69T+qJlP/xDoD
nl4Cw2a+sNmqkbDEaar/xtq72yIe/eAb9T2+1FIf2pwTEE8+rUnZZ9pO51fcY9AS
5IRITsUvoG6jwH5DujYyd/V4dDIoql5X+rVJ0XaGqLLyKfzGlMZ/7hDiku3HDk5e
u+zqdv0sSxg+EB+07f9RmCBVn98FvwZnofbt2oUAXWNVZ/NfUy2ml42Wfgwq++DD
QC0dwZiwO1wTKn5OwRAhH1sBtVLW3/C1NziaiRP3FulwRG4kTGZ77X17CC+y+IhF
IgMoho0y09rY9pd+A3AQE9m7OSqbCvHkI06Iqgk1DRcyJ+LCh1jiVVnDE+B9SQ82
XGYKYW7wSeTTbDAU+Ae3pm+RBVe5zUAEDmMLA5jYXnhJsN2xJ17xoGLIWOOCtpPv
E3RuTR/UpLxzOvi9G4t7Twrg/ozKLKyF6nCORoauOdhsxqQirXwbwz7t5Oa+koST
EUwBwdgMJmaON6K68W8nA2NgUMA7LkYYG0fVTrEbxJihv0XXDaY4f/v3p+grqUrg
eSoKhkdoq1j0F/0wfjWdfx/6PklIsSftGaIjvJlZyBIz9qWCUodDk5zvBzeOw0oH
slZreCgePhksDg4rutTtRwHg5B7VrLEUeBC+RZ5iKNLEwx6Nw5TnBB81ma1EjcGk
KjiGjcyCNO3HaATAbgxoXPqyVx9uQE89wnKVMh2aSZTQ4YgSQ6gfeFTOjZ3gPxvn
tpOkEKgT1IX5223OLn6lZlQFBl5uoLJaJ1ZUVJUUv6ueNqnn2OxYbSLb4O52PUA+
pA3u8usZfMGSGdAl5SEG7NT593zBNEsnebDicS5UKqZV5hOkMUwziQmAWksH2p6Q
CsE/tuhQs2i5DIx+QxBAEetCN/i4TEwhJ5XBRscsquFEvmQfnSip7LQ/9av+z2zS
4hVtrt8RLMYyLlTwbQmMNoms/fIWot2dnjxZkEL+ZlPvzARjPsUmdJZC/ZmOhLY3
DYBH+nowdnuA/gOFBt/WbXjc5NH4rNGEOevOHduZfuRi4mKBprJUUZEZcRiMtDzr
qMnQaN5xHVjUmC923YaFxAj0ig3HoGAICzjLve7BKkPvD5mgSlEnzUQ3iy/ylMQ6
nu15JTQBB/ooi3gSc9TGn9SP6AJRJO9XTCveanUq5dKiiyTRQ0sQYlYQX9nIjSZV
9paKNZEueAODSzsZqyNKgTbep+Xc3Vo/GhLKhp6gSGnWlFOBsnRwoQPDw1Oqe1Fc
+1GWtWaiDcSJt3vWKBl3a9GMYXFzqIpXOASHtSLo5k9kt9V1qLygWUsRYYx6KERb
MXj7AZToK/fp6hf9XfqAzvBrjwWaqhKlJIbFYKZ9hKuw18/EEq+kLSjIEZLe8pX2
WYSuFro2zocbq5VEyi3kcjxeJjTpd/WJbDzfIt8+n4NXRa6MhIv3mi7zI5xVvc+u
X/KfBTR5D5g+9sOtnq3x8QnRSNW20aEGGOt+hQw6fOdbYnyUWrH0pNk/ODuqL1/x
YSlh4+DD9Mp/lb4qNOsFBqSiEZuCcdLyzrQ9ip/WWFpS37Hx9MdmWNhzwVkhupvv
tvsU+Ztzk0pTp+Q05nfgDmvPwsbI67kZ+SYYihRMyCoknJIgcd1O8bPvAxgeka38
C5R5t0Zqi+05X/JI0zMZ9GohFGb+skSwP0Ab0JSKdP3rQrC7t9yqjuXJCwIBWKFR
fWtPfz0jnB8VnQnTvjKxNN1V58rxlGy2weLxiQFxwjaSisyDrih3PlTu/ezsX0jd
wB7DvV9JlGshet1TxGQYu9NNHd4oVL5+ut0Krrv7rQEkyyHXIM+/rIKB5Aq+O7Qr
f21vE1ZnsPSzAOilRVr1OqlTHR/arIZsP8FWR9PFzaYUlra4b24B8Mp/6j4fKyXZ
/YpSL0QrY6YC3Fp7Zy7Nxg5lTAhDeVDWowNw6XmUGD/mTlC9JQnMWQPUjTipRiUj
flheVNMfIfeb7deeLdpsbQ54dSK3zcIiauet456kNhhhS2FF4b0scyYm4IvFUqHC
S0wC4SLlrGW/UeAc+pNfPhJwNTT9EnyZjixsNOdBfYgDhwJJddk5B8QsZkf0no2f
3RypKBAMyEDxKEq3Jzd7yB1dAa7C7/nhjqdwAq67LEBtLWTjrtx1zGbbhPEZUUue
hBffo+9coLIJ4dd29JP2jCEsl2SCi9Rnso5NpRc+ssC+vWJbHXzgeB48sjEE1Sye
5UYytktRgTw8KksuDOlxBpI7i34hNyvOEilsrnWehqDTiGnN21sM1eXyDFwd+Pzh
6DQKLr3qqrgZWr+LE9vozI7zA4z5Ne7XwwrcM2DiQsDRApBc3PEOsS9M5s2DCgjo
pCiV3uSHZu/PhdexjoJzgMJsXRSHNk0lgxFqk4wRw5q+goGpeJPw0hgt2v8EO+tM
uoD1CHuMWIAb9D4oI5Uf2mTzlEw/Y8xtmoNNLL0lJO4hIeeAR0ALSS7/h2Nska11
vsHuLc+oHWVKXmlpjlKnUm8l3pQXGEX3HcN8VaMi4XC0M/MC5sHSDzkbeBTXAFcu
FsbRlrDAjbYPkS3jUdWyEHO6Z8Hq3Uvq1CQeJ7laN6hRspNK4S2rZDe5VksTq69b
hMc49zVze+JYYFbvFFI4REGLFdZS0ZvdWJvFAq/t2sBkniGsYHIvKB35cCDUUZyS
KiL7oAq9lvwx0RicwkrKUNSf0Y9lvopwDZbYJpuZX6xotNm/S3ESibOBew9L/Vkk
WB8y5Ojf6arNYiRy+HmNgz85PWxY+8HSG7sH1Nqa2BmoXad8optbW0rfiMzsKciC
sR8NrbQiTOl7U1DsYz8U66B5tfeZVWsH9VhsUxf2lzN2ZuD6qJnQndObO78y8LLW
ipM0xGMEO0fxk7lT5W78F89JWe1hYZykFvQvkybHkCmzuDd1qsFJ2rCEdXzgxFXL
UmOJDKMC9ch5Hv1AjjMX0A6jRhzU9TZsh6Y2SafunyToZENFsuSS9YpX/WFpQhRE
iZ/6aMl8guzEXHg7MtxhzACg4bk0KaBnktKjPg6oA1s7/zVGJl00YjRYfIc7t39R
PR6chotMiNW59xZzAdWC5ome3qeCx98B6AlWeevtiqbwT7tM6sJPOnVVxJKoVJoz
fRUICDQ3V8YztOCDlwenPCt4LKPLvIHr/3HJKdRkzo8pShD84OQ1oyKywRUeZXLZ
aXCbB4k7J2Os0FqrfGgwnE6GnntTp7q/Fu5aV2Aq+8f/Bu5dr54Wp/7iHQQnyc5M
YpArTqNAuqpi7ceHipCR35y/Gy4HawdkqehLu44LXdZKLtoNtirAtU5Di9vgM5tu
hKQ/mUfY0smIgP1HzL+7WyAZ2iaNiKO3YQMPatpxbiYOjlbr9wfLV0KmsK0hIlUJ
NmY8VJQlq37Llh4gacRh5ZQd+4aEgl1iismCZlJujmNJfFvTyiUeuZqMU7HdKwdt
Y9rq39BHABZzRscfTEbAaBxctQpFUBTKJw2rIVcm1Ax6KhaFMPuphOfgff/XkSHe
Md+PJYTppC3oJb1J7kweTqNAEpcXDlOabe1joc+tw1+5vrtVxVCAnrwksBoAaNpo
COXMJxCG1W0+kwpaEF1+zmdJsy0YiVwQ2maeBOry5FhST2TyES0vEMYqbmGR0WYC
EzzYsygifwakbKjpEIY/rM2zaL4jQW6icfsCA6Pf3pFmvIj6wD5b93mjJCAboZe6
zOWqn3dW8aoN7z0gfsebElt7JC5fnoMtlPX/yMDQgC6Q3jZcC15CBN5hDv88n+lU
zkTwf6OiQ/8etwV944K/lbgeVSNPO/ppGkiH4B5Thi+1fXi4uxo44EMlk3mrgW2X
grhisCM+fOJsLwv7Bxq8xn65xeFqSHZ19r1hFXR59zIiacVii65c++rPXRKe+1s9
kqXYxZPUFL3DIY1HfWEDdSvtpUMcsyLi/lfatZAMT8JlcY3N94Z4HVckIzalGF19
/b0p7KG8gkrPavqCv6wAQGXo0vajuMMA378gp5qfDY85VUMww/932VsAz29yXWdR
Rs9ovIhUVqEq33/D3ht9TtQ5ijLnKHXtThTbKcPZofchuBGNkVY0JkB/qOe3GxG4
13Rnv/YWTqtmBQ1JOD1xDbhA8iCLEqvPckN8MvZilcTS/HnTVZlIGtskXPbKlk93
XHPM+dySp2GSJwt+fjJvnOYD8Wk0nzdzVEKAztBiEZLmX/wxBa5f4ZjGGBA39I2y
GZQw7c2bYQa9tKJ93P1VXrxDwGUqcB5o5M/F99msOg9sf814TlSZ/DmvRQQuq46k
0kqBa5KcPeJMS/+2EWtOtguAuBL+wdpoG1xwP2nTMuoXidsdXCncbSsqsHYuzOsx
zBZPE0LQaPUuctWjJdNmSeI/LgBpW6Zqw98akahG+kB55paSaOYJZCkdDsegFYVU
LfCSyNOCGf/ihBJmtdnqDw2qWxIalLZ0u/lz4HMAzEH6pgK4A9nQS3VfPMu9jL9Y
Or3B1qgcVDW6hUXHGv3w9vWykjtyRwMDjz271wLeK/DDYy3+2upEKvgZI/QYjJIg
L2fygT1uHh2kVESR8DWQvIt5QtbUr7pBIcGdHyOaa1d83zPcWUDONJKd82Xu8eeE
RGJlX5VUAiX9LGHG9t72dFfdOgsBbDlYGsmBAiKi5HS/9t97jhdANLEdPTdJH489
qj+1AEojuP3oX2ckC0IphxX5YwgA3OM9nDZoQ6G+isJHgEGv22SAAqZoakUBpxvW
zyZvOZogIiRZ8M5AqeTA8uBoXpI4cHwIFnsVJaag7NMYQfrtkTUVZzw6RUHITEJN
whryl6D1WGRpvmPiajbNJ3derHir//SytvX9V3Z9EBqqzEXTwXTg7QtO86WU9XoQ
WQHL5UnnZYJLh4DSvvuUpqxumNXfDGbVVzp3WuCmZbVANFnNuLsVnuItJzgCkMax
UDhQfW42Jt9KOKh0IVZTJTg+fvQFIVF3ZAQ6LaMGmibDGl4bnSybFLGNgFQwoud5
8kTED9Z4Y3hRD9URhhHUVrgOVPtBQ7khKQlXsBd3hHszEl2Rbe13SzjpvJWA0OYs
XX0qvOlvhk0tkkq7HkXTIpEG6X4cKOUdC0g2YKmlLZqskePwpFc/MAlhE2h1IKao
bkqrP3XyoNuIGO9KAfunux4M8LiisM+4GolWWmdPi3YOYxJzsd3H0+8fk/YZyq2f
vG1ol/DLlAUtvwZHxhF7miFmheWuaLgZly4BnCQO12Jf3cM8G5aRVemqEt6FhfYD
tBSsca8aIeQIlFg+wHeoLtjYTFohgggBqAtTesR8b0R7aYuMdF30xerZToaZUegb
BWPTvnsHDVbddfpuNvFLpzdGyZPh5DaP14scsgcNJVywhQvEflmMK6Z5eaDf+RJC
KJNz+dEq440WWd7BZomzF29KndyK6tprpBFbU3GvfL6YoiuhC4zvZhLY80eYqzx/
TVFHzdn+/kAEvrOwMIEqF1ggnX+geCWbAEv/oxSDsE3KpzSeJzdOL7fLaZi6B+EU
nB8FkLXQvqRGhuVkyFuGOwUYBD+hYfYhUT1HXcTUlV7FdoWI97m5Gi6u/ppVEl0n
nk5ZhIaLl23AppKR3RwuK5hsb8Gvps1G6Rnzu+WoEC5rSGEP5OyOuZ1QHb8UODzg
JCgrmwUN7UcF+hMqKC9wyhFF6EHfyAvDP0jyxeP4A1hw7NjXfzw7B9gl9IYstog6
fSHU+GYWuDvbfBJZ1CIIEVLX+2ZFmGYHXFUh2bftyCZ6+vtwbkW1BfuTDcUZGgbG
Fo5C0SU6i17XT9hJ4DFfdj7pToZZsiuffLLci11jJZlILwGkx8FEUw5r3Px9bZ1e
NnTLvv0vbJXG/elfPSPLKROhjHLbE1RNd2FO6f4/RiOMIKGcJrejUqmh2Iop9f58
xzOgG28L6b2qErhjbjr6rxLvoxWiAqmvC4XscT+FzrGaeKhXWgYHodC54LLOgz5V
GvOEGamSGFYHsRKHo3Bf7EiLTnd9V4ghQURsNLqnY3dF51zgv8iRz5uALLScXSyY
le23WB7xUbfsThoVBWgh7Qi+LcgoQU+LbN8xPB1V6g7y6sVcmDh7X/1Gb9ZIOPaB
62MbUthWkKJMXzazeAvORrJgV52vSkRv0LE7zZieZVmePw8tvm4uszR/4FtTuFfE
B7E1LHQWSG+FXJDfEBPzz6pa46cUFoyWthPZWROCW0dcrt5rb+KH2HI9rDlCcgLY
VpX0BnLsTklym/IxX/0qSFx2hPEyjJnH+5j8EpgF832/vd3PvYmbvA8lijo/y//I
F52yu+d7C7urqaPZ3GQ+rgU/Yv4yQvVWSR3ap1b0+JCGzy1v/3IAo3//pLv5PkfS
BeXa1lACgO8ZzAlRky/8aoWSlJjjlBmX7LuIQoRnAcDcf9unzdUUm3f+1/FvUaa/
f+SPUtNmiuhUXpswJXWaCeMD9xrxYQ3pYk/kE8o0klvlW3VT8PGEhzPcMTkD6L1I
ELf78QJdk4tReYFCcTPpJVxZr7U+XqztbgKCu7oM7uPH5o2VGK/gWEVdUYCvHZzf
7BSai2CC/aXy8aorv7yudtSJuz3DiIHUl4L7G6pYaY4rbBqAKqNsLWsZpCekRqDH
9pvEFu+Lqfy8gHZpBulXMDWSaCEPZI4W6zadrQv5+MZgChBKApAU7kAP5rRtifVK
6ZMr+nyZ0zp+w3KCRwXtKuwRSxydJ8P/HxrUMROd4p2wq67QACyALphzz9S2NJAg
grkkTqSU+xjLwWYKmAR8rVEM67Whdi/MHtydScI46JTsePe46nnSKMTBdoEQCBl8
uYFd7mwWWdhUGTjd0LQngCCZjfQL3xIz5fCsgTyU/jV3WIgYM41jb7Xyl4PRx130
PD7wuwjoDC3w89eRxeKW2VN6e4WFK/Y7o+S0Z1FJYwUmJxA+SFLWzre6BDeH9TXt
FieOhVVwHDh7neP8sAgCrVfc9Mi4CvouZQMB5r6FeDyx8Oht5j/mKaUXDNEsRJMT
UzBWBlCTuN2Yk3hZ3gArCOl3CFPgRR8J2fgZvjp5zs2gIdX5ZOl3RDNsat9xVmbg
nckRlpuXmAME/C1ApHOzXji0PPuSeVO6w848+OJ8yO0TSbbQ7lLuz973WAYoHOI5
GZESdDVg7zWR1P5YtiK4TIsV90Ogr2LBWIFwg9P1Gv1hDm0fvPnGhaghwfhtBdaF
waYiHrksBgMmE8kv5taewZ3frUwPDKAQYY5ugyDk0KBzuaCKlAkeIg388RU+KL4q
YStzr20BSNM2YrZsAD6yU71T0DAJcZpXENqdsEi9YN7Xmva1E/iuKmG93xCpr8Ug
668YS6ZToS8uOZaSXLVLr7Mb7g8jwwIZfWiAeNnDBALEtiayZKQfk07AvzFwRbtU
9grqws72CF59R6PgQ6g1kVZ6xOD6f77qTUtuwh2E5ZnWcr/99d5mLtUj+FcHgyax
xWtHW8QNvEA11UiewoW3AUCEO26vUQLwIlBetVa9zpBb1B5hVowR2HgEQH7NPfw9
YZ9nLDyfy14TO9xDQnXv9wz+aBpvYEwgK5AHaRFhdAMjWlhgXFrVSpwPLzzIGrpR
eqzm9Iu6Mz/P2W8p5WTCzKtHBRt3VA+gv3dtGxQo99wxzGDQOuxC6wdz/fh3VhTt
JJ/nx6kyFcZxQa8MjPBiEJhhal0eLTcukev843uuRa9cVxoLwCkdaOpG2x4o2q2L
rLtX6XadJyBcj0QwQlTIEb39eVKLwdKr0YnmTfLNI3fcUHZSE+BUm1LQXFLxAYwd
mthWltTWbu63rZdm1QBAN/TYwjmg3dSRRdZRPteiNleoXnY0jYW3k2uBDVlcRBHD
vERJlSIKYMk8Y2xF1t0NvQxcQG9vEfUpyCDLu2GYggHi9N28wR1jMo6WJH2HpqSA
8OTmH+PgcZ5LAXHpHXc3Q9kRUoEWg8J4PXRHI2yegKxujm5k7cUEYTGNYzeDUMf7
TrF1MZWdwGGdum9rwvvTaAEMfebYWKRuETwsG+mnW9Lv/9Nd4NAI/aNEOdoBocyq
cwNmbS8Cp9IFgWN6F6wSmBV0W94tAG7tK7i+aj3A1u0bXApOL5MUF3lm2R3lKkM0
H9j6JTTySSgdaTRRlxfHryhMgPfBao4jtxA42pthmrtW7W0+BBYdYAHBCmoek0dU
GWbKuaC1TWNTBb0TvrJVhO/o2iBJ4/3rYKEYLm2t6eYv7+oC/fiTQF+LnE+1/oMi
n9ox1ZxgbkesaCu/2LnfwNF9ws6toUIzGij+WA9LdAUoBGnxohm6A4Wt+fMIgEO/
JXO/PgSJwqb8QGZJ+P/FAZFVMi0RMfZW1e9oQOADDZzhiKeUtHV6V6og+78w1alx
RtO2W2tHv3PkmsshyqEKQxkzw/TNjFcLcu6chCX4Z2yy/lBNgpIIBUHGa5dqK3Qw
PH1ASti+pdzljR/VkqQIDp8TeBGX1dOI+IReIJAI4W2QFN4COmtYRXwpDECwZF2P
UdVeqbyV+8+tPOSywi9OTLZ400ekDRMOBOqoFjgVVpjLa2VHoJFE8Ez1jtP6j7vl
x/4Xr0XWYcURCOB2ZryMfZZdmanDvGfbECTVdPLx2UNS1no4JU0qly5jwIxFHRcQ
A5dxBEZCKQfRcJ82abzbYQ/d6mAdKYuDAET6Hlao6pL7DkbDUVsivp2uzF3qVWjr
gLC/hB6IMoSn5AJn5CXnIjFO4Ewgand9bf7Wfindls69DMr7a6BES3AqjhTBgC/p
axRACOEZ94WNnUs9w6j6XnKua6wFu2AVrhC9cFmhUdoi0Fzsk0YIHJMozDeErtKx
VLzt7XFLfMP2jUziAnYTd7ob+uwhkyMRorCN2b8mhnCKyVWn3sahTzK4U6phhiIX
SEmtZv4oBJLZ3OBgx00IZ95niOeCUG/hPJ4pdy4d2mh5LYrpf7O3zvu1BjW5cQwp
xeL6KQEijelPf4tB/ysFPakjtbUhUibt4DOckmc+MeW8pIMvfsa4k+SIu5RlZTXh
qwigHzLJV+5kQ7IAbuFrKZFPiMaAvZ6TdEGDB1VSrpj1h5i00qJTwRQQXEOm9evs
9kALC7eVrHmIDnJH6zE+YLxH7lkrGX3MbR8qyyS8QHJq1k2MofKHrT7EdxDz6Hta
FgssV+JgPWQ8JSDb+vPrUNQCm/MCCTlL7xbk0urcM9war+4k3nzJVcRiXz0PvyR4
zAIRdz1MEM+W5od8cVGa+c46z0bQq1Yf93GgrcMg4D8274T7GcqFp/JdrfyFYTAa
Sg2fIKCJ3d/6vWyGI5RX8xiAq+qmqW4M1/+ZIBhxUKABQjsUaeqBA1nkJ9RY4DUE
KDColoyud1hlIYs8ITl0Wxu7VDNPnft06NYT0VQmEP3K8Hmgnaep0ovAYCRSAhwv
wF/i13guOb9cvLT5nQAvLdBppzoHnoUETfuDCtRZlCkKze1bxLKHUZoSZea07yXg
dBwE66+wOqe3DpR1er/BSbGVfptNESs/Dg9dfI+5+OYqrKKoeAxL2gSqEc57Z2Kx
0SMI4c82VYOnkAiAA756nbx602cFprCix20+hP3vThon2YRXdIdDOY3iQ7HsIfxZ
RHuQFk+0zMrQ9FGdiCSZCAh9Zf8sbwqXVWdhqF61ea82rkrzdoPUq37V8gs7SXyv
OVwgm+OGG43KjEBwZZRGHsvNeDehW83riobGzw2b74XEqcbuIsslOTUPT34EtEeR
ZSw25uFihdZGGwQ06TbnAIGJNHVTvzTGwCqI6OLo4VYIjeZ/ItlMDJVcq/t5b/rQ
U5H/dCYDlJ2K8RY6i8CrCYGNcSeMiTyR8mzJyE5NHdkF7EtBCu6WuHPLuE7QEJJV
9041XQSEFD6GhJl0zzIGMtUkX9dH7WmRIhtCof2HJkKqZYgORJiFXjKfpU71eUCH
cGMWwuDPoMa51cRiVgrJc2agUMRlosaHUV9KwWU7tu1j3VpI2BGCEV/zTStTqRtP
OHBhJHj7KKuvtBtUO0awwCkX4hgEjEXIOCSY74tbPRGaX5bX9x/3fmqnyTTF0GSJ
AlXBoMwWBGSF/UBqL2EPB0N704FVpfOErgGCYNh1EAPQn1dpPZEs5kRdCISRBlJU
bO133Qhr/Yfc3+FsOndeGo/vilLI+mbo2PG6dgqWwtU472usPyChGvy8rw+dXYZK
/ANAcXuzkZQzqW50Cvl13PNASiwYhGR24nUjcr43hMjKbrLfDASN/T5K17RJkK68
jfvWL/TkEoY+sDS3+DhArvyf0Cu8L3F2Z53cTR66xyGhudb9RzQNYxPwloHNMjiF
YazcK/1Y7L40ZLb4gKLi3YA9js5FJ98r6B9i1d4LavzzAbO8yAGaKkqTysayaRlK
6kRPRS1bqBzNg+IMRC34dKvvvyvM/KdcFVNrxbtvYy8bFDhsUZvZtInAeBCCORSV
nirYk5mTxEWOtPHmqQsPtP6OysJ1DVtJFlPZckUGCj3Wzqw+EaXaYFJWvMfdSoIs
viUFeh8X8ZDHXNp1OEYR4Kb0ZgdvU2rHZtJOGiLHvxis4hUrO+oMXr18WsNZGycS
AMFYJgUgsMSPiokc22yaaZ1oIs/hmDriZaTQa+jgsNyfcNRY8wxgWglKkCFQ8Ybt
83CfVE2StGObxICN5spHW/6NtR5reNprL3sbHtJlxDBUdLWcAIMNlkW1SOOtzvt8
Jt5X2Gt46TyVtwKnUm6sBfHoj3bc0yQrt4LPE2cjiM9X96oTj05kmgzVSvCREY5p
n2M/12BeG0kD4x7RyaxKCZqwEuAKrNsK3isUgs8pMB6/2XuD77AYq0WUF9UZ/hBj
/b1rwOy0ogNLissGCZQ/PRSX6n2iKZW01tUjJ1DGUwJg0RHo/C3hZESUI9nLqidn
N+U6qrgv25qhO1vG8fHBGHheSrVO7apfsHnWgcxf6oMMl8JW8MzPCqraeKHcnRqe
IDgT+gBysyx+dH64S+oaL/doub1cqXRoVDbISW0aX1x5IBWIadndHYPREF63y2jt
W7Lnt/ciAcvsNzBCFuWsvSDtS+gk3VxNvqZiewI9hALcJamtopFhbRBWMaZ965wu
y0dvwwbgqV0FBmTAQWq5p4K8nSkAvEMSXkq73pu2W55l7CffKucEVXCH1EWrDmlF
NgJTy2Ih1dGKqkOqFg+NGQ1YMljHZlF59m4ibRNaSlNToBpsguQiVKsLCy+Hb4lu
soKXz9vgaAvvhunXpQMVGSIYRvJVhCbQVmzn3D65I6iSKh51sSOgl9FmIcQRP4c4
m4V7S5rNzgRjPhRVZ8JLg4fCc4AWODi7kg33yzwPcEPMkavxQtJ6j/WLsCKmQvnA
yM3aYfIvfn8AqPzq2G/bT8RHFMJnnS2x3y0lxKxRMwRsgYb7w6QIs9J4LW1A0vUO
Y4/JlCMdMeVAmVj45IurO4cm9bqQbULpn6DG1rWi4np5e5gYCZM8p3rUT0Y2pAUZ
r89EZIryKCnVoCLJsXGAEQ49Iq4ZxjRzglHHimuBWxo8Fp1uAHJYSk44aULle7dk
QmOg3llP2s9eEfVbBC3P6FQehDY2nTk5YLnNUIeZEBMzSZdVCCfB84KfESxmJYxv
bRw4SguEDaTccCGLC22ymZbwrfEAqeVIMSZgGE88qt2N/f+9cKTrtn2fqqwaEjWf
foAF3ZHEcAuOvwYiYrxl2h7QulzP9bto8LsT4mU/7uMUMmuvVrUtY04qNhrgzoV5
ZkMW3RrB/qxLju8VffuQ5c82ri2mCgJTSK5gG59dIsxdyelu18BvMEtkgvv1vROw
LayVMRVLZaC9rDhfoOTE73njp1GfiIKZzjihMBVUAPxSmBrhN2UrPXzzD4ZaDqSd
yomaaqPQEIqXqJBioOgfYdwaF4tecldbFe1lI8Qp/vVG1FdgRjosNLatfK1cc0+O
buXwzTCoMZldZxkNTMLC55PbnI1UTtL/H5Rn58ilqjjeJakLkcydp5dm3Fn08XqS
YRr8TYPDJKFQwUUpEykqAXICU5kjpacdH2+F078iQDyrtZf+Jr+goIJYDdKSta+M
MkTjioxL6iDsaqtvNKSkI/Thabk3xLOG40NQZmd8kV5Q+exth17v0WbKkUmJzZ08
XOuejAWcaPajNcq+iOWBylL5fkub0FlH2RN8D7iU28J7uqOcbGsoWoyT4OaYOAga
nPHHyjYz+2rT1iqW7PgREA1wTnbA4gupk8+VNwr5H9H8B5gLfmdr9k126w94QQ5A
qblp+ZBpItKv2qjN6GWS1G4FuabkjqVwD5FyNiEpQ8eBNU6k4iY1HXTrKeUnhTW8
G9k9/jZUiOsP0Gkl0YHiqSzKnc8CI3d/OfhwMUFl0YSJDMUDNrlovUHAmSW+Lrsy
VEyTxFJ4TbBTYsn39UZC7Ct+TuVkJK1wj0PR7G+dR9kHdX8i/iFJrLVE3UyhJPRO
ODHHBQHWMFQMtMqGwDM0JpdZPvBFH+15ssX31Wgn+1A//cNdK1Y//E4v2H9QwJi3
mWSt/oiowho+sLADUx4NAVckJmG1U727sfR3VZc0g+OPRrENNFb2nD/qESGB6GmJ
JsE3OEp+NJ10X62zpPi6NAhIU5sv/0Uv5zHMdlHvDlrNVwZesFw63rtvGPhkUpjI
LD1kBKH3Jk+hFTMb0jkCdFueqNUCL24t5+kYotK9qAe4IpiqHuT/a2By4/2tlYSr
/cXoqxBPkL/05u8GisBPnu9Ba1mkkrf7oV2poR+caE4eNwVgcdMd2oqQZt/Q0vpz
+g5C0RaNPFWyruU51M4lh/qOxexyx/GbM1h5KmjOlaWsPr/LQGE0EujtEf3Ws/cq
DQnhHp3/5n0ySs3AwxgRZ9ZTyVLtoLLwkQcr32odfr7OhpnuJGmc5Gs/yqMkGSnA
7JdM+GavKPdPLy3swwst5FjCUmWTfrITsWrh6gA/dkuj0S/N9FBBNBmmRPruKOOp
sMDCRXVW6RpAHZBJWFCdAyl1aCXColaP5WEGD2gZBk8WJYw8OsaUTbsg9IcA5Uuu
xjStHVmxLxWFw6bmhPibTGgd6frui2wiCQU29vgu8JRJOl0ZUII22n5l7qqw8jA+
EzMnQLLrR56vnB8+AnpdKXWt3qIYeRUYFV/+s5cfFHE4ls/y6YoD+tE7ffbqfRPb
7zFhf2A3dFHTB0h4RAidRzTGbi1IZU3Du3txjSHQqrbrdY79QWzBz98JcaYypIJJ
cWIv6AhOYaFnGcWRrAE4TmXRdJ9uUb8v879JGuV35xGCs4RVQSRYnRZvnKdVlUut
Q2aDXRptWFDD5wPDGM78lEgvoUjb1j5BF1xMuz7r6PtgShtZFE7mKmp+ajufiRNM
/BPCK5OQNlW52HGxmChpr3MkV11enBFqSQz4qcPcNXhaIwpBkzm9i0N4pLkn+XKP
Q6X1yFq3Kq5nInOucl+DmoRR13ptYPxviCf4xGKwzGOSjC46T8/bE2wnI5bh9PxD
m9pQzo9zdJnhvjBkyYiCEJ+0HRw4b0KMbxp/Pehc1WRrvK4pzdUpQ3aB2TahY7i7
boj+SniZp4SmvSInqhUnmaKXuBPx2zHGUm1AvZdFVL8UBUewDySeuXaTAxvsnoPr
H9Xi9dzQo5Ntuh65myjNU+YETv9yUYketdg+sSjiUT1I7KiSEifVdelyB0lxAuPZ
US1sW+WPILxzszhqxNJ7TjrxW/YWD1sj6sAiSW4Vjaqn/4g7cASoC7rb4YOZVV3w
5AYvxH6MsW3B3KuI8aOT9Ny5fTuJVDj3Iea2rZOLNVJ2z4X9QzFjKoOP/7zKhZ/e
81/IxZG7cq3dXBs/LLqB/RFtGNvORo3LZZlLsc4lgWxMjgw1Naf2PqTkwXiiQag4
qI+zWuFfK2eI4INtH3liUCemVxsNgy7gn8mBr+LZ5lbQVG/EVYnJfQAdqLfAsko7
74Ewdsdb5v5i6v+KF/DqTlq7aOUp3PPh/YSDxb8At0uiHy3MZCU3n4Srbljy+17R
dJCmQ6FfcQu4Ku4bPE9th2fy+9t1WLcfgQcjWY8schmss19mVx7/Lc0d3B9WXB5q
QIlLvHRYrNhTONB51wdI23xi6kn0viaPY79TUWtb95fgECxpklbgPjquXk8Cy1Zm
F8d5FajVcVUWWxHC8WMF/pIS/x6irEdfaPMpO9hUV3vF20ztoI6QKOiTDNjL8OIP
wCCKNGiraAxOf/kWisuEQd0vLP8qk+mZu87myn0PRtrMu3gPxwS7sD4Tc4XMpzQ5
qDxuzuB0w6ptK0JfWeKYOM5IOXefWv4kEu+JJebETRjur9Ru46ZDgKj+fpFD19jO
EqnbS30NLHEzJoju3VJPGN25gtw2sRHbpP99JvCedRmV2ahOaObCkMpvgXGVvEHk
LC4q9ssMmZahqhIlHv+6uW0KEq0OnURhJl7AO1xXLdUIuJcs1gIiBYFK4wZEHAXt
LaM3BbKcr6PuJasEpH1IedCH51Y6jEP6VussEe1g1yMrZ18KPgWYkg9l4aDErOAT
b8gc0FdtRhsCBkGarS9eh212ZEERJomVkC+OhX03embFxrJLZ/7i/bdgEnqqLPtC
a3fAXbe2Qlc4k60uTavErhjiZQ5nyqb1b/1cdhA0lH7ho1rGatF2GO9Nyu8S1mVY
vLFpTmR6WoKwHhk6mNNRxIXKVSUwLbgapO/Wxvur3TbzL8A2mE+JVLYnbk1KkuQe
2vVLNb0bhLCHWk4Y468Q7vxx/O7aZ8NcxOqw70NlgzCU9bo8/dnFXfC5D6UC49BR
mmE6Oyeydi1GBUvE8cbamaP0U/R+6OcF0YA6E7Bh7M945D/EeWkKpcqWWwd78XFg
7sjDS9xu+Kj7HroyF7DIUYZpl9aBE5A5Ni1qapKhXRycAyJ39X5oF2hWZU+Q8or8
efY0QoaFli/nLOdD+cNJo+4jw9GC1KJT7PP4WZ9A9gbTaxldLS8D6sXKSh3Krx3H
ExSAryw1uzWUDQXVkP7CcZ8eJDE7qQZYIBjzmd6GZCqUtMsxqd6MhDYhMZ2LGOyI
FqxW5ubTTJkv+X538TOCVLZGrF4YuJTTPltwQozE5FKXmzBktglM5BmMUiOg4wLm
CV4qm5HDM0fZeIfRuS/r8TLwLhhzDu0HpOI430c73/e6yUPOI+CkBL5QFKpgh14j
EzC8vF/0/PjIOnQ9tIT43rSVR0qlqx4FzK+k1VVEYdkYv5A/yXGos37TMBaUrhpn
Fa3NVVDErrcVDMEtcrOPAvxcdancsD03ZaUFa91ZAevPwLV/29d0w4gUv4Ty1jOT
tOGdmVathh2hnx79TJr3G2eubdFfnCpDqOeaQegeYf3WYjp1L8goKzgR7qvIsCdr
bAwZvlwdgOoNhCLkclW40ngm9D28eh+hcb7YyTskSnRgjiuNMB5giUvCkuu5GZIi
xGwT95PaViYK7IZddcGSL0wvJvV85uYpc8lwrPN+612LYQHk0gAi55Qsg5UWM+fv
H99B+qvrNcWsCO8xQFDlwHIEa3IKUC0cheLT9fNNsi4MgUuAa7VB5NWLMJSmiXCw
nuf9od4KOQYQwewBJvSxDh03pD7PNNEGe48K/3OsfAUQcKecCswRvPTz07DXTFeP
J2INuPkhbW+f1UzwYWiN/XqIODQHsm+rfQ+fSimUaYfF/8ahW3D4pdOumyeu6cpz
2ndggeENUqH94I1slxcZL9OUzfRsdtgNToOFS+flyPjEAVAh3+f+mRucIbKBUGKu
uCu/auSAw4qBT8/CLIfv/kaJIZMp/my9iT5zODMbkYMBZaWwVj4IrDXqv8XbCJYH
OCx/8vYCNFKhYfetV/JpjWG0Ou1GFzEJpBFNTfXP8NSNyG/UjpnYqVEVtFYwu/TL
EcYZHQZHF01i4khNnoUAtpTB2nbVL7s+MyNqmPrNIYNSyY46CmvPD2CaQ8eYeJp8
EF4q4dIdc9r7FZIfFNiYONjRQmkcwM74wMle9//mFYCiLAHqjSMzGQB6XgB9IU8S
i1z/WRw3i7V8E9M+PAlbRk1jd2h/NQSULIBhndea2QAaxleca5OMHmPu519lNMq6
xnAhUqFVLhvoXE9Tm4KdZt9KwSppC6LBmeOpbDhTU1Z7JGyQKTOW5XQpaMCNfI7p
9MUM6/sKMIIbbHXW0M6GivzuyHhqVD5WtMeuA7cvrjhgoaH11VRauepBbYnmQ2Su
Lv7u7jps+UKeQlHUWsMBjas68yJl1BT06ljopCSQaPzHZ94455oDqBWHbb0v72Mh
HkfAj+ZHU7kyX7rUL7akYUWxDEjvRusQmdj+V9XuTaQ1yVL1tNmjhEATL3gg2snK
sJfKfrAwxgNkfUIUiGXKO2hB5264n94GSiNCJmxArUgBGGBAvN0giMpNX0UpGxtY
pCRbVYIYXT8HYhw7FFgGMqzKtDP/QU45983qzK6rb8vPJFG2eo2DhdSku2GLXPYS
WqVoPzSRYUg5x6mg1akQv9h1ECk/6vuOzIyBFPFk0Y2rR+o+ymGVW9Mwl2Pr4POA
LJCcis42lDsVsanHiqcYbPLFnFsCgggExZbR7v+86IQ/J72OxfOD2iIUqOKWTdZ+
61qJELEBXHWHJa5kJ7NkYJO6gEWlSJLojkQyGkRYpHxROzEzNi7kkcmnXGO9NLY1
vsDuso1IBJwIqnEJwt3JQCrAICpqS6UOYyq9+NDN2S3rkGLGs88BgipDBrfkSqbg
Jdb9GCYpBT76zjMpiumnl6Ps5NGMHQj18cJfWWKC0NQ/XVdd5gbuXfg0K88VO0Rw
erVh+fGf8/ZJtEE1lLtLNxxMRQJ2IV5ic9e9fkmY/MVuxix69X3ZEtSy0Mx70m82
h7/AzLdD+3e2Tz2io1qGnQdjQyM7t0V7gXmZ5TievKy0tPzDmgqxL8l0pXGCEG2F
P5re7XpQyzg3Q+t+l1rWRQHqycKOqXfpS89rbXw072QJyvvnIwyLkpXmh6Rpedlb
xIeLvcZLyCNquvwTCVrmBWN0ycMH80ys81iFtiVBEiTPKHM+F2PNdWRgJVIN5x7c
/IX19xldnJnUDdWd4DWrqMIMGX3sJDFtahIh0GWjFFbFKbK9QPnWgG9rvRANlww/
sULOMBrFOB3xwW86q2dRqQtyl3iqvHHQfUjYxa/s/mcNqNNofbVi26NSKeiZ+BI+
KpkeyjO5vyqzqpFmF9lgseqsp03cgBg4TW1zI57ZXv/lv4ABHHELI5wEV/zw1Jog
xUfDh77WrjjMq6/vV6tiOA+GNlIcEmPXt39AOpjC4VdgrMt7BgFPYG5MhT2v/B/q
pjPb2jGJVJd2xQeBtDsqzX6sifqDyOjTAEuKxxmSEB7SqvgYT/mFPr6hel7W4UsX
CBwS5pyi7Z7aZAwFLxPB9eMfQH2YNZHbd/6jrvpOpDfXAkx1ulN8faGdmXX+nl7g
UocwyWWIClvIb+e958AVtK+tm6bqQKmJLRIYg9Q8vFk9DBuOAjU/X+DuQrPtXN/P
1OgCftBIDlX93/pbDjyKIh9QQT6uAKp25rGVfVCZlxGbsus2iFRwVI0mC+N5/wRI
yd+lLBlhYc5gZgLhE/yqQf14XqVhVykQJDzKf1s9c7qKpCDky3LvNp7YNUeiTOEI
EF9Lxi+5IKofzd83UH7StugmJgSBBxVJVh9+DCw3Yq9R5u1ifwTqb30ocHSpXHTH
BbptPlq6V82QYq1vyX3Oe253yAdNm4MGOMzkK4wkZire5+bFwDMPVwBDsBnrmBkg
nxoYiLqZjr0tl5NTyK+GRXna+b4Ms8LI3iEKYI/JZ2+gWIcqGg+t1kdg0gn/bYfP
XONxbeupRxZyxYZkxMDlShr4U1GABqzbqU1o1JOR33SNbU7BWTs8wD7mu/nRjrzy
oL1VWgnrgNFBhSr5z/g/CpC9sYwj9OO76gXutms65uDDUJSgui81Yx2o6xDKMwA9
oA+3vF56Al6RMBAMfqKrU6C0kD9pI/ysWu4p5rEIbt56kaEYLBIZiPSLAzDAXb4M
qA3SEY20PgG23q3sBNg5Hg3SZnRt8zF0iYFZqiqq9iGy6oHr+cH71XAkt0hZ5aMD
WPIxAN3r3nOnPA0xmnM1Y86maWyBsdCa7jaV2pt1b9eg/GSoMe2/b/rsQ3dP2gC1
vT4Jbm6+0Y/egJ/9fouSWIuS1Hm9bfbPQxOE/401m/kLQLm1dGO9PkSuA+KKQop0
XkPIG60V7EVPYDQPj2huREW404OWsZVYVV7IeC9Ly8JKxkJdI8Pm6BkGiw1kShd0
LkmUlnDjrcevofj2f5IrK+ez0ZK0zrjISw1M0lO6V2r5xW9uYZ5ODnXYF4sDf95S
WsHdnuLjNQU1t8bHSeEf5Ic+fzO2JbthJp0JKdMuzeEDACUkE5JwERVCPtK8+Rlw
qRQSBhBz6OtgAaBo0+fW5rWWU2RT+5V7oQTLA/c9H/Mu83F4BVTZjS6RVQvt2m/e
LOtDICDJ8MQSdxHVFyMKR/7rVhg6AqBwkJ4P4AU87agBad8VeKbiaxfqqNz+DocL
ex/VNE89VpfOmQe3gd48XP1tcxPyKBfvlJmh1phdG6w5YFSXdeSDCbcyMXB43srU
kfJxerE3VkCjNWOuaG4h/ZxShFeJVuz9Ki+y6y/OypGPlkZaYzC8HQlFohk/Z/rq
OY61/pkZkUwGqVe0YDRbmu7HXcHtXzB4SdDsrT/Ad1M5QvkVOUJwa6VuG3P3JJGt
nJtM83B2P9Jo9M5CeDLvTGkrDFa3NHZ217otAFbneyavu2cu0WBuMWej6GsjNphj
3cxEdramdXMg6Qlo4vyZrBKjwidwRtTAjKCSvPs3puxbUf9SDePTSOJC6RrNQP3a
9NVEkYOGkOxaq/qwP0To6+TVKKuaeSOgR0mH7U9qY63pUnFRddplm6pfSMisPZKM
6+5hODpG8dWhyfiN17zvgjBBbZmVZQ/TWkAAV471rhKk86+PTlHqMl0sxlZwLSit
+k5mldoGr20q4FSRgFZ0KAOaNizJEJyGUdO0sE4KxYPnuvkZY25227Nz5LUHJ9vk
dNsVj70ORY6mGgjOP5pieOmCfZab0wSjsx+m5H71lm8BjgOWyuhbcwMsHIxcZ7rx
3cJQdCrAkSPJxlO6rOpcqDNqSNBXBvbx3hgIjb9UP34tHz2Hztoy4k2sSiiVWUgQ
EFcnp/UUS7nl5JI8H/BL2WxtUzOqC5hqu2BJrfWCWwcakFZrowsDX05q9s0zYctQ
7QFj0cYwWqhkQCYcUB51bI/VzWZebMxy2JfSGrXvqUhJM3HwADBAj0rLu/oGaMw5
DiKS7K2xB+2sppF7+OG0HG0u8Inl4fplpD2HL4eaygW8K4OHZw45D7bcDnowT4H2
uZqWWSxKJELZjLkIaBYqAlA6gCe1EeRs2NMvNGLN1oc/w8Fb0uphk5sjThLGh/Z/
UZ0uC9PtgKeAlTm2ssqXUomBkjyGisxLe8SJO0HCGjPTxPWP06+Y6fSuAaCqwH+c
PQd7Mqr9hlL9V5VLi1TYfSHLoqPqM81HD9JVsh15n59DLf5z/A86Kx/MiwH7ohs9
tYomCVIpL8ALvVzsaNfAWlAuh1euocQ39W9hSUI1zpdIQr+dBa5HFtw+2c9y3j8+
ddZdp9C/O45PXgibpefOTQMipFv3eMO0tncPLAeOwKyRzy9eOWwZehuJZCrMZOoT
u3zxUE7opxuhA9aqIu7Vt0+FDpvOfmGehpym5iUWQVSJXqdAUcpnzeBF9OO2Milu
9hiHGCgCQQczM6jOe86gRq86PpbO2j6pWHLTW+B8+3/v4uPfNhfbfkAVZVVbeK2z
THiAO1s2a/Bc/NBh3Za5nbak6z541kSa2594HczzU+SSqf3LOPozo/rLFyx4xrSp
C90ydTXCfWLopsepwv6/Ru1Vq4+6fE/yl0qRH9j1QDmzNO0xO2jrWhr8ZfTtEXQG
Y2SRP0KwBzHAvdaq49M9nB4URo/849C2r+BsiqBGPopdX2vAZEQZuK7t6dyv8rD3
7WPnNHUVIfKbwHSfKfvumlgdlS4DwVcEV3Z5JkHGNOO4ViUesmDwRXMf1GFQDER0
hhUqsZKejXl6PIihbReB6Fj1H+B2KPydL7VE1Tb3NqgTJrtjKzYoM2SBR88tu6Qu
IurgAEy2dMkYg5W6wZDmXpRYx6jynr6J3N83kK1Prkb4EHmYx7Fhfb5qb27ytdn8
l8vURlH3VV6GzWlPV8HUUPJ9yHBEijbE2tFsnsUgxmkLaLXD84kHLZO5d6aD+J1k
t0wJ6GDL3UPfJb41Mv7Ik40Aiw41dgYy0TxrQcDOPpUPghfZUABOkmj1/bwQ86Vx
aHbAq/xz1GiSAqJ5FWe3dORr227nb7aCV11JcSFEjshyCtqhcN6CNSHCxSq4Qe27
iToVOke/SqXYD4VamMCMmI8MJjDWB608khnDJmHNT5EE9YpF8htyEW/lzis8YR2p
5Gua1xB9prI0tWxiJJGsfg6nmrboRmLXtno9V5+yHp2jWuAprx7Y0CdoldWKFiDL
ALrvgGLlpDCQXD1JA03pmPxylzQ8tRdEGjnfIyWVaTcv/2BymK6uRuFPObT3KBuP
eS7J4v5jW8zcLSZDFcpWyvr99+LM0WDknSreoTdfTd6hspq0mo7CqeZNOpLqOT2a
bSIE4td7Wq9fgGTNY+jn+GXpGJg+t7SY4ruR9nZI3+WvzH7II/6LUW4eIohXItuH
ZvVIkVR5rspLnu+XhPXd7a8KrIaRp1s1K8GSS9EysUlDS8pXGMGmPiNxd8203sNG
lkK5I0thhwu3MYenfmFIj7FbHA7HtkbFD/6OxSnGDof2nbUd1h8ZnxqpFR7erdZS
Li0ZvxBoQl8gePGlF0SwZKEzA+pjaxZPZyZvQIlkXtiVccghsmgJq5WulYzFiazR
Dz7NAJWs2/vL8QlZ1RRs7Kar+OrawKw4ii31B2JyKSaSHW2LOaaXWl1WygzGoKV5
wqv7Hqyi5MCBtuuFIujVYte0m09hK8GtJ84WMLtw//dFKas0JHk+oCACTVE73Hl8
zLs4RYmgGjnQY98ONVb3W7HUunS5GpFuGiPNds4Dx8QFbQS3ixL6ydbUPdsrv8CI
9/COhrXZAdvatMeMkpeKJsi+iLKRXSG3wCbgeGuCRk96xEHZ5wjdWazXoWIe68Nw
lCxe0CGqTKx7BkMPBQ8FD09ln8sdB+APu+lZLGqT8Pcf9lOa8vgPfdmWlWMhMH1P
7snQEioSa11RHd98S34re/ZGL6DrUfucf+9+Di9f5V0fY1P3pA4lHlhfVMf9ajtU
/VohFbIDxRqkkjlSgwb5HhLhnLQKN+iuu/fBIg4Wis9bsL1HJCsdM7PaZ82aRY83
iue5fgyMXUMYtMYoAkFR8HDgO7U9ChdrvQKCSd346mOLLao9zm79EX/OVeyugCL1
yoF7JEQjGlzvGv+OFFjnNb/5q4R67AgXrYLwYkIG22+CcAaCJHrFuux1wwBiUv0+
jVXLMvieXHEc/ZiTCv4Hg2MqKz1PGZFiAtoGm59jxyjwA+rG6BO4uxuqLVfrU67q
LVxK+BdSj0k2vvwQwr0/Xob7hfg0K/VgfrigmONvl72xPlY+8DKlB/fX/8o9R+OT
eB78MOs4uy5vI7QUSkytSzsF9VZUKo/cgG78PRJc2S+iGQfvGkUVwpTBKxlfYo34
5Q7d+pvcMLQ6YVdFHONJz2KgN5BqdoSKp5cYoT0bENLOqMwKtHjEi5Kh9gtfgHvg
pyQ6fLwQ/dLwZzjYo6MwPk++acE5fdm5ztGVT4wW6g2AVxAAeuuB+bMmKvdmOCkR
2Z4rHTZnBOOUklXVg8XqAYSiyAwCytQU2Ql3TZsu0t60WpHBwlGDGrQU/1TOFTMY
eJLIWWDUG6p2JCSrfVitCe4C8Zf14Lx+KuRDmWWs1LE7ouUXRbBfGvO4mGpyPuKI
2QsIxvBH1Rm+IgGCfGaxJCWqNUOWEFShcW9DnTNGRPxYPqOcFiIlcisg+MyNeoDD
g4W9HkLiWkiRlPdlL52xN0x/Eh/b7WeLVZ0lzczD0Mkwd1KaXzn7zcfAGZl4KiPG
p6asmayRf0Z4bAJ6i1+/vHcJHHN19mVUrIC7cMyeQcrtOqd6bnFN/bWmg5FpqQU2
sONSMD5Ognldb+T3ooLXWpM/dfmtoZtbyKlpLmK0c31ROnQGeB5lzF+BOVf5bqXK
oLJWQ4En4rmpj53iN5PcLpjMzHOhj2i+7TIFP12xKDyJSn4RyvVe7U2mwxfbS7Oq
MpeSeZSx8iXT3fNynk8CwPlelnvmYqTK7mRsGlcC7+MmohvGJ5PHR0OL6VwDqBA2
GfMnNuEIvYTdfGJGWud2NavhLSj/GVErru/IpXZrkkBq28v19L5sE062/MPkkaCk
2kTljM3WnZinP5awo4ep08lBG3EfGeDlMfYyxvGLV5FCTYUt7IFeL3eltKyxNsls
be23IeNQYEY93RibLpa4wO8NcP4J4MP8Wm9aTBNL7ihPczxM8SNUwx7/hJaA3nr8
3CeS07SUKbaqVNTQfr8MguwOK4m2xAMWOeNAf9Ea0vMQ6g+yYVwC2hhk4fLFHh0U
YTN0/Lh2zjjEOm2+aELUee42fyLXYAzIelgK7oHiV8qqnfXJLvcIEOFvAOTBDnpE
wVZgdauWccRMl1gvgckOXRlesdngv6FWEN5qHXgSJnT2mhWtHr0WmGvtbZWtV4z/
arIHNvyiXlwaREbai5Dgkvu77kiqfwtOnhYM2Cr4HD9M7T4ieAbzc+uz3d6lkfnc
uyKVy8LIBqWjxwV5a7tf5yGEdxP0bNRrwX1mxJYCE9SnjSaD4OJ4HecgehoCHhFG
xgjfdK3AtlWeN8yejE5WlZ3ul6oyJw5NC/om4r5X+TLBVmXHg1if2hrlbR3j1RwB
2WJjIgqDZTsoR1Ao4IJy6DaqpP5xETKug5H6GjkEX/flQJaIF/09RMBRSQFCAkQe
UpRzR81zB9cJfmLqMS+ZeIBjnebVPPGVuZg662Mimo9tx8SDDj/XietoJP7Vm0lf
Uiv9iek8nHodi6s/HB25vCxEXt7Ec08rW9Lbr+lDXux8pZjKvJabZp421EqHHhF+
ukBQVNoWA/7nZFPgPkvvULxjLkq+BF4yP7mBpRqbBeBREkaPL8so1wBlmghjYf09
ZSJl04ziKZ4XfrS39HjrS9HEiJh4h7LVQJ2GRDHCnZFFgcK7R+zES/x+7i0tyGyi
C4GMFiFJiWNTV95q1wxIyX8jBOWyPZAhvEhrJawi8i8mnWgraP5AzP1jc5LIN26j
2ZA7G8jLolVQCSL5tJav+Wd49556bAKc1MDSRYKcsr7WqhadSxOa46nrU2QBAZGp
p4PXEaz6VZ+jlvtQwRVwhD12n2umd8U+H8LlM+FGpN80lyhK6i1YLH6vJei4d1+n
vZty+pOB0sOeKcsgJ7eCHRyvDY7pkFDw6S8VCWaqn4PIQVpKgvZNEvCxU5Q7xF53
5knWoYAD+bQrJveJ+HzGQkQ1sHRvt2qQ1ZjKH6HvF4yKWSQwMaG7YyLPoI/5OdKX
DNcvY4HJ33W2fEnkGLauNgh4feWkCFKZNdrd0JyOp1k/C4XuFBfBurc6DzLpzXFf
0jU9TMyGZ6CVw+gCbVl5LoKIOxlM+jXiPUmbCWvdSjS2EC4dp6ZCtJJdcpp4H0Zz
obt1ZtfOkMh7NjCc6tdRZ2n2FFvHsimChn1V8M/bq+qFeWyolnzULLsQpHIan12H
GUoHLS8wNdUzBje/O1ABzlFbDLpIUTw1KrKHU9cMOxWAhNpA5/QpSMZpxmnMZx01
H4kl5FE9q7ydqHhqgDu80LJyhQsvaGZuGs6cG8qNW9CA6Ra//wi7XaTgwUBSlDrL
7/ArHDEVlxf14vwGo4iORJrLtmNQRkhxhpL6jxWc7ssWe+swzeRJXDQiAkVsTjq6
aMybbHZnBIZm6JmxPNWAPduDKLoDXnHrg4wFpUckzQ5badc1opnW8LROj8/CzZBz
MLS2Zz3R7olujT2nAlxHSNC1TIJMfzSCQUcvgP3bSvwUHlgPBSHtp1S06NAQjIDt
+Qe3+GL1F4B56F365umRl9Om65Wc60nltSpZSwR6yct1sMtOMioFMgkoF/SWMr8m
/ZSD/6DCNUPCSlLOpC6jqmJNWmsU5DnWYHk6ZYWYQhBcxth7pSaDYMKqV0GboSbU
ts5MajDn/vqdfDWdRW8E5sJHCDJ1923SF/gPOs7KEYPsKHapY7Rqy05jncxvjU7/
05JqdWc4iRPQlWTbDcJvfU8ovjQtWJ5mM5uqSAZ+sEGh9j6U91cV/joP+0qjpEKL
5QgWaP1h3frOn4pJ0f9JGUThjC8kLBwr6NmWpvOyljluKIIKCWbaZn5y3Lvr7PVE
nGiWghwHq8MS7NYufePhRtizbkvrCaC8FDDh0VL/B0NPhuXO/TQP+gTw4Zho8n55
fatkpg0bEpRyF2Hoxshr2arL3UlctbawKK2GKbHUbSvvG5yB7b1gq5DUlMPR3xYl
vHzjV49aAUJeJe/+RO/VeRYiVJkf4ctEPj9xFE5IPsEtRsdR1HOCmKu94X1blBln
9zZ2swUr3K+UOXc7MdKjFTMHpsEzFyxXh4gPC1DK2KXyAjGKCvq9vpEBobPQv/6r
BvopurloyK1HKc/tZEgW7uuF1SN/wFpaOOr2OPvyMDCiLLk7jId5GmWuJyo+4uoH
pp4UZSi+b1B7sCAc+WJb1XJ0OTHyW6gmhEmZeJ4hAGWLmwMB6yyEmUfh+Byzh8Ke
Uy/WWcTCUc/nW6JJY7lBzKYMYNhLQZSCxS0seTD0KNa25mgwcEKsmI93q3tQyTix
opdO5WTjGtczS3JIR7J/zIFi6wIqT+rUsYnTCft5nJr/fxce3ChySILjq8HfPYCp
/e2iDUhfA+Q8vjCvXhrYHiRzaYsUcFjG6rnoT9Qk1CPj562vZlDRPZt5o1zpE/0n
0DdUiNL9FdWspyJHb5IsnI+DEhhJapKRkkIwDLBza1VcAo2twERPaT/CohPprXbk
Mw3WYq+E/4M6IqrkUQ1wTSV5fftVTFkAZ7YOjFqvd5JCpaKc0d70KdTcTqD2vR/P
OsvzZap1gKypWd95T+vmARkTHM6IxVm/czrEja8dEOJlsggdIJ0YxLPaNdDNr8SD
ZcV1/qtNqAqrADWdRoaSRW/GUF8AC8Zmb0SBIV7H8CcYZyYcdDfNCIcK+6YwGKjG
iDh0lLvJdv53DkSoYm/SZa9QrTDXvfrhFseAUMJHu2bSgckYEYSJIZd/ACknh2Uq
46ZU+YVzsyuYhhXt5pJ/bINZncVM4GUpE/1Mrbq6eRxqVtmVwTBPQ8dWjIkZ0f9T
lMneaZeoO7ulbMbbkz9iLolSJTv4J6I1nH7+9t71K/moHaHgNKN/rnzlv5cWV4lp
3LVOmkv5LTZwTAG9k8tLHTuoBn0q0HnzlrM1hZAspd13fKES9Mj7fLOeu5zU3uRX
+DLfOBWp33iUuOwo3Vvvs++8s58Oat5ubRMqcC/xXr847UxnQM+DEUY9y1cxC2tR
/TQRFIdP6c4rYsB7Apm9TIC9Ko2qahw+keWTr+yitpRkMAQjL+ojWSfA1JmrOjd5
1rr6TlKGXkJXQgDZRN9e/FMAC1iioxJUFvHVJVnw61rF+cDxmRxOEUXHwxkQ98e0
TTJFozCBzuHjgNa3mm/8/NtYTUZBlxBVlq5Ik14EfuGDOQ8ppbifBLoK2UvEh0JM
dxh/hqY/B2JKNq+V47hWLc0pH53KCmQx0/8aAUqCoPjgOhWw0pbp+VMaGUZuTpTx
XOQoxkBPtQvAEcg4bCByBsdyFQ8HkE0Tw2F9WzUrmTAXWLjBx2Mxjprc1Z73yhh+
93lK7/fkFiCQaWi99u38ovb+LGksgnccK7+i8lmUrGrMShhE8LhRUKGEODKg6Eyk
/b0fHmvYVgtdbCxgweIFomgDVoEMlTfMblh12+0iI3cBN8zM1E9tq4/WMEf8SqKF
hsOCGvFmCphC9S4Y55Ajkq98XAN/4DlIY1BPnnYq+niv16FI5K9jrJGHbmkKjg0W
QRs2MctKRFNOTZH4wzqNTaIqsFilkON2u7OwTSfmAeGKnuFbo0lBWA1eNae2rrce
nM4XL+I11Yz4LteyHWYZpvpSbvZxdALET7ugsAQ7/JL4Vzqg4x4fH7SYUHws/jtD
00om5ZUxyFj265VQ020WOgJu/FXxMwd8MUs7qQIg3V8D3L4JKKhhXpbjW41gdrq4
CZ7kSJ1PPSuYmC+a+akl792AudBaJRvjJX62G9EwApwjzXwr9pAhCXcnWKpUNHD8
ji2Zo04O4bA+PwHYJh0htUZd9OPb3291S9egwxt5BmlMMGLaDNqY1T8uTVSXDSTR
7ZL/RllE0Ise5tfs4u4PSwMZ6SOi0s0AJ9N3Q/Pj9eK0Dp8WhcqFw+g8KObKHwe+
wSy5M83aw5+IozvSteedl1YoTDx9/RUdo3WKxGOWrATgB+OwOiV1v5c9QXWFtSB1
XJS/dz8zNdUdeY4zyIl++rSGIKe18yCJqidsUvi3gTtxgysw5POK9HqcQEG8K/b7
BKLxPetpzZPP3NXtlmDn6Y2M2UfJ2qzb7iilIaBWL9mqHLBZ0rTnobt5gMO9jmIe
LtbuiDyMMZsXDw2UGxfU4D3X9nvcdTCWyK+cMZKdoJ5ATopDTta4UczGVYEEt+J8
CAZHecpl3H4ShiVcoa7ifIm1m101cuiWbJmN1e3dG1cj1iPnLVaff8Srr7SAJBOM
oX+NyNBnoi+O6tsBe1KEVovP/S3daQe5xInSiguMpOyTxMprgxH184g/PuaDanRo
lgyQaCWRS3QIzjXKX5siOKvWVy6GkdCef5E2H9nLWm4Q4QGVN1b2X2Lx7buwg40b
JWGlnnwLYaVUvV4ouQPH/UoFvP8B+N1HrN+w17/C+pnM4Tx9r2yxp2mnrLzqQFHn
PJYGRndLPcXn2X7BQ+jyzWJBYAfExYP+6eiDsdBgW4PyQl4R5J+npT+ZAyC8Qjc2
8yBP2PBBv7eHjXc0hpfkqyP6XcoaWdrK9ABPOQbTRapFce5C5CqVuuFVB4Q9dI1u
pNNGyhBNnY6dS+r1puxSoBEl42U3zqNzbYpVXiB8yL3OKBDRYQbihKb7jQLPFFPQ
U5hjoAnLxB2L2qjHZs/Mx2+70zLnAa5FHb5JcI3yHaDqm3pcm9tA5RFCzdEtgEet
NtZfHDmXK110WzPk3PngSDJ21wZ4OSWJ9ulBWfzEZLjyWaR6KLY3vJGARZQiza2/
RUT6/nkAuGhiWKz2c7flzRMP0Ix0mZRkNCebr1GmcG1JL09oE+SN2aNGH2NVwSAo
te1rCpnEO8hkkqkUbUEU7rI6vRIievAebD1PyWKpT+8og8GoBLFcqHRLzL0ofcy3
m+ZmGPwYazah5PjFGz1lGnUhKYMsXVfyIMXHGhJcVejvi3yG8xZY4hM/6F/gk+eL
DoZCZC1pKenaw+Ou9y2EAv6SAgxh0/TNpE5m5cMdFyJfzOya+mSGn7j9jYiBmhLJ
Z+a6HwNgB/6ScGQd4Nk8qH+9LRh7sqHKrjU7EXHpsGUeU2M8ADnGgVt4m25pDkLm
+pllyhrzLx4U3QGbIZ9T9F5yvrvFAg1hVZSPdYAN6RSYYilxLhL1hZl+sERVBPoO
5eBJeevFWbrJBtozW5bVqaa/hxo4E0N9AP3QuyAHRMO6A5raqPYZMGaonlI6anNU
ZDS8eT2gO5GOCucr73jDgk0b3Msxlth0APQDBDFsu+ZX0CGGSF66JuiQlSQ/pTql
w0C92zkTfznvYIdgoDO0gxxHinlwy21nhJ7/AZWRSMwDGp6Hz5+o9QDZa+7XQaM+
kOj9PPfB6JCSsv2yCZvK8cLV1GO5GRcQF3DVb2x8EeYegpMUr1tf097+YpW6qI6a
6mnd5WUZStLmyLZhWp2uRsB+xdRMjm8MZqm0KN3TlpZIhU8zF70+jNf3Q1Qm8qNz
qvWeS1cnkJaj3CWcjXeSc1VtMhgtdttSiKvmf9aciihzbrppk/HAzXiZ8d7H1dIJ
eZASmjk5EWpOYKL8ZXczZvUuUQt3tlnEZWnuvx4dUKgEYAKqGAUbzbMSg9A2qFEZ
X0TIDO7WxC1SAhD2NfanoFHyqM5pwnIHshSeyXg2IsrdmdBXzA0WWHipu/VCXF2T
HpTz4J1Tu2fcz8hgELN782n28bZIFazKA1dCMm40yxPqxvSmVVUxNBUN0yiphB4q
54h9qwQ6eu8mqXq+r0WFnjEwYL/n7m9oXpOPapFTzRRe/KcMUIt3RJw3DGcw3oNO
e28yBPG4+k5kd//WPu7QAt7+7/3OiqsAL3D2r3P6YDL3u1Q8ss4lp3wSxevY93ea
Uv/Dh/xlzLgW5G9aFHfYUzK9w1JKo3MmgC7bj5RW09S1UcGvFIv3eVm4nTTb08cD
URjOYClOlSdaawlTGQG7jvPJe18HkPv+oJeGLLIX+zYmWBjYVQFHrMiTERYuOYr+
PJDJbiPHtqzw7JY777L0XewcjNB+Fyb1Uk6LEGOeZftOtcjCTlL2eHGmGAmRo+TD
1JmXpxbmy9jnJ+2kRKwSdu0pjRHRo5p4dXhWpuM9+imFQfkGYI3xROvQCGNie3vm
XyomT8xTJQy/8lCHGXFeQuhwVx235rlwGME228NsLuDgt6YteB76MUnF4R7nGhdw
uQFfNXIUa19wYJSr+2g1skT7g49vk/z5zefcjmGKLXmC22j6ZVrB/2ikgBiWhU6o
oqi597/t+TbiQgxJmeWhXOYnhw6j97UO9nCBWrCh16Nbr5Gf2XR8VnjIN0tVcpvw
iEvlZJjJNYadG76fyxVNBtTBmKwfJJZehu7S5izpXXGcLjKOb7bXJPrWkwEaJjcC
qOEJT8+u0I7AZIFU7rYy925TRH4lGCC4n0YiZKIHEkIKsckhGyyrKXM6yPo6DWY8
ak4Oj3Z3yxGleBn9VVaH3bD3A7qKBpCoKtTQQG8l/dtokPAmYOOoy80aNNtb9l2F
LZ08R26bLhvMsHmIjjFw/QBqZvAr6GSU3GIf+K8fqXxf/ERXLsAOwTqXeO/F8Ezf
qzW03xmRVdEtyqYgPabXi3oy1v+9XivgIJ5GlNaliFArgfip+JztbW5o+nqQOOgn
JykJH3htfruxJOcSLKYKWZ0k+NX9tfEVwM5JwY5IlNm1uje5k5NAG6SqacjRdU6R
HBJ7lPfVHxRxOGhP0UDZLuqjw2Jh5YDAh4KpBFG7sTWD9iicUV9EWKS+1XnHw1ce
BezkpTXGCKsIw3IyCt/gh+NVjBF44VIDt/7nS6Bq/2l934WJBkhUWP7EMfisU1Qy
RiRV5N6EiXGpX2G020FNqFGwmnFCOMtWsVK5XuSV5lXgfDphiMSTfL9jUa/d1DkH
fId7E2IPJKtda5lykSyX+rBATvzKCvI5UBbx0Lk4b8LdUj9uUdZ1fqlIIvBTlrUU
Xx5i1AahKE2MHbSgX8b1RITtSqPQWP/oHTXz8DqRDcbTTAMrWnuwPjWDoajANHMu
+UKqNKS4Us572i0BHfWZzHF8nFTIkFNkjJaOFoGVqzw0uQH8WM/yK88vrmVspywV
4KjSdDXPveEmfJjMKIP8CmIrkAQm7yhfHMxlOnSe6McETL/9zViKEbdKPzKacDtx
uCThquvJiZhUtvRJ2lfefs5nwm94PtvoKAUpBn2ag6qbg5O4MAU16bcxq5lS5jQ2
4Ntgk/ebAxFh0KcYpvtNxGD1QA9yH6fD8vRhcztpiCMjQcfvIPGeGMh8QO/uZjDp
0qwau0Umew5bPXf79x9yNP1oxRelIoWmXBVSGhcB7SuN5fXb79Pm3DSZJR1dyOIw
wXGugTvJADcPFfiNiPGxot1kHvnDM+vxaROFKHVAcPnMkBQcoZ1NQmbDLTZFcdkt
SjKx0wKBdC7lULzr9BmVZRVnUjQ0o9CH35sA0aSCNDnxj14UQ7PzQ/MFnPlVkuit
jCLW0EdMnILEdDxZhwhRdv76RQWM7EnGXPyTlk5fzJ4I80unHqtHTiH7S+6FUfkr
CrA5kkMgoCDa5yQuWGUmi1CCy9utOqf8oe27ruyMj/PKSabgwIqjEaD/y4/CnSPH
E5YgK4ETEzvLq8Wz/6cBRkWymwXDGrd0rBfIFsZzvHtr40enmqsy8z8HvXq5XbfZ
Sm0WUBKwP+BhMztC7hHLrR6cMjlt7x5a+CzOaQLW6X8ua6rEOTaWFui82O3ygoaX
9FZPPS/GtxPxTHdPq/sfACPM0G0tW3LXkJLnn0BbumBLxDuv2tRv7OyirLpykIZU
wqV4jxbVy0aRE0ouim44FyjEbvKSRfqBZ5a1VLpBFGzv2YzECqawLLk5Ppfox6mo
w3xJSPj0Uy7BWI0zc2sb8HzzEi56VQTgCxz6XYahyAaKriD+SWj/Jc9L481N8wc6
s3UO6SF34xlsg3AUvkVqXWT+MHw21xgwKXp5dV7+FB8a69atbpbuiBDyH0tBoJBa
91ir6GBa2SztuFfgT268MTpFeYRr//TJDdwB1nLz3C3m7R2roBRqtV76RJMKd+lL
k29h/PFDDmL/DXbqt/lnKwomytE0SqnAYc3ZUrP4EipOzPErOKYwipz/JUGSmxsz
/F/I3Y39Ry+FoWItlnzJ6HsWIczakzY/3F2QXAQoXJYS85RLeatDJXdHQc+qtSFE
Kxul6mzmi0hNnJRGPqAkvk5S+WxRfSbSWalHHMzSnL2Cfq8WYlptElNJdZfqo35Z
XTOPLfTeRVreoDFJBss4FoiDBupNnpTh16JVBLykPPFPFIATrrI+KBAmLcSelBPJ
qepfeK01GwsyhwTiWdEvLO0NTYDuUyGkF6oCkUiOVMjNvfip4xcoUm9+I4j30D4i
EDRQDBEok5R6v9TzE7d5VWwg2CtX/sqXXNDy+/Ykv7H30/UZV9GP+lLm3rdE1WD4
DoVrmV5Ab2vfnXePd+cLSI0LoJ13gQxs3fZlhJt0s+/1IVu7KbbNDiT6fwekME8s
tsuHjmcmYKQxZpF4CD1TN2osNrteGDfQggzGQEry13s3jRotE2BxxaZp5nA3dTln
fml2R+9rhxPA55f+JRrzNOy087sRtBsWBEk5gnvtVNKKuTFlOXxNQQRcCHN3cGg8
gyjCkpjwQjlBuYnCzUQ+EiqxZpfj4GiDkG1RQIFM8YfyjdNoFfjtqh7GHLdZuXTS
y0UXbsN0GtE0BVACLXYTd8zvBbcjKnaOl6mIAI3wl6yVYy+3wXTfGPmYL+jAZxUU
UY5GaBBGyT3NHCEoZSoMFzUy148QNfmwGsuIi4UMoZNMNiNKXFVm3LVlnvu14wwO
fQnkyjbYcDV6utFiQDtONxON0jBsCY7y6bUWlkrTtQiU7/JEvibiRza+KrmJO0Hk
FKpoP7UN1I1ejo4FlPM0ClW6gy3Iw8UWrmFx1Cj/cOqi5gFKxV2QiEtafjd8tHbi
e7gmeKKWZuv9/dot3cW98MHg/NO3YozhsikR/JWaTrWSfDNp7KQ1K+uXlHyNc149
F94s2+fKZ8f8XorJHyYlLpLMJlOsQHfLFbUzTajwMiF7Wo9kMjs8NYvPjb5sjRi0
J6rGLEHGoc81o6R+8tNOnM4wddaP26OGgxDwfeNW5oSyt33uUwNXiEoGFsyIhYex
pZSk44J0S9DIGK/6wOx0focuULiEQYluygoAG3rah8SXz2vZx5jxJtOK0jIsEZn6
/YaUrCp2XWaqJHuK0VGpXyChoLiRzUcmC81DDCtOf/CHTDxFY7Lzi2qfBUxDoT/q
fDAu9e45ZNn1Ho0S2OY3LLYvHFpXgC4o60pyOD9btBVKtmUFRvVn7E3Ob1XS3zxc
cBC09wTPRmkzWaJyCiXFdFG8Bea3ntx9i8t3JH3XMCXhBRpY2/lNanwKjdGobVCT
EdzbXwPvtmGD7aOrS/FSPZ+jMuWAyvWdanGrkSbJ0DQEb35jCBqy+7pafgODPFsb
toN+H0/baxxm99IKRfuN1WfLSuhQaXVpuIdeRTJIRhnYpOFm3hpMNAfYudH0Jchu
4cQHvXjtW320yInRhH8KQOJdRWpMm7Qg0g84YflE6q21jngNDNO+wUvb/A6Y120K
fjnAIT4M45EqAw9jzd4qgqXOpkIKHV6CoqXdxJ+UY+9lxtyY/w1+g/bTOlJuGeGy
RqHOnEtkdgsXWk9HXoN7KLfIpqBohd+cj+vIR4yCdTHypJK+31zk3Ypi3I/4TK2B
zoQHS3UNR+63ke/eiMZjonI0f8oGWS3QAfSYAzZleVlRhLDA7Df7bE9VQU/TXZ/Q
JQ4KQilB7YCwspGJ0hkm3FliKH72Q+ykO3I9GkOnWXkcdFpQkCenqGAz5uwHPaYL
fSbw5hSM4eBfmFzs89aOkEEiIJSzp69yytZ5374Sqe1jlxC102A3E7GQPuRG29/3
9sWZBeWFSy6nySR9Hun54YKtNgmP53XtJX2ZxCedlLjDH85f+h/Tni0GQdgyBKDY
KEQWTb7AJ6JWWg3Lh8zAJrBJESMRfBlSUQ3ticfLyVz3WkT72sU9Huqh2hyGYMni
H90vowaL1Jb2UqsfwGw77JLITk5Pq+WaoSPpIbxYpJnqaeJZrVRi+L8mIWJGW35T
jgL3pe3wLFVoUX0Uib3HEy4vRvpd7hylCWrm8atjtYNPnwzM30dJD2j7jzSBTRVs
btmFIAlV7SFMC/gSnsL+VFE6SBZKd7RYBRtHPkvqDgwfyxS+xAblqFF+FPU6OdfZ
fv0SgM8Mb9W8dF41CXBqBNMvI0rXGbQG12L3L1nx5jMoCiDU+thEM2WYrj950Ezl
Rdg44sMS19/pXD+vCUqZUvWEvuKpjQniEeyNbBDFgPCBfYQT5JP/RhDyNv3L0SuV
5AGrIp3K1SevpCYRFHDyMwBp95Ph3fCxnuMYnqSsjJgVRf7STtrpSEmX7nLevsqm
eyxn6iqFgB90M2bGl6IIzoGVs0rKF2/DWb0bobXhqFt/zOP7AWO6B+NBQW6kFB8h
k6ZBTqLbGK+0vsh8AGGqbup+K5Ilpdh7g/3NhGz5H8MfxZjzFwEc/0wmDo9WdWvZ
cxtsvadvUzkuOWh6ZszSePs5iYWuoMiVp6wNtHCQ5eb4y9vRJFXklvS74G3/T8cD
nSRhjbTvhBdq+HAalg0o78ihr44oRBr5pKHNklmYNjnEFJdsVaFm4gw9/8FbWKxh
7a8q+OIRloaO/nUPGTIorS9sagRchU5XxloYRCr0BP0yeQK2Zj3LIiZ9Y5GV0ykn
UFyRUHr2LjyVvld/Z+8hr7Ex7q84tW4qLMEcEhJM/+P/hchhlihTn+uC4TvijNm7
wSu446oBuO0IAmQuVL0dKJ7yGVkW48oLBpEaum0xBkAp3zeZxX4GFs1MWJA+wssZ
lJHHtm1wkmP5Rl3QioAHxDNjbxqhKCmfsMVLlDn1wgx5q8qjTYFgr7VXAsNX5uGJ
Elm299p8Ku3WRf8UZXAgigYQTOOmgUN5EeyJBgD7cYdN4lofLuBjUozR8AOXyC6J
6Il4XS8qLiNY490U07CRoKUx9qutm815Xe7iAX2nBKweG3hWlp27pfj9WnoktqKD
rCW/YrbQzX5qZk/3PzUdqyJ+zzMWs5tnBBhIvgZyRu+Ac8fxrWaw0qPOgCMTk3WD
sHCQkH+A9arYIHh+ool+TjBqzoQW9nSLQK/P++eawATDPEzgYmM/BItneFqIrLRH
5a+Dh+4BDHzLICj3n7qtEQBVqsHkb9XFoY8w4WxBZ/tazAxOUD1SZ8Qc6WRe5LZ3
9Cf1/h1IuI5sYyLw0J2jN96SOTmMTAMuovUWmch1gkCWlRsQipaYN0ZAj4l5Hxzz
7Rg1zxeyC9YvQU4NCu1LhDEIs6RuAXeU1ca6zu0eyLHFOTjCjLmcuNvGOReUjVxL
DjtfXm8GQa3BoouAYycCrxss8RPu+7VoT8zImL8NZfXhxxUKLCD7yid4JLHJjrkO
ZjcLXo3bL8JCFFJrqD/A1Do5naAqoXcp2mzr144J3MjPEWriF7Aye4E3cYpmBVx6
dcyFvzq9R4zK9ILM4QnXNK/axL926OEtZ6qL8negRuyxt6j7hTQavXaj6BLr2yGP
fyPAI6AVO1qAClsJoZV3la6lc82SJ21YWGnXPe2/6e5cVEnf9HXaoVuZbdBS6yAu
kmo4Bld99WX90c2TYzkt3SH5sXXaOy0QreDasu/GgVOR4B5Lr9jHOv6XWsrN8VUz
lp4T6HjbononMt9jPFH0tmfyN0S1Z/mG/V1a6dKK41kt+vVmqaDg/5ZPVtQuRelz
76VAvtgeA0iuSd+aa/+jOYsmKdu7dIFkqnURtRdTzrS88sQKtxHNAIaTOe6w/VXP
sNntWlFuEeKz7aWYV5JnJM+8jiXJ47iGQTOKF/tO/7qdlacxzOd6Dncz+XYq3j0W
qCqtS+FfsreR6K7h1cXka+0kj6ftW3hDoSRyz0ynnsUqNmoERFuo2u4lsWY++IWR
gvPc2GrBSd4F/7vBI7IsvV3EHqB+faAER1Ry58SwK1LRsVf7qjZo5WSMQYnqAsBw
A6NKvf7fsG75jwRXGU7UD7wfxdM9hEUqoMmn23mbhzQFd32Ouedagq3xzySjklPA
kzGhjU5Getv7qvdu5f+3MvGyAXrJmIMuqccW9ptxx96MfdpE3kVLSUOvb5U4ZAb9
wInKaUODfwal9sqeDCFkSUpXvC8HovsfRae18yVF+ONI7VwwTXT+1oGzcduF1xFC
C1OvnHoQbIsukTgw7e82sXsAByCXgnoxhETYm8rWvFXbUe9XNtyyR7pHYjXTZyYp
eeh19vSqr1F3Z0+6tSNvkDIVz3OH1HrG8FsU/25dcmICElrMmdGIg6jz43nDFy69
09eA6ktESTWQnMZJnYbg0ZLHZarnafm9/UVozByo1hKTYeg2g498zuXyOimh/ymM
JFh1OYAMQJrBSCGinI2py9vHkj8cNgsj3pWOL/ewVNPYN2Dt3GKy/8deR3Ud134Y
/DOXnw1cYtpJv1jeGvZ/RSpsjeksx+iJTPVUFkgRTQ3aHdtrW3sMSmF00C8enKJg
FEaBovW6KZV0eSxkPZXPrchRGPPcn190F5AopignfTcKDF4Dzdqk8pDL5qdHKVrt
WGEyOwIGf1HGyc/HMsQ8dzLDT1dIdfgg404D3cmHnQScBW0HO+CG0oNHag7p7ZWW
4pY1hOx6iTPWeonzxiHjeRAksw59AY1TYhiYb3Ndb0AwnQ/eIAm3mC6oLeuPIGiq
qGwjIfAey0e1MX8FSr0AlryRVb0H7QZaHFNqIImCXvAOTSlsmThHLqeXHeOs2XPe
jbPjAGQsOagPbkU3hVeFxBjyf820mVR5gt8/scuUMpMA0e9D2/a4Kkn25sYMj/fj
Px6RedHnvpzuChscG82z+igGXGpZvkkxexSoOdoPM3hsUBnLqlWMVaQB3b3fDxq8
SinRmUHxNcvILkK7AvCgOtfqKHQh8rjeD2j7iwjG+ormUkl8Wx8iWZzF06CpFazo
hrmwYT/lRtL4ceK9ZkoK8SNPLdqfsgTNx/ukWPO2tlg6tRZkVb4UNSQo6N7VLteV
zuBvGbW+GmFp4Yld01N2nShHQ/PW4jEdfaATWNsD8JZ1vRx7OvB2fygCV2y/IVre
46h9p/3ZPiUCKhtb3Df2TP32WjL71lJspJU6bVn46MZfEVFVUDwRw5VYO2/pl85e
SD7qdH/McoGxLfNiotRhiJ2t/DKBdxuSfbdTp613najYIrdUx4evclSOV+EGjGyF
cXBBJTkeZho4SGsus/wQM7lo/WnjtH+NW+yxm9KN8tX3K14O+dz8kM7E2Tiyv8Ss
QZ89D6RxmXmNE2oS+yqL3/9F8nPCmKjmykPjEg2jR4OqdTNl+1rThIJWx+3HmA6Q
IfY2RRT5ay9WYOHxPxe3VWEOuaZAlZopcQZdWZmosMwp7yPCwtvhxMKi+IQjoWO4
jNLMULteLQJs5D136D8J50jUXHDnuX+CBu8tPeXLkGmI/iGEnRVv02qlMlC2AzBF
pVo2PTMFyzXIQKwU+ytd9HKjA95OoaUInQmAJSWBYAG98fEbsxeKi7vhcVfFCtvZ
d/obo7BKuAd5Z13JWqj18zL1HBHycx434zT+sW/P2s0myINwbIuD35aAasQrJ3ks
AN1bjSEMTGSb2KFz6H0exTTXaPuXisoHh+Fg/Uuyp6yUKB7MRb5X/a9+rN/f6ryJ
Kq4MRSBQnwyP6x3NwU9HJnQY6ebiC+vCxMWJDqrpoobncOp0xiTcvtNGC1rbqd7p
JXCznPbRgDbHsBt44N7qfQiRPJKSSVXUPLly2xDhiU6mQQ8uMWUwydU0hAtsVlHt
W1dIxv6cvBhdRIEkeHy0d/oDNqKhNfR1ioQv5hEFgNsqJdnlWhBRJA9ad07xYAhm
df/qd8zlhmTQZP25c6GgyWZIBVUEjUL2/g/VwKPsRvIJdOncHagfVRsNnMcJklCg
dxWzv6h3Q/EQ607VPBVL0HMU0LQT31SG4EESPz74NSfbeyHedtbokYRkS/GOiQNn
PLIb6qTHgrWEoTC9ofr9JlSyCSBTXs1AfqNffg9I+WmFQsmhTbVdlBbkRk82kzkY
qWuE2C7EXZnrne3oubH47vtJjNRxiHww9Luzwr7xEOWEN2aODd/Dhek6TVcYnst/
Uv2yL5PNDv57sZa1mLI9CX3kwUstWp3/RzeODE6C071mSyH38x2qKQtFIyK67X3O
A/SZHlCgfEw2piewfbcxSzhLB6mdxf/jMAIkjIeylx9GyMbh+2jcuQ1IOzkCdrwV
w2aKlZeiQWZPAZrsA1P8ceVcT5qYs1nAoehzz8yzN9E7lzEbLrm2JH2ipFJInSsm
OcP5lqAqDYyidC+cCNkkV2kozq/ysBZk7nxhBzlpEB5++kq4N4CkT8Ml7GxLTX5G
GNg+niQLwYwSp7CGMyHFfRskObTyki0OHqDWNjnAN0xRWANTV0wf8QKhjPN20+Y3
E2xcGnbmcO6ai0B8j5sllMD4sRxXjtk4Q8heKtd/vOnIxvAvKuR9PYsj7YcZA6RA
vUl/nELwKYa+HaYQaZLaBWWAihbAq6/jWu8yp5eiNZ7Mr83O8p9du2aJI5+b56Az
yHrcv9cPyrUW4BuuGyxxhVHJ2u9hoUGDXE5dQNivaoMmeT5qZsL891mYcQBD2dho
Zb1T1Zi6pAd7k2EaF5384LsYRvCzf5CK5jpLW4tBvO/J52a6B6enetrfWgkunbyB
wtNS2wYqLNsl5aQQrxEH2vLGkiHucb6JQ2nfDXycafgxeBRMNz8/qi7mw4NlrW+t
CMi64vm8IKzyTkJP1d1qGpfUVyGRjceb6giss33EG2de1PRMe/akMX67IqJraKPm
Ur5KwSzgwcL87z+lqfRYWIJT09v3Awbb3Io2WAnnMoSPGPViyVjVB8e9UJKE2N73
5YeQynGGvgQ7vC1N56eRcon7FDIx5yDB5i+Zltt+7LqxrhP1U9WNqANrhxADx5VD
BdhVHSxeiYraq7Iy/BFDzkdz0C4Jrb76xdiEqC+yS0XE6+z6KfbMqRujxPUSYB2D
e1N80999ImdCyrCX2mfW3u0191LxId/hXEZhEUZs6tAqhjpWOcS99ohvmyUeKWt4
Ge7Iv41gg6Qn16DucVMGjLx0i/4FLCeCZTP2jKeZgyc/0nIreSxOzL27DCCs4eBe
Ve/mXuFackpySAdlFBvHYOIH8qUPt0owSDuHS55u28mPo4+PRPRSCwXTnCVeQCGB
YfDCRMgPeV2NqY5FHc6DQZ3A3pVq5vrMnqJ/U/1CsUjtpVnKJwYTvBFqel+4lbsL
X5+bu6FMl5jQUrVXzp7VPU+UU6EHvQfkN9pMmTIWTcbMoc5XH+Ag8JCT0I3zMQgt
mWJLAnDbrMU8D/b/sZuE1i1wId+RlfUMQWnkzoA4j5InFhHoTnqLyn3GZAtPTGbq
WF+LXHqLWGgQV+V3ocYK+aMfvl8dvnRDKSezz160XNVrUYvHWe0Y6LB2JQT9G4q2
2niyKEW2bYCGz+Shxyrf8Dm3OzngdYp1eQXg5YoXBbgnD1VWRIOjiqeAMuQOzmzA
jT4QEiFRJbq1M+8ymRdQ6J90/ZQrth92dfgjMUJ/0/suod9Z1wRkAQCLlCpNmXz3
mXT65gb+nhj6Af0h5r2Jm13d+Dod4c+bc12NK8ECOKPWcwZOrgmzLnRBJZRHXief
Pt7hcvqkSoo+fX/U9nvcAKp/0OHvBD3i5Sfv/8E8LIetwirpz2CeyDLFkAww/FxN
MX5m4jM/0YLcrvuv8dO1iB0CUIMmbyn201Zf4jgGps8rhPgyeMDI4h1DwC/7Pgh4
w/6Cqh5vvuDnTYrmtckq5zT6Oz3LJloM8JYhoN2iTc+ahiXdG5eD8bot5KAquFBq
vL+0T0PkRlN3bcApXpqVYno5nGeADwwQ6ktN+URv+1M4Fki7LrGBUFAMiX/ZRCdr
6OuBayUVPlHTre1WBE3bMGNjkuHlpd2WL/4k/1GB+ODxILLjjZlClfbrbYOGVbNe
JiRYkF5Hk6FLPRE6O2WG/j9GEynea1rdGyc7kC3U9lL9xn3dAEC0VX56QjmTNexo
YTcqt/uhUZrDOSmc68cBK8uM3fmPrNXStd6bn2fW3cNJ+d9letRQuoDHOwpfQjnz
wNWY/1QhNg9ffjmLRPmh/08ivZmKZIfSC6hN0SM76GBQR1DTVqpvgtvkjVL7KLUE
Er1BtMravDgtlmVjri8PUPeq4UP5elgSSEtP3gDp/EeGWA73CjJ2n1bL4+gNGIhi
aovbZX74a+W9NGcbs0YTJWi25gVC0SsH5j85nKk8Qye4/JCYo+O3LUUj1LaBVm4I
sBt/9R03hixfZA5Z1Io90Q7FlA28LLeyjm6ckdgZ2IjQv/h39G2WPQfCd5NKczOp
LVRBlx0jHvw5/fcKAdXOBu5h0i9gNDykIGzJhUpNB75QHd7vdWcPUogLlD0Z5Pqv
fhHd6PHtbwg/IKN5DcC9cSHDz85VE2iGTqQ6lV3TMjXbyhNrJi7k5bU0EY00r7Lc
oxu/Z6RW2XQe4uVj5b+EX1eO7fK2OK4OZJ0MhvnKD3LUXFb7jI5Cd02jl4S/+yMr
uTRYR1o7tArSurtkqpCZyl0FZutluSjtt29p1N91bx9kFZ6fyJ0rFCTAXvw9twRl
Mcm6vfbg4DmtfA52GRLvO5gCklJbITQzJLfEMZ1rF6DEzf8Ig6QqjSLZL93M0FUD
tfIKFgnS15g+jikXS+JzKonsIKmiY9iTdBAlGJoBQmQCpLRuKDF9InSxl9a0LubP
GLDf4siNLwf1NG8CtLsEFuh447b6sKDGkIgTXmqy+d41xJc+aUIkitxn1F/lJmjr
jxGA/ubGNMqDX7zdqs2D++naF7yCNxgnoUwvf7W8N9EwBrTghtYe2R6ZPMhe6OKf
rRaxJO1NJrqhhQdzy9Bk8UPSoEDYKfbmNwPZUHH1diDOzv1elyDzT/LSdg6YH8Di
P67VSmpyqOmjWDRjJ1kgYF16PSkur/0dvK04hIV41g8Ps2muC5tC90wsHoVPxHXZ
h871XCVWoplBPCReeB69n5pJN5o26ol1ddgvkc/D/9Mk4BXR2CQ708zDHCGMrDzF
l121eVem3W2c6bgRBMscbfSpL/5YdEu2D+E5Kfs0PzBVJVAuWCpqtxriXCptAIxj
lhFI+5ObTSatFpAfcNwOyDGs/dL3NfhvcggdQZ8S+NSd20XG8Zhwng3/dAyZXKEk
rorVk/A/BJ+mHJovaWeFpu9oFuIrDrqqdv6MLyCl11zXN/MCEYDkedEIy2cPl64D
sqfIeINFIOUwG4LVK3D8SXPfoXpdm9lysnmr3FwQfd0qqObaS8eC7HgRSgO1wAPg
y3b5+fzFmzq2t/PVeQ4cMhQMngr9MbAnwgC1kUXoXPYP0XFFn8t6Clt5kYt/27Ru
0ITmgmpcQwZF0PHTvrDJIZQEu5I9CmGSoooyw/eSkT4wdsFpVEK45hbn0Fll2I4m
wHoLAAEa0kHeVrOSMRgntL+S/c+0Gw7oDVUymwRRHq15aAj/Cpfk1H8+HnW8aTxZ
cLKDk+VCX+EaOxsa38w1PYQCQCLlnkzYpJQuzHiqVobsAGTMnksBR65DbE4ybhlc
18/jxzycrQTkzAhjzDmFnYnZF+43UFWTJdh7LqWdzGCA4PpllsqdDg21efe2KC+o
z6NcrQeGCUrJtwWX0VbVmZb9tydA+0nDxE9OpBLgoUY+Q4m71xj/5Ezxh1qj2yn/
5hzjsgSY8wPOkzyfofPDM6gScYT+DbF92sj9xjtTuJh+ID6zjTaZtN+3gmS2HRfn
JPE1BzY3bPlOZwJ5aujPsgW8tVFL3IL2LKwKKVMO9ZI3TD7j9XheQ3rjViKuIhW4
TncdUB0j7p+bDRUIMIR1d7IUP/YOMms0eKf1elx+YG/VFUyxAwNX0VITQ+HJn7ce
id7+R4DsUAy70+VYZcJGUWM10ENB5Hy1ciM9DEY0QKgx3cxTArtcXHBEM6IIiQOA
dJ2MXe8XI6oIIGqCjNJilS/MDiT14BfF2AJ9f56SiJK1VYJGumRta6zw32XHw6Fe
kgrtJDIbloLYKwqhkZLVZplgQOZuKAOtI5GvBoKsSh7FdRSz1LqPb/3xQQMkNIT/
QaZavxPBEJHzythiQSasMJXgJ2U9Bzj5GGkK0rB9EV6tobo6CATuGkcsGftHfBwu
nBiAHX3gMY+jnYlKsT4cFpiHbPwJ1HIQxjxZMc/r0534eERFjIZjyE2NhS20+dHy
TfdEoCNKuVzi56f0VcmI2nl2ukHymqMjyKQcID3sUBcCrOPqrZLqhdVYvS9FWWrO
ZVw/kNSGz4FJ0jZtuSoo1C7LhMhtRX7RHu3KRE4ZCj3yoReg4HiEodjKDGg2uwLx
lrlvWK4m/t7hxnj2PcJtgSxRRXbnE7yo/SaCukKIemMkbWV+RT5TZG1xhsXYVnS5
1C50JlmibqB0HlEVIE1V9kc080PFpRu2V+YihmHRQ0WSMRkSske9taJ/5Ui+ym31
1m3L+VuxYoFssKJaFM44y7s9vd4aFgPp/aNHAKNn+JCfkcfeCMs/Hg81z/s2WSxc
4rn1FDhTA9IynH+W+n7rJAiDNHsTdNqOzOv0T5BgJY/2NMVFm79tVyS7VOPWdQTL
5a48AjfSlK1EiGkI0WaAvXQTyrLDBO+3Dj81iT8vJIaRAL69Jm4iv9SZiOCuepVV
M5F3mRXjGKJjN8R4s4dhzm9uMvSl/NHEhKgd9Zgpx9WPLllcApCdNUHIdj/EWLIO
izCch0ZWgW0VdLEHLpddNvr3cb1iWx+gi+bYLRWfzDYLx3U5xUR/5hRsh9N3qa1Y
mD3Pfo1g+SBgPxvngH/s4YKWU+rEi3nGNGxObssgMMiTKxN227CPbBVYEz/EGMQB
5zXBfE3UP2dncmeKKbtNtlBLKwmsoSI9SMu7nevfA1kkwLHidM/b4r81nyDP4uPC
CBevCTwfhhw/AfCaNy8HzMyZRSmH+pDjuJTn+8UXxBD/cwukXcAs/Yy9cs8BSDBF
K4kKZ41Lp2KeEQ1ZRSrSLsJPo9q0RVseca+Ix8zsBbq1mIDpu229rcHhuYD3Hg8T
yQQpMMIYYG6ywd3I1welvh+dNcUf9YhMMupPZDGnwu398vUxv3uTmlQQxQgmRrxK
EMFgkCQTqCZQh/zRbXweQf2HjgpebXCkd8izmZ1AQhjWpj38MLAlmazoPjknBYV3
IN3X05+vg5dC1i7PZspBoGDF1CC4SQm2qekYwJkKab6wxIgAzd165D6/Ua2eqdk7
Zb2pPN+jelSVlDvgIjo4hyFrEHDBED5lSyk5/sDFfLM46VqIRJR4/RdQ88Kp3EK+
8Yjt+CZD5aYsS9k7IDNNb0c40WTw5f6QqQK8PPH4EzFjcIBH+9fspRyZe9SG7meU
DWq4MsTppXr9eYDoCF9F+G8BLPmQ29KK6mx/oBW45eCNJ8DUqrSLUydZUSCJGJA1
ecoO+uN4N9O57TY20Mfn/eP/eqs00amBRXG/D2GpuISqUamIN2bcd5Uy09g7vkg1
RlglDF0LOouR/glq8JS9QbpZQU9ExanuiIWOo/TI90AbzlIWZkdJoypFOOzvVH+b
Gt9b/nsTxzs+/BWe2nUD7OaOaPO0hbyi7iLFuvT6qVRY2P3Aea0ol/MM9Zfi2tDM
4uMC6QRWid6L/y8AoQB60DroV6T9+MW9oIibRldckcReP5RKe4m+a7gsZ6CVhZ84
vzksPttag/WBV/TnykguO5BURnk9DGSd+gNLUJzGOfBuO4ERf/SEZemuUQbNfVCa
ln4GcKMKJeys9/FwEjOwtVng7T1q+AnS87wxdJk3JDUcILpmCrqpUbI0b6bPBK5X
3bcw+6mAbEJi2mdL4vnKKGdob41uG9uxBglsaidVHtitsJmMtSAPDe0gUxSrRxqu
01LaDlfr9LiJ79tvK3N4ensSPR6IvsFxDama09/xDQIBoKkvQ6hF5GKVlyJj1sUs
v/wLpSV+kITxH/jQsU3oqSTwM6Qp09g5nDQsUuOmGKCLVG9fmiaoG76OIjzBJZfx
tl1o+zrqZ8RPVl9i1JaajNWRHMyjDsMci2iTzMNI3q72H0wAsD/d6A4kv31A53O3
dMsU+GU3o/iB9DufuUz2Ev3X48gQMzt6eAGmF3SzhDgpQFrG3BXOaF6KBtsPmrDR
EBfohO+7UtON1g3642/qs5WEsAMXZkrFRgbZ8WBwwoCA60XdfUqHbzRGPwb3krkq
cTpmXhSsRK93eWISez9Mbkce8Wr5QgyQnqTfN5CglIRSjykl4y+7F0Eot1dXSck2
zrif1JCKLnMKcYVMI2HUONLrzk+a9l3KjIfD6VnV3YEnVhRz+L4DQm39hvabSPID
9+1MqVI6LFk13dYVbv947jPfC1HMOl78H4XK1Pqmfhau4zdbTRVERriFtdKQDV4s
ME9zLoG8NMyodFT/2vQOOzs4LNZWNQvxgE+x2SFKSMbJy/cnIrLBMzXvH74/onOM
kUQW33lzcIUttYUFXefkeCwroipSA5JGx+WeTWDvbM9TVM+/woWhBrVqdxGsIpQP
YL+95M8roJ6qkhMU7tAPeoMHwDciYCzqjL6P0vjsZw2c0pnL/3sKE8++MrRwdsTJ
T9tIBiPOz+PIHPrMixiuo6rQ5Ju1QHAziUQUSPQyc6EXjXzviHeUhAs7LH65S24V
5dV6nizYQzIoazBS6KKrV1X+PbMV01h0AG1iV2FHFVttUJTiakW6iUH2saRk1SsL
I/UrRvOobRuFavKOT7vCCkBExas846GKf+yA/1fXRn6tkq46x7jwCaizFmKOGDz4
Ha6nwdXYLwEOotXPikQrC3Hnb18p7moF3m8fFLmClJp5K7PTjzQw0ylAz9GO/EF7
PSI19LxGKRnlRDR2CnQ1xRwzLImDzaZBwlfSEa1N6SJ/rJ7L7S29n+Pq0v9ntVH8
qRh0aQ71wVO0Z5Li0I2Oyhjn5k+cgOy51P29sUGGpmDoiLopfVt4RqVSjMlEMKUJ
c6aaLDmn3vWGybPFgYmDewOARORE4KvjJY8Da4RraUGJdxzzxBeDtcrxUSTS/79m
YEV0bdm5QlQKJ7ELlwGeoK98jrRMgiwOxydU9nYZPqfjBOMTb/dSwtIldUSNBRW7
DE84UyYn3JaNbXXOqVSFq5eC6hUpzXEFIktvA5F3GJzeBnV3eqkOxwZBkBeFuLxl
93xLyxBFWziyGoJhu0SfDGN7ZYRiMGe0Q1Ok3LrozDeM4OrV9nXTUv9JFz3CEZ9c
+Mn3KFFG9nN6EPXsSXdEbS8ky3jY8iVFYnZzhoFJkVpZe0I5GAwulvW5QflStJ6e
5VJhbvWL+S/NVF0ROrQdChWzsjgCsklCEoPaT7XBzbkJvtCyI17DUsVNrsNyy2TW
rItwcdx6nar/a0aoSMF86emPbva4tjVKUkTXYvCkqCIfTM3AsygMxXCIPuRe3zsv
W8zwL0T0FWoFydiVfctmWXbpVB/MAnasqsgq2peWs0yFtuEVaH8yNQPf8Y5msJMA
jKmI0G0HcUrJ/Jp1eny85f1UtxGpsSzHTiUs2/HR7JAFFAFddj9Rz8EugJAFkQJT
1jGQBqRoXlFCKb8Q+OHmbjC7TvPw6AOCdaGFmwEi6E0+Xmv5ebDQ/9+P3cd9UNQ2
vCQU4VQ1P4OTQq67HI0mL5+0zbQoxKxK2Cc5z1uLiL9ZUYYKMECfmj1DtbJOe4V/
psaXdmMQ5d3qIPDXUam5a90AtcRaWRJ5rFZykrKNme1UqcQG1NxooJk3qwlPZqa3
TPmvszh74639rXkz6ZFLnRHL/05rtBtvBWJ5FXvp7Kzfpis6hySfpBpy/dGuFVsS
UqqYMTZfFR4Z8WeNUNCEPXSInm4MwDq5TQsqTvxDIRR5EOk9J2Hhst1S4/CMGhCU
ESsVwm/03w20g8P+B+pGerZjejVj+qKu108P2fs/5e9kkMDucnZHmiEakSu3B+2z
5OBZ715sXtN6XuGabAinqz2AwfSUjuy8C6dKGlPOpl1WZ4+UNLlOz2u3mLO+V2Rc
n5CaZfpa3+/t2sq7uNO6TS33Br1Cbn+0hPu84TMklhSoG307wOD2Uo2mCpjLQoI4
OTXBh+AQONEN7s6Cp366CNAhSOOjmGQcgV1EoRHGi93q+vF9/HhnsHKpe+Hd6Dli
RVkaqGyNgizWkx9hGz22vJF+ekQ05f3zF34MF4FVOrC7NWx/UmVUTpUek2kRCX+A
X3mGteKTQSXVhG8udthrcjTXphryK3UdhP8kzpnF8rZSVuLsNRGMG6azmTl6SE9y
xlUlPW45Hd06OCaKldpqF8tmh3u4PP2ApjaAdhKE93o8DNMdVSmHZdzI3+Ek9yBh
EYAlnzxklHx5zOkitQQnxQTPTzZqckFoyAJB6PwqbK9LSyV/2pGrkcvDEo4HGnE6
B7OZrmRAVN3AD9q+PmOB0QlC1UX+mvVtW2d+qShRscgycBUjeQTmrqLRt4e+ZQQy
mvqmaGHWA9hUSLGbXIMehURxd79i9GP4VvSIcraMd6vcvmSEPTk9JZLgtc+nAa3v
hKTgqLTRbRTzGaOGbXoba8grv3pL0KBHPEkkIZJLy9Y23Mv7yhQEyMkv28u5WELD
+lwkGl2V9HpeHUV20Y/b8xNLpYPI7OPAqL2DQ2OA4dt9VMqt6BhkLdlo6nsMbE/X
du5BeeWy/Dq8l3pgo22Oqv4vhZJiRb7Czelo4tAlcud8hm1lQqvycjgSeN/crcmN
iT5uiLaA9NOabdkIDMkLQsqYXvu1ivqzl6HEJspG26bGncZ4hjzRBxtf6s7TI7Iv
cRBzmCaU3B1CHLdBfXMCJx/2/kycspAdQVTMA2Vv95yTUocdqSBzzNYb+hMHs+k5
q9VdDryabFjV0SqSUXw2QkPNOuyqupbMhE4lsniWFP7xPMj1EmmCL1o9sDKkELs/
s/1MjTZo2COp/hlB1nx5slpwva+XrSwCJLnmVDFG/tOnwiRdcl1lmRcoLafdv17i
d2np0XTPxYEnCR0Vg/Bb3zS72xWa30OcFb/fwJSsy7xeimpaHkqKBESD5DEIVlGa
fZ6/SZNDE36nehB+ihEVndf7peiPtCz4kYU+vw5GA+IMuEpdYQUg2GhPyxtptGbe
FyWJThL021HyEy98+dnLwmZMr3LJqOGF3ZDIlJPO4vX/TcdA3mDbK5AB+taGVBiP
sJAeY9DW3ERPlLFK3VJ060FWR7gc4B9X4a/zO/Xs+fH2HV3ZLQ0S7g1SQ2qx5FEY
/hffe1kaKT6OKUjk0W+7jXP2gxTPq8xuem2Ugz12X9IcXxBj+1Q+SvCHzmMZOgCP
cWI5626HQbjx1/95WpN3hNSK0sNtI0DtEia09eUxeBEzJC2u/7Nxrpv/Ugi8danD
180KnLjBQpTEeUsTizHGf1Fcg8qF7Xqgx0toy3+iwVheKD3d7Dhqd+Djgubu1cw0
Fuu+nPDflBJBhX+7kHgCIKQw8Rqtek8m6JvORoX4JA5CpycTKaHgCxA8iJibL0jj
Zn/hUqmqP9S1UxIKu+j1iO/NmxfKBp5aQjCk+YmtdJWsdYk0pqm5izUvIhR5vXau
znUUoerx8AgasYhb3gdP08bXRH745Edc9i/UWzjCUgxUvcjDj4pKdcVSHXSGbYLs
IdRO5WqALK5Hc7+Mh8ErvR9/0asas3B8GukwaKPIoBPtCKSLmgk1KhotXas89jla
l3JMCqbT6FnFJANjvagOp7OYfqGiu3nfJYdyyM+kMw/WSAY3rjVdXtDjT8O2tAtD
uOuNzI77jPlxQjRfv2YQhNYgkkV7YvcErE6X617BjCj+gjTK6VYZWl8y4fiwUZu+
1ykRtWPBIIN7ssqtERw3ZWlSsrYRR7oGxLaruAHgt1yziRRAkKpqViV+P86CkBt0
Y1uD9HZQZqFKoC7LFOoIS11jnzfbWdSIIhB4mOilXAsK2c6KZLhCjggnbiCc/YzP
cnNqFvbfy9tMiTCrT3xhiV9BDf6cChSqROCJqx84UDH82uqN5Fo/klBk9QcrYU2F
3zcetxPV4zg4NzyTobUGYn209b5p7v+12V/CgNpIVUy70C/FE94IGjB1RKBARIEs
5wuOWbTNK0Y+j22TThHdgXX6scyo0YxyoaDGwUz6tx+/yp9f2Jwhx+K7M3A0CKjQ
BEvLrXR2qSdpdeYcQR1QphxFnRCA9kJBsKNL+qODcxkvd+4wl70YWxe9yY9/RG/h
bEUvN1E3raDvoRbyqB3m+R5lyGgF1d/BlzpHMNkCgwHLDrJIkxNvrCkQ7g6kywSs
vP/COz719z8/egNYlr8fxu5wkEcWtL8mX/V3RbTtmx2gG80Vv5yMTzR2KsKgw8QQ
quDqhxqZUASFDvHsjKeaEtgydEsQQmzW/Y0ho9UyKYkA3w+YB9zQ6CG3ZH/HlC5/
SGCnXH/vaPSLMpIda4LSRdhdPNCLnvGO/3jQi03XvpPplf00KTPLNt3fsBA5gBSB
ZCPnEOo4eYzCv1aRy3AB6GI9382Vkf0Lk75oCUlxv1mZ4yguNzZ0IxaaQ320d7Nc
m7504RBIei83P6zIK83pNjLWQdRjHIxMGXtiymuinBaCl1XH8TicF58f/EgAExnJ
EQTO47Lnqpi3X7mNbMhljj7ww7sI+n7ALdzDQ0cvabwt+AGZGJf1oNIB5NCGgIF+
SUceceVWQDGIUp6ja6DI5cuTBb0+z0sRFzI/eagkEZvAK6EVVzwHJGzi09b3eucC
aL4nNbINrf5rJpvUvcz1hkiq5iUlpVbfIHwMlgKZgDCuJTYBJTy053IUiRyJMbKJ
lNY4tZZKbgIV+fsQUsevYVdxkYOg97cJEqMgumeF/ntz89Q1xLNQW3RIbfxjP1dv
QTt0cD70UZkwwMlc4T/FNOl8NjdXBaoVKhH+lBFjpZ1ER9QZA3G9BZMssB7P2K8I
ldc/pLYCuRY5+/aT7Yds6MmyqOLjEMrhlE78eX6ioA2XVwtge6xbyPC9qOD+1FiW
o1sjoiYJ0N0R/jFPwT/nTPzDRSu/kHNsYmSSIg7n36rROGlLTtchu/WOoekKaZqZ
NHgsG4J5Z/YOCh+DGUUDU7YaaK2caqYZnpkOUS81bF2d4qe5WT4oKEP6N1Ew0bza
YUPqfU3XZHbMT5r7WomqfrLpWK1WownjPaU1J4L2k1DQP9TcJluvdkgGTZ0pkspm
uxfM4h6TvmBhQybpDQb/LMzuZkzyWN0RUtRJUhxFqboD1gKr+r7fZDkaIYieS4MJ
qMQpJURLvX+YyfJAcFNOYb8zWycXLpvfr6JXBQ/8z1wiJ+XlpWP25iyKaiQCysua
k+80ktSoEIR1xBdd8DpO8x/A5kTM9l4V09uVhvqQ9/6glhu3+19kAlhO8Q5esmp2
lMjoELze9Nbm7elSdtTSC0iGr5JTY/0qa1FNHoOI/o21nR0+KWzMXEyDBiJdUPBl
JtR7QYgMEOBd0jvwWSVltJUdAyPytuFGmF0FJayNqjlEuPt2HONR7FAOQ9K3qb24
MkLq8S63LRsNtxCh+zM/7w9rqKV6Ev0Q5CqqlgvXwdq5zZFtSuYWpXoW80J28lJI
kD/8ncpVrrQMwLQMeUinsSjhLr6v/egf3oTTQo6K61aTbdepmHD7WrWyIBPIfKOF
NX/O3t3uz/ejO+Ck7ZblRit+JJZXrgx0/TvXGADM44InClwPEitIiVE9ThsvedLn
XtkfLQ4pcJNvdl7+aeKbgnYSJunARErTYNbmglzPLSP9jPk3DuKp+ash/6MDObhx
6EKjm5XlzDrotFwZPLR5oYKJ7IXSGHJUqmpIeCsJg9lDGEtGQJTVtrxK7sc1dEmV
hcIQM+gVOHldaPgcJ9fDznEx9d5oNaiC0/K9MTBYkrvdKLzqeBftjsAJ+gLcpRx1
EMdPPjTkizkBU76gwlMzy0D5U01BfG/YW86SHqbQY/ovtrc4YnA6zckypcYOyC+I
+Wykh1Tp5RF9l6DNYFTaJK8G9uvZpJebzuzVBbcHeaWaj6mzoo0SJ5chOfCCivzA
Ryqr+qTTOfT3A/Za+RFz6XdNJjxRYc0YLb13qcOMn82OXysQp77bIYs+l30mHoZp
K0S4bHPtjCLGl+KEIRS+R+ASNJHXW3Nfq09w9vZJg2f5fTTEV/Bbl2kXzfx3l40L
wadRdHYp4U5r7Mvcm7DzA4zFMsFBMJVYavBOcCmIbD1FhFaNGaZqZL6jGIIwI4+O
X9YMbc+R/sZy58mlq+0HepNKXeEdQKdnJS4znWqsg2rkx4MEhIK5pYYaytFyCHcK
x09o90/IzrwO0WVqthPB3T4WugBW7vBvqdvvIjNxOgCVQfTgaYXTSLnKJW8BM448
siHZV+W3ny+8UCckfAc/Ol5EHTMZUJPf/npJKj5UM3SmOnhR+H3XHRenlrjLVLfw
xkV0VAP9YtE39nRsSqpWI1bvE2z7IUrVjWfgfPmtSvallWzkwF8ZyGO5WFq+jZKy
/7pgPt2jqAlSybST0/sTAXv2sB8ZymPQFpJSqFUTielMQlkLQMgI8TrlxkKi62iy
sxp0IYNWyDrHeRQ6u4sgoC9dy8nRWITDTJM3fhV8C6O+sPNRyZe8BA5cVKSWI9lF
xP2Ewk2A18R3unovNZsWqdyOCC4ffjq5ohLFIFiAOJiGrU/JLjy7QV2gkhsy1gnw
0GQrJzjxHa7wT6vtGuaTVrSuNaaVbX33zRXtNn9GsmoZxR1HTyIXYCFS46qL8GMb
2IprqwxT+Mnl+pjmlzjBcCNGb0m/z1ordceQMSZ96UiBGrFVJ8xKMuNwAZzK4+TF
TreKJWls8bvKdBhLrYrCZFYcAA2ol8Ve39d1X9GwBOcW/cobH2PCg20zryAZa8WY
vpU9y0KvV4ZgcoNQR8n4g8lGl/bQIWW9cGiuy7wpE3PhhOaK3OYKFYR0RljD+PvK
RNiSn9o7mrwSrUGnpqutfS9cGARQCz/tojnBfdmvSZpkltXGu30szBlM7z7KiWWw
KNGgbHs0CfTpXKcUxBst3A6IKxfsqT8prTZQjOWhlyjJp/xVRxL92zu0Bx8yFFjo
di9ezNu6BLqhI7s8Loei7yHEZ7o2zxck4Y0Jzx3vQuaUB4ZyBVJPzygtnVKARRTY
RzJ03yDfK/4KH0+3ssfiQlMMaIBFYGoUhbW7l/SQUTW7wnaUljxGlZi/qRhejScG
bNtieW2i7MrFYKQOD6KK+THVKU1M623ZslP1Ej+P5HK0qIVZ2J3sDm7IDbwLoJIb
Um6CZ7xUQNxK/0V8hRw7WhSyMIaMWxCgKADSG2kH5/onyyh+2ZxUNSyxE5KqItMS
XZ0olIHrf5xW3ZhhW8yPsNNXrcxGQWS04hYcy1huR4Mpoaon/lanKFNN4kBboHwJ
SYWR1X/hyIHs7W6gEZUvwjssqryO01UpsXwcSf8ESiHrv29Da8KLQaEJB9R3DCGf
LPMSorGCbeIYDs3YoD4gh2QWfBN7q6ibwSkpFeh0LQP88L6yeGnKkvsfcm81adeq
ICWEQi1jCJ+nHtCZXofEdW0YVfBbU7tg5cMYGsZdmd3RCGvCGzT2DolqhhwpfJXL
kSKbeMER3j+BswirIQFin02P+IS+0qhBgscOAfLcD7M7VhNK64F6LbZ6WsPQEFVB
SDK1U/YRI6opTnKodxxqygt2/Oyv3lE4wrwez0cXQNHEBxCOAdVU/lxTAlmOx5yO
SnVjVamCwTRndCTouzoq/74wVFw6jvP9b9Q4rc82M1obL8EGoBnrlJs8zjJaqI+f
f0AmYv0gDdxP8fd36xT+aG34dugr3t32qNHxVSao6e6EYOmNizOIvwURZJ1Clq1g
r7vg/B3X7XRgkOE3D10Uu/Jm/xhd4ya6RQNHEMlCIkVXos+Lk6G+qJMixx0l+G0j
Ldhn7ZS2G0b5vFN2QWs6117BrWWPCjVVL1rgwv1va/KsLYdpD9Fb8pMVzcTceT0G
+r5MD+JbTdDp1szNawlnoM8Q0hm1bY1HXWgUElAlSQ7OLVcfp4Fcwd+cBvx2MTYT
v3i/rB3JZPQEpGt5F2DTwhha9jZfi4bHOeOnZC6UqhjZAJKMcOsoXUgGW91YTKun
Y+SX0zpRRxy4UZBv54Cu2kaML7+1pCTYjsXuvRv6ww7opLYSuhA14unKfeJSdwuh
ilgXiC1MGRnN/4VJcETKXlUaR0MmwpZ1Dv24VxDk2WQ2acovj28NjePk/t0ti5Bk
k/Km/F/HCwFJoMpJmZJsic8NCYygruWayrb8yRwcWjabfImPvlDI3EFiJg9kpzXj
p9CkAleMD9syi2p8CrHW+fDhpksBXpjbeYZ2Y3dicJBud1iF1LnMLUkJpOZmJn/z
euMafmj5LR7WyW2Y1F6Uyb21yY88a4C4sEEmFRhMqXqntTdFZud5skLVgn3ff6l5
jxhYy0klIYGyluwZJxlNqq2jRHMU100byfxb2cTmhdLQeqJYiVaJr7NbfdMwAisQ
2ffOWwcHe6Wzz1TmWvK6vmD5MirVRXWB8Dx9fXVAZH3iGsKu33JB1lP+GGLay530
8X+YTLF5+BeXFrrRbIuKnGCmxE/vS3kJPqSUpzwlFKEpK0jd5zvDf4VZpt5e5svD
uM/tn4nJac/IQL3bnY4AgyKsZnL6ZQtcOovKIktDzpm6AkpUZXeqXPqasgUXHIhg
58LDqbekFMGcau8p96Lv7uK8nfbsv/DGBiA3lg6qNq83iaTkEU9DyW2PNm4vwC3T
gMPKtBH4nwjb2etAdIxWqXS7/ovJ0eOwfsb0zTs6jdKF5gJ6CZsXA4WlZGeuAP8L
xDf1VXfUnBeEVHoFYfxaEcZW2f7XvNBszex0tO07jG3yfpGSgXj5tOvWaQnpujSJ
i0v7Z73almZ6EBwRU7R09nGVEdsrW8lTtAaOoHIIUG1Y68ggWWNndPrh/EoMhKIR
8TG+mrc1L7z3ZHIKsXpkJd3Z/Csqgabx4np8g1JGnAYq7GV4//CiGmTM5LGyobO3
yWidEwFyCewpnaDpXs7JZPpuXb/HwbS2S6SE+3dRUiVdh/lmkll3y8EFa1QVKF81
FHSBYESUTSZOYpvZA2qr4yLdx8M1EXinK8Yuu0hzRE1iEVKJODQSDRPE4BNl/lGR
qpMOPpfk64jebriWZIfEtugnfXf09AhzjEjr4sHlHrNS2+1Yj83CWnyqtAWnB778
MowT/pwjX7beSfbnC0Yhbji9HeZ/zI0JcZLfpWXpYmHsHN5sjQEUwTW9gklWFo1S
HE2j/SaZKYe+5EuwuYX5gwh3Q04LoS3+liXTaVE1dwVOqqDeZgycnBK2BwfpgBF9
/Bueb0Yndqc+jm3IeKwktZ4NGUESFTfzd5nMJwH7QeCDm8Z2/rmDrs/hBow2lvRB
z1WuMuIEIVVP4uA8Ue2/iB3ySMGkgMsUZydsdvZoLgooeO5rWV9kwNUYEgf7DkIZ
bCPsFRmOmfvRG3lMfGjafoZKMcPCy4iqa0FJpM3WawNWRKaVi1qtANGGHQKgHzAE
ogqkjftRNswMDzZk8J6/R7UBjEhxuem70Cd0czKCu0yaso8C2QmHr8rtOK81aclJ
hg7Pf9reqvUJKVclxjk27e378qg70Z+cOOoTTIwVK2lHo2NjKiAhGwmN/j14vMP1
6EoGkuG1C/JtWcs9AGrHKidI/JneZ7OogxRNCZmAArVWGbxxiLy790mogO1qnAi7
dWrMpiSzuP3rBTYGNBDbZyiZHMSbwIOEwFztuD2Bgc1cTCMjKKaS8oDv6EsjzN0a
aZpSheWuEtfwndH1mL/uo9RTzYg8+m/1Ag9XjcHEBmpvR/NWH+Yh/xulgBT5VurY
MTUiTzK38Z5767n0krFw8D+cTR9ZSzTfDojbiF90v6tAiVJ+fftLV2wnUQNB1/0B
Ap5H+7H16d8ukCuKM2ZaTPIP8vcore5LrTuDSlv6L7+EWnkbRe54Oa2sJ8NQY+ik
ZIFDUQjx1DFn1wxFfTRXNbUuW0X5QdkMKXTUwDmHUh30mbBtp2MJWqUlljVNK5uU
ANmhHIHk7k6xOsKygMgInt5PD0X8H7cuHJS4HlUku/M2/1DyWvtcZb8zElA5RQAr
N6zNRuXAxSiaAxabeLwqV1k95fzkXjR3P0mayxJXBOKhbEPOk7NpZ9nqHSck+S1M
hgfZ8r0+8/NmKn0Y5sWIfFYdNh/4+u2HvLhxzA4/Zo6JkjI6ptKJH0WRG2UUhkKP
dK5g8ph9ALWtZ1+xtpNX2i1x2I4nlqdQdwCai++sTlLqko01LKPojGUwRZSZ3tCt
+JwrBBQNOAIpWeh6xzgPECT1st/SPU9HU8Zdj9gZIYqnT/2FJJffX3wEj+A0NXCm
958wQdljOomBkFUNt7WgEiaqMP2chSGk3cy27bRgIV2xgO9FNJWAowW35UnMYiFn
ShtAaDSv3D2hO05T/uMBMRLwbRKHXyC4iJQSmtGRhbb+ZcX8kHNWdegGMEsf8cvt
pLNGRHP3ReRAgieUJIbMg3S78YMfTto97LmI7vfdDpSf+Sn3ESoc9H/3deHoXQ9y
18s/b8/Lc0IFCw4oI0v1H5VFFIt8axyE1BXr+107FjjhZ9p+nqH/ILXpPwDAszgk
dCCVj5Z9Mb62hOz97fpTOK5ntH5jvCqZA8GAesM6/Jh5qEunZsLkWPw2PckDIrtM
iFuoKFXHhxz4u81+RVKAKM5TX8U642T9wF/Ap7MrfPcO57m5ff2NQyJQ96aIo4nr
8Co7yWTQDZnd/2n8REMcIM8xdCSugcmM5urQ4YTSf8Dl4Y2WXDdudFKUjIDwnHSw
VqGRfWIsj3XHx01C22xUtHzejnZ3BNNcF7Wi4mb3wCbVi8+Bxu0vZLGo8YZ88ioA
NCZ6KY+IdkOenUWD+wAUVU94GEzwDwFxsHM9KPtBDVnIWPIXu659RGYaeXt2ckCQ
M9lpNQqrXyPYcfOY/8V/3MWqy1Dtet3FMkQbwQ+PWo7KUHI+ZDnxR+h2M+Sx0T0z
/ukTGgbefU2yD3b+kmoKCSvQ+3m9NyKNYZt8qcPsyVbJipcS5g+cW8Nq+wVJw3bW
3l4vugvfXf/O//1aSr9YD54iD5HPmX2+CdReqB27IgWdjdrQO9rZONx16HPSW7Bv
VzOsoiF8e6YnpaWeCZQCGvgpgbfYePsFxfUWNHd6CSANB1uvm7KOQsOpzhBS1CcE
pCSrdi4GGFvhCppdDOyF5ZTeDyjuiuYTe1q+M6SXBd+38SR7yB7SxOku7oMJFoJO
rVkS5IYCgFs0iA3otSzdw0dxbQps6MrerER68ujjXbYTLJjkYh7h7hukWqt4k/7g
NetrrhQRuVSavjxjd0qTih1xBPB79snm5OxUs21NPkFVTrMu1b1I+E93mtEjulAq
LHKxlMgZnho55bw14/St9h0je0E+5RT0+XV+QxQVGJvVNcn7ta+G1JgqexjmoU1N
Ue9pvcoBijMcl2fLMy8eyk+sOFaQcQXyKzxKD7Ut8fu4tsS592CA2iJ7PkzA1hWs
iXWFn/Jo9SBK04HWPIfTc3DQYjOFNIocw6hGrM9IR6G+i7ef6tV7pcuemO/AP+wl
o4FXULZOGiO5TmmoJqWcsd+apoG9kdY4DIEuJpEL7GlStkX6X5lboYflDWGsFfu0
k+tfL/v9YsBFufhBapy3txaPvx9uChPQfQYHz7bFJ5iHaXSUpPh3R6GOAVkGY45f
sCJeRh7E/Ng4focDElhB3EYishvPZCgME3M6eejCWW7LAp/5tR3bwxZafAbISqJR
25p3ia6+X5jfLSAIKIwp7rv2qwrI1tKervyJ2wAiiUiasNOhFzNZA75lClKfRtNW
FkERLl9jVej6jfoW1hAPWjvRX40MQnXmVXrLMSwRcGxpMTqrdUtb8Oq6/LMJir52
hmLfE1GEbBMjEi64lnzj3Sfa10u4npTXPWji9MeFtdoTmLLk2VDOKIbfUrrzD+WN
s3JQojQY8DhVFQsua3+rXTaOjONd4zPcYvhmv0RzZWMRzigwfONiP7WT7S7ex90J
0IB+7cF13zFdQYBNEC3ex97SJR+6x74U+uyQiM4L/REhjYulJBnUNOVShZhn39yG
e+L9dqdPyOwJ0mWBNVwhXvWnZtvamz1PP4xRpFmyUcmL+X+PpASRULinF6/nSDgA
DW9pxc+KVOsx4jfekJh/n40h0rFuwvSVROKkqfhYuFtnExwutwbBx4BXzVNu3CqQ
s3C4GAaR1uQfVDdaDrLnncPrsYzrBNem5uhYkYtPbZFi1s/wIno5H+yKzVPipK1J
dtz8/D1pSDvnwvTab0Ee2tAOw60Q2pALNiA+HW3TSCZMvMVYnkeSpuSlkCY+D4pA
qp0LqG3gnaeSXN2+BmnGCFf79klrQOPwpfmzI79OnUwyH73i1rW0eaa3yYmdvl1d
zdJDzlLL2vU8oA3fPcKBWCA81e9Y806lzh4QO5i0/vVQqWJsAUF27aaMTrdFKx98
dSLc87QL7PbOFmEQDf4tLGY3RTJ1pj7+jmUxgtdSUoIqcRQuRkEwY9c3Jzn2KdDF
3GpC4pXhPJv5S5HQl2QR8ts2h3a2Q0N/pAUyJtHnI9LTm/1ezXOEer2LCJB49Ocv
P2VRBk2a9et2UT9mZJ8+60dADlTbGmOhAs17KKPySQYcUoOt44kRMUmTPd3l9x/L
Xwh6oEnD/ywJOvB/4rMNvxJCz0Crf9VHH/xsUTBZapBh58pI49ls+QCyVBmAzhpO
jaIckA39JuZVWuKDIx7GW74vgz9uH6RSO8SEy1GWvfRFb2E7owbG+Fn4bXwe//nd
N774raOsD4GQ4q0h+c2WeiSEVI2una9+KIeyv6YCzBrAkikz3p30v4Ol+t/uTcJa
l5nPyHqFofvZtCmQv5c1fkIKkF7b6iIfA5XIRNOse8QVPS2finv9DTihPDI8g/y/
qK9NZKDmtRhROX2v7lnTkcakymhJNv257YJup7uDJgYXgBfyvqOchm+sG3sqZROY
B+5C5f4ABSX0MVe7CPqAllje6CkTNBx3D5ZL0kalWgggcK/kjL8mEDr+E1hF4FHJ
VMbfSM3v6xJsgxsM8P8TwVrPOeyRxyolv+UR4zLCC3KtBxSKo9NzBuC2DE3fugl1
7HtOICdIsTwljeO9eIzsoKYaDWkH5P97HKSn1gbqtQJsVZNCO3RXPfj7eJBicv1d
tgkV5cnNuvz/RGdjEaFg+w3rdq1RxbzaFg7SOIKWB1zg5s9otq+r57xQsGYBlsc/
tfAgWEbP1Y43kyGwkQht1ertAFVR2hqpZHvEKZw9xNHQKTAmSvAP+pQENv4Tc2Xv
uIBj29Hbbw3uJoS4COEtAFQk65CigtkMa6tQWHRw1QZ69hJfPx/qh/ZbbTtxBBFN
14WUJn4ltSF2sah+0BNPOLF//ueAisJuZL4XcrfyPJfcL3Mfa9c+tyTdN0fGQmhU
Bnsfn4VW8fk1aZD2CbZUAIOu7qi1Jr+r16t8NJ2jVf1zhmlKdRaSXgz3WwthRXaK
7HZbZTH/sori8+RJVFw5NO6zjcnR+w3r49gFQJg+oxjB0IVGqqeIXk/iguKoB7lk
VFmWwMnVH5iKv2WEM9iT0Z4LYzRyx7JHnM+BNz5N0zwt070OmzGK/9/ExrWeB/18
4zBk7KGvPK0Zsupje0SXF39k7N3GaGI1IKI9OKQlMfKOtsutQawNOqdoIiQpdJ8E
3AD+RdSV/9M5oOGlYBnQRoJzRvVlbHp6he/6QIwoYMDuTu3CR6xK2ThERhUE9/I7
XgiRMtSnWJ6r5HqB5hGvlWetEIXVbwzJ4AjV05+CFIabWZTs1y5ZeHwiciEX36/M
mBq08e4gj6OCf0vdcNQZfgQmYhtCBexwSJFOsrGyPq+9Jiy/6v/X/wb8cRnA3BN/
I04p4LSuX7QMYR9c4FvHwlJqkHSRcFa615yru6QUweBhCiAnA0OB2KzFqBCRc4Je
HgKbCsCZgxPfWex2X6owKHIyxp51rukzpFTXlcvMa1qCYa89ryZdk43CgmZEbCIE
Er61qywIsbgx4YDCIu2D6tgGNmF16bYr9g4UXpeJqk6ruagBE3cucpguuq3PktOp
WyqOojqWtN69zNOi5fckP9bQWeXpHtsrCUyENfD+3LioM9B5X10kKNvFxnE1vWbW
DOpO8o0XMm8w7CKFhBxqQbxp8Nxhr+PK4ksbek9EvjN6RBH8WJqVIHMa65GWVmDG
93hPDhbRhUtLAsynLJdbHkRSQu567A9SoelYtES60xyogJKxU4g8TIyxmlQyV287
NAUuLlYmXrsbgKb/MviN3RbN7lJlFcxAE+CBzkBV3XQhR0SN9eOe4ObjJdpdjVfu
ioQXLcDiXZTselk28k6zIt1E86Q7T3jiTahSMH223S6loiOwzUxZZH+wZBiYaBQV
/lym1eXm/hcY3dkqjqshN4BiQTn2jyKfm3wYH7s0XygQ5W2lezqFrMvhaE5s1ZgU
5R2LZV01acBgbL5iTJi+4FXPCr6vCaMYFY2NkqcdmEkaxu4hBJmjEVFGxjZO4Wp4
ZFB6VK1WxsMUZnbtpA7zyB26obmOlSWSha34BQadS7iDj7rXohRybWWzVQ9KpENN
9ijuMF5g2/AjvZ6Cgydxo0ZAqUn0ivVPVR6lMnb9Xom3c50L/gILgcopUTQOSKa1
CbniD1XYfmkWPFPvjbMoJqAOKWkhGxIw5TmJNhmuPx3rrRasF3fPLskAD2xYyHTL
wgHio68XRe6ST3zm8guPyD4Z5+oiEleAViMi1azLiuGfbOd0yI+vmOTm1I72DONR
3K8/wEvzVvbt2ryPNc+ktFaDW4thlE1QNOXNZtxC9zvX64kYhGHMtpAsppdRdrmZ
xAJvnwGVT06hHpKTs2ha64VWOhHpzeMrJBJLLHAQMJMiwXvMk7Js//mRdCM/3wRJ
V5EsPin/Y+CI4Pj0szpYphOIQDdvK3LsCU5nYzrbIU41qBXjXrOxZtZV3Md07H/2
LwkXN3oBzGw8EtXRTadCAvy1cshag1rzZttI9zqtbm2E5b7L1LAAN0SAjKXzckIT
HkIDefDOuW427URRPylHDez6vUC1EDbEboUEKnlWwT/zI6QX1IFfpNquSMJRmQE5
pTVa7I+BM6i792MmeCHotwQMCcMpGod1noq7Gqye7vO3jTzp4cWcjzacnvesJC+V
8PLR/i+8ZTN1/rt8xwxnj1FCUhvPUm7fTSRr/FqJUC05Tr/HOxiwSoSh1FwvFNMw
wwAD2XBxSHgptX9zS/mzm5j8Dd3i94c5Kd1pe0WkcPkIXDnWWunFXfKS/z+vQp7s
U9pyi5o58dRgPgoTLRMHDf28u/irA9HjONVqxs31oNWyTNAcLKxqNeeP776CWY8k
YoY4UhOAWIMEDBOjgUACdIRdgniE4oQSc63jIDwkTrrrbXqiVmnCyEPxmZIsWciZ
YrehIEsFkFLpLSLkekcIHQaDQzpv2o3IvQMVQ3DcUG8r73s4uO2//othFMEmcGFu
ZrbGj635pChzrktt5a/txvUMCJXuOGCYdUnGTw2ugrwfPnyadmITc2CFR7i+jeWl
evo5xb9kzylwMEePJB2wTBt/Es5WIpBOChwkQ6k+zZDRAbhrbnpHUdp6gulrak9v
xpfXnQRo6NpjTR2eg5DL98vMwd6QxPw/gPHInbATerX5fjkFDw+WXb4Alte0++UO
dvpCeXwTpVA0kcuX+fqrgEqkOJ+S+BDmgGTsbLjDDee+/5EBECK8suL/+dAZMtNJ
jCCunitQoYtu5tRAIsYrMHUh4znfeZlHIutGUr6r24m3oMUj7499PR4W16G89V6W
CrBII9xodtM05Vpnaen2YzyFDpuYZ/xxXgnVfzu7E06wNYGH6pU2y+uj03gH7UHj
ke9Fsst9GsUSz8GFjnPIck3Bh8A/dnyCU+279YqpEHQvJkfsRsNYx94YjCFb9ep+
ZIK4Hr9DcRPOxbbWe9w7jMzIpPyzR0CXq26mvq5glq5owNowLTJK4CraF8Ndk2Uh
sWaK3Wl6uo5NRJqaoYNYpz708WmhKIH6mU/MbASjT7YRCAB4UZNhybWrijJs5Otj
855S3iDEPl9f0GXGHNx0ss6g2LIMv4Nd8Xyqe7zp5CFXF1v4ktu/IghwbjkcbBGh
/b9ThKK5vmX2GG3JasSpz8r4CeVv2Hel2XfyJgxeEZatnFY61HirwKvtlzgDHPmi
s7xSQcDsZbkWPwEL0Ejm36y7SgGxe5YLCScy2o+AUaEdQ2SOvR9vETw8pdVAGHbM
skR8g4M3wOZO0cF+yZmJAzB1NEGIN3/TdFWgJYpsyR2C0UGtUjAQKDu+Y3ISS1Rq
Qg/Rkk9Q2NCQTDHoClawFtIPz6nBcs5bIgEZ5+4wP0WPpVmfnznnvjLMaNhicK0V
FZapOA9x0kslsiveSfGV1O8UsSwKv+vfpFhoCIjdPx1u0QLxJflscYzSNc6cdCc9
6itXXwargRBdURvksQmnatvAR/yY/jXwsBZfZfa2aozCiRAmnHeTsMvUTPcJrx76
k01TeZa3U3oVHOgjnWIruv6LBSBuu943XayDPvAHaN4+IlRjvlFBx3G4BF52CW8j
v5KbnTZarn18OCFff2KyUuar+62xdfWrusYOwuF0LUyaFVCHkh8ihHmi9sowfqef
dkW71c/S6NbJq7s3JoqbDJnlmIBcGWWGlzWNwOFPLscQWIa+x25ucbjo11DcxahN
f6O74yGaBYO/VYeckoc9BvM28TbuU/GsVzGg60PLbYSChShos77r9O03T0T48RFS
EVN2uvUduLAmlOd6jQTPP7hsrn5cBFl/I/SC79BQD/4ZNSWnU67vJEiTwa7Lo3Gg
mwlZQv59etmE1kIn5BzIULH+49GxVAD43mzW5h8U7Dby0AcgnL7Ur8838xd3TpOg
+xXMhydkw+fdaVIkcb6XOxB/QpD93oRP8D+WNVbjGdNbpsR9yl5YOLUt7n5O1IqY
6MskzMN1AuzVe0ruyd5tOVqs/Fmgt9CO5qiiPTxvurDqQ93/SqJeBKx2UOCjQQK6
KSGKr6+IwIU96CX1tWXbaY1gvoBqNwPw/Z/kRxO6zaSyGrKQnhUpakR8gT8T5e9T
7SzTH67Hi6hfNkHB61nAHABDO15LJDyuT3tfk1sKVObGD637AAUNZRSgR0icHu+N
AWjfVE+q12Qni/N5FwA4FiFC/19ZnUOi++RjivIBsa/bVlj0rAIJzdTqy7BV6ICQ
W86mxtAU/c7p7Xpnklwtm2SZxWk6r3w3PLseHhljVKWab/mO3beaWmE5xU1NZ5xB
7rBPwjz/cZxQxXvs/5hM9VR0fB64cn9rMhWdo9XqCSmKCLF/bAJmiF1PScRDF3dZ
cxJ15D75hBz2ggZo2+WV8Zn5unVj/WzvBEOctiDK2cOo2fgX9tIrB7E/mYjrvqBI
qT8JsIZ7WAdwlKyXOUFeO/tVmhJr8c37Yp4sIBSt0Xh5Yo/yQfNdn7DFFAieQuYf
3D5fTzkLHOEM8/oeZWy9YdV6xvQ7n/hBXcCf5RM5+l0Ah4tjLatOpqREqDFw5sG0
fShwVVu/mfDixkcACxty6SGzYpgqLgD24QYeox9L4UF9hM9ddJ6VMF7SKTGfjxWV
qJOegkIZVgPrG1GdvXY8OrpowfJICZwbd11iO9fGRkg2hXkI4KKl4U3lg2UM+usb
RA5UfEnfLQHgzJd/zT7f8L9FnWmmu2HvOS78pfW2WsAsXl05Z14Ur5xb8Uhv5THP
XjmMv+Pp1rpC/lnAvlvG7mwMx+VEaFcAvxrK+MdkaIhKGQfqokdsTlL2sX9skUDP
pzaH0eN1Gpr9Ny4CDDOirKq/DjvEbyxcJ1gvKEpuL/XJxEEtAX1pv+YdJMyGwXLm
p8PgjTvbw8m4SAi8vlRNQ1DJsPJh68WjjL6Xx7oGFLfLSxENas0mbz9oiMHUK1qx
A8Fy+rGLQV0arkk46NxuWkS8CdPDwyWtsm88BTUWZ2b9mDnTh90wun1geh99IKeR
z7xI7PQowkZzG5VkK4kZTOJuQfTg7M4fbrxB56CZ/+mWfSmW2Xlo3kmdXoLEcoXH
q6nO1h8eD4WAyJn3MjTsypP1v8x9bW6pdfoCUBrfj6No5P0qA5aSKhF7aUex3FBg
RMlwpGDpT2O+A8XDmr4mHRN2XfnrAY3R7h8S63JeIr21Fxk/ZrjzT6SyWKNgBFfW
WLlOuJY3cVQA8w3jcrUas1/y7hf/BYzgSIGIKoYiv65C7h1/CCPo1nCbxwD+pVbp
8tmlWg6YP6HgAa00eGij2Q6ozoMsA1Bm12bfQyIsMVH1ZVZI6NQFSqlfXOMyH9/1
9yiriYkqXWG/roKyyHbja/NmoNTNZf5BEoN2X82cUzJrFKMS5Gz844buOPC11GkD
10Le67ixeZY85W2ooXWhbmm9ZTbcsUsit6VxSDThn6wb8xL/0b8CJml4jvISSVGS
uZTaZq9Lgqud1WX6ozW/C5mI8cAMPMj6N2cfxNiLn2VWXfx/OrQTUgEvu+uKBi8P
pjGMuYydUYfnXy/KGtu5tFdiZng1UQlmEZ0D7pSHrwYdRzhmS+RjaieVfioRXk/e
RfBPQMQjDu6NjR9SWEZB967morC/YbKeO5oPbSxjhHD4W+aWmSyRcpu6XgHuRi/i
u11QhkehELob1PgUkhfXs4Y4ifkmMITXe0MYxXa/8lgO+P44HQN1AHOWurl400bs
WvIK36QiT5cQn0KL4fiTS1KhR8f5fqbtEuLTK1WOPx19BiOCqfOMUF+GlKNLvlm+
2+T3iZlV1h7kmBTexrVs4eMIz0YJwjZQYRS1Inkgv4NTkDCkeASQ1yxmr+QTZ01L
zVQ+ar+P2HxE+xgA0UB2KEKqJpSGE9RzHZ1LSmY4v/FyPPhDSZZhBcfDbAGQEkl6
IgWMUS111CO6JlCAOELCI4QvtSSBATodMFQvYHApxzSEAq/QQ2x13gwDxH+xChES
q5QgB+JfKr9IN5zFTqt1nnmPCGaz87h+GFrZNwGmXLoxBRHTYaaQhZoRUwjBb+rh
yOHaNmZfvUZDdVub4e7G4VQhRwLlbuF1beajKgZTRLPHjWTgVNSqjBBiPaWICCyH
kfV24Zb4JTCdJus4F4Wzwzf9oQNA3UieNvM6iwQM9yU/MwadIGKMS7Tl2Zk85F6i
FNG417pfhf4RMDfIwWEBdgAAjw+lU2MCkZN3eMy+Tn86CTld23dNDyspjW0opiwJ
NjaodTS+nMbzw91a9lyGoIpHF5yZC1RetTIX0bZ0az43pJpvSUYWr7JwzkeZwo4f
kq95NCzyEnd6YRr7pxExVuz/vPZUiyBHP8ORGRZIZsMxzb5hFu8pvOqccvua2Cz3
ddW+exrvXNJruXuLMEMiDdG9c4a2RoeqtcbgWIHqdxxVfZwcmRwP/SHIGXZ9gqek
Aw5TXNnnuaYPYKQsDp2pyWitymWZ2tDKn5H9xtC5wK+3i5/DKLYrXlERU8dEAyBM
JXsgwjUSxjBK483GJu07nvBZOwD67UjqACU3zYw7Ov8TYtMAzEdBWsjJLr1qlgtG
cUrVFs5clZeTGLjVvMTrey9k8k6/K3eDLDMzqyfNB8FCf+/9ycOMnhQFX3PDaJXF
SI2MsBYbzbOTG7HlPvToo/cFZJYBFdlILPDUfxF/vup8ex8jvgEEFGbAv2+/NRtg
O5CsCGzUmqOif2CANUJMb1qocDtxuuX/iD+xEiOFr5qE7dwb6vaA96UdrzIteRXV
7/L8vaeBLNjxlZdt1AROU2tKGPSvCWC8a4nZEJfMvZqZlyinBj1WGBco0n4v0wc1
dMioCEaGsw/LkTL2lT8ldrKJ7vnqCnER/hPEzz9iJJ57aVtsfkxwV0XJciie0aIf
JuWAI3+6BlHdwbOZaInFJhoeXG/DvJWsAODm88Teer6JLJ+W5kudBl2vLyS5tZyW
tKjBVpdp6AJi6qnE/673lXvLN6KEzqwHtA2Z+54mfCpichLOXP/UyyeuB/kKWH2c
1ZhlSXLpGQM0q57Xe3f8QbimJWdJXTzO29x7Ut8h3x04ulq5ZbKfWkyaqwXm4L8J
5toOZPgVyurE8jDyMG7/fFO3eoh8ByvNF6U7D+Yg3LG1m/CzWuZMZrT19Kh76edq
5NSrNaqukH5Toqcx2YtozQGRhnn7LN5wn0E4FZWDINEtZZy3+sVzgDGC5lwbCMa+
ajZ5aHG6YYmqpZa5BrfXEyKDOwuDo2/UD771vLN+0g5MlxMSkUjadZz7hqg2Kkwt
53qKAwPQ1zCZORAE2icqrbpIANxLmF1c5GQnWMVXRPKXTfGR/kXSeLD2UVWRDxoL
j2PviadJT7szE46uANQoM2bOewFSR/g2w4PqLWxvEB6znUy00ztAZ/+GFDIUFASr
2tRoGjqEgE2ZoI1iIEI3gsqDwENszXS76/j43ZU6fQaSnDpegbQ1V8XWnXNx1FCm
rtiRFePH9KB2Hr07JBulx/gCLigCkFeDEyJt5uG5kPoQZ3M37tz06pT6XzpC1pP0
JmS6odO49iuGYt4lExbv3urz57lCCy9Asz+ukmqWdNDeJ42gm830OgANO4hZIDE8
szxFLFdhg0b+pQ0LbG2WKXE1zsXPfhpjY62CwHPrhVnWsCkg9xoRn/3xExedYrch
h+4twsCAHmQFPc7ryQ9zlgkBCSPfc7sAYAUgL5FcWPbkPOYL7GwsdTlQse6S2niC
xCJorqMA8lgAvEEocV4WBECqHFIY2hDiJxmH3Mq95E5vmkaPQIXjMMfuRFgngxxf
zEoI7B/YD85+OezmzNKOY2JuTw0l//4rGpdlj8UrHqC6ROQ567/6bQhE3j5v0S0W
nGTAw9/hzbm2ZEJUYkLziw6SU9t8TWvAbCSeHJuMRiLfB66GPhOQll+SXMFa7KSw
ZHA+FHSJTQ8f/e/ChNkLFJLxNe+2cyfZipe86kwTZ5K+77GRB9yczWiFAgnbNUD1
HNMjPJJGYQ7OX5pjcijetNqdyOjd46IfL7JRmh9NTDUz9GuO6trUupNlE09ncwPF
op+wPHyKZBnbpBhXRAk+K45oY6kYECD7Rh067hDxrOh5LKQXzzf68D/qnqc6qHsz
1+q5UdrTwRSDwkeWRnAvdvqSOHTBp9Eew+XIZwKN4W7nwT5XiYOfX1nRrrndrDTx
gN6PtyrK5bYNPcaZMakTDscu2y/+Juie7nBSVoHhrNv9eNBIfnuR6Hz80vDU7+9o
jG5Bgj4fe1i/FTVqdGjJ9lDQCM1YD36aDaID1rYq4YkQzuBWQ4HYhfm/e9S6OwhT
lMDUNtM+BY9KnbiQ0tKOsFYQLG8az6mNYMhVk8lDlZHoGVNv/y4HFc/cVGJ47IAP
ndpb8CaEvWIMl1uZPA5T7jn5zxe0F8q2ar0NKwSX1dyF607ZlPTCNAyf+I4skEUB
lovALY+6SHP7DaCaEROE6BhxvrmPPNvW1FWc0nTOMiqF2MMvvlfN/SXzeZFzPQSU
9I2dV1eGbb6PNlV+Zvsx4nquCVxYnhH8yRsRpG72q96Bet+rCv87xqgLixfB1dZ8
PSfLYYLKai62OzBNGYllXuABi2LZtPX/1TnTeiqVSi3TRmKoGX0LBMv3cgh4Glwf
gs/2GQ9yT01A4KFhitxkO0aEbMBS9OTd+iHkv46UiGce+dIp8dV7WuZLZeRDxOPQ
3zEYPb/QTh8NXjGErXx6Otm4eG8CpbFPQ25Xv2Q7DjBmf7N/SLR57dJc5+anefG7
4AuAO0njGTnbdvGssQrxyF7k+fuuqONn7lzVx54orqF85TAsMzFeL87RGUbhjNQK
TvI/HIH/AEKwoA4ZVDVIQ4FoIWJQG90WuFhibBrjarC3HLQ31WpXs7gp11tam8Hn
gB94IXbyNyc9hHeHe15ZgiRB82UdQFYJO0gKRSYE1urOcupUPWFzSlKYcgoAvX/6
tPcP0AqKWS4FITiafDxmvNb0FxgZb8vAa3LwBjOJOKnqR4PV9at8bpOGgyQLY5ON
4iVAyRkndslAksToWqjlY5Z5Z/ulWnwW5mmmwtKTomZ43AwtKpoiVfo0271EqijB
iCqsEDHPLUdKShW2LcBy0XzXuDiLT76gt6hWvQRIZoF7dNwW0gNajD8vFIrSPmKF
gKlk6beLhU0LBPL+IPyhdL10qDVmIKU0q77k4Y6SnKjS7qf95Y0b1AX+aE0NMyC8
ul8+wfF+XRBKGeSD/XmT3njHP0ti/d6B84QTVg1xhEKTodat5qN/BBoEsgusge9e
HcfBHSRWstt/hKkpktxT7gV29+fNjtv+Qjn7TCgYVBG9pf3m/Qq7ihVaSreQx+WL
YdIJEHSbR3NuGSyNv8LUGBjxzjpEIVpn9QGliwHbO35H8Z6qtVXw6QtYNCWNy+yR
gSFli6Acp74HsL8eggMQgU6a5LD+OxSd1XRqSZO39JFr8reD0mexhbsIKsXWB8vi
ypdJ0ZE3bNs95jKqEJQlJchQWp2o/A4cgylwlQEQMmJb+oguUU8JL9Grhu/+Hcjm
fsrzoIfM/78d4OnkPNbFdyLOpbdu+Psa8F4PpRDh9KhHeZv7fvIY4KNQxtgT+9k7
0T0AWdLU9LPeMLXqf7dznHYF7FA8BZkGcq3nsGPCBSrmGgavXSQTLrKMUYzUPxjU
WMx7iRXnAO2VlacinupqA/TH9rvt8j6lnBK7S+h2wNDgqSayB9u2JBOL/t9GOwF6
GSKxquvLvFT2FVeAyMEuo1l2icg/7KXKqkmREdhY48/KNEPcSkGi0eBHEPzIsnmR
v+N14E7BiCPebNeMl9BM/gMYf5w/oQkKZFsJ1dtnVD9taQnLobd0G2k+qHpaTAhm
UI0UlO2GptXeUfzXz/6v8PNO3E5YN2dulIWszIYnFgz3iChHmIQYeFPYz7nwfeYN
KSGe1B1GxGoDlZV+bIMmprK1lu764BgMvox74A+x9H8ut+tPXs97VfDakHIbBX2u
Vw7duA7UnaIAWcpY55Vc9fXMVJ9U9kUYds5xmWh6og4yildA9b5IZCFDwAVOiooQ
iXhn81YmdXZRYHYlH4DTwHVqD53+1oo9rXxCGcVqB4aEZvCBEIg3WcvALy6fAssT
VHlEXI4jfhrqLw/l//8qlHrZsTzC9C4y8k1X+klNPe9+RaN5oC3x//T40M0thgpR
++kzLQCWgl/QxNgY2cpNfu7jaM/MBnaQ9OefR+tvSaGMwn2VQuxqGcsMreGj6JVK
nLHI6jA35Ao4q73f19NpynByJCHu67+0tSer/D9ncmGNCLyGz5s2Db5+FV9hZwOJ
5MM1OeFJ0o02tcSxlQczOUPuO+9l67p9tZunnSS73XbsdPsCgolnuMxDWAp80Jgl
CsHNYIwv0xeRV9uvrU21+bYr3/ljFyRlXQ8giJazdHAWP/6UaoWaMq3yeFFegMk1
H4SX7C6lMCGHJPq+w9WTfo10yMgV3v1sfDOhobHK8rBExJP9srshuX0QdJUNe0uS
pAUkq5sfuTHyRPWjLzYMxUVBLf88YBfReWxANqRkuR2Z1nQEmz0tm31ShS6bgIaP
FCSb7+EHqu0dhHGnISpK99TRZmZhMDF1BrX7pB4tITRhCu9FbKuSNGajMmAzVt0y
/58LXe/Bkz24S290R7E0YAg9GVkTCwBfX/Cajqu0ilAScxKPKcE5599eJ85YQIhT
JGyY0WjABm6oW+njGK9Qw8Cf8slOhhk9xj5E/+O3+oQUMvaMqdbXEOgH+6809tq1
1F46K8JuAsYzcF1RFQgcW2bKMNGfYDld0/AlkTjTd/CfVJNhDb8KaFLYvP7e086B
LnWp6Lz/KW5bkaqNoCZIpx4TCpmaRTT+eM88MamT/DPCLON2u1jI/aHxyv+qtKxm
CXatqp3F+/9vFUHPBoWlWTpZc4T9iPnkOLOhZLcwZ0MyAWJR3fcp0UqqkdgNviFJ
VYiobqzdUBpsEbKkkctnYzJVll1dd8o4rNwHCoyQwfHElmaXOYW22wZQPMX+gVqr
XyS9aqVRydiiHHgRUTrOACs37FMcCksV3U1DjvqnqeTix3APxvnU2WSNvsvZpuSd
Qk3UJLAIBTgYhB/Cjd6/tN9ukwqsavpGQqA+vZNy7tuKG0BnvxFQLmhGoENGqrrM
IoEkzWv7Ax0cRsqoDcgmMOQ6/TXLD4sYdZGR4WILLLe2sWBTqp7AEmutCgPjCmZV
5+R5o/XeRtr+Mct4dhvG0qmGuXGE+hv6TYHcGKXXsjVLpFwWAe+SMzEbZ4n+qlm9
XQtVx/Yz6Y4mvFpT3AN1VnEBYKE4c7H/S+kCvHCvIsVQ1qBOLny0uHewg4FsHMh/
vrXAMMgoZ3yXlMAD9pXEhlPzOWbD4hMgOP4LIsubHOGF+SfasF6t/IBIE+HWjZlU
jQ7c4f7ydxE3CAVnovPIn4k0kPPJbv39FiyWn28atHZFWDXjLgw439j1y2zwcmjz
JqFxFvvRnzo8841lwqBQyQx4ryXAbtkT0cTLnRjq2vX/VIRoyDdN6FB7/f9LjdVQ
sVDZszQRkBMsASXbCux8MZS+CkYoNBgi8tnceGRohRvWzAPwF99NSeyezSZLpbVB
w+iD9/XmMmpxQzXyr+GjJLjsX9YkL13EoWLQYw7oRmcBpcZJxxUfDy+jcQTgzPaH
7JF05jvZQVMUdH8NORpUfZ9JF1b4KZUGOnLsxtKPr2syafrKIv/seIRl5aorKupT
bQMqGigq/4fscS2wR7bdqf78MQuQzj3LnNGbq9GwVylrFRAjo2mFrfeLo03BMmRa
iR7b6VNcdD5LycYEkNqpJDrLZnkEqSxl7MEdOBu1FsizOGNT020uTcAg1GqbNUpL
2DbHz/yzIBEu8XUvnF3CGVy/xJ1AHdCdm+5p3yyYvZmBO0CqLjP3KqtiGzcifIy9
8+DEGXXAwMEP9US1gBet1ISfsN28Ou28acWCA9+IPyE1JrVQZmdwk1EgWbCSRGVH
0H0Oymfvw+RlusAUhcESBmLGGNwlbbrqZqzsEIDUbZheuy/aNio/aGTmBy23JKwz
p0gOQ2x6XXQnFEnSODf3BwJwZR1BWWkes7yekaLUVts7s6kgwiMmWHbFH/wwqsA/
MpzvFmINjCwGTOItfmsI4sS/BMli3qrQLF2Ea6eCXPz1RffaDIMbwHD+U9LNmXMP
nS6SeOZbYXWnT9djvzbMYQmKwXV1zcUrzVGirSUndBqSNzn3wPkr+2UrXmSSR30R
0J/avvqyuh+A1XG2KRop/bQVyPvMcrO0Ya/t2hKhcrXBr5CrjeCfpdG6t4/bFFhv
zmd//ppk2748u5O49a+5nYlmnd4KZ27Qk7sByvky9q5dlR/ha97mdLTvOBZ2Qs7Q
wSxeBWR3HGf0wERWEokLtfXslGYCZShyFewuhWvFa8idKIU9wM4Vu7X8SQVyc/RX
7qNuf+TZ5I6mpJ1qvYkGZNPOreSjGnfJ8VEkWaGIrhlCc+MvCqr7pShha8bis4G1
1XszBPRnUd0ZCpNG4F6ylY4qYpWFW1oAIxUKKviryMXnOHzbjQcuOOAkbYn0mFLY
1C4cZ2sNzMubkT3lUcTN+qgt2IG0EbsFbjgbAW0IevWjUkv7qo+kpvUwFyeolHkZ
mUw2DFDSs/DbcQR401IK28yaQ6azuoJtv8VDUSnzgzPypjl4PF5UG5iBt++nU+5R
lvaSH80bDq0WuLJOJXqnHCRAXJw8cGi1iDcyCGbnXk1jcbtdLgWnoE2smkG/kFvb
8KPnCNaMXiJlSyIjbJBDruBihydme5i2/W1uTijw/jK6ivHFLYQtqFCVp9Wo3zsq
xOtw75jPN5/SsGxT4aQ5DE3QP9ipZ7e7QhNhF2qJClx2rOSb2uphBpnc922rFrbg
5Yk7v9L3rqHJX9EHPGHFUKVSqCRM5889DpR6O4iPbaLfuOrSgb/Of3oWvEwzEet7
yV0mt5A4yfk2I2qJnt/BlRr4ntCp8ktYGSzpOwam3LD951NMZMPgcBAx6i8OCFPD
ZQuIjQ2SjsnijT74ITOyzx0qbuMI1VSWaCx9aJuR0ZiC0UOm4KlBB0fca5byX3x0
rmEy8tfAMK5B4ydmCBft1jQ5PieOJihd+FUr8ttwhoiPRpJ335y2hQItRLcn75u8
0E4BhFZAM86w4DKoF7kP68kzyo70PYnrMO2xeyqFXLyy0kpdW/pVFHNN9lIH073c
7jky+3h93qCSW+EU0MMhOgGUMxX6RjXvJp1jaL8TKOICCog8RcdhjPhHfEIR+v7b
LkMWpiEqS4a7dVfhhBgH0F9dIYUhVC3qpv0n2UoopqnzQFBrdyyGAi+bsnAAFn8V
sBtAt2uKlx8Oem7X6USZ9L5vppt/ADupZT4pO1PfL0GLwD/OQAAt42viHhXlljdq
oly8VxznZ0tlIvLGX1/bIcrCfk5Co2H+ki+XqDyXU/X3ikmqjVGWRrc8z4gFsEWX
B4BgC4NL7LeCSmex3Ga87VyKNI9HmJKrtRUI9Ku/aTkqTqYVAUoq2Qt9MzHvKax6
khJoRm+Z0FZ8KVsLd+b0KkZSUYa2zi9QxWpdRpW5ARhddrxoIsfukJiDV/9Dbq7C
sEZP+poyxvDFlyEUSYwh4PC4pP7dDL5eFxM7QFGP+S/fCd11s7Q4uLKtF7Z5VHMP
1hfd/wDthunmpP2P7mmif8uQdLuZlJ/67Katj2ALL79W05iChQM5+XK3dbn2pdFZ
fr3JozClelIsIUm+3jo8bKNoVar6sazD2Gq5qZZl1pisPlKsjQcN4w2QCoMERzjv
suS5tsnP4kUEU9dx8gpawQ8xQqZBYGUN2OHtXI8YZb9USHjAjQp18VfU4C1ZPHcS
3y4apb2ddCEy/oceHAMHNolcEdLBh5VbaYeEtyT3+VAnOybGahX0YreGvxr0rSNz
mcVZZnm8kPWyy6RmUZ8zo33s52yWf745s/RxnmCoiQ3EJMRmC6OhjVejaU4M8M/p
dii0XjT7TpsD2ySx2qIpAqFhsvOTHfDJtweNb72VZwpbSIYhXjARnzU0QI8oUuoa
ADxKTwRsauo9UTT9SsBvC1BY92/OQ1yIqMJpN1E0n7lsuo+IDfZwIsZo9KS5MB5l
BNRomanH47lYcWLG297sKEvojzzTD7aW+4leWJBy5PyZkNqv4kZkakUmML9wvnGz
qdYMbA9F6n8bZWziUHoYERbFSI2ZsAKMfHV3YZUjlMpFIMT+YJbOz13W5Atr9Esb
zdvZychY3Nklrpg6hWSECvMnaqilZopdksvn56XTaYv+HjNXTXYB6Ym+lwrGuhH9
9X/+/hUtCUBWBqF2TUIfJ57p7AAE/v4OE6k9R/1+nqy6VOl7Kuqws3Px/zmJAgDo
6EgXQJos3gOaT/Eps4US6BdaambsGeo8kFrnkxLOWpX3vEhU6aaIFvFbmanT/7gp
NjXpDKlXiI1KINFhdp/Okwm4pU8Wg2XCQdvjykEMpJlSq8gMlnHZQcxPOKAMPpNA
kqHFtJSRRPIrRIG2kPohgEfHSRVIed8jZTupycnFGhZyXdgwQBnuGgoRowhiF28A
oMllhARqgCzO4C6nt/qLs8uU4xYL7GRnUvPGs/OLxmIP6UATRYcRjV3+wKj4A4mx
SSFVw53vwsSCQ+pcYPqpONFuqhZmD2xsyuEkNS3P7RJs/xrybJAiYSJIzke5Pyfm
ns3H1efbVO5mVlsHOX6VzTMGHpFMPGGamlnt5Ul99SKpmmyatDK1g7/AleXAdE8A
H8p36bVDrvhy0y7SaZVPdBTv0vkKRIV0IqVirgMz9VBrgryRXSsXcAo333UcBpcj
iofHN27t34oM4mo4axPgziXA779a9XCex3YN2fH5Q88ubIjYfaWK4mhV50xsDeZo
4hAsaF283jFfFXqR3EF9HXJ+jrCBNqHTAsZbkmzmeGJUSJL/0vrv9IFc/koJLDSZ
jcYC7I9OpjKACzfe7VJqNHJL8SHMPGKt0l+Br6EEId34hCMy0peJlAsp+kr1/QXF
0sK/mIX8thwj+l1cNfkosQUhTg8ktvOOZrG2JlYU4nrbG5eShPCdMPC1Fje/CJGg
P9B53pRv8RdEaCmaRwKRAlRyOnmulHGGvQcAR+I3Oj6zcD01QKYv4l6uCvG6Muys
QQAGfgXCh1v5b+cnkS5lJvFfJFoUxxOCkgE7LvPz0n3y1JZoDJ+QIsySOWD8ZYy+
4OdprEJFiRpGnqu30ahEqnYkw98lXloIHWaFTOElTwHbo6uTjoUePtTLLlGUf/Nl
yVso0eaiumZBRqAikRGeYkkd0OU8i+C0Dcf4N5PhukNA5K4syOWzsT2JpDmXdtJv
0RFTdF/dxa+3SXKSQerQTbvRXfMfiuDYhBHmjyZX/Au+K0OmKC2JyxH9fAi8b+gF
GdhfaQ6alvlnP8zWTuFZjpQTD7q4kdeSEuniGI1ntesl8sOjiKv6On0rZxx7vIKh
sUScgoiJ0tjIxPPdxGVBtBMMNZCE9bA1Ll2litAXi864mIzKrrmFIXoAU2tQc88n
wRieBNEkDA+qoPs5FmuXkcTF3EeK/OZtP0S7yW4ATJLZ+LeB9p3JHqJP6NgEnwRY
EdT+5WixLRbWc9/mF4NE2HDXrmAakDVGR92Rff9MMG+htNsKyyBb11rCoIBLXAEV
aU50Lo4rR2XWEcY8SfjBWaAU9rhCnZCdM05RU1ujP85dMBbpep28qdkvyH38ImL5
36kRofq8J3o9zo0DwSJSHQKfZb3IyGzP/DIa4faMD7XcOf+E7+78KV8prMBYT1f+
sOChwKeEzmpJuaPVQuRwwdTIrOCI+YTgTR1Lw5Rn29swC0ITHx75774tf3orCgax
vN22P9ym0kW4f+4W53Zs0uFZ1mXVeG8VrI7243cw/8N7PNlOSZj8vHAwZsyEWbU7
BQbO7PHjSuScBYV1KmnWHQVvycYmkOgnN8t/8V6VuGLMkPAfBDGqfDzf4plutcQS
oQpo+U/IJD59wWmZAng3Niz7s0zWlMYqIYf3vgJN4q/eefdxrhpOh/mdDVdVxjGS
O1mZXCnUUxQzjQyeXpPYFaaZ8yKp/F0Rf1kwxZBAR/IpTi5uZ6KxUW5j9dUSm/Av
9g8eeR/ovLcQonaozEgZnqBSKKmotmZFmukQWlazSPRnZvndmtsIQv6ImmNUYisg
Wp7zgFXDCmC340seC5kyabcv5AHxX8m0+/8uOTTo+huupzHYsviX6SjA3sjoxTms
9WDAOSO1PRl89W6CZ7Zh8umgxt6Jf5vZ/yKhWol7LKvvc/mdepP+l9okgyqeTi6z
Uq8jE2ZrR/02+MTRwLbA2OGgodtV8kvoD/bONgmEtF5SwRkGaQrM8EBP4fIuiY4Y
Ap26fXLmF6l3x6vRcTbdQwPI3D6XCTCbW4LZtnZfwhm/kzxUqJ7Ersd51RqnRZpI
BGNA4d3D7bTSGaidbFoqmJAwjmuE6pZz9c31WRNCwuBpzvfg5+n5KhMdH6IDLlHD
S1eicOZusMXWhk4mi4qvTXQgloqWU7LtkANTsvENfZc23eR+dXWGJMvqWBBIVs9w
sOazQTJRFZDB4sh6j/bidUklo0/AixKYM2vN7jlkhSoQy2d0voSVRWTuUZP9G6yn
AGuY2ZX0BnM+FcfCJknOl9m2ICvxAZhJygbCYIEF7NqugDoHKUji7E/y9diqKunI
c8k2zcYezfH8MiqOmw7XQay4yj3AAAVVKyLJEbRwmZsPjFygwuQjgW3aCWb9hg/G
qq/Ep/cCakh6sqL4cYTwzxgvCtHicpAFel6Pf9yL2ncqiMBHuzlBbK195iTwxDR9
8M748ij69VrI4B6fZgN0RCXGWxGGeeRJS5Qzkj3aYTYCdTgC8coWqxPBUcjryAtm
4LRyk7Zew3lRikpBDbambzA1HAj4ISWEYYc6jT9Zp/phFMZmWrYIakQ6GJId5EUI
Iu9S4CjU2BcQknDs1ZT7QCDKwLDReoUd0yBUee3Vly0a4DtlRg7st76yaTQYtOxt
xeLldsyxw+EebIGe2HExAgzjQRa8gZ+m9i6H892VCqPGLak+QksiFRJ+iGB5TA+/
TWw0xOn4LTMFmbegHSWP+e3jT8hIUWHCfR+ONYtqwibyP1bzxUKFGzlWUexcTK4Z
Hf86BFqjAlHroGzbCWxEVzLCBfEOugvvGGXT0uOl8MtlFZ0Zmt6OcNhOnCK3/Lsq
3icEENWn2All4o3ARDXOiWdZ1ReJIRedZV1Kk247uY/Gks2NzIumQSOYWrQmRwqZ
mDZlkp15Sb4OIazptXke74moVxkPtj+7eOQg0j5Nc7yoSu6Akb8OZqXqpXAJFWX3
2amcKrLqE7ZWD7Rv+pBOlI1X16qlS5QUZ6vv3ECg02bGu9lTMXUEID30TFJroRU5
CJGDaBxLZrZGAKierVvISn2x+GgpCOJZNo8oA1sb7d1FsNUaxgF+PyFQ2PX8bfTc
lukLzAa6lHY0KtKuuJCkphq1fmNLWnrNtp8YfbPgAMsDlD+YPYeI7zEpUxtCjqCs
kldKsedogMBTUucL7TX2LUiMKJsHVoR0Ths2TJZ+JHNLDGDPUij5mp6nasFd/E+x
sjMiV8Ufr5Q/8mieFHJZdqGMhX1ViOOCoO2gq7g8N8mQPlGfu4H4O3SViLbm5Bfq
97b1kgJcI2Yn76WdzNyisfRWWsoC9SHV/U5DgoTNl9s0hrBFjKNORyrw3U47SsRB
iNtrjq5JPjcasjq/fJ50CYHC5pUedOrdOLjWxOhvce4EDJ5wUqCQ45vMzJ/je4mj
OTZ+/kyIvnF5oxvlQh+u0/JJhI2bTtpakMa+pb95fUMRzQYgXRnkSVo2violgDhC
HW3D/GlwO3ZqEr48pyvWSXAllCldr9231sCM8c4vgAZRl4PjL54A2cHVu4a1cklX
KtDYxD7mglAhxWlGFvU5XBfNKgUaO6uSybHLB+dUDQIO8PzrzPEMu3R3fn1Lg17L
xoco/K1Lfy03RoISKIs3mzbNBt8XlYmyi53SUCA8WkdQIu5/+fYlHoKNU5gVjPZp
F2bVkb2OObjK7Q2w3l1ApDQuu6NZeTuE2c7KnIxo4umYdf4BKvKOzI8VrCWIy2e8
JJhurojWHpqNIiKpG1Et/vj0WmLVDNrsSe4s6pf3ymUPSWkv6bYx8NFKLrIRWX72
JBL+eaaiWmPKhvT/bo7sxetFZiDRp1T3y4wb49mR/9WGkr8xq6BqVH2jjaLAZoib
g3paur27S+cU4IPSWwjP4puzaBGmmVlv0dMHOlGE6qSk0EKckAroP1T9HBNxktFC
YtNlY7wsnt2JOR3rT+mNYpd6S8oatD0zFaS9O5Zwj3AbXh8SOM04ngDcS7yj/lYq
HlhS0HI9vmCysHeUSgEeXZSs1w3iJEBt1n375kYNIyBQmbbmQca78C4iilCYxcgK
QNU05cPUHHnuv2vc03oaECsUZz6TVExsjg7dQ3csbQXGqmts0LcU7BXv1fBJ2UaK
/47CJ3LxAc+NvJzfqZH+fFLBv/k2saBNp6mILDkzE78Z/j4nK6B41FraLz2C5KYK
8nypRy9BF5iFPKkUX8icKRka2Gt7uA/JjJlQiCKbXVg44kq4N7hVIwbriFTv8eIk
TX+dhDBojsKH7brXYFEYxP/6lCEftl4C59Qp/e0XK13uvAwv3QpJ8QnHwMP5JWKl
6mXBizm+PgAIurMqQhM0Lx8MMgRS4hc5SI23zyj6FbdNRebbb1XEYJ4FRp7KIyr0
Gwkvd1YX306PscL1G/8hnvTvttvdWnBWsN5wI2/Hx+aC0BK/lh3KWXtwCwNcngV7
o+6a8MG/mUjrhdhMDlgIWC9o2UA05+zelXXFgzklKitNX+hz1h+NcluosL3VwJGD
jbGicQxMbVTsyxdQPpyVRKCIIXqLMlLRKKznPc6LyoDznjUjMku27nurOB7m6On/
zkQ4eTLgGTznL2HREadBKh08rCuEpeAAkokBlD7mSdfyoQ5o0XpcgzQdOVUHZVS+
ENLpFQsTq+Ps2hGM6JsnG+8cshPl9ljEfUuEx+ZYBsjKueVvfp+1IQSwX9j06QRN
rxjCpQ+1AETlx129c874pNrtzS0alekGAWJyvtzIZJjMBl2FKvwzz8K8+W+knBEo
N9L7Uo+4hriNVNRJdB11rj89OgK0THFBz5n/1Zr6OlgrywcDoa7ZvWTbxGeC3LzI
W65BNj41XSQa62KBcLGdlX3y7bIfNjB06yGp5zZF6+1ThihvrkI0sH0FtKjBbLou
M6Oi5sTbtSkV+4Z55oCBMlOj+3mJtg3BBkvNlNb0+SWvDlQAEoRddbmlhMlOXNN+
O6olbyNOdLOILwEzjm/CYgNwEkVqd+aH8pU4fH3PmW5fO5bsp9cCoLOxw1PR3F4y
JCvjxRyDZM3NzvU/+bvMMDouCJXLy6GXIatzx+ITU0zU5BLwy8dha6hihKufTRTq
WVnPKoDLUfzXykbnxyTxPqmf25xB9ytAAdRoO4qVt51xKiaUAdiUIdvUAsQ34Ykc
cw21JK+T7yy1Ut7rbya1yayj3WkJ9jM8nCdfUiUSjhvIJ1gLcJYVSMWkMtcAeXje
uk3MLn20jV+E4dgDLj4qA/cnXlmCLcsQ/OSne4G1SrUCnNWGpsJub4Rq9q1fVHKW
A7lESEfVtXtf06yXZiKtSXgOlgtn7BVoNUssa35ZMuT4GRq+knl1i6N9hqUZ5QbW
lzKqKpkNr4txSRPEhHIpaucp0W7uKAtYH8a92nTLvrREElAKDzWRN+hpwNKc58d4
oqGl4L7D36EUB/6eMWBwagjHSSeR/x/gq1oLEPmbDDMSncS0bJXukfcLan/q0rcU
C4WaaE72toYq41LB4WQ0J/RYykvkmzLq96D9IDt3f1LS9NLORDR9D/fn7SALnaJw
JiBpm3sK4w/rYn/wG0KcyPSBG6IyeELMGXFP7AFa1ja+uciMjzoM8X+vzToYaAzs
M7mj5HXuAfyu6/PtKW95iscOdpoOSBJxvc0bdJQsetmRIGksxH8kOasHgtYDzPz7
D6S8pP6JnWP9VatmDrbeysA/35OmonMe7H/VxCSK1A7o2kgF9noDnEkUTLK6L24l
rW7whNVu0EewCJVQX6W8Zh4wqL1dxPm5ZviwQrICYgnRZ9T+4S5MQhnOTmb1xj24
dJ7xhfQxLtXSZjAxNZSP8iVxwRme3uobO6O0FoBsN+chpahuukUTpSuQq4+vpiGX
ZsSFEXbhmM4b2J0egIJ2u/nq/i46hBzVNTHMWoepECeaR/RDLcOdGNRzcFybazVb
a1Kp/n0I+enHxM9zx8r7LqNSKey4uPpj0kQ/pGI1sAFCqSPhbZcEARG06ucIYlEY
RX4WWj2SA9C9htJyWhbyUYuG5xfY6dNFoHba+1eugyu92FkRhauEMq066VhkWpx8
mph3XZkAa6wEJ7c70SOIDRJ5WH8qevSzvzMgwPYpeqHzXM1OTeihysKPSmoAI7Zl
xSbpZVDZd1bG4nZZ2XAq6gat8OfqGbuq/R4edKJNcrK7TD/7Z+FRXPIqU3v/5UMZ
AXJCoxlR7B68xIk9+FRbOB9faei7ce/zl4X4vJWMR1oir28pG6175qN0VS0X8JQj
/mL2V9mcDcIUwRxaziQ3x1wcmvve0hOKt6xElz7ESjjk5y4WUvh7n7bQ/T2vGvwK
e81y6bU2HrWZe2glhVDzLY9sYt/2RlNF2Zqnzn8bPvAUDSNxuP7HdwPb5lxLFGeK
c016SbtNVkyyKptmNpvsGAEShB3SLIg9XYrNme4B5Sv6wZ1jS44D34S9fJlc6IFR
7l8KG2uU0qJkboLJkSlnzhgM7qRQu2DTcI4SwHpUNiAng7FdNV6IsR+eh5GekndJ
nlNKqiM7yS0xltA4Y98UwnrXcFIteKSq0Wx9EYOi0voih0iwus0TzRUHvy9ingoD
JuAYkwsn2Dv/eaKIWtztBpdx4DDXsMdAClHeWpR/PwDBsBE6Tr4uFU55G0tazptY
ku6gT2B9fpelGN+2jmRqwMTXHUTsBPlJBgAzGd8De5WsjzH8jYO3V4luf5i0wxCM
fAoyueEpYHwwBU7FytTYxQMCEU9cPYbVB5t2Uk5UWxqBVfMHMJ2zLjQ0MnBe2h9g
9DipiCx1VoSLFX6QHGE3It/21Vp7T9nDZAmVoVVChg0Bb7MSq+1gFKBisijls9FQ
nJnD8ow6A7qjMTGnRT60mtloDJcCUNjb3EJxlPgT3gjP30SGV6LkXguvbw8Q4wV6
t0oglZ1uXqJGgi7lLK7OiuCj12h/5yB0JTzyFpCNLSl373tALextg8otk2msrmIk
uBcixfHI2VS3QunE034J7dnakPrLI+3LIneUGTF1X8dkJX+/h1bospYOXjmg7XoO
p1s/WhXWGBDQHEjkmvM5L8O5HnSDBvOHkZAKOmZu3fRXq1hXTCl7HBuIFhDWTJfv
D6nDo5hXs8it/dcBQTHf8TZRDr2wJt0HecnD1CX8M31MYViwzHIMqw/b/Bke0yos
zAeYbIaxGgjY7HfB9etFEfl9/9Cgs8QjsclEum+1ZOEuQlLbgeVoLEIVsDPTyhAA
cgVC/8AzfVn2zwq7IcJPqoifEvLrH97reSLtY2u8AzXw0D5n9GNTvf0zp75zeXoq
hve/6b31nN6LTWR2OH2Esu/HoBYRfNTYHhU6hp3Omy42c6ZvQ4EORjN6VfQEQMEa
wXa8xMAHx2J3/labWQnbmzrsTzb4/2X5Az65BFavdvjcdP0o3PQLo6lvsCODvXdo
mv3qMRiieqwlS5JQJ3VUFxwnFCHFVP+ZG49F/CJkq57QhqurDocvOL1SoxSeLjss
qkNGmo7EV9uKqn0Whj3smYJL8sDWZJ2C6SOnPm0SA3hSprx+0S+ZNR6blNV2HATg
jdQdzAd8lEribvQnCvvtZyRRAsj191TwDuyn1IVRkcbmG9Urr89UcQ9+gBQ7eEQW
duXh0K3V9/GKtNeh0qDQA6xbyLOjrT/XdD4c1kUAFKZ5nLPELeSh2fO8E0kOyPay
hGF+lR6zLaiB8hhvl7k2sANq8Qsjh0qaLKTw9HMpu9z/Eb5P+GXaEgCrr53kC/SU
cKwVuSFDAqjBYbhNuMWpebqwcVKKiWVnF0nCNDiGtKHGPsmZJNMj6hVFIaCbS9IH
s7d/FjScl1DgRvL/pRNXj6CyUCYQ8aKVYxoyU3bfts6jRkpNNkqxTvUE+yzU3u9Q
zBTITJ/pwOBp/38EFJ5AbGlDd6JcKLijfxVSCq9w100hCoDN6huwxAJ8q8ktLjUG
+op7nOQOBZw2n12PZKqQ56F66j/XBPoxf4oRll37MMXTkeBVi350n9XZocXsY8JI
ZFGr/TAbYstFEdIBg80ON7skk2h0USjRWoFnrDBF/u9I4Hs6s/kLmhV3oZws4kOf
Ywk8EN8VNHkwcyGkw0LJKl2f6WzBLUwTpC1YLGK9+k+E8z/S/+JxAtXSHk2IDNG1
mlfbnqIKMFMunyiUiUeKcMcitTsykW2nLmnKKQCDkroIYkmMjGzUC2tQTdlnKLos
LR0Puyv+9Vicj4ZdjdURNuJ7QO0CZ8C2+oZuI5cVmZkYjDqD3Zx6MM/BR6xyWK9e
+Ck3BMqltZ2Z+3sY7hWCc2C8DvurLfB/QxuUfya/TOtRFB0DhVdYjC059EKn2Bmq
I7Z+UXRpc0KzRwLycn39cEKm1rYCDMddTDm6/0NdoqQ+IAbP+3uvhVGL8ucxF3f5
SL5iT+4Q0V5LsoR4dQfne1f0bg+aJhg4foaNeg76W3zWM5cAtiF3yRA75P1kuV7o
aPCA5zGyFEMoqlgLcMClMtEDIEDh+w4554SzZ3j19/0dG52M4YWv0xJiShdG0zP2
HUICHfHtJ/8hk+2ErDo+OzLKKvnoo4z0xqNzsn45RJ3VzZbNYHRwFlUdMnKPeF+6
Gc2nL+appmk7QGUKL8HC9BZdbTYHeNvgU9XIfU76+lf/MMysBBWm+/cuzVLhfRZQ
/Faglti870yNMSiBfmGUwpnILueBwLlBpbN9T7ADkzkvqhdP9PP16JVu3X1SjVMw
8wuZwhk7TPy73m6E+BAQwff3/X4O2om04WMW0UHQDwk0/IyV12Zcztw1jfhn4LzF
9TfT35s110Fsx77epkvuZRmiOAAKvp9Puf1y4jAFVkfDLAphRAqg2zyFX4dDudMt
jwu45cHyizXq73ZmNYvpBs6uIRIZCTztGpaXBiJbfWIKO1tbBeRVo8NTWuIUkPs3
FP6UvvawjXko5EnVUKyFh4exoVAxKtrzayGXRBz3A5b8BITQtRfLKGJAyBn2GdX8
XAUd/Uf3GOuNKT2A+YMU9tEumgBVBJ8j/BrPA7cv5kkSd/4jm/5HRuJRLQOqmTEY
qXErKDOpuczl0teAoEoPY2HBp1I3LH48100pQdF7/IO8fS/JO/jQ0nmXCW4P0GDp
3oBmh2DBGnBBEdz4trgHIce3EIoM7JYpgaSEWWvD8AO6KBU2mjYLi3HX9OIrUTc/
I1ZGWWpRQ3naO44Stk+yOea/TM2dQ/y2EqB5ekKA1isiP3VV56GZBrM8y5i7Qh1Q
Am7Evp7yC/LfUzhZ+S7kZtmHDjTwImbW/oOo00ncGDw0dLTROkIRfc1lIeuUpgkt
VDyxDs3EhaJgtEWswkHdHWhJc93wiqBnU4AZECKvdEhr23TabhUtUH+0OiaWKE/6
1XXTVilcfFcSKJ4qqyXMCJ+EMJ4jnyMQo9aVRKCAJ8K++bBuIBjQ1TaS8E19WAcO
7ekvaJ867apzDbRongzgZQthwvL/DnlJOsYVFQEj+Rs05Y9X80EgZnKLimzf+y6n
86w98nn6aC7EUe3iBkEXoN3D7b+19lT4Si0N9I+hZheLsxqwxJ5WiFRPq1Xxsxn+
i6JVJMNEARw2YlTX7iJ9KLmSsbXBF9N9qAFo//CEDQrdtPAwodVy7WW4+knA5bsA
5rMGVg72AcoxhCi2P9+BqbX1Ax+xQSyqZLiARbE7Kc/150bwGHuNL0WRsKCCvBvW
+TtEdfGKOdUOgSxr40SH3zyJtouUFV8RMw9LWy5uMAhcuRig4XgrJKWNPRzTyt9y
HEmL7hTRLFi8CTJABnsFpdDpr0YJb9UeK6tmqv06Sm3bxe/j/8UGIvwitLEPoHu6
2nD0rIL6Co68a2IzNMdlkI1MBG9FUtw7xNKdnpewhhtt9zwfZ0R9HKYKa3IEHRc5
e6zJhyWe/7tK9AQ7sEdVTKGVLnLg1Ji7oZLBCcG3fucNq3I6YeeU11Ek4XZi05O7
gULZfnNgEnxZYrO1J1Hkp6yNe7wJcYNVhpsb5uFf37a4kuGYn93oJHXEe+10BYgd
59PUvWceTFY0ZMZ1DmjPDxcyWCVt/E7qkyjqDheEc3/OgICdKaW1qJhDf4XryjfK
J3Lvg2otoTj9TfHXlRNwV/9LXzo2SX+SNQtsAhnNbEreDPkw36ZppP278mSFWgVJ
9pOWPeoDPcmmvTwTPTOYP6v856i2kPKGhzfsIQJIsohGxQvVsG1YgQa65Al/4iJI
PDbd6vG+rqPgc9lKEri2q60TwwKH6L29L8fJT7TWl6fYsfzss4+X4rrLrF0brmzS
QUMJfCIWpOkGZtDAh/iVVNEa6ecxrWxeHtz7yNIIunzKLjJRZzXhvvtnk29PkAqE
JcgOBVXm7vLdNHaoMnNVeGADE/E+fFFylSEfLJFhpDqEq9wdPwiL+l1OxsmRU+tw
mHCXytsji9N21AStgEEvfYv+W9olhynkxuTmaJglzeGuIcRq/Wx5dt80MWvtv3TC
R1UCvPhokGgeZcLCz41NQkpaFnuVbXD995XFgKJyPb4nqyjIl+PNefWbf0hDCvpq
WG61hQ9sWujMmKO37wQN5PC627fD9r+FGTLd8PN6xiHm+iZ59DHRj8pH3AJ4mUvL
uBNWTtO9yfU+tVw9FTF3yie19ZD4kIbA7hWhd5RzY/EH2E/SB0jvy7kOlla1WyrC
U9ikKBxU6SFH2XF1L55EGmLSIExlM0iHIFhN8K10OdVPcCzWOWctWCW5InvYRbip
KyisG9UwCWq+oQlPMc6gEyq4PPcx8MbJugJ75rfAqsR/MXOeqCDVQCxBpIzDgGoX
yNvu6LZP1omtqVOtNKUWIH6FS6KmpVg0c2i2UIa4HRVjNSwoSZGcj6S8w5P6TXje
LuAxFH43AfLCkPGqCCooZMpS+sCTWrG8BmVd+hN8iJ0t+4apnWwFe6FCWIAKERn4
EvOOYc64Hu2tR+83eptGZPZEvu155w6KUF0jo+u4ElNqVIuAx0vKG7Sex5XDM7pV
gC/NxeZYfFlpbvfeLcIhh+2S7ag5bPe/4LtVZP7FCDYxMOyu7GekpHjOGPBvqA+A
9jCAzckbGA4ch6M3ojUoL9iB6dIm1RFx5wpMj6iuZU88m2Wosg+br1Rb8MlbcwGu
hjhpGLyZili84iNAlmemQ89k2KpXQTyS2STBbgfUkNcdIZgYleCeHmqCUs3oKK59
fPqyd1utMOH+5RyVo+my17KrcbUxn4UPBqYzSFiujSDefqhGIYj+/kKkPIlj52K5
y8843l19Vgny5CFeWFiQpQwCT7DuwXjw5zLRrxaNEOOsp04QE4849b2SvmwbPfKV
Z1xt5SlFFYlH5jUjvcKB1VhLrMs6dPaIJ+nfnzs7s7/ss3fNbEIBtSQwUUdrcFkM
/W1+3a8fpVe4+de388jt6os4CRQup6XYkteWSJhuGyaKIr3VBcsqTwH1kjmaoeib
uW/LCVVThjp4jAA6u38LG6BdbqTBYS5xPZ8GyU2HgC+BXax4sFCdQZrY0INjQRju
bQEltbVaPirAJZYm94N4KSiyEFCUpmrU6B1DhcR/FSj4vxXDvqfG/Yw7NHq4KYMU
U4wNSlkzQadS4W9oZME0hauj6j3gC3RUy003xFmkAtRFwxiFDM0oDcVlThfp2xxu
caDVgBMFBjCPhVWWoRoHVr+Q4euWRH60HaXXVOjuK2QOuW/s5Rdo4GptcXqRwPTv
wBz9SMhC01xIq7bgU+Nz7uDto+cqYpY8STd92PY/Y7ZH92rEW3KJYqHHSiCsvo6o
DU+xGbi6aNFoBWF8Q5dVOSFRHfZgucG5QBRCgN/JUBh8mg2vN0iYfsIx4TEnqhcs
kM1tm4/oABHHTPZqU8klmBcQ1f5wPozxwFSKw8PfGj6epjAskAn33h5OO1eFVzI7
0TdFCeegogfPb9Y12fvCCwyFp+7kZWXtQRvLy37t9mJ2dz5zIymnDtNPeiZlukNW
uxht12iLPDg3uVi3NEKWrUkF/TM105dSgYIGvzGpEbZQvFD3+QVHByHMR0OrmvKd
1cThH8RDbuQdc7S+09/0a6/xJYQylkG1exJ3L/jIzvxIgxrJCFAjhMZPpjP9ADFw
ckpb9LO4scIvzf89bE0fzzUVIbiptHbCKg7WT061izRi2U5NEtwKwRxzlXrfFooS
463dVIt3CZmZMXlfpStlXwpOWr9YTRC/Gkvuy/188vUf8bUDRm5d8W/gLeHwOJF5
2i6ujlmBPCDeZWPpkcuQLHOHU5iaQpVGr9xFchkun/ldJqc3fKtLUF9OTzBmyI8E
tgzSdhcKgXuZmKJMumVS3LrA2WSOtiytwGg0y41Vs8vNCwkxpnPEtg8Ry9ydhrGh
R3lhsPFJSQFu5PqWHQmFed07khUl2r7rbrWdcbBaskFalf6IrXTq8Ez01fLe2XBa
6tTiom1BCRpgTt0ok+2GLNrdo2t8FLaLMVeOGY0ukFvurIHHFtuoBjlEXWMr+s/L
A2UODF8ZsyXC2dVtYa6T6VoXy6AsL1YQq3TIWLpj7nytZmJ0vGqLChS7k4n90HXz
guDc4soHqeLggGILvHCemV9SsM/DAX39/SRJpCyMkeoZ4nlYvKSam9ynhYy/plTb
2Ms3/ZnAgH8kph2fPleTuoaJKVCrtrJLNCrDY21HFG1uJYRPjx5STMIPOopUqxl0
qpLxwsveJ0V4AYpL27pNZzc7dPtvkP0thm8oLzhbrYoAQGRxJN3pt2NSoTQUNVY4
EsDcwRIrU5Q7O+D32OL/pbyluPdJtIKw9GZRxDVu8LRWe27swQlLQN3XT9rKn4GG
fexiulaxNAasm4YPDKE9tLG6XkhtQOUgp6KoDgV3IXFTLs+G9ptU2+1aYMObXqxl
Fp5jdGQW2+/b/MbCpOBtRgzNJHZ7dn6K/ij3JJBxIzZ+ZKWWQFVX//3YyRT7L0dB
dSfLOxVFjxWei5uydddm16edYDmehmZ9iMYzG6AhpHF6MEdqV4VAMZySlgcnrzfl
JOGq2zaxUWSOrfqkUBclhveSS8g657RPJiGb53Puay64Z+W5Z4BEsi49caR6WEJG
Phrpw42GA7WPx2MMBCv5qDEhMIldp8cUWmD8AJXxgWZ3ddxEg7rpZ5cW6/NCGEsh
JfEsUkVaC3GYTBokyhyvqxJY5bEnN+Un3sMQEXz8SJswprumGG5gf43K/UUN2UMN
pqHT1c+izE9Znec5J/lj0XiaMaAYYUrd1LhmjLjF74gVm+Yx0EvS/4AHRBARxEvn
8Q+O+Fvxk+OCNyG568teW4tWcVqBTrRHL8elj2XXpLLRtCgmRx3t2B25dLgbR1t6
mKg3JR4PUqlrmefPMAPcbA5aZegMOV/mJXib81u2VC7UvmMS/MYMEU7g9c05c/bI
lkUjUo1pLySeIgL08OBEi9jRP5jHfk9Diwfc99KQwVK393uo+wrmFGxYcftsgbTw
okrxO5CANLKoIAOnilVEGLoj+Z3teZpPj3lgBcI7iyG6VOGNv+eqsgi4A+yCctZS
VDBwACE60S/RtbEYnCoiax9TcGmCAG2VNUzScBVYlsl17kr1lN5TzwLCNx84Qpp+
AJdweYQd0NLGu/sgJkvUaAAmhXPbBM7qtVNNN7FKk9VW8mzhQZwSaS2fsKIRmbxo
LJqeuHBfATGZl6cxIRJ3O/OnBz8Hitx0iYbiVsJ/yypMzQxqEccbeE83fQGpmjoO
4D+488RgY8rIgceaXOhHea4kOAj63moB/joMA9oovgUKg1x9TIR3f0mjJkv5rQzt
CDaiNY+QWtMEeLfcl3m2cwZv2XRnFYo6KLbm+E+IsS5vzkvsvYDhHBULx2cHssOv
ZdyAPMXtQd610XRa+9AMVmXLOmS8i4TyT82bB/ASPARCc8UME8F2Ixv46hKEIS0a
jvVzncSpz+RBoxFi4isfrXtdKC/lJnr/p1a0fuWgBOB2dBzDtZQbHer4I4+2Hezo
DOr5uEnIf8TRzZ3bP9gO8V+2AGEeUPqe5OtuTV0MnfdavGGBVpFp792XlE5mvVli
UQzI2LupjOSFraE1xGL/chzF65A+GGgzmZMl2470K6WWwSrG+FoA1HtZaXJYfTGj
T9FirylUBET3vaVa3c+QekksAZPb+3QcmAPpvwsfSqMOeE1sdTTpuX/GAEHo3SgY
ThIj2pdnNvBWuG4kpRUJ3nejDQwgzh/lZUnGP8jM/B11YwUfid1AjCs4MK4dpBC6
hoWS2bid4KvF240sqgsooqGW2bvu1I1jg6Shk4UnHp6hvIK3SNE8Obzv5RKbRwr1
ByLc6C3QBnRLiHWjZaqWQWOSG764Onqw1P3Q14r1KWO+1nZdE53try0yiEeXJCal
ycpYjMzvM2kg5KsagzkxhWhGgEMszQUCu2FzwhpAsfhTCtt4pVTSNXrjkBpd3pse
5jGKz/Oezhli+/+uKBuxt1g7NVRCTEuUHKQZixOze+8a7qJdjdOHjwNzhNysyoDf
HnIC2j57Csam2nkvtruwhQ4F0rZPbMaaZLS0KlZYMigXIdXFePf7zPRjP3q7MMcH
Hkg+QKLbdTyxGxke+8E9AenhjMaqawome9O2yjQahB4G+gHcWvch3lTy/dBB3cOM
aIZUYeZvE+JSo2rv6fkivQWfyUSVQ1VSqOxRctWPwRuuz76iyMJx0CAQiFcsmoKg
/FlnsmhoYMrGivu11dJvD8zBLvU3ePyVr6cCHiz8LcnEhXkOOUkNAIPx8WzM+qzq
1LrK/A9oVXlJiJXJepTjDAPiu8XzN1oNgiOAwdmawB5Fn4U4NsIpxnWRgSRLoM/Z
Zrm7IDa1j0zyXUboasnaoZpolHWvNnN5G1vKqZCbSgLM4w+5EAMdLGFS0T+2ltLL
VTB1WDE442K7KzZQ2Azunplp4JAjTWQh1u2MYcXjX85J+F+fZSF+iWBbgk/GT8CO
49FoFq6miwb77qmAzhGPSTAi5KRLMqqJPBFOzIzpGAq3iCR2LKOX2qRj+x50LqPN
PiMhgg8wKbN39BuPVcUryUXS+hVfbb+rzWDGkUIZ+9sZ0I9YaR+ZKU9CHyl4AAiD
woC7A3yew7mA2U0qEgvI81oarhLu7llM9oZkLv0Wd9sIY+Kl9O7XeOelTa++sgSN
XGhVFIBi1cxlc9sRGQWomXxCSiWDAWnqlKiwgzsvd6lsPz7WyX6MpmgfHk+/dgMv
xWSofRJBZKIu9+DMyMsWr/YTCtiBXmTdyngLt/VZPX0efffwdOsGiR75sIDKHh3V
lpuuZhpH+YdMWjQQAoJw2dTWIR0i3z8BKLW51CW/O9TPdmlCePKXZaZ/Qe4tJDir
xyAAsHABpDK14zia9MLNZxvpxToZiM0D4N1JGfVMNfUkwAgp9s4j/gScMLORsSjG
PiZ8NJKyAZlADABq2reeu+nOuzerLtWPyTRWHwoSu49vHhMmeCratk2Ns9XmHeRA
ymLGCi5AwGlHyS7MrWBL76raVMKrG2BCE8u1mRC1QUwIh3KyxO2C7yVyZ8dtS7zw
S3yDgdvkij6A9/A+XSsYLVZckxByDRMxlVr7ndZT0U3aCB0vzO9q6i8H2FcIjOoO
nq8Qrs61LZs0OTc36A7LncYtF5wnte8VvuIE8CETMltu3tRbVeRtBGzmdbll5/SK
URA1+6QBIGAbs03x+PpkEsq0YRZjQvKKzAsqOkliMuL6d5tY9Z/wDvfekO79ZvUX
znlpgXJqptymkix0AOJT8SoGycTa1TPPBHIDwB0kanivlXXCNNEx1L05ZtwKa3bj
vEtmyVrFtbZshyMu0Wkt8UwkAoFC885Uf3nOgYQ/jzxWPrG+bI/ERy9oenz6Bxj+
HZmIuYvUKaUCBpCe/ER16hkW1GcNZc27WrrGVNumSwExiYuplUkA/njvQjShxMXP
cLKRFpevORaqq/UwO3xApasuJOebf0Cw5AV/6RD3ZkQz9TsBYGXaSX3sIH5W44J3
P3+jj7AVnA/1hTv98LYMPzcJw+1jmLEYRxLaafE8Rfdf1XrUd63vpRQ7YKHYICbO
FpGUceAAYzEzkjwQnGqAk6qUJwGwV3v4gAJfPvE+eyrcpm0Ru3EcytZq9qNswl40
AlzjE1FfvXhIDHsuI0Omayun7YxFPzOznHu2MMcIIlzPqY6p7ck0Munx/qs1Q6Hp
aCrGQWX3jiAuDPTsJimfRRDgp5TlF14bIvR7Uw0epQzAKq9ZzFOzzYSN+We7u94f
fczXuyObcD5txT/k+iXlFLRp9x3DZBv26HGqmxUDvf3hXXgLu/Ay/f0P5kA0u9KG
/gt3oxXSA+WpVczcj2VUpyoxxY1lWwT1Gz2P+ITUBsNp7lmXXwxOktngSPzlxJVj
yHo5fbbQvFY4HSlwKn+L1VMLvnBjttlfolB9h3XEOjOFnN/NO+oQGwYla7iYlrGf
2qAwJrJDX9UKi5ivfFxe/lmMlfNO8BsqeI95ORU+9+0U+pzIObiOpKE2SWpTW/gm
Dam2IOpTO1r5+uK4IE2c+Qwiku0I7n7ucfHxjQm65DuZPoXPUE+IChG8jM6OFxao
sUNmGeDwr8w+/KWTngCTbrP+HZd1HC5TIHeDnu22FDWwX6FeuTG7TMKddgZFVNOz
CRNSOTbBIefY7iZTftCDc/BAZcbLIGWpWhG6/RR2WcH0wjfCmXEmEmiaNPE6e8AX
0qQyuNbfgjC/puLQaXd9n0wSLfRQEu7b5aE6ORQ4qs5zbfSkewlVi5+nlj8OYV2I
utirleVzo4sr4BcdW9H6m2GVbv7goNtx/qhW0lt1eYUUkzfmwzxWL4lVlix7AKVm
aMsFCi2bKMpNxbRTurNCd6yuHIh4zUOEinfcEIm17FPEt1Od3byEcOY5uVoC8058
VDq/D+LMVmDcz52ZmHwyJG+dtwFRomQOkPgZXHkSC1z6KXYZJJhzi31QGD2ZpSi0
0P0SFyzR3N2uJcvshYG50fIuC3HeIIiqPs31FJaTZc1Mc2uu/onr7o30nm9Zzckf
JgzovgHpBBQZqzZcAec3HF2BSpOKTxqRuBZcoWgIet8cnCAPaSo6Ms149onXlZ6+
eZH4MZGm+aL+KzEF4SpjsV2NB0uT2Qaxlp2VUrhpEA1mrh3MIERbtLqc0U/pTJsj
0k3tWcEmKorI1FtNsjBu8dRMLp+yEwVy+oiZGy/jGPtam44vtPgjxAaNADgWmX53
23zDWIL8K6fF+UO1zzrJ64aW3CqSekR1/p8/SewLEzJRfVY0TDF9ccxSZ+hd0s7E
7+5bK9wOf1F7jGLc++md3Q2uhc1RTRWitAa0TgyWznQ4S2jdkYiUjjxaWpYQ02x0
BS4iw6sotu8wLi2HXmO9QBLU+foC4bNCxKO7pAIofYM8m/fI6+5ZtrPSHwWRPiBt
XMep40n+xRKWSQD0EH/EiWOhWQ4N7xXhVb7JFfOT3IknoEwcy27jznY9MS2rDa6A
wepWqOCK/fGSvHgd3GksMJTviPFk8k9w9JvIM7qeXTBd7N7gNpH9eXKpCAiZmdnP
pDGIF9yVOy49BaJKFCEwUIY5lvsiz+f83lDQ+5Ob+T2mcC5S+Ln4fVHWeFpAAUh/
LyuaICalFYL5TK7l8iT07NodTnNaFp2Y+Hdj+tac8747k7CSK4GxUCGB9q+9hMwV
PJeRgBAWt32AdrgTUFvRWVbbPuANIsJopAY0sEyCq2s5P+jj256wL0qPjTWfPSJT
ttqOEcaBk2PoWSdbkBkcWuovKlBZZrL1KMA3G3WAP3Aw+8cYx4+soVJBjMGSdAZB
MqGmIfp53DaG/0qie3eqTyz5Hf3lSY5PQupyhguE80fj9F6ih/Oi7bjYQNTMa90n
ldIz1wuIJ+FJZZuL3vV3cmzkQUImWWYNvDMgBeunBi4+9IJDzGxEaFUkJIyYuu8x
tvzujFuwVxeGWvU9+boOobN38wQwdbH7uV0aVu/OM5SwbwHZZFmMz9j1T0onkKIw
t39O33NU5d4CARXCLAtWFwmRl2h4l0jjyF5WCfFonUwJbCDcxa5wI0ezpSkO3fIB
mGpA9Beg58gUzY6LgKZi6qH0q+pjdNfJuv7BNMN0iTIkuzZ74EWdd+sHBpLpVmp2
8IxVed32xJA93E7rauYqa5cqRqiLs7bP78Fu+bUWoJfDKhQxz5JOAGQNPrtetenx
DDokMxu4J0Fciz76Bhg1hCt4GGVzBDr9tIK89LLccPF0XyB1U7yx7xJtHC3pqEUg
/5LBpRv039p1jRH0ZrHf2XPsXIfysvbdvGLPLmeJBl8aHBaA61WKa7FacQHCTLLJ
7q4p2nQodT4vK0/KYreSp/DfIEBgxg8jaaeglfhO5L8nOhHC1Xe73XUwwycD1Dp8
ZZmSaDYywKWKWNYavR7PMlU5S+rPAszQOIi30EBlEDZioqsuIkRPSYUeZpJvcJBM
U/v1wKi/acgUaIGDysEJr5EFPB7IgA+NlKXOHcE1xHIkRYjEMES6FBHwdilpKoxL
5iqJZaUODJ4z0UFT7UqSU+b1IWsr75DE9OSvb5zOexurz1J1Sfgtsy+RlyFb6GQ/
X5DrSBtCw+efZEJI4wGADxTKPEtyXgStagSi7DA526v598+856fpU4fiSw5v4+Eh
WwuRdAuCTY/of684WiLeZ5qqNbjGLhFv9jCR8I/og0/5fA0XYYh3RfJT8lwVRAtF
+Vs/updtTuuALWC9w3TswzKY+Z2CslPnp15ZrFPo5GmN7ETfo3LRWYvRPDIzIs5P
bJobx38AVzrJge3ePcgYkBKkm3sFFh2r+EJBQLCulp7T6tmoVzoe1lTibmTbhket
1EgTI/Idqfir39KCR1uR0feHf6SeVoZFp9RPAdnh+hoKuLKHpWvlYtI1VJLH0YKu
Gn+6s5dCCWtyEDB9i7THRBAUyQCW4pV4B0sP3GwKT1KGwqkDbhERkFnCN5EGxW7D
1ovkvs7YRQefg1WHLhAlLZciJsRXDd4kQEYP39NXRmvAgNcZIAvEQvffibHxlW6z
pDZQsDTR5/+8u+i++vQ0tDKo4NgoKj30uHPcALzyv3K24rD/QoE4mX97Uf4ze5Fi
80uftAy6dbVBbNdX453Oy7M1tdb8RzxrBl0yKjD82JLfbDOwEG5hYJlDgYvMIVhv
I5a82tvaZ405nlPM7QB8DsIBVARS25njxyhBFKn5Nu+JMIHHivyFdTLN9cjNT4dP
6o5aJ2IvfvZ9SfzhfKekwOiKCg8DN7u4I1Q5oxh+BvIwUjU7IaEuntLs22yDLPsI
T3+3MHh6Cc5kvOwJLQvLPGSCiPZjWmU/sS12MgQUcxqyI5LNfxxRcHt2t7mchqH2
jjleLqQdKRQhZpedSD0sNK8XcVTNqCKu9XQ+/0p1donxbErKtk/Db0uZ3He6E9g4
HTwIw31NjJuUeL4xDmSjoGSqpOPfFXx3O3dm7cAUI6+IHD4QPjAvD/ZeR2G9OB/0
g1eCPFbLE+NcWBZ0SdI3VvmLO76MkQ1dqxEWA89ukbSCJQNiSO9bzs+bRmYeTEk7
WqgU0tkoTa19cpOn2VVoM26v2mxeTXb1mc2axVrudc70w0sSs0cuQfFlUJVyENpy
DpFkdRtJywapmSU6ddb9UVgP4ZAa2cj7NkbeeV4KO1ww7hHsm+LBM7ZveTtT71qf
P1IBWeFC87HVNw7cdwiM7PlXUPjG0ROmSlM9ft9luhTgzxBObyx1Un0rerA65mdq
MFmFlQXN8BSfo9XMmzbbcYn+G8DhF75qIRW2lf6j3YhI2mUJHiVFrQAOoA1fG6RI
nEqQW8kPohAPnXPiJDGdggK4UaHnohvw7YQLTvJJHwkCwEDyukxCWBPGtZ76M/d4
bGCez1+cD72Xy4afJxWgCdjYsnvk2UoNT6iJztKASGmOm5ap3VEqRZmRzT5yv/NS
tO3glfhVguPDr2NWnA8iLPRrej3PXihN7CoKA7apPbpOAT6m2hTEzhaHKxjofrXQ
dwth+/uzOcXTVYn7y6ipP6rW+0ri/Z7r1N+GqNIU5fEZWm5Cew6TNIcm9v0eBX6g
g0rzQ5bnngKaNUyK6iDk62Y2ZrbkniTcCGNwvUO5uV+S8MKDP2MZUBkDeMekszpv
bHn6m0YXYXE9wS1eLVGqZiGSQHoDYzCu33QG64zZFYmfyoCPrVeELldrn2YyHr+M
2LZaf3AZ22a3PjWGbX0icKR7Cg/bS8xOFL3esILwpAqzRUPKAwLOtRUz59ShRN/4
SjVETiHtRxYO+tV0e3xlr2N6rOSAD1ZbsgU4I1GtDwoWFkeI8lKB1jCqjNAD/9FB
A7jpPRercK+LrNgObHeATHpvLTRCEaMPJdLiL9AkTRrpp+a16ReLrOVgcNP2PJcf
0CspQ3mqROdiMBLqRHP9xmvVIcZYmAdo/2YOEglPzzfNDqUs2lDoBX8J5pMe5M2E
MmeUGrlDw8K3grIKHcS0WTinmmMv31tUEhbPTb7mpwidmhYAe97BilK56H0LVGto
5XTwvlLjE5UEgjB8KbwJOMFEiir6U7Qg9xmQaWdjldfFt5OJPSd1NaBVLZ5a9UMZ
+9tAasLQ/7KBlM9KVAeuV1TkzBGmHSNcO2iiHoZT9vmfcrquwkTdQVl6NWAdIkRO
bix80HzkDkAQYlcBROIGdMJMq48nYErPEY+UQC6MZ8TvtWEMtNNcrpd/WSOIQDnF
RnQv/FlwvW7ot8uduhJCMUeo1ZNkNRxLP+z+jTUhtHKXXiW7f9aNTishrSJB+RnP
zeu+ypSlxZT+xxkuFtG9wMDtVhWdg4farvKfqCWNSmxIeODpkvxGgkgUBNgx9Kyu
TcIpfot/FtqRGFgIkkxkVwqKh7ibYdByECSNhhqM+rUus8kas7x5KpbQpjbL8Fp6
dJof6TPCNpFVTN+LbkBbyn/7GWCeA7NxOnpmxCfwunqDPwStTPKCdBsc82lU84t9
+vIVxtSCt4xzuFOpRRqkBK+KFLm/OTQXUqgRJO4dTqffbUiZ9x94kMHzZ1wHk7vY
ueGtS4FBd5F6vCO+N2nVAwaqdiCl02lEjLTdYaONe12G+jzO+Rn8VOUmoWI5zDKc
cMavE3d0+qYBjGwNzf0yKC+aD8OkKypSF8K/iI4rsqPj4CH6kpw6+LN5LKCiDgEV
PYWOphCdqicRKVew564YSsGA5eAaVaS7QW3Pprerz7M87gsBfggGSAOzy8kcUHxT
eFa15rURItRs7cgZPlqg2pde0W5Tn4uR1FLLCpmDCW1LzLRERu2TKcVueIfF3uno
B6wFF/s1/K2U0e8ESac1sygJd5eS313l9pWYXf8sNuxV2YYoIyCUMZCGmdqZ/lYB
k0Jw+nB4+C/wT56dPhyomctQJwBJhGCWBpIZ4LL8/m8KUpQty8YTtNI9khVdqh8q
7T+vRm8J67pjZROHc6oiFOSLQcGm5zS15t/aHXdcZpH1CUw4DT92rKVU5+jOfmP3
7FBbFG9cM70CBVIrK1xJeSIxAg24A1DLzOqrkOaCkGbDhuap1LAPPTmKPUi8Ku2o
vkoHjjTOze+dysXbC7jiW/zvf4GuO8B7Ouwdk8LwkaTPnWw1tjXFqcoEMlhbCdzo
lt4q+1EFhxvsn6683HKNQffo0GRv27jVp0/pb8W8Fd+bLSP6QpKE59PyhCHFIt19
VgeOn+e0gTJynjEvPtYbH01D/957jZ3n9d5hDK/kR33ScKvhrhazTqCAYCnIZrJO
ZMk78foSayVw5s+zjA7pL8RlKJ4TyNr3FCxE3awXlG441QWVwEuj0WwOJf2ws71G
du8aoEGXs4tTHLM/xoglDUvAcbJtOc6vvyoc51x37GDRTi1bchpvhtI/y00L5rLE
cs3j/Y/ZmD2P1sV8vZ0FQY8ST2aJjqJOVXK929ix73rjf+t4Yu6hF8XB/UU9Ik1y
teARO065n7VAZtUETZCz+D+HzqaL03c7eR5spIjQLiHfi89JTNCvG2Eplw+twH0s
pUgyJBWgk6SiRaT8vf64fM5CFK3enSVVekGT2Rn2mA0rBSWiXKJZmJMka8pXgTkZ
nOJZHvSEsArYWhVN9zpcVspO9vewKHtnB2BSKHKTcWAykComh0qn/Y8cdRtwglK5
vVkkTibPLgZhKOaIW3fmM2z5q/5IOW3tzZSBlW8N+BdKAf3iqTttcGhyTzhYxC2t
xK5f/nY48S6uOxiNctoqUKVSeRCx5hDvt2ze2C5bDd4tWGMbUMBtt7UuWgC5KKKa
qf3FHClRgt76DTzNuHRs5wY6dSuX5Cl2SyhjDf9neRTCDE3Cb90OFgWdx1f2lUu4
GbBLYGDzYj8BZwfgf8/FYQJ4Vn6Bb5e4taMMlH+bI+Shq0fv9Z3qN/kQneoKsVXq
vWi+4fk3iIPPCZ8ZQX/kt7oCWF1WLp/ow1wCDa2nAa9hgtVwhHE9EqX54e1+XOaF
A62sBXT6JQkPuqxTx6O/SjveCXa0swPf4+Q1+HU0yYP0lASjgGBvxaqSfmssSsYa
Nbc2JdPI23aSzVWbDJ4pdI0rehGOX+qVMsvwiZqDWT50m6QRVoiJh0ckuNkSuO+M
KNiXkiSA+1NBqdfL5sBVV4e+qFdk1G8LIP6KA1/xD2cvZUGPVdFx+A8MU1nq/A9f
0+ZRfa6u3PH7pPj2cDiZYYpyCI7GRlPz/MlFrn5dRqN1A+VQU1uFOp65jI+mhxCU
tmDr5idYUUGqDXA3847pFTkSn2s9t0DZen2PX92p1t8yupXplH8nC1Wo1E6RPbIQ
yg0+0B30dbEwYoCqEFSF2JQRlACuU706sgolOZM7unRJL9NOfOumv7bYjEZvNPmb
O6JQb2mjZAj8e25YWa2iMHoVWFgpEZByYx0raox3JG1Sf8vx056JZJzL/AB2HUYc
aw3inI8joyU0Jbh+IhDqs5U53T6gNR31xML0U0ynHJIfmdbNROfiqk3u9IJBVhXO
j2LFpu4+eYS94b6yrhTgV4vc8HILVPAXOzUSF2w0XZjROd5nIHuiqmh7owSPQbB8
UGWaeQA4hG28bly/QB9EaIDKILq4PipAS/Sk0OUicltBEd23SzuPLKsdJ5JMx/5V
H88ILkDRHtbwwe4jXhQ6X9Yp8J5OpmgMGqW1sj2nuw66j8JuGWIvwbYwKYv4M1N4
eeGgYWaM5ekPThvsUupvyjO3NMCNV1AmP1OEDs5oda/fdvYaPHdvsnIq6AApPYNE
eyoQDeV/shHrqpfgZoDBPgFCLng9bHBlh6sntgPrmmDfJ+J1i1ccp7l7+wR6mmM3
/Xj0hrJGgQODHXShtoZBrdXccDGDX1VuhnpB2slDn1xGiR1tXv0hjT8oHizKwWUP
qDq1Ve+uYnutXN2qN+4mqIwVTuQDzH2d+k2ujF005bAZY85aetfRHXTeieKZUSAH
MZOg/8nLEVqrxb4G3kS1Jj5iWwUTXJ5F0cOf56cMilgIXiJNlilz54E4+kYUJsIn
aHTFV9e8/dk7zLcQefKsYT+nmqBBG1YVDy55eUOyjCGU6JR/Yls6DYFw0KM4SAwk
7rp2mc3szSorfBrjuI2Hr2aRQ0Rn6bIuf3V8eTvUZbAEmmXFLt+/Kz4G83W1PO4O
U3T3d9BViH2reb2t5akFuOvcfcgWpVZheRUwuKW7reX/Qe6kL7OMfy2B7XwHq9au
+CN58N3BljirQXTr99uLc6zToD93LK23n2SWIzDzwvrFOwXkyRgSWPfFnZVRlJ7K
1alzT6I3Rn9v9KBbk+Od9ed2T26yQVo8w6HCaQZ3A8C68mIAbBfIjtwz6lyEGDUK
ulcsyQj4pRJ8QQmeFs3HPLWz5WlfULQGRoIXMhuEVbsB67g0YhF6/idz4sihojXF
qiwOjL/EAIvapVOXmY3m5aX8K3wwudJBg7qBFHsZFPjbam35PLLM/QvBOE0reyv0
HgGSJmnKixHklkN5yk0ufK7murjAAgC93DmuXfw3vUOruD5jTdpmT0kOtSwef4Tv
D+Vl6KB7YNo/Zzsp9pzgoSqbod2bRsVjnQJzgY3ulmhNkS2tdhz5x1mmLwlDJSk5
FjXum1nmnhVRSSS+Vrk6DPeD5tg7cJGqHLOQbyRo6+jAubiOKP2EggbELbio81o5
CMfSZSrFU7A4Vy23XgL4x+sCUm+JthSdBepMQvF+4Nl0MhWh623W9OPOJfGAPL4H
GIgrSsrPRKbNjNdspJNQQGHrsCbEPQi7vG6FHMaGAd9KCDwUwG5eao/st1vRs4Xb
4tbHYbiejj4iJTl7Bs832uCnwhOzmBksqHFzSBqPxu+e9EWGCMa1ScXDwUfGEcN2
MOrDDZoUsdxn52KjB2ERrp7r15fEd9cqfHRMcB39hu7EocGpQHxUKtGwhu+rSmCJ
feOPZPdiCo3/0P8TcG05izxdCYKNNV7WJhgMXHTqhYpSXmOHB1F1lBaao42PCcD7
bAIoGzjAoRBi3hX2KUYVKO1a6Mih+c0icLZDOL7Bf9XDhLk+BR08zX+BGjTt6O6j
4g9mWUMmkGmkbHig6u8tbGL0vdR7Ljrt4IqyN3DxYVNezrUic4JQYFyCRPu5P/aa
DWY0Tzqua6hDW/CSUyg4jviBrcg553531ELdOnTCYbsubXoCWeHCVHQD5GcSoBTt
G0Ts9IrINCLUU+ui4414WIZaKvL7mpev0ShpWDMabjZuLus0Gk6q59ZXgvTyveq1
KUsVuqrC4Jlk923y8N+3Q1m2ypCg2xf3HVcxK274vtyUo+5zABnWYedwdKPcnaHZ
QkAMk1lia3Of8pNOGxAE2V74fiG8IO1uWmXDmH1ew414L2abgEnv5H6fBgrYg1nM
AgtC7S9+cfZJruPMVYvHix+gV2xvAZbIOsj1i7Er3W/fq23ezZtxJySnGj0KsrEX
gEP2dZI4p+RGONz4NVp+moVkRkygcnelRe/plz4kf4xmR7QX6FWLamDYaCOT3+I2
p0N+IAt/rRuXS8y7A+1kn3IM9CttUMmvxDrfA+349FiemU8F73wfPsCTruU5ZCef
bfPiJVe0FTQOpgBf9eyQb1/C836p9U0+tcuAsBr25T4hJSIYUt7NfSmpuYEg97G9
NCiDfa4Pjc+5oR+pFkek50K48KNbab6ODfAbzNYgojqMmWVtxIw0k0c20II/8O7B
3ZGGxzwqnICPNUdMPGruQqWJ18Rhk3O8tdxOsaT3eePqRzxYEWEdfu2kecSXO45z
M4+7zJi0MBkG7/XFlB0Gmp1Ugo5N/IZJy+20lJiXohFw/xO7SXp50RKuKoOQsVos
rh95OWp4qvhRVXNKGALL6fRqrdfGJWua+hs1nB4jupEsCwAGxxwHn6ra+np0qfo2
NOXhzHXUt0oTAv2k8YXVIUAriLx6Nwy/9+aGWOI22uZvj5NRxTZ/xCuf/pWVOjzS
U90aS00f0oxIkW2MF0GHOoDByOcRFrmmL21K5u6HM/Dpepc0qJYlELp3Y8peQAqD
AhlclYAZ3W58YyvzvlvtOo5Stsln7UrqpDoZKS+hD4oMC7eCcMGmYwDs4dk+Q0HM
qP+mMMltfCHGUJJKRsXHDLVvSJk6d4Wln6N9RrngoTkNIx/pL3xwpw4dnztMnE6w
cNCKQg478odyln7/EhZir3hTq2Zj+/8k/jO50nTBEyEnCkIiUnGz3fgzHrFF2Avw
RcPqMo60w07pWTEW6Qc8qJ2zqXOXmZxKsa8l+dhEH37vRsU4Fvxr0T5PKh1DjCul
KcdpmsRpeeLuX45IK4a6Uw7VenNfpu9dnL4xvgQBbecjKhhZwFr5dHrxCy43QELE
JBS+SWBSvqB4kWIYn66y8REVf8pN5g6FwApaD7nDy344K+Ib2kjntnYJ/j6uZBnU
WGJWoQZMO4e+AOjq/e2E2BQdlW2GXwv3LPJwXxEXp1/6v8JSSsGc92Y5PhQVvUHK
WeNb2PAqBPF3tggXvlhIAhWCyy/4aEdSNYgBUs88Va+Xl21nQ/i26q/E4LaEnK3E
pmShy2Q6+ngRE6qErxk9tX/1+6+TU7u5sPt1S0xJ47cbAwNMHfQLcg5E6yj/xdvW
WlTiIe2RsAsttlP1FEvlfXB0aiGOKqYgGdhdJD+xvlAINxGiDd4aB0uVqfKJStma
BNZUYaLfdE/yE/o1vBGb1g3quk40Q7ouKLnpIZ1mJSs5pBTcw/LIeELRhCrPxgKK
UDAnjeHcNhPrH999v23nmiZ6tVG1mJdpA5tlmmi/fkuvBp1CRA1jr82OELnIdqEM
SCZZtwBzvMeunWJTzBCEx+VWxVpJyy1Wsz9lvh5O1xS1qHnd5pGWm2xkLDaTSHol
oHIj37xdmJa+FV79KftMPzCHb4syIp1LOaZyUoKlFhrzQ4CgWYWua4uMrTD5lipr
iF+ukwtxHfOFiU93OLv8UI8bPDF2qgjX8Ij377nn1pDDKvkVvt5I9ZPNx7xZnc5V
zQXxuiIIQO0ET/fW+OPfzFYnyi7J+r8fUwM8tmoIaONgcVBj77Z6q1yYiP7AvHDl
s8RfVFjGRYfMi4zajKCUYemmQSkqJA8Ncj9FdFXge+bv+GVJ07kR7mG8B3o6/D4q
DuRfNFVsYr+8vQZIMYNAD3IqPBkn8dLX+lWnfra8RJTAAsTnC9TmcaR9bEQYF312
VunHHFvS9K4y9TO5v2TUJIvsoGk8Ot5NFHhPK/UGyQaIOVYM/21a3q3d05kn8coa
lNwY2fAs4MCSDlyfnnaGsJIK1a0mCYJGsuB25mSgGTW0FnQSFhpjTOv1Ro/LZ/Kn
rxYygHqOpbXan5qd/JlBcHZAoLSqJ77U/Z35jJdBvLB5niqRy2dgLmmsLWXgha7L
WD2nPTwYY6MsA2+0Dx+toBiAm0/0sPM1ALE1CjeYoggxT1rz+opmrZpRKfJeQ7yZ
gPxLk3ii5Ugu3+W8JRzqJzn6Kbw6CDzwDusTeZQVBdl5hp34wQNyR3JqNciILGod
3fGAVJ7FesGYkxvVTpibC+RQ+XXogG78MkmYsNh+E0HhU8kDeqsDnCTdbG/Btbpq
XMnLZ1miQlMN0i5UXPluW5dltdV/Ic36GyQkBbesXLzr3wKzA7xYHVczkfc4wSBM
dG2qCyr9uLQK81S/WUlJsFTJHp+FuxMV4QJDnEzKZ5rIjoGcY8pgypnuDy1Ewwqv
XSZVKPUcEeefm/CexOcznBDVcgytYwDCmszUxk968b9MDUBlUEJ9GpTz8YXAvy/K
CqF3775N/mObFdtzgvY4ij7CJeOfCKyPZGL+0e5/J1OIR3ZmofnPwYR+IEPzcs8y
oK/xu/NZLwUAXJ9bjFZfbzlvocie+3m/qzCiW85uM/v5MzzFD89L1IL5ZGhcC4E2
hX7EadOsifYqRujsZEcWWnqoRsTqHYJ5LJYnl47AFhnyug8pW3DygTvxkEDqAbDB
XMbNLG5kUfW+OlN4o4Oa/ME4PE93O4diqhnmBlF47O+GvQIhzSCmZ+TWUa5ecCJN
l3B+MGWis9n+G3qUU1Ar2e+mK+qTKNcJxmDi57bXi8Gf2D4wpXKjXieSlk8lsREU
SJUPz41VFlVmafVRD/3kkuVTsKTAFto7mXcu6gcN+FuTOlJjP9LJdXsv5E1AUQNN
R1mV7K35D/ZwNUHEW/j/yRXOzfCaOpJMn2zNiL/cEf5emWapyTQcOnSxUU5ovv+O
/+Tw+FH0hVr8CsFG2NXVYUSuBASJlDJ4K9FfsohLJkpBtyn/7X8XnDLAhLV7e+Ik
BuhfU5D9zeUV1z2akkD8VcBFKBB92i9x/gUGjY6rSqpSFnHFZiZbD3bHSb9dQXXo
uq+QYpwJCWZ4fuRkP0ZPLrh25MqIjZKctHptxm35TPUKNZ8VnspitoDGVXPd/OcN
7/EYO7E8zAVpqswodEuXIOOGIzdPEupDzWVWsL5BLLglo5slVmJ67eOPRcwcORa1
QTRADSVngAe+gBsZrsJkIdPLdDT4WMDVJP+AD0aD8YdiHxDmL8Yfr2uzapnzz4Bi
ObOGGk43gUYjVb7aLivMyZXTFoN0xY71SxioMZqR+F8JBj+Slu7llnkWG9EDcK10
S9Ag1CPLIcaMjaO9oXhkT+Vc60MZvbAGQXE6v7WGnL2L7pYERi52pFbeKDQGjK2i
9itNo5vFk9uTtQW5JRBklICl45W+MjGEiGnX5EaOHqa90TlMBgqpCaj17HM5BdxT
c/5tiM0u72bPxyyoZMfOtVHeKkG7Q2UFF3X6BkjVXtM0mGlW28MPPaqTaTaDg81s
RNHQacDWNZfzl4wn0O3XKzlD8jr65ZobEyP4SUyRx4ZbAdQbBEQwylNnmv8nf259
i3j4Yl0wOOtQlqmSnfVQklWh08LoYrWw4ZgOrB6a9QYcefVD3louc2R201k0N0cT
7im9/PVfFWLxpfsA6kqMshHdd7DFr9G9vLZXxr2EdIZ4MKJNnlApxFHOLDwRYnuc
VfWXBw1x1rg0ut3hMKpVE+KajtoXZIXu6fN5I+VP/IlgsTAJqySAHjU/0b8Q1B2e
5ceCZnblAbQAMzBO2UoxeXLd2rVuj4/uRWRaFIshOweghTNnefa/NtQCWdVzKwLD
DXXuSRpfEbeoVRs6sfjjoYa6sgSVr06ae8oFt0xulG09q1GRiiyoPKcI9azVtjzw
fv+VfvLDn3SGiEcWRzbUskt9iDb3qSSWtH1q7u/3EOoDkVS7g0MBKlMqkqrpfS5J
TvPo/BEDUkcTi3cDt0tKbf4LoDF4H7yyehsz2fl8ykXyIxaoUKzAlzRxXnw2LGEo
IdjPsY716ACIy1kOlyyLFPM0xA2BVR/rP4HdmFQ/NGMba3EQo7h6+RtRgUEq6D2Y
4vyTg5eBiwXfykHRuWm6TTZG+W0NZyQB/RxfyvWdbAHHOxAeRc4RW2lP8qHi42c9
a1lclzT6vgH5PtzPikdFGio3G1igDEvJ3jPREpwHUY9+3VtWYyKOL5wVAdlj0izq
JseFOFIABiC0T9LR5Qar23sJfDtnqxPxDZmHNk7u2NSDvsQJDOup32gIqxNOP0S5
DnY6hh/P8x+1rr5GK6JHsmDQtUtv4Kt/ruaA5IS7yhV+oxr+jKFUcQgfMRfdc6a1
bARuvEEAlw/1cjmhacKDHCymeZL5dvVU/Wpvq71T/5EIaOJZ7WoyjcFkyq6gMAoT
Ri3PI8az2lbldEIPt8EtVprJjNKrLfjDwa4Jd1JehyElOBfmSEPepvAimVR6zk/D
s3W+eQrE23TMqAnyAqEzbEODUIMlXsqlqeeAFtej6XtJwr//1iE4eJ+Jxr7A6wT+
lVknZ41+wEI/W5F1gRTdXaYe5YEmuP3tzxQSgHquEPz3ann3VAou5OkRQrimcPD/
kTa/AK/vdr9ggu4un5GkatN8rbhzLAeRfsPrVb70b7LhXKnVmuMyN8cQ486x09NB
pJG2pz/HpIZFiRufociQgKFVzT5ZK9bQKglbwK6Mo1RLIQLBqoqzwmp33ZaeFBcS
1gl13B2998Ig75oD8FgQXgY6Y5UyGHG0l61ESJAsKuowDhAtICT9ybvu3uLPYth0
5E7XlgD5Y2StI/la8RgOwgHnrO5Ncq1Ado92q2Sk1+/VLHFhkXaDqPd38/u1qwMG
WzA7K5jKzarvAcfuNHvJYxg75hjjzqYr8H5vBiSnL2w42LRlSE5pS7Lr5gbY7Eev
Mrnp7xOVBIIBWVYvnGypncpYWWOwk/XCtuG6S4BhtsGc234PVQ7I/vhrDE5eNTeH
pARCUZ93tgluhAVjfvmVw+Ac5pn6m0gbkz9a7+FI8fTIPRj5GpncmZS/uM1FqItA
gskrJ1uRzysCqXv5oAmgJ8jEcMClRBxbjSIVha/4u1UbAV75CTLMk51aGX2f6Ix3
NT1ZD2G6kA18ZsYQ/rtjC3vIQbigrwaWQJx8M/L9niwYrmlsR+mqEcDD6ZnxKKNN
0uLZgguWY+fiI3adTY6kivFBfYZVBWKsqCUtZUD1nS7ZOBy22O4xTfKOwDI+/BQ7
FtRa4JMPJELCvsoeWC4KAokFaZMxgq8wtMeTqEKA8suMax9XTeE7i35lsOG/3vwl
dbVmf5yDDDW0/ZykFT/t/59GQ04/C7EL1OnVXCZvi+hkAkiowHxrFFLFtFgwPPZu
SJX8e/9ovqJlQsq13y0uEp+GkKxG3+jnFC0Lzw4txxMSTcNJv4J4PmWsACruVY+a
fnY17VqgXkB02cgQLL22EifeckgnGRD+TJ4F6Q6VodDX2Z5yvWPVovmHJwGX16C/
NQZ6UvIHpIjqLjTuBvFREG/XAUdqQHNDVtW1r2wgDDa92OPm+ZMUWL4hEsOfhJAT
5g+GMFXszlHm2uVtpDtwr5gFohiyOESQRGUYn6JP1QdEDQoGoa9qd/7rmif0yGFJ
8hpdPrPxaAeel0+Gdw/uY6MWI70bznU8yWxEznhz+dn1RUzUR+Ff7sOq6K/m/Qb6
8EfRinRSW+xQRqVxawkvy5JCaTrpLGKJuAYT7UukmyKINSX3jo6s63NyJ9IvtQC7
2xLETRSLwO1YTjrFxIQkt22LFmHAGzldil9wcKWVivMCGhIFv9/nSGqTl8ab3BC9
CCxdRIlDZo739SqRxVYnRJrgwrznd115TzvmbOCv3BQZSHlUJrnVGNxvzRFo1i7q
okLH3OhOwlQrZoe9ZomjmoNjrL/pjs1Itl5MdwdWWcS2ZlC9IeZ5mW2ZPmHhzJ9O
aNvqCY0n/Nizvw3VcKHkSlWTrF06v8/zGeJUVoDRs4bIcbL4MET2somE0YQ7qyBm
3MLGlDTvMA1BO3GwOF+/ho/gxkEJGYvhjjEoAbouUxdZqhEgzHMaqh2g6T0YNUqY
l9jlVSOVrafStWAXdRKAU2aHLDOjSjoD81u0CPKg3txLfCvP59jyq6/vXNBZtW3t
uCy1I4Gpis0FXt2EuDq18Zw8IAaar1/pdchMvFV/yYXyrcMJ5oDsubhMxOy9KSZD
Jm9Kn7ShHgcbev5bGgCnp7ck48rzXjMce6EngG8uuLYuHH71xuJ+RHdMaM0coRI5
BWJ5RLCAis/kiHGjWPBeg+NoHk4CB/KZL5rBPounIRTnJ2ITb61Fh3itQ1QByif3
RMsQfcilInQrSxhdNBXsC295+Ade3DRolQGq18pMG0OEYf6PhB07Sk8P0swIZ9vc
H90NxXrMdBvTPAsRlNa2HXM8zPhmLH20gbz+BPvbJOBnjKE/yy9d2HQbY2VJ18jX
4cHVMtfd/Jm3KJdDN0EctvJwBz2cRouBd1noS0c0gPM2kNyDeiZC9tna0ERQ2H6D
L29GKPNmSSzLl6JV/I9jN5TI/ZVfc8A19xe83DdL+s3Jl/Ek+eIvT9o6weQJaDF4
VAQmbWb/VR0+YOFIw4CIPL/hNRM5+GaoXC1VgsswVVFvSvI/Lfq3qKaZSuvaGCFc
vf09r+r2TCqwdh/EkiSVeUbB8C7RsdIwYWJVr+Z5a8KYUbyrQARNqw8UJXnfBeun
NZbWck8s4Tbp2ZxOFsKwH1Lbl2iujUT9eqJ1bJAES88kRyBN7QnL5/bXfX6UkTZn
RatVqRAOiOOJpP3nagJ2C0c6UAPbiJP3ZQG+YbtuXhNkrqQvKPXxsf/E4bevpzVY
xsA3gJ7chYKsvcoIQdEePbenUQTDuz1/pNCvFsXetM6JVBkRnyaJATcd8af3hCk7
bc1+mpiAt2w3HOqrescxH9z2dfMN6km3UKayO+IwZiOZ/DzFWkuj6X+eOaFlpdXH
4gb3CurZ7+7jaBnir8u3kiOMzoeWFQtk7gwXbKx5tDmpnFTtHEjag5EMbNy+CgzT
Vigt64uMJhUU5lfwS+bakJmNg5TC6XxlaLZjPt1kZ5ODzRgqAXqUKUGsOmgu5lpf
p1FDSwVv0XwLV1FOtbvSIw1UwGaIGkEAG22tnHbVi81scv2bXhIpFJvuKSdOQYVu
jBY18lMkTaQ1iMVTehWpGBV2/RCLttiLyTdIqks3BL1b+ElR0yCrmAJehHvgqRiR
KuKcQIByGwCVRjRKbRojBeufoWXUDTLmLykvjp319sJMMHBmDZbIPHF+bW4i3txp
SNUdOeKLgJTOLEYFykO5bnr8QsqkZUDHNvtJA7khsA2i4g8IUF7Vv418691mldAl
W9fdBmzcCxVC7Np7sQhNbqmLrauDCizVZBA/EyWNuNNoj5uk3F8XBmZrFoxIbknj
bUrOC+mm7OdIJ7+TLGq4N8D1xPFfasVNCgwVm01fn6sb+zGtkKrqvh7ylI5x9OwU
R67Ip96WjrxwSpoFMj05PGc9dSReDphYUWcn7iE7BJ3oR7dRTzPr71iQkg428djW
ae8uZhsIUsYznlCtckR1NmMePhcohTY5V2iQnCjkN4CXJQ9jPORa1RXaahZ8ZEkd
erXkwjS5DLPpYXz32GNVsYVgy6jo4ztlAz+Jew4Quy6WwIvxNYQZQHe5zNw8AbAp
cBqO5eegnwG+6Jz83PDemNOiZTv3Vt+Wjr9Jbi+OGMznnhg3u7OKWwjpk3KsH+Lq
T9QfE9z+14BGwoGQGRYsn/Oj96xb00dqkqIvXM2CyaunX9Z5XoAY0Uj9urPLpID2
ZrE2tYim5p/5W95qe3ctLY+SJL9ij7OFqEfGHgkDokus8ilI0i5YlN/gt/XZ1iCE
UodODXtLj+7ET+JbUq0t49Y7zRZHQE6RKOSyB5GH7/r04d+JiOCJ+bcd1OdLceUQ
2q4IoRIFnUNY8282F4eEK5xV8mYGdXo9azhnND2MiEyuc8dEyCIzSKlbZg2ziwdz
b99G+oag4v3idmq/awKlBnqNyOmkQmCSpgCeDsLZumC7nr1pxQFIORQv/Ac8uxMD
rB9YLhEi8WZrGrxmyV+i8f4wAxNh/l1jJbIBi4Fv4FsmLZpPZAL50o4ayOeWlfIf
dvAEUxBL22tCNRxCBaBpkEc/gso9gdgnWfyEs2RQA7S3+WYSh9briZ+lMCE2VXiM
UF41qXoYpXEUyKZqWa9MogN++N+VVVS5AuZH7Ehh8ruQjRUnGjjNRRpaIh2QQ1vm
//lMSi0AlDjHEWjDoUnI3Z3RZeBuUXC3veLMM9zg32+DDQkLr1zgde5Ut2vM96Ik
O821uLtqLMT4dfBsFz/wLlyaVS3Qwy8lbAU0gfYxRfWRTfwYkYkEO94r6KjjHEv2
OuFX4ckJ13eMaK1e6YcCGSv4iLFQrD1LT5QUMj8lBwle5EjIsW1fWhogiKQrYnmw
A3dqBa0uqRqCcND9hYAgVwfghIjLvYBB1YBzROW79tHwo4epDua9y7Kt1z3QRLbc
3Bg867o9VbnMSuPnRDGD66PTdLjmRaZkcGPc+vrhJAdXTb7lFr8VBO42Gn/EeTO3
rbo+LP8T2U75SeQNg3pN/sy5d8F+1pmM+u/mB9hmnthB5e8hmvwrMhECRlXum4+u
xhBMm15qo6PeONkgmR8oS/qEkIqOW5V25CUbZPQCRhUKVZkBczH0umaWIMN3w6Xt
vPqKuJxPfmhP9RCa4u1EGRaDGBMupB7knDT7KtQmsnufvI6BNNqqniBkw6S5dkv0
Stu/sfDrrDZv4S2GawiJOqVtDfuvRd8cftrSqJWiK3s07CP8SoDe2HEh+2003iCz
nucrSsOMwRVJvCW5Q55UjTbFbP6mZOzKQ10x5hLHKMViFUPT2XUYlANQrFGyZKqD
Itxzy4l7tFLaeRd9Vjbrftz4JcaB8+2HdUsPzlbSzyTuZc0O1c1lt4ru8Gd1K3ZM
QSa0u5SrXp/YU+F/DUt+NF1Ku4AH09eeNZTZLrlZPRMNgTy9evKjBEk11ZjBHstl
7t09PrbPwJOvbdcFEiAq6zETcvlCiWuMu28Vx1LqAzbhrfg41+QHNc8cdxsz+BO5
6ADJXUNC4JOfFIt1H1l9gqrmq8pBygl8EJ//k5KkBevGeisiVNadQP8L0Q867hvw
xw63Ss3vn6Q6i97lBoeigS8kuTYKNvfTQrj6spr6/MXCIj0qPZCi2gWv6tCntqG6
/vM5XsMepXwGOJ4Zd/I5GLhLyxfz++DTd/cf2JbpbjBNO9Mog1DThVCZA0L9zc6k
EdcKPhvnKp1JIKxVicDb4Z46Frr3HiRjFXmmXxD6zGMcDpWMxZdroLJ7h2jBtbut
t/JArkvKw/9YjSOnT92h7k/dCiwVozBk+v4XdVrqVW330AITpvYOAZQX/troCRZh
Hp5O3wkU4PoCFfqTZLBXq9rJT9/uutUkEJUkTQMZePdYVRaQQd55GrMY+yahihMx
MsHeUTBEPj/sPhBqUUXS0zcO0tKqzOvRFmtdYlx1fj+tmOeYdRVPzKqc4Sdg9rer
mq+EJKhdWZbR1qzNcJOK7vZahC1AbPZCPm4oIPqQurEoLPHccq2fKTDUcx/v2SkL
Y6NxoOEOLjMLrcdIK6aJsO7/H1L9WPTt+FrSNw6eEMuxWhXceZz4Zji+Hb48nEPt
KhpsGc3X8c1pFL6yorlUg6TwEK7Sy8pGPh+ey/d3oPbLIGpQyPKS2y9bmxb+DgYz
zMQReercWVrTuEg92smVbSvF6iIQT8R/7eHTOCl+rn0RIRvo6obK6knPIdRpNqZU
y7NJbcD+KCyElB3Y7VrPrPZOkqLFV2wUkjKvTFlFTTMzz1SbDTNha/ClstGvnFDm
rKfMEldFAqzi88CHALw/IzdNN49Nc3QV0dgOqaneczfZXhnhIldkEjSJzVdkvLiE
XZS6uvb6O3GD4oFVtTaX6g4MTpKqF1sIOSJ5TPdSNyCouIbH7B1aplCi+KyuJ1qD
KluamE/SpotZQFxC5UxmZjc9MObeORrcVBi0AOSru2aQulls5ecvuKZ80BDopYz8
lvw5wPMdIP13nBWykiieGrEgz29hwZKTQBdi8opolMMOwee/Com2pmgobkQZyAhP
oEAQT4LS+4Cu6hHOjaLa5qkrmiGIbn3QkWurA+UiHTgx5lYxLTewTvnSiwErug26
O/Zv7J3PrYEhZDrmuEp0ZgaP6lmszK7eDkuo1yjlqSetlt0h/a+F6WW6Vfvdv/xJ
IwcYEg2D9cMr5h9zxlS+xuh+r0kMkExAP2R84ObH/WcBVTpEL37i/mj+CxW7/0+j
ovqvrZROi0V+NHvJyIUwWlMbRSlQbpC56KNo01wqO1AtuEwUM6zIEQ1/2LHhY4Mw
VnFDC7CyF0dmSH+06NVFiXdTCExt7zgb7xN5+3I57tI3v+4gHzV/oiHjfmJJ0Zho
rTRLA4z1T5cr8DP2AE8YcN5afwdDmp1iwu2ty0fpV79lzqhT4HxI5FnyNkAOv3lj
73upf8WKPs24gQTX/yUha/4/47vRq6pMQfNL/ljGy4ta2ItvqCKBsA0SY9LKsUQe
4KfFsDMa3SucutsuduKGxci/jqWctqI3aMum+Piih2XZwIiaOaYb5AKjDVZxip2P
sN0HUL4PzKXHjUmfD15Vw9XRv7fJC09IRwtVjQYvEndlFsYiIksx/uEAjdR8NQYG
7nT4oh/5nZuZG0xi6DFQf0IZ90pv+4aGAMjYLnr5bpZXPigAR0m53NLYpJNXTDlX
T529i7h4FueP3E4VwL5mv70hVJmJHV7mT6n/G+kNVjCWxh5Rg6jEYgaTfux/mdoR
kvAYXQCLO9vkQA/mfqLdiHfvRnjlcmNwjdoJ9djjjyl3nJJQeTjLgq/Cv6T2SLzu
RIJILWugEYk8tt4rpy2BtPaWjaBqQ55/CSR4u1EZENJUgYX3dMwjgEaMnGCC/D/z
vKlTwkJnQfDlEsdTdOM4ytbGpaHkitu3r6/KKT+aZdaWE+CZW18yQImrLQgDnpIf
gsIVcwcD1DXWc447yScVS8wwMDGYw6slJkVh53dWWPXE9VDArthzauOfwucDZGnH
+arX+AkzLh78MwN4e1fOuLvbXRS9M2V9gfvpVmdrLPZlvHVmg8vaRQ7GXYUW255V
IEBsbwZz4FvDGYqAKRyvt4TCx/cJMQkt7Tkv5JwQAOUdDvHP7/tS8s2ZFsXJNqKN
X5vTJeUA+5+uHYsIYLjwX8hXkdJqZsa9QxBBkfxW36JWhw34gkU3twGwD7wojLD0
9l9+vmN8si1c9jC7zsdryjzK9sAqq5yWIEd+0Y0UUfgcsFEcBHrSfB6KXXvPjyC4
KehqEJVawp2/Wg04pKZG9cozyqMg583kl+q6aF6USRQZDQC3WQZ2SktutBquErJY
8zS0llQxmwKQN8eZTnocQbod++AlUzZ6xL8lmKMkYLzG0efeLDheZTWqQ+b2hD8U
fKp06Ws5HEiwOEkSW6Zb05eZrpYgd2Q3D/uuHIt29grKE59izcGmrHQyUe3HPvWT
O5/Oi0q6odpkWJ284EyUkHeh8+YgVSUpd89qVc1GXaVnEi1BBvy1xI8J8QubuzH/
bSAILxkfJj1ZqdGbnGUs80xJnsCoF1FGsy2B4pLOkhDCNEljoUVGJvN0LYVKx+Va
D1snZfGXU09NAFuGtsE5Z6wHZ2gL/C0wPHu+sgvN4FffV9lmG1Psaa/z1Us2XRwv
oMsNmo7YQQuKbkbHeOEviT4nvIhkEvQcVWbom1tm4gHQxSbWauTsNHhC5DgEvoq8
n1dD7qQBUAkQB+dKtHfObnKAB/JWEquqgof5ib2D2F4pysLtn4qS/VexXtC0UuY8
nbmUoG4bFAfMYsEm8UTULYDsVFbFc+qxSExDxc5RyTtILt0uBnA4dY4gW/inftbd
j8JQUKyowoTWvrWstg9uzCzeEMDr11EXQ2fzzaaiUnJtfxYFYhBoxzk6jTNXKUfy
vCJrCgTThCjexK7mfCEB9gZySXtkhNj+16f5g5vgyzTx+hajIKEX2qGnjD6MysiS
8+YswlMNl9rP4HH7oBnNmqHMBUX3jrBK1rjxuH4lAObxmySVb81M7dn+6ICrbVZt
bJcBCh/92O1KrLC7MIxxj3RHl8uGSBh30K+ikBs4ToB9xqTCV6AfFqnJT3Lz9uRf
v40i8FJ1SSm72SjHOHui5k3UdSjMXXLglY6M2aTkWRTKTJdSm9zR9ewxQyJPJgk5
Dcwt1JqZwdsez/gaDat3bMHZ1gysBA34jImn7o0BqV+T1xK00tWDJ6uZoOIFXG4/
81PI0OXT4d8dhlxZFYEusDLeqDq3llpa8GL23Qqna4mOslzIhesuLYxy8L3i9CHd
pH2kg6zZ60qKwpAkw6yaoBQND0PKezYxkkjaVUkpbmxDFaPieDbNNAXemtcRfQwV
ZuCfzzhA2PfiX8F/cuNusEd7hSMFlQ47+0StBv+EyYAP4F4UyKMN/x+UT2MwjTVM
gQIBPGNpqsdTKY+jYjJyW8FmP35mfy5t1dnBufXASfUYUejBZ1iQJ00HQgIw1GYz
xDovL6e1bWRrv71kLlNFxS+wAYWQwug1r4mPzQhUO15m2ctjJ8dpxQZSsDXVpEKY
pckQ8U167a+ZLVJP/zv/JvSiOo0cDn4mzVW42wqjtydiI1lJ8ffxnANXmv3GqIRY
DF0DwD7z9QrL25AX5q5Xo/Hsu4aTZGg7C16Ij30RAs6nfwgzenvx4+EOiEM/ja+Y
/dmch5Fxvlcru4PIpdTPxBeHs+fLh4NQO/Ni7vhQpsMF2CSiI83SiXafmlmI7Ht4
dhHQfdtXW5H+VSVUizUqO0a8Z88BzWNonlZIrGcsUgGHRJhXDIvvyjb5R9vJne7y
Qbsde5KSsgF8QWu7rGb3L4aH2NQMTZGq+U6If+C0xzufReMk1pcFjipIUhqkzk3M
y8nOdSfiEv4VrK1qeJjpskDiEit89AfoPSuHb9kKWkzSFapE30wch2TC2gj/dDqQ
+vH70zMysK1WXogqS3MOoxpzd/55uUvnFBqUyHVbH+waEQolYHHpsnPvLwvuMDuq
QTss4+LJEXUVFe/nNR5uVn829MSUiMy21h7H0DKDrrd+9Sg6kQvfczxpXoaTQWth
XKlWcgrvI0ymwSg21Y1b/CQne4rfAOAa1o5nvFgNmYsNOThcRPXpFnb2FzLLAVvj
/CAQXmMg7DWjYmxH8E6C8yKXOIYsAB2AwVz1ILStiCsXBRBCNfIkNADQPtmRHMHd
/1/arpjWDaJEI0dkGY+ZLoQzb6RckkdZvBLnfb6Tqkx6jlm6tXo5MhsKEzbqNmY0
6PtCzR1vFMzcTZPcJf4Xqdwr9twQ5Ik2MzZOypqPzJ5aZw7r28bGRY5S3UYPXNKC
GKV2Atlxbd31zAEdfD3GuEN2zs7D+IXxoTvjSyB2kfNUnX8lWcGzvqaqC3L8rnYl
kTS/nWo7RgzRbvyflJMx2a8PkRYKnA4XgN/ZcQXHcK4RPjm4tgnhKqb38jrdBqTB
VcLTCD8UKCtRx06nsfo7GSr6zdCS9gmc/LOuuXDmpQaD1oQHvdy1njGaIg7gPxdT
8rSENkiGb+X+b/+3MgrAhsogQD0sbKDLeCMtM4YyNS6tNbTXZkbb7B/bQ52kImyx
rjNPQ+7l3vL4EbikT9PrbIyXg6LgU1MVsSVC2xg5k6tP98owjuwy4IwfkFZrmys/
uhqIU5YAbYjWANCiOVEFe6gscdeC7kPKnn9t3+lqbPfna2OhDc2vOaJGFETrbufs
bR+5Sdwx4TZxT+vn8bYq1T20plUHoLFajnMCvc1ylwtkvg7sw1zu/Gexvh+g/itu
3BRvOm+jT/S+zESgG4QzCCLWzWcTPwknnaTjIf+PIdkqSY7tz+IQAr2AYGtJbHqO
TcgHkTywhDnacNB1MGq5ApbMGt2wXahOzAQW7pdXVnmvdFz1lLsLXDk/Tp2kbxrP
cqUjJaLvpD39EKI8ApaLT7cR+DTMM2PUh8w21Iki4EH5eFrgUGGO7bB1wTxu8cR3
MH5Z/zttI0tzV1kOWplyrVzMmagrEUV7BQ02nSpCEPgCfCnsJFtM79G58jFGNMFU
4NYw7NMWGKONNBqljS3XnUnD0CrJVs36aIvO2AYFCifwX5gvJvmqTtBBb1NCKAcL
QDAmgBXFYci8HdogZV5pJmZ3Sv0wmKwxTlhmwxEP5/dohjO5MDWBvzn33vt+yF0m
4mAPZa5omt0Ep9UKpIklDZb/l9kp4V69iRgEVqog5gmlPLUgVAKDCz0NmiCB/Dzk
xOflLnIwj4rwH7PsAGXe0yvg6gmTC/mpyoktl2d7fYG9U3P8oThZwNg1DTc/ccqn
fWWKp/qy5r3HkFli4D7bxlgr2fXW0jVtFfiecElQ1SPuvUx/IQzW8Gx8h83xgcIe
oaJkZjVYVEBnbosonr7UkttF91VqDeQkC2unu0XDDHOB/M00R4HfUZJvNGOVc5xn
HyfIrTLufMKFUGQetERJfx/pfF49R5MvqlqXszpBsp9+4c3rYi2bPWD8o1R1ZeBu
W1Pt4bvt94AvDual9hyWGqLm3ebyjoR0RaFnXLJ/P66ojjYsnCgMwOSMXcBMfYk2
/UTpa/wQhysjQOu83M92NMJxcLigGBYdTKvvN2Yff+Sy6QQlL4fV4HCUKER8v7ld
TezsieLDSAQK4RkBH0Qycvs8xE3OOnvQbo2yUbNYrP953a64Z1xNFRqjeSTRSQaS
6ozZKZrnA3b2LuZwBcYewRzYpxT4n91lkFdKVcDgymkiE/Nmxcv+Duu/LCl3XJdH
weag3T8eR8gTsYpkBcqsQ2UK8td234kZxFdDeybHUECDXY/WjjX+seiJuJQ0V1+v
+9qWK3Mwf1ivLi/rI19YUEcw36z/WhHa6/O85hQvhbP1iqQPpCJVKOzkvJKO9FMe
tSkGGJGqj6f90hfe7jMexg01vNZpGGzfLoy1Q3j52Jsjci0lmdGe/XUZguLvBSbd
JLCgmYihlKvqFq84qjJ//i5N+SLQkqU+/8SW7woTf0JtGDEpFFM6CTsxmyO/T8SJ
uXHSwGbHODkLDtu23wj2TaM18wzrrBNo+prx59+XU5q0TQGCqf5B4Eff0cbMi6ah
XxunwpL0dBjJ8qhPk6SXJmOr3LiMFyeW3duGVK3H7teriKxQq1tQCqSnmNJtOPpr
/WQi67gOP5GWvlBUG4byvnldyoAWg/Q+erhYMS/4pttkf0JonO3B/voKGmF1Bj5y
JRtbJqTMyxCCCFpRdvSfwynKj9/lf6rIMuRa8g9nCjXiadi3/8kUw3CNkkF9gswW
bUHlnZEzIZyRTGdJYqjx8qPWx/DchbRsTS9MDp6kMdiBj2y/m6jGAEapWfvsj1Ac
eWWDxKodPqRgsg6EgReSAI6qJ92Lvyylc2TDoBF/CDbZ9AZvlrrUUyv1XCE5goBW
AguA9uLkrOOTnVwAwfPBwWHK6Mxa9LT6THICpWncpZa5EBrrAMw2E1XjR+MYMTqW
CihvNxuqkfXZ6/e7HQo4ZlqbXVmVCdbivGHFMC13rCee0oMocW5j9HN/oPRzyr9h
wlWxfJvjLX5yeN73rxNcMt+Qd2aPM7VrO/VJ6Wrzaak0YLPmxY9I2Nb0o9U7GEJr
ae8x6BOJYiiZ28XdscJqDHMJbL78yAgV7yEOHZQAOoOnl8l8V2Z4aigeOLtgRFvY
lUIsUJIYNDIw4MGN/yBNDrtKTlz6CwduC9eIV/0CQtmFPAolpiisPOC9Cb0BiXtp
yYJq5mw25NW93pbfMHoMP3oL3DATKeBWmefYNLBpINLJPd8mSLfo8/ZW8VrwcmbU
nAAmlmJnNIJtND0qQyaZS7+u5RGLwaAGUFZhgCkqW1Cy6ks4BpEoxjSGRhygR12N
eb4arokZQTK0Y0gbGgqlrOCQ9yMge1JPe7haDjgmKKW31Z1BJzOhKcSlFYpj9J6O
vu41XpyxXbZ4zeREx0iEUv3cI4+zWVm5oW/O22ReJqyz60GKnoGvTG8n/SLqRXi+
K75O3U2e315yaOQR71L4c0mRjdBk7UmkH0a5ldyk+aXCbWKhOGZUMMhB5Ex/vkCv
Gm18KV82CUNLzu56CZaWvkshm+AqDzq0gs9x+O0njJpQKFk03aZqJyRshzJe02aY
M0id6ep0iqP1zgv6NJQTvPbPIQmHyYgnbdz92m7wxE9sW087T4u2t8O03UaBd7p4
ZTMSAm/RXeB4DQus3n9jWtKxe3Y3YdEzD3WkTgSDMVc/wI1vGbRqjtGAe9g4CEHH
jy4O/768M1zSWS8dOCY8U6bHQXcKVrz9ZlUXvuVA62a5LRVdXlnSROmE7Xu81L92
s319zEq/wY0ZdeHmJ7s71uoCCWKwwlO9TLcdGXnYIQaU1muUIs+WZ0RAl4ukhkZk
708q4SkIvKfnOkYI/WC5/FZvmW1upqIiMSYTGTqSf1WrixL+7SZzL/XHa26nSvHY
5XAKTZqfDStyA9o/V5rmLoGuzcU8CvzYi8xoiC/QblXBCepaGLqQPEOis8RmP/N6
s+N7ydc4hVGxCn9W7MOqWS7ZBH2BHKOfMmqoA9V68O/3I/3CSQMlClpevINmrHr9
LR8WXiRCdVO4cv881oIGkEQ+sTMswRokEyt7e2w9Ix0QXzZP5oMix74vJVD+Bpzp
8SrZWmAOpD3G5dRyjMbaWdtj4JPVzf+tLjCcPEy2P1pTBRW/SDKJ9v/Apz5I1CKD
exbxewHXYQ9Fg8LP8CSkH5YZQmE/15DSfbrPNBLScEDR26uN85kuvZTkvqxnr7et
HjC9hT6hx2sQihPizO6/XdvF58h+g2yJ/Dt8miVzImUKCHIBSG5WK/2MI96cUQJb
AeU6pMdGdXjXk4kOEQAvKVbmtIMfvcOVUlkr1vMsYh5kQtunoOyFC+xraI+GJP7y
esc7/xp2jlDr1atgqPzmRbEJZm1KmpmbUyZA4nnNzY8zNsc7rlgDeAhbCQDK8ZpC
9Cw1CufW1Z/n5ZzSl5P/DMMH/4ymix4tpTKg8IdmGEVdigQts/IzeJFIvT9NccQo
iOhMAWQJhQiW00QiFI3pECORBD5pwrwmMclQ8snheO+YV0wvLDti1apXlAEMJJRA
vjEvzBtUm/ipVlRwABfy1pVK7PO8e5uC2iDHevudZnWPWIZBYw0iDfSd98rb39d6
o96E4q95V1s1kaNi7HPAJHYUBxJOIdN0I00zwadI2e1wZCgy2WzZ+f3m2J4XUTtb
1e1W+ITrst/qIcXPEEUfpOaCP1AyE9Qy+TfuP17Kj8Da8U3W2JFpN07lPUGbC/eo
q/YpT2uRNMkNGFykq1yFFFubjw4esqQzJ3JqdHjBTeicFEELYqrXNIEXfVHbBYNC
tSJ44tlealk8dfnjko8d2guXJO9bV+5FLwdqHeQefBVTo8tMOgBIcavrhJRZAtqi
ewzgtIO4USMmEL8ytz6kB4bH48Lw7OzfaFW/TjVcO4nhweVY5oUH4hn0G8AifTPU
uZglPRsNr7cq9WYn5/pgqhL+TNl78FTBylDRIXTFt2O5FfebrirZw3Q7+oO/R2Ur
xPaYHlNIAzM9FQHRG8pFVEtUahq1fWg2t60W8p6drCt8OG9joskgAYs5UquWkLIf
hPWpLvX1u5gRyv/RtaNiNrKiSDjPN6ywIDVRftiwr0sY0YcB74Kq7QOR1CvGw8e2
upy6e3r/jojvC0epojXNl4eDGE+Uz6/DPYtTiVnO4MFYT9DvP6LWa9+vq+rWOXOJ
Fkv/OuK489eYBxZ+MSpVw+xaCLrBvp1BOKBW8Wj3PESoAV3dTMyLNetDweGxxwJc
dJ9UJfLUBGRDQE4r4ojRmpGOTv7NtSXEqm3Z7Fu7uT3UKB0RtSc5RCD/G6528L3Q
bwuCvp8sQPW4qnQGic9O3p/VTu/kcvBcLUkeAi3ueVwiwWFZ2NCUS93l/rY8rabz
3az5RnfHsDULCOq6Gn8uvZC9Ava2Xpu31BIOqkpcCqk2o76aD9uz1MubS29YSuoH
QvwVTLPnzlrmiGoodEZkISghKR4Rzsg9r2ZWN0hgrbwRNao6i8Ym28Jw3eOHNK6N
31W5JujDq98MiiWfrNikFeDvd1yJCsJ1+4hfDoMg1nB2boBC+Lkx8sDpsrVlQx2+
pJZswsqM+4y06OQvlSyjFIzeHKkQarO6POIoeG8LlOKT/hqbl1HjJdBEXq3j2HP9
tY8ZX1iRLKn6Vf9+jCzSuF/nvp8uk0VdI9kRdHVL+MUvN6iCz6Osf7nLvsxYOZNu
44MmB5xYNLQfHGdai8LUa7jC6+OvEjWcwRZ8YKFgvq1+aq+MfvW7ackf5El/Wtid
VsaQL32BMCIr2cp961pL/u+j6ZPPK9NSjVhYx+JwyWt/OiCEmw2PjWf99XZjXtSP
R8GNwHYT6a08qtI7UfXRXV0DjomL2jF+xgTvvw+9YD3O2LIkEp8gU5v84UsjJmHH
pGEhQe6Rt6FEXIlEJ97bqH93N8lQM0s9YOwfk7pLWbulTse6dUASPMRVI+ZsWnHo
tf8O/hXB8MGGTa6RYgNqkVnKvXKYOKOrhcomnhWEWtneQde7oXX6S48WkIXKNUvU
Uuau5qna3F+/BBXnC4IBCyQ0zSXoUI7gQB6al7HDvaFyGOd2TlURPy3al2yvNMWf
e5dJBwPdUGFmZtNubRu0ygGZxHm9OBJkgmh0AauKKmRhF4EhD4974EtH24ELpFmS
zcwNJ+rf/hRH3row94XCDGeQbPuC3LSTdE7qk/xrauoLNJpbvjDBUS+5Ax3gYbES
luGdtNwzBl2We1Ml3ZTchQxHz8AObKXd0FXkSTn59xfbPdamFET2esROBfHnJOMv
RPGmstQ+zFrV30gjOybxFvWY1opKdUxrNcLnWchydKyJO5rRz/HRrePhnzm7RfCF
G1Fqyq26rmAZ+Li+RKL/S9JXZt2pg3mvCHFpgPMaUGofvf9L98zdfDYFMLbb5GTu
jIUoGvG7RWFGQgQGH9UaXugCzjlY00zemuaKTxSMhMUffR8+BdY/5GpDseHLPffm
vuNQ192MgQ0mIixjz9J6mcuoOBKwekt7s2rKN2kgtqfYxsCxUnw0difY6y5Fd+t6
l9KBtB092mxXMCioct/FtsVvH5EPpGT4Mh2ktoLM75GVazriyiTFjrt4wESZqUA6
JLqOGh5kTzxoKOE76GzHbZlVVEYWLYh6s49++0VqJ9J6jzFB67la57mGd6kf90Hh
VzXoNlE/bVZWtvH9Gm3hrNWIH652BL7AxDKkmLob498Ig8Xg5Ln0WhT8qMM6UVu7
SpOibC66wd6nTi6SjVxCBivUYNhWBsEx3WWcigpcRe3BGzjdKnECccP2E5bLUx9U
110nbfCEUnAoyMUjQOzw7BPazxzPYfNHHLk+3CJ9kgDxJRcjJH7t1zJb0sn5ihPb
V8B5HkHpKH8Hhkra95tgAhzuvOBhxprJV7HJvtV8wxJ4gXdx0eTtziTdnpVPULvR
ddrzwPZhDTqTukmIBotyIzPMDqbhloMVlZw0Nj7qIhVJpYquMQoV4690WZ087iol
PYxuImqVOmXgo4BpmMG8OvOxEtkNd81+60C/y+V6o58gNFYpt0VvrL92Mea9x+Bv
CncT8BPTytAF7e3vvjlz2klQAsuiMtbimBtgKI2NPw+GQT++V7CqRmOuGm7yP+ub
QNOzof/x0PSj1I/cHbxt6LbEgKv616rCa3k8AueKlRo69nKhgUxHK1GweoEzrUKp
wfksrfzPkMZBCvrCg6PTXOR2K4THGZxUS+Xq4DQQyVlsOkoJd4FZtz70ednnFcay
7XwC3D1AX9WY6Yd0d+j/mjB9SUiJANTIpEKOaqu8OnLmD7Nry1pGfqmA2dVMoMWz
pOIodOLFV/v4AtoauggKWODenb8W74lPsVvnJL1dVpXjyZC4sl/YPgZ3IfjeRzTR
ntzbCxtfaZ1/xLShVKqbQg3cBKl79rkuoQhNwFdC1ocFvWuzJk2GlzFiiw1K5Kfl
qvf0PpNVptxmSzbEa0zLqtT9bwzCQRr0AbQBQGQRkRUL6LH7UBRnD4mkT8rN76XG
aqhazIWdI6hNdxNi6Hn/d0+lcS3T/Y6MsBOXuscqxQnKBtCAehnuosh1ZwccMDBP
CsSmd86YCHQQoB4no5bs/rx5/J+a5xGLfzjt5r2CUhfRaupX07JypOTEg+tYK9K8
FLtVyWYlX9qZm6hWDnGWc2mhlTbCttr9ZnHN9C1+QIw66zlqWv1RzLvOG7f7d6EE
qGbj4QkAl+FcclBxMlURkMC0C+xJFzK2ZhhmFMpMDmSyUcmD5yc6/zk/SV2GjQQP
1c5ZxOphFpQAc0iA+ECnuQ4DxQhGirBkGDtcyyOjNnaNdpfCo0wvXED8pCqBaHQz
/Clh1Y0pjQZDrLP/rGnzsGpqqHPxATpu2zieUs278ygX5FKLyGLqH+LjZ9MTfN7R
2GrFAXWZ6SSfboFR0Gpv2ZWIGN8BIrPSC/ePKZmeqXeQVS1cgjRcL8XH5YZSDuu/
ir/q9dMh80hf60uysDBkpPlDPpXln4ip5Ov5tohcAiafSSavKJDEfwnyt288Opol
CaiUFDfLY1lEmeM+gLLryl80rve4BQO8cSA4b/W0wqmgNZJ9C62tVzfrN0Yg3vjy
q/fsnxMa5yzK6a+PGhkh/8UFsf64iRMzzMMyCHE98tYlAr5t0qEtI/mgEFjGgaDM
ywqfdrqQ0aT5ayhav7oah648t+shgmEwTNTqlTEpkZToszE/qqv+IP9NlTXhpFnT
L2UqI2B9+RH5fgA0uhhYhGSLmYL7WkkRuMNTKQuAmoC33kTwkZVP5JdOTAZ3+vF/
wImLE+B4wSoIFzPD4a0CmOhyNbNE7AJ6JegyjoSrdjVxBVd2dxVUC27UXvRUnZFY
8XzkVrfI0LFLMGa1erICZQ1H6fxRv6ObNIZhI5y9Nc7DbicXLjgBO+nTypv4bU7e
2Eu6rqqZRa8DDDNiDGhhiWBeVbwtQRQV36XLir6HHkmRc6ddArZ7rnE2xYRRQTlC
zgG40jb27J+jozSGNfasOSkV1Ng3iZxsPgh6IfZhOHOQXNp1Q+LWtIYT9J4Iz5in
8XJJjIX6+WOGDzVbm5MddMMbaKT6x1UKMyzADa4BUpO880MzJt6SMLFt71l5cm9O
Npgg1p9yG4MdOUyST5CO7O7GTPP2VkQWvdsFbPttW9hZ9BlwIitnEqdtM33M2B+9
ixNtLV1r+YKzsmjVglvzrefes+JdqZxX85f92r5fcPxrTW4hVZQH6GJppt4piHZE
nQPbRMmP8UJZMbmt+WzbCBR/M75dquSMUv7W9PYjCNX5sAZ2zMoz/sSAeKUHj8VV
bUhFScvc/dfu2tR0m3R94x/eaFDrak/BKTWMK6i7AmctnzBnYTgeW0DfODXjdS0p
uNhB0eBFG4ne+rioxkwY2n72mK+kZaKT1d7nINSwEIl+MTbhuLQXi5qODP91IR4O
yC5bPqrEu02XsI2InBSKoQv04idfKR+Oelq3fiIRvGHtv+iebxs7gdaEnccUg+Bn
v0wWu2AgwAREhkYEXPzOfPCk/VBQbFTki74ToJ0q4MooY0tvFAUhnZsRJPF17mWT
vrQ2CpdkboK+5DupA+FOpNTjNIxKN1IPX6V+xwmxJHJQZByCMUDHFyyoPU3v61zB
3d/bFMZ0M8wxebOin10L8IHVvLPRkuIFT5V8aZipMGDrjdwwhDmZtzb6vj0lwL/P
70UDpBXVfr3P40LLLbxHB3RCKkkweRdp19leZMzNnNDXoI4AWBzspse80hdInu+O
s6n0XipxcilO8ngmvn9DVmaJCY7gW+iDK5RzU71vtOFvTQsaiab2hSVN1AL3lnlF
bva8HnGm96hnmM295P013ZDCp1x9p2wXN/yX0Icu6ONbR8F2/dxsFdrFayFM7yvu
uQ66xNkQ9IsJ8NjmjSzCsoVdKrvyp86YSuV08IGrw72H2xu2/vZanXICMTzK6qmo
6l+UgUjXs8FoKBixAzogWFWc1Jl3SeQExryypvOxuB9jk0beHGZQMYb2DjuBDWZe
M3kWKo7lpWT4Y7lZAiKSvDWePm+iGlTIhNJDzLMG4QET9lvwn7H726m99nDrh3iH
wNKz4aCrLHh02RBCOXPygZW0udE702MmZjpQt4HaD3TAKp831wzKTMdq9DOhtcP4
5QOJWIroppPo0Ri/i2pgl2RLx3WooFIxSlkhFYAP/0UhE2RNhqIQ72fi+ARgKstS
ZcJIVcwkZJIRzJXXh00L7MwEWmtMMHjt346ZZ4jNgDpRrLa1mltyfMa+aszcPMim
zqJqNdUy1OEV6uG0G+s2nULrJnzAAziYbZ8cHcg8m//ACnJpDImaD3njrcPe3ohK
VG2XtdE1gLbAuFqRVpZ4J6NSeH1q5OBzjOhS0Ej1JdHkqxP12Rj5gbBo+/LbnQmo
kGIBIW/5pTPAiCPPwvLRnxi7lGkuXXckk7uNBXip+sjXwNvgJo5VmBMJGnOI0j1F
bIKRUGcOfHecrv/kVTOqSROwMjqK3N0fARfStZcUvE/gddscqwxbFvI/prDbXAZR
88ZOSRdSik/4tY7JQxPnIIMbJOlBMkASaJoCVGxiz9wrt0Y9mkkoh6E2OXw79ZiU
tNnmCediiUo+jCH/Mof72oYCortV0s/hNuejzfR9IEvWd7d3v+xkhs1k4NdNfbyO
9/LOwj2okpikV6W7Z00rw1+eBWl0MAqCCLL2jkbbcGFOjczs8ycyHbIN4hL1RjxM
SQcEq2meE54za/r4oQHAaNhhk+AcTGjfmPBvkVhZiK6eys4TG2nMFQdHuiWlCEh4
kOrmvcrHt2dar7wCY9MvXOP0FBe6o+hHT6PSSyLwDCZwcteGKXFOcc4ukIdVhK0G
Vvs9GCQoByIQhvVc0nmgD6b2FRTO7p2figIJp56Y/NEDheCfes9yXAyrGKTOz3cR
x6DZOCvKq1nKeAJW6bQKI/8otVhoeNs2vZSeQEvuHSE6GFpTuHenIWhrjz8B+aC6
NOxHWk2igLaAXQmZzh3gotMB8bLfLlLs6scGdqiVjmvMRWadVLh4sqRBFn5ZZ5+K
bHw71d6Ou4EqA6F47GzvuP0FlxwUhMKZeVJddVqnzXlVImMPPm/TjxN2plf/QhCN
vCqKsG8yuVVSseitlKtzShZu4DipGz1yg4+MZxyMvOHAoGvBRPWlV30TLQFGBjup
fUlq5Yb+IwaraYWgXxH+CA2DS70We8+xoCsZ9mmhXc3p32uJokLmKhlGfgsVxa9C
D1OAuUv7uPD8DMeUP0p0n8jNDQ4bneoVQtRumRHIrK6KG8mHI+uLwqqTOi6iaiuQ
yMACWCQN8ra/T/U64SJi5JxvMmpALyXBhe48DXBiI4sWLmCCktiORdoOf7uYJ1eb
PggoWg7Kp3TybinMgde2kUUQlYLFH0wLShPoH3cVkD9efIN1LSVLWqEsFBHSEIgK
UUrBipV18ukpHqk6ul7YgqhKkmAo/PxMpUPsYU9zNekEmunr+5o9vPSKa24cdWfS
h40KiNgy07hBrZrUeO3w8rpe+/nM662RdsCe6BbKDjD4UOeIKCi+gIQy8VECWlbc
QmqjHcfZ1QJg1ZOxxNSfekbH7QuXbYPjdvd+KohVKFZwDyRzm7miXgirt/N4Qq+m
6/94qwW1yBeJ4WOAgqzSc9DmQhUxhgzlelt3/spyaGbMPjze7UUHc/GbB8WVRdgc
5u7Chlur01pUJfnItKukdmOMIH4gL9YQKu1NeRzsLE2ffnAYWqDbQT3AYG1xWBjY
gmPHXyrdgasmWELTwzRw2gvxFXVzy47TjQAuQAzvLtZnzFd/2n6wujzyWhmbMe7A
bK8b6QbZWrMC/4tPIpHJoUDHeaRUqdVqpfnLuSRqTXovzrPwcKvXm5+IYoT+Rdw/
j6Gye4bCbZR6QnHPPnzTPveakD0jf4LpUDyzInQYDBgx1+4RiT3n2kjz/CfcQf8g
6mGMMlCekKIQjrIi3nkBfbCmt5M6kwvG22oA+8S2BVXiC4gBRfE4clvyE7lBsS6I
yCDovN0vmazcOdGkHZ8m2q3GjT0gzTNqrSb0yrcY5B4BVkkViq2gqlg9W8PBXZnE
PeP8ZWY9pkkywzMgWngi/PpzM9IEDFNpfUzB76sccAMy+d1oBjqjO/XCOOwVa8KL
4wifpwmEqyFRrFQqkCO/7FeiMKFUdPNffm+THGyo0F2ibeM3+wdlovLgwqME1+OH
aSXstmZrvXLpqTZQcJvksqnK8V70UUV42hoUjHV7BLuFohJxPFQAjG8X2ygo1wqn
emDgeEVh4Plkn4Sw+fG9rfaE0yRevJK5vOZf516PYgUcS9bUpU+gV8uRGD/U6M+Z
t3mGcb3zTVhk9qSIgpzfPmP1lYYDavo8yI8Pve31dn2MiPxOZVQY5sFDS98OwF3r
W1qlSUlDkMkmzE3qLfe+Dl/UW1kQhKk8lNQyQInTAep2gB5XLnBLNkptez4LUa6r
PSZk/BrwUijyiYo9Rvnou5bG+d7FT6HVIGu0A1zMpmJHrYFTLGb/Kne8nsmB0a6v
fDpOlOtklMiRpJv8dY5Yn/zk42VQ0ZaiCRfhunPPjUCYTFWo0CtjOjfGw6Rrm5gq
3vdIGo5NsvTiD+Y5KZJE4r/IVuLlgHYWtWyRkb1vJfemWFyUaBcByzZmuLkWfCIJ
tvKDf+s4YWSAmkJf6GgDjr8CmV1RTyZzp6vo/bk7cnzPRE9aG8RjynZe9zvvXV9g
9DFPkG7auDecSG0ltRI/YiWwczqnsgfTpWgoh8gtKQb8W+ZfniNYHKu9deQEJFlU
CgEcJpn+OI5IpAuA/Bu7U/OEaVL/xf9xsNVxa9CKuapswxsQ8ZOSo86Gwb6VPKdS
yF5D9uICC0d69mxazUfu/IisJqVFAmTTNAG8x+z+aQ/E4k7+1Klm6Uq+Bxz3uphG
p+7N09uAiSwCuV9PgCS8TMC6GtC9VWbDPctRTVMIk5sYxu569BqhzFiGIn/QdmyS
c33YPLQS46snMf3fv0pHZHUkwaL/rMSC58WBP1eRMuJDTEsrF0CM2xcdcHzxQAYw
q/jd1AxDwqPThVSenXUbcMWavaqOGGYP5OoV/LTywGGt7udKz5wnkdHXwM0o+R3b
29tNHh87weeOAz2Tj3g4ZARg/ja7AHX5PkxRAL2qz2D631ZvJCSk8pHH9KnK0/yr
yqg1GjhSHci1bV/wh05w+PbG3xIFtUqrSSRbFwRjRvCTgnfNP4vlg/HikAIsX1z8
+SYjyAmULuw2+7xHzQvkzkx9dTlftlHKlJY166TPv7byZw9kEI2L8gDY3o1hvk/X
KvoB5u+IYabKDr1a3AiSJ4K0I4h0KnrgnqlxsDOAT94gkYixzP+u89a0Q/fDJUiN
Y2YI14MnMW2KQaL2J9jJJjoMsTU0UfVDmeQXifKCs6hWxrbzZ9BMnk4JqMVea5Hq
7NBQ4Z01zxcQItnRDxMSuspg2TJWMJcVXM4SyBzd+jH3o8TVHJgTZKiW+SheRgYS
4ai3w+RwUnlg8JCjI9F2r4967T3+4poGe0BY1RKNPtHbl8/mwE3nVwUS+AR3FK1v
3oeXPw+HwL1w429eSDLiXPn+29hB4+mbDNGXL0qz6Bn5v/n4FXAO68s2ETqQDghB
YGRdWfG7Ka+mpRMPQ0/PMz+KkNsRjsvkkvsDflvgEybk7YqT7x4dZlp1W3e/ypnM
+dBLIy68Lpvka+eZ5T5VISSqtPrwitGDCSuArYZ0+DMD8QhqtlvCtibvEVunrKhT
mLnkUhdYYDa/YYzVcJgsgtW0hhkbe5NjABBHCLVz4Abrp8ycHkJhbOVE352z33QR
UyKRD2uhVSauQ43FcOSxLLtiDDUHE+a2h2F4pKyYidKcQxm82qgqD5yvJoS+BiDi
+NprbKCpuQI7uHK6AoV/8ZzJChwtvrVIYxik8JyELYNk+C0yMt1iPf1idtGoXtEx
bOLNlE0oin3TtdUbNCF4uDcGpOF+5RICD8R53HK6AxucRmo3+NHPuF8wrQkrKM/d
lxHcPrcH/N0Nsug+Eu2ABZGDCAZAp/ilhGvJc1Ki3MHUmsuU0pqvcLENVYJRql6U
ybg7ptQ9nakfR4hdHg9gfnv2CJdMEc8aBpozDxATJlrfQ7KMFbcDX2s0NBmR8pwz
dbQyVtn0Mj1jMvpZA80or8ChfvXH/gTeKHjFl1y6BIHhJhiaRj/rzsCpQgLjJX5+
0eXWa7yfgJ+6ADIslPn6Y7WlfvGg4KdWRzy+VUocLOPfbhs/EdyEFWX5qGSwy3r5
PNYSz3I2LTbf/VsDtNBkHQXGLzTVrSVn218P6WL3UzBZlP3LGvAJPhFo9p2WOXLA
+G/mNX1DuNQ/h1b8vPUDoGaxjxdA65NTDIUvhZHK7AVgwDzBycwtpZTCdd5C7z3y
jIYwYxHGuT0KCI6ZuhcwBCtVhUyAEi2zgH6SgCR176AdFVwZl+VXZYmnIbQnQGYi
cKe6SpEcqJN4KKHW1mSZ86IFbbTQEt59XrmBgY+Fmompv+AqImnO6mbYZS62haOM
3w9ClB3usGxJiDTEfFZVbHicyI5BOJ6ILBsns2g9/sCMeeekeZzylYDfbeeobxCG
Y+skv+SwdTpP/PV2hBlryHMu2wPqhAGiLIC7lzfSVIsEFyQIa38uXDAHJV+QPXc/
Mq40MndQ9Ymo6x/KxYdGuQNjIZl8YJAQ4IxoCdlzbLH0MfusJqT7OAFGjNgdXjnV
J975dSLd8CI7HrGUx8uICj5MxhMfOuTNbKGUZb+SnM0pVerYOZDfwyt40OsRDwFE
7iMxKEDNsdeXqpC1IuA52KQvOxfJvH4+7vlJH3x84PWEMUx2FAH1huImf+BYbRwq
gR8KgTgr/opp3vADEgBHejxIEZc9a7kGvbUZMuB5FAF+lJz44FeC+Zxj1lBSSUBA
KG6cK4a30SEVrlyClf8MpSo46ewe8yKgeVxymqtJ6pYuS1+dUrydslF8NGNWBsnn
MnlS01PJFqjZmAjPIGIy7bIOwpx3jU9v1h0T7svluVYOHNzGBZYTX1KXiHBRCXns
6bNKiqnHh+OURGcRvYgQUMOjoAe4VdXGHp5URyeBpVokVxCbIqU3SDIQIbgJu5LS
BLZ26SSbmVghnX3kSKJ8KXrNMAxZvfMv4ALbHc6/kk1FZJs1rJ4lGpyv0vbnvQv3
YAb1JltgnM538rJnGLDPnjsCv95GYt5sDCTJ42nYIr5aFsA90Au7XwrjZoU30sph
BVyOK3UAZPHW/D0TFrnWJqvfTxWx9Mned0BJ5UmQcvmEuZwt7rPJqO0y60gFs7lB
1ZTcxrAa9P2M46IwdyxT7Gih+/aLzpUvLvL+zmXf+FgHlT+qdHLrRWCKE5nEo37W
MuoWPKD/pn9Go6wzlLaL4T65C7lqh4Ma6HHDaOehlnU9TN1SaCExrradBLAaXHRj
QDRhr/1lyVrYRd8/blFQlEtKFtdNFUHbjxuJBoFsFH9SIbPLvEEhHjZzwYjdbp7+
+7Hu+Jj88iNSYhwhHpunJZKTKyEZEuCFMV//r1uOV3PNwLK5dp/jSHLZmFQY5BaX
rG/fCGPl3NFZ2ON5rLM+DmfunL1UPmhHkL37Bw5swAjk6CLcIXKbdNbFt28gDd5a
bEFuDXsaA5CvFb21AE9FXv7N5tNiTaTqv1sNPmCOmbtJUlA8iiTP1r2InFh52OID
HeAm3p0QXDoNGzZsjzWDHcmjzuAyLfd/fJkdKIuGh6pi5WLwp0Muj6D0Vg9WyFtS
RcHfos5+7IN7ylQghPmP3Wl6uPEZe3p9Lt8muMLZJoSPYBtsfq9feKYNnvhBiNRz
Sd6IPHWOAFJwdwHKsump//3LJDNyPQuDKugfSsW4LbDUiRK66tPr9oFvSUGLW28C
Cdv8lUXFcr9L1doqIE0fqae0+/CPJkfU7LgzVDZzUX2lLtZWz88KGPKE8xg2/Rxh
j3S5fuSNIdAJohUArNY9aYTga8GWQGNzBiz6Vf1O+Zz+Z+Faq5btLzVYoDBtbgKV
bECxFoygG1/9C42kMDugXob4XZdxZR22gfpDVPETsZEYsWNjJBBgMO0Vw0GisiEP
//JQBRUPIcFlm1B3TRqFkKO0RYPnshuMZ8jTRjtip0z5witwUFnPruUhbr9pq0oz
lFj4xYuCxVfuWtC1XJKjzqQ89OWE8m6CwOdzFi0iRDHl3saLYP0SQJpU3EfEZdEs
gNhcshgOYkiQgofupyskpA5aWDMqc+nSBAO15OUM0F1ay287TN+vaJ3jUDgNytm6
2d+yRnilQkUbZslUU5b8AkCg5Ft/ZW/j/UgiJtygig08nSz0Xw9y9EFm+eUx7dwe
gbM37cRTMFJlN8aIJuu1qRs8Xy5SW6H7Wko7iM1BsnfEiYEoN36FixeEiSlleJAO
GZsGkOs4Ooks/1JpR3XuldtJ5JJQLJR7XXpTTBQsowvgOBQ5RZpepyH0USh0JgwO
VJByLyuwfm+zdEXJtfFSNu6IzQMFVXle1nhzCHASF9eFi4lkR6Ka+dYPAuHmtCeA
vy8JNqhrtcWxeQxaDU5gnJ3aodLVJGTUrhkvGIO+rwC6rCZsC37eURHs/Oprj/7X
XI0azJdoKVekpIeONaGdaMGU3ahWxtEC/R0iUi2ib36INZcTi3y7Y5KbZqGv0ART
wGyNadh2Lj+m6718lL67zXu2FNRJ281+Y9/l7PCWYfDZWbhXm767tkr6tfv001rw
R8VkUlypxjPV9aRsvxGpg0IoXr4XjExLSD+pyw74+Qd8gj8em68XDYoqIIJ4aQaF
ywm/DX95+HtZaLAHszwoLfblksdt2YPdf/AStnmi8ATLsUfYw8emk1iLcld1pcL3
KMDqJtk4RHSJIGhn8qG3cPweny1Vc2gXeshpgKsb4jA06+SXsGM8+nqsOezNHJW1
/we23qtCFM5Rgopt3Q5TQSULqEVDz8X6e/1ed90cIadGkNVKMIY18WtWMg5gjyXY
T4bCN8ndUbMAfb9NKO+DwM+Hj04shRmv7fd9b6AknrpEDqBNLbAvi7KHhRkfTDEU
CboUv6sfdjkJ8nFqI5e7wZxQu+86MLIQ6QIp2egAfJKISyHAzaZnTINhZGpLxSvA
u4ytDTmeIp5uYrLQkGRSk8jJwHnP2+Km1hWyOQCK/tardSqxI8gySSwAGE11NNnH
spz2FpUvvH0mTMqgCOnJwhDxPvq+ieHflYxUyJaPhvarCLDG0R9xCSjR9F9Aa8C3
xauSshv9eX8KGZY6LOJkpADXT3fAaN3afHwu6WYntujDRVo6vN1KIgvrJwa7vAyE
Sht7iNqJn2NH34Qw6v8GYfiVOgIGECtVA7iTD3ym2t+1L/wRwg9d6UTt5qRUozGP
/q+oXpU62GBAGC0UbgXCH87RzGzTWR10fd8/xDODnDkYgu6pWvCNBAoee0D7Xgf/
Q8HfBk9R/sVwC7KGJeaXcn1scryvCvzMnecsOtWYczVvkBHgBvmKJxDQoLOsCf8q
RJaRGxPVmSWMgjrGPb81pir8tLBb09puWenNCPuwqmyQJe/cJYa9xbEHmHAuiQiY
bW1nIf7+2IfZiXy8IwkftFLcl9aJdcxx2LjZnEOxEzZoRTRFZWcqZri9wUNzMzSZ
HL4mrEFsEqPol7xMkshT6yB3kUjYzm9WOaJyalLf0TsfpriC/uY+ZOq2po5xXSR+
UMMKyv5sGYJCYwrSEGuCGbQW4Um7T0kJZ3w9YvwXmGag8N0i/fc5PHy53t/V2C+5
1oHKr1fh1xWCMOf+DA3HycgNwkXkUkYXh1XjT/sjikSj+q9RE9KXW75JFzKNj528
9XlgBVqwxtl6w2MTE1Z+hH4LHSp+kRdd0X1lRHamJO04tnaU6Kp4RFlQ83aqbUb4
ce0wVUCSdloSNcpSZNLVUWmCyZfwUu9VgXIluzFUN2W7r6B5dtxy0cD6tGEGvGFq
7ax4Ap/rhUtORdTHjHxizM7MvjiDGAw/D5u2gfZESK51fMI40g86Uc/esF8PawxS
4M6RDiJIKGUd9uMVCEDIVKbu5LJ85gIO0tLwNMDJbKEyNHKSOSCpV6U5uHa5sa8/
2DCFwIQ36Xn0sgbTjQj5j/RoPiIatWogkbDk8Nyh/G4Rq8Fp+gvw+tZny5Gbi8MP
qm9U3BlGMPKf+9CpX91wnYgk7Sl0ccBchDpGZasCRJjDdQD1uNajCxOa2krMusLi
2GIOn1tn5oZ8AYUp/vZBUJhbg7ZPJASEbjXI4nt2onkFw3JMqYhq54dGsla8OsW9
fXhpv7QDw+uIcu8vvTrNwuTTohWYyDEfexk3h9C8lry6fxx4OCqnSqdLQ62Pmwza
ErP6vJ7VehCB5Z6aeLK9wHD5Z/B/0P4SOTEWcMfR4ixa9FqIxoCf9Dkay7XE4qZu
0STWNdu/QP4H8S8Qz0Kj4PxW7DeWN0enpxTT9wYv4C1HJaNjc7T8kdGgB70sLjVJ
xHx43btOiqp9fvDB1iVH/eBhxCOgLg9q9sICB//b/mSik7HNkWr88aqNViH/vYCb
Fyfp+whubS80ULJ/VKwWASz+OVxPZj4wP3E/CwDFG2e2j3IbuaENHH59XopUtG3M
Nk22+x6+F7+HXtdCz8EIIPeHW3sBpplJ+DV+uklO+h3b+firpo/pApfKIpAMa2tF
2Q+y00a+HSL+Sn9T+AQF0/XiotSSgjT3CMlqDlgH8+pWT5PFVkQZY/ZA+iXUIxCk
FfCP856OOLqc0OQW1nzAWeOnytY7OgyP2cAhs9ZqlfJ61MUHweW+cNWfwUSgMAuc
J3Vs9i04lk1/6OAD+nt4yqCU8z8ZbOB05/6s/XiwAoKsUORb1DwDNvNj330OSyEW
10395jPf9UlIpriduKGF0zBsk2u45eh5O1kOgh2cnBbGhWJF1qUpib7ze2Hr6aBW
gPDH9O23Hhe41v5rYZrscpYW4H55gnN/GEzngNr/9HcmEckB3945JoB15ao8UIjk
JUC6HFchMPszYAk6bjfh/5bPLxjfaHSIBLVpapFX63IhWihn6+FK4AK4DC0Zqgwg
B1GYTG7o4243dLJ4pstqYFzkI0ZVAUZm2rgeVSnSISO0i0JzHa99NwWH6l9xvlAd
FQ0aOd4VZcdjJ4ImMIWfBidWLIJ+SYO5MdDc/pLmRHKDTaQ0Tkn266NPytBfgWx8
wnsByBOA1qPBI6OHI6sMoZtf2gizU49YtqHhLt3nGb0puJBgUgcZ7vf6VICbu8Ut
Vs6KCoQqKcLFP7rE+CTwyP+j7WW9xjerknplkHVuf+ac5sUEi3E4XhjkZ8gw5rMG
ww9I2hgJmggiiGKNyibNJvuoIZ7Q+3xEbvfC9gVQh2b+pJAucOJFoP80XUqWILDH
kOJOkVNYA33zjC6DS9ock3jseW23svprpdVkbVqG7UnLFSfGi7g6S7HCBboWnXvQ
9E2CkmSrRGno5Wx6ymFz/9UerVH97CSMX0qUKHKu2ewdjonEKBAUz8FUKLUpwC8f
9HfdWGax8Dw99txuLmzHV1mUVRq2qCaPvEISFTIWrbI1ZFACFUNTBJngLIvia0er
U3xbws3VB37sVvhqW5y/TvMvRldRm+YO37nUsfbDyNZqB1YrfM6TxuV+jzhgNzn+
aZM8DJ3nDbhloroabyvnP8EQox2vOzMDNixmKb5O8+rgB7EOl99IOYXW+I2JczQT
dRINXB3gjTLTSV0mbUc9VHWhJFkDQsFQ7wcLZ5x0IUsx6pKX3ny0xtL8HAhSVD8D
gLkjDKI7Rmf6DJdJr7s8fEq9Zb8SWRNqLVoUKQxrjuJRaTBB3tFNBxK7WvKKDqWs
DhGLEMkHLqCv4CmxTa1FaRzV05nbdqGQbJ/F3po5cLOqYg4PRHhbL91wAKPNjypV
TDbrghj96EhHKhf/1qUuABmFh27/gDY4oDlAtregBLhMiMBeG8ldj0PhUvQxYyKk
j8Mx5HGH6CFbnMYbjCKVa4JJ+VG0nbcYV2JLgGHBZdouTt/Hzz2clZaHhb/CYJkM
K3GIe8sxsPmbEAVlKnK7REWVMLHbUwC67PA0918Mk8vDsds/bCZxsF+CkpOlI6bN
5b46zNh7z1bqA33bsloiLjby8UaQqFzGoag2mL042xIrdBGu3YWaFCzoJdm+qLGa
8CCivROoOEq7OS1sIprQrocBMXmLhcdvHLpiy9Q4Kh/IwsQxDuVg1oUatwhR7AEE
bvW4fkjm3fchnuJ9fa1pzoEavU5gG/WWA2BbbXXWskCAzfB+KiCKiNGt+tipRc5g
X+uTeQYAbP0yyQD0BoIoepsJGgPBhLrDTWSLODUyqvKZO444BWta6EIF52gwEtCC
gdEUjTKAUq88jkZPbqM4/dI/7hVJnQsiT08785D5j5D45K9vaIpS6B7+Lis0nUMe
vxmb458WcISNMIAh/g6cTxM5hY8hgIzisSCs8BMTVhcXzProfTYrltiF9Eyo9E/2
izxIIYZejl4Io32ZmlNOeYvsKXs5Cmu0rVp7Uk9TElDj4ni15Db7qtlRpVGZzIoN
hdo7VUG7xphNLS1+34gTuYpfqvZ30KfhEvgqcRdVbOad+gxlvAO7CNiWQso+1V1W
/+Cwp3fGf+89+KCIyQxRLxPgRyILEpKseDKULBVtUTNgAepyLND/BnfJYjSR0u0w
tnILmugChB1ZwDxKS2PnhW7jUIeywEsLt51njygnE9NeWJdDeH/71aJUxH7gEvlB
Dyx+2XHbqpUMYIHX0YdYEKsJ8cHl+XD3XJ/evv8LgcAAx3cMVofD55qmEdJMmyx4
rjqd6jbs581ZutX/6uFAxce5Vvke0PJNmtKcqJcvZct5NYK+xm+XoLmfPDjTzDsl
8v43V8gfYKfq1w53O+VqX0Et1YUfi3C+5dEDUn1GLEWdAk4PuHeypJFEdCu4ucpw
KqNjPC7Vv7g4hrEDfe94ovAbV06sSp3vd8Ufl+oAXhveqVYbbwqz/1PHzEC0ZEjt
UCcYJ7ocqfhswTNAnA5EKLjw1brTUc3Ov1X9hGEoihCuR5wJqA9wgWTdwMp9mAbi
XhkJIUkl/HqGZKgWoLepvJ0Uk2S+dkt1hSpTEBSqPuD6bS7avHwbzWeBoq9vWV4u
45+4o9eXC1OQz0M6+RuZHvdLl2Jfm+Ulv9RlvTSGnbWV0Z5QPnuTRKGXzeP22VY1
XE3GLpiUQROX+8mdUi/22snnrD7dWdK5sLmMOrHlkY5jZwegMJIvl9Y2nEWT1MLh
qEHjnd7HSQTNvbb36NF8Fo50DWt1Y/6pvSdpSDIB3AEBFXITxA+6xjO3RGKeBnLX
Z2Z9dBjyUKEDUydvPVsTMIvSPREbOo0EPgDXgllEBP9NkpzL9ptGiTWRGyrDcA0u
7KLkqw5g/2IbRlfw7MUg8FtgfgkZLF0s6SuNxe3etajakLAApa/4o6xvmdKKkSfb
6JzYm7cavsmuv3XPJ+cMXgVzSiz+g5s+IrEha4Q7kZlYaU9qwzTmXPQcYvtV2T++
A1/LzpUH4kOnarFfxYqgGXQ52/L2ewRXfMhVZ+HBD4lt1uyQVR5733DsYzwJFd8J
LY1ukXJgDC4uaS/bnJcT/tpF2eZ2guzrNLsTrAkFSc8UK9b5VbVdCiO1JF+EEuUM
SdegNswYWCuPyNWNvloicLEgVr3DjLS+td1YA36ORsAd8hcc2b56mqJddzEnGmBD
a83woTeisUPJymsB1g9kNigT1s4GouspjraZhnGbaymRCZvZ2SgTvFKiUkOH13ev
TptZ7/Kk2aGxu8nHUgXJeEWa9hxcDvb86eCSAi2UqwaKt7VlsaxGaFEoRsq7hP1X
69z8DN21xnNgV4KV+RCvzaDI4OydBq3onEdv3g8+o8er7Nw8qEwDq+MTAntBxpqk
m+yd0sdR/DhbT+ai1KHJRr71bV+UhhInMLf2IIQp6cY/DmvM868jf1sViqyO9QuQ
REj9x2bJgikLlsRvO7DfjIEL36REmTSQMfLj27Id6SKcg+aCZVe9z7VKChl6VSjN
jchOel13aZMTn1Rd+BAcZXxWtgtnqg68RjThDxrGVhDRV623ZCUg4c2xtesdbmZf
wwcmSIuAt8uGyd9yzo/nsGMrFLP8jAoB8FqfhjTwafNu/J/Ui7NmRC4Fr7K95Ycp
VCeBNr7lOdPzwNM9Ub6oITT5hDTuZX3lLy/lB36d61qtfl6eQlLByUJzdkKkGgS0
ghtkdeNYyaaSO1d4zA2U8CZISf74I8LIs1CHMDOaiiZEU+ZqdoxZhBZffuGkT+hC
5mz6wcABPkRZdiOanTMFPNCy55rI02uLzPwl4+YnD38I2uQeZZQ9SIn8+C41tlGo
ZfZ7NFlrTV7bQ3EA0BAebKwnpSwBYOeaNpFBf/OWwKTnwEY2bXBEJ5NaJt7PLBca
f3wjZVZaUqhCdjhJf+H8/iOSPUgZt1oJnSwWBYcK3QdAWSqgIvZW0Rma6ammmvOX
HzLt7ZGU85I2WA1b1pTWJxWj4nS470dLM8Y7+0HV6HkhdwLnLyU8PREUuC2XwjCa
t3hq02SuuBHhZWOZGmWACvrmkJju1CfbY+ZP6cQMvKLjdZMifZ/vgn84ChhvxtDz
oBpovzu5Zj5D6LT4nEjX6EdkDHmi/qVbwKE0K470ccsPkG0FCD418h+quRwb72i8
UL3QE3oXdBV444cgLFbennjinKCsC+HSRKZxMKUbKj+j9ameib0Kp1vrVDACDamy
Glsz+G7I05hZXhT510+npuR+e4kqgJcnfADDsAvEkMqIdNqMns5jrvZYFBS67Eio
mu8uSAb2zBwkz8QvuPY6aBOhCFCSSGng3XTSMiBXeb9ZalA2uHomyaTJVMNELgPW
xj16KBPcrEYz7rebIyhtH595BZHiQgLRY1BuXFk4W5gNPddoFmeQysPoOI+VCZfQ
J8Ij/xOH2sWv7hVL8FwgW62uqc1hu21DADmvBvln+GVQJZyyL5ecpZMh7iXX6MK8
VO2Tehyih5PbEmrGOIYX/wL1k0dcBO8gFTFWShJxd18zO8VPFGWqdLcV+fhtzbd7
cUDUhrKW5Kg0RC3eVSpM4+UwrBWzLE/IMbDZ9Mf9oUkgF+qCNSKZ4cwb0WNLqUkQ
2UfFDu9wrcGUTtQSmtZjdkrfY0iwNQ8EIuANsdlhKyRXCdG+Z3Ws532yvnIbtFJr
3YT2S7NjfV1DM6CqcU3MdWokr5QBG7IT4i2/SMDisfStHz1RvBExkxQhirCMPAjf
w3Tdo88ueiZ2kC2rP8tw6U12dt7eSS+tN5D1pacOu7GFSUmD+tQE7Y/7y9TSh+4X
b0q7pKjBQnYCtq3p4tqQPKwjN/2Z1jwAHYZCOkJSxg1LIwub2P0dp8EWdzb7q02q
CtcZerTkino8CaXZcNlFaTN+ZSp93IeBY14M5d3dA/fiM8fn80TYLDXjt+uPMVZl
yA2E6ShkhevdUQaVo3GYdKHMH813Oe/r2GqPJlRWEhsZHd4HHED6hmGn7yeU1Yvp
048eUxwCqCUuSHYNwJcQ5qgpGw48OKmkNvZ+1ToSBmXQ/mqVTbvwguuR4sExdVCP
buDVoT+mAWRreCqM8ZbAl9RdSiUIdVp+qDlXgxnEhi60p/L3DOF6LJg8G/Uxms86
BHNJseLXUzmzbwJx2XXWgPo31baPyO/kkCc1wOsw+Dp/z9yu99mhb4SBkLrBnDQ+
CWA0IYdfhtiB7xTWU6TmA/x0AKOQQDDbfrNNzVfTtqGVMxOmfdQgjXD5tNCbofLI
BFHrb2iVb2F6TpnH2FYxKLHSn74gEUV4Z026jwUHxzpjlRtHu5k1J3BO3ZOv9YY3
v12Ns7tnX8uzqKqhEXrXTc3whMkDY0hGwjsAbgFBrCaZZu6YMWP78PySOA5Z90Xb
9EzsXPCcMtlGoI633zSUZZJUjV2Qe1lhW422tBojkT6Rd6TJ2O/Fzdn5ds582H3z
7F/M7Joqcz/5FCXxTIsrOlpPypkhZDxPIIhvNt+vCm8i8yOZCntXkCCWFB1Of6RI
ujq/EoMpJdpUUpePVjPdGtvmuJQATzwYkIqVA++vaEH3pBjBnZUX7OdKB8cuu8/r
mQzbfPTnrLkcEecwjmDoOEKV3Yq0wPmQlcOyQBZ4ggeWTDEUaHG8/4M0jomAu7kY
2fv0mvL3gtxDREg8MeUABd620+yIfPnYi+S+iL1cUhKJ4MtZAEmxlrU+C9jPOa6e
Q+D7pRsoG8TCciySGr6IghCOt5vqSD0izlKtJVmm63z0Hnqx2Y7AEn0SWNsK/ia1
nj4BW0NUzOZBdCMKjqdVd1Ek9H9hGs1x27oQ7iV2UIApLV3p6A7++mbQgM7V+fGL
azFmEmIdfCRMDJ0zlVm5gETWMQT0f1PiRPvabJ2PtgMuJs7TJQmZ4pQW8qst+7zU
CSNhOnRKptTXrwNXvlHvVAxQ3h5uqI5z5eBeIf/xJjA/M/vaXiS/plsSlu+yzSSa
FG/LuiyBuhD4Kb7fMCrpo6VF6hn3IocL50+Ag1FEs0aUj09tKtSiuaNFlTPJBcfU
b4qGOg74Y+Rz4N1JIWgGPYpm444EBwQr1EdcweAZXqYLMYaN4vlQ4KagH6S9i1/W
zs/XjyYLYR0Iy5HiBLLmvXvs0aPFJV2Dc7mPuyC3Ot15jl+/XeI392z7ROpomVmy
qppVs7UfzDdyoOKctddp8xtp0PQkYC+GHef1VvoxHrXgFViH2mLPRF2sXAh6+5AC
Mn/fJsskCUduDhoerqfWJHVFXuNZ46jIhiwus/HNkXhui1OWy4ZZr19rGq2FMJkX
pGWdt1sJL20MPke1npQdzrjLmM+IOpNihkgDXBGdXusqj6KdwD3+hDfVYStWoeff
NmZ8NRNnvDJyfgODgcYQh3b+zygbOukpsBBST9PkMlqDQuCpRCdm+jmtYNgSwyW+
JhdNjq6rpXfbIlrojzgv7L/2VOjnq0jZLV4tSXS/lfgvexMIhxpWF8J7yBAJXSIM
T0LG5pVRsIwEr+t0Ppv+fDvjL8N6dBH6Xv+HKSwOzm8kyH+c1+ekxMpCQQPGiA7E
s5Zzp0Fph7s0+60+R75bM4rU5ygSrWfEkHZKotEVVG9TXn5FHSsLa41lMrxuygrP
phR51PeRoZXH8C+Nbp1UhdFys/k54vb1Ur8+yNdXQ2r7iHwZoJn0pVwXLx+rwj45
rB/wu276m79kmOjUzc7tVh/Cj4whEfJVEJ6d4ePpQQrymPe+hONuwRFYn4IBYT3r
MfjjHcqIaw3XnnStvrAtLRtI7QtyaDfENOpFZrJtUOJx+vsaG9IFrPTcyj/zvE15
8McuOn5eO8Q4YM0P0iD9sIyMR/MKd9dhQrCcjRZxzFiPDCFWhGhXGNrnwc1LrEQw
99UhV2LWhIYkyku6UT78wrOKDD5VZHIoHdpgkjko4szbC9iofw/h79DvFMj6CFkh
tiehjGdadqkBk2/9W9v/qFK6kkTGkHHtjmuyrAHFqNdkqP7WutWLSGmpFJ864nla
DyKwsYVFbV/LE3FGSmPzrgzT29SoxDvAJT8urVQ1YcOwUJ0MSAR3lOLEI5RiX13m
MoXudmblC0Ec7fFWLSRzOI3pnUwxB5/WZKv2pL/KnEIyg/7EUhRn9d3ORNcXpOjn
cHZreXR+W/fE3QHCaPcSeg/0DVbQnFAOwglPe9hiFKLbHn0slWe9kAJGzyZl5Gt9
e1fC71gP/9nFgg26gnEYC7ZBXC7QvwhdPhAcOGZhLibeQnbvHDPRac+cu5pS7x9p
yOgTigTXSfuwbs78PlvJ82gBpdXk9tEIi2eOhm9gr/rUu1lWUm/el8JGhiEImgdu
8MsvCdQQh054kowhh+Sj6up87Hd8qydAQIZevoExiaKqw8gBEi4r0cThuPJVdSO9
/T/5fEdnpSd0bNMyGRPKONkidc+YKhNUzJYhRdYI+xYGwm1SN499nS27jpNTniRy
pkRHtSelMoV2xrNK2udPMP+NwhyBxJ33jhLkZmcJEc4mOtxXSzw2WfvKfj40+ZzU
Lz1WgB4eQOWkXJKOvj+NGuEPPUCLqfHtipq4GGEqw8AvwsC/1wBoQgMaQhqNysU/
69dfRGCMpkmFB15I7s+8Y5xCb69qLKIqERp+8psnrEOvJfadYipSEgdCrpEluEmB
+yjyKeO8p/eBvYMu9FX8IG/4qJhF2ZzVMg47ESGh2onCnJtIY4QZYCDMjscCusfe
QkxS3zaVzyWW+Ks/5IA4k+S0nzribzSx4es1vn/BUqCq8utEugY3cWJCI1ngipfZ
4xnesjpPQrumAtAiR5CP6GCnucJOCjCVVxwk3nZzSos4MP/5TNqlVlm00kQ/Ak+J
BCSlmPTkK3g3DOP89Q/ItE/MeMoftUVB4zFZyVlpEXlqHDsMNJemOfmkVhKLgHda
MiuVWfEMmfkrrKsCN7wi3T5Y1AdNhKiLSOkAdQ+Ij+ViRcrUL6SxIC0+sjVthXxw
q+RH/0MIzaY5k6Lk/bQQDSGT+j4kibEOvQ5kvoP+MCDiZyRj34JbsGt8RZjiHJqe
i+xFhxvWe7LCp7nF9Q7KgXWVdUkH6G+8xtCdSvHX/DDD+V5utOV9/nuv4TZ4PnuP
YmDI3GpoxPIMTqF6UVQ2YPAEN3Y+qj36fTJzu8REISBbSJXwjUm8ID0AvFspNxSJ
RfldGuK4j72l9eJdnPSGgA5W3AlfRaon36TsnySW/wlHygEOwxVs1aDtivP6qybm
MoBDm9SIIz1RbAJMmZoJTtbBBDfIR006WB3X2Q6TxgfwyAtxy13HP5n4HWWkc2RK
xXVuyN814SGcN3zpF6S08V+no+PUurXccpLEv1pjlHIbx2Skml8ttByLycEZHETJ
HUSoZwxnGT9Sj7f+SavNaK9RY8pc0Sd01gg63SxXdVF01Z5bSenJBMBiTpVvjQNc
CCzdI/Ebf6LVFd9184MRbRmFaLjfIvwg07FNliuB1gSfDzP2vbSj9JuOW647C9hC
OUFw4A1e775+3kzcjnrlBJU5KCzk3A4QIGtNBVnm2RVTf/mhaejUyM5KzIaljwun
hrYjA2gREygdyOd6S/bbb+hAGOdixigy2vDnMPXVgjJvMF5naUae6dlAj9wZjgDP
wPnQt4+l+f9KayETkgfIpUuQvsBFuUQb7TLtg4e7FjzKX0L0AABJ8d/4fkJsZglm
YVv8ZIVEzCDrzhsQR/EQ7546jJYFIG70TzE/8TbGu0IuVDdYYrmlEBVuthbNUAXy
Chr8YOqqydJak/Rs/tjrydzoBJWS1OLjEPt55BqB5wb1VPZuWe0fJsCeCGeD12vQ
dQ8FavQi5VoT1s51h+JsgzBxgteFyuJ2g3/8rRkNWhAm8ckufKjdjtFaQG6PIN2g
+Gj4aW6J2zN4QWNrJsHLnte9wwsnVi0rXkObxGni4+gFA3zHgBN16aziuE+0ttS+
Fx8Pr0UA7xJlnSGNUa5RsT6xC/4CDJLR8X2dwRlguUxZ+DKlejAf+PfQ4TlDme4R
VXYHBkM0n8l6PtFFtFyBQFVE5H6/mRshJ89gtnGlwyo6952K8v4lJOoRzxT4T8by
yDBvKBleRKVdvyLtRkl10j1ibyEC09k+/YWRe6U2aHrSMqPROFdTGBu+N6DvpH3y
Mc9VOrqxUbkJ35Dssk3ZbF4KvTpeb5DtwKDdAN698Ly5188S2xz6Ow6ib2rGtEdl
QkDiqe7OTM4Jwf04bkQOflsBnbDq7nC2VehygaLmgyR7nTfkn587MllzuIbaiZTj
iZD5nl7SPUgg4qYJSJBsmkA9Qm0PtJuCKKuzHKemW7fqW2LtpljeO2hXLT6rRgJD
m3SK4G1yXXbzzd41RtFCKCNXeeuDs8MbcDHfPutr7En6qj/AvWeOD1kd4IZ7/DBe
bOolLLQ/cc37wsrMnzCADEodbOWMY2y3TJiWunPff7Apg5htXbHxMF/6aAXZFM0z
lMpdfwHIXNrSRNSQZIWEywvEPdy4DDqtaoHLRxnqN4SS+bDYRWXH6qRwaeIF7b6w
wCd5MU5guZaAyEkGEqv63kR4r42wykfV/EEKxWPSoqzlunkPEY2X7S7AaEo15ivu
cvh+IXyDR876LYfahODNCRZ7x8NbMfBOEmvJI4y/4VyuwsUVYkC3s6+df4Xo2bNg
tOlFgHD6PcBNVtK2PvXegcI5A7ZfQVisAzY9OmsD3mO/GjIphMLyKrQxi+TaygDi
b1sP0iwx+FHWiUjPbpU97yrGbOW+iBqDh94lrMZ90y8n33GPeyLhLnDyisxcrbe+
2/4XZp8Er7jkLfxDAYQL0Pvt8zjbnl2pu4YGnC1Wswoqm1LezJ1InzcqUhh1V85Q
nM128rDYDrdDNquc8QfrcdMtqhbU3Iqg8DvdS/bdKII3m40MJd1P9UiqYz61gYQg
2UwHvVYJlXjY7peSnnXpMS3QVIgmMKxZdhdcH0qwRobJGXcopyP/08Ae98dpHdax
2rLZ0K6/u+fIE1S84EaHkukYiQsxkhWBGTK8Cc6meVSYW5EcyYXimC4wLLQgShX6
ldFufb950Mtp+ZInhZJqf27yM8AeHiWS2YU8Cdwm4+Nb/6cO6HJlMoCmiOdK2Euz
EHgbvjRRGk3zJ0qieE7ZI1Nb0GCC4urny0bCEq4oaH0l/wgCWFgs9+TQN+MuiEpa
cfxDZgOt11skeq2RrTSv61icaaifxtzu5R9EBmifJjSIOo+Eu4IHQoNAkCIrqduS
llbJqpIZodyGCLsF+1lFYp96IaQZse0v39SUrJCE/v/d+kLnTzsYVYbLPsfH79zp
7XmDhwBPRG3kxscOmRVo3R9g+73GSVV4m+coKQKvLBPFvt35T66BVqPgsbvpXT4w
W8qu66kopzqm2P/hvH18mCIpnBwqito6PN7mkm400REQ752xOy5Y5e68pxW0/6b2
nN2TCB7TC6Wn4RYoWoA+HT2oT2pklUjKXi/cQZ7sqdIhCRxBt/md11GmGTIK1it1
+dUF4UgnP5cG+JxqSUYYfnyw7MVK7x1/fT5zDDCJzfk+m4u54PLZ8pgbguvsF81/
3sJ3i/cjkxax5OFD2/qcsJngOwoggiI9Ny53QvEOkVMQHWjN5xOn7dO9kMgnKS5e
BJuQAIrNhV9ly+3qESprTZQK8FxGCivUXWS/nbaefsUgNoxbq0dFfXjXm6i5ZlKW
iNBdd5IaaaI5d2FzWBobVZ4telXQlahBEfhpUuAxv3P0ZpBb95nG8WP18MBKJaJr
G9Ty/OpPl3LyjlXXqCbvoi+m/0qyEBJVFPMINmUquhfZ565Lf6nLT7aRnKuuMj3T
uc5zGCMhtGCZTEAXWZ9etFC6NOraQQI+YqJvKk+e1v22qL9klt9cb1G1ZjenutE/
IXuhwpFKGhFYcDasYJVXDM+n02wHw5y5cUsasTcfIX3NNPk2/HUj/HnGho3h9kst
XMWo4uwqIB8x9B/1u+pAFjLS+DyDNns8aRUdCetTvuQ8G7SPI2BFedDB9VO7Ly0w
lJ0lYJTfUeZAUeSzfqdUa68cyYTb6W7BXu6coAH+50MYA83l7nBorWGlQM83yNvi
qglQqcTO02TB0vS0RMK7IIGUceGEybw/pAEUiOmU0/dM2wU/pdYvL7FoXZYFbk/V
NRgLiBUlgHlHLns4sj58rsBUQf+HACWLHGM2aKpZSmNR42YGbvEQ4fhm53DhmoHy
VWv+oDDF7HtbNPBeC4/bXX1qMsLdtPH/LC2zQ7jggAFIJIa7rf0AREsOp3PD7AT/
gFyKg2V7ySAczhS0/V5HIbKxpVhnTbweJQsFYGRS9MF752jR3YiuaEUNZ6Ymdy6R
/aFoxMHexwr8MxSGmj95mNXSOtGh8Q1/5G5beG3N3cFnaReddvmc0O33GQbUPtCR
uPSVn87oUQYfGikHyOOmtGSxOd4JBOK2eUxAi7ahcYk7D66oGWzH3RCVYaTaTCY1
v233tnl/OjK0DUkXhYwoiE4nGfFyDe+hbmNY/2PHlYujuE8X4Z8TRxn/OBmVVy59
H9JsPbx2ncHIDTjM75Qqdb1XAZ8345NS0GNH7UAwnPOONVZXD+JO3ZSqYTnq32Bf
31huJtrEnDe8m99QAZ9QLja++/iL1EDwfkJS+EpeZVbTt8+7+5+SFBB1KKv9WM/I
gwLKhi8gviTHdVYbXq5hnseXaQ8LPh+W2elaYPxYVP5HHTOjqUEPOBQL/C5hQTUi
L5XU491Cc0R2Q2X3OQm7z/fd59dr4zbRJby8s+thb3KM98ShshC97NkJYT6Kxe1e
rCfSmSq6NJZV6lCv1XsHLS5/H+4aEKvIF9mGTKfinSPxbsQfz0KRZ2UMTcYfjaaG
4izTxmu88544dvi+XFsjmd2bC5t1rlRtD7ceG1vNSNERffsG+yN5rwKCQ2vndWt6
jqCjxK6BWmFqzz3jT9/X6rIvrGUtBTdpUXVXp6UAphoo+/wTdJ74EujBFs0Hx2iw
9xORcQVbxb76wewsXa0iZbZB9typ+ucScTtcr/jsLD+NHT8O5Oqyo6LhUHf3HfA7
QhhGXGagciMBJi8qanHY3JW8yoVkc5lm1/rhpLA4a/kVTrOJq6BQb9M7Ao7bpvs7
j+8yc5M7LzGXf7SL7+kWcv1EiKSud0F6KcDfZ39V5GuFJlNWC8MD04i+S5X+zc9F
vsQVH3GUeAw/fPZ8qMJ8EopyXqNb7l79qaZmzENaocheP4tjYfpFxY8mZWlV1kia
WYbphxVkDhLQkL2juHtczGy2laXGzMsvjJxpdVaMo+xMlEq/DDRbdRMay/4Zkasg
QfRFhmkGn8PTv5zSA2Mnl2GtwTzTKBgTTig9Ynd339FTvSPs7aeTp/oaTD+wYOZV
d/INlo31NMsPfOs/tAgsVLtf+HoV5ru9l8LZvFghblyoA04hYyIQsU+4XTVIpQuD
bkM7zm2wks855sTdji9oUaYgjnkx64G2ZpIvKceE4j8YMyJoMLnZzVLoX4ziv7xJ
wBZWK+633Ad4ZPnsrd4aKIqnRVeCsDT3ySzPza81WC1igrmCnqmG787n4FWcbvC+
iodEK5ibJfpPKi3OOWq7stav4ZwPpbjZma3JdipmDPO2pveooZ3nB05iTuaqTPI2
GW1bix0DY6COSF4MoMhTmL6hbFaNYu0jw53atyK3Ih92GYujiy9nQ8diLnV5OPXS
neFGTYtoKgesNkmmAZLktUN7SyBdbzfyjd+cTXCCw+Vleu3/TTwndrPjvg2s7ZSE
YF3CZk/r/svRph5/w+Dqsjc9nu98PFG1Rv+Kq1rb+S6Q6Ek1YeUiZRq3v4RR2VHq
MHQxDBhPnmQMA19y9qAk/tOsCFCibcZDSfk58AkbO+rNDaK57iR+yfuSaEjP1Cah
h8ZSBDQAywPZ18mu/MjOy7XTuDWlktJ+e3V1YlLPSRJhax4o3OzFv0VIayI586Vt
DaZe+2f9c2DThXqbe9S97Xc1bKOnlXGUvlUiqXsbeD+vtT88xu790RXK5/8YXyfy
ZllRObmpxLPj6My03N2WyaJlYBMRtJ+5sUNXg74DDkIjQ/k8oJ98C5UO5oICFmg4
vMR6bgE32y7YAeFitlIQnQsk42zcXHOlPMGin8RwoUGF6kHymyjfSbVOyoqiZbHD
/PhDxQHTfqFwzLT/EQmWDCVQJBvx9EIOThQ0c5tu0/Yts/2OMWj8Ob3Nl9EPCazP
7uyf+Ff7I0/fmPMumPH91hwRpTzzUL+Qiy9NLuoLwihm8wUlu8NUFcmVP0JltXGH
qK44DUzHIBaW4gBFTpVkpehnixQYqmsli3f3Qg/vb+USWnASdkgwhefYM72xG+YI
4uNxg2tarXfxObIlGvjdkrVvULqQeY6iDtMFunrI8gHCKfR9kUAHtAkfzCz9pdVq
9UOZhjezU5pk49ZawEX9qIu7gZsf2vKDa/aDbaho4FNw/lCRPVxCmx0WenblsmQo
klp3Tm5STJS2Lnwgy1B+AJQgwPHZPtZPKbbXeRk5Wsxwx+0mEkHllG/Z9luh3P6L
DQ+Ja2j1/FYeZeUrn1p094ckLJ9geLj06sIm2tO33xESqv9PmoiC+14AJhJLtgBa
UNEcnKVakXhaljlb+Oukl/HiFI53jNKwHU7fK3KPo0q6LCwGoOxK/pdxeA3jqpO1
teY5UtZQTh3trjHvnhEjywM6+EFsHx8+exiYj2phJdPLluqr+oVje0lvqLDOX/np
dbP6fUnAy/8asbRKmOjxYu9fItGeKIwAgO65ScO1P9Yr123eeMoQcmdPh1a8tRai
V5DAvkQD1Vxx3zHYtrJCQjMhm1LB2NwtsA4QmZxPcOxo40s0O0IsozqrnuTN2dat
6xO6OXakR5RoFptlKJ3f9Ns842DExImB1McsUvfEArSiV8PJnvDP9hS0yUpTahmZ
8BVwyXA4JXF6ZUz8RogGIVcppiku7FUluktzN0U/4GnceZti+37QA6gkPt31EuAE
NZL3Miz8bZ6xC93x63WHpuNz9Om7J3d2QcHoNvp5L0bvcb3vMchdmhH9Laqv44hR
TKJNZ8ZYMm95gJkYiT1t95uDqboCYzceDheOwlcuHmTZk7W4ED4U0FBKUMyL9Ypj
5/+UqkSLOFEMKJ3xzS5WIN98EjfZaSbUxeI+F1ST1T4jLW4veP9A0edyXFni5ljG
JFpcKGhm3ba00H2sdtw98/6Pe+KUfU7PvGRGH9RZGQZSOkLqYn25Zy9+2StZvCxI
ngW9bfes2yjGpZUcqgu/BI9wqnWpcFkxBS2/ONIn6X9mqD+rsbyKwIpEfHuOalDF
0JXm+tiPmSuJIbEkuezcyvK8GyOSfXJD00rbeaGHprhNBp2Fffx+bIStP0Q+D0xs
Y7iPyFSZsak9QD3HVhy+CPCfWn/g6Hb6v9XybZZT1gdtxzldcVnJarZDEU6CrGVs
sVnb5DSzAI/DDYafDTuzHdJwz18ouOIoyKkkmGseGC+/yH4RwAOkek9UuxdxUU34
SSqxIMWcjmSEZ6N6G8AEwdKQmHmeD4fj9EaSbEC3zKd3fJrGmCVAmMXqKeOH1lZH
hxhhb+tzD5OvRWF5dotPrXj9tE+u+gSGRnnGxtUxb0f9fBF379FU5vqT+6YuqRkh
jCWYMiSvy4h66Fhz7Q3tWaLi4vHk6/Z8G8n+AOQ4t85Ei/Mg2vgPi/Rk52mAKq94
T8rRvORorBszhwclWhtUY3gtDPo85FgR7jOUqMLcEufR9Ql5zU5oD6bpS7mgVr4B
1NjRgJg6hwR6oQMXbQVGzXAgsN4HLqpAgkN0yy/CdCwblm6MZUiNRXu36reMfwmT
7itpHCS0qG2yFE3uPojAM43rC/mFf4xGRptMb5VlL1effSr6z+N9XW5DFmsgE1P/
PAdI5H09h94/qxgdv7KhQUT0yef66MswtRV5n+WZNE3AkMOUpG/Ft1Se3flOXQB/
TvEhbq8yojH+J05nuZGaMVi8nDLw0I5onxi79TlFNiCHMJTEBjBShHUWpBZw1ves
lHCMy1rinN0qJL7OpnlTjUyu67j3ycWmuH0oqZmdhx9VgNHiDQFYcRE0QuVo53y2
1P19ZUiIuh/3qP9b80bjjavsIxNQOnGYZLHmTg/x4tFTacPXLg1vxl1PlKu6QB/J
LRTvYVkI502RzOVAZFrZ+WqWiEZYrrVwnmkAplpo9yjyZ76J5q5VLao6oR6j7+/o
uXR4U1M7fOMLR+Tlw828iZ73qIeaLEpqErO1l+9jUy13h1kmWqAjuKeG5DkgOufq
v2xnHkY7ubCQUiTe6CrB+KAxY1JCqN2FiyTncZdq4X2FMElpKcR8DL5YF4NgxUXh
ZGdX1mqn6WQzcs1oEe2nJ9FPDlitEUlqLHPdHXmPvbZa/2MTGdSzsgCoK93T82vL
8pTsRmbABoqxmZSzQrlluTzoAnDv4gISVqjo40u/IDXOCiZVTM66UUjY0PJBTxst
/eKxa9zI99KxTpDMridt6zNCDwpo+sw2cDvHGdVV8jXh7xOKc+HOlNHn6+KAivWi
R9Ub5DEe/rfIg9siVvTOb02X3ermTuhKe3lgUY0KURXZsbFVowkskc3EomvM4xP5
66wi12HmK6kocd6I9ghXlzBEbnR4Asws+vl0t/CI6KIXxd7A+MBIo6/CGPbttsCY
7JyooWD23/6iI4VORN6tFOJMxeko490Kzf15CBmyI+INhnCMTCZtFCapqJ5VZfTO
9tHMx6hHnKeq2XIUdcIIRzMXMKEyuXcjLoVMbW69dzPVoTWoF3ADRhpA7Lw80IVu
Tc6id/5CkuR2Nb0n09S3So8arU2dfcKhOPPk+RA17IMG9QPVGfDbiJxiIddmn/ws
a4Cl04mFsEjuhL/RBuYvcOUABLh67nxSQiVUDOWX/6sXdMD7Eb3uOcXE3284/jW2
5CsVXlEoI7MAKOU6wjYQRCpN4l2ImisU99NCegNNm4Cf7k2oHZLNLHePJwPe+tIA
Cv4XOyusYBG5nNVdhaJa5uM4uOcAjU5XcJ/F6J0g2Z55g4mBcrO4pN2EUj0Jo5Ra
3d7SaHzF54oGjmSJB30oJEykolODWcoepy/kx1sO4nLoRwZISsa3LYrT06SHLH8w
kN58jAJBItTR1K88nkRXmuQ45mN2yrGqm2zx+BTL57cscmD0jJ2KlSBGR8Cr+i7a
Wx+knj1T5YSoIJSOr6yGCn4pt5wyjWHK3fh8FjS2GGmU2reZz42zawYCmVDxXu35
FXCJY1VrS8kv479lRrGmDmVy8k9CrYZtKSA7dEZ1ORe4kwuLTOgM7nmSwC9KOw14
XaiVvyOQXB5N+a7EX9Qn/A1qxeYy6axP/bPaI+QAlENaSysKGijs+hHKDSjqgsoA
2rCQhT6kdmqkbWteTp8JMuft1ejoZ6Ng7RXfH3exmyIQReGAouiEc3K2ZoBFmEic
PHAOMoXp9PFiewFnPZu0lO4UAlKuboHZLbAmPcW4hiHpFNVSO9zSeqXR1vl7deJC
mK3qNqpU8bWLqXqO/qQNyug/Sv/urnpNrWqfUQ+Znke9RD/IfwJT32PFfkNx472Z
/ToZ03V+j2v4YASRguhz+CUzlpgRZ86wbDqkgt4sjKKE6RvJxRMgUY+bkOHOed6u
hv11HM9safoPI70/AFOl3hWciu3Ufvv1J9hr4HawmRP4kRs5GS39xIdbRC2GmDm6
YbBehWQeFYqxMtPBEf+r8HVvokgkOHobPcOkS0Pxc9uZTf8tIBf/eml+mN8veQj4
0jquLcvax75bJ4rrLYYwJ3qgpRRwUgJp78eu8kNzEWo9oIHoqjVhSxLEEbgZMmIr
3hEVXHXfwD3OMtiHhgGjCIlQm9ijLgmwBDdHh1t72i119Bn+lDrHdzV0+w4F/5hD
JuM0eOLyzOOwwk2IKDM4sTI8dsYSi7rXpLR1/cg9LHtsYd3AcJO1jCu83Ufbharo
DiCMlpl+/3ZFVejEQlnipbhVdym3PNuSWNKK5+q61auEovXStDNRugUm/77JGWUB
q9Tk2EKOoMZwIgh2PJPfCLp3k4+hGEeuabMw4pZ7zdZDj12jDFGRm0xVMXQDCwZb
UJGFJl8qvCTwcWZYsmBEI5HMDHrbCTiCQgmEKS3vnxHv267VyPsODhcwvheDo0ZR
ir4eVRM8HEwgGuOuq6jHqutj6qr7q9O+0Hi5XxHoeVm8E+ujrJJKfRl/EMYiDpX3
bW0RFSIZBwSlO/6/WENTQaqmg3SolUOhpheliJdEwjZS4FosrPtNLWEx0ynFWY+4
U+WOC21kWSg0DkQnqrA+j628J9ZITid8DCECy8OnI6C8eZKk4KRY95yriJzngT9g
eIaU8LSLCCl3lQWZkSHpvxOMV+HytqnkqwcNR8X+LwjLVoEM1Jsmp4D9+no+Rxpm
o5Nl6yubjc5OkhfUl0xtxTu/6gg3N0rSFRnCfGUH/6dBehn1xJcImXvoFLqeINz2
vELjUaSbfoOoZYzIETN/jS9JTFh/naCjNVRn2ein8NnCUlqQ7PCSOLwEdRZOjfDh
3NtY2AMER8Is8O/r0uyt/wiGYYO4ysZ2RNoF9FbS/PTZoBR6hXhBiECEElduLtAn
m2U8Iuygt82wX81GC98J8UX2yclS2AzDwzpV12DCMJn4+CMLB5rcRLpLk6rYXF37
Y4s+DQ1bO2CdpDpYVyXJg7gYt+++VMoDGDuqQWo1Mem+dpQpyTVCHPFGEozO9OHi
s7FpG00Qu6jhbcryoeuzQ17kPDLEg+WqTgviDO/R+2p+OTc3UYgJiAWg0u+LRFCz
a1raLnbvapJVu4KCltXQdn1pD0G27zXLMRG2MR+Pnb5zxI64I9wPW/0R7M2iokuc
Y6vNM+b7gx7RnHNZxfcRXRFmvAl3BW+1H0/EglYqd+14LerHN0ilQVWnPYx/L5vF
zVfodiICGTXKE0yqUE3rBXhRD+sPhIINPF/EC+zyIGg0NAP6UIhKqUc8v/r3irqC
eJnVZ1RhjpKhYnBY4WW7RAfajlKsDJ0E/BVzW+4l+zKDFnCgsscDn7VPpWA4zVzc
bcwzJbLsUbXG/WeR56lhMkU2ml3Mzyh/Wll9YyOBSPu1fmmazj25GrYUCdls+zHg
mMiAX1HWcTLwz22Hib/UNzgsYCieBw09vkjA69b6WXCP/R6On4aiEUW2CmB9dq0I
JNjWWAz7gNj3lgiDaAvNvRUlS/77r9yrQIyPVQ1x7ha6XnKBdHUISJa+WmncJp7b
TS9LL5+H0sgnWJVZ7r6qXoJ84amFhjccN2Zvys0G+bBe7KiL1c5mFem/IjG9DmiA
7xNdP46aGijN1Cp0Xu+6Vw4PdLME/5EtPvTxbujlHFanDz1wV8GaE05dDKUml7Jj
uHh+89qv0smXw4iNSKKMVAxRPGBHjaoRT3Nz26TJTueSO/mnyXoOn3MW8u0xOEKQ
Te/bZIvo0OQzJDzy6cFTcAU/YVMV/5mokSf0oNViauH9f6mH5EvRFaGK0OLWMrfr
aaw0azmvsow92Ym8yTe26FGcFtYu1FA4FSu7l4w8Kk4JQUPl6mkRPU50iKPZO+MZ
tsuDq4ZxLI90M4T+QCdlhbC58qI7uw9HTOzkFn6faW+rI/dbtjsmoKaIym2nsHOj
iHgBg83dKoQ/4+O1/tdkOHwRhRlJuSuMqZqbyX/SJ5X3xFYJvoNjEj1UPP4Rb6KQ
hp7P6fuDkQxuyyNfA7i+XqHKUbloecM+KshV54wJ1h5MiEHpxPwaMcDnMy4D/+Kc
VVErnkSDPcPcmQMm09dMW6dBH+dPAedvaubreQrKEz2oMbMknd6EwItps8Zbxu8z
OsIB5I0gVjxzKqT2g7f1agNGrRvrOetic6vOp2s5Rgii0l0egv+9WDREhnW9mWwp
t439A4ATJ1YnKcz1wwigbM+U65lghadewCERaOEVcKmhmc/ysD6H3etWuzC83aJ7
uluBJwTt52OhKSvxfKgEAj2+qgcTaOmS303dSgKNbIi9BAXGtfWGkWO596LwuHSb
1wvfqUvZrmN1im9NJ32Uwqj9EHSq+RTpas6gdlQHqQiWEvEqqiSBroQkIBw7lila
PdSfAnVpg+wGFD4z79ooYJUpOzxN9JCtnLfOFUg0oYTEp2zeW1LEREjq4pCFH1EX
TFU/9X0cwv445yv0vGfYMcgwh2g0p2PGRgAq7W+5DcEYK0H1pRWUHoo01J9/dHvU
S/duXbEJV1Ip0lumASm6FTabxy9GbvvbHsBJKz1EZu/Ee4oAYd5i/nVEvJVSDtDS
P1gXlflAmLVDgCI+ykIODGIAQiG8g4cY3CwfYdHPIKDEC3fLmtjHq4syM6LAZmxa
5Casf1Y+/L/NFkhMl419liNtKNRiQ5fHLk+tQSNTxlqHemwi0SygOOshjbH1/XjJ
15HP12wy/9FpjhCJYaw422DStQM8qppzHMCwFBiYDMjslAWXuQO1VZ5+Fxah1p79
ehvKIOqRZ8Tn2C2p+iB0UMRSPfFkRn2nAYI3hoVBRAHKE6re35BT/YSmBJhDOzzY
V4XURVjUKcq/4ouH5MPLKoHpA2HU66dR2svF1OkIgmRz+8EOaGWt6VcF1pvV5xBi
kDotuzNq5EwgkzVYg8G0FrL3M37SgC9M9x//hWk9zSmDTNpjQDPq6bucW+mHNRAQ
qeIZQuVxPeJFPpXCCwL5vSBU2oVK9nsfRIlcxjnEopKZsdfsDIZk6ClTh8faz89l
DfsNe7u8kAueVD8a+GtGrqWCKeHWlmfZH5DNGGbBZxxKOqyT5u9IHT1LG5CgTsFp
5lESC1bdXsndj9xjc/6Cva3lDrA30cXvynPlrg9c/zcZIZka1YTe5agmCchkerRK
v54LHWSjiaCvdlRqiJPDSdi4lCLq1MVMGyEoEZsybrVy8vJg67BckGMg2/oV1Zeu
cXYPCDcjZs2rLk4GwZwrsZUq2EzRjhr12LSULGELjEfRooYQLcb+Sk/4QmS2AfBS
amn8lxkiB+dHJyRAhpC4FnrIIO7mITBtxku4CbyEGxbFTSTx9tW1PFgfZj4sXFrk
Q5Sbhpl1OfMb5kepUTh0ubVzLtbUrzLnd2um6ii4Y19kBQNnHkeeZzs80CgLQ7pr
Mo59VWyYMvecyIa6f5Qm7EDflV5MbqUfaBCB8Gz3gR3/XM3ERBINW95qHe7VmDoj
lLpgZrvzCRnj2n0zSpAA9dZDdab2rG1K+LW383Bu1R0fG6B22oMI8XZMeTa+Ah45
hhRCkX3F8xZOgLtyLMo9G9ju6/IVhit032epp3MF4R6Y+1CFMnlBWClQle35jNcU
Zceb2Q1yjKOu3jxQrAWJb6wVBJChgn4vCeAW576BPelGIHr+IEcDb7Te0u/qzcud
DeAfmqg/MSbm19YgisW4uw09buKh5+ESx1IW2gd8Hzblo4O62pi3gI0yQr97n7O7
iLDOWeOJ/7NXPSHk5CL9sfLSiTIyk63WU1teXN3J/4Iz9okMikUZVx0PZXORK9NE
NcULHu1KbWESDg14POV4XN0cMiDlsfs2uS0/f70jLZlai1llpYCHMWrZr0+L0IEF
cJMeMF+1PMaBz9prhEUW6FcaJ63CKhw+RmYWDnyxhvY7W2JvA9hkBEs5NznaapG5
0g6xIzNA74g2S3X9UbeSKU0LqDRgpiFQBEB7afvU23BCKWUC3P9MJHoKNMCSAIJA
Xc8j4CsRVBP596R/NZJwBmCEmpvfSB+l7MJe20HPzmHyKdD7uxAsFjiDUiZE1j5D
FsLrhHbdTdaCtZW6ai1elu01ad0y0grSvFaIM8wVnezGxX3uuhqd0hItX79hHW54
Clh92lNRd4gpohUv2Y/uW64c4bCPB1QnwKj/QZ35pX5d3km8ybRdpSQ/RhIdxCru
QRSh1DNo+CyZxVMRpQofX5IuuQGLz9EyH6+WkED+lQv5IYBVoxpnBoz/PhvLOOcU
yGrtQO+kbc+nhkMR+h4rutJPnKUGDK4VExIYOVHcjBaaURaKaelub8NlR4kpqA5p
n8iVDUGELLBHja4PPGdGBz3cFoKPvwnM0NYe1Dj3K6s2iu9RygqBh1YGKwD/1nqh
T0b1uplag+u0w1XbWnTYcoX4VsAKs3wMnEeLw+TAlCA7Il0acTY4uH1Gf3Hn6bUo
s4jx2gfPPOnNzL43U9+JnnCcgb3bcm4boJcim2C0Wd5cCqbxtjK8qmtV4biT9kfa
LyFBcVe1nFyWbjPulmFG0WnxOC11sY/NTQBocWLOEgKgI4xdQoqtcfDM29ZE5Fud
U7TIfupXdOX0Gvqt3hu+QFS6TMi8XdQwp3k8YhylwmtDAgfCvPiyI6uATZze5Mu7
U0RAUDuPm2NGywT44nOp9BCqwbrJymX+f5HcbuUHlmW0nftU01P30wR5/qu4wrTO
jP5OabkSof1t+DyIUxW+jN2LF5E3zB8FIYkqRqTCS/y/vVXT6fI4WMzZyOIULuJ5
pp7TCzQrPYQBVVxEMx8D2tyYqHHn3POId3o5/PfINGWd3N+b4va/rsA3BIReYzMn
qlbWoFNvt0mdzXoGJWlRIifsovLm28GDQyHbb90HzQyDJwCDlbrUUcbXyv1P5DbE
7Qy+xX/44M1HnURZkYDcw7KU1Cnf/mstUNkledP5TE1ir5DqNK/pgpbFwh1/wZme
Ct4MSJTpFjhQdLC7RiXZdfGgia/vWdZ54xF5ODbHwTO09I4LcabKVIdlEZlXzq8B
aj+5zRlv9qvbr0kYVOh8KIYpZLxWlt6I2kwYtqE96CY298N++tgTVK5ONWKXQFgO
tcOQ7ajc8DYJQ9P3jCJDu3L/VThh/OMOTC+EZM4zbzLRMYUkUire8LYGrTXLaqyY
39YQcbtpdvCbLgGrlFuYMYE/MZMfnamRwP9eGxvOjEiS91BFKTXrTY7uVswtbFen
A14y3o3B77OJnNeT4raQjNKOYKnSmlW3oz3hAdT9+2x3+MjBGNDP0VKOsK914g2f
MO8MZXv/jjjKTzKkr2s9k9VtWBFfZeLWRKCG2G0uG7ycyUiJHrNEXQo4BSDjL0Xt
C+tLI/rB/M8rgXAEHLqSQDYFxgRqzztA/Wh1eRUvk4KoxQHQO6BSou3M78keyeKk
3Tb/OX3amg8ElpAze5uCOcw5NTRGoF6iihF8FeUMS/Kpj2+vlJ0BEMItOGwCxsBG
l1ZLufsmsZmYGp9tbeYl7P1WmHJb30QTXXYoqgS12dIGNtfy4WrZA32T307+8wRA
dieFkRoUUi1qy5UJhkrqu/PPhrjJEU5csnOR4rnTsZdbOucHs6FrurNYlBSUuN/M
k+2VLYR2JnqFnzrSz1AXGDNKCDh0NLpoOwJoHgtjZHqGqZrWWtlEdJhd3CzzE7C5
FLKxH37meW0MX6hEdjCAhZ0IHg46JLgyyAwp5CDTk/3UNw/zemZfSq9/CAyxiDfw
i1FvavSpGSVpOqiEFQWMQ2ZWRd5Sr38k/v26vL/g5xqHWGs31T+aKzmeiFlwJ7nK
zkOthwnVLQaoWdVRS3OJsZteAEnVdJu6gH332dreekzsWD9znhrI1x0ZWikT+wHm
LrQLKSmGQaOsc6dTqYtpXEc3OO0qJ+6TNaPsb9JDQvCxm1dL3CEYpCJW6g+zJKBn
vao9pU/7wFbUgRZxl33KOzhPCOlumAC7uu7FOpM64yNl98ofaXzxlSgueQDTrRtW
5vcGtoNWhvjTDJv92KZGUjyoCgDr9ERa7ECsMz5/RUMU4LrL69tXpeCGb12w+9cr
IKl403I92u4oHLHl0GOlKsBNmdEEajJn6HifySfueQz5dvrFnuot/SX99hReukXl
mjRvN+wWEV8PuI7o/ydGlh2/JvDZa8qVjy5ZWP7FTO7l0RYt176OO9LaHn1kXUHg
1LszH9Rl40advBU5VfZYRh8TwOXogNX6/FB4FBH3LjW7egfrH7Owt32l4sEg7hmI
U6f/hTEqsqGmSH2dfrXlZo1WwJTs1YQshW0Qpnm2Sq7KMTJ6tlM2uK4ZG1CsElv7
xfctArTT9Yg9jXlOYrDl0XuHGIwebAzf+Y7Hgx3L0T7wmvAP8Xp/G0FSAFLf+r86
DLl0cxYNAshw4pnkmlAgGxy5FL8HNb6aKh0LA9nMT3luZhEmTC49xJVpKTaEw/p7
PUiLZBaBkPSCxgrbGWtAmGZ6v9CcNcOX9S1JNGEtzatq9jRF1N52L7VDc3Pv3r5f
YlnDvS7HuucjpR92ad1pDmGs9rCTdI77fX+8usuXfFD0nGZiRz4APK/U9peOFwkF
HcbkAo43NtEQgcKii/2ssb9d8R6XuTYRjpGgi/zZCgEjIOneWyrLjyrWK4uONHY8
x5qVdwZLEMEAjk6uMllVJKabV6INFtE2SqRNarXeQdn7SgbQfkw/yMMPTOenoztG
cfHLUErPGAyv3YXZJsGUBk8f6n6OR/oZjPyq6LjGUnaBI/UYr0VfgP4ASJb8ePEx
KmJM9XNxJNxU2Vj0kDk6aCXffT0VuCAKllHCGyC/3CVlHY3IAMsbGLEQjMSk4V+l
VwlOoWY36pUqMvxvV8yeRkZrsgA0sA+EuFsYrBjcl47KThvijcPgciz7SaVqA7w+
G9HDOanoz1S4OkK1Q3CxtgN9oNubJX3/+pTcYjY2ffM1IBQtIcqcXfD9pLZdHJaB
j1p/WK9tpx8YRP2hE3j1o+23vt/qvUgsN6SA8iV7YzHH6V6X7HiEzMjpHaG1UQRd
sRc16c0kmUgdD6G4eFfKlnjhW2GvUSuHD2MH3n64PmbE8FMiVUMzDIsCzCEdJ9VY
1bWgL6yBTE0Nf5XIqduOQkYsCUPybQt0/b2qnnbI93hyjDTtcPBAGpzuidrvR9V6
E31h+XC1sAGhwBKiOLKlhKYWxFbRWg8sDAqT7r8YsEhJ6B4T4jiFEZbguBW07GUm
RFzH9bVUjPrxSfpkx+CgCJZhhWWz8izmsFB8awJxgnkf9Wy+LbZ8JZKZkB1HhazK
fZqBc2BSeBbCu7/Na4DVyxXdB5N9KjwISU0K5SVhBZ28ENT8MYZsYcItsBolV7IS
SxAV6UtynnwzFDwCy5PWbkowMjr/kRAyAczwNIf+GrGLSrPpz8hke78L15kcA585
o0wgVR2uiIobtx2PgHGqURiax+bvGXNcaIGvxxe+p9/F1PLIFlgGE65+pYsH7RKq
4BZTNPpzC40+AKl9frd377M4b0eIGYUlwma++j29u5Lc7FRSxCe72yeT9eX2Jey/
+e65GecfW10qtzw1uH6EU73sFHykyLoiXOO3kWTz0P1ozoiU2Fcc+BD36N2P9h60
hJEmlOHlCsgfxwHluQ+V7xNTi+XseRHLb8Qe1fbtjQ5BmCZBjPJvWqukLE0IWOhk
hydvj147wMoLv2QrUPxLU+5ncIpkmAi30mwvXEGkNc8+RzT9Vk1FUQjauJcDNDIK
PQtMdp4WXamWQqXwwpulj6u7ikhLwqjNWz7EsYUPw8dQxS7Y62NzVt8y0YqHZiZa
WUsxliMb0mMt14aLswJgpY50nszBnJFwcftLyX6Aye45z4dME0bMJbVVnNSb580q
AQ28cmakbNpLn0UEFnC83/R9cnCWjPI0fd8y73kooiH7qM7yCurJwQKpSLda5OUl
w1Q2kd3mTGTqE+7akKkU+bz7bJZ5+3eQQ0vgDC3T4oLqcS+X9w1aduSEbvmusQKZ
LxufmB1r14ulIe8SDg1FJ7SwFA3y/45R8ZdV7c7LXE9hCegc4g8Drwz2ciqBkKiK
BB3ltZMjT5QtsYtbdnzxkUUZg2esWhPVQAyiIR6HHESPwOOuJCh6BAmxNBKHaAsV
lAFSkpsvJULfa6747XTEg8EHI4u+vjQEsAr2GhcBB7fGCWjn5y4Hactuo0LrPM7v
NYGbLoDQioA4U5qtbrYQdZhTK7f5oYlqzYcT4prp7gx0+RObJUNpQ194W+/iF8Z/
wyhPuuGgRc6oaf7FfodAWaPCxtpZx1pr9XUvVpnkLuW1IZGZloqup7J3iMwWNZOy
KgsXnTD60GHR0h1dGWObhGlEqVrqC4XcUKoAZ7O/Sm5bkDHh6ooXzssIVpCepJLW
UESSMgHBgzlZWsIChyHUDmVmgEhbWeAGSgKMZMsKXQczoN0Y8NZltrmThz0WevbQ
ICsXRRoXV8kPsjf85zIo/T92asJt1gYg8phEiGfL7K1g31pYoIEKtt36HTuYHV4w
/+MVM+tjO1cxDS1oQf+LHCNg4ddEdWE7fWzx3wA+qRJLAIqHr3FMTwlGTNe8Wu/6
8Qw1Za6I4InNlxPQ8eGXy9xeejTUJY68y4Ye+afymaE+WbIsvNT+rwTUuXivzSeb
eLzm+0RViziXOAC/Ahzk6c0/eg9FvWaRFJfAHP4BBik2iYL/VN1rgot3/YfoXSw/
orAib/Droo4DSue1go6kNHIs8na6r6kOOWJN9RqF469S17Um7qFe+gIUY1Rh+P63
QUckt3GGtVUvmLhbqi52gx6GM3reJhZx30r8uLOjCsqTipXEDGijdu0Qe7cTZCD1
wi3DZPiiKEQzvwUFxDbT4+WuouGW+Y7089tLrrUDhjhn0lgTeni92nbYF1goWHfv
jyjOjvlVlgHcyaA2Y0Q4yybHyWmgoiT2V367ssJZGb1nHmEm13kRJH8ekyJpB38A
82hSz5dqYVNVxzJi9p/qNMzusV+9+n6E5Lq0J7X0nXniPJuRC5A5cE6YuXBuf5iY
LxnwI6Df8txp0p3grMJsCUUXO26qe1WMQ/MfY7YhE0YRBYMvH30dhl4hlJVlT5tL
rDvtbpuCaGO8kHEsfkvyBH6eBL1z68xEmJlw7NFNs2XII55TXrDiu6i3FSxBmiPj
z8z/bjbOOStuyJxQ4+8xjN4QjRdG3ImXmKjgFQJBVDIKIIiWz31GVPRlEzEmY2p9
fkOgaqk1nUKWxGAe+EcCiXjqwVDy+XnjCOxUe+3ftgsi1gsEDsZemk8F9xJrCvza
VjQIXMZok6Z5xWTXywlsFAvwpg9Xvh3KbczAjxXBETfryf2Mf25pw4OL12JZk4Lh
SC+l2T9Uu5YEAgevS+TLP5NMj3GrxMV/ZRS50+YlIPcmBtsNfJ8haJbOGeUbEc1H
injzxMxpWvlA9z0qfopzf6iWjhCVRoxU74KAAhwh/qOaig0VZJTkVZKvNb9p1cKT
HP9TRixGwZ+D4nJxlWOtfWTENP+Lb2rbkFD9bvyhKFDrq5m2batu9Y8NnLhOhsv4
8bBK2D10GiSlMp//OYouNmxbuoE+pq9Hd9NDtTs+5e0lS4T6fXRF3qBm/uv1BV2b
W9ugWLNB9RDtqiK/66e3Sel9Nnh1VxHP/y1jRB9Az+Is+KEWSDjunUyB6zH4SlXO
XkKPHUCoRKtz1u0JznvVSfymkB50RAPPzXV/bKsRP8mTR2ziiOoGZBMSLmlf7NGB
b4Iua+Mew1YnVeakEFjB3vuWMIejsoybmOslYvIIDgL8d6ZGBd3J6aSfgGIHcg9W
CWZcQXhPxZentJCz4+90RLNYhxbAxZa+snIdZLTxLf3iZHsToJk38p+yLi+Q5ujA
5Y5q+GIXI0j566JV3VaWsf4pIOBQQV7e3SMunwED5K1z2vGo0Gusu6bnM8t/ROHp
InUMaKs006ERE+tOjDDePO7E8Hpus1H/cozhbyiEK/jiXMrH/vlRHzuPT60S195j
/5SKEVuZoUZwwvhPD/6Ee/RjwSRFwanfs1WXGj+8YboJ5D+B/9dsuXTC22LfcelR
BneOxC7pzQ7gtNuSaMEwWj68n/Qh3ZJ1d2kyEZMFjwVTNrBdRlFpkET6wgO78F4+
F/a0MrKtxFg4W3ArUpSuO/t7zw14ycMSKl5GVgxabXa3EbHFkM8sVnCJ7tGsTCQu
0pkidCkkDNfaoC8KArxKQ22WkeN10/vKweE5v8B7l2HDtvYvC/oeddqFeSbBT39+
4bepjBYTL2DyMQQB4Ufn4KVFCiQwjh4a6/OzFxi4LWQb+hxl3kLa1pfwK5H2SL6R
oBupktMff4QyVrwNNH0RAhwUWI6jWPQAt3tlbB7Pbqgo/9+2q3g89BI1O1ACZNu/
k1oYTLdxXNYvoFT+eLXpd27QGS1ri8fblOOStjmAeQ6FsZ/srKOD1Z+siCGGgegM
fsHLD6h3fnzmvUFZBHFPi2zC6iym74kVnk2XIZD/juODBUlEr4k5AvxZW+3h5Mu2
68mztjlyDxWhpURcAKS1585OpCeTw6GeDNtJx6l/lAdODsNdYry0qcxdeZh6xUNy
PcP03sxT4uOTLfk7d4AesYaapbkUagTXCr5rlhDKkORsvuyNm4KBHZgpRCRKWcfD
uAfgOlnjKPL6naveIoG54c/GLl2GTEmmszYY0tONwHxGSd2mTVNsA85MG+Jm8AcG
A50Xbppl8NwNfl3OAajoukWmBrAC9vI9m5H4tRvwkKuSwbuyT7AprGU4JBCppkFT
8Exa1TW7b262NMDgzD2FcGHSb5naDIWFSeOokgWF23SGxHFO+gmYKTDa/7G+Cvxi
UohWWhw/bOfVauZrWalZYbIvd/CY/N5ZV3v6zgwo8/jC/JEeo0ItXfDh9s/DZ3Ke
rsXhShFrfm/ohwGjrB/6n5jppIPJ4pdzG6rqC0T2EK0ta+OKrGeQpNfr3uecbL7s
/YvL71gt1qZlXTvH+P1Z1l2aeudQEvM47f8MOkEePsYExZKQyj8E1grD1c66DQqF
dG/lGREwgWPWuv9dhnhefbpZV9sPscszR6MlnuYBlnQl4zwZ9I4/w8HDG9mx/7XW
vsMnvkVW00BQCSYZoQMldGZKPEGLKq/fkPvD13vSXaNd7t3Ou/bGVciubsudLkv2
PESi1KkCN/gbQ1KG/SG0YWMRZp2zxKzNoxhFIzdFMU4VuH82CyjdU6wPleftB+sR
Mpaaf1DCo1e9L444+rU0vFY9+sJlltJ8NebmOkGSQh95YAnecLTVMSNxba+jJ57e
M89dJEVH8kOJci+Uzs35wICF2tO6xDzf5qMeTW+XFXkMkChXzPeRDZt2mtZBwCSa
ZWJsInqPfywJdvXGsbac0teO7WZJuP8NtkmPj/KX3zrT4b8fHbasslEBqhOFSMWj
uq6qqkmRDZo99Ii3vyXUhBlSNwkGu5Vq1sQvmz9xvrB0CU5iR8bXnbJSs82pPR9K
RF+5X7+DrtZWpLI/CKvNPRAeav/K56p9vIofA36n8CJpSg0YBcGiYhWPwgayfkZA
6pZ5qDqyppFyYA7w3N5iW0c9Oc3h0yYNqq99v1xurOd/VqmNueIexe4QBXz/4CQK
RZCtH9DkAdRk2gP3bjuJaU+ZBbA/dfMYAAzLLuMHI7gThyuKzBjVY+7ebCVzi+r+
i7WtZGb9l+bcJPxTrOBEJhh6iWRdNBWCkvxLMB3UiiIR0r0j9vR5tZ1GLc8fwiQI
m28I6GzPCWNlwBxc8CoxQ2hdIomRSw7sSYFszIsvSkbhDzGDhBY1KZdNVdyJoxOB
xktan6nMGGSUah0GogW1oudO+tYCzknew7P3/t7WM+pKn6Q2hJOS7Pr3ZXk4usMC
Yh8MHmUyVnnb96cd9xu8izVgE5eWZwe6pQLNy5dHNgyHWWnadwglD+W7QB2heOdN
9iCJlmbbp22YuNKKIn1gzjoOorjNNffyfRMHuHTa5LBtpNKpkGF/2+NF0f8xYVYd
aKlJn6tZrNlobnrAa+W1DW/deHYdfQx4dY4qBtPyELyF0RLeF2yZAtyq82uCGmVx
9k1fIwRpIC9a++7wshCyiq8HlxE7DyzF/hsNwGR5fNp+C+YBMCvaqfLRqRN5/OUZ
1nzS6gBGXcXWybFPi+Kdqnfi0QGP0lbOwo2jy0OCrKm6q4MrPeB8d4fQHC1iW+A9
DxmrPqsa6zMBvXasW6Z+c78fvbFhPOuWftBMAFol2HNJ57fBJ4KjJTKzNGrrzF+M
1V6xcr/eE6xs7cQcfWugbbqL/GYpwdvCbRCEJ0hvIXlDnHUc00U9buhvQiiuN7kV
BDI2IJAiK2mqaQkkmU3P+vwE0vMU4pLUTBRRld8qZsLSv9LoJAVCrwLoXHqtzJh0
9CII5KrGkCiqRCKDW/6g90/Jby9Ou52bmxEjrVGIbFx+AG+CJEl/844XfROWgkrK
AHflBTTS1MSItUGYgHhyx8wI173V1/E10Fh4UyD9K/qP+xzqVmep8cSRrcLP3Po8
HzMhYWcdYyRyXINtLwvL3e8fcf8P91+NmzPsOVNObAWiEtguGZ1IgGKik5ERrk4X
0rssp3hP4hTRsFokkbkIgIuxERhiNyHEx/O++Dq+m7oEt0UwkF5WAoyNSiCsDpE4
vUi3YVJd3dMwyogN30dZpFOeNTlJP6V/5fq+jafu/mk30TKc0v1jdbeHMS26rv4Q
xJnaMO0d1N+6Uv/SCeejY2HjwKSAK+OVBZS+v1bOWzdJPrlN3jpAxefzJEdw20cu
sSe609/Hr64xkdSAR5HNJMBxcHANBdxMu2BR4/2BPqC8OsHhTQ6BNZvADP/R+YrT
VBKsVqpjlRX5O7Z4HebXE/nvm9wGAtuSRPHa5FTtEXFNlW67EE/rV7N6OM/AM+S+
J4XEhhmKv7huI9YEB2q6JbP+JUf/ulRQcyRKE9aYcZ5PEpa3jg6Bfzu4OKEgcwBa
J08TmnFEC53DHiNH/4mQbdaIxX8JWBDbSs6l06fckM0+dSjlkaz3PwXBhVrrbh0N
Tv1Z5aZ6dqTxv7jot+9RMOi5RSOZTjE9P+oGAhCBF8eH59OIzZWIsoebf13+F63V
5bBkRa3bT4u+/IigNvmKda6RyNJCGKqgQPgs3CCm6X/0TeNxRHFD5d3NA/rkh7iD
0FqIVIOKJxMeGAAGNMAwE2rHx5Fb7Qn6XwtLuS8ZEnsaiCHGk/qePVlkVMrtWEoG
iw/Ea14bUjNqgHOrbFDkTfVrWCtP7uex1F8zIzLv3cga2/SqMMJW1+RQh/SmkAVV
BnSAd23sOcAKvEki6CFREk22YOblHvs/Mo1N05EkAIAktPjDK4cZWzncbhIYHsFU
Zkyve5aap8V0zgfAVU6v/sj4DZs5xSpEcdZmPUAouTgjDavfrU7U6DSGHMLhs2Xi
Ud4YLToa6ha1aRIlKxHh2lIAHDMRwSG5uMDSGQVqJwD8mmPNuGDyHDT5oKEg9fLV
1FKDQBDgJJcoe/xOU+UcTE6qfF6w3gtKyZWbPknsJ+NwMbcCWedtUohucN5QF6yE
/5H22Py5yGO8F/xc2Go/rANZu83YbCImy5YN6nibqT1GiFQGaXHg5X7niEKYbG02
EZNzcvDg4Mulid6HI5xoV0fpdYvDi3JilhDlVT9Gv62YVVykG6/YOHQYry0fEFhk
+0z38uNeUKuZ9kdqfdRK0KvL3UTrdR9lT5ZLZ34insGBIaoPaqfISXXNmjUGw2GN
eyFjHvhCqLL6YWAhMvzCOqR6cWpFBGNFVhpl2Q3MTDDGjzcBeorEgHLCL3LHsAio
P9E7a0NQa3kxxfuTbua9X9QlXrMrrWeAkKEpMfl5AnkQjQniuvHmATl1auhn3JVw
IqJ4Hjsfb7FdWafqayDLPW1qg1g5pvL0oueK6tzNGDfr+9aPeX9WH2y0lSzd6RSd
TcW5L5Tp/AgrdqqrUhLLmUw3JRm++9YXTAfBTUA0azaBGXRawlqclcheKjTdWkxM
jkcnK0q9ZwvcDY46y7BM+ygI/46KJHldxnUUTt76gLgSWle/H36JNNU5T286xInB
IcWuR3H1NgfUsHgu33MXrhZgKVLqEkUA1zFVzjGBmpX9Or7tFSEYjKLbpqjtsvaz
eqvfR2NIrvfhm4Qu5kCWD5ZvgqMzZojr9/vr+ojfqjbQdiJQ+eVJcvliw0C7QSc3
JhblE9TCgYOPeuHU7lTtYxYs0gYcuwQxnGt/pDk4CDuS3vC6+c/XiDFreX07l0nd
AgWummvXdPyKCDW6okuesTzHiCJU5P+g5LhN/+GO/RrMoSFnkol5ZoRJg7RmXIHM
hIka3p7FV3+Lr2cGa6O6FrzWfMdNZQowKE9P60dP/A4w5cnZ8DeisB791+G9wsG8
WP8zFQkGrYKzWL1lscu6gsj4J8kYn7QDMmPqJfgjWWUiUXBITcboieLfBXQnEsiS
zY9PHqneQN9LRNFysg4aBHW7soZ8ySLmfIXElSvZyFvQKguqtyCNubU8ou+5f/3q
aBBbRgn3tYce7Bx9K+nW+SY+HA6SYh+XQwGRsbhFoW9ilOl1s+ckJukv24FnA3uP
rRns3py0oBwgkebIIxMoDDvK3UeSP/cmWZvDC5nw82PSU7iUuGeSyiX+bcibTb6O
Isve0lUpxTArdqHw1O5n0PIb/AehuRxNtW6tNUQgyjtcCiDtW5zSeixcPdeP3u3M
cY4vWtLibYzCA6jCDMxtwClDSX0xj3ybFEtyRhrcKztsXpZekekPaCq4DMDqJIso
HD2uIP2M3sH+kL3UrC5BOgJiAbadm6nsdfIhDlFzlidSNH4TBhglxGOIpmuDFq+K
tkk5omrtbifL7I6yMbIpX0thshDDcHmVsTONXUHNY1q7WM/aphlDgBWBRsifq0Rj
YOMmQ7BIUHR1GXKBPjID2+XC527qASduVyjh+yr1T0HRr2yBYY0IovOXNWmQSz4M
IYgi7ed0JTe2eYuaI+5G2Bz/ma4pXmQC04h01p3QS2hSZnhEkvMjmdd8maIHJrkU
VZCi19EbPs4O6omeQJ09FDoDK8K20JqVEKXcqek5PIkxr7yxEhimqpB+p7Y8gPiQ
Zf9Kq6z6Y3Ys2rFHAu3Ss6QREl19phfEMhbN6tnkRHAabiSc61AOyGJtYC7VYgzQ
FM68rhtZNduMfU7mdQwoHhbPjw7LsER8zGAT9P2ZOKNKqMpvAQt9qc1jDDcE86Tb
3aM6HVAIxxz99ypyUZuxqvhjGtbYHIpP1uuA5Z8YiukYV4FsRliiEEd6Y4dXVvYn
PQI4l2+18PTp1j1Bu3MvSI9G9RDIb9QyNmkDyMjE7pV+akqfyXpl6UY/0QD8V11P
iAZUjDsoGg+xAwSAu1O+yJ4kAyxeUJzpiQh5eArFbHGX0yyLnGnDBiURR6qz5AML
P2S/5HyOdP5hloN9NyZKlC8xllvUEhoaYZpYH5heviJ5T4U28DOv97VusTptZCLd
tHumpcI046K7v/xsGlwRsHEXfW1MYrsF2zR8boJG8do50veyO6t8cDu34ThriFN/
n2/Hcaknoj7xKy3ixOfzoDwRFdfiS7Ll1HoC2aSUCp4ym+68V6OPL1Jz5/7jdhXS
+GJbr8TDpRt1+BwBa2cJKBjhZk/rPGPbCZT94nhzff2zWcu7ctWJecYpfLf1kkma
txepVAIQZkck7TmcAD7qpzt6NlMVxuhZr+X/alJWzta4RAHnalYSNQdjPsuhHPSS
aOEEEL71f9tZX7oRIctwbHJg7zC5GOGUIj/PNvD6yBZ5h7U/4rSCmD4qL4pSfHlE
3k87CAiDH/g2sYAQ6KxAc/F0aiEbccfXckFcW4da74HWYkBkW2FyN6tpg4Kks8dB
DwxvoNnsmtRhbqbxYGPwcnSBSdIu7ej8v7ug2JaqxdyWL9P8fIf92plScbuWl3iB
cbuefb545gwDVhfQ1UEaAm1psUaqnKQ/LN+rkNa4fL9+uP0rSaplxisp/oMApW49
KpfGyCu17bKm2J8cVyoR05NfptlxtoEBhiYoAtz85eBm4OLZnFJ+E6Fec7uGt9n2
1a7TUoXd4nkRMGFuvupXtfjriG1GwbDbQRKkejJA6MgVfnOW8jicKVR7Jqe3eg1+
UcqEpePuj3A461yEtXUXG5BG1T844FAHfNwMqij4PMqCkKNwWe0fE3ufsrlKrdw1
z1mohhXywMK9x9UNupo+yO6DZZVr/qjaiO04bmTmnsTtkylnHF+A683PmnB0ttCQ
7iGeS1ORrxifQHAfDga6VFwZU+nntB72ejh0Lx4InLOf8T/Hkv/RyNLcEMymr+mR
hWV5vxQcXz6Wf/7dktVGHABu83tLYQRs9+3F6N9fh7hRAy+pAvjkXB4sv4dlY3mZ
L8lThKQwDenqMzwD89clpatsengt+wHzNk60bXhBSqFzbfqWjQq8G7gqPak1u1AA
m1EOaY2USk/75gh4rLW3oumfx5uPXEPDxuS6XDTgF9SqcexnBbZk/czkSiwh4lZN
RUV3Qde33KXk/eC+PuJf0aqxTR3lY4Qb8dkw0W0Sf3qHLHas5jAtCmZyIS9p+o3z
jsKl1vQC/mEYaScR7f+4lelY5pdfLIqgwzveHoJrgpSJwXlI/qa69tEjQUYFADpZ
YPqX6ojfEEJe6jJoUXjYdntI2GKb9ECGIWsyEyma2t0ONFOywl5VifsnS8Ecuk6D
ZgzjwmPMoYjDiJVQGsWheq6LryLo2JGnmiCXM8Q8DznxeiFk1G1PxKyARU94IIv0
V79EQQAOp9eTfTHPaaYfIkyPbG/ZPipJVunxBjpz/J10KNjKYHW1sN+D+71RoxMK
f9Ej0eBdZnHJPlVVQgnJ25hmBf/Opi/Q0AdILFq9kzbypGMxpGQJHtqkvQExxKWr
4IRR9arvFSdINovyYEMKV0jDuVKYSsv5TYqNZwWk0hGRb4D8zBYbWPTxOuEZENM+
ywlKdG2N3JnMiUSip5s4gcZdaZaMFS+oM9cwUYH3sWuDrrRhGQzOXZ2LOeOY+zHV
EfytHpspclbQrFxzBC/a5vO0AKwQ5AOzNu5Sf2Ntvmyxp0dn9spWQ4XeoHjW+3n8
aWVumjWHrtDTMljEbd3/Sj0I0xQshpHkNb6SWYUEHv3flseHYF97H+WXo3KIwT82
WNisdaCZK+VMnj1Wu8Zi74mNKnWn9j5KJQh5GVEUSLyI9qP+eS8RTMGneFFGMycG
yapvI78H6aff+UFWnLK2oHP/ScmfxeMj95aqgXVQeTX0mRpxaBvicGzkBwB+gN7v
51dli1BhN4aFETzu98BFRK+VjNt33Du6Q9q35mJYkKUw2yfPn+vo2Au3NjKi4j94
9irwtH5GL+mvyWUoazAE4gjmrHss/u1zFe3tmfWoqyga0SHxO8Z7WtFR1xYKiL9n
RuGQQcweRMEcuv3hthL3AslxId/X2VMey1hJisukAQblTH0nDdbn+nbBL0jzFC4J
1KRnPHfXJVGlZM1IBlV5lF9Ea/0HdyIf3rsO178Y99mWaRRprSu/7mKP469YUEHM
QFkY41RJ6d37NLOAWOQxB1c21ODZZDc/T9IWaqZjIIMqa6dQ4PiVJy9YMlIB2bXU
Bowh1ZK7tRDwSV21M3TFE1ZGJAlx9MH66/8iSRjpKJXKYCEwZ4G5+VWvUz0OKTKz
mw0jpI3HywFsDDBzwTLoNRvzWXKf9waTA4IJdPTKWC+PZQFaH0/Cnc3T6sVh6+7X
bQ3PKQW8WV7FKH4H+//uqzsDnmaqdQbVNFibdDohV59vRb3rso/QmoBvLAtTvnCl
cNJjGfladc6eN88ViPoAPM0UiJ9vTx2Ob5eQSgsCjJKFq1LmLu2jRMCqGJA6/V+e
RC+R8dYnB59e4V7IaYOt+PT3xrzTBjb7doPLi4pQojIUh6m/jYXk8o1FUN6VFXhV
M4b2I76/KVwFZm12faU2zAeRyNng0DyzcoGcKmCUFbeTIiota1CpI6dC5oY+RE4K
mDOpS0KHEKONYKtk1UPznvFOeT3jS1sLmG9iqgBkM+rVPMbJnmSJaJlO4vudPZWP
iIweRQ76gJQ3w/Xtf84yMqODFjgn8gdUOQhX9dUEcGghCFHbbDoGaFk/29bYqpXl
5vT7aS3tAkdsg0U0542M7VilLP6Walkn2XaTxFC8H9aHZEiQ6NTgxFjzzfIpowl1
nRdl3SvYevv8qtcUTN8mQROCVGf3uM5WCHPDvNyGHog56mCLTqU2PaWGfLewcQrO
LKaxZKuFN9GRJnjZCtbkixNPJh5GIHOyBqFV4/yoX6gjHFkAdBy/ILbciWWzZOWn
ZOIgANaWuPtjjKvZ58Tr1psHLeQvLMfVk3L1qCNSVDnIEE9l282Zk845RP3SKIkk
Yo2rJ9L7TEsYG0ZtXIMfe+uugTbKmy8EB0chMCgS9ikYVxuH0+oRhQQnGiKwdmsu
M2/qLuph+FW7HAZmP+iyb1mSsfKL+ZUML1Uge/bZsOpNoTwz9EPp3FoKo0RWoy1P
FHa4gsntdCzerkkUcS6N98TDmMazXWdE0HXKR14PEDihNVkcKegxACCUn159c45D
J02/keyT6cCNVOgV6IXOiK/BsKS5cY9/cHg8kcRJlTxG7nJW387rFf1usZBp7hmY
xfkKkYBjNWMLAhQF3DcrGhhgDFIn5V7wKmQxS6dScdzeMX0ilhhEE5kgi/8ACv5o
sRCdAgzLWzfJt/obE188zE0jQJ+LR7p0vwjh+HZMoF4/6u3SnR9l8WIdZ6dpAhZE
tGJxKhnzc1+yY/kS+EfIthSdjD7p2yCjsrotoE2Il9ftzrVeopWVp36YSNYE63SF
J870JfC11mXDnCLVLCm4xCiRhUQdELFKtN08r0CcjC5gsRTLeQ8zlgN2mT4iAEzy
XX35O5xM2W4n5GJINr5UhEvPu0U2JRj4EYnyFM266cL4pS7BvVs5P9hCOzHt4Pdv
kSoRHrH9OqnzluKgpwiBF0HF5yTJOEUDpTplQchbWtaXuVfvtq8VrliUQ2k+Re2x
mEgGQVkC3hcQSNEKQMhyH+1smK0nEjdI6n5PjWTzTDxuH0rOdfHjHEyK8KTrTYqd
LvazO9clnpoGzR4/oaP+UgxUKvdItHH+A893yqHyzCGsXsXdXuDBPGd2a6KeBv2J
h6k/Qotu8wPFDoPmrmyJamSx+19z/RDXiBQ6//ojqXWBrRu/Z6HoyE8EpdGg+Cwl
rskkpCV4zea7arUhDjxW4XLtFAbsBuFW2HGC66KOk2BQIiqnQ4/JG3TgFmbDkza9
1+jvtjWRWNA9/APw1X70Su6lmFRf4WGRIQtH00cUNLBDWVnCt5cM5AfILANBI/dV
uVzBA18ZhdGyjNts4lYJikgxHDS4TNiPj9oU2wL8iy8F/7ZBn59B6mIpM89FBNZN
brUbcMXBb4SW/tY7sWvfWfSkKi8I6axyrRBgVK6rqL4qjv/6Eo2A7lANg+iauirR
q3OrQoo+ZAUUy1MaXuXn48yWZ9m+g3epkbzzMs+qk/xA7Z38G3DQglwfti4wHNak
wgYLQ6wHqVfashloKNY4BukVOUVqLmxy/kAoHY4Hbwo6EJyYQaIK/6AwqPxjmQHj
ToNKNQKdTo1JeU6En1gCYH55ljIyXKPRSWLtz1HGuhgngEPVvtUPJrPVEX7itMBD
KVS5vul7m3oO5r6fVTCGZfrcObw+y9B4hyNYe6ZRCGh8gDIRSore+lSPIOuzSoJB
0ssBEA4tNQ9n0TvFsPI3ZoKbzTCOuYTa4m4+MhMOO1Wg37w5dorAfdzLkEw6DT1l
SLZRkBD1KZlWYtUF2fcqWvKxLCSLTNtaiquOiUpJiaFUwAuhT/JaSayCOqVfN6Eh
hZs8UxXZ+Nx5BmWWFEroU6iEBE1QaRsEL1+pm+yBNH7GcPhrQo9SXmFXPvoArhtI
2v4/ERABMTMQvKnoXRozOKFlxHGQRaCuHJoiSvVPvRqvTKOadb4R+eyMv07zR+jk
HonxEkjfvl34p5rwSBXxztaQbpQyY6Xhx/MBGQYc6wSags2f3XrC6tQAIqE1FWYo
nT8HPevhX98ZuLnav7XexitbqeuIoItlHwYqzbZ3Ta+oGBGEFbIDFQ36qYuP66JF
oJgugg7BHIaxa+z4sZhIkFdnY7X+rvcSgSKF45/NOZU7c5BXSDVeAC85x/WVMk30
Y5NSsTdc2xK+OJQEKXb8X6nBycXczcDtSAfqhKkNC0QmlW8MKOrmCcPbw+e8sy/Y
zntwHEMRi4IaGsBDM9tZ7y16SMIHlGlqMUmn04I8lziwD+9H5XCBnmuIckNjBfbJ
CR5fJi28Of1PLFCYV6XLYIjYh5zBD1PjjKcKbN+6FgVSg4Dy5snjS2DCSr4C1biH
E04GBmln6kGCGsyGregUD0atUpTiUBbaUuO5nKFQG0KS38wv0G4Hz0ZUkjis0oZ3
WBmQ55cUzEJXEQtR09xfZP8Xt0R0p2ooSdk0R5REjwD7Vq1RsQOt6HdFhf+NbFO5
AOHU4cHSoCOWygAC2t3Bog29WW1bNQ5r36uQyRzL3i0vvdFMPTK1m2wIxI0vtwo/
z+LscudO6eVK25OdI4NDnt9pWpKOnyBmXmFz6zMNWUIG5fa/Rm4mNZoT8101fZg1
dqfj0ipHVzMv0sO8fspczow8AliSa+tleRKMT1AT11sZYiRakJLCJre9L1S1xeKn
+32wUoVt1y1Os5jf+M5bVg8fh9FrUg75YmNzcjsSOmEDhtW8LZq6ZqiYUGibW42j
DXblZTEXSM8uXNA5RF4awbhhnJz7wphLXdG8E0NNkeWARsGCkCYOTbNtzmeQ94Q0
sU0aZBGAQpx/w2TNpCBmm5BNBrObz7HVzoJl5JlRRP772R63c0ztcBkAYkZDBFNm
t3NfV2j8RNXlwSvFaVI1nK9mBACmrlniTpFP8jL1dZOInwbSLA2QBOeOsqT0yne8
GuPCFGIr4+csFAmcQnSnb7ShOBwEIKIGdeqm94QZHDBU20XIPiiRtF4Thm1SFq0X
T23XlTFfFF8TDtSMeYZeyKQRFUjC/cx67senZUkUvvJGjNAFVVVyYgPVzirM3rCr
cSjY9BHYYnFqj9iqKJ3j2jGLmmG1pEL/XuRd24KSWApcNZyokEhyPrMk8uDkMIBq
6jpzVwvlC4aG5XF1OYdcKw1oOCXKf/kqndI0JmTesA7x0njlZP8qjerkO3M+PvmD
Rqh3a5iQaFeHlkGHo9VQ4FvGvYRiefhpfem5KWXPsfiMeIJlYUsxlCtTSt9wjGi5
nTQ847LKT/K5uyPzUNM8ikrgIYE3bRxGhtLXONoVlVa5Pte+9//n1wAi+vRnEqjV
nF8CKZ9Z4Rkmij0J5XniN6Yre3eCdJBgRb7McIsD9e5ki+TTJHLob7lqGdP65ba/
ArdNduavCH264MagL07eL8tsEuKvwqcd240PA5iQKHZ7vPupvGS3W8yS4L1i1mdD
cKiHIUTYQfHM9oIuPqRlgq8kLB8ww1BkSd5sXPcujK9VyuRHg3Th/OATP8c4ptSq
/Vc6s5CleAu+LLEwRO4r3Uu40dbgUA3EWwejxTjj6UuofAZVWimsY5a96AEeeIZM
OtrN8SYLee2kM2J1h1cQLezqm8vv3bhihFEgWb3nBM4rGYw5UIfTzweM/exgv0On
BCyqq28xHcRoJqPuFbLBI7PPO2YIUGbLi/I+7RX+vAZeGpqpy/ByWu/lkRXo7dyX
6f0n/nYJcaEiTOan6tCaXg/772qVl7naBcfZ3Xd2P2lQ6r7Lf/L9n/PnN5sUjgwr
VWd92Y4rRvzQssnAW7cqUwtAiXrphDePRR6cTEo1uk8U/aP80xpGT4ZDlbpFfULO
H4HoDzfxMlx7bwhP7Ni8YdES16Bn3IS0nFRn83pPZUSlTpKav3u3yyrLk4weJFX9
bk1rgWc60tLMbMIk9VdZzbS2eQJ1BTsO4AlGA+pKlBcwVAU+jyKbVkwia+zRT9Xk
60W0o7bCFKjPVe1WU7CEwesYtdQ+bfMFZQbRHcu3sMOBHrQFCQx8Jisg30t+5t6t
lgzXGI7LS6mCmE93BcjqiNKSvxQLQRPG87ydmGlcbu4atC98OXylqycIzrWT3AIB
xoDJlfq4S7NMP0n6OewZISq/XElsVrKK5mZn1SH+t88a/jHTsmQbzLTQK9Q+tBze
qkiztILvwDM8ZpkD9yldiv+HulKAmWIj+u8Y2Qy2P0XOyI2DHJO9jVMWYc5HzKfG
O+A0C82SzzBbKgShRbptFar0jfSD56ZMinix2ZMdanVm3zJtR9HU7AlZa50sY1wu
K7IJnKVtbkkOFPrUA5coVsQdjq5ghghAfFAnfRclRhSSo7YBkOvnY3+l+iK0oR4Z
K+RxIa7r458K8skHuVIw2lL34n4ElJi4Osz59mhCMGlRYpLJFXd4Cj0DIGtEeFjL
roCjcd6ASRE9l0oq9QkPppwFfOse/f3AOUSu9pgRRWMtiP7vjThqcgp5BMWSLHw/
uDJKUlzMRjg9GaY0G1ALWiGVE4xfeUv+WLbIERT49CsYRarmJLdHGRc6zrATWCFg
nU3o6j0fGHZdDNffe0TpM3HR4KtxzAEYoGi61/SpA/jDFzskMuXGDFiNCE1tdir7
8CmboZ1NBWYtfuzUoqgWgUOeXVuxAEih02Q34N6S7HMmT+51nX+ECH9JDCFwmIia
UaCLXVAsFN/6jzmAtt/7xxa5ulNglavrY9Vi8Gz2OOHH6AQ1TYtFmRbGWMIlfRaK
uPoLcVfqFy0rzUYGQUI3mjRZbIeSDUYWbm0/oLn5MUuakfpiVYTWvPtbMnTbNP+6
G6BPv99+xoeUf8Alhr3dWGQJvsPQ+LnM+jD+8pzrD1VgbA8fHbwH6XsjerS46ArR
RejEq4R3uRtGYU9ddWxD3ZbakI1raLCbA3IQS+owFhD09ptK21cdEa8hGjIZ7RTV
+qpBzhyqc30OPYoxpHwbkBWatciQoh9sNTgOio9vR0arfvHiibRCV7xxipiUjeAt
0glsDuWqMPCDSpM1d1Mj/XXxvqife0mXNSdXCh06gFg4FxhevgDzRhH93/F/Uryv
ZJj4JoMGDRZVzIVDXwsUMo4mlgbadJY3BubImMGgyboT2RKpXUcrXGaQJdO+GDIM
EUmd3sCUrEcW8IM+ckUW/jGNkzjQXfqlYIEWDfMgSwosEHONFZOewcXT7l8mWpB/
qMlrcTPBNV7f+Z0W65FFnGLJgI90P28A5urc0W6jih9T49He8NB4TTuu94F0KbiE
liB6jPyau+GtbLfad/hFM6phe6ElgcM2CmiUbcQcdZ3zkzjsovuE9z/4uXsa1GTT
+4lf1RP7GX/Adny9w9Ula/KXtGLS6c/i8YPnCUYBT/zorZbEmRgOW1ZovVK068cc
5NnfWTxfyvo4SSjHBkJVnIu6TWHxia8Pq/bwGhEro6Jp+1HzFtMb+Ysg0EZiB0jg
11+jA8tabq++bvKkQlxilSS5Xno2p98Z3vZ0dnFXankxNZuw/khYvop/3e4i6Pa6
aK0vWlFNlRIi56SXfnUZ8uwiZqYdwAD3ghruy/ArUB8lo7rOCUbX4yY4XLRBQaJp
jAz+NTK0XULqbg4+sJ/ebYN7LlM9byu3fNQtMFbkCEiWyNcwcp2I1We5uzp2zQ/9
2KPY6ZxTgrEtCjmJ19eshGQVE2povM9+9oxf3vtTmq8T6VyEhWr5E3cfW+hEbA7h
4JfuTC3wP3YTfC5ovvy4UcD7NdU4hBs67jzzsQzdforMlgbYN8Sl5VWjax8IFb+P
dbjYJDGGjsxfXN1l0qmb38i3glzm4btbfJwRfrsDgwvj5ApERKVjEnqSLCLhJv+g
1M9jNT9cFFhyT65Mrkao6QjPk+Vewa1qjh4/LXjtvwK5RadFaQCol479FDBsovbE
t+imUOWvAARP4TwzifVD5GufgQVysE1CgS/My6iKuyInOuSqugKop7lo6ZNPh8wV
wwOmb4WxEMPN5J4CkK4Lf04pBLBVx9n7fgMl7FtmZnBPoT/AIlQf4CbjQgpwSv1O
mFD5tVikWt4hZZw7KKtTL68DQPaixbl0KQ6PiMtPU1TuNk+BAK1nOwkoZWNfOqPV
qW0roPQh8CK1OG9uOEydoJpINIdfYqUbeAKrXHtgoMAViavvXfWSvoMMDM75ksQV
RQ67eg8RQyztbKumrzE9CxQK/94tFEJ580pC6rvSFQBeCw9Li5/G39PWRh1MOv4V
NDahY2N02JC24nw5mz5DmiPe/eciMFXN/z7i0ApmjQqiv0h2YyvAGWcb1QH3svK4
lqlgqWsdbxGi3+nYxi1FMlep4VVTMrenYBQ4OpXcFj1gyFs4oR/lk+NbnkruTXwj
ZspzxUtPwiV5M0bqd7PGbS/6kdvRkBdgW+NMKuLjW6Xy4WVH7l+cb8GV7ZftePOZ
+0d0wHYl61fOcFxF/xeoy5PC/0Ek9IKAAoLrYgx31vik2e22Yw7SuumwqbI+JQ7h
vqN3W1Oi/jQkZAb8ha+deoDA2AzyaqK9LAHNtwTdAvcohBycNNumpj7KWnaL2J3A
uN0HbVyoVVlp+wwxJqSOr4K3soIpIUXerO/7zhstMm6QNh1pCmaq/XuV/x6wrDaM
oiDD+YjsN4v3bsxI1cKuhIbRRyT6CaUnL5GS1HqQQE8V/pw5bzAqSRBlPck4aUI3
NSM+tiFWWX9tdPUzaW+ws1hp6TA/SvucNooMDC82BWMlYfjPiQUNS6kCNO6aZ/Ll
PYFLl57FnxeELjnL0l68mfkXz7DxOSu9YBn4AQ/foEFlkn8bbitCzoStPtHKm9WV
hSGArrwTKZYyIVFieqmTD4EDEF6rJ/nD9KPn9eo6JXmMYG99l4RVStSWg80iB3Zt
BhBCBE1LS6qC6QRVD75t8wRBoEbGsI3+BmiN8ViU68d1S8SBlg5UqiO8WfUNkWme
oiiCqMYzmGs1CNLnEo1k+7OtFPBt0TiNG9+SDv/Rm9BuTDn0xsGxkCflcuLlrHVX
aM4Vinu0jLhtpSiQ2+nz9yfLIG8ZJwrJN9x0kvmQ6jOQIo/k5qkzqIfuwy0vSzUU
xX2mKwTb2payQQ6t9sL/QZAtnUjqelQ3cjt44Gwj8aS0pjJWXQN1YUk3ZLe6muLv
J0jl4NBmolxNPDkFMyh+igy4S4hTr7HB9NXwHD9BEjZxbkQK5So2CjLbITW2oZT8
PmmA0wUQGkkrvlxMBfGkYsiZ5CQmTNABrrFQ8Zotnh/d39O5l1M21R1/Oiw0PhWF
H2JAXSMl1V6Eu4qy1ymYm7UKzIAHoBFgfSCCCvBS4cD/iw8HSp9wsCp9lTlRK8OF
NKBCMNYHsU6S4CLZLxScIMW8Q4kTOEccyYVbwk3emIEg97vYLo+5UlnaNeAtnguz
VAb0kiT3hPahdEiIHACq+BZ8l2RRemPtvqdKGYLob9f+moTfSlCx3mJViDyWmYdV
x9lwE6vifIzXPX5NIe7WcxPzoIVaPEPlYa4Z/rxncS9su8APKsR8wcM1ekrFn/BR
gxfYTCNiiFsJjIJ3ZSYCu2BXpQPs46kXRVndG5Bxk6Kj3oTYDt6dPV/g54H0OpcZ
yJJdSyhQTILOINPbsRfv3QvYq9n+qB19i6YB2CkwewtsmaYdmNuEsDCUtrkRNucQ
+wEsvbdY0EpCT6YSB14+refmmfAmgoakWxgKtXQ4jhwt7V8wCrR7sbSPiBpVe1J0
wD5AB351/ZjWO/kgfu+3FhN5DAVreweIyHv/FwNvQMgzjQp+r4hKncmyav0/hZdZ
OsAfhhw6EJhPWIrHShfUg9jat0qMQ3Vbj4uqEmY/+0jO2sv+HPTsZMYIGYEW/KFE
NT7D3LujqocP56ercCE99BwR5xFMeSvml0ZmmdwLUJNfmEhdL2xjDGuMJmVFibKz
19f+bppWQ6k5xZbSGje+J29q8oiIblRrcCoWekTTg8Belfgi1XdSseFg7UqnbHmy
bICfgw8Ka36jG6lELklW7B3qOJvg5vpAIzrZ2DjDXMwYKbTNynqxJNw6G0dBIDgI
NCvA3LAdNFdW8wtapJW4kuKhOP1eVz8h4+Of8qEf8TtWEDZ2luwvRWhwDzkjPRD4
4rDCw/Mm6eC8b6jrHoL1cpCokngapBeF0U/H+kmh4oAjfm5KYp1J74//5uHzao41
Y6RsBhVOX2ZcQB67EG//8XzJ0FDvHTuvk2Zld7soDcfoNFUymYivJlfo6Vc8BoZx
xTzPMrnuBGTJjC4F0ta0ZuOnbrgZZRxwKASqAWiQJPjfrnRiN2pN7f5vWPB5AJsh
MaLlaCMauI6yd1oUqkgkn35Cy7Lk0ccdTqlGgwk3X2nTUT6HxbVLc0WdC0UjAkdB
S7cQWxgSmZD/3uD5A7smRzPZ+YnNBMVK/PUgu6dNiNodfQUHqilV3aKRWEB4cI6Y
/ajeCDZUs2DfHRD11Xm0LipKQUAVmALqG3eMK0DvzBuMYE5+a0iknod9IfW1/ieo
qxa31KVrP+Dd4FMPAE2WduvTsfA4ERhdRNKJmidPhb4RRuMi7E4vqJ2V4ICzSIW6
9qI600v25IuTJ+4RJMiT1bi4bkUElmlvjeILp2yVePhIf6Kz+PAAjVLoI8GbAaEa
azHV5aNAPO3HerDaIsGSyMbCY37FdCyts/hVbkm5wapeLmoRDR+4tL5QBL1SiFms
n9Lvq4lt30f8CptSfX9kjfLsDqMDIfDiTF9G/vx+1mok4WN9w/wXXYgzeYC1zQ0d
LxMjH208B22ybRZgKln5Roy4s80gs4pv0/KuI8omMTI0RcQt5SE5H60zQW+qLxbE
5ADTuOvl7P1Ps+eS16M92AySv9kHAdGuU6cvp87j5oN8Q2DewcV5c3Nt4J1M2Qkr
vSjJ5oF11bLysnDPOqwOvzTQZ10Cgkew68r7MdCfHdpGzQfZuBmgtOvaFkP/kflC
ZVCJ8toaKaZgfuLHsC6IuMoJWKTnRZl0UeA9Q1UtgcfYkvrg2PTdwNiTZyIIfIAM
c47HrKdCKsubMnu3nqT7PN+c6ZzuYENNu1cj8szxc0/Puai2gViHS8jMpkuaN4dx
Vo6trfZd9OLTiJ34Dtap5jh3IkDbm7YHUC426Fwip3g0QnuOSDH6jWvZ0UmlYahv
HiwimwHftdnSceBDl5eqTH84HMTEQrRjsgA4acO8WS51P1cEnlE8vFlU3lw3KwQR
KA+LuNY7YP1bfNMCFnkhJ8Uw6ptWDQX+MF4gqhTeXXdng7BDvpppggBmJeNy5d4q
S8StZCZzvgzjWCe5fhGC8GgvsgHo0s3fG6bWHfmv3ncIcPomTQtGO7aeGqr+X/mW
j04HaNMGoETlJ5zWsdyVlx+mkHYgfeMJ9FUQhqh3QoKvwO/w2tBCYjG5thK+9DmP
xee9ZG1IeW+ZnIRGG7uK0wdEFj4sPrXnWyybt6QiHndJb5z2QugAR6X6phHwBYsj
nIKzjISkEQ4r3hG6sExfqsnPEOLQjdRG48/EQVpaDY31QINC42tazI8oKnEkZnMP
H88WjYlvQzLcs+t/P8hLW0j+24AxDDObuWWZLUDFJdjgYKvxS2jzBLCVFCd0vyVn
iq0BmtBEPVjw5U+MNQxf8p4VNg3/AqO5tXqlusl5QTgr4Gd0bWKBffO0RJyEGssd
TwL8W7ac9SraaQVJ9xtIY2ixbMX3CwDWkgvlHOXwTnVCKjG7rU/Z5PLPjSJX6zBC
ScGozZZHDfldYFAN3CZ32ZZoKs73UR5d728Vngj75ZKjrB30NHIpTftAsIrpRess
QYx2AW/1RbPykivIN4d/RpsUK5FDi4Q0FyaRKtybEFGYoVCXiul/mX7Q9WZ8XcZQ
HeU/WUYoJOG/rMMGXAOJ3aOT0xEJe2r2R2B3wOFa9KcKcwiklW9h2xGpZ+x6y+ij
Ej+syHDf6UNP0VuvBJAVH+pcXjO+1eEdu9zMMU7kY+TXULbtV1VFVI/ouMC9Pd8N
7R+4wJbDRDkc0NsEhnFAxM8h8JJLTxCP2vm+x/b8xzoTr0wiC152chihw5jWoJGO
w2L1JswsrAziQF0gQTTxrI4hcjNURnG3IZ9iRBJvOpgCd0sAWSLFQ0rlnfB4ZOV6
OHCW1ERSgcpYdT6WwYjwKx26fvKjaOcdwJD7Uj8HVOxmmQJ33yefVnX/5RaMFfxp
vjEC18jn+I5HL2DcCfIZMVKs3Tzx+dXJNn4rtHEMatTtKECb4DqoIockoD/di6ZC
jpDKvLMbd1cgN0Q53pnfHV9oNGhyC7mYK2VtJdNHrijRdfdWmH8MUeWCFqxxoHtp
91HSdWWmzDriE3ARwOlVNH/g1Fhr71B/v/Grki4cs2IkisZ6iKRrF5zLrHu9DZEW
HmOpw8MgBNBqR7cwy2rUiwMy32e8yQ/evO/1ndhRd9RtsM0Z6gFdIkxcx0HUbgDS
jBm4PnPpOhwLWHp1vjmbrTNFMl2t/5Pl/qjCpNnPXi/a0QRXcWmoo3T+t1jzE1tE
f5diDS5ZDuprFuRd7n+mS2NuQF9yuM42O6N1G0UGjWAqjVOmrNIju2dnLskEVfhc
P+oxXfvQlUUlpUGmj5B9jskdwMvnhSzN9aBPE5wCzlIIeH2JIhJUULYGCY7Ljdcy
T3llASWn2k3g5DMmgD1SCQhhSYaIk4HmZTGrDXUuLmAi9z9657l4uKobWAXxKuDx
/8naGvV9fh3v8pCO1IrG5Oj+9emnUrmbUVuznAdPiVbBmJjsNOzM1oyQF+Q6Dqh6
kkkwrK0Qt82jAE0ZKnS3g28mrDIkTP+qYehUVLF4uDkKZz956Trbh/RaPPmcFIRF
iJA5kqdXX9fA7iTCrZXr/XpZnjDm8k06YHbPBQWMDtOVU4iUd50NoRmSq7Hq1wQS
/ev9a+NAr2jkOm1z/YM296am4kwnVp8w8/6EPABajObXaA2McPajja37qSlEScRn
Okds/x6fyIS+02yVzRHr7A+VnqIdahMWW0Ry5O5NfZgigB2G3dbOtABD74cxj7w/
AvoirXHVg2UoIiyp3j1oCe8cYQlJoMwZUmhsDAJVCbxucDRww2RQhLZwRznGEIOA
KOjhjP2MsH91OJTlJcyUeukVpDvuFILlI0MFwppjqydCgPh+1Md7XWLDOGj51TKT
1rS9Xfh7mjgvb6RUREtEBToC/HI4nwkY837FcXNyhXKbygVt7dbW/4A6NhYMX3CJ
Ilfs2QP6hsDvgfWUZDW0cVnPKdzR6h3fgPFlm6OrC2lcNua4K7aoW3SsGKV7x0EA
aW46zfWyQGM2tk9oQ0LbNre8KKlN5iI/bSpYjdeucE+X1fVikmTZflc6Y6hFhRzU
LHw/6zYsv11R8rGZ1eH9cN5iC7SBh5BTjw8wa3ZYvDbykXOmbv9GZbv8rp/YOM23
zaHCUZKMrAqP4SAu4gUeH7XKDuHNn4E82fMG4kBxaRq4D2oxlzcFyyxvZ9eGBymm
2yqoKc6+P7H9XunQMVUkg7ADJ0C5BrhXjL3B6lEun+2LPVuSQLdfoEFSQvagV8r+
RcTt+XFTQBP4K8GLreuM1N0l4hQk6Rutep/SIzjR1nWk1HuVo704Y4W6/UoOrp7i
5UVa/fEfI9zfcn8r/taICGDSgKgelQ6vz7oQ/VTfUfJrWLHVUafQ4uLn+l96pdiH
rAWufr6WaShpH6qXyZUxsS/Hsjg49qP0iGG7THxKdUM1XnYa+zVLu7kAjGaRk8kL
sGbg6iKVDrdjwwDRM2Ncpg0GEUjceKvHmzPRDjIHE9nwXtuQTcrNR8gtToA5gzHY
AtEZoX2IMxKGgrqxoHxuciyf8dRlTqn/WBV/3c7DJyNdqLyue0xEd6wDS/mtG20t
raDyYH3QOZOG+lFBXjBo/schWn0VNKGT7p1GE9ZZ9BsAPOXbQ6OY/NpX+UIqKqMJ
qUhik5YWBBy7igogE+JfPDghhaXf1jZ/CdvHT1LOTzBWoQB+TuqqfYpWQxFy+8FB
kOLftdelykqQSdhqSrMLVPiAMQnJ81/u46o3C0BFaIfy6698+14ChMWuuKI5J8+J
my1J0sMfmRq9MxkE3XBQabHrn50IRoDAYk0GnHxPuVCTUd4XQySNE5ltNlesmEwJ
yvPkXst7b04FrfEvF707ViV8I4axVS45i1soAXxhJj454IWjiRYCytIf33UkECVG
lcdAbyD2z8cGu8wTZE1QcMwkY1mKeoeqMWo5i7x1yZl0v5khqR8tDow7wbWYBeci
eMB8YSEZkiIEtsOdHsIJE+RqQyeOgB0d6GkJ0uRlh5vpiXNQUFMbFbzjwBG9X7xj
aRrYjzNIfmrzWIhW1i2yYOn2QhhOn6X80TkDNptl7hj22m8LnaU8/xlRUS99zgsL
+NUib2AA8cuoUnWhjtnkhoA6zFAeqIRBJXc2JS1tfe5HpMqYXIgT6n+WXEvN/m28
ns/ZpMj7kij2xKQmG3CXJrnrIaHJ7A70AVY6QiHZRmhQun/e5/Q435ddJX2swWib
U4+SVGAnrHJburJ6gdaeLr8XGmJd6ra+bt7GxulZYeOrZDGDZj1YBTBKRyTKkMPP
8k1qbq7XJW30pY3CgWwt1nYqPXju1zu5d+uExpIDCKKTOc7soDw9yLvA6jrRtbid
cEcSeVarsOUQ5KEdGNDu67v4bg7JNWqZV1a/LbxLipoXbSo+q+Bka7VroSf1N86x
vBgSHz4I/LMHhD20QHYU/0BQPdAlLUxY5YhQrRAGVAgT3RmUbLUu80aN3gnZwiEr
ScZToq6XeKaiMRuAgwPy5RFI9mBPGno2diZSGhSz18dBuFnLwhbK5L8ey5vXnbXt
/Pf6zV34kuzCMiiVxPqeD/vSMt1A7/VyUTIJzHQzpO/tM6abMC436sqXKkI9WUKX
Tunb6qZqAfDOqsWIk/cIir9enYB+f5i1ko85eskrXdHite7u02jaJeAXuwooKKBT
Wi53pasQ0BS7zdhTeUanijKuaN73UOAgRdovU8voKhLcS/y9OYXG+aAk2syDjK1l
14J604xot2QsQtoLm3OpV1IHs122qblXP535Q8NnKeY+YhwFrN5AaEYapRyH/RZQ
SlgwAuHJUQTFmEjcKkLPtZYw30068076lzaz5smAQsgO05/ig7O1tTX1B3n/VNkh
ZoJV1XnzUi/zfDFHHJHMCUmUSkIKOznxiilIkLrbnChHQpW2CW9FlMQsyqJFn6Yn
t/Wrjq2v7gJe0OYE2VueHtjByO8B+0GoVA7eygAkHJK+kHcEVA57fbxlPDXXXXll
ApAKoXoD41CzkivKuFup1rqnwEAeHNpM0dHo34/A4k+yHzzAhsW5mI5xGSjIM3ne
bHXpPIGv0crOEVEClHM2BoLLB9HXVhkQXTrlv1JEXJI4mtYZN3o1eiQG7Ee5XvYB
HYv3C8eRI5KSoXZ+Fv7QGfgVJNumCcsW13N7METl6oR5GkyjVottBzjd0dvgWc7Z
EScp6lFTgFpC9ih9yb99om/avIJmBE+XZ7w7cH1lFGLQbMCO8opJ2IpNsU5aP79H
uhZzmPqA6qRkllCBkKa659bksIiF3NfDr196SOQVOrcjJt+7j5UNMwirkD1/pvjL
8q86gzu0aPDW13Z/TODAw2abnLlC7+2d8LdItK2WBnzBzewEff4JOQqyhkrgw/GO
D3l6pNhw8Gf0nBVEwzUMTP1k25Lorlin1zeWNBecVv51posByB1aB5lnKA3edxb7
5j7zfe80Ymu6KQKQ/NWjzzHUHHwglUsVPvo0TGnkFDCAO4zJ22AavQz+k+mb3qQX
P5YroSPsdxSMjbE1w1H8UP7IC4IoR9hVtoBeinSd4wwcJYkJD9aKugJqoam+EJkP
vqgbJXnxMrOC/y4AxsNQVNpE4rpoZT07WpbR4eqt0JyOy9hCGKgg69LGn3v92lJc
0TW80BQD9+wBDSDaBjyMti4UscICJQ7QGw/fwKzcOSelCE2OyuQPcHlgysI69yGL
Ghio9oPXtr0pVVBNk9ER1n0TkCtndPP95c+f7nvrmSf3filjApJWZ0JJd/pG6Sup
t/fwDzIqm6U5U9vCDm1CrGAKzVZ0Yxjz5sARlvFkjUQCijC/oHY9UCIC+nHEhTao
ZT/CdkwdlBzRQzu4gjmy3xmIQou9+83moVV0KyP+q1ij55wW/hHsqghyj3QaKKRA
s0a1dEOQMbymKAmQBiaZUekcvmNrZDoJm2n3UpWwEEjxevt1Vfk9C/Mb/gsoxOtP
Dcm34zPr/6PKte9vQ94q8TTfaHiJwMfdXdK5ffEsaRPi9Ln+EMIOpilJ5dc6KBT+
1naxm0guQbsPQrSvkjiJEtgRK02dcaQioRt67As6hJV7cR19PUb1RtuRD6xqJCgB
rno34eQeu+l2s+zylmcfrI2qUeIfFUKLbp3u/2hMMWqDW2PSPOhROMymnfeHwerZ
F04lqAiJa4Z+ZtYTI/6FuydLtYU9ntqy/zYKM7XjzHgUUBQZ+Zrz8GC1Z3g2Qkch
gL7xC50dhb+pgK34rWfw+GuqbB+FDecr15LBNRJ1yTCYUC3wMyoLLbX1Mv+GMFE8
jX8dFD9E8005CcPolMCd1qy7uydzn8kNv4tqAh9vNPW6U1kkw5Ia5DO62vCD6J2P
a7jKA5XOzrwvdBtxN7HqAVnYZoqU8kbFYriYwgWk4s9rFTKe9wMXfbPtQUrnuGoJ
2Mdl9Hjyy2zEAaQGGldSE1R5HGHcT+OXc3PIEbRULxFvUYB3/RuD9zDuM8CItV+8
Sh2uriof5ib+EAx0Ot/71agBVSPwMbR3hqVSHHmIvXjGKQ6U8zFmmEQGUN3i8RGc
JwM+ZUPRFQjyLdJKOAz6A5iEcPPdIBLPRNmHCnxYut2CYztArfJDobhyJdiNCIzF
TQ7avEA3amrT5tDR2XghFf0mCG9tkU8W1kN9vCAlNEBkdQEB6L/Eyo3Dp3wwNwOX
LBBCboAdrwWx/e7+cPCO598xDd6OGUTZ33nH1bBkL2rEAifJjTqSQjR683kG0eed
ixpcoCB0tluIiIT6RQzuOin7WogOIblLR7ceGTDrrTXxch+LNqvKPcZJxPExEry9
bRsbkUAQ6YSH//12sfAxhVh74hn/WMdeMMbAC3FbvT1UBb7L0CU0YPHBRCdebWiC
082Vi9qvZU6TqmAob6rzO2mGeSVgpCDP9l7DopvNh1qzPdg0mGkcp1c/ph6K3mMs
BnoNAiOkf0ltg/ul5NN/Y7KsrOCUsyxR+Zboz2E52oRsklcR6NmOS6lRmx55tT/b
FDCwNOgOSHnVWfTAcxMspjV0bCFRkjEY4xpkCn9+90Rf/2dFLcB8InvgGG4pifb2
zF8PvcJs4JtCVVdJVl+q/bLZjO0uqxl53OD4uF98JqEyoTvrHtsyJcDwUk6RwZE3
HBR0ID2d21Atv7TzmF428qYg184yxXVYgCrTnZCr2wDb+LsLr9Aoi8JmBqJr7URG
FnwIzBMWRthkfvcGMu7B77Ln1Hs51Q2zognoZ5Hsp8dxCmtI7+HCtrVGWM2zmfje
DWNRcbFeECw7h9ayav8kVodNXwtCboOjBZyiPYE5y0GmYRzLz5UZRTML3sbdbb6e
QrTwbsx+vyrd5slDiCmh3Tm6rJKSTD0kZ7fa/VGm2lk059rUaznv+863gMm4eZ3B
EOEyAQeR7i+MgyF58b37piTvs5lCrUvhtvK/w/rLmeflTYKla6YEtHoGOTjNVamK
Za10PQAKNULlGfgnv/HXQdYab12UoWTieSl7AeSeUcd4EU2fiFpsPUiJ03N8iIE3
TCYktwiZ/0Rnq5Kzyx64K+Wy358J47U2l9BIGwhKPE+gGgqLe06o2ibtDx36F65v
E9XdNaoeA+6dwP/c7vluLTqYx8VnYA9EHRzWaAtiMy614P4NWMzVBUDulnNelD63
Y02Xj/WQp6kPDgM+pmq0gOhG13b75yfLMG0l+BHn++Xxe3pjLNZqCWKDO0hW+tX2
DdA5kSjuDyjoFKE83+XZ18S4KU4/DTicxfyldgcE7lmiy7+3frb8e60HpTnpZU8a
OtLVb8F5msEoAaJrzGEMURVHM+OSyEHdaAQxBYcSqo7G4sHLFp40UWZo/mAdzGgC
OCC+zqGvcDrOpPLGUor+xXlLi2bLmDsfalN20g0hVIJY1p2gc+kPdeBF2iKIy1Gq
hsbKnOxrkcQ/nO+rfiJohMrpbyNtP65BhBs86aBinhCjAPF6cI7U4u3Ev3JAw9ae
SJ/TOfTEeWVaCKTEemzNO8gEyww31ecqz/4gXpmw6M2mJP9UfE6EcnA9Bxw2kyTI
ztWSOICYI3CvJMHkLOvrgsMFl4cOkSh4uxKnN7SjcaNMfDJzuNM41+ygooVTvkKQ
NJvLwjjiEX8rLCAzJrKgB7JzTsf5kgPOM87g7ZgfjEytlIa1fVmDFagFiPkKlPsP
UVCMHSymp3bnTi6lOlgHsLHDjbdk7Jv7S5IscTC+vVdSFvyC3m9XWX4gNxVj962F
XWaBEqzk7aUuOHLMjsAaRiDKv1JORZNO1OB9zVw2MDirDei4nWLUMB+NmsV/3sIY
+bPS6LLjVY2eHWAktcy6TFPPdVFOq0DZZ47mGnb9Z4vAsTgu2KzSpIltttg+NUlD
40GyCHSO4TYalYsMJfnEitAY3f6gOguVTWEQXlgYr8r4I5++adxA/p/kqn3YxZnh
VVsN15jsegvmdjZS3vPVc0XMFwAqpc8DfadF+z6PsgfR8Lvv0GEXLpSz9XYFl09l
OFJ6Hpl65hm61aPYJsFAUylQtDjVH/YHjpRAlXnAzDTxevC9iZoWqnQ0t6GlxLb/
r0S0XyIY9VFZ9U7lWRrucWJ3SlYq3bpB/UXi65F+jYvXw+I5ArqKyA0yLaG6IhJ/
qnLBqwBp7wcbWMe0A0UXQIgk3I6KiuEYvDr/4puf9T+PZMolz0nTy+WWisimyyYB
jlU+xbhRlrEgvwXdK2v7LcRCnKeEdCZ8AF633nLDbxEgLmUfkvZYzqVZP6m6MQ0F
jLFSEJgxrfBbzfjG4Yn22P54y+LhNssiFSwsv9XZRfg21AFkqpNz3UOxdcOUNwES
SKQ3G/I73URvUigMwMApZPYAGW6Abn8gmyh1Fz/VnSrVpyam4hxQgFUKk/4KS7Xf
RBRbNr85I5C5ne//mIZFyi4oU/++vCcY7h85KZ+nirwe1gfxin+9ximlG7FZ+wg6
S6xksmVrvku6E4mKPkbfwopDIhPk5BUgxeceG/i9M6BDKWTEqTfZGLTggPErrDN7
JuaSBtjKNSBOr301FWQeIuyvdpjOMXJfWmYkxbNPX2uCOBQrDaj0nRgRCqKjqAgh
x6X2wGiQoNQYHAiaLg4x4Sx6iq/SpLnplQzzBMYugqpKnH9Do8rQumky3CAuNLEQ
6lkQMp0zumw613IG3mKIgOkwT1a63hhSFG+KE6o90hZYEnJc3a0dlhNGK3EzkJ6u
rcBs83VwGPqii7+oR0MUFyLwceqbQvxzT3GJf1swwp0b2SVz1IkGCO6WQpdOWXK2
TItSKzKujlHOhg6FnNiye2ndM1cjBySyw8U46p53e22a9aCLnYlXNZWR216ME7wN
dSjsL5rZy57VpqjvqkXYJfuG00RIcz5Rw5Tgzz18M9P/ZH+ovUekvZF6Io0px9BR
OCZAhd2CTByYPwItq8gRW8KOGJwoJ4iZzrO/MnEML/yyEAjwdGT+HOjQRV9UtAms
LscmaZfL7REp4x++UxLP8JAzKLvTOHOadb9GDZWlRRYc0ECCm076AGwrbkr2ZEA8
qSNBOQ6OFGLHm3FS8K4nwCHHEvxF+5iE+10du/tpwh0jnrlLbGCJvvve+hvAIUho
il8lOhR7FP+ufhY1CphhmbwEjt0thJSIAnxx49YRlS2EVnqRochdXbTOqDnLTDaj
7MY25wIaCxMSOl8WvCGqHuedebDkpbmvRS4IyJLbnHos2JJcBEuYMBfsSKyvr2wP
xdML1MRDfmmV/k+4PuKrmwqt6rVxzEn9yBdnjvaPwicAW4lvQr+LjTFC/wf4brtz
xYVtfvbvT5VWPFbTmOQegHTxzBRXhoUwK87C7uh8o/L/gKHwfg4Cqe46mEVx1kDI
wPMIOeIAG1S9WEdOtf+bGBUkji5fU4f8P5s6mFaOwuUPWq4xCERPZRVV15CikVZL
kP0PTYDgKI9e1NKmhgt96i5TMclOmCtgDYF++C0vh4jglWZTKmRy47OUZtRKtR8A
DYAB+aMfyLPmWIJe8dokZeLLCOFKj60o/fQsWdXjP/PT+2lvN00BJMMJdNJwKhNJ
Idy/vU0QixfziT0VcPdb62PuqjVIAAF74Hwzr6SQ20tuqsFuMuEjjwQXZ0wQV/Sh
IoQkBPGD0bMjisXVsAp8NwhsjX6QDu5BTTwTITd6lvPH+C8XrTAfzf+apJXaVPXd
c4wEakPBEJAkJPj2ZU1GgoW/v7pnLnTvIi/otrD9SqCn8SMVQzwPdD4poKYQjZDq
ery1O2X4xmjJAS04a5DrkTWBjGBESV5XadNTcfWBJl6u26caa7DDUHtHkGNNhkyW
JlHGgZAch1vtw+TLEVdwVzaDSflLjGDAhF9Gmu9yFIMV4QeVZSBN5qMqCCE/EAzH
LtLIeEd+Um1heN0LemYi9/GXXKsZJYddI6TW6mVTO0WVclvUXetvsNN18ubBXgWx
FgywFv0qaxtQk/ShxgC0+ei4xLj5g4UySXQ+rtFJM8fcD7X4J+RxjoN1AzvWTiFu
Nq9MJEqij+2mqkl8EKYOjKacH0OL8Bu3JQrRvnf3E4trIpSEOZhaU20UycCpgjit
DI6DcjV6wT9FK7U9dE1VKLNeyGl1x84BWZw5v0mb7vV9SNsHhsNxPP427MFNz85l
mohrbGwUUYNvu74t+L1PbpFXk1Wwo31jDollWvGUS6miJF13E2eQSz7QVPl+7G7V
xd6KjQbon3LBfqD+mOINMLz3+pxYe7LswpPwjXZCngHxyKBxoHQEKXuPGRYIs3oQ
7l7YEeIrPheiSqfWqEu4ByQ2HdJAnrn638/TgJcDOntUnD6xdnFEUD4PEsvj/J5b
sn5n1L4E9SkG0y79KZ3l8XUC2beKrIKctDBpyjVVyzVLuLJ5mLTvuX7CyLvcCGTp
VG51uXM3FYWuMXmuNFiP8ljBn0W4y/x2gltQoAnbXvdORQ6lbfb36XT4bdugxy0f
PCVd9vNQau4P3q7B03hF2aqCPLoBOIT2UISKt+/7KcCQmdpYY8MskRJJhOxuQdBS
8DomQuE6lLTYE1VUzJZbl2oyQM/wg/rviRzyvECViMNOv6FBrd6Ek2DZvLJpiyYP
0ys6gZqgPvkQsjS/uOVoDb6CCCXmOh9npVNyM+Myiz/SNV7aZMDhpawO+bK3dpwJ
cmErU7kecZC/6ZRyke8bLVZPjsv+Apx5pqjLTqkpDrynm3U1kJ/FN9VQZNbLs3Nq
DCFg+219fWJV4hBNnFvKqeSU34+CkGCqbhc0TTH2QdQESU6/BaD2Kh+vYeuG8DwO
SsIQbomfjDnii59ewVgOfSUsMKBs7qdMpqrNaUR+iaElzVo6w6VxRwyXv8fqRhnv
vU3MG/WdR3fFRX3UV85yJpC7BGRCkqrRGUqZoF+n3SBABHXN/ivaE76eo6mlcsmL
d09zdksLiTIYvIDvFgydCHOurI+8zk81xshg+oh7JAWr9JKZv7hkItuIDyLNNQRB
/X1P7I0nqgGG/1rT9x2UHzlRPTgOY0JVtF8JwPRlnpDEFT7E4mYYzqbX5ohtdyVg
9mUWV8UK/6z9BQUc38lw+FrUU1bzvnh3TfgoNJpRN9KeBLci79jK4jbaTMrLW+pO
1G125zqFezp98c0DHeN5O57jBBSsm82bPJJIV8O2/v3+83fPs4QpcgmQ3nf8suuG
asVmJMxLAMCK8adpIHRFNePQN44aUTvbwlO0yU8chxxFJ6MlxU+IEuqOj68+ml08
F5pCmAu7uY62Yz0C3TCkHKW9Q1S8Gu3OrfvIjeOAMocJFZsBhz2hcnKx4DQR0qSA
fgvWklbTyiu9lXMW7tWLFqOgM4cNGvzAxCD2uMhu04jxQd2Wt0VLK3LNlMgeEoTm
D7ArOYuqYnj3Bm/IFjtJQtOAgjcWu0xM0NURXNU5/fBz6paP2Dj/uOJ16hMA5bU5
8N9V7U2n/XuFkYN9D3Lw/Dahn7TFOyBWQ8pnn3IB01zVErqpS/6wO9S9V5yX9+Km
UD2U2VWUtNwatpQqQS7Yr44alYCHxJDQ9E7OcIRNweKJpTBmrHvuzNtP7UuA202x
NYwTHWCHFWT7qPv86y/gPuHYJg4QgJz2i5kaljAR59qW90/qVj2dpr3hi3b++t1x
Zw9aWs9z3l/43qIfx2J9de9XsI8V4oDKiiKNqCUY2poMhEQm1qzX4jSPCmp/4fx+
lhHr4V00yntbqUVbjlpEkeMLwe9wYdX3XhquSrrSeo+RffKSPbSeZc7TpijFNhxN
dlI9I3v7xAWhLKcQAHfZJlbTViUtjmE2AeHzr+AWQss+QTyA+KI2yJ9NBMyqjthv
ImQOxzxPoYSX/MHSIIzhLF1tRheWny696VgiHqKEJtWHxtqHrzbG3Otb0ljctUpo
ddV2wdRXOsbPenxj2VyZqRY00Zl0UOGQzeCq5wWyUeVZNG/lPCAkkhUKPrTj7Oan
mKaIDdnC1CAGsHsTjFCoLiT88E2WlnvUfItioe5zbHIUy+B8wnACcI071jbNNB+h
Sn8PLxDCI76TjSyOtrquLvXPgdrb6ASliJcu9qnfDJbmCexSMcZ0GK650Sq72KaP
bDzSaV3LZ3ZG78gbAUvG26zyZ5W5ObuyDcSVDv1GDPSWGZMZ6mDNaIyYX/F+BhYJ
MqiUEcqY1Raw9o3jZTAjoyib7cgNS5kId0jv5erVr8sGFf5kUpamY7xkc8W7mi9n
/JIIxtjNDELXc3mwUtlyliHtCCg4mbwb6YXlkoGXKe/5X+F7Fjv/qbFo/EOvEEvQ
5penjeW9Dcpp3Rwx6mBAggMOaJrUS8GPcwM4UBnzXNT+bDR/OmCv7sB1KfDVerzs
RrlhsxVGs7594/ttaWYOZjG4zM+x+lwt9XsZB2IHNgN+dBfP85LUKYaZ1H68MChj
bKCo5sybGehEI9jgKx6h8Uij+DXiyWOyYAneMB8iwTUUKiY0UcVxvFyI17sy2Hx+
J0wz4/TOT3X9Pnd3MkpcuFU+JlpQwVNiWELWKLpxQ0aCJT+bjeXoSUJbfJjz+RaL
DHDjxfdB5Mfj0bugb9fxRU4HfTtL6V+8RnujWvGZoDdEAJmtMbJv2x7Pa6HT3ggj
VUWmiLs/GNocQ4nPjqs664L8N1jSDoBcM6domb2L8AZcGvGkjnAen5Cd/DH28UvB
AGodM0T4J8igKzzpGOSdnOtUsW9144RB1kyHhv5a9aoUCu+mUtqLd9nIVkc4eYKg
F7kJ4sudIUh7MCcrhiVt40qMCXKxNyclOhMH5Hz2YGJbqTOgMJVFqw3yeJC1bWWG
M4ON4aDEH3/0uz9lsb1q5/CwFMQ86waJsvnHqLT5YOZYLXuAkSAELXfnuprYU+QI
0GcqGExz6ZijLjE4uWkmzqShGY/91WKnl/7kc8qGf6f8eHRcSm+QVVN4wNNWYHCB
CvvWH2M5MvX9FCYhPt3Yqc0JBaLNAlY57nwqMma5mfKNS01uniRQgY5w931TtfcA
F1QSuG0KqdwhD0tSm491umaXdkaNILEUQjHUw3M0uZI71eizEaD8Ot+RopZvHf4w
1GTb+UPAi7o6BIOX0L3OzMEOyZJsHatuXYExwIosFjRtcNrCNW7dwd9M831DFlk5
CK6fM8RFRj6rQkZg15rLw8yvGUgrwU4W3nwUeIsjCo+RSykbgCj3X76LFi4bnQaW
58Y49K8etnuUbFv1YwLw2b4h1yIqEJc4++xNTGs4SyRIbw1SnVv1AXpk+f7XQGED
BR+gLZXIbnKXAwSeMjDHffUzpjYLF8iaXVcF6ub1pG8+uUTWBZW15cf+vM+HKnGn
WjoNIAdyrrhnFNz5dQGC3xe6/8wimsLi4IapyVle+ST0Hkzl0Ltn9IlwkNCnY6xY
K2uCNCMKoqxweER75LJDyj26XMG5eB0sQrwAoHNCBqqhufp6jKLHAwx3NRTTUfgC
K9XGp1RzXEm1FXwYCoOxakqbdzpR/QIQDX+yikZhsIcXR/MmflHq+CbqbF8Tp7xE
cgWS3fsDYHoR4yq3wZtYRtaJQwkKN+gOw3JAzShJLX/mJzDoQHmuFHN1QTuGrK0w
i9+Bl+BqV6noQyl1sbv0pmCOpt/jzEUA/F/YgGHEivFGttYk3UWiyrc7FV6EoUbm
IDNOHgOF4gqRXd4442C3CTVzCp2S6LGfoSg+JkmNQYPA5afQF3IT1ZetJvqR0oK3
LgxyDazjU5dgvgboVoA/toMhR/g4kBIQoEvjW+CLvYa5RSwTT487VT9iaozRe78H
2sxP9vkCQ3fxfy3ymjHBnM8IFT243kxfX/e+asX3H5TTJN3pMMya4PAz3xkbMW73
nyCghPTrQdYbQzwO+Zp1xcRzwzKyLnKBWybUNdHK/t57Tsp9N0k45j4gd1La6WKG
cXh9XLCtjug39k3+vqNTbZr4TdNBT6Fx3vz3meGF5iGlRSgchAAFAoHoss/oKSPw
expX9YPElQUGEZG3tD/gMLzE+EUulx2AQmHdQWmkbjYgx+RHsPyNA74MP8ILG5xk
ghx6vnwqQVB8oNLrzBwdBvEKLx1T935X9bxAXaXaGjgx4bdSNpzm2pVg54qXhbWY
WY8Gb3B4HT21RdqSIyC00/jywoc3FU++rP3jB3eBB1dy8D3Nrs26rxfKMB0pKRC+
jmy3lZCRjanhgW1JlI4XLnCcoUharAzqffNamCcWbs0NJ1GEcamxvNq3RghyEMhQ
C+tKF95LQTp5YAJdBwYqyLzM+buG/o8piQeTi+UevunrnSbrGbsnWRA+1Th7aEjm
dNmIW4xiDBy0UkFWulF2kwt2Z0zGd9DkC9scf61vc9OKN45JQW6Uo21U03bHHYFk
3ntCfPyigo9zZz99R28A5FcFcDd8GT5Ls2TYEgj5wzErloNeiBWuC2tgwjCv7w+p
DuJwCcaK9Y6fMErChPFa96IQyuikuqiSuH8NemcgPnapCmo+wob+jaLN6GYnm5F1
QgtRKAEXOZIIUNBOHneCcV1jIuxinZLA2sJhSIVP5px03BjJZBh4jp8Rx2jTIgKP
h6Xqe2eu/7ut4kaUV3IS98dmhUKrhhkCjKViegHcKFVk7wjm4sG9EugdcScfTFLN
ymCLB7Fk5HCQrb3/8uFyGr3x3ZJlnUeGHBcullZ2OJZU6IXfZHJkKi2k1UJ0bls6
MfzSXimARJIVaCTO2tfSzw7v37/Rap4l0rGpowYpZ6TRyU/jW1lpjQaFOcDafDB2
W3oDlX8RFMZsTIOBpyKfzDdP0wm8A9SzTlqCXzMwmuPfQM19OMG84J1VSGycqBsx
5ggBTv4lAqww6w9HKpPrnukkk8as8iZeehTMA3Lswv8hmQocBbb565y6/F+lcv2Z
Qz8ksOewoM//tb9SlTlN6i64hW89VUWwiKiHQIGpWTOpdqmyL/VlD4Y4gY+msNc7
Rn5wBcmC/iCyE5GQJyFW94hHKHB42zxewuzky650ZY8taI2/F1hVodo+ZblpXyt5
J0yNmYhc3Fbc15I1IqKMGjmy7OBIHCbp/eHflyQuEi8sM5wjsO9DO+RSEcJGmuXH
Hg6f7b4LFiEAQjCTdKKwEdy6CUW5d7E1SlnZ2lqKN9eZ8yBvUPbq//uL6RGr7ECt
uB4fXImciRhd5VNJiPxiFKiOMhSj6Ai/uEmcBv3w4HavF61kDE1zeldj4WHtnpUK
p3Gi/4mc+7UAylQAXtVyBJqWC+XtDgCFtHiEX9g7sVgNXH+CnYToCf3Ub35+SDb4
Oj4+hziG+msmz7bXGYlTtpna/9rhNnS0CFz+QXweqt5F5Oi0TQowWIsW8r/GasPC
f7kKB3Pw0haQ2MJSeqKug/jzGhFeRCISX6uSYv6PEHyJBgBmkpss6l4FtVnQsjy0
bu5baVfqtiDTOkIyBcBoI3ocsaMgRR8LBz0sq3EcqMztjKjY1Tl0vb/Cm05kMXT3
uX/g7+0tT59XDJbEiiyvI4VOqIr78AeynrwcT4naAB66wKtm+omDxV/D7ZNRrTws
G8XL7gyogkX7yqhO6KXETzJyD6GV93mEDXQUZ7WLt6MTqf+VB+UaYwmI/kJ4vZ16
IZRCIEGo4mho/OEDclLfVQwwRFFm/IBqg/XKukM15pYVed8dSROJUiCXq2nmHHkD
ko3S0R6oqXQlg2Uk8nE2X+fcXlCPM3cTgU8RXWEXf4QQV5eaJAWfVfZcrzDel9u3
4EDXlrIWuxQteWid1Mnj4ykBlYAqPbOnSpaAy9TwGm5/0OTqXr3hvAMsPkUEwide
gwVfdD4AMseEJF9bdvjZ1jjdsoxPIJfsalR5c3yitW4KhFPvaoVqwYhTP3fdYY8A
wA1GkUSUszLPhb0cJzb1wvoWqL7lfIdLNspZ5Vec6UVZiqKStbJBLWL2wHi6aGVf
5/pF4limEPw8zdwYZVexsXMAaOxU6qbUl8WL2f2UPZtAlacXdArDC5aCLpNRaGTb
S0XpYJP73QwKxdn9njbqv9eFYlSLY0g690tC9E4IP0Q04ud9xcVeeRYEQJPHWGDi
jR8k7lFrzOXNowwHCNs6BV2NslB2OEwcKFodIH4DRVSOU4M47ZQMbd2BSvpekdSk
K22cT4uQ38i9KQlLp4SKQ09+kb9GyyrKc7NPhZ0W5diy1C/zpYqQp6jbgq9BJaz5
rYEF/OG78k2DpJpn3hiq1pjxh4gniHcHiweMdLXlkDcv6YBo9kH3aZ3kul7d26tF
qDFntImucdj/nSE0VY7yEFsOIUzrZsP7BqaN1Q0cZdB6s5k9FY0PhTDeiCmBc9BE
Zwg/2PB/3F5yDfmR72KeUWrl/MY5yQxH/bK1f0Aeagdu32zzvmsgZFBu7soLGiKU
XZZZx320V7RJGncVJ2Ub76uV9F4hcGHU9tn/7Hpob9IKEadkfyPzgbXdh6WIWZey
pgcY8SI0pGVPRMYG1BK5eqhReT3FQRRkY+SsetkXtQMOA3tLLMj/HxFDqzlrAhZD
HOpG0O+10JUdDuky9RgWlPBR6uaGfpq2+ORUljv89JiDwIOSyY8x9Xys4+WyODZr
zi6tgoGhVB27SMf1ePmcPRwCPt44/y/k4ilYF6dtD1EjP/i2Vm6Lv9n1qOyqmNhh
UNG4H6EB2wCPmf4yS4raglOTPELVMfPm6aerOrOJ0oW6tRNAisllqOnONPrsnrCe
fDLzLTuUK7GjKCQX2gPBaaZNC3EdnZJ+Gcj8JmZE/Meyw1IwDLnvSuLNcZjExyQM
tZ0ctq5M0fxhqQvuigDy2JMxoOHcDDJy1Ycc5j1xGu6ZeduMDKx6KCDSo98Vv6gk
BGCW1cfhOZP9QcfUaFQyTRFUX26PFWlb6MvjLrBFVJTlA1yXzNe1hN0wAcpQE506
2Wwn9OlvTPALuZ5wrSlouWi6cCI/ZuWh/7U5mIe8VETxlZDHz3a166qsO2VaQ6ns
9DcPlSmn8FZdCACi89fPouTdr761LbdzW9dSHwxaHd6llq4kOHhzWksWwl9If3/9
mTWAS8AzouZsuQola+LystKH4Hj0OMXj1rYeglJJQHLPuR/ETzo4S8ykvW6fVh/s
l0PLKp4ILi8VkpXqH11BoaTtEpnk0jCRqyI96TIJdatshOOyJeksPcJVCNN4+4Cd
UjqFvJkJi4wNyljt2Pj4bboMuMSXnoCk9dVpqndRI0TaLBZxBwUarn4iLOjS5Ioy
4GGVWbCo7kmcWNQNKJVC0wBNFQciYg25vjkJnGWtcXaPHi0k6BAfDPFJlUtm9pHV
mYKi8pbO6z9Ukj+DSA8f180NAn7sBdzImuLwxb94Wot3ppBJAmi5nFdaHdMEsUeO
3Nd6DBpMsa7cCXODUd7MOvtSp0eemGL5gZcjuwJ8Kh6PRAr+s7P4NvhJxv+tswSO
qHLilo93atg/o3Cctig3wpJlTthDLGUaNQ55wMyx8D2wCwCxAdufbWzyzAS+sRWl
xPfYOsxeZLiiDme0TI+F8FT2BDdVx6eWM15pJiNKgL8XaYT4wGTt9MK5s4dMQLcp
R5rO+JSkSLzq5gr51Yc8TBSPawqVxxty0rAmDhrmyNUYaB6l7lseih6MYsO/fqld
3Bv/QZbWPJzvInHS6rYRTNgYO6YQIVasbyAOaihbVVjCo6zNVl1M35KJUuu3yf4V
pHW5N4tExhMNHIlaJD6UZAsGxZiBa/+3fwoEVlBjeBwHZkSXLcdk4a36Uwsaeg1/
w2QIoZnY65ppFpu4/agw/MBR23BRh9esY8a3Vv9sJu1UeeST0/Hofi3FZMNSym8V
ClKQISiQgLnhwPCbhDMk0s6gvAmKwc2FpQUWn1+OqnDZEZqDr9mL65KS/EhSc02g
nksjuek9C9Mh0j5UBLkMlKWNDLpxWbClMPQLX1/I3SBc8vzBNUor9w+g2A7MCaPl
N8rRtZCHYlu+OEWgB3RHlZFqAOelneHWMQiR0iVN+4c/0eHAp8OXiqCgjXMI8SU7
6kOkwE4dKYnHLGqTF+XXhcfl4Cfi76NvI/Nx9tX1eRsusU818wlkB4S9Bq8qHqMa
/Mwb4X7G7SFEZHR/CxX8h5md+K1WzBlDnG+FcUgnGBraD9byBLGOW4gm0OWGBg53
YM/2T019s2myIUiSNbzbnE9UCspc40sv8ModUqS5Zx6SUgOgvtdNUAT/aK1A9NnH
2ViQ8GrNlzHbolcOYg7A4k0aypggPeiLoOt7QMdD01Z9/AO2oBdUFCGqcKF32/cL
GwcdvdyWPDI258wMycIRveM5H4WOqwFouP3cUiJeNBtc0oTQ71jKZY259FNTb0X+
INdj0QyDdNPDT8NEGiXchSyXJmh0yEMEXP3ZraRXDDf65eAIXJh5LfXNZteZWGvg
VdS8e92g+mIJVL4XmtUnahjce5qf4GrG/RGc+rovrDsK2UNvZYbI/E4o1ZyOxjOW
MGrRnvfpiQLli6Q82J/OSVVZ9CZjMeraCV7GZ+n5HywKmwCDm3JmjnaRsTrxunvg
hG9O018dpJlfKzS9/6G7gk5oWTn+oOFuHmh131MZRKR7kWI2UA27rc4cJQ2w8wb3
DlHSxPKz7KehR51vJwLr4AyDnIFH83epb2uRJTRiPJn/889Xg2kGprTmGdJIk8Bf
VOGo+yJA1VgAGl+XyP6GCq2eEklor2kFmkqW4giOu37dUOfhvi7cT6dHwtjgWuMs
KrVyRKs/WV+kY1ujA+YO3tgx6rTPGZ6dJiA5FZ1/SAwiRcV2pShom3pq8DTCMyWx
sBdB2mXltIqhPLh97wH/PQc12vy3k1jAT/u34P4p402K22bCIPWjVH8y0WVeiLhF
Ftmkjs88Od2BM3c2mV9WvpdQIntrtT70YysyIDiUak+fGmM/MuhBQG9CJM69p8Pa
A1rlNrbFvMPOVDvRZ6jerxycFUQPM2t+vHaAMaJnyCQLIck+arPdYU1mjY5XDqtA
WUe6JOKUYGIJRb3KizB+0bUcGlvQa4De7k/DZl3k8uV+8PtzHBeiYanAhx6UGvTm
39mM9fnBNdMI4QK7VKJpyVq3tjnsGV2kHlVIkVq3nuojClcyCeVTzaf4moODWwuV
8bz8BmoiVPsR2bvp0M1+yzdtPjQMan4xTMlagOpM572OaonDDR3keyQN1xqP+uD+
pXcluHslHD9jweFYsAkHAoWKTOl+BYBb5twJeE4Goprooc7hd5NDy2DJGDN0bFf1
hEJbAxW5O95nF8tAtgN+mB+7HXfiMziZRRDXNIfcAPhk5qq0S2q65KFAVdjzsm2a
zWb2w++pNH32krIRH7qUpFUl0n6BFGwxDwEoVfcKVUG95q9M3pq+6weak0u6/GQx
IySPEAU3OzMzJ+ynLsxP1JWHZmWZYngllxEOJkcUWDzWNz6wmDZ9ayNBfIzZL9WC
udulYWthOzc+ea8a+17vhg8GxEJQb4qsrvRkOlxLJX4PMYil8x7wB6S1FgY7Mayf
e7ZTZlXrDwPYze1SpuNIW4S/SwvBETL0E+zqpYFFOpsvQNUiOZytZ1zjAjiiy84i
b52p60n0MlrGXurb2k0eF+fJiGa1RpJfE3kPlccL1y1zFLp4sPUQW7AR7WULRAEV
w9+ckDYY+XTwCQLidbVSrOseiM71BCxRtqL5YXSUEg720dI1NQNwMyxS19qZ66cr
HAc8836Ui9gCXALRubQL1wFMrF/QWV5ZiHR17M+1jRKFrCU0UMdyydgGrhdSL6qr
y4Qsrxu1mp/Mvm7YPO0lF9IXJ9Vq7FvymkPyQe9/3csgWJrg7f/qdMR6Vz7XWuKV
c+GRaTbl6fl1ztTL+rGA3sX3X2hEZuNdMamkd6KVTHcV1GTD++5mpp43wxeTC/zc
pTjD60OZh0kYXaZe4W+3fw8Cwt9iIlDLHTIehC3E43hvMsrey8dTr16NXHPnp2ID
l+s1f8oyJjEIv6QlM9fD/W1Y1nb0IfNC7aT9QvO3bf7KARooITiGFRVopqERqfTq
NbI9BZV4emXNYKb3h/xU1fUkIinOjRvayN+OMl0qs5H0qN1dzL44VJVC6KPzlcui
pqQYG5wNkYYPWCGs0nwXliLz69xZ153rpYL35Mygmmj7lTl3Ez1nOoGsZ7WaOP4G
wUbeu2r+wMqLQ0yvee0p6oPw7YtSBrO1FCS9OSQcz3W8yKvmbQt4eqb5GsoC2OOK
9DIZKRGtmgoEARGBcjDuRL3AqiDodrNHz+xMN+RV9mTdDpGvF8AhiQ7lFWZUL2oC
erR1Y2KGoWTmiu6JiJyPm8oe2KyPRTLJ/fKUIeGQuc/NbiF4CnZA6dyLE1bkGIll
qVfSIaYRUhqSPz+IqodzWnM2ZNNLPjWZWWbnu2FGKVimwcv2Ozl3EfSoYdM6dUXw
z64Tr+lqsjB5KkXZvpk07jnLIpDtDErZFSMIfQcFGXL16LmYqxiPVTN1GWv6+7i8
Y/OkUH7ICwhVaURIgQ1vGz0dUcHYi5zJmQlvPb/muzsbNNdfSiJBozbHFpfdubjC
3Rr3P0rGcZH1nh4kNNDUtGWN290xE5UgNHt+jw7LCdvoBkA6KEheNGSrihB2CACK
gSo/AqSNbSR1OQbftrjUKmokbuBsJEFMi/+401wmDIibTiBv8NYvCcYh2OZcdHBX
XRVMFF/g2VQyn0J+U0+X5F7YuO8CW5HciUx/3Szxn0QKSwrSEgBLLENUOTB9acOP
iidoQ+LX+7GJcgAQBc1gpRKROo1MT0jRLwXfV/RbiaiFdwBdZ1lmk3spa4IxFLFc
0/ym0DFuf1qtLRlNsODky9Xc3N+z55e9jQrZZHIk/IR4g2m9nNnndYs5wNWRIZxS
a5GLFu+nexIGNWhtqVdV7kkpOdWiOL27p2Hq0XlzBEcVK/uiNjHDkyD4IJHljeZ9
5zRYpK18cEDj+UoSsr8CDHUyeoKjzK3JSsuOFQ6djoH2tOi9x1TEW3i6VbGMmMZe
eETLv6jI4nOUBIsGy01m77Kws5JlLjrVEt7EoYhK3wOZD1j3j2W/xnyayeh0Y4rW
eNT9iw2hvTda1Gir1EQOqnd8dBJHXZf8uxo1Zq38vcRkzGPGB5RxU5pAVmuWq86G
Phx9DlQvOkgQxQZWHTOj+m9OyM6qyhahdN/lbtpyiER2DDe0spaXtXj6MC51MpVc
Yp7xTXYzfNZIsnPuUk7C+QvGCYqeYYfqm7bsjRv4nwtiz1oCEupqb2mAzoIMeuLa
erAmPL9V8IR2S8FupZnmcg/eIkQ7SLe+s8iOzawi3AKtfX43W2SFhwfrBcxtT54D
LxYkct0BISadprRPgY4XUF5nYiH7zcgyXyk/YJA7Dutx0boajGk+mwjs2tmp+CqH
sV6Q5o91tlMuWKLjjwV20EscUc7IGddU0Wkb81KI9Y8ETF2pUlbowUdaX1opYYFb
G0BGqddA9RvTR0EEDT62jPv1sGHW7xuGtPkwvMNH79g29JGaoAnkQZVOl6PS6dy8
4C4/H2GFCuZUR1N1t5m3bBueR5cbFwtX7DEE3dJxkjixOzo90brodDvpW4Bw6s3a
saQnXraLfy3a/ntNClLS3NN/x0tPTnXV6UrlTSlUEdVGT0Yz6Y5n/T7Dsn3PUDnr
z0K42p2n5Q/3YkKiOlDNcc6aC71mHKOIlBzQhDl02xzFPTNaFPpAtQNqIhteFcU0
4kVOQdNqeA0JnUYinmY7jfd49Qg0slHVIYlTkvJYX+xGFKbvupdyef6usZoiLlMp
ofKE1zWmsyY2G0sjoUHv0VPg38UCVneB0QJd1G2IQwH+lPhtcnjFV+ynJFDqpuWS
Hw+82BEK9ZzThMYLY3GbPh7/K/w/RuztCMmhMQj484GiRRpD1ELmEKG2c9/fgS4h
b8maMHUd95wDu1F9F3xuDpwN6A2wFjcoGdRDLjojztBBm3pMcs5+DBFA94XjEfOW
iJkcKZ/AEr43SOoRTSj+XJ076wNuQm0Y2ZpDFbdCPL98DMsslzOpMl/AvAFUPjhd
ia3x15E3aFNCuHGcAMoPINXKiQ6Nd8hAJ3qrHu2r0roK19IJWumg2ftEF0cnz/J8
2JeR+3rvweN6SaUJP4RL+lVq/Jn9lVyERX6vmowB7VZQrAxULoWd6RLwdiRWwcpY
+YUgWaNESihgeAafy/lKoR6rYBXfSFDAQV05kxbz9ExqT73m+Zo5ZhPN8LYLA7iW
AP1yY08FQ7eBoufWF3je2fwAdNTI6PlqpGACZXvIqx3+MVTpCRVY8rTt849ge/IN
SuByMNxReg1KKFHEmQJlVnNGF4AENe/D4dPBOJ/aIH4vQjTLucJNpqOcLuxRhErr
Ti1XsRZY5gofj0BO8PrID4lCE8MrFnQAwXU3nIk8QRa213oOEuv/A9a8E5UTYrjs
N++X4jR/kVUYMNbXsMvs9GmJrCUo5HMXXbwL+qP67YViKnPO4YmkVn9h3/w889cx
an8OKaPc27JS66Bpu8YLuayUwG1tKeKM/9npjIoiQqb/uH8QDp1oSpw6SFSxgM8/
09uPrYfQHXdGawbDzFUbOnsyVJ45uAf1gtEU8TrL+2bro3G5Q4G/pVIZ+l13zy1F
dVznZx5PLtsrcdJef5EvmDagyttioR7/M2Fn9yQoXeQXk8i0UBnBmxqbFPHLxiMp
bLumxrj23BC4ZaKRPDmf6fGO6rwFjGDoWWx39KSLvxX0W9HCQhIbZHaDuLSlogDe
KrgzCAm3m+d9dba/UkoNEYa/G/wLVzlDT9f6Ojp5cELJzI6XMo6oh6MqQKyk8q03
3CgSI92gcN19SisYQ7x2Vl02X7nD92hkcwOqXvtn9dpXF4gvWJPjfPYLTL45NRfu
XZK+I/thZAmKvMDyrQLmUXFErFoivq3doMANdaGkMSFxKgRwaBo4yojSKdKYu5wP
Z0Hw4pYmFtkjFIyZgSwz9NdMluMr2JwPn/2GVOJy2FiGOixFB2rV/PDdbHRh8/w5
QlJ04q0QRo1WDIs0bRpjOG4eRle9iGyvgPNbImdVy+ij56jggu3wsagJScTXzCuC
XKSJNeXHs849LP+0HaD1i8K1BewCTeQbtRVJj6OAChnyjkMdqNNct6io+gMsZZED
6opwA8x9IrI4rDqHpDjnjwCnnHB7oazNLhxcp9QDCPkfj1GdxAVMn3kjr2wtOtiZ
f2T2g+sYxXa6fhUEKt8tSeq7y4PcyaYZw1HgwtJHFQfY5QL6TQQCb6LnMwp1fMt/
g99Hks77KjDRgTIBePS4hxuer0mp4cVYgXAzLAf9Kva36VXynlQtgDtQQESb+xI0
wMm57m5rNtG7ZLSzPb4HczXMSdsqT0riZL8VW78G6edLatQJeO5aQgUUVt+Uq4Fj
piPftyehH9pRIppWEqN/GDrjq9x2KnmrqEVZxGj8YuKcfe9kJFod7yhtcXtdLEk2
Dw70IPNLrQ2kVTUFXZ9SKJ1ltctCpj+2tNCGQYIaRwC/kgyBC3oq3TwGPC1D4xKK
+hPELTppS/VugPn47+m8HWq7Miw8f/oekLYTdhHB/QGSU0dCmq33F7HUbV6N56FT
ROe7trV8do8eFlk3KpWFeOXP/wDjDLP80z23LIbqNQ4odbu4QDAjDyTG7tualS5h
IYbJGv8pJeHIjYYmKlFoU4SGYXRusMx/Dzq/d6DQdwoEivVpCzn3/ZrZuR6Pq3sD
oDrGC2SpH8aBBp7aichRl+Bd8uwuWD/cQBgJVIcUd3yknJrpC7u8XKq4uR8dl8Nt
XcECh09CVGLDcEzlQFj7rcm9v5C3WmMcv0Isan+ZEFpvk71wy8+TyaKLaZCidvuY
CM1pz/sa0IY579081KWzZ4/nuTI6Smj+4uE7g3wp8IVcGrSZKbSeekLUVHEUf5cB
e2h8X64lIQZ250FVAye6Sop2qC4oSIoubPDE9Bmi1WOhn+DJlMp8xAWpfYVQS/II
/vCVq9MJN269tNIxtmVNfHTDjZRgztNipABCX8J7q61W3mVmEamvcFiOd8GOjU7z
qgg4VFlvIhcjf+guoPSDIZ0WbU3WJ7rXwIyRr9JtSmmCDAxSSJRmIFfcNYMGh2Z5
4g2LevjtLl9wV3Ust1yN0H1KNv2t5Z3qY8T0NTdrZHbam3lbOUHjtDxyxeBTzxCk
3Bh1YVDbwY/C8ZbDTpJBI/uOTdvmX/5dk49goYf/YrggrzO1A3p6lOZsr9c+Lfxy
8EgZN4dtjf70UX/ijLfnyCBRwPKLEPbQkZDd7OTKv+VQ4TS3NXzbje/2fAckmi2f
wX9CHByMRU5RzRn4r9dq4fI56wb53l/Mvxl5PDq0NqcCjQoyhFuOhBrHAluRwNIe
k1QoyDHh7cVaH8uXO6fkUO5k+V0cIXxsVIzaZ1uiNqoAn5eS+9V2ngALt6dLmiiR
wMJPEFQvXe547Zg+Qx34UlAOkCJHw6HGPzLsNcmpMhsRmvSpznNk3nhebk75/sp6
yOmIxSOsVWl7nQ6lUt/UMWIkyuYVao5NPfElSmxtobgOAKJuYZhN94Wh4f72KB61
d53fC9i0IWWSKHZ32Acqg7bYsNzeRLVorKhOV+238QCojvFxktqDCiPWU0XIGYuP
1MuCw3at+QlGRzR3o6pc5w95ODxm5pJVczYumzaLzr1EeksLSh/pbVRCTzlyh6NX
vpUuK4anCPUGo0rjJjnEf3jKkk4AXkmj+A5dEv3ToNovknpjHY7W85WmimPkJhj6
4sTTqLxc2nD1BwCp0j0Fkw7d5CLwd4FxhTqp7HJdypYnx78sIKGDisDRXFPQ11s2
wRkYW0kQvYJEmbkJd7aI6E2rT4qJnfXfH660bRPEBL3+hM3WLZ4NXULlkk4dBt1F
EOYmukcJ5cry+skqN22yc45utlyR3ayTJ1ue4u44vzElSEWAFMO3zKWPbTUNssRY
4dquSEhfQoxDiqxUOlckSaUUpJSGy6G/Hhk0F4Bq7oXPWsgwBq7/YkC98kshRpBr
IMWRFPKCIxBWBFIuyWJPX5CDBIJyS6/BQ7VqaHHnnsDdHHS9V630FEwTxfI7DplM
pVvuKdMYj5Hj2jW/57obuo3pP3pHJczUIGNiFthMZ2RcQaAPOEF2qlqlN2l/ARa0
sRBNLyVQLBw2BGX5VneLMkbLTbvwj4/I8VYvIZWptJy3EfhQcTHS/qrUVfR9Xy5q
r8jPNzeklNnBmFphCucfnMfFZGA0SmjDynF0oDMng1GwH0957BtY0bW6dDKDo940
/5QXCITnKB80FdYEcbSqrMymGqmL1E0Y8SZMVPhrt1kymAJzMc8O/euEr3iBsuOg
+xq2G27OiqIetP3l92vmdMVW/CbK0xP1cLsaknS+H/c9u20pXhVbYtlpOvhjQD6V
bnEo/SetYDsgUsv0IgqYNNqzWPZB3HJScgSFCXnNyHEgwxj1cVmzDPe7OgBeg/q3
uk/gNtEOSjhP79erqWhB9oOEEQ8zYDwuJk+uqfTn2lS6vLHKGQZkATKHWiQeP7/r
JpWh4d/rGr0cNepAxd+euKHmJjgeFhsQy9SoNwqb9kMQgOXATTkkPEIMD/8YPF74
gOjGUHguTVMktf2XHn/RHWL2hIVbJnJsknVdIkRzm+uzT9LkOX53Q5YtpSvN6p4A
ZPVuwHfXjOWX0NWk8Pp+KIwimDqRiLKdSUxXHC10UkZLARKvRlQMvMnWbbFw7Ub/
XKVo/wDat8C0jyaS6MNaXyGqLPFW7hghJ5tUla0aI9sLT6rkM0Nl95fUr+Y0y3Sw
06xRp5XxQLTkzZqesgps6ubgY7u6uiPr+fHvcFhjvlGLcj6nVDlIzV4ESbn8Fnre
6w3XnvJ0pgWEgN8H0ACJSqYKp72rpZJZx9OCmFHpMXeYoz1CiqDzk42zcWGqXUmL
wJ4Am6JVWXSZdBOhRBkJ/48Eav2Ub54/2O2gT5nfB8avvZraItIUr6qiGP7tEZxG
mVIo4294rjKxHgR3Vy8xm/Cv9Z+Ny2LZ60/La/SlaGaAxfWedpnXsVVXsbUVo42w
PY7mL6PfD5BBw97krFuwlENryCMKVrJNTWs2LAfKV7tXnwIaTBQYV/VE29Fvn20K
LdK5WXNqZu+LseXwFBzP+HwVELbUEvrD7YIBqaF2nnVectYIBcJEu4tJz8sUTZsS
ZofycsOWpatsIhczv46Vv1vFwv2UCZ7+ZJUlEspWgzCgjKkylKqdg7WW46+nsAPG
65cShnRC+KSpvoWD2e6Ow8OMzWc3XEaaMEFyOA8Z0lfvDQfUi77Q/9pkb9Xkez+D
rXTJ3frQ90Mftnsr8bxpfKkFQ9lYEo2fisbdRxYx5ichb7R9a6MUISFQwiie1tjm
1qLAie4zigfhe09f9NZIjqyLtguzbaDTcj3VDZ5mFuLjXWkbzERhN1XQdJRIP7bU
02f/nzonXe3Ruj5viTX02HmOJ0nJsifxwd+dNheov0h0xl1DuWsQREZyY54CkRkY
uz/S4K637FJMCfrteP/PxhZu5HA3kS7JVat85CHo1d/T0T88bCp0wrG93qHBfFOs
hs/gTVzo2cqnfzOGkT1jSg8mL6J33hZHXcWm3GgJyDE8HZN/jagadGdVXz/W50lz
aoUBh6GlWyZefFd32NoM2usmlCAF4U/dR78JEnRA4TR9F4+3YOhFrwhU19g1y/Lp
GL9+AQCst5o71BGS1jBrkZ0LdXSfPNLssuJ0htHxQf5U5PyhlSpYpB5OObdgAhgS
WbN2LckXtETvKfia00uQ3f0w/cSAnjmNoX7cenmMCZMpj2mOVX5U9REgZ0U8TtAX
c3ueN2yR/U4xkxhOTA+950BnB09cDkZnZ4PJjqRFxhR5Ngq7ScN7Bwb7IJyuNGTg
nQ/q18nsNntF5NIcO7YkUVTBD/KOwHajXr/r3Yxo3AupIlgEaFeBCzuwHimCTq9T
3tpRfwdf12tNcTxjOUXuJ/VcVK3S15bpE48dz6iKxppJO1pUfnh203GYqf1wo7GO
hSE0X0q6uAL/Gyfq1iXDqa9C0nzxqTYUVfuY5rQD3MRU3lIZpK4T03xeUOsYb0ID
9p1PkY+//w8IxED1xJ9FAzWarCkU/OQ+Ua29H/uGhozWaEMiOyc8sQBlEYg3z5t5
yfvgRKg5hgFdZVt2sCjQ807nA43ZuZPUtReXLjXzVSiHqwp26ehaAyP2iJ+3nRVB
YH+B/AwwwheIa4iXXt3l2P48D/t37eFSED3hJfonLrDgJlkNsvnk49BC+6aQ7Xq5
SnNMYqnwKtAuuBodYGDK5KoLUgs+FI7SCUrEsyJG/FsHB4Rk0zPWixZcrTJ5w53y
JW2cGyVxlU/swkso81V5WspGrNnPAOflD0+IXlVj15PjhjNU0BZfraXma/fFjXYR
hc12q8+mK5+ISQfjmNuVaaM0QqgNIiHC76EPRm+fJ/B1N5kMVcldfJY+xtxJ+GK5
NsovHQutDGWetwpFvTeaPanpZU/+nnd4LVWD2AaTLfzZhFjSWZ+CP5hqjnmObeAz
ihO4EWDlfz0MSlQv+E4IIo8fRCkNeXtPl2W0UBH0OKycBjyS0og1laets8nPDzcW
KRkwf9Z/FuGGrwxW23KLf8xnm9i4B09LOiGJbZC7xyON75cWfLKk0U0soioVc/qx
MTgfz+BmC4d7//rvbkjsModpSZAcx2fuCkrHBaFRCyDGnR4z1B7GMu4hQat16+6o
ow3nBb4Aab8arKVHzfwZ2JWjrEiZmOBdgS8EjILDfIQDXi6OLSJuUo+tYH+rp2BW
/1+vW+ypRyrej44VpyW4VRr0aoV654wRrjNlxFOVMrrxLfE9cs74cE6fZpBgWRmS
QiXweBjMY9cMpc4O8hs9ViribIicGpoXdO7UkEwUhVPeywZcTfdEEeHUuA68OdSx
b1SnDAh/TVb2nhCH4y+15CJLitzvbVPxIMjzfBll3F7grtp1FlILWx/J1Ihvy/oO
x857gezaA2uiCdb4m1NV3Ua6+dtQt4YdNHzOOyBg2ti+SfJ29vH1khxn3IThnwgv
5BfhImShQRirpqamINRk22zufjnEbsYs8LIrdtt+OjUXDLrARHiTFMvYz2H6TRfX
5h7YgbWbMyw2h5jubuFq5dMSzw7n0QdlH7QJdAitnlkxn3wTlM2jQaRddcL16Vyc
hsngjDuc8agPBNB/Eij0PhZvRZRCfrEdatf+fUgQ/ydUtFx6R2RLc+F5TBSLhyCg
rtT0vpXCUZousv+lhrDFnxTo9A8Go7Oa6aKWvV0PrP1TiMLHrsZOqL6CXMmFMode
WJcln9oQ6LqUq900gdNSukhmAkBzTxVNFJ6z1eJ5+MBXgxTDAkwsFtYirdcfDRgK
khFClcDX58MxQejNu/ampCPIMXXA4mmDq7gUuoDvSWEjuBzHG6pBa8cNI3TOqkaf
Ov/le6XMjIt73sD+y1vUDiYKuekzpD4AqUjR+FVOYJ5y3CuPo7mzaxHzfgtBTg2j
rL0dTynWeSbzq3Wud3Bk5SunCAttyLuDquCIMLrKvtF6nBtNFft3s9B21XReNLJj
q4eWVKhJciK1R+c1JzT6bj77LWnDdwHx03E9xJox53uh0i3vbqT+aCGw97rOpaOp
wg57rZYGN36HtW87VpdAsocVN9O+PZuSN1y68fP+nQeAebeICj76pZW2hyCz0v7R
jnFgzUvDWlZNQk6/fYgW1LQ3OPyZi14I+Nc0CCltFYdjH5N6timNj8Mf051BcPmg
VooaSWvgicYIC2ENrbErW8+po2iSQVOYqE2dJFEptltS506U5P+f8syuUVlMIWRj
YLseolqXG+s+L8deP50n+26de5WyR8hNIUy94qcg7O9Y7KB8uKH9XApi72gSdNgJ
tIPYRryWwS9IPd1wDYqnQey2z8b0adg78RMquOH95OFjF8ybjMBdw+uBMVnqWoUs
n7FdlVe7SGFk2DxWFdIlY+mUOHj3nzEMYjTWUprVP+WGqMj8q6mKsqjERrMCy9jz
2+T6LaGgubv4wSrZPEawUwWLWHC3SYHrWxk6Cw8LhF/HoDdBPc7djPxORkv6m8jk
CxqXtJzuHng3/YMAqiNt6LlYKQJkettRMAAlB4dKVFKMbFQRkNfHlFkhHwcy+/uq
j9wb8UxSpuxZuQi0lq5cCUnsTIbS/Bv3SNC/CRdbew1ZoqDqsIbcDsDv26NVlpMW
MTlzvJo5VCxZjPfIzFn8K7vPJ7Sazqf0H2M7QE5zMDy4oe8gswuH61mjyaHkdid3
J3ZGA24ZxVzTfOQysCjCp+Z8CJxcSA9ORSNV8DFM8L5AY43anMhAkSqGjE0AYn+p
D/JfUOmm/wuZ7Bg4zPmc072cAqfURMs8+orej4XubNFZ1Qc2htN89mP966of1Y+l
Q33zkZUiMmcMqLzV5PoNItbPdei1JEIdA6LoaeZIZTgU9kZT0EJJG9mD6ssOSPxR
Qf2X4r4FgLRf/KuD3QHmDWFdDJLZLK7y8A6bmxGxnQOeE+0WQOZxxR8ssfHnCUOO
d4nbw6VV/aB4akKmzrd73bZZZX5R0Je306tDi+3YQjW2/Eq2z+fvDGqwY+ZK0ktQ
L0B7Q/wjJUxLpeiXh+RVyTRGO96LkyZj9krMAlY+Lfp/GpA93mkAA1Nhk/KyPZNH
nS1V0ZHPUyEXHJFnbzjfNP1nR6sX02q2pOZa1vruf6bi0clMe62TrRRdNHBFAByG
I4PYRDE7E2YRc3cXtivNEsVsIkpQ3gLc8n8r59TKs0iYhBPtcClWT848vrvdi+m3
9OJvUqNqQqtX3umdVI7mvlXsUYfEo4VLjUH633hfVIYSIBV6Ac82KeEz8I96jbAT
LLQ/VwsOYJOKRQULLdIq1FCvGJdBBxuDFZ5P8UnyTtqxYivDUamThb9IGxv/H7P/
OL5K40auXbjlJW0PeY2oJbRivZJ69+Z5v4rFeOBAOIWRogiuYwjjKpAOKJ8ASf8s
BqmXKPr6R0J3taAhbCDFAIBGmZBztrxw3BPuSSRDvexVdjxGu7YUf+EWenS3CWwg
kBYRfx0xkDHYUKDJuJkHUWhq392SsAl1fKWRcZSFa5kmCMiL7jlVfqhwFHQ3P10M
L4S08awZVGSraTw8pzXcj5b7oo2fHeucVI/H1mqliuw8DsfxJOMmDoDFki8gKkSB
7IcP1Wvt0f5sZbve2Yn1hJBaERfHIo+NNJFfLeObih9UuaF6B3uHDVGFTAaZ2Lem
0FkYrC/ZUuqfn9prpRuxsf/eoAmT3sHtK5rSmNHF2rISKXSLjoevRR3uoZD6alhR
fWMwI8FDRwcyuI77NYogF4rnIBLNa2APtHT97VaK4my0wtUBUIh9QBfmsvuKGgLK
hEBCkSpkOO9OvqVpM7ApwihbApaCWkQOj69tfsAvSCLGTEBTkLr7bnxyoM1Cz0wl
mahh+7lJBc+tzLpwhljMHyDsTdUeUQeEDJ51IytblVS+FXvyGCuSgCfHM/syCQiS
GRFp9976vU8UmzX+XtzuYTrD67NHaH5VMgiB67iNErSdKqkcQpdwODf8N1E18JyN
IQ/GGakJG/L8ItsL45qbzIivcn53dnkbksj/vO3hkn79oYEVfdhcEIQfy3U4i1Se
te8aFgTCgMTX5aNWhfPe3wrTqahA2PG3kSBPkdwQnmSM76ju0uKiOsaKRT6+iXEv
1h0X4Y8ERCK1IjVeUlp9AEGIqURMwOlw6ejoZ4dFjn4OxBLekWpBbCStosxyaVVf
1hILAecuecVIeBLTCIobEZ+8mjKniVv04GIuHhOJD5Ooa2zPipvY5wFsitcX3D2p
BL/AjM7pXnHVoRlP3qFX0AmhqZ3WFcp8tj1mLOPqGt8Wsi6yrRm4KsC/MOxey0e5
0/4FuqxrSZaCge4M106nAhF7TR1Qcb7ARm/mw1/xaexRneXSg/AFD4o0RflrMdYJ
78tjYE5s190kPQiKwJtKj15WLUnbJJFnQZ659nDfv1tXf+MmznDMDoxxMLuIAOFZ
ibPCsdg+8cRptFS1WPZYvWs8vjMeel/GV8mhjBckoRUS4TPxZ/hZ8fI7Eriuw9bE
b+YMu5UxrPea42+Ox4x6eG27Ek6xMJYGWDJfeIhG95rKb7JgHu6n79AzhQElnU37
sP6YugByUXmeQQAeKlL7/wpfFhfxCddb/u8CSLV/W5pPNoOgc218aOlW+I+OfrSP
RQCKR1STwncOzY8za+MKJ81Lx49QNpeq+wqJsBzLvDqZNA+G84YCyGvhcELdmS0B
TnFFuMgLkplAsSGVNXNi26QTA+1+/hNpwP73FuhwzrQG0ZM8XdRzL6dGXMyEI7Mj
6R0ndwg79r9Iy3G/CzXTwvBeyPxIwKwj9IYce6ykk+XIemWMIuHJcGcyL8w40Grh
SxmuIc2FVXqq6tKjiwPEJqZHf0YuiuT2HpsJlVAyYp6yqmj/Meyggrj9+VASi1EU
nIkyi4HsnPzx+9svBtR0y4c8u1qZaBtNzfvPFdjrIbYcZy1J4jSkJSB1rpY76i8f
bzhTBTKy6sKGymvSmy00D8vDwmDKvVX2YyRstZe9GnQOJ/K3k5yFrv3wml04ok34
B0WB5ctVQoR/3aaQhLlsFG+3k48+HEyx/oBwmbAV95LAheRm5Jte3qstoy9yA6AH
0cJsFPOFdG801YtriPKmjMLKnfNMBOMR0WSB8/ebEYd2OxLT8WpoIlyY3wJHQzZe
ydFq3yD5Lq67K574wMrJu/mfcZ6Co+9jOPzSYFqOuyuU2HZg2c+i8IjnP8RqI4+s
cdneJEuipH7BJjHbzpcbHJSmvBvtSnpqbHQZxPtoZzar/lm54cZjT66lRVu8c4PN
SamrV1H+n+h5FnTqCLpIMahcZI3oTWAttKKYiqHqk5QIvz/TQ8J2Anxf3JyLxB1E
cnhjRCZXojjyFApp28r7qQWZ50lpAHoOlr6csmhqyNI2Dw7ky/FbelYUNdLnbeUB
V6MM83IADewJPdiJy7Cp3tnLv4695/TLyfYX184vqma+fThGj9ceCmJh0AjgB7av
fhQvvnA+xSmXulUggeZ13M13pLF8hPPd0sQ7ZOom6yDCN+BAaWedxyTNIv0kHGhc
zoCBBpzMmGRqR5KDgM7+uLDBIMAqh24K+zO9lrDEs63SFaAzGlc8aNUMtOCd47hX
+ictZeKkmuCv4S7v2BSj4pcRNPKay30r0UQR++t/9/0xdWuSrNi7ToylZtsxmtW9
J2bDrftxZdphcojlqpRkeXu504CLtph1V+gt19bY+QHaLsb4sM5RMj5Tpj6m9sGW
ZmArKbWnki1hSlRMlXQGxYR9xlS2TTAIYL2cYw9qthStaOp5q28/J1iAnn4pZ5po
B8i9iwC3teLIUyqCfCNVI3EeCrd9sKCMSgdgqFpy8JohrEang2iVMrb147GdTx4t
R3aentjw5mOe8L/MoLyddPbl2O1Ifq1H7X9BYPzFPNyQ22hFoXkyn8YGJixQAkQZ
s/XbpuTeNF0VijeQJSHWCZUH3c1J2E0Crsu25EWfSknb+uf76R7EfdwRqmfJQgck
i4VK6+ObxPcYJ9tQzROEOPfWVmG4Sb298BFE+QhTzbTccrDyh/HM8O0Lt3kPcfW/
+K8+QxVMA8uqdjF/7LcwgkONf5/tNvOIEpSVpvJoA+7Di+7+xzwfYTTa0Tm50ufK
+wNyCHGN++I/sapyqnUxbjxooTTnV38NfqbAJQLoNqYBVnt3C21OvhXvbHdLrX80
lbi1Owai44pBBMbub/8Q76/UNLxv9uYBwab5t5hQLkUNw3PvNu4dUaIVtCVmDcNR
CnoRBWefEZFbpS+KuD0atzSVVXiTxfc+brr8xWW8gLLdlbNvdMDle3Ucs4dVJKVg
QUDlBJLDIjR5NEnfW+BTKFxgz67DudHhHFvsEZmbN6oPF8pqcHLwsNNexmuCenVv
rA3cDa8l86tALK8/R08miwmm5DsYVPGF/yvq3Bd9Y7uEWaI8v7576JYOY+bEsTKk
JEqDpRoJCBkf8YYLdkaTv0iAhfYz2YEvNhbzwOFWmqLrj/XQeevg+RCnK9e8Z6IB
l0Qod4LSNI9QyJe+vF+SeIlUCZ4kHhLnJ0igZkvTtWczkbDdNiIrNVzcZK2A0Cyp
ockhMU97kwGmVMjiENonXarxx3RjNHZcx8Ag8ldQiykCEiv8kUTsazQmZ3C/a4BJ
gACbwrUSv9Kz6gvqqOOtIPFN5sxw7PpGLUWCJ1KFRoEgfpVS5QbFf3UdE6otjHhK
6GZU/nX6Pa0bFsG+ykqLXaMCHsh/a8VI/zhDVyzLiZRsHYXiSfNDXz7rmmidkU4x
yZy96/lR4cryndYqJ0QmNw21f2K/n7cEpU8xTSTN27TlgAjEvmz24LxZvlyeE4U5
+e1CepYEpqyNTNKNVy9cFT5lH9jJBRo+oK9ZEPbYm+WgQxDc9g68MIQlHlojWlBF
Jo9YZaWdJ3tPjaFZ4up7RMDmaIcm2HrP+yJ1Wf/IDc1owcDO3VhMbx02MQ6pQKuP
FMVcHDKmbkLEVoRl84kCGszsxCqhUTE2dfEWzdkgVNFm58B4wbq8PFyKdyvmJbW0
9nKOwetdDj3aGTmt9GF33g2BBhpaXkZovRZrMDmmfHNl0a00HJhuoNiWXN8jyTYg
fFw9ZNeVzM2nnyfqrU7fkNxyLtABlzBGXOoQZFXfEQxgRBfgNQN0HU+qkz2lIiqM
iAisFykXuUloNUL/0CpVKJ0ByYr9n9JPEIYhUYuNJwjgWT479QiH6glw/WwVMXmO
soCJkWRElToslA2QP6mrlNjEaI/xsi3zzWND5ITKO3EGoMbBFktuWxh9xJTXzx9F
3kUBq7g2smBkWPIyxEFOlEQ8uwpCD36Jmryx3Gh+qCYwWgT7xDpXQSJuGHt4DlyW
o+72MUJ6lRuBLO5e++KwNCeZHESJ4w5EL1bgb+fq5QSuoupQ+sLU4hKMCZRHVR6b
6Szg+gCInfh3NMV0Fy+NUuWRhpO+Koh/ZLvxRgAqhsChhb5yBh6CQbAp1TcGIpmG
mAFO5JDiz7Ow5JIpDGU8gpfxJFY1qYytY6VHzx6/rg3HiV2nSRTCS3+8i35OWuMy
bElHwSFoCuW2stzvoLtFBmRmbYVU5P7A+5S+5Xqh9idZ51zCtOw4Sjtjl179//T8
ZcwJK44h+mYsP0/QKRxi4oWAoszQjXJj+fLqbqG7cidyWlcUsOcPKv88frptI8aT
b7x3Ca+QazCspggU1i5rkSr8RzzUZanku4E2YNGRJiLMybcrBvZcSSLqRhdCmaXU
7uC5cNPuRYxq/yx1AGqoiaujpCPEC50v7y0132cS2qYjnTvJXvKTCNCI/bjKqJrJ
eGRkDaDT3biILoIR425afB4wUwfmbEyJmWWBEwPFObucrdvzb60DbFu2/cCoSLOV
eYf18GcZAsWCQpt7X6nfv1x/dMJTIrmb1XwZRCnLXrMjkIKephYZpxRgvdKkQ/F7
4D0ubRVx43KmxUQG0Efl9t0aRKODxyhHzQ8ELeorMHi+vNvz/CZbVxOAGFL/lnIS
ABHqVBv/I6DW0ZjLCFoibzBgIh3uN9UK+Se7uSEUttdJFdDzcIEfVkvl0KN+wbQl
vfpNf5PzKFz1J67gok0wnrLDRw6wh4QtUmpjtfrUqnl9h2GzfkDUkVAc9m710Nzu
X53FVBj6GY4QDHtkgylW3t3RlQ+ROIMZxROjxSub9+/Is9m2zZU74NEMz/kA4Hpd
A6e9zG65RY8aK5nikY23zqC1Jj8XAO85ZH0Ynri3U8c7mGpOmNUVvGlCViSfsEL7
Z0OOKHMvXHzojoL9mY8FY/J9bIkj3BDAPzcZBE38Nl7HiPa2f60uchFl24cGh4ib
7Auj6uk/nqOv9GfuCGdRDekYrNIuObUsQh2TqSgokfie44XfQA2SYgvfcpZwt72o
dqC/UkVU/qM/eTIzhVvFcB56udhD1aU4cOMd2RPm8jUKt3OvMjoYFV5O2yq/H9Sb
eJagL4LEQETiTSanWPTwbUelgG3HmzvB7KrwqbCSwWapLNIB7DeUuSSCxPw8FefA
CW90CuuXcWzc+I2bLm1FR1RWszfaP21oTUVQT9CK4xDUYwsXCWPVGlUknSZYu3vq
S4LoK+6fgJ6d5hxs+dnP2r3Gue+zIRJS116W/OUS8a2SpMJWevt6yL29IWBnwgWf
VCjtlnjLgY660eEZ1JkkaUcUkBm0CQXt7tnrX4BWhLo09Syted1nLedCQWaOMSAR
k6VSQkU4Irjzw/nOp6N5TlqfaNjIXfAJuKSIwsElYYgWKVcYUrOcgaRAk1dVqzq3
cVLV6GcH/S4rgV0jYQtRY4OPnSaMqFq3G0+5E/jN5g5LJlTwAPwy2C4cC4/PFyaU
rZQPtZzT/bCw6s/13abkVdTrxOfoPMOqjDCgWl1AyY41566BW7PteR3g48HfNcrh
r4GgHM3O/rZRda6XR13K/vkit0ehHnWvZDeUb8D/x4T3n8NMR2M0suzLDuG32zjv
d0eW3cqFM94mQC6gR02FRI8vEy0NvBkK0RQ7q9cHB016WhWse4fUD9Zhrlz7r2CN
HZElvg5Gf/RhwC7P7ZO25ybrjujvE20UBwejPYxbTLmzPZc+0GyxtCc15rCXJdLt
d03+gDzGeRTfC1Qao2Ff8rKyU2fXgBEGLPHknNh2+ZLCCV5cRuFLyi6YxxXEaI6g
I8QtlutuXtK0dYumwLo27pP/BaKneEDZpsmo0wxnNiiAooOBvTqzlhITf8CFUOfv
R01OnYW+eOIn1BII7O6GA/atmdpBEqOBCIAksu2FFwmHDH1cXirE6ZLU2VmscrWP
Cz6nzIXBguemnfONoekkg6oaUXepl8OKxL+7sTJ60oscJvwJJcCKhbcM+f+6+rKQ
Bh5Cnjefi7WlleHt5K9KTWJn0DikI3j0VtjDcBwkO1Z68QrbK5Eoj9daI1BCwEFG
/MQcHGpiH1YdP9E/7Gmnj1b2E8MTy3dvJXHuYGGG0k4KKE4mQZyire6fylPDsYFF
6aXZUkh44D7xQzH0iGvGSyHWmrXAiWkllLS5dVTSaBqpX+lEr1gdjERMefMbDavC
QYao8hf8kfDDfYSPP3Whp/Rwjuiz2PCBMMQQV4hZeKrSgXBdHty2zD/8LcFAveKo
I7begygJ/H75vksamKOV0p8bWQaoQm/iunj4BlMURU6hai4kRXRaNSSFycKXYq4v
mB08oMXVvqSh4Md4RQXmY+l96tc8yeappDqtTGlrszloEW6I/pfLgFSJWj2G+8Ms
BtmLrPeNG3vTOfwGuaTuAT+uX8Nj8HyK6TFbzGdMx5Jchqvt91gbgjRzCn2fX+DE
4jFFeMQg8mdfIEiY02mn8vL43gWxeF1duXpIEdwhv1Vg1dCR6O1w8rt5ieWD1nFq
KUYvYzpR+fAa5ADX1Xrqu/KK3rMLgkdIEWFjCPjx0tBS5zxA6X/3dpsqNjL5dJXM
vnQJrW6dny+8nrXXptsv3JhbxL4W1zQllhXeHyi1XeZce9BfaYMpRzdBkHgmEzu7
U4RFcR+tsWcQXE/rt+kH+IUoLFrzJJN8IGkxZ9LZQuBYeoMxK1oftkQP//aI3f9h
UaycPVs2B0oNVORZ13+kFbvLios8OXHCowgz6zxMAuAFeUTpnPDVWzeJTpIcVJku
sTUkDQKGr+Kd4LY/0MjByK9uKNKxX0SGAncJ6e9fKlVzBDA5DYpDiHRxj4kJJIG2
qU9G0wEWZc8Yi69Gyg0zQz8EXwj/bz9aiCjnnv3c2g8RsBnmjDGm3OWHr2MUoA1x
cCUWLU84RZsXFYTunIHwiLsTbxEnUcLhkoz+RSb3bfL7cZXX9c0RUmR5D2JfXhuk
NpquI14XfR9Zec4lzoY8djNyl1aDxOM+NC5RTaUNDISTmGNhvzWS/fs4rEdhFBC+
otCWOYp+D9iHh/T8lnsBodqqvIG/kdYj/az7Iq/wHETy2gGio6bnQXPs6MNywhAU
J3yic3VOqmzoyJeI5+2sJ23qKuQ2W9FBxQx7yA8sXA2A+Rk0bnNw0sSnbmue1pdH
xvVhsoZIBa3qywfG0lQfR/X/ZhWZ4Orgw0vi21qqLfMubQjm3AHJ5kdOXUSz+xLh
PogZ2AV3b25rxEk9m3GoKnk8/vOwCPfKEz0GJf7BCMXtzb3cYkpmhZ9ypFQCIcZf
5DAbdnPm2u0WZKjQi6uBvHhvuo2fsyLfSO3nlIw1jVWpiZBHI9VFqK5dHWm9AKKX
+Qtw0r80hiRnC4Eh1iOgmuTQs31xzJnceyo5o3i8ofmUIxsn0WakV0nS6UVpGWzZ
r/02ElNKxqgx4kwTpw4OqLFYldFJHNO93HazVv8CLBjzMncUBCWkXFp2jDcnDw0D
qaPS5lXC/RGkcF69Fc+PvlIqioO6ZJ/ztA4WOw+7flsun35GsKTA5j5gZnp1OLh2
fGPb8bu2gRzR7vUDg73oLuNlImtlAhav4p5AXT9NpHmuPlVACkL27GbBJAlAmC0B
hnYdQiUBhdvvxRO5f94K7BGpq0QzHbW3czr14wf2EzMFFHDnyffkn38v7nAmhv6l
oYBO6M5AODUW/lb+7j8QlyDXEy7qndJw2BUxiUlXNA5E8UsyreTTV44eMKlWu+tT
2fNh7wrWHIFjSpPNu99+yJrOH51kaOo6ERG9bgVs/xuKaxoTo55MFSAejZ044+cX
fQ8fzuS9YoO996DPB5Y5uzn98BL9VGMSUYdDJwugEVycF7sLj8r8U1m/koWHwhEa
Kx9Gw9Tdvqf2chvyLWQUKgCQNubgEMO1U3tDqCTSuaVYG7v7rR2BjPYs/A/QLZ/q
WqNG5kB3BjAGxSF6r58TO9/XWeIA2/c3wmGlhO1Cc2+hC87qFOf3D1QEUesd9bpM
Z0NC8/N+YrmhEqAWG9BhJHTNtgRvshJlrPAg7iURsy2nIqT3IsJkfbNW27nm465K
QU8Q/ygAExsycHuQWZIEuwdgp0lCgvErp2q6cd5cHhXEytum4Dt4FFdTFr1ieO/q
57tFYRWBiJVsqOBg9RwMHhWCROF3JQmQ7zZXVW/m2XaKpfbMYATjdrARudtb7x/N
qhomtb6PZtRdAZ3MYEp3dHtYVWPixoskVw4kxK0eIHM44X5VAuM0l5L8r3+WOhnH
qzNP4Uk+L7h82AZTHafKAzGAeG/+azvhpoih5DhvB6Plg+BPcE2qp1O43cDHiHqB
xKawQ+FUQO8byOI06msmTgS0Dwf8Uj5T6Mi1NydWshGgH9jd+OxI2GuEPwJ2wLnO
TUCbm5As1dM1v13IKUdnOZG7Uq99ERJd2NDLzqIHF/ZEDlsiWVr4CsBspudbEu+H
obQ+dQB0wkvzn4ZGEMZVkb4hdKeoL8VOgz05pPxRV+E1cjVfRnZhK9HpvMZUI6Zx
SBFjP0ia2PjQPzIjiiYeOkQ+4HuwX1DRA5j6bLBOvOh/HLmLl2RdlgQEJQpS9Hp+
2YR2DAQBx6zUIQeJJJ1Tv3cpuAMtLLVmghrfF6U6eVEIVSBptYcg9ynHkv9Haz+5
sXe8EGhiOGXoJmCVqvc3dUjqMyiDiQH/Kc9bti+eZ+QbtrKad8hxZ5+cbdaHuaTJ
xCS2yQ4PXw6hRGIPZMXXYOtcivVCpTyPFoqeAZtuL6ZbvZEJ5AJHv56T50Uo/Kdr
kJU9Od0S23xqhVoqXhqdwvdYF7vIBir6gqhkOV5IS+3HEzOBFjJREBuibIM6QJTe
NUaJpvJAOtcZNn+uY1J3zacOi677mzCO7rB9Fu65ZBIWJ8MHV9YPaZqu8+ZCCP5c
SyfP7K2dVpDDhnk6luDR+qY3ztYdW2fwfKgbXzZW3O40uorSX2vK+cRoWx4StWfd
t2eZSNRKMmp7ieR4Ox7yTXgWAQrdDEFmSb8Y99zTdyoVCrLLe3X1Dby5cHO14ZP3
/Os2yBHgGbt/K5Xcf6gcNMbuBY8DjYR1E6B6sdsKPnnC7Yts3rNarV5p6MbbnDDx
Ey9FvQ2cihEU6CxU3SF2uGCOKPQUf+ytws5AabGx+wWYj7kfXILZea9T4k1jLNp4
nJeIxZRPZN2SrW8+sM/OHK0teEKvUPs3FOIfI1oEg0W2Sph/zPbl7Jhf8aWG10nI
EGeqvAj87oALeRCjfFkGXKYXgS2HF13F+QsKo3RchQPGxdw/uL/x5nDi/rYhitQZ
GC0w4tw4DKY9Hl542tUOZm3xK2Gt9UTFRXHLmqiM5BSy2Vk7bzFBmUYj++wJhRpM
HMwFj2KxJgtvopRVbXTuHbtwr/Xmdk2NHUO9ehe44yH6OUdVlnoVzKcJNCi8yvr3
KnstPfFOM357Ebd9gQkLJu1UyfN1FJ5l8COlJIpE3Y4J+PnZMaKElN2jqeef6ffV
Ja8TXVagFXeG45hQDpn5ishBPZf9R6KIzVUxGvnjRogIXzav1l6nRAjOuVX2WoXY
nGK2jnCWmYbpH/pUvTfaHnmAIHlVlGv3MGFjNTI0XdjHYgWr4OaPVMpFtpxJMtRq
hmtXA69Ncu8SwqdhEqCP0A89x1uPnqw6YSETmmrDfkw9iQmDZJyTY+kIybDmvNn/
cewHOijX2zoeF7CetWep9X1c22UmdL1iDNC5nBnSlWd2Q3llEFYJV18FpLJnm9h6
71kMlQIAh+mQvDv77Gg4HaTZVhf5IYMESEgoJzya68xB4xx8XKJhPBS7BvVQWBJL
GoxjEQY58Yxn3VTz+qBALZJPEq6r0i2lNvwzNZL3o8ou81fDqP6DI1Jt6heNJsw6
xWalgMwt1soqA/uq08HlQI5ufEo9zqznqtiMl+9b9It7ihJQrguSQk3tR/P90irB
WBSL4iH5mvcaBHxN34ANMZ8XRL4pZhPjLsFyLwOoyaxqjnRtBx33WrnWeQJK5xY0
jLdN87tybxpYXk3i6/oncsPLTgerEKuhxwlHybb+NgNSGF3YbishqlZqB2d5l812
I2ZPaW9Uq39Zn92Oo8ymqTWV/nNtltbttkO5pgYbAM0vf2rZQ4tAC0etCD8Pji0C
Cxhp1GFQc75wnWk/8j4vOudiAm54/vdad8YgmRpPg4Vy7Ai88jBIm/rwMzqP+ry3
GM0zXriTK0GoOdv6Pdl0CwgdlyfX/LbHOUNEHwfOQqXUSSz+UO6yO5xWjSuKZyl0
1U2PtTvjvpA25BgGL0PNxlNWZJtR/h0yuSXv8E1IkprfBlPrRD76pdE1aTLJRvFs
xuupVPh3etyU+8nNB0iG1N1vz91zxCXSWZ5Usgo0NnY6VIwwnT2hSwlzPfQWuabf
hO6y2+r6ueJVoCfIjwIfpz+h3jDPP1Y0cCKaczInxOJ1vEG7sryzLbrWbA/fIcZz
oqXPBPKx09jtqrZgDTTKsLLas5njB4OEEUwlx0uBwSBtdcs07OF876J0RrtHFVE6
eUEUgyywzTzlqPE9aWFidex7QuqbBnFT92HGbOlrHXfGAG5v/Rdh2JtQk9fKktf9
qvjFBOn4UgxpbpWb+FctFB2FDtsRp1MVYzkcl7GrEUHWntbO6QO6a7OiduB0UxpM
FmlFKjwk6su1QSKGrwDbXUvuD9tGZRa5OgZca5whrA/YF0sHOBgFICxig8Y/lkEc
FmKkEdY8zH3CmseVlU3GwX3EE92v2CJy58dmUlYTkLUaLufelZh/L/T8agc2Uect
nvGkNRa4s3acH7NdirP0gJnHU+v02ozRECyqkusVohpV0EAeBT26NbCVmmqZNxY2
vLQy/V1H17hNP00C/tkuWbw+utONNfYIkyEap/XqU5JiaAI61b05T14P8Qbs2Bfm
ehTqcYXqjn+N5uzVJBpMvodZ09iDCmf+5zxk367CQ7oC5srO3b+TMgFFwzzyCP1K
CvRE7G62LCkkfvA/et5PjGayC79MSqZnVxYRi1cWW4rxDbokCczS+vDZOEdbQrwZ
4Jpu1g9f0Dk86+EGgMwEMg5ss6m/yVEkw0iaUE3pq19FvVfrPuMbZ/eXjCoeo2cm
C/+f9g35KXd79j6YY1LpvOIDlMUi5cukv/zeV6B93gRa4nvp1Gy8hH+T5ez44Cus
XEsvaSiioFFb27eskDYQ0K1nNiSn0GPBX84Ah0bx0QwW9RgUpqEPBYKIwryQ0Bod
MR1JMVKE+nSkXJIA3UkPXSD2XCanivx6Koas/6VPe+NEnRuL2yUasrC+/jVBMTcB
VKY1ErxBZyR/nTYMfs59TBuEpKF5UJGkc9TrudD97umfZlab0wGkUAiX0h0X+co3
VUnE+AQv1cHKlJb94iDo8AE892r4FgHfzzvXOUdu1mIHH4Qv46UKCshtRVG4o3ab
sneckjJAW1ZyZiZNueLPHjPyrfr9f/voglpHzwWujumkTpd+w7h/HqDBgDuFB6GQ
hoE/DYdapDq+REzHJZ+oRoO8sYqDPwNDJfYMz1BJQjLlfJrNWrq+xHcehFE58GR1
OaJDwb6T0R+xToml1Vp7EKkatWca0yMZbF/gG+g40IOwX0mch4UU9HX6VVN1beqT
TJ/zLr2vhE2e8mKQ0uK8q2oaMGz/O03f5yG2Rkgz37jZ7Eph/BwDu/yU7SzazOGM
y3wu7aZ0zozC7ga2G7Sg+ptuhEMWgfanob0aSq5+ur5p3iw06A9S4RGz4hsLDuGy
+VHe6UlZC1NN2XqXuABa1psA9OwChcVD6BE9JajzZwQazLu55IwnfsS5FCRUeVAP
iszcn5Yhh4lmQB/olhcyNzKNYajI1x5tWVeyVQqkUF+AG1ID5JOZgEJ+Evj6AtLw
GDX9GIfRUvXffmVbM+QYrcCLTezI24qEtVhylIDPxn1cl7EyGuVPjJdBCvdQO2YP
PMwkHwUJQWW5o7LtLgIhZwyzTdLOADutBE/Pn9ZJqHaFB6f9XX+wRaDC/+VKpTVe
1VKN+mum90xb4ZIyNt/AAFhusWAo7vwj75H/t56vdb/EmFPVwd1kjLc7VgAJEOL3
BFgdfYEK67yJyFbRpjtS9HFxDoNXi8eRj28bwPFreKL0Ixfw1smtDBHDjBwrrCdV
3npNmXqaJl5WGC3KsDbFnFtCOwq9X1/pWR2Bz5BgewFKG+Xs8d6zfetoJd3hFhcn
M0h7k2A9slHaM7J4yZJbKcLye8N3aIe2kOBEbFeJw6zlzQi8NV43px3Qonj9d+rd
0MdibBhrr9lRdrxJGtac7dYFo6e5LbHt33UNcG9k8Qqn+M99qSkJGHzFqtp9niFv
CXBsCXnymn/Z6zNml/XsoXLap09yvadef0BFq3QqamrO4REVN9IIUXFAFeSvIZCP
0bufavLF/4igmG+Cx0ABZeyHaykKdUvIep95HEnkqva1BjYuHowSKEaScK36e6Ku
0j/vRFqaGhlyq80lS1V1dBMStmr6Hs9OyD14SB+evwNhmzHmal3SKSuh7XnBAegj
dNXISl/tM8PiytVE5r0GW8MRAnc/lwtfJPl2It5dWMCIXxxeGYxRQdT6cQBZ00I2
xj8kLFQNOYPcbFlhhDlt6RLy96Q7dLirF8E73Tgz3fWpk+jN6mlfNTCjuZYbXiwd
88aU4a7WPqhAZf8fuowvb5qUdmOwjVNu0MoQC2eLz6na42eeDYa/nI+lx3w0fcR6
qYkMFlddEoZ688WYAvkwX7xuatxFMhY+x+72bkl+BDHc2meaS4Gh0Sxj9WjHNfp3
i0569+yeyfhaVMuzqamY1bUsVnqKHpTp4e/X58pCO06HeUo336K8FvYZdRrUL1+l
tfq9nLCw5NWCPsGSO9BMwFLX8x/3wB7cADTCGSH6/8Tj4iT3G4G7qO91iYE+SDSd
SoQXU8MSKxuRFnSchBoYYxASxZ16fTL2Pxt4j+bs9Fuy8USPLlbbIN1mZVdo+1cU
QryJIj6NIOJpdmLoXZBBzR1J7Z6olXookNoD1a+vGAtE5XearxZca3NQ7z8LNVgE
utvvEczU05HBpmxKAxK08jV6BXRuA9jSHk8KLuso+nIJTN88ehgsdx1fmANufLRM
ypJs8zio90kFijC+Kax81JKMJFU5pFOzVmd6C51ZabOtsd0vQy2u2qA3dFiJTvAN
TsxWb7LoC4MzrqEqfUo0EDMa8CoMxRuxEsw1FU7DvByA7BRs3BtJ6mb9Sb43vZrP
UnPE1xZ82nmtE/LBYJxrz4lB/NHHjR+lq/9htBRdt/1DvmTi7r7vtMfthBX0ulms
wiezX571r3ZPks/+4sTGni61DysPJ+dYOPJTwSmKs1SNvEI+cg9Udc2mlhmRLqwr
4ANrUn5k/+ShiqU9qYv2tWfS+R5XGX/FlYfQtLMdrppWmB68iyDI5q/Ck9AgihSo
kOqy25XdU4olVCovuuChMqCDIKwtVrrQ9SPFeF4az1kXY3F45w3VYTyHhkQKbbL1
6HrSWSlI03MFAKX7tyVf/p0SnX0MJ91A3saqA+ILc5dcSyu2tXTHjIkaoS+BODnp
cuJ5SPaluzOOrJjvE2jsJkbSTOF3CWI2JXtz46HU4FEyjRoLto7V5mG0+x6xbueC
ewM64FHIXpz/B3zn6Hso3De1vYNCpnSxMClkTsDcq9JCRW5UeCxi776jyF0Hpl0k
bgJXozEFprP7xoPyuvRcZZSUrtBFzTngf6SiJ0t5+B+HH2qFSRlcj28hrvoXCYiX
EhigYz9ykWT5aMPmZ87kRwB8tBBaRuAgSr1gbAvlVXLifGXvAI8/MyNkbtj8autQ
SvflBwBzKrYrcwjRH7SzsCtYrgz43jziRJ9wIkFv4kuov6NQQP5WOcHPKtV5ss/H
wc7npfX4RTXaLHHtirQrJxtSCkx8SwUkglWZjdZ6iTuRLJhGYi6/87WRq63N3zzG
qc4X2IEUu91WvCMUmC9dmDURuLQ+DlFsvqK8COvEfWhHDXreooaJNsbxkWqLOjo6
lJv4ZmBVncqt2sEtUA6hsPQY+uxjzTzxtxzmPd1tn40nhdnmK6Hmp1TrTZXGSgil
9ZBxkiM14DzJZp8zvgH4gto2pKfo6trUg3oZdz+yZ7ikvx42zP+7uSlZ1tupoSKW
lSDwwZUguAU5KEZMemcnooQvDqj0p1wqGdI11Q8wQtKqSt4k7wexXdPWozTTWaEp
YUTlHsToX47fC2Af+Je+0mjZ+w25U30vPcxAscQTeyptRv+tbMxGHQo8jHd6dYxf
+eOoHV+1HksQF8A5gudKFwfbsev49hU023RlmwkErCjudt/hP718KSwwTg+95TrI
BhVJzoRnkNYkdAi6HrHT7Oa+AP9B0mFhOgRu1BwP3tWX89AU1H7JCnuvjTRG8VR+
hgkEEnNMCZhinrTaQIlII3M11+QFSeCyDspLE/YU8m9Xytq2/vPo1i4xyBCXW0ds
0+gUhWnH/wS/SHfLnlBeyHLHQB9OGd47jj+5dU3NZYWppMkT8n5DYVBJyM3CRMfA
M11Jsuu9q5CuZcl9A3rt6sp4B7eP9vQskanrUoH0X+FhEZTk2aEbcF4Mh25u89jP
cTdbpBa6lcHVi+P3LO+eJf6VbchvTFU2ptmAaXrAaDfCz9HQnSYURzLFN1kVuPE9
OhKvSs0AT4oZikR5yBaPXlmNuoVz3a0mBxHSPZQsgtGONGqQW5Z9nKtMUN8Tklsy
UOJK+d1ZgWKb7jwnb55qs2d4IwzpnF1we+4Drgyj4vWWX9pYCeaUQeEoaSi7QDCk
hsxtolzplU+HtHmnVQNU7XjZjvzZciwNFYXGg6YokAy3bCUn2r5T/BcPRzIINCdf
iFTWtiUkV5cClC9xmxEAh7K6qk67cW65GmV3btrc8xHU9K6lsBLA1V+az+PTKh+B
eNa2BgCPiDXArqS59Vzl4FFlUgn0Fgb9iYpE9QwouMyPnIl8JgiwXyObGtlN+qIS
b7doAT5+iSZR3Tqs/GEtoHH/E/amDZjQ4GGR7RO7wSmFPMolOU7+7olq02laaSKO
HzSFt41UyVR/58xSbkZFIryHtMOfrnoEP3jlwItOjxS0oreH82JUHRy/VyRsbjCR
A0e+Wtb/OEX7tsWC/KW9AEMH4XAWGgfTJCZWvjKOaRqqXtF0K3oYGoYy3DrnWryr
ooVdwinZthldjjpBk2lkufzmsCTU3HxzDdrTBQ+3MthIoWGx1LklZ/L3pXcNU2B7
n4f2efEg/RAN99OBf6E0/Kcax1V9cfty5iOshwgpjShZZe15N2D3FKizFB4hEWpB
6rU36ic4ZUOTe+7vkE3uNGAvNwrwrJBtPVrTNzgQP8inI0SPG2bn4+qTfuC0Xtrw
8CNmvli305BTNuKBk4xQvcyZRN8YlcmfVIr//MgbUjA/EHeko99YoGTKzpUXD9ZW
gWDic4Gu01Hp7pe0rHh7aIbIlXYi+zWMUggjr22Q+kXn98RhY+9Z6pkjwKUYWNu4
1LlDGgZFHw7RwzZ5eHyfTk5rstC8aiwQiPmunHiNYxr6Ui0GYxQ6DBK0C2vUWWhK
S/Euyi43FWi35KvTXAgl2KPSny6z+35T1BGv7FmJdlePt1y6ydjCELeOyo9PGl4i
NwyRryxcF8S5TwSWWJtjDVRAEhg+TwPIJ55sH4COzeBMGMUEE5zhzVymPOGIG0EN
ci9UH0bCUdoONGGJot7Lw6mtOEed1o6/1FnfJ2Bzwrg+TPAPL1s0Yc0RIcS611XW
ZuVff8fyUqQo7RkuQ8utb4qElE+sxEDFRv6wyz792k43JVYMM00Mmr980pbU3zwZ
d710VP4Nm49q3EdY5Y12ltzOULut94iXIKZ3q25Y4JL1s2g40SLErautSpn0S/K+
S3zyGFhingnwdVdasZZxidAfwR58Fdwhpab/l4zx1XdpVGfO4ma8rfoeU9OvHLit
z88yOUiCzCbWjsNRPaawycgDK1KlqvBqUAoRlxGap1DwapG46OfEWddLaG0f8Ybt
lZTGROyZWCJbUYKzfcIBJHPVXWTn2lQfzfPebdKxuv4A1l+9rfoxQ2RqDrgbZl3D
4u5WtoXO5IMMC2mKqSK0tJirSZTME/qgsyyEMmmGGuQndbCyJaT2qa6xRfkFBtZf
rfFFlmVEg2eGfG29Ka/ZbpJC8i9Fbw7sF1Sy9E3CLR4W6yZyxyZ/mGd486nS2D/I
cugsAYBGPWnRx/rHNw05ybd0wRTWRWob2zGDYPyK6UE7DtIHzc5i4p3liwmJsIUP
WsRSmD052pwKA6O+C9aTC0kBeJPFifvl4AQaO4Go8q1Lkt+muJLvDeDbSM/VbesZ
tdtWyTS4A1dwBXxtYQc0moBmaj1V/sOoevffU8MFp+lh3IhrdJqqUiuwPTIYQKbk
6YdL4Q4n67/HybIkd2p1PqG0qVHIRwlGw5JykV3FiAaf3dTw9iP7objOyIRyS7Bw
CqwcDNr8tbeQ84FFhrPJ8A+lIBdGTFedVMCBDIQ1ibLGvw0qo0TMWuz3eLo9xfPb
GD0oj9pU4A66+0lNQkjozDSiJfTmlSOPQc3gmLIA1Ov7rO26SFegjgGONnoqbSuv
H0YE5UE7Vg0bN6ljvpFUDRbUk0apDJqxuLNaYeU6CwuzM4G9FsQNjLS0YUkL0prN
mJnTBsK7w1O6NwMuv7nGBQ/sFNCaFQx2BePBdtjmmmXHyxRbh+Xj981P9T23sO7u
SX8Uz0Smj969EZIv269c/yP2d3ylMQ277vo8v5DGJOpTaf2pBJPT2MnH7XxomfOC
oKitytySGmgQY075mNVNFeByqGhL/xHfMuFjZ8wRvuBrj2KJo7uKzQryz33kuLhr
MZRPiBrUy4yn63QD/tgHdiSXkOuhkf9WeDFE9w5Zj+MtgAJg3cfmyveX01+tzKQk
qfTYphKZIzZAD5JBL5WfeO15xa9VZIOMF9kMaR0VqWodugSNZIo0i/Nvq1M3VpdI
W6FFxluv8iWlTGy9AqdDeGpI3kJNi4D4RozYKl1vtQOLnT6uRY6zwE9D+3j+SdfT
TnwuTCSX+DVOz7coJEJuaOT1Mi5xJXO743yPDM3MAJCQaSDEvTVtxk0B+24mnujD
jlk7sYJR6auhoyttfqjkcf6IfoucZfHRgodKmw83mH5LGsc1Tg4XfxJSH0I4hBpv
+9i2esCvGAH3O5uWiU5OH48Od/rLcxTeO3Ynjq13YdENd5pTPKJ7jOuPqwCfnV7g
epThetpWouw2z2BNT4mOg5+bSSsd2u6d2f+7cGvz/cQx3Wt39yGezOAKBaLzxfr3
yd/SABw3NypiGXgO0d3sN2lJ42PjJnrmDsir/hXp4WqiEPyrFuAnr465Pr0ekN+Y
Gu4tMi4cL/fhhPc6LkVl34l7x5ooCVrU+ZeDz5hVqGFZVLQIvEzVG3HFUaz0er7J
R9IJlLpnc4ZaPt45COFmqsiy/1BcUL4Zn9N7Q1W5n2/v6oDTjTaPOApiS5qpOOS4
ne2XRZY+U8BeMQ7UX+ATX6YdiLzj6j6ZfrY0SgWQlI02Iq+VNRiQ2LTRa5xLw340
3Bs7h5J2ggVgUY1nSge8qPVTkagBkDgMOG8D/tzp3UVyyP5vTsp91el81KFEwqHj
SFa6heIeEBtLwdeCYeG8vpCeoGFB9PApCZDBF9XZWze1t1Jgy4sQgpX5PfccGLb1
LOdt9nDoKLGc3sdL6Z0mgJ10hUvWlE0kr2ZEfFcC8pcq4cGgDdEYs38vCUUwZZ6J
+MUtfqO3NQ2+9Ehnb4VXkQkLdLcJJXfAB/vwiTGFtMzNmPIZQN9prY82crMRQcf9
bu80pJ1Czv6sy4nEF/DcAP85UypkhWjNf5l/nM0cfqozv7j0gFLQVqWfBDL2pLlp
FONnjsSZwFeLh7SWCwi2pg6jjpjv91n16/1oFSn2sLLmgddNOB0GtGHJdmhUS0yN
Mruwb+Zem87Wwr6gV54eJaFY8hNNwhD53xm+VdfuzpHqTYcJR+DJTd4uENaTpJ3S
z8t/qqmu9SSeJqemQ16YzSZdWpRaBXmp8ojVx97d6cynBsfO9sScxN9jPikmmj3c
jalooxz+Gm1vvdDsdFLWi8CeM0YbKyh5N7z+OOIDJINUphEnds92LMsVtrsYFYqd
iShSiDtl47983yRaqaFCjhrM/bVweNSo43Na7eOPgkKm7Bg335fjUAp2hvBef9e+
OMOjX0BP9V3UEnC4J+h8t3t+44RTRhG+wAJiiXj5DIkwvBv0wc/ZMPCiC3duUppi
nNmoj961XvnLVcOB6MypZAYRm9KTH/WB5oE2AwLtm9NinOTrqcabn9Bu6pt63m8T
5rRZMBwIFZwt8QGndzpo/sP+5/1FzA+q59X3ccrAxuYKHqCDJOjlJX6NzZtmntWP
xeTU+LNTZf0zMOj88gcWkUGF3NRdBsa79MTb8mmOxI9URVjcKQ+G+mMUHgttOdcw
xOTqmeY+R+HDgRCN8uxgCKnqCsh8TENHMNM6IDUToJlvvvzgN2Rr52183j1PH4yD
JI5JlTjsqSsGo8OKQBW01cizFGTX3rhu8KPT9uTE6KmM1aRWi698hSjJdTvZpO78
Nb6A/yz4jPn1ystONOh7rfMtBM7103kTCOzhaxOMFwri0l90QtiHYEkYQt9BbV9y
fadk3lHqoAnb7a0qIfirVtc9ptmKGqCMyxJYKR6GqWOBARZEkqgQVhinUU1xskW6
kflUslHMLnwFVKZuEwb/8qgqq+rWlweCqQWuP+MsDlz8ILEY1yQrno0aW1rk2N1z
MPdKL/K7F2d11Ru3WcGx19Kg1XvY8QJNqFIBpOtwlNbCa3T638CS7mQViFotZWSZ
KFiIKWiA7kQij2Wym5kcnjzp/SvTHL1oxl8NZ1qdLpXRSxo4EwsUa+d80VlLq/g/
fC7+HvsMEborlU9YDqD+krALtxTdgSGxfO0OaF0a5HpDymX2gJhSUnsNwc3tugDg
hLbDRNwe9Onmi+p+p78ahgs4DjKNS4562m1L76p2AE/LbPEP9oJNiBEDkaorj+0y
W4HiW1efUIAlXH5Rl5qa1pQz+1cTWbuXXjFdDZ1AQh/emBk8p6vYSZzYeg6BMesl
HzuMMBVb1YHQCU7spr/T7vdfpMsRbLV7toRplDDm7e4CB2um3KkERXviGHBapfat
dstRfbnihMog/M3H7lbNKBJWgil6PS+u5ZXZ6Rd3OmB5iDV/Rsk5T+1OcX8AIOVq
SsvoEwGA13wQ/UwNgckhLgn02OmMifUD7X6Bhs9G3vEj/KmmNp7Fl6lZIe0taXAw
xE0i49hLiQEUvSVSmATGE54IyhZXNNr9uIJavlkjETZ5L1mrkGqwghKzk0V2u8sk
cIyIfsTmkV65ol9pF5INcSOp63ojcMPU0FkvePZ9CSHRU1IrLspKXBveNkB+RqTE
/7TLWFKSE/5/2bC8k1NU6zmIuOnLzm4/VxLfUoqKI6CZ8/vikigwuAtkSQK7NXxC
KvDXOqoAAkGts+lAwb02ZIVzHvwYJD5UboT2qUDHodeCUAuTfUjxN/VD7TGeNbMe
e8wwZbaKCc3iL6n6CnlOCyVef1sqWJHgqAZHAw3iq4KG8vAeqkfYoXViS7uonK1Q
Elov9ldsNbyH5v49tPWcJ4THShIU1kP8ewqvwNNNvNW4mLqRSB6JrUffNG1Dgfie
6ESZ1rvg3xoVF2zqDSevztc3bAwdZsdMiPQvO5HF6thXZ1RrtHjXnCSu6gZmWDKX
vJvXwDFdtXUqIxunDg8JsvspHW+cNPgX5YrgoXdumqUJdZNiZCQPRjbnx9/ttKnx
cbiNtedTQjWsIzgshYJtKUd7kOnNN/TFk/haL2TQwSS3cDsyPUVZbDErpytqXtQr
HGlTjXsoAfYqGPxbIF9BG4+SQGUkfL59wPG7CqEWJgmDaNZ7ontFn65cnjv+4cYI
rJ24UAyoRa0xQz1Eqrf8/04rKygroicpKHRjkH+ZI6ePDTCX8UDJuFrWzGhBLavV
zGFn7YqB+PyX8HbLt6Wy3R/aFW2PisFd7Wt/TV+ACkBrAhF1JRSGNIwkI9QCzuCo
vSFHv0spJkg45F1MT+MvDQDQygg0cW/MJQDTvRMxtgHFQO/gGug06oOtqISGDDtB
ax+tA2aSpIgS2c2O1SrcJU99g7F1xCHo8abPjU3nE3nr3/sAk33cJEqJfKeoiu3U
GqJ0n2yy4K86HaOPlLYNGWnT0zuWZoQXwNbWBPIjpHXmzaDhDjcd+FboLgKLPr7j
pSWHRkqy5QS0NmRXLfJgHyFZ7lHpB04qJydPiubwnQE2YG4a6PuqRzXusrL7U/O4
jRhKddtfqvIyfr82cqHSs3ncKk2s+h0eod044lOvmHAAKyLxTwpkmwmLTVIrqrBo
7eao9A6pQYO373K2iQ0Qi5qTVrwd5/MsyPgI9sdooAvMIWj3b+BbuzpD7OaKwu67
marBqUGqDVCNq7xQQyAwellSjAjdtOxkY2akEAS/o74BTzMySJhNoIuSmw5Xw7Jd
rdTQdMAh84Q5L2mDjod/n+OqlQlF6Ao9in+nPeU81A/mqfAh+BoRx6TlXiRSgPMs
3Wmy7tDwaraG6PJZ1dOq+mNqo1XCbuXyCTkMfYJBIuhUIvfMz4fpS81lAlJZU6yA
rlT5rfRltaU5kyKitD7h7TeQ+/25eogetz3Q/5sVVN22zwPf9GikrQoap/+Pja8Q
ZZ11D4HY+WthYYpcSGlaYChZQf+rHlsu7LjIjcc0VB9rnwJpChy8+RnLCsAET2dq
AGU+kKgmyzJ362mtOBhM3Yk35K/d9hqWTn3QFBgOSXGusSHzz+H6/Yqd+/eXNGo+
i1xtQWawTvOwXN8t33dSHB/dHgT5Z0ZtnENFseS47Klr9zQTM5PcseK4k5KW76Oj
zSiSaNm6KoKbQfofdH0pTmxEBovt+KkhQmqApEhnHja+5O/NuCmaa4urSXP4i67f
Ljwv4wPpFZX8F2aCtNVMQsFqVkEp08Inbe2zuqDvYY1mQhdSPUDczBV80pS09r26
vS2suGmWGG3Qrl4L4Uqu6TjZl4uL4hDF2lZs8DLH74zpx11EmwGpnFEkaPaz3sKN
njFWWga97JoFObHeq8jSD5BDpf7rrmPLbDznrLLbL6My+PwmjESxfRDMB0n+wZX4
apQmmIC+zFoCCWFqn0r6jAIPFGUb/hk+TsAdxQ98kWp6Rn7u1smZnUjsHBUreuPi
HA8/82AypOm4sphfPzg7LtyyDQ1NDI26SgrtULtLN0IblW8J38v7txPvPLEu7n5g
l34XWVAW4oc83UKtmbLdji6tvPRg4imyMlrmTc5exuYbBSF5PzY7gnWv++Hafutt
SmRgFajBgm4lTtjtjFoq+WZiIVaDrMimowYGzmAb6EoHDCpUjSCQXApT9elajwaz
wxRaFoMfU0OXNjCKUmfGOFyrUD6evisKlW1N5rNL34Wcwl8zR/ETupyAYldXBOaJ
B441Z9Rr1RZ00g/FNe+BrnEMiAA6qZfgn8PpJ+oqhqCaCY9sM184ZRMEwoTAQgZr
W5N/Jsj8No8tCxHwMzLi9dexTrm/5m33jxce7ZymA75lJtiF2nMTuDj7w76MCnBQ
gCVtiDZl4oKt+TOMXCg9dv1J148QkzRfeakXeBUmh2t1zVDk1fv+Aoy8JeAdOyWt
C6gGLULuQ7OPPFRSwkcyTgz2+0U7uxY0Oqco5Mv2cIe8jUXhwiXwulB8Bt4xG2d1
UjTl+m+GyE2Av69LeHKZ7hWBIjGTi2Fn0fDGLS1fDrsD6whFLarw75GAoXebvl5+
wcLjzu+DlGtFsObmqvoNYonvgII3OQBed4uGlz0YGX85GXL/1xsIKgMQlvdmo8c9
79BEKgH3FvKWHHg56CEqDnHC5DYhgCIL3vCfD2QTza+HKsMQFej6AyKFu9BPM8PC
ySpnOujYCtLTo3fjh9xiMRyJaqH40nAUxvcfCUOqkzg2DuyYeXNdfM2GXQWFsNr7
zuCwRDXEQH/ji/paNAFhDlVi37EM0hTd82TSks4rEce+5KICkxKkLta+yDcACcyp
NZpP7N8B1xt01N15inUU7EP4v4PNiemJZVfLcWAhOX+bKFwPvHS/Uhbo3Db7kebJ
Zg9YZs2TnohRhXgHqsVg+mXCL2E65y1cA0ynx63akhTZd0zkO89WQv5ixe8Kn46a
xSuwXydyDbLQQtKX/PrtOUOCG9waNNAxiDz/Vw62NTJnBBrDjRWgkLt/8jBuftxd
6nWISmdyVBLk44LUuWcAn7UP5XZxRnF1ejtRR3pknmjY+WqNe+VXQvKNsIbYj/fM
+YAg0lPyhVhT2suSX/mn+utU+CyfU23A1yeefvvLrV2IX/2RaPXLrJ2vLSoobsMS
VwJPLxQmkG+wRXhSWRWMGfKQCxMRXcmA7oTKw1U0anigsdv/rnbARFizG0lOOWrR
O+NHhdMNBXCnSNhLfIiu5VRLqP1kU5+OtjNDYAo2YGrFdKlXiQ8eOLwVmZJsThra
x2SLU+mpz1h8mraGFlYUI+imOMxwD+cBuXSQ/8FSFyv7ONp93jA7l2TFF8hyIBvL
9M1ButvVJ83M+BhVtOBqdTEdv8fg5lzMbaH2BMzMGfW7QjGrTJWlLbQXsAVuBvYj
1mkpPebmiiJ0ex1ZeLusa8ZI7q5sj3LlBVZsB2EpJBxUjaqb2SagoTE5kwY7j41e
zYthCoyRUOoneyfcIhQ10uw1bUxROnzzzwRtyAL1YwmFPr3yucA/suKPn1IXpGLy
HHGkrdaerEhL8bOC4wC8wci420Bps6oHSY51pzstdesBfI9oc9dBznD9Dr6LlgxF
ZUeKnGFWb4wjaLMOkkahP0Sr4JegUj3VehggQj29xg8HQcJri+gFVFyMx/AzotFf
kTsOUnKefhXbdqudt2CMw99rR0qpCJ+NfAYa5V0LkhkM6m5PKIU0tOjNsuKlpNts
BpCtrvuw0G536zLCCtrr4UU1zNwBlFLpv4fDPHbkfK6YgGd7IiCpNt/WIrHQ9b0Q
1uys1CGu+sHInxRtgCLGxyABQEBxhvHMixZ6z318Yk3s+MGj/wgnvqzBwPUdZwjH
bECsWgPgfz6VdARv6RYVRpcwAGWEyW/awkTfnwRdTc6IaEQ3nJFOGdpVFzmtnePD
qM9tq/CieqFFCjXTrVWeXMdxgv4oSyTnV72Tahq+ED4qKz9U2GDANYtBQFFFwTZX
uzBGGAm5p7ur/6oqGwcrY6jP/pc+kJaeuHgrvOzPvzcDSD7KiTtqiGKjT0WSs6ia
phCCHrNYdwjiLvVqroXzK5W2sUTA7D1gZyNswSnYk0H4G4q3NJi9Lm8dKPfRN408
wdOgbKdcRYAhKM1hhn6JEazkI/InCl9rz7UX/zYrCekblwCYE+nzxu1UIvJZeuWx
Y0rgFy3DGN7qIMoDxRNiVtFMbpYEn0UL/7JPcgnlxNviMHNbOJIwiJ8uKBn4Ertk
Rm7c0FL4E/FlcVC6wBUsKYCTIN1D528h0a2w/TGQGUZSnFgIckEPJWL1Wt31mdVt
16WsD4GgpTk4k2T+VXaqi44mkay14QGzQJQ/PJDTnKdGEHM4eq+nx+HqtsFeJwNc
1tNGsjdfYFcC1zu5VKylrj9Z8a9WSxC+peov5l7MpHUCGjsgCGvyX8Efn7C/Uj+N
Fb9IE2whVyQjwjO4M3TytGpJXvuuAM/jvhSnXrCKD99tbszq7c8JWMrPIeQ5exim
PAdVoF8mOoFiU/RwUmjhPHzcU+AbvvWdUiVW7Afr5UcPGFUBE2a7g3+wHUWK0I3W
IviudJR/Rk4MelcoGlXdcMuLdfcQOZDcW/Rz82vgGEhQQHH+omHoU8eas6Nbe/cV
bI5GohV5HrLJ1tL5H0caUfy4iq62eJ6nS5fFoQC2x+0ZYAzcnY9rXPSFsoPUwzf6
iCP7eWVGLVeZJ6kLuDfyljqNY+WkLEUUkUgV2wo8W4idn24eZXj7HU4OCGg+sPdR
K09u7dmvSC5hrtUkGHdnheihT4yjWhjoEb+86aGIo20Ce7ogYh9WpBN86fCgcJ3M
SlkK5wYWOSrnlb0OEzhR1QZPhKvqdsT9ElQJwOmDunBkJAqWaKETohP6V1fQ99dD
5P7W02u+PahFsIMWaufyDz5QgOXgmxW9kQ/GV9LR2QLgEQaDM0+NBvqmAnapugVm
UtdfWY3xIpOSYE2P/2W3dxVi6SRXBP8ThCnFNysYSwuy2xiaRb0HeYWvUqceBFZE
Nxk5e38hRj1eZ8SxYbXlD8oa5SXtgKCDmPUd1N7QDExSlp3grl89j4Sp8ynX/lUI
DmrEsjCnOwofU/wED2D/fHsqyXufdzQtXroCmsPatxaZ1jW1PqyQmsGvGz1QVE4O
Wjr7+bde00c85qMn7Cp/N5g6jqPjszB0I3+flAO2SagD/wA3eGfcbEKpICNAi90X
4SL3GM/34zOCxhvhdsbROCFjXzEkrgnBbjNfEZ5bAV0VqkmnW+POTA9t5wJf3bMf
JjhDqJkMxJW0LDULdlvgpnl+JkY81cZq4FOZXWjvN8cDHnyDYqraLjcA9sm24Mvk
Y6q89V9SGGX/q86CRpKIlQBUrZsIOdflAoBv+6icPB2Nlmfa/emeqG+Hpgf9J83L
Bu2HmULYE1qJMQmf0ZEwTJkakfQeAuhWs5U13SsT1HnK4WmOjDVglZesJkAz7Xy8
Q7tyFVnwvM0VSN3np4AtfqtZPQdTqswQVGV7H74vNGXoymQL9sxgCzlcwumlt2bb
n70D4r75DA0Oskg0zVpc5pYIi6tkTIdFEAf8iBdpjTKlPKiiSTcppehvEGplvxu0
ettoJN6UyAvoMuAIRUCdhEKy0csC+Sda8MF195vvBjkafItvp64ESjx5lpAQBUH0
HovTfLEEzAkrGet7e+sc2MA29/EjTl4krjZcJTnaIqzPBAgtIZsVTHYXPXLiqzyJ
2/EwK0B4Dolc3Lz646/9ODgucbRURHH1UyGb+42XndwxH4BCi6GDtA8oQivNPsBG
WPe2xWBkkz3wa5V45EhU8eJy5Q5/7wDz7TeURnNwAeX6r3MpMJnT18b6dLb1Zt0p
ElMaehUNsBwJM+K7ZtpNk/zCuUJL/RdeUx8b/vCZCpm/oP7f3sJ7pPElmx3m926z
QwGG/ysf28jFLxoHzWDlBqHe0sxc4QQO79F3pZuP4TPMfSNswV6Trg0DLfgCz8ZC
DbanSzCV2GIH/Ov/oZBM/75g258dVz9Ic9oJ32Mr0+O884wme1y4CF80Fmjsy0Vj
rZRG2UDbV9dmwkRckwV8ALyohtnfj4NU3K7wSpMDYHi66YPPhFrA457cCsi1f45d
RIeCU2FZUf2PM+Tg8VxeRHJWxL2EzuSusDVYxdj6G/QvuHwl16MMerGj674BXkYe
SPzdBPfAWOf+qa+spzjSHycSTZuiPm/iC6FwBMb7noIBo72Ng/q4pklVaoB2pYgE
1ANJGVEhwYHrAy5HlhAQIa67Q4ih+83zGXvTemcSlS4Qa93g1LyzpEAcgj1pxPt2
zddFiylIKSJtF3aZWnoFLuybZA+Vi07YicKWTfowQnfBYgKBZEwY0NU47EW/bIl6
aqyOcZ2KIClGtY5rk5dMJKVQqFZwYKKoHrUroy4toHU/LpCpSo5685cAD39ekGnX
JYE/2n9EjhfwIjtFZjBrgcs6zgxzPW7ikXZyCeS0HunbjHRs3QHqd6v2R6+S+rQL
5Eo21Op4Wobm2GLftcbEONavkyNaA2TUEAKC+BVIshuNe7qo3RjW2OJ2U9JFUWn6
x60HdIl8KmSblrevZ81v3QpjnfixwZ3rY8wzMGameneug0XUHvyPeoTG0nKgvUdu
ZScSizFJZu5ge5AXEwxNVojJ8+Velbz4yVct2wlpCy9eweszz3pQiE4+tyL+XO0j
h/nvmt/JO6bpgic64fbQyxKN0Wvw00nAqHsy+MkJ4vCtiP6EInX+LGtJLYVTr5CK
s3sKj2t3prml0JVtZjUfevcLPynQJtX+Th+PudPduX6GN5MXNPcBSUTx6f+hg32l
5P/VH4Ab2S55LbLb9Nl9R27kGfGK7F2Z1/4av733At6oX5qtHlP9IBEilE8WOBxW
KfSP6Fz1PeowPmeV0hRc8QRFwaijX+NC83leoAy0aY20aS7Si79UP5QGB85MgLfw
6xyIIQpD6CqUvAwYZgXNv+E7hG0PLnt6R+vZ202j1xke+hGsEaf7/Mwe+sPOrKSR
2CNZproDr/xi+V/tKsDH9fabluUf8WsWI3nI9SjXPTJzRRHDQfrTqKBV7oAb44D/
87BSn1jeyxAi5LL1HXg+14VOZufEv6V1SElv2mRz0T8SpU2bG2TP/xzCyw/UnZlK
SGB4NSm6GWLqmgDo/4WhWVSSsERsco3fRlzwUnWOslAJ7zCL8tjQ4Bx+LtJQ2PxX
mbe+Y/V4FTb4xAEkwVhsF+A/JdEpvW7HLp9g5rxnnrr+0ZzN+1i4+DI13G8OpW2Q
J4D1VFGmpfaWiecLJMILyPNXGECzaYOVqIJUO8LbHqhfPynzy2Cw91GuvJ59HbDK
BMLvXTrVKMpLDkmZCO6A65mMqqYaRemXWKPT+b7DsFPxF2rzpWgSx0F8IILhrsiM
Y5rGjgSBEUlh7WxSTGLEMmnXXdJCyvsFUqR2Cgqh+NYp0JEiGS1ZsXOjjsixHStN
6QI40ILM9AP13PDUWTTp6Estz4tdvgTc63uXQo+KXTbXp/6ux5FbZM6MYwPwlDH0
NghLgJNQ9bifAYSGk4J2w32TykIq1SshH97k6p6gCLpThmSwUScofHK++ABVyvpW
wx/3Obb003+0AymI18ZyyrKbvGYpX+Y8vIGqsG/jUJrRoaFLHEoxxSgKXGO+tsU+
24bXiBK0Qk6q15rZoZsUa6QF/4PH7vozHqVJL/r99hZpgBTIuJvTnL2yPQz+FGeM
0BT1V3E6M2bETSJdIDS6oDv1sQLtc5doQungjNoTpHbi3MvWkPhFZkZgMuz237kr
ulel+rnZkTBjDu2CYJW6i1Gp9fSbVM5h+HMgaEKp+zKXJKs1nllioSZTJ6YWqgm5
Osa8sfJ9S+42yZHW9HaenICQSEiZgzZYnphZdbKUIyiv7zC5h8zsmzjrlLVnmKPZ
oV47E6NNudF6Qxg5QGHk4CnVWwUkvb4M7eZO466XXWp2bbDkhSf//GrSDexTBuUO
x7RBblG/sRayT5TzBJbyj6qHmYafxIdpgkBT0s5O2Hl/QfZ3+5xbTPatK/6jcYFc
zyogQEciMqckzkmLmXNnhGuwodXOHD+A+vcSQa/sHxZNtkDvv18wL+81nymmSZeF
Qk8vYMEaTIa716Bw99ZwGhaXbmISJZUFPDFSIUqwtlj/qEdjDULSBFYkfeMtPcnK
jFh6SPa0QE2cMKZt3dMd7OPKEwzSV3oAVZYAReuyiZeNMYFIQhzG6W3pe++Ldfh3
e2AyQnkNxZkd6hD4zoPXexablsg6uKGtH+wBs63c18uwnR0TpfPxBeaTnEHBu3q0
F1xjYmrc/oPzwtXDk9yzuf+OmwA92jd2RQ1wgr4+zOR2+OynV2idmSlSDi3LrTph
wPAO1AArZqx+LHiAFMJoXPCgtGk1XlzTDNatRF0Oa65p0PbcV+qm2jOVzHRIXiWP
QCuY703bT2c50Od5RdWF64Hc0ac/SEaJyspVqspa0fQm/vlpfCd6dJ/E5G09gDyO
MYvRlKYtzzUfduY08iFy1jLThGvt6Po419ih4Fk1pjM9u30DlGNAP0u3kcYO2XrT
p02Sw6MGzkvFXIJwfq+mKILTUeDi4xDDNXG9DIbRpYmevCNL8dmxEdq/G1TEJ1mD
9kCX0ivSH+glkXlC3ignBA61TUcZ55PKTwMOAbvOEnB6bcU9yhF7vjcN4zgXLWm6
iQhRZPhf0CvXi5jD9WRIcWB7B4emY5D0hWSUULXbBd4aMBI9GPc9o8fJtEPOeB3W
7uKxuncwbODmNs0pTrFHvAbFGaz3N+gEYDKzPh+tFBxxjO3EQpOA9bS+TUtNZ7bV
o9H8OHLBhqku641EAimSHr+6nJq/qOMpodbFS5lonnKoQyYqA2HTuTz3UtxxJAR+
wixYimYOumxtAyHHoyp+eAa0xfyod1yE5uJyUqMBcO5VWjAJ5ESB2YNU1X/S0Rk2
BMwRps4ewHG0PmhajCy3gbpFesouAC6JQQRM+X+pvrw51khFPpz714b6i18lbXbb
jyavT76JNcc4sDbOtN27xEldTf31nenTHrcfkYC06Q6rky1JiYZyRELgsy+T3l44
xx+c/QYAF097VnxfSENfeppBw51vXbggKp2/wYCCqoUu31EO1/mssJeq+jof4de4
Nm90fMUfzrzbLSjgQlqOA6lkYqXN2SJeklIe2aQgQiw4dlTSiOhtcr6NDOQlgrIi
/Q8iuJ3gjCb5ZE4m/x2QW1vpvOYnAdOYfKjM8QihxwoTOcu4WKbQfa+DHyGuwF90
nTBx+x3VjI+bDyQoFPn/2197H5z0cJb551qt67axyT7CKqkVolcAGPjGHVpxpJhe
VV9MTn3LwVBegbu3Ki8bdGciHqWI8Z3qpmt0JA2g8q5Z2VK57S7qqQATEZ65Pyp/
isOzfCFfOtSqaBfhV0UIGSc4WL+ocUuqXl2gWZOre1N7jSLpX9Oq+0h/P8Ox3IUl
IsvvGQg4o/Vobhw9NvRfD0glKo3wVvAWBY+pa/gdvMf901Pi9soWHf9JARTvVWTz
YlriN1PS2QiIyevIpYmsMH01FKhp13T8c6sdv8/wc7ZY95gMU9CNgyQe4/uYVOj2
htY4fCnrp/Tr9Beq8WQ3rxkkXKtufZoVANJKC60wtLbvy/uKOmmqCHFVf2RZtpp0
4i+n3xeoVJutORjytvtE2omKGwiuDVorX7KesvzZPE/qZDBFfxn4PaUm4QpCEJQC
8/IwvWvU+gY/rN7NJNFmL4c8T4pWwfHTdmxVc1NWA5NGY7O2mghs3pcyJWrVIiPs
Bdb4afJveuX9WmzzJCJryD/HIjmkfGJvBESb7pFUCRNet9M0rWQhdZ/aLOYFX9TY
Ms36xjOJp3+hq7hNJRxekpJ2IHSX4dm1nf+z3uUUHnDJlP/QnqrGUA+P/lyUcEpO
Qf5kVyVIxLErK8mh2TsmnL7OcacpiMgEb+giH3GqLATjF2N/8sG5R9nyMr7w7lTQ
89NyvbP2TWw5X3/oakNsCqqnE7fiAhARFbRwoSaVhD6uqfK32knOrcIs4f6iM9LX
klKGLAjEnPJUtaw209goxKXmeK2WYbQ1nnuUCbujpLjNdGnFKG14Ydw/jUh1QEcC
cEskCyr5U4Vm775NK0w9QNt9UiHFJsmxIoo/prNVafn0w9Mj6UTILysaMINxtmFn
eVa5jNP8LKs8XPTr7vn/43wTKNUbct6VIsUnAJzVGuYUjYun2bIUtbOz3UxFsJlI
FEavJrkb8kjngUdouHxPSNtp1JbK8NHs+fOM9GQ/UB+WSxwxXhw0S0p1SKqUqM6E
ZsKH/OAXp0G+X5VTzd4eWxl6V1CJCmdhthAO2La1KslVQkBGh3wEJmOD9xlQLE7I
2FJEZNCQeo+ZAuYVVd/fclpko6vVMj/+Zavz0/+6E4YYGWrFd5wMVR1BLWbyJlvH
KbAhxBUTVpBlRq2DwBCKd9+1r0wb+MIW0y8YfCeLDhGClZQiti2Erimkb/HK8Cq6
9n9bjBVp++cIF6zTQoCnedCqrcXmmFdeUhvaHpUt2sT69XmwT+jVZZf70T0JvdDl
+UuBGBSV93x5QRsrR6+uF9xllIa5U3Q/z40iqR5N3kkB7J4d6jPG09RPmG34eTUP
dKA3wSwHar28Og9gDbPw4zj+CvIQuYLPytyM2aCs0F8AOCNVhrf6h6xpmdjSCgRJ
YKYFfLVUD9Qn8t9rsGR5jjLOb9I3qreOjjBXbNsDVWtbNyJzxsapbg2YLELGyBSl
dnOhkkqb5q5CDEsRIVB2KERj5n9omd7GZd1NuFlEu8AUvSoZCdu5xO0mjaZb/T3S
tuQ4YOKpJas5jC5UWPEUfOwJ2ryRuiTl7KgrwixYytyheGgIvIA+VLJCbUuR9NI8
BOBkGCctOB5LqL3gvuRfdhJEbICfseqABrKxiCJLmVlhNel7Vx2l04w8Rd8QsTEm
nBp7KVIjyXRbAFnuo0AQe7TrZNG7uV9kmO1rKFsusi3n5f9wQm4Io9RZHl1Jl472
IID8Gnl5x6tBClX0ftnMP/uYg6hU5nkyFzSXY36DX99bqo1ep3wVZ9MEl9sI/2E1
CC5N0B2DfwuMKxsD8CjJIzWhhFG2hJJD5IrHbLnwDqifmA0cH9adglqS2GjtNT3D
LuAsV/YxIV609onD6XSh0Xivs0XmCRLu2XteMhkcaRTqpSw9nN8eHUi4G/YjQHn+
4FxiiDQhMI0hZjV4UE6/xK8IUxBXIVP15RyKFc6/dMiOQslX5G9CyLXVHzkmHunW
hu/5wIrrQzn+bAp66M+DgIf/+L9sTO5JiMTo0DrKT6KMT4oztI6jniulzT8PlnmS
F/Cj+zK5d2HkTl1OScL4tXE5fcuhaZIgT0hBwAd6D3/Tg0I59Dn4oQhJqjUgWnyk
nqlVTCAwZy85iO0rALljDwl9wm9eIoLRS+eSjteVLSNM+RlwyActd9qxOSsTDxiH
ORVf9ENk89G6OXsOFWE7RwwC6M7rKWAYo3oOHtJ88Or/kveFb52RB/cllu58A7na
eM0o56UZCrodU1/AmQz0zzIDf6HiG3vQG2MHPzM60d8oWdgixhMTXFsui/msmGow
JWvDpFEoK9CpXO+RQukfZ98WbcpmzsCKQAtX0fZlxjmaRYirK8JxyNWCsLm+znjg
LIud33rVNYL5WRCG9cGSzJ1djKbok3bWg78hLyudb2IyCX6hyiDuTw4S1BdzN2CQ
U+AHe9tbjlTwW4Ts8afY/Vw60N9FARQRoU6Hfx50HNVccd41JyV1whEFp8V0DQXe
X8vYk7c+KiSiOYmSOkuw7DW8+kC+Zqqn2l8WEXa2QELm9WauUMnX/TFOK3vjDwLc
iIS6QRXJ0ZPO7RPr1vCqF7tRbLLH3quUmxT0wEy11jOzNjzIJQdGLkyCfLijRKyU
sMffx5Hu8CANqrgKcsyZQXEGvaQxElWkAPOsC/esYkK+7tSBo0viMECWtCD3GUtF
X12zfg39RhvoXEU7C8cfArgM6IZUtA4VJty+wTMtt25vmEfPTSEIOdJjwvWjwasC
AkUlB6Q6RjoZM4do1JnEpkgAaMIDpTE24j8Ie8PASCjJ52vzrX9HCTRVf1/4nyuR
dGXLpsH+DfzT7SpAJgXBfbdyeGCheeM1XMQs8l/flcGOxyhxGSOfQv+PLHUgL8Bx
0Ufst3qNDF1jSMFM+5cvf+g74Tjtbpmb6MzyLLlUT/8Yy3CfLdyPqh01sK+CiWTE
LdA+hREV8NViAssE4mGX1KBUpWQfYlwJSPiGx7KaYxKFlTuJ/VbNjhMZkEGzlzPF
8Yes6Aee1yz9ijCJlLb2gkq5YgmtMOQ5YAShFvL9B6RVOJTv44tJr8kglyeMac/Z
TRjSFZm6G8GEwxpzBsYaZzUMYcOp7HneFYpn/3Xf/k/PGteMkDfSxzQ8thoLwlHP
yBqWAgo415SDH7Gy/h20sRXCkh3lenMVytpO2EgUzVRwHlfWWt46LOYMiX83ZqHj
ODIe0rjX4VatbW6vpUpeXG0XN3n+JiapZCTT+aNNpUaOk5N9+cNt0oIyysY+3Fkl
HJ/fRKDkqiPw4OBYc+GY/XMWUcs1MzQ0/FL8NQtzlbjs0wMAu1gZIPaOY0TRYmq6
h9YuJY7F0Mur12zRhhKI1YjdIAVVNRuiC5lQwPz+v0JNLaQAA+TFyOJwZS5cuAPZ
7a7fRwh08ccM1N+kVXpHz0egxQHU3L79xgQVxaZeYMvyJ7pDucLQTLOp7Z+bTfnU
fadTfwxEw3ciyc7Ghs6sVx/887LFIH1FcEBJKA/eemz0p+aDpo5NRfroQVb1EKxB
TheYUb6UwqLALBG+M6orMYqX0UPlx06naLHFFDKcozGYE0b2lH9wBSIQKoFmhkYs
N/uj0YWmePAhXW1v3JElfQ8v/H2mRV5H/w+kkm/uMFoSZJDUIvR1YE2a8MzncwUu
w4UojgdClyIyyU7MXS4Tmcp0brNhkEnN8DmRuay/S8rQAfYsAnp5RLAOuv6yErLi
yRLCtChATjAoMR8KnmutRED+E/Qt42+pCJ7HIBh+jEpdlVN7en/RHXiWLJs3ulYJ
0cTPOpyOvDI+67CJQ/C0n5cEepymHNIkmCMCNA/aPaUUGWcZy2BquzIGvbW9ikdv
/5Oaqd1xvOckXWMSeYBDgJo4seKg7+NujxTA7P0ZO2LX59sAZnaupoXTbs4s8jDt
e+3xjZ3dP4vFr8YhFutNJW7WNh0QHHTE4i0VU5wRV1uv8QjvjiL3sWHJDCarJVmc
t4XEi+bmO9MZWbcz3+Zy0XJegIe9x4kZu2asPJO4/szlw7NNZ2S14JwzzIyrE1xE
VIRVcmUdboE2P5qGT+beXR8FCuwPVGyq/NAdR0NxyaXo/IAu4F0e0IoXHVdK41ZV
epPK74NOtdyM6IErXUbwqntd+hWVTqieytjn/idHbe6QmgReJBeGp4JQmXlufPkx
DCiKXwVRj05KKivjWuUQldgCRWvxnBaBwTKArR7EpjElwab602SZQ6ip7e6Lt0B6
Fvro28c7BmF6DDlPTxBsoHKnYuING0ZfahxzaI7KTtZZDfdhJoXj76Igp7YiRfHd
JEg5i9DeCwBzlQQpU5QZmDE8xGih7/rmVTrMOiIaK22iA0Eo+7gW5yaHD3XymnO/
cKwiGWjUdGMqaNCPOREPsow8ClxoHuOAkRJrI0i1Kyrpw3nP/e39aHngEK5f/pBw
w8/cIjX/BiOyRorE33DGWdYJRP8zBLBkbrX8ce1XsGEjDrE+WecPBDF0EJh+Gv9N
x7VddttdCAyx0Fp9Hj/6JKrb8cU651S4Lo+uA24b9nS/E/K6QqJl5P5gaxe+0xAa
v8nbF8tcgqyByu0bk7jW33+5ZLLbM0nqT297DuXHPBbdRpm94jYsGh+IOSd1CmtV
CkZDuoQ9DKJKlXGSJW6Z9KwP8PutwFGIuhuiKmvFXdk5yRKBzZi68EPUTKkicT4N
S6cp3tjs/4I67bJ19oYQJdR96DcaK28oM334t83W0NSnlOh2DvQjoNG655/IDFc5
kPT4XK6qew2QnAKs+fxqFrrJfPAltEFgmnOoiz5QyM6BZ9Ji4oXgIrxt7bBkvBuT
X2TNbbyFMLNT1tWoEYmJOQOI82S0q6MenTtkbJC5591fK89n7csi+sC+6wF5OiMK
13Cmi+H8r2Ep0GJKRBVSYDDY/mjZKjBbqwH4u89955Mefn8UBXYqlwlb36Yb6njl
dmYYUVP3amc5NHl30rwmeJihqSGMJNXWi3y4IKRTI8eg29SxALdqaylhfZMotA4H
NXHm3bdj3Qe8zDqx0VydtnaegdYotJpQAXcYqD67AmmaKnTm4WbtSW7y0SccSYbi
sfdiEZYaqU/NxLFJfGBwS0tvud3AQgnhGiM6rc8InnC9eZrb7mm3LUz9BPKB1WJq
6dcRHDZurvFbMlpb/oewOSj8N1saflGK2H6CyoybAkPrQ6B7aeTAhFPLPANjdVXw
ETKdzJW3HWtjI5MtII1h0qHr7L+g+KbtsQHCIlpK2mWZZYjZm7MM8ar8AQAROpXE
pkeoRGot7a1/kD+nfht9y7tzUshSmekVytJI5soteOG3cRc5Cf3wmWWrLB65g/8V
dZkQdaJBJkI41blKeHns5B0gShIFlG4orBPGvGZoCR6qxeIh0mrIHbNB6q8/nBJp
hRGGmwmidUZTJ9jvaeV029clN+R1b4i9bsJAyHL+v5pbrhoZYeerX5YrpJzxekkH
mCWGdpEdgBx3ZTrDUKnz1BgFizYpPl6Tpc+6AXrFgKE3fRgFjQu5qjCO5sgQ2fk3
y8hKUWDkYQ+AxLKg7p/0yAZGwjsDEeBZlbU/2I4VE8POHCrgOLtJgBP1fZys3zv8
g4CQBjGUnL2TG+Gh4sWDoyMvzBVrP00v+MRmDFqj+v/AtKwVLth8d7HNxwdWdQ9V
RK2O8KQTbmyCC574aVpToleiYTRC8mXpoLNgAPMLlBjdj3rsCDuqUaeN9RrxwT5p
bHJz0xT9GRa3bTdPFJ7fZmEajFF+uz9bIHj5KYoW8M8tCahZd/x8KAvF73/OFxJq
p7p4G6D8wtDTTccD9FEAezzualTLRRXWCHQ/tG0V7vkuNTWEf2RRZ+6QtTKlUKq6
K3AhLqT7qY/zv+fvjmcY2EcfiQMFtMnQx+UFNeT2hT9I5tAADVBeIufAmoV4crwU
ab8jiCLkcSuE4m/cWoUiV/eHiaOUuM+7+vEKI89D2xIfyPJ1KZIFZzRWQ/ZJq76i
yXWkRtjEAuRdfMRKn2aTTdUKNYrMq2IwuFnivWEeX7wPaTuXpYHaJkXyTgYlvD7z
v0QFXEJoDZfNuiKm1ycxFyV9CzLpx8Ox4BoSawnJH5YAFif6U5Oq4rQ4z4LdMRyN
SBujD3FwSh5nxmoPI1x1861hMQ2H/3lbOlo5d1m8UouXXcOEkSF2eJOWXyRtl5Cy
0cqT2conEiIPhT1ocEL9gmrTCLbDdISKjJ4CVryXexcdiqbLXWeNvQfbunmK9iuD
ppSiXvNXJQFSAcWJ+1eCGVhmI5dGkhWhlYiZWW5/Q/EEWc7jkX6zWkNgsbf4C3Qb
lyAUuDRQflysTlp+kgxk9ZoqD6vKiXpUM0245RMRQPOwPCviBnb8c9J7pejjX2eU
z/hsEYCatU4hv86VOFvJg/mYAB4xKBpHVbvsNFp9ZcnyKqhk0G0TikqWF7/UEE4g
alfFD0KSYK8vtdfjQCFgfSLLMBMxFbF+XHEPypF+moKiFjRPb34uQ9sgWDQXQhCN
/v2S5HervKqsg8C67ZqXSIteNRVnhV6k+lWLAXJ/5sWRp6lJwuPey9XiXcsL/EJ4
9g0+8piVN0d/LNpu3HHzTfCwkmGjD+Q6Qdwral/HLOIJ1aMMJNyt9G3wRnDWT53S
RWKzjeNs3ZE9RK2s9tVAmOxn3iNSdFEd25Js72+591bxKmUL6UvuDze7tcMcvnY8
WiTyJGAw5yHDfgPfYEmkBS9WDnh4zeVReh3+8qNr/zTb6cE74o5upFKggaBre/of
Ciqi2AbQIoXMs89yw4RsGoJJgrggh7BrdfWgVbxTjI0Ro6qziOI2lrRt6gH0b7Ks
HTSsXrM1tNOO7YGaCJurlK0XKRVkYwka2OTKlyka6Xetjp2/NU8fMAeXdj5O7i6j
4ELLDzuHAODk8lJRoUq94S/B8Podr3IMSYrt/rmkMuzsKRZG6zKo1IajDzebl3k0
eD8B/7IRh+aeL0FdABpJLioPktyZpoE5UDSCIpB5KrYUdU+2MKF2caCqRvAdZcW5
FIs7XkcOBy/sg0e+4YLOTMf9ePJMufmmSPRT3jlueXDrN7TH7LduSjLTUpKEMdz5
gu+FKcXsgNxWzDDu5kmzbYrrUvk9my6cIg148tXNm17YhGBEMpu6taQ2KRKKD8w6
EyK+LGgS5h7iE72KnOaJYoaeLr/KAK0f45j0VpscqNLXzPSW9in3NbZ1pEFp5Dei
yhVtfrnBvZJTgXlmo1avdRHrbIGv+PMDSOiZ8+u77MpEWRszNd4l2L8LZ6hIcDrc
rLnG343+MlHMwTFvNFxXe0thvHj2eg1iccGMCl3OOrhui1Q92UL5Sm8M+oG1GaTE
96O9EIA9Dggh1xUpUjA17kEjrV9rBQVzP9U0XspzLBHIqBBP5LctL1GgO9gNbMb0
O+ljDvcN5gUSglPvy9ZqGxLKF9bX06XK1oOTyPLf5NSElx1fu8u37IzXjt46hoeU
y90XSZnD8NdoBF/qCQ2x6L2WLVIREfgX2tlR8kjiCmWlIFbc0APK0wrkZHAt5KbQ
iJu/IrUkVBjAugSgaMv5SB2IY1z/hX712AoglFMpFani1BkZubPtweDL0Os4PApb
x1ftCRSvzTCUUgjIMhGXRbZX/7mNRRtRm+Yz2OY3UFUrk80i/+0QY+NOiWhLpZe7
ZXzdtVQgdsZCcKBN46+/qodUBuM8UXFBAEb2rfE/H/xfeqQNvh8XExiUQEGu5Kb7
KHbQz7YmquNOwB29xUaYsNLRvOiyR0SscAXY2E2uNiIAMHy5gzfFuUBHXTs4Awf7
RMDVmB/XKG16RkgNca0eOgJL4ra8XzhB70tywLIMtGk2slVK7tZgS9coHCpklDWn
ca/BVWBL4NuZBbdyH8Q3PFtBEhWx666lGSg9JfnyhVYimHps5P8vmUbrBQ+3fPBi
2jalN+Mkw+RxX5LrRqQ3c7DIAfzAREusnMokelABCWFBeEZSIPYshHL06ljuHpgq
nbPqaokMu+5CbSeyPg/bOi0Gn5ym5JvF4aiuOr79mIVro240vxBj/6Is78Kk0ymD
rrtgeHRmYJqVikxEpBzHfcmXv97weoVHw7IJ0Yr3V2+K0FPKP3zhEbZcRw6sAp2f
usYYP/I7e2lxGciY2o7I7cwESrKd4d5tCXnMjDls9MCQaw6HvSZ46vgDG0AjvdYi
fUqj00QFoDw4GM45qBsNItDJYcatIsQ/f0tQQAZEulgqvsF/doxJnLdY3uTXbd5H
8wg4cFqUnPYBYW5Jrv76d00PgviRxyEfkh6tkwO42jK5W62sp1FbOg5IF5axK78W
PTZ+j4OHs4VMswWyz/YjuZaXMIkpqvEqpcM3l36oLp2MVE5TID+uTBwq1I6ww/W9
mXZXln0B4Dj/DEFM+ODBhbpFWjkWPCVawBIb44xgU65YUmgZgoTRvBaCVKHKzaU7
9yl6zoivOqLu8Ol9e2eFiBjoo131te9LBPK2YiOdpPs1U6HqoREnIfvWL1nZqgDf
5vQzkwVgHME9nBMvQCV9+vzSv9sk96L7vCAqqghc+DZotSo3bphp9dTynCC4GWs4
aI+u0HWxs/MXFeBzaQunSmMKgZued7z0DKoZcy12HP34rwR8xIKwinEO3utg1MHi
jrvqkk2CsLDrzBKDm+3tShUq5zHio+802DKmlnjVttusmqyO92PrciyfePiVgat1
yWevVLYn3J0EdAMWQyid7VzwFk+QlvM4t9K0mjoR4PLgaG9lsquGa3APZD/LgtdD
gtitUVtqqq6P0su6TEZGa6tEQdx5tVPefdZodOYpYJLKzRaoXKZ0R6k+At/zcK/v
d+MdWm/WzbNFwgDUmpvmZ+ugPC9nshMhTw+RUdwrJerBV/KCI+0SgrJHFziAG/ij
dTonRknlZZq9Jzu551tTE4NWxEttEHTguF+4cABJ/COvzefIEdaSqHbEGqxv4B4y
8MmWD8qxueOnpPksgbFmhMoRG8NSyeVRBIw5W2Li/twTbvDXU7k0vng4JIG/3dLf
+gpeDr5yr5gOVDCKNfVT0/D0vErwE0sk3d8Jkc9Y4iB1kWvC+POqw5Dr/wCVCaN5
e3UTFCFfeKTdM2oPRhZ0Jthx1s7hSzEpP7i+yT5yMrz6We+7H3NgqHAIwjRmL605
25UujT7jT7PCKe4tSDVhSwpv/SceGFMvjud0FGECVFtT5K0MP3eI419BFY4QoTVo
ZEP9yhzREQVrO42ln+XRoDdXOeQKN4bynJN0cranQljRO56gqlMYTJSrRouXabv7
LWCSB4r5oyrlCoYabYg4Lb7stV7HCf14OAfZWeEb8VbebVYip82KJ8XOjCxQWM9P
ukPNR6Gn9dgMDGGCNeDVdZ+KaH90Ouxljrt5LYzOvY/LxxUAcvD5fgq1aCH5KMtW
JkY71gpNznVUINg3EvVPQQgALrFhk5xpFwDCR9luQvrNZ+CSmTN7xBN3xXs52VTm
xMwtFLXK14sChWfeg2x5GOxLEXMHgT5dDT2ofbW9AlgWzx5XV8rWwEicz/rF/Z/C
wvUEXSVglhJVcUoIb0UNNJBlD0APtotbfrISq5imnuuHtTGNcv36tJjryKXX7Ut1
2gEmRqf+Iqhi5usB2MxtwnpdD1hJX9LDDyIjqDNKtDgS7x7767NLwrjmPllBOgBx
K85sDQ4HzAqDqX72mXafIwGIHRm4f/5A0huLGJzmitdfl206SHlFcGsq18T8s2qB
lEkgNa5gkcZnp1zeYK1g/xUZlNkN2VBVbyuCdep17/ntdQ/w3iHgWhUjQ59vAqbn
82O7WFEERkV44P/qNf83b7dc98JuTPkerCRUxKeCOWSUChfTl4c9WJBY8mg65T4r
uq+EFay/Er1pxKxbQYq9vjtxMQrmlpzmV7y6CZhAp4oKHEEzUYpo599JkmLkiwx8
azI2lkdB+l2Kzlh2mIHlNIYTmOl0GtVwwnplD3YX+DPVju2i8bMAdfIgYuzv4C4j
MahaXg6BZiBTwXA6VGhPNUHnGyQDHIx3629tT4EP8w3IgIfOzMZUb42CraYTuCJx
OwadHlDzlM6bwlmW8QmctqRfQeHWZ+CPNse3wH2YBRFPJOEh4EK/4K+k34jXHaNb
1EjdATeWV8POiF/TBn1k/fOjAtMTMfV2b+BbSWf+T1HI+fA1HoA+1xzKf5N3rpSh
RbWq4KzHfFRmfRdOfFRRQq818ICZqbYt/mEy57aEaqJy5fZ+YsErk+M4/DHIoMPJ
6WdPbJZZmNqTkKDuee5RZTmjRfgPLqZhf61t8ixIq9HXY4/M6aW39BysoVh2bmS6
1m73s3Zcj5bfmbYDR2vKxfyxDRUfZ9k9vYVx0wwajR0Ov5aA60Nf3guhZPbcUeeK
wM1psbvxkfMbF6erg/bOek24loTFsLxiS1MskObTkacoHYTZubJ4Xy4rsSKJjORb
FKsaxbHGoRIxR04btJIVO3m8trLurspnQMgNvYCWYQmj4FxDQey3sUSOBWD3HReh
AM6ZSByv4oKx/p+RlQlomT+MtWHBZg4gqRGvSMrePas0HgR30Z86OfBF9tTuvI5j
7c2GDJB61w81qmY1+Av4dbzrLb9kjT4O1zomoqX+bNTNE/l++LA2YNILDcXh9oAv
cC00FI4ZHKWey4HlhtoQYu+iz4cblt0TAjFujfOeHboPG8aZ5jxitrG79jylVGJn
I+4vcXzrWcIGjIh2HAn7BSNvyvfFQv7mTb8Lsn6Y0IhChpZiw2KMuTgKiKfiVBMQ
GSlEuE0ROt+vtUiMJcWB1rqyEBue6ufhgUGCkuPPu0eJwL+c1VRhO93cKA4xyTHV
a2zbWSPYTTMRcDMJ3zKk6mi4GNVNKWbN5HFmBFsYupAxF/XRFILSCjv8sBZAPuh+
T7M5r3/WrlGmUzJGUGJwtSceCmobxlHxSPSEQ+5zot9T90V2wpHyIrGhmrjF4dID
eEP3ennJg95ISomao8t77JtAxfxfTiXBXf18JWGIm8egXiP1gcm7T8rmH+ttM7D3
Ml5f7k2f8GUXyWKdKt7g+P2TnRGRy25moHcHDTmUD51u50LKNPHXc56RSC/YlFZN
ahY2ofk/+CY/3Hv5dDN5EiTh15dFxGCmeve9XcG7wcBap/9DTKbR2AP3p6UOfICJ
uXprx9hDEhRWsHO+f/2d+wSs02qqo0Ig0Ok5Nz1iK52YT4EQLPjgPGKIQF22KtBf
f/AZCQAXzyOfd54kOHS77A7AxYeFjcd85B2p4JuW9MJWUEzujxBFtgdQmPDxbjzT
TBmzRQo6mJ75Yc8WWbqClYnnmqp1L8qDbB1lMCgAtC6ldb0zNt6UNwPa7ScL4A4D
yiL8DeG+jUMYuOWefohjCmCq6p2ewthZZoWxD1mm3MX7KJRtqUhnavqmytjrWbO3
SCN+TB+3ydC//DnraUxPZsd4gnoIXFSiNQ98703yFV3veSRVWSfL2HaW1EjjAbxn
haLx6gzTbDKC+xaAfYi2h0MrVblR+WpUh/5rWGiNt7uXHJlL5QO3PexL3jX1daT3
Mq/uM0nmrQZkYB/RZLi1QtGUZkKHU2ycmteVQJM2mlgEih/Dhpd3kzOjrVNXtEC+
7wbJZw47R3dAf7Cn0rPesp546Rm4owRSUf9o/7srvO2m+oh3MX1hnAbT76jFmb2t
7hlRdR/Z38VI5J+JRsdyhGMwyRa6bb6MT3ovDrepNYpiG1nhLl80jIRJR93bvV4d
xb61tvLqK1tD4JSch4rQnC2DyMQPPf6v5un3mNWou0wTTEyumPovNXJdjYRVVDCF
ypjUftMoCcLmlwcoMn+CUzSWpzFXEZrf6jPJhlQDH0Rasgmz30dcxMXKgkPUCpIg
rtjqyyBdbrb4e8ujyvm4HDPO0V3pZZh+C5Os1UFaFoIt8+ZlXk00qMcOZ/rly0wJ
IoQN/GslBqo6+Kn681LNzUSY1JDtM0cdq5v5o67Sui2Ze1l/JH4eDWl9vIjQ7aI1
40TplOMosGMjTQe5Z/cS8H+LEM9tjufV+CCYCYyAtGf//hwNFWmaanApfr3qvJ2p
CSjV+hMQNwQ8YdUDGXfNl/e+QHwglnEPqFoVL6a4dbW6bGKkWqQgjXiYVfKaL2aV
SVY7UpEMwCXgbhTCMLM1lI3cwWFFaG2JXlCQDxihT8mOJhLOS+Sb8beWKKMxIEJn
lRmOitwqztKAjv4f7lCqtFj4UQayyZpBl09Lx4SJDYkOx0qMyIWE8Cc74j7Y6y91
06XDsyIyQM4ZLbeZwep+BSC2trA80kDs1queARCPanPbtc45SQbg/Mll0yfuz5FG
xSIEE2t/egNPEIg2SXBuyMyqOePYYvV+phqDRySgLHnf4NZIwXbC+cvYjblGZfkZ
Y0yI0jSIqc5S3M39pATXpt+etCi2S5Llvq6p9hl0gC7yGP95dTeek3uA5F1RKdUY
vfs7KmIaFSIqeegV5p5r8owHkQ6TpfPtxZw4kkCv1ipYTEWPSd/URuQg2zrB3yga
u0IxPkxhcxrbVXTROIPzdmaLL8ZqMz2v9QYIiCl6K4RYgx9tfmk0VffJJFIlqRO4
6ddOjdLfxwZnXnaEfaCpPvAt7oJ6f+QccjeW2y7l7oLV2I0Y4qXqzknTFTIYliIw
YJc/IBKJpsjItgT3nXsZxkNaCZpxwYE6ZS7qWgo6NHtI8Muc4FIzGpRB96LEO2tF
TmQ3ynmHw7iquuV1H7mBQur2aSr6V7s5YaxNGaksHDxP0xXGIErV53h6XNfrTBIj
UQIh6GAuGGerr6GMElc6ETpr/ELlIVuxKLMHDuX9iTHCwMD4fz6UCteWTtqXEt9I
q7kkOCqsvJXJiThkj3fjcooIQKUkS8P1ecDd1hIshEifhdhugBqnlEh7oD+WYoQB
uBBGHJyS3InhXFRSgLMHaq/z5NQx3K3VkJKqncYU2LniSM66NKZMIOBz6NtyZa5C
pjmF9LPmsGkJunettr7Mk/9DUeCubgx/8bjQz9XpdBziHayKm+rzDpqcLqO8nR30
z3399u5kc72krl06GHrsS89i4+p0kAbjvsix5cIbp12pmcZbJ1bhKxWl8dbS6F/a
YgfzNsYc6P0rDgst880vZZ7fGPqkKKI1zXcBBzKT1NpkGD6zOn1s0mor3P0kYq1J
4iM7ZeyOeVDbbRAR2amNB/cVk5zJ4tYzpHFvctmt4TIIAF8a3vs6O5a8STajrEtF
a0L5LJ+Q+tf7eboECmD16wc4dL1HHjyH0He51rWIVwXKO/N45C3qoBxxuVeXmvVn
vUWeluwIR200O73vjMcuUiPhBWEPfNlcfsdhkTLImTt1KpUBdu3KFWaVt2hMTl0I
mpFEgVKmBw9StfsZekudWyWVek45OPEd5bTklye063foqpHztS5Czo2v0NMRB5yp
xCJ6sDVyUIBs52fgHRMN3lOxoPTIBrkSscUFVEtX4z+eb8qV5KF28nT/zYqSVdsb
tHAi7xYtPX/bnRap4brPBdW/9x2BdpEa4nHfM6UDLWuFchLoWg6ldxrFy+QxwFns
rcDhMxYbykSUaxCA6gnApGl9J5NQvyzKtzE9e4GuUhziOmTKksduZ7ZJ5PURFutI
EUXubuHqUMKFSd7zKlowOP7Q0uzwnXBylskioAyggpolCQsQU7dfstLrW2S2V/8N
7jvPXd870AwuzdxjF4h1CvBnZi7KhcTfVNP7rsfr8OmGmzGjNk5Y2HxPCLPGhn3K
/s9RLrtVrVUR/bzT01/J9CwjRXDGZBff703MvTOUcxvRTl/IPGUAo6ZQIlBT0YrI
DsPzkfRSt5hI+yhG7Z42rY4ZSrrqrD7XYadOj8eDcOtZtgR25jwQC+sYAIBSPeNv
SPTYF2w2OrJmDpOZ/E2DexZ49q2bGOxz2bouB40yLxP332djDYW17A15RNJDAwy0
VOAjK7yifJPGu7KCfzzj+Pk2vkhdnH++BdiNzRW5jQYSW20d+d0qHW/Jo9fg7TU8
DKCQ/I41gh3fPVUQdOXBpHahiBzJpABhoL+MC0vJOUkPwaH1nJ8PEWLCii+GfTwE
BT51x3OoRTXz2lOSbp9HcncD5gVW86kbpkS7Jh6xZPDnMy/GcJVwK1m63bQdk4HI
ETaxCNFOjXCgImUHw7gan39MB9aSwIVRxfeIptGkj/L912vhQmRoLuXdInYPntLP
wDThA0hue+ejrBs70Xwg8COlv5TyHjQ/OkI4vVmmHhShNNBxqsNOm7gG5wlaMCtI
rO2z2vw/LxmeDL+WoZBxB4HOeQp3ZTObVig32eFslKVGIEMFqGMgc4GgXIyfGu4z
Vk7eX5+WLW3bfxQL08TydvYkU0oPRA5AojqPCu2WR1F6fgs/X3sEzXZHS4huuY3S
AUhys/bcxErle1Ucnd54SFlc7YzbDGBkMAYtCYgEKdvgUzbDlujaK56RD1lMZqaN
o60sV7YzNg05HPzcfMbbNP2yD6fawnpiEe38gTlhFR/Vk7Vh2+TDz40tsd6N/tVv
cTL1EE3WaYUMdPECeMdaoRWSVaNLJlDdUh4OvSyeSRXIa2fT75A0qjPm4byzwpNQ
oRz/5sQcqWNR5ZPoqCgnkcQNhd02514aZ/NlKE8SAg3mrvbcb2GJal86QK9Otm16
yE7XVI3uUqtIsgqs1Bm2Pi98dUzhcjPsw0SIjzQi9ExNdMoxk/2ZXbg0EDGkm0cL
7+OU+b1bCkErHb+6TX5yNYnoW3VG3XS3DromZx9fOUsolPTop+KCKT1TMFxKXOG6
9PsG3Tzh5FJXfjucwEUnIUoGPBQs8tlJgh/K8aWMt5XyhAQ/cwB1PbsWfYLZAeT/
yhkqSq57Vj0kMyBtjxJEqGAklMtoIHjHCXcqYus1fsA5ZW+Dn03x5ncVFfFrvkVW
smAYBsZuiHFi408NHuyJKG7rxyY/jtlXQeiEJKGWwoJmGK0oVrYm3TA5KuUsucra
wjX6ioW3XQR6gJNUCs249eBkizokkw+5SIU6ddte7O6bjj4dUmhspKUbXA32QOWq
4LbxeTSr9XxI4rZjhNogzxSdaJhmz5PrShUpnDDMMzIj+8KoLNTum0HhBpXdO0sz
v7/B1sxFhvLc6TpAzaKx4j8PqjUOXalF8T66R2kF4naDmzdUDh0IDTxfPO25pYJj
TZx13or43ps7IDP/ckoQue5t+vcuxb/1nMTsXJ00cBMDx8XmznwUtdknozMj7QDA
f1IxrBKvIkuCyDznRD5cas6i+ZEJNG3T4FUlaqEyW69TaDfc6Wm2wRjR9iFledsj
Ps60qa9w1sRpWzgNxFb2zgZuwFGNoL5PlsQiENFG7Q4db8lE8Se1MYI0nTANDfUB
JUEvWF3M1PAruc40koWSS/uPgElyLEioPfD29YCq0MdLwqDO98NrFGerZIPEoOoB
xhU7R7F7bv+cHeH3UKsMxqW990xgdaW+6npycdW39YcUp166ZvVRsCoogXNOY4Hs
8hWzOGJkxpTKPVjlSp/3cYnMtarxTufU4vKaC+jrwktEf45rn2jVfdIF9GbSpzc0
CRwkExROK2FemPbvNKHpb/DqgrHecFDI3GT5Kt18unU+nGAtEH5eBlqFYGSi/ALt
WAoGi91W2fJdIwAQv58unz5jdfjGn6/rCLI75W2OB7sjJSOXf8zJUVvE17ifvuKd
DuhOcUnjq3h3YN5LfzeUvozqg4x3Ro+QOPQ6BiFNdbWKAet7SUafp6SEkQdqaN+l
f4lDmVaZHaJdmYEPpkxmvgqU+qlFNdsiYONYEukfLE23NQKtyyfTYmU8H3xPJb5S
hoYRzpBSE7r3Q9xbdTbWUtGWR6tJ9L8p9taCpYw/FyiGn2ADpC5lPSbS/AFNoW7I
ZfMS+i2irHwzlFGsWaMVWwb9kcUdV8/bW2Ts7MwFjoR4mAlyCbeJ+wdiVEEBkb8V
o1GGfD/VgGAVA2gvGDNAlyY1Tmk0txJn54yIMEo1MYKx8jltV9pVut37qqn0vxPX
xm2P9zr6812ky5BxGBHwhuYPWFvmXqCinvv/gQC5TNsKrEZwusDWQca7XgeJf7Gi
V2Prxi7borEHlDmFup17v2zl3AVfAzYbTmKUIRgSrwKWJDjVOQ2qJJ3zJuAtLz8T
v/1tddpPISapYCkF58dd6zu1Ds2yFQlCrOfL6UptI2AU7H7VKbBaXVHXqCJME0n/
mIWuhFRrJTfVfhsheUgxLbkFmK+JSfI3b3iVNudsm+AFo22LkNPuZHOIRCkq74+u
j57jsb+L+7+O+QqHub5C0SX1/PT6ww9B6fPSG2/w4eNKBIFLb//8H0BWU9rR3EdZ
zjyL9uyHuI3nlHpdW9rRbJBzeyRUq9DWOTAPe6vc0IoOZRqTrPm+uPYVz5XXTnVe
r3SHw8K+VxoO0AMYFUt6HJ/EF//PuqE+cYX2XWQl1NOpSvvJagzGB4NA3FZrxCPw
FTLay/tcSL3EWSlbLvuaCMnG+Awphj/PjojMApsRSa6snkdA/OF7H3MW62S1+ZtN
fYJ7tn9ZAY5gO5/myYA14W5JN3sq0wME5rfPyfoMMB/blYrXeWWybq6L+5HKM7sR
gB5IDtSs9bGvOeX3nMD8bxBZ9BifHAoBTNp3uUdX4MPxGEk+ATSk5qaGw1PtJQ0t
vz7+quzpuoHjJxTGdHsJEHZbmiKbfcvkBP2fp0JtWKFWD0XdXmjFA2T38KQpNkLX
H5zIhSp42vUErOKk3A0GMARSMA09C15RAlGl6eiTt0vKgTX8XGa5l6YFNAh8r/0Z
CrYXIFxZHTXveJO4o4YIpc//+xju10RLq39pMRnB7pJZuJXNWdxZ8BrJ2ptDp/p7
vEF6EhGtl8nlER+BCUv4roCuAUIl824xiv1ivKUpse4nq9lZrrhBNoWzJJqYSH6d
o/lxjq5px/giGkxnDplAvfPzpmY/Y9RmmV7siG7/gbZzy3/8zermNBW2eDPgjeSE
Nn9LyQ/sg/beVcCw1y61tsr8a1+Mva9G6lqgfCTOazVKJidcwaIC4Wbqg6V/0f+6
J60J9S5dn/MDY5m3imPVO4RHaPcEIOYcuXAF7Hb+ufF4PpABk9t4CB4HNS3VuYjq
r0GSnE+YsqfQYLzAog/ch2RsO9uGJBixK/JnkCK4AtSkMK0gPVAbCb0Z8GDYbLv3
iY/8dI7JYn0EQMQLGJfAGxpS6UQB5EEuOEQ0gCgTWjUSctqPSFSZ5jQ0bI1QuXjX
yK+LfjYi5ob92y4umSqAs5x+YCoI+xJX1UUxPTPk2GPlIN1ZzUWzQ/at+0tm8/Ob
2iPvvGEMnhaD9jTaxP/YIGsY+4Mso4+qjDf/GW2dZAgz5/7BTu0KtdoKVHNgKYc1
v6PcaAzVFwP9fWjt6Rh/JfiIQWzkGjf5yU8r9gjAwZ++Y105N1e9mihDeUf44BdM
BrLOZ9LKACRPRKgCzTrQeNuuJ1H6JfMWnOuLCtJplLxmP/GKQvHKu0/CVVc8Pi+q
C22cZ010yLzc1OEwguVGMiVUrg6j+emKCPhT2+3PIonk2mCXhVIOthsOD9FSkMjf
KrGtG0F6RjlJcDZ3Q1xYdQ/MoE1ALlXqJNPZaUaCsdhhVP1SWGCxzwn1UFrFfeJT
zf/uTRkdOP8MqEGAMiHZyqmJb6Uns7MhR/0L7BIIQudEWqOePaTxi6n5RR7+1KJc
CpoxHch4LK5EadDUGxUL5Uut3mEa1kPQrceqEc/2pqXjo2FNUb8l1Ohw9uzA6edo
xt1FyH/t8wPaRHF3gMTKjFS9UG3BTgd2zLIwxX3S1oTkuv/fB0RPLcYuQXgUDKaO
z+KQliYex3Tap44VPnfNb5z3IraMSVfuGhmZuFPLhlH8erNHx8yOQ1C4s+dz+fmU
UPVqCaC6c7YBlXPuKoQRdXOZPnrCy7fTpNfW7X57Jrf90jZlZhYlZqFrl/JdLnz1
QvRqUtUHHx3MOJ60YmyIJ1iz5g4iBaoWxfVcuYxfz/0Ac7X3PiZLPcXAf9BZB5bG
wQbv3QwVF3zoopecLNT34tyodfjlB+i3mXC9dcNsEAIIG0EmFxWLEHlvrgytsmTZ
Yq6nhEHrwIjpwWEtNydckAaCdtVQHgP6d4/9mW1MwzkqaO8Qj9tJzz1fV1mDyuQz
6UhTT4mdnAW8ReHuVFcAv+r7tmX67B3FvHujUEIn+jA6jeEWssdLhgbxKh0+ynw4
bRMa1PE3tvkJ1YNHP2IxF3Ym0j7NH5IJcNNcdZ6ZX6Lvky1jKFMxWmuPrT2WASE/
lmDqJDI+mqMz9K4+pxN705fMlEmEOf+EICoOy0eL0or8OyzjZzTONSBwu3uoURze
oS6JVc/1opOz5L10e9me0M1PBVhiK2Zc9l76s9P/C3VFcLzhb9KMBIPFgkxjJlEB
jCUXYKMcIMwrBnf6Sk84D/kmlH8yUGqkP9ZZhCU5OvVvf3e/uosdbsLV79c3dCcg
UYFX3VIqBdG+mrjgPf7CLjlg4Jj+w8JDrPyUDUL+urMNA4x2f3Wue7iSdgBDbivA
wnmAc9xnsPT634XnxKKxlRNa1gdjgg2fKxcc6Ed+hugFVgi2g/xBaoLguQOtDCdl
bLV6ZL4j1QYxCSAm/dfBcPOfBHfxz3ughFYlY4/WCUbC7nuFPGf1bSRvdupZgmaS
xwUCCAlNODthXAPLcNdiVQuesCh2PAjQb3og4DQcxbGBG6aBIzUizfJX84Sa5mmQ
erpoOLHenHAs+U52a9dLFqm0Q6/is40ZY6LiQ3zVEHm5vqRYbxusIhVPCjTznxwq
6F8J1tWYlSfb8iBFKKhlZI07wLfmIZqTfuuLABAthi2QpqhEyLG/nF9rrnJCwWAR
csU4kVa83bSapo/ur4HLspZpOCqzv5nVih38ACCDFUcPv4j6UUhp7TlvveQKwYF0
1a35jxQ10X4UL4ZbxSy9wiUb6Bk+WqpkfgPYpN9PGEEsQtxRPemBQ8MdN6RPo7Jx
aTCs+FffIVJaSiiY/IhArmoHB5vbMgdI7vvygxbaPVfZPaAVWZ/etI+bB4hHeBk4
8sH0/zQ/OWEKkr030n9tby/P7ge0JORx1G9jqsQAug8iPv++1Hb7m6o73pww4P5Y
i/ZDFzj3lzEvelR5LLRItbTk+VwG4URm2McG34wYyMMiZ6fvCtkBeSiwRV1d91RK
k/j5Q3OldzP84YF9wguBw1bUzR/IYpJn8oGTK/SjDxK7F7HZgILvC0T7PLHw97rv
9gqMiEkcTAua6XDM04BeM07qoSu65KKDEM1sNxQtlbsyE+AWcdeP2BgYbVSHBNlp
oRTIdZPU2HA0e2OleJTB8pLdCT4ERSofy3XUJS1k0DKM7Bp7g001Wk/XMkkm0rv6
tiuPVwGxqkYZyytW8oXexO5/bxFyh/sWsyg56qv/+17sk2PA9jWBdq8vn+WEwLkN
gPzigKTR7D6Jw3GKEfGUC0jFs8sU+hPvWRasKzuv6PbfprmVk/NP2hdhXyH1/m0b
yFDGhEEQyZgR/j3INPNl3BI+vX9EN0Il+xCvNAaKot7jGPVys63h8Hv2EwZAu4Iv
bRWGyU+3/SD2Hj7c240CwkLFmu+v/nKsZjnUeS5b+U/DT4gge3sqjA9sKyN//YQG
P+vvSk9uY67LEL4lpM6p0yO0IsMMHI4P1ISz0dbRDrAa0jSE9UXEJ9AGy5+XuuoC
lAgapEpN90kzFNK3yrqqOzb7FmpvoRg3YIE0mffliSjUq2xLlorDG4gRXoKrYUDY
BNsi9waNbWI6SgwueHnWBp15Tod4U4CjNkl1NuSJb/qXWIm/ENS+VxOwamCITHlx
EuMfIRGwMGJhIgX59sjXf/T2gAwqBNW1aZH/fVuFtrgcEduspqr4MMopeUMG36Pv
3qOkl9RohwVqwqcADJBmT8qMxyaV4/Ii64Ft4IrvUBL4hg7AljrrtULcL3x60vs/
Ine4swtsGeblB6DHJsJOJheFRHKX/wD2Fpqi/9HFzB6AFCrZW0yynhflFYzne5sj
hyR+KOwScfpacxsHpa5P8HWstDxmI4wcKD2ISRxD9YZmlWy6YfCe4NFA46D+vBJ4
LvZ8r0KQt+lVngcskZDO5mcjevSaFFMymXFtuxrtZbIIS+U/WRtWvTSD5/BG3mU9
YFsFE3t1lsSu3gernkPnOfkzDOMGLNUBp2JTk+nN4m4hQxrhTw0E2tObHCgBGFtD
KE9N+uQ0P6gAM9lX1RNLzN370tFzoO70Bjfk7WlYq3F2nLZ2sj5OuAHCx/t3SLd+
5usiXbV4VmK9j6XwxsYty5zgamyDPC/cFzhHnJVYOBQUm5lhB2zvXgDaiMV28S37
r4t55LaCL74gA74K0ZjhKT8VjEAEyN0+SgXhED8/CtXGYFtc7OEhwN0A7CCyDwqe
kqrNWVZUTVEM1CJGKB0fb+1wCs6ADiOkH87VtFvTGpnacdgO5v5ddH1LvI2UKXMg
4enU2t5VoXNsCzun4d3rJchZbdP27VvOBQ9p6ANRVoGz3HO88xe5ffJ47T9L0WL5
Q7FhFJpcxzgJvG+Zfb2jmX1+cvMkPf+kkGfNx5BIKbcXzNlA6dxHp7fezuVyKY9B
x12SwboEj9XQtsAJu/DPVdsoI3rRGA0bOzaSUIing8GjDzUp18UE55TI2vp5czzj
9iqsY/r1o1rGlOdKCU/PjPEJUr95kX5rNgwHCCe+LXmd4dYbENAxNR6TKlR+MUsK
U48BRMiHFx/homAFQjqy25ffn8xblwZmgrmgZOPjWXe7Bw8109QnJE1vD3KT4X56
Lhf1wTgXRX7WS6G61CSnaQCvmbk3gdbPaYTYF7GQ6Q8gAIIIONMelXA01QtgjVzD
ZcdJV0edv3ABrB8hVE6e/g7YrXnQm0Q6HyQDf+LzH4giGocrocdUV5MoMi89wjJC
OCxx0KjH4yn0QqWs8O1w+7Wawfmbn48qyOT4+h1Mu6oJinDvHRALxMnHRmfpjsUk
t6cw36DgDtjYgL1vo2+LFUYnzFtEryuO1JOLx3gWCdNVweBNQNsdH++47zyYt+oi
iJaAPs+44u8nQtuFKSv/4AbfQImLc9X1yy4B0BBr6TR6Gafu0/P5Fu0tBN4UjEAS
HNlbXGvxZg+Onrsq4/7FhUxXGgadRDSvrg6lgPS8Zn3dQiLo+p40nMyk156Lm2S7
dW+7fRE3qjpfXVab0B7b4p6KA5sog8PzSalynKajMfz4qtro2adA5hKRNFZNqO9L
MO3sdGv6liucaudckZOX1+RIf5eUt4qC7ylD1CsYlooUFyXsSd1e3KuZpOm3lMQt
Vr4h8+SzmlBE5iIsfvF/W4cnubgAKzxGQzxjKZ2mxtz/H2G4GAmaTfvw2P2C5Ccn
78/b6LFDZ5++C0Y7yOL//KoZN66Hpq2rpp3iqMoWnXGar+xTrnOboKy9YLmLviIo
g2ZyA5LdOzzYd84tCE6Gthiv6cwcwRa4mXjAiAa7UtJT4VAthmyiU2u9lqRRGRHi
KUWWiHkWZaNAruaCOzihP0eXN7jFEoS8ykm+7LcpjF2LWNUg35G720FMhgVPRwZX
E0d7dGiVVXFByknrFwKTBRT1zVvScD1i39x48kw4p7tJvq0JiqZctKw9cuXnkmHP
K/X7VzF6pTZQt/t5+kzutll7mSjz+4Reoy9CJRfT+Iere9Z7GnXFImOsMV3+rx/P
pjZfQTeujvHiZAIEeJJI6VQ6TuqmkaRltFOXKPQ1WbVp4bD14nLt3ROkuOEyvqEF
WEqdTrIlIUF8IdfDHthftVeNikA+gbvWueMOIzhU97eTWuHm7DwpJeF7AnxkvKeR
5T5PKQgkRyLsnrY+tYfNQs6D8GQd/9Qa157N5cfOyvBgVgYoUEpYrPj0HgwMSX5i
KbI/1ikc+pul1ml+fy/kNb3ylwAjn8M23F7tN7gDfGTr4xv9Lb5AUkZ2WJBllGYM
rhxeLxS1JhGGWd67uMEJYMy2PARSD3MRrBtLbQrgE0QfInm0wFzJpW2cpefo32yd
cXe8j+3u9GGIbAugYvHkp549vRP2act6gjIZsbMSTI17b5GDAq0xaYUWceChnCeB
sr4GXenIkJ+9LRHcJAqr8+KNDzoXzVjpSxznQsAP/gNRrMFFl1IpyarKQe3wMv+o
A26B0tjARYbSsBf/Z1f9HqlBrcp3X5dvKSTMz/ak+cms//tibZM75gVOM9UV40CN
7c9SQH6JnHGm+DNYbL+xnVxpbzrGOdgIRTXaROmnYJR+XocjUwM/nUpqjOdw8VlU
Kl03rB3knr6/J0M/Y/sCfO0k1DiZb385uR3Opg7XsQzY8QoXjBDZsujpQSJbBaFo
zeqlrVIGZZA1Lpsul4Bekc5ntO5x/8alycCZSND58COSyts9Swue4NcTgzGfO7vk
ZdUtc7RFB9N22su8SZNzNTp0hasrCYXS6sktkus2W+/nCG6hqyNNo8TQ17HWRUKg
zlupthqGiuOd4BASXcV0maAj0NlG9cuRR5Cl5WZmubv4mJQDVVkps/OT6YFpYnHp
VGWrMUGrJtdU/OWEJIj0JvhUvhOCjgflRGX+37xxctJEFhUOs5U6vqtXEwvATIvb
ZmRI8QnuWcC+vZDDNBwqAqjrbTb5U4Jagmq/bjMGP90iwarHxxCDnNh/eSwNyy6g
/lx97RvjjxvwVs5duHTpjxniervx8FAuFUXKHJHt/3ker7a37tIw7fCV0zsmYz/X
GdYSCFuU78AwAI9RQYvvXdYC5ozVGW3p7N2z4LZVS9Yb8lfgJ8DiGg+1Tj4eWmw5
M1RsSA30AFHqmfVUVQufSmQgLQga5DbQSu4fslCvKZEbtPiz1u/hlRzWcE60vC9m
MuI76DulDSyWZPDQXAbh+PUBs10sGSKVIRYjmlK7gw9YfzgPbFmIiIyQu+KwHR9D
OfviQ2cB5VLVbxjw7yP9gfaa6XdvgsZaV6YBafBtCCDWQKppYP9Kb/VdUQokvJMI
h5FrDlOhr9lbNfN0FZPFk7HiaORhjdkHrwRLR+mndz8Zn9sxrfWgQc7dGvkHal9p
gY/pxk7w2PqFxB9JAVbPiJUCk8L8dedXUcEPlY/LKSbEv97FFbWuAj9LTQe35J8p
0Q2wb90z/XUYWSyLAE0npptjeDJDuv7GP3b8uCVr96/mBQ+1/GzwJB5v3jiSyloM
pilq/C6kClAkSOFHRQRbCApemoNrJjOInX5ro+VDWmIP88d0cVKSIn8GJFbdgwZQ
9FVNfzKKSyosbdL3DazIw6yHxYXp8PL9lUINuH7W/sEiyLjcB5ZQsMrnL0TL01ZH
um0V9fdjpC+mFd6+SyXEGdOdlWsK2aHEhsc6Y6jMoBpdOvZLSuRUKy98pXymMLZq
Xp9ZWoGSM/tDbdaJ2CtA3n0MPUKguA1kw+IwO7m1Dn7qSBvXR1xYh/mZJe1UbQlq
1i41LYG1yRzMJ5KDUfI/QO7cGZr2O+QQtvwBSeZohPjGYOfY0u/vuo75oOBV2SIE
2g3AggPFYdKEJ7c7yncLXEWat5AXqMsqj3iL7m5tcyD+r0vNhKZXbZ/298gb84NV
Pa2eJCWgIuGQZRfTIJw0gst1KodNbSPvso7ADQu4vMhNXnTpxcUFPybw/hY9CXlP
gTTT6w+szobewwvh6tmefoGJykkw5vrnd5sygaMksxwA5uhp/pVTigP8kRTuQVuk
44HBhMsmBAKvI5EUTJN8JnqPhgo+sWEd8F9B3h8HRB5c8rf7aMrgE1TA49PzaX36
bI8xf/kUNm7RoMj6LpXIFCe1bUKLtE5pS06LJ0s3hD+Q4Y5C+eLvKSAN8iYQoniG
dOtIwyKlBoqN9hviytw6dBP0kZIfZrjy/HoISeObpaY7mPVr2bNrQ3JY/Gvw2GEm
bL0/3LQPnaeYLKx+lqYb5CsZi2S7gnNM9di1KhYtnNOC/cE3mIbvzmlNjUxF8TuB
NIlPVoOgaEyDEeYpmu2UrddMCARvcMXLMXo/oPKdK3dvabBattU2GhmzPMx8OIO0
TVbdgQ3SGv+lhIGbzJ0I6oruEBBq64UyiqbGAm8dk4LSSvTGdjwA7JUcboSR36+r
lNO64ndrQZboDm0xsYwF+AU90sb+1Q95Y8+RYZGls6g71bfJNbQM0R2qXmWhBu/e
hkVBCjX1TEeHN6ZnfyX5JPGuup1y5/vOO9e3xF2OBLZPBqRvURs89ipUH9bO3ipy
30NV1VF/6cWGsCm7hiAF936RMxmIMIdQ4gj5QnX4dY53GrAzJ0qys4jGUB2YDAiq
PT9KeKtgPeDphm6o4aN4JJLtcGul7GGpn7haN28y7RGyhtoLTotlwNJ00vgxhLWH
MSO7RENvm8IILgT39Rudzp4G4mdDbhG4Cx0gS3Qq2YaGnPmB8fUURK3vp21Ypy3D
2fl2Y/F/1Dt4ymwTSJoEwb8WXihxEtsmtQACqlQkVgm6xDn9zgAEayU6dlazvN96
ONds97d+nAwRgetFKNxRWnb6C5JT+wJYpp/3QQJETd4mMCrmqu6XUXPPcQ4XmlFJ
aAvjp5wJKDfbEuUa256BDvL0z1Xgr9kW36fjCZPD43sLThdb5la9sc1D7+1ou5FC
GWPNmum70CrjxlaFs4n+veMivuIlMb247Dj8srwo4IorQh2mNl2FOnNwJSvjB/ue
Zb2COubHIz41Wia4r2HlTHjBCfoC5zjDmHizxPpdOWJSOTVOYFq8xPi3jcKZneHw
H0s28LfdrrU+EVc7K5Su4ZR+SalL7w1MHKj5cblKp2rqXr7M9F+gKadoFhECzZN8
v82C5QFJdwPhxwlRl2vdkTlNv5glUkgM5btH3blwE35QUJTdT4fnBD8Qe31m96lf
1zVnTGCJksDElGcOakAoEgz24VFaRvPoltoPwKbEKowNqHUX6mRLFXu4jSIrtoaW
Xwos/8Uk5P3UoeSkXDDB/t0SQDyTQJiXvK0+bjQ6yLfZ5xrJUVPAwKE68exqaq7X
/7hf9ljfXdoqueN9X+qm7TnFVSBkb/MEqFVMxoqd+7Xaz+A/QWWneBFjUKXSSMUr
RgAbUgd0mHQR0mMf6kkcr40DuNZOsYktd95SgSNZU3r6PrUT9pyA8YbGNIqSQDNl
XENjgMQUwD52qEthKGFgK7DGEBhoaCuAvSIGocrKvPIq8nDQSY9YLsMwfC/unshE
k9IiaNYKtZPjoyMpN9lgnrZM3WCoDWqNAZ0VTn+gMiJPaW3FLHKdWa6wRGZtUG3Y
Nm2BK4SEJE00QotovNkcDyNfncUqwS975ewc+/0ElnTIBonGHOX0B2KsBcFD7rpq
mYZOIwkfcHUFg5mXoi5V2RYqX/vnaV0+B57qPktRZr8O1y7v8uONX9tgO5Y9axPZ
HRd67PeG/BzdNzZjw3eT6AJPPV4oeoerIpGxS/lpaGDB3qmMWltfrM77NeAYCVpX
hhA87TG3pJMJqabLwhDcOond+2xOWQtZ+KRWz1HrFZnN1PdVIC97nx4pAA6HQT68
LP4MyWG3068Yy12BRmjgmzkctb5CpxGisra0TiceEtIWEgGor/92RM0FpdVoKJ0K
hwQXQTojtx97IEgJHPrTD8vqwJuA1yl7dyoM+nMRA7J/V1ZIOjF2tZ0V5/aUt0at
YBrJ6z/FsdsUs11f9VNKLM9u5ZP9OQAZVnHX7EfamJ0pztNbNIRRN8eXaXI7EA9/
QxaGI6J91O670H/6gfy1JvIUFOFOj4ivUhn2TA8G8vQKa6ipJx9NNwX71tMNRe4z
gvATwRWnOZ008iXXXBdVllsp9Lcyi0mGTudA8xU19rl0FyM089GvE1wNo8bglMQm
Knl6xrtPTuIJlpUkSZHSzOVctyf+v7ieOS0OJYLHP7fyZBQPDNxUGRxLSrpQoEAu
qHNlb8hpcunNmf170jVe2ITqbreJUMBoSWdqQ6uH9+q91nEJ+YxELil2A1qxigWa
AyhE5pZanWQP3ZoHJLYEtt1FFizvwF0WiyZgzoD9et8dUoZXd4veU514agtxuIDw
YDeoZ+3DYQRZ6p8HoSjo885fLw6ph/FYzD+qhHM9WH8owWX87pOHPsyQ8tBS2rl4
v9JkGiWhkjhWNySNHC11ut/6/yTm0+pdtB9ZW3mpGlww5yR040JqgG0IwbBCaxp3
VvjJ/P8wQUrcW0XIXu79rje0CGwl0Sqt/ilVQWu89lQCZ/A8zZA6hVhJ+BMvJNTn
88HkIhCrJxuLmCdVDCN3OdObO1WyxgGmqJoT48greqiAACg4jgGLkDP/HbbU2bzM
XEiJqELLRUtGSLKn8AO2oESpBUAFyCF4KC5zaLwip0FZJl5vtPKU7CCrGqzsm95O
t2cxjMN8FmCCi5NEuRHqvGWPASEtaoCbNjERkyG87gJWnprOCzTwCJuSPC9F2ksB
H85NWCfVkF1K29CobLJ9O1roTKftg0tegsMOnwLmcX6yRXwN/whVkCp57EogUU9z
8zj+RHTwXAzfXA1HTeeLnHFwN0CNRsODYFtn+2wvTZBcZLRryiclFNp+jxz8bh7n
8YDv2lB454Fbu+dqWdwkioWPcsb2l7bl7fuf5pWnxBZfe0nqApd6AEzGga99UHvo
G6qbpGZObI80OXWcvDM+5l2yTLtvrJ6pwiNT98E7i57XT6d2sFL3WjuwrzLGqWtP
IgEXkYtYQPVBs4UyIAVwG2ZLG3KxFpo7O9pwHR4qUQbL4yhSWYOkSt7i7X6ixFU4
DgC8rjcSP+8Wf/d0oGRKwbrz1W6VukUZjF+P4rD9py7haPpCL9s4rvPfl1fxiIkm
aIraEhkKP6K3iJLryGXn6NyqNVQkww6vxvxcNHL95eID5Lxyg0Wcy7oypqiPd19O
6/hXPzs8L0sdd2UNUgpIcYeYME6HMhWivQN1T1tuE1WSEhzsQT4gt3EXykegdXc1
FTFwFfWATswaXUMKXJJmSLPyaZjwbjkyAC93ih+xgSXdP1c+1IQcs4uOLpKvzdFo
fNO7z4sPrUfe7Oni+JUmN3IGZIE/tLk8lvM4P8xWJbZ1P2F/8jcLwvp46qeNJ1bR
r9IxT1yvSXlBQyajjaLxXQUP6T09L/2dGkRyobcVsjgD9AYla42uR4mjv0bbrVVA
UV0+6dJoui6YJbH3Vg/UTwzO5zwN7NjzCmHoz/yjZp5fiLCwm+3XaJ197HCS3JPy
lab+Rs93rB3sFdxBjSa6xwCgd1cdQjdgCCAYAQ/6pAXzL1HoJohct/YGNTcRTRuM
LZRU31DrWUOKrjkQ2DTJ7pW5QL/bPWtO4+TX1Tpr06x/lwjDE1NmzQRgYr2Jf7GI
IWM8/Lm9Kd79+LSSPPcCEaZJo5jQp8q7PguPrMG3u/Mb5X193vu0HXVEyFY9k970
JwaVhpiBYi4kJcfH5cXQ51v2nBcNbcSx1SGhlryX1feBXh0oi8rUySLP3JDCHBKe
1MLseSaZ1yERCR1zWX4FS15Bh4dyNWyg+RGpSTMNI7c/M4jK3a6WZlYYffPSFRF5
eabPPA7Q9jwh6Yh4Hrbm7TQpFy1jJTepd8kW1OAUv0PJx725PN3A5vRdKAbA50AV
hkwyBzs5JJPvZmo8tteMVOaSgQPcBVtvpqcmYYsVConeAG6+KdVFF4O1SYKT7vOk
G3yiEncZw9Eh00RE5zbuqlyw21Gte6lheeV7Z0ojMziLQuQOBgkG2UZANVHveYgY
6BF+5+BbF+6fKXv3hcmjKsMwQCR4NAFTLZfb6EOovBlVW2b+mhWDdGncJXncvK+b
VJ4sW0Dd9NcpAfzkvDk3qosfjJyzVnJaFEvLCclz2TaeK1XYczmk+lilmojMlCna
ProDyOTpv4+UYvjcIuAIeJUTrBElibhpkosI5EL03z2hYKgnrxJykNfYs8FnoiKF
NijpgwCXc5zu8JBB6YmuphjQhYIqnGgKERImNP90vyEcrryw4OEtJeWYLXOxigA1
g4JEHTbavGJK99Vg3wXqW1ZUqRINjmLtwa0qwcAqmB/JF9eC6LN7XcUBkTUZEOFv
pODGmX0M9nU5THfpVGi3dcNc6kzBGX2JftWXrWQFAlBaMmIe5pqdB7kA456bni9X
fHexA+txfLlGqvFLRcDrFkoS9q1NI4KpVs4mFOCbtCrdvKyvwALqAdQJUgYiEDE3
S1GWixeuv+wUjiDrMJzXYq6Maw17pn0gTYwTl5h6Zx1fy8k2+v5Y8V8O9LCa1JzB
6Zuz8FjDmCDIDpajSdfYty2Qv48mD0p7VX6gxtpMdsRj7V+dIFLEssGXTTaTsQO5
8vXeyB0A6L1mFVQFHoeoB8R+Fw7EGjJjbLpzrODZa6HT9xBsILr1kwCRmihG0ph7
5UqgN4I2/Vt2i45rd5Zopnz1vVSWO2TJM2SKVSMrw7FTayWtKq9lGJX5gSsO+4qU
IdTP5arv1aCoWIcZ3LXJF98vOlOXREYIBPcFIhvcoUS6f9OZP6CxrS9JXPp06n8I
VgPL/ibNaIamW77ngJSBsmd8WheXNIsJzvKpuD8Gb/1vOfI4Csm2QZkPkb/2SH+u
IMchwIIII2apFmo3BKjZnp+MimhoIAvzhpsUu/CjKS+0TCP0QUeoDORDbxB/KPfo
ozsN2YZDFvqXjFCTcv0JgAMqjEhcIyIR7T37MX7rB2YwCSEAz5tEy79qBi5rbOF1
FBXHIueLdM6A+2AbatiC7rW8kVGlLYmCuS8Q5ub8OdelN5SSoXRElbazzlOTYzIx
5mEXFb1DnP1l3w8ZvlXZTcgCGEqR5aMrXTInZytQRPL7ZIDasvi8NpxX8HXOUAyc
lm57buK0Js9QA+L78LfZvKS0o2bbAOHM2OYLAQiCAstkMVf1Cv6D1iTIOWH4RhOY
oeerEIiyFYvoaY/Od08Ku2Ow4pBombHcn96WDC59S13tk2hgBG21G617/vE2Mk1/
7JwcMLtmTIhrAyQJTM9NrHEf8F/NfqyaVXrtozLUPs4gVOYn45diPz23knW53l6E
Bu0F8BZXnMs+9mmOibMEjTF/tjnzgbhLRp1aohxPqcsjtREtlWXa5j+3ce8l24pm
/NDlXMQ6sDjTTNHGNkLczCJ91oJzQuy+U3Asr/gDJc/UqURw++1pXelkIEMEHeKe
qRLbhWzQN8dqX0WjugB8bD15oSf028RnN7rDCrhvPpmwZhRyl1sPjHc7rnEX1Uyt
p82dn2CCNQIfCG9EBRKlw7ZXT6EJXS+vuCFlA62GPbCIekJWc3oTsd39yJNQtbzp
oD14CIoxHk1JK7z5gtfqeJijUxkTOQd2S95y7STG7D34znBLoVt9Xo2bKx8hZwG6
eWv6Yf928wNskkoGilO2nvaA8L2x47T50R828vAuugezNO8DF6ljQOKyGQSVAcYf
BF5xuArHBmmWOJh3GEmCffqNIcEjzp3bBoSjteE4z6XeJUY4FxSnaDTq2Yd2Q3MO
QWqPtc3aNx8CHnbjYDzE7drCyCFV3hmPIPEg74uC4FwaLRQ2fBSlUUt+fgnmtVhx
980FbTgIwx8MG7JIS47N68Ch3d+VK7To1QCZUOtrGXcTXumbB/VTkWJXwdzPTyEA
3g5JNTkd9cpaJoNU24GbK/xo9cwUtbViLK0Lf1ZZrPc7AR1kJg0FXTeHs5Olfg+q
l6oCPfL2tz+06QQTQ0KumE5ChH6G85CUtWDUqYVqAvM/fDlOg+R1H1BI+frtmhen
6B6TZlOXhzMaCWaxfpPb3dFxfuS6L4QdLjgEMJBhiUJoWecRSl9V3xi0JasBqhA0
xhI+cZTtm5tQwVnpMzTCwYqyyKGKy7lfutbZu6eYe1uEXGmPbbHmJo8YA4DKChYN
CSbMAlFMPOPHdsyUH3hKnMp/2FI5TEeHsAsvjoaktPiibUpH/bAfR8eEy+FqcTid
uesEAQ1pzTRDs7mbujxSVbLv1RUjc8a+LndXwmqjg598+E7kr4U7KnXlqHd3xBx0
/KPi52kXm1MKAQxkPweTUBYwEBRb7rHKYdESNCTvGiTXwGWAxfSXPsmu94NMhFEb
xtrk+cTxWbug93vLbenMaquuWO5H1B9IePoY0Ca0C4M380F3uh2A7s27unh3tnAh
UZydbEIx3AVq4EYUYreB4zhhjdzGfdQJX7QmjQ5D32GgL0lWQXk7VVJzpJZoXuPX
Tzi6YfrpgQShCiVps7LOZSpsSAZSVrfa4qQiATqnmjD2fAVwZIu/fIxM533jEoAw
QIm9wK4jowde048wUN0S+CaInKgjJtFBBl1zIdxkAT7nNapOlhdIF+RunZ9GKPRm
DmcC9xIs1RijMLqzv9LfsKXy7IO+K/Qs+84HbdP6dqg/ScH6YKN1hMnAjjlRQm27
2vA4v2mKm3MfCl3g5yF4A6WYswarezm9J7xIPBQkLU78grr6uf6twmW0YSuRqZAI
lF6+4wSkPs5FN43uWtQiRThS8QQcm6VZ2VBjI6N2syXuIyJPbwaRrEa5A89J7c0X
zr+Lg58fVAPt/P+xKlJrhTrloxkN6HBW4l9RnWkBnwH5ll8eE0xnxAFPxIqBm3DY
Y3TCh5Z8JDdLv/ygA6fFuReXnrQuCZ/p66IjEWWz3gOn8KLNCg/vqYWuOqVVgfHZ
SNct4D6XA+Nb145gatzJtY0dDjuqe9/9XgLWv06PItUCFM36w5rSETFgu5NtQ1GF
RMv4QIkgTJch9pjBfAxRMjlw/77FMtPhaaNl7cJkhE4u6c3tLwwVPa3tKZmQYD4r
K65ePAI0BG2eAmmhQmp8yTAK/pU9ZNfoi97c9TCgYmqSaeVW9iQfk8WzCj+2FNCw
FPokTek8XpeJOtFWt9QTfkx3y3+FRlYp/sMvRatJDWMwYdI8zUPrJ4749nrGO8F+
d3xyCaMFXjUqPAf+cDaXwrthdIb2a0wG9/FMjsYDS4tKklEbsDLBxVYXaeTCHtI5
lKahzgI0336ZgeW6I485xak2ZHhRNubpYe77qq0fkUR4GipQHWTGfQ7mvm7nbBV3
4EGXJ4PJIGabIyfHJfq4SdIXh0j1jYnQS+GSNLJDYSA4EwttipT4C17jpoCiE2UM
rWoBQybvx0p8ErbTZ0jG66oKlcD/O6AFzNMX5gEVD7gszc9+qU048NE6vTV6rLB2
+DSy2YuJfbgK1X9q/OFrlZjxeeJ+X7fVgx+6G9YarkdCVrdi6qmX1dzfHUDnvtiL
HMRdNcomg3qsAj4alV062orL7C1TeT14mWjpoA1UqUMdImVunwQe1oI30wRqQmJy
g5NaPiQz86rU9aiSM4HoCh627aqfz58UkkP7HXvIAa468bWx1gj0x4RVw60WMD3Q
MMDoxcpPY8O03rPjSoF6cLR7lVycPQpqlUJUDs6FGPq9ARxljEWCht3BaBqvoWwY
GJjyY2i6HczBPRTX03y0eF517q8ttLOWP5Gxktnn/L6ZZR3lZgfh3aOp9g07EZYc
QNbIiMzxWuJg+4Z4t5ru1gMkovH/D/tnu6zwpsopBZrRGaXoVN/X1BAcJ3I1Bhkl
WCR4iDPuTd03f5Ult8DkQlcwNNC4xdQ2QpPcVlVMUOcjeCwhnZH5y4oF5/snU8KI
bVXdX1yv6Iz4jkqc1zOXQH6TWvZvSoZhn5YElG/XYRuLQD3xC8iyMferxZlpUBKA
XCuwKBoGf2ezE90FSJuILmFlfZ9ZCPTZLUTCpGhtt5z4PKLjcYnRrDI3UKWnqPMH
jyGNmEvR6YT2hJBeh+h0snFXVg8tf1RcsPOM+bsNp06aLybV0MEPC0JDFCsVlw12
lEHMz1AoR5kFvZ4tHSsFDFhJMiylGdIP4p9WOFg7U6vt8CsPbMHIHmWMnwf4zAiI
NDHmLLDKVNdphsf4sHSDqWhePV0UVt0tsqRj2GFfvHVuqekcyOZ7DGFxzoIaHFsv
vqbqSBlHEkBckQz4aUCp0SZYMJJsOTlxUaFXR3lt6Mm4Oy+nD2oVneIDQav6Ja0Z
iKPqXaSYQeBmJ7CvlTzeAtR961aaleLCTK6Sg5Gn+2TNJPqVLhTymIgdFOFb685d
GM0plcsYFBgoBUOqRplk3Vs1BN/EoPDdwAH/2oBPdFIJg4iEvuwknReJ5a+MwO98
dItQRiNPsOfCOo4uaSzsb/n9+PbnJ/gdmaKLq7pYa9quWGTP9akrrGjACJyZcP4E
hGDYZtUBbR+/ES0c8r6peaZKp7CnFkvcUsOUkIRab0Tz82VjXZzOKPf3/RGNxUdR
AkOW1XfkoAuiAP7STCeJXwZMt2NP61gU82vdSV/oOQzEX9ifykif6tWHJ0CQFPRx
eYNc+19fPMkHV/GxPXnmmlF1gm25B7b3c2wUCgR68Gfghx1rk9mS5NYk/kmwZh1B
DoQUaTp7AWLWM2k8Z8ds2zXWB53B5hr7/vI/HVHttEIX11jrtDgS35sUNzEVKRTo
+RKANWsJUg73YGi5sYMXwb7NUQrmVzVWKyyFevEvoBv/esQCN0wgoDoN71Fr/d7N
3EnoC8mD68HFadrhNBfsFIxgwQwwaUoNAC2ryrCiSG0nVTXiPBwbH2SvV2V5yFao
K47GlOioWaQYrYomfuIzTm12MBSgJU1BydeCCGdIv5M80WUAt92TnrYZaEOYvKD7
8uxoFcs0ECteRJfmAljoNwgBb638nZYpbHBKP4mkynANPpgkIX6xyM0YtlJCTM+o
pF6e1mfBoSW5pebLa16YXuIj0nmRwwg4A1Yt2GOtTQZXHb7UpJf6lBp1+sDKttqw
39BSuDl5abeT0+QOL9xztb/TrRSf2lIIOo8Tzs4HDQi9bgeK2dCBD2q8DJ9K7e3h
/thuEf3rRj2SW2kOjM880fZvKNaZhHLFlzjNE+tZ2fLzGjoFqa2pt4GS97zIHs1V
5gIVweam03HHttzFwp81afch23SKvVDHIxp2J6/jSbHlMnfBSdLHnzmgBP6Q8Kc5
TidMcrsti/LdoTkQrAjww95d3COZr3PKE3U7CFPuhvlV2Aapd+orwkJ8hvqmvgKn
hldJsfZW3OZ30ccCOroaXhIJT08F9F88dovkLvWh1iCfeJ1Nzq1kBUo1pIzJXkln
l0eaZogHV9BkLGMOW25pNIhRvJGyNVCcnkqZFIIxNLyBzhDYpIcJQLq09dS7W4/r
i9nKFJGozhVSxzl2rx4TQDFSC0fMc+hUU7t0JD/zXsHk1uIP8TeCzDurppqz4KUi
BXxc4HJ8XXhyZy0ddYsLQCAlTQt5Vvi/pBCA6CSxxhXt7PwtmzdDQjRmw+ZMKmW2
f5/9FHai+3Ebqst36dCQokFmq8JOlZuDuwRjpAllA1iPXNraYZiSwBtwXfJUEfA+
dBGg5rt9KH+Up+XZw3SQVkIMbODdJN9vS81M4C6pBYLUyq1+uHAS6Pl7u84AM+0C
4TnljcMZ9+3QckHMhtJ2G2182pNaYdX7IrYv3LeiYOWETv0dnhord+EZ6Ve3/GNz
PiKr73r7lvs/t9hJ5F4iInSTjbpUadlr5VWdnZ2Ifbqd0qCyNnlV+Axf0mcfTwuh
foXCl+oNJUzsatxP+NrWHRYFmPO/BkwCQxARaexWhPJI6o4I5iuYxNnVvtKa3BKM
/GSu7xC+qxXtKyUitugjrGfJ1efSz2vVAoLwvnDeOK3a2W+b70INfH5wtvYH2sza
IcHBw4wYPhbh7zEo6pFenb21ZzFXBaZTRzmnwXdwDLu+d0fyU9HT1HfYpy0RAXDT
YRTTmtw+HiogOBUffvwdpv4I7cN0Np6D50mDkClOHvnH4eh8YKr+PTAjx9b6qSMt
PtGBMuYcM/i+j3yIKncbiAlHHUcLSR8cnzFjEeF5VnDHKWVEvHsjE26aYTDIPP5i
6/nZzMA24EeMy1EsMfb/wfH3Nw7tRANXlovsaSi+fGnROULwptJCCrwM/mcA/Nml
2QuPDpLAPkD7qWn89aUpboPK5xtfLAtwaaiT71f4F3/obRaT0I6FVHoakH7CCeZt
hEGrFAxtduDQqh5xpS9Mzm+jvT7ipwjmcsR7Gt+01mG7NgzOT37BQQI6nOoJFtuB
NPhrOgdQAhqq6Ve2IM8cLVjDM7cj4+1zhWGJ1TmKVqchzj2pJUN6baE/Ue/m0BAO
e6uxbdBLPSkEAV7TkvRED4QWIrcn/3qb/2kwyCGPoSuCnX2p4HT/2DhvA7NqGZiR
se6qyiLDsqL534qPHQSBxfl94ukA+yPyaMYchFruWGYAqeI/cXjOTsy6odzuIP9V
wWAPLAieYuCoZhb8XwiuTsD4hcST1yiBgfPNeiOr7lUuNabaDBrjvz2ytjlzEkO0
FKqf/5fefuSixjXlx18qJAioDoKxrksIdvlk0wOsibpKBobJZCttKx1Se269+CTD
+E4F3idMjsuQauTDOU9i8h3C1VWivDIGEP0Sr5+EIwK5cue3uhi3zrxxM1DW8Q1J
/aw/5R+l/fjXVFsPsu0/2QQ93QYs9YBPIJZeKeuUHUldN/6MI/cmCK4O3athWboi
8+ZpfmkEGvGEBFMp4MncC/QQcubyoDmu6iYayZ0XxAsMXLhwkrtQxyrmrv+LtXUs
/DqZDaP7n4vywQyw5QKIftdI7GaeGoDn0zhj7NiCPz2MXfliqXJiu8JbQscTbWMr
fdXQVe4vh/JImQw5OfKRHRbh9BkFNp4QX2/S4vEQ8ctIZQHMi1yXBU9DPFfvyjMv
q3i299qHMHX6FnGgsV2AqgT5SnOewAJbwuZ5ChF8ZlsBj56MJ1Bi80vMzUbjAdYo
YNkyfd/RpbYpSx3CgIzwpcpH657VAQyWuwSnZJCAW3jBCK2ejDKbKgxXG8yyfoAH
gLLUMMAqMLItoAuC7cWnqq/l38vJ4dNOFZczwLbEkR1cVEFuwQ/8tQQNy+/IDooj
cNt1W0PwOgc8lls0NCPOlvpo7T/aYK71w3qtItotjMLYI6d1CkgFz6tWS67wtUrQ
usNd0jV1DGoitGTQAn7aUCk5EAocxHqP1M3u5+pknMmKS6m1oACMFCYOcRHEq438
qKgH5AC/6Mf2PMzZ0vVU6HzFSx/R0ADnP/sgoKiRDBtGAU3S0bqjsvF+fj9jz1lV
wgqkneglTNkMupxbvV/hgY3AS2jMWbE4JrANhn0BV9486N8Jxch4SZrhySqZRqvh
QleyiSdZce8XxB4Cej4Xva2wK+/pzi57bFNg4phd1cJs5WxdPhhld6Nx4N8Tdm7S
w5XFx56dch++CD3q186RKMBRZUc8f8Nc6o+BQr9eHB6omUyicdKdNmi77U0zydIJ
afpjG1xctCOaejFGZb/wZ44Qaa6ZWA8W2ePkAePd5B2wcig1LfE7bk86NrORtuZV
8yiaHGNE46rnLJb3qAVnMv+JtIrS2iWnYNQbxKbEM14tiRVNkN+5TmuvOimqTJi2
ckIWyyk9nV903ShAD0uh/gz51RlfhOeR2aq3Zm+5DnpuqvfxoUYUL6ULJYD0PhWJ
Sw5VrYfjKMjkFXprSA0H2iqSi1go6GielY049TuveVR2LBGw4tdJq2PcAv7CSA7c
h1qtO7GcvDv4QlzBxBdwryOMxwwghcgFNv2v0HVBKKtXDZITXTx8A4GBL/D62IFo
8e9bUKVcJDNxXK+gR5L0ZPACKq66ZOHtdhYx/MFgUG08JmfM5gvcyJw8ggjVMRF4
3d0HtlarQNgVq8EfzRUoCk++AiVqgjyemhjiE+NTpXAJI0ortM2yfFYlYgMve62u
mrMPnj0qdrm+9Hwvj9+/8aq3dSz9qntKO5zGHuALVjWBlGGw/ZS6cPgl3roMGpYd
i8tjX8yfuN3k32tPeVxjUXmiE3SkhG0LTrPWJ6VOJ32510vcOOtVYBCD9fWF1r6p
vfa9d44YZxZug73PXr17a9F+qzUkkDNA67qt3ky+WEegctWJOxgY/X/99dzdbvTt
VzX8xqRFVkLh2dIAdxd6zU6J4RdGzv5KrS0cCOd4VwbAc/6MrQBRXdjw71PD78z1
OYdpdimcw7EmsQLLFgHd4dvE83yFsMFfkEeAMovb3wyOHvqqeyEU1+gBgKuqgLOR
UXiB765nQFL5/88rFF5EV4+6ja1Mm2tC5k623ntx+llL5IwUpIEcozrFucT4Mh7o
vWwsX8Y/A/V0IX6ogdnNM3yr1tiGcN0Y+6W5BtduL/kEcWHV3ICp8xSqJlGUi5eU
gpdO1a7b5Sj/9I8HcLqYoAq7KapHS4WBo8F2t7MknnwwdWphjfmD/AmIQLChahWX
WKn9rvwIJhrH9PG7jnEbKiK2BGwa7TA2HYmSiTs801LzNisqpOKuA1XotX0G+rQZ
JBdH8dk1mCx+2/DDPIb0PX8Vcb/uCXJYxHDggRNGXz+tXjg/bgRzPfkCMWMU0qgM
i5BbdaeFtV7ox8cHhCr4NZTj7tEwPzKXU+8SqrwbaAa6obORGY6q8JOs4Qv21N2B
3rgZgOFfzWmestfof/Z0Vt0O1hZVYHJtNFyRyF1pLKpnincl20OuV9WHFKxWb9Rc
m3VQobXQPMYoU6WuVnBrAAqMMOBchigkNQAdp+6ETBcoR3c34l8cV1BHnOqNl95B
3JPiHu4LOE+EzoYqnoH4xCWFwEjLS1eozg2g/H6Dx9gde1CEKp+h+vQxBiT9JJbi
34HGpn/tBGaYuZTJvQXdIA7jUwKu3/jnF0UEubvF1U3Lo56bYEc9HTPHCtmJpAt6
oMFmkSsBvO65pwhjCOWy8CujHef/LYUbv7p/rrBMrg3jsPJpus43KxjGSmN136Of
DoIVZ/MT9fXxvQaK4ZL9Kat1PX/bY+jsSMvWVQmWk+yUw5vtXdZm88MECptcxzkJ
MeskAYwsYgex/+k0QVg2jo3evoUlMRYBcxDcDNQFJW1A5HEa2wK35TAMcLHXqNLx
cy3Zlc8RQk+6FNJ0xZqZWbKXspQQsOCnZobbeaQIbcR8FxmIDyhhGiluZsRsOLWX
9Y0GMlUeRSxISJBIkmV8NHq8w7EhJE5tdl1XymYjvO/Qz/ruSpHNovYjKnFaVply
CFrVQpVz2euq/dHMyB6wuwIYqcYWp6R7LAo91EclWkFmikAYz1Su6mJD3BDnqBxL
I/YqHNGBhIuAKNM/gs39fNHDzm3UKZrm0GGsgpDbjh5tQmGKZmoGXmLv+gaYHiOv
sZB/TvBJujivbJsge60G/l2R+YphDzKFx0O72h7jYjvxt6cw/7gYQofPGGRJ2MSL
ckfDitNmKJLPzDYlO6A9MchelE+LgAOeY8HMTB+IZA6imBB/li6KQRgLbNhjMn4i
D2o4zvRLwbBwNrVtGDnhXIX4uUECd1WAve9CBzARs5h8z9eCT3J2qncuDRVHcC9/
ISKPawPZfRIMGliSdX82jh4qt8GjEzOk+cJqbWBtuvwtWtlVvESwdkHAnNmeE2f3
yVUGi1ZrdhplflXMGo9oBbJwN08yfkRWBiFraja3+6XpFsWtab+k040jSnEmPtKB
sf7TLCa6Nu2oceSwSmK42b8N7sXM7Ivr3Ok6/ovtH3mB/JERBUgdBZ+sGbLR0D+U
+EATmsHyy9ff6Ct9y4F7SZTYodyiXfQ7yqOCqP+9EfY1k51kVesDAwMbNSgnQvuz
JY5gHfRgnFQ6cVO91HtjwaIYwKkpHIoNfWyo4xnUAyHK/S8EULaOJZhZtS103ixg
wfYTxU5O+S+9qlOcuU3lxlyXslSuSTbZCg2cbJ3BScRXInlxOX+aF1JxKnhoeBs6
nuu8D9HZ/Vj+GKmJzRLPyr2uShKEtAcsdAxIvEoRpvbidyc88DAsMfqbm1FPxTit
MZa3xdKudnGcxIRSgmlr76KYuWgZwxqpbFz/xtpCz61FjjctyWbOpa+gDdfCvV63
pOSmKt81vCTbh+83RHZybnbupEkV5hILfGIqB4Y4XaFLmHSGZXYPKWZVxaK4g3Ww
Uh/+z7smYeIaCLjzDoJuGxP+1JyNw4hrOT97vHc3OM6dPCgOizKaZqA6ruRHTWic
PUE03xcIsTMD/tvd0K4SrZdHUObdNBkP/4GzmN224tIzQwI4uDm/eYfc7ylp+tkF
HDRNowO2iPbebLJwF+K1+qfm0zW0DMCCbxAZGk0EO5Z+6RovD1TUU8Ea0+WhRPr9
tTHJ1Z8CY3Y42meP5hB6dUWhtiTHOQpRv7vpvMWE58fCvmR/IOSiSicgi/+2ZAuQ
I9y/eVp/TwtOGD9/7y4dSH4dtVkbhMppyFA2S9Q0Z6QjxizWmSvUBwrAF0ZXmoRn
HBqA7riFJZveiT/hA5k1jAGPHZnn+YzCRk2epMxffz6SCOsRmb6ABzsVLVG8KFIr
hTJgMf6JzeJ0ZvszUIE/sBO8w2OpWdcH+T4UUEj4TcAhcI0cii7XHUvBZmkHiv/C
DCeZdBqwBKo4wmtuH6L88gSIH3GHVRo5mUgyZwcw70qddhfWJVLNPXXnevaQShA1
5URC35wNB5fbycr681czsdAc1MSDMydITS+OC7HCvw1AlOhkA1xoYEvYxMSoPszw
2gujya8GDvVOV/BFj+uSqBrGnVljkmVHdJM1zNyAJuSb5XBRpmBuMpE4QTs4myy5
1PQtiIqr9IAwKZv1z0GTAQvaCKIrKs++f8jmCx7dI0DzyN7m0/0kslPDj3cz9YKk
d9iRP6QLHP8ElY+XUO/vkpCRZhFwfdiTsPAcpzFl/x1DPnHmk+eV1qfRrMKU2Rfj
nFyKGzLbfpIoIMbRZrWQB5VAyhOZKK5hLfYnc5Qu6VMrtxCgHqx06rcDSilW3CjC
kz5uDkU5mBClhEHbp/4JIQQNSuYkGCezxxUkQ1ov0UqJXIyKPKOz5i6C1VMZASdz
IcBAqdQwYr5whwTL5iyvVGfvhJDkj9vxhQCWu3T9XyXnxAzc6pPyF5h40AiQq7+c
wcMVXcxXGt++D1BRuW9RHBuVQopLdhcZYwccskwVNmX3W5DcCWsWLWhLBF+cXmTp
1qwsYFwo3GORR2lFHWMQjCd4ugm3akfYYdgcx+/1up9cxpPuOnpJC3WoOPaZd0sC
t+2gMsbMBT+UNYdTNwQmw2H6sDJbZQYjcRnz+p2K6+IyHepmWF+peSu7rQ2196Tv
xmQbAy3omLTlES5Kb84yTtX3kq1rK3/hAEmndvO4ohArbrt0p3nVeNZNDyKvbiRo
BI2kr6ARYi6JBPkRasmAT9HuEVeZQ1MxQsetzW1AeKolF94FMT9d5iPNyKS4TcpC
JdJkS2mNdJp9ULOo5OddldNM1r/WApEo7wAxp0WcaREIWYXB3yeud7lQOUtkYkPd
I58aEWhBRYXxK2NKjlBTAq/droGJziVXO7fcMM3xM67/YA2XPoPpBUfqGAJEJJ2c
9l035hf2c1RrpIb7HyASgf+3ReMk7F/ORWo1Tjy2t4gkBfAFqWy4xcULYvv+/+V3
oFzboJ4UveLgzST3E9IgJXQZoTAefC0Fccpa7Q2f5DlhrCS4KQo4xLXYIemGjiqc
YbAUFt93kZ9z7sHIeWJlLHQrHqJtdyU+uzI82Fe+S5GwRY4TOKIaIR5heZR2N1N8
eGc7o/74JZ7uEPg5d5HgYgzez7nkUItVj9mq3qPatZwHTS/nysk1Z0xSMXoA+LW6
pKkuEICez+HWGHPVWdsvFdbYlMafGasHsDVPKjxrjY9EyMMEWt0CCOuYZ2KDVLkT
GdA9KobYoJ9Wzd/t6nWXZQi48XypZxqQEICJgqsO9/9TpLPvgs4NBrh/iAfmzJyy
PAeT4KkL82ePDplR9iz0BcMmengJ02qWWQ+fk7adne2TCEWcMsDGqUDmoCy4OXZU
NRl01z3oTMeuvWPqkOYdTRB+tzueuDUY3a+mXOQMUUjzZ4XLxMEyBoZ3L2Agtetc
WgVaSvSv/UNSG52nzbVJVDEtnMR+/W6U1WDRwDBIbss7G/xxRrzexV2DApSyCFO3
8+pq8maTcBiYYGgONj5FhzrzfyCSpqkxwFuz1P+6GPqkAWgL49UQ1s8ltPr3MUt7
3mVDKC7fOEsuNbpesnWp0EiqEtoQlLqYfQ//9SRkeW8I2UR4zxQM5dZxUPII2y32
rwISeUfl8s89Nn1T5lU2uABiHfOqKCu+o6/usSwbcwa8c2Mig6nGcfT0cu6H9Eu8
YwAzZAb1hfT3oQAvScfyUOe15H7EnoZorbVWNt5K6C8pLzW2D7VGMAJWZsBgHrVt
bf6pqcEhxXY3cB13lqbKZyKzLmoP9wFKh2OtUtvcrDbKWIgmHiw4HMC1fNBsbcow
/FFYOQCFh97R9YWf7jKO2gjPgIvO/YLXSOLXa3dBRu5ppqjCePbgWf7a13WQN5TI
2wAT+AUoDtFM/BVJHKmwxzSvmwAWgGXrhVB7HMY1WjVPg6TyJzlAMUP7uNvXpnxu
9IxHUVLKrbJyW+FMjvAA26MlomXCmiWknEU7IA9/ZI5moD+rK/3YdESTHHHt6byY
VcaWCg6OZLMjXcXiBh4Gb59XwZd69CoG5n7Bg1s3xQA4n8KSB02bs8wq6Z6pEFRx
YcfxZRvytbZqqF+EV1EBus1N+aVKXhPvjt99CKTAkmqxXtr9pBJdgKCRW9+VWd8O
zZlXsO6p0K6oen1oA0nU3rpTtehQEQhFe16b2dlmeTqeCyDV1hYHYTdyGJ1LjfYS
AWMpUOTfgbpP29cdThAu+xm1HhaZxq5bpXBp5dQxkojS/ZTm/b06/divNapiKxCK
+z5CjELrOubHcrLBqQPBdG/331aTXikHMQRA3PuicPz95VIFc0boAQ10C9VWTdh4
8haLT+gGAkg+J00LxXi646Jm24ZY9nBYxt//Piwu4Vz3LytY3HKZc9gDfCvIJw89
4/GWFr4dIhf6s/Iy5MHr5i8G0k/iyoGt15JqqA4f+akQ4k4eJ4wAeMV6eJVTxHQl
Tu/AzqFN3F3Nlqca+ihZvneE9By3+pBzy93rk6jpjifwmuCIi3LHOWSz6ut5kQp/
CTyqmG7/Br7X+7cO0cAS2T7ETO1nZCDVLstJ+cTv8uApVh5LEn+QX0R/v2n13GeP
C/oYIOgQvlW2Q8VfWxQn50BYnNkl87h6QjEMMQVFKRWmDR7VKnYeXZxVYaNUsUaF
fzwEICr54HX/HJ/VYSx7VFjcxr6PU/dhKQFpTzNL5yod4e14EVGikuLaw/UZnLl0
rJ8HLACMuU6mB0s7ghecHexkQ+MTdtQ5D/li+lLsxYx2whj7ctMvy/3gxzWc0pGu
2/xpHwWXqITD1DSh5vEJOUFbpfuvE+xdOQT6GVddXl3OIWIoHOnRMxjUe7/YeGLT
NPpIz29SE3oljNPUXBLa3Gvns3p9T9iK3EyZIltXnmsZjevwxfP5oG2VTgQACwxN
loOPHbVnBSaZe7zGU/4gFb14qmZgo87PgfH7HuWiB/GCA6Rxd06VIA02Ld6rI1qg
goQPDM9a85kfZF8BVZlmf1dHBZZvaVeQIS8VueVu31CJD6KqsrdoWQyJLePpydoz
02nDjIS/fz8xuX08Iakl/pprZHD/dA2cTZXKt5oNvusXAjBtRoyxYQuM4RyDgf05
h/06pIre4bBFZddvNVfYtZ8NdokvBzyG70ni7TFJOqbcQjmoew96s0pPfvQmTMcB
Fa7h0Gyt3EoNLu/nsFVvoizOvKBJWEylO9Q3OCDoDblzs6VBtjnpmfWkq4sEGJiU
ws5neTg0fvAO1vUq8L6G8IAJnCVoQAlOHDgdj5nanWwHaN1K2dSqubEa/11yR4AS
8tDON8j5JBGSokSyjSuIGgLF3fupesR4dNIzan24q8K4ZFwuce5PfLzmUISvLbgX
QAI95QN5pPxQiHHn13qRkKlX63y0CcmB41pFjjdOp/bjFMHJ0ML9QuykSWmnUrh5
z2tiyZJtmPtBnbfHTjzIdEm0WrCsK0tMGe8X525X2WNQ77xg4xTiVPfTz1PERiyL
Gd71TOSfLq+qzhIJqEFeP2hM+/dbI4UeJl5pLJmIvHo66WLQLlF9ffO+QJHzINIl
/D2IOBGDK1aPST5KqbDq+ExWNH0jeuWoLX8YBS57lXsJ1a2HuIHY92Fl/DKzERmk
DjzJenutG4JVcooCCFfaYnB+aIvGqhlQreCS4FkkhAGgpPBaBSTgh7dXCYK2MeeE
QFlG2ALYOca66i59Jtp7iUa4v/DTXXK3/fATt4gPcYuJuS+gQEbFCnoMToGT8FTu
MpwFhE8siG6IMAGIZNAWpNkvlWOtFG0yyyl50J1A7AVuAAY7shtn2eAR3ExOVjHj
K0nFn5XyenpgIwoQPPA4xqPJWOuVtnMbPR8ObPEN6QjaIl3TUL5Vj/gMc49EbP73
KrgFV9UsKaA3IG7X9v5B4xXKRKt36OgNvRSHA12L1xPosDUiD/3fLSJmzCyVunuX
0Z5zW1VaHNH+xd/M31UrOjt6aCivn3VbvuqaLsqNHCsaGWkk0XQ6zz+Y9J8mCtHR
M8U5dtwk19xKvReLIas9OXg9dfNPlwlw0yqn9hEIqaFO8bo9lvUjpmiWse+f2fBs
vuP3yfEhe/zFHT89iFOsfnZS18+qZ23aovWj4WGea83E27n7UNRxzPm/DN7avgk1
d+glhSjHHlrBE6xykJtoSeA0VrYmWdMlq1gIySwnhxuzyWqKMuHRdEKXzlCcKpVf
VGfL30tBAJRpqM64GVSzGIWEcMcQFqUZZXqcVQEQkUUufdeIJyO7MvhD8GxmiSWD
CeBAX2FHLLkvttAXxKZt+HjYyEp2zEZurmaZXck53PTff6Qo0+pOCGAG84fQrHL+
qz/7UofZ7BH4JXeLgTVlIffrbHVV1jXUV+I9v9kV/eh9gaFwJxm9zwsfKb8nvEQy
r7qWvFtB+Td5JOhgZwRW7mUtU6+FsSBfclAaUruKFFV2Wgy3teM8zCEpfPNWys6G
tIoSmzt1CTD8Z4ZVRLzmy4g95O2ZVSCkTE4yt7hjkqhL0UKRXEc5lD8bKqS4AtYS
DazFo/WX3cUQv6u2aLduG7N+hZMVonvpdK2Iml/u8G8qJvX13zLaRGII8ut4LGcN
QMGOkA8Y3daIDgMTJbJN3G2cVOTTWxTTfW1+EAgvPS9s/GFbNwHII41r9Qxb2HoY
UAFVMkf7/Ix++TT0St4gO4lUBwt7SxQn5W8BcAuOMpCuEk64FbtQRLpvo0VN85lG
SrZYhgqkGeg3mLkSyXKli9pmLD4Yvp9fSqk5ujCvcBKskhgU3+12/7sSwQYeAjiJ
0flppN938KweZQErPaQaIPcPvi1g5hKgtvpXkW4aE/cgVUqv+F5d/6X3FxY/HUKZ
S1DSy9ibJMOw6QmVqtr0IqxbAFgffdQeRPCzzTIhJuXeOdt3wI1hJNX1K7nPhLr4
4CBD3GH7oHAg17EeYXdQxsbpnf5mXVlDtzcRNN+g83tA9Wv3br9fB7aIggC/zR22
jhz0vNtqHL/7zxlWu7sWPY+Ff6Z4QewzFXuUoBZtAD7r0E0NeQiXOevYqsOIQPt0
lKE/PZahcoQpvxYJs9fidzN5LzRnSQipMKv44fTRZXHtavfyiIzQ65fn+zuBcyFV
p5itEHFNqw1ajyMNT/RMklDG5Gntqchk8H6/TGnPzjFVx4xvxGfFW1bikf9lAFyH
/U0ETCK1g5jWD51YY6c+pl1NqPGFw+ONb8ZYXRxa5Snv2Gi7izVDg83b/9keNsED
bwhZqtO5crpN6io6t/RhN5zuCcFd7kFmu/0Lp3x7VgRg+ALAUtVOfELdR76q6uN0
YXPnyCTijI3r/4ZorLuZX798lAsnb2xcfgoDDFOkDLk2SZV9i8GePskmw/7wkzTe
u59mZ456iSWQBIrXbZkKpWQDLiqn7XqBSqBi+5V4yzQvm4fne+JcZX0bq7HuXgLA
8qZB5EA1PR4H8IdWen3FRLiIRm6P5YDp8WpOryzfXXEITL225oGZCyM56tR3dGQi
jk3XE9NGXjKsvVJMYLmmhlYbNjP9DPfIDqmA1KqNFiB6z4bKsh7Bb+esLgKUyHpk
pv9RcHuhOxrXA9bCtkSqJF8US7rU2O5HVa9RAQwlLhTpSf12zKPpYi3Mq4QTAa1a
pUrSL/rScYNQsFlYytGZ7CMWuSx/EUbFvXh29sktXV8AQcwHBt5z6fnnRSvjqM74
a/ZM0V9Rn74Vah5Z238arBhVOIKBbeHPnZV6je8jS7YhlMotY6lFVym/e1DTTZqL
jGr7SZ9BHBQ6iHL/wMLjjgEEc8k9JgczHty5SXFTKwSMnlkk27AH0xKZ0NqHmz9w
pa0RYQT3us6/pBCU+tIdJyDWR5OXGFyYLjzaUi3NEd/8BQeXaNh3DwAecGqwVhZL
LjLmPiZqc9tzfk8MJAQ15b4H4i7PS7TU6qOCTj4/l1qoe0tmPTOY3+w4mdBhppo9
XfsIvLVmk8Oy+idUMkj+kxpBZbSQ6fdXR1+y1YfN4Jafhentm7Ru1T1OEGnupQCp
Eq5qjujlU4QHtPNdhHryc62L0SrQ4CdBpwIOIy/Z4Yvaq40xHGAcNXFpSebbCKsI
tq76iPbCVenbyyyb77Kbw8BflCAj89QGUx5F4/8iSYSu9kMqJwqoiXiT5C9+Yk/B
qvtgXW1yPz/TGHZH08ApRaKdVa+bJNwP4WZc28sGPp4ZS1bckvjLKZ21xE2lrtcE
6TXScVlE6IajKovGa40FD5hE5QbfD7cx50YTavuNdDWOwEmGrsMfmictk4eZDyyT
/nKL2FylrZViFPBYc9rPSoFLR0Vg7IoW5FUjKF+5Fqu3Z88BZojAfIBA6n9tu9Bf
wiweiZ2ypEFTpHnYk0ZCgIl5CvQQVs9veqLaMdVSYw6gQFTEMFcxgZQIHrdL+qCP
GNr0BO3/vtTi4KRn6vaG1YyNAF4xYzygzNuepymAFNkH7lJNKV4ypTysTNqeqbTS
3qsGlSY3GrcVE/qk4aT18y4iYLl3gsdJ6wiKGvBdwyhPiDlQIvWsV0v/uweVIbPf
M7Cnyv+kfXIWuu5rv2vIobm4vuHhJe/38VWQYuLwtMK5/BxWz+65yB6u9pbDoTKB
+XdH5RNsebcfnX4t5LR0Vr7c+XXQ8wLrbMTMSsjqysqPpA3cAjG1cgBT389iO9Ub
eKcD9No2PPH5DNiIqT+tiz073vxqgqrU4V5hQyuL1CbMsCzAE686eStVvsxN2X6f
bwXkm2uysMk7wdbnc3ShT+dsM4vf9EyE2opr+fbfMSpCEdrrgnMRLqtzJ2vlnsmw
iZtXCPt1NonixjzMBUZZE41ObjNwg0H0Rfvyn2w0dgWlzgWi9/yAh9qnSnVh/aLd
zK8xfpXGI15vO2RF5QTHv27KPcssrurMlb+sJwnojNUwwG5eNxDIlYmGN2IMVWAb
ZWBuh2XhblJ6tRVKzU3puN0gQOZcxlgwfhAeVoQdVLCtp2co/7/yHzMDJWqRwlHG
rL2UwJ76+sKwRPV2dTsQplMr0RTylMNdRo8f0P/u5J9xv2IVqSuMwDRmubPGiZKh
iCkEHQYu1Bzz7JeYKxzSDhqRzSEJMCDQFP16XEHHSFUvN0BwYxVFUCASFZT5SIRu
nLTsQ8IA7INUJ8OCp20mf2yWTt0afcPwmZXCm2BO79WJH9N5/oMmkCb7mXNzl9lI
VgGIkGqn3aN0EUZOiCBMW5bY+6HaQu/F8q2OV69JLDZMkFEXqcgHYTD6UOdOugej
2qe9FLTYgDv+CJ9vYNBfdnAytAAY0xagxgkW2RT+QM70HD98aIqEwwQvOqplGYDw
s6Z1lX0rN8ZCOJ+Jr77/hkEtiaNbDnr9/CJb7nrvoKG9InoSLIsK7GK+lScyiQdf
uE8YJ0P/C8wA/8VKQg8/npbMb9/ywT8Elp2tCTdz3VdzYTenTkdW3i20Jv4CLohL
0LdhILhO2xNh2b10egK7bvj/qqLOP/zv9zlJ0COp455b3SV+golrGs4jBm2d8uq2
aN9PzqMZnW+N/5ZqWFaXKJh8eQeG1eiqCP9DPOiXU1jTmpWCpk1WoGrDkGWVA/yR
Etyx0LQ/Ul6mlGdXDpIEBB0VRby8jZM01efVssZnn3F1/HIExByOobuUGBeLOyFW
T5oECzBCB1/zA64VrenDwkrl7RrlBfzFCxhkNXZHRW6ZX/7pX3cvmjXpMoPy2WQ1
u60vt3qkw9C/wzkDqZ4eA/tZoqfWS+TpsI9+qlJgyGngCmRxqfwY9OJIfUa0+jA3
CaGcuZ25IneqiA8KpqTfh0S4qHYRLB/sC5eF3tjVJP+4M4J8jU06R3ShgGXf7d/j
fzgTz7tYVZln+gmER+7pezWelpVjWUDcwVFhTdUHJsY84JYgLQ8onVk7i6zhFkJh
UXvU5gEx9Lmu/YfDxCjeb0AugmNMSbBpzskMqmzcFnLd+5uWGe2FcHlf/anABUNY
v7mjNRm3hqDGwSQVQi4dr0uwBMFhrHaN4rXG0aDXZaPeFDUFUtEuxZhT5nLNd0Q2
cnMe5jsDffxT/aTdY8qn2td09L7jsyyWPLlfzUseVa7arfBjx0cTD++G8FKnGGQl
AaO/5P257IKvRYTc1cgGrzXAm+mFJ2q6U0F+79Cgc0lz8S024QhwlfcWvs5mIhMo
RdNKId3p0SBnvhCXzPXks19sbct9WhpzlFgQn4nzZYzL/Rked4LdmQTQfNQiX7AI
yjpnqWjjjoDjmrB9+Grq/shKvMyXQlzyHopJd2r20Dk3LxZnPekhTx2Dm1umlr4t
UBqomdVTGl82pi5cwdkWBfkrmJ8oklx1hjNVjGyGN6Nt6QjeqhXOeXkFsza8SSnK
b8WMOWRRbuTkZ9Vcsqx/YYMTaARVHaTooYGfyqbI4NcIn0PqBJTsEfLhwHG69r5i
2SHfK/9Rgx4ornD5Omrzi+wunk5thNo/GZ439CvdNpgZMi4Qi8CMWU5AsBmLsmqo
xworZ8xsAJKYp9ETW2JJecSv63iRgtn/YjF4+HZCJR3OK+JwHK8QSyX/pCM3T9ZA
S54mfbmJyZeqJJpB8SCCVzlq7FvrUTFmhfkllaV+heOfm2nCFQtpu1hyaaRotEXW
9/ArKsZroMiywIxkMUP9UkicDOebqkBqNixtzia65fvzKjAeaG+5Sa/k4EiSkWu5
j7xiolPRTjtoNTKkViR+UkrCRpnlrg/FlUXwWIHKnd7TFAmJheYH76N78SV8uUGX
tR3NJOV78u3on7eG9Q0tnddC9Z73MtGteZNmla3GMwzDfkBy3G2wAGsrV2wZqPLd
eVBBZReb/GJtDBoJhnlCG/6rzlDrzZbWAtjqA3BMuLPgvvNTz91OnJEhMf2tNafb
RIqAIAbLEFp9BfnkaMc8ONwU4LgsLVKIHVL+xc7ZgItFsXEwE503EPR4xahm1+SQ
hXipdPQjrHEWa7XfcLLmIS4QBsgHGaQi/0W5PJnU2xzLCinBgBq/bpmhAckXWhyw
4WPQ4B7tfnd33knm0QMyaB1GSFOP7ltfmcqmdMGTayhycPcqHe5peRiasWMz/ydJ
wp+G2ZbUOjvRm0JoMZ+jmtThgTejw28KkBcJIJHwx3Jkh0A39tl57e9rwaIzkYl7
ur2w8DjgGo3JeRyuELSwpFDqnkvSh56Ar5lFkgtWMz7Yn8Du2hFPeZNuy7RW3weM
1b9ClwZlaMhMlbN9NlSSwveStjzOlXoA37pRVEFDPAawYxdZ4p+cuakmgvHpCcA+
MqVpnx5X97xRD6hfca3qOCGBg+A7Hy8UouK7yuhINAOqhNku61JdnEFgsEuqAfg1
cMMqGGk4rgG94e5EuhZxPJ1GD7Hh7QbPwUbetTitGfb0KJax8SEF+SkBzeTJQ9yN
Sd8LPuuY3u/PzsiDDtq3ASNan2whLo+alWtPSCR8JgWYLCyiEIfvekx8OsppBirr
0fZ9qoYscT5ncPmGmTH2ZeG6OwlSzvj/sC0Azsa0/FqgdJAijHxltFKdnbDqsM9x
GIZu9UqU+RLeMCpvHYSsaP0xUVQ4J/3aiWXE2EfAUsnQm59UtAyhz3c3h9fuY2kp
46SSIoiwsQimyelQE5f6BDHgxJ5qmgiLMpVZSSisuWNAgDn9AufBqAVQ8CU2Xw1N
f+MyUsf2NpcpUGrERIMlr0089W24UcedjFYRJ8/h1Te57r7q4mRav+lL23RaanU4
B6xQjFFxM6h2Rp9Tygf/usw8W/qoRFOBf8tkWd07w+TlkDkld0ezMZHu3bH/MJ82
OkOkcmm/ZdLbEg1islp9QF2k7IgePdywJR7FhRmWz9DedLRnQ+9yEVnu/cfYjlj2
VMygjCUyl/qkHct4IMrmI38X6Z3vRl6tspbaANqJMrq0yExZ3t811v7Ea38YXJAx
iOYrKlusvui5rdlTsF96QCltiHhhr2sCjlL9+tj92mIqy2g9O4mI29z9Yb5Zvsnx
TucA9A+13tOH34zibhAivEDGS1Nb5bR9ML/NP+bt76xETW10SSanVd9oQoT8yS9t
BUkkiy2LxDCJx92zS/PtJbVXmIfg2YyjaM99X7yfsWMj93UTZEy7/9NbYTftn2Hz
ImmTla8fST3UL63wOxbayU5NSEH+JsAkOKvb4vD3Iqq/ac2IcMusv0HTvhALEYpJ
a3Xpgc9ocdVMNllLIM86LSCQEKeesuWVVAjHoNrOJMJ9pNGZ9rfeMbXz3A7MCO1k
YOFzTpubFrHaImc0o0GDYdVVKVCzRlXFMbjV0P6on+JJOSRaOx0ey35gS/OEQbD4
haU6Fas216vS1X7Nl0Dk+Uu3o82mEgKiYFH1LwsuAjbhKzRH5cLf5mTZ7BroFVOT
VaL2ayvF4eQwu64SnatorimBZJ6v7RCisTLfNgbcNXnGy7kkkCV2E7Fi3EQ5oJCi
Fus+4yYlJ0FsVY4fTHH5fIf7stWgXQNaI7iFA8wpLB63HhfR9wbOOfh2QrJR2eh0
C0iBrkQWzo/57CpeAymspkNCY0nnie+sDTDHyL793R3nswDGIn9Pusdua77evBio
cR59MMhXNNEmQ5xDR/FP3NvY8ST3HOeNPzjSR52yRUQe3F+Ebo99G5Cw1+T0ITxx
xH+xTfvjy4ookLbsNnyu7mCbP9eM/zGFdjto7JSqOUh0WWYH+PB/iXvF+CdcTcxK
5TVeqCck4yhxyk20UNJxEzHLE7HQhawVYgufQXEy3KMJZC0LP8YCF5u1taXPAiBx
lXAI2Ltsz1YX0oB1M36UIG5Eh6cE7reA/VCXI7exkLlExF/kbF6D4YV8GzeAkHb1
eX8sWFRYXju0pGvnPDxbC5GahQXF7Zj3CV0GZl93peOtETRhFuXIyrw1GPZ/5usR
TRwn297yvF4JFbdOIFDU41hRPKEpZr8gyF/yWcmJyxCF0D++ZghfDCIM6obE2gBR
+1j73CQh+6VDuSAQYZwdsqCSqXRohNChvsDCImON2KMRVCoRwk1SOc+mJDTr6e1C
K7Z+FskPL6IvtiLdykzLsCvAlrOLV6uZOl1za8p0kI5w5bt5mM93KK+EuU/KyyNK
YTrR63ohXojRcd/k0OSGAgmt/v6ShCsaBhTOCDMjOwKf+JjXaxsSMxetywgyhIg8
fiofD4AsTKXM+rM/vUglZzILGXKepY8JLpxno0nIdzzDNoll0i8XYgml/SDejZQr
e4TVxJi3+0TmYQG9iej2TwyWGYd+OWThHoEFSoLPB2gF1gzC6tZO+6PFrMvKOrdX
nqpic2xwTZ+5+6q7aMX0I75Ye8EAuJwp+k0KLpPSew9I1rYKX3rypI7XQqFX/wPD
l1ukppDZgGICz1UUAvGLSL4Dq8AAqCDDlfo71nUxvPqw/yju/+Czihv4kB67mSIR
Imbdc7xV6sgCJp0OTsHPYSaivt0GUgkzGmx0C1YuKo8ANIwVAaXYDxnSEx82mM2/
Uxv/0W73CcvgtXN4pbHaEfCklnHH3eifDMtwY0L9+U6YcI6XIiebPR5L6cqr3nxH
s5z/BESdxmaWqdvHdFQxfKEElCjLRqSljenY+WOLgptbkUOElfN1w6jnCwbAa88l
OAftW69Ol7C58RG4fSafwKKNUPjk3SGTQ98OTB2CCC8mnreYUgL5uWP9BEa2kWnE
ADWWK3PUFa4e+gdOqwbsRoYy3G2mVRK+muar70VwHioKVQtvp/CGinJM/ryd2otq
GD8Swl/eedefGAAaSrAhT6188QCMkLED1VMt3BKROxLfmYbFx0dG9fQZPxdqFqDf
Wfd/K4O0poK8ymRrqWumCrsRzX+1jy5a1j1HsTLJlzWEKsEjUVKJbuanJxR1T/JK
TrRR2Jz+CHIeA+jlZH0on+pvE9iWZ3iwD/DeezIwWcxtnUpaYcrOTf7EpXPXIjYm
IzPevTG3d87u+8ql3MbCV7j3KaxOkLCcqk4EzRvpQLzdWpV2dNcdmSq3AHL4btZ3
C6rHXN5CEMOTEo0ZhgPCX/ixjuCtWNP3o+SceMOESBB+MzU49LD+MjBivNT2b2fq
R7VBnyFs28kDtsbJzNxKBv5y/+p0u0REoySSeGqPwjNl6DLuEyq0Tq6jiVwZxpnT
BwpEqt8W+xizeLrH/uiLCmoKtTtklNtZHTnWpmhHTlpYiqSBHMNJoKw2THXiWuta
ROVn8Micgnh7pUGGw92HJnO+vA4AqX52FVG+Heou8mQVwHEhD+rnDBWs50yePu8q
VDFFXkfso6yd7bG1IF+dijoJuPQuDo+dXnwoKxXCkSWRa3KmD1nMkMCJBtRdwTgY
weHmM1YCZYThkQBF4Edf7dRQDTTTjT8GsztYfYitda2LbDv+6D6xM9rnBXnHgFbS
sFBkKkK0FaTORRhJRfzxEa02Tw2G+dTLJilm7UGzxebuckeEuVBLFflmtZbGP7Rp
qzx9nwuCJ7Sf5hvXO4483E5e3UURLkgDJSyOXBDz1/cVwQRUlD0tDq+bum1+Y81H
A45kN4z2k1lahDjWf9xOMhpV9W900zdJElporFzmaICzli/G679n+BKZqRLLzM58
iw9hZ02uIO9caJXzA95KOBEQlu0IZ0EGKilSzL/pm46moJihdJAGC2vW1rUmXRzR
nciHTufIvAvA+je8t1vj//mVp9ttdcdOYwlHbU3tIsvY1hzou8qz60ZPF5NrSfH5
VvzZioujcI6yR7eIMlFDdIyz+SKZGkMb6aOw51OXgP7Q7cv9eZHrJBJL172UStpG
FYfZU4lijL07JqZJW8JwoNgCUnk3EXujgvTgJd9wwytU3W/Uuj6lnF9whVas3Qyy
pxTrfYb+SGkedG22VwyTO/OM/y5Kn9kGeFX3MTOeyTrrYKNe9wIve4XyfmMhIePX
4C8ppwwCsD+mtY0ZMe8Eu48sLJwzgQ+NrQYL2MK0h3oSp/Xvpqv/xMKPtdpUNdNR
/gn/E32AkCnCfddD5DFoWzjDWsDLchY2ahKUdIgpGqIFybFLWCCxMBeBZZYN7Gr3
6A1gD7iGEf4tjsmmaTDMtDIDtXk2PmwkRGM/Fw8PeD/1x6SAOexec4KX9zOQKoqV
fxxoOvhjY2fTtWBaixkLRrOSDzP4W59n+vh0fBAFwsYMr2CrMBy5HzvsujWiZLXK
Dm5TYALd1f5Wr5hSh3wfW4E4fFCKxjzVVTG7vCBpjX10CodRhCREpx2nj2htH10z
b76B4/SYbhD118kNwalASX8ircwcDBp2aC3lyNG3lU09OoIYGFPX0PqFq8m5e+/3
1cFJasstBFqru75sykUo1xWxig8Dox8CzEje5IJMPN7hvrDm8naWVOapIurWXB5k
5gNvCJMb2MpLHuaGMszbFxS5bvpVp6XV00Pk12FTGrsKnJP8DpDv0Lu8mUEH3HcK
/MZfRE1iUKpPV1EWfaHnvsVftjag1OymT4PFxulZon2Qe4iz3lT5fhtucPTUC29A
nQBr6GzBlpIbrAlYHHK+4f5N/hjd28YXbRxyN+0eEFiAnjhJls4i2Z4tzIyt9vO3
69Y+L+pPV9HhJE6UOnHOqetQRn8CYT87yE7RZB3Sd2JKBOKmysPxoDUxL73MknPi
M8l9HW/L0z3itQwi/zO0oni4wJmmgpNttCNJAc4RgK14RICvs/P0WD71/tf0vona
TcxUIn580jOrBIiJ/wsRjd1OuegvLVtgCiIlOUEYHNcJQ6pv/0+fI+5lP8AexCPu
7SEIUDqG7ktcU45k+8XrrpT9DEPzbtC4pDYyjgF81BnHsmAcdUG5Izc95Xgka6sI
7IOTfbxqfsuFXoevcYVKyGZl2Ry7W7JVUHeyYDcc6QzRRqTf+Z1R6qsVmhAeH3NE
LdNW2qDUf4vokmA0XRJT/Kl7KYmycyKadgLEBdch9EeF64rtNEGXxI4B18AvDwWg
aT3qeKjFDNKozPnvVAmp6fmPka8eRHFtkOuk58dXkaf19LdEE+wRsEUhahL7BIeG
0ErIOvtkpQ1L7l+RO6jXDNpVT2MjxZ+wA1+eR8hMY+g0oG7Xd2Pg1yb1VgEAw0Tz
u2v08Ap0oxhZN3AeC+pCAytedMMPpc5NvKWFV8Gf3LOHHfsCWOdBELPk+9fZxRh0
UEC6njwESY9R0sCa9zct4WMoY8tqupYWnn5452dI9K8FVQnHsGWG5i3QGEtR5oTD
8z/qz+lmEgLHHbS/LCLK6oyihj6/OEsvAY9OWoR3TaR1HcUsG8TT2Rc+0SPwaKyY
YpM4TlOFlfglCnp15azhCVoREKT/pPqT4mMUaYY+Fz8Jxvik1ycgEl5jGhb0vZ+E
WTVQfopaztAjzGUt+XMilyTRczef8OiQVQqKPVk/KzhM35iLVarwuWAc92McIhdR
ylJJZL+jbb5in6Cb+9VdRgbRxL1lczSdRIOUUlto2Qs9xEbVBpIJKfLCIWI0HfRE
5S9PRwqvXPNPJusjYNQOrex5VMY7ZsixhypBEF2a3uvwp4/U7smWNepcYoYaoU6a
RhqxFxoLxt4AaU9dbnNNq0GrmVs24WnZMYOcSSTx0Z+dibXNGem3KifSl14+KXKl
RI9Nwnkiuo8eVdeLzOZa5k8PpzzxqtCReQrqBJXAiW2rYcBmESTXOPyFa65JsmSL
fZXNRYNAxUZJTLqP/ux52y4Qt9nd5gNsUHQHr6wKr/JcebcENRArHejsNxlOhZaX
2bbD0iYvUsd6BLQh1NMdwyUPMptJCfxbv/lgwXLP0OzhmGWdJnC/mXvUnFt4r3RU
WFZ2BswlZ1waXq58c4tj0n8wvmulqGsmLD6ulPlOrpWbWh8x00E64PpmrLulAQdv
fR8xP519i/r46oI7rl1CEPkyXLJd+iClKqxueTdCzfSG+bt8NqD391v2LTnVcxlK
Cm75XsdG81scYCwMlo3imU++gCsf2uPGFTU9+kcoJe3PzhurSL6JPvx/lO+ZSafM
d4GGvbYlvXJTSFFkZvnrwx6edSxUOkOZDVxqIZj5i4jI94KAeC3UkeX4WL8CIMO/
ct3FpA+RLzeaoGYq3KtY/RRX01xTz28FylQYW5jMXg1mn++4JTb229zLgT9eHgAN
+KVw4qqOUeqjDY4Ls/mACgEN077mKd50ej20U3hQqHja+8HhnsqEA1dblInZpNwW
gdozQUsbeaQ16VQe1Vl9IO42w3jRoVgER30YWw/3x+nx6XlWF/Eyd/K87X2+lTPO
WHiDiH41zuFQj3HmVGk6aqlnarPHuCJBacAZP9W96OnN2q84MWl/yNuWZbr0l3di
luOT73kELJca5BjIGlhZnMO0PVpQL3llsl39nLzg/2Q7MlGJ8CXUAZY7QNA1eWqv
MhR8utzFqtwKuGwguLhJXlptqaorcDlgAVT8Ruqg6k8BOdPBqlrs8pIzLzFLzFbL
13GGDJ/AodqpA3YvluLNOvbhb1Tg4cw9z9/FIlI8ZqTDmRhr89E55/QabPFP5gkw
7m3S//qrzAKZu0HeLJobj/egPzP42LDziFNaznJRd/sx753uEWiq1ACsAAt3vLHM
1uUDp7/S1/r06xEYLGsvN+MmYi+CfErsDydFEb6yOAdYOgZa6TWAWSoBHgCO8Eah
GpCdyi9K84EHGOfPHDFdSHBhtEme6T7NwF+13E/y2IKoh+7cRlt99Btflj3YnQYl
CIAEv+MZEOw+iBwQecE19L2LG95BS2C5GmaQeU9/xHjSCcCkvDTqAD6GpvPJPCuW
KsqTEcVsZWAYfuigFBymwi4Mj0W2tlwLQnuvT+erFYLtkFDY4EA6K24fqKt20Onh
Ess+2US/obEzxNQ6GMJKcU+9E21J4nb5kcTuC1/lWaP+iJP2cHOuN3Nnd2YpH7zK
uLnjC2zgtwSNEI941Trtl38RTjreTff/+sIWNpn3UeuwtXUIwkM1bRKFkCR0Ps5W
vusz6FkrzOtA5M/M01vCZALvkX58vHqVLcRR2jP7zR+cqj+iSoVfha7Rd4B7Fzju
k93LSDGwhp1ERxF4DXbFaLCJ2Qo9AwBv5QTkfGHvg36XR7O/0v/2mYVWQE/16Ul9
oim0202I0OCIOA7K+h0tytFqQAI6UNcfaqjHbocv3k9VXDqaxb7HZAYnium7p40x
s+RYRInYLfS1/Q5xp8SZFozS161oogK9KQgv3Yh9fqjZXwyk7YIzMvpm527BvDxR
VbMjzGtE/S9HRLuPnUPNGRpsHu22FHAGhQ9AegFLppv+Bfdte2+WbHK5UwD4Z+Dc
KUmTmQO+CfGUduLz/JFbVx6noCmNRkO78HAjJBwYbwaDfagYZ8FnoHP5gUaiUdQz
ml8BJ4gy4RFoA41viykuc9yWSbpLnlaQEkz7VaRuLZ2tMIbaTbWV4Md+PEQNToLh
ptOIbGOfZ9v2jxhh5rCWqu0RSJB44pS3dgSuo5jRcyerKfN1u9OPLU6mT/0ptwxL
H4oAgsIVl9i+GEUCYw9kA7b3Gby1EAIP/L5C5huiZV1yxcuVx4aPLMb+zxG3+dQs
8GMRetDfDDmq+Gxwl1/S8ClbZQl8muR6IZkMvxevnWARtHiClyp0D/VQEOKDsQTi
gSuv3saeEXkGE/z9PYdTfLqrN/soihmM/DjwEMS/eLAbI3pnEtK6esTwURDnohwH
euCWgMnhpIyqKIS9OIMr9MLfE08e/MIsRHpDkYghrJwjpHOerKTWKQwaR8GlSlcF
/X5TI2FaAkcfEjUbLpzm/RhcvyLy1V524dK7rw/rgBVzeuUHAnw8FgBYgJztL8vJ
A/jrbmUj7qWLQWk/2X2wtkrJxlNhCpW2nr3Q39dCD1v9SO4p+q/icZblLIz2UQtF
/Dd7bIpHPE41UAxe8YWXZbqYjpxtU0QUqUPHHcfOV1DwBQfLNKnx5evW8jDQ3u9W
emLyBoae/jsZSNJt7CiowahJW1AL1bvSg0Z/VNsKkFd+ZjpT0kFF2voXZvLgf+9R
Trm3qERbL2FoMQSPizOY73RGkno6FNKlN282GRdGBliHULhYgGjhQC9YmsZ8dSJz
lgMsdZCSbcboZDmncOJMLtFcNiXiGdaqqnT82vGXR3ypNORLnYCrWPErYbm/UaLr
GHIMAjrvJAgNM6VY1HbzxPhq5cHafAMDKUhCpcVbf+Oji41CV+rflwrrjukbHt9c
XJ0yplXY86h9RjECHexboQSeKJJ5OFgPYKAxCVhLkqSzyWMYJrKWd7fJDwmyfg9q
p28KyG49/foj1C3jIFGk9l/nU0XZJSn+IvvqyySfdE8AueoBrIDkHZIA1/L43vtE
zsv8/vrXgjte/rmK8Bol0xnFBCjrq9xoKKAFgoi+/FKhMIclBLWonWEkOkD93ckV
zUlEg6V1b4XMJC9UNIiD0GcU/SAOJZaF1suPE/gVpa5Q3samxeuHy94C8b+sqebe
Pdq0MQCvSI3jsq0dv3mo8A/zmBvYOb7KL9LQP6zixheWebbo3XpI/qr4i4mmb7hp
GGogRahrIBB3uqmWcK8CeCaXKfzVb68vrWbY8ZKeFhoh3P92UUYTbdIQItM4MsC3
IiHwE5JSDJ91s5xbzmGNW8U+lxrRmdudFsZebrpOkz2s6m5KBChGzHbKiiicQ90/
yGiBF2PxvbapT9LK4UmW3N0aTBEB6YYO4rU4l9oOSk2Mk9xW754SoeUgjvYPbljX
fKqb1wUy+pBS1q8vvEySpvcL3InYaclP6ZNfgyf2mQWMCg++CAnDKR+k+0EbJnYW
d14mHws+Bd2wLyfSp3NJ9Opi4Eb9NfDEQ8oTcNdNRqpBsMCFrUC9bB1Xq8LN/ckz
RNl4Ellc62B7pl35ktt970yZv6lbtHdmLYQWQ0JvC+AuTgkQI9jwv6MNAY2NzXT+
XIOi87Y99/dpk81KEFeuCRR9Cj5Zse/I1YD4wuhX055KN8bJldwG55eDbkeg6mfi
YqxSxE2wvEeQIqa8wJACGTzKCWQl18Xsym0u7Swhz1EkJDjQOtnHMAJlSMR5MXg2
oYDL2oiHklEFirftvA/L7AkSgMYH8FRvyVTVTh781G5WDDiW/cGfFtU1C+K6164L
w0uF1i97dwk1zGJKUEa+A17ep9nuCvC3w/OawfBlVjuvrwBHM/aqxq/F+bExAmqd
IJBnVcuInPWObqnLTzxXrwywsT19UsiyAyY3H1w5uAPNr5bj7Dx25bIr+QlnqFQZ
g6x2ZU4HvMqA8nLbJPsIJGMojslpCyNcz23U5wybCbLQ/HpR4OvAxNZNvZmJ6I8l
zRXOe3WVfz6dvRNx7VJjir7ESJre5iJKZfByDeIjl8h46hvaMjMetsTtICs5qDGS
hCm8g8Qi7Mu3IiZirae00C+Zh+wlzEByVKP2EM+PkAoRPtGONAMF/Rn9HcP/0a1a
jTlrMgDCK2VWKCDFpwhNY3S5WB9ASVUIEJbx7qREaNDT0g4nBS8XMBefogZzAASX
rduXVdYOe98/EcE1DQzh7wMoa9QNm1hBj9jsBXL4ZIEEt6YjDmNp/9c6qp2KvVph
jJsBiLzMJo/IHVNX0egGlQKcgLv6PmT5rTJF3IrA4b/soIBJzh9+mCkSH3WsRnqv
4nq70IkKxqmgv9qxyI/igCC3rdlNvgCdMadGraBlQejW9Iewkku+nYRzSwLE3Lgb
6EZtVkMYX8mOp/NTtMYCFo2MpU7cxPRx5Q2Ddi9Hae3na99RS+6vMuYBQH0wPrKZ
hDJvRqhn+KLQLWb1uwWyRlF3Ad1S3YhdcUY1emwW9ixVyc/x8eEGHLU/p2ESxnvO
NSeJHpJ3JHWjOlugi3LfNwPlqJNtgG/E5SU0l9oef0RQ9fTXXWxkcVPSeg3maejd
XbnPR0t2trFZ77/+xefzsAQxsvHoxQFyFUqVkkOKo5WZpYT/Dl697WE7Y+8QgW4A
Y9EVAeiM0JcqR3WwtJUmPiXSbR1nTJ4ZyJnC3WIBITEFakNYEUOXPGZNrjuH8C68
KTVvoOB+Hfm7ZBw4L2VOylSVjwu+r7ZGmM/nvex2bL41V4Hm1dABqY6RZahiAiDv
Rv8VAg25P9/AsDb3trnz3YmMJyEefIiSJ8j3eynjLVXGDbEoHBjcw/kU/gCLoF4E
dsh0lJ03/JE02xjb/XANHhj4Bi2fdBpp9C048tvRk11q50/UtZAL5bCo1i+5NNvK
MC80A+3+bZoHDbT+apCcs/v4vVXrs9tMxU2n7sa9NUiipQ8pYhlwiktJyK5w6NFj
Mr1KSTiOmhWeiN35h+eXI+dio2L5Jbq7dYVKXHLSAIUmF6RK2KXQyzzW7wPLQ/7g
8MZTri0k4J6eRDehXkmMSc+/PwQSdqZCj3QiW0zclbChQvk9pVYeJNoo+P484COW
/EWnGMyNOefvAE0cqrv913B+tdO9gHaLXZI8zQJMqw7YitVeHjxHTF3IkhJbZ8WQ
9eypOFgVJN0JxefHiNNTRKufk8AdoPmoWvGiKU4VGpodA1OOrv0N6ReBbdZu0Q6j
5/kkEsTRgYUyF1YI24k2pD/UsLg3WQmX1uG8F1N+s9MmlUfuA9bGvTe08PbYN+L/
j2sij5+j6hsQDU5gExvg9oXTYmUesU555Gafl9wbtfpF7JueV1nzKgNgs455uf+d
HSNtKSJZce1u/Ez0l4uTLcbgGTMPLVXYHemLu9Y46dY9hU6dMt1sjG+JwMTEq0L7
AksDOmeb9oQkF3SukOUvzlY6f1+ksb8fO8RoTI4XCUxCqKVHhD8yzFnCGiTS77o5
2ioWsb2rewQyKGtAhtG9iHQBb0jYtvmV9TI1M5+SBiZre30jb3nA36Ti+DaM63Hd
4xwNCZJWgXPGHLHoz+7oB1H5SD8LtNKmmijw0RI1HQeGGy/Frc9nV54QgPUSO2YT
VvN2aNyGKV5MfDPeDHsVZTNsBrCWZolFXDrhU1TJCfnql/GDC4jEYYW7k8UOB/6B
/FZfyEWxKmeXFiftFEalsmPzbADw3f4+zhSlqZEMrcRNJvd5DAQf2udUpYCHpj02
fJ4GeGgYfIrPI56v1ULbhRx0gKG7pbrRp3hw+MoOg1t+UXz+zf6EjNXFa1tQtZ6h
1Fq5oNYHf1JWI+wrX+VNMgTaVm5+Qzl2lKPBgQ9VWTK13+G7fFjbJwTrbZOaZn/c
eA1CxVv8ONNiHfX6XHjBL75G6TAL47qb4eAewFvV0QNM/v09Iimshp+E72XFP1AQ
vais8Hu2hJiPGL5hh2RZphaxgSrteicXLDRcCVT5pM0wAmzahgh7SNo3k+6I3ObF
Zn5hF7bIVGnF4fLy4B0ooOOUvrvc/EyAsgLgYd6MUmhnIA1LdmftHzHGRYt38SDy
Ys6d7STUh1hNuLop3IdwLqwzIhPg9cGpvBz9E3Q/4gLdwBLLVIBP6imbiIYCT4ue
EkPN0WYPDW8Fry1ZopTScYouP9AMs2BnviSLPgvMsXta2lt2GwH2/81g2K246cWb
+793x3HQlRkwAAH6iIAk1xGkg1C3q70U1ZH/mg3IEaTm/xamZKfRS7GOJaWgbtMq
FHTRzUuZyvA8rCLu49cYJEYsfZ0l8VuPBiXubmopn2QyiXkuKj4e0QxQLVJMLdCY
YNsyKJG1Co+H9Dzq+loJp92Jco2/2Ilr4wZdf6EHwuRtG0lG/Tftwnqp/7z7/zR8
OUgiA7awjAIXACXSNbFAj4pahmJdOKv8N2eqE5nTk0ul0DiwTh6UwbCDxWx9g0CZ
JzxQS6sXJhUoXquoAejRqkM6fDiIpIfhvx53uyb/xOWlYC+pjN3qPkRmTrgR+RUB
gcbv5OrVWM5LCLi4Jcd1cTCbv68YkUtRn/9LcfUX68o5/C3mAIyfDGd6jBX8TrDq
qHHqzpl+NQL8+9KAAiih+SAY1QgP1X0Hxmt7jV5BOJcQqYPhsoN64FbQ1C8h4IpQ
+Gd2RvJidn+sKh1oIQl/JJj5HNTe47n+SqwlX9qsh192QMjDd/S2VACyw/HNAj3g
APlE47a9JuaAfIf4726aSIX92sZBBSWSIArAQu19zWsVek8qDC/0KxXKaFDQC6sQ
ggLN+zWFv+wQXuJ6NjtM+bbocvQs87+nZuD0zV+p7tYI9Jsqc/c+/E8iZwwArjx0
WRGtm0UYhKcAhnCDvFNanhwbD/2fE3Fy1l2eHRR7mT+dICZ/Bgiwxyt507aNomnh
xqdERqs+oa+Pm2SzUZsMzeOIaeq6n5PfPCX4G6LmT3h+jP/6teFftAgnaI3N0k4o
L/f9NFueRdoBSCDiKEq5zdNBx/H2OCcN8veuXrv2ty4HJ3JxsAiewnvDpROUZq0U
Prmh8WkuSetIqmnWKxGzBnGaXTj5T0UAca+Ary9Ugcb9c3yzBcJNqo0HmtZDo0io
ooVKXo4hdJ/NghgUgEnyffFVRzN0eEO8gPz+/TC7VJTQtm0D0gv/K4MlwB1ZrgXs
Lq4hJkcPJ1xx1BxgseLIhwcyc5JsrN+LqOfI/dcfPntDsS95cxDc6CpyTdyHE1kp
tpZ8vsj35C+Bl/0v5o0t7lx7ClcyjJontDVuQpkeakxX7Oe/J127EHoI4Rwk2erV
eR25aipA6PJ6xb71AdpDL2KDdbl0g1TB3nEYi1XANO+EkG/HIuhugBifBTEEcuUY
Q4HAdBWc0PWSMACeAyRs+Uv0Yq7dZrDZhe1hxOfUDlMVygQaB9tHOkmeFDcXLyWx
hzmMQkaz4H4z6dKNFPxPgw10G3ss6L9pKSvY8Hb2xDlE+NoP0ZP5UQn/0fO0vXIf
0q4znMgXKO294RXx+dGK+Mij8NWC/9rhhCWrrWmXAwQ8GN6IPBxYD78lgem2zrde
zbJL5cbtFHNJHmWQNnbrJY586xHwDxk0Jg/bsZykfq2W8b/hA4UnKxFxFW2BvDVi
OxujI34Q5kF021tIVlqh2n2+C8xPnsIaABNvc35ljOl7iuOdE8Fc2sBdirT/9OYn
E5Sims2TkZeAdpxaIWNADJcGVtE6WlzFTcJZ2QabGMUG5pIhsCVb3cvX7s5uzIz+
OgnOWuEHNrf7z56oznJJnb3aoBloo+703sipaUa+Y8DDxqgLD8n8VymmRHIr5b+9
bsfkAiTtDwgLdXoPFKD20XnuIs8xzUuD/CHRTgnb4JmloaAcIZML0RS8hHUv9aS7
7u7zqK+RoBOaWYTxReI07PhaPrJADkyVJKudm2oDSX6fvu9e9W/hXInGRRVKOIaO
5W87U52BPM2p5ND7pOdygOCTPTLDiAbDyTdRkbQ3eUsdeOyyjXd4eUKYtMPYMy3N
q+LvZ+egIErjAgA2+tDRwNw8+xSeU/EF5/UzGeHfGFp/vR4jqSMpg1s/JNvI6j/A
frLs40dtkUrn0s12U0btEOKSye53DbYj8RHP72xtsLfEfW69kATs/ukg1qjqP/bX
OCEG/TPJtTORhS9i6gfwqI1MWKPiII0OI92G4sv4lT8Lr1p3T9ySmSt6JxvqDjmP
4/42WNBRGY27FMJwG2cYsOAIXfKJZxFCbGwuPVgvxmtPb4oPS2AgQM9G8TJ4BsrA
hkyaoGOtIe4EUDIoS670eMXURF0+TUo+TooY/+lyAiviUMLd1iQkU/LVCwoEZjsE
qCEyjZr8I5j8aBDf9Twm+21Bm/G3vs3X/D93SmBgpKWAdFkQwpT5v/OucxXt0FfK
JVQbkLf+8RYUtWEGWWou14wKgyjveA5yYXUivP6qisgiy+UKAM6CxGQ48YiN6C7I
D9kKN/BonpemfC2dJd+KGT9DI19mf5xhL3c4zhfqm3dKCgl5aXbaUQ/wMqu6wy0i
lXxkZP3nFA4cNLPawa7CQtn49OaQ3RfCcTES3IoZT98wPKcoW8kYk3r2gAXgZE+k
s5anDCrVCBxRSYc6ryEYGMhZiBw8UeOVI41fW4gloh2poVCfvhkbxg50dJpt7jOl
yIZsC2WDMUpjW7f8sRGlQHZtUKF72xkjVB1R16v4Ghd8vHmCVlbVjRoPwmWPADws
CmuQOq0nVc6NNILqIgntrXmQl17G+kUCscZGWPbrYbjNMEzFytgC8jNZcB9o3kON
Douh2QmS3FXVO35XMtpXSW5fz3fTY6HYOjQ2wjFvbNp9GnfEpQgZ+iLsVqFixD0x
FWqYjlw8i8IMSnE/lrZSYSWhSU2EpY1aO6l1jgxLGqjYz5mVEOSelG8Wqw2bZJfi
TDiZLXFyw6vpX0lEBlyB6u3XGMrqj7UQQlvxrpDb9G5J810FVIiaz+GvSTD1cPKy
FNFHTTeChVJ8YRhwUS2gzw/y4nBebN3yLeZNnvXbloQQh2PRrcY5cXF0gN432ENa
a85RF+mSaXCJUmExXKGj53xikJWd3Ev8M9ihgzBeuCn/DAbXJbII/5vBgONvXt9E
XuH9jpLUFWKWmZmrQDiCRB8RZHOJLbeSZq4i2+/EB13uKQbCDcBP3Zp2lLoJqyMj
3NoBAEXocsGQUUnNB2QQCeWtActM3ymmeWlcDgSIVYCHy8g5+cHQggQX4yjtQDVg
GudiNi1ufTKyxDFj5xI2z3hzybYzU2w1EYHIQp33jhlG6HP/TvgfsVac1ODSfpxo
yaIUaKettEnLgU2ezoVtEskohk+KNf5TQGA6M+KtDrLY+2HJL34LIU99Q7ppC/6G
HZpcfTA6FA7x4UyC3H2T/6TMrKjEQiurP4kABwEj8eVBrujanNIioorXQwH/Tba3
lxujzbfTeDaC41mfG4LcnUqgxP7MLVd37Ku9BhU+9cSdMKcplcJgADJGgPw7uK+B
WjO1hX53iYtVGDjHyUarqrjKPNzy+ILwV46GyUDuJ4BbHxTy0/8RkIh2EBU2uKsO
Qir9JDau3S66RYgmFtSNO3eUq/ZxBYsmMqCL3liRgIqeBo7gNvygivrHvlnL21IW
ypR12En3peCY7Ob69m2d+AOe6wuF5G2XI6awX3dFtN22MPGRG4KsBv+A6/C2tGJE
1QQc2dhkFsmv18TqXtews3mxEz9KL0a4YinS+ZLODsB/X2zrJIItsxwE7/SFMyhH
ZpkDUfYK2aer+ja1cqlM7FJ/EPoK8J6QWTG7OURiyJ5Jcsq9d/ksznPHv7f3UFjm
I4maAlGtK+HjAm5olKaMneir+2ApTyTgE1pBaD4z/YeDl2XM6RnLdsrxaDJZmesK
vYbq7+WobXGkHID8m2TuUirbmP/0VQGF+NUPLkX9QLyGi4TzwryGCOyuNcF6Txvr
LngOW1ds8tL9ZPyXYgAkD+tsTnmsJd5XYyjRweJaK8rlaUNjylfWgyf02VAY3/lT
Ccxe+GbdEUOQp5bjpespJ3icDeDPL+hkp9Cywxi3Ffs+fDBVO7mP8fJjQpKyeIJP
aHjAx/t0OqsjWTqYShRSH/zI3YAd51p8lwjsnYgZQpOOA8aunVQe+N/3kkiHa8Yn
LFgzooHnREaoOxlzeo9nNKSkTXQcjhkwL2prKXkFlQFd0WusTSotGKAtMT3nApD0
CXvBvuLy1R4SKvm0kTIaTlxAn4Vz0iynEJoWUVr+6Zwo5TbJ2G9HUFhwpRWBwXMb
QD9jQhLHnjD52SxOoZF7TcdVB5auiPdM2RjZF5G63eNWRxbtdlEdbhwMifgNo4V3
omQTLxxml2uyiC8pw8a0Jn4wzU/9PmzaBxcAAFdMm0B9hblena81qGJYWCUc/6j4
9ycvrL75ic6g6WH5UfY2PRb2ergfA8LeF86g/p++sjZZnijfrmLSm4pcqpjVzaUn
mabOWsxc87iF7Quv2GlUJM1KhRSVF5CgJTHGQIRqjVO8Y/083s8ooJHq3QqTVoiH
IqL8HRu57aFVPORWKEIktLm1Gl2IH2MmAU14SROCYGHcpCjJNAmhhubWLCsNcwI+
59/9wz3lw21RyljnnlhYGCTEJfx7zqAEiK29HVxFsH/gGeGo30zRPCJnYv6IuQHe
ri8uawSAV3BCEh3EdfZrpd5o6juK/GYrh5To6/gBweWsD0LgMJSsS3mppPm9abrI
d5PGs8k84lt5CkPhe3kjtcF2F19fOHdBIIYAKloYAA6MsjL2FXnk3Suv5UHfy/PX
bmxhcWWquMcQ/wd43k529wKps8f/cLt2u1OfMByMJBgJ7IkufN0zCMwE2/GGkqnK
Vdf9qb4cLFmffLknKdO/uyOhZQyGcc4EBip8eVxDMLQLgUxkGvEcTcVwCF+Zteh8
Dkds+dC1UHMwwd6zqwM5rv72Dn6/lDciMbI6aYkBbexcFsVvYBT7FAmG1b7pNy9q
OnuKSEJsV570eUCSo94Cl1eDOLzUbsil7qDp8Xf+EkLvaf3u7tSZkkrxijvIW7/P
arwfw6m6RWHgVVY4U3+IpKBG5kzvmcrhc5T2nFUDLSJHq1TImRFoEtUIi+wrvtLV
pJiOWt/1vvDcjhK5+2AomW0zeyy75P9Q0762Aoj7lCzcddCL2pLtCPhTNGEezYyQ
OWG8H2yJc3U3PFjet//gm+qY/UjzMkYP9ynegRTAwkP7ICacSH/1O6lRCkkGVYbK
8zqZ7YY+NYG100fHzE8p3XvF1B8K1DvxhJ/D+E1shtAfBzXgHIZZyQ99sZmIjHY8
+07CFR0xyk3vdRdx80o+HdDazDB8iUKj1vWStyLWp/J0gcK4TkIoB0nOSkcbWUWt
A7BgWvWHJPA2TM8WLEhmRMFS6ZpO41OnEjkxrahhyR9E80m3R6dwIeIx9hxf9pY1
sKjb0xBxEBxyS5nU0S2yRAxhyaK49Vf8J8+U9BjiLbuAvKlDz0bVUaCoKt1yt1kt
forGb0Z6HazX4VclJMGCdODw8A+MEEPtb1FljDVJwTkbLhOM0VYwNIiLG+dLdYQD
wQrWQw/nLRhwSaCMAN5J2vXItuSa0+sdCpl67+kTfMmZgjpaCvp46+SiZVv9+P7d
6EVU6aZkdRHZDMXwwa+xtV2quHYdwW6B8Zr11vTAg5S7N0tTz0bDfkyz1aZlnCOe
Nqya9Q+RPfuX+pOhUU3RxaimnTvdtHHpvJtq+1JgDYvvpb7CHnj5dCvFFcwZ0fqt
T0MhmxTquPYrJrb3L5VSZHDzWp9zwM2OQcd/ElDpX1KKeikVVXY+g9LWrAkbvrDb
plPMCwAXo43TJ1RH1R7nCDk02jAFhoabknrSunFJiMufOo9XAz3ipEn+dHw1bGph
aU+Hb3TggpVNwq8chr9hFEOs3xRe1lveFk4UzpzRlQSflC/S+7RObqLFB5/wZY54
64oEKM0AU+2TS1BeyF2yFCIFB+SEMkNoRqL0k/GpG9U3o7Q5A+ixPvW0VV2UdibT
rFKUIlxo8watxWpJR/a/7p8ZPPR+AzgoBeAYMaQNAJU93YmcoAPA0St2foR6n6H0
5CnjwrxyNs5QNrHbLXA1BRXpRaBwHG5JknyXIXbpUEhOO4SklKwyVgQ173JSGB87
NachYfEs50VadPUWGJizKVTVJok3QM+K8NVpT+kv7ki8HyYd4FwA50Vj46UJ4Y9J
0NvfpsDtRnFUQ+G985Vy/8dEto5r8AfvydiKUxCE3CdNcUhbiYP6BXYQQbLb1sMY
4ItFb6nE5mX3nDEVa9b2AfBVw7BWT+C1PNzHVBbo+WMYnTx4d+8D7G1gP0QySOUo
kPghxtXiyfD7lrX7M2dbr5xCTyAlzvjCnsesasHAkbtUxpSiik1zIsmG7Rs/SMdC
JxKojMidlkkNf9WfRirrIiXOumS6gKPKSfeb1QGsnj1QNbCKvJ5iUn5kLTUsk+HB
hJfYKyOEvAbuocTxNJ4z/ksp2bPY3VI7R1f11ALa/NRqVDgx48ttbFXhi5UPbK7f
rTqkKy/zweRtJSPYimJOqWTerTktlk9Nr4XdND+dQwBvx/60CDiaeP01jjebktIz
FzDoLdC1XD83pvJteX/vAdwE8ZfwDX3g5h1bec59XRPU70a1p79I+CFLWokNtJ1P
61urlJCyc1Orw/NFvkcZ+5ZW7OYLxf9fQepk+MH+R+uHdSl97mZHhyJurh7akAuf
n0dx21UUbYlBNFlvDnsCN6ctVUUHjkLuIzc6fsr63/cjKzAlkQ2WNf4u7kRYSI9Z
9WaKn5zIKQdBDZhd7KNiyW0hIv6ZQrsT4/YOo9NZ/Wf5T4a/vYNPEsBeAP18M0Vk
vgTIGnfXOo6gqt4jxC/ZwqgoecxK/oYi0pSHd1A04E91kG9JnbZLdxEfWjPHx/Z/
9Z6aJoR9NfI4KgCHTsaQRMXEJQNSTcPieWihA3QknwNUXxGxj9wKcvEUHm5XgduI
FFFMoBGYJmLgb74k9aUiwbMuByTizhYOT1VmK9RUo4QUptfbhdCLpv/9ve3vJGmK
S1nb+jtP+FIjX320Yw5Zx29Zf99806RKSLwMWfPUPRYIOMetlwxzGr05oBKPWcW0
6iDw4FWnty+H7yBJyWH0hC3WAIaF6kKRSO9niAg0iqLTcMjUEE5Dibn6zF6Zod1U
nM8BFzgSijDIgnnYi8LVfew0mKcs4yiINx5+K22GkIH/kgNbiRNnDep2AT6EfzLs
vIuO7nf/e+3PSzaG7zuJwPiSVPyGXYZ+vT24hyJtN2vKygvqWd0ZV0HQIZALRIw1
L9/L/w12JWRLPWMLcEzsdwmyPmpDkbWDegDk3zbyrcsGr2mCXCcKnOwfDenoKZsL
ydcoO5NSZonS6uHSlboIVw2v+R5VMjk1SAXUCkjg/SFTRM/pCYBT3h3cZ60cOhi8
cSckglQ0xfbtSpJoRzWa1/NmWZXmTU4+dGZxWjeLZtU3pEz9IU8YO/6Kg9lLWcH7
DX9J6KiSZHOZxplArnUs8Wy0wpkTeQ4MOUF5BbW6zYaNfrxlRFtxzW08pq4rhmn5
LL/isGbMeUSS5Pcc4Iq+xxFeogPaEf99D1ObINzqAU55JNJtKcqyHo8yzIop3uKw
JHoD6DSkN0UxD2PSj6A8Mm2xmU8ryYAdJUxd1qr9NY+GFfHZjHr0lwyavq8s1Esx
2XgJGZG308f9FZXKQHCv+4C3WtHS87JUUAV4aJdUWnz6gh4KCLQywct/II5/90O3
xFBxsL0q8+SBT7fFTBTzgqAKF2nmnJRWFpSQ/DdrR3JSxy5a22sxsMpW/Ln4U4R8
invO2S1GQwow6snZgy0oP8cBAGotBmAxapqjH//SQFzKfS/Ym9MOJvrFEEhPXkFr
O8Om0EOSvGzx7TEpGGSEwbRFDbL3MMKV9kTCOP00YAJbsKTuaobBbr5ihp5YtRUw
6a8pggYzIYqBNN+8lZygJ2fvfas6gJW4g60mOyJ/zyBj3UvlC+MmsBMyJicU4DVy
Wh9tzQ13BU8fudJosr+58USBqPvV6qeXE+udCWxtn6K7cNJaTaCZ7ICB1AoJVpuM
TnoM/FNpKfeWdUIJaeckZQ2MEeBNS5mkmZTEGQlnsLalH+m7k51rIQ3FnafhZKn/
WPZ6YIx8rRYGCh+fwRtHcqrRBixzctxHdKcXHsPiVkOjpRuQgYcSF+wpxvyw71OQ
7kHvt75/recz/l1Q2Okjmme1UuoR+G5nB6PglsiokjlfI7kYjJ3Y2VtgCNlRHyz0
2WGckPpNy8VjL1thfAPipF2GpvH21/xeLsgzsqdMAuJQ7exCnbJlnNqPGziWTJtz
UiJ/NZ3mngfDAhUsnVLZEXRqz93l9GDVgluclss6Y/g3Iq4LkQmm+J1cYVcObLC/
YkDYRGZdSjBdwP2QYXGBUw5+bTStq4h5HXvKWzHVvW/VBRNsOIVabHTANBA6aq2e
tydQYA90SABf1qCIR63el3uDT8OP+kPfLq47GC1g31mj1MVgoKClE4XiAC9opZUL
E18i2HsW/xdogYxtaCmYRP3lErEOMf9RwkRQAuQOnxxZuO9TL0JdEdUvxZe77uj1
fECAu8XZHlkHTxaoiU+JbYwQ4gXNhyE/eNVSxqFNFQysPcj6oTYNph1zIbrt710+
Jwa5XFrE9gkjWNvGT+Omaq4EfEYqAUsCpBPdcAtDf3mWvW7BcCu4jUgf5rU5JVBo
pwbgBjxhO5i/N/4PzoMD1UiP5DrYiwY9kwjSpPY+p0C4la4yCa8KStvwRPdyr9cE
NHhfBhuE/JHmlqlA2I6OkwoE0RYzseBhjELY/1OzQUAgpSStT32W5z0xEA70LIeD
GEzI0NS61SyfKRfUPtuZlqh6H/JRRahf2lWm8CW+sLltU2WD/3FNBmTAybxHu4Qh
fVwi8eZ63/F7GDdVabiPtwIWnObpYCOSMu7Ir9NhM4Oc52IMjJrqdIOAgHOq3T7O
56M0IiqQySmVg/4y1EOAi6B42J5z1lRnq+bcnB087wM2U725xURjPqwPofBWMEQi
MIwb4xJFP0H0X4Q9mTrhgImaFrqQ55+owSPG+GO71SsOOI59WXntVrcUZVXWrkZp
GyyMKoXO0jHUGV5s0IxXUQ5rdR9mkNq6P+MME+ZvnfWejk02cln7WS6/cLv5JFP4
C2S3XD65YxVgy5SUCyrgYCNXR9SMdb3LkjOlZcgVQLWUjnphLKF46JVeNx6rXUOc
7wDpV64iKc4Lt773atn0EqZGQkrfIZHMIIGKt4UnGkIT4/E+/KCWkjp5JgzS611D
dj349lO8hcScQmWhc0CT0ev+mkeihMbZiGfbhb949wsROJHOPtlCfarBMNm1TJUu
R0FtiOrkLMMbOzWLWpnJJBm/tDQvKRRBaWuriFYfGeIR9NwuNdACFKJvmGqpE5d2
fIDgXey2ZPFGEFMdR+fxQ7OiQpjUlhNTJddgPecuowa+4EZU+0VsLzcOR1ZKCiGI
BuMgAweoR1KAxuZamXvQLmJgIHAxVaA/UKozguW8tRxNk0CjuUY+y9w5pkJXRJfH
Jdu2ZSrprb6UIze3wN42CHzWBdxup18x7Lkz36jCZ0cB3EW8A3X9H0spR/oJNH7I
FC3igP8bUtjMS5A5Os9sCd3TqJ23I46imwF/ueiit47r1eMSFV019NIqKClAb5B6
RH16ZKw/qVooB6gfOniIHdJQi+UQItoWYYicDQXmbf2EKbOiiJikbCxk2cvc7JXx
xdEIqt4yKgEs+Bnu6a+kIwdL74YbTUtOrccxHAnjz2VUTPOE+XCr1yj+hyFlzmom
dWkixME6if/IWtmD77uT+R6rZrQLGDvauYmsZCQ4nDAMeBxGBu+brsM0G+QWrJP9
7U5+9sGqCjfQws4VuKjMYxbd5qxWlQXZ9FRS7ccnL+VVR75WHAoqxTEnCjo6erfG
eMTKIQxx6biSKzDPFVcnne2icZk7j5E5XErCfaoo6j90NjGp8Ft5zkwOZdINSnkF
VuyCrvL5QhWlCHNG878YpIfnQen4jCLJ57Enm7zdylW3p6Rq2s5XqtCr1OvISjbB
6awXVmty1qKLQI3plm2zABJ+RXVEagbe+BOm4R4FuUtccbvlJAsL/KZwMinRh74o
+M9ir2yXJ4N6A1NpcxrTMuX9S0ARWXMvVUkyPy1r9l39YbHtmT4emZ3RDxFuArnQ
bB0ymw6v5NwYXdmMyu7kGY5f5jZiQiCKD/NUmFohZus9CwzfgMrm6VC83mrkFgb/
8ehspAZ6yof9XREgDhM0PgqFyzTvDZnIyEbS/wt4nPZJlKaOUk1ZROxIHJRP0Df0
RkwsVKnJH6ENZwIWGbSoZvhX57FgL0fyh0MjsgphqdIz+mhpoEOBFZZBe3AKl0vx
L632CDz99OyRFdoWKAdqh+zqHfWEu1wl4XpObTXTHv9N+XYj1vOBVC3V7t5BkfbX
TtK+0CBVbkAUws4tgik6um2LaUZARFkTD9uGwK64fdRJNbhokTgSdskZcnsi00pU
MW3qScoA03vk2XXjCAhySdyjhfKwNKcpxyHw4gjvl35Ih9o2H52+2nC9+PrWt28P
qfr4DhAfanIWyS2ZbXEB6GEqTyQj8X1YFuCta/0OkWyNo0RmqysBw93mMF5vC5os
2FO6iZqaboe2QrDA6xUV0IeOu8IxVhb6N+A+RGQn2FEPKZJL9zi8TGVt33zKs963
uYEAB1D2NG0/pHbkYhjwDTzKtjC1zie4iFAHc7ZrMcxEzmexztSOdLHnfKhSWBlS
oXpx2WSqrgptIuu7VcgNSiJfpmTrRnCgSn4rE1YNZYuVwKhT84SHsMXxJEubPeXD
LMvQ6LFvicN+r76qWI2SWgzx0ZatN0mNl/bwLV/sPvQzkvIiLjqG4l0vk0gPJr07
DzYZ14de6+5eTlh/vURhGpipU+P7UE4UF6SPOApDxTKiVqwKCVduWug/MgePhzf5
JbD2J3UlmIT45RKAzESoy9hoVMsviJcveyCFJrMZimBFULOg60TSi10BTWpwKG/S
dhvU4io26CUT7c/EKfCQDvsiTTn8WsKqcHQtHXGmnz1/upGIMAL8e9whx0J8xCnB
vMKcwCVGyY2+22YZwYadyiTuni9YxM02QdnpFpvd1zs5jadTp0hoh7PaHKDjqH3x
tzbrRjoC9nN9hH98UHxveYgxI6n49kVChrI4D1qKMw2u9bCu1sKu807FMDroi9i/
rGYRnqvzVctJEW/48BI5jRMoIxG3czlJ3DPSw7KQX9zAKGDBc/Srm9a78DNWhsw7
exRVHY5ZFhANkZIh4vquO5hlRvucZXz5X1t7WgRmRfeG4Xhf2Purzy4LZaRJB9fh
voT6P5DFKadvzmefC16G/bILCc2Xle1gqumbUGVjtgGOczeauALoI+olfIhou6pk
Do9/8yUrOiHI4wzDuDr/F1KzCd9tctddpNChvO6VWc3kfnqbRtJiW2aQklc41HdP
Zy37b9Mt8BGI8tr8NwA9vYCChkRg2SQekQ7zniHAzjVgKvrYXEs73R9dP1yIU6E6
ii85Q+KWralTyNAVmqn8HM0jBTWoOD9gM05QKAW28FFb8cIXbfTQO+Qc4dSH0ouG
4U16MQeObS0BsTM3bWPc/4DBuXD4DNebVtXbwpcUeRfgeMnTP7r5c66lipK6g/kD
QqT54U0f0xs5slydNxAe/UyadCS2FBFhNI2EoHkfPBtgZfWu9gkpS0+YcgXHTTnz
CEb3hNS4LE4hhwTk5dry0p6Xu3McKPJDPayyuMHp+Tp2M5dpV3+kVJXpwkhsZW2V
+GKXONIXjg4YvR1N+9JaaKo7pWxAG1l4F2c6+8J3cdufftzPN1f/xN2hoP/WKls0
PCoXbGQtN72t2ZAiR4SOydVE/eMOKQBamYzVVjVqTooi6vZ3FU68pb0SUsKMVclY
Cl6hmfXFhKCwgghzW4jrVc9xQ0BLrr/Ak0gbgInYsQwS0ljq/os4VqEa4o4kMrmz
2gSdpzT8tNO2TiFn87iAS/sDIUyVnLOXVi31kEtNpAfOpozw7rmovp+I679ZM7Fd
xjQSRYYZPEAAQoa2etSKyjojhANRNu+srW5xH69XvwTL4FcDfNPcts3lFsuvs90l
tOrUFcpChqoS5xXdUEymWqbY6i/2TUXchxC+jlgrKF4R192d/AYgrjy0xlP+mmmU
4Ri4XA2iaBeOwvjoUT/u/hOyJJSQElUC/Hn97TkYAUzvbVIIUIjj6kecQoJA9dsS
L7QhHD9EwOXHdvSDRfW+hwmJvUNvs1irDXTQCbTQwhx9h95R73NUPe534m/M8vCX
Ndk3Os+9lZIAnzDezfYcYYFv4l4AExMUszYYxTN7BHwiRmvG75WSYe+gSW8GJ4NA
eNrDoQ4n1+mrYbUn1cpslgz2ZR4P/o6cAvbPGnVa+C8hVH2nMWs0zXgRzM4QDujF
xMOg0U78WX+iqJVTMbfBMhFMZeaqBI3jWFKgnMupMKqmaBuhtlAU6Un8aLVWDkAD
Nkq/v65ZAuE/8NUDPPXlADn5CIb/G5yuCIX8RO4gDP+Zgw/htkKGFY8huZwNpEFF
Gg0aJj9BjQx/FYypm1BBs8Ao8kCqPDPaoOt20t2uF7+TJ/hm4FzjNTaIoe/p2qRP
YJ9nQQlv7EBL47oHAuoKrHDrD678VETWEhxbNi2kBTYt5wCrlAVO8oa/rnVdin25
lFZBUkUXJnhVnE9XW34SejbCE6yGd7F9TJ3eeQcVaRKlgRZlj6sUMhS23HLaUkkx
LWIVAxS4GqzeXKKpqbYUjIUxpcMa1gexvz9ICs8LTXnZzIXu2jY5aLLlSCkDoCIp
4XUXlY2H+PjnYLSyQXfNsr7sW2KLGyTrBvf0Dq8BIZXdFJ3znaiYprY5tfoaRLfV
q5W9usQUtNTn72tmGOflWNvBrKP++69xi4TU8PXqkoAEx/uvsYWb3rQFnEd10jw9
jNsE8yb/3Hp2U35ZU8qKsbncLRGLwIRX/i/19bmpGOrjuD9Fdw5jvnaifCvb2h8D
SkrrBldI34HOIn7II8H6Yj1yA3dqTjNExhcgsYWbHH6qtUNoZFqJGcEEdurxkVHa
jwaSHDaBvCwljWfGZzOg0gdhtCLZcxuxoIEBoID2r/saZIgs2nzYlZat0otK/3X7
F31loCiTII3GDFYzyUhBUs8DE2/7pD0Z30DwdjqAcbwJ9p/eiSvt5/i+G/KMHT0V
nbKF3F0VdvURWWjGHszmx1wPZP96oAMJxklsMotjLoepcT1Vu7kO8Qy8eE2MIW41
xK7w/qeUxyOz8DlZgD0iwImQ6ZXGheH5dAz0XpmEHqRterz3lvZ6nffKIPWGX0RM
Cuv0+WsKQf/7kTO5BHd/vNr249+RKDqsi1i4F8RjTwPZrKiJcpMq6c7IrgYbTM4g
AKHusiQhkXi2himii4SrWsLmIdxHQW2lLmYWEoo0ZgfOSNWemjNg+zfROKWT7r/w
DojXchO0ZaRM4VibpvLRTOsfFJcQ+xKfY3eUmSW209GXF9P8QHKv3phz6ccBaz8o
FlI6LJouYYSJDWiK8Cxyr2jkxVEqps0BqJ5FyYBlboCKULJ1k5e56nCgDvtP9zv2
I0Bxh9zVM8gdz2ytvhRkadsrlXlvqTiu4sheqQSCLyCgPK2S0tct5FAMvVn/C9KA
HnsCh+2jVz52WvlBOJ+Cr+LLYNHOONtWOnB2Tngqv4+f2T34mhKnXYwf5de52nkw
yMgI8jDCtUSRXjTM0heB1pC205fy8Q8ljk+hu2kpGCFzGrNpoo/pCcRhiPbQVar4
g2dM+a+DRdKU10OxFlLSeujWmpaY0uTmDApC+Pz1Yd4i/ymF/MGJtKpfYWZnnGle
NDfxAJMTvN1ViHcsmzyXM1UE1UnT9TuMwZLqtDHwWcFBiXZyJXdt2MP81WDEXjoH
irOBHnWKOyB/rNz1BJ/GfDTYsXPK8Tr2ZMO6utTS3m0p1u7+PT5beFUdjgEWxBNx
llHu1RN6yw8jTwEpQlYefJHP7g5B3uN8Mm2A+amngMHlcVdrFQ6OwdM342i73vgf
0YX0vSISFraLUcE6McH/e+6FfkkkUj4dTqhmmPsKROC4R5xddMWPpqBtz2GCqPsk
HUSlhsCVmFsLPpAM5AvWYwwi0TRrBRj4DMLWADi7z4+IkaZfW6UgOyxk268rsa42
HSAYlHdzHHGdAl3R2qtUzpsBxKc2fuIMa8nQXlkL8JZouTUN+tGLT8aFfRMfNLwR
AW7shGnPGsBBSfVm1lqsWYHcLnuaxbYqrZq89+blpuE5tn1rT2405WbPLIvsQuQX
vo4mU50D9VsemyeTl1I3RKQ+izjqUYCEhGmAl8VzhNNfxfb0adPTKAnC1kMwL+F1
0gQw0kpWAhvBZXiq+CXoO38+q+hK7dZemOcPvspWLNpwuKte6xa90B+udBcDjNCU
ZH0Cn/QeS/Q2iTGqOwXodIMscslBNvLc6l/gNfsA2ep+yXsROZmIfPEkIaurEVvm
SNBOOkZCN+5eKq+woVndQ96XA+K++3FTHbcqFp86tG4wW2XX1kKMtYglMLGeVign
64eGPp+VFhAzb1cNGDfGKxHJS42lwkyUzW/wWG1io8KeJbzXNgjyOpIHjhX87GfH
IoRQBYy/eyKq4Yz4xagJsiDrm7abKonw1KcS9mu969LdSJ59aOek8Jx38fs9AMXW
kBAoxx1K2RjjNRUBUuk2De1k1aRsh/i4FuWm+rwAyYHl01Z5aBkdIltxYHLhkkP3
3WNuuJLJmt5wuDbxwVpWOupTxQ79ws39YJOTmUL4GKgmI3SDwx0VoI8IN2EDEgo3
chc+YZiTgOLy5Jfa6+MuCULHuDRIfJG2ODCC5MemTbIt/IgF95ydErmXmGFRmWUY
ibvZiiM7piMPCKEa14to51Gj1kLGXtnXv/hoy3M0QGMlAr5nw3DhC3VXQ+Endj7H
MzPJxnWsq31wF0asLgM/u+M1yDyuXVNkjzuKV4g6682qko5EjnaGU6GjjiEvnxFP
UKTTmy67zSWXvQssDEdXM23Dd4+d1HU/LRNb9gZwnwfcdSokd3mOHMkYe23Lmwna
YdXbxdYNIYlfnn1ywarimuLs98LNT0wqWLpiJwXRYZHzYRIRbv1hzrINUI6Pvvny
zx7IXvVdEnDxiVI+H1sI/lrYW7FaSEd9BzgxRz4LwXftuDtDA2t9tCbuQm/O4AUx
NFiOluhc6k4Ri2mrnYfFQLR0DSljfK9tASZbmRXhAaGvh7toLXRlLHDESt+rGmyH
InlKFfA2fL4iMjYcyL8lI63WSuzZIHgOKmmQoGQO4IbgI38gqk/OwP/Te5JF9nU7
MgLCLIehXPGtf+By9VFh3CaIzriBtPRVmeSCmktAf+3J2+m3D1ei9jF2gIAZiJWE
1Xuh3al5GRXBC6N8uTnfT9gf7KFiIdYnswQW+ooUSO8sf6yVb9hFQAsNZ7Z+F/E9
xl9sUnm39D86eZT5PE0REqMweZ/Omt4HQvVYjKNuBbYUhKftSsm991695Pg9nPaJ
Whw6dUQrAk/GFBL549iX6X59RuLzU4NieI4+EBzKU35Y5vsq+kzC7KVRibtsaGMc
zeETY0rkcB+igCXVMcXEaR5xThjc3tRUT2dgzEVBfp82hL0xVj34TNX3/Av3H0r/
kLp7Xj+rSQ3Kv9D7yvG89erBjW13zikSkggZykO/KIFL+3ZrEViALopqeUqlGWbK
rbZwaRJ08IE3otdkJS5dUnCWbnrzlFVgUOZqiIVlsA+q3D4ug873gWzpjNl2mfqj
+tO6RsSa1EFv8wdHDXK5A87iz9uACyGWUBWpCIyue6vGde9tU7Ef0Z9TzwUykAeK
05E63j9NVQ4g7O2Pzg54YtySBlYP2x1i1WG9w+WXqTVlRMQITfJLE4ocH3DRFcL5
g9YAsCJ23wtk65WZUzWaFSIJgCD7te+WWW7EzVEGOcNsfAZkw9oVnj0fzVmJ/CaK
JBx7i4k0DRzsWlkv84EVQ9fQf4og68/12btY6nrHeFGOwpIAeR3Tjj8LlMWpUxdH
csixH71uF1BrBBqYIxBJCKi6356SABcMYP64gngK1mIP/TyFyZ5i6dcXFX1CauIW
yfhauVNIXBNRVvira14+XjC0lcQQDKlwVZbToJS4+Us1H/cZBiKbX0aIkL8TMOtg
Y8bi5yo3TuCzNoIDfz3DJUlZ7beODUcKC5Q4ReONoGA0bk5BmaQIxnPjtYEOou8z
+huYFiws9s1DiqcI6Pph1GrXnTPaUx6rTGZxvS7u93uHiCl0qSgsCJ6ZRZJDvRM4
rBfQ1w64GUmzgTTzz4Kyk4FvKlnpB91oIX5nBvwSZ5xr4iTvW+jp+9rLSvsCQMpG
pmeiGpmx4gXmHOfY7F6YkvyPWNGlFzdclFhRyLRxFNYd6scYuG69TttR/cDOzBTB
hkOcaW2n/jk6Q3TtgN1GJKEJ6xEYISlQFLPLM5hG/gVmBGrYNqucPmO3q3LQcjU/
Q+pR5/YK1MaBFA6rmSseTeOFtk2Ldq3Gk4zgZ08bqhYYfxflSRjSxwLtqhwZqD4r
4u9m+nD2lTQ0zTv0nAttEuEjaQ3ThYLaneNc4W7K/pYB7et3fjVZ4pRfdS9ZIelo
9VjTDo4P1iXGMuxpAvacy9TrU1N2N/ICJUPX+cePnOGrjH+hEixbMzGtF0H+LIlI
1XgQUIiDuCoielzAdTgidm+w3yQZypt2DL7X58pOEfo+ahE/S+W4hHtN5PFfy2dQ
A5sqrcv48lN0AhEOEzMToFvPdvFkEfRP+epNOmbFJXCmse1J4wsM7tP0SnGIjLsv
M2RLfmcUr62gzK6mA9ozE1eaUoqRs3S1tdVKu4GYzfaiEhaqmbN76ChHU5BIpnaE
Aj8t2GaJwzg1pc3oXoJeneJ0tq+hx/wuJmQJAfV4JYes1ywVwI+YhmKtCYIG/BIj
s6k2eVpIs66zWhTH2xIG7B0hCSCYveEzrA8NFzja71kICccEHKgoyfcR0r0VZ9Su
4uA/8pouqEwMa9cZWk5Vym90ixB2/JnkYg4+qAQ0sl3QaabGjCrk/4YfUu42pv5s
pe6BSbMU2pOhigAAxcqs2zdGkb4B218FQTowuAseETkToNguG3iLge1corfIPROw
PN49zz6R3JHzVtbADVkVkL45yfwuUmKfiHPfAwjcKmjPEP1PEa+bXrFns1PH2PM1
ylsq42gPw/eB9/J8StaQVpBYzKD3Ty+36hzsg5FfJmDU/Maj1QNlSwkfN/SXY1N9
f++KNKSY+PQYGHIwhIzSMpfXU4aiQ/uQQzTwUuHzTfxWVCk1qQ/c05hITak6UwLZ
Y1Ud9Avey54kZhC4vAVBuzBFUyLzRaS+q1nb/k+mcqKTMrCwDw9p4AFvy+qy0336
40h3Vp6Vv6cl/dfBE5Zz9PgyZcqAnx6k+Bc8l++++dOnWTAZvaBcskYFO74nAt5s
ZWiBwmsmvOs6rOe/dxb1XPk+R6eDn5TYfmF0YDhmYYapwj3k/zcYyqLF4Gw6VWVE
EZvmy6juAXWvD56j6N7nrNOIsj6qSzkmFwxhb7Svxzdxbiw2oXwRdym3CuVPVCTD
o+uHbn58iomlBT/IXkhhzFkd6+eo8wDjMyGdsbngTt07vKKqJnmCrc94mFG1I0V8
DkLPl7tTKDo5veBODjZTRIoXLETIQkqYq0NiJwkxL9LBReyiKgXM/cFmd/C6gOO4
/j4wogPdlkTCjmON50Rd5zWp+BuqWQe1O/yj2+VAKjapoMS3g+6DzjDWtLpdK7G+
o8ZO/qSvCWaXNVt4B5wrRcZU6PLr7tFvUD6w8tDSjfbknip5x4dJg0s5c5w2HMEF
u2kYnGtf6cFpYjSvYFQyp7Eov1oQKcz10sCsqOlua6DSr4pGZn6OqOb3ROqDChEQ
qilXsz0+G+wV/Eo3CnjFSh1fQUl3EpkEAXjkGJzxuzj87lQn1+BPWb74ztEe5ocD
FBYICUt4QaV2N8Wxuxj0OAspaOhfJgFIObs1DvelyZuEnkU6qZZTGuxk3KmGJl/x
9Nnx1mz0D0hFIscoqRenuw/aXpQ0NlaQNBhaa9Q6NXr4vqxyY9V2mihg/pTolwhk
dZXwTD/jNe2flbEQiJgKzkCYbNVka5ynIrQZZjht0N+ManV6gj1jKsUMC3dMHneD
xq3pHVa6CFJIJ2c5VcvbK2FEVZ8Km4hHXM4/5N2yOXv4F1+I95DvNERMf1YcLN5X
pZN+rbXv2p/fFSywbedT/ph8xEL4o8zG+Nym8IsPfVE7yAt9thpzps5QhCAU3Cc/
LqYH7iShiaB8AM48SjZuxEyag10Gl3gK3x+IK7NaNixjmr7eWBk2cEIY5LE73Dyh
ks5UwKeZxrJ/nMaDfkEjhtZ9tzequKun8ptQPLqqc7RSLtXeDbdZ5CBd3Qwmizz0
i4nyQHEbd03RHQo3f2EIRO1GDofNqKDlrU+pYmQNXeFJvhboncgawVp7barga8d+
7EOGz79TJGY0g7Nhnp/BHRQ8+RKpXKlSlxbETvjDV0/EP10zuR8Db15rmIBCRr1v
I2fG5eFtUuhalWEK0iMJDwmKVzg9ZIGGhViBcDyYYmQOBZSnre7p+3pPtvtObObZ
2Pw2paDZMdPxp8uIm00Vq8u5gcuV3EdiIghqApbIcXSbWsvKMCQxgNdFlx8UoYzW
S/3iJUwpyEuxCyynxjS3dZYS9qmE6MhCiraJTzjmp5FxoMbhMmeAEF3friukuM/m
NPLu86F3/oPD1Yjkib9X07F1ciqFZ/KIsYhEeTrMqWYeDe4wljSGSb3xlloMoi+r
F1TZhm9QEYIVr/oWACWS5m5Wd44Hznj5mUP7hhATwk/zZyoR1TrCzxHv0BHtDZ/2
mOfmjgBmeW2QTRvidfqyzeQ0N9DjNdoRoB93/hd/dv3dcxdWUIbFFPxneE3pmXur
BYoEcm8G7HRalC+nU3cqw4jhj+qlR+cwB3uaOtap0Irh42gmn9rxGWPK2OjdN1Xh
4X92byAc0KTZtNNLuYZiW40JAedJj79bG7T10C7h6hlPXFaOt7zMUyov+4ie6hZc
oKW1gq4IC3/8Od3tnMd0gdS1QEuV08tncQUU6fCW2D/w+9zmhW+FV5YVYgRw9SRD
+5ZDUCJHZey3uHLOfRsV8zR8HOxKacIIDXz2hBVPv6EY3yxM+r4Qw/k1YcdzMC9f
rhgFmfDOoAwHSQ6aRcdU3XV/ma1zOftU1rg88LPk70TDUqnDo2p2otFsmnZkAi/v
6/J7djr2Xa3K8/MIcmNTO+/+gXo30JcwsjxruTdynRKiMLFX6B1u3W97Qljdrmct
RJClOhUCnlymaFf6Ljd8WwDd0jweaRF/n7uEMvTKl70BAeCaEC7imskCqzX/xWFb
EGtGrErp1zxv9eQ4KEnXa6fHlUTHI8E3jdvG6OQQV50y6iGnRtzTTQ0MtjCYmONo
D2iQkxN2v90cc6C+Ue/UZUK4yzHWHROgFRyCiuN23ysEfn4f6V912f4DNPoL5IoX
yIR7NhiQ2hkSG/IanHTBV6HqbE8PwPh3Pkw5zRAhdfYXUEZdRWawAaSD5Vo0L0kY
C4RO41EBMrzY/C5BEVNSPcENfykt6MYkO1ydWK3x4PqnlVC94v7pluzISKUaJViQ
XZM8UCfBUXgM1IujtBwD+vKj9cGn+jZSMti51qMVkRNq3PSSbn3+BmJET/oVvJUY
F5XWgOrPpgIVLtAHBWMFD1Wd6ji0S/DQUJr2UwiZePlC5I8SmNne9s5qfzS+C/9m
fzbRGT3PLBwj5lgl8D5JSm0LLu5vgWp0XmolBuIC91PdHMvd0SFc62FQf96Z3vI3
v8xRnU2qmFs8EH0pLfLjV5tHWGfG3jDPtVkUNBpa69TnKE3K6IFr0ZuGVdYB5OFF
lxtxelqmmJZ0kipyNKIZmW+9uIZbW0oLGrzY0fTr4YAGvjmj73hjojfOCqHKDSwn
kZ1mZFEs+AJQxhhrpAO/tcQjOYPzR0hbh7GWSE7vl+iIQ7H7PhYqx50Tvc+7v7zy
vfiUiDphhLXTMG0uotdYMk+KeC+XlY7SenFJ2JI8UdQYRnSYeVpYUoCWRXK0xvLz
3bPljiY/BbPM1o7czbgt8ZoSE5LEkWXqVQLQhoax/7slM3hGiBWlpfcU152nD6P8
ewse+z9qxLeL1cHT0FACx0T1XfD+h0vjy6EDwtjUVsNsXm6WXJi021cGpVpPPL9c
sMVy5RPgrA14GquaOMVy9poc92JGmCBihQkEUZHHjKKr+22ReQL69t07gBlsFUuV
ysjVC+8TIXqlAOFD8ms2oJkG0D9vL/E57iPFbHTEwdUjh5pl4TKYjqdub+BQYGqU
leYlorVUPiuWSAw2kDvQ1OCHSraLFGEq8G9NMsxU/5gYHVObKFIdqIKu4vzpFxRL
/HtERA3xnDgyXRrj0BqFQK3lKQ6pxr+rFnpytwtaETZArJtRL+EbEijdKhHYlLrO
J0MW7zb/dNWuxKHDNDGBrMXLty7rx9tVo6nBfZNuuzC9GfZDJdOcSJRRgSQf9HVs
uw3JzrjpsLomCJJ44BA8wcFcFkI+cemaVh8vdY5+k7fbWZpYaXDV3iY1BOtw6VON
u8/0wSOQImNWduzzDGY3L4bUeGK9a3lvgsQ85svWf7C7ORe9Bq96BMV3roacMGyv
2AjUh5i0kUFqQ1VRktBVwZY9vuFnhxTQUsGcLCrGaO7FskZbfpfvkmzQc6uH8Qmz
BxJISHC1rtZ9/NVwlfswcrpUhwvtU3p1SgycFz3ACgCpXz3VXCVeuOln9c6Xpuf1
JFz17Djg40fffQjN4nSMOJfTf2fcfvrVKHVOhulH0PU61xSBoaiN3wvjUJzloJJf
8QmCc23B2ZmVU1XBe2hILZT2igu7indlHHqqdBfmYYGeRl0NqurSeeyBW071PCdW
Ij+Ma1BvX4v7Oc6ky5kO+diTfhwB40TD4Buc6ag7TfRpQNIZ6b2LZ2eVFgrmi+tA
Hr7HY28RD5PMS5PY66VpNEERIKTMqeSCWYWT8eYdZjLncJbkgG12oKMG9Z5ne2cJ
DRFyxvxMGRqCAlUnz8mhbYpg4uf11KqrBU5pjY2EGossPk2/sI9id8MWRQ/PUQve
nfU0mn8MtqyTj/09yvV21cDU/zNLGESbXYApyH6ls3VWX14/vNViACPgcXTTemRQ
yGenN4T28vDd6BezvkNxkPNYz53R77jtZciv608/shz4uQSXqlWGWc49upbTmq1O
4rrXXqLYREtdmvFGFA079552GPvFT594MjSYdEmtVUodncOZtfesB0HKbAGE2hX0
uai6rIBGz8+kk/3lnSHnOHkgMUdY+7kGRJ4IStF7Wxc+jnfoHalKTY0AAYKyGums
udrgBwBNwNc0MUN7LjOxaeJbN9ANEHk70hQlgu2+ysEw9y7aZLr0dYXKgeMDeRQ3
LsZc6iVO1ojVHxF7ZxQUunU6+3M828UH3rTm2M+e3dHrw8vCbCQMM3n6+gXzfO/i
qfvGA5tgYB2I/JRwCa5XmNrB5m62Oc2ikra4KmUfT57I4i6ODVo/nz5NmOBq57Z6
sLui9zJxL1d2a/j5S4BAdL/TE7QVIiKhgAZiFE7HayelL72MWahsZtiFsN2Ao8qz
hmNT54UoZylFgQzfNsEb2RzL7qNyBteYUKJBoBjwApuILqDFrhMf4HXoAU2xs4SX
H+y0Akz75xFGxEYhekr8LSzFb2YWpvFOHV7O3wBCTvKaoYyX6UoRT/ZQHty1hkco
wYe9sBKIgnUNPKLAYbeXVDn/LwqcEDJtsCcFWzzEQqEwUdCkFl1JpwDKZMSkbq2M
L0nlJbZVQWTUVU+fQ7+nCsLzdgs/aMOtz5dSpNOSk/X/PWfvk3wevQgwR4/4+kI9
mBrj0+bFbvJmMUFs5ba3Tnx4iqcDnN/YfnlN+LrRVDOWT1yBKrCcoy4+6b2ivIgM
PatM0yFhPbVNggIRJTcHkRuC+j8vmMOS1tulsmVffiecaQqvBwWLBT9xapRJVG27
6js++0gmQ0YEPnEf/lH/JqqLltGyIrnqcSskfFzJUT3sjDIfKJpuUmKhfiYiUssm
zctrjlkxJbyc7X/OaoJClCkIpwFYv95x39Z/odCAzfKd6I54LFAGvBFpJ8RFkWfE
aZCNwOTXRwFCyDDiFLCOh3PLloiQCj/n5o0/z/FXEe5lB36PmrqM830zi1zvbus0
c8FPYnNFB6AW3hcjXWAmT6xod/2RE7Z9OUziP9p9tKkJryLwl5G7RvgwD1aZMO6W
7YzFBvCC0id0UuuJOV5aYkIHP3ioReAMooyuz9qKqmc5h7XyTVZt/bQWcF+daeRE
akKwjbXFu/8GXZQVxAFelwdl4ruWCsIQ6Q3M4k4LBzFgS9nIg/rNroPdbekTYvXa
IPJa7n6Rw5wFUydR0hqKjtm2noaY/XZ+pBTwrhxe9svmzAJwZpFFlImI+qJOsXIT
71/L31Wy//lr7xYuHFnQa8O1zP9+IEZGJaTwyNwyNmQ2cl2N3V4QtIUJn4HHT+AC
MFEH//tG3Uwflk3jeWOT+1usUiXwxTVVZSj18m/H2NOuc2KdTXAMBD/OkpOy0h+q
KDpwBfWeDtVL+mySEiUHr4Lu6yEyRKu4yGiThY5tZqjGtzBGfmy40U3ID1C/W5No
r+2xoAGFXLZn6YlQjZlc25dK8i8GIS6vHAGcPtl2+AS9Hih/avgLP3mrirtyy7gA
PDtnn/Lq3kpWU4FWRHqAUnBbY0LAVl1TaCGxuhr+QVrQJ8ymw8C5AAwpScPqwTFS
Napoe6IMb95oakOH6oKIQf8LZiVtwQAPX1s5eHtoiIOalHc/AchNxH65KE/q5RYB
tTk0Aqvxxs9c7uezoxuJJCNxcvpGJqqXO6Ulb0X3zxYg2C7rq99tSRktAjfojHcF
Z1i6F5jZJpqOv6Zro8d8y9oTUeIh/DYvW4IkLl3gyUcuirhXuIzpmGh5A+cB6Ciy
m0v/KxkUDvj+2YeW98kTHmjUK2bVUEDibPYj8NNa9vW/cuVqibN5Sx353ZFAUsHc
iG2wkhqrHbC1oKSvESkgyFdvhdleqrivXGDtgZV/QCzHPtoaUFZHwC3bUVJU9z2q
dDmbJe1MfGiAOG6PdPuJNQvLEfIBon79nlg6O46+632n6O9CVQNvjmQRHX8CLRWm
0HGcVjLglHrsfX7PAA2ZzcLhQsQY6JCO3gzCeRDc9CYO+vRm7+cpq/hzzMBdkL18
lFDDoSBXjgErVJ3LHvqVydKxn9QVpF1x/VND50G/U0EF3KHkE2tkTP3RK1llnsvL
rqYndQaJw4i4YwDWG+UAyC1yYgqI6gxkEGvjAQe8haTe14dfG4IHQEf6ustrSRCD
+/Y/v6WSpLYaZsjjt8XwRnzkKbzCgBXytsCp43v6TKKpljvwxxnVqmb/EZ5czbKn
xv+bFxA0WrsZilkPpnhD3nrwdNl06ul0Rk0tnFZfQPZR3EGE9nhAgHiIWNIBNJkr
xFzo5PzG0MHzh4rzOjRefd4++DqJL4rchn2rLmSRgELPbYeGSn7SgwTLwNeixutl
sf+8xL7CqXftdTBFoKuPZYqb0N3J7gvFQFA9KUrlTnWODzaaPaeAWkL42BqYNn3K
XqW34NCDoudXAKwXqLKiaKaW3R8MgPI7NmLYxGdbJGwtOmkIjx03xZDaDdkBYMST
nheuVCu3Kl7FhD5CaO26VkJfuGQQKZtzsLI8TY3TryqMAQVsjPZ1bHE98SwThVGU
RXIe2mjqtNjtoqvjREKaPLnUVUra1TglzSWpuW0CqBSD4Cr7b0wfidOATzsVE6Jj
Lew/2X2h50wo7S7QR5/2FT9WsB+vhvSmGWbhNNo/yHf2nkOx83RyOeTKH5aSdG7g
G5ieBWxWWfr1zLM7xnkMy+EuwKeN5g6FHiS5tZDLuS7qbBPhhPr69KQ/Pukcr+Xk
QkBN+5kDQ1x6J4EPhQnVHcXPsWcOReTR8RP1dpYm4Vp68QsdIHjEWSCY+fa5gOaA
b4tVvLbaruc37ZaNF929jy6Ragm79OS7iNY/I2biYiQ3j/NBAeGZZdaGjdRBevRe
OSQb8TKBXErZsPbOO7tukYSdq0CKFdTT7bQMv01yRLvx3NFNaJcAkNyEx/xj3h78
n221wt+CAPYR33ctXV/8B9wiVLTOyrrzmNxcMVXfAOwmmBENYGkW0nttruSCN4AH
5w2Z06rjXglnrNfK/1AvDaOS+PXLgD0UsiVnqtp7ITQbgMH4ss/prsp8cM0kFXM1
h3FYjh3BO9fcD35cMb7D6g2efuOAo2goK5Q7vLDsuuCfDSiHMPd1mNoixq8ueezv
yo/pGksdLyBH6auqBVV9DdLGUkwsZ3rEjykkj11082PQ0FQ10Rl7/y5fYVTiZ9Zk
k4ylZMeEesOWMm3IjJocPFKiCdcNAxyIfiULyHb5kp5PcM8u9Wo26Kmpu6dwVYUv
ZeiyLpjHCODzXnA1v/vFDjv5bSpjd8Z/aeGN8PfKH5Gp2bqz45CVTp1I11xfu72i
LKtnU1R0XxrlwhhVqWTjy22Dw+GCjKyGogI7j3k4jyRRvnuLrexMDYs49+gd8/ZX
e1dJu3muh78IgfcCh65J/NqeormpbjQhz2YjBS/R8qz7i2aHalz07L6zzYnh115p
mjFI+yyJl+kn1TWBqZZlO8MoFsgW9IYTazT9rXeNDwlqlupKeLtvijl7K4SN3c/+
azHCltKXL++ybYkKRKZyiJdky/OefzsNZuRGfjtGgOvBLpNk6VF//+Nh2A/50lnd
ifdyh0zENFNCELQ/KzlBuyjjWC1bm13TT5pmu8fahDGPiryxECa7vk1GwIK6vWNK
T57QjVpINLuz8Tqn6P33KTXgUm2X9MumjZcAyIaeO5DASdqVfQp23uPt4J1tzTcd
BHreL2/7G8oJSS4+fKS3mH893pIP3GHiCiF5Nzskwmii6L0vDBI3OJux6B2TwDc9
m8vAc2gxiPUgWRY4gAqBEcY7z4QhNgPZ0AMi4Wq48hdIhZ6QEF1g9YbtdUkqk8WK
8i8Oparudami0kmIV7z1AWjclG4+84JhWIfJCOVYR23kJ9egAgxt4DJa06RCn7Wr
/u4z//nmc7QQ+qo3qu1aurGfuG5Nx00R2ykVu+2s7m34oT3umSHhWTnOPtgzF0ya
ZYT/wJwppE/FupJEK6zkxiBOr9ikHaLWxBBnO0JXnQptjIU0zLIqT1FYX6hu2jf3
FEGgCowKG5Eg8YbdyzR3O/76YS1FkUh0pL7HxXINbIlGmphqtJp5Uc8WHBOemTbL
cqy9ank2lWL80lf6m7vVINCZUCfAdnqw4RAZRlL148xMVfHFgDkXd8+qssHo84ZZ
CuK/qSLf5VfSVcBFSswFgo2FCyMW56g0A1/mgf55WC7EkQycksfginMbfPwY9O1B
h6tf9DMmTOnTDin17wfwKHuDjff6Cuo75IEYevm1fR6jzc9O2tdyzq39CJTt5dxy
+zEuI2/6ZKkMdlTGjRtvNTsG+kuDPGcBz/P8PaIS0XaZO1CJUU45lJypsm84RIUd
3T0UhENrZuuWWj1N4BA1nPq84uPVSkyUT+4dZXJkgrkLVF5T4pOrq0/4/5WYhdAA
qgkgTP16D+Kj4gaLCmUEM+AkUK1Qa/ENinLUQq3/BQvyzHkLq62lEWzG7/2j7J8/
n+9qjKsOTFUFlK6lDaRsF/L9zAKp7Z/eG7lEOV5c5Ar39v0qx8L05vjMhDOMENqp
gOTTT1vPs1OQOnOJFDOwUGxI54Vz10DiRIkT4jNH16rlgWxXxW2t3fMvQ2aBwyXw
yWa9ADA102ZTcbSPzPSGyrOj2hRvtdKV94GbYL/b6uUfhiyWm7RLdNbWZKVyVvRp
cgaC80Etk42iIJH1RdyFXmVG9WETQrFh5JN4Jv1J3gOzvxP90wQY/2oQbVxZHSOF
oMaPRVWOT/ffGJU7wd9szYS0BsCSY33pjqvx3OXyOePgS3Nj8zNDbZ3O9aPZiKhZ
VdFVZm+52IbaqDPYZ/8NLqfDsB/KJSdVtIzXYCoNF1LNdMgwPAGm5Ss09IhNtOrS
NNP+cGW3o2Sq6bkd+TPeprxYWhYkioQdhDDmmzFAZ7yjHLdryMzaLR0Jbj+flhpO
CwkOVvElFoYaFONBuG5kClDRAguZE8WZHBawqTs2dUC4unqIv4F76yWiAaW81ERL
Yt6P5tkn05r8gYZrH/q1d9r0m6sEC9wjPDB3ywzveQRDDwDQyih9Tl6Q5nbZpTZm
q9K/0Vy9MPtgboTfg/t83ij2VsjKwOMvlVLw7owYA2mDTJs6KS+BHBnx1A3Cxqvp
EQKOG4Iv885YGM4cjCfURY96fXEjqtMSjARFO6BGlZj4x5t0ABL1PB4n7kJ41gkC
ahxK1SVr4izq0Ql8KF3O7Etv+2Dws5jHMJZDMiTISjnEJk/dM27gP77GdHdIMBEv
ZmT0BP8uTRKEu+rEdArDZA9U495V05wXv/ZdIQhYF2D4jyNWKb6pffTNbd4gjsBf
N/Y1+H+KAOGz9x3w/XcW6MEfOl1xmQI8LNZwJXaJD7199Ino3LcJUupn8CONeIMh
l78ys1VBgWXg6Nn2eED/TlaW5zwxQvCk5AawOZwUHqNB0hIoywfua82bMDuhDDfK
g0cVsiVv9dpLI3Z3E6xKLcV8+D9vtleyhutWPLP4+16dyk/E/1d33NWsIJ3/HY14
9Wb4wB7r2WR2elt49HhFkNcCt7ZBccNmYHf6G8RSTrs6zjqnqXM9W3vT1Ben2voK
Z8fZg/QaSAYyCC2c8Ye71wYrkXE9rCC+vpEEkmfS2k0wuD/6bXeyMmb9TRA+TCXa
2wp1/MjQ4+txdDgD7vsiv4HbM0wU5imaPnG0Nf2DpfY75UQlG2OPRRy79Z7hhYWK
wZGi28CCJCj+Gm5EyGImhpz12EslTyVT4nC55MlWgztgoHLJa3JzrheNAwyCO70H
j9JEskrPowEL+m5nD+tA/Pq04bL91FIQ9KzKVSL92HoI9FwjkKcMXHxNhdTZcZZk
i7Oq574UiPvgArm/y/ktHVpFIzhpVKesYXsVwWqNl3maS2fGhGetQzz9h5w915Lv
8gaWqBqgPlFVZlg86DfsT+x7e/6s2wes+z5Ge/sp+vL1LefOXceBYZiVyaE3cWFp
/MhSt3A7f6+i8PDPTKwQlUP9EsgO5E+zROsGB1gwpLnP1FCSz7M04OOxd4PdzJNJ
caLe+FwWeo7aSVeioPPZVmUl3ooXKRZqQdFQ/QTmib0LFyGPShKTRgILA1VYreU1
AoKW4f1tG07Fp3ANECZMmXfgU9AfGruwVzrZUgQoly1RL4CCCCYKLR5e03pG7C3J
rddk602fH+4oz1mZXTgve5QaWolB7jqwgF7r4KlcwWYeCJvxmd+097FeufrvKNnD
xVt/4fLD07wvcEd5/4v/coeJgnWoOjWMs4nckc51l8MJl2KkVsNiDBY63cMUAiX8
CWh+4d9Z5tqMKQwQvZSosn7KUgHqXitju43C6EMPBQdyNbVCgcOYy0j75SDmz3jq
0QE5fWW4OqbCnFG2GM1QTWF1DTTp8Dy2gzLViUlqXdAEMmoZKb9nI1a2VEdx7NTB
8zV81VIbG8deyNfHvqYVO71U3b234jLFt/CSInwgje9MMDQcbup904AtNaTAApVQ
NxAvCzgHHR5MIunsg+d+CY9waQaPWnQO5eEHKG38bvGSz9RuF5BjdOtHDF9qY4Ed
khWEoOLPcAHeSK03AGG8GBYTyX4phLYA0HwGWAwLZVZRjdMg3j5YRC41/T9Ry0FC
VuX7QDOkqcYVyx+dvr6E2U8em2NMbslDlWIuU3Oub2jg0gO1JhJzzEYqEW7+0LO1
AqW37AbP+kqX3e5RZCo4y8WGvg185BBwc2ocbARGIRo+xbCn3fBpObzi3H6DbDUI
FJoHCRoS0raWRbpFnB+yZ4QYThaceCoJkMxuemxYffhZmY/JrI5MAI0ByrPH8zp5
TqBKG52JihrL1+8b9ynJ+p/SbGH7YFPxUmQWZa1tnoShIWO2NK0StnE1a3n4TjG2
HfIVCHEECB//6rri38kKovrWILwonp5iCKeoSy0ma+lB2byFwngCHYbm+e1eUUc+
1j6Mv4BEgy5Tysj6RHLeFMPtc2XW5/dYkpRfY0bO7apCKyjEf5A1WoxbsjsWpBQG
3W/z5mVJIva4FpoLjJ9t++8p7Cw3GL5/AoBhaDoeFSJSF7gn6Xv6F60yOoePxZGC
dzFLqfRfIdjrvVBru8ShLGyfVkn/BAsZkY5tgUqb3rloVPPsDrW6oUfjbuMVkrud
DFWPEKq5LrfXu1as/kn9xJPHDs0OzzLnQSVfpjmLbZCnUIN9cWvbn978kle8Apj3
TxzPstEsGgXTD2NRkKoEl/o9gt3CODI3yrxaRp2E0LQyUK0v8eB9KkVRyZXPeR1t
wQe1FvmqLibu9MmOmSbwmG+uTtX8j90MTEGPm8E1jJPeLwQ4IzjN9HBznCnFtiA5
n9/4vjRIBHVFVOzc/jkZ/FsKb0gPOarRgcJX0FriUpGoCPzLH7wVzP92Wht5Ew0u
/Bij/UOxVu6X+y8lUjlB165v1F3+hWw7OFpSd3X6l2rFyb/oAgayToKVBnPJfUi4
MKXT2cDECnMsLjeRFxAIf8syK0H4URTtafSA98dJc0yCOmHTKbFmASD+NicLk0vf
qEDMHhRvZsguyKYzhTkmsulWLWQLqpgKSDG0UXKfQW9WRN1jmo9j+cUS6l3RNQwA
WwzIlSX9GhI52uleNqIWzEVWq/6zb0nCT2rjQUxkSaTBslOIY/4ORbg2qnfRlMb0
nqSk4HksDerUjd3wcCcLK+xXpfHaJ9g76M63yrlIwmSpO3WBqmerKD9Fiz8KOG/w
ChJUUU8Wo16zx2JgHGhFDjpz2kyMPKotyXALOt80QTAZer3d599+33Qk1Mrv3owP
RUu2as9culfM0BzcrmAjwEfvu2/pKB/B0HwUa6rUJVealWzDVsJ52W9Kh96vDPFK
iKn6iRXa/tW52b5iIvCKPkRlM1t0eXfUzNr/iF6u34nc5zVCHc7PeyJ0QO/XH0+R
+AsBQcVgWtSv87Oq0vtKQzUcx+i4HTkAGVs657WeT7WRq666JD+oKrL415SAcaNW
uz/TZQdvAimR/DkV6MAmD9DBs9gq7ObXs+E7tnqriMXrUQnn+bxzSj4XztSvYDgj
F9z0BVRKd8S4cTsn76OFWO2sMQH4NAsQh78/gsQwXBwZENjl6GOwygrLBaUtkziJ
8eKa9Nxqs6eyXJ2iDTiBu330Ib1LkobzWlWV/8rVHgEKmmy9PRVoB8JmRTvtAaGv
ZWeR0lnmPO3Fq+TsaJ52Qg5JhLo/QN0r7tGexq3+wjnJ8wth/01Z9l0Ptc25SvFc
0VdZYnIr8yu12h8alfEiB3+tXynssaSPSgUl3cIDkc0xQUuLin9NzA5VxMqu5pG7
rlmyClZSyfJltejkgmIvr0Bw80pYlZKov5cDSKUAO+a6i9sl9nXm3dTZSyt8eZ01
FFy3bRDg8wBY536svLOAlRlk7CHWU7yns5WiAdrhvIoT1ZMBr6G2nWLkC6R4s2h6
kyp3DlVzHuahfcVwOHoycbbcRA/wACVqL1uaVHKJ+MA+De1NHJK2axl6024F8EgY
TLDxLJPQshX2CLKHP4YwirHjLHXETIXAyHPsg5UkFYeop2IGcfAYV4yIHSZXBDX6
FoUGzNhnIL0xAbJeR1qYbrfG77eEC3K7YaM3PpBSQANQPXl9OSLSNu9ng8xqaLQk
0STQzHkRzVCN68nzTuuASai4LBp+7fAT7unVV26hoalshbZvJuKzPvKuWOdUqT6d
gCROZMOVLz/0YU6O85EmK7bryQo1SOgI62EordL7qc9qtnm43dJWPor+Y750I/lz
FrBt11U2YJ+POCmMrdNNnbCwA/pRmla/LWNhLwBHzLWwWPRBy53AQS6JLOL7F8Ar
xS1o7I4kb6JyDBSxlfhhZ5CvB2NHex5cfk48oKEYM5w/tJ305TRoocFZvo8F5oa0
O0f4RThIcjSGlKm+0bie2W7TTOFXXVQjKuP/ZPs+QApNnFHgHE3XouwIbjfFoCwm
ziAVYuxGdaYRYKZN8EQEDTxsCM7ZMLFR/iQcNWWh+YGzoriMhRLLrPhu3oRSPHzc
cOb8TvtGLvvJI2A2vwAtH1ViK+oONuTiub2haBNna9muNvE3E1fPBVdpoydhnY7J
IftCZjiKsOE1eFB2k8/fD5L26McSCTECEAToi0WudU5ZWHri11Exb81N5q6yZJRX
B2YA2QdjNzpz8nLrcDhjiYMpAIMuyoDfsBcmorBtOXqU4l4VY+SAYldsOtp89NO0
xZy+0Jszy6SxJGlGQDvYMWOs+VYIXENAl1S0CByLaC691Yu9SXs5W3p/TorgYEDM
HhjLUYi1LWxnWTIH5cAPiPdnW8YJwUyUHxCW7FO/8y519bot1FqRxdm+VpPgcsIT
m3t/Dzb8+SFXrfaVVHz2Q3nihqEXwDTM3lTaqELCsKGlJ/Mp+h/AhFVD9HtFhoA3
r2e4P/Dqk+O7tj4CXm3Y1yjU+ZcwSM7L0vQrnhHvmTRg8AxHx/v2pGSuHNv/vs2b
mK0V9Nk6uK08fP3PvY+QoXOFtutzw04mYti8iQoBU75RJmlFvFRnsQbiPVFS/8Kf
QY8BGHZ3xu8xQM7L7sdUuZcMDeebKByil2lWcK8OJGLNBbVEC0dmty4cL1yaCOO9
b+2fGpyeiUd6pROs2nX54FgvrzAnWNHBTxhffJkiMNxa5rfhaZZU+I5HZVre6RmA
+aQPA1V6HO5+CvYu9Pr1CWFQHjTbsvWqg57oP/+6XjL4PKgLLQX4u4+yLcS/vVqc
+B9/GSY1TWfN9vn8KtRTFhI/Dyu86mybHjS2cXrT1X1nMqhMTpxcva49z1D72tN7
z5pcoNCORhNhbglloUX3YmY9O/L32BJo9aJFut4ESz+02jFvKrKmpLTYIKksZuOY
ErE9eJ/yPpaWEHlxE2QdeVSXC63Ol5cL+qqLQveIB9doC2+k6r2pI0suvNSk1S3R
uYY+AeQRhe9uxagDDBAvM95kIBeLat9uXQYh4ZNnagOnr0MXgN4g3Fn9/Ygnbi69
68+jEfWiJp3COXWvwpb7ULHPtY2/f6/+i3dwH+xVeW1qr6lI/crK7c+riP9FNKuf
kVxwrDfuVSnkoGG8O46+pweez2h+aasoEcYRLFrrqP1CANfQmMSkfgnCgq1PTa9D
/4d7NgwwAkD9Me51UtuLOfDL/7cDkA1hsdjPoI5YoAZj/gD2H11pgVRbvatnQmbN
+7ZpOqOBuUxrF3kQ8noujwRfDAophId8v5p/DgOogKRm0vLtzoDMriFi/Ta81EvZ
AbMIGYRajzHqmrxVJx1DhS8+nBj0lMsEtb/+XZcejIEz1iaURlITmDdXH5L3LyxP
V6QXqMYjc/mN4H2+47CFi7B8mvnKLI/BXGyih2Z8i8b/4zenwVXA0/rSPhS0KTen
wANkYxK5O87ZYQXhck1t3gkWOg2M07ysr2hcZAyV5/89HirUDRL6i0dtrJhQD8cH
KDgzRDIcX/zav/KHZUk7l7I6+r1X7WUOSV1ArhR7B7qSG+cGYXZp98f9dUVHTxmA
OUlYrQy3KB+uU2EPXrvjKsFGdSPA4VDMxbH6ttnIoGf8fJ9ufokJsDBJd+lcipdX
cxpDLYftE4N91oeZYUzp3Z/70PJSF4Mz30zdrN2vI6MCB3SwWq1ymOVIINqsAYat
TH6RPh7x4rTuzZaiBWiqdccPHRr9heAry5tyaF81o9emQ1I2nZ8VBzDc/1M6asfh
YRVcYMnTc9p+REJrp6VhwnItFFr/I5frXAdW+8hm6JCQskSwX8o9sVKlxTLOQOwu
c8EWWiLrDmUkaCk0EDeOWfytHxB6As6FOz1olgAjcbThw2LAwmdvkrQgfVe0IO5A
UCdK8Vs1WVu71KX4wP5eNJtAYGpaGs8oNT6rhf2takdxJCIFAwwiXW2wedQXUhYU
j8eCcLhAnUGc4bPSpFCHk09nAjbFDEjcSix2n1jTZhF7iPMF8brOqGZKdjQOJEcf
xgtbE709phPAvQ24ISKx0wMlgENDf4Z09+v9qf5rtWBHdSm4N6GoF84+KSpZynJA
4F3g3wRnA5b1eT1N5HzCl7cBsckRisMQ5hDg0YIOeZXlcdiZAk8FwowM4hIpziWI
wgt5bqRWpCO6pnuSYQl02KmnWiQkS96yrGLoqeakqaC3Zqbf7Yez/9yYXTpEIqkN
0dOtNfHiwq/Ms9S+pmgysQZHoZRrdFUwMeOPFGzTZy/1CWv1Mpp2ps+8tVw06y/J
diZrgAYydbji6j66bmH5N+Li+9DDOpwUhBXfoB8rn004YlHYrFrZSRoZxBrTYoeT
o7MfddPGXdbxU5Nh1BDoHbUJ5t/UukPJMuSEnC4B2TEhRGBLQoWjSDEKILBkNuoN
xV0tuuR78yAdSqRgPJvW8jyNglPsJPFm1cTKa3P+6deYbytpHCZIO5kEuftjC0R8
ISE9npUuuF8M53fb883NgPShNkk+vv9CY6RGTjdQXZcq4G22TDUud+NLBa3ey1sK
+drfMqG1V1897+660/zYpYHPaYJw4c9Ey7s0qT3vKR0aKFR6i8Y878rNaqNinVjs
R2tXd8t03yglE4JXbuF76MDQAz5kvFEML9OAKM6D7NbQGVNylP1Fb7zhP137C41W
O6fGVqkS2FZ+PvpoV1Zkq2q2B7FBZga2Tn+xSOCyulfoLlZ/n30qygjJCln1oHLI
tqfW0OVltCX0dB4Uis608V1U1FmPg8/4I+OsHE+qdW7W6w33a9MSBGsqEZxH9KG8
jOnHCFHR+iH9Gn5ur2fFv7OlVq6VNM+BYMOBOuNznvT81cT+g9cJb76/oAcRc1sJ
OUGqSW7T1aBS7QnxojsJfXmtrdpcm7b3Oqxk7WVs9XlxMhMwmAKSW1w9eHmghPol
ZvEC0HQbNvLE/fuD3BieZWqDzoTkyOBW9Cp5TcnwHLC0l12At6eXCNrlJ585jS2F
3KtInoh/qSMNIVdu2HYSOTEZMB87NpavhBQAd9WkndyPYZOvTYOMCK13M+8or1qF
zK+oZyRBHQ5O6nqyAYpE30sAh9TTXz88KSNGjAyyrgfqmnRhOZ6cFmVzqfCmdqOF
aaeWwbQ7OCWDP+C7uWCcslg5r7yAQkSILCqZCVoOSomxn8Qq8t15Bz+83MHsCXhg
WRLqOeJIV37nSAoyxPvuSM3YT6G2aUZeLSKQB+nYwxLCXwSzsq3HyTkpA9+QAa0c
0i8uEOMRv8lY0jCpbMBHHfdRoPdPbdKDVuhCB3NW/XVtr9luv9Ot24Xg2ybFw/fj
6PlIkqRHTPPtyjDzyU03T6gU+bRl6vyiQrMfJV7KhNP5FvO2eig8YwIruv/R00zs
xNnpt0Ij3qaFAs3gz4kPAGzzNjHtExvxkJl99s8y6bY10YS+QBrtSGCVTfoZPBe6
UiL+tLhKosJDF52VgcDs+c2rKG0i4mVqc9FAiyHzJh+n9A3f3uS07lPo1aeUeDTZ
XkSFp5KX4sdy+ltazvjAMylVWzx1n6G/h3n5wr9e9wEjM7fu7aiyf/JfrvwCCowz
k1Q9XJqwxCtjbVKOi8TyWF4LwOHhwxINthDuB7E4NcQzuhpBbkckVhM0siMWk411
k4hOTUCJ316hjGYW71BCOwLVg8cqhg76jKJu9cUXM+hex0QH6eOyDVUfJJm0TnSm
S5vcf1QZUT0TYJ/Z1zuQTkiXuaZnK2TNzm+/g3aKanQOqN+UGoMe1nGg87miCK00
fDRMR5ZPi/KAiGg/80Fisl53/Oecjkjcn6Au8lMAoCLpDxVzjj4GMSbYrLcRwe0+
9qjXQGeKRQPnaO81x9k1Z8PiSur4ALL/QCqCBR9Ot1wNSyPeSdx7SGCuWeY9aiSY
guZuw40V3UxRR/LvwrbWmzAnadT7QCfqDMQ1Wn7FSynCHgnTUE8R6w31T1cz4+BL
AMJDMo8whRPtOq14z/1lkkJwTZ7nfmRcrb3EDVloWsXnWF2dvYSGV9Oam1Be4jF/
1xEWQg7Rwd8iIe2q8u9xD2P9T6GH4NkhjAhdaYKDw3/K4F/+ZvZSJKlBOTpA2vOD
k+Uk4zfTkemsCOFoav3E/TrlbCxT+5BjTOViVo1PamyWauLcM1E49+0G7mMz0HIv
3q7SPTCLg1FmyjRv7q+J9Uobt2MFTG3zqJna4b8UO6oJKK7mRRd8EjNdaYAg7ndS
DRDWivkUSZyaYY2KHdovx0av99bHmh/tA/LKBJP7PAe9RAY0Q6h0nmEdVLzwCXYE
e+CC8jmvG4E8VIi5yO2NUNctFRFta/RD033QDt8Fep78xicdhGiHg73UF6t0G0Tu
mslSettRWZXg+NuMyhhKCu+Vz6BVvX43Zgs5YBU87df0VJXe3cIM82pWZwdB87H2
gN0lggeEFx+Q2xhI18RNfFpJHidvQqjA685xajbdQmUEccQjsFcXhw0P2drUUIZi
3CBKmGsxkPP7aAByLL23r8XlF+wxO3t75Wy9yQ7tRprcS3hHXUCu408QHlRjnLsG
SffVbGhqXlkQ/r1Z4f7UZCRDagjoP6lp0BBTuLtxE09x9JlaKS+PMvLNoLqg0bhq
TNkdIhObD1xwcILU9Tv6EaoJezv+ciJs8s0tlNzXSxnbPdCIFk3KvMEq5SY0D+uX
vvhkEc8Ef4Pa3V6zJeAy+vJBEFrNXcrJlYhtAwvQ79HbHvv6iEPlpyvWgCiUUzDN
cAcZLA1rworWJWpJNKmlRnA89roDpp8/Nio6MMH0hv0+1xBgSssiAJ57+XJC6Mqv
oWAR/WEnCf9qR/3lApp83I8nW2XN7r/4D1bus1jzKmdiaiTDy7TwOMe8jLxzfa/w
FEBH4VlWZA7X0Zy2CNVN00GizBFrp6SmrdCnF+dkjPrhy6RaTZg6mJH/zDq0e48U
tDqMETrtz2voeSAbraUeHXQ5pxtasz38kH/8vG4xT8ZTarM+SSa+15GcHUEWfSyL
RAkxDOuvgxAYx5eYEG7PkxSXFgcmzhBxrrk6xbnFFP/wFj7lErT0qWcD5k9bfe23
hDWYVeNsb5xokaMmxODVdSp4qsHbEZoUroMWJRWUbeUcsh0GrLFQJf1UhbWyb6dr
Kwg7iAt1gvxOnD3QvBipRW+6ElHJm98kITM8QIWV1YYpIpsF2YviZbHZ/L0V9Gt/
/rvwnpWk/jgVGQqDi3z2Ua5EKU46ohDiZLxQcNK4OgyrLRF2Dr+F1Ve6BCOfA4Mc
69VU2BA4j1Rm94Sc5r/y1liYID9NQHHPAYEIgh1sbB1xOBLxCpyVCgNlLhaNSmHe
JBvj4fusTIRtBDrl2EaJDxXLVlp9naZpKvaPDmGz31adjzGkUSznSNmLpqB1i9KU
mVcEUuCMz5AAXMKiBVDPYVpkBBrrS69on0UpIQjQMN6YgHqzFcjULX9eLouCOQrO
ujlgDEUtAkaC2XZHkdUu9WAiwFTpGxVi9QAn1NkkX6X8jox7+lb6XNzB5t5zdYuA
4ReKBkyawy3mZKl01KOVi1BNPtt0+tAPIkkHwftB5SyVbg45ElbFnZVMgojog6V3
2P9K+SnHIaxAAxltpoXdEUz7xHdDEJvOe1KE960TdmVFhYtomdxeJgqZYV0cwQW3
zYFvpGEAkxLH+Wu3YAWFiuazWIe+SrqfCJp5QPzY9gruVVjoylzTYn/27mDzO9HQ
u9vggjubMSdqrn0ETCjA1fFRsKZKs7GtBwNw0zcizPP4reiapVHBXqjmNa2w8ZxH
lMpGwP+ZuFOvQk0sij94I99xP2h0xqHyJijux7k0ixOdnTIbQsPAt2Yuy4WcUyaI
2wxJwJuUqzi+E/WGtSNsUxRcerXJ8T/P5onRE1QFQxqlmiYyw9tu18Gu8ySf8zdZ
wLbGuSQiZajl8bcOZPGWfosMP/ms3gWo6QeDKxUnWEhaqM0I80EvFwD72r9gzJOs
9d6+uuuYA4A79Qo+hXckPWeOq0KB8vf5KpbtKRxUuXLio0fwiBVzTyaRnFyjcEq2
woGrYWbGH0CcI+y9Orpw91uEG5GqaXLClDtUTm8lbjkOfbhoMoC4y2MjAfyxi/f+
MoEcuN6coaWDCYF4zynumAUbApvUVEQzeKJDaEK5HrGMtbbpeW5qIkk7D021o8rF
JevCzDDdwjqDZI4ZgxdneyIyQi6YfJmMDgDTgw6cGcgSb8JG3YkWrkDjS2603VXJ
uKy++U+FukBTDN7iW6k6u/FzPWjrqVG2I83WPVbNz1Ph4caaAlkFFeTtIavooVhy
4PaHN6I4fu5nky/dOytCq+0656Y3gH9ofVfURaGp4R2CHxsK3PqDWieLlcTQJjvE
tgVSK84AvqqKHNkqtVhiYLG98cKD1yrru8S8fS2uOKXrZ/JPR0B9dUaGI+K6Np04
0WTfTFZkod9lAU1/v9FS5GiRukeiKAEHehjBOJ16JTDaxqnmriMI2EYZ+xNZj/bR
gsa+d46zm6iocsiGIGNWYMb8D912cXX5ZXyXNgNwEYRpM727ExvAjQIRjpTq14tp
5DD+PCR1d73eTzF3xXnCEBPN2HHsOEn1LxvrYAVhV/2Gcyh9c8ivKEHUU+7HiH0W
7AxYNgauVNMQf+Tsgk1AIKwV09F1cnozZPxrY6ZMEamXdYefb6JAgqta+huBeXp/
05f0zFi+C7Ld5HduPn793q4Nl0tVBm55/W0P78jjvz4aUW5iAE3gcRiU+Fc6uYQb
3MUHmZi8JjzwZUALuV5ZUgmPz0a7yBUcXTgxsVjylQn+7QPVpIypRfomjimMtvtO
w2kdUWbVZU5o6NGPMAfI4DaOeNxWlnsrlVSLKMYvCqgBxekISAhd7R8Y2XTbeWOA
65vGv3JXlQ+yJH8FUoi6P42jAjeFNOPMfdBdqdgw/tQSHQhJ31c/mdWhfqhNVrtD
5AZ/IzFE1EZFBeZejp6hZ4+HGAYJeLZjRuSO2M6BoE2V5OJQPZ3Roc3/4B31Izh3
ijYC+eQHOh5VoYEFfzDZ7N7AQiQx8mFPwndghAM65yVq8DtrmZ8Ax2Ckj8cO1qt5
gPnU9DT8EXGSlNWTTtAKVh/9WcaagA0IlyIsAFMa77SdyKVeo3Gy3g5MSXgm4RDx
zodQZG4+U5B2PYGOl93ZrwSrsKFis9pNR8QaygwPltDXJsTwXwX9w4u8pOUYgvt1
DkNa+3q6SE+BX87t2tbZ+p8aNbHVZmwIVVnNwhP6vZzsmnCb8jpE5RYP3Pmnlp0/
q2fclenPuHoMkv7BtGqElmtgVXGMQOuXWPGt6NpEG/svPGK/ZnMBT37BPwo8CEjN
IlwpZxoFb+3dJV8RGIiv0IwOhR7iM8olsUJvBgV6JsxLS5BVmOz240+dYeFF17Nm
1xHqJ2v0tf3a2P2fcYoKEXv+bwCbPtarKkCIYo9DvjDcKJ778IWNnqg6D5AGe1BR
4TPQvbo92JgjxZXWs9y0p/hMCI2Nrta/BwP+8+SDzkxfWfXzQqFoIRq3oYvH8ont
PdqVNduo2gTTE9AADzWELIWnLKiTRWND7KRwn6whvmCKQIXsoD8XXWXVkRHIZsmw
FjpHeZB7wTATnRiEAwaI9suxCdrnmKGDL4RNCCOaxZXAvOBnD2LqILFekDQTmX6i
V/iOTPWg/kgT0VS4AADAqvTbG/cGp6FyPO97ODIdxY7r64SGOifsL8E30Pq71Hm9
BQv8hXrd54UJKrnGrmwFvq6zI4pGpYbRhMkjJ4e0VoTdAKlCt7Azz13PKjmjNlL9
cy/Wd7bASkKi/dvzjdi/8Qa+SmQ0gweHGCF8f/l6CylwTIDfTfq1qqptqVLjf4oo
SkiH/KCFIknuCekAgcU19De5SYjQlhxL8Zbf6/MOL9+JWi2N5nrFJoAz31I2dQFK
7y+8udEkHTbJ1bRLliX2xfdnOIH1zBUl1uyUs+czTUo0FPEJ/0UaWCVf4Pc9Cxue
EqTulnVPb5nyplG6XcDjvVueX366qST+u8NoXlkh6eNuhgcp4JnDWmaXq9XlNwHm
yb8QCIYWOykEb8pN3d0KS3QvobqwVCSCatK3ZJNI30EcZieRatcUgNdgqJUtcC6G
NN83jyV9Lpc6AGmxjc7CPoXX0maMgbOgYSvBDLJSJBtXldy2yaKjnGkDBgQFnQ4A
KDTjs9CHAVpk2eUFE7D+oYYrYovNFpMtxhbFkDJxiyJ5TKEbDBDO/vJH1omf78Q0
gPAczIskl3pZV063IvjzSyZ0N5Pt6OBq+NnXUScssVVbyZzAUdifKUBlkiHF2piN
Ah8gX8he5dI6vNo8H0KIKVho2wpjXmiovrPQzcfcIB0zObxe/IIVMzAkXRfoyQZZ
zHOQI8KVN5P57ZYhJaMCXiQlsEdlF0EOVabzkXG2G2Wft1lt3yf9m5N0dXBb5Vpq
Ti6bJAHmyIDFJZAEM5zpFJOKxXiANROPIbK0hpp1JOEg5AiFTflJiYhnmgse5Bum
APcA3MHT7rIaQ6K7JQxIB0gF7aAdGqe/nWzIKsjsxpC25hmeWtJL4ljLXN7SuwoN
94+o8dtFA97cf4f8XQ9Un65cKnnvrVqQPYtGDMkKZQuiK0FGMZ8z6opQmmk9ik2z
FFwfFObTEtbP4IOidUDu89PEsbYptmYITSIVM2MPh40ga/n4EssLH56j4oQQRFZy
koTYfuOH3ywElJk83bNnF1Q4coHEScav8K/KfeiA7xlr5EvkhLklW6aUKeBTACzi
r8IZ3XoSxZWx02BCOkMcR7hAMtwrPAoMBV4XBGIQ7SUzZMlq+wRl9Ivu3SXBg7uC
uDlaSPN0DMZhZE0N+WH3KozeuaQMRtpYb4o2pOCst3OdMcHA/JlVsGVI2GUR8XHI
YYwhxznzq+ESUwP1tf5bitZjF1rEYnvrhcWTBQ1g778I0SC2xC77muhKpAW9/kEd
pQmZcm508djB282k9d9yuZF76ks5JOZOXFIYlylyQ/Jq2eJ3rdGxL5b9clMiaOey
WqK5TGtcQZhobjrcDkVCwmKBNQfEbbCCkMrR38n5e/zvYG7r28FYIj1VnDpOIZrs
DKaK6rraQ+rvSiZZSADBFXyut1jI1Hi4UToiF19Tft/2QgMpzptVSCMFGzV8iiDi
/pR4foQS7DTOQsie2McGcaz5qeQ0SCX+IqcfbuPsCfMEQjWNn+yF35g/QGrpG9hI
j3uI7Uy815ubXvr6vaGmFWHFr1bFZhOal1FoZD/BYytQUCi07jiBvMpokBosKQlt
BEWLJtwDFw6h084f0xZN3jQNUx6n5yH7UvghEnbnifZcT00ID+Vkg3nygenAYo1v
fmUFc+kLAlT/OAKmWm6o3zZNwTYjs0DBj7HCBwJHoG8uYGxhjzeZaWmq43bH7gAF
0AhSyqIj/yYOkBtyxeV+UdIFobcZyht2Fa9Gt5yF0jhJPGMu3mRgw7GegPzr47r1
1TagtAYPbXNu3dl5QTHkvCjEnD5ECulvROTi+GhtlkOOO+WjP/VZu5u2EnIJMz+w
ApzooGraix25MLXb+dyWtyrObUKfdU0IEbPG84pjK2tC4z7+vhru/zpjBp237sGS
gRHDXldeuPs6X5RFNAPgn6ebVqjGc7TWiWaXR6MkTgjBiiQw2Mn0ky0B61X9bXx3
CT401MRvaGBdlnqEjLA1T06h1NlasnesBE7/JNJ58D/dunZCYJC5LBYJ3g8Z3tME
qmqS648POWHXanFICB9VXbEm1IsXIGsLukDFKkKkJU/W+1dM5lCvLFOPvrRqjOkw
hdPB/DY+xkZBaVKgsKg+UAEvDLur0geRpIzRSxYcBsR8POmkqGXhUz3hZu0FeaHu
Um13HXkXNCtVg3s5TNEgCC8RZ3FBNvaVVi4JicOi9l3tDWuIMTaicFLnS0ntD06Q
46/HS+BbLE83T+EwXCtPFEzTejf7sO/Lz9+8m/G+Q3sg8AtWOArVxabR4PHw7kVq
PHUL98gueCt6TI15fN/deAsnVmISTBIG6kc13sHlD5FlwJ14MYy00qXp/0dyVNQ/
TNKATXuB0RO3lFzEUa+k93ZbqhA8jHU4qE8GeIIZKsGjnHwojQVyouaE5LrDKbUE
8uJQiu9ef/8jfqsvIwB8Ejy51zQM0W4kifwA7yKYfyknjYboxqfNjbkShU9en8Y4
m4FuiUWDQPvtwVkREv2JGF4SDagMoz6RGUzdZUsX2VqF4Jr8uogSLWwwWHvQpmAc
hwHntW5TTX9tc+KMjqjSx5GEQhQKgjza7khdIplWsuP3WlJpj42L6n4CHquREy15
8rQ5KP1g67wtNErvJiVPBkQ14GTyz67MsqDGRKa68JI5rpQK/qiy1648MLiOcAsV
qzd1gI8xOplvuq0Oo1+vGusjPQX+sG/FZY5k+sqEumwpAdiv46UjmNvED7Zab9iA
TTD8pQQcLAQF5cSlzsX6gKO0Ffdrx0OHE6GA2NqMDruA63aZhzxfN8M+N2g7bnBm
RfxFyfcmVqrgEblNBTzlHZ+zua+ckqIbPIVrUpWwE7m2jhf+0iOjJ8qUVnbaI4fg
GVIe7EaYa+E/84Lqnzw4Gb7+kHp6Qmdba9OqkRqC169RDQ1LsHAUmZ2KK9DvFNUK
rWgrwyu3OgI2wow0uWsKrPCWy/EO0Fjqo48+dT0tG136eh0tYj2an3gnlBt+oTgg
Y8ko3U9Hr9vjOWLr3wp/pvKe1zS0unE1VLsdicVfqcTx7YAK9Sb26x7EzjWoL278
VdWQ9/pVHsRC3OhN+EHzORA6Ebi8HGKfBoBylhKHMbIQYP2eQW7pKgAJja5TOToJ
A4BeTnbdubKH9CSEUPIaCfuUOoKe4KmJdpmar53xU0S9ePPuFHszIlztSoG95yWr
Y/tceDp5HAiTKpEyNfu/gKChDi2LghiEf3tQ8sX5wYj2bcp9w81F1qqsW3LmpaQb
hW3cQ0Du2QAVOsOJv2cwIE7ayxkILMvN0pOh99tOguPNfmm8pTlTmQh0vBPysOzl
oicaracBeQOW82L2V28jskSeNg5EjhsZkTgu8k2CZkAmoJ8bAUyglFDifmyaO/mG
yeCRkHdgNOUogRMEiTcsIgbHJPNHGXg+h6PUvULU3kpydivsjGmtwTDRifB6Kzjf
vEnweyrtkUl+w1IaCmaYsxbWrRcjelrMvaBN6ZCuLLelwX8iaPIGFU3HcX+VGz5v
93LU9xTXlKLniJbWoJVb0gn/RIOcpNRaTNnYObr1Ur9U82ZsCJBKDwTdMpQ0iHRa
1pPt/OdVFJPpmM59Tj08uQSnBBgRYU5OTAHRmOounars3erJtSUP4DpahTgOTP+I
Wp+adr1iEdeUVlYbqPQnjt61ga+uMSDwaTOUNGDt/N9Xf7k3Q9hOff9NyJZ0r777
tnz58rEUuank16GNQHoWL6d51I+wVL+aLW9DK08Nz8nExlUOTC1WaH7fj1DGNAyu
eJu5oOhajigDKxnm2mkZaxrOcMXPagfnBc1cZ82b43xwaYKo8yLzOFm8aKBX8d9u
FvztuSck72xtDdRhtwQmXTBbQGTroTlZbPnBmGLhYs8nUehfGjfYTFm5PGeBMkM2
sB9CGZc3IfVDrzY46nAXzjBYLnGnDX80AxcP4feBHM0UxwrSWWUEKwZRLL0D/0zK
QKmUD7B5NfazCmwHq7yeTRzHD7R08dtqL+ZwC/3pElAZnoVKQDP9YY1QlNHOUHkF
wLU2mp6txKwcuLX6L1DD/by93yALcR6ano3errB8gtOKZ9kXuv3cX3hQlf2H6RQF
8PIW//Uh8pYdT35KHDZmpEGSBt9uz5/4pjdfBKe0p1qBY0onbMl+PXU4tNv85mAR
k6NesoSYF9+o0JvYOrIheLr2o/yhB7Vr8GrJxVlnklun1+nhHBKVex9wBo4Bfnw1
laz+R92qAWFUDvpT7qKbWLXRVOketgcXXFi6a/Fmef6sR0r3lyE6uWSkyJU4UNi0
VjiIPANMwyuVNWQxCR6UNzZGpUYM/Ctok3HRKLgeLNlpZV4fKOEodtYkRwMKF0D+
YNSlia6tSJAL4eHt6cgYO1Ykqm9aHchrXOq/4gZzFSa1WuIUyRnUGtq0LgmpSaVO
GVJFRTEAwaXjzVwNfeyWmSZOSAgX2B/OIJBSELTKv3k0BUCwUqJDUuRyc56NVBdN
SQoz+brDxcYe4/l7ZpO7YdV9QpQJNonFear6XURCwAP2zENMIajhKQsvxn7bkHnt
oELOj+1YxbQJVgYd0c3xtnlvmu8Ms2kb9rgmUS/HOqqDKUcsAoIgrxDseC70wtbl
bSa7gw0sKG49OXfP/+HJELdgToQsmxO3QSl/nJ3Og7JyjSooFgeZCgNuhWTMotIz
l9+b0yViS1oFU9XOXHAbeUx8ESdIEGIMxNTmYfIGJ4+XWPb0iZlN0F1NRFFpkqD0
AdaTGnRZvN3DJLuJXelPaNfos3P2J0mrGkxRYfM6FE3FxBjJCTvaPWJYPxhLsQrC
/gJEb3TpL6fPrWYo1usYcevtkuOYbIFC2t1IqPsWL8wxlji7JARCqM/RzZ3+UIlJ
pcSCN2zR4R8m+YsLX+rvb2vJALV/+ZmBRP06rPGzfRM3Wp9lci1XhFEIQOfYSK46
PcPMjlw3uTsNatp6L68bwgixkVLdZAvKyzoP7xybetFJVv60212Ncwsfo0A7SpAd
m4hRlzNVxxu0CnnrQh0b19m8ID77XNNNpT/aLpI0w2T/Woc88dsas2K/HJWEYF4S
ub3pYe5jw07w0/2spwu6ohnefOcwnELdU0DCCxRgXhbkGUcTwXtIxdUWW73ajsK9
Yr4REDVvE3SDUyKEOy7NzlInJdnViMsD+fMx/2umFbwrCAqAg7uxA4DqZ+c5QcOu
rlhrjbeqsNCjm8f412Buwsap7moF1gcD5T+kR/H4O9srEYas3DfRSVReZ7LdTKmG
2R3iL5ed9yTAc/blH6VgLUwdrs5fBZzgOaqB6mqT56tawrHSyiUj863uqgzWF+En
uzcVnAtaTYab5m4GYW8WBhN64gbPQb1QFOTB7IaqkbYC7cz2kHha3Gkb+SDm/1kW
2QGEmtaj33zd885AnEXGGMxKZne4fXclHeIRdDXTVV53utP2x10SNboWVlocEYv2
8ULDGgOGLZzi90kXzMpqEQxz6JqxPRxX0dP5tEX5t+jWS/wEZTJF/kEHATA4waR7
ov49XhfZ+hNY28lW2hNrdJyDs4pJEsW8ZhLTr9B1ijAxt4+JvG7K6KVvHDYLMS//
8Q9UMQNsUsA1367QjWdFpj4ZM4qAPGDC57mhP6XUqbgkUoGK15p76BKgDtPXsIy7
HIQs9IFSjwf0sf0k0uXyi6oyLfGovW7BUnTYJuQK/e9tingA8J/XxfDXgz7B/Lx9
kTAszUkhzqQcd5g2wFQ61WZE4MK91DLT68u1+selMuTPbg/Qk7exJr1dGPFGydrH
vnhowW+nF910kr5OSe6CNxuB7xP0zBqYNh26MXODVzj5dp8w1Lh5VvhEla9Gh+Xt
MshRdQRsEskZu2Xnd6Q6ggCvniU6o5WPcMnu1uiJyCcS7LDzR+HaqwfWKrgFJR6c
92g+FsDnOAkzZSkSWoPsbSs52n7f8Eoq8sbGf3ZYEqkso/jaSe6cMHEkPVchTdOp
sP8mKyZk/FPlF55kBqToq6OD83ITHjhY+1APfIDr3Up1Lc4O62uRMyL6YR2/waI8
V5nq6/xXtmMR8phTnlU9xlZ9nKRmABVIi713vf6bTm9ND62XQwX4qy7EwVU32zoV
o/855lDPQLHuG2j+7Vi2ZrB2Z/lk9Jb10aidXhPA4Msbn2VaxD9hsU9OML6IxFtD
qV3o3pE6WomOQPENvUTPMd/mv1o9BnDTONL2/XxlnFpZBL3KDFrgk7511bsq09Rw
A3WUgfgBAnRE9ZgXRkUdx8AX7ix9ynC526mQdk0qalZs0T9R6rhpCYItIYUC5RWO
qbojYu1uMPx4eyDkQyOkTS1UItUJJcaaHn6GFBcez1wTiOSvcCB5OM/ck7jemwwX
qMdUJG6BkkDAfM37L7jIVvU2Gn4VslmbuK1PnPECbIgRjwzT67hdDxiISF8icNx+
7PcRXTE096MZhx9mfsuQLn+D7zSKhI6yuhqIQ9x76pt71bRvCe9eoGLcFZjhrimF
ahGlsQ+yXToIAkBpb7h1EMX4T/0zTT41ueLsRj/h6jvdlFh/NQiPyYruzP8lZtyc
S2SS2bhmc9muChbNlevGCgVzXAoIjsiZdbnvN3wiZCk30bCjlqhGAdzaoTsRnfcF
TXSHRlyuSoFrI8Cq/ErHtOA3eGr395US84o2cxZWB8Rqhn2bondJzhQpmfLqpLRk
tr8z1g3OddxKKoAk94sK5WF6scsOqUhKwCF2GlEv4cM7n1Jjz8ySj8QGc2ihCw2l
XQP/vtrznQa8UD1btKmzeQ3iMO7sGsiPwNmKAUTmpZXXN6oOZGQpfvlHVKTuOsl9
znrnmXGAo8Tdre5fWmpjEKj8uFFtaT0n9Haa74Jl+MNR9DzjWXIYM1Lgqqi9FxEM
ApZZtiB2CTg1a/DCV/W2qtaxZZJT3Z9BCyzFTbnBQukiJt8yeDb+77iBNzl2Dxck
OSJEFswPU238ZvqEKbnZ8Luw+ILA1wnQ1itYiF7yphS2+t+K/UM90h8uSqcUXWWe
aMWNviTgbOoHXYm5qvsy9G+NL2oY8aJGXj/Dd5TxB0lzKbDCDk+OFjvbkHfaljiJ
47e+BopBk30lIajCGkD+iqqEQuip9JFIhyCwEumzUyzhko/kIldbeU1qCwGVXdsC
yUocwfuIFviGs6arYCKUwn2skcEKHxj9hGaWD8++ydH7eI2IDRlzoFAKVw9FKeTp
5Yvo2UXU0OLRUdyw2EF+leJVJDqskOaNk9jOK/ABUfeqvojFTgjcPTi/IuMqm2gO
mul//bZcg8QuqlQpyp5HlOhd6YW8no8lbXss9oO7lQlEITBZZ0l6schhf6ybq0os
iQV3enrqmV6f0xzxmtGOpqkM5V3I3FScAYOUfWXCqYBzIiYGBrbd8W6VKBSukqsy
nDXFSXeKFZujKwmu3zLw1XKtWn02BIrFfR9RY+Yg6ts0ON0c8MzPku45ppd65tx6
1NBWAnZ50E8mY9IrNiY23IwF33jlaO5BAyXTZs3atUIR80qu445wKuQapxTpNBj8
FI+9qkky8nRCpDN2mYw3LnoOv79uoAWWXM3INRIU/63IhYiomqtW6n33/5io9aqx
bCEbknG4QMLfCxOkkO+5BT4PK9KVW5fObrtx7X3FqgS7Fj94Q2qpwTj2WmEhhxQc
YkTcUeBxCHrJTMlacTVddcVhrbJtsEaCV/qhHqZCgkfk2liYD8TL610Q13iiMNI9
9jtotlB8tUUMGOXq7dnNrroZL63YtlDB/QMYX8FIsFFL1cRJu0KH8G4ZXoxO0+Cr
YyCRktzXkXHR6HiyMt4/i4UHxeD307fAzr6w/rjqmr2V3jY6s3OcQIRy+GV9DyrS
6oVN0jGmckUrBQSecQ0iR4Ul8eIgH4S59xqS12wsGRVwiA9MhUbGj2HWXy3EBeLh
dj0vS/90/5y2YkNoFajueV4OcRGfENbUpa5ALvxafFyWmO5tVEXph4nv+rLguWw6
CekixhRzUYYddG0M3rLJCPbbo1Tj5HQGeh2ykr1KxvW1EAtwweRNFoFgic6QxcbL
TBOcrxy0wG6zk/XlbzaZo/cSY2TiyWx8dBjciy3vzs3HkOmO4Be6pWyDND2eyyYm
NEW68ltHzxWc88x1TpV1FxrkmScCvTWg/TQDe6DtHjfeLkeYOnbygNmn2nmqsbWK
twCQQDtqvkSAxvIgAWj4looCZFIoTqeH/GUL42TRDwCX59xdVwYvUQkE/BSXrLKd
NTvxqH2aZj0InTtKXOmm1jNK5Pp/g/0B53qQ07S1Jhe25ZgpWaArwd4U1l4E8A1o
mXMtnqoKvIdLaGkiZodvJ8GgZVhY6QezYq6P1qGtNWUHPomFKkShpXDClsJLi4Do
rusfC59u7FvPK7M+8AprBn3QWFm/tmmJ8nSsIvvxxwNeI0CcBdZNDVWzwzjAAJ7B
FyDTKLdTLeApV0xQoptaIMKM8kfjLTWoSnaTAVk8Ysv9e1aSJ6oW3plh6kaw26vv
GhY9OdJHefkQH+KgUXHWqk4CrIuornLBAvUZ5NEeWlN5uprvNgft4e4IKPcOZzsU
y2Of8UUxvhkDUIoIEmTshoaOlOKW48zvc1MHn8BJvSpWHfpuJKJhD3iNq5Rdp5ot
fQjgKKiJo87SLXzSHf2Ag9MxxW36powKv21XUDHlUXrgjqZ56iml4aufAB9H0tQZ
B9Mv2IaiIrtoiLOxOu0GhtDVOMaidnfgKp0pNOuvGmyHwnb+YPaypIcNPI7/a6wo
uwwP5ilrSwd+qo82V1ffOyLstwKdlT9PpGX2TEsuOT400vlO4W89+JEwpdMUvm3f
0+idFJCswWdj2LIDawVN3taqC3aOOzbh4ifdubI6K69FhUGRYjVUnJtyIbbZBvuC
dNC37SBumHSKjQUn5fNiwdJT3xLQDrdpib3utu8mi/MJ02Pppgi1/6AKP95pMPsm
AtSeuJ5wwkXi4Z6U4SG8q6YvrHJ/y7ZrAi5NWeUHHfa7v8ubXA+vgKwkbZMLS518
ckoh28dyD9+IOjkYeX7t6Q72/7DgdCMdBOaWSmXrxhsuqFzhVXEbM2TDqxJSKgvM
jClD0+97Q0mGXUPvsfyB5iMvBbrQ2AVW6fq8YpCoIjHU0UY0dF+i7bn1hEsa9htw
H51xMqnC6hL/9mZ478A9zAkh5Ufh/bAyJ62g8BATYr4bFVLN6zRmcA3Msrs/kAfU
uGHg7cD6BMfJitrTLNsWCecVG8sY+q9M0iekcl+HZI0Q5UFWmlgNWa7JybHRDw4R
bnDxchVeIHgInxnHvIFl7c9fQcAGGbDFyLknBc023+orO4JC7I4qcOHo5Yly02ok
nRfbaZfVMkxScdiEX4V9JxW5lmxuGcKLpYVBp4q7Yb4Wio5yp+vl9UZwuOpsB5MU
dZPVZ3EM0cvYVtWeLKrjlXzYLF3GraMyg38cEPfZSbb9BVK1tGLBka/nXcGj+wdK
JcG1k6UlZOWmGB/l/xAG3L2qSgvb8RTFx2DyR25nRlARJc2SwIovZeiNX2nq7Rio
LeUwDQ4+1FweTKYkKxCYTkxJeRWQKpLsn+cyWuyp2x1dPBIHU0Gqk8Hg84jfNhKf
QuN5wG2PM4cBnG+p9ln7Dl1AkmVGV0InCcQmI40p6supjvVB+/oCOqng2kTeMAE3
bt+cmvgDA0ThKTJ6UPzV4GAJoX21byNylpZ59gd5UdV9WINWeBMJqijb8nIGuZSY
A9maskSWxKObXk+F1c/bImrfoCBCmqZAdBBx5a22v0Qo2BR5o5xDA8nInv4TuEgO
Ek8V0vN0fjqc0Fm0s9OEgB6U3OPvUb7Su5HbklDcQr0N5/XRaSnwCNOYyoDLvaPP
ILxBXi/p5TKNXQny+6cAnVlnbLT6awuusfkxRsvb9TXboZ0hYtuT9ZShWAej3e5s
UqxaPS9t9wUprZo93y2OMcqgh/zsHf4lUGP7mFbCcA5T2Bnl1FsFY/Oe5DN62LPh
L6uSpl759Z/QqnAo6ti0O1p+MyZn3daHHj2rbq+GCBN0mxFNOAV4eUWZdGx0KPLv
TLNzdtrUsnFT21lEQPCg5+mgZVHFefhLEGcBiKMnFlP3fW1clU0JfEd7Qnu5DvI5
87LZH9cOvIcCUB4DckgyraOlLXCRndQrQ8aGvzhLdPP+pL/L1qwRm5RkN20be2TK
YVKCCtx85zmDkFi+8WSUZYk5t2fUS+2KQlRIz7JYaRso//0KO7ECIqOehVHU2dZp
lNNYRYYkYe0G4BIpsuERysf5R+QCUuoGuvAZXA1QGIm95eJocq7tCj+awk3NooUm
gIeW/YCMc0cPk9DOQZ+YtxS9KalpqUu/fS0SvxDj1mASkaBE/OKefwHuCtHUdweS
j49gYpOjDT5PyUmzKJ6jCLgG6WrzqvESlQjXFb9P3dg+wdAEDRRY8k+lg9Ebc1xQ
toKxLbyiLFH/AWlxDSO/+50Ws066IkFBVNvB5YkNB34US7sZRVMLwj4SeXRZENnS
5ltICjgcWZg7q5T8wIgIkJXbVWpobTTOPTIv7pgC724XPgOsq08uMqdkJVmWL+Mg
lPeGZ1JDqEe0EJJeLrjqB6JYjfq0BqdmCakd51hT3y8OWjfP6DIKPd88HudRMd7U
JUKpqAdykaMjBs/zhZn++efVS4zmWsnXaKzYb5qgVd3pnhm2EOtKjUonbohKVrbb
k5rY4MXz9DlCj6OA143SqGVP1tcVUFIuZnqDFV1yS1gDDF22GTxBL06iio0UbNIT
mpXSeP7wMOqB9MT/4PqQW2Nf0MqOITLUdM2xjrRf/P8Q/hG8F/JiCf333ZnX4HfA
8EFkxU0dJa/2HqUxifa4McQNwb0UHTPPDzQyfXAi2cDT0S9GJgkds3MpS2bhkRjl
bgdJHLvGfR/cJkocUP9Pk2ro6rrDSMNVVhx5MoP4ofXsoLdyQW0w76LCN2+E/ceT
DTPD+e4yvbYQg08VpsahG2Rq5zyDzsUcFvyWLUKoxbc6+6y/6Xz2bktZFKi3snT3
Hk1VHXO77mQZGi8WrpLpxrzxh3OnAYpWYDClIm+eYA9FFjgsllI+VvFvNLxdvgbE
15o+3mZZTufQWKRf/CW6Am7Zt66uGFwFvcUVfhpQ7fFWtzz8bz1ybIlRbNf2wWXl
ZANZ5MkWaxgu1ceG03NW1qiwwwhRoGHUuHXlhAU2FepzX/Sk4zhca1iLdJQ0D5aF
dB70opWFXWtjI2ZyWTMDE54w/i077gg3k/yT4ZDnjv7hk/a54NW9aWwsWBYQtrEY
w1qNZhyFGI58ELKa37dwDqExE9kPeilGMkmy7PKxInrDPj0ZskUn09kPLo1kYsnV
HVHHw/2kc3OWXdD6EphGyPZwn1VtqjAHBqIB7QkgpFx9leqF2j16vds3QNSl1bgT
VfHJDDXw2Nzf8NaKdqAYPO8OlFVr9y9ac3bDlGscozhr8VVnPy1w1UPKWHiNxFN/
JABBZ1UThuwcrrQSGhaduStojVfTHCjwpPpaoeODZgCJivlafIJ8IY8b2sYSQvct
DM7yA6WuxoZd54nkfJ/8FuAjSffwyDOiH3PejukjDSy9UWuCtAjjnOiP5pddbxjC
PaTYSUys1DCMofEPB6vMWrDUpqIWInZlwSprriFWYMS8K7ma5CcG/UZCOvZKeN1O
A0gBwQGJiLOHzGETFBfVsN+7YXmWtZb0TKaX/Vdd2vK/v5m3Ih62kfxDZHpUGan+
SrMs3GBV+T1Woqos4NRq9CibdX7uwp31Tdfoy7gIcVC0rvZdGUZSgEXBRX4MO+Lh
qSTNMYcHbRU9kugTNl2OLfi2jsMp9Yydq/9bkqBDfc5snv2hDBPJPHYGOBxXmed2
5sQxuXW8Rt4ptJuTZd+zDAnTTOvt1e6AfmrGPRq2HwvVBjueFACENZ9JClwg2Lqf
R7NP7R3k+UAuq1wIcYaEzj+QjeuJdkLuMAEQXTVYz8gtxc+wT1H/8MmPVDi4V8LI
YOzfnk9yJzVdBSU3OEnqpE2w/8Ex0cVAFWMtieSrNp/yi1iI702P/wpEPkoq7XRp
S0mXLxCUse92/4XNUSNb+n89wLUys6mNMvWRArHXXLJ4JqGRf+xJxK4GJ+Fbuq84
viSoflWdTFSe6yrnF4bTkVH2M9C4U784pJ0PUoeNK4Oz3naTHCx3ShNbH73DfQNV
ZqFmSPtW786dcRjr7LKnMc/w9qNsSzsSG+Pd2+TzlWdbIWquMmVW2emR1SkvQ+OO
2VxZzJgGmTIqOe2ypTNz/bK2/edSnTlMidM4Qhkbr9+noighAhqpBpCeB2pHuk8U
MSPy3VLX0uNxvCIFPRvGuDFnvP8fwgyrHokJcd3eEer2izGRqEywuGgGXOjaH60t
e5hjYZESis5RKkELyXov/SgYVCj9hsJzNIF50Yb23pjmHxp4EQgO8mT1ZO7WKPIF
SUC/GoSRh8xxnplUwb5UNjQJAvSvuY31L7RYw0az3OYGjSqEsFCpp6vptv4yGiNZ
iO0eMWuERuQWHAfx+8F4D1WdedCnxVaLQ0Tgovzxr2CZI5iDiEtvoqLASpANHU8A
jlJcUm6zUFj1Kr6ONOGtJXZYeeasv4kMeR4GboReq82rhVGMOpQeGeAyC4AFlNFV
wWX5Qsd3JhRzpzaYwLGwAffwQc3lrdTh7IK2ti6gQWOcAbqTMM+cHL/422Cg1iyK
74vN+lS4AVMInkqEw67hzcbaAEPlLkA8e26QBA/0vyumSewnOuGkZv5SJZ5NjlTv
LlTmHO0bVLBQZywmLhxEaYtufNHRgNVEZaxI92VeoSGaGjwAtSjcX426QMWWAO8s
e89Ocpooc0gWVQKRYrZ5ijWzo2K15czJfkaiLQrvWscabRXKH/w//4SoamDUNfTS
Lk9+Hn9VH22g59hdNSoHy7hMeIJRQ35Y/fegt7OROi+tHUzZ71ZTxkvA3c8FaX6n
INKQrRtQPSll85CMk0QayDz26MhIWsoW0Fhigho3nbtMxPowoV0iO6mLXHTqDoh3
up0wEvpbEdhFAImKU25XvzQ21I0Nmk96pkFfxAubfuuTwUqiTkoRTYEdu+GzpU6L
23DgCHNCt8Jd/iW4abTYOClH8YU7Yt0PmEQaTRue3e9y/QXu6uUlato1uL08sz12
N4V7+CebqD78iSHXTcr3qdfdVnJTbGiSSnE4CJaVAImBbca/i9ZsjUc4jXIdEo1g
qCDtaXXhOGjtdhgNZ363ww1QyVj6cQUm9NTI2uDMJ68Q8EDPOuhvOQC/TQynLAkb
b0H60gijYHYRE4HzOcAC6BVPYtYl/cpjihw8g/MsWGxOpwLGwZUrQnJ1JvFxM3cY
KAIR+PYnL6LylyTesVubdz8wkZfG9qR9ovxFYB/k9b7c2A5hCIoYl/jeW9qU+tUd
uMFGdluAMxo38oMMO6mpD3kC/CizN/tw//sA34kHJXvddhmiuHW4eP4xyw3eH17N
g7YgN6KmPcvEcNxOEVzfbyQ/Rd9MC9RbgUkR1AcQYbRurdDR27yCv3y6uwLeqZ1f
aAm2FK6ALisPM2BsMMbGpxEfYC8qNIipdJJtoXnKlW83Vsaf2G4Y2K4KdfksZ1dt
xkBnlpzwTD3kF8wDOxGK//crlDsbxab61eAMYcEDdPGJfKmxR4OrDHIhI6F2vQoY
4tNkYqD8Lpxa/HBU86jL9Eu7ukVZZKrV7urbJNyaMhjqkHS0Zx2+V3sym0sHfbZ0
t7+j7AF82DvWsjqmzx0Z8Ti3LN+5E6Fd7PlYW3hw1pSDg0kaBtcoiwouIUkvkQFp
RuPHDOVwIuVKTk2axnJ6RwXEwJDnKYiCTNSSFfLPMJTkPt7vZNnemK1Emy6wPctB
AxfK0IAgi1Qi7vrlHC6MR0oFc13TwY+BBKClFOrPGCLCCtljVT3zsA53e/oBX3AF
e93G66rl2MRVFEedMY8267N+lvGkzLIS8+NID71URYJO9rpsOK8Naf/hVC3rT1P9
zqluXuUirA1oeAsC782KMCSNwu/xLjTenPLhPC0TuXvJsc6NvIXSgbhH/6Pf6iOs
YjgP8RDrAjVAeUnYBmqdnI3OtZ8xhxWA4HJkEHWC6ZNgK448ZZoALMsjdo080KcI
Q3mySpKoS6WoCvH20xINNa6IN/swczMFrTGdW04P33agDg4JNdvvYGIG0SQvdZCr
cME6Aag2Vdy2tKQ+fqnrLIQTCGz3etmKBsQpCZixCDW627xVNKdNoxi2QyhpQ+2K
9g1C0CaloyW9NHJ+dYFzA4pT42MZbkXE1s0UZe1Blqpcjn8TXphZzZfoN4oLNLyd
faGR+QmaC6AfLi1QSwcTjS+7N2RZ26rs3cGwT4BzFqNlec4dip9qI3l67XFKGuD3
xAG7jiI6Ecy1dfUj/Pwlm91fF96nsrhdNKV0v5gF+Hk+1y1xTlKuYL1i1J9YNJYv
VY6fyjmZVi54yYeQpqDHHygj1cc9s0m57HLAytavPzUyFNegXwUYd+XDW/tDTeUW
v6hXSm50j+SKHIGtqxHJqYey9un0gx6X8+Hhoqx6nJ1K/mgDFWiSkKnBLwdiq078
ZmhrNtJND+IKnG6ZW9OCntW5YN1PGyaHVBmxvYV3pC13LxgeyLh8H4dpkY50vEOH
QOSUhFZBvup+3TNdpBOsM8yz2pjwqTkq1eaPIbBMjfwtjHUAImLxdmAOirYzkP0D
K1lvDNlm1pyQSSsj9tJFY6h89NrSnwIvPibXEzABKaapj8VuLd/WL4OIpqBLbZLV
KfwDaurPXpdFFlh+l5NOd2RYfHPwLdvxnueVkZNdiFEYtmgmfeOjm9RuUoAKQq5X
/AwGW68fnVd7/K2bvuRjIy7+SuXNQpfJlxQvSfZI7/nDPTQtTYWTY3XbnTR7yai9
zXvHNOm1U1cX8oVdYxlUpTHgU4AccMWMmIubSKK7zQyK7hAKnUlcrcnFQGPIpu94
37w353Avif3D7nQP6UvjyBYDPgJGO3scMTYhbaOLBy0EQUq/OW+Qb3WjQ7fQGRX7
2P+hyQtGPLDd6vuv8jUATKlrq/rjqbv239Nt4uL32ivRJIdkFDky3qSZkPQATOVJ
ffd9s7Pv6PEo5mDO7X9Iohm85vmRG6EmVSdl32alOPBtgZga3fFRdpVsT7M9qWGo
AE9P0jM/NkQ7idL+dHTRsQSj8zY1G5jEwWk23vWP5eQIOU5csP4dWoUk92s4sWpp
abycqZVC2lO4SSCb0YyUYBdyPCQAKvnQ3cBcnf8Bg8QpPVZ4bx40c4AXLf6Wy0Zk
am6xCOX4BeMMN/E1ghjrN4GbdOILmGfpValgJBgeBAbc4SkC4ccrPbQhWiofCppe
65kD4uWlWd6Zm/DIt10DO8KytR0BDFyhAmURVZWPzokSIMmZKOn1nnW0rk8qyVnj
1ihYvIiiudS5dm3E/XV2P9YohnbTUNVTLJrtQ2A1rRt3vGA0zdw5EyyUJJRv/mqY
qzKs7aDWZjaY24v1Gc4oo64Dp1hFhi8LgvBv37WQDiZRWrQgEyNYW9DIfs9+mZbz
1wdVOr9uIC9wdrsoZKArBNDduZMG4AIqB+oPDxMW4pEoR3v02XpGFMA3iHWHyqV6
zKfwXgvg3thDQV9tQ8sB98WEwSOTcEoC4eot4d9tpd2SP76BdAjyBuQ9goywzZxi
rnjuV+3KbVm/D6qFPZ+XiVWM5HxXQwcj3ILOu+K/srXwYg8SKyrT04B39Gj+cP5m
doCTECk16es+eLjN7SSc5s5+9Ic3Yn5tjyUMYaUJpef+E+v1KoGiNGxbITW7ZNJ/
OrSKdi5dgptLwu7ld+lcWtehrZHk88kfh+gArdk0DaWveVrT/k5zBYs6TEvcd7fI
6zejtiMSfhZ8ZZ24GZnnb/h/0GDN8Fh0TjOHQChdnjQqyQKlpF3VoDpfRncvWQOR
zZtD+aSyYPY3Vhv9O8tcmMpt4P5XeI19BijT1QxjV1NGP/IaJOr1Kxtnhl84cx53
S3Og6gEqz0bTGWtjm2k31ak/epOmlADT4vfV0HawUD/GxSe5CfBYDDC5T8piPC3C
2d/WtJYDCTLxwUYGSJKub74IXwb+UO5bnlLFxDK8NQdHY7TjXcjzTJ6BVC8yewnO
wxADPQgcYsfi5AvU4NSkQa+Xt3m4KUbvh/jbWRBWcivTJmVAK2hrnAbu1W0Ab0G7
NbLXGFRIuDu16PFJIDU2xjsJKh6y2gw+TXyzrsDiFHCYkB8xt3kO7mEX8MUfN7k4
qIUtBMcZJMc08PJepYsJx52WUPk6TV+Z+eVqTbdGCHZsf+hl+P+Q253JPgE8uUP7
DIi8LqC+CYleqGLHpBnc/oxXJld3ewlpde8mU6A3/pcd2zn64CHBUpPCFAQiHMZM
uQTYslMvaMhdTNJkHRjptNBBu2JiRzVNiX/etLF2/YtYTtzMWns+U7iYKFWhH236
ZBplBW0zPQnu8hWz0hDqdx41KR7hiYNkObJ3iHFFIQoS/QJKvumZaTOdFyjRDlpm
ASF7AkCVIq0rGtHOinAdzhDOQdQqhEWIZ5C/cPan7l5J6XTi+odoASr3O/hFlELF
7RFNKXwKreXIk/b40kst2X/5/12rpQRe/qvIg0WXUIB3Pv65BNg16aSH+ajEUGqN
Dd5AdaHU5Tdwp9w/gTBHwBqHwlUL9BpsLXzFwpDr8/hNAbNDOf9zU+27d7GAEd/q
eBrab9f6NIAGApLIueQaV/3bV0eW1lRB4oFWT2+UqSAVKDcebJfP/KIMxoQChbc6
kSY3AgraRcWqme4Mb55LGoRo9mqniyK1i/+sAM4jvFbzsGuU6h86r8e7im5hXO+D
cZhhgnu0NR8LAOh95HB8CCStRK0evj2voEHXvKhhUK8uN4dNi4c679j25z9KUohc
OBYfsjBPUqfaWL5MGCbonQN639neb1QvBCGk+x4jnmMbQZJqAhbYb7arOIBCkV5A
dQqAm/OHNIA2+DMUL4hAnq41u3iv22fBmtr+puIWoHiXUPWVYyzj/aHyZAzZfWVa
bvhnINOQITVxnsksxvMyOzaeQTRT6rcNfjCtUUlb+MeOlPrmeie5NVT3E+YLbtA6
+D4+qaHlRawG+ClFozwextBq5hnys5bjyPkz1ihSvd71/fn0ynmRcYBajsYF9HFl
gD6N0SalxnHB3smJ3PiCE+4ILyq9ho49RRO8c0qu5XXCus3YLJGHDzmcCrc/O04f
hV+x5MtTHTEaiF1PlWtc4A2NPZlMyH+mSALybAI1SWsLQvkjz0g7wRCAehWa/8Ig
f1uHLiuvOYUgWMsBJfoZ+146pK9DfBRhiO3T9aI8QynM1Wccnok4lLuH5r1Hs2FM
Y1hB7gpKCVc6IAS/Y2SMi3p56QFnJFUnNsEhMgP7romLtp6wliIGK6rNQ+lVg6/c
TYJSgf4Zny5+MQtGf2QcRWMBcm1LhK7IBdl81CATh2GiqIHNIpmV2MqyAzhCrZci
340y2lVM+LmPe7rAveaLIyPFlI0+N9aWlr1miB0YgXDmVF7sk7wqA/lh1IMcoNdH
8rTMLLbB4lO4RkzJ9lyfKQeo3Nv3WWclwwvELjejZHFjBFnnXrDv3rqEQutaRVML
mle+reEY5xu0VyE42ayUZBBTtjRpDqzb5rmKMPpyyKzyZrKexXqAaPHotXMYD02i
oNCQBJPIP2EKbrpvq7CX5PCUR6aSQFIq5/ZqiM3201O+lVystCjwAvPkey7LRGJN
2h2IcNCQjawWlWcc8HjZuzZxa5BCgiXS0iVgthRoC0XgAHTPs/dom0gQiI/FrrO4
AcCW+2yHIRVALC/CuSeQ0gWcJCqQ3Ev2b3HCxNKtUGb4XG+qPPK+py/pWk90ZlC1
oX/jw+NHHuejBKNWXCh2+ZS7KQaSbJ9EtfKl3JZSGxTbY/4TJ9QXw0ZPijRVohu4
jj6/PnWcdl7vYFPePa/nRs4Rv5BzucQgohcyiF639TTP5dklcJA/rhCS25PW8lXz
myAoKNUL1uiN4saOkGd2za4og4Z1UO8lA+Htgywx00Xof7yDn5jq2RRWWSOJmAID
2LOI1W6901rbq2fB8KUu8Ni5qfDgqIM7EhDppM3whAOsRHH385uo8JnDfp167VFW
WgkCGVo0thivsUMZXSJUu2Kg1XNaIJE3yRJQ9nsTkEDhT73fnDgBmSlV1sqF/Cpx
+FlAUuCcm2enOvm44+KIdZZi6MUzM4YKnRnnamsrstIWKruFQwrH0U+Ym9lwgGqv
PGR2KEilRlkY29sXIGb60P71AwwmDO0z0Fte4/1E0Wnms1F2wZ4DTIg1YPZBwiqQ
aWbyoodh68P0yN+Y75pBv4skuaD7HAgwHZJiM+OqqupcyIRF5c0Onb6kgv8tfOKN
1Pm8TC5NoqaeiM+12JJHBwrw7FjNRJnLdb+pGFl8LxR+4Vl1BhPlZdwVuqEb219o
LFtNEZRLEqYAEF5lvZESg+TFI2VT9eAqePV4HNO3cgzOhDiao37id4KJ1dlCDnBi
73drrzkg9H3j0QK28a/iWnDgTE7QdRcYYyp/R5XlId5eSRCGc2oQe/pchMwHQw2a
7DfhoOFdnwJOC188PF35DiY9RKeSwmNjxWNzSe2uLZe6dL7ybFwMpeea05HWPa+3
T7iyVKsGX2e3yuUU3fvrbly1u+w9KukhIa39YYC/wvGCOurxtvvQoFAYAGJWODjD
DsTYYRhKOBkcQAbZL88z67wkGvQ+0HSHW/k/CaN6mHkhBkLr5yjQqycKmCKoqUW5
bCvT0OT1MAiZ98+CDqqeXM1QqZdm4bHU819WF2KzUtY3r9EFM+IL+nzJrz287wcH
KNYwooBZ4BZDlXLFaNDJ6NsSZwN/zOnjEdjwqFB9/RCtslE+oXEq/Ful/3DjURXB
ksujKoLOAQX1Oq5CD7SMXSEhd3o7YXJFWxwm6ZmpztaAms/fGpeOd/3X0wsGlge8
trS3bK0HqJ7eHVUkRsTVQzgJ3ZKUCJhr/iXVy5F0hAtsRV+nDkPUK1+/rNhG6NpB
Zn+jieU5nRqy/g6nMiz8Vdfp1Pu+u7kJuLse00vL1FFDMZ8IovYjAOpD8wMFvbZw
Kw6I35AbLb1qSnjW65auOfsGisP7V+LgkvsSkxbaiwpqNY7Z7rYTFo9UOXgn9Z1x
F/tRgMH4vBUls0yzHdZBMtt680qz58bY6ZbSQsnP6mf8Jl5+FNyBx6UmT4SyiGp6
lEES9lCffHE/sHuXxlbIL2k6HVjEBwClTYyqlJ23bqGpSth37ttRk8XgLUWyynS8
7ZuWa9Ejv8bL9kUMJPzXGJ6uxubwFzgBx9n8kK3b1PbmZg1DJZgMutwhULQ4YPre
GW7Tt2zqFKKciuhOQSLrE/8iCKMxsS7JgHWK6cya8uPS2IjxGkCZIe/vIGOri6ly
nwPL1wDg8Opvu0ZD41baMh0VLHkelRkrFwt5Am9mWPKrK9x8SgiWXPy5XlStX8cv
t5Ykw9BfySDDfdI5rSIYZKSJm02XqA33M1l8w5skejP8v1f8zUIxFCng4BmL2KNb
+PZMSUuogkkpPI0oLJ3muVe6GvEwEhirPa7rWwghPcaRkIyBFBhP9toser0LeuUb
0Apy2usXzvjfI+nq/yyjolhkobjD9Hl7ZtkHpvJblUKyo193irVi8ffCjJtCIgNn
KIqmj1aqkM6ZIaDj3FS+7QWnEpRRYmPK4U1FZjOpVtqErixFYpYe0D3WvLsl+1e3
EX3CkoKhzXS4rKtqTVWr9hT4KYykmMDqhtvQ2MgMli5EynGWsNYTrQrW7UBdMQ2L
8je50aut9KS0AGtzBw53sGA+PRFvMs3YYgtSOEGGqslgzPvVZhhT37fA6Bcsl3T4
n/ljLABzhrk9wOiTXb0p0mtBT9MwQbNuyhmxN0lb3zh2v6Od26e2rGK48k9aBxwg
AngRrLffPImWSB0GNejUkpF/sw2O1cMiJiyKPFEDalCeSbA6iOn5cv0QbCELT9b1
98XI2YLxlLUnnPa08MlSbclxePm4+j4kZmXq/Z8nQZPhXYOPYwZYG7gfWBRpR6bU
KhFsTzOhwVbUGsoQDvejBMdnElVnA84IzVDn8aJUEwIqaLza9kErbh5msGXQt3r0
lV/JvIPPmNoYZtz5bFto7jcb7OT+n6JVOCH6T4TyFi7DVxT4AnR/VvIbycMYxJUA
TYCLNMyZ4h08xPYdzTgrVx1KhDJj88xS3g2mYpGShT/4ZWmh8l02oFJhu29CfcW2
v8yCdtsFOKN4FHDfjHOYtTa5mOITL0CgoWBoUBLbEh9QHrwVvx5zWwjxNoVCyUCD
kSzny3uWPjZ47qZXdhWtvLhp0wCsu2DAYX/z/nkbfoQ7zx+//g+DdGZhtbT4VI5Y
LP41S62/c38A8TAX6QsKg2Gx5K11DyyryzDyuW7ExgNDTo9TGKPxNL1nwT6tjU8u
o5hU4tGppRtqDHcZINKOVGGBun3KblrxiX4BeLpgkrtKyLfa1F0HZTXghGO9tGxa
AV0PTqYwaA+vXV+/OeFQo5zA4/37Gg/SF31bhhiBRq2GLaoFnZ/Gua7+Nr7rnLir
dSjs/qh8o0CJKmmFeTN2V1GW8sVaPZZkARHMgNBChNhRU023YGF+bIZKmmQGbkqk
+jvfRR08PgxJBgf0fLE5D3F0UoZwR1UHuEjPMHSHvQRopUxzD5+DjwncXVkDyi/Z
/8VyqjMzjUeZgZ61+ExmBeM6+n+OrHrYEbH/XetQkCnhzO9YH3Ehdj40yHMdsy7T
O88TvYTjB6K2u9qZI8mu02m1rC3L76/iNyQmDkvwZB2dm8z7ZQfR+GPzSz3xhZg8
VdMDjTQCjrXrm7CoodsFlG5Noz5+JpFuYYWpKfTJx86r934IOji+v9FqL/FKJjgx
qV8MXbD6W/1dvIOmp7YExJzuJWx/D9nPZnpXdRynjfEcEf6iqPCyKs/xzFuX2K2V
WfwamUxSa8NB9xFrf/PJAhb553/io0TicxMmHXSQIpnZPKvaE56uEhOmUlYcEbii
21ZO3WQnP8dV7owRuE6kbx3N0DIF804jC3SK2qAfmnjyValKM3pL5q3iTcqBhCob
hKDytOQ8UyZ+ngjgvTTJuLsGj3BQhOKpBOH5N+aEpdHRLuflT9RxEtUcON2BiVA5
JIFYgSRIVSkeV36SHSwmgSoLd7l2AmgEldcThxki8o0Uxuh6AAIi/Aw7Ne9urzaR
lTJZY/00bFLfN88TpudBrBk181shzzG4NFlvQX75NPQo9DN5d55S02wpBIAS85hQ
JWLAC5PSICK/GOSHMnA/w/kPodClxKSC8xn3VthLhM/JXmCDYhR7nCcKV8aoItPq
mAiTLqg0J0na07RB3jgN/Ip0Vn5QhYkLi9IQOXab3fPQtuBKh8HulFK+3c6HuGBA
2dx78RDyQzNsKnBMn840Nwh+4CUG3/pbtrXFxl+I9Et0dzt3VMfjX/CPdE44UL++
i1M8qfIHnE9xwL9yfc72wl1TGyOWSi8tGy8FsxlNlpodizCAAA70qBhSoa6yHXDd
YTp7ZY2HyoBkWNIkZSR+HIe9SKvDh8qaX2yYdIJMZVVgQ+lbXxfYGivphdXvuu/U
tA2YdeDURh6PXoNtDgOnwNUqoQYi+EaBWGw81ZfyoWIT9qiD0/uZkM8RgUUCymod
Fxz6QogZna6S+OJHN0aq5gZKhgoj0grW9ILw23TOsPznuoU1t88aPmLItreUO0n5
NnRCzX+xsLEd5QW+UA+eh6xjWEHDHtovT4Jv0el861zF+DMS8J5lnaEq1Pd9LXg3
2e6Er5MdQ5P0jKv5gBBXgO7qFjf3IA2vit3m5OKR9H9kQZufwcIolPrxkZxlXYe9
Bz/SdfMmBbOZrDRcqAcI4IoTblYgn+AMhYBndIb6E1zcuvC8Dujek+NKXXr83P0y
fDlNT3+gSRWPQSLOfu+Jff2dwVKY6YegUluoLI2X41zAvuopVOrSNXfXuSrzTjcU
Oh24ChZMXGKX1GZ2wR+Jl41tadOYCNeUMPRfF3TbJsf+cC51OrsN1+bX6uGfU5Hv
ttIHzrziCUA6mdKBPaifXekFnATxK9AOLufMpNHjfFu5r1nacyJkYJN1OW+gUnG4
3TKM5gKplhUgCoa626U2KHVsZo5EMJTldyfDeI7oQvkQcKX72pDerjhryf69+dDw
H08fB0eQ7fCBPbCzQmnG2msbBURxVmPw1vwIAeO7QxV4zS9FPE04cLWIfafVdhID
XyQ7ckRkSL74cUreTftiMJplUW+feuDZ4vMiTVEtDP8JDOEeMUn1H4i9YeoMnVPy
Kkl84N+S9c5PYvulMxLY0OGTfdejX/hJ8cAcoDrinGmuxS3ADA9iVr3/HDGhmn6S
fwDiKUJQpZOjArN0TWLV1ZvBePCboO6YIfSl/6/ZYukUtNMkm5I+cUyRKoUfWX9E
+ClgFx2ONNh/xp7QaKNG5z6KoXVEtAEGdVFGXi86cOtZGD6jj6mWkKM6XN1ibI67
Z3IxMiX4ijL5XyAf2XFUUS29SG/ILxr+2qGdl7lQtoJiyjTMa6vP78JzicxyyDnr
UuYmYCm7C2WRQXxX+vvpUAqNst0VVMx/WpWfUta8XmlycXWyht5uyBb4BWZqHnkK
mJZtLTXCfpO99Bnre+kNyZjydpNTSThn7Z7YWzVoso6MtmOPtvwazqU9qlUk4D20
1JgsEpRTGRMc19p+63Q4RP6y2cV4U/6dZPY+cV/sgUB/v3+XdRFboBv8xNeRUnbT
GXLdznaQBS38dcKYOE+yCpFDkz4oH4+k/vzq6JsOv3OMlbX6wHy7U/eGVHC+Tu2m
hlqmeZXqtRNq39vsUSZHWHtUvfW6R1vMndklNI/LXtOaP6V5U3uKzVOaozEp8mxr
2RuVKkmiX2Pj/C8vTOSyHA94A52DcunirCzMRz7Nz+zWMW6gLKmXNK1VbSb1DVoa
c7mwyHWrYqV2IW2ILsZzxBooasVJ4Ygt3v/upd84iS+iFwPitEoy9s8wGT/es3s3
ytN4mlz8LB1ALw079UhJi0OZ6arLdze3b+jJVgrSwN8A/j8bZZr5vTNn+Gx3gOYX
YxECSTBeZIxOgUynGTuO/AvBiOJdOvYX0YeJ2TsfyGcl12cxLuvqFUk7xTpS1RIK
oxH9UXdTbKceTzZr8xf+0eWsk3Gi0flqtkueyH2F35Kjf9do9v51LR6nOBO4vD3a
6TKh45wJzIcPxTEfJtvCRt6Ou5ANZXcd3T5X68VpSgtOVj6hn7wOLWhzRNgCVC86
ukqZMKfDb718w5pInRswmedY5sQAYvb8tIJ7jP69vXprSprTqqKBsCPWF7pc9jxQ
c7SVKbg0NVjUbnvvr5Ux/gF7UfurNlikWtwHh3PGS6NCDoorZjLTkqwsbBMxRwiE
IklOgzM+i+K4wgqN8I40KdraS0qgfPATIn6fEfb9IUWh5FUMxALu8+ZRI9+ASkAA
V35SEbBqHdxd+wRQxbvSdhYCAZp22XzHES0k57j5YSd7qBJ8SsJqfTwqfjxw2O79
KYx16MySewYL4SNF1UM+ZS3/lQUefAIq8Xg502caF+37vC1RBVzS+cB3b6EDLC5B
0M+uDzKCk31agmUrihEEmdG9mBOnpEF87RW1S90S8fxTiuFACRZImpuGAK86Z7j0
4V/Z3OWDONTb9Cz3hQlJXAj+09t1cYWM5/KkHYf0ftL9s7Lw+uh2awSK4a6lvhlb
P6KLqTw3wIuHNxnK/TZo6uaIl6RQMY9NClu8PyDJTWHTpILz5fFixr1s4XgzibJ3
ld80W0iCp/BEffV3xLVi4/2fQNyuv75gGBzD+5cM+wpU9bd+ZtAeTMhQgxBwe2Ea
3RacPEHleQa5iuYhzaKIPXAzHaEjVdN/vWkGgJURshcjYi8rFRdDsmDjkfis0PYw
1SRLGZu8BtapfdHy1BvkXw+Bz1bAOAUy62h/zD6mDQZXNyDt9u6eD7sfIfMGzfgV
1rfb61RbrfjKSl//F9QJczcwWiIslHS7KorJ7b4CxIQpFVO7EOfakxANa7Qff0B7
z8vs8S+sWlCA9Dmhv8EUrdeVOnHJbrgH3QspkCNrjYkio7RY/DFX7LAvKTcqNbc0
x+3Tlc1ad3KfCeLN5jV/7ZH1kwwhk+dDMDjGSIqv9NDi1GXeWmPlxMyX3Vmt0tMc
lRmCWCt0PhjtCqDsQUVVdt6ZXfNVilDZ8QSJIWtck/GCNA0mG8HJE77GceSby7yb
fnXZeXfVNT9FR9HndVd4vYjzTCmqTBhIJpKzuF5MnLFubpcO5OklyoCYlbtfm56p
p5XRAyr50crwsawlwTn3Sn6NJPYobpl0D25iabqvM7xbBo1VJ3bbfADkrhR83I3T
rBExHM6uI5nzdsw8o2jhdyFdrjmujSh1LbY2ACBB1o22/t+wJQ+F0sW7NufiywQ2
4Iu+w4N5UEK40YJof+quQiiLF7GUwTsI+/jVcEKm5vl6lyD0WfsuhITbJL4O0/i6
JaiyKj61kKRGV6QnLsY9+R3XCoQ6I8lul4bXxl61q2EiYd5xgKK20YHB95/xppia
cAgV/lZZ/T2WOAump5z/X27mSgVuJZyV2EH2q2R/mfPrtESYy+PdMkFyBdW1lUeA
HAwAsEIYDSMJlGZqavXJsxmeLCsUotc9VJJ79SenwlcfuJcTrSf72kYG5bLM0QmB
u0S1UgdrsliHUMkDZDonvBQLBZ6DlErnHG24EUK0fH6GxmP/62XA9DQtJ78n9Zzk
e9robMhKqdkyTWxXgCOnQvpoiaA6TfNmVWWXRjM9lw8hVip1EOlsD/Rtz5eb8KIW
4iiksnzvr3kM1lpDQ8NoL++lYMlEaHtAE8ZE+HfpEJ7S/WQgVRloHxBA3KxfKMWO
sm3dZP9xdES6Tv+b7g9dtYQkmMFpKpQWW3E+K5d5quUl6TXppyd/o7gyKUE+RC4g
JIK6mPhyrLqNgSvEjxalW0/h50G7PAsc3KL6fGjttZQjm6wcLNPOFny9a9R7PUek
o2uyFnJRxwi6aoDgcxmI97udQxWysca6dgqh3UHOjYYAkJ4wNDKPUg/+AyN8h+jL
jUnuGMR6wNYvQa7HUHxekObgyDbqfHBPaq4Ynlshhy5uoMZ4Op2/Sa8AdSc9jw2c
XInpFSAeaA0fJwq0VJAaihMTyfv/zkXDHkv9WEl2Pg9uasytZvlWHB9Ygf/rMF6x
rxoGFglWATUt/gXmwk4C2rddqwIKKVsZJshTxH8d86YZnJsoQMZpRaT0/rI7VzZk
Lvjl4JLDr/w6fb8oK8rdbyBkmf1uf663latW0Q+g3r2HwJjEjxpN6oK95XAeDKLO
WgwqcpKIc9CGJzfJJvTFPaP1Mk/bye9GvirwG7GyYYO4iY/PORUZPbpa4HeI1kXS
Om4Ikiut3ZdIi/fa4uF9nYQ53Z51oFtnfwu881FPsCBvwBl2n63Xr7o1GuH5FAB0
yrOGJKXYwOA3Y/m6N2eQLrwixRe04xlF9BGnCV9tFVpyZf4tmkahMq3QKPsmBmZj
la4XxvaCyhlRFSI6GC65Vha9+vgQs5S+cM5XZf8+IBuOd6edeqRGzrC1qqUsbPzR
anNAGrPKWfhBrjoxJfKYTV+I5TEBaoLGUPsY3L6/HLNFnsXnqxbV7JaTOKNC00/L
b4rX3LpLI/2lUtGSjUv2XBdcVQYsQFeNAPHOhHgDHdnXfkJ/rymUSeOO4BAWSyHY
IEQVuY2sQWVuam2anPBjF/SAEqRCcmAVcA/2IyoT9m+Wc0RWFETNKNYnmuaDZdNW
DAV0DG+VC00+2QCcqIl487vsDLgiKQIDEK3zNzogkjuUfS2uhkcc2gQRT6WCDL6j
KslKqbuyZ0BUzKG+RLgs5h/4QBYs9ofTxg4CdHox4zOzlFXfWyxH4d65ghSJGBIw
BLJOjQ+9FCBvXP6jQ0aq2d9LV0EZPpOUgoQ33H+xPIF41YlPKNLnCLPSGEctwGf0
gR7fwvm+9EvLtQPXBbCjJgW8rOkOBbLMX0i2lqPQCIpUSKnefslZ1WyUUg8nBU/g
MM0DwOEsLS0oZkaLlSUYvvYIA663fMIhmKdsHZdwu9FMeRpRWnxYuV34bWH/UuyW
osbSGOBHfcMFHDsyy9Fm6Q4XEaOHG+xkBCgUO0T4a/0FCuQIFfF81vnSKd6IfLyU
aJCVV9QpuJ9FR/6JSiPirP4ly23GHXEL++yTLvSgKtrEK+e8FB4h6Lina+YpGAI0
L4kbDPqDR0s1LxnIGt7a0byvypV6tQBoKjaS9PkU+FgqIYXlWCEP1DxBzHfymvAf
V81Edzc5H0YPQsWjiXk4yukbnAcKiZvdvUOwK1jciHrQq7QAPw5x4BbsGsiob3B6
cmQPuKxd7U9Fgga7nJTRHlNKoFq3B5gQb1EU2EPbwg26dfNFlw1oIFa7l3WtFR5g
lxmvLExESBhT8ilrMKZZO5zzyPRaoIMvVeAr/gDmsAKhUgraAdVX4FZ7GKOPymPO
D4BwLpP2xjTIF+8fu83wGJ6PnTOBvOeD95mUCmiLoj/zsm5voZsZniFMJcYC4Ejl
a3PC2uempl/iDl9mfe/QgODTup8j8hSPnJnsUnmniUxOshM37M2bVQejbW+ulSCD
AMnhJY7GChTAXT9m1mHKEPKeZ7bEKa29Zl2kR0f40XFN55i2GIbeRX+gnJjHuzZ5
+e6fQvKNv6KZUV6IcWVp39vmOrzNtUmr9VFkK+KY5sZQcVzBQ3G0jKuxP04FOSh/
i/k+z999OlZqKqAMErlGkmoQe/YppGqpejY5Fxw/3lYz+jNWLiMvRcP0nZcnKtn3
disOCFs5wttDh57vNp8/035VPjj/PhrDOzTUboLRr2taPHXgG7EcwAMCE4Ap7G8x
QcEQrP+rjUiFdRAeyTFIom5An1sr9ivFGxYjRvLDsRV5Hb/ATINXT5z33+/32owz
yXjbhZb6CqHVm4KoABf1TYYRjBE45XTS0+fF74vrhrSIi+m7JKIFsnRnf1aLk4a7
YsgVHKET0FLGD3cFMi/iMCpM8EsnGUH+8uM1jp/qE4HTUEodFvOQI4zysnb+dj0W
EkFvnYIHsuUTybdsuYzhtFYFZBfSHv9+8awnfgacRNQzuHNa7kGYboJ8d5KEItUZ
EIRBIProY5Wy4O2fb61HaJ9kvRapUDlSHjBXDLuB6ccItT81DyW9YoYzwJCMHFAQ
hUoRwxORT/S2weRPIDH/dta+XfL16jRVnGnsvLN+x/8yhfUnhb4wcBhycjBoGjqh
CYLGjL38iKvVLrQZL4PB1XSQtlRoLQTSzihB9sh8l7MfmMmTeQPjUPzsZFU1VD6e
KshamnJFuNdGO6HC/oZ+1tVLWCUogWYnCkxaFUQ42FtRa1gKAhJ0MjVG3cxPjGr/
qFinSjjE+VH519cz3e3v7GGCOXyDTYUvGIwpG/RDbd4TeN4YPr4c/+hE5JkjsjDU
CjLT2JfjX0+hyWBOQU315GCWWT+RwZeMRJeIimAfoNxE6ubd2CoTUILdLWsR2wh8
jXwq95jvjujfvJOwYLKLn/7dPysXvz7m5iNcQpU0WJ5J/0gJ9rmqjrtnPxBDFHrZ
2GpaEFcOPimslMAGE4PIQ5+0dcSDQRJn1NPEQALEJa8wnG1Rx4oW+gjs0f7dV2i2
zQSAUleOwHcxbHukVrRTNZSPaHFHvdcvMZn9V1PWhJzG7oJ8Ef20fgJMxL8223dd
tGVl8m9hEb74CmvMfeQO6EWsYBWYwgQ5xzkhUXb2+RImWHCcvTlT69rhzR1ZoDRr
ezb9FldeRRc47gcbFBvzPh6jsw4m//uUFc8HK5KG9WM19KlAhBMGXLrLEnCJ5U/i
7BMq6GMrjJlGwstuOCvZpuh9RRHltPr/zwpfDHvdhptc2kXENmuPmqQWODlJAe3y
ToO+17zH8HI2t7UVjjmyV1r+OO3uASRHXSdrRhvVukPq7trm6eDDmuBAvSteRdGb
HqeK7Sl2frNzOWt8o3pjDh3XbYNhC435x1Yeteu7o+hlGbRWL69LzlijTjX5S8Wf
h5/yZsUlDMHgVlj0RWqzVccv8OtZ12Z2odJ9ok8i9RymY19VrLz/1Z4Aw8Sx3tdE
ZLdRYzzZtXuQIuwp7QJWKl0/vcBX8RQ4HFAdF8ybIudcdwg15I3A29+LJCj+SOS9
hhxcJsqyO189srtldCx1KAKhbaLLLMjsBWC5D2ujIgpYSMLw5XFWdHG8ZhO4PtGo
RdjpKH+rtY5DRZeboPOweUdnszhPSJRgtZcKqWTB+hM18U86UWyPssr8Nz3CUIZr
2qq4MgGGBIOiN5iTskIN6e4ueZRj/9DuuDEsvojA7MnehWWnTcR2w86Kd34R9cON
2RLXh53pasbslO5zJkNpViRwgk6t/X2PQ6bvA72LJSuYMw4QTfrvNTzpCNDppRYT
8LD7MQ2YdYXI+qYe8H+hiKc4NTnf2DiubcDvgHchJxZFUVYrumnkNUXYAdCbXA7Q
dbSyncwjH/DFgDQuZtazB1dZZzf7ilR7gfwKzby11CyB5gVbh6kA/9AjgdupVqm3
R9CburXd+dpZ4upUexObZXzA89d5DbxGzwl8+WlQ5c1IF+YVppEAOz3wrNJogKa2
pTCFG1KBz4795z5gJnkwhTT0qv90ynJ2gQcObD54jOIqQEhtYS8hCetcNmGrny57
YAbelRvzG346AnOhwNpkhz/KUqL9USCd8lAF+pa/DB5QWyBB+YRSnsLoHIVkHPee
e125+CRlgP5/Z7/4gLBuHmOwNy1jdh6ugpq3sdvVRqBG/ZuUSH+acckrE9WELcW+
a9gCVgOX0DmS95PBfvV8fymq6O0g/DUTJa8za8WHmBclNejSPDXGxku2v9GIX9/s
VvK6DMA8JIcdYpKgAes7Qu+jW3JbkCgEWEXirkIpj+vjNtoMZf3NB0NMLIz2NXDO
+9bAT7W4zAyhskjDdsLVtL21c4tn/H18AF3SDPbdttNBf/VuQkAYP5gab/UuLaGr
qVsdzCZI5J76ccuh2h9aHJnGbPBt5D3amTrozLJTfVOIZtP6DieVmzlrg7VQtmzG
14dNzQhN+VwDzbQmgICQMsdNmz+K1Fe1Btw7CiJMs2CqVc8GB5++6WeRNvJrCLDt
T/5ZBhb6PAlPBQDdJtDlUpCiV0nLwcl8URU5ASg0XVbPbrTNymnWU9Y95RBU7yvt
0xLY6C/F+8dcNZZqjfovz64/OzpxGqCa/eI80ZtIL6Wpud5ZGqIKQwsOMnn+Gzki
Oxpw+AsFc2WMHPzUkcTsmp7Fdgt3XEGfOyKwMMkjJVArG5W+OEI77wzzYdBmvjzt
0HOyflyY7fZTKl9yNURAnIRQdvgiauXycvcvujsRmzfRdUDr5EuDS4z0Gu/Ocd17
4W7CHLsfMw+VFsN4vUwVpmEFXsSAL6hgdYKiF/uc6PNLddlhv9jvSwjV3LwrUI8B
aJEsYXdSBIQX4NHoZFRI8wrV6HMlxCLvZCN97nM+oH95QQW7SPOjjrm/rX2JxbF9
dL79lP75NnPLXHRvlc9Iii65+/60yCrHVN0qU7zX8gmiplh3dy9m+FqYSXyImCss
xgg6gvqbILzcE52HYKk0gUFXdMG7njaJ2nhX4mYJI4HFz6x8TSkq3alk2o46n/fh
YGSYhA5K/uc2M3U93DDLPFsIrb9AAb3T0LVsga5gD+U3adZTy+tdoZQJCseBvsOQ
xw/GtAry/5Xo4/ZFsyJKQQGnl6BphJ7F7hFsHsvc3d5B6/1QbbEcvDcafoyVXAxo
yBhOtOPeTrA//LGwM0sWgkwxS/zVLkj6K5ojXyUPHe6BTZxjxw3ivJrP/UPEqdY+
P1q1BR2FkHUmb5RS22sh+9vnGfD1mI2HBKPEGdvU/f57jO2f9cdK+Nja+wn6H2+M
cbpC+d6N+6Dyr2JjJWJX1laGRTCR3y+EJB8t/4rJbL58qWXIxvW3bBK1z1a0aMiO
w1aEoOoaqb54ndt0M2DXpF4wP3jX14Ow5ZfrxJSD2pFRd6IwsrrnQSUR0i5o/Dg5
Tx/ltuDtEmwCWk/er9EvUuNsEaGW+3xuU3gtkB6ZHHnZenAGWIqtu8Xm7tFl7dM2
Dyje0Bg9c3u2SuwCT+NrlRLkSBVHpt+TFs06MHjXwKI5OSkCPznK6thKlC1EYVw5
FDAV2ef+zQDEg4NBDPeLcurCJuXjXbgk7pF2Z2JxDOUmQcWIcm1ZdDKTuc2fyunc
V/zcuGFebAEOArsuFRqrAQuX/mNcztvbay8deHzmoVFKSz6jMELA/rHd/46tn2PG
AR86/KNQL3lcnSkERMzosbDZS6h8dNgLbehf21lSG4sZr8h+zEq2ksQZzh2TfckO
uUChWnSCH0K4331waUL7Ny1h95dKwm+L1lgujQsf4Hn6EjzEMBd1bR0gb0jCKo0W
53hYu75J63bmeXEAqXudkBG7uk4AS8yE7Aim1VEybmLcqhA6pa1TGdZXmyo6CgSs
3BzTvKbwJuJrCR+ecy+QW99/p0TIwkpjG6EMK8HfHArdYVILuP2ZhIfgkTrOe4nD
8bAhkyRyPncoRQd6oi2JxNQYrcfQlDX/ATGVMtYurk/+Rju7wur2/7y5hBIIYTPI
TfOZuBJ5cpAs9//+FX/lW9DMMSwCtO61dI+IJOqUaZB6PuzwTnrsYqgJt54BM7W8
C4+ZDXAXgDFuirq3Q0Wxlp0b6SSrDykYRLyESZnYOWUKn7YwSQEXMIHYBxZJ2xoM
ZtWGzKIBntTYl9jA7zy4kUqwey5/gJJ//S8nyA2vl5QLqtpdPkeEJuoVfUPZNl8G
nsCBdkxu+k8w0nTXq7YaWzcR58j+SoZTff/tbekuXbkGC76UumAz1qMrQRNn32rH
tSt3i8/cdTIyQ9pnfOy7yua1snaybf8KWL6LOk0PNyLK8Qpmx63/n1HyQafG9QM6
fFyJytl25gm+wBQDndlugKIBWME0SlgDTWbUY7Pm68xqIR/Pqwa6ftXXDoabINth
z96RbAo/wuOCNZsXv5GCDsCuthh1UAusk2YTVGhDiBeK7f1xp8LszCMyhNwzWn5L
6q7l3ZcKov9pAP0LrzCrRN0pIGNxzNp728CKE71VpR081Bi0Ku8wfFqV+JlRypHz
PdpiDFVa6IVh/ZkHQNY+Q5/JmxdynYe7sxRyLG7oG6X5Z+jBX126X/l8lNs531ch
oPGFpXgkPYKF+GLjk4UEof0UzCl+t3CmJPbi1fmoNKbGZLYFTrStcmqxJ9IxjiiR
sWHYuwvNU9ZGAywbrVQmn6WP0cRSHl/v2G/oN7FZnfhGRg7z9ybohOFKoolEiEDe
pz1oZAXH/sUEcVeaVnKyrZDWR6wUCvXBQ29cDBlAFx/wRDdTvml0PmY1sexUUnue
mt9Hzhs6dbGThjGHzR3LHV3bs/crRviEMWXQ7cSTZqPMf1aDyOQuURnyKQXHp1F+
MqwgmEtJgL8jhJLlnCuD6x1PPXDhtvqlwXtzd667cmAffCPszVcDTyzaGv7b+lKf
me4hIkTQvIx2hAzwuZiN8DGRzTZ4NSN5y6aDNvnTUgcxFp2TkaPAuB+eWmBJkZny
FWlLGE/m0ksSiCdGFwig/K0g4V6xS9kLqBgq+o5wv31IFd65mJBxm5vaEtBiE0mb
qAQC02s/yCF1RULITYz5OkGhPeFk41OR+0l1BzJNfN+JH37W/wi5mPJv/GRgJFTZ
hQyR7+m/ckgsrsg1XMxjl6zhg0y7y+qQfhnFcWMqT1LHFtCVXNpRQtx2UKhXr3BY
BogYJs+YT63gEI8ydMEFEl7PoM53Ac/apwn4uIsyS87VaG+IbmPz0r3e/F4DOXFZ
RfImVh7QhVyt9LRia60urnMVODJ4O/EYfcuScOfADqi7wbIczmHrzHqZPrvfVnA7
kOYu1HJEfJtYDz7Un6o3uDJ4qYRpdNigap7PpOAr6hgvfWzWe4Wx0xbYhnJljxWY
mVt4Okei+81hC7Iwcqp2fud23mHMfJqA+9Kx9d8BmrendTb92Vk78zfq51t/3VQP
S61OM653WT1pj193VYJQ2GeWgkU7E43VVkmoFoi+7M2goDlfPKdXleiKuz2WZnoF
urh8O2mbgsILbaPj1FRiMMpEEoLsC8UgGSc4x5H2AS0QwiTn2U3gdX9jsAXGSQUu
7/NZudh5ZCdfM6NYtOHB1X8fdNcVogGQCdZMJLVUTcVMMuq+1iUmRPYc7jJQmKgl
1HCO3DsHFDK6eUXgd7wHJFWmoyftCoQ6gyrHDTfEN0En/hrP1bmI9/mH6PVaxHro
+ms/mYKeHI9gLKUI1sPI72KPyO7KNzDksidhra0jYZELktMqaJobXaQhIB4O1YVA
RF6xdDde3hw4v9yMSFSMvB1lDg4sGV3ZWu6am7WB3A4E3R+fSbH5/uLZrONjgYi0
E7WLlU1r+RENs2TVPobBVHr7wJVjJKJq7+bpTDgj5A8aQv0ig6M8idFMYZ0MOIpl
iNj2I1e6mH5Mw2EeTxbpCSlsucc+lCISVFuo+yK9yrLvKGFx0gXrKF5xpNpdJhob
MglMMlgFqu/GPAmwkdXdHDPFwM9ASM6xXE9/jAJsT1r61xdu3wS8mlH8XBwqkIA8
OabCHpKqw8xdHznusa9s9eRGH0qcRoTMcKIAsAn4SuVLc4noxDG/k7fHiRwO4hB/
v/j1QESed0O6f/P/GkMXGC60yrYjNt/QvJqW+/tBLLcVGixRlwa68YIZpnxu/pJz
fuCj1aSLwTfc6oc0oZlBXgnmO2GIQOkM0LDfLDyWva3MbEF+sznLoT3VjJyWCKyx
NUQi/4vxN185cdNk6oc7DZA7hQfrm7A9b8HjiHt4OOunJkpR7FNRpgWn+HouUZMa
o8xu1dUWdoKcXRr9IqOuq+YQSuSa/nuMjoTRMuCn6zhrDjv8d/0ETYes2gOBZ4ou
JnYcTvv3xa4VL//yIgOWesiYOhvlV5LjbfpaRD9DoFRDXVDx71WjGwm0kBXXx17F
AMNl3i7sGDjBGPYc3Fg+KNREU62PayInv6pd2VB0Bp7ino5HoVGlso1LO4umnMUN
qKMQBhYHihzSvC3FV8Knl4bhaJdJJl6KV13QXHjXiwxX6wx0BiTQpUCx55Ddzgu9
qeFXV2KVvg7C5Zu2XbtL1F8iL93cDi36yz1N9FrBgxVQH1W+uLbMW2s8BpmfYVG1
m5d/qF0MJuGO82qXhZCMWLG1/7xCkcDNnqjLU7UL0cbh6NipHf+Iuzw6CWpVTMrg
4R2tMXOHiwvbjKH1URxBJNHs/PlhERnBZVyVtYMDQCmGNBbue2W3lGWU1v/Ymdvt
Y9odGnJ/JIvCGpsf+7lVPeXhSztXpju1Zk3ijdlqkAt503OuWTKxavKnvBDSpg5N
Ik7ddxPOxnAH1pM+p0HD/07mgrdUO3xcbxangrRo4E87QyReom+1hpb8wd6y955Z
9kIxDMHBiy+h+ttqzCbGNCUNj+PMTX9/iSkKVHCX5771eSl9SUsDpD3O4a1SImG8
Ys5YDfpscSVqBfd8bwrkKtpvJgKQG0yuIcIytsA0VOZ/UciDR71fFT2y/u0GT1xa
UPRbkIdbqlDr2rs5WL+qJtmEoq5TV9wz/vZSx/H4B5X6i6AJqWPjNJ6XhXkUplnB
B+AiFiqk2vgrvVzzYBUKD+z1he4KFbGzo7VlA7jmVbWy8lAyhqhc0GRwpuL8noSo
ainNMoVvwyC4Lg5ka30gnCUtvHy5APkVVJ5LRn6tjr4JtYxoOfxCUzXBKq8GunQN
o8XERJkgUSblm7itXTadbyZjjD31zZkswJn5kQJyQeEgmjrkxaYDmCbgWuyyMAie
fp0ZI3zeLHLveNFHTlVsRyJ/bEQWmOXcByK9E30xeh5HPfv3VfOYGf7y2m9BfM4f
vJlzEXHxcJHl945thUHKXeV+yNSTYPwXcyGUlQjALL6/pFhYFqsJnrQucyAJcLY1
jsD0O5yNfOosSwTbScbs6rgKKbL3k2f/CLTapCvxTMTSg1qQcB0lIHyl46kbxi3e
dRRTQ+lF1qFgAsWP2LIwNIwpbQBcpMMP3RO5/71rBnE/bDcAJ2y2oJEqAtcgPPT2
AA+ITKOuTGRS2gLrncNOsWj2JvRPXB0NLz8cvZy/ordIXVvU34j51sOtbzsy8nrb
IPLaWN3ZMfPgmuGt+1wEj1fChH8XcLgGIK9iS3x13r2+mDxe34W7WL6wU2MixATz
mkVidq/D5MK+0Lno3XRN/dNs6Vaqhxuk24BWgMDGWkzY6duH9WaMgrUk0uy6oYRK
h2L855lXZw1nvdLH+3QMGuBZwdzMyJ1Ff7l19Hd21aun+AZyG+x4QhYyoVl2q0F5
2s6tjeUsbYs4RV4O8Fila70FJ6AezbEkjmCnifNJpOEUaKJlVFn/jMHwCKkr9XCT
WLnPBGm9j0FVKesIZYIPYVpjm0QobAmi6CmNyiJzNjNFpGg8LbXSVyXoTri3jBdr
g1PZOtPziFiTUV4VSonq7hd0r02wajkeSlI7njGNIpOd+iYLVV4A+00DuPCoSmWa
Zqem55GgdcgahA/Uq9qhTqaNaHoNT232BfLiWPQSZ+f+sGOg3PBwIaKSg50kOeoM
+1/+YmawDbv2gz9K1UmQCun7mw8Tz9inU/puqcR4FxFd93vhXn0aD+SU3fS/Tjq3
fEBCWJCseqztIwywQrspZW5qZu/6KVt257ShiDU9SBpDydizLPCvf8BmcZpSAbrW
vULgDaS8q9MKaGTRCLS5/F4xYPY1wdzsmtXi8xh2f+68fJcgohYeAkMgwawHBMmY
B7AALR2+2+D2vkLDNkZYGpEDRJQS7ZRl0JXqsd/9lkXGZ746/fsc+wQdN4rCsD71
y1Ne2wbn4+NLLpGivSWkuODiLeFOVUTMkS6wLgLC0CmGqPe47N9AP3fgQMoleURg
K+WpQc0Rx2M4wpE3FQhtwWBP5x+sIRjnRAmYoLhSQmw07TS60RdpjTebCoQCT4lU
+FRrgzb2dUnBExypfLk0Gk2jyNZ01KMjr3408gJ8L+5pE9uBdZvPFvUVrwddAWTC
M0Gggdt+VTiCrZOvtUk9lK4xEH2fIESK2glCbP1oKCgTLEjIAbPEs/SH20tuOgkY
x7Z2I4fszXucp3lzOe3jQEHOeTKHeRosdOUzgI06c0V7h6e9y4ctGyskLvff58mW
VYaM+xPEuhWb4p8Ql/NsP/xUKYnhz+5XWqMF85A4JwcwV8md7/4Oc07fJpIByB3d
ePqXHpQ9DXYaS1cVTfGt5gucKJ1A/rtAzHJDow0SmxR4L3minivV4KdG7V7PxXvl
IWl18WMxpGcprWZITI2hiQbxqWv2N173QoUnc/i32tN+VYTIenORDEKnzmQ4Znde
n6JlxiR2shMbASX0jxklvVdp6d26juY9cMn/bNX3N8wvU32y+TP9NI9Sb72SGYE9
6+cFP/fv/o6VgOxkOdyXp4fJ4tr68g3OFUaAnRHEpg5h5C8XtcxLeHJgrQMpDBW+
eazsQqPW7tZF61a/gK3ULqwcJE3Ebml5BR3UOyTvJgbN34iZi6WH8si9AmblyVoW
Rj9F1JWDwzo0zmuImenmDEtvUjmlSwAfIekGv4EI2RWv8m2T5BHGTl9GcNyDkhmy
snEEaUKfqmb0zpySBkwU4HIotx5oML5GuY9wd5uh3dhDFwZtydW8hM7JZ1LTO3ix
zR6b+7OFACkD6Cdj2jYp1wYFItkJ44K65zwFiEK/wB7VZiZhLsSuoGQ2CuicKriK
gepGSnhnEbZAPraxmrTXTsupxCJonjS9iL8JNEJ43DnmN5Y26DI1JS1WprZxpvV2
mgwzsdr2+eBmxXD3S4nuDbHBHzAc7ZQGUaufRvkU141oncXP2XJBXpOlf4SQUumU
Z6RbM8VDEV9iGHWvLaJtNbb8162NvVJC6FWRQr66xnA2rgWthvdShVqR5fh8nn94
ok49+bMfuVXm2FQkWAH+ptqHGjRoEhaPm1sqGgKIgLdguZJh6MTDsFD38ObR0r0P
E3qTqFgNFQEcVO0uSEi1fcVkwj3dIM/Uy3vWVlJcWOH8PwkHPhuhousncLB05TxR
Qp2rwWuww1d+SGi6B5pDHrjq8TRixdchXp3dSuUdmWOEJaX2ak+N9cU+1NyPVK26
SjYe2NbpKQBY1EZDudg37Hn7aY2gDtIRQ52miOb4Wr+F9ayGj/P1s6uiV0Lm7xQ7
KPIxDp1BMPJRfE7K4TdtusrKsWi6d/G3togNiCUbABn9Dj1tKT0rY6IKO3xEnXpV
qmURF7qQ7qlvC8a04IciCAN1grYlD4AL2zNbjliTP+tIjbtLBnSekCgGxkb4W3Ir
OR4P8j+mF4HXb3WrrKuxNW9P+KTAvJTYCe4RcfcTYy+dXK7Oiq1ELvRJ0+HTat3q
I2oMl1uMHVlGR/m89Vq8IMbxXg7aOqCx8W9I51jhAS9DyFCb6DpEbl/xqcvr5xWE
4p302262i6pAtAkH/OPkAnd9fk2eyMTI/lDlXUE8yLdSSIaijaImqI2xUyQIkKcT
y/xx6lxCPmKaCZfNpu8qtzLHMTwXICLgErw2f0lDD2b+5MOW+HVCgz7s2feUSKTl
DTtV7d03im/iBDmu3i0DcJv5voJiyKSt/uw2hCu0cddE50lER9Xgt3Sw1nsv26yO
uqJJ9K+dW34qSK12pcJi44d7O/Z7QFQP5kPByWI9c5/RsF+oVAEbqOYWRUnUgcyS
RnY0IOHwhLufzTeQs1D2yNtD/0g/l33dHwJcCJMAEPS+AX3loKbEaqcgYPIhEddy
fW2q2UivIvjfgCW0eo3EMLyWJ6aOAUv5TKLF6kwvMPB+7lQacpkueLqoBcP6YzkC
VCyBmaXy1TTfErw/Uw66MKjpGiEY5DPU5jk+DpDlrMetyhEZ0fvVLFFb7PwAUqOM
n6Cj0uS6kpeaysRBpZLMXj6GoF0yvCQG20ZdAzyT0zJsg+lvwTgmbPfWLF9vDonp
qgbFKCKTh0nwQxgCjuy1pHzIwJSNJtvGQJzSV695Az5o7fYp64th9gw76m6fTSOz
D+dMjKem7OxF8YB9KPAty95nO7/8khtYG2mj9UbcGrqiY+zKrohy9+B7tk5p3taQ
tNYxpJv5vFCtcGm6Hyp+eAQa7r8sF33QXiOGbIvqKMUopGvkZ74ygfiGKdYDR1lg
510lef1i2NOHN24mx0KaVNDqomhP7XOJhTyMjkGzFRlhVVXm0Wakm7iaGyvAzQcT
bPq4H3v1m6x0BQ3BFHVY/Mkdu1kXozsoxq7jXdYwNhsuDC+WP6JVUcJqkYT93bWu
SSlGGNUzeq+oLkXQDZUmhNyXpp6lVjAWFtnK0sO4qChjFh4rPwEG0xY4PkudhLUA
P8IRf6ZTmwXxD8NhUHJQ7HqDjHEL/Eie3sYuzI+L1iqqQLpwdtXjWH1YWR/YFL2j
mD1eXV9qGFIOHVrw3oSRosOINSQD1C/P7rPDd6BPVau+4j62LS9+JmtvQoFV3Jwd
Qu0/3DoElXWpWlo3uuqyHMrHzn8SnTRiW1dTQbdLzBtbx+JhWbAAQrux5twy3VuL
KtK1kS0nXN+yRhkJ3o73/uvD6c2OCyBh7oQfrmazzS1pOTqdHx4zTrxhp5+BG7W5
+WFJgLMfwpE4RPaE6vy3Sjhpjg8obsl4zERGIcECmfItHpYOWresvmppfZOjPjXv
7HEKF/kxW5OLQJrLptLwH5wgcen+g6OJRHO4wVq9/JTta+iX7T2xx3BS19jBXNhG
idKu6DJWetIKjRHzyBqvVITDxkQKcncO/G/GYjdd8rOqyO1zsY4c2XmhqdyHUEix
x8cUlVPFzzMVlT3IcSQMLSbCsaE3aaw2VNliMHtsIeEoGlNfkTMD5Ts14v8Naguu
YJcymQojM8wDemER4WzzM+Wzwm4Nq3/ElgGUR7x531ILtXqNyLv38IwzSnmK7X2J
DnGzWmo/FSQg6nuHgy3WL0Y1a2pyLq8a+F7FJOe9yM8ZcASQfKi9MhJBD5VTIQNN
P8cHHJOT4JkiXf1YleSzE96ROO0tiTJ/D5DLFJrJZOHtauMEHdCx/UUrzhBKxuDX
CjGnTVpV51oJ39jpqynQNZZPKwzVTVgm/g7wJz/nV/M3oFFBZR8q8smpFhsaxmkP
l/4oDAZq8XuhG5Y9aL0mE0RdChI/TSo3zWcbESCs+rlmHgwKAhnwJiq7UQ6f/juW
LDOK0QuI/SRCRRFJfkUhVwi/kvx8o1T+0Amvuviaw0Vfh6wzPe1XISPYaTIstphQ
EyzXBUSqQu+6kplBcvr7pSPMfJVLvdVL15k+4cyzCjvONfF+bZUgqczg1xCKTR+X
oL6aJKyzaeJURUUgb/54qLSRgKOKMf55yvHRsRQRgBqV/cgRAPKLHxEFQ5At1XeP
FTujU+hBsTPr671VUdo0TU9M+eklGuX4D+34/LoA7csz3tTPtsMmWGABP7gkVc4K
SRqiOeQGt8A7o2d8kriwwnUF4eyFlpehg4zLASM5oYRPebSXgys+OzvQUEvmpxDx
ZZngfZWDwr3TTHOyyVmtKc91emT1O4whj9uyjRdd6cyJzoWuq+JmUQ3T2Bgukj6M
B2PP+C+nH6DMs3N9Cv6KEIbeaPU061cs2g2CZVmbGfytZikQ/bRgkt7dp47Z1xND
YVFMHA9UQaAqIFU0z0+Inor46TU9YlRD/9OEM4FBBC7VYrKMSHRYZdppOX0Al9/S
TtZHNdbXJ+HsL3yhvVVCOZNBqIoS6jpMtAWLhtE6aEDrwEDIeGP6n5Ti/PKniKEf
QegK1PhSmVcxDU8+lz1bAFBIuF2A7ORO358ez/6ON2zne4edjnr3bHhypnD0qKTq
TNDBktOZxFrPJys4YhZmS/2bZ6WfmZ4Sl/m40N3xEF+gSMwFqLKDLDS0ywWRHVlA
fxQKfV0Xmtw5cVfKMtwz6Fdv198lGpV+4INr69oL4O8hjeSJSybfQe7so31oYV76
T5tQ2oQ2nXj0n2WjnpfTlPAGhzfNDl4O7ngVON5hWGoyFkKKHVWN791EwXyw7Mrv
rHRBjzPTIYOCe1KExsQIrmefeg96DsB1Tu70evtJz+2uAS8xihQHjqx+1fzeI8jL
YdTM2rnSDq/Y7yxEZvZZpqIBNZ9RMdRPz2l/smBugVxwisZCX8uQDUrHXTkiyUKd
o2/YPw+OdEpuif773o4rjm1uxytEa7H00o+vZTGWqrUhiwNTo9EDY1AYafVsw8N4
b+e4AZaYoGLKAkVsYBL/EBZTRhh9q4RSD6AOPaQf7I0uahWV9ysFMAFCqWTHEf4t
ED8QkWcb93NvvTiXZ6o071FgCKblcFW3KcyWx8g3+j37FZkuu1xaQsFQSQpeWFYb
7q1I6x9X052/kT+n5XQLpxXMOFjzCgGiLf1xj2VQD19rUnica4i4kuAAT4dMpvbh
JDFTHuIzRsEHChKZdO53UTxd60nNTKnNVp7g4EKQcHTOARvpRYTbhhgDdauuPpss
9dFMfTpGoCYNfhigQHz8Ww84PZdGDqn2Hv/qi99weKbdWhqQqx8zmF1aGklZMJ0X
Y8EZJJ6qVKD84Ydmk5ARXqz5SuqapEsyKNcgbW78e6XL023YWx5521yR//PHygos
/sPmr70yGdIn1rDNrjc69s79jZ3RYamIrP6u0bMzVGNrItyvrNnoM6EMVhQ8NyJF
6NSl2DQicdIyavt4KNXVBT05/SHjTH54QCqt5dloS8LKQLkrDRZx6Zdm/RNGsOm0
O4UMgtOkND2JRDwZinvtd79B0t4vRRiVJkQQ86dx8oonRGJejO76/JteV9/Gg/gl
TDzLiGDg+evqRbGtxhrhSvVoGn/OUSxA+iHDx3EOrEoF4QPmnAFYz3oJOaTiLkIJ
UK8Xgi36HlE/v0WzueILbcojXpHQecEP5AIHtrQ/d/+vGgojyEX4USdWYgcc5cU5
7p+OgpXTBkDOe6xHc7tiOZ8tJ3j6O2TfCyo44Xi2KblFwx5dvMESgDRDoK3+UEVX
hRgeORO1y3f6y2NkTUlQ7s8Zh/GrQk1vd3biGSIVl6CzteEGIXawq3HMZpUeVeIZ
7qr3mg8h4WTRdTu48AY1Bf6zxuTbqh/3kyxU+CLdcWXfpWwJoskZrDSQJSHq/lrg
ChMpOiNtAEn+m7dgalPiefRZ1L5I9P6gv9+MQWJX8jboi3n5e7HAZmzAJXEFRzLy
Jtjv238EdRSFiUmHvkeYoWCxPqYqJudvI8zxH/5pXd+f3DC0zsKqiIgNZau9CXTn
S3QWOMfmY4KctgTjTlm2LLfZ2cE4//PeVT4aMk7AKEMDghqTYP8xx6mLCPYDRP16
H/Qr31VrZotJ2xdDMRC1TQ1kusDW6HvUFgHy4kpzI07PY6fcoGlYaMVLK4Jgs5Pv
AOD96cgteXPZamYgylC3PluzF3iIBFxz3qftDoVkaq0UyIKd3bZoygWmhRmvg0QA
T/6OLrFGspR2qKxrK0Bgl1B5r2+qZ5przdohdwl3ZTqOLq1GS2sMOPyNb3OtZRyZ
uiezV60CMtZmzpkL+pa9VxBjM/JTUCajxKk4A60o493UH0DnD36XREgwtQecTsDg
4tvpGV94S5Cz64eobrm7DHHGBHdYpRzrHYNY7oXMldCnSrB034IBbKId+jP9H40r
TwYrW9PSPPJ9g4dl1gn18ywbNDIUrXW+B50jMIcuJxc112ofAYhe4xlM5kp7RV9c
hZQ2+FHJrHXUWJOLGXVPHJMXtErrXSibJkZHOrwI1fHlfcJp2S0dgkdvCZ9NTY1u
mrBqSkSiDhI+qgZTnzht0OMgPsw+GMEEAoCn1twJPCGr7PuF11j5vCYZgHyfCDAj
J4RLc3C64LWvvLnY1WMbjIRWly2hW4UqVL67h9md2ghtcPMOZdcrVjaJ4yApGGiw
YncuZqWDqycrLN3JfPgkPGoHwE/cgP5x2C9dw3oyX24sdux02/YMyEMk57uPUvUk
5YO60xlNES0mb6cJhVBvRItaNyu51CI8L0knN6NLf70OAQ42zvdrf5BehjtQdlN6
i1Zdz4WRZv+1xq3R7Abgasi4Qu/lai9+hm2zj8n79E/5uiQY4PTM4xtRRDiWUX29
VyVH+wIBW86hkQ+hsn8NUV8XI9KtiNHvviOvvCZ1eMbZvx2RAoI20qr/0+3w08H3
RO6VS+uUF+EWBNFYIi9x2d0d4bbEqwIAFx37GjA3AxrGwZcGMbnv7SWgGIslM7/L
c5SV6OqtaNpPIoUp03rNmwrYs70TsWa9BkK0a7tPEJ3J+zq+FBs/Litv/Fd8EFDZ
K7ETwt7rPg+4+os+fVBmz+c75v3JBo0seXmAhNzTQjKrN8AZrqrVRQPLGT7E/DJt
40BZZ+W4LtaHkXmjhdyxU7bHp/iNdBZ3TphJ0sSKHhE5I87XGBYilz+P2r98vqD2
/wsIN0p25gZHi6sOdwEniodNo5N6DItER9dIL3zL+Us+78a9YJYwnzObtpq/PmcA
C/Z43yg9HD7BCWs0rm7YmioFj+HGxw5Vi2Y3o32wScdLIB5Vb0x9w3kTWRSYzOtg
AOnIsMK4cPX4fKwXAwhEiN6Q1isC9fD/VygWV+AsDMxhyNqZ7/xd8EkJqiK4jlTD
lzjwvJtKN5AsTVC8vO7qAeHqsncJ3p+CTzU3sPG1KnzCFNZF8GYkt9l9+smvhoL5
32Wp4UXJwtSZvDPskMn7kR376OitX/rfhocRKe1Dd6HMNyXRJSSNXfVYLeptrAx4
RY6/Iq04X8g6JzgLrRkMMhi0vP0AuPIwh/jVxP6PLfqMlnhWOFOPj5c+l1TLAh0W
rbItKqiT2elhLlQku30tNIIl5Hy+S0TPryRofJ1GUNh17I3we4XrZschJYKLrPWu
l2KOzhs3v2nFuhVQqbyj/nDqQe7oE+NE1AJpzsgvIghPWU8/nE/w/rvDf13AHX2D
X70vjarTS9Bdl4PUs1kWG8pXwuWdHoav+TVUbx++InaCgqctroKgLGe7Hg6PisyX
iC7N4dufTyFs282Sv/pDKtQxQX/+j4skys0kXg4AraRTbk0pC35V0tynPVRsKbbF
j09pX2ZD4EXJwToZ8zYpzpOv5NmiwzUahPhDlyT/zTVSPC2MAUCzIhsm+Qdh/9xP
3ImmRmR5QqP1HCw9oE+pUozQBDa6MJ8qyAc5F+2wS9HTk+/NZwLjUP6I4Jb+9v/F
68fyvreoas/YVJfdl/BXSyiqnbP/4pK12zBLcr/kry2ZCXCzlS3Gu5LGT+I80D/C
FkGr4FatUc0LoFL0w5pAyIh04jOByQQyHkmfAF6al6uGknNLyLyuGlDJToCb7GyY
cQxapeCV26NoVvjXLQ2HHPW/u1lWZhRZefSnVO16zbmDAxCu3CT+7+9vrJaulqyO
i3HhiYDgN5DzU/RdPilvokdN7qU0jjvU8fE8AulsP0T3NiUJ7pfrhK1daEOz5aKr
jqlAHZ5slsLuKsjDjWMHbiVMHecFmoCqGVGR/oZeEshhs3Z2PbZ3WxCmMWf6sTXo
CSyhAy3SjIwUdcqilCcrFldSSbEKbnYmQyexDsa1VzsmPCs3I75R0ZY1hJLQkwZE
MbRu2Gh5TaNo3KUOlUKm6Hv0z1S5PstAayfXcaMyiDSVH57bXlJ3PyYSrz1flvMs
Y9PIqJDxRcZleACs6fd2ZxMwrcTD4LeWanqTd2sCPWXqk7Eq2b4Gl/WdI9Xjgrmx
Ilh6NfEVO3pMvjsR7AKu+peBpnL/lN+Tp49bCfrCixGJGpYsYOBvKVjaN68X0egy
qMz3+RCVw/zlDGetE2lA6Vv67Ki/7yb+WO1rRA3FQ74Hfg+9RgwH/5NuGfXN2/KH
OoZHIwMz4PtyF0Y7qpnwCiepiNAheV/Ho+L+xvNabq9Jrve30J9XbzMeFmYw6wQX
ZTDzqdZDA4xG1ap72cRBgA11FaxjQjJfqb9tYMiduene/2KqZp3xFqRqTT9E61hh
iQMdkbpyaapCm5kp31338RfrDkCuAjU1WNjKjv9cHIl6deT1jfSo0Cs6dYCc77tK
Y4n5H1Ks5bmrQTaojG/oS1dA6UbCYHuRoljWfsWjShlCdEUU7yb8/DB5bBQvTUzk
s8mT58G99gNGAlG8D+gaZPhBvoJZMsjlP7seThJm0NmQfcWjeR+hodTGysVRKe26
g8Y2E3fNm1CLscafGy5mV8um/bIZ14guXv7Y3aVWBcN9hCb6VDsz9g7uQhq9x4k7
q5LPIlUXzWsOhX/cbJPl5c9CDwkgAjhseCTU8DUVZzsEIQ4m0jWDVEbIhRzYsiMO
/8Zdf4FlJ230KlDM/pXeeVorPo6mvVXhmOc63L2O2u9rgRhqljjC/ZjfVj9hsUtI
ax8UrJoqoTMYxap5hay6GbiPERE3V7Yj43MLFwpQ9KpdqQUcgxb/tpoE+aJhR4iG
io8X0ApeXfnqxJe0e9xzAD8J71aPUOgvYb8fLaaS05dNOrvsI8Bi1z5tu5cKrZc5
+RaK//PPYC/0rQTrHbPof0Oi8OaydNA9XPHmIEsF5uBk+mgkSR9oJWgcCALiifkh
GpucN6G0XRsn7W+zTDRtd0kvp1oEXezRw+woMqVB3CHOUwFOaqlHOcqn+7Hs4cCz
iLcfvSUjI6eKtDYgmjGx2VqKjoTGNYCJGTVxodoxP0EFDAxjht6C08WUOJvpo5nb
UwNqbTPrIlWAtf87ncjVLW6kqnsbc6tDLUc0eZ/9k6ZmiWAyNCpegcVrKA7X2qV/
RLJ9dj327k/At54CBnF2akdgsstY9o8ClS5wszrn4Yn0yyfVt7mkG01nz1Ar/d1B
uNrN3wCBQMa34LgOh4jRqsCZuuuqrCx6o/ZFHtJiQAY3NF5vHzQcJOxSfdvaYhTD
NEHXKABoVnD8oGf+F9I58FDnwa7nzAN8NKdkov8VDmY9SBQRHpKqbe0GdvoBhA+P
jbM7NYAmnnAqMDl5G7R+yXCBtVCWSlRr/VNE58gH0xZXF6d1Bc3pPcytbutLPevo
0f6/pxojZsgaww+BjdgKafEalBzoInn9Q4Hy6i3NZqKGkTrrcOTgd22zH56OaSbW
+CmkWSYCbnIVtLfOtCAex/zS6SuP6Dq1U6h1GaCngH5vOkXdnZyntndQLh5SWQTb
CF0EBAF86awotpGHVP5M+1jqePjb9xA/buqSCXHOYtJ4EtW/e99R6R9qAz9rLWGb
2qyIsJ8oR8rQyi0AE7qFj9C80Gq9td0ELqpyHDTlwm+rg05rPVeSvdkYcn/V8C3m
JKs+tG8PWe+CcWyMM8LQyujIW+1j4cVdHkpLuuMItPofYo8bIPOTwgYzFEKDYPoT
XCj2Wo1ZHJqSW2L42wygInTqYzsTh0hsR/ZCgM/iuqaTyauZyD7+MsuLvB0sscCR
ZP4R6mP5zlhPby/sNKdzTZfLmhWIJdBVA1ZeY13F6WS/myG+7GOj48iqgrIDIQYY
T0b8arIwEFkLtmEZ92+/ibk60twbgLrfHK/gYqcI7z3U6JDNOmjp8m6hScsmf3wT
y/1fPmrdinPhnrUXp6ip7SpMpEty2HLUMRczfPxrtogMVnKRkkxGCppPP6t2Kfjh
ueTveM67mi1H/u6e66adOV+3dkdx96ncAm/yJBf1PccztJX6iSZbOBRY0hL4ablS
eHkN56zl3UyRiD5ZjW2pZ61e+iTI1HYCVxxRjVWpZQ2VGbr9Gjo40pRcbXjHmWr4
nDST02BTIAVVTSJWntDOl6zZ+gYmVBAQyX0fnP1ucDjtiwFuikHl8ToktiLvs1N7
2kAVbbYQg6/t0oXdaKn65ULmREo57pirL0LPUSA2hKcIFNekwnadXDF5XfYI2Gcf
qQ/8qToiZIXTieaMajJZATIgJTCTCXlCGpk6TyV8hhOJf5U1b/gZ/+MWB63lrVHR
niejUmn72osiT4NfW7zQZnEXsoyhB/RQwUaMl7yuQ3xKIWuxaIGWwqHa/DWh7gc9
PhlkGiZFAdrKOteiaRYa6Rsa8IQKEQWwoGW+7pSryZaBBMfScaa0iVtToLrvRoP2
+xG4U4HDI3wPyOMkoM1xLxWKGjqmVveP0xGAYPOz+ODPI66OudoCjQunZ6LMEBih
YCM1+nzcqHWIA19t7Pn6JCgK8IYZWUP8dv1arhn8bq3fZv8D54vYcZzwqHHjdcz2
lEcl2H4bRTFgC3NrxJwHbYk/7FYnJd32/XGG6tZK/oZyN2/uJ+MUg5Tc5nYMpoGu
VIOOvIUqApEmRVSidjrGP0Nopy0uTjqkxxhVv2xzWYORdSM3ODZCC5t+/7C9JZ88
HT6azMLf6fJETR8Xf3ItH9tlT5B64qBAHC6emP3dd4R3FiKHKN+yxKuqms1QFvWC
wbaaPDrWtPCmI2vIJK6PSDAz04xHquUbyozn/wnXU+q66HAP6cIGV7mWT0pKFKOP
sxzyJULyD8EbHpeGSPmHRyYwNZakopWsPCQpa0JKGDYGCmC9ug8iEUWmMhkKkpC8
2zMlPbDl7Q2gJXoKYBq6MeV+zhKonbun7PKUys8o4QMS96W/l2mdqv8AdCoNbEXE
SmgcvBytVaeiz0AaZfn3tKYsAaWap9NKqjTmu9TjfXx2s9+OjTWO8E8lZtEmObvs
iLoCOcAGOy0SP6fCM4Fv3F3eJZO8Kb3PvAWVA9WARV78E4dU4nl0iWPnDlrojRPU
CdveM9H3R89wuO4S2odxl10p2nzAUJI5KMA0QNbXnhuvceRZaq2E3b6boO29wsT0
O7fnER0saNGWsNn7RCgL5XwzoW/WajPiEo5jAwDZxJLyJ28oFrwYZryVJlsO/Klr
16pYglm42pAUdUBQbTZQyDYGg56qAlS7YcnIUAxsBaHwXsRy4mdv9BpdKBqH6fSA
btVQ5i3aJwN20nOxJjai9Yvnp9ueTq0/XfojSWd/qbUU5SzRzelalq3gZwplWD3n
Rt7MIf8LI+NXUvHG6a0bHnmufWcFkFM+uLP+eV8RfClqWj4G6IJiybCKREDi8tVe
53LUFBXVVRwoLv6lULkG8PW8i7/4QX6Uf0QBSZi/gBZ33br7pljAnMI1uzv6VHez
b+dwBI/KXY8M278WABvBRkpkGwuXUmuwZqd+/HGaWFOR+3Ge0wt1IHK1C7UCVUI3
QbeyHdwxPuzruzaiyMFAvTygD/Ps63OoDZCfUoyJuc0NUN87LQLnyiFTe7Whv5JB
WXq++29+/BY56XuJr5u8dOQKTEfdl/DUHlW4E0RuFVASMNOJ5p8LE0b7yrQP62u2
IAY7dAU7Ns9V680yDIfyrclXrHnhtqTLrHV63NoNjpTbV537inqLu1tjyKFgZ5L4
giyUUwHImg288is6F2Ofh/NnFf8uxYW3L2jT7AKuRYLkioFquvAnT9sfU/YSmuvw
MxgI5rFUpGB/y4S+p6Ai2tvRJf9nKVB8I2Vz1SdulW52Z0PdWOQNgg4QtqidbvkF
5NTrnzyx0n3adMgxaYjTrAA8xCaJw7Zi9ngiELr65KNPjlBhARfWdGdkiP0AjIEW
EVzrwyIjfplh2X9zE/KLgzWJ9rEDfu2fq68EPmaDCZYo6gDrjkiJHnOkI9VZF6Kw
HraI/FO57Rv1ljkt3kg4214dI5ZjaB0KkeBBmajQNTOTRnbBHRb95P1OGHUKx7iX
w3IklcKHec8/wEbSkCc2c9zZGZvojzvmBRMYAjLBCA88tSzJSaYxe8D7793GmWEN
FXGWACpo0jisFH06mNcWi0TPJFUw6IMZHgRWpBrSkh/HKI+I0MGEXnWs78/qxfPc
IwY1ayrRNFN8XR22FaEpijudCjAyTwqOpDsw/I6LHahccyhwGJ2+N3JJA5UKCFNd
HxD6Knf9P35Rn43lA8V2oIqGUzI8EV5CHc3EHG0FdXrASVnzp7kX1ix8GVfizFaH
ITZYvNnHTW5l70RHCdYjrxBe3gDfnutaVsVgsmnGVfAy6FcVeeglLVVGzoXJ9nhk
U2ZMb2vFPwu7JRUlWN8CQ5FhYXiioXggJnwLS74WQpQFJ3ZjKD8MYu0+E3fVoXD6
9Ib4ROM4nYS8a1N8/pEjDfjhhohdRz1LEMzJP7q0wfTsBh42Fd/L/cgnuZXpvXGT
VwShqsU85qh4MKn2o96Clj5gm2OsVxEbjStOlRgUhY2S2/aAAi57JrqqyIE/zQNh
mcHZF7yRQCtbFCoJyTN7YZyclS2mExS5wtuYqwCjTXTSjtKUyrYXKm+aLGPGMHfh
UjtRrwM6UuZ2pMHJ10Gf4ii68P/rfFTDE65ZHEdIwWQ2BD47XdXVjxZR1o+3JrEn
4OuyQgjFBcjSv16b4K7mRo/AZxS9ceNLtR2SMIPouvb92Q4Ktd044w9EZsM0wvcO
mgorAUoHxHoDJCMnwNo4Is/WcilnQMEAbExZkahNLmjqxPY0vJX4U6SmWO1jmmf5
c3YgiiuyXx+UYwK4t0YmooQ22TvZCLkbZrR8v43cPxWnIdB2v46GOpnFnkBJDPCG
F9df1Ea/+imig91bes7qNHODli9FlQMWstqeS+PCmqz8F7KFLp/DDJX76uymTV+j
RqqOPovntnTuLopojEmTyjHI6mM5vHhtqwuR1wzteS9PqpAkJojk3PoMvWDDRRsG
AqEy8LO63k6VNA+xwqRa+X/3cZMrJQJurm1Z8bxvOP5AxqnsPndJh2eNvnJOK2XU
DCaUpCBRONlYj9gtPc/s82MsSOb4xY/uYvTUowvrLqNEZjlfDBHG0Cno5EkGqptK
maslanJwvbSilFjHhpF8xtfYeB8Id/Cc/c+53tGNE75/1wKiSsgY0EJL/v4rRg5I
0e4IFSToN9m72hsybbvHZ8yyK/AEqC3Mo6F799DtLdeDIp0BxqcpiMOWvYp/Pk8G
GKDdID7acmNHqpOgRzq7eTOWmFTP7PDHVa3hFQhXL/GvrNCaQJxFpbSXLJmEJVXB
8iPRo9DiCsjlke0LL++gArLTVuT7fT2dmkYWSu8NV2YlZhXYTMNCUBe+w61lhZfd
BqNyI2ViRMn0v3bfAEosQSZPGVvhSU5CWJtQaafpGZtORbZHO6ojFS1F+ff45Qvf
8Kn9nKoZL+uMjFprjxQceTwnFGJKCzrZlmAFo9Nf9vcgzQKp7f+PcwKA+zw7aIjB
Relr0VVzXg2UQuhTM5+gs3t5Q7NjK7JYI6kKfX4nDDp0usXikDw267WFb+LpWugZ
a6xvWmicVqvM2fd2ELmcypzXXQB6OuTXMMNejYbFtTyN/Axb7HU81BdRdqUxyv4v
/4k2X/bFkKSJxKZIGMmCNWDDnDi58fRVORoU9v3fZ3PZIPSb4YZYETNSZ9MvUoNj
nCwO2s/FW+uxHib4rRPOoyqm3UlpVbSHEaBjVkTGSqoaL1zWeRhN6jCWeUx3kFai
NkuxAFibRuK0dYhgG2aFFnt+SOkZhx4ii5h78HYVJsnTePWw3oWdqvfQcmX8pKAN
ZBiMZ13vQv/7aQyt7+G/iBRoyoBHXvwO/M9SJbladmQg9lLLakJWt2FdUTbwAFkI
jAh4DEJCl8bFg6wDlKNmFoJdn0WND+EN5S2TwHfq4ycRAaetphK11CXAS8P/X0zx
00MdHaw94k/hdoyuIeHlREJQWIsBGGX48oIsRD5a1K91cliLV/sml4kzEqmO5IGt
eE+0UJ8qZtzu2vvxCYsWUDXLhIZSLqXPlOMbRyDzdZrWUJPJ0R2IXesyfvMJxyaE
YE8L3eFeDF1V3eCIbzEAvYqwoK0YKWhgyaQU+/jXtawLfiqS9pSgA3DJ0w2RrPcm
k0qQrfV0AZwg0OYbRfUzjT8TSl1P+yODg24Qp1R2Ll4Y/qyjWfhhzE967mU1tMzy
ChU2OPNccno4LUhNuvRsEDWvPePyUiiwV/1vJ0472ZFh3qs+dEvaHm1hPvJxpjeq
xyxJWMh4c6yhj8TpTNLX2NP62B25XJP7bSFGbvKU7gUJPoeowNnynbH1UZkEH/Ws
s3+k/5fVn2PJwS/4axaBzDrHKJV7O4+Yu76DgtQcaIfdiSJOD3I3lFgzYo23j2F3
zfmVfvp1epSVe98ACOoQaRhGyJF8BdyC+ZHmuLL1W6FCjYwSp3jstkwC+xsa5RZT
1ASl4CoQieyuyPEw/lltIE018fH9cwkNOkZGlyaMgBG/fvC/h4Q+qy9mBUB1OruI
cDs9nNt5lolo+rtzhrCpQRv5aliOZW3WLcNImlFj75HC0Wqb3DuHJOinFzBIcl8G
AjQWkjVb3WdfjJA/Ij0SSPE08UFcVTGNyW/r7ulb6ia1b18F0JPw9S4mfkU1Wp++
PtODlL1IteHjP4DzFyA2QiAy6I9xxBdIX3jQ8Cn1tFdF6A9i407e94kiEjhXe896
Xhfn0GIAzI8flHwipyeQHdpG39+I1HtgApZyfWPtg/73Zb60Y+dQpRhJJ+G3qwUs
C3ph8V2AJOSWKTu5fEh7VLMTFRmF6UXJJyStqtHxQXDDKGAOR95QRvmLeYkHT2Mq
EbP3MW5Z73moooilijyimPq7BakIqZOLzEIqTlNZRwO+ugN4F//109lQLokVA6kw
fE8sZ2QTHS+8DmSwVuD0UNi3+vdIxs57SKW0UwOIrlhT5nyoDJ0w5Zg7OfJXrWQp
sHEdDvtgqfW+MzSeco+Z/hl7uh8UnOQOHh08sLiAu5gaNBSFoLWQ7SBc0o4LfElc
2t3/tknTaV8spp+ifXnFWNc3Zl8vy4FrT7+B5GM+3q+vOnoFt/TmdkNq8ySoTQda
Kl6pqd1+kbdZJnWNgdIQxNLis0P4NWBAmlDGu7CAAm7/f/MtSm96IO9Kpbx7ci7i
RykuvKDxRUIIDgQYfb6Z5olNAcL7+qLoK4If1y1ocsZhv3Mr7j3dQN4nzOiqBPEB
f1BvmitOaoXmXHwEB6LFojoVNLBoaEoAbQ+IK9y2ILDsWPTa+B5IzOttR2bxCrGc
muy3/l0ZBixTGnmrW92x6rSo00GWhmb0oCQboqPyWUWRzKpu4FrXsRYBP7BfcQVp
YKNGVx4BoAb/QFHoqX2kEcnLrLYVhPdEldKW9Qcw/lfeQXWyiYmOb8o3b0RnmdQ4
iif1WCVwynnUrTBQZygg1Hh01cTjWfXECiQHBKnWWMtMbGp2RORwtEIRRI3esiQt
kMmQUVHJXy/gm7ZxfJ308wmXF9hVkNbNIMvieCR9JFgAYYtDJXQt5Ns0HSx/+YcB
Vs7dTsqnwvQ4sClNYALR87Gqgfr1Dt6OtyQFL0LOd7QUo8H4r+Ba4Avxns8eMEWA
edBwd6MVSQxOG32Wd//q//RU5vvLz1LH4vi/7NyCpSFKrA2SJBqLiq42rNCcOqh/
AR8zWJ/VNkYpN1ezc9PmAMrCQjrQu14UovAjDnyrXx8+W4NqZy16p0mtBAo5cbB2
XO9XCJE3OJDHodjpdzstJeomibaMBjI/roVCRqdsTI/7qygox0E9yZoQfVzwOMPy
rJLcOy2fdVzquYlb8TAfHWl6V22mWcexcfyp5n5pDkJLnMVqo6DcCz+q1J7kjZBi
sWw4VIc3uhVORjJUVO11A6+VpI5bKWQRA/oPGuWtH7wetS3hUq9NcXkg1O3hSAUD
mEHVyGyVfamVKmMTuCTCiViZxSiCwwEwC/HahriH5CjBYWbJuHKgJLRNFMU+tde9
6jo+LC1n6RR3Lh/ctHOJ4TyQYIexqTJnbJ74juI5ST1ajedX8H6cQWPqTEnDAjp4
Oq0rXj8fJfk/4m7zIHo6Gq8TMt0yzP/cLRHeXHKHn/Gw8iDn2qUqdtVV9YY4Po3r
kpzoYrvhTLF90xml3Aj3fO3nGQHGohuzWU9Z9SziW9Rb4QkNoiJR74qVh4gx2CDW
3GzsXSg4+JYNKjyosFqjbOcllftzIict8J61ap6kmb8n83P3zfhfaoNDJYaA2V6C
JswQPAhsPnluFnIW9glvOaI1VgIxPdMsoLJEQkk+dqHPhOF/cqWQmBXs/STHDMAl
/vT0ydoWousqIKaC7y6xD84QOLMfHoInDpugUZH7kaIbytjn8/9ppOAPI3vnSvK7
NzzrIvizNVB0zmWQ4SHvu3+HtCMm4nJiqyGpoHM3sD5d2o9R7aJSOXfCf+wHrf3t
0jHSI11TH9FH7oNZbqNYCN94T8d3GJxkYshnqZ0UIwx5JiXDJLKt1cRR43SIAg/g
bWiQedWxA8MXuGZC7Q3wqDiOuk2Fho/TRma8YNu4gSA/JGR0/tfVyNAo13TKdQ51
o3BhirkIPglWfsWDqU1WV2ZfSkkjN+2NWiI4QchjOrOQFHSMInhy8yGXCHInOwgE
xQBgMmoJ9y5JnbMourszX3/ZRbOM3VSzQVdiRmq4lVz0NCRSDtMA6Sri7rm+HhXK
Q2jqQ0VKtRAPITEhJuW3ffmsdYqthp84eUDCZs4upEm9gw7IvYOgwXR/5oxH/dQM
LlxH3kBtL1bkdiiEMeb1UVl9vwXQSpdWIJMtbktIm7ud9XGnSFTkabstO5jgYbIq
pNICXNerGrkxAU3s5i2C3Oatu1s92/z0XwgbBsX7Z6sU7z1ayh6xqyQqTLaJCTqI
7A2g+iicnD7maRIsm+3rHCk6rdFp+XbWzbo83rUWJkqwC8p7ttBNJ0FCVxzjoG2M
s6C+IlWF+gqUFymCJb+J8oCDltcFkm5czUNYiKXpgF+c+UWcq9p+AiVAn9w3mB2U
5aOKX8bOeLqnUUNfNBS+s4p+rAa1eNPX6pQYVkxZgM/Q+r2kDHKf+uOTdYcvx0iz
xRUAqntmCH5GXyjDDObd/sFvkPS7sDzZ4NtN3em7SI1mGhI3xSfzRKaAcWfonEZ+
WNMcc13LDxK16asT90hciVqDi9IHW2Wl6C5fcIQeKZ9p+ATK32K7IMszJa50/gKp
MBc0gBd719EIemdgr68yfAwgmv6q6aRqQmUtj+yJHg5UxionwJ71jx9W+TmcYK+3
ANu7uLb65v7hUeh0b87MHiN17uv6bekxMKL8SnUwM0T0FovJ4c0GQa/4R3o0keMy
P1u79DtrzoJhNMQnnijLc9AoD5toLC5/rfZxsD8LHXrmlgvYbl6I9jWq9TpY3JfA
a5MZKgTwrdTcGh6vomgzsVRlVizqaUDKH1nLt9eDttKZujniYcu/ouS6ZOHdb4Mi
YTPVd75ONgSsciTHWza3DmbJW4JsoB62Z6agChZfA8XK4IOykPm2h5HoyiHXpMo+
Q6qOkA1uezQ6ESh2xp9XdSwfNE6n8t9GKmUTGMOWUp5p1caRyIOenMjXvguIstls
V6WBgQPZvizJyca4QUBhsZ4taFGFOKnDVxjudR97iFjshTsgo+3q3RSWxnAoKqQt
g42PU+CBDjwV5wItJXYlPgSk9xAb5wbxzN+FU4sb47MEo7U2rY4nPot/vEUA9Cf3
GUnxZg8VkPfipzWLnZvIuQDUpBGtbxrL8qKUGvXCnCSttW9n6mrWLGSQNb7Kuptv
kuNbjX9JBL+nDuBzsXGUJKiZAV5nQY5o8Oj3INNJYTzPoQU2O8CKdQQqZmZegBmB
t6aJOh2zIcBQ0kZoI4TavhVvqNzVxirYpMr8/WlZcHfpROI4yOFN86lz/LEIHJLz
2WZWOkVCyPbPPhpAE+KXxlcIb2eQjCs++gfvRxXwv6gqvcZKW03odMqt8286EP7U
pauVjiaArHNQzcA8VlP6dxBxkqN+Ox+XzwCH744ufwDEASLa4PNKwwXv4YoLCUWZ
Ci/uzXBnPkvWLcOL7NaA4S/bhumn3pIzt4vI9eGON08tqx0pry+gLKanvh3O+8ak
/8jbaz5GJ9Orz6kD7YGeucMiCgyMyIh5hF5RDNy6tvcWULl2Dzlo8R8CZ/DVgrJ3
NS9Oy1av/Czj4Ydi5Zs03dLWFvV/6RVBzRFMcfC+iyWkQlGiR/ITBpEYVHrNmYgT
An4vkv/KoufxQc6mlSA6o7/4AoxY3Wm6PVTEK6GQ4xgRdFWpNG1UK6hSYFSJCNeU
JMhQ10t1G+iY2JTHTgroOl3N9/TO76O6axNhPIH7rOm30Ikk4cCUiQJrOt40oRht
x7xlQUkZlYIHuRk4mwNGLhDKwfAHC7zwui1xfuGvzPSxD8j89L8BLrhMNEiFxsAn
C8OCYuzvBr/ASxShW/AX0ivyyljev9sOH64K+n0sc2svqH4jHkihejxORkyTXqdk
jC0IrgV1PUeFWKsltXw0dLDpNkEdotRUOG3OF2g8Lj9+s7FWPdJ+fnfjrZTEA8Pa
5GEtyKq9lV+G7A3s3DC+L9jdiBz982ECTKN2g9iCnmReMmYH/m4vr0O39rxDok+v
MH97B4neoNqMr9CrBKPNuyKwhJI9uVy0O1cgtFIGtAhHDos+ZEiQdOoUS26XT3Iu
BT2Wkw/7AbZAZHNDkEnGTwiZdpuRw85zI35+xGywrk9GG7EcKh8liaYL2Kgcr7qE
n6yLZdKPJgcmwHF+4HqXBxbm0jJ0VremnHpChs7JWA0KvCN3/YrDwT16IzuYrLuQ
FzJA9t3F+HIsMwCT1hGvIQ1BHGLPNM6+P4oG+cPGpsKCn9q/CIUDrJYJ0PJJCRJ3
seGUQ6A2Y9pppWI7NTtYbkIXopTGldzAf1OoLrhyvorDKQpZRZlAtxomEdy5xy3A
YdJ0SZlHlZLOUnTlc1jmnBZTCVxVBCFjZrSKnBSI0Iaj3svLX3U1LswW96xrQXQR
s8IQWk/oEJ29WEYit7bKbOiOut6dh3qwNiWaJkKyykFFRa5G/3vgtd5oyLji1QpE
UKuOTydw9b5mFaWiOOhHzYCjZQcGoURS8AVYQKq/qQaSk/huQ79F5FBscVH5Pr5g
y8P1k7IFetfp7ScSxnyXMHERcsDaSnMSl9X+bazV+17HpCPq5dtqu9PFYNPcIwCB
av236xQbwAnURtpr35fZpKWVatk0RTLT5pHUhRQKek/T8bbE4+8yBr+B5Rr8CnfO
001gtLfhadnCVESFMEEpkWW5G5lCAnNwqnZOgGjP0gMeoFw+dchhxV4nRaqHfmfS
RW8ynVh9wgDzaVCX5et5ilPAyYoD+6//jr20972MAk94BoNydt5QkoGQKA1WnMHv
YWGAvYEhmSro3SNFBLIJBtiHIRpj1PA8MQT80VvMqx7UBnsGTZtvjV+EWc5tq7TP
tMR0aAzrDaZq20eMxtFJoJPrqL4MsnszH0uC1mEZ0nHsY3QEZmI8bOrJVUIrZCsJ
TAjA8GzMRSrGMrpqR8YxgD6ish19vVG0WgjI3IH33MRO7gqvv3gfVAhoRCsbzA3K
YrWvDiFH2R2WlQHmSJT/6a7XK8un68kM/zvD4gEY5CbucU85yaevEVO41mlUIxIe
pnHyS2mZCsmlMBdv3lZChF1AsPMH36rXtCiBWR7x/yJ6HM6JGds0KCvnEIvDeAJY
lcxUWrHmYjdvfaNgFkReWHnC94U0ff9RYSAm1YeNSJSA7K3Rr4XFcE0ZRH4+E5V/
btJRRPv9JgmPigsb1V3fMhDEffR2ISo/GKaWBmXDPpVWNe5ZsiHxPW7y1AWhfzkb
OV5r2wMGCEfW8BUgSgBRpNr9G5UfvMlCyTRQxoxt60/8mnZGsr0DIHg5chs+ATPK
SeFfQ3JH5ce+64bzF4NIyuvpwKrYasfq+wSP+CixblAVuETRU/7XgIUxOakkCeEJ
UHOC6NtSjcwmU7Hn4Q60GWcjKbJO6aIvUfYzYNjiGhq4ngexSNe/Vh5YAZxV195a
4K6hC7n0bjSXEJRIckVUL4GgWh3OfFpQhShn9CmLaqarvNjyDVLP8yO+Y0oPL8hH
FZrtpyBDe9qVEs155ieVCopamScAlsNdaiHtg5ZDBtySD0zyYmWQ9sv1YQEgmu6A
NeOUgEr7p4Irzsw1RM+aB3uCLndhKCWFA1MyaXInNXzcwBmnzyzFkFrL16jnjCql
943tlviMXPsEgQUrTZvFCNHd9ovLXNjyDseje3P/w3zoQ5mQClGw7NC5JqoLGZYr
guDyu8CjqhKPd9udwychRCswQ5R73BR30EF5Zx0MB6qJTwRmIB8Eg5fuoNTbF4sU
IKtOFVFuEjdsaBoOZcLePYkdaEO0NzoHOYnVnKZ+Noc/7duhwA+qJYNe2b2VlWlr
Lz/NJtZ/yR+fmTiNjzaGLEhGHmp3d7P/hE5L/F9LI5wRjqNUklD5Qywl+Em08JPL
J8Qauz8Zl+Lh+abAhlE8f2pK/JCB7cl/VlxOWKX8/R0K0Nuju1kRd9isksN4DHuT
TJO1m0C6LYmfoWQd1GVrkFZwOOi57VDyhOg8DL5lRTjtza8CjbZUXfrwjlMuTdbJ
4JUIUrsR4c+mpjiKn5drktx+GzS2/3FWu5gLbf2E3of5KjnT2jDR34F8tdUNVbtL
vxHRlTAAxTomUAm19tiXxB0GGRrQXSGaQPa2s+deZ4YmLflTB16kBy+lRJPkcMTU
1viSf+E4XgjTDzhuMnTl8J/i5JjE+D6m4DE63Ezlq1kXMil9FTHLDadNpWq/PMCI
PbQim2FWkry8J8B0JuYwnXvyUE2zatvtKG6gRH+seglSoEEM+UD5lmHPfpmEuRpr
f9tZd+02JmmWrJJqgZQJ9uNE59O7pkaId8eIHqS+PFS7mc9qMxZeFha32ehvUw5D
+bM13vu0LVfePjClxzk1i3NZx2e15ke30eCRLbCGb3PR7ziL/ZvwxYLqyz//z6eu
G6fXUP1vibgq8XPliKOY7AAxRx2jDiH0jJaW/Xjks8WlnTz6v3l3cRRiCaWmBmtG
g95g/4GX2BDo+49sEaKKcbKmzO+xRW/kFiKL9pBQR3TR2aEarhGzTm6IUdV6iKnb
5TWW6gayxIK/4Qul5EEFmJqnibB3bMftm1uGHjwgoGArnSboIIjLL1WMT4xNvwPC
WXKTPEuHC2/3myys6Z71PdYUgWE08AsgBZiUkIChrmx38tGiqvsaJ+XSz1zKTbmh
B12gmjdlWWQosO+hCpPLg9wcVXvGKzOUqLGEb72puGTdJwUiucmG0FE5c+SBAHEH
k4yh7EQZH1PvAi9NW5E7sHUnd4ZMiZZhyAILKH9YMsf9KXqGz9z6JuBQzR5Nv05/
eIng0hMlfbK3+rEwqKC0ZuKXjuMnO1R9pnptO9ThX4MYKr+XGEF+63HQmDN9tuha
2/y11Aq1ZVi/DBpoxjVu2LrNqZLDNXFDnknIGzstrd6esie3koWwYiq4W0MT59mY
QwAKQmIc4JAa0tLEOiRDe4h+sJZWaocZ2+EPyN34BUcxh1eUbKt9q2D8z2hKChZ6
jIRsKVA6wkNXBWd89o6Lc64+0DZkVguZ2vzIVRPXFGdDDaHnpOs1RKx97dOkqqcW
3GwZ9JhbQjiNdpFb8MekU9/EUIj/BEjyJh68AZzA7f7IACQ87zSOgJA44gxT8TPn
SF86nnUo5urYnprGWubjKxkaZsxMkFXwEfiDdeR3ssOT3mb/WfSFcy9cLFF9+856
1LQQ62B9ZFvwMo7fWHhD0khisvhQ6uHB5eglbFZGU0PagmfuAOfvRO5RyKf2yDn1
vUcJNKUkXz3RrvScqOQql8aCzbSjq5q2PxKnG17XB5q6bPP/0J+lRAsXRihie339
rGu8meLle81K/r/gd/BNisoxSiex0HxRRmVOKEZzvyT9+6ZU6XmAi2hOoykVZvYL
pMN9+LIw2SPKlohiKkJRgfqwkqjZtMbHHafPKrWpfWhdpV9rnyL0E0+UVZ21zbGe
rORCzbl6ZsAG4C5FYuScwyLXVQgHnUSrBNCWDMZ2R40WwrQSk0WLf4c0AJL7937u
RvtsGqcArqXE2bLFJ7/YwMZYJnhMeuBrJFSKygniy232mkyzuQICi5S3HQ2TE3bI
BT0zQogV7oa31Sd88hP4q7bGEJDMY1+qdkkGmjsVbl9JdYXV/eN4JTTEt93v/x7Y
96nhK5c6pFBknTAt4p47HkaUCjseHB4WlNfZDc/5GHp4JPLPSd0PcTvkam8h5VpK
HCO9gKTabH6NjhwL5h37K1JKfiZr99vlgNXTYf3FHW4iTyR3AgS+txt2olxJN/Lg
AVAioOj4EAiQgN1Ql2r3ubyP/NhwNkq8ODFuWmdiH94kfhFa6oX3NSxBMxYUw8+K
ap72M5pypE8xtGgBQUCbGcQZ5jhCBpBgknY8hs5U4I/LoJexw6i3Cq554mWUDxSS
b+HO6I/9xISE5AR9BrrkpaSGXfK0Uoycx4q6vgaDE6DXI26RR5J9bp+P0BURszCo
/Z2DoIhFRUUO2uO95J8a7gnGyK7cCyFRSz+Ye5ZkEv4gEo2zfhPvN7QBmlEDwopb
ZRI9DNMMv4A7cE+u/BRe4YtvbWovEYrtDLw0au1JvUFJqqyS4O1x1qzKr3TnYYNT
G2Ne2H4S8qO0lFpKY3uRK1shCczJXYCOaH6wLuIBKEa/GydM8WERF3Wdl3xxdjtY
dbkpwwH3hV0gwFU5vNrUvpqjB3Gc7AnryIxzGIes3W/t86NLC6ItY+Nn0Kf8ypwc
e98inzZHaD7zQ2JbUYzHQq5U41nPg2+cdJEn5ntDNRMGv38ji2+ssBkgTc9OOrDp
5ewzT7FTZRaNYWdr3kQ1ox0fCwQcUIt4D6Fx3SwYv1CT++XRwyH/H8C5SFDSmJeY
Nqn0lvwbFK+Ps1KKD/PZWC3tjCkietge8vlpWSpM/vICjQ3fBPJF2/L60dR2gGHs
8FprDv55Q7aHpi2XqQcqDnE7WdP90cdkxkxottEQ/omw5ADdw3BIy0nR83OHtRPH
sQnmIRRzPBdR5Za76cAA/UipX+CKGjtASq9AvjPF9Z7BsJqnnN0BTnF7XfRZHL+8
7xhMiWEzslchCdPhNKNZ5vNeKNV6Kb7x2mLkkGkawmHSNzM9pFuA6ThPCQDYoogv
wZ4O3Sxc5gaHRE44mxSam2uehJC/Xvj8sAhrskYTGJufSl3kAsIRqcZeNFth+18k
icHc/5BGg91Ek3JkzEfUbNVHLNaWtaAd+kDsTNdAFNdQh/RiuyrTcO2wt7Fp6o2g
sMit423asta7v1uu3SkOBa0+q6PK54WL7rCTXGNbi0hm6NjEohBnqKZerRiWTY76
COSsdNISJXpo3RXKJXF8tahFl4YTH9mgrBqizXc9lVags9jmcgMtAkHTIST98bPV
fdRQKJudd+aARF1c73jFylycxrZ7Mw1SCKd+W3dhMmLOlzoI2Ydtchij+TcEiFzp
T2+4MqQ06YWPcvUfkKk46Q4pxCbJCRGWnzQ5vokEx8NjoIxN0FRD6YuPqEbUrTVg
Fdl36moxMZgZ3NjOO+oB/oC2gZM2qHk8kF+ryV5saP04oCU88ESp2DRuBuHAVOov
U5j7ASKQjb3SzFNuTQ755/EowgbJoo7RgsNQwCG90ZRXuYR0oW/IjqcyHW7L/v3V
XpRzuqtyw5HNYPNcQ+0gzNZlzviCB9UsIinSnGXahqOJZFX2Qz6+2FGx9G+xCR/x
uxBbn9+QC8bxKipO93O8yM2camQLTEKKBZbztUwc2pn/n4dy7Ht0jNkqy8TN8o5v
zRGlm7RzcuqngIyv1l2Pd2HYYxP3iqaUPMtDP6gFS+mn2q43Gl+ZXVY9hjtIFkjw
tJI6WiVEhvQfI1XnAddpQttoCy7kZnxMEcNwZeS47Q+gri7teEM3X5TjTOI+HH+2
lilYVD9n4vl5g5/TSUTPSWGLNzC9E1wFTlS6MOF6XeuwG9fHnmU8nTAcxucYOwcW
LMMY7xhYEGqrTIpdqnQm3yxXuqBFqHbKgZDerJk0JdN7NlTVlFVMWVMzfKmWmkq7
BUQYFeWzWcAFMQZ3AKrX6JAb4+T8qpMPws9X+10BW80+DfjKxp/aMC6R2DhbXMYv
5cVRHxP7yEZtSSeKMjNhD+3VnXLbtovUkW0wj/uspZAyXSp2+RfJrrzvKBDWJbit
GqZ6Y6I3DF3bxJuoKMDDjAu/JONNoqmqeDXHwHkHo0Tq2lIMAD+bq8JELQQJuhHr
BN1Lji3oMMDHklOIE/RuJ8JU6XDAznCfF69u0MHbXD1fbrR8PWVabvmvtFEGz02q
icQXE/ZdKdS0u+7ianeJtBdGE+gW4tdlbYukkfc4ue55T3S64LQVh21RW7k8TDey
6lQ8qeRLt+PpuCRo10aHiz6DF/W9PTLIu0Cl7cxzHifn+PwL9VrnULH/X0hisCFE
HECYmzhlsqjh8UIL6POYZotxWLVXTrPsr9s0CXjp1zC93gpyffe732yJUx2kdkKF
HD6R08YjnySugfUy0askmhFsQM7kJx7CHN+VdWLXbwoK+GEnqCzqZ/dOFusxWW4w
3nMdu4mijF/EYFOfKHRF10D9GzR7lDd451Ajr+3phYun5Fue3Yoeu3hfP3onlJ84
jiiPWLfki8eYVKffWt4bG85TagNfZWYp8Q5Tt3ArbAUq6Vx6U3hL4IXsbF6jxcKo
GXhj5K2rdJQ92q4P9fzIRQzJXPRhwGGYXSacpmjTRWIjh02wfGFdLLDGQkt64aB/
wppMumGhQ20AvxoGDoxoP13aENfcqp8kXSIauQieKROfXlU3kYMH30Qh3R00QRgX
Q6RC97qrZkIjn+Pj3zyOtaXVUTxXM1QjbbUqyS4jbXEJdB5dPr/ifh3kE5M0CBJ5
PGPCv7ftbH1RBBnPctMowjS+xNo+luhaJaX8vhvUV6OmgQJDLry5pI+aKd4pBQQp
1IuLr8e3fhVaCJXFJRcTuf3cFDhSH4O4SKhncf0fDEJ2hfQsAVRap0yeRzw/GINz
n5DBYyNShr2TcF30256TuNISPgKZLq039DjIwpWQjJ0DKIpx4Jw9Mg963iukPYst
chN8ze+4Ao7QYeg+7t3K/eYvo81p1GgvpxZhmiFcR6Jgu/Dhtk9mVKgkL4+LRoMI
MN+BMIBMCcdMjgIdT3+UfCRoMnUU5G6uVsA8PR7KSJmdar8dFxNK33B7MKUowtj8
uXLh5uH/0Cl2QuKjevgOT81DMd48ltNjvcsOXsr3qTIlHtB3CW4V38HFHsO40XAM
tfb0+HJIuk51XkerfsYoHUaTG0YnYODY5alJMIvhpUIIVSUBFCGo26ivaFhuAqbh
7aw+S2gAf4hT9KIKKMf/4VPs6fXTteh7xVe42gMnbXiHcJfY2MZTU4Miul0d5CKL
gLhTBkc1mwgDhF7BFZwhm1yXN6QCjmQ8DUhaIhflJh0vNi0AUh9DzShRbRaaxFQw
3OlJdkS8Nw2OKEKzYiGHZO1+l/zk+3BcTDb1FfRtjSxMnnV/fx25Sill/aLD1TQd
dkyrW/eZBIflqKjfSetukHizSwfaDGscmqtxtIFWNc2f5g8yLvn2YT291d+lPPvq
kpAQtbIjifyUC0G/osJVOefOiQL4cus8dRx1xhF/hNYeaWK49BnTke39XPD5Fnhr
nxVgfev1FQuiLYifYSIJrBsTMUN5iRuWX+ilUbBYeLVIpqiNzK51wOCg2i9qWCjA
0HU1zVQgJba+snuioSV9HMKftVpCDI86ZAXnF7UJXr5dvZkT7ZcgSLEkNQHs60Lq
LjzO0lMNGZ9tC03WXVKjNqN6VR3hjEwSTkqSkEYdAp89Tj6Rjdpcqub3tz6s2fn6
Qh9vPjhwvcNxEblytxUHge66KOz4M43f4uz86pKFIuyNdLhaIg6CB+SDO2Sf9t9Y
kzY5LKBzqVIbCNxbZ6psaJKb2NhZ1IWx3pDENNDhnoKRIz+s3U7llW7hxwmeGv8q
SKrolLkgxumceTPtNd3wHBqahYbLymxKXLCKF2cNXdIsy5hcctlUGtM8dqgwtvqR
uU92m5x0IbGh/JyB/+szehniBCe+grsH/IChdoSOEbzf4RRLpRTIG7xJSHlWC5mm
27iOGf5DGMS9qu6S/pG+uELg6aYrUGyj3ovqXULEVVY+HfJtqOL7MKZL5o6XMBqk
2IIz9og5fskTnsqFjzogI4tlL5WEmRem54cvqNdHorb8s9/DDgRRWVRHnlRQYtSH
rMUrYu1wIQb8I4u5migghnjGumuoy9ThooojC7ZHotBFoXug6kdbwKREeaoOtMzN
ZgnmkslzOmBAtKIGhqoBWvIyrEnUFK+VmCeqtiJuH25A/0I60jGdN6ZkM8pQ1ZlJ
5zABleoCehZZ4gqYPaTPGG/asNr9q5dnLlxs2Lp2yYfz+0c9Sg42tLNBlTtIvZJm
dHpy63iyP+TWQ6e5mT46DLBxgiXPN6Z3XTbXDWq+8KpZAtM/AcMhfW9b0ZCVT1xK
bzU0kHzUfCAs5RzF6YXZ7jzV9ucv725un+VgyA4MbZwHFGiLcBqYzFXIL4ku3DFZ
NCie/X8ajko6nMHCO78EVVNOzA/yXXGVBnzMTIxVgFfBVuhclXSVM3G+5j8nia3E
bD6vDHFW4DUZ5DUNj51OKah4HfND4dSF7PH1doFUQEhs+Kzydpt8USd0MwAgwxCm
2eI+2+hVaZ2FFLTRiL2ykl4t1jxpVK1oWRGWzfdAy7rzSgZ3TlnYgXARzCu++b3t
23hZU+Vxi3yJz6XzcdiUBw1aAEBFFIf3Aj0AikXp5IjXW/x4q0kM/GvYxAehxVeP
61vpD5nhXKDQrmC9z6u9uijJwa0dF64QWOBIMXSc9YXeKQuq5bMVqtPbOimpbveg
vT0fxyy86HRXx4TeXS52cA7Z3ub2mQSoXs1zO+hoxsCbupTujhlUZFCuRAlcDV5t
OvrFr80L4zy/4YtjO5LNkgB/RccaLhHw8qDpB9BJgSAiLJW0EjoUIIpdOK3vmmtW
mc63WVkKTz0M8Y+SJ7gVGIhNgjph/pfykjyO9hu6Rw8mvcZbrRO0Y1D34rwgGajd
O1K30TMZdqMBgi4N7hdSgVj+fMEqBesAIXqt+1uJP4618Pta3UVLTOFIyBviV0m3
k1DKrVDa+qh693qWN4zcR2FBTRbEykYnIt1/F48KHhU1HxlKIrbjoKJvcOlnuvdc
3KKNZjFopgBGEvJOVtV8QgTNazzKmJnn1OrroUcMPWamEtLuaOGphCijIRuj1CD5
ZUQ11i3Z1AMRRgHnbqOm1MEmRQImwYR6pNa9GPCrmhUnOcF/tfqyMameRlpDbkF9
sqGLvtT2AcBY8iKYXOztlhd+lTQZAgCEQ3KumugHp8QXjxgtbgKnOwsJ8KEC3h7J
L7pVr9oyZJaczlHCvjo3lrSTICRfNKv0rKlatj70nNeubp+1FfaZH90Mt9ODDKh2
9PitLiKS4M+msCxSU2yv9QrmDiD8BZQ+JrXNuWVm6ZTleq7U7sjkWFMth3sOqBph
u8siXNYqkyp8ruiPij11lyKWucMDWh8/3Dsxs9QgDx28TGee1K2Lz26c+Fo9Mgna
un/FXShOsvwRG7b274RZ3P2MmLJWCwIrP7m5A3x8/VFxa3SSsWKaYa+u15xnPWYm
vr0kXr9Sur6XVjfhxUhnOs+5/LZnJ83VxK6u6we3LdXJeAvmhoYnMyP9aFtiPVnY
J4HFngi5ok/YWbaxpbH0OKX2rxCwqISLEYlC3xVgjsZDfYZj8A5ffDQk8oF3L59C
NtRyMFbyqRCWEtcOgUPWRfeTngQpe8CNE2XI7GcafB5nb2Pka9wnsgCQk2OqcYc2
jWypXitKT1HOylFp+T6+sR+cQ97msKie4Jo6ixc3nTeT9BEkZ93KFUlGnw0LWqVb
o1jpzW7Mh+1QWeBr7OzeMK/ltoYQS76GbmCUaOuVgMf4vmrmx0bfMNfys9RO+aj9
7pIYXRrbffKWvaFvTFLF+c/oVp0a0bE0UerxGTJa/Gty878rfHveiwvS6utDkR1o
Kt3DQ3jp8rNItpKfcCYm4AImq6Z8eTvula1I77c0enrwdeHl0D1bfc2SWwadwDu2
ORqtaaYY72Fg09lGVn4bQHwaopBsuvTyl4jPRX84rXOx7M59NlNsBx+LdH9Ujiea
XuX3IPGAl4/BFSN2cG9r5E8tM2MIr08L9ATLxj1z40k8qFiwgwH5YjXR3zIxUrPb
5sg4JZdngYc3VOeK1FRK8VRxNnMusECHsQoJSRf5FIi1iheKxDfPbQk2KRDLpxEz
DTHtGyAfzHLLQkhBLfEownlGjPHGKohXMOW4jwrTryYn6uOp/ZkyviSxg/Dfb+kE
wXkla4tUofEVJjZ6Za1hLQsZN29nPCLi4AHm8eaQoMt7Wk49tMzuR0j864VWitus
D4eroKcInCaH9U4zDntHnT2mAurZ7TuBukWFtEZ+aFM+a9bXBOZ/zyxy4laBckyq
UsdoNB8mQaGnM4UHZ+9Az/nKUd84dj6EfFjUdfVWaRaeXQBG7vPC9WWKVPYykAEH
Rw8uL0aU7srpTkivT42kIg78tn6hfGZDd7A8GPYmUa3msogkTn+m99DC+bkYxsSq
vuMxHsVbqXoGBkHgGm/I3uuulcCP3DAQe4avvo7C5rrj0ZtHv+xb4m0Rv0Fy715h
m9L0RYB5+fGkpzIdeOYUXoHcKEulCqCtdxo3+8HlsnG8Gm/uTAMNUPCrGSHnM8Sx
kjnUfFqspXtBtyrhU4F+XSfalyZ6P0EZ12QLd91aG1bKCKXdgT6Q0BNjPL+hO1Yv
7SwB+83cKW0vJz6Wca6dh4KUHWc6g8xtXM96pc2OQhmv/1S+6Uehps3G+hgYenfW
AbOk20z6xIQn/4TXsXlAZHYNZ+7AcZ2wxep1dWnlOpM7XfXVFF7LpOkFOfk5139D
wTVW31V68jz1CazbwsGwUk5kmBSvkfut8cYS9F2NMM3iC2HtExIEMUswP0iARF7C
jTiAHJPhFRcPeztyeiza9u1acikpHFRBTeDNbmJNkRDZYGZoPUQ772rQq8/b6DDe
Q2EbbXIdgHH6zDbHf1Z7O9sozcpknnfrT+PWwLcfbfoFS8XX5IMkQAzbxrXftdeb
zm0ABV10BPwCOJJ+mGsLfc6oz/OJq3T5M5dl9R2G+PTSXMMjMfP87rJP/azfTgYV
2EibSHzhtCTuammfpW6szYAGazG8rJAVivDQgqwvYmfIVZKBgANZ+8nI3w54f2Hl
GJcJfbTKqEroAjXndMPgGqaZLrmq3DfHnpLgf0hqXSRZm0Fyen0mqRozayaa8qzL
CVKFuEOgaw6oJtaAPo+6uSmOXKR49s7IVAzJWycCeAPKRK4bst3h3v3THhAki5In
lVo1TbtpPGJcELB9tm+Stt9EjZCp7qwGQCn6UX/I2bNwQMw//iEgUt6iw+/jPdTE
/5+6CIFtsjNI+95+yYo97vz4C8Y/ReQFpa0zhHgLeFYH3oAiIBzt7QBGl1uO61Mr
Lvmzx/3iVjroeSNz2SawZdk5Eb6fOa8KS0+0mklHMqqtyd9JArd810DQn0joyUY0
x0DB+RaPSufvPOLboalmZv29X4cHpAt1i94i8gucn+osXAc7COe8vh5YsJA9Dp97
bWFB8PL/Rzep5eUVXLWdTktPt/uYfozAnNxF6p7Ht7/5ggSuEdtPB2hvpwU0AvVS
fhoBJ+kqXax706kxcbw9YtATYwCcnonRCE92hkO/Kiw1k9kIUaZs/7834gXztlWg
OhjFBERRd4SmgMVH67c7+V/amye4/EhttyDHy079wgMVfTFycxvlGjY2eSPTaIEZ
d1PTG7FlbGGzhhCsGkWkksgfCVfULjy15bzxjrogJgO+KUkbJPC34n1V+kV1SiTW
mDo3v1MzAAsY+FS2iirHXdawHdT2UjQfiwjKA+VWx3zecE0nBS06cPI/IelmSXzx
fSUSRtjOr1U7ZdwNFmAhPB3bADsIP7Nq45/awxlZL0PtmDWmbCcNX/jqws4gTifQ
a7umrGM5iOtnOdzMPM+wQbWSLK3zzrI5YHSTzNsjacXgqmjJmevQD89RnfS0U5pu
Wm24BgkUDnmYtaqPfky+hD0Cv9cEgwq2KFm1LuVw9Jvd8NGuweRGFpIBjKSMShDJ
jPc2TpxbvV2iNffIbdMdibBQAiZYcT1Bh4YgO4zUztYFIWlVF+7O3MKRdpR7M5DT
iB7T4RSOIgaWr70CqcjcLZcU7gHzOAuT1mMggZI8KEGZurykNJUcIBW61wI0QIOa
EnHaI1+G4Y7SowEvLM8mMWt4SU97hrQ1FgHnrRzGsfrQdaPMcQa3+fuVkqJlzlEt
bnFb2372L8Qzwkc1J3KVXLUWYcJ1zfB8/M+CBoW1wriE7YujGX1woQXndurk0alE
no3S/dCfT6r8weQqA5RTGkQGUcv9+oWQDxG5DvK6iFysbVo/5hiXZcmjaqbUMdsV
M8cF3siNA4ZYCvwmlwCAV2HtRONlZc4P/FzgKTxJgeR1N/1QGS7ytrUDGRsiyFFj
MLjNG4xwJsYFyMiszBCgRhJgTbvrRFe0iB36XDNGwTOHaOwkugaKJwjn77+P3ZtC
qN3+s5hPzBNxsjNXSVZe7K8+NHG29w9KpQ3WaTTPAOAHw2QKS4N8C1JX9ab5IxPB
ftJNFDPJoUOyDV4cHRrcY7gw1yGOGXNo6QOzRaVjRNbj9kHlG1HvAQT/D7K42tnN
AIUVLxvDg0xkqE+UMNElOASwiewVU1FzAmzL7l/9f+D/C/tWAE0YBuRP79/vVtRx
R22lcZq1THXJqyt7wTwfF5f1Fgx+O/n7xbAf9ZxTLGGZhwNveieVK4Vb5hSnD6sH
EZrSvh4FQXGYmKFetedQ/PAJBQ19no2vZYT7XiyG/vLfq6de+D4ABd+RURLOQxDd
+W/fESaPyhlrK2jqP04QNXbtaCz3bVG6EBz7jDTC3Tx7BGOm4V4eqdZRdezvvw2l
F+DJ+EOOTrXwf0y48X0HVawiUSguoSDH0tlFWMciUzNq82pv/jlxScQIhl0RxHCz
5eAtsOX00L1GytnM6L8S5xrHewBwzBtZEiG5GB23z1MP/m3Y2soQsJeEbd7yOJWU
6aoGffYJtZHpsAMyFA2+1gyNjnfV0DC5gQZmejaQ5PBXoCJHHxdta6Le+gRAFMqf
o1BjdHXI56UlE9R9o6DvkbvAUw8yeuiRyPyh1wBrzbYdlk/O5oiqoEYgEp+e5AxM
UQniVjckpSgeRCQx+dClKpZGpq7eHLcKdNqzaa/RuGtkFexDnPbOz54KkgU8C5Zq
AB9iQejgUsUl8YU4DN8D7LICv4iso5I8me+0FvyhSjYv5VxGGeN5N067RLrQ9cSo
pE2rxCLUKPVCvACzWFrKlHkZuVjymOaUEKq4tm3Y2cPzZw5xLBoIOuTDSr8D5qry
NNPU1j5wTo+HyQyhUa5OK1Ixgs+g340Rco/b4YGjIfXxooRAJjOKPX0+Ne4DclBB
IANfb0BqIQyPe1IOnmxHBRYP6Mkudn952uhoWjNw11E1283fC/9H42QEeMbiLebv
CI4i2KQCaXJyeHgxmQiVOPO+9SN/DmDUdmVMWxBfWYjR0gpceIbGsMg2+yB/Jbaz
saymHSNpTsa7PxAhEtEA8GwJiDtsf7eHH9MKhrGnAOyUqcC1HZcZoFb6/n9TpE0i
8e2+ZumlgFG6CR+XEv+dPhILV5MyKwv0rmwrLdE2m43mok12NnTd6EpzpAwMpaYy
j++LkUywb+eCIfSXmUXqKckMMUuE1EXUjBlXG3Ng6bN71eOjYFPeG1b6DktO47Cx
ETzKzP05Cz2aHNuqJnpk2rw7UskSyohv//Oium0vks4rvg3ntR57bcsIlzkLf+Sh
g8QP82NyzHSE86FY++gpDyj+sz2B1S3dYOuTfCOuC0RIq+BxMcEMKO28N7RyDX58
4FEYBTIe9+U5muO/I41xPnz7OMQnYf9veq73Xoi3hrcUIv3Xq1vjv35ukNN9uxhW
jtl0iZ5uaQI354pNDDpUNS0Nvv9UfiKWmmaVQXKPN5+mSDe5sSAz4yC1sAQWEKNx
Yau7/mNO0LQTYHIfpD6cbFsaBcMwpG5d3+XSJMO5wj0T3yhVKhfd/4fELnKyfeP4
j15V1kwEAeNrXD38j2qxXt2lS8W6wKHyEB7lZyxa7G6hkDjbcRZDnM5FhChnHzh6
ktWdbSTEjpTqcxGm9C0Vcpe8kv8z18n5Dcdu0xsxOAFx7kujNUcvLCyFeMunPFTp
CEf6KOYfDkSMjo76Pr0PHaiw8QefPPpdyTZYtMNksl5Dga5U2lrPktdnDIQzJqUx
u+lcgmgA5zkpx2Z7J2LlVNgRCPkgye5MnGnG2DF3zXWq0vmEoWuOyfM6j41x2HdC
aAzsCFVsKZMQqjP9HKFKXPQxAdoV0fO+IgglynHwGBIG7UJ7vd3wMXhoe4Mtlc2m
YFT9SGa/M48M2l7y2bmgxJpwSO9sSXYPxLJY7snwLO9lJSvVhvM2v+gx3YJEBVGQ
51YwDQYcdL4rN7ixmT+4CdtQv+vofFJ476ZQFtfnVUZqrcnUw+ezf2SdEsiI4BHv
Jt8F5AOYlLWz0G0sLKFKztgX3hI4mDND46KbX09jCRpZTOgknC+RVcf9ExfjKgsz
Z/IyEdkW1RmZ85SkfSv4t3VIPvX7hUoceP531Tk6rR01YbraW7NRyceWfEjXYmyp
zRu8r1U27fSNnTyReFJ8sZ+pZWVuA6MjhbMLpJ4+67WFeH3mgOIUKOXQxJ/dKyZy
PHDjHzn2w1mTr512MAhRUP7HBKE1wiBZAYz3J1NBSjLTCqEJo2G1V/2tWxpwQ0st
td6BBNO6UF5S0uR3zAOECaTIi+IXxDaRFIwHhiG80lZ372GYmFAF+nd8ED7d54SD
2mp0paSmQikkgu+OSSV9BPz/bDAG9QqZYR2n/eH2fTumDFk9gtJE4A7y9bSTSFad
9kYKyuGMWeBFPIhv7b/u8FbnXYsPKTjo5KeblyWSajVLQgAPfz01BwyBGGNG8DRM
Sj5JCwPk23UpEClgXHx2vr8Qye3i9V3oY7KQVFEWxGCJyKVM1jpZrECBGGXjGyc/
zN4uiEhzUieVI5KZY4V/W9npokQTz42RTO94EgWPIbwTnp6AyCj3HYv42a2+XmTo
ainITXcx+zOc94GXyFwNI/wYL217J2jn2GxGZaRLWItVyH1UnhMaSDoimubqZr3f
lx4ey5EnSLahBeCDNOklesOCEV0mmV0okVt9s9g2jQwphcM0L5fH1WliNTob29wu
ohd2xYlYOHKeRn9D8ynFbTM97v/H9drvHOBVboFkmTRmkIVHO/KSBOH/rwW/CXlV
Gypu7WulIXkH62GA4ogNPy7CnPap396pliayIKedEH3LpIUX96Lv7PkZ58OS4xCX
NkwAiX+ZZrTD8OMSjN4GmcyG5hkyJsrVT6odFmiMr0kI1c/Nto8wmL73BBY4i3rd
ioJM7WOXVDBPxTCyhXznBCz9H8c8T8DRbxCSh3bItDpo9cCVzlCRfo50+FUB0y6u
Aayhr/WI734Ab8PMTAbSmdmPMudNRNMHbDmXaWcyenrYQgai4no6+mMW05zUv8ce
ko0VFdUVQqrvB4EdrvzeHZ5P0S4+cc/nb3fMSaW0iOzr3kxsHJFQ801KOKMmSIZ6
nd3y28Dr9YlCzH0CyKWcg8PO4Cfhyfpf5dysPyJgZe3jkKfyZ6I/xBnf/kEejvCG
L46IlvENILFxbRiK8NeGv0ExYwldwoTPK8g43ZiZtJ+0Os/C3yL0xiR6UaYEViIo
gvx50k8SkW+Xffr4qrNBGwUgMI0VPTws2w/qaSHozBSThZsViKpIT7ofsFPphc8q
mPPYQoOgjdChxlEART1c4FR4nYkCYStZW2Ah13ksSoJd1tMUua92D0KGwSiW+wsR
zHzG34NVMRP9PLR0nRXf8dewEk8rW+zlrznPzmxFHvf+bYakkTSXzEmlqtDVhQ1C
jX+t/5iySf1qDR/qRWtLnog7Zq/n/ROMYCMPXptuhTy2L6hHSsjak0OVYMi8uD6t
VGKzC3JQY8Ozu8X7uTKQYmN/0Rqujm+ogmRfDMzNsP4nunJBZEhFEBsQMT27WFjy
0r6InUA3Mem57VLYtsi0cqYEfxCf0gAv3n5TaP/GEIHlRJRsnKcZNEBqSRuP33s9
cmfwmwjWJGRTB8cqPvTjwl/0UqVwCvpbLTVGoqHivDFH6io3pixSo6s39OP3hTGd
71lAlhb/hvWGI/1ZrI6hwsLZvO5vFxn+EvBc6Fno99q5D436UK0fORdABbptIY9F
xgA/cgwqaI9fgVEwDeoGGm8nusrbwgleB9ljaQ3mMHhorhyTC6JnvV3l5PbisCnK
lU5i8Fos8EHYMJcKu+GYAh726Cg4teli14NyPVIe4xsU5K1ykmhYwIKcsCTmKXMk
nkIf+Ke74XaNZk5MK271wk9Ki2t3MQ303IdDz4AuaM2VVUNcLNxuijBoM38LreFW
IEOZ8LDnAQbOfDenDbwz7IN+bmQAjLm6S1KdJk6jZa563NBmA/juuuZ06bNEO7Gy
oQ7flnlG/o3IRLpdK/c9DzJajnaDdnmNnbsWIgbSvqEiYGlYNQ6uFTAlaMIpygOZ
1JD26VBkViJYNM28QhSPTuKtwY1DJYDCV5b424/7MHgkQ+tpycux6Gh1483qZdl4
swXXXv5VXX7jxRBQO36xqOK8E1QUXo2GDZp0sG0NlKBBx416Tl4pqFgsn9CQk51E
74O9fFDorPVz08Oc3yDJuJKUV8yy5duFLntQarzmFrZMZxFf6ktHGz7ZqAQEMjXC
soABZlSK0N//i5SInpWMWXLsygycV1D7v0X5KdJXR750DBlRj3TyyjWajkjkgrmn
Ax6soWgIb0+KP8r537fMQ08mlKrn5wQ50k7R8Qy6JB6OX5eFixY+AqJ+2AVcj76F
8gOCz8WFXKHkIpKqPY+0WDwWGhUKGb4FRt6hDhLIJq2yAn4ANl9ukHnMm7ojURgH
g5angHaImJGopT2EjU2COowbc5ZZ4Tpe/uu/xAOPGusVu0lx2LcjvDILA+PxoxrP
XGQFq9WHtb9fw7WwlnNrARaxXUhDs/0u2wFXtmJJBHqbrTYmXHxfTYRZW5zuG/fO
egKY+uKvhZKu5QX1EJtNV5QgKHIPgApFmJkyi+ZYJ2a2C0uBZ6IDc0+NNh7KrXo0
lbGzm+t/AWBz8tqCzoGg9qV+b9CHOi3drKsNivOGqFD3Jst6YB9X05XL6FnFApnv
RwTZnSOjiboEknndVyWebR4mss0qO2E4DOft/RKaP+vRwg7MQPviGK33PyVMVGDt
27ebqLcDrLsDfbGfCY06U1Udo51fXYk7VDpKcC9Z5HcqvRpDep6xwN/ZoYiBD/6F
n8ObWFVSrLiV+IXUXcezV3PkFlqUIlcmybEebTeCH7sMMtwsgA+38zZFTaVgKNAT
gdp/CLmlN77ZGUDT2jt/uqVFouTHF9qeNyEm+gA4H6yncq8WBRD2Av1vJ+ywwCfT
np2vsOI1GhUmnQCl4AelUuL+I10RKb3sM6c52eyMHjr/U/3YHnNvenoBVLWv1xdD
BGGjDeefX3wAWioebkywjXxjz/1Zad6/sR/gVLafxckT+vh25j7oU1RixEwQtIyO
nWGVoG50Go36LoVQMIoEfdfsXAiGwwrlEHDuNz6OjSq1BESl31qHfsN9ctb32+sO
zXNE3qxoEm6L8aEovNrdyv1gOGq8W0QvDDDSx+u9ktJZBCNbaZsrlG62yTFf0uE5
4Q0GBZuCnJMob3dVTBXVU0x9rxX0yjzW67KXjZnP5qynyKzILS4QvtNEUvzhsLuX
kYjS8NfekitzD2wi6BfYD4elSLAYAcaFTPBK/t5wxfJQzcJUQ+AHQ+Zn4tH3CEEm
ttFmPshR4MfnNZ3hyOvIUFjDBYMWjZ7YKY8vR9RE/I1D9JSY52y4Qfe38PWTid0L
lJD4xcvSHtN+rYXhF3TQMRdUyQGw+a9bWBx0KckF6gQGRdSNi6ZRsVc4WbYcR9AC
Y00dC+w1dyc9GpIBPfom1KeObhwW76mNMZMaJrhIkWDLcXVZfRcrN6ByRyfIY3U5
BXXzPWE6ynhIq177srFrLouT2ljkTXq626ykG4k3EnLi6BhqKmRk9l1BMHWy8Pcb
+w5CK8KKKFeMibmGsjTD7Ivf02kC05VaK83yc4uN4VOPG4sQ5RzmcrupegCsuS21
OSfmqPhh+joSFDaWwjobfdFQRYTkMsN59JlhN1+yAfw2Z9hWN3SOzIvdwN6Uy3id
Ml9ZI7QjFtA/uin37CTMXz46soLrckHgLbVYu8kAXq5eg5vesoDuHiEXV3wao1Zx
nHb0/zAdj9CySwq69p0JmYr/LHj/UZcw7kXSTBUCVobPtAi4PsRuhwhwLIRBOVhG
gJjZmwxH7/5QfrxpbdGKKLTyWfbymzpjRy65vP/1pYCYGuEGHNoTIYH79yej+sjq
7808ejsa+pPdHLLj2H4I15Qv3Qe5TLMuqhS08Ni9Xq/HsDZu/Q46+JWce79J9qS5
KCbEAwvFTxyy2oNy8PZQoqb994daL4qMYwnLwfsmwWFBwZf6Cv8uLt5tMGg7S1xd
KfDIj5y3HPWl3vERZffAayWQTXU3LqGSSqfZwMFyDFcAKfi4yN3c3ucIX8sb7oMx
7gsPadOZw9vfocJg+9nwcCKpLK9gG7NyXPFk7QoJXwcMPA0NBW3X0AdERDBz7dP6
zChh2j+NEISulwJsZokLzYH1swKI1XHWdXroc7duTF1c9drpo8H0xG352++1HT4B
fki/T/9vlNGll8QfSBoWyLa5lKh8C5kpSjzDHIyd2hlpTZDpCb9kZJ80D4j7ls14
qmEYm6QDQWqla/7tFC1jFfpW7Ae9kmSAfVqtHaqUpEI41a+l+sq1eRrZLE6oo1E9
hR+KcQsoDg+cPfk6A3ZkVGZ01UZOuv9AWOyLWKX7ly/quk+642PbfAsp7yK7Tg6m
6cxsJ/v/ucPaom9K4ekXYTH0BeiIrGA7XkjKhtMUpotDHUWT6d6lP2mZF4EarXuC
Za5Ju7dqUUDFMqCo+pPMtZIT/AfNDvmdsj8QsdNIaul3Y/6ajWaF6MARtsfbTfkc
CKejMvzAavm7J3PJ4bKBRndWMZoQfc5m94bLpSeu3ZB/75zn66T0J9J/HiUT9Iy1
WbfAi5s9s/I55d9gxYc7R/aFS4XSu5s4V4aNXHvf92Ko8z7LQ0ze1L+SZ19rH1HH
YzO0IqPgXCcrLS3o8Anj3C37rL3lx0zm9kMWiwbnSIUIzA55Srhw5L7z6GojH0H/
DORIWD8oaxEXdseXaotjFYcyNt/C871sKdmLuuuMNwPHYntsBxN3vxUVntWVxzXu
j18ngjmpHjl6lx3SkBRig25EeSM4mbRIMuo56rk4nzkbpjlNQ/iIllvgEDO30LCg
T7qfqHfhEbsKXwBBG+OPXQgeU8YLF4GdG6ooO9K9ic2JeKkbgWwxRCaH9MAyPv8w
0XZPn32Q7hc67Nk8sPLRcP6e12jjhXEn+VZrMLY1iaWqus1qfTzvUjtdxPCeFMnf
1jbj4btR1bhIZkF6039ybeYGWSCM4xv5CC2vkmS0ShedqvKRaghVjAKwpn+LsPPt
up1sEszfiRCesxlmJt8t91gLTh7Iw+HHB88N0esyd+sPVIy1ojGyjOUCYFy1iPmM
92I84vvwqXbab1twCqwo79HHIEcrBviur7iUkKYH56z2yL3F2o8hXcl9MYlVb7os
2VaRDzDby4aoM+JtKvGfuzMwH7DQo9VuOTk7wekqVipiOLM+qXrsPrBiOU7y8mtW
si4CQgnVmSfTkatPHAi1gaPX3OZPetfFpoUL2cIwKb+YGefXyZP3z62Dfxgl05Lm
fCHzc99Ojfzz2eBTWGnrqbM0RHBl2tCJohVR2t7FpEDRb/fqb+w63CfEDAZ3o9/p
xr33PtyewuGgEPMq/0QkO6j7bMxjkNbswvjNm3stE1sJ7CbiObBB+sa+GiCAgyw0
Gcs2cybZde2JNvdLq4Y5qLCWvyhOF2FqU2XTYuEd4t1mCczMSgrYvT6dncTL2bZg
fWZ512iYpKlxtUm2Rkccmi/zVV0G2I9yDhVLI2c59e0RQfqt5LCGkUC3WuEHzMdb
Z1mLx0rZmAJAud0Ft/KF37JQgxH8SHCv0XmcstzIXud9BLE4q+A4HE6tv9df8piv
fpTuNuQNW6dxfevGI6NlvMHDG3G82rI3rlnoPBNDYhuMNATUmYp9WWaiwAp2naMi
OGZbAkS8OpIeDgKylOIJjj8Ic0DwJskBMw9UIxuZUB0beMHo6YTBFhL6r6uC1bxk
HJEi97cJF6TE2cyywj0dE9w5EDoqy1WkzOniLs16guudRU4fuv0lnMjfwj0TWOvw
yD9REIVH4NzRDHigOEDlcnPfy4cjA5RoHrzaMyNEn+Wi4LH279NLKPrgxK43RyAk
gH9dbFcLk049Q3+eTIjwvIRdAyC/SjQJAvxQ0PgHoaqEttRlCoGEkeJlOH6o1H6e
7s1Yv8QE5GZIRTlCNWNv2Mq9nL1pbXl6yWrmKve4Mj0ELvOxPOrsXPdR+dzk3yM6
wOgA1pipvegyq4SPg5mzThCev6Tu+T4s+vhosC8WKrF1ocLWulvQvnFWl06NcY2v
D52boP5iExJwHcdVL7DuNDE9LcmNQCr+wK0RJubWKklAesDU5eA5gnuPJOtVK4wG
/VDjHbIzT1K7jpzQPm1YkYCYzxpd7XTtaN6+E6CbeIeWkRWC2m1ykcyGZN7oIMcv
BUID+9AMetgGaWL4uvbqJkiBVGiWGP0jWf4l2fHZ7078YphZ8q8ivtoTpUUrgj51
Y5BiTybQblPy4FRlAFO5qtdMsiC+zXkB41pPvbfb1UrJQ8Vp36Si2pIlY+wLB2A6
glGoDzwpBIGl9A7GoPUsDyyNJ2lw/q01v28+an1ceSVD4t7DiOC+CAbrSH8BZ1vJ
kWTGNNlzCSVVxnYPr5hIByRuuw7IvfclqYTUqtjSnyzoQzUCP1rjl6jtgdtk/N5U
fKJmS0aBO+UagrWmy6tpDmycBuUSidjmfe8yBxyriNjWd/92Uyy6hQ6xdkiYyIG1
7RXKanKc1q9dmI7Hn0E0VMQ89BAALrXThC+qZ2OFfTJM2VRwnowKTjUyWNuAwRZZ
fopNOhF1ktT4qfqvQ6RTL0dwzTTtKH1s+oMYKVY/ITjdcDp4nGgfSwV3y8viQRVR
LaSMHfl7Q4uNlk5+hNZ6PiTBsQtTYFjY2u4MsAOTHG4yrJxjQNEUoCQs0+VewjSh
xx6Rlgw+9sj4g0Cg4EWdiL5If9ordw9qlQuxiKxowc0k0XKvCkJZKX4CaZU41q9m
NIIkC3a5oQ5ex0wDh113TyhwJt/IaDnAWW1kdClEiYKomyRsB+jBkf6l9sBaUPne
qqH1/X0YZK+fBM98MuIfCVmHRZY9+R7qXYwKC65iJKNvtBiwvHNw2BM3WTYjnPbq
geiEiiWHsSlVel8z0daj2Nvlw3gVy4XMXx8GHTlyrIhwCih4HmMt31s4k2wDubcu
anIGzzGpPZ4F2Bb75tCXRIc1S1MuBc4S8w8FAlgfN5X15ow32l4hLw9T02Hr16w9
81sl/nHi+bI1gDF886ioApOX5mlpfzjqm0EdbkqZc3KK+kGmW4UlLG64apMbAwQj
p+i0p/vyVBSqtfre2TIhxCoVLHwpfzIfMijGobheHKbvMyxxto1g8DXwTfcrGPlU
riAOut+DFgbVzK7PjmAFSUYJ7CufxB9GjLA86EeesA4H6Q8ZroOBDpGJl7+9h7Y6
F9rf1ZLOSaHIt393PXaLjMLHawTT77XtsOc7QMA/S8M5oFOP3/b2XYqfJH7LRM7A
Tw8ZBj/HcfX+J9cRgPKzr1x9PNJkjAUi1e58wphNUKIDcOeHCsfA3qAQe7aKjLAJ
uVRr6aNn0MhmJ4JZhSQi6hD8PKMHhu6U/3+BeK6Lsdy1Wi3qDduYsGf7c4WJb36H
IHyaCy/CXUjki7/0CMoXOiuydk9YFcSZorffUA0o6lMj2BtxtwxBD9TUPPzVO0fy
/uXtX7UK2WvQRuuJ9S2TqvT3XXhdier5hTN8T7srAkwgdQ8HZ22/TNveORah87aE
akX7fPJZtC9xSnUs9rqcCAKRYR1bzdBuFpcHTnymc0V0t9gPm7G+3dr0QGQBCZZc
2EFljBZidF/TMJ7IxIGt6VhLy6nnKPgtUVRXPP26LH5GNTeIxyPIkeD9fROIGGZW
H+FYyH9E7ECfrHXjGEoSXETaslTZItxnAQIjzrQrc84YfmMWL9WoeWUeBrcri1We
9g7K1FxsNVSX4YmpdHGJV2m+KSJhX3u6XoufClAZC71veD1YQlXtdz6tjShKcUzc
69pa6OKSq3FNgnnz1TXYzClWVxapehnlLSdzgvk7ISeIJQd2IfIzi7FSxSbIg3K4
KVbEp8c7iQYimuT3JtAF1ffnk/Q/fAZXp7HUcOFbGQkh2q9VXMJtsCprOYgVDEHd
U+xB9k0IdxLl2OdavL0Kwj4+hojbvPghKqio9yiZGiFNy1xNYv+4BdhaVH03B6x7
/zIa1PBmkoQYym+kyD1+Z1UUtWahxiqBbRG+ob8Y+EIHP6YrKtvE4S1pZvWxDtty
1TXyi5gsI6ZkceNfZy3LHMG8Jz6mRWIZp5mOu+lP8cJDnJcIkoBPKkWN/ksxSdxO
fzGmD1GMj2AAnDpfMvERvIbFkWQVsYKZmb0pvqZQ4ANwBmerbifDoOjWvKzGNfRl
BwbDpC0W77XOwCPCtcQ+7hMRUd82TSEaw0u7iEwB5Do8MSEI+2PXCpI2EJZXwatj
QBOn6SavN4wvtx6H8wn62jKVrYzACEU9GE8yq8jUfYtNTv7zXmDGfZhY6hYUJf2L
jAI1vNw2+Uj1Uj/zQfhs0kWSEeKc15pHXicHO8nPdWVyobNoc1kLCEKk2ybV4faQ
MwIXdr75XvxaqhkDQiMQwfaQdEmRYwX5rl5hnhgYblvVFdreCOcns20QVGyPPQ5y
TsUVhh976vveqEPbAksR36+O9G/6lXsZcww+BVtG+Z1Bmk45ItrEqwozxUwOmXdP
KUbzgRE2zT0oGvVnuAVTRiwSxBmsmZf6frfiiMIE/QmLK3Ys3Qm9S1JYcaXEYCTX
hMK07NJd/dHFXMFFwUT4uVZ3qQnNyrxqieSTMoIVxuyNpR4BuzXf+DQxGLOKrlQR
UuuG319QZEQo9iNvVGeePiaY0cQgLibqG+64aoSIx8AI79ripDE+mxgjg9ea1l9z
3v/hFL7lpc9i2bXL0tamf+zS41PJrmr4DnBPs+Fi7QW55MyKWocOtY9V8hS2xBXl
6z2jbqoa670YT7Mz8asGYGQJznG4XLWZU721XRtpEcGczKsKb6y9/RZbIhOE9a2V
J6PVth5i9ll5wcQ4beCS4gQzXSPUpzNeIq4tyYcWaCFqofBIBOIL301GCHhOvXYm
13TpOMCOzAWdBY0v54W/1LjKJOcfdUb+fEBKa+d0wfX4qmYp2GcVpwpQQQ3ZA5Me
8Ue/QbXNOD/3W480a4YLYvAvN5YsxNIZYTJ7bm4bq59z6R1+r9fnkLOFOsVGMEyc
WNacUWKEg0NncQ+fOkAvUujmOmV7v07Y207htm6EiHC5+1GPPe1LghOYL6cBG1rK
imx8V80cZGyr8KsoUZ/C6+Zz7L862vTdeqly9bj0QB1bGmO41MD23elaqzVH0zku
oCB4GFJT56DWD4sZ113NsDiRdy6+ljg4g4q8XZI504zVcNHfr2cA5U1gKq4axfv2
t/T2h7QWMn5/03T8M3RA5Wbxm6i+YYwCgqboZDPgvqxHLqkoMp9t7MN7aJhOkUXf
oHW+7GI8lFehkf6VFkGdfAuNFYG060x5JcuyzedrZQJMZeNj8yhjB8rAg6kqP507
gbdfJYt5sq9/6vVvQJEHvI+f99elCj3+MNTDGVDpktksPUCnbA1dfxXS9DnlNy43
XC0eh0KILPA20e98SHxK/XBhh/cHEDZTzFTwgBDkhcaKh1+wd5NEh+oIQrbvIfmD
Ncbj7TqHP6l8t/aVQ1SE3Oocr0c2NxXIYOF0hN7ojYIpRNXwgqDT3AZvX8iw0bot
tVWFIofkW0oWl2Cgt7T3uU+lED6PIMfZ9YZXDfVWL5Jy6FXkZCsll+bJF60J1lm5
Ok5X9au9wPWhkaDYA3HM9ADCcIjmPD3J9G5JT9RGLMwqyVlcN4/fivhLHdHWU71v
VaiEzy7RSFLwodZ3lfpk/ycZSBjOuZyj7jVFOyDZYXf7mk1JZqikjYvSPuM5rwXq
bbkitdGnNCLtIlP0mol2oG6ejLcXFK3Hu3Ir2tDK+caoqlKWnAWWEghM7BqlBz3i
3KNoT63n0Cujd9igEGZ09RcFc6eGIYoS8DbicenSLIM1KslFddoInIEFIjZBOgQH
oQQ9j4Y9M0HVsKPdR1co8HTz9MEMjXheSQM49RLhkCRpaELXqsLrYXoYGIpgSCTK
g5IVTWzYRT/YO+q36jMn9Aug+5S5bBGwE7tNfiuuIZ5ckH/cCJqstHKLf38C3JpX
60VXj6ff38Qe0gPe4kE6A774DMKfNoBflCbJSba6TRF52pwZvzr1Ufoomq80Scii
S6jK8sPwpMLleqlsltsNPPsAJH1ucj368IFJNg4sO07UNq2peLp0nCGxTCAMjBfv
nSWr2aU39P8SKwcEF9AUTbEK7MqXGssO+l8j26PYKO62O1gT1UCK+qyvvY/tLWr9
587oAemljib01Vse6pQaxSjN56JJnT+TZPWmVBCd8ZppjlbzIjeuSdJuOf1cBHJx
zPzYKOC5x50R8t/uSNXnMuJS/fOYZXHDjgWt49ZSQuPKD++zzCOt1u8sEI4xSLn+
RUNz53pprJ4G/SDu7FNfu0Sxvc7HbAKnn7xgpxJ8PKqTPI1oCDDcM3Iwg6WXi2uH
ts3zcgGTXsAlI4+2Jc7jkxK7wGbSe4CxsmjCRQolcu//hRWcojbbWXD8Jjqf7cDl
5aKjbAoUWke05oAF1f+awYkLF9xi0PKp/Odlwj+AGe53gTma9rkO55UiaUTO+OcQ
JsmO/Qcw7hYQ6DLNA75s5Q5YAfwnDeDGmyRSy91jjz+uTxhaNRtZZIvfTo5VdDtQ
pExD6XxUmsDgbzbF3LXgz+5bUP1nz+BAaxoZ2GzgeXBZicvaaWIJkRTdmjcay6Dv
1IXUIqEe/hKc926z6Q25DyRQjV0bb7BVuCYprDfSFn3/1K7uE4LNeLzaROzq/7Fg
bYMKWKqJu0bB+5li/J1kf2ceL9CGXqOcL5kO89C96FjZ4IlO4U/awzRvsOqGSDHC
HXzcqKrcCPK8/aocP+Z2AbgxQrO3sNabCMTgOmLBasyJPHdh87pTw4k13uYSD9WO
m2dY7FpP4b1Yra7fpG5ReVUXvmwrB6gF+rsMBNJsgodQMK2bWu9JB31rDYNuLupI
J447NcBn32kx9TM0tA076GyNntNHZ7qnxlVz/lrP+nh289k3Uo5sjVqTdZnDf0rn
EuRTxgPCvb1IOTqgh2tcKNIckEzU21byvNwW4eE6SjR4LHzsDi/XZm1eFGgAOUkH
2MbTSLhGlAmNv1cPfcVQQVcGlrTrfU5NxBqM+/DQHOUMX/uwKB99S5xoFJynr8WA
3ABJRa95eGH3KYaw4sNv1MQNIfcT+oE0QPID1E/nbzY0tGO4XwLSY84B2zoLRoPF
trc6AI8lboxQ1tlnbdN7Z7jj3SjSnD8kzzlS0ylySDiaZ1KMwh1W0TL9mH8LWMGG
I5v76TL6xPmLfY19Sm5QZhPgHhQ6FYNMSMkJLZ+VrXm5/hlhvusDPrX/3rhVqBUc
MGlpdJIOnmaA43Z6DTSOxbVAqvWrEcefNX+8OWg0tvmuBwDNy6SzXdeNd5pOvggH
NxKT6OUf93VyVW3W7Wwlu7WD3nzhhR7xmkmr1Tqmeuc4FQ2tqwFXkQxD5YHEeN3Y
IZquDEmzl0aOSUmc3e5T/OFMx5RoIFw0MzfohHDSX2ykzArKK6aCfkaxp5gxoOD8
Y74Ynrmb7mWacpK1RDcpZwZ1ZkwO2w6Iix9G/YIjyTeYlfjENd07MNFFK40riAWc
WxGofzqhPfb2N4lk0BUZTpMmTggliPaOH5SaEujVI9Hr9yaF9Nt0g6YvadoHoXAF
uFUq5AFTt9DsEQwRmMsZ5CaEIlmuexyZ+o06i5BPX7VD7k9OC6gUg9vLCuE1QX0n
siVuwC5KPZJGhZ0VYdWI6m+CySshBa0aHPXUFzPdu3pVPeX1Z74Ez+eEVqZCnlDG
i7dbKPWAICZn0/AAp6U5rPZU+Nkmxa67waZHuQk8jRbeH6PHIMxfsBfuEs7YMBX3
gwPrc8bt+Yu2h/cDBVpSwIiZyI1NhtGvRayjKUMdqqKVwTciHtmPxWDvVxpQ7AdO
zWjKEYglGxt4A0OXztPBxuXz6ot7VZxrah9DIq2HFW5dK272yvjCBv+663mSoU85
dEE7PGTyt0H8x/ThTHI4k8Se0MvCo4WSYUlfegXZfYB/3fno+w+z0vDyzKKs0ewW
JnTas324peX0B9PRN1F1juPCb7S2hShLu2P7VkbE6KoZg6xY+7Q0nVlbflS9T0nb
33LP7ks7dVg2iFgROjvZ/JMIeMgrtzbaqG5Qe6r36v2dxgO/uf6c3tkvZJToFJMv
CCFSAvwnhKhF7iIQ2fcpn4VZRHS8N4ZchNqPTs0kEppKTMahGKlo98mtbUt/VALF
3aNXZG521LCzgQR8iYPnhZsxjLp+SUYWOKcCBTpXE2e/8tSqDe6h1b2Bik4BsB7Q
QCoRsy8O/EGj/GQgUkF65BUm8qCFYKUxLDYSJctpL5Cd6tEfQQsBJklMt20LxwtP
Nfc/G8Lsz+4sR9jnbLORKA9KOFs8RxUZ0iwVhVXoTH06Q3HCxzj8kN0hzCvfYtAM
t2olzIG6S5p/K3cnIauSJfaKZSXL62/+h3I+lKtHmJRdbtyQj7/T/s5bJMckJB4E
w2NXkImFByZypPr2k+jxkLtRlWIo66zgtOdOuxpznteDCMidE7lQJxtDNZsX7kDX
QwyPuG7y7E/9JdTHCkleM5D9GwUM3rtsMgEG5EnULzYPYs/b3AHLhx3y9pvtjtuh
Ju9is46WZpVeOS0JY8nHO6g2WgnUW75kib87TmCYLQ6B1jWdBtDsq77ki4FTKdPQ
eCQoBNt7OXm4Dg6kD4jqgNrdOQw2v1nBSp9YaEbRNqpivfIZf90aFtvCbyGWXtYT
2+zCVd0MJ6WQZ5EDPemodPh/7k/PD5BzjHGQ+t2MvN/SnaG4/ucsPPmv8TRLx7Ps
HNLOSmbt+rRCBjZ+B7O7g+eVWB5/neZz9IaVcUo7tLtqUoWZ+aOa0yWuK+2OFjuB
6amrR4Z/0p03OpSrFr7rDQkOdHhoLU9tvy9eQds87a/kQfKgnsWfSywivg/uwc6P
PaXD88AKda5GJPb42co8NAdxh1fBLpaqPhXsiGp2t1+69K9CIt4iV7U7skr/kpvi
rrgtuW8gENCkY5hcS0iAHbUSODcWKtr+0Pxqn5YkA/apPU93281fJFb4O03HuWi1
iKnXBGwHWpk1upO9dCozqwIkg/Opl41qp5F/bhvbEORaLiM3S7iKDIm7hteRCqjv
dVm/rIr7BK3XAksEXI8rEy7XgfWXQOTPAZh/nQnEr1z+z5q6cjxQ/WemSL2fVDsx
qyHBmXpqi15JPkcLHzI2ZLK2JfxU7panFXJDQyN6VdcAQ/WZQg9NsgpaH0AHU+ac
kUXDDTwWxgmjGIt0+XuwEShN6HRxY2ajVfbYlloDjZHl5cN1qj5uOXYqYfE/Fs1W
qiZFG4ED9sgVzRjHmwQi6XYCeBT5PWTMFfC94zxC7mvzirYZdhjkuS+KatQiCflx
qdpUYS9YB2za/MnTbi6SYmR520Llv32wbqyjb49W7PzfgRsUyFNQgAWWVgznH/VC
BKuz8pxD09T90v8IML/0ITBLU7c08gximjH2bxdf1LKxs8h2Q+43V0LTKRsl5BQ6
UNwyPughvxCm5I8OorYS/aR0QyK0FVT06liVYm5O375eBZPIyMVR85LzahogWxwd
2Ur3sB94p2FfPVEoVijjnYKdsUWJODzaBqY9/pndKP5BdOJbGYFxxvrKsveQcP+m
1b0YNBUhrJG7ceC6y+tF1zC63bSomj+kPeAaeVtDsnKrmsd+tdJUDgA4nQPJKMd4
y7QoSXyw/grTaQH6NKT3OyC7M3H3lPSIgrdXc3lAeBq4nm7HPK4vQ5aQIkFIxU8q
KCiHLUksF460NEPbIXynKhkUqmdr8ko4SBVdbWivrCfsSfJoKemGAQBIE6w4lk3L
y4EU4SaT15q9hG2/AIuCWwq1uRPQKaPdVYRh2FNEqyBXd53oMh+7WI5k60Qfrkic
X+jBS4LP8mZU4fXDmWnbvNT0cPaHT+Kl4Wp8aPa7Zds0wWtWYEJOJ2/4nko6qFHW
7jQ+dGvu8Hvt+st7kEw+Jdqdcr3CK0vOGUImgP+FdaMHKzaLKO0NWqcYZP8UBmzt
8OFEqUBEtSUirvkPMD8ddhDND+3HxL5UJEat5zozaEWbDuwjueSwJQjq8Vo3Bc+p
iUbANQGWEnaX3+hwXd4QSQvHoFv7bES0GgELeotpAy/r3yiUVJIevpuIoM2yQPPJ
oJCf93OMk+TaTAPCh4tpjJDZW46KLtROxZS8+sQdcNF48clwozN7j2tLlc/Tc9Pg
bL7NIkDlpbzm955X0H5O9TQ2OBgTcqlSlNGnZV/qg/0kFUHDq7aQFMMRRFhss5Nm
8FO74d3AMMI2nh7DsjF37ROpTUvPbsGb8aFXxEpu4Rz555KLmR94Cwszw3iBXeRH
YjA0iYZ80AwrYlWEjRv28EW+oc+ngsBVvWw7oKtZ896VGFlH6zGOaczkQX1PqNHk
XvNFcLY2UPU8ghyajix9SQ/hBQ8vXm8xt/6Is8nNNrib3cI2sOgsxCmtMAi017ji
JIUmdg95Zkc+KJgfSOIpiilqO9O53R/JTPeEIae/gCF1CEydBsKlSMKZjtz14OCU
zb37AZbWqLZ85TMve0KIn9Q5V60rk7CCzemFfekxKyAvdqIvyCUxohMYpxky93xH
eHlavAeybnzrWOnafuy8tWPLucKJEYY8qxEPA+ys/rANj7A6cwN/FnaHbm6Ftscl
hV0UuPbdldLJCf5fRJOkSLmCZ1VyRFIHOtbGUIuyHu3lB1uZLFT6i8yZTTsUgrUW
IE9Uak06Ch6VYMESJ6LYzEQTw+gweiw4bgmHPlHP9vjcN81Ck1ImMKePSwJbiuK9
1KvhZmq/t1R+MvIgtM5UpDIOCkn/TAQ42UElm5A+pgpmFCesTVAJ0MvnDkSpB037
iuyezh6dsJrNO+SxVIWM6bbX+XldZF59LJmcyUX9C6Q+ZQ2Mn4NjF0JyIkVcoFbp
OGsqwqdcTj1YakvFn+gakTGWmL0+nMQREiYzsHVYJ1kYBIRXiCPu62d2TNyrladi
KYGCmRkJIF+dL6rEW15d3T79kXIFJVDqeLa1z6ZRVIDiC6k75dzpdudwvFXFrIuW
+RUAIHs2sIOnaLgpca+ojl6I2wcl+aXwG6mTJSacqE6hvrYc/r9b+j3Nn7RM0k0c
1+rn+nbzVQC8r4cxLHhyys3LPQ1mTcBdPyFFb2mPy8dYIIUv+9EBotIUdtitgTiF
oThYTQqs54nH3GObxVBvNhPAk/W5P0o3pcMv8/Eu/LUwX0tQcbEUKV4nkQB3kgjW
QgErfkhMycdHZtDCtSfCVweobbyjkTAOk+9ajb/SELWVYVSDZ51jxWsddRUn3WV7
JmWoAIGXJq9c3VVxkSqI6HBQUHnKlDw8Ls1CaiakkiOqQTkjqh8E3QO6wFDi5FGd
kMxwt8CBsuoaIpZ7EV0YJnpeZgp6cyd52DbVuP/PaUU/uyYEqd4PjD2GdKszcPAx
B5cTO6IueJXL03ZxXcpkvGRBJyanBZKtf3/bEtglf1c34pyKbFmpsMHQDiyINrQS
r47cpeH/DusYidIimcY/iSDSOQ2E+GK3zIfQO+dN4i8cr6KRg47Ztrrcj/o4c/je
AWizA2sBIl9lkemBqL4PLNaOCjPpOcPhBB18BxH2DNwGcceZpjC3wYH/6AU69nS6
P0lKQgDPvsEgK5a75Mo7oBc7RiP69W0l6v4OpqY2KRZqz3X83AJj7TtW7HXpj25s
YcIpD4Z2/fVjJSiEDyEO9wkSZm6k4cFBRs2O4NgR3SHSph3GBSbvEf+MWyLhEM3q
TwdxW2U4qImvLB6v9+0EM2gP5FsJibjtBguB+T1Bls4Vkom6Gn0IuCg6S2gzL4uB
yzWod3npbWH24BVeju85bVgHSET2duabKTyx7BDRd42UX9oeTjbliOS6x5J2zq+4
K2B43HCrq6ONACMfhW3TX56UmpcwL1QZH3HzstnjQ2ZhxXaBP+nr7kbvLLU7+QDL
o9l/6c8CU0F7T3sFngsGCPNuzmjEeC9p5AbEN9waGpfwrBxdlBlcr7sVbxLtchZN
W8scGSDZDX8K1xNhwiCQ/hqBLTJY43w0ymDeVo+JL195p8vwnIOK25Z1g8uZp3Ta
ZxhLPjDq4ak40Uvvtsf765lKY1L26HSo88FfQbNYoTGMASebLEB9jFNNdo+QgMGl
mzCniARhjD93Rj1otMM9W7Xbxzqpx68bUjdUV5SevRAjTu8KkZQ4+B4ZCaSnA1Y7
hwhpOQmdg8t4XTN/hX7551Ds9bitbSkzDtkSqZipAJz5HlzFZz8U+cG/XKji+DlJ
iBCAMuIFHHpKAoGhIEWwR37ed2N5CB4pdc1AH8OxPO3u80C/Oj3Jp3YgeVBurMm0
kQtNCzrfddZq6JRQ8XQDAfq9275FALiu2dytULd7h0PHCu3Y0IvHb4fgjDt1TRyQ
8JkNuF7h9WZsK+VpOoPFsseuh+xkCTNFevIsWg2rzT9pgIOP2ZhzcGIfRTCGH9r+
juNCAigOXA+fPITC1CnXzx1SWwHrEHcClUAO/g2HDu53YYAKNdX6m1W35SNPj7r+
3ZJqqfXf3IYik3lWO8GKMpnsNuYfKgzW/AfFvKIBTDNfvqjZ8AjXlGyWz82tEXFI
XinA0UgLjWERlJgHjPsQVVL7rlT3gUSNh9OCKAkSbJky5OfK+xT5/mxIJKeVdZlE
NkHASN0rdBnNgA1lIovw7o7AE2NhkaoPAoCqh4vAtXr9RNLXbrgxKlD5U43VEks9
GJh8PVk6YTB8qu8desfEM9I63J4nHcEdg0Otfw0jclcxZ5uOReSQ8oNrIIrJ0wd+
g+Wz5MUmrT2+G15h8JdFbzhfbPZjD+xC8FMV0rIB1NuLJfFp0nrM3vpKnhWmqmb5
+KN4f30Xvb60SA4dpAG+1Ki0leHTr5VLgyXwVga86GHOrDlJExpk/cy8TJVpmqcl
KzRrbHUSjq6z3gSnQ54GaTWVPtwacs1uOeKYO2VXisA8nWebBw83SHEhHFThEiFk
Kbjy1/Wu1ZV3DEss5M57VfP+UnkChwd8cBbqJMqonV/BMsj5jG1umxfY7YfF/9MJ
RyW9nmo3HWSVkpV1yYcV/+6OU2Hj8Bl3YH0Cstl3+FuyURvdbWC2zysfhHYMJy/d
sPy9Tct3ckElx/W1w2cqDxnLGYg+GVDZPJg/6iimgC+GYoH6exSYwmRX05h+rsoh
O8CyO+sfSDlOshNJXi7u7WNKpZsagvZVkysG5pawuSnL8TsAJpmI1RgfQ9qGia/H
E/uYEVAXmyUS3oLAVfstygAnga0M4T79lKw7zxKty3hWVr0/v/Dhnz7zNlN91Bqx
1JWi16McssF+it8/GNKgNIzafVwbj4QCSsH1GmeFkRDwR+gpSqXVdFKQ1yGTBWKb
ju2kuPpQVdWIeh1UFC14FmJFNZXC4Sg79Ym1MWgkrXGyz68f+1PQH+0ANATYkR7h
69n4UmlxVIO6cNPhlEKuWz42gXOZJ7RFsmGc+EnQpKR1muZql1zgikcQombE1rPw
WoioHoSr4A6PS32GMuTF3DaIibyClvpLrqhj7xDaiBIqkCao+pgPoRfiG0PEBTsD
Z/uIgWb9OEKEP09V02iZatAmV/wKA3RFRZIjaUoU+sCMsyPUTYaKxsz3MwqvJja8
LvTjQGmdXKwlayBJILiPFJVkAdnerzIEEkCkBRckIO1j9QZjXC1Temgg2XTKSrom
WRNehCkVHaIai9+cAG9N1eDhAgmqFee0zDMTfn/CS/r+Z+JEgwt8zLz5OcSoxrA7
TbNhMW+MYjlcfNsNKOIgiEb/Xsx+p/ZYnS2PMJplg9o9ob1bia2O2mlKQ2mgsDXb
v7cS53Z1UF8ZJae/JJh+epDAxDS/bshJ5yHRRhol8JLRDi8e8nYlkkUMYDHYZYTF
3TgCiMSuTGz6/tfR11v+b9AVS2GjnRWzClke3iPa8rlFsxRd2zwbBxzraDUydJar
vSVcpCx7vHr4Xq35XMdM9vvUaXx118oGgBoMcduV9ig3mkAlXJGFs/wDlocDSoSW
oexvYqvcHp6kahlCcfeZAm4q+xsIsNjy4Nx5akkzUWjjPJbF4n4gojvpZyW/qKyL
fH7LCidmDa3JezxExfrArM5uX5quNrpJ0yECq3bI34+nNlcOOUNKeIh9XCYHQRBD
nrcU1tR27d47J4mkmwMrpGhCSh1ybQ5/YonL8GNoBR+ONx95njRrfmwgegAu8R++
AcEmbcg7VXImKBqFv4+7Be/OWOTo+ph4miuHvAtieNKczuqaEIzf6znGG0Y8lG/m
rSr8OdoGOsgb+6/IBg4EherKGbOEue5u9M9BAgmZiPJgh/A5eQJD77s1hz3qC0+b
F9vI9R70PeWM5EjjwXJtbVo8E8hS2ge8uPXkKigk19lO/2YpfzAB5kfgpy6QUIwH
JK7YtWINjaCVO4JyL1zITumzt7X1orASeJnWBJ5ce5Mq9UuRkyu6ilUts69+uPtG
YR+PO9Bzba27Hnx5iLZTJRCPhwhB7ynTSQlrKv5y+A7YiTB901dQn7hBPQcOgyCi
mq3Q+lGXXCv7gPMHSzTgv6g5uEmd0FM9jVetWaQPuRnboqBByKtA3vaNH5+wCt8a
3p++RXZs2M63qY+7JZJef7OF/kqAQCPhja8TaH0QVwaiy7AYaDEACBQGlZsMq4ah
G7CJoAGifqF/MPRqk2IgyTZUL8kFkkAZeQNGXgUshQq6x4EZ9fRey2Gvw38kq4nQ
TPvX3sVaRrDYkBKLL7AvV3WaLBPf6Pmginq/s+t0HHIvJ03453yoN6kZDQhXA9KO
PUoWUY32+rodcCaJCTpYzBZLZkaqD31SYdxUngUiEwApfJ6ij9Ed5I7axU6Xlpkj
h0BtJHwb3g4rqQSnI9jbJBWuQPRQzFQo8G5R/BNASmP7yivBopx7/RwRulDyp4cA
EsCYmcnqmuO6V23ncYgC0iKP6tSToQ0pOMhcyu8tqUoCbGP3RubuXI8p7xUEYE9P
y6HfiyrMzkpF5QRzX39na5FrkddEP01peIi8mhxNVhEhkqHcwL8cPj0XBa3RXxnA
Gc3sSPjYU7/jj6VaGZuaydtw4FeCjEjitNyOjl08kkl9WFksTSn16IbkEx5e0Qa3
pcOjIniuZrHKnvpKenLS6akY8GYCCPi1G3oyuALop0NQnPH16D0PWwl1piUgld+g
XGg2TUTd8Ptq5mVSSxUy3uniCOu9h9kubJAFeRNeDOIJqtB3px4Saja0SAAUrYyd
oT3VcjdM/1VEcvTnue+691ISpdl3QPHTOcHX1pB8+No/mij1aAXE+N5Fuk9djPKl
UJibtbpdVx2qI0Iy22m62LZKwp287GkvjOJiB2RRSlQUIFvQIBfAGcSjzjkoEym2
ercnboLmGb46n/cbWaMICJ6SU5k44RhwMwAI3OVVTCejrbLesx8TkYhJ9PSE7NEO
Pum7Me6ocgu1xHHlWY1zrBosFpmpk4dMWSYY1gKnVUF/SJjxw01yxFUrhyHiZe2z
dmxYxOAcpEqCIo9Exkpmatkp853G/1ZUaS9ctOn5tz5amRGvaP9Wj1Ed1Z6Lg4hb
ISDO20RQ/QG5sTqFk3DphKsLc8hBOiPj/NCi6nDvwu9J/5n8fJ/gxXcNXHlb9pqT
A5opH45u+d1icgevPZvFZUY8YZu4VqHewlnHpB90AiPrRM+VNPCSuIKemcRo94Wk
ael5tQ9btzaPzp1UMM4X4HRQA4djkjWy82T5scHlfuvXm7ajP0o76Ce90VaiunMS
VtQZWv5kfRDDg7GDagLU0uslKGSy4iiqtZucci/wyxS4c6A5r5umoxonewhGxzhU
CztoI86wy93wFkEyqj/9r6AL4Z7H0D1HCPsuRCp9C9nTGm4BuOQFjTzuMOkmjvYj
qV6OStbP4m9yrImVVjGDTSNPnjQuvm1USiL8W7xVqfAmro5St75OQ1iewwx5dLo2
rhbHE8yZXstwh/alLfVmaK5ldVLoRPQeirii1Ven/bbNUf7ZOkdS1ZdSDfMiKNgo
KPAq60c7CJTjNi/4dT3E95tghzZO2MG6JLPaxj4cAfNzMMC29dm3izFIB61J9cd4
J6nYkbfKtQpkCiBUOw1/SYUcq+Y+5okrdKo04IW6gD91AhnKACBQCjQGUeXr1ON7
rVTVLzL5C4zmsgCMO0KCi6sH9OzfpCO0xitB1IIxe9tZp0oD4lxarLRg9gJg4dN6
0VF68MlCwiVbosZueIAkPiCCa5V1Af48crBVowtgp8/+XReyXc2eYo6Xs3alTbyJ
3waFC9rWjrgvFAoy0h6nx2wJaEGE4Hvd3Xh4YmN6QXgAAw2sfqpYyN0hJgx+y22j
5VOhQilXWvIu7sl8e9bfws5mLaVk7LVFrcV8Ye2SPV3gAMzDHsUh+rYsYiblvDMr
Pxn5igYqXjTG9nPmRxbdGBmpdxip+FH1tIF+O1IMtdlOxWIJWnGD8rz56U5SMhXm
4nptBJUuWW1OVPRgdQCjTSQqAP0uDSnaB+8vHN+4dTCUxIt+mbPKvfEaX/+jS7Rv
ldjqxlKJr7JSt8ccC9JV6gyyGhQ3i6fqwifb7hxXSGrV+rvrTHQFFabUY1K7Ukrk
32NiCpnPRY91currdXr6I2mJ12Re/tkjmnA//x124RPlQDXtkSNyQZsUFeTa8ugq
gIgj6cWhHbncpA1GfnEknrUmUflu2amENltGtESDXf4MhAKuTsRZriB2UDnNJESF
dfI3hm40gKhBz7ZBF7EV1Hek5SmV1H6S79T9xmsgivi2H/kYnp4h179fuXFpQ15/
hwMaCIIJu5vTq1KQtLOYbip9u3gSLnym91eq3X9VdLWi3Sw7utY3VFSLlOfteZkA
NepkqRBxxaSkYxzH8IgvO3kPcpjazuTLq+ipVvYtOxPZi3nTR5PjAR9ccm774zQu
rlS41ASnaKErOLfhM5oGDgFzLQRHU8Ww87DgWLkn+YEqc8bNoAjFoaNia+iVmWrb
WVXZTfQHv7ZAbOr8+tKqCEDAhLV7ot0P974vdG9gyc8/AYzAccGMTlbi54HuUxKE
7vLaWPXqBoiPQu9cwS9KKqGSYFWpdFDIICVKRaLOabD/51tSB4A0zTFelO2A8cI2
Mf1EtWJEGRdehP8+PbfK6ITXjdznuso2wAEVVfzMeKrkvT+wWWSYB3LnzGI51s0z
ytupEWmvRb83rU5NNibbsyFSyUyAb0OP/KdgEkon1ApiqGTsG/vpHLzP7yStmuzF
GKAjZ4QweK7Gx7eSe4Q1B+JBYRlI7s9ob9X4uLVSOILLZR2LpVGggxl3TdYYrp1E
1OpFIZ87hlHfSFz46iJiXQ5jlhwhTB/feBARwt1GTk0TUoTAnrdBAcOTpbzVy0wQ
0KySz2MvUBSGU80f9W5yXSfkyxiLdCNgDI4UYtXSPOrsRrX40w6cpqnMAuEobqtp
X1qkg2FQSm6JKHoQ7FnRb7jrRUTxKyyJvlgR8jwOMQ5zq5+41Mfzv8GbHS7DqUbE
B/wfC+LguixuRLI6aVMRBXn+IGuHsU5PzPE6xoWquaY655vE0SYFPyrSse9j6zpH
OwAJ8ukrvJkKoD4hIaRHEH2vM06aWOh8io43l8H1ZipCxzLP3tamujnUX4orLohO
rGb8y1yp5/0dD7sL0AoAQqXgiuq++oWzbC/0xDeEfyAS2NxHtDwBM2+6ZokV+gWy
h+USFkH24983w69+Col6Ozab98YnAdSqA4yF1TnSeqeoyqmxRLBhtt9JWeKZAcLm
4G8qv0lLtm/thJVtiCEcRyMIVAuLJVDLcgWK38r9f1n+DqqrImuoxl8vIRf++mOf
alMRChFXdexz6U3LyN/BEEj8pY5SAACTxiW+9Nw/gAB+SJICn6S27Npq95BPM0tK
6DOuizIoRz+G42HzNJY68/ilMFXHEKW9isftMPr9sKK+zcJw2BvkyKnVHXdKnrlD
g2m4DGC6t3cLxhtPaDoRW/7WB5XjoQBpcxk1eUWGlVkdhRtha/hawPR/pyt5YtjX
zfN/rtjawOL4LDJcQ4j3OiZl6ddppa1lsEK9fGs01tw/miSxlFUhG7lehMeyDLG3
3HfoKHY5GtMo+yqie2CGFgX63um3cY+rdeyFsGf9ccTMrQ4Lydz/KLaAHCZk7Wjn
gAIlsHu7A7QFTDU+2zHIom4V+ZIKbesQFhhVt+I+sGWM3Ek3dNolH5vViUWBAGtt
+yUd3nGARJqTw9jOtW3t/qkhd1XIF6ZXZ7XQMQwBthaIrymIWX884lGC2tt7MdbM
B2yvbtZGXKFf4IVvg7vEEMvyut41lX81C9Qdb17MekJige3vO2zWcu0wllaOekkU
1TZKTbQMQGHATayECLYS3osMH0z3jwq/ZdMj9fLNWzDDKIyAXznzyvCwmjr5wv54
QyrIln4bhMYd2+MZd5Sq9LSr/TBXTPcI3jsEyAqo5dZUcinrxihBRgYDn6PCefj0
5reTv9njklK6evadlnlJ9AjUtB4jz8uJ4DYmp0gTuLjC+1GAaH2XTmktk4K1IeYQ
Dz64MnQ2ajiHfKZwAIUQMRMoRKym1OKBJ1Ma4/NApzitz7pCcUna2kxzJ0/lc6Cl
aJqn0WLTyMbQkesh7TSJ+3oTIhSjtovWzSZOTj9h8YeFItRg+YTwOBE/o6QRyMNM
jzwKMj9zMXDZghIawoHm+jgplNWM/bSEBxpsuhGBjF8pP3sMrGM5XLKy/Wr1TUQB
vucsdX1nOhurVzxa/4sXGZDgMBiLA7enb8AZb7Es/z1s5ibHyWN6noxnMxuQL4FZ
+ZH94AYFpQ0McjmulbbM7pnwEzcpA87gXzl9BTMlMfpAuinDOYcLDmqd6wwzpSPQ
yK3k0H8SYJB/x9Q5ESR0inQAMjLtLrc/Hr+u3fDLBvC715u0nvJJE4qI0cD6v1rF
fgKK/HmjZ9lqCFrA7PFXyoFhFKRxh3Y6V7+Dj+03UnIvCsTupdsX1+MN8gtZruHO
xoyx4zcI1R2Yw7ikpN5nDXWHg55yAUglFCFfK83O5L2RRdidzIGEI/FYzqobWjJD
ba+UYbQC6WRthVqE+GKi6DiYZgaq/cZjkriLk1IYJGDP8rckSimA9nUvSEddTlFy
XDtNVsfQm7CmrZA5I9n5qxED9RA2BKDMkMGXi+f5OjaQO01yJKK/cPoD0SmOzKJp
Ue+SDXtiTV644iijEs/MEs8JRS9CZnlklZFORptMdY9ERIgc7iTQtqk4zNZlbRIr
GR9kjH5Dw5n5QcIRJpoA5UsHMMiSwxSBA+dXt5O5Wb5exYw2reHLCY+vC8nyvwzE
YetEN3g6vGLKW6qHmtaNBCCVlAq/XA4o3zpmwwin7CcDnlebwAUSjHoR90cPvlRq
TyeQOS85riw8ZA5e9G2Gg0SBpKk3HW4ISWVdjDQ1L1emSztuVUmmBrYxsl4cIA9F
UFeYsDtFywzKOHDEj97Rwa/qWSw3vXCjO6vjGyuAcFYU/ieaz3jHDf9BpCPJa1k1
x0MctZDCJE5PleQ0NYOKYnY7hI4KVwmaR/eTF8H/c6b0gXBQk79pG9xPQMU5JlZa
X9l75i7AdkF9dv2WhkUcXnVirYytV6hH0sahY5M1A/dnI0qXFkYpyeTSkIZx4Dev
ESWTPufB/oBetFlvbu2IxbIuYTGce++LoGjj2X3ltVTXDxUkWQ17KTmOPkX3oedn
XrYR2AfbERFMfDr/28q2LVYxqq5ESy5S6SRAuSi5Yk6aCNHwvX45OBXKQguHrhRc
nmo3F/voNYy6bC14vzVmBI73x9rwBfALCRkxonlk3TobiGtGQdcrUA8N0xKrqrMU
b6LY/Zg5QqyYaO93gS+AaWL4ITfksj62izPDcMx7Ykl1WbAxjTQtLwGRTa/Mp1UH
YWoM7Rc+b4l4BnQWz53WqagB4hSXYu9JxmXO2m83BuV8BoHIOwII7F2gzgyxyvst
cXzfrUY89e1xDdCsix9ORv6Zj3mV3w3/WBq2ewnKg/jaxTXO1WzWevFwdOXmcTaR
UK6Lv5YIXjxPWBv7WaLzqefFItq3lKeMjtTHH/4aikTXkcaYuf+q2qBOCGD3XkjQ
IK3y9WHts5yiyFmuU6g9/OBXMHODviV5KcJYdy7Pdw3LWSZXBoO8XzUF7YpSreWc
CNkGDQhcPdNhJdzF8boq3coJOmQRdAlvywG1nDkz/F6wAIX1aPeBoGQd+T0pyw6Q
JomH/JpHTRJiv5krKan41SVx7Q0ztt3MOIH6S1/qV2fftDNyzYZflCFbzrwAfjPn
a5+oS69Mwn/wZW8X28sgg/a2w/mJro8B4Y4exid0SftqDQMyA6Pc/9WxvOI+pHxg
PeMD4z7tw3LMDMkdKg9/Fa1oyF8P1BXYG8HJoDab7Epdww0pOxKJWMmUYlf0eCmE
VZqE0B8hOzvUWNmXNKIZl/WpDD56OcclqT48DgcsYU9Ver8C65i60aSZ0CKy7blU
zKYu1X4lqPZH1uBFmkTec+ehz/b32q0YP5PPh36Rt/sV+Bjkr/veTTPtqKsP3alO
yTUsqQ5prjf4mVzX5HIq6Tf+/Sr5Y/Mn3gwqXCiCnPCEQENdX9jQnlBTqxjM1+lX
CO/uyw19ND9bt5m+WjBoXs8lLd0EcxHMy+RlNQnInbWmDBe5bwamOOa0qnyAWjUN
KzkAdJZ9h11TeIN3bzIWtjSzHyALi9ZsK7oDK5daQl9QpzljkImaF88RXDwyKdsk
w+ZfzQcsBc2ED2yrF0xdHX+SteOKZHHsQtJiT6XGz9IC2i9VH/KRjZ8njpP4TtSf
geK2j+I2HFE8mkexDE94iJCfwqxJOgmX0iGwGcHVVxUqJK8tJQ6Q+9Zp5KtUDmOd
850V31ipy10GPux1rixOffTdof2JAuKUYYFBv5FedpTYDzdeD05g29WAFeRIX3Fp
QcZ808qv9tadRLUd+gL2DEhPqDpJKiTIS73XdIWsx8VZSREp28ucXcFXmQ5RUcEm
AGL6n1Yhr7bhG8Ih0ExYOAIVYHaa0q0tKtWwmVrGtYo+K5xipWb/qNyLr16cn53M
/c3gDBySLq73V/PB02GndqUMIgW5Z5qWGxo+ktC8hNKiZoxOjJlp9MvGfWDGqUes
w97qug/a7SshNxsJZSJ7NyFcbTKtVhyRoJ/i6a4s8xuv/gO85AMQzoSVhVt1sWew
kfKtofHx/Y7xYSo/1VWQYUdTsM1MpscIJzW6C6Bg5oHHA7LSuoMC3NIKzvPCyXi6
lWZs28fS0I80HFlYCpzPdfjpH6wvqbpxNiOp3vkjrKhiHiueD8lk1AiGrZXx1OQX
f+E6PxxmVaEROiMAR0gc4/MG8SCKgDOSI/MqpbwTKqxGKpiuiGIzxmqG0i9C8hot
C3SI4XWDZT4fZuqmWOeP4dXWUk71O8ngxiHfZLvh2VWeOLtR9xa3RtAkwxq+L7zH
kp5bp0Q19gg96PuMGKc3ZTWP+oRC4x2tMhMjQkfEYSNcZ/ccn66sNKVOboWxXvrp
KK1/DLV7IfysgisIzqKvZB+Ea19DkaR6vB71pSwX+f/jsY9OF8aePYf6ydxyLT3b
7CGYA6IxAu/YXHtalN3EtmpIJtN6EgBK32BRezDg6qYtKbEGpxXequ6rbWjru0zH
zHWRECphlUSHTHYn62Q2zUdZVLbaeH2qJv+Iopll6GR1r5Cr5YchURP95OC4jSKt
LwdWU054lqDVN5GK5gUeFkDn8r6uxyVWvZzwJl6nBEDHwBn20gNXWHnD5Gibr7zq
UDA/eLvnWdIAG5Nmefq1OgOQ9uHmrU3dPYe9828CARauRdNmsKvIrsnLXvhuUXw+
gRNSuGez2B8GWq6FM0lnQpQuNgzH/KFRstfP92BFzHNAx/Sw9H43V54xvwMHIaTT
kd33dJ3agsQRtOeZ7LVhwe0zHj91fgaRhx5fThMARrCmKTVS4NR3OCJWrOLonW8s
HhPJpbw7QXKFKfEsenRotf98gZqz+mwrBJvSlblcXPWxdzsXj01pp3rd0EmexXeg
fL8Hh4NMtr9YEdKDaapxH4cea8Znj66d6u7hz3vsAFY2n57mu6UNsv2HSIembuHY
JWW+iTfa0w/+n2gpi+ayMYG//TKmGSJoYOStk31uxLKRpS27yWr6udhrKLex8nfp
4UDC9tw3/wRB+t+cNuptIiA8U0tROPX38WTGlzn/NC96EY3R/AL2/WMr/I1wUw9N
chEI2yN/wEEG/5S50kKR5x1nPKVd1xVxbnIHvw0vBmm2ab9iDuTo2gw/3lywTmPC
Hhh8iLB/T3Gr0Ruqv+oMAxT2PpbnchUHJpRJhGTJlFaGUzKzMCXV7i4HI1yAGKK5
/D4QItKHB0vLmwCnKbnDMpMtFeTsH1s1RSFSd2pjpdtWG1BAMP3MKrXlf7OoanUY
/ozrpIAvWDN/Fz0f2Z5oDt0gBZTAfn2GgYNsvkDJ1hC2uF+ZqIh9bYDxzDUUK0ta
odD3FSECWsPYO+yCyb/t4Flw/atWzawKt1VRraFIHDMTB3ROAm164cOHIwbeE2BB
LnvlFMq/f2/kYGiAL0ZbLW+Cyoy/KnSx+hKRKPc5UOB64vzzli+KBlroaa1wR7mo
wlG4iLL7uIT/F4YQ+YX2i/dxQB0nkTsQP4ycqiel/dfVXbLBVsCjYaYeCWli5Srh
++9AByqxwtLUnrvjHT3JJwsGxZ/IXC0idpI5HRV7X339b9XYH0F0rd0+hRg4i/uT
sEYGCa/mEeE/LGS9FAAq9aZ/R2uFFIefBDqD2IAul4Zv+40H9adPAV3w33YkcbG0
nAYa+KHptBboZNr9I+lEqQjGOtmqb2kcarBGT0uB4Ib0d3SubOKTv4bGuFoio17G
GXTzuxTPxATQSEO4CXPzDRJpggIeJG5FMOESthmwkrZghj+pkrvTV3YHhkplNDbt
Ix8T3TYA2X+8F1XisnV/o1kl/9QHgNDPSRjF1nzjf17KoT0UQ9zbrdqt/R4B+xEo
kMHrmccSTPz9sCy4whHzcwtnHoVGBI05FoID3mLbpPN6LGawuQ/m7UakBr2Sxgau
H2mho8dmFPNjmlXe3qkFJV7txqnWE9Qc1ZczAK+tSz+MCiwhk7xiTBq4Tu4TnWNu
TGkNdTbxwln5eZfUzuggkCpCHk7x3aGLpyNTNQmrBHQlz1qhdgKOV7Lbf1p+EGCa
8tjZ+DFILFEefksZrFKe5kCCBwxhujWiRhM3b12G3OcQkm6pGBfoBGtgmZqbyWKb
MHZ5NWQEi9lIUVD+S3Zh4Frqq2Asa7uC3+eVUaZSnmVfxRsS94dkB5Ue0J3WGkVG
qyuuH2TkvzUb348r1VZGqJxB0fgjV+9oInKR/adXIEhsTFI2YEoxo3bzVDj9Kmws
aXtGZu7V/VSlWW2a3jA4AMT2t5bP5Uh+DmFZPmV+fF41pMRY/tr2YnjPbBYhUZUF
+aJQLMpoFX/EgBBnmWgd1jElOK329EJUBLAlUk12fwzAs6EE0O9CDfji69zUGg82
p7SM5pxat9HC4MaELZ94Ly7K9Hgxko+q+hSxlOQ4Pt0VUSLyghVyeCmonvLfqD27
FBAY14D/qwKLztdDbFdJYWiy1QVb+dsq4IMDsF4oGUmEMdcDoLQumuUVYY09D1xb
rHqabf0tXY3H87NFLLvoetEEvJUIikZ2IsszYDNhcv/r0rpLVATCxFTNmm0v/2IO
pYh0ZSn6MYoCAnkPkKuMEGy3EFSE8O7L9aME+qeypxEKRMOiF4QnKcmSvelfnRf2
kPeG8Eo9B7MIxD+9eSwAwfiRxfPqQRTMIDu1LO4EIEqPNmpXfco/onZZugVzR/kV
zJ6btLxzFtwxG4A5BnxLzMKgywhH9aG0N3PzT+mamIbPtb7j/cMAD1CjFj5Ejh3a
6RNH4HSLGap/McbqmY6M2nwvzkI8h7ybz4rHfVyv3zQmoTW/BE+Cwnv1T3vJIVux
rbZBSDbuhncLJYpofM33B48zFZ4wGP8M6PeJmQbE03qp72/NL3TZXxYjdL0FBLEf
2LJmD/9R6A05nFbmo48IJLYtFgQrsifvtoiCDWT/VkG9hxu1vw4zlWODAJ7z+jfA
HX/ja/dZ5bCPt4lkcflFbGvlV7e/VIO2dwNZhe0gEyktP1TB03GVre6AgejOR9wU
M8VyRSoS/3bYbB5nc5aizSdmYZuxHh0S+mmg4VWABdfNFjTfupG/HMkGrfazxZjs
mrbm2lwgC1CzTpvKXqwqf5V+Sc4O1gsTwzNqiC9vYnV9CPfVfZurb22H/SPj7WQO
EZLd+ptOmUECQX65OobxGqMRcexuSYJu3XKUnyMc4mOmJ5Rqg8KZiq8FWNOC9nJs
I5COUkKL2IB/WluhuSZJ9mpqokzpjqmsAq9q0wJd4Iqe0tdfnz4eFj2ArNOaDbip
9h5vJQZX9yYfgAmBReB2z7SxtxrfpVwnTLyfzD3vnM8Y0txm71ZvbYlZ3i3kdgXC
sVz9LfUDEE7A/dAvqqqKGyI1K+cRfmDlNQa4JLHeA9nHB72V94NBs3YPPlay0wDn
QUIJkrNVakmui8kQCIRLaVkZ/SjQsM2bOhdaj7E4pnx//+Sld9kw0Ev5/b0S2Eoj
9hkzvT5byha1s03IdObeJeaLPCHI/sD8lxubzSYl3+M09jGXVXir/ydpAICQRhWz
z89PPI18G1UwdP8T5ox+JNsDxauRI+B3EQBCfJovoBxTjbXayZchlq4fg4ucfeNq
PLa1WhXPs3HSuUMgQwTGDVq6whySe4n+loIpIHE67FxvuEZaQxE80xG2hxCYhBqU
xw82cNPHIiSY5HdWVfoMC8LgC4LN3rXh8zW9bwRco9eHmDlyQIEfYQ9iodTnWhyY
/kSDSZHDhkR00oUMI4jIXChMal+tFe0zJp7iKnmRYVIV12XWHB/LeYxIIIakCYZ2
DfRnibVEBtvgvwzj0l5JnVAibSnmucrd7yp227X912ZATEB8zK2Tv8OZslEdkHwq
Tepwknj7ubpEdpQrXuKbNCcGFbT9YS0/Cg4GGB10pfPZqUAOEr7QeUAovQ5s+1D0
vbZKBkx5lir3FaPBHyKCfxBFgjSV25HGPV0g9JsG3cufp4qQGi86r6nRhW9a8EyQ
bFnCiXO6nXfedfYI3Ut38h0WzqJ7yO1Fd9FqE1PbHHZJfDBDVS+PKZtqnrmqopt5
RnLNfFrcC/32jY7nUeu6MsupI2Ntr6ZBp9QmRYwo5DsBqt3tOKyVJWfodmYlSsjP
ipyLYK8qFvPsJRUry3AK/yrBcHsFRxrczXC8e6tZ5UU7hsVg+78unPcOIOP19ZqE
/l4/e6P2958Cv2bjVrRms7RrrH1daa4qkEBVFdICAMOxMAJDxalfkfIG0VCFbwuF
/Qwsodz08Ibp9andUk2+fh9KH4A33l7K8YNjRd0qBf3v3naTgu0U/9LlLpjhvSdl
HgF8D5au5kZ2Uww4vVxKFh3rCi6rIGRcguMRErKogEU4UZzOX+TjeBcjRZr/SGD1
FdwI7v0iwIyhBXU5GzLuOW9C8YicmbP25rJoRuV5/7vgKaRYgpmDZkmj/DHbU5K+
cnwkBy2JAuflUE7WdnsOLS3Va6892bkZiFr6YlYOCMJAap7A6U8kHeon5FTczoPm
+NItUr8Ksql3A2iqG9M3PA+fZ4tOEbqB/aRYEWm96V7Jqeq5k3TYZlwEKYtfTsnr
XuoIeynAVhErqhE+2qtglLeKzqWst/Bz5GZQGvjguiJheOPSuO+M/W87yoxrQ3Gh
03cq6WA6OfHF5Mki7luzh8ZmGYFd8wBYR/bwICJMrp8cOqFh4esyHFQcyJbR10Ks
sq4pFImt74HBqMtP55hka4oBNV0o1kqMonbpFa1MByNUl+TuAp5nEWMXPfr7Acza
yUkTq3PcQzKNU5y6IFkvQ3WlNufIf5EqpCrYQlK8qMbFKU9TCkgc31HOXfsICWym
2nmgkm+DC2JmzdjrxqI3ahUqn94Lz/myya+6ABMLjylUYvFJDwmB8gf+A4wRbyhi
Iqf712pRAbR5Yhr4TQBO67hpMe56KpI0RcrqoBM8OTHMVO4TeReSiAgjvKjHlc8T
vQTayJ+f6enmUv4oCxdo1yCrjsYBrBCW6IDZcNtIY5ntbDB1Oxt9PLL3oRYAxEUx
QLN3mcja4rPV4UpQXdV8ykp8tY/hEhnLsMi7oXKKP7baVOSLucYSUuQBRa8tl/5l
z8nHUyRKjoRHJfSzTKgFyQIcVLJ2d1H5f1QHeC2FYsBMktTduft30/jRQNeJQb8h
6ygJ6yQ8lFId5zNAInYPAFx+ALzKFlXVw0X6X+6xFdGnElGAKMvsP9/O1/WdU+Pd
Nl5bNWCJDy2hUjzx5K+oAGCylFv1FKmO11KMVVDBCHDrKnPDkq96TafOhJg8wCj/
QvyuZwjrOw9xbzP0xmeAhLV/j+HraFgtI2+HiieU9n3pW4H5YZ1GnuUWJGxwOhEk
hhCaUhvXrr8rrXUt+dzOFhCMIzDTka519LWcoBSA+TdExFDTWZvTFaQguV53SaW4
JFdeQmQKr7Bbvft7BqEUM1R7sj0k1BSkG3vuhkVoKS9MCSt4wcFLLJxQu3csv0Oc
q7wu0fmofjPytz+S2WbURpZ9QkyWzdx4XFD02mLvFRUtl7Q87cfTi926bB5kyvzu
4tsD52HNaVdmrTlELdaZaIw3XAbZKkoGShrimnIxBL0klY0OPofv2XTxxA2HAVBK
2Qss82hY5uSZ76L/eNxA54h/xrhXYLEgJ8C9wJI5T4+shXVcW6Mp+6E5xR87SjRh
Q9saWd+bc/czyk30TjGdqk1uLksW9z0mG2PTEAHgvldEYbVkNhbR4ZNsZvWT07WE
qtPq83Xwanq5Dql2Re/VeKcgJ0k/Ki2uLwp7aN9i9mGpCZTOJDcC8svTgCsNrha2
k7p2w0b2zl706vU/Qh2LEWBp6BPXZ5JpW4MxoHkvvCqD2VLaFaTr2n/8pn/EG3DN
dVuvR4dgzQLuAdl6yv9Q7QfvH0DwS+5159zIoNIlWH/iwpxZj3J+IB1xNd+J0A2s
d2vU0TUqXbJHrrhGC7sytZluOSVTyUH1KRwAV1j1WH/Iw589jhDFdMoZ5CIZRcmQ
ZWGTGgGSTHSvQvNIJIzTQhkFxvLOGl/tb0LcFHy76Z1ADO3hplhXUNcJo/4Z3pXc
2cqA+xQpbetR4UEnWTLl/bvqWft+QJ1LYSENLNTAUkscH77n6Z3YBjWqeuF67YL8
QU8/uu9pQXSxCKuFd8+s2pOj5ZRthYH/aPG7ZWurVw9plxGq1sVl3ls0zBdi1O/N
eyyOLqB4sRonmzxvM1a6qpmYRmAy9Xe53/tFVwNEnsdgcCxuJV99vXpIO/5Q8s7W
ZTOrS3+gq76dN9xvexGBZPq9HuPk6evrKsy5Z8zi5ZciIMNm2MCZobzHuu9RHn+n
2JAlgh84IHQ3r/+WpKVLrLqEEh1T9zKwXrbMpx6sF1ts6THmg8oVGFL1o1bL+kbV
wJq+mzvfnYOsmpjXJnS1QnagWqQ+9T95dFcKOU2j000v0hXrM/cA9pmrxtXc5k1t
KH3OAILYuDPGCYOaiCESQJYf1saNhe5X0Novz6CuAA/svvqjcjRFDePtO+RR/w+M
Xvz1doD+35CCQZCQr2mRA7lSO3U/Yq3ugtSe9woSHjmizABU4EeJp1Gl3exdY4FQ
krxSSATXD9WD2finKrY0nKCUPXyBbM6rPObLGIa7aBJ9xytELle8X2+XU0m0NP4P
k6+UryHxZJ4mtzW9SXuis/S+Gwwu0j6QCixXgKQtBrbYbfWcgpFhA0fKXXAwRdJJ
SdfvGoWWuT6gseTCrMV2CrlKa0Hzj2XJgTsBHY2xSIylGkHPqts08/GjroL9/cfx
HsdvS3ZvHXqnep/kPt4LtRDb2mpw1gpZfkNc9Uo03br14bhIAKcnxzNv2yGc2ilv
LU48AkvLvSh8/LeE3BMCOVq2vNE9cD/949yOIWDjj5yr0go+zpRabGOEb6Cp9NfG
1lVEESjtmrWIFdRi967Bl2BzBDfevff9Dk6H1g8OmElh3ng8ArLmnnbOEUbnu5c8
UHDWeGUWsCEdTGmOMJ/OV7Ufkq65Lpv/WpYLS1GQnFXKk2YASWdCXa77mD/nWJ2n
fZCVrYrW0ROHH0K8iAHXdsW4tRZIG2adorll7TzfZB9NA5fCFfgWTw6f32+p1zRn
25VXZpI8vxX/MC14wbKkj4JtmDpqL9nOyIr52oNZAmjdZoFLYdtuYPQgpvTog6lL
5pDJDcqIdqU83iJ/f07jYthY5UWEWM5GaqoBR7eiQ3X4txEhWxyIxvzb7jDuqS1S
kt7GVKTw4t2nCk19IDd4oaJLnfY06Q71sTaEJI/ioKvl97WyEwcg3n94SfssXXKa
l3FF8JcdJ/zXHd3Ft/BWIJNfZtJ9NJAv9KnLNSA9CGhJCOh0nsc38/SHGsd9AIxg
OMfYATaQ6Hn850UAMaMirz683LfctcuUEkSLfL+LwCgzVnKDl4vymVGKTEVcpzDn
wApkEvsSh1ju2DNoKN2cBG+DfXJjJA4hL7ReQkx7hmvMtp/PoLekld2cSmBJ3FXb
gIlL+bTPiiJRkPObz00T8dG/SWCB+X+6uoKiM9bovZy+8Gt/ViG0JTGx8bZGLNmc
M3ZxvoMYCOfzC2CL9B/8LzQTmRuq/qUk/+aqVYvNApyoHxi2BZbO228cX6u/WMNN
ZE8mLWGi2NwHUvub/2QQBQnvF2fTpJwPvtGS/GGjcjXyc0DQDEwrvwsBprBJeoWA
yJVqXHe3gQ+5vu3BDKjwPzqMj1cAru4pIfN3IAskYRbOncHBQjFuG5ahHf33mF0Y
6lOpyxb2g1FxRmYhBihGyh0zQ4aveg7EtFLr1JpU9P5n16PftrGrhxcKlXg4FmY4
8H8FG0NSVjKVhUCfHHzvJ2pRg7TcxJrIdJthp61GnDFq0Qwqj1R7SQR2Q6MaAEjm
soPty8PyJjwmw7kUMo6ZXm+LjDzva8ps7TuiIWAJ3qnzW4wUJEjw0wu7k7QXyaEL
Zd71iLnAOLj1ObhHg+9v2pTnpskbfVQYsT1jM4SU75/IK1xGvC4CJIaMowkp4SnI
1oOoDwR8i9qD/RF6euxMiDhz3hxvSDsyR8GEZ5F1mJpqI2D8IbmqF9cikJRkcDEX
FmcgkdSZ9s2eGQ8A8hqMAuH+pwBS1eCqoN9RRmaHGFUJwVrRKbtFsRmtDGL+nIV6
QKI84oHVQA4A4C7bfu7GExLUOVs2d5IcW0clrV+Yp5+ATRRQ0YbAWUtpzubkrpzI
LEKp6N67Zb5Rt9gGMu/bO5K1NW/27ULHCSVz2OtrYrKelSI6wJMwKs+FgT9EVSUC
EIdiMIJLZaTXJRwqfU9uHAcdpJ9Ng/6xdoiaAB449XgmPMPACYWl81I4ueH+DAT2
mDDK6UkfXABk/wszKLkXIfqNOqTUH1m26iISHdeoCepPBLEJz4t97I9g1yEDxQcm
XFiLbipLco/OBPB4P7eJvzY5mvzSstiGm8+yjXokhtKriCAyfUM6zt2q6moxRqiQ
Bojm7gksij0aQV4QPRQc1tPGiyC7W6h+jtGINocDvZCYEJ8PSdoV5iwGIlmQjHdL
i3dMaevc5sfxrPBY10iDDZ9CjuvEHZMnrTavLbAq0uRv6Sl2fYxgk/9dl5O+znrE
ZFBF6FvdhOkiwBoaMXrxys6jVxGb10Ihl39rCG5CjU9kEa1OeQG9XvJPNyiKXsZO
EXEvd9csep4xSDyY9CsTy3eKrb0HP3BM0nzKFHmUwwONCuHsgcMdgIgD72Lxxy9+
Tr65urVmGLVpcIWX3mO6yWMrgNQ+ZmRx0kI58obCOQHoxT6WVNa25ZaTQtu9wNQ0
unkEOV1Am6bELhJ1ayuhPq9C18Hw3J3iiUNzoTtSBiA51vMPt7QAMvObq+axqpur
PupONFzx1qtzbcBrdi/iTJT6Ew7Y6I/j2ISEsqDaus8kkT8q3xhk9M08knH+pNh9
y+/VlmCN75NpYfzop4so51ybZncr027bYZ0Hip60YOzuhPw19n0MegWiMpfNPoCw
7Ra0OFx5BV+gMpyOLlFTDItqFSWn4TwBJ47pxWALPgG/ZcNlk+E6Q7JB8CF/iw9h
DhNkbxcqPjtmfi5Jps1GXM/xGvqTLQxGj6QzZoUwg24UcrJ+9R2UosHZ/XJ6fkhf
57u3d+Chqq8/bBMJ1anxl8SrGuEOswSMoQH8wF6ThPR00uLDGSBxBVuJTbMGOYm5
lpYl3taeCVAmbR91lMP7UuditXV7CRSxYoLgN8FPfaKnubkGJIouC4Cnd2Mh0Rl3
29jsN3hXeQloZUHuE9rSn+PpnfBA2VTWisktajDUI0v427yzJmhcnj3HT0eeZLXu
clHrP4qxMRvjqyVcaXfdq5b4fd0bHIB72UifXGHkTVXDqeOUhu3lvz7VA0ai0eDP
zRj8AmyZreGht07Nn6GxatWjUqw/Hs0cam9++noMJddK1yVvuGkMcPB302v4P0aT
SaDCyJ9vufnfB7WsYNt/u3ChGQEzsjLR75rNqC2DAOOkfjuqXvMH++gak2wFG9Qt
lcEMi3CVEsV+1bMAMsN5g1ABSOB87RXU9yODpgFDmF4o5b2Mmm3DOAFmjFu19v9D
0qNDXgsAxMFbZw+G5qaTeYbSYhXi0KF24XUpfIMcyfuwPf4E6131ui7SldGzIQbi
S04TJEjJHpqPe7isuIUQZMkPL5bgKf6g7vnHpA02sfPijMmAm0CzrkqMmQjM8kxG
h7d48zX/bB/BWv0LJfsE0FA3aTMeF7JGquaC3XCuXycRtEa4RlNUncyIZFh8BH8k
NM9P7aE97+iCuPpHJrIKCXLrl3y0ncfzG4APM8XHBHndKPes8QV81M2SqNmBjUl5
Ej/2hrAiNY7WpdJoggxpApMmlMx6xFnA/G4RHRJHjZ0sdvQ9DflfJLnvIndNB4q3
CP0cFP8PaghNrcru4Djo7vopZYtGOUcmd3OhLQCOQ5567lBvL6fxRak6lLkDvEWk
qh7zepj+sB44Z1B+U+thB5mRNKiumht4G3qf3sR/VOb/ZftwT5oxmEc86tVtdznV
y+fj7DkNyHwZgbYZLX6075css1Qw0SNQby4bcNbTuMitmWWNWcDQ6tvRl14x79te
Urgb3iR0pjQ5+5TLc21sexI63y6GHQhd+g3UeU64QV1eDav89TWMdibnuUJOA9jn
S7FEjT97pW7ohvDRwz1gd+k3mO7VA5ZB6abrOSVrVVOJenxUU5dcV4rVBjD4/cR5
vOiPPypzHy950q9wz3sc6jBN+BwUbxXhkIXKFGnq6q2IqxmehAi3zSklYUfN7bqn
s3vj1XPbe7MLOUJptxdUo4KWdVmP/GIIMk17Ai7BumYbJgfo1cYaBlOvDrKAjqKj
FtTbxcP45JJAeOppDtotlZUoyIxqR6F2ZC/zu9iMR5AahG+nHVvMIrdOimKnVczd
X3jq7NJpBTEp1pH4yutrk7n+U4dehvUkNMQ6abX42l2BKT3SgxdlK4zqp3qRDbXm
eI+s6q6Hs4/Vg08d54dPbgje2CiUkTHyy49zlk2dGEzdxyubwLIfQ86SJhq9Splc
ZKiu1wJYvX3K5Z+Jr1ivs1tArqTtHmOc8AvgEpkEgpAZklLfEY6z2OATUPVK8ASt
fS1s1odio0gTtZs5LuZAnUoBRZGNioyYw89yw8wdbu9FQyUL5Wp1rsil5V/lJtWX
vqkuWYPd4gPj9ab9wZwD/FtDoPN4aLBIrbkN00SN+QOznYOSGAzcBPVTF/55Eldy
0O1jcv7sSKgTzD2U+aCGwZvafWGnCC6Il43+5lEnVae9ofLIiJ20Yo59Ft2BZW5a
ofNeSqoDH13Es56QCBwVzv7p2mZD2w3xa+ysNQKmLV6aoigUOqXrx8SlqSkIrmrt
vWixIO1tqnoGnsPUZswrPbIRxN+qIpzJ2N4Hof2+hVlViWvOiy1HcLzSohcecJ1q
p8UuRj3WV2VUwLsdXrk3cAHtLV7fjDcttydxt2rtd3FKr3CY+k+ENa3tgom8P5l3
MNKPGmmLZw8JQIe6wTtSrgk96g4L9frn0KhJKHHnzXRFAQZQdXDGs0IP7VgrEov9
OUNZusmNdi/gqnJmrbd+KqG/eoyR2o3uoBrjZPm96IquqBPJEjv8AtjbshFlrHPG
RqYj/odRljWbOH4v6++5ikEPENGBWRLVs4E9sXpiduCO37VdOWu0xO0F7mLbDyOr
jsALMfvhcBwoNo7cN1VfBqCbPjJA/ZS70gJeYuHeLL76lSqc6xdsZz+Y7Zb+CJ3E
VrbRt65cl7Y4juFki8yMYG+1HoSh42vH/Ws0wkWul42XnaX/hbNA21m69L6r2ict
oGgFdCFQGPaVux17O6w099IUmkVFBQqn67aPwnEFeTXdfQrlLAg2OstugD/S5MDQ
Pg1IhEsMf0PvF3TjNvCjbjy7AbD9BMI1GmCxs3HCekcqnmoD8t7o/XdpKQ2RZug+
HkMZziFDIAUuz/WxZXS82zqU5lXaD9MRjuPIv0/FuSyyrJxsPnZnR9nAcq4WxsDn
1rZMc10Amt6NoWhV0zyyqx3Yuo5jM/26q6cRfIC/K/7rCN/QVOItdNh5VJfICLux
ZqmV9dUI3V+hdWZdvwrgzYTxOVwoKLo749/FZ2Ycvrfpfflrgx3zf8q11vaa0vG9
XywFQrcLTIEwRmHczIqj5M8Dpn1FQMhitvDgUD2rXFyJg2Mir7TbxeMTVwaoKrIz
cg0cotcEJkrSkvDQoyMhyqK0iwQd4wVynSHPFPmwDp/ptfgCwoneMdJjO2CHmQ/6
sGyJgdfrSgUJClF2M6gPiXqmDEDDsS93QxY7TOoIAKan1gee8Hs0DOhyRabX5Y/3
5CZzcOmsJvTP2q1zLW8ZdG9Gzv4TU/ycdJUxkSazHX74/dKmAbdg7h0lWV5SrgfY
nyfpZA/gS7y8w/GOc7aZhmNkx3BNcXJo7t41NGwHTpl1pEcLHK2ZLp7RUJkjlSMA
17mKn4bS7HM55PRzItykspWpkIAwhLWdd9B6AcrqLo2YMwbiYXTzSlmkLRjqibRc
dGxg1zt/GHXHnbiNpe9nFL04FHVlwDoRzxf3sz1NKyOQK8i6yF3JMDC8Kdw+sfG8
af78nS8GE/p4BnCCsPIca/Yj40Qk/VB3ji/wkAjZ3T4fNAYOw+XsW1pZai7PUqMI
gq/e3co8RBTk4J47R5vzPNf+kZsVeL2q59giC1mCGEDkshJbI4A71mXIHzJy2L+B
Dsi7HRwQb0kKPTf4rI/xCDzR8yomomo6+zJVU87ZnWTRbW6G9jrSrv9H85/+Qnc/
l+2o/55vw1eShxwUILfM1NPlPHxaM4Lr2qSXlr+/kKKPAdNpsKzz+eP++oO2uicp
jaT4I18ctJARV2SLzfu1rhC7+feGNawWvrRtfBtyd5J2XxQOtfeRgv2Ia5YakSIC
7ghzLWobB9fw+8Zemdb7WJcJWvh3jUcrbnxLU8zbBQVD4puslmQkZWNW3eAZ70kg
4h43KIOtmX1BWT9qGmbjhN0tVY9P9Zw45D+79/uJyeZUrcJcFym51+7i+Ue70sni
a7fQCDstbQQEPo6XjHjy3y5iIAu9TXzZ70MXuC3AK5W6UORBz5OXOUv+xB96la35
q2vWzRaYsGnfeVKiYQPQyQJ1qhLjISN9k/EUY9AlNc7HYOVLGDKA2Nyy3oI2K1RM
5KXeSumfw5AnTHur9qBLvUIB1RMUqeh9cXDLuEGG4fQ7NEecvI8yeFqBtC9D/XX5
27I9hb9y5MDefOR5JiRbt8t713k7NmuNohpmxeUntCvTe8QH288v5IktiklA+3bJ
4IlPIbiyZkDIp4jHZb0Vl//9dmHileiYgDrNd8j05sgrKHVD7bWvjUYLMOzQ2B15
epIhwj8FwwppWs0AnUoNiX2Fhy5ldfyrhgvVjpS+BXKAv3JBWP7Ebc3w8WlWJa90
0L3BbLIA6qn8smNEnMB1DBHNyOcdMQZdu4ABMlI48p0TkiASB1Ls6D5T91e4hhLj
+40Vg/T+mDohnDkl3Lps19/fGYGV1ykIBhBBNAQeBRYnsI04Aj7LNPJDa1pwsDzI
N9JwupB8Q4aqU7+wqGZ5Qbe5kZDqW/nnjXCMvIe00/h3V6s1KNYn3DatZcbAYaHV
BwSKxXeHn9/BfJZYgCD55C4NISoSBssj0mRkHYC7nqQLZho3WYnD5VqSW6qVV9KR
+5pfplmDvz5Q4F90JmeMLroV2MrpVDVesNpjELDUqQdmn4yEYVxnjduFkiHqD/MP
lMW+w4uIF5Km/BK7kJ+fqdpJ8Clpj3ftbuQyX9gu76JWzAZ+QqONLLiEud3pEaQs
PTO9tmpq9NJ4gHSoVPsiw/nz7FMIx2z6FOjRnkJtHYbeeqrDyi4tale/q+JAT2cw
tVcw5IPiAyd05RF4PLgi7bQImndMPVRNnKrilrLpNWYrT8tlHiPk3o8f5wXhBCSx
zK1sztubajOVX9DxxywbHx0pYfw4xdxu58xjEOj5S+7jHgw799cY7jg6eVAxY++1
qqOOKNG+QB4oUww/qxB9eKK1MPIqkBZpV1SaE8W2DbxUUwDERmNYFoXvPA2ejRLB
4fP2E6GKA1JCx590/dm6cndmQA3qQdHfICte8WoZrhbqr/9aJcGDZx5WrRy1HZf1
RXpY8bC/+H22t8njROjUw3lDSRXA1o6RTWDcTfhOYnrR2Dz9wjlOjwHXeuN070AD
0JWwFceVr5EaGXJxS/xRn93fIoStLKZSlnKVj4XvfJ9VtiYc898il0Gfr6ApWN1T
WYsYzBYsAVoJCMcogFtXhmHsRYtMgYK91tKhQAzT26hEGfGTNcqaagnfWzktsF9m
QzUBghavi4vRTi6csPj9xEj/j6ytzKbdY8yg4Aix/DyPLtxXwhdo6rw5az8AzE6D
z2+WNrSUJuQPL9Ac6PHsC1bj5dtr9i4ca1E0BiYDq8+qC0m/SsOxqOPUu3IXgWEM
x0KDXzTrDstBbI5eV2mkPCtla2hLiKJNVgtigkj0MKQicLa2gA5gymRhN3KOrQU+
Qa/JZgHAWYVCbQqPOobwmbAKcBDxNC80XHBXnYetDZW8ACAnLj7IsqeN2N/ckPp1
nA8tH4yWkLDQ9vXfuou9/RzRrfUrzhikYs9alu/woKRekqk679fhKsVNq3aydgnN
ZPr33wvF0tr2EL/FjTiN6gqc0DKNaeHUHUbMQNfJsGdBSD5LRmTAv7GXFqlL2ALm
iPcXrEieYaJhx+uLK7EYsQKpfcp+jNiZR7Bjo525fyF4Bc20AWiIur0g20h2sYxw
ddJ/3nM7YwNliTKM21mYm7CxRfh+idiwY4b3tFVaq+wdv7tz4mGcj/FZiES9xGFC
10geOhrvZ2+IeEdooTrfjcgzY0Vy+4q12h4FFey/omQvN4MVzBzT42K4IXINsafl
kZG3X116ra8Tu8iK2X69kUcR0HowxE+7xVZDSAiH46nNmneH7rFbCArAUeK4O9wH
2EpItW2JDphvDp/FbX6Hky9S17St28f4Aq5cKPnp0EDjN24YxD1sruvX5RI4jDZc
zUuF8uulc0EZJk93ds3aa9IABcksAVbmPLxcpYYjxEu6ugWPyJxXEajXi5fqlu6w
S3WeGE8BMEhobbVvl4gBTXU0sUwRpcASVTK7JSPr6m6UhiqWmFerRBmwlHnXZ1Uw
ReaivDIn9I0LTNgxQtlw0M3GnA/iDejVewwmPhVwtvX539XMd+u1MD6/DWLi/Rpg
7K51AjBZFAavhom5n76P2MpuiuACm621pwV2AzGjz9TSVbSV2rBt9Vc05x/JrluM
W8kjy4FvGT8obftKS/avZ/Nh/ubC6jEpgumNBJfgXXT9k1z1eQh5dJE4f1K8N0Td
7HjMRjqtFBPlF0bhNnjvg0QR5eTAsD8AvZBX1Wcf6fXl0ZhzQxXQLdWrYt2REYZZ
GEXy3VfgUmpPKDjQvvW/woDTBxJDHg5iZw3oREFMwFuIHafbSvqq5QgaDU2B3FwH
z83LZMnbDDEKxbjkLYHfFyC4rRwz8VRL2ezc9J14jA1UKax/H+6y/gbaCKOaAf40
/DOENL0Bvk/LFL2wxGXFHzrJpeeb0QOkivL69gXLQP66ne6Y9bUvsT/EiEsf5zAg
Lu0EwpQFWc6iO1rx3bCNL5pN4AHK8CMk4cw5m14qeLAscDaUSkp1mGk/jcg4OeV6
FxS/ZL7Vx2BbczsbxpJ8hpLaSOP4tI32IV6DB0PA03jhnhqtHQ0EQUCSrVBo6reL
Es2VSbpQrnpzPxOxqkFxHAgpvzI3oabU7kiPtYelGlq/9my2hT+Bi1yvZxqaxZ5c
7AsVIp7xIZUz0bcN93bI6vSWlOcCDMpSwYsaPF+qLg14hX87Kh5SKaWRbUE/hCLb
XPztVRt0lS9n8qzJc9zYq0Nwyi+rccMxrajsBVfWIglPbF24LcfQxCBuQEQ0/W4R
CJWvivsRJAmN8TvEYq60mtviBRBYdx6yxrA69Msnilfhj7rj3UWmZzk5pDCTS39C
/aMe1MG6kQI+FZkGHaS/hX0gTdaEi4XkbW4j+67Y3jqqTzSL4yWVilL33qBD1sYy
pKYbzf0q+p+4pG1zR1cjDROrRIQm/3kZjDAcM7MSPNSGaMqiQSvGdpHVRxv9Zjhm
hmcPGXepwXkk0E4tBmcZwEBlzgp/k/GILT/AcHGXh85ixY4UfYMbgKBnTcq/vl7u
77xOUT1nnjgmebHhESddHF38vrYOa63Sivz47RDl7qqkuoQtAPPriNPfyxY0r36x
9y5TVb4g60jLle54NZa8wI3ht+Z5oeNsnKJYMw91n/zQLCU7TEmoEKmQ5d6rceqV
mroun4/65CVhwewrlGYJu8VYRXbwJmh8QYqog6+6Aqceld2/JQqvNIrijUGurZNK
tO/jlJ4/jo5oSaSHqHtLRv9D9x9/U19qAtdz/XoDUQc/H0FR4CAYAgSd1LpVRhTs
m9SzVpCneppgqfphV4aw/kKzxj20CT8/6GxeyXejnMG+WwvVXQ3mZOCzeNKaMCho
nZ5fTKyOnBdOIHuJe1T/sES5j0lhF2xp/jkwWA6gMmSKhHpa7hl/EgD6ImMOjtqr
UGymiK71rvlLXq8M7VzsArYqwrCRrIHdJ2RFDLpbsTpIRWEjawt9xmCu8RFxN4jf
ZmHFgS3qjL39IMpkaIrbuIfelWPNQ2aVNPK1qcCV5rrODmtE1u5ug05Ukp6U+e9J
aWwquqD+Bn8OOabf0I5/uaH8Sr8toPS9p+B+3PMyPjiyBizHgapbg3H9aoCGPGiS
TJJEt82UekISnHhJWwidmcWLMmoCu1inlK2HIv7KdfOMykC9ru6/vSshkuqGDAYA
6D4Odue9qQxFXYHHAK0D0vuiLSRwPwuWMrKzsouQgOCyty/cKsupjf4OntpFb+6w
WAqZioci0wizJwhJ5eTHoZY5LVDaCF7B35F6kdGEWLAovUsHBmRw2K7AJnPt+7FX
2BI94pD6BtJuBXmzAxKbX2cET7W4+/IC6yY9CHgALstikA6p0ezeFwPo13JyRZza
pu4J2nzEWMuirnb5OTx4I3XJ3Kd7XWQKEfeXuNxCbLpSx2v0AD30WrYU7+WPk6gm
3e31+kPXgTcYUK0Bd5swHYHZqOH3u3dDuN3M4Ebe9Ed/T1+Mwcf+FHCDbbWJO6o3
0NKQoM4/xRqzQKA7Vjz7I+AfmBwzL3t3qwebqoYitg1XgFWcRE36E8cRNHK51UVa
tixOxdLib0HfWV4D0cBQPPwbsrt752+kvPavtd79p1s/O1A9ZJE/G98/LGsBWxll
DXIhbPhi+Pc/WGXOLz1ZoZHscUpxGz1Oazgcg5K0YAZDlda+Guk4aVAIQhrFSXP5
m4OPlGkSY3jj2HBgdsyCRXA0ZYkzej7jwD7dOygmyG7GBzYmr+1iBtZUYffMTBQB
qSPsS+7d5LoIWl37ZMlpL4ueBQv+a3hnRnd7vIRR/3L7C4gCtxLtFO7uifyegMC0
95ZyKaOR302fAuxAXNiSIut6WQyRrPZ8wJd2MrudYeOYsGYO82nw5/zb6/eV/KmL
qt4wfJ1bPKojcix7obgH5P1c7drmJxM74HA04fa818J+Vl44FxMY/f1owl33OuH/
zXl6uVNfccRBuYEXQVou7aeEWDw5bgNnkThyVu01BV+LMf3qMFsVHGnq+Dy1xJXI
ZfInvF9B2PqfD4L1CvX218UEHQGJdQlDg+40jDkLUeDR1IKlYWZjvg9hy2SUDcBS
J89HtXhE0zBMjdhWNZgMT5iG47thVMZWinS1EhL0SykWtlNEXawULUZWjXyIkWIf
468UI2hW5c0SMhHeF4+xl511wP7abYfX1KvLLLzwruUPAeZ0wgRE9lmXNuw4kObq
u/9Qb8s/a1BAn/uGn02Z8G50BgXrGk5MObqGAFHBvxaL39vOpR2UHkiBaiKOJdLC
sEy5CIPyeV+loovfjAgqmjwZRwXx2j1/2Y6pNr4zMZWJk9N7D1fyVsqz5sJJlxIK
EGxr0JJa6L+zsvKl8bhxUu3zOJDhty2Qswwr/jtcnNEc5lOsjsC8nquClGpC2gNj
R1sCCpGLdxbpYHBFZsil0hcYcPcoy92mMibrHYjaKt31XETIM3RgEnvnB/1kuUyQ
xn1QU94cPo+HJ6Q2QgAVHGX4FtbU/CHKJsvYnbjU6KVLPIABQZIQ04yGbHqU+MOb
7kmoLdlqd+jGOChbhQ8meiWYP9xII0U5K6O+NFgkhaqhXBdg/S83PiLeb+is6ff4
CrgUEz9CzIb8M5QTyQ4XbG24UGcQQ/0Gh0LkYhw5IzOgc5kmPI/4T3qBN/po98pE
S/4ef8nq+xf8nHrm4R7u1BmVMjZ6TKy7kSufhpShzqEHK7ayKPDlKCUcGcZA6rcD
Ys5WD6YppsCF70KRzktGZEAGypKVaN4YWrUoAiPQ7A6183PPYjD912NvW4X4ZN2o
isOlqcsfn2CBKYJVS6NCbEiXqDjJQHAFa/D5ZwRq9ODfP8Q2byqe8+Uga1SkNUgC
Mq7RzlAjyCcum/wkF+nmRcykyysIrVDd0qDPDa2sgcXBQkLDpMpDvp9GzWbD9bxs
j2bjeMafzV34g7TeH9pORcit1PEzYqmOt7R0TkcWWJWPYDlAsqr9P2Sxd4kpDPxY
/0fnHma8zxGx+QBtJBcqWgNOgKfQF+uUscsJXPQKo5I47rVi3cPXdmpDl4Thwy3P
Sh/bY5n3daGyUArKZEdR0aDPQdPeBTuhztgYUK97VgT/8MnnvCQus+6ZRTvPjQBT
0WwNSJPnMjACbQ4jv4dLWV1BMhPcd3cmwn6GTusZWmVs7L8rplY8XNiOwsyp3dL/
qjupkbUUja+4uIQSq+FGz+yV8P8rnTxmzcUX59nkhOXLn6avabsxbjGv6R6tfU0F
ks6KBFSci/2VAZN+addzKw1ToOF3PZ5AyGweAzwQLfxWbALiOmSzXrgVfWKxktWI
TkBHwhVewNPq38q2b3o1s79Jqa0SYqXLNdabHnang/wzFUnxBjBI6YROOyoLMA3R
aWidZfdaQZBkz19mCcaxDYeCpAPoh3kZwalzL+AsWuRIjEW3oRc6zEztChUeAPAr
kSWyphpqM0bShYPOUtBHhx3MvwS8lvUE1BRCKVmC2ZudJt6gtW7Yf2l/Ro0DocqR
qC/8dutX+EyL1L3kXXPhyEcvbgOxHuvhm08vbXeuCSQPIIVtzYy+KEYsvf1+vS8d
EpykWNk6GjLYecbLasbtebMrShcB24Ej2HS+SpbxyCjNn8BBS8YUu9eYNHoMZfyq
j72H+dx3WuoUKPK1VKtxTVQ+5EB2i6DJufT4RiKu1FsYrrpnsUuKD8jRek+jaARV
cSSBWfT5KyEm3XVFhYCFreE4WjdADVXaXeJeCfHsGVpkhrcdol0/vfMLMoHCyEwz
3KFRCi1C5AFtnCVbVIDPOdJuYPSi3zmXQ4lNvXSzr90gTmPerSzEwhE7TMQAKVOd
oXP3rW5BSuJ3UNw3Z64IZ4+y88g5eC9ToVDHtmxCj4N4TQWLzv2bkrWJZp4P/bdv
WrP1x9cezb0GjO3tGX+BVKhr4DL/6UyLCeRTS8Tlr6T3WsjOUfLmLjznnZ3xqqzG
9s6lJMWHF/jOhhqHSXYgKQz7DWRWSjJMGjWpfh4X28zfmbjxxRE0omK/oZBHPmTL
zZy2TAoeShLvjUzPOlzFMxfEtXSGCWaFGh5Gfz93O0geukLqzBrGDbnMhlarT1gT
+cjLcMhwA3g9CDCx59ibnNdNyPQIMFpeVWxqflM/0eCELFYm6oaa+Afrw0ukzt1n
Qk4cwvwEhbPSdjQdl1S2bw4HFBqkXeTycQSdk/agq0Cf3k93AuX6bvCBDkjkbfDb
2U5KjaMzdF/H4PCo3b3ZxN144jMrHb7uL+eUOb2KdDYgNpd/M5IApY6ENdFyG9Eo
y7jatT7ztAlkAHolvQD4tzOfS8BcPnzJFp4yT+8Bpzq3mE1e/duEbZIdyJpad2ot
n9n+6GGge3qW+5ssJCKL4EyXYsDlZuidkURAqBL7lKVFD6L3sQmFKmx8nC2vs/Sl
YZZWl9hV8Lejq6sDjTr19/O+CsHBSykKnOC+JgLOuqnUdXHMKXoLzc5Z0sn7o1Ed
p/uRn9427vLHywPpdtwoKLAf5DcH91+G4Qhov1tUVzA5SMAW9dohTcsTC1qmNC2v
qN/Sy/xMH9Lc7jOrTUZdZ5gcz/klInoUZNjGpXCKyfr3xSAnp9CFJknZ6/EtQWRC
Z30tVsPFCOyuh4XVh3FR5NiczApPzJUKkm+aPkRgVVlgyrYhihmCBQKLHkQWwqcK
HM0RLjQB26NjJULMYsQFl2KQVEosGN76c4wvBrvomS05BT+1WSSEtpRSmuWY0Tsq
xFdGAucs5/9fEMUc1EktkFIUrcuSfNzUbemRBpK1WYIZPDQd+aFsk2Ly9uWP8ncg
u3Zp7bNn54FhOotdtuwmTCv+vysz8Ew2GY+2FzfYAdxYWXJZtqhM6fZnmC6Z9y2A
1em5CEqX9vxt5qmrP3/xutBDEu7URTjh+cr1PBKGeVdr6Ejk/hCmq7PQhq3cwHik
qjZRYRjgHsPftRWNQBjKfmg0Ijyh4w706xGy5X+idBV/nGxo5EluB4WM2RFCojQg
jfbu3oS+kbn/C3bTZembB2VzXB1a+dOvhmExNSpWofmBD27cCCXgF51hSAwrx8R1
qsEYyMtJvuICpA64ZP7UUxi8jRZ1QR83EIo5ul85cbAZXh/ZkG/tTDoyfptV3mzQ
c41yOOI0MhNl43HSucFHOgo0UAE9ZRaQKZfPYZbHAgKYcf+XkJhAiCxpQXqwmpB6
1/RpknKQIdVycwFmjSTpLeXewK3BGywsg1P08L6qc8nW8EgEkaGKu6BfcFUvCJpM
b/BhcY49hWX9KZA7EOYARq/IrkrarGkf71I7QVX3k369h0gpv8WssRsUmKrC0XwH
H4GI8dgt8zTqV9rNN7A9qOdPmyl4ZfpuhApY10nueG8XfBw9PLRoTYk6n72dOh0J
FbqNqT2cxklGR/Jc7oNegzFlEKyQ0vYwdAYBEDUpIytQ8ZxQiTdRCqNQNJW+6d0I
vf/mAWlqsxRiFoWvkXzjnWY4Tvu0sp42vGLR9YIYscKC/nM2MvX1cs0djCJ4dZRw
F2TmjUKBKX5fULpSBRsYIcr6UT16asXnUUJrkmq7+sXGiZzBsVAVxw0Htr9t97Me
WEwKH7SJcUyzqKJyZ81neAcBAwuqrHKoe3CjLgEHJkJuPa5GX8unNLognbawTNEu
UID3SbfyU7jUclYYRr+xi3pm5eCibFyChGeF6KVzXEdm8cUXF30APDXyoAwa5akZ
J2UYGj+PRTHo5jYMFBHBQf9qKcT+A138CtHJDWg0A9gG9mJPG8GaL7Bn0y5c/sNZ
cyn1T+vcxaKhQ2jHln/zAVxl6bnQrBAv81pXd/RNtswK5J8n1a+aFkKvdNFVqhrV
ML5dVdtJ4T6tbIpo3nEOnfj8J7qzvd3I1HzaJ1w16uYTsMHdF1RgUBPoR/TbtK18
P4CfFnxsDMCsaRQlNuP5qthYJH7tchHeZHdpQQrHYuvHbd+4uMQols9oeJTNWRIb
Ea9EOy4j4UXwh+aXVu4WIvML2WTG3TOMBC6yz0QJ8TZr5aq7E6XZdAVcTKlzd/jU
bpf23xRao8nWiKi5DE6PECve3xiOiGL33G5r1atPjANBaL4qMHTCF45plLqc9fQD
mGpqa+4aW73/f/6qHKCxMvys9eNFXb0tnVGJ199lqNUChkFa/T6y8cyuk0/7+uDb
fqvRbLC6Tb6/VqHdzex52Gry75aWBOjRuHq3J0sBZN+2FSIPsbXpUtkaPbr1CV2v
7eCGRMUob6G2GmUD7kMAYfsLPbmnZhC03SaM6ttKtg1YiTfhUCITpVsHfInjJFlO
3ghpJAGrYGo0r3GnlwyY7qYUAoZ2x62HLXbLmjJpZawbgShrNsrpDLirnvc5ksAH
lr8e+nHb+C7oc/Irt0W2iEiQSuzfYaObWDiHeb/bQAkcuweZriTfSeIb9pAuUkOK
QJUTf+d4xq4SN3+0gE7oMTfoXnO8MzziA6k9tPgnWNSY/LOdlhAfXLLR7GbQC+VK
IbilTZoNv5R+rxsJ4tnNN+C5VrjFZcBkn/jabNjoX6ryKVxo9X3tmgbVnWBMN4XN
4pK4OxlUxxMzUXrrT8z1Mo/XLejqrYEp8+b/GvPBtP6SF96ESCEixfK7JpIpvZ0v
IaGKyXPYCsYJS9BMsO4d3J0VKDLZXY7exkwBswRQLbfjlXVxZ9Yy+bdJgWh0BZzO
SE3AHVqRi0Kwnzl+1d2idq4usIzjyBR3X4FRckDEK/dUzjO/CZRynos1EMAgnaC8
Ncr8/WSS7VcOg5DfdJVPW4O+9W8mt2UX0xiChyPfXzfO+4G7PW9EuPyTU8i37Aof
bOnO71qI4psMiFXhXH6+a/x5CgZw6AmfDgCWS98C+o1ftqP1Jqw5CRL+YerUU1Pv
GzIXwA8b060R9Gv6qxrh8unj5MqnTRZRf1RtWP2iQyRj4JoLUGYpxz/OLgLbJ9La
CeOf1WIGDrYODHyxbaUJoMn1sD5utvLIWlnuQHVnyQTq+QupPEce0KKv+/qUhm1i
p+jyC/+hOu2kpyHTgrT4SldgXiViOYC+lM/9dNfZZ+uiuYqGt6f0rA5ObhMjKnYQ
Ni6bWy00QE1TGUj98kbNPLV8IWAUYTtq/cxOuWXYu/uXsA4U2gIj1dGhmrkjbEiO
Az/TSi1yYyzvWfHtmQd5xrKhhKAzIJ8tSCivLCeDfrNBD+rGxgczB6A1L9v0tCEb
ouf2NDBYNQIyJWbtwCwkCr6SJc3LUq65rECLoc+/R+cjQiEaFnqKuMlQt1mJOVmZ
MV19EUKv7G6I8kjfAY/yS4GhDfL68isHADId5hKtbnG3u/n2Ij6DMuuwMeWAlnMl
1O/jCjS8bdbykZCiGYBriRgi6XSqc4rYHjXdlzJUyyzXjDBY2v79wZE/pd7xq4Mq
iCGSXulrY30Pl/ndYMEfE2vExNZNyFhA1ltQJsObkAaDzxLOQZ640Si17Knxx1aZ
Enunc1iakdHP+mxrf38FVSd1bgW41/KAw0KmxZlXXh2pZ2UBG368bPk9emzs1f3w
yja3QmMb43JJherCTfiz/IuJRqtXs5RtOHhtZFK5NflJ2U8CKlWtqKi1P6foMXfK
yNSCH908TKC/J5vSM3VF3NBIdeYh5GXSJdiYZRAeqF2L6VI80wwjml4c6VeK3pnz
QtNgNGT9vo+vgUSAJZ2KpYxJsYSZpEwtmfhObMIPW7YFd/37IZUcYNQ3WBgqyaGc
gv62emDmD74r5r/J/9onTZXi15BriLHXkiYtkJz2QDkc7hIZri7FpSzuqMCItxxw
2yo7XPB/wxYmTm99onD5iqXpqFnQc5bzVbIsxptty12BucTLntJ4Erx6uGCZxfpQ
bfesTueDTN8sDsPfAf3CjPQ6mZUEf+wxL6lbkcVf2kgEsMbjkeXsgVcYoM1HWdSS
63S2vtvzjkmwFVyMXmFD/SFAeMnvXXoLDLmimDmupu27ghpTaDOZdkOEd/Z/jW+6
/DtqmL+xcI35+frt/x8g7+GoLAJOsP86/l6E/86pXh/xz2O2wr2hCskj6DgOURUW
tJIDbsz1yiEUht8L4D5r5oZ5vfpJNFkykwpOsS0/8799YAXLjm6EI0BoElvfp091
hD4Ya+nckjaSVsMvxr4dnw9nkqgrnrml2LXr76qRLGJA8G7p8h54EubmPwtjTQho
8ou+MrltWjSsHueeITIQJbimP3V8KROz5ecdd8ewAokbD5PaazNujzz7d7ybFKTS
PawbZrSaRr4BdUP9VHKsUrMsJ/PZs1QHLylfuU8ivjJt9LPAuLzo31Y9MuuX9baU
Uf8cXfbuQwaphAgSf4JMytfLOzSezr7woqxsS3ATPupIYiYQwX0OaO4BV/lbKJxu
iK6eRbBGNozyKMKUI2yceXA6Xk82z/H8B25QO7M1stpg4OHnLcr2iXNGBARks8pK
rG4LnWTZX44UgmEVS5P3IUBHr07pAzeY1jrp6DK78Sa2yx/N3z3fADB80z4If04l
GJX5HYnMYhkjNvmazWy45/K/Ubp160uhBvoXNh7uvijfhKq5SyDxKkdPCmf1dviP
9dfkdiePtEzkEDCG9t2cGQwLB9ajSB2aWnavtMxO/oTxyIpkZe05QkDCjtDSSBCb
4FfBUClu7OiC7k8ZX6fZVLDffi9iLGCcCqZT+wZMROgDL71aXd/39byl2zfrHnsP
7G7ydjdIsvHfn0dWhyVCcx3TN9z7bXI4j2o3RdTFfV/8+6+KJM6SU3SO5GNbgGGU
r/zK/xMAJ4Dh6sNJzAMSj6bX7xE/iyNmuvczbzRzjaGq90+XA7YUQaHRJNOgGNBx
qRm3iCUPK5LEXqByyC14vbzmD647oZ9ErvQ2UJcCHOnpMKS3o1os4OZUXrjcbZWJ
MDKYjAxDwM3JM7uv/l+15IWYDYecSe4djnoiu5c3ZHcjfwCz3KyWjyTEgpLWg4AT
vKe0VJKXsxBAy7jWEf0woLvKbhRAaxjwf2xa3XQafF4ccpYnqsfG1ClCF3q3NF6G
2UXxaYBz9BzXCkifwBVi9Lx+rKO7oKb0QPVtSll1/k4MNERlOUHxAeYmYWcEBWjA
pkfN7j5xAzXL3ZLQIwarKV/OtLy+YnerxVGZBJxJv4sfXEhnRV1giP/vVIGxLJXe
tXJ4htx/KCXtmxcAXgWRsA9/RSkeJHwdc8yVPO2iCc+wq+9jGIh/j4eNRzIz8V2s
vgcRQOhm2OkOqJX6lCsE/kvWVRzjraaMY9KAoRIq+JqFRJuOI3UO55QT/uyjpYi9
9Gr66bCQ/mQExjHwcUPaQL5hnKHE+7VMs78ZaemfOqkQZ119SNBB12Mi81wPG07w
wcpwaCXv8Kzp4Qauqr+qLQRYd1SftTeVtss8m/Nds9dOTQwgNwSGJpt8oKS/FxOH
J90fc7YM/02tLoJJJGX7PettUywu0YkWMAdRlMbedbPaHW92B+CQV6l9feW/AsSz
lQuo+vVw+rlaji8mYcSjaYK33oeW7rlIDj90rTlP+9Ma0c3Z4LKfJ06XXwLOhBpB
50hxg25DLoPtQGpxiMnmmqs8DejbgG1zFJc5havVIol31RkI6UZ+lw2AVStDnnVC
F6czJWYOq3c9KxojBxXG0WL1D1eqZxpRGij6DIej7R6kDFpsmHbegjYcRsmqzFkw
Yb2qRQSMS94gH3tpfI/wvvC4pm0RmShP8XwZlj13ZYjHuLptI7cfsAB7oQV5v01A
2B7GkjBqHCo28gzElJSalQM8PWps78NnXeBZGkw0zPe4Rs6G6UadxtJzOa8cZ1VX
c7jvkEFmQVe9ELIjMWFIrrR7AQHWavc0monG+hyNECyeMKVJTRBjLA2mgCoSviBM
vY2o8UVRvP0CvaOXpSYYVnXjR3hQTZgLyOL3zORKlZvvxpkYxAQ4Z/GJcn7OGVfB
XgdYt7hNfW4n82I5hbJNkp+tf1Panan83/+z7EQ/SWpoIfGrgnKZmUbaTeg7s1Ye
90mQAk/o9CsGNtpuQnG2ykat3t+TfOKGX2yAvK2ZQJZVCuWtHu//6999fjhP3Uf7
OG1OXel+dnXoBOLnACjH55Ur55ZqEAjHp5ugk1wVPLzbZQTtDqYiP43pvHysfswZ
5jSJpYK2YkYkQgw8HB8KSG5GnzY5xrRP4VDpWm47SDad6SA5YSjFOZakkokLnVcp
d2Gd+y7t0vzC72V4hRTpqsxcSB2Mz1mJuHhewtsCAxOV+TjYX7SqpIwDCOQnJby+
N6jIjqG3CAfXXwuDAmsw0ZzLHhnl2Cth4rgJG/7+f/qXAqXWsvWmV+gFWEtOuLzq
/VKQQmeuVB5Xx7Zy2ir9AwX7byeQZEOKA7oE4opt4zGcDkL0XLUnN5R1b6up4Dy9
qbjSV/sRk4H674FcOwNCfL7rgc3XO04IcXVogjfZwOKttwx2pth77iT9JsGs3Bc4
pL6m2dK201X1p/X+PMtGSQDTX2GnFBAA9KZHZpyieca/ZaMVPFJ+ey1lDw4mKc+e
NmFHC/I1ofR+PBwsNZmSYuSDjy2Y44i5IUSsIhe5j++sAOHAhmlq6y2APfSgcVkd
ZdiKPxnhCWvx+cRuWnLZtUuRKZ3jFa9SoYlLNQRVeQmoJYS38lE9Rp4p5qzYTCBU
b9yu2Nmh55jp0vliYifbJDvZ+yg45w3FxMbDzVn9ka4+sWvKfrzDW7QP1perGCaJ
xyVRXefbhRDkR29MlTkzvjGGdQeZYarSjoJYR6WOdAFB0fuHExD1aydbygHkoEp9
69XWkgoOjXEpXBYfz3XHbAWPazZQd9puOMNQHnJQqGuDaGP/cT9VULoiq9LRxRqS
GvBRdh8XoGctdtIB9hsLvmfy8FAQFJXGKp7qRR0BoBvdNJIc5QtHflDAyVbKeF/X
5HsjL3XjGDoxDKOWN9k+EA5iwYoccl0SZfYg/0b/As0tXqpwqZxWz0GlPz5IYe5r
859saMFJRmRAPLsc3a40n3bogVF5Bjb1zKGJm4xvC1jDwTdSbsnnqz8bk73gpdb7
hUBlZY9gaFBLPVRdQz/EK0NKxPnZrL+LG5MNPMppH0sux3pHWPl/7kidBxXfBb5X
s6YLuh2BEg25B2DKzCfNZJ707CKzlWHuxpskJRfAAD/HxUoVd/rilmf/qa8xqa+R
11KQLtCzokI4wn4vwxopE1FFtaxXGzYVTuImH7FIFb8G7vH49qkHTXptWldAmCR2
/mKmnnMN+9VuVOvSue2R6vlFXJpe2XimDsGx35l51mR6zNuE/X01UoMRHlI+cb7I
ffuNttlljAXysIZOU2M4ZtGWt+s1XCrckDgkvL2+sdmT3YeUQI3mJa9QWuwXruxi
124fXpukwt5b+xQSXFmS79iIXQf2OkguYMYb4Nd/3BvHr5+Z+CuHZf+7TZaeaCRW
fG1ulClyP60Cg4qF9/esdVJGjIyKPgIdB6jKE9PRWXIru8yajKYjIEMfWodOc53h
HIwCXk7xcbmyoPQx08kVhYWZehiXa6x+yekJgaIueBgKtsJePuwuo4Ds12aNwhmr
bPDC7iQU8z1JQdNgQzqxohJztGxeqASkuowsBd/IN1EeIrdg26LNAVyeTLxoLqrV
4/CJhXmWTwiJG+2dTRlL49tVyhGkgwyDBOl87HMrC2Hs2x/TPkUu8Zlp2lPx5F+B
/V96eI1TgBRwOQdycHL/zKqCHIKi71XQyWcRHW7avzc2z9ZzGns4/CnZ6uIQL5XE
CayBd1aO8nU1gTGLV5XbCpQBZzQEbIKffZDiPN6aktQ4KxwlMZv75ZQsWd/nFgIR
6TsrwKrF7qbxJaXwA0UWuX5aupV5xiKYyqld5o58TRa/2gj631VhJVuS1fQJ6FRt
muuYIxQCfQHX3OHn4WmbjV/Ks8h4lQb45qaR7UkxY1tT+LX4leVVqozba4rmS7ag
rKYv86SQgHJJQ4INT5s6NYHAjzK+GtgttX1xxdRMfT8PU73t1K5arRNfIweSp/nY
JsHfeigB1rZO+gFSO3WgxJhVx04l0rSStIjSjiTKXDqECzLzpJ9LGO/gxwJQbkYr
w8hOzrZhbfK6k/OhmhTH+4Sz8q/IEKKAx7s71VO47D4VaY5KUMr1fuZU0v0aDYE3
7Cp38duyIT9g9Q9wGqvKoq6kfhlmHH+UyVGixml19MZjN5RooR2VmFuIGNmpJ7jZ
HTMUE7rWJY5t6bQ9N4HpTMOr4QhQxgkpLp24HRBjSAIntH/bmUPpRjoDjkJRIr3x
GEn7AwxCJX86x+YP6jzF4GCId0CkhAvNK2GQ7xz+vhrtHzliMzb/FV/ULn13DX92
2AjtMFVeGOcWyphOG5uc0iPqlPq/wDbDRBvjLbxtCdjk/bdJTVg7/UKA3oKzs7No
QrpgGFpiJ2IZeX9mUOHe9NT/UhVgT5y8H8wZeOpxlUlCp0eOgmNpV5OgfpHlxnPQ
Gq12Gbb9XDt0es6frhP7mrHhH+8kLqSAuUf3XvnvryVrhT5QtDj0foeYEOo31S85
ZQucddEzurOQFjQGvz5PV0cA2UmrP/3+10sknAgf5RY4FrHpvtwPpTGZ/8Q+kJMV
0573dv6XFwmLxUoJxGZb4jGvLHHFwH4Lk+6KMIxDNSsP03XHeQcHvtLVERoBgLn3
uECMn+C5vNrPyv/n6trpjbH/kJzZPyATeMJ6jfaU8rsHSjh4TrUYn/U4mm3CdniK
2c3ZFaK4hmkQMrGmWzn5NC7jOxzF/3oF9+ENP89sdULe5e2MnnqBoearokZIJk5p
/ypy1e6H4zTed4EPx0+EeKnpZF4bTKDImnKElKhpxaZh37Gwy5Hg85F1Kzse13j1
cVcIUctYQ4d71hH+28secXNhs/cvnizxmfzQtLi2LpU8xwBE32UbjuTusX6JvE8A
b3CpQmoxR6B0xnbR7dPoKDOcydL5uOH3i/hq+Soit7OA4gyaQIVVufqaDoX35tp8
O1iUexfcXF1K0YMRFL5odlxzABadjaQWmbo1QYYHb4AFRnN/9oJ9fyFjI29gVyWY
hZWzjYqAyzhOKzciAdhTbcpItPitwMGDJ/+Vc38qY1wn+vTRGdzn7Rx9z4lG+nd4
GxJv/Y88n+ssBy1G5xssuQYkDSJd9KEEUOyfKKI+3bRFQKIj/0AMIkaB5w3ciCM0
NeBhBpI5txa+h/ftGVc8nihDlw0POWWaNnsne9KF8hhcI8Fx8QENAGOn0fuoHAj4
Fuo/nUskW5EUCjeU7kfpTr+70ifLnbHrljmm7y+MGXbswwx97RM22kI/NWZOMXP8
78wfdGeP/xsd/Y+29p34JUw3EnaIVl67G3ply5PrUQ+H3ZmdGZtDFMpgFt10AeM2
IFQtI40jsiXlxLTTqlvhy3dBWGy3e9wWwe4i4oZoI77FWs6AcGfvvlCJ4tHeHrOH
dy55RSgJ2rA1kBW4EU1tgq0AUC5HACZBFut3vzmTRSvjtxPK5SMBqzO1GGDvqI6k
K6In/dVXaRClpSYajUx9Cw1LW8zuRKOFwDOFzD3zmaIgvdY4luxz3Kyg/rcdllt7
nE4MW/k949Z1GawV6QEBDT8+fD50TCyHwFL/W4bESTYIQAprNteb8kLxsAh4wHp/
X0t/55zSFEOzC6JnC9XrJ2yApeAHG9e4NbO2qIOaMNt8FI+6qWJ+3ui1/AejBZw2
cEO2x77PNtIRn9Fhj/UF6qRYhGNrI6g23o0+kjECmvu7oOy2TA7x+JMSUUVAYsJT
NOnt8NzBMQ9a7V3xL7QqymihUlGhvAxmZcAfYAxZDOOXC4so7uKmYXIuDIL6yj5a
Q33+Ei/pWbDAW0CyxrrxgqWk365IE0BgC0jAWxV9RK5kWVbpUz6iftza+FhnGjDy
LT1hrk+ShDYna+8QOElcjgGxe/IUUVcz2i/2dLYiGYV3+tMpCHl7QGPkIcJzi8MW
DIDksukO87+w7EaKv0sL2NbSHk+pBxEluQVLsDBOOOnAOjwS8HXQQNoHxVsg27Dt
IFepu4J2aNS0x0YyE8MUzBZCCxSvBJn94ZEJhqf75ZYkSXWCnVTuSdZZjwkBi9Vq
zJx5S+ve4r8sFJm8tK1u3Uq7mOGvA2xVdfpSOLJr/SG6ItOP+7h6vRJxwqZv6Nk+
+aMRG3T7f2F1lXPiJBLr7YIotyRltH5W3IpNu+LGlI+HByyeBjqPsIEdTAETlbON
cfiZHRfHbGLGRglWecDQqja8utaE4sQ/y3/qzi6ieS9liMQKD8sqUFs5quqhxhjS
mfemstTlXw7TdX/UlTUnCXG2WGnUYRRDTb4saTllor+4tnj5fDwfI6KaHhqwvh/m
bLHYniN5pNnMTRDsq3ai+ITU6FcIMSl9772Dr729t3o6aW+9l3eosHCMKCRdyWN+
DSF9B4zGwyP1pFQuEo/+QwxBXpENZ1TrEU/KzGYSqcd23B0O2qZW3X14+/03sQea
9Lnimi9a6FSyPYzt8nKtjEAhbenFY+uy2+Ca7wK1aw359aJMk92YgCujiXVsWlxm
qbV89u3YKRl/mj1qEAjsqieyCbXH3ti+7NCtZRFu1/RLyIGasHrMj6Il3RU+dIJW
uEJ3n92IEU0cYL3gMQ/CzRBer75UR2XXp9/uADJHu9gQ+mmYUJqPq5H09/0ng6kY
ODypt/YIG7J5gO1yyqsHuURnNZiItJK+qul1B3W6tYyZZJPWcaXzHb8krOxiPLS3
Au1t7cw77ds2oLzjTID724UL2l/7U4mMLQbWh7uHNBPNO8At3zLFDTAEVMM+QO55
JA2pEkHcZ1eGa6k25JhTSf4Y+9J19z2TCq9SG4/WUNWXVUE/uF+8E4CX3hdy/WRn
VK2Kd/gdwyaChnBnq90jpn6J1aE1EvCgcspUV5eW8e+BtC6bWtYGCevImEsZh8XC
Tjp3vrWcZpAi8M9FehVU4cEbz5r3zdG96O/xSFfsj9d/d2J4ZG5UO50FSKIL67wF
as+x2mY55AAN26g3WWJ4vIdDFmeeQOfB+27WiSEy5Fus0VjdR4gbvIJK3u8rImVl
5hJ3cwdQiDDP30IRNkOtvOT52YtSFKpIe+n568TcUjDT+22v4cq/Fd5EA1Ybxa6S
rslFPai/c8ozni8FN4NYf00MYT7tNUYBHj3/83ToiXrBVQiAzd55MaMOaBMp6t7O
rXSLp89k0yUCpV7wDCRsOrUdmPoIJT7wxPTtAk9cmeqmADrB3veMKJbSXkzAtNBa
RtkVnlRt9rU0opgf+1PHJudM64t6SidZtTZa12GND36Rtj94+u0F+Za3EfL6J3NZ
ziMtleB393Fjrs6Ggys1O/SdxXVf9gRiDjjpvALVe1idgPeNPEOumysJCMAQ4Op4
Pq9+826yFD/Xzm3jwievCdpKziqGx6NZ8jpUBJbwVeops7nu1ntmMfXVjtwhQ3sy
iMQqBOMTk2LoLbWbXeQpK6PCH47wenKVgvCCUUlMvEcGlqpasaWtaowdbvughsOy
fu8v1q2/nd7ym8MZuDOZ0ZOk2Q9se2FuoBREtXEEVn3E64885Rzzw7rymZyT5mHW
QDpvGHzT+QCG5bU2AfMG/k6SByRTYWiCRqD0mbN2vS6/9TCxrHJA/cTQejnqRb4G
CbhC/cOWoQgDnvyrDBadek5SzNrtoTmB2GtrMzDvBxaqcvzxJivGdASGiIBGKI/Y
SfveRu9A5qukEX3gnm7UA5ATvtH0o2L13hBHfRLhExblNEi8pA22dB0zf0L4PcwW
g25NoyHEzqX27fAt0fhbnIM8ZZgAbBqzKLJ2llCCbhKEw0jJU2UanAGEfJ5Ol/4k
VsjBxKxB8ieVX1hFNCvvQLjd6mR2jT4nbmTgi1feyix0OuANz8RpOAN0yHJ65ewz
Ua2LmRTrR98h0JA2KUvH1eJcu3fDLJV4TZtvH0HGGPAbnC7JURoZqMI2fdgNvJv0
APOB+s84f8pyoZIwvzIiNVxy4z4G9OwWCE3taY+o2vvYiN2GdhXPmvDrkDQzCgy1
itC2hJGV7j9kTAEq+qnr0jw4pQdYNiUG6Qz683QCm55cqdXxgeY7PnJus15DO9wr
wzBtnndrbuEyQ3DkKnyo8QDHuVmxtKEL0MgPbz/0BFkALp+q7hSrk5M0D0tDx+oA
CCDZdwv0zbkvJ5efS9McDAAtK4AyzQ5teYI9S4rSUG24+Zds69e4OJ/b3OhS7Z19
QfTOB0vaJXhphrWMsjj37maSRS7CXB8AuP7aulo8MeusFwBQ9zPqLjfhXrYAWEYu
PLlPp33u5f758JrEWYRvXA7+4jQlC+p7+JSXK4FeP3gaswBnF8mLOnWdM6Z9xI2Y
ISHMBC2k4rxNeTFEc6hhJtMaXguUFpMPrx5sfq79h6KaQY29GKIIWNNDpv24KdOA
casjfrKfMpcYQkCgXbkG0F+Z3v040sz+4qrjS/DeX/KaoiW1rcO7G0455Txbn32U
aIWr9MgjZdP4cSOM3CVjKVfO4yxuXwc2PmljBzLEUhR/kuRAGV+VojWLlmAsInCq
ilLFtRh5cCk+e54kxvX6Kezr/GljldNtS4IQpGt6dVOyXPUyYbaFrVwiHU3dZZaH
oO4kcrolHMoBMtTZsi0xbuFJX/hzp4wwrLHeL7l+1qOm06ayzNe8ww/nAlRGCABu
Eow15Z16YV3Y6cwsTplMqKfnp/krWeAV3T1ORg/vaN9Bycc1NmjARKd2HfbXuvyi
IsIhFvY3f/AaqF5LcLa4EZjEaPwgF7eQBA+0K9znM6ArtcA8Tl7LioaHX523p031
GrOaF4p8ZfQivDn4q7Pv14E9Ydk8NMiEGd1oN5IoxZl+5rd2UkF86TXNAW8BIM/q
kfIzx1yr6TBYacT5iPNx9cMrD4EuDxOLKL26Bl/mrVDDYr40nitQRGX+qzfRHYNK
CG0FsVB8ck1qj0vpSnflk44hq1zc0El3LFoZ4WbeBo0rULtd7L5ogTBDWEJPQsFe
mO8XumG0ZteKMRn+AelJV7kJGOdyh0tl5gEQ0i1gciw19gCPupnpCP/dshMBljD1
kDUG5W/XHIx3PBorZ8xQdwFIWJgInj6F0WhDIwI95na+bswTH0dvvIRUmjMedjY/
Q6MZekAp1tSX0i3Nj9s5RJanKAwJeRwj+qfn8qLVlAE2FZA7GJu46iX0Huot93Ov
3WLm+j87sIBvd87Z1/Q8JZaEw5rCFkjtDUmcbPBFqvRcZOGrxFSAoZAY2qrmjgNZ
MiaNKt8WZnuG31nPakPWsGzeqgtfyebhv1Zrt/1z3cvqZuG2u+Q7sC1jeRbM6bF3
VqHXZ6w1YuvV7Yuhfmrttna+aUSKdHlgnYXt2meRDoFS8mjjq4Pmgy0zd8Ra1l+D
HC9LxyGIvbI35lHTdTlWIxKk/MsGVcynv6D8GWdt3gBbz7q11iryoD3PDh/rD4Xl
X2PNMHkUX5H4kmOy5F9pfn16IY1SLYdT6cRY/AmLKsImCbeVuuvtG7+SC/4bkJiB
bBu0bsCXieXmTIxl6p5rEbC91xoDNEB/OL4OrawnTd9myvnm/eeRPwsFGeBhDV8I
pdob+8R7Zv/RXSrrktJt7CNc3rEk8Q/qsgrQUvzOuHacm2TMV5RtJajg65kMTUm6
b7P3vUsyuozgpJmAwYVXMhdJvfrb3DCsu5T3dlfgBvTyOhNzw3PL5m+Njd0kh4BK
Rd9BZMfpL0C9+b467IzZUrkXFTgMFkZmHcS6qZ8XzUEaWD9GNyUYelUJ+ygtqE9k
l7gk5LKY/dGLYqkbKA702MrqzhwU+UJIBjtVi9t2PNtSPPkLWor/MsRgo953M0ok
TAuWzkO9iURoRcz0WZeO5eEWA2Ek2vRqJHOV3td3xFDXwDzFsqKWbla4qWXLavNU
r+3rIkyv29n6GQm5UvYXuJE5b2fqMmPoO+2NqFkTJf+f/5q/M3CQAlyQVwyG/u2V
Md+zcSlTAvrRgHqmnReFIeHOuKMDBgdfUJQ/cm6dFMV4y0bPyHGyL3YY16lu00PI
wSFp0+2oC/EhkT3FWAYUZW8HCRbhOznNoOK4/AlbsEjWVVtrtaAGSjmpfiHkTVnY
BEvrgE4ETReJxjFTY9ibhMgz8fbyS8bZZ9kYCQcHRtT9677MdGAtpW96R7iPJRGj
RKstKt9a02vuGeNpVRTDh7jhqlHgmSygJImZ532oubN8kBQ9quBhkrftr3g+BAvv
0NEH4qyILa4l7MZ+gdoEl8/AKSn8juqQXZIqYlgRurprT72NiuLE5zpSMsHtPIcc
FUI4n02B308LfKl+fwp++L4KWcmbwsHxKswIucCnar90f+SJpEXIyWodg7ZZNBl8
uOiPNRTuxE+GLZbIc0S2GsKTwVmA58ijgdqM0fnrXaTBnBqnSm5VZ9T/pP5IJo+q
0tN+MywNqmZ7IYJM99gaOZUpxpvVJaBRF8fi+qLFoztyW6waK6rtTu+Tdzw9G316
jq2We+BnWaqpmJut9TBSIffJUJu954MKVS0lSSNk24aj2eyZJMd7wfoea385nWgJ
4upAsjaTvhJ9NDLy5nSVqsxPljo0CUrmpo7+8ly+eW0xBtE+FxWEUCh984hyPduU
DjJJAtaRQD9l+0oFRp/q2JExN2d9IJp9OKOUlk5hHIybenQtRQX9VzfrE0HEU3Cn
lcu8qSxZbaHho5oorxWIotRli4zD3NXquWhM0Rqjyu6uxBE5s0TKzjszrAVQmEg6
5xx7YA9mC9gTMtZLAXYSb1unbl+BticXoLKPRTeUoW5x1Mrx5SkgLKbz6QII8Oa+
P6MxSysqYsBypHT0JO1IcVj6k/E3pkXGfVNSNL+3tmXCDRsuL25oVJ0P5Z/VF7Ix
M/REzSxzyC/XMx9+YDzK5TnMj73xX0cVAc72LLIoVpmb7ORiGt7CaJDBXIcv7uM6
xOxaZEafEQ+VUxoKv6F1BBIfhq/mZLjvZk9/MRrKiLxGxvUG4meq47CIj1n8cpy9
ZVd7djmFdN25qSGLZ5PBXik3XG7ipP6wwlf40O9nIKRqFyeyOtWK5w2Qw9llr5am
FX33cGv0Mvvfb9984ZzADQ1dIuar2kT8YdLP7D0V9DsRKuETP3hDh/eLABllTOtW
uQGVJQxbtm4VPYZB7VANKZAUgTZdnvhAzMN6xrmcGHybWyZpy6DQzJ3iQoCyhb1c
IRR9mgtQfz5litzIfpxtFxhYaNd2JFaLYVxIzVWuvhQip4qzsXp0SwWITuSViH09
fR/+MglwRdG0vXu94ljoIM+EDVshD0ZPW7gtKD8rINGpcP86ZpQV0vtWsEa1vqOd
XaWUgyuCgQN7C995hXaHX0tT1tgEFlKLiKx0SuKZb6gFDoGdTdJigjHn8Uw50wD6
gsdqB7tmn3zfwoyDX6eGWEa4mQ6/+Xb8ZidcSRoU66ZpbBISYeRxjbLxz64H13hq
HLtV25yUk8i4vskkzlbygcrveTVJwYu+CSvnPSpCNUWXNtNERNp2oRp/lTcW3oRi
mFw6101yRo3jmGcksjFO53tuN2ku8/WMU1TmF9eQhwkODhYnL4jWCgBLapFaWq+a
/hEzcdLnSdXASu3Lb5Eb2gpxKBHQuuPQnMCDfftIMVIecWrscsdsfChRyQBEN9RV
bf/+kO2bNZmzCc0lo4xEy862q7AObVZcFO5WKJf4NLp/T1TRNN7BFQ0tmcc6ZKR5
McS19Oq0kziWuRCkY2SrXsE2JJHqNYeFEVvRttLLb6hSktlozmQ4dKnu8ekLcD5V
f55fv2vNuYv4ADNLQCYsLdSElBD939SF7LOlZI8rWPSVkSNSH27dtZN9l+NS4bLO
Ld4AOWuruGHV7aa3DfKMBeyelrrHFoKQ1MtI7UT+iTrBDoLt3EcIxpWW1aulPyaH
WoZDl12I+xrqNsvwSAec1MqJ3eF7IjTSkrzQYbzLl90BeQs4Jp7C3CJN8CgAy7Zi
wKAojuXdqM2A4QcncChQX6YcpvqOaoxVMBmQvMsrIJnDT96kqrD8XuNZvVolB8jq
tezbJCGFp1BaDigTV9GYmLQJ78aPhIHKgFHlI79ZyEAt8fJg9ZzoBC61hllw2QZk
OHOI6ynUWsB0vN+f5bWzqFTuMQ9FSshqrx+DtYqO1SxkyUMjj0ymOtmVA6K5D1jp
ALtJqICwWK86EWompffgCxA5RhYqrkFoRZCA/IxIrI9gMHe9c1rfRiGw5KtplGUy
VrXXtlyBt/u4snR4mRe1WfvX8heT+eX6hQ2opImlQk9Xg1RFcmDlLr6EgxftCKFz
/4OnnMOyHB9HeMS45cDTR3EbyfD7AaQuZpHg+zRI7FjKIeKGyPN/hIeTwroi90ye
FLC07IJUW+5KMDCJ/TDGfXmIvHOE4M/B6kMGn5HJMEeUDE9pmQuM6Zwyt+9zNF51
n3jz0zz+1PeLXPU9oelXTK4hfuHVwoYfwAy2+BXM4IRWXvq2c1znhYdEi/e4uq/O
ZSSCsvCE4zXMQ8ClVtsZPkPgHRI0poCFYxKUDqqHkgp1Fq16r+SpvPi3R6IpXE5w
8Kw0yFfpTJsBpsQLZzETo7CN+ezQeq2TOmcIrJQv5ah1FN9lDMzOtsTXcH+lcI+U
ki7Zo34jVtNgxeTcT16hi0hOM/Gozvz3VBf7S0eRRgUnQnvebgTPmvdU5nVL5Fms
fdeVEDdVjEbIwi5+hmBJgZIMnAGHYixTi51oddrKHge0ycyCZryrXr9xbW1K2lm4
l98gWIi5S1IPP9Y8tBhWA3AfMyi5QQanm5peWuWMulhqgAKkvoVhar/PMkyk8X0Y
3Ny/NG+JKbBE8RJncXfcqg0NMaMKbckVazkCuiL+hr8fDTttS2nV83qVRfEMu9Is
zSY+6Mci9AA6mAqiMPoy0fyYqohI+iWxnT17UFlMsi9gc/gMc5bUfUO+PTxMtpd+
RdqHxUSM7tSsdxBII587Pu1/DUj8DkgHfBzB7o0/nVWE4r+nZeA+vNa6ejnzHOK/
F8aYZWI0l6/yT3NIdehBaDtU544UEKj0kIjajt5hJhT8pfMCVPp8bHUwtO3P4Hkd
DnOwKPglyjXpr8bLpd8guhOBZY6engCGqf9sTqS+xuyBG2KWT6T0l1ihwV6jd4XB
VWPRISwKMAodmrw2hImOymbtAZoqIqVGqG0cdYXashVQ6UA4zFTLqg80qgCgfxsw
qvrlJKavykTNMoVlsNdqSCM5lWM7Ac4tUiFcF2/W+Rft1bGLJJr8JRWr6v9YbnpK
KdqiRnFbRExPfCG94Dwqhz2XjAuK2SVlPJYl9VWOn3URWJeJ7pp6aisOkeS4PTQc
OFW+rxVks3/lMG5V0bdyPBHK5V2EtqiXYzpXXY5eQfe16FIaI30jqY0uazYZU1rO
yqoOPSU+JKPJkfQcsn5wZiuyTpP/gbMsbLcbQ1nVzxWjiO1OhmS4Phsf4WqXjM4C
ISbOK1RzBpqFyOS4awz6Lg8XpTmNQDh87Yiy5e5LWEM8oTm/zPCkc1359z8U1Z2f
iZLaa9Gs8di8nUNZfS1YyPoksYaXpLvEpQW0qE9shy98kIJBseabdKQt4ebg0VZE
hroXxrPL72rCsBHZ+Ekaz0IpSFGeZbmYGb0jA0ppbmCPFDf9elFWZWPb88YQHtjR
JjMfv3o0u+k3v685a6CAz/FGXJFjg6khRafititwuM0y/1+oTJKigQTjU0dhlqz5
elyyowCy8Najbu5aOhgEkSw0VjvDaNwZGxgu0kxtdQXMiNJaNnCry0Y/Wfum/G+n
WxTdo80YZk+UpnOn9E/vXgjBHD8LzUBY+zRZGiYKs30C/nV9Nz9wslN7KDL8uRjV
UFGIoax83viPwZ4iRszWHcIW09dPEAQPyGd0YcRiRI+YW+lCh0TIS8eRL0hYZmxV
N0xWtDP2zfWK9Q16BULDUHh1Bf0BYizGISxszihgtsqhFmnNm2dgVt/pIarVKoOh
z0Th8wPUPJetNYKAwkbt9Nm7lndAg0/rCgVgFymMzuR0m1mWm1mekNRvu48A4boA
8midwF729fFzVjdtxA3OT6+aO3zD7FxynIVDq9HL2jLBV6C5vgtvuNK6FrFpebxN
EmN4cbdRUoIObLQ6V8rTEEA+faUNHvTwV4d/LF5o5Qugx6rAojjxfUiLG7ONZWA+
kIYGiPu86GF/0t4YfxdnY0kdidqEFpJjcPg7QuhavXMuE9BpLgPaay0TkdZs9Azp
PJRqtcGJslkPAHIQy3U78vTGXE4LwCT3T2L/PfEuhznGrGE5PwAyJnMxe/ZnHjTp
UNZ5rbGgwMTfYM9LfJm4G2c0odGVxJcN8iolJuojagB0jgdmzLHXnCgWIPShrt75
znrcTZMsl+y5RXE2I8KPmcD9G8zItAtcmzbWMOqOVEZ+Mx7vJpoLzgVEuQJlq6y9
KjF5RRBA4qHS0EpxVpd7u0o2iq8iYpQvYmDCmcM2lsAiR69SQjxvW4VTZJUv7NgA
jVdt2KCM7ksk9bS/HYnj3c+LrWdvnqn8QUhoEqUF+MXZLnmvzG3Y3AHjGIUowJlV
EYZj3GC64FHmkr21d7sGWmRht8e3PndeFqjuyKogBwKVJYc4gv63mB/wugGlMRnq
C5b+OAKEZ5bYjxIq9wUsKOQowqgwgojuJ2p8XjBWkniGEPWfDvoDPmH/rNHFhPv1
fQiwyyeXDIouBRkCrriLA81KUbWLsa62CgCRxzcjWyddAkvmLKyt4DB6JfCB/n0r
2SbfTrqbD2Fb2r9jKXPPvlxrgFzBZMH74SwytupkonsPjryXnhHOJHBXQ/YYQRg9
avirhxVWxtvJuVefpfTDK2f/eJGzECHgwfTvPBt+RNsZlxaDeWNMyJHxFvdO6ns4
749QQ9BsuCg0eWrZcn1SeFtEwhQZFWS32VSmgEiK8RYEjLFgw+qzyJTXU8Q56HnH
MCciwKRT2D+iPAFlji/wEzT8bT7m4LL3o3Kb8KhPuRagt/HZY7XhmJ0i4Zk63We3
wLQtSZolJpyJ9JC/GBLkkAFBqJQiTqhOAK6YYgWyrh7StdooJJuiRsWs0hvUh2bv
GLjh4RYffq2hy6SabnR8gCVdi6tfFyuHoPrKg5a52FUW7Wz2NO/NcbwLVLiiqHgV
qpgUdB7B/Hkzaf6ZPm43OeITj+6sguvpcV643rZtv/ZmARPK7sOlRL4iJTVoHkc2
qp34u97TBqya2Qi9vnFTVPF3+eV3Xc95i7k5AMRQ81A8EAM0awbguaZRRqFQzhtP
woNjh4MtyHRU52tnvxxEPgd4bd6FyODrU4ZIGu3DK81hE3oLTVgYEJSW7oDw/3ZD
OhyBZV4PcHolHYzuPRitFmTNRmdf86fxhXrw02T4x19Hycs4NBpQplzxKpAjvLDS
GERT31SKb67O/+8wZ16MrKMAA8gwOqOGw3O9gE5FpbUZUtbqIeCBMP1DNzmibrf2
HSPLgmrTHhXZ9xc2oHW7jBx4fBCvb4mNiZRoZpcUhB7UzDzp7LDsVzbJbILWGFoc
/TqudGTrmUarOwasLsqp/szqvHaxHHLYqxN4U+QeLoDqLRfOatGi8giTk5Q5m3c3
mAYu5IRNXN7ElLIP8GwHCBm4Ksh/wzIaTg+OX90ohBSmzDTMhjnbMD7v+pBOw4GY
h3qOwk/yhfqU+XK26BqUFjhr57nqPvdh5/Pk1zwzKWGFK9xjkgUAqM6UZlsVhBpN
JRjtEo3RyPrHsoW1af/AO/rti7ekXVBZim6cPkoxeJPB4VFupJBOUw0cXbc6Tmg2
XLD8nJUFRHBWEAbx0aTLyubgUuX5Lxg/ip1B6Kvs6/EMGqVAVfw77OrHo/3aH/vD
c2IUXXVcsaUl5JiiZYGvOEdNX1ckvQ5n4ctOsLj3YVllWCMIo1QZpl/cU02u2kNT
ntpbg/YdkUlTn8ei+gW2qv3Fg1O1RHujgM1LCUY/IocZV7jI0Pps772RUHwSJ5Xa
F/wXPfVKii+sEJqP8h29C8z1X7Bju5QhGTx9Juh+7ZswfDd/QZo/suEQ9GPDHMDP
u1b8PAn4zKYiCRxT34sChhvdx8lecvvaVdJGBtPwutTIBjA6dtbHInshJ9aOcWB0
s54vUBZeUqhHJl+5K1I3Wrvdbi9XvCk6ctmpC2pvt50e7JBO+4PCpmezZbvNM+n7
WoL9Y+b/VC8Shcj4LEot2D2KHIUXIYchzoP4fT5JUXztuCYTGLz6xUlNRBuXEVgz
ZHSrEzKn8WvYDoIy8tgu8tPLwQXyIhriAhhJRSq+34qsKL/xF684pNnocBCdGBXI
aXoxkKqwtezU3/1oHhYARKcw8uRmafOIUClHvTg3+2tfOjqoM5KT1bSvnMDmvH8A
QCpEv8135oAm/YxDLuTu7fy8OfM3akjJlHu4Km/THAjgmC2zULmJ/IisFkYOhxGg
wSZoNN9nBdXwZ9FTa0PRvBYp9PuRMceXoRAoZL4zfGiwRuimd/Fb0uD1ldvXaXrW
6BTbPIhSmFS1ZGoggXrpcW+t0XLO6zqIj973X3nhUBC37Ejfzhao/WsLvW1xeFuG
rNKuzQJZOaR1sRjelKnDHY9OstZ3dPqdDGZhU9kYkr4zRtGtoetl9z5UW6/luCZW
VrHYbxmUdO3QPA2CVd+pCe2gzv07IRYdq7pM4zhTKCgIda3SC6CH305Io0NPBjsW
2H5rUdwMMoj5VKnjn3t3FtYL6Wey5MrN4VWYSfjSfSTk2VyLjyKrESBVTxSmUTqD
pKGPptsIVpkjqbJY1LC1srHn5B8wCVhGw5R4m4y+6YbIdEKIR2n85hTWNIBibtCz
M+eOstMODM1PdoJoenUD6Dm6rdgC0V1810ya8TyqhFOWleTjxEbea0Qe4J56Fyz9
lv7iclCOGyUbkktGIFU7CSPpAp8q91iYjranf307DmmWna5YxM6sp9cjKkPof8x6
8qYX2siSj+SpdEeqY5u+KN7ClVy0XNDKnGqGxnrF3XeOSMwJaxF5JuehSAJ01D82
P9ntVMrnCpM5MlvV3/07iWtAJamVic8UNUd9N412BhLlAQvG/l+immcQVEzb3N+/
HpgXW81YAe1ozJslcRK1oSw5STOvGwGAFqwNacNnaNI+yufjZE4c2UqHm8XksuvV
PEXzoZrZg+KaJAH475BcAll/Qr15LTrUOwKHhaS16dOxIJ3yK+s2xJ/OR/yx62IB
OuoRqG0+2o4uHv5I4r8UNH6XMGbky2sOqeKq6Op2H4wdCXn1mCLyV61OnaN2ePXk
GV+Nt51wrwCdE60X1sXvBjFeFUzkrbXzAjicTdTLOb2/kKxCKTe+3/7b7slSRRZb
VLdf5S/NXzrICKOzwtCWoG2QHmG9h/rLUnMwG5oVZLD30Qtb7nbY5AO3i7JXnhnI
RHMnkpwAXSvM07n9tBspeHMKzEkrB0wThMYd2duzB7TmoT6EnF0vvGpeNyQeo1Yu
eNpiTUs5yDf29n4NdgIFOVcTBFGvpv+RIF38YPEoTPRLBA7yeN5vD7sCzagUE0En
6WyE4Fr/9RaThhGU1PFHJw4DKKr5/Ih1Bu4pB45a96OfojCoVXzZU4kZahcP56oA
GoMJ8KMCEE+INMU3vMu5EHrTNz/UqD1fTKCyaFVf0kaP0Rv1nC5N61zb6Vs8KNKF
RG437TuNulAyJxoKyyUd0tbqgvuva8GHEfNTpZy/NmNHF0cWT9WPWsY+OrNDO+Wt
/Eovj1gLJx8LR64OE1HFRiwhxRoHd3i/r9EFH+aHEPo3eY8AYsZnRJXVHESE/is0
k2XalLvUw0EN3gkTWVBwIl7gAZ7aBPrhFX0uCOViEXdxAIGwz6pERKdvd6WURMBX
Wl5meEih0Hd8wXUvujuj44GzEf9+oELssZefJSBoNO/djtHzBdlLDj/U9daNjT60
Bz9hUriQ1qhqeVQosF0IBE5CgeAL3kHMTEpjGAK6omiMLPaZV6aeSYC6dj3cGlqb
dFsbxDw8iC/IZW9vrypPJf2Z9Tr6JsyyNtEJknd3xAVg5RmgAwJEV+wFTiZhMOx+
1jUVH9rxi8lDBvxRJyILXOmoh+s3XF264jyhKLHDVjBv2HnP72tCow6h8hsrQAZW
Pyudene/ZNzhL3Q90zeRZ2Eaz4zSQ8jBYj1uKOguAIhXg3q6aEaUBZG8iRxyQ7qg
rY8kb6/www70nr3Lsw3ah2vZBfFmJq2cLIkHf0a4LV5IucYAL1olVAgmkSHnS76f
NUWjvBP4tE/m0PMy8SjLIWgcEkJZ0r+ah89asFbiILhBAOXIwxQDAfGpQIFv38Fe
ebOPXvyFiYOB2j2gHg7EK9keSkPhv9inR8mZXpMVy2Iq54AHSrdwu5yakaxIp81t
tDmgK+ciB+0NokzXpz4t8wJumjjmxsiXETcIu4ecOz2pPOG7WhPmC8P0FtxjOgp5
Ob4Q0+TvFaVa9XeDJ9tEDQrXt5roCSU6DDEN3aUwWMuXRgTHKlsIclTbkw5vsQpT
zVWai0Ymhipe8Ehg8bCXcDNk2hSHs7ZIIoqtUXiNzWLuAfqIwkWQQ4LZziuKuina
B2xiFTfgR/ZfyFOXCCKs7XSaKNfhJge7KSEwIdJibRLILr6aAu/v9cvu1bG3dF1X
QehwLXWuMpeE03FioEtLclEgLyxGheGE5V5Lt7PqvRqFtQjxAXtcu/pdoFhByEPj
LkEkqXgTk8E7Hb0vUtXizHNEcx4+cZ8/6Y/ezd1I6oWAAnAc13//wsQin7wJmNRa
DdcTF7F4bX9JvbMYqd+7YVALaHjoOmRc92V15C7t1aZS0XX0SAWo9V8XdDsOq9DY
OMmObBBPqI8/5nnjX1LItGaZV/icQluUW0jTCcFg2HmARHaqUV9ZtL+TInbs/4Zd
n7zbC/6GwZ1cBaipbUMzz62jb5SkjVocX/2bH2L7VmzCgWGY8xnwIzHqP2MfaWtE
8jWNLpWidOzgcAQZfuOswIZ9GEnffzNtoTfKt/TnKoXBNIU3GgtRIen8myXy8gyV
+TxAqbu3zqfRQT/7FRONB2Crk7oQ+xeIgizuYxfMy1tOdWY/TCYzQOt18fY8aMmS
UkAaWjpPL3qamIJNGyPL8lrxO5RLEidSisKS7kpe/MJEI/WAgqrAL17k2MFNgBIK
Op88sByJ3BmjAd8O7EZDUXIbmG3WV//BypolNEOoSJYlWBRoaEMVAA3NlP08kaLx
vDN49f3DpVGBIW+7Fp1pDUatcCvc2+zp/TCpklTJbKqoSNBGn7bJ6mRuXrC8N+82
8XSppsJgFjN/hg7fyuBOexJb6RRUA8O1f7MpHPy63litBBaZZXyjBYjJWv54AIwL
yVxW7MsYlzB1vMfw/uIvd0rEyoDx39RHXPBAMvDu1Nm9Y189rBsF5tX80I18or0S
27rH62I1Ep+gqMF7uHwtpRsDePwZOLpo5H/tgAOWrWKz0wb5oCblWQzohIzlBm0u
J0wVwVpCrVHQDO3nSY5craTqE5JJ1REWgSAO5fayuYNC4Sqyw5cL6I1VvqWQsGm2
T7ASFr/DTBFV+ybsqFYYQK2mQmiKsm/CKhiBJ8MpF1kxbre8wW/F4jp6yWThYfmE
mO8vUv4Tkj2qPfqQJ2r8CWf6vmWOG1Y6O4+6+dULZFRzRjBK6J/1E4FPLHMhCN1K
uuQkPYHWe+3LmkjCcUKcsecWrwWG/Bsnwkq5TeEgHPr7e4v+nKpDO3Zj5V5urAlX
Wskb9hi+v1+/NYecAd2UShC0Z+181DZfzexeTVIO8Ml7Z1o9t7Db74H+Gh148ujv
j0tnfIhiMhmfZrG1DbloPatE1EP0RAY82AgRO8otgzRrmlvWOrT1yfoSO1Nr47a9
NpU2agLutSo3IGOEoB6IjOxTdTcDhApYJg7WYMdoa6ERUDmJYzxzjjsBqJHkPXc8
bs03nM0/ik/rNdQCq83q0XQjO4wI0xzGmYr1QonxaMo5SFwQ2Wuoikex7KXXZiTr
4+5IqL1BFrMkqGCauWpkq3t3CI87PQp3nos8Dn1ckWVO8m+r1e4jaztoxkFnSCPA
/vDpmt/gV3lxwhxyKrRl3y5j/1IvJh72ajaa49F2MpZr04Z65LTnr3CZKowuZuUD
1suRLq7+NqRKNpo80BiqcmITsL3LpzmK4aHoxEOpV1Er5OR+ghCh/TEewqT35jJf
Wgz0Nk3NWSsJpIQK4A4aj0CEvn0bEdGM7NI3yRgT2Lnl7u/3UCn+IcNsSJZ43Whv
qwSOQu42Yt++AekinGLjttgjicZgGc0plu9/m+XxpTSRoEnPggcrdVhEayWIAii+
2dWS5bb4deGRvHQ6kY3jLW8WQLi44eaJuATUYyYdiCFm7+/w7bIUtIoEsdJUj1Gf
d1sqnrwEzQ7S33EzNgwro5vy4TKrZkkbCnkHamk6R31ET8oEuNyjZ0x8Fbh13Eff
KWYsOnjY0DDUaig0znq6QIchDS975ZWZPQSRMIWcIThxSa85AbWJxAybI7fpt4L/
oC0uKkR5r4koBwYsO1O8gyInpM3tjxalcYwXQ45kQJWiOwldlARrrdqGK+WeKsD0
Sh2S2WEMI8iqy9ZYLHOcC9TJ98DueLujIdAw2/Ezs5GAxe78YejaT/SFE3fRCFaQ
g5ecEz9Pt9irTubK/j8HGPiBpw0KqD1VYYga+npN5CuVZnXXIpQ9ZFP8KGpZ/TNe
X9gjou+Mp48woDMsGgA/YlFlVutVoOz/mWylUtdkKohpFOIVSCnPN8dX1b0VtWCu
fdz067wmuMcUFSCjkGPIXCgNyHga8QKRqQnWg4N8qknpDS0uKRowouSXDyTUCqPG
IdcVJlOwxsbcHSMqbm0zW2aaPOPQoqOdYiZ/2+BjdY/StDMJwjBoynAzt35T2VfW
P8svRds6u53MJ4nAQnPGUL8lbNtq3gPXUWKVrI8n3lLC61tZnOc3RhwNKUw55Jpd
CbBpeQhdOyEeEQAGUL4NVz0tP263d1npDW8htX8sws4hIarw5SPQtCD7eh7rKoUi
G6AunPLpD/0lssAIJThqGcXHqIWo5MTAkdpBbLiPyqME6pZmpGxxIoWrDlXmcd/2
uJkYlnhFXm+JLUR6uCggCZkm3lJP9WklBuJ0wf8nNtIBeKZl7I33exFMJPVxF+In
h/xwpAfe4Ysqsj+p/pxZnnPkRRlrkreP49I8lsDindLiw9ioTK4XyxOUcjLaPGB8
gberi+nVxFugAkenKaVtTIFu0c+HetYNw+bi0TBHL8DkK/Lmd5tNuKzu9vu/4z23
6xlZIr2Q9tLW6UFGAk0fR6ec5+NR8cjYmJSzEDJgSaIZ4NhumH5BuSh5Lu+VqFph
9zpD3yJXsUoGEY9OH/FhnfnAmPgdZ4We2c+YLEwe0Zf4/FXiSFYsLIqWKyq8bQOE
jXN99dcNXinTkpwYbdjXY9TBrK5izjPzapprT4FJ1PLfQHemW2r7XbQLar9x8j3B
jgQydCbxFuxTwiw6GMnWCZMBzghuu1AtDhKVLHoTTeaCyA+KCL7LjggGwj4FN13X
YhEAFuExEnr9r5MpTAowtHczS6So7q/Ybg+eQYeYRmxMDIJ60aTXoX42aHFmBcnN
+Lh52eT4E2FZ8aJrfHa4XHpYaHBAn9dDdDV/mr6dtimDPHdZaMGS5F5XLfe86CQn
tWnQu14pKL3TWug7lPguhBU3L1v0yh3iAmlESAkqGnU7Mjho7ylqvEpNtar21P6A
k8Hl1qGHRZ3eDI1oTE1dIWo2yHG98D5PfLvUNKYVO5uOevgoZ3Glzv8zNiPe1GFb
JFxidMp0AuJwLNvxfCTckRrenHDi1xryf/VyPhM/aeUH3DSiZTPj9UHHMW4rslCY
x2r3v6utrbcr+WFgij3mC7nO3cQFnoCzrKkSPp75QQcirMzdYiZimzXq+ZznDquz
CAtnoF7btEI1eGp5nC+rhulkxVDGLf8O15X7B8ADV9v5Xv33Xa5Vmy+Dug9QDAdl
5blYQjEU+RQrqQbjfn8D1jCIfI5OuYCMCEcNLfrZZKxnwOdGmznR31VHgGRPJBoS
OP1NegHNbXfY4lfERGIrHDG9EFErH7LiAcUuoXPj6YdeIY6jbEuqkglwWxBaJQ57
8VwZvIMHSYKooF2ELI6HIwKix9o7x/nQi6hQPl4ytHrBWypFDydWHknVuwXj59gs
yn2oSYXAld27ynnt1lovUvjQSFt2PdX8s7RbF+mX0dLW0N804uo+1dO+4NGW7A+9
vOq8IQbd/Be81vl/PB7GXHTz2qMxLxRSkWhMY5IUbUScurl1NiHYXFjdGp8VpJpB
1/TdXy9oDkXTYt3YkkNgMsnJkl0UADAyrk7G2luTYw+RpatdvYMVnLIoAxUqTF2h
427PhIEmHtMUI8lZl8HPDTEuj3SJeymKzFW6viAxqC+q+VqwwxqFLDI2R2yJ4cYt
Sarhrdda0EYubVJNv30BPBHyh0Pp9r4dRBl5J7QnudcMxhMLXm/sW+FQAzu7O6cX
yA3IcNf3fIOft+ZnzNzugc85Y65gmoUj0rUzLwNXGykMIF9xP/nxw0ruaIyTAaJ/
dFJ4Sr+J6woWw5BVAJ0mig34b0nIdX2n5BiY686btajcUtYx2l/R5EcLm8RbXL4t
ZnUS2bGR8BM4ISg/L8Hd0OEm/reUh7DkQOt7Pe24g2k/rgXR8JLCoWgSsA751iCo
d/Nj2V+Wq6agPfOCEOcD96XTe7wXHsMZzgrZW7lqrLPwCaGj/EcWyo+wtlXbLLXg
X/ekUB3A/b5Rw5Z2ilEm2r5WIHHOhkEDOka7Iqie7Os3Jh7Qs9dvCCxFGG9P/0O0
Sz+7D3JYE4llC8qB10qde5dhHM2a6QfKNYVgKCA5jr4SHipRLgM7EluQ30GUz6Vq
OY3HLm8L/9mXsz4+xMICZ54W2GyXzYA+RCtS/ZsONoI7+h+KFpzbj6+YSoPXml4+
xrXLhD58V0V/oIyUX/XMN+JEjpD0uJTnMunqGMcO310XizpExjYx4KdU2pTr3M67
J7THVROZqgci1wRkvQ5KhyTcSccj1zOLhOrBTu2nUS4uM/BRh9+YPS7RB9Ni11V3
eCEE1EMcIliUVLjFNa42r4s/UvpkyHYEZfcz5MDdZ7FxisU6xEGRx0kb+kOEcjJs
bNzS8xOkpbTlU+57b55PK/K5ClMpBskrowkkTIcc498UuJWIucDz920UzA6D36k6
MoI5qeD+QIhtmkjWAPFGiz05vbJU/mP45HVqy7Gu1blqn+F7oAaH/yIzvEw9LuO3
nifO4iw21OXhp/sF+9PblLhXCrUyg2fls6dEeCUkNh9NXfWS3Q3gtt3HpWSDHpYV
2+BU+r5kSensuuZVZ5DewChmby9BC67cl1UCEbBK5wu5T/yGElHKsfYOe1sQ9X27
harimBtbX/opqvvY6BjHHj8KQ/GYtRZ87ykaop/lbktQxi2z8vq08aQx3UqTMjls
a9sITvLwDZBn25CxhAX5HboXWXtNHP2oRVIbuyfN6tB4BW7na9tvp9T55UXJpfUu
jlmWRah+YtCau4erumr/469LS/zBAakqjfwPBrzEZ8w4vYGwiCvKl9xP9do5vvbD
apjMYaRvlrtqMEFrfu9o21EAl/W99uIamHFJnpCVI3hbmKEbd70gxAXVILWGWOUj
S+3Wa3Rpr+TCoIQXiBFuPiCH6oZx9fx1iKLWNxfUEQz0Iw2PmcBnCfHfUF1/37nC
A8mKn+upZvlXdUKagBmMZtTw3vY8PlinCkiv2uAjaav87gpxLDjsWB08YbezoCOy
MPt6kj/ofCKnVptSObijSNlF2c0f2OlwXk9ACKV4bt0sPuKkxNBCc6I3mmwLtAet
JmskNH+7TmUWrcFR4IMs2JSeNZ65Uiw7Stf0YxR0RsBeYdXMvjqpKfAX0ZrZMjRy
Ne4MRI/6eBvo19SfcRJixVthbWuuiXLPhRqhLhV1nKcR6sNphfo4cDoSgEY1gg42
Darv4jCmrK6pQ6Q7nnbX2YT4wLOQ8L3yXISXsqM0LtAlSOfVsGGlLHd3hq0mZlc+
RQynow1aOJNbQGyBTDs2NWATi/i+O7EVlxmrqvqkCAr4CFxkxL8Dgq+8J44cSYGI
kSW2x9bZ3nS4zC5iEivmhG5+B0IQjbiorv4aoPLlVl00brqeypEPVG5AKqa5iiaP
0dPFx+t/2xDqQ4rHqQWfLx0rTI7bYHn35Ia2jNxcupKscL9BB4iUY2c8nF9xn+kI
MmqMac+xltl2e4yRNeYxr5FtLgJRa4appSC7xQ9kEK0wQH58iBWF62RA1BNTWfLC
nbtwxYuz88Wr/s81asCjMYQ7L2i9gN45GwYo5iZ2CF7RH6SjEHafw0mUFZXu1dm/
k7s1Aa4wCOJ5uIGhlmiUxB92eNzboD8wgcvbZvSHyHe8zXIvWe+nwQfu1vtzbDu2
0/WTBKBK0gyal03Tj/tNZkMpzEsz9dQrDBmiReh8Ya4z9Pdk4OP9Wevhmv9Fhx0D
fnXsHAuiTi1fLfQATpRIlMviQpzfPv0ralHqPoXHABgh5DRWZn+Rxa285o8NSTeB
iqA96gbnOkcJzRPEvpNUYhOUFKUrWa94D3UhZrx84nZTVrjThhvimfiHd+2Ll2ig
J+IlTVQlWDJbt1Nep9pK+65ORUPFsWkD3Ttkasq6pkqBPjawLIQxYFiYAL6Pm8LN
9IVC1bPD0q1d9CKcWgxc/mHOPwUCgZab3wGU3ZMQarm6zFmydJ3fy+AtEtgaJX+e
iqxqpz5IrzVhACOFIPPM+yr6RDInDtPNPeSKsM806tJgazrwWCW3iRqi1lF+H0iA
psPMdN0N7m5COFM4AH49vGpGpTrGeGMmvsS237eUrWBHAfYMteXtfVPAXCDSZwRw
skRo20Lt7Z043WttI61TixoTdpOHHI3FsyPJ4C6WsEwkRZblAv5mj7tmGAH24wS+
3n4IjwFICB3gnH6YAaQF5HwdzDDCgmR2UHlG0C8dhhxA75R9TKRDN8g6U+oNsiBz
G/eT1Uibvb3PoxvmtCSDMkquAYLsrwoH6/zy6LnIMKwBEPUZuY/lwLjFHKOMcJ1G
eZpXodAIP/1NVB1A+K4b4vZDhA9f653iWu6l7UlCJff0tlcy6i0a7kZm15z1y41g
UnuXjQybxcazi1R+wAse/C40fKTQ9KMTa7wk8Cy/sfzOtquIdvLPAYcdJs2I3weR
HhhI8jmL2KtV+HZ39NUfITXLHTh3gCMCv8k5Ygdx6BBSv5UarelG++DY17q+Zloi
XZsmbU/VgjwiMF5rFos+90XFZyYC9PIvNEACwwKjYOugScjloA8m3BHjDFVuepSP
Que/6z3fbGs7H8Fvt0plDVjLnIdiUltqcuTUrktdf15qjCTqDFkcKfLfTSUskbVA
h2oY+mgYbCN1G1XVY9WhW+xP0KLjJ+QCmPmyapUxglMotPlmAWQRjVgJM+Aeu3UO
7Zo8p1wQ7ptHfIDYgT2fXau+m5CzVOnlitvWnrFyrYkiTnSwgCNaFEBTEfyKFC2C
oZ+zdIC19zcXK08/58FHXEGF4pi3x8oSNf4dTXJtqf8vnf2yomFusfSmQbXTNtYJ
G0MwXnCmJuZTC//QVbUqYWqolQKgt3KmxLAJ08afEuOsMDjwsgFDqpiNUClqneEF
UFkTN6oJTbk6Y10D1WQQH+m516G0owjKcp7V79VrYo7G6Rvw+haBdBqhKHs8Tavv
FXS4eVrHtF/yDqqIEGGCJCRlRnPiplvkoJyoT2Paxp1tfQMGBCB7X+BDJn7wVAN4
PABmiPEdogFWcuaJVDWG1hNURaw3RuzVqTDRm72fCWGvlydc5p3I00TWa+ANe8I8
XXbIBtUpSf06iI18ULzncT6xo1eKTCdP8iZPgo7GnB1bdRMUrFqKtsRelga+2JKX
GlM+oSL864oWJs0dveRrgvm2wPDp/zZV1T0lLRB36fRv37M51hxshZNoJEUnPjJk
sVA2ThZ0FXCm1CRvdYUI//wF7nkD6fY8mnD+WxvMsuspMazKZRB6o1GHkZJ8+QFl
ZNyI8Z6yHuvJw8YOExki7d+IX7gHXDJ8LXmQNOYBC2KxWNYrfcfTBIeTD+jDnRGv
7dx3QeVYJ5r/TizCJDMBF2/rrG+IMm39QN68Mzy73IXII6iOfwBVBBvKj4YpjgEi
9AgRfEcdWQr1mfANVOMpsspTKPunpB0LFsOlS07oPPbREjex/N7MwSowD/aGm8Ff
Nawp2fULhuFcVlez8RMzsrnhD+Nf5w5n/GW2hMsTDWA2EGM8uMO1+hz/dGw79/QD
yB+8drVPBBGxJDN+z1yWswar4plwcTof1oXPcrLuk8AZd9tn/CpdzmPczeRdx1do
OpCsi6D7rGVX/hE66+Q7bqYz9u75VcruWuyPPNVeA/XXH+bWP06IDz3XgMRhYh6U
9wx8TgkJPKZKCxjjU1T1gpQPK87s2iW3wLkw+L9KCJNJww4qXlkARXxH4p+VdaIV
h+c6kxn6MsrYJf+8lZa4bv9bluhWsZonNVKJVV3Mds8JHxm7VQa+f1n2znt+e87D
ypcojLI36oRvCS0IEaUgxE8I6HJLcIhPJyai57yTdXFqM+6+LZ099861Tb7qTGKR
dli5Ull0IGPX0hPjPLeqpsCFS09+kr36s8HKp2aNxk+TD42ybSmx8hPQZ1WPR4NL
0G21oKHjBq0J/sLJ7fiUy6n0M8LzAXQtJky+f10Ge1OrDxpJmEAoieh2CGlUzWhm
KG6WxdsDM7bmpkCdQi2QBd/MawcEh/qBbjxplbqOiYhhAWVCXEO3aIeNIqB5ZJF5
dhrYFyEv3WWsb8wK/u+NWIhy7ey9csMg/dQ6Yyciz3dPBD9K5Fw4AO13B0Cm/0zI
+uGzTpxQYV5HK09E03YbNAhRxyZty/3X4Mqw2It9d5MZWWi6La+GDCuAlC5hAc2v
Y20bpvhPuzvSxT88Sv4nj3MyiHNbpi8ctnTsxzYZVtYeeWsvWq4amQJGKX8T9yvU
QCIV0ychKifeAu5AtUVqIqdyEgaWalIyqfXbRiEahmnfKYauXbgFBWd4eYCiIyiy
B6+C3XQEGWuI8bdVCzFJ5H04BU96uKO+D1wSaQJZqDwIxZF4mK1iM1MeVillfy18
diAJdxEVLMgKcLqsnGB2X11YFEJa9vuUsHO075+UEB0szJnrBgebW2qujPL17wUl
DPzyG6WGBQbPozD5SuTgf5Wj/sRxWhbxIE7mL48OLjYjt+8AH/LVVh748fW0Ewfi
2DZf38ktz2r8fIMY8tFcbSMasgKVm8L/3bygYP/oICTaMK/t7J561iJy2+sk6Xxr
X93yWIb3QhbVefIuC8K4RrHCQh+uMXl/eNzlUYW8RkXtABWzPPnK5nVFsL5wcUgi
z6DnkfKFGv6GbbgkpFwBAnECLvtM50evwBfye3OtQ6A2sI0zE6VZ/vVSvbAV6qtU
/OkCOvbWJgACalvI2sIm8ft9/xnXE73lMizmZbpFKTuejxtd3xVJi5KMPF+P1u+o
pYr2HbqIBPlPmy3cgmdr9Ae7/MRck37M4YrZUCdDSBfjaZcjy9Dwx0WlC69BvsIA
iY1PhflCtPTGaK9b4L3MbWCEY2hH9zZfVxDjI7YES4Pme+t/mTDxdhk9SPe+fMDJ
le2jXbWnDnJ4b5ELxuKSGihV+vvL1e+ZJghe3m3vuk1TO2lzJJO4pGWZXsRTtNyB
FVR4dYyx916S+pYwF+MULZ0muKWxGvMZFK/Bok8yaOLMDSvIam3+AjoeflkfXJP7
AkesaEIndhUgzYVI3V6sq1LoFwtoHB3iNMwYdfuZcrbiBSE+OumLMw0t9RM5TRGp
O9ADxI4xv/GatbFYOZ2U28D8zNjHjuQk19wqXrEfECXQrx3wnOyjTNIyxCeaS3HH
NwdPftxZ1ikePMIwfMqtRpiODWMzqWa90fn3UTvY4qJcrqQ7YM4HWlGAxCQV7WfY
rLdFcRJWyvxUk2BRbXyAFvPhV2ZF/oMWWbyubme9Bg/Dt6MZa3xcWRvqBMIvc+0K
LVAF8304LIbJkhrFfxpXrRTKXdqWfgH0JsiLYE+X/+Kr6z5qWGtP/0fXBOZ5UNTA
XG9TsSCRl7F3d4aGXXeLSADEX9heM3RZc2vZMVyHIbzoaaNqO9jgK53lVDlsoxOc
91bc4n6fsugAppW/siCepUSQHaKLdHETSiR1KVsrcJx2ogv6dxS19jayg2aaJUC4
ti0O7RTEealzfO9+Xa8b5hrZiwWUhfYyDH0BifHW1323dl5IE73FRlgzz+4QFmx2
HwjUgfI2P3D8PYgk2+xdJD41td/N+2kX0deZHQBMpIHe/PhLuaNhIg+nzcuQ1+3A
qyg5jjjGXMwdzQjhjyXvY44QAvqmd4LhFg1FIZelipIGZPexcmUFEoRklg2zu+W/
GBsCQmEGKOsi4uQMVtadHiAJh0jvyIAyZG4sTNPVLSxF9+OjOje0FKP32n5STiqq
5vvnlRCZyojRSwGykwlYq4YzJYk3WV7TPNf/4TBzq7ESu86boXsWT5uMDgLystJO
j4GFKQ5XDaNrjytCAl5ucSAy2bvPcT59NeEyWyIdpJuap2SS0WAdoDjiresvjjkV
VXs5jABqTFcOTjL+6hM61WmZN3vgq9vnokGQYQUPrU1njLmSuejR12CQG8E6Xtdq
S240aBIKqIXbHuX2Vm4xTf9yTnEs99l2i3jKKbIdW2v+ASv0xxF8ho3HtK4lRih5
WLRLZpWyQcUzPCSiCHqBkPAsO8mauLHf17AUsWlGWhHhmBcvb/bgQXCpOvwTfTK9
X1/KMHGCOk3dz4AARKdSCuYcM/y9ArwrxJxrpELaNuAamx80BUoSnVCmpBgomZKD
dpsmEECyySRwhZX4Ur/3CVc849EcPlH+2PFoU7ZgVw3VditHEqCPnul4qne71aNM
mZfAJWWVJP2B9XlVptluDKq3EnxJ7Zi2jn/TqeOmmTrM97gLpqUct9yJ4oPs2zKT
FaXD6UwpUMthdcEeY2SbFO8rAIyLjuLa99RZGP54RDlbzybj+N7ve6K/bwF7ujjC
tSoxglMF25jdsjy8sOEGnm3qOP/Xrso0ufamTZha0zoxX0oxkfTDnDFcA1YjNkLX
dbR6FcjCo5KuplJzoTQOhhfd5/LeolVl5okWpupfWb5caw9etzxUHCNV8QFyTaGa
0D7DOjDz2CeqWFVkBm/MEgpqUCs5lat6k2uiwjntxRC8x2QHTwtqUa08rSCdGOQR
Vy4ckECZOgdIW4jQmGUD3AGpffy7oROXlgcpDg9TWOzMpltv2m13L1a46NocEoxh
+6Ax7g7WVlfWdEkNPQbqc7iVtr8QBBPoUNxInT9hg30uZU+nLNPcT69DyjzQvU2Y
y1lfBk+oXsZ1obhTVX3wSHneOKwDy4n3eAmT6jDyZsFmectzsxBjeZsOxXciECD/
HgfDgG4Exhsd4LkUIcJ7tVhI4Jsef2iRLyooG9RQmic3w6WH1ObvGvXZUgXrPwi2
41IVlMncX7HIZIz27KMY3rzwWErr4HyN7dvJDn7yMMKFqvuO3VcVbwurEP4eibSa
nMy2YWf+P4DYTQERYXSSINO7ZnttYTFEK+gonOqLUCTF7dFmEv7Xy43rfUYaPHct
s/oFObZijwr/W5V8ZYlFY+VNslBk5EUwl8C1ehuzMVpZEjtmruxLB+WhnRUHnNS7
LZJUrRh1JULeY30/L6qPdbII0K2DIAWfHJFytmPqNFUKrQhnWofe8oHd272cXITN
FiVSazf6pQV+lWRNJx7akDiVFV/bS3Zq5kqdUt7zGa4QM5KRKvi2mJ88bkqjllr7
FGYDLCNr90pgapI1JtPNFAaS1DsXqWI+X/ezk1zUXbIrlAhQuczLrOfm06rCCKDN
aN6s73/lH+kJ8u4FLeS64GjvXCujXsW1Z+0YCWS4yUvddKFE8dnTNVBDA5HRcuRP
82ALQY372Pn0oWmnV6goSXONHFVlSzhLeRCTX7O5lPdUMlNlCZyOiI7HCz/rQtub
hgVTlZNq3xr37aE9UqOmEaOkRWrytsAdErlN9Rm1gdbcPMO5NOqcLU/9NhNwK0va
wfHE1QbWDMfQXPAeo0s4LU8ZDt4ve6hDTmi+7RJtQpnTJyls/dQ+Kxle5bQ7Fger
RR0cezOz/7ZuU8zbhaumBgj8Zqks8oH2njFx9c18PX3Z44B2ZTs0DNfrTvsFPctA
yzsqIBR9fV/uYg6C4RGL3Oc430Lk+1n3TU7kcVTYdvA3Q7JckN6b+soNbOu5r55m
8QmxMXf0Xbig6nItASXMCbV+qQJSxRtdekt9qiqZbzev5aQj0I/hjIquzTvL5KyX
MtRT3/BjpQZOzB4EIkHrZ4OijlfT9hPWiDoLGNLsO6WYjwICO3crw9mvZqQU9UZN
DFx0hxgLqnnpd4NaTw3ULcQgmL3QNZfwNH2+c7Lznn3iVUDD0kpYRe01KmZoaGnQ
02dOWKdsHSKnOGALFisxHTA6esl335TmxNgriMFlUL7uJvaBG1w6BFn5ew2zpt0G
eAvzqS0y0GrXQleSAIsd7Q3XKjL3HZtkGw4dixs0M+ypYCG4SE0oP/AI+1jOwDg5
uEG63L1sN8o9HmWuKWDOQ/CO4d4yTnT1353oI4erKry/hiqw2wUEFsWI4pWNxmiD
xULpmqkjF6ZtuGlHwnUXly6g696gor+Xa9CyIqFTt/vNuzhQZxE9MwAoP2krYuA5
DKXKUncbratnMO9S7wzuWcOkCW5Wy1pkjCGpP34B5/HmVBAZn9JzPXg+mhKKhgv2
pJTfyCJoYq3dVQ9Sa2TYQYV/alAGWSPzYv/UTQLoTRpuesIUYPPRceBh8yhqjGZt
SVG//gonxVnt7In1Vk3fQ5voDkrGEfihwd99Wd6/r0DONApCol2So2ctV1jlXORL
w3W3PQB+7gDtk5ThD7qnAUyDKbqnUHIdqP41MnvLLjARk9uAphgBXQRd8UE6TSn5
g/knFeK1gPQBYomi5DHbMBADEwdyhxPwC+stfyNOEEiKJ4yi3SKjGf2fX3EQE1nR
SlmZnJmV8GTf4PzbCMHCT3y9YnHVAZ1aLPUPYb0i0kmhOlF9jmGhGmqJfQ8U2Xbc
0Mdo8Qlu/tUMkmgfdDGuafAZmR5Wcx/EJQookFejmB56iNOTxg1XBXDj1XKP+e4C
oohlDHNSiHS5nqfR5ylSvwbHidVXWoLKrXtCiDsjxKf+UyDk1kOAAohIstWGBfa1
S1DsF92xtHqimUyaxRUTOpsTL2d2kp62IRy1+TZrS9aEdLLNtYMv/5rh6fF6gJ/A
bfVTtOUKrp27+onkL4wYi3LQBZ4uxx2iA6hIRrOnSxietMlwM1iw3DXgATFO8DiC
oE+psN3LB5/EonzL8erlTRr7hay6uTYknNHfTCMl4ER+QXJi462FaZyk4wNx5e6P
KMw0POPBX34pj2fuvLdqfvtnDhGzCW6FbCOrh9TcwBkiUnmIkJ8N7+tDqwFXhZy2
ZjFedK+MBc6DO2nUlwHr4/IzcxwmZvnCRU8Mi8Bt9k6U3VcguWlLn0TZZ3k+VLVr
byN265XUiMUp3vkkeSBFaO3L9gU0FC4Oq4hIQ6JLB6UxfbtbEyY0zLzBtJetEGBN
avEB60U857i+j42qNhIJrZ+YPhLRS69TOjnvQmpsfjMb5H7OJdPG7kOjjvKGwzLP
AoV1eh+uO+YLbikqsmWFkepp/lyy/P6otPxPQY1mPPzGP+tnKtUG8dY7I289K0ib
2lCHGOrpGbza9pJpJmQ8qPpAEvPZ11cX5tyluzVkdQXI9/9I1zoa8gooGnfradGO
9yGs1m/kEsoJvTbF+8tI4N3ZLi40rBTDCpyDm9NNnm+L9WlxsReKd+Tprtu8V3Nn
fu150tY4moa/tpnZ6ST0NNb1C1n6qIzgokmF1kkOA7KUfYrpel3XnlgtY9VAIjHC
5KM4OjyfPaZkOh4QzAkqx/KJcxGWs56uF2mUOlWYYSMjvkiQ0hZgkyUnj3Uw3rss
4PWnTqUD173tB4dhhDUtVjFM9horySQ5zHIUEhg/5p1wMlA6GwKT5Ne1+rWQRZFr
lhy5zQBJk/+NxHS43ClKfG7jvWVMHuSs5o7vX9QkimKln5Tf7zpOIeho6yC+Vh0o
JphSaXMfZMrsJL4LN3kkZSqftNV311NADxo4BwdlWXWBEkUfrXpojJ5UunrjhgpN
K0lGIWlbA4oTQvpCVZxBWYbymWvsRfXJFq6erzVBjhr9wLGXkw85sHDv5nVjvO28
gEcOH5nFIAPIE1uCGYKtZDAealbCxVR7m5B1C5GhX4+d/CoI0IOwDFltdr/K3lN8
Tmsxl3lpM0brB1ma3312/Q1r/dzT6MA+cY2Qg+PQ1ZpdO4d3iJHsE7BcsQF07j+q
pizde03NGKcLlqIS/YP7kxsN4z4xtkyvq9y3+drVV1V2g9ZAZ/pkxa7ZWxkN+efr
gpmuMLuNcp7g3PzBTUTxX5Be31l7CSvkDQ7kO/XFT4ranJjVI2Quc/wIvDnSW83c
Qh6Tb61wjuRbQKyLyDSLERPkOmvGN5tNBrCEeuOzdGJu+jw+KSEbE6FH2vLHhYEM
/IGEZBhTPK7Bl7j90NdFF3BgNse7DOda9q206por783Al1wwYra8M78X4lDbJJEH
E8RhngTVx4yQHFLaYZxTaV22JVzBlrMTwTmt/mE0RC2o/haIy+tW0mymo2nHuiHJ
BkxV9mFfpkXRdigmucZlXzgYhRRqfuAF539HpgGTtFc8wGf3WYf6pv4pKdXTbE/y
ePuxoDsSb+L/LE8eQ6ZJfxD6IWLcstr6Bkp6PQSmKFhCIs67j7/s8L9oKwDy/cdr
GwMkyF+urAxSg+NB4wMeNz/+rDBZ2oVuTSlH57bvBvODc5gFpOjILOgIkxSjR3mm
6PX71Wmcr0E2fWG5E/7uKWymVhWnoVgEAhm1L2OlN104i43ca1rHHvc9Men9P6pd
5yOnh5R6zOUNMwd2jfsQWUHh0fZiuiMyy0M//uJz8w6TuGIQ6CC8nrD9xvKp5iwj
WY365rCA8trVtO2Lt7j6sUaX57rG9J7QOeJHzA3UzWT70ATzOTTkuuEtO2Y91PIm
9+SyQCcqPXMAGMU0kowuRIjJn3o0oxZ+DNBpuAMICu7sNsKbmTGgb0GKCUG9nZJy
tcGaDIWyZwO/3VRIb2Zk7vnhyzk7WbDS/l6mhpamQxx6/xZYYHqYgE10tQ4gLTWR
eYwT6YUxa9FPoy1+XJKeN8EeO9a93ISJN1IkpthfGQbfpcJRd9S5yR5d+V3Qn54g
YUd1IrURwgLEN2w2KHTw3t8Hykw4oK1exBIbbmYeU47pRD4Vnz1iLapjUq3Vs015
1BjcCWcmdIDtFwF1ojEKadWUS35AhCy6GHHXqpSyE4fcLmpqhVMRQ5+a7sgprgSP
17b+Ba3/QvxPFBWnohzgTcdSRPN2mxwcXRByKt7jwa8SjiqzGedDDtqoyfYqt7pV
UPd7fQ7FfMeOI6wJuW4dP93hMNo4ToZ47VmMC70jckxX3ZZX+BY3NPyNTU1xrCY5
o0ngYzfqkQUFBPO31KTdXiT2O+BazmDjqO3cyflTxGFYO8PeaJmr+R0hCJAVs2x5
V6jJ0UvRfI0+Zsi9vTpY66cnhXzGWGnryHCdVfq2QG+X6nJ7iNewb3mfuf4Je3Uf
jl9RyKNbE2rDw7eolgtaB353voFduPpyN22zbDCAq7mjB4A0tTP/WRELk4RQw6Rt
eA/FOgip/0pNq1eEEql6DxwGHwivNlmvhw21Jenny+z3SJHg3LS1qt1FsqmE3h3S
dd9o81La3RsXTUZDTh+btKw+FE1HPwmuJ86BZrt0aZfWkQzDuCMEW9cfuBrUf9YW
C02veznopV52oE8yyZFOenCs0ey6fyKmXSM/H/KjeWnfTpCrh6GndJkBIXySgV8L
LFLN+4jcB+YZV6BIh3kuxhSV2tDRO1xrjuy21s3WWZLFDsnM33kfHWkOPKA4mA4f
ei4RgV6uK9LwEgGbaTiK1sxhQmDSufeQ+eP2B8mujxE7SEAbbJB6KkmbQ41MfpnI
ROZLVtJiQ+G1Nua8kZ79bYOf2XJ3ypwVf1k82/W8H96t5bqDvL5a2ibNf8QsonhQ
Vi3NwZQhMjHRG8ferfGI6SkhfTH4OhRmcjUuPnladb0BmizI8zfijlHAqNiZHFEE
y0pwBSE0AmX7NDak2OTaTUuGoxvk9DGEmx0nyeHzFGZaxJ2a7sAaRLj2CUGqRVN9
CN2EOpbqdmIwHrHl7EDVRReTayE+1Jei3NTYBBTOVtk7I8FLxGcvk+9TDFFo+RSy
qbajgdR/DLc34yCSL24iPoi7dYM0LZlWHgAKVvAUB/neH682hj4AShE5xIeVDLd4
xIkibzjd2Mwt7tGWjj/cBhjdBAkBQ19f0H7deILDt2drao+vOrQS3Uix3kaB+bH+
KWeFswZeKOmDWmMI+ltCc3b9sw1q+p3geFDRW1BomFTt/ZyCi3pgPmgC5GuuqL9I
sDXYUsQ3SNfFYiHkD3Cpowxdia3+ljbGwh41JU39ekPcaPqvObEYVM1goLVToEss
TYtFU3JWga1YFkgoQTn8G+jDwE/Jp7gYHwJsJ26JZXxAoMKjuVYaHHhy8SvO+vLT
EAdj+X6gmHCXK7Yux2XqqwfSqeZ7EzxIzj1B/We2F4h5Ft65z2byCd3EIYKIqQhg
BgoX6tuwAj1J1vmmFLKYOccDBPmIEQVcuYQv9GQrWTUyrGcIq2ZEunlafY8afdFo
DHpHHwCsCXNk+R5aWGaRFcV6m+YxovwHIfEGiAhykNcsAut2btYNk7woqJ3aAFol
fLsf0gCbJ628muHm3a/YxUnXZjcukP66EUCayZ3yZbW1/PLY42nvfj0Y9nb11G2w
wrwyGEnjaV0jmTARigcwkkp4CluhrCXbbdHcB2kqHnBz1FKFbbhox1Okr9o/iaqK
rwPWoYauT9xOXQCsqPjnPLUXtMpCP7k1gkJaXesl9/JBOTgL1Oar7DraMoTZ2ZeQ
6J12NKcckYm8tWp2IuZ0F0nG3ZipNvsVS064ncj3ZicEptE5HqsI9c2Rs/Zcfv8Y
xhwkgYJboQueNSc+cTBTBg0DX86H9V3o+cC8asX2gQLmprA6JBW8/MvLQ8vMEPVq
XFteSbe+HBCzoGOCrjc2tav3G0bgbzifAeJCXIqlrP8MphwGO8pIeMXddBxAqKKN
Ipi12XNPrwY19m8BohFoSBMpm/Kx472TVh+375mZp0nwbL9y1sVtDeJvKQ13N4DU
KFl7221kHpmhMUEn1qUPWQKV7RzjCfekPRjtLz2zP9WZMwYcNH6s/GuSfxoiFlIW
3X4/ZKv3JLG4p7ryY/OrsczYx2gIPzQ8HxVolRYYNPud5iR/UWrYNw5FZlqgOW9G
OJNp9ejfn+VEbkM+83X2LZOijdBuH9PawOzuN23GvWYqPVPLjW137joDvEW59KeX
GgwRMzMDWsREso42aIHbbFo6WzJ3nrlTu97Pgx/OLjF5s7EJJ/BAIa+4AH1Yb6Dq
GOWQ8fjEhdv8nV75haaOKdUVsCNXhGVuSnq+pAVlgSrUfzCZsqrF8tp6XgQ63Bht
8cSgyJ5VcaAp1MC/TWQou87i7GMYpyLPL5BdsnMhDU0OtsBOONCVC9DmVVYi8wtE
fimip/0uQZnQs5xgrHMb43uNi5okxSZWGj8KQsOMqCnDT3kP4/zGdxtYtzlHSqT5
HF0RS4/BcWKv3qOzOrX4Hso6zxJJGHBJVnC0O6iEIGrjHsrUrltw0hsgH0YNA9Pw
x/NuKvxHiI24dCYISF9lSKzkppIL4qxOWW51VkD2sc9M2HLL+9CFi3CuCqhOd+PX
eR6AmDYL3Gk7WzV5OUMhRkOZaRHxFHrLtcZVsu+KRWOBzsE935ZYR2acZ4donYYY
NUjz9S2wPMHJlWB7+a4qOdAnRIJWkr+NAxpWE32VBk5hsgssCgx2HZu2u6OxRUnR
5/rBotA3Yvh27MdBTqpBRPwz0DU7JEt0JN509+nj1VEhTUfK4KsPW3aYXmyGmvpQ
XGZHnSYx+QF9t0vSA5LGLC0s3F9sdldrWPHRBrm2DLZDkRp6T369/CHaSap+yfQO
MFI3Z+wcwOWtuZTn0JbjjywxoFv+fFnalNPnX0knleKRaJsxac3k505TskELKSvJ
2XH9d5C+jPkxLx5w9dSu84B3jfE93sF28cGUoDvGMC6BEoHJz/CKoN/FLscxRs+r
tLKWbRdHvd19LGwXCHVFOL1lcSIEL6ZB+3pTIZdq/TKPIxfLI8TOSSzF0Ryiwkz4
6XBLVy+Bvt6mIRQRYVF2q3w97YsjVh1OdRdzmWYyPA8LhENgqlCYaUtE8sCQZdIH
/kmDn7CUa9uZhhLGx8p5z4fkj0Bzl/hkWilwfjzYKHmepD2hL7SMXaW9jv8PoT/c
HyMVRSTkfGYJ9atGAXfkiKoPQjnos3Zzf2BVTtQCCIkn+WLygm2WuwjByh+BtAwb
ETJRT3Kn3w1Zsx/o5w14t2aYOI0DPjRE8eqJPnY1mgiAmysMSFIhKDySAkg4zvjQ
+8ecEaAAo+hEaqqgg515WbisvgE38crRn7ZR4njz2i9h3KZvbXPivDoaAALTIYsO
8uzIb5qS9Lu0IqPLFpNEFFwGRx+RcQEf4Y8skoGKlmwidEORQfQvE5GQioYIEqWD
+c8tKup2deKhJDGIdwbNioaltqwSywAHyGstHbErHlnDYpGnO/fXyknIGxVlv1KL
NaXLDR1j3lyqpoNtKVFACUShwe17ZkfANAqVoT59YBsJaT/tUrY+RuMoc34THl7W
Ht6RIrIi1IUHMjDjq0l2GYIIPujo4od5yQxTq4YUG1ZsYC/GejntE2t/UViHIajj
MTnNZXSDH2mn7jqWqBXKmYtYm3e5JICuOfgJNz2w2L4jTa0ff+MfmVCNbHA2x8kC
ZDNpqSlNtvWUGC6ZFKDZwZX6Ehw8RZKltE2WVYq5cfSqGrBEQIqXOwDfYh5t9/W8
9X7lZbnAyE5RDLWfZE41VLPJia9Q/rpqVoXNzCBR1YlyBJLcu/tHdrXwRBxTL21f
dnph2kEtzIb2jgCIIWT5Ssz5wClxBhmqDL4yh50eToB3y1o6nvshj1rtZQ+I7teI
gWhg5W+pjLzI0Kt7czx6M+CF9XV+nYjQWvKIEmRff9itIk7W0RyCmdsyt0uV/DJb
gzuFu5DkKrcx6vekir9iOwS2PAyYFEpsU6k3ghqGfbbt9kq1BB1DqNecVTklS7at
d4uPwjB1yWE+0nGhbxafzaDuO2mOLi4rD8lHR/vDezOuAk9WhJPe4NASNDtKjO4g
7mjgxh7/fEEjR3HBM8OKgZxWY3n3OiC/Ip+Tisimn3fhnzx5vWkheUcq5C4pwKZQ
d4uPNJhus+SLBcGpY6bkC3LzFV/Z1LbaFRYr4yK2BvtJ8N8mT6xnr3m7Dm9tof23
wCna/Z/KOVz+6yS1hP9JbAxdtMkxsh6b3Tetw5+oLvZssI97aHQYDGcC8B26cqP4
qBGVSv1u12kBiMm5l0OsHjYa1FdmsqL4bhSU0AHbVW30yTCrZAUPbCx/JU/KyTC2
QrisQ0/iKx0RJuu9qV1aX9ylfYF9O+ySYHvDVzFdZB7gE9zykA2uO7ejR+97UAON
EhggqaI/CufRmcPKvyqTPxH8nwMOUAlkRRNyo5SS51phstRakPUyrGkaGk5M3slR
V2cyslLY/tjoqF41CY2P/hGa4QaNcUgMB9KgbR9IRtU9uQ9CoNN6se2jRLi9abK1
7JXEsIL3a6fLqUP5Jv+DmOqRq8xgIwuNfEt9byMcfEB/KxUZMwhp/I0RqMoFWZO+
wOzyu1Xyd1oqPEpV4owH5hrCUl0qkryGeHNBv2+F704ludVJ47Kpx+SfUK2XjQYe
H10fnO/wvsq7P+eJ3QNH5+nNXZayy9cpBH2X2UDYs+3/P3DldfF/RoWzD1PiHin2
GD/3OUUZfRWfrMR5TE2lTMex8XxTTxCAiTjPgrj/zD5I3b+jPlA4i/y9N6I+yhgK
4GFwNKqE0xUQWWAv3bja0jNQpXtRgo3DnBt4Wudo/SpwTKxNe9q2BOTOG3IN7aW1
lveiPV06+c11ersIxaUDVmoljxTSsF8IvSuRnvUaDJyuxm5KyjDoKPIocS3r94Fp
fhOkb3XtICh4yDGpT9OI5AaTJoxKe8tc2cXlGupaExNCILO6cLo4xjXBTGtejsie
Xds1nuPSS5+cpmE0jRpIy9x0osE9zRUYkTEw6r333EOz1+yMewwBOX8sxBtMikCZ
+uZzoghZZjZQY/O9OkvdVjcHmmSpFhTxwj0MTPhwNjq7gbyUrkxyTgVQ/NoLdGUu
LtJelqcoeM5bhHv8eDv/zS91A1QwZcLiZs0FVJ5pwz73R0VPTZqdlHIPp02ltbNT
j6tBmNtpbgV1oN0PUKg0ky2wsjwDFJwj35v7bAsoeg0NpPGnrks36uKZS+gLWeF5
nw7Ah5t1PIXEmYgyppOrnyikqwLdIdUoGu7AZXr3AI3QRVdxvFF7M4LtL5dfc9J9
LYwB7qy8UqlrdJwfjTy6e9ZAU5lOXFeAZ6evIGK6EmhK+0+LtIZNA4ASmhGlPyeL
BY/eQw3ANW4Fg0O0clPVMtuSrfdV6RhY0L8VvnittN1FRqkXPjQ5b+VygkABPDSK
FIEUQX5EUZW2kmQMcl+MnWLsedyFes/ugxkDm9vnFLx30s7HNu4S7SXFTI6NAFQe
Q6C1s2WkJRgxv4axpnzL3uv4FFyp0JVUuDrn7mtAIIXYUxsx4w2WLny3/8+vUHIt
rlDmyOpRZIyM96SsaPNCiFo+MXmp82rrab26f9vKH1PViMX9t/mKufdZALY7tI5r
YfTQyTi89VmkBq5U8GXHamYpXTJFeghapKirXZuGPpUMfn99Vnr+z18T7KUBd32F
3IqvjbgtdAifzRt+n5/mAHBc4/5LqFBOw9eoPlQoZQ1z2jXfNFCkKPzlCeSMXF5f
oPcsI5h0Ue2d3CiYpwkF/kKX42CvPK1XyzEWRY9/3tlK4ulD19fXleteGkOkaJt6
xSwJ3HO2W+m4Dvwu62O9hLIv8knDL2nO78+OXyVjWdifbFdRWzLY9COegIU0fK8B
1RoCKd6HQRIURKuTH9ol/uN32pkasJ9E8/VkZLfpgp/0BmyKg5fl+39nwGWxkl2f
JyfQ+KqcGfO/fdn8wgT+vOShzBpS11+YQgBmXCISGJUhES4ei4lKdjU4elE18p/D
LDWI67yJVnoNDf90rrviHBKhYU7IS+vCQ3Ajgr+fwo1gTHtVVinbKxm57iJLu2PL
6XbaHZ0n8vOPL6jHYpNBMGY3eSOQ+E8+3pBIirOnmeo5j8CxorL6Z0YXrWG4b8Rm
MvCrKSTQHMTBCmObyZPVtht5VEicD/x3aL89MxAObCRcMPSBwBweW3pjI9/MkjLL
D3lglY8JR9nnLe8QKi7j6/n6BnU1kpjC2jWXDvlkM4+QkJT5U+2oFymjxidoLeiQ
eG7AlCL1HmMC1Mpb74f//SUqcaKJc0rcuf788vVH3ufMEyAwIrReGuGCxJYskKMG
xoZThUkEtddQQ9UrKESOdYqw8HZ2WDuIm+ZjLGo+Rl2oHuLa0/X9bvh956USpdeH
x4IUqpcgQ7nh/2cugkYTpQq2MkeZRPC8EPwlzWgLaw0dI2T775tkl2A9e/l4CIfb
SjasOhMk7riRMotumDWgoBO3wiFIYMJAFqgD0tk42DLGu1VS1eaPw+rCKD+vgoDt
AiRvG0Lbpv/MQGpuNJY2Tnf0nlTgmfKCj0dRDL9sgtu5AWJCfK0dYxz301WHamsB
Xg+gH0Ec2T6iN2UBFbIF9I/7BuIrYy0PV2LZLZUud4yMtjDOyXSVOu5lIICd46Z5
qHxYiIj5+4JvsohF9bXA3pIcucyi0XeognxbQ+SpQaKaph+egFixVwSG0exGTXKx
xLpWl4OVbV/hkFMz9Pja1D0JDYJM8/6uIbWP380wyXxdhyT2zWsOLXmWQrCkrMl5
7zUZDQMyS9y/YnbFDch35zUPt6hvS25u1QOty7pLqUzedLX2q9aYHLPA1YIi2IKf
70fvesdE1kyEeGo3JvucNuf7fIiLUBfP985ZOLwJ3EqMLUZY04NPkXhBHFk28euF
4pZmqMu5kpp5CaJglqn5eUc5kRQS9WL9RbXn361rkSpK+dm+dCubgwkfxxHv5elE
YDVdNY2TH8BL8EcZr6C+1aqCEIQeBJ0LivCBWO81SrhIyRKwTLi8cviOTUR8U0tM
1mN47dq8ul7pTOy3nnCt+wYHMl9uLcfuArzRIAKg3auYgODE3Tr8SnVmWBt7Ovr9
+zn8nV1rogxe1R1YS7UGp2TFB7ESJfbTdAPiQt+FtEVI5chIq9BZb6EzQ7naWs4/
QTarPt9OhfhV1LsdG+7pjp1f6jK2W9nJcHzmnDIKQ8JAYJYuCSzvuny0WoiQfOK2
aAuaW6UCHwLj/lYaLjmKqgcpg0HYe4EDUlDp3cAFs0WAElPS4cmndMXBJqXvYPgo
GPpN3qUunYUz4j2HFXZdBpgFfWyWKIhT+fg86dj5Qrg4ZpHLdsZMLuOZoM1+H7rg
xeczKUDSbUDaEd+fTUv8YILSQtN7P1xOi6byukv9mYN7bc3onfZQK6NUWoNmDOhy
yV6updk8bDNqmjPi8FvojgvkLBQbPzQMXlcoxR2lbQsyT4xLlo20vbVPp63UU1aT
uBHgK+boQqyVaLo6m2Rm6WsZ5STuTkpkLs3eyLohAgUjz34JvWcGQjgsJACPdHF5
eK9JYu0e4A3UJQsr4TBb4MXH4xD8wYwQD5jCJZhJS2anSYJGp4ZVWkcvs0iovohi
6OBQNwTIx9uuABFxedXuDyZmJIosrldIi6BlMtW4O528h9JQOicHNaHtbOFUrfLh
gymEG4ST9jLBE0fho6Av15aNsUPUOojzreEpOLWvcMtT1hVj/IZ9FJd2aZSDrecv
5rJRCqSuHp/DLW2IQjhzjKBcI1h0YHLVc6VXFtMfAshMxhAxu3YunBP6KT3pyzUY
CFGpcaYKIf6TyxAvWSdT6pPZSbOUyX8mAeN7v9Ri7o9Old7ixNYZg4gVxsb63prP
AI6jAf/YYBay6y20hItTohp+5eltXSf1mBrgxmrvj+4O7jSrXeXmBl3lK+DCLiRx
I5cnQQP6wctG+YwvDtlUcrmdWRwIzxK3vwe7oZaWEs+v9C9XI+a+9vtJC4Coi3eS
jy0GLCnJm22O/sGJQ0bl8/9qJ9ycBaELew1mcQwfGBrIjtmEaavF5xOuncpQlfYS
YDa1IWZm/doiezY2JXBrWW8xFd9KlSWc1wpMD3MeXW/y4dJisSxGmwXiQ4WvlB38
qgVfs//GU7Jhdx/X/Oni822tJUQpBLYLzFjn+CTddxf4A2L6wAs3V08910lmJY+G
NSIjGadmMbjRV/W4yqa6KpxSwelxm/C82+6zAWy0w69fgzZHwRd1B7v7RaekrIHh
A62aIKTHkcyU9+V4dOfoVyImbOeesDpppJY0oB+q3p7Rjs62nimSYvlUBbYVSEhy
A22+pzjyVMJCoI7IB4xwCBjm3kjZzu5NBgJd/1OS6RqgkZ+3FS+MqFPP5ZPCn7B9
0KTzmpMKpnvu3UlFBwQbfSGuTqnK6jNGWR9nqbbhlbQ+yHFDKn9YMkaohBUTCa2N
HI6yDgUUT/LRJArJjwzrEzOSuGt3ewlOeuN3rEJdPyseZL6DBRxfqApwEB0AG7zg
1gCR/WcqTKjAPTbsuvxSZyHUL/QHet2Vtoi94tslVtykQIS795xkd/8vKtw/nl00
u3SQtMuaKtDIvHM616u8M+lJ8uM3vznriSdzf9kzkIatW5SBbwYbQ8YOX4/g2kqJ
zO8J+z5X4reT9H5UkWh8cUvBb7peyiHvqPiK09+UYXFZZJWq8+QdAHlQtBH1uoNZ
RMrjsfvn3adRBYQB83ymstJ3kryCcaZJ+eL4ANgFc+CYvvbCZmTMbIPTV7y+Bcer
Cscxjh9TIE4mJNvV2+dwho3eEt+Z/6V8X5QaCCJIyOcPTnW5Fs+QIbJVtIpGFGhv
m0V0t3aWLUPVV8fXNwBd0OHG0e2DE07mOVPqSBdqRhb5JodpNSHzuGemcg2BSDAv
LgRka4qSO31kaAkZ82wZEsoGCLg6AYOSFCr3kudPVeqi4Mg7ZXlpLjJQugZlwW2x
JU+v8aT5OLjx5vkIkix5IIwZ2OZHLGmNee2RXTxvQq16urQ8Y5E8WcRABIZenyS+
Qxn/vZRU3PZKsCK5UrdZprvZJLUFcbQg+HdcySR3sZYRvXaV0crMFjkpJ05qFetd
JbWpvJ3rEnVB971ExI14/jKI/qblCoHWuG/lbLBqaSrz9KbrVJPm5XigO9eBJayv
A/5g5JkC/8CprxrMSP0Rmx/yi3O9lZnsBTiiLa0psCDrgUpo2+56hZyQNSDDuX9u
7t3h39r6b0cGn0VOXCwEeEpKJcER+Q15sjIYtqOunY+5U6pxYhdo/B3R7lPUA2jN
johYTfeOK7meeLHweh5KMftyN6ivCjt9dgRRJ/lrgd3c/PrhvYSwDH3F3Je0wxwI
rv4tcMDgrZNQm8upgYoNxz8efGYJwauY1fvRyQPsP0FbL6cOsG37XxxDWz/bwBsA
42PrZECk6exTQIDZKTpnU/zBQAVdOG5l4yUtuPIgAebvT1qlRGIprwn0s75rpsxk
YCTmwFA3MQY4bMmILyQL1jb09NDAqtUYUASEieT7WksLLcRMfy6V1TOnA6YvpQi1
b53SEoeM8rHaVf2aj3TA054kDroj4+s4ME6D1bjFqfK0PM+0/sTQg/jamTV0iPTf
r3xkP1LroAHPHYOK94AUfWNksLOqIE32xD7agUgsRN5JZghctu2L0zaGalnHvk8V
skxTg4W7SxOqNpBWhcDSIvIj/DbTwsFUxVUSsI+kalHDvZjoQxd+9nZ7x0g40Qc3
JaY8fJS0NXcGLFgNdCvNmar9443TqNv75uYOAwzxbcuDexnZMqpGwerQYUhjrc3t
2ZrNyM+QvRUP8NDTkc18RnHXzQkSL1HlFb8fUnLsCYERr1F8XVP6ARhoHD0OAsQu
QL1pSVH0mVzuzwEFPyRLcmIXXDBuTHexbxilskgxBpl+mQhBBX5NIRA7EZA2qiiP
clDMCk8+CtnnKmvzeokCizAr0J7Cowc1ONpPSFBjP2TBhHpAsKjdx+yYK13aLqV+
fz5Ddtv5xACn3LAJhoE52cKGeBI+bhnAhXpOuy5iSDBWSuiF0X1ApDT4SrLYPaZK
wiJyBtkL+fsMdNsNbfXRRsf5ysN6xKQTAyg7IZH6+ebNpTUsirm3tLoX89Yv1V4Y
N7lLJ5V0vngiB4PUJYH3r/cPBC4XiDtOZ4wcW9tGPAIVCUQgp/5xCDB77ffxeI1J
dL4i6p1u/YBJ5uvFHrlk5awbhpfhQzGoG++Z5jfOvmpi+Pec5mhiPycP6KxTNymS
wpRhu224/dGOuJUuja2jzEeur7jlSIQq4HCKpub7Ognoje66sEqqS8p5dDwx6QC8
Hub2X1WHWs1iiQK1x1nd/OqsZ/G1pjwiAsogChuXewyjInHfwRYOxef+5J4aQR4v
pacaQu9mjKwisG7WsEDEWoVj4zLwI/b5bYcWMKsami5502YfZW7Vd1QOj/1gQYbY
GeMKvsKfk7eivytTjGm8L9F0qmByPuECQenKDXWBW+WnmKuWbgTQ/KYRhX9Dk+PN
89pjl5WHFaoG/9uAbSMVkogNbWLzwTiMBi77Ooj2xEB3IcCeA/rX1TkyZQNV5blQ
m6+NSmsAhn6J991TvyK2nH2IzrSPHfYcgoypqnI9Raoa+NU0rwd48s7kfbOUqQ9b
VBrumSH2m/YpLN7xmiS4+FNZvNcTkPe2mSipetMeWj7eQV+8/REjclcUG4CyYDYA
79PsOlbZN8vDMV9I57UIAFnXaCKpJEQcx34oPt9QzQ7DWj3a7x1JVawggM0clsfw
UBJAhS5WcU9oHr5nFgizr3aK6FvIn8/bixRPTs+cpJwbMBezbiEm6eWsW8mue55h
0RSSQeAnXWzj8GY1UDFQDkKkzO3p5XZiXeKOfnQq2gCrVQ4vPzoDhxrTGBiudxsh
fSBzjO44KFw3JfYXoPgR2ceJDkD2+ukriQHYdzbVfpkeJCKQOa+a1E09jmMy6CUM
MHFIe1rC1jmO8xIu9WibQE6hcH8I3QLw20UKf6vzsq9avtAnfy0CuQs4H9IfB3nf
tkhpWqbDxWU2IWjnHh1v7AR3fxTeut8yogUmxJVZcW3akmLxNRCmVOwK+HjQJiI6
PCFJKgp2XOCgbFqm64YdDigrlK1Xj93AK0XAHoJHMFq+7ugOIO4OyRHpltNyKtV9
yNzFXgZCOvWmf9Jo5Z36DODO0iC1dnZge6TwPk2+fQ4R0slW+gBk3T1H9PXGDyCT
o+iCe99xwO6URuxbzKbFraC9ZH15Sb5qVl+/CwTpXaPqiO8RqxzCG4pS2Zbxk+kR
ZznED+M0816gQRq6vHLGS7W0t2otsnHbKn5q4ZTXq3r9o8ki7f6MBcseZ/xWrERR
wO1WuiAcocQDdmmarU0OPvXlX2bj5pao/5pVQSTjOvbuE1kMfeUiAsRXMDvhvxsb
JpLom3lnIVIkOwZo37g1rljeh22K+b+QBxOgNsuukLeZCCqsdauU8Coqjr29sLGx
sVVjXAIQioTekQBpZns927mGSF4grUyjgpWUQwD67B/dNDJv35S5lla2a4WJKldg
yfE726PS76N9W+oKmaccc9vNhu4m3t8HUuazB3tLh98wXct8ucfUUp0icZ9f/2z5
5Hy08riigiIKF+CsdE1hcgOU9S4EIPB2KcnM8Rl+XaxSGxGhFRVL3BFEErS0Xm1R
p1CYbG9H4PblqZVyZm+uFbSs7R+ZJ3K04o9BAccguk657XO3L0rEBBP1k1spiHYC
doSwZvbDupjDq6OYYlA+urXzDuUCVX5S+lucjHXReEu6k1u1hhuzAuQFQsVGQ2TF
eXdQXDZStedYnFONAP1w2uDIMYhfA2U8GyxcOhmzsrEaBmWguEzTkBu4v+vCfepV
pk0bZyPmLsqSl+l0Cheo4RHbF/8K2T3WP7q2SYdiFoCZE9JJA37lI0sTC/a4wZ4I
ayMMHrJF4pmbukAQMiYjb+PyKbObhMpuzdf9RrvnmdXvcsXmyo0YL4h+0L4o0ex6
nbnbQMnzgFBXFNyqsrOc3nDRRd7Cz/Ifp540Gd0J744mnsqJUz56BqrPhbhVtaBH
nCVvsdtskwR4yzKrMJzjl7UitG2uSh4vBa69lApcLvM3XZAUnmSB6SGw6g+DVfi8
1SLZ8pj3McBIYVfg1a4VjLBOy2s+H7pjjGee9zKXhsQ+R3e+axaommpWqam6LJ6L
Dmfk3Gg2130GxVvemCzY1+X1Cxx2St3JY1I7tC4j4ENUzycuwS/2LctXwejmLFf2
nQv+e2iasXNMUjEZrUJN+ro+t9VwRbRmS2yhtW4gI2MbNh+DMYHf2zvhcBbNQKt1
qoXDJXoc1VRvVoU1Lkc+vqDtArtycZpK9zgvEz4yHuxuDLl4x7XEC0wWXudHbEIH
ViLL6Ycnr6kCRCZy8aXyiNzIM+/GQBpAp1fCpEZUA6cqMztRQVeECUcEfrIITVh5
V3KljdFrfcaPdMZInmP3ggt7Q9Ff66p+cFQd6EmVbG0Bj5dT2NsDwZg4NOvgbjU0
5FyzBCCVXgFfcG+hYNk2w+rgVCueSNt2VObeSPDBkebzqY2YGclQ+7kFlmxUF5QH
WmReMHccJ3Ktk+B1mVJX2eJ4vuOpeEegS2lPPpAXugU9xR2d4C/lpO5r7eaKjE8b
5vXZ1X+TZftvd1VnR+Fx2qGVr+ZILEEstKkaz1jU2FCM6p6NxFDFZUdYTeatIqgY
3j4YQuIpV4c5MbzW2Beim025jRDZVOIYnHAoz1PrSTKGBxjqkNugi3L45h374c7z
Ie1kbMQCDmr7hCOn9ETD+3SX2Mx5ot95QxKvpGDUYhZlcL/uzWchiNxaFgWhV99l
Uhqb1Jb7E4mlxxTjFtyVrFHqG4BlCPvxO22h4K9yT070XDceOCSuup7xrHr9vKsd
xUT92FGmGr9W/noaSSwxVUEC36lMnjRb6F0KW0ixNpm9i65UG0JPeVC6wgH8BxLf
deCdwD9eIhBE4Chg6n4PJlaWi30ZlNepD5wNi+8BD32fEP8JZKzHaSCtdzbOswaY
nA/Ol2+R5AcBuLPWyfOXSMB3Uj6RgSJxCNewdFHwacWcQB/TsGqZZRtwzpXRjAIN
D85ii+SLhD5bl3s0GZCanc2mrLFEQYCAcTNBws2v0gEa3Sw8ltIau0aQ7aaomSYi
Xwqnpyt7DlkccJhrYWburevNZMWXOf3Jrk3CW+98Byez1GUCyX2DYRjScw/pb/YQ
ejBtuvDow7GPD5WIWjwfw5uLf5TgkVs5ZMKareNt7EDrJPUB923ZqEU1I4PsambH
qhO2ViBjfWAc4x5la7lPo6Gu4L/MfK3FHROzfJtIemsTQIGfKSx2ooAmelo0R8n9
fsIvnFC1CNSW1uGlLHZRUwIFaLDNIkLtIroVh4Iyb/7bLfdMqJSQ+J5bxmZbpQTn
cSg5XEIn2mj2bcLyu2rbv8xHG0NH9pYXJiaEwruTWDLRtjwWp36e4Oa5TwLaEIPF
D4k1dsqRI5BxPddNZMXapb98IvnFIgItt0RzAan7kHo0FLymba48+sQ39u6VeoTN
giZLp6I0qmY4uG/5gA/R/VuKIPm1cycgBKiPlScJSoHY2Tsm2YkjW94kZ2xfAQ05
I4IGPY485rIqDqoS18UoQblGQy2arqcMd53RvtNNqgf/o7ogzzh29uOQkIX94NpM
DX8HxKD+2obfkN905IxAtqIUIKGbnCMgE1jSIxMf5VeFupYYb0wVpMeyxUEZqMbk
IUv0sMKxvn2r1LBnkYappzkNUq6tdlQ8EGV0WxazGWfzBoU0w9KYdRYTQR3zChUH
6T0DwWl2s1w8kH5yuKQJ0QDYOvb4tSvYYr9Od91dj2Skmim7MDiFrwcM9qKGDBvR
XNxlkuOATwdG7ySUE0fgI7CbD8UnBaTrzQFwO17EXNS02iyUq52avUjOB1yfyNiN
BG8x77ujeAa1BuHCLMcOKNh+KD+4ft5J/FnC3tteLJHhf6hVHzz100qWs0geNAR4
fM+LcBT8siuT0EXf9Bhi1xJMiuIuqKrZHwSzME5cVUF0NZdRHhX5yXTBTu8Ylcfk
1NV3VCdeWfKxBa72KzigGhY/hTyMyw+xnn5HjS/L3LwxO08RuhEDScUbc+uuRubO
gey1Xow65nk13h94o/GRe+XQIC+i5zRIT21KOcyTxvTPHMGX3onDPYUhuf9dguoQ
T7yVaOGolqGUczS0+JYzRMGA2aDydq0vqopbhYxaKfV/YbSPJPJUjt/Yi0bNMIue
d+hjiF18XsufR1MKtyIAPp0v5e0GezmbkOypsli2N2KTbZ4tNGxIepK2kGA2JcnG
Am9C9+5wRPXEnc/ajOQ4+UrfO551Dxk5aaVameOMs70U+LgF6qHNEMnz7xJyrcYl
Sx9auJinlvg+0lCdITrN4KB8hL3XvD9j8HESpV5rFLky2eHv7ZrQr26OeCv4hyrL
NVlIBnNKtfboGVHbd1SEXq4fmBBCxU1BxK9ggS0bhEf+mRsIv9nwQx1kfNxxbrvK
9p+eAUrX5VTb453Vp4Rj4SCrLT5BMkUmS+PrAWFIx5Yr+jVGAAP0DSD2Z3gceVc8
7V6A6VLXgrtQxasZCqiNLt169tJM5F0NuXOTQrEEW6msAl2C3nptkHGY2uiPV6ta
wA4FrcPqTVNxUvxrrfXcNanjCEIi8N0IMkpvs6o6plnT9v/xgIQZgX9++w2TrNWs
wVsPEH/obC2i9U6FEWOMTJ89FFR98zWSla4VLMZ5UiAYwM16xG3SiyJQ/2gq2IjH
vTmcZ/YwASypFTyrnHqNKec/5atN7EOlggOKZ4skMij0zspeuukDOTFzCTnonlXj
69WGykUPT4yEdyRNdsKGp2+Gw7ihXq5jR+y9VUy0sZBtcgs6WiGAMmCD4CRVcYGq
XZ0aTxwCWGRrb7p3ZBouQDU8RUskAfefCZjwHy89W4wcB3MFxlcAbGmXd+6R67iE
+rJpA0earFw0rtGi/wxrxyjDVQSK4Tt4zUhT0f/VujenbVOnwL80bC3NBN11Kw/F
qOHr/NaEU5r4ONuHFsAW1oTnszImqidv5W92xl9N67eUdlDQUxSNGyW6Wn/ihgzs
QV3QqVsFLyxVrI9N1oJSC59yjQBqfNUf8k0owBbCMYTS+Rw78cqDj7dQaEVeJpDS
ApKvCXhguf1K/+ePjuUoxnISkmp7sSc07EE6x3qVOuFctouiZTNs8ImE/GO3thv0
RN/DIZkIsWYJwUuPI+0uR5jlotQquzLeVlJRAfkIFXwH43YjpS8KFs3ZfG3rOx7I
0JdN9VTMthe7RGfgVskWxoFNlE+nqoiY9sJ80vGOYDYSUQpnXEBm9INvcWOyWfC3
wb+CFKc72+UeLlzygiV4xxOStXA9C2TPuncYFP8TTY4451mfy40ZKWaTVt6MjtUv
sRJ6mxEISIN4pJ+xgDcNGcnVZbeTfQ8UXwx+DNzDmJoNcNly/J/sGGGntZlAlvze
Su28/01dnFCy/zPelyqTEEC2THPMD9xkczZrf1E+WEpII+zqT5qsoVC1Cy9VonNL
fyuRlntc6e1nPhqCkvpWHsncNjRa0aDpCWToSdc9eMtx6RHXNR4qltHDb+8GNlOw
UxfbWMkqNA4npSJ4XwQWkLzkIpDN3ctDICbqZO4LzVrCLbgtZ4R/M8ChYrDX6Iv2
AUfL0HnfymTSuMZQx+KxeRNLald5jwue/w+lVLdu0lSz5Rb/QoPsTJ+vtLQTigsM
Ha8gxbPVIOyXCSCIa4qQ3fjcQDAc4So3WrwEyUk4efL75HoZ1U9rjTdvN0HTh8Qj
PPTiA12ZlMvNXVAvTPBIfuOBhBC4kwpC7bq4RBJIYoMeAm8Px4CdUETYV+WFX4NM
fLay2gCjDSsN0VYH6D53SASAmxmDqyTNtndW/ycPPOTWJshZ6AAV4izESvdnEFrD
/B4EugZQ42JRS/YYbrywOoCyoO6rQfWO33vT7GMQ64WfAtCCfRP4vzilLo9sslEK
SQbPC7lsWjNjQIdoZyAq7AUz7eQNVP0DIToLbHxGMvHDZ0RzUGE3Zj4PtByoymdb
OLLR3JTDKnBmiYy24RlOvHkwqTLqN3gTCXce7SC2OBvwqdeOkbtmcIHrR9B07HFY
Ye+VtrdOg636zf3UOL7dgd/NRW/J7s3WMYq4BO6ak41BBbuYYIF4wzQY7O3jk1JD
NaHU/bvmmFjfeqBENoSvtx5YTPO16qoFVBt4tC1XiepX6fdHVo/QWKaqbMxmcb9o
gvKS9IylKTUR/4dCKZNR6g3B5ASzBWslz/HjoG3TLWhvDTxdqk3WsItrIk8W2jRd
8OBZI+IuVl0aoGPpBX6G/NqmyL80Vaeh8/Q/NxL0jFbxNaB2oA2J3qMQxAXJy3FZ
XFpQv0GFMGkZ6JxoW0GrC024dwf37bvUdKX9ajL8xmUrddA1caQI2a+EvVGxUYc+
UuSk7r4lICEWmODqmSrmVeLV2GFB9dDOcqyRUs2F8yMReTa4YuxBVsskcSpK43Rp
DZ46uOBZ1tlf7UODY3ywC0LBLBX2N4Zf5niXKKK0pkDZsRReFu6w1IOD85+C7uWi
JqObSRNcplKwnBi9ZMEBQ0W+PdRTeIpKe4Y29UoKIBReNnx1WDR5EaApjlnPh9sK
OyMPF7zccLE3JFdaEziZcLUNU2yXyi3gIzbyyd39BTcp2QjU9SE23F+IrLRlqHgx
8CVHcJdZTpMcnFTD3QPXC3C3soUU2aNPWhkt6f2PkzIJO94+WPfV7wvSHOBM5wav
B9CnL1uRAnqGxsni1LehwFSnz+AQE0LD4BHs5KF5DKxvcLeyiecURCW9AE9cV0EH
mGmPaGyT2fgt+yLNaj3m3dvgMNa4SGIccuKUaaS3tnQQpDJFy42y9qPPgEykUOjZ
RZ/e749aqeRXhRehWbAl51nBMA+MH3RSiyYoGnorhD9CdZTFWNZhfsT8rukar5+Z
qthyOuSoTWYuOh5tLtuQiCj9VNjoXhRc8h+wj7+4B46usZ5KFt9IVWnVV2h8EnAe
x+ECvhTxMt3Dg9oZECDlqNzW8rReQ/FGYENDVYcvyi6+TXMzvqf4qGavQ10jTCpn
gWVEIxiia2/XBeV+8uOnnJJGSNe+U39Ve/t2qyHC4Csx0I7J+izQHRx2lazufd9z
Ut49BLhAZd34TK1syYgCGNODfPeNPt4CSriUnpCwGUJnuGZAd5xPe5/rFLQSVRV7
pAr6fkPC3Q5pJAsYC+/yFzhjU0onbgrX4KP1vPKZWp74RcE0Pa9jlGi/tvcKp0nO
b3oahACWtB/FR2BgwxNS2m12C2AT0yL2e2J1j4uaV7fVuABs9FJN86bZ2cyEsQ8h
92TYqHOGKUWePtGCYxybNoVTPvMV02nig9bzEyHLAKHtOOKn/ZIzz6D+Gnv134hj
XdbXaO80X3XccOxYz7HDX3EaKPTZOOzJ37RPEa8AqqnYfETvVE0SkJdPGG/ShPfS
Q30PFoVIlmNhfJSfVTYhLBJIT5wZyoIWWukdIkzaFzAtBuDSi8GN+Wl51HJI4eXF
D+/e+vB0Lx37yL3DAWv1G8ZAsb9Q704fhJaFIr4hSLrww/CbIPRIemvmBWp/xNk9
GkFY+hVHzGou/7Sw2JvEciAdb1hxzFTV3EAkIlcgc79YDWTz+8i/U2hKczBLJLA+
wTxSCis0h/G+SjhMVsYuSYg4zaVYh7wPvOBswze2omqTTJOROOegx7PayUAiGbTt
JF24oFJEL4vXdD+D72DK3L9siJhx54QLC25mq9/OMlk1qLsZtWSb6zrWI9bIRVgq
LOygOJf0Mv2UyJW4b2ZJT+wWje8QVIf4udWorLPh/zm/ksFG3XhtNk85lVcUe0In
UeTX0RbBsMN6wl/QboWOn2tZMbDf2TTaPMKhPVPT5eIFCSm5XnuRLSH15mM/8n4D
AJbFQHMV5duWmZk3bKnH26u5YPjMTlYTL4o7RWcKVYToHkGlTcYe3hn5Pz9Dst+E
aixF8NTdc9MPitlh2hLklKRIO44f8OfrzaKLkFL1d1rgRzsjVpIjUwukZZwvIt6N
TqwerqTHZSFVsSE7ZjGmnAdLcjAPMhCZlbX9oPVpKRN8Opeo4rnXFbSJpEeGf3iU
qq9xCK8dZhM7abjNUWgb/6+LjaVFEJI4Y/jY+Ki4IHphtPVYtdLVeqFa/SUVvihw
V4MZwECrzyw34i4H24P9/zSLqeppeYxy9dH1OvCH6WunDtT1eFOBRynSeA4BEQYN
0A8rfaP/B4GW4aKvSn3FjwJcc5gB6ulILcRNy2KpogawKiRCysQXHtUcDF9TqaqW
BalFDIMsYxEQPCH+TLWQQWsPMJJGm9hbATZFCg0168caFzhp6WU0DV7yIJRsEbTS
q8Nss+B+QP24bG5mYAXRUeXIUpPqUSX15OZWee/KsVqyN/WrjegqU/lOHFyKOfh5
rcidqF9PwBajgxFXljRQf7v945EsUAlt8kkbxzVBWb6prFpiy9WSRfiBMtzxm6Vw
mxdYPGwrEw3PZnIR2+RzRGbPMoj/qxS1gX7q1s7pJ6OuF+pO+moXRcHY8iaJRf3d
8cbep6RMjwnbyXEpZ7ApiLLHtbZ5nBA7YcgZEjLSgMcjq8zblsyhnWyJmggG2drp
tVVNcLBSxPpTwwYVOj5U2q/D3c6I+8N6ZeRKXweQ/Ht25Gnz9NCV43/G4pr7it0O
St6CorbT2OfcJ0TevRcxIMGYGmkSx3JxyY+O7shVrL8ahJGSB5PHQeI5nMlYxFOE
NTpOEp5PHDdWQIL6/9viBPaofVCxts3Tpi/mVS4CFtP9WIzFIomv2aaOWWrqh6Pj
aCpEEe7Tc9r/r8VdjuKofaEEBTqG+MFH4apqYuFy0QJpTU2cjGs/mOeqh5XNtL1i
NkkZURIWApL4xXY43/Vdm6Yhp1cRYGrsRQajHedB4abG2PtaSQyQS/awIpR1id0l
dWDYbPHEl0PAfQ+SDPkgSg3CM81gDj8L0xpybVbjQRN0rAYw39af4HB2rcJXWDv+
N7/280/WEnnZlbX1dJ4W46KrO4Sph2VPlY7eZGmaUO9BvAqWL+5D/9twCDDyk0n4
iw4W3xH90h94eLMajcgZZjgnuw7OkV6Q4XWUtQ2mhDJs8CztWa9S94sdDwofvbrP
R/CmcLjk5vwnEvE15ogvcNJj90HRf75OE3DZEnW49J6HTSrV+wl1Ab/UU3WW/Xau
tOqGR4Ku6qj790se7RdkeqzoK2Stzb4VT+uAvzxszNBjLFJikYiycC10zt3GilVT
kNkgr7jiD3naFp+ELk3bNIQj4y9Yj02u0hB2I+Lmi9voCcc1DIkkqOkRaBVSeMRp
Pl56fqArZWzlzcg3Yc/EIsNtE4OTLJBgLWeStHZaiHSoHM7irbXSL4QWlxIIaynz
9/FzZzphb4M+1B1Wlx2eOO0WXM28Io1G+51XG6vvcE4n4JgCLArgVpmT80upHhyR
lUdt8eNj/MqYlWgZQU+itK5BbOKQhSRfbQK4iu4IsnNvt22WPKt2ZIPreqms1yHr
wGUs2oP8su6T3S69QAQSXwB0UTDGVDo5Oywd13oHHbYL1SlSndQHtnB6jlXRKc4x
10lreIqsWvikpEbZnSFGi9PloJPe/now9zIPxZZGqu1odx2G4y1hp6I91ejxllP4
vTpo2m8I3gv5bK2vgek+TJKqlPn3E6+H6l0tN0IHXYiR3mOqAmC8/VKOr7HZ0CFc
e6WddQdZlH0nSmW0AkgR2RNQ+wqI9M88gHrMlSaowkTVruvMoLHpYcbOWf6d4Q/i
0aOIr00l1elN2ew9tu7dM6yw1nglZXt1IOVEpeZPI6bfMMgmPAt1PsltCsj9Biyh
34u9N0pT2wZy7jzsA1bDrYxJxKYL3c9KQJmxL9cj0fWOrLNI5W3A3vv9ozoxmkPW
B46DybpokXk0uKEMmQIUw+SeivO4F4AUi5s9EbRdTIuA4LAM+IlCe6OecE9gFYiL
UUIrDr89wNbJ6TBkjRAVDZmZPhwDUrKijzDwyRhg1+IpkNaQ00KX5axrzE1XFpEb
3IusJKSpYfUj7vmxamUqSIYO8JZb1+DWjJ7P2Awjt8wOfh7MkCx90dwhtzphCbVu
xx2CGDnCv0gCuPgGZmIQgPGDQsjHYBt/2Rgosxts90J4CWrOO+0Dcvrym2Xs6vxR
4GB6rnAsXyRnjGOcdJuI8RH2lW7vp54ixJ/yR7rJ6OjEM5cx8bUYl7sOLjXhIjHg
U5K++Ij6ZZh56SKnyYEeEeHVlvTqkNsYhMqNe0wjrzY78exHSXxZQKQng1B+blb7
l6viToMRaXqBResLz35XvGOmQunhPny/RxNC3ulCvkU4/fhcfx3DYp1ZFDCtJ81d
PbxRviKBRARdPgL/fNNFfzZbAbVPkzG7SqrBql4GM3BkMhBG/APyrD4ji3Yxi+TR
jZQLJMAh4fL7YPQc+eO1yYbsk3qcuzM/l7sC+kqVMxkqGNTYgJFG9sHvbpGbsG4Q
tlLfQuOIgzMbrqZHcILJRTRISliieL0A48do5vG2JR6Leh/qI+DN0hxtQaYRrNrm
1sMUbNkWF6R08xlwDJW/3b98QWV5scAWAY8amFkP1kUV3OdgCk2dtRLi1M79huM1
5TAbxjDyHZxTsyHTS6PLUBCTwzOLK8JmbYu5Nis1GZhm7FTEFtHO2yonbNBsMtFQ
XcX9B0K828KP8QwQEBovL6hJKQdpAEFcgGvnb5XTEh5ZTS7uaQEE8QR8lexohCt2
ZTwR+H4/sa59HmsuARbPFy9WO6cgx8eDpFiARSJHng57pkcEBdu/dSZbGuAMhz3o
sFosRMcYB0hAvLIz0tg+v0YteP+evQrh4orloscJVbdmQPcpTAwejfVkBUp7C1rN
qoTJ0MBbzOim/vAFHSXnb3f6LD8ixloLHe1OuvSj2tqfrdpgVmQStwTPcT5QupSC
zrRdd7Sa6DUNHC9KnhDBqHxuIG13jPnpgCNSHLirUuBAKCSI4cGxpykbShzCEGx5
2srDdzOfeFciIZXseRp+po4XmFNpOT96C9NbYKGSFJFwKGAT0JT4+hItzr4VVkFY
mY64IUFUpcxpgLgzmSpB+WjN5VUmtVNGmgImR1zIjl4zCK373Qi5gatvwQoK+r5h
V3BHirl+adgOH997p/hpDs0QGhJIOMDSV//x0zLz2u2n9oh/VWb/7vDDV8J3y3EC
2iWKH0w9lRBNOvyCHKS98SCPp0VUqOQlwog3zPw+lSl2Cpi25dRqgCHW9J7I2O5M
uQe62BtObaEr5b0xYOMIohUILIE2GbpItmlvMrS+8M8jfUXlC5KFDrykWOLgAv4h
CxKRDUOZpKDwnqu4yIY3Py3qUPMRsoyiG6mGorPPRvS5x5XDHuWLxOit4t1S2OYO
Xvfutzu4/hsW/801uJZj2c05CXtRASao5tmk8dy0pwGJbIt29G5TAHog+pUerzXV
qH4jD5HzKp5yCEaGbAGyi/L62gK2o1njcBKib9iaYfrf6dHOACT1NAyAQ9YNCY8w
pI9xyX3P2EuloEcEilahdXALvr8Hd+kZg5M5soJ04DMmjHe2d+opEawcXQ4Z2+Sb
wNLjwjrI/OVrwb1qwthqsE9fJXjc5TfUg8qZ14ycg44ZMfoRHr4X6F6Q7YRhUBgR
pUL7XScdj5zb9Gs1RXph6brpy4G3SWpuckxDrdvQlR80B0/U9n0zjmEMa2Yeguej
zF9S/jz+HFSpZHFz4vnOMQl4hff+6pNeo41b8RkQ+MCLNZBX1Hb8+UJ4vh2TSjyZ
SMaPxboMQPaaaa8ySnBkV1p15Oulbq0FllTGfLjhzIAU0RHiIbbln2llMNBexrDm
q6fUlHwnPZEhLwgey5j9E/wotaAXeq/IspLF/7Co/7xAC3uBIwZ5QQjwqB6GvLcC
T1IvuN2w+wahrj+XkbYbm5cS9IZ7rcCZFiTMnLNBcYoBt7SosPgcToR0hRAz03Am
Xk8Zpo7KwzVLCSmpLcmucmvbeXBU5da3kdBrKPZzSPVx+99P9FXq0JIw8AKOB5qJ
6kJWOVA+TCbveVhFXSxNj0z//YCn3Jo8X+0GZVHlP5YFVqZSA3vOReXfyKwuN++U
3fx8Yp3DWuMWFs7XvMxwKieJSK+Kjqs8QycaHjIZN19NkUQJGRj+toTTdYRYrQo/
aNHBjKSvao8fbv4RyVGwVRTClD9mSQcifsNkC29gSA+CI9xjB0HRtAW9eZCx16uH
QFPh9+iSGfY7HLteBgQGz44B2TeTtFYb/iVfiaXTyZD4Ny+cx4rxFPZuF66PgX4Y
rWHJxraVuK8lnkfzxZC6+QhQSq1cCXwKt2i8BN3sJKCLQSgHTs3Vp0JP+bC0turw
lt3U/4fZdmP0S4xC433+In5XdpCJNIxnJDfMH/hof1kApQ/FLu7ohqlcTfh5t39Q
OtAS5K0L2qDk75YS6f7L9DerVkPDB+VB/vP4BnPjPLf/5fTYGoTdFhj+dPuypLph
htt8A8oV7MOUlBF48KCMGslXCiBDckZa6asAypbM0xYaGajBtp/48YT7hkVG84ue
AczzwBrKItnlCm5UoMEeapQfVIl+jHo2fwOFewosJDfSW87DgqvGb7rnigVy3FxC
hNslDxltoqp5V3Sa3l9m93AE34h72SMBiCO8HdAFMf53DI06bs+Iy14vFaArLAYN
HJzgu3lNyBmbGWNvz0V6gLH70QjV1PUQr6QxvYHfp7RsfrXhj7nw2bm1yUyKkl1u
cmgt49WvmG4Hhj/MM9/H6nR6lMxNEDQlr/TKLZip3QRR5ZfjsynBRhrsMQsKgwrG
b2nAlvedZmGVS21YgRRe49XOvcyfKY+NS4i0AglwTcSHO6BcdBXqzbr4gRPhz4xA
p2ugRKPy+GWcH27iQX+C6HgqQqYvzx8bo14IhdGOtf+1DDWFoRk4K72P/TbyjJEl
WIuPZxpPSoJrCCRu5xwdReXYZvrAYMJx87Pzby8w9O37IV1MbRBO8YkTtw1hh7Y3
Ry5oksvOmOUuGsOgrBqm/zeizrTXOHEw9KOyeTQ9u00o5XXLjeCfLqaC5Yeqr9OY
ZO2GkYAqdnzRvCfYccdg2EmFNgcO8bWEmfAt2On5fEcTtlLbfY9r9Ppab2JMRGPF
GmtrsvMmumb68+fiaxSn3gZ6y29p4YY7uTdzc5PEvLEniK7sjk/8nCRTFwFaKqnB
QB92gRmOyvWtx9h9WJFwV7ZO9JgzZEkImaSLjQHfIQDEtkdNh1tj0BuJGAHLUk2h
YseqJaYRVjK3/CEkzj6ciDu5bzfi8Hz5/aO7uZxHd2IMjtLwEkMfXEWQ/JGVr7vx
dPCAz3/a/Zeb2eyuy3OBzh+/E2JBGtzYGI+kpuvweuK+sw48d7jyOQS1zSqboujb
2LQARfOi8jqhDfC62c3UgP8kwlTnfViSQxHTG+4hxfhIFLTnf76L5ktf32+KbKlb
q86DENaJMTDeUNw0g+HRnxiAzH1/Cg04KekmdAhGEcXGSoIGTraubUH/gvMR5dWW
hjts8s4pm5tjZFiS0o7GsmTNdNvxUAx6Imyx0CVjGBEwsN7FDpj6ezY2+yKKW/D7
MdSoBMzMs9Syn/yAif3nbzsxXiF+Ga9yWB5aezHmgfKbRvfTN4OL2ugxVANqasHJ
F2zno7U4TRllAfdhJ22GmgrZb4pz/TG+Y1BLdQ4hODYjGIY+rK+PhqjOReQDQTC/
wyXb+aDgZaOPyJfuwexhxOuHrKOClqShkqloL7lXYVWNr3JyiuczoYMdgsAKwGTj
hl0GeVGWD6SnVhuk0Beo/MxINpZPRQmDrhCFiViB7djniLtIg5MgqhAKY0arK41P
w6AgbTrhLiJ8+WtAmeq1csOOngmDQ7TA3cS517askUwYBB0Sp2L3kcNsjeZ2NVaM
Y2ExHXEHrmISMh2OLJyp4/t3nN47edxW+K3HbmDICx5yntyNEHCdww7ELcEPEEg9
H3bGHdv2iiDTfiQ16aWnQyDvHOR1KK3i+sk4xSm0zCOpndYg8JfCvUhM7lRm0wIM
Yu1R1bo0SP6z10hSZmUKHBaYzz1mtcfrIAF/uTHgfFbsfXRQInR4zf9n5uuSU5Hl
QUovdjxghrsJfOVY1Q59As/3neiuPzTfYSAz/fFEgo0MGyHY/9V4ncx9utvWvrcj
J6x6iMoLqSg/vMpMcJuMyBZ0djPB8f8eud/v45yQOXX+4q8ow0ifiqWjooCHp2O2
8uzYNKi5SVJgYxMsZ1JEjhYczRcIJhEGSZen6vJxLvy2ORH39Bbp/MEm/PxIFaZK
hTb3k+P+3sKMKHZ9scUJo9Ch5lKRqNtl+8cDw5znKRevw9GO3zuST7jhj0P586wF
6rPh9alsQw+iO4+nNYmw7Y6g/vJkfDpygX4KGjWkbADPop2NOPA0QsSrXrHTeDRx
fQhPe5Iagvf8DkhlW7Qun6YH2bs+eJbWq4EgHOeXaeOsr9ti+1ksHXSJZ145HtZ1
gy8gJYWmZCUFMhLP0gl8N3pL3P+UbNHJ/fm1q+HsfJIY61IMoNx/PeO2o8j1wROd
n8xt4iP2y1c7pgDr2RJx4mvveZjrZGK6IXMCoBlYzhmxAtuXsy0kjUcwdrZGKDMn
3oVBDXvOv2v7GDQZf2aCXzGuLvCI49cgShBS1PIlSphRN2SnrXigMA03GIygmKHa
dCm62eYgAdYB7FivrVyh3s5h2M/nlEUd4eK9yu5DinX50tzY6kgk+ME2VIJeMAcD
QbG5sa7Rcvsf74U4iLi9MPmn8ITa1kQdvfisy0m8ryhXESOYlIGFq9JjaZPcE4iQ
D3Ybqv1CIsLJokkhGnKGSkOmlff3MnG5w/nqgQaY3qxZNCJjDhok1AzNyCz8OlY6
IJu1dcIMiQ3TwmBlqfRW4+RvIxJz/Q6MxS+mWdHNOGlQb36otE0r9P6W8MvEurmr
Tr0JVVsQv2k7WAB6YqLZlIdYJhjCZ2EcAwzUT7HIewkHQZoFKEewxpE4J4P/8uRz
DTZOivWPdCv081e0gGZ7eqH0Oyfx2IgNN0bnO1UexSi5Qif99mSPs3yYE6ifVt9N
Cdg8RooXd7guc1MftdtN1vnlAC8aWKMNN52B5bEb6pC3qgaoQmbnqL/i2mMLIM2J
LiImff98kw+Kq7uut0KAVYWoV89E18hKglkpF2upZTZPbkPLV7K9/5TuwhZKdNKP
5Q9pEfkpUqHs/5FdGTqs4uIFk9alMDKecgQ9Pi2uFmsTX/NyZnDHSZ0I858ivfFz
TYD6HklV3Ws/p6Qd67g+t9YeREWYNyzYLEord913ktAfQRl+uSLNnKw4t0u2xwbY
rkUoPvsH2vM1RwGBr9qN4zDIwlXCMQUM9gNOUuAN2jmDQEWzCPOjsTLm0qc8URSa
I0vepFjBFD9Y2ZEQccjd/ih+hZg0dnTC2z8s9YFeTLtZDcTv5T7rtojoiw272H+C
I1RtPXy2Y/4Ck/WUOOvnyUAsI1ygrMtjHlnS+9dRHofChyUTHYMSkqYgEi6gMj3n
jk6Xw36BcQrwSrvoYXUcFwvwQExbXCFogiYPChA7nEQe1fGzVj+UKyjG8g1faMi8
RG7r5h9uj/hQmJhEOWyuHj7yb7R8tPhSWKpFSP18ZWyeSojqar8PHBexW1ILCOuN
4WhQJsiBQaLKBOn5c5lD8pYCsOiV2zlvMIoDHyWrLGHMvy5aPl+syUSwbAyPq3+C
9raSrXzX8kmYvRXuModwEgVDYTJNZDx9w8idWJSlL/I7fsNToHqATIPjVyCylWj4
sssGIgqinkxm2fDVOvpqxw8rWruGYykBlHKYLpS2rEP8LNqamdtEMWaq2gsh73Tb
59XwQw0XdMFnuhGPiUoDkcHWFsiQEl5VFJ9w4Mb681LfzaoQyNuq0JDx8hY8dl8A
PB55mkswWUYXH2RZcMhBWHTETLmgSPT5J5V5uZE+a+6W5GT5hTDBB9N0fLfNrkLJ
MQWoIn3h61etIXgSFKHjkabG5Qs6YaegqgI2PPmH/aBJhtJ1ZK1eOOuXp3J1nztw
eOH4QGwpO1IWkf0SGFXcyDbxoeT7g9r3HZ5toucbMp7Hcxr55itPWPJG229eRDTb
K8NsX3Hv0ZuKpZm48R3uiqqf0zZSuzb2BiT7gmwJj3ZB++bA0piE7dC8rjKadzvn
SDmR9yvmn3zYjzRykH9dElEyPTIFgSimqTNTQufSCOVsGyU7K4YYgT5AHYYOOhD3
GMOGr7tKQ2O3nTU036K04ui73B10ixJBPaCFeVxEto75yr4Y439KcNeoat41W56E
Fil/2Y6A+ZdyB3lAw9SpZ/ZzvthEY2p9zNq2i1dGXYAKOIrgcesllf+XbqzW4nsX
enOFZYozscMHLehI9suSJHVVkwbcxMW4N9FkHmLzUu71yN8lswaQcBk7cDh19EuX
o9RMGo52fJPGzEMG2Ia0LuUDNZPddgXKm+FmIejIEJjfho0zbLW9BNaf/Wdy3fdF
X4EkEq4WoXzHFLubXqekoO4weN6K+uz/8YhmLcXr8rbcOy/bOy60kj/y6wjNuImS
4aAseK38zyyRp8C9jFNXwGmKVQ2hrc/SVuMvpOaYflyzjRSIiIUgKzPXunZGhKe0
Ro7/RsD2oKPRKQuDUFdwQA7QzNVARgNwVSAOr+uq4PvvhSgPCeoURylYNha31kkI
S4zoWUSGBbd97mrkDDKVO36HhX+knR93nMPq6SUguZtbJt6GWoeQl4jGugx7XmQS
oZsJ7bOqUn7PgoJgG8OF08aaPA/aEnayX5Y1w34vhjVceyfLW6uiVMv4sKtaaZsA
jpUk9DbkE2l4e8pMc2uH3OnUPS3lXGCTjxMbGERWlkp6SdGAVIZkqFft69b/nLCY
B3bc6eEN+ppy2Gdr9eUH8jlyKjuXDoYmakoYf9EOadXeKD4cws/WVrtHvYZuyyQB
fhX5PQ5ynUHUdsKh/rdtb4vECWlhqh3bhuT8VP1bC2NFtegG33F2a+0sbye1PTUU
LkXUdUaD7NrdhdSOMG2nrrMYJ8YJsuPkmp/u34pTjC1QCVWOvyYDOf/MbAljSX4Q
l62fGdrezJb2po+dxekTx+TgLmnFQpmHCM3ShxjnPgZ1sdQQ3qFa+kihUgLVvgml
xnxF1GC0MRJH6uN56RaJ+jcx5D6uaetRBYc1emQ4T3Mr+/a02YmnUFzpGocXeml8
ZRDyXJSoX9W/7Gt7xXFBt6B9klv/dQ1AO+/zLpMazi94EyqZxn/RyHMN2VEKOb1O
NmhklKOzkfcwETsUWGAeVQ5ukTqhsf/3dTgmtH/HNU3/NEHndt+syaPytxY3A8pC
1gpizh0gNTu70t1dMEAtI7811Y8IEcAuIfp4ELA1ApmDr6AuAa3Dvsrqw5TjlK4J
UR5fomHq2wE+ibwUfxVhvtFdEujutHTgdFuNABbVOmkdQT6onLRHn4R8T4kIOSdd
xTC7gh/9VcoBI+EQAz3jfD9YxHDdpkqRYG/Fhow0fo1pB+n2fJVs+umWmL3uuef5
PXsfkKEhvfvuGhr+5qTNl7+HskQ2ITO/6gDEUYK9Zi3RnkZi1jT2h/BNMcooXljJ
SeeQPku23minE1C6SFxYLEN2Zt/skoK7q//OU4gnlizAGD8mhJGqK/abmz5nHvLL
C5rtFKkEtjBaEM7gyfa37pr0uvxOp0RHFwWyFz/KAG2qTHtRjLVF536IJ4DdI8gJ
E3nK24joZ0Twy3jE8ZU9jpMsvWVEsOMy93dAOB8ONeuk3o8XcWgAsQE2ITpup+tz
fmDgl/ElQyvNuKE5s7phTnM5GR6n4oy0LNETW5nAvb6OTaNQvuV9wUQuLHS9vc4e
Qx/t+w4tAHYbIVEtiRBC3oD+JRR2LpLQlBK+Lkg7U7UMT2PthT3ZY5TWeStOw/KM
NfTGY1STuty5d/LxMiINvKBFeBgn4bWj7k/8yJW7t/9Yrw61TcQUOQIZby3ZxKTd
yJ0oWHv36CtRs469v84yk1hzvQCv5GTmx5Da7ZVyyCQHWJJb5wQ2ezKoHrcxbPJt
c4W0VkNjSWD2EjOJ18wBD7/dpPFzxw0qC+VsfQ5VDv+b+zKtVSmIlfiUQMMkd/dD
YBVkUd6FfhFZlteY2T4U28PO1mxgjaElYQSnb0rwHognqyqm6ElsPq9opVNVes1d
MIXO+MwJr3CyZi/dz9ApfzaV2mZzaxvd7+liIYGHMvfXXRDVXclVULALW/OmpnKo
szvlK6hn80VwoHqYABkqcf+JqdHEBLhtkAdohj5xky5oVHKCMfR/Tqo1HZ1fM/WR
dFBrfgZfvQ/1MTMtPMOrx/uIr3ZIEWAmOY413ZIPyxZ0zPGDS2zbgsN9TW0sGS3c
eY07Ap7Q1FSJwMGAqe3pIDR/gcNm+Gk7+fTIq54NXTLnub5BBf/Rpl+h5QXbv+Fk
q3VP9e1wle7vJ1Un6AoaoqJAX2WuAI8YYUyrrDmdPcSBhQIe38/gx+1k84NjH20M
EmqZ+2W4lLJW/p2+OOsbHjKLF0XJE57vwKZ6uGrjzAwr69VHT4Vgx46B15svF4Ex
0CojK/C67efG8ndbC6WDfdldza8jSPjrGf0MuSy6RUfTwzF8m1o5f6RODMM1+HaH
6ukx/DpFxeTkAlB9jOfH0rX0jpsipkKUlV0OBss6HehJj84ydMFZmBNh88NOFnMF
heeesHDzcscljynowUMljoerDwVigGZDJ6ZXzZ6F5xS1DCPIipZSoxzFH7Dth+XO
OYEXs+fr+UqNNLf2GbjgamHMWN2Fl5wLVayOGgG2ftlwN/OHq3ZAI2TVAi1LSX0y
Q3iFRfpjFzhD/O8htOPU2r8k7AKsEfn4b62Sz4ouoLCJV9KLsQDNgrPT9yNuO0jN
YA3974WekWyy4IyDpxcN6Ku3NOxJwL32r6xIliZXTCFajRUISdqhVD+wvr53t3KA
O8rNlr+9Xs9QZowhuBUA3oraHT+V2QUr8mlwMA/iLhMwzkseMmQGgXJsy89dBpgh
Smn7ZQuD6FrNW9kwPEuiIv36GXkAKuQL/3kEon4Qgvc7y2tbOwT9fElphp6iIDbA
rX/CWKU2pQL1MQ7ZDvdmgc/yXWZjgt9zXbEb7C7AYbCAJyX4T5cZTquAj8rqaB9e
5IEWaNMriVR6wBWhVcGHg+ORFfZ8CpctzJVFRD50ZRavYX3QVekIi2IMDR6OLTPp
gkKTzpExgRVRZ8VWEO6vMvS2O97GpOt3l21YRnWA4SqxpjCys1Xs1pLlr/lNf0I/
IfeAZsfi0a8VijrZnmTY2uPm7/fgDu+/mDwQ/TSdduTOCWFVaWZgrP02Cwe6hbgA
zLCx885dQI8cihOddNt95//Xef2Z4EyTYEZdKHLKkYUAxKgJ3f7oxUIw+BGz3K9D
dCCvDiEQEafmOy20ByTm3vZEE7I7o2erjrkbCIeydrQdFSpBdKWW15RNllNiNpqR
TzciA18sKSJHQG2i1SklYVy0VASroFP1JBUQkPkhMIiKO2f7GrBdNeYL6vXRbnSY
XQ1ZyPfxmEc/sOpvWcMpjBZCq+RgOYhdeq31k913czmGDm236nMrtWFsL1V03CEl
CP/ZZzMwsD0lhbe1OyWFBRqtgnZlL5fJ+X64ilqImlZgCoK6eTs3ryUibHMy9U2B
HkxlsVvUh/iNEZVYjBOPrc8Ye99gnT7+RfkZR4tbLSA4/7IGGRalPjWhHQc/P5sv
x6h98lEG0mmZtIZLPdHQY+M6FXIMm8hcPoXEPer+r1X7zhG2anOLxw2iiFyLqXIJ
VVspz1SbU+vJWymY4DH2COWjAKtvudFABqFE/1NrVpPqOTWptDz+1ogb0itJ+waq
tqsVZV4SgJQVgCRKAyBHTjNxFRQxCciuGtoI2CHB8BhpvC+hIUZdNWuzblgwL1w4
705uX6YAWR/gJXLFcyT4KKtiwAyFuWSiraXtMjGUh3Su6ua0zHNCW3sVCRxDx7A5
7XbVsp1jhpPtg4a5Yaqz9iLahTMn5ypES17PUKH6XPTj4mg/lx+5KL9DeRIHfwEP
yxsdVoOnmvYhS8q7W7nQQyeg/IrbrhNc8LKb60M37kGL/Hijreq+yAWpAUOVAoJA
kqAvg9NH91p2kqcUkvOapKr2NGqiRgtrZ8In9SN09+b/HoVAtHFQJA9ZUUyYBlPL
JaKv51MbgBRyZ51Dwt96f4+w+VD6dhKGy5RgMJPkw7AGRuFh5mySiYtJYodiEINS
+Q+u/CRPQYUTrMx3W8proTn2Sm6fsQRXqSwNK33NVlVf/aUdwCtWCXUKov/dkJkp
cCZP7PPNdpvgAewBBFoJuLp3yKZA7L7jsWVcAb0jYsw7UbKL+IkRvRzzIIs+4McG
cOgHI8ESDIwBQ8qIOvWrPzlexT7dhyxAvV7NJyoxzIgxT45R2BEH6Oa7JJ3NE4/B
jlKNTLcmBN6cfa9tT0qyaRCIUNj1T7iDrLWxPbWMqdoG6aWQwChZHKcbPbvPKN50
4T4rV1Q8UUkWq/26iJ/AdNBgL9PxsYlw5xNlEwnILsLzHOSuiu03SWKiBzfUbxNF
WALHg4e8feFm5fuY1+yKbjVDKzpW8HPHxxCrc9Fj8rzX2itw1TjuWuOdW3i6lvce
x5++8whfeuPd8QUfrUecBP8E5UQwXySSN7WIuwErR8X4f+bqIn4pQGG7voYK0Hqr
/lc9OqKMMkt0byIJvBfw+52ONr9Wmwv4ViBVV+ypLq4I8H9rjTOjL2OLJqoZVf6k
cMHuKlQh/6aHVMQv9+zHawQOiKUqW5s0uRFsvOAprTxjys0jbxtFyfpRSHaITTa2
x+1FZOFBcskvtx1G3L8/o+VzgiMn0D9JIz7x6jU7ytKl5Y5qnhB5dc3OO6Wc6+Rh
+j3UJ3A0Jjd1n1qsIDIm5YHJAF/PoblVKZ3Z5XtIS25r8/mqsVxYYpz2mPQnm8QS
Iux5GmMF7S3pqtcgzfmx2E7XeJZWDNdcM6XdxrUfKrHu9c0xCRKeWtG7ruDoh40k
oW9MKBydSh1Tv8wnjPvZo+I+iYxDkKkasBSI3aVMgby9igfAi37M4Tc6DlGlsU8z
Ha5OfBuIdPvMxU4KhB8yWwvQYlQneP5TweK0c40aPPwIuc4EnOMlSVld0qmuWu/2
4JSo6px7MCUAWFyj2CVjgcmuSZIaaU/wlqMSdyeV1nXgY2s81rHOHDCaIUUN6BvA
N/9AqH794Q3nz8OKgucW15sb0u54X+d/XyodtInuMz9Pbl0Skkvb2GomKJKm4bWn
f1BncukV5T2Dt83eKcoFHsvvGiM+U0k43tQCT+MVOdMKG8c6KiShWV1tVmCsKrQx
KwflPIqCIO+2BDlztTzC28VdiwGrrJIVg8U6F5BzSHxMRy1sGZWOgXE17YLYI8Kd
Gc3HHmweEABN+jvJtcvOQqMTpVYS6x4OkFrqjXUC1R8Jo+xBs3igBS4bDCRMUukb
QcdUSuIMKb/6S5B4hpipQPUgWHhL/1JCASToZjdmNTgN5yMWac1FGmwhrVd7qakA
b3stpuGF1DdAC1Rh8/LVDI5/LPEDueY3TwEx/rxkdJmOrfGCodJQjepvIgNtmu5Z
21Np9U4US0NrlNuAIF6OchRGH7+Gh2C97nSNuQEgKruu67sS6W2c3tImIfALUjn8
AGb/oHNsUGXuejMWN9isfkbONcH9tonbE3ce/0Nqfo+RKdekEuXywDhY3ycfyDIr
ma0J2PYtnOSDp3FC0Ux1Rg/kX60JI2qvCI0JvPqJ1oHiASd7mTN5O0VXe5EVhfPG
QPhdrucg10eN6dHQMQq9IMEe6HvM3U/mRjVjSA3aE0rWYslMJcjIeR5vaEl75Hmb
QjSUGquAWgzDcnLfZs/Zng8u5D4nxdAk551/jrXbGuhfh5joInqiuGTuaAXz7Dxw
sAWvxre38FZcoO0YBz6o3pBV1/HmMyVHsGv8YkaryC5DRJC5flz33CIfBb6HQbxl
Hjkts8oYgCW/NjHS2kB2FPpqacKbwILVZgZDWyAUUqXEb3lKm2x8HCFJXxOrPz3d
Ob03/xMc8nyZN/3FuMURnnyCzpLMEDhr+lFe4M9fmfcC0zJmGqS0UWfl8fS8WCq6
9u9SmXuIKOhs6xeULeYM/MB8YIA5/ZIO/QykVaHtitF9D5lZnM8fa8IwhohhAtQD
BHz+3eZFwKg9J3wMyT1Dt2u7CtFuwdv+PQqKeYisHWTmmth1LxlZ26VtiXUnVMKv
fDG3Q0Qs1Po1P3fSBcK+TP74oRpVrBPxQbEGl5Wrr5uiz49xr0vFEgpR2o2wO/1+
YCdRqNK90JgJf7NKWXAHtK+3lK2XPjclYpBVhueMRNxYGYXVroycC+O4Co6D6Sq/
VxBqpu5U3QOsOYOtgdbM8reD3TJ6SVxT36OumHoWStVNDAiYw3BgLkrrDLKEfAOo
nVCC38mjV7mjiKwWxNB9mxP+ThUTe2MpuSYDehwqcq7rPggjb6toJ1f+CGaW0xkf
rrICpfVPDkBkSCzukqPtElfhqZQZhMEa+ieu4Zgb9tspNM7AtVEVy0wOKHz7a1er
DGIJxn/pVR3jAvdv194qwU/JW7TLqkqt52HbJysRpTiMK0NsvMyCmJ4YJNCFKqko
YpUV+RftImWvogSwnZWfdjeYOangUjovxVZ6qhZWqDpeNRnLElGzs3w3ivGg/vho
7Om47/3gAWOPYn5defognN7T95hY/nzmou1nRDgfjrAVjN/P1slE30TML/DwO2LS
GF4lzYJif26jGJClSNn7Ocz4akoLFGUMQ9oSNGoByYpziRsDeKjqXnFKU3AX/fL6
nK/vlRevtxCCuqBPQRs4r37tqB4TKMzJkTC4EG4g133i05Fbc0Jc0wBmciW4i4JQ
ka4yhSNDVPx2oA7VZm523LawZFdXE2hiIOp5frJDVj9hy/aJB6Rn+VWzUEV4/Mwb
LMgLYjV6kF9YMJsa23Qk5Q8G1zqJsqMOUMYU0RN1E5r5jvRHulSy8wKMeXi+GqBG
PWMsQ+iKXukTDjkIhiEPA4+miAmNM5lAAE44NmZyPRGYXSNIEza8ku6WhKg5NBTB
hgQ1NVVLO88d5O0tZmqWl+W2h4jOevg1Sskn6dQ/B4T7RGU2tqw9/I5e7H/JrOLq
l+rVCgJss2tb6bdo2NNanSgsw7Awpz1OxuhDWNuAyTG7PDOxeslWrqRor32nyQGq
Ze6tY+HA92q/g0KBNCGgdMlW/5zN5gWTtPJ4NMZtdpqHcnYieC6INkMBAYikIoUq
xD70lioP03/EGi/2rqwq9SCTDB6PgKdGX434Ejg7n8Xl4FRKpMCmJ3gayir6clbo
Fp/U50rSY5hi+vDu76bHHIhl0AOn5QCZxbWJSR6ekEqal/iRSMxnwb0Q8EI7XlQf
aJk8PdlZMIMOwWJQVwwadwxxC4JwbAclRvclsMEIS/y6WqtH+lFnsvcgkd6LWEbc
2QGN4A/q3gt1T+gRLcJDJrUixOvgcF4KT0l1NAyYwY+NSIVMMVcBz7KlGJk9HwJt
wYeeLb/W6upnR2ZqK4uo4psige3yo8fxi1EyegN4pYFJJ9tf38jaSm4EQyqSwHC1
KlEQKu6zJ3lC7qPIPtIntyaAwZNOc7goORXZowu650gUSXhaX11dexE39U8zFF73
VOQ5RdZ6BTEcxH98TGfPoeGD7g5ag+YStcWCvIInMYqoQHL+9D8u9BpuRfRs70q8
RYRnLAFfmtYT0+YEvP0vXsvL5O7D/8MhL/CpjDSdnuo0MxrpfQvTtP4zO8/zQEIt
nwn2vjMML/UK4FwPJsAEY0i/fsbraR7SuWmT/5dnwjsxPpglXBb68toFZo1TfJ7f
HxmE3bSEetzXUFqCGip9PHh44bubkzW8M2FrSHuat0u31/S7161KAEUgn0lXjLx7
KNl2UEfbQ/3jA8uOkjwFClry+l8iFAP2MwzKw56wi4jJuvB0Ef1Rujk0VBcfW6un
kiFj2jxOpnK1NwfG6woqgS82QKVpDGEfUl8clza84Ka1LqiixrwlfcB3vrENJD/0
3BCqQM0Zo1yj67KvXY7hykafGmwutw6UX/VsDk90/m4x19AbhoKqBVouD/XU5+Ry
UJZOcoau4yFMh5plBSZc83gr0B5+Y5URjhdA6RAEZ0TdJx8bDRzjJ9cTPhBZhXJ9
b44/A2cZTJap0AGfXHnFbcYn63OKviF0kcq/sZ66+XT+A27/0PY/jOndVgxjsdZ1
WKQ3kNRJl8tJo8ZdtuMj1TBVa601D7iC+m1DYpko2h59co7YELDmG31RLUf9xFfT
Shd26PlbORmJPuEy0C97Pvrlaee0tmYJv3oAsMjff/a00fnwU/HfxWlOETa+/gEP
mie9HAjrHrXxo8hWr9G0IJZNRFU6nBOQDLt4NXaWg79R9pL0wRvGvZQZAWxp6qeC
sXP9mivDzgxc1LpdoI3i4pm2kAX+PDKbD9rPRY5qgpu2qbcAHerJJkjOqc0braZf
5spXca8femxjNgZGERE+Ur3xm2WTKiSwIgvmvV/EuYAdW9QTpHyl1y72AMrLBolx
Nkuq/OsNnziPHZZMTQTFO/+7SxQzlwmgC0Ljn8o4+tAAGDxIiI5QizvCLac2t4RC
UIYZo0yBL4BrQ8UKR8V5vz7zGbs32LuouXMKKmCvhycZnOJ78u7DwT5G8g9NQief
8YuDE7Zts9OM9hVp9UZQpubNX8cJqOWQcnFKf6rLToH4kVTECczM2YnGoBnsosVz
+V6AHhO8AVDmxhjl6e0yp0EsI8d0QtN+3dOLBGbPJKJvSSAqrEHK1vzqMtWG/Bba
CC+QRGxBoIukhSjwKrWLq2yqIrTf0IRWnPJ75XkbzX/P1rotgA67zDktgjSZp4vu
zsCc3VBEtTnoEJPSJN5llyPkDz3UgnY4SPDaQ4ZVrudCDVZxRhab+VC6bk9N+w61
I+s1xfzBy9lx692FakqSi+F3SRf3vWDpPf+TVetzs8apBClzZYIQaue+m9cFtXTT
YiD7R5ss1bGXfsoSaTLFTDc9PbgxKfkPBtiSEaVyG1Y5O+SpM4zJngufdblZbSO0
cebapwY5tWb57U4vb5YC4A12ljrxjsjJA304dRTZpVVzJxHTvPPt1QBTnoxSpGdM
wyK1Jiq16jEUFyq14F139RXEyrjmWzRqNXgWmVpMfgOA2VLXoNdhTIVk9b37plNi
UsKWsrvkVnVconOuTuej+k+OgEIp4pDih0tcYZRIpe6lzYIA9C8uovjHt9bERo9m
hfIfKcLOH8XXqmBNaXWhUaehy/BNGyWMOmkuHStxXdKGYsFK9nVpTBc8J6D61C9g
tV59Cmme9Ff3C9Ki6UWSd3NSc+Ou1VNaFmfxP8yTTDxpAp5DObk53dPb7rbBiR3U
tINULEhFwJGq+YG0eDxjYFIaD2PFmmbvWOdFzlOMfcE3KkbC8a+nwWcpkV2zRg2Z
pBGZsWXEL1j7k0jkQXZr2XSr+BnEZnpjj7ChPVX/Zl+UHzwJroYudkYuGPeAZ1GK
aupAdrtbBsShLDx2c4FJQQyYapxS9QQYUveWuO5e1hWW4TXXJ5Q/DdYkTCbCbyjt
nGi9XdBjgR7UoSJ4XWwEGpOe3wjSUvhTVZWiCRxh6x3KIPTXJ216+3xy4iE+LSW3
yqjVr1cebd6VVzyXkn3R9LFVZ4dlFYPhXnk6N/+v3DTayuEVtEL14LWIt0QFVN4L
BLmDT5RkmxsmELKqefrIiQTzTQr4vzOEExQEqR/ACbTm47BQx+Jm92c68m+JwBUk
H8QF4vi2t7N0yVYNupkfMqR9c7YtuddDA30o9b8pSUsdXSYkJtdQPtgW80/+Gc34
i7giihxrE2nwVddbC6dZQ1xNEpe8oPEJ0zz7ATFA0dhPig5X5jk2EY9pZkq3L0vx
mv/JmPM+JAwexYiOVkqmIm69qu1Q56M7XDxUeGnEftzHTxcHZy7aLKX2DkO45NfJ
+aPwwldxBWbXBHhxSZXXkkmdMCogHoQOJoRUvYwDQ3bh81mCxVVNUzVchmB13j1F
sVEzGPT/61DoibJmuDO/OR3R6GGzg/Jh1YD0UUiNF7tplknHsqweWnhsvUoleS5j
Eu8vyfmV1DojROqOrkEf6PnheWcJD/XQPO9a7bvnOKjtflXQwRHuGVHdYy/uPlvV
SW3HVzh/p4j7SG++yfFo12h9dJpL5UIjoEjT3aYE6GWqRiX6kdGPHuYLvO20nZff
UNwoYAb8quB5S8I0pYJH3cAjvR9qfdwKPyRp+qpz9GK+aTD4hS+fVEFN09XDZa2B
SvsHzohD6FOgFy46Ps5w/jybVUyJTxsAvvN67AjSWrvRqcI9yAhwbbOQkDC6OXXP
ioL16m5/U8Tc/YkjCiClNHYPCrr7iZipqCB236RjRgUf7PpQDln7NkOzmjXhCuDn
g02T8+qIgVdprNZPf7a8tzIQxMmFq/hdFi6HhO/UPqWUArNkfR1NcOC8cCNOCc3N
PivVUX1Vyv0MIrvO2ZkY5hBXv1EQ75Zmq/nbATxSMHIIQCGeny67BmcGkVumY0zv
rruSzowbtpSQ5urW4ac3rutSQY0C+B56xm9iw0P9T4oQ5pePr6xBE3P+64Eqv/TG
b4cyDhXeyRcS0QQX5nfV3HrTOQg3kyy6iILSFXlEXOsNkPjct6CQYYr1ri5m3CyM
AaNbUqQrCGYeDEb3z4gRn8PiIXCTnjvtmi7Jeotqqu6FeHefT44UwLguki/IZg6h
ej4kLG7G/JzfdgiIB4plk/sXHJ4okuQqNtDwU01XjSxguEEvbaSMWszxH3/TE+re
lLmN0xCTD/Kb+aDis2xfuA4noZIK2KpM/ZbZMvPCgx58Ig+CCKQVU58B/rDT/OpQ
vD8S+31QXe7pVJUR/sZFZ141udlUeQu8JE50VUyJjlbVdLq4sW+0xoWYEJ13A5gD
62voztm1LVk2INQ7ih+iwpuCmFvSyiSgCySWg0OPEkv/NC4ksuIm317K4yfWH53t
7E6WgT2mswmw6uv2MA8FSIRxjqjpzUtjd1ekHS7E8z4EuyXONk1liLnBWzoOBevU
TFdNW3xmJC9+vvvkxd5aLsWoSo6m0vdTjRlHB3Y2zDV+nb99RlCaCwtgUgJdEH0O
GpoNoBNHWMkdqDcx1LxmpVhi11pWjP6A9JczmCfdAsD+j9LnUhItEuJeRMByUT4C
Rlf/D/eYKtsia3HMkqjwZBLx5IPZpDUwy6qs+1LhhGXeyPjF84n5Cp76828zDsG8
WdFOGXb4lU4zXKCy3WQ1gkHyDjI0wso7fRIPfzclQG9gX2BsJxoLiBjroUKOq0ju
wCnbo9IXg//4DWX7XKTiCEoITZHnv0bQumndxHh72hRhI2Au2obBuDcC8OnaLT0q
mQ6xyK1qi6ubrTmOT6f+M8UIUfWmCErKhLoFSprWoNcY9o9rsH84Yf0FTUTyhjtE
N8PRBXeN3zX1v3dpPa1LrNH6o83+tLQ0Estz7gspzZ7EVbobkBUQ2lbEMe4vX75B
MmF+JrDL81ByNCZAWi3qDy+6MknG5JqVqpFXV+vKLZFKiStjORYeDnp98SSTIAAx
4dSD0xoQy78eNEjyg4T1eAb3ysmcZqaiXjMZ1ofQ2Teb4XXZKGQdeA9fNcFn0Xmg
LFlSJL9LzO04ERV12MAYVC3rDGJmE1xNrqNFQoIj/S8WNS3SyYy1ljdp4z/3ZhOE
nWX0D92j1d3L5PTKOCENrWvlZGDxvXzbd9I8VhWG+H6XVE1nF5GMXMCOO5DGXIcv
2+YxZQbOqFleLmh2CmH7gzDoSaA2/zDmpJh/axwHWITDsk9UYGOG8fUBR3PtGA9U
6lrYoyiFV2APqELAYm0ZcnhBDT9sCqDVn9S45XzjVhFWKubUtQq7RRgCocVbNY1A
2o6G6yVYJAi4PMxnF9DAFGlLHqbzb6UXWNTE2KgT4MbwpVuTYG7vMbcatb3mCzSR
PRVQ6cdzRaOwjeJUpTWmn0FoP/sCEAhDI8wzw6qydB37ogOuXDPomyiRKCe4mTUD
Guoez7Cr4BMKlotbJQRNvppDsNhGUaliKCdFhmQ529QG+CWmPjjkuxsXe3T0D+RW
3u8hZCfxDCbvIN4i8BDW1MB0ioW0ZSTjuzO5fhtsWxqtvBqZ5jYoqkJQqsoaMm4D
yoPcY6ePJ4nsQFkj8e1kbRM/HiKxGjPOoSCoqCxXDGK4G9sggy4vDUFwIRlWelMN
GPHe/WjjBKw69RvF7loAcTzJXz+Gz5KOc8xb+HEzXUVbn4LnywzDsblY+0qjk8PA
Ch1agqSMUL3u282B5DsXmquxX/D+K4N+5QUtxJjB1v9nQIMV/NC/R3BvMHz8j9il
pWEV7QI574sxcLXmRloppkQb84DBTrD5LIcEMMIu8CULDlqUCOt+JDahZDx/DW7j
0+ycMm/pBzkunSyTe2LwXgKpZBA3AHz+pwGVYU/RWNEXko1F2a37Z5ab8jRodREE
49Fj49aPVVm4ZdeXA7Rse0lA3DUSnxVIxcRHAHCuy7uEXhXtI7q05Dnrijnu6dpH
qLl0oUwQKk2BCLJVvxm1BSuNi8SIeLa5OjTFF+o9KBMhE80TZJVfbwUFCRpMeElw
Cl+z7opsG/YkI+SRKX3hIdaDQjeQaOTRuXA3+PhzuuqGZ0nOA1NHrpfjtXDSQjR4
FERaFwaTf5t2plSLtEA0D5LgqUfchj6nbh+jenaio93P6Kz/gip7b8IuE8AlzjRo
Q6Nw7ngvrgLWdqAbc2175tmY6U3lAEXJuUptwivbq/Kr22KwfDeMdTJq+XxDoaXT
v1aFxXsQqbsHimiB8ZIQ5xhmSf4RqpXqusIYR7NwfnOlPzSMScMDfWDuSwdFAHh2
/H7SHq5gWmY+SZO/ss9tFaPOXG7q08jID5xPUxL+8ECoytUBn3GW4TOKlIes8vaO
e+IRY086Zt64WMpb/SuYTk3iHH7KBEwDaSNVLENpTtAdFT3/7lQUisncfgC7xKKj
E+YWfJfJ6w+KEpZUxZmK3FDlECDncSuezRGmlXXjqXKnB4+gP+F21PJYQ80ZgB54
P/6ZcwukazEQ8lLFjmC1NjvDR8KavGBeNPtqGxFWyaLzisgejcikPeV2KamOwlc7
pXZMEHbTBNHdzrXZAG1F7R5kI7my4Kfbp8LWxMMg+5Xxu8FTnGKedVVWe5M7AAIE
+seKYxtOaeMf5YR4WDJE4dKHdTLA04LNBNJDMm/0MvhcLHwAu85HSXDdHgDITRWA
yhz/BHwUorp0bCiDXzhia/9GxlSakzQy3/2voA7Nhpw+K6nhu3QuYacIRnqMxV95
QEyHrVqcvxwmeWNUFicO7KjQv6Cri8ws/ZC+ad4VOxemY8jKrZYeiHja5Oy16OpF
Qk8z9oPi0gvuGmXHiHQDJbj4cHWYrzTxSybUZ9FpFXIjj/9Kif6mXmu898RibCmx
vMJQySyz2O6W0pxZyenBCMjrIvYyLcR/2+egXwEe5hPrc095K8y27nfg5GI/a7Mj
rHXLs30NiFQ6J3TTSnA4l9bKquBMSIXn88RfOMje64ruo0iikZpa1FyKIcggHS6y
Pb73DueYdC0j2ns9E9Sd2ws3K5sOYPE+7mWO1ITdp5lOv1DRIo/0iOPbYToXLwEM
s3tBZRboyTSQyeYy1Q09+QyUOCoY8IqiB6AUOYgWRBQOJeGA3JgenzhFGzig4dqb
8UYWW7XXfZeZ6hoJiyTMtwtpR1sreZNWGy1aX2CGi2Vu0sycljWgBoE3I40shj3d
suU7kVPfelqd6rqxhOT2PwaPhb6dhWLW0hOAdzhDBmfdI9/aSSUVg2fXuObAcyUp
KdnvkqMIbytJlNkQ7TF65YYIjvFljGAtnlM51ia75KejNQMR2sqL1svGdzc/sNv2
DTxZiB5ncxCe6UcPUN2xk12Kaa8zm2EVDTJpPX7mojHu7x+Ae6uLI0cTbB7cNhJh
aW7VvPw7SHe8BiuyPO8jY8jG8dJnN6Q1opTeBV/I65NmL7+iXuV82vRSWb2Mu67z
XlGbYsuzJSjuCtZXt6uvjNAT5TsgbnIzmMoWanszTq3oGUjSgP6aOdoizH24cNd4
2LvhE/21Qb5sMFDgcMLojhq5m8sB/HDQM1HQ1seP9gUfkZJ2zLMIYTQFCvYVbcfs
Fp2qRcLKoBmrllvUnaZqiInXOuRD+SPtd1FpGJOdXJVDKDGevHf0z7JplvqJvqWt
LCX2KMquWqtqY5pJfGXjOs1ONflhtRbPE3Jet+p1uNUS3jXM1R8oLoBrEqRwdTmm
OaFApzyonxgMjC2HIwRsg9uDj3OWiNzxO1X3TKepY9Z7WC20o4nA2oQ/G+356KIH
wqbyyPlosqgIAbX5Mv4aUPd6cHewa5Hv2Nhh/V18xewx37tgHj/GdpQwrkZ5UtM7
gdzayZoxqM5lOA8srwvQhg5G1ta+gzvHb12vbJ5NmtZC9OlrvkqFbTOxVgt4a42I
sN71pRQjnos0WpCs+71Fwl/BAtUjINO7JZu4yw9mF0fzvmVlpc/EZa947Pf4CUHm
b+gsY7mtOex4Q5UlGH/QARKYIudgaf2SAVc5DCZzFC3OusJCFYBMW5drLUGJH5ly
6zyf7nTGCiv8tFy5H6XGy/tW6w/gCzVVVpitchGMNZNXPp5ILKgo5w2L9OS/5+Uk
I5f8igdogRzJGUiM0AaQb5TbamiTDvR1WvQKy89kW3fgp7torcvaouMqxGbTm6C8
IzIy/6ylstm3uWEgzlS+XBqkz3jbZlVKu5asyerknPowEqAtPZgJDdk7ig1OmDWv
ate+L8qYnEmNgw63WtOvMW3gE/TgbhtAXNEYd4sg61HUDU0rBJFkwQQ9oKmoPIRM
hCZQLAv8m7P1AXGKn+1IWXv9HIf68+7+DjSpQ0FBs5CLi/0rDz66cVo1lLP9SxQP
Vk+QlLZDDwTgvpK9ioNTJyRgKxo5fNkwwLlLK2h+QbAO5SbU7pd1vVhQCyJr56I0
SDk3dbHusi7ZI9laHZGlo6y5yXPHMrtLpyuKLVPtXg1lbkDSBU1OdVz+A5Q8JNc6
hE3E+M/pan+jfnLJJUYmXrfPVHCM2IAglb4Dexae9v9Lg/+nMhCXl1x6LWap92L8
6vkZLN3xndgZhGcOGcXubRU46HTjNCXmqmACf1FJD0IOv9okz0KdpOypk1RHEPaU
p3zAgnVm1UAzXRovxHswvvq8FQk9JdXTYnOZMs3nXMFUJXQwMR1vTOXg5+cJsrpy
FjkWL6Ac5ve9nDHLGvFQtIAlHZx80yYplWd9avzYz5LIILEYP9uNlNyv4oGHuKFt
F2oMKtGxE56QR5jHtZGHK8KPObfCSu4jqjVET2L12Bkwy6113v+5E+cvsDK5EPyA
rxUsOtAV8YkOGzLGgd/iN4av8PyZqR0vfK2mcGk8xlf/vFuGcwbzy7Xw8Ut+eAtM
l5dzulYSTk4bPPHDBtPvmbF8XAaDEiJzM7DFDDApcUxC/2ramRvPGg2DPoKG30Pg
X1zJb3lhq4A0jcQhEJOXUJUkUaz1b5Z4THkzctQPU1u2x3pC2Zr3zF5q1VWFquG3
W1ealuMHoxp09OfPwsLVE3pP7PaIC7R+3ydsnJIU0Vbllx217Mc8dujgaWPzt8BQ
qwtxRguxV6mQh1T3CFh9BOvNLi24RMBUfowuAbZjsgzcO4Ez/t4dfKcBU1KD3ygh
uFfZnL0VhD3EEbPtjSIpLLBt0ovVifwQ+2g5INyIK7FhtjUCx2BkdoRHox4GYQe+
HYqKEkQO2ceNrD2LiGmocvDNrCP2iQcRSx9S0JXf79ENHdEV1mTW2qElhCDYfxEj
4JBQbmm+nPgO0Lp1VRVZVn2yqaxSl4959ob9SQ/YUINBbVwWAfSHalQEYPTtJtXY
0P7o+TH8syuvx8b1m2l7gMLlQRUpwF6z0nZ/KYxAgvqy2ezFmCIvkY0CUFekDgZ3
PpgoGHeDGTMQuucsCl2LFOa7VP7AjyVRv9OmcRGknqUV9eYnu1EvMlXce18UJ9JX
rPAPilpDL5YrShsryW2iwOKXy+JlOzltE93i0gixs8UJTgJx725W2A7899UO7Eri
hzj4goaNZ/MiG9Zq60DTly+iFffV2HWlKVEZLw6MutYDtZqNHTZATaEUaWBeih+0
hU/vk1D2V2zxebfwe/WjQz7ugDjkha3Eppopr4oRV6UTuyEZl7R8iW1YydMWQ6OZ
tu/deYo/Uirmd3OdvQwKX1NYNI/0WasLVogqb8ur74alzJGwmXwS+2n2TxhxDH1l
BOkmwIbi2PIrQxtbsWLc/RqxByU8D1xKGg/hbA2Xg5Hx1K0kJrowpPvZr1LtQtFq
OnbzsoQoaaXWzRm9JZrbHAdIAXQ4BXPIj13gbCQIzHVuikzrGxEi7tSbWGl2/6SS
hxHo8TteziYLWHFDC2goWRcPEGwoLokptDWhEB52AW+D764P9LuKGQtRYkPhu7o+
E+NHJ5Hybuf2A7E9smLZoC101wBQ+2Rl5ouKP/LOYYfQyTALE1O6krcPHQaN0NFe
GKR8+BViylbU3y8w6MVN2e9yYZW1eu7dK95yj8NqdYUfZZ1qSif09LtJfx9z3NAx
bxEdMFJYUHmQe4zDjcN5ognDT1f2NHgaOED5nKpju1RdAo2Ppaffx0PVyWbbdZnc
Ng7VrPdRhK5kOcQyx4vI4kXezGIvqZ8WuoV7zyb4IDVZ6204s7IPOG5iGkHRWaBz
REVBWcQz3PPpZ9oKp6dhYL5oxFZ1JQEN0O6HcebpIWCj7VZOTFuAymtSP8+yZy7h
aGLPLDs/ggBTzAkSqxrRmpVD2MRzCpOz5X+gQmwOsb+zqNbIHBMLKiPO06c9ISnq
bn/tVTtg1qongwE4ODJoe8lnl7E1poSAaEn8SyoXMwJKyi8yqj596iQOh3mROlCZ
kICBSNoxkKdBsNxC104PswNA6QeajCCjdRh7NG9AQUV7DC/BbToD/vws0RMKeGa7
hqm1BirQ0+718d2oj5HhrCQG6zrCqYRG+S5Vh0SrCrFHvLx2ySAiK5geMgo6Gmyt
hSIxqqeww0xbxq0fA4oVbPL8Ob1XdHOXMve6Ic4x8ujSlu/FzsSsR1jqUISR4YUn
Y/B2rbrnfKN50rNWEkb63H9I60JBP75IQ1wsGRrS2rqOAtwVJXVQmjaBNRSQTU5z
qRLTMPKBDlT672ol0xVByM6cllW2v6OEvU+a3Gq9VvrvWBEBiEwqfnuyOsqr7/UD
nJpKm3Gb/kgajqlEOIYiKGXf6p/quakw1SBEefVUG6YamjVHB8k5MdSa8lnjqz95
7HLs2BVcDmcfzVg6aZnPkAp8krb5tLYtKW+KitOpmDLibqlnfS39Iexp138N1/te
pYAdn4rujKuHEjK69Du11s3c05hVJkpxheLUEUQBgU95bkm3jePQ+SwhmkHYqCIs
ZdIE0OirGDGnlKoTPOS1Kkm0tELzYgVeS+s5KXJSaX6OkpUc+Y7QOqUof0CYMUWt
JD7Ufe7D3YKvErsZEkVQ9VBztol2oLzAG+SE3fkALpj71zFvPBteDdz3wI0fZPNH
fhT/BUn1IX7P68lO4xo2MeCfaLXomaXPvd1oCkHwB5/qTEWX6xvAFNivZXpInoJP
mAh88qNEfVIp16Ws1Ghs9YcggFvv2DhLlLgl1eJMiVj/2JeAg+c6T9D1VhMZLbjZ
LPAcNEcmhpLfMZLrg9uI/W4qVCmklMBMKzQPyUpqCb1C4mBRwFY1g6aKP/MbE4u0
yZ78imjNj+wbtLdnQqgdx9irCAoMxXeTE4CFlQSJtvHNJ3blYOd5in8IxEEqTCpM
GhkEcFdR9uatz27vLCMmnjcDnwP7s9YRtJ28ludPWyWDcMwvYw4lGFW+8hQwYban
HIxEX6Pii4ll4G59vp3DG3xNbcj/uMmVe3RSx1ZnLLOzNcyTYPXEV1B74iDS1X4K
5zoR/GARWHanuW4ARCpUuzLGYzbOu+mTGPZ2T7WfOUr5dyLr44wrjRJTXcPrXmTW
yhUmA+Ag5RkxAuScKNUystMiiUssvxF7UHYSj/HfYJ06c4PhP0KPsy5NRvf/r3bl
m+62gmDO5xO/iBKSOKcLypwL4aFcxyk3XwAl4tNp4XiDzaAIBP7Yo3uaqCY7fFQB
9I5otBnuQ3yY6sr8XRg1tJdB6rdKIWGPbeZld5xtFzpYvpD6Ccw1vjV5P02tSL4m
rPfl5BZxmQ2MyC1A+lEQA4DzHQNjO6qkngmWlFvbt9RRPvzWLBSJFn2Roi76qT3P
08eJVGgI2l/DMMsr5Q+Wfbz4rmBj9WD8Oj4tB/zw0wOD5VnXpptJNDpr9Xx2AmW+
wsI7hDe6DLnhoRMsHNNtmUqDrOYCAIig8rI1nHfFEUoVt6qEGFQT5hFS0AWCmteg
czKQoHFpiioyP9AuUcbn6loNqP98MjRHHbmiHqxO8RjKVAjlrJRHPSzG7bQcQkWj
EWOmC68+Z2bSYqwc1l4QNgj3GInS7KDTGtLoorr/VZTNYEmyoCDgPruAhJ80QZGw
iJEMFXl5rylzpn5GGeHzqxmSYa8L9PQzin24l+/iNrZpXIDZl2c7SZKaEXwDB7Bj
0qlzq4dqDH5QzqvKL0MdTur4fte3G/ax4gelCGt8pmj3u3ebCYdB2o+XsJaftSd/
yI27++tXGSuvUvcswdbhk0KtQo+bubdorlCwcUcUAfa4VfCYwG6FeeE9nw/X6Cdj
dqmshdHid5Tb1bbmoAKmEEMNCAVQ51TlPXvxIijUCkW4nfssNflv/d+pdfGE2Afd
TBEsBAPhOBEuJyKlwkqUHB8lIu5HHHaUl6FwbXEjMDqI27XI2rwYIKYnWzmjJ5fH
2mJ2Bcdki/0xW1Gp7AxH123q5omHQsiMkk5zYRKVv4oMVDcxFBuegtu1X9FXD8hB
bE/K6469qE2xIOt4O+eCIY8FV3gqKLCwhy2px81iSNlPJkqhhzXdFkkhSylWcIeR
g5ARY7kC3DQvWmjPR2SkN7Yh4JbSU7h/aEoZgQ8SUUayB2BIcg/9whsN3jCM/Ugg
f3+Fnn2UQpOk0XuCI1uJKE5054fSeY7q38vC+5UuHgxdJBA1Ru6dDgwZz3wg0hKT
4HtsHrxmFfvalG2FFBsFL3JWKDsV1AJ7wPKHNcJo25uEbp/AJtXCQdQdaDeXkm5t
8OYUc5JnlpnXxiq9ujkx3gEVVJTNFWIH0TJ+vb8HNZ7Ho//eEVNQU6A06Q3K0p8A
cLBTVBdRUfmex6kZufaSpzIMNt+ZnCk2df/lug+V6iYpVsh7tIUt+FopdCICxtuK
VslhIb2F8/xpXrgahO0MC3mIf8bTXLbvO1jDCL2bGBbXM/5F74eY6bkE2m9GkfMF
W/hnT2z39FNhWWqUQ9D+zAGtFlf0HCE3/wINCQihNK4/qwJAoIjNMZOPVDWP59q/
9zgxIUHIu1uueXqHt43Mvx07IStqjhr4LcT0ELRHKoO6SqgPBjyrjjfmip7fgndC
DssVIZ9PIMwpG6/K3vkjW24R3OX4EcAM9WqFEaXXnHZNbQcJPfwRKB/6Dc70Qy0W
kFuZrl/vUg110w+7EBeDPUaDSxik2How18jOpX7KPPX3VLVvnUrZrjU7Y6kqSQFn
nlDHTcSIiyXImF+ZM/329wXh+dsqL7SpZr7zBPlK/sWQ4eD7Xz2tlOTuHlcGTROs
YBTr/AN/BF2v09OUasYuROKnQySSe1RV3/sYVYji+dNCQ0SBYHLxLlqSAuytv52H
4wXA3lBIWOPnkg9Zr2Rb52vpHkkF3/h5x9AY6DaxxFaO/wh1ezMYoyaYxokoMvz4
oMZ/mDdcPYF4BqkQ7mi63gE8egXACjFxXY1xKraiyeeFvyW88ij/H807XAJ28meN
NkJD6b8EoJ+wcb9KvYVVohSywzLx0MS9bOzg7derJ0Tg96gfeLia5KIra3Rn9B37
Y5YhiIazfVw2Zp5a6HW6N1jozNA0+YMglm4rLkKZqgIa6sLF0qer0SeyArn60p8o
8GYxweXtqy13n7BHL+dYHUuLPp8ouSGRwnLNpz3Dcp+NY9Qb6kbQoFJcxB0aWYZA
YxjS3tRm7oDwrMung13pgnRhMopIkyv9HsjoSDepFXXT941JNqsW+UTRQjTNJMFg
UvekvAiPL1GsWe4Gj0+iFEG5pKu0wxfrrxrojOh5SO55K/VzXyVUXfrn/IuXgGvS
zgH7dCyRJ0dNba+9vzJTo1CF0EaxyRfXrmF2MlTaqD4OFB43EdARDXVYYFB6k4ZU
ugUiTXCQa21WOBDVXr7htQQWFrKCzw2D2A90+TiG4ADM1+70q0mzwQ2cGJeTtQan
N3jkTen35tgUZVz82aX5POa9QK5ai3hbVIptJ1tUhDsuF+dgkOOYt5OtsYBDK5iA
dhD0BSHEnnF5+b4hPcDBKCJh6tW0SYAjbCtjECoOzP3mlPIm3+6Nath8V5XgMjPN
gUEqVWXLbSJjgzQk9wR6LvGuhBn/8chSIDmFJGRlI2+BwOHySfHNAuDpe4P5yvv8
x3SYzzYGyDlkc688uOm5ljC5TIIgXFX/AX/790hI2uMg//mS/9CBcuk0/1YBVoX7
cWnlJAR+Eb1tT8t1uWqJZCP4l4etsQn1y42GgVjgiOnOyQEPVNTLTDscw4V376FB
rQLUngrWewUbZiRr+Z3On5N2NL3iHoAayo1C9w4Sz+aSFd9QvNNmzWVRrywG35vV
v6UHbQG8d9hGddP9RHKqHVXGfE+sQ5KdaSZNZKCJ+CzVO+H1E5lpcyPYbSGSlKHR
zwYZklN0W6rkoaOAqkeh1+dBiXZOXkGKulX8od2qHZLBu0RYEEZALSYpRSNdDiWs
LWHfB35BQhfc4bhs8efyS4qY1quVG7xqGwya7qQE5PtteWCCKoGVGksqlqYCf5WO
jf7ET0KSt+lh7kcVHGESv4SDDgU6Xq0csmGnhic8JyNEgt8lFoiOo8nrF3z7EF0m
9bXVxup72oFWVNnza7ACL031iH9bplHmOgzBqXQmwyCnphFiUELK4jLz38RJbZXy
yx1DTFRXmy2md/vg49q/pHpUCjCK6FLBt4E0vTd12JQJKTLFMRNrweA7hU6uk87V
p0G/XL+GfS/+HAavuuvTZiGlAq7DR0l2y/YgQsQj6KggjMFp9+W7q3+jP37huKoF
ifD40AnYt6xbg8CPJL/pSYJ8p1xhuSZkgh5f0hYDy3t73Qc4bwLyPCQe4sFFthML
rQGOToyDuxhAj6+cYSfj2lNiILSb7jzWqQGmPGwRdkM2vnu+POgM/Hc1df/edWxG
4tLH4xio289ereUUD7HSQRh2wkJI9Ms8eWB3D/Hutha6as6n0zCNjpkhcbRvVo6C
y8WZfqnZAto01QQLiRMNd9xwi/tqpj69QVGOPMwv2mGAHd2COHkQQZsbf3iwlUXN
jQAM0ecpL/U0cukaob8kBvH21jhDZjTRXTyb+qEzM3r9xeCiZe9YqQk9uazDTRsV
fkyjPGNbwXYSdirbOfSOU9et4ZnTJJ1NCWQ6c9sM7murh5Cq0j4onOukUGU957/o
gBB5TWDSQ6joTKtzrMRWW+CB87MKuV8FZ0JVVCKmta8bCcCrmbsShbGXjpP1ZwrK
bAs5lP2Idq9x6Bvi2Ab+4lbdxXPJ7WnmMP/Kid5q274E9jsCdahPwZW+yZv/nyHB
Ulf/aB4/9CrjsMBn7ySAnOVmbtKtyNRUP2KP1xIfJp8F7dem4KAuMXa7zobvc0hS
+GwxO8zRO6VAfGpqKsA46OZzKZCW5v3KnwfWOxwSfHtB1fQHowNd40Guvzu1BEyj
ST2xG90LRLkF8rHxawHyaJ81B0Ghkug6q4EwJVupocjRLv22zXzwS96myatn9RH1
i86qgFBdTQlTj1fX+sSfHsnyDP2zcs7iiLrrF5LLIAVB8PPtn7mlQThMVsDhEKI5
amMHO4MhKJSHLiDzFwb+QFEUS1Ba7v8lbUwqQhjXueGnUnfC3hrXMVQiEQRXVINa
qrRGRt5sKZNquXUy6zVLsBt6RC+CNP8dIR3St1VBpX9R0EVjqK35QCRkciYv7ded
k0q9AMssR48PAxtbObnzvIXGIxYc4bIVBP2ZUWFl7GcjFWu28eKfoiY0EcNCGyJU
gb26cKuD9lHH2E0/WGQ3/8zCQZx2zH1DTBQuFS6vLux2w0ZsSwQAMapmJlgN7H6k
x8C5w+vK6JE4qjpdVeZvv9IJfi32Qze9wgBZptlStVOKcuKsC/A7CJt3SpaMSIbb
Tkv1zlBlHhQSrJf9xh61B8XTZ/D43mo3tRZKoFlclUbTT+SAOiDgaQ272A6MJNxi
7SZnEPm4zlMUz0vbKLvkUZm5wNNPIsyl/oFDCMOs4TotTjlUCoAL8JLwK7F8MVYV
XWQpg/9ce0X0wguUvnypa6FWzLuOBZIoCmMIS9FUlYSUL+okOCFBYCV8BvPIHl4M
E+NsvHBiZnLTFrkAludGX++EM2/ddnWe3Z+OOa06x4MhoqMtMmBdUgyqP3vqWG6e
89Ap4trM6dC2Qo1hJHxx21Hx3+v14hgtzLo3TaTwNKAFCo9Ax5yLxipQXJ3On028
jGKCm9agtTjlUgDMJVizN53uClLp+ObTBIZX/XiWgjdlPnYPll1HHbmXNMhvMH0J
LcPW6+JJbWo811FUXyRfVZR6wJGbBQc7da7wQq7oSZ3/tgbv0I5m0WWS3EtJhu87
ciq5Q6Tf8WH5opzvEnnrBJjswcm/noiQNPyFMbCLbZldE0TSTM6Rq0r06dlmvLM1
azFFwyVyLKSYXWQTCi6h6pFbjSZkbXxUn9yCjFVTbCm61FLaJMGDPNooOt1aXFeO
7us/60/gXjufrJIGwnANlnwDtFvf2qZkr9RChnAGVfr1sVFVClKTWKCDrHAZHjA6
QUaQYXFq6Netgz9P2Mg/To9dt29lqm821bywFwfsTBTUOGWH7pHNhz2su0EbyUTn
BsiRoP4YrnyjKrjfhEVRE25hOxUDZ3pbQg7N5h/o48k+6rO+5LKOTD0lMntiKlmS
yz/hnAzejgT2dAVy3I6fQsNhsrcABXTPGD36YqLiWoKxoLOc59af3glmONWvbmkb
2cZxvSpQrTFYU6RlP2vTkA4lveutS5V36BUaqwvsxJAtXZOKuThw3lZwNP7LawHB
xtYADkEO5wdyr5XqLkrrbsMREB+TByls/x8EXsX4USzNmHnwZb/Cl8qXb9ykE/vp
sJkyEGvD1FScWBCWPJM1cnhmjiBvMSjx2V5tlnwDxjvwsbBNUZCDWrgbNMUKNl/G
ijUNJVRuOxCg87pMP23O6AFyfRpxxx4zStnFgWatn4yhFLsU8pMn1uPGaA+wETXu
hA7LGofoe6qp7AcPpidc9qPOFtpSfBe0U8SgBsHQumg3sPXPmXNT1bejs0HdWyLX
xbkk8trYzTGx1YYxtbrAykRdBDYpLxIGJ5tW2yLT8lrMm08O1YQlPuvnXlvyrn/a
e5l6zHRNj/+5HWnYuZBgc8yxLn2ZOnABX04dt9jMX/rZ2EPSwg0gD0S3Tsbuu1WW
C9wwE2pLO6yKKoqTxgl69PzhuDEQ3tki9JLa9epsSuy4gKDtbdS9Tt1reQKw6jaD
9YAYVbV2hEq/IE9pYMVjo+qJHFLztZWteLZYdxZPkLXFPnOu7qlxieAhLQgNmAcr
vnrJegyrvXkih6IKhZkwkxfstQJ2lldjOzQ5H6IAXM5quxLw18RltQ8Hu+4+kyHO
tHXVleMt3nbodZKAPJXzSaLWbitABYfR786wO04DdT94NOJfQ67ePcuwYCtdV2oJ
L4hDkxIcynvr1MOg5QeT2jNJyneEWuxcS1z/6LkanmVoBtWehpze6PXF2ERNAfGz
S4a818RVLe/9Ogk3czd4B9G8/FGd6vErGEUr1QSwfyS95N8ZlCnyxDC4oxvCyeSu
+DAfkNRA7JanfbBJyi81frDzzjbeZsXzoK8LlL90b2IP3mJOplMpGb0xvNQFMF2H
ALDFse4w0trpoca/ZtD4z3jFKCvEG873lohgJqLLT9mSDKt5I8nfIOnITmj4E2P7
s/JQsioRgM1/pWOlh7q03sk1ygh8VPgb86x4+xdu+ksNYsC24V4itGWE3NPbPiqB
xMGA9/qyBW7aUSGERX6CYwKxSI6LFHdWLw5lx01WVGjfZcDFBi3/okYMHvhfc14D
yCJFtmIQH8LWSrrngP4Y9/3jM9bKdL6vILcL86KnHjkywUBV0MME14uGwTog3Di4
3QLkllAsLsUxDtnFj5ZY0v1962dIPUgwt4XrkY2qYLzJkf83rXWu11aur3CAV90s
TbV/pBvZYyBFUNxcj4mmY6FdMjGCGJWEajtcpfr5SunT2nKpsUyEF6sDZOHEQAIC
w7Ghk4w8U/8mJ/y0gcyEofNwpxtFZRy/kPmRSu4/8SKEQvO0afa8janeyQJvmzTo
OZbyVQGPQsp2xbV7OIfNsbJ8ZnqYKqtfDyfGiYe94nSb6kh1SiyWH4QtIwEu2eHb
42VTJSgRZmwpnCCAAzgCkpeeBfEBRk+ApUNZ6ljzw+FvO1lyAhsUYkkicHMOBeH3
2ibwFQxnB0STnL7H5jcslLxOaK7IYzJz9366GyLBP5tx7kScDR6QigJPSTyVZc+T
NwY/9Y/DYyAZ41z0gx/d7Is23RE6n+eDcUBx5cWlClxjevHKmizXCGi+P3G2r0bR
7rc2orLPzpqaJi5Cb6m2K+k4bvUdbmHlgL4j5bUNy5JyaWYJ7e/JiQFIFS9MSYy6
fAdqDIxW5y0sHt8dWFi6VBDeRJtGW/XaxOgdRVuK+IQOi6VTGwEcJfolDUdWNS9u
yCs/h+s3WPVjWSCImu+J24rsgB7zZI3xU/PgG5PzjkWp0zL8l/yiYF1pO0rnejjn
A6t+YIJLlMLoZmhQj2U9xue7/UhU5cVF5IhFghPjbSTVD1d7qk8GdXmRUbmflFE9
jiDs5PciVxfWqDatNB8T8dPWNAo7eTGinasXMXKxI6krhw0lSTnoLNPNmYsPW/KG
H7HdhkJnfO/yGaEcN/0NouZ6CW3vqKmSqIohC2yP1adYzJwMLsGQn8DSoF4roWuc
WgFQbcPRMGRV45swi58VvSmLh6sLQMxMkniSoI10jM6X8OSnOXR1kN8ZGDknXJEy
g/s1XSmn6lTMfaqPsILgJu917idh1z699hem/OyMcFwBqMeR3RswwGxUu6cTi6B+
j3Lem26Q72nSSntagmHvSrvUw/WocPyA0d07AWp5zRt2Q58CSQNaAcXOpGr2SfCY
VW9u7+AUYnKGZNuhqdPd/NUJumBihql3biLv2BTVao7NIM59VxksZpKZaHmTJTQ3
Hb00KFUd9c2AGOe7d9CrBUy6hte99ZWawabHuI23l99hB/IDN8z2WE1y/E2Ds5ux
R8idLQRAAqOSIH4EcHF5Ji/aHv4eUBKa/F/dA5hVNDuYn8mKzcKQAk42XXRj6Y3w
ON6EOaz0pPjCAk04tWt6kkv7zylZpmjw9CmkoX0c5Oz64KHXqn6czosZVN+RC38P
XHFfYxzldAgJr9e7ToVPCSMtsVFuOtowsqlUMt/eJanhny/VpjLUGkg2oBKSW6il
8B2pBsYGwckxv2hvoAtHQuKDMcb7Cuor3xHZLj6krjoiTltwxXrbMIc2FFnOyfy/
yNGPBsj2LftRB6ymZ1H3CzprC5UrDgSWZ2bR87XKWKJMYeWebMKNjD8WAKgyj9AD
W4H/no4zGOqxE9lh0ZUa8ZvU+uXzHvv3srdKeh5LnG03/lGUW65hSae5jAgpFGqd
0/pyUmjY2YS579+LoomGyYdL/nqNoApzOb/NaHJiQjKMB+YZpZU8fh/emsttm+Dy
WwOkHF0NTz1ifLmu2JyItz/ru336xR5ZetGvcl9ljfnq9KEiVrf/8wEUIYKPyCZ+
UPhOnYWjuWulwpRsG0/BjL9C01XuReciLbNiZNEGS1j1xSTNa4Lx2e+rNfsvvZzh
Rz1sJYWkpUARxYo2g6+R5ppx9m9tQ7HaL9nyPpWD2K2mHRkbb5E2jirL409VAMQ6
/PwXz7eD8eadIjbYfmpqZShmmA+chmmqktO6aZcz14Wqwne+rHusKOHXr/RGjmh7
vhs/6CqMqDZg2skuqWFztiKIn/VPhptIblaWQhshFoxV6H2fah8XpjF3Q8azhdJ1
1ZeKPYiDZngRWzVfb/G8Bii1WAf/M01pGyCCFkAyGqF4Hc2wySCOowwuyUiZNo03
974mZcHcAgi/q6fXgsoHNOeqHVTImuo6v3RX0GLdtlRc/hlZIxq+vHAx8J1NCJcE
0OkykXJTlRLMMMrBLHNutwCXiXUKJGdSw8OmIxaOHgn98zz8z6OO6mivBzVm/ZI8
puYmvzEOC+cB/pzUFm4XpqOsVc8kc6acHNvzU5yotmhFjs70ZXClpuvRuRzli/yL
ypI5PcCFCK7suvleXd0q2tPnPGHR7JdadAcMLv6lpYQkM5NEl27D8MgIv3R8+9zu
Cryct6I8+VG7F6zu6Cs/IU1ij0ey0LZ5AO9hBvJ/nprPoeFXaDyBb7sbOBZ6X2py
3Q/t2XVazA1G2RGW9FuSTLf7g8eGuXZ6+weomsAEe7Fsip2hOxuxaaD0gAhcpGHE
KkyP44WOOwW5yJschiU0dplZ/F2SJcf+3Gc0N2etKgAfRDIT+ILa+G/rgFv6NfMY
PHFOy7Jd/C2byUESzu1r56e8fB+nkI2emjhfjXABBCM5hSlrXHnwxXA0fjJyOAeG
4mlJnKRtOf7C2r9z7Yu+0/METGcFEHzwBD7XKYl1RG11MsK5xHsh4/otqu7BC+vh
ec0Mf+9gfyOH26kV0BSBb5pNTgX5HPzlGOWWxHWchJwLl8lMkVCHdqeUIuSidItp
qxRavSnZ353+Qkx0IwlTmjr65C1tJmFxmXtiVV514KGo8ryEFlAIZIK/GUe//Sy0
1airWHme0VtYgofaIJHLRBaw07d56T2Aue24fo9JuAUzgvlmck0KySmom7hDygu2
FYV4T61BGNvs8g+KwUtpDP+I0eRKOKFr2HDI/B/YM1hek34axhltk3CAAhlVV574
4smaNnbWJEjcozZdiLEgTiQ5tro/rE8REf7XGM4bsZvLAbF0NFTOmx0IDLT3DM2b
cogQ1UzxOzirsBZlBRQaiwOH9ViCY/X0WzQDbs8JzfmsZ7k2CQ7R6cylMtNMmJHQ
dvzwkSYU0hkusF72ILdo+5g7GDfWNJd/sW6ZTOZ5lRREb9tobhcOhICxyOMVB8t0
oLZWNaR1id1C07x51vXSOePdQiLTl+jbVK65GS0MCdDs+HYgejg0NDyf5fOfZldm
3Mlvw7WO9pT9ej8O95vedeKlgdw1oDIJXe78x49arW/rDIaDBNxn4d/cHXQN/nZM
1kWHQMS9chZ6LKVRN2GD0iEsJ91EEoO/wFSgIVUX8ekXE8mv5TibU74MewQTwckS
bWkXH9U8Mg/uhjaYA/xucL7gftjurnWVAmKKMpApZpyoNL7Dunn71UhWXssu9W1y
wIIZL4Tyk3yUdHducynXASo33KVxPdJ0izmirTMGOOKn9F4VsmnLdyYtyQUBnflc
DwX5YBWg9C+VsjWgZAIcCHsiLa5+HH15h9uq1GBj0N+x13bXVTz+3ITQ/8vIVcOx
V6DImVkmqZgG2hTaIhTmMVds/okyDuIYKMZnDweYKm9ssbZhfmoKb4OQPuEpSgLK
UDxbZu2WgCFICaxu+6vV2yYKpGSOR6gPX7QTolLAAOIROwj9IJvlUeoVldFbzRGU
fxeof3XoOlD/Dm+WuPIUQGYzWjXeMOWDFlW2UqGV4Km8NhNFxaYGvyjKRYUKqUH3
PuOPX3ZiB50CZjNICIxQC4Z4tsRvP/q3IDJMfl2Hgu/ShuP1MoYc3orljDkUVQ7s
nr5b1QEzYqI4xSbBiy5OPMEUO5sfh9E+y2Sz2e6KP0uqQY6+DoT0J3R29hJHudfU
kSGDkMuXYKyib5Czhfl2RUQMe9+bMl8oMs0LyI5y2kVcRgMbnFS0GSKheF7ZyXMF
dMutoBovUK61XkJsP1drjcZ0ZRuotXzU/rCdHfdFnJwtzTO00JnWRWWh/4YQRwJe
F7h2UUI9Xx+IoLZLIIwwk86hCH9w9JMmfn8RkBKqrTzgPbxQxFuG/dCRh/maSFfX
tLWxJ/rbEtA2GkYlpbqsYa1VObT3XAU/NEZJ1oLEUH43N9l8VlmYghTsSQnW6IBX
M6hzwneiVjgdfZSf9qXuBgUI7C0djNG5mmLktq6K+oIPnZBN2721uS/XijFAinjD
VS0SlGMX3eTyzBZTJ16nw49FV6zhsDehjHkRmLTEseFNthee3G13JeDjeDfMPsVE
v7xPoHX4uzzo5ediDddBTieNR6blpoJQk+iWqQlPA8Z17V9OGpsuH/DTmLnH7f3+
zAy0PaQpV4apIxX3egnH4e86NSQqtxvI7u7tUBEmVCgSHWzjirkk9qNuhFufmP6q
0wRIEAY88La6go5sl6CDVS7OGo8nIxJm3Hho4yuVJMGb8JFQ7RvFPD4dZSUAAX7L
KgXW4o2ElKIOzMpDjqxYLhFPjDIlCVtrLXDckCGOEtWSsHwJmhXqP4e2YTl1rK2f
dIGm1gdungwFLb3R6n0CjQVBCGqfuMvfff+ZVc3ZsDJsZS+2v68Q+R4Ik1IJj/74
C7+LI4WMuat17C7xJvUGlmhlMWzTcNGM7VmpODwM09ikSwVWHI13sZV2TVyLC0ag
N/xRgREe7dOha1wft42eE7VS3o4Vm5+KCefNv3EzKI/zaTlBxKBC/CSKUF0ASSoB
PlauJ24RKBHVaymXLSkfC0WMoXUYWMKZ1aXKXLv42enfGjHfBIRs9DQKiS7FPLaU
Ex2udvYquQNTDQEDlwU1KA2e7q8VhPDNhdFwqALsyjyrKCY+E4jzbCiQcvNLDDkN
0LRvLLsUEjbbkBLKEeI6dxXfgnzMzkXe/QEZxOGWmEdL8P+dPmA+nvP+AcOCb5Fw
3E+c9yL+YQ0zwMM8gwhEO5ylNfwz/RKKAUMY1yTaFcvx6wgdJrqyIKHbWdcXLDKk
A4tfauhOg4nmsXVjwLBfDsDoj1T7vrUttkQsOWcGSt4Zx3vVutn0rL1UQJJpLYLP
mWCILq7ABDJaUEculkOLYSvfsQJ/zCEg6Zm0BggwCYEjCwkSOqTIGgyDmUqhaF6d
7roj0dEDZC9RDOBXQ/4S3TxpyLPlRQmt9cpzZdFr4SN4OJRWldXl/lYW3kDIvImt
8IN9vHloxzMGMplkf+kQZCgDD+MUxuFY8cb1anh5zKoi4qPeIcZVFudVqqdBwHyn
CBTyb5hJqgTmGQYnL9R7sU7r7HvALxRKMPWuBtJZKLRttSEb0GvqsKu4mNoTVPc0
ex1d8Ad7MJOgwZuLS3Wf2rxsPT3lGEW23OxDASgN/UpBEXK9RycAps2CTstrHnoj
9tyO8ivJnLIuvFWiSFa/tRQT5BSPvioFZGg9yPUPSwdH47Am9WOrwKTq/qSXtA5w
uENcRCvCskN/uEQ0eOR0C80MWE7MqB17Fnile0pmgSvKJ/f5fNk8FQ+0j5xDRH7W
SgL5hJfmrFhSAjmWLLeTNNBaY6mtTUinVPbTH1i2uCGqbTGro6MXdjBAmQjMJPtz
sQ4BGaYPVY40uVo5HoUns6mWc7pp6zQ54Cqa0cX0VgWxPMb9KiIG4yGEWqYMjUFt
tqeRkCp/HzJInn4a/c5GTgACK8PWzgo0q8xPfDAws3ZFLz5BuKhraWoHKDyxJhAk
oY3ZPYIYTCCvo5qOrb1XK00OeD+YWJH0CJrmrgmR/ihhltzFeiw6S/evUVK5FUQc
GDdoqaFxtxqv/eKWgj9og1V+iL5QEtzZDgRTvT+Qqr2GfhLuObcrl/bqpv6rIqpx
lwajGbNma/Ix+fKdNS4AftjqIeNKhFY8lEG9TbSsH0/ZfH4dn+aWqmqJNDcxCSRZ
H0P1cPCCBuMaYGNLBCy9AUC/2Ctel4OkqC8952pQ5pBdNSvAx8waEFtRceqevqec
8zYKx6rhYyDyvuGcHuso7J7fNkQ1YUBR7Gc6WjBthpluFfnXliCzI3MpoOuZcd9V
8gP1LCcpFm3XTIMgr1AnSqVE4HL7ur3va1A3XG4ykE3ddMpP5GxWvUnRYjKtPapD
fYMOYW1J3W0p3g/0C0hEcbZkYZVTE4MfPdkwssDIRPLelv6JqDLMRWmyawLXfHBe
OXfMKqKq+YAmAvN9xH5hIdz+zgPiTitxBCsahCwj4axBaWfLHJwlNQbAX5NVsD8z
qMnwgmPrpeCu/wDz9nXPT2GuVkeUGjaWNz05HFBlbJucIUs9BogsXWjCjYu8dgOy
06hRSzJ9z4Y1KeWezSWYEOUylXwvDqZHOpPFsznuoZZlZXzI3qJWUwirLfx0Bwo7
s4tcbLVwP8eLnI8WXV0+HOlxjY0i7ShG43C6vCMwVGxARoL5LtsGwrABvuityMB0
z2tRkAV1C0Ls9p4SW5C9OlSdLEWS1VnALJwSQZni9+YvvMMH1xxfsqAmbUZWc4H4
fCu8rHaPDxk7rSpLhPAY49CwYyzGzviknl/1LdVXwGt3jlsMXDsFm7+OimVRpfAd
YtCYa/a8W3Pv/yuNpMHdVHsl8M0ozzMjQNCyWJ5477i6iOhe/ZDW+wAfCv2vwA9d
05DmydJjyDhPGsOJRQKaGPc36tEBRKdkPRfuMUSc7BDQZbGlKLCQEPA3XvQSsdhb
gr0LdIIvBYzBCBQRd8l5LBfbapscUp9Ma6jkJ9yvcsH6l0imsfHILY/533hiI4H/
Qowuer3IjBXm7rpEUcNc7jRugjgZ1CkhG+5wIY9FhoPqqNJssrRe9yN6jBBhAAyR
Zq/CS0+mpl4WTyeT/RqPCYM14/vH3xCNeY7WOZYn0YgZb+yX/rGRC2e1DjwaBrfX
xwseT50J9iP9DzxmlIYVZxpPgM46WSX+l58Jqd2Ify8I9WQnu5aAqTCyuXQOIOic
ospyiDTrSXcw5o/j8+0vlk4SuDnAdMiIcI64qFoUt4w+X+BcMenpFM6LCRi/MfZG
jpnYvxonLCB96nun6/ao5DIXe/M6gnNrWx37lZRx+Ot4sA0GambYvTYylHHFH/jH
vMDVSdt62hHf8JZkZhgmXIF0PewFK5bM7t2s6390rkJ+2i2sQSuBjHT8RGO8ZJ6i
S1TATqEJVrmSRrbGPEmwhkGkcx7+nmNZa0qRKpfJ3ZX0lHqyHbhXgoTOokJWcFJJ
m6Gu2vwAiv50WbKUPXCoJO700TQ1chpy9ascSOpmSBBZp6Q/PyBDTiM7mcVcAqUZ
d48wRipMUWFZd8WBRN4HYWo0WKkV+7Auaj9bKY9sfrqqhrtk8XEGanxjzrP3CU4T
5a5JKcKYKXDpJWYOcVNzl5fFRlb0ufE5t1HnVaDbvwiRQP5jMMK7IKscRV+rvuvb
yTNkoqxpgxvaZ7ikvoUyqLR0y516gD27R0ugGZE0pmQe9s+gcCGKF5ZqI8BNoMMh
015LjWhozgKDKIZq2p9XodP+HmP3w1X3bUTtUPMuiixGrkj1w3gbCf13fs2SqUge
vcPKwA22huTVDOdizEMHjH/3Mdwa8U0N58UXw0sjkTxgR3H3E3XdW7Y3fOLvdcaY
qf5EYF6AOC/9PtVlP7S4T/xMeEpBu7JDmAGib0JssrkrrDrAYK/2VR2cpQYNGOyo
PElwgj0o/z2sgKyrICVpzfYYxdNMEXvvmiQaf3KRM2wyfRYWIoAN7Npsc5PFFWP5
pVbEHTnBinaFVMUTdwvGEOnyuhEy0fowZ7bIJ3FKEhQsbdJmry2lSK6xufGhlPWl
4ykhrpA2aCvZZCz/8gvRfmTIkZN9D1N1lnx33bTedvA7SZyr7ZzFqvdq1ugsf08R
+ZFtYXQGwqsxBOx1Z+Ep+oQREsjflOtPD91YUOiVYVLafOfJx7aMOtlA36ruyIAw
LSET8zOJNJ1kcZmmi5GDQ9dcOA+ZD0CjcFtVkzDZn23vv2YMK0BA4YownZbufLKI
8fg3xCcREwAPM2bSYY4z32bqMtjB8PeaXVLCU+vGjj/LC19b3y4g8jUiKrtW7Zk4
FuH8NkMrfkGEPVZqbUa3BJUptqg11vZ5hUAq0bYIeeNr76qnRdLBnJSi/JoLjkfv
O+XBrIwNc67NlHrPIBJuHWavRGtvyS5dVb+J+VXWFEf0kgFuWkTv3dWnUqf9SDY8
yzDeG6dQzX8icy4CVBt5WAPheui5NjJwOyimNQCQxuGFg7IWs7fKSLN57J7LyR1I
HRN5kKaTU/VngWUV1/yR2gUk5oYapV9stcvjdf+QzPR2QjB3BoTE3kokf9BvRDgi
CaJmZ4liFmntRd/nh/JDOnDMHlj3TG948c74Z3YIE5mnAJGti1FWBV7rAOjEoA3k
qjDCOPEtJL4ZJEcgn3DoVQx3XpBV9PNoYjTNUqKxaGdrdM19mM1o8PY2z474hPNj
fcLXRZSMD3Zp+lxJI6KLxnZWIIsjFV71A7ty2AMUTY/QLG3c50rRPa4LoxGCZ+Sw
rCHBDyV1v2k0zsza0CgcE+B4gid2ZBvTdCJ6h05jpKWAmi3o+a+q4Eqfv8TxJJJC
+L31qlDBnYcbABtkOaze+rk8n28wk5QyMbQeFZpnYkqDD3UF6TYHbuP7sX0v4Foi
zHxbRsUBZcU6GWpkHhL1XTA2TcOHzQ7SCUCzwaYaezqPO12fl2JL3N3YDyWo0B1v
2vtJkIrsNWlGf/76saBwNioJI/86ddBq5xxHYVhdcUjyDkj0VBiVVI4MVlI6Jsvi
gxt7Yfpgjv1JuHPLdz24Iru2wPCMzPOMkDwI6swpSTWTW95TmxRI7Dx6Zy5uqia1
maQikVmyo6YRgrmGnIJeIYHgqWWgYeOCZKRba6d43mP4mVZtJTXHvf6koWtojds8
NitsGghHlSGtInfjVjghu4R5LVbFXBXnllMYHnQxZRpS4vX/ZYHKRtwZYbigP6tL
JHFtgTjvc34GQa6BbFfCWEWg5Zrvduar1udp8s+ZnNnOtSYSTntgCKSVx4W8bw0H
BIbKEq54bNeyHGqgHLqdG29XfaLBmiKas0LK337CyAAUNiQcFdLkF8kEBv83kd5R
aiWLUnEU0dgOxclKFMP5olfnISwkFPOZIH5NiMWm9GJ9BxF0TYIuc+Uvjl7kdQof
MGgNCu+rVeyPSN5y5CcB8qQvLHBfi80gxWpECHQ5WlWPeRVgP0jvqRyx3NcI6VbK
5FWgso2vytusSd18fQPmaonOa6eNz/7UIKu4HYxjRD/4QcoPVhAY3joiLGdYz6VR
kQGHnYvVVOD0H/mbmz5lnU8clS+d0TdVa7pmtxmBChAY6Mt1IwP/KaZVaUxb74OC
zIdMRL/eDb6+aWBil7buzg0c8K9lVH+BmYTHYTp9prESJuL5s9E7adkZM/AT0ghW
ooc7g6CGjGZE5uFr4n5vGMXMBwaxiK8EOQvTiTXXdgAYUVlQYIy1vkYG67FEpYg1
8DwsthOe/a4oMTyG2wq3OlDD5O8Kuy9C04ntL58zh8dCftqqY/dC7b7apV5rZRuF
9ka4p1a+bM4i4ms4hmZ2QJ1bAHqLW5kUOtGPTF6s+iLvNthS7xmSnmWMhxNnnhyZ
uM4+qYDs92YnSVc4HeqVSFWAGBaZOm3s8SvohkUFOmhGlG98VkW/2j6ffurLart1
0RkdG/Cdx/C1C1d2EQxVvEW+BlAuYbVupck1e+lIK9qkX0yseMeksuumtrTlx5Qm
l7yl55r530mQ/B/WJeTTXctsNsZtowbPQzNraJbhwn/oyMk8jx04QOXsaZhydoHC
4Wrk5jNhffGA+A1PCbfeABnVmtnH7H5ighk/HdS+P5lJO31oXWMeD9ghiNsd2gYD
+NmdV4HpDwdQ8uTxj1VKUwLAA9CRR9ge0BEg3XELhNjKJIJfJ6FhBsmbQdbr6xjo
dW+U2eysRX+CeQiqZnRnidJShQoYtgbKOYhepT0izdHsqO8475xyx518Nit4AjXz
RbN1Q2Cm9VDpqVN+1fq3YtUo5yGdQc4th7vjTB1qOF4zBaPn0H8oikmXkn/ZCy6P
eAHwLBJB9L5FXvoNKKvoguCBCoF1LUwwARPrIkPX5T0LvnL9RQhppab0felyA4tx
8+P0HoHlGdID38gM/SKkcUn3l1inzWF5jaBFRtyGK3h4wQEecUPNBcxqJqrJfxZj
9HvuHzUQlmKjvInFirEpKrE9eGYOhyMhkVWP7wlWEtLkpHMzkqdDFrk6lF6HX7OD
pt9l1o3ln8RSLhlpsyaxFJW/mmrBwTE4LIN8ANZyRpD2g0g+2YHD3hW0bSnkarqM
UZLR+jN3GDofGjtQiatzKj5D2Plx30CPoxMDg9rpRdm5OrKrNHo1EpaQzZShxewK
YwuQo/KD5eAYgGqomlNGvmHsvxcfUzZz/fKc68fVT1iLwvTwxHqpxP1cn8mcgR9G
g6m8pAwrjbXAVxvGW5ggpOELQGqZyyPW7mCkoguWXObfglTQ5ACuIuKVqC3qGTdV
B9Mk7o2A5rD/PuGXYYOWfF21cedgLIMaptOhfLodv+K+64f2209aoCaONTMxIJV3
DOnjTk06OXQe+EGkx8qec0dElelULfW2x/yk/AnkDk/lRUEAXGEwLDJeUAsCIBn6
yfkmj47L/MVRIynnehpssMgaqcHNeiAeDfLvbYtc+kVUOcX4A9anEVTSMSLty9fn
A098v275mBS8bZsJajNk//HR07/ucZWlESbVC78rJ30kQwsWLtTqB/VyC9+l59AE
GgNK/dLUOYAl4MnpQw2hFvIYQMGlbJVR+iMEnsDTrUvMFbsh5XVaG55HVlQnM248
F7VhzuB0F/7KR68msp8rvhmmXrk7MP8YwPVZ3x85fv3uBAEQW4qngxoX2DNnf3Bl
n2Kgsip5Q2ukQgfp47VZoprPe+X5cC6p9ZuG72D3hcmOkFpomay1QixVpC4/WUci
maKzVh+ZApvpWrxtYOEXZfq1Vrhrj9jl9YvaPRN0Q7c8+WIctTqcKgwci9+ojGbJ
WHy0kWNJgqjQ11mjFIN4ghduPwVSTu645WKcVu+ouwhRS32SOGQyjRmDg+HWnHA8
UfscieWj5IzFrleOe7lATn7I8dt9G9gyEJXy48pDpZP4xs1AO+nr6P3fPacEuC3a
YjavsSMiC8ze2gHire5H3fn+BXxvcpwSvajqpySUhK1sayJQsBSDsI5I3CETO69N
NPYF6ODyc6dF8O++tYog+j4+N0dlSHtEDpDQ+7y7Egdq3ZI279E/PS3GfNs+CmpF
uuYDyJ75tYSr8+fvPEUKVJY6WejiIvc80ykoviVYJtJeFjFg1hiiXE9dwPNSgchO
vAaUgTQ7KBWzIkGqgZ+5g0/hLj9lH+NigxDnIYVQfdysdgx8Pc7L2y1o7xUho4Ug
PafakHsuU5UV86PVbyWetmFo0FaBN/7f1bZNuq5lDaSvDPxgyvGNq5kUCW0LOtBH
z86XURsRtuO1iDwmgS2NnE1sekW1HAZDWNWRIFPEk722Dnn9dbbs4QiHTx1A7cHR
Gy7zXZWmoA0QU0Xs4tcCRHUqJEcf4TIJg4Y6/0O1r84e58NVNn3VMLPGV/wRNJi+
szVtxEQ2D+47n2gp8C3ZS55A8QsA/AZ73dSb5tTBuMgajA49ENiPfs2D3btAQy8S
ElbT19wAuQEMVQORlS/Q7n3hbNr0GQ/SSv8mGXlpL4NCYBfSsgG/213cS7nVSg4Q
BAEIyTR7uiW9L/6RLdHIFv1+Yxyr2OhrqQLz6lf9gHCq/kP4WDGD6Bzj798TZimz
EpDmc4YheeFM6AWzApGNFRk7BtD+pCuzU8Wzukah/hILfpnLTXlgj+3D8IEwOg/t
KNV/vq7MTG7LsNZJsr5q0XDnT+CgJCoUcErkfZZ7mIDWVf5uSANkfwCYrPsaOJ0W
TqEFAE8IHIpSDx/XGBzvh4mFTDgPRRE+gWxDwz3vKo0ZZswbRdDJjaTh34CofIaR
+h4JaEdclTtyN3o8KvOWrF8kq3/zkFY5skxcD5WtGA57ONS0W+pqvW19oeDKnFo0
ZBNxggo9Y/qhDX2Z0pSicpQLUZg+aOvQ+eAxSAI5ZZWHzI5W6cnnGZFCRTyQ42ek
MswParFTMED8/RgHFz7yuAWLevKReEO3kRjpsMSrcn/fxj1/BfzbluvEvBoRfeV+
LZSFTwdZrZBg3JU37Qg/i56c9NUiBtrICW4dsL8hLLeSW2MwT3ZfezkGsEENHyAu
oIJ6ELUJdjcvWlpADvbOQBzOAb+/voK934bWx4ReQCjKnFNs0v0X9D0rOQaDb585
6CRHnZ+Mwk0c0L0Vi+/6FrjIsRtyz+XtbhUV6uvH4bHUyQrBMa645V4UkTAFRiLA
zyZJ1Cl+FG3jJ37J8GqR2eIMMtsR1hwqOWyHddGD4726gcJpalGrbqaCtVzteF2+
P4qzIrSNOS0w7imVz0no3gNMM7PVaDWXpfYAqkOunz3YSDHY0fGc/wmaRGezLEcL
szF6ZlNTTN3F4m6VNe92D8XC9u3ihyai4rHMMt8lrAmSffIw5cKW0k3wIq9IV2xH
uhR4yeT49ZDo1VfXZWX5ECZQwOLP6/zbc3sUkZ4nwcg1dmew0gfk7I4z5x9pyLj3
la1yCKKnW/Pr8dVhFqtJx6cYDL431yczzTvfuhQ3VHebuO7qaubIgKk1GnqExGi8
erBA6ZpkaSf5S1Nybs+PnQOdEwZiOz0QMDxvXoQIQXI35Csmf4/q2Y5JFvZs42Re
uxfnxTZ7AVoPk9nuMLXGTs9rS55x7QXO0B4r+K+ZHx2FOwo8EisuReuyXY147fRx
FZYKKcg7Q7trZW8fx0+F07XZRn8+lL+WcF94OG1h0DSeRA/LaxJZUAwDmbypfm6/
n/rqgj69CJPFozx7KtoKENyvT1VmS0FY+uVD5nx0+UUpy68Bg2CPpHtrLRn+by/W
CtzaKExX5OWoVZTk7MBtcUngpa36llR+fk4uApyWSEvD9XlGOculNFfhQxuV1GkZ
WYH7yaQWYRDaglI5gXslodcxCWVEL9mSPA1LyNPje7JrrCwvGhN/IogoOSOclDNu
WjcbD+8jUsJKQV387cMzuDqpnjSfCfof5RKuZ0WjjnS/eWSnbLf7FFmuPGZqmfoI
NEK5wj/kpHVZRN3g6Wsle+ZmHvYYBPbBf2yPPkls02vHlR7Ey9rsy1PiFsYaaBim
MTOFKRK1KZpIyiiiCtUyhmYvRzqnXGMuhwjJAGua8mS31lzTu4zcAfnqR/1KDKB/
lIsB4O3NOnxGwBUkdigD+f4cxXMu+PEHkKEKymTxwbeR6ody6li5Vb4jzEIfYNe0
KoKZ0PkH2lbDpkR9xU5Fo3AUnxt7TByAIXspkhryutpXsg1i1o7deUGLFvo/6OTN
uwBQ1i+QTeOy7KDnBmKvKZ9mCLfF3s8dJ7+OFy+ppLjU7ylXKPz1Qg/4iCfsnFeO
Bq4c3BiOPdgNJWnIxROe+426J9zl3MJXkKbZ0ulRBNNXSFq5sVoLyPoZpy763xku
CjvPGQX00vIxEe0Fb/EnCXCENHf4/R72LzopR6uc66Tj+xYhgAQkOXGL2ksEQZHo
dTzpRexOKMaIELefxEy3R6+1iH3qAdmevyzDG17+U94VafLyIqkXZpCthJf0es81
OfOpA40OjpNIBLPwmJmaxCPgA8t8k9mN5Yae0dy7/nVw82xPDZL9hlY6fJeEtmqm
XBjpi71G9g3/1y+efxvwE1QJ1zXjADuclU1YC4P4CHh6zN/sTePehqxVXM/gE15b
i0D2EVukM7f5TR6pCy3sJv+QqRxKEojNS0sESPGYO7SQ+vcqvoU9hhKh9EnI5++e
75n2pINjfRXEGNpgwh5lV34vnAdr4M3f0phN1X+sId6gQ/QUoA4BVfnDOVq0ple6
xWfkS54e9TfKkl9vsMc1ebjDbEGsZoxKyDQuqvLRZMV7/KVVwqZ0ttLHQmabon7a
guPb3/3PODY+lvbI7p/GUgnbDtvhsHJSi/LcUDSVvUpT/QOVqJbYr+8b+qP8R9xk
ukNYL0CaYhfbDKks+exhjoGPLq11JEIEUm5KVUIWrn/w1kxobH9W/IaJ6GwcIakj
9iCOutM8rebc9ACiVScJ0bt1J4eUG7UM+b4NDfZQlO4ycW4uNm7WHwfkJStdViwU
7FqNs66mMB22MUDlig8DNeyrB1ZUA90ZwG2CsdXt0YXlOUR4jVyEsQH2R8M8ld5h
LMJdMWZN7WawAHh6ECyoDl4Ufx12I6P5p/eNrfHIhw9INoWheEhHrXC3GlH3YF7W
USmFB9lTRxO/mJAY7L9U9wN+MnHpn6AlwRHzBrTToGXfrZTX1XNoXFIRbxxL1P9n
QbFq3aClazYn1IJjdoVTGnztU/HAwbxY8K1ioJdt/YzsgZUvmqaV2nvPzafaTPpK
TiWOSVHrcyeT02snSlWZbrTIkoi+EP2xLqqS4zPFoqhEA7OqWH/7T+HYYcGp8Aye
pt3we8JHX64psaqe6o5fFXp1MvzTNJ+IWF755sLy6iIRpVj9qds4GofKM6rLzQZ/
y/74+l4TWCSTyv2mQaxDZ2KtXJu6IysQYZ/zsAV619kyO+C1EeWWvzYr7sSwbW7x
f8stjqbmWsNp3pOqhPgVdIt21dOoUB8Zvt383cO3nKo1hSOLiBDZduhIeKw7d9Ut
bOVvHhWRG42NuFoBHoQxDnkYCCOAmni55aFq1RlUQPkz0gNM6LdZqGqFRWEdt4Wk
9f43OpDNOYqCIQ2XZBuKNlxheaLsXSmJ+jidTITy/BxtrgCNGVmPN/9zkuCmF04o
S51zDIqqBId9IcqrCyOxc4zDUkzTgUdKwKOW0LlPCnWHCPjgo9cbT2WHi5VlCxM5
bhoU48iOg4wjDiWNGGLTgZFFm0THgr2MsM9xLF3HXsdR+ZToR485tB58nsVNSJv4
WwcpV8LueNqjNPwLj/qvXStj+e92PVygDp5EYEtXohp6/ElbqKfX1jYHObB6epE8
FhiZYRd1IQdEYGmJlPGkfnwtohcgVqaggYcnLrk+lI3+BehcTGxDhjcS5WpKU1z/
vJnRF9+CPcPjKCer61dJNknnCM+bx88KwoaK5514eqzLJgtDHifWzt+2AunU/fF7
3i23Kry/tagB7+UJzPoi3AFtevCkdwabb0naxBeEuqzCJvBGO5P92RGX796xNoe9
7ryXSPyQSuq5qPSkkWqKIYtgalv4RmxnzX59Ujh2P6MfsxYEd0IPOXneTsnobmms
cN120x45T9xSN01CczxZY8G3+ULbWyGVa2RwkJ37N6xjW4ZGaG0BbCxWhV6rtJ0a
GUHeox1/XkTzFjit+3v+SzAZmiKOd1FBDAXWu+ERZ2yqJLTgEbuOjHpWthV3Ybg4
XUCimnwWM9QDVkKcNaOk8eF28QlX6qKVw7Sgfx4jAWKEytCjePb1erQDAfN/Gvf1
a0b/cFQBr7xki9t8SE5LA1yT5+KGHvR5Fzl23tzy2BrgUZru6z0AQc5L1qXfJAcW
PfZCi/Cwl0yCj0WX6SCFgtJwn5+7Ty65D3S3Zis2its5+5d+TLdzJKes7EMctifB
GCKmwgbcJRSScxe1WdrZei0lO4XBrUgh2rXMiGzVEqZQo7jx1utLEcsgksSHry9a
rlGhPTkSs27ITL6iXhj0JbF1tFCFOyUD/h5LdtEdSnf+/WMpI8b2IFzYjlF7IUrE
6jVPsND43OHSN5teXjVF3Y+vNA6le7MTF/vqHk1Ccza+Jt6XX3xYHyBTC29UvP0O
ic6Ory+anmYmloSF9ziPejOpJ4FhWmq2wtuz34BPwspRwWbzddU0TnPzinUz9JaK
INXkNF9uOEw96HiuTmrj/vZ6wW9Y/q79ljMKJ4r8gScXc8tzio21fV8V1Tlkm3Tn
NIKycBZiqKTKR2HDwHHWsOSN8vL5XIJk4MNCBlskdoFk+Grazlt0+5ysLSmiLe5d
HSzDkuVnWa/ZBHnjOfq65pw8DbVIBCVXa829Foa/Nvm+SRUJYXB1K1nFNE8YGLxS
z3AdjBnEC9ZybxPaFVDsYe6Qu61RmR5NvnxjpRfb2M3I0+n8G+Zz8KP5VZsEFhZh
12l57dBPvtKjkXa9G5TqGICbxbbw/HudVcJLIlTk08njdU+PNoXxQ4tNq75k8FTm
QR8BY+kRBbA9ud82rVR9rMmtAJcie5lv0DPxP80UWJSNRaZgWoW7jmRh+pdxcJkM
o6UvcLo4D0Kfd7zVzX+19QUCMNUcm2gi7vZzXao0PunqwcZCFA8+KwnVAmozilwc
Pgq1AkA2LJLNRgU3Nrmtu/5c6a4F7IGZ1VX2u4Ubn0Lhv6/hVVjaNS6y/n4IJUyM
MZLcOFdCvfk8YFbATI6GtIVGHKQVNngYjksb4Y8188D+G10WsX7aKVvUm0SILt8f
npHJW/nfSqvLSeqMfr30gxUklezjo/ZwY8qsC053qy252YI2gQjFX7HPJrtMW2bv
G00AmEVWE8+8krMe5fVO34xwRKNCHmpHqtv8/qMt+NUZ+njwHCCR/cMDJkkhOwKG
8aIlxT4Ev8tIzx006mNub3GDoFd6C4+pP6WXtoCjf18Y9fjx6+/8MvnTYemITL2B
7f6jsGkzaO39eGoTiWpOKQR5IOI3TzzWCB8L4XzTqNKvoli7Bo8Ecgq8JIWJb1tH
oe5UK2gW2QW2+tutOx3ZzU8MYF6sO1ztaHYfKhZbt3NbP7PEkRUrxS20lHAMjHC+
O/ycwoeYhWvSWwRTi2ucevt9hnGTTeAPpiKubOrittVjJjmcpjKUf5zh9gCxTORH
CP0nFc3sKjpLrYRPvwAQ+8SWoZPeWzxgvIAePGvoxEjKjqJmR9MQMMOlw3W4ZUfU
q505gKjy3wnY/Wzn68Otr0TkCUOctlVPAtuWxNG/taLNxmUmS7pVobFF9VowLvJh
cheNQt7Ebfz1obv+w6DqibkOgChyCz3fyqhv61l6B78DWxqsMv4XbuHG5Fgc7JRi
y5JqpJykIQQU+ksfyk8mjW+o0mkfWrk90CKYA9Ok0rN5giXm5/wCmQK/YOcMpfqX
jiu/vANrFlRr/58QkTyUdciumeSpjkoHBeEzJV63wKCCA0PC5LzE3IE/h0uG4pe3
VioNd/FhqZ/D9ewOSCyC3SICW7yzLLnOk27tOT9soaaDvwYdZLlNTUVU60aAiV/8
fJWeNrGJmJSlFxyghYsSFCUfQgS5vx7WUYm89OTkfMMMl/E4veO+Y/drp4ut4EEg
JzJFp3mj1JLZ+r1dT+rq/Mi3ut/ipVjavOpLYU+tA/nMg9TPKKfCP3lZhhXrl2qy
QCNwMLXiuKC+S+9aESM9jcWILQgllkwZiLFkcHckqQ4zQRiJEdx2895qcS9xei7e
ALIz7d0k66B8vUlFaYROJnyxWQMWrgMPLORALxEmGFZncDsmP3m0DmhRjzmc+zo9
fyH8Z3o1FL7LOtqlQWSTOBb6MxeTfV3I7z55hqJ+nrCziAOvTkR93DjuiDUlC3KO
+PiHEo7WQ/z6fzSeG1s7Tggghi0VcfEnPDFNV7tmzFw/+mVOiIS53RnmsOlQpfmW
hHG4Dp4ERNQEfC9gWJ9sqfw2heQxKccfkOTsFpsFTsByveHiZ30JxM7Hl6Ii3fjR
Duu60zKFcpFfp20sIz+ITZ+b1Ms7/1/+jTnSTyG20xbclTPeH6iwOR/XWEytEMB8
GAK3m2ykGqv6WbEv+zPFlUVqTAdxwKoQSRJL/8JtTkly0b9S19QqFEncDS4Me8nz
prU2+akn36een24bP6C2FUUUwcw217Lo5V7eL6Ga6+QVfAdCe8MIlNrUuZ7tcvlX
Il55a6NRAn9mI6I0zTkAHDXKPhw+2QvTlxTvgtvEYKFZI0T/njoxwsjdHU18AeAt
XWcmmJPHj54sx62Z/Wd8uVgUuKgj8QuX0301igEBg4w3nyYm9csI+7tgacw6Wh+5
02xiY2CPlOhlW6At1kzFmBCy/+5kcntcFZaUeYhPHrklXN/RSfxalKHbFQTvYDR/
b2EJUjtqcW433Kg3i/8cvDMZBKpSVIFxDGMz8a26/Vumuo1hVPaTT8wL1WhuK7gQ
ZLBzIJD3WYuSZp9ldLATm5GYYUd5Rimua61ZyquT3eTWd0bUjVBQHPZbeEWnfUA4
7bFWy8k60yOX8kZadWprJm60aDGUGKP8Ei/BYQtdrIN3wUfyguJ7OKXOAX4aP3tc
efsd/dhzM0RUITIY/v5HJtkeap62/wRVAxLSjcQYaDEQMpHtJqo2JiPAF+chdvwd
aMCn4OUYVNpdxv++/lDBPSBa99bvMGlVF/3si0jRpVTJPfE4Pr12ML7mEk0wla79
w+5s1e4g04cHcHCWkECmbfykCV90fEWKz0BOXQeDRgfOBpgBnBMPJeshho5U2ok6
oFV6wysNHJJnWg0yo/Znz2iJmXkEdK3bpkAhLpOfBS1huvmXEq0UjUslEJ9/mn65
VNdfTONFmM/Md5XJAqPyiiKrQ7c/x1RFrbxXyU+40edQ3FTTeund4gKfavg5zcHh
FThQ2lIoyIdYsXHr8XoM19y1aRGATKBhPEFkQ7vwinWUWMmN3ikjMhIBxuYb3fVZ
pDKWLJY/Gbowq7EDrn8YCXG8kitLzQYZybjRkpK44oz0H9RyUobuBqDW7q8qpL9c
8hI1bTkXlf9M0+i4fAUGols32nmWbd3JPmeBnm1eRTWbkalwvRA5y2C2TCyanuFD
cJK4SYR0f7n8RLfVYXU8gGqZghmlS6hKZQgmFueoLxxJVr4Jym8uwLLOMUqhhzlW
HVv+zSwATvn78TZC8177pvaJRPSdPcfjCsPmNShjWEMcdjHrwT45xHXehnIwYRss
7QqoocR6jma3M7xbNgomGMM0nPxlb4Ey7PWeY7tXeRASn1X2dMY/8IgCgSjgvak7
geYypuAafQGMr8k9PMBH4qY4JoU/fH38XjHOv1vrs672xpQGqdBl/iWeJsVhUaPP
rU84EABXOp8kZafCsOuspMLkDGQDrW6WfYz/Ac0C13D5MrIuvdJCZZ6ELmxS2uKq
kDYdPkbH2Xb3duX3JNOIhcUmePEbJsRtnlv9kso47jmfpcH1hUQev3yCYiN1KxDJ
rCg3p+3Oox0Pf4yc7o2wqizlbE/PuSqmN6bRJJ/gjNmxJS2wAJMgLlvI/Yd9q7IK
t7I6Q+a8Wb+cy2z6Hy4uQaZ0R6/bb8DND6Uq3VeMvPteRLRPNWliUFX5a5SCDctT
3WQCCBPbc8yx0nj54igWnHofruEP1qr9xeEy8/mjYOcWf2FFM4cpJnVSCSBAECOE
Nsliv1tFvdB5yw5Mqz3g3kJl6Nz8hIiG5Edxwid6MM5WnNjlOyNfNRC0Aa5qN6Ht
fpEOyiblipo+rRuQVXkNb8X3fPmcRxJnOhRbsG3p5KUl8ARGTrM7bBTKQ0xpu32v
kEnT/ZWgR++KrBxTv+QjxFIQzjSsB/xdp4NvHLUSmUgvZ8uoKyhciXmmuM8alYM/
ofsG0Vt2Sy3otHSWBSpJ7R8wWzfCEwQNXkPho+68JKP7adZ885Gf2DXhBxrCfDOO
X/CdvlfedrfKktmNx6kLgLh/FEqVME1V8n8lYZY2+fUWizEbLsOLkTSNLlKdmapQ
thxayAuCyOcSDduK24tzApj3LxUUEip5mF9604hEQ1sd2axeMDs0N6lV/wgsQhRp
KcFI6CuwN6Jsvh+cVDO0MQUPgCThPt+YxZTf+5EAlh1uRu6qXvUtFjGCISV5GRn2
4ydH9ZeyoK795W4WlzrZbN1bqqMP15CKyFMzgrSmZb5m1K2tT31Sr5Hfgt+tHtHe
S1UkXEiS5q5R3BIidpUZJ3WIpYUvAwYyy6fxeIp7pVbk7fRyTD19+frKicCKOHDO
+K+S+ABPnQ9B+QdBu5kOs/2dcdOaZOM1lkX14lG/GE6WDhwEvpync2dVNBPS2ubB
qi8xvqrdCgBVKQzyx26Iz0ihIfhtIHnWTzfz0Q+WT6SaWviDCj2uaohjVvTBDMPy
Mba2pWj1ZqZVohrDddzf3c8am7gGh7vk87YNiBQxaBjOmQ56RIRmkuy5QfDFA98m
flwBQcVgnL8KHqrJTvWeT1rsVd4KaiqK+1P8d2XL3WCGDgmMgG+1v83V9m+FKg0M
L2GDa+xEDUzQJucg+PFbmZ0CGo1QCzsZU+B/OLevcNMDvblGyr8lJOJs0J0Dq2RV
xK1SqRkCfAeFzhapn0ws0B1f5rH+pmb88YzVfDi14fQwhVN6Z5qFEL2qxMN2/hZU
sv+9bkPBS8+yqoTHxyZDxiaNVxVzr6JtW563V09v5cNAbuEO7nAke1boFaRUfROW
HSCiIZAN7Lv43YcbQ4wN5AH9buUMtRWJFZRGJndrMe5A/Dgff4quf96uokDbk4c+
XTRxJ2U5VLSlRNs3ELqcYk7/WQkxE0vBeT4YBY7JBm58ZW15Di90FnWLs+hU8tbT
BtGmW9vJgFPMhRJMd2Z2o/glC/i333J3x2jJbILKnPb23firVm9NgToYbKMtGWz/
lGF/kyKb74EF5137/xt5HVyX1eCsFk/gZQGGqX9t4vAakg3VsYLj4XukYFQzrkNY
y2HBirfpvtTd9siB2bh2oLg6VaqjCwn1O70B8AIP0obRuuwqYi298aGa7xNCOZsg
oN+IBkVS8rAYs7M1maLs45XJXeic898dOnMgxSvQcCzsx+EnnLbva4js1mBX8M71
r+iK3a5ae7NwxpnBi9syJMD0tAu4ytDAo3WLVR9QNfzVLRzqGd/0DitxRVhDpezZ
NIWC4z2BkESOyv04Y4inGF/gb8eanuOjO57W77tPM8T3Rw6UNs8IY0d+N/Ghr4kz
QfWNiCVtqvCkdoFc/1/NWHh6pGPeE0j72htFa9BvasnVSjlMf67guNm012EPOxQ9
RrstmFxx1unQDAPW5gLdAxsIw7GsK5P+hD+JUkso/SxXWnYZe0z7qpABNg/MdX6e
D4hROKb7y4MtgA+RAck74MD9hZPeMR/4KyNzrVt9XPj7YH8fQWvEd4NhEmjC3XGF
56ZfOdn54tSNIv056VJYnrElvuMEtQCp7/XeanFrywodYft+ZbcuKPHl23Q79Vna
d79Zfw3OgDjqpisv4Ggj27ld9hNyq4AHBbeJ9wBcuCkBD8jQT5tI2IYj6nXZDD4u
NfrXZSptH64Pe+UHBCw0fQwFLfTpGOkVBt+LnBRDbDs7jBOTsmOdDN+kWqwWeAKB
LFyGoQkBuDBeYVV4gdviU9drZxYgzNUirDUh5fCzZmN2UtEWe7Ya5NnzYpVM148G
dFLtTSKAQin8s6oZU/o9NLffnrENF5yPXNeaBt2qzsPoyBz4duwtPLxJCpTVcBMh
MoBcZlC9dEzuBoDDg3WlyNn65hIooOFKcw9cZ70gtMnrW7CD33attSfIhzc/+0zn
zZsKfhu1fnEkcOUnby4vlkOhzIJ2KwdNbKPCHWg7BVAT6DjidAVBPH4KLnaRptXP
L5POhgXxZfs5KHUO4q40GHC3AtYJh63QyfyUu1tNpTxZonjPkQUCHpdcS3xvQdt5
nA3AAdv8JQlJ3JS2iyL94TqP35ak1mCGiNjjq7eBEalEnPUGsN7QOFvG5Or9fZNe
urNKvxmZre9xje9WfZGIaMZ2/6rl1nEOni18Wm7ixAV0jpdH5/EQxAKHmU5z4RNZ
IxucdIHT+QWzoYWezVDL/sZp2VCgrx0Qzjkd/VLFjT5S5iqb6lVVd4g3BCYWfxss
gvWJ7ojwT/6Yp/Nx2EmvuO2m6EqDrnk52zvg7Engfyl9VdK38zWKVXUpR6K6Kmcs
zwRGWuWYxXx+mVrVdpZMEKI2eS+72T1V2YkJiSloazeIhXgMfOQA8UMP/rv2kOFc
8oPz9E9ajM4/+fHBzXJfGM8YPcA6ybgpzZfjiO5G4Nfcl3cdofUtcyjYAGP9cxT8
8kfHtNGb97Jk7PZGHBrlYRzAtKvPYQ4bk6LUEgh5o/froCwJzBentrD4wpNs6r6p
Sz8g9nlSyVs1KNPS7Xeb5aVKA0PNz8m48Y1FlxtvJ1BQeRo3Hi5SoWyvEL4sJtk5
5H5MDHR+TszojS0JL4FPzOXjIjaOx7UQ2pxMIT6fdSAq6PDKrl1s3aBH8oqfsoE1
epebWJcVmZ0mMJzHvIp+djUJ2h3dYC8htpXHySmNNfPojPI89/4+nq/4G2YDnX/J
dGmf4xmlw0VRzI4izrNni0Tv7qa0IRNmxwo/v5qEO2QzuimjW3ScCnX1V4mQmS1C
9mwLf0vQWVkiuSA0+CIvpj1SF8aSCTtCdeFcaDR2F5F6AAonZMvu+RAB8ysFlLne
UBdjPxUgQk6lJkUf4Qd7yBrHo+aYSufoq+eCVLPmmws5OL/eXcaZI0auwNxhKLLt
nF8TVqUzosSkL+JSrnjGXLWVnag8zL7H795j4gPCtbIAGk3TU8g/q/yHn+h41tsp
oaP4h5uNaVqKIgbp3wW2GB2jfMy/aQ4syF/5QIxTkInBdmW8i2n7yd3Ke+pjygDS
L5RQrFC3pDFMsXNi/atoL8/hbaj4WD8nGRJTrImraJNSmu6QJGVJSMmAitpE7tJ9
EgcHYslU1iZRB28V3hcRWY1tzttLclDQwVOLAokkXtKfdX9KM8G7z+Zt1zqGWDTV
pFUorNq3FmKUfnvheoIcfYyFSHE9WtxjfB8u5MrnHSFKGXcHAOtNjwqHJ9VM4g+k
BEwnw6VzJRDsPQH0loTN6ucHaQNWWO3Eu7vgpgbfs6h5Z1lKj9WluHdI1L0hSC4M
8mOnvPJdemSnYa0B5h+6NGKXAx/aUaDbjq0CaAjOz4dT3TIsSvOXOjZw/Vej9Vej
ubIEQxZmmVMOtVXDJci/7/OT6ngwdwMMf/FkTyno7wlb+ANnoRLyBnGsHAwcWnv4
x86Fj0yr4HJfyv9U/3mss3ff78XATOOANnjSljnb83+MKuh8lkFoSsQ7SGypT4c9
H23L5umAagY38oBvFyfT1BKYCfXEbIewOxTyF1AWnrEIFQ6d7xUYcaXehgMMbz96
u2VY+LgXcmBKgkrEBWGJRBLCn2RmV/u2AfRPmrh6qZsmOPTwSwgQQ8KLQQx5ucq3
njBDtQ1Jgkrn8tUPaKf+CH6VFPGUa2poEXUVPQw1r9QWVhx3hYtyKULN9CrF2kEk
Vqr1SejnPe1nPmGxPZ/eT7VGcp3G27NABupNOj0QuY5AkcT/G6JC4ER5A2Bce3jH
1Lh20dmdx7XeRYKLNQLglHx6GF5SNXBjvi99Rk/DGxM/c8thz/1HeJvVhDtB5yFO
zOEefPvZ+8RtgjywrumKODXTPgdZc6huAq9Vnqo75K4wR1as/kaSPfiQKZTtP313
eSy09SSBgVgJRLAupKyBksZyL3qre4gPReYJCN8otMmv46wm6a8McxwtlCymYPh+
nstnAPxntmSiSqtQg8FGc27GrdbEHh0xo/fFOP4/wKK2149/k32dYKonDwav48Ig
Ng24Mv0ubYtR86AMmb0MYQ3bGB0JiiKL/kaKdNVcuNhjAbH1/7JAWWfGwckv4ju4
JTkNUUWCIxShFuuidgKiCia0gc/MR4kGpA4OR82PghQpPsyqoZJ3IMTDu2svBUJn
sP8UrkgV/cPB7oniWJkKtYpxDHSHzRzTJg7XzKIkNVxgH2rlJ8ehXZmw8RrWdeuD
maF8YIwbGOTK1g2NhWA1GBZtwXK6r9gLup2Tx5tD44c+YEzscegQdgbw4t3i5s0p
/XAhxNn1xI08Oigop7gA0ZI4hI0q3nq0QkjceD1TxoUQN9rHrRSrN1D/4FcJHFbO
7xR0olw9sOVKcwcAaubWA12GvsVi4qkrxjrATjBmLyzxot7osG+BFwg/O0BmxM7r
391Duo2EVK95xKSWD1fTTjJvpmQhzqhFje8IXIXP3/0iV2UNqgMxiAXZBuGjJdAy
EXaoDfVbiuiP4y6JfUPZ3uEt/lwtN0VRu07uttvK+qcckASV9G066h//fb9NypBC
dJWEgJ1ObOdFcAxli2J4RwuvhN7MEUx00HtVkSvRGNZwsYKKortZPIU8AcT+joaz
nEmQyaJ/olcLG804dcjklYvVJzvm7zT/KrltxKzXz5IzJaNdWgdul/ae875G91Oz
rnF0/YqXCKP1FPOZHOAuWpZmMNCsIYKJyh0m7cwP22yJHXdKHmH/87MOPioR89QL
iYP0G8zE9kqvD+2QngYgV0mc4ook5Xu4l8vOzyOWbyKp69+yU2HLA5TQSNgRqhld
q6ua/mwuQCnNYxrgI1RKtgaArn1uqF/+qbdP4sTRQpR0X8ONRIanRFraohf2SbjK
TknMK6glUKHGb3R1uXhvwWphGb7k+y54vf4iPohOfg+eCj8awcMnlz6Y+SdTWM2L
UZRt4auZR7WRHX+xl8gasQ1dDcVTeXm7PeljkbCm+DOKpPBnpW8KlD8YFSu8Tpsf
GMcYu7siobYCY9oDqxLgcpQuTTzEv0cmY45LEpgQ5JDQqWG1l86RYfjKjaw6Xy0s
F9NA2TwsAA3HulXOeAX6WQQSBybnumr7CSnNpe9hMo1Xy+2rUIwPuu5Cm23z8jM/
eCmiHrprRFlA6juXkI2SDFy95D520BvcZU8PR9L3LnjkS1YjaJPr4oQ91I3lUQxU
lIIjSXORxjoXjuDkO98LQghVeHY3FkkBkBMlVSigoS8GJjCSDg3t6z+EE2MhucQL
mGF9+2nVWwnOGY+atYCeg0TpVgGykTlARdF0VUrpzDLL29yJg6rWbYr9HIuqJG3o
YGl5qwRlmWnsgypdMYaqZ1SRKoFh24EXcT7uqhJ05l2ec5gGGbqAbs5IRMvBtIjT
FQb4cEgXT1nH0DJ3wmVnZDuOy8JQ/De1m9ru4yF5yB7TxFDmsHMx7zjCDsYFO2GM
N+sFy7Zsw/Q83GPoUi2NSmihRB9xOBi3XPzeZn1ywU817GDKmIuuRfZtymX/xBIo
QR1F9MKhpvaeY2IUSoCow9SwOQdrvNn4nqr2pkBfpKBWsOQJsc1AUiTCX+fXx41A
XeMINW0elFecjaZy3LMKW1ecCYrjBXEZp50s5K6qmBoNVO+QPiRe2Nco1jNERi+/
1xS7qsYUIc+u3jPUMNRQiAWysXRAbstcGjQdRLDCQWeSFOMikHQH+AiUC5Df9Il+
4pX7E1EAkrtl0Srrz+vtW5UX7Du9FWY4y688sscoIaZ6GbWZs3qG7lrMoncCcH9m
K1MvHD4FdS9zQC/CUCm3eEN/3H/1PElyHlbMW1g7lx5VIlFF/xDdLRN4KmJT4lZQ
iujz7a1ua2r0APmFwnFmGsa9oKI52j/VkZa1O26M+z6ABiLWdkcjTwQrn/hFFggL
vkWxpPr4vdbSbpp0Pw66mn4WxYa1Xqj0S6qhD1cyU5oSzQOMPv1TyvGv/C4E6R8m
rntZLsWSeNuKpT10JacH5FLkUhhhgaf9EpF/81hZCcWlQaGgGKLNyjngVRwcklBf
OJuxy/ITOnZtoPtqQKK/aGFe0UxR1R27d9adYGe9kKz2qBUokZrPTeP2Y0ilYsGO
SxTFOxLdwVM0qnSVPi8PbpFH+Y8HG1CxdmZZpkpW2zcWro1wmmq+fHCYPxcn/5Qc
L+/9iZN0TUCVKzhz2RgfW76mY9kVM86l/lGUWhJwZLPmtfvVk5oY4nd8xYtnZE1H
aBnyhBDtfGjbXYZWO8JNIyrKkWWkYJdWjTcCcbh5bLnC7RFfUbB0iAGfcoB9eaDo
BPqrPcyZRi21WJ09ZEaiioa+ZMCjI0gvwOrIpXnC+LqGDjQIxTJDj5kChF1b9WvK
z2U9/oe8GQy5SAXIS0GFcy/R0M5HRFDKwctSat8CuP0Zchm4CYAF93SYblNuQy4p
sclDMymkksOPRjs71WF9n5GnP10yB7P4/mkQAQOywWN8OKtCybPYc1r1etnpDRgs
tcPxh7l2AfiIlFibGr5JjOphpRIvXBENF44e6ClA/WUYsPIhr9rwDxVtQpX3SvW8
FI0RBImYEI96D65arPFcYUCKyagadJ41hdAwN5EaGSRBQHlXyVPlr7CQ0uVgif+o
eiKxBDgLGI2Z1KwetrHvr9NUuE1od1eTl1MCYfnSSP7pVvRQuJYnug4i9fr7NcdZ
qZstFepD8ko/gyM83qaBvdHXr2luU32sHEor97XgFtrcn3Cx2J08CD8LiKSnoJPe
VlJj25XEElJwmBsF5H4gbe72uoib7aBejnnFZAEKBJVdFwhVsKOMJjFM+7maU8C7
W0NWPc6y6UM75dZJTC0qJLL+B7VdyNzGxyiGAMKuHUriDPcL9gGNSOBB3sgIaWrm
4hmfWxEXVb+gUXrFyAFcJ/hesRld2nbCphMcOgM9NdkyrrjiDUYD+Or9ORowlaBV
OA+gfmnUTG6taOcfcNo1LA67p1YlAS9YcfH0aRsHzloHmQ8DBJW2U1iEdvfBKLhc
96W2CLWiPdkcXGYgJQswZr7xYdK/kvDuOoiZeri23C4RbUNKO1j2QuTjD1uvxUCl
kdLj+6z5Y3xj8TPdzqTPLXT3yYDMQQiHp1PUeAWCz+WK0d16S10b83euV0Gq2VgC
3fVp9YD2uZo802qw7O6+dLEFXn1utguEWVgO57KDWIaEYc0bi0GI7mXgCqL51zZF
RS0f0SLRlbnRpS+PwsDpujKJ8hA3cGCN1d3xziSabTGeD10ov53gk0ESx+Pk0j52
RGKYdNdK2cQY1UzDBYszm/EP2JA0TZJVL7fXzA7PJXP5rSUk/NHRvYIgbSOKalKk
+TYZp6jkIHAo26KaAqmEZAx8uS8OyziFI93skReVccLqsJcvEkeYn2IFCpzuIq7a
EWpl4XduzJHkAjiPniCSqqxuVhHE+WM/CGL89ZrRgyoQ3kquTZIwVFE6Co2zcX2g
3h8VgEJ/KyFPCdKcvvSktBOF+bYRJx6iVolYVBu9i2WVLfG05Bg8JhgMPDflE0Pf
FK9lNp+frAaAB6JdZm4YeX0LkhOoa2uZ0mxwSdsQEDQTJ8SeEqCyEt24PlzdcTqS
0Ba7zLQURoEm4imNl7/bqAy/czV4grhqh2RsdJfg/lssyY5l7DI6z4F8bx1qNaIG
e+gAlUwX8LMUPZscHa9C51y+LRCjqF4zzfBcMW6ibE2i8T81PQnVoPf1c8VLmlyu
6IotNGtwFgChgNU1jEJy9wLMhMXsLAPa64knT6oQfCh4f1W5UF6uRArgpcAssTRU
ZVMfsc/03HXondQRHfVIiMnKewr46UaopyByNeKybJJ7QQ/htEQ4cQyg0KHrJ/t5
Z1EkEbGfQupxKGi2vO8Rmpnf4suNZ/gkKLfZla8qMg0EhnLTzK19Meco651c5dEN
ohTlRy+AoVACwDdh3MsYjhUD+VX5jWqXEwQqTkjkk2POjICs+rhD9bWln06cMVuy
Ignm3OcEupezBqkU0aZg8bP1qW4eBKBOoaCZn13yOUfrNNxKQyDJ75Zask3V7ET1
KwVjA7hyBIO4zPtV5xMZ4MHE53wLOkPJNJnqdr+qJ89zP34V1KS7qkmasQYIbLYJ
CBU4ePT/7xfbh/C0VOGdQusMOKj6YC8GHs84MsePAlDUAM2M5fHEWCCTSWtwDwjD
eLcS70ghuPgEecxRGt6NZmILsMLPP+ZAs2hzrnJXQVTZbB23SsThC1BEAGE0HLPt
Sb7I840G8lBwZ+c7AMbabMPAx+sR5ojYFzuJN4K5SrbggXR/XpPswr2idX7xrZFX
eXlQ/oiM+e3KefDNP2M26HXMlrKpzPQwljJU/VU4Y29jqejtcv7mmpPrMP4pJbzf
zDEcG1I7SNp9QDGJJnTNMoax4GxVt7rZvR05OA5oC4xThAXK7xSF8BWzhb2IsRJ/
FchDoavjrydlLTmgWl0CqASCWk4yVmldlwUfy3h3kD5TPaojvzXqdSz52H8Bh+p9
gGCX9yK0++XQaUEUWz+4yKX2zdTBPFZ00k/gCRFWAw1VHBCXtlTzLokTDHKR/3Ca
6c5B5acwdCNMXhl0mPfUsTtexjGNp7tpdg2lmeosJUMYeE0+QbBMn3k9nEMwat78
hoF69j9W4v5mtfGf6x+hWW8GuW+v+nL+BWtIPYqOc9tcCym/oFuUN1UY/7jEkvFV
m8ddDnRH4HIrba8GEXrL46rz2KTIrQW5b4LGpnV2ADzifqsXatUpwi3FFKJbxQZl
bWpjNEFZ1Tn/CwvtdLgeuYRy6HFzl6T5VCnxnruuM7sd7X+2Ue2zrOsTNs7VGJ4j
AaCp+lObmA7DHnd7zjXTFz4L3Flbv4Wacn/eOFYOv1oNdGfO2lb1AGsNVTX9nrtz
pDR1xgAaHaBqUZiCwoKmIftbNJYpzp+XVqcNjA5Wyf9CwWpy40t9eBDQ9ze5tnbM
8mbneOgyqBUz0hfQahDMo8syrQgB+QrV8cYp3cYUWgGBCjOCISghmNk1HCIoVj4Q
4gu5ThjzIGeg/pzm6beyDFDpPnZlAXRQyFIEbumBVYjRkYz915taSZGo5DuYH09H
xobfO6ms4iz89XERpuW2gb1qn9WIQbj1DzFQkEqFACG6y0M/PaVfNUZCqN4IuxGq
iL2k4G0JdD4lTC/dllnVLiWAyYk8br6lJ+xEIe88PzXaG8r+RU2mE3KvFLAUPI3Q
lBbNG9k7lurr8g3C2D75nosAxCx5rBqpoIXBfE6sj/oeW0U4/v6gifxysU4Wr1/F
xO4BmtAfWDW65NfFVY6IqzW4wDiAlcg5OawFnQo62i31Ww1oUylJeUv77fWqZkdC
a2xJFyRxz5yAc0z5hr9jwT3CGFkPEHBc/brFxaMoLXkqExZ0Tq0YE6R6PNbXEPLm
6nzeaICbumseHLmBD/wNTUZZWkAWBtJGUH8sdDHRmjlD3HQP+JfidSHOm07wpi/e
6K9/nADVs/hOlwbobEfKQ8lolwfdE/2Ms95UL0sPLXVYVp+k6KcWtB0rZ8CfFMlW
hPV4yQOtT6sxuGOOVpoIw5VEw087EPxd7KeB2GlKuqduoJP2OcdMBcy7zQu5gpiu
h6TmgePutZVJ0Ghk3nJNosQI1CKPeYoV6+1jkabawxvVqAWkd1nivV5faTeyRs3P
rHWy3FMKHd1MvPsfJuhaY7fMcKoCtyCN4P0SH8TQqifpnbfXJoADf4hiFTBz4Mpl
bZSkbT5IHEVe3K11I/aa5aBZgjbLieiPJFHuMD6Q0OW/UVJw/ri2YlMjoW2mt+1d
Nt3KoQCXt0YpXXztrLGDasnk7o9nO7HV0UH956vbeR7bO9dzaCDVwTDwxzLRcohU
+CdvSL5HJAejAeRx50QPVHJaJ7EADYn5ampyb20tl2o8b+D5oKPLsYusQI951a/m
q4/4J2Ce0Da7EliAwytarcLr6kJmKwruCDou3og4bbNXlgEaH3XMzlYDSdZTQKMq
APg8w1rFJHGpcfDWEI2hD/kyp/l9uSp+oeUttspYytF42uo3yhmOP269wT2D8VvZ
pcTp0a2ps1tACUlfkcqby5mSSvPApMT5i5qxEFmcNBiJAgV34Ngiv4/B14WQFKu8
GhjEB0m3C3fxJv2xfSuAAcT57/Wv2ZLBhraO+J+0hgtIFw1RrVXUP2mVF5YUjWg9
aaMHw+je6ALqjl5XSw/UN340+EoLve0rDoY767rN6TqNATp6RNOW5cAbqyizY9vL
WJhnKbk1NHBD3w9vLlTE6i0BU0kCGFfjpx909SYdAJFifErLpnk+RK6tmRARfEEN
JDdFdql13/ddAx978GwXhmiSIpUrJfHJlTH2/Y3GSZSvqx4WVIRkh2b1TOFLIWIp
HmIE0zkJd4bRKkwDG2P9ww7fwBFSpLEdPhJ3/c4Pjno391dZqR4a7IhVQ4mqir1l
A+1hPYGeL1vNygx4AbUJF0Jr0V5UX8G9L1WmXdNU4VsVwuBlh7CSkX8c9jXBRQST
lnV+FZsRLetTdNbRZ5QR8PRH5lukrAVXOcsAwgsS6BF6iLf33j0YXm0kxoF2/CUA
LZh1gNTLXxBdagtVKBkOPlQNxph03yJczsbNg2RJmJpSTS121NVMIxb0KWNBCuRV
gTmZcB9H0Xg56w/tDNzNNZ7eVWt9cbEGRjJ7SV4LsrOuxqunG/zu27MbI7S0AhKr
oRgBvDcuq10wbGevY9xHOniy5ufiGXUF4Mcc68j+Cvfq5wvKic9Nl+qVI1m1dbLu
d/0BNLDwnZVj2rgGx5rAixBu3LBl2lPOYNkkxk5FThzJ5m1HtbjHuRNBHPjzL0l8
pqdHTBW4FxLdbWZiV7/GLTnyug11KwrJm2x/GyoZbGHKmKrFf3CghsuYC2GXmpsw
8ff9WOvHgwLfr5AzBD0zcFW3TnktK9Y0SHtAlHaZKz4/gxZxdR26GJKeBTCAgFA2
F+meNsGWzSrsLtvk1qeHHh13V+C8buFwlAtl0OsEaddTG6X5bsvkCCGfI1g6xpbT
IrfxBD+ZvoKR7VbwkAMDlr8S6UYWvlbReHbueXdRYg/qMnzNLeqOJ7ZrHuA6lO+K
cpZxFkhovM+OyRAgNtXNMm/zKWmq/QPJVPCV4POg8D8VtNerPmqW5RRE2sKT8Rxs
rqltUWy4khXZZG8DZTJ74yLu9KY1tkWWPfDIGeReoN5jnf4U3t262YZbEX2BlHT5
TRPJPEXyIFS49Q0WE7Si7chsBRuui4hF7haYGuwAMxDVzZ+EveeDLJ30NhFMYNM3
7TgQratLYsKRQGBP7G4LW4TN/iOml8Tkopj3ddbpEPzrw+4aj6enhh1/FAxz10Yp
w/dfPN+jIu77HKVIZZFG3JqpFaFovT0VPngjJHBlNSg2kTxNL0UJ6icE7R/teoLX
GE0b2y2jpG3u5u5L4ClnAqiGLR0vYS6tJK0cp0PfEqFRoBGGoEzFuBbghd2ERf6X
bJZxvU8ea82yIxyY/ick7bq3oTd9hiybD4PKFuKRkmISXXBp0aUrm06fj5m9J/gk
FVDRFKWWfjQ2XUhNuw7DJWeDEtapJ1qgGgfcnLUpEHx7gn/lzC+bW2L0qpu9dyU5
EZz3jg2FwvLYUbP839PNGJyLWig/QXwCxegVJsNqZqkTGv3tEI+Qjy1RqtJY0+pT
B2nVQg12kpywo0wmEQfaUyvk3JcHbCV7doGqF2hkkkWY57UtKjc/32gH58Wbj5Ou
sGSvn0L96q+1H5gU8gXaoptTNPzExX4FK3F1bUKKIOGdInmHJseKUXk21Ir8AYfL
gqz7XW0DeDTd903VcEf0qxmF6Azc24kPOkjnCVAsM2EeSQaLRmh6AyLadq7bIeEF
ifmHq4qC13mL0XfcqktV+hKwlLLGAHHn2I7AQkTGzdqnj/o4Mh7xnEv+XUk44qc1
s8ONIZj9PmmehRqg6yv6tmB9Sqqt1yFHdF7XcWIv/O4CA7+UdseHh25mYFVN529S
ndyWrg8EJWAJRtei4grPPWEne2A2pL0LA42Teins8zLyIP1fDGBvofWvFJ4N1QJQ
5nx2gn1XQW9rhN7Vy8WRsttzfu+c7TK9JqO+rBGNvR+iCyn5EI8/HaEeV3szgOmD
hGJC3c2/EWCE16K4fcr7fL6ufBoEMYMnBHVds4gO6NfoL+Coe10lU05v+MAEBy8a
OZIDEQU1Og7oCqWfxuc3wb4YXtzV/xZDUqBUX/xYdIMZe01bnJp/j9I4jwlMVnPP
fPjuR/sDyA6Me0UlX+nyt9OduRuik4Ep+UwjeLEVzVujvLKcfT3EuOu1cJsNuPig
hInfG+2FwVmDHiFYpxLjJ0C9NTebM6o7BsHFnhr/trvnYdq7xW6mkl7qrToQ4LZN
C4IN9XEMiqBJqNnz3TPJypOZdQKi/m9QccMGSLQbFKLfhHaQGceXXYA2p/EJT7vl
QPGiFNGE3gyHZlgGba0dRL8qw7GeTo73FXneFqepuWbLpVxX1ldsU3tmqhPOFLN7
L3JB7Uwu+tgVAn0iBc8KD1YClxszVrk5/1TQXwMgy3PPbFl1EM2rX5nHn+YTw8xt
Unn0J2D7F5Y67K+Ls5LSD4aZMiZt5pALlLvfp4NgvH870d6y5R4g12m7n6+cig03
oEeNezdTVeu5lpq/VuWq/dqjuW33S27UXZetQ3qSwq3Z91hcGhGCx8xVZzybtrgg
5t2CDqHqo2AEpPi37PM7pPSwuAXi6mSGCEVB/N0qNkmJ0/oq+YLb0C9JGrDQ/pT1
8eAKlkTB+kUi+6KBu8ALNRNQcobKuKs4AAn1Ve6uccg+7NKKNT/+skOGUIq7HP0+
Qw5fh50605XKJ73TciAcf5PAk0/1Yz5TxLmX/tqM0/RuHK7ct7x6H4QjN0X4d5A0
kXtzjx2AX1lwBlDXhtfuQLb+aavplND7K68gPX7w1ivj2ZV8v/dYIiLgOkkmRFtr
CrlXuvDnYWpCSzuC7XLnEcD+6y1/VdFbcVOJIdZyc2ZhPen7NX9cAdkg02FUU3ck
6c0YcuCik0hGHy9ejCR2Skl34+mkR2U/bMm6kzKrN/0Do+4PwzgHlysOl363n7Jj
B9odK5i0hCdhEgNDCOdqUQdGrNeF8qSPOixrYiaba8MZo/egaEe5o8NuUpjUAyQd
KQ7bnF9Qy/h9mokGir2gSO4QV7aPFg91Rt/b7ZMLFAzgmjHah3sszK71V8SXGu8E
EifpBhOUu57FZ+BV8Kbv/sWufchxgS7yq65oSUTV8LEKGSJKbOAZhNOUcVyTVbXi
xSh8G7AQms0HApE4vSy9MEACSzISDAZtGcWwiNRL329wLWuV+GIsr7ptezMlVioz
RR7gUSyZqHLVyFRZoq9ISCmOCOgScx2QX852pgZ3nzCP8/Lc7iraIsw/DHA81BsY
U87bUDn0BI9hQp3JyYaYQgrc9hZsCfqTZKn7M2VO2hAZewSaEWMGZGld5qgQOdRm
3gJiBJzLcwgzqXP5pX5ij7TcSWCbtcbDTFuax95kB5gZSyNJHlwEyhYgiqP/ZUC3
lWOnyOAGMGwBtjKBMRuaw70htglTdUetZNFayyFDs8U3xjZwLZpi7gNcy+teBIZJ
8bqeVKOwxeX1LvDge3KdeQH+8SslLorCGegltA8CtWtKNMhRt49vUCCXAdB/IxNW
tmDXyI5V/Ifs3JzeG1pNw/bfYVBSyGCqfh0OcAdhDIY9d19mB3QcNnG+X1rR37L7
TsLTrq2Po7GABjzMm/SCqZSEcB4dLPn+K/46//h1Ga2KeEML2bmlW+rSQaO/oJfW
p7zB7DlRTxZ5bLwdNmKAIyKGTVPNK+RLsX1+00A5eaUoptzMUN5UHOVM9Lp0kr7m
s6/FswdF/2K6UWGoDK1KxOrScj35T8CBaDBl4lUWbd3GvUyZuU+uHNd4wcu/B/M9
d/ib/wFDmO5m4zJzCCpoKrzx+ZfkvoffECV4Sc/j7ZycDcCkhhCPcczOqbYB0cu1
ckGmG/IfuVjiHB/uOdsEiEaW41V453e78+oTfQTg5zByMIQM/9sE50oj3RcS4wo3
N1+ngO5r4DBFT0t/aZXSQqA+qB8FvxX/GSde/K7wHfjHyY013qEjFYjSyON5vR7c
D3gvG19N4e6B79YoPIkG0b8snUumXumxPItBGVRbEp/28Ai+iqu+Q4bB7jvLpqBB
/4JFRBA4/3v/NX2aFpjGwKnM5VzjI2TSfTaQwNT8LekjWX2+YBI1i/rFEsUOAE6l
4uS/kjUnb7Br2ZzRmXLPIHTWk0o6XTnPhlHVDzJBMjBT8wWm0KxZ5Nf3zIvpepJ/
Oza6pQ6U4PliY0dewkBZ9cloYWuwKgPDnlwShmlZANqK7gmwiPgrEpADVmL7sFxs
sY7910hWcbQ5dLCnbS//3clcwiFqNPHUg/1u+QdvAzGSCBN4r7keXWoTZ1QjiS5c
WMDN60PBf5z194GMpOc/jzQ3mDvAFikbYZHcsyubr+FoOkNlE1L6rdhHPkGsUuIb
w3VJ3tn+08gZfzaMYqbFL0N/9u3VvbhSciZ7CPZ+lEuPu6yfHPbTfvZ6EGdD8JXG
o4Mln68z/NFnce92cW/oFPLGD6hoyqxdyCJ8sMKMKfaUMeSlE+Od05eGCTjjWZTr
oaJ5Yf4xsmhi+xKIBsO0gC8f+ix6lzCcLJnaHQ1KKinOhWToGLmzMaL3ZcQqH1q6
ZmJpnxX8L7mCVDwx0uA1wXVaUVAyFeKbSRiPUR7EE/Iu4NMxGv6+OUdrrxRrus+U
CNanSrm3JEWuw2OuTeRfaj+6vwF9/7F7odQ6A3sKcgg5OttzXarPrc8yqHfnLljB
aGrr3DIJe68Gwz2gcnWZsLCrX1mLPXv3IwOaPCaNW95KmlRxzwO+BA+wFka6EiN7
e/3d9V+uRlArGf70mp4OVxnr9g4okJNzQMnrXK5064rLSZSCdZEh6aqItrcnus8R
OYa/Wq7L0RWOBDoV6u6LmtdGjKOMLVH5oKjFDV7tVDrP9pe3VNGMw9s5gqxyKWHD
9n1maYIQmB+bKFHPEU0s1KBT6N9badyI1QP2BSjrGiNYhRu+uqBSqPo9cUy+2QVv
/+wVHbEeP3HJme29SrgPmAkt6oFUndPJfrs6Vwg89poL5U8+H/Dbi6uSz069HdBg
3ApSn5yQBPxaCM6+fsTfr/xnVaCCDw1FhCjQRKUfeHponmfUnQsrlg5LjBcyn9gG
JTToQRCr5x7ISh2YHR6X+VTuj0HxVUwnzcVimEadjP+jpkgf6fwJOqdaTK5mN43c
CE+mkffJgyVroTbAou3voK/aouCZbKelszjzz2TODIb+dxoolp28pvEio+mQ85Mm
oU4FaWeCcIqMsUa4RnumPs4nSSv63/5pVYU6nZhsvQ4+jV3UK9IgQxhyQpZ3R7X1
nbTHmhb2Ezu5Z/u04gFVLKFRlnKqn9rZkSX6+vvuhvNKY+8B5YCuWB+C/J5B4sJT
Vo4PUacWl7HMjvinRqSlOcwzJNjTPwSRw7LpZA9bv45/MHR7+owwvpRazKnbU16K
7wMa63QT4lg9K51KeSY9tpVrQxyOlYLtswS13ji/SkJmvNQB2/zQ/iKEC67czSAf
jsylhEBq2c61rkVrTl5D7o1Ygglk2JebJjHEm6AjD/MkY52ZZH8hSRANbU0tHfPD
BNbk9zXZ4tHpaO5pnHz2qTPwAhnlYejx5RV8Ei2LcuEmFE01DrlAiWM+OpLRylC/
jzlwIn2fbJdcAACY2+rWqQWWjpYZnVc0ZfNHZEMtlOQp3mKfwgtZ8gMQq/yb2cdQ
yUeOWPLwEemlYLwFyWUHDlQpd2toOReCmGMUv1yvXhtLM3r3tfbZzDsz5ysdOTdi
5p3YwVlLfXGHUPtB7Roj1Ruyb83ItrZrKR0ARnNJbmubYpMaBE29Et4oiOOSC7nk
U2GKrK0xQFM2ysfuy9Fm1G7nDGqtuTF5cqTkEmh7HZhVoA0UAmfMzjxoDfR19LwW
h8uv697S0WkTD5jCJQ6tONwruVSn2AhyUbW/gY+CsED1Rh44eJzGQgFF+ESGckgN
3X3qXjXhR/GThO4edxY/wu7kIUZZsbO78Aa3mZw3ulnvg8/foLVXRN5MdGdv7EF3
cLIb3PXlcWs/koMA9A+i0BGiyEVQ06GDwyOijucqtBcy1lm4ya45/jeKT68iqJBA
43hj9ylRAz6tOKHsDYJm1DYqC37xK+YYMuxC55Wbf0WZRoZGvHW0b9lbDiQ84lWq
B5KyZeGbeK7qYoo10YG01PMcAlMkjxF1gi3app40DuKDAPKAoUgwWEM2XGYvU+FJ
wOFuU7xqyCXoijAMYUwf6VxarJnscua8r1xpi2eOTjvsuXnMNhDNjbc2J7jc3ltq
8ZSx+LBkl+lMRme83vv/zpgCaIuU504xCPKnQivvVMVDFCElFlF3I5jgy7hQnB6A
4IVdgH8YHxvzUrrAqSfF1cYSQnkjUD7gbHh/GJclj5r8d9C0NtyH05oe+ATn5C5Z
P55+1lMuTHR8nGdOlOwPbhMO0zreM5ZPQ4PeDqF0ExTC4uUV0QoWOKWtKg9nNMAJ
t3KKZxNstdnl16GCWyVR9qxfGV9WfPlzx1p6xptRPruvPk17aN2ebXyMAAzRcpc4
PlKOqcQlEgtC8DNwYE8kZFtjTy0gNPu8+jAG2C9X2Hva7lV7o+H6MCTyCAExDe1z
/WyZJensgC42blvtJJvBZwkS6dC91kI8muV/JhvAelSG6KB9sNX9WR/+X+Asmu7S
m/30r40doCwmuulBvXTHXFpujiahbWAugW5UAhxnnQ0B4P/OW6fY04+cCqS8LqrU
UMVVnX+AqxBsf9q6lGPlvgBfE9rZFsQYy127v00TywTGYrmM/rvSlhHVFDRfFljs
2k+65FINo1HYQw6OdDdJMW89VYkFnfHlwoxxCYjCpcHEegno/v5ai9PjG8KK/HRJ
HTOu/q4kwu9cuntiE3RrM2DhBxjOHlyCpv10b5tZ02VGU0xVN8sgAbTCEhSx+sQW
UMivEmiYFFuIDjyS9hIsRw+CvK/teMT7LaZ/hb+eDwcwYc57QafbdQpUWRBMQK4b
QBPHm2HH/PuOFeju3iyUI77IBhoz1hB2l1MZy80fl/MMs6Sag0fZGuHX+Boojnth
WgFA5eHB5solVwt462wPUCeapZ0xqULsAwUuAjTd5Kx1neX3W9u/YvtI4kvL9tbP
7yh/nLJsVDAsa3NCwItoEJtnVprDOPTxvoUJA2fwoAy7n8hGD9KIkkf836+Nc+XA
aOGR8qovHyFNd+kwMfX3RF5vhX4u97I27OYa7lHeHccyrMxx7rHMNvUPCP/bFzvC
2CK+Ee2QGdEt+zsxXxFflsUivCY2Rh103hp6DLQFRnwgviVicTeaUQWMjG3WUDx/
EJuSgOyTLzr3g0RKTnWhUz1lwjpx3Zo8PaGaFx7EiUeaV9nwPRG0rNUbwq2JPv0J
eOyLuCM7fcJ+ltsmbazICbrt3Fw5du0igQvwE/ichxB5FLlSM7NwnSExoeLOiVKM
EN342+3zO0m8/r4MJebLIaXNBAQw5Uxuz3q0AUUxcV3SBFkO02NTbXGi4s7jeI38
6JWTr94MpljD57btgJeTyQBK1Th14H1uNENHIkh876yNY3c+xc0PSvPn18wgAawc
gH0gJvUFhKvdo60Bn+0tNcrLvnR1BJ/D+YQGhcOUDti93WlhIjxFsrRSKr7w6ZZC
saxU9DRGuDrf/OZY0+Nc5mJfeoKwBpXarmiOACXLgS+jNxw+bQim8fVgDBklzcMC
tdItwxVXfMTOQj5N4DmhO8ttiv+r6D0fFXXNg9xqNAV1znazcJXcWJLAR7O5zoom
cvqWuuA8nInTQo7zJilojcV7LBm16rSsxFqOggwz8RX7X94La2dbYORF0gmochaZ
4V5re66mwXDv367jp2LMPHpqwxRYy0EKNdLxZikJOSOTp24jX3Wh8h1sQTuqxybN
ZZIBe0JtqelCp+Gx8mBj2CpvLrybCz1VEoIBonw1GgPEGk3kpxTzOrZ49+iOM3S4
EpqA12GjZBUhBZWLszFk0Kk+5IiU9Y+BdlvwL7PCB0PyXTRJbgHW1hXX2N/5OJbR
rXGY/KuWMw7ofyObErp8P2n96wsuTCeK5gPYELqAhIgaSqRwkCciI8LwLzpGMZPe
ZQx+ShBW/LZSDbhdxrhEXArG4TZmMpkxvSlIBkQQC5I5pIspTsIaiGlHjF3+VGDQ
X/YisbYNpV3aADxKT2XpOeY0Daw7AJOFIirJJq57e0iwKXcee1GM9hd3HN3T1zbv
CjxuvngI0wDj3eWhWYGQFBkVUKDz1AhcKN/hX/CGgOL4sB8piVLlWvpqdTiUj0jX
VDFA25lQfI7BuAZ3l8y9IxzFvJuNnSLEXGfZ48IBGpQ7Kq8vEGqSE3+9CKI7xQJ0
D2D5mpT8doJ9Vchs3+p969IYNcfpdUr49wuDmwWo4YO57O2F0leS9Juxt/IWY3bA
U+r/Ng96pLoHAheDz/0d9M5uVD4bMISUpBN6NkpjNEvZ3ryTtAXlsFODAw1TcbQk
wI6JVYYRUIFAVrV5F+CJ96QIWh5CdBQTQTy2FUU0sW3JaEoiVhFiyy5GgErr9WkO
+MEZ2AJFtBhKRRrs+XfzBqRPYYbuKWSgRBuN6FFqeHnPKD2mzm95w173/x8ddv9l
E5yLkUxjLTDeF02rCyEJRvbRKwMTELClt+5tGPl/NuABM7C7V/KRMXCneHQh42Gt
kGhcC/sCmip2sBnicejCcn677IjwIH0U+igrzAYfH83QfevR8mJ+Tb0PeFVO4eVg
iipthMdGWuczVjkhMA4Dt+XIockk30a55Dd4MB9iW0gN5SFI1YlhELcToMGODx0W
r1+l4VH9eTwJ7yMCj2l89Xe/tH8a+jAnZAkSwfHZgRP8gKGf3R/F1iZ+J6I9/pUi
EPdJROr1IYwLD36NLlVdk3/eEkDvXFNxxNUWCWWt4gleXFdjky9QvkvB54VxAzAI
Waf/CWwwQdhVdeSN2tH0In2uHSqYh2X25ylEu87Jfjxfcow1GTyMUxYHnl7tf/wY
XOPRlamz/Wo9VMZP1q0s85gv3AS4awY2R3m6Kl1YLWbYonYBsilJJqRaMqFgWQ6h
1UmrVjATSRcAvYUU73IjszbmOwSCZlFctRdyJG/njXmER79GkDBDK5qho/Z1Q8jl
FCPxwlW0ztdfpJJbXaDkEhVE3JZP3EbrLM6F4k8p5FczTiY0y3Xc5HQQVQXbcCIo
ai+7XP1o68xBMrmvkeihunIXkShL73pAfuBx/e2CTJlyrZEKghnMYlDs4kNwyGSu
yoeRKHKWxe6i54FDxlVgyAzLTwMJUXQFNgaTUbtLyPuIZ933BX1XoWGCtjRJZ1Z2
wEvA02tZSWSB7LlPZyjvTSxYzWr1sBUrlI8Z08BxBqOc/fUdtjyZeZG5DPcDEOXY
Fjn1YD1DULOBGgG4dioxGlGv/AJv86EiblB22xCiSIOod9YdAMTZnG3dkskHfbPr
3+d5eEoyghx7qKVa+L+H1eNvYkXYzNRTj0onCjdO53vQB3mUOCmJc9iyyjG9ozrS
2dU/dWHMZgmLtQ1OY0ZWMFr/wu/ozl2LzKW928nkEV+jZUlkWWwYH8EqJ9dUDfi6
5aLCetCR3VUKk8doY7ycUtl+/JJzx0nGG1MgCVixvn9IA1nwZt1bQZD7C7ZRDviK
Rlt7DcV8md2x8/8LP9WyTRR3BAWtItFrrnAE12w6WpGk0oFUgAw39o3sfcfobKuW
dEbxeG+sKCLOupmD+l0QIMdPBCAtHBeVzzl3i5n3V3GOcV6I5hA+cnDe4IRRSZJV
v84ZVmAMyUWW2r+J0MRtod3+BAbDes/9Lnl/lMFtC9Ir9VPlzKoPDXwN81OqCacX
q57QODTzG6S4HY3peipcDXNkNxoWU7JiDAAajp1q9B8sYKzYEL8HA3I1KkHPcCu+
yWNiU68jp4fAV8nkVx0rBKLz4ZqJAPvYkiuDp5gJxK2VYD1FkzxqmvwUy7FDBcOx
mZVXRdrZ2dvM6GJh55jcHJp9NjA34j/enrKCHBWlJojlqsxw4kJxJ1bBzY8LCloJ
sc+2cR2zdedvliPy29GPGPtRl+OzC0neGyHLztHUJIR4o3DuQBjAwREor5bp37Fq
lhig+bEy5mrvngejUe2KSRBeHs8cQr7wbAb5w76Opm45ULgE0NuPr62l3mek+6aR
rYhPi07Kp+uZz3wfHGQ73qUFPNRZCZjxZicl0GPsuG9/rHVCL+kzOwRYfU2UWX3H
gMdE/Zcb9LmqAfzh6Qqmhfk1laJ2i3ChzVLNLTq/UT2ny7cRl1r3rcm8lSQ7QWBa
kD4m1vl13WdOuoBU3DtlNOipU1LsJOGYx5owRIa6EIPQb7zQI1Ceh46DxEb319RZ
j8DgpwAnEKx1JRqU12jeKT/4TYwcFlMPIAVBEyxZlephe1RV812rv8PkHWkjsVDV
Sp4X7w325XFSVHdXOnGDh8aM50Rs5EtSPNzP7y2jsfydPIq0Yi4DTKN7/xE2K5Yj
skkHTdl2LXGuDI+Jf9yHq+WIEyi37I6asmFlRz6mgE423pVp+ggdjOiuj37Cwanf
pDZeTEfaOZ1fgtS3SshXN9Sc3eB+D4sH3lRl2N9YT3K2wG91hHpXT+PxZcqPC0lf
JRtN6SReWO+SDM+mQ05aF1cQrkjnkhoZo32VGVcEuuvqxOabSf63vCQ8YcztY+CV
ViJKneue4qBXu9FVT4mszk6WK9CdO/W453jhkMSf9OMaj+CgnIFzIigRy3ib+CH+
UjsnGC7MjRW5SZ/gqTGdXIwoPOpTqT/soIoUuzEN45/uyLb6sGuxMbvOvsmeEsVQ
RdAtZp0l7/HouVCe54srLHHd6iX2swtp62nq6vYQbYxniy41m2WptaIQ3PixOpBM
kqB7Qet09vVYslsGG1mIZc0SlxbU1/w35cy+WQhFMuQwEMDCbuJs8jR9a0ivrTco
ijYWwaL/h732KawD1cIs9z8yqeO87lEeMbTZD0M/etlPD5oHRsg0jZI6eiUVOOyt
0ugvQDU0/OnOLSSmTkWJLFdoYJt56YrYC8RUY3mwUZJOg4HchKDAgURVn1Vhkaby
tq+t2+APK6Z+RwEeSW8dyqx2ad/FI7hwzBAUG8o2um5g9kIGwGHue7ao/jT/Brbz
v1OasUmYOFDVP3fEpeHdlo7b7xz7wTK7WNKoazoEF7PjODSS8GEgx3gm+kMO4INi
gQ5Na8jDJobmC9FbNGp1Duimw8uFAQ5XnPu/vzKnl93Wv6mm3XMKHDUx+l4rQfgP
6YIbcBVbr+KGczaEQwZHTiBK/8ivx8VPUzcE0XDA9KPRcyqC+cIIT/TgbUROztwt
O/gxQh/VEcIodgwFq+0/Vrykx8jj3BflHzkRuiSo9Z65o0ryHifOz5XwGsd/xZsf
y3w001znxSTg3di5BSAxQuUduFbZqyueYfRnxdqXx856xsZS9AsNhQKztipYxUKN
zQA370Zq1ZBeckQ/7e2TpKSuqQ0saHOtc6m7gDKiL7RtFViM5Nskn01ia2cb7gxH
EqtLcYZ+jz+pu4KZBNq0UI4aGcQ6y/iJcTwZAmssiBtLq1E8wgZMk+5SUkscSrZn
16dp9o6LOdgP4G2/VmHNn/HpXnrM/yyxn1HthWOYj4FGaG3DvJSwtb8tqruHbLkd
kCYZtA5ppuHV/cuOfHxJiUCmSyl2vOiOwzcVTRihbSGQ7UFnfZTv59+SHJ9xi+eb
5rPfHJJHMoCrCpf5yMKOliPin4bFhkhBRbSuCKOwu36FzOEUBH5ixrueU4HrzFk4
J2HvqH1S8xdLVoriNImVFuASLWLUbB5OCzc8z0HjUEX0gagbOKCVOiORrHut7y1i
vNzx8JhxeEkCtZ6n7PTRi3taKabp0nJsca/D6tGaNzmlMATpW5EDDxsjUD3+GnWp
DYoLY+h1pmyT4J2CpVupWcm4vB5rCnD92LkqCfhmM6AuAj5LiNRHf61nddnv+X2P
NURQMnOOTK9CKarWrXqclWbY9L68gXe0WUDONneIewwzkbV4ssjYpXR45aR8JEDC
VUBec/918BD51OOxiDLKcodGYZbgTjqV5yRzzJN3zmd05+BJ1gnKzb60qAFjCP2P
H37FFaW4Qd4jDJFuMKM+8q33sqSGk7iWmfU69HcEUXapfT5gM4l9BW/v1nLcEAMX
NyvSbBdCNXv6454o+MzXAv0s7zvmhOqJsZeFiZvd0WAGGGtcDWospXf3XMgfNnBG
Lbuwtn6MBjdMaoG0Jd7rIvzEgpEN/G4M1zxS7IsMG2VlQbOdU3Py2j7KUaK0u57V
Pz+g3BFF0UkSK/i0at3hrYAYynEaHkoO31qRHQmjnlfMZPfH4qBwLMycWh/Ragns
OL9neHv4/Wuznc/PrfRdXFp+8DLAAgLaxJZPHxSKxO7B+GS26Fxe5csRN47vwVOs
P46TRM9oc0N0WevfUKaBp3ayyAYcKGaG74tnxzYNMfibfV6tnYC6fsp4KaZO7576
VQ7iKIMwE0NyJetKIhgm4Az0Mr3iOZW/r7/qTwJ+2uOZOV5sBzuDeE1qWFvrgjel
1KZJjTkYawFLcGawrkjjiaBfwh2v15EOsfoXCv3nf/w+Lg8ml06ps/d3j8HhbB+G
H5sqM0OVwULp1CLRWnbf8kWIYR7+bgeV+mGv4IaXMoGv6+N73SUV6s32y3iIEqOH
R718zplSN1EyMFAh5gDWuujOrpV8dYx37eTXxFrTXYC6xWNxUQ6sQ5nC1G8t17i4
L1rHYSZfEFZcUBp1KsLnY56oZt1uRTU/rQcX1NLYQq0495SbJV3WCYshR1tNPQeT
g9fUUMYUEba1M5WQNASnOyNLaruR72KIvXBkzEz77j5r4P1a6j9+3zcBZYhfFz3d
fvCYqRTEfnaT53DNWjtqCPPb0LLITLZ9zxBSy8a2B8e+j6J7WnChOc9TyjC6GBq0
cPU39V+FZ/GJleOKeDw95bMxJVn9VQHV8RCVUNARgRVgPRfUuKDVNwvrVFAXpUqE
h80uobH0iAvJ95PFNMcbjnelbu1fpQA5IqcvYj9UMSESl2Fh6pk2iureglLj8VMJ
k0UIUygJQUzcvmUoz/YO0V/P0OabwwB7KF1wUZtEEgq4jNolhQgxOnaTGJYWBg79
9rO6dyP/TGhgkcHQXdh+IJnnQK9uGtVyYMEq2ZRnRYcaKnws71h7uSibdzxl9q6O
uh0Vj0605wwjTqd/GLlhcOL6Kr4qNh8ambtek3nJetwTt6QlCHWcMcI6eXPEsVR/
AwuDzRfPN+NrOdwNmZZthRw6bsHP+OVnXEWrv951zxMppyZPrTeW6DPms7oeXdLS
eO80aYkXUzRKE2a7HRXQf1mp8phvsgElGhdka7+ktGdoOzg9eXNZvQLHo9ZdVNeC
EAMIELboB6zG8WmZgv1R6jP8CVqnhaiBizjmDS7Rje6TqsSc5WfuS8ak86aNLQ+i
jUoviLxawJj6HGddIkWXOUj2upBN+ecpkgJH+vZg5siEUztT51pdwtvjKYjhs3Zp
PDz6fem3H3teojbdaydkQnUYwkYODs/62TYWMyDZuIjUGHWNWk3Hunexkax0/+8/
CitR5e0ueDN0T4WLq4UIlAUsrbfY6GtNNhWwt2GftazOLZWtRqELVRy4JyVSx5sa
0z7IS8cBA/pVKpxcAtk8otLguX/MVUJlEhOBhI2WJoO22hNWLEjH84rr0PkNb5U4
R1jObHsN/vbAsDeAYlptZ43vuDdDTFxanOlOMypGj3dO9x4o/jXI8WpBY5B0FnkF
FPbEIbcl1cvuFHEYoDI/ci99FzvEfbvhwvUN7CTc3zjW8DDWTdHaHSpBBJ9tQhYi
aTuYQKeSbAe2GQb18YaF5qDrCManIEg1b5FaO/dCMpywbJpn272eTdQJ55mvv8BN
HanRW9nNBhgs7gwmV5By0vUEKvSs75umOjjK0SDOdHEdtKZ7wdfypw3208NQldxo
Zj1KqILrTIxjmlU96YIqnOJMYXuRYJUQSKhC1BaZS9n+OjyCbDfetzbCk1ekoIwi
4wuExi9KCN78QUldg8u1iwe9Qqh0qA4CsC+qDMGZ0+fOsmfK7DYOLvqtnfg7YwjJ
ocMzQDbYoFvq9pCJoWAljj3BTRoR1UePqGkeoy3F1MhpI9hV3L6TwV6wmdfhlTZY
MnmlDBp3MiVvamk0TBdRFg5fTOzUJBhStfZhat+oWboDrQ9hP2IhoFwvp41uY4dJ
DAoIQly+WmZa5w1kg8BBGgM17dlxgg5MIHW/Aw6FP9TNth3bcjh+LT/SO9a/yIRe
Yl3ZshkVHq2hsQK13HIO5YFY6gkVzQYzRBbxku3F3PH7WGnXCieI9sUxTVJADjff
NxmgPUajEe0U2nhqEo5Duxv0TzKHodl/oTX8IVq1uYRLpvlvEsT6RhPAbd1MNFht
Ch9gT66uaHnIRyptCXemTozlqhk/p2fMjCTaO8BZLIi7rO85E+NnRKT3o7ShCoZq
U2tTdzgKJN8lBz8btypbm/0MFkdiUd4PIkoEcHEDl/ioKaKEkYqAdJx2tuPtK8IF
6tk3HhWigh5j4sObGzy6AAp8s94ComJne2qUebALp7zpGs2R7qyBF1UqfkEc7svT
zyxu4QdZUDupenPb3f3uy8x2eCL+AUeGYv9IUdzfVSUKGqwU5spG8DlmpqkHCZRj
+3uvynjB+n1gZq/bc/gt8ulzAwBw60xhj6UYIRpZzXBe1Zd5uIkc1d2ecYjmKtpN
wIYC+t1tmRi7GDKnT2JSM0IhVc87UC3jX2GlmynG3nF9nX941zvYVZy7kFWkBnDP
3bWPua+tArIt++EU7U6i8Id4+k8nF6KMgjIg+l4ak4qW45Yav082jZCJXLit1Ipz
OBUu8+KrUPg2JmHQpOI2HBttFrhq6j82bqaynJBCMrQN4sMVeBqIO4IIy2uazwsE
3BuQzMpWQhUyQriCddB1tu6uAskdlHBj8Tx2UvpXEDfGjF6M/q1FyIfhQm2WlBtX
qIR7ZrQEjJGe4cU9vgXeu3FicTmWcDE7BYoqAMg0NnYx7wqcHy3FcKu0ac6u5pI1
WZbeO0Lq9slyZ/UlZxOGLDJgfKKcP1WNPPglFZuHt7JfmJGyxv5mBf6isXXhrRsZ
OHkuSr3SyMQq+LoXWiZ1mn8RJb2RrE7Lt+63FEdRHbT9KD7mq69dtYiN1nSTXoyl
bucLZm/26PaFrKbJN6Qy8GyKDlHajeTr8vQjRtof0k47U1CVYmZSBoh9h56eXrd3
2mTLEb52XlO01iI+cp5qlvKEXK4zGzCdiSHHiHkK4/UAFkSo4rEFbZiGFVvN1MKG
u0lv1Kxnnyb3ZYw8obhgjgSU35PGHXCrTxz09L0PhIOapUxM8xP7lbBld3eA3GHA
LjGfCELZCBNaWxSCa8ARTyWYufgTvm7Y1WY89qj6NpGK0+Op7qV11t+b3pDu7u7l
wgwrtuxKQPnpp+NbzF2qNyy21WwScU59pbFrk6O1p1i8PY3OAcrp2l/Hq6Tm3S4K
z0ZRoyGW89yxQ8g4HFwpBWToIWnFq9ZGaodoMy7YX0LzMKrAQQ/8Xah3r12jxlcG
O06K5adjpP2ip2LRUxtVR/8UWFQ/sEV4wFik+3kGcVGxfjvl/XecuXnFoG6OZ7zG
6yXl2kwK7hIniDRA9c26aPrhzwWr9DFzUxfyBlpXUwoGBApc3Pr5pO8in2Qg2ev7
+HZZlhOiQsHTmHUYIUg2HxSFmShqK1OHORx0fpER/Zg6nW9Tb0rt+htgiYLgHmCx
WHDSnW+tn5PdFqtRbMkbdbZp5ic0dBnylRU82r17CFswOSFlRcMsPtrpk8Wk372w
umCGG8A0MzaB6q6zg5+1fXeFyOexKgBaOBdA9w7pBSNREEZD32nSSxHjEsoz8htg
gPdDQ3jhPltYHN05rVrvFdx4vKVAiSFop63lD3APhkSXebaU4Qj7UiReYCdwM5aT
57ng+IqV1MTfimd4rH8599hQuj8xOp/z50w/CF29dUw4vAxeb1VieG88EaYlk5JZ
pL26BJ8YEZ7W5LnkzbeI+PUDJSw870LOAA0z6WThErtPzTSStpcfMxymQuw0rcbw
jX5jE1Z5j1d4VmAPvI7PEkbOjtBnIDmva9H+T051coJtUHCz0Cus2R7/qpKbiwUU
CTybWKvsus14/CjsDMcR4dXay2mfdvE+vOm+ZtP34ZuJENmV0Jpln0Zgs3q4ob6E
a2qvrL5L+shl7mzTmTnC0vQrxYucJynrzE6lfRNkll1RGQZDbodOaMiW45Mxa2Y5
7V9QSqgdS05bOaEGmYAOA4zw+tr89OO/Bc4tO2Ecism72J0K/YSgF0ikYNrUIdE7
tKndPChIs+NF1G+UObN5vqSxn22cHuTx4W39IvnmhDPq/TLowy5eLqcH5jLkpVbI
42UmO1VXSewA2bYqYIPeRICnF4iFt5StHUC9FgprLh6ihgrzc/V4NHMixHYs5xq6
ttcDjkCCgFS8SxTkiTQr4B9a5R+8axyTmX0/yMd3MJh9nXS+RI8gMnUVeZ/8WeBi
pxzQhR8iG0NhA7ZeOOneUfIZeSmb34OOQEg1vNf32fKDIYa6J83eCtnhnLhXisUW
tiiHjAnkbg6spOSQrvSCotIf9qsSs8ts3jUiKDdtDwjsDbCOZAEWtfFCXAsG3aoM
EXV6pXp55/KRPLLCdEI/2NgKdxz79AbQxErylz/f1XdHSGUeOPBztQMg3rfcsPQD
GhtbRaeio7iveLOhvao4Jv6SDpP8FTW9wfx7F8rQ6s11y6yvGedhn9TWLwuxhg2w
0Hto2UrrXu5MyuaNrcu4zUJ0YpY0IVCLvCIEU+DLm5nPI0Sd+zqftEmmQ0Bcd8Ut
kbo913xmORfwXAvtdklf9zvHHETi2dHYR0Ymy2zEptLx49ocZRqPb7tFOnPJM6Gx
rTqQYlHiHJY/Dwx6CHBMc1cln+NlujG4SJfWoT2F7z0XgIFQ3FOLsFMbfJlv+C1g
eeRt8W9I1rlyY8ErUUQihZA3ysaj5bE80oRNFKvuh7Ecma7IbJ0J2zYg0moj9vHu
HBZwWKil5S4XtpNKimArbN7E14zU8uZjt9UBWkR5HSnpsUWAeCvwBc5pPvugkVur
N0DnGqtG6uTrGXO+vPPVvSbi4LIonk1Qp8OiM0NfeLE7gYNX2OYNh10cmA2eJvpe
tEoesWeNxNvIBQEsx8LXxuUkpuCKOs44FcdufpOdEpvGUzAk5SApoYtHEPnDxQvb
ZiPgiQBj9uLCR2CRuIGCjd2GFZjXiB+1iLzuE8ad3I2Gv6hJE4xAtnFzSnYhfj/u
qxx87DunCpoDGi6SNHnZ6HhVuDMQRJZcWr3D3dMxUZMEHK1CZAlUqFoborVFYsKb
u02Ts3B8Wo9GehVCd/5lTNfL9gT2MAJG4xDPOW6nNaYLECYQbHLFTDh9wTTqk785
nP6yhgZFztj1U8GeO1P+ZRJkZwb5qBVEbnJbFKHLmPOxjoAWStbngAWVoF2q7s7X
F1FqCuLFExVdflqsTMj4j1tO76Vp2/KkFZB8NH+b58UyhD0Ft8+N1RjbMSrXHhcc
9xVOax6OH08BmFQi+cRT67ce29YplMzY35jid6eoLbyUIZOZOUfSUnLjx6kHWiMj
hfYrs3OnhodtXWs1SLvSQUHzZ19/3dlF9/hG5mRjcDwFacZNqW90Q/tuHMjfM8XE
Jsrp/mWT24MmFlc9/sEIoC7esm19VXr+JaFc7AjEwxaZAgjkGlHCWy+MTFt/KKh8
3yVC7bQQ0Ucd7Quo0KYjOAgl32R9RZt7vDZz8DOZ2WQjfpjlMWWTq4LSa7G0XJ22
iBRRJm4hBpqXBgXxgw2voBi4H4MuY6yCGgvWFVMJ6TCUeedvPuistnImtgX6Cz5d
SoTebr18P5BHbCR7q8CC5rAHq8zIFn0u3Dwu1W43kmvRqoneXGbCW65CDV+BNgT+
BAeA7kYDSnpf8o27iTHR+q6KL/Fyl5hL8P9sws6elHONKvYruttxoeKm9rfdGK3B
wFYKVZpS+70yYOm5oIZqUepOT9T8boDvMji2gfJfc89X9EL9jR3VmZZJkV53u27S
6a0qJi3dRIcZ//GplJzHgh0lXTWvjSmhWPr/Ids5uFJ4hWKkBLkzX4DtHPuhF+VZ
OL5fF4tMmWJy8woW3c7Cz3vNgP9YJ4zTY6lOFh9eFuyrKsBKSILLMpPmFvZAc//S
s+W2t9BRsGPc9208kCrc6kO13gzq6k8hjX9E7MgGmLMbJzsbreFUX1UWez5E/L2W
edU6Opdj7cGtUD1aKerpivtJ2Q//f9Zxy3OOSOUSVp+Wi9RtgDhuvvwOxTzx7sVz
U1yKC5TFPXGML6Lq0UCVwDlLx2XUygyH19mA6qvpAI4JRVnepzMfjes5fps/EwQ9
nbq3KUgJY/Orp4wWbWHVqZmGmLSF4yU0fQsmod9igvnIHPJC1mi6yuTHQAGJG9cq
Du/8keJfwUHLvWZEJi2f1c8ZadKYWodWoO0j0l+xpye7XVPYdFCNNktn1TSRXJR0
iIGwoxwWG0bgFd1JDgdKwpQHUfDqwDuKg9qr5G//ly6DiWkRJQciB9S+zAp+Hr7R
MHJfu1a/cVRpbxQQ/hqiY79rQkzqGgvOt9eI/YXIdUiHPXxEjcr3S+ykgLTtcEFI
c5+8kr8iLCwkaR92vgJ+f4+9eKxVte8ut3yZnXTd6sPbcVQ2UtlNwzil1NPBwuae
4sCnscBqc7M8bIxKH0x57kGB2WoXVdvKo0MWCsk2V0d8cf1W1lY2dQwXJEQMyXkz
ATmpayldyNFDMRG9WjVGDAVlogB/LbVz7Mo9LmUZ4Iw0bh8+lUurHAAP7McDj0Dc
+4je+6Yj5Ak02pGLqlaav65TsBbbZMsLKKv3KI1CtUR/jTPXtZOSE2K6zV+55Csj
hnpHFIAYTyWdTHZUMlmD4fmq1huNCb2wVTy1O8uhLvlxuJzIDDzxP7xFNRMIIbcE
oP8vhcweVLna4S9r92D8V546AEgBZz3Ob8Lf6wMGV0KaJqmGW7WZLK1jjbDtsfbV
dbcIlfPp4eM6LWS7lcjB51HVKNWB/YTHjhLwkk3mMp4y+8S46icZ5Ku8HtlZHTD8
0pBVFBvWOELMFHcrtoMYJ0YUP+Hkiqw0m4NhEQ/zMisuv2TFkW/XbgtBfGmwHQ8I
meBRTQlFft3Kk3BckG8KNxBqrIq2+PuCSxizuetJGQenAgKZJNJsw5QTRzhTly3h
kJVBIglGDlAU+jaRxvhvA9AJelZagzjB0S5UwokDykQDdDUZQeIz9MsjqZuMAoGQ
XpJcYdzHSlHDPEpn7RZ9/IUbM7imY42q2oRG8KRUr+VqLoeleNj+//OYkaFDQsng
7GQN2vuoFjZrNWV6l/12UMKZG5QhE5zv7TuBY+Kz1+px9YxosNiyvGYvK9bCqZyI
T1J621qHV6tijDsOtg0jtGNcETt0d4N8INkNKtlgc7t7yihfneaixH20ViLJr4It
T6VN2Xo9OB99CElbJYe8Ued30ZiFUDKD7l3aqiMLXMGseq3qdnb3i/fyYJNItenN
8n5tisHyxiTxrbPh4I9BgT0nsOQCfpyyVErH21lI+z+p3gVL2ZnnT7QQLMuRV6kJ
pV0yJA50Mi7M1Hk+YOs4eXenwzWL8zvvIlef5hgsYa2mFgP6MU+85Tffs4VrUQGP
gzLkQhDPQFpQrBD6BFG3BUhTJF+/ucuGtDaUBg/9sfBgJmdHm6vDD1ZeWaAwLwa+
xztUdmes620ykzsazyc/8CYXfJXAuccmzzfJOXCyO7ZD2dG3xW/WAk/0jVI7QJrO
rNfyRpBAABCd6nNhmZeRcAtt6DGantc+LZ0gK2niKUyvXzc6e1DJ1YP8GRQRJzC1
xOF/FW95SgqKHU2GvOkEUmQeNX1g2OCFhDa20CK8ukovfR12BF0bKEpLLLG7Hm8T
UPwpjKMRMgoTF7nYLj1ZTYzmcDbHMD6kjxypa/7divx1+yh+BpKWc9VhDDQMnJ2V
mXfN6yJVAvBslxneLg+x89zQbks7PEDu1f4qNs8D/fhlgYnIEvsRCKptc+tpewGk
TRTgrg9qdTqThwdYs2MXLzxLGbYPXIUrpWHsa3eqUkQYDHb5x6NoPLiNz4fHteTa
bPg2sd7CSAIlrQqBqdfNPqCmvxTBNTXVvpEaVoiTi/8aSm2Z20dWPYLwTmyEdbAV
S/3vLRCZ1YwOv5szAvGDTcrjboMc66ahmECZZ0H+JWK52sbCUMzkVWqfhZ2GVXFf
Elxt1S1SihZgpFMnb+osKKSfOq3Ude+Y9DkSBJJtO066vwLtqq7qJVyG/ucVICys
zC0xOGwtvtiPnYySxp51F9JE6JyvxA7M5pkW7vX3JO8DMFHBtcVWmDFr4AAz4Jkf
THKjYU9wEjPebdaTJ1BXOl/2WudVDGdaUGqGklju8I2XCpOCtvN4ut50+VntUid/
cwwP7J2pj9lP7Fp6YGy8dSV5SKfMWYwj+aMkHjfJOB92HuS7u+bBlsvAllIz+tXK
fRGevvYgTZBRQoFn39wdCyRQ84zYTO1Hhznk1t203gmrc8ci3SNTFdboRgtCnJty
woCvHEX2TuJ/IXNNEX7mNkFqhYjkHTzbK72ze4qVKKZcccPhyX2kSr2rcKoCefLa
4gEIUrhnnVW6r19edBHSr4+EFPy+col+f7IKKQf+nXftM64/51H/TXHniSiSXwPr
JgQiIUxa5xq90Ln0As3lqrf3MFj5I2yU6aMWrjEFASaAk0031h22iAZT1zI22EYg
ApldU0sRaGAYbfDyHPlDlHdfOMWrLylIojiIStGWX3TuZXzq4MmWVO/N5sFH038X
upihzmvomsCd5sfG6XUDuvQEXYiZIb/kYPnQd1+GKumMwbj0xHZ+5S8oYOKryBya
clw/HodBDbEAEBIA0kSPAjHTur2E8pmGBOVn349iBgRHYBGsvBjGj/xHR5E3SobJ
aCwnhIUHJ+l0zc14TwBA23UyJWecSrB6lLRBrkEZjv4bSZ6LzLDohCCuYdUDoWnZ
1+ZDILJxaE8uTA5YHBN1wCufx4I8/9XXKESQPyNFHGcsBkLz6Aqns8cpkjDh0oAH
rJNYWK5NEkGRWBP6y7122eju1CV8a0BTi8ytFoAjcVGiSdTvR5cvYyufoUu7gQUb
xgwYWaCLtkCFbby0uqsA6wwfZoMZUTkh/U5LxSU5bnCUBtCTQYk7Mkj9heoO5jQY
ItLs0QLIt8lPKUQZe6pTToIfHevShAoaySDgV7xLU1gef/PhLe4zyPQ3TH2PL+Lc
pOPqL52rxqC9usrgDZHxrneH0i0ZpKt3d4Z75V7A8IqLsGLYH6WzceZE/r11dr3I
SP06W60g4wsSizsO9AwbnMzCeU0xim1ZGoGEVryf8NZyk2sCooEGR1eYlAAk3J2Q
g1V0JT1mCgQaCqKmjHia5Zoz0dFWZ3Uffe871eA2/b8vSjg/3chsx78A6C4m9dkr
RlZNi35pxTyXB4ZedfC1X9mcPWS4mWHwq1ztH6Mn2oG9YOZU2iDJfBJh26kyq2zz
EX1wmFt3u86hNcgjEK5NVpQqiyq2dQTyK/xF4lEDaB2La6VAI3j3eFHiUqJmZDkK
JdpY3VzXmTr7dyacKzJhPxupXTqyzab5k9ekgGwqMEi1PxTHsuBxCYnkNSfeQ1l1
Oauqw6S5HQzTthae1usCrYl+McZtS8K8Jnf3oya2O+jrteaM3y0/INym72I2G21O
L1DqroXRO9b5u1XQAWcMnmUSuuQJFYp68lnHCzAll6T/vSgbpBzePS9m9bhCqGM8
OW4SH0WCtU79Fo9AVE1OQwTWRCuOlyS8WoxgwMByVBHfelT+TrVVGMHdr9oDw3X6
Ub7CknfH9DOobIe8BFfjiSI/Y5Io2dYOS3TYiWoLSclH/nPkFkjP5ztB8Dn/lRpg
K7f9FgucT4GSU0WEmSs8uDObKPagBuD6zi/RsgE3oU3AQ9tFsV3aqh6h3JWCXcEH
Ez0L/Q2bqmXlBi6JGfU4VpgCaUkEiIbXXT/KsnQ1QtTwZRgYM+x7uMQ0LK1yKJCC
JhcWpIHcJNF0hJs3msqDihm3BMIXsAyeKKuZ8nbSI1JkDKBlIzQB2SGEC/bk4TTI
2Tq1qJIWOWYkaZpp6nF+X79x1TY01i9lFQwotnc3HVikJRth6bLYZx8Uf3+lWEt9
uUCm4XsxDOBBzTnv7MRtqhsNaRP7PMIxlrzVdxcSO+3QGzpWV8C19DFEAMXFioYh
FK3dYIpcJ6LMu+yOspHkTL/GKQumh5O5bWmJHPKrepl5yN1U9hg/G+x8XyBSEelY
blxMo4RexkojDXJvTqwedA8l8tddmZlia4/5mRZTZ/BSHo/Aqcan8+lgTrQ2JS0B
eqbB8qZPan7zxhJfVjclStYZ5JxmguoY9kmCzNdAV7Aw2ET8iwnfj4wyF+xHxeVY
412M+FNoRdhUZ34tIY/6ctfg7HxdPEJfgHJ9rt2jwLN/QX+4ssQILfWeIHfD5Qu2
e3VdIy+29/TZPyeo895Oc+M3969hT9NB9hs7K7lxtfvD+waFHAFFZ8+T/WI/j0DZ
OmucCjrVHFwkWtRnLQzvOJXYagemiOM7DBtZEk50R7+ggbTiV5hrgzd+DdByg9T9
8wn3UiDqe/A2du+XmlJsBrtuyN3xirxfpI0u2y8woYsIg18Rkfam72Y8CQmsouay
AT871k/3Dgwz9twidT1qGrxJH/Ev6ovLHvKMVwWDUcXRtQbErJwoNGPISKiH8Bfg
RLsqQkpxNuxTpyKMyfpT/HmiJELVrBcppn9coTFHqcF9ZgznulfjWwVOJvNsKbua
H9O+MG2CqkdgUJzOoraaZnghkmNhqY3v+s4lTwQG25nzvTirQDPLjTsmZAz7hZDk
owVGxpnVB5HTdWgszBAd/OpGdW32334Auomfwj1CrmqAhZo19772mkojpLpVmO8h
wgiBhV9H2JXkYGhMvRU5KUKAZERiWMIUqb2WUW6Ehk3p8fJiaJQ/BvWda2+QjwxB
0+p/fKfaRumMYxtATeCICzldTJkS3zs7KcpYzaYr0aoyYFHpA3UftpuO3r6X30WW
zfOPKe560Oh1V7ckMhta2pdxueAnRWztCWDEXXAyFhOjFJQnO5MUafOrvEEX+f5b
slRio/2bYu0hJsC22Mfec5Dxgxk7Ls7Bc7rdUUv2zWsZDHULBykYaVNTxQZYmhLf
L2WR3xNgLvzc7GgZ22Orz4XgmdDo5cNKz61kEUs2WP70B5MRMAzL960DYQicr2yT
FLyxC7PwkmYU+simuBpMdogxr1tFj6+dwa54mHnNx3MO0Rk/9Ok3nPmpSvXOeYWk
WifnG3t75KYF/aL80yYHv1g9yfgKGjIyb25YOEvOMtLOI+d3ltHmFlyd6joyKQda
/mXg8WP20K223XxnX58kEE9FqXUKqF7W8bs2/p7+CXpqJGwBC1UqGId0Ip6IKgk+
A56M+BD7MePHrAgluhbR8AL5dULXCIHvse3n/lov+BEZk7LEERMO3Cb9ECowjtQ+
cT5ec9ONVaitAdVN/4DDTRo1Q5hZwp4ILkmp5FWcybnpMuI2Echpde+d7BTTPwWX
kwmWOrm+OuSPukM3Tfc3aYVDHDr0vPA2uqrKrfA0+L9L6BydDeGt6KigqxtW4rhq
KGCNMqBR+uU9bGxlgqzaKqm11WtIqhWsZyKF9pdGhE/Yb+Is4lJ1jB39nhj5SmYo
u5c3VOCs7MW7lQE84cpTOXGmhT7mokJfKvBtGZbcGevWHZ6muwz7jHRhWGreb9u7
2w2S5VgJXKlGA+//eFlE0bOyxq0N5uTNjT2eCV292UL9/HXEphBnxuSb4cd7oNkI
2Ux+M5cHUNDZShOCrfM8bvumfMb+dW8W6Hm+7+5ko8AKvSefwB7VK8VhMBd7zmRP
vOqIdqYViVfGAibxKz0Md+qN4n3Sln6jRFi4T4jzG8JedxtlCLfDrhpMyPtEtrno
bw3wJ+tQVTps2mGpYdsIIhDJbEabjwXl29GqLYD8pfT1dk9hlfEPvpfG5L1+73tn
GSDcgMpHuVlH3J0tBeXqKdqr7P22z3XdEhAcOijWyA8NBYNLNmVOUV4JMHodS8ax
EkUzHepNTQX/yAaUOtlKocWoyxTtSzEnq5gl89eDBuB6IyTuSZFC3enE+gKQfybA
+UQtMkaMgG63HMKiw5j9wvdze99bghm39excM84XESN0+eNmUNtGjqjCADWUbUbh
go6+qh10OmLM+R7TiCk2X68VUxi/gqKdWKE0h+ZNr13CpNVJmBoyhAOn/U9yYg60
3NvY2+XguMAc8Wvm0q7kLIgS2OUx1T0mbd11Z1dhsbsM3qhYY23iLx11KREHfKf8
dYsav2AwZG/c7rqFaSvPlH6IKFD20QpUNe/fn4k256V0tfR/CgMP3DqqCYXjNl5T
DbcWCUAmdAtrk7bsd+jtqXZ0xnFEVrx7fCa5FUAneRPTftM2ExMTNqhOUNPew8A7
D0Vg9jXLUDGEe5aV/4NuHdRQ0Ao7jhJmpBcMxkseIya8jBxGNniMHkE9Rd4B2gyf
0oTPFdoBODOgKP1y5lgL7qBjJ2x9xMkzJ2wN1uTyePUVrYMv+mB2CiQtC63K5pMA
IpiaAfnc1THD37tVbs/wXLqJb/Dte3RgLpBnh30BvWoch9OaD2kbHoHFMPNl1yYi
rc0UhqBnFcXYXPqivaCUkgD0/Bqr4vdQs9UxhoN5yy6FwbWvcLHH2d02oWiHIBsq
edX/r4fblEiJauyLgseliK5yrcmyJawRd85hQNUskREaubLfMj9lJy/LAAxFW3Fd
rvF5cC7xqKmS6KFDn0n3WHWmW7MatrbMi9x42BKR4gHiHXlnZ7mPpN7dDsuiZ3pd
J9VkMvEbdIYKaZU4nQNmOuc7S7H7y4A2junhWHH0YuBvVR0JII+JQuf+4TrgTUfb
Melks9HQEmMqUteTqBkUC8n+S6QENkrlHwAoUrwJGyyo3YyF6ujaqDVwtPm/Jp5h
yVsRcB+9mjJwbJxn6qpfNs2o6i30A2KoPNdL8jEplDUnW4/1aYTbnS6z0D7knXbC
mCD7no9LFwBQWdLElrW5828UDZsBHkU02LH9YL/EwM0oH2fuAeG/wn9fZrdqgOB9
zRY9SvF9G8EcFMxKKczHSDaUyAOPyDcS/xmOqP/hkL2671nGZtXTA7T7LfwuFrFR
NHJaz3b4CWn3XuVbIAPCF8QiS9SaoDAoRRgDsnbssWY7gYB7kXJOsRyartaK/GB6
oKjLoJnc75BQZgiiEvlvPwqAZrdxhKNULvSyGAZB0yLiv/X6dmLuiC8BdUoIlDXC
d2ZeBUwEFCy2zM/bygwCyUy8keDJqOPzgVFSYUF/8xdi/+xBWD5WypahyItkCKJ7
0DC4LfXx3J6ede6s+3l5cR4ihznkP4aru38kFj+yvvrY8S/1gtwJbZ90q7UTTaUo
vVrk+NU8n8ji0x7957Cz6eWYX36+sQH1NJJzjSmHanVRH4y92ci7SWLNazPshvhk
1nqt99HBTz1FEyprdXlx35XFFuSOeCVru0c7xgDC3hHlJIByjoJfN1igFHE3KWak
QohiyVdo0Sv0oFjRBX1KyqtgFOln+oai6WFSfiOeKoy7FDXQWRVjV1qyR8HlxnLs
hxZd5ja8Fe95nFDWbYwljrN2dGgojfLVla4E2IdN+gUhnfIriq7GSYm7o3vxi9y4
e4JmBmPIFWP1p4QQC7XaSLKtI+LRWKMADQwbtXhQXo/vgmfMWpDaeS9JYcHe1iZl
JidJ9IyRzxC8TxPbiojL6c92+MMApFsOUynWjB1+WKBVOKwQGqgHUX6oxASogZf1
vJBKDVDy2Ct6I966YKqZl8WbE56erlzmN8o9lGbCA3IrVqdx9uavC7xOMAbl2hnk
JY53kyHOqSTFKMxAn44NEYxXx83SOTeYwt1fj79sU5vXBWiP1WX3CUtGqq02+sIv
eV/kYZRM2mBC+DkLON6vn7p7kDSwEEKNMnm8YdLrtC9SpqV5vk0zRH/4eAeo5zWL
AOBB5FmgFK5J6SzaaF0tArawdOB2KTGAC56i+7XrzHWyBoY93KfdA+PHbAG2ATxz
6s5+/ytZECaAJ062dbRLRtqecYKJAiw0LQENJz567HnxGiCVq+um2XlDkqTo93uF
0D1/0Vn55hwl8IQhqeSlyjv2D19atCPvcRtkCjgTQwiJTPH+Edd3FF+WapFlPeT7
Fh/M5h3ivEXFXQ1ZYxLdtcWMgtYUZbAt29dO8UKhFfvBPYyvn/AsJSofuCP1BIkb
eaIYKSYr15OM069Dvft+sASFwDfICn4sEciAqDaPWKPcq8VNoHaMVhyEWAUmiygL
WltNe1lj5j6ZGGAuXPrbZ7cPK7P0kD13irKGx3Yuuu3QxZyaWrYkU1iQdRpUrKwc
A2SXLC17wBnVKPBTZ82yP9fBivpxkcqp0awNb6zoVHsrnhy3ROsSgZySA62zKIs8
Xr5CC8cqsAh9srxmf+ci0BMmjOfxhVayAFJ8yyxdDvZoU4hzj4yuVfAW+8vkdJow
bD+Sf2xD1/qty/zTQ4kyNeC31iM8LX/FCbxamEI1QY/ALDfUBBHt+SbV2k/v1y0m
AfaaEcIWwUi8WWXM2lji9CqrGfpZhXvAgzsXBkf5WrMVddMDy6bm+9FRneU3fmm8
ZjXa3AgQAlxkHqg22r01Q1lVrJs1fAuaWZzbIfv7AmGGdxDMBOEG/wozkiRp/myj
H5AkJ/wnqUxVRfUcdPklxtJyH6Q67+m8GItFEolfyYe3SeMBA4f1lbqK+ng8iMOd
4c4hgCTZytAPZ+QOPeCnMsrlhaA2/9Jpmsv1+HIKYqO4DP1aXWMKIjraneIqa7XR
cj1Vn8bjOfGW4yO8jmlRhsI2aSEmu4R0qz6hbjM5Sah7UEkjRjCuRRsL7uh57hH/
+rZvGNGi2YBLZN9piDV0r+ToxuKvsrD/0c+s9TJ3hgm648lT9toOfAPiPRfqFv+g
yJCBlXzY/C+OsAchvzNHZGhBCTwTpw5CVSRKTuXmmwZssuBscPmdeva8gKhzzxg+
lgDr9h6JAjoS0tEoXRpvMTW3EAqt6zOEMrzMkfaIzKdJ5RBH/XZEmfF1plbpbY4y
bb9QfQCrRjzRhxDCO+QumBJRdOnpUeoBg6GU0QBtwwD4NQbQ1xnVX+N1vyp2w+VY
/O/ey+BiD+e7i6XwJOXioSmRZ3J63lAxXiKFLz3vQjt304kJfeqa6maofOF6zMan
LDe3/p0eroO9Df9tcX7eOIXPxGyZDVEgPWHqd5kowh6RcjaaBYs9X3prKPjcUjFX
ALg8yePEJB2oeRJmL4Uwxonu0Px01JIoEyYrqijXvJTWC9ABb3c2PN4MqAZxwSPj
BQIaMpJKRrppoD0Ph4KssgtquPNbhDAu5L/ZRffmpvFz6XV1sUkeCCMPRVLTWIoy
zVnNTQmjWjfVrRxAr86prJ21Whjkr7CUF8EaVhZV18LDtMcA/2OKcmTvZu3geBW+
mOqnR0QR/9GdH7+pjpfmCtgrgjBq6nBjCnwBeXEwkpG2vBKzgMf6gd5KB9XWnD+Z
eLwExe354U8Rah/ohEA0EagJuoWHKrf9e+Pe8grSaDqwJszeUv4r36IJmZ0Oi7+s
ZoKJXcgg7s69bGI8TYboA+66hEAMbl/p4II+ny+R2uDrO60jS4l0Vb02nuArIgX8
Ye9C24VNQbEH+iMg8abKmJEpjfRiD/if/jHqOtgOrnaVtzTeCOd1csvpRFaUPICW
xz9rOCuguWSlHUuyQYkiI+S36vvHVR3IlI0zO/zeq8JlYQ0uSNAUbCb3j5Sbuz7s
OHW0qow4jmyXawsfBOohJLRq5D8ob68ctKM+kqNSa0Uy4WdAwv8mYtpoRMD+n0Eb
kyG45wx9UyK/LQXoN5ofZLG1JeETV1XWiWCakLBqvL7gnLnGOYDHZv+zo3T3ZF0Y
JVXCFmqS67NPlFWVG0ZLgwEGFnbXb5SyN85NzIIOquOLEvXolkZ5Q+F3yv84uaO2
i7P3jVnYzxJ9FFR+hBU9JJ/sEZ/H7Q42SXgVWnaut6hZf6bFeTvGEZQ2kjMBCZfl
Osb4AhgL+PAA7jMVn1Htg3J6X6d8Wap7vR/XbvRvk/PRSOivbXVF/JYV4JBfO5Vq
UsJD3DHp1rDUUfCiIFDtGTfnr0kXhSjsv5n5BM4ljI4X+/C5zztQ0kXdsTVvbNb8
8711e9cUjAl8LBWsKmexORFPEq+v9CZ9H0ii1yv02MHr6DYAG6WqhDm0U0CguOox
O2kbqCxS0utiGP6MinGu0LHEUQy5HF+qhHqo9vEzNxXewsBVi3UP9yBgn0xtiVba
9D1oolnvHbjM+jLTZQlzXYPCvEwKXDTRRgIccxVmtKOT3WvVV+QvLK8dEgtQZyBz
1JBTwXmX+CJl+ZH/CtRdF2kqoKsu4yqZaKgFhwkFZhZ469/HElVzrzvgTJW6Tlqx
lytqDRW8HQPbD5DH1aOEZ+/zeF54ByRtUkhQMt5nvFr5C3FfjCFjdZhY5m24jdKM
k1lw2Lc2PpE2rtThXEOLSVfsk7lX2mJjPmiWjawwqxOMeILh57wYkpgXRCpnU1pM
KJ9ii8m9cUELYVgig/UXvc8awnW53nCiBBNwAavoPKAkEydstXRqScmtHxmw0XUP
t2wCXjSx/s0dKSqL+f4qaQBwSwutNruUQwMP0UI7C5QZu2kH/Ww215NmTsr1ZxI1
F//H8HJKojuZuBmJGkDiV5z5RYMb/95lXx2W0Wgv082VJ67bTJ2/DQaZMvYz8Oes
SWGf1tJ7jbW9IhtNk5BDy900fKQPa4qkQFXPdSblDMCR1/aQxy32FTxDYgCcA+md
jN4S/KPXn7D1f7mTFLmV3a1tRMbBy8t47sBExcRPGuoN8gr5K82Bu5KCsItFDNye
/E64JZ+uwI4alzFbuA9qjWjvVdgtUKQpSnAm/08K+0Ou7r0hql6vqC1kSNolxr57
OGF3G6Sx/XhdYSiUwFSIDeBly5dF4UDJcQBiisqLXVBr0aqYl4+C4sxCy+qzfqGi
Req39O6zzRVoA9BsRfUCMp8HWSU3mK+AoD4MOMMRAihcSiBjqbXGWeKeKb+h/M1T
rRjXw6KQod2V4YC98Iel0Q94VpkX57rc+wd+SlGzPeH218vog3H/bcP27nzzW5f2
G/cBGlmf0Bc50WbOLvkObUPpoPF06uco+0/emdZFNdhdOI+6gJfezpMXpOiJvpbr
DVQSkitnztSjdyQBGPZ5caVR2r6B8ZC1738WrHYtrpV7xxlONLn3rF7lKp2eMlmX
8IwXoVKDgvqVCJV4pRIYYF8d8pW6C3HWI6jC8a/frW7iV6x9WSVE5b6xbbS2DzQs
qOkyTvt5LH3RYb9CCuSPZay30psHcq/AtHlJBbZGTPDyY3h2a9dJ/r7SAMHUo3t6
FxJSuNf3udg11Qi/RrQNIdYTKNBUzH6GhUZn05BSnwdyIa8fkQXIuDoeCh8yiGLA
nWXQqj2Hb0vgvUZfpjlFD4f/Ki+ROpZezzVyv/OpF2iFojI5XFGjtafO4wc9s3Ml
p3J90jUzrKj+xZu+R0JkKwt+QgYZ2BAzvvotIs5wxRJEjML/VEfZtX/jXs/gZ2pm
bKkvbw+Fh1ZEzc03IXEyjrPCO7zhmDaWhacIu2rZ9Z1UiJTI5QBzr+HPyAeCvi6x
6ONLvb/1UGstp5am1bosr81ItW8rlnl7iYjV3pz0h+R6oiayJPn3MJKrUenXIj42
58krjaOM8OEnAHcPIha9xGlx3muX5Ik0iDBYb/aXNPRUuY1W77ql6o+NpmBaP/W0
XpLsNmI8FcqzIxeza+tSxPoo1H7VbP9jz3jEh/zOwZdZcZTbURoITBsQfrtCEjdX
loH5Ae9zjhxD4fH4Bn4mlR3o7yVZujW+TZeNEwjdBP0Ujnmvo/lF1j32qBw2G+Gg
MM6rgZL46ww13cC4eIWAOmMkVyFqKneYIHXlD9Nxs4Lsz0Q+aG0VSTACQ2IR05S3
bzWpYUXKOAK2xlksG39yOH7m40goiVLvAVVP4TuseomE9RhVceOEqB2GO+z/3la2
CZ1hLO92L8jOsR2CwoeXib8ytzZAaUb3q8f+qK6z6elN6TPLcOUfLWrTGVshQ/eX
qOFRkwk0WqGOi0NVbOH0a8SXdHj55L2Rf/tIuULQo+uB9+NtHf9i7C49LlZ6qFv3
j/7UsZujeAzvjq/ncjFMri9FuIfHdMrj0/G+VPsAhslj6NzA99fI0vJFa3wwmmmc
O25XUQ8mbwsHbo3pDmOE2uj1PiWl8iTKRMH23JTwn0fDg3mwvz110rE8EBz4pVTu
OQZDx4bqt9bg7u5PwRRgY5KcaUGstyAR2m3AE5f4WTaCaQQpXrdfcl+bG1Alf3hH
i5BbBzcJEvWHA8WcNqzA3VKLWLvCAkXaGKW2v8O1GfrIrR0/1K0rKDqXZyZTQKzL
NrqPx6HXdvhWZNFBjSynbXACcBChXPrjbG1ir0+l7q2swXo6hopZOdslEZPwfclh
a4BWhBC8kNtvjExo5T5K1WPKJE0r0Rb0mKVtXRK/48g0Awxtj59AIRFWYQEadPpG
5411NAjqcb966ztLh/wyu1KM3qqFFoqiR++2M82TlSFyZkWuXom3g9k5Ct404HyW
BSPDEMa5avx3zEGANqA/dfdJBe9QMcUxGSqAoBaQB6hkEhb2DblW2cBhdJsI9Fwg
F0BxZnh2T8vAv7XxWKqRUS3/H/aXiuHPohNC5qwH6tG1g77w5yyARy86XmXG80Nr
Tzv5tk60uxqdFFjoRpC5ymdTsgTpRgyVovOOfBIpX7Tw39xZ7hxXk6m70tE+56c/
xGN0YCHa4LTLh/hsj3RJD+nhye7qKbpQUkpwxy/zG2MilzyzwFhKaXNpCAT48N2E
T8P7+FGLMGNdqIJK2moc/ogw31cDAlSi4QnegI4SkjFJtGSqj1zSfZ7wfpuNjxPo
ssJn36cBi3vCvxPssUgnezCeC2IahjPZk3VJd6Jegc9NmFgSZq0rVzOUjdqDF8DE
OR5xhxrfxTFAwhd0+Cp67z/oYmfkWjIWgYKi9QYvAK5QbqeC4fDiGfU9zXlajORG
ApyRIcxQkbR2LIOfpQNRm200Ylhp96rGBsgXH0qMXgVJLN8mouCCzeZkHHyiVqyz
Os2b46LDzxr7/vM2zrTJPb0OcQMUP24GNP72CfrxBzrg67uihurCpNd992dvWt+5
id0IU29lUyA0W8lFWv8HJ/7ONsvS+dZ3IAD+2qVenlCZeI6/WaxgUKG9irnmZ8fh
EplYiCixK/bXg0Jh8gyqkOxTILUl3m7q44wAYeeKYvqadnB3zbsuMWKzwAHMrBGX
O9Yd/vRVneMYbOwQfpkdPk1PdcA7phoXSndYrsEBSD7v/PzR79qrV3rey5zrwby6
vAAd1OZzTBBJryabBUO1lxyjzWpRdvL9Rb8FRxR40d7JusINtxP8yp4M8qprUHSc
f/3pmIVxNT2drNdi51dV16gldb97QhhaT+Varza1lNmi+4a96iqONgbnVXf3lEsB
0X93Wn0g/387S2chX5yPWiTXqU/gP3TvynXuNgmiqHAE4EIfwDlnOnv7gk96zAoS
6Tz/KY2HzVdfLma+1NTmG2a9dHTt3egPsXdkatwKn16ShSkYtmd0DCEdxDuJXuZ/
/4BvvfcVIIx1XrRJ2i8yyUp55CeKoV5Vj0xeov3dpnVXSG9OaLYawhFthmEpyTN1
Jp1Xrf7yQgPzSNq2NETeoyp9GJYCfdy+WWJ1YRGwyhnq6j8kMv4cVnUXBGMDs+Ht
8PrNDuKjIUc3sK5QwkzyVKmTON+R0VN4Lb8ae3lsmowNaHTV+kz52quIPNShmbKy
+P57g6d6Qsuos/vmxsxe+o/IMhMbdwBoxMYB1M14wM+4yYiT9os9DhZaHsZiFUCE
qJfhMpVEjyUN8B5X2ivnEOGq1z/HQ20ZWb5dMuZnNKm6KrzyIBdQx89gaiQq7k/W
iV20kFyyHwA+LS8rTem4ujDVO/BZmPUDaVYZD8aSD4fLDhgmOaoAxmlCT173kuFG
VNJcpsJ4Kr1LCe6+kwN2yDQ4JcERqgZdrgiI7SUWuJdP/zKTSxADA7M3YESZdOxS
taf8ZUGbXqg8WnEY9h0Lh/2vJ4r2bDFXo7uY85A8rULQSwxyuLToe9a3/F2GrM3L
fPHGABDbU+EtRH25v6oyNQx5AStwuqCwsTawXdKBX/mEAU61ZTVqVzDurerQft6f
sim/itFy9TaicgQSinZf4qojoQ49nXN53JtwnAjLRxPCThYuUcc5p1aZMSKnOt2y
GrfWTekNS3lWBpdn8szuSy90WO6DOAMDxCyEkMimH6eTFpdMscVg4tJCiwyMaEOy
LFubgvK6yCYgpORXg4b9/D9mLf7C7d/1lczbi93YCNa8sfyo5wMDq1NG+ebclZ8z
vrZAH5GO8i3kqnPKTy6Rkab9o/poKA7Cl05uy/jGp2w7q1bVgGAzA8Sl9p8a6zA0
DbTIGdTRcQQot3inaYn3tZ5DoADxGDnrMCv0ENZDMDaAoIzS6k0B5yjm0Bj1J/t7
F7t6EbENXXvN0OgBwA7PTonhJW4MbMhpryw/cINHXZEY72cm79cNJKlZjXzE9ypf
L/wVOiVNuf/oQow/06/py4mlJmMAfu/4u6lej1AffYer+hZDHMFp3kk6P4E6yOfL
nP+YoR0qyLQvpTrXEnKZhd8/q/azDpTg4z8kITnBUvugpR9ZR/7hVTiYqeL6qCAE
WYt2CHp/Gdds9ctMazNlTiyBYOLCSHDSnQWX5ExB5bUnZpjF1ank7pw+0fsuggoa
01tkIu8lYZvGmTEZJiT5wydYyInYayDbRKG16+Zv+9DH7QY78cjHvhvAAPcvWg9W
b7xDE4Y/ZuatpvPRivKJn4IO7gPejPp5C1j28L2Y+4Lq9zZ4Q4VT7Qe1e5LeeXrs
OTNq8SEon0Bm47VnlbF7GpnymRDfS2hwD/muwSgXGGHBV30EkLwc2bf74uyundh6
rJ96oFntgH6Z3+krudjTopMBAFTq30fBBKwEr2eCy5iVqbC7lwRS5BHTbjN32GFd
2LWrFCBSgd3Go8NQMQD1w47nd/zALlD4USaRMUeH/7lD0YrzMjSHzkpEbYUHyHH9
fqo2yTAAqj+UnskSd2gFc1RLLTFZ46JKqPPgVwlflJm+yJ98/dsc+9sMN3Dk+g4K
U8a9zXbWs2hW37l8MqbqUsNUdH98t9bQhZl+RwTGsnd/LKsAXp2gpec9dcMCyt46
LxunyT2aVtsV1bRF8ULawgLxDPByI5o4trdbeuOSlbhbyRa/H/KKEq3Z2JN2bi1G
NptLJIqD8DzPeFddis+Dtw+3FFhsQs2vEpEd1fRpLnImNKHSZw9rcbD+hm1fz09X
t4WyYsZUlZcUgjbY+7xRAbPgErDyQ3G+uhiMg2PJ5ohXJjCr4jvMsLUudbU3DofW
u5zdJpaLp6dxJD05OvnKmLxFooQbrGFzBpvS3PwK4i7KmQkRBd9DtKVJHk8VQuqo
2KPpiH1wcqfweHp2sb7ddWu9Zz/i5YCBwGsEuvq1DpNw8OpTrMJkny+V7QWZ7Sfn
aIZgePfMOOYymIQ9f/L3SDFypT20ICREeqTL6DWUmELUYRdPH0XrVMj4u/HCS+Kb
FRtNc2kJNANNNIGNpCQzps0zZD6i1w/ycMDqGuoz1XyZNLw8LpMuZB1w8ffhNPtQ
FuzkEiaVdprnh4XJvFSG0Vd/8Rajbyj1luMY9Ymz1bcZ2A6bCkLK1p/xhwIrf0lm
nd2fqxWQ/7078pMUlnPNOvH57ncAqjTU+h6FT84hua5ydiNapn5rQyKh8zdNDpjc
FKtSijM1XTFUGafSRSH6KPlEek+iQK+VtnQ9mzn9Qe8K3NMU7SLlJ8jxzWgfuE2Y
X53BkYPMvZjHHamGIB+g6nIQzeq3ftSSodcr4EzAYpNh1srFbRLmiv/S5krQw7Px
jg9FLwnrwWMsE9kjYbvkNG+b43p7VtjmVJKtysP70FC4I3NT8afSvNhxOwcf54CX
CNY/6vWhut02iRwbKRbaZ9jT125mQBvK+ilovebMY4+BoUoOzy5dEBhuDdIqhbZB
u3ImTfkXLSJpvWjd+jtafpaXOCgC23HVKXhrlvFIse8FpG1tMc4fNGOsE4eO1i9Q
kBdSXzBx/6YFHxXIPvCPrBxn0FMMTN9c8XSPe6zIr9b9Cjub7g5ln5aT71ggfIPe
cmI7pkl6F5KYPXT5/OmzLLSmS0ySh4Nbg5XGBPN9WrkgIqDPgXpdmMXRfuqIohQW
kb1A27vIMaFR2JZ9H7rpXrdIGdFQdWK5L6fR/OOqel8iiU6xaUM3BqCCmsfP6pcP
Ku4q93JrqhBcqxYz9vvIQbH6eqpKuIkIebrgmYgjntJr56dmiDTc2iy176cqnWpq
ZXCapSEU/Bx7nCVapGPbqQg8295VfvK8t0fZR9OjdAZ+03ipzdmsmjrig7uks9OX
A2Xh/lCcF09xN3HEt+HmX91lfVHUuAnxwUKC/FyYBRWeAgDFPXxvVZIc0wG/KHcU
uyzkFUd/4EB6MJKqbUkvpBKr3XEShei6OuEe8fDdsm+XYNewK+Db4j8v5Qrg9e6w
kdojqmAR3RDbvJo/6PnvOPVlPdUxvPmFKwtwjRUtVZw75Iq/t4jvMz64wplCTYNn
/YcRio1vnT0BKRDb96oROedDLiGwun4YpaH2lnVj/ubXK/bYY3V5i8eb2pq4wK5f
UAOiot10I72W/7qPt+pqeY8BXFaUjZema3TmVvSGxwME+aC39VvxAGrhbRk+2pFc
UeD0exwQAoxa2/QRPb5MG2Wmbm0QljQLmpwerTJM5lHyxc9sDG2DhJ/tKv5Obg/Z
b4s4O0Z4jw3POcVZ3VlExBEsz3LFyqlaCMxHryiKZ/Glx9Ncb55DVFvN8ETAhwpO
LP3JRSID1iyyXV3twPskZ0MI32ka1+7X2fLsIC/VohCUWk2i7nOi41/skEn+iZz8
+TNSO7jlj3pNpKo29VvapqLz1R/YCS5d3D9oYW46gTE0uhEeyw7HfJgxkyWbFcu5
Zx0G24BjdGf0ZgauZJkcRHQaD3QoRIEmi3qro/cM7ETRWiOv2dQADCGLz2/SG+vJ
9GODCbaK4+/z3PT9Yzt2cQ5bp9qrHnsbTZCC1EFF68ZLMGw3UwhaZJd5QFvaJHGN
njK5vDM3w6weR5Z/jttI1+3nhJOp0DJRWvUq0rIJcZXUTbbzGSed8d3Q+q7eL//1
cdBvWPpPXpeO6L5MyXSaOb0Iacl3hGlNXzCUmmJ8cW1Ib9dwNf6FPc270syWU5wY
CU5SXKhtXnbdZAE6Et3SUnPnWX88NSGDd24S5BCWJi9ZVeFNFWNF3w3/890yra/x
Iyvb7WXi/kmUnXW4zgUFc8dX6WbYos4oObglimdIfl+jEaX+AWNEY1BKOb1//rKv
6wZ4nnUiZOvK51+e+E6xfIagwKOxLRm67LfL6zqYOJdAXgFA9cbftqvOzPCGzpdg
gt90xO86GDJHWQSkeBSkNzp7HoEDa1gZfrgdib8VR0HBL0HIds4LRB2VB0siHjxr
e8YwH4GEegActaQA4q2o6qK3UsOJADj//NNhEO3LUiEpEj/6bFYqfnXqmY0sPrto
F5RYFANyv5uwP+VOPpPWtly+XLXgB9zTSNkfLdsxCiRoHQ+siqWotoKcMnIU+RK7
eNGFgsj2QNuoeZAVP1hYjSm0r9ba/+EV+2m7B8wOk20rdwQnjtGhVou7YMwhOrQR
Uim118H+tA2S/xKtjM8c5CKxnC3BsvzEaYx5UooaUb13WNpoRO8RrBmK0DuwKHhK
vB86rOL7XBKAfZHPOUUMiHb13qVg41MRsKt4+RVg1P1yQb/cFeSErXDjSbcBIP7H
jMWnkdz5xBfa8V1wMuY9G0QBHgq8k6LXUyVrn2LhXT4dZ+GdXf8Me/ePdjkrpDWu
agQVaj2rZxQxV2iqMf22imZ7zLrzZ/7gzC/Ekd0oR6/CN0kHzQ2rgW/1b0Lt2K2E
WZFsaBYQUQfpXjOh5GRH36cqUaZSIsq1YsmWqPQZJriLc/9g3ty4c6nOUxAEPs+G
b5upHD2eVbqoXDRdqOzjaV6j+Gt3JWSuzLmHPptayAuR4d9svn53iI6/6Wj7kzJu
5TN56uflkbPAxnhcOJiTcYKbvY477RqXb6S6u9nRNdwHgUt3yrCfsFV/8tQrcYyK
qS2iIdYJLP1jRMhmK7Su6925jrmsxcV8Sgst5YzZRUy+mCK0I7OerVdQB/BXigk+
bA6963Xh5PKgo3U1WscRkMTE6p6BQfhvE1F0ps0jiAlwCVgMo6Ik9B9rHcrHgaB/
1PWGMRZEEttI2ymXX7dOxHFi1V36Dw7i3qja0WcSbI0XsSAHNBlCDqITyJyuPLD1
JG4RkCxPg4wOWl4eNNDRRa569GStPeGFZPyKHo7U83ztWiM0nEmyZ/XhdGOrqwcq
aCi4rMExb+p4UcGPD0rsdE9iUsxUxPjfQa/W2kcQOmjWhj57SzmzLCpLD8xjvpUq
aePfs8bY6atTQ4ipOYepp8CZ0PM7o8xFgWZMkY4VKysknVp1ZQKYxqrcTYcUNbkg
2l1Q/NiHnAOLMxOFTkSUdHteBY0erjn3eHuFvs6NH3Lwdz8O4seO9pzNo7f2bohX
Y2aQRK1Fqeh45VBphWnas4yoqDu4FHUIoWqP1TEpTx0lZFuHf4FLh/7fxJvHdTwJ
gIi34EebDruOaLn5kWmxDsQklqPcUhZjarxxrr1FfM2GPoqOECFFeSW6LKOtBiTF
n1+WkiVBPkIVS4n+CP3VtmM/lylebaCTzFQiky0hgnsf8F695aQyaH9Vl9MKG5oR
/+f73ges8zjLDoxz6iY98j5BvjlD8swDyfsXVvDMYknWJPPjIRCjhou3+uIOVr7g
gTahat8A1EGGJuHyL6CeiM7Yh6KZV0ousUbczKkEcojaAl9NCnore29sZ7BAMl7k
4FV3olX66h4JS5YiRFcOtLxvQT02eWFUwq0bPjhhvZZATg8DSzp+tgwVbLesH9Z4
FIqMGQ7/4G0cRUqgNOnCP/2XkZFzD7QFlMMzF9iZMfk6FAEucoSBTX05Pot2qX14
QvXGCE/N5w4MGMaaaWVFbZbL5EfLcORQixSihhYw9+4r0etavRuGq7Qsdj096+CH
ZucGbaw2D5yglS85SR9lO/+ennTr4VcmTv35jlbXcKKSDpaR76UTH7A11NbYXkT+
1mvFV5aUv/o8PUwgqJxZscMgQ1i/JP9rsk/6sPQyiMhtitNee+sgoEznrG7Oao37
LsZLX3vlmx5VVI1/pZrTK7qANDXJOBGjhwvFbKXtgb2vsY1Fo6W++UUco40Yn4z1
nxEg9RRI3xovpovXqpIBJePlGF2ATkZCAISAknErhB0SmIhB9OQVSs/u09VCwiCD
uet3eWV4qnHFdPP+8+8e4U5isjdz9lzo2zSzaoWPDPe6ix22VizcGz1qY2mHij86
v5P/iv7U0K8qJCVtits3YomDSre1ytFbPmyKHDJTgg/NvO6o59X24jcFK3d58ox6
3X2eGKvmv/Mb0ZfYfio+PZfpxw/c7dGYvcg4uBqaY32FuYDCX+1uZwUr8aaIjdW/
gUzY9F28UeLLhJm1SJcmWBcUdS9EyGyf+KdTiW97zDHIVtbZTGAQsYSJ+lWJatUR
JBruilH9w8VVIqf41RGeij7ZH4XqJL05GBg0joDGzUE5RJY8AvyyYcVNajod1nDP
UQSImXLMIgFfKG66GwW916D4r7ijKMGQcTVtKHp9WGET6n45Yl3Eczf5eGMDlZOR
Uz5lTStlXCWj3TQYbZbBkZnKcvRVzVhbhKyX0kxhQDIV/mac8x88Pr2hxaR/KVZV
YwDcTRpZspoTJsTn/ScXkIBMZK0xHnFHgeEsVlXT0AwvodxdPEaoDXDzvHJIN+fc
Q3MjFbJSnoswVQsSSlBwqwZ34u0hpeO+fwQfrotksldZC3DFC8kbouSuJKgnNwGC
c6Xsy8GbBkAhtOTqxK1w2TfKzEnxRAmlOkGM+KP/DRe1/fyhLPaH0RxcGHeOle/g
++LGDAW+TgHePnLrn/gDUCW1QgI1SlE/4T5NnNbbWs+w+J/3n96SaA5B8akCN9Px
1rxMkq8r66ORNGyidc/mL0VAxVcx+mhGvdFc5Nq3ioQtgZX6G/VwqgvBKpfp6gVb
jD7/Vse/2axMReDN5O+ZyZrLI6BwBCAAnTHMxwh1LNhRXCrW75lk4vDqoSEfHJyB
NhplEwbQtWrb/h++JWKx31ToAdB/BOlJiah/ei4Jq+iOu8/28rWG8FwcqXz//A4x
qjXtS/+dqY+thXif97NOQoSRwg+Xnlq9C/BZtnrW4vhTHAO8BnchfyTg5ONiksed
2Vy2DKmcPRsbfiU3k6yWt1kCuh2w9dJXjNh920OFmZWwZ0RiA+l3oLkH4xU/SzSy
5CfG8VwXqCfDBsdXILQt+HgGz6zwU2thsYbmNjIrnSqXhgN2ex+FbvQLSRW+WmJM
+oFCT9LiBgICprAP6qcZ8Imibd2V0gJCOFHJ1TuP/xSdjvCYQLn/vv5osVg8WwlP
gKjHDTeAnayC0nTcxCTcgFA71FpSSNElYWqweNsd9FY8SpzPsuEF0Dem/XEPNEkG
3erogNRqISGrO3om2oiO56Gfs/4FIkeiHe2f3ppX76daoatHgl3LxAkXDIxZ4npA
wazu15ar48uzgpoiseNsptwIYSEQQi0uPUqcA8NwKDnKFEpUWrBLbO6lvALJEu5q
wiFhpD9mX+f899HMyP3y9seQ7gvipw2PvXWjqRX3kKDBEcDm662qcmqNWegERbnX
uk9NDbTKJOd8TTUK5HR+WxOeS2ix4JVIdwE5Nm/c+g+853C7fHlr+XNqLGup6kLS
GzIO6KVbykkQ5s1u+/ap8/TCCTgvvK/oWQzj/ykiOMdQZ8qM6v5xd3g/pb5LfUHM
mSS6tU5aO5/vs0N6DhestpKE5ASTlgkPNv2JzAtvpKgtpJYEOdQNVZnKRDpE25Mf
RT6OgXf9jXpIoq4AM4XMjYf5MeqeZodYrKRISyV6v+Yg0W2f7VJ+TBxjplE9Nu+l
k5mNslCAc8gV7lSFwLjrM3AYrtUrT+ucAvXhCewmPrfHFrs35pAVK6egxnGfL2nQ
ebVnH9vXfIylBmN/zC/u9GY+YfTaJg8ChCoKvsWU/1Zg9bFL6JgZ9MGRBcKmt9VS
Ly+D6254C3Jv4tmyocyDycJguuW3+dvYxPxhhVax7jPVsuWnqh2ROu3FcjRRIAeg
edwKXs88cjm/mrcavOaxWLVeoN9hhqszwqxdB9cxOKpmSzUygq4T+pvycldXme7K
XUF6dV/TY5YZ3VUDrS0nhfg5ixNHv8Kf3rVSFACbf4+M04UAurwfAkJvbQFYIP7X
6PMpIdXMa57M15RuawcsxoYOxnpkAi1pl9ZQqmLU7e0Vp09HIcSKFik/nPynOWjs
FPFPMM4jex0s895BVYlLriiTEza2kCAyybXlgZTaVljiOdRHMbhQkQPrHm8pYAly
Te5UspAHMUMw2ATJCXSP7NLBqdoffoE9BANOjGxh/tElbFV/vUkvk40WUIIIW0lc
+Tg3R6BbujcBvbTJTDwO4HUTH1xXpM3b9Jo6iVo5tQtChhe2tYFs5paTv+C5L2d4
4x+jfb71Czk2cN+11wvSJzE4VMpPx+cXvaq4e1LKe4F5o0FJCjeuwyPkolL5Y9q1
oL0BwscL41GJrASNHU8QZrki3WQOK+mYQLMjA8wgq4YDiQLxI0QQ6yON3/IdwNxo
8S6NMlh7d3q6c4Ap3UcS5BgDHpNVHQ5c/1HXzXVmG/bjqCMut6w0w4zrMHS4JTof
2bx6QzJ8APYXNzjl1gVFQc0Bv4GNRZFoMJR2QlA1qNh/Cri6LuGb9U0N2NwlVeYw
NmEZIBGlCTMw+jvs9CpSu02AYUByhNTF70J+y93Bjn1pF8xczIgyeeeTtFHBMPo9
NU2ykUYZM08Pjy2817u3bDe+SueWaCkPETMTlTxDwekv8tcrtaJK7B+BZjYgJmoD
c/srJYBdk/26JmRHUCSyQtxhZitcS5bglOJYyNwQtug0rMxKKvj+3o7vHggWIg7X
K3k+7hIJmfzWAaK2wGZ7XizHhORLALU1QOt30f1CG/9hxUE2dn7jQfw3KfS0LD6x
lxBHwsWek9ZyP6geTabl1RgN/W9nrJy4NYCUsJXq2vX6fKX45bwHXTDsMAkt6l0g
LLkLVKUrttJwc59upwMNLSwmTIEl73XHaqoZllZHa3+PN5T6iiuECTYhADRH26FS
JmgJkH/YzYEDy+6zmLtvQOjfEOTCxx8Two/oF9YtJ37IrYC6OEgmMY+WnPStg7Jd
+YhxcU8pTJWaMFM28WXwCDRE7wdAFopB6U8wGk1purOBM7EeUNUamVA3bNm6VGCU
6EzPi+BQosbAectGxklqc8/krZGP8IILojASltHmoXrEurdRgd9/5tS2LU7dQce6
8PjVMyYilhdOx4w7J583LuRt16gYWmBqe3zAP7xl/ZnnakEGvF9TOfhrow7WZBS3
sK7D1N27PAJggYveiCJe9v63eBsw5J/ZlL+lX5EkWozY6DyV32OTYYDZkSVnAKUu
F+woO14fB41wtLjW1i3d/cDI173uT87WYiiTiEDVcPBb/b6TeDcDF1I/PCeAPnNZ
QwubJ7+qT24IEFs/FGpXeRCce+c/HHjggyOdzapzK5hQul2eN1SPbjJSe8cfnIGx
d4UyzsW3pvQqm+g9Kujrk0lxSF+iJYzQ6fGFzU/I7Cpz8cNqO+Z5lTob/A9fjtYS
46psIbb/amjsPnki9duc6hPfMKhE9HC+tWgxYjGMIojF/Efs4YNWeSGQDxBY96d/
Ficm2ZVs4b04zOtwT5bvF+8YWDKHbmNU+v0vd0KeKg0I27zt3kf0QLsFzFJregII
uGtpdss/bqjyCzQhOuRqxkSL3pQTvUKwQZ6skSBGofG6Kt9sfmrqjSLDtfCQEEIC
RRSN04dfkQdd2GF7kuNnJrN9qG/tJvehStJoYLaWQSkn5BcNClnfHJB+edtVAi/h
91uGIkQlLLMDAhsAL2ywWq1G8cOlEpBD0YBF7ZODAVHS2TX0xJMILiz0EXG19Agy
HovVJrHSRLREkYdB2pwGaHClW+bAu6K+SyHW9oe3bSufoN4lH0SnJ/GUR5r4q5gY
ef8eg+Oerp1g2cfKhuuE4LnuwuY1Fy2p++QNcVxIkQ958j3wsLtngyPvMxA1S71p
mMx8tpZJvO3n3vaBQfjAMDM3JDhnNZbEXcxhjfe3oH6OOe/Gs7Sl+2zXkVbs8Ll8
00UFmOazG+LA+5Zwf+yr+MGtGjDxQD3H3A3D/5NVw4Wy0CYt+4nGM/35nmKBwIE5
xiu38+k7mtkryEc9mihOsmudXGomuh3jYtDOjqW+zi2XIzEOrWtMv9UpHlakmPDO
1zWYHs87K+JQvdlCImvbx44nZrzjzxGhveh11LS5CT0wOH/oQybt1qARU/a/Bx33
RDHgXZy3iHjiJSM/6VOA7n5tT10NRmfwAXxB42GI8bSO0tNCmBO/uPoazP9fAu0E
QEw4Vwe1aUS3qWjV8TpHTrdzaM03/rVqGeUNTnIKIi67+XyvjHQFophqW2XfsiMu
Wo2R6sHReXOBroVd+1hCmJJWKNeKUd4J3FbEsx/pghdR9lO2Pj17Lo4SUbroMW92
7Hd+JTGJ5bP5ceFt0Js7NGwYM009awrI1GWeR5VonfpYcwOMa+p2m38RD9NqyPUE
Wp/vQmPPnEFH4Eehl/VE7Bn9P9bzs1U6CDAALbdfmCkpsxhDxaIkt9zeuZPOECph
mMkOHhAYT9zVT3CcZ41/RiMZnKDCtVmVD+GFD/H9uRQnY2+CB9KJhQCQG5CP2Ity
w7Np9aFnGyUvCBr6cR2TLzI80qwmAGaIvXjYHaFZzrrxAzQDlXj5CXBO2d8z9yxl
3sUVQNFHZNtAgTtpOu6FyxEo0zWs2krjRy1Vw1CzVFodYHVbrklxYEIGuez5ghaq
x4xrJm8/YjWI9o42tWrVm1FOd3ZBCQO5E9CghSHUfMsT3urAVHCGZuo7RVMWZNx1
d2eXfxzWyZnARxgDKa8zS/6t3dhnYoKfYuMTnQHuzeEJygGu3umlZfVny+NI+xVB
SYUjxXTSE0MqND4Id3ZZF/H6jh7kzBzvmJOXQwb7Gqg1ChKe9I6p+arKH+qdT/vY
1prNoDmaiew51hcUyp4xerIvOBxBeyxuB4MM16ZyG7RJfZQd29B/Cb2n+9GMxI/+
EGr5ylt9y/Tits8imaccF4U4TfiM3FANPk+N/4L0qa3O6K8BSwokAQ7zmrKTp+fC
aYEPhlcci57m6adMi+9Syp3zyU0zcPzYfgXHPj6Oawe4JwOX/KUM0LxUm968FPjC
69+fEhkz/OD2KFuGUL6NrUnOvqTUZ83DJvJl0Md4ThQAfZGRqMcPWYkVHFbss6s3
VRnOmnQ3iXV6e3PIklBAlprY/m02H/n7YAj50rbOfQI3Yuii7a9LGenPte6jITxq
kxAnVdljLqROjZT2sPywvs6ppIiFwKpVDBVOGZfSCE611qIM3LePMp54OKtV4Po0
fGgYMb6Yul0QY05gUdrucyk5E28lgQakOIN5AkEI5QUjJ05fWFYujN1CapxPTv6S
tGVl9/hJwcRc+TIux14PoIh/870MRv0UK5LGVLKfytZ4k1xLEuhSr7adM+5HqPBi
xk/2XroV2ENqSxu+WKW1fyROgjJoGtWmYvsz8cWs7S4wVtfdRZ2Z5wydL1Kt9jUT
g9+mA0g9SLuDrwGa6oK+YVrN7sEzG6E7WH3h/Oky829Lz+jCbfkjHA1KF+cJPoQU
TIySyJ0thUuRFsrFRI8sytIBI+yCQmVwt77QCQTNqdu3AnzCmWe52MXV2MSah2x8
5sQ58R28dPkaxhpxweETmICjJQjRNxJ/L1uhNWZY8zTpuCyef8v7bD2BbetK2lvi
vfy5Y55sCsvFUp+E2CFdskhYn+7xu1q4GcDiotmUJ9k/pzp9LToISkqYdpSE6mGG
xM4cr+ycW/f23V0yd/4btMcIY+m25o+2mA4rYj71GgXMhuH70oOMP2VqKukLpyAT
Ypdlh5I8lYNYKtKNSzzVqe/FuaoN+zrLEOtNWcZwB5HPLk8p7C+QjNrlb8oO5WXH
hpxG6L+2/8AQtdghYO5L9dqBfhKPevAka3MvLQFh+MTYPeZBtCnijkSxqXG6Mtpm
wZaVtYdXSP+TzPqckDJUCvPPuOQ8PWBuZtvu0ARzqC0GZx9tBHhaFoFm1jcVwRzb
R95Lr+omHI0IXgOqoKZDjW32zpkdwDKgPzKi7U8++cA/Vqk+898Vtq8HqSRbi+o1
rgNcOdJUS6jdk2/W0DFzoR0s+8fJAgW2vRnFVe1em59FdF6UpjVF9jgj/sjmpdZl
VyTdFp/B6EqI4N/iS+LcjwmAeJ/xgh61XUI6ggN6r4KHfPPMrizfLKtaeGJbAi3d
En1EUNrxKg1svtujyc5Qq+qfvQ6OzTKHpuYolJO3+9TEhIOTd06NTt4UX+9uGkkg
s/WsFBygA6oCmqzvj+4CUSPlWh4vHa7yQTX8OraTVsrXL3UB3QP4Jwr6N9bzIRdE
gIa/ySoaXJLePABfROfI7pcJiSow/dMBgmsvuv0Xsaujr348oDxZ4EPTOhg1UChh
SaCs8NHsmBKQVqmxPJAAvW93ml57mQz5QCmUnarjqn2lX4vD+n82aJDvj3siePlO
DsEYY9VXtCWV8pjDotsHu3kuLxo8jMO6V+bGIZwDz8MFHtKWGU7RMBIwMhY+P19x
ed466zjyPBv8xZFGZ2E+JzcZWI3nuG/XoqTPP0wGr5H5/V/e24AZWvK9732HxbG0
+h7MrP0DHhyfksHN/8OqbiGwuaIUCWVmZuCK8+1zVIEDITVUHhpAtWxo5OiioMf/
Dqo9Uj6qr3qiMDCdcbOhYhNxvIYruHo5qSGLUYOsSGroEEJXFNstQMbeey4pv1Po
jG74LPlcVvHcwXSHRslcFkb8KMbDEmhd03ku5vHVi15w8SThOlKaUrDuwPUvqkET
6Sv0sXHzp7tZD3O1r9J0RHlxj4E4JR28HyEQpXzaeQgYp2Pl8ZtL8Lk2xO1qWZwb
Ex6aTVzo9wH+9neSXcGnB+kxg1y/TUziuwZywihJNV+jc1kORSNjGhPcn2fiS0Hb
wK3yEal0XWM+vzVX5s6859SEKgM4tE/Fnk0COj1e8BbCdgyySXbdasnC5iOCHbb2
y63+sfl/NEI54Mcrekb62PjlAhIJA2YJOa+bzZqLJeDwl0CEVjbuzjNUNc+Adh2N
ndO3NuYFMqXNq+geAznUr2vwqgaRsFqsJaDuvFr7p5D5v8HbeJpBPu50KHK5YBPg
v3tIe8eZvSKTFL0zIDg35l4IHFxixXBh32BOUbrHBJpKPi0sBMmeJzImcrYdhZSf
Y+PB43UkjtW/zRRNxea25sPYKoK0evXv3HrhCLWwHIA+AwxTMfe7KaHJxCwMXa2Y
hh084u6sW5g7Aszkw+T+SLszEjTNLyyitJwDx537D9iCp3shdTGLFKJdV8VtXaYh
VtUpIe1T4sYVpKdmXQ1lDna/ZHLzv2ewt8AlqaXG3KTIwz6vOxlfmxlOTlwzHHg7
ZIygBwVOJ3UOgu59Gvf7sJGshI+9cAStGuJTt9hT3Rea4L9AsrjFWCL91NMuN9Dt
ajOgOLdcUyQvZYlDmdzYX+s3QY8Lickt8cQw1iBTxowUK9u+EEpu4zVIHXO224Sw
zReGByMoVl2LXl7QkgkqsrPw/XK7IbVzopDDHFYnBvHm3uABrdcP6PkNolxFbeIc
oM0OwxmR39+43jKG9aLO5Vu7+jaQnRXQPzHbMwkxIsxxPgPyqnQNvYdan/sW5Nn5
UjC5k+c24nixv37wZi6qTJM4fveoZzP50zkv8/hdaxDecATNxDIbJqgE/RykeHLB
G6BhVbqf6q06bBYExBXubngsB2kq3BJdsRnuVQWPRAQ7IKrKr91Q4lLyfNGb64YQ
zhKfQUmP8GAVxxzdGnv8Rc4yhLZbfTtzN7JeC/J0iZUVXoNtR33C1uY7upO5s5Wi
KSzgXXhVe2ia84JfNVCPC+UVjRxYlUsvi9rf9L2K/Ic6yzzwjbYtoV6r/vvEd4By
2d0xgx8px6QEFPdpO/Z4/xWLmB8pMymJdNpEOKdkMpYBabnsN1LF1WZ2Nn/0FxSu
X8Eb/bpqp1AQ3LPdeS2C9AgU4QcIHWuCqr94EJmG7L/tmU/COjCgBCQD+SDOGNg9
SEGEmC4ykW1qEsgSsp4NTLvtyt9fWaQNXl4yvGJaseVxqj+GY4WYTl4iqciHNwWX
bn3bFhUx1xCEEoVmejBwKTNbT2SYRjSx+P45x0ij/2ojKmTeyZbfhwMkcbAAtOsz
G/U+NU4V8LpwL06b9dLILee7Ycf+J167goYlr1pu6EHEKTr/n1dkYN0VQ9JtRIQH
pywSRVXurSVUKXMzA6FGrzWerECwJUyLSOK+oMvaGruLZvWumMbR/el/2xMmznkn
ShsHEHQMPPl4qsa+lYAVyU2ONcZkPEqd2MENppH/iS6qNvAAZBWYW5+0EDiNR50c
54n1lriqNpKSeyXAyC10OnUSMANokenUOwv0ZA/4M7riQkbRB1LISTh5L04UuF7n
/OeyK6xSYWaOGX76HwMS0dwQ13SF9PIMUPxVj+wk0uIuf+T0h+6Qc8nMe3rESpT3
VYVddtwvG4iZhcVbi7utqZI3NDkrsuDOkTgAjnD5qao3RzqxTmE8kI2iybbtYtRq
MxPX/rRve9d5CKTEtEu+cSBRirgMhh+o5/oB/UYPDQmMmlX7hVGPw/WFidMKC3YL
IcgYT74xKSEjIRF63E+/gfbNIM+7GN4dwFFrpqb5l1WLPJkblp3OOlcFiXIJoiOZ
l97lyy/YYvFlUIewka1hPIIrqCPHVAjQ0VLksFrjDAb3dOARFwuXtuNrRi1IGo4T
nQdLAw10TiaclVTeb4bQY2XIMWsKhGO2UlTFQJ9nbrzRBByyyeA6LZhDXZqamqsp
r8ib9WlLX7Yd6MjPEcpQGSaydE7Cis/C69A70r4kM/vTx8tYofLYpF0D6WOQMjuD
aFbto/GiRZxGYlR5cOhLWbO2yHNnDFDU4sRcTTGHGRsSNopQwjLwpPSoCS+sQ3Ep
M7dBbMkq+yDVdvan7ggE98zKYAXhfxinUxVpWlZQCwezUhv26Ih8a568XFr5kqbY
1RSqs2G6jNWLGkUOgWQjmDaMDOO0QucNS/NFIjmSdHBxM9CkcDAgHj1n4rJGGqak
AkAw8mRoM6FwF0gVjf8VjioybUpnsCb8v0bk9boFVSVw+4A4pkEHz94HFcYkNjMY
6vOA/2EOUWC6FnF1ZObvxpkt5V/FK8fkGDI+96X94kZOxUtuk/ps9ncn2XaAZV4o
bc4ySc8Cqju4Rib7rEGfUESZrxFdoG0zcS60i/GCFIfGemYuJgHigRHYCONzADSl
/qkXouZZ+/AKpeHW8wOFZWi2S3g3xCbBVqEF+KqAuU9VDpeID0tY9xZSUhj3/5Nm
zelsK7rTEKibjv2filYTpECThwBd46NJxCviXhWYkZgUfSwm4eqVW5d7po9PC8fm
Oqbuu5m//vgPen5IUMYI695tK06kMiLezeEvaH8AEIF3ULP2GPLUNLpPCV8dhfw3
fyyoQcHrMRrT5aQDOdMkkSYug4lUcXvH/eglbiVbp8ZoX4sSTGCeH8LVHnZN3uti
yIwiXwqnYYrm2p5kfvuvyJ22Xk/TP7gpivcDqQEUxO95eWU0eTHVpvMjnDPIXz0F
AzenFGKnjm/eo1u3E3pxC9N+OPJPRvVxpxNgXpUz4d3FN6rXSdWiTBvpCuK4ZPJi
x+sDMMh1iBv83tNMDdNnMjv7HS7Pxs99HD4c+/1Nt5D5md6vMeGQAeHkFfKKZoz0
/PyzXuQ//2HlfukW+cUD2wFjYAUFckSQXGxOTFbR3StfDaErIR1N6ojpwtETVnLi
2hGcYcUAC8qU/FLbWfTVowzE/BsjFdYkZYLaPvSgwbNQw7BCqW3JpGQQe4CnHgcK
IZleJxaEMKYgQu0gXnrEtPhb4RF5h+2J6RwybPZml4yqy4EgFeCbOk2Dih/bSjR+
6y6F5H6Hdg/3jh/+Bi7Wp5MbwGhj41SwYGGpN3zGWYP8BzJrKB+5wFCBOILA8lN/
sR7aZaeIJBdd+ABf3aBahDPy/IgLm+bosdo3VFHt0uO0Xzs0vv7TudUUq0gIDqhP
Wti/X3F3+5w9K+oFmdpGCha9DGEBs+RMkLO1OaM03UyGJrq/sPjC9JaDpyJTFSX3
aPbFS+YIWa1zmBZYWghaQJFHvGfZHEHaL5Xz6o86wKpjlxjs8jUXanOf9+C0GGbP
Qa+XRYR65Bzcz+Alq/8vgCeHyx8Vzy0tjN730picWRlg/4M7r81PjXqbOjZf3VBA
KTIuaE2t6NfviJgoqqnWE0oOCapbCyG2ewDgDNUxbB7Vq9gTxwINnxHA6NPDMkBY
qKq+beqki0JDPVMs9Za/WQg7YUDdR9khc4CkUvkCDcZ2LXrLXlioHx3pwa7FageB
GTD2zoE7iZIzqbWirt/F0a/z+oWQ9/phCfmi2G8Oy386wN5r9b/vq7j7Bh7GD5e6
NOMqSQv2PRmu15nFdcoNVybdfOmGjgEmLX2OwePoXMUj8pD1cAM+qGleTq4M7ey0
TsdXe0GK9ETKoMaQOk8jBS4VouN6mMRkNKB9MVN9paWBCGeMMbEHRClapD1VutWO
Iih8wonCdPVKiYqU/yzFeQpiCDCKGxH3g3Mc8ERXWnC5WjgGK20RSBAVbGtjyfa9
x2bsc/8JSWaZi3sKkVz1ZnjxO/LewW+F5rPbbEVaQuAawnZfo8bHsWokhzVJlQ/H
5qnN25v6DFgha10QvX+0+w2tCY9pQ8GiqtYNiGd+ZfgBGekt3x40GbczZvuJo0zr
B8cGnlh9emSsoZ2v3DAzeyWjno2bW1N5egqEsqcnXT08VMYV6xaYA6q15MFBS2PM
TiBz2yF5sylXPdEyEXKJBr7ewYZGJrH9Ul4TwRmCtEgB2mpBImq8BatV4fEzLclY
dLj8pKRFk2LkjKwYpQd70Lvzl8e5r/rOFnbBTjqGq223vG+WRZrZEkyxESXp8/tg
kVxSRlZMN3ayUSF74ANPItolhFRC67jjfRtK8xV1hwEdD7v4PFLjRflmjan01RD5
Ezc69Nap6amq7i66i30zqu/mxpfNrzt26TNUejztzskoekFSNaMsCwtYVnSAAaOr
FfvxBg1G8OsLhyCUwdc2a25t2Tv6WS4gXFy+Ky9Fsl3A8+Og8WD4XYhFbHVU9zNT
/4CBwuPVcLzpWSG6BJe0W/9oV3S4UO1UfwiMNlN9FCXe4W/Hs0YR4CXlD+VYwKMG
o/IGLao3OdDGwrKFM3cjLmIpLs7xhFSiXjZ+RmEZIcJBH+OkciDVZXd0AFKDz7jA
5BXbBF/VoOIO8VMCxc0/m+IP20/zQfzctZFdS5gg7J0Eqh17L5BW9EbNmCvCr7ei
6ezalt7gH4+yEnw6RiJRTtV/i62ZkDTqtYi9gEXM1zZiUP+6h0wvQHX2QP27JlVA
ygXRtUyajuHO9bZBxv/GM92HBi6V/sO891nwyXQPFYJAXDA6ZSWcSybyA5hBnyxA
65tsmQoafsYrSmXqu7oKhnpW9il4OqQdXH1mD30w8enDD41GAY6RzUsk6BaZERbU
yJnxx4U2kKHjn4oJJr5GOMq2UFtHwKHtrDeelgHE4fiK5Em/XuxWsIPE/T8q1sdz
ilGAwT8f18krsbjnci0oatLB5/ttLgo7T0On8k2LsOt21up5EZxBP1tEUkO2iwA9
JOl+HlZHHUtJ+bWS0INqQIL1YtJmKubDDOqzNZWRrF12CWOnX4HoN1O2/X4BtKIw
upy+/BSHmRtuzRN7BxJIYOpJYE8MF+9I8YHIfC3jV3LugDGTiYIFbDsEUKQ1pw5i
hj5oPTF0Xh6iSxcL+TUkZqx492Yyfkuo8FBKfqmu+vpQdlZfpfSpxgV2/FPQ91/0
U8Z3vqG4iZ76zep/vWOAzTEk0VcJR3H085kQldhLJoSCbYPq4sg5azJZs7Yrg6/m
JcKOAXSbIRmpvIA66nyUemckt/z6F9AYBPZU4/t6qKYTtzFvgAHlK2Kqi20IS6Cg
MeAvBfrh9CDJEizwyTaAUIg6RHE4oy6TQhgcWSE2LUZ7J3kJe1UqijvDn5genKjL
VJ5vr5OLS6KnXnuLBNI5QwDfimyL4ofNNsSq8SJdahFJjunZjBviWb7lrBZFDeXc
8rWsKhRm+FYLSPTD5Pou8jOf/rNNoynXmcyTSOY2+xCO2WfO4xivyVLDGPYi90z2
4ke7UmgmdywUIVPHt97Tqrppi2LZPgUxGkW6yJsLvZrl1PprsOpKJxOEBxkEqq1y
0gQ4qPSFETVL/XVVGrD6Wk0+eAr5m184kVWUepwHwm+BAFntEikVUC9VdcCFZgJy
7ezAGl5Ri0YUNMs+KEarjntXoRCMYv9aq+Jr1hpkKt4fIVs0qKc5OpB6oDmx7Hdc
lJaIDdKsgeoF5N6HlVEAHEhS8t2TgSIG4EIRqAjXNnltxWt2p2dzqGdY1mbvhuTc
3wOEEnVnOqFqlyc2iU0g6m8QRfKLMQTqjPppntzRVaYY95rHR/pBv2ux8qOjABhe
NK0ae9Ib2oPy1n8rtW7T8gaQqDJFHFymhbP6uG4T+2nAXPfZwdYlgq2NGXz/7Frq
StZ7Wol7IT6izEfGo/fX2NZuT7bu0XPYTIB6+5wEMy1YG1vwQPAAHCHZoiHVRKtB
agfLgl5xYW3mKyJNazNAbo+GR+XsdHuqlYXDdiUBgS+SIjPs1gctGLz48LrAlyg7
duThbjbs7A2aBw46Mnc9ZSMykXmrKPwV7+P2K34qitnf2RhAV9aKPNXIYQmmU8hQ
fAf9Cl0l+jdQxPLMC7rfsg5Q6/JHii8toVY8n1W7/ILnNikbjPghlGR8b38uTtzb
huk97siytebPoqtRouxWGq3dFzHxYS/dMYYzff3gWJxkSr0rM29u1h0AZSuY0geT
JIoT00d2GP9D8WBeEkodJSbq1scn/CdWjoMmFIBY1WyMmbwyYRKN6eE41NYkwV3X
xxCxPAyTJoekRTFRwt06o99tWsVZ6yu0AhwFgBwkvu+xzF6TY2G1d8Yvw1aecGnO
PWYIoIQHWUwygdLlc3s2irOoDJZciFvprLBsSaIodvpr+qFn02WlUs8Vui7+k82c
JiRe/dZdlfAkeOAVgVSGrpJR8B/g3YmOxOW91qiA26pitsLz7iTizDqNG1peHLH1
Nss/Rl3N3QXqHsvBQcaekh+zCJCGLIq6btpQOw1xswxLNZjY1gE5w+1ffgHROYiO
BDsWVdhqOOHlaEZfAjPYUriVbvoCrrV2zYCmUaZmr43pjOF2iSMVwAg5b7MpXiZz
mwTZmIPglHRugof6o/0sFX79rIBqmX7E0I6jC1qXiRO0Hi49rSZRaq76q5yfzWTF
cbl4xif5XPbSy/RqVIVryU2hj/7zu9ll2MAg+Uj4wGZr/Pb/zjYCShYPPXGzODA9
5AgKBxtry1pBWltFKaK+2NlJL2IgvB8hVXwUmJeV7yRWDeYjxfBzQhB0/dGLbFF8
ZVA32fIGK94fcRZX74oI/+K3OySNPsWPbjU4mgLDXlOvmQyMw5+TJLknySw8owtS
zplfGKhcH4oupDticffaHbZGnK6GaHWz7xSt1unLz5vmvchYns6/5i7zs18KXg6o
ARnboELx10KPRVEjD+fM55RS6yQcGCPIMVTcI6fyjzaZzyHcfw/qtf72GVaHdz0J
mkaGuoeVjpIKiugzv6fSGeB0WP2SGgK7attlZwcnq18RotoBRE0h9hbO9lSQeCrh
pgyg0RwRB1O2fAMWxW4sHX/oF8rfhNwy/YUoWa3WEy3hcqT/Srxfb5j/+DOUIBq2
ri6aukBUz+mH2sGExsYOdrc/OmKUbOzAralhVz5oA9VuFAv8EcwNO5vrDNVdXvLF
WwrCh9cXUzlApbYeXph3gfwwUwXGl9HQoGqPREs/S+TOiDthpEk6kZMO86e7ZOxt
n0NYHWa0cNjZXsLO+jQtsbvU/flFQZAFa5wA8x7eE2hUblGR9RZJcQXk7TF2bjVk
FEQSUqvIZhGpITs1Jr6hO8NnqnQ5ePaeM5Vh5qwBvTYcU/JJAUwYG6uLZZcgf7GJ
5Sjgfi7gzD+YTX1c/pfyM7A1CgpIgCoo0ewuBXWsxYjgykm1rzv5Cgop7tsYM4t9
Boh5jlhG94DwHgW9Hp+BH8qvDy/lijGbKU3dSX+dH0Yhyn3Whv2fVlo+lAQaAmc4
DnWv6JLAYbthItlUDQ/p4c0zix/0QRFZIL5FgSzZUHP0C20m0MtNTeWDUJ9JsnNh
2xzjm+zfzVVF6shCIAS+m0Lph4tS7GmUNvAIByGkLkiEYX+W+/R4Prx45A58doQY
MFX+4pgoo7d37n96mmeeXa2kaV920I0qryd9lmUC1c2pa82tu3T9RfiR8oSqT5ys
Ky8QTm/1zpVcy2P2fAC9bgbQSlfOPibWCEvugEq4xOMY91URiDo2ENh873o4uhHR
J7/i0zEy1wXTck9mcopf8/XJbKgQ1CYoUMqEFNbqr8B5sylKFSZHoY1oKcPuuVAv
/6ix79YxilIfp/3mEAxq5Tvn38l9g+HIOLEZaXsYzBp/FxFCjc7Iv2wH495rCE0I
f25kVvRoINn7c5Q1zIskizi7aBhtSI2GxzjXMmat8EI1J/pxI4MXp2b/+GRifeVO
d+UQCLjyFbw3qE1sxxCiB1P6XqeskYQD8r6IrT6MlQy7IW2MsdBv2I2NwsvTMAjQ
VcuND7dY2UJHgxTuhK3S7efbBdUGixBALpb4sGjcn3vm99Hr+WhVQvG0sJQpUW7D
vDGX392UKK68D0uPfY9/JVOECVOWejmf1ILu+WbrYSDW8aCcLjCHksUUMMgQ8IN6
Ucrq4+CqELgRZaiyjTKnVJS+8KKuhOeI1E5ygQ6GyDuYGPGclcT61KmE0UJ+Mqm4
CiOYtREeVgkE25if76WRFqJyOJJlq5AsTlwk5UWhiL8HMy1v8p717h+zUTJElpQ/
4WyT4UFzF8kF0oolLAG/Eu2NOVf1B9uG3NEvHEvS46pxTMISmcJ96nIwBknfhamp
SUyT5RhRKVcpm03W78Yxc/VIyGktbZpjvcw03mB/2GfT+qAYha56Z6BoV3wkLG9j
9bIWPvHVjOmH3iU3t1E/KJuq0+y1CN2kRqTu1u6snv1fu+igcne47Im9p1mbEPXG
LOa91u7rzyrjg8CV5rgsF01CsSWyrnOVFuMlgi7j19ZTtcbP4bauw3cSycSvIzkj
E1DDPhEt+xe5ZreWCZzWtA+rG51UaYY7EQKZVvS2ME2BJm9sGNlJRGhzkWFUzQhH
Vmq6CZemHPAwxd2DxFYFavjrvB+ML9coOHC5mM9vQBBRyN831Y3al+PLGxV2QDbR
CoU2Ci/y3LM2fFcDrUALmGjeu3GHaH7B6COaN0UQcGXIB+86jH26Bf/JiTww6vto
Nw9sSLjjSgzGwRfoRDT7I90f+nbZ2BKRqEzj2LT13OhL9g+pljzK+l5DLVQLJQVj
SAYCd/ax4aoHnd8B4sm3/p7ndle71JDZMNvafTep07gnJmJAHtZfDHqJ6HMXLD06
ES8ymjgJn5ll9Thq+w+3MkVzbbphH383xgEGjS/s+mutxYdcUEjR9Pg6jvzwF86S
+sVwCcAFQ6ANS3DUoV8To4FNkzvzHITAdFSPF2HPfrHPqO999dRekZzelBimlCGq
gglUeJEFt6Pt9V09j+/ntQAHtrf7VvSc2YRNanDcalzqtvNt4clAyoJ0SOMYInP2
wMbGAmjwvjrSMxVxkiDxw4ckGpOPDWiAosW3uGaHwypsaemE7d/MFlbEm5fZX9M8
0XfsBBqvpVSrjgaRixdP0OLU0B3stXY+NPpO30ExQv6gz7jzhRENIab877rngAMl
X0b8sLH/HinpoynPMBF5goSxJcbdytsDu7eMXwUKsYVNSFDmWfSOMDTJfUasHdU1
yzzGUtSq76m3y5kzmQVfmyrsUPFjvFLMLPxCupAPVlGsvFIsUSxpRJ6U5Yu0x8rZ
UHT/NBbwyzIaHuRKsBQM0D1ODnPRQO5VTardbeshcAtYtVtW9QfGJu9regwHc7bw
yaVRoqGu4ujrsAd6RgKNB2l7shslyqGlHg8/f8uQrs6pi1vpVaYICDbEF9rHUSVZ
6tYS78QPXxi/lDu7gk+OkJsYoepOTCHJy99q9ZRS7/ULRXwbyJuzc1+XzUPjnFBJ
a5TbPG8LWLEfQZfC5Pk07YyKFCDFOMlIJsmfukAPtmNTobLGJDlmwACatomUtjwf
DnBwp+YXiGqw+uQPL645PER7ZUu6zpSWPsP93MyxTwRY2ImCKi/UH7wjm3srKJaa
81rCrToPN8Of4jxpvQnYjVaZC7MFNYVWVSSL17EuANoX0PtjAWuCtcIYjN7idSuA
/jk3M0XwhK1cKzq7yWwQ+AE5m2vD1Njzs91TOELp/g3S1a+Od91Yut5ulv/rbKr7
Vsq6mD2P37aMaY1Kd2uuTdh9bScAnvnACv5Nbz1r6YP4oD8pP5TNlGzK11C00WaM
ckBIsDXAG6LD7+YTNLvdxULJuc2dQnnuYPLTuV93CBxBhUZho4Nci754mtF/T4+B
WCrHjlvjWiOipd46F677d0nA+dTamKlBEW1dFNZLPZXPly5vHhDgtQCTaKDQXl4h
owZPZljah+hrWaQMxot8tD76om/bLuIcW0oxGLRYpc8j+4asKtsda1Kr2ucgxajR
BG30ttT/zXdUZMo7qrMyURK2vVik+fkgtdYVOZIIOsVPceJ/kknoLtbY3M/JzeKo
NWB3C//viGl9Uv42EilzrZlpHne396nRaNqGpTMIEJnXbnH4ieU8CVX5PjayYt+p
vQLERltiE5YQUkhH9ZN8Tp7HMYLQig2bPzi5S+81ARINKNOz50HbI1Eash8Z9e1f
ekDnI9dHEZYUa9O3V4XasM+Aj5cqiFxaMfbZ6VqToWNm9sq0H0cD1sHg6P2yFPyh
ytyc58FRFM7fY2IU2qVuWFfyalGrc7pIOcx43aR4k6RV1Z9Nm4IbaUZYY9b0BEjg
cYqTEALe7VcaJ+AovqTtylpsNy9FapHfKHd17p3mgqGD8NPso90q9dhDqnuQqDZF
+pBHF5c/ZNrGX4cl0NnfE+qetIUnUad7pYM4KTbdXpTLrnrH5m9IcbhgdaitNsQy
Uudrds/fSofuTNmc6VYH8BWvofAoaVorENgd9+UIS6FCwlYzCn7P5wCQ4+RX+K/W
S9Aj26AE3lk6SzShj7p2JLU4ZlGvmqKn3bWSqu1ATMGGKHh2gfDluLSE92kBfwy2
qiS7JlgyjMIEHbvYGoK4SkjANDmdR6Q7TB40Kp2u+kQsLZTdcv659ti3HoWOBqMW
xz8srLNKEnwlOdP5sr/kbP/Tjw5+PD7jS5Q5EuKVWrljXDJ2B+7SyfRcI31Ntp46
4zbbU0hMB09cFDxrhMUR1XdH/Q3rjaGjs8qfN7COE8xdn261G5M/7TQ9e8MKjcHV
JAVogyT2PUxNlmciwk1zyAdd8zjFrHc6ADPvQlg9n2EdDvuRMIR0LG1M4RlJfEBg
6lTrOfa/GvtY37ShNvrP8FJ64D0HKDh+YoB+xwIzrHSzrbocanEH4PgqRFsrBRyU
bfgK7lDSTyQEqRMSwKdKoUB6mOs8GsfZ3GGFM8OORxHW5McCxNASd1hxkGdEi6lL
HShj4rktYE9uRKl8Guyjjcl+Zdg5MYuopf1sNwpG53hfctdwXBp8bCFCLLLjOtZa
54y/VE2/UlorPWiLilIDJqf2Eg5hlkv4Jv++VR1m4bdV1f+l1WV2Q49ljCcZSfRh
pHI6+teBlg9pLywk3lZggNL0SAKYBZjTf/Yn4qLwou33ySjUcqbuzdjYF5mDxdDp
xVzWWkfhoWj7MPXy9wPOv5RsNSV4J/3IRAkiu+yMyRj78Nf+bd7CA+mLErtCW3ms
iyMhgLMqM58czU0/BpOoiCr2u/gKzBHSdoh17X1BdAg4GFc3bBD9agBmJbC/Cdpe
NtTkFZq/tTfCVDRYo16Vz2MUtbQGbR9OhCh8wOhvamCaBKGzVEvWLk6awxJuJDPg
J1v34ChkgRkAVxeYiesYhTsDD+vqkqbbKDJQhOM64jh5T2WFT5X6/XmTBuGdTDQk
lBUT/XRxkxUaKvgP+BVBv+em+MAZ/jTgK3LcG8SZ1PECuiq5gB3IgzNI6VtHuhjQ
bObGA11ES8ut4hmv/Yg9ZhtbyZwKGJTK/8pVQI2u3KI+ZDCLALQyY94bkEN5Eiqe
bz1Gx+RdBimKKvb4qsnYILMXr4n4aiRvIO/RhkUR2vcpmcxl/5U5LqRomWCIsCEN
nlHrZgIhH19Pe+8CRe242QcBDGQstSneg1ljwi1k6YwVbNx+rg1sF6Hn44A7Dp09
0OJ2/bQXriUiSNdUqTyx62HI/fKNbQJ42aPynMHyJAFFgmh81fvqucl4B8zjEqsG
RSMsbhrCZzzzBE3Ar/kWcIWbmErZcmvLmZjfOClqgOQKGJY8A9bA8gG84YH7NTgF
nlQynCij205RLJd1JfxHg4H86SO7SXhTR9cgZYlQh3jaUoPF80bxK5Qov0K0UwsE
bqvKbJ4SPuWNjxsBKad0lqm7SlNpW+jtvjPPBc9MBWXBhQl7dn9catc+qsXgVgtB
hACT3TEHKVTVvUDohgQqr9ipj4SHWgQrZgO52SUvduMo1dfdmZk9kJkM660u0U74
djtVSxpva5YTJw+8BOHgivooNNGggp8X4XaOQ/sW3E8cmz0q17kx5xjdufVoHJ9j
qUqFslbOn0TR1eNSV819gxAcq7ISvFVGwpk4fOACOdHD2VilnLb2l2RkdP7WXw2H
0b651+FWLg+ex4S3aU8cXdzw7ef1TVVrZVSgmcQrebvBSVrNltoQ7NE9FiKr7CZm
z3eIbKhMBni6GLM8l0Fufy+8AHMgq91o5FL/xajtJ98OV7TxP71+L0JkrLiP9MtX
27uQqLxo/zg/zQWOIvanJYu+b1HKvab/ybQUabetwFv4GuGNyievjEdwhBTIqQ1N
6QgWNbmWyWsranY158cm2r/JJ1wJZeNepsNqHn6JBcOBt28o3USybyMTG6V6o650
aWSOWWEG6oEERWdgEA6vhgBGGCkuQsgGLpmMtarneO3naG6AFupowaaJGhZXB8/q
qQHZgJXiEfHroHYtTxTzSxTQxdPSeDPAIw1LMH7kE79mcevVAwAaiBMj1EQrOsFi
6LvdJrGWC9XnKEmq8jGIs3K2kYV2Ud7MLUPBE0T1rg9R0paX3VaTa2bu0hCScywn
UXLh8TXnIq67lioKTpVVmGKcac9jD1LAUP0UDFoz1UhqrJotWiE7A/NzLFMe/gmX
CwDoeKAqzj0SfLJuUNGKA4mkYjadg+wu3y/4hRh0hzvHA8S4XeKcgruzfUhIKEnm
J1x92KCRt+2DS5jyX+6f/LA0NFEzdEcdclojTl02/Q9NiFqqyFsOw+dJDlIuP4xz
0C5xcPxlqfKDqzLeECDS3mwHBM+smLdW6ceOPItFdNEzwN1FCJs5DzKt9der2gBE
8asuLLKJoacigZecDZPhRsllb85/8BanLzDeSJ+qjTWGiNAggaemWLm5gf3zM+rS
WmhaU7Irt7GJnEAgP+aSCGwC3xq0jQBBZR4gR50lpHtwIF7G+Aqw1TyIEId+taHl
+yBwUMCv7A2JGUHEUYUUInSpcGwvUzsdXV3TS1N0MgmUjJURAuobPMYeYo/EnesV
r9bd9CTtj6jv4Uof6bTZoFxKjE4+OmxJFZ12sd9XfCt9kdQwQJLoQMPD/sTD3K9w
sZaO01SGC3toSyGm2K8K1Fw2mBzq57aqRxuMpUbxJ4ovnOEkQvqp18wncfRUluRK
v4eDsddPQQqU16zp9yCOV12hGlh+z9+kiDVJK5CZkPjpDGHy/BZM4VP2TSiFDEAN
a1QnNlpyCjolr20pX1jlBH8qTll6Cyp3TaQXIokvdNlhdFbGZ/DXtPNGpSx3FgU3
Usf4EH+2TKVsuvGzArALV8pYNymf1l5PIdX+LFIe2bKSZhslvKjuc6fU7ekS+XRM
pz/HW9WL8kji62sJ1qta4YN93dvvXoJuiqWsce/9Bt0RHkG8ThYWQITLTqRUCHfX
Q8BBdYEJJUf/XQ6B9dKMloE4kye0NeKOBZPMgad+9+OXg00+IGLwmlLULXvTpg9V
t/wFJk/+MWQ8u8+F8bNhzokTqTHqvNyKX+PI9khfMi6PgouwCGifIakNL1LY5tnv
gAAatIloH7SdkyVt/FKaBqtYMWsefxoy31YFd+L3K9P3nV7EQ3cVtOrkh7AzRABy
A2M+EEbEwoLXW5X0Htg8pTol7cpNgCdBO6zg5kfKkpizgJ++EW3nLnnIzlW7XdHJ
DCJLCkzP+rr+sgK2nNdg9c2LEdloKgbsd+vdeBD8FNZy+zSLAw+k2dFUeLUQRtbI
Swck4hvjlB4+/0TUv/hwX5Zr+LuCkrOmDh81xL1wZRXkh3WOButR1hhIuhJ7ty9T
EnlbpU8YKbfk/gGrkU3LU91RwR1J6rHKkodHlcxyXNr3izL5VJ9arvByINuW81Nh
iPjiBCn0JoV9f8+Bd2zceHydRGbXUs6PeUiT4PgxS6xP9+vD3PjwA++gtmhCnt0I
RVNjcPmfE+KazM7rOC55NTSI6D5k9bi9HOm0/7C3EApp8bUtMp74D1dMonNub8WS
Fi83XU1D2PdpFYi6lnu6VQb9dW3tj6GhwnQRCZG71mQiWe8J3hzIm32hDyfdAuDx
OSptDegadhVzc4P0vaQP4E1TuAoMiPQ7e6kIUhawVE75//Qv6qURm6KAv2smmGmj
U1c1oiQRryXqPeV6x67raUvk8ePDl7BD4JuPRdaufbW+uaYanZ/iGFlNNTjctzb9
u/Cic23OwEU2km9omoHczZmdZemJDYyuk1ptS1pWSpTMfO5LPByuwAolSkosKGWN
5gNlus5MKXcoKJ846yrZKZlZmjUIH5A62/r3Pz64ssk3uA+19vE+J7Zhm5ijI8du
vaU5ClfQ4xgfnK+YwH+2DCbFVSZ9SSyX9UWTsSBQczOIts/9yS2N/mLv8jfma/Mx
6ltQ8+W9WGqG/7qBVdRGwjfej5OMGBvtPfG+MY6tbuHyJBApzHZ82oVjXFRUI/VR
R2+nILWf2SXhk5o+d/cfTuzabPb8CWznAAqOn5Y+ONUGBBjDa8Y3U2UVndRuE0V1
lBMWYOnzuNzJ1J9jYsnhXOPDqjiUP+WGmp3UcScMyHmSSuulSQjCC9gj2A3/5hEn
8DPmZ782me12S9PKtkbfpn8X0eAr2WdDWmPi9vR5B300OUkPUg+4WX6Z0uLiRAGu
TC0DTC/lztVvaCAkkE1OJvHZSgAk8+P1DfLu00lCkY0wnR6BVbw6rzcyCy8zFiDN
ZSCOYEFmjHYkWxGjVq92o7ApJHASeLBzOWbhGm22T/ZxMDI5x4LUHCXe1GMp6z/j
uGS5ha9ndyz07PuPqBIvAM1w/0D278H4LPhdk4nVhzz/3pT0uAwYqwx3b9kKLLlp
TgrLCYCEsTDv6W0xuMir5jYF6LVWJUQ9lt0tlz9PsB+VR2ukhhtTiukFh2zto9YZ
1+53gfAXV+doH/hubYVvYfGWV1TOcyZl5TvcWRjKLl6XON4Elw6onkrlQagTjImc
uxXWEh0jxX70AUqdz1b8j29hcmSIMr+NrfXuMeJCv8NnkBd82KQySF1edPBAwS1n
wcMtBHd0o/LJnuozMlOrjZq9ZKpneTKXBqnNKc+QxpvAuQtGnX6/mKvYTEpNuicf
+HkWGt2dRzDAVgguBib+6VZUAdSe6r9WTfe1j0HRHFoYNfsrBHQ7P0ZW7O0iCja/
lQAVXZMc3KVEX0zRtRn5ACqaaa62Hf+PYwScmIxweS1YR1UdQWcOKH9bJdP+WOxM
Is20PCYH3PPBPU43ZbrQm7rnKQFr/uCq8mpgR85fn+ITrJyGEK2ZNdQO+QKOr3w8
gZLp8I5slVfRp4cAYOtibfDxcgMSS5dqcJjSZZgL6KUyecL8yY1KqZi5I63Y6Ckf
fwpdcNUhOBctJNXY1wphzGTPczaNKm6u1PzX1qKzPn3DtCZFzBUWqGQssi5rRp38
dfGg8GcNgMSN1Kqz3EbuicHakThjZg8O2IZG1vGnQtnyUE4cH7cRUx0hWUk3BooD
OFFahCgrbDbOaDWz50EFDwdBMYijqzkZzEPkVsLrWViSHU6HuthcRHBM142iOWpc
MryxUEk4QG4Lf/e+D7jg/C6G4sf04jVxiHpPXHHyq2yHWACVAUCxxTtL91P1XpyS
AXsuW8iPcKcSSmcuGyomnwFpSK/UyaQ3orgiaO/I8AVZ21acbae9cVi5cwtRkL4u
RBrUQHqBsSKDbNXPXGh8pOcu24vaA2ePuFmzJah/8GuOudwDpaV3DKl7GdgSSwHw
iVmhqwAUO7yLeWL6nMqFcSF60zr0RnVNcXKxjRk6HeE2VXFvQbolHdCNlPiPEMgT
O4qYk8uaAz70CA1wccnmCwH0nkD7PphwbzcpyJrhIxhZ0jqA8w2Qyokf47+cP4A1
zNsFB+hb8e9C8BbLU4iBCrQVzqDwbHH/tHQ+wNUls0Zav5CUqKEQKhphP8odBlv7
aDn9Wz4S9b+LWrPaiW3fRUcdNslTnaorT2z3GB0qPpXFxGuQIWuq1/DX+7QmHCP7
HNMg/+HxbGpN8Wcm34BEiUtGiKWsJuISGWQYckhqhAkuRHAofFC/CbDoEQo0sd+9
xoYIIoIfUdyTB0xuA0y5dqwI5E1d8P+RrSJnGD7VvHT5P+qwLPt3B9IuTiwUK1Dh
KHXHv4J1oVM0005sFCLglmJWwDzTEgm0W48cIN34h/ekE9VZWOo2Bsuqgg7Auy2j
PDIeeUGQe7IM/AuHg0CX4s4ZOAqGF7192UnSVQAAQQ2DFA9pyVXEowpwFTmcA+U6
LNcD0CZKR41c3m9V9ujOOsLu4T1UNawg3J3VRYVVexMsITOkhc3aLesxcwz6SDZo
nijrt8t/PiTl1qCbjqm0Q0/JhXg3emY+nqNCtmydT744cz4CbBol7qAHJtX3d75A
9ONn/gFX8/HZ4oqafVDet54rvZEsRGUGrjjCkPCVRU8RW73xzhLJLepyj8zgzduR
7ZmnH1WI2bY30BuOAzSYFb+1WRiyLjJqDRxcZ+S1eGNx5uSrQyFCADnX7hIdmF53
hLr7Yevj/pXtyQh7fkcbpPpjpWiLRTdpdOq/KvnYQIADGGEuIv5Zs5aQuPxF+kiw
dPHd6rIl90W+MlX+ho1Z4qI5xNLaP7/4i1UNheThArkh11dFRKfPeNo65qHUX1xw
lIcBOviwxTw8lGxxXYNZoKGarkFeq6Zl/9WpZu7nqVp1kqcbC+N1DKfp00d4HY4g
M6jIiJUvK6Xd2fj/SHvVo6U5sGEfhCyOPRTYhfkhlJ3hbYmOUobp0JW/qMXE6Xzf
hr0XYS/jb8/B+KQYtunylOrVi/i6iHD1Bu1Aj+XKE1JXDDEm/Se3qL3flgGCCqmT
IaEPunBccubjtek3O+TqW3HFfMQf6xFy8y03+l82DdJva26Xb+q1j+qTqv74gCFK
86jFTxanU/zn80X2y8UUgT+05fD8rMx6PZQO0MGEYVlTCxQBuSymNxAAhoFWnHDg
FJQzfEMTFtc5H1VjXAsC9DB9hS6k+fx55XyVnge6a+zGXkQPUjukwYmWDHWfFYVS
0PnMOm4F0rSQGT5K1HAPCxeJSQErk0Vv3P+RwixQVDXeFhD7CA/nhm/Lh1yqqo0m
WOeOj8CYlGjLisM5lIh/gpmJR4fxz9Atx87R+Ow8ZZ7HO48+2Nn7HIaChsTxfJXG
ybVULhwd3uqRh42GCrs1yhMOdkoXksn+u/J+JmDfNrNwNy3wkwGrSSiZ73sMp/dr
QGmylIirsQkHOIs5eUrM1kPwgNrmPJnSCcAH+HHT6nG5LT9m9jV7uZ1Uci+S+Zwn
ZPUd4fZtv7UoRZMKnMfFVvZkPe1x6LcqpIfAIp5ZDnbgmuv8kd36bXggkpoUsv43
KUceP4cgZGpEGK/XnCROW+dw8z0co28MLiYu1kExTrgfXdWPR8gpP27HDVOzewSF
tTCjY0MU5ghIUMnfbWhRANs/LOLP5rtVUDkzNcSZOJqSV2GKn6302tvxtrbMOVLZ
hjsY8AnnxPEc89OHLLlnOsKDAANhi145yErAiT+wH2pgfLMFm7ApL8Om3hzKS1e5
wmf+Ov1wtBEMwsPxIj64Pldg5w4MrYMaVT/neUTXl8v7Nhkhl1aTEF1ThPuWfUR1
sAuNaxbPAY98ROsxd5ScnyTodmXh6FuC6kHU8SQruxGBo9ZheWGcXfkDIG+E+bN/
GMYdubj/pM2PEW2z1H2XTS/n4XjtR6c+c2jAzPHqFQ8g7sfPJrZg08BJsOe5h17B
Ad3UeKHoCgevKHkxtut08VTMPhJcWenb6fCl5fOK+UGEiL+URzvah07k6tu5y9Wr
pJiqU3exwrgtk5wA6sLAvKTeccKRWFb+LRF05TYflV03l1WcM11o1rXp3FOzOudA
+f5uduFN79vzXWq+ZmPBU572Nxc65Y0qxo0g7N6rpxyo0t/n/rqvFeHc9m2ZT3sb
+pZtWfBqEN2OJ8ZoUIy93eRB9tLhZcl71KxhTKc1TwV1ONeckUT/iMTNusigFeFU
JUlxejQrirSlnwvhFxJCPqbsWVuYnzj/IcwWAg1Qb5dh7YsRFJ7IzqTyCV2aaH1Z
G+E0iZXDA3+oFeZZdAjk+mEPP2KvW/oGf8Lxn4lcnX3eoN0rMrtN0J2ddqi5b6OV
0Qu6xoD+n/R8TbMcL69DJLrJItpMhIRyW+5WRoeSKzVUmHgqhloeLwkBJeAgWUf6
WH3QIrKINta95dqVKTJuUYchOXhbX2nRGwgeB0z9GTH8xHLmVRoCL5n3e/+hhCqX
t1UJzc5C/+Fqn+xRQCHn1a5GdU6sxEBt79hXoZnkrP+S44uk4+s/U53D3MVAGsA6
EG1faQujbF8XlKALBHr/Rsytl/8jz17M9LQcigDbq7SnmtDLZFKK6VkfvymuQYo6
efwQ7sn7Y+qIM7nPHqE8DXBqoT6LaDs+eFYvi4E2tm8NLyB4EbcQnHyi6n+joiiv
TC7Raf1k1SuHzY7EpK6Z7J9QFO5Dz2+m5RD2bv/TP5ekUZu/czVd0TmE024/eC6c
GDINGJn3FSaGq5yFc9cFT2VlWBHE0O5rmcUNeTqGmD/vxGkowdZd+RblyWzh7MRW
A+oVkYtJOz+TmUROYUOaqLKRxAnTDZ0qLHIM/Ecu1Z5W0iIx4GQqeB6a39vqlB6/
BkmKbe2B1eZjdJdHMhbZXi8RR5ezOWlNFH4jCDT+iC1scYazHhkffj5Mebvbe8uE
SWyQ+2JomAcCQcy62BC4UljgHpWgRpuIg+A1SYMqA0vW5GnC2TiCPZ9w/oeVMayG
x/tanDnuQ96UQ0uQpGyqP5soYZ9KvPBSUv2+Gc9+XaZnstb10x7zMBq3EvuDacs5
PEXdQE5vkabmIqpCGbc01GiVbXeCGsE4v6CN3UCCdk7x/Zj1MRam16/ITJNCfnET
3gsdGc/O4JoXGwKDGqYJk20vKRW9z0dDuelVnLVdgVzeFdqovp17zOW5oSEFl5RQ
5UJyl4QkcQv9ix0SbCdI9ltgrZQj6UN0VmNWlXGeLVmNaSKHyRViTdElP5i4lw7h
Ww/u9atwHBEuDL9g1eTJgsMTtImmkY4H4lXf2a4Z2Xwcvf5u4FJkLIFHZ6mWolV3
KUQdXcwarc+Q4Va1160JG7oSnfB7xvtu5YCtbGuk0zMxx3Yew0FIJi01SrdKBIJv
8RoPOaV9zoslDrhOCyJ4QFozQoxjDohLab7m2Go71MtQuD9ZmW/zNd7uTRkSLyF7
mlriIydKvtRjW3e0yWMyEK7+5/KIDYY6X2z3we3vDqGv4JC32cxbKdknVcwZmdSw
38oMh+PLjmIY3I8l16i5ww3L3pg84yaJBB18ckBu5NuW6fVAKvWoDPrCfDDB0heB
4KDg/9QKamR9Ux7dT4AGsUiz7oWQqSW+WiCHCvMKX8MtY5aEZ+lQzVqTTRwXhOK7
UGraznahWH1UHoJ+biEzBcDIbjZZzP4JWMYqsaJPrSk2e0JK8SFCCd9qMtY7MOaO
npLCFYSucZ/rZ+iCZks1dvHfQ4TK+KxwhFLz/Att65QGnbcmShHgs0OEF/m2bLz4
nt6giI2MVeT92u6RhoiJMIhUY17GfNejr+JDcjyUK8jZyZbUN9QkoVyFi1LiQFF7
1XpW0f4Ov/jcl/6NdXrvRcPRdg5Bp1iCrt72BCBzCNUAGokZIoibfk2QB37Ex6vM
aa96+b4+ZgueOM8edTBkfkXlw5XmrlciJvDL5/8/Vb0ARvF8LAti6n4JNJ7J6cTB
LHPp4pz1UfaOrOBgzRcWnx96LCu3AysAq2CE+6lK16PNXsNeY49QMweJhC2EhwJM
WNqlUQbxpenveqdxvEQYmzRm/shqjLQjWx2o8Y8jyo54LuvcpcQ4YbLo7NDl/+cw
8kjS/hQDxXX/I+B0SrX9iMKpt5Jm210UVG8FKu09UpBP1BsCJ1WFPo3AkRVVHqkp
bkvxBuK/95QX2xjmVDEW4VEqYTimpkLkP8tOcqhX+EmEQ8jYj3Q6JNV8vsKaJypP
+n5LTxms0JT49mTrSxjZJZlh0rRJc2x7afHl5AkI/wqsENIo1d9ODYWJJ6/3/PpU
4q2Vsga1Hy4NHy1UkL2coqWGHLbWKILrhTd2gu+yH3GvDAoGiS8EtNGrx3Yp5B2Y
XGBobpwLiBpim4NyjVdEXbvg0YwyTimXODXxCZDL36ngFq7ptdpFCOOOEzCGQ9gc
FYM7DNZoV6uo67Hwn+qmrCo5/Tj0xW3+Hn3nxZeyi0yfvIzERxs9bEio//etJXGf
Lme2EoTPxVe0D5IWVVzA8f2Si0gk/mC0mX7XcaHAFdbIzEc3fzYAU3bGLXy/fV+4
iV7KoGMZkuogpUqwVBThH2BUqaie2iYxnfjkHAumUQsnvMUd//8xhUL1gSkmPc/1
MtB2VdILAOJ+89/2w/WA+ybQ+Rpd0Z/rFvYzmK1Z1sGsiGHIoe/CQW2Jx1KjWwC8
UBRLY2M5JARqYOdry47n1cYkwcNiJzRteAJOIjqLjP/dexTgfQvkzVfe+PfhKZrA
1aAsbTjvLTw+MarFGF2dXOFoOQ5G4SW7a4FMe/E21E+zuCZvUgsMgg3B+6HO0tyt
eE0lGkxwv0cRfngRF/dUQGqd8DDNLb/d0ev2xgr66k4/J/Lrv1rIiWtsWkc40Ahu
pCv4T0dYeUzE5RbJzoRtBb1I/qIKLj1dE3vLk68xxnuuG4Io3EGu8DT0En3G+gyZ
LFMUEKr2GgyBI8H7L4c2adHcIRwIQx6La4t4DWm86HJ7KN0n2Jw/pfjp+82vnw8Y
OTnRrQ/foIGYH2gtp/6I4V7gP8w5hXzbmBOjH6cMkuTzeom4789zAFdbAFLpIZ8x
Cvm7lh/7OeeUBchk91QTYtANQ3jLSpsbjAD8N0oNYM5J6OQGpdQDDwFyhkS6vEQv
oocImrc4oMI2wVhLVkaLgYgi4aPFPSfIvtJLtsYXpUIkzoiHhbkrRLpgClR6aPew
skfRfXcFugKNpV4RNWePOb67Puz3/gpphQpwX4qXsADamBroxyKlz4fHpLgl7G4H
ChSI+iI4jQ1YGeG7lruycHEDn9IKSvczaksfq+1lp5pmndfNTpaXhd0ZNyM1aop4
nYA+g8vF6VsaaG2vdngRyNVicgasb6Lr9YgNMzTdQ3Hg+Md7KOxoJN82noJPLcAm
ZqYMeBYj4VJZpSXB+M+RITuBkREOIaUw0xa4f+d4T8prCLn5J5lAuH022LwVALXR
AqjoSw6RVW3ha+L0IVufwqMqVJ2BikJTCEHRZzNTWhgjfa6Bg9lzIzlWm4CGf+gR
SoHY4TmTnCk9om/tdNOe/T9TRO35JsPsxlAfJdDX37MuQMhkdRZTMqoW/tWfhNvt
2rCKNbkPZmJg8+lZB95n/rZpF5+7XxVCaDtfWsIBI8+OU+6LGMomsZ7cxtDbD2d1
FVVTUxFTXbfZ1DqWhAHlwmZ4vWDMxMGGwv3Z/+K0vCvvJ9k3Qh+l36yoJv7pbzNA
GDe5axzPxik3nS7V1V5sJK11CV/Kd7lSkhjnYY63yEiVrWcjfOoSgQJBo6ydD7tm
kuNy/FB4TfEsPN0+VbmEdj+u+uLkjx7LJy0AliDZNAt6f48Wws9boUzx/VD5L41g
DPN00hw6CNIzXLIrnlyoFQsrcItICas2dVWSJrpNtAxPiMlz8t8BSpPtfhSVHGJ1
BcHd900pcWptYPYJ2TWeDohadxT7XnqjKW9TvfZLPJQUoZ8yM2X90mrjuALFth2C
GqBaisUc4mmfhl6P3r1YZq01AfV8lgJlICE313kHxamnSLPAJycKxKlwugMmIFsm
qGYInQcyn67VexXcL21L2F8mvGA3FXRL+2yTRUGYAXH8yrwn/7V5Myw2WudNUm2O
a9BE4TngqALrkXcX1Xa46kbd7/JBtX/yMOOz1/2FMv5aWfctz8n+0GsI8jUJIqOg
J62/IzLKZMSQNoMuUxBlhuSbTebddfF8ybuPwt/YzsaAlu+cPwj5pPV4Li7mpAyC
It/bknqwQ90JGhLSnz3khZB+F8uhlCFyH9kJdKOV0NuQhFpa2f/uofjDhXNpbE7o
YhwDaqwHIARYLLXpkm73/EnvOtSZdEuKzPceQ8p0fHfvwODv5jPehdc17aEmKOen
GqCcj6OOKwy6YO+glcHqPNQXEcvFh1sRKGe8coN5k81TWU7sywZzy5FbhU1SJdDF
73qGOekwpdc4BRnUlp6Qsugvt3aeSl4EbZ30R/jnze2vEPlQvP3EJUdH1o4JdE/B
AUcduOHpi3dlyaVUoA1F+ZaVaeM5cln3Gs5TP9361deOHoJmCrgbcwM0wVrWVrYO
tyvE0r3+LTdBS+3ncAPvwLbMzcPX+XXOMkTzob70s9NnPcJfANuYwgqE1c+GiJZA
6Q1UPaO77ayqw5bHry3NoN6shPFGOVKas+52beTCC9aNIPsiyoc3rG7xG3PuKhAd
T17MS9uoKI6IdqtRjSODVSAdIrXwRsiNM1IkQRzuu6LIiyi3rXr69O1EtZnZn1HH
rdXZPRdvfMs3JF44Dtjq76S41+oLq4675InS9DdPNn/lEtzmUuv/T5KktscUw6AI
Io0tKZiTfBi7MY1Ul254ulaPj+huiqAPN7aGi8yPPT0xjFCwMhUKUZizG94ag0eH
cCPhkIcyLqF1zBa2NZgeNqWTbmyHiLEL1nROIS+yYyYAp7EPH6v3S4hEfw7s/7oX
03FXsKssUBKZEV5YQAdaKLNblCjVCi9DnF6rnFChEUbo8NGBt8X9v0+t1bV3aFP1
k9ExQmFTbO8hc4GlbaS+u+tJ8w3fUBwE4Tem3RMBJh5XOOQ7fU+vJqG5Rh3dQINs
X+6PVbt3T9bB7ixUQdMTDuHr2Fzj/WPGr35VAaSMzmlvClOvukDrxJYBzXbSHNSu
BxPIzhmd98qYPYPmGanHI0895qc2/yTiuAwrgjl5OefkzbMrdyZ/HHZHltjmoHAv
8Mm+rJJK4NFHi0DBP55HArsZl7JokcA4CRrZEGANK7lyT3fDLzjVG3AdBjt8YWVC
bWemXm7wk8tEnmQ6L3mxZsotd7UTGITFCZwP/UlbsNziSyb+wnQubE7p0S1vjjMf
Otovv6wjFSVVb9bEAj8VN8EU852p3o7cLNPA/8ZWqKxH1X9Dfc3czgas5XG6XWa/
xJhogkDbyRJpNhg6m0cMTxcEHixA3RoToex09wDBHjjHgN6/QHSLXNFpkhu7OqLR
6jGcIu4DjuCev9GWv1GBPPSypJ83K00YyaAjHtf0FPlSyS0mYptJyiLdMDJtXBbj
/nNYv9sO589APqQVhE+NEplJ2AfnWVqjETT2wgiy2MCB7GBiduAUn8cclkz7e2Rn
hLXeQahhZwIj5IJPVKp740foB43s7F6bcSu3xY2zV8dNZ/M4ACFMTjk9dHPLpSRV
ShL2FZWHMC/w+d+N1ViSI26OuBC0ewbItv+mSx+PexschUJVpsNYwCYqa8p5l4qP
O+bNZ1ztqA0rnoBGiwuloRzhnzvzLCVQQ+1PZF1fo++GPyG61SbypKZ6cIsKNQbB
ZzQRjyy3FdUC96GdtBVcb0ZK1S00e+0DFjcrrOi3pWBPcABSv1aN9MlrxOLETknw
FtiplcgzyerlQWUHBOu1gjIR16Ss6RELYt7m3XFriREf2qB+e60p4dE2VrpQbz0+
C9KFVJpu6s9O+gehraQYzrWDHom1+BnGETxRnjpDjVNMjqEg/WQqn0fqZxrVwZ1C
0tvqdXux8Lpsq3Kfwq4o3pvUftBelKQiO/fNwuqBlafSxO45YKWDGH5XYsYJ3k6O
66JZ4eHWvoZ/rIP7c/wXxeKwqufUk5E9CK766xwUQcNMlDi+tD99zdxb0hlG4ILw
qwwQEXiHaA1dcQi1A2sHvMQOfhNqwifC1NlEeQ+DNMYYFhgWOzNGbossdu9Ma6xI
v7H1t7KUt6XdHkxcAq1RYnKvayYdMtOOrX/6LX8s4BKUJBAqFlJfbd2JqYjr/FwI
0zNLX+TiTE56rHiT1NqsWL0GqcgA2bsQPgZvMIwY7PfgWSgfIQx26tJGg3Sf86wF
23OlNNYvRlhbwvT2iWywClNq7YbrzK/FQ+f5sgfnIPeM6OGwYFary/azCj+l/Cig
mpPIAsgNDuT1cPDnAnKGFr1txBtCzU24H/JLmqqmaTQBWf8crOK2625V71T6qRF0
8kPn7SpTxZpR73VwAvYRe5AYYJVv878dFBhSO/lIR7cCiX29+SJwF/7tgru78FoA
GD9IuIWAdCcKUqyZ4FxtEjPheOjX/fKjLaHyZ/2OsKLUV9T0e/0JKrT6UUc0M2VT
gmNs2cwoAfk2A2TyGNpGHlOBZ7htKe8nCrw1hA4MW3wUsvzhq7YPZ/a9rEKFTAJ7
q5W7DpIUHhnOFhEPcf8dEh8qcc6mGsV8EfwZKkovk7Lzj3wp2WyE2oxU8gJGzYHM
Fv9CPyr5Ql3qHhi641d3Nd6o4QiRa9zo/su3huhbgzAR7iA3WOiPBhsP3jbGCsCr
DdY+XSdmPCqZ9p56M+ma9XSZpNVr88ZTrq+VVg4R9GZgWic9DwglLpwgmBycFzlS
VjtYS3iRPp1zhTRqec5g3HcN4op4e0ru36qcE+tvscFn0kmVMimkOCkXGnuchN78
sp8N7WFXxKB+7+daYt+zydmGE2LDZOs9INtcA6FTta6CNDqmmNChwetk+WJzMkc0
kyx7Yn/cqXzSYKWauVjo3VekR55G21lUgOuwhfOMaFXdTLRm3p1SrboORWSymeSE
RpV7YHBSGy4PF2dYYREa3peNO8UoXUaNUtTRKjbdla8zEyF9mU7yCrAS7j8Zd1GA
fbXQ7a0bhiUhARuQMfjH+mHaVjDcojf1dgs7qOgpJ4aB4PbpD/hqt6kclGIs/4Jt
sEX33h65FTGjj709mlyMSQCtmybf/aFgnPFtGseK7w55jL0Hb7SCr1iBMCXTAxWv
cCwMnPaE+7wUztgx1k1Aeedn5qTZXnOkevA5fqQNUG2dw3MIpn7swz/JIjrWdDJa
n9FkFae6Yx0ASKkieOhNU7WaEyoEl6kLwIW7J9aefy7Lqz9LtOl3Eg0qwr2pWWoL
SrYjlakxvMpsyVxPaNhcjFdVHPq0L3XhGOocavMIGdoBatc6UhtUGNUZcDAILVde
bFTVmJgoU5eB9gfGmjWHnmEPijUwkRbkd8UvaZ0YX0FouT+j7C7VyQf1uSSDiElo
sMmuAjBiKXMAiKn22j8Mb4AOuKc+6lBw7SSpksJYY175UYQKZgWm4QGVsOJ/Y6c6
xl/uRjX99+JSJumc5/O9/VWagJnorNea0JSszQWOlQbaca331c6OOq4NTlT1SEre
cHR24mUCalb90X35iE6RwR6Vi4dmbDvsJ4xogiUwlKPPzKRoXN19zC9OAcjI8idG
zS0RRZxbWXWakq9uGvAUWXi0qkxAD00RbGr9i5bcZBcHO9WcSbjXyt4NpJZJde8P
/YVBjF+Kuhm+OjmWZP9erzvQc+KIG1clf/ddr+02wbH/i80w+WTuRBRlY1snuUJu
CAZrwDQRBHac1OS2DqqEW44s7+0Pbka0GP29cgdwpQWI6VYwx5beG0V/yHny7EZG
RF3mIUKDuAhp5ndNP1JbmAZMEZwWg6ytC0OMom5k1+lVh5cQB/6QcKVMyK9+jOE3
yOQbec7y0uMBkYEnJWBk5fSDAGsmbFGZL/aDsIN1kiWFuA23JpNtjg23/C+q4UWD
j85ymUGJ/E7Lkp0yUD22BfpzBPpp04Cq0R8v6hKLeQ7v0B2eKjGZpFW3hkK5gEZ8
W4nEx88QJy2bDUfreOIF8ODFYYkfMohrmFhTag4z+dkDzrTWaia1u2gRpY12om1n
jEbCJGn/PCUi+/+zFPMzGYsZq+tt03XwR0fqppUw0yB1Nqm6CRV4+r2WuWi8GsTB
fuNpg+Ucx1yQF9nXGpp7bOCTZNbJKiuGmkgipCCBV3FI5HFawpGjsR8FPUC68CFB
DGTG7hFT31q7sPM79Gncfh6QgSnwj5QyLEv60hkeCjFyfp35CSZxCiJDXLXQGACF
KRYCu17meQlOEGYPzcWBkIsp729BYYOQGyHyzP/PROHMEuyrE+1FIsZ/R+RwFKiP
E4G0ANYirRHBkPXxgGa1DBPy4/lxeYtHh7cBcMqfnej7ckXWMdWKzH3wuzm0scTd
/1LApDLbNgAO3nhjp0s3OkpCfmak67AsZAXpJcjobVGxgHA7eZ1z01WjVLwvLYGI
uZ7f1lonXUDiV7N6mkniaiJ1d3/av4LeKSN7ag+obswc37CYBxI/FQNfWlJbqSJx
IZJ2KqgDJ++8CySmun0js4la4fRFicbjGRdiR8dutfyFf3iGx35cMUfHjKjFu/Uz
lgsllKidwfEc25IohKDEY29uhhzGC915b8hn5SMebUkeGAK2tWMoRwhx+CeYxbpW
G20hoakO/ENUCc6dMZXzDMh2oDYZ0PMJy3ExF8Yiv/TmBg/p+G3ZrfX02G0uSYhV
+31XGBj2+tvrSCXQ2wnpmt2niP5Yz2xZHgEU2sV0ksStPAR1nYsSNca5pwvfh8vy
XkjtVjwVtXbmKW11Cny+Ey1ECYizGEyV4rOpcB3YEXdbBO++kO8s+RnUjzw5daHh
vikNnqlbPIcFCJ1fmkzxXcGTR/ys6f+2uLVwEwlGRidyIgjH6m+riiXp6MaF3mIA
e6784FSyA5OBaPzDxgMwQ0lKbqAaG8Zx6TpGd7luT3HuiOGP/9FbX147bS+BcVR/
dmIKSWKaE3BRHv9VYLGhciQROv8wtbRW60aK78dzFLGcM+D45suhIYBg1IC9zx6F
ghGirJZLtRNxgnqwUo/sRkfd8wiXa39FGA1CAyMBLqq3U6GVNjPfDzmDqm1Ng4X+
bSZzficRJu0vB9A9Psj71hbJRCcMArrO2ISOIo7/s+GJNfI1a/HUSJcijSCa5Jih
djl+L2Ux4WaHzT68szliS0w7df5u9uTNverKvj2kMd/nuJqLneyp1xJ5jWKQIJ4+
voKqAywSlMC41fTQUOzTh349uUu5eB6O3E6SfG/yGMODhDgPfiJO3qP2gCX+HL0n
0iJUVkPzwo7L/cDEu5+M2Z7JUfak425sQRpY0rzGL/g7es42aCGT6sRZb0Ay+PMv
fE35UpHpdn4/suKrS6VMIXOEqcGcoufyhKjCuR0aJYEkWsD8wfik2vAFYmxh3Fl7
xQxES4uJovi0Tlan80mEvErCJ3TWkaJVn6zSp5o0Dy0dOtBibiP6Oo9Ls/iN8oah
7JEKlPG9Z/x9BJfQkV4no7B1vCrBLHycBbyJQ05imkOY+DU58GK26VxAMo2Llm+E
e6OrDN4UoiapPwKGu3QxTpuOtkv0E6TDOu7cnGCR/T4VMP58NYAciXlrLBag53kq
slWTbASurDzjW0vVu9fmsBPwDbC5OFtB9Nrmx4uudcIhiqDADGbnPN8TF0wxsxUT
ssC5QhJS8dQAUlUEhEYT6nnvb22XBXb41crmLdlK0YQKZqx00MDKxAJ3d8wrq36s
DXqet4o0DUWiSU6Z0iAUpuVKfsk2nDo/WdfP1yrTx2Ol3j0AMhdmm3bonKViCoHn
G4Ip6+kDs0SAe4ERR454H1OzyDM6rRCl0gkjMjks81WaA9/yKAidQv8+D9btVyQh
ILL1kySDvL9wSLeT6jTbSyf24YGbDMUq+5FhV8YgcY2VLL+ZC5QqEpAwgZloaGTH
pL3eQXSjQR7QKZ20cY9Fhc1E1jJDToXd5QsYsWnG+y7iFFvIUoN0nCNzjle3WD1E
KY2e30EJx3uoRiv5wgUGSg7xxyRljXbWY4aMfLvYxZ7Q2NmtCZzxMpRHbGpXaJNq
VNOfTbCIwwvEaWfoEdhP282dy2J+cLsysdsfzhyM0EiYssJQL6uYdv+DQMM2bc/m
pTQ98azuYPccpcPOc0rJxwAHdXDtoTXV2RflgH9Fl+JizZGhDwiLwpy7ldRLIrb4
tH5pr4bI1Ja3Q34ny03nGm5DFPeo1pxW7YDQBUddLOfZndHqdD1906KXxzk+os4V
3dPp9qqOMno1LiR8RB9FGwQhdHlEAmhXMzTZ/UUVZ/h0/oFEIFbuD2nw6o9w0jRH
VzFUGivAvqLzmIl3ude/1BeV+rjkNBEIc5jHht6qedzjFl15E/a3ZjHf4Rss2pxx
jg6mF9+vklfLIQ+VAWsQc+sB5yrd7hXRQkgYlXXMpdYt9Ssos/4jTn2Fq6njh/ZW
xdGRdQR4geC/p/cSg10AQRaviwCWIoIlhUqWyMvp54A1QbPge8tLA7XHrJcOarft
Zis3RpaGfQfK83VM2E8t6OKRHrH2hA9oB1uWcnyctwDGoUdIFLs69b/vVJHGJ0XA
5FidXzfmm6LcMJa6HDrZq3g2y2ZCJZb74yy3VGj9jDi26KG/Pv7M9qHaegkvYn94
Wpn9uCqA5ZMJEAfv4ipD46gYUXnmyxBGMQ422nXZuja7N1lklhxXn7c97Tf/44Ar
/fejuCbtKwwMiEnke3xuouvB9gO7pD2MpTueqMYcgHxV78N8/qucHiJbUCqckKC1
3g0WhtuTrS1QeIkuHTAGz7Jw2IHaNXnFgHs4gLph5bb9c1XIp5aLQhzGtrytSV6K
Bk4elxzCV/7eSICmfK04xlovUOjLID7e+2rZJcDCv9uK6sIsAc6OWZZgPTooNKbg
BaqwL2B4uEweJq6Cvf45yKSOYcb5H4C+MtbMjo1b18vXI7Jl4FpwWmqAG2orz3sh
nP+6WEeTqmW3OZNYMNK9ubNp5/3HuGZvJ2KzSaE3lIjfYxbeMQIjqvhAxFDbyfxg
3dSiWOB/GCdm8Y7AicYIEXN0vhQJKa7/q50F9eWmvI5a6DUS3xih1xeIvGEALgEp
XyI4dKCJZdfS/mdTOmxpml4PjoKhPQM80l7f96XDPopVUx/823AOeYKpYmge4qCB
YhNU36yhtQBfB73ZnV4iW12eRTsJPJXiSBqizUHHxPS+Ys4vi/4ljA53RClTb/JU
0wAJ+Ct2VRbCz/wkhGGW95tM7+KH2cZGlWJ6Kr7jNp87WTcRBrTSkPhCv+sTwOUv
lCyokR1rCoukvO1Zic0K1Ro7hapIcYIuRkpiJeIStC80CDjTFlOthAX0qQbGD5FV
J1KwzRFOHqU9YneMVgNsjTZUP/f4BRe2vnxbfG42+bdkR3gngDAv8QYZiMYKfdjH
NJ7wnOPcfLM5oedTkVOouBpwET4heGU/OGWl6GgCE6YY9H07TweA0cOLWEi+I0uR
x+iOcPFq6go17q0b7ccfz+2RIOVJ5FUesb5lu/lSKTQpSsV5C80D9EmEpatbSwLG
aU95TyGVkhfy/gb0ZbQUjWTlRkzDfIzd82s6BF20FrxQPLHwF4wAD9wfoI8sCoXE
pDxgWAyGvNleUYewCtY/CpYIKA6OxCM+J9yIuhnCy7tM35X3xDCt+F0nm978mFXe
U+FgEmcg+nOxHlqs+5eAwVkG/A1lxGLa+9Yp1sKrhqyI0qnJkGHpaAMzTkjDm0SD
5S56+sGkuiA5IMoR8fTdr5DqCLKf1j6ClvBykN92+MuIHR6gkOF3/bLFN1gmz0mB
hKiyjiKc2K8rmZcv91zJPcuiqA92rPMNtv3KPuYSOU3vZCT7B5y8rMiYkJQtOgBA
DjNmiHoPUNtQDIHJqIFpM2W9HSeVjxsSq9y3NfPNvNLqdDYUSj5GGBoC0+EZsF3X
HukSrtnT9JTlJ1tm8E4mo8Y0T6qFgABoMf4dbJ+AxaYsG99dQ7IU8actPLIzMWqy
lqegu/bisO8DSd/ea6tzwzNyQW/z61lLIwgJh+C5yzgpcztXSR+cU4KjM9MJRIsA
eSmuzrY2ZeRMjquz9pBeBU47bQniGr6CNxtPkFH0bhpmfWN8vLh0C/82IHXViUx3
j8HGXBBBsgg2cZcZ02bPW5HcDbuRGeNiSQgIpEOnzvWvuFjh7kUN8jPeEmwchf5N
LcAokaCUhIH8rHIgUwPHNtv5c0vFQGWOioPgY+UrZpcfqeKJpKtlJoQ0vmZpnj2F
JBk6Ceey3wypyOYHLFLqQvk7L0KUN4WWSJNYuD9LepTLd2Z1ftjd8d16ryiI8SQy
lTeQR95GQQKhColKHOdHb6jeujTgr+nKH0iqGB+5DAFGsC7TqddGUXY30lPUZR4q
+arDETHMxNeXHCpqdzSboak392ducx6o7zJFZxszCX6Qapcc6VEXrmxtVYEULkAm
NYADn5bj8VYF4tDnOvmDa297ycwrdPRceScU7Y/sqX810btv0rT3JvQJ+zCIhcR4
X9ybsvhpndVh9JQO3jC5KcY8c21SOxaP5NyrDgbQF93r15Ql7UG5LSVlsRRL+CZx
zsza/bOlaxn4asQW0WN9WWmejSa/AF3ivBI8YJMiniY5X90YMoci9j/Hvu+bHlfK
E6jiMndvipdG8HFb/njA7Zbyl3m+XFn8T+azjSZ7MpOmYaakTV7K2GV49cECZo2G
Rtu0fOuGxUcBt6nemhuOYi4jk/Iv5HoebQJZPm082Z+/JgMWttX7PxUeBBUrXcdq
faNc7RZKnf8yXVeL8YsL5TrqyxUbKFQ/TyrH7fYlwkGsxHnIeyu/kpkbv/X27A3N
A2ZbHDCsLB31Unki47GF4EVQhInInKD8UzmHWShB1/Z4PZynlLs1qQRbXHXaP8OA
fpfIyGxHXDVQZ0t287P5oqmzxZBRs+aOJE6XFPOIhNDRpJQAzeo7dHRrXAyjiI3F
QFRapJCU+8BA+R2wGY/H3jqJjzvyQRoX6oz6ohfK4IXhxrkfK+CbwQ59qgErKQNI
EyBs2wfoelu0jfo8cv8pu66y1ZlwI9QWU6s0ZH+1nYhVc5H2bBtI62wqAxfby3f0
w2OMGN6Ue8F/rBfivLFbXOeyXSKIoltEBZziKMaeWU8z6Kb3mo7C1MT66o/XX3kw
b0PAsw5rVM6OfkCWiLrsBvqzvBF8ZqqKaDE/Uq2DFA1aXZ27iN8wKaODCNVWK5gM
ToB7dG7AmKK61HQ+q7OG/nt9piSwo2yk/tpAok/l1M3+pE/Jc/ps4Uf/Sgqwv2d7
mRFMbNvW4d11G9vt5QJh7XVAVLoCjB8FcjSg8kZHbWzn2qxvyOLTlpjUl2tsLMMT
xJZAtdJuXiymeSHRQ74MZStfkFzgIFviXBdXBc7Ot310kL1/vVxORa9dQDBM4aqV
PZQSP3Aomdu2AQzXxVqKwHvVJ8oCRzYo15sD8jH9GmKjFNzn3CQsZQ715Vm91rJh
iBJyrnqeZdLN6a9V2A/8VjJqiyaoL1goG3Swf0GlMeRHq9JNiWrVFy4Kg2mwzeq8
mcl/KS3zqTFMXcOncZuru9qXZ3zlGxCKJAUNjwRPXJ2cJZ35ieJyTDDoZSrocBIz
wcDd40VglyeIMzCJpO45NFdGPQroexMaZ7hvd4aNCBktU5+j8Kzvz1Dq1zQeWeQB
tHYlROlwFkWvIc3qNaHsFftAQTtPEq8/BaoDw0nypnnfs54B4fm1I/pbexlIxVEY
VkASL9QL+O764sI6DOXNIQYiBuFeSZ9VPJWSzB0KmWg0PBG2YUl6I8Ue+1pkCvKR
eErgCiAAMGky7rbQLfh8HFmvf88TbDsmyvgCD0wQE90fg1zqBuCc3vSY8D46fjIP
TuVnA3D10wYf+jW7F6oFJ2BIWX99jw4AvLAwnTKCeV9J5DgSFlgK4CSx7+HLtzyE
9bd+JF5+TZThmovpkZj3BUDRCsCcgfnvouhBeb6EocHrCZ0LuiWYt1Ob8D/61C33
ThacIwxqMZO9Nx6kd7xEDdQfT6u1uUcoAwb47Zaku3TiOO9pqvDygmlQon7/bPhK
a777MlABmPIuQ8SQBqABs7CTje7od0s+e988ih1CeR8Q0JPXjgOX4Rg1e5UBf4V5
vnAznqGHq1fgItfDOtCs+ADRjbAQGOxc6WerkawnWwbmcBUczn8rdKmWFF3cwEim
Kk5EHHoTv5xhMAyKW3Ev4b12sVZXbuFUO2XhGKsvKEGzDofj+dg5Z1929pBdzkMM
jQorpCsk3R5dBhF+aPr+/uQ334+9aLAmIN6uQdsmR/ld/GWZfryrqqqy7qTqcHMo
+KdopTpgvhzTIrVCzblPflzDsKaHIsfJiMEv1lRp+QdE42XdclGYzi2Q6oRLKohK
ZnWIdX5sbseJ5UmJPOuSHCr3U9qQR3B0MsaVeRc1Hr400IryXQx2LKrYbD12cK+b
5EDLR//wkSx0F2RmalU1LV0XTfa/nBcoHw/DK36ngKwckOhfBE/ydcgJuJsZkutz
bo8NWkhD56uN6Pvq6eQCNSQbFsLoVbGNkj6JXTjPBMzKhzICAuTer//8R0/FO+0q
+zi8NII9Cri1FiKV6lgZhTRsFuQygr+jOpitvhlTfuPjk0duAuIBj5aq2Z74Oywf
8PsNox6yP1AcHQjDfgW9EADghBt26GgfQKsth+taurgwvOclDEltABUDqj2HrNBB
7lVboIoEhiR0tGyXmR/HxQ/OJGrYhYRaKKWXtC40eVeLKLkYjhHz63atms1WTHK8
rldYOBjYCUrXIlgVG6X4d/lC5WiqyxcPLFOXfHSG+apJiR09Ime6jK5dPJU3d5Sp
bKPE5GUOfRhpSAcX2betYRUPr3c9nele53sJe3u+jf025BDIL5dDLQ0x6+wZizh7
K7hUMowwAf9b3DIDn4XahRB6s/j03u9nUFo2oAP+5ENQGRwyrp3pweWS5WlwGgqC
K+LFAPCNSzH/NNHv83VhEnKwUf6zc3ju26x8AI9tru2bDNfpqSY4JBGdlRgf7wYD
ATxLyRLkWCsxx5XwsSfsHV9QLCD1L3p/U7/Z6dzUW7PZ1+0h4i6r2g9IG/XDj1N8
jYN9A2WyQwVZmVs8buXVWL0Uo0u37mUWfyxdfXhxo8OCkPOASXqZJzHq42tRas2P
MxWq7jg0aR9MgxhoJbVIvfVJ8w6lE0KhKplK4jf98ziCCYlDt7e3O7pLGcf7g2jF
SDhaW01kdz0K+SGXIsSWItq7BfsZGzrDNEFyHrDdyXfC2UTKXFzIw6FFQSGA6dch
M8chRORVEfSU/xd7sUn+emZxn+iPAy7rVmiLo+S8wFcg9PiNCYfvuJ2ZPuUijxCC
/MmRM86HPq5d3TyYwYS5/uVuKp6qxvQ19k3HFwcZiOXCAJra6ICjJLv0ynYwIsqw
FdVkzIF1279/pmaH73xAlyZyZrgARlr3Lcqfl+CvWRzyyqLNl4R0ipg4hclJLC3b
Dq0rXLdvSYj5bU8Fl1qpXWq9wip4Wy2lOzaGqMBpqmzoSBigyO+Cuv7JI7ZiQ27L
VkeFembF8jIe2kFYviUr4nige8FDjnS7P2AITC6QgWgNEXrQF5ZihLZePQtBO9JD
WFST939cq35en6NHsPpBuJnZXEazLPHnSWL3YEnZGu+lbK4/pUnm1s2egHWSlpp5
1abaM4JuS59B9tnkj8Rggtoll1JXcUEPtN97I5LfSusl/nfYAwY9V2o26FJl+arn
v7oLVykOr+8c3pLY8cdfWWUSyl7rnB94Ote5MNy5HBE6LuHQhnnca5u3GONal0Sb
qxc6sq0xQpH1CXNMcGaqEHDCs1V61l4y++qkpJh8pGBiIxelluTUVRzPiaqBGYYj
CHJNWRWuTCvLn/eozkBftpVEA8GIUJufpoi/an03lzUljYbERgO9y6QffKXtPocL
hCSsM7yYm00Y06Hi7H6FPlzoHiZZZ7PgRcw8PNbUstJAFpdzE5T9DxJXag1P3daH
WWVyvAR+moCVmDQT/dCKd09lsLZkIYY8RxgVa2jyHn1vV6s4iNA1YDL+4rc6k/Ua
50/8uzV/ehp3ufH6Rrp8gChV/ml9IWeGI8ZnYRS0MPNoDSg7dKJZeukjWIsfE0px
fLoNwcV5qMM7b2d4PE4ZYRoTewsE+zkp6SHVCMsC5UWfe/aGH3wT4qB+3qrgXZyG
4IwVIYfhgK5D8UkicxgbLfG6+D/ffTrCsj+MBBx1lnkroY2YntS5PUQZXWz1sRzR
raTgWm03oaP6GYG7h9p8wSdJzDpnSvjaSCVxTERfL3Wy2C4psmbMZAZaDoalJ8oA
QJqb+Hvd32Fvv8G4j0lFdOMwAcs+WdgfaV9TdTxuimlroe3O1WoM4/KswqnMKC3Q
d/4H2bcmRkcSSBLZS0ZqManifJhWxp76zM4duRxzEfBHFwivWHsLKHIfNbGN8mjY
6zv7M8LjjSetBZGVHZs7/3iNYsZUUAj+51Ri6F2i0qZrAbOZb0HVAY1qWoK+wwPF
S+Lkkcsz1rncvTTUjFEcLDvJW253+NfCnf9xRELRmlZCcTX+9QZbsXsa6n/ut87k
hTwN9aFONfUm7VrpvrdAoEuBulY7KXMJc2a+hewn80u4aD0KBuIQu2KoPZuNPZ19
4xMkvvXalVPtIJ67CK00tMGdAZEnpmfm6ouK/S1Jz0S/0tZsDpxgB4+6Y16aG+np
yTIb/6aALRs4Ux0c7VYr5kPZYXzspSxsQfU0OlkvEFfpfkH4SJwa+q+80qciEFas
JPCNXvAhLlOmf4d9ZLO15DpN5cQXrLG7rAJfHnZ55AoS/ATy1TkgwbmCi3s+MIqO
XLEk3Iorze0t8ndH91J/xoNzCknm7Ao2sKGZHBr34l5SrxBUtt+ldw7qRsLr8Fgj
sByYH7lMUKmr1KB0bX4p8lltnbDV3bXiNIAMJmDgLawJwllW9zrpksWEQsjoKJ6v
VTZx1N0wNf1n0BInfy2pB3h8ywB5eHd9wqCb4GecqkUmTWhlkXIK2xdBXURbocfr
wb0JnzosfkT5fHTeJgiKJpFi5ooegPCUbEMf49i2oPpx9tnqCUlGuiYn+9ZAnFgG
IdmXka1pJeGjG8nv3+lXDHvuu70xEabomhiJg3QR9sDB4iCAnOlX5cafWm6QLKt+
n4uMDDWs1L8JSHsc9IWpjMRVRH+zdSEZ0ZUakMqNLrKKK+YmWjKCvu/q+aU9x157
Loxd+yyvf+g/+TcNiPimSuh1nJ8wPbSVqXXm5Dc4rnqe6Nf427y+UyV3qptaRaLk
9Ugg2sZq1HUi/9EeSJHcFj4TZZBlGyHaCavnqz/HjkgHkaHdGz/wCH4QBQjzPmQ8
jeypsUrdDP0Vzk3kDi+FTM7BgxBs13OK69Ongk7AitAT6MH+UlD3wrPaYNdwIjel
RJEMbBTbtQbtFGPYxfH4EaIHjd76zFamAJswWfxxjm2JCdhqpJ82wTQl4lh0zywM
/yFkmQTyGe+ozXS6E7xXCw9ECk2qgEaM5D7pladK2KMJXYx0nmsls9LRqwdwLaKg
3acqttTr6Hm2gXNSTh1d9NJ29y5XLYnbJxkTFrIhDcQD5eCmHgCcWDbI+VTrAK3t
2Lqz38+t5lkv8JDXMzJoBGA9bQnsovQyW38adcDfbqCWqZMBcjMsoorMGCZmN/GE
YOwhqDJwA/kWjEqw73lsPbq1DuKm/UlYe6FfNXfVNzAFub3LlyU6zZ53kYr3XByz
eyhcSyDvjUCV8SeMjwXtE4DbTxziXVWjVdHXRtVMdpisLPT0T1nbM/4/htsgKmI1
cd7hIIobD5SWZTGxKSQKSdIUiQJ8xTB1pKWfaFakSBzrPaFdySqRWz5mb+X4Iw37
eqjqkJxegbV8WKz3YzpwoqcxGwMO2g0z5amlaW0xcxsCxgoiEJj7AIQF4EMCjO/4
csOP+PRncCVUAC3UGuYq6k2Dn6IpcSKCaryzw5youbeIwxRC4EenhE5Cac9tf6ce
r/bPuhC4o5pNJUlE53Mg+eDF+e7W7zEv4IGZHvv4DbvSgVoofzYP5VHaNlQiyYbe
1ZIfKC009r7IkjX2lm3gNppM5feWN4FRZxp5TglE/+EL0rsMdg5wa9UHX5wyWE1E
VXBokkk9kBxSvueGI67cWv3AQijSu/TpehRx4gsb4Z1fyXm4FFw7w0eVZTspifh+
2rBnkJNxwqQSNOgIwnbwnaH9KpgpP+qrmkrxEvbzoD2h7J/Gh2GzlcCWsevI0tIC
FMwPliTetKfEj3V46OF5HyDnmNGP6kXPb2ME79AuA65/2eKlB84fE2v+cYNh9hJr
ZN9/8F+CBApLQ+A3oGFXy4kQH1HX3HhazFlQe7BRlMcsnAgnsnJjh5pg3OJIEiIL
2Xk/4OmFvWkkJCbp6FiEx3H9MoMu/noZiUIsZN2W2a0GTRglMbnaQ3v0Xk2ES0ro
lt5nY1poDeuUHdszQrh48tTMpHv63U7JBRFEQ8kKpd1g9QbxQCDnS3+/CSJ4uyJZ
MZR282SmFNuF51VA/XfbzmjbSSpndlax+FRBqLMlvPqxXgn2Qj5/nuBeeRIolcXo
2j5y8D/RrV+WA6WmXQ7UnJWNn07UHCxChPhZTCfwAJJ8ADlaglycCLcrw97oC75l
ZMShL8eTe9HZ3a4sFmZnu003pWC+zzmbav/20edCCa1BFNp6Pq8QhJUT5J8gd0/N
4AT/0VPzQVEEcIrwlGjHbEEv1jpkdlIEgozx1zqpZqIxgQXZH3BF4opu0qqQvrPU
8qr5juCMHUD1/kqknugsCv0bFaL/iwUjImP3vduTq4JIjSCB3IS4l27ezB0MHsM7
Yv0rF/8uauW1YWMlmz/cdCOjfcVO927qoH/1WK6gM8XPVD0sfOMwgr8lgu7aV+ss
iB+p9yIzDplIux+1awwAS8uYEApf1naloB65wLQDq7ko+MgYZtwjZ3aEesGuN3Xs
X/aSwLx7sFTCHoNWu0eLDUOqlK0rRFbjO6vA6BIZWNEOguxOsd92bpo+a6yvuZK6
6CTM8hgovYdrugX8Wg2W59LOAV3EJYJc+CiWkOyJpAjID7h6scIfQ91kKPwrqPUc
MOqlMDmM9ck4GbUBAdqu6hqN8iVg3lGS9F2VaZzulaFy715LR8+3+IYa6G24Ycqy
qz1fa1B1EcLwjPF8P4P2rkps5cz7u5MSgnFZTxqqaGfFoFFJaDZ/JKNeTILYuf8b
tiDWRtWr7BNK5MuGinl3VB86hPcJg4QbnprM3NjdtjIlzI1eRpFfQHKD5LZHs1yf
PbjXsVblPGKP8vVqqDDAjaf+ZOTWBIkgZ02hUZgEQKkeyGtAvPF599CkgIK20nBP
gG4wIgp7HjS7KDreJu7771EZ+YrLKhuCLwJ0Ygs7+y7OQOO01t9LNwrxfre1BszR
RYi2+xsO4iwfffozh0hsydU8SuKFH1uOHCsj6fCOESOEuLF7tx/24QhaCxMAMmpW
rjhbVw+lx1t4EC/BrZ0byGqO9hiJZXpX8gi/YZHUpbh3UivkB01aPDYnoI63kwWk
eRdnMoi0dozMefiOQxlAb3ulPz0ERTevwPNYm0Tn3OGownse2edtY5GOQfmzqzRw
emyNWp7LfQ/CjxsYfBB2mqdRVpWQP0a/EcjLj3dTa/liOMsQIkFGego7xLhoEP7L
CBJ+Lur8mf4Y0K00eb6Hvs7+cEs5QpDj/Vs1W1tFIF3ZIIF+DpS+QqfYftA/8Mpe
skx9n8TuPJPE7q0yS9ntSYQStfdw31AeSa1hjghHPn2G7Mo0Psjd7yhn9QGBcM73
Hk+SmFGpPPlYjOB5G4iDUNNTthf1dpU5hGpKSrRQ7ClYia7oSTUC1tH8u4ZCsE1E
iRr8DM+btLy9IO5A/BD+1BrChpeyx87Bz7z+0JKWq41qMnzcBMrQIHrI5PjJ0tfQ
Jts2db81LzPdf4l01SyG4+oVDR7am7gCOzq7Vc5esAaZPTKGmvonfU01nqjhtXbH
QokEdMC4JtTSoAUBft3LVLkTIjX+u1GefsFGYVlcCeqx5wjKUvtczkhHjBS3j8KI
PPDS0urB7/0wdTEttR0dGaBiPU0mO+6s9+ZcxgGtvfHnNiJG90szGMdQAR/Z2o4z
DZQdy8d8aXSFntmoZ5GmEqZI9tNA0Z5mYzHkgFNA1znzYRAaWzdRf/PoJs5bsfhn
nyyFLuqxMWpijAdn2/CD2Q9bLvwuDoSjy42ydHEkWZEMNlWeq9BVqtRGEzmvccXU
EOslIrA6q3PaFi6cKmpZM6i962gY4TJ6RomUZSFADFUnbYJNpO1TIveCPuz6CUZN
9U6SeNR7eyZKqfpT22Wu92W8Xda/fdibenrUuWsORUYPkrNg50+1DOb2AhKN8FrF
Oc815WY1zj9LewRJKxFPNmOf4eSkvZ+rS/zzZcZEKVGlTNKrZ5KptAFlBiqNdXXT
klAwESquo5rQxO6YD0xO1u0OrdMGBW9CMnun7fMt/W6agbUu+AEAe+wumHsmbOCG
nZt0AyqKKcXN3Qt2VxObuq5ZRwRIcmRWiRh/FCzwUXbOF30kZq2u9RiYNN/FN1hT
7zsSaiIZZXbHvU1rr7LhZ40mNiDY9uKe2n5Gj0QxmpISygefQuHlNC4h3R1IfAPs
XDS3RrdgDGWzMPtNzyyKTYKGyVB7ICgmf2mciuGm0dtbaqmze/VG3MNw7G/qS668
XeokSgCVt7LS5JFpGmqWH6nBiaYb1Fcy37UWkysW338hZuyEBHQzOP/hqTXIkYVh
k9ujfg5VULf7g10Sb3HU+WvERY7XiZhS5wF/suc9Q/8LfGQ0Df05+xUaz07zUv+W
/KfeHNa2EcB7R9SM37Bzbxhp/GV44HQCFhUrSMky1DlFCt+jxx0jyRPdP5bEiNPY
RAYjE7SsmlZZ663IsYysiy2wrgSWm2QIdqYz+2liQiPXIb8ZCsrVUISOEQOm8VUL
wSzi2VCXO+sT3cnqgFhf8mPjOaYftqgcp/P6Y5fDttgqW9aZ5nPQpuMApBDVFQhV
Ly7djm4iiKC0n7E54XCHQbh0zG0acWK5IcVOg3dwS+u0GJV5BH55jKXQmwx7aNEF
ye//9/i+hmuK3CmA02z8g4jzKLukRjW9Tf9sxAN1Sqlsjl6um+nIlVptQNRsvRcX
ysyiNoky0pXf+g3BmScUbvXAE49iLoDDs7XMeScF4AhZYsy2OjH+gRYQirzEOw9M
wHaiyH1IaBZu+7jK/heUxyZ+EyO6e7c0MNXN6FVqGfNuMmeJ+JmxMbgIMqCb+V73
q4KQYWEOQ1UsQ1Ec/0TFKUQPDkcKDq5xtz5rnl39AF/p0WsHohOP1njlkYEYmqlG
rzv6xY6mDdvfJMiXehEB/Vcjw6haK/hfTK3XWmhQnIJSjnIf9s0JtIAWNV1+D/wd
K3p/m8VyuRX2vV3BwRl+X06C4mNEoe6NffEJ/5UnyOGv967Wa/hVNHZE41mZ2Q4w
f5UC2nVe/j3gjJkShIbkprbEIRRCh7K2WJAdb8Q1hAWMxRK6EpG2qt6aHaEWyKqT
DNcZPDbnJcfwAWI3VUEXUR39TTMN463+T9b4kIg/NJSES4wWtIAlUF5SMn3XZYKg
sR0MqeM5d6P0Jw5lpM11dMx/oJL3niC3/LPi5PLV1G32EyVSKLrJpmMKcpMMTXs2
TPJEQ3dz2eFkcNfEHt03Wex7hiicSaFZ+MAkJqF/Hqi/ysvCcI6uLGfh8biSYJd6
ovr8DB/PaFFg++j5gtbBFe4PNu/7PDoWHYfAJ+ct7uQFadu+1XN0PKHZlnCzHiLW
8DFzS4iKVavIE6Vksuq2/oygeW4EyeYuwdiofo8g575WDaq/SgsmwHaos6dbO5FT
VfH19MrJSTXbV1oeLt68Mu9/flCZcWLY/KpEWd8AYDZXWaFxmPZabMYBMPg3JOl+
0cayJ/jpJkV8LVozCc1pqVyBtn9asNAqAyaOfGxzaJyS//FL5Qpnf/oh+jtM0Evp
gQ5TeZX6rZHHKrIqt3xnx9As00hPcQTbZpHezgV+utscxqngkqyxkcqWemje5Ayd
EWtkbxlJxAG9ieZHHyUMDrITapP4SlpSDRLyy4LVKqemz9pQM0mOO9f3jHQZ8lTl
clzymlS2JtuV3J2SaCG5BeH5UQkskZcMeZ87xydYbL0ABPEjfLn4TUDagkHodkDU
Eq4x1CdYQjy5obRm/aK0Lh0P89wfQW7Yo+KXOov2veUd3GFxVudlj8C9eBJPgydC
gGQv7b3Tsw+jk3O+M6P1eZ+Oy6Fq7NyQ3QXHwr2rEIxUq3rBRYvrIY114Jxjl9zz
IJOr4UeFijin/LF4NwQlTsyMnTgEGn2bsReqAOemdvIyV2waZRvEgxPIVamIuCn8
qotILJLJejPRs8njWn36B/OUtLMjVOM0SgFS+vNN9aK3E6ufLcICaNLyd5hfWQZW
cWEgloUSFtyPUULhacigPgaD+5NpEQMFuo5lRwbmExgiLGHUyyFRkNlwZYTMLLgo
3VD/01To3sq58iG+TVAkabVAf827VjHKBlSMiCjjGlPx8dHMY5W02hc97yV3rBH8
2DWzBeLCnsubkf0J0i9Ea02nuxc+dl9bL6gdZWUfF//i7+j8FK1n2Qg0Q18/RSo5
su5GmJjPHJdPDRv6iEZVrwcUpMBG7uhjO5T+5cidR1AzlBpLa4RvThCuAiOIh2kS
TcZaQtj40Kynz/nFX2k5Mf76oCi+ASx2HcqNMu8yVRVo8oTf/wCdgxRcrQMyGhJy
hgHO+ctaF7ChIFTmjHMc8WQXcKrK9Q1GvxvQjrlkCeJ5FN8IYYoaT+kPr9elRho8
te8V1xjkjdOOLJfWXcvZqggnijAI6dXJa327yYdJdnLrevF5rJn2vZoAQw2qGbeL
i+/WntBbVNu3K0pdoE876juRFOUAspffNdIHxnW+rb1BCWvRIsoXa11uCQTCgF0u
M6NecFTtumRD0I8H0QfcsoKRlCKlKzip5QOV6FwSu7yjlE40rgmJDCHUaWgNhZoz
qReT9HrPwfMgvSttCYlNyHoX7PsQ9/vkIBu7W8jJhv8Akco62ad2av6eOYKFEBaA
3+8qJLF9cwxm6yaL1KTf3rD7lzM9h7Lyawf7V0bx6hZ96KaSq8JB+66bmKahczV8
hcj74tthB30A2l8VrMcq1K09SFY2+tg5aH+xjknaWbyDhfePRsbZDBlSyGltS8X0
XxyQ3/sM7rHK0mfdSuyOreFc443jiW/0qbvQX1j6ZTO4O6hcAIRu2MmYzMhNLNHm
wfuCgza3mMX1YfjesMg3GmgclTdYDmF0tR9tpV7MsA8tOHmJIQDFEJMzjGwzFMgI
RuzpfTsRh51Sr8MSal8/BGzfd5cQ8JbLBoYWZTLk25DFt3G5L1pGBwXe9QqU50Qv
HNp7/EICq+SgCqGMhSG1KclB5WpoESXnRnnpWtzkYmzou+HyslKwoTuxhr8cLgMX
IXBNuH22Xjb9N1RSKqFmk3z9ww4E8F874tcqazQVK55V8sYzXbga4BESZH7cNuvw
20T3HPbo/vANtzEPwGSpZsotXQJDX1Pn4u/Nyi2Hd6VrCQu7ODq45KQOnumtAvMe
PfaPieNCoMwUp08d7h25K2WMv8uQ+msp+7gKrrVyBqObCEONYBrSR3F0og5DyshI
6eQtMIYwH7QZ3QN1ClU3RrBSYchobuMCOprwT4snbHomOVzqz2zPrCrxvIvS1sVT
DKjni5p7yuFw/GCEknTknvd/8Gp2cf5bnZIDUci0gvqsjYR4g3dAP50EseAcoqZA
cj/gmpVbEgrN8jBA0XaYWdV4ireRG2cOdJ/42Kh+urgmJyRagT6k/JsD5KT0CsO1
FKcnXWpfuGQiUaLJbdfc+PdnMnbMpOurwalCsgJTXc44KknIJ0HgL549kK+rWy8N
Deh5vJarC+6ejFBZGcUEbGTm7a0DGhv3Js7MS4GbiWdfEjVTEqOWiwNOP/6+ZiPD
tJIbx0KLPl7akKi8Ap5/hhwU2sYwAr9hvp8WYUVfLykBfaR+5mNgjY2FTsdDKYyo
a7vDVfMUcnX7fC9+FEw68s+hgy0qnl/KLL8i/PV2a2GJimuETrFsA4giSDYo26R8
d3oY1FyPOUFgsLzOEE4BSG4SXrf/9XuNUbMUIjsA4KeE4AnySlfr3CiIIJAd8fan
f4qmDu+CQctzyC1BfvLhL/wpRcEryyoQZ3hzG/O2KKHj0SVO9YSAcm5hlRPzlfCT
RDJuv3davTi7RvzJVh9q1GTBcEVfSxi9dEHXG07SPv4Uabv3F184xQLPDTIbTVhM
VzrU7micQeCJj7OPSdbFlvYVyCYpIruzXhPBuh1VDpeeaJND6kCTqEIcxYJaVqKc
L2sqf0mxl0J9rmmCD1PT9ssquviLwmqH827K7y6AkTZALyRx2/lgmoARL8E1tQH2
g1Bdd+//MSzXWV1a6cJ7EkRDkm1yLOF8wyy06MvcKu5idnjCNRNtfMPqnXv028VY
By+jpV/87no2rn2rWKT0mTqtj0BIq8l8DzV/vBxiv37aEhUrwbJQtn+3G+lzzgh/
77PuTPTJ5YmyLl5py9VITLxf+wf52Q/mwLBfQS9eOqjYjRww3xX4nXNLDa8QL+3N
CiG5xI0A4Iy961nBTdPp3Jz5etDF4R59UsF4VIgginGVl1fGmFKoxhKCJX1axZbA
R0fCP0bWI+4IYPDIzF6I0VEryIVoZgABiBqBWU280/CbaZpQYLq9jKt7UmUhF/mW
W+zoxvcRRXz6u9bUTo/3b9FtHc05gW0SD+cPhOoHQrS3QPp7j6qrXmy5cZOdOEMW
VErFQA7vUH87OqLWHVrdud0ZhHlYvi34wqyceLZmVeeWu+zrjm5RI1tj2VX1MA2D
invGH3oisfPTg8hbkU9/izU26z0KsWt50LC4b9qm4QtvOo+k4qXlf9VWIibO/DaL
X5AY7qIHtX3+Ld4HfUElK22CtChwTtZDtt2/zPaAf08FgAZeYfUrMxzwi0T6FSPI
9On+kbVnI0vCeQO1LigzapwLaQ22k1kxHr0Sf0bn9LIuHkp4jcluO8kcMrKu7Pu1
gvLHzi0B50K6bVtX4nbDgVk73NGpfD33lelPRLqrUFuve1ZvYTS6agtHCrlOEImO
S7/fXd6ZISAjWASoeIosKD7+f/k+zUlf9NX/TVATIGbsJphp+ZbGh+NLnpsyICz6
pAq7muZyTqhlAPM4S8iSPzBBczZ68VyM/BGs+CFlueNeZL33Zephh+cwazzl0pvu
d7SW2yLv7WPYUYa2PBU214tijl9OxVT+BAKnKVKgYBFgo/nmXuyssM8vWsuTplzx
xTNQPvT8z6S7zGVeVQkrHpxK476bb9a7cY8sEny7UO8Z16Tf6okLhNQF+1KZLQu3
zft3lfmuRJM/CownjFJkw4snief7aLlUOO+lo8UcV35oRdAuXlqUuY61ltJ8x427
/AMEY2YVceTZkCp/m1Ya0t+2YAc8xncNGbfIzwp7mESOJc8FEb9KjNQleWpw+c2I
sD1U1nBnwXEITCJmuvdaFrVmZ8/tjmEkZFko28VgCnA3XuNqWkdEs5cJAbPWytzP
uDBhdbNbOxazpbTmRhh/A/QLEu+BJi2A2dx4BxB3wF1aGCixpQBjhiB3a2qaKobF
YZCfNxl+5aJRXMROY0KiSelFRVPqFwcIV7T7YbUiQfV5nWlNEyhAJ1Xnk6aExJmr
ioP/RLYembpp1+F1yoz3v90IXiWtnUeVTJsAPh6VNLKNKO4no5EJboxg47ILV14Y
qw3ZXfKiNP/Gj8C374cHje/MEIr2CqskttGNULSUSDwPT5U76zUY53syjNU94Pug
GmNUKx2i94mh4HedlfqYBoSIeSGWAUY2JF0kWg564/rdJZBfxQANeIaUQC2Eny0A
hSs2/w/lF5AKbYyfbOxUuR4mhEMBXLA/fBDqRq1ii2L9PJSQwmb0T9Bs/5lVFSXi
oAN/KuMTzKe+V7D4vwckcMGloRwdB4whRvXn0Vq4vF37+0yB4va1qqZ3WZReKCw6
/mX5qewnuzAbZmpVMSe19t+Evd2kqBOy5/afpy43ORMhQEP7F3h6ggenwJ+Vn4II
/b2aq+14kS88CfqumiH+udacETQ+ZIpwmee2I1aJn5dLmUoe8Nd/DTNr3JxkcDhd
Brphh6PJZHgwYrmCig5j7mSeBoo0jNiTnU83XMx4wb2Q4hmiQGBmsxOzW7E7y3kv
g0KTX+Cl8ZsjBM9aSb9jxwI0q9cdQFSCKWSmtL/CreTXh3Ut3JAAyoT95QQ3VpVA
SEY00tHp+N+w+KN23mjz614TC4JRknfCW/6yg0vXE4yAlE3y8avVjwYEqWbczW9b
AjTSGu4R51QbTPtdDGD9MRKsyrfLWWFivpL7W6nkg7eJ3PQUE4zOO4/1aFIxcql+
IsUglYxnQW4BEBvt9geRkHK7EO8KlhtL0mT2YZHiW/VNSmJu0vti3wNIcQk34nK/
M9s5oasoK8XnBfvG7SNmiFGtC8RKMLoPxLD3XMjeb1z0kC7RUirDUgdbfLE3uhOd
Ns0qjVqt9KUe/K9l5aYNgD2Xc+c6c+gTc5rPwpQab22sYEpgK3e5v6ragP5L1pPX
aCl/Soudwv05/GpS7ptdyCX5DZCjYz1Vb40UsiM/rpwdBP/3mmz76VgJrpqIskw9
Tg3LsV+g9X6yt5Kj+C08OLspVfVXxIopjVb3vvRB1j66BN11SgTD2ZALM02BNRnB
d7cuGnBImxbnwEfith8IV2ofM/Qgp6wY+OeaXzaST68XWCh080Yd1fZ4pR4I30j5
HLqCaSrEtucmYWMtivK0ESnQgyuwtgF4+j5gAGr5GauQ5ovvCbMlNTgPg3SKUG6C
rX1HrlXaTeA4S+5BjuDxSe5846wDWYc5S07euIf065ewdZVHS2IAwFaaQ7yLP3o7
2jbfgD10SpafOnHEGuYp/Oe8GydvqErtXOpN8LZRZODzOtf9L/jeZGWjomPiYBx3
lorasYTMeZpTAxHq6xyVtPnNeB6qsTpwzy7qBcKTWQ6Qvre8bxoTS/o+kFEMwkIU
BuLWKFUcYcQ62IO72u3J141TwIkYKhBu8gOlKpjwm/XECUzF5taYePSphJGmAbCR
Pkh3zKg6qd6Nn1cENx5uubnTY4IFiWcrt9ThrCI4sGmNG14NgXcj5jj8rhhmpjxb
g/4qk5CFPeThUc0PXaWmG30eYa10DLhIJOl1F4L43D86zTTu4uMMeq4E27X0amLx
jrX1LWkCRSMucgTyMkKSvag3304WSN8x60WoL1T8RQAfc4NqfJq63rnxqiTM43P1
r/8aboeYYrbEQpXnSxGwTvMKQ0SWrp3TYvLb6l+ZRzPs//RTEYNVywoXK09yCIUb
pkR6o/jfwQBkisZB3wAONmGTirLhCkH4sg6SUelwu7D6eSd3DGVDD9u6GPf7em4E
i72NtxxfTMUjQ7rNfWfLoEosaS42lR9AiuU7rfLpCmvGVLQMzxly1ZvvdaH3l16E
2k3WYbYshOMVHvhu9nlSy5jrhomTpxTvZVFPxN14maoiKEekX2FEFbE4c6sunL66
i2mTF+JlHyWUiODTEXpJ4yfVAH3jx8TfB7wnjjQcVTvx+ynj1EAFhNak6E0m+zDd
XbIgAQ0iAwehw87bW2i7LN2jtmJHnNKWGAoXi/e1GkFJX619BCYVOBaYh10FY7pZ
MTBbVEeaxYzjiGheuQf/ygvykalLcnCfziT9j6hbpP7kScWVWYGUDjSpaQEKtHKA
OHRhlaa+XIqCLaOAN5wIYsWxHfdkjqlAxXDGsUWMd7zfibUJEqXSi3UdDfkaiYWf
kZGwJv9nzUJgQAV4Ex65gVPcHIbg6srQj6zbUPaI3gXEdsMgqABkbSyYGbQtwj4X
mZvVTUcPleWXHgD0szyIv/59Gop1NfrEqVevr2DG/uDp0oRbA7+tZqML3EmAMgmF
YfKGpAH6c4QWOS1g7kykUdLMYNTTkugXQ2tj2Iv4ryzlgsUoY0/fW+dRI7UU26aD
jEF6zTSX64baL1BMpesaY3/1HgD01S0Vr3VdqlcfAgKZDrFKZesY/gDIaU0oIyOi
mgT6SXuyKwJywi184IbQrcZ1Z00KWJtJ0uUR7Ap0vL2JzdHERU5YIXHzWidiYSPb
EU3fMcKjmriCIW1Lhhq4dgWiDWBZpzE1XvyKTGcwiw00uA0HBWgllu7DXbN1Em2q
c91fVohe4TP++MhijM2yqcaYilLPnSp39MCviy4bbhfYQFS6f/S9fhK3PspAqQU4
2BUY96y6U1QQ8W+yG2+slPvWN6KCB/Kt5iyWp4L7RZUS9HTI1sVwLir8K4ERZ5kz
gJiAZJaF2jpqmq/K9J0G3yLiibM0ovBqov+cJU5csRr47QLTjE4qMEqBgVc5RLeT
nqqfzu+yZe8ltRLmlupWrU/iY49Ht4MRXHnge7Vj7+UX1DcVXdiSzabO0nBeLa6D
7NX3bUTDfdoj2AwTm1C4dlV3IE1MSniPhFRP05JmF2lWH239gAsG4m4FKmGSDiOo
UMErauhFhQpk50ioTw+8bHAfnzjtKvrnZQ5jx6yFaCED/alRiE5OuB4/T3w8ljqQ
uNF679eS6c+Xsv6psaAFr2FA0cIlmEkf2Ge2rEDXJOqgVZXVju8gntf8QnNl13Tt
9flaT6+F4OfbWYoZIwwodLMiPbZuXc+7MZuJMompUC1QgwG8PR9LUQghTegYw+IU
Qmp8oxqiIEiLPr+uE4qpAIJC0cO4Fn9MMNc0tXw1EsgvMuTQdp4iky9HiNZddA4E
D+tQaEb51p9WUJjXkYoVW3rFV7x/Idydt23V8SRJfJSLoO4lqvXysy7TEkfyAoP9
h3VjIo0bOe8KllApTYGLeGkPJCfuvPWvUonVfBnzs+x7qt/xrIxgtNnZxPtzyoz0
/mqm4FSIQ023rqvGBEGMaS1urkKzoleqhTcrv8Ev9OQ4CtArNRwTfp7w+gubLrXC
78ulVqXhihWb+Vvqe7Ro1Clk61fy5dBO6h5rPApWB37rucLvbE58Jf6WIzEIIGv4
riFNl/MlP2EBGEWmT0pFqXUuVhv8A0oY9KSkLsdpvXbe0dVfUH5GdDDM6IEHaARr
0bMl3vbxzF2qpzTGQTj68PZVsT5sgoFRFTefQJ4zFAV9o/28TIoWUWZhacJHnaw7
p/NLBjf0ChkerIiSwIAurU7Ufp7lGpXr535L50tAKG6y+j9dr6IuKeDNig+mcsTx
z2I6bR8ZhJ5xFdNwEtkjwFV0jpd8FgXd+SvyLn0fAPUDCbN7m8Sg5bGLEjrepzX6
RcpbQN7RwGBVnkZdJNZ1RF9PQw5himW1+zmO/t8KskV4Tf394lO9xnZsUJSqfyp8
8kro4pGrQBLucsTTmnnkaONaY1zcjScp+OEY88oImUtUwxMJPtIIIY4QyPPwIFxR
/0ce+e+jZ3f4T29CPCfmlhAPV72/rv65V7AZC2959YdY+RFrmtESMHH/vdaAHS5Z
5UrzpYTJbomeMxEFOs7wzF1TbEA/au3No6xt2dwRuRNJ3ImCdsLvhkhw28Fbma8A
blL28H0456EaEgM/QHLnubLQTcI9szZIH+guBDrRZC56hErqWmFiZMqHVBeO6etw
3H95bfuzvkgdEKG+UpzO55F0NJhuLWfj5TeDrj+fmo+KHLeEwAAsARL3BH5tgac3
XbeTC2heqxLKrQogNXxDNLsEL6tkKpghF4GblX4celYigp5F4cu0uKmFbRAGXAD4
ioJxxRkl+svbiDZj0A4BESQY92fwmdWdh902B5qoGGSJHjgR2JhzIr9JYV47m7DS
RHJV1Wq2UskAVdUlUvMj4sQo+wA8HHlv4wMsMCV/xPWDEz/FacCrfT6NAgLYXeVW
ZsmZM9v4hr8aE/EjArzFB6xd6bdBY8/rYMj7meCYpdPsXdVM7S4i7bMFU44CeB1I
T2xm+pPp1CW9ZqbHM63tP6grjf6ZWR+6hOjUnZmLwZYFABC7evoN6ra5Vl6DdM3P
5OqBMQKFfe2Cmh+8NgWxUZ55ftsZxdT4afatvEfW/NO4p3wUbrotYesvtS8J7lkU
kNXGaLz2qQKqJ0jWnoP+Z5g03/kzjqbDt5ebEA2ahNtaJL3IT35061SNai+Nf9Cm
bqHmeT3PyrnStXjGOzltq6mBoHVWKuw31mrvkpPjnN1gMgDRJwvq3YqlLvPna0PQ
qXRgbmHJkVgDUfthoO9jLMGF20rgxxDKFHvkoHYqyGEd8bj7ww6jQRGcslwNXzVF
k02u7HnbR8PNxtJf6yDiT7DBGGmfzjDlQlXleedOWtHght32W10s/Vk5C+dSS2Io
EvLDkBf5hIRrvg2CMbBBhvZc6USbbpsE3pJ9UYc3UgIVV+vEtzwzO4SbtGGEn5Ec
Xr7DElVZ8QiXluKcJ3YGC2Mju977sEdd0zqwNEdSizzKsXy+hAkRy3OVTLpWAYFZ
cZb7V1ybFbGp2KShQ2wJ+uZycZ+p3YAD8qyK9irU+4TQxvOfwALo8+mtFjlReBjp
9XKt9EwW5kgt55IF2u4yqQIpytORplk3AcxvZ6gndvrBw6pcQyoCqaukiEHGRAXW
KSDZLNfKlTG+HLBsE9MlJVdwCE35owb7WVSKLRoydtrNpS8+uHNjtE3QUO8/yDEw
RDRIFSE8MaEm5+olewYoNcyozN32uA2RYLLhGsQcZzzatUNfz9HUHjOFCSlh8HGd
9xJtzQ5wWO2upCTS4R58GG438ueVxlfldXvJDS976VX0o7uZBVzA6QIG0SaFoU5h
wAvT/bMY5qc7opHmv399EPxTb/juIBp4Yw8Kg7xIFa5/x2EQjmCrWFMmhW1sQCyQ
BEgx/ct5PCg7Jk3QV2JipsNLtb73qpM8Gfa3Ui17n9US48FyAXz0oiG2n6NzvDsK
Li8Hp1hrNZUsKV57adau49Cy9ElcIPpUxBhr+oYwshvu9GznqcFGpexaXZGbH79m
tdIiTv913NnVBGQ/RUfNYCI16ruAdHVXsVPhAlacJGxvk5C5JcFQKpvEUdID+rJa
TlFUwL+Vjbr7xtZ2wD/pCycedHty1r8plXjoYaXJkT6cMqWSM/QfMaIQfSLDQqCu
oKIN7ZjnByg9WNpP6GDpVkrsbBuK3s6Ky/qwPZyxGiyklHqiYvi0WRfO/k0zKbDK
0ubLW/NgPSl6I222JpWMrIoILXZeSAtoj3CbZ1ddp1Ad05UZP6R+XWpq1LKenz4m
/x7yi/58+Y284/KH6Bc4CWGgTq8GR9eg7dlujGxaO2QfkP/IgsJjQ7aNk7HIkjU2
Gp/jypDP4zU5kSFGUPCnvQavEL5Tc9FkFieqX+EZb59dcggsh/SY7BJx1NUhz4SK
964kw5O5jrA5SyDa1svIRa7sNGbn4fqpbYsuT9/VaoaUzF2mlnmD5ffkJsCg5x20
SYOVR/s+gsM36WmCvtzOXK+HHY3TIa1YPBc0+GyWY3tNt0TQZgew4SSjbnjifXTT
xGy02HwOL7e0jhp5Y/1zmcddzGpPXSo8lm8mvh15NB/LehSF3ibxMGdK/p+J8M8x
gTD9NGv675CNmVoK1t72dt0ZfRzxC2AYP0HjR4KHbncV/AD4YXPqEyEWMnoNC9E+
PNl4zc53ZL3aVM7HOE3VkH5UyTlpt80asj01+xdg3C6sFDILSs5iRRcHI4s2P4dk
6E5r4VRAbZm+c2cDgY41YKcOXei6MM6GZ+1d8BeAOQ5lcgZYhVzYvsVDdQcAUxrV
g3QpW2ZdI1dlrjDxA1jSDSWbWBFqgqXekpVq2UpZ7WZZC+EnfB64g4aCy65x2S0p
U08GOJzmpXwpPoNkTJ613sm+TttszDty/2W9iNOBJAjgSOxBX6jXJYfzVhodZrKi
29cKb5NHCzfdKhgvFB/j/XUwQRRXMGoWWw4G++xfJL3INw/n0GH/LRr6QDfR5BT7
YOmNuQVRaHSemZgtUOzooMdKvuTOX6VyYjDL62ju/9pN7+WO2H+jzHE29QiC3529
LnpT6viny9asf6w6gP1uxhVaStEDH92nJVOLTZ/Mk/gNEDjLQpGHammW9CAcCKAD
nW7n/tWe2OC1NqIhEvHgzWh/SKKxlOaISJZ59lELT5G4/n9rJ5Kkrs/kljvYYYbm
dTlCvx/vonNin2M7GDB0B0dY3+5siwdpPPzBID4jYlCMkjDwTiK9H5mVxJm2YbVX
J/Cn6RzuyERBa6hmyuOYtIzfRkQnkzWvTSzgH985UqnfUusF/QdonKo5gZIFy7xc
5L8Swg/cLx5dhAJGQcnPfd9W9bNHE6FAj/4Wh+tcJ/dP1cwLFdmYuFcfcdYYLwZa
U0dCwfw+0vMnLNu+SKha10ThJbHyT/sKOefHwwRTrpTzRHYtw/tcnCpE52qY+/fz
TI4VLohPl+vwd4X2iM49NPACnhDVeaD904J597rRuYeethStl2DKhN0EP3JJ0U6/
FLjKj8+7vqQnxbrUG/SYJwqAYe2/pnEXTCGtYq+/gHQk8Y4RtPSROO7XvWGKb/FY
Nk81cjXzwVHno3/sw8Q0sKsxKBakMacy/aNyHc00qi9DDLodyHKSoyanIgDdat25
qU84wFbhyIXMB2W03alJUja05s445rngYtuKkvHYsJ/Xz6dQFGUVEZ4C+20MuIey
twOhViwWvgZaAN5HixspOirD0Zv5slaPrKD2Kh2U8TuVIzGbsuZzeEJRe9FOr9ii
x2wyX8RWsZIjJFcQpuyunNz8Ias0QshdA9okg98d/58sb0WaNGMex4Jwp8N0CRz+
9xhbfYarYW7PvmSDlqWoeSTDo4fUrYPSahQz+2wIFR/uVTIvmOFhTp7HX67JSRBE
+ca0hx34eSv+M2WlJ3LdaN6byvKIaniCGERfumcHOrOChA0JgMXf4tmI4SSJAroc
lvUJvnY/Yl9vy/jQA9OBRP1Q7UM3WIPNxwU/zUzchewsx9UB5+oRY9sL/DaB5lDc
TJvbLxcxl0RqtA0u/gcPkDF50kPWWXayTDVYUKe5GS/fqCc6xdX7nSozCskqYpaV
bG2pU7nDHUQksxpEtgAFnthS0t3DqixIhMsEVck9saj+3g6MQ5s8HdvtfUQn6z8M
oiDY2iZuSqHTLEzRns5yzD/HTZmmnb/RIQ76L+ep4JFdbEVVbAzUNi+MXgjMZ8Hh
UWoiRIzF/E6KuFADdnRtgA3MWqE9IrKNrkIrfu/TGsyb33GSWzSy05NrjY7B/gX5
FWmL5sAsUnRd5CrC1eBPcqfcBLTV41v9aItNATFr1RZ5ycZKX0izjtT8jlgBxezW
wC7oRSDw0Z3ir++4KpVwebIfre5a54XLBYw6UX7KQpbaKEjGXAUSkzD6oOwD3jrb
myaoTnyID+oPjr0VxwrV0rM7QIkkenFaNXRnr4OW7CzYyyFI06QodTJeto7Kv4zy
vsk14p/efC9r0XbhH2tErxLd2VIEcZpaMuLsYlySjcUqYqZYvM2+Ns7UqLK0Teej
Wh32XwE7tVfw79PDRNgdfeRSLWSU6JFcskSjeLYUDDAaTq1BEA7lcE8uEEzrBYVr
1ClhZwUGDEgsdImqguzFNY6Y9SU9D7ZmZXcZ7MTrUPWJzP+zIBMwGPI1VA30cJSq
j61xt2irnfnXhiu5uFixo+fXH0dqf/qyGVuSefO89E54utW6tCheFJjXhAyleNc8
OfzDkGOZwEqFLAksZOJs4xtXllFLwE9s79JZAZuPQJD4Y5jwQjAirozrFqUAKvtv
qBEe+SLOwrHZ+xrZ0vgimsLdjJQ6uGQ0l3AqJy3pJOmJGClnThseLbUi+sWhTsUU
vXN3GvQMV+kj35rfqI9nInx4ga8ZYULtk65xjNCo/nMQrAEYdILug1VpdfU7QWZN
b8t+Y9wh7lysoa6nct1MlyQsuQG5145Mfb+AQmtm2/QKTkRAujUkbKjfaqYdLCjL
izMLRaVe1ltJP8QddXE2fc6PC9u9HUIMQVUAgSWpHAbUWhb0c9+3twV3nu/10gKu
hLRK/IsuIbptNPFcwtLkc5sDwfrWCMLLw8ZU3UFUy9q4rGdBVs4S6xrTXCylNjWF
mJOCxtf6peT9qZHiF/SmDGOd/I4pnRaNXHt0AS3IxsYSOeB/f5/rH3TMQ7jwj69V
IxgpB15HnDgqNRvGrjvY0VZ+p+CY5aMyUPbmfyouAwG1tYvuRYNkFotLKs24iPTV
go89cinSvlqfij7xis7AXcXhPwHObIZFuHzOyChBBfyrMsvMff+QYmcY4Jk/ApJV
cOL1Xds+e5xSfK+Tdc48BhyRL0rtKHyRZ+iEFbJWhRHe5wmzv/NQG49XWfwZj9n/
7r5DXORWxLg8br9gT9EbZV1Vucf1i4ICX0G0Pje3ziYyBF9cBNMcq6aVtljfF7z5
209XgheqxQyM0J9y8AK1xV/vtlSlhkomCUSfJtAbDOnCjBKXGRrbkSaJFnqWsj1a
Jz+5dc5Xxwl+XUkvdVy95q8EVwd3ZWCM1EsXFxSRWD3d2zK7rLcZknmgssi8ggcp
kEBqiJc5rQBZ4AhhLqA4+V0jarn1QaZ7GPYZoLZhryZzulTjqjR/HaD1fOV1IcW8
q96El4pPN90Rkq2sdp9yhv+y64XVhln91YDGBo43yVmUHCTcoV78IQp74nc9cvOE
lYyXCayJoU73KroY4D+8kAjIesNyYODZo2Qs9gJghWwOFUeL0hb6/mlBa891n+BG
7NIAXLTmHz+YC3GvxIh/dX1aCm1FSr/XIWDHKPEp62MsY5DvjdlARHk0O9LqKiiw
rO38bOVyPobp8g5d36UwKpWIA52hz54MkqyTRLdXHi34tkJYsdTrUgudVu+TzWQc
x1rBRO1FEIccfv27Z2TislHUqk40F/0jIMe25r0zyjfFL2UkEYilFH6z8YNHmYw4
mLy3CY7VoHmEgWLiD/jluQ+TR8JfIj2tg8S0g6MrYf8g6ynKgfTUuqIs4GR/rDi1
dSYzD+gWWRI00PUNtIfOnBHWfu7f2GQ6M83tch154tM1tWDuiPM8mc+ahyIiiKAm
zCKniPvKiB8uEVMPsvDejLMQkL5AZbV4Kibe/WZ9Ko1zuESWDd4yZIfCSKgJwpC3
PoPvev4Bf15vVO9xVcQrmpN+gMWgFx+xJCq2pNE7R/P3YqivV+x/E+U/ZfYoQ8Pv
IZTdiR1nObbwT0AoLf4KBxiH0XjNOW8hVrJTJdLFYHBclt+6298d28q+uFfCS7VP
1iYba5PhHqZfy54W/rG8N1YBvwSOTekVrhMjg/qrjhO+nXM3XXQJprA2pPXiasPa
Hd3Wp6amIDM8gQhKwZmgQ13SUFZINIMSyZBnbKg8jV8k2qKYd4+Msq8hYp3ET0Ux
aRU9j3I1AVC6jFmOJ0I7PGZoDjctc0IRouE0DnwbRr+So9lz0uUUUMMi0UmjjNHJ
rCZRYIfMqvqDOIeHZlDlDDVFQGtKedfqHFJJpB+GouHS2AKjm+QCNUDkulf1erTw
VjUOaiv3KFRGUqPQ72MO9IfmoCYk5fqcZwBNQbAzJZVzR1hjraEV6VPHzdxifZNd
Zi+R11ADrLPnX0ooxIUM3lFI0i+5Mxqyt/jHLOYR1X+cGapZf2tS0cvhKr96viys
EwSCGrBwjYFz2dPAvYggGPXa/ztMEHwYPaNeQXWFLofoOMi7QHzXFiBSB+2yXbsw
FkBCJYKFMPk7cRyKe+2wHLW3O3GkLAhkwvazrlbuLtzB2EmlH34QOIn0lc/Z+xkt
ECzxzSV3JRvGRZ5lVQ7+pB1m980fykJ9MBHQyWM+l1NE79tgNmllIgKmPRs5xgjE
oQqtWfjNOk4I7LB4KYRJCzb4U1OgY7E2tvFtQyrBM7xuCAWHTBhGZ8Wq3hhzAlnh
409LkRCuD0K2bKzB3G0PPNtspWmf7FcMnja+l1a5Nka2tsFx5cKhPF6LN6ODcWW5
r2eiesi+XVkEFYX9NaiLPcnQ0Sfj5UYNcopy7dOxL93wxTZSxiCxMs7NTxRAgHDi
F+AIJKMBlG/BvoNCDOTtfe/I/+Qa7LUoz/OaM8oUJZMu5fDU02FT7v+L884gGCoS
GA1n3zP+x3REMAG5S2/CmU+P10vX1MJvIbPPxb56SlKd4y5c7weU6qSLfqNgjDaj
XV/Uco84iQjV33HEDzWOaxSpK2adGtOUjY1uquCuRQanhx7HpEZVl3z4AfY06rPQ
XGmQvWa/BDAxGihp5d5vFO3Xj24hM2IWLEY7dXeOCG9t7sxbMhwhLorPrWc2ZCrE
VlXkqDDT1eckL3Vni23+Y29RYVUa/cnZW5X09gpTDXN+mErPj3RmFsBiGpptWn5A
hVePVClBOsG2PnAzs47p7pv+d9+WE3HtatOkdWqusAiJEvGer2bN6xAOWxakrtJ7
BAakQuAUaArMShJDuxB1Pmm4oGuJYnd+BHHziqtM7FLvMCS9t9khp3/KLuyYI/ZO
A44Qk3S01A3Dx4qDiYowt4nEAQP/9v40v7czhoIzTScu7WPTvqbBkHl0kEgpt5e9
s5dn9gkfh5oEQWwCRJqCjMTBWKCMVqDFG74o7Yfthumgqt9Tn51huK8lMj4IEruM
ISmRMSs+Hea+/jPxC/AISXNvzK6RVD8C4JTDV0iBKFHV7tRnPMbcPhB7XeWtCcuF
eWPXDQImes+2NmkxvyKqEdvbzP4Gz/HZSrogRw4t11V56j+/N31kCmEkiCg7Glbv
vSgPggJo/m1CqvISyEvXvrF17h7uq6Q7aCKQTVqxPmOgAs0lc80l5C8+VH/IA/WA
KfTCgKESVedL4TkQr6jhVutpkPfkZY25xZriZm2k4LFb4c7Xlm6f8So2Sw8FqD+S
Dc9NXEjXRY+V3+u9um0vsh2L/LFBO26y/Az+DGZOyYcer+G4t1G2lC0SIOnAPrSY
YgPqOVpXjOQwrVyXOHgLJMpZsDyZoNSsMktlzQK7vPZRhuT5WgbXyh+6wUCnYZgy
8aWQ2ecL1SCRSHl9yCgZ2LVXyBk2ymgBbuubEFPB+oO4RT6EzgcBN41kK2e/bpXm
u2hCC6815PmA1Muazd9iikxQC2OLnsz08T0brh1APJmbQhrqGZzYXZUYr9ZY+2O/
M7MUjSBZUOLN8oO7GwwQcZfxTpiSeIFhgH73RiPhflRY7o7mWkNTLJncJ8rh4z9z
WH/cCjCFAvGQJDSLOD9Wal4DykJ+qS2G8VWDbquaSw9tTMtIM9EsFFDvseMTSo0w
REDOFCALMatLfUjUNzpc+CCWUPIxtNBfQsLszqS+1zSApUQdqmJCaCtLxRdAD6Vv
cLZ0Qbi/yBzy6ORBcdTd28aCwYIRhy0l/+advFP2JiQpmU0maOdMz5tAmS27udP2
NEBGey+QJVOxYw6jhOq4ZHDEFxJI5gwj07TaP/4KZrCz9JGMAs8dgmcNE0kz/UJw
Vhj7+Y4mGJwsveyYdsy9a159B/h2rJsill+aS7cB5Yt/WB4i4ixNgWjTmmWICKE4
IBFrfU/+emdZTS89DgT65tQGl+h494XUZVYooGnP6fMaaV0DcoZcGz0R0T8Mucur
jCe3gkot5YkgtFjW4nnmrE/8qc7rl7bWvOTO9MsEL1yTHN5twzF32R93dwCneaib
gQ8WzbJ46pDdH/9r0Ut6QLDt7p6ejUrxtNLhPuXBt6bsA3EsVkECbNu8bm7mMejr
KjedUJZZx3mS7qGiemlmV4kv1JdO+eqBlZcHrQHijALJXHyJpBrGkMrGPnkfEVM+
zanrc24WctrUhKJg/4G+4Na3gTFsxU8fq4L+PGWtJe+uXEu+CvU+17k9lf760T6x
cpMOFNBH6dRG9A9oqROEtjdfBQh6epKUYJJtuQ3YOxesXnSC6GDGaD2xsctkC+wC
NnYedr01qN0Fo8N4WeyKa1qT1+2a+vQNvFsIMFcsP26OSVf+QUoeGjyaXWFRZF9O
iEP6S7NKIDyRcVpHe6KVOhrGwlx1SSQxU9W643BEL45+seKJoeXbeH4NP9cNBpGs
s6ZRRylUrGPBinwM5UxYnUn05/q9qd+aFm88wyevPTRHhrTos5oEVCIFLMAV+jnn
I6UFM5uto2G/8EVdzFrnYzwG8kVMV/gD/PnRnVFXpeeA0h2T+XyduTTgautFkzhJ
yMAMFmQ161VwKXEk03+QAzgI+zrH4UCHd9L6ebFZ58PGl1fzNEEha0OHTV/bvRTp
JSIYH5bTFQG5o/mhbSz6f8dng3lKRY3kSUhT9EoqNVazHpsuPl2EV7V+GSVujKXT
CdSnS3uqmzRbHRs8LVNG4q/mzd9ntiyTVUGb+N2BZu+sxHz0RzUs+ZcaldmT017z
0MZDFCl0VD59KjqNbxSUPHVE6/410ZiN5P40ePlNJdDEM1+PdOVRPDUnxoCrl3NY
bHAcK7JW+lRNqAh5L13IsuAzl+xqIP2sVRbRekt1F0oFw8uBHjwfWYrjrcd5sMb0
mz2+8drNOYNzHolTGU2Zy3yvCVUAkYx3odRjj8EyV64XMev3E0hCCAwfphwGJayj
knU6aEUteRodOFOVkHdHUPp/nL0nSESaKLaMukMnLbrnmPNPdLTbVZ1amH8LLTi2
MweVuYcfRkltGitZdOnLIVXIGue2HTRaYVIlpeg0seKhwo1/eD3g1Oa3BpexQRVU
hTIyBeMTK12qR0FmhaneLKak4N9Yyw7Yu9Ak+qpsNtYN1CkeKfmhecODcZtv5GBW
m1dJWNPgz0CDYlt7e5LdICiHTmP8mKwPcIbGwqhTlxdfPVZjCbXUqCnDoMkH3Ael
JER9kCWXn3cq346KH1h73kwdhiGSfn0rdngGVJUwgcRmyZvdLSc8D1GwWdzJ/ok+
fWKRNG9m74aIODXi9jTDc5Y2aPlZe5Ii3jfq+mcl4NCVt1FTp+GFX4IpeqFF8vin
m4LBftmUihHHxmfH6Zy49+vG9isLV4mst6ripVCDZLhm2KsjRjcU878WY9yw4QzF
2mJdz9jJ9scRa83feKYlcl72rVnqXlIuW23hAif5WtUAWFQDe+hsffLSHdrqxJD0
X5AEpXAkyX9XAQsW9NBiZgGvXfizKOb8HjaiGCedK4D+fj777C50ZvbCzhLOCagR
vMx7RCW1jQhQzGQgXxGsOfenz19pWcwdT6DdnATxliBRxiUhnZXKBR+C0e09YlwC
Nn6LigIN0mJWZnUkyx+U8EVOPKVWyVSRhvSnS6GYRLzOi3GN+VgnczHoHhXDjyqL
vKvv8uxUu312RBz4slSqLB1vxW5GBXslzJLzCsw01MoRKp3JiW13FJCfwSgPoW8E
1UdAsPRfClOqMj/xnrDlOHheadMyj263iY3IoeBAO5wo12gVXh5jthmTgEfmnl0I
5CQGVLS13hw74hTLo1xWAI9aAhq0yKCeVKAYLT8Gwfu29q6fs/DAyRY8iswkKbWo
qqAlrBF3oA3sSRk0cwZWgtpu84nbW//y8QXBGPtliaIgAMBZVT4VCxHFEw9HUiMi
SwsuOS1lxwnYPFWPryBf7Zi6Xd1ScD92g4UMj0rsL4OWVfS7rGwfDe1xz5hqiZIG
SS0TP+wPIB5tbvyA42Pzunr7rf9oM9rD2CnwIMObyiwOPBV1wRY11klvtG4T5PNc
bMv/onImR82XEjpBKPsuzpCN+0sksA4uho07v+d6+f4CBXwetQjNj5lDkT273bE8
a5krrb8fDp+FlSaiHIf+d3LLOiyrNbuW/Mlk8zqR4r62LPuHoyMYSLwDS6QRPn+/
K/wKiT0u3CFC3cnE+qMAc/XLFC/txFlLSXKDssITi1mQ7feY2+++7XgMQzzlQ+ZF
8Mv+vZk2/IlIJcno40OCkPiz7uNUq8OAldzlrzsSH9i3x/c94h56BRmFRxwwttrx
y11tar96XpXHlmTRCoyorTR4l0K8W956O//pe+MV0OSHeXzIXHEgBCdknJ+5r5wG
KpOW1MOa3QEeYH9NXql4J/mJsSHEFASTfOMDG4Ul6wVGo35Gp9/KdUH9yJ2WN9vc
FaGtW7mFAPzkrcgnr62QnHHgJ8fjtFqA07S6iCWaYYH3UenBrA6YnHjgYZlYMQO/
2oz5WAKwvFlBXIWi4wnjULYHqOY55X8khOghPNIxH3+xjtiwi4xbyIVuDfNDe67u
gT6dfLZZuaEx4/Pa1EtXi9O5l23O7iOaEtogN8yLN+i3ZVgtQhljNxF2DDcTf/fh
E+Qu3e7zgr7ko4Z3zHmHgapyPlfdV0lJf7mrkiCfexwbaYuBDXew8zI1wn4o2JEc
1GHyirC4JU7v35M+4zWvcpk8K0fjp3huiC2mME9lVwLPRwTGXJ3Gb4XXQA6p8Hrh
2T0gTLhZsZIHVzCJPCYt5nnf+3MMlvVnbtAR442TShccUMyaVlwzpntfagB5Wt60
gdnlorEih8ZwGjC6IOv+GYtliQzLkWPToIbjBHPN/zOSFQDol88ApOt6SP4leAsq
kFfky5JmaRPgZ+DWeBImZ8Zi3sBtM24e09c/8eOfkSwQdzeS9i0qM5vhqM+JpqeR
B6XhhpMyaStBCaQzvFtVvCY/1qyTu4K1g/vdRgKM5ysQy0NIiThyyGiATfUqKd8s
SRpgdZVLlzjQfVSSApLd5+znMYQCUhXcZKRHWXbCvTjTws0CoP5V1ldISKtKWzso
/5zfNlSyBu4Yre0ZRwIsmPWSEo/ZuSFgj/Tw8ndyKaP+4r/fXhyRtO9IczwJJrn3
VsEP8+PcKSGxD++x6ZTUvCN0GcAP3dLgdRcpydxQTfm9OkxNhQh0l+rCE46JMUyU
FOSAGSOUHlSdBoZ0+tXLYgUVfuun3Wy2S0894EB94l3iqlBgU0b1m1gmkg/Jagr8
k+GBNabacLJgs7AGRuss/QQsKWLvo5CiTUBz0A0FjIsSoPA+K1MmFxqsVr5OO0Lk
O6hd97EJbAVboHQXJ2sIisOGRFSCwQcVajLDFWWc1v2XC1CWVGoXDFLHBEmXxs6W
eP+t8keBUt3znuMO4Erv4qWyp3OhSE89BH13dtG/sdaboQBc2ACN4zDA+7HPTXRa
uKGlMbOXQFwdVxDlSvIB3UapTsfmnxIPo6mOwyUxwvJ+83aZ5/mpbjD5F30pL0cz
ITJ3CyO02RI5bc2es9eFk6XPCBRg6Cyn6U2IAQZdnN7xO4OpFL2P+QSiqj22+Njf
mWO2U7YTgEs5JkZhr57WawIDEhoNzTFgdkiEkQj/ziC2bk5jj/raA8FyYdoB1neE
KEBNI1WhthIp41S3sZBoix+7k5zQ3O1gy7Bc78q3b8YswJLlloguH602BrYU+Pps
6BSdHgKY2VPJY/vFLWNVB26okhAv5ekeiKZbe0yElQwSGpx2XSqD+ZO+mYWogcf1
Y076s6tdm+Be2ihEuFCW/QMS6z+lim27nc3Pb5TaHUdygKKqgrn/iYDiCHNZhSfA
rT4ljSYoP9Zk0KPKgTdEuLY6dgJK7vqe2yFu+RSlUi0HYwtkfWJpAMPHjaVBO04w
i3Y/g+J4QeraqRFkrIpEBqxM2AJdEH7A1j0UHe/u32kc3xCc8+2uiTOlBFHd3Fzu
QsSwNVRAT3z+u/0hc4Y6o2o/4wGLgITDb7BqFSRSDtOYb00s80QBFUXASwXC4gCW
Bx5N7LhDPzGkJlUb1OSpiKUV3ijmLJxKxhrHpkrn9+JH6YSRtGFvC7HuXYAjnBwH
CDYVCqlkP93hlT7fsgZCPa7ivqAPOvl5FC6J3t57ipy/oQg2x1EAFfGwuN1Q7oxF
3xds1E91cqWljW1kdgW+KvbzKkI3sKQwponqjd/l7ZvoRX+kS0Q36pjoE0TPwqeJ
cQTWY22vIxaMwjs6uAyU4eVq0y+a1pzznGm47tvTnF+RzoLpQDDde4nHZ6RRONpe
nRiOsdgzn39Krgy+031sHfRKhQLVWCA92IHlQXPGK6x1lqsrlRH6PfafBqknZWW1
GRrPZlRlRz4e1T0PK8bnkhVpq1pjSvifN7K9O6RWPFue7IRPh9jM3SKWRJXpuq4g
Pkjclgs1fwiI9Lu0GxbYqilMGS8BsjYhpMlJ8i3Q4/uXsCwKyXRhTXt8Gs9w9nRH
SFyOCsrB6x6AAXbyYFOrLHvCo/nK6K9wPQPfEREGLfC45eXfmrdqGrlYF6iqP9aO
m9VNfwXaXz+JE7hRKFwVnG73DvKa63LQGxMkNl5oqhaWbCvOkO4jf83phZ7c68Gk
qQtZoP4eX5QKriYhLHxILfDH7prSV0sZaTgwmgtqP5JVrffY4BdtjlOqke9uy+Ba
fIy7Hx2hK6BIbpeX1ZkMyBqbaUBJHPqXhBP39qhM9GfAIEh9DQ3J8vncPNRlM45+
OOqAD6vQDmv/KUD2y81DDMtxV0SRRFnPT8HYQ0xnBKEyaId0ZUsexy6nyGKPuUa+
TZ7w2IycVfanJfruZZE2rp6xlCrrmCh1itP+RZa8tPNolUxha18Pclb55U+sRVuO
ZYTaxTXcuwWFVSLKYRFNDhLxDCQ8CnNzungaMEtjHNTL8Fm62V727Ik9r3Giq3m6
rSOD8TuEpp464lM+j7O6O92gAzu8jK1g3t5Rqzj+NkVM1l6HGRHaUrCAxbPulFAx
sHR15ARSO2AUPyjUhnz1FTPXCjbfeuqSg3vhUDHPJG6X12UzknwwPEQxmBES4JgN
tGbfcxTtmKbFNlIxJ1VJq3sO8oUTnAI35VijDD9U31RDcA4eEaQZyBocolwBysmt
XtnMX8TjlkIMqX1HjxyBRg3wuPHOS+fk2XMm/UxUqF+p2Edyb6cFiQWAqu/R0b5u
qPIkh1wreRT3ugTkZZMpLmVde459xb/glLcW+J0AGB5ZPPK3a331K8tIzSYOvbaM
HEx6fGcPtXPseyMtdvBKUsP7C6CM640vG9NwjNKb2OpwfQdD5wHNHcUksd9j7n6h
eV758+CFKWqdaceV4QrnKlqopQ1TcFecfYHdyO7t+NyARtlOnTfioNCo+o3HeLQg
7kVRNoS8q25yFDAYt7oYDV34LnjBDtBma4TapE4F8Tq6RvsJ9Zo+klzmtV2eimpd
KQvOOgFdBfvWuLlp74Xu5j1RcwU7FDxL3UMvPdhuE/3t0qkCQFjKsAcVeHz8P/yZ
urH3YAD20MutIcQNO/kS3iQ1X7Y+nQ9YtcqlT72lrQoo1HiduwH9MiMfNyAcY3Vz
yUoOCFqFAlg3YfTEOHuy7zs7XrtQSeZZ9DrcKx7Y0D7LN/7ePuxEIaUECi4xMn4i
06zPYK5d03+Xte8EEypFY1G5h/OB4eIeRZtQ/IvktAm6oenMULPPoRrvOPOjJL6B
w7rNHGSrEgOw1ff6KF08o0nyPMNyOFtPihmj/fSmDGtuKrReuemdNOmXzCa+NQUd
xSnfgr3fDeHTr3LmiIcL/Qrg4Nzx2YyY2EEe0WHPy5XKBqAB5QP5C/vPUi8lw0aB
eOAOA4hIU6hIXc/wVNhP+PdAXd17znj6KD6KcykXTHTSqM359fuX3ufcM0suTb7o
thDwqj7y1yS18bQwfnMfQ/DJWnq7N/WNA7DBjpTnwds4BofnsdMzfM3/qNaxcocW
q8iDnwKiDr46uIpDFONnPAYPYNfRuwrAKsL1osCTX9Kppc3n+lYWczT4iiM0PDs6
OX313Qlayk5MjugtjsyBwG8APvQ8qrjIUIqhghnzZoq1GoQOfyvbnnWOC/ylFv0B
7HhiI/Q/3PsSNqcZEkjAd3xgDTM9M304PIoe1tALo3LI7y4RX7XRM5aeXyFGb97E
2asDlibRciS4Z9ULOlZwDTH+WPImZBeZ6Iny+J38d1i9D+vrKWPXu+baPVqGw50y
p3LpgvxuifA9zV7aklrHaGvo2jzp7NMQpn1pWsrSmbEvi5Lh186o0hLZnzeyXFle
I/3XoRbjSyOY0/podaGevOl3ZiXlBAmn/Rec8VQh9FThdT/tpD6Y2vJf6kK+iO2A
WFxDOuGrZarFO/LnZ8mart5+CJH/qyfk/2RsTuQSB81bQbzFkwi42mksEvLNd5jM
fXRws6xxSYdQgGmvHBYZ1C/sc01ncZhkr76JQ9O8xwqWrZc8vcz/DyugZ7B5Mdaz
Ze5vwx6WkfIjb3Htb42WQxAGbO4Z6jJr2yVpJ+rnXY+mWNmc0isQPmEvpDBUD5Vc
3a/9i4B8vnM1PZIeoP9b6hkssO55n6ycxepPGBVADOrVP6HunAEU4y71bp4oHAB+
PW4rUJlvILTgRAyLuvwhBcyMwFTTRYeDxg44qK79uKm31b2hoae5QNlzLd2x8G/N
f6aDT2R4AyPhiyWaHE75QocBNgzin1G7DtvYHC1VdufpF3gio8TYeXqaTt9CgRIi
PCi9FSUr40KARZwXRHiVHoYuf0gwMpxqvgzRJzbLK5lHTvzi14FkH+RXDiHzT9tB
E6cjb5Wx0x0hG9Wp/x+XrGxStFDk+Hrn/F4Xn4IsyNDC5IjDtAQHP9rJzgKXpKfn
ad+/m7X7v75MS8RrrZIzb6GDqdLgGnnPhEZLjpGmwGO1socfnM3vFUJiI70pDBX+
z/pn259j+dJ7agVlxT51WCZvbX7M+SX0JlttzcTRzkIb1eTtBCyzCpc0t5FrnJ9H
SkBFD1DE6iRNseEX7094/xUYO3t0L+qkjB88Hb21o8IFQHYuAEVqSFYrxmOGJ5ms
y+oNN/WBVkpXavIoiRYTMrYN2Y72SeDhSItRPl3cBsmIYbkUPvMRfkiD3O91/7Nc
i+22KJxN12T8Ypjf9IvdO0+EXryAusMlM8g6awvfKS+K91I3LQmDgwPlzkEhqRrB
H28uhQvjVd2hGt2NhFfCFa0Vvl6YQNutKK2hjIL9bILqFNPn+OJbjk6NpMN8ryRF
utiLZkBZHODLwyYwKvG/1yBeumvSqeGZ9dg2l5k2g33HEd2JQ3tUqtkwg5AS/Shg
aFx0PQK7P1/sG6kPitjVyuJU/A6q5ZmYPsTTfGfsWNikU6fAUfKn0dSfhsZeRnTp
7W9Ixwbmp/hJS4JsBTTsTwkoK4AWGAjqiNHgpZjQCUhebR+Ux9gD2hMiNhCk+nl5
Yzh4FPficgHdGi9fw6pQvm9BL0iJJIsGcQAuDGJnvssb0SDvPKKruczbTNBNOYOj
X6fAI52hR1JN0z2qCvJB4YU6ZTDyprADsAOQbJB2ylv1zD4/60kyiY1/ZonET98T
i9JXqMo+u6ZNo92By22T6r9MLJbnTIo+6yD6ieZWoYkbi7K+HqfudfZDuSn9hqVM
0Nw4nZD2Gvn1kYJlKvMN35BZT3PcuAgMlG1eaKuc2eNTddb9vu/WSert3nv7xehR
SwrTjnCNuBEmtOvuLHlpNUwqTjrlUMHv8JLPqfamomaZafD54jVu0G6sAXiOkj57
TEHZDkqXqZ2DCAYF6TnZMfz+VodlbYTvuyV3yhFSTGJsd/DICSVdHCijAvJ70ewl
uYnDtEtZXXcSWLnA89T0eucgn3PypuO+kXDFEiPMfdy9aYN/C81aYrWyMrh2WQtz
CKme7zJNaYIN28AO+QGhBJ0kFT7Y+DyomYpLgWEgkyAiKieq3xB6ADEAx76JiBGJ
qaIdUgeAiVKh/37x1pogAHkCpNDhOuUnllZI6LZdDKBYId2xl4MTftYecnv5yVSB
YY8eantDaL/pe/ZPDSM/SI3RqFyVTXbdRPdKqS6OG9hOpsxcaSoAhFH4aP6Zo6CE
TKq4vFmH9bllnGc5H5DdI1WJ4s42szFQsBiRg+k/o1zF9Jykvi6eFgiVgH6Vxvpl
VbQSmcMNUFaTdbT1Z1s6jq+3eagXZ6ySCqE4UUB6GmNTtO46ZNCCZJxyKP+a33u+
+H/RDW8ija6YpfAq4ICtZAqjWPitjClnm/ztit9+XEvjD6EEiHTroCbV5hW4tM2H
+Wq4cTe+2WLeVf3CvnzaDcI+9IBQZxjzw9qzJlc9TZtvQiUa6UkgU43LJZ/9SApf
GcBmYl5ctWXej0kjZwzg3wWP5f4BxJ0ihMv7A08nINnE8wVKJABBesXHe8RmWjm1
ka+YFcN3UoLJNBq4nmXCDxCfcDOd32ge6L1lQClBoNxWAGbk6BPWjf/+5hpn7GXA
Hh/EmfiO+lD3QGcPhhtNINOa4WDHdPn52euaDwOsuK0A/nsG2bQcIOl1GMj1qZ+R
gTpw1Um+NKT392M+vVVJMY6OSGc2JiDyQvo7o4ByrH9gHBsS0YKHDchLPLEZbDWG
Rbr5A0UmiJHlwOB+spoF0GeQp/xWTX8maCm1wikZGE/KELCjJqThtv7kk78mX2Nh
3+nFY89YSdvdfXlWReCQbDkGE4JfNqFLILvuJl169KLzI0mPqwXR/YcyjvX7R7eW
4H4276eerXhIi/7HJYdNxsc75XSE4Vq8bD0uZTrmApDhTmnhjKDw3YMaS5UH5+pG
qy1f+YzWq8T7UrrFJdZXZdXgKM8/Q9RLTnrDZMpYXLGFy+b9aE+sZmVfysxmcmsW
lFQBqY1SnUVlAYfYjD+MrRsLeC3mkdWC1H91VM4kIQ9ptEtSFi/1tomnYp8K+5fy
60LA80AC9yJJxOlz3mqqAXBeXS+RfHfXuBbqMvG8e/FMK7Ez3pdHSUMHVdhup1FS
mDxcIQhU3hynf8O+FMxxfK7AF0U9pjuoreMM+J/13yeamvNswvEKZj3JeDTqBiKF
3MGIzONhBRj25e5u3EFqNyZq5cklJ/4VE/dNg14xTiD7Q/v0k9yCkD4JV0MD5tOp
+Hg7Z5/LeMxOHvdm0JuOvI5zWlS/Vr8x41XShCd6jQLtxHgTDEoUv14giOOk3fkL
Af6r3rlz3K0z9ByhP7zBev8ME15CQUD4NheYI9qpAv3Ajjg6tKJ1h+DO+bRiJ1/c
IM2DY/h9/HWt//+f9MljjPQVT7JwjHdAj2rjDsjKIR8T/8xbtqmbF/9ftnTP91hO
n3P4OcTr3Dbrmeru33DSgkbwVe2SyKB2HyHTABHZX7fQNPgO3+TP7JHoYMObtdPU
2QgW4HZcYlU2c0oSRHEIOwjfyZiQTO4JdLHH1H3aP5tl29AI7Fr/mQ3BFPe7Xdl3
q2H0Hx3IWtbvA5CGM4AYFqRhYHxv/TdIE2BXPtjejTFkk4KVTbiye+K9qM4yBWwY
6VUm2tEjVAmST2KNFTEfBFC9C0qLWY35+epVOHD1OSH+1KZjEzF9UiyaWFfpNvXL
cubb8e7Wrnnas9hGKLFFA1ETOl6fUTuos1O380Qx37p/Rm2duTLHkbijX8GqRY5J
VuGGIra0ep/720HFfUHkEjYwLyRTzy/lXs4Ko7VGBZ1AyyyfhCdx2me7CjOuIHn2
+/QQHCuGIhaKb6UEpEG3gw6antIIdmaVRQmz+bMeeo1dkbssF+9R95y6Of6iMT91
BOipbT8ESH9Yabg4btSr8k52OLuth8JwfH1lyHh6si8zTvK+UT/3jxysdoTQoOru
hoU21MfW6u+JiPWr3KkgxvC7/6tDPgChR40acJbpag18rIqG7gSaZHhRxeyDBJNZ
23KXlyNZhMUw/sF60uAya6akpN5xQFH7ylxh8oJykWQE/Iv1daxlC+vq7I/lLAgi
lpxQd35i+yWiqzSTVHVcJb9wR+IVIox2L12XH1mfyT4Qu9Rgoj/lOC86hznD5B76
dGs1fUGAcpmXSb2CRcPmAwiXkEyYAierxYmd3pc7QVCkmKi+XOjCzKGfknuQu9HW
hSeVMR7TQRp9sEjogsWysK/N+GYRmce1PcfCO1zA8c1Ul6aoRFros8+5RAEr86X/
97QGR3Wwe8sUb+MgOJPMSnfGL7eKz5jzrxin8gUt71m5LX+mpmMcamUgHBcDFXEL
ZlRf0WOXBZfnSwOFj+Q+rZEh5j8noaCSEN5kWtt6Ujj9bY4jjSjzCdrkr5yPsK6S
uNcPZFky7fJ6Bpodp4YY8x6Oiz588SWhJJImO8IvXtcFz4XomQg4JuE7xa5FirML
U2HmxEZoYKTiLXPik3HFVEIsi4IEhoGesDOe6qrTxJp8ykNuushanX5sWg5YhrXM
Vl0EPYoUuLKXdq8V1h6Icv5ALKpPIf+FEzXenoI/XIhCnzT3RoB6Sz698mRJKpZ3
PrNUn9hxBoX2anY+tiS/PbALrGX3++4m6frUFGx806mvHPVu0r2LV7TYMafvGUJV
e6lGguMgNMJVrtN0In+qgmCCmJeEyg7hozFlvIlzOEPvSZiEW1HcYdX/V6XEtFp4
MTF3xxIfJTOK8QOEl47KaP4rwkw6kpkJCzTHW51h4hi5hGqeL+8EugEybd8ot9HO
zcoMbXYlzOgR58M90qfIOecoaA1Mm3h/yVw/X9m/NkL2W8voKaxH9EnfKPP0jegc
b99qyy6aI4Mz96WFXylSoReQnabTCFMNOAT/O4ZKJ8109XQuPWSMOgt5+4TA996w
iJSiOl8rO+CKmiiA7lWPRBOUbtS253+1PxMnjmWxzvpXTd80XCflC2QFP6fbcoLt
VarYEPdQrQYFiDO8/XjUUcMvIr8G6Pcu94hKhKlpPSiCp9bsF/KIfRzVcOFqEMR1
qms0YkqQ4NcUDyp4p9XX8wLY8Fd8rJ5ZnqqtOqKSO+7Enntg2V3OpHIUOZjbmGkM
SZMTwf+ctghCvNGt+Gi+a4wY6JhRnCkj5Ojkmwaqs+wmG2/U//Sm917gUhbqG2A4
C8OjmFKOnIOw7N77tck5gUE6+d65YZDTQwvu0GTr/654O9fE91ZUWDz0+7JQLDSk
mlf9TfZWvgjXD6QH1b0JczkRK/TAk9Km2EhEjN2HgoxblkhZQflI0fypK+3vWNGZ
Ie8crqOFL9/HyLWwzOAFaa1Nr1jnN1o/qjm0IITg7TsQM1nQ/ix5wOqhM3mik8pV
wherg3Ih80J8Ta0osgrwpyfhpM9oKgcwwcyCo88seOFbA5yxXDKlPwWmty1Nb5Vy
vdWzq8kWPbrJ7OnNOXCzc9Dx271Z5W6yfOT24BvthMtFprHUg3hwULqwAytZ2q+I
vNfc6csWOA1sKpqIlOT7249VkBNsErk+FkxPYwNUtkd2/Qr3myUPtHlVYiPgr+KI
laMa2LwHCuoLM/elsmXNoaCGBp5LjZXc4JF/0RqaHiK9JVtorjoJSDxAE5/uJEGd
MQJzWxzW/NhmNSgSQDjfZ4Pf5yYtEPgCAC/zZVW0uDHcTk+1RjGeKXhwUlwWB13B
L9dsTrMvLpcE7otn7ujsc+5ih2fB3MOfZ6mbbVOMeaBK7Ueso0lfhfRjq1EUnAcV
ZAubR8dmNnKKFSBQAEVUlGPb/V0U5/QTSeNZIr65dOj7StEsDZb9o6LodvuKI5dZ
ajaim4Xv87Ji/PK8c7cAH2/3F0Uspp0am0foCOGY8Cxy3qJKHuN6vBtpJnZ08gWf
rBCbMNRTrzw61r8x16rZJhIHZfPciCOjt0YN4L4WQ1Iv07FRu/iaw90a0yTqGpjf
+RCu3I42XcIOlvkSnoUTid6iFED6FTt7g/4iLibN3ZJM6/xJr+y9AReBM6yR8eng
MQOVgFObhfRXX8TpZWp8F0lbzpGaag7kok5fGq9etlw1P7H9D43iY+IzAFDZz+w5
HcNjNs+xpqb8wOM0wrJGKrfO7lrP2KGpSZl1hmdBiiy8WEIfFOqgHv3HCKs2sZ4L
A4zNhtGQEba0I6xSAi4teIflNYQKJxePQoRf+5wrpOEBi8mZPgFI8/RXALsbM43n
IgslGxOOW7hNivZHywuYfPj01omRWSeurdbsKdlQat7V6nw1xladdk8PGT73ZDzd
HkyrU+DdiZhAnZioH3ysi7lVy5cMxq6sqT51NPS1shlhFFSzEMrUs+UlEvZ5x6sS
Xitlctzy4S113jgHffuzmA3QCfSPa4bA8agxfkzoN+Z+/J7SSTH/H11tkC5tGyfp
JUyj4XOhdA/xqVSoat9z2BOcPuBrg4wJqxrgLNWyiiipi5qM/gw3TCYQT6QnEc9O
uhW5090acmbgY39O0o943PmtV0dbLlMd/9rhP6SPnmz48VU0SwfSxU6onR6OtQSn
ENC1p04MzmuPKCVAvIo79drSDXFuW6yXWIvoZus3NEryXEf9mh5W2nU/+SlTcXwT
ENB2B8tJzQC4ZfStjQIOQ3NHYRa2MvPGpgZqTkiy01Tl4Ot8vF5XU3U5R6k2tzVy
yVjx78b2oOJ85YkLwsOVx6LwnAIiqptiygubw3hWW3aqUXwtOGyAXAGoCyD/zxqU
iEHwl+7jCSkM0F3pVDJ/XPl46utNoVuZLqyLgu7RZ9yqHHv2a2KEiAHIabL/OgsS
d5YYe8B07bQIzr+6irwAhiq4HYIq/KsOcGnWd6K5+zlg028jNRaaGP+aHHyIHGGR
mEFLAc4IfK8pspUG0HBAy4xZ5lfBpY0yCnKLbLaYd7yl5fa8pyfOXGHH6IgVBT5X
GPFgxA7H1yn+dDyZQDSIr8g3P0dBdeDVwBTUd0nD8JyLQANR9+JoYMiR85hgM+Q+
Jpy6K4mgYaywcEOudW+Ai/iBzzdw/XfY5DT918KHUz1Qe3OW4uCCnOtO4v5bvHue
yEpkBbMwRlyu/yKysuGadvMa+fYa9FMRH9MWltbo31ke3XWGDyCoulKS7mfEWNu4
UTFW5u/bJb9aw0/KuY7kgQ0lrKNnc+PYSsmAMTpL7Oba0qirs7fuLYrdNYYm+UV6
H4pi0Pu8zDJ/D5EzEXuilkEgl1yB21lG2uS/naRZnWDYrVg5fiIyKp7r9ZIcIdZA
KQo6ctYTR8k7golDkUcvJA9ZBT9wkuLYRh8QwAhofbFDF5aupzZ0KAinuSr3d16n
BtCy+jG3l3KLSslZWxF1to0paJ8b1T4/X0CTpvPVdFTAsIseTRUwzNK/765ZtcYk
xT0FTbZ74EcXsu1p4Thubew2h1JCDfw+3n1enbuvua0KrxRf0V29mT65oQlL1Wxk
wbiPQmUGQOKRHTq+Tlp95dc82dTRhoH9OdXCs/h/wr6QJKdnKQUe7astCbltOTem
ItpVhX+JnbEbUJCQ2W4vCAvxy69uwgC4cNEN+qO3d9vhttbbPISVrc3W8UTrcfow
9kI6Sq3gvM8no3EFk7gzBLSglnrjUm0NA0baIN7Vz+MhS1kKyTnXazQ4UhxUcYsM
9RxRHfmEASk2ovNRig/+hdIVJO7TsvM+vDzjleEVbFVKRdHIhx32lAGZC85leTSF
doiufQKpV1XjbS+vOXKDVBCU5A24ItrJeSBLsIlNnCiAkTnjbTvBNL7wvcrNTG/x
4CNu/aUyM9+H1FKb3sDFr4ZdzAcYorY+glinYLURxW2AlpaqG90yPi5pXboqHocq
O4sTSlAorDgLL8HPFuoeBYMrPtdBvwTxdKxVRdqoI/UVC0OxmgPZxJIHRHg795Mv
UFbpQvqC7kqts2G/1Uvqwk/iz1cDmw2Mhdcbh+xY0zXkDvRD0zWBDDn2o5jZtzyi
etHfl5hYNYBcBACj4svK0I8j1M2mXVBl72XMlVP1Xh1sUWJ0bEEJ9+YAZWQ0XFgQ
5qo+Bv5wQewEAC0/sX0Gfy8ZNq7uqKPbU7Dm3aEgxr9XU1j+cXw3agmzDqNM2gHx
79vdw5c8FBt8XjUmvSPPPITE/XMj1pmX+kQwXcUXRlH/9oMb++7UG+/KE31tVmR/
A6fUs0EuJDs+o5Otur3z6czpms/HeUX4hLzgtwpwYXAfLVMFGLy870cFWq1gTC49
CWInrFZR3BPmU5nEN6+0Hnq/JGHPtiQZuhlx5QeizCRXElmT6cU4J9GXY3PbmcVM
M+iO8JUl32yr8MGearewwYgQhaeYSR2qMFpPb2o2FIZtEn7Kcw6bt4Le+qNT0Nkk
sTWqKSOsiuEBALNjyNuPewcO+XAWNS7EWJ82BP8kd4+4BRQmiBrCX6F0bYlvlabA
wrsBM/LBahjFBqL/pGmyfFRXgyCiKjm1whBJ6nQ4GvnoiugBs0+RkZiZ8MX81Mk9
9ndewCkH4vje7LcOGpadBRo/+b5K/7lQ07X0MjbGqHpDUFC7Hvs2bNRBK3Z2ePgS
pQANUK3QaP09zsyPzqSmFyJIt9bfov/UUvwIjxguwFgQGOzpBwDyAKs3Q4eaOb03
sE3GboN6hxHKbFJ1WULrfrJYlBRuakD+deBuxH3CjStDW4ypPdarZKRV2ZHPt8D6
oWC41/JbJ8ZV2cppQb9AVnYlGkIRIC3e5sa+GCVdPoI6cjyyYTCHlbUp6k0i4Z0f
1uGHNKYAsHTaQURfuXIUG0LUjtfn4WCGDo0RgDLgOw5KuuKdYhKM/Eki30jJ8+T2
+RfHQf1lvQIwKOya5RW4i3sgJiUJ33Eo/oCpp7206gcNpmy8A6Irf9sYS7W3dN+T
PKe9E0npDAFeyoBTjAugk9vPxAs/8Ti1s47B0QTXcq9sId7z0PiKr+L5PUjDfaxE
Fd8fBePfu4eKAMr9U8i4ybyN4w6Q5whVL16Me1XfV3cR3GqLnneTgNHjEMJmQw/1
3uQ/4PPCxBb6Q8ib5sQB0VnkG15e5T+C9gMbYAoxlYs0o5dAnwX0TX3Re8d9DSdR
1a4BZZH+5X1UP441Hyojh0i/kn6A+d9BqUnrupjVZ55s90SFmdAtPeVc6n9nq8NI
jz1vMJURQ/HYGW8fPShZfvyRYQrPheijhh3RU4Dcz0CJzWVtg8Bqp2JzynKbcamD
ANUeK6e3OViXKU2IpKlC4+J5SEZ4niIPuR+o5HyC4aTLchKf1oixUkXFaL9E4UBM
u08QpsP6R9FdFhj3pd3of1paUfoWKv0tbnzlY1z3bDDGjcbjno3qTbyoKktCHscX
zdCsCOqz4OD6xJ4my8/xpiywiTr1xs0rSHPUizpW/Y8TEE7IIXM3DGLNXuGh1kkP
B9TwUTCLRmN2k34UFLClbv8CeWWkFsHyVRUe4K129MMoeXEIm3wqdCLZr+4q2lm2
SNsMQUtVFNTpM2oDh/cVWoQszUfaNTlr8OnM9OEa2sf1msoTKIFm63V4iYBIIQgc
+qVnW4AhFWg/O0zjWPtQn2RZqL3zoILyjFpDH6M53HWTwXEVArSwqR8Ijoj4FojL
Q9tXN7v4dMmUHiBM2kMvbfQs+EVCwYXCoJDvUqNXzrcaSOYQD+S0EE4ImD71lQai
nYw2L15g73//BT9R7vIIoCw+RFuvg+wiQqHKUqk3CB/42I5VLmX5TTPkIlM+36q4
8VZqwvWtqv0odXX/GDu+Q6skO3AK/b/jlQyciE30gPOeiBkayDvUz1kxzgFJifp6
Syks7QJHCoFTGzCs+3MPv7ud4MH9+tYPYS0S0vkcI2B0WZshpTp2yy8ColHLSwkR
3MD1lQyrhGmtuftfWqIlXVgxYJjx37G1pweHnNJoaFuCyQ16TQCjcr+vHEIGmnyL
TtcqF6nKc2iTWONHEHzqnAn5VPAxPu4fWSwD82SnYqesvER05tBVF9dNISkUl5oG
8AFXn37lRREPR0JYrhZJweLvqyyVRGmz9qSBEXvkUxWe7EmmPGGWlWKgpcX4q+cQ
M4GLG6zbojWzoRL71E+8dL1ua8RLpKxFrzoBwzzFmAAyKNyTu0TDTJojqEbSp/yq
NcbIeQjzbvqw4Nr8UZcx8EQgHq+zP0Dd25nwmAhVEXm5xKVoIUBljhFmvWQVoZhv
Rswubgw/HSqFVNgyf5LHev/Gj1/5ELXmDVZx8zJOaVK32AoCpmWbZrzraGYnUwRT
XkPZus+WHseN2ef2yH9Mji6aPb2DzQGQaGTNMI/Zm1zC1qrh/kTFjwWqRyJPpiOe
Ook2KJ0NhHx4iMPCMeZOx5c05bCy+jcW2n/qzbtJH/KUXz4rfNRYyB4LYt2BwAPj
FkqrOeKDgGuseNibk5IdhnHC0FmnSuvbarmP8fqULzKrmy3kmDjn9YJnBIlW7lrB
vMZpGJ+sdQZ2KZ2KkYo+f3VTQFCx+8tbPEzX325OCenuOy+6OLUjs+ReOhV9lZ/R
1A9K+UzdDf/IqfA5XwHa8DiOMzhJNDRQftQhw4f0CgfkoU3utbecMUtIwkBawHJ5
XqDtFefsmre6mcZpO2VbkoqZPP0vkmviSZl1hMOHNv1yEfv4TLEeb52BjejWTg42
szoRzKP4IESCeQzYawDHfRkOHOmoiCqSuREOi83/z8N92/3qirTdOGw4BgH41sV9
dSQuqJTjmrcclqebiZgqgXGp6OVOj8k1F7pInN9ZrwzYkRZPaHUH9QVM5Ke2hhP8
DjRwBHGNAbdF1o5PgJjNeHp1BG7T1J6N89vOOKp2pMXjSgqg74msxiiOV8rVqt+V
jgYGLSW6suNf3WprV3iR+64O3UoJzqc59dl6NwpAGD65sqNKgIz15xuqomnGk1VQ
Ev2NWfzomo1vvSfCAJ3zen1b6olL0lP+sc1zx2uesHu6u4GGntgGMpl1jhaqPMcu
zWWOEyIDNR4qYjoWILD9kkNjAiXEkQLrW1HayryyzDTystk0/mXzvpw1/70kSWwS
6YBbiVWyMauGBzVkLKQe2RkYKH0jLoSC2xDGL6wMF6IUnzmSY+lXW3Ve/tSxSJDx
LjY2sOApE+L/xP23LCXkoc9ZLIzMK1b5dvdYYxRlkMTV1BEIb2knUhhCRAcYNTV2
k+FNCtnmToqFnOQoFwyluKjXhcKG9yZZj/T+xXpwJ65VNhh0ePJyJ4OT4q36fGZu
dQ85PKhnKki7z7apDzXXgPQ6GXupvy5X269MaML1g96Byiks9Gx0G44G0SIqQybq
3zBbJqXmTyoqdBQEh8LocNyIUh2rsFcNl7ADE7SxGDDvwz/ibwRThE8oDCRZJkFX
lAV6bWsCXL/L7NlzOiVf37mFGXo2MwXb0q0vnhZA9x2r5+cWwMsTHcXYHkfs21NP
bq2mbYSV3u0gU02ZOQG3zc/3lCN04tapL1zjluHiigIWp+PLkndZP1n2Ys3GrJaE
gFZSG5uGdrV/SgCDqWI/K6BUQET+wkAhr8I0NwS6wI/Zh1eByH12TOTRyCKM0K7h
Rb8+7xUqm4zgVUcC1It66uRiUKLxO8Zso+TeUkEiDojMucvZmX5XNEQlEtIyfmfj
sm1pFpsMoF4iUIYE036i4jQS+1iTX7jYqoo71Fm4XVv7G6MR/GBWdAhISGK33ecY
45xaH4WoRDbsLBf1z5e8D87x8hOSgih4STOmeroNDcb+GFFirCnePWJOc1BdD3uL
iDl5DqvSnlHLQoEDbrrltkLRJn+QSs+aWCGBuWpgGkUOmsJpttIo+GXmojrHcCyn
eKex18Ef0115yZmEnpvG/oWQG6uOUOv0+O3UQNM3i+udMeYGW2FIRDggBfql4L0N
aRdchMBe9P05HvatBrpuNYpbsx2V9L6d37YGjLs3ZoPotEO0Nl/XMVm0HVY4icb9
egwreYfrVwiEfV7tkJjNtFnosFaNgIil1pGtLNTik8yxsLtwfvX1kzwSfspZqoZJ
kiKUGyBxMppAAQsDyElpk7Cs6GXmX8Gpd3dUSoLn4QPvM7zZ1VM5cnR6SPnVKW+B
EgA4GVujXBlxzxTWUx/1u0URCnN8+qu1qnljbqR38fNzvjCendtGGCoKav/tQZTf
605r4DGyclss9t0HJ2jquXCL2500ZVS5aIJ14anu0FgfBduIDixCVt4HYEHrviCx
BRCD2UfHoc/RHNW5QOb2nahZZxe81BLCfdcFwH+wD4fQVg/vQMHsSkgqAshEI2J8
fVOhO28qXNOJqMO4IiGmCo/ilY+iHqu4ZKyn2lQLQQkAcl0UX9mo6SfrnYExZG44
nToJW7dIFJVPwi3b2ZDT8XZuyHDRyqVA2CrZPV37bQ1Q0Y5rx7B2r/QXjq5wp3F2
8zmTa5tWZIKH6lZ/RjnY6SFGeziL+uY5w++CWTM2NOC5Rib+Oxy/v8opVQiOlobl
G6F48MvkcVauBGZiPWn8kco3tBUxxcdJ6dE6I/mQ2DKEGdPc9+FQp0apI1QhNj4K
XUTavepeqzutOIPHrmTbncr1Jcwa86iPCXqXpynzhwdY0/mN8JPu9bnkxNRO32CH
bDe+YiCgItOpsv/XMkGZbc3JCrW6iTowDqx6yMDCv6dfddDFJVj01pGMM+mh8B8W
B9tb/AHnqTBumFdLf7pN0jJPOw5+D8jYOgzvwMd0kXEajfR7cMW2IibdWUn4uCkm
LpGvZpSTpsLq/hBIFEPZJySro5gp6VkmH/WE3d9g8NPoncf/wbcYchugMnh3Sm8K
9jVzIvyyHRCCPrGMj+5cyxmj2dosSpzyo/Hi8GwdS5GPr9Tw/s2NhjWEtucK7o0m
+NDg3j/YQz6ZGdlBeDvj3FZaJLDws9d2Yj8DYJQUf8ns99IxK79WbpzOLVe3hFTh
StFgtmwn2hWhKrHQBoPtBjKOo05gfTq2flVfWMvMiJ/NRhLS0nv4ig3RAC9IzlSz
+e9NBEbg4/8Mf3KX/lXz8s+N73uiSEUVYZnqBap5DbyLY61aylaiaXAJY8VZFqAq
6oSmm7epMSmwehrQ+hw1JKYzQrFxgkfGTIEit0LjuQrhfJ7bjDf6tTfmNDKfyIvR
fvemb/BK3yXcPgcx8FZzyE/sSmzjubbp9a/rxUIU4jzCEX1K8QeqTXRp5YZWmLyP
tsBX+gK/K30wpMSXHmR1CLHk7oJZ/TZaTclZ40d3oe6hoNtQfyBPJr2uE1LZgfLo
OvvEc8C8dvSi6h0LfbVPcrQ5b3wdgpyMd9WLwBscT13f75UI4t3K4EhP+txyYSQr
Xo53c5JQYYDrl8DZofpkEkkxqmykIqsJc/wkbFlYBZS8dfNHQycDz2zgBJc9CWet
FTnxOptqnH8WsCnallU5rCTnyvoR/QNQ0Y7WJbRK5ukvuhoTVvLe13pv+Jv8nhWc
dl6uYkzQt0+uIxt0lST+sMhvbnhb7VBj122zkKlnA16Kt4OHSROMo6ZmZA+p43rc
xtv+L/T7GXBJfS2bMQBcG2Zxd/IA6tJlzdfpkMHqz/ey1v3Mk6qR6z4N7ZDJSv5X
m3MotuWDASIfjKlzvRyoy+QS1apXLawEzKAQticZDawt5mm7PAHJeuMq+asDNqxl
++CgUt18VW8g5OsPQ3HgcBiRkICPhfA9RQFyJsj/BcaycK2C3vkCyYKMq59zKOw2
jHy68x5jBKEFlpFP98hXBYI1vktp8TnkmLnBKIsUDYm4jBc7LY6lsimwTY2YgwkO
dgNfixYkfj2IN48hZoHOzfW+GVJ4/eVAgHBpRtpUEkvIkDNf9JuYbCBC6fAXzEb0
FJYPWVNJA2oSqqKx6N9kA3+HYfvEx5ae2PnS7z+o7D6HLMrHJQX1A/qR9MAg6VxT
OAWBaej7j+/4t7NCZQBkrKTeGQF4pi28nO1d7fPP+cRzmGH+DXsISJtle1t0CH7f
Sb05xHJWDhVuXcIeL4cy749hD/dfyxkQi68rF2WnJEj1pgTxNhFX0r7vP0uWAGUU
VVoQYXCGHXB7kM0pXICEHE7iBVSMtZuDtuLZmzGK3dZNAORkqHl0O0vPY+zXPM/4
zrW6yDp6axCDHGsRgzesL6hV2FlI0GxL4mLznNMnDdBRLoi2mlME7JOc8fsXvxV9
dXnL+VHS1LU9JIlqBWwb7AmgTgBRBW85w5A85Gkbf0/lNWJghi0sTiIRVYsK+/3D
sshTHytbfGSRZeB5PekVD+0rpaCunBJijM4v/gfwkuurMwwfqy4yV8uVV7nvfPtO
20ctjXJYqqRZQltwGORoq2CboTqjqMSn1LgHJ6iErjL3y3LC9wUa0gdRCcNsXLCB
dqjO9Iqb+lBrROyx8detCMP5V09GAdf9pp3ELlOlw79sbR9PYAEpu/zm+PCboyoJ
yKKJaI7U1Q7XqC+y+d4fp0cq7CMD24CflLBZxaCAX+aMz9X1Y5Vqw0Ll2LRxLWYk
F3rt9xOrJkd8hc0edYa5Sox0tU/H2WQhU2K3o+BugOsHHk+D/8iU3C0yr38nh6fa
CR5ryT+qmWjLs1mSCq2ryUx4GfagxP5p+xuwd7W3fUbTgs9x500tOlNOMkux8Skh
9yNDf8/EOfpl+08Qdi/iQ62NRt2ivf9DtFE4j8I8Pk9iEwKLSzpzgUTvgkRmSHHw
CUMwIki9XtbjS7WJznjEUEEfhwygMqkAqf0QrPdFNZSoHOsdyqp8EoJ/7kMCVLVh
ZlFAQmFCfVaxuKBtMWUxUzPVgDg8rHWlrjsr2xh+KUp2hsyvR9Eeo27OotN0NG+s
zs8EFqQLTXKNPkk+e7bLqiY5lJzfZwctLMmWBgWCjVN0AggCBFp6ZXRyIIn76//h
BanPErKmpk3RQZXCreoWz5munP1cpU2E9DSfZjTrGatuh0LyCeSySoR0r7BYtcZf
uUeXLhL/dxGMyIhpTHE2KbF+H3bfexcVxhfiVPK0bJo/1itGWrDDjMsqU8j1XWJw
hs8PWKvOhzkAMIg5D/t1jysVlPE6Cd4wd7NwgwP9x25OE1icCsc4pNgCgYtWtv5j
VkfpVwg13O1M5Uh3zd3E3BROB5hFoTizYS6vwAiOU3jQ27kbIWZN4m02LnTtn3sh
2o7X9jTE5XyeNNHX8zNeBxCQwFhyFfe6gOYvEMJjjmPEGVDVCKwI8GgQ6bgwMr+S
eG6iktCmHhHAgUNJLoPCLT7iu7BbgkUte5yGSTib7zebuBjtmYY5W2lODEAm0Z8C
wamupU8t9CofAYdFTkx4bxK/u8A62pZVxgR5ihdGFez7IyuA0cxxEBnU34YJ5Igi
hTb016eAjV1kQtwfE2LCtgHz/5XjGlxOYltaCVrqEOUxqhZNia5l7xwmrFbePdqn
GQyjKmZ8v+3j2VsrZn4B0cTgOb5sUoMSyFu0mcJhhwt4BMDTOgC6CVemKDEaQcZ6
Flf0tzGsrb0TZHQ6ibHOplPL1g6UvHe/sp2huaXDs3McgiPSyRD++ODP7OvNxB2D
ISYGC9Wx6EmJ1yopjsyW6kLwliwrbVhvZTtvi5EgVcb7+41Nkyaji7+CFwFhBCO6
AWuw4bMX4FJ0fIUHxzsiG6k/MiE3KWE2jN590D/FTYED8R0DtVnVxjN+2Tv4EGK3
et/g7mSPM1oFuftYRriiR8I5g15km0aS7otRFk5mUSVFBgDcIXf6Fgh2yLXtUd2m
CKYBY+9sx/b6qBudBg2jIx6GDuS9tsgFJfBEDQKILknyqklIREz0wpm7nAMmbOYn
ZivZhNbY04kM9jcygODNxXA8g3FCf90ljO8fF7bGozvK3NZfaf1TQGjr/KDe+2wC
EOgAg8QgXO4aXu0n4D3BWbVQapc8hZ3dGaYxgdBMVU0lahX0KRda2Fz6yOw0NsWa
ZeX61KOz31IX/LZ7H2mYxbHWPwyjz4uLd4wWD2Qr7rnodGRd2Ibup7rtjLgQDTcL
hr51RUnmhAzAMf9ILUj7G31T5OU+D8seuoFc0CD5K4h9tzsYt89J0eiCyX+4m0ry
E2QVHZnBeU1pe7cOlTut3mfyfyA/OtH4RR6JGNota3PyZsCK9hiUpkySltR5LiaS
BCvteEpUQC2Ksl+Xxr1lw05O4G78rzo8tV+R7DN98lEknBDesPR9Z6Sgmt7TEt8y
TmYPPljusBcYxyzDDKH+IniuJMfVd/niBzS9H647GlzR6VgyqUkG6R72qgTLeaIp
9II515/rxlYebooNepC6zStJ1lCceBV9Id+nYlJognZ17eEUw6xzNjfbDSPQ1+jG
iQyErr59ElQGXIAZC9xf/e5H7GY4SD+BSxo+mfw6w9OtIRE5e/aqSXIsn1aHqb5G
lMgLndQL1jcDk7BzawcqTYxfUNR/Kaes74rXZJnL7KCiVBC39OSTv5rUrB0E+zz5
6KKPgoHfwVCIfQaBaICq4NKc9Aud6PM+1gGTxi1U/iBI8OxJM/vRGYX89Ci0QrHX
iY8/z/JkXzr5uXOi3ZV5j6KbEsmZJquMHVvbKHFoOqaqTPMklFVoB/5UtAoJXwfA
WHB+aUijmACwryoP6AeO2z4kCfhCjdyCHZg2zvytnKWQbZ6a3RuT4F1VG4NXeiS0
HOuXo6kWeoiD6bTcGHjT+EHaldI7dsem+OJkvUJaKEGdIczFxq+4eDwPsG5VuQ1e
pIq9pNTaJlKCzMPG9G19f3bPGHyS9FCnigjWgJMvvsMMO9iAx6pgUood9IxUMYKN
L6U04aqjIm9jlSUjyGxPmCIGEZFigfg55cVu5xETJ2qU7WdSBY2pBC6e1F1H4ClC
JTuk97A8NYKkvcUDB6pso+xQhqjCTFhhknr4x/UuQiOy9kFSOsgj1rdHrDgI8WIp
DAePjoYXiXeqA/1jAhOrbbkatlqJeiMHh7wMW7RmDiMiXsyPbwFPYvOt3Zp64ze4
XnCzCR26zmRs6plS3y//oaauvWrtHEqgzPLVdLPrCerRn+wFYb/UyXXHk8H6X5XY
vLh7rDljPnrdEpX4ZkTKGQDGU7T1yWfD6tSOh5eiURjRF63P3XIYbdDxVPqBNV7H
ouYNNH1sacWEBHjEuL0zKajst9GEV6fa4gYev531XB1FSBng6I3weoHj9tLBniqR
qYDIrvkN/jBWU2uW9Fc/ka9ZUUiONMbFdLpUgFqxsuisIhIeL5FVsndBNpySNqZn
8MzhwmP3aEFmrrhZWLkebXPAgYFv9VNgK3NiFq+kctZjXiy82he0Lz5GKClBhjQa
kUg4E8RghRyga+ivgFRAlBxMHJWy+2XgUSdhn8rP4jZptONuM8UVJy4X0MxBkOhq
AxXWoOBnZ5l/igFILcbqSPuh56uAhOIl5hIhKkf8xkdqu3C37jjCTeDH8+mN7r/U
8na7SrtgZ2qUPKiJTKo9gq0YXreUBEc1ra5/g8FzoVG2F4ntwwhpAf317iWkhDv1
1ElSAJIBVEjD479I+R1uME+UJi1CpxIpvlIYzubXqkfaxoOjl/o31U+CA8nmQ7UE
0808dX10Hi0/Jdpn88YS86e8MUIfc5fJqaqYvw+XSu87zIwkpaQHPz5pBIO4W2dU
0KUvu6Rf7AzIUdWgi79UK9M3/tIFTb9xYhmYg69NBTgJYJ8Tno33mJg76wsQ0Cv9
cgxdXNHe7kn1rrAv9cUtOJRGb8Ge2WegQTiRcuaA7J9KsNIU3iNqCnxeovaxG53T
4j7bxbVgZs2O7W+YjJbIsv5aSALStz4euBvUdNzBZXqSAQD8TAI802GDk3+avCu4
roa0akRTz5pTKNdSEHImSBwz+CkdEL8COxEbkkshhUTPM+QdRbYGAcnOSKiMjOs8
lI9/gIxE1tOGGJ6lp5gf57pz7lvnqELmYstO0wgammZp0Gn57EWiJAm5JvTilqNK
ZkLtNndlH+klR4/bf/uKGSWPBD+CZjynAPE5Tsmu4lirnQsryLEiq2Us+1fHW8dj
w+xTfatglftE6sng0eGb1RGhn/sjbKqMzEy0/b0GIZ1gG8xLoCKMLU+CLt4wrb9Y
aFg4pZaAiMknwv6seJQtqjT+gGcHXjgHJy8oxsJQQNj2Ti8Dr/gJnOlyB2XpSgrl
OeQtbn3kBOtErJm5yDf2YT/KjunMaMsbTtcN5YpIUbL60aYqnHpPpz5f3n09CiZz
qxSiyzVGmfgjNks9mVZ1Yy/gO1VGzdfXKDZrBPNvAkDGHQQcV07U7Ix6Lk+1qZFB
Flaq90vskq30PYtV54O4HpJrWdOTMPOb+bnCsGm0oWQSzxiUPdzCgzn9JHi4ufj+
De0qKikTaYzY8zSKZqxpvZ3yR4hmTcSa2OZCve8Xf19XxSpo2lhpoFQNK1fONA+w
ZSXvjfi3pO3Ds4lhvCTX6UT730xYlOM8fx01rRg1N2XnFeO1lO8cQgz0TyKp40py
Lgp50WrXnX2xTNGLQCY/Giwr6SsHs8t2wB4rilZ9a+VDtqJ/g3R/oDcQLv5F1in9
hxIiXieIdEomVvw4LW0wxyGD7b4qGHuuGJ9HrwOVeKqF7yt33U6fg1TD6K2tzLxM
dShO0ufWKDyUqJKrbzLqQPQoyvfC0fsvZhx36vBEIjBVs/YdZxOz3FlxpXHx3lxK
MntdiXHKCjxP7RJSWDxMkk6QrY9zFtcF1BQkuScAMk9HfBLQTaLLecbqq3IjkFj4
hw8yRgSdTY/wXh5P/UY72Jx405FXKUln8ALFhcI4xcG+bIqBfndmVKoYTulSXK4g
hBhc28qbX5NzYyxMEnJlDuIml6JMXnd6qF6Mod0OzDetgP3m2gD7v8V1N9ycTZeE
uXcvps62fF27JstZV/onDrrcwNi0zepNrklN9ji3zyXohMJ4eVZE2eOL47iQbMGq
a66PtBXbWDd9q78z42sM+rwDbWtO07oi4oSWExewjEHTMVrbgCNcKZ1UOTbKlnQW
+leGB1ycWga+1AStZ2vlYXDmI+mECKcH7kKF5vEAUk/yFJSgA5jl6zyJJOSEhPZ7
KAqY/9ROWUEckrQcutZX7zqDFDdENQTBG0qFf/GnxyfVlbReACVKxe8y9L2enGxo
newNCL3uswALD2irJNvzwj/E31L85LirpZf4cN6XNMslag5wUNEH8F5akcpdEHp0
BTNk4DmGnlHpUWRmPXWykWOqgUEdBHAwJ3Zvmnc7vNvLcSDUGs6L9HEEsFgOelu5
/3rP/YTSIGT34uNClzTZAVUKZ1PSsBROHCPfEVLnmYiFoHNWbiyz5G7exGELXVQl
1Wb36CEnKRDlPnupkGOj8YTJs5qKMFkxaf3+4KWUvlfZXv8iih9eSgK3PF+AlN/8
b+cxJAIfykHkZ/HhrWYBQDSq66DTd3gUzDPRc9yti7dvmw7RPW58xiZFu+wix26E
bp7Bl7ZvYGVX0sp4U8ZH6Wsoiz0mRQKt5zlb/ALmY/Ci2Ahc5/7ssR9el3OBdGe9
sex2Umhb5Op1MfgrrF+w88yEYZZ0ZkysQCURIPVj3nukxPuoQvmxvpjwAfxR0JqW
7pyLxARC9BEphXZRyp16WhOTGb2uRd/CHwd6+Db0QdLVp/PwCzNkFas45ihfCU17
2LPbixe40n7BY2ADAWiju0okJQR2Y13l6gt3nEH0AbvPBuFgCc7T7QEKenOKnEmV
cPnu9CpF4xN503rJc1la/bkBnTik4xqg0jJrkltu+r3eITe6tiGEY+STTLXwu3dB
QPI6Ky9jQnitV9XAa/eLrxy5TBat28jCUj1QyPdw8bwgBtM+K7pLd/ZQTdZiL7bo
d9NdgMe+KqLlc4pqOsFY2x1KdFH70jXHDiuNvh4eMS2RUs1M9BdVwpvZPey29zD4
oCtLNNETt5PLnCBWacLDzuN2odjgrEHdqcoeJzXhnxj8mzRrmEniQ3ebk+u7W+zW
5Q5pfp9cr8+5d6/MXwA1tEfg12HO/0+9fBfYjgks2dhd95HULHy/Be00+OWIVknN
090vvTS0uRiaEKaHxsdQNJWXshwcwjnVOgaPM7oDj4fjoZvD9Ab+ZP4gpvE4Iugv
38RvHWgtc5AqJXFfg8d78XHJvG0H/PoUGoiArmQ2PFGJf54qBHUWvukCJCNtnL6q
wo6RqFZufA0KXzENmK33j8JQFgerG27UPRD/mm9xWhD0IKwdC7bHko1vdwC61jxN
syw7Wk6QR6MYyzzgKZ6zLgqUfPGzlgdRW3AIJonXolKbzp2eVHX/w4ZEpit4sjTQ
6jf4boZVTlRGR3dPh2jOijPBDQWGzlCdCdygAYdI2bHZ3RYcCSMFO+bsZ82zckSB
V2Ls87BnJCGurKGR0kLZv910noxsOCGr/nzzEpjJusj6BQWd19vFjSvExsOS8+X5
Eaa6Fb4EwhqFsuEyGG++iuFi41UIRT5ICTyIt+BwzkeNFtJvo31Tzr3jouJILwdp
G/iLwR4dGidTkiTa+5WPOypXHYo25lm47agREUGN70Pw2yT+JdjkSna5tRIfwFrz
wIHEFBe9DhHJ6N+JjVRHyL2MbWv9sXc0Z/4KPbdvcSTMpUKxocedGBRa+YQlGWJG
SXIF3p1BakwxyHnkaHi4HqyfJmQobodA/MIK9o30ynjrIL70hfqbO64TgR1BWi2P
fyJIRZvwrGcpdwUew9PCCJued82ftHU9a9DRHUmzC8ovHxpveTclD6aF+2Tf8BJ8
E5STUNVXIob5LzL4oQYy8w4SnD/ZJZYU/ll8gt7NEATDqpxkLVs2MUmps7yVGZtU
iOo85/Ptg4X+RvlAyT6ho2CDAWna1M1wn+2Pl46NfmoI/p3yNnd/HkixkKMgP0kk
iUf9+vXb0TyDMInrAbZpf/OB2+Pjfe/vpE5OikNRE2Slev9SJvNldNsbGUIRoyM5
dxejs3AP4FQJ6Z6L0OdhL4qJt94UwZuW1EhEtkAS6LDbzNyQVsfBoBnij0XAgxYS
7HobSAoeh1MT5x10MfMuPAmIdEnHFGwTO1MpaSHz9w2DN0T+pdIGJCs2FrzyfCoI
Wjcm1iOCVFY95xaojJYhL0ttzZZs1C74CLNmRqlaJ3O1MCgSxZDXeiUXD/JqCiLA
BUWgl1/PGOMRJJ6+YVcnejaIyi7ImRwMm0emDdvz+pxdzjjoSXYUgQ/c75ITfMG0
XRD4tmRiHKUC/R5EzIJ7TT5+aDHc0zH8h2wfZSvXqKOaHJ6JWEhGBTqRnP1e1cef
7C4DbDyAN+G3cO8oJOex1yjEcPSCuCDN1AoqemBkV+mCBNs22a4hXfdTqXUr4jYa
Zd6dxZYwiXrLaWVJXTIaXP5/DG5B5kqogqA9Fqlnrb4mOY41NGl9F4rNV15d8SpZ
15d2uLfuYA0Y84c5IkkE1sc0X8AFEm/A1VfTyGtYqF73OgyqlyH7MQQqOfutQa2C
McBmzWl3DM1JwS2BAczgrol2phD3reEl9uZWPf6tBNLMQNkRJpZzWm48wT5s8cPy
uDGzvUwZgiusitdW38RgX3ZAYz6u5ktLUJhYDKtSkT3n5gKJ+g1Dn44HwueuJ5l7
X1H8gJcZvqOB+rTA3Ovh96/pNwuoWo7HzuAhNDiT0624URAvNt23QhujuIxY6oJ6
HC5pc/tTM6N2UhUdIpr5Bf2UIgYIm9NnhoHsS3h7i3palCM+yeoLBEdMo3rpUvUz
D8SLf23rMWjJNj3EEyzOSArOA1nd3aIIdoKRn0HhReGcXKxIAWSlv2lEme66X5GL
slQB6vQU5uOdIWnR2CQuZsYiKQE6whScVscJDsfndxUl21vKzkSVFCsTsRXtGcsy
V5gYnh/9JU18cFHqdrMG2ypSHNR4DIWV8b4tk4h54NViSCXHoijRrnNfeDOyglZV
TWddew0wyPceDrEAugnzrPZsjTqkAlOLNazO6XCFWvjKen4/IXDYwnkA3KC+Da5p
YSr2KmBJKjvVVImVuw+FJwHmOpyO6T/D8oGx/3TWHjVaU8ybBx+A4u+i59opVTUv
HXVVrvo8XuFoA0BF+km0xMhmr6Xh6vEzzQa9brr0FcRut6qUUaW87DNHPEc1Zxn3
rhAr8bdL4E1K8TAZPbNHc32RvqlqKvPeCTMRDGH33hGJ0nPwN6uWFBQtqdrkbixp
tdfcd1+n3fCD5mkLLrNdM+O5N4H8WEpS/VEiXFBs60Mw8H1tk3kkwz2/jBk098Sy
5ejzPJUqB0XMtJvYBeOdaGQvF7g3NNHfJLdKaRShwT+mkXGxLGEc0qd7uXv0/q+a
d8AWJ6nv72rCXIUWuu+ahY+J5qZz9smoY7pCd4RthPlFwqjmHRBx3PdaK93j3KF0
1yqvEX4HguWPu8yJtf8Jd5N4X3v5zfIGNU6aqwgnAuYR4DJ2AhmIFuPDPiyWzLvU
wfZGk/slc8BMKYMFTwTbuSqNgaFNHWziufdRPYdTzzGZq86Od/RswSJbbb4KWlUz
mH7BMUUzYHKvAEyvMY0kiQrMiFnHCRsW3tq6r+OShpHOnSjpW+EALrdvDi/lUbhj
ZZrPesRBgTRQT5NtNL8cCiTBo7dJRhxN7bpp3SUBVgeZ4igeGvfQRlEMwpCe4ugY
efJUhj42aBFPLc+PJJnhufduVYf3ipq4oWol6o9mPcurZXcRdOwvr5DRUstvfhKL
EwKHeGyRqOuPXsipYR9fNEGVN7TEeJfQAZRad5CDKHZfkr0Dtk930EobiqrUEDPj
mS8AeYVDFyT7zqD/q38Cdb6QOUzTLlJ1s5ceA2Z3+1ESgEMA+BVqjFCIaWCt1IzU
Ube0yJvJ2RZTHBCVdZne0RqmsZVhXdPBAC/5uR9FY9bFqSaSIH1zoBZfBjboOuGO
WeGVX+jIFnUL5X7E24g2rwFM+acnpEMfmBJgG3bYUxjF8qrxcRwcx4ouNT/OHsH5
bhZpa6ATRdwccLc3fLf8vhQ5zHqmW4qVSR7oiUX8m807JAi4Wcudl6TLmnSgorl5
wPigKtw/eBny5IVtAM7qslAnWoVwRgSTrHbW/Olkv+YEEX91H/z/x/3hTUztGhmk
Po7k5/x+YbnbTkLmitzMatHQ7r1e6n2ZO6DGKe7NFzk02tRJn7YsZ3ETRWgRYEkn
0C9KLP2xKhtLgARS4/e1DsPKYtfFB0jfQHBg3AxN1jzrkTJ69yjSUXbQME8BZUPN
QD3CIFJk9IRgZcNC4DYvZ/KDCd+qn6hBs22s4wXK/stM1DdAXM3sqTvtTBrigdCt
OjX57a3xyEzQjBZ4rGitP4s6qj6YlqkUbS5/k40ChhlyqPaQErP42s2/477nUj8b
jeoyyUn9bFCm/I7o+ZbsQ3sCcvKqyIagY2dhZ273GFhRyDjOF2xmQgBgeDl56duq
Aju/qIE01u35dhnOLm+yxIlmRilJcn9m8BEnQQAXRoz8LREvqpVHbpJEEqU1TtEy
aLJvErdzgxUcj1GXfaOtmIcFBvduWFGHEQM9EpXF9sIgUXTdJ3LnZCd+HMCWZkj/
T5dUMLxuyEOsnyAZy4X+TdGs1aeUEswdAR8XLUitN3ykb5rpi5YGSvUoH0gRf5F8
etHXvbXedhyJ23F7yqMVIv2pcGk402aeaw8iEdEVipYSd2n3gbSfp7L98ckcMnnF
jTGps14f9xsYHzjRym0NzqCc4T1VdwVy5zntFYebN5TGQarPBRYNGbm/STMPHQBx
XbAl3OlWUID7pPYDW/fLlqThftoQqgr3gZM6YIc8SE+V/N2zGXlmKYc4hSqcvdGX
tGTYyMxBAQZdCh6i91MCV2LYImLrHsffp81Gp0eOLzFYrHskFutSuI15cb8tVnzl
7P/v0IaTWRR+tQWQT70Ey3I3TstIDI0ybZ70mtJLw9grPlDRe4joRfbDqcfxc+mJ
X2F9QHSBtrFvxvAbcmv+1BsiIhHQMRuMW+EqP4BCVvOvZiVRnL/KlSQbcpRZs13h
S7vODF879y6uDO2GmSgL9mVNylmbTiAtsvb/PmxJ5BtcC2N8cJzTewiXNJtdXjqt
nVdZoepYB47AXyT0z1QHmfb3GLcXqCAcJEbG6mDmrlA+dZv2n1IA9ETenb3Ie5Fs
7wvBGtW0wUvS8sEcXA9KAd0ytw5rrz/N9wsyLb4XgNH95J4t/ySGN4Mpx4wfkLpu
7/59Hslpi82z92AzROCuW3fNIADmBIHysqjubYfpWlcvmghRYYYcR9bi/7shhTit
bwgEPQYz88xpqf56LSsnX1JhXdUJOKqNWvo+IHD/cBOIOjWdVLmsxI7pgeSnUZRP
sHabM00mcmTVPTsEU8198zGi0VuC4Wo7aOtd8eeYGW52MiH9N1X7mJgphxQJP9/P
LoZ1zekXUSfACiHlWycDD2YhR8HfAkh+T29jOK8dlzg2meE9TaKty4L0IVzNyNRH
am6bDehNw8/oCj5CwXboQbODFHsR8MMEz/laGF8WjSlu5oohxmONQ1Yp8/K7kBZ9
1uaPzn1IJwEhk2R5iTYM3MpMg+rUM5ss/dzRgo+0vqqcKbvyAdevDu+eR4A4MTgV
oDLLvIM9BuGCqddTn0LfSCZrP7Eui2He0I+PIQeIFUp91Sh9PxEzJcB4trDxFCYo
YC80CuTrPLhhQ33v/VtuL/1yfda/kdEUjI0fJqcOpbZYFtiNkJH9r9+w9dUjdywe
EsbJSSO0Yxs8J9W9gmqgchcE3m7HkHJOmcOc6KTY1AsQdapTufy62UFe3t97M/z6
6eJSZNYNS7jweoUOLuEUX1kR4aXvdMvT0w691r9TwHWWv5ZW0cbiOp+oxQ3Rzprp
Pu12bo8dH0j8SZwQ82e4rRWyw36rO3DMHOwJtdRm780E2+KJ1YtcYo6TUMqxCY1b
yl2gvQ+TsstyHxMPTKVDFdvxSjkJvvIFsL1P/b3bvs/lNM40JMd3HH69/ruIhA/L
KTkBgVwKvj2j53xS80XsJ8pw/U9kpJf1keOqWuVH7C2zgcPCuhm6cIZRV5fffATm
cqfIK509UUWaFhG/1zdCyM5FEQQmWPMzaNsCU5SiOyI13QSnADryd2X3WhXYCu+5
xwY2zL8wp9lOxkL9df55f41JWl9lMVUozaQ6AKM15BXS3ETqApdm/+z8c6gTA3oq
/wHM/4YIj1gfJDFte83CQ9oHUfV3w/sIBErf1EvV6lG/bY1+XXxkNG5IK3ED9Z2u
WKEwH5HYCHaV408iwLve7BqIo9CLGuICYsgK9J1YO5SqKhQI52Oa6Ytdf0zjBVTd
AR5CY+Eu0J8yrRTbtn/61vVDOknaJtJRMZP6+RM2Zz+n42DHtiYgviw04SXwNaBJ
LY1vOAfnsvqgEclzXbtCDK7V1eRZcTfl4b3tCdc711MuHTEppImugpa5El5bCszi
BPUgAZPhORg+3gXyntSRBsIYji+lIiF++prZRV2Lo1Cpx6bPBm/yzH8O62HxT+vC
JanLo6QjZID6UXKvRpdvub8yB8QOAHZaY4+/FAiUvJtNNNCtyyNqcRYSt4ayBN3E
4emEl1AHlJGd6rwhqHAZObhEA7dLwGmCDUZlSN+zwyDf4LqgLlEaqMrDN63y5C5b
VHaCOHqnFmuMkO4TFOsLd+/EAbYwCcq3/cqsM97Xlx2xMCQDqL8rULm5DvSnpOZJ
B+u0+C6BsmplGUba0CBSpVvqpgCBImIZbOKwYMyAyB2v7VFIpcQkbasiJlIgQ84R
cJusb3ymz6OgVkUvDmynVLqem2Q1iu8P+329qbnlbFpKKA2Dts5R1sTSzr8RHaQb
D18ta31NqihOUaJQWxczKU/M2/SryW/a+geW4JDafGYYZ+Bt+H6VxN3JpthXnTRD
y79dQgI5SgwXdRRP0lvdpTB+yt+sid7TaPg+jnvk0iR0OnoWfkIRfae3Fxh+ls8R
8kBfoA6CsnGQRHVJSKm0VHFuFHYYUybUOy3HUR1pyvIBW0GtTsdng3Pl2ucqYKxD
g1GgBJ9x79RJ9ewty658cJ4pwcWH31NBVV4xWH117Ix1oLIJzCyc5W7aM+d4i2qT
u6Ncijs0YcdbyBf3+8acybuqJRoYtqSkR696wjrxD3l3E7bnJP31hbQ5TwNetUj8
3eD4N2tPabWuf1Axswt+qa8fUTAryVHT8aWFj7jgm6fdgT5hiDzLVrG7U/UPp1/Y
oIOILIqKrBop072SRvt7g+YoFUxwH8cSCz2IE6mhFokIgABvO41bQghuCBYsO2UT
262D53UH62VTZqm1pyIPiJEqjoml6koBjHEOiHbyCsBAC0Kpj9yDo3m3o0v8Isfd
ZlmHsVswAIviSqy9Lck8nOlqdbGEaGOIJpF6OllM7YanBjoFHiq3lUIXa1XOpoRe
L+gbynVTyo3THykiDJh9Z1y6jtu2fsqqcY7nJAmcAbR9TNaay3QYhOOngQaX/c5V
bbWgjzXzRh86D64tQ5HZgnTQ8Tts6HPI+tTQ6wwAuRdpPI6nyLA09iInGcCD32P/
nON6vN+FgOWemWsoeJI2QVF7sAsJ+w8R8nJHvwQH2DlvAC5sta4hjfatJWFb4phM
u++1L2kx9U0z1ALE+QCj5Ov7KVESgcrB9YKuywxJT8oebrDrlADvkMy2gromID1u
bO7i0LwACWbMZ6So6/n26agHnA0XhkFkSZwJkLiotIPkwgNdEYshVTIczq0Uy5tH
d2Dd/p8eNGcBonmhebR3vDDePMxZkEuk6rtZEtJaOHgr87/n/ipdwgkIgJhGHw/J
t0ifpIieycIGH0K48AIu5AMZFUdeasGCWt6hJF3jUrWjgKLeGBMy4DfyqBvG9an8
/PqljPAYhV4C4c6DZVNQeeTK+i1giWPBt5BDH9jQiVtRLPJpooEm0Viqh4Vs99jh
z7OE90oFK8D+2QEZxwfLXWw9vVOHakpL3dZ2a4b0RAHYYzG1b550gyFLVcfs2lXH
ztpiIQyCys6dnW3fe9NT131ESfs+IwKC+81JNGzIunNyVLadEEp2M9hUgPozSczk
M6oHJuO7y1Mn0yQ/8iUYV8jyLuNdRerRtaXmbRB6oM/sBl3Is/B9Lb9arohb+7lP
HtHoPj3gBNhQXdKU4BX6cp+CGSSRX8OFZqmN2bMS8KHXAMo9UiU1vmZMMc9xs8kS
T5wOG/96sLymnss8bLV84qVHy+gATsgOaiIH+e81UcEwTd6srv4cSEQEQN0UEAqy
3vE+RTLyytwxzGagjB46NK3vZ+As2gnxHR/40oUyH+uQTepHdKzMU4GinwWzuxoR
S6YNUFmhtspQoomCxCjtq9Ktc/tXEa0X/F+myf3J23lHnFWoDdX0yJrjJeNtAYn4
g5BGG0x+yOVtHEOkk5Ubz7m2/yMS44Fz/MrvZnD2UAhQiFMpFNyfnyYkPbifzIId
bYy65F6W4LWFJC4z8Bu4SeR4DnXqxYtIAWFbPDEWKZ3KZZIAA3LbDHX6GHZ2y6Xx
rZryGYpTiTiTbZzyrI5Y9m3IZRF16mTOTWEA3eBrbAHgeJQGBLwNrUIqQQe6ayAK
Mkjt6DyELnTUInJ6rwCdHTc44bkxTJMnGr4115t4hcCk0N5sWLeqbpVYnO677j7w
Wwe+heJuB2FJBJgdoK9cP/l8QfWNxQlNmlNSB7HBWy0YxRdHMAf2FNJ+KWSN46eK
GryFWpt8KNDhDIBe8YWsF0+AZOhlbUNsB2t8DVxbOvho321WhJvNFbp3UCP0qr87
0Cv/ib7SR8j2z4I/RTzGMGPW91BhTAfgHM9ArhbyCw29BXSxptqFBD7qPIaG2Ken
GdG8+jwux/qr2H+pJb6UoZbvIu1es4akfrU9QyTZ32VVT3mi5sJsik9b+97fRsnC
Nbrzru9B6ofi9qTg7eHoaqo5oAQoXkx6Wz6XOGwk/s9h0RcC/aT8/1JJlTnSlB5K
QGzoOsSyB4UxiAu+dnlsv69ktwK4aQWotM4SYYIkhiTjN1ZirMRIVD1u7zfpuMlc
ZLB6T5KCijUvvQRAsKGRxz0HeHOK9yvC0qbfQ5aexui8Jq3wdmdsAsM88+2cmret
Rm+5NQKyoq2M8LuRNO2uoG6P1/3hRLf99t3LaDFGxNTHMFCad/esBBtA03EujmF/
1PsxNSXVmm7AXMI7CC3JXnKjV3rVjsakNGve5QJq/vzroYB5ARzAlPe1gk2V3+8l
n1Azjz8v41P5H/rlmJTfVPHsaT9yGCmfYAXe9JnhDzPP1c382edllRuvqHVTGKnf
8ggVuQ8ExkTBpXj+82og2YUpn8ABiD7fWLXTdNhgR2oGK1iln5XyE/9my+eLqlcM
CdBtRhZXoEEyemUAkpUkQDXL+L67Yf8FPeOSOH+LdGGu0CPoxJrRWyZwqmy0AUdd
5tiH2aAT+RUwqUwV1OxtOCMK2H/pSy8YeolV38kP4deK4VWVllXTchWICo4ZeYMt
TcE62bGC4fGRJuKdJOlUZm1ULj0YvITHmBEHzmxueToZRiURpp4ChQ3OouilNT9J
+5rzgplu8Gly+AjihZ2ZlLbp/+f9rHKDgPH8/uSMiB8oaKKpdF+VmWuLpQiaJYMF
pOmvHg2+0v4V4dwvAgOkXz2K76/PMo4FUxEEvi3L6bEFp8fcleQDQejQ0ayynETh
hwdJoMkJ6wHNQUqHtmDNhglBPxE689qUvD+LdBy9iRVX0yJ4GBbTx+9aYpYwdGGY
bG195QpIGZBoDAOztnKjuS8qoeZQJETNHhvVioKHNlX0BMEFhHkF45uWg3sCY/Ba
teZj6xub8EPzrqejzEGYztBotsTZqvGfwBEm1O7xF4pcGFMiXrCLrnYpwm7paxZA
HcPAxF19D3chuhqOviBFkyYcJY7oIOiP4kknfa0hJ+8IiQwC5g8HIIZv4u49Ujpo
IHRzJHLeGpQcnqWn+TWahsvHzqDlDgZazUmmaK1RYTA9JTaBkbvb9ii1VRMoOqxR
3X+/pmIYyU3POvjjZoDI+bConguMJoccToZSw8Jd0BymkEEfr0JzHEdIR8238b+k
ErJMzFITGdt4JRMp4wx5PJ1/Lyrc0hgCXkUiqPFNL9yj62zHz9oky0GDpHdpvZGo
cT3Kz+3hzQYd2NGODHPwv09dmBmJkNEq7cRzB4ysMoz/iZ97OXvfaVCzOUQw8CwY
sN231+BVfykQk3oXjEA6KCsh+NcohJSrYMgYymeXqHYaEXxGizMBuXR4AqFJp2Cb
ks4cPDKNo7+kHDkI4KVB5KWxIudBQ0Z008J8K0Ssspo5WkTJnkKHcXr8IuvIHCXM
ADaLIAAFyVDcWcnDlk3npNETtTLwq5jcoKqESablEDP2PwLlXd7PCMTA//42kzRT
36IWCxylyx3uhVs1mDB0cqLoV192a2Q4GQesEcy+I1PIWncvMGUAkjQQWJg7svzc
6RMWgIfosRRRtczpsa1h9j+MncfIsLvNgbaVTOG7V7WtQZPQ/KsUwT9HK82v/W/u
nOq2NCzBgqBEPwNM5csdr96XNjGnTNFGyFd8y+q2QnNItnrh0r7cuu0dS4WAmMtw
xkvzdjTtNv8RZy2eOESGpV1v5RzGJEBP9aNpaJCk/FsM3ngjDiH4uWzr4sZYVn2O
ZFQN7NPnk4Bo7qn8qjNg/5lfMt5imjB99EtSJ6Z+17J19xEv2ZhjX9IiB5k9RpJ5
SZKw+ZDYyj0ZgDH9s6kaTmpPyq2Q+Q1Ya/lgTuTq17urn02W+1Y7IuGQVPEb+MdW
QySftkuccWNuK6leRxJUdYHiGlDa+5CL1/qHOM+Z1JACABFYwAbge0avEGoQhWaG
Iw3mtJam1w1lIt2PVrKQnHF+hOwvmjAnQ1M7qXGDA3gV4vVbY5enjJEqh1+l33Ao
A53bhTnEPnIuyW03qR49PO/L6Av4eTzkjMp2sp6+0Gmq+ndngUpKGNECJOFFmcxi
JnDUHUebRt72Xx1wnp6Sw1H/9WppMpowZkvB5zgvsjklSjrUxXj18nM7QL94l21A
moosCTEGQbkmiNHkzn0FgobO8rOeo71WEZDfjwrVR2Jwct5VdBb5KqptkdQ5htB9
QKrPgfEIFWKe+6GtZfxdzsIhNDWTzsAFDqn+kihnYUd1YOegLdINkqtB7Ki55VM3
QOH9EQEolVj7TMAzACrB/Um2HFL+B6/rLWgCEkYhoUvGU0tkEjZVJxpdVQf1BV26
/jcAscGG3NZEA9p9zxRdqDfFGnY8GoVaGrXUkdOWsxx5oM02/hauN1cYvALs9AYy
WWqEhiaTK2KHrR3r0XU0/8wTOU1JMM0dn7+4AFzwn19eX8IsZ4NZ2i17oTuUQ5Kc
/Y4ochYogcDwKYCKni7LgtlXQeZIMnP76exx6Vi1lRFBABemRZd3BedbXi/j/tTo
HUNIVmWGJSoxvlvYpbebkJUvlxmHACImMbmDGxsl9RXl7eNijovHzd86odbraUMD
9UGBGEV9m6CPxS3WKgflEcVRiF6w+TaIxBN20/lmJs5FSOfGv2MIuIG8jv6eUkj8
/ShwyMbBMp02s5+mFCp9FsKjsZvVbAxNJ6Xpwc76ORHKgxetCzoU06Eu+kp6ArVF
OSts94eQjD/mXC4piD7IXN1Sjo2a7sUoLRnhjbNV6vvsqy+OuYrwXB+6aVmOpAkY
6+MGF0/6Y/RgGgyl4JXcb4kUXqBuwrRQvXBPqQTHh3KdQlwXdmljud/xwaqbId2m
tNYPVyd1M0dbveBwJSTmKF2tOCRzunExFLIVDSpAYEU4VM9FNSXvJ+5B8cREU+uG
bi947LXQKFe+P0CFW7JvvRExIRpmMFmqucZnkwhfd5nhBJXUIw9m5cZuRmLxCkh9
GX+XaH0gA2wqUyj4pNJk7+jTilSpa5Fp1rF9PNNDBzv95rA6KDaaY0fnu5H41dpd
9cNtUF5gAFNwpvjZTqbOIYSRCslATWt0ReGA7iAufKMqeDzXw5VJR3FSAQwT8JDY
i+bhXKcO/KyErcoIDIH34sGxb8VGodP6QfyEwv+w0a7KVXarxJ2SyL68b8vYRUJi
am0d7AXvxDluJcf1TPiHQMvB3/p+6KVN7E45TV+1BcmagRDHFtWw20SGBMLDZwiV
Fycr6/6TQ5SPpxdQETa+c8MwL1DmVUQ8kUwg5oS74UZnZIxrsAFdDhu/BN2GxjU/
tsgy/BUrrzaWH8N8yhzqAjDrKHG/TOmChgJQV5MXAgm0wemZpvZHAEy0MtgZtsQV
VDhKEVIVNeyujQOMKeqIDNi0/iXG5RRoNdG07Mv8qui/UTg2nIboWMNn4r7b9Tq7
EXiquR9Tq/27jCbABpTVEICxCXDCQb83CBckFzs2qAzxEgikOL0/nzzviGq/Un3w
Ef08BvUv+MEf72pir3B3TUc36v9SWqx9615JZ/Ti124la5etUb7rXU7NIFZ09b/M
MZ1G7qXk3Qsi1ISuZkC/+UmcKDwLxXfki702d3KniNN2BfxFy0BvsdhVT0+evJ2d
5fKke8Fz7JknrL0UOr83SL2fV7McWTXLxz3Xnj5BmhokUw6JsfTfkYWugJuR7dpw
yaPPsP4KpRI6A+oiyb6zlUcZ2ZlGsub3T/nLd6o/9N+ETGHpXHc3tAAQo3beKlzm
MYMmFCulOaoEPjPFnuJg3OvXNLzcU+rKIr+EL2fcA0lVjLA4BKrvL1szCPyJRkxy
p8Sd2W5IIMblY46av22XIhm5K5XIPljksa2BjRNXIbL4YTuGHu3jDkf9tisTuunC
ZceV9lopHGLXWQUyRtNKYsUKpjSF6DIGuQ0dbEG9w4UV9uoAjbxKP59vv986TiNO
38XSlXM6IT+uE32xGgP47dM2H5VylqMJcEj0mOtPbTsdNqTqEQmn/d9Q5SoefkeQ
xR48eYpaURU2e+3SHbJU0G5QHDxc303R6kYkxfiaLtS8p9ljHrT5MFtBAYxOODKP
n5MaVAqG2SBZQBLVCr56ZUzYuC5zdauI390Hwy+VBKMjWIbwr+HF+/OceDPxJyDt
cdEuAWnVhKBSMu6ohBsRDyvPtpW9IlTfMPDoDc9+NNojAlUzt9WGuupjSaQHAIoq
tbx84/MGVec1GOEw5oMQZc/ThytNWOorvji1cUXGtaMqDofX70miheUK0fsLlBu5
qOmNiPJfxah1PSJhZTO6L8KVhxK/y32T2fNKwTWfXqO+9Gyw2Eok01ifoJ8o+3yb
7HhDo3TkBEpaPB2Y1/FjtLApBL1IWWyEath3n90/T2u5IP3TUBMrXYnYNvpIK5sJ
uiXOYvb75nZxOMuxPyDtD0Ks3ngoDy42448LffvodQjSClNaL2JwWhnWt8Otjf/A
O8WxNEAWUHh46zcNju51FwGjGZYP08XQ8Ov25UdRmQjmrg2c8cjDlq/dWh+myuSM
ZGpiMk6A5tGd/Qp3HkgOxqwQe/W7yDbvRdgKyvQM73wZtcoDQZQIpyoYKjXlHtzv
sNI9E0gIiDGQcAE+qBpPvDkDuG6yGtCd6o/WU02gDVyYYi2/JLJC18WmeCLXZRbq
ieodDAs99ZfOjmZ56Mn2GQxpYwMqzMmsfAJaVvMJN7K/G0aPfqsVohH9m3cb8hj/
9OiIdVtZus99Ep19DoQZf2TZUDebTU0X1WsOHsUA5gSTAY55Gb8hLX8zrNc3RQMF
V90JaePxw9vjVLP5cy8yhGf2DSMqSVxYFvIyE8K8lcjDZMT8zj0USM+TzPLpcNT1
szBLE28zlxSAdZOzabmNzpgLzChrK8/IZ9uxowb2TH2Ix06AixUmSeA3fZudJaON
H6WuQxmpRRInC8KRXjRIa15LG5ADadCZdt/yGoU+FJcEk1OkSrnoeqGb1VJ5v0fZ
AsmfulA38HhbDXvyBID6JbZGFRNDsPECsKpnCNa3xJgpU3tJZf4PqSjUu9kgrpsL
ObLFYOP7XhJqEmOTbLWLK5p/Bwk/17Pcl2SRbBplGwCUS1v8kxoFbTypyMVpA2c2
vVtuV9PNf4g7xp7DO97dtG4QlqOx8g3edonT9yWda45aJt48dF1Uk8hDmqyLW7ya
ZeiB483utLXpgTdtgS7Y7xrJEMD/30Te+4bFllzClrIYCkrA3qYwWyeIhqw3pcLd
iWXCl4LW1DatbIhKXnd2tRNDiBjK5K6m36h9oKlA6aoVed6jyeC/G8+Enutn90IH
6dgo7kOqIHuyvEzXxriGXK0c3pFtwQ+BLVn/JcG1pYnfHkmqVQIsC19WkDGqGTh1
7BskSIMwXjYlfXIVV/lCgqmn0t0qQPBNhZE3B/wREQWDsSCkQRvsQzd8gb4nCb1F
gcPq3CHQsRc5c6GQZ2jmE/S8E9AK1g78YBi9ENPnXD+FfgeLPOoC21p0DiA8F5R6
2/xRXHyLB40HLm/lXZs3Y2R4DYPcYpw6SfQH3c6wkwpff2aysFVAvmuA5EOdh9jc
KTfpyXQrLJXjyXFNIpmIqFzxo+jcUeHD0UQA9j7BtyzZU7pmjCJHMyRnXs3D2Bd3
hjPzOUveJWsTLpuBy7LEispgXpi01NJuaUhnL6S2uZeIX5kDdojKF28wp0q0uqFn
UsxLGLleTdNGRYuvl0pwODgs1YbITrOqE/jPUG6m02EsCytp/+Xk1xkfmXIPAQ02
fwuOJd0raUKzEdnaY1DudbTEXgQzWzPglTwTycM8/psuTCW0VNIXvblAdTTT/BMX
QyFYQu6FX41AUM1oZplhNU3cTdFL+Eacj1RqYfSLM9YdLvxz5XtoZtnkICuu0k+k
t1dXy47T6cwVC8uWo4lZ24M0xWG8gkJHLhlFFRFQLgE9zMMewJ/72FlTOwc66Bk0
mrg45V+IgxlI0LnU7lEEA0FciLiOB8Xe8lCcE0IHChXDchwm/YDK4jjaDvQMpwuj
UYUU8EqCTJbLf4JI/EGlzShhM40F32dDOyFv1Fr55yiV7fSxdbrmMCM+Y5mxAQYl
ktO35J7VST0N2njqzTZY2UOWjf75qDLMMCuT+1tWgtldqUyUP85bq/6DVe9yWWCF
HZV1uxdXnWMettZlEjZd66xpgLLje35WWYai9bDFrHGhiLA1hng+zhUYZ9eL6j/m
5jATu6f6IPb8t3Gw060HFT1oYT2BRhW9jNYSrLalzeSxA7IzpwVWdHqy6UsEfp9y
K0sEhv8KJsiumUG2DVm0qGG4AltTQMdZ6d4vT4RmCAvj7Kw2PqcF3D79yP9safRd
CpQP8XcXIztIfOlYTpcYEiacCn3oXB5Dec8wp7YSTrVw66kx37GAYNf5lUuWTKrE
oHUKYoFAkxxG4I/73nHwx0/FyBIdeBhph+lGLDL3ASZYjJDV+vDObxEh68q2Dg6q
6xXlApAe+mp/8MyYQnHhwj9Ta/SqrM4j2xF/2ZYGKDF4wjvq+gpjxOCmcFKWeM64
6EkitrC4ssZa1CR3T3z8YX60E7ZUklu6gGzViTW4bYDCno5QpyHOJl2eus3iBAQb
w+8WS2ygnwGHxZBvK9Zx2ZaQ/8o0MJJuqEurjA3kObz2UqpDgBxIASEKTmbcMcrs
fWQLZWC58D5NEykTtxtKeq9+aLm59yiNwS4FDj/1KJoHT7tC1HEjZ0yKGDRvS1gs
sw2gPqZiVhBTzen7hlOlk67KdcpKW/gAkMoxCoY3z76W8lR1k7QN8dz+y+zY/r8h
LBZCnQsmMPRxUWELXt8+Vsd7w7ylKaQy+oRxQnx7PaOFznMFiRmlhTJdhMdoQDvE
KR4eUOnISCRJGN9Q1nhX+SHfzeS6rW4u0ZwuKd718xCvohZf3dzb2KhPixSQ0Yqn
FALlt8KZSaPoX+Br6SM7MgvtTON7UJ3yDu8MhE4wQDv4+g0K6PCFJVzmZ6GxK+AA
UMWpNP2ZDx+okoJg2oPr0qE2qsO7wFuOOjZN0pS/1p9h52dALrv+dDShIiIWS50k
LFywfA4jpP41EBihtJ/jYLWKPW//DnpP1LDNgnJMO4Lrjn5HQbE07c54Ho6MzdcS
s9V8yFe/yYFcycZVrIgs3q4uYotA48YOJjwcnkxmOcYDi+Usg0u1uYj53wTpOfui
pkHyzz7SgQGAWwyo5ZTztxncKvP0jm0/YGutUlSD2cFds8zrJeX5dbiOtMMqGQQx
DZ/+7wPPdIwg/kc7HpeMt76eCSxVi85sc1wl/IsuA+DUebv5PBqgoizK5jGzBS9n
0idtTt1fWeoLAMZmFiiyJ1otrTH+7k5nNttAh0knrnitIJzwNjxSk43bvjWBaSuX
7P7NdtTOPr3XVNKL1DS0rDN5lAVFvZHnWHwwH4gnAS1P+ZEXZ+cAUuzuVSRHj6G3
gLwvn9MgP83lWaBqTAwkX3LZAXcmGUq/Z30nSXk6ebSaZoe04nsi1a5si9NY1X8V
VC1F5gG3mJO1yg2XwpFTBJ4E8CzZxjUKnu7bzz5TwZrLj9Rn8c/jOjuDpDjFLf6a
sJtx0yFCCIVwvNlXXUOT3mlakyEKiUJAam4ae4a67d2czEP9ZuPw2YOMGLEeyC9k
NhA/2b9fJAu5LAYdtU5EvxDcmXSaM9zTEiDjodSf3PMwy3qLy7zh/X+HtHU9vw7g
/rfjNsKUeBAUTmzYnnvHIf4tLtj//OrELbKk6BTJ5WqexBCjGpf4zFS0dtG8ivfF
Ex1WIm0MNnCUeoYCgj8Ryr9ivC9PsDYk1k1H1V55AwzYlbQa2ed7BfnofTvgpdFE
b4RsMehsS+nhM2ItzJ8nHADs/Uz6vIdb3QA4MeYrilBaCKuIqj9+VuhN7EzDcfOg
E7OgwTni67DwWECtoMlEHVwvngb+en4i6DMGzyem1FuQhcy+mPbhc6xAvm79HjK6
GWKk6CGqb646VqrGpzAnHmo/t1kK95hjn+c/Ebdt3L+LeQAmIbtBki4LQDK13RHn
xXJva73PKXDUNCfPu7C+dk2ZSSQ21xKgN4H8zTgi44/cE26iZR+N8sxNNgIJaJL+
XS360pwW/TwQaL+8l+ApBMkGVhnfBhLLRzZNK4bDqJOc8NzlhriUElmPC07UHV6Y
SdWCI6sy9zC+VcrORtr4vRlmKzAcK0JaOGV9q71XeyR0Vri+euF7SRb4qQPE76sP
iyORlGRSQlPsCtAHsebQiLItfXfiolWPs8g1BZfbNvYeFr4teOJpRXy4bcKPrqWa
6I2vtjYlFykfRAeusXXLXb9Hxyiz/x9tj7GpkhS5F1wLlJPpPscx2GWMpSvM8KTv
ZUgM53SEjeDZ2FnGouJaiCDtFgj9WOspenfNcO+qEfHbFuBKeA+ZFgpqsVHrSxBj
2QpxpXsTwlizPLFTyE6GsLqBvYiB14oL4RMI9UrOW0QXTx2ABbBHCsPOEScdz8Wz
tSMR4LyiNzA+yNeAWlKOW8GznpGyDZb9u0/EGED5pvSLYFxOj51G7RxgEBlwjEMR
OEHbfliiwB8LX7ffjRiLeu9QVIKYrgqO/bgjm6CXRRw3+8C4JgWX09S+b7qjWiHv
c2b2VY330oiKTkkBhd430aTjWcPWVtaTs2DqqQ5Xn9i5dN1jWFMh4FMoMl8tgVAx
GMeByepL8Q2UrBtC0MrYRaLwQJR1JtxlNUzLnpucgqSl5B9ldxb28Trfb4OSfEtu
rlJ2NOGUpvzFtrbQid8u8OcNsJemG/oalHCsjcuQwlbkr6VAEhbi2GQUSjpoTJnf
qfbl//1K725fhhCWpXN1IyNyMApP3zEmR0qIoSmbxFvS+r/+5gBahVZJ/sC418Iq
d8HkhZOrmA7MbSDD/6hiYuu9ERPpKZvWewROf8M2J5TN9EsbNywWXrdx7tBZVBRg
FRl/Vg4bvEumns3XvB9O3UBoagP1cyz4gxr2vUwRWIzCyQ2AYMCwq0sEvv3aRL8y
QTQawJJ6oFZpe7XBLwo9TZJtRJXD5n3ivShV9MJB1BTHQxpvbO3/9lcBai1MGRnz
hoK3xjbkfZ2DslHdvQbSYpqEHFMzTns2R/q0XegORt5z9GGUIbVNk8OsDxRi1gAG
7iMyX6RgwHCwwsqXQpaJAddqlZ5PyKddrfMMcGmXQKgkNZg64eI8ERfRdLNZs7H4
mEJmHAYb8WsDSykAVU/coU281tIWkv4KDdGn2oAyHYroyy3E8ISTWKL9NHy/e5jT
n2iiF6UrKJJ+AoP1M1pPVbdSo690cd4WHYWsfEwm3Ufo2ANX6ky3p7DDnu+EyVn3
rwtXjYa+ZjihvB6Rc65wM5EhVhfX7BZka9AH0iWI0Whmm9gbb2eeV+o6Zr6DFI/b
igF+Tr7Xr1kG7J5r3Rcvy3Z+jN4tXnlFH4OrtrJ1hrv/C2VxAP38Rg5ASlzcSkqO
Q8+Xu4KTwj3IYT/F3JL5bwaJyszJQ7OJJwU0Kd1AgHYG8txkcpi+4gi7S2KaDUGP
0O7fv6mwGJds+ojU16TGKZ4MsrQgKv6DL7qZwLuWGfynCHSJyUbRvxjvZLdP9e5P
kp7Rj/bSu9NKPdMis4WUE/tTiIvzcVhjN4tTPaO9jkmzhvJCl5MAfoRFO8IY8oHU
pOmqSfoT7EuI/d44NDPKLhJlGXS36uN7X93jIsd8+mukWL45muVZfSuJpgbw/j1z
DA/i05T/hWAxjw5lqUUpX7gi/GRBZcC1JdiIgzdHcCvCgtCPIUzkN8fAYyH2NrOy
JylkoX9EMaaGoitu+PfYlrMgIHOV8M0Fw0oQ4iPaeB0ph/ZXBJyx5Rx9YAwcGOhC
avmqnC2oXtiP+N6BZdhG12+rOpbDDiLaljPLSfjDzjESqaRv8JJncrKHnVZEGEph
TZnTHN3GmuPGG6M7eq01aCDUrT1UD+besK0r5M5dOyGlMhaiTlaZdrXCjDPiOVqv
TcHg/OdiaC+Mgt8bQUxI8vHaAj3JHxj9jKRW9aVMU2a7IJ7ekaFnZHx0N+iF7L3L
qmnEYHdDDC2L5/a1UZSJlNWjQ3CiiIvXCN7SbunKB7S6WWRCcf1JBV9SkeEmm2Qe
nm4jwxgNC0if2QsjAVI8pUI3Irli6Bg683Ghuae1GalGxrwiISN+LEwkd2jvUPbC
D8WLGJCQe34wW1q8pXyCqolLFSyjL2OpVQu260krXSQajRYAStSJRVFPrIZ3tiG4
dXnqrN07gVIjIgVocFnzL0RCuTX6nl6atWb5fN6fUw4vS1WGuO3o8lb62r+/8BvK
FlrvUbFxW2s1qz/si0a3bz2yPLjUFEjYjQwqNLsrKsehmNI1a6wDPtLivE+0GYIQ
OR0+NJFY2H8FZAfDHpZNNwelqPJ6unQzmL+9/6IreycePI/lfvXzo4dm4jPgl/FB
s69fJO3iJKYsTCOp4rMyUv1wrBgYFGQxwvvzlBUIUjw48ku/G1D1/f23tWR9bYwD
z6BxLAjjibVk3nMigZGzzCsHaStxMdfgzjUreWQgpnLXKEVST/AEOe8rCSaoc4Zy
Gem3PQaMyC5fPpoh8SUe94O4sCaLefTblfF32F1LM5Bif0f3HgOBXJcerpd2wDU4
BWD7YYlV9KkGLgiSUx2u0Yj9uSdrFClzAM6MK+Dg2defbpg7//xz0KjY11RrkGZk
khl1S94sHG6hh1vB/gvWVfrdq7YnuggT3y7+e4u9BLj1tnsgGc6RA1OKq4GYRSrO
7F175L6rFIVzs2AFjhinrXyqCG4U8alNExmsdBjKFGi56iQgpN+DqFcHEeMHpU9G
m9f864tolh5eJYp6csOtjMB7yl4aMBQL5nfjPXarr0JHOIf0JeEGECo3T/9tBx8G
zHLaDw3UtvpSncJpUQC2gOGOdm0AQpa2ArWInzHQ6fJcfBrS8zKP6iPwcL1uivkY
E3/CG67YAF01x78bnEVAbVvpnw4hIH6eDcDDrp+m/QN1FkGD8hSsFFH6iCvr7EzP
vIWbrA1FvWrBpwYHKwZMERGbKIqxI9vIpwFOzRflNbiUAA9UesrS7bsXXTFQX6mQ
t9NXB/cTop/7kt4WhBEJU0zBV26mZ/GuHmIv+JfgnEOqxfRfW2oiNSFdeOs+EaVx
gT91txA3iZP4iGvs2vk5eFTxLFs25iR6j8HFBpHdu2yLvB4Kuzi9kkNJPMQG4CzX
OPRSQ2Xuk7FvMRj2EM50+e5Au+XE4hWoaffdSbdwV2Mz2vWeQlbQbujNGOIZ3zrZ
NcjeBJrc0iObhlzX509dMdvPwLVbaywatc4I15bQHMDLx9R7cIscUSspKZssyW2k
OMVJcnKTIwcjuI8tu3Umn4DKXGTieOQ1oGwgVafVGdFrn4s1zfyV5ZjOMSDzKiEc
ORmuoZIHhwhLhcnK4et+hXaFzP4zlmv97AZmTRcd1eSV6IXKSkBwZcsJQ70O2DmN
TMYgqcyCYdAbkQ91pLSxB3lRZSpETcZKY397f9DMIlYhaERGexEKZuQNbjNN2ojt
0YBAJrmaVIA+2VgB33FYS24e9qs6SgIafhDYVOmfmHM3LPRxWUvY1q7zGnQzwh9u
qla25ApaEpElkQ5YP+gCazrOyvLoFZE3LfdAmf29tuGRbisbzXMgyL0W/i2+xyue
Za1J4Aoaq5scu0d0LIw46Km/8Na2pF5lTD5Cvgv9lkF43nr01pY93/G24NdKR6kL
kr0dJCYScmz/rCYgd6gQ87KhI4lK8VdBEkuqZZhn4m1SwRcS2hyJEXb/sclZPJNu
J6mmxg52XCB37P05tWFDPyHdLeH5xBXDxND/v/gw9TxzHsoLJlCDxdL1zbMsGZzZ
gI07gEQvN/KSoTR0lTYSPBp7M9DlYW9Wq/+4O08ZxVSJNzftERi2n3AhAKPVH+2p
ZMvE5JzP2bR164iG2f7RkVKeEeivKfl9Ya48kWmIi671CwNC28FVF+eCqWGGrisz
IKTZcIw1WMMVg8SZ4KF2ST5rLAcKcomRApi/aHcHLZiYYDHVXYvj4k1jx5w0TtsM
F9CLdSZ+4KeF8XZM8M/XGcyxMPZKEJtazXpXcZQ0MBY3GNbVO2Pm1tTEVtqr3IQw
GuZDNsFSafiiUN29nWwfKVN4bGW6Hu2ySwstgB7FpxHZGKYsHTSKyi7SJ+4sVfF9
dH44Dd3f3mmlAJ7BqJbfzNiPAy/CO8UhIsDQNIf47slif2lyc16ehpQaH/qdpAS8
eor8QNVoMsDD3A/n5StWXmFGo/UkAjpX/LnKdQbPgFxTXn8HaYFuxxUy+d9X0/r1
fcew4FbrIo0E0rEGxwSHIffkpCpPqLSZdbUIgQ2cG5Og7yUa/rxhplbC8GKu8Uae
XaEB/qgOTMCohlL/tw/mPwRQj31YvzVscBHs3jlAVr8KGjxDHsnKudyXO5RfRqrL
FvGXKdmdZn2JiMMXoN2C6Do4ePHHYr7lyba7BQfx0rKw+OL5ixuA98VoTInzyKDu
ECGvBypltk5ImAAqHG3A+xWoiE44vxMOUwVny0GNdiRmdq2yxAYqHZFGJCgIj1Hs
EoxsNdAovX8iJU3Wr38xHbVpZkyk06KgeowxlX+WeJlXmC3PUaMLuQSRYTpV9wmM
8dI5c2NQcwFQAuuWqmfkuTDHgG0zZTtTx2RjfyWPb+FFhrKcXY3Hald88qai6D00
ZD5Tsb2nRpITMfg8piGqfoSz8COEQ5nkbtu4i+pUQOn2n8Wb22qkgLC+X7GI11vU
BLgYdsedbpgT2jI96i3Qf33aqxcQBNyFKt6DVLO3zcCIWHQXDraUwLZTl3Cy5XkY
tuAgtEfHSsBSvmLPnk23qctHL3GSEOtklARRSQcgjepDT1iYioV/mJwaAXq8e9Bn
QLe86F9GUS8PN5sTYJY8etnrMduDXjg+A2Pl+6dT/IS3ptyjZVAWValKtb0z683n
iwJ9riPbxM1rtUq+zUAfkpI3Kms7Ib9bm9c378sTw9TSfE1higviEp4wi2EU8hoi
PJQ+JZBDcOq06vYy/mofImbvkRBmNMq61HOx5VqQ6O+m1GoXlY2OhdqY0gh1DcSV
vBB+DGa3bvWStuJLX4UHG37jQu5MYH9mU3mtO5v/tald1ssyG9WgxwNLUWtdW5KY
tdrMZplLu4WPV2GyyLKMM4eTCgMpAD418QW9LrZl0T9k8spLumLY6KpTP5M4K46L
46LeMYwvJY53GEYs/WbvgcWB2SJ2Xpyq0agm4670aKk7nZONOp9FRZylM93UFt70
1DX0HP57q+haXiIXYqVh0GpamB/rq4HfGDDk8JgIE+jOLziUuCfE7YqrmzEidYmA
yLOK8Nm2sq7GIJU8pVmORArNjK++oyWUkvUVt2Aeah6v4JDb3F6II3JXLeC5kqp9
ldqONHyb95pPF6P3dHk/F03YwNm/NXvPEWXR/mfBm3WE75NPuWvDhqallZ9yzHV4
wLNpbzLaeq7+Qy4T7vQdVfuelhD60rfW6bWKfo27ARdnZ+Gw3/y3/e2lDGzPSulG
w+tLLtEW5CVAEfDTZ5NYxNbKOk51OzBoQWB5N6poXiwMcJnz/ZiTNvuijdRhR731
bnN/HBeHcLoExGKxX28pq0N3dW+oY0UyzFVVX4JDrtKDWGyj/zzra0jMtxZN6Mvc
7baX02wa0oGPE+JEOkNwjWFKmeJ9avso21i7IOWNQA1emcmoSYHpoIH6vwEtGRST
PcbCsegf/n39hB9CFxloKYBzwqrilvJ/EVnxTev5i/ugXydoMH6vCZaQc/8vX9Eu
Wyj433SQ+ZdpEaJWPs7VKFnp2QAcfZM/udIRPMdeSoF8ZT8WOZnheRXYBQ0NRLlG
p3NYNPblTp7KRpFNcolTcE3IeIF8JK8SPc0WhVPKSevT2k9BzcjWhVbvaEk2dvXb
gJxQUzPjrxcjkXuKguIY8qCkLOjpDCzDBmkQQUm6H6gWuS/FPZlzWG+wRYcKX4ZA
Ktcn0y18/sbrAjjjSVpRD1pIxpi5/KpR+u9rYiqiaQ6q3tot6wUJC/aPxtb74pCi
ftdd+lt2HZqkDsejs0WlTcJ4uhYJwU+7gHxubYnayLvv8JGUzcvlMp38tbpwLSGQ
f3j47eIHNBUh9Cj4OqS/RzWt4WbCO4ISYHSJd2wz8yBqLdNsfwSiRwGc4Vxw5oOY
EthheOhEOG8MMZQcdKPQ3eRQqZQ50m/EB9sbxCUTjhr4YBmY2jCI00o727SP4Cvo
nu3U4N81oXQY73CANMyy+N800fCzJtPiUZs03Vxn1wEKx+bbCbBdA10spvi3jsEZ
M9YNYq3bEiIx0hNBYaPT3B3ptDqvOU2XhUoFh2IAYhiLy1a2p+0EHxClfaYJF+UB
hRaB09Uj0BNQXx9mM9dBxnu9PDHBCdXTizEJuPLs+Sx3HDBjOqdwTGUb9+h6K6o3
OktydGmug3HIHLWcSXHwY6nH3q487mh9QZ/CNFvshep1ffe4ItjaZZiuFdHbB49S
qED+9a43Oow2Pjc3+gHTj2/8hu4hJlpVAOEbDctNISFIpZjLqNXYfvVYi5ljqIuD
3oNohpcmiy+bSgq1dFpuQc8ApphqmZt3pb+/5W3LEe+6xk6xVzm4uMArSb/CTCiF
+Q2nkCvD8ZPp1tfKKJbVeof/VG0uFS714yWRTkLg8lSdzltoMGNaDt6rPsRgpmG/
Yhpx/D8RfOdBjxBG/axe3ExUBwU+1bbX4k6zP1l09Uxq3+/KqhqPOgjjumxGII7o
obg+cPaCku1jqg1deTXzOZLX8hG/vJHVLqPa8/nN7EmCgIx+Qt/FM2AWkFZjxMNq
4BgNh7uBGDy3Ts8ZzGqq5kiiKpNRVOCmkqXjBTIG1UZ9qcotMMpTwrFSnJ6+qEl3
vbOU3QKLCyX+gkzJRXE6qhQQlasWRJ8OPud6EQJ+WME9lsT9YznKpc+seD0wqHGn
3lrTd84T7Ch7hE5oPTNO/f5lOFR52QL/g4M4L3WZSMlDLgDZcrBaOxF9TDhAVwcH
0tcD/t+/Ju9dOgsHvJ6WlJLGo1po71AK7HSvWPgcsEkTi0Na5eKZRBB0RpCCYzLn
wsRlykDCdnlLQZMDc6XT0Q4ctWwyPzbaGolzd2iO07z25SnL2TQ0vHuN2K/bitAN
CEhgB8inhITulOAoRFwJfnF9T9iTSlE2ktzoc215OdLmT5eflE3HmQFpHTjz9x5U
aW0l7COpbVdEd9Pmpp2sDc0QFizAn2BdSJvf/02l7fRWurxnqqUL6ZCv72pPjdhf
HnvxfLsON4R5eTipNHRdre8ijnEZCDPkZ4U19gkn0MgstQkKvF0X+XMvgvngCwbb
zeDrsbod4HdaUr8obJH6wt9/WwS8XtYhom5UdQS48je27X52TsEXoaNQLRuc2p/k
9gfraLsmPbz9f4X1ET1fvUVkgxS9r9fgS3i6jxWkLi1cUQJ25ty86aVPVZ738Z5k
CiKtNyfKpnPBs5DAEL0gyTGzNauK9UH8bHbmB+c6Mcom+xlAaw94MBom/Ip07/Ns
IRg2umnjzipFipUf1LHOrLrV6rVBaHgsqlERTJ4GnWWQJdhFEFsgmfT00GCpEund
XNzxlNhSQ4G0Xy3DHO5Z4I6Gcn5MYng2ujh7d8K48g4UnrM/zBYYizS0Ro3MvZMd
ybfYylwHHYOBNVYmjVIlfoYhtmNbf8Z6JrrwqTzrKSmM3F1oil/1iaIAPaPmAtWE
7niQO3KrxNKraPpboCATAUBBHJzuBr1Td9pzSjG1ZVQiXTxNx6cDJrJ2k+EhHaSg
x8jxpX/75hR7qOIcoBp4iTB4RFjT3KHJFEAkzCwcLYOgL6rhQtNy0gPRbESRNV24
EmBkHhfMU4uvrmjdnJCuTatZERdA3xmoKDqWPQnyEmVxMAX7+DN8VD4PShmIazW0
QzWxOfiFBw0MQEtURw3sZFfKTsmg0YKElZOTVSkuPIE6JJM3TizqSo5xYFD5jqYH
yr1tvZu408kX0UmVXGZTh/UF9RkgrjscxNX1a99+PWQuxlhNt6CKeEzaV4y/ckdU
OIEt+yoUyDFkb0Cb/A1MM2M2OXbyaJV8WhcVXLHV0O9BNB2xq4qfr0IwaekppbrJ
vlVn23YJpkmP7DU4EAGv8njdphoeb2q72I7aY+Dhx8PRsL6gBORzQiVzYoNuMSky
F4J11dizn099XqvLF/thlRUpY251BWXxUp7DA6kOkejzPNVsPhYhq61OVoTysexQ
gMCMjibvX4FFuGgcDK21UcaO9AxYUZ900F2By8XbQuf1R6TbsP3pTSEP6MZtD3u1
mrQIJTfBo7uSDajujSZUGvj7i0scZm/Bb4hXI/6L3qZsoFYzRhxy7h6Hyqo8SSTu
G/V3s//0FZwo8c6GYyF/0Pd75OKGf4qPSAcO6+lVM3Iv66dZiq4se+gusOTjby5H
LAmSqoYPd+dhKMj2MgPh1iqhHDk0bg+b6MjWdvfi8CeTtMfGUD5VL6GvKWtKDvZp
XGsxhVoHQI01uYeNyH6N/hGe1UPvaKbsvmJDc3dOKWAL+yoWBtc38B8cNJm6p+jo
iH7ACE1N4W6j1+osKTmLT5szXNd2KkP9OG3e/LUtjZ7E3dOrQiy+7wQt59+jaUd/
j85RyOk6b7S4IbVGgmM1VvWreRBohowCKo5t3a6vgz1FbIMbZsRESOQ8CNh+pvk5
VcgIrf+Lu1UBNQTd+kEfnZq/JZ9OjZvl5N6abgyI7akt9X0EvnVv2xy3BBOts8gg
om3ll74yDKvZTrREHRWziggTI/dBEDEYb3jqtKIrsr7uCeJYn9uGGgF59d1XjI/Z
vkfiYf0btO2T8UwUVF82HTZWljaXTSttUdo5o3vQnqIgXsb15H+UjUe1PsUFyRtX
YFqCc8hmStKoJy/838Uh4nXVq5iOQYYeLqU/mz00EFDs2fKHzIv1zkWvyEm+Ebd4
z3ucCfoc0Q8+pTRAc6XgWILSqcNTR0WCm52sdFMIhDjyd4GOtl2hQgj7hmR0TU/K
w1S0nvlPf4w86di2A53rlmN4X/EskllPG8f4EmLW7YZLZPG9yqLT+Sj/aSi3DKOO
DgEyf/VEIrulSmhCSjxx+EmBRy7kE0MH6tifLk5Ne7FBAk8XFBEHjbOsmSdMvI/v
NncgpnsqNYv5tjpwZ/Ux1p4mmULJIGE1DiofzsfgKtEVgfZWRwO8k5rTLLn6MXbU
SWDOi0kLIqKBbxuNq+O5cjNwNV87rmy/y5PkULB1LQDo8NsTOpfufzV/CcILx0s5
VWS5sIgoXrXkEAdkJ0JE/SkmzBXpCrxv2Fg9wujgqxg/wsnMfWoi/RneMBYtWnuH
Ti3a8T2PgrMlkN6w0nsbwoXyMDR0hg9Pxfhd+VAR72ZnFJeRABkLtGfYTyxtuoEA
BThP9QeW6K1FXDSQrKs9+yMkTZv7bdWwp5vPk1PGLgaZ4KVoYZAliKHICKM2I79+
PgvviX87n4j+axlwUpDVwfTXGejwsYXIXt2er7xC/vVm1whfB2S6IHo+XYOZAgR5
SuW58ZDmB6vKC0gfYWsziPa4GyoZ5w5NvDDPJ2u0EpIDNZxYMuZbIQqA7QBsIhOk
HB+5Iu9o1/iOnq35xT+lg2etwHkayRjlFWZqiOTqq2JnP7sMjk8Y0ijqKJSBKUmO
a7I6dU+Pr0fk3Q30+iUdLNtZEPjRM3KYLdjueDticsyYykKZfOF5MW289ArjAMXX
/a4QxeYAJI7NwFm0Ur+tKgvRAoItUs0ga9iZnqNBOXK0kI/AKGAYzTNBg5BGxlIT
dJvOpJx0NHaK8KqFGhLwDOJQ5ErwhHRZdaA1AxBYedDDyqrI4fK9Gvt99U3CaBTR
xli1yJZrF9CJXpZhaVol/5euymRl1ZcUPTfdSYG+gWMobHOzZLe1psEw7v3JLDLz
tUxpDeqNgzvhLXH/kzATZsij/laPRUKOeDo5APrh6AxiOzJBVTDwUcTkChtsfIuO
UNEOOMtiYKFUkQzTc9jhHbqQydUhP1J3EG9so0LYd/6lcIToUQjRL5/UIr/OqWIC
qidYXZcvvc6WJJ2timh8anMgwXPke0EoNsMSC3yorNkGcv8l8kxUaAKxarmR6awW
taNqBsO0FvL01Z0oGaxCRJUeCxcOC4SlECYhx3FCm4QDqnKAWK+DLVAbfmd9foBe
WNhZZh0ErBRlGBiGHI2+zNsCPAnl4LRAwa02Gklrji8CTlenM7cZDXRaVqVhjkAR
JH7Q/JQ4OCHzN/iSkkceuf5MuN5QOTcENpqjPyd5bfBi7tRs1IjEpYkt8yBsj9I7
EU5pUudFUfwm8Fia9XK1Kjmyu24iAIc3nahN+AmHa9Xgf6Ba9w1LuizPjrBBRF91
CWTDp7yCaKtBDYpzVWnhyAWbMx0ljA3fy17mW9hOW6K45F+JmhpfeWzdKvAEu2Cn
EV+N3gzkMvozo9tZfWD+gFrEa/6IpGdJGfieQ0AHFB+oXK7g66/ESMk8Rzbdu8If
eVVlV+9fkO3JEiXH1+RnF5E6B+EtOzYqFzwiCZfdeUDwaT96neVX+Rbpk5fHRYFd
YSavMMua8whTNPNZMD8MImo8Kp5kOfsL02u+UKG/IvGHEv7soa1SlXI3epLVgOpz
3vS2LRcfELvJyHyx4VI9UoyRbAI2Domes1NjCYO5pRXldFH1D2wEFOZlf3AX3Tzr
vFvNd0Ka0mBlM5L4c6axij8iw21c0KMKF6WIRbcIPc16t21eH3GofbVX2/oUxIK9
byyz3eOjmoXApbUKBD01CaV5aoHbWB0JgjTN5wWJTO9UDqP45JgMl52bH+AgKb5D
iNyPb4+eSNaoTqFhEbEU514ZKuy4gaOexGq+TqIMp+EUBvza4FpN1+u1Kt0YXb8i
4ge9RAHEKluko4l+f/tVI+hgj8cNqkvuGNVulNlPAIJzXupOItDxoEgDOvVTUGke
ceekG8f9Y/bTSRoWxDcPw6O6MTcJ4ahRfvE+cRWFliPtcM6Fcl5nawEsFd6B8jHp
ZC1LY729MpCQWthTpwAfju4GdQqkWDprOLWfMI9iZ4V6IWWnLG8g2Et92I8gF5Q8
wZytL63hbv6EY+BLf8hmtwjspwiVKzqx2PHeTqPRpsedXd/3qamg6C8SVM0dRdPH
zTjOcFToNNiAi180Z7HBrtGrA+JqiL0KlrNh/+gol8noNChFTKSVqtZtdljg32cX
rwl1j2up2kQLVU8SxmGMNlz1MDmP7uWCIxuJoUR3t7YOoZNHkPXsjWeVduzGMlHf
s/9ZSjvQjXPEqWOQucGkpX/hVEaAaDytbYOnNlhgO/d91E+FJlVafrD/6i4bE1Uk
o90HwuxcFFcLc0PVY66VeNr58a47XUFFmTXkFKMmTKBYd5c8oG9f940PVmfQHZ3E
pWFhWr9C4bIlEQUPv+13SPMi/xW7/wrFS8w4A5FzuPUZC7FdnwuYIcKs/VuDrzvV
8d3l8TExHQLKpYLQ0yoAvSCBlHDgsIwIrALubRcwEjnHSOqlnaV1cX0P+cptWp6O
uaiaTGnzoaozx1MSdf/P7rdUYoFf4V+6RtLpRf8dAKdSJfMzDBQd1LIXxhnJKvjX
Ff7Py2K7JyxAVm9v5OUzzVzRe1pHIbezlDMylc7tn5V28JTGND+8GdhGUeAr2wSZ
fcc6X9kEy9s27/S2i6ZH7A6T1ThPs5X0yppqdwCZEq7zLyiyxOtOkdqX8IFFcIp2
JemunP1WrhN1nRcR7tSdks4dCLbFZBcU+OigthnIaPKLQlSNHjAJHx/CmNDPvEEV
EaDVijwmA2D0ZWBSReqPSlRXHh61biPACJo7Lc/YbaAWdLMRwBGc7jjFn2+Bj2bs
fVNVagtko5u+BoVWwkFAKL3A1M0eo77UwEsdKWEvNFDEymtbNSLyUHJCRWYnzTxN
AG0Zok+van7R479OcwyvTBZG/yx2TxLKrApQb6BqoFoSO7GeinG7UQ3disfH0jF8
qx3N7Zwfkwl8UtxRQkC69i3J2xWmyzjEoN2Iq77+vF2yU2GkL1c1FyLIDCkNKg//
z2SpNzwAoeF0D/Iv1ekK2q9FlizMS6/zOGCfIQeh9t1DwIQ89K/5gBRgc/ECZKDM
Eeo+OWiLifULCeu3L5VVUtSx86cwCMjqsVMOo8F3ux55XUheigeUg3rlcBeLM8KI
cIdz/qz7p3zoI+I9Hp3VHnGiizYpJOTcAARVd6Ctza9qUnZvW80AAtGcPFSIKRAZ
KQVtQ+OGHCkwsAEwiwfDT94mho2vwMvoT4lMNBcuFToTIFXE3Esn9N4taQFWXbTU
b09UOgHhvOUHe3/CVpGmQyUBPfAGar1T7XWSQRR7iFWzaJxu3CosaP4q3WY+0igD
2NA9P1JcwK6MooJ3ezJ7uNRRcC/uv2XbVUvyPMnShm0BBx34hKOawyjSkyhPUVIJ
GtWnK8IrTA9fTghF3zqtQos3i7W8KXUVp83p62S94cZWn0pRdOk33mbr0sdgPYKw
0+wb1poKfxRRsPRquNwdf5gkAChMgFLTb0pq2WJTDPJs2XS+lims4jl0Rmr/venL
dKOJkRa+IwtGklZ/790zq/GvSSuMLiF5JY6+hUqpPxYlE15mcvArwhiH03NiN/+O
Pq11YLPZDD67lKi0LYb8qucPG/fLwcT2VG0H6kd5X23X3i9NWKa74+cvYs88hrbm
SI3R7DH7CMk0ak/JioaSzxpkcXtYL8cTFhHwau/dhbkkng48S2uaE+gBEOl1ZeBm
UTwp9kAaxbcSwkjQ4PhbW2/Z794DR+8WvBI4Ga/OT17LDbuo2FOLNQP70CsG8jsR
WShsGzOLACiYZEdd3+VT92iDpOV1V7n3a1QB3Vw/hHy/WqgrXDFV/CLOnOOm2zOt
HK6iQqkAMg83nQWUAoWy6p/ozXz+axCWTjUXYncsBb1Xlp7wl/6EIAFOD5fd0g0p
FrI1i0iD2ZQwO/Scw3kCvBZu4ZWyz36JmELa9RfCacUaS/gKcmQMw3eUyP1hFBSM
+w95TcNlXL3ZcwGVcSVDmnveiTH2FXftKMTk+MFG/cIHy50FsMBS9DSmBCE7F1H+
vmio0vY9ntF7reCjzBDXJEzSms39PLdfkD1z1fWCHT0ifrLZyHZDt/rwSmg/E1gZ
R6kgZKI7hp0sT9t8Ae/74BITyN+aRfehHTVNi2ViZqghprSfSSTVVa9EPL6edUKD
hh2/b5DKkEYHEsAQKzNyvai5zYjeJG+553ADmpuHGEj8acsiM7JkTDGzFj9La3aE
8YlHq1EGbGOJGBVG61MQZQcW7GE5lqAleCQQobBOWWocb7v/+U5d4sj/9ygLmDTX
zFMcR4Vd3Vz5n+t3OgNsxkdUzemGJSZm/z46NtZTaSDKRGnI7Cr/kSOJndau0Yae
7lLH5LF2GJYKrt/0haW7L4HXRYvFRH0nptjuhSIPomasHYs/CuSx2Ew7R2ZwGCzW
vZOo+UH+dzvaYFub09O+lZlR3V+tT3a+GKUB1W0nxMNHy/9V+m4X+1Kp4mn3bPkG
teT8ENReExIe8kcH985flztBKqzjaY6gwwI/0qOVIaTTMjJznr02/3ooNfJ2XeDi
fPTjunnpP5HLCq/4E/6IgiGFl80HhZLWE9m8BQU43AcETpVeTS15vjG0vcUXLt0D
NJ7qjj9/3AqXuvHXqNLKFOOBdTvJmN7cPOhO/WvfD55gLfd18fOZC/llyyitCOgj
MCxXtrNbZApf41FWPxY3fN9q3B7Mfz3k+3pQ4OiBonmDGfj8u5pJYByKdO2HKtdG
JwDzNNq79euX89sr0A+DlI6qiZbypZ5tlKC4/mldMVA0WmI8qTg8xGAS8deOzoyY
xbdxJmQGDgX0T12mCjPOQPVzx4O3I+F0ffCmjARvAAWhzv7KxHi+lXVe7PoxfmmT
WD9LnZPfP1J8AxtzRjSkb0rqYEOC3M0TzYV02eS5D2nbNcsTjx4VWCJ/ShxC1Ym1
L7cokk7kmKRLv3fAUCiy0bk5vkozPi2U+Yc9eYL0ALIBbUy0IPgOy0KWWgHlPfw+
cHHFRd87Mzfdyf6FbyexfRkzX5hhH1EEkUUm8S2+E1UMG+TrXL0L62NVyrYMcZGO
W6UDzsM6m1AxMpKXtpCKMA9hEiuUYihK5yNw6bCbdFPvlEjj7dnlLPetbCGYlm47
O4JNPBNGyU8rOTnX4VuQN88YUQLb2e8szw2PoV834TgXaVPcQ7v2c9YK/bXgPitJ
70NXSfgg2DQ/lx66gzhiGPUDuk2mpTaQjklXHpzJUj7Y4xFmzhQMARKeXiHAqnmW
DKVBjD87D2fZwQFx9quJeoebaNDwSFqsYX+CRDmqbtHSGoWeiQiwEmLVVHRjc5Oz
wreqsQdWtWJd9/QYzR1LRdWzTPYyuxhFUfsSNUgWqvQ6jnxPoSFjWAs9rWvMJuaB
YJM+OL9Hnv0+x2M10ew+dtWoNSeVVKwNr2Jt45KPotzcLm6vJFv4MPhraOi2y6tD
Ff+d/8M1dbJL3zPIE4NFMxnoY3dKeHP/Zfx5/8H0XQTr/RBBnoQC9iYEN8iwbI1v
QDbam+495mHdPzr71Fbm8W43z60/rMSu/yob1paJWMabQX9MlgoP4TzhmnEguaxF
zxVGyJa7BwaTyYHquQSyGgg2AmbRfqAKCXN5T0VxR/H9o8jM/6upMQ0Cv0lpbQiP
gYS8FkS4zP/jotfV0VT+iNwae/D0xNjwB1O9Vz71om0w4MZmyb57EHZ7a08+68mU
ATp7tu5EPTCExea6xN5L19eOZajLV/1w01yLh5YvqdP2XED7P3b1dtKcsjx8IvbV
hb/BhRwOtfDxAHeSaVedqnghsKDqTaXa0lh3L2o9sYoj3e+qlTOS9jCx3FmErKNc
aSDfq24o/CoexSelWcph9JcN4Uqy2eVaFhpT2/4dc/lGwkFtPrVOVrHcm0x3+9XK
VFBg95QGs2i5qYVYKE3BlCNzBNddKzXhXraUD/qvxAawiCi0ZNnzYVCvLLaC52Tb
rGkTz3BhUvSl8j8emzMMdLmbTyXXdlgnlexBxEyNEJHx2wAE9yTxjfah2jArMv5X
jkncyGC7bxSA/ahoR/ZFHji1cfRBy1wwlmlp/ueHFD3snen1adkWXzsYO61Fvxiq
EKWuYlETHRQfP3jU9gzSBX4CyShyCQQR2PNq31+4jAlYHtuVYJ4ENaa9Ewv41J5J
skz25E5HjB81rIchOUjHRwvaDUtFQlafGywafgHMLPDZAadT1VQgsfVgFlYmjeqp
50DdL9xdlgkETAj/7oIv451KV5TKPeXuK/1xlOcrV9R8eMd7eX05jZlmf6ilLZ28
rQWkWtYvWVd4GkwNcf9eTaH28XGIHRNt8xH2OPnACT+nLhjkJgphXWMvXDz7WEc+
t7eiEtv2I4mVy9xJGnLDKjT7cCIuzDpP1Um+GvmxueLI1OC1+ZzgveR+cRcUbE0b
mNX6kOItgug924kwiBududBeeEkOw1lS6gSqzX4T1stOr1RB3ASk7KdE1HPN3SXj
gL9B9dNRicS4gccQhZsjoFwxe2lAlMmnX92oq2nE4kAYfATQl3++gfkLr6lGIxlh
OX4ATJ98Saly9ywXX5gV6xN9QF9qbtNf9mKNBB/ye/306oXufnvQL1f9UrD1czvf
xY1+GUYTiLfBrZHv0tLdJYY2afQ2p57muSkYj8U8Gnl3KHT0t6pqjzS7E3VMbTjJ
L21Zj43FGh0CqpTy7Mho8Y2YQdIDr8dfe4daCHTfc0rF2INi2OXh99xX75oiBlUJ
p2H8OLhPh5ezW1cpdL9TsNPSF+OaRBzNK6Z7CQQ7gYSYduvOmircIXzjeHdrjazC
jseKXmhAIpL4Ul0d8GyQ11Ffeygc4O5jBmX6zwJqqGs6ZwZjiF7KCey6cp891+oE
DtpsPWGY08Cf8wWO6ONgFW4qUxE/wv3MGbQOTcrWXzbefCyI5B4qNvgfFyjQAqLT
rNU/UGO9tGpB70S4DQIXMiQtRZ/HUfUPyu6Qpwsrh7WEcxDuXTV+tITJ7BNbTY/n
5McUgMjaCrGNj8CzzJMYeKJXLU+xcJfhzR0EHoOz9l9ralSbzbMF7Upo6C+WG5YY
ZO0aD7WFY+pd0179yt0QX00+bUSrbdVvG88TgN+edGY4AABqITpwJn4gJMaoSTmv
U/c67Th/eoEgtvomqM6hijIoojOHSTucqsdhkAfHisK8JFcOpBDwO5umUXns0zVs
POT/UTEGR4dfPerjUqrwYSAER+OSITCXZ39S5t1OFRZIA72rTxHSdW9fOc9lvVPQ
xyV2aAXpVVWxMHU6bmKO80JDawGex8oF7A/ICMw1uSSLf//qVTqjkChjKIWzQWxc
1KEAFjSNtrjCNxu7X729Vb0YYDdq2+3bpMLZ5qp+s49uKTrRqt3h88Oek4dnuMyV
/eP7SAzuB1o2DfXdy2KxT8+5PitPZpZkA8fbTKYRMn308qcyc5A1l9WiSFToaspS
DoXy3k/4TzjDOb6IVb51yKjoUaauXoqpyGkpS83dyuEMCtqyPPnfiZ9Hh7SUtOy7
6gxJt3/olojzZNxbbw4/r8Rxly5qx83ajtHlR1HvdIQNasI8D6LJQMfNhQ+roeYl
s3N8+enQPpW2U85aCNnGZltQcUkxUaX3XKJ4Yu8JZsViFNoOrlvCum4oDmO/hZ+R
Er5rh+ecfaWgGy0sz7fzJTFEEBjFqLk0lsuHt8p+/4Nd9es7KmD3zn9DBxk4cjzM
09pU/2pYhWCOftfFwMso5HeqmkhfX7GrMqlhJH3x3iyrzBY1bPm6lb2F1IC/Xqln
ubZtON1fWEMiTxHrGixKGUNWul0x1YeoBqKP1m+Pr0f65eBSf0xHQh56/IndZ+C2
SGo27M45rg2SJTsFWSFRQptzWQ8dM2p9680wtyCUK+d/XUV4Ke9N/E48YfXlrTQ+
85Z7JMfInUtJktKzTskME2k0zjzodCsd4ClwWT+kExGbT1yXtTO6D60GnrUv1jU+
9wUa7DC9TuKlPP0T81q9y2tZFUSd2xElXau3zUFIDgHsJUdoV6Hi9P9bptHBeBoU
yZ8hEDOKpwHobw3UjvfS2Nx56mMZkd5OyyaarUDoKkAFxx+ZhKyoz6l3fAXTTBqc
W/F3cf+SxI1AoxgSWooORBD0DuyE+0YmtxqXQi82NMLV46CHTDJCLoSHwf7fByCX
74+wxNIn7bRfwUcP2FZI0oIzqnpgFxuNNZyTqO3ohOhWZduoz7B7SGE+ORwcIJBO
YeomWClsbcIqtOWzndnfXSNNhIo6gxYlljzh8udt+TfHhZEfCumB5Q9jjjnCi0jh
OQmvMjqWoqBw1/+UEyuKeqMMcTRsUst//HloPFqdYpqSODvPcKUxb1+JRQkWebUU
IXu0tXKAzAOywWXvoe6W1pvm+WvcoqIormf+6OijeZ9tskDGx1aqc1PZ1im9hqWc
8jhM3DwTbSsMP9C44p68i/YUfN5tXOU5i5r9gN772obUMqRznFAjpc3dGWpEoNly
Lb6IUw8NnhgS2cn+JHkyyEnqdqseKFxNL7MOCQ6fXdAn3Lpr98CrT47mrLWagaLa
7HkFS17KGVF2dwFGdPiB3uuCGXJ8SKKlVoPrbNi141rWZET4VhbLRXlJ1zAFPycj
hWhCjBH3sGIVaTy+7efC+RwOuqY6qTtXWpBP4sVk9GNj/pNjDPESlykwfwKGw+rX
20mxpvM3HeUIXqK47NroZTQjo5/AloZH3Pok1SJrkOf8yWS/4aZNhwVyYhOY5KcF
rOnz/iEKGZoj2+WiV3Ai42J/ILRyp7YZjl6yPbz3/mzrrtKnFouZ1zuZQ/9CwjoR
8aOy2RuKbzOmtMkPjse1izegM8+VmRIC4cr7AntxqbLWLUL/q8VbRsOGqP1J4Bpc
QKHJOI7QP9Y0TF1SOmqM1s7ytJeoVzeYD66lwX3E1zY+YYHGsVUwGkihYwipUcd4
8YIBFLKE6JedKwcHv6WaXwg0irCp+kHc0YL9WCk5N5Ltf3GV5o2pTDIZQ9zvG0XR
PEWMB7dGE4XGSpUMXUVi4DLOzt5SY0ZziMiLxV0SyF6OVBPHpz6B3PYylZcgbfmN
SFZ+W3c0e/t4T/I+DdPIZ23Oy2+bTx1vwvujAJaDu5iQsZOTlTPoYzDymZ0afv+o
C/H8H0c/NmAfZ3t1/zwFWxZD3us0Xsgx4uTJatBUuX/+5EU4yLdtUi0sOsbgKIBq
pr0nRSBXH2yjmXjmQ/YzpnuCp7iVoVI5NdmmftiCN+BrPIKegy/Shq4ciitu1X5J
reQxhfevB08ZpjKPXDdABNnsLeFRMdRNyiBvf49e/zCaDl9aFtmqATf45YBNFHNo
Mfkh+7a/aOC3xcGIWrvQ4jaRSKhgfJEMstammJKAt53nRf59jvmHWohvJcHOn175
y7d8pdPj93c9Q7uYYJp8kcMzYtO4Y+AUdemX4ENF58rO2lzI5REuMuxl/ydpAVxp
nBSr+tbm0bsq4c9MyNcy+ySyjby+GsXxoEsvdyELOfGOOyJEuLgCCzNfef65A4M+
VOXD+eBcui+66R9DiyZoI4N0yk9lV4wZVBFafIgfPM0tGA5Ni45LzmHKrVDqCQLj
Shqjr5S4vzurc+1s9qbWSnZ33LgvKNCTj5SgUtAxp3QY9eb/NzLKTH+irSPrDeE8
sAVpaQxS9WFOESIEu48NlXfV6ZrJDHsov5JkYbWL97yFhwbTNu/5KfOHuP4yyfXC
qE1jzeAN4Ssp+ROdymJys3CH7pZCAT6TlhwZ2XlHkhHAFHqYDJMjx1Ism6y1ijC8
OYuGFxEw24Dla84OmC9Z/2m/QZQ4PXRSfwYb/SSbe+nokCAOdqp8bydh7vYJqatA
e1nTBGie6SNXc7wT9U89/q/h7ZiZBt+1HvJnnILqz618lHq+kGJ6xC9wA9G7jYW4
Xo1yLUwJ45+16i27ZR5r30WrynUe16jcH8VVrcDQLqfpxZK1NiYSHOO2BWbnWnhT
vJH1GmI9VL6njfyuHz6pss6YAjm5aV9P+xWOZ41iwFwToWtGGKGr32hK+HdEX567
elaso5kB3uEg2MSDotT9yg6ou3ozFJzcnOsxoiSdq7HyDEc6kWPEZGaPzVlvhxof
JnZe3diQY6qBtMcU79h8eGx17XQ29qc8M+Tqy8P4SlAydKqlg3c+3Fsj2unx2Iux
BhWtw5Yif1wH9UypWZb8dsq2iCHQwzMZKTXxoR1UDhMDWyly1R29mfR/FcK9C6dZ
6NkFeUjDRf5uqNYdm9NTEC4mVECciec0w6QCGXKUVU2jL3w8RarNAuqqTDQQuaZj
n96ejlKH/zxUkbTz4ezqSw3ICAVRSYTMjxnSuMdm3/4SPvnHVVOQyhNouDUbDnyp
9x6dEpDRGodQysqH75ak+wGf2/UxTelx1NmqF7ZxYaOkQ1zNCANAbXOuY7m4Ffpd
jZC6a4L3KU5FidpAVm8zr4lA4JsFKVNFiI48vT5V/TicscqM6sf3qRtwUMZGZX2w
641/l8C3Y76WrTmCScvcK36TORF7XlJfSRiq5ngIf2rfnsbVYkwdhuiknn8oLpvE
7oJ+csZrGyb4hEZjuasAp4Hz8piaLRJnFwLGhQ0/HapLXGCdrf3uGTBQwVkrv9ky
Qynd0aVkxyL0asmmne7RtBQdvSKBYHp3QRu4Cb+kt+EHi/RGdNH/09QCt9MTZYxX
C8Eos2UPoj/5yI13+ZMBiwxXnghTaQHkd+mmwx7sIBDQvvWM4gS7AsSgHMTJmGuV
cvNgRbJsCur82svaUeZ8k4GKGt2fsOZAX83Zki6ukkI3AICKVOqj7TOEGLesNCMd
uz1t1dcB+fdcO88fBulSRNvgno2wa0Eqb+VWwviF1mXEiTV3kAQlbhYlzQ1Ekcwu
37jpXkYvuNo6iFGnMZ22zKF5okRBCXyh78y4ILLwfF932WptLthsN7ryvn0BnbVB
UtaedV0LRnNQDHdgyksuwaNWPvZZB4yNq+lraR/PunipxGinoVKGSY2432GPD7VH
etZVEVkNy6SmvhJL1ZDYP/XEyx/GhaloafbNZrazZq87REhQu7KxDbOt43m0o8dh
+/jBIRWJixAZy9/s5F+wVsY8n+NDjiRdaJbeCV//gkepCLeStBpjCG0BJj47mljV
x2RKAEzgMl+3jdHDOxuGKT/gZ/O9qB/rzT1pMs1sJk+S6YsGDsvjgOdTqzJMReiY
PhPwkQ7TBBHYV53mrsoIuK0/xorJcknh1XNJ7XSoolwSo9NUw4NeZhR9Kh2WvAQK
zmPZfQ74AM/7q6W9imTno/0ts6tLL/aOZsd0pkde7yjbZggoc7AIbg3+xksIJQPV
zqalv0/9LuJ9LQjQHJKqMV2bzrk4FrgKrPbgTPJUzz49upSNNLmDeOUdfokQHx1a
ufWh7YqVi1FnhW5dYvDZbAOy/ah7fcQdAMROhtU/lToPkBYT2AVgab//eWJknecS
e3jDquoXgrlLUIQ6f8/NPOqUg3KaHNMQ4YHeF+lVjITrriicJ2SkbJFhR4FOiL34
MJLNAGuMZ3WHzmRoCmdbfXh+U0FE4y6IUpbK/LSwUTR5EXoipdrTSPqWNjRG9AGy
0hwVY/O7za3hnTfAljDYocTOIIZkUFXHpady7niCoa1dEtMjcB4Y1I4xVdmEcugC
0arljAUESsiOSGo2P/lVdwwxCM5IMkTj2AqObY68RHymKwwcB1jnnPCEiYSuoaV3
UTmXc0IAm1JVpTRka2bD/9mC5uKOP6KIWd7wWmpXEW7unWe5EnAOKFDw82kVCtPU
IkjyzBNyvz0g9COwixyLzbvhEKXzIxwnALL4nvCU3fN7HeCy+bwMh7IQsXrAki+o
aYQYXGkCB9iiyEHz8FWqqwKN9DShsYxkGevpH+Kch9BtdpYCJT0fA1r8uwqjwBDk
jsOEDiNYlFut7Ees6chGhKldlsFd1KZcXdR77GhK/rdOiKY33zyfMrsp3PLYwmBY
E+TU3VjT+24i5HszQYNgvyuJUJWI4C95hH0ockDe3tqprzyyCS0wrrjMNH6C6kBT
LbvGbs36nkCJ7vBcRitw0imf/buU8k11NZfqmoLmPtzLLmzdsXFDuqK3DnSbHGzY
MExSfHeIjMYg6BBmetuF9PO0YIxJe7zKAcNluUYlrUIYSRt8v/1ZzxEp46O5ciKQ
DC127yR+0iYONAp2oMXYVFj5tUMLzZxbNjQnNIw0Mp8taXaiR9dvfr2wai0HmW/m
mISSltw+dmG7hdGfSZq2m+i18ruQbHlqZWUa1k1rR4Twp+Dkc/E5fA/SJT+bzAqs
2LHo6Qfyh+/aDs9syhUGXuaAdVEEwTDiN6BiRq1O+aqES5rip7A6iuaIM8Vryc6H
2I4HU0Fd8/Lq4NaG+ebqzxRkMQ2Ffg79bOQ4yz7G9OCOF9NZXpbU8OJYr37e8xvB
FkoKSBScDPsUxFAh/uDOmsIafBk1WLyGnjRZF3FU4lerApIpJbWKLY7/E6u1vsz/
K7zx5JrrqsAwkHx/jcoSCqC4puw0vPaPbzh+NnTkhShV4gutm6LygjKyfRpAnqys
RyQHcFGG/rsBDpJmMDInQFp5tYeCNwMMNmkiEOqxnUwiYE6zIQZxj9JJBFZ1FSbB
eFmHrMdsxYMOI0DIdwywHJ54FOu96AP+SQKS2IyZWV3ElytlLoKP6bFEyGFhQakX
jlLHBekeUL4xjSUsV8MRmSgregnSYCHEoniXJY7L7d2TQ8mjza+wQSNP4+eMCS7k
QFS6G/wvWJNPeFY7Ym1UNbZxJMXbibHKKjfaUlnhYMgY7aZ+HKJ7QEzDjtpgxHq8
Vu3wFSE+Rv5cwz52vvnAqCbC0xdj3p+zPMj/Xq0N6M0Z3UgAHubidBTABWFl6uRJ
ItR428piqDuBlBLVfoHX1auhZ1ESAOmFZiWzBBHbO2cDc5BjyC/ATEnRec46HfUc
Ec5uld9+znE6gcEQRrZQ3d80/P1SqD/BIq4z5qpeOP0GZZN+6rFbgL4JPxMV0EXY
3B7wuD5/4YjsXvI2/XJWFyUr1j016neKV9QslO7GVD5gVjWe94t3HvxoQ9HOly8n
IvMopP95sarcupZHWRtEx0t6VzYD21LH18cN0//t02a/00sRmmQpZLYfXOAVU+iO
hKCnfizDHNKTB3W3d+01tde+w56AYSXRuEW1ccD0VaHVLRXDZgNmdNL3mLk2as9o
J/Qz1bS40YzM7MRF/HG5WIFVhA6XhMradWvENFQMDWsqiy4ShIVi9Yg4HfCLDGQo
tYmYi8Pwjysp4LOHfvDW3bwmd0aEHB3DArSGk8K2c+BKmmWbXnB5zPI85wz0v6vD
N4uKIFlHPkJ4OAEjtG78QCdSh6ePI4A8BsVjczQfezZ/E56nmvHdnDG2ZyQ0HKo7
lT6AlGDZFFUnbv6OEoYWN9Z19zfttTOiDm5zwyuH5KBLe6jiZxLY86KUZ2sfpWEj
xsV8MYQDCNuN5fYEhD1G9+JEDjKkR1FV4RZ/Q15BvJxGNgSnRp7G3ywrmR6VVTnD
Kd+fptW52UeEnkZdDIFChO0cp2NQO+xkPejM07mWIBzDMP8/VG/2KteFOrkVj9D9
42FG14nNzn3pZo84vjSsoTx2a1W9BbpzlbEN9fGuOeEiLBieHd8KSdJzdlvTowSd
PUckmg3VNlyy5RGSXW226erUrvX/1XBOagt49+GSTAVp3AB+0PtpzjSxjfTXLfeU
uqSMAvunG+hEzkbvQqIer2GXuxb6Jy6348ohxa/b0Zv3c31NEBDrx8JCgWwOuNOY
M8jsgZNmAK9FVAPqoubYtiu5hBADm6JwrXkJeRksECmAcTRdVjHk6wIpfNGfSfah
LnKLQl1k7nE7FW8YC8RxT9wfa+Z/eeGdQoqZmjixThK38ea6syWb74r3+Dcq1Lm8
yBx0nvmRoltRk9jBmzoBnRgvkBGqPhg/e3X7C9OxYu5ediCt8FzC0M50QYxyl1lE
9oD4g6SyvdcibriMkeD4JYJNlp+CYxqfLEf7KuMRN3Rvh4/9akzGL1CnMzYgkaCP
e/fHf6hSmG9d47N8h8Uues7NbwP9miAHX1A474YVNm50KoTWgK1g/vpXmOYhcP0T
5fUmBxlTsIUdQjUrV5xBAHNw5fWu6pcIk7p2Yge+Q0XcYYWIvu2+2VWG5yy8M6Ya
AGjytYHRmmOOH1W+TK7S6nD3T6GupvzAgkTttngWKVPYnRbAg9jZ6ErZey4DrQHn
mIH1CmpeshS7WDKivdJeR/OnPx11gQd8f6d5tBz2nOpeOukkbvFsg+zI4RK4P6mo
heSRj6p91a03zQ33z/iwojJZ0OkKMGNWjRqOVzVAtZpIQJoHMnqSnhtZVEGQ3Kj7
V5sGI08X1Mw0S1UVPy35/hOr1DsQFxt32C/MDT0MiUr+GXUuC9QtM0qIRltOIEf1
/UB8YHdERc9q70RQc3V9hGkzvgtkQC3jk+SKJcecLfSisozNRACa/63fYHFMDDzh
9Tglt2nQrttO5mqlh0WciPeSS6iXTpgnTRASSWZJqPFfP6tTX65zHc6CmYyhDTPF
pU5giz0Nc3KgB0oS8evraOsDRMfoJq158c+ooxYZ+ELWnNrKNj1NCF/9F9Bjn421
zB+HIVu06xz/vSd/qMIL3WBWTbWlDP0b1pXC7sckThJM8pYGUfBVEHSjouzPIpgz
8DzOPR6sWSyCbdYwQoXsNyS6TLKW5tUqij84j5jSaj0/G8h+3tnB/ZfVGxoviXU+
a9tstxf+3TMlZCmt19HjMclT4vRIhSojzPf3Agpz/ABM1cBpFlauAwa5GLErACJU
l3DR3LOr1TTiyEshUPA00ooGNNxxNjRKq0KQyZ2Z9Lz/oD1bRJgAap7u0Y3XXXOc
WIW3JJHgTsEdWO7H8gfIbFCH+dT7wW6KLskATaUwmsm5/rWCcc87aYD5bqDkXm4y
2XeuJaNC3qy2jafjThazg1iDp7DMbQTABruKgs4IvnVbslcWVRDy91EaEoM6Iljt
hSjdXI+SlM3NaZktCIvjtAvb8JWQrJI07pDCXbSNvQTQyqhn/Kj7thLXGLAHLFuU
dtaJ8GPPeGS0/THgRF2j/p1dZcQy2dGL8zK9x1PSkQ7tuirs7abOdaV1A2a2R0a1
Dv4mSXrgtrW8xFazkByb0HXbjVkDsP7L5MOmDS59OprTrvPdmxhSA7C8Q3NJuZ8G
Mu6HaKn6hFGeG3qAtRdhz+XHQxfIm6iGn7iizV+eCEr6ro3CuJUcXXVmrVBg7XlW
GN8z+EkypuJIMfERY5Ra3hMMJBHCxBjqM9BpT0P1LC8I6t506cvF6FSgWcO+zjVA
hNm9sBobFn8+8Harn8IdHDYmdKBndB6nR9l3+9G6jVip1Ctfm6urE2oRxBZkI89x
mV6CJeaynfA3rvl9zHf3e/shatpmXpKd3izONuFwtZweOV0whkW602xSxfL3FDca
L8EDoiGQGGh8JPJwBL98r9SBbh50iFDtbIWydbMs/Dd9QHQV48txXlYXKYZY4TJf
Z+I+ud6UTer0A3jvxge/ZQxHoewzg9C/gYd9AVL8K3EjWx1EFo7byPhZMI4/jX1g
qORF2MoxMwgnJ8P0gO3vYM3LIpOraU2V5yLnCYMDc7KSH98/vKlq3Exy9ch/i+T/
9Vn++yXnRILSzru72dcfg0PDaTXQfiQApc28KbAW+Kxm8PcUUNXmL9nulRrVlSoI
kNfgIJ0knUd2LtNaQCCnXF1Xc1+RYERdGp0qJA5xR3Yk7XLd9NOMx+kgSeRCp1iN
u1wXFYpffxGPYPn5KisQATlDZfU0i3xAQOnWhTIGQYlIxaCCYTkztIXbuuSMcLib
6oxY0aPOUgMOV/CpJZ2MJvsz8aEhOXu2q4Wk6DQAw9InO6pAXNwcgDB786UbK2e0
ROlb+JZ5ICoHQzFu9BTcl9YrxGinsXXS0sniSCib1PpeUT/y05rFnATMYGG3mlno
fK79T1aAy6UyIvdCo9WCZoDu2gWvUK/tiLVr2JM3XM+34oOAln2JZDHaNVTYmTGu
nxkkytmxyphFdPLq49L4p0jVF6hq+ck1m0ekc2TMIMBjuxdQRpQEYYeo05WKRdiW
Jo9oUoP/M9q409aB4Rwp6xWQ+CxKBkmOWszMedo9C+gTqMwMiSNAGfdiqVWkZwQu
yeMvBn5EIdCdbjMPSQ9+oOxoWWwaeBiICkLyyL9TQ1OoLrkfTDti9/UpW1YD3w7+
EjAi1caePX52Tih3qOSIKUu404w5Qlh+OKXzhKl5FDFkA9H0lbmNN0dbKgWU9WLP
dsuZWuzOJ5qh8DG07FwzK60oiSbJ1LVPrOPUVHZx5RUoc8xFpKQhbWkn5OYDA5B/
1BxNv+guOBFU4/rDD+KsyypgbH+RAohW9r8r7cySYnMDnhijEb45gEmbPV5jpLsX
XaHo5pa26VkaNh9KHTShyF7g4JSslpt0bg3ofiDfQku9KfiU/QeYYFjK4TohMDUi
D3gySg3oupL9XaZFmGCtn275mASjp8MDIQV/e5L+UDoCLaGPebmTzMK+QB5sun1n
wek73m/YHVLWhFrnGTz4KRV4AyWc1+Eg5Yrq4y8RuDzQcQJcxr/mVuLHsqJGwkiK
64f6LqrN40IwKcsFKJBiO9MLE1va43dBA8Y6v3opBPT3CNssvh9zsAglrCNTWhap
JfvsE8XHgdJzVqAphA0jm038PLGLTMkbKl7wcJTgz38wjWbIzdst5bsu8G5mbN4Q
IXxX7CH5XjtWRWM0TO7fiOzMvjeyjoZ499hWmn3GX5S9JgbBdppyIKs53ERudxME
N/QWPZFK5+q2jexuLs2ewLr1Cd7jmZXV+POrskd18fBQZNerJoeID6lRPrJMgeCK
tDFnaoXsLWIlI8ZU5ZXkCL7khF4fhMLrjUY2eDCcEGIt1zfu9yHjUOgcCufwI/bY
QyOQoVSg2iI0/ofOb+bfT9DabQqcpfRhnlnvhHvWK73DlPErUlYgDVggsa1LPLPl
9Q/DP40+J0Qs9FqJ93c3WM2I/38Y9ZQctOJ+rp+1zg2LOH068bi7etH5bTdqLJjo
JtZdfV2IQsXBFs2CiZV35fNC9h9YsWh3gs2Wr/aoVlZ13ST66cpJXFOxPrLCEWXv
holaB2Z1akPrTEWMVoy5CNItoJVkvTr40KuprwzQZRVIdAUnodZsphlJRFnY/g/e
TL2T7doVJA31EZLoe3696cygF4QHY3HKBcxp9CIImSd7B0OkIyAXhat7oRfW4FAM
WziJFBSqKmNFyUqg2i38AINwWWS2o6B5qjDL6YaC0Y3HkChlqtYs8fHWGDcFHC7N
TXmrow9PzRwUttmK4ygNW6C1psBYMQzqS1e7FEKBKJIkJ7wMsdE2tQ6n+UF297jy
mqr6rTM2Hck96MkISHed3AT2ciuWmA3Vwh+KcpELsXx8vhwC92Ykvv8+qraUAB1o
aG5iSG7qWrNx64RgAknL6v5PGk9XqE5oIyBlQ9UnrCgEQ9NQbTTsUei7m5GzDXj9
Qswy7NZuVfYHtGLm7xG+khkH7gZEBQQ+jS1Md0gLq01u01WmPz43jV+/oTFwDNqy
/6/dne2eRuI+1MOAD9oCQvL0omOmmLuThGnc5FHJl0Uf7TIsjVZtVpCsOvB8vB5i
Lqbwn1eoe5cplWq5dDIGLd9X82lNe69+TU3g9NX6W0eKJP/SvCCPY4eS6ZDoMMgW
R1Ta2rCO26s/vbS4GJW58bFxn3Q+MLhCHMpx/r/2hwa5nT/x5m9UT+euYK0u/pD6
kvOS1tekjbuj4wkf0bj0p0UOCvrSadVSEcFzHG5BrBVreRDzb1ckTpzXb8x0tL6r
BkojpU979hmTrY/HxW40jPpvUFe5GlKpA0CXSXMaW9cHesk1WqnnkbElylL4WeVh
YfeicN1suuskOra5DS/IqIvpYkKt+MBHA+sRnUu8w23wwFv+WuWw2pOesVQjfNfj
mmqN1aXyzkIaOvRUbNgDRN7wEW9RJpGAuuJOZ8D2CfYI/8lvkdra1GEApYPNmuaI
LEEY8ACpMMc1vjM8zRkSsyt832xGmP1Gm+kx7xq+IDyUxPCkGsEruFvZ3Cn/xV0a
U4Hf4aAJPrwI6cKRsBi4jorC5dmKXIYYe5ORJuWz2TZmQsnqDkORHldjwcDcQf32
yi2ZpjwyJsTl3dW4xYuTW5LVF1HoUA2j+a+PYlBwtP06DJdqgSIDdX924+L9riG8
xBNJN+rfP1B5JjIGpNM/tvfcJOCZA0cOG5deh7Fnrt/uL8M00+S2Neu9uJtQlkNk
Rl2+DkDAy+1CmWStBz39Fr2cS5hYAaFFOz/MCiL6FW+Y4BgKX/YPrVMd8Bfn1dYs
BeAanirGk3totA5V4FNmB8LiiBXXKyBnkyGWuGiLdqK144Coyt4X1t9qurN2v+iR
WkQC7tnrdU6APPD1dxczf6EKvEj/IrVAz8qGWEVMRFc9sG9dEQTfH6NZqHn13uIZ
6fv7qtlH7gsAc7MRi3QVXtsg1eMQdUzz3n6ysryRvAFjURvl/cg5HzvvIpSG1/ui
GRgNz6Aco6Wvn/HaH5JreiOE/CJO5XilSxEb5qel5i5fzGg8Uk83KOC4k4PL75NL
Bi4CCYDql2waJ2Q+uNbbtc7352PnzGISfuQDsRFvaD1Dr3Dgk7peVlx4lzdW+KU4
xWBePLLmJViiPF+3P2WGiD/hb7UvpnCWsdoQVPUp+xySN8yeDhJGQhAh78vP1+Ms
3lhIsNZVUtIIytnS1C5MUuA/Kf7pmlPjxH3lZiEKuKZvnaOXnJ8dTonlIPZbjfX/
UqL5/XYPD/PYJ4RSLZn6BfuE9hhyIn112MdTlhriHhkJz8nEtqVZcLCCj3c+Bm0R
DhiYDwqCgDC4YDpCqTaafius+KH+CaauZ7KXnuvj1lemvQIjm58vd1d8yFG8L9PX
FZlJu1mCwotMHpQG97IBUbLejNIi4MlCqgYY9WJMoN6vVAxf0sehm1XMENsGSA6M
zKt9I2FLwpD3xmVvfxokHQ5PMlF1nhT3B0GkTqXUBN3U5rlBz6yTNHo1FV3IyiCa
lbwBhaqrCX8hQdonEgPHtncx08IHiH0Zmy9sLv5CmIk+CJ0dPPL4a09rPmRxjVfd
HLbmdCBM8EYrgBHxETNYkk/JVG98kHeRQlfnTjdJzBtMJ29/jMn1gRrx/V6O8AJe
fvNCUxVZqSd9ytqCHLdlhZw4V5PO7QaSjN+8PxYkbjfIjkr0EaywX4KA1C/QEp4I
bc4RNGLoYdPftMEVtsH3GdtmJuXSKU86TdWqlp2QiLouDTX4OMv8ezRNxQYKtk8L
0J1tKrarEvmNZKywdB3m3iPMJppa361HP63atVhYUkWm1FXhlwrucZ5AJTFoUaTu
dSDxyhZ6dHdrYc713bb12xpQfbSdhVYSaJrKB3TCAimlu75qVxMCR0GbgcwSzyCx
e17W7bzPiMHSgva6kz70gwZ2U9yOApU1E/I8ifj/rHrcAEN9jYfG5wT/UX1sOk99
lrS+PHjC/EoCxikAc3kuxGzJjA55bXFA9qnBz8U/+LurTUfFFgoE8h1E0PiRw8zb
bU0ZH+rjmZIB9hRbbE/oWAzG3h40wRBXfSBLXT8zd7Iguul2OYrObtYJDKn0wOng
k5vjR/gGoAi979fOpv9Gj6Qs3+48s/rpDI2UsrFBCk+mjOpGZnrBfI4KQ2TgFELd
5/ytqFdk7LPTdhx464nVe+2nWSzWnUC8jIR/lPsDCPIUXB2WccmQWESVKKpqnPZP
yYvWDPSzhfjIVMbYL6g6VcLmEaBOlF/deCsgjmw4Mty0m2uNXW3rnrH8osn0RUi2
gBxaAAERKTR8fFGi9RKvyw9RFUQs72tn93ye4+In2qLS+bzrTlgL7nsXdTnpzk7n
1Mj2Vqh/OsAG1rC9QLXbdWp7xdaC7BiTFOt3iSYVFNIZy56Kx9tTXUH+n10hoYZg
BY4xEh2XNWBZRvlnNF0SFERtAEBlirJ0mnwf8PBqVg6Z6bWOCs7fa2bKLzPpcj3R
/2AdRvnURqcbYRmcX9nI0RhPgmVRoFjPl99lNwSMoKaJ/E4SFAv+SkS+tl1viy78
OP4GOoeb7jWrmswS0wxfm8vEyGopAwL9YFPiHhBf9WhLFbLJFZY5wN5UU4SiLV+9
Xrt7GrALgLFaJhcnLreGHg4cpr+2lD99qglu23YOV8sZ3cojNQlw09X4x5OtgHY7
eky8YvUME8EN5X84b9sFpCLdPA7EiNa9PhOtgupq3/EZRz0VNfKNNd90c9FvXdFx
I4SmeDf1R0zAT6aNHtxyYBdAMNUqb2OR4uS+jsr6pw6V6i5ovNeqM4kOPBmNh+XR
+5UJb+ataDcxL5Y7chklaWCFAEXrQUlXY3TzZRTrqEQVqcP7KqCZZZHCR4rVSgWm
8ZM1dtvDx4iEFMAWa6AKCZ39ep2vlu76pMgEJ4z3Z/5HEXXElBZ4UW32bUrsiti1
I2dGe7Tl5M4y0MbCv3p2suWeuh3+sixwvqU+L1P+zfDKEkVx5K0fB0S8zu/+hU4x
uPYWzeryn2+7cME3Wvp81AcP66P6xj6BcU6gTp+hQGfMKmvYSHKnHOag8gthFsWZ
mXCDqz6ETB7hfro009/mKbg1qFeGXHfYcQiLg7Ooa8z5kxFpkZk3OdAT25gOlJLl
jNvebvWtIOL5aSaDQrWCs3xEO5lT1VR7SO4Wn4crBP1Hscv5+V8iIXeWxR9bDNhE
4KzlY4ve1DliByjBNRvVhINqew8btonaFEuWuc2VSVmvW/3LngDZWnoHk7LVKe7y
sjLgDLa6Z8Er94DXj7dSmo2cZb5OuxpJUhxBNAYcPriRfdsW6VJdOzuDAxw6sV0z
XGgJ+GSK5Vny9BWu8yXw1/2i9cGwQRBVoUm3mVJYNFIf3lY3rUOg8l0TbxaAWvz/
zQdy7Eje83L0EeLj8DLLd8eEJy7T49yjM6LoJrTzHPhQYNGu7LQmGqu7CUmS+1aZ
wUh03ZWnvxU6cL/93RILQyyrmsH7HpNJjuACk0pJ6Ia8G5yZB9UDSgb7Z/ZCNa04
psjbQ0BtlVkonQga/B5wyktcDJ8IsEIpbUNecA3k/XfoMz9lWvnAG9b1XQvo1ZDf
ZP650VtUvXIRpmKWxtEgbDfcLMC9Y5DjNZMJMy5ouvuA+gplyaqQk1+HeTvWVfPl
0PKr3cg/dPSpDIWqpgzN/oqtX0Hc8Cx3Up4p3UllCcCWGQ9jHRtnpgQFOb90nLfI
N7XtKnCMmWWLywnLv1Z3/ZreD7NYfNJTlO+xEmmsGUBA8n47kARxMUXQ/L+25cQg
FFj1vrrIEaAgzOe394ZJQ1ION2EoDORF/EcuTwKdgJ58xDmncso3LcIel4RT+fvu
GzRTL/trhXglfSu5g3N92KB0EXk0QOo3NU6RYttlty923JW5O2Vrz06PeODmUgtu
Gkz6R1YO0vXpHzfOYmbqRG+GV6WYbJDCOLKgmoAA7L/bpfmL9iLpYDO3Bd4sC2ED
05lgq5dnV5p5QslQikgd8T90vCYslo/ZJ5ChLN/l01AW+yYhXCF0pOKn97diop+d
1PU1hNXcAPLAkLhIQ/QAsfX13HOZE8GBs64C+nFc7MZ8dtUP9FlpSG1GDU7183CZ
GZ/UAyZFJfMDIVCOJLqf9V1Sn4IUPVZ/bqJ3D2hhXC/ITlWeysJ+n8WJN7EAptt+
WqIG2ekwaNUwkWpWVXp9k5d2TL0dVE44LBSUFn+3vCh9UL3i6ovF3BcpZsOolKRs
sBYCpygqNyMQWDkg/0A8tNxplyQAIkFREXrIsFiMQqDok70Ai0imgStDv9sribA0
f5b2viNA5gVqxs6oNa/QbqbHWJyZWPkeyUHnqcWbYtf5Ohww+OZgHS2N9P60HqzF
vquDx0AfahutPTLfobrG2qgC+jIMDOCDy55hVT68KqYg8Vz3ggTX3ZAvxueoxTan
N7Eph2W9auM1JTizbOGNlb2P+O+6dfHCkhYJhzSEepn0oAjYKKWnap008VlXJs+V
RgzyaO7yMiw+vzXo+U5PnMduFCns1fY2Cawfp0TFFQhcrwQ/D2lhG6MJxNxfCHgt
eCScR94hmIR4E8o1JMlH1iHZnSaWrGjRGhIqPufKYoqAqmOkltITiz6gKXr3CsZe
/mK4mvC6neIhaVshnCt4KGKOQVQocx2OcgPZ+uvE1y+F2j2W6m1MkU8YnXGMVbvt
H/mdN/9eDnKwQjuSvp22sh1wrY3S09+XUNaFuLSjfHXTZOJDgKpjL1SHz3kRfjTw
N0qApZNIY5FNgjWhB4h4HkfQjOo553bH36gbdr4MDJcEjEY3yVJN2PCzTGYuE83M
qNfhGdlzkN3Rk4mPGi0WUzRYMlNURDQrNrC6B4CPjcuiBykeQT3Y3N1e0DlBY3T6
7Db0oXVuLtYBYhBrQqwIBkLLnWovEUFRq6j3J4jrTSTj5LHevlBYYBMj/D2BSmTs
3bwc6NSYNv8QZLXrkLqY/jZXwIcLS+SDBlyKaXd7wDD9ihYFWvshXirJ3cyPRQYl
FcH8443/FOcL/n2k5JwTyJFFopSmt9oALYdb8SGKYLr75vORAObzx+inbFtDgNA7
gWhoyt4dTtkW8k5keg5Hd9W2AGywh6tF7eCgU8gKAynLd5D+5QPEHSjlF/X/l3fO
F2Xf0B0Ypvr4DUFCPVNxHJc8jgiSZSkIs7JE8AdLQqlshAcOfi24JGDa3wc8Z7RL
1S4ZAP9cNTrL7ZBmIfoo6E0B4mTpSerSHIzImTKXyAAIwQYJEvqYpntj2HvDyAp+
D4IQk8qJWYPkEuhu5uU14bLYdEjHX7+fslPw3hd1HLhjqTlRADgYbXk7lQseeDjQ
Np0cPHbN9HjyI8t1h4JVchH0ZF1WYCG/5czGKgKFUI7F15c7ewL3L4dUyKX77xvd
bZrFvHdTyjRPPEwVlsgkCsj5ThQzQMX66s6N9lB4iVEYhtOdhXgKg+TZgaApoXAe
2zeBxfYgNEPZ28L8BrqH2D7VugEQQtcOwGF8SursOd/UktTv8bTXwdMh0CGw+rPQ
/Rpml+N2A7PO3iRV2M4LSJRutH0YxiJzuRr6kS7O794Znn0DIcDfu2FRr8fJDWxQ
9+JFnD5JycUKg/quCR3E0xh1Q+A1BX6FJBViG6XT5/8/fUdfeA9HRIVhBgFWRn5H
u+TLVLTsDitqrPHKxDHLwpthGIrD9bKXRywe8d1kYxg6l7KvTIZkcnkY4kkj0lT0
LMo3OG9ymIqyl/lyoLDTAMBntsVOgRZSyBkwzF1iNETWWrR0GB1042vnxRiHE/Ap
SfMoUDCjAA92QQFw0/73aVnpw9RYdEmi4rbVF73Y3A2oidR9IgtvrueT7fQqDJ0d
DLncusFHuXLMhjHW0E3Yy1hZlM12z/TIj6M1wa9/yMNArt/wuxUXclxW7yK3IPpW
b1DQiGFZPAfv4WovZDJyTDh8BSo7Q581n/Tj4lEUSBU+q/xndTncu4bBp0p2L/fG
hVUmxrhwOg5w/Piih5fh6xT96GulaiLc1HG8gFwiKFKFLA1X2XnAi9la6R/h/P6E
cYNDe2R++GYrBlRglZ50HsHs+X8V7OrokCiQ8AvGbbcvd/VtwwwMWhH0oKeCMVKO
rpkOoIlTfyfNL3HsDERw6DIZlx/+zGLoXAQJy7DdmS/ZV+Ju//iRMjcRaSY+4uWO
lwFQ4vxHGWk90rN8FdZBcHDjM6u+XZxrJoLWi+nTqRZaAet8Oa8l1JX43IamCYUT
SFBMeU3iRCgrInIWPCsnyJScwYo/EkE/+KTCfpZjtj/RUzYXJHKt///7l8xiuctl
izP2U9EVSC8f1c3mVMBSwjMM8u/cj25xm0EWghT62ly30fwpTunPyNRZ4gYbkP/i
YmpIv+o2aUKYgym8hlraj8XjV2Qu2RkmgeB6h7d/dnh7bFo8RBy8CiKeHLFn9I76
Wq15tqXSK/HsIs6fQJgYRnfiGSoR4BHEhfszzwxVG/pD3r5i6Dib97PsIjw2PXTz
RMxlsDtQO6Nhd7Wa6uS/wNSWRWBIQUiaiA5yQD4BOyX6UMUc+N8QgSWh4NuxGjoE
yBRbhAv3MwZrKQtcQcYK2WlshhXW92tMcnOkv9B8NHHdyyTEprD+dTo6arpZCPn4
5/jXbwFBwCUSqbanpv+rED9cqrhyiz8L7yF+C7blR8zv4EP8cZmOhyg765RP07VD
Xw9gBVK7E/jKRUD59kBpsg7yDUFgPOab7DBjI8t56kl664qbjsICRa+Aq11Qm0vY
yFoztaq2+uqD0zuyfSQN0BYcrqCZn40RA+Kdf1C+FVBfg9teviJ/ggbxNaSh3mfL
p5gZUwdevv7QeaC/5P8UkhYG6+GYpSzrnSVSjbhXWVy/l8X3sJIHasIYlaFVLeKj
w/KR92RobDWQWCjJdOP5RJoYHXVyt3x/HbTZxnoNcnSJvLc8dec2iE+aC7rjVhJ6
mEky/ElNqEAtSVECkTBntH5xWB0LvwsoQIWZPJObOKcUXRJs1SEdtOOK7D4Zm7zA
JwkQc8Y5II6DL1rsksbwxCE/YrxYY+UlMiOApXBWswD0LuMEqFUyFOS6AfrQsEbE
8jF41HewW9yDcgHy6uWjvzysL7IMc8hbqvNdVzgIhc+IY8c5/bsVMKUXEBky5x+d
+AlK377MQYymNCteqOkZQHRV/Na9McwOhlOESANqbpDRMzfdLZiP8u/AdRjCtZsn
JCVDz0gCVg0Uo3cbMcPEf+5iaHB8vdcpAsYo43lkIJ4X3Dc0DP2zTzXZa6NAn0NI
PgM5Q+MsXCkZ7QQ6GENPaAYyT38i21rwLvNSqXKNfzd/6HYaAqLg5JNhv5IMP66p
Rk/57FLrG0gh9mah8osgzvHPHrgWTnJU3mJtVw3eUhLJPl1qY8htgsZpMplFmO54
1KfxppUQxlXIT3lYv3JlDX7y2niew5GhBUjlGd7W9lBehVvcLsbf65gwk0a46O3Q
K5+AH3UQZFqFPMBs30V6BoIKX7B4mQ2jLfRlvwQC4v5Tp+t53VPLa/hez/jK4N3m
vuGrv4ua5gDNjSHMcRZza2Kzq5XkGyVJsqJlmvyCWyVtGvQENVtwqyVl9RbVS5mA
lQqb7jQ0GFoutOkgL7w/JOV6BwzjOOpotcNmqRSWxgnW9XYhygfc7kj7ZoPO077q
Th3mYzMydFFV2fyYmizc6m9UV/5JqW79STwLepqTvAEBIgEFzYmD9/s6wV0oTtVz
cldlQ2mcyePXKWInClE55yLCXrSAY7EcnlacMblbcyaaMcMtd+KB6I5H2PVKi3jK
jKx68sogLr+nlTCqoUr58kBUrxyqkKEI1jJtjFRDkhI9KMsB6h3+gkFmVFtQcigS
NCOsbIgD2pCE0h8C8suHnG08zodxtVCZEGDVS4H5XxdJKBa+ykvF51frKqMCVaPk
0peQos/cBj7RAKOfyA8FgoCrRHpf8/aQXtRo7pmmYHaKNxMYIs00X1njGcMop2XN
kVxsqDIqOSlJiGBjAUyjeUWylzvDT3UnKV04VaU//4IjqKP9IR2hRb6VX4KGHg0Y
03x52NxIRkvH2mHp0GtbgxS7DXE/E4VOMxdHIMO3GNwQaWUKqNejKvbIphtSFxmZ
ooPmHe8Om09C96XXq2SHESm/0RZhj3UPi9Fy/iW0BBeohOO74+xsWaVUjJJlgv64
eu4eKtGGtCSQ962CkgXxfwNlsHOVLsDGbSOcS9wt8idatJOyjVWj0WZO4/rDI0cf
iQzy7lgTzRxlO1Zd65Mq1ZWnwnRLX+yywRaxB+dsCNNOKr6nAL1u/ZXlNzhS65kT
uxCjehj7Fm++LsJETa6KTV/R0wCZWIBKM3Lbegxtym6CnyBPYfAwhQQF5gCGVwzq
FI4wEnnwnan/V6R8yI7+3j/fAp+/k4lJn0HMZ6t6u/VphgioC5hhTDD/Z2pN0YxV
WKmJAOjlPYoTrDZgUuwItbN08S3Q4ZuLFEUJVqO6GxXipzarLFuNpo4xRYnaoXPj
lkctVZLvnc88uha2vGnQLrUSv0EMcf4FbNFCU7ofLQR8MF/xlBm6DqkPsG+9ypRB
ugaIrnvL7ZzqhzmmlSu0GZuLBrvKhrysV/ROY2J92YYPzRTmyMiiIbf5kyaXp6vl
C9FLD2UeieKR4cL5Ly1ZR2U1ceLYCCrSCih4QMzj4XaAXD0zCpivNZxDMf4OuCAC
tBT4TMN030JzO2tgvJqbj8djQmyLG7nnbaI4fnyYUIYZof/iS4XknzHYdVP6kfBz
yD+T2yigvvhlpA0SLbFL0smY8XI7jp7LM1pLvBkBlp+qXD53fLxkoYUak930TOPO
nroUlWOFKlHkQVEpNQCRVYox7NJSr4isoklNu2rW7D59QzEK3/+e41cNXYl0XIFg
uhKMsadbMqiA/m/8TqQRWa82/gN6KObGRyTc3Uz9vlpvqbhKAlUgLcaCAUUN3hH3
vjzAXAQZIEmUGonHMbqiokS2v+D7Z3wMJ9VJtWBwTMNPlGbmYJcTNwZUB6ItBF0C
6D3VTqdRWexEL+eGJcGmuiHKWrZVT5N6Gi8qQPoS3sjQF0hwNDRUESmk40dLXWMq
dVi+mTfAqCPBOZ6ObYtDxtduTP2LeyWAGLk2ZV5tUOeCtXLJyEMb+hC9kUyKWYEK
sY+YKQIEamjjDpt1UVNHj/5HU3HZcsAA2SXCg3+2SZ+XXlvs7SwAXvjhqBry2eCX
tN91L1OLHrXTT2CFhFjV8clYf/jem6ru4DcPUh5ZCNusbV2BnioJ41BhFsAIWt5i
V4LwkW+SFW9GuwdUC/14zDWW76zXFqf5pJhvT3+QjGB5YJLAUiEcxTV+eT0ecLY0
+q0POyDHhanvZUHeydBnQoGLHkarY2gU76QfJr+3jb8K/RxmFCsvyacucHsnubVn
HN4w5muF4pzfY0XWBwh/zJ18KPLohEOcAW9NigXXDYizNhYwMpmZ1jWffj7GNd2j
mYLOMa35k/U+HB8KAMV8S6bTtXpUxeNOOkoC++WJR9TDjQSfHGrsX2hmEPPCya3E
7KaYFaz9i6eAv4rgDYNT7jSe1ZGeilPb6Kb0v5fRcLUYdhsm57zEzHErLquf3W/6
CgwTY7Ew+dHOl1Bs7nqzDpXWXpDWv2jMtTObdLEOongKrk5ckzZycVhBFdB9xSMl
/HM/mJh7hnY1XfQ1KQ7W8snquMxi4tBYZbqbU53vLX4/NwhNvuDOYBphZLB8Enkj
n/G9ETml0Ho477by8OlK3Q4rrUww5F+qUx5UlBERtHiatC0kIkPtb4YB+Rq6qfGh
Av6SQPrFdU6+OAOiTEZlxBSCPqGA/3nMGInGwzYSPmlG4la2AuliSPGJhfcOawvL
Urj8VO9Pj7HDG6Q3uN/+Ej2JSl4NyLq1ScuX9fdoqoRGhjHM/cNffWBepUFCE/zt
su0lmx21agPDDXhwOFY9zEmvA5YOyLvp+ZuAKj7SzIKHsX+vIISZzGxTRxzihzPw
5Hk/YWnKLshm9iX2pXJHIG48oxc0s1nE/g4we4gX7If4zLhA6BTBzyXVwXT+yiES
t+Wz2pFUQnq3MvzuXEcQrWb+tV9K+jrTSZ8T8ux6G3+XBFjUPiHDfIojyQ3grrTo
gZv9D1Z+GBLZ7MFsvlQ0slqZCJW/9lLcMqnXjCjyTkTMlDc1t6KfjzFfLNlnsCWH
AvscQt+lIk1RuqJAMS0iBxrPqr8g3J1lfr7s5RwC6r4VFF7Q1F/tz8HJ5o6gK+V8
ZXJv8VafLsta4tuSzRzo7qX3nXSWRGf00IJPEVYDQcQXjzvRSU3zOPcMQhdu5Zk5
MydPwFW1luihh4DJ+mnOZXHZDZ0hjf+8RNqrKezyPWp2pCHFEaVcyqbIAfMaEwsY
vIkWRkb9v7QFMaoWQUVMeeM2w5xk7clpYmkXWT6Da2ctkb41oVBEhOf+PDJZnZ62
Y2Vb9DR7/DZn3/nv9XKtUxCOwvXpqf6op8bD+OvCyb2u7OOSSciRl6lejxrgWrcF
YXLgx1wEEeIGOKx4zmHGKoYjsUXuUR45yNReCfNuSVekxcPH7wTzrxx8e3rWCchv
4n1zN/PV4ouLFPk7qhwh7Xz1Uidxx65giAySC6eGQjsR2dvwyjMEbfzRoSsU9GpU
RX1ShVEtP1fNW1mxIctJeC9OxKUWfV6bDkxSKsdpYfAS8JgMOJ2ur9sM8Oj/BGAM
6bvq4dyAyEKnS95BIFUtS1nE4ISPydHCfiDBTu1ZM9SLCosouOPpeBJmBRFcAGVF
xw7gN7rRWYCJGFSro8M6v2heBfQYrLmGWB84+29+TYd+qKMZMEIaZCLvaUgxEZ+t
wKBeUd8NymBQa0F6dloufE/01nLQP998UsR6GuIta55CV3v51ROIHayxHI5DnKSe
4DKMK/5p7GU5tDC42UNSVOOnBmspfj9cON/7/kQWOSIxzXqtFc+qj5zawyWVRgvK
wwJdqwoG+Mp3p7yBmjWX4Pqc5N5uDVvEoBT9sq3CV9mFJk1ggB2Ide1wmwSOWmcR
NfQ8GyuFHMY4XN+KJcV318dQvNCBAnDEK6F8mDx8wpjherhWHwR6FI9ZcYHOAujx
FK/CHqZckG+DMBveCiYarXcDftyOP+txIFQl4scPT9jdZoKqdz9yl9M4Ut6oC5Qr
HUCDlc+WPNsC+As4UwJ7jlk6Wj8hS16QA18JvHtdIbfqjnlqMx1XMyKT/U7RZHpR
sAgLTlEP+Ks7G1AyPWFXAdttmDfLnpDPUjKsLklY7mNQKzHiazdjZGkeFLYlUlTm
a2EpwOyIRvzhvmIGTqH4OzWLyjJDGrNwu7l7/STJH8erH+om6CskxumxnCbG9Ha1
DiUBjexGdi2baT2qHCksg63Hz0pFkcbvbYPbTeXl9eHdl1WQcCfMrwG+HKGUQZ3b
2dkArvtCaL5kenpTTzxuZCMIKrExsPK/DaC8794ToZnKHfQ6gHEDNT5M+CgatFQY
5RQMB9K58+LLpixuII+knO4C73MEuDTUGrPs/GS+M8a1hlPfBO+PColRna/PtsQg
yX18MZ76kIc9e0qK+KdIs/vSmkDyHymDOsqHYpsppSC57i+SBb2hhVL2nbSL+DFB
IBuevA6lE8fRWhoHpTPQWoSH0RNfb/3OPgp/18uys5f/JuR3uvIFngZNrwL54QMK
Zno9pPhpkUZlEXeHdFV0WwhANsj7Q1SMGvlie8NT1lhfkKnDg0j7tCcYdwhW2uH/
qbBdACvg6DIQqzVMndFuKah/snKNJ0CoyzYcB0NYbkt+SwxXonyPX2JpIhOuig1L
zsoc5oF7cTk7ijsawLGIkgWuTEhfC/9r/zRCKQL6zTh2hTF77SyVRS6yTxWxn0jb
BynK16Pv2wJeS31HNrGUzfZYEeZHxm/DwJ1j3zVK0r6lPs1RCKp89yokze6XEaaw
OqzIuyT1BS3VVeeizlwZtc8jie0LigN5YHKbvUaL1BN6b2qSg7GWEXXP/YTkYQZS
EonH4coa2H8ZuTI1kd2X9ZpcVJjNUhQt23gHVcEeCEjc+LifbOwz2Bd9xmRQ41Ib
Pjy02zF5qZW9ZxHjzRgRxgdQNd+g7Lszc3Cv2lP+dfM7Eu3Fxw6iMgMh5WRwBwOm
pWNf+fXtNeJEcxgOFSi1Yuc02QV4ZAlLt/Cy18hD4XGv8KKxKfP0KUgYXmZ8jr4c
Db7LtO+svhujvp1F/GoAr6OeRsEIj/bBLEY5aDFG0Yrzckl1bJ1a/4t0jbBrEbJK
kOQ1xOZGONfEpwaiL5xQkIt+huvR+6lr/U0iyIk5sB5Y9Fe2FQ8PM/J5Rqi3oV48
uMkvKX7SuVjlHnzz1EFawwgjQ5wHhrZ3G9uaclzE7wzqk8H87AD9Gnu/BIAVfRNP
jI5H6yMbOInvgQjBkD+DPbVi7BD1MV4xi7ZuSvxP19MMsn3GSctncM/dM0uTH/97
r6yTMlVJ16HMWDIOsI4dGhDHshQm0mZO1DP1bjxYNElSNd6FAcf6c33dBez8W8iS
LH3Dd4pYQc3KJZjah5dmi7O8KDbqYSd6yTxqAGfVl7C6c7l8/ip4CtnjgV0KYELv
bD1pCaY+25deKF8X4NEadcT/kLS9YIjwCqNHIiqGBAXpPjCKZYUAa5U0LB7zcFnC
V87WwPbk+6VeuV/GAEtp1IE6LLA8e/LA0DnggwQrFS8LBCuv4r1NfQ4anJE0Wwt+
39PhVxWXI2Yye4TZkRix0I5X8CIu9PihU6x6NFKeh5KY1wyXUGo+RxCWPqcYjB7/
qB8TFLed0bgSqH91EBga4rr8kLi/Rl53eDAu7yBBC1SLciIS5ply2U8GKtYMyeLz
dMmWGpVdwAEnSml4WkvuZrcg0rnfV2IBMqGcXvIJVOgvuziZncjc9DApw4leMATY
syvIHQoeW6qXaleFceVrJm1njd3WdTw+Y2VKlQg9hK5ZY1Kz5vT7/ZYXfoksYqtt
TL0511XSw5SEmVslPiIlGpcUsTMKALlVe0uNv5bbvcptc3OY4syOogEusJOGL9G5
CM3XaZ40m9d5d7DFqOUluebTimg3TUUvPn6mjRmkGBIguxIKgLTOEf8ZkTk8Jqpa
vG+o9qKYa/uDlU5ouXBVLG3v3h2rvsAtxkj88hjzv87YDMewbAciUnPCR9XnPvVE
IV3DtGb2Xp121hZgYj8v9gcRzFcw1NNCak7osRz+gSjGak1nrzoeH8NPAeE2CV1e
oD1Mr59d3ufMzg+68Jz1qeOhuL216VLmm7NpyzYxsMZOYMeMQXmz5MS7LiU41Gfg
XCmFLpfPSIRgAPppjE92xfjHJBw231Q1NqDFMzvY0mPtDphIJ6uqBdeYerlqidvB
MY9MnzpjaJiNmxGAZjF29prP6m78RRv3muRtWnO8zSZc4RPZUkrCakRKFYRoxab0
bc0ANMasWNvarePzhLEAYLl+nasluQbgjUQeCil922Qj5dtmv3Nw1J2jRxJNS4Uz
clfxjC9y1PNmqKQMOhUJ5ZZCZs2a2tZH6k/RbvfS3ngpckg0XoMwoiopmr2GNuOP
AoEiGHEEgpYMz/jjRki2U9EBjb4DIl1jGeu4nIkE26WTTsJxsfMdL8YiKHOYgeyt
G85YeGnvSpIar/17rBBSeFUMLTIdIuDpZYeU1PN9BRFdMqXWMNRl1g4BWJR7V0+p
+uBZTxqpzv7dxDU5F8wuN7N851dvsbQ63xrgHH8/O/KFqrjVcI2oTFSQO/IW6lNA
o9ftUCGbtNOpFkJPpgHVBvBhmsxQ6C5yuCdeb/hMfZ1BLyHARXqUWCL5zgej1TaV
mYxFaaq5w3LfkGDJ8XUP3+10DykVRHNFUDcOVYZ2qaxvj24X6rdsr5UAvfZL0EwX
4cYMRJjEvRjPzfN+9w5gKDVNgvMYnPKIOXpAf7gj4qNr4mMW70Ctgr6qa2qwlBe9
5iq8yAUS0yhw1JgyLd2dwKEcuNJwQrAptT7dKCq4QmJAP2vKDxZByN8xq2e5fQGf
MOcFCk9XuQbAdOydJaPogxWw2MGh7PEWpypCzaCP/RgJtDUvnYn5ybWY+6ukmHrp
JkvF3PbfTWg6Jdd9Z19hEzlYPAkciw19/0BGTDUTxsvnGqXTo4mS5PUTQheNQpcT
VcWWERnowCIT5hfVmlxtNEgKVN3KUAnkz+0XXi00XmvftgV2G+kMs5tB96sGiCHU
Pe5kNKBlKwajNTP3PowqGYU5uExF+PeDTS+V15OIIhlFiTu6E9Znc7hkoxoUZF/C
0q/IOtZrKXfNizuUhYcBq+PZeCLGbyR4GZSmibHN2yVXwxtqkYKjcM93whjPIfhH
KqnFlHm+pOiWqU2Kp8nmuo/3LQeExx2ysA4gAoFnfmII6g/MWO4h6h5asIx8ohyG
ki+hbE7QJ97fPnKwcmIux97yjkWqSdnh0TdOLpbyuZ+U7HSbICfuOzCY9k/nzk3o
QvILD1DjwoyG1Z/Ku4Ip1/DZqTwqaYNUdSjBzdkHf8bxeoMYiQG3HHaxpTQZtC7B
DaOTCbdKiLnBd6zJTlgbC3SdEuK3lC3ypcq/aoynZ1sPsKjoKCDwQEQ9rjz9h8mG
ilZBC9/DdOhqcscOPT5SXQ0AdfBDRFlZCBDzZ3/JYzmedmlBcTjUUeyLJ+zn9Kwu
KhluvSflRA/eUzdBOS1N4TfhNV/VYzambmZpQLxinMFFIp576IAWjIRCXdXbMjxC
qmtIatlJgIUYjuCdFa60ytJeyi5d304R0D53ZZMKhM7oO5hjjNfPfWBPXNEIIqYH
dVpgSCqTCo3KybH8pNxMCaIeg7gSCYk1znRyVGriXOAN7D5q1RvcPTxyRjjT3TU/
xinZgQo8Y5C3prHXAbIH6wDJVXPIi8N745HCK5IcLP+5A2thdb/49HuWaoSdQ9Iz
q5n45/ixG3409ZndoXEtrxCKKSyM7VOthEAawMzHyEUOk8Xj7pxpgVlDoKKa4TIo
PjFTQUu2HP0lJ1U2NdoWwgKptPHJfXlYDNdg3CxSxOwGuI4l9wzQO7xo3megv0Tv
axA2QE/YQ4YDOGqSz+aqWuLTHucyfeLmZs70tlAGAy1PT8ptvNCbcyq6+vML/d19
7Zr1HQ5CctAiCYfagy0QPkcy+ZmQzv+wXLUgyjScLwtCnMR6VQQ79kuPGZjZUfcX
a2UCHRTr4aCjWI56fXjJUvNCTbamvK90erBp8q5wiRSXfIeGLBe07HRihQEeE6+R
p+TrPrXZxcXu8AcICfXPdeqXMstfpq7BcNHQ5Twq/tByssMUn2frEJ+sYtnifjPL
i0hyWfnz/hr4ZYdl+6/TZ+bKcFYDtR4E4OcP03W/pBdegwQglK6nF0IdRSymNnP6
2EYmeyKBKZ0U475iJd86NBYHCHefcae/3wa72q8uAZ2Xb413mBW9tFd21hRuuh0y
sWNmXywS0fzikZBS/Q4Q++HubDv+oThHEJoTjzxv8bnoozjHOqKlTpdLRd4cJM1j
/JtcIg4ElAC0CeeWVP6TsLvsvym1FqpHvUI+XCriE+Gv3LqqfsDWZz1uantnEYe5
/fkgewCS7N/yyEXU8jUFXY4Vdu5dEwtY2GPPM19QXcQMwPN+L4MDjDm1VWpdM9yE
HmDi0lFOUVDoKFu3FijFgKv46qCcaQDRMGqxjDD7aVDq9/SxlNeR73aQUxb6Uom2
OUlzWJza2DHmZbFbKHHy0vuN7qzaaskvSgNNupQdTzQLReZua3NFd4E+TdegwIhC
i2FLwG0JwkUJ4fa3bLw0gtCXJ5MCAQ8ScBNloojKValntJC9E+Brx/tzPgHrQBia
EeoEfU3cFJpTQVPxLPJnNpAMn6+YUCxeezC/78vHUjA3jNBDE7A9HkBX3dRqUA2E
W/9nFGag9aRkbdPUb80MTL9XS/ISSdC7+y27egdCTDAF8k12Q4t6BpX3yTCsxiYc
TixLPHhL0KZh5gWvLai9Zeq6HsMfPWflLwxYFLqT57lkKYlmWTRT6f2L9R8u9+zr
eUq+3h7ANdr3T44E6fOL/0XX+spuRAI2PWuNFBdA0IyDdX5kV0Zb/I9Kh8aNvvxM
VoO/CLTjFjyIAWy4PXm6Mp3vG1Vz/OTjp6wYMpOszQxURZANGezpgiRvDZWB42Yu
WLU9YPbMSk8A7nj/zmRyE9bEMmCtlAjSPreyoQE9be8MwV8XiOY57VByQQbx5SIs
Hawgkk0xSBFKfqJQg7bylfJMnOJkb9GJopzMVWbhAJmywT5QdUNjV6pJnMEi8T4C
36ERMotRmxj75a1yNm7ti/3klhY2NJw4v+6OSozDilwF5d8h4bvpzISPiwyOz0JE
I6vdQjACzdFnRfV+BCyzXz39GxFfj44AzH50c05yUbCxbqa7Qpf2zNa3ycG7RHI8
gKrFSNKPg1oJKpUK58WBpBexulLMztBamSnj7Fut2cImG3gtMdfdtYqz2+KgNtkh
OgYLtQDXGzJxWq8n2+afhp2SM77mCqYYo9aDHMH1eOmcCRhvp8/kDe0eVfi6bVXL
InJmvK+Uzh/pputRycCNLD2sW9zvfnGuV63uA4MT/d7P44hCUOUMgByCTsB3+Q0U
q+CxR5toGIRfXT8xSW6NfFXjzm+2TFDPKiXh8dHDv6vv/P67PifIGdfLkx2fSoJN
bsO0QTp1Uh7hE9HEaUjsjn7vq8hHrNAxGNZo8SVUcohFinRTzPYwDgYLXR5xha/E
8E6JZM3t+gBl16e3fdo0OTId0n7BUB05UcwjCoADe0dVerF3twGWzlpGAoXI2q0A
MJAGhiDlbVUD5pFdDLawDewS1F2ToOHFj3P78ryexecCq6Dnwyaz1oZeTvpo5ZIX
BvaDn+wNDn1PkAkttaIR5eOJ1//cwQShq/fPeVN+Vs0N6I9R/eriTOfrez9vIZTD
o0lKHlkN4eiHb5KWtCvJu5WtcEu4OqbnqEQREYzbBZ2egk/8QhHAczn0P82tmvs6
/gwguELFNymt6J2fH6uG2wH8rrJnLvIDUF1zAP+Lx7MA6Ox+aNaLa92+XECf1xft
7Oe/Sa9nSkGm0pkneGPtpPoyQ20gMgw4T+pEqwd529ir6eO0NcCqVOnVBFZpVe2/
cVV0e0jxBuSzp3uoSXPk4WLgcflpl1qhcgqqAqgBHuoql712MkI86j5QgAE8Kcju
H8tlGri3AeRZHFW3Xe6su+9ktD4l/1tBCS9jtmkzmKv4GZqQy0gokYDOe2Bw/1WH
MBtzxEQENjE1z74SadhukoRE3FN8iIxrbG+4J2u/5+8mymikOl36KSzeeqexLHRF
Krq5gb1fQO4kJ+ezcpCpAwEUtLPT2XNNxlY3K5i3ztgr5bcnNRq//Dil4mww8iZZ
rymUlLuYpIBEh4BMAZMTkt3xyl7r7yqlk+47hddVTNn5IbYWW6eUsU7S/f2Dnsus
eCyHJ5Usgqc+02LRh7+wuWmSOmaH90/g1LQxxVsOyJ/mcnhOZAlvY+fV0HqcoUaj
6Hh/ZTMCTUhqTji32pu7Ieh7cbAi4lzy1WUbx/dfl+KIJmD/ZvFL3CBoH25WEOCz
RuDJ+KUwbI2IIxQWrAeOWncd/OJaD7eN/P8lIfzu5lq+naX7B89GLPqUZO6ZXfl2
uWgDbyRBplNqJb2X4c9qbR2+Wd78QK31NU+k/wUCOaByFUjHvJsSL6ZTabhiil4n
IG0q4viNjTzdqwbmlWjl2vrODRkEotL3WLd4IlFakCsjn3VXxDD1vHJxghUq7vea
a7YCQ9dGYiUjTK0poup0uxRVNknJ5AIIbJ+P1Rs4/vc6YW/F+3rCclgodIVgas63
0AvkCDtN1a5B/5BSOoaI+xobjNOyW135Bkwh+5lx66iG9Jy1lhrobY7QcAmG7oEG
kaH3LD9UzI7kcUmj58IdjS/Iay9jcPCxFQBOBF6G1W/LGDEyy9ImEDDRZi6KBP4G
Me6wQNKwGNx+wLuL0xMWgHSBddbuYGkzSpqCUdGcHLHUSYYq+G99veEVatI9WU+B
UbjfEMqrrfqQCBmYEYJJmY4xX0gN07S11MENWJvAf1AiIGL2W1IIBfZ8zEhhi7+4
BBv5wodZQhmCYo8dOUMBIjtRDtaSukn5dMmIVQuQOeuhjNkWmPy88CwKRO1P8IiJ
Fby1OhNt6LDT44jQgj1rU71Wiq/8YQuSKA+OQo1ol9rXOCkN/QoWsTk0mZHEIF91
8cYgFk4ZJernHGCEtB2I2m/9lPt7xn7vZ3fw4XYJjOUGqAWsxYjUdReb504tfiNf
EPgcbsOhZFL16WP8kdI9CGQd7H4+r2A/QVRkRYsResK7DSVBkRmvKsOX4bza6HY0
AjdkfWnvwBcXhgj9iPo4WMBvkhXABSvx5/UIf/qtDVzGzo1wwA5U3rqdyjiD+Tei
JhRpX8TD+GO075ymFz/MGZ5+Wbn/fxZKc+Q0/dvjvMYGM5xo6/sLbNN7Yro4nV/k
IKj0MA6ypRygH10ki/+waFqhQxfJt0c2uPr/fz5I0eGCf5CCTL2cg6Cu/2C5wXbM
es6+8BpyMFxgLH4k6qvnAKCYELslTGaHNWe4FVrrbBpKvNZUnNsa3KT1TCB59rah
8VzpfLoBK3s9EG3X3m4qRtcYb2pDKUuSP/MzhW2kSi0Em5IF02mTED9kEuf4+NSr
7VX7yP2N4OPCULtHTlLv6PlyIpNWN9o6i7qnQp/VujcyFq99I1eNT/pl0c3pFCxb
V52SkCD9WhNdHcsDcZaHjb4+3Nk/nDYypgdqnyHtbpzZJCx7WA5mRQi6KwzMfESe
/G7ZfmZLELL6RPqfNtVe0JULtmt/lDMFbAxJd+lR7h/f53wCQIKE8CCRvH69SRJJ
NRrEILbeHmDmrM0mp34qACn6p5bjkZPybgZg1W/uTfZnBBbh2VcsUxIxCaVDUpl7
GJXJU/q3aXkCK9zholZhKrWRCLS/4+uZFsW3ABBLHWTk15KaXhHDsZ4+QqpFNold
/qtz65it7lrGSvRG1FisAeKiVVbsUBz4taBoOCno1DKr6uy7KP2WUaPahrOgMs2V
uZ3khr6hym8l5RQbz6ZjMVaXrq3eiEQL05XVxgTWFdJv04joovFKIBaj4Fj6+HGl
sxGej67SF8l+bdzlZOvShLtl0n9/TrifXzdaLyZi5qtX8gImrIJUzRT9252gSj2v
WLfBtrECViCIR7IhBwJkwWVzj0Vn8w3e+Ibqb1swIeweIDRZhdFNh6+X692s0bAY
UjeMIxjY0OVxE6TLFy7Z+pMynYAQAXKDpgYSj/nzlMCBLT9FkCja9ZC5KerYdJ9l
WjXg2oLH+XxxT/5yCFSIGBJdeXrG/64Gt3VXQ7GttvHuE9/QJOY6NmB429NEOYbu
ShADk7mBTFFfJcl7wAvH3SMIxbZpaFFGrPrTTT5vRoZeJdabAaXj7Oxt11WRYWVI
DLP7D9i56actPWhhBsteIZyYo+9IGptZTX4hqKQe9p+5bBqnHuQH/vjLTAPVMQym
PyaowPRAQ21LQhfWTF3ZnJXT0bswfZwNKsoxX3MXdNLLVwvT+jCL2NF15cP8PQQq
/okJB5tBJc5X1guAkzBWpzk52YKyr+P1qEpAon0uiZ5h4XG+O9F37SVKwSJWg9jb
T4O4Ta5pn/N4tznc0zYE6NHMQxicQ3T+WsM1xdA56SwncOk8W8Iql8AlHvvy4VYx
n6pWRpGvudtTGkQhlRfrgbytIUJJSldJhz3h5lysMKcvkuqvYGmGVIpRHhDh7weA
b4Gp1d34puZ/1ZiXD+A9pw2OqumQXJW8QfVYjm1DF3NSRNcf8JpQv8YCG8p4Jw/o
aqRzBtmc5d1mmVj5Pa3vrDdHa9XZV1MHjmCjOXdpMBRzN05Ys66SuM/BfNYNdrBw
ahlHfCoBdK08CfLbkuHjvyaOosCacgNzLEBykN+Adkqb9Ulhrf/jxQU/kCpBa1ix
aD/N9xw/UnJfe5Ud5CmKo8GM4c9zkufDduJRR7mEXFNVpawPESr1hMP5CyNgdG4F
chgeYL0RILIJ0gNCjIhmUB/lDu/q8oifSUIMMUmnM1i4nPwsqDOZw9WfrYnG1GJs
/xwgh4JegJ6Ikk+EVAGhhthONXAwCyUmfPtSW+g9Cfl9eICpGgJhlt8IlOpzKxHn
k2b+RVZMLWDG76euMa4iJ/WWhpcHE0kxWcbRqEFi/kyFcqkfA0KjbP+xQ0bqcYor
ntejs0+r8D8tfDboISZ+/5MtdIx1N50Hr9ikZs+OTJPJoJsHDacsq61T/6HVs3pJ
5h61KI8jmSxZv9bnUiJgMUOa3alYNVlo94Fgi/WWH/nlgT9xUzOnB4PO2tSvQhKM
13BbTVYDFOFXs1yvT7dRmQa4vuHMh8mtWLFKpbJSXm7qgPnJnCIyRhjJp1J+QrPl
RPCSRTBr7z/SZdLgDaylPNPh9VmG33MN/ZmuHQ6chfj6nYmKSXalIdsiadH46zs5
uhEs74aMzmcVssuZFJfv2cIvs77S/iuEVVMPkLctmN9cxM/2a+iSCmmG+sX4Ogre
lkA1luIFOyoDIJi/9jKc0F6suWmlLIjTUvSOYGcQG2FvWBOZp1M/V3pLvBGEJQ6Z
xbhY/dcNNgvIHJxaYhwcP0lViq8NCQIISkzxKmNIHqe2R+Sp0t7PL4svaUCWCnfr
yLK2hMIjJR5R3209ST0mYZ5f3NbuSHGEPUFQDvcLXt6IRBfhsqnRCrXd9rIUtEk3
fQOOixJT2yfLAJ34l2jeDMRvfUTd0QW3u6g6HvAb3ezcUEKVHA2zps8ZT0Ycv30M
78yMiyNgmbFL46Vlkr8wkPH+oaFj76mZ5Sk77frxLonIAvnpvPhdjVaJ/4YXDsfA
wfx+dj5FuKHiIH2OiYoDEB86Ox9SK3QZM2ZBjnhTX+AVAdtRo92qhR4+XvO4PNH/
ZsEPvkmk3WQtvLWq+ZM6Zsc1VXYVAPuqLld0GxO5p8starEDgceWvpzGplhvW1pB
9gJq09xz1RT6WGptND7/k8gtYxSREDRAYNdI6B0QyMAwAmuVTQUoARbotiy5tyo5
5CjNYPC19dDuFkzhCwS/Z30bxFUW43Fh1nonnJ8URZ46hSJVD+AqUM3OpNHWZqgt
F1NiiIkD1Xd9V22j4PCoJe+7YVevtJLhn3CpOk0NiQt3qZ934t715W4v83cAQLCk
BtSXhuatVpkK6B4xnHSWVGgW664rDehUc4NNryk9TWZrIRCIo0UoDnPksh0do36e
yYXYHamwFBtia+DgeJJkZZAwNKTtbcL9Ce11DxZnefsAcv/Sbk6kQF7p4Q2kPV6T
oKaQmx3Q3llpVYjFYdHC61aXk+mt78hp6oYOEasXaoP3FOitmHAHF6VADHHU4AwA
LsT5gSC5YuqchF2T0knNtXI5kzOZrlSoNjsvrk3tce7XB8ga48nsjRrA0d+QXr/+
RETmTiwytDvrhPuHAgooxzYCz++wm5revMNw/BQdPfa2mRDp1BtyaW1zBtZVSySM
ejS4avVvTwngV1ApV8Le7iN6SVQz4EPwG03VGWhtWDVRIs8+CyKssYyifvnCh5J7
PJhQqK8bigsEx0EeFCLV1ZBzu60g2K4U6ocp4szSGN0vNthnUsx/pFuqOIo1ie4Q
3p4ff3FtDHJHhRYm4QzHao/8wurpHxf5H3baNnvC4wQISEtN9AeVIhJDDtbsE6m5
w1SLM4xiSomYT4ZtWSwWGc5+LIYz9b39yjvA3Aju8aT9lByA4lHJmBN+s5W93SQX
FJoURUiD+3d2aChkxlglxPuwPCApeybiOxN4D3bSR3GnG9yuTIA31eVLJ0SNy3tU
Sw0Oi8zyOgXjKj6BB58DhCVFUmfPLZgJM34VlYADhS2t/GGapb/TBbDmsl1CaH6S
QzRO16NDzfCJvKOyxI9qXFsknlmsSJhfCIorlA+BWtQVxuW2+T526Jp7FHLqyaxq
bbRIsItFYrfOqC7H6BcJjnHN/TpKKUR0w/iiGlfkLiaF2ZcSbTsbK5WbdW5IrMJb
Nu77uTn76HsimTDVohGwTFwAQOkGWPnBSxmnCg/zy1ntukdA6w50zLoBj71kTU22
fKNxipoA7lRt0YxELvJ98oi1ljElZMsRZAABCKxgR+ElKxV6RnFOqCEr0pW0kbGY
nQGamUCEV6wn/hIXyMe3/KSAZT8svnP6vLuS1+of59VEnxZtxG0eoPGXG4uLaLf5
v6qGUNs08b4tTy9qEjcb/+2v2uZuQ2vvn38bJxAqaqn0jUouUlBBgZwvUjPCpkTF
lcKCvpERX3Qa1jflvKMrhbOszQwR9lkNXGP85QN6K6TAZgP+nGLVP35kl/MgmhtQ
KGFAb8lGIkqcftuabkSNV7FZIBlCpos0o1I3FKYQZHx5xVJFerOH01eOPVfF2MjS
/go1ZdDu0rrVeSat0PINRZJJg5GFcLvvRpe1IdVSKunT7JA57vq85nwCucwrG/ob
CSOlg8gySRHhwDP2lamEgqRX9ANnp5tGomLl4Dx70LhGJMndg1zCfC2pzkDyas/f
mpaDgx4TrCv9UljrzNSFWl8pTq42K7JOAI5CgtYHV8OTGaT86PvXXg/J5LQZDSPH
4Th0tJ2xLtSrVyaI7aiQ8GzdS3UaJhhr6IDbEUQ/cLop1qInC5g+L/XiTQj2l+n4
ERH4JALn7Mqd9lrDNh3n+yrJDjA3eQBZKPuj871SLzd3EdyYcSig9Q/7vGVUmsOq
3Lhn/M17k+vjYY4McqlBkHzyA4HCzsIC922wjD+elOxInJaT4qIFlESqduo+MgkD
fubqtGHDpe6bjMlXMcyPKX7RIApGRcz8l6hEWqYkzbjrEbcwpn8NE4ggn/iy1mqF
mkZPmZyOf+0CpMFhIuKvry74Y3/+uWjt4KPzljOleWptFBc9YK2wnxUWQrkgc5h6
+FsY/WYbD1r4xJfiF5MbQXuBQt4v2qhkuOM/Ofk7UOQQCIGr/naJlehpiBayQgxb
rt9p1lzE/VLa31UjjBJs3CXsCaIAESwhTMtLqZ5o3SCFriBnG4CU6trbbBmHRz7K
214FomlPoSUax9trLA4s6tljniUUyjAzkKE9F1Bb+En7p4VWAAmGuQ5yKyh4LpyT
dJZGmiXUFtaKo8/+modyuLfG2iffESvGJ++V98TjvTbfFnhUYTrzd+AmYojpxuwr
WXQNliG8mczEougLbq9k93SCnPP/OTR+GlDtSYtMaW1wSaxDpquURizaO/0TGGVz
MoOebFF6wsU5ImTcbZDFwAgKl7DxLjqaObnxn/I6+FtoW9RJwpgshTShETn9Bdqb
G3dv9OD4hZC8Ua4sEF8iRWShQnsfXO/BCdz8cG7SSXajXndscEvuTgyJ2DIFHiFR
h37Lf82hmCWnx5c2mA+PlrA1+NDug500T7S9c8D2RY4SMb6rlYccDoNUTfsyX8u6
zs2X9WehreHG3jBgCXJc6fnWpPLmYyAk1zaZisKfi0excQaR/0FswhThz9KlO+va
0jOpOayX8Xkr+4dpJ704/5R/PB5KsQkkYicFd2RYgEwxfiqrhsjccHhfI2RuevdV
r5tVhnOl6DAoHC33dXmyqpQ/UQqREj/Bh3EKYVqqMzHyVhXD7WuJV3eUPzThAegr
r1WrJjhUpJTZIOXLkOSadrvVnPKEIAPIqCgo9ZCc+sH55+Mu6zrW8J8ybNbPrqdP
Sv/fGbkdaNhQgMv1pFdueUSnX7k+YWlhoHBcDhWjsRJnZctxe4MYIW8T17azhFyu
ZXOZ3ZC4T9LA0FpRwqNQ89li63/h9BUODKuNNMqnzmpGkFNDePK0f1z3RXoj19tl
4wxcCFHgFiN+Orczr4BddR2ltLlhJWiZLL6Kpo/vlPAGUoVjDCJjjrC6QRURY0kq
bXmSxpL31cXfciJftLQYi8IJvcoFxUfrYzLUzAfL22lEoQggNexZ2tgH+Xcm3X6x
gaAdnLTGiEdQBJI8x6L0af/QBz4NmLZgnutPayh9EKzpkSsVMjKqKrSvSAtRnCq6
O+PcgMUHvDP1aw6N6Eb42X4tZcWEXVgSkMyLafEFSYmpDn2r7w5zChRauJlmpaYH
eOK34tcLE2BveYdpR5y+tPyJMhD7vcRGJfUnF4wctY6OwFdeCocbB2OKSIXMfCkR
ekyyBQJIOkRf6WIFJ8BPMoCVng7A/5t5qmcWFEw5iqPzpZYgGkqZweIz+gdx8DD+
YxnCFYgCrHrxOw6yy60pXtnfmtnt2edDCkc6g8vVcXrwL0BxZp6iHH//Wa1Y6Z+b
P8lfQRg43p5CJW/o+ykZoJTctmm+EZWmBfTI0rijMXgFjP59MKJYEDgJQwNVfsxH
mVpjZMKHaXBKCy8EkdqHrSCnB383PSqMlu3dwvFMjjG/gsJWIHTqaPjNcpXeQv3R
En5zkSh52vUjKSexNhBUL+1+GqQIGuzsxbQI3Cyp5+GsBBMS8IB+refsxqboUQUs
sk5fGEvi5dwJ8BEisg5Lkigv4Xs+U/BgMxBCAWg/gTKp0kT+HnfYZjO3E8TYl3xp
xSLXK+bkDgzhEkxGXt8UY1Q0A2LKkPZ0H+zGCN3uSkyJI3DlwjfsLpPvDg2tELoS
PWbcqy/3PTyYmQk0Q99SograP9rCuG6ujy5+zTKtI1KnyYMIQGHODorV4rF2hP5B
9t2DI6tJJSsv6vwW0kYoeR1UL5mF4M4XCs4qaO6vLzIFibya555k+bYRTRXC7d+s
JVxzeB3bP0jNtiUPgBySJ/8Rwi6gAef0rkffr6dTDcK+Tj0pN9zg8I2orWHNQJmP
Oy0z59X40iesZDHFNbPzZ6CEOGjgXX7xbsK2D5x3L5Vqy70HvyN4r0SLg7Ac2b3p
mXQqcPo+Pcj9vWrItP09buXi59ifGuhM4zFuRLCa12Vfuq9umGKl6u6YrZo/ZeHn
+kwsy5gLPS4Ml50+Y2Cinkm7VgvIWwIi2Do8nUjekq3NLkpc7Kuw2tcDAjAWet/i
7sTFenEjNtD5lvrxkbDAzdxekTgBrBEXaaXBhFrhCHe7XMxIS+xu+S2FdK9YMUte
AqEUtbCEKV3bVuwEFccb3xxVqRIp35QlGRvoVaUFSEpljaquDX425antpsT8kDsL
bgJuuvYCO7HQ5wQTItC2lnU2QBTIQ7uOHONWRXpHfdTTGZ6XU9P0J3NGqS4lWPpB
iJbGuJoHYdbGhLY/jpsKDB4dioVszTo+vFuPryXeXYy/M5DbLL9fcHG2brhDz1J3
jTNY1UG1L4zTrIaKS/L64R3Y6/QVWNEzjDGacW6kdl5aTvg2h4YVI+3LfUlOfzW6
jr4Z0wTDgaESfmh7aFt5lRjD5UTulxF6w33SpyOVP146sMYJBBnnxPsDd37q39oq
lTI+tFRquwPa2YMYz/A2rWvfC6NoBiHRZBkwHrBCn2o6+QQ49NFHwtbj+Ue0+bro
/yWVa1zddJfhm479hnItCHhZlLgWdBglZ0cfOXfuqAY/iY8UwKMgj19IZaboM0sF
SiYRd1lHgVe48Y8pQmkemT6xxWpMwIhkXWsiC2JYvcSPqJfG2L1JCR8sQGSF9TaB
blP048EFS81Ls4IawNj8dGEJO7ECp2zGaJY93Rn2DE+iS28iDYdcVh152aBrcl8E
AbTj3iy0H3/rR3FkF6JCpzHSgrJfAmMtM/7z41tXz5lEKHN2Rjj9CKJe+HcvQI8Q
6kw09d8eKA5UT0x/vVlsaXho2RiHjkbWog2GeMxxnxF1vJ/f85oOqLpX04zx3bOF
yExZlY00BcUo7gNiNtwcBJaOlZDCmdtM5p0UYGszEtWwlUt7fm5zisbS6rAyK/ms
azqLEs6JDKsUKAi+Uw97BflumERBV0jqm+3jMtMpbXrJPlrfCCzBrTaq2iUtEKS0
4ncIMLbesgkolQgXqnuMMb+CSmfnypEdDVqO/zeO9FpPea6sNEmOney7vLt18PdW
TiMzK+RZXyAx+DzntKCrGuZKP98bnjrkLUzkl9tRMjZrlV8NN6Owcx6nr0XuzL4A
xtwNL3x7aQI43DGoLCTvxTaf6BV/7VpCS/niPuVV4AGCk8bNjqwhlQrN7tgn/MUH
UcAl9Fla3XRHpz+hMhSV6MYPUMSHEaXaJ9nMDHIg/ISnPss73rwsQ7zRjV04fm/q
+QK/r17SeJb6bzkoGiGeXF3mV7Yz7wpeyeIgBfe9TpMMwye3aUX4f6ubieez2CDe
ugL0gEG4BqUFEWhqLHxLByrRMmjHScHBQ+qzGzaadHmFyxNpRNXW6JISmnpVnGPv
UJO6DCvXykMesiRed23qHoTwuDYg6T9+TC3Qa1AE/aLGaqKLdLmwn7eR/Wawcawp
3SQKph/SvwX2cESZB8ay3kQYTzOhrEKVEXoh9RyO8Eb+OFGhkd6bBMxKBiXZhbTe
//aIQbjVT6qaz5ct67FwHiFwgtgiw2LZD8vU5yvhFU1z/IAGx8tYUWg6l/hCC6CE
MdhnYqfYZHG7zNxxAmu+5sxLQZ11uvnwt+h4IwhMTteMedyaZJ5XnfYGq85LXTm9
A7OYvZVSuq1n3lUIHyhzveikh5uasHDfxnxYJhrjmVdffFheY/Z/acYQwp7RWZQ7
He5/V752tzVpKhxpoJ8anXL5R31wozlsWkMpecZzGoDiS7j0JIuG5DzIfwic1BFO
RHhtXqWMpArK2Kx6/BE118RIhuQcMUhX5xc7yCrLcahEWGaLVRU96fC354L4dZ57
uT1/CFD0p4j53lWugOXXBHvgLJpuOuKaZv/Kmm7Lr3ngPQEG2yIk/2N0w8rrDbNn
7nKRbbW7yTAAc/dl0zXmn0rQ0FHa/C3wqx3Fc4WQ4PZfKFBz8oYRURvCiE7vfkje
qeEFmXtVoNUg2zC9NHa/ObR9nNgEVmj5drJy40awZh/9svObArwOK/4L6OInaE5e
YYdeld7F4GyALZovLE+uGywMOMzVNF7rKl9bI3SbfLevpdHX6mS9XZ8CMjWNtmY6
SmzafnwsFKQE5BRx2IFrp+U/lcsFfd9/RCBHE1lZn9hMB9I+00XKlxLykXOqMBrF
PH/J2ajZKtBZhSjMOz5ekUyU43IRo9lUtq2YMj1hQXmJgKNvikavjS7xy73WgMQO
iYa7GMD67TMAK9DXfYFqlbO+tiHfA1bDNMRIkggnzIXlsJHEeIUOu25v9fkGddLZ
1Z5wYpzsWSM5jIeYXM+Y7Ni/2xVk0z/7UtZmM38knD1E9Zdfsud7u1qZgPd1AA0h
qTB7WKQuR3pyhVOMkqFBpSfi4yqv4i2nws9ULHohtORFvi2F/j3X69HXkAaqVT2Q
cgGzHYQdNlwNdHbr4FpX/xeT5O4J8AzDzsbL65NO2cqTPAzJ9hz3qeFt478GOHxj
xb2KcaGyzYfKa9DOpscL66uhH/4AsXOVDfKkLTe03ck/yW1sLuKQyOeB9QI32X6C
cWfwHb2Iltp6n0fTT3ILmVgkBKQ0NwyemB5b/WdyMJwUBY0Pu/H3eGV0L8dOrPBB
eOYNdQhc2bXoUg9vVUV2ZvM3UZzervABB4TleSYpy7IsZDq1D8y5H7c6Tm+YtVKS
egeiiVCpnq4tpahW9Kdv88aOzm27spZ3aZeyw0eWC2VMSIXk1w8lSAGw86b9ZNe7
iRD6p5I+3VjNfqHZcuj+F/MvY60BeNjKBWGWorv5OnhwKApNwyeVg2ZKZzXo2VtU
YTkYx/uhaL1Ha/NuWvz8RoaJARn1geY0EM3HxruFytDtFbj60uj3UphdHGZuDeM2
57eNxCVnoryLOY3CRUmiLpzfDXER882Xfl2JK4mAUWQKaRKsvtLBWzCgnU/FRmHe
UTHHwgu+6dPlUOJ7CPXpV5T624hkeOCeNJcCxpsfjx2ZNM4abSzMnFNXNHH2zBVD
8JYQ2FJrQjHsCbqXZjQRNdWGW8CvI8KcaZFuWa0JyVv2t8kjbAw4ykXWt+c6/8P8
/Hfs4E2ESf0JY36vmIFKmgdWEjT2MUnnV7AdUKxM97n0E9GhB1tZYRhUWIDrClQO
SB0GHX6Z0uwvfsNimmReS6faUIFgm6/UrUDAwMnflZp44UZWC4tQc5J4fnmQh7eE
DnSFliCWWk5LIiLNa6rMjGRPCO/o8mmH2VRHcaJRxpwBs8BZFIUb8OnuXxotIYMi
G/e22Z1nsgXQTu4BUOSBRXxlIiBjBQYL8Q/lBcfnKyyOUr0ZolcOu1ZorqGkJmkh
hIphlFf7q0ycWaIEVCbqoV3XkHm82ff0eAnuqNXXz0lm88jt/wiyIzLI1/bQhP/R
Lvn4B91Jw0AHOnsiBilMiODhrk7YmiS8DtXqy4i0srmM6LraBMfIR35BfH0X6iYe
ylkA/5DxOCXod3pj7uHM16lONhqCMM0p2Z+PcRDkKuOAqGwIO8mLmyTJ2SwemQ7K
qAMXLPLEdVrOVZPm5/T8FPSE9DE/y9Iy7FVv7lFxeo3OU00oIcccLOIbMy1s5S4o
BPm1Jrv5EUOGD6AqWdk3jGwp0UiXrzw5Aw26yOeJZLGJb6wLNUwIT2SwNAJMDtsq
Z7YEEHhBuXenEBrjEnFsGkOXKGGXmbkylXrZ/nSXCwh/TVNvdJzzsmgwn98iZO42
P8GA/ywC0NLneDj/boCjdHZQL37KKdKHoDhS1ly0vUbXn20GfRDZBuAhNMQ3BHOx
V6OR4NUnnI5vgzJlmJZlfsyie4o6+rXcluIHt234R1ZBhPMy6ujvDjlywgDwftyv
nvGkhaKmcVoNqEuOUSuAWeaOg2JIeeROwYxKUUQ30T6E/vWVlVCg4QuTg4p64UWR
Iwy7jjFtbi89fXch06mR4YBVyR1aYulhepj2TZeCXX+d8LgLimgp4doQbiILkVU7
QD4RNB2vZQR4TRXniNFEgsyZIV/a7N99Z40imDvYBaxTM9itKRJU7nsoRlEkPKWI
kOjvBJgVFhqgBveur6530wyRPB2/L+wYXDA7ezLtlNe6ppXkiLssMFnlgQT98QfV
5jYtOmaya64l0HuoHpB30WWRhRVM3KBKrp02vsC7k6QJYkiDZXY8+mrGFlCr0/te
Gzos26zwOelXrdymZRZLyoRuneb09tIb9DYH2OzDzF9BFB4ouBzQb+1jeZQPdK7I
j8eidzc7tWEcObHpyhFOQZi4ErO1vz8YU+TOWGlgfMNWE8rDGbUfudqszEBFnh34
KvNhcKtIBGgwSkp+IlseX91HJ8mflCzSdbA7EzfQ+S3qoDjJoNt2KV3WemVTJ2l/
YRhjTHX8DTM+1YDzSBHTuAmZK7CTrWS75D95VNCyw3ZPwWUGExHc7qMZizF1ZwWl
JoKSEdYrnMEtgAASZbiMC8aF+OGrFBJ/WZZtM0RqHmxTdLbPwdZvp+FGOP7qah9u
okuuBKuxgu3IjWijej6T/MzmYb25yMrHVBoOzTQquSNCMUiF5DwMPQriWcLnXyoZ
3oNpLXgyPV94/e6QB/vk1R7Zxthm3LpqA0jOnK1ZbOffXQsRw9uAGV2woeHS6PVp
6WWsefQqfVjF+DabH8a2MEN1uE8MtWWNvPzLNJdKs2YgxsjcfBTCRYuyzwITtFwz
lOkU6U2e4vpBhXSkihIEkcFq3XQx2Yav1uc59LvMN4QDkL1THYraikfRoIzK51CV
DBEsv28V/5V8sYQEMq/RLWAQODPDKFBJnSe8nHiSsKW5oZgNA5D8R0HmznqyvJSd
nNBZBNfmIewWu8L7qCRahAuFUoSvG5pCehZ54M1VSWf5swe0mdQ1TdtBiIwzOXsN
fQJL9gCT8KFH8OUEefv3UHTto3d874UKwnKGgGtfyaWmwarfcKX+yPBvenZMl3k9
hclqNNrHthA0F/QFHQf0Ihbp9gY5UGwh/F5GrAOCkNkmtVWzAZtyeGhKCnCu+v/O
OQZ14IB5oF52OdvLS6k4LqCqwVIzO9xVhL+GtiQpyEG4oZaWNFnuZ25+vJQxwtPd
7nVmMhVcJdi4xmedWd8e8HKSlgOn1sbmTjbW5McyClaSBBZq8d9fIXwR1DzLcCvp
ytYGhD69K9lV4jpqZCv3iJWIB8acefXcG0vLiwgEJlvfJLwReGbKbNR+gp0fc4zc
Paq+d/4wg0WdS+6WiqiML3LMhiCxkbiQdUP4cZZlnOPr6HjDNagexn6cqpcOA1a7
psGLB8YLQVEoMA938Jg3FbRzIBOXnSYu7psg+pTt9uMK/2Knio55+aJhbSMrHFid
hYMiZ9NproCDtl5YqtpJmdN3NiN/b/3PIWCp4sT9Ho0BB4rAnMp3lUmJx5AIfRsJ
dfAspFyw2qsxcMtMNZ0Cm/s51jVnfoFvu43d8v7xpfzTvLPNgIhhUxjqlACIQUp1
QC3UqMmO+LTJpg5MkrcHE/Term+PYuC0uNwF5hVffMXJBiVYnrem67tWUPWk6JQe
bvnlrRinHYrq9O0iCkegtuM0kJaL6yEg6pGOGfC4FEpgWPh8ItNOKHNuzb/4eJFn
GZ239+l3gc+WDJhdi2qKLtj9nyBI+L33tIP0VK2tOfZPKcHx2orLN2fXwMBOL9lD
bZoTzlZr4PmCbO1g6AzLNegwF2qN7tRkDUzctVi4k9ymS/Xz6ZSs6yn3amcE/Q49
BuC9Hg7mCYpe3idVYOBqITM1ykLbr1p6p6tXbdkFIfmgEcUNglF+8ENe0/HU9lEx
AMXdqGiPUHGfb65OoJP2RjDYEDIpCIWqwfLiihs0Q992CUC7mOTDVyi/XVzhQHhU
qN60R+A52KJf8ukbM9X9IA/iaaFe65DFnI12bPSmX65r+X/t/FBsBBnr90Cyqtkz
oTg3hMfCW8q0la/oj9US9JFR5/X9ylxuAPmQBIT8lpPPxqQ1A9kAiMVuObAlH3xX
Px+kH/ZwYZTTorNPK+HFH0tgkREd/4RybynbT1IOqDTbsqoGRp0kDwuiJsOjA0aa
sBtukkStVv0R8ZeUH75ufhuoCI7uads7BD6BLAEkuB4NnvMotzzg0DfeIRCJj+t0
a2P2PkybJyQR/rd0USdqFgDj19rvGsadeobksFm2Y0eWU/lMjucD5IXFQFrPgUBO
Qnz9L+QnOHG+R75RlR5HVnDD91gD65yQTVSpUtX2jXTYgEBumZ5rNmWrPAAeQOFo
rubCickUSc97vjXOAV9/LLwJ3GwpwDpHXQ0ojKdwpOvOzh80Ss5WMiybUhGAfxeP
kzvyXBtxpvDyPpOPip7qDxw5sOKgN5hY/cu9h3Ewvdy34wQwq20N84pNXZ0m7ztJ
4KXC0QN4eREaeSjY0kKNTTz3i435XwIIx5NlWbWFrK+BKjId6A3+3ZrIyt5gdFwR
QXm59UEsVlljdMxsIJDtLeADWZiFAxEQ0F8yC7xJs6l9LSknsPvPNU/c6vRKdjyb
Gdx8QNg3K7RWHTPmafd+NbbivSuo9KRxiWy2HKDe7kikwUSIJTvg7xNPAGXP+6lW
tEVC/YAPOsRIHU1w+xCSaOuODGDdvwZhl/VqBIFSJ3BCXKe/fRwT3gdM/LXyc4yA
eFuUfQGl/dDy02IBjxoMKCTe8eRMcvoWpXj62Tu9dOaS5YJKs3gFNrTw+6iQznyC
il2m38pBFDB0Uo4EtfLlfDAUgHfrsFO5nnFVQmmCEX/cJx0mS1wdzrxZs0I0VJPO
BCn/Bljtta5D8TK2kB/vm7r7P1Ts4A95oEOktHsyocxFIP2e7yEd8efrY4HdI77t
/T3jDjpbmBM3zicxDG4ZKmiGTVoYORXrQQQN+rEI+FS/4wCUXAZshAJCoKvw2GeV
M0lyQrAjn0C4i3woWdVj5b0klzIIE2NSy3kIsrAiDLzKX/9BN8AGmEb7upDnpZgv
SjN48KFLq/JMP/ghcmVeK5WNP0V8jn+QLI4iw/VlG8n7uPN19YqDBQx0ytA4K5ck
OUoAH6/UsheNiK++d96ppognRI2JW9qMqp3pv6H9KBduRk42pnOIrOCPNmEACjk0
lizG5kQGeGu5APxbrYT2UMy8phjcf86tbwC2ktZ2q2I9ulDflEhNfeUqBzgNTUJR
+h2PvJB1Ehs5BFqWgwGSFWLs0q4PfqQT49G9UbZtHYjiTUXyW2ZR08T8+SyquakR
2txdwD5Lt+iBLj4FtlJCWg9lZp1U3nsC3kYE1R0z/v10aGQPs4E8dSGfC0SD0U7O
vZmvoSLm4t8B0VHxF+Ce/1BFKz/RQYlKpknUtOZsNR2Orz9XMn5AwPH4DCSd1exf
qjv/5mXEJPjhp5qVR0jNvyJJCa+d4xbP8CJ2Gx4AjVIJXFoJ9qewR8O9zvukO5Xh
Y5yiHw39rS9VRzIjR2DuUxcDA79FI+Z3PjCMwAkNrXSMtG5piTWBP9t5H22UIeIb
hAV+EdN2KqhNe6yqemgbNDsZhgQM8iUyNjOHZIo/mSXBMIEA3Uc5zZK0FO71IaIA
oxBswuIS92H4oY7+WKtt4GoODW0VVD22Lq51auZzgrN+fRn/ScM9mNSAQqZEUvp/
cdS9ykr2/RqQ2SC8D/RNeBHtQXnFE/VPKXo7OAeXDffNGQea5AYJ6KLczlPL6dcN
u2AhG7EXLBQqGQ7tZJqGrV4tWxWwJqRqcAClfdnZdOl8g9HU2KFbG1gwAURWilkR
HuIfOUdHxeDS3v0caap15Q+tXrtZGhxbQbqhGEiAEgHvcw9Clc8jhhFN/8jiU9H6
zyAJ4Jz9BGs3O8mBThdz7D/1j3y5EotCjPfNkdaNOi4/e9AVY5y2r8u8iMGo2e1O
jODlr1O4G+snzqNrT4VLv72GranVTfk14Gqmlf5qvgrdGWuIVkuIejWFjP3iU9Tv
8HkauMYuecjLNdUalI9YpwQcNd/R0LtXa2iwdSOzAhmMRu9ZH2LnHevaLYZolJ3k
5bWr6i8t/AxFPjd/NobTAQ9sd3HzINLC3WM8wZ2aWNmUtv3r88XyLcb9KeaAPj87
QYz28XbQF9T/PmqFEjhqFRV+VY476fMmzYSq2zzj7OlwY2BGj790bRAB2YXY4poG
OqS3Tg5dZ93lH/Dahnay2+iU490nc7NvWIpwG41bHKDDbXseQkaFAA2YMTCvZIup
p5Wgw6yJvPiHKkvpsVNnQeOtN4NstoMgM2eXqToA6P8/T9zj28KXcrBpEToqhNaI
sndi0UhOcgfhGzSz721flSHued6RSUclKOPZZbMwJn3vSV3MaYKBuKgljZSxibCc
Mnjx6gZcHap/M/uao3W/piloAvfJLqb3Hj+2WZ3Z6sdZtsNvXagEOuzsbSHyA9yv
u02pgfcb6QBBxI+lk4pOc6y1mzSD++rIfSAJ2mcAZj1SWvLsjzPb11pl0U3UzZWZ
SIVQIDMIzWOFAjo5wRdRPwCk70te/eCPXwcLQGpzmpYM5raagDUdqwlxsAk8HTPT
ih5M+2PFnmPiSbAsGikvQ2ZDEgXyzS3UN5L58Kmh0PTwN39Amlwy3GzbHPhkj8KF
7LILJHJKHYEeSyVcRejgXrMieZKRNt07/1IF85ucFQeOEGzClLu1YUS9xfkxl3SE
voRohx/nlpRxKLBCbTheBzRcMYz37TN84mWyDnchrnK4alZqOxS3eGFn7eQguVXQ
zuYR4i4w4eWxAKTqssjh6UdPC6KNSrmqV1JnfHORygg/km2E8XSnSafgqsHUoq3P
44sFUt37i1tPbSgSw85ofwbSUMnf+1EVxtUozOoKQ6m2/V7tnKMjVLjwQ8jIzZgJ
FkWa3bKWCLBRZwKQMPAejpMH0tf7ys9uYIYCrYEeIKtklkkiO8J8jK/IDOzpKUNE
AY1VYIc7w6OymuLa7XDokxBWszzHZEWEEl4Np+Rs+72wM0g5CxKM3M5a+9rupJZA
N0uzMbELir3E7O719WfRDZusjN9/333b2qTnFVglnQcUdIbEN7ZF7gLOy8Ug4O2f
zYtwsKsV3dwlqkfNslZFcq5Vywd9rRCmtKCiTgyUn2NJPgYjtI8CARZizIFYcIk1
k2V2ztg4jIu9rSHWyKABf0Kd64Qk1GBn9Lth2/c/7cxW/1ZxqfV8Ntj/vndV3urj
RVbpeDI+pWjZNI+KsMcUBdZOQpUl4RN9h8YBkyD5av+ThtBnBEDukAiywtjs0atO
m4W9vh9kkEH7qzHK8wjkLfbgk0vBhZa1iVn0UO+hFkK1SbC41eOZuk6dVgld+PQR
jWOekF551xgz9/uvwGtxQdtLucPSFpsvvqEIMgYeM5+5Dk1Bq9+iI+d6g+h8XG+N
sSXKxS3eI2C8r/+3ZlAHfViOvuRL5uNeRf8Rysu/UAbdmamc738SqnCeRjO9piZB
OCRtd1QZZhJ7FJdd2Xeu5LLeejDgDEnVmgw1LPLgfsnggCGp9I4GfLINl37M3luv
1D+2jBlvAjDKm592okpvCdFJMwj1t59SNqoOpm9Gfu7eC/N/rPh6Izmg0rP5g8L/
jb75uSYUS0yz2Pf39ThdvY8Wq8adVIErJuJbzgZN6lKlYT+ptMrYC4p6dmpNDDq5
uILRnL/MUqnWuuHYaqo7Z41exh6WPrdLyDkdrIvY92ZGqL1kVO1dfk3646kxuDiW
PMXmpKBLu2rfI+btUXqqkZ7AyYC844D5maDEa9Yb9P/wFAcOXp5o7vMeMx0P6MnV
8nZRja5zoY2Hpr0fYLCx9JyLoKQn2L6ZDsIQJdN7DP7HCRNkMZV//ILvrl+/T8ca
aK54SqAEOeMSSoZTjf33CTc4BE4r++37VTGmQp9xLBL4gwDD8wAWaPbh1N9/QgqK
8tZ/atruCSp7jihuSFJGR4J/0svhm+O07S2jyzy8WDcIYXsm4bLslEBWKs7oOsKW
D/wn3RLVzdZRqlq0bzLc5pygYSUC/XT/3/T2Qkf8O3KT+ABuZEaEEqQNsDiks3Vh
mZW2dzStURpBfbTG2/cxKEYn0egrUcbaFCbieOe4Vm4UkGJs1YDduMwhZgbm8OoD
63TiD53nIrE1lDqjc1TahCDJIJCs4s7AabIdKwc1w+SV806RROTx9nhF3OWJSqxn
kVSR0F67R6TIJ58UX8xaWS54L9h7WQhzZF+dKD/LUStit+nJrKY3kmlgaR0JB+0D
FjxwscnwEBz4fz+/QltyDyWFomRIsLRyUwFMcKtiwwnMAflli6eEkIDXBOgNl39B
iaO7KcnOnMf4FyRjgBX9JymNqSWUXb5z2YHSSHsdwrpyYsNYWYfriP+6tb4jVPly
L848mgbL3pdqdQ17HubxD5X5xE5QVsHbeJ4XpkbIl61gAE7geIW4rc0caNE9iEXs
fxxJicasvqpTP9UvyXxd1IeJiSfz4TMqKGuC+SmW/FkN3Il63P+44HnHyphtug8w
RVV6+sTCPl1yx1B9cVQffiWZboA3f+8W+3VE+jsmyeaWhisBxWwf7lLwKbrnz9nY
Bu6dTgWDTXQhFZLN5MRCznWUESdXXd+18Gyaa8ox6GgT4wB3vrTclx3+L10QRPbO
XBon5fludzGpPXkRpNjzjv+2Xuu4mOiqicV6IK5WBdVr2FazNUQB9LGVOOMueK0l
g23EmEwcdl325Zx5Wp351k9RRZARc9mtEnluL/FXLQ0vlGnW6k4E6B/wiqDlR9vH
41ozf0h7c2wIUB2VSL3/WWQUXkFgqiT939Nc7GLT1L7UJROipDjRA/tRCcO0zcRH
FWP1tFntItFDvHlVHBknU1bV4pOGKu9xgVyt/lkZVFKKC4O6mpbORc/6iCbKR1qt
ngrARUXZ3SNxXHaSBlK3zGzD+GGQ74znGuC1dN4rNvHz9WxgdH0ao/fPr0XOwlEU
qsSsqtkUtiKQrDegAzdYj6kAc1VObTh98CEPWDRXMWYBp29gt1ox+q7sDFeP83Q8
Jsuciic8oaIQzEV459zCvLb1Rtj+LuWxGeCvO9q2/fUdBL0vAcgHDbmuNCEt7qhR
kXkfVk++k1WC99PdlmEY3v+ApsWyoMvJaz7QDtMJXxxmi14Y6gQ9a6w5qagt4L/H
4SwigIDhRyBz3JKuyayg97uFvy+KMOHw5NARH5dWZDKHmiNoY7/Ao/ZmjBE5YY9c
2vvGF+610rViV7Gt/ld4LXAcm6Q3F9av6EIiNpy4QYscbkYA3UGDVu2/dpheZc5W
iFz84G615OPcSd0/JEIAEccoyVnOFHDWwBpAASBN3wPaU48T/zx6XTU9UYh/zDqf
jLroXRdQUsU+dtGaUvPOl0G4nkUpRUk/IaSV2YK+m18MSOMALjtFzBOT1MWSCrea
36Yee7XJv1RMwEouToK01v3rVFlZ99HhHSA9jfKT9k7uEG1Fs/z80fgE/qSKxsre
WRyJHLI6TvzjbTfdHMXTr5ddVlPfhzd16MMu8gmN4LyW5COeqUXPJaQnS+9K+R9W
uJXwTZGRUTb/BSH26oTc3+qftGyTb/pHq4CXJYSlGAxkq4o4qQYx5PXisffdkMvv
sxwDKLJBYjUxVcxgULG5bu2fJEIrTJMxLtnqHNWRyfFMIJEAmHvn7ZqZBaMHIios
1Qts40Emu/PGepjd7OgGmHfxHzPk8Y9yI9Bl9DrEGTTsTxntL4Vo1YIBaFsduZJO
hvPp1kVK4BNdkUMWcgdUrlLl3Z7/okEPEijt0z9/2eP3kZW6yAPoQe7z4yVxam35
vANgG5SCZO2rojrOfTDhMmqCxNXWSc2OvTETbbRbsW8sTJ4imK0rrm4Ro8wdWRu4
HhI8ACc5f/l+lpvMfJeHWr1XGtKf3xKubcIrxHdnO8WpUl1CvdYfeAVFlbJB6PrG
F6zmsu4aa7+IkPdcilAGMVaPqKJDTYdELIw780tNyHXQNhdqeQ+vrExMOpGG0ZPw
jDl45Rhk9u99M/DuzLVMXdrb5+wtag1smYQLQjlbOKBp7PbZEzg2AnU9ryEzBTXs
V/qamoFzh66w+r6yHyeiHIqE8Crq4Mad2rcsrcCMV8ESKoq0YYJhzlgFifEtIfry
+t/WjSxYBjuc+ibgp/HtxWKVUQBgiKbuvxBZ6cgm83DHqnzhdJMMxdbAIsCKdXtQ
dU1dZXhoy0g4TsxTFDKU0lrkdnBGmojGHdE3SUhVcVtjU+zVoKQpQqdekdMLQtUM
uKf5OUf0s57dJpZxKQEraHv3k/n6RFym21gh0Qab40c0Oli22XraQ0HMJKN6PTUZ
zVj/elWlXw60EvK5LDk3cNMVv4xmSBTqnGDDPDzRGvpe7B5cm3J7JNHr4fpKtZ9O
CU5h/Zf8YhuaJt3oo5kSXagQGt+OXCuq7w5zfIZncRtGqUoOSwA4oz2GohdsLFV+
P49n6n8A3Mkn16xr7IcmL4q1tW/yjhZ9DfW8WAVzHUzpTLeqmqvGKIls/ENguHpY
AK25DUeiCt38cQ5AYqiRP63DRdoAR+j0PzYBzxnkled6yl1oiZcDI9UayCFu+KrG
HkqngIxbp5b8yXvH1PRlhG/ydUY67kcr/S3afBAwuS0uynmLEUKv91KwXNBnwKnU
Pet/SlaMl/7VylIcsM37Py7xMDoO/iV/t9iDn0jT2fQfxB19k3NUvEl//EnDGAc/
RNB41MOoZuSpFLNAwUAg+8o/+oV/zUeez8OT+nRJcbPLVbTmulD0so+jp/Xsgsif
fZdMoBBhggyWVYDiGVRirXijImj/QM4NwJrSn7sp/oVx5ll0r5io+LDsReY7tP4f
ozJfZ1RHw5rN3JUdG48TUC5kn4Ky0pXF9kTaXvGLDHavgZ3zcBhstZyeBgkp2i7L
TBrDbB++gtGjSYlvDSpHMmEg3S6/x+t+pZBWD6HXS/Nkd+RKvHXfYwGcXse/CDoQ
i8yDjBYRvUZI8OePv/jv4INWocRjVOEtlFeRMoTt2TKtyDu2mnQMqsV7JqnxbACR
dWmOt82/x6GnuiyI4L5M0fIPUA+Waov2MlyoTHR9n30mpoE1T3O8r8uUALVeUJUh
Nc8FMFAVATwiKrGlznK1IG92pMsGQsIZRcoAANy+Vagf112nkh7g1c2r7gxjxwxT
inRMR1OnDSpuX1gabVP8astIhID7LmdogKnpaDuvmUwe6Muu5q3/b0uBMpA/zvlb
+LkvjqMzxW/V94dARxfGCkcNPOLXypWDRONYcr9vu4FCPpGG87PYOfFATDGL7OY0
0jSKodOZPSyY95+lUjvLJuhxSmVzrg9FWLUm6OFUyusMaEgcbfyNsDrqzOFMSSyA
if6JEeBz1Ndion7lua9vbdjTooitTqX/zhhNX0fW3cjL4Yyl6/4a/rDzlYPWLalK
wMmja2iauWiO5JkvmhR8LrVYxO6FiCbUYQA7saRvQNFGLhHecO28fa6itAxJzLo/
OeW0mZML/hpngUM9XWKDR5bWq+54mzquSTA4Kfc8w2LwjWtQzYHU6djKLnZNghLQ
/dWYFpqemJJvOk+P+wvrzu+K9VvFrSIzWFmKmt2BHt5D4EFtMN/+BlBZhg+y3Gd3
cIfvFejAo3RUFtwyZlDgAzJA6tFAFmxZStgwkdJCIixpEUmZ7fk4/bOf+uOtjBrW
TyPPH1Lg4hyQ77IqnxrI+vQ1G+kC7ypTNOxIdXa0AZpmjaIhtWuFRoqxiv6IoBfM
hCvDcbVig7fHA8BSE6FkIj1Ux6U0QU/B3tKLu8PljS3F6aQUhSARQjBIMh5Pfbk1
1djGPrH07dZHnf3+nNatCLQRl0fjbzebHx7KclggrEpXk+w3oN6VJnVGWJT8F+wB
88QsQF7sAl+fjW+Drdvt+xb4ZLahfMT3//EgUfphcJFjvnLK5nq5WBqr85QjpG7u
m+DsYFuWu3uQHP2V0LQYlvWi9BPw3cOP01gYv1fvA2CCRmd4vpmbhm2sWadlAzMS
/7aIm0abo72eAXSgaCGhdJ6ztBkIb+YCv9/hiE6Y/2iaIZozyw4TWnMqZlp9LXGm
Xhg6eCP1gbc7LzPT5SFoFWeYzKGSwCL8x8kkb8Ysyb3CiMIIn2mkN77YZpRXL72l
j4nq/iv45gctqrF4Udr6wPhNl79bVWZDbzhaOS367wyPneHofurw1iTVo4bnsb3+
/DbIECQuTTMsv8fxb9b3pMNUejnJDvIugRqFJiEg9G25e8108yXqgELjli/rT90Y
AqyPJcCvzcaSH8KOCsCRRuimyv3sKGbGEU48C7U0DHTqdvdzy5+vARGAkvSKe1v1
I2/46UcA30XkZDjHdiP1ftq+nE4T31voCJcBirqIgi0XSFlbMkb2fLCJFGA3kBzD
Twis6FMAxvuwWRNpvThbfIRL5PfwCCTbKfgiejBwEjEfbiX7YIKXF/j+oGAuRj/N
I2rFCOQGG4Q7gJbPJRgyYgmtZb3yAJaqkFzU0W845Uym98dQmI34b14pYTQWcWM5
fEnA24CmTMATGyBtKjtzXPT3nbpzU36CE0ZoodNLOWnVvoDZQq4+mjXZWaA/f3pJ
aNURe8CyVXQzxW1SZ+Tbp6sWGg7NHrlB42TKAz4yTMruP+NYSu3s5mYfTF9e/4Kp
Ot9OWF4wy/TUbpA9A/wJqhYLtJj8pr3md8cQSxXltat6En+LW2MwK5WNvllsJuPL
gLu2TH7lufNfunFaOysBcJIEaANITWQ5abl6znhmlzAcJgUAdMpfVvPQR3VxrZ50
VGd986rkr239j5BClaMoHClT4tBteVw/85gAfnn2dhMBVJ5MqGzljtwjrJ+tdxM2
3Cqspe1UhZ4/dIMVz3anjJJaWV3PWBI3cN/cxcYQItPbHkxb737W0tDPwUjWoWUK
u8+lmi442g+9ukr3XrNUMPCPCT+YC4e92YNf+b4/XX8zl3kTocSee8plxZN97lcL
mCn4bWGihbXIAOCWe0wg/LpQOfQk9g+vnEQ2naiYvSmBA2qS5WFIjwRuGFw1i5HD
NoXMfMEzn6QsNCGspa7oK9y9n/g1ebIk11gdqE9MtRMzK7HmSKKyI/aL5yQtA4ds
r9vL8IMJ4+oeXn3x3j0C8uWvfhfvExesL/0Bw6GlWe7zk8Z1I4GuF+ucklPOn0rv
b7EexoD3jPI8wHTmgMbyKMxKh2jsIn7+Jniy7i1GrGmOzXfd1LYuD9hOiB/wKZVi
/O7HLPI8YBlCAZo55ZLT/hUuFt+4SwZLqHmtjG0pdHNGsRwu5CbuTQ9M31jl1lJr
YoyNGABNCebvzDiHwIsANMd+0GJEbXnBhbkQM/R0iM2frq3ZSeF1VHnmEdIO1/o9
dTnO3zzNWePUGkbKHHaY8Jaqa7eVc1PbQulg8V6rnSopD+mU+jjKyikS85cHMCu6
UO5JL+FYQSwqcsNACwBQFdlR194QI7M05FiHXOJoYKdOqbF998ZJqMe1iBKO/X1E
Q6ytWZF0yaLqfWzXwmijKmQeE8/q97Pc495tnQ5Mejh59ZCUOrXpt86DBVq/flYA
/Oxex1GFh/WrIbJ0pqm9UK03Rekw/St943bN4gmOV4q4iNCUZUzK22qd4D226BX5
8MWXK/JemOgVJ9JcS0Jb4CzJzvifOaq+JifHsi2Tjnz5G6cbZ4a8lJ9qob1VQN8s
7vo8L8QKH09cazRMP7vK684xaWKWpnByjWkkkI2eNPOM0W2JMALNTXA9Nydya3K2
761XME27GKYIGDGJLQsa8iZ3pw9eZRNs8LNfnm+atMiC+Pxl8e2FrmMX9HcoTNuP
FjNSR0WfuEFUN5eT8hoJJdvCJnmZmBvnnK4sh98Pf/HTi8dHt1Lxqwz+2COw6bA4
fIFs+gyVHiHmvdnHeKnFZZ6wDY8renqTnuq0wFbvOxpW4TFnGSvCmlth/bLHMlAT
wO/j6MVJ6aDCjH4wW/7xiFV83FdiYkwloE/dgAW+kWjwOxhG9RZFqnDDZt/XPFJC
eGjBT9M9Q+Q9QEXn8GeTIlhbnIdD+EX65HyKJJ6zPukVPHGU/Vo/s3c6FRuzi/4M
joNRguZLWNKGJeF7hMMriCmA6yYfCRYEPBBKCH7zepd80qNxDItLrDV0fMGnT8UJ
04KRvMUBwkNn4jyrGgxcciH2r5qmktvpHlmZxBh/uFU1sx78ueC2iPIpafthxi5/
q6MfcZmxsFTwHmhk0qwAZ2qv3CLH6grg72O6FgHKGmpjNvO+bVCZaCxiDUDAQ8UA
yWw/5rU4P06/7+jmExuflpF6BgQpDRru9f+UJNyv7eHZgMPd061vhOw7twQOTxNY
dlQ72BhjF77miaCLhwbsVg5vl13fib5F/qE3NvhH4WMY1JO27qkJ9PexJpGxHiMw
uekh5/y4jGrjGQeWBQZWd3cJkzTYBwQzAEHN3qdiThtnpSrseaSFunHbj0vOlo7o
Cxm/Fhb95qHcZayaW5sNQv0FJiK6K+zkjfZmjAoCeD9K0rYSoSZ134fRKzW4mTbM
SBh+2E6HGSk+ASvnWaQF5CyrMn/TqgGFDMKo2aG75lIfXH+DMyiVxiA/eKkeg3En
0kbuaehzkCc04xT2r6NWKSN356RxJnk0m22dGrMymk7xZEAC0D3kKSmqADqvbBA2
jTnRD1C0zK87rhEi2ykLySw721OevnvAlRuhrz4OMibK3b3IoOJN00Y+rlyV0KEB
bkZeEbA/LDlz0mcEtDdjDTmiJiJp34sD+nXb4RHPEx33zR3ZKKVBrq2YwNIlJdBu
TYpoxzntWknskSspUizq/3TV4qwGMu5AF0ABjvOeGnbcuObwi+Z31mtUilDYbHfw
qeb1iqWHhh6Qdx/0mWcE0S5TUJF7ZLOhB00Z6jgWhmgHSKZg0siXNEImt4YjDRd/
4xBleIKG9UXcYox+ZMoH0e9xeGIQk5sUkiwhlRjjYb7OQLPC6C789vGI+RrnZGKZ
1W/wXED66zXqOEK8zp1Bivtf4FPUk6s2iiKn19mQbom2SylWcl5doWQgGUm5YlYK
NKKiCRxVEG6X7IoSqU2FLKegbdPcRgjZX9qpdSGHkLomlUQTYT9Hmpzw6FJpR4tR
MiX2YZ1i6B3Bad8v9MCbdmAI8YyhelZCnFJNXLt4q4T5HEffHobt2fITdxMcPK5V
KQXfT46ctdrDdLg4uj6tdiZwghr5W4cH3XkgjaNmSd0EVEhsgSdN8ilFZHZPc24e
cZpXtv1MqJu443sF2wIZ+suB8BK/bbXAsBcm4oMmRFFOU/lQQjHR8LCK3rgXhAzc
SSaSKL8a63fjZdlOFRnK53U7gabv7on+rch+kl6MlH+DJ2zDa4JfSTjObKE/liAf
J4MlJal3iQsUza/pl5ID+sPCtJa+IKgyF6a12WEVl7ktLBMTovhSdkGYcnAQuWQw
pOEgwiLVb8np7Coo3QbqH+iTOXRPrpKQnPeBgfv4pcxIqfKFR7+8+Jpz+nYVZhMG
PsUJswFkctTxWXMwQ+wPL52v+D3cXKMTFPpfqrFpEnT83D5fHClyiz9DQdI8i5eG
DaGCKqxbJZAuHb9+hApjLfo5O4NOZY+q0moPVb6RBK+hcbLU3bhh/OysX4hKw3IZ
L92rBXvmWB2wTAl1PRSI08etd4jF3+Fw7CtU0hLc2dgyi5U5fvWx1S1U+pr8HCpi
SUnmkP5SNRZRNuuq9GOdZcCp2yn2zhNmWoTy05eFl4hD7kYZPlMRBk8qaEghmEiK
cCvkMOkL0LIBfpGzMC0KYZ2AyNSMjEyECmeYxa67NsbHVfHvLiqo0uSgxFk0I1iv
EEQsyZe8wiTlMYPmchGfDt7xhxMh5we9cGJ28mCaWj5xbfgnxDjMQZSYoQEmtVcA
hUpU6gSSfJSx0jgm5IfQu8FlWIDRulhyniquxoqyzNxBE2MK0dj+ylrdzjpqlBWB
8oVrG4k3NmSibJsvDfc+l/f3Zo+wgV5gK0KU3Gn2hKOMfrTAXsXCTn9eGDT6o1pK
7DH2RXGshmhrh6Uo8qxUxWV8bphYVun2arrwmZLRDP/hfKy8RPBpM5xulQ0j7HYN
vN9vfyosFYuS4pjRRBVg61hJtC7gKlhBNa5ey2Q4U5iEi2gDoziRF2O1mWVCMqNS
DnlkefEpARGdL1Jm5W0ychMiRvQBKkh3sKsl8t7F/beMnYBqqw8ykKp3n1lYrRZ8
Z1Bd8844649QgTCGtWtKsgJ3MQ2c1Yx70g0N+drmBeZ1+zITAo8rDKZlgQcCO8vz
4kcbbHF4uffNMJwfpCG2lCIfJXRY7jcEQDEVmnZM77IuYG8fWW9Zq9soEjdudHUD
5CbxsB+GHzmO3nCd900Yma5QZYeqYme184gaRMW+DT0okBORuM1Xt4/HmVn68ouv
rIBXgrihk+5Odvvl/9TM1Ob2+ILP4YsJmzSLSzZH1BKalRqsA5hh6i0Ymna8YAGC
wEXjDT15IEBRKQl5NI8pGrbQeSa/tExXM/y2Q8eoCqo8qmwqZNd++bRFq9p1bK/o
jb0h/123ZNftlHvsdXk0rHyI1Njn8iMzcwXWf0JY/sKlr+xCMRXpqBJeC0I5+ILf
pRb0/rOLlxu3EOfPI6+jw5sjw7niA4sThXzcT8lQ5aPGrh0Pd2tfBwUr7PelPol/
lVmyjlUmClpW9CVjhswkc7Hhh5Po/nk8fJ1j7pOD545jlWL9aidm89Y8Nw0RtnUW
EoeEWw5MeoWCjAT0T0j15OTIz0KW5JqmyXdsgw+KZW8fwqcllGBPU1NVxYOoKdT7
IE4JRk8Jc3X6dOR+OhAfvEQWck00gWkbm8FG4X/9tKFiNX8OYgt6eMFToJAx/ZTF
vYWLrqFWeX0NoXnCD4gD78FrVLJQUnSCv7fmNsC1goR4LcCuPbZo66OEz8uNNz8e
xhHdsIWXD8ri/dUDdqzwzgUQT/O9nBadLpqIe80nH2sYhwUqQmmXMVomw01evrIv
wWUh5K9XgCG3s718AS06lYl3gG7NPRVJr7+17orJM/lX1lgVJD7rtlMFZA1b1SAS
660gwqTC0KZpHPYplEQqI/bYzseRiyFtBYfp/vb8Tdmrn4U9UHRSwM4pirUb5khF
wnE3zhI3FNOU10eeD6szudZVjYU/rQ+sXH318mbCPCdL/YX4kUFELrGzdvdsAc40
OZyVxw/daay56Ta/EyDbBl0cGiYdq83x6owQCvmz66s9APqyUoLMTVudbrMTEYOz
i9iovjuHjl78GqfjmjPFwJAcv496YIeYcvyLkK0aVTZD6Ta1w6FWItOWAJAcQtLC
zMouDNRditBXgLbMt08CrGTkNC5YTBFJfPnfzhOjGWbMyOr+opTa2vnUg9/owVld
jic8Jb+5Uea5kIR6Qys2IpKShpRE/GqfLXm1lwyzTSlGw8MsaA+ct25wxbONfsUy
X2Vv+wp0Vxc/9cos/Bfedvyjb0zGJSz8z1VOLH33BlSC3Hx+OZdQi+JctZGOrOBh
TJESF41K6FKSTmXqljAY1FaXoppvFBqaemgS2f8AN8A3jeVU8U6Z+jP4ldkZOI7L
+VCzN4kcXLFYFmrDK9jOLMavEBAhyDM4AtEszDQpqF8iJHs9YfsY4Tqnu8r+jqXg
qIBBLKlJMGgKuobxOEMhpq2M4aXLsyKo8V+eoZKJT04NvTUvM2ql+kU4IoHTCiB3
qaBKOE3nsX78euEXgCsNgwDWP8isOUev2Sm2jZgFyar/U/dghlysAvJxdC7p4enB
gY/bNGI5NoYiju70FZ1ddgfoonXiUQ9qeGteWa9UlChRKgKF6VZn2Quo1Kae4OGA
AknLeX189vHuJQWC4EkDv6+ZWqjNmvRACKEEffVT9nOkaKlBvQgR5L/WPLYkhwjl
QqxiLwoc6rRIjWNZypLMIVCFf0jBppA0uaYVZHUU4xXkqEBRfT5lKqv4yhLIEMOR
C5W3BOXTJ2sHt4aZimLhDejKKRqaLAqjYavs5lXhW1KeFvNJz/qZQBDLGohEEqj2
L6FaDQnuS0AzjOynvpC6afkN6nyzFHoaGdvxX/DLfR++kwsmT7JOMBhZ621Gzaqd
WeTRlL1kQpF6xU3yJApIg7cR7j74lRwQIv7kzJb3pPHsEg9dr9ZGpkwhvsUSQpaW
UwIMLC6FQyhi9pBl/d2mQ1gfbPOWBwVrTKdzGvhZVt5zjUApB+AUkDNHHwBD4dYw
bz2jcp65YFg056ZJ9PwDQNOUlBmZDEo1bKIhW/HrX4bLVRPtjQjxyREPCSnY+v+2
3yqBRTnI7JvArJBZlxciVVs2MP4vJQr/RKSS+EDq4bgItCDibjpMIWouPU8WA8rl
DKLdP2+juOamaqc5ZRHE1V4Ifepmamnq7HJBl4R7WKNVncegy3RnY2Cn+2idHZNU
s7hSYfT1TNLjgnj7R9si2KNzSHryqdY/WbWJGBKA+5sp7+V2e75Ncxr1IS4F6r2y
2qRyZAZ6hnongLm/1lWyGrwOKeTm+lMxTsV5mrtuqRARfBDnKWo37QR3M5WdKeCH
ocqVke96WPsMQPSlo3NZ01eW4882H4wjX/npPEawIoPWi/WIUUWVPnfkbC7/QNr8
T1woWTrYJWJb9K2UXukNGO+JivTaKXXqPTTe+YYngNAtPIZwmHGeSi31XANfS+SZ
02eWu51xLvf8NkJ9aWhsrV7SiUx3cZ7rYinbcZSf/RwwxEMR5b6gx/dV6szpPVdq
O9s2Y3sJrlzASzdexOmkE4cP40gwZqQnzAUvWBZoxEQDM3xmlguzeHM9Y7NQ0fCK
s9prGospbGpHgZaOLVufnWrMCMRG4ejh3puXQKjA9ZCr8LKFCx1Xla0D+wYif9KE
yNPO+26MFAUKo1UVv8/pbM6mEIAUbUZBOMPqki0u4ctq6S6pYAz05qexdyvNQ+Ur
N9EHjHXpbs5iqYxrGkREIfCMgP+3lOEiSo6pMkGr2BCtynAfZdgI+9kyx5Pz1kgr
8PEIYMvoHT6v8A7mWz9rMp9tqZXDxXsfxq1DKgDzMk9wo23d09/KT9E1s19WLVZe
sDI6W34oEtaL+l09FnZaDFDQgCaT4m1CqC4FDW13Hten0cgmKj6cee1hcJqwr+so
3OjZC8h8LzWnHtKbq7nZUS4w0UfDOXuSYh7WMqkGLBhP0Wp49iodv3/LqJ/mWsQg
OCaglxWnm6Q99L3DhG641Xu3zyKDAm/BpZg0YEJ1Zi6pTFKlujD2EvBFRl5/WoKe
+gJXiCotG/lGwrjAVAwjr9cCaFyQWrTfZJXe0QezpGOzniBnTeoPHKOo65G/PgT0
zaKpCEe4TG+eRr6xdwW3e8SAHkmWR/ooKNk6r8xOyCXnFrLutVt6t+ZM8ngpk8c0
/2bE3IJKgbtidoshXUa86PeSQbe1kUmE1cGeRbVleS2/C5+DI+ZJTrwkuF9EWRMa
GrU1jqxEpTS/lSRtTj/FgVsY+jLnZ1x5TEbf+IIjpCOEdskgNniIrx7ms6Oy0ylc
/fsT2gxdhdFyDh+VNMYtPanXocGuFt5JHO+lphvpxQWAKnixNtb1NGActFAwY9fT
sP6jJbj/L/BHmzBG71UTjRGmqpCTrJ49SnM6FpuHvcs75zo4Ubov1WnI/peJGXYV
FgF0II5nlm5Mv7cBy4cBEFHhJ48CZ6zFSB8uWhxWJmX41YiPYJcdk+Fu1g2+c0cg
miNfq0Z4lQgLFVeekvKfko7ZURXAInWIraGdReQK+etTgJxYwBYVREvFsdSy2D8A
SDHE5JCt/vEB5NeoojJXmeUXbtrq9a0XW5l+fjn/Vm7PFOvGhS8RUd7w7WD8Wg1N
x75oIS1v9uNP/nVmex93Cz5x3CHPG06IOZQ331TJnZLvv7evfYUjR92HuxNBd4yA
6TdEW9szlDBnXJipDJjfCjeIK49mFbQS0833CuInZKG7sEnLK1lUCT4/VFytVkdZ
ngczW3oZ5f05I3a+L/sArIsGgkMoCcBSG+ifr7G9TyKmakpaj2NXBuUkv7YvOhih
eVX+5jysXJ4zXtEpmCGEdyyv8tJb+KVXbuy8rY+03Mh5PtdpFswqsqpS34JaNTwq
+PDmADDIezpa9aCnOTf1O4LOf1ea8Ou/B8nrEExSZ1sVWVMvqlZfQkeTPYF2DZIb
AIfiKNNtmCzsQil2340O6RK9j2+z4J8y0qFHyQJkLYOf6kA0elGULZbz92uVjzyV
vs4VGRSqRfsTCaR43f4WlwlMxtYEzbSzpJj9KlhflNQHIk//ukpKCIgBBL+BXC5T
ZWa24IPFeEH4mMjRhQWIce8fNvHuih58ibuek3iLQOkpR960GJunmpK3fkmjQ63d
KTzXTkJLuofqhrv+xVmmi40HYRTdUItb8sRBMzdpdbXRB43ezdyEw7q3woZXhtIF
BS1FYW4yskG7u0SNhxHtQngqNqK34qPYzZgg59xy+DJKkLjwChztdzYQ0a1QGXr2
Z6hJwTUdGJjk6vuD0ipBoV4rgZbzgNzO7ehNLM/ho+WIx41xqYYqSAUKOrnrniKm
7+jlUH++r4NlV2PrtNDhdCMudgXzOwZido7vMOsNTj5eHsxejOaTbS+eViMy3FU/
EBTdRB6/90qSgux+ZH4EIDsXgeaDxc8NVuBLaESe6aYnJvoKfWWJg2PPfHzkL7Q3
tkHfPB3DSAxI9Vn1XeXPdmhnO7kEX8iWtPvrMpiiaZU0GZvppTmM8sixzsLrQmzH
9Tnv3yykl7O7atul3+9ktYkqRDUL79m4k1JFji23WDdIvSanYAlrA3d+Izy8zpff
1Ww8HPtVO23vHUeR8PgzGiMmLJHD10W9S9na/q9GRVWILK76rhGYclyspPw7cSzG
Xynceic8ZQre35EJxwl+giCJ+zUI2aPI3CUiwZOLqJiX7zzZxhjgmkhCinuHCYHT
pve309cD8igk4z5aUjGVc9IT1Fw6bQC9OUvgbo32EXb4Etqro3xBZL9SjykFJIlP
ATr9jvKSdpsHoP6w7qBedinIFvbqMf5npdpapQ40YazAHxpl0Rcw0KPrtbGAAgos
/zPx2wflEeMcyzSmi8L6svtPQjw0QO7+Y0zTfpnCX0KnmClKrIitWNzpmdouVUPV
Yr8Me0Q5fwJ9W+1QZYwbucHrVSM6IXyrUEPXKl/VEjfJWx+kVT07F2V12l+itha0
VCMIK8n3LrigsT3gOGYMtcCIbKwwZ1p6vkoV/S0H6aLa8s6bUAkUO90GxLirGSr9
XMVLehJkuXyBFP8MUTdlPuG35OsjRSE+W2CvzP9d2Y6F3Y7PMUspvPGJHnufE3WL
WlyxKvhplR2HFgrXsJ0H0d736YWT7ER6M/xyMAbdAa1khQHtd2yydC5x1TspKpOE
EkFjOo/srxpKg+v9NGbyQpxAPr+FHj2aKXzK6vHGT2TT7z1TH8uR3x1tMdh9sy3c
AAaMu5AxrSBjl478gv2y5RRiyYwpsTDCnh2yD69y0YA5Y+DBM6d/ZvsJdhNR2LIs
vQtwWj2zrTs5zKM5aTb+MYASSGiSpYNa4nr+LzfQTCqyypTzcdDkRkrZnVBK3RMB
uE5OU+1BNV09IkUbwVgFo4mdfo8hHGE4unxmH6wTfJYohpECP6QKgaoENYJK4Nwj
zPTFXeWMVMm2vqHGme8TkJpB25x1aDZ8TXZyWXmoiBZnG4bdTbWd+pSS0qJGlQ9e
n09Vb6azWI8zcnK2IKTWW78gcynJ2TC4pSA3FKgvj3vqrpb3hXuNVuQ62dge2HvU
Jb4yV1E4tZpPtFZ/F9WTHWi+lJ8iwpviyZaqwlpRPNuvuuYGeSzdrZ7ruMy+sCu/
lBDJNSDHlkXhU0+C2s5S2x8uY417V9/KOjx8LLs50GZhIxksunXNfW8/ufDzyKBQ
dseqTVMsxQNytZrDb4jjOXB4uYeQELyYHhFVcQ71UPQzcQqzwdz6jny076vADMHI
mxMVfW48VSoHEb0AU/NjFI2cJbTNkytpQn8RPDRpN49InKUkyy0M8rg+MAiTGj+P
2WqtCkZtiziDBqxJkJ8fK/SuMmu/uk1+Bc/WzCjw/WC/6BrQaOUqeyMkrimNjODH
9QJEu3M8pPGnyhurjKRhI2/n0uD2GrukG2Z5+NhLJnei6838/2vrcuRdSiiHVqIy
1SPdaO2pswDonfZ1p2EBFsU30TAqA0uPsPoAEJagBuu9vvKwaOHRNcx794RSVWzK
l8wiNjVJLZ/Bp5EU5QGwyHYrxlWrWua0hLfncujPutloJsxEJ8GZ3blDkfSOMHMc
CSPMVtOSqdFLQY4To7SWhmANerv9Tq6aqPBKj334iLkXMe9dwhM0RfWOkwLyb50Z
k11kY2FPnHF//eP1xl7iopv4HLVJnJPDGSnGZwVlR278BSA9laBkrw/hJU0paKv4
en/Vm3JUb9Fh/Q0jJkT3Q/syKNe2ZNjiBIxf2NsaIz83F00Uple8E0DLkDsRnytv
KLfBM6h68+1pwVxOCFlVokeO0twFxUF26ocBIR7RrOFFo1UtRRXzP0UaBMODSEkS
aGIDAsEG8neKhtqQCF96ndzl7u7JIIjr/8yXXuICgP6Mla7V2I/veZfp7fS1FT8G
F2owEVLpcdLO7eDsf+QkLQR+5jKYnbz+avWhzd7sav7Hys3wllwUdhhF1ITzukry
lQtxANaWnxYyLBgkjQpIjaHlzsjyOCvk71TA2UqycK6SegZpQyPD9nsAt64Oe/EM
g0OYsLS7phdQ3hjf82fzE9gkoHyDIiFv4DiuZgY3B58Mf+ornghUxLTpkwY7oE+r
i/XO5ZjAPrhzdXw3feiUXZf6dZtIv2rGFT+RhQQuxiPp8Xq0fGOjTUbWbgKDXDPl
+TwO89h/5CmaZ3WSA9fQi6bGjtYxHpoW8fG+3YSRjpjF6y9NlfN3nGNvNcco0qa+
3yWlP1haHjJnVV1aYfHd5DVtyrrVZS71lp6n8vjxARA+vVeaBKTFm+F3qoGFJyOG
RP8t/13vAFhBpTF44JrSoUTnJL2dl6gSu1uXAwiyl45cmFnSV48I1+GrjIv5JOEv
taf8H6qO5GMIgnJjEcVD/Fzt2X8dz2IHJrKxDzhk0E45pLUfDsiN01zDVN3oQaob
xm4lMKzNzR/sBojAin+MiNLcC3QCEluEOdrIvc/RBXywpO6GDT+iXf66jjK1CCkW
Y1Q7VJ6mhDg4gqs66DoXNgxXnhN5NyubgU9/dfbbapcSHNlEpeVrlhKWmYBB8u3W
OsdR/t64GfcOXUkMrxiLAk/x5EOCrk86v4Ki9fuKeeGXpYPwJUom4VsR2RxumQUN
Ss0oz1eUIpKsNRz+t1Px+7pR97SvfYg85VSy5jrO2J3NGWDRyWF4DsHYuYuE0aG3
20D7+0nj+4/KwxaWrvJ4/tFoqUVzi9FBJrKIAxDuNOs+cb1x0Yn3f+4+Xbqy4MDi
3VATqr56+aqMLU/p1sgKOJQ0qO67jxjF2XyXzSpyHi+cd/GRvT/yXm5OYvyCSmVL
mp80moxHjk+ar69UdBeMYVAU3wGq8cj6RkCS1xdOmlqr9X79ElW+LfW/K/m84VNO
+L1Jg1lAm5QTYqaMA7fC1DeHKyYAEM0p03E4cF0yeXTG4Nu7W5bzleIxXXZKf034
ei2Ag/wgG3vY+ctqkPRe2IyDpIv1ccCu4ZzWGrY7151u2kXqI9HKnwqzPXlV9QAp
f11MyfvMtWDWePnPcrAkOMoBM/SJmqiNokRfu8B24RJckO125WJsytLYSpnrO2LL
rXpgDiD4dhrAsw1lNP1tnDUJLdPSn0lqulcz5pYBE4XJlMGfup/kuL60VC2tWBWN
o2TiUb5eC+gGnSHtr/QbudEWp8ltUza+o1DOKW6PgEtze0EEXkS6qls9JVilA9Hl
sbX+dZ2N2tzjYIN0iKYvpGL/sMCe5gfxD1PSC5oPagWmGlLMISA7lkG6YN2o+Y0P
P53zpA3JW7ZuOzNoQLk4yT4SSlK+1mMMBsRqIgClSIF/oFJDHEX2knGMpJhN+GFf
GTJyUj8hmZ2K9ytXog4qgs/B0qgkq20+OdjTieY4dMG7bOzU/NJvaI8BKqIcujFT
p6VigSP9BSOZz9dKgcY65M+lK8SDmNOJ2AfFnGCUwZZEZRZ2UEq5zGs7Xuk22QDe
OZpGTEmr680A0cfVTlGuZC2PdZliPJH1LBowQ0K+58dN1g54nYCvUV+g88/VbNAE
lXIPfy69jGwG3zZjKHQ7FDcFVyt1jSsprTvWkhaUe832pAhBdjcf+pr2lqsoasQS
KcS8xaSPdTjqa65Xxs5GOy7dkUzec8FFwohV1yVj4HsjJIRTdjLP3aIFReK7gpQA
ucLaVMfeUnz2AUarEoWje+rF2zXJySpHvDA5joTNmsIr4TjZtRazOGeawmJRO4/T
JpEr7Vs57FWoF0snbHBjq676aCd/BnfHCPEOOHCCmW9x7bFJ2jL+XS/MkVI3LtCD
MSEgO1cYLw3kf+dkY3fcoeb7x5uV2HVR9J6CsMburn+GUUu8z+w9YXkYad22CLLQ
5T1Ao6lcvqQnQRTXg7nrmBF9yoMZZxcxIL0L12YI/FenNVOeLW1JTgyKL8DDVwNS
qxenZOjQTHe/otfWlCezjx8zuaW9rsedi3Yh3wNfNc7RV+HQdb/k8ZxLdR0v1YEU
gF12xci7qWrq/L0N8bs7MfA0lL0KIy7Btj8Y9HTjU0eUAK+QYQB0lSXs+JQGNLaW
S08ZOA4+rcOdgvdr32VFYB2bpS6fr8QnP+TdHxqmbtlHjXbrRjtwalIPU6Ycx77y
wjpNe21jRMLNEt5Ey2S7ijTbeHyDJqOvYMFYMOphX/RnFZx1lY+YUzlAttDZbqFA
bEjlVYU6gyDEi4eOmNpM9axRzUg+dVQcFjMp/ImW7LSjQpwP79c51VuQu3sQ0G0Z
D7CBN3NcnSRtWP9aQi6mYt+JhrwGUYsWfB1JLFe8pzHfGHbS1O+awrTgIhKsMnRP
UCLyI5wBwW921LDYwaqMngCxx+WJk8CEn2TTsinXSLF/SAEWIpWxlzA4xHxurmzn
8YYEyvs6oSvYnoorJUaebZIWEWFDv8wef6vBEMDlctSNEh1mMFKa8RDs7CqpZIfr
8W+MMGop7iWPLAHQfa2BpbVm8aXXmgXXjXy+zD3/4qatw52dHEAv6+U+cZKlj/x0
VmyCe72il2C7Uv2qYK5GBD3ZB2x9yiUeN/TgdRMSm6+yYErKw2wnm3ves7Z+IfSa
4xa7Z9YrsUfmq/Mi7pX5krMg537Sy8vhDlkUY+0VrYh+zN+QVO0+JaDgE/NjdG5N
PY47NjTBAN6tNChsjC6uhgw9+6ToqxXJB9XlcG3GuY1sk9ZRf76YtedsheFbXQo9
66Ff4Q3yjHboMpTTKLaZl4H6MLHfH8HQjkhbz1Na355YxIJmmSu/H84IzGBEDSK4
OG0Sxk4lTJWnrxLN7PRusF9m8oxFg8lGtCi43flMP5DChKUgFn4F1q5veKo2Kukp
LUoJsDnH3nGNags3aHzGAEFGsK+2Kr/HddX3bTJPA8vYhOI3uY6pumN+sMRIGwj7
yzd/Bjhgl9qxk+1pIKCYEJDht1yUfBFT9B22RZG/2xNy9i4bUvZmy5ZP2uDHKVu2
AOLqliD1UzKsHLb3ph74KGJQprY2m9hVyx8o/ADJZe366/lBomJRuS/XSLDX2PrG
O27tuQV7gd0n/L2WrNy9N0A5atSv2wE1MTxWmvlsompb8s4E4PvbkFfCwP1lvcBp
pkoGYycci6hkD1Jd3DdcjqMDMSZAZ6GpgvqbHX9Tw/SmMo6Mh7ZcQq4qQy9cdmNJ
yvLDTTFIjSh3Gec23ZG2wC3WaefQUNLlp9s0KgRRVq/9KGh2ZFxGfjMMbxdKmSjn
FJFn0CG/Lx0/b720i4HGIFKg8l2VQ1j9tx9rdVVz++YQj5jjP0GDBF6bQDHs4scT
cuPH00c+PSd2gcK6rSvhDeHB1pwiMzhrbDP469uUemmdiKPbeYiLcp59/ktAwMoK
L+bL/myi8dcLdM71FGbA0KtcQUWNSQqWtKMd4gS66KVKESOj20SxAXUUULIVHYZF
yAOE6TRQr8Yxf2PedZrLeudOJvzXzCazpO6W4N3C0eFPM9NZTyDfHFH3z1g4VxyR
E9c4JAS3qsS365mUrgX0NFbvr4EVW2pHk7wcSzkSoOk7Fc3RsTxS93Dw3i3AQ+EW
TXgzpThLPfMHX4RMGJ2p7yj4/iJ1jos2Sxy3TUe5AJUkVNv5qvL0M7XcrcjZmDmA
oqftjTLwoz6z+ZEAuwjPQ6hk1U8Bf4FyHp2O2X28wvcbGFLi/uCeIepjKo2qR6NA
u0tgMy87lNwVeUiFT5XSsqdDlzdZQ/iBxo+5avqSnh7YeoRTUsuABxkkxPF2YFVe
ARcuoUrr4NVbqigtrsYk8Ahz9MNcMy90sdxiB+g/w3PZ+TxXMuihfb8z4PLs37v9
r320b2uOFs0AsLOuDWFvb+Hqlg+wyLkduasHyajFO7/LToTG6w+GUsI/s/uXZ8Zm
0YbbMXUsQDUHAQyIeL4LM4GAagqrlNSBZOB3xb9zdYlBC+LMQGtMiNsMGF5b7BXu
ILYq3BTdCv8fWOASBvyzGqQBws9m6RGAaQgsY0wcwZoFjsNcUidpEccY0AwwE8Ua
AdUWhvUYA1cHVzZWL22cb5nqEZtvP6sNKjUxXHhJP0AkmkjwGuFozg0irhLsq37q
+cmJTlzif7zsnTjDITYzXi43Il3kg1nOAotAMjx2FsQB/CxVkuk0liN/BxtW+qbk
E+c2k19ixBkT3ROTT3eABpLjbbrm9SOfp61i5+ps5A3NHH4mWPbTLg3/jWxNNLew
emHSsrA3wtAKbWkxM/UBzXOf7zSKuD5Shq8X6p0kjXyZZe7K3CPYjqtOp+V2pwUv
X9QASTT7Zf3VZk/bYsXTssHsSbgEqt3sE0L0VElgXqR+5Ct+h1yKUPdna52taACs
JSTcRdG2dtdu+LyXtpRl490mERygbyPUPb0HwrU2rvJWR5P4dj/uqwJXh5kE2Fu+
gesdi90MCeJrkzl/mF3KY/Ez65jmZHfnQWjXMlJwi+euCyKanhykfwFYS0bmXFJy
/uLxcH2v/jT/HoMYg2ZbGVu40dpIAzN4T1vD4jVBYCvvOLAjIjpqnvs4FdsIkPZ+
Mo0Pp6dKNMV+6tMYqs/Sw5/6BeLUzBoFrkq99plCRHy3aN5JB1w9VLMl2VO6inrO
HVvcMR94nSTShiLJaPCH81DVi2n5qEQsuVVfli+FKKQUbr0SKJntDSB/DCKlKbGa
nMnWCTb5aMrvm+3JbRVxS04AM0vk+nTq2wAPRwhDoJ2XIj8gkbP31aWbp15n0q3+
2f144Mf4n14P1m45k87FkYWI+639/K/kBZR3hjKYP/HA7To8NRuVSjx+dd1/+LtU
UeSaZpT5hGIW4hiabTBIJ0AOvvyM0HlH+G/fZg8X/RLD+cSODGQpBgPPYjqT+zRi
vVcf1TBZjOk8V8Ni0YpQ9tpahUQZwkPBTrzxXIfXXEPkCoS8TaM+Wo/wAumbcJY5
/NfEEBdmtZfKit7ijNM4NZYfw2u+5nPOWf1EXy6YCad48irLlI2ACBa6wwXXW8dw
ZOSj6RoJ2JsTeyd4oryablSShjmbqxNC1ImBh1rVIcm62hJHq++qtWb18MXypUuC
/DK43oNNwayU31+L2+qbIQURu3hmk0vbFJcqiHnLvsJUvrgvL/F6TE7JhSe1N0qv
Y80Ky5ALdvAbc0rHHfcJCxpZnY9HNB87sMPWtrL7fSSBrwHgWGwzQ4EKoJo8poGc
XO9Dp9z1rJPi+7PbHakaUZ+OEt7LJPwgjt+t18fVpnu+AF/g697/7/XNCChTsblI
ZM22AW6+Io7MbHT5d+lyJtPFBu8LZbFEVJrF7UgTotqbF7we4Ku5HyDakSMuX95N
o6dYkDk08KpJb9AaCog8Kus0pGXRwdJHaD6AZVEJf8/2O9W0fDzsRV0mV31PWTit
GKmBvqzcqzDYdffAT+04N0ovIyPzyR9tBomH3xgbirzg46Eo5bxaBG/qDsdDck17
5Eknza0Jbj35y02NXk9mj3QupGf1nHcj4PfNY2dTHI6Yjl7cZCacmhakFTiIGMRQ
JgSru27O2jEcmwnQ9HbunLVWhyw2RtPND7lMxf4efAFJX79orT2ciEYwsEcnth+7
wK1dQS86wr06DIYTiOo/sBjnCpAPXMPWGYUrjtTRoaQG5D5Yc9PzBKTDk5lpQQXa
QOwNPG4lqqKsXqiixX2mfqA1R2RtPtIBxFJK1yGbAVjW+RzrxxqoHf1E1JUC95Fw
8tjrLAdkfs6bxHqQDaBjhKOHGwzG2eQPDs0x3Bn1t8hMg5XOeT7qjg4NXJqcp8mI
iFObUwkhc7R46hzsshiOZCwxqy2nNifIHHQbNoQKiHM65w4yt2WK5u8P17jPNMQv
HB1G7qcT2TUYQoz1Ww4RBrhANUzoqI7PO1dLJ/fahXOfDOmKKliL/dUqUCyQ1a1X
9q7oS+281P6kwv+dRGHXFgiZhSHAytaH9s6kvfIw7R8N6G//8eDIxAq0ngYszTKT
c8ksB27ldD5hQPBlnFhj8RiDbVmacjWCBFN68WVMq/ASsG+ck3R/mSOleFUj7j75
kxNZfOqQnrUtckMfdsImVHTVM5qyVOkJ09vklKS7QeYIydVcFAvKJ3k/tUBif6Wt
i4alZ7s5wJ54qFQ2y9zP9YIDie6TqhMmZc2XrRrtZnMp0y3GKEkmSXYs0D9ScooR
Wo9pNLB1mzqSplXM8rAyf8+KrVw61H/EbLvYqR2f+IIQcTBeySNZovtX64U9eimm
+JtO2ozNnMa7V/DNsZpNQRRDLQHR7OBg7mM6RFNwYFmKc8clLDM3Ox7z2AeBpZLI
Ij9IOP26ZCks8jkWL+TEdFJ8sadi5+OE15V1BOYg9XSs2aEELRwqoNSa42IQoPJj
XoRE4MKgWbZRQkKkjmT8DSO1Fe9dMYcCEGzTjvpx2ozeKx0097n8ohBDcO8tNkLI
jgQRjqc6yCHxhuVEiuKdWcSdu4NszmG1yfR/rc0ZvWJnkWYsuFJSz3c2pNVl/14o
qS1cf+NTYKTsadU8cbgd4j65m+ALmrBOmZ9hEaJpG4kQ+FIte502c+rLtEIibJlb
AFZEAaht9ovVV2A01R1/URy5FApDcoKVKiWw/HP0cayfDZyscVO9rqQPtvP8xDst
b6Fxg8WWLw2MHVXw7KZR+ZZ+lS3bKC9lTkHIFvgjitoPPQxfT9THQw18DwGyef8Z
zfIXGu2QEnYRqe2ZTfNytnCI8pc+GEufLzHPdRKm4IBw5H9qjD3fZEOhqFhuDFoJ
FzNnDmDRpsuxToGS8HN5AShsww6nUHlb0KsN4XvODF4APMpVmn6dHgHIj9qRrlFx
CA0pku/VoJTUoxzbj1QxR9hLh5p5v/xH6LIVZhrTE4pSJCN2mr3vLhPw1Xx/xYFR
vHnikvZdYAW6r1KzYQ6VXv3alyRHbonYZh1CYSI3rjkJacXGyibef5BZxOnfZ/07
qq0IkZ6pkIyCdbp+ezhZ3OrurhzkZ6pJss9CBRhh6Ilj+OpBLk1Wcg5adVjo9euq
suNK1M8Z1+ls8nRqfdgr7OEKjGvi6xh3hOGpzsmN6VhIAoipO9H1rA2hxs0xlVC7
DhBVszY/Wt9pDluF0Uh7NVfRGh6TvVAk7EjzeeSuVRMbYlPHABNWcVaZKaPJ2PdV
MgA3SwhAak765clXgptku+amVj4MejmR33Pbfwtw+8u0LZ93hZx+dWZvHjIAqVjp
0QCGdQtZt1d5918PAfVVuCBPW2zQoTsSdtsaRiHz61O0Iek9iv2DIhOkmiTs/taQ
Qb3lANkKEL/X6IQfoZ9KgelWJ7A/IEHcz5nA5iZNvDbibDsP6qlTaSmxsfbxTtp6
FI0H3QO8eO4Pv5S+TafZj+5vz5zpSE/EVhkXB3N1Wd6PLhnu8pPs1VHavgqaGRfY
fKXStrpoyZ787BbDue9uA9tayImoVof7oVvEDIp55DCcfQquqpZmZ6fNDsoK4FTo
CrDHHJ4LvWjuk4tKwLsbcj0kfCLQNrnz2q+hsrOVLYFZmxBdkerpRY+P2TvibElq
Ufine9Dsrf7lRwo5GgLvw9OHp6+0j7RBR5k3fedQPz4+j8MHUWaowfIfGg3rMqu2
b5mBCiDjkw6lQigY+5vqIgikvxS0x6sfR8j302Y7mS5V569L8M2tD87CKhd8o/gn
Qe+yBaXldtcOUc9ke0ybnjEHMtg0GanQl0zyZA62eZjYiJBcbiQTTqIWBX5RwLOu
QGqzUBSV+qV9i7E88R5bZFdDHx1KM7VJoBVeA2yvRoJVEOiGbmYBN8uQwhtrszcr
juoG9R7BQFh4+EUf3bxTXEXFhU74r3Iz1UvMIN5htHfD0JRrMGzO5jg5tYb+DtTU
8hEBuoL4kzdBui9QRJqPX4zbAMqhapS6viJeljf86RdbTj1ACnS7dWfeqEa3v6yj
EjPqpFgfUc0ngwwkbzccldHGG7SfRFeaxfP+g5403aKS/a3tC2QJ9rOq2d3cMgr2
51R1dzGmQJe7dxk+w3SnrfumHfEwAfbTq/oVHE6FjiGNS1KXUitNkTLvuNjIh5F1
F9k+vQQmwnYeutNPdTkZFxCFBSPG9Zad/05NTHw/jBnVT/kKz1rW3YWN2xPBjGnd
1vxyP3yxWGYsVz30hdzjjSU6svvQ6cdLV8TQBw0TeyzKcey/gdw/QoTaux8zOejf
K8/ERZ6nNIHgZSGMyRNRo2vw0EdVYAM1/fL6NSnHyfbQ6uVgYNhbTKZdbz2n7KuT
gGWdn/+o8PZil7I0Nhw/43xi6uERZ2rT0cZ641aATXO10MGwEtPjw1NR+UfGkfSC
NXRvaU8bE8gP+CNEP0N9YNig+GM8JwyXibBL9c2AY7chDNL3jKzXjOdCXr1u0XKI
TQb5tD8QWyupVM/1zjHRXWuulnxnLLOeJCUblSjKCNBBXIh3lRk4+1dgDyitEMhq
wKaPXtoHDpS4wSYAA+fSi/1TD/FwNbw1YoG8rbs8gEq2CaoEp57LLR1I4JWmzjHw
oxe2joN2KMzE7dsQy+4TOgpcDGDbi+i+EQdz11Wb4pGy0SN/r+VBwC/SSRHQ6i+g
r5Sn9UQhudjFX/Pg4iWLnohkW4IC2671vSav81bsZ16wvn7LUVyf/LJ/ICwv481C
3gw80DvoauqpwjOrjPfcm7I8xuu4QlxlaQbTRn4aoijYYxksuI+r0RG1EyIztY66
cAxHfeEWxFamHT4agTNDqU0KWQXX4+x7tfGCkfuqVYF5NLhRNb+O6xj9Rtc+SAoW
QvPG7gHCJFVbeeIopxMjDmlpoJRmWPSdJSaUsILHrbzRKtEdEB4H0B0QdnC4aGfi
sV3lc6HWo0b3goN3pCN/DkELnNTqqq5MDzM46CcaIOHRgSSqZpeO4FDI8efX89yg
lACHJJFiw6cMfhxCbyTdgA1vdMA2GIHH3W62D5WZUMJicTQSixerfaD0W0WJDPbG
pc3f/w5yKokytPi4bf4rLZ2N7asXhqM367KgM/uGp27zAp2CevduWzF92GT6u9pG
QJ/vezNUEEPOkcgZzSQ85Rkj0nlMCQszogZS1C4ZH+PHUk1mGKcfRHtK7fXShfU7
E2lIfyevUjT5LmG7NwSKRFOqiwKsLdwPDoK2FFJJzGneU1xAYkXiZeBN+uAtpmMg
TQ/Kjlwm3QLTCDWIAz/afcvsKv5GRrNEfUde6jceRmuLasuBeYgZLWtKUO+lWhdo
ZE6/jRysvnBus3FZLBf514t+rD+2ZDu3XNugygNoiEG7QywLWHHeBgfh27YM/JhE
lBgaWn8sG6fKKXGsSCwnAboN3Hyln0JkGdpVNyEFqKYLVKLHe+OMITln9uqDNgE9
Myi+FsUQlUGrei/xAhWiRB5z3OeU8IpPEjQudcBiks0AriqBAnXtUi4FA6QtsGU5
5UV6bpVLW2EHWlT9D/PXXb+rxWomIshSQ6XfLVeKeNSo+la7FQk/C6MbAE4JIKfA
hbnNGKb+ltbJmU3cuc9KmrPa2x20/CeCU4smHWbFXLTaSu50+OQAHHxtqeoumfoS
Jvt2KooKJsuniY2MkkgCub/48Bj5CTGGPCF8srrrCO4uYWXBDkpL9/cIkGgrihsR
oOCC1pv0tCy0S00kla3slIvGsFfORIgTAzXZm8niK1Qp0Z/HHl61FZIvwraVYB6v
un3LijeDVlfE00B922bXO9n5zUxeIbl51CcA4B8WU41zz3e+kRIbGEyUmXpszYNC
dljv15YCVhcQMtQB11TMllNnrX+rtTkPVLs12u04pQFvib4v7SGXOyvWnEtvs3jv
pdCcUi2u/jqyFJW76fwcvkdQkFvDUlL1af7oJa3zi7aYeUF4OViXp8dN3MSJQB5d
NRQAME1NskiV1Zzdb5snnkp5lHfRmJdiUROfSkq5vDS3zOdv8ZuZjkSkckhEfBmA
LyCPI6KWPoeJA1fF0ikzdtkKmYSdjIw87uI4ZJ5xdB5yERoQe+3XG4E0RcosQ5df
qQyEbGlxHvyGjoXuEx07ikRBwQ4TKrjbbbJzl8ln0dB5RJlS3660OKKwVJB7FV7b
17aWKD6qDsdKZkSaqQ+wlhwBWt1WBUceW82C0C5b/5ehrKwXgpq4O6obSI/3c2IX
hEtg2uVT4U+ZTpsFXnWRfEpypqyHrYY52ZXkAuChXUu5hxKaLuOtADIl5+rxY1Zo
laMjucr/AWTeQ9h6KmHdHr9eJ4mwhX7qnvy+pJTeZgjTZJ+XUTDX4veBme/IzLLZ
mEgovf7r2gf2A9kLRV1y+TPy6nMkieUAB5gHHMKNhajzDhDAWj3doIxKwljTbDrf
y91w8w4iUdacqbEmnmXENYKXckzySf/qOmMeB2SNU/yZBme+wwen6zZAhmo4pfHv
Egjhi3deeGTu8wqFJS7ojRIQ41CPts3IjDYzTQEq8auhHNQyD9+oqgox6DVs+xZv
lQN1xeNCXamD6Sm59OEv9GP3hO1sVTP2QEgBUiTB/u8vEdYaZh7/ewtt+8bGo6hd
Rr4usJRwbNao/NqDWMRkDxFRn0maWJ/xgvEUyAyqK9N2hvM4jMdeqsHvIpq7mzjj
trd6dJvIzffdPJHMCOQ63wjN8g8cD9ay/UVxFO97GEnlzYQ/585j4mDzlUZd2yfC
Xr6ovYp4HX71j2JzvNObmIB0YP/MHgpwZWvKxR7AatjLJlRgYPlYAcIG4Aqpfqt5
qX/O0smZXBZyxYqwlB4P8f8gr3NYznA7Cdg3koFHPhfb1Q/OEP3gA9GTT1uIiV33
PRa3esUA5zMSfMgF3aBzJPxoaALcCZEVsPMbbGOZRUVY1STLBHpo9zLOY1LgPiRE
xdATTGVlAPVjxOCCGOlrrX7IsoHBrwbfofqkV9diRBVKMkBNqTNRXmv5nkuy+sno
QSqdW1Xjlzj9PTbCfUA9HnmdIBuy3HQlOgHdRQ+NxZ3ghQJpGYR1/pMFb+KZM0HN
XLhqxVm7VC+Cu6NHuRKOj2nAe4w15+Cz/IWbxmxMC6/ZZN2+EB7a9KcBIIyaImGn
cI01Fqqd4BNgS1IjcFrDXM1sQzuW+ztY0WLeYFGPcOGdVF9ejglbm5wsOGZLeTY4
vIF9oEm0YdE4mcRl18EPRzlqRXeh/7KH0uH4LPB97gUK9Fk3MmX9aA1LukHnkdky
zdSj4rNIpTsu1CUgnXEdL+mJt/+XN0EwpCoi9R1+0JjklkoQ27j8wIXaRYnJT6ew
AqmMw6n1W2QWlEtFoXv7/ZZpP77mSuusnlis8J9KT9eLuSOan+mT6GgO3HuOo/SC
c09GhoZDEjMtzs8QeClQqMoHI80pDygf8upFRmvllUeSkKDbo/58XxdDDfWRIPOV
ksZEJYem5bNZSJfx4nShMStgPJ9OzbNG8i/U7g8bMT1ASW5ib4FQz+5liRuIs/Wb
/Lw3HwYO3YUoKbyOSnyAE4cIRUBvLd28RBILsHf+9Nk5TJX00hW+ABbTUMHg23VP
75Zg9KwB3B9OF0S3vktVe2gGmyXirkzzt0YI5kmL2DyJ11S9bCbGl7TzIye15Kw+
sTksQZU9F6q6iZiV2i3413Ql5mkqrSxoxfgMqj2d16tgutQQnRAyWth7+f7LkW9S
GIX3VqTqofAKlmFzm0VYg0SunAcwWEN4LZenFlMhfHbbsjNdK/0sxkQswqsn0EcR
ciPIT7XwRrDZX7vCogfbC0siwF+2lM7JzFt5SypaoQAyEaWOTo3aDzt5RzQQjjnx
sve5YgDWEWgv8iSPBYXfyAu9SvCC5Issk6ayAI+Ctwy7Fom+jSFXHW9e6B+j3rW5
LGClpVDcQ4N53kTKnqih27C+4PuzFWFotMiO+ifZhqjgdEHfYtAvf7yQHMpT3nQd
vZV0lipNcv6E5tADd63vxdcfWZC97HH7fEBtxN+rOMxW8bnEFtCVhPhUfYKxOA47
KphnKSqqE14fy2ArPQD2oTDO+u8jXULmIPfImtpCOQdWsdASieeFSJjBh+km8KJD
PgwtzLGgfPEK6hh5wndk59lf/hI+1IGeVuiLUOTGhnFc98ipLXjIyEu5yuZ6sNV+
dGkbwyD3Bt2hamZaIJptM12pdd9ncoy1RYIO14uw71sqMf41nbUSK5yH5KfaFNSy
+KO1+lB4PPXO8zQON/He2Op/ILaQntng+LF/jn+Q4NxIVXH52eIH3TkmIiH2LYCf
VIz6Du/McR86DX0rEzxSCXCtszlV/9/mPDQMynN78hHdt3Of0OEzeXujiHyrLO88
bND+tyA3/Y6U19XnCrgx8qEIl7yRjxnNvU767eTjR+pZfUEdWhNFB+y4mOhH8UyB
qduYwQrtvJR7FjMS7+dLVGbZaoDtz/jMBnJCZFXp2Sdfky1pa5mon4guxuGuoR9G
f+lPG16ndX6ysm453mhS1CPcuwwhXkjVnWodOmDrpTnlotyfyGnu61lEPq8mZ8em
IT3NJuS7/AFm50ERjHv+778vLuvjg0z+aTH26wfAXpWbwlaPdprXZPu9/JEP2ECC
S5VEgSd7G9lMEUZHbM1CumvdE6rOLFsx5DFiG6Rv4rnVuKneN1ch/cMy4Hjh8REj
m5bi1CjUfCT3GCGVeRRJ74TZ/0jARwpH85ShjY88jwW7lwI+lr4E9zksUbEB6u0M
yDJH7qIEjVj17SlMqrg3rcRo0i0iWjW2jBouF3IvJdi7WfdklbmA81IE/ul0m5B7
edIcOI/as1bsy2907t+anfRsydOzKaxxFUGsCILzJD+ecZiNK7Bmyy1AFUaBR4Lg
EmJ0ptdwvgm9I++idlSiJIjJZTU03tjuHPjg8b1gwcd3fV5RgBLdniONsiZxW7ot
kMdBKV6duauVXn+yAEHwWpMOVwSb9ldMebsGoF9v/xWzuZ1nvY12pAPioATdHIvz
n20mp9sJF1Ec6P1wAgQNRC9DLxFQt2xlOH/OuNxXcTAxVnOlaDmiW4zrGjJh5IAU
nkr3IN8DtLpnAuV0j0we4EtZLcI/siUcDS0fRQ+0tFm+YU9WRuAXqlqH4zTAMVzr
+lCnRc650ucDt2Hs7O8/iGzdF6Q5pUeu2ZI6AjemqKsLh3dq0KE+l6k5Fzp68AZc
L20M5Kpuhvjj0tfVNjQFq1Rigf3xoyD8DRFSbBQJg+VpV/aW2jAOyS+1TGLHYVFN
X8ouqH6jgQbXJytqUD1Lxc/hcMF7yvMxq7/KBM95MJ2PQ6F0XLm5+62bvpp1qtuk
CP4Y8WY9p8pGM3d06NUdQ12EfRLwgfeFf/F+43zFyLmrOQ0zx9TZUnjAOwrLLvBw
4AZOHKZ7cl/d3ldHQQc+5VTT0UNzo+vKo+Ngxbjw+GWfOGSSQWYW61eIfeoBgh1U
yVpzs9LEuendpLJSnX7g7dpCUH4A3TXTpxJykad+9RKx57C+Imut/Yc1AZcm71++
mgJb1tKRopwJlfBuPY9F2xYH2+7vr+zv2xhgMOvPl6gs1pexm725SL5UZ3fdZ5Ax
pVqyQ1wm5LXFtW+oDyqAt8/dYtJUh4qTLYjXNPgpUjN//cE4w0Y4nCXmCv5+RQKX
Y1/uLfO42JBlvG+pIDnNzwYW7cvmTp+0Jx/WHU1ePLeUe0vXnlIeNexrZbWA9XAF
Z1fSbWNzP08bQRZzD9+ZMDgg/jInek8ACAF2dSINi+LEiaY0qHTI0pI/6ddeTGKe
J5FPRH0MnCiC2e6YLq+bOHyWiyVTq2QaMsTauzzoPzY9Y1jocwIubXRyCdxxF4Ax
u2iZg2i+19GMwuEtggYZZoEIDYiP3/M8z1YVQq8xCJMllpxzA/KcuG+TtXRZplgu
JpXHRXJFzKS+jDlgqIV8mGyRhc5Bixs1kjJxHLzfgy/ihSZgjNFObPs4JkMBvtTV
BAGmjYxt5q0liLqpaMaqpSaroNIJcbx1hqQp83syGoXDGdkpTsm5Ypk7FChTkqz4
FtpCWfT2KRCrdquzN3PtrtfrSOcfwnOZoi77X59E9+fS0X3pgifdZ+W4tvodxw7B
1RmJqm4UsKFC6C1FoEuUfm4u+ZaAl4tPmyusZpUoihTig6PnMh4cfYj7TzqWSP3/
YpKbdVb92n5K8DRUyGVqhZXNI9dZ6brZ5wnRncDE7xX/M/KKd1TVtdDdDFdGCVwK
RO2WvvC25i+8SFs/w/eM/bK/ts0i+OgZpEZXddph3O9gxiKbGPCRhcx89eTZ91aH
nUKaIz2CuWFrd7dStH02LIAR7nup40czhxo40uZmY203T3Ke1aywIPYgsxYijTk+
C6tGc4QefxcJZfLtWYU2cRyb0ky2cVqH+ByAV2Yj6ZA9wK8lOUN8v/oGW1Xl4t4g
Wa2RFg63BuBFkFiD5g3hsy3iBCtS3w90YWQBi1UCZ8dUTJG3m8uFpxzBPLJdtaTB
lhGueTgC+6o6Om/6n9NJ92nIw9jM79izXeTjnnG6NaJlJvHMZ5V0BdTVdhWa5Qa8
yEOcMBHhzogl+/AZXtHJwDVd8GOHTfASC1tJ8NPXUG/Ooy5IPHYghaJYVGOQinsz
nrcedE9xP53R7duOd6HfzbWI0LBxscazWJXSlhQnh7LzAUYVdDXbr5hK5cKXIxCl
s4RX0wRkQ9Rft2lGIlZucZ1MeJwGRF6+50gOPGQy+RgZHchXkX7HucPmPWO0BK+b
QXnwOYJaFURCGgT3GfFF5smhLJtbNbC1GkHju0k+hIfPlc3Q7VSZ70XeaaKfxAnj
WWw1zdXRg/SAaihl7V9z3HEA4x55kNaYbIE9TAILTdVCXMhdGNnuRy0n5evkXrHf
4ykvqFreLkozfPPBiOQdC1C5jLqz0MR4ADObsY+4/9nZlFQSxgEIIuc4N/r5nJ56
KNBxy7fvIxvjAgvEBmPpHxSuKLY8lsje2HXNzV43ThuZ82G3lyHaHu9BCbDs+xrE
9BWa9k6ht9+oGpheEcFIAdkEy9PyaL7as/91VfD6vrt5PGtUbZn4QvZFZlKE2J8N
fJLks0PPHdL7g9i0wvXuIwdynIvCS1YDptSU9axMUMlVw/MVlEQ+SesO0F+alfuI
g33AglGsOT95vHBAr0fFJwY+wGIm8RbQMeB6YIw0QDfyO2lapW/3yGBjxvFskET6
IAfa8zLAVQW8BzUC2zC3EJZGtdMzNIV5Zyg2Zu5vq/Y8lsenZawJa/s5/r+X5Tuc
WNAYK8zyB2R8KW48xdH+UZrfxmnJ7zGmIEetccbdUVuVRkfAU7Y8Ak1PnkbXdeT3
5TsqfAA8Zarb2n0/gXcQceAIh0TmWgYwu8jXx8/Ahm3fcO9YIzxZ123En49mqkNx
xA+GyVwONGmfXPjt0vbV4+jLFjeBHHG6L3Ohy/bYpvJHsNAxJqZY8zBXhw6gUPWg
Iue5kob3k7U57rGKLd3LLLp0TEhUL+dzaiwhDg6T2sKuqUi4LBO0MXvwm7eq/A1l
YifMArrtR10yAQe3vj3Wwa6d+EjlIkOJQgws/opmnNRBlv7QZio/wdlU7lMR1ph6
6QuIbtTah7RVnHUEuHvnmNdUDemHb4MtqXPAQrAD+blIP/Hs8YEx4cJqeWwBxBXX
gh00m+YNb9f0r70DblC5E+qiAZExNNvAX3CK0lpRO0KP7gtmtfU1iJAeeJ5DHRSF
6FiPjp4bJV4iFdUAKR8uMOC6oTnlROOJ6BnoSmhYaykSP/otrCKHUh28ITtwJW/P
A3nXyDKITKY1M14BuHe52oCzIZ6pEoKcGkNMtX/YJDYXDgCTzMwyHeRmyKCq8qsl
cjrzHhoos/CrSs3fAkIjZgdSXRvceOSjwKHcqPhgvZGvt0SYBPs7aAH9bDXmh70y
7nuMdzyD37WAFnNdFx3LIlS7miSxNWdJ2CCI/gu4ZLVauM77oW7fp9qmZbV86iD6
rrKpQd5czRI5gNNZQbmWzJpdl+J8jSGu/ne2VcErQZl5irm5eNH4/4+ajLs5QqKs
/TkArrQT/JiZeJdWouK7O+WUiWPlgsVf0F8H9oAhxZWlNBPISpl0xR7mevS+BvnZ
QnFfwk2U9nSEirKi2WfqixYzokKZ55A140x1KVl8rBr37CVt+VYC34LIPmuU0hy1
JdLiyWzw8mwizeObel2bJugENrawx3BrPc3MWpc6680FzYx7Z87eNy7iBQstWJJn
8lShNbq5/GU2uqbbtDsFtWMQcJSuew57CmXEl8IkCBngX3nqzYvF4fcY/5XnkY/i
nSTyLYFREV04tjo8IM44rKgrYd4iLkVgWMOh9lCNVrOf/irn7aHs3LMGgqBJZ1uu
lURLUOYoW758kixawrTz7kScTZRvxEQyTEy7xeqSVkUEaqblbazb14vnIrIcBEhd
kE1kcP/5SoevL1EtGO+QzxYFVdPFKlPA8LG6UKRob6Da9gdRVYDCliQzLWJFNh9j
6RmongXs1HuVMe5iRpx8f1GWz5m/WSWTuDP0KoDiyuDgPZUFUcYQMGTC2dSBDtlg
c6KXBUYM0T4lwhAo70fzzXSH6aN2u93KQxor4gvwX+tD0A9PXsGF0k6GloLQxoNW
IwCxbMMT9w2e1okDSMjjGIyEiVvw65NuNEyNUelJh02v3lMRozjpNd26nIbWhYr8
N9Rw3NSKE2HudYjutazXzucsoYy4h8Ri9mpQQjPc8XhZLHbqbsxSTCl5I0KA3LRz
hICVSzuex4LV46c6yy7ly7reYTtSlpz5QrF+gE9zeUoQGx7d1J2ApICOs7i1posp
FvlWFJawIqDJF4BZ9X3rfNi/7eFDIvI/CSkvkKqxdS9hlfc0ZVobXaFZcl1Nuw3I
2tGx4KHLFY/szRIXKr3ZQP9gB6SK0ENYR1zzSsxdg252ZAmKsS5/XWJfEmagv38X
8ipOjHRzi76oNTVFzfCLPDIHhyHGSeZbCuCsxXm7vrSM6W3yzdL6kT8Pju0ckdEm
XtPBTJtypgi+onriGQdeCsz9cddQJ5iwB61/hfohcjJshd5qIVSQ8xf7UL0KTirP
Vdyc9ZYODHszn4zc3rNdZ825easLyeOfxKcLIxlRBSL+iAcAFzEIFYIaLGQn2vd4
X//KMGHpKkCWAh5LyIHV1GpnJHM1JYCp9huLwaW1jnvuISpCfjR+R8iB7ui7yMoS
fcQfC+TyxnkgwPXH3V5ox0PgoHFuAfrRpdyN+Cp0Gs6sB5Wl4icLEKryL9o3+6Uw
vo2+8yhnaXy6It41KZV3V0oaj4BpUCZR+3YjUuWD/y2WRQqyg1iOGWl9ps1dMi7z
6Nhd9LXVTHxgLknwvzY9/3UCqYDE1W2JPKiUXeMCPKANwzOP0mwayejTh/EvZB6l
KLUAPo4AHvO8vdVPqKMG4Hl92jVWoRVW4GmAcjFrMnseN6UcreAt/cMSpNvRAnG1
Jc+WHQSUvO7UCHKHEsVo6/mzxETX4+CmcggNH7/f/IWlkHZbyzMfgAmwk2kYGYun
fcFG6esnqQNSr7DKwYQsFN38v0JXacco56Vd7gh8jwxBmdEPVjg5Ek2kvWc/6RbL
LFWHiyakBRsDLmB9FxOtR+3Kuj/fwKaGF95GYgHB+xBzJd1hakI9y2lK18gvysAk
y2nABRtBctz4d+i24Gv6a17ytpogN4ZqiTzY+HV9EQqZpl/Tl8meGoDUp0upA6nY
K52oXRaAgnPADEkR9jH06FQQu3r2k2ZZbhmQ44JaN9ayAWhljFd8CwY6qp284T5u
VQAusGsvXYeTHhLYsARz6JtEZMO16DwSF3RbiLMpt1zyjxiR5+dFwOQ+KucSp75+
Yr2wqjp01AKr0Kbyy/UHzcY7Zea0jwsMRhEaulDO8VLthNIHhOGTnJ8zkcow0zNN
eTlAMIvznpcK1hZXimv9iJ4Wnw5I7Qn6sKS5bgdByeyh/IpwVrCWjUnybP0Li2MB
W+BoCWNUlapis/MZfbhtqD+dBtuTm1xdtYeui4hC1hgw/oy1A2zDlpRGbLj8KAcX
YreGZG/nd6LSnpzkaZvTJI1eFPz2KiDGfq0xHcG07x8BUD5f2TBrwbDlhXedcNZr
39VuTkpgeswzHr9w8eEYMTjPMDS8btPsrircUztk+dyz3wyR4Z0RMB1omHEJgcJu
y1xQebS54jKGIJx7BX7SrKSmyqEEP+o2+GRQBse9EirzwDwZenVBTPgFiTc3zC5B
FnxdX+WMTPkifOKN8o18xOdIp2/WklgLAWAKqaQcQ1qzPV01ZyotigeLnTbFPH7n
6fdi8oP9JYDl4u1/dne1SHw+VbZFy+gUS+lR7mDzfGKA3XsKgFNImv6Hh3IVHuUg
V4AhPGlc43YdOFq++fwMcZthDeRvaol/vTCio1R5rVjJ2UshJxyB43qUWzrq3ML5
qb/tizw7vXsBJuLWG9KWFwav87eaFnR9L1qqe0ESiB9bL9KMp82krEWDB0ekY9O+
RTRsbVVYR/rqfjkxzEfw4McTXeIPdL+HjkFKt6MWVmTeTmLSP4DxAketw6fueulY
YdSO8k2RFXvaa7j/kNjhsxSckd1UsI2Xq7+I47Tyn0YI/NTmb/I43mWJZPZ7WZL/
LkL8XwbP6/pvoXPXrKUHwJOy7Z2I5lV/5rFoc7cgOu5ERB3fJSXBPIpzve6d0/WG
oDqs6hUKPA4nsDch49N3eXVeI+yOuJll45/sUtEwtR9Wsbffl66hYDXh3yVN1/Ed
7oSV9C24c70FhYL8rtuw85/YAN/YaiLKUav9cb2G7/jGYQihXLOG7bXZor4FQK4b
w1v/C7Y+n99h0NLe8pnKacdWwuTm8/dJXHhtQA6eA2QvuBx3QJOTGhqXMw2B4SZP
djaFCCzU1g/lOg8v98ZU2dd28EtorEgT69JowgNuXfKig3IbN36DJXgLIuBXTE15
1ZG2esU19iuSG8sXjOWM9jT978tV4ZDhfAOL6OqSZhvDp7zgzgCYyw2svOQYT5TK
hOwWv5THc0/ihXv4LmpZJUlKZuIzq5AvOAmWwYimC+MRqiZ8hOltvIzaMjrsdrkq
nX0yNj4Fk4qX2doDC34TNoCJq7S3l5HrPeJPKvmvAdv9nVnKKJ7LfPKST+ns5ruT
Jt6NxLcBwCh8irkCJMQ88jUoZxq79vldKVKyncAAbGr7df7kGghGK6z2vcPw/sMc
zyavYzwCHSK9gIioaY7tseusGPOgSvQ+1nTp+mgjU6RUH3J8p6xA7cOML/A+OwyK
3FDsPHau++kZFuUI3BgTkkst2GWu+eM4rpcVyQ7uPbeyPPOugy00nFj9+qXqVkIE
9GRokfoAuER5yVqcv96Z8sx85crrevtMLk6FHgDrRrSlMy/j+AmF8DVIUKo4KwuZ
y55qK1/d7lqp8u0+sYoO7eVqmDwjikX7Z5/H+OArcLjBWksUCpsacx4/AVQ7jUKU
KluNMs5cNX7MbWQUEeQlKSKAqbsaQqCqYZywiunGFj6oo+24u4G4OFo202TrRhoM
8zyGaNUYkC7ypwttYAxSithVL+o9DLmvhz2d2Hlj9JUoqSqGgRDhmOdSAsDiBtC+
8eru3BKkX68GQIeLzTHS4lep3U2V83AMwFWXycmw6HzdQb4RQFSL2nTxDXSjXso+
3Q3WhKAffy+kogfY6fCVTqTCuu4WH5FM2slH6IEBfEtqkJtwiHwrFA35rdB3bsmS
pIlbhBLZS7eiIZUZAyiDheKMYAeziigPhPKQIqmjz0sH3m8xPPp24jkIiTuF/GJy
KtQLvCbiD4aOLqocfGYFxCDuyDUI+WuuHLzAfsoKeFcHWxUildjLgGqyTI8wUaCl
TjH3E26oYGXQNTOJbYEXljFEbR/e3sevGN00dL+dHYoC3y/42yAKWW5SnNAGWgbZ
bApvXUURizLn8NNWbwLc00caPzc9QXqWCQcmvQsOH2GXTAV7cJQMZsck6YehbBWj
z8YJ/COZAqQuKvCLAOK7Uq1+UgXAiiBS3Mt+h8hjoXk9q0BsW63g3y++ZdfNjOIO
aOboTN/WXhzg98tUkhA7xrUszXT7LGiipyK/70d++pPGZsr53VJbZERQTiXye+Rz
aK8cbsVMCf7AFFz+JRMjaxWx8WN/6YTmv9MAKGXjnAjzAp2zOQktInTXsjJvQode
lhE2sx0XGk79j+JxdbJyH3FbpxVWSZrL79oG5ufvL3mNazeW9zt2U3+NXfOAuFVv
ipNk34h+dhJzUsM9a8Sro1czOfTTN5WLC3XeePQLbOoZ9bzjHJHraFofj/TDnlOx
OoLTd2gq5AFfgB3/p0lvWE7MSiqU/xWzLOc4YJbJrJ7bAPHIi/lfJCmKeOjodS3c
bAD+4BiG7fLL3rGjVSywN9NJXWoGKJpXzQgBvR1z/u5gryBXN7njSBrklHyTDJty
G0xVdvHvR3UiFCa9Tqy8+6qX6ejVGjKxhI4a+tG/UYuAsZKTburT3NoYaoTKRET+
NaMM48q/qHmb2Pqiy2uxA8YMOipn0KYhDRdY9ylchB8XRm5arnVizu8Q0W42ddsI
qEdps32Rb9Trg8kIGvHGNkJMnr5fV4zJXnWAuHhL+GGhG2pB4yKK8KWLnI+FgQKn
7/y+LC0a17AKp64NDaop153Cb73ckjBWfD2POBqMt4Ebxcx/I4kOiiOHjGARTg31
FSRR0ukqIAPJGnvSFXGjliS0xWvzBYnwI+a3x6iAmwgqfMPdS75lvLYnRJhGPKrj
gO10AiRtzxG9T6QuCP6rXY2Na+rph6vPcaqHNi1rqQFTRYg26lv6kfnTeJTmk4DK
UpH2bmxrmLddOMDDLmev5AF6VE9Sa1SVPaq5VLGymKV8Ka+NPMTfZFGKJZtDBRU7
Doyb8X+tPFLQDackSPApTWJSbYFNAdcUMzWRifMbESmnM9Eo7HsjTlC9xm9P+MVL
LPvqnq/pC4jC7Y0vPnPcnr3iGxFXLKdDW4rT+MLsgjQ7CUyfWQGmFWGZOxhH7TxA
QNpKXpHrJm+kv0BgIP9a3xAWSU7JY4jOVpT0Vr7LzakcJ3Pp5HUsPVZDIu9qWVWX
IfvFUfqltRLiDGiYcY/yDM4WEQkqz0Fj4VFlxBkIMaSb/6JURqhtzDm1gJZZYOOQ
tnmcVMLYGnLrpU5L8WV5x8mXDxxUpNFg+FvNHFKYAtQICBx90/zwq8KwkDAn3/E/
Aoa4ylzzC7f2eVYLJFK9TThnfOUh8puZZ5zHJHwUXY+JybouvMtWSu6bYO3nrXj5
SNALq3Ng1OdONwpPbOWEPYBxnMmbUgORovsEdvz0EULPn+k1oj48P1mGVocwotzS
o0qXVgprAl3UyETZqNpDGLNFhbOCTKW/cVSsWCjuiwJJ73MwUnVNqKXbc+RZHqwF
pCBhgbw3tv2LaX0SpMd597YfuJ2GK8HW/Q7RP2spsv6wNVxkfmbPttR5ZWGzc0G3
xuHPjGvpR0WODaSgoh1LDTKrqwRUNGKtRwz8/YR07laj2s9p2jVqvXiVXX4An/xb
atk/jCzrnfazw4G3HooH0m0VhBHDUcqJoTm9hMyJI+OF2DoyXvnZlbEM+jefWjHy
XUBkErkav/b5sOV/LV3bgQKl/8iZQWR5SFTexxeN05nd189g5HteDVsYofAYjOEz
cuJglGF8hv2Juk6bfbvWTsQRmgxx+DIErc0nuar7LyVFsq1DExjChtxJetwV9B4k
MhDvQ0kaSbmB5JLdKuy20BnhELJZR0xNZVUMMcv0AR1FK1kF5KznNVAKwrtGwWEo
5hm2H0xaKUIdUEJN+nV/r5h4ekqKcbrb6I4JxW8g1+x6ORJGdP4l4QxaksxZ7GY1
+LKoE30l5XRkIqmFaBntWp4zpXbxXetEyIKiVHWgQU1afVqgSZmF15P4aRCswWlV
8kKyo7Gj67BqeqIWT6ZfBBJHVeGQqiNAtpslQdlRCPsb5DVTJvWKgzvI0fagn9QV
d0eGlQAJW++Z2b5bcom2t6CYpTuMNokkxmh/dxtwLa/ZqH83uj4mJlNJ6B+eulL+
Au0KGzszJtvBKKFSas63D11zVvh8CxEIUutHEP8MCZ+Y7Kidv9dzYGV9f5Lo2n5B
+iIdkfBSbJrlBhzLWypD2ylIgI7BjtWZF7uO9unguO8PCbEYX5N7nf5CoKp/+O/D
wLB2h7fmUlycSds20XYcOzssSfDM9tw1GzjFVg8pjjzQlHq7R74+rjvRzFK02PSL
4k/ECReVwdvEWQGNtraUMzo/C0QVLWmHD+G5DyI0G3M9WZAwhggpgG7ibipHNe3D
cVrwEzu+9TsSvcme+/wQAUon+bUV4MunJDu3k4/IKfJvot9tGz42tcn+R+nWZ5XN
svwocfLJT2Y5bvSKtK5wbuvevpN4PF7DeA512SNT06+UtYBWdX9PBl5fYaXJ7ygP
YQ73u29ODfKW2zuB+7gKMiwGpwkuenJWJW47gKJkuof07QYEdL3AgaXRPWQSV9zN
E2j7UcbUHoDUPORT2HlZNOJqsItp0FFQgAPT8cJOAtH8nPEEsKXSwRwmeL2uTeKf
yiWRyEEVpoRl68AWT8oUeWb0kzFo729X7ae8579P9mSUpCaqMIbaUYXhEs7tj+He
qX/k7RcqJqBbm3X6SCBm878YghUuddb2yGpY+xI7GCbfuTGBuW8XfLuDUTA7j8Jk
9cwdhjxdISPBuQH+xqPiGSuLG/01zYayGHfwfjhjmeNC3Cr18NG0VgcHSS6goUll
GwNnh3xNqwT8tRYdqcXWgNsfFZJnTSWqAIeNb3bKzc0opF1MrNsmIa6JQXEq9tnG
6W2sg4/5Yxy06aOdbEgl8B26fJIhQg4URpdSQkoPKaH8OuBCMakGTtMUMGEwuLTl
rYpa9C6O+HKEjVZFcXrtNd2OPQD0gsgtz+LbX804hjvEvO9E/nP2BhRxA1HzeJyX
mbC7/Jsm176QwWRsIeDuZNESdevOIWcrGEmgSQ9GbHvodvRzi/K3xcaiCVdX02Yo
wNm/1jUb5KrozMCqGLa7mFX3tMwMA8x/OjqW4Z/7G/z/SadCIdPfRE0WP26EPoka
YW16lxYxr8GsACmzILaL1isRLlPxrhgkna4dOOd9Me0JAEMgWPszHHcE66aE7dAb
CWcXDBXYhSAyTLZpB81Q/iBuN994+0iQ1tvrE7NQRXocx0LbfIHhUC35uSlTiax7
vL4ZYuZUtvYw5IL/Kl1sgQJcPNgPJIJIVkH1qtg2+ancBywJmX/ARse0cOp+nYH0
WZhBdAdxsBKnjVkxa9V2a0fUXTJaUS8AOD2kmkh6CpYyYx1rz0s9rkfsqADyYYXN
lRq5Yzajy+LeGqdOVOM0y2b04NRzE650R6u9vKKuFhs76JoJKLd2VEYgHY9ubhYt
EmRzGKulIIWE7qRzJ3MO2KGaZGNl7v5oa8DtlVPstwFH39IcFYpir5wm555IbnAJ
PVhBtVrPgAh/PD+hpmUrOyQqD/bL6UyT7O0YRaUtcqHPpZpwA00aP5YWV1UEstr+
guBvczC2cdSHizcpVACxnZN+aNtc6zWIMF0btjLR7Grt0Vss0BVJa9rzcaAgZIRi
jlRfYFI+Q/RtrO/DX5bQ9kteuc57StT2LhfZ4JYXlWvVda0LZaXTcmAkMznzYMyZ
RVsNAXxAWIxY9mGj0roOQLyZlbQkX83AmUj+qIvcjvfQWTo6WT3idnf7zm1YrCOA
q10s3CExyHCP6iQEWY63NhsLeBI5YDEjQiuGErMz/oCcylMm6WOQlSmG6R+0L9kw
5LtxPuud99g8NZoGIIVF2lDQYtXQ9nUv7VLvg43B5Jupe8DSfbj1R/tfznk9XmEi
ibeDbEvHseq68P0HpC/VoNWMJDudSn+DVQ00/YuqWQ4XBXDZhLRycDQRBCxqkynA
G+Y+CoNhIWbo+r7vO1exI0z9088vtUpExVGu+unCRom6tN0sKBMCvB+gm96hAjLH
SUoS/c3uMvqXEPqf3kPcN7xkf4LOapOxKqj2pIWZ7nbSHekxiCl3q60oJ5jYWT61
RM0PSESfuhXLCZd0RPN1eQIcuNi4C0hXZ6cgb+XA6GXMd6Dkj2ZsgjCFgfooFMaD
TSA6l0CDWG9qpykD0tvdHsbBXfWvyg7R/+QBmQcrwd/Ll7wPM0Dbmrmksyd4CG4L
qnwVlFep5Us1I079R8r0IKRGtagmBGSFP065i13JnM4TczqcIVAWHJ29rkM+ROda
DEAmrHGPOszQZCDMftPHALlk5dGsbcQ+AMxkna7m79ewJo2bv+yOTvcrl2nHle4R
7MlvuK51un6xGppT7wB7WGDSZ0D3P1W5sIZWI7RPYy4g1Eh1GpZDo0o0MhqjvSCh
c0vVrtWfSdz+rO+dd8fLOm1tUtqyfSFppi/4xIVVqyIsmsZ+Q1eQjTgxz00HtzDf
wAzoc2yeJqELEoge1pfUl667LF6H7xGz6OXPjU6k0A+FhBrnJKgRZSaUKwpBxbta
/gK1QW/BQeIH7jLtlrvOW++SI/Tfn6clWeV4VSq4HIrPPDO8VK50mFiM4/CJbvDS
uILdP/y8FM4ikl3QJM88XGuGuipJvtWJxk/cv/YLMMiCRVzSmy5rQVMitWk1Gt+Q
IirPLdnk6t9F2ZXeeECW7d28bLaEw5mQP9zIptqvkS6mbcTwq1A1Qd3RdLd5CeBT
YXkZpyb7QVaavSiRN+O66u32boXKWb0NirIkdTK7N/QsRUWsj+o/RiHbnGCNQvDk
N9gosm6IQoXTNDDsvPm13v6IjskXFgK9F1hBHkYh3KKoWCE2DAwjtwAOXw6eD1jL
cNQlmzf+O2Hw94EcmaOZGPrHi7huJq/gb6WUiJsxsW5hMyFpfRXn0IwGYXOUk2gT
WxksomZMr+/A/79T4D8Agt+5kMyfAvZhG/NMss1QGNiTRUdtDCw5nq1FfeARIeC+
pgtHkxUt0VwtJRrrLOctIgb7Zw3AbmrV3oaRwNUAanUTzSJ8VaLdP3mvv7vCwo7v
TC5zCL41Jfp7U1sfeMcwshuMpuBpldBnXea9SCK2GLCyObVciF+nfpYkEecYqjrc
qChQSXl3FDBl3NtY3XCF4oV9RuQHcMDOAYf8S1P0ikTvkFR9DR8VZbdCIdtfjOAK
XSe9b0c43lrMvmxLmr+5k+oH7LBZw5s3PCwstkIt28sLv7qsfCR3MKR74uLCI+gt
7ZsUeA5Zm/fHTfuErKPG0aL7Va8b9I2qMoDczMqvsoFhVsfeGbk/hX+7+NGGhHHg
8CjMnkcAQGt2VTg8x0mY8cRHoE+2T4B0aZDijpeSbLkFwQkWVxRKaP9pcQgufXdX
SWF+vBgcLzvE90AEcJJpVat69pWuPqjNnPayb11mlpeeYcxChVuunvVE9PCBc3TX
ncSfiHP7JUG3WiA8nQl1hnqgjjaPj8+miPH+mSWd1QTFbHPm8A96O4M5OnWnSGWf
p6jw/Nt3afIQ1lHJLtr87Qsp/mFzW4sSv8KbPvgYOsqpkE178laDQBVGKrMBdzgs
5ks/2jMMMTEzg5DDUXIWZgF5bvWll3dF8B1STsBoSsn23gedZXAOxDqtnn1uxIg6
/vb//wqoB0cH1hOGKMD5hKOBxAx+36RWKOXI/wWPbbd3gd31sdF8sRhO8uAdFD5f
0ZjEx2/dgCICju7UX4LUA3HZ+tQleR67UkbXOPUhSinRrBl0ZN/G7rVTqwrjqKQ6
IJW0X0PnOqUSMtYNSUcHI7fW/LE7Q/cRpP63IkXdVRX16BbcwXYldiPlLWkQf04w
4dJio4z8TYLKvVpyBaRYR6xixfS1dulOLW7uporzj9ZHPHerjJxYSvhkeS2sNsPv
TlZVDHtkUiWVL1YN9ANCBu7L1Y4Sc5chPJJZzs9TMu0SK7TDvacudQTZ7/TWvtu2
V4xgV/z8AZ+5qWc6lPSJDUfXmgi5Uamm3Zu7fvaNUQKQj8g/EotZ66sXfG5SIKJA
Cpk4ZbCfCxENHopcSo5dh8Q3YYSqpi8HryEBp44ZAGLFD59LwFt+3QysNUcsJWZj
n7vi0hvRybyfGXzoRUcD6X1jsxnVID6lzDhdlJHAhT5PXzPxaRl7/MyKYM98I0hX
QKsFhsd6rfvY71uJYDMBdCnRklmWKrTx01JDMZnrW9RonAi/jQhxz+ITaycD04K9
3fldSU/E+mPI0ZmxCPJB15XuM92ZjpTjoDDzhxu8yj1Iv81ITRroWO+Zwzm/qMUt
hSbtcp4n2e3M4j9JLM9vdUHSTvwbe5+9/2uPNKEN6vhmg8DLTk6EjvycH7jnHiDv
8eYaS8orz6BAcQuHnV+JBJlr4FrUfKx6pB5T9KLNr3pO4FgSCDQWMvGmMlQ+8/ao
Kb2VnIr/qAAbYq/4K6McScOdVgng8SHXpqUI4ANMFWWUOKIeCy+FFmU4R53f/VHi
Upu0dhxLPjxvTRRDjVHmwbJOCGvVL3ffbvzvT31wXmqj9UjespvZJvXJsH9VYzcC
913IziL4ePKlNX1zBgiO+vyp3xCXKF7f79VQ/4exNDgnRU1zLBD9r8CSxQcaT7pP
BIFmzq4iGJFwuAjvOdNq4BBMfWbAhkdHqZBW0sNU9OcysmxbAu3/F+tXQfAY9yqC
aFaOYOMXgw0cn8lPU4tToQxjMvnA4WhimuYFxQejjPZBSWJ5pVX0ioKuAqV2lw5l
8P20NyZW0sx5PtRqVM1eZP+x6RYg+syZeJpn61f1vbu6WiPlQLMEU2CbDiu3ATR9
BSz8rj6z8+rm9KQUse2YPj0ZBkT16RwRg0uKB1iTgx+4u4BvgaTdEdVqftBuEFpn
jNmRgukZDR93IIKILUWksrlj2uJrbM2MWM9vVhw6Cn+JcF5CPvpYjewM5qx3S3ve
DMGLe8bn+RL7P25GD0Qj9E2D5w0g1ubOwGcHrMMPlmrUkWVG6AmNVaux089LZ/j4
hni7uwtGjQeJ6DfwJ/kLs9kChFh1f2E/quxZJoJ6uuTvwOW6Yz2c4EqY5MVXUieC
U+qjFSI08xp1CSpO3q7wBO9JD+XaylQBBaDVdLAX591ywz4FGdqzF/h46lEGFE+D
LwM4xfN6qbVS0mbTiFoQf9nfHa3Q1Sd8V5dsspcgvbNxsJichQn2fqtZRTNXUqR1
mH2mI4QLGIf3Xttr5naE+3JpqaWPMpVLhVKXq3wjhGk4eitAzMKL1qyeJg09rU+4
u3u8/J6rDI51dv4IQvO9m2Lk8gNEXBFU/9sz/bvszBDpkvzZqCJXxdiRDiZd9RYN
2GYj44cWxLm+VMNl4EnYtpGODkQk8yxTASShHD4W/o+iPYrd8ohLNhiG3XA02vtx
U3whcaNcWkptP4FIfOjIYRFs3MzLL525QkSqc6Y2CuCGFEPNqxBMMyKbx7dYiktT
e/DFBkCaPmt4d/8LAabE9h3ZYlAwMj2Wxwr4mwIC1Ie4lqEd+pcRzb+Pe8HHkDtn
Ke1k3ZAWZKeO/Y6lWyYZD+sG8KZ5KM84VMblyWAn5W/HkRPJp55no/Qr7Vc7KCsN
+3Rvn3DYOgrNsyMNaH1IJyTshFQr9uxM9lPr5y85pI/LowkLd7tiN4PvU36VADcs
EHMwvq4Me0zg8qkibS7JRfEjQhWMWYFwh0SNi9e/yDZRdvodzgAdtl+K0kj81P+h
xUlAf7zVWNzDsSxwVMPf6QE3r1vJsRD3TQeKhqCR6RxW6agTyTrZF0oAoblr4Jsb
iEw4VmM3aiMOKWj5vhb0hsCJKzVec/D2/5Mat1lWr8Rm0etkfFYxI2YZJKbxASPL
bV7UXCA2aQDGwRocJDEDuRxD3hee9Yeb4a8S27MJb6OXZziFf9mmCAXEw0S07GGI
OUuM601hfKy61+LevncXdlgFITtQHR0N412/+Ng7dHHbjBCxg8JfJMlZvm4l2mCI
qDWiQsVkt6ZL2SMIX7y1M0vLFlGJhcL9uULK+9JyIaoTkA/FdkUbLYAKkKOyZ5pe
7YyoM7gW/GL55wChnWr3SzRrKQ8jwyrZp5es5sPSJlhd4bCb2jKJMteIMjnIfBB8
MqxyYLzwgZrnBUccXuIm2PTQ5sw4+AGvloK9LZHVBCrX81XAxR2XX+hCbXW/uQHW
zb0Z+R5HT51u95EsYTONgbOnc7Yf5XfNrRBHuRzRnr4oa66/FL0viYWcLY6V2LL+
xyS1Es/39YpFIf9XLYnSrkG+9xF+2lCaF9P7wixjE6f6m6n6V09ESRLyndYHBEDA
hY1bcVnQ9fXi+2iPa8QgMBTIgcY+p7/KelW0t78fzjip3YmQxpVMX9t1iZ+CRLPP
naadou/FYYri3aC7oFYqJOZib+4mgB7fFvto2NJPfSIhbxc9oXJuiGWluGqUtbuD
ChLbYgytKghx/DQn/fY3Tx4EM7p8ogiaXgv0giTcKZLbsx7PquVvLg+K9blSayS+
0h8Wu/aGedwKz8EwIovcrQ09H8lQaaZ03DvkKHnC6uh3nd8DthnLUAxpd0tXIt3A
RGDPa1wrM1kDLPx8Ig873yHYrYPscc1FiLpZ3YXiFCpxShFB8MQpFQN2TKKRigxK
LvH/VLdjGkK9EEuT99YbEphwQvpMN7eMyOtJPItrFBKUss5mz1fiD4Vso5HVuBJq
a2CwOv09mQ8YG2eGrXcifdQQszGJhDxOJmzFq/7U0VAzRozCjirxFcAKbHKp+xiB
Rb7y/KQ6oPChQVyokZKmW9xQslN65DVCZumOCOFnzBdLebGWdooHFHHpLmqwvtee
0CBz863G/Mlpe0+L/i1rkx0LqZ8LBv8OF+cQUqQMW9/zyJqrzbArDTH5ErYPjC7r
Y+tcBvtcGOHHPhHAmxG91WSeBvzxjxiJXZc0mClAqgsC44IOI5cgD/UnoKExZTFn
bGP2YS89azpuyTUmbMZtyCyxNZStv6Gu80sy3kHWB+MkCsx0aAjgglWT0gm3Hdwq
NVQ7lc5noK3rAAAbE2Jf21WGgl0UbTnmsnvn8fe+SlTH0DSS7rbd2Xysg3byv/MQ
7f3jD5b9rmKDaGumf/25DTuIvkVk/MAXXoTZFxoFedztnkPV37L5+CMrf6sV56CR
GcwQxguj7h72k4WJpCTblrth+4qqWTkrfiI8g9y8NE00lUdbllVR/eI4A1lF9KFc
lwQpLxl6qr0RRDbCJqJG/vJXMJIqXD9GieUP3MRc2JWt6Oawk0npbuX0XPI8qi/h
VYK1Ue4uDYA+wcTy1ji5alg+uuLdITnwiPSkJ90aIBCo2mF2cdjfO2apJkCRhk/u
xvMbKRakFbvGWMJ+DR/BJvDZMGdZTdc8tC6V6dbD87XnsFmBEBs1+3ryXvWBCzl0
xHP+egYG8hjaAZdGgXPiHBKvXu81xqaqvB6+e2dj+L4FIkbKhA64Dd/KSam8/fGg
iYStUKO6Ry6A2cwDTflQPYa9mhQnecKRTgyKcAXte9MqSgyiuHsEoKv7ogETU2tC
y4ECSTKowkyQqKcZOwxGnnYNkGSnwiQe7Y6cg0aHfTQLo0bMCYvNPnG5SXxT0f9A
BJYMd3la4vv8Lj0UHaaEA4e2pLrSLL9tcdfyH/jveE2LnaHmvYQBXo4JDxN5tOsh
sdz8dry0Mlmc8GpqF/pJz0O5Yf/82LppOh/fZ+JcXXpRCycl+uQLkKNCEqjJwnni
T53FYs6de4WitJ3WMumS5eR4zZGm6KgDX2tKrpCRXVtSy42m8hO6mgUU/dHcPigX
gbcxpocMIMyA5dDQiqutjHpXduxC1nnDjtas91enzAnJOtu0fi++bkzWahgX73+Y
fnvE07QWzr5CAPPy3cAN5kSU+JuRz1U93atTxXr0A1kw7/AEgQJgDfUplXFigV5y
nJxHoQs86Og5BqyX0p3NOWomywbqzmYP5IrfqgLaViM8ymIZFFt74cwMchFyD/nB
t9c9IFGgcLfsSb+0h0AjyQ5ykYewdnfXKJ31uHKTyS5IAe+Xq8QDUTLchChvfAPG
LUvJiax3VVf4KnW2dQoUah/n5nd/FHruxam8bbn2qadPoLAK2Rf+GGz7pi1sZqMc
5B3t9xSqWU2p8HMo2YLzGuegjp6XoTqeANZUhWDyOyE3cIwXRmPDj+flX6QR2XSP
ZuBKVuBpMZ+Ruc60gLN+Q6xyQdzL9WmcM7f6M27o8g7e30el7+T4Y89mjklLwQyx
lZE6H7LNsD5eNY7eJLxwnLDSeXlJPmbaKiBkjaxxQxjVEdsJsQPjHblg00+a62s8
wGd07sYpNYFXNxHKlx8ynXDpa2vTGbOXK2QCzdKqrUndkhjah/sdjR+HePyZev/N
Nq/jHT4lWRnF/sWaMsuRhA3YoNjmj9RwbXQRzinayYpfJTLVw7B5JnhZRp2AhDsj
LHZzJdbEsLe2XgIbEA+K/IeIohIiRBGmEw1ez8aeI4ts3xLaedeHIEuFf/fttaui
mUwM0ZRkMPf2OFSYFTsXq03VZ8M/rqCJrledW0XWYzWA+ldV+swHQbzV0Tj36/Tl
NpVt4bDEq+JVvn5wK0UeIxwR232raVHCVAdErUxpbhPZDM5hDRqzYE9Fexkz37Uf
ckcmE5NV+9E+8O58XwtTeFjan/lKi/IwapKn3iFDsgcCsMNKrzI49DUHG20fkSLb
8l6EcnmdRYHqsUprkdVlIel2oq/8hTCCsHP8ZcmHypZVGc1iucWiJ/sSO/1D3Dg+
qao864c2lB/zZYvltYvnhBrEPxv2k8XgfadR6HR887Qgl6PV04YEAKTUuy39mLcu
qeLAcJyvuCrjfdvEasFXTsnOGWM1lKDK7UjI7JIYdKYtIq16X9pWOs39xDOFy6oc
7MS6avpOJjJXNo11jGOKFgX8Tv16j6wH4Mob9nfnBKRS8yNw3e+azuuT31JLMRE7
s8SoRThLcgbMyKYnGPpnACkAWQAT1fpLs3byJZRCfMuyCkUom9tyz58UbKv6NDGL
XwcwZYfSsI95DKp2SC5S9sNr3uGmhC02wcimiWvYfe+HfK0FVtcca9qr6giZ5lJH
bEObjbXh8pbLtr2fbiRAqVHkNub+psvso5WT+qETq83FnP5xEoIMzwBvRYH0WS44
1QPmWJSZuwu0eAiQUQP/pgn2iYMRiiLfv0wUPSmaLE35RPlMkmzDSK3QChHUDUqG
SoslSzSeqRQBD+a7IE9wTC8rKbB6J4Aw2VvphAS8Whj8k0ONK8J+vSgwr2VUuFh6
Wp4X6VEFh8rEbojCp20dC1PwWNVf4mwXprpcnb7PNDqxMCGOl7UetGymYz9kxvSj
h6noORjGbG0keqUwRAJYT/mG7mlvK5r3ctfiqf1x9ro+M2W3V3b5ywnwB9LTjjYK
i1ZIK3SEwphXyTrLq13RfJ1+Lw0JmfGuqMPMKz5w+8WfNLrKNNnYUM6HROsg+sbO
tU1KnLTnHvwMUkrtcUYBkjuL6+j+tp/VSpPaMHSoFSr30MDMBcoLj8KBLqJtizbv
XWPNv7GUwpaSKWgt7cFa4/JyrNM2ciT8nhORdoovfX2gexcMQjddBMAjxSFM2FYA
XBUJkf/uuEpShIcD0COMtJrJBP5Af1+WsbTivOGxDwNP3WHBToIPLEiH66U4j6e/
f99ya1zXnq/kTNWh0sfIFzGm+x+D8bCRhiiAHrNm6oNaZbrwpI8w7pP0bOUev98J
666A6uGRJqvdN91tDintw4ALd5l+W3TlJxbmNX0PrzyrS/8I5wTXx5vVmVLIxRJ4
bUnUaxKbR9ALE1wC7J0GRgZ5DYakuY4qFTfDgU2MFmq5L5fEOXaCEmgiL2X8+YY/
+qnGEJUphSXtapAuZizpA0Q30AgnsWv4mC7RUw4HfR3rc51RMt2GgRGWh6fFVklG
CwhwvWjWKuHluOobjBVhYjuGnukM5LgQT8IjtV8J8M+L58Uht5VS5QVWgYPic1wR
0OG9zeIgRUNtx9PTLR4mgpKfZ9SP5q/Gsh7yydGLNxFJy9NYGRunp8CE80DB1tMZ
r//P+UCHuNF+t10DCpm8LrgDVs3ZxVC01AOxkfVuZVFSrgTwkV+wrTCCxcEzMPbs
egnTGYaC7RvJtkGaV0NeLJXF7+PH4/SA11fT3lj/zWN507KWzW3YT8OnYit/36OB
Q6Sv+arnh7wUDG3aoORVgwlhnwvbJqABOq+ypH91r33j9qa2RdEiknS2B2k/WYmK
V+Wsf8Qny3DSrdCBaEQIlzjwLDlTd1ksq/OOAiAdMDHw8n8PActJAz1gstLat6hf
ugv9LltmNUrsdOIQELAmAM8ZAO9HXjWjayHN7rX/KLqNT5t5x8RY7qf/2SiL11FH
fwf7E6drLzNW4QPK6J8W6suuMf3mcP7PJlG84fnIhIhQMwQIEjJrsEG7JOb6qXNY
aynj3s6OHv5rc1S5s5018/PNgJ/bJJjrpXVzaiXgTMGVhKwFz1YJ1pF+3Xb5I5bK
trtVw97ZpbO8BnNs3iAzhnEzA/S4x/edakx17b10OERBTzjEDyvQJ5sTdHHEuxhX
/qHO9e114MWYAeAmJzD3K+Kmsjeb47sBKbs65HwzmCM5ZB/PMx3V4J6EYUqHSWwG
MqMOkfZCmItsMJJdmFcUgd4feT+eRE/DLDiKlLpnM6z8VpK8APYRKW3gl5hE9/KP
jzHuvKeeTQuYpuBCMS+4EetU5yPRV9mpXJzDL1Mr3DLG7TB69n5O3m6F0cB3iQcC
/C3Y5o8dh5Rc1hD7jfHcTbB87Mtjw5MGkdf9tzrQMmBE0F7x5XqLV2TFdj+vCt3R
dgpq+7W55kUzrPoYjbBUr56OWV4vbfHBY9xJe75gESq0IYuPmwMlkZ0M6epr7oAd
WWpDfL3zPE0RLdm2epcviuLiTeOVTUW713xt0+MSkWlPZ+QGZNkQ92aS1GFWrNUi
pMA9EwAgFFdSpNz7PKPQsji0gGgIZhzDpLrJEo+uoEmJgJsTQyBEExRDVZdpb3IK
I//Sa+WFrBX8uzqi7S7rz5iHA3nPabSGH7pTo6jX46ag4bxFURtcoLnlU7EinDCn
zAwvRi8DgClcUu3epGQ7yptlcLFb+LARsJu1sXRXYIf0fJgy6w14mc8wc+dwu0Em
gnMWXW3a5pFr8Q3r6ncchx3UBPjqhoOerjrs1ycY3ujfj/1MAXQTEBnEiM9U6bk/
Nu8Ct+bnmjDGd3SwykzNDHG6ql+2xGBMdjoOeD9Al+Jvb37nXPE24uUL7V8QM3C6
Kva2vVA8UTqhm9cwNdcV2M16eyXsZJ7leESCe4dj7KqukF6NGCrA+5fSJfw1DCmq
YshnmfImA4LDsMqg23y+IBq0s1a5eKEWf0xL2RGwNRzw7iyEKymCH190HujoGS8q
J1WSAw0ka+KKkLG/xq4NFXPuKEzuxCX+YKSSr37NT8RA65E/Qf85gbqN8429c798
8+o6h7/Zw555p6TpBo6UZvggF++KK+atnCzNLV4zYl34R39vCF2UYntC6zhJmIMJ
vH/NH7p/pKevWlRYOomdbYosWtoD8LlgUR1mqENCHEPQvB0vGOis+C97oVm+hkzF
UMEMg2OmVTwgbBznnH1eOxJJeU6GYY3MuJ/U6O0ELE+iBx+Cd8bUxFX11QUdrmT0
glgZGGPboP6TvYNuyQM3je2yL5Y6Kc5E1bKVWFN7WGK0aSfrurYOGmxF4nlrfjfm
JOeNyTQfw4H55ricYrsnjFoqv29ewLqUig+QmxYYtTbU1/p7wNcIITEfrIyoXuyY
uqoLgLbebbLSzkdE2zWYyhWzPLKO4QdwPJ2/niHlZGfK1ll4KM2cGa3EVneewSR0
ytUAO2UneIOKoe8Jqw2iWvDdYT0RN2l7ZKqlgszL8w2jTZxoDjntl8f+GF9mlfmR
+r4BqP2PRuyqlMjRbdNMk1tdah0BOcz7hWZFX9NznEVr2ddU95ahj8SxWwFjMSZF
wmjUqvWph24ra+Qj4+AXsGexbQK9lRrw075aRVZuxDnI8jRphM36KRrVVK9E6kDL
J9Yv6m1Ni7F4BsA59VNhtZbMqq+d+OPNKzQ96dn6ylcKCjIBhUuqdAF1OqiHk6bV
VkFOKpPzxFnXPrqMNtICHIzPLjRTbav6F0B0mrQfzpJaHLbsoyGd2+FEnhvFEjbn
PTzauHi4aODHjVm+Ab1aQeFrkD5jB/zrCbP1OO4IkuEY0ERnTIQ+MyXvQ+Ncf713
rjfZrj2JuwAJ+h7zXXVRiXOK6b9/5OZqXTqaGSqda+mWCypkPq+TTpcCCrDSNPaX
J9x6nx7krLJRk/+AlEwNwNv5vD0bn7hg1kwjqxjd6NxQkhWryJKPZ2TW+aPWkLGj
sPwU3V3hO2sLldyfCAtXbbKVOo3uE3brFwV4/WVpqxTTS6EDmmyZBRadUOF4wVxV
Z9llUbRa9NuMAGx+STcoTLeX2rVIFYrLC72aIDfCgvdWzTbh0pm9hTvZN+2RyeIu
lxsL031V1gVvzZn27XcZyrEDTbQq/HETiYIxaF8iZEfQoPqFMGV0kxWipDJ+5GAJ
/YN1ytD7WgIVVfiJ41LxmpCNsCuSTUFGtdblM4j40Qkk2UI1BOXAHKR4lcbS7doq
hJnIuqyhiat1MlaNslwRyaR8PBLcIxjwH9Y0wPqU2Stt6gLgJ3ysq6k2S3JfQyvO
iNm8I4Bt34kXdsQuD55pnQi7TJJvGQZEqA+eSAXSKbTDs7h55McZw0pq/8Y2RaCD
MUgPMsjO+dlmQbIyAA8nEnXEFESpeTyMvZ0B2Lw610YRTP+NTeeOvRcLlxdRL7iB
VAG1zI3s8DUM4nIJVDMwK18vTfpX27Ni9sqL0awJEn0BSMbD2YePt1L5Frt6HQwn
iG60NM1sjuHPxo1r+DDUmtXKt7XHN/jjmqaQaaQhzt06tI4RsRo62kdtxe1LXCZ5
/n7X/E67fjO6IJVgPFZs1KPBQfX7P+m4n0gMFxkaHck6xJKIQyPjEmBDmKPSm0HJ
MZsosJPeF7+d5XsHAiGM5zmtN0LZJe+FJ8tD6xEGIE5QBcRGnMMmrQkhxc/Irroj
2zLlKLSGGORi50H1DsfItxf6gbWjEhLOyAU1E4OCtVhwOfcRU/MdXnDEBrwA5jtD
nj5sdYSGDax4o2l29h9LkWRNvO+/gExl0/Pqw5ieL4qMtItKnbl+igEU+9IkSBUZ
yuRkH8NnD2IPVlu11tXeBvxv9o7QwTAVpg7Quzix8QRBOpYh2iQzOTlQaPR6AXxT
EpTc0VyYngtkpaD/1nE1MI6cZZoc5AvMbXbvqP6dYMLW042ddTcTPFr5jzIlGDYw
tn2r3apqP3lb7mY357pBC+QbSNHjoyUCmUXP4+zX0gVmnTJFFJ5uGZAjYR3kBVBG
8irPAC9YHVslxTDMjohlDmJkumr+gyr3S4PWirpRSqJLIojS/N7rz6AWOlifx8lh
BPXopanguODpTVr53ZXt8v7fNHD1OiPIcY2chLtmL9TdF7Da/L9OKR/RoBhZcVdA
2ahLIXMM6bGlhRfDnM2wuNi7iUr56MHqUE4eAPAfRpR6J2kClZ+ZcODOGKS55mDO
7N06Rv71lgXx0mKvQkGkODci0AE1LcUb/Th8MzhkknUKTt6H7Q740T2NciGMWiqD
5EpqxiXiS8ib80iX50CncG+VPqLCnQeuDGFBr9b7LwkjskMJ312Dtqsk5t+KCMKH
fl8ufbhgPCqVMV96bgjQlyY+0Shj7alohK3EjKjAwq3aCfRFuVfmpAn2JnEPvAPU
Rti3yA3nMrLcaQgCaNtvZ+drffmQqz+L6eyr6hJPdxDlpd4BlY5g6Wj87Kv4frNf
2xWmJm3/RJkDubq2gtFPn0whZvYNkBf5WVvGvn5sb9MMzTjg6WKfDYXpqrfo0QN9
v2N32LpIqG4YOOu0kHSAtqFacJTY4u4o0V62CHGdbmGUanLdIo1Nt0g/e7nmRBIk
8MDWdUlk7N6D5dlwa1wkJv9QbTOiik9xpWRx7aMc5rithhaGwbyyARBzIXbeOWsB
6xu7Sg6Q1Ud5ycyn7nEN2kRurF/Z4dRSt/DKkKdAdnbRHtUnEPbSBYr2NnqkfyT7
pKD2elUkKa64vafMa9B5ARxN1rJsoljvxV1MFqQ9XZpwD0loZtsyhl2JLOgIIvDZ
WpzyPgFHjpHDR5wnLJTY9zYZlJi+AHxx3tPPsZMXNiW8eaAzqZHro167os2+A/9h
ITW21ofEVFbNrJIDUhYvv2TvhhzqCSYTr/r7ThhI+yASnss9+jgP/YygaQCXx363
GKQvDbkVpVhyMrSVNiVAcYUC7NgidxWh/e8SvC87EZnp5mDe251mfCtbTyVeTzLl
nQu7nqa5NnwVt5lrz9zYoVKxw/WmjAV4ud0AF0lS3KBHpxiu1qo2dtNDzQ7cHL8h
fpgp/MceyrxL+VkJrCbpNbQzCumP6aBs8cEhdbauTLzAIXEJTUICluT8fVUk2M26
9QNHnmORU5DR1M71KRcfQGzdd9F2Qo7DOZCCNkXzmfG1OlfS001NnPyaKwcqAufF
zrgLcK36JybrhuF9alav/nc9kTwxOYugUfpCrttdhn5Dm5m300tI5pYDlBmArv+G
fOy2iheXhTNix093wq4NX948qwrg7KFkrorIqehGiw36Mc2KXpiwnPmxmY2FwLV9
om1rTisEThDA4Ax8FtkRyV2shD6i7bj2tTHvdair2PwYYsRPluYCCTKSQBPkrw9x
ecq2pfeyY3sz2Aqa3dO0oOQvA9uJMWqsoOwqnMDp7cd0+ZpDL8FgV61ki1KCY9+t
BLTRYoH+Mpg8ZhLmhd9TdotgUHklcKFGuh4cfiJppzhc25hCwmGrlEX7lIHITNz2
Z+97qWx4rx9n8iBLHjSOdCgZC3BfQs0H6AX8H3hBhXfkwUVvJ3Rn6P4sT+Vj9E73
LQSIyXOKbIwUi5DV5qaH4VcAnZXT5KowyHHdwnH0Qw7eBdmdnllPTQ8NwpmdWDna
EuvlmM5VJoMd9ELNeHgX3vFgZm2Ss0p2d0dI55mo+2lk/zNZSTOORU8zT8sL8/RC
A0JZNaf5PiMl9tzpRoQjmTAV1XiOFZXkwMq1VW2fTHjZliE7qwLeQrXOY858HlFG
JDxizKrRAEe9xt1Oe7t+v4qbEjVZYGBILagsIkmIzzs1yfNlHxDeWgXgCo76fSg/
hg5OP5ip0KBJgNpIS8ODmEOaneFl2aD8pKK9V79pSqQcsm5npeRx09YRoDTc5H+A
lEb+7j4o0KIUHvKGznFdiVuEFUxNwQfQZ7GwLFurGX7t3gPifUdI1PLMNom1QC06
4ZDABWRsv0ukAMgFtnkDH9wfXMpNJ+ufAP8lQcmbrkVX++1sz9J2xpGHizp2gxx4
apJR2GJBEPqzXvWM0KpNqFQOG4Qsak+DL2LOT6cnAq5OeTJY+Ilvq8e36ya7uBfl
IIIkX7x+wXPM8iF+gZUPQCdH8gIKa1gpyDAu7AVWarQZH5I5IoK/jtNos0WBMMYQ
kiO0WBoUWzqcqT64h+c9A5OxIIJdwVUWKcdcGR9NcpEXL7rO2nUNXJlZ4EipjOVJ
gWJeMVzJuH/90CwtqLsfuVIk7or0s368l1cKDFK+fwP9Y6p3g7iBE5lPXjK0CZbo
tCS6ltPOLE8bJMNHX3NaTaqRhR7DYSrl+0h/SVJoRoP+oR/yUtDMgcdTSo3HB8nO
YOGLKvax8ILn56t1fVyms5HH3UzmaDByfB7DhHneu5qonHZ4VMEFI3S/gqHEN4lh
f+UCAHetzlJwP39iC16/Dj1Hmyh9tkia7r+ddHOE+jcIM+5Fvnqy1uvBekhtbxHj
rW7XuSi5oJjTPHqXAp6+Xh7yU/s/eG8yvn0adnsB9v6HuVxCa+sMaaj14kH6Nqox
v/Xcppe2qtVoVNkxhQwMUqZY7Ne0gslIRTlXZEGyDQNgh8pluot6XXd+q386Q1BR
7fWk2Yb6DPKu0T6zJ7IDkIe+m5qeBDqFvOLvxW4ZlKDzlYkIz1jhuIEo5mWwVrHd
IN2HTZt4jccy+9RzuqQ7tKbBxiN7hbWPdRChQYBBEgey/TLtUeQq6E7QLAcKuGv4
EuYIkiM5E7KjhBX6/MBotT6KlITzJ0btclvWodrG1lPH8xFXYhHzvx9y61CnbIoA
fqZj7bT24I+0E2ddwbeiRiDpqgkW7Yek0aO7mp6zzYdzECeXwF6lrKtO7Aer7T7X
G63VOYrFCPOrVfoH97ewrrP32wWvmihgvcfDih1fOOCTPiDwtf1AVIiU6RjCwNwS
2QyoGVTtuiDKXaok6h1k767hwSMOPvCOo/KPzde292vU5ZIhA1Xx74GU4yNtGmMH
qKW44jn02n15s91RzSPENThRaaGJ2QRh+rWgL5Dc4Q8skl84vQ3O7B3K2BkRCUo2
ZSeese5ZCRUOkZkwTP/XNGdX6z35SDcRD2pGj4KmrIOAYWnkTNnJhir1scAVqsKD
hCIrNwUqpsRf9yBuC6pj899Rr8bS31uR2RTy0sd7AZdEaVwUPDkzelDkc+utm6Vv
V2m6GHVn+jMZScitkzRtUPOd53cxTHQRHpywYV+6PyoE7UfDhcdpFxXjMZrQKy5P
8sRJTgxmKfK+N3WuF9AkcdjJ51QJX50A/ZyrLK3gpUOp0abT1ZSaVoCN7Z4Sb0tD
GAPZ4Ajrnt7G9v25sSOD283xi5HA84+tYXyj1N/uvP4aVvwkuNt02LukKTfkKSOW
qMOcPG+qeWhqVAXFh6Lk3Yg9aEkMyb8hu327J7QYheZMLc00FcoxNYcxez5FLzbl
B0VEeROch/GvgVSNCs4SgVjUH8dFhfFy2XSf/JDiftoe5RR+96/D0l8hjiJfHbzu
3s0/7uMTH1H7IJl/SW35YNul6NhSci7wCksvA2dgMazl5P4cIZJYwueLrXykrV+y
poIw5BhOq0QCJiFwtHLLr+BO/yuqHwsjjivyaPzKUTFK0s+9kXeFTWxd/gGXo0zM
lY3aQoxn+Tx4URodFqiiSulTb4MS4XLaw0BwyHrTO/h0yiTCun31HhdYRaATUqJm
ySdk4xd3q8O7q5u+Q/dn6BCcNkSURbI+s1m+4ckqzLFlcNX7ITKUMQ1vBe+Ky1K3
LJ0whivHXFmfu43rKWASZM6BwuNqS3mRj3KmUFPmlKGnM/JiZ8UZDAddEt4ek4dx
EWrxUcOYT8RnfI7qPLuFa5inhBI7QUEFvEjwMYdcWoDVsvlTACNG/iGtSLZrE9pM
PD9iXVwzBmclpLNb9DBJLGT91xGPTUP4Ju41QLNCa0g+3vLzLxGX11zwnBGHYGl1
aXG9+KAD+UZtp1HZMGyIIdtzqLcRxFjD7Thgzy/qllMjiM4Zt9swqrdqVjz8RD1u
6Maj++t1AzZPm6w2wT36DCOnFbkgL1P6FEjJHV8dPlzs9du/tOTVK/YLsArSJ15D
LojEIMRMztoPx8BC8Kh8LiRiVa5FD/VC64oAdCwoMJ7aKu3fNySRBJlC/Hr0sF9N
w1MLB4RRxzJvxzKRWvPm4DWIi6DrNbkPA9xn0oyLjeeI5QLFwIjKG/6oO4oZMgoP
WfPPPL0pNom4GyFpl8aOqbPO3V70ccTLKL4jyyV9y4NwIurvYbq+AZDFvRDNLQo3
OwbUmAiKblrZJ90YSbt4g00j2cq7AavDXWlRpJpJWjly5DBbgmsAwy+tVYugn3C3
UUnCj8hkvH9hiYM/xe/JU4XBCpTKyhUT6yhvspGYcJWez80JVo+UiNZVqvLZO6/0
7Mm8VJ7QJOz4C6O64zWbLGwDMkQ3qtnD+bmLswcvEtr3L73HNBYI5KpMO8D+VXzA
DYhUozQFNrvlIvnWZ207nrek0HrdXo2mYphML+9oieFqW+CzYvWT1lk7fb9Nzui2
vnfLSYIwPd2JBP/m9+HuT3cPF5XbAj6NnHJ7B6MV5V/WNElM6Td6ArGsT9sO0a+M
MaJEx+dr9Mo7idJtAKdBZKZhblDLSv2yUvleIZdyPezQuLjun2rGIoYuN4GnhJoT
Nli1cpa82JQnrfxkeWM23naDUOBnAkQgoXqki1AOzVOH7cOcrhWuso9uoRkphIDQ
F0WAGhJtw4KVOZuso5i0NSot+B0pdW1eb3Pkl3wI1DCm07CYM87NHCkOjdyiTGr5
7muIU8MnGOKVp3RtercJEeyrn6oTZWICZsCn0kft+cIHoCl+aaqqZtY0Vme31vRc
9ESIig2kiu9boU0F9DvibJy4+diFwWmeCM8xeqneLD8LSBRKdhK8fyxuGTp5paF/
gtTCHV0P17zI+wqTb/yKWnWgnrozspIsIs2Qjg9A4IfFJ9cty1XPIMgzJM4NS+GX
LKz2VrmVlZuN7FRiKpz1DRA45xF5Ab22mduHsVVtZJWcm+USt0gGAyx14IR2lird
C8kv9o/I26nPn8QyaDnFTL0PMeF9BqI86z3GK/OEjJ9bjXOeB1hP1gcAKSYqTfxX
PwYptwj33dU69TT9+tWWeuqsXXJTxdwdrwycZa9zbLpgFFO70Ndid9SG3r0neOzL
wtPmXmhPIErxO2SRAWQepu3lcriTaIixVsOOWL1M5KSaH8Oe1IN7ygGYx/ugTjnQ
8eh+zV7SzTFBKtjQEiMF2TFzFz80jur1D7z2xkG2pGqExYc4b7gHsrm2lwixzSiG
JAPXVXJopK56Dtwyyct/m1vSr+76W4ifl7GwMKyMuy9ybttB4JjOnAxWY3Jhftax
Uotp90CHHHvjlfltEBW+8mQnhCUV1QNsGffe1CXNxcKKRvkrk/gnlrlsyAAA2bNO
d4EaDJ/9Ta05V7Nbk/NQXEYAPW7VA+hH4dCEjRFtphi6rJFoV+TPKqEYXjWbOGsn
yRiQ4mKdMXTRqfOxCOwN0BW2Lj1aEA8YxAjSeU1WH4nBhvRMZ6BIzcBGf75VtwI8
f4wCl1/Pn1hINDOiHpyl4yOAIBYSy2O1aNJYyq1+Mk0oQP0nHumtQOj8oNAHivsf
lmGdmKBSgDytDyzbYuGjX+e7LMBlAw3abGGdgWmjYeMY6janlSwwtfTo2400Te4X
zAzWmTI7zLAWJQqlOsY41xT6cnGuKaMM9q63tnywheinOM38rgDJGiCFUbPAB0ED
fKhTkBUJuiIdK86LxoXIeQPI8/R9rlPg8nReoLfVVKo7xMFLeLLCg+hTjyLdUIVZ
ImfokSDcMm1VEMCNW2oqi3pAyqWvPAmxv2jdjjnd/JD17CR6L22yiEhMGfoMK203
LhodmsyroUVXiRlpjBsaHQnDE/Fp31d6QFvjcMe7GoFwkHEx753tSb21W6+BEDbA
ATTCkTQ3KlvN7QpqboaWjf8wqD9XlDXd916q/1hiD5E2NqBwoUJeRcf6xbVSfu94
8tOjUENbn3djwujgGylU4i/PMMmSYmMDGX/WODUuJPeFoU+T735awu+lKZTCjOKA
qn1cYb1p0jcOh6e7eNGb0DrFiHUCfyVfMgg+z7A7uWk3opOtNfLZG/3ih+8W1Aju
WSz7vd7PM5NLVAsH/zdp2JT8Nzoq+8zQlVRHSX4MfmVD67LtLQu+HkrAc4iMlnNJ
yPfPYdk1owOEbM4NlWdjavfKW1N1sG8HEprX9OudViNz5bEliMUaoQVUAVIlyKBk
Mu0/Dh4eTGDblXIslvstjZMw2o2LCmzuCrGZlAJ6vxVnb+UY1A22DY7Er3YX/KtU
SrFjzlzF13R2men++Dm+WMDzZt9Wqma58xsTpJWZGyhcwXREeLiTHohEAFcm9+i/
5B88w/FINovAedTu31NCbZ4KH/d1xf21uoI8GIA8gLvePAXADBi+x2dM7yIP199r
Xi1A60OcoMuFU7LgXKPQ4X3RlyKdLsTQdDCQV+7BlE1Z3xj0n/1LByvYqhGJlbtD
Eb+XjPy86dI8HW0dys9g4Xsk/rjh/1RDe6scfXDc6kmfXGsr72snv3bLtbFP9kjo
KnPV4MjlJHDQB4cIzf9RaDqThqccxS2KEW3wHLIWvDnkPnf7AuC9j6QieYABPEpz
w97zN1Ez9ALhl6ZhA6Vsa2R6v7/eH+UKw39/KdX7Me8+CKaDrJ0twhsET+5sG9c2
p7uvQbtzpHXjXVUhl1cnreLjFOhmmyygOnz/vjbQYZEtd55iKV24Ah8vE1Y56g4u
50EG90kOTL8isunsRTJ47siC3/RDiZhxw17KorueANT2cUztE1gwv5WSJstYNXgT
hQqZ2ofaBeOXP8EOkt3keyN3mRMD9htPgcSyN+ii95sekl6Wgtz/TzKwNqpjCtPR
vyMMN1k8/V55ZgTg0gEWZEhHrooP8/uMV/noEx2PrRQMfZGnvUwJmZW3RB8zKu/d
MRJ8LTiGVYQe/m/DsvcLkbb8j65+l4XZvhPkVR3EO5V9vLTw8v9mJjrpxcV2tPGD
aClYhwNT4G0HeHv8R8iZD4hb+51tmPtrfoiCV5ftYs+YvlTWUaSDVLiwXBso4JeP
lAxC6e5275uqS0xdPk5VijHIoaNWSveimO+bkPu/x2MGKzBrBKy62xwPXCvBIlcP
az0VPHa1nM8oqjqjfy+2YAggXwC7lBD9CTe2+W5huelItlstksIDF7bA8dzi3IuA
SOnsuv4me2fffWBQxa3/QZf+y/jELhkS94QwuRRy4ZKgrZ3KCLsqokHxbkqojf64
Zi1VPpjz/3nTY9SZReNKnY4wROh+Va4VCD8phHqKa69mHcDjpCfLUsUd7wVEhPFi
X7XgSSa4TsqETVXpRlHUH2xlHaFXoOb7ayuNtNCX30n1u5IDGdPBfEqSwLWo0E3K
N+NRBReCabCiIC5EdQEuN1/huwgMlsZIIuamLa7D4EM8Eqg2p+rDZzfwm7VWZUpb
4xxIgGxv84b1x3ocR5MhMhxIED6+QXBvf0nyaxClCzhISH66LRW8DFpIQHpNtBS9
X/BsDtjNo0dsEgcUvfACSD3PeFCuKnp19HU0JBSrGDmmYixdNuRylimvsge5pifs
EtOyjHmxOWVmLpiralGelQ98LyIA/gUfLRE/g21tdVXxvVBgRYMf7wQmfDPKnkWq
g9HJehiVmmCTZYs8Hx4SDlK9sLUEUOEM716rCOfGjMIobRQgik3udWpciNPuc0X2
oB0H1KZzwJ8ZpA63pBl81c9SA/x0dLRmA81tZJ91g+RF6SvZcWTQrKgfreNskz+c
s9ZG/aGbq3nNEgjyu4vvxNVqokZJxpAntofi3J8CWOIx5rU0eix0QLdAnimrah5P
dCBfG3w+Vr1pmjAkPrtxYCgy8/Q3FtprU5W+/BrhAfe4e98cn4Rbvaz3v9eYBJC3
c7sl33PZ3mZfzugzetpE23QK/D3Zjdsg5EwPjaU4HACUIcdITUENV6ld96lHc6PG
Thaxvxcv4Le9EQqpqez44cNrYF2FIgdiGUDO5CnF4PXr+22ef52zab7YMJszHPYz
mgvP4HY/Oy3lA4YOV5eqBsPCQwdXDDPefCkjr0jfe4qAKgKyoiAp0uaVDyS9qFMy
buSObqEjsl5s5yyx/sy7SbaLGccfIRGDOVLcK9snfvRgp0gV16aQcWryWo/BXMwc
Z0/YWtJO6njmcFkOchlrf6tSoz77J7bQx5ebEPD/qGm3W+fwtRnvxewB0upvSzUs
p4/oPsCTG3tgBWGfsvMVynRsQkv8IulxgdVtK1mcrk7s3iEWjsX3f4GLSSP5ZxEV
nK60PfbrIrybIa/P9xnN8lFiPoFqiPLK5ryn0wqSkQwLBHehVGo8y9xZq5oyQ7GX
ccJ1zIk2SyzCPzZ3Grg4+qAhXJeo7mwcV9v2h7CnpAIjUssfwEjnrt+DUX+nKZ9/
QGAnYPpCkjLerXLCxYlWvK1ZcxD3gXkC2t3x4L0lKYDEGcK0mG2ukAC6Feo1cxY7
x5Y7fd6VdbTmu2go1MO0wArSVXuhwFgMe+dtyDqDuuDzK4eU2Z8Td6ao5QExwskZ
o1zPh7xd1D/gtR/J5AnlO37FVMgXAR+k/i6SwdWgtLAImmckDGz4O+CRQgvFfHcx
oE7lH35D+l407QsFQTJGetedgVKYv3F0MwrtSNOeEoaonPJlPX06+79Z/JpcC/0G
V4spaQ7L6J3M7IS0JKFSgVpk4kROw0m3fdbu7VtGtOm/A+aNw2hS2rFE5upkLY2D
wmLGFZ5xXq8sQBphB1lxISMwKWG3CqQFuSnAPMV1ApjHAClvwh67ehBz/4BIYttL
mebGudzOmozyL6cQZdIDjWZGbZB3vwd+F+BME2YcEKOsX0riGK0Q6Enjw+VuqWPH
Rp4LzNFq5bFWcQvOYHQbO10/14bJ4U32yl3Gd6mbUVmEyzoNdd6bVrwWbWObPdDg
ujKeqGMXgIZ4omNd6DmrNCBMdFFxIs0n1SQlTJ0ROCvrkrqyIke51OUzf8WLKtlj
mQ4RGGwF/vvXMzcH0rDRTJhjE+r4007P/XToseeT0GaMGrQ5DSqE990vudyNKVdb
lx0Ush5zHOiOD7Lzx6J1NxZ0gKPwqMO7vlPwtL9OJuZskbH3pC9mBFuo9t2b2gP7
NgfNUx2ZvtgUO8KNXuNs1lGrdTgmXnD3uv28+lukfPydLWjUgqKUfT0II01+ZtEK
5B9zfqYtlZN0g8Q6Ghs9TeZiwONrpIu5ZRgdsnrA5g7JFJqkgEUFIkzt68a/zvHQ
9QFnkgJGO4pAzwX30zqYqQ6p1Vj0My3/YcJqaC8wlS6XBvffrqm5NgFwt5j2NZ0G
yVzGvGyseEgOFBTSmWG1awQKuETa26NyZX13Php7bHQyVn8wez3haVtM8boj02Zb
P0MalufIGDdScABVVUKVmhXP8QqqTo1g+5aq2ZxgV7Yn4ndXc3MZahZCTIKoZNkO
VkrLPc9na5a5tyYC5SzofAltLQmosUfTfu7VxS/B4sldaBHZOJ4khX+PcPEWhGiB
EG0dVJXSk3Sqzf17i42lS42jEBKVnFrWGFBTIBQ5CNg0ziAv637M7lz5hXIbsyKL
uKam35onELKtbE1Ou9h/2zIGh+QRrY2Yie1BzsYGAx3dJDLtg/TWW/7rnUdEdxCd
MliYRx/27mPPX55r04hJ2+edEoy4Gb38IX6yIfNBe0rz4vAp7VvAzNCUizvL17cA
CTeq/ao2j78kjMLlVXbN3jDqOlQWPVAiICyL1mNDs58AdXgndjKHr5R9vtQkZKbV
77kkU0X9kvO7lz728FLR9+gEMYuc86boS2kzK4zV8zrTJ1M7xu5LjEQ0gaulF1aq
j8y8sCwcjfj6sWdboBuQzbUYb1JaLg6ZhF+kvjVQYLPvYBtOm4uWbyeudwYt8DlZ
WV+R4TfbY5l5iqN04mENPVXNM6ZRepp7Naxb5921bfWCxG8nz6wB6JhRKXwBRMAb
qWmFiAiN0BDZzCqu08MQibJEFeafUjrm1cnTMxOV81YeunCt9v1oTdojObwM45nm
WBkIgvcDEffMCCjKyDwJl3Dkqx9wxMwtIahvLjDN9ijfMob6vczT1pYIPRE2YnK4
xpC8Qn3iZBvkFKPxOpuatvhYTzWnkGsl3G6yN+Eam1NgxwmetPkV4lTOm+bXcCYd
bEegUq4rtNOK/Vu5IZjoLT+iOhdvCxmB/KD3VuHZ7JHQPbFoh56oBELqSoZ7AZd5
y8PyCztvaznD70qJEt47qRzYudYctiVhz9gh9VLg+Pj5bm8nvCoxqAW9P0+07IUM
dDc92wScNB2asHaIc/zH3oMNCuePp5So0zx1+AEyJT30Oe3sfXr4wedRDd9qxnKb
JN1kRIon90UJhuGpG5GvWM3Je5DeE/U1TDyLT8mY5CT/APRv92SC9xmTAz7SIzr4
1FgxEd6XyPqAlEE3wculllIreQYI8L3lnX7IxkVfW7q6KQRwQeJiPK+p/X5dJnIq
0PjQ4pJo6o/gqIPbNqe3a+PSx3lH6GTIEUcYESdbDSUoWCPqq+i+phlfVuSGfQTr
+JLfhIvreA5i/ghfLGgYhOGEU1rM6hEoxqOhUuspvneFIo1gT5MCr6j6d8hlhUqn
fCI8b7Gkq7elXqwKhExPLxEXz6j2X4Pm+NxXPeBNYw55uSzWSTuzZVYr6oxu9B83
l4Pj5P1lMye2mqMMIgn0HzJli7kULGhHgBhdi/BQo/RmeXEyepGJ4bBg/mjfLB4z
Y06vXpMTAnUbEN+14jAefIesWHm8T5Pp2kg0uFFScWaOx6/bVhWnJRgZV8fSentU
cFGnozlj+2ZA8YQF+Wp1jgb0tJGJOM6F55PdYVkJHDye0o4+uZbOAx9hqQOmrkDM
pqeDgK/zOA1AZYhFrVmGCdpJA5tiIwupzBSO8J8xUrMI6NLbxtMFv3+U1orTtZx2
YMGa5QRuyeTGylkHkKDoUS7R0s5ZexnBV0YnccjF/IJ2It4u3IgiiACZKIJLy72l
h4gxFtS6vaOmRsLLsi5bC7PSPKGNH/PJA4fkuIXndTeXiMGlIk6gfkzOAccxn4nw
ovtzQ4Bxoqk7nmm506lMFBg+bo6xGX7Ce9FxxPUiWI7Qza60l1hEldkM2G0dLYfG
xUteobFfudCzvzNoIpyr+lN/kxjE9BGt4rFwhPMO7l6SVcvcvS3mYpGKYGADKxCw
d4X2w2SVfamE5o8tAA3Sk27aPgF1s1MwwvqLlCD4XLPhQhKdmlvn9DpiHK6PBuJ7
y8/Or89TnCcoOBF2ogjppCvmUFDwEEjmqFeJp/EaawNGlP+IlKAU+ExtwdUHHNlH
f5NVjk5AEY0wFtqQ1rOFsvCn7o/ZPQ4vGHPza2ukrB549NENk5fe2y5eXn591TW9
WUa/cQM4aNQl14GEnacKwwOxQE1LjqalYG1zG2/JCOQO2u6EU/DcrLwf+TRduOoW
pEd9ZzyiSK+e+yM4fg1lYD+VA0voi4VE1zrzVMEz82MUJ7EXMcwKriRxvbgEIaRm
FRpa59omCnB33kIn7RemdUfn02ajlDIf24l2MGcJgec/Sit0EMJqJ8J0Czcl5H0B
6tWg6KaAcTFV5w7NPZrFKe+8MePPM5jDWaADODt1jZue18ZwshmBqa/t/zNCA0xt
CUQckV2R9gGYOGEpzP21cabtcHlfuoBHACR8qf5esN90+OX+8qlYE1WBKCTG0GV+
xBPo77t339+P6d5RnM6PIVGuevQaFMxjzMR1dN9XqK1xj2UUZ/xn791QXSRK81G8
gJ6zc0o/t9Kwz65Hg+grtKIWZLYt+pwND5hDmHIOFipQl4BpBtS8gcIjut5X6GEx
m6dm52tyGqtDioiPAXHEWAdLhDHxdas3X5XnZmBQFpzoFTDQSTG0mFr7WKqJERPu
9VwaMnQrNzIB+lXE3WSegpU1WJCmth9fcqOorpm9gYdi+kN+/QH5vhNRT2qNYiTj
RBQ+T6lzjg+LypDb6O/VyuuZzlQmgrlVlQjMUFVCmmH+ClNZh5atBPFIjD4ToZtm
o8oGCa2Tq4I8PcqLcnKvKuX5B5OdPkV56dyr6MvU8/M5QeQn7MskqEyM5hSzbkBs
PYigDqFhuS+eO3219f0sSnhr18DM/wCzHAa/oAcDOdmdHZzHdliXCtdoON7Njb69
DdawsA8/fk3+ObCXwWw8YNPoA5VBtXz6XW2oJ3TPXioJ6mIgqQi/PfxORVIrRlGQ
LqHRe3YqfC/38ie1Jrw8KyaxlgZGkwRu6NBHofHWa/ObUPXUaltiYHpJrmgCGJDH
oTvMewawRHNBcVkdeQDz2DwMnVJ1ygASSrkKMofaFwujA8817aMHW907HUJYeHfT
UAHU3GVmRM6R/43a/b3yIX1VW4SaLpZdtphUuk9cVW++0ix71F4LewJ65v+75lwS
qSwI9v68uAvuOGy6+vVA+zX/LAbLEJNkDH/sa6075syijKmLgX3rYRkVpEvNJjEN
FnABAE6wRfjTEcBMXYC2HF6o9+7RKloDHtQfsCpbMvk8YpBECxJggD6hJ1yd42te
2FQPrsw9jAKnX7/mOBD4o1jcaXB58LL/wrD6pgEB0wEN/NV2o6/WspB6DBEcSL4c
KagT+z6DKJh9KesbKfepr8ECksXBQpw5wizTK5bOI3DAuaZxWrnWmJMa8mQLgOHX
kHN0HoUUA4N8ieLN9EvlLNtHEttYgmqdzxkrVS/7dTWygMBjuj/AQAq7aaRNGsHG
IwC+wAXlsTM7MT9Cs+LJimwqLosKiJ5M+7lqMYfbiX6SK7ddlrlfNQ/MkhI0XOyI
KnFSfGWRc0TZCCBaxKl52DjjzIVAdMY7bzq6jLqcJVXbZzk9+zixXIXAh5IOlE16
ec4xvlAH0rwUGsmSkhTCaZ51rc+ljBaMdvDmgfIB09exwCpND4Ch/HLL+4S19WXc
5Ix2/0k7l7FMEAaWO+CMMPZsmALSpDqs1RGL8F6oD70u249Cvqzniq1XN5948v2W
o7b5j298wx3jsfgQMa9qTYi37cQfylABgIES5BBaYbRP8Y7LGJYofpO6CQ/4ZkZ+
J1WGsHttlq/XDGvuSDd641F0Ht4TiPL6arD7S0siJLVWVCT94uV5/gHUIUVJx5c+
oz9LKflnAoCO9c8o/5bNThWOtZYLGY5JMgmDIb17ovCNmKWl5AdRX8J0XG9lrxTT
M6Zi/v4+4CxJp/TVPE17bmdh1jXvXYMuEInBb4Zu7vkpgl2EhEx3Viw1RtrgwfqF
3mZe8dBPjA4zuLoWAxbIKGgGCS7E0D7he3eZ739kintRjB3dYDMn+YabMmdM5psd
58qa8cZTS4fkZpjG6WTy+9vsuPMLuQgd44RvPeNpyBe2AK6bEDBWnSURv2xbmisy
xLTfOjwK/SfN4yGhfqbn0N4ZZezVRa+0OVozxTHrouuQhWIBmkqll0535CJZzdBB
8XYu0Iq55J/4yH/dM0Zy+K788sTViOZ77EhVZ0i6He9kSuBtdUWRdVM2gLGJ6WzE
l0P9J3khm9YjlDw/0vjwW4L++NWoiHKcS9UfP1rI1dEY09n6+2qgU7gk47EPdG+s
8ljxDKBnwTk4QV2tGfEQrj/xQ5b+fAaHuDbx9/MAP5OmPQAnvNaXThvPIDSTFw+/
6o4brj/S76gAa/QbcOXfEWI9Ec2n7VqSMJSyS5x8tuOdpkxRAPJkvXxz7cBtEdYE
kqIDLMNByxXVF5gpxI1vAqkdHuXQgNW5JoX9TAQeaDMWwvfdPb1aw7BOQm1kBiYD
8jc5GQbNhNWdFePpcbDsqFJKxghCwoTImOobozCDWuZizMtgtL9w/2pQMTq/BLsW
x7lcthAUnTeV9nMN5BYvh+aAyVEkn60RuLcfcpvechImu+nUdO6pFhRgGbQ3b6qq
ezj6dXO2Zsn69iEVnP+x3CbUpzBW0ODjYoTx5ZbqyyGTLJPuyVyi1lE2TQgUt0pq
dqnsEsCfr3QmybxKl7h4/Sj5uev278iR9YcTZKnyDnnrYb+AeCip89EAgN/ta4Q4
D9YkVrvVobN2YQiS1mnleYoaK9wXNaWSDGQNFLYGsO2exG7agbqjl+IjXWPMXTb8
ZdveZncUd5h11WPPbfwSHHmEl5o2FDRSQnh0AKIaIRwK3ko/TVQeyBCcPWWYfz4I
Yj5C8DoAzsnFCMROX8yW7OdXkcqvK2id8GU/R+XPLyBjmT8CzOkcpr89A0CVC63A
jlRHoT6OHWCYVQvh6RAk7HW6xntnwei2wBRZwuH6gyC8Tq48WQM+q4V2w7gN44/T
xgHK8WpyPCqYwyy/fQv3njbLQdf2cbJKU2ZSqw444fM4Xmx4rEl2uItdXj+5sJF5
KQXY1/5li3Ta04iXja2IQkVK+Us7lx3lLCoVcr+zMDxG4M9v7KGlFmq7CohRUWoJ
DCJ9iJBOjhrKEbJXPFj4f3WlpZVc8BAbJavt8SLd1l5Z+BGfP/2EyFLRLO3Yj9nT
Vm1iwO39AN56YXHECQg8xpqIvhjddmHmFVxHfkvy+y/+8xLlfgd3fVZreGkWDj8K
nDmmvCAbxJcTmj2VEJyFdaB2v+OoDozQ5vudkzP0dd+fHZiOJ6lNf/Ez1owdULUe
Y5k9+rGz/YtIutFDVgcXRur852wZO2PG2Jx5XftpAqaxKKEwCxrpb6/u6mho6Oxz
sjCex+l1dwvmC6kY8UPOnJJO7GjAa/kJJjs0tbShscQG2iARiKFHHCoGeZ6c8A/C
rFClnkXWNoLmfgpYQXTOjRSkK+vDLJMsMkN07+ir3H0OfKoEn++wt75ihkRYNR7n
Y4Km/5V+IJ9ZpE+BzHxwl9vsTab+epgyPi+3Ty326eLx6jx64qyfmKB4wGbCCrhb
Ty9olKW8SwjjfZGSZuiVyeaHDHZg/aHtmhFD8TiDpE9xgcA/zsKhfGcaRgbDI1PG
sgZytvA4gtlHxiLgQjF1z1chhBwaKS6rGXAEJfJzbczkWsqXGAiXq7Vf91av92wc
m+VDkbldptIFVcB2PIl8CYaVTEsy5qhOk/3UFd/B4O9SkawiqZj/E9yXhsCtQWUh
SyILpz0WKgf5kbSn3lhiRCeGMF/DtqiIwcuPGskaVYcnT5ybBvMcyGxgLRUv+mUg
HELKcFgdcVQbXfSCVNL12eANOFMT3AHfpos6mK5Xmm4zCVA7aCCogd0zsgCd+tqi
/iGdPKGLPhSGihKo3VaXEKgj9sq/9EkJgegqNQQqfr29wwaMc5GvgF4g4XcA2h1T
vTknQDFd2S9G2Rt1fTPUYYZACtRdkugxEt0SFhdaQPA1I/YAR/1QAy9FwJlU9chi
OI7cFMLaY2jSvx7GjWAjDEEMb44DWZp8exK5C6MlyzL3oK3lKNRbVJD4H0tadU0S
fSYztBvuBN+I5yMVGysLVqcHoKOsC7ODGLQGFQrkGDJR4B/7oipj//+7xDzb9Lm+
lQqr7kZUmtkX2Xx4UuDLtB00akd+Z7SUPgKtPLi0BAnGki6oo5/fu+74Hck1uvnW
Q+lL08houzXuvtpUfkz2kuVgGUvx7O4IexELD88oSpdtR8LUSIXq5TgCK9mZI1ca
Qw5hqIM8x7zf3dvDbaxSfTbUu/zIYn5Ut86wvJY2ljBORkoP+8hqYMYkqEH+yrMg
jMx8i01K3SXUMlaUIKlxaU/HDM6upGqivQLg3JXZpT1gOdPDE/8jm0uUnJtgt8Ng
9PyhCobwd9zBqKtzJahRpkcl1iFTsCftPTp9ZYs4LH7H1yxSqe2sqdTHVD4+w06R
Ru1yVI+PO28OT8xae4+q1CWhZjAhhE1XrtcWtYeWTVy85Acx1mNWJqW5pqtq1aXz
l8qMMBxVf+TAsefeHMKS+5r1Mc7CnLNPI4NEkuRo6fpd0itVAFS2/WkpU7Gemk1G
VOHhj3RpFXXqULdqSQOOSvJ0h3BHZsclsjvS8/yTedENpj4lCw5CrVSFLBI7+YUt
3VgAOFFCGSLtsRAr9adMVH4vN7x/5F+GnbRObHnLskEbqeXxbXm3hRcNZcdJl3GZ
PPXSoNgpQzpLlZIf8/Rwkr9Z7qKXlu4eVlZlu5DODA1lnszSIcZdgtrK0hRYRL14
skO6FGeJIZVtBPgxKdMZwLwjrOqEkk3XDHHDlX3Q4WAM/VJcSVo17pMBDlY+E75M
Vq0l1CzShkj74oVHRHviNkC+im/KyWOhiuBo2CmrwAOL3I7XKVjOIarf5PiYyovF
tLAArNPj4omcSOVfdGd+7h8YJPCbReZS/1IpGXadyBLEX1qtoJGixa7+LZj68RmR
6gawlt9sUp0qo4KQFxRu2XAI1pkloUevj4pS5bDa6JeP3mFV6zyoXcGzChI2IRiA
tQncM8XFI3vYrg5MP+M1sEnDI27p4rl1wJUGHsNnE0hrkwwmj++WC8VyebyngjPV
aEzENTIU2fqmYJPDprDI94p2UEB3UdojOzP1u9kkEOwz4/l0XNM2TJJNSo7ILCMY
CFZZTuF/VbFhMZZgYIj2UvuPjzFw2SAzK58zkPmVCePIjDwaL+APCprMaFvi1Lco
NbzflLMQ5T4QxxsheEZvE2usC723K3wzimusQDoda3mNFpm9nby1HUDmdHKyTQUb
B+2oT02BphTgzPKwcoO3XwC51uXBghrLAUdetLEt2jV3iQDlfF3Vnz5qiFnjp/+Y
YoBNGVvrqOBaAz1J7hQMnCBlzzaGfbtpTJENAWJ+pjPfbA0jQGDAkIhsqdZNUeYI
JT68kn0TGYJ9enI1obqubIcshOMfL+ACbX2s48Cslj8dDIMdr8nBS8yMC5pm044j
f/LBWrhGgmwM4nv5KwcH9GzAm3XEsu5OdjZketk+3nQ1KK12c6mQUIJXrGdq26Vo
a6Feql5QtQYncksr4AukaCbcXQx7R95/y3OgOWfe+PjYtb7KCMsz3yv2fn32YNHj
1gLHfCiq5774V+q68wWuACS1oHfXjeZPFhOQIyw5aiLZ+ec3T0CxwhYsUlA+cTC4
+XnNB371yY7UF1brnmeJAjMBniVBB8zNhK53uAzeN4NHaMW4dX8MatHkALx/TFjO
1Stmefg+vcg/xFRASI9RPDiNkuAFC5yGllEzCejOSe7YCcZx3QaDcrJsneh9y1fi
aBrtYmhyB5abqw2NjzSxaC1KLPRQmZmOwrUSd7DaWbcp8xzSgc4K8wfka9CblesN
PPDefEpw3a7xMaevr2s5zn6sdI7nD3IP1MY8XXw3IA7ofuLh/6bQB+q5HLfA+7zo
hNGIpYMuorjUyCmB1S9ksIrGbfSDXx8mR+zfOIqiOswmKtIYfzBkxmRsa1VG3cNc
nrAs8pFKeI2AYapyqvt2HXm7wH6ste/7ku69vrhRjrCVtWKDVp1D+w93ijUYqqjt
TJKB8WWYVv8cq0XBNT1bNxI+7KzUGX/jF3nWbJtk+mG1BwjxHWntX91+ygTtETzL
WCHfFBXFAfgN95q9J2/DBOCbVvttuKOLINVW60lpTpoT+z+v4SMu+aC160mvFKN3
DwVZkPtT2rDhW2CRkCgmh1ul1Yxa0C7TdbPxWxUahG/FRvn6wYzPTZQhH5skdNzN
W5hChpre3D1aPvc34mhkmOWkO3OFOQ7UIwjhT2Bh614gokSpmVQatodB060UYLZ3
K+cHycq+wn2cGORrZ9q1LCFGLatpM51KJRiyT0kKjwJLZdGcuVai8ESNVashxVoU
4aZ2phpvegwTuyc8jBYFKl0kXUCpYaQrUhZcSSBfQjX4nFmSTAbev+sgt9xp0oLV
z3wUbGkEsOqzvgVgya0UFbBMSSjlnICl9Igmi7Uh3jypS51yvY61EdtyWzaXnlKo
ic2+fm/xayVasrXaULO+pVhhKC50gYCC6Bg/afanoaQBIG/oCawi8SsrhPK+KAlb
i52l9e7fiCxEaeQcSlBb++grQZtS5xnUbUe1KpNkK8JCeU1WC4YO/YodslFiqk6T
ZYC8+4wjEBx7qi8zaq613awptMxzOtm+EvrGvyH6GecfCfSFqL3SLFgPsc6tCKrw
psPKpK3TuwdEyapPq3cooX4DbYfNB4RC4K0zdg90wbgcDwZA5ZRO9cTD79F1GYRf
4/szWcWNPzvMr48o8KJcyW2if5IB0nVpom7Nu/PB8SvipyJqPPRoPYx6ekM12vPn
iFEbcaABvmjZZbrtSGU66pM3wJ+z4U3mLEbFPqrQq9GP9upSYIla3yUKHhdQearh
qDczjnqFVlX6B6GM9wybTqbNlqyDtHO6IdzlBvm4usEB2RKJ4mOn5k1KceYzU3fm
Sda8C8WLxtZ9NiRnDKvjJKR+fB1Ca9s0rJ0VW12FpA/L/GqdJPx7hfKr20QA9CA2
MjCRn6dAFkJnpca+uoJrWWqQLUngihhbXY0japLxmSJD6kDvkYhPRzbp3NlNyV9F
6x9nIvtbsJsVRxixxGLLttTelj0yBsR95KRAMum1n7HUMByv+LPpDQuKawPnEzaW
7AMRLNL9qGUnrWU9krBd40LDA4b6Bv9Aw3YbcCKik1LJS9oX2DhChbldL4RDhbvn
ertMF7voKtU5nTB6QM2Fq16Kc4lUaq2Zh3EF1DWmhGdEoWO19ztLZaA6ciq13c2Q
ivMo8FKSHR7O/UCWm+91oiZMjk1OeN4/h5l3RotkPt+d7IfZ8S1aWMM0fVcDdphC
OhD0Y5gHBWuXOeAif3YL3nfO8LZjqz2MPdja/gS4xLCnoSZkhNxC2qFh4P1dw9dU
zYqmCwj/oPNbHWp1ArZst7yw4u8E94t/cYXOSxLNN+x8Qe9zaCg2IMkXfho1FtYr
muP/nBJX61u4eOrE45ooMB50fnw13pOQELXDHnYcK6PNN/KLQW11opAMAfnM8CmO
6gmYWd3OHz3w15JWYaf6GuRB2DaT+nouSMVNXNrfNq6dLMnRR12n4MI54t9jB6JH
ydaC1LtzdBmc3u9axF5CRyn8kegf9hF0e/Maoxc5WlaARMV8mhnhaDDJwne9SCUY
lwlaqV5TlJuLQUrh2GhjBRHWrqrkICAq9siyW67e8B4WbCNhb3i3XHhh1TN+fR8P
MWwn6J98shhrykQtUNcZCZoedN3PC56hDYbzi/2nC4TrheWcvPmrexM2y8rzAh2l
Nxu2r1EGOIzDa4G91ch+sAoS9K6kH22h8ziqf+FhUx6ssk2/8pUIgYK2d3p8xZHh
ie83AGhHioaLXUv16TPJvzFzqrQ1d1H+e765tGo4q5lT+CRe1bOxH4Fjcnp2w7Pc
MTmzleYfY2FLVA6KFhsfFgbatsWeTzzS2Zr4fj5zK3LOILSwmv2OGjPQ6RK3tbw/
QtCs1aWMOzy8lWygAGv98OMkaf0h7DqxlZTGbcgCLYLpjg1OUynj6BGGh+3Wmci2
chFRD/RRlcJvN6rS2ycatMYWSOwN09obATI6kZvb/K/YFiHPDYurifDQkQyZL+dd
Y9PUerqmFRZUCFOdw4fLqB+xvnTqDTVSGLB6No72mAR/I5eMDuNsSeotVTKOQi6D
RVyZq6PV6vgPLKUaPEACTKX84XEOsuwrbWb+pnHq3eDRmOrRGOf6hyiIHr19LGV/
x+VHnCgWmnMhJUmKayyC31yQu/FgLK/pI+W7uP7d5B32RE+rgdRNEUvzn3cU8lpW
btbW0zV8xH4Y9HVqAVwvHR3eS4VxswtzCEffUuSYRDWQIBfy0i4aIvWlpPQrhpeV
Ew+GEXT59JBAxOhDk4Ko5+UPz5b/i/2im/5MzylBahJix2Zte2alpqjbJm0hSqch
FqauaZYXc/I4Ug3c0EOxUjQ8jqBT2x3rQSteMK5fbP2c+iS54efAMilgjy7K67K/
gGDygQ9a9ynVjxZ7ktSExaJNak4jCRv71orU4o3tAFD2DSG6iMkZdAC2PxC2WCGM
eooPSTUHiB8qgBNZHBxUMVLuzD4IWmmmuV8rNbXXQBbMhX9d5KHqxrNi0wgVX148
UF/3AKzhRZgd9A/PH2xRxBGdnTBg6eKYgQ8YcjLcnw9uMjI1UYsRLHFrS3s10oCF
8f5sSOfjdfdhqeDoGY1DRRgRfopPOwl3KgZ+FWLVuCdgK3OlAo5IHYpMvLpyq8Yl
5iV0WM2QCa0fmtfa0fTkXM/yX/7jqamQryaX9lFKf0uOPmwzeVC+I2hQdRxDdXd9
E3zG+YSyoNI7W9h1jt+iehjusypvxLN92Juxqhcbu8DvbwwpeAc6/MLH+8MBeYsh
ilepqmVq0A0940g3P35xgR3UymeqzCIJ3iwRQ1e9jalslUoqckrrBvhDb67qbHCu
fFOb9O1saHLdfk1aSRRbmdZNKYsqX6VVP5/7THu/IQqwKNdUF5XEPENA/uBXRnnY
2SkGCb2QbGyPrZsE+6gN91qHYys80Irxe4RGegq53f46NYZus1BSg0dHQjC8xuw+
++pNICUeHAmwEdD+4DykiJHQEFYbknmPPr9qd19Q8yxROWBJPVdh129WrajQ9oHU
PmnoL+du3dehmiHhLAwIaBDBWCePXWFjmpuxa9+cM36CYfHWaX5tw4OagHbbjkQb
U3CTLn+OR1DUrvE0Z2CpqEVBrL8qe8z6s3gYNyEjgrcOst8C1angtjdrcWd/qbD5
cYofDZGq9lYV3txwVfzIWsQxBYQbkeQH/Q1YEEX/0GevgkqzC1jHGOqNT+kHB8VS
1RfpHvkYvxyQUbUsc+f3wqWvxycth1hffQ4eJGRCyLbJ7YzqGp2qtG1X8+EfwGhL
J8LhMd4suZCVE8mJA3FmnUKn8Or7RI4albhDSVC3fS5zhp78gyJedAGxa1Z6BmqT
/7Hmnt0uduXrB5thLaBSIkWTRHa18CXfLUofFXzEs5VjmRpr7V1e75KTjhQfQdcC
1qkPZLtXLP87gaMhOTmQoAA1J68/LSykIANRXXwwvn6yFOM3r99IE2q7fezXPhgZ
k0lTwv7oLrBgu2ypZIc8gQ+oGLyArSSbZydUAlG9IIGvGJ+5y4MY5fYdnOzBMq2R
vX5aBPbOaAh9gfNPZEqRBezk5rhYfXN1jGTSIRK45y1T2Fa2aBfs3OIW9+hPKYnp
Mff++GMsvE2Q2wIftAiXvMYQVREWqht3Ds60W7rMVmjpr/XSQuneXSJrkMBDC4cS
M9tQBo2qBD/8XUEyr+Zy4W2SqrfQXfNTTUpHR/FuxjI8wR4mTIbbR/Qr5TXLeY1p
4J4IaYVMvrsN/H8urcwbwZAh05418X7+NakU7TeZQ43m4BXjGPwa0ejDP6B9+Vp4
2ONCtTxiI3VjddXKKCol24TY3ay4Oj8JzVM6arDTV6vFJww9EtA2y2n0T3QwgM2+
xqcEQM0yUa0jNPfX9ue3d7TmoQQz30RK13/CEF3jVR7u9Cu/WLedkKMPfax4LHep
Ce3Eud2fGuKv1wK5+VsCPwODZ1xADJvyBBlplHdJ4Iv6G91oBTi5ZoM6ie7c6i3t
2QcTrH/4naeYCDWc+27ZrLiOwpXQtf9MSgJvsEbwK7e6u9fJfW4SHZ3rg5lwPpxV
7yOL9qeVjrFbiemkodSfTNrI4G5Fwk8VQZagwxJW0dn6Hi6fhjPy4LKmrCZEaBuJ
JSYluJFVKGBAPyy87SbwNXuMZlBYiOOTVTE6dKKJA5Lhn5oRXHOlnbymxfcsxokZ
rMNs0yjesJvcQi8gMvN5oN7FyD8ZNUUsOWCN3V4JuSfgZQPoeKDI9McRWNVVaiuO
EQJg8lmQ3oLcb+Pe6+rItY4DkXvygg0Uaogrg18qkZM23ixMCRg6sJ3dsVXlrcI6
gv5y9xLMetm/Wkj/HED4fczAGnJTAktCMWP7wtVIsBWkBt/y7m5mzh3l4QfeiHXj
3rek0tlUtKPePCO2HXoLZPtsqmRybSvCfuo9NFUxdv2XeA/glHMCJVZIQfUWAPGn
Oe2vX+h5LZ5aziL2wemBpjYzHZkJ0kvueS1RdkxcGYf5k5HRYAw3fkTB3dNHw7tM
pDqNBlVRUGD59CnHd50lEt0IqDo0LHVoGj8ZwFBm1oNpUPZkTc3ghsqtjehiTXRV
pOUc1Dyl4CMvEm+zudMIw/ar3GB1+oXH0Nq2W4nUGz9qjgR4imW1Sg0LEEeYFf2o
U9CmZWZ9332VY+8WraTsQ8FpMOL6JooAtVUMxXkSmiJy75Rcy1GLncF06TDDs5GP
O4JRLuXrrIU27e5Pn/mhDsz7Pp+DBP/9/9q5P8ueJS98BkqYzINyVxPaWB7xJuIY
iqHwgZ9ToSfc5ONqyPd/L3f5Dnot7aOA5paSkDOYpa99TDkXOulZvYNka1+gNUT0
IWmeqVucEs5WVUgF3RK4fUBiAf4nLCRCUGb9J9tVU3LM0LcNx0mYUPUCB6wW34sr
YAUk0e8gMvfx6pLGDQlc/NomR1duzYl5O21ySSPlOtfN7Pa7HrrzRSAeuyC0NEAL
oBj1fEvZB2qBb5l+n8XsbhQ/zbEzUnoMOor2wAM5dRtI9hTqGHxyY9V4pweMu7Dn
lZ/ZbLQYvblDGX4xlE5rHyuzaWW6z2CxorYk+QNuzvscNHpWBXLY1C1gI7F5WOJJ
qR48HjLLGiz8cFvURyWIcePC/Eh8ISVVKHtxWOKi40KlPcZP3lRvSKgbg8dbGjtf
f++yLGSqRbtqwgi/zculcRdGbcZofczZIqDqzuUFImOE6FL/DVvEptMc9SuZ5We3
tC8A6oDbszpHJDj3twuzq2PhNgR00Ap/zWRVVDG0sCwyxYNjwRdpEfPNQfsIKqlD
OtvFCpv6U9OyXr+zbcv+gz487gHVvxgsrcW9XELecjPDSfndTzhy3XO3j3qcpTwH
CkilRVl0yDXfpF8kK24LCA8tCzdwfO6DCvl1GggOWiIaJEHSk7E03aUM7lwyomto
jVoe0rK3UZLnebUZ8TBEs2OycfEjcJkAi5vUazxlvax4s24RTeS+52xUHUugsc6r
vwBFsldlZ5SQ7DyYKc1RujZF81KlM4OBeUMy/Lej329rItap7bMdVSkv9CILxF9x
i+8OreX3hdPMwbbz531+vtHO0LO30VLB255Lv+eNmCdKfwHHImptOKYnjrQXAGhL
fNXdGurFWKiwMbktbGcpSUY0Hr7AkvZD3h+48gqS/+w+hlXbQI/wpIYhMoZIte+2
3RkvDaCZgbrWjDNm9bEGxjz4KqumuLp6IPWaltNF+3E/fOtPplukslLpqTVO3q9y
l7WeiQZ2nD3+tVbFUazY6Q/bbBii7MIB9SeXq6BsWkrKYvYma8hEv3DeOmDmSycz
6FGsUsjzVpGQM2BnZtztN8A//ay6vpmWqDQv+U4xZSJJwwL4D5mxfnUaiu7Ioxd3
tnA0eErQkw7GrkqV+vJSU4rl/UjG9Y9rumWjX3e7YADRrbv/K1yPi3ZIk0oMlOeU
1nxiTUvEsw+mC8mZIBM/Pmw8ahtx86bRbOWtu/VL/3UpiUIa9etYqb2ue+FW+rlH
raAj19uMNNIru418NtMHupg64Zpzo8HHFI+6FqXwJ78IWdWuunB6OA5oMuRtJN7m
ZmodOH5GpOtmqGfsCjxGiGCK9i14dxrrDpwDXvnzkmJd60uPMBSIhplUd0pTngPf
7D9iB3NziOJqI+o50RsBjDHVp2DdDC2Ef3XMlnGdcjE+YUba5chHaMD/iwgmv1Q7
NVOVFMoMAg8L7sw/NkxfR5a0BIvzkkTFbxp2Ihobx0+wBgK35zd3RO1LBZXoJG2w
mNLOyWyFHzzNlCntzVJ3Jc0Vvn3ON2rBTt+XIQrD1s3KBJrlxEgoEtftnhTGEAF2
ZY+kG99W/N2q2v/dFAhpn7EEDxGZx19bK6qyLuM+uTJZOIOk7cG2eQfwdx0104tC
JS0Q3aMbOtrVYtHA35J9HQN/fcKh2fm0PLrgKFAMu7tTPePZLrsTdL8fpwS53DDG
ATJpVO0O8DyUWae/kAV4cBRWgcd8sxLgiVvYOideZIBEaQHIk04RWvrezhTsHD1/
R/G29aBdGmT5OVBa3GjcURCYV4bpYpWIOx2Ha68DYn6ob3dNRIo9/VuRUbLog0Wm
8bVAANXikfmmdxb6oEoFqjgwDDEfJzDbeyqrBFxigN7rLgjdz9wHwy0a1NR5ffuP
GMEqCPpKsE0xmD9T0JQ4TIuwwzjJu8IueDa+9/RqlmxfFhTktxr9KKGG4sE8qwsT
Wp6WQc34TUMVD5rw9zhwJL/3D1OTmp0WZuRNMfsFjccBceMGGxar/rdzvza0q/v5
w6dvTFOx7xUnlAivp9caEoMjruuftqvlypot16P5Oc3AcSD/wHKgm90UlwMEayip
bz7vKXD6SnjjvV0X7EPadmZ6kba7sDX1EY/71HgAMdDAbJN5gQqWA/asnHMQocT4
Bz+ac33lAlOamaL98qJbE1nnDuA61zQsO+k9KndAiQ8TuvY6XFSC1JQa9AiV63tn
t4DvuvIiQBkMjQRMQNEahvCjAvQUCK2Zjri6ej8YxnChG1iikNAXf+cjS2MRnaBb
jPGQ3VQr1mPqwtrlLPzh+ljZ1C4oKJMmHaVx1XUmZt2+Jo1xUaFO3B3+83OuJXtj
fFABNht1gehb4+KcCmqLJ8f7VinqEvniNuWtMQwxq08RfADAgk0nbnqv7zmEOmlS
Soa/tzb0a/02MnGj5n0ptsJimCbzu58MXaThUBKoYB1DQR2SSHhBP4e4oHB8nhp7
XxCVy1mufD+aVevAflTh/ajN0RMhr8KkvGPbCK/rb3NeCzeMad8GbTpzWdOf+J7b
vNfhveNQH1gjZ4DPUwdGDTGPhRSF+IFSnSE8yynruL2UnW1ZyD9ELvNVjER97qKO
u0Kez5ma2P6AtzGzzLBNTo3yVJnmvd3o4hMMuOisFtf6crD62+LyMP0JdK4fG4C4
vCeo/2IFvypGVlQw0i1kYxR56T5TJjQVt9KjEoUnfktnIzhVV6S+pN2F2qUAdMbG
hCvg/5AkVNT5XQys0gxcTaz7+dhsIoXkGXWxaA+9JIe84rsy+TyjBrlc7156O29o
uUGUF7778gcDzELIDR6Qh0Objrir4B4GykJM6v2COEQI6/cmbCOJhzMyPky2poqM
5vgzpRaa16fE5jKo2NtrfsZg/1zvnaikEF0rJknPOWCqmXbYzWzUaWYeEcgwgFqR
k/fdKbWYE50tLZHc2RRLQ4MUVoi/q4740r/VN5a5Ryk/3vF/hWCMr76PDwLJYeSD
lsV7W3xvk1KRgKuXTC6Pgrsw73PqxiLjSlDZ5RW0J72w4vQaWkpwb/K0L3nFXHem
8iXk7Z/L00WLi7bwVCDTj64UHFYmxTbh65Owewm0VjhKE8VVZ/RNmgrIxI5NV1dx
ltvF/UfWe53JmXQc1DfieeKsUen7rV3DM/IWR27T+g281f2x89ydU4nlZ6/vDIVy
MKOIGtj69Hln0Lo9z8yO7Vfrl3UScdhPmVcMtCObGHKXshuTzyZTgjc19Jk1B+Yx
uQ4fl+EybjS7iGkf15VwfQ6kI5avivwTUu7vba64kMJDygq2iUWheN91WSj9sAHa
Fofz/aggECZ3DIRw9fUj9IaH3vOhcXFWdR0v0JuvBNURNAbaU5ubnLJnUAQCNkcl
70ACba0J+bPT7ZCjvAUfacSo/FhIHzv2LkxjdaNj/ussSt7h+PC+IIZ3e+teji6T
Ha+CKoOy1vW9O6cq8UqAsi7CcIlJfIht+qgEjeV8Kx5MvEI1bh4o1/gq41Rp0CPi
ubq+35E+4kLUwqCJzHDjy+51dHH+W21OjqYO2/OpSbYA7ZbpdEj/+gF4uuQI5o0C
4/H2beuoSRYObTjlHiGNtZ2a8Pt4gB5R6PgV3SZOko4jNgC1N3uKgGXkaZPaTVAe
HUU+czV7eIN5FJNk6DR9DWg1suNIaztT5iA2jT/x1e/zWKc8dwrst3WMmPBkQPyT
mnHIgoniLMKeIzXSEaSkqqc0gvio/2rB2wPyDFGGaFsgMdUxpHkXUuGRdeayAa0s
qRKCHju2SbVVOLsaXdbgqqhGEA6C9yUQ4VRkP7PTa3oF3rYo/jtog/HfFSUtK+Mw
I6ADhpJ6gPPjyUcisBEewikwohw42BSbjX1Vctbtlhm0t2M8EBo2MLoh4xI6W2Wq
WaijrH5+OME2lLVi7JZvpNA9rXHkDL7iLDh+jZCdYnBzFYUbq48583zU3Z2GN88o
99Wieop1zo4NkM45BHv8AfmuQ08Up2LSY3Krtw7XqhG5azf3VGy+9zLBo+HFTdOy
2ezPFoG/wxmRJlbXlpgLZR+cwfzekBoAcXF1zi0LJNVMw/DAqyL9fpelvhUE/vSS
PV+EE+UBLxWBqxliLyUjnP86AYEKlOaA/N0ISUNnI9b8aU3gUI77TRxwX8c/TztV
ifv+DGPK15OhWZiX/iHpP0rjKrDQ4AnWXvxuN2YAtDgSIKj7Owj0hxhYZ98Kw46Z
D8Hpzm8udSLWjLF3hBNcW2c1RAhYdMBhkwOblqn9M5zG3N0ZJtdNgd/XqAcZjvsX
1hs/WjYUfLHxVdiZHYbjYMM/QrLWL047Pc8i2Tyk5V/VSdotT27GWGKbE6C4dWfB
ZEdir/uqQK+QhjLCBBRAPf+60dRhxwZY5LwEcM/uGoxcSZjbNQBIZIxg3Gv69p08
EuxXsVTBYbCrw2Wgk32rHIYLNOOm26N1LGJC5B5HA8s/oNGIj/xEo6tgwF2e1iUV
41uxtSGz0EQHje3fzPQvvu0jv/BdK4UV7COoH/OFHHGE7Xl3AN8GhzHK6gw7y3tC
UghqlsvMxCWHie64yRHUwfJp3OKSltQOw/9phWZLo3yi/w6HsCEryYjNxQLinOSL
SfTlA8/xzD/tnGlsQayNdNt3YYbMBwYM2xE8xEL4F0H/85CByunQy+TONsiLbsY+
JuvkG/eOF6Ybl2dmw/sMuFhLxxwmaWnSicvE5zKssNSPWbQPB0Zi1XUmgsgRmtzS
Fzi4/OWTvr/GYaCkJ0jiv2ymAgrV9xrAL9sno/bZf40TGwHK3Lsq9ma0Dmabt/dk
nw6sbosIRmx1xih7Cd4Chd37m7efw+DFEMzGR4C3CbgmXAdTMONIvu0/2Et2jEaK
9prwwk5UM20m55Lak9ObYiaBi58T/CB9nLHkM/YRcNBgKBigZ8MuMj57uMvpnx1N
TaijUZklF92aOrxenbNQbVaTB1NroeK3paQxVcrBxxsPF1PqtxIM7qpKjbKv/bmw
ezVQ2oKTc3cl2BEMWlIxgwewaN/E/ko+Tkqo/Qzn2qgW5KZMuQWITVefWoxpxfBh
wVQ5u51Fj32ro4C+6EnOGbA0vjBkncjsoijArVtxMunk+IOc1akLH92W6e+w/Pnx
UKK1GHRJpmMvpwRNEAltvvMFWNhr3TnnwW/yVx42cm9x2HVAgZaBInz2kJd7YOpI
ann4xCMkgjYxDw5c4eBUxXfFbBzRm1mNJaWa77HRpXKU9zBmYh9sJARGe0jEtUgY
yP2uCJBUQcOwbGh9GpIXFGbNor42MbrzCCyFvBCqVNjXBd52s76KWIou0L0u/vLy
m9QJO97zVci8yfeah034wZbvyciRacrITLhK6nyY5c0xFyw+uGdasU6gjsb+f2c0
QAmcOgCZK27JvggpIfFtKzt7TeMSiQO+lYF3NC/CSprQXvNAW0DXbBlqS30OSjZl
Ixs3vZrQ09zfZCbQx19X2t3OwS+cgjJMmXkLDjPs5Y/gJbbpoVnC5zEdZRxv1zJW
dAQVfYZXLz2of6si3yIfH1kCuK+nRgBefa8h8p6loGQkDNC+v3WRatrYtVQFVrZO
zayQ3enjPfoOtuFySvB7PAk7PfjB9/iiTkU/H+xZsK4UOinSj5fmWNY+V03XkROY
jhUIS16cOq8up3qi0H7DYahHZqUmstY0r1lE7KR7t9yJeg/Z9xQY1NqAE2y5S4j8
q9qMa0GTYp826sLmVpGq5h/AHSEXIhivveoHfQGsoS2lNJT3n3ComXkfc5C9hJ6o
tGs1EHNbMfWW7yLCfL3wpGj9egpmg2Mjd72gjv1E0qqlWe4LfiCd63nrrLota8AE
10XtIhia5wiQ8E8MsIfen+HHMc+B70pVddc/Zy/Q0wQ+hPdhhBIETUaX3pOAQr1c
eu26V/iJjPWzptJyULC8bdgLAu1MyVeocIrJuJNKAOGKzlE8B/4xRrnAheVj/VK+
hf4rJILbyvGpUVvW40QvGHPiki/ZFxRaR5Ser7vcEud9KZS1EIhTlFIyG6cOKajt
orA8vMezX/u9l2bok2Dq4dlxRsKaLUq33I0houWR3rXE5xeTh/ZL3ifdonAQsIiL
bQ7e57A8RV4tGCjD+dnYi1ZK02biLCuzlSMwmUyo+/cGvVkAr6vJwW0E+nJBeYCz
4oX3mOj3O3gNEV8ZH6zRj0oYSwMg79szFjwTjcFwi0zCw/ikYJabyw1YZKiR5ZGx
xP755wa2+nYWWPXEwx9O5IaygSy0kaHnUOD7ZzaDQF2canUWepP+O8D0Sod1zSL8
YhlTGxBdvug7/Hnd02MDacRotjzhPoetZzRmgZ1+iE32TzQXrU5CEGBhrT4UrmKj
CvHpAI7dR9RKvA56+AxbTmyIzq+8q4HHuO00NcE0wpt0Q/K4QVhGaTsgFqGErVNe
pc186gFiUTYA64mlkJOdI30BFH4qhK+0n14v6X1SfvBrhw9x40qChCGOMW8lARQ9
ZqFbVoZFwXUOK7EP7rQtJ9o8QCgWxy3G3UV96wjybt9ypJ44XNmiEZTcvVCwCC8Z
iCAdOTmI0MqhyOhrahnJNeipB8LWO5XB4f6ktiYfHLGhdpTNlS7P8pxIrPUgGJ8k
sI6dXxM9wbhY5VyoVpoMpI5i0A0qIHUHr7nVYSJH3TONXAntm9rxPT7gnxTQsO7+
ZZq5ou1LRa1cPQOr4HKaa335MqDqkFsx4ZgbYQLXqM+S+sAjwuYSXW/TnxvSC555
s5kwLH74Iqf6RvxLwHExDOdalExeioXPZgbc6ZjrXhtOOQxZUfS0DrPBeIqHPWMx
n0k1mtJQN8XDGRAFO6mP3EJazptTpknATWe4qwrTLr0MHetBeP2Vj/tN8PsnvoRH
w0dLZlGXRz9G2lLaRLy0TrzciScWNFm0lKHWQ9bicKu03EB4PAU1BGs4eXtAHEVm
CimxiarNunnOo2ASnIMKZVBM5ywL/I1fjXlBnKLcl8PVLh5P6feTvsfEQv65nt0H
xekBP3yzdex9Svms6/f8a2WdilmCGibz/F1kPsluH1WjKjr+LXuR5uvxKnF58044
kHuYhVXNz3YqavAvXWM3ov903YLcZ4CD4rSNJruZwWwn+qlWjrfs67WLSB3+uI/Y
Gu9ByMOZSL+cqWM13qTwGzBbR4Pk8eLC+Cekj5ro90YvHZQEnzSFCduPvxHCTj8a
751Ag7ZX6q66uO/1kSDA8GV1QjAUcOCcrSmvGASIiknfyMf0GOnpwTMe7UdwDx+D
bza+dc0kX9mRtCFtIwldGe6jmW5SM043bakyB3WwNz7oU/3h6vjZZ5fWNVMLCXjT
nPEMsjztv3JQowoJnoJV03D37MbTbaDoHjFv/p4zTsH2Mp0eWdrdHU5bp05OdZqg
FOm4fb2OLlqcaQ/Os09uh55Gk0OscE3uRpX2Layv4p5Tokg78WF7ENe3f1LwSdpn
yMFf33JNAy12rTrJKG+HFIzC3mx+7wPl1udPozSWhx7C3K8C+QqBxLJJ5v2iLdIA
JQzIlnl1k+45q2rQbsA6nhAsCbD2i+3W6rC/4YLdvSTAqJl5q4CearcUP2OYNf7g
MV3kgZJb1cIgCMD03ua78WNS/1j3MKFistv5tKaMoX1XEyJ0Df0DjkvHNn9HGCen
dUaW8OiuxI8Do+Sz52NqU9ccs7Bz2YI8Bak9m8bqQo7BXNRyRws0e1t3wK6nfjrA
db7XVj4wC7fgk2shuJ/Ak0H4r2kd22LhPS5gFoL6pEjKddjtmKlc91aido0be293
T8ejXWRsDXMUV+MPkMtreYTQmi/7ZdCzrlU2Ils0wFXHHqoXiWV++m3EKHR52BYW
vw94mZ72ZXx89Tqtxvjj0Ffk8aLIYW8ssJQnZJNQP8FIlb7VWxtNvAlytSxKg+CH
Qb6LEHRdZiOySBTkYLKOMheJFaA+gzrAFjkYxMc/e8aJVYkEkzt7vLjpk5/Djg2A
v8ahJ3aROM+y3iO+DoniCHX39kWfnfZP1BgtEGcxAiARWxl2oHYEE2WXk6gy0Nmy
d/dOlgs7l1e363IFZX/GlIVd61LsXw3p5t/iPROg7tgRVq45Z5y01RUYKLgRW5aK
QR+qPu/EQ+JirALfcPsuLZ9lTGuuoX6JVYmJD6nnbR2XjoM9ShtB8AoMnINk1fki
8X4Sqik0LcC60OzTQbSPjkEhJ6nGbsszNIDpckTCCHkE41x6v2kRW0WKTegB1i59
cq9p2mE+z3FgYHKrhxit8LL57r+f1iUu6G4R/yjP+1XwbKIbv8LUWzd0vZmANvyX
+yDzbuxVgR5z+XiM9xVpvnCZaYb+9o4N5lyP5Y/nSjuo8cPz1jqPB84Mb7WMSnbl
3iF4j5wQvuPOoFAB+QG66980f1n4Ys4/EFJZPmDVhgjlBqVU/zVLKSOCvrtmhEOl
PG0gTc9UusDkSWXXy3S1mFHVNQZ4dAPak7i8Gz/26gL4J2eEJFzPj70CTOtgtCz/
rSfFm5VWesyIOoAI1KB9cYgS/ihZZl0V4Ua9SB5jcqKuC5cxCOI0GIxmVAI0O9bJ
VFnYx87QOA7sS3mBsCktLBu3Yz+V1iz6y55M3rh2EwJjO8zeUHasKDg2syJzKe/X
tjDCe8wmPR24NrhOrK/VA0lDr+8tAXKUlGUhOgCEog4kQGoKxQNdiNVD+WeJ+i0w
9s3GDJPJVsMe0+J+u0kDn/LsiXo6f3r52CsIsmwDDYhl1vGIgu+dyH8qRNHw4qNw
ONcR1RLnlBxi9V91ETSZYoHCOfd+5EsCMfk8c0ADaO0hpt9wVNn3lk/JD/FMLNGQ
Ovgyf1YpHAfiujRN6r4O/x43h7lGq6zpMZ5qHXcrVF0qpfLIPVfTtzzj1i22RzyV
z0cTqgJAjGm3bLDlWosp+jkPDnHhpsbNOwZT6jB0GHFj2fLljv5Vyye4leTfcXDe
wN1xC6e6GpZcroUSRAowsY1UBV5HYaEHmWWegtyX/ejDVkCfp1whtY8xFRs7ar/v
SAYd3BBfRBugTkXRnd0ok84faGTgmAkK5cHwR43HNvjI3wlnfL5j6bYTpfN7VSTD
YEXigJr1X1YBWqQDIB/bmno4HHp8FWVZwB95bvzT0F4Tl3FrREUcZfM41A4W353Z
iN5a5ifAX2seh9Zvi6wyQD5Ut+y55KKwAW7cwqInep6d6skSalTkqoclws/wPDwb
e9NKipZ0dc4rLBSKAj9RVYYAcBhZ9ptRdNO98QhLVUI9QimV3iEB7Fr+bdgBpDg7
kMGADHHvJx16BrRecnhXWvW3auWn444JoRYPLD1EkWTDudMPq2lO+tdl1uAV2pIP
/EaK07afd20xrXHdwyllN+R55tjftzE8T9Mk5mdSTHkMU3kxowMa/POgtD46FmcN
BAVdRrllXUUyqJDQmrjm8oVmGh+lvPgoHVhw2dgl9Gzmyi5/2j8sUMQHadjTuppD
6DRk6ysjTIOd4/4J9ijVMcRRJL3C5+saL71PBpIDT7o4KjVUvOB47okQ+hTulS0q
wjogl/mZBZD4g5zR2YDnWGL6Icil65XhDu0JWWDksyAzs+8Ydwk8I1OzzlxvftzC
RUiNx9XNYfQO8JGaqLf5OcUqfEUiImth1yufR+4HMZ3GGxm+xl/bBIYexhGJ2Rv0
mjhBofzWlVc19xWKQ83rMloYARsYzlhSCKWjkP8+kQSMB+eE22It8N6mwsqFKrAM
wUj/sdzfMYKFLMNx/thkdRvPyOfykxk/LTQcrpYiO2LURVfV/W23NSqcsWAWawzs
yhRho/PZdJDss8CYhemT2t1Q2bHcIV4Ur3rAiWByNIVZZ1XNkrsvdfLFXm+WN4Em
0iofE9tkXBjRM4Cx24vKBZO5Z1cpnn2xIIcKLW9El+va/SZ12WOBrU1D3GF6ziyR
H6w+PYUkrggRBrT2/RcRdPS9NzevwCdB0ROq5GNU9RD4bmF6nGLc8WynHIFzyiqz
/M1B77ggqACF08YTKnrDSSR6jp67rmLO0QIjMrUm+cAHxkp6mh+y4FBAiwRxfFwY
aokymiWJUHLQ2TowAwPmi1RbVv80QLej/CO6WvDS6BvvOaBwa+I6eoOuixAT0yOg
2AgIXlzXYWakvQKN/50+s8faBGNvrRhDR+0Ec7sYQ1zxf3CprXCd0XddF5RfcbBt
+aABDD0qGU1WomqmvJHifGuGphOU+eXnCyEojSgcjq3Vpxqu27xTogwgzEsOLa6Z
6VZAFIIP3DbXqDqDCfn22Ed5f2Tnw98+N9t9n1syQMGz2acmiz7yfwbdY0suAdmx
Fz07uB7vmh6dQF32iMp2BAyvj/lgT80nikUyjiHZQAphQsQrD9qrrFjXD/+OzuJL
m0E8Wch04Atqz8HozLY2RAGbR3/rw5FjEekFpDX02dti7ibqnP6xcxiMcqSRcJGn
stt/5yveENOXEIxxlxKZaS2vDHbonvinzX/X4R27asNxtba1ZzziVfyjNWciKE5Q
3XL1QEF8aoG4UafjVCryKwyohgtKOGV4+aNaCxgYFnVAGv71OZDd5CYVt1IH8d/S
fGSKP8O7dj5hz0LTHX+/20Ti1cLDW4Ga8oQ+rnCUK7BenlmaygMxhXQAKf+l8U+U
A7ItnIxwkVE2Nsc5e7HCol0Ghxkr+TpqABJ6a6dEsuaCeHfGgDsZdXwlMtiXr6oO
yWoN4I3EpAe7VqUtaeQCM1E8qYKDiDqhVJKN7QPlNDpEpsELYRIMDlXyuB3AlPr2
8qESYmZyFTjTpOf9dRiqVB8oSoT6SuRCbd4qsYwMUnk8zQaQnNPqbgbdKnN2Dcd/
quy+xKICbFetE/wvwl+7tU7KEHQFkAEyEOV1QNdb7zTMkG129XKQDZLoR6vwSRTM
TSDWRNkkzRN0XkD8EsDqA/jY3mA4xCh//6L23y40kKMccP3dwsTv5Xwfn++lSCKe
wrvhShjqXOpcu8eeSHaJLBdo+tg4L5PWsCIZtB5PDXqA8ZhQU9hbNl4bb1sh33WP
fPl02Cc3KoWxP/NwiXB3vFwd9D/b4k7FlM89jF0moFgLP1H155P23rHCJZrMhR/R
fn2o0WcSNAFd7tmcsS/TgBStwztWIKGsSN/X5Js/62nQoa+qrZtrWCp4h3ubCZF9
9q407IkKsarvG/WZWf8n/cHE4Hnq9bnhKKpnyn1++9w3Ix2cHD3wtjgZ7d6Q7wvN
NmYkPna6BibQA8fwBOhPKR9QgGWii8iWnNcLQtO65aPxAOOYi+icyVo2kFtTNUfD
hwmtZd8zZ36SVBQlU2BY4BuYyappgoDIXk7fO/YIopUC+M+XUOLYEAVW6Gqu8C9u
vBXB7zQZ64/x9wJHaPb2+v6AcyPFr3+saEnsjohs0mRLNsu6Or3FWy20prDtIvkE
oSluJKLI/x128Duuw1KFaVP4IifMxdFKVJroXafUTpvuqVpytXRIYL2Kao9s3UYo
IKSCYK0M2axZ6g9Z/L+PzvqcBX1vA2dSdWhKUp2p2hJ57NpxqMjBQe73CyM+ibM/
Xr67Ku/IBYKzUtW04YW0OHLKCFIHazlhkMerjlox/7KHekWQQIUV99SYLl7lXU16
CwPc7BKqIZkGeR7+mHejxeqYbTUqOXaENl15O799Jy9JK45QJ3vaSUHpjXLwq98+
wKS0bX359qgiCwSOxGhjKJnJpXlTFc/0ys6T/DFDWy0+FtIiHc0kwxccR0abn0rO
H4njGUPk2fP/gBFp3lBxnEKdRmV/1aPXYOcbAVhIkEfpf8kboQGvxgIiiAB5Sdb4
0dsAwy3XM/0b2Q3aZ20l2GuFzMeevxcX/D7yjgOeYcXDZ8SjQYdBSFT7XqdDzFNZ
5cJTie5xuCdJcPe2c1Y9hu3BmkisZ/uxwove0iHj9ZpRQsEakhPUtrnHcT0vmzjd
Zzbjka6ip0HvodilfyQ5fHmphIHRpfpT4A0TW+xlXNAxbGZpGQ9Jp6MYw2zxCZoA
MlZpsMqttDlANbCEbUw1muuoL8xMtoTXiMg9fhLo24nR16E2wF4bJ8RMEUGNZLIa
79hNQ9wNJSt/l6w1YkkkeCVu/G+rPfYCo57tkIOpzJtUMYJTYbWoYbG1rP7rWkSg
2iWUvmrfM3TfPQiQtj4EvuER2yo1ktfxXJPQBpVBJAkXAeCo0JuiQJJHxqoUyWes
uf7tY7UnkRWoTuEqvU5Lj6vmmi2gavRcbE6iWP8wmpk3O/cxPzzsau4N2TlOAJnx
7Cgyxy3YteGszHY96pFDsxZV5MznSeTXMGdkQOzKpMW/lZ1aIfaE44b7o+aj9RIg
dmRBeUL1zdWOmWFLipL3BlPvQmrFvTYqNg+6hmc0dtqqiR+7IJY8foiupJJ/nLXk
o6QIzXmKoFvTVBg8usN+ix/hBDtqVby1SSMrH+sDnD9Br9syaik/hwR1Iv/aKqbc
5K+eiZnJnpWcPlwdBXVshK1YfJhF/AH73wmdyyW6ESBGai6zMmaumddF5ENF1ZO0
xbkdymfB6Hl3ZDnZqyZVnvjyf4Eb5jKPYXmT7WvGynqM0MN9Ba/0PxXh3j+1fFpK
fw9heSY0MzmJcTjGOvq6BhrEecWL2YSde93sE2P1ExtPseq/Pblk7hd7K9WmEw1l
Wyzt3adYvjBlAe7CO1mQUyskBwzS8VYSeoHAkO/uPpNQLw7nohGy3iXdQoCKJwxL
wNfucYNYib1IjY2OFO1bsYHjgwiWcsRx8qZgJnVPpNI7Sxq7iFeMXHnQbPNV+vIM
o3PA7nbi2jGUkgIHs729ox6bE+p+4yjIwitFNfuJ/XfcUibfw9ytCRvwSg67G/2C
tdaVpUYPHXFv5ahS6gFb7sH8nvp30iqjJdBdyrdYjfWoEF/PTSWxOBYSPwpq7pS+
s7fq6/P40pOuGiwMTBXMEGJ0OOX0wwoDtfzhNAOJNOgGzAntk055cUoizhCL8rMU
wf6OewgWVVtmWY1Om9GP1t2I+YVFlsLcCZfQzoSmaH4lhaVkuO3LM8HNphb3+0wd
C0sUTEKeKRH2TF3X2mdvdiX2bnOGdc6ZKAWSkhECE2Fv+BuOFrlMC+OzYmQ+37rr
SYDmZ9JpPaB+MFE3wJQjt593KrVx0dNpoGSMn4wunsbivBSA3uoCCcDnwplQr5bQ
R9AAA7uR6BdUtxfZZTLac+z/eKB029Eg6DIl9/Tx8yclGGEOoHye75kyWW+0Z44x
PpR6xyV+iqJP/JHLwEsS0/EwxFC0jOWPLXEfmXmHN3Rr7SN3HlaO3vL7iLjnW2IB
bBQuqi/6aXuEIKleWgptcWE/9osE0tiEwKLl3mbJoa7yNGFIPAGA5h/kpJcYfsFO
4rMKDO+5xmYVNqFdikuTtzE0NdFbxkXvfrcoQqNacjQh6EfMi6ajqFbxM+3a/J4j
BNZny1QRTIwAFJfzd7jnusHBuD0+FZczXu2n5U7gFIysFdRIMu4KR0XU5I+ksloh
LKNcW1kmBc2hDt2Dvi0M7+bj4K/v9ZIQyzaB5CrggHoQtvfEdM4hWCdc7dYJdkD1
tQkOBTHCvt5QeR5cL6azkrLbXRvMkunma/EIB6ztER/o6FHrkkPt6Mc/PjiqAy4d
BTL7rBS+N65kzxrtrUG18CO/h6Csx/qx13X0Rrdp1c/5yI17mIC6JiuP5ZaSuOKL
vyjIEyjrFmimIwm8DvH4Gt5gaQ8Fu7MSPD4f0HfyprTeSV+VHIUblbUAxjH1eLqM
2wbfz1HHerelFnNDMf1xdYxhk713fW9FzZBNAFamsND8vaUHjrmvwJlFQGP19Oz5
wMdVehAUaKw0zFkqftzgleRuYCQT3h6g1ubj9g3HoBQQVg3wmDTzOYwQUaxyH+ky
z3vx7oYEWt2/x96ZAReEVM8q3SVa2y6K9LL849VkOITXhBHxjjodbaWszMaJ7zXf
l80XblASMIw5esM94OREOttnGJ8fYnPz6J/xVXbyEzEQLjqk0PKZyycLyb3Orozt
LWXO3DEsjUb37b6ug4A/7cOAKfzGQIRJ6bAiBRj0Q1ubvOE9LoX451N/v2Kd798w
p0tkLonDpF9KpYhY08E0kPxYmCaPPE5lkFHcef31OClAnLQUTTqssfGMya3HpWIc
7rtmusEIPWdZiFEUo8ZfAtb9h3I5f03VBiHrLOy/TvyqchGc/hB6eJOmecRlYVlX
/F4z3ps9DX8U7pAc6beRyhJPYVFxT3obHuz0oi/yNxAcUo33o9ShY7nraQlDMwFM
j1d/QrTnO0+dunIHDtTlf6C1maMgPqoFxkoVp9p1ExfpT0wMUisEYFLhX8ejqns8
Q+ySI1DQqR8dVHYOVKgyXAMbNGdb/0DDq0FL6RElhAmx4ugOQSoVcN/xnDG+yvyl
xfR0ZIsqEGDGteprTzMeWZC7XjTY3OtmNG5ml8fehNSI5rHHhywdW5y3XJYkQ7Pf
9szIKpdmZN3XVHs6xEwLMbV8CtJsD14XbZxiEVbTuMO60GNPcGnztBgWOR5Aicgg
TeUkNHJv8gtYdH75O7DSgyWJz6SwRSPiQhcXd/nW1dqtaib4pe4dYjjBMziQrSQK
qVPqTu3I57FQGvJ2ggIczHynVlzgbFcNkcy9Z8mhyblyLJvXPx4fmGNvQvwdZP1p
XjOS/Y7s/Ujvoii97sfZJiZIew6118BRKRYu9xaySWXucHk41pdIgn7l0Yj5vEPJ
JnuDoNsed+rRtg9VGkwAj8iLNoInIWN+CD/bsATSgVO22IsYC60kWZYqp0W3Jdfg
GRhWNhJTZG/0IjeJxsA9+mhbBj+69HFC5M9eqrm7W1H93QuoWDgx+pT/9hENWQ79
EmAahlgP4cpyc4fqzBOX4ZBv4hUCNX/di4TUIvFXbbp4nKs32zXugpcFBeLnEqy6
ttBJ6UufWLAfoRRKvkwUglbnhXkEXyLP4Jg+BtW8Rw1CghMeA+dVImv8Z8BMgZ6a
TYGlnJpvZoRcjc49nlmNQRdVkEu8EFSQTpxbX8esT0Vpp28U47I9mMxUbRNQrlxo
OkzLw/U6+QL3bVEXP+sEntBmYZbYX6L7zdC9TOA4wSpaaYjk6Mjz2aXHLSv88occ
4Cx8SplNSm6RFajf4wNVmw/NJplDmSEV/dJEGY7Dgb+dCc7T2nhelf90RyGsR+F8
Vwo3+8PYN11RpGLK5nNI/LIgLV7Pw3qY/Ha070aGBlzLuBGdhPBDlGtNHQVIBatR
MZuLWX4fR2v7DsqwAW/1hbOphiyrhcjrO4gjp34Az7Pa5jK2qGMe41ErTkc70gB7
f4o7yh4dwpUb5zgwGkCU6ggxVoo/J8wLTpkPm+S6Lwg4AeFiSdY8nUAaKNtCVWp3
H4Z4Ca9tODfYNCOHA07s2obbMcvOJMggyjrRFzn3dGobG4VaoB0g/tLXvEJUJ8YI
fpqDcj1PD1hz3Bx8rz6v+Yy1IsZrWg9MhGnHJbvnmNjTyKmI3ojQpOBNq7o7KQSZ
Gkejnh/NmFDIdUh0Mv1nogpynvGQ4cuV7JpaxhqDTQLjdTNVlGJ7E2jZaJe/8QfR
FkSKxMNrHvm25V6LfnrGZwRuKKE7SrHcN87UHd1hUtwTyAwhjInwLnsBW0OI7YGW
foAqaTQNXQ8oyq/Y7vPG4BkKIzXXvamadsVCij1kqh6jA5qZ/E+xk9IPw3ttZBOj
yvq2ugiCYIJD/+l9eBz3ZZ39HC5ebBOW/VYlQsxJxp42F1RCbb3UDfcEiZKBqW/4
wYrjphtf7b40ow6jqe0Jqp15z2YWCaPv9ctYclM20vaYGnyt6/k66QMHwRLSruEI
5f7GC3Oh7bExeaIC23tzEkh98vhuBzrghB/d1OlzR5fWdogDO15MIWzur8c/u0Xv
If3Jl5RY6P3MvFaWKjCjs4MFL1d/V64KvqrBxUHc37S2aSj46g1FheN2jo1MRxdw
VpnxI8HJjI8YOp8c9hr2zEq09Q8n+NbMXeGtPq+WODRwBs8Q2pVijS9hZ4BeiWnY
WjGTMOzgzEm8omUqbKLZ55UnmoKDidM1eLySA+jyAbknH5CBgN9BNWGU6EqRhauD
Bl/yJ8l5OInP8jO14XcqvwYx1o8u04NvcaIiydSmw4oneWOWbeHgliGowpKcvtkY
osm/06z0c38s+v4XTr0lF/gh9/hLLvaKzvP5PxjMYSYUhdv5jaawwDIVLEFZKdC7
ADmSAyQi2m5lBV8kg3BP8UMGvpiuPl2HN/669oZbyAA0xqVYk3qibPLDtdwh3QsW
xxokZFFHgSCVD0RA5sYiuLgkjgB4WcvQcua5u023xOCr4TkT1BjoqU0lwsWMuvnq
ej+TBGT3sYvwz5kJO+PrAnn7v9LUGBdiuC8v7TwMj4f0FZtVOG9kcuR75Vc5qiRu
kxg1zBUiPX4ae0LgMu5iqGb7f+e7np1L1294NB1jQJ7ZC35k8C9FcGF4gLCSiS+S
iy7w9w2g4Yx+AkgcDfA1fFIm2TFo5nhtbVtD3YlMu5hzEh6vlLWnfvoU7/DoVO0t
IG604h5pvgiu30oDXVK0mnh6w/IEsGPmgYDh9qDtyPl+NHWlTD7wVVMDXMt8rRIz
Gpaxgqz9hSOVnEQspKVyGVGDcUxPWq1v2xmUBi9fkRJLM7opjanayR7u7htP4VOf
A8E2vRhZ+yu3r+hYb57M/fq84qRcJqDpOPyvyM7WAA95Nt2wBzeQ29hVH9ZhIhcB
p1JetioQu/azvLe8JvjG4+8zBFP9stdjKRtWvXWPxlqHklJ1TK9B7UWkRrkDoZyI
BkiiOGPTQA4QJRBI9wjY1+BM6mY14CiATVOOjK1ceXlCsbHhOOQR3oMXyV6dkTiK
l3vcH8mSRusdFWAXq8syxntGJ/lZkmVGGzVDGewtR9VLJiwg++cbuqILz7FOBqNt
stHLkbvfzXi9E7dZ1kpnl5UWyHtPPjtopqg22QRi/e5d/kOZJf/MkT/W7Cb4TEIm
KZ0/rIEtYpcBsbsa164RN+LXQ9VOM9YCHdRsNOMrAumUZvnVB1S3pRnvUvhlOp/e
bYC+PFSaagO+h6ENOb5SH1euA4ay7wdASVP/hrkVCu2guAyxMdYRAuLA+40A/G0j
vsjJavqEAYo8Ru8ozoWzXUpTqPxSlyM1HOKKlZS7HktOlMoIpLUX5dusuggMsgJK
yp3mmdtmgLdqWuVxEP+siCpvYTkbHrR38/RiErOEnVIo1EViYIQmIS/Ee6YhLQ+L
Wm/aizBkfmgppPJxdlfFdVkbalCwJaYYXTjQsw8u8Ex09KVnXMeoJaB9iH7kymFf
NJlq/EGoEswnHgnS2c+rwfwezTkDo478mWFvvuylGsZa6vXmwIU2ynwkstSMCJsi
mfkXyoC7PX3dWGMbBRwviV7a8K2igHjCNx9INpg0OqBOM5Hvq6DIhiNq5OKRjys6
/+CjnbCy09mEHxCNUiClVAVuVMnNc4qZ5yfgD1ja4hoqgy+OCOMrvpMRqq+UnNzp
QZ6EkBW/b/UsKTB8WcYk/xwmj1xoGstloNpw769dLJQiX5CAgYvaRKHtyDYi77+h
V+kMtHRJf+5ahlQSoknF12vtNApDIMbYjpjmOaFSEZX/GKUFHpwqqcXq7bQZ0jGE
KlwwsLr0Y/yQhv3knCrQ7SrNKlQ+KhEQmfEVo36SOJL6vDLATz273vIr9A0DrCgc
T4w0xxt1Ek+hV77dxZgP1xa2yQfXlY53a9hCBV3CGAPJd/YxiP9/0qCA69/ddw8a
0ucoDfWOl4KWZQi32kAlzl+5E9LpOlI3cq5v6PYlKl7cqufERVFHXfNytDZjN++P
zi7fWwDTdl3Ar9bgc2m59dYNXBsjLfRNUb5QoQXO9sMHPK/Ee3PN8OYmj4BKTY18
hG9hA+6xtc2DjVxwMOkWNccfvgjRyvSWJWGxaEfHJJZjI9whJ9Ni7iiK2n/DIc5f
F5zRef6BZzVRwCAWFAAcG/Vk60HJdSLAbfOzeY1S1uur7TkidlH1dpMQh+SZGWH2
YQJ0ctYz3OkQrXPaRy3eqD3c7NT9xcY8PympvspMCWsE+eAjJyfmKFgPF2hS8IS2
8gS++TkIMw1kco7oLaQLVS66whKWcIO5GLpwN/Fygd5sklZAGer1ggmhEmErIo82
BNfESMNqZ/dGditchePC1taVLiL5Wl5QMFtAcj4QT/74GYZfXFxb6TSyx/WG7URG
qlu+EQcSglig7PP3GUrR1UOi85u2s/Q5+ca53ColQU1SsYnm7rrjfYKaJER4E0jQ
BQw9jchU97jXgKGa5Dz4j6lmTIOtt67nky7986pxlMjXzP2PSz8pSTsa52HD5Rqo
s0aZ1lRCxv1pDn4q/HVVAOVsXFFa+/1MkGidJ4yc+fU8XukphJ6Rd8DFsONnBbvO
eLkDa2UlUDrtrzHytkmwPvNvuPfkWDX/IF/B35lq2oG3Yv3G1+A/we8tFMzg+SFS
1zZRxwA8doy86RFQzPJZqlbe8BIJosexSPhfSsZ1m7b7Zwwu6xJ4beRrxCt7W3zd
Si3nCyZYPBlEdGqGhrW9fsChvkU14q4xSQr98JIz8Yx3fc9XX2CsrZTnIp4I5HXV
MGU9o7akTmELpcV2WKsT4CzHHHqeyuAWz3je9a2HHCYwuqrRACdihbSGMrIBWZEu
CMyngw46ceH+4AzQ93hz2kF2CL2YLMtJB7+TYpKZrA8+HWTEBt70SJFVVuP5MDFd
jbNW/1+8ewwh8Bmlaqv3RN5NSqmIVgLSTisWVFmhwBTObpsQGoU4jU6kfW1wFOPD
NKQq2jbfvSAUWv/dFCGHzHvHxWcWrKjJ7VihrIzQPEMQrsZO5R4da9WVktq96vp6
oeiaatDF0FVqOnaLz+8MU+xhZID2FHNidI3aVe33Pk6V9jK07iO+NrWMmriDCT0o
avvfT8cG8+RXD3Ef1H901aWcHW05tqe4oVVGN9jZy9/Lc8Nd5eRIzr+l7b1cwDKG
e09YBiR0CYfW4TMTEtlPSF5upOVj/yVINnepNuGgy+c1gOv19YrHUhDtAZ/Gh5HH
SaOpYmZ9D8KRg0GiVsOtxAooswRzkPPHqoR2qvj6Dr0/G6oTLEXrB1DCKEPDgey9
8R0rF3UZX+ml7j5yvQ1glNiO8SNSyBStri0cmJa8Hl2bj1S5t0EgeNiOtxTwr73F
xrLJ1ol+Q2ntmts+8PlurcBi11vEzWmECcykGOECHzWwZQU2av3mom0gL10JBiaK
/lp26vsEWGb2xCjOm+uuyZ43zZmJmlivLqPMiaRWAH4DsB/MDlMB5LDInhKRMf22
9njrPyU8jvlw3iYQX1+QYR/r/aYpGsY+L7XKXent6reNhuPyxgNVorm8J4WauuJO
uORjUXGyfp+ihk9jjygtwuZKeg/ZKo5yvnw80SSdkefXIojTvxs7giGHZQZx7hp+
22TdGxpUE4xgClRaXbXehttCEckrGyXh6kzlvfs2RsCkdxRX3ow4+6/kiCik7bvh
hWfblSK5GuiUPt5yMREND5HWnxsZyg9SXKz0IOOMZIQ7z+KyT9TNBD/TFcRR7oWZ
ix8FVPq9ympXuq9ONcc5cz0x6iLnb1TFMGTi+/FV5F4O8J8xvko/8pHDRB8ySzbO
D4n/OGK1yNgNLxidU/Kfh+l4iFp/0nmq4dfJXN2AeffjAn/tK+oTHfzEGsPusogK
86f1QU/OVU9vKbFpy/srpWCeN3nJaCkLaD4D/gg0sYIKpz2y9veCbONDsWszts60
Ekonl75JJaDi1JUEmcRJMeM3aF8Or5D+dP1+PjJyW4Ka6MkU2rXNTFEYcvrPg3kk
6efVjcVSmrfzB5YJSVG53OuRIbV+M+OlCMTIxs8DGk2Jnxhw/ja7ihA5pdHgot9E
DXR2A3hnQBcZMBq8jlU4ayMst1UPMj/VJ6HnbFBmo7r9TifrM8yEYMv0lIaAQLSz
0rqIzvxE/wTTp6bwcBm6Nim2pso7Uua7oJCwaTeTJo79zTDYKCrzl+CK0qD5d1Rf
Ku1sCEHbd+4Ebv07CBqDRVN+9MwkilFfHHrZumwSu0M8a3NKK68Fg4c58FZOSEjC
ntiH0PXgcs+1q1nUCJHYpAoFzB9uxaY/Y6GHjN/YYK+ol4LSuzSyq3J1Sz7OlJWH
zqjPPXEr3ZGcqOkwfyl8hZGiFn2RojV2HwD6u5bSv5Vv5/WS1nYAC6yoeQDEqAcZ
mhhsjTOCP3M1htWBeV2EwnseLwOwNXqkadsLnyBjYIw8ydi6aw+3wf8wHlbu5Rbk
26sWCsc+HFeJrt6MA4621EOTIRyAlDWddWmcfcxNacPxhD9pdaG8sgNLH6PCO0z3
J8gtDKW7/n/QcRcMQ6i9hWsJf2w4r72yK+h9c+ex7+vXMycSpLBs8m9uekTeyvKU
C1fKfkskXO5gDL6zQAoFS7q69K0ru2C8JvKMkOryzun/VH0RV9bN5ypoDgRmGXis
mjExB3KfTOwpdakgthT2hST8lhciWSDF4kMpR7RB1cBXytuoYgT6CgruV+7Z/czb
XfpN8id9mEklS3z54dBRIxOAjhD4RKxaCspTf/RAiRAmSay2ThAlJNtWLsOAx57K
lCa4C2YdHI8DP+rZK8MDy9DjM5VSxbWeEx0yA5CcinwcksqWGbrUrap3P53V4k9S
Zhcr6+scfpWh/+AG9wCc7iqjIOqi/OsH/20oTzM9lWLESzTI/Xs/wpUajLYMI8Ur
SUT28quMP+bdjTyk0p+8XZjxLfUtVnuk031WdVW1CrYlrDic8hFgyjO1IOOwTSgD
EQmvrNqUH13mc/wNU/I6C2sywaGwGgoDTtQwwizyws1xLhqsVvrmbCucfuGDHeG6
OG5ISbFd1/Dl2sDA0WYY/bCrRKmrlrY9Ui6CrmcpNcCyTZbUBmecmiV9EK7Xsq/e
h8TCOMp/H3NN+MvreI2HVMavPi7qUahmPKjcIejZ0wa6Ku3ZG2G2wXcje+vN4RTn
RmFnWVCECfsu1IkoWYWHTeLdbb9rQL26qh+SAI1lTaYEtgArkPl80SSmbaw4lqai
HMXeIBADhjyMpf/zsH0UIC/Zoly1jDmoVR8aHnJI9/vlxbSbXYqYMB3nKNcNoBCx
oFhJOaYhH0mneG1agVRttALDysV965utA+OG+8Gp7VCGV9JaSy4JFHz+eXiq2YV9
wyAx4PypWF3tzBkxb8p00BaB9MT/iKoDYX0jEGauS8isBQhn01fqTKcn9lf9ALBW
MvfSXQdHC7mcdQQg44tJWjOcR0Y/+A+OsiAMJJ6WumosJ0WfA0QgEULkT82SJwud
dwmkX0z/V2wDxJppK0qGrcXW8F0O6xEHLMcS6ZdW/U/kCaJdl7L/n2/yuP8uaSnj
x6tPazDpA70R27Qb6Y+v3jtLaKpIjOAxpwH+0e8CXbGniSWKbFWi5DEefgpY7pQF
gg+pzce62J8IdtpkugdTgKtfi/6MITt1v/FbZG/UK4eBtjiBhCcNI8/Jy8VHfAmE
SYcYCNEQ3w5s6nt16VSmNYX3BIz2leZq/uJm+6AqhqXJD14taGKLhPrkrlCUMk/E
pOvwrwz0jV2mA+e4aWdePj8jmAoV2u0mwMJ9Axgnnd+s29pWJzy7sphXI8wQuAPk
H91JgTgB8ou0IXPVbXcbQOWBgiyApHzlJsR2DFPUKwa7cmB1aXu1zNYbDEnJFUEd
i5WUulpmcW1GB/GpcFWoTgQV9oUQ2kPdCaWE8yjUyd7m8DITRS0OzAX1sYkykeNI
X1ROQH5D3MkxZFYRBELWDHtH1Q3SBj5jg5umJoUy0y1K8G45k0DjjlkMANbDcI18
orjIIL2L7Eiil8F6+S7ZL1YTMyLMH0zbbNR+7MPp/ROjDeBqrM5uv9+n/ook+HZC
VNnMJNgifkICv+zUhjRUxIALCX092y7/wBA+RfstK6zUXPlc2fc8jK165jXGnshJ
99cBmuD1W0Pcz7SeHqJaPgMpPQ1LOBA6TF6+OvibPqlp4crIeLWFaKcR0wGdTgFZ
s4LqSuFlZmHyQCceFGudamr2fPkO2vCpTJXtfmz8zLcdUopXfCXgoUcEt+j+rM2y
jz9tg9QtYW4GyNHDelW7c9dDBMD+P/sfmh9vvvAFy7pqoGY6XW1SZ5rYPblmQiyh
lCU83lApsMj9ci3i4Je76pUNFNYJQ+2KF6VQAObcuk215wcnyCEIBX/UeQ6gVy6c
DpabDMqs8dNk6uLBCBq1x9/dqUB8f9CUzzlanUYTXAp2y0r4WulF3fEJPdHVhwGW
jtXpOt5/QvhPpKXk2Kq2qZRfk9Zj1a4Z4SEHuHi8g7aBb0X33XT9YYS6hPHEIsVU
PD6Cnqb8smhgCvA9J6JXPAwENje0TN//1eA0Sgi6dN46n/B8ppc2szbWIJJZhGUE
hyfR46a203y7za6Fa6lLcAnFNjst3pWFwwGfQ+BdsloXQ+b2bm4BxxC6XSrgDRXp
dAbLjXzEcXSwp28r3NS9dmV/0d5PmbkybeN/cVZgjepqV6mqAPMDq8ohsN9Y1CMq
xkCR198pNsC8gXPMKEgFme2qmOUqlZ+GbTuPPcAGtdK8kKUa6xV6JeStncEqDVpB
fN9ZGasHjiTngrhJ1gRTwSDxLx2YBuhqyRDnYXp8aBXRN/9mx7sr4MgBA57uFCf2
4tnl6sNuC0YniTD6PjAaobykOT9RG+iriWdMOtJN4YpcDMRVi1kvFQRUbe1/zvQz
EYhKVKev5QSKe+e1wLLDTjQGNboBSUGDRed3Pt+4NkpxUMaZrhs/zUHsWd8VXNG4
WW0pPYg+3JQQVcO7mkvaQqoMMGxd56XUEPKOwFur3ezy+XeAlZBiGWOdyZEb5EPy
ktzc7508TqTSysa4bhsB9DyfaMllXiSLKh1urAUflReT0MmBFHC+WGH2vEEwCdCw
CxV2E8wgmQN/G8qRPiWRxpwr0jDcU9WVNP0NftAt/bPY+tgy6Ci3rG+/o8g3bUvR
dc7vd3d7Fk4yjBW8151dN6OQxPVcdCUBwGIHqA7d6widws2vAqt7fp3P18aQOjqF
nwGHNKQC1DFb9xniulA3+DXhcnjE2pp+f2bvHvonIH6n2P4pEeFPrCPEUKv9xEoD
YjvCFMKVj74/hEngILNW/ANm3xqwXDZ/H+5EI1N7voqQ7tiAjHUSi+Db8WivXWrM
8hpc/fHBr56U6ibW09n5lXFl7gdvBdAjVlbe1/vIB2mba4QFDmbJe5idCjbuZpPn
3X3z1gxkXUiPZzCALS2HoJOCf8phPu05CH6Z4uO5tPszrVfUIshknRKfuDng1yRE
L2Ekl3/aVunCE4xc00tzuYxm3PWfUJsDLsS1twsdfimrj5FhXO+3RM56+jp5KrhN
8+Sy1a14KiVAfnAyeFuc51BKox18xiysksDH5kPtqTiWHc0pmOrayvs0YeLItzTt
PSf7GAybhSH3ka6VPigUVfdhjSW9TugYiJVWnDkC4ffNsjpLtqoG+++0qv1hPbr2
GhlfLnVl2Sw7Zyyh4MXFRFK1WQ8YMBMBzaYwOfLHtjkjjbMkM3Yk31AjHyo2r8V2
yWCvHs5EdDM+GB+yoW/h7VxCl0i5FRfqSvaJsRGC7JiepjMDn5Ssyh5YBejZlEkn
L/gKpjGiARcsk0CZNv0ctF9YUVFt+o6OF5grIRryQKDJnIWWTc9l0t4NNvz/rjlO
58RI06PciTYQ9DHfr1Ov4TFEEhVgNL7WHP4dSknt2nyNPiEpf/wo+vXxfm00sRvC
/XezEHf8QgAr2NdsBmRSCcIqabmVxVGYcSwjtmJBTr4H/uH0PRPA24UQeVKL9ufJ
iZxtTiAm8Tt1BFTTuIAxJ240CUJ24u2LuJilkefUTKyXVTTjbu/heemT3wdK+pIk
kGF1IOoqeYKCk1NOytmIED4jIK+Y7NOx16fWYDSMDPPQkYdJ9jWYslCBttVlz574
oPzDo21E5WmPTiGSiwFMnJRXxnRZESPKviNtQaUSEa2fMgz+wTGqXLsw3M2fz3tG
JFV940S9oDOd6KN4y0Ii2Z65QXqSA7CZqlDaqZ/nQ/ayNDc92Oo3/HKUMVlHIb5E
hCV25mKi8xIF4WnfvP1DWwhOjKmmNd6BFaYsoVgpAvWrFlP7P/Bp7wJJLJi0RMQ3
2f27jof7D620R/ECF3tSVRTRhQL9pWPpa+XhBzp7VWHr8XjGH9ii4h3t0fRqBRq1
7MtCQpyFKrY8OFaIUQgq3Krgysb8vfYNJJzeXJsNpisjW5rgQv6QqyM/jyETWIwU
mfb2WLxtMgfLUij4l2vOLcZudHDkCiNNf+vFfsLWEzCT+xxhOP0wlis2G3zneQji
hYu8kS+0OiwjcITm1ukb/M4hn6lsbgVnciDGfMHcoOuruYS0wo5oCkeOTIOvkcRr
X3imKZdUuoAMAq4g7y2+d+ZJPE9SNVBZAxNhnt7qK3ujfUgzsRhSyIUsiBaVJs97
Sk3O/ZCRA7g+qZokLHWc7tYYvI6VDC9K0F7a+qZbu/PSgrxDDtrKe/9itYur+gk3
+aPGGJ7IG329dgR6J3sR5TSi7TNC7/GWAna0HAont0XEagIV2itqb+yCQFXwtMal
9ZPGN7pV6fXUYfDo6jEu/i9aImAEn8DHNWm+4LUxVDr6L91maGcdN7EfzJq3ESCw
yux62Nn2mMf8/z0tCLgc3n5M/bx52wRzdtvv3u50GVgAD9HD9hFGY0392XaauN+V
mLaYnPbDSj6mhERCecSk/R7sptx3xKve64SOkWLEvzNeZKAMQZdoki8nFVh4LzuV
SSt3lW2XmJaMoNN/ePcfnTm6Tij3RVUbZ1tMU7Bw7FhHxvvfVVfAW26RK/Qaj8wb
j9plkKZIqFLZkcl76n6IyvE/3Vh4zVsmqXixCQDYNarebW3irQJUouW+mdq37/Ds
sgQccPOdPc5lgFLgpNav94BIjgtt/6bEfQ7AUAxZokYJhCXtNakz9Yse7pf7n4PX
yJE/1q6Mnq9nDsiVnnfwDDn622JO7i2pbz2GUHc6wlffFl2OZ68Uj2hPY6wka/Zw
RFaagpteSmVxniS1UfNbZerOWUhCBmQZXIk1lOF+NTEElpGFWoXjccUwu1fO/HCG
3pCaw6A3SapkIKWJf2IdjZksJOKGGwK2Rfczj2Cp9lnBPvrer4P0JeBnR8TnSb1K
iEfnrT77XcP1uPlYZ57dQwQyaEpxr6aspNGcTZThum5AjLGf9xzMLIly5Y3bW3nG
3BqrLyBCon0gBnSCUilciOjB/YeRrzWMWackrB3NfDdAlBK43bDJmQPG+AMUm0K4
jzhBmrt4PjfgOjl5q3D447R1FQAEhPTVNb8lmVM31NXNgiDhgg+/zy4lOoomGr4Q
Siq/zaKbFe0U4CiwfMYijjXMfAXw0TP/g22QjsOz/pIB72CQe8VGWcFc8pUmiQYN
cGGnX/+DXa4ASlDUdwNYsPCOz8DArUx3/O+b5ujPAC0u0IwgFMpbhujFRmEBa6Pd
iLmwX/XAWLZsMjsExVVVvJbr1V08fLnnNQZ3u87qmBpD1NtfNia56dAEp40BpI87
ZBxhSPoDVJgyaf6ZnCi9Sz6Agu9YTDNATIMUfImCzmXK2SB91Wn60M/awLGc2HPU
bT7JrWAz/0bdmU/eD1sJ005VA2SnfJJZldPFbxF3cakSEKBR48jq/XHcwnhH93Lq
X7NDUEXCihu5hqvv3oKpjR7hy4whNP7vYlRSRlfEbdPvjdIM49wVJLE9/+IjFpML
OndQAQgm9JIipxAMCDGgcyR1aObr0rdDyNbKi9MarndBK15bi/xfPuyF8/KF//oj
HZf/4/u6J4tWNmKW8gEcUGf5IOqjJ1EyIC6IKyyW3ERjAgVITYJSZJreJSJ8YpzO
9rSlx2z/xKOp9M7eOL4lDKgHZ0pQUNdLnJ7heOP1ZiyoBdljnpl3hFklQTevIOaL
v8Jtrynn2fzb3jmFomt3jRIlj6Ga5ZDR7HHBlHX2fORWHGo4Z/wm+EEkoyetkJYj
IOUbiwx/OHOju8NHsN8gTQ2FLIy+0Ic3olmfRf6KHEZeys1hsVJa/x2kBhkNSBBU
nPM135dVGhiNV7wxA35LsD2GQeZ7tjXLBjboavRiF4O1uTD6dPu3PeDNPZhY5xhf
gqKaYVICES0Z9Rxze9Yi23KayrIdcJTKVYRSxEe+HLo5JZxXMfQtMb+5IiDm6i4E
IubSTCBwJ8uUiDi1S/m6uRzMxMh1idXMUkXlTfythlLW55XP20FJP4R+eDccPasH
16BNzUIfX5EcUwSiEkcQphRsjxXNLJqVhAyn4Hqn0vgrLaDrTE5zzd7jYj02fcOO
vtjm199Rnh7vgmyxFpbuyVKTKQKT/d5EHycgH1ZvvofZqSe03fshA1PDrSsxIw0G
GSfyPc0RgfR7/9dOWASelHkSvEa4BhFMeDfpAf+6GKwh8dLOj/pe/fBnUSGyJJ8h
r5ytQfmsfJZrR2NMUMt5Mv6FbTHwnVQ6YK0r3mDHKD+TbkLVqXbMF0gcLfax1zrm
ftJVqg48Vs/UuMH5MZoecOJsxTFXV4x8hW+d7UeVgNztq2Agx6DWT2P/MmPg8heC
ncq6SDcKqWRadDTDebN//UeHCgQ7tx17/l9D00BNEAiSNARYcF3pBUxhSl+sl+fv
NA5Wn5z1aXS4lcqJ+WyDvyGXSyMlUnbZKSbtb3SANT2AA9BxoXizrf0kkp419B37
wFCi/qnCgAyGbY8eO+lrV6eehGlrZEeEn28chvSI53iUpC9Kh+NBGdDHyA/YC4j/
hsP+fs2vwNvw9z2b8CUZwnbEwrV6VXTSGDvBNKpvaeDSqtmNfS77zzkhuxq34FMs
a4lERFeiiqRls8qwgbC2ApcCAC5GtOhbI5CedejYkjoqCrPiX6V7SyK1frHMu8ed
ROkn1MIgF6T0ldgGCtAG4AAMoLeoLZkI5VjxnpOSkxSvS2BRufZkQXRD1ZBgxW4D
m1smo+SV18iZ8xskeqQYdXzkZWugS2gQLBGRgt4JxwKkP2dNZ8V1BZPq4tsx5fAf
qWj94tdglKVwFmYmzj31/+VZHIO1E13q17lpryb3+rCYz52KT96QWNUdy0DxDrMB
jsXUGCtPNiBVOyddOnc/jUF3bNfP9TJaX0Z6EWDwUBCoxFXmvjR99cKWFgT7sZZ9
BDAFrZax7TpvcHCMAvg2paXF4L0hoAmqo8gnqYxU4K+uKgXr4kI18nSh3Ui+g1/E
GpQXKhyc4uorF0gK/eRsvW1VEUq/N/i7EoHTyuLMh6K0gVqnnlbZgtJz9Khf2S7K
hGjXnzyZAZhK3tGDrTNMvwoOEkP9C8s8dhj/tJ8NuL7c5TJDKeaYIE/DqPSmAuPE
VmpldZtXn8LPmshpFGxAej3bib0I8TER1XAy0zc/sOVGY9A062V+f/37Nin4xHqf
DgkTU7SpGAVCmN2gO87U6ny0/xHefbbQbNUxl7FbgadmduP++GHqenEEzI/W8/AI
TEpv76L8IHU1z2EDddJjp3aqEKm3mPKZhHjTzOnzF6agMttwNFletYz/dZubMjgY
HYLzE2FTvydRUDIwKJ4PGvSs1Tfo5QUFb+Swz1dVc4CA49en4ZeZTuEOVSYCofe9
MDo7Ia6LGYU9bFDpH0NJO1IqUcpuYDtVzDr7Nv4jy48AO5SldRIkwOy+Fnz0wQ2W
v4wGmXZ6BkTUnlEczZ02kA6CDN6cZR/A9G/uaGrAXgIbtdz2DEbNnvhhSEUt5qtn
5hWM6I3dXv1Tzt0ch7h/fa9sjobmwgA7ec1W/ObfZHbRsayUmZ5YXrRkG3t6Ndlw
UPifXI0cA5Ka+hHzeecyZ2fg/0eyrn3uyerBM6PjVR+CLnciISL/PSVzuVPrE1LO
R35crR/0kzOdCoA31nE0XWrh7gwIaPeEuiJ6/3ELNZlaHihgyRh+pv87RVYUmmdV
qK0+sVYuJ5ZRpXeF9WG2A91lVD+24kYUuB0qo1XyV4Lr70KLBcYb7E85z+QkQK2f
kBv+d9KUnJcxjL0Xm5vF3dsPihTx7T8bokp2KKRiASqMIuVBHu2mWlTXKrH71B6v
SxY7XIAKqRVpiPvxN2o+UCRn+mHAU1aXT4RAeAxWrj4zp5BUd55tjRiIT2FJqiIq
/6Bt3v1YVadqQm0JuKOmE0PBHYyPy0zLLNLfEtj+M8Q8kM9AaPBo4zhryTBBhCA5
p8p5B6/CkIDWgV68lWfw+uOdfsFVkrgs5wM+/Vyf25P4CxYyuaxaBQXW/9URj9OY
kr8oCQ5lbhRbuvJ25Fqcs5jlA4AFED11lmS2diqWh2CNDGU7b/6ZcmRuKTmbLy3v
HkxkwjjIfw5wd84pynnOhScmCrJJ+YHVHZ79M4SLjSy7/+yZnaXpt6pwb1Q3h0Yf
dkGr5KwK9bUe6eZl0hpQY7xterCUNMciWVAT/WayOVXcXiHiD+F6mXE8cPbxu32V
smGRY+nk7g/f4HDET6t7BxKrDJsKlp71wun0JATZN+lT6DQVKn92U9FL3OnFTyqf
TC56r3GAFAUFtWTrAc3l8H80whoGKL57hYpvWdoQhQhfzKQCgFA4mRNyqLqqUgIy
L+QluCTefz0A585KyxknvQEkviOYN7nVcTf49ho1XIhEVd1zZzQASLW0m+ZWi2lJ
KbszYE+hF/CxZr654elhNFkIgw6cCrfxC7w0nxSf0O2zwwNit6acqe/O+pcSKjLo
m9J1eXMxfEZTimvZiQPgi03G0teqPGxZUN30SA0Mm9fxcVTryaN5rmIBL4r/rGjY
RINbX/y1iSzwLENXCYAIyVsVFF16no1qBoSFmMVW1V44/94kMUv3mVNg17zFlHMV
b6GAEcj7qU5X3GL+GwlvOFSBrrGSPP9Efdxkk506+1eRN9odcvoP17HK6UEIctKm
vgQJTuCV4OcaQTbejoZk/LmBFJ0sIHTuXAz0iC8PRwRNgRRvjXkwhpNE+DMYuJme
xjGvRhawICSZYsXTqZ/xQiC68/Bga8JmjzugY9Khoyyw2JnbDaDhIDEUl3QTsJqj
Wwks6hiD65E8wWMnc5PihLoyruo6b5zfoMXzi3kM9olcW+PPBg+GyzMDMMp15cHm
w0g/jY+OjBP5zLa0ojMHa7J9iMiVpR7KY5tcig/mHdjjEwOVeXZ2S8+fFTieIJyL
UmxhZ+JSo/Ocr4ungfPS27Nrc7Z+3xaWxDa9OTFzJabwujaVpPAy3ZoMr/keWqHC
Of5kXYlM/Runng7k+f60LxiioVokBRb29dnYHqXJU51kIpFapwcaRnhPas3tTZR4
CvuSXYSMpes3byy0jL2rQ64CL5I9wj2r/Af68+nzmxXbFHg0T25Lj46iDb24ceak
PWIyXJNg3wzSR2qs4q/Eg4yRbdUzoujVXrUy9zVEvoydza3o5w6N+Q5slv8cn19m
H4VfHHqtUmE/a1ZOM9KP0yy9ZZlnA6cBMiRkqkSBS5ogr6CTOdIh8R4sNtyj4t8m
ifoGXewOrksCvnTlP4r+69Puam9hLFmTan/fHBLUvuqElx5lsg50cC+jLR81cvgX
A54ZVRAJ6U7Vyxk7Uyt/Uo0CX7ZiCSwXTfp/QFK8G5mjJ7H20p466A5Ub4sQajQA
2oYKCeC7ooMQ8Akq5bzHClcurMyeoddezbjU+Xup2hEggOe1GwiiAoRA7QgcNR3d
BbkkqGpxY+4s32/LQXjMjFr5F8d+qNSB/1qsGm6sdw0plWnphnFycKPSeiDnQ/wZ
I/FpZhZwNOhyMdNTxnnsk4/MHgkJDXYtxUHAl4aTMV7QVMd1Is5Mf2cq14Ed7+Dc
FTGrV2GNARpS0ogkoNWN9rMIZoxzFCgEHJTUB7U/foIs+QJWg0mmdpoAGIx5PpxE
Ciqt+MlgQs6D0iPHRr9PHyKmgkhlzEsRZ4UH8zmo2/C2zIg2tsc5wi08bwdQd6I3
/RBE3+yvItzEgFEnFsb05e+WWe7u0io5kKjvrgBedtlVi5Xv0WSGyh2PkqmvplsB
NjpmlP/u6eWNU4WlJmFXys2bnloQZ3FD7fC09eeMvUZPjPmjAAPFUt/3zw8kHsDx
2UuOup2WnWsSOgQDs4DIFP+1emkmRggvg2xFMyZP1jEH7Se+qHAB+hawMErOKi8m
OgdGyVL8OFeGGrQ+oAE0ZiYnt+/KR9HjHXw592w0bBimGcPXt1+eGpBXRe3+SRPi
nE8HnZtTpC+Ps05UJmuyv7FmdRpIzmCUpHgOo2LsLU0zpB1qY5UH3TRhAYzbbKhY
UMKUPsoKql79/qldgsMAFQFSHxJp++kvdxkb/3+/EuE434ChlTLF9z0MQh2GDWg3
+9jHAWXtXjgWHbfDRnRzsHbrzY54blV9EXBGNbRIemt6K18iqajEQC5Z7+OCQEEa
fAoQChAvGJ0FtFUH8DQACG4tZO1yqOK5a/OJIBfZ6cuy/E8UVXPiuxbq383nutSL
9iBfMaXaYxhpPSwQJG7jVHY32B57NCzDrmNz/2J1bvPeQXIVw5GkzoJmuLVvZ72Y
jejEQ8jnOXGsb34pxEPxa3Jl8Y1ZayVHwz+vBMMWDEKi1ou2fexJVKAKdVSZzY/4
4OHvY2VhkCliEIxuPgUulnp9AqFt3U9JHUsFGh7QAjq68tnJvHTKdjOvlMnlOHb2
y5Cdc6eSHIRLfwZsu0GS1rAEwyvbfn8P1Uub6yWiiBWN6UsDwMUgBT63VOFX3QKM
kWpprgdhuHNbXcXZYevIzvvMXe6OsVXxJgI+T6zi6wnw9ZsezxnCFE+tf0L0X7Ad
6nb1a5TQSN6hVmP6ESc3lmGCgJDH8a/1MuYr+IMzlCZ+QTB/GTJanR2+FBgiV7/I
wBqmasSU9rhWnkvVVjcjh568znvWn77lzzUR7i4pkrY6EOblOp3t3wcG1186lC8V
IYXrR0RkZtKkbIITZsLjKUlDDx1lKLLvN8+0JfbidCY5GA3yQpRuZlB6YvaG+Nfa
eA6QfoB1QqWYb1RbbhTaOpztKs7yJ4csGVpv7sUboQii5PHujJfwjze0MLaaXSoh
r5TxZa2KyRuZZtoRFpIBkiSfNGXecfCLj/1/KDWrc7duDVhkwPC1jaU7kcGo0I+Q
852Ffsdp3Wq8ppPvdbBxor7osH8a5lSl2NT9iTwHO5PTDa84OP9d9hkQ3ty17jOZ
HjDMeJdTGm/KWm/YzGNbLrRRJmkxOmPjfSqXV6uePn4lqSBkj6qSAZsh2jixN9V9
hRSQoo8TDhShi8zXYNecTxMg2rk7aHEmcgawcXoIcMtOSX2MqlkrigD8chZnb5Il
BDE63sQ0/i3gQy0fqdI0oyndlBtIt6OrLpQTsxlLBaf5IiUj8R1OmGHm+2VINwjk
W8AGLDUxPiNp4qLsn+v54c6wLpA4qKiuiKTizz0GQSu4xa92gkmt5vQiK0QR7ZnA
a2Ykq5XTEHp+Qsw8Fbw5wVIjWnC8MyWMZMntAH4QwCHGiJJwdueUn0L3TJ+Zfj+8
rQ7tdC07aNAgLZXUYg42wQF6Kq30BAhj2X8GlXubTkk67BaycGRHfb3MvpKCMFGF
wI4bFnQLdEYRkZgwA67gBohMsJihfwt98inzyokJtZ7AODm9C5u5XgLoC8cGFE3y
+XhzaM3J1ibsIvqN5hHbcjACKq5eCsLhHSjL1ARh/oVRjD83U/igyRh8DaREIN1d
q7Yq/vO092jTuxwxxhRKdpsxsH2hWk2ExVzYAii2d/n9vmjD6gQDTF1Ue0l7YO6g
+bibWvXBwL1HZ3hascZn6H1/uD9jOiCvgyRDSyRm3OjuaoJF+us0qrwY9Usia039
TeCSWLFvEo344DzSeUF6foK/AQA745hg7NWraoAraEsndBwVq0pkehxhtKd+MxXG
LMCF/oi18Y0yHaZMceIbDsJRykD5vT3m4QaE9sdjir3trd5fmDUwdt+ZzTK06Y0o
pojw6vfP51ODXQyK7Hn240c9R0I2HpYEa2T/TSFjOAbgBRYffaF2uyC8BVReBfzk
c6Ivqj5S+MxbDavloJoNGfkteNZj+ixjh9m854DBzTyhiCJSQVFxYXFaJRIwD6RC
OnF6dRlchYESq3UgZJRJlagO032/H5P/y5vHTIZYH8jvOX4ATKdJcaiOIs0v0pRu
sYjc5/Aeavi4seW5zeXOPKtbBquTCYN0BT4iW8ttsOUZAJSXL+/Up1N1NRS+RKFO
XgrUNLrRY121ipllt1pFU3fJqYOteLUOHYkIUeW/UbTdmcnCNpt0nxiVkfQzVe+H
63FbzXPT3dJScAe6RjLtcU1zSAAhDNsXliqew7/akq8FcF6meFCNkGLlRzdiMcAK
POkCz6Drb6kARAlTr17ViFczOUWWiQDealHx++f5CBA7gt9mSY3xwQ7R6CVsGE5B
YBXEGLpao0snefVgKWmBJAJse1CvJ0IuFGoo2lNfoJaxGPa1URUwQPXxPAq/9yNZ
j5FMhSBVcNuVhFqYvIr0GsA2UW0c+MlJ0uO+BLtGctG+fON28OxxKSsMsPyT2ip8
88ZkXbUxNa21jXarekabszePPSm9Qt6/DDEblmDxzAYYhtdJHYPkzMk//U6yBMt9
mCKV55flYIN91OQm2sKw3RM+vGO+NT1Rz2Z2MUhxHwPt1zNt1wJdPoby4bnFIe9N
gT6/uxUjPjlF9ych3MC1qXekmTCy+tdwm4yglKcJLZ9hziBgp5MqeyYN3xg+vuxA
WOwKFsX2LQYAOqWsYmSFukC4BLXdfdS395n5fsECa3AhFF5R5ntS1CTObqqFi3mo
glWc6dOLHYtF8sEoXxt97Nb70grmmScaS6j3JMKlayA5uTjQLKHYUBUeTUEdoZJU
ClVUrC2rOVthtQ4KUFHtjlN3/M7sjqxW+mXqnAbuatzAFyoe6YeK8B9KefrKrXMp
Ooe6mmktN4oWo6Kk2nYOuZ+Y5yZ+HhEeU+f6XPbBhYN+lvxvHpcLf0bCWI1/XbMJ
Cryi5EDskVXsU8e5W0e7HMIQYbXuKLpEX/c4eIUYGMaOg3my40H7BEaiLO3vMQDN
Fvx66lBu5L3a5WwUB9QMdEgie7uV6r+dTmiuVgsctHnz26nRh7UPt1ckBL2lnvcH
Dkur8rVrgj/QaPJ3qac54lvDjYPQeDJYs4mh8RL27SaMQqDBTCwFVQq9Bn1Kw4BY
RWXpwIr9E9hCnd8Oa9xj1qZVyKjFc6tRtKq3aUU8/BtfZ3ftUCP0mq6QE1DQBJrF
G8cnYKtayWNP3QURPCTvCuqUbT3NU8slzi+0JWJ3VEQFVuiQYiE5c3JZQhCOC+CC
3qn7dgPf6Ym7ZNjnuCJalBBcS7ljnbVckLDBye2oF+35hxI9SZgpBnbKlibvJNxJ
ffeaJOuD1omHVI1LX8BDLKg9GUqiAolu7IzGMy2aawgmOa54QgVPyQkTOxL7Z/d3
jzYrwHpscm65UUNslCdUSJSoDJ8J9sKbsJYA+uwDbA347xTkpGKMuBGjxjgcKQHj
DbYkzhdvshvonfcQP1OrjBWYbLncbor8lPkibtQfITGM9BLzTCB6G3WTMstA5LVD
RuPzJfRce5tZpcI8q4ot/bEysanEIzbTmYWwXl8IgWCsqYVd5YG9MjJl4z6/g296
KT1R2ZEn97mNcxfFlf92IAvOTr/FRM00P7C26v4ukDNrxy2Bi84ncPzEMyt1VDEL
8tbOanuGASmD942YXzQapu8OsKNjwqrvlu+ZTuRyqv9PdJGYJ1N2H2M72TlcIcRi
hR4OHV2kG8k5YWWUiiIpPKZ6vF8fji373fYXTjUg+Vgz7lQzuPsybm6ytKdncuJ3
S21z0rYVxUSKW8YR+ZACntwi0JM9jIs/45opRYhyOHKL0BeNxZiwl3wxGbwcxkUT
DV1bJUJXNeezeUAZJli9mFRKXCJR5gMbwDxekJOeTMLm8+Mu/2U0GK+7a+jlj60l
qdhembH1Vf4KOi3UalugmkJoQ3QsQdJ449WJp8EEk0LohVclmAZDCnWJnc2jXEHM
JwCNtDiecJxlWhY2UUJh1DkrQuHapJ+2IihupiSrlKTmEEf7bJE4BcLnbo16+WhX
y0jzoDtHJNYuSx8cHXevDEFr5IycZkJt8fNkMNPu+PXcn++vhJV5Mo5GPz3WJbuu
aLLY5MQ0EVMaDxZ3p3L2OpIy+pa0zRh10C4PEMQ24v48ZB3bidODrp8Du2bjf5eq
6vcjGS1GN4iR+tT7yYdSvU1ZzGNkHM5BIk3gYDVRlTeUwE3/IFPfb0tf3PqH11Rr
sz4u3BBPz9qCaQ1A/X8HI73l8GeTHJi8Yh3D+jFlxpu3f7LAwj/73tUoZwPVejc4
48kDhnnd3WHYmnsVtrwLiMXIc/oN7DCLC/Hmtttyr+TjSubna2USi2qy1WjtmTjs
6t64WTheCWtzAhl/l0ugQq+k/mNrVCec1FNH4zsEd+eJ9+lLp53QxDJj2lAP9CRa
a6GNaHInAIgOMxBdX1gkIYrsv4Kmo583VoMyQ1vfyrdenEqTJQl1RLvx3ivcrp8P
dD2BLbOHfk2x59oEdROFXXkf0SDxKg6uSCeLAzsYVD1LNmb9b7OIO4LQMVSExZIH
2IpBVvBasTk40zV805aQT6DM3BNRPwR+ZIf3n6LBTurHg9USOvsnOkX79SeWMbJF
vZoV+J2oazbyPajsNhL2iQtUcc7LnbTShkC66ZNqiz+OhMFyg7l7XEurcv7jPBKr
uwkmD4JpE6JVpcVoytZHo1SnjkdktjhRJbwISvQWkzjcZXgqDr98j/T9M+2OO64N
5neM9SkuRO03JXmkYf5KVgS4JlQNjnDEmA8aQTwUobCzNUom7LYrAHUl5DbUaCBM
1BfqJf7Ip458rwsWABYVW3weiol75C8Zz1E/O7KbdVCXEkbaP2mt3QLi4lJDe4XQ
6sjyFPR+UNtwBcz+1XhV3lph4E9d5e0+QXAtZMJyWvPCKvQJAG/p5/5t8PwH9QyC
RidwJVJU0U/n37/7D23HJoKcsY0PaWAVb4nSl4Jnr/E08NhmG8lRIbEWxtincY1X
ZWoUSFgrHL5hcZy09bJNoScWWBFNCAQaX1icrUiwNdpp/a5M3Mr0Aii2YzflNlab
x3Jbs+REIBTdP+Ii/6WfxYA1AprWO7s7qoXaEEgBbD/a69NIGGIsnGur9hkvXKeL
lQ+FkuNwfO39ZkWxouMrZCpYfphjgdIXcMqNZIEgtUPIFDWlwzUrsfvWTd0efvfW
iNF5cxAF8cjJKAaUaQIheVNmt2itM9yVOQdIwQldP/mdd0JmLOhniWOlfAal0m9l
vShZfZnPMDvN9NwTQBn6+ct59z2ncyucqDbxChS290neBMSrO4hz2RRF6Dvg/Cn1
k/ofO7LSzir66G/6gyohkwyd/G4NErI0L5L4oAP0X8jnhNPd54C9PdqxfFmV9exr
QmBIbEiksDSkum4kxkTAiHrCBlLXgRROWrsKDTwdAjREba0apJbxFNC596BAfLub
cs9iP+VKpuwEbC4z/z62zR1Uim3yMU8XgQOQmkporh+fLRAQWn7mCAlr2valklin
/1Qh5RmPQCgvckRb1B232TUUwY16y5h4QE0eouc5rmWIwQFOV60DXTPWLzP5ww3i
QLTLxRa9xgz/SWaRVbMXOX56C48WjcEWaJLOswOQspdXnwVQiM6IIGFnPiyNaAp8
YCVT118EOQysRYfz6Dq6BVykpcnLXX3MAq0BThEN6hd9YKHgN9EY4x3/jP8PEq6T
IVkf4WV50NaLz0t8zhAu3WPOqEhlZaM2rCqWUP2gZrWS8Tm/+ogExmOlm9z9Gh3O
iePnny8zkfJcJSHCm5jrE80W1voX4LDyoq3c4qtOdDib6rpOwwWTyrIe8s1wnRV+
RnYQpq1dw9HjgSYqRSWHG2vttnFBSdphm2jODgUW3NmoJmw1/7LC98YG6SIrLGFf
1IuxIlhecnZuxlK3qlqZWqC5YCFvnFP8Umb4+xEUGkOGPRWgzKY74J/9JZsk9y3D
vfTAx+x4j0G4qzdQQMcpc81Fz5ABo4tCIrq7sqpdludzswmoSUKyLrj7IHvTakUP
zGRpvoeRpQGxMbZdTjvp+hvh2z1wZdz2FDSMurI2AtiFd2T2RHX6gl0FUpyaWmRX
St22a1bn0Lcu71g0VoQYuZsVI6Qy0yaw5iCQphtuEl899tLAycLpi24Rkz+fHucs
+yPOrmGKp1WiteRFujfK+XO1+4DYIPZN4VVBYx+WwOIQzn+wQ+2ny6LCtbrzoZvs
KdxEGJMacZHrThjCGjIxP2cMYRT7+9CkrKWKYhgDr4ptMLZ+IRi+EtZG0rintqCw
iLWa0xxIBfl3xEta6auXM+pmxgWHLTYpgSkX4L/7C9ebXvAD72kO97PMPmcN+vE7
ZC5vFzDxAgRcWD6/c89GoPbM5HB289kZzLXy+TR/ScFz6Dp77m78XIxNMxZo+OZ5
ZFTtCEgPxZkys/q1PuFyXA6W2n0TaajSyr2HxctRXLXLXBqXf4eGVHL1qLxAYFGu
nruX8b0cBgab+286RxwiVMCv5SA7LThNizI+AYzg0IFq4/UrpsKmOPVPmriTubdn
MPErPhVKBRg6wAndixwROkpxXOfq26rb5NplcaNC2cqJRnia1e2u4cKCOHb67fyl
LazyfYYKcJOd0k9fD+BllBKZ8shlFjoYpt5KEg1HQRATGFPUAHgMgxD/AmzUyLTE
9M62dUQLjP1sXy4pdqYBZYXAIWcKs/C1VHB8uO1dBKRliVmhQt1Ld/tRPu/wFGWi
YB5+lShOBzIIAc+Tan2r9LjCl+etLCg6coLmr64LUB/RooN5h7nmQy3XUYWWMQ1X
KJIdvKTaecE4XdhKuRcGYtEUiJZVMNMqhNfiMz3Jv0YD3VzMgMmZb2Sq+yoDULOl
bUNm3qUL+DJvUOmys8npFYs/QSUiwMPjjJ2OzEmPDEv+IiL++CVnpdbkLbcUt0Ov
IDMuPi0IskJX6oAA4Aat8m26FgLyFPUpt3S5qiWcakHpEmQZvM+h4wQN/64GjhMF
9p641+6VlGvyxAH8lwCjiGq2afFWaYyKaCetVNdI+IjZ5fXDcFF/DoSR7eSkEaOj
kj9ESm47fQc+G0oGtFRI7RFzQcGIYUMQOuzKajYOLFHl+4Xd0SoqFdljoWdpqyrO
ZaDkcLR/+u/TIlh6Ct6BsTaaC3Im4UAqX9JqEd2NTch3K+aISsKRiEUrIFBulPFF
tJVIGzGgtVNfPj/26MKfehH8VfxyRwLxcQkKpGVD/V5oBLLPkwvByvXEgJ+Gv2Gt
pc4Pc5XMI8VKVX/yGZxKcPvu5SN7NE6+mY1IfmiUcTP+ui+ZK+OXHi+Rk5YmLrG4
MRM3rIxuYJc/9GDZOfBvxvmuS8VKohLQ/amLRFCVeybrvxdWhf7qjcrRkb00c093
SMLVLmvE9QHPzfL8q64OeR6amv3q8SoSLH/9xDBb+ap6kZ7j4UcPaZTfDc3h8i+i
9oUYt7j7Xc6nC3MJjzhXKiQobm03CNjOa8WIa3rsgYISjr2bOflvS9LJI1+Pab/o
wYfjK/eE1D3pTK4sYsGex9DP1qeXc9uX52k/aweu7lGwEeXuJV0b6y70yvwDlf3F
OWGv4/x5GMoh88Ql9O2vLz1WEoGzrjg6fixk0hWnxOGihYeBL01c4vuA22uP8gL7
JG+6qkR0FLaKq40GTlofIThm8fszLz86/VghEEK1uD9tr5MLyXJbiN8lSgDfegrj
F/Em+7QmeV6ADO8Xi/wyNa59Ynz5+qtto7j/4Z5SmTnksB9e6wXE5jkpi2BwZcjG
hpvt62NQVqmJs52IBb93NF5fevuB4MSJRVhEt0zpQgEsxgylnlkc5JNFPf/yjw5L
Vnxce8BOS0pmvEIyyk0IY0rZX3FiFTglbptRl6J+92EBmhwv4o2eC9MfuUTMPIaT
I8m847vSzo5ItvA4lo6u3H++4Zg5uFPJTwphrzjkTXcKFUmgZsmDeUz4Pra2GcaA
gJunbfc+qDdlQ8qsZGTdQDVFauhByGxcPTtcpF+RKcc6MPUAId7/Ebrt29/FoKb+
FO5A/BampHFZeM8Fsm5GWEvHNe1YgUlxlCu199GT85AFKrUz8aQftr1b+MSPd4ms
VxtD9Drasht5tn0ZpVXrBLWpJebI/dcR3KfmRUZ934W6Xm8PPIITUMgzFg3ZVKpJ
brFvyfsRU/VIJhIU+zZ74B1gb7B+tw3abPeT8XrlM3HlE2IiqbbGuKtZVelevaej
Jo5GVoWY0BoLtRHDf3tTvrrUHHOL+DN5yS4ByiSvPZOGMWVy4blLpR/kBthQsFPi
Ue6uzKBXZGLVxExiAJsWKEO3ng/d32kX5XV6uzvK9u76Wp5oDmKb1/t4kOcnRy/d
05eBFouXei+jzdY52DlxN3rAFZ7T2Xjw1VsHSUdKimdeQ91IHMsEgOQ5SahJ90V7
7tr5NjOykTYZHhMFxhvjtR0+BhjjH29TiojE/W1/FEEBpMuQrKOoi0OXIGm8P10w
GOg6/JxmTT/ALcNnsDaA3YkzETxzzH+MyaN+xiAgyVVEllm7q04GYcOLqdeN6QQk
UNUxWII8SqXck8v+t4n5z2gnq+YZVrV481qK6JYx5USSmqG2BnqSbN6ccP/bqe3h
sL7pBKJ8oG7OGUYOXyRNffTikV/9OZZAHou3PDbfy8IIQyyrkdMiIp6bHHtawXKV
R70krjnz+FZ2K0s4F5B6nct8LlLb5qSD4X36Q3Un8SrOssy1Gwg5eZ1Pv5PpySXX
VQjL14Ben+k1zVa21FXDrxNCzYDyLUDlZ8Y5xjkMSwC2wQmdI5RLxN50ZOLw0ghK
8spb0HHuRmNhkMofmR70uo1WNkNxBld1QmFBdtZI9kI/cHVbbXUbb8QZtOXSSM3f
ChoNtURqbkYDQIloYrt4GIWl9DUX9zpY6yc/YRgUHPMF8I+FiJ8xXp/zXF36jjs2
4TVXdsh6PXWorvYhXuVvwMuwdZosI4966+xXBpcKZI5ucLsyMNRKD6rzwBwJsOMC
FN6qTh+DnqN4DKaQpvDBLa9SwF9x7pna3HyQz3CxqIz3b5dqbRX0FDNMPfl2zjdJ
7roGAxEr9fTZeMBnSDGO91THaDSmQ92+1NiJFJJJyXn+VETW68D0DcokL0Mm9BO7
9FP6wrSoklh9IhmawAOoKTH+vbEUOOk4C33uqQdveyb5CXgHOoRCJQ3lPtgj8QRd
94L4tV/lpJPkbln/P6BVDi7Zug3baEDHtO0YNWWCEgwAR2WfCqZX84J+HFI1EaCi
ovC/H0JMrc2btPkAopuBhqmCr7zpCkr10gOt9KT3GrCGO5GFb4iF7LQ1tmkP0dFt
DEjay9iYBw7YC3HGBJB+rLTGr1vxRjie+5J3aNMbZ8FFoQprdjwJFW8LpY1Y9CIp
jf13bZTr+rB1QKlb3y2vvl1P3pGQsvjPu4lM3yXX+kAToK3qB9KurtCgoqILgTtf
ZZP06n+pgI+la0G1LJTb/nVKNqgUVTrzHZmIuSwQFo2UgA9ucJyhnt6uA/JGDKlh
AFw67c7Zv25n3iVgIZanka0NUFjaVuaqhB0KwHwTAayziibak7oAvsUHtOJ4/MMk
ShGFb2sNlJDZCUTlXTcR2ujJd4coIbR82FmnX1dNgNTMnk7F3OxI1mBKBanlfnmQ
Cj9niBEV3I+cS1PLBJSwIBmuMnMVvmbU5jW+13B/OilRxFJLVPOufiuCcZj97RZ9
QlEhJUm3bNY9VylW9WSijtfkJZbnkPf6lzpHf00tpccfsa1T3UQRTswZGZprbVxF
0/sseDPeA3L/syWzvjmspx6Nz8pEY4z3LBDgpA7FbkwHHQ0eMcns3t1KOvGOHAdr
/pR0KrnbrMSHdmecPukjBr4549c5k14qZBGyTi80RRuwpBi7W1fATTlwWOVb3kpF
z/ReHQ6roE3QFZRah3ZfX+3iB24LLwGRbVup1Qqs+GEnRQrUyQn1yCmIm4K9Wbp4
/2j3/tIL7ZDA3eAuZUJRrFTDj6FOSw08woF3LnZUU10ZFiYhdOEK5q/770HuFgwG
AUS9w12+pPfqoCvjCmBz0IZ7tfLOaz/g77tTotr8WhBUNDwOzpw45MyvavMdei5e
30qbdhrNBQe5igRA3DfLet2QvSZa+fw9pgHE6uxoSekEvoOjhk/g6+KZc3Nk1tCz
87PNaIQadGOIvUCii91q9diqnvNaKNTgv83GhsUo8bNnXZIwn8IwOx7jcGlf198s
ADadN17QPaqEiu4cDPbiXJi+thZYrcoyLskAUM/9T2tSYm054iEb4PJfEJCsVq1B
IpwjPe+WvgaE5r0NJ5J8JsQyB73cLcSlEJu2UHUO8EDhsnAkV7ioPL/vaSxzAMpl
AB/E2uqpz6cITa0y2BfAzbzmKdCMUGe9QwTyJX+ryfxdaDeYktmHfAbQSQga6Gh3
x4xczFZrKjdYyAKqo+EcOMCP88t2YubVi3xIJD6j933YT/UkfGQEOLXx0Y7V+A3s
8hVHvqVoUIPOT73rbXUIR/inX07zk3xJ6qiWMGGx6NcchhqRlboP/EewO5oDG3/u
etQjEg3kntcCCkj/Nd+UyOu34/A7JXc8WVpc2LpPhvuvGh01RrXpr45gjWctJeu2
MEHnoPw6Ni74QjK1ZaDKCnBgx1PK8w33sKUs8cHgSBkM7aUBqBy3oTWA5GRdlS2F
DzIyMoSBlUAZ4lYF/fqGmT71w0WGBiyCNn+sygOJeO0q4yyPzfgPvMmd0xva+TK1
egpRQg2ZqdP9vFTSb9qIB1w8nKUmSDCvY6gYIEpMV5s0REdMwBDiTNcZjad4Carz
H6Y+lN+UJ9AyAVAmSLjxB4IGpEa5AjHrjVNMdEXNv4EGsSRTw337dcg+7Fp4fLJb
EpczUvBNuDrbDiWv7327DKHRfJoxtAXUAISh1AreN2z2Wzfj6dZdOOzgPlxvyZr7
G39zInwpiz6jyoRnJcUXWN82VZpzw8Y9sYHK5mkTaHEpDRRSWH7TYQFoGNdBc1b+
TboUfs//jbovGekXbtHZTMioZN420xhMUPhnApJBa3KQ126/4AOxtOU1ghjv5rUV
l0K+8zLjJ/sB5nzMrzM5PQa6ajlMQqhzq2m5AVwbsdJBQVAr2yipH1LyplJD3Jue
zaHKW0tfg1/YUTSpjQ1qAa6AZBxoZAKFmKdtFjNu1lZr/KWrHLZBn8sgD5guHMy1
yNZl7j/XLuPhFzNcu+8A/sGbisjnTYgzulaUSdhYH5gE9ba3kFEiTe3EZuF10Qco
NfJA+DrJHF+Izhtgu96N1dJls1MWqUQXvMZ3SIFJ73lrAuzZh72rB3bqHwezNmIJ
JqgSK0Y2VJmrOoh/rVEIYBEcm/X5ez8fIPOVT/6dlSfb3cQxh34/PJ4NFL/P0OBK
IeNiAGf0/vzTHD+R44nuF5Q6/nZtax6c0xmYyTsPYTviy8YgL5/+lL+Gin9u6gjS
qzGD8/klpi870zZ6kaxZkceH+XPxYy6bzmWkjXSMzrnErnlbn7aHrsdGd+dkxGCT
AlCVxVQA+77+IVUURkwgHXPBsgcwGLmr7eRQuHDzvu5s4tBcca0MHL8O4+W5b6tH
LLlQ6rQjh5X0aFL4TPdB6fs+9aI1ANSp4KN5OcCLQya7pZym+9bG+8SPTSG4oW0g
Lx05giaM64aJOp9UrX/IWch+J6WjRxgvt4CwOEePHWLm2rYcDDZb6tug2qfObSO2
ZUnpvVraPxlDc750c+NDiQv7CXo6fNIveX9k1rjPIdct792/zEBdgsFzX0Cn3phP
OM7VTi4Cfa2Sc6KewSusOICePv6Qm8JC6gtG64HQklsxlLYON/gtfutlhlqEn9oE
zwC71GcVqkfqnOeXj03NZoMm6LEvrq1MvMe1FOLsEBlZ6XV3/TCo29oyE4gyCW+5
O0O8LHLkamhKvOozJXZcAkq0psDC4iP5LWPCE0dmLg7EnInc8KK4OlDgs7G+NLdz
aBkof5TuMsvDL8hybOAU7WqKouUGJihFEU3YUht4Yf+kYycoFx/h0glVLOAdKsD1
D2POcRHpEtlv1kIP65N2mRG0vAk71dfItDKBbOgh98qvrWJ0mtHpgQfaxW9RjYPJ
AP0ft/V2YTcRnv6DpMnEl9N8FmbN3/piDZVHqR1zKYK365CiOS17zs++ZMKzjoV/
Jsg8DFtfcPFTMSr/+cmFGIAhkRjwNl83pucpnwCuWBWBDwW7uELdXSqkB81lwA2h
VQ0yJV7uImQ3NKFvwm5O4OowSozRvMnlywOYz+D/l/HfZ0uVVA4RnnUn0U7v7myb
zPRPHVecLJnBNineWv1kjVie0p28SLicYBrAUKS1khCJKAPJROqIwgQOn5IcyVhC
aWwbNoMkcpj+RCa9hvKRoU5JF1uCbY4HQVNN69FGorPPcEDzidfSrgeOm21ZyWmY
qt0+jrX7g79Ta6J+ajxdQwPESYKYDY3FYRE/yV5xrCWcpXH9Opoa3IzLXZZtKEWW
mQbwkw6BC6E7hhAsTXCnyQUZrNmDNP8vEHfMPoaewr+M3hrXM7bxRTyH3fea05CQ
jSvJINYPLzvSOZH9llzm2dWTPHwsWyKRCmuo4wWVx34LuVFSPqMcU1aowktlfbCO
hbHEC9hr1yQuBWv2OPkZO2kp8ErAeV/ClpPfPwbKqVokZRtCxCyVZUM2T1XVhdKv
G27UfVYjOnNwocH1ZhZbqq1REcqDbNKOqFijfXoeh1t5dri9PDA1z81R/X0bibXq
3QeQliZ47cbOewmu07FeY8egiCZuXPz1TxFBl8EzZakal64FvL0snQ671aABr22j
yznzal+jgfc47HrNPt84KY/+QPFUPkUfXd5JXs613bWYoQx5s/wcv4aWDGGV0scr
nv0r2jugf5206fxyGMCAMMXwYJvENsVcmr3IFjxlFjr2G6spKjPyvGKqzD+eZeLB
xx9Kn2BaTjx3wci96LRkzLq3noSHtVFBCjQI70FR6yhZkUyPd5lWzyQqJmqlNn/b
rHcxCVAMVh7hl7/JPMWwW5wkYSVP/dhjXg5hAvlIShf3KioENy8I+dvkyUg00mee
K8jPAQJY1sZQcJmJB71dBfcBO/gB6AfUPrw72dFSNykUmoOkSmN2jukRUTz5/IWf
RgwZzGZIsYVv8+qD79m0qQzkptZ3EyLny2X/+xQRQtBTIwkeZkkSj5dFLyQhwmvk
SD6QmSzlRC8HoWwWEvTtW3c1ZI2Bglli0RECHKBw1eS0ts2jr8B4/4112IIniBmR
9QGgLzxBJPgu6rMtstosDcDg1eoVxRcuivV6dk3VyK4tK24NHWC+cACeqy7KEvlU
P66lp4Ep064rqDHSJwwLR1liM9TJv2q2CMIx/xAdSLh39n0Kqa9HD8B3KL/EzzMA
ea/L9uK5BxaYIfSPHvYWwv8kBY37aKOurl6vILS6z8OsvaWGUFItDQ6fD+LjVZlP
iYv7Go/PJR6RBLjMWIFwlvbCS9Jih4r4mBwBBpQAN1cxQVZMF9/GOLUfm/0r+mwD
Y5wZBXG4lbo0a4xqUv2o+geE2yKzl56sVM0cOz8yOjYbJGNZiGAfEJvzfpaBa0ev
7i6Ih91TZ1Mo3+9PNdwcj/8KeLG+taq5Lr2dNxZq+/YpWYV03/XgQ+LxDTnHO/Lr
iR6TTzeK3kz8Htc1pq73mCQphW7STozacvW4ZWDTUU3btN4KvwbXmFpcPxtDb8TO
Rj8PKCABJgiglgfgT1KS6XwUEV1iNIjlP13nBaW83eHxklrIL7yCn5CfcfZyt3pV
wJUESv4CEGzJCCF2PrTE94wqODLazTLtq0JQFhoGGvyTZIsaQLt283LovXjQsXZ5
zQXu4TpusY640qHZNyI/3rJe9hj/ASuOk1VB+4eFYkYofLBBF6zhyLp8C6+uYXt2
FwFkA6COLfJIZtW/NLbcy/Y6B6kzgRcNn32p2TyHCPBMzdwH78SIFfZw4FItA0Oj
dwel9+nf39UiH5QR0q7sGK5ZE/74ZzjTXcACQa+bHuWy0Ov/i9SdfgfUePCtAKJp
C7SFQjVFQcHbb9PikwY/UcpIt/4MTz9l7VQkMrm5JEQKsQZemZkRmM7vQNxJ1SoT
aw/sf12/CYaysdMt69AzkATGt9QeLWmT7DBGh0ioRC5EpizrBKcgdvi0Smo1P6BQ
5LKSbV47lSb/vTOc3azDcxtD8ZGELCoiqItBaVLSL3ISly3f6W0hRUuGaqqwZ/fk
ZjtwZA+r60jD3oAWVdOJ1aqj6WhFQ07zZAKWsgDf+ZfV9K+CcfjvIlFi2+iST+Kg
cYMdRWcimTtiLBxo6c6o8x2bV9tau+SPlxVmX4wpdtZ5bpFSJBAuFUSsCD76OdQV
u9VC2crQaXcvSXqKvW3YYN04X0FUzCbgMF4hKpVijFNdccYD1EpbjP1FheKFHL33
gJnrik7u1Rffhn/8o4A5vwY/4/a2sNJkgjBSFAlnnd5hLbJy2jyRE0u2CgDATDq4
eG4PjI7Wny+35vpmSSOz8E6jt/5nlxhcnh9rSc/s+qPAK9XdMber5kD/I8PVPMn2
QhwE0Ki0jyM9nxRRe+59cyl8T+Jb75RY+BCNsYu2pW7NgLSTQQBKChoBm/igxMhd
iGI5dmwrtqB2/VMpL6qe/5Y723v8TZm4NezSOmRhXmQ+brbOy0dNsFSXtYfhEY0K
+I7G21gzweFrsmlhQGBXeMLb0SapIQyZgporxtVFT9N7xeM2dSjSsZu4efOvfpkd
JB3DbwYVTh6OOcvveT28G4ySC6QzKx2CgYlHvdSAX5hXgo+QmC2Gvnw2lUOHrPvB
GDFJokSZJuqXyAl/08PAeo++wYoD2d0oyEYp0zHUJAqfC+4RAfiKjzOv2nlgNzmw
dg4XcvnmZtZdhgSOT2TtJ5Y/5CKhPHL+SJ4vhntzGOgnuUzHhbqnVjP/uHqLREe3
VFkywA2CUtmvG8YpHh2K8P/NmNm8qn5q4jNxtxJb7T82RhCBe2LUn+n/RHtpVE/+
lYsCYCqDXEuLcTSkxscKqdB/cjaUqGqmFJ1QAy5Tv3b9LtOlqvatIRfdrtRxjzOI
jba3igWhR45nrlghcgd26jJ1doXB7a7UjohvP5aOTBphg9XY7YErP2LYh9A8RQgh
64fRof7ATPr4JQH3IYlF05bQrevOmMdya9Rjc/TIEmWqqg9Ki8REK1Kn+NXVFPqv
i7dTrRO1aTjqrNB/Zg3vdL/KITs8Ncow1gnlZiHmToAhyTIUdvZpEv26gGcL8vCr
vLlAQkXvRNxCjS+lZt8o1xA7Lv++WdJSjZrgO4hbMkqfjqlkCUJ7cWfp821dRTpW
Sj4vPWUdNMWNovzmJ7APY955zNgpMDKcfyYGpx7IUDe0EjEDZcTXMOsm8V5HW/Dh
a1yqSwvcbE50oPsSIk9mDFSFHc6kEd13u6b6WjSPkwCV35V+ycjzefSy/vzSBX0Z
Ba9552f/rFnV3jg8d2bBc0OWtY+z4O55Ujqhp0oWBx0OLRtYFxiwlRd/kUwU7aWy
1uZqC8nA8TK4LU2+r73WntwGfDYhuJonQubDJdjw7IuKc2EsF9O3d4puGr0MuqPB
p3BnTC+AQpg66+10zvAdY43CvbBq0jQaVusrcSsJ3dU4xSnoyF/sVz9uFP1250hk
FyuClElAZQTVfrLSP++qOmYVIoAIIcOBTXH2ftClCrs9Lr01VUEDNbZnMc92sHbU
w5wiBMJK0r/rFp689BapY9YHyhIWqDSef+KGcmFVt5gsIQkuygMDSyRyTRRXulHE
Rd12uIBUVEg0xAw8HjIXawY0VRU4so1/2F6tX7DHhzDdqAhHtnHe8bUUCzxPG1Zs
r3PI5/eHhGr1ieqPgZxY4IyxxJy/OMiOgnwCmZl9cwll8ATaDmZBUHYrYVHpc2KF
SjJIXXcWgk3ijWty5WW6YbByK8+Rcz+HGaz3BVAaF65Czs5dnEQrBR4uUunoL0Il
NN1CXwVncMaBKFpNjPi9POJB0hem6EwoQ43hH6vDwM8aPZgv+Xvv0Y8o+iK4JF0A
U2wPRkRP1Ojhs4ADH0dy5aXi/gofPCctU0tm6v1XFiIpuo92/qJRIbjzN5oWgXKh
zr2WtSIsGoPWivvkQGjn8HPnOeywR+iF+E1xAw0I4+/9EjGw/wPcQMK16yGdIBXz
4Hl2ZfxoOEqLiEVjUg0rnEC5BWV53SLfeBDqvaVDCNcJNgqecnpMo/2D5wxs7RBo
je0H6tXVwbhITfTkokhoAayzzlwzmVROXzLYCKFbtC4+TgQGOLur64gTaQoappGD
h3pNZimgNYdCFIAdUjy4BbzncpqSB8YcDaLp/91gAGY1FBw0kKlmAPI+XflLaEKI
Jz74/hDBa+22MCDg9+kFKmQwND3IbVuDJtYlMWDspgffRw8Sg1MjDGYz5KFXx2bV
ngfOoRHHDcxhCk7BJZLiZX8Thykd+O56ZmHJAbfOJtzRBqWP5p4FNby5ZsvDrNnA
d8TZSdyCkx7urJzdP4MQXH00jP9lFolQpw12Ytx6HsTIImRY3zKqUwdx3QFHYVGK
v/vgEf7VOSA7owUM0UzemGYHv3mcLReW6fR/OllvzppRkDcSbWVvxW17/qUjxUSk
IfIRu1iogmJAxH5VzUfInIme1gNw7EZXBPUETtABy/cKAYV/FwSkfP1LX6XsdyfC
vJlJAHLxOLLiRbunfHigYLipYpd5hXvIXyI4DM9IltwgRDX0X24EcXF/Z974+yjn
WEwgsYlsEVOVx9mSIAhOvc2nCxS/4glmfViEdLr7gfNvvB9WJ8uK9Jlq9kEpUvrz
2bvhYt45RcoshIBHI9LkKeBbOTlQZg2wLOFmesi6XwmxzcUO7gaZ1l/A/WwQpgTb
XKf/xCEIQW13RTHGfJzxapVA3O8fJCetuVBdNtoDGc90qH7CFzxrHId1S50jqnx7
I8KbgbkeCTqXmE9rHT4765keTOE0QbIMO43Y+2CB6jxjtOD8sHk9D5SIYvn1hhjJ
C/H6qV9eRJ7o/UZgX3DE0J25APiMdTFBLeNyMMlOAnLIfF5WCfSPnqlrbXspLSOh
4Nc1pXd20R65RR1eTO5hf1iPL9eh9hqC+bR3b83p0zcrmYMcvybT5b7puA9JJbWR
aNRwXEbkI9gdva1sArHR8gzsAKGHUOGOCYbzkL1FrqiDbnOlowKWR+TcW5uNeNa6
Ziq9D7j7JpUkVb2MguB9RzjZEZtNXN2hVpyTSRjlEW+hmWuqM4c8LEWDuWLHDBbl
vPyGstBtHX3URcpKdME1evyzk6xaZXOP/JM9RgsPItL1t8hc33UbSTwrM41rQPI0
6tQSmlH6xf4NWRAiGwMcUfcZo8j3uq9U5BWymCksEQgP1fY5mamNwI9fhzbYBxC7
57o4e1PxE0owYFUidroZ7/IbQwF6q5XYdu3+suEapmab5wfxFXqp5g0dQVz4wuMm
Tf2HOxZxsXRaXlfH5a82horqY17mPkgbDycOZgvTTgXlfvYe1hGZbZHWqgeRe8OO
VTjaTqIJmGXwjkubLmdQgXJw/cSwBHqxOyHvwScHbonPB2snh46fTAwQOU67Xaoi
+wSogH1S+RftL35Por61+llXeAwtH5xR8Cmlvhd9nZ3ul+DEItBPpWHUlSIoyQO8
HYz/aGrhC0WlMTO3vj7E/nYmXATh/YYV7/Hx7V4bfnjJLuRUPgms0lZMTWyU5+Hd
URpW11vHdHPMKqBNVCLtPBo3VnrfBkekWwNPZd9zh4/khbse0r46ROS1czH8z/Mw
4f6QfE0fXx3qUZrU82aIR9a9LSPUj9P5GftI9Owa358IAngF1EFyyExh+PMh/jq1
HRnCzUIJxT7YjsNV5Zd/QYUJ8piSfAfbV30/dyaVJD6m+PYWREUt9N1nzkcFrhc4
XUCTozklyNnkwIqNe95VXHDyJPF0N1eZIFnekFUIheTCnkhtflT5xt7r/48Ay6mq
V0th+n0aUeyoyOrB5Os7fQKYIbiHiJtm3h0YgV4n/b87JPsXL8/Kz7dTo/qy5X5i
J1PeoNsSUYQHpQZidSWrzJRMlVe2xq2UJv7PzohzB/UTmThUPMhHOP+l8ZUvkXkw
TIGfxapXZchXscIxv7fKr9dMdY9hvtpKN6Vh+P7hNOi3udCG5KhYrHn1Xgd5bxw6
GwZGKFtlLDvkje9VxurZSrfFdQVMtQqGRBvskK4QaVlGOx16szr+GrijOVjyp4cn
STqYPqkVKXpU9HOYvgsotRuoNnkMAoHleWrFF5avkvnCjOFMpHzzMaiOWdUJJK2+
qSnTarTDuZ6w79gge8+HNMC/Lp17eAKPnQW6gyER+zKMlUpRqNYY91MOSrZMNgdC
s48bXOd0exci9lwhQPHsbeb9Ed9ndP0Y7zhgMR5gPs9n+265+lJ/hbK6T/W72xW4
Wu8Wm6zULCizA7LknnjtsxzMhlfOeyROMDZZaHj7KbvSEwfxQYBhBl1L+xKkpfLD
Qpwpez1UiKxpl7i4HJxsZmh1QFV2wmUnTItjIl71+nkZ1Jjsp2lF+k/nGcMlsz/o
izLiLaPmgHlgWHWYIMG25KZTdbj9iTeFQX7RqG4eurwsbyAD3HVqTaHqO73huikJ
YjW1wHK1LDqoqyYbAoxJJYkPGzgt4qiNN3vw/foDRMuoZmAb8jUe6vwmOudHWZ06
F55vjcmRqCRhNano9vi4uM2+9EyvSUThc7rWULazKEr3AmN8P0mr3w57SxrCPuLb
+JIULzmXO3H8+0knFL3LLnGXr8UznKrUdbDmI2SrRLJCmAycWfN52TEj5IAFXVcV
96KZLBamjU+rYOjxn29K9x8HVbDDAsbasQennAJr7uAtFl0XKaXTt32W3bfu2O3O
rdGnTccYcMaO1vk5hoPAUKYXwnKor+i4UVUzXGzVz18mLiCa+QA2latfLIv5RcB3
GNQOiHUSitWvPjhrcyTU46i6PYzc3ZubsiiMJLNdl6DoJtn6VypIMAnSZ3u7PUJA
UVVb6fj/5VSMfYKE0A/S/YMtSeOU+82WGBqww5wFARhRpPP1w0pO93BN8beHoRgb
kB0sPY/oaeJQesaNP+74uFm/d+kpH6LvcfiBsEgKOtZhzQ2PpCKpGpiElKECpjTg
PsBiZqRezL3TZ45wzk+RkT7BTyCM7NFVAXDAninlMhq5wxtCkX03SApAccu6TyQG
l8fYG5GNwlSjnl9iLMJMy+y8cleqnjxb2mvYP4YN0n+7lAT3xY4RC1YzJIo5ovNz
2NPbG2W3kMT/BDIiV87uBiB0D9TMez0erGPigrVJL62F2OrBusquJRt9GG42I10t
WZ8GpWaJBXXeo3VuUZ8RQQugdW7LjhEAsmVbAcYOVNa4kVO7X+ks9Z2e+IR7hnYp
qwHhjTmEW5+V8fHUTZ59JH/VKAUMkXVd42qrCti8H3l/EVUHBc49HoXAGBMj3TEs
bajLmGi8pO3/I6VxpkFNCF6HUWX33n6VMI27mbeXjoqZqcjHJseC5U4vOP3O1wdW
t+lolD8nyEf12WsRd87c6leLq/yYuYMZtOnPFt+sgBucQHpo6ebZFABPyxZfHyVc
aJH3LLOquMWF8xY1XMU0QaC29g0QAW1vyFJffRCjP/a4//v3ZpHHuu+NTFjegId4
18xNEmHu3wsPZonvPxikOuzMjSa5BpGv2mXOhVBfyR/xNj+3gX81MrM+0HF4Gjuk
Y4PJRTucHRT/O7GnhDRS7wjaYUFKklWkkBOVS0YkThVkAeSCKcSTG5IRuqtZsA8F
HNB2RGEq1hFEg8UyWeEBT62/ULEWuLh9ImaAamqDJUbTpvs0pk1n2YinyrUmo1c0
eE0EHgp8qPf2j04k2mK7HM16TFM4cekkJ8jpjVWFgfJEWmZM1IXThOBWsT2zHJhw
o0Mzejd88A4nM+ulfV1b6MEu8y0yVFeeC9jPzu+aodCEOUSU68ZG7y4ZE6B9xNkv
m83h6e6/lw3bZrYcocah4yeIutZM1/XxBDRUPacBCuiLnb7xy1hyPP3/Fc5AwUZK
jc1CqGesX5JzV9y1dTpNUqXPoovLiTYlDLKTETEG7LYzZBfCeVr4rSVSIhqQv5RJ
C/j0PK+r4hBmZZcnd99qVu3WME3VEItRUKRqoREinV/f1zzRgMaKFSeIIGOzighY
/mG9CaZR7L87Wpn5DurUQL53Gh02ccU+5LEtK1f5Jp621ghl6xAJKl/z1H5mqb0/
qibIi3s6SX5PNmqgpaAqRxpv1HKDLs6tpg1hE6mv2ptk3L/VH0k6/PTpjCzLJttk
L36Q35eKUg9VczpSwYIjxTp3TPVBbzsPMurhDou1TcpTDhf4kOOFMk0lY8eIax6w
tojNRydIrqnCZTHHF49h5An62jOMINBVdk0ioarBplV6a+WcD1rV/iZJrUhr0vYQ
La0+VhMv6M7hCj8t9owoF3TgsgfNbIFrRkdN3Ehw56lk9Gwf4uLc48j0OzkCp/Fm
Pbzfvfwnrey5Rq4RXmFAHKRsW8P8VZOx+YsojyZDyZEbc8j1nt1LTXMpCPqEkSFV
qPbprym8SQHM+QIQeJHfY/W3QAxpij1ubU4EE0vkNRD6w2kNvqngABpQSr3iNH/q
4Umj2VFD08iasvBWJ0nPh2nLfUulNpyHJcGLSBUPZYGc6BAIL+1NbgAzjAxAJGeY
ykbCliYXjYUoo8x2LhQknr1Dzl/xXv7OYAa0gTkyoenG5gB4EqfhS0f5a/CzVs1y
TB7fEEqlmR3iV5RhA0wsSbfDsOpdKZRRU8prpHomlonLD1esPvMcJkH3HLLnULBC
FchEYhWn+d/qNZFiFAhVclkm70Air3ScMBWHI83syhBAPH6BILr2XwXlj8udYg34
PniibTVTMwdcasoUGBKMv3EJZkDPTEPNhukklEI5TAFLr/FXTpRaYYCWkNrNW+Wz
A9kDIdRxWF5VE6tHSGnUBNSubcTIx1OvrNYYAmFmKmghrk3Np7jHZ/Df1bl8l7pL
G8VZwWu8V0j3Eh50WhzwiCR8AbwC2z0u1m92eqI0nI0vsqBbB9Y4jutjqLO9psEc
PKEPM7etGLTS5owmKzBANbh+GNObItAamWDfjxXiwUXVLwggozt3yh28tb+KjII3
vCd+608+5dSzQZDfc+lwSygizAEzTvID+U/CO9LCyX5N7ryRV8pGbVYF0deo0ONo
u8MneFblpkDHJH8UmjzIyHPVo6B0TtPcmKMDO9VLmGrhX2U+zgWkKsWynoDe2K/u
cLE3+5YYYt1dnaf58bXnNdp2kLQkh/iwbjYxChQuKTUcc1lghOh6F0xjMRgA+Gr4
2PKBg4C1W2S4TGZ5otXyAdagqm7/fm8BrXWGP+CLAtmA8yFiBehC0Ur+UbuxI0az
UuDzz2lBZlXRpbPAiVh1AshHGJJS9j1jdWg8st20Wj8w00WnnAH1ZJoN1xZDSVXD
8OwbRv/uNzzwiIciutCG34opcM9nrnuptiwJuCa9JZPYtcCYpwlSpQ1hxNXRq+ki
eoaHuP7aV5BbIXtzUqxiHNVQR5ec88b2+pnWHpNy7bm01qMCccISGMciqsou82De
1wMYpG0lLTMedsoggZGs6jMwIHwS2Bux462+QBN+Y+PWoRDadJMbEHyjkhKK/cad
Of2hQixtgougrd3ieggL7zRqynrYzj+mQUf+SrdkOkX7txsAuXbMnVpolMYEG6ah
0p39qdppCOxRN/UHlv4GP6MYX1xACDz1LXHVrrObTaaqml56O0tdjjy9Z90u62qI
/FJymWdYi0k96UIZbKTF646dFaFoHVacCTMn4jOL6SsWJJiV2vrRs5xkRTQmNd4l
7G6YuNlBGVp2OwI6Ea3JD9P1c7Ha7BnsdQDWsuimj4eQzH1AckKasbAyRy6cMu31
2gpDjkA6Bo+9jbq6dYfo0RxoQZb9GhbuNhfJT5FrKfa3UY9MO0Pfhk+9p/L6jXoO
QhmmTUj+KEXnOOVS1GuMH4UwUWRZ85KgJffabDmvvQvJVuArVA5G/zT7TaGDCKdr
oy3692WlCY7KYbuMVnoPr11vmvwGPq0GtnOmIUVH6ha4TttGnkPX2zNWIA3b6ChC
tzTSlYkfgtGGIKrotMwyiuFINAjasJbl4GfLmEncQHAYAphC8/k7xAmkrQaSLQUx
Y+hnL09CwiUN/Pr2cU8pJbcBVv/uyXkFtFLIMsmEKnHpzlq2/wEv0KYtUaPCZuQg
TYLaq0BRTstBKXU8hAje+9yGBARO293/u6XURD+b9FGWL8cIl/Le21JKMFW00BSd
FnBLVQFofatYam6FrdK4ynTSWWP8y7vjxlhJ6M/xwlU9Je06MX25cFjBSPtHsRY3
LYX4rFzeP8ppAEY2SQcua2gftbnOWLJ9GUkpEwM/aGohRncrO1Vh3yYt64G/VC25
bjQ7Bz5XV+hV9UITlUmqxM/zPxP2inJ0M7MVqKhiWLSAhV2rpLb7Xqb6sM+nIthe
kIkhPM45+wJ6oW5K6Y8L2q/4cp0teETE0YRKL9rzM219dSwxiLFRMWyXIEXSGOyO
cgjL34xs4I5gXiq9lncSrhwC199i2Xa7OG1rmMyGQ5H62P6gPqQ7PxZD8jGDpdE5
12Rd+rhE5FPxfOxSfjtmd+VDpZs3dm5c/kvsXvCKxmm5Gxg3GJ8QuZ1KrT6aVeB1
+L5Pfxnpb8FO7XtJIQ+rA7gJXN/8WkOcF+LuUQLF2dlgpPE1P4tLGn4bZk1gKYyu
v3qrT7zZl0k9qqm0T4PkdO2ahnXdPaY5UN2ZfOH8385NVFKXB7q2sxVM8dpHMOF6
yAoSQIpRJhZzxdDNQa0SB62M0WRZ5wgZmzai1EYXbwlNVapu7oq8v0ZfxapjPRor
dmdl8OVWXslYip9zA652dmkJIsJJid2esDsNCIZJBdzZbBA8+1gzhnaWoZ+njcaB
lnv8aOGdWgvIXzmACxpxKecwJ8XvPrBpccP45fPAc+0MEU7Fqg60LYLgizejHQiu
43V6lZUNr5EAqUug/ydb0B7qLfZbgkeIJ6shD8/n7kduGQS/nNLPN4YhPPGkcSF1
tnP45N4lQ0VRS2QhFNi9lEw7EuNy4z9TpBpKpDBB6QAO2d5FEPH7Ahr93ruEFyVq
111UOgBVWXwCr1IxDrEByBJJczA/yhQnv5zmFqQH0f6mWKv4ncWqoBgyxn1f+VDG
bMeXyS991jikSGZV4NmFdqR8gUrPZxKnfmATpEbQnufC+CF4UUxCxmRja0sQRKef
+L2NJYPR3uFb9voUcu0m/ArHompSyWhx3gyknAa+7V50rqrOljoxD8qUUi10+8Or
09+5lDF6H5iAK4xUlnWQWFZxCUx09owXL249EVKcdHB0Avy+wEDQwi7FZy2P3eL6
54FL6WXr3lu4DIXqnmM1tP9c0LLulb6fSvnsIH9eoH2gBK86NxNAW3i3KyD96SEb
QocCvmD1+23K+99Gl2A9r3eSzOD8F/4oqt7A5vqC9ESyfBVBL/IpnC55agom2Gen
s/bg44LET+2aycOkB/EAg1Tv0CiiZo7ig5Ri8IeGiyFH8qMROOZmwlNLTgEfq2Jz
rrM6xYXSPNmC92ujFquqWuFgSj4kvKFjQeeymbfJQzap1JnyiI33fDjkcdT0IsCB
27OfyscfGranTr1R0AIaMVqB2NdTQoD0cHEn7Q9aFzEE2TR+xsvHvVBghTTc93XE
5dvYiKz+tR9MLmkSCjiHi/QQye2n6bnsm/YIiA6bW3IoBDAMuq0MxEy6UaGuA6K1
+7ATN8Py1tNgaLy73v43s5BKRMo7NlJ+6k4qSQ1LEBXsV5WII2lAH8duquQuMu/e
zEIzWQ31mSMq0kJ1umHKtCknnzCVzV2h6L4pATEkautLh5TJrzwnGlsHOLgddMlv
OELb0UocbmwhTXmK6JYGAKVxVffGBqOLhcZgPPZkufEqA2s8Dsffc4SHgGpkhw8L
agua9b92V0nZ0EC4EgCLoAlneIv7Qu52M5fS+0JSJn5LjsbuqjmECZebHfMjVtxw
3ecYNH5DQguXS+hRLpU/RaCJDfNGMK1le2cyxajRT8F9OiuQfpfnN4L+ULWjtbrR
cEf4+nQpl1Bv1i41+XERPIm1FWyhHVVt5YYgVCtAJKcUBbdY8jTW/qbJ0fmszN5U
JtWU9P1/X0OsdfK2DpxB5M+E61WPswcs+oHGm/JACbXa2OT6VWw5ssJeSfvQk2O9
usOqpOr6YDCPovbv83+TgnJ/abPoFrnfaFvvtoDdz2/b4PDNZUX3s/OfAOIWtF0W
HzLsij8+/AuEz2zeGYjZj7Fy6bk3+m6HU3PKGpCk+8gNKY9rzL0b2RFtlxt/GLkk
AzvP4BxpCXsc0WeOhXRV0wg6qT/cXfk9uAnMFp1Rh1/PNLSvcgOHbBvXt0bfnvs3
z1UQ6Z+XjclWQGbNmclw/Jjo2sM+X6ZGzI5PuSnI6DG6DukMoHBYmU4AeMacKOnK
eejm5vBp3475eDwz1WT1GkY1TwNqqQsW7p7HFwzAX7Sbm7UCIgodcW4TOSSysaqB
HkL1iqaeUc/on/LweSCsjwz+FFb9Zfs+iyciBvy/+robCYMvXif+G5MhlDiIYHNh
acJF7Ut0Pence08amnWM3qVHQaMG6ZaWuRRNWv3oDZR3niFfyvBNTcID8Z7+q+55
gij9IHT95IdzIQdR7AmA6B4NVc2hWqjL4hhYHzohYNwQT4Y9a9IdDftXKh86W8PD
/ZvhAe/pDTZO/qYSyzSrefuZZ+e7QiYVwfGSS6+Gsg1vv2o+J8L3G7JcTb/j3FwG
wSAHpR9/ZGvZb0a5PqP4yGkG2vESeY2FGAYNZFlfZWjCOh1SXKsFD3xB/BzeCNi2
zDRglkD1uNxkopb06oWwVSYU1artv44uezDb7Jdh6gy9BJmlYv6lQpAfVmH7n8TL
KAz2jHmmBDt2dB+ecGnqKiIzb/weioQqsxOpBY6rOdBGh4kPkod0GlDd8CO37uyi
xkvFPIH1hiQ4WCxxt9oJUm6gP1FSxYD3ivLDC3NdUFqUUxI30if6u5uPCElsVJ+8
f//Jji95JebQuagKvblv5qdxvDBihd4Rxp02a170mgws10jcUYal3kxonHFKrOGR
+wyVag1sPpW9lD6dJjKC++RfJfVoOFt1yya3TdU65MoCfpDrbgiJatse/eQpmHmL
NTq0kIaVSURu9Q5iUocrVH0gsqC16JKm0cYnYModJrB0gA4sSekgsbBI+1a3IkAs
FCILGe5xVv62tS8kFxJh5eI9yhKmxy9Zd4Hf4Hk/BqgeCsrF5ILhaYIf/J23lSWU
ZYKYzK2zkb1qDZXxNhZfHv1yMKKsNGh4InMMlTNHb/6GYwbzh2GeHAnvnD9lGiYK
wJmQvm8UYAZJoVn7wSik+SnaxyluLuuxEKF7QUcnca0VSIX5CP0pmfwYlkk2MmJH
17jVUC9j3MlVp73G5XuzJfRZ2SCcIl5jOIUSfnmrKBWM1jEhdig2vRXVXCuJx6sb
pI3hGAiKVWwPV4KTSe7ttcj4CsxSqA2fT7RFaLPGbpARUOuqyd/lE0zJLWHtNMVp
a1vp8Qu+c22HWLFoGXfFCQ1DtAg6EGq+wR1+m80pXzQp6r5BrDIgtuufn8uW4dU+
PPIgVRWtfd6joEH/KuQf8oAbzXuCt2s24Xj+71qLliWifVfsut7L/wrjokigoRJ0
v+m+YqjRJxmKL+7g9RYZCqsXJeOsduE9+9j/3vqW8Rb4i0Gj/de9SymEVSv5TjQn
t7caLYIPfG15EqLFDqNp0NGGmJtulev43edgmlU5ix2ohZ+tpV5hIgDoyPCBk9Wg
SNZNyQ5LEOcpaTkGBZ/L21lIDR+Z4Yl0Dgtxk/NWzn+6wkJhRVLccrYoIDmj4eOz
LvPcWNBlkfG3w6RqorzLwdiC3Na9qoNlfthB0gNmr2LRAYNNW8biYJk0GrfItU8S
kGDV+8+bEfghPtwCnVnE/cxt/bAFtk240zOCFupvXM37wlambTSjs6MVqd4I43IL
QF/SnfV6GE0Lq1yu2fBNZM8Z+pxrE1f1Q9n/ajR4ez/r6pHYgrw8b/7XEZ/ccXkn
iWQVmmZ3AvWBx7pl7cmyKv/fFg1oxtFXtzFT+N/0VUeCI0GhzAYx85C0abpmQQB6
Ft9/FyPskum1ULqUOPeQjFEii7qfo2E37D4kPDKRdGGLM2aXoJLbn3O3+bhGh6X5
Z9oYCRThffr3wSHgZzMjsNE9MxssJgI2SsMFLcLCZNiX0ZR4sc1Y8f5oIzbXiYds
gnaY0LvayIryuk76MkpUqACI5VJwEWdjf+/gW+s5frJMmr3kcjwAm7CL8vlzQNhj
JZSrnH9avxCajFYFTp8i2f1TNp9M6On7wVnUmciezQA+RMJzl+tp1DhMwcrbcohO
v4i0hsVwhaK8JQxjEGJ/zbDDMYO+kZ0CPI3mGB5FaU1ZeA+VtUgoawUQs3uHee5h
iC/C5gfr+oa8Xg5dbmUVciO72VzpjmDTseNCPBORCd8hkETJiM4TtJbYoq+kJuvz
o/UD0LvKbOlDLFiEOaKDkS7CMVjAYLEneG9xV08fKx6D/Ytb3iF8rtDtQoTTMalQ
CnubEle2EbCUgL69kQM0v1iUa+4jRtLNreyVYUq2UPTVLBkGlLo00fhfnCRvfgkm
r41+dw0NFNYoi/ygagfsBn/JDuFJPNQH720fIc6PX9izSlRpVfyZTzXOY06OzCkx
nlb75dLYvSz1YzEoQEbmdLJ18662uiyp0AsBky/h2DJrpc9v79R7HUh4QCJ+UPHK
dtCxdnf0Ok/I7m7DRaFtBexGS13emaI5DRqEy5Eeda8Q4YW10qcVQytch39edenx
blXFt2eR/9odYFKN8MoxOeWSVtkAD80/854aDch3vJqTFAjek6KKkUCrO0MzMEH7
/92DOzXZlXXKDvdUn6Q+5GRkpfkgttV2AMY4X5Aeh3cVEbPXg110kLShcCpi2hxa
TL53+LKhGgWoNA4JMydKDO9H7tV7dIfvUXI507AWwoNEP96Jjhj5PEQFr250rH3g
LvyRQ2l6voITHRC3gJ5I+ZXU70JAGpnY5BNpTah8ZZghedHpZ4m25eIv1e3C8DE6
5/0Gm/VAS8UEyioKUNmMYvfLssjNRLadLDgoqArE825IqJW/NhOyfjQgatY4WzWf
QxWw2qQb2K1if7XaGyhhLp0RU6ZxXkQEpRLrk5tAQ7+oixqtV7598NTfcjsvqWKv
XMT/16Hk2SDsI0Nq0MuVfTg+1R8Ckf/m7VDkJSwnobto7n/Yvm/zjH4duRjSOrBy
NXtdlyhm1GrH/9NBxXQLgEkjgkH0ZrvNCi9ekClm4KanbljJD05TRGIpf4YWhfkZ
cTMiXfOSu4xvHjG01KYQBZblZ3G2whjWD9oOBs2Hewjue+45dO4/qydLnqQgLAJk
1ip/gZDnT2fJ8slTemFFr8FLTAoXODdM4wJwzFQt+bkUvT/4rg4yCRCjsAJ+bRRF
n+pkwqmtwBODhZihqFjCfDH8NqawXbavRDVFwQcy4L1ukChRbrHwVWQce7mwfioX
0lSq+BnvSK9WsllKBlHigeZtOc2oe5HLv8pTe/p149hrlvWA0PzuVfHj4TJdu9ZE
H+H4YyCRZK00/9S0EPWm8Z9EkCsCmtcSunstCdjt20eY5JVDlNcEwLDBMiurxh1f
t/uFajnQGJqHkS+9RsqB5KObBbypVx8nHt5B9Fh2Pdehm4ShJqpwXREGtRBatVx1
RxHqM704n+xu5DGw/O5ttFq1De3sE2m/4Ok2w9fINWTZ9rgBgqOxc6KgCWQPB83k
WjSNYq2RFMPr4ZDE5rXpdCHfnYLlR0BNIMFt8vl6OnnX/mqCmS+9eq2YqEar7mDF
Y3tfwh/x/t0phISvK73YoYxz+ih7W8YjGXu3Y3r9qDVbz6CUcJaUSbO5JNXzeSTz
jK21VyxZvuzDM+v+mA3oh6Tk8iAONga+zqxNrChOqoxgZpRf5USmFGoK9AxBiNpJ
RZL7nV3Vm+KEb5GYjiKzPiUGLULHqZz53M1x7wySLE16hWZVmZWrvKlJoXgQ1m5q
UF5gwDd1g0vx4iKwBVLNjMWGyrd7uCPsnAY75DxxRzqBqYgNW0h32UXx58/0euGS
88sUGTsURaR9We8V9g065ZZ9wZyFZPbVutecsE+6ynVR4Y8bBHKARVFZgSJr/Vqy
iIx7s3tj70lmsdqf1UZGCQvMoOE+IImkgwU8dG/rs8NL0ym9rskPr/3WMNXU2jan
K81ZShrTcglGR81xvuT2jFb8qQ+c67v3X/yLy4Q3iypoYuJPO6oPWf6HR7BiArln
tUshF1jyLsgxydh4YUlNnrIeH+z75OBpLQjgIKu6mvs3gmsfBCt3q/6pe789Mga/
yXLBfMG+0Q4mEzEPwfFt47nalys5hh8bb2Y8W4jdp9C5VQODN1u5lAO/wVGaY73K
XLCp+b5tyS/EujECjuAB9cOKjDxhHiLyEdfoPJX3MuiGE7nIHDUEsUDIfAILnWhc
7dZMEz5BnodgnjTQocR/FG6lw0qP2jT6iLoOY+HuVPHzi4SJvfuY9ObT/802a5Fx
qDg32SlqzwPhDwku03bwNedgho3ah8b1epVF488Vxx1hAhid74d07Bz1OkCH6IW/
Dg45Nh6nv8YQzy+J/KPFMLUv/HMUZNiB+EHnkZkephAeISez9FdeYP1Lu+JG3PqT
GKJTdbNJ3rgcR0RaNogmriFVftcalHVyL0gzG1Rm/XFHpNzLPvUV1KRh2Y32lQOL
9k/IOH0GSxb8Kgrj2ZyMJqVOZRkUmfty2RAav1koa6KphlEDTbNWs7upXN2E+Brg
mzcxA+JXQ1JBHQft3SQQ3sJ3t5noP8DEYdVzIODVcxb0iiQu2zYfKg72kJwGPJA/
17FT+pFOQJEYlHj4vanYqbY4QKOAhO/04IpZBJCGPtzb/GIHQ7HtT+P0BmbWEKuj
XLEnRoUlyoGjvT65cK3snPlNq6HzR+gP/rGh3tVkEy5ROJ87RiwVqQ/x2H/h/K5N
+DbVKb3LNxeF4ltgPkDh3+384AndXWIvz/faMAdE8VZeYmSvGN4QZWEhL84s8Gfb
K5Rh0Nc5J/q+ZESwUvqykvBe2GYTDhSLfmkkxfRPEs0RDCgioZFNnqszpJ4DKzo8
s0OpHa7JWLdD/TEDsHoa7jzEAtRA22Z7sjCq3zDan5IfMafA+O2czZHJwHpW6Al4
+pFlXu/MwZ+ylLliI9qTtowwVYvVuYYd3r/hr7mOobZ7oZe0pCScvGyU4i3j2qIQ
5cYpuYVU5JnX6XVWCSvAtsAIq4lXPlo7h9aRhriQ/0T8uEC+4uEauZkMFhNzluw+
La8wN6iPFJOCJw3xuXXeR7DfPdWzeUhB7H7yZ8vgzgInwhGmxKR136epk1kSU0PP
t6RZQIRekmJ2HkzA+9QkDsTtMDDgLq8LggpWzEVXMnYMCNT5YS32P3/c6wB5QHbq
8i6dkaAAtADK9rHhiXjUFX93T5Xu3BH+yX9yEryKWW5TK4EzNcw89Ms1tDIAwi8d
zXI9hXp9ycwU3ZMEfqRmTkNDvl4Lvvw2+uE4g20pyoBD519yKpAGjDiyAGm629t0
L6kcrDTIcJ8UQATxdFClphfgWvGb+rTbKgW/r2DOMM6axKtaJ58krexRzazBHzk8
R5K5B/5k0UgEjSFLsTdE7kbnfQ3eYJ2Wi/s6kL6bSDfWjYxDLXBLLGElsX9DKS/8
T0a3JjyLvV/9pCG4snwslnsAtrr7tiDtcbcuUVjCivxbhI4TBeYRxMEUFToRIAgL
M5lJGOUz1OGhZV7Nm++7Q/Ce/ZyuRhdpfmPBbdQWT4CBiBp9IL0EAvOvrJZs77pI
i+9eP0Wmk9063BJkt84ht4QSKretRrLFHu7p2KwPW0wH6+qSTnazWopxlYapgMXH
p+t0BvIPEwNhzBIEaIiyxNXfRlJ5apKRRbrOrm/Rpmfvyq3YxQ3AHMJXybL6O83Y
Ny0MMOYECW+kIz+BqGIqzuSumyfFqXdy6+o2K0DzFmbvMVZtVkc13zayb6fxmQeo
YRcvHV2t7oNtmlf12c4KDppTs28E8WCCQbdG1GM0JZvnpHsu0R7ziNCgwDReg51T
iucgDUDneuWPUhQLrD9wWirgU1z+52Xq8ROuHvLcRjG0pv3PMHZ6B4+azcU8bemv
wa72h6lSI1GaJx+MHCJppnT9pW13DX+rd/Ov0TvO5lNGiumFjHV70q/fry4sii65
fwMugiB+3brlIHz0LTYwZ8zppQs2PLTN1bnt6aKpYwvgeZDemTW4FhZibl8Y9iyz
iXTCss/scK+pZQ8OhjQbCU8syuVqDYjoaNn26iGDZpotOOR780cBPdGe3o35cBDH
Fb9LMoFG24DBoX5gKI2KwQKT2V2m/7M5RQD9IaKlCuw45DVz6gQj3f+oeZYptRN6
DYLIpuFpGwXsLaXAGdxr5QX+LGSD7ibkE5ST5xCNlFzSewwoyzlj0BIYvLGcHcsi
f/x74lxJlBG2BKJN2p0SAASBarmYBkGSS4mbDx4xycBUSVR8VxVo1gwR2jKK+lil
2Bg4avmIFuZ1xMGsK/h91GpKe52iyVVn4LEMoweFULYuL2z1DXPpHpbhZtxnvt7V
iVBNktlHRvYOdtaKDWlfSSL4lgjkESGMq25bhhnpEGjZr6GFsiTRrqdUHUKEvLH7
6tKZZHm11D2rYtQf7snZUIWRxBygLeuxf6GQl7Rdp1KUsf9B9RJTDH/jOuVkFlLJ
C0gRhRi/3fB+UQY7dJBCdm/9yeicKE0d1Qsc63nLGE+ZfuW6VfCknesX69DxId/B
6ICUTKNyiODkOKsJIvQfI1PYmgQtBDYvPkS0gCy2E367fYm3fmwb9WYWGq7IhS11
pyMIQbUA24Lrty5kPduuTRxqJgWAM39LkF5z3sQ+kwZbyRYLX5IV2Rnp547Vzelf
D29xrG06OjEzA3D2guXr9YEHwHyUD4Lgpn2PTmydTQapeoLPXzxiw7CcfqbuvxgR
HFFuT8SD0yRW4TGJSimSZK84dbiPNKItbWSXIujRok/3bKm2aezryN88+tlpLkFh
wOA7zWKqjzLVS+40LohmE7w0q19NZXK5gy/qHiul/bZhRlmuvpKdVCM8/XvkH/Pb
TE2d7a8pHtDnbEaMhHj21gPRt97kGYh2WkOuDsX6Fs/jm4E7oy+mCr+IzANaxY4W
gCAh2XrjqpN02s1T2OYJXAI3alcTub3W/W/50ClHU2pCOis2lrop29lbHgid15Y0
OYaQNPRbCyHgF1Dr27N3LNUn1mxcQ4VW2NcSP3Od743D3nrZrhQuDCj0vede1Mm3
4ItTLSzhnQ2FfCb2aF35zk//dAd9jXRukWRp77+jX3WZc2lhtFXj5UFsGXps7SGb
PrugH8awJDBYWxEqfRqD5+US9n3OVuYeiOhK9caxrpLEJjiRaVsHQU6256FiGDip
TPWgr2+JK2YqVmDP21dl0NRB7tIDTOPPLe6ALHwWduneem7goKbbdm0Llkbaq5Oj
rr0HC8NfDgd8FiCqz0GVETGebAhc4YYkbQMv190I28IySgX6zrR8rklKRSq17i7G
N3399wh7tj++rPasD8tLxMz9km7iHa6ePziu1DhGUZiuTlm9rvjG8g0JBmEkKr8y
kS0q0OlHLMfI/c+httOYAH0dlFZKCfT2ysOaYmBfHg6Vs0C+Z7WagNRwgwrjOvWu
x9fjGmPBRvMPojBDQggn6ZRTN0J2jhahy24j6GYTwwEalth/bfKFD928Zr4+WgAF
0ZyK9/Fv1GUEhE79gszyByS0OY+KWMfhUEG+hT5TS/qa9laiILbrzynVrtRWLqB3
81A5RldKRYfdjWjZhJ6vSCyslRFWn1geCZ/WSXV/zb22Ko7lH2RJvoBm0WTaL0zl
TuyWFVFWSOXxjFjjQDQt4qLR380UMQa1ecSXWjvsk9GfefdX0bNjB0+zLmYqvSic
00DXzYwN2Bw4aCk6yEwzlCqcBDWrwJ2jLOvSkEcjoKpCtjxr58XL82OZgjY5CCsw
aZqpPFYxCypf3BuQOpUSkLjL9Fvc1Dx38e6+r/9kbM7XFEiS9mlwtQAYz+BXmt4E
ELWS4OBbYEANSPW33G9SqOAh6UMChgG5t0vaixKxfrzQ60z3g57jS8s+/bd5q7jC
EGP3IKmLMUvU7KPRhq9wTPTouIqOv+iCjc/tqpVwouTyKZDf8ztJpt8EgAyvUBvk
0i0WHOfhfmsM9CXLdlzqhAEPcFoeQin5Z9rGGmmnDQvbFHgEgoPAe/N9Wqh1/iD3
ayygn+5j/AtCj7+3/LbX/kfMhuO7Q6DhGO0YBiGVpycJKuvDxTm3GNDcVVddEDcd
wiI5dphAoib/A+GiXTvCqRab2IcirfaAvn671Rl5oVJIP/WwcvsDrif3KhPfvF26
wH5CE64eZz7cAOn8YlHAl0TxuEdFykYYsdCY7VIrT8yhnLbrPDOHBp661NVOVpTf
BxiKHNzeww/T8DutKSNufulXICmuBJ+DYiYIu06d+0DGw3wVWzKJHz8YpA87eUxE
nKPu06OLNkeu6k2OfsNw5bu3v46IZ7rd/+mqQ/vZMGvjwDWSOH43/oPqiAANUbBT
8t7MA249ehEe60NqmBSAM1UC+RBZA0FPPuBzjNNPtt2zxRxzEWDnPgjTjz3/vS7S
3DIFZfHbIxAj2JS0q1112HHnQeKueB+9F/xs5or/RqHwB7wLJIbwo8pmyqiNwUX6
5NKF3loiHpV/srtnthV14jTM+RGNhR8oqzh0ng3GLBVijm/Vu2PTZHVWCb78/pVx
/30mH9KvMDs9++ynXxsGh3bXr8JwvkijTP3gfVbGc2xAAv9WGW3FMEdvO0sv7NLO
4rPCtvHkAEQAUMfuiA+hpqv6ElsKPS/hz3mQVohIwMS9XZCxz/JMEm4//Uo27JYe
2hdL5bbtckvIDdj/IJvgd0YNYGV8xhu+B4/MjR2sTxUzWHtaWG3ZsGqADbl2EHhs
ovl4nj60RsJNsWMuUAsf4i/8Sr4Ne/T5sF7adh2yoJ5WCsAUu3IJRD3jYRpRutrH
GZ9LDeRTgjM0WPnkUt3bwaRz0X+ExkxwUTrRS1MFuhUAyWa3ojkZWMGa2EiixuYJ
wOV0qDZ8P8lclwU/zDd2QFheFpvZjwkrhHNBVRNBjzAf3q4Ju14RRokg//fYVzfW
ZR8mDS0eCSGGrXXcWtIKtR9ufUfeqEzN+tzilnaGN2oOW8BKnhsgqOPQ1Fzk3qDf
ntt/E3GkwKwSUS2KvPJPiik81rHH99jcY4kSZ0TYtKeiju5jYY5fzbh0lJELP6KU
szwsxwDDyoRj+EzCqckTCz2oh21hco6dAY29OReFsV/UTtblVoxI7CQKs7HIjDov
PPEfSUwrIOGj+zzHXM913JEV7aIrQauQsu3K8B9CE1nfzUOXLMaxuWaqR9zm3FVg
3KwNKAGrRx2XQo4qkLgkIbz8BlbNfBuSAilJ0sf87F7IRJcuK5uC06+D7kztcheS
tXo/cwBP38HoddCdY82wbbWvK0Lj58Ndoz5bEeseuasQsonBIjG1f2kFZlXpSNf3
uIhRObjGYRrKsqcWR6bC6vT62Bx2pDL/UVH0j3egRIZ3MbCgfEA4AssvSablPrHo
0pYLj79tVQpmbAXkWFFHKoqArNqZphMpl/b5itSBKSmSH51bzti1JOl55R99PMfo
XOsr14I1FujzfeHAfE9UEK1yy75UygyfDVTaR6QfZU8HSx9+LTxB4BnZDbMYCVbR
mTSWnLonkPgISbGAxTNC8lm7keVHajiWBR+CwDTyXFb+fb0MQ2T+veI20oKE0so7
dgmpxeDrR1imdxax6N9WLxZVaEmqbdGlpJik4chwaz0Ne+18d+BZxLtNN5IWEatj
D4PpNEY5rjp5nE7aq/o5nYO2FxxNI6wk/t4mIReMSHCnTs+W8kDLKB+BDg2qrADp
d3vxQJLrebvHOlEqn37vHMGRMXLwtYZmevytVOChW9hHF/aoNh7Xf1U0C5Gz4ZpQ
1y/8cKWJU+uIoMTFIcLiTHqsCTKlstzIaVS0ec3o0DvBHegnhT2ohy4BnHTxMn1H
pr8lKCpH9d8SznkudD96vGwVbNeuGT+QFXTxyOHBJWCPvVBUjRA4PIpqYCahmXTQ
QZn3SFM5H/wIbRcAihRx8rZhoAtWsCms3B1NjbgWJU5I75dqPq4wwjGWXhiVKSd+
+mCL/sS8pv1WhGcBsvboSor8LVHOKyGDwyG+X4/Nk+3AHWFOoZxgF2l3PFmgGteI
dTHnQ60AOaJnXE/7pjyJuyHVGg8bQVo/N9LQ7nA7hh8hCk5bqH6gYtYu/HYdxC4U
sZqmxNyiapu81XJZ8KFMdzproPnxhCk9Tsx1dfGxW1TSENFYNQgoY3nyVaGd1B4r
O0ZgiWpn4GyM3U5QVQiFo1s1X+Zb1F+bpW8kTjfL5rHVG8dPiuXFv+QPmScF2BnT
oZ0MApoQSFNGlYUhfhmp2APbyuxUevULcp5D2Wq0t7+RUAnu8DIGzDFbMS1nBK43
0Hx3kZNtPn6XYBirPG0tJhgUch2z0t+hT0ywNBpya6zihyiwT1I/tCsSHcMFLygE
iQgiatfIc+7EVzXusRsPJYgWn2EHPDLoCsbjSWviIhDv1o3shIgdxMLP3VAwdty8
xU//V50OvtdovW/vlygqmlxGunSMDhiAFi4Xwl+hqhgMXgWr8Yq95kThGCDH1scY
X++vtqaP9EBNvhQ9nfGCxt7KTgT4973h+MFmpbQ6Y62k0dxxE1LZztqlQqX0I+st
nbYvnF+S+toFkvLN3nIT9Bxhsx7AqtnY78tKKZgVX/0T2/wBhzXNJW/gKHkjVdXa
JGWNCGCfXIUm00uT21b0v1u2iWvZZV2L6PAR7M26ZP/WxJLYMoKPCYmzc+a6LDU1
odzQeAEWW41WBwpD8ojBA3yo8ChqLixre+Ts0ZtRC7zv4XGJituqqojGRcMjLZPg
ymNTz8X2vVeEl6ZCte0Up2CE8uADsIM2YXrPIxdwJsTY9WYFBRg2Xat3N1Bx7z0Q
FhJv9kuP68VaVGxThizGFlFUOm6na6c4+3EslN0YvgVphiGqMg36oYnpHnkCVxlo
tfFhTda6ybVWSCcStuuq9JBRZS34IF3DM5g49JqUhJXuIhN8bXd65b1GGxFO/IUE
oYMdfzXqTmnoiOFx71Z6Huy7BNCR9aeEPbRRSp+s58Apq2qMPO9zPPrFoMAQ0msC
sb3+VRtuFFqNPG3cksPBbWc8+W+QNZ3lVkOlfuRKb+s/nppIUO4TIhvmBkJcachn
wj+uWfP3sRM4mHVbWwRzzdFhWtPsVlRzT02KenRQdcAtTOkBFErvtt/3DyLeCIH6
RU9lysP5dHfBQNb7PpHGDjQcvV80RsenjQnxf0widnuJhN5pw/fChCNGEUuiIAtx
ECg+txpw0zKAxi0jTZYh5JV5PWRwVYvjBI8q8euof6ee5ntpHjDKCRu6i1+vNi1v
2siUpC7wkA4ImbABb/JlOAgiz4Hw0k24q4lehkJZWiGv3q53V8rCEkDjhiZEuSHl
iFTvaILUCdlNwQ895NbHO5lVe6//b/E6l8pL6XldQ6gsJ39HhrX8lxMYro5iO7MA
SCJcEpFa14mQcIdU5cGvLEJK6Aooj4iqJ9C1qabCMqc7AvWdKl9ft5xXvr3pitef
k61AjSbF85XykhlNl1PLKqBmbGruoesp20sUI+JIYqzYsrl0E7MeLjEUKZo8ONC2
46lseWoglwmMaScifHkLSrtWOY/4UPiMfVPQplF490bTnzL+HzhvvFCE27+KILxO
W6uYIOxbPIMJk7ZYgw3sHaEInYVRhEMdYNVEGBqqAV7pgRQ9c2mBFb7WqpBDTob9
aZ2UtshYVAcavioVmf439iaQdbzKjI15+Uvq/9yL3U4kwEuLrd5PSt7g34MXeg1q
FvAUh7w6s3oXRRri9Ueu0EitClg2tbW5FWYXmKT0dh4uewavlPRmRJ7VmKEVj523
7f0HkBf15gL+eI3PDCZXEECFrXvfPc8bv1ZP7sUjfLhVioTIT5R/3w2n/2Y/pXLL
RYEcO/4bAFm0nD519cuZi02UEBGH93RXuY3+n5WNzsc6Qt6dYRB8fye4SUdHxBPb
G6MijkOKwlTTOxGv2i7CEAgK8Bo4mXoAEtwCwMAVx/H8+nvlakpAzGi5kcWGCV6c
BZi+0OjpOsDnYFewLAXYz0dIx4Ak/5NXu9DAzk2Wp62RZL1rMxH6Bw1/wDe1gQ9q
Twazzi0Md3BQG1rb3/37JTqnT5DeHHmd171ugfU3I0G18a+9NK3tEZXdWeTMKt5T
CBWXjcseuR6jQxw0xgRRwssJv9h7vK/mZwTaFuUx+4jEcuYtgIqVJYP4UcBsBDbG
y+jS3cCRo9rJGQxr4Wg5bLACnaNChK73F7ZSjpILUE8iHVPfr7S7XdxJB/eYfHrN
JqTUAA/0t63PnE/vpExAHC9KnjzaqILmeNBfI3LYNO01ugFM0axrH6vDozQLFdo1
spGZ+NrO/rwbTFuWHMspTNwybdmJR5Uhl/gIsfv3KwOL519FfUtYsSgQqmAxLiKn
5UmGj1MvTZn6y1F1CsMvQdbsXMHCSfkxaKS3G4/HBNjUW6cyHr7mOz4VU8T+vwjQ
XMFOn64f485yZA/Ykg5gmQf9HtgoncSfaU+a1S3GKySkdjsstppBLCtAHDThNGBs
czGBCbVsm1AGsA+/OUpGWT11Qr9SuAKQffeGMs0no6m0X7Vz81JhnOnsZn6sPfzu
TdX4cCBwA7OgfdvJcribeZUM/3GNT6vOmNMcnoUA7fnKQZgIhcQlmiJeImeznmV/
TbOWKX9PGxT9lZLoN7vsBkH1UZXT24lcKCkOvbI4LG+LUk4cU0jZOB68GAIrtARP
AsVJYHDtARVTBvlYJi7G+wxPsZbaeUJZqjAv0CqpOQ3UIVD60OeTUeW1aQoCMRDQ
lXiVx2hm7sKLGVo5BxcwnVROEDLIwXXgJmn1I2q6bDVVZf4G+IyQB3OvPl4f95Ri
V+sJMoePDAT7yHatUyx3fKP9UuArxNtWo6LhcMaaxSuDvjT4EwmI/l8XFCuBo9p0
3wpqDEtJFBSTj9yxTGk60NrVo911zJL4J9rZLCLE4Nu9rg2c7lSHrtLGg/AHZ6n+
QjQo5rzFI9uMn2NP/P7aml9kRAklt0zw10OnexC3F/XyCPyQ7aWN2Ec0bU6qwvQL
LK1ORGnkk493ioXmy3HAPR1TKdA/oCP1ZNX5Bm4qQhY+7UOJ723aPJo/wyTMe452
qJL35X6eS1YpJw76gBDxbEu05lnaBCARyy8G+apvHXJtOtTad9hLmkk2l9OgF7Sh
hJa5bRRVbOSJwUkgawIOU5E92nOdtXSvNgeFhTRq4W3CZ09G2Pcid8xUp/3OqBCW
UeDeNnTVhQwQLNo6b/d0kOATG/qglemA9RvOhQH7hm6McMFkwewzyzVmtMFZjys/
XLEQPt4cBcm0sO043ujtHWLI+QKbpjLyMUvTvxKpqjOVOHXqbzEQX0rHCSxe/6g5
b9SqC+g+Tu0b8F02EBJsPrMN3IeSRkSwYM7uXyi2UH0knc/vjBcr60Jba7f93rQC
Yo3VaEJnt589xJsOEVc2svjPEibPvLMHqyQhQbB/deCqDCa8HTZ1Wad83A5EQ1f7
gajYXPnO9Iaf5nr49uGkp35j+R3Qo7vriypT8YOfFnGWTMOx6F967NeBxpmeoJHT
EDCO4sd/gzBxc4vyH3XbOF7k2tMZvRwE2TRQ7/QAu2cFvj9AD9S+SAKmrhi7k8TM
9IpXJXB2vVF+jEuNIgnAUIRDWfuNbzYr7eavSt92Ngty5qwVaU0rtoAV35WgJ+Iq
83FhPyh7D7LjBTPxBkGnGxl8/cq1q44CYlsHF7C9/fpCJ+jBnSVo9ea7ziyjcFzO
gMQU528aOYO9TepQAOy33fYFzYtBLp7DA3ABZ22YVmsfKCj1DU/XyEIgvJUfBjub
8YDO19UXEQoZyzPmCooIA3qgnkva+9wnxf8952GCIrKIk55EIz8nGC2Xwa5qUx4S
Tn/DZfGuYP6cmOxEM2MoXnEHo2EZOh5oEWUAGOxmNU9aQoI/VC7jNGyDCpzThWzr
Ztw8ojPiFyw/HdURdEsSJVt9YUOf3D1umEp7GsS1wEuyCD0ZNophSvG6z5RfHni/
Qo4+A+rWPLnzfsAfdS7vyYnCkQJ1alYp0h/9vaIM9GjtO1lHNw6hqn2UpSdnhxjR
g7EtLM4KpIaI3gcrH8gK68tmscBCkzq+Xa6silrWmZ0cDu5/yZbo76kB2r34b9Ih
LbIFYQVtDf5QBw+tHsNV9r1UXUIGCQhwHqL8dcFxKBpaJxdOMjUUaEdXYnzPMZjf
P7xozcq1TVMELaBmcnSCiRKFMu0y9SgG+bTcaIMaiwVgJuXrtPozAOsx01FQa5hY
qW+LKXcBEU3XQDxLW7Yu1P0+y/H+l68YQE9i55GVvCi5iSHudlM9l/X/g8OuQLTC
MbM6cXzoQI2W0NwkCiyza/9zLvUEQQMNOFnSLlD0R7aFZ64KGpVnj1xiLKbsZ0It
gulUvDX8b9f5z7HY+XzEn2VzqQsyDBtIiUDR6jjDVNba3sQqAz7hByTfX8+0llVU
lJFVl1Xh0eQihgOJpK3ORjWUitgeo/3f6iKhh7x/VAUP5HSby2u14rBsj21JG3pH
OVkpTYMp4K9NHrdKPnUfNJ3oBq6MvGUHQKpjLwxANEhH1M0a++Qzqtu1Ca99JOeI
1H09sX+dlLzcvr9XwXps8ufA00BJtLh59zXeKIkISVO7qOzBe0YdE2QDAXAzOujb
6pYTxEpFk3mjQ6CS9tAlNn81LjAG/o30kGDEWqvwGROqzOnipa+R+US1+4NNf8lm
QBTw0QAIYGxLl8OxQwnur5vGZgfSfFIk7YMXK22c4lnRJX/m894pY0ZricnLzI5G
xGtRt48ZjL2fFX1v6/Dvnj6iZAGPFqU80kWaoMFDXVpn14OcjVWyeA462VQXBOSt
+cU/sAnDXyyBXK7nj9+PwD8kHhNUitrF+GvembB9cxqD64DdcSJ1OIOIA52tXIEK
kU8n9RPdHJGodpkA2TqgkT0Ukrzhd2MQIPsezvGXBqdt1hW30pbl8bgiOPgdbYvP
FqAWLI99LAKv4HB/wxpvwKOpwpDu4/e0pc4vsjxDwqVqtBg/j+MUDkIsdIGSO+op
ZnII+tea+C2Gukg4H1YMNyfoUhE3vNVhkGvFiXUhXtsQmwhEUuDoIDli4wmW17zw
4WXKHmknV3j45fGb6p4AqG3dLini+sFzVtqIDdTI6k/Awk4doBBnaLAVofBw/Oa6
aTtP1ci3l4YQYhsOTaD2JM9CaHzwOSQwBR+e6eCO+Hfnc9+DyuVQ1ewG+STua4wM
9YYh4Qj6DWT02ls+X7gRx0QMTTG9ZfoIWSx6gh8iha84SKHGVXCpWJYcGqY5FuvL
kEBErx46KjNij2OgteiYw5GmtYZpVcxx7GK87/Hy4tj3ATBB7lefiXUBNlDkaOTK
ppCmoPNmqEEHvxPxS+9BjUXqBWewLSBUqGbv4JKcnIj7+WC4ty4pxlrqzXdRrTRk
Ncj9Q0+DBEB9DXTtMGFbXxniJKSHS/lSWW6V+npJ2yymCpgDD9uc1IXXh4DG8uXr
m+uBBakPIvJx6d2IMqfdb6rKSZYm8dLgBPDxi2mpUVUVJYfSUy+QMbs0kEM4yGRZ
yb2EP+6bAFUqTIL2K3AgV0lb7lYoxSDuC/kCU2ntDHPOY/qpHisBWknk2l4+koS5
IZSPlJFXoe1XHLJYbk7Mzm0GCP/dnFcurHiPpFXB+CV5NITRR2rR0we3O5M16++p
km3GfSzoSLRivhbjQg6pRBsPsQHhyANtVlmy1PI8ELPf9V/KxqLdX8uQ9jfRiH/a
ftPOkHwC9VM92G91/vTBaZQSfBetoT7OMmww5SFprX5QPkfnNQgHrFi92Bd2qkHb
047UPcjKKr/T43FuGBHiW8pcfffFSpWleUFSj9eV968jS6Pcx5AzjgY0mOErTiPq
ZAy/blg/AZqldnTPwS8VVQfAn62uhZw4zVXQ8g/ZYa3sJkGY/T61KohEfLOogYVq
EDvFJOhP04H5eXQFn6RhxwO40JtIupKccH+elQTICWe0ViGrqwdA8oyfd2DcgGb4
4a98UG1KdXglNCWkFaut+rLmbCjVKPPaf7KJbyv0QbWwHqaLp1ydZxLLTW20JWU5
OGn12XTbWSSuj1JFks34msPRq8JuvjlXq/kriQh4gOMN+y8pE160g5zLD38AtkqS
q52H3ZgKKnTDzZsgP3M4fIGvpGH0yvu1ApqttnIfWbMwrR0ssFmaXMhWc3T4ZXxC
DFvikfiDiDjvIYQ1+lr6cR5A0u0ewnwluxvxJFL+mBQDEAc6FxzdAiKT5+NknmxF
d6jbZu23DtG9kdJ5Z3crzyXtlTlS7uQnrgVCCKuGWAj6kD2v6iJ6aHRFdKh2BHp4
jN/Il1Js9+u6XfiXzTVUo7F/R1syMQZV92idbLnldEe1sTpfu+y7hZ31RzWOW8pU
mfLv+BoQc1DKsJ/CDCbZ6e+rpz1iyWz/yNUk+W+ObOMasXZHBvCX4aMunAQiAmy7
DHzRTEcPZPVg4WqXyPzKjAYwyGAZ4uLV1/m+cZPk110PziEi6PrJ/xuRNzGi49il
WFxtM2eggrheaXjc8RmsxxE3DaoIESrZx12V7VYQfpUJhvQ7It3K8xqkDENQIwb+
Hh4gry5+no/Az4aEnDTkwyxJ+HBFJG1UrvyLc7ibWdzpKL1dUwo5UoIT6h7Gi5HC
XtD+cxDBfNBN2O2ICSwxOKl0C7fdznHR0PSzCpJbX/IZGv18AN5bWWeHdPbsvBlM
Mn9W8zoauD3xq4xSg7GTpY3UytxOYcFnwlFk8ZNtIRKbphsG/AJVXwoTHdXufk25
JyeyZ0sTz9sdCpOFYM11Y7jztQeRwjrwvOqh/uKRUfAemIu+zWEjg+aOgBGgoD87
h4oXCPx4miv3MNySUIojjKfWk6WA8lx4nixQWyagQHDxr42IUKfotKjpDC9rR6+u
V2XozVCrLMVBITNBd5ITChMAiNyRTbhinDFxxs9tX+alLlZf2k9c4/44+uEjS7w4
AGdBtx4Rpw31ofZMyAY78viCgSGtv3oOZcaB1llztHlSjRU938w1lKaEhkMPDLwT
/jcQ9WjtddB4vwXP+YfOW1C7Et6pofVi31a22Uie0Iqvh7WIVkqTdJxVPF+JEBLT
R8wLs5sEDoETo71uljXpSXss/dwChh3IRK2RHoo8My3DxsW84OCgmX7sqN/EsRu0
TSXpSGwasK4De0fjbOeKsV9of5LgOT2Dh/ceVaBMci0b4y8XJLgjsaNvLK7qJKeT
F5R539bG3IParL/ma0eUjiPvLJLtt3RChdA/cFyV0ZN8XQ3m6xFzAoWTKyvZUJNT
vlHZdyGYOHXvl+0oLksi6BTzUDP/tu35DlYWZBtJVonxihSSV5i3XPMZS0wpl32A
8v63Re9B1BcDb70UBNG8N5g6ZAVQ0YbpCTyGfMD5y0NSUfD0WfHeO8GxKqi0okeU
pY/lNS88+kTynNvUN8aFJhOeE56By6LhpmdJIybCSfSkya7q8P+Hai3jIZ4kNnHf
hlJHJBbQmbC5txetdSW+M6uWn9x8DCZjd3RNXdcfpcsHcf75eovWaRbb06N26rSn
iptRGwsMMeOzK81xDllm8zLzypGuvarpO6Yt1hjuiRPpz3ecBhdnXFo9RTjAjprp
hg/NTHIpm1sRbWOrqHKrUweg5t5xKf9A9qcb27yvH7BeoHTSTkWc9k9Z15XxoiOL
2DbVqaz3RiaVsb2R/ZYB2HT6YbGSUYMK8ObDfElePtQalN8SU5g39bTdjnzB9p7Y
BEK5+BuoehHY7tjVg/2iEIU9cQcHhbdPkM35RhEGuiTkmuSYAkZSHjjxz2kO4tuR
TjGcYYhE+g+vmeGThZf9raTB0MHyc1Vl7Fdwa7l4JELXCkYbGaW9Ka0evlNcuZLX
/6xXnEiara9gDjrjhxI2rljg4Hkwf7oYbppJQupig9Ue0P7ZglACzzFsgKVYM4Fc
WJrJBbcr34Q3rVVZdPS5nC6Tke2CSGRLENqreqB/b5NRFTNSjhgYNUjw83dstwL5
HVrKoQeE9cKJQKeq5uEdy4hhSkWuL4xmK3t6eLiNO7rCjSP1uigsSLFHVVmGD3zZ
9sfkB3389++6ZFVKO4XOHtQTGSlrvCBCCqkh3pA7UFeTsZD9JT9bnok0dg2QL0fT
YSH6LbXJ5r0kmn3vLhV3MJ1JIOebLP13FQWY9BPsIEla4ttJfOroXpYv5HKGTwig
7XBmK5Hm/4H+31McTSl1tN6f7xILIa0/+7H5pZwVQQ8yV7ZgdHmg6Xv/PqtehyNo
aJs75Skz4jvDIyNizWgoHwKMAEoAOkgIRv+cnyZvhSxHZLDWDwZRNIcH6twOMKJo
tKUBVrjeRuq4EfndUkj51KB7gF+s7YivVAnO1X4EIW7dbgUAL4ZKkBxSveYyi0Z3
hRtSBBCEbjytpntJZJ/b2iSGA3OcKTDzbPe41UWKTWxDYIvcbZY9B4GIekqXV9as
fYcJxu+VqN3i0sTlvpVPmRGsZ7/Md+Ol+HE4dCzaKhy8ZKbeiYqFgu7vnPAPtT+i
jsMMOYyuNF8tjEHGJiNuC5hrf2lk3OGON7CdmvSdNOtTxLfDz4AMODeZKTb2Mprg
nzDNErjUU8+YFM3NPoC3/uGJUCfZz5dEulj20i2Y6mZT7GySrABPaIKkNkSqB4JG
a88x9pHZNXiWfa4ogrVD1lCi0O0tKDjq7XABRrpYV66fIuGfhahX8fom2tnxbL5O
BqbqRRnPn5gbEAUvyZhPoxgmTlhuishaLSpoh/zzVENGXIJa1hLIFDMc1bth9Af+
Tk3LkMXGu/+gctfNCcPzVDHcup0R8TKK/fJxq60VXRAx4+byH/riGNT1Gf46kvNh
kzgwj1ZIiop2IzymI6NPzttjA3MUn5yIjYwJrKOnv50aK6U9NbKopytqXBiXh/in
HQjxibmewE2MSU0KvUF8EAYqKbEvPTNWAsadAVNChBPO/SIj7gHohKcsfANQuMgN
CzdpsdGBnAv0B7TPnfxCrzq3GjEX8qeo+daEdKIlv6q4uia1FH4cjMx5DxB5lCI0
cnBY0onis4UwopCNCBSde4t4p2vcpZZEXQAKSN5wK+GlpflOb7zmRXipW5Wa/pWW
HD8XuHYxxHccLtBAkXGczAeT73pLw/+wyYZKdULgWPsvr8iFxrUxm1x6Mes4GOjg
SwgDww4lpLWszwWzDmn9hIZs8VBBEt7ZxIaoKbA4VPVvOihBJXVtYzN8u92cOQya
jexTgD013kNU26Cgb12A9uVJtswbbvdN3t0oHfwhG4Pcahy0pIQN7LUOsBSyj8uW
bU5U312Je74ZAKgrJ0Mw4GBCkiJH5o96iPHr6M3yK0fZ22E5KiHmBb1VG21TfF09
yASSUcnWiOtSY7TjnIgGd4OI1A0QhYWeuE+2pWpcMaUv4xxIyjZ8GujX+R4YXcpK
vBTQb+sdwe3ZhcDjQRndx6crGpghMczFLq1kpw/AGXONMQy40iNBlGXnV7QUiRBl
HZM+NFMc//jocHU4phQaY2vvCjlrOGmpE4jCFlnRsTXP0aY3MjFgrbtBMY6yXtek
h2J3CZ8CFRNjFkJIeajzEY3otphhBKwETczuZsEf4K+Z50IaUCTsXY/X/I6gnXQj
zzOZyXxmmpEpskcNQYo5XRQSnpNlUKBTMjFelBG5W3R1o1vXAuLBtbZWpfRMbWs+
X4f5D74jP46SL19dRdTv6tWTvxJlC2HE1lwPwNSOGBmF5f9fkcbkLGLtJIE3qTAJ
EK9j4ajc7M9Z15X+LTDTISyIWyfXr18B1hHCXB7pW27gzF7yc556NjkfwqLLDa2Y
UUyR79dL8jq84/gIFyYf/z8MBoJLczoYT40eiEtrwzwul837XJmXDtkU/vPdcS3Q
SoLS+0LaMRJ5lv/cRlHOOOvRtoj0+BNcBb4wrDYR46AyAEaTqSu3eNbKBIB3uajz
hmnKfnuYVsF/RQYycElGdOeV2vmrcJxqG1tdEGk2MHh2p1jCGOQ3FwbOUhG+j1fy
grL43KgnI6nldHb9/EPv5coUFm2V6wFDFuWD3fLFfOFTxxqBNMb05YcdA8GOlZRl
OoP4XhNuk8TSRc1ZpBZJAHuy2UZCmRm+6o1e/aoe6PYMCqRdAq6yH+ctOgjfDM4F
SJ9WJTIM8gMgq35Xf9sJ/nSQMDKwRHyntnKIkyuv1AY/v9ZsmdkbhJzEEzYmyDId
pZHvafx4q2IlIU9PN3K/P9mJDFA8N4xNSuTwqgUh3t3cpLx4olBQDDrBDuQ4O3Mu
D7ykVSZcguRXcuexXnwAm0YP2uemM5LydPOOe/GR3hGS5nxAS/zH6Lu2GWWbmjUr
3to70Wd2vKuwYWVdIYnH8B3YSOQHFAl9tO9MI6/NBkZkgA9EH3jUC5zn1qg48g8S
K4Vx5QARz44N+GIMCWu1HPEbZs73ZasyZlF/56SlRZwub5u9ZyUqLR3USMTqGlRj
4/Dkw2rT0u+wUknRcVb6cV0Z5tWq+KnsgryWOXv0nSIoEtXcVx/5YU3gz0y+P3av
AUSBfeItmilCq/Q5mloVgswGG+RxKLdwjRagEWTG5vngcNj4cAKVuj36u/UP08fN
oESC+hoOjxCVPxz4o6B+K8MzS9f4rwhqs92D8P5VzfEi52iPSUYpxXgXsswbSYxS
U21g5ev650krYDVPp1gr27QXSpZcuDVL1TeGGV+gKy1Al2cGRoWz8PtHvDefh3zn
49+cRC7D5TSNDcBNljXZbznffeCtvBAY8GVhDMYHgLA1k20Xv+cRZch9BESqoM+V
67JpI2Y7W+spTB+5zIk/TlOkh5LViK9DiW/QL549r4zP/2AdIMGPoESmcXjtV827
ouzk4WIusVeATzBBdLAxpToo/mVUprchMpsVULD7B5z7vYx23natEfzQVp+AhQGx
m6n3862WFAcTgKoDRbQ20qSIaz3BEkc1bGrGkNuaUIXtJHpCRw/awoEKWAJDGIFY
B/zUEWAENhWuumv7mY0nmTBhtjB/wc8ISe9ee2bEJvNIWLiVJ9I99bmMVup48+5q
teHf0fft4O4LMwwY4oVvX99g9qfTRDCroja2lGo5SER2dk2rV65OcMQoMZfwJPxJ
fCF3ZIWWgDEmSOwwppaI4VbcvH5UPtEeVaukCXD1vqQ6MYJCNDDTook6H+A/yaVB
whBpMWAXNEkQyEkQq35qOgckms7OFigzhT8KXd07+grV02HgwUWfbJOsbD/RBrXJ
Q/Kcy6xWkaxHMtjyFUt6g/7zxrM+ZqBa8hOv9cdl7xwxViVZrq9aH9T6t4AglfUc
hG40dftBgLLfDVia3Yuy5x3vXiy2/GPFXPD6K4E49vpNJYQ8MmXBnq3OJgwsA0eW
5TJNrYM69MWrPQqBuTr8gIFGSPhjh50D9OGmsL3iPUq9Zej5ckuiqPrIG/0UALGe
USV8e/TCd/h0P1biMOY3hA36wmJE6aXlKr8XikO0KBkuNDJNgThv3DWS2tAqbrTb
gA9pp3Z+8C0KdWhW8DksmatXSSA/PtJk/DLm14azLX+nEcbjtWLZv03U2VVMGJNC
mM820i8PJKhOfTUS7/91/+tgyWMWDOixA6MXeeufFxCubC7OqRnoudGOqMsz8BwE
PmztAe0BnBluKr8JIGZm5H+hzqvmaUXt5vi58NOB/nY0YF9gIRCW1/KsmykWutAD
kbFq/3ZJx41KpTYfO0LYnUVO7ydoB4RxQtwrAo5ftQYuCVX+uEXzWPAbP2eOcxnp
BC/lPPob5ycueAEmVQtmMZujqmrk1mVYxNMEFVkCsWm2GJeN/1IZoyNorOJqjWPz
ecYnqosEeZmBHkKI69sX7DBtcffV4R3UXzSuq5nHergpElzExJBYya4kmUxrVaBC
HyN6RZNnI17mWxVXP4+fASf/bblGTVDY3W3Z7XGVLlBuOyRnH9S3f5Gaw0D9FjXg
/+DB030oi99IIfktIJ6Twwr0a/o35Pv5zLJgShKMQC9WyS+qqckuNrAcS7pSsTQ6
1hRYSgUd+vOugDw/s+dXXXmLtLJtqmtltjp6bNoC//FtvT22I41uz7jLWJzrm5FY
bVs1QwUt15yiVtMWyOJ26KzSzb+E+ukB468t+k/iLatxiS3eTILl9EJI/1EVWydd
X0OlnFmZyn7yakTwwwtepmtdcJHagXGZXtBU9NMhafRXeafh8P6jWjE1ZWgKrm6W
QyIyqYZX7yEzH/oB/F88XpL2PRYtt2vwGpd5F1h5JGxE+jJ+o2rJhlqKa4QKwrIy
ZCZ8ORKoTm3JhEQLXrTeyWSmev+FrNwsh7RMDE5Qud8y93/6apVjrcDQsCEMb883
P/oQNPHCcbu5zAvpDw4Jp9fRHyJaJyBc5X6LwogPiCkda1ygtzoUQXp0n5sesLaq
B89mByD6tyJS6hGNmP9R5Cy9mdILnf07sa2TOwFBMCt3nf+ry+SVIQ3zhZwP0/lR
lXKCnu0m82X9+/q7oBd4RIYxGQrw1Nw06eSm4MzES4Gm16yoJiPL8ZiVUdv12BN6
hs+ef0ZhHlDbhxdlsudnIK9AdlzI+bPQ5jkrZfCAuqQ6oph5HddWcUDq3BwVRIT8
kI5R3R28+TQ/NwRLPXt/HrI8HBLXWIN4WUBDwRCnz0PqPKTmZ/dUqHiPw0gDrCGg
4S6A/F69OuvjcEpyJ/A0kqROqmalRcCHMHUaSRJYGD247C3Fw4UqVrGxUA6eJFhW
iD8e640NaoW5/z7VI4F4z7dT/9PEPmbt4VzBjDwoUm7528CDUC8as0xCYRXWSbu4
yJSgajaCv6rNOnEIrVcr5VbJcxltFgrFqfjqMy4b8sOQ88mLv3HJZ0cw7K5JS6Nf
IzG0lXXPxlKWDL1urRM/tO5KUcmoOhlI2KePZFP96STQ8wD+DJFFTjICU/y6nqAm
nTQrU+TXORGTHktAxaxvpMQoDrv5JVXyqxvcMcHNo0CzYQSHBTIamLO8gLVxb0Zc
1wUoyQJ3i2zQDgUT5vNZwoB/4QtBvlWDGfjsdTkHpuLJjqQM1D0WCrQFLbUGE6bn
ni411nSW49wrBZGyvUWH9RhbnkBOdYBVR4/0lVf/lFzSwNtnNYYQmggHIXc0dney
Kn8VIV8l9paBmSnB63ZbHcd/iE8hpnTomnq7X76p5PMflMLPxJUqGgez5As+LJhT
itViqy/X37O3O38H5dh4nV1sDS9YC3UIQEeTjxMi88IxKGYMnwrOBNNQ9JPaGBNW
Lxa+cjraUmSQmhUS7qMLZmsaSw7oTNAk7kUZSJQFNaUNIidFcOi58tyFLz0WgrEz
LO4fErpjYVWHMYeoZ4IyHYtKV7bH6xB7UN3xM9RWxk+H+P4gvdy8CSI5yXoVxPOl
135Ev5ewdLi5qee6Z2QpClKJVechyaQ2pqfkkRmuv5JJHdCImx2aGPhFfQ2rwhOG
qRL8t6es1vihI6bJt3MQK0YsVLwTbxk+KD91l49ZhKcomh/0JAfwEY9cKLpn8B1B
TBZYiK2EwrWHyQNNqQA3XPbAJpIVwwf9kVgNZFrDGKGNROwsWR7ve3RZNulS7TWT
m7IdWHhHVLXJf4kIovRQhgRzZfk/XLmK0hNaXKzkobFlON2eJEdgoMpkCItcsrxV
p7KQEzV9/LczZnioejjC/i1NCc87SBxviuM7XsbQ+6hN5y3m4GrZJ39/sl4VF9JQ
8s6k2f0ck84d1N6rRQmgNx3vDRSonFUDcGOgRbGbUVcvaEKKOn3Rp/cAObEICdZs
/M/QMK53kicUPjQP3qhcC1gpjzz5qJUpY4smWtkwBKIUKcasRRjIUyxjNp3YFacU
xlCK1F/4ODkjl7bLPqQnq4zmy9lPC4nvLm8SKiC9MWD3Lp+ESFXqKlKzw9U2Zify
Yz/Lx+OaqPwn3rfrF33cHNgy5b5GkbefxogXyB2Z4WCSnNWDvYDQVe1BLZqnGyIy
NEVm8rxivjv89Qw7qHcQMdbYPTG2yyWe/9uZLhGmPE+zI2wr0Cr06boxqTJ72xNm
Q6HGo9DwsQesieg20csxQ4LeyXt6nCCyqnPGjWt7ZbXJeggtVyU/4ut+pLjhq4Jy
1QKbIcvnZg9LAKSSFgdBsoLflC4V4x+f1JQhAZjZ1KEVlOEgFVCErCMLwEOS4yPV
EO2hT8BDYLH44Ua6+JXDX4BIHeaweWxtIrwZRj8Z24ZDCkmezaWE62NiKMTlD5uK
vmZ42C0F5ganhZMV4I54Xke6/cwvijUdkD9JBqFMDoxFITcs1o+hlv/umfGHO7+5
C6zfgFdtl47iRh/sG3/u1hKjmXH79LeYGZ8ncRAZ/vcyPw8EBhFrmBfHdgCD6rNG
5Lt6/2ATa9iNrCRefmnHZO5LzB63e70HzCDU8a9dnQ7DaqInaBSExkbGjKKyOkvB
eFyQJIu2SsIpe1Vi4oGCnfozaI2iFuFN2eH/DA/PvOLf9T/RLX8GDpBFrj6IduHM
0NiQrl0qMci+qnsBKkhRzSGIPPCBxk3VQEr9Mxc42He4yKzSzFyHbAzyRPxVKMbZ
TnOsqltqIMaeTmIWP3Tq94pDgXOSqTXnOGYuRoONU2wMrX3BB2TRhpuYhlMU6r2Y
P6hFRAnt0vPIQ3Q+0K0OKQclKKnVPQ0YZ33BA0E189oBij9QVKuJADDb7wdJ/B5V
9kyOxLqIKgYFtXclY43NxuB7AZuqYRD6Jhhel4sM/ONZ5albzb0XNVOX9ok0D9y5
DgNnUxb3vt5ZYtMyuiXRyjgSg7Hm/Yr4jtoqJ90wcLUR9iim0NlxgR3x19iJ8UGX
91f3/zne1HRL8V8uxksi8QOmUQXRBIN6sOf/4ik8lCsSWb2wL6ie8djC6p7IhPW+
5ZMy8jf4/qwCHCw9e8nO/S4kkqFQg2kGRbuu5IoPJyGaFKxlQDv/QXUEVy528pEk
tPSuYCtR4eTFylM0xUf2l2r6hjykuiu1t6bh3RCh/4QM/OjILZe0ojtq9NbHqCGM
hGwbP8L+GJ4uDGnLfgWWZQvjBDCzwGzjXsYoDqBpiifQ0hIwHioHmng0rKr2O+0c
ayVYgh/DUawr0JVt/MHppvR13YZTDlWA1m94ClFubnyGCW+58w+qhnWVOqJwYbUC
a12lMm0gCnlRw+wOMtxPCPX6UhbxRktlSSlL4Avq9NGgIkAE7/O1ZKvL1v2FpexA
euzpTp2pTOFBza54BWXjtcAmnLW4sdbJ72kKRwBFBXupcYW3PMAuDrgxq9TJEhe3
t7PF2lHnuW95S46/SaO7CZa2n4cw1c7aLFx0qirpiLVipmpkM8zFbPS7t1CgF3P/
TMyLJbJqkeT4R0KiJev7i4J3XTOMT7o/E1kpnNgjhJ4eTwLC1HKynWvTgCSo9gi2
aakhHDqoO9nvn7No2oKSpwfr8cb7DI51oGxjapNv7NTVnYUFcgOM6CPQVXujrcJY
12MFLOL4j0X2eNzuIjwctYzIm1rQgW4bWMJn3r6UH9U2H7KdwAbnKCshAP8mMbzl
vwD79/56+c/fYkjmE2NI8GDMLTU7408pCrfQ1+42j9JjbfeI/jlEuboHSAhPX3RK
vvFkuViTZ6yaTZDmVjbyrdPEs5E3hNg6nNZ/43fD4LriNN/K8KZSbjPzEvk6Kch6
00Pt53RvTogtQ69MVxsGcPa24B1BFz/JT2JsLDILYQJSdg51oomDY6SjKL5Ejgum
xwEVdpp3t5O8Vo8PPlEGpp8o9cu9iO/+DuOrP6u67dI3EbYDTKUSPhwv04uecu6O
JmL9ZLXJWRPFTB3wlWRalVKS9qcyjs+YswaodBbtyaDuu2t8Ab6DWWCyr8dLokaj
Rk3Lt7zbF8F+r2zrqu8f9AMf9+UOyxFs+Tb5Iuj1SFa3PsjtqYGqgYLFDrJ0dvni
m4V2OxUqG+CtBsL6Rwzf8AfrlgyYQLuyH8uoPMPp6BW3SNXvxEA2Zg7/Lt/E5yHM
93E/C6BlxZWT8irdTcf8nHzND+W29elc8JkI7yZCriqRH9H1upRRggS59i+Qil1q
kgv7tMQsQNorRcCTcTD0l2RcIAZKfAd//F661SRlNf/qdzbMwdn3eyRvanfxBjuf
IDGrYS2KlGP3K+ptdmvcHAoQp1lSXA5Er4UvwU9Ke75Z2vjHlhmSVHEmiktNYU8+
QxvqewLyvgHU8eI9sXRv84/eBF4etSSpYD0m5OwQNYc5TtX11f2TIPktlGSLg47c
O12rIwCv7YKVR49xBoipL/eGbO4FrVAU8xX9d2i3Z+guk2CN6sS275ZCoig/dYKf
3comPR76fJUmSMOFuEAXPFDGHPoHixutpW+GgBh6rwoC2lhirdJeU9wDU8SkpyIa
4zHGOck420N35dewWGbGUsv2Z64B/A+20AOdfzWW+lQ15F3bXV8204jMqwM/3jKR
b1Q3gDGPIclszFSHU5792+DXfdICtLoXp5ivZ9kCKQcYz79fp4vE0T6lkMb7yss3
IFphuOIg8he1lo3VtW8UFTcjriXm4r868lDUVne3rV1XAaoUizV53CfjHpGjT4Np
Y3st2aDrjCwHxt9vpU2KTelQM/KUjN4NvS3vWGEC3q0UerPI/vNI14d0LsaxU+ja
xpgcE75iALvt6qSx6LkyWweJ0RAr8S7ItyVPCBR5t+KmxG04pFjo3mZlYNPAJ7em
RDXpSWaf+rZG+c+t78YyswzN/gAfsKRaIcltRaTQTLQEq3FCXZ6kVL80EIjs5YOI
ofI//IRg3sSx60Oh8G//XIS+PmRNM3KYwudx6nPwa1h9uLQdi3AbsMjCieNatXo1
jzdqvctn9k2Inw2h8mKI2v0Ffm7/3QmZeaF0HDyQv2D9tK4u5fnoKf/R0/NF7hi9
nbGa5Pgxy2cu+BrAHzvMhnl/rWk3koSziWIWCGLVRhkgeOSpbvRfMU7AEhGnMstt
jXpjXZu0aaRAsyXjqn0hsfroRrsE3UwQU+vhY9ZGKflp3J7+sZlUPxhaeLlsPE+S
R0DRIJ8augJU41yhPvmZHLBrHbWto3t2QHKKtBQUeq3igrXoWmRmLA//SpuzLCZz
mZp52WgsvI3gCRbsJbHt2Lj9VvlKdj9qmM1yP2ZumkTp8YbqHB+U5kb9qprnlE5G
KV7fd/6nngQ23xgFTYiYQ9V0ScFTKF1ybUW7qx8c+Q1pz+HDtPwItey+J6R1WUE6
tnwrUjjML/UNm9bgxE04j8FimzEciisKkDi+AmZWLpWpC7u+4dcuCH1B4fWBTjfT
QJffcJEq9NxWosn9zLCRLPp3m+NGWoheeEDkxizPOTVT+uAXXNO0We1MTjd1ox6r
nw7ZG0DSxTh8h7p9eoHFa948AMo1BfbVhPQ6bG/LPU5rS6cu4JSMx5SoVaWQz9KA
ZYDY2WZslKXchcB6qhRZRHg/azSnzrGhZWiadMpYjd5D0A8qcMkIbc2ILm3V0m80
RlH06xwkGQXiUJuU4OjqnQnhZp8z+RJm1DUJU3KbdcrlGR3B/wjGV3XPhgfjcvEx
JbWshXdDbH83YyB/qH8zfWUtbIHafp359WaJT0Z36nfKQ61vrrwwGcjZRFkwGmHE
fmvuEClMITNNasOJj1mNWyiI6yiWpcTyjw+AG3bFnh2lLRIsRlQUm0d9iJEUf31y
VerfuQieuL89P0TavIGfkIkebOwePW3ftR235U17YuQ5cQ8wpWPQK6MB6DRWtdRX
M6kMFUDrx4eWye+TNJ4FhXHagEKMpf+CevR124xlOSkaxqaJ19Qwn87g09KxMA8r
xMTZJF8Yd8xEoXOvqEEMAkI/saInTn8DXQzy/5CLIzU0i6+bCVctc4sgdN0vxuxA
gv9PbvsvqaM2TRwPySHetePP5BX7maKBGKQ6RbwSiQyCG+8miLVGewteNEHfVhpB
FPDolu/jZairYAULgLyy5xvlqx30Wr97PhK4MMRKbdDPWOIDD8OhfptM8QctPqCX
/JnfJNY1mbO25gMbOHQaaLOfoYWePMlguHss8JsViq0hzBzQ/1YW2sCe7Fb8Qkgn
AquetwS0mHNs3Dh73YiXH5aXdRvGQVjxyAIVOspk0Kq+6wbqygOycptUJdVCmbfP
hWYUIUCtXcCk+QRGZKRigbfjtpNTQkvxvVHeCEBFKQRdpeqwgdGVgN60OtBstH0Q
GGacCUROSmx4lJ5Jqkg8bKFS8GudF/k95VoLhIZDCQ6z8Yn1dHLBHV/TKrY8KaVN
ecx47nry9pCTjq3xyUeQgvVdlf0PUGEEG3cisfKWj331atacx+HkkSnQ+yTa9ez3
L75ShUA0fMFOpLpmtJQvDUOnrcWU70pmIOHEei9JCgF2Lk1tzOzATebNc6b4zHvV
jwVnzeJOB6TYvFYXlSt0tcl0qOlDSrFyIgWJFppJRbuoCeDWASwmG5WAeoleYuzH
p6lmPqZeLT75QCkfIzJJgt9rDpihVyAD5mte6YUDRlNe/MRjVPK+vc3Mng+tNtF9
NOWkTEPoCpHkoc81VckzFoXdWy8XX2mF3rynh3rAQnBd3HNm0FDRsDl3k4+MfO0+
tHZUqdfqvBAkh5ojo2YRFtfGKELpxadEKTCUAbNxrOPG0L7HlXmy3Ij4RI/Squhh
qCnSD6ivjo2f+/9OUJe37cSQ81lWvxXUx8EgHo2mMJt/rTVJdASa3iRuVp/EnnrD
xUyU/7fIjYpN1kVPgqfJG3LQ0Ct5QQzaTVLH+dgNs6BryAXsOd7bKuEDyWA8AaRD
Z44+fwh7hnmQ3J580nGDeNC5cky6/fKL+zwMSsli9XUYLuGfvKydKxJLd4CeyW3Q
KWQHIvpP8sxi/lNpQzpiCgaXFgzeq0qsdrZK39neWEW5dgy7TJebeX1oAvyalOdO
g/6oH8uHhtisUZstnBoPpKi/1bUcp8xepWr+fKDF47lO17LqnNpP9Jff2IXXI7EG
XVLOeMfmD58hed6BjMABOlBnoQfGZuBKeaJAb/383lHXPNhjHVV1KTIf0di0beX0
Uw/X9UxNYCVt5oJtv+pLb7GRnXNtkzqZ/BJV7+j+v84iR3hIEb3zhQG53FzT5Bcg
ikqDrU4mtsC3ovxsSIM9n4DsQWDzJ5R/datH5wM18nhylCTw0i/QEeyBBCnDRHVk
UiIButYrptjbR1rHXQBI9KojJn6jFYDZWPKV3OnGxuemF16+Ttekb6nK83HZ6CwZ
z9le41XDE2s9d+B1XKuOaA7Ah1t9pFtJurPb0eEIdbhkSKPs8fK+HRsMJroYU7M6
yqlSrhWxttTiHtWdL77tYmGgP8gZcZa4zglYXI+ATTIcSxvklo0EqzEgUnQ3BnZp
TPIUldLpxac7GA65o6W9qIeuqQ8/XYq6hRYoeSYe3Rcb8GGgOOIJ82Bl7xCGYTFt
L4Uqm1fSYU35WE8CQ2SEV8ltICtQL7DfgpAzeCwpfhQKJZYBOrzmhNXBIzXZ9p/D
YtvGRKGyWF/8E+jI8Wcw5eMj/DZdKtGjmS7le+kAnwSef1dFm3tWGP0fkrSVDEn9
jIJLWk9KEKs6FaqKKK4ApWFf+4M9qE/Gby/+ECSkiugSr7mnXgKJfv30ITa+EZ0k
qbXq2eyE9KtrMGp6EdgEd1xjdaK43v5oJnyS2BDEUTdLJALmml4YL1XqKaZCkFIf
BTpPokID6vdLidD0nhkDG/g1tX1gZjvEzEh/XCr0phAQYVNJo7x6kFiPECUM723c
rufpCulOGH3/WHuOgxMhBo4YccGAoDL0Vneq4B36wTMCG0du2murKAm7gUWsGfQd
rvsBJcqgLXHIainQQTaYeGHMcs53aud20YrgQc9n4zxMc3lLoJGBC6Qmyp6zDAny
zXAbITBv/wO7uHdsY9Tx9XjkCOcMsQF4M+423w5UWwn4GPmPepKF4y0UV/ptu8FP
nZkbYxMfY794rN6IcFudBy+NOFZhew4wAL2Sxu7zFg2OpSeHTnuHz8PGAZO5DKXe
5YxJH2AlWhYwhPfKMQQfO0b9P/pCDUz2Jj3vCNNsqmlYalBQz6SvbVfXcqnLVsVy
NpKJmiPoR5EKFR190snQi65nvU1thiz8MAS3MCHAW5/uUI4lhk4YmbkVBmfYxSaA
Zbs/SkW+wa7E3tCuUsO1esSTRHDBFIUkOgFivuKr38Z22ftWYSYSHwLf+EK7m2LV
UgwVNQkyv7tifsP4PUKVM2+q2LFS6QM3MduLTby6qhi2/ghKp19inh9Wyen8Y+cm
xCR6WgTXJ2wmpSEvQskmlDocNqcvm8BPWkiVAV98EZ4iBBO5X+JuNqKOJul+b7Q/
PF0fKq9OkL3kaO1ywunqdVZfS2R3OlWDaNAh2k0+IAliduK/mONqUBLQk5XpPFWs
Rlp6aengYp/Own3jgFCf3rGQO6PNRL7VfFEdmBr5m+4FHQIRTOMJsigM+ml3Cooq
smJ/rP2jW6BQ/y1n3Nw1m1pnx/O8Fzcanuz3PeAv70EkUmsly+omF5RnXpQiofFj
DI/LWSlVFivUyAeKX/jZ1F+Tzdk5y01j49kIEIgUeFemrB2UzQtIraCWpM9OqPtN
hb9KKh8tXAsigm/6coknv2eTxgH/klovoiip8nh3TIxQIGoahLHKWc455vT5GyvP
sHrs30tLeIFSz2RzCDEu+Z1XvhUwD+8BNKkZiUQ/2UrcC40OJnPADoMlupHuEZxk
RGGFW7XXkSAtrJ7EOivQppb1GeRfTLMrxrHfzKIIcrbBgG7BRGR0iaiK8qV9cqNO
y1Qcz0WLi2g61oEW/JRaUXPc3FbZk48aw8KKSDsYpvCm3ykiBGTpvp47mLdBy8fB
VH7awEVrntHreN3khHc2qVBY9D0X4htJznqKQMh/2YlDc4zbOUpJ/b0Pcewg6TAh
N+I0fjiKV+cZ2G5BFoBZ4+XrYXSDZprqb0xMct0QUGWvRH5p3nL8bVIV88DQhJk6
I/ZDv/qcl7nYzWQ5SJXMUCnlG2MXoonimyve/OZxcs3XX3flUNWwrjths31j5dVI
ZHMapbsbynxLAgYM7hcz5bAAS8VvGDs3W3eLVxA8GcuBm4moFnQxXPQDEELmrcRb
Fl4vO9zbBENpVGJpkG4Uim66hepVOxHg49VrrKuMAi1L8u6jWD8dSYUrH8W+whKm
NmX65GEEUL9HzNiY3gVeHJv05EN23mhjmH7lwjfW7VY8b2p9lbKwa2dRj+FeWWEn
Po60Kqew7A1y/pHUKLDxYQeGfc/4q8/3gJI5e2YCBTeW1hoa2Ug16ktVPCK0tYbW
Li5wL/OKnm85SR4aqbpJdBi/pezA9SPDuIeIIK6yieKPDzTLkqHSCfYYIuA3N1tK
rfEgjClG/83OqIP+NNA1S7CMwVL2v5LPtbTh1mIZwBpYec76aQDSak/w6TeuGWcy
pb3cY+E130oapsAyVKFdWuQ/vVzDQNp0TNRP9PPYIrhbYE1EeXM+wvCqljv5Lp02
Xc3ymxsL6N48J38Zk6Xs6u75ReUxyE5lSA759ypbSiZL067q8RXQGkf8fsDCKD8z
kT4vdG0f8lPLnqQnIX2v3ekG3PrBAq8XN6tToNvcHma+RpijxXPkVGO/xPEPpZ4J
xRKriGnMUmsX6ZnH43lAtWKV5dbR+Eolnxe5B7gONTwd/MvZKm7cnlTRAGAwUGfV
XzMc1wX2E6yQctOpvZaj5O0eBugXkjzfWzYyJ+X2Q7lQPm3/BaAwhTpwHA4EP5z9
DoLvriW6D46zcufzDWJe2ZdT2bFxeULRXERjsvvO3M1+omZOxShteOSLjoG+e1gx
EZW3RbynaEHyKwqq22rkweTYa0x+IS5aaMSXku9JeYB0hcuvOEG7oWhKFT8wvBdN
mHJvp2rvsIaJ6F3+PFxVvxsm2XH9DZyNDi4XY/EDyGgbduyDDTD1ZdYX1fsIUOC/
hnd8igtvqMifM9F9qzEdgsvc2fkaNMEHqdvqiJ6WKmWKE6WoB1t7o8bg6TeznsM9
Uma7epIAZO1D8x/5xSGnt3a76s9H5ytTdlpPkh5i/buo1E54kCRY3YovaKH8g9Fx
22TXpJ0fAlDYTV0TfyRSrcVZmz8sYejOEoDwI6xtwAPfRw9KFJsuso8tzuxECMDY
k32BKdN5KT6lEqgtEhiVluZoeBpK2SZu5Py56S2iIXRqWTl/eTCLLL2fjduioE8J
c/JEtaI+Kj/WqONJUgVTA8hly3+mFpifKop+XyF7bFQjdnVDIBaH8k6u9px/Th8M
YNN2YdGNg8p+SH9ykeFOz4lblhtjgKXgksUWuEs844u5nEQe89D2vETEjKYv+8L0
jpbBzvST5uTMc9FQ3j+gsokHFgT5MN429MgnWvBDlfUlxru/DTgrP3aW9ARUIbfO
kYCC6OU+CBpW37PdT48/2kKjYcZwVqT1U2uty3egSz/gpjomNtK7uEwkcdADqSRE
OrV9ovLX9fNwwZKASgck/bW0qwcq3N1FSjaCIZqAijYSL0lu+RQQynRUsT2CjTN/
me6xeO/CGjyQsmhdhlDA28+j+u1I2VTiRFXyjjbCPAPacLRWgmrZqmA2QwbBrHGS
iSqjZU1V3jJSjz8w3kynCPFCQnfRn0XvQf7gwR6u4resgW99hoEdE5/jTAuZ4Mcg
r7esiCnLvwDiJTiwqj/evvpDGunHtw5hWbS0X2LJXOhEbn+1Mrt3g49izoMbSFUd
1fR7TIrJxjzbBA3RmsCZZAPJow+OhAIOChKyppr5jbvyG/faUsHQqq0+sYVJSvH8
stRKlhxgYuAbYu6lfASznZelUYXt7DGgh1W1DXfsXwUR20/9kKnq2nTO07vokF4N
M0RfSRVQrl5fdOJPgN7D0YWH6sY7RxAj6TRxCTM8geYGSipP9W6Vwr3hAy97V/c2
hEBLu4Yl+zLlEph/UiOv3UXZJYOWty4uolh8SJWtc2g8ZY3j1xPFAVhc7GTRRSX7
1maLSVueteCImBj7RfesbROBbHG3u2sGaQr4qChOH4hUmcSiH7TtservGcrnI4/T
+bz1WlGcMHO5Z9CwruPjCI5UbRXt3CDvUnuoYJ6uz10dNCttNliXwq/RqXy92RSv
BBnJb4A2Y2kZ67fO/rJZxtHmxDC64pByrN2Zl7GgmKldmfqzaMuminuwlNe8AZ2V
N00YGH617cAi3To1tFzLiE1EHBcKRiYN2DlLHq+x00/GLBnXGDDTxUApnYgVtt2I
FbfiL9Gj1rrEj7bRn1EVSCIPK+wMNUdquz0Octr9sBaO6R9iVhUI/wNFJqRBgRJC
a6dEz+J0U90i7NrSLfazkVL5t5iptGbM3AXKFbCESPwbSKBIVoMre9TAebO3kdd6
cQF9++u/wqLfLZGOSdJ8n1smiyXBRyuoGQGldpQdxCIAXGOMTMuOLMNd8fcFL3fh
9BPPlM1jviPUVgIK5lJN+dDAuD5IhgEGo2CrzAhTnhlYWLSqU08Jz3ArqoQ5Jp3a
0r7uNiEcgoq1WvAjxAcDLE6IP3//2ZSJwzWiiHU9nR+Sf5Y0zZeT1700WgBmaJ7k
Ek0Gey4WV3QXaqRPDoNAydinsswBNggzN8cxgbMW+51kIJ+5eCf4BxXowa/Shzpv
wmfLaSRBCeXnmWOx1fZO8cdyw3K2F2+FDz5NOW3GZhbS6SXZHvZTCgxjZcjHkU5J
yEVeZJRPmXqihd/BQju10B153UH8VI4rViZAHtUAwE4HQv8GTf5ho3K79yiDqD8j
ozcD74yXrgfBhIGxZ2twPWB/GmDRhzbPTRpyFc1F4ZtDHmdoHNeiSDeqTqcN6WF4
eMbMC18bHSCHs0Wk98oLyliRBCre5M6zP7RMnkivdU4DgaeegGavmmtgOLCNvOdM
n++e/0F3bXsti18HtW4zFIYXbmZxqN/zS2z/8MnnyuHx9LAQ2xlZH2wsLnT5pA8K
CphSF09n96ur09H+J4hJ8liwGI9IzRRCTCOCOj30jWjuTzdNqKl5JJlTXXG0YVit
r9+a/W+bqE134d1F72lA7Xx5WGyXverqL2blr1rvHIDb/f+33j5vyjD1NQXezTHZ
n/GLZKRIfU7TpJhCeBhrveQIc40te1keFKYEzGUewcE42Wc1a+B1W92NlokS0Rxv
vkxO61GO6uvzFNU6NMoOzr7pB5CzMli++vJ8ikYSkvpu+eL/k/OoPkFs8GqgPRBT
VC4s30AtcpyfsfAGzWJqpPrvnZVP104vYJ+tci62kNWQFSfdZY1mX0auVPdbGwok
KZy+P+61jXQjsuhZkI29JqeZn6niab/NN3Bv0S5QpwKa3lPaxHDjZqopYTm+1kMD
iifgQ2WpIsa8ktnxbYoNtwuEOp1yGV+R561vrLT0S8Ap2Vr/B6y2IB9CHgza30G1
HQE7KbI5mz4s/DFgqvlQcKhAkHdf3O+iUniHIYXhxcEz9k+Uk6wUnDni79DT7BAL
l+UyBcFNuepe0RQuh92msySYAimmL0da/IUnXlpMQnHF7TmrU10wwIHXXjgBBGeB
TLHujX5PfzLc2dWDjSA0Xaumv18qhG6fCtZnWSQJUT36NY/yoxtpuN+wKf/hpAhT
z7KbkISEDnXWt4k+FttHd8olgqGSjC61448bzHt2D1okAKptzQE8HrDbDEcESZbi
S5k7zQWEToRkjLp93pOqR5BRIlUcH8WTWIECXD9eYPgSMyqtXBt4Lk0odd0Q6ykA
Qat9pVi81GKt9Z0dkhBp+bCAgbkBTGC+o6biVvxHNsOziJ7321ItTm1sQWLjuQRm
/m6VQIE3UiHLHyxWqZei6B+ueWxM26Iowtdrnmzmg61A+nsO/i/G8MvOkZfo48J0
CUZ73avKJehy7CU5lOJ1kWNRacrXioww4YkqJoI6TiP91jde1bsroNW0gx1HmpN9
sXjIrwa5kBhcqcozmsSrnJpFRnp+7U9p29JszNGoCXnXY8QmT/XjIXQJLv+ETzPx
WDDrIirfGU2l7+MVIhZdrpaEGLllorfQjsxhST+7ltXVj/pYwIXEPwadShbH5RoT
+3imxDWUQjrZegBSDic0SQmLKHg8ZaUG9b1dCU0o1IqzcOVF3aOKHagEpgzK/VyE
FLaJNsgDoo0reSyiimm1/VVyg6/cf6E+59Wtq2UvQRPEg+k2gXMP0msUWWz8mRZH
HxcvBbineBb47+VnPI00q4TJLFxFKXzUCxDPR5Emf6ZV8sgDLBR9ya1Iw5O6wS2k
qfDhrPnG2N2MgTXInVijy4o2Tvc2YkjriB2qvi6GmodtyiUqUIVezSofDoaxQT1Y
8B5SHEkjsFijrlor5HZxNAqFZtk5+M1SFB+xNsdr88LPQd4pnteVT2fg7HQM63wl
92icfd/rk7hpzuCR4dwKw8eyjGPvxMEVuD1w1Piah5P0eulIr5G1V9ZupBTsMIwe
UzDSglnIL4Aeh0v1LbPaeuYyoWAse+RpEDB/LZVi4ZYBezAEY3qey0sR2mpK/TJ0
exNXLjt3ZN/c4mI7h29RUgNio6ACKK2z7hZtTM/9IzAz7Xq8OwJuRUAANey/vCTd
QfNbgCGpOhuiFwoMpcY7bxddd77HDc/BxAZ496xADuLtSoQhP1514gcnugga+Cag
xV8AXDv18ti2LdUxHEBvUh+sBYyMEaI+JpIZZXal0G+8frxd0fr6YrxWDKu54dc9
XJwtmAXsNDbs71s1pGRsFxqD5X3zjdW8iKLeOKrVOog+UkgrjGAPfIvLag5molAT
8WymW3ItiHl8+8SKykRM8Tx+l6DH/HX0ll3+hIVGvO3hkB/1oMzHog5durzhzf9Q
SyHQtUUNR/r2JW5GeJqBlHxXZF7DZh4cKehOWGF/APDhwqyl7/57wT/DDvz3r3jN
XGWF6yyxpJNiT5TG4yE7yK5+ohdb416EhlAvDZ75VJtAlrU69gtXz4F4CbF3kW8a
DjV9ILOFHQ0t/l7578+ePR0VtM5DwCR9eiZCh8DkCrGo3uqpTA3ELpHbRRA/urOb
/8VpWoOujGV1jcAQKKB/EDxEkAj+fY/TgD2doqk8GSz23IfSLYu13EOtVXheAPeu
bL3jCkubbm8etNQNE1VOGo0Rvh8v7r76OVuM0Nn+JIcaK+wM2y76/ARC62XG27Ql
XvOJGedXSTkXcw8Mkfh6FhBqSb5Xtt9MEdF7MirWMQqqxA7VpkAmUws1WRlgLJOk
ZKpP+3gY5CBukJTUDMHp+FVvvzeOvSrNnwDH06LVcJy5sGscbAUrNgZoCfM0qTmE
qPidfXPFO/gwNhik+xbOgMmYDZeNhZSUdfSa6E3i0OoMw6I6wcxa5q5lscVqkxf4
Rwso+6Ig4fsLQsGsIJ0hTia+N1xcf6B1Gu0/yEg72/+D6zOElop9K91q9sARBD8a
kxyIDGoXgIolniQobV2KrTS3Q+BrVjuDDbn1PAd9NidcSebGl18Q6weYq+5mXxwD
QBOY61y8yz7o+wFtsmQkFaYPPSg04VaA5v1PTi7g3ygUbJsjXg2Vw7tSBLmfxDOa
w2wkKE6nekVWSUp0bNTOZM702LfYOULO2bZTSKSDN0JH/Yubb0pA+gcSAUYou+wF
5k69n2VojoMQIuoFGQyCBI8wAwdbscnyYLJNtERFOwCmfrMSmuYBXqsHYLtfjydQ
nbpx3yf8ToRbR3MCI5LnjbRAtkCS9Ivts/GE5fIekPwpywomCjXzOXvw34JhJngJ
aZzbs6DCFRZrYqMNN3e874HoisPOMY+gEeAEC7TwW9jOxx+D4/bbX6Tw82f/oEbR
r+B4HTRy5ag7HwDDoOWwM5+ClVeWSD517iRFv9aP5OFmq+1JROoV8FZ3Bo27YPo3
qJrHUhAJrlAxCK6fBwnhL8ljeI+uTMe45S5lyAja6D7PkJx4ozAQHhhF90FozIEe
a8h2ULsE5jOc698BUhJ1N4gM9snOM7LO43X5l1nYMtCw77ybnBI/A1FEIoFuvmqa
cjzb0YXRfwBYBfmM2mvUas/++tcjTtCi/8Mtep5WE+72qWTEh0QW9PQXKnP7Y5Gj
pl5b6/2anlCHbFUlWk3KCKCYR8QOQOQNpPkTkT3omQcWk4h6JY/nX8sJk9HDcto3
2srd6xDwiAt+qVET4cvbemVjGzzSHh7QvusAcuQL+PCNRNbq0t7oIBrUrwAw1B9c
hMQxb4xGSebid34D1PnQXbh4JFVF/YFrDxdleEDSp/wWVIL4h8E0NpVca/sCFsc0
KofcT5FcGiBd0J7dG82s09DON9kdXwEhx6quwLupIxE1LNRw+4BpSjm3Q4lUaO7T
BRmBaE+X791AzVO11wtmyd8ZHuMwBujvg8kaFabkE8fEixHdw5uQuyObUTKV7dU3
KJ/VauVy0TgHg0bps3G/MA0XGvViAuGmm1vUrCSthm90ABt7+l2JHmrDir8w1Lxa
WHqRsJvdc+RfHQfiizpo9sbR4YxiowIqaGIbrO7EdKAMZGnbM0RHwctUYEw2PeYP
jZwSZGugBKCGlRyKxKPjpDOjAZvHFQPJdaMNO/bIHIznbiAYwCx5d1UfwMwGp/0n
aJ1YDYHoELFPAv/k7AyoUqk2MdNdmiK5H4sP7rVWRaeBug3V1k7I8Y26oSjCN3Ka
CyEzig3SkKQXiFdqCiHLffxi6L6wjEZX1IZY0CrSJyrYNCIIAVaJYK24KzwF4NVH
/dIL48Nq3TIpeQIYQ3bzBYAH80qIReT7Xs3V0DpRQbH4+Wfw4fj6NNz53E+eXtPT
cJxHvQu0Ed0NqEOggmRwLvFKe9K/RbgaXH16jcy/DeS1PEmIp3zJeZgwaXTD1tud
bO851AUm1GIYzT3rOTyI3i3fYlXwsvudhMbgwT4GzMDpVDbGopFdTZT/MjmocOJS
k8zvJcFJWpUx2KJmaRmqHB3Nu25fJJ6EqtyOwb7zo6oIDgoRUVO6/bzSJlXfH/3F
qXNu0aYVl1FkDgKAT+2NRTQl8vv/NFvnAZrVj5G9QTpeQBapYm/XV09UwxmITyuy
aBqROxz4hQcp9AzXJhGqbyFPmJ5IY1oLHS0UuXvnWgRb5cLvbgxZPnmKAnmWXH7C
HlyerjpCaLA3BvfWqU6XJxivH5oQPhovF1RuoBaubPxRTf42aJEgCpIaFy1NvrE4
ImomjdxfqSxi4/xjxkp9f51IOipzTXpc0T9vQGx3madibQa7XEY1xOLXQWK/NPDW
gGyst8BZLZOptzfAtMcV1cHHxkbE//3xBDNFXeo4jH5IAz4tfoGWB3wsSSHVyiVW
eFQ6aO7p1f0Uy6ZTQ8HNT6l2C00rwgOk9pKTwO5BYk5izUBMz0K9GVACGZm8zqGY
wQ9O3P8qV88LxJObxmA0Cq6LUJCYYnEQ5W3ycq3ZQ2p2VJUPPH3hH4ig8Dbw7Ocd
XKXVpn7avyS1/z/e/exONYNuBMF9RX3yY5EWdrCYpNHB5SMMGS+3hvNh6m4hjk8x
nqfSSxxOAzI9sukrXvITDvq/IIh/1uE0NXYIWU52VkNrsSuOd+66/5+7ohgMm6+8
UGpiFyikz+OWEbxEMSKRTMW1iHLODBpjoj7j4mJJ97u7ujH4iJOp2b6o6xvJDBJr
xnvIoN6fHbmvtFF6phhgu4Q9Sbog9kty2PdSPPiCV0Vlijr0z+kRFV/VjfAbZWkD
gt8oqIcldT0NHYM7EDqblFVQI7nOLYEg621VAVHilTVjjscevAhPFUmCnohjFtk6
hdxFyirUH0DNUzCtkMVAojPxv9Z/GcR6xzCgcWSJHbB3/R/Juk5yZq8Sdd4/0423
ZO4SnDSjX4TGmI4r3fEukFE1en0G2u6t1BsNLJLfCNNzozrMtl//R+KfwkbL/VFA
X2JuIXA/wwWjmKWeSIaT0h/krMEwZ3sRFhN30kcIEnbS2r0gwv1XsR/JsQhwfcc0
8JVnWzwqoSiJ7ce1qVDk7oa5l1ZN7XIubGm0spQZEFFamcu1yrZYN/XtnuXZqNOb
VMKXhpvwBqSnqear6rbqYtJ7oMYLSirgdULAP4TMA7g3GOPtyaMBqn3bb//Wz9V7
OdFGjLS+ArZvDA2s9zq+KcQ/maClQT+N3gqNR4eRhKBuGcK+IOCjFvEiLV4XUWOg
5DMmFA5j6U1cWziDBLuFZVGcqRcmSwOOSs3uukUaz8koK7Up8vrnTjI3OCx246sf
8mEpok9z9MODDT0tKhawW13aurmkK0qzGoeD+lhbn5KrSxWeFnRsB2g33f8i1wIh
26qaFy9R9e9SVn7yfscJBAuNtZJQia1vm7EZjvS86ucU5hTt66bvNvbGvduLDjNM
92BjxnbKiX76R2s2zx8Qc2jUwg66gMs9XaaCui7XRBzHDjrJG7EiWveRHCWvfaMk
O56QT2RO2qqYINFn4v1xxWcJFQTAHzlNbjYG71PKC2JpLB/tuDcdexe74OXx+A88
qt9HiKS4FRNmjKNmbg5arlQCirL4m80X9P2+KtVq08HZDHL/ubC+0QnAgcRurY9L
XlsW2FMY67+ylZHrsKHwfJewMPS27dBDT1Ib7N+as/mh8GiQIQRlYrq2zz2WntZp
W1uakPjk4zsF+mQx8sBPlKl6+f4382mGGLzq2UgB6f5AuVyoGVv2qcxVXxIpmoYb
EBUlroPfk0EedfmX7BqdeG/gCMxqj8w1KhOI4Y93xsjjKY+g3njKxSIIebbkekT+
9ZTkOM9EUaYebsGSOUU22QGhZUfV0BhKnobA1Ez36Gh6LZf9qCwbw+5VElYJBtAd
Lspv1aN14jqMDcPk8JbmSo+d0fjHL6+Nv76fR76RFvdrwu+sbgLCIOLd5V3M5Rkq
wyvamwfaE+oBBf4i3O90NJZJp5xsbAn9mGBZF2HpTGgCxFInI4o7ShjhJIPLeQej
JxeezY3KnZV8XtPRtTvb2oesYEBWJaWMRdWT+6Txx1SnguyObTveGG1kEI3omLuK
RL2x5HV0yGOoCieQEOePemUtmyegg2CvfapHuddFNpUQC3cq9u0611P+CqG9xPG0
6stXelSytpRfN4cm2+j/5cgx1tDOr6wJiF9+MyYgpL6MtSopHksRsp9qWdgrN5qL
zKd1nOcj9KD0mDyxJoeyfIoDzN8E3zjeIKcXEBtlvaoc0XywEEd6ykcJgaiioaUK
BipFMU19fhgLuDV00gCatwtiWuA+D5t2HepXX6grqHTfW8THbelXyoC2pLQrn+fB
art/xVjFm123JdE3DSvkAyo2GnCkina0WZtuzZfHM543VsZAe7OzECNRKW2hHKdZ
YHr8WNhQSYu/p0+ge2uuMCdULzIaOX3DmW9k4ztLyUmqOBuniVQt3in5ywWHdY1c
q37kY0hvK7EmnepQBlmAo/LLgw27XGffeeWUuE/XhCPpIigq2tzqCRXvfn2jagA4
7VwN4Duhsp8S/8YNzBEQlGX6yQ0CfXyJ4il7GiPWG+dueOTa6e5a+rirF1uQMHiC
vc2btNLmSoeZ2QsWr9SXzfS54nCbpUp0svsWo1yox1AOIwgv93gDXsHgdzuHdEnw
zKaOSkDza4RDCo5uKgwLYexwLCTNoMGa7dAwe5hpSVr0HJrjQ1wPmIf26kktmLGa
O/0NuDjtuEjH+JG+pMIkM+XhYFkmSN/UXmf56aD38G9RcIShzMrKMznQ2hqwBFEH
8QIh2PcEbYWC6DBW21QhVPsxIYm/v1OvXPUEOljwrNgQDGIFzG1S/ScheDYivcfN
n6ERj6cm8Bm5imDJRReDn4GnrXFuPxGqUKhXPc+bYpVNxPHqVEDo/M/sJoOs7ZD5
Y4+cvm8yOGHXk0gP8GMVtW7Pwx7mpd40RHfQjHA5EzZf3eICxfKJA7UKEWql1yo+
b+GsA6Mb5fX3xeJzmQFWoTv2VxTphrzufWkcKwRV6ucjp8Mv3Qc4qizBlEFHq0CE
ULQ9ZR57uM7QSOe77PJMUoLsN+f1x9ODQ5gVhBf1qCZsdwdWUjSZbOufk1K5oyKr
mSM2pFVl3KtKCdj9diws4fkDCaGj/I5S71EW6npNY9n9hTC4DJAO6diYiolqm+Xh
ko53qASt98h3hKw95TrOIJM9m1gLvD+SUAVKxUeO2xKvoYMZkNCw8mD5jO3VhaRB
nQUmbyLOmpB42ttx3awV5Ym8P3PeUJJYH9U9zZUU43+UVI5qEs/6VbBsbuiJ6O+3
irkaHoP6dh2Nba9e6synLgwwc1DKioMjNxMQSJZWI2jCrGMqoHTuwtTf7ku8DujN
1ZeL+Z6Rim9zZ+VJwg3X2L4eznMg3IWoa1JqV9FRZ849UPVzlFZUQ7NS5Hla4YwP
P45INdbwDIl6WOOOzVtwPHBAwllkaVo3k5txg/zu372PZmjYyn0TcMA2+y1B7dXy
n4AglZArM6STVGBaxIFEX+iGJxQjGCdn/bbzFXElquwfbvFRWXFNAbuo8o9Z2KMu
OwMic2rQEmiumcPXqqNp5KTL79pdNEj3BW0/mL1/bJooVTA7T6QD1hsFRkLtYSqQ
w9w1M3Pa7D6hDU0WHy2paJxXgnMJrg6w3w8LlvZlSzzYZThlr1e0y/KUmbSyaAoE
rethCPHC27X2WVMenuePSs3m5Pb7PeHZtv0xF4MXnWa6GgOvCypnnddcrFodmYyg
/EiJnwCqmU9qLEntUZx6zAbSnzBPxSyhO+f2qBDQnVM8gFLem9NIz6E8S+gmZDQz
y4A/NRphPiFmJT6noUgh8BAbfpQ1g0ZJiFJxDf/kKo2KywZoDBw7vUUnyrPCNgnt
+La99LnwZSdndDGwof+LlZyb+vTPV1uOCx+/pZksWvSSJSknHM9B2CkNhJoQrPWp
BCjChfOIHzNSjAzHsvFqqx9WwHXNqzd07YZnMYTVEhY4NzeKqfy9toXm/Sw4S3Oi
+TAKoAzb6nifzxav90DfjS1MBIBBZ1eN8oTJIFsoqtmPX11h6T/PJB1okdopocBH
6BDGzFcfutCfp7RhIRsng4AoqmrjsSaW2lxYSmXbUZT4d4DAYF29g7L60ZfTGJMa
lxxJf7Uq4zMVUW9ur/BCC9zI1odbn1SPV0gXWYYndZSsGC9ipP/hajgPVeSd5HdH
5BknYB2MWo9d7pUjKSU8rTY9iojYmn9bo56gKzai8ZGOTMbRnWh7oTo3Cke719tU
0lxHAZ39BaP4rPNjWQrS7J6OtRSjozszLnqr/2LQq7HHrOnWp4um3noL0FImMcJz
HcAZ7Yxfighwx/b8U2SZwzNr1UPkqIO/8zmxses9j45BuURkv0BCCGgx4n+wU8Ww
fWJVXkJHr08Kmzff/DZDUho39pg6wv9HCNkmInyxvcm2CcGpnJ7GvXWPWnnPcY81
zJirA4HrBWHYRgJKCoJsQbuZv9ykvfvFR9P48ZvPd/3sTaiNzs3wdPxf5cxL6dpr
mZcaE8FVEQi/6LcKAFGPSpU95ioH7YUx9JkAVDjlnJJ38qoDFobt/ACGDP+NhTDr
vTwu8F7dmPtB3ztIC5vPfLSABPPhlyRcZcRtlrFQEE59Myzj3ilANnInDaY9g64F
/c1Tq8WwED+Jghu6ZSTv7Dr1japli2vchyvgkl6P7GYFC9io00TuE1pNthl0t/c8
4prPVL9R8/mW1EdVOYzqIIUGmN5BP5P+EIAP+G00Rz4IHchubPxvilMoLEPKYiMP
Ril6BvIDTp7DFJ1ivNuyPT9s88WczfV9/S5I+rkcqCQmbZdVPNCoSzrhmhW6ViQB
O2MhJl5G+mhCe2sIFB/kzYayS2kjhXv69jOsCYa/wsimHk4ndCh/cvdN8UIKSxkL
2o/1YmR/X7MpEm4H4mNrefIPfUwreiMID8UB5K0scZkLdaDriZM7JSkCPdzMUv98
hhgpXmGKfzg8sz4j5wpHH+pPFGMzu7PIKJlmJAjXrukoE3LiW2UqLZnYdE2D3mDo
lfdnNfL57uwYAl98NzG9EmP/z8tTeOjkgyd4xGvGnAIqoMU9KqvTWxbEEXWgsn9b
AcDjoZn7jYo5jDq/Emujy3vxVCJ1jGQpbGqjB3e5Lf0U7+JruMPaI5Dk9VMasO6j
CswDrvzgdfDQg/Ygk6iZne5bYY7u6K7tuwOEhm7GcJi8GxLqnoN4jNNc58E0AxmQ
NZoF0N1e3r9+bCl4S7sncusCbL7xZ3AuaKgqcvZHDSWdACGB49mnQbDdrLPWyMJH
DOaU2/+NrvTXOQYmGmHFAM8Q4e/zFxJhPCTiPWhHqJtWss/jZuA1IX3YOTGGN5dW
OeHi4l4LE3wOExVqHtPmnWh8gUjBgWW1wGqhd3drAIRctC0i/qZl6HNyKuGSYizU
A1nnehTp7F9IJn2KCZ6srULmtnXCVTpzFeJ2Au4/f+G3UKuErqBq0He+vqGKozSP
6nuUA9W0hl7lTYWYljsDIFK4T5a0dKsZ8jC48nvRFhzfGKEEezI8rtXnL43A6EUu
rQbxixzGfKl8ZkzYMt7J7+yHVZQrqvAZcqsmgfyAjpnO14ecfi4M0YFD9nPZW59c
P/B0UmE1mFlBvnJvrNPDDCeUb3EDioLoU3nAvJO2mP+zHeF2kTJYVkR/RJ0TzYNa
Kfonp1uoh2P9wDFSDkpKtxtwqoODpE+kXHUppSzDNSm3OwazIa+pbiaMSrE/7k0y
gofCs7iRSCHl0oXfKR+Cdqs14A4X/ZTiS2d7Ynwt7xCN3cyvpisgnia1d+p437bJ
ycGUwG6fhkKtyn9m05B04dYtCE/WuHv+kKPhGKIyZO11R7npj/SZCpBIubUGTDQd
STP0pnf7YmoxEipc4Pat00q6sNKX0OblruQnDEYyRxyWaY02U6vByyA41B2WUqe8
KY1k0Uyoo/g47FWJC43Ke3dr5fCEH9dqeRX1OFc4Nrat8tOYGusrhbCmixvS7IqO
wBDKQzNQe+wR5GuMtFJA3SZdhjVUil99ZiBR6jaxoH7Lqfw3akIRxlBMSkpHtYtI
JRdkiY2JlspkRVeCfJLdAwgHKgdrYMq9CcDJEqYd604BtzO0qldY1nqIdliCuuPG
nbhA0TLJSWABzSl4yPZjK2HCP3pGFDcGPDvGTqImhmiTsmC7gjvtWONDKa+gmsLL
2Wm4dxrS5lxJLTWNPR6H5MRPC0v37vDRicscHGt/GWHssgOfennAsYA/imlnKTke
WuvGlzsCl2REKVaHZUjWIIJkS1ZSTXMFlQELtPfQJfiCioAbiLIeQsDcHmi21Zqf
fuk4+7U/t8IeL2LyUfWPUMzyvT8fvU9A7WRHQ67aG0hI2PmtOQinKJJbfNhXCBjN
AYJQJS6eCX0ZTifEyQzZ/f+kDGGcWZcMpPSqVbYtTzPPqGzan2y4jIDZczNmNfkZ
YU9nbeBbOjZHPRpTMQafNQlHxS7GC1HPH3wPOIZAmNZ4OGBKu9BEAAdG/qArF5ra
uNQhEIl1cMveIsUsAWvqjgOu06e0hIiHznbddIx7zVrp0FwBVZSSo9VzJSSzmQ12
z6xMc9XHb66Zm4SBfivv4EO8vs/tsewu+buTjIQ5rWf7fAl4D+InCwXoLswNX/44
KW0ed6DlXWCTig0MwulSyk/nbHGlb5HypU2oXOSJZuwEb0W2jUsFrxs88X/ie+ir
9Y5j0E/sJpgdIrKq5BEG44swR4d/HZxrq5E7PHuzmjv20rXa7MQVTi6hFBOeRVCK
8w7AaxfEK60ROXmi/0qmYXzhvAXSsJlKUR6At92+6by669ZhapqIURUc03OnILKc
M5HZHS+DuumyCdoBNUqt2v/YNnLM/MJNgjqlTlZETFMFBJIg8aYt8GoqXOY6edb5
3r5WUeFF7jkBa3HzLiSHSauz4S4JhlTAqlLvXsY032cIkNkz3rIR/WiBI2wufzWy
NIP+kPaoFMVgXTrkNxoRO7N4fDEX7IueJMNNQqVxLxKyZ6BbFVpPJQnyk+o28EUt
VWVI/2XhgXjVRlL3ds7PKhxAictic7jXLmCDXS8OUDjuQlQlL5w1aqbjvnMw59VR
s78YTgrHENoaC/BVjgwSSOnArcIMQQKfX2Y3mwx1Nb8ulGm8QTVUvS22PXGytp16
0e9+CskDMDUQWfokRCSfXdmqSH50uPNsT2cGkmpkB2yo19nC281vRXb4YfUNmvsl
iDoZ0meOLwY4JOjR8WNvhPG5tBMFTCAJiTAotc60h+6gkXHUjaSJW1CQhcn44QLd
X2dhTar3bFyHmeZ2+cb9niHh4eHK5CdzX06gHsIGN4zTI5RfiFUWhDnvcJP5Xd7i
6qNJiw7CRaA2C37i+SdgKX6kFxGIMhUdD3M3ZGEkIFdS5o1yf3ut04ExjbKBhGQ6
4bJNqUG0KCBWlSTklld6ljaaDAdu5SMfkw5lvJ7Bi+RI7gEcqTFpshAfktlzNkPC
5ZZlEb5TDGs2/NHP6BCcRLoS0dszf/NBFXau/rLviNG6pW67Vza0fIbq8/syOp9U
XAuNNc5whQdwjNE/qPTbfLHi8hCIhA/fThq7tnzH2YfsR7hl1iZw8NtdWRADCHBZ
wZ1rvZLtX9YwgVJTo/kx0f4+gDIPxBAv0Iao+qvyaoRUUS84NEk4Klbt4ORe3yAA
5PkYhamExOe7wsghLY88ZURtWVTfszbky89dgfC7WaYgcWJEKYQ/h64w4hshx03R
ZAAVHtgBwTnpBvXDYP5J+IjK5sT+Tz6KUYObdrIHEWz8Ya1tEKpvL+RS+x7glmWF
6fZRLDTZVQOJB4qfAQDzzRwA7t0a2NIfgsVIKNl6Io6svf9VHhbH2Wxan+c8pdNr
gGOzVWoW6B3OyYY45fuidk6yC+RnfjdcdFPfECCQsZEd6zt5VRVSwlfH1ktRrMYw
BHu6Xxki1QEpqOL5oyJpC5QtthFPsYO0uVlhFwu+3UJmpaTHT+elObtMhJAbKvwq
JzTBjqzHganITQUgfdvTbaIDGViWibSYk7SKs2H8993G4f0PloVgStlgzhAET00i
OQyOpcxT1zOTz1ivbCQXjO0X4+flipWwxtD1yey8RnIQNTfTyyJfaaObOrSGmQYd
Hyze2c3WL39js8fchWv/n+ADztnDBRoWkMgoDMhbtaYuMOupxJjm0I7Xc7ah31sH
BPATdnK9ozNRfSM5rcL5+dQ9JI9z/sQHmf/pAQh0t6iEmmHy5sKHrIMf3IRUxlXs
LHMlBbSOyitPwhlujUQufkBZOgPmWjm96sdYjf3DzQlmBWvnjtA8fi/bRICmlMFR
EaRliY9UW+KcoS+dl1u0GVus5zW2xmOCn6xvAMak2+ntWcWHFswMiIHID+Lgfb8f
ofi1DhS+1LffxP9DVDRhz1KbV6ovk2wxba3r5w+Uq5fdNxtTk7qRuIwxJuNSHCHf
vK2kZWcp/I3UoOnndQfR6Hk1x797GGEwLOocdxvLCLGA3+3GmwQTewtmzNIdK7tX
nlop5XzLzzYbjVXRAOG/DIvu3OzVtl5EK/5j4x8HhMGzg5ZZC1P5ycCCVRf7uvyw
uurioIpjKLZqtjPT5vYm+GUy6mOq9u1+FfD+35pXAVSR3l8HisykzbIU32xWhS4C
YC/o2O4DonERZGpePwR7hzhvu7tnDjA7a3eqJhYwaGHx4f9epTfT9AIhniIMWLMs
lIT4+1o08QXwdhfMNBuLmaOWKx5+gkztJ/WoNFlUcIEpq3Zv11NbHLML1ppZ9V1A
paDFlKi7vWQUkVpisqNdohDKvEAuMn7jwQ50cZrM6Fg3mho7As8U1CQhfJxqdHr6
8TN7Scl3nll8MAFZbT1cm/uQXMieAEZ6fpKKY4+80vzEpnk7c4HWaTr0SAxi4OlV
MsAPhQ/vYZGhxxu8Jz0nRenb+DMsckCluVUu9mV/8Q+WVPs16L8x2wqIC7uHXCFO
j/nTK/YdtnZVTLl6mzFUwPNX+bFVa48qAg2u5dmt7sOrz/lw43VnC57VqeznFxT1
hjVNBvei9u81HHiWAJiK40gGWP7EY7Ozjo8fqQchydX+pjpJyecTfL3kALgzPUOO
LI6goUG1AgkcSkKn7d9cJZsBJ+6gszHImBNK4gteaf9T1PpeBVsqLu6ESySWuTEf
5/ASszoto/gK7/ZwJxkxn+LeK07l5VQA03caavzyB/IiTSMj7Dpi14LdSIJ7XLtt
6iU32Z5dBoWwhBKmuohUYjmXuG1JZn5aWSChYuw4d0j9gVSeSRe2aQEk2IPALLCj
VW5Mxl5zrnqrIHWdS2tPsRJCV0xcCzzp72RRsXtEwEFDmEwuOr0cHMoAtonmtTaN
j+w/xG0f9wm4B5sMtk+VAcGRPc8RnGgFmCvw7eGIhV16ijMBzHjVRSDH1R3LFP/W
5LriYmx4ufvcox3wHipT1GAJ9a71sBm2oKVfBsuJZZOOA+1Wqn5C7SNFNELdm5aG
31Ime14UVEX+fgPzKBy+56VRtl7JkGj7MFFttRB06kkL1Qb7+D0Q+4CO8ovjYwKW
kvwe3yt611rehcWBkoseRvyV4rBXsoZPayT2y8OmrbBtmwfknTCcxuUwHIBpV31Z
pZLs39DgCCv7h5g4gfLw0ZSTXGezpK34Ws2FGSUBwuakQwsSrP8gW8qv1cXbZbWq
KbWkbAxQB0Xxov/djHl23zrlgAM7FMMT6fg3ydz2lB184B/6nw11RqSaxpjmMkFy
qNpHT5SNe1N9j/CAesrrFW/clWBbOZ1gXnb3oo1WZ3ms/FkpTafptN2NJrXaajAf
DghL15eCc+HRZKUj2tyMby/rEzot76PYq8EtrTTJm5hH5eXwnSAeB3gva3t3EYld
UCibYSrec/Iy1JJRSeUIgLsYetmwWUGfavNLLNfMJS400Tv4oJ/XI33DD3JyQE1a
BPENQLzGdd7BdDohuLiElX3iEjZi7EM67lVajxWRe8grybzPm1kCsZ7qiTQnw0fJ
2vWSWAaUDfs6QHkxbdVxGfv3y0tyMRC0Nm14ZBF3tETN/73L9sZC2S4e9ytf4/LU
lvS3IjVYCrhu6trCdiGq1n7DkWyXqN6PgqFsDpfCXzK+zw7VdvOTd0C/8KaXDyV1
E1Rls28u8XqrjijN8asxK/Fa2nz9HJapxH3Xh36PN6oRrRPtZR+8uEwrZAe8bytS
lP5+cv2CX5it0xf+uPaIr9PgPgTqS7f13Pm2BLiMagOE/gSPc4N9BytT66WZSmoW
lGaZEBh9OQY7zUvfRCZFeLT047seqbowVznTjRpOYNI9GE3AJOZ4RjT6BUA/IObK
zEdj6j0nKu60SSYzH7cJNSh+44HQv+jO0uuI255mwcpgx9cAoJvmPKVZJcSMqd+v
kSqXomCBY68qOnI9oAgkTFep4wDZDE68rLsZWdINw8U2bKo+qQ+M7BtZ4Mb9s1oa
X+xypWfMXoYF7hbDEDBlZe0Tx0XplWYp2kGY0AQI/wQHhqGheY4jxtw4sGS0yezh
nJ4wKWhbaSo1HxW62gTPVlCpkoUpKs99h5tUnzmYJnYgPY0OPFmv+O2EErh1VNHx
esMpoBpH14BHO4gLFboLT0XG3rO14QmRlWQZZj+oyGeA6h1Z/4E8YDoDRRlgbFkO
+bNBQZYXNsDDotdboUPPnxJ84IZmy1FFCP/wmiwvNM9ksqQ3QwnLbEdEPAhy3Yad
KrSpU1rUno/wANL0L9bAmaZvMIwaIPEwPg3f4wcVkTGVbhNcONs5X7cF8BjzwO6M
xOKvQaO2PsIucq5Xk9LFkQBTc+KNN5OqOxC3t+0DvtUrpzCuJICrzARtR1vArd45
m035tB5JGzmBkRPLOFM5libv4gJJceMv9W9SMnbCgT8kgrVydhQWJcr0zQ/OFm/Y
wYd8++GE9uLbb/YJDEUOsPdl60vQ2OytP4lu9UVTFLE3cQCBVkxPZNheIN6J6Gm6
psi2jh6tuI7MjdgzOh9uvXcIIqr0HS8SrIER6UMl4k2JPh1QxTRoOUKiZ+MEs5vM
+sp8HMq4Ff9y/Onze/7puovdo2vsxUqPxvNF/P21jsUFlljo08CnJQmiq2x67bpF
BcvQG9X0Z2RupKzBypcUvct4raUT8Of14DG8cNWx+LlaIY1WHii8XjHiXYCBnFBF
LFH3XP2T4v+6lVkUY8jx9lwMDWDW55K+PgWf3SKdzSfwTpRRxzcqsrE2K0h7wJOq
MCzLJClyy5rthDzCdKsS3wiR6TnD2O5VHjC7+ZHheKTMxPMk03Fhiq0RU852g5WV
oXcsAEoDKj3m2AJhNFaURVruQ3SMP9QmbDF5LxBJgfwisyhfdur2ZnL1p3iB8tdt
ExYGjJ29uWSxMaRX4IHAgrkHcff4OPS04bvgjAlms8rWOCNZeA1Cjs2CowsxpSlH
1hJiL7gf7NBPD5UoVMYprO8L6v2tmD6r7s6+8e7jUXDfYYBhK8Rq67QFY0Isw6oA
MmqK7eW8CcwWJwBIWB9++t+RI8b+tXPAtbZqzRyP4r/ByPhBXScNXYCorwoGLg49
fHxXDbJDFYK1nXhXnkEVhi5xpo3gIPUvWIMcK+skjVkRrULRGe2q1bvjvOz3P2Tn
NtwZG3Ls10H5iLljZ3DLbaoi4oB6GwfQu/OeDL2oR1iPRI+gFL/32InjHth1QeEY
XpCQlFEy/H0MgzwjHZ0fGfFWbd7iWXQG5BAdhwfcyPs+X+nyt91/nV6dLzv1aVyg
Yi3MUVzVMf0GGJFlncq8wcvN9x4FacZCFd1meMHtfD9H4mwPlksji1YE07tMDr0q
WiO5Xp5iOz2i13z9JhxLsXcnynh4pIQXSf21aGX5YoGqNvMNYyAZFO3kExgRM7L5
azeg8bvYFT7yYRrPVACMohvIHmg0gpqBVhNZHYUGtuWNASg2WXGL1ZQmDUqe4YAO
DTUCno6vuyQuHNaAvgwlHBzQwbvKNm/01SklNerxFOhtxDuNb0hGwIdbPyC9vyL6
Uxw7RSXmOt/8aYp2C6tmw/ZAbXIJ17paaKKyPq2TTt4++0G/FLLZIAWkCZMwXMMb
arjde340YQiR8Pb+Eo2t7jGnq+lZEyQE7uT+tnpBeiLXY6TRRj2lGK7k2SeC0RGn
tpyf5riQG3P/0376TjlzWhG8VghNvyZiXUuKSkTPW/mVSgNdZ+9CZb1JIIUuCpif
kzIq9sz04y6nsgOjdjXGu6Dt3p00EbnnXfvcZFQOcziIvcmL0MjtR/Q49tplmWQf
mwHdnUv1o2JwUQ3oKW4HJ+UGaXbTdBn+zmmNIrLxtro8eRCTHLV5K12I+5YxIUBG
lk49NhdXs/TdneVFJXMPN1Vmu8eaKx/nF1Tiyt84/Q4IlTgGOnkMOzU65dn899+x
PPBVRrFz9YLfDw53XdYPSiVrJiZqUOTEXFclX/9Zv4cS8bd9bi152yi6F2Ir2UFF
KWZgslQSzoaIJhXDMKRtdi54yTOrJMADgb7j2RWM0Lk5wnICQ3RSsi/5BmHfPCTB
Fsi1pF3DAd8VSn8IKZflHcNOxEb46tVpMukU8EP7O8XhMQyW2ZqksMDu2FvLZhZ2
Y94yxN3ylxClE89Sle2fjBPsB8oZ//bCv7O9MVp3vLpxlGpGV3kRkiDxtHKESdKj
Gwkr0bsVRW7FNWyBrZbPRQeb9p9m4RFQOBzfLkfhWCNMk+YHGTVbQiGHArY/evcn
HpALBkTNDAwmbXEJRzuw8Qclxyb0ZoODPnu9AhA70361AD0wulMXIhegRq4H/s27
TSkpDWVoTJSN5adg4wDNc+8TTfmngeor/H2dqzCgQz56iN7JzaSeezPsnqhgEqaz
6qiBvWPvXfZZ6L8Hael2YqGfXGji55eMy9Gh505pLblsSur0bKjPjiyKmARou1qa
VP7j+akKMYKpkL3FZQ0VmGc2G1kHn/Rgh7/egom8fmW8tK9NVwYY8xcs3e/iEWjC
hRsNDXuwIroGkz5YI3fRR3TS8IPgj81ukbFkzk92h9IwiJOZZTiQJAJZTP2Rmj0T
b/MCcfCAgO6EcncxVBZKeRQ9UiJsi5nIqstJ0bNaM5n/KZGbqOp/50g2LJfxjBTh
ewTyIgyRJDqblZR7ZYMhPN36X6akAyOPK+X08MF07T6BSXxMHQT5pECnTuBftUJG
9C3Ba3GIA7e5j5am5qgMUKIw2Eqt8GkDKsFebAaFMG6cLdJ6vuaO4WzICmiizqZQ
AddkJgzBpeh80IvTTLZ3bvsUzHGGK5zvIuZ7hihCtJjooUMEsbTvcMNUFhPgE99/
pewY52LmTNTTt97BYG8wpgrQCxhDDsz2aHKWaZKQvMrHr6cxCembqA2OlPH2PmBE
1yF8hpQM4RwktAaHsXqsT5tbSHsDA6ESCKSgH6IdxIOAYHf341qbYBovUOHvZBOg
DIA/vRltYwi4lf0V+cGmbvBFGEzVO0apuFGO2v0TK5w8bIYjfCR4w5nfbDlIUxzL
SJhWb1a6KM9V3IkbJ4T3lyq1vrF4y/1a1ENgZbWqTwwRXjMSSPVItbovziIj8KxO
96Pv4mcQfTRqJ0Ih21aq/8GKd9NNq0WTu/SD1C26uqVo8NlgVASr9ALnzMEF4sy7
65Xcb5Tk1TjPmkyEgmcjt2kf9SVNZPPhiQToOleAOycF6jJelyRXqxMfiJ/RctBE
fedVOsbfqdWWNvz3UdJOusd8e0cK9yz2oqzZTK5KntQq8cqJiazKS1I5kRbqH/bp
59KRxOA99K23hfZOpJjC9M9qstPQo7A8sY+kZmC4x5vW1sP9UBgKstAqHFLWggII
UiQjNRYu5egvc73K7jRz5azcOVKxJeLqLBy6cCLLmJkOVX4T5P87pVOCGXr8f1nK
xO30SJMCInnQdHZStFweM/AyXJXM9H0t6redzkonLrBUI/rMvUnLT4ydjPeN3WHy
tfjY5bEVxpBoqzM/YAAfIohwsPq9ugcMo35Xz+9YvN39nTIOmR36F9vOtZhgOWSI
tNYaq5iid4klgCZSsNyiIg5gk1xxD+mq2NeHxYpTOBiGVhspp89BnNQu444Ws1zz
sat7UnLsJc6GTKtp9MhxdWQXrnqspohiRHSIpoXmJ40h1zX7JEXsV3BlTAphQSS7
bvk9mbICF9dUCi2i0/l83HEron9CY/6t2Ni8H3SWXeG+32TaJdG6n8idD+tETKUF
wmF0TAKzqCj2K3iWCOg7No5SoZgy+qZMpAITIudzSpleQHKVdjkqyjorCAbu0dS8
IPHzEPk/6lqwBafTzmzzWulUF39e/YQSoR0a5gCAfnO84u31fmfszengaZGvI0d8
v5bJw9AAO2rTLm5uAM4aEqS2aRMi3wFSx87pMppsQzSDikQpNP/sJb0MW+HACqKV
uhWK/xOhMcGwukx67wceZaqHInQPlOBL2t60tL1ukIIlp/5bvgR5vdSaXnDr0qSq
TMCx3cbbVWbPdqhcr5blqvjYs+uarV2jm0eia/uFavEcmSab9AmDMTIaTQKNKTfB
4pisG030Ii0WFjQ2cFak7bWC5Im6rUO7MRR6v92mX0I0C5RwsaT+CEdfP3+/z2Cq
7eoJ+wjdgtXNmZar2x2RnbNGYrBugzv90DhhCYnvDAJ2DZJj0n0ZmXSivLY/lXpt
BEzVF101GNkLFXMirE1FSK2vtJc4gPKKHkaUK+XgUzHHq1pBV1AcsB9zpylsTwYZ
AF/byKfnl/IFGg4x6Fr7zJ0tm5j19fbcwLjdRNKRyFNjt74epOmY7iVrHTjRmkym
fa6ysmQWRtTSBRoW5q/Pli9TVkdKB+72fV4cwLggrh+U435YlShPTKEuQEdz0/uo
P9CObbVUNypu//JX1UKhtnoXOUO+xKV8SBa9idWAjb9BNcpBz+spbkoa7GtdBGa6
OZl6foBLoNzN3EQFAMv5xqJpmZDjTK8RSV18b6UKGNwWIx3HULhkDo5jlUn6fzbE
VY4Z62u/xwsqFHFOTt5kSw0vQ8h1f4BtvdfoB9wrsDThVTGI1QyzANvZuqGx3NWk
6LYGXiMV4YSzPXvsI6MYC8SROs1lvP2rVaGXpq94KUx2RNLh6i0XTSKZLApujcJv
+mmomi5j7mb580sZS1xnxWRIDhTjWGzFkz6uam+A1A30uB1NdU0CUr/ubICR1GpU
dQFD5sPiTo4R0tb8kA5K41aOQsLoA/JSc66y5e2Ih1Rxf3/mkdrpJ0l2VD36W0ae
Pk4TIZ9be7Yf5sqmOhYOUvhlU4Qen05YMCwF0ZbogQvSeLfxJmkVFqJ3X8toNCVy
5R8yf/FugTpPu8kiHmTZXaYeL10iCymaYvf88TonnNFMjjmXP0yUalb8tK37q/7O
TFjyx1vz0RHxjIrstIhqta8OdgEk+UoFX3mUiJ3wLdqlcPwRMWALuGG9fp3hFotj
r7jiABZWFuCjQSC18xp19jz/042VxX/kpGjwG4pJEUQyfBp9XFl1YtzNanIzrO9b
2/raPI9KCqT9fknKxrhlrmoCEKCp2w9mBPvmOOT/OlK/gaHWtF3/nfBltsOjZtJI
AoPVPV2wfWvawJkuFGIg2QNANvHesPz+CIKr79MKKAWzok4bVXPG0LNLxWE7KQH0
zAsbYcCcxeOTRpKFwuW3Mc/SErZ3xkO928et3wNW+BYzHu+CgM3O4AbmKnjqnlsj
35sqv0OFEPibphV9V1qqjjqwXtGKqoKn4nKaWOj2Ob8oabYn7JOx9bP/ndIqePgk
yH7kmjNiVOhVJqXyeqZwGyNZf0I/xtVUPV4N1ml/jtlf6VNym8qmuC4G1t7Mj3PB
jmvKdP43i0wMM9Ub/yIl2RF/5KOgPl9Tp3kdJc+PJNQOQLS2FKb+NfWq0rYkkEhq
85JY3eSET+JU7edEuRZncrQs1/PkgI/fgYCVI80IScLn1ZzORicEfEiSDHhDP9oB
yp/OVJ/W32a6l2F+A3jRH0X8GHj2xN4ecUlGtiL4P0R9r3epiwMt1PTkmQlw59+6
9wIpSBiHnx+HqxnxtOFk792h92ee+7tYu8cqVWMh/ATzXn9fXWysJjJAEh1VUgbU
kBy9Ebqz6pFepuxl8eSefW1cYJ8crWTroB13cr1kNfypcoh7iQxVI618NLIgAZju
blcvzfH65nkhX1iXgqYIPSPq3RKjU9uPRrR3w9MaJSq56Td1YJw57D76Go7fCeOw
hwZoN0NXSllUbb9DqTS2a6DCnerPLug7JamWOySUEOxDXpPP55gCuO5zXqGr8/+g
Aw2Ocyn08/rADQrk8RNjw2tMIA9FFy2I7lFyeH2MTpSkiWm+F8L5fggnbgzCfpBE
HQcuAbJRP+wMi2RWSTVhkhWVOZwBA2Eo3C0jQLR0Aj/2G5uF9IOsWMl2aVvwHaYS
vgpKxxZ5ndRgluajAwPC53mx22XEV5c6uPrtWXBsHPk/YB4hyM6A7oqsk9Jxn/ct
kdAyioLv+z3G1Zn0LW6a7bJHm8tMzbntuMzYgeCHhD3WycLskMK7mh3JYMR/kz3/
/Q+6eU+rMNTEaLOoJxaHhvSI5hhx1OPlvmi/DhhUG4QJJctmSYZVnJXAv7kPeix2
JsCrJ6KNv5TfEJWFNvQdbXqF7IoAZ9NzJOFjC4v6XNybd60mNTX9RRubmaXPk4c8
fghDJ+0lLfhySW4DIQLb/CVBXRX58zwPqR+8nAIQtqHAnAuACltAGbMLLlfyqzPl
feJPdEGBrJTQIdoBMTmx1I0BRnGMWHrjXO6M/+M21c2JlJB58NZiYt4R+hsXYOZF
vYCs89dUxdNLEpuevy66EAauzM1nlImTfaIda/qcQ9XRb3K+/cCoorW2HPgpw29j
jWytABbBEVYJrPBBT7EZzlkM8avberPKlwdAiEnJgNstGH3T5U9ehJy12huvwerL
2L1/UbOoxIOGPifljvuYdhQoWAz+415ftxGBRCgW2YtuD4gvxYI9HmFHYW0v83bm
IbIC4fkedxwxOkU/VtaiQGk7Tm4pAeYLAdK+oWOKMXM8oisHTlT/LlA4GEU6slpC
otwp6jOrgKt2BasIUis8GBcf79kmZWDwZD9Pt2pOyBov/DsO4bG5G1VFVBwGnOmL
wf1IXJZm9mWwAn51/5SN04oR/wOek4cdQzLvGLlEYg0m2h33Pre7g5e5ZEBC2uC9
hCn0HfpzZYVWpA7fI9YVv+0Vb6pgMcTo3vMXwlw72D5tbC7J7TbxEdomtO36Sr7m
p7jlllCpyC7DvuGH2jONbxxWaOicpQcwuplRgmX2xBHhIXek3ZcfPSKfMahkhAV2
U4pIjX7BsYLVvtLa8ObnEC/a3JLOSo5WZaYxhgNlXN51U1MtYyxkxXcd9b7q7i18
m+pvf2uqeOyXT6NmcaO4SsXJoY8L+R+04IyIdOGsnn9DX7Cror8sYSP7DHbB8dY2
E7xxeYTL8A2ct5GOIsKqw/2WEwAu34wGXrJaKAiXCjAQUZZsr0gF6qKQi/hiqil1
6+IrNSGtzbF7PICtTa2O1DnGj6tBAF7Df8cvRZr+BXGF1+bVLznfGH3LVhIcTVV+
MJ0CWbHG/5k6Q2oStrWHhBGYbEUtdy61I7Z/+QHQVSjg64AXd58EJ85SCDB+e4OV
GxaJcFMAkOHGmhfIvDNk8Ph0uuOR+qSFLDmCtYgij4KAIX+hF7FGzTS9eES+Up+9
iYd/z1wSNPGvFwlm8bjOdV33QWdbr/zB2LuuaapVyJQS6mjBxZyjYpqvbfUcdSXd
Qk7d6zRN1Hkktg/xtOFjtz1uCKmAgMcu3giM47+XjwBZHBLT+6KwmbnaT43HBfXR
5OiWSFH+iYPXjgQMjl6ZPCJ7f15MZCCaqV9+qHTqQW0xDL9a7B3htQDtOm07mzsF
wAo2w/gI1qpF7BxqdaZKb1vD04gDHZf8YJaXcALZhGviCbKk0e5OKZ9gTH4KLJa5
j9ylv78KW0+SM6vOfvmz9b4cEd7PksCoBNRHqDQmGesUav9Do27hboRbyR+MZRcu
VcQ08sbU3sujO9crQ9UFymNev45PSpIq8GjoRXttNkNZNZwptCfolySLKcwWLOJ2
0Fa6OStFKUlIwtp7GuSVguLyE36u5e6r9hrf0xyG9zWDJ0VgjN4aXqnhXR8to4ES
4vYWuceoyEQz+Ky8gFX4Ek0FFKHIF/Ht4xf//5wzBBjvQzcaUsrsuqZbni4FpACk
iDCeGjyexfP8Esn402uI2+oDDrQ5/HVRQbv241P8/su3GT1lkxo9h+54RW2WdgPZ
esO8Jo2EGsyCrmIbkHnqab8pSfKzUwVwUlWwpTATP+s9fp7TGq2dPOKYHudE9T4f
Pdzlpn855F07zIVKsymgX4UM3cIOcJt5mrVXJrMLY6p172H94cLJKXszOyogBf8s
IyKg63TFjhMNjWnm+XryGF74kxMMU81oM18zGDRMOweWc2rBaGpIZlc9MCFbmqsg
FRURoIs5GUZ+6cBD3i32IIPfO+zsOetLdVdfzU//nl8TXKDXS4GKvoPE2sEt6jWy
CMbG56T0elQDjxWrwPYNG0fvoYH/EIPHoDgBpmdjfU2oUVpD7jE4JFxNOIF0LfkC
VeYhYIrN6oKWRqAH/PYQRDBMVal0kMBlmMiexLfhyflbdPWNiAEDgfK4kSrDWnIK
YtmURfHpl2w+YoN5ixCQ4HqTR4CRhZ2tHwX6D4L8sPvyAyys2n44A7qqYxzGyWAF
xv38LVe79260gSlNiJDr2YV0Jq02AfMEjdr15MEIkk51z3Sh5ycOWKODlX6SgYD6
df6CyOYGOKyDxGVWKRqPdjtwNq5NKhAYS9q5lREEA/0p8Dk/1TkDmpYO1gwLAd8d
KuGJjig46dQlAsYxvKkCZJKdTN/1ujDiHtUyYUrmCs3U9csrm1mK2/ztEz8ySqyp
0vHyWJzCfWJox5zGwQnDr2gdvwsHNpZRzZYUYZDKy3Pf8zH9GwXpSjIRXePHdgMh
5k/eauY9n3QZsZVgkzmvTiYBPGv0bHE07SVK3Iyf/MZQXlS7Rv6lPL23o5jAlghw
KvJ8qJJzm5TQQKppGTHcQJzetxg3+Ry5ATBk35nO4ZrexCPzmj34Ha0Gn5kCmkBA
QBxH63yd8TJihVex72QsCAlG/vfMiK7Ga8OOtmsN2GdsnktPirJvjesww1UU4RjA
A/NB8xp8VbzPBwJlL32DLR2IWTuZCIlD9c0f1zrg4kYPwvp9MDn4n8uF6bP3RPMm
UBFckQoRed0WAMVlZCAFueOpj2260vN/NoGohisOkgcYlX5Ry04a6WlzpoCrEu9J
mF60PY+SA0UgqgZbUGseLAz0dqo5C/exDTXuRF8l7THj/5S7Inajrkj9lZYYEWlj
tqI2Zy2lLFETv5QIaidS5cCQC1xDez1E2P+1a284OaH8HVL41v1bchalBomcYSnB
gg/1vRKb0GeOc/hXnOj/ZCsBRO6+F812DWMoDEL+0ym7c3gUDjEPeAFvQ0GzZB2+
yN2GD9EmnZfZNWgoanVkg8mbShJc4IzbSw30ZDtUQTBWb9WuNk5p5WCoxBfztL38
InQfykNZDKkDsSsTUrqBfut0hVbQ4R9BOsT64zCBHWmAXvw0s3Isic5h22xaVKwd
3KcGQLssML7Ja0m3zelVrK8JeEVYXFhdcmDpUlma4UV1PghRAruNRSZW4y2mjg8N
NU77m7PtFTeOd34tzPLra+gDoyumMV0qzuyyQarKLAXDiohuHkGr8d8TvCW4RwzL
zg/wpJCy2X1pGb7YC+BihPdBnap+sTQ0GOyZnp9HCWpiDPjgxUkxhSbyKShigHv7
o8QwoN0X0qc0s1XXlG7F1gBFqariCsRojPpm2oO6BhvgUeBbGt39uFuvb396Qv41
5XQGAypa24d9kVB2cMvaaa8pdrFTDvN6/E+ClDQYrrYx/BhdQrg0jc8JZbmZaVU6
e42ItgvZt9ba+nPwl45jfuPbGmNec6eXUft1Q0dARR50MZlJekC9Kednqc/awV/u
ZmLNKOsNeKdac+FhPPNX9auNWzXtAaOYl1fgRVkoS7rMFBQeD3YdjNb4tvx1oqI5
9LnhSwBpWcA2CoTeW6u8xw4zIwTu1MNN2p58Bf87JfzSFg8piOuaDIhx+iWeb/dG
vlZHp0FhEezrdvUxRlT5EEYolb1cxsM4hK4LxRpyShAfLtsAPDU1uDulMWTpsO+E
PwYfDqn/5XHR1ja6Snp98mBkgeerPqi6TSHLv4e+m4MHD9tskBY5gSRfG2WAtpiW
jB3bgDUINqEey/WmNqETXSCA474UK+Luvy5fCXJosDgv2GBbv73W5g91Rg7JMwx/
9C+PCyEy3G/ok0cxFV3kCSwqvFEp8nltcvENygfw7gG5dSJ/oNhWK3/aeJfizUzN
BpDhkt69ixxYAr8JwkecqLLCKDzR69HVTaScbPxn7mfw0R9/NtgATtiz+lO1xZcI
eDxwHsK/GHLk4VgK78Zj/5aMMhCfwjfBCpLmhM0B8ER13GuWc1IElckaNmnOqWam
ZceGdoKa1WZQblKuBmBmk8OJB/oBvoVdKqq3qOoEXDDYSdzj7PDJyRzrctJHgLXV
mA5LJx0GMXilKWVlmfdMhdlM9gxetPH/u7YP+q1HpfFXLhvjnwLj+L9/FOS9QymI
VP8/q1n1UeUjwTdEMAxnln/rYswdzu7uSWXPgxBjLi3w0k7QDL9dIRzvMI+77zqd
ByMXAV/cXH2cpkZYzfTpYwYGPxSrBbG9nCyV63Qm2UlszzMc8UGt6Av4VJzGf5HN
FJ7vDD/gntnvMEu7LgBADclbh2sPsA7tV2rIoMOtzlJQxhRYxnkaTq/0f4xMbGuW
VNo1fHbsmPaRCLAyFzZjQeMz9YsFjczIOZKC7K9kweIvefvb+ZbUKrXG8gha5hI9
r5wswKBBxI3eNiZqBoMXvH/5g9nX4DiAzHD6Aw5TdeRKmRBaWPlTuik72rZ1GBVt
BWwD7l1faJECdAxg7w5WqxsEMBL2eXSbku5Fv67nUdhqvwjWzO/k89ldfs2LfZYB
I9cqh4gg55wFPU1Sa9/T7rDAIXM5L0Lxm2GloB4uJCt8AbYmO/RFYkUIMHyqDJhl
9IjvtJwhsiaEXNjV48guWdTGqrb8HtBS1U8m59II7qriOyAxbnfXVk3YK8W8JJqP
0Xz+kC1xndvEnVqpqQ4gD+MmGB3k3JSauXQ1PpqYJQRDEO+Ivf14obLfYTHvioDL
o9TT/1ifMiHNNjHvOBJsC/w8WsgipmclzsF8VlVnMIgI4vRUIo2P3Uvr67i3gLMV
e++qu3edgbp3kIe4YVdXQj8pSByOGBUiB0YgiboXDN09p1ODeJL82aO/4GQfhdz3
NvBH7cwxgi62pCMejq4kisJpWE4Jfsz4UGUPT2QY5yJC9JjLSndCjJucmqyHqrwm
+cNVz9exNujoDy9qundyhSnaAk6oSBU0JHW1tu0BAltPa+vmq28hv8Dei/I//Fgx
BuECvV2MJ5C+7v+M9xqy6eNl3QuIGAikDljqGkYsnOarzSJOi0cjzFFCDpYDXWH5
wzTipld1gh5q4MSUUzzkx3r7rgaPYrJG284b/3QYzZdewEP3FACdXiQjNxoBj3Hl
caNIn6Cd8uA4v443bdhjdRYf841u2GB8jrx1t5pi/wN/z3tDhK3m1MTPLqpdKoeh
O5sgjGZ7gcyMl7FDMInMX1rOo/BDvKhELSZKKrzpelthQLrzxXdGkPGFKkv+gDfz
vbEmkrR4R4hfLrT5nZ7Md5IrP2msffP8Winis4sGuNezkOGxvBFx/X8NBM1GntP3
ezme9l0BP1dFS+sl4rNr/7njkfRC0C2WlPoaW/VHwUZQ3mIURYiZyP9QdrvLli8b
E4aYowvkjMDbVNNXaiH1MYbzHH9JR8a0yvL/wUsF2n93DpvUuoL8WLhHnY54jNFr
mv4pAwxgvM9RcNlpspmhM1go8czBbAu/AgOIfNYM9ZtPYiZlUhYs+PUzC1cXWDEc
rXATzQidGTmKdcSQxJqXvqh8OrngGy9RCoa5NMzsCaAHZHpAWENPjHBMZbsESs8w
Cak4C/mQvPOHvwJbeM9CebvqlXYMnyrljeoF+Pb/LBG1lOFmwEPBfTvxzEsxiDZI
EVmY8JnyG7WY5TRGjzx/sH6MDU18sXCbXJt692zQy0HDs98Gnq2YY+YIECjENzSZ
1ST4WT3RFzrRnWfTW+3oFYvCU3vL/gq6VtzHImXF1rFcvGSf8OIrHAJxT3D1L4tj
+f5alnmujM524bas6HAD+XUbdIE3JLHoZxpwN3eZV90kehPOeraKZXQsjH8zH5Gn
n0srgm27GXNP6ebdFgiTzDB3yVcxgjjVgQm50E32o2do3iOntX1tkiLyAZUr7d8K
qttU2Qr8KVOXhnb2BE7awS3CbWJJoFcfFeFxetHmk8tJyXmqsScD467eRFYvdHP3
mwc8u0/e3MFijjBG7npug4WAIswR5evsM/CYTrWcFoFdJwwByJSRVgaorX8yQI8M
xqW7+ciLb7EAFDj4rm5/V+8VTe0wLexMysjGRwyWU9GGsXWmax7T62aMqnJbB/6F
4QoazFwrlfJ6hD/4GHRRBTQJ3L+HcV26D8JZU3pD8vt59K1j+sdZbTcR1vnr9eim
bFrROHBQhrovc5t5JCcFhigVSSkEl0mlxmlhR/ioiq5ZUhok2lxB69gDeArv4JoL
c9TgJw12Cu9W2d+16P+Dt5uWwWJH1jTaL29sKehzHNANijujRgluReRQqv1Anrpl
SbXQruP/MN4r924RznCbae9MfOwAy+4zUsK4rKSmhYDDhsJYrw2wm4N9LGErUkYO
ykev5nJvrG0uD41YiQEa1Aq9j7U8rsCUJZlzdTaZr2HwYKcxG1WrpBfBDzQIbvUO
UVKzwaqwTe4IfdRg0i/FB8tETz525UHX9aRvLyn8rrIAZJt9i8xcGRhh6JLEYXIy
AKOnGCy7DN+Qq5IhXYSkGhtupnX1Fbf0aqZi++wE+1sUbV2VJwchw5kcIXoKP9rm
nOazZ2+4Xhka/bB1diIC9pTMH3M8UG+BiRm8LoSOWI6ntx4+PbbwsJZETOlTSlnB
tROxNtf7WpDwD5hqSM8Ks27bRjF4D3a+Ww858lnz4M9aLAhEoRtN3E+MyPxqHItV
FmWAhOoJ55cp2h/xhUPXmvY+DJScT3FQ64wX3A6msupG9pUxabfghA2rJuvdQMJc
hD4zfq5cBJH/eIawBGjcx0eVfD8ZvnChL1V566w4mw0/RUYihvm5BJ27ibFB/WR3
oAWbET1heNUGtZE3mrzCvI427H+bdtpj1EY8rh8s5C4nANx8A4X9V5VahAS50KKm
M32d/r5fiQXue9LTfMkUKuAHDX4N390MyeQCYzYEBmetczBFlLUAQ9IhtiESaMzZ
qsHKFk6rd7mke880z/3hCCOoRG92Y1BYA47BVWGOuZiYRwZ8JxM0nr18jTjalRAS
ksrRrpi4XqGZ2qOURfZTIrzxL2+q4eBwUvE7yqiOfEqwM5snn97sgHGKXrdqEnU0
+Ho4z4Yo7O8mBe5bXEwf84zjNEUuJnnaNT3vU/FyGoetGrJ90IbFGaLDKC5S76qd
NHilExst30CmAmZpUvW/RRzMoDfyEnZGaM+KAO9lIZfV6lWqUksbKRX3oWQJvJBT
Rvo29UVqJmp1kz3WsTbtSZeO78c0pEFhmOT3OIo4mnNzMtaDHB8LdhSD9B0DZjV1
GR9biTfFlhCYX0MVUl0bdCJebYX2HoV0UwQUpKVYg1sIuqaHj+9w2gKRzoPnibme
BYF3fDSd29B9BdLDQm3hyQsWFiSZj8NrnpZ5HF63b+wJ0Xp2sfGMNhqEdBa1rfKc
/oR/zlNMxxHcX6n0vkebLhRrUIznaQfNb5Sxq5XyA1Lg1JqboP0+vHIhzLd2gWUY
uOoI+XD4S2/WUrqzeoWWQTBLu0nUWa20QB/X/k2ef8z6qXTdjKR8CO9chZyzz5X1
u4XjSUAiCAb7qlf9UKwoj+FMYL6V29kRpSOyIvAOKkVf3DD4YruWYuUsO1EY2EU+
PxcfxNWvJa0NFLgJ0aTO50xWLxVZG5wFjAwic6POYQLutPSB9j4eMGDC5XrnOEWY
KtgLFlsAF/XKOLqEvZGYEIPPZ3rXj0jmv1KSAs4dDX+N8aBzjMxx1qZTeSiYSc8+
k9gjcc3VV+SII33zc7R2ZvQtxq2W+dNNwplirZFyGUxtC7hcTb0RX2BwDMqjw6eZ
QiABAZNyY4L1UFHdgFWBY3+HJ6/9K70aa5mU+KlyZnqSOFkJovpyMXiCH3S4TAAP
uYUdXDbsyooKD2vpn1gb5PvMtpuk6uBCjGwor9Gid67rmi+vLBNzssi9hgVKGrJl
H25zxuw3vo2sfZ8ZBaidqeJ+TCtdLGP95vHqCATaRjBew4y8G+vQvVuSPwfOolwL
4PCVVbY33sEy15Yp3xUKghFzlcOyavGchFpCsqhZMHE4Yrv1f817y1R7EkqVCWtP
5y6oIcrcB9KqL43URKHHvlOWAG91JEKSjphE6X0hylX56XyAPZf3Tu/wU67XS4S+
cU7198BuJ45ll1QUd3d6XOCo4tdOb2A05kQgzl0NMyGwUXRfX9r9B3+sVyyiuk6T
R/2+1N7vO91T5K1Ds8M2muh16ijY+YBkaMRkE9pm3T1ZMqYhr47j2x8n8SabLrWn
LPGDC2ntUtb7AvMALiYq0431OtFqBVEClt99UA4LW0bBrLrU8AY3y+K2TxLN0ko5
0dnjvubYR67sYAoOliQ9h7DrabETj1Hl7XO/cdw/og9jW6BscONH8XJ6+V70DM0v
mlWhx6RhJkgj/Xfq4WlGvqopfeP5mJKW1I5Sjziyr/pjE1l6IGK4IhcO1G197Riy
MRhuhdQZIpS28fuxEIIawPCUUVmt3UqthboBpVU9px8k87C7W36XpE8MHlBcH2AF
kx2X2So9lrYBDZ8eKfaJqD43w+tWr4w2I0Acysa2occZFA5wpLi6tPW4tgvRJo82
9sGebsLCfZHakZVWBmL5oy7SSK5lRfFTYj/YmvfNbqxtYwm0NG6lO2AqOADhpnCg
4UIOeqZhzjbXIeqTDyx88bHtwxkSq3PLiUZWY3bo0z8aQcHtZz+KSK/ikOKqXVCm
wrdNEwp4n+wnQhUNdq9VGBCkWlcQq1UlIaShWJX4orKxVyE+b4jsIcjkgTV0GD4j
tXy51Ad1/CM1Wb7NAsdpGHo22+qn89SFB867A/i8Oc5JWOMOo2ZVk0UYIrvBQkRh
eXG9fgolLFSc8/Omcfj0VS5C7AjocRYk3XnhRLD5UHGBRc0btlMU4dS3coQUpPWS
T6Jibjn151HNz8Ck1UAV04RwIkTIpbjIP8ywOm1kJ4PI4fxcLGy2cxqP6TxgElNq
ICG0MclhjEq4J7zeA+lsUDQxx9t6Mqip0T2IIDsDu/AqTXqLsG2EyO6SuKQZCpMw
IDajhPfBdfQse+uUwbSatX0B5yL9ucP0FuoXnoWS1SriZpT76nYDfktilu4SZrzA
5rJHkM8zZwJY5nFoxIUeKJH1ZwruIn8AKoSXM+nuYMVAYc3AM3wmEqyMV5nTs9ms
QL3+f71qa/r2JKYHT6TWLGh5ui5K3znoiVxcXXjhhzt2co2UerloZ0OJZn1K5V3d
sktdhlOYJzI4fYD03RDuuzvwax1HtFSeOZJ9UbFlDSDXZ37O/tQDXcYfgSWyrr/D
zstiJkjN2WDszOXzPnVTx+rnUaiDk7ULhY1XasNhV471qs1pXespS90xmw8/eddu
B3g4sHJnK2U9VNVMWxRp9h/Ng9PLfVsluCyAE8wDvyqzliVZf0JPbfzfICS6eT1d
gI3BPSmln2LeihAaxuaMF7hDmDzJFiy8Ob0Xzz6pj56OjNGCl0dP275V79yiG7Y/
EZAztiju+o45EJEvCN0OQX3oAok1+EqcI2f4mha67ftKTMKHpRjtqnUAuGgvcAEA
elDNifF0KduhQvAAhnU8pQ8z5+Gce51jZ7Qm1Gjvkh5q0uoNrG32Jw2PcKjPJB28
HORbTSF0vIehHEzeXQBfB3gHWaQG7uezlFijNLhMLzvVpoC6pB2rSIGijDMu/Xov
DQWddYwUD/mOkHLkIA1Vx13xDM0ieYa6vuumNUZHr6i68Kdiy3sd0FT/7aJ9iL/o
mVULVdqNqnTN2JvpSRZJ0i3z6rrgpruPoiyRajjTsQujJtCweGxs1gxZEOhMXkXb
2CJqkYFc/ji0YRBo/9yI6CjxlHzerIjM2ZOrhEo9GtgM97yhQxOEyZkq+lsHfqwv
FmEf6ogYdtNVf3mixLrcrFc8hzNjFJE0gKpGXBKdF/NKlmDQyHeb9IomNy6lPA+v
SdPtfbNsxWQkcJqcMMrq1jJow1AjbxEATgHh34Y50qjpoUxmbarox+XzhRHa1VCe
GtKofAjz7xas/d3iM8aGOKN2OFwOLaEIBERWwuAFTpSTehNj8aNI6UVM/4X+yC7d
J0GwGNP1/wgj4QUrFHLF63pqYopDQSWtSKfA+oXlhsoud9KPMi1CKHuYcBD+cc50
0CTCDW6JNLDUMqy9OKTw0tq54ZgYAxq5FSrKgXgoQGWqZl/82HHK6w8MsntxXuD1
RAyTJDj454SNd0u8tZNxJIS7WCnhc2v3JBcm69x+f9ds5RmQ7MNSVX5hZZaJ/XEr
n8v0IaOOqK5lHf2tPzajKYd7DR/SaIk56FZBzxDsKZYHRpLTIUp8bXAY7AsznQhg
W0Q5gcKbQIElruSnFqhWJu59d4muPz3JFRFESjhr7mGyXRser63cMS1FpeJLJHSK
I1lAM8FS2blRaaNyrRp1VtZrqORGgu0TFdUxHSlYEZ3xn3T60H8Uc7MXOcvfvu6q
VGfLz0msONy3OPQhVXs7WlSD9jwSz4TBCDqzc65M11FTRgpWe3IZZ3YaNNiOjpI6
AYQrjURFPy6SxRFBh/02KjVjvUj3Me54isA5WE3P62M3OEro0K9MdXpi1qLWV2C6
nQzU6pt1rEjjy/F2pkeGHCs8UvQIIGClnsF15imypHPglWpAYUQlDiaJeKvm78xV
07P5fFAk/WjyZOjlipfehKeG3YhvFoNuEq+FoGo1e6Lo3oLVCIRxVBYyqzraWeJE
Qv9UfYlODNhPQAI+WnqQTrbRYibpLhrurt/As1YAWJ4HjT3pS6FCRZS/bcaYsAff
7hcIFxh9ojWtcvPS3A/wYiEfiamz3SzwDWXTyF7owsSnqKn6bz+sJm23y5DHmpKq
g41T1bdiZKjaHhDdUcJaHH85gl8xbTQ3jZ5p/LfDlP8wjF+PxAScusczTcjpNNnt
q0RgLlqfH1FO/StTC6QGZxJ1R5wkXHgoRegwyncMmANG0OLlejgSWQoLXGcO/zGU
PqiWSEf2yd+1J87238MoWOfscEF4tRnL9h6hTlUbrBIkaa1LZhtbDV59JrtSuiW8
nwDo5NrsZEPWWoShFU2O0ZQdSk4UTNOA+5MdHsGV4TSCTzEnQtSBDCdhlQ0kmks9
9rC4eJ9BaMn0Dzh0Ki8MPOQKHOxnPGcDbW5tC3kfAkM3ASX1DmNrPzjX0kqLA8K9
jzIyiw2PyG6OQHYgV8VZoN6OCcGQqw8+Fd+ZrxNja6BcdbkFM50YG1pJGy3ZdQe6
2SIXqG6N6BuQ+4EpxEKXJ9zefu+Mx2+QiO0IZILExn9lPWaUH+iY78MyYzow2I5S
GZP4ylcnKwsTBWc7IQM3JDGPHMELvKkbr3JWWfSZRlh9DE9PdfjbZmaUbM0pIYks
tQXoXr2fQ3X7xjl4UwzZtz2PctzQO6dsc9y4ID0bxH9vVYLA+m/db+l3HSwLWdx5
f5IWo9e/X6vlKkHnWKTQUqAnldN8N35SsviUGgVucqLAGQn8H8JKri2npuO7vQIa
Va94ba5Tv33HFW7FNQjd49JC8qwqU9IOhWtuJG86k9GsGsKCLh/OSXW3kevR+BkE
yN9HEQFFhO3e5rb++DDKS9K4n7Lqkk7L7QCwZGYFl4W8xGaEOFlcn2/Qx8XfAIZR
J6EZdzVfijwAjttE6yTDM96FnVncub17fzSYtpBetKkKGnYvK3P9pausnH566OKY
ZuIWne05nswoKAuN5ghaWz4ZroLe+0b2pXru/Sx4c9fLgUgmXDw2d5GPyoAJytIQ
SSB1exW06zUdY0LKpWYugOjuN6UkltWhgaLSmodVKuXrDSRnh4gb8a91IV6Ufc72
pYBDCf47YDcpQrACCnwUJGPU3gs0IG5D1cgCnPndTOn1f3gED2rbUOXey0yL7Ujd
Tr9tUAa15amL9ROUwkLIktLp5e0XggwjyGf3uk1IiggGiDiROKdaacprVu35DjNn
VjEqzTZRtXTRz/lYkD3JavvR2OARkWjWTepv0+7T2BaeJ+/RK6ls4rHOQoauxsjX
xvYeQQfa6LQXkeLIKKdYQJHjq/LduWhfeGXf+zH1cdrhbYabmMU7GAmDig87/giN
JLCziJoObpjUGKhQjOvJD/ltUawk0UQuffuqu1c623c7lFIGnqmBGUs0W+IRol2x
ClxgrTgjnoAhqYfO2c2QDqHHm2bFfdwT0QMVe/CMLPvjgbaBV4YBivTlIL0hoF5Q
0qENH8eAI1Xs4dilDnLbcuTH4DbkPqn4iMYRUlyqf2n80NMlyAFUlAan1WQiGzQI
v5wz/PkJpmnI88A+B/sU+THkTILcn4LNzPeh5zKHraHl4l3grQohIY2k8nCX/oSt
Usr8lL9wMMXyoRucuU3We/IuwqAPkPZnY3CavxreJFgdBV6wCw+J/dIqTb6/J6z8
IdxcdKpdwl5u9VPzRnkTl/NZETTG6CUlmxVyyzd6kq/GEj7J5uj3YMKHuKhfndXz
1S/fQL4NXprr7dhYLemGcBcBENdOZDJ5xoTGPydH7DRxQ2XNkf4j3ug5QFacUVSu
dMsJg9Gqby5gVpxQdMWxKxQrSwyN8lESyoVMJyYiMNzSwya6uTu4D4l3HtQoZDj2
5Iy0awcaoPep+RhL5/2WE9ZLwUa6TaOeeYK/kxMCAH3OJJOY2dZOX3FPA0pSlsaq
VwJlszk62tf+tO8dzkvVHt5HGfMzFHr+c7ZopMEgjQAfC9wZIq9nuTj07Op2Dca0
V9tWD7I5F0Zl/syrnPkPNEj1CpvZ2CKcfhJ0ZSWBqWovtNr9rzG5fsYvxdPGA5TO
g1GgleNIBtC9zNnoNGED0MLg2FNjJXzezSwscymdF3wj3Ao+FwoS167HtEad6N12
sv64f001SHTgXPxTowle/ZjrMZ1MLFQ++GdS0/rw7Cc6gNGtJR+Z0q0GC//qX/qi
Iflvb5sAcr2YQB0f6eBvG9YJx10/sH6jN26eqMT/JWKI9/7KFn0HGoZpXvHbQ9Qz
ca5a+4l2GfYKyWrvQyJmHdacCEExksrQtfmYb4XeBuW0AuhiMtoi1pwjmJ5vz2T/
EEhCJZwxXnp/9vRUQi4JGaYqh9r++3iK3k3lwL5amMRaisHh5KlPNMYZq2Ep6TOn
/mf7YUfvNTU+J7hNFa6XLmNr3kKWL/foaVSkg2tnBLlyeVVcKW81oMVUND8XMCOh
mlyJ73QFA6iSwqIH5OqWk0u5tAD8ZpMbdFbPvs5jgYEzW/hGjp0CpGutxhUmy9B/
YF9eYRvRBFQyejtYlRX640giVYct/Zyv59DL+2Y8rCc9Ao0rSOkouLjhgL4hU4Z0
NLY9FCQsqWBDXmA6asRVynpZv7lMDZIcMBTEJoM8m/bezBj4AIy6QY5wkpXpVRBM
S4b8UOEYRR7FmOf0SviZN0yPapMPrbWJm8+oGe3tDYiVipM5wwDxw3iNIa7Z8vmR
bfeGUN3bfzPcANOy2o9V6LHgVzU07DP82qyjYRmwhhhpiHs/Sut06Bq5JcHTVzYL
pFVT+ubITa/yK4iphJWIao/kga8itcBbo5AYevIqZgXAfWhK9vqmKn5xXy1TfnSM
XFvSDRMXnPpIrHgOnZ3Lbsx/4fhGd/CWDgjf1/477+luKsa4KX2P/GjuCCf7ztrP
eaZKIcx58kBcIPx6HX1tmoVlL/KQw8aFLcTtbxxVuGIXghl+VIq/SG9OyCJHYL38
BCg3CrJLXL7h3z1toWkzLELauKVnx4Pj/qVcdzw8nbEHoYeg6eRiP8185/C9Hn5B
ciyPLTzi8a6c4JDRQkS61ZoVAEs6S5WYBuchLEBR9DsxyIEXPyaiASZqdTaSaU9V
28QCLCzbb9UHNxbjwk6gnPIca2pQ732A8z7W58gYBJKocKJ27OfZpXpWLQ5z62Rq
bIXxX+SJMpstAdsUjtrtBkerJ0ZtRU8DdR4ceE6h3BIdsuDWnpOrNVAAjtf9RTBt
z5bGFwcJrluYs9sEYwroz7dpqoKAE+FDWzaxBddbST7zmKcj7U7B9jjWV+EwiYb9
fY3JOKa5ooPBxV4ky3eutOtoziYLE/JgpjGmgNHTVj56Dh0Hq9tkJcQsAQlR+Isa
mzR/KM/U3OrUMSj6NgEoI+31/Cn4pZkXZjDa1RalOnHYRYLkzHqGj0GPyblFzzWw
WV2+Y3xVBGdz46b5AKCJFBPTVlshpA2qRJGdQuZ7su9kHjQe8I7Zcg6RhegEFnL1
VcNYQX4/XY5cUBgFk86wqQDDzc9AKyJk2aU8umIcywN46X5Z17Mvg9oUp2H1kE68
9dGV6M4CiUz1ED8McqwVPjp+Gbr+IX6TGOnwg+WA9wZTH96Eaf811CF+VaQ4iTjm
bPS+Oc/VsLgbkJCfRWsCF5qX0cRRdk7ZSz7BxJEVbQVAFqdPY0eOD1Os/bANEMlO
g+yY8JYgQC7rH+X1KZToSYut0QR+tXYBKABFTgp3UK0h28pmayC0L54jHuRSiasO
/91URGTtqvFkSePdrOhohLq1ucZ4Ha375IcOXfxqYU0TAxa4oxNNfd1ai7jcrV8H
EdLyrNVtLJAJDBOFyYOqlU+gY0S+OrUHpaqem50S3i8eNljiSC9qijSMQdLZzUAB
50ad50Qp21buim/a3aKdGPhfTdiywaHwOBa3FrmAUqfVYE2uW4OZFTjnprVNobmH
f+hR79CyLL/IIMEdZR/znSepGbj88qGE7Q+9Tl8JVHNiicNvzkZ6PKigVawdXg4s
E8GgwTxlELk/lOvdzuoTdBu5mjOlvdfazQePzzPgs45qHHmkhZIEUMVwPUkykMDx
tYpwsUmhSsb2jTzkuX/f2CRp100dHM7pFqG/yhWJLJrIAtTNAoAI4gk8pNU11EPi
1YSoiUB/K6qha/V7X88hnSDI/yrMxa5nlbAOVC01twInPMi9/l4CNkAr6sFfTL2p
KufiKcPvLXR1yinKSyjn+e/rlFqTPm25NFHDvsbyz0Grd69sdaRgrXwaY10b5f7E
dEbEXZR/WEML3p7yUzvwMjKorFYKTXxcYNI37u82aQWMlU4gx1u2S+kj9/UAIZp9
n5AoVXps/ji2Zv5verOVyb5qbFdVL7cd1udzomoJuPRbuHDjNZURy2LSLQgNusF/
q6vrybSl79pEHTBeVpzQ9fmo0Zb4pdFVS3LdqAB/FDx2O4Y8EgYYSkEhtZNF5iKI
YbNgcKYiBVD1CUFEDC8y/5Gt1UAG1Er2lY0lmlskP6NzY9ulXnruUk+qzQNnxeMA
yZEiQAQ/aDKoyQxbNHQ3YOR65uHvmFfGRhkbIpHYNogITq11ezJJHYRs4heoL8/e
rpdiRQaTBblAT0OIAeSyQ1pEzXs7LBoMfS9jKRPi0ulTawsCUk+GopIzztxksk3J
tEdpveN1yNBu+rU38b1Uz4d9D9i35a8Xob0/rotK2+D6zYxKOhZQIk6vMltMRIns
m5hImaRhxBzfGJCGUX3JNmJ6wPO5qnXNoT74ICEkEm/nVI1SKkjTkDOxQdbzDlCE
A+mEU9HMAoahi5SW2RNz1Kb2QFj+qSoLsSEdYS/pxaAxAtkr9UMIcDE8zy08XuIB
cXx64os4TdDiiaPUV4z4+EBYnkJSCuaXmmftY6Y4QTA65u/gGxqVLSHOsxB5MIpt
G447g17ecLgFF69MzITe5FG5Juw68G6qdeaEhT99xp+YSIPRFdyWEAkkwIrKxDn5
0XWB1S9oFVKEe8Rb/2iZ0DbVNhprKP9teldTErHjGeyn97aYlpzXI8L2e879iclW
9j1XSY1SeURHmAUxbG/g9izK51i4xYQbs6dxzi4caJTLeURYEDOEi4ykYOWSQsNQ
svaaaMnn3o7Ygn1HZu9WY/QUn2rPfsiyAJc/4ApUYa4Me9UqwSzw6sNvTEDa9bsO
Sy26Qg4mokFoSGN2Kj+UAcGXCPhY0XOOv8Jx0zSqQjOESc/HihlnbF/YTihwUgWn
PqDjuNbAf6B+yqo+6BKQWishWNKNeWurM0lH2irYnuh1DZFH27duSDf7kKu+k1VN
+n2voAzsUI/sz6LWZ6O1H8Sj519jYncz4nLRgtHdZifOjFtEYc/O5+pfkGqJYcGj
us3d27lVpFrGBSNbgW9Tp0ZoCDmNEW3Vmhf4Y6ydL1R0ve17YmvoQaTOfIMJLizL
QTr2aYU/buIiOM0buLCXuqPd+YdEV1hASnjqBaTz06gVGLY7U4IvsWWmvzAe1h3T
3HL4CsWc0XoK59l5uKzV1KkM+bCOb1qjINh5alVJr5Y3j60nHvI13VsNAUUPerMq
5iiuzSvlHjFTn4pJAutayq13PROSenR2urIFc+8J7CWQlxX++960uT+HaAD9PJMe
xZupavwovmxIbtfhwi4nfrS+W5qAdUKJG1TjPTCIIw9UlH0i3oM+C5n8seL02gRr
h03JWtr/7XYuBVkzHbOvNCOYXWtnqXwG23XGLSl4gFi56encBSjXSpWRWm3aGAJd
vrczv3hBrD68/hBEshr4/t7x0YDGgAcb5sV91EjXpR3zSs+k/x8xR8kDP17Ft3ZM
yekMvOiEkvamXV5Vxi0q8kEur06t380I500/w0Iyb8qfoSnvVLfEutkMLRpVjekH
+lhVxKUJAcI/FcJixHegMRScTEzpOeVOqjsPp5r4HJFA5STTZI0YwaJ8upxzAa5M
/qT5MhRxPA2Bo+8FhMZ1vupXuPzn8zuIr4Hbr7xThB4MI/3l/FH7uorrv70H354O
ZUY+nO55xhjS3x8t0Br+wWArL84SO1lRBpw/0AGFNMdGOOZWEh4lffuF38wyKgoA
FIZaqDymmz45Z3CKu2QShC+4wqRAgrUGixw6D7sNVmIiVGSwP8pfKdUvHySfHq5w
d7h1ICEOpFMpd0Hb4Wn5obfkq8qemQFRoAg8y1T7C3Kzz5FRryCwpBl7+IHO1DxT
lhmfrfqYnjtY1G0+TkohitHdJTdBe5FinjR8dk+SFuAALDnGA/fty2lnJtjuhldH
/zGMk6MfdS6Ww8qhxTpalxWGNkGuD8zvQy/seElDLUPlLCygM2MNM4MLmsDv35lm
ff8lwFubdsxzj5hHbRjZrtc0N32AvijuKdnzcJ6F0cq3iaDzdeEWkRSq4/YjHJZ5
B6jKgl0PhrEzWZrUdTNmHNh5/k4PNf8P8F3y2nYOZWrzrHAw5X18V+UVadVEpS2k
E1YS5uTq+30amVWVcfQhxezQlrUCRnE+UJvgD3d59r2UeB+YyaEzRhnuQM/6EDkw
MZjoiT+8hT0xsbBf0S4YYfGJC5enAjzPsZ8TjOqr57AL70CEsNIGSKBkgQ7cH3wB
z8HTKjCVCNEri6OId9QXJHmYroE5B9I1qxEgT3yd2Wvx39QppWeHt25ZRi6P1gbp
yVEyF49TWpWuWNnBYNXjHRnUa/cUlxR6p9uUQ++g1uWLf4bgj+PR1iKZPqd9ZJH4
Gc22WX0RuqSVdz1KBRKcI8LhWDMQho0tl1NpDI3YKwXP4bbr7vBPayAyKZjYeaiz
10ZQHKpQoxu8VdLz8vr0rRQ7q0KRIF8hY09LdfZS9GRPV4P1VXwifSLm4KQbAZDe
oJQQjftUKsa1Etgu+ZBx04eVVxuAx3HwmbVaKm5MR+Zdwu1eyQqXo5btrPJlEHU4
OvdtsOPxCrO2crSXJXwAFYovWWxThR/FRbJePrJXUUuzug+Gkf1Vhr4fgH4zM7Mg
TgOoK0zmgF2Lgofj1GTiYOu9hof/uMdeaIvN5Hds04rk2VmjgY6ag+zuaSLuJ2Xq
yY4cshGhgte+wTgrU44Cc9sJJRgCAj9QGtLdmqg4qF08ED9USeaIGrSlpfmWqppJ
UYq3NYgKqOkJGIlUDpxb1FtMOY4DUsBmpx9rGQxYemsUPNolUgyfRwsnXIRJ5ZUb
GEtn4xryiPZ4SiGTLjbCAg2Olk/LSgAP87WKC4Kiof7/gMOXjYdD7ann+bPKoPyu
DShutsaDoszvtH8pPIVDPRPqc1nU3G6JY8thXF4nnhr/2QSo5mu5ZVVTrXv3/M4i
aGeb58BfjibPSBrAJ4m/vQZ3GXEJg/jJR9QSsl/X5TP9TeVyr9NjFkznHU+lB1W0
AeCQX0H/h/NF3T9JaN61yQZX9aUQ7uBGCpz/awbNz0/sQj1CNv9dV4v/92pWQvfv
6UY0XFOKcladwAZ8TyqKNmggDNdh5A/jE5mB0momAg9cwIJ0+/OFQoEShznRVEBR
Dcho4xYgWBLFncFtY3MdYAI1qiMuk12vStNOLflKV0hUkhFrbdh1nVZqE37r54yq
4XoqU0ws0Kb+er4DzK+fvNLbglDmVMYKjXr24fvbBJmDRG726Pbwt7+6X+Z0NMuJ
eYgVFSoCqbQpbZ8LxI86jijIC9ZQo0ivLraQW7LH+apjZ4rTLh9GqKWUETi9XJpc
3m+Ap/90WNIFf9MmrasZecazKP+kUFj3gIlV67Avds2JNu6rbbYl+PVFJkvld06O
khvDRPBMTmlzeXxqnR/iTZV+Lng764/Oybshfz3ZMMxKFsoJWVowjeBkek75iGat
ZPCJzwghQ9hYVPm0P8KvMX6yD20sjhLhplI7a9U54KfiR6vE78y3+kKMi566yqDg
9eDp3IPwZfJP5438VIBcxk73E5mO4HrpuBIsMSkitDo7lh+2tTFE0GhrUlnXI9Gy
yRktUeGnzRk/BD8WpgTCq2OlT9l/DswQ/aLYgxgHGW/o/7q1Z9kTL9sJTTEJ2gGM
d1avlFgVbGGAWdIvTt7JdyBzjR+j6kc4p7TAQUUxROg+dQ8dwSfC7sqPA+k/TkGL
fDoffYBk94kvzFihqzygDxEZJyqoKOPGGQJiv5xhXjbQ2P0sI8Lz9ZxtGal24X7H
W+5Buox/Y+RAbzOwiQUj0rYeAnG2aYF7TqhdWGx/PoyK6oc8f1/v1TalN+HalsQD
WlxSezvZEaN2Auu0Cv/FFAFKrMP6jleNMK96Sqe0omXBgwDwYzBKCm91D/QrFo3s
JDpRuu5Qo05Ptyd4GQuZDFuZtNV5/0CtmFZNcEOOWTpJYilGyJ/vMn9JYvAc94jw
KUxGnEjUkARBCsH3fCDM70LhghlYB0YdKDXAJ7woinciQyW68P60xARBzyCFbfQk
kowusg1rC5XbF+pPNnLYFS4mwmeZBtLMFzgwNKhw/QGSGQabRrgd52vaJ48ZQ76V
mIXbppxldZ9cKCNMOZFF43zMFXPb6kE+9NNVqiAcveNFrm4OF1JR2kvMHgLEIcUA
3ffrCYJ5vlICA/GqY/TdfXparhurKc8Y9QBKjEe4cwJtS6h3/BQedNVM+A7cYsSf
1mT66Y/wYMBbKnxTtdyV5ua4mW8DtNf39Cd+P+CpPLok1RzIvntfpqzDt5wWRdoG
49WL3NClkCq+ovbtJH+5yL5ruaXT8ko8JLoBwtMKf54MQ7J4teABb+AWnkRaKeFV
N5iIKBgRWvRnYLyNy6QLDEbILtPqUDuegaQr2c3rZvdY3FXOy6YEC7KPYdlVB1ao
8HtZh3YL47OJU3saEiXAbHx2QMKVI12JnC+f75ArbOrzX7MA1sXIeJzstJBva4u9
0nS3RvxM9wc9N+x4MbyDYN612vLZgJ7sGZuuFxpOWYg+De4h6CLsJzIlxGbMedcz
U8wMnqz+ofPeS+jwnEUz+6HrlQB6n3+8IP3K76jH7Ul+90av9p39FBPjSh889Bho
ZYxjRRjtNZax22dm42wQWDwQUtGpiAQrbW6ggtRLNFKGuA/yonqKymnHZFcObqHs
wi/NwvKTHUpOHSpUXn0kdW8Be4uIqkI18L7UMQvu1Rg7J/bLECXpPNuPL3WTQOlZ
HD2XZtot81YNSgsA+XZiNIrMl7MAGbT5wZPDcJZ4jWk2z9FiSnuetOsGlSxt8ASt
RmSqKaZr+kJekJw1908nbYYckCPGbEAb7MdV1MCSIqymL2bo901p26cM2ji9Heyg
6GLcKanWIQZ5OP25LbLhxw29Ycs6iNJ9La//uGe2eiF+A0VxQdUR/f71OaEdGNYn
oQs2tvKWXSf4Y4PVdB4g2aSPOGGfE20r7cn8UH8/EI7wpIBckwVKhoaC7+h5OgKp
nyZQLDkxxa2cUXgOgk9/xiVkp0mr3sIuZ260d6HzuqTOr3B7xiksS8Pvm8n8m0KO
erG0kKvpQPryVJzB42lXDeHh6qwjyIbrQ/lnEmzjV3xcYjpHd7g8MBX1twB2QZ1e
YsjDeM6wS9tl821GWqz6OrRL6f+DRMz3AzoAZtvio89+Rs84zuUdom4/SSZm2fIH
GYjGI0oX1l08qqWY31spyGIsbfoM6oTObq2XOp8o1btybiijeGzH1jolif0wDcAP
u7t1yCmrH26UJK0sauslLiwA0y8alsR9eCw0A/yRf7FZiwvbVOsl2tnrHhibof2J
60/bKTYJ1ZXWU6WjKSJRrcYT3LGFMYaXlRW2+1uk/yLp+9GIuk/A+FM6YwQnciEX
1JclgsRd1NN/ZW+2HR6O46v6SmcKXpFOcXQ+RJJdc/EylCY5glOuUJWqfW+avvR9
uBwLzSm/bbWa4hRD/zPmLbTGsVuw9uq1pV2ysDUPswk8ZvrNv/pbe4LccOGL84VJ
tCT7Qt6JxswkfO9NVH6FO1Kiff6KP+WAohKu75n4wvEcRXHe2HaY2XLQIAVFiblJ
lBt0oPxf73mdMrEDFr3oqOVo0yAg6qn7bqfrYfXi9ULlhIrWHW3Tbheb+SQCKT8V
dASh7hljNvkatbuEC2ZfXJ8ABha8udJUWHLZlkVLZCG3gEXO5AOyIkdF+d1jfuBm
wIBRx+vWAx/jvE2BHcqCA59RxBfgBeAyeoV6wSSkzSGIpCxxjHjCB8RGuf6oHH+Z
33kBRO8LOXr7P8qf+sLx4isr8Zkf3Hd4ZruZErjd0gRaceEHCdYpwLo6ieKnP+vp
Wd+h7T4XmqSKTWeXC02inOnDxarnE1RkNB/Pqs9TRtX/icHgMTWT7BdsrGXNVK9M
OnX51nwBvdY17CZd9DLqFpuGSdsj91aL+OI6lkTB24S/NW7CDtKflZRtzWZ4I4Ie
sb7e25iRvf3k5X5mheNw5wbr/9p94XYcAibwABn++5qEq2uPyzrDkEEDsdg2AcRz
s1rJp2BHEdmkGbC9ls85n3mWFgkkpPffjRcZGeJGsNG3xzqNhKavSYQDGj29uTJT
rDidZ4N34WmaONgKQXsEJJHEwcE6EVPQ8pvUcSrYaIoXIofErEr/+535Ow46oNei
zyF8K0q21pvNdVlmibKsQ/vfJF1UxaURRhqwgE06fqfeuD37mrPQ4bpqS2hSSC0N
g4/DomTksuUbV/HL4C+az8Z1KVE4be4rnJ12IobkpMRjAt8PQ2tf/77Wi/YK5UrK
nB+gMJppVQq6ILDF0TD1hZoUHXVccMAux5PI8NOSoBpMndkHD/jzqfNUmokmK+bN
NoEBIgOb2qpCjhZ9Lvrs2HTukF08F06Na2b6g/eEpMsTvlENvxosNnH19Os3Cm+r
6YsyX70T3gDU+BP3mwAyBa1gbTOBq/INtwxoZ2E8X0WCi+w5zZpSulDpyG8SMOjq
Hjhat5W61cH+eANomoOeWKlF1wJsFkcD0NBqrx+pEa2Kg6pVC6NOdnS+vLCfnFTF
qP7AwSsFxd2JeT2UeAO95IcM0GuT8Nq1SkIPfpzBT/U4Tx2xc0tZHe6gm/mECDv1
po6Am3rOu9ryAg1XYR3fFAxE4MAB99qIANjK+f9mBW2qAn7f825sLSQyxUPGt6E9
ddxhSqQ721nMKtJ92U3iH4V1n5DsDv5KPZ+jKfBLkXuI8aX1jrQCl0EWgGlTIuyc
xbSDr7YaS8D3DCU/OImARr7Q56ju043pNdZeAXzxOojhjZszMDrs5J8BQp8iT4rR
VY3PIvT8AZTbbwwJLA2KHIh4jXBe2eI/cai4M0iUnnffQxGJxyHUcO5Cd7aLqGi7
9lktxQ2qjyo6964QwKlrWtpNRRKi2+1nvBo9xTxoR0Yl6vbp5UyLYmZB/jZvZfa3
kvu4jq0L9SdurcHcMVfUt7dMkAvgh4vqYXl2SeH5K/qsxOPG5YxtGRAm56Pr25BG
Ck6ddnqmT/TVvFLnRpVM0y8dhdTlf8wey3N/fISS/NTGMimLOOWvPh1c+Tkp05VW
M0/z8AAn3aUoztVskjCp7q+RnVTmmYwQVqWHmJOab8mTvRU8bbHPRATEPlFVjqI0
0upwCtbp1HL6YdjlpQimRbp6Aj+H6ySdyXRfOpz7SrXtysMRvIJuePbGsqPZUv9b
CNGLZW4HfW3r144GobXZPkgHnsasXBVbaub3UE8tcM3tmEBQ+2ROkH2ubnbnrKoz
lXCWfolgkDptNVtPSsdC3rApJY73/XknTpWIkBTLMGvAxQpjP0VIfJr9ciH1zuvV
/jmpfw1b39cZ6DA94P9EECwY7D0rx7g1enKAOBqy/DohuHLbnWwZCNTgmu+e7zGv
nUB067h33/6+OVvtdTlGCispL02AM7epsdqMDceJjga4IyE6RnLpV3Iv9DVS5Ra8
V+U8D2+f7Xz6T9qDTaJxHKVjVr/zRdMkonr9zg4Mi7V+2GcOBquXSZMQ0JfuA4gK
Tx/0ZHrYtVP4mAk6T1kL042vdRbKPt4uxDYVMIafG+wYwTlTsdv3yhncRFlWgmPO
mQ7PA1nUp/nzmNCGnjJdfYhla7AqivD2cxAEipntTgIKPhzAONJ6iAhMVGjyG1w/
4SRSUT8P5FQjZLc8ha0TLX/GPajtKuG3Fk0TAa4AoQQ2kLboVpC7g04QdNI8FAf7
sgUarDCokauuALXGBvcfqELk0f3LMrV3SJ6EH67Zi5GUsZyPOEOBN7kEjDpBaNvd
O/8UBvmbvsG85uEkiMh5wc104to+4JsE5EpOXgrOMrFeVRQIeHPvhv5s0x51KgxZ
zW002JUL4T0/HN41REddTpnfgpmGSJKFZX+Xux8fJkFOCC84vTzE8lvFdlrLMese
udTxH5lbNg3kucDjXFBiW9z4v0Sleq3n2kWDi3UJwij1ov49kp3wqpLWb6lvTbM6
U/0S+kUdoHvVVjzWMhLSx44L2nbYevIV/H32cKsyGqn8EJbP/Uh5Xn9rgE4vb8Fv
aJxu4ptKrImhuCLRBArfyKrVUDtAXeXFDEZiTyrCzPAVnntmRsuarWd3qtusDrwx
RX55isExWiMmt7lVHYHKDdFPffZG7uUxGijzsMvhPdDR7rsQvtpveBmCcnkmg3hg
ro4opXNGxc/77Y6AQFzOn/y0zO14/SAdGBJowvBEYOphrpkQ63cvuAZAcsAW+SyQ
K2fNcGs8XfGajDpHhvtQ1uPO/KH0TDlGoGi7uhdKsK9/zqWkLUUSL2EjGbp0ylq5
apYsfy7FzIwxRln06QsKjUAgGWZ6Cbn5VcQqTjPXMy2hSyYBGRdK74yI6kNMx21X
TqSCdg1U12aAOBVbwqwI2boGBI35mRcHPOoyK/d9KxcDKkrVNIpM/BA/lCNV/Ukh
7cDkEM+2RTFAAB0rq7N4mX+kHFT2d2aoUwq331nZ4jXgPge79uLjheblEZovfDlx
nf9600claFq+3fK3+XuJxzVotyEgmdI4aZ85Ro0r6knR8LzCoPJkP3cfao6clgAg
swdctvPDoOc1bAHD8bpWinGNsNDGFj59sa43yqarlk//GEpYHongHb5E3JdCU+9N
TgDx7kZgqpd1nLQbLf3N28gQmSDpI66jn4/Iylups4GpRf9vzjxDde2bcoihp1TB
RPuHkZiQSb1MVAenadrEbwtGoulQfwFzljJyFO+60KTwQRDByj0coG06z6t3lB4R
0zMJFyXFQN8ss472z9PhI8T81SAK5e2xVV/byPP4bW0TrWdh00HwBYs4ixIWKT7L
p3VAfMXO4txpfLDwV64LIzNCGKvebkXMeGgRMQl9CknQ5OTpQdxj5XEGNH08KOMf
iXAb0hf93/o1X/P6XjgdLqaPiO4DHSxnVuHxa62W5t+kWM3je8H8D7ARQM6fbQlQ
rNU7zLIBWIwy189PinkPrc/+3Qs66+3WSshPfiTxGx3XrHlx9PTS5PfSiqm4vDs+
vjftXAgPqA0tL3CVUgZyO+zx/NJKKVvsTiDMa6cEaKBmyoyVOFh21NfUM0AblxLT
UmeqfEjKryIMDITgfv4mrV/bgkqIn9HIbHt2dUdB0+hHP2EeI1A5R3n7czbkihCO
Ht7bglPELEWSe/y/LpCGTdthrNcz5DKZtHUabiQWfAeTECrW+2dEF5UMjKVhI6W+
PGjGKWwGIferg1N/XA51auGRGsvEd5SwRt1biQxWlq8K1qOTgUMEyLC9ksdqSWOI
4ACAI+0ksroV2ba0nyMARR/IBA+tHmAx11dgZcWLOXEl6zZTNGP4+xzjXJe9sKsF
+ErVDnSMaLl1RcwvBoRHBl3r5ZjYkxb74Nay5apeDUAKDGuLVGBwKBc8iMVnAZVG
sd07jqByDHMKaMCCTQBKRiwYV21ftT0WMPVo+uJr/0CiMe9G/19gJl5y5iS7ToZL
MGSq/WBxBgzmZPwxgyRzzrAxD4sCnm7LwiJY0bZoEpuLf20z1WPsrqmpeXgMkQ4P
HjJ0RId5Mb5cAmbuSqNQjp4Z8V/8uU0josoEtkEnv8ZvYwIBrcXN2xBRvIYFXxQK
vPrj4qtiZ5x/HB+uOwYWMfD+KBdt56FVZg+QAcTvubNDGU3iEAn1DHsEdyZZb4Hm
uTZAfwV39FJe0Y2ZtIwxQnVEkKjgO3h8czn0Szb73i9rB3M+es7ydrx3I/T3hFHj
ejf73o8vZIwSfCDmtrD2gSvwzeuw6l8F1S8Pqv+oHiWQ9RqDJ7aByDr4RC91iF12
CwwRratF/RlN3EePlSY1/T53rg0rd2NI39wSs2eZuSd5o+s2cO+xh3hD2tJ1rrTh
+B7QQN2h1b0R0R3Kv3au34sNlMsxb3Xn9oRWqB0T164srmmmVFBdmZrL+xALYNGH
GbP10sAj8TSdlzygSgCKLDH4yCrvFSgkxZ1w1LB60ADAv5XNa7lt8MVa9ig8dViC
4QVjIq90uMrpeR28Jexkn1F//CBDy05XOYGXIscpOO71M/XGJLPyDzYtmuD+pe1d
sgarC4xLdocWvMAfVDXhUzEecQR3zzUQjAhhcbc4cEQTCopPDgXKuAiFJG5XWYiY
24Sf4LIszWYpCJbqw7wta3H717UXQqAsILG/8XbltvUNJ1x702BkxFx/z1O8+mym
gAvyiwgPRnp2OI+cAtrzuU754VnFJjkBPx3Vp2lHy2dFZAXdML4qTg2XAGqrPtXh
+xwaDSgjEUutxOP1G0Zxfw/8OVLvYF3L2U7lK0E/GOLVWMenZUVi/4opXyodI8bS
Bc+DdBVAPyOP8pVSJ9DDT5OgptfcvI7WFzpQMwwNLCdyURp4sNqVm4WqfU1WVIWT
cdL4zeSS9s9aq6/kNopzDucbs1ZdakBzpngsBQfOEEY9y+UkOBZvqaLII+oOC9jT
cQpjZGt0+K1VrJNp6CG2BRDjtANa3Kt9KF9jZdJ1vbMmPd3C6XA6Qd0FNamklwYq
HW/biuvJGyQU0o0McBIMCQjsnK0ODd9mSYKiw1WrG8Hnic/DwfmslZ7FRFlRweRn
2vMIin+O2zhuX81xdAoL7Jd6cHJpombDXpuBJB6FMNqyWE8BuH8tmmB3cQIS0uM3
G+vPOAYHRimwe82FhsCZd0XbkjIjrufsKnbOH3ZhrjgPHCpV4uh2MzM1zqqhB9b/
RSnGt4B4ORx9hc1A7HNFMfelNUTMl20fgwuT3XdM+KdGA0lyDJC278Zj3JOwHIBW
8KVXt33RIS9O15Mz/FMJVAh9Li4oLl8My0xpj5K4BFNB5tr0LVUq5l5Gn75p+zLF
uKAz8LZfvtXl58esfy22kebj4qwvJ9Luiyz4ug6Rem5KFqI01DTLySRjIk3w2QLo
THTBk8NCBNg7TRvbgtP/n6X1dlnAIpdiGKLLsSkZYH3Hvbh0W44y30mpt1ik/jcw
OArLnTVpAYE4Xc2uMOArvGff22ttgNbIxKZ9hXDcty4e9pmgGTeamikKVy3o+yCb
H3IYGltCmKsNtMht1IhpXeODs5lS453wS9TcikbXUB60K3XFoxzuTzLD28Xls/DI
xQY3S1kOeNRljL6e3OkCwBCh2EGYLLafDtaiDrRa4dEPHLyyH5CgPCJ99kcdh2Jb
nwCjo7FpccIPUhlDM/Br4eZwCyLBFg/LsUdtOMl3IQwzQIMv9640PJIj58V6SHem
e/9EVYVhzHF0/LZhRRFu2+RxDFxCDcVkOukYKvVyhrZE11hCqtvkb68Uwx+S8HFw
ucIggnRIFm19Jv1GvmbUFiwa7dUbHWwA8BWvJsUnmlfPvz+mDSFDEeSNmRpCZiqD
d/vux4FBu/HYHPzyxADE1Y4wt6ThXmPuKZK8CAWHx07+gInrnw4N9gf3bITs8rSu
5fvw7QYah6OUX7Br4MbMv1xPr/iRoSJNrPjeRg6dCQH0s0GLQJX1MuBJ/cqQeKwQ
H+O3a+9NtgfAdgkS5AjUNuG2ptJ0v7QOuy/Mn3tUQ+kZ/c3OUwRoQbCtdM2zN2zL
0WKPeNuOgkLuk/wdGjzeQGt9XR93jRJyJJ8xTD6fJk2QGt6gEMQE9jUftglIUKkL
vqZHB2mtPN59ie7PoMIrrXn5G+gMB3DqyJLZGBGBpRMHSCV7nxO9e4z4pHyQY99b
QbScHqTvaKR/EcpHBQ6GOrBq4WjbQFKoBr8WkE7uehHEt9bpLlwkks8kd9nYB4V6
qNusMVd+WxdrsXwf+LSVic3aIEoNV7NF49AelgHazxdClU6iVszgsXqZ9yMskG9i
kwVspnCTM84BhMM75VhNXhDscarUlau7qqiq0gYhYqEq++iNqirHHHiZM2RCEHs3
+IF8sSjl+QHt5W0cCoPnQGj3r50EO6wkv/1yu+gqD1222pmaLDegxU8T4iYrIr7q
Q2YoksRbm3yxIKN1kXdReY1UZYar1fd1iRPajP5zRhxdrHQmibWOkFufAuncQAp8
km2GRrfs0s11j0iPOnfmdMvKCNVnEwkqNJtYHD7OAvunB2WyEOw665LHOvxYA6oI
tiUTWPEXflMbherhGt6PfVr/mh2KkFFlvo7dhsxYky4F9nOt4Yi5X2L3a/zIRUZn
Ph/Z5JM3tbEVZCVRmmvkQ500bI28AL5MlpQdUWC/G0O4WddoS2vmrZ83AtOcvWSv
I0ght4vKWOHwCaAuSh1cx+56PgTP+OnHZuciSH4QXV4ojcpKbl20lDekIMHtbAlV
q6Ca/JHOFxqJ9sYuLnta3ZpId1PFdrLFEJ2uM7spy+1VmZBCGZ+9J82ityzt2FRP
/0Lo5xNU/0HL9FrU83xafk3iTX7k28q8Eo0VaIVr0Zwv9pYctdjxhY6LhgAncv0o
7m9kT7Ylb06FpYKaLZinG4WRogSB57n1QnWLjlTh00xXU29ofovjmD1UtkORtU7o
Yjb7zA17ip7bUT57Lo/hrqVK308rDVd83yOchymJ9VourKp02OHJwfXv4mWGvDBD
c321qSVa2LnvUKY7qPb8S4ZCxMLCRb9eNCuoAkT/9iFTw9YODz9uu86FFv6Y+FSm
pj7CTCdhgMoM8KvU8kAC2Vppp+/HAtqJNmyEm66O35Xdb3c8l4VRQxdv+7DEKSVz
BKZVmXRNO+VFsYGR/m3quexaLju8dzIPfK7qnZ7twUaJw8GHHKuKt4rrf8UhB0Sn
ZxvzDvXJCP7uoXKrVNiXH9sSKQVWGcW9YMahj47/7x7Elw6m0wWmAdYbeFb3/Smh
6uFdmGnMGzON7Slk3VQ4AVfJBjy0HngFQF78pu+B/H0NXP7PyE73yG8ERTCfAvLr
31Huw+Rcf1/8YuFK0C30c7TEP9GOdFw/lE2s2zVE7iru16aGTWGSM0aSkXPSsQYW
1/Sm8jy932lGFFbHvwoZUo54auYPGzXKLEg1n0IjHJbnolQM2MCSBz/IuMNhE4u+
1QbAkxzGTwU4CygBbvtqJcHef9mK+7z0N1QPCt/XwUX80SWI4pr+GgmeVZJVGuR9
WrjvdGhi2Hyn9T9XbeEw+fcPA5GZmu2CVo52xv6vzpabj6EtJgh2Em5x1mpCThCM
iQPYByjE9vZd9TGnlDaVujjpMbmCL9K+HVh7ZPpSMFzwdZX3ouynsAr4KDi/2hhA
AxxPW8Xbj96t5M7G70ZdkowARBnSQZ+qBSpQGaGqKB/wG7tA835cuy7LdO/9Z3XN
hKHpakw+tZOhTlCbxq6KqyhyRBgd9N1MfUxdZs+KRN0dp5WQiehqWNyE9yWqn7Ks
bgcai7SAsjdR8wABn2qZWbh7wucMCfiN6izljC7F63sUDYXplV+tOCOR+55/4zl6
QmAemMprOlxl+kadooY6ieb+3eiYDdBSCXaJD7xzRsa7LIdfiB4P9s0jAWcejOah
t3ptDuDJ+/jCbYQWtN2yQJxjLmGOkxNwovp+qeM4fC/nG7LLorf4b1KOjiqGjV3f
+/XJHeYIF5kXuZyR7wu7zizw+zNuY21qnKxLHO6Zut5LMSFmdNt7NhQ9feD2ivmN
XLAqZPbygtJktb1uq6jRTmiTlBsx8wCvp7Nsj/42BWDWErjllPSX1wb4YiAGNVzm
Z/CiKEbFroYwZDAqYk6Gcnyj5eUkC4pKpZWSHIjvt4lJMC71QJUibVe2udOOs5qg
isyVuLOTejWb+at4wt+dHMqmEBF/e3N43UEk/Yoq5ChiAAdWEkGLv5QFQwfO4Y+J
ayBRzARmTa/SdCbqLgDS/BAKonITwX/Rsg4pUxGBliYnFgd1+Evqr/UqHd5EDOfG
04tZ6FBct+NG7ilSb2MgDUiMV4g6qaRigKluBYP+0j9gQMxBFJ/4llSP5qgRVRMv
oYHrmcmVPd+FPnnXWSvQHiKrkJ076P7nvtVz4vEKQ4wHF79jpylsb5HWN7HLDYUu
GvEejYJYJ9z7Sp5XX94e0nvgUjL2tUnteV4890t7CqPjSNeB9oFmrv2BGhnb9UdI
sGGf3J/Zg70IA1WtXRoHsP2Rr2Vj0IMxviz7jcpYWXc5feLJTGRfPPfPqmIpUprw
CmnticK2ByvfeAmLfgfhDEXLjTXj/5cJVCo/czO6w4o5/vkqiSFDIFwhiNlF+eh4
m8GyfTLzyzTHlXtMaXzdnUwrCI5iUUcAG9LgQXGn/WPgriSWq5gU9dhZd0oZ3YLa
B4955+DBJkO8SxjTH4st56TMvTEG6M0omlNhlLDU9Okm8SsAzvotENPFxkdMqVC7
wSXqRuAC6hoYDsTTAnUfAJAJiXMpgcD6nzObsibLPhBM+EMXXypoMJzG6VdudzwB
ABmfFMskXI6kPYgdOuDh/t/XBqICQL+70Mk8hk3HpAQkneKCT25MCW6YGPmtV7dv
yES4Y3HtVZazZ3G4/Ay6/ftxaIb/ZZtJCeHPsOTM40a9EqZDdcudbDIMBBWV1LZW
/uf91oz5f6rhm0hGWmfmqhhRPWsQ3EK1PTCiLbUXVONi3a6Uu5tYbWgPM1DtU0ua
MMfpAJG6Sn5LKfj8syy2cLIVeOxCZDT59nkLXUGAekMrEXVpv2ipdxGTUvzhT7F9
PXAg7pLpOQ40D13xgMk6emZwOvbTbZ7SuNKZSVxmmFgoVO5F45w5tkxpk1SxISA2
hE1cFAGXwHzXjeTBocRwZWtgxr/HeEd9rlde5ToxnvOsRZmdNt7bP+N96nZgjeL1
BmBLXKVzTNpM/BZ6pbxWFtK7CdxF45uNxEyZYfpdKMsFY/gxihdU7wCMFUHCTpvg
vcQtMHTt3QCxXr493OzVHP84vp3JPbvkA32ApcSfy6O9CMrZfq/HTvkTc2gX05Un
qTTUhJDS0/EM2XFOMCoZx88UfDQM9I+ZCc2sM7+TJNtJD0j39GtzUW3dHvgubgHd
DdQHj99nUpGgTi688vIjwNVT+p9Q1Ys5S+4mhvXDuMUeDNMGko4BT+S1Ct60vUsS
yN2VIrKjDXfANUhk/OGjfbfRD/LeaDbWfFVjWtM1NBh5OluYpzR3gx6JfsLxs9dc
V4JJGnvDFGZnbFJ/mMYphbHlFysXHUgQELvQX6Nrs57tEt5xpLmhGn3hFQuHmjIM
tonq3iXsgZmha1JfqxmgVar9DuFqG8vnyDiY8fB3CQVPNzjTMW9kGCabh9uaVmOj
X0Zjoql/jGbm9oxDyeOajiLr3JfYB2igF9xPhnLLwPXvQ9EMGD5eVhcpsw3jw8Dd
VokAJiPqxqBgeUSu6Du3SFVQJ7HR+Tv381YgDJ8fY2q/nZ+K1rHJ8mN1ndgTSbjc
SEgxUrOg4lI6bGmRFHWY71x7sYxF9Qax/g01If8vVNzvfIzXlNso9J25kLb9YZNp
RPHTKH5wkfrs2F4Qo6G606odhly3LqKQ3VsvzLvWvJBOiiwNFvrHYezYsM9HsgqJ
ymNznK3My4naj9KO694EbRSpW9U/hDaETDtR9Ct5ca9FhjzyJsjqXQSqwf66RvGd
5umfcd9cnqNbN6WEZGND3qZ5o7RWmYltIjVg2Y1vN+gp/MFaJujsFZ4tEMtsfJiS
PSfQqsjf8VPdjyTgo/FWBjzIuwJsgDD2G85wXzdN5bwkReFsRm/pPpVXuUziphYQ
riCgpsrQ7X5QBkEiThA8csWTpMwJtUjspenyFHKPercolh2Ul6pOYhq+ZIf16sfs
mxNsdsiIvbtTgD51PRNvhfjZnqMvWv/EahrH14U5IcBZyqQw7IDDCObP5BEBcRvo
4eDNcUpYbv/6GQKTZcLX2cp5oUMrCqzy2jGUrk/0w1m+Jxoya3wgKTwhgOu0Xy4k
oSuxIC0UOHb/WwKdXe1VYMtPwbjVVxDUHYikRpf83Joc0nHkA1ld/KJkpUE9HNq1
dS0A35q8JxG5jqR2//cmJtYgBAULgYwfdoBjmaU+Nwr9az77Bcvmvqip1VFZkpMM
CzZ2um9dRcpkWvSAs4ZlBUARqKXJhbde/a1ndC4frz6rjwc6ImLwcn074FmAQzvg
9ml4oGhzw4OpycZl/AFaBx2AFGuVExWLV17yPEpo17FPlXzy9558NzucDAFKdU6W
PBW8YJpYGflEacFeFLeHI6ND9dImzHZNSn8kX4+s/s4hEVVkHUKtgRBHfiP0pqQU
7SnRooZ2YCXI0MTPPXrz8BHbNZR2QL6QMLs0nZBVhfMLD2BT9dAiRl9G8XSghrx1
VGbL8sqsIvWGonW0msMIDJdkjDrNA90J0gVrd4+MTVJOKklX9r/pxSW+YkUB8Wec
Ipe+JnhUHluQzs1cGelgkxYO84iorOdLdd1bXbuP6FerdEibo/ttWvvEtWSDb5iJ
qYMZ4OUWzmappP3yeB66UzEP2Gco3g3vZyL9mXDZiD2ziQNqRWnELlaHN1p2ZP1i
DssNoTVAjPIvncI8ttpSGUrhiLXbSvD8YD8ossjTYcOIsQ4FLYPalmtTTwdncEfS
YiAVfBIqEKmYpUcEsmavIgdBNfB1HbeqwXINBKdpqj3sEDVyHR9oOJCikGtcET0s
oUyE8DcpypAS1RU0QjTPWuK6HRJv1AeecbTbGWKJxFcxIHzXJIA5esvvRqIy/K6S
n/nWEf6ZWwfZvDauNhhmh17NAlbrPvtRjrrnqsoE0G5KRP50VC3rrvPC5U5RjcH+
uxse8DQmUz7f9CNZK1VRvLGmmA+X9urKR5n3l3J4i/b9e/gerRcDS27B4h+yUAoZ
gBmLYJsBMJd3VhZ9cBCk1446NDXfV8JoUiYm1dJcnurfzFOrVGjiPXXaXHrcYvmQ
L6M3Tpmy5FubsRExPPJchrPsCw0ND9XZySnpurMEXfSIvr/9jfWhDv/jrItEu/mO
8RiBcLKL6pzVZ63dB0YdIIp0T7T/IcPDZbRAlEJdeBPoYKclnZCYpQsPWqbfL6DM
ePmPr0DkivqYKyEZr4SxZ1W/8zTusosMzW7L0XssYsRXfWOazzqN0E0bQNSvr5Ba
0o3hAMeAi4/tMetBbbQkP+mIdHhw7Qu70HAvg4PI7TVDdP/9hlIS9klMnpjVkiiC
OxOb7GFpAwWGvU1C7sqcdd6qFaTq0C0k/F5L1809y47Etfv9d6+yrcnFXcdhJiJS
e5pCEjyNBAaog2tyqD+5M65qVSMPs5Pi7iwVA9kq+bTPb+BlFSiTY2hzafw01K4x
/LJW/LAgp3xgIGwbeym8Zfb+Tpx6u32tUu7aN/uKlDnnkli2Gq79ob2jrC+1JN/I
EgVJpOMILR+wUaCPg6DG47lPyonS3yrDq43m8ZdzdwULlf8adXaK0mfQfChtZ/Ql
45bsTPZcap3pM68vj12lcMuCM/8obXw3B3NillsxANXLsrDcwkZSt1HGktbTTIc8
8lJpY1LJ0deOY4NF1J9Nipy+lqHapFQWvRlatMjHxl0+9pUkg0ekWHrGyxO7K3Ts
/ddqR25d796GIdu6rEnVPw92J1bpvhR1Sjl4a4pEphsrp+CG/Kf7MG5sdcaSI47z
Ekcp2kWXUJ3cpa14Gqk8J2Q7sbajTYHF9ZFSakp4+D/fyVB3FZYSPHP7vnvYMMGV
H2qcNj+jlIPqiFETjn53T0f+JWKikJ2vcrnDKTuqT7+k/AKmxiJMpE6RpkCFwJPp
xarwoLR58E4xFVsprIUmmxeEmgS49/2OEXARkgnL7fwow3pfrn7M3/2m+ElYYra5
XWUAVSQ157w/JfAKUz+IMnGZPByD2dmcHZ4oTX2f9wb0YO2Jd3xM2fHol3LztOhB
4Xms5NvXJq6MeDBdMX7tU8/UOHoE8DGLYUENkWFt+F4lch7nuoRFHiLRHiDpUh9G
KLK7IJSMjmFXaRTLkdqcrqZ5mCW+KEAcIiJCem5m0+rLWxF9zz9KWrwM5A/FLbNw
bqz1njOeKwuOVlsmTvFuO8ABhFj7s72Nxw7phcDMFF8xmu8tMH2qB9PHBVGx8r9/
4sX63RlOapMvVS7WgGmW25XK3N+UqrURkUtRR9XMH+WSEWPKuKdKur068t3Bsp2A
MflqeQDHQnFOATcfuPArpuABzh1ayLRPSB+e96eV7F5aLWN2r+/9lQJ62GwcIhT5
AlrhvzA0EbxUlBdYIBrVbOsL3BdWZ1b+v2U4JrOK0+a+KqhwjoFETLlZR1mWxZNu
hEm7XOPhEg0uwzEPoFbsQwryo6JiLBeMOVLyoId3kE+pVLcZqvUR2EjvKbxC9t14
2/4MOnOFeM2sk0rOw+PnIatVExCOvd0iH5YQbQcIrWZsLWcV7XJvVqqZKemw+yfN
MD2SQLNkhGlXkmFCpvKWH4y+K2IrU6AI1FA1VzumCR6evRI+cTT1hXjs6u59v6RB
C62eW399sN1rlyyvtE+7eajILvnEo1venakJJLmZ6of3A5hg2xctzJnXoXUxmkFX
ebzDWP12wy2zwygbSup63f4PeLOK9QWg6idotQZuCP8LXEU6G+uhcR8hh7iNPxHF
Nkw+FiVzXKABIpVKkn4cGmtiWMZDLXt2kMmewpWvfP0Bte19kqs/kKNSy7K99PpT
EBrw0gRvOkmVHBp+RJijsSl+39lJ64zPVmy5CAsjnXEH97msfjAIr5Jzqg6ymKmb
mZOsSlju1gTvn2obDriwPx+sAVX/1IlE17eAU4lDBHo6kLpX2IQxALdDfwIA9Zy+
fsa3F+WW+TVCXx6yNmq39OZI/nlYcm1BC5H78Cf2ZWRUBmiTs9BXUnZthQIibCri
E/yB1T0dvoj8R5ZfQvtIrtRR1sqUeQG4JXffXwFlzKdtzSESOjfL5+RgISHQwgs/
vg4wCsefLqAq3Ztm897Q7JDBnButf73JnZyZ5JsL5wsZgbwpNk2i2viYc+1qKnd4
KWqnqpN0/+uD3qNnUyghSIN6t+ZRJ8uKJ/ZzHftKewQZKO7/SeM4Dh2de9TAMK0p
Pe4QuodCr8rvdd6DXS9EpaCUhA1NzV3nwz4sZwNjwOnsI/PKa3Xuzhhl6CSOzGXS
DHebuLg6Fh+xnOJG6/mP2gIkHVXa104OevzZn3RmH8FpkHbq4ftA9bKfx48ENP7e
X4D5OBnYfCttf01eE1UngDEEtb0Pv7qr4f/IGrOvBz6tE9eD2Bj9Vf2ru2SdMs0I
cYCwSsWKiFv5gZWbeaXVp3mjHMsF3frgugkdGMtBJjeMsf5lFEBvnXHB9ZUMAZTr
Rn1AGIc8yApD4bcqWeSnv9pvhflfM24gsFhYwe+3ttK2tjuU92LYXuQOJVJHZBtS
5b9hh+lNRKt1Ouu3k9XSmgseM8g9if1mzffvKwC7dHTXt/9NotcnrXNNuAM2xUXY
OhMV3K22BUFRtEq3CEzH7BZ7zjeUDphItUUSpQl++rykerZOaaQ+uClX/Sx+dNUt
f2hVv6yIJVTpbEoyUDjYjS0a4ClWi3ehihRq/vBkadcIl3CGQs+VUEsMOoi16aJr
5LU/Qd+Ha7e6AtbKFheFFgzIEdqZEB2hTWZ2qK92xOGm/r3yGIgMSBkRhlcY1BzX
L4BVHcG3xFZIy6eDCHEDN6UDcxqoraDZDHjnunGU09+7x0aK4SXLaWd39EUmZtmr
V5YjOImqMMrenkn4CGJHhQ5GkVJ32s7jyoVw/pM4JQKxSyjWk8ZX+stDTv1KWc9W
1JWvYxEQk53pneu6oGM2WxUMaUredU4Mu0BFwsofxtwqCx2VnGZqwto8DgFD6td9
/gBB3saZACuONndOWiciZYBZ1Zbhn7MNJJ+Bt45X2mX/Fb82To40fPQ95QgycAld
RpryyKp9qQ0PregaOAiYZFgnHHYeO0TtBm6m3RgwosakbRyop+bwNng/fhJeaoa0
bAY/rSclETU2HtOPObatQlmqHcWkzq07ofwrvFd8b9kXIc90PqRJrTr7tjDWm342
tkKBU1lyqjlGpRNow8mpSRerl3HptRpkE/KEMYcxV8MymfJutgUcB7rFVuVEPT+x
9Az9CLtm78obLX9rlhUULPr0BjztILYhVQ1nnuTjFxzBWkN8YNReE+g0hoUOTPcK
zXlda0NubFd2SZukYu0HZXtUH8lz8VAn7XiNzV7DY4fBa9+ki1/NjYkT7Jg4LruD
MV2pFVTxJeaiWk4LuHNESKiUOzOPjqrVZEnZY7Ps19uRNMthaY+d9YZjqgVzJ4lX
dQKb5+b5xhTRG0CfoNpjBhSzMWqEQBpzhdGpu6A/r521eRrWAmMJeSIo1509Fp3y
5wmgxP4NXXIKXKPw+SsrRHRM72/GIJOFRqkjRR8eFBkZBxhQx9hQrD7HnQHOx+I4
LqzhTKUBBhzsL82YAsuk5B4j7ClZoiaICuEvJirpij20D4JyYUdywaN37n3PweaD
C7yWCIU/EewSdZfEfmcLf0tMzGak4gJPBlRGdyNPAinnX6T2LflhSWUBrprrrz6D
yn06HMFxW510NgaPZJY07nHDKE9IioWDb0TILWuR4F/c9yEZrbaQzvAAR3wEGUQZ
ELmf9nvz1Pqki0PHOvECXcM4CosWn5IVsisLQK4jwEH6vs+f73zm/HcNpI6Zzuhx
stjLvPTFLDMz7lxtA+uFgOFiZbUVnhWQEmH35OngU6OThmcSkZdPB1MsRrTyP0ZA
lVU4mofinifXcp7jcrIX9EFJdmLlcxPg08Ma0XBLeVgUTwvoWMnuBY6bmkK2De5j
5QMgPgIh3kENA9FnJuKWzRZObgzPsV4NvzWf7R1gyToAmjf4AFp2datsOW/GLv8S
pQO8NDPcJ7QAcdPX07UcDO2Co/eDGr1BG4DXJDvzbf++7/EuCeu3D11nuQerx1VA
F+qBnRXLz/wXmamdGDAteTuvLhVUkyR/mTLK4ctgGrixMP1Y6pBCxmQbk/nfgMkK
Qu8B8f/raFFOjbOEOKK6havDkeGqVCVxC4z12innfQcW+M6fPvAI5w90LhdFP19J
pCiwBGlUyWshu9xE0l6RGslQhInUFV6RSSEYgW4BcIpkc1ig28uGBGeYbZ+p5kuL
txtYRQazfQNp13b/V5DQ/Flh78eZJxkOI87GCMiFlbGGopM0Hd9Eb4p7Mg4wkzIC
LGcWdn67gNDRBhomnavkMDs5TEXJiKzjfFAiS0S4NkPTCprmDdqwIgfO/3ndDuFa
0zyBuwc5h1ShTVjCugD01qIZDm7mqUQ81GacTEFnIMiBt4tK2FBy4Mo1aEcqQ+W4
kgBTOyiZ6Q9WKJGJa2whwEHPj+s0cXS8rZWIwc/Ak5tNpk7JChjJrJUma8vhnk92
GDTChPxMsGr4Fc5kvNfeEfvI1BHcEeHtRBa/rc3CQsSvJ9Vour5T9/K71C0dWJKF
xUVpFmeRzsNQU8/PIW+YX+9KVmM6to84NJzJCwqujM/vSQA5b3Tid6fV/Cj1Qa0v
UrwcXxFoKp2rmmBZAUGzQahsjKXegMaYsd3uf2YuRTu0JhLyco0VwsV580u2Z+B9
KO3hyfr7h+AhN8PT93RiclMqlQSn4n2ZPPUF+qFQ6VEkWwRXIfjB+QNoaBIfHpfY
X8osd7L3+uicWXJbdE3p0W1nxBtAXNn86gpRnF0RejIpxNVYwb+p/Prg0+vVy/zo
Cbm6ag6e0BwIDE9y5K+Vq/RosIkd/Ox+CI/QZq606QMa8RNvnIg2M5c6mXOsf3IH
9cz58NypZ8Wo+vu+LCWdssYOxlZQk8Er/S+1EaXikvrOgyYzm7Q1dLMwSEMQ6xzB
mZkOaw/rMgDSG8KBjZYz2NU4kU4rObB0R7vANjT8EdbqW87u7F4xgfGpWoCtOSVc
uJhFMKarzM6Fsg/LkYclZqRhH1AbrP40YuhzrytmOnKxvpBQfzEMLoX/6x+QtIGn
w42Nh3Vwsqf2JZb0XeRmKSfEfDQ0n6jIJ00ebe+N2lHjcFPmdS/5VIFVw0C4bHVZ
zo98V8+lxyEKmWKlqS1TSntl5xXHKNBQaZmrBT96q8J+2MNepQi2CKUcfjDjWDmc
pQJJ+z/yMG3EeZGC762LzNm0qt8tM4X3of+9lAKL3lNNKqulOzM4AGMJSuyHeBkV
TECiaR7jYtQRjC/aDqulA6rLiq+h8oxVE666KwNHLTi2YLF7AwZVRDXsav3FWmtV
nXvR9ipdnIv+1axrrDKPHspCZkZTtw6cJdA9Gr/Dw95nPBE8dLTuyEYcWxJBVs4P
GogfTSsCA22etcrO6jarfEP+3MOLaTTeH2e2QThIUXl004hl8N+z+DHLGK18qks6
mDzQvwhdi7Id5oY0jgbPv4oc93pCNl4CPwGNZ48hmXHPYWLr1IAUyxaWkHfNjQhc
41wCshgiyJwsKJUi+dpwr0g6YsXdTKSjSqzmLViorxi+Kp5Wff6PxEhrL/28zons
DZeSABape68ega43txezK2OhEpYYbwqJbW6D3Hrw3+it7+hAm55wD+vERYNCI6MG
TDMHIOg9j4c6SP+i/BwtVodPDJM8Z2hhQkKtyI+fZAbU7ifKZ2XjSxsS4kK7Cl+T
R78lparvBbFEPz5pdFy6pml7LcH9OE1sLNreeOXsObdYNrj754kl0M0dZAbUdvc1
Myo+9w27Scir0I3M+ErvV/PAOaXVUQksl6E+i9p/XzERZyUo5WnxYkXZMWwnUFAr
0PWQOcJzDRw1cypSGW9muBWRcF4PQSdpdaatWB6+sVbxUKPeuvU7M4leWoRWdCfo
VqbebuKspKJRDHXjdsqXlsOVFcRachDsYzgkNofTibOzlWKLar9vKrrfxb8Zsgvi
6Ow1LBzVZCElb5SRAhpxUnD7bDDBLUfLWZReWFlnL0M4JNO/WY1d0ff/rIATvhq1
LskJJn/6+GIVhRYebvCFqi7iNL5x15rL4t6YlrtFZBFDRvET4XZz+QjLQeC48P1R
GHRGzhmaaC9wxLZNUbgzvazVof+kt9MVkXYcQqR5s+kTDMMJLFEIjiQV0zCa8dly
HSNMfsVV20wuYKVXDWdQ1LBKmgoojGBywF2L8lW/IfZf3eOB7KDl4niEHnxaTt5X
pfBGd4kyWVRXGHomrXK2Hd5b2a4ISeWGfTvP1pALZXXDpuiXMl7ZDsaLwOGCvKtY
vnDwQuT6Rf/05bHH9/UHTBl1+r3x3bd3TrtdWEz0qY1BJ0eH8F3Hz3FqKwG++kHe
5Bjt7YW2LhGQbWJC7ndnqw15y66PcvehFTFhUZRfwd/KBkAaTcA6OXOkOCh0lBwI
jFwySjPAYXV4h9WUkpsgGcxjnUUuDQsMWRRAAi+4lr/KE1Sl2li80oSveNB8hwA2
035Bo9nAYRgJMjMT6zCmmA3AN18s9Hbs0/rwZIaRs6QYUpK/gVpaq1Eqh1xPElM3
8aG3waKYkJPBp8oIrtnmqEa2KLQo/GBYCT4S3TAKgoFcoOuVdZ+mF6L0S/IR/ELk
i8+d6MuYnYj5E9zS8QyQuMI7AcdokZtaJsRGU8G7JgBDrswpOATcuGBxkwfrAEuI
98S/VvQTFb+GYGOGWQol0r9Rl/uAVVPx/fJdhtdVfN9U2ON6r5RkLmbH2AKAaBG2
AUBEq7cBgxPaEn5LJbGSiTEbPnjN1J8jgZalCmJY8cpxnKooPZAflwC6iExmfWcO
aeTZBZqiFVaVTz50jF/UMsqfgJzLoi6kt33Zjj0zEeUWXMkAafHvTGIRs6lZNQye
YnTSdvrh7lUweb1HLJdWawQ2ijR5BHJG7E8rN1vhgAaWLB67pkr6lsTTghxSGbiq
sJclBSn+nCd5yHC/e6JCSz0bEt9g6DEIlsen1Kc2GhAZSW5cfC0+O/If6Mf9y9jV
/Wgr+/7PjP4HxHHsd+/vUvovmIcIGxSJgGQOxy6tyU5c6j7fgRJjJRK/TaNwL7uM
DZsoHjs454LXmJfr14YQ+GwtjktrQbxpZFO0dUGVivTwpCjk7eob0+kqSwCPGyWh
NZz4MdqCr/dqUog/OdWXcD/GAn5dD65NZxyaGTzbc/Lahyb8gCnlFLiA8lLowCGz
dPy8nD2hGNVjiVcCjoRXi3G4E02gzhlgSQSmLNu+VN1pLb0rAVqQO/uTtN/k99tS
8FjpDd5PgrQQy4zT15yo15zty7fKhKBuC5hPQcPODf9kF+EzokEQYjeXirT9xFxK
HHmTAoz8GKHT+Lm7uo6+r3wBfE4HUEQs45/PlushyEGqdH7fUu1UCLR48CB4D6kv
+EPmjIkbuQYL9o7Ik7uq70It5cN4KYJ3zRxkNwuOBVLj8z0i1RrPzx/f9XlYzW8C
Iift5moSW3x+LtxAxJGFyKc4Xpkyc1opWkgH0mtwHUIpkksXwSguf7XkFLiAnxzt
0jz4iC44OjzC6zCdbR8W5FPgV2ZHbQbEgPBUaVbin86WMU7GJs5IDzr8l9OjZ5jw
RCvkb3iStfssDVt01linwmUXAVqKfGDgYCw2MW0HVmHQl9nUV/6hqSf2zNC62oPX
1aZ9rmnx8UBE9qW3Ww3HsXmActqcq6tvURWKjNKWUubQ5a8wjMhdql3R1trmQteO
mwrpHlKhaa95SXfwCmm23MrpZejgPQbDhdU2sJM/tp27Fdvk+KTdELLpwBLSHl/L
jHKvvtqvvl3rc4OHHiFNezb3y5SpNPyfZG5PwrgYdWbgPTSskGsxa9Qo4GGwp1r1
WFEMVmyWV/mB5mf7XgjR5wVLiV8ei1W9ZRFCKVivGAdL5I8kvTOh4tT5ie6iacwO
1UQNrUeTWHkHrlypiqCgro2/S23IERSBhaXD9Sh3vBEBi7HG7wdyQG9nX3yI7OB9
60OYdAX3nhf7didnkBTdOLykaq9LIUgICxtWepsImAQI+k5lgJvAqhyV9+/9yS63
AAOUTD+Jzpv9K/7101KrI7pqnbedV85o0NErQ+6n/3mYWPWewBe8iYrW0x5XAu2z
mGsXpXmBbGTMo8D2JOsDFxrTxXZlnfpUXK7zHwMo3f1xPwJmDB5NGuQreWA8kqTE
u4ZSioyV2MWjTHsBttRbhSzgWSC5lUjPT6zB7WK6pmgMocW96N88/P4vLJLhlvTB
Uu1MRA9N1GON0QuEQQ07pytmd0N4jyse+5ZHN7ULqcYqX4rCQuOIY/K+tORzKLnA
BpUnj1TczUvXyD0Xaf7Xr9Lqs/sUOGBmTPtWDOmgPXkVx1wpgxnB0Klpn8JLCgnI
f5tnbokAYaO6wHICElgOQUQX+nNniCHKCBOv6MJswOeL3qWSCiK1Jy6d7EHvETej
40WYGAAydghiPE++8YEHw80fy9Q2Hjk+Sftm3CNTOC9KIMZZsD8qQHB6x1iXsWgD
kqU7Pb2BI/ryZ2q2IaVefl4M0Ew6itF00xVQnCyR8xJpg4871lQPvfV+SeSMLTiS
pIAZFaY7oeIk/Iwdd4K2tHU8mT1TXis8w7tPCdHt8LrO8e3XiCXkdcXUvRzUoYLm
vxEOF+9zpPbFGK9JIPPlWASY/syvKvJl988N0zlg+YlCceLRZaqrxdRP4u5x5oJs
kGnapOBOxq44kx7V+4xLhqdfzoPKUJtAZpvDfbSto6vW/B7Af6m/W1Dkyf7Pepll
0x6leN8z2cfdL61K+5Dh5U7TTQQlKS7V3jETL5ZfufTTOL2GjK2G1NvqSQ2Dwhyv
FrGinJcKYgZlRBjFxWpSITuvkCoIT4jzywalOnSB1vmaWHNhkZ0ytm5iaPgA+8HK
cFRf4kRIlsu55nSBvewlY7+JtVyEUDmvbSxXCKX2GM4CMVZ+60C1InfDYaJdl9ip
UCwPH0fha57JRywx1CcmgJOqkusAFsqM+K9Q4XUgxThlctTZ1dKmI367LYtybG2B
bjQqnfBaFdc24IBfhfIMjixWv8x5HdQY3C4SxaM4LStyV8c9xB4fems63eulRdU1
gDMptj6GJIksjcNTif3GIO2KhcyFlvhIErktIkxDqrJkQlwiR1iLr88ygn6UXlGa
XEI+wnkRNW2ngJGmlqDpWSpdgUOGMJMI+pt6Ll4DbWzwmmufDUkJkKLG9fP2E/Lv
hmH9iuik2+BJ/LHqoXUVAIMNs+svdf9CyOs6pTRVd5P64nyG/82/mcZxX6HRE/Gk
Fi9MPMv1hJGyZZcH9d/Cr2amlRG0MrhWGHQXf5XCqFjWKmGe0rJYrw959aYIRMIw
IQzyvZRdGY5SBUTz+mge2to0YD/NYsgwRsqB1GXVMrp9quv5fLTNKUctJxiobniJ
UDDTlD3ZYjeOWyvHoFcu0iIDaF5wUnpy5aolZ//oOp30PhfaujOQZ8FniaWUCVa2
skEsbKLg387uS4ErOc8ACtx/meCGAMST4paDs/PAHvUFDrzL0gfbADbRYY+XeQmk
L3guoCyYd+FlBQyyThWQu9BevpqoE6IM1qIpDMAoBFUYdpfd8y6tde59GWmxaa57
V24bX89HTY2Jl6/C5JqORneeoHlguf4U9nYHskrkcp4atv+QmU9vfMVIS8z0nKUq
rnH2G0EqYe5FWPRugqal6UWpJdk/qI0MPJCPeQ5ec4QUFuihni8ExWoPSEVll9qu
W1oXZroTBD+7tMVqwcO+QaoZvQgzE0U/mwUJMLA0djB3F5hO+jqEHomgmQAakwR6
DFiHXkEjZ/P+tffCXcvyDvNVB3Whk7709jctWgV4m2vPP2ifRVCS+EYcU4jcmhlh
37s8sXvqDt1yRZuzMHWYIscOiyVRT0vknjLNWfJjZBuZKgIcvXjUSP0Vbor92uAs
htCIoXVaGU4jrOK57tmwJx+BANuf28MF2N2LpIzhlc493sY/5UCEg7f1Mf4GR3db
Y1+rQZyknoMgeYjtv7InzCq+UMNP0Gr13EfaKhCRpIKpFiyiYUp6Pgnz6aXX7//o
PDO5J8CS7ILmFjQSP1T98BjngVdQFCahUVcc2nzWpMFiHdhI6Y93FnZP7d010R2z
kdtWFVsqy51Z3jRpouHoES1fGh53tqAMCsu2uWbCrt3hUtatS8c0WARQnhz3KtQ4
7aY2Cy8M7+fNJopklnVCMO6g9G5A800YHlCkMlTHTevoZlMRjQcFPyU+uuX+r7aX
BTWPN2s9OsJRVvvB+pg1/e4vWZiMZf3VMJwqFYpS29x4mog/BwRyOSnIwAXLN7ft
6gbVkXWfmG8HD+vA7NX1O4XdfGlF3FbDFVf7S1CMOmelcz3AewosdDbLgmA0Nhgn
UkdYLuT1iiEAwJROdfGTKmbjDyI5y/n/ndK0tx8sJmCLvPBy9hTWWxeJPMqQoaWI
3rmKQjar+vSTj4bCxi23MVveE7Xh7VBkdrmTEK7wjedPoEBOEiyvL3s5A6QXFILM
2N+Ggso5NtggQi3159iQDBdJs9glKR5GhmMWYBg5HOHoMJT6ZuDGrzpi3tOQ6Jct
9PUWJXOK8WslSWTPamTjXIVJoaMtfdBxMjGiWtRVX1WLthfVsPKvIQyGKJ98W798
F57rYi4nFSDcGftRILMZxhDohbdcLwKAWqafSM3dRYHrsgrU+/8GjcFxBmc/M1Qr
GwOdvI+pZ1ww6pkfN/BRfBI5pS9F2kYZVkSNfz27DQNgk/LM96vUMWhHNJ59hAFg
0L/WqRUB8mgQQ+NZ/g3KRBoiMUupXdTydep8gprKIspUWzlE7Vzo02biCx8QuE/F
2Gtm92UCWw9eEtxfFAv1Lfv8uNFtOTue0b/cEWIY3c1uE/HRTVn8KGWxKBeTXrNz
y+LCMF68PnLRuOvD4S82CrXSfmnfQ03EysJUcODHgmc2GdzRC2CGSp+cGVrii2KH
d30/NZY65Zus9XZ1o8Np+VpdC5Mrf8Uvo3wk9UlbD2VwcU2oadrtWyv8QNhMNj85
ugDJ4BnrI+whsAwUCuVPmhdL7+qyg/d3WId/046O3Z418IUYJW4snZ6gBZq+7hex
WJvD/biiY5X1uwc2GLAry7+DSqgqiQoryRqrJURW/esER1zo21LLWME4hp02dY9D
5ByZ0QiHQBOB4qxmHV/qJhWCZVZvrg2DaV0GmCAZLBPKpSEH2Mvb7n789G3kCtVr
wYGpSPpswVCJP4wDpodRIlm6yGQTFy0GsXeIlSFG9ZmThp7rU8RuC3eVFaTCT1hL
GvPJOeLvoRJ09zWwGdCb1BTfgE106oD5SDI7aL4w1th3oZeNAjMpKc7TTMHc8e1Y
oE8Dyqt4JyLGXuNIRx7PAx/b4onFRK6BhnH4JzJez0oYF8yq/RNIvV4g5b9VQvTD
NBzQIcHIQTXkzcR9ADMO9lWBVphULm8SYK0jCT7snf+TkQ6pmn6uETde7xKkXGXI
iIz8gxbWetpRy27Xnd5SaJkzxqUjLRsB9t/qZykdnj//TZ/aFwUc1xdkhNhRTcd8
wSkmjctyCSpkFFQpZJ5PTopwALiiFFmro/d9+Gmh+GPmc+x+rnxqycf92dS2dKJo
BOIaxSptVGIaH5chxeSiU+s4GoOMB16j/bMLFrjfzXVllA13Qg2HBqcV1BmDLmP1
8/J47WzCtMua7gXiz9lmfgw4AhtxhwH4fnIjpD4Hj1aUe1svqZVVM/VcipTxvz6R
mq7xD+GTbCm5nhhRtMscbQaE/JD8uGE7kfph1zg8CZSCa7pjQiTxLTVIg5uNm4W7
NBCdiMEVnLOcB36Q5FK31wjxWYHPQvPAISHVVlCziLSt3/6NZ2rh+lrVMIPoNAbm
N/t8jUztpHHsiT49ufgLWazhK4nfwdDBWPWtG+fho0NZQve/9KycuBWnSLyv+8GQ
eiEBKDcQDbNRalMWeLbDnLQIcKhepLeJ7uSuIyVlmCooczZz1GzibPXMxE86DvoP
/BpXsW9eui8cbBIVixZcsg/UW1oQlfjLLAt7cvklWwUjo5dxtqnKfBgsoV0XUL6K
l3Kldyvx2URlD37ZkjpJcBg36RQfmevDpee9pZVESWecklyb6vVMCUVai0ojGpHY
39mtGFDPrJIQTUisCjjUrBO4Isbn/mKF6JiRDW+QeBL478CYvGjObqSDOH+0Lf2l
qWNRfIK8y8co5AD7Ie2lExqcsv+9pIJkY3zlGxQ+hP/KGmD+yisEl7wcyBiRoteg
sDxEiIp9RdzrhnruAlsCxchAja3q2w4/uRqD1fN8NlXgDkzCka9arMuv0HVb3lJT
30Wbq2389DwTTAPhtnR/jpOVRGgsxkSUELu4Yxblk9zu7vV9f18DMJ37a84+lXwo
tUJu7pNe0QMuPz/Jfpv41+Cnxd6hqxdNaH54ZvXrpeXB68u5f3Mk+0TevyFbMjoB
to88Wtum0if+Ecv20yE3DiGn+MrUDaxVpigjMmyCc99ZfafJjrjUwDhKMioJk8/5
GfZaQMGeizgFQ+QyaaqV2VuZ3B2hleqWaVk7vF5j4k+cGS7E7FGsELqV5xbUz/jC
g2TiybtfBs8XDXZckT7q4PsB9fk8a7JQQS4Fe90yVRF7YxmS0YeIcwZ1th8Y4/pZ
Va7LguScFXmyBrVfzAOLBPYlVeDyaobVX5Il76pISdTZAaXmo4L/TQyvyAgJ3EIs
WZjuD3P2KlZ4KZU7CdzaksGv+jZ8EoZ/IMdaW/nGds5pkG3nAP40foT808LprmMY
Chw5IvtBaovHXqvQfR66DZ+FGmkVcEGJA1yfsfwH1Q2bUMPM7p0JymGdf/cpdlqR
xSmwsn7A4CF34IG2GkJ04GnCr/z48foARde8yK31tqlAQNRgPrWV2hnPc7JL/peb
Y131mPs5+j/PhMOflG5vcgzX+WAGwr6qWVvv+I6SjVOK1gTs352ikIpKE49PY1rJ
wtanXxUxF88hMVAp42iryUJIaBqzH8tbVeVri3RID0I1nRjO7PWEimRaB4nIY7ns
TtOEOvzHokBdfpFUrjAzMetD8ItrU5akWkTINELJMVd1ApFSancKZYT3x3Wa1xgh
27rPchirreCJHlXvw+9sE8teE1rlwo7ZheIRnPR2+5FMFUSws153HFSuA4sjrkr5
UCkla2sQlG4dI06ntyPf5D1gAN+Jj45rdUH0/bYwK1wM8IkGyuBKRjLsfCrnrTKB
si5OPb34t8cg23OzXD7lmyQ4T7S4g1WSbE/DL2kSivd0p6hClysLgqdGGdwSWCe7
7jELLTqOX1GvWEY7OlY5uTfIdRfrUlEHS5AkoK54CL/hc9GXq29uhojf7hGPRNwY
NnMQ90w0U1x0kPCzUgfbih7STLFIz+MxAZepCMnnRpmy8NZ3Q7R0kKv+wPsDRKfZ
aKs+0qMeT4rkL5sHOCSYv2oVSWELMwGS14w7B5I8a9xfd213cBkL7sKPHXMyWYNB
+9rq8XL4nvonfz+l4GZ/N6zvLhXwbJirVJRLjcFrNfeOI39HnECtBZDOCXPQYMwN
5wsTh/q8484+w+GDrFoA98WM/XeS+irdqpCF0UGWoMTtFAw2mT3afeYWUz8Ra0tU
0vMDlTFKRVMp5mPMVXRlU59jI5q7kTaYLSYV6RcY8SdlsdkKJNsTT84tFaX/Y+5j
GZGlIslz8jLX5KkZ2FcrntC1UJ0SNw43+cdk+c428niMFCzRUYeOg1QXCb0DpQZK
6zMKdNUh6esy0OjTSAp2X4H1KWqjDn8nuADUyr0ETzHCwBj45ZJ41ZE2/vNfMCSb
FI/wawx3olBXuuParnpvXqvDLNwf1xJt6+1Azw4nODgZQp7db7j3M08cavQnInjg
i7XHe1XtXDFT9E4Ax9zk0wVLfr1ryEYlY5qsP9ugvBHO6Myo0nYZ4gZ+1anTOAe/
NEWtxGZOy7P2sf8/ZzxrubrIu4GGbUgwzar3/xT91l90su/FGWDKFVddG5Vf+5Kf
xkXM+0EfPrg3due507X5FR7mArFJa3o1C5ettjvGTuPyh9/DDhmfHNF/t5km6WPn
vkgOkrshnnqL8tTUpyg0YjZs+sOSOZ57iWT/gcWK+zftjpk1VCuf4TqBIesf8AOx
MXZEs7jnVFmTUScBeDMMPXyOOh23+G28znU2I0eW5PaZi0jHXovXDvLyhtv8gKFs
PqObliy2WApdEP2XmXLgF5o3/W4t9uwrHJ1Z8Q5PlrTdXJ4Wq3nM8aO31nDe7VLJ
NSDDun3maPUqWw2D/WTAZXLZgkdzDkHNIM7aCls04qcmMLOf+nDlzqONLX1/EL+n
MycO3NVHv6xKcvOQpMiT1kx+0XVSxGY1gEJ0ZpF5VJtQeVfZ0DzbtD624i0fUSCH
5kaULhbudtSs2RYFg1mqM2fDCDcmIAboGjIDM+wooRgCgX+LP5P2OrXRz88Jvy+Q
oMszxFLmXGuAlCU8BIdTOplYJZrB3Ik/4bcVWb5TQHGf2QA5qWalGHTxkaYweCK8
G9qKujkNRfXI3XZ/lS/L6RGdCANgiRFwgqlPYQx7rZooFgdnTJN26sqKK+DQugES
MOfg0fzQUyFxWCU4JKJ3h+n62L1jnLzT7maGr06SCdZd0oe4HGwPWkn7o6N/C1hG
Iqiy90tCcTP/KFmuE69ORxHtCID4iKZwZu1vHUrvDZhBsdPSrJ1BKew7a/pBDCRJ
254ZOe0djJ8QYamiR8EVZ/YbBp5/PKaUwnvyGxfBcWwrKvzgLDGyk8YjKFekr+Yv
r8xeDOy6GhSe1aEnCK3GJBsEDic7dq7Mb6jT6aclZSNMaL8ffbmXcnQNJP2BNhKC
YAFZe6Kk/N/y0teNRGKThZjGLYWy1B7e6kVEoiXvP8cEiMnA1p2LORonJDfzeZM5
dLIIiN+2A+uGIobPxjziVjPufr81X1NzEVhmo3pcrc431w6wOlq9nt0TzA8ivpe0
ovWJbjnoSGFQCUSEoQ4fcJrFh+7M2sYGYEAgAFn1jvjb0PNpNWof8aoY2eZ1iYY+
g0yDfQZacS+FxV7dvtRiMq9pcT1fQyGq9QH2OvZxgcT/nZfUm7fc2NORXfjnOWDN
2TVes59LOYduSInLvHQeAb5QdnTn7CZaCdsRwEX7oAyFhqPJ8j8LX28DRI90fl0C
JGI+9Sd5AGEeixQwMplxb/n47BTCVu2uZkK9FjoQSTgsC1etDaT9yCFddvJ55CQu
kZU+WOh7MCbCedoeoK9nFKk3NLB2TCM4IkU0chf1mbx3Ym4w19L/MfCOcmv/D3Bi
1i9C3AGh1lXMb8LtvvQx3ssnfkzGJK39y2RQ29HpE+SPrX8w9l5G9aWrbryT+Nmn
tMPaYtcWicdLdZVzYzOn8RvyiZSXszTtc43rVhqj4gh4lFDlRrLcoSgFSRVXLcTK
Ip99flztLy4Agy5+P+ulxC71zm84wm33cehv3PFZrw3kFAYrHizMEVbMQgHUTco0
j9FqAhXxoXJaKmDTnm2k5Vke2GNa25D4P0TC9qDxfnwQPAoqDD5UyFJ7Oyy0eVA4
dz3OcYnAqgvIaX/T7vIaS7dwSniNVYAb2kAU6HkH1503muubEbKW+cR+5zIyTs2Y
FtNSYLgBlmfczP4e92vSuTIuMpPp+p0Niu4RvX9Rkxha2+2+VaQGhd16YVvpqNOr
Qep/jcsdhRKDKoswiVmhMGhfiqmrZcUFDLe4vBBIdomw96f2pGzeso4GvaSz29S7
sxIVu4EKaz+SVBDzNegvKl+1jQx97yOH84plg83E5rInvAqSv0BK+Y+lVqUles1t
riZmAyLm12IZZthcfAz+K1BFnaVQbD8izbKBp1JBP8oTssumhcNVFe5ipDZU46oT
d+/DS6JPGjXOPunnL3oZJ4tQaPeTqyh22tHMxOGy7FEmkgbcRJJm8DKe7UpQkCQc
jR4oiUGhLO6zm9oZyv+KaEy48wAXh4VOqxOiLvCUXqnXUqHGo2kIuGgUlEpBWhb9
d+JEVI2fdoEyDdCUFT/iEghdQDQe2gpMNGQ44ED3J/8wHq/NZPFwxRZrqD7GSdJp
TbunXVZxto0u/BM0oaksFeO44OR0I/8uOnYFVl3coP9nB8vks/k42vOCqvHTzGXV
s0q7M6GElUUBRlj9iGHY3J2HG6SboBymLYFKLf0Go2OC3SVX98DtoOX1+hynv9Dj
Lrpm3HP9D8Qft0KAFEvwY/p+5J7YiWKw5lXvHd7M6n6mAazjxiSnPmiLKOEp8gUp
gGtXFUWth8SIuQ3EaUpWSVtlxxQDJeqT22x8st5yaKmfypAlikZLML+giskihVbL
9E5t1bEe/8TPyLRymjLF/uzJYdfDHJ4Ipb58DKdytgieRJeKyeQ9rQSry5q7EQi1
naSeyrkuUVRpF2HX2CYwj8GXupzv9ne2Isynj9NvFm4pIHTivHqYClrYbAIELDf7
HdZZV9A8M+kyN3Yn1t7coRq04vJqe2mNLcA8S+f1TYUoZz1+DphNKGxvLtXyjal9
SZT+++3Tfn7NQNU+Fh3vE0ompGE152LcJELgtvdO5g+pRiZbLAqcDYeFimaolRgl
he76/3mOhKs9PwDk6r8j7fysTXBhlOc4BjgsUzwsq5GfwWYL/b5kazzQc4kb5v5+
IYqqLfZcSa3w3CuI3wy+mksBFNkbLhwl6Y72z1TdY24HMk8BHsf0IaB6aLvmJ+ZL
X5n4FIXEr1VXzZDnrhjDckuXj/pz3j/kVUaCUa4HiqXFyc3u6e7W6WGaKWMi+Epc
1pl1Mj2vVYmEfwiG5r/BKFVVSu9hnyoHZkqMib+WyeMjI9sG9kO8KN6GuWSq/BOn
raO2lUUlBmeI9Uoz+62EfG3stFkuqBdDU0EdjBSzTRQ3ALFF6X/8bMQZs++Z32Wb
Dul4/Fx+OktKcMZY3G07bRAINJ+V+HTu/8H9q8w6ggQwElCLlzil+TYeyKxjL3BV
CfPakEow/Jmy1/Ks757AO5ohIp1PYcJ8VX9OOSvSOzE5v2rf7k40SS66or37T4mQ
NdRhVGNESQ4vAAgonlhFxqBmEhqsbrRfBHDwFIcTy5E+XIhDoF2/qsK2j15RQoo8
KGf2xJBEZqeeV9V9ELtwWFQ7JDJ1yfnj+50TThuaCZyKFdPv8H3kdrqe+52RYigx
akgrnHcaIov+FGlNZqqvMvVye3iWn5UvaQujKstxRund7StNFB4xCy6TO1h8lEqI
7QEX3Yfum1T62CEo+EHpPDzWh8PQOeM3w6NWu9n2vZKBlfllicxynKevK+URnXNY
m+QDB1HloU4B3ZThQ3uMRjb6f2orKIwv1WLSyocnRztsT0aAReJ2PNoRk5DCt6AK
GjFQdC7DP5TEXwut8/JZife+2NPZGaq3/5H3i18+jiVCJUNjMTF9BB5SUT9cXm6V
q2q06ALtIgID9kDBZlEfWGeQqKk2eRcMzzvp80eUw1vHr/0EhuiuYmTZOoV7nMMd
T+k43XfrvVMnHY+QYLf9V6QsNumYH/mbVIz8jvAcMqMyl4xPn6QcFUS06nzky0Jn
Atct3TFDZFcULOfYWRH+caesvp8dxCotEQlY2pCtpSYhnroC74488mY9wl7OXL9S
v4OtrbKpCgj8k5IHpKCDnOnYathI6PJfy1ex1npmpsukVU6Z+Nrp9fuKS3bnziT2
sE8k+mxk2fxIIGSmcY709CPbB6Oq0i8+5yP9LUitxPdo2Rn2gchF4gTesY4Mpq/o
rBJBdfNqXk0NoTal79jwNfocOomveWfeiydnK/euLbGE9AP9QWVbJqOcCNxPD8Dh
mdAjK72pTCPuobOd2Vl4KC6ehWjNn1/T1HfrvcZexAQETdSH7uKcXISnKybiSY5Z
rsPCbxl7/XhXS1n2yxDJk682t7oKL7XZjL0NbYIFi+DtAwlohM+L/Den3qelO6dx
57U0jitquO4lyFfnEG0PKKGSiGpmta7xxLeyaEcI3YLtmZD3eu6+802dQcin0vNm
uPa7lKJmBa+HqAra9CFYUWiaxoOk9bwSzzofBU67zdf2vXpx+UEpRIdQ1bHRplp+
1ojilNQ5dZ4S4plPzxN2E/KZ4pFe0S13pJ7/EJX9XQ/8iv8/1klTniyIGTaykR8W
C745nFJsg6kH7+aeUD0ZnuwXK6JY0ZA/D5yVMeK7oXLryq3fCUnsIyiqgO+gqnpy
rpK8DYkJ0ysde+C3216ovEbv9y+4xKheXrBIRjZjM+QTLT3UGOBaP5Av2zMC1nat
5XSVmWRTd09jyREHjhueOEk+mM5WXOzpcmiSJIRxGdXzMPwd07cwpAbc2F45IXvo
tOEKRd8o79rxSXMZPwQel5eaenCxHYfPErWyOKagevDqd+x6EmmSOZdZ7RiUnnL1
yS3QWlwI6GdRHEQlHUmEcU8278rCF9tWqQ3GJUH2pbi5C8g996Tzr1epJhf3d3Rm
BWrR4/53/R8OtUkGye/UIMh74B8TAOkaO9G3YeIoRMT4xY1SbHLKhyA+NJeWg5SV
w2Wkombx3SybAsWJTYXPFk6wHJGgbCLpB3LbE34nSeM3yRItco/DzZ7ezNvdGVQy
/M0J9EUuCjX0Post20p4dkpMkWnmesHlVznly40c7xJkITl3qjacBGavthrIZPzc
MqhMyttHztmUiJiEZBZty4e7+rNzlAmxuP674erhuCi7hZKEqwm1sPkRK0S/X+Wu
hNIqfxvSt1mlZ2XhltSnGFwIYHEJpbl6B86pxu1BFLMgoiKsxJy/s/SpsR19qpAX
16rXOSomygEw6XB0qpyLuNMg7nzli1Ooz4yvSjPCuscqx876npgVsfmZ4cEo6Zor
ueQS6/wp74g2fJzE7YPXkZyNqvQvh+63qPpnYBxyq+BR9x9l8BKlzwfKLSEDzd36
6JdKet51eVM32NEcmojThEWBNmo8cgj8ZlkFIvCINR8DejKqmzjud0r5LQ8Ifr79
my4MQSvmwTXPefgdSHjDNDb8Fil5Wfa1LSghGo57KN7ZFDHMcpzB5jG5T51ZmLDj
134Vv+W4CBcQdTmy+Mki007csCo5t6JJpd5N5HcuclNWs1i7glrIXepaRghUB3uK
RPdk9K9C/DvKZ23azJIcvz1fhaHgf24DMDxMAsA+lNHP/xofmJ1KYFuSE2MxT/We
eTuPxC1Wacxz/vCvhH11T7nAHcRPeku6NV7qanzlr/Wu8J2NVi7P79cS4VpS5ig0
f9TRJpfu76yCwIxqbpbIY+UM2l99zGRM74dM2BXey82joBpH1QvW5ytplHGs0Moy
9gK/g69fe3bk9txKJfi20puDpJXyOhOPnCiZeI85wvACZ7y6GjwBLsP+JO2kBY2b
yoh57C8AyWBLQ0PAANiTQr6/5E1MikD70eg9QcPPYRamks3RCDptxfRLYGkkgA0C
FBc3ZcIF1xV6YvYl1yILKUYwVHTV0KeH55sBEML53A8TUtqphdg5BTUCfJnWHig8
91FyGkxH6fWqlzc93OcJQRvnKbrC9wkX/gP7mq7cvtxZZFaW1ebqahxhMHQpCtRJ
YwKXJemSUI6cAT21uGzXZhFyBmP3K18FTyqiOnBY8P82ZJDSLmA7us/z5kv2+sCe
P1QlCszzWalJOOkDLHShVUfaAEVZ0sCaxT0aivrCWTyQdQ1AAAn9N7uMgiIoAXda
NHMrAF76/krZtSveHcOqc98GK3wXyXOagDorIl8Uo1NqmDSFT12GpdfDsY1i92Sd
ZJZHkW3nH5/lHyPkIZcL0K0eYwFNAD3xwqucq0AmcECldZf5aoDWnreQNfY/LqPe
yO0z4kyqDjT7aBgPphvQ53xY3B9mSC/HQMNUFRP03mzpf5vbii3jWoXR23Lw7GOR
fyuSiBohwS529U7irOti9v2PWYz6nqVIw0OZphIX6ZnZy9ZZ2M5h+SE5fb+OSWox
zsQiNjB6IvJam26sxN8jJ7mzzsPyh2YfDwBXm1pOn5l0vX6O7PTZlvR1LSeMaEuP
7wK/Sl9GwbWL6gQKOF4EgTX+hByT2Td3QO+B2frYPuMRYVNNLpqJ1pf40d0IsY1k
8dzm6hiRHmT6EcjT83/hWfUfZW00zm2ADW4eBn2mozFzJfpiiSOn8MzVd17WCuXv
ULEfr4P/dEOcVQhAd7E/qfc83HYN2+1vPFNKayZ2M72ESY38FSE1glbJOnd91bEs
czZs/W9w8MtTyUmpSUmCSwvji1o0vL1He/aUkgW39/y//knM4TPAzvO0o194Q+qt
N/C7tmwWfSs8uPhBIu0kt60Xb9CQxNKR8VBpAWyuN4LghDKLXBWIFtDqEEb1pfGc
4GNgy4kd7aLy2yKtpBHCiN5RgEIX06THz4aGwPFfdwwnkoHlrwjja+b04SzdO5fM
0etaDZXDqi8m4DTLdcCTIqdebYMnojikOb0j/Tw4jfKTt13znSPLr+rhE0/g3iqw
J1QS2hWIr9H1HjFCOL9WNOXYhrkaCAIpNqoZhRen+3891PFqbMiQAt81oOpHGF7m
6ofrHBAYJLXCfAtuyH4vBT6+oYXfQ1B1SkNGDVoE8XOHg4yVk1HJKaEvUlmbra51
orgGROaB9B/9VLfmK4wIcZiiCLXQswggyURMKztSXZ4TWCe7Cq3fR4zpAQWaXIei
cuVEdHZSXUTWYMP5tuRoiu2KFaSKJ1gjb53hBbm88rmvmUnFZ1bz/myM9MihvOa4
iS7N0wkFs60Aj8AqekM/+uwrphn4SQGk5B9iuZnESpOiLfH0JChUKcrczr6d0l60
bpL0V0Wh+6KXkdaj/IEEu1Lki0BUG1aDi1VEwCwVI12yK/PtjpiUsPnzOmWgpoFU
xGXttS1L0Vosuqb4Ps+1IaDjBXN6yMpzP2Rd68ZyV/0ER0gdlMC0DyMM5lrNP/SX
RPl9oJATsgq/UOuXuEZThbs4GVNCzp580MoDOxO5DJwscs0Hd4siTDF2SjFB1ZrU
WeJ1HcIyhNtwhLu1yd3VvdrCHyMNnlUbDBxusChwD0RIjb3VPCD79MU/7x1hIWqW
X7yvGP9hh+fGLmmN7xzGSVl+E0RvjuKIr8rpR5BfRfwO+1weUfyOCKi2nJTToZ6J
U8IBx32bkCc9g2DZM8UnAiXN1WyamuQIzYqnt9ada1Y4E+TgaMsCcEIqoLCSxuEa
S91UZuWfdh38qg5X+9rejph3RrypsNvcV/iP8Zqv7fJHEOCw3iXhZIE3rkzO0WLx
RRhiGLnftmEVzV+UdOmhqrC8zU6lff2+BKYgXe3OyJsuDYdvbA4ySKBV+Iy42dYJ
tTiuhCv8uUeno0JqsIgQ2mRG0taLu2NiUcn5SIrg4yB8lDeO28LOHC0aK1XFmdp4
lr1glwOemKtXVw5fB1mwgDnbbHk3p4drDoEMV5F3loScQ4fHU3tTYrJ2TgsF1QnB
B+IcsnzIUZaXgocd7ROsHa8W9JJFta11q6y1G4yyxUXcs9Loeh9YTXNm8AEvgBUY
yTONq1bsAoLWqqE9qvM+CpC15Z3tlZ1lJ2GcKCH9cQYMaoe4d/U7o8cXv0rar0BT
W60RpIFoY/QBaopy//76SAtvxiSV1z0CRvubxN8ZUTv7vbfuZ0CM3pqcmhWEbmjv
vMAAC/fSquGTwHJuPbHwd5ar3CpiAOaic/yTa33j5RcVgz/Q97IXyq2yGVM5MvmH
DTQbaIdcpxr23zRCKSocOYmW/ypO1/YpLRIxFlsKL9H1UwAsKBYPd3iHKQtlNWL+
FaLICMCyVLuCPhnd5/X+4RKoIdkJb3j4SYbs8RpXXnVeSYGzFLGSWHL6y1/pXhFP
YCBA4dK36tpAkO33DkNVFn96UzDl9gPSsHu6I2RjC5HU6M+GBgLCtNi3J4lplXk9
5xBrvY7gq3Bt9IC3uebV2BqUBpZyuocRKldO2DJOY+gKNtrVd2tDfegnYFfGPnpz
qrQ5S2kKkB2M9sDu+g6UuqS2d1VPrnbhg2vI/jrVrV3oEJlMTE5Vojkj1PGnbfO9
88SO54/Z3IYfGLUKKE8RQ/5rKXMljI2vn/j2fUdRQ8mvtjxg5uVWUcwV8aMQfHvP
Fhy1A2tqfSFKa+ZkjzRJhYRzsIf5wed0JRtsCC5sA2EKf19aA26+f/bWWroO5HEL
G5vGWk0cYA0q7MDz+BXXGS2xyRXx7CcgxF+kpb5vKY6JeiIXaAN3DnsDkh9km9tN
BmIIM8DYwg89G6O0FoZrCNhGZ+X9c/GnY8hTuzrA6wEFlzhlBB0ILnAkqbWsuWik
o6tzW8Tl+E+jjyDYKoTCwu0fvAdKDxPlE0Gl1rLJvx1/yDqrnoTIbRXAKgaJlpWQ
aPJjrlfcnreVyw/A069cAu17dX38/68QiGnlCoTmUjZXJ+l3IqoWRN8YQgYH4LVP
/F8C0qwWVg9sZyqPwahLj4t1xncnmhMGMjRqfoiMF/ZO6lCo+QWfOQJzFbTur9d3
54As1pHFhqgkQ0blQqGzcNxtg0kRfD7y4TAbikTmwnEI4MPzN/jf2Y8+VJUlwOLk
0nemvaiVKEZCTp7HYj3hmrga0Ia0Z6UvVyLW4rLfeMxaTF61lN9oURYUT/bEVU0y
f8VlUtZE93qlHUwznBpgc3Vz3/m7bzA68Ibv3hqzb34FxAwwBGTq4GJXseBVj7Nd
cLsoJ3Ex3uFibA4edY/9aZYg+lXoaPVRmI2oiUQ7fPiivwW9hxmS3PbJXyBhH7uH
VAy/mfWRIjzqb82WL3ChU2TLFLyuP54yCAu3gZv0NgU45OYqf9ODGEQDZKkZIfkS
KSHtAsv9ymD5+MkxjwrzZrkucQ1jGDwyhlxfDMhbZ0dnY3QNKjPP+022Kmsi0m+P
sv6tIHoxrIfww2tYjxVU7oOTtCTaa8D4udh6g+LtBYIeZMw2i/qrPXHCi9CKYani
/03kum9VB8KWtRGX7nhlikylpgr6HJtPS2gAIk7WY/cin7vcytS9NIRqIqYhfWOK
HzVkMo9SbXm6fEe/5VtsexJ0eeE61HM3zhPjmoPkb26Lc246vQbe4HIacO/IlWc1
e0BVxa+d9VI6O3uHan/tIqL8rtsbmVlvU7NIekHTQAv9bCw1jB+8puj8c/XsPlgW
hlyGLhuqKhs1WiOHbwcyNdNxr6LGzfz7/D2UqeV9pvEv7ao4YvCibqKqOYZdlF8u
B/M9W79aoizEjSdXRNT+VGeT3zs3A1P6IV+S9+Z29KKLEMKQCWN41T8xIAMaKJcC
FX7mdrkeWL1C3Dmr0JnzGrWqOb2LVCXADQIq11u23MsoS16GNIb8S7OIixd9aK0h
oIGuVjsK9/iMXce3hzYtj7AxMPm7ivmdLfgvO9pxoIwRu5NtR/Iwy69GYOBmV2z/
lp0orTkkN3TWizlwTSAc12g0/UmnKW7acyN2C4GSPb+XDReR1192nASew1SPQmKf
9yO7RKSbD7fpxXdmIKVzuFVAh+BOpy3K1Ah2m9eMC98JELB2JpNZk7wkq63jQdM+
uSKZrJvFr3epZipRgkbyqnpiBpwa2vG59/tIpd5+1/YpJHZjeLqme7E2Oh8MpAGG
TSR7UPC8oP1Pp3w17jFu5Eaz2TM8ygYB61iUPs6Ywmsdqx16DsMBLPEfu+aCYm24
OmhEc2rEm5aWm/LNa6eg9waKkwW+o4Hf1De4rKSuh5qceBCR1jNfc43K6OuWeIxb
lWmJJ7O6fywVC7xLRSwOfgxyOrGZuZoOeJabYbHoMbVc7TaAYLrWjfHPSZi/AY8A
rvsym335n/KuBCwSyfr2bgxB7sgMi3akeDC1ckO2v1X6dsRM+4KHwUquq0vRyIaP
NScHYtaVPwgnTJLDZ2beEN7sOqnntqbBS/EudON7wSilyhqenmolS+rJZZ8SyyuY
ofaY2bl+XryEB0a404SeRJYWAJwiaL/99ARytezxOklohDB1NkyimWQL5Ol2Byvc
6cTiwtyIbKmk4OofMAKJS3OuRId4c7RQlAS9fQ/guxSY4MmPmphzHIw6XTpPD4CJ
ZQV7qEW278obZyDO9+wt777KIV5zQZ/RNQ1mu8Lzxwy4r0WJLGzltK5Vo6KNyuPv
lNf8JWd9julVSwFCljozo7Ymn/vPWicQQ0Y6bRDaMGKhjInMTstTA7V6tUuzFuOD
y9G6isYMcsbdQ/umUL0gJUxE2U3rm/d5c0FofMUaHyTA6zGr+ScJXXIVSLNzvyJF
RTpc3dlZiM+ZU0iaidKTYepVaq7dO+BlKD1F28LSvUZLUNssWcv/4Gqig46iueUM
oqtnN1SUMXPe4svkV9EFNEb9axltjrfalGyeShKr+6UN7zDiznSYyj504GCprmKY
sHv3ofJC5qJ0z32BBW2ErGmA52Efo1lAWObq/Ml+xmY6oIOoFmhbD3/BDA7VWuCY
Ra6MFxwfGaxtBPjYBVdbUmfr9F3VErl7GufHTPY9sCIcdYTQlPnMx8fwXVn3/At5
mSeJjZxmZpCltzNQxvvvFXMdPhI8hIRrBfMIMEtweJO2Oicv05nvR1S11K++SvtH
Bbz4v5nJDusH0XNq0hSbHUpP0/NY0RbRMxrv3M44QWZESHDoSiY5wuKPjNl5QlLS
v1p3VlCVghQvCs6/y0/Qvy+UV5soC/piCKCfvkR+i6Nul+mBnXZtz5XFr+VXag2S
YVcJylFjSLpWB7YETmfZ0MXvS7t1Mrzb4EQTLjIb7XSjWnAABQduUSrdqN1USU2L
cxQAdezmon4NpjHg/DFdDsyZBQ8PIks0/puDsdgzoMJYfkopXhAchhWsD/k1VC8f
GD2tB3LpuLDiVAWY1grOlPkhnyZeU3sjqBAeSpI+CNsxzbLjxPpBTEAG5kN7ys42
AP69wVRo6bnZE1x0bzKrE8I0KcscCcDGvP9kiKOe1NKSMtC774cAB2O0Kvl722TO
kp3ew2QosDuXiw+8ij5ycAjhiYOJuwJLARdae7F+HolVuLJHtGO/wZLgju0Xfnay
QGOQkD/sMzr5jE2rrpJk3unbNVU9JnKGj3QkqqtIOjhh95SWBjDbg3Qzm1wmRRgx
czVwcq/ACTwnFKTds5ngGA8/f7TKjOpnsybQ+IK62TTBQtdnXwrAXmNqa/oLwcve
fMuMzX7wl5cY0t5I6S/+wPHNL5uLRDmlNnc8wd5M+s7iws+SNxzEzEktXgeh2tL+
obsrBCGpNbXZ5SI/owY0aKLyUghTHZ5GeuB3bNQU5OftdPtFzk3fM2UFgvDsBfKS
E3qNSI58V3Vi0FFqOBooU6AKTmloRN568fsHu06rhbkGdcJW0+o9ej6s85oA80OJ
PNYE+v6YBvWbIMVnQF4N3wnE3s6xZgtWjvYNwtO6u9autO2GxpiQKiUVdKRJHHpP
LFjQ0thhVcPZUqSajco/ux/L6Vc4ExsC1gEX87jyR5qpZRvw5GIkB5AjIADCl1bN
FqR78I+NCwuXd3F2kuodJyGhKyz8qlbuhSaPEDAq06tp2IDzm4+eqfAOlJNpwOyP
shalnKkqCFwD/VbHS15pvc0FPsCUUBDQSOC2Az/CHjWJ7IFlU8VqRKWxB9D2TWGL
qmoeaRzovLXxaCamOkQnLmV2VnEb2JefDfobrO6rkGUulg6jWaXHbgnmnrWcz3py
iUbLvFrEdUQxANZTT63tUue/TtKNgrJSk0LQGjDkXlmRPBa0Nu6d6aSekb8PGYa/
odjKjYdZ0X7CuDWXQuOT8xZGodcqOrJQDSgs5iii1W7U4AADNN41hjAJt7p1p65u
AUXEeYGIl+CTYxWRM/BiFqa1/I4my4FHlSKsHBLKRU0xJJ2/R1vpnhQiP+BAcuRO
5dSrXmuO5pp30hZutzTf/D1li2oCy4AKa0RYoG/T0vxqxjOu7GDM20wurSoBU7TX
e8QECGArEZKvBfZrDKzF+OypmZs2QLA0mwt3UX9TQ3ayW34r0cU4yyIxje4zUpCo
JJf4NBmUsVHjUFzB9ZOBIeUwLAaPWw1EOLphSw12OEnHPWZSMmSXhpZAzr2aAyd1
d8OcvN+u3aXJlkc3Z8ey7mZ5VxSAATlqvL0/Fi1HdOfCOagXjjrNpJXRYJesKR3n
7TI9Oc/NiVC/wAu9iY/IU6dvqUqAjAy68+OgRRxqzb0vLDLfO4MNdpVplmIomTs/
2xTxus4cYycHb3DEaCjz4e0eLoVJJOotGBmhcjbnHhLERxwzb7iIOkojLNxdNmUF
R0+1whNanA/t/SaIBCwZjqOP5ChfLngaB46y2VsiBcYfVMor3b3iL3hCZu8Kh0Fj
nJuKpINEvK+uMcy1CX56InZSBfaoZakhhVbIfSdaXldYF1hJ2pWrn5XxmzM4NdM+
kUOtYA4H4Y8Zv1d7ynoYFS7IUqMUNVA6/25T+62zcyRqe2I8JIQ4SpYeFrFbyy1J
3nPePYDyMMW9koJNi6Xw3/sGxgmdZKw6OKMXqO9OiDfFrJNnU77BF+bT1oIRxYak
H1NwQWRJJi6zgQoEdEYofQnYJbLxKhg/T3+u0hjelLqqs+WOlDiBMNZMBAF0F6bg
dscExQRYYWre/vAr4d7ntUOzHqHqzhDsQcHnWNUEYT6TtDUBeZDCe3qSVqvXq7cs
kE3bzu1j5EEVu+dG3j7m7omB7berofgDII5T4N1O71Rp/AGsA7S2S5ZqMG4zwaVl
nXx1zM8gj+y4KC3xtS+kfONVLamA3H0OIdMWTYKYLakyFHMwLqUs7JtHmtXJuG/a
nnEOtW8N+777TB7gBr4399J5l9VGdLHCwuxuNw6TFnnht4lXM2AjZBKDRD2gQIt7
prkR/YuFXgd+FQ9oBSHUs2QSTyGn4jkGfBVziUpOQd4So8WfZHNCZEwKX8MQEBel
weaUG7T6uj1VBEFjYbribVdUGIGeM18coQXUWd2w+48RKqrhkRPD8mA3gkslT5nR
XirzxDr29YYcNOqnrCNJZ2KVCDDY6M/I56GRFkOnkABsD1BU+8+rBb12KBfUTGow
rn8r0GO3qiF4mwmFpMgVB+AnA+DWtl+XZ1lPMO3C8I63b1K5AQM/9SCXBBE3RsoR
jhPVfbdvQCUvrfqGpfeOj4Ej1ZThhgSiQpgeWCy1sIANKPxsziMuyDA4rVv8kB5K
c64Z/6wqSn7FpCEi9Z1rLq+QmHmRlOAmudkLa8HUeoF2LTyxpicR7+9LW/aiFzCm
i8U+DC2MsU+v1xu4qTSvsB91ITV/ObsWFUUvXpZnwKlWVimCztBC8L7uzC657GDi
vAyogxWTFhsCedhX8qntfc4+F7/NNt42fwOkH4a2LZWpf5FTykZVlEQsDXI5hW1a
2Tl4Yhv0gKdrOmGLQsuFKpDF4qhBRfQdd59pMNF4jcauX0uNCyCX7IpC/Ji4f2XF
7ghlv1uQukK1eVZ6e2iEwYgGsWVeW1rfvK/m9Y/lsrmDxyrRlZPO4veXovpXGfBn
TJI4ajJDB7Z9ZUyuiZpHHdg77aKSSWeOQ2jADxmq85tEtePuwe9MFY/muHTmqqtL
T9XOshJ5FdENzJLRU3IWpSY4qmU5B2rQO8/O8NerLvWfdRib5OljnP5vi+clk95m
q+ZWbHkPU3IC9wDq64fMYkDfo4dbMTrZqTbtpIGDfETQ/MQObDUiSOPTNqZjkDiW
WJEiNN/cI4hcp1Op3fXWF9m9utmwHfJp39EkdW3i8JszfnqKP1ulnxbSnpGfmzFn
SVrnc/+JhiSDjVYRqCIjtFFThRw+iaqM3yhWL5vWyv/QTUiX9equ6GbP6DT1cijG
d4SLBp0OuhWg7RpReJ2hlafIjRs+97I87qOQgL8Dkh46e30yzan+lXg9GdMHiGA9
QEMG+rTlKd0FotFeqpi11oy3UpwwXkvx0KZ5/W5hsZG8e7a9IgsCuhGD894fuVco
cBSRP02sLtMOER8AYuVQoXJ8xzs+s8z5YOX8Y57DIsu4rd8U1yRwmiVbSiaTPlGH
C5FdnnXzlceJASb9CqTKymoinUf5qIQ3DZ4vMJhQAKrnlYRtQGBj+OVQdahKZnNv
JNPc2+/1wFs1YrWS/VDoDfQPX0Ie8xHUzSo5o1PFzOZ2HIU/wWk+Urzb4Q3o4l7/
sBXKDRwD3XZAYXJmEcN+aVYWSiKp5/iCjno/ZVD7jL6TzHyUBGLMieqIItJiBCzW
Spk+NErUePBQz4JDaRWuUZXZSqaeEjWmed6T5cVI5TcIkXswRmtmktb611e8w1I9
nTf5uuzx+E9MxwdeQYT0PHq92lD1+XAmstcpKnLmEIRy7lTVkmSzFvHv98FuGM5O
dAVKceeLO6cCQkplO2mAF3dkUm2VMeZVEBHj6Jhj3vxJkgcNJ40coImZJoeWSpQ6
k83iAAyWVa5O3cEzujUyMvsFNIocbrx+7TM0dHacsR6IginmWJ2f5eWmjtwdNCQt
eSmFtkXw8+NGyO2Uy62OgXWODBrlctFSG/1dkzgsutvg5tldHV6UQj8hR227Ffvw
aSkJPqkou6wL1SuSfm8ii+TQU78Liu/wmxT3dwo4+lGMAkIH5hVZqqdnM1KHXkmq
PfkFBWzVff+EvlXsfiQPB6779KySrfD2nmuAMVCDE8VHUAg9A+sQKvP35LI7X91j
pnu2DfAg4J3BwYaBYA+7Kq3TNIkth5iZSTLYRePZgSFYrbGwQF4JqI02bxYoa7Nq
3TsuQ42IcksGzgAadFvj4tdGzPgxKG0PE1ghaT33vpY0H78Ld7C21d5xWQ3J3kdr
R1E5+B06p0P2TGmNmhu85fO/QdTY9uDV4ifRRI1nFTqsCKJAjabxu6KJEGu9Gts5
HgP16227Fzf30JG1brMQGTLmrPijUbNe68otQJi8//tyea8ffGPwb7wIZICinzDL
n++XLNBv5y9YoquvDiGxuEChHyy5KRf0vL+72xlfSsBmzzNgOOyQeGuzKY0XOsVi
sMsfACGhY6Fsp27Mrl9xNwywH/ymWf8QxpO48uSDbw0tYcvKmacHqu6F5vTF90C1
IpbIIC6FpweMFPU5t4Gd1WApj3541Jb+NEK+5moX277Pvq95wGgo/ZG8WR6jnp/g
yzGtQURA6/MUceoDOb/557gS4cmGRvq4vs28kduAG7lssIf4OUrAG68Z9yZDl4Cj
Tv3mjgkLTmAT8kmo3mscf+epxpxcyLCozbeCu20eKWebGoJsSyKlMnflMo/SEQeD
UM4GfIDJ0LvhWhY+i+AuKG4WXkV3RQ7v97kWmJoWNyDFu9gdyK8uLLb3/ZtOaMPT
lZLhprb2JFu9eKSSaLqsnj5jRTBcbG9vJf/8xFCZ39N1DMNC/d3JeS2cOKxh/a4b
ag/2Bgl3QshGjDUZpaDBcMBKNgkccmWQLsjstpltWBo6AN98rJaxs7cShqODa0qy
7BMh3TKmv0fW/RVM9r04EhMRu3zm5VGGxUk4niApYdIb4qyID5LwylTX14x/akY+
g9pYKX464yR5O1icGCt6Z0reEkYTvRJoM2ito1Wfe99fghlJ5D9v4fj7X/yHjYT4
QaLiTdlwq8QC3zzkjMwDN21KX70M4gS6mHWTbkeQnyJAdFmdeAqzsLR+uaXwAcJ0
BlKgZm2l/t2zIFu10brpv+y6K3DwSb47hpAbz4eFA969C+AetB06rcbOVNJUp9OP
ykYACTxCzXbjFSP7jInvr0O8tK7x+t3klDCkhO1bojqVE+67Mh2F2vVcw7GqRT4D
bIuZK/WOBhU2AtrrrHTL3EMyNGm607WUSW1M3sgA0ONqNMob9DBmnusliGniHGyz
5W5JuGG2X/olleCUh0pt1Ta1h5aPYStD4QsuDjFhpHoq6UFncraHwohO+KbkI54r
Rl29JoL0/1B46LXOHHxspHmXTeBFIc+73BBgdQFbNmCYleZJMDj2AVy802GQv2gZ
PGRrQVE1Wy4vlsdRR1wPEu4cWf7fOydgSiokFL0Y657lR/IO9mQqa478qbaGJQ7N
FmdqFLoQlRbaWZguNQIFQCzCLPhA4JY/WyJ/vX1p9HkZCFId5x/Lyzq74f8V3J71
d2LDlIqtGZZtoYpSX6jyQPxeuYzix45nUJo/Qv5ckJ1Gd7l7lKgaqg4pGObxMjSz
ioZEt2ILhLVtjSc9O04vE61Sw2fxcvDsl7bPE11gc5gY4Din9Q2IOejTl5JBAoeJ
bvlx1TIxK+MtFucx7j8rXXq0/EpmGznPi8USYskHwtYSgf46xujJ6opaBMoCC2YL
BINVizt2e/2HxOao3S0hMRD/1Kl7ArGZMPBRXN54iMXVEEQ0MhOh4qClLJMSxNwY
fkH54y8fsN7SaxbCnmpTrUgnqYtWmnhHBnEdKm++LKTSn4etMVRLFk4+rrBGX3Vp
SBCLwmbKykgTmgLWDPGAdr9HKk9I0wHqieGXHjLLJsRWLWml9zIuTG9KG4gbo5Xj
1WvxlHmBiWiTS6X4wNxhSK6j8raBJloXo0w6r70SIFLjvqlWzjrXG/BtyLMNKbZa
eSzfjbcJanHb6LuvrioSWXYf+AzEkyNgeBjOVIbc7vJJWp5tYm4NOG/nYMFBYJnj
M9ai3vlsDFpNRgM8zJc6VgmD9+7QQo3FzS1h8c+PmJsZRHqXjhcv114nmnsoqRN2
Mijf/eN1I/xGIOUEdZ8dHCblFdPROA6ZBxP0bLmud4rOsOokjMV2P7W7UfFh09Tz
lcNVAfuvgZWDYB8xIUJRPqGTh8CWcc4ZPtLW3SELHutMm3b3w56oCpwGRxMrurv6
W+iwm5paifZEJp1GjIILHV2nK7cotUpm/NRwmsnWjVWhOB8C4n5hy3zBKnu3+ECp
nMVnEJcsuo4S8hmN99WF03ifN70QTf2wGT7ZTwJgzpko/fn08k5bDdTJGsC9Yx40
Eq7tdwaia6f7GKLyLeB74P4cGcC7PWEX+6leUMYvL0CtnWKLQZEw8eweAJrW/hwz
cLWPfyZLYHeEBJ8y42CnFCFODISVuiXR3U1aP5ap71vWs47vxmHlLZQ51xBcbQOj
S6MLkZ309CSpEuA+hNlXRZIxzNaOQEHjPGg1Yw02W5iHoyyaxoNZN2+LYBwISozi
zqNiWeKKnzzhozedEUhVQMk/DVyJo7lpE2KBjXiP9Vf1nQblTWfb0YiCRBFA4kyi
GlLyyj+3vhghWYkeCkV6tj91GDbCMD8UT/utJovgelJsYIZwST8K04RjT832pYbJ
5bDMR4PD941z488JnVxxjWINlNqMbDIeMiKCouP8uGgN5cGprDeBxzVcJK2e+IMx
We5v+WvPQAzufC1XvQm8qJG7kbcbTNA6GN8/TGmwVRRiH7cQFey5+qum8SuUnD42
AM43GW86MbcNAYRwplmBYlGbNrchITn4fGtshryR1GKgtKJ4JjmoKA9Hxuz0zMcY
DSB6BRZ4BinFWE0qSg896Uk4gLYZMMAEgMj/o2J2bVeckV3tXFStTSaJ37pxXGdx
p512anMDhHhxRx/YIoc5DCD+edkgutFl1H46gstZ6RXtwSXR9M/iMtH/3UdkpyK+
ZwbMGUVVvhdDwbEgfqN3Yzxg9YrOGYjYD3HsooLjJM2Y7rQ+IPQEG6k++vC9QCzH
xXtd7Oosq5znSXDsFzaarj2oj/KodhQEso8iIci2GGReD8o5qxUmmLJogLYun8vV
DJvQBhOa7gD1OW2hgXvJ8mxTcPNJvQ0o2hAXBzScBdzexlKAMbJbs62AqWM8Wcs0
TLWLXyGUROnS6zz43C9oM08N8gTxoR1foT8lg2gp7HReMjgitvrvpw3v1q/ZA8DT
zlgHQPbKeoSR1DNMlysgE1+uIk0zPm4nNBFO8IYZIKpSEInA9ra8XdeeBUKEkYjn
ame/HgizQ1Xozo9TDlLeAY/nzGTXlyIkpCSp05eWu+KC4Z8/C+jW+K67j8u2jf/V
oroQQ4w/B6z/y+MKjlZmfV0nn2IZxcnbV6B0EKAV7kaVWiH/Nk7blof8E63qoDBS
MID+5AFjledrq9qYDRKMNuQNheLiHK78YkJcDUTueDSV32W+0ki3uG/Ohqawvovc
928JxAOxu0ykJeQIq1IrLSc4WI+rTVKEPrtlRuonKrmCLbh1HJWUJ4cWFFr0vTWH
SwjgGlS7Whsesl5F5cDvBwljftZQaz7bd6Aj4hLYSOi/lMu2vCmn/7tofCfyUESs
wtlvyvI8fZAxOACQUmQ4Cpr/7Lz+BJvzOFiUin5a1QdjHb2rrUWR5Uo+k2TTdWuu
3FT+T5aEFERvGXre9xQ7+kkDzQCBLsVY5BFTJn2BJVqlcbHo73j2b1a+sHKUB2xj
jAzu/unFYfn94K92lhIHZay7Z3Q5MvrHBV1eEd4lAL+AvTyRK+ChhFWViabtAk9/
ZknNwEYw54pmD5GuEZjn29zxSysNozwj230ivsYp0fR/jBPGw1kAkJIRHrjTRBSH
oW+5GGe85DfTxTrPirlsmk6dn0Dea/Ayy2iCV6GdPYt/MnORK3uzyyJf83QEKYNd
FEWE/NnoVMBR6kTskm9FARlD/WfGwOyvZI5SqgWbnGBz5ZzJ7rtZUq+e/+KMAPdC
MX8KVKhaDAW/lVNbsD7ikK7KWVJLWBkVQ6jCegEnjpkJkBMPTWuaCDJBsJCzGTrN
OsUFPLMVynZ6l4q4KHvUfO3oH2zjWnmD50wdmR6kvsdTsBLArE98s4quvRmK60Js
HeluCJZCFO+zkMUA4W6GXLEt4UkwiAWEYaSND/SLsVa64K6iBUVoDvHFCLqOXXai
L3kUrJrzbEweHcgPFmdGjf9Cu8g5XFBrlPan+naj5mkqNpg2Je/iLou/p15w6DS4
NGmN1NZG6BihyiOvDyHwS4+uWAdl5jvG+6jT10IHeM4mGmdWZy/+Nly8OBV/zlGp
xgReTbU/kkh8vahd5tmMRaqHEglfsnyZ3RLJuWz7TDu2N0CVirbRNkl+WZudVxYw
iwA5hy0NVnSeTlSICE0PWIDgOzfNnMi7+gEJJXVQqmt1eqJpzMvTVsWcY3d+RSOM
ec0thigLhpMnwdDOvSnjoj+bwR8GReu4dvD/e6JBtciTbyUnFI5iWbNZkAcs+woK
eAhOoNjZ43nUkLutnzSeUZfMjQISCug7OULwZfc+CtVXxSLROI5pvCLiOgk+foYu
XYzFa7yTbRRHe3jucWMBArtwjab65cMaPRDHCIEKHjdgRjQ3OzwxOKbOiV3sc2fm
zsiaDyo4j2tq6Vj7YSSMX/534DkyenpeR9HxhkiJ8+cSCaRfyZVxtkHKFElfw9cb
oj8V8JXzr4L0WuXD+Va8EnIVOs/PFjpbVuYF8qMFE1EbyUPym1BXdLwHe65i/zR1
k+TneTHENB6nTU3KpfyuVNJzB9I8fJprzqnWZJHo37xGD8i6vX21K+I4HNtlAmaf
KHGPr7RgFptDJEIk5xV/1kqYsv+Dj25bIjBPXYWXSy39xm5b/ilby74Cltvx1bGx
I6mXxlLyfwU6ngZASGs9IAW2Tgd7LHxL8hv5mDh8FLIMUTst5/4E/CZKFM2tAPWO
iADUMvMtYpt/1pE65nZdDwJsBupNIvV1Q+Uag47zDpjlyYTsaajuhhWYz1bxmirG
IxrpqNjVaQkMTNIjb/IPfW6vx96Qpgb2XOnbmnZd7giP/LYaR0WVhU8rM37gRqKm
j1vMOnwmTIBspv+td3WH4ouO6aNDpUjFv1AVdAWIvOgqrAtzQ+rqHkFoJ5+W0L98
EnCUy9eV+Fg2jJO/oB+8Wwwjw3H7EWPdw33hDDymKgqPQD8Wi4vdfJVzEqqOk+rg
2efUBHodWSZQDZnlTZiuow/wIIt5ZvxUcwj9WrwGIqi146EcE9X8Nmt4C0qy9+Rr
H333/oHH1QvT7NR/gQnef9VRSr3TMGpjekmePOHLqna6jDOq/QV/pn79uBu2IauW
WL3O8NRkC6DoXZvAJ7SmxTxPOXcGkg5A4xmtD6H49dkp2Wr1dfedmzwTPi8wqDiE
r3eqhk/G4QngJs55wdKRVyoZYgIDtXnBi2xraW5quBS1DcwT/bFbRKM3Q8o9QId7
MhNC94aC1pkKZpM55ZE2GQWzK4leTtpqsXNhUBn5lRN/ALFbIKNmEVtO2hkT+bZf
vDJUJNm1tGJtheNvIE3d8GTR1INk+NYYTQwn10p6DEB3aE+iblRkNDXBq4soVDH5
9VemgyQy3uxBGGxxuMVSYJ/faLJ1JcWUy0s9F1AWWG2z9XU3N46zm5WNv2gT7CnE
TWiGW33HujtAIrlLlfLTHLNi/6jS4aOJdVVJarpXN1ZL8671Hs4GkyLWaDgqVW8x
JUQxRnNvozK/rpDaVpo3XpVpKXNzlu2WtkmN3VCTNfRpPMeX48zK4SsyfxGJlz6I
junWYvKSfqogTVg4kq8O24NGwgbx8XvYUpuWwwKS7TGTjtgL6vSIPhD0jfoEiFqN
VS76aVEhWa8a/r1cFI7oTl2JVR7IMxSU2W8WuSOaqokvHywHrM230Oo54bMjS3yV
jJCCrd5otj8w9AVf+eCWvLCMYRluBgqLWIbUU7DWWmzvSVNPPNs95nkHzr175OZu
1MLoapRjPLFhACIv3VBANPu31+XYN8z+HpW5X3dWIwsi5JSEbo3d31kKdyxwFTHn
gKruBR2jaodZFVpMo6tJjyGDEO/e4wJxJom+bsSj9I3awVaceb6LXbPR9hezh6Lf
UNmxX+h8mdXg9PQs7upeHNS4+PZ+q0NqKye4TNnfva65H9ucan1O0TVYr0+swNK2
EVLQfeQpzSvB4j2Nc+lAtmZy7soMfnW1Vd0OM5lAV0FhWxUEqFZRb3dY6Rpx9gGl
SOWsr2zAKBKwKsdx4gZqGPbI8ZtddY6H9EMdsalO6mqT+nlMw/wudRhthyR8tfy+
fpkdw20NQZSkFcYDA54Ito7mvTyChhU5Igyrvh7vBMP1Uk9Sz/76xUsRWxa7KWk+
Vwb1BmJXRbhCcKdw+a2/q0sbK1NzetNq15X9ynzhdrsQAOVqf3esYMK7Admh469T
35gj3Wv3sN/1H7ZixdHfXx9Ld1GV/UNdJE8D3sWLo9F8WdBO0AmpjlhSFRXa9Oxj
sOpKmzOaYB5x0BcmEuYpz311quCF31mnDTPX/BOFFlobD7cnHziMrY9aiSBu7iIM
3VLxR4wQ7UE8KUCdCJslxaZMfPkWypMNPuvRC/9EGwCJLh7BoOeuu9lW6TzBCdau
sD8whPOdrcjoAYdL7PBtp+VgLm7bvqb6HgKRHBINvnNF7VVSZTmMoLzLn6dCAWxK
I7XTXVdYAb1Pn2j2ci7mijHfvty/+F/cm7tlmwRUpcxctRZ4s3BA4C8v5sbkmyFH
cRXSbsP9LkljPiXM8LVjTGvNVHM0evn6tL1K8r+L80oUkldsyBav7JhiGE9X83cK
fASyVgPx/XmNgscS3M/wS+SErqzlqWrj0s8yFtQ1PPISjCP8DqG27y5ZKBDAaRIr
c68+7vyny3rycPd5S0e/15jJPvlqq6mGJaf8pVf0z62Qy9uUgJmxTm3+BqItoOJy
kb8E+aJNKnkXH/3lg+qOr025c65xvvVN2lbFKWvjO+sMA+eO7zNahSHf+IkDXRQV
bVi1Y4UjLaev6gKTUNxhA8HfhpxWlmLuQCM/+WvSYYGs6ke2pLjovWv2nQ/Dcxl0
qYEpJV9QxhskDwYRw8VhjgAPh4RliudijsOP647XMoCcOMa9SXo4KYBSN+Oz2aOa
SBAImXMzr7iVyPJBT//QBnetskLpL/PgYH46ztux+NoGmZqScjR7pOFNVHlkD43Q
tv8mNAPePmOi0M0htPaCve3CU6bcQJwyn759YTgmQNrHaeh6QnGXUPCbTObdu8Ct
E8eL+eIUK8RiP2kXwSrQhuRb59eV87Awwh1856C4DqQd0g4qV2fgGgc1QS5zlH9z
cpuomt00MIqUlry2trReNcUi8VFduz4ZWHP1SvPXYOvKJ8TmzGbj0KKDUhAzKoie
oOb+/KvtWUX2477H4UWqUonuOQAK5kJoLX78zOBr+sY52Wkzj0XLr571XF+WP68f
DV8byD+YssFcCIfFHI4Z816KzgwbDChHal+qB1X+KjKA7t0o7NMixfOU35+Y/9is
5BDRjligsUrV2cl+JcvQom0H3vCBsGcArCexlDAzm8jgfnNHdrDVfr4G5IJOXhmD
i5f3q5N0PmuPzeY0pjj1jX3+G2A6jFnJsiHn9ylJYH5xQuBaEGSlAiPie00KXmHQ
g9Pi5im2JvKOjhhdkyTdDzjyFt09HJh4H0doLYB/iVAnSG3Fkp/f0jdUnNGDiXTF
XGYuaNSA9CrP/jVg+Ah4qFe9qNi+glNf+F1oZSXdwdX6ywrmxLErkpTdmswrwb20
AOQkrQa5U5LJ+FUe4MZ0WlABYDNrg9QINJErUbKUcBc79OQ8UkYaBhGTFZMTj9RV
T0zKPFFBCzH8ZeFNvKCemX63nhw/XKo9oe8SM/gN54bsTkctsAmpzAyZkOyrjZ8u
zJawmBH/+Dos1DL4m50huyC66c/jk0+/Dg48shSjWjGyjtDqcIEJ5y7nypdT3TWC
/Oc4+zbF7/0dTas4CGfq/V4t/a21MYIumOADWWpOb6xjLTjVSkHjTHfU9DLovlaX
FT64UcJaOvkd+wr8u8vRkD3PdblGTI8AvAstkFVBIm+IjQ8ZbEU0DPjItm3lMvJ/
PK2JzObjpnTl+x4+rPn6TMxLjE4cpvUGtfyEw3Eq0eA/bWKdO4YchA/A/MGXANGe
fb9urBzSp4tYZe4cYOnLRUksK2fRDmJ6Uh3K71XxVTT+0v1JzXhx5PF3lML8uLAg
tXKYYFJe56ydjXsXMcaGmNaWdllFT9fJOBtrIy/zbRsd9a1Kh/ZKSZP/iWCx9pRV
wUQOY803S+6AzEQoEZnHJnmLZbN9XKVPM+MtnMMibyl/i+6vFC7pEmXjnWpZEU6i
slP+kOvQfZ/mJRMrr6WmakhIsmx5H7bud3j+Q+e8DeK31Q/m6Hlcj19MK9wemjNR
CqDA2ngO5wTgaYXIx0Ihyp8+7jz2kMw7wHPn941fNJmsu6XJxc8HoCkjIinRDqss
26TX5a6Q6lE5rJ8vLolY6FZ63tsprHhWMc96vzeDoRd5wvIb1X1DoVkxkBEx75g6
wUjY7sW5GXGTuoM8DSGUssbK9bsH/HI+pGmn4AXUnz/UtJbtVQJI6KVNakKC0nqe
AD4mfVzizKxtyayntnxtY1CIva8vNCVgAqPnR+Z5rTQW6/rQXABZzcqaXUm8juul
MJqoCO1NOXWiW4ojpsLg4JeBXm892ZuM5ynVD1r23poSxi9TLHt1My/J4RHjLLh+
bMrmmTIusl33hsNNNn6q81OgvqO7nwx6BNHP/3daNRc5f1/sX5id2TNIzxPV4Cp4
biJfy6WI44nlv1dlxSl8+DIeyRGgaupS39GbxmjzU776M0lkLx/9uJgRJWxsgGsc
3JXqIqxMpx+2JcDQucJsEonFGAErUad7TW0QuEOtP+9gXmmZ55f+x5KzQloeuOcJ
3cm156R9DTbswOZsNf8fo4Zv+hA59cStXnTmw3NzFpmbivHfujFNjcUJoUScIsJH
d9oAcXPrEPqX2GIRNTmnFBak1QEW26mzqwLTB2vqytEdyQWv+YVL//7zKdvOhwqR
PA3W+ECLb4B6WBd+QeS0+WHWwrxNGQlKvLq05PPzAcVrE3mMwfZq7Oa8e972puYf
KKjE11JuMt1O2tUCLeJKv9z+dXK+cRmaKWEcpmcyWxPdkhvzz6SsIUboyBjswKNQ
5tnxFc+K4zwLhDNwCM5pVpiiSM/nF/XuKEcauHky/Jria0YIpCRJzYet3jL/Jbnk
cDQ2WFduCqwGsFjdxruQq5qtLWwLo4vMAkEht6XS5OYSVZRJbzQuw0919O0HuJrM
c6/wiWNgsSV26lfHgyhRJXEy32wrZCiUdbCfJYn5ODr0OCewXI2CtHMZ8xCSipgQ
lVku/2Q8jNcm32DResOdPxoDbwC2CfQuQDrjR2WWp1wAi+9u834/d2IJIpYLUcZq
IvwHYIF6Wmilr9gE5665lLk10x4d98Am5ItwtArHZ10rVTAXZGckOT0Vv4JXUaK9
aYj/IIByhgx8gJ/0tBzG8JxKspFQMSXsWuW38Lo/cnSW9pgYRuqParSqMe/gc6/6
wcODNnz6XMCSrufOY81biVaPPFTpBBKwWRRQpsnlwQgJi3U9Je1f1HaNaiPCvMwk
RfOIXGISDQjvpBq8M/55jRZVQr5WHN9pvG+HVK3xuaWplCeTSkbs9X6P2G0Elq4M
BsJGsdsVdvW8wTEnASCQCCBe4rkircwqtAitR+0p5O7Amk4iv55gU4UbqjUkZm0Q
IyVr2nYZmfRJwB6G0hCy3NoCryYb9lnUirbfllyZ2CBLUu1bs0Op0tVoOrQpmVQb
MXVHB0P5vFLcQtkfx9PSj3I+F/pv/e3VP2ZO9jjI9eUuS0Iy3y+bFT9QEojW4o1A
iCp1LMYhJfOXMvcoN7jBcWzJQ0pnymIDW2UykMFdPnmF777RPT6RvjBqDUFNqTxI
v3zl+UqqPKDjMCEKD2iyn7OpgOobrPYM8EdiM3cvFCxVhnZ0UxDv5ZL4HHzi/SAE
Nd+gcFiLSF+7L8+HFtX3DRnCPc1C27sz0m3KIaiBDNqK6viidXl5sGjke8ZuVNj+
UbAHHm7Dc6out1crw/0Rznt3umB2EQBi4l7jFy3VbiN5ZcwBbR3IlPe3QScvT6mO
/GVXupD1Qj79VL4LKHBIdkG+0LIpglCyJ9luJc0dN6CrRbYmp2pSWbFzrKQAt0sl
ijJMQp5IBQvem48nFKnQmctoJ/0WtoeF4kwEGG1b1S8Lr9FeuB7ODhms39e3JIe/
Dwjw75ajNxHt0cdwm/tyAcd5vtI8Sa3CHz/+Soq0UdYTeONcTzLyQqSZE6ls4Ung
aWifpt6tunyQpK5uIGgSnOUWbkU4xZsxain2DEPXUy5lLGr9Tc7iJibdEmjng7mz
IbXpzZxMc2W41JFUEAvPsl37Y4JfDWkHjWuay/3Rm9IZxpXriSYLzBysJ91HDgy4
VIGeHlNp/R9qavqyUmFhdHcUUmGO9gFOezJX5G4tJIdT9qt2dokWzOrPAfW7035E
piEES6veW3Zp2pt5z5yOGTfnMx+6f9CZ6fTSHEggFtvuMYbqFcC1+gWu7g4KyNXX
To2lOYjsYh2+m67P7+P9K2ooryHU6N+aJqdEHdjfXJy8hOtm48UdXRzBswqHg1FF
TOJ9UQQ83nyo/d6UPz5SyHYj5xzqS/tHMQPPJ5EaDgUP30K042skXBTt1WRlWuRO
RvPENhhVccIkFhoz6ijcQmR8gf67A66MiwJNQIjiuqjwfMXoersSB//eTVeNKmCS
tcMCnyMgw1CSzWBq5PM6sFkDB501OK3Zvt8VKTZpM82B0WLl8DlFi5a4ALm7Woy2
6fxzpnJ9Yf4VoTdOlup/IY4wXXTFfovBPR2oyQcpWlrduuOHjTh0eidoTUIcfkkk
EX3Nsj1e8M7X3nFFtrngFIbpiRf8TqsL14Ds1ZoYkxTv2UrgA43uehN5ZZJGG0N9
FVY8XHl8YDnXSm6DrWJ6rk3YubLdr/u2nA4n7j/g8zldV2FfMMzbcXcAqaZcMrod
ciD7S2Yg9rOFMNU5qfzwx/sXhuFHWc6S2MIVKau75DUzGzWtRpVbNJIb4yG3HRMl
PabbrZmH69Sre2ckhNEod2DqEVnVLhV1rU4dC+YZCiaorzfQl4grbW2dWDnpg4pS
FSyC3L5k2dpdVZWTA+9xGZFx0XsCfI9zpxJUqYL7MWeo/gwQRTECndUkwlx3oqQz
AZewUkBEF0NjiWDY25oNqObCDjn0/odA0hTTKSQNrBmoi1Jafzolvnh66s76k/fY
KVFrrf5vkqFitBc4HBxwKMY37gz6qv9CHMVSprHrSfvgh6Y3q3v0V1spNAJmaDuz
Cd+CBd6tUMv5rAboTVRUQFbel3STCb+GLi8ErU9jLHzl8wYqTcNFMZGaOgofsr0g
pnsbk16s9+rUYC+LaTtVKTx6pg6mwkQKsigHpR1HzWEDGq1rP+j8kNBvaig+ORB4
0VjZy61/PDRt4AxPK5gQ63czjuVDfqnOUCUJmS499dtElgsTxlgEqf+INn8VbAzh
ZEFhSJOczpZQe5uoULLioUu7uKfp414Pkc8c+jiWKurebVFXesjqYQ03dhwguLa4
mGb6G19tfWz+2sHYQJ3bKSn3TciLPO2BNeK7eSSnYUQksqnNcf583hsO4Y7LBUkY
ojFuwGzNXuVYArZvfB5LEHwICFaYMQSC8EWP9WNGOOmh9dpSQsdc7DPlcxwzVV8I
v7SSToeoXXhcNujVDt7meTXW4b2+rKsMzUwXmoGc72JSkxnAM5Ka4hEfnkSY6qOK
rFqBSX8n/GPPVkN+dETdzNLyo8+Q9v5ofYhm8JVQpEITGyeNK/FuXkDbjWPpi3O3
RgTXRA3N4PcjM7seV/4b5izgWxnJ9FMD8MM4njvIOOYaWEPGATovIPuBxNM+2vWp
1s73wOYGbZ5eFWBi8wLnF/yZKH8FHpFH4hsD+4en5trz8fJh9Z2H85ttzFg8B2zV
p2dyjGfNB3dr/FgAQ0s18/HMeI7aH4plHzwnA1/FUCB9RyPHKNFt/x/fUFAyyy7r
a0U2Zzao18F1+JImh9Pxnl8A+Cbji5f0kq4sUPloFq7N0Jd1b6oze4LBzsdV/9Mt
kpt6+I+SVs+i2oL0aVONzaaaH9K7RSQnn3vLsquEnYcma7FiY7wHEJ35xywLn/lC
ZqbVQ/KyuXDgEwicBC593nsscbQkv65lQfAKqF0nOen9FNlbvCt/reoh2PYne5jg
l7laYE/yOnWqLybDNOkW5Cv9KMLmEGWYgkqNo8fsxjnwuLJ5mSJWIOkjAgSfMlil
H5t8V+Iyb92TpIh7pRWMPE3KcKziKc0Qy44zm2yRAA1SIUsOH+oL/GhXmiy8qMZ5
9CiYxeC1282Nk6GToIQt2tJt9Nj+nWsSPfof4kYGoiZ0ePJ7BYvlWUmtBAY/PRj7
LkZGeld8JfhcExIzoIb6Tv2RifiGWgI/tc4IjmNwrUtOXFRw+zj146eFTdkwYpFM
kC5Y8Fvnb0CAzq3dD5D0D4E/KhsmRmFOIRfSXt+w7Kt7w7ZbskLDz2T747lYfm4S
cfzsVmhp3Z7C1SByLF7+rIH5nZPmD3n2By7viBvbe5OdrDzx3AoZZR1Z5Aq+UCSK
EsX+B5/xVzkqkpXYz0604/7hk6L8bu3khlhAwPkterwKmFSAqfougApKYsdlCI69
rCGTMK4MiSC2gyB+NruuQvqf653r9o6BT7MhiMOj/w+UG2fI8l7Aur7q2oqeUNsm
2dQhpELB1K83f00DWZsTEbIr+lHegURjBA8RzQMZKl3Rlf242ateFr3ACrm6Is4O
XyaK8KhtC/LLQjYQPa0BC8GogIno3tHY2svHnLx7LHeKCuklXn0HxWo9Xbbaq/TV
eqT9gBhXNW2dF4U2a7ySyZ9zfw/vc+P4Pk/OJxf/qDhjDj0x2GntlLAe6DDuyG5E
94rNFG18NteatkSICksMoJOX02TRzr5N9y0U7fkPc/v7ouxyxbRajPEjRKzwMifq
2+5FTn0JAuIffCt/TVekzIkXl7d65SyW5ImNpYQNJiNWrWM9iYYbfz4I46Qxap7P
7k1fI9B8KjU2SYDLNjQngjzozDbsSrAHUILTSHnZizgv1Tk9c52J4TbvONhs5H00
d4HXplA96/pXivsmNkAlR7a5MyWgc+Iumlc2LYLNJQbQyObtIns71uMx07pKqYm+
kUfIiRR+DxWDyY13rgjZUEHxMUmTRPOV4appsKM4SqFp95D0kgnxXPV3H1AK4x/M
HSdbh3J3bAOjpSsU6AOqqTJghXcowby222WO8Fs+RAuGsfxADfPul2yRrLUHpGpd
E3kGFEU6IXbp8hisx+Dpz/JC1e4rZ7pIKXIYz/2EYGZxIFfzK0ExLERpHwpeaFVy
RA2PW8UVovf9+sX7+e5SriBPAW7TJ8ilZZiLE3Lkr8b5rQn0hmWwu4qjkH9S3SlS
aDfQMI3zvH1aBCUTnHtzm8JwiYe42OWH7hppVENX937jYYPBj3ko8gQtqAP7KnDD
GOICRbx/0M6Hp3ZAQmvJRCh5W4esQA8skqeqz92uYaphBgj5W599Z9TqOQowV+mS
C1ffWKmHEzZdJrCH1v7MH6VCNq17juR5XN2AOOPEeQY67Gxl2SKzfeVscCAZd3QA
iTy44qxyMewVJEUJ+qp7CTq+XLB8sU0qvbBbYyO/r3GMFZzj/5YuRIt7zoJt6z0g
IdY876SK+U8ZpTxdbNbZo0SUERk6zYPnsDLbaY35DOnwlGGs540ci6xcAkgl1lF2
YwAI4IbmxW9cs+Xw3urPl85ePAV4DUBuyC0VgC5h53Ly1xrJO+sVjkVO6/EBgHSq
Z2S7g4L5tDfunKHIArbg6995r50PzfGpcT7NEHhT6RCkPSoW2+tYesvqRYauG1+D
bjVZd1g286eDkCysx28KVIoEFGTlTuyi/LN9tx5R7nPjZC7VazYYXedBRn7+3i9C
OhPf4LHhPGCJB2tqkO3/qH+2L0sx2fNkA6W2JhohJwvyBGY3VcqK2eJzvAK8OVJz
YXQF+t+7kYB9pLuA14Wms6W67/2Q7OYh4qBxvTbRazlU8Brh/VwKdsW/YwEFH8Mj
uB3jxrHydmrDaxOes1sMsutZsAJ7DbkunmXUnXsN/fNKNM38CzxNev5ivWJz35+m
ogECEHlhsU3kIM9HEhmX/YLMFWxu8gvV44ewS2vwzoOhjX0M6QkUomAM0CvRq5br
n+cicCqd5ZFRvV4xVsQ4W3Cus/nfYwnM+rXjb9Hw1lEApSZEjZKGJnVDh5m4F/No
4pZh/gsRuZ2pmWWQWebFIE41P4FVA1Wk+tyqIpSHSMH8s+7xh3EcVKlj/Vs94ZfQ
HpndPhPv2BZSN4IJPWUH8vNtAUB5k4l/p8vFPobD0VkOdAshgzq8yMocwepp1uVd
Si490BcbWvnXoamRW9xXMyngJfTt7XvIGT/pC83Srub607Nv1sja5hjZYDHbsN79
V3c50A2/NqumoXtsNL5dmv2FX/v/dg0zW8gov4uJGRKuWkgmMpWVEItrEUSIaI9T
voP2nwbyHCqXBy2Rz0JHnloKkr0l0SanF3DmSNQNpcJFdrpDRWoAFM6e9BRPid/u
HSd1jAcN01pv9zM+M5dtJaHqGGzxPSVu+tiGwPvFH6T9pQOSAmspjknOv82NLU+t
V3YGDMWw7gcDR6K9uTqn8xEUSlTLRUQro7tKM1mRtFpqQrNrGrphQy9rMARnBUcP
hkjuHhjxvy5t3ZNX9LZtvbW+NMPkQn/yiwPJ1spm6DaNV0geXHdg+jDrvp6myy6Y
/hHTKIoIFI5fCHM34vGV8kW1vlHe+H+VVydBg6zG2qO2TuD0VfZqTVxVnNWfoyl3
eroFeLmbirSugRrASUvyOADkw51GBZ1WfspU9zZFVeWRJPk1mxcfovxGj5/c0JT8
RXurL23jgl6wVONapohsi9JfrMF9nR30sOQdISB0WXXAD81QMM7hnYHtxGcSYMCX
IG9gNbN6rUsVxxAbRFg4xeyHuASED3JjAy9n4RGHJOl8G9cwcC/0e1XBY8e+fy+s
QA/KiF0+Xrwk7VbMl8plYMa1RerJbkKPH+1WodNX7lj6RfNLOMMUCIFBHbQ4dHdC
ljRK/ZEFBTS6+yO6awkDOH4whrRvitNhDNakUmgvnWWCriiRKsh5KJ1z84G2AQcV
Yw7h9DrrfuStMmjfw3ctM9pmptPIvu/IwkuSanKA8Aof6Pso56OXmY6ZYf7W12hH
18mE6FuJpDXXjRRL+D2wctCFkQniNegOIN8ybb5mKOQbuZZrV5DUnLuteM/zAjyK
xW2t7CdTFzWrnsP/b1FJCkSL9pS60Dmdp58SdO7NSoLNl3CWvlFRzwKZpDThtIPw
OpLezFU9d5JCbv8b8e0KOnPITp6Dl6kwIE854zSs9tigXUgO2rjloPa+IsQAKMKQ
CUmmyjc2b4ZQ+43d03LoGAjvtEN9Tn6p4ENfpFfdJvmLObAMmtVQjpYIs8rDSWgV
bcJxUU993F6Fs+Wbx9c3l/RCioWTrxX5ay2fOs7f4AV4kEaJB+sl7HgiCPiYmhp7
3Ar0kflgvu6W+Fe9eMmk/JB5vB/bw9Ko1ZrXXJJss8xVpELtoVF7jMESA+3/2NvW
86KmluEJ0GZvN6LR0F46vuRULXrWLz1/DeSez70imZfmcKH7XcwwqzrhlULvlODY
CfrVIYUPLiXOqzx9k07wB/DHTbFqFKwcq0pS3inri6eOE2BcQ7EAKKpHQjJto7yF
kH5fGGWfBvOPKozxI+cOv80/Lcw1nke4v64ivfuXvbTqFX/8ldZBkPIfv8AvgkoI
2V87+yP4811DPDnQEQjyvycDmUqgPk2iUClctqtN6bZLRxojFsCmHBWnoCEiDlFb
PE2iTUGRwFP1M/x2IP6fTf1VfbI9xXoIJHLqRfHw/ntqedrZXyHegeCrMmfC1cJd
r78/66PaY8V9Sb0oA19ddyFqdVPv1QF2nwjcm9Tg86fKrXB3X4BXdW+27So5cGOz
d3FBby9wN7uuG7gIW1dwbZRBWjGsAgeG+ts5Oh5Iv31O49rAXCxUnpt48cBYGZRu
zXff+NsUr7cMjgdicjdBK8aXZTFIdIxTz9zYAB52HHTl/8r9N0DB9YFRWaROcvTr
Zx/C/DykAJ9IfLn7OFFjRcMh5ul+vveAdGBK6lj7vv/NwQYZ1oaOehfhalE5R9fE
y8Svv1cYBcuCgQgky9nsUgP5+ffmE54FzYQJzLOqluT7fWoIYvbsbqRyQPgH+NQj
J77321YJ3ClEhyGZT2ZcgGibDzs/ByDseA9qzU8pORe7qq15nFiTDIMc5SJPzWVg
3aGXgb3y3E0uRx6Wn/X6aKftU6hrPDMOQPUQtXrjuE96142wk0PSr+xvAniwH2Px
nBqJt1R3cmnvApSgdkI0n7vjlhNkTJUAS+T0k2RslQKkHMJHhaH0pBjGqG3Yw7sB
TZAstQn62oVO4zy3H/EnFqvVdnfLLlRUkCgSCTPfdvckMEKsR51dh5/aHg8N4nEo
9GknWldggDoQUpb16pGoZyCN0YLiB1tnXXrFL+wb4zOU7jD5+0dameUMXCYmJNgP
whNcw2hCYDZrYWjtx4oAyW2QugJsvNB6zTyEHL/PLC0leh+UrJb9PGB2Bx6e0zsX
VMRXl6iFef3kuVFjf3nWsuIJCmqc3AD2ThVcn5d9HEwEQyOwNdS6sL96h79sYrxF
yd/ZCpsKIpTnnV0maRLtKtNEyN/qkhP3U1vHZvlrUJBgXQZRtTPoNKkTGi1PzIsR
vS1tHtw29RoKpZgkkR7Jo54J19dJvsFAbmhXaGDg0dYMACck0SkHFYlJ/aKNDvve
8XW1DvDGe6Y5YL0kPBtdn/PddhMNj4P8x0J8iHPDK9t81JYeN/6l4dYcD4n+BsDA
JIZgVvV5bAJpxJZHwBB2L2Sj/9A1NL+m+sQ4/yO0uOGZXtpZQnH2WgERHHPX9Vf/
+rc8xFTRPCfUElyrmHaWicJBd4TcK4f0By2W3I6+qLw7Kg9EkhFMU++JsdljD6qy
hT5O9Wfiw8PTvadZyXqnqp6Duc16qgzvQO8udRnaMTNw8r5lfqVl6UhZ67mnYwcB
eWP4Y0kz0PUTew3WA0eppZddYsaCtO+zI1/uexxEBVL6/7yoHFyUSh8Ox/KByzYz
CbN5yDhDDTzGujVff1EeZTCNy2w8PegkvwnyF3wQDvoXzntYkhkyn4hCEg116ewA
rycvzf0+iEZiIH7gFLnDQHqxx3jOuxj11U8RCg8r/7iGTCQgXhipqF/trvtzPDyg
TOi1y0c6SB9OQhVU5h8SvI7d9KMB+K0vbJYPh5LZkEe3wX3aShI7Xv0wE5kaAR2X
DCwdOmEavhgSH5vc1Wy2G9djKkCbP9nIqUUVLa3bnRe7DZadPZLvVVHC1bAH3B0v
Zo3x7VRIYsbzKM2HVII3Vu1wRYo4VUu3Kkel/lmPRzgCGoZCIg6Rzkr3r6RgcYVz
l3XT5zf5ese47/jJyg3V+AWWe77F/Rv/GPha1NzQ1npnGVhJw5s8SHXHNwu96lSB
HkhzwNqLmagiTrHVM5UQkOz4t+yKmvyr3BVmuGW7tVV8CyoSZDZHQ8/oQYwG8Th5
FgoS+sA4rQ1WOnXlHmlIOTFOeoO+oGBm7yOEqZsSR8u4bp/+aVunErvEvZ7DWpoF
xljSHfGVyfhDY7+O0osbzsmS4ddbC9ElTm6+UzSeEb2+kUbB9GOXQN/ZrUipmQ2M
FjhO9TkHbSka/pv1pOV2TixphIv75ztLERa3ziTEZ2EpFcC3Mbbb7auWYymDrq+/
YB0gOF+Wlr2l1ytcsBOApGuUgKLMgx4ChZV4doH2vrl1UAZ2cTBsbnDB9t9wNoo/
Sx9MTiHLg72DyXskFNmFvS07agtDC6hzrzTmh8hPs+CAZvbwNzDS5yhLKyHdoj4x
0gh9flJB4uGqKo4Y6rfIvPAugKLizkCpVlnK51ORZRzTvTYg/1p3dQ9hFvZaG5Sn
HY5xKaxw7GkI4Zly2iARnDKW6QnhLV7JExxvcGq4ifz6Zjdi7PVfAJcfm87ehlZw
Ay25S9K7csm20QnRw8RsaJe7qgQKWez6z+Vn03ECMgi/9JvvFYE5UMOn3Gtv2Wnn
dp+3sTqXUrIXobX4JP+iphNDFWjiwBo2YrZqkaiyB2x5bNuQddZtuAYjtmAtb2vq
wjI7fHCMBih7+H9iLjrVq9uCOdPTIJG4JvIY2A1tpcxPSATf9GFjNZneK90+TB2V
IXA+nQmwG5ZndvTvKe3uL/TVKu+lqKtARWloSZnvotWuisJ51wnlnJj868tuyJa7
t4EsNtiGOdbQ9Iqrbm5iuzo6CUhcxWB4ffW2JR3yFz9eagDTl9a9tO0Qb/dOmpp1
gNNpTTXWvM5uBbamncyU1lenWo11QwEnkAygBa7OKqjVhzFatIJ3XAUpnQs4v+6d
8awkqQYJE4GXebm7BSH+PoiJt+ef0E71kmr1vaCUfLv72ntBb5t+EgNGUqPy0CYc
0AEp5qvfdWyc9r/0UrWyeSfYq/cRaddPFQhSy6J2FPXJag8KwtS++j4Ps4hiZPHn
JIyVa4y/OdcIRvXXnyp0wNVsLvjskT7uL3tg7fFMUX8CAIWwmaJzNpcTPENkWVvy
lOf5fvbuJnH1KGK7G6QNWBm7rsC8ld0jUzJ+X91LfBHhPZAHkHibtSiYCEEl+vrs
8H3HdUkO5zb31eigbKptYNBokHz0uBsE0cKY5DExYndxGo21fpWCoTMC/8jJywnW
yGo9+4LoQr2ta5h3LvDxRctk1U0/X+DUmgXsXCitOK+tld63CNfhOnsq+WoPrx/U
DkKtnwo04VNoEnXIBi9QwOUHpaRnnkMKY1H8OOBBT08a3jV0qc3W+u7Ie1LaPqbc
AacG5aeJKMxzOcKNEN2tdtp6RhBfzHYxp9GNlvB+OMJ8s3KA6k8cuiN6MyNMcY73
kmBkg9PTqYpypmLdpiZD8++3nnRDWUWKfIqNPCzgi6ZDcXvJY6eJ+FYYIg64jC+A
U6bPZoAYnIKYCdMp+gxj30rcBWd0KGqgty5JPgWNJWlaVMbqI5/w6NzCx22qWOoA
rZdlstKlqqPhc/+BXeKnxKUiurj2ezrBNY+nzqH2el1W/KBFD8ucOKHbxbBFUwJA
MVxbbvuEvwjnMki4VCG/+RZG+lOM9oebPjX3Ix3hoMTWX1SXg8lAAWGVNEbvBfvW
vceMoX0k17RFf6o/EeKj4jEEBWqdADBJMnqRgPueRcDU2MyNg/Ppc1EYrA0ull+G
pmERmqonc3gLZTO+YzE29yl5xm+/E8pBDEyjb1OKSl6VqeYOsj+OFJunWZxSDp+z
Q+qsfFQyt0gzo8UvO4s16b07Fe3f6spaKY6wOp2z/+dQNat130jGVbvZS1dn1pgw
DMcU9OZR95RjbMUIA/TVjikgoBEL1+Vkjya/qLO+U0FsaNla34PTmn/NGsZDgJVE
4oHF2Xu+gYGykd+u90QiFjGtnheW8GyipxF38jzWSfuxS7LIB0hE5xvfn7iybalK
Wuf2SzHlD5Imoe4GFSZBtch1cBiyRO+4GYripdnNvzvad7yTMgRFOzqEhNwzlGay
twu9Ltlb5eq+G55UBMNlH89fFbkiNEbfYnKhelR465uHy5+dBFNvP5nX5iaHAVKb
YSOANTSPskaSQFW7IY7Q4FYox3Kixd9wVhOxlL4mO+U18XABX0O6pHzvV8yXyPEp
WnfanNPMPu6zLp63uwzn/h/er43qXTtQYPRKuKH7LjAgfmpW83oGkUxJtRicSH53
jRa0+8IQYQhBqo47BAtsSP6BbUotq4BK2/2bsxS/E+Pa/CAozdO2FvDbm2xURBjJ
rdM7+LKXUah5tfBHYkXv/ecFnRrLpep+tQAaFuohmCLjiCISg2yn0YSh3vRYXBsd
YKgVPPCc60k5wDoQtePiUn4Oj3PsFkC78emZsr9FmFdrOBHTYY5k16bfbxlfvodq
L4XGbjImV0ibIlxUdo6rrQjjt0U3EWviUkSvP9P0h/V0snsBE7c/JTl2QFW4nfj9
jWhuXUsomrA81VOHpqS/+xEkr5ObT2aCRU+qm3mgyeJfPIRwG0wR/3UHSbohC+T5
YGVa8mP2MgQYxq39y6pMTN24LRnlZplpWwZdHoyBvdNb5I31Na2CKK8IkLIrPVri
lxrN8AziXuqnGF5VEyUvjP4oc80gvkTWUwUbLg1GQ3qDwOptwmORbsQs/ynxh/7N
uAamwCYsSszrYJHu6hiVxHJ0Wx5yOyTwsC4B1WWim1PkYa+e3McnxMHC59e8jlLZ
sMkAI1KZqH8tdBOk4ht8Ip/1QsRUxyU2zoPo49yOFryO46Dj0HHl8QCscxYnbhk6
AawYGp1njyYjijBEQT/2kAGfoLtoPWAab6VuyRBKPr6kVKih/GGCiz0oLzw/BFZe
qliWAznVZRX7/T2GTbC++P8ADCSmVtOej8uJtzv0YWThIpSqFtJqp9FG4TDX95T4
ySiMAltAus94YQhZ+jau9YW5Bzd6oYnLOvDQ3knvp3Xq+nsj54wQWbOJQp/JcOpD
vnfpa04XBVf3SxXk9z4USkUazS3NQsU3DzitdnGopvddpk48x1RW2Z16PhrYqhNy
90DDHECh3JYUkm97e6Qb+z3v0DTD0UIUYstmGe3rLH0wdvTA5ptLsKiFiBrUym0N
QjUPEYMHDhK4lzVoFkNEs+YZhWDvCbAaJSPU/44wRtJfJFPxGmBzOZCAAIVZBJeS
Pao8SDOf1ZHZfjpI7934+3Shk9C7oVGh4yG5nxhLZZhqA+MCnS+V3QNh6H/ZIK2A
41IYcajDhjLb1fzdwpz5Ns+bHlcILDDAjgl+BU9xnBFMew2Z8H5olTUgtr2ig+ov
Gp/uP0oIbAbaZqm+460O6QIYxw8/v9R2tddG1rAvwnLL2xmCOipVypHwIXJ44JPs
p8ByRDtPYpaoyrHNy/lW/UXIOaCY/PDmlrTfrkXDBjR4C4UKIxMD+E5BKX5tPY4a
rwUllsqa3JHhSTMQxmAIGk75svGzRK7UiD8oXQCiuLxKHfAX9qK6GWC2u/EkpAF/
2ZxL8hECCuZvZb1nRTEuH+eWgGbV/PD4EnVKKh+AlCUzGkgSAsIqcpP9At7FwRUk
DJ94ks8NFjQRzGN5ATTNLHCHjXfTfw4ZjqgRSd5kzhLO0TpQYeyidkxA+LHBDdN+
OKQRFZMZszqZWtLPIC7ZpTwnSruVunrS2yBOqHoSkzBD9dsorjsPdlsgp5G7NnXd
RPn6UgjsJlbETXtutvwH/YQD633FcNX8O9Vt7MHxwjQQiMUnHbloTmNyxZpcfBPV
zJcX9oer9ecFFbA+dLqja1EgGFQn0Re9oghA6miy5zFH8NVqeMEX85BGz66yuxm2
4eE1tXTOGQRDtvz/TdyFogGn+ySOmpcDnD7Bjgl4W1s06+wIQpQrSyvEvCOvy8ii
OMFTY6GdyrSWBaKRapJCiJ59P2D4cjpuay68hok8+veRMS3JnPVGvxThirqxKRhr
plniv8nUWp9ouCqolCOVmSOC6dhSyrQntZBsWI86vNdpWqFsmBP2bhD5KcUKgzoj
UlMsicZKUHlQj4gDpZAQQTJuLFa1vchXYRgDilE74DifV7slMrx5W6Wp7KgQah0Y
FZbrBGhKDS0HYP5K9Cj4Y+VNVlXKxCsE9xttNcFAeBRilX/BaWQmVWKP1YncZYqx
xB+YrdB/zxpB1snkNsQILGjBMHNal+0W1oLfL6p5qF3Km7lN3qgdOd7PLGsMKrYm
HbeLIiWPXUXvOt3g6hJJao/VmKYc6S11VKCPz+NMk4WBi8FeJySGkNpGV5jBzf8t
wUxvBTeSz2zr0jL4BUoRGslnp7zaFhpyHcE1yB57P3GZmuz1oB9bDvGEtMDg4cjf
vmXMQisjCpwA/Z4hXr8Rj215pSzudTQMZWOduYn+eqDMrX1hUI9P7qdpp7nM02iX
3PdwvisWLPPDG1SllcVj4E8s+Aa4wdRLps+5lnke5sE12cyCaRNxf6NFeELfUkEH
R8q+I49QEIXUKIawrAPl6L91vLp08W92e8N6j/0orOdZEY0wUSoTvTTNy9M1eMQt
Ai2IVJ6zaEE1EMWg/Jm+yT+ynalhgp3DJG/vdk7JgQ3D6XQqWTW/Vmst4ZYX+YBe
GpQR1wB5uDYuWVAdpkz6BRaslxUeaY8QxcBFQT2ETjQQ23Bb6YQvmWbkJznQD3E0
4DiQlx/DXvmi53AUmYcSsw1l40ocZqnc/cmeDrqVcCAwNvcHlwRgVflpMMi9hu2A
381IStetV2IRGO+wQnT++jsMH5llFoswQm3GCDho3dU7h7gP6jyPzU8R9lkCYb3h
ZVMzDvyFRqd7KUfKHk+g0zm1kwDg/cLJHO/5XmpsMaTnf/4d9PzIZi7wYvkWQCvp
K20zL8jgg7TzWBmMUwPeXWayrr0PjXhfVAbbHUqzvPv/LuDwf3YqFV+nlmnsH1+H
bYIAq6tFoFkMHjEYVO96pQU4wYT2wWA0gdWqlvsTVN+BqpmkAY9t0UFKRqDrGCM3
UzOdOcQgInS31k9250OlvTp7Ds8zRw6R58WxhMlLPMSbm1fDpacbC50t8pljyCfW
Fy4go1xNk9lzYk1ILT7Yc17RdakSPAXTMug/8s0RcyYztNSRVhUQTHBZPgZC8lkU
Dhfvi5goEYKSlCQrKVsEwDq2ct/Xnum9HvkOfO2RT5e5YhuUrQhes4Nf9Zu1vx82
UJfI2iprP1C8Hc/cpCBk4BZp4lVYxnZrGTxsx4f8Xs3xx1WADGsyZPxY9rYLztnW
eRyIboycLealxvoxobDNBWKNKvk439dB0qoNY8XdAfVoajGtt+Hsmhd4eHAU601z
dfOdBd4rpdZ3l5n9g9Fh/qc7aQnARZnX6hXaQbZdKivX3EHdq4tTMl2+FqWq4hec
w2QN8uGiSOQohaeTf+0U3ZonZeSoo2UysF1YeJ+fXxyeAZlOWtS+mC0gHHr7gsmq
Og+34J5DyBgTdTb0jpWMi5ktB3p7WBowQdNpqD65kmyHwpsFzbtDaCDCpQIBpctQ
qRYkYgtn/Hqhpt9H88CesSPsZs7qQPd92w38x9ygo1pYWTjkLuawEuPuIHRakdWX
37AVpQ5//AGkl4HKa8QKzfGzuHMQVs7OrAlIscevkA55AssY0RWAjudjiPv4wmze
2NM3V1guQMk61XiZ2pkA/phdfKJj1NXjRk/fuL6F/FhPAMdTfYviY/N+NzMc6Bq1
XHQhuLAZqvikSdwNqKlyjRzhajjKpDMDmC2aNzY6wXBa82L9+PB5/k9By3jTZprn
i1hHXGcstnRcH7eNAmOUW3Chu9PRN3xEnHNdd8wrOi7w3gO2w0/OxHSOm0pFeCH1
3b8SSD2XmhmpymscatQ1JFinGpZu8L3FFdTPhgk0/eOnUOBIksUh4mV+vdKVpnGJ
QULG7PnXR+hnGanL5rteKH96etbTH58rjwomgGfZdA0/o9s/HVzds3+W+8CXT3KH
RyfVusiMiXw0btQdSWkrnnHDSxZwmNdCQP/W/tN8cbh83zVlhvLzjwqxLYJ1Zdvy
itvAIO1ArpGvwOnSJTIOUJffrXNJxO7kY/63J8g1Lm7HlFhxA2rshaae6rcJhMz3
pXHmOZdFQF+ooKmneVbQWUrZuEpQdMX2DEIDq7ZSzj+OwTqP+2uPQhkLKRBVV85n
+m+FetT3NxFJoRAWGJSSsJaWukQGpkMGke6yWD5CdDoVda23KYWUv/MgeY3oSkXc
4k8FRoPe8B39Cz/2f1cgjEBOrcmfVN+7XhJQXE2mCyVAe81MwNT1C3d3P/m5nb/c
eWyGUfg50fD2L/X0hSISxeWpC3fiGRVLo2iGE80KN0E2SBEMsuvALwCt07JrgXV+
XF/Pv10BnAUTAS+0HhPOIlwzOkMDF3ZEE5j81jnSn5H97i+tMjMgQaShadh1/AQf
jNUxz4Mfk1zBUIbhZct5xlbh26bCuKZM35JHGDf0hs1Hcxn8Cw04r2XhbD0kdjp0
47IZQtW4ytDGuZ0ihCnJFVVCBndhhRceWWYWRYIg9gUFzzT7M6pEmujpepa66CfX
+rekc3o7n2cRls9l6hIhvVjJa0O+mPIiZEYiq+SjGCEPrRtg/4x0ddy2fCrrdbwH
AVMLD+Hqxv5ty0eqLlfzfag1zLE1vpy3lX0Vy2XqqjMbsBM9d6x1Mm55wg+ood/6
qD/xuQ1b7rSQTJDMdfyFFAEYZNPuWp3J7UGgLQVKCFTjRQeyYRmkVol2cDy6zq2i
6mFLNNzkU2QVvGFMa8x6bca13tiXuMzoTuQPX0Uz1wSXfQ5b5pGMOGvufUgyIei+
gn9c5fRFbYDju31sqVp52OD5NMl9lXasGhPCPEhTGVKHrM70ngUN7YyxH/fRQhF1
z8DeVACMHI2CJmi7PcAGkgxcbjnth+Zw0eLHvfEvduqGSj/17jcF7I4Xf2GPtoA8
k91ftY+ZxW1cgtEgWvrfDmon9Zymn5DaDzT+w2I1idP/WJQ4lRGc7oUoEMiXi6QK
Mg6Bd9qZuTci3xcoo69A/nO2hSnIk8ujurJTuWgTjyXSJ+LyMdBoBjdGBtgc67Z9
xTeYwCp7ZZg4roQZ3hEdJ/LFCmoxiMLzZPsRhFuRKK7MjeMCvJmNdERjOWsc5nTl
nbL45KoI27nRXS6mp7I5phC2viJuqdfabxI26S476M2sTTY98nR0uKT1RvlLwAY9
SaGPlWgFllID/Fk5vlUlpJrRo/UWmjNfjPcweUp0ILooLQyVPlaBqYkjYWEr3SRG
8+wiREweGQRIw8sOBuVohPDegT53sgXYxKOCKG9pQ+BoEvHMHP/UcEoDRLCjm4rN
6sSly57tnUqyEcwU5ryIfAx+c2BjlsMRDHiihzwGKkmHyFKSp+M9x87G8fBgegWl
txnlZjni9Q+g9Yr/pWryxqTC9O8h7xa74xlvt8y/4MXFmneCQc9zgYj8RcZwxZpi
/PZnNFh6FIqDBBFIbC524C3L5PLmnexyG966Ce48buEck4q9fI1hdRkoWvlJD0fV
tFSYCDVumVp+2ByHj9CJ0hHci5sU1wZBI5WtYkfC2IuEmzxQaAmTmxSPFIY06NL/
a3/MambqdXhyYJzYmPkDDA1YyfUKq5gE6V1NSjd4N2QSlvIfugK1/dMBInj6au/8
WuXgrDs0Gq6k+0pEjCKxGZ9l/BDoHjj2OS8vp1KHPq9zetSbO2u6pMughMS69uDL
NAHyTgegBoCgQapVtz/UrE/TnGvI8H0FnuHLTMvcls3/6zQRkpD+0yrl20Yw9jhj
+WdvDFVw1MsnGziOd8JR+VffPZHwjJ89G2uyRPJyVImCjWdwF2GUdQ7WZKmlM9tF
upDf0YDnvWlJGyQ0hz9eGszlLKPY6ePgRVyti8XzUGTDEtKRrxyVP6EaSkwm1X2r
+/VYLaBOuQT8ynd3EpXQyDlVMN4KRCEiH+fwNWORjkXThMDMwEDQBct0GcXXgxTw
+aWwgdYrBcRFb4HamzD3B9Eow1I25dK40M6GogA+xR4vvVTYOQ+UrPYEOuQ6l8Is
vtj7PW/v34+wjNyNm8vJ7byMtjYdoKtYAMDxCIM5gwRSv76gG/B7cKhDcr2gRwI3
o/8ZyYMr67PXhRjBsUVkEavByGY+guat7bmDvjQgI8Wsc8EHhTOTA5aIKPJyFXRh
hNMc0B6TDDEAOBhML13nsENrJho8ZcyONolYgJeu9O7ac4tKOfXTcr3W/I1CU3C4
U2LLDwrY4Lcev9ksBhvPoVt8RVKLN2eXokzi+ipj2sEwPjUHzHCbTNNFhCz8v/Np
nyjlFrz3+UrYCMrOt7VY7iHqu25rNeDKw/rx+di3TbwDQY9lDNjJUj7dETclRpkB
6STbJs3Lf8FD/VMYP0hoZjpmETZ/9BgZTVYC9wJyVYnINFsisRkg2ZFf31VeZJ/Y
Yl2m/1/Ocu3K2CILhFvOYtpa6Z9zKk/mXjMmPhDQteuQjikbT5scHvZadf9E54la
e2CqSudX0EIGVSlvCOHSx0u9HxpZIqW/7I7PpmfiHWiWDQFN7yjSe8Uf5wG+ht17
4xVTLxXopBLsXvPeVJfP3fzrkfEfsYTdcyG4z2fG/ZOZkNaBxdDCMs3TcjvSq/9f
dvoX9zIKAO1nlpHjlkDaTzgdxTH4moEmbeDsgOoLmzgSjUw377eltPMcrXvESRbN
hSEghfgdGNXE1dIJtp0+QGOy5nnJGTcKzsEDiBqjHBBiICq7rkCVagL5f4jYSSr1
iwcI1xcI7uMmC0S+K568i1mZxqLG/fw5tyOyHzXAGEsVqX1f8J/JOS7rK/CbUvQD
SacGp3FMsBup/NJlaX6NruPQMqat9ruH+9cnu+YWBfzv+ga30PSR+/+Z1d6bQ+Hu
y71HuoE7SjzVLUgsDc6EFYq0gN9irwI+z7Odn/CvYxW938qhBHCAV81PlLlxcUAb
o7Gqu+KsVU5RsXo9Ta4ymEK/OmRNoFtdPVdF2YSEzp+vQLmsLRm7B7Qk/l2AX4wk
YkOoQLPQF/naafzTC3P9cl4JZZfcnX3fPj6RQSG3zIauUBtYjY0o803znaNTL0zf
km72iccUxLx2AharDtDnoB/pH8IlYHEs+/R9ChQYdCrNEMFYr4aTNY9k7ONNTmjb
M9DOlisAFPG1kshvN1KWgrx/aiYm7YuWXD7AXrTbYSLkDKAV8c8LaDVrz0KNWfRW
BO222KVUQoAnr0A5Rn70uilgjO7vPU3ZpoRqu1Hpl8AhTwZtFTDZk/gceEGvjYgU
ur66u/IQSd0iYmZkSUkCuun60G6MryXqv5XARGn/hWp33bO2XfsTRGqPc6Ga0Uv0
Vh/4UQmcs8qx07Z8vhekRz8lnhcSTcX68iJwK0Mcx66RSSd65BfbsEBlMTg/Mctp
ZJjkT/MsLTb2hCNjqIq4DrXk88NSmTZz9BJwGjB5gHZLLVf2+919ZJ79rWLyjy6L
TDTOf/SzZLke25zr9b8FSclml2CYi4Loao3kNV4A5k0wqGV+26ce2OKV+fKcP1gl
hC/6xtChkXLNmS/QoAZIt7yAZhRyJAETMeaAP0qWIyaKnVIWsgfbHWXcWRV+/77V
B+GccpCyOWV4LKRUXjJDn0rKHa0hfDm5ZKTGgB9NAa0zUq3CbNBfAWI7dh1E1Dmv
FpKRFXGjzeym+umuYebNIeoxIXlIYo8jKXP+AwvNfQt6RZD3GLDoKng9UeWBTRuN
uCcZUkMHh4wRJGI8OltGhYi+pTcI6tpl8xsGdZCgxFYV4Qv9RDaUXWd0AFcoaUyp
oXwiol0SbOIiN0BYGDTJvqfldgdzB6CPvWQNXDdXbbvLdPWl6jYNGExVTD38X0rS
9jzLX+YIW6+D4FTEV/f9rSojMjU/PG+ix0hHYhzs6ZekKMx10vtWJQL2a/JA+GUU
o6LOAqAa7yyNv5yH5vcQEclWhIzqY5mlQWyBwZsi6pX2/N5KoS+V0WSAkxFrH9MH
g6tajGRVheLCqg+4s6XxY8vlSzSEtXCLi2AXF8c5YRq6DSYe2dWNhyemYNfpnQGM
FMviFqD+jdjvE1tKJvO/KDWpcDkRgxzkKscN6M5iOKWDgR/e+ZCaAhwp7EWZLQuI
oC2kmKlMIvFVw5bEdi+IrSQ5wFPsaDuecMLWO7+u7Ptiio9FtJegzBDGXec7IadX
q2jd4ejqcXGMJzx1yMTOTEz76D7022QcMNaRATz6/wMYYX44V33UThH7hbPQXEc/
zOcT4CbadBjEdXZSPOQ2jJoJWV31yOF/SVE32FqBE6tZ8dutOq9rIFr5JJfFuShy
gHC1PVP5AB63SCT6UEQB13tf9N3ZTSle3jUkTYgCU6rFpv8JrgMiVsOoT3eS0aTg
K25gl6oVSybhnihtgZE6hbcxRAUCWqJDq8yalccwXTbmcucw99hoiAYpzWdfzai6
HaHqbk+7I1SEMANaynOtstVwGc9HrE3bk1XkwZidmnh4ra2zqIIOLcn8mpygP7X0
NsSvMkNbpi5yAqrTnWnyPpSVFhf7TY7hNZmyTEVX6muyJwoKanClAQLESfFJl8r0
rlDuiTLb0ZBiBNj5M31Qw/foF2NgADoEZTSZW3oWGftnZ2o/33AxYx+tnkXCW49/
uZbL4rnPZK2v3JCpxxHD0FWgx6akfG++E4sICNuOFreYSfil7ZvaSQL283bRn59o
XwxIbvdIkd3EbDOZydaTv0na8XlrNrOwEoyl0/F3kQZ8XPTRq85DZsSjKEsslNpC
xD9tM7oCzGAERIK7lpSGDx/2jYgr4v2TNqRta2rs7dlqdkDt+LYgP+61zh9GUD1l
Ck3/55QRglAEtHiDj21M+oWh14TyBrSgy8VThHCZ2urVy8r6C6bFKRq8atB1tZmB
4sm9Q0Sr1dmKt62RAHLsxgggtBTt65bvB1TQ9VazPZZMkgBS+uo6z1VVXAxc31Ni
iAwCw2BKZFxz/DX0f62XusH3yPZ5WXvuWlwu99xJ9I0N7S+k+9fqPfdkjS/6xEAE
ckpzSpWp9+jVxXP5nFDpqwOV/sdBB9we3s0m770Jae5x1e6IPFZtGuIzZ5JXuVqW
t+2RalA3MiZ6av//8gI2TGdV0ss4sxQgPl36vdcWUh+D87zGStmRu6ttFGxNF9Vp
ukE/PFtSie+mp7Lb/j/RYXPzwVc0GW8PeyLotxE41Z+C+aT0G7hV1lCR1RvTJeFr
KAue1PtiLaYWLcNpjj21fn8YQha922oSCSd7hlPTjkKppauSkBAbdYYMXOPdm+oQ
B2c/+5KmoyWNqJFUueBo0IxDUO6ab/WYqZhlZ69g5EseaXMYVrLJDcaT7bG5ztIn
Fxsy5eHeFrUecMn4K0CPiIsGxZpe7cpWJdwDzPYB8i2QYi/K4W+tSPttCnnX52ov
uyyiXs9aEb72tZkFnWNo3iLXiKPGRMYRR+9GNZ7ET8DjIchUqht4V/KMQNmJrnzU
KATLRfoTi/HHlFXtYyzgZu5M/KAA0KPdcPaphqlmiN3f0ofh1LCaDZt60ijn4Ggn
gFlHqMNt3LUbPutQBHkPXmB7THz4LOe5mmPayUqn+hKJQYp2nDM+LlmYC91AA21v
1W2wUslHy7H+wPYKRAkPlu4Y4Ff3k1172+Ix8IM3fZpLHs8X+eBoFpPNmVDefwlT
NKNSkLhWdwCAx7RZ2HrciIiaq/5OXcROQnvXQRa6GacfbG59XIstf4E+XhguTY5E
pmEvwISkzLt13XxSFh1jlYehx5eHZhn4OilmrWtCdnTvz1ai0kSbtFn2fR14F43w
wRTvn1/tppevpY/0c+XM/jIQDkFguEPhD1ccQ/mNokNnHUaZB3tC9FCaRLXVnLjp
I8SkkaEzWM9CUZ6IOtfPnWcOqs841bqQB5wWx046Si74k2SAr62GxKwNoyWdHQi8
mOw8NZDGHZ1kcuPwqFRny1q1WlsQws/3/TyQmAyfAK+6d2PVs+JEZOq7c1QnTYBH
mthPe3x4nIp072u1XYd+11PpEdUgugzt81QlM3jWRTdxf5KkEFQlT/4y+mIETo6u
PspY0JJ66xrniO7X4bd9C4rzwE2jQfJRXHokIfzjy/tH8rVJ840yxLNguGxuuPam
jVw2Xjs6zvGcxan4HbGgRiYyziVtRhGfQkQTEAsAHDVN81cz4I5mxBEwpWOxyO4+
ipA0cmqREIgtMsl/3k41P1hJjXU8HRICYtSn35TMNZD5xeZVaIW7dZy9w2SN61v6
nk/eM1up0Ej3+gZ+7qgAjUvII8SR67iDU48QQBLZMYpkrYgs3Qvs0nMWkOxgnavl
DiOS/f8FyY7HC0mwQV0CEacgU6HcU/zuyBGeJmPYhs7GAg5Db82bRsQi+GMYtZ02
9oy/1Yd0oNeWKqMVLdmQInADcqH9b9Wv1nSfbStpSj47CtQFAaBXTeNM0ZB36tcW
3q5MLvPCJyIBmNtl1NUkqRGd81/HpRS8DgXgFGkBNNcEre0UgPVqpFq6GXhq5D8a
A/vQcyJOlmaG6kHx0/1z9kFpP/dQ5RZGMDsK22vTd9FYf97FwFBvHWnXohKv3mR/
RyHb/WcEx2rImS3PRA+sjulvxQAlFKBwufPo6/yDyYlXJAEF945loFQHle9Onybu
k6DIC8W3g8uFiQib8bMz9Egtw5exxFl7UI78CKGq12hCvLOHHxvJ1GdR9rvVJEnr
aUWaYE9ygoQF2jr2L2jOJ//uTkvI8XUX5yAgNTCh7TQROUYvQpZdjQgx2r7uOiqB
BEgPu8MHD5Sh8MM5hy7AVWCPTmPzYxR4gQQ+aLOyBNmjM1yw81HMkusOe8WdtOAM
PW9zKFUlZWoijnQbC1nHBYAWNlHJKyBHAKy7FXupatHO/9KMEBJq31Er+ZGov8Nk
S0wJekG51e3DM1pEC6McHmHb82KCW1hsnFjsCQMDdsHm50zfzOr9v+XBAcw3zNRg
xBg/t0tXTh3VuSaxeqQmLrPx2BTzREGBk2Z3HIJE2KzJyQCGj8kt+3tGf1uNRYlZ
s/i4tRqssBamShiughCPjKB3pS3673iLXSTMaLODgw6/9Jgcb4A8REnfX6HMOYii
FrevhO1t9G3tYwyPq1B+8Gyy0gdJ+iUeKWBkPc4WTCE+AIyRlkVNO9ob62YRn0Bb
NhCli/Z1WgIKPCuv2mZ6OPSVyBt3BRawAaxtgLk4ZS6BJ5PEu5/Qk12t+DGDlSrw
CKRjuqLZoFCsoRYAlmrjSKVCV58luzlbxjwPn5WxhUhu54Jw1ZqjSRds1sj+XIqq
ZjidCY8/kO1d3V320B+gx0N0IYh2KZ/bu9Tz8G4s/tWe4gqEXurmnU7Cnlo8Ef+u
4ivM7yCFfQXCI58E/LQH+tCsCNRn5CPqHvWzlg9DQcCJSdM0UWVpcRGLjHQqrt8k
IwWbIueng3vX03J7O5iVZVUROVP/ndHA7ptqzHhokEuIXYeMvt5w7lVxEBKFAjGC
1eHsq6LCnXPoSZX//PMvcFTXsycjJyictpgvwEKtel/8y2RM3MEGAzTGPUEMQfK1
+63lrijnCDYNgxRY9BWO868NRojwu9cwq2V/6ajOorB4uMF3GqjnKJiM8Q6jJo7z
Ii0M4uPV5tSkFq+0dcxqB7orWOnmgUJp917u9+o9sR0M3RIXz2CRRjecbzpQTtGx
g3iug2c3HqSYsuBXeSFqj9mmeK17j2/zD6o6SrBKpXrKLWjN9CiZGYV9qnZy+fM9
Yc3dbUA0aZpSLCaPC4MgtcT5JQMGh3GqnXGi2umPLbMPDpyFxxmt3E34MAY+L84b
Xht//LD+YEO9LsBD1Uj1CNrIfdWTEL9XPz167FY4jRKbixTcV5IShUe7UyTPPbV7
r6v9zFiY73iAhgIWJr+A+RqRDwV5w3Tlvj/Mg9AwbVmZHl43tVAkgNnKQShMJhxD
bmjB7PZxkMTdJ1ztQvVbC1pemontJdav97NZjUjZjP9Fn8u58rM6Hk/L16zKOM4h
qxPt3e0JqroSzuOBbdY+ATH9gs9c7Qwzv55Gk5z2OD6tztm7b8NeiUzO5wHaDZe/
o7i+t0Din+/5bzjITlnnB1zNBY/mdFn18LJFt34FxpqFxQ60nAJdf7R1VfSHQOnh
jVkVlZR+RJx0oqek+9iV/6ozmMMM3aVOjT4YdCICDKXmKe79JAG4xYxjavarz+0/
ECsZDifdrqPFekpK+nsgnrnNj24y6tjuIT9323Ec1vusoRh0v7mWHtl35juN00I0
mCu4iX+hSOfB6wC6Bh54RcKVrPEIr+uMK8ArttjfZ8PVlD9zFF7Q8YdzdBQcpZS+
B4ucg7zJQdc5mztFYarP0n9IaPk3sMWYMoxDm6Rdn4TbkxOKYwRM6ZpPJA6cxcOl
oKiNFitsu9yM/hpQFgCBdMVn6L2kBqIcdq2/+pfw9k03oqNw19l4no17PTW7dZZY
iwTnyRYAlNn7H92JExnzpI9W6FCT0pw3YzY9+QCU4+66Moh3JaX40yh1LFCTIFEv
sDX4gospeJ1DQPd06ikGaSv4gRjzSvgaTCRyNAQukvVJ+0O4nTr6BTqu4y/ISxAJ
IhmUepdLUQxgqsElA47hZFdIC1uSISalVs2Ao8HE4aC6C51tqy0O1QVsolaFoRB3
qdu1dv8sCr5xn3TL2SudcGzR6p2KoS/9TloHgukeayyOU5cnelVlblixRtI/aWza
dcslS5gFqwhq57lNYCzIZrbcQQpJG0Ufcz0xWVHNHVZlFS5ZsIvWPhqZS9wA5Zls
pW4pqeKEB1gKNgksCww/CWjEJxVRovK7DuYN9IRSQqvXr+JiS1B4GzH444P+04oj
pHC78bAxBRNSnDM4cdJK3pQZ8kXyrzVBEimDs3VEeIF40Hps3jg7WwIwbYx31eBg
fiW4IO24t4a1n3s8Bx0DCUSTUN4oBNNBzcl2d4nt/uk3cgkUJs9DLGSG9ibABCKc
sTa1gd1wWa1PkESTcaqDA+g89i2ixXQ1G9rwgZEwTu1rWPEK6AejvMRwQfIKU+8+
USlpYZ48X1z649Ceh+vpl8xomDx8Tmzjwy/RrFOFw3wddL1CkOc1yR5wzsljZa+E
+5Wev3S8GtO41Aud/b/h46X5Jul4RmLoVP1WNlmN5ZI4WksPOKiBoWTD58/CcRtC
sdGnF8biQ+B1qcS1zLd0hhcsj51T79p9RouCA0gBsaeI3E5A+nl+ZxEYxKEycTIP
daV8ILYx9uDayRt2c1wXUM/grOscuwT7aHZKv7wLG4VaaxWTKQ3c8v7C08U328/+
FSjS8q3YXkpzXcGlFkS9KdkKQQIGlbsdYcX9/XLK/ZxO1hY/5H0yyGWxZRw7sVZF
rI09mvGvcFsz2jJkXX9dl/BB2LG1nbgzLvrOSXUhd5XSzEMIgf6k+kdztDAzcDKf
ZMhlnteHr6q3PE0ppKXwBga0t+cndVFmQ6h9tHtsnZAUGbXfCPoo951gZ9dP5BQ7
q0DFK3kYGuj5cJ1nAhk+k7pfbG9Svnrogftdcl/5DGC057A5S6kq+ST6zGraJvLb
zWxBwCQwanYu/AF5Bffi2uyxQBLZSnVSuYG7Myitz6fyyQBMp7y67Af8hTpvExTZ
LWbgv0t0xWc+41UF93ZR3OI4JnqeuUtjybU0z9B7M2WojczuZcZAogmP7oxFS2hL
Kkc0DBqyC5kFWjrPF6bHSKrEjkIJYV+XhZEBHfvmxD9fzGFAMvc0WolgsGFzsael
/nZzjCDuMpyYjQ7Hgb/DaFsj7csKEhe8xkk7cJl3u3W2jRhkZns2mwM7DgxDsW43
k9AcHS5ItwDKN4wNKfrlusi3gw7juN0hw0w0baR2cRCe/u+fMNmZxwUaKFi2RJS5
fLIkIp7TnAUgQ5XtG4HCrIwpGN1Q0X+Z0aK5oysAFsHKvVKvIkqGrYBWL8lC/ZwX
ZdKYwLFnB91Yq/QL4IE9xVFB99Grk7kNQrTTzLiYwrq2G1PLnc4ueqzW8i5Oak5i
o+hKNy9pRmtxq9HyXy/FPJH8EPp+OjWX2TfFA8wcUjieCcJePP98D2CyWfwqWyrc
2QHZ5Mi4GZ47cYoBzUHZ5Nih9AxFZjrcKhyucJ5fd6g4jx4OSdsMu1yvMLdJx68j
cbw7dSwds9c8n8KbN6Mz1gdYSjdXYk6qI7mTQacaG83ku7b6HRqxK9t5QGtF5RYG
xKWdvONg9NbfbZ/NqvwIR1/MyV4ytQx+zDzUqN6xMWc4DoEQCF+95a9B51Fk7klu
HxzGW6CyLtU6j16BsJgFsxRWLpi6dD0KMGtAUiJ8blq454LqkZEuKRvL2RphbHsl
/6wr7WVXLbZuGNNMJOma2+4sXsB2GWgvcq7v7xrZ2xS7Ro9Zw1+EiI4YmkaDIAp5
0BNHWawdKyDstVGrxrpjfF1D5oTcf8svHrDdCNshjH9kKemQnbk4v8UKMGXMY36K
7h1XV6VWt3n/+41RUz/0cLEBHHHvLjQQl++719ifXGeq/CDke76rMvVj6fduE73K
uyLVo4XJIwzSn1b4GqtOEe+qVvGDp0pGtoVBSEXKhJd3/pfTRDQZMTrg5VgxeoZk
H0nGZ2nvMbd0OudDLucB5RRFNhsqHHPNI6+r0WKce3bt5i8Di8QZdA2ICFD3wSy0
qQOPPrKIHel5xxLYgX9DlXMJsEPRjg/5szB1t6U5g059S/7ug5xWB+zMFuEawHFY
Uw69QZyX4cR0s6ze9hUqZoYombD30GcwU3IlxSTxU29Ob6qkK3DGxrDLU3Gip68M
2TDN7/QouGzezJE7qStKaTuqa2FZFlKZ4WF5NJA9PKkk4ltE0EOWLmq+2Bq4ATDH
jsA2ISrw074zDFgQUikNbdIKiaxx55zqpRlc2neDZ/7avEDQ7RYZHWUhWMxf55zj
J+0h8OTI/3fUzPvQcAhlqlyhZYyYqaWbhqGtyBMVlL2BoZ6TREosjGUjQ0MQTZCq
QaEf3mLSJCRIOR2cKIVgcCBKZCaK2d7LU7CQAKI+06yVXyUFvOFZo9DRBkVw5EhH
V+rCg8UkqqmGlkI45gKXP5w4QXWnRQ286SxYWBKYPekvXZ1Frn9VeYNlZaj3HGCw
gznNnsBa2hiZaXbUXCTyaxCWcG+6XoebObbjwBJFNjtjDcIAeQD+4EdPFlTq8O4W
ySj2vLtMZh6QMx8cKpBCxkiaLW3n5moJsIql6LnEO/IObBZ5A/fhlMFgumJEN2ub
g9LwITWcwfkgJpV2peSsKhtIkVtQCHKlNEUmrYRvfZ2NVg0FybBWPUxq1v/Jd+9A
tiLLdmrV/n+Q4zCQHYrJaF4BySO/H99BXakivnirSxT3X/5HmLmRSc1nkXZR3+Iu
zfyldF5vjK7uAU0Vk+UyzICnt0ZHrZL6nSTyDToLn9xT2CtBBjbM1ELNxJOAn3az
DHJfp+GBrws3lwdDFlc2fh9wiRyBGZ2QT3yETHDE3eg/WEwALHUotfaPtp8Qsu3Z
e5nuATNSwbDusA+1CE0zQye3QE3LDb6HuAAJcYQUQr2v/BDW8vd7UY648ahOlvQl
ZvQqv3lkUkPuU62pfL53HMdEApxc0E9fpMV1cpSWyb+Aa25PczZVR1RkH0Z/tNHN
gzxx7/91pDqMbrcXX2a1Zu0SaAlEBB++wyVg7smS0M9BusfnW6sMb5qg5lGaAEgu
bGj4jTGkwXxDzr5C3/xZ53kvMJF8Nf/ubLvleBS42Rd3I/Ro2509bwp6lhP026Si
sbqLK4/iBd5ZiWYI57krIffmtMt8utWTD7vYKlWY39SreNLKMBqkivPbLmFeCVCZ
MnPv0kYVOF/RXN/cDAVdXEK+1fq35u1CaQjOdR9yZ24sCQLINKMR2Dr5rooRFL3y
XZ6znataJvk9Q2jINdjXm0CeeetpmHmclHMYZJf2gaCTtf220aEjx0VG1HG0GOym
ATL7urKTthTj0g/v8e9AkVJzuhxgJdr/43Xy5MPjgeL0EkMzani+oB8fBCuSfwT2
eA6K+M7SmDFdr8R5yLiG0xdjv38icSqMRHYlRmj3SKws94+DLYOQyQQMV22c6O7m
sFTrBT0EyrOG1BMR5TW3HqgFmGbxcvt30HttYlL7EhmCcoHdq2EdPmU3Im3oQJ1w
PgIW7I5clukHrPthgDtD94oI2us0s68ybaemZQTClxmFZB+wbBwVlBKMZSRV5xBc
SUdHRQtzOeemXPVVJ/ZWNPRb5KVDv3Rbaw3C4rzIaik1BIR0XT0VAUatwT4o2GPD
YDQhFWy9erAjGgKRrPRo0LYDhhrgHrtAc46CzBcdc1WzyGS0WIeHMZbP8BFjKiaC
dYvkw7y1FPgbXfsq6y288gscnOX7u0Y8R7dq19gH6/3o1PtZf7OGfqY2kOB70rMN
s8kTtllvIu9b0auBbXnOunhm7lrZB64DZKliNmDOOSvdEFAvoCSUz4hdzsAJLKEm
rtmW8wAR3LcBmn7r4UjQHiwv8S2Sca6OZYm/eGNmZ3HwveUcyposTu9kJxHKXShr
Tv3CQEyjGYeCXgPKKODygKtfoZ9I2Pq7+EXuPsoUiHaT4FtockwvRtGtA3GoTKkt
vQdslQKwrWj5SjYN+SYgBfv1MXawn9xtYV0Wd6RZH657/z92pEH1BkCWcGowLHV1
4zevKbHW9dz1omnstF/9WSvJTq3jwe7DRhEE2JM0hedPB8hU4nf1vu+M0UtE15Nn
QPHaw+Kokjn+SDIswazuU0EBQFKeflZ+xyTkznEgBGmfhyO2CJqHnZnuweYxG/gs
oCCZXv/qwi7Pxwj+z4hPRvK4MeBMcs9rbNDL/pA70NDdFXjpJsYNBGDyXsfq4Gq+
2E7vKC28bd4bOnkdI67qMoiDZdN3U1pOcluN7rfIPJb4wmBBJfmQlzc+VCeNXA7U
l8Xu0rSFSZqfVN1G7r1CyQqQMrOK2KrxUl6B4qdpbS5L6d5Bwv9jQiCoGhX1/Eta
F7DSshz87xg7XQr4VtW3ProJmTFEc4gqf4kukqN0tD3hAOaiRpTgUrFR9ZIVYk4f
NjnHCOM+Lltbmzf/GNKhwlnqiLD39GOn7aPpw0RvbMed3qxkbnrUofekIGoM3CTb
Fsnr5auZprpVF0a2BEu/yDNbCI1jWJEqh1tuOmoTE3ezqu3mirJq91ET6IZcjSWn
0PRY5m7PBRdRqZflv+E0DtX3WvEMkot5CfwKni1ktGab7q7JgsuYxbOj7oWjfZzT
/pKpGF+0wrpK+E1qJvR4LxVXRrgTpcYrS2E7ZTUowpHSlGIL3PaeoU+i+jAS4k5Y
aBgURErM//9zavrtdbdjaXJ9MzizHuseiN+p6Au7cM8JEFP0fXi1BaCow1bt4oEu
nH43txwmKE1RGDrJK/9yhOmIKuD4bDXOP5Uw9X8q8Z6uSxkz0QiVG0OGZdqEbJ2T
/VhfwcpPJp7Kj4emdPC/l75Pi5Y/+m4Nide/c+wbIHUSDTgA9XbQtmLvT3Ffw57o
SmKMV5FugLbKl9avaIEJv3P5ishJ3c5HWgyxfI8X5oTCv1vwaWUUOd3s2O0/MYS8
N3djyNngIGgSe0ELWr/3+HHjWLdj83TSoQt0ZrirI6MW3levuTT9trB5vAr+tOCU
+Cogb/hWbDpeIIjqVZRgaQPYHUHc2j4KyoJB52NnX+SjLgKSsrlG26hUu/9efc9V
eNdFOFtTxenm7HCdN56ckEMJFzWAsEqAW5WXja8oVpIN/ilmM4suP/3KdJDD/sn6
dr4Eq8D/s2a7OlMd1NTUMaftZf4cSfoN7/KoD9qkgQp5sSmRYRnSsiXU+c2ddMHc
EIStqIH7Je4lBPG2h8n1kvR2kPrG5Pv8+mf6hmCgR0ajuFuq+JJKpC6YjNf5lGZT
WaIRi6XaylnbbJaFNqE+8RSRbS9dgWouorX0qlbzOfj+/K9gOn9OKiVpInzSc5Eo
xtfST1QvS6qLrONyhMVi0R0x5VCWuaxXPsvT6rRpOkKVUFyClVAjS93gcyDp/Obj
MSM7T/rjdjrocM6YTX/R0iK1q56ByLLsMdq/zNU1IoykyoS0sMIHQpGNsoqhZHCo
lWh/sbvFRdxzFfbf3mzP5GeQAL1fvZ0YSEmkvgBIhpuC4SVlDl7Ugqcy+0WQOI5P
vscocGCR498hPSwwTqNh7by8r6k72lPQ9gLMWUSK5WFwzY3l9Q+AecmxNuxt4vE+
1Zpsx06lobBAZuTesAYHkdbcv6iYJwNt6lo4xT/u45Srb/xSCBr161fnY+BhI9jr
0YJBURcrRGQ5LWZdUa243AhZyR2n1Njn83mu+1wKFBDp1OS5K/a5GJx1wULR/bWZ
R1U741sQK7EESplCUf5DxpNGb6lOHbrb5S52RGnMr0k/cO6qTKDjTm8bKFF8reO/
x3DUtP0vh6LJ5N5MDzjA957qQwqEQGShMexkh48PyNyInAxgA4EXv64BhlX33UjK
emh9+UT54AqUZAe6Ghfi9uYnVgLesQRfCLlfAPl98SgymcH8nGplU9Z0JiO5oKbN
FJEdVGrfeOlupYw30BvXcrnwQx0Bmgfd6jT1psGCMPEQBdZhQiwr2IXBC6U2Azdk
p2+QLTTmhx2Brs9f13jWHfUHmkGi2ulnpg7HET5Eo5B/z7ctPng4oqWBm/A6dJaU
eq/5Zsd1xbGHZeA8q/ohc6+3tIcmUKMAuRJ+9BT0KY9pLBAI4IlVu2uPFTrswAMU
kfroFdyNOGjQu2T6zqejXcJBiz8MdA4KMXl4D5fHjxMwMO/M8CAauCNMIO89kVgu
zlhE2iGj4Pbz0rcrrNA7ileiPXJtKbSGzoVncuWIOeXg0cvBtT5LLzC7slhmgxRs
nLQkrI5ZU3t3CQegIFD2ACTmbzNtMFFfb5PLQHskf6AyRziPl8Cg41vrmqDhX1/w
GxO1ldQGn+mPm218qkmr22OltDzeah9b3qvU92IBcT30urK5+l3sU7+ARdcV9vCa
7qC89H/jtVsE7KjMvdGphXmarrF1AQ/sYO3RW7c2+pBZGaQZquy8Uvv5Lo6Gz8kD
oYWHPVUfqZE9bEXta52Wp7TY61KjWvbcXQoc2jzSf4TzFLdUmXfO21ZyZjAX3BeO
h20KhgCoASbgs9YXPoV6Kh6+ckFR3wMp79vkkgBdeLfRFT/hmHuzhELfXi29QyB1
pLeumw5389mkL3BRaJFnQ2664++y6gbwWu7lOYeU63RO1jUVvJ82BLZeduJK9fh3
vzTFr4wFfxXp76XvHbM88kyXjt0Zk58Q3EW8ZhwtCr40WPKkaij+Jfoh22e4sK66
XB4Xic63YhNGAMTD5JkCgBkVMg1bgSKH6ivMrUdu0rWz73xU6KtPgIgcNl05qGfa
4xjXX5B33f6sFuz3Nms55rSADYvYX4fHLRGMNu0nkeCW7bEoJVvO1kKtcsekltcC
uOIMJ6eh4llkMgzurOaD5wLiIbT0ZKt0cIMMBcN+TczHpNihJF9s/GKNZtWEkj7L
URMRg53n+wjneSz1fVh+dqGnq+uLReIaJOGoCxHctysZOUbX0Z1P1UEFYVivwBTQ
t0x7bLiDQi9llkDDZst+r6ZoDX1ykBtW142JWRiIjHFMmxMKLHsPD91W+13Jf0S5
0iYn7KJwZNNBY7FKgn5x/3CUj/yuN7FGTXyJfiavE1/VjjdrKiyzKQXYzQiIYlSj
WXbl5HSNfOWzP0SfL7mWhNnd+1sQHf9f4FYwI4kg2OtWfi+1H6+u5ldE683MSQHn
2s24OX5wDIveOkaHVFpUcLdYgp1jjMJ1qcLjeVNy5hwQtFtogsmEaZme6OOXmkX6
ni6cHCPH4F7rDn2o9yw4dlW2rXi/Kpr0WDoojNPF8fajXNa02qj1TvCB2sEn3Zak
ldY45QT9GVg87oumOBTVohHNlXjOrdqaM3uzZ8tjDWHRpwfi5f8gifxVrPmNnt4s
bmwHJptOqIz32Gf1eHWmALGOIs89GCdBIZdDFLitaB7MvZdRX/ozq3s21pgi0zQX
AGLbOnnBNS75SzNrswY31Kx2D1fh+1ZB6uZjxO7d+C0A4c0JLKoX6o3xd53gCYKE
NFldHoNZ5GJzIxHUVc1C2hlBElzSKF/hv4fe7LMjLmTfLv9fQY7zWCPMdBF6ErwD
NRxnxcj1UfaOimHaWu+YKu52tpV/gBOdPKJgAwU/alMLEsrGfQ2YDBsYgE65NHLK
jgnpnSz7+sqHGBJum9e4e/lCIqUrIl29hSJtpiKPTYxj4DDkK7Rnpprt8s26GBml
UoIWVLGJWPWMlWiWzhsxcVI/VIUoQpBS4dAv0kDxerzD3bxdagrHbg00UQbzwSYz
SBkdAK8W75Tl5R8Wr67p6lszqVe9gT82ChB/EZvKfYU2PZsUW83kEfVmnx22Xj3m
BJNNNT3DjSkBkaM8GJxx7fK8v1Xfhv1yEmF/QDHbjjvqJmJg9RuDgIDxP+24w264
44SSTdpeEIf/C7hz8u+/QjgF6+gt2TfMf4j1gIZqxZszQ5OeELB8CRGjzVcsSs/l
3QOVDXj+jDLCGDuvw3KTOzlRQbuLh2xDoxTB2I2eS2YpKnpIjaDnXrrYC8OBHB5W
WzxbPiCRH8tHf9cV3n2IO3/g+ygVhPsJAUHUc1H5V2HFmmTVMYUXOwoxAbNaHfyo
KTWxgg/tqNR+G25b+kkThYxYMf2HHPHlS/DJosSvA+GneqprmEtFsJuH0SkvihKb
RxGZuP8FT2XQD6D9PUyYoW/8koDkxgEsrMGtBht79W64u5RdY/MygkxDlfnSuaQG
FPbZfMxweIYeRoSvPWhR/+ogXizYNUHXdD6J3eOOuCJUjja6AF4wy/5BUm8bXuV+
tZQ+nII8XTn8mOZIOPM7RZLuyAUTDpHfMlVQhN8+n302XKnEIj2rs8NuhFsaQnv6
iNtTNUIInrvrZ14RU87yWoSh7oGUx7VzgBc24Y5EnLFB8QuUOeUQio2GIKaswGAe
HCagdofqvK/SSyXCnTa7h2FeLgh2J9w6aRNyV/l7kdoDGzM+1qCiwdkpCSSqwQ0L
OFU77ghDEFpZTVPe/TRZXa3Edm2vksH/+E36kvbRnPl7tvdagQAS0V+jFZAyemuV
giAb90IKvao7VmKTgI9hMeDAK3uSJL9FFGFXMP8r1OiPfCIWAU+2MjYAzVxSpeeD
7fhK/pCpf+3dF5qNFP6gM0m7RQllSqhu48F3MYAFrSLQLGWc+9t1BuMxHrWLY9au
gyRfgcmuIMpZhphT+8I8k6+ulCSpauhPHFe3WHmtTbe3y5NlLCijdpbUWQgx1bp/
91mpcD+ho9qGT8N9NdhaI/BPtojbohXIzjpC1gasUsMkQONQrhNPA7U61IVSo9kZ
obEG0VZcxd0vVflY+9H0e57IQZh8Tkik9dldKnp94s0PQkRbSyCNCurprNHwEi/8
xxPdRdIY1ZhXCs3I3C+XMwtoJnYVm30fIVH+HkD2UQL28ztrP2oyEUBd7WDNs+tg
j7j2B2mRZZenHEvWjF4xG9odBc+YegNHg1IGQUglr/+Mhe+BaUjLVEPmNVaIBl0g
rdjJkzH5GK1dr2JbiIzxODpadxccCK4QZrOKBOuOtWkcAye0iFo4wy19fxL6sgjy
WAXulwXAXKj51FMlAfdzvFztghtrALGr2afFuYPpMD3Qwj49P2A7G+EV5hFKHuFe
6b2apLH16yq/jLbmHAEN9LMrMTwzQF+v7heAVMLoVUaVL5xsOd/J3zZNDEb/lW1l
xuxA7f45MnglQIDG7UEsR19mGaRU3A9bHMv0a/gPplXkVA//o1M52TPN9UWlHc3R
vyBr2Iekf0ERxecfwWuTre2qaBOPeIZlpqh1ASxsEcfqf8FpHzQtrSkKs3toquzA
9EJ6DrZuqzJ0IxJJM2UPrxq5LgVjN933YTz3skuYiuxsJk1UAIqLupH49Dh7e3uH
OTK0eEsGoe/I1PMR5C4uxtgyxangjVQjhTv201Kuy22ECgjAQttKwioNjrPvTF5s
loS+nvBcif9Adtnfdu29AyOPxcoPG0MH6Vu9tBHINC5KoqaKd7lxUhLTAlm7wrMC
vc3mWhii7LLQWTLuQeQVyukhAcxsoR7ix0H2gk85z7lkMetSNmNkB0MqlLIk/hZq
yB6Nw1TaqydZT6LNSoYGuma4kCkuM+b+ji+pi+h3AeVpSuAV1t2oe6PbXHRtAcGk
GF/0uMnXIFkt3w8DOW/xcpLrjjlsLMFRG3/bEkHFbcY0deaAwN51mdwnTBnTTpWh
8V85U5aXZ5rYvzWVm53hbe4QmXVwKlf5WXlc0PQlJew79nJ+8bs5jgktjosNh30C
2N96CAeAcQ6HVilx+JzEk0ing+FL714F9TDQrFLTX4Gxw8XOph3lf1/pT7Ge5aQ/
0zq0bsAmyZjJqcg9ni9eCBC6vdWgMtKV42u2/LrtVNJFCgA1qK2RMLgwEH4ZJ+KX
pc+ZC8LxNGREzHVzEGvsy3g/1nnKTcwe0hVVi6ODe8rYN3dV4kiiKdfKhfrdu10S
b+cdWd1e2zEsnc12q2WTm4DOz1rubjWWCmghEYI3AcW7CvuB8GhpRPODU22YbxYe
IU7kkF1XwQpL8Qa+aGioiX3QYve0fiPfOdh2AjwXTs5WSqVW1W4HreAQtGK6+Y4m
7cV3MTnAcPRxGjpsLuOCE86GWZojq23CxYSH0b37DVlIqqy2jT4KW7JKBDlEsRV7
ngItfT5NPnjx1m0ePYgF19I0xwAjUZA1z2x8KTLsroOeN3tn32bLxtk/zYaPT3Rf
PdannWaZbJWm3Ry02ehSc8ZTrqbax7ObcgFtKZmjUSy0+wx4w0igAnQ7aojH3+2o
6LQaMtLQ5KXuMlIK/PLMY84eTpp0WwQAB1O3GnOTI0WhCrqWKZDlOtUvmUTEsMfy
oj7qumSxlcZqb1fU9RcBnx1VMJkgwFCeQuXuLqEQ3zMVuNpn9ikPAixUizCcXSt5
P1m3D6AdlbWYzWaNZBHLBzvS4cC95PZ12rQbroUx12bFnzgwqeEDOYFbjegTm2yW
ADnDURjqv3TroYKuEWTe6OMCYGrRqiHVrdv7igyl2XH9YINist8x75lJ1o76Qm4W
YsP6F4VlY8dukif4lhIHfWGQNXIPN8Tzl1RKATsNH4g4hOxnNnx+NN6dYGCGKBH+
pGRCXx2mSqOpbVZd2uoNU9ofncqBOVakQfpb0ic1hU+6aONPMrJgutUXBJfNXj6v
BMyJe1qi5FlyINIDvTt0k2YDhnTELRjPct9sL02hyyBGlBybFAICNABcw5hCk9dC
6ynMa3wdu6frme6/dZMwcbr+vmlrxtawSjnemB9envB6TTUuK+57EMQO4wYj6+9J
q5LXQZLFUk/q5eHVbv6WZCJkk5HVLO5utp3X0/Nqhysnd8oNuxnyPurhidBKnLnq
w3sOhKfdMU6m6bxLpDPpJch+YM9+flpIM0UhACmBG5yFn+xmdT5qX+0jNPvZD5G0
Q6dDxfrYBC0eNC5TQ/ByY7vdB4z3YhUaBDFnvEDrkH15ObubSr0HTlCvkknyCgks
MUC0Zk7gsyvrO5jdTTSc34st7cxd//eK1p9nFsi7NgoQ4SV5em8DlJ+EBS0PPj7V
VY1Rju/3DUdgE2eirouRegx6VCQvmrFoBLOT+3UFF7rJn05T7s2Gt04qgv6uDLz1
FezhU6ubFkR0kMQKLyEz54ZO2l82WrJKxmiETNTRKrCNTLQIdWRxqCme3ejE0bpo
YsqTtZEfozeVptsCmkwYXHGvsbjhs5mWp0KHTmqJIp2dYu3tAcsvzZ4vyB5xudY+
DPgGGMut8jGSl9d8i2vmkDdbPqDpuk5tF3yUH4R6T2XMUrJt+eO7qln3zhaKih0c
4j9Xe/1hN3kSJPFaClawXpSzh/V5ngLLYl8mGlCjvTMcZdC3J2bkVTl2Y7+V+D5v
nbZUlgE4dQxoV7jLr6Uc0ipU8Eeh/Wv9/W6bcLLZLbTIIAwRAldFMsViRmQdfV78
4M1BbnGIA8LaULw/sDgVyeHvJRLKFfsHOuZIyMnsOFC2U1obm0QIKwZ3UlVFQREu
/q6iRCTzrkqidS3sfwws67h7pEmxw2Ce49qUHtiZ7QTCh3vhtpCzIARbqgBRXrDg
nn5wk1ta2ACSoe0JG1kdPIEM6PmeTusCJFhhylRyhCkdy94eMy/1FKzG/awGEkcA
j7tk1X4Khrz4XdETdSpOv0upNgyQF+99jMpHGpDtlBPqKjNQepDt0aM0UDIpOtDM
+Aq7nO2ks6uJapm1iydxxGLwRrG4KAKJ4qKkTXllv7IMr0Auh1i8EYPSoJof4A5h
Hu5mexjXPg2g+LWqLSyg9GS9KaDkoAWZ4chFsMudsoFpoXCmCqrRaL1fQyQrdMDg
qqVrlFoS9MScJM63WL1tRgyZRET+bV4KAuI2l3PvztwiG0ePrqnl9A7u0XH04aYj
ylmYhuFmxrPt/JmgZD3bBioAa6560x5veUhjUjDRci4oXfTwCoOyGvoictzA5AKU
tkT3kqeaVkreoTvA1drZuvG3Ha33lrM//p2GRHJROd0ns39A38PhvgtyLK9X/MmR
ibmGkG6ntC0ywSkcXT2hmC0c767/NxJV+cuNNfBfzLGpuKJAL3KWu6MklJwWL4IC
Lxq3cqUHW4fuMAJoPWJJDC1UV5+Wrg4puMSFKQBQ0xzgJn4qolawSgfxnoZnJVVI
corqvDxnbbhHCaVC9iH0jkIRNYyHpLrq8WJw8XsIGXx/XDFc+X1m6GpyVdpJ/Zjk
/W1s/0fATGlzAwAdXqYRNGCAC56zKVf1A942G0pS5b4ZXoUK+Xr4CHfBQZEcm7u8
rO+Pfhyizla1r7FFUSFsDg4i8cEITWQqqLz2FMBWZgLycdaqz9XEDwBJ8UsNk0yW
y3SJ1Ogfl6gX0ajIkSK49hjBCW5WrJ6jGSG8q3XY/0Suq0FksFwaensbMqOpdnK2
jutQW3VXjXZxYMQavGUz0l6CXm0QHqFRzsJLfqkJntiBd7lK/Z7yE2nrImwWl6WX
zo+nqIA3KCOcjfVggJT5lWJmShunfGv/QtI9kgTPByZvFZ8jpYDnRAzVfoMsQp+K
hWQljksK2vYMIxrjFRcT/xX+5DYxrtiOXsNhZ11/E0Np10UzqoFKXo7LtCqz4YV5
Zv297nprftMOoheTitWbedOMKwU4VWm3eNC2hkT0YECi3c5XbR9g8D2crAxYvrxO
E1vep/yHGyqrdMoO6w4adQ8iDWKvPetyP4bdRokqGyC9IhaZiCcLtcjJmDPW9mOU
SCSAfLiTV8eYeGKBunodvKfoOUhRwmPYMekWbBCkWS9ySdrG9nq1qCwGtRdEoNKB
5xeuy+J4/bRK74DSmh/fCHc02mrFk5bn2dM5qv17UA2Rkc1WOMi7LBcjd1sReAGP
KaJsY0q5ZOa+uZGvnbn6nnsqyDyjDAgPkrJeT3djlFzkBxicOGM50Kpvvc9rWMy8
UTR14c1yiV95idBzswFgUatE71kZb5LmG1OQQHbLsqio5ZG6sCqq9Ik3qxIM6iNU
U1ktBT46YmGFEOphuL8S+jZhYedHcNy69G6B64pNhyDU4O2pUxdoqqn2Em79yk7s
iuY1BevcAdSxb9usRTFzXcBVp2XpiSgXfKJGtW23eDXM32WvN6KPqqZzQ1BmLq2B
l4bDX83Wjle487wLiocije7KKSoXqbJCT1WHbzbqqEp0C+L9SHkhitOG9I+E2F4Y
8P8ERQdzUEHpXcoG6CenlRBG0heGseS4jYhWyeJ3gJ0GdvsTcMYGS7BxAKLd7s6h
SHujECe86sHll9oGfrBq3dGG4OGZ/gjCFC/PKbE0sjFXkjdKrrdJcNf8XxY+A4io
SSSZO8LASD8NHg54GIWDYxdfTJTcsTjadXQYE3/v7ATd8M5mSD5+dZggFGkAO98w
t0fV4igSd9C0FkZaWPufGRI4t3gHOUoGvzx5GBAS4+KVhLSejlqwBs4Iyn9mD0UA
6ZlZase6KN9U8MyMt4f3HfK7ZhA4eT6wN2TFzy8HwL55bHMAKgS8UgRP1IixMoux
Q0sQjwvtmKWrxzuch/kYbxftDVsSN+5+C0QDB67+FnAvfKbLELCURLUYoPQiYkA8
UJYXddauzeiiDfSMlmDx1wQV/K/0sW0NarmbQarZxJlhxVLwHcBAnOSAUoGiUQbr
kM7/7xiLVR7t8UKueRNMZqPO/2zSFuq3tsIV4+QzC0z4UaxJfEGIeaqf39PcGkG5
obzCPFNAzYz7h3oN9Dsjrg55qC5LzUsf3WpSmde0NpBdxjMdEA76zeULmfhi8zfX
1xuyXD4sldX2Jwm8AQw6AAv30JWAutsQZzUfC/uJ9U830q50bObjOT4w5ZWDCzSt
gRxBlyUeuOeyZ0wOW5OpMOvvHuQ9k3M1WujkuP6eJvPFZ03tnM7iA1LVwSBtDEV4
ifE2EeZnk4iLmvyRUZWirRcitxK/tQH4PYomiTxbbHmQU1aDAijEEHvpO7ZQLZ53
m2aJRLZtPvmYOts3kAkEBFvmmTNXOefr4TC0DetKyGcX0fD2V066sNzGP2Gz17sB
h+RTAh2uLmA0pLLzC2DJnxKI5r3I3Blp4jCjOuSJbHPNEYQQi//+tmvEvXgz14gk
6IEQy039XaetKEyo2p/zOCV27RGFV/eKxpomFrywTfe+C2flsdda/zd7QypE3FLH
N+H1ZYPaX4PgUN9WE36jwXESuv6WFrc2nnUl2yRSBHniFVQ5B3EG0Z/113UFSD/z
DAlPyOdfXN0fuAj7e/Q5b87W0Ikl0xcPysO6u38fgxnIZ169cfypzgmiW2vErrD/
OxP3Ztf8aEdaEt4ekaBS+wNbyjE4r4Dd7ZBOp2nloTKbJWsoSxXMPbqnCERWrfoJ
Dxvl3TM82Y56nVgCsXWyR1oSgyE8BerhOCQETnVDbY4vzWaSw9/SEOnSZ3lymojL
FHh3KhLedFDBGOMVTag4Q4XLf93tVtH2GzqEi+/ZKIqsUnGKJwf3kIydsvzoaIkt
DF5eQHJquhtqXzgVPT1XrK9IAj1fgwR0isUiEVNP6x6dmUYw4rPYLGZPdOQp/tmk
yS4aDFITCQ8NmnUcehLodyQGckqj8Q2b9Dm85aowbGTSODLKa28DpSRNLOi/3C9F
9vaLRyfG3dbhnLbH/Fttyt3ulb/pAxs6rxNxkuPkM91ATD0naf2mWbrxAGZichg3
J4NjbtHMEjgBBz7QwrrDoEaRD2moMWuC9iXdUob71QTUO3TukfdtsJkd8FExv54H
UMh2gCExkOQXjGuzf54bo3xZ8RKVejkJZdcnz1mYboLOdHJcEZopvfhEdgXxTNb5
oRjtwKrT1JGOwHrVIDpe+eVxIkAtBRAYXVwW1ahJnDE5DzJT/bmXlHi7BpZYzTKK
YCkUKC70zyKgZbecXvoQGNJt8X7j88vGXHE3ewXYGK5I+F4GUxi4tEBrwZUivL88
ak3xR7cOSHrMD2wocOqJfIDJTZyozpN+cfvEt6rC3WknM9DLnsbOzWRCF5Paze3N
o/rdbShpEpvkGkCNWnGZH6EBHyBIswM2F6MRpNTssOPp7ltcxoIHraA6JpPQY/fQ
p//lDVaAEce0N3rbLCZt8OpQG0HH8mpNDY0QMgP7Ms8KKTAgBxm/kIfjUql8q0S/
n/z6RdYb2Ocm8fsWLxpm7iUIV7Cz6ohSw+tlHgb6HvKriSZqODCuJ2NylU5JCgMM
Tpq4rkYLs69m8iDU5XMbVBZZX92NY8X5q8aKJJ8sl0SEJ3mL2F/U3c1TPSPfxSMW
aZrME4A0jEfgtXGL/nPppnXUWtiaISXq4i6V0U87i9i7g8EgMeSXZQFPkl4TMe7C
K8JInSPWIjfE2TvLWk5yLJrw8Lo2E5/SOdVtmMnWMvKZvBZ7uZ6N07p/vk+jg2EX
EWeHjIAXgyrZHWYG8kIYaPdSpQ8dLn4gPHtkf4qH3YG1Gcxu6HXNjvIV96ppAI0D
RL//zz1iv1LClNaDwJ29JMtmqMLnGR4+xHFE+5+eFGUWdusyIrgZ5cy97AxW0o3g
f/fcFmuInH8Ts9enqKYBB8l+gRpfwZAepar7qa5AhTcjw+00V1xRXoTGPN47ZY1o
hVmRHEWb+zCz0BUfP+7IZ8nTDz08aypKdEMekfBPo1K7EJQgeY4vEI4H0qlrtnyU
0GPfCPXl3N2ErmqZWBh+5HEd53+Kq9wsLG5fNIKl9S/qzj15CgJw/QxH1rqrdFv7
t3PREw07wYsvWz3nTgKFlnL3arJ4NqE4h7M9B7ikuR7h5zkXr+EP7YbTuNa4f1rU
poPnIw8KAaIokzuAJD6IObtKyaPxNCL8cSAedtloCN34UXzTB+3hWmH7zO7DYj2r
cU4U7Q2rQc2Z9BlTywyuPibl9dZb1Ao37lwUq+p41CQ8vwgO3PG4shZpvrf0lBdz
kF+fs8lBghb9YfVB3MBl9MFtGvCvXiDIelTF4xKlCkE2rHoflnlYUp94ZZ2Ki5iE
paYHWWdsnoOtQxSLtA5e3514ei4dVUl5UY9NNJYDZ9qK5+XNm9gY9mX/Iodf9C7q
4IgMoP0eyCcxs3cmdtKaUw4a28iHHbF+Yw/lCXp5zpCx+oywA777Vnwx8SEZcrxK
pPxCm+yTj3gGtUhbHOSKmsrIZAztg9bApAnrs05vLdfg1gBAx9RMwH0Ac588vGtT
GJYXlFMeuRO32WZA9+Lb+UWLEzFKhBZalxNDDEOPzns2tqftWQavZIhpIMOfH77H
RIUyC0uZEAWj7SgFtm7UrU/uyE5F64lBOSmQmJBdaYRMxgR8peX1f8FZwBuyesSl
59BIm5tgOnMZqMIzHolD8Seas4hF3sLbt0Ca0mdYKktteQif+OanUMaXL4xcpoFp
aAAkqZLREF6y0gOyJmmEAXlbSVZrQEBppRhJO1kYpry/Bi5AKYBOOzHzMQmf4MCH
KudppUlV+rK5oclnH8BsJnN1Y/lD63GBfB+Aiwgxq2U3UJ6XB33+9qr5YZTn7Lm1
IK1OeEVpTlQVj6t/Oei1HUfqZhYPBNqXOSyBj6ZIuiZ+UekYjp7QLlXcJSUomZ1d
0FqbrhsKaJQmsKjlYsE+wqujANBotqOYXWnWis7xO2+UKTmlsvaZsldzVeP5kHc1
Rd6IhrCpFqjXdooTPsHAEAVJZKm7RhyrdZh+xHd4d8YtcWnJXSDKgntKoZ1ZqEn+
B+YgveMtgXXDgA5i78+8eW7mrYhBhR44kq6ao1GoKntDWQOYGplIh2jzLnOivKXn
1XZelKCZSBfmLq4pJGUChWSSmYUL+RdOtzhEl2vNPqEqLHjjBpQtq9vEzIIkwAWG
IebzsnTniRcad98X7Y0YCX8cmtHySt1+eqDIvLo4Uq8DEPTtoDXNzAiHQEhbL6J8
nVjM6uSyqn+zd/n3ct3HVXtqbrtrcukfSZTMh4b3WF6nhJe5OdleazDMguk2/41h
khc1vXZEU/9tiFYwyBp0WEF6WdrGBXb70vnV1h6ticj7hVPb9hCs/xYj3i1Gk0JC
8vEUn6wAiA+MmwerQhaC0Fb6ya+FX9BVsHfKLnzWM0LJ14gfTGYNDTIB7o8IKmVv
QpWsKU3ftQjl8VVZd6g3SRN1GNn/SjYxWrCeBCV5f8PdDthaOfS5CgAZR+Pv1zvY
H99qfQEVAzk9CzHsKenE5xcu6SagpInrY3GwgOp+zRXbBX/iXhx2/Bg7Q3wYcrgM
NNR2uLPwvFuLUlaUmHElTpFtFaEwO+9d649kMS4rug96F7dSf6cNOxzgOReL8ewA
0FvSQtyPlvgo5KncYXTIGFMtMv11iNGoHWrHoFrsas1M6Cqi/V3A+yj+fhafy59M
webKz6zf4uVxrKwZ/FcQKskkGHd+JsAUJJouKEuVgOo/zjnemGK7pb5gRlp07nGg
LLdLpBQ6V3775MjO615v9e4KreXOa6EhdbJihwgTrO3mucBgMf89So8OIzmNsdp2
OsUJdsC3qarJtVxf8wWBzwVXV/uIXr8dUqL4TyKSsqrXieuyKVRy561XXzf9DpD9
jVoKGLJH+47TSeQrw72VxJCNgfIcHPGXwWPT2GjwYz25tUPVdwHTAXJTK8F/tNpQ
GjItABBLeNX1Q2v68O25CAqTriPLbpr0S//wXdq2Na4uZuQgbWtTqp5IG38Owl+R
dySXzRrsW9RTLaqyvI0xl5wPBQx41nDchDzPZpu/ojwWqIgGEzv6YL2+CTFImMHJ
VsXydqieCPMpyTeERRP3TRNZOk5yqPeWn3iPwt9eTYZsQQdSYfaJtIzm207oXNMh
hIK+dYLiW5SHAJcqg2UTWSmoBAfBqx9ruKqjkqRa/Ic0xqZTzChOOcNUMveNHEJ4
nOxhSVO1vff6h+v960lbBKNUTKg3RWdOd+L2tRaWTtdX2zAQg+OqRWfia3RJVmRo
s6eQvZtI2KdMT74uTK3I4dxQyPcPMLjQZd+zXqRq8yj8CY40+UXt5P4BpxNBHm0x
1vQW2vhgE2eJL+5ygzUpoZUHmNGUE6upzyuLJhtGqyadvU9zKY+VmL7gV7ENi//V
LVdW0sHsJHAuWI9mhSa1I65U5o1X4DkTj2XZWEh7FWigthCpFnIOfmIrlTyLtmPY
jjwGD9x07dqz9B1u/ETd2SXJsDDqTs5FRITdwj0qCm9CHgDa2z64Zm4z01qTYOtb
i4t4FabSz8NKJyTOHew3UJsbdpyptMnyD251yFy97I+Y5jvvRjrQwQMzmzl/6Btu
1zzWHO/oZLR1plv05+NHJNrQpKRKmF8PECsoJ+Gp8ntYz8xvtMZd4L0KCJ3v7Ka3
cAYgdcMFsWnnqYnvuV3gBCgIKyhJY9BbBqs4LVb+kx4KKdTOtnWS2wT8oJbJ+ldh
VmdAMiWh1m6xBDlNI8O84XZ3xZb10nuyBdQzpOXn2g4NElAJP6uO0AL3dqC0KFKP
mkr9Gj86+lhk4Z6LA4PQxLUMyMEcp2Pqe1mgiai8qx6w6fi10pMHuHgf8h5CmdaF
gOfp7AibeCbS7O9XwABu3sjh9ZVlewfpGARsebQHl6guvgEzg/dRgU79wvNtflLq
H02xtM1dWpLi8XGBphFRoWJ/7fKgjVIHODWuG6D5xSso7orYS76YOUyVlEvPuaq/
hlVVfnRZuCY83APuuAvWHqhA8hqDV+477iDBm4vYz95xls7U17G3SXuvn+0Ulb9c
I0sV++AvBk/izXomgZeq9Ott0TIlicPMZ6so/tiZEClbORbBa+18LSQORaEEVn4E
XZiiZGrxYnYFnGgXCCxZPPR3wXS/u6JIxraoJqq792fKARN9yzlS/Rt2hHhsIPyf
32FaC4IR/lzsNAQ6+yqDFbp/Ojpvz6o0yuEU6TTZE1E+n1cGuqVKcvk2bSn6RQyc
/vtd8obdEo1Y1dWBpr+TZTa+BkKIee9MNE4SZpi+BahxbawVcz7W9zHJX72dq/G8
IpNl+n/kerZgkX7Wag6bSV3H/0mlDr/Ccntp9C7PAb12kebPbHRjwRvgJdgXzFV3
dzYuT6LeXnuoa43mf66OjiFbNHWp0MJf2dsCiZUj79NIEbnijtUZq47Th7aagtvm
oT+YFC16RdWz/2dd+k6SgOoDUYOBlUcE4TwyPdbg4QSkDY77crrARfe4bW8PJQwZ
vLOxoDgHNs7LQITZL5vNJCsjrp5drQ+4sKBlv00/cGF67p6rqKhRruSTxUP7NyRj
+kBv/U4HZAlXCMGMX8yYlWwZg4L3+dCCUqsY6+NxxzjFkeU+Aiaa9UN6Q5IuH+fw
DHMrbC52WC9ei2wp9KFcmL2+Jpvgq+hXjRlI/RiuZR/b0nGrv0K6i1TcKi0B/0dL
u0TZ9kkVnwS7vHBuqT5QJbCY0uNOBabiTfW6o1CdgylkIFEjYxky9Hcrq3i4Yyvu
JU8ckpd9Qiy3PZ04VdSegMZlpIigOgDeCLBGPbCwxipZJBuektOVq24FX8xYgWT/
4akK9SNNdn8u6eBeltGHS0KVnxR3sU71TNepI7uFqbkbDkYa7MWg9ao9BMpbZAPJ
exWJTolGJgsMxz+8iwGzVLE3sC5H7c5b3n1w75uBBrTMKpi2BYw+V6Yx8HJ1OliX
pxvNVsecfe0H2wRoXwAQ4xD6XocZiii1tGilezv57lJn24O3QCQW3f1T3C+uhX0v
C2i6A9jNE6vW7rXYB9yXUMfhXYlsqhX3UCCjEz8ncXGQXdvnRb5Y4W8sL4hJWs2Z
aiSimOQS3DKYCb0K2ItTV8lpah/wuR80n9gk58+k/kdVTZJZGowHNQ9t8ZvtPe1r
bt0lNsz06cH12WMNP1E69j1u3DJkxIPtEjVaOCqc5yNJs4XyJ/X/TJlCH1y1JqZu
4d1mlDahhhfel5eCOCPkPPUk7t0U+n4D0lVzG9vLqxXmbFyDDqNJy4t8TZurzuOB
CYVJVtFklvYakWnAmMY+Yp6fy8xpeiscpHLyome6NJzgFJ76vH06fnwsEfwAFCWv
YrQ/usahDCLhgFmmaB3EmXSFPJmqEZUCM3I8usyOLUtLGcy2KK4iWiTJ68GYL2OT
S950J1J4dRg9uyx5VXVD6D7+qRgxdOEVFenrgDeJHN1g2pfZ+uY9qwEvYReFmHll
Gmdj7SHqHiP/5yoNKg+HFSM2ELCcAEhfKdCcnDqe8FLoU1xG+KA0DcQetZBfLjmq
9x/xQNSvnWZ4nj9tJuMHrDnLDDB0rUDU/ihzBq5/FSl/NmAcXNqMztB2Kz99k/f/
RnZBpgflq5xB+jMtMUfKtouJ2SisFIcNFP9WRexDjb2t9NicCO8PL/eiJ+SEFsXS
AFOhKgKokqeB/NsPJYHPV/SGpa+jWBb7YnewhJBXRSQx5ddX7efFiR6gDxp324dU
Ywr3HH6gIrKREJOGZqm6HPWTUw3yMI1x19RWiYihLEIPBnCeXRP91S8431sI99HR
xitsLOWhuy+C8X3r4xGCIX1yPbo5xhQPtomMhjC92SyPj+g2nNCA8aeSn+RZEQ5V
cQhzCO/5dyVn4G3C1fH6GgtX6Q6zw2TadfOabH7rTsG5dsPbr1ONJFhE4wUE9QmC
RJHo1hVWEw2al9u4NzLJvdDx5HKGJ2LdI+DBHcXYFHqCyefndRBQRtKWI+2DU0qg
M53BGIonKCVOwJ2V4iR4/ZwKf3Jw2EzfH7s3cyVrnHdbLVNvqhwJSzzWp9s02qkg
G3uEQuORSTSe56VtC8IoL5H9TFjdqTvIEbmDoMFYBH1uE/wEGRMMlffRyLxLivKQ
quDTO3ZE+gU81rwcC+NcgR/41Tn8wS0Uk41OLtIUDStmZjvf3JPBGudODbQRBr2N
fzHgnZU66g5lNKnc4jYNl1XdvCSYCwI0IbkeRMG2bKIYSgSuTsEIMi+8McfpcwtE
lIkURFE8weMKaNtFjzk5XxRZRd4fdn5pCVuP+lEWQ1/uM2VdUgAVhSDYbln/xNgA
TmNuprGZJKs8bteBoaHI/LvxwlOBs2x0gmkETpAFlR+WB0rkiY5X+oXCGummXse0
QdcQbV9czQ2458k5pypnaUmrW6R9rIOhdIbAe51a4C9vng3q+8MdrN05GX3Fl2k1
0hz8RrAsihL3G3GAorZH1+cZ4SilABsnSu2kZwTlpa50M4eRb9SVEFm9xdJArXtc
ArhbBOyXY3NFVV/56p8BPjzXeiYMNKqYCqA/gv9Te7+A+nMPaipxuCYaGDtIDDTe
8CS/KMWQ8SisrCo8TP4fZoHKkhbf51y1xZkKJzGBGWlaEcBUo7sX9XIO+nhWfoUx
74SUegQfKLibHZeHcbA2+DI0k+cFaKpyCx1Uiu/H+Rmr3fcDZ/HEVTafFzudhKvJ
spSfthqBnxzlLOBKjS2eS7m23AfV8ZSgYKmmCrQPJS2mg2TeJPTSU5M5TvBkPgDE
Ivu7aGfAqPUzNMjAiBnutI/SkP7Q+sw3if2zTUGUhxEpvUfDL9Yclwg4AFyaPlbw
FvInxrxWsoz33lnhh2tRYW5+ZZP5haYbWr7LZHF8Dj1umYIdpwRta0k7qiZqibE5
cvl8ERLm3f5txE32oHya0RPd3mpOwf3gdjH02CmvcG7elfaAtHJlf7YxpxkymqKT
rgr07N7D1KCTo23qtc00ARxSSPrFU8L3p3dtgsaR9W9zTddbRuv+qprCh7wJKwv9
MhvcUuvWTtJZa6j0cGwCJtApBx2ESTyFq7RpAIkS2fIvAoHrkge0YACkIV8dRgjB
YBfJet7oW4sM5ECD1OORMbkmf4zMwcUeC3NiyMAUGWGaP1VuZrWWbXeEtP0oLJwe
ylAy298sQrVX/iL2wFKbDzf0Pm3HKP9iEolgRWdN/3mtM66weKo0w61nUvM/fNm0
3eEi3j3+Adps4Ha8A0fUDToSnuxqALPTnwkNes73BdjGFCqDbEfHbrdKEIMEj8ml
ep7uCGMx5JcN+5Nwk6/oqUFR87o02/WYE2gAgm9nIRA5+NE781ad12m00UIXDS9M
+B0JhMC6z9UQZvgsUP49YL3U/IRgcCYitpQzqhUMLMnzLO7QhWvOgsOJkL+0MPz6
wtbpze3n4xtTb9oADqZNimAX9ON6w50Aw3L/o7OgTcvYN5Ze/oXYzD/Xx+ki8b1Q
Jhi1OTDvmWTaqrFEHd2nPhbVkdC4RMb1EkxBcWI/7Iy9f52BXszlHS+3iLW2fmLd
njEFwpCjW6UYzBd3So5bOhUgD14iTCawzsT92t7ph//WOdeW0hCxyvnsHjI6yeRh
M9gFItYK+xQ17E6KMmomKGyPD8rAIOSsuUDJ22j42tTvmgGxJOvTBGtMXS8Q0DDX
skRuAlkwt+vR/AcFsbraSHiDNad4k4pU8qVCo6QwwwTomkdsV9yaWple0E+CXldE
AmxIQP+hyYeupRwxnmk7PXjT1EdMmAt7y5Nx2+nseuIwcOAxNDeIj+4FaJHp/jBk
0bshOY2R7+8tR56I8M7O/Azx9AGbNVMkdBrVB4MDsHhr515fkiBRCZ4ul6YpQCND
ZkTZ+qutHNr4Q9MpZgGXgeooOl8HV6fFJrZ2qwZt7T9sI1WMgSNTtm4oKUFP3nlJ
eitjLD0EGiATfknx2vfhcdVr73FE+Dj6STAqs7J4vA2yXaKkW09VK0oTlbS7qNI4
kycr2qbTWYHtgrha2UMkB2Ya7Fwaz+Rx39lzxjskWL9Jwtf+yarl1rZBi9nk0MeV
C8Nom09sQlULjc8RRuhIlkONAjItXEu/OB0r54qjr/b/NKzuokupvJcHusQJ5b+P
UpSFp1YbdrFO3iMiWXHma/QZkBSKoreMifwrzfxE1csV+1f6qQ/UpJkBmsOY75Gp
2sx+66eEEhiPCurB101XWnc87pzhOWAsegeJqIDVLIv1NulyxBIwo8eYFejOfaLd
q2/qWhIhaj9GtK8uzMtWVDsf58k/0PbZp6Yi82LKRqNsTq3JPJCMBD+0v+AmAcJu
GM1aX+xNTIqml/Df4aBVTDELfawnD+Fz9pKvffD/cIFIBuPHNP2x2DD1UhsuqpKt
8oa25A9ev2VqCB/0R/2KQ+EhZE7UcCt5MqZWKnw0ijDkM5J/GfUZnmZZh3wk6EuK
Qm2QR1V3iwJOeGGVxVTTcdL++MUdHYfwFDSFL+Yfg1OW96buOECrqhaJgWhej7hu
GVaX3Gz+pqctm8tqYNrafGaEvBlK5fCCrFyN9ooKyEKO0IAPhakBJSXVCshnKrlR
01unI1crRHnP6uanolWGR5qo7iET1tC+pyOnvKYR01gVTvU1Dz9iWLYWX9PucYiC
8+RW/d30Yut0QDApju4CtNIgHMHeqkqZRmGzSDdX9umQf73N+xr52vq+UcFmbcHB
cu9WrMvIQ5hOGQMJ1AAhOOdxuFCBdTinUapv+3q9c5IwimnzAcmBnjbW6mAnKUij
xhYPCTLjyQg9WTPKK7ZW9CUXAikxAGLIHVwBdcCFJ+s7yke4AZuPZcz36T2hLvKF
IohwHpus/iXvzv26GPnTrgIU0rqq37yu8pVlvneUtHKO3r7Er7ZUdxyH2c7jqfpj
z6oQpZc12Tn5xmXXru7eriXlM6E/UT424obvjii/0VRgIlUM3HDGeKSgEYncKB4U
s6eIHFwPKeIAuL+9vV59dvdzuPq5b7lunugn1kseBBv+ES73mgrl9afY9hWp8vp3
bjwfKS7+3pR5TmP/EMEGZ/5jGRJUASOVbr0ZNssqFlaBEU8A8dSZbyf5XH3gv4M8
ii/7KZZ+2M4Zq36WEtS/YKkbtJs8L+WawSD+9Sd3PaQVauVKTTdmUMkyu3nmcInY
eVTOTw/CHdUfkLZPU1+YSSsOF6gnd6Lgo/1QN6UyCnNaLthnCpqGn6TUKH7cxkhH
Dmln2S5CQORgn/H+crtir9lz8MbxsoubUBFhz35NL5rUcPl2fBeugWIT13A623p6
+nEMfwA7vDfbWACAJBbVo06mK1ChZp7xLFgoOKs6jrbCrdX7EF3VMUjklqx6jONp
En/oD8VLRjHK/OtN/WdtCOt36qzdPaTA5ejsKAgsAIgWjbs3Zen0shpEO1UdCC+Z
P4zdwC4hXjR2EkZK2z6c7SLIDf1Mb2qWHHk+VlFjj2DakB6xbgzbcXLso/g5M6CE
TOi4SK1McnbKiGPP+jo7wENdxx4XDYC+bMnOy4r3jIcoeRiA9GkHK+WySJjBf+qP
4N9BKVEy2aHKNW/fBwJxAgy8QHoL+hsrXVrH8BizQjhRR9NZpn3lARHRyB+9P0dL
f6dCISvzIziWQpsDR9/eGC3O3H94q2DidtAy/k365jIAam9J8WCv4Rlad9Np84Mh
YsmUgSVoJcyZfSh79wzKxz78z8IfKsLSHSheeMEZ5KkrV7LGamMpzIvNko0h+qIu
BjDnUV6ShcljlXfJRDBt3sSnSJdXnd7LUXlrO59e2TLny0bQAVbDRk10hFzUd1j7
w9eHWTgSzA9q95mHxFDILPcrxrsMalMBIhjmxGM2RBQPt66cmcQyzbKuo0atlK9t
hfCgbmJ718fodAnWDQI9vuErhVWRJz14LS5NusFPIqkvHwTQhjDkNnQa+FwCtJSK
qbGSYTN21XMeJYSf5Bxxyzo86xsDLf+ZRblfj0Xf3WTstlEeMHZHOTwa/V030pX8
MTNWy+gCJTgGVfAZjkAIn3YOlEH3/cwXn2LV+SLG7BJwQUMnzB+u6Zr1DFQ4j18k
v4Kcp8KZgaAOYcFi6khSiTcY1Q194Kz/KsZw42Lo5Vql+enaHxLV8ts6BZlpZlJ4
RinjiZzlSSpB7cX9I6+iATu/FwbkTAX1c7KozloRL1LbJzJCqULtxqcCQV0T8RV0
jRgfvTaV/5vM+xGLkwrqbr+MRqH/CWbfcolSUX11l70zVNX9C8Sg10deKLcL/zk7
76WDbHzIMezJgRCqECqynPhM/4bR1sCKd421DkxtxYzilFuTMWi7zAUxyfp5v4vH
oRQ+Ee971ZMwBIfEd2cb1gKRNuEoAuUugzazBGLtRuXVi8v6OZuJQihRchGY354J
Yr/Bog2lezzZJ4ttZScYCShm6kPUqYGOeZAn+W0C41PqswT2xzOjDDd9IUl2g2hc
IhXTb3w/fBByVMSwYroKQdRAR/OP/W2snC/AOIHy3NpD6CBJZqueLHdtUqQocpgq
vLMOIDDgNHYfzASba65oyrKKjZXJLO6/XHWlWsWTpKTS9P72khIyr+j//SBwcFP+
y7l8jT4eaxo548U/2CZ3DCC7/FaINzyYOAAsKr4kNpTzOdg+a9Avw1DcvoRafMlL
2+Ai83nYy229cFf0FE8f7Jsup1J0kkUE8o/iVb44MCe47r2EwK77MDy3Ni1JujjF
76tW+VsAd+g+BJ2sjYAijfwIa5D+RPk1SFYR0htiWKuB2r7lLjs31qStNOsSsFHs
tHqZrBkRFqR8TZXodahVxNNIRZhNviBMVKUG7bPCiDo0nbHInq5NLxK0vdcU1eo2
nYc70YWKRtnXRHfCFCCpKgCW6mDOcgRiIevDXMRv8kuKR+NMHxXKKNYVLqkCfaSK
CxFpn66FQL/N0MSgpPLd+ObiTEcVDDROnm4dKrMtRIFrZO7nyyPm9o1pt7tGbWDR
zp7hLuTYi4q0477QTh2WEzlKL/NM31110za1tdH+7y7C7O2tToK/e68a7K5vRFwY
TsRviphN2HZ96gNGRNom3gVOTXfBY9WqpjpnkWOnhpUjvkVf0OffwZik4OVqMxGv
leFdj/JEHj+oilkt7ocdHG5vfnegsfjYqO9sUFMQYrR/vsqvsolsgaYOQRGHH/7j
WQNpErjfW+/x9WC9O5T4MxoTInb1Fw8uPbMbajasPoGD6/nsNEEEh/NMD/zAcMA9
V/iMC3s4luG8ckr+ms6eBmEmNtO/YHqgnb6O/pvW96Kd43w+jOCQXRDAF9Vte4lX
h8huwGNBSj35SBrE4pMdBlPKv5QiLcZ5RTbRBSYYyd0ybuxgt/fTEAVN+s0XAVzp
qgLr6St22G+dbXidipbFvoYrESlcHRmtrNI50OJN6wX2q5IvGy0aTkIyu1T+3hIE
DwH07VRDtGbxsfgxOsuIB+qihRXDgcsc8rGOii0cZvP5v1zLt+sD4IU0VoJMRexj
nuZlu7Ty/SOIVzFA3kYNUEDpwX7VkErKjkCJi+AznVsZJb15xP3XDpFEDHApt3dR
bprmi5TYyKrkO1DM4L4ysrgMdQ/gAsISj24OU3CNmfvGMEGH1myTjOQlaU13lw9o
rEcDbIkk9/2RanlfD7JwtBcK3n0EwjMERDm0MNUvR4X/UW3eojHGn5/V5d4h+sPs
iKbOGm4n6ibTjwMy9C2ozLIBPpbZfuHsO/psA/N9a63iqlOeCTKTKRNHupSKrKQ3
DJk1kEkC9JcsMrn6dUmx0dtNiw6qA4G2IUqtwnBZNk1miuDXeKE3cMdQJx70fdCu
QzuUhpaPu43GHcpXz+Wi2vzGXsN9/Fx7WlAbljaWZd96K5A1WdH/peSdC9vM2PFe
fnJ7I5yZwTpg+EOVIO3Ry2QbKPY9eTw1zd/GEzbpmMMVAaGPdapMWkqLYHppIDvW
5pJxktvhWt43A6oF2YTQV6+l6PvzAQ+1TAUM5e86ccp4hnJRAS4ZktMwfQyCY6Mk
HhN7KkcIVZtbeJ0ksXAI5HKQq1BBQ5fNd4aysgouaMYjhPU3K6NzhCh340ipMKZr
77Z4mv9FlR55+fzeRVQ607peIokY1ldIzFRRLqsjxfZm24JJY/uswOJ7w3Ou4huR
cHcJZh4ipTcdIZhPkEC4ybU1GIEHs/pN5k5WIUDe0f5Q6p19CtVzO5QiPAMrObTV
zVVwabjPnYmsJlvQB6r5Z392vHWyO4vozaWwwK94eYtryLV8Aoj1Pt/BscWTM5KA
7EhacWN7zwyBYtiUBydh3Pf45L/0MwsMuWJ9HPWedALfwXicmMNX7OA2j28jqqFz
bqM0xGU+XBZ+JRDvUSb/seXQK9TD/iSyRVjABEq4FBgU3gMilavM/3XSW8Ahkkpd
ITR9J46XQuqtao/zlmnVxQYctLIVZ65PJln2goMy59Dec8iaBJNeuJPYNWYPGq9b
Ku5Oe3DRF0eAMuE/bqGKsBTMSVl8BzRoWlVu+s85sMXVZ4EnraXHmfwJ9Uvo1Lyj
PsyKJKTR0cAQbyqSvR/nCJ54Jy4FpS2XtGS4uVYbks1oHP+NM5QEvGGnZn0L2+e5
yY4DIrv91Mq6EcuRQconX+xbghg/MQrVNujSuaM+YH+rGXqnVpZXJjJSz9bLELGy
6kX42eY0TraIdEGp9tamSiUVPhrmI2rmmm4dnBJPQIiyHEUOWfQjQ14G7WhuSxZs
IleJplgE/1gfxPW5G8uuB/w2QofkDDJmGluNfDQyXIFis/rZ4wNuLX7hnJpb5yRd
HGIvPOw3dGgDR+L0uE1voXesub8A6o0hsrlUekV3FTyJoirEni9r7ZldAiVs6fRE
tJl1CmWAecG12jRMyLOR0s9LqLTIsW61awufnW1FQ2HN2MqIDA48bRYSFrvdE75N
IEjdU7RFBdlVKhdIaeAQepsgB/BV12snjYqZXVtdLB5wgnleqe8NRn11aC1H4Zcc
BFrHBpqgphElv8Ln/MOIHxiY9MHMWz+6WgHeTP9dRl7Th6eN53CNWv0d0tEviwvR
gaIHmyQf/713Bd7ulcHeDIdq+UW6LphvjYeAAbVIyVqUsI4J43y/C5BvM2mkE6Mg
x/ZoKpcI8hIoXnqH/OgO69Z2HomwHys8cf6MGlxAHcMBeFKvVpsqEs9CLTSwbt4c
mtSga9cQdqfKPSshiZ3isL6LJDbp5o8oylFInGxSKu+sI5n3AKzAaKRVCC9JfYNm
kahjBJT+A8r0XEw4DUtvvnVMBivzpiGFPHU9+QWZkTns8GLGqPssUJM0yMRFrEdL
C8G9J3/TXyCXWSI3flFsR/ogOm0QDN0+0iAOFoKMJvmHWnSKa/Id5PXtTefgRiAr
vOw9T5VdmpyXxeUIGPN+ZcgHaPX3UnK85hReQ0mseBsW1QkXAgW9KhiI9K9gb2as
aZC6qCpFNpl6g3+W5J14a607ltysFX6XIy1aBiPA1pXUNe0SQZm9cLmBxjAm+HWM
Rjc09+k8ikKBsmAdObJBQEN4KjC7vNiEX4+cILhjmRlBV+7qOTzAVC4bOv5LRD4B
Nr3NWUTHn0TgQ9Oh81niEQ/zSmfs3oep67RsDMWtRpVH2H8kZbwEdJ4UFCmsIbjD
5Z2mx78ahpRbknAQ1jJsiXSj/cGLc58isIUO800YNR3c0/QDvGXil286UqDH9kS2
iyd9gW2+zzaOTzrw3lpL0iTHo7BFj42M22AEWvW4oBVJtBIt3h8JckL+/E3nygxf
ZZfp1dhLxH5JilbSEgbu45PtCymdmazFiklMmYUgV1IgOV8vR0SpcRlu7ZyZtkf4
PecIv+LxMqFHCPaFlcrbSEaUwjo75Lojd5qPbwG99UmcHFjKEY5HtFHPYt+jASqu
gTP7UWyKHeXkLyW4feOXhViyzrotfN16VDINRKd85MOti4M52zMFKJxeYmVAhLh9
W8BgctfiofvW3QQe+KYLUqVb8/JYRx58uAvXyLPda9a4Dcit4bSlx61e6D2k5OXU
2dzj84L8V+dl0wd/8ioP9jHzcuJVHpquGj170H+Gi/alrK3wlXqqqrQn21EZ1ASC
3IxpfKHO4Z2ck60VB7GyR9MhnULoA8D9+hBDbKjwz9wpIyjtb8S8qn4Lcmahmooo
K2I0SSDB7HCJRDMdu14tD6YL+ZVwmRhgyMecZ9+q1AR9fjaKz/SNMCwqdRLU7V1Z
3s2TLHQq7OJS0Aya+h4HbOgqANfrpyyJxFOTW6jinzFhC/laeWVbTKh3KpGJX7sF
Bxh1e8mGoyuwVBrLcS4+18NOLgUfkHwrU1EW6MhXteunHIVFtnrVBrNUshaY2LEx
SglSMJbimE75wdET9zj3vEQREmNZWlK0HFSNiWKhz82lyP89zM1gBQIU/CkmsJb6
aR/PlqJAVc6TPTpAMkjWxxf8LVjE+Sl4FlHICTA3Uc6MKkqt54hLt1esbqxFrY/t
943bklvTWsm0tN91wWKY54RfiMd4orZG/c4RtiWzvLPkMqH2KRi8BDJxmm3d/0a9
7knIoYQDGhpybt/nssb/TwEUHUalniZorrERoAQjuxvhyjyzDMmrsnZExm6C5ko5
vbBz1BSHZY+7DrfzayuzAwSEMkdH/LQg70pQ0VmReeGWy15DhkpMhzkmQQdGIbYQ
ADIw7NJq2h1SR2wpEl08+rdoIG8neuJX9HxopVwKJuyViRt5qfcrx91ZNh6VGHNb
3MyOk5Krd+bkCgBp45voXv/ebNjXUXHJ1nB5U6IECYV5B4Js19CWxKYL8eDCeUFu
m8LJy4CXttDs5vCLSzzD8PopyCCnmS3yMnLAmM0+0oiH2ZAwyFYY2/AOnpXzjR4Z
lmaPxoEqkeZDzYahw3zVB+QW+PQax6HKdCuNX73H4NVARaz90Wr3aD/EZ8QGtovt
rXQ6g6LqzoMNBCsfuRulXkw6lxvdWmBWqgJWCjDZKjogpVau3V0pi1WKLpQSOCro
POPYNOKZ13nWaWpSmCfTtFispjsDKp1S/SZlZug8U2WfKx8mhAbnNBJ5CXm3WCoW
8tWaj2gZVmsJXYGBq2vLsgKikAUs1yoRMyhH5Pv8hofbzbHbYULli0ALDdfb6oeX
X3uVYsZ0l9IMs6poXSWLktAf+ZSR9aZYFtahwiMGSj4Twlp0lt7ingk4f5XDsOs3
3l5npBKou9aBsbod0l+BKrCSF7sLxV5HG+8fmWCpn1TSq8h10mbQDCI0oanqmqYu
PGoyaaJ/RAlsaAFNJT92yCPpy2piDr9Tc7LMT1aemv8h2SwWLJKAyPeOygWdcpOR
tghPye8QnuDD+H0shCu16NqwqZKoNq4o8yXaNOm2gImIAwiXD09HqFur52tff+sP
zbdZgeHGD87d8XdChxnCnzHe6GDrO6YbBH2NrHTbZGgTaRngymOBMSZNsfH0dHw9
AweOvaHbz6ENBuC94ZsfeJGbgJOL7/sZ4IYIEuGT8GOcgz3gvI5yWzdR9+9EKKzU
kYPxZVNn+eEwYL9u4gvfQ8DokJDmyZI0Tk4Tnz8mKPpf4HHxiHbW/pNnJJniPBXe
lVBXit78OWUJuAhnBhNHxjHjBbNbHGvmm05zlF3NEzbMOwf6gj81MCtIzKsZJZ6X
BIVVVxh/3SjALw62wbkqQFnDiDdpm7wnTAdyZziAoDO5PyeTVXiRVBUEor75V9he
8kORkTFPC1IQIsiWQaa3ad1DjrFM7JTE3fGkQsHo3rd7d4vwK9gmlOmUlC/Dynoj
GK6UA9ZGry/zQWV+MK2zG/OP0qCNEqb7i/rflxet7dZ5uSj5lheqeYF0N08LwMHC
rUgUtaq0PmsHJtQg4alHfL5Y2aM+aSn6t0sHIMGfkwTGCKTLDdQgOAGyO5JNoYvh
1zDZpE2Qo5N6bxK6QD4d+Pcei5yVP/2MD2K26Ctl9La+mlaNVhmvoPc9zCbfQQID
U1hIzM2rZgk9fFD5DBh8LB0IrR+MEpnjonq07wugcmNl0bXzlJOvPyldqhzcbOZx
CSsKP80biGbFNcKn4i3kI9+EOxCnBR43yO1yDaKOKT1Rz7Iluu8VsvkYBaTrEL4b
cLfc5ABPVZKI5gKXHdm90YVnoeBWfC0nDGZ2ONxS0wwfCV4ANS831FbOdKqNQ4lu
qKWY+4ZvksKISHOTRqBRmbetwA/6OZOgQxivfell9inXt0g7H4Q9NvPYkoYH0hvg
ndHT0Cxs01XFz9xTD1UKhW7AIhXD1Qv3jZzxfjsiSQG8ZnKCenQX3zmkzTOHj/fe
LBQZF2otsesSjQZahq2T68MSHhwxOqFh8p587cRmKtZmq9KRXAUaJuu28n+HE7Nq
iqoQdTxgJEJmv9AuzyohXsDJbPm7sM4oeupGP5BKzjSM+FmVeC66SjUDU6Js/ynh
LWmhmdcpNfzlYqxfLAdk5rI05paRdGNd2h3IzM+br50T7qWSz6C8ymxY5emURfpz
hdzdDY0mwSrYSx4bR5rITPcNTkznvPF3secCxmc6k9iFKx1GZ2bN+xRDcBMHXykF
Qqr8iAgK2bJ6uFX1CTMAyUi+AeNP0lP38dSW0V4uYGysKjuTSsG6n01fj558nqFC
dwdJKpe8GgZkZ0Arah7gs0DLn+eqDVglgN7iti5wXq5uYnOTVktq8UJADAfESBON
bTVYk5P/JGUc73HDTA9vEm2xfTv5YS0Zbu6t1nYCqgfYWrpwd0ME3C8II8Ra3GuA
UffoDEto4hTJ7OucZkqqFTG8FenE6gWWHgfZ7MHBCAZmBDF8/PryqcEEDH97SwoZ
jg2AIaC19v2ZGlN9u/x0doXKgywcgcqVhgBUG7g+MyFEXL2mVgcn2BUY0sw1PWZh
f4zlGnnfbJ00+2ZTP56bGNMupBdGzot4Hjve1ohN75eV4MtlxeL37YGmGjO86Ht7
q05D754zxz94sBrO7QfqAnpGodXbyamxAWF6sFUrckHR3VqencXRnhj7R3tUSK/i
VduxXz5/ZHyEYtu5EW1Sibbv1RlqhsJ6tTZ/6TC4o5yiqCB5LeYx++/orrvFRLgP
jxKc0PYt0lSjwuTWAJ9BNoJqt38/9IytbdDW/T3H/UHqzhenQjuGtAcK2gm4Jd+E
nvPXwd1m0AVvFd+pIOT7012niVFqsCoZlNXXH0sbOI1VkhwBWSdKADeLk6mJlJI2
cawvH6hVtcmvhcXCmGQiRq67v7MvfAjvw07Nf4/nm6qaZGk3kJHP49+R8cPf39Ga
83jqQcpeQynUGHzT2EOK8Y45kll2E4eTnqRAJfpRS1+JAeizkMmeE33k7f4d5KSl
DXxXonG2/tUkyjOXGybUIBQbsrkUDtxTfP1/2qA7OUniGQsBhczhXMeyNqovUCd/
8JeuqqAdh24U81lxmYUUaTNZQdYwfHIwZpzfKUs4+kgTPSTM37v3DY0YasgriRiD
O9CL6PbfMbdHD1x5av0ItRsEGgOSPjwMGXoVxYN7Eg46f5IE4Nn13ApGuu++tmzg
IRkkiXinUW5aXUUgbv0mudKp4GlS03eUVBVoYA+LfBLL/ylIvnmYl+TBLIOzAHih
2nHaVQTA5/ERFdw3/9KqzWYLW2YrfrsTnObRGCSsjSrQP4tJlX+JfuVWSwSQjYDI
wiBRG8vwI+iSgxMlYjayD/3qrDxS1HnHW5IBLt0DureuHqFR8JOQLpo+a0VFO9eF
X1pC8aJQoRsyUE45YgzH03prADInOkV5W+Zsy1q8IFdlWZfWh9A2wzIS/jsP32TU
qP3lWRqBBufPpNv17BjFAC5QJOLG6ERpZMN5OmWPn4ZA7+3k7ZZPCHnbk0tpH08x
G7/83RkMOaWLVVttSz/VcixoQ1Fvqx2+kcIT8glPH/lnpRQqDpAMepY3Wu7oSWb1
lTPVfrbC7vTi/Xm6+9aeP7fxHNAUcaGhqSQKeDKL5otg6lRMeLDhu4Zjr5JllQdp
Kr+50xNr7aLLTZaMkOO+L4/GWYqZicmhpp+QYvHITGevzhBy7LghHbnxz2/Wy0Tj
jSe4jnq43tHed1pLsjmGZsCE1gyqyBQJehh1zNkBvsOi2Y/8alI1phHrvMSsTGoT
KjnJ0Z1QWmz9oYt7MudOrtTYYuGlo3Y5hQNSaetsh1yuTHTiqfizV6s6OnQjRlWc
rwtJwAtu1JTbgzaNtT+TVZjLEbgHWuEtImENNvVEq+nGaNkM+lX3tcFn4Vznv6hn
BmxUX4JV0DzBtsIkm7KU4F87Y4CdrimKFC5FJOcfuJVrwRsPL3U1U+esigRpQ/rO
NjQh+13YT7ZXAc3YjEEtwpRmyiT1bixlVv8tetabkO2vv+PD7vT3fE2JNBztPIGn
Htks4FIVrzTYId1Vwr6zQCKGfOMiNG8tWgwqmwJwucKDHx6o9LDbCTbqy9KleVOV
z49SdyrfoMlCqKewVUmEip0tLanWLv0Pppn1eSeEy0MxJwjawatqSTASmSILC0kE
U3wVSVVdvNBMHj6sl8B30z689o3IdaXo0n5jfZa8cr6Rwms6G2zSum3dIbkHMax3
owqnqKesbx8bmWjEGWgpDNs31MplNFhqVw8DLpYDwD8UxJCUTYF0XEFnckAA8yC6
PMN3VM9yyf1mSjrvZklBJTFWjBy4NEKB7V95ZdaH1s06OhacndEhhCPO0eiU6sC8
RCXwoaPuW0KVf28iZYZkATfiW2zXUe5x6/RcemDyOjmuBAk/Nv58WjzJ5jh1cUsu
AA48OKMLNHJHvTwe0zvWXkqIkcRFK2pNd71qLu0vpgX91yKheZz/cyRlQpzY8bpo
4wdCPyV3QJymlUnEG5ZlpKtw1/U5BvS0f6og162s7PsnrDbysvey+RfiDt+dJY4y
W4rqZ4+icQg76+05dPIywSwP+Z5rfNPdp8OXViVsgLFjXq/RwRYMVmM+PAz7j+fB
EXcwcGzfqMjlv1bf9E5fo9MOBl0t3NLFZ99clwtBEPx2Jq1ltCZU9wSfMnQ6VKF8
eUr8rZK/oUOllim1pfWnyq4ur3BCMSpHfVuXRzXJsEsRD6TrCwS6yynOj9Px4T18
YrgGGDXSbOgaiJB5DklO69Dmq4wuhCUfuAmUQnbq9mPkqSgM+KAHodMLaeh5NXV3
LQAoP7XqchsMddddLe1/1a8gBqewTbsbfJn0+hiOOTI6BW/he03HWlcGBtV9dJmW
naFQnkwvDLLYN+JLAoNblh/4m0n/yKs/trsUv4M3yrm6oCZCxOiThPVzRa/CG+c0
NDKVe5g9kL3PLieAe+TYUz0FfLISxRIeoRpk4nhAMuIgZxhYB2R7HBzyMhOTjp9S
VHXXYt+6tikAAHjN03/Tk3YxndbGVHgnqSFsU3vCnP4t8ZCxE0ypMwjeCtvYr+FA
CMJrMqPjBTLM5xXoHSUnFgEa9YOEuleQqE4Y54AnuH2H/eNMaAEhUBJe/zCbS0vd
Oolc2E9t02yIoWSEcVhGevKaFOmIQhcaQDN2GGk8LDtP+GE4qoKt+PRRjQeSz9Ea
1hYRQ4vzOFJIvbZxse4l9zsU7QWEfidH3h0Bj8tdP1f8UnlYKcd6Khzd0NUVP4Xt
pkrEicEjVs60aAmQOeXJZF6wLMFkUqDzp/yLGMel/4gtPOY1wMwfiMLkM+Hf1Xc6
Vz0K8NcDSTv8v/H5vtUS97IrKgkULe9mQX+To9Xqd9sHJALVuEmebFGwBIlusERK
frVn9LZtAzSq29s1ipM/3T86HS1qydecO/qwtoaIrOamuvbjxEGrOmAKbc2awrqB
39r0FCPqjYdRqL3toK0xC2KCSi7PkeTFw1MfoyD20HCcFcW4OM/AgNfeyVJMDXKq
mcjuNfICrXaDr58FJ8lbQLU7U7iDanjGE+v9QyElCiZ8I3Q8LPH6wX7ziKUMpqlr
McSXsYG4QDpwqUOlPQ9sqqjBr9IoEtVXufb9GzrK7CgUPP6sjQLv7mkSAOtydoHh
yS22mwZKTz9YabWavWdF5SrEUXPT5gvna35rGhlva2gEJ3F5vC93PErW4oOfMjXq
I4Gg1KLs173tNHpkvY8l1Ra55MmaPbKc4bJ99cV5vl8U4H5GBxTeFNXS/dWnpj+P
kC/vrj+5AAOsJzV8kbyD9yE3t5/JigN0In6oRFXdZiH7AB3n3Mxak/UP6tkTtVk1
ZxUjEXg4b1gsoGu0GW8v+Xn6ZO4CWWUEahrIzO9YeTQMtJPdQffUkJZBTX7VRVVu
kV4y7sA2/iq9fzK2sLUtJy7PgiG0UVbCqG7IcvvwgFC/4Qsq+VlCXbTzaLUkgAy6
4R58i+JoiHfz4CJkrG2OceagUjPotnOFXWP8EXtbLgKyz6zzLD0qIl1Eup/uHzLc
sDdoouW6RAebiZUrq/fBjG0tt41GO6dmKVJlvLYY1z8L+gx73UAsFOyZP9DkcBa8
9DXBCTw4v3DY6Fj8QljOsb9iasAvdDFZc7PMJfh0GrjUM3FFSKKMJQZd1XDKYHpr
uSYhSPVFN9PlzL/kYYM106CjORmdnsjvDcJVmBAP60PItoIO2H+e7c//+shQlCRZ
QqRkz/4bkgl8QiltwllDdkNYwix5iUeny5Tw2WakDMPc2ZvtKp8BJXP+bxiKXKgW
3DMUPrPNku1hpMjd9jPJCcxURd5215y+mu0ut2utsKIY8fpp9RpXdKyHKwP2Livo
uo2yCk78tmg1nfOqSNykP0nim4rLVEpnAD1YtQtE/P7y6hi8rva6JqCXrPVu/4WB
beLEv7YNoGky71d4ZB7ZnGgogA8LAyOK5x54RPlIItmbdc7KTHn9eQ45CDhuQoPn
NhfF+y6tnDMaB4fKF6Ots+mkzwcgHTk88wvvR/X1fRjJGL42T3Zm4vGRQ6vRhffH
J+rjZWo0hFoX09C8HlsHOf/+Z9q+lGk0cRPapaNPQX1iVWTZNuH4RcPzihMs6Uny
SIG3mZnBwqwyH3JLEY37QeGfake01CFnGLi1VTi7zwM85sSpbG15XQkfekUkdHaz
gHpPyN9L6jX61pEWLDPek6YVtLLPJnrtfETlUKNwFvMPzZjQLYerw1I6Obl2zgNH
kvgYKEdlvbbdWn47AAmDp7u3vpjtRWmU8dXebtDbhkADEtLzJuovAY+vFShlq3qf
Q63XkrYPyViYJTlwKFUS14QMemN9/uCgB5xmV3HgAa217SZ/yAcr2zpFWG3NsQK6
j6IKvi5Ri7pykkhXVoR3+k/+uguARzJ6cMqd5zR7w8IZhxGtXvjBtRPJryaqTJqZ
3pkvjOVAH7JZGOg3Ttjg7uLAQEB/lADI+0Iru+f2HJpx5AmcETGM9V+pXJHzMbwc
tE/NbYGcebY9aecBtzZhfcub0EnLBQEubE+NbYVx3e5BSihgdTthQnzM8zh40Yv7
FLfFxXmPK+tf4S32dPNKa1WB1NtvRalUp2zmARcmXbIuAXDDuBOfu/2l7BRP5mJZ
HXhfmFAbdH0Ef3ch9NM6m0dWeh28OTWpogXvgLgw5Bd39CU0UnW32D2Gddg4vGc0
Sr6UIEBhmN6MC1c4Lbe+c4EhkVAYk6arwsG4r98+OSv9c/F1MaZWvRPr6bdF6U0F
jg+Fm8hHqnA1OM8amFv7tAJPsjAPqkHykNfIDVs1CAP9fA+Uol6GF3CXtuPvQFkA
RQq5E6ANvc9c1Kv/+vHBlh5ax+LJNfu8fwRqUV/7AEcP3iWM+zor5wZtwLJb2YXH
ou534wYQPbN5rIEOBM7iWkv6t+f3B5rB372v0xkT0rKJSFzgtF+GxmFd4iUGEkwM
0GDsQMLOamFyJw7X3GOmEs0AMiBUQcnIfse2kax3mNsHrDfYfqTaxqU1w0onveqF
IPJM67j+7OUJVvn767Matfs5Knlqt5AMO0J41Xeo1X+2MVMMvkG70dg4NdPDylqe
ufVx7aZNTLOK/LyfuoluQE/Ze1Q5g8GfCrjGReEaMqwlPlp3k+qDM5SYLrvIU9su
6x9bW+S2ASpNo4jJF7G/aTXuomqgIFUlesqNVX9jrM02snxoUoTrbGV7OpPTOGsC
eMzn9wFJOz1fy1mq9oiJM0DhjIQ2mEH6dyoIRLtwh7xb0Us/UUNmZOKWD5osfi0h
5gOC+6rMV09xqqD7JMFkYQ7me+mdh6tzVmn9wK/SaIsKJvQm+6mWziY8ggMByu0y
aJmRTc93OCMaV8D+BHCnzI0R24qhP3hO557URlCnoCOddyEroRXb09x03B3YCsuA
sUsounDADD+4YS4f/V+LPQAVrbwsBtwMoasm4ws8MvNumZ8WizJmY9556Iz8HMe1
PIa8/mwhbrrw42+zSlfLf3/ncXUvtD/tGzJam/gwIH7FlBcc2AbtjPAgKtOkWIv9
ja8HClwFMbqGDrp/LAF8tK1FZCASBYASIDQacaO/30mEsTKm2mgjnoCVh8JNv14Q
xZeA6/7okYAIgva9L5KJbrwpC0Um36GP3rmgBDgyJKN+gMUFbToBg06afw9wXJVt
FfEjgBjR1S/Z2aVd6EZPp9Yk2fHY23gR1HLtAPwPHCx6W7pXI3NmMRMxHCLgxUhS
ONYre0jdnZcUWAyBrQjJPoJ5xdLbvU1TvY7wLNPBRJGPmgOSdN4CsBr+ODKQLKGN
YfH1n/mCvaKq4xo68JmjrdTbWN7iTAibxoHDxNt66+pfAapvyIghWoUOj6Zyl/oD
+RMneJ8QbBj6Otbwt8r1iXFzp9+ApEq8SzTgzIKnoRlFu4trAl5fCnXAJ9LwfO6Q
MlnpUDx3fmoLSUmLejKSRH6+TMr9lT/5S6c/A/yRgAjrxuYkdUoIGa5sr+RdTpfH
feZ5ygtitAj9tC/MmqYB0GQKB6h1NPvrzQFrDgZY5qQPcPCCe+WlwuPoBgNrHUX9
XFeK6S4dnjmcrW+VFWKKGuIW0RI70RDPecBrnPkrFTx9Fw160dc24TSM2+ZeLXS+
scNNXmzU5KmPob7YNnYH/JFZfjjed7pLk8T5op2n92lsNrWdmK+Uo8Ivi2bl1ujC
6ho39gRR0YZrFyks1mysw5TCpDXphoeWbKTg0wvw68zIaNFwOgWkIVaRRgKKZ7GD
Yd8X4Al8KJ8JJR7lrxZ9bD5Q2dQj2/X7ybrGXxVBEANjR19s+HggtrZpXesrAzj4
OA3LXUP0Aw2Tm4BZvNUSfZbHfuHc/3lt5jeyADCauC4pyn1zIpSEkmdJVEeOlP77
3AQJoXAoH23Nl+KpH1Hm7Vb77KZES7ELD1igVc9+TyO3LEACK+TM0ORwjsz2NjVm
Nn4p+kXWxX5YH6l12jDUx8T0gLmOco2W6n1lrQ8Mysep2+n9+O0LLEz40BX6/eyJ
5Oe+4BpSlUKsRowFvh21iyyAYFDrUARTU0z4qgNnuHJemVZD+iW/+F7B8/cy/JD2
Urh/sQNLWuomMFVvirSuCYAOTVDFe2ByWPYHlng/J9ZbucxqPlaHoS7b2us3yU4A
V8q29Maw5JPVNvxTsrgs9oeam8T9GuFGpEdxODlXJJb7GZPQmHgbu5RSg+PfRrF4
KQYbHXR1wRp99KNI7gTvJaymxwrfB9lEnixfuS47xZtD4XQG7NtS4OEQ+Y48hYwI
yacAdYhgwHbFu9rmcptJnjTKJgbHjLniqYNymjEYNSolJFDbadOJ+RY9OkcL0sYl
gRrUFlcskDh79g3ZdmAE24rO0g0MmxOKMrfwHujeZG0UqAjtpBcWd7CgqEjC7k6x
W9cHGv9vj/7ZPxTmYSxqdFFZsj2x6cSnNYf0JpewazijcEo9ir+yxKwuNgxg4NtJ
aaBXBQoCvpM2RTyDSEV6WgH9X2rfsdlguO3ra7IO11leecpvC+1XtpDeMRPqForJ
dmiOzcAQvyxeYD20upuA6j4axe6OYk6KlRT712M6duNaybv48WwDY8cUbGBy5CKQ
Af7s9ufafxxstOkfJK2CQU2NXCLv2+NarMPbSgYFl4z3TXhYqjXAIxPt4nvkdJjm
qmbRYsQnWsKAfLtrCB9qDupg45Ujd7qruPcEjmkcVzmYlviYcHOwQMTeVqPAx2/t
Hq+yr8K0qjIn3FGnBBg5qekCC6UZszmSzN/WR4tERF6z2ZsV9zDlYXUyFMlaGnQi
dGpiNLscR17x10RJdlG6do0yZ3cfgs54uecBnFifpKmEh6hNPk0jTYuwWLTq/qv/
S+LunAqL+4CyLtGu/pF0x+8lJd/8vgzKwd6zaNdnFhjdUggwiEI5sj2P5lIEcbCr
pdqtm2ly7TbAZig5bSAXY6Y1SnG9yjiY5OPuea21kqhgoqj1aNvjG4ZTlASiIcSy
OCN6Ksf7txyHCl1iI1zUMXiGsO48VIb0t4EOdWzi7M3q9d8Et8b23yb0V4NBt2NB
x3iZeJIrtSdnOKid2fyl7qnBMuZb99G2gzjLRLh55M7HP1obLmVHG9lFO4LpAjky
JMDfZ8E8guBb24n1/gqyqlX+IxCBKlUpLi5Xolwoxaj10PQZLzEHooE7bT/1ZFI9
ArkY0ZxCdm5OJatarzv2VTgc9uON2JtAfELQVk8Lgxzz80waUxziFlXpbb1hBSAt
+vdaVQ4Rg9X3G7QPAW6igiHhExclF4pM7waXyeY/RrpqvWZUqqr+JkwMxc7+IU6p
VoBT7BwIHO7vundKB74z8qLof54J0dLPhizmMd40foFbNFjN139qhN9y3+fivVYa
mOiPmLFhFoN/VjVoJ4UIFVG+YU42NAOA99K4qNfPHwDVcGHNx+bNd5u9LHOSToqX
7R7ffl8YHE3XhGa1pv9MPBVUEDkM8IpZHZw3HOZ4UtCFfhL7jkptP7mEmkHBgujR
S5l/oBttP3LovC7ohPiHT6ZwINHzT1EtWUHJqBAwxH+bGCUbaSrKYTHqCQXDxP8N
AVVbEtC7Vm1dGJcnM8/QvKjx0nvWxuZ1hH4LOFrfgmq5tsr/E++4HOQ2USAmwZOj
EGU/oMGCmwWKWoab17eCanFiK3anzGAs4FBrEbx03cFA8YRR4+UOs5ZT7iONg0tl
Pt938LEljepw4o5ime9VxBaN3W7rO2Pu1p055qg7Puwl0efh0tdg8i2I8M0Nwza+
4QkXVMBs4i2BsxR2Vk8QV4ZAnklikmteL3Gb77N9RrRanX8895znLUJLgb63fUJv
+qt+NJUyia89AM6ZNQ2poSYyPntVuUm20bOTfJfkaldRPesiO/K+sKG3P0LqhqgD
3Zi3Hw0gO0APqUuzv8DcDjsNBqUc5zu/5wahu94Bq4HkXGNLyK8tMSQlxVI6dtTh
IlLbwt42qK8zc9lB9X9R9g8flzP7DxMl/q9iu0dkFscw4mcoJxlWct2Fgf1GDYQ6
K7gnD+3JSoPgYHJWw8XooghtsGvKzl40JRVTZW5vbGbtL5Sl6BYwJhtLKT8ITx42
oCQDU+yLOzr++giIFLj2br0QZ3sMGd8Qo/RskBs1VQehp//l8alrdo0R2x7bHxLt
FutaZTqMy59XTJbD7VRjSaQ04htXV4EqQ214FMAVAXJp35m6CoBmOXoztTgi4xj6
5+qzazpWQbM3xymZ7Ws1hm+29IhYm60fHVa6lDrgI32YubqA4N7zL6nZUmkZrFO6
9GPPkkRrSBINcLJbP7Qj1zOo2Bmsz8RYKb7loFyLKY6p+15mhlqIzJC9i3MyLXzh
B32OQBQ8k6PZAoOimmE6oNluVBRF6QaNumHk48qbZt9k5uwwP7hDzOcCf3wXgqbG
0orkl8ZgZkD6ZGsWixHRU8zY8Q6s/CK+aWR+bhe321vbcFAcaaP1gCQSolwyU8MO
k8ZhJw03/lB76iectApyzckDJwRmeFlXmlYIGQPh3m+SdolMsXxXugPD4XNkr748
H/l5ADHHJJuyYE/huLeKUDq4OiScDgMovD/ccXhTidjsqy5EI2bbZmmlYYcZFZG7
5a3s/2o/l5qfdHZbVkqDqo8wV5Y+p9Za1fGVbFQ094URsh+14qtt9AIga1TRIrC1
RZPTOUkZO/uS3k0bv8q147+Ht2chaEhBRviWnZ2ZXoLjVW6S5E936UYDtXyaTC3y
PMSiLmv8v9tX1qrtJjZdEA2q8AcLlLZhXiGrh6GO2IA0GHKoPPQh80WZpddpKaEO
usWNaQtQoX97sDUrVEj0r5FMMj5MVddZ0HLzNadt/LX5MSGkkOM6RXztlr08Crdy
4i0yKukQmxNijWtP5XhfTqTZqgUZMJ6mulamndvnnot+iIkM1I/ntaakYd6Ut9EH
nQ6wA/0pygRLKwl/N/otmQHEOx6QUUK3Ljy1BMyTx/8+snCGstyXoqn6p8zCKdfp
kCrvotTMupJQSDMm/3cT2VaxMPW9w7YzH/EtQRqL3pBKhS4+ggAXfrImjt+IPPJK
FGW6wc47aqU+h9iScPQzZjkaLQ3ppwyWA71OVywhuSq4fvCjuYnQ4B9fUnIbcZQH
VUx2nF7qPmLtxGnPstcWKhdPrz2XA+xb+3BCs3Z6vXIhLhhqDGH2D/FDasFF0xbL
nKEP4DtEBg/7tMllOCx86qtH/hyMr551E4XmpPhE2H9ViAzfK1Is1vrODBq7Wtcw
8Nj5HbJSFHJk8gxwJS2L0ijjnVcxqouuXotYQGG0ebK6GOTsJaE73JXDjo3CTaVs
/VltR7bi7xXUD2FdtUmm4eGQErU77q9DpF4fKqNpE975iMia8RAdPd4s5j6cVbej
xGSaxHc/4HMOg4FnkNHTsmMUtnYPFKO+MwrOPmgNSP2prmq0N7Cvs6r+pSR5R0Ni
hxVdYJZ49QCWo0O4CGazfKPi1dkorfk75FFY3LDV7exl18hCnCAZ17RuH4Py0tn2
efXc22xpZ/Lz5G7sid8Xm30yqCXyv8PdwddEd8Aj5rqh/gWzDv3Y7gJduhWCfPxU
B/DT56i5dA1ZRRv4N+PYFyop3WNsTWLsZfiOPGHkfXp0UOTX5WgvMXW6ew5Ycjjr
T8yNUpn4eeVNUUz02IV108Me0dSJtxjF2oJJ5UfT6geOcHeERt4DC+kSD4vdKW8h
LGOhTfFWLDAxYUgTdava1kfuSsmGjiuaaLcSs/pE2OVAtdTDNauAzlIbfm0eKFlG
HW7vWDH6zqsUd/gFFlRAho+OdqSSMHah29pJf6t3K54EVGAULuv6LAXosKTnWpjL
XEpVJXhqS5bfJRT+2RxDV7mlTJSlpTq2FZzXpuwbd88MJeDt62E5qM0uOOl8Y29y
JjiiZ8ckJsuee+Db23G2YtOFs5R7Ekc0/Qa7P6B5znUpRFgrLhRUswaqXQCEch5d
F8U/LvOEgaeOPwcSMrZHkReykncvpdU+ffhwqRHH+T/EUG1ft2Za9G00uwNk/SpY
5m3H7uXQXyhZbbyb9rwv4DUUGc/Zr6g5rC4BhtgqgEqed1+FJ7bENFgvsYu6tKxT
ZcqPvSsHhh+v2pPYO1ARLANfPDzEm7CIP0YwJ4Zl34EmOQB0q3uK9rN1iOW+Husi
F8vtecbAdSgkW3od/sHziSlRWgqX4dAnsQ6l0OfyRrGmsBzncsgt/pCIzLENBgxu
4oFSR4D3IjnNitMW4np7gtzJ+nzQ67LYXDvuFGSRFO7fBe1r9vEti7v0HsbviQdy
0fmi56d11BVg9auTyuK2zHargIwBxLPQUqbz2vxAdTqZhpUzqvGenDDTYtONZdxu
iy78s6FQw3igi5PdtuZIyLnmmoOXF4gKGN7tS71J4lD8GX9Ey1on4HZTPGcrSuAK
4/ZM/TFYRw2U/DhQgqJ5FVIH8z9K3HlA78d9xP0EOoeRQW7alNo5IAJbGV7GSUGS
hvjt5XVjYEomQPeYnUpmo88zqTd3tq5NIQvutq2xfq0bZGljsoxC+Fk3Y+h3hylQ
SxdCzdca3R4XdIrex66lXw261pHNlUdRPln5gS8L2LAJZVVY38QHc16fCQY8CklL
T12k6fkYCNpYw3hBU/I1WA+N9ET+adC6EsiEXFC5R/poGpv68/U7Fqe6avkTEohy
iYwztNfBuht2gCbt1vMIhijdRKd3fqN3VGB9rHOVBSRoCOwCTUI4fskJHcHqrfSJ
bC+d6KeOwAo7UtAIMTH9hbyEihKWyJIAw4tkap5MU2JwyFGh8P9wII8CboQXTUeo
oZ76Fh7IfOEPb8L+gmjqY7VsWzrC/i3y0YlRv21JCf+65bASePXgfl2faQW9HLhX
LK6X2DoStEkdJVniw+FboYhMfcXcC8tn9s8AHyunI7gdknUvsiPbcqweg9kdFaM0
ey0Hmy8+oHy3C3ahlXSU8WMLOlQFkYlCYd4xdCvyyG2ANLZD/EhIWZXvI/hcy2Gh
HMG3zzC4+Izq8DrblsAnBXPIvxis/Z2lHlU+/I3Nyq8oT7L2On/+OD09etUIc2I/
0niAmojo/ArO9slGS3moQUcE06fBh3hlqRXnVECnm9LqUk7xGmFlDe2H39/7rAgi
FQuLD8/G8qDhdkAfko4v9cuhTI1HtOtXMJIxRvi8fZRQdiHnP6+BOdIbyIWx03cS
u4ekGhl5m2UlXJqgcqekOTSjLELCf56vq67XUW6KnhrwIp0bZctBEwU+TCpzpPFT
q/w39lwUmBPQQv5E+kc55a3yUynoIEd6H+iOorkX3h9SxcvokiyTRbZ1zNUe3AnS
IJglsP/spDM8rIkPSgbbqGI9Uta8D0Y6F1Fdv0estC9gT0jX+rlCjUUVd2FLBn8K
z8hvINg2WvLAENNdqlDaJTRc7ab/B3SQvfkDEHyi4NXa6DYHhaDu8L+fD03hRJNC
eWfJjFxTPZ7uUKLCpiYXtR7HdjVttp5kZO2psv3vbVe9wjdKHM+bDzUqlwucwGM/
INL97E2LowHWyULG5Sh9KUGLXfsA0Cw/SKBJWyjnmSOuR4U/6c6yZBmIq48wB/eO
vt+dMXvPA1xA0dZ5Pc+H1pWYyqjJ6+lB6gB3aHbKfWHsCwlJhIBW2fPDVBfCPCtF
3iCdDddgH6xaeSJAzfAGgWNeaTpKTZrP8zXeBi5XdSsWw7x7ps4uX/06vXUAiCIm
m1Een4V7JikswHV0suG7DSVVeZZOGVNqk/1zabmY1GF+zbc6My6n0K5+N++2FFFy
yy+vuNcIKteAq739c+p0KcdtZs7jcthIIEEq72pvXoEN+A5c05Wbzl7wJ7fq4VcH
hX9Ku0hyRinNaDs5q/H8vmwxJBNPLbUkejFDt5Rql8N+jGTggudJyu5I8VhSWWMW
MEW7Z+/NPx0nBkMM9RwM6bFLEhDSU7SDUJBgSpJ36wGyO6NO1QBolsrHLA4As3W3
lI/0/0ORYYCpYYoTuv0kAHOFKCY9R2nPyqrLAhxlQKlQJZqaNNrbiLUPf2bGRBT9
IXMvqD6AQQUztWvkUsy5pcQLZ1egHbUji35KGbKenXfAqYnl2oo4TdBbv5tzbRKI
mpAjcVb/rsmCcgeHIvlEQqy6KyOU9hjEDBNwhZz0gQVAbbkEXsOH3jupFOIkCqVv
RqrJC508cPYEcZpWgl+5rwHsLQGIdkBQyuKzLbuUmPMhTKDIbOa+d2s4z7srlQbC
HcxCS5SiuWrJYQDb6VuQVgOGliKjuSsiVFpS5NOkGGoi0Vh5BbncwMM17AD1BSL3
Xv2+v6WaPoqsJG4MX6wIYcCeYOjnk+CsFLJ+zZUiJNrSb5r/Ib0lEmNwPgkxN5AK
x4G3uoJB4VxyNBcWSoW3SlS4x3hGepLpMPxCiywhjSEWl3BdAhGlJbwVik+pywel
qTyV7Slb1iQtdjpjY2gj1istMENP8BMWSM1yv62PUVn0MeKZbvD4Nv+wg1Gh6pJE
7cqE6/KmBkEQlsADX98TjcvHolXDVxSsllgO2YQjWEOSC6uUq+gEbN1lJKTw/ffO
mJdWokuzAQ8xbxwcgHVnTakxtb4bR8snvDpBgNr3Pl+N/toaImYO8Khjz5HKBjur
YJdDbcCNsQkyuFh1DNV9jhul4G21uwaYTcp2W6k8KOB8lxpIpbGBdNJRpgm4OEnv
jOiE6wyD4Fp5hb2pQZErOoQBNddSiV05dHgMBZnVakeD4VHgNlNKcJx7hfCqhmgz
4yEy+qM9PIjyu7BnmDVHkkF/xDwm03KXwFPYP/8YNZks7KpN0rTvohKdkxyIqUvG
q1X7blS0nVg6EyCRkFi2Q9T9JvnRErci8rGd0XP+Ru60ygawJMYOU2Z7s1Ls9WnY
5KSxfax7FL95SSgxxmoVrKdx5tVWynyovkJR5Kzg6zhzjO4WxTGRG5Jz6vKaBc/L
p+4JyoM8EJVoNOm+gz53MLbrSLgbu0pL9cDmKK3/oT6FC8mFJdslv9RlgUGCcfyc
94ea8wKw0xXi4C8RXhUZpXsLr3vZQqWEI1rXLc4+gcxxsc3BpYTFuYd28VEQnWIz
C7bMXXLHAbFSptk1CWzhE1oyF00a3IR/1hjbPggKAouRu4wkB+cr+bExHw6rBr/H
gUXuTQ/xFLuX1vqUn79PgfInJMee6Saw4aD16SH7MtkXsWMLPkNQARG5uAhoTn/I
rO7GlNqAercFz13XUJx3jXr/HzG2Tbz5Y+9OG5po2s/YjQqAmoUGUoQk6LbNEj4b
5OVKUDvy8mHqOWXbLVjVH+NPENELCknFG/zGEp4x7NTaOBbe+MeV2+yeHQuI17zS
KmJwN6AooDtJNO4MRAUoxdiKGe+baQ+OzFUCv/1VGjyLwldtCmKP3aCTM2VBOc/n
D9XEv0X+lFCYYK20Z0CwDHHeVg3I1b6lR8W42xndglcUv81LSb9sJ5U+n5RhmkWS
Sw5U9KMym8qXL1yrwrU/N7rd3o3DppXV9dAxEDrHD5t4rUJE1cd4H1PP4iLxDAFp
6hDg9n3Rhv+2xTyBbRFOWqXAJaFY4amDKqbuoK1VYAulwF0gFyWZCgGpXFJ0gEdN
fUUYwAiq1wo7wB4RmPM3MyQwxu82QUnFL8y0FqfOxcd6y7l1s43HDckAQ2Hr2Aey
LHxkZ8LC7d/4u9+H5HEo9gcmcItJDkvPtMHAJ+5rBP1fT9h33S1oEJdUpU6HjUBB
VkFkYatjZLzNbXzzulejS2vRqjSKRcAL94sX9PLaiRGX9MCfz9XlLK49hj1HnQMV
nUzouIRGsfDaLZTs6LHbxFCxy75F64ImnUFOz2/6XPvsOXedZxRR76djLH6ZcKHx
fsS+Xr51093N2eCH0sfV1cKDEwgWRotsT5vUSxUxAoEphAAm3d2URLH/bTnxY5op
NXJoAjslk7XMNTBmVkYNdiPz2Foj8LpWC6Ov329rgf5NvHdf2ZMMaFQTOifLCigU
qiFH/AwoFajaPnXoAq9b4aT5uNtgDUWcMUK1FRfhb4rpiUItBBlDPMWcDYX62uI8
QRbg2tZ11w2qeeFZHTBpZPTw5HaXSOoTeoqz6V3y7lDDA4ZzTocuKrfGEgBRRdm5
6Bz8S4WBglPMa0tGn6yXhbzq1tRFArkQxaE5/jbmsRY8/djYM3sbABRmKz+1HtBP
K7dpwe7eYlxVzgiGXdyjePieDhmqlXxLQ614uE2WA7UwfmPaZQMdehUY22vhV41f
51RIMGp/KJqgfP0Up4vXyRIk9Qmy8RJXXfwyiJ+FbUW/irknzSnZKJ2q9DG0QuTJ
o7C+w6CwViilN9QjsE5zZhgX13uBKT6aM65wQmSUMk58zvxLelClWmARUqKD0Q2a
aBI0GrL8tYBcsgoDnIihEysfYUd5y3umjVGOYFJUDl8NnTqq1nBbYqr4QTRGM9+m
uCbL8cnhngPLOtMrNGMiXNwHpCJG4wPIhGjQmBp1k5O4AM85q/2c1WPRn8I8cJNh
x3QpVe/vWRcCUFGmi2F8L7f2v5fgkdW1LYWSbRw6kCYN3PkZ2jNJJkOE1LMRKFdc
R9dDoy5aZ89pajdScx/uv4bCbR4lkDMknu2UtwD0ApRFTC3QJxKRLiqe0zX+TfQr
yYhewVTJa3qrLdf6QTPeO+Ncl9rcKr3ZASY92YqhsmOsIq8TwyB22NYW3sXrksq+
gyB21j4voHAAa9Qn7ECIQyr9yZr60Ezv6YlBud6ZnHf067MGe8JEu29mCzQqVA7l
R50tsUDoqr4pAcJSdSzfW/Plz+9gTrgnAh/LWqGowpJzHcwoSUUunG5KR00/y9IC
BFTWDnfRxD4K6qmY4dZNiRO7pnCgsVLq2cHkitUd4WaxFwAwYxXpIcKdCqWSywlH
0awtvYJHjzoh8qCrj1jjNyirnAOppfJCG6xP3bsmXbA/jK/6c/23OPKRJULg5vbp
veXqM29x5OulgMyq8Dt2F2IC/YQSV/G9kXpS/t875c0H7ze+qFIDJ96Zvcifuhmd
KXRlHHF+26nQTYvrpbkLBh8lkInhw3mbiYvyFjfnp8+dZ+ZohLeVu5fmQC+3ivLo
qj/nxHi9Tg9zi3OR40vhPOtZs76Q4CfCORQn+gEaZbvptHQGQ4Kr4THJYYonDdR8
4A8gr54ofjB7MQujrhUK72LcRr9UgK3klWOFHCb3X8TwANNPJT1mRe7rL14McLvT
PGpnUmWB1kaGVpo2/s1lI8ZySXYka1pt4Sg0bcSOHn5Vvn0A5KCVcbv3tXrhQIBa
X9ju76Ez2RDrwWXRMPyTy/bIDexW5/+L1sEIsP85VFTOz0pdeAzZOUU99GHty2RG
r6DqnJEXCx7jNfDVz6AaNSgfNEXhd/yLCSjTVUaayCNWQ4wmJ6yB2glivpj/ZIBL
jcnAHKkstrwdfYahgwIU71kCCR2r5ptakgSzMIq8v5HGi0Rn2cQNDmnJlmhQlig2
XFfG3RukvFOL007U8dvJabozghZFqLRahTVju0u98EG+Du/+RXNeTCMHc2mOfjqK
kZ2siy8lqTcqMqSPd1O5+KsmOEGybHB6t8fnBpg4o4zYEvE0X+n6KJNMYlrnnlOd
Q6+m4cfYzJZDLTvo1jK/mgK7UTJ914nHAfzQdoWK9RVs+tvEpW8e8JHFdWAre92B
k5QEHDIjWz+iwldGgFUSQ6BB9QhF+SzQLFuQcx2Ln4sEfUystI96v9jNWtNXYZ2/
aQMB0XFsZkddBroqDXWeZGxi4D2ffaL3VD71ZbHd+f9y2ss8/MAiRYqUHtnTSOjV
VfXU/w4pcmMqvKrAuX0Zed9HTvgq1E3qciKPtpet5+QUxMRcrgtVssz2U1Re5/Ss
8BZjVFJLamvEoWjP+S1yYgHeYikqj8o8QO9pWBJP5rTuOFlDRPL1qp5yI0dgiBHO
7WOvkCND+XsU7yxKZDr2sAk+Njet6hM5CDY/s+vLxGPzzSpJTj0zf0eH4+Sm0w3O
gamJGaB++EUZRyXCUdPgqDeQfVwhfTYDe8eXYjamwYf/4J+KE11SLMqCYlh1moSV
N6syreriYzLkbm3eok4XAeupSB+zCm8mKzF7ZRqSHsVyyz4RtZhUL7oVUBpiye9a
p0+qgWvQov6GYt9GOiJusS2nkS4znkIQ78N6cStImAFlhE86wGUNkUuqZLwf5XZa
kONKFeE3Ezo/OyZ+QjIgOvtLuk7BUxH4NfJA9g7PkWE5qIgSPCqNvcE3orQIPytn
yyB9PkTIIvc+MGodhINJX75YAgvn+F5ovTLSeHNA8YHZRb7Du7otDsGLJVE+4wCA
I24uDTnpzOJ8nD1kYRb3DExQiQQQDd2LhwEO2e48IEzgRsvCZwL1x5ZJ5AJ6eUSu
oscPfvSzanHFV2T6ayFDxSUaHQMSGD0S6/+MX831jmnMrSsIaWRxv5NxLs8VugNS
WJSOCjO6xukOhC1yrDAeKvKg4ZxG6rhMofuVxo5lpHzwy0nPoV8VkMAvqdsjTC5V
NQmEFNg1oWVGizsBSxox8Mb/tJgC6k5ngyAR4Ezp2IRtWfkObPq4SVjQrKBqhPQF
XX70PmZROcYvpxWzgUXjEzkLne6o2wec24BQDYlo+NrK/vfijPaPl8x0sSi8aHhg
HuU91KzTr7aXnS9xAJV5c8c39KVuuzrNE2xzx+2NGJ97c7quP7BQvhdgRESRxptb
hYkIj4kpry0kGFBTrwJ3Gq9hQaGVUn9ifpOCh+pEWGbIcc353igOb7MATD565IAH
AxoUZMuil7KAtK5TsBlpnCgjhMfGrUFyQuNVz4TWwaxekSdF1dZ+9yQXRQoLgnHM
+sgccXdTdMi7DUdtPxYw7QETGBOqIScUR6sNngqj51Lk3X5eYluxX+o9m4KOG9TV
w/GC3L2izH5/tx4J9MaRPvIWcWhLWSS05xfLBunPn+9Q4Q8w83lhetbkvpaxAMUX
zfUswbrdQgaIwP9FiEdaIqnbX558jgWPKjX5LTZCYhXtpX1gzO1AucTTq11SWdn1
LKcc7XvJx+UccacRcduj9x3HFpSqJ1+Y40ldN9ajJu8HnnlvNvMY3MwIt1USB1fI
YsavmGGS/KzmuCkPJmNcltsLSJh/uxYKtDaHDR/glMpp3LZS8QKLiiMi+PBZ8SKr
KAP0V8QSxGXmPdJQ+fQzi9kGYamLx/D8UKEz3ETRL14lJrN/ZBmgTnvTYqppJu0f
mSeWOkfvEsvMxwanti1uewbLduKS4A9qTKSGl2B24dGVvsm/8FBqDm2JRrNdFYEL
yMAWFYmxtz/xT8fg9s73FMBZOZVNeTbnj5zFHBjrgRVY65nSxn1ggw3jnRVehBS+
wIHkVG4segJAlbk75k3pTXNtKREDPruM9CSjO8dp+CXquDTZoTZis5Qxra4ELWvB
YRS02jp+1xXux+bmXi0pKgdAiUaJrNEAawfZNWt3EInaaraaO5xnDuUTFAvZkkX1
lgKKDgT9fWur3EzdGeRYUL46LnspbpauA4yMeu41/WK8p3VvLJ+iOHO5BwbWSwRi
Bh5NQk5yqpj/Ku+f30EAKmMOoB5/Xf51NQDizkqaiX1MACHro7zTJc4MvluTvLS5
A1GQRO14YUI3+ptUYQSQAFJRF0+F2m5YYEXjnCnnzSSsL6EsH24DscYJF/EeS8No
d6K8jqvw/Q02iPVUB1o1tKk5CFXT8cqB1lgH+xhgXj0sGBoV2caS/aGCSU3Mf/wJ
NYOIsImf+Jdd0UC4M/Cbpv7usOIfxhE3SASp2BgJkrGjusQMSGP6qCTuo+31QWwq
wO62kHsd2HK62bPV2Zc0/gFDHYFBMIVbotFdSQQb79RM+W32jYpPaNICBh5HWdeW
b6RdTPxWiwY30Ug4J6qlhkra4kF6PI9TrkbzkocBT5RGND5N+buTZad7FPl6hdBZ
hwsj8AMKZrTnkUfehci8OrFYh/y35ql/4J0KmLLHj/ZNDv3+odgqBFMmXLuWTyK3
ct2zKRmLHdg2/PIMmRxc1DEReJPdQDFCXyTsrkVrfikXMze2IooMlPzJnqr01/HT
buQXnFPyPesLVAeG7fTxLXepOc+ikwDYEHCTkCC4+EZaKLhF6HDJ7lpP9GDj4x1U
FyEi2T0IixBaUsjft5t3RRGsJUFVsP/hhiyxEeZb2N8tTO2n3XBS2GCq3B6g36Jb
pKSix8/LlQd0voru53f1gvz/FIRfwpysFaEGexRor9lcuSSAJjv75K6IsiTRJTXy
TTlQ9iI2lrMDSHlxdziqbPPFNe+BPwCVqjZauSwrgukg/+Cl5SFB0vDY4A3xbi0+
xamqrBF+uYlaX8/f4SOA0ZyR+GzThWGDb9mWT0liskilIUn+tEae2k2B41Y5XGVL
LJ/z9tishNRs67/xksq9QBDHwVCbuc3CUb3+VdqhaRgBFRMY7HrEvV5TDgHmtW5o
LOAXezAzk+r/xn2u6qp0wl/h6p8R246j4jgznamnqsk37qH290fBIsjLRlyJ4/4k
zWmxKDX0dAfGCQq7js39UMXF0rn7WVtBHIVM+atKmaUn/op94EPKSupGz7vZ2atO
bFOnj8a85PHbsrhdnhs+yi3ucz3hhomVtCwpJqTWJIZbyWxz53vWtV4z+TWlgGKH
TOsG1E6O/N9bGN7M8GE2MT0GtnM96SYy7JF9YinZghRSy0ty9cTttK2JQVBvp+pA
4ELdARJzYZzqRtxkFrXUo9MeUIOj0BOwmbPBmU8J6/+k2DDAczTrIASfmaKtAJAG
1CAEqXtJpTa9RCcwldnrUziQwgp+1JwDNP0wPdN1kBti2vXUsqxqhPNv41/LoMe0
VvZ4hg4YJWGakKsj6QE8N82Mou4hOq7AaHhUkzkC1SfCbCr0QoNrLrIt4bDokyLQ
O+gn5XoO4jdgTBppn944NafvXBNHJhHHdJLL9262iisiGUL3G8fEIocng/jIZ1hX
yrT/A9oNaOXO76z//Up2e6LeJ0Zs5ddWLFY3fPh7MWrufbFSzmmwlJYih3A86l2L
ZtW15rQFUV7eqkyfu3kyd7nXiZ7d4lQ0JZ3ndYb4nG/UCXfDD+hNeOfReYSODW+C
sxZGMk3a4VE/2AlifSy3kMdwfLnCRGH176d8+J4lvBAfOuI5U9Nngxpdn0LO7k5u
Fp0QMmSJxDOhjeqPGAwaeZ0yKEF2SUJtl6d9TMzyoE2ShjtKIF0bHo3p61OqqYpP
4iwNran/arXE193Y7b+jealDmN3yaYsruunPpVY9boVBZ7aQIEDd/tYbou+nmYfJ
GENaVOXrh+ddY29BJ9XbkOK7cBSiy8iVtZYKvxtEMJ+JpEsSgBcmSgelZSfdd8DL
/XxP6zNBVcbxz+4ZxJbVW8TM4JrX2dHsr0RgnfYmapqq/PTcqILTt2tuq19vP9p7
nSJP1UAobRrlap10MfoZZQbwVVMtwCwy9j6HsSn8I7rvGoPvfGRxUJls+qtYYylB
X0outwwRGDb3bWsAWqNW61n/vg8HYEVYe63yQxxn//xsqHrGRWBPqccuxbdq00h2
aJJvYPByAmxLqI4TIykeZCVWo5/nZsVFPBnfdE5NIuJtDy5UVcRa0N8UMrbzSJ+m
qL4FUZ2zdBuoOPvAAovHq0V0TH0TcbR59j6Ieq01RXeYJQzKolVokeuzb+IxPH7m
sj03z/xNXzoolMxFooB5q24gIp6Z0CQIRXW1as6yJYqlMpmQA+sO5to+JuH2ARc/
t34vZ7YAv4k7BAh624Zpi5PjclznQxfFb2z/2FeuSXh7SSyUKdYaPF20zCnfo5b1
mfM+RotYkxJ2WAgvGH33OnKqdEoANAlTiVyUqpPjnNIlVwwmoc6mtSoLYhAPEySu
SnAUiAhidwnRGd5egiWe3+Ay974ZUdCdtogVik6+78lMuAQV9XcXm3IgMeItf54b
jGjM8ci51N9NklMirdXTq5UIw+EJwvQFDxtnaIZMyxnL/dqJDWlHXaBcpJZxpvbV
P/o6A/+KTfv+mW9+4pOkuX8zi33fOtnTm5AtJHpNIUSKqFZFumLMr9XYXR9O8nLJ
rc1V4uPUOJPwsbbpcqY8CrsIGHH9rtpKzqiwJ1phL+nf1QpVue1x4VHp0eAdJ1BS
7B0QxopzKoHCwSE6OvctLbdyJfBamqnVLR1WxTsL0k4QhtC45jQv6hxIIjgSQTO5
WCTi7Ckwdf/f92cDnbwRBtT+Rsk8asJQvpFplNMcgdgjYAF4oM0J1a/L9mvEWnFz
0mn2mmDLDWgQdez3AQtSv8a+zDbKRxsdzDaxfB/gylimk9f/yYdpfsoJ8QuC55cD
9ITph83Ltysjt/DKhtNRqd7ayJ+X+O/3DgKqsITTJh7CAYVszwb4M/q9FoFBuJ9y
aoGhsld8i9JWy2CHIp2gjK91AGI74x9i9lArx5xUCMleRuasNe5DCS3L2i57WiZH
e3FCbtohqO8lkvFWWzkl0BaYMtfhVb14kT7gEC4k1Zy93Uu/tk+IL/WghthahrkX
MHNuJD+mE/PQJ23hZMXwiXbVvnzS9otHoVxn3W5Igdf9RSA4YeAoGJhe8p2GuV5I
Lhrn4ZGTYkvbtisuN7kDJMCC6oGNOUrygja1sdXtzgj6aJEclb/F/Xx/UdgxyOm/
DHOHMqKt3urfgAnDmkd4uGrLXMjg1LYa3q831MBpbXyXJzrUyT2xTWuEOf0FxBuv
RMfq18LBU9AwO+LieNMUlhBG1lTcVlP08qS7TWXh5sC28HyGJNMoLIbCOdxsLZME
rk/2/x/g831ZrThj9bQw+2pr1SuhJbzrNJ2vSuWIyOBd3MIkkZ81QBNiAe4bSG1u
sjyhOp87tOeZ5mZXwNyCg/cGhsRBItbPR8j/TlhYkiKJowMXJPWV2nc0rqC1BfZl
6qkJJ12Zdk2LhHZjuQkeBjg7cMKoiRJgamiDqXG62elvkHh+Vt6Y1vSe8F13Aqbp
w116xKPx0aEA33uDERBHDblh4WrJxIhDRswZ+FJL5NXHZIwU0jd5rt38ebyB6u20
QvpUANtzH5EHGrWZi5v1w9vl+RxrRLw2XHks+dWI2sOnxET5hvpHQIeWIyoAHG2q
whOmwBzlzC+isvb8XPFPwFA6aZWaQGuAiJ2TwQKrxCX2PRbkf7QDRJrXzRR5OjtM
fCMbmX/fPeZxJdZ2+TmeloUutoTkWzrxGsh0th/hIqYVCBb8Rakjgx4RBSmj0gNu
BI6jLMGkABReVyMdZmk6q0VcU40Pw+/hzu/5Z+iAhtxlw05oVirtfuwZEv2y3iS7
oxCmUN3i04A0+eO0iLKUNEhK+31RaKtj2/dbCYYHrqjFxuZNpBM10M8g/OxzIUdw
g3SIvaKzLiZ9212mtUwzU8Zx/hPjEAH8EZzlEXsHONrB67kqD+2hpVB0FMokPJL3
TzTpepBqfZuvqatBVE5E3X5oYZk/PIc40Zw731H7wcyLhqEDB8j/vhg43/I+lQAR
0LA8sUJHh8VER6uZUEl6zFFEwxYzaAb6RfsnCng+0dozx2Xnh36Io3s/SWscrD3L
+ZclRnGB8P8N6Z28tWcN9N+c1Z4zBC3YgQ2OUqbPKHGW3j7HSxK+VGHK0RwkNUvs
ZtdBgCvXK9B234SzlvwEtSURdpZZ92v13zckSu5f4ieRlpefl/PiNzodV60oGOc9
LI/zb8zB3X5ORxEY3+ZbmbtCVuUkiUhsijdzvaF4TaKDks5oqc1++OS+GpDxIPO6
Ias4GBIQ3IvVXupeNoQWmILTgNdr6MPQouDaQmm9CoNp8q/zsMC9pmAe23vImFkN
RBP1RaNVGJbge0k5XRh6WvVKMzK0xoCTuLrLC2QEMpXZ9SDcn7mSFdJq3LPE48KR
Qf56yJY9Su7Eb4C2dlGyLTL3qd01ARzDa86V9nzXlITeZSeuRmA6s+PSwmfSOfyk
OlyY3gByuTqZ28h6gBLSBwHGaxml0HdUbfjLkvpOZdg2Im+n2IyVYn2J1IKXF+94
lu5wscXRIpMASvPGZizx/WMvjmIwc+ZzJP1UENJ7NDp1nSo0lfFfgpUpvFQgQWVj
fdhO/yQVQRNUCGRbttOdOZvA26dhoY5RI7vOUN73RytTC8Ji/UF2xaCUgj/pRdOZ
+idkzBxParJTaxkK3zJ2d5VFA5FK+n0xg4AZJIbEN8g/ruhcbBegWO59bmfou0Xp
k63o8xKEZm3kzIew5NGsDKPeBTfHKKLOzbxx2H3w/kRHXb7C3MQ/9j06oOXFfb1T
+XRPPdlUNUVRSOIRyhviLiZpFtTT4HwF4ZvGpU65AD98MKfEHYGPc6DSTOhD2F4S
A4poLWP4ZJcG2buVf69aPq1G+dAHN5W7ZU4Dc5Eh2SJnAsfoR2iiNW6xnbeZln3r
bGpVwzFbeYSQ9Ov9139PBCBcofndwoEGCsrz9pOH5VWJ0mnYAuYYnfuRF0T41oz0
uhWCtFYKXCjLp8hgGHkpzfmbive7M9Vihf6auX3OyYQhWUYD/3mxHu7+4hYdrQoy
KXM8NykBNgmbd7vQfKUNJCsLH4V1kia865WNmsfmGW6ShBkH6VDnUAfzngkyAiji
n4Fyjx0AM3vc8qzpTX57HKTVg/Lib3ouMqjdIlcpSMxp4+OmR6/U1k755gKqrny4
t3pnSCm8OZrCDFukNJQkmjKRqZcvLcI1UCtXDPYjEtOS5nFi15epZ6z5Yhs/GADl
ctwpfNwtMp/eImhGO0qKhbTkPZlYziktA1S47aKySpwqHp9fm0YD0vGA/7LThTXS
HYxkQEjtdAwe/gdrTCOmddzZdoyH1PxqTDv4OQmz2lBr5r2QumxNA38EbYnZW+em
L5qnrlKNZosjAzLdHzUX9pEx4rLzbve1DMj0xpayobA4o1n3aFj11H1Uo42NTm7W
RI1Yk5BYN2vYeOOeiVM+qtjVt71rq9VrFbQ2ubS0+964P9Eyy+yGpkp5fVY65Zzt
zRka+L45cDG+BGWfI5XOWMURGIcB9ZMyLU9hCRxzkNGNmsMTwadYKD2fJfPLJEn8
BkIwEnjgFfYQxtZLmjTMMBZO2kUUhfAPLnYD043WxisR8ZmTPzzAvgU+B1AXaMDy
hInN93hKGxg0pmjHg8u2/uC2CCRmjdk5zoqT3738QYZVxK5QbVntuuqBUszVF5eM
71/OwaUp6BN0Ksg2XD1CmLLNVYMgFLddV76e+5KSTmef8Oa+jOp4Rh/BZapAU943
EgLZOpVpJo5mbea+g+eFv3wDR32G/y+ZsXx00+QlzsQvCMPuae54RrowSvfg/0f9
ZboZucMb0xiHiS/yfhCFM6tIJIjDDjoUHjjCyYOyzgtmKT9rupTLbKhqXRmliv/e
DTtHsnI/6eqiW6M+aZKvPH866H+kHfnYtnHIO4NtVqpaG6BT6zmaQF29ism3hX7X
SMd2DQLPcrSvkIFygiMIhBVJcD3NqZRXcY2dn9o557rw783h6K+mfcPKn62hPg6B
SS7FNFUve18QECD61o9ymo5W2xJaAPXv8geKVFj25UzHgtyiv7WEYkOubhQMZtL0
+14+T0bwithyyxFFDvPTOWG1k++ggTs/2pS+JYfu54VUrSuQWMyKpVatYjhwVNll
JxMVVsIlCnecX6E4zf5+5xBc49AbCdFIBT1a6KLjJuQ9UExf4UzclE2uKoyNiiHl
us8AfhA863CsAokSHqTFS1PgRDCnFlDyMShz67Jef2Zewdf+vRmgNB3Oyn5bu3Nu
ChiC7B47Z1TLY6QqtF4xe0+zwMgab1It8Oj/ieZVaHm9tzEHUiMcC7U8j753u8OC
gcqWGvFtT/7lbuuoseEwsq/5EUfZ37hBe37Xvc2+lQidFQVTxo7EaL4/0RMn5NiU
Rw1mxNsC731FKJ0993AkK+t+s1W1lqMDkQQuPf7WMtvG6lByuGVybzmxoe4dBBdB
sXkl1Tyn7wFXH4ykMbc+dvp6kZNRWzBUzhh4I7Gj42UfMmj1N3L4GskXSEV16FXL
M9k0xjjU8HaAIf80grewHAhf9I3bgREDaa0wZrOOeq/Vf7jS7VUTay52Pi1moi4W
86uW26mml6j6Uk/0jpXz9SK94HDsdjLlTmEXM59Edoa2N7h+LWE3y35GLAvvESiA
VufdKBzdVvOSEf5l9CwPaIo2bbygfOdSUp3/e+FYcOtS5LDTYkXnY/HXQt513Gr7
zxAPTOfD/brjX+hnp9fNjr26mNClVS3IHyH9Hxr/X3jpgjLF6SnhXcfSwrr6vjVC
MKyv95qS02Ct42KiuKrHVoD9L35gkqll0S2EquILhrSm/nA9pbhAR0OrsQbGNu6T
rXkvWfZCjt9iezp6laGkPGegTPJQsY9v9fWOPJVEewtKhsRBK2NN9Tz9a6KUj+ZV
XEkXm0w9Qu1D9K5LU0To5PR/finWnoLyTf4puNhrEXrj89dV5feeW6fc6tfir8wB
ITxYAviSlCjUYucurtLZ9Loctw6iZa1CZuNi1+tCRuO2H3DEQl5sMjW1Dgtdji4g
iK527wM0abGK3XQChGH6SkyWC+f/abqdxZgahT1K1FEb+1aJw29w2gFHKrHm59BX
1REpHzKbX56SF02stmdPP2S7sMT46OBfKSY2QHyI9gfIPUvn87LVZfXIc1cGOxk+
kklBR6D3NppNx6zX01SKxrzdFbM2QbW63x1uZZFlUB8xEmO3EUQzxBBCCRWQxB0/
e3Bqi/ehVDCDFznzOg8Y8goTcvn2fY13nZMdYfMH8SYujm8s8yLkO+elBtO15oiO
s0LKCnHR7jdVLquooQhxg6BAiwqPee3OtTGIC7yghWrKuN3X4LEaEKrKfIBqU4wf
DxL3h/uGPb4fUGbl0EdChE3CjXFrR5EXYtLOB0xP2HQ2KFVDcj/FoMnWVv4NCmKW
n2YkNnaBRxthbmOIldjYh3Gv9jVrzBDFfnjrXEx3KNIHCrSsbPkSuFz3WUcUl7ys
JeYDqOM42rQyRXnAx2zjagrXMg5lIOeESKwe7HRbn0EVtFml7wtNzx+6S9uY8hcs
K+ySjwflQHQqct0Dk6sRx6HPWcI1fyy/2LErZy2K7+Q3utvnd7gvkd+xxIsZzy9Z
I55n9mnjsaQzpQdjnQR1pBks2xYw5KXTZyYVFpu2dRMvQ80ys0taDajMalhDMlTK
7sQB8RNB7C2MVX+YcL3jvprdRo9b5XQV33wurgIR5e0ko7LVQXR2fG39NgbRQEOK
KVYKXYmoCV77qKmYkbkCntqGKtjsrQN1hQ7AGAkLBC3XtIA86K9viheLRJ5Jy9Yu
6xYAT+kiaLFOGiZ2seLWkWd2jlCauRITpVfUvFNDNmM2fUsuwOMuPWT2gtcnRDOg
hX0h/FmR+5yHfA1PTWb+2eF4HnRmFeiBSVh2ua3aFLKvGbkMpVof35cv25dBWpXi
/Y4JtQiKQ3mbnw2rKqp2FlqfZqUwBeSXZrzuCbFOEb7cjOnchFvfkn/DZqWn1bxV
7lTClvX3KuO6qpCyWKt+tuquk2RJmSyhQNSJBoqHeUGa02J4lq9XXmVHOkvfFZOs
FJtj5wj8iNYh7xx3Rn6BpTTtYUHxEr5iLCTH9bYTrUZn0VWLSaIBKO2LKm9xGt/1
z0baecMxYIZbKocfXXvQSWVSDTBr9lA0h4S1o2xJdIEDdPBuF2yofbPZIDsku7Yf
CiU/grWZNguf1nCGy8YQKmYUJTLfuyvnXR/7h330Yz2R16vffzFsyyFuwlS2dafX
FGyhxKB1j1E0Ki3SN7rfUrf21jGZOc7qimse/orfBeRUaggzc3gCEvSmVK7qsa4Q
Ig3jcQ3wA05jYqROHDW+A8baiubAxWzeSfogEkpnhpgp/G/hUMXDY0eEUjCB4ZHk
cBFmyFBJ0RVtcJQg+15qeRx4B6FE6KjFdyXdweHEDiULJTWB9P9MNlaIt4lO+5z5
5M2vavVsbNzVhkYkJIvFogKE7Yb4DSChggHM+MpstJv5KKEGkWo/iAnE7DYthvY2
qz1rFehOPHJQ81t2xB2KN8hL1SBFlOr+zeiQFrAY3vBC4oPGCZKsJnNXG0F1G4P6
2Dniv9+JgXX2wh9sXNVZYE/QN6NAVTBW25Jpkom1SSeP2hD/ubJIW2p6GKOgoktK
lnDmdTyXNu4VTy0zZ+Rd3kpkcPBIwCRbzC4jz4GwddKPNC2r5UNvaBhW6AaPJ2wd
YqZqKm7mfin5O7rBoab+eM/oiDRAKWoSLtkZJg6DYx3AYUZ2G7oYUUEOz2XrqtIS
SEqrOzEkmrtikLNtnSla0COl+sidZbIGv1zhcg/NgeT/XbdQoD7muOe6kWbodOId
hdkv06i2hfAOdkpcdv7+IwrwK+4/TzHeLllMgxWeNkAq7+C0uhLLGqsj/zbTfZXo
E5Z8La0UcytuVu9QCo/0tyP9v/aTUZxHFhFHdEEoSGpmeKysFFaBVpo4KYbvc7dn
TXoboDdO/n1r/bB4/3Y07ibsU+KLgm8D6InMO+1XFYwQhda8m/abRxPm8iNNsIHH
6B0q088G329XAL99u9t+NWTrGCigndd3AgovLDHXFr0ZCKbzMH1gQTf6PpHF+FFp
2674AYugRi6Y7jb7xHVwzGCpCSV7mCFdZ3DxO07oOZLQzx0sq2OF4WGftY5Lbiqq
NHw1DOs10OEaEwDHTLi8FcUmeuIEcZHWyhYO5LBNTu/m7B6hlWS1v3FdZTTEgl6C
VUqVox5D6Syj5Mh9AoVgm8Env5EuM8kkGbaoNLskKeujPZSPlghLlivqHT6inMJR
hslTI9SWuwLRFtTuCdUQdx5dJgl+ZJiXTtAX77ULkSKJHl2fOwGQoUpfMNALkejo
vZwvQ1j4ol6s+lamAywA50n7byY9y9tTNvAYOt06idJW1whwec/yhepCmG4NB8B7
NUd80lg9I9EqivmOBjPLWwU9aV9yKq25zJqbc5X5MCCLresHxUNrHd0B0j+2iK2W
rgM2lrgRJ6B2CJgASUzyiHTvd87lF0Mee0dZ3Rij/s9bXFvd/1D4PnOL0qNxSywM
ecNu07+jTSwTx4yuiSy3xj0r2Di+bN5PzhP5iYL/6iACtR0l+SmzAVW0ZNnOlF2r
Sa9Imqff4E5dwF8ZFwtbhz/ifSvbn85EFyumldP5qh05Ad/5Mmt3ennpmIgTaYHm
EF/MBhB/TzjRSml0WjjW2jB+oOGpr74M9Vm4F5+oBjeQhtXgQpWM2p1JxHjHO5bw
yTJRKSdJn5Dhwoz0nbIo4VMmAeUuwPUMGs567qzMhKvDdvL9RWFt9qcKxNxQZ2ZS
rsGAzZ4+j7Vw8XI46wlz7EF+3+nUASWw1Ot4hod0RplMc9LGsQkgsxAowe2ka3KF
z0HamyaS1gl8w0HuRzMAGdL0eobq0sm2s/UEFxyT2vs4D57HZnkZK3wV7bPmubv1
ftLGMLY6aIWXSRBvxb/AXEtQDn1+gkGQ56sZ5WOtxDHOTFMFoWmxBnwwywOKusAj
ZX6+axcDCUPQ48drCkaMS48Ac3tgZp410XY+I/Js7Lhgo7V+OWsTq4hzEvzpdAVg
jFGgIFYyHEB+o3AWyoTaMwciZR85pGm0rEyRvdzwV0ZrEIkLfCL6rwn8mN3b5ceb
dD3G0u09LkVz+FBYKcp4WkVSS7FRSvkOvjhdpk3Ah5iOAu1I0/wsCmyiG7LMvdvc
CC9aiWXAXk/766xTKAD3qFudTtgyvT8qeaEFCOFSLpWVLPwW13l+aeUuECoN1NrO
L/Jvj9oFpBQ7PWlrti38etkLRCqyQYDNOY/f/a0724+PhfHxbmX5yvI6K6CVasYS
7sb0ENGo/1RpqpvsTRRvwb5g4pInp7VL1LH/3+XOzJSE/SK9YyoHasSYAJedRQMK
PYg098Q/1Y3efq67ZJrRrMLqoZnBxV2f0JxMVEXwxNPZkNOyUrvgFFgoijX1Mr3b
Af5wQJQozvAhN3qF37ZeREGq3VP8BnFjypDJ2FbYZK4eBk5/hXHwSF0/KU5DZcYR
vugFXZgoiAgJerSvAdUlYxM5g8TMKwBhCLRNIG9b+8kCbSzOQx68R3ERVGrkJ2j5
b3ombGMugqxz1mGxPkxqITJlkih6cZVHESuAfYOLsc+dnEFoUznkOs3jOQx+E+aH
2Fq43gY8OCVlmofM53STg0jX7QeMChb8wrjnvYvGIXtXPyy3Pg3rNVCtOggGOMJO
PmC7/WyuZPg7OqQ2u9oAW4aOdvYh3Cn7bnwj7tEu5eBuXdDdVNNgYsSYuXp9MWOR
aJeXStpcDYLtZih3xqF2tyIW831xzU+V4bD1nYthbL3KFb78zRyQipGSNHKziobP
PsxRN5e7T8xwba2ib43p+WH+C57ExBYukDuOmXH4J9aRg1e5cWbFLpd4DQ3rSyWC
JNHlrT+3+IaksawaDo7cB3bFRvBV5C8ckHuB6o0zPHa6eq81y2stSOZ0zBh9TBmZ
QO1dP35LEd9LhyxWxZQQcwXyt5nnhmMx/fFduzd/HdCMGbUqijjFdxui9Jkrxxf+
usfk7TBX8LhhAOOZG3Kf/k4yjZVWpdxMeSozl25uGTQqFrw5izusikO/rvhxURHN
V4qUfcUe9dDqQzuc8DgiOKulCewggPU5MBR0efirxIYwcMTJ/UvYUuaerpWNlQdc
Vh17ruNP4rewxR5LcAC0wHy68mFH6BayY2Ld6V1KM4dKsNLHKHwkSpohmJdVJdDo
Ghfze0dILPF2n8BD2eCftrdE6H3l5k509hf5wbMuM3YNtbK4KukIj5TfzgfS8gPA
eLARmUyjtO2WKSMVO7V4CfggMgmtlCEkZ49O2sI3TnmoQcoYuFOWOIQnywpvSiDn
ew+9iiQXASNNjrhnyntxeFeIyYPfh3Es6ps8aoj7UuVE77zVRN8jq4wV1i9vZ4jE
d63urcl9UBYT3w0MODDygNHAJBFNCzfjyaDTfCWv1n/9x09msHhXfvqVsK4I7FaL
v+Y21zJZZW4lIKW9sRDzJj2b50OzpYNpIhGf7wOScnCxXN8u/5Q7IYBQEXxn5NWk
A9lYqW3TOA+JiqAg7vN9Ya7xhU5US1iss3Mf9LW7ggCVn+JwTbIctFqQZ3xM2BTm
7SfG0xnVzubvZWCWlN8eHKAFWs8QP23arlJcP00Owmg2jE58tq4IkWjA5F9XUlsD
pB03hgkaNHj8ToB5XY94nhLLGoDcVl3oD6Atftn2RBix1HVpTcFJomSd1UbG0xvl
wgN/nDkluw38NxXFLhW3eomgvTq3Nwe0ETjYNcmx2FI2SKVqPcxth+xWqc8KJJ8U
SyP3PBW3PN3vew3EdGL+RfEvx3YQXZuNutyPl+E2tHdgn7jqsYYOLmBEYLJx0MpH
uMU/Z+1X7RKyvS6PEfsQeJVTGM+MR2Gmx1O6d1RjVMAC+f8hih+bzC/nbY3HwM6a
L3k22sHOosut1nUYjxigZR32sE3OBoqzAdbAed7RrbiizckNDYEOk5lMhXavYrlI
67ChTKdZzw+HhPg+1GIS6WM06v1wJOiSIylShCvBhRcMbbpVTcP4mGKTvvHNhvR2
qGIkhYwOi4W4lDLopj2LWLaBphLsekTpM9MX331TcITApVfnZOpOzoCApKoCH9dO
OfYEJgV3fzj/+4xOneK3PRD3WGSclLdDWW1qcRxoA4RZogVJp2AUV9NrWzfi4IKN
24XU1giAA047R3ERUzmspLcok+U0jRlbH4JK6CMi4fz3iMtceK2Sya4Ij/Q8p2oc
Qfpe0G+Jjb+6Paei8Mz4TzU4dTI+GIHxNmsRpbUqF2ro15sy5FI8WTnaUe2Ez+dW
36knFPmXgnERMHI4VBO5N0YTyCLncUG672hgWF29Lgd1fxXhIJxEDntm/Mr7ZZgL
IhV+HPAReS1TwBLlL978tnQ+hLiX610PbRk36YUsV5FZLk3mXLNYkpp35baOe9Jh
xzdoKIx08ltGIoy1xFnAkHaw16hz+3o1SdUGfuHqUDH+W4jhyKpa+owrvrI60Ugc
oU163Ec76FHJ70r5R7/+9cdY0EvgxIhI1MBMYqa3H0ZqDuqHnQ09za7js4W4+rCz
I2XeHQa5z8B5dm6wOTk7TndAjZb2tA7W5ISaY5uPK6mWpV8oIfOyrQ6v4Zrxc1qk
VqBzqc7FQ527wS3YhSfLjyvf6x1kkniAmDL8e8A9EOxLGanUfA112yYO0TKk6GiX
To585h7/KtGsvWc3Auca14PXVWijhlwvR5AFqTR5GM24Q/FTUFKDjRBMP9EaF5EJ
TJsOr4OHlbJ8ryTqbV1BCBD9IT41j6Vzpz9DTAofXoZJE2ryTVaObq8cqgguKMGZ
BRBuRaOQ20MOXvtpiAI1ASMt4tENZ3zbZ6nTDk0ejvOAIjopHx+FAeFDVpE3ifGk
nLBONk4kzFnku3YMLafhf/7W+EArmtgtK30/SWrL4IRjLKteBBampPOyWPM6xgM6
V7r90G+ZCaUX3FRQVrluYgNADoCcIKjKC5YACnbAAsRGH8MeBAfyEPExgc41Yl8Y
rT+o9tGUD76rf6vO931BD/LAVVkzCtIhfuAh2qoa1wIIei18zp0/dfjDmNcMiSZu
msZwgL6yq1PTieaV4cqQBCcCnA23FfrUYN+4K4CCi7qUUWToov+ue5P+iagLo8Eg
J7OYDT+COgUCpQ8gWWnuVtTbks47032IwfbcsmIpWwTVDV6PTpnkGdZErbtUY1Xk
11BOHrf8hibKJ1dUkNNykv0PrcZD95pyp4eSKUzKEqJd09pdOiTl+LVsN54Vo8i2
zMsqTCX+NnSy0FrGQfhl3aV1cO63ugt6xS907pqGWmJij1w/t9a7GFFtg8qbxKQw
g4O7X+mz5+H7WWfh2MAhpJcuQviO2LgmbLtwIOV+6Me/hzSwdT9og9hkSfdEzsCI
2/yOxA2XTrUbi6d+Mi5roQnklFpj/om8FX38yDwSotAen2S3bsN+O5ig3bF4eCym
LXQQOLnk+p+khotvThlr56x/JCKv5TYmJbyzSwRdL3RLhpsxjL66Wqeynl7N++nu
tfumhLp4tmj1/RyTzikePVmPv58sm4cxcIvcmapPgX3+7whJHP/t0BKGC/BTR/ks
82uQDFKPm8YC7ObE5yKPep6gumNfpxj3Y2JCjgrCzpq/Gi6i1e7zcaYAi8viiqVx
u1U1R5ezKjeJgJKki+vLHlCjNsTbds7owmfKajjvoOmhnvynub88o6MarPWq7i/S
TbzDzIHjEUXYVIlghOyoQEWZ6cywwnOZWdR9YCCheqDE35DnVLBfrydUIonYfC5E
lSsN8SjTraHn+yUg3XzzNzUPTjHgtHjcUXLF8jAmdsqhOcuktO7MSIXDOhQrjlTF
ZYom/p8I9fnsO9EhwGJuKpZY+O2LuGk4V9cWoYl8EKfYdI+tC7pWZmOUqIUzDXMn
n6s5HkEMOUzdGo4Lf5IZhdKeNGmC966DXBXUwN1qHalweTWuTBLz4Q/j/zgfWFUj
XmbI50LA7wxdDLH0ddjo5H3D9VBprHw5pyH9hdTcX/za+phEDsOOOW1Sj/u0p/4D
VPsIUa/GoGmjcJtARNyY8uM7ISfcdtN3150xcfe3cj6TCLJtbtUxBksBX9R9l0Xm
rvThbOjcNv+p+lIIm0JihrNfiHTc043u+8uwqD8KaB7TnGj4all05ZU9ccL4QcHj
YIxF6EMJxLyajG77Ug6F8plzCOr0dOcxAKlL4Zq46UU4tvn2RMNEQg2YWuSm7bFT
QAxdAONhTAF2IeIpxwdDEDXr2R6BHDdb0Vb4PUxdeSYinZjspIAX/GjJ1lfWiFK4
c6uR6FapHQYhoZ9EvYcofJ2zzSi6rc86MTIgep5AAKEES0Q3N7vGfDwAYL15AifM
QZMzdT4kTfxduqe6hn8pUvu9YckO2H81kaRTubSHOqiYKPivSuvBqiEszDzu3dh1
UKFzDnAbe9p7CvHZj5pgyQl5hRhpEd6LluHaQBVaP8tA3Gzy1VQcDRtFimFfi8My
kUZNlfx3RaNsCiq00TNYrvcePfnpPC3LwQvxAUZTrbgrb6Xak970tsbARw/v3DSG
adsnTPJ2f+YrJzjnpa2PkqCmMK434iwdKCvsclQya8T8DblWH9rkHecw2YRQubzb
soC5ixJdtTFiOvxVONa9D4U+1udGvKjV+Uk1bV3XC2FyCm+khzb8DJxx8ZNclyUe
uVUw3wyOlILoqsIa8PQNsgdFVEx+NcFmumRJo40Lrg0kNKSOgc5m8R254yeGoLo0
fQcbq7Vvg6hFvRabp0OjFAyuK2SjJhikGPa5MYQGHfnrT0pczn8OaD6OZNr66fX0
oWJd9amJ8YM/yLo6ASAu1iEOTiUxbfJQ1S7IfDddsxBeG28TbDwEAMqoTQGvVbb6
4tvMnIGdud25bKz0SBIFfkRDLehUK6renrK6NWoidctneVftsodJB8r9ZOB0B/CL
C9Mso7c3Ko24es9YZQ9idPbeyRcosj1zgFDLj58vqJX9h4B7NR+Y5XqtWJG8qego
3VceCXcfgjtZPHj7E61965fvvSsUiS1xHGJ8+RT2TaV5Jy+nTgTvCMk4hNEq/2Nn
DzFaxFgp7C64AVLDUrbc9VhXuz+qlpFDqClCQh2eYr0mlbYwnqe9j0dkj/6M89EX
z/AMPXyotxSJvTnMkFH4BFjBdXZAnofKS04S/Ycp0NvM+83CI2as4oZ2rI/grWat
UyC/xog1EA2ZuBo2Vk/y5oVcRQhGr7wPfklcBXDg9BBO5KEviJ2ENGKJdsDKGkCP
DXfPJlEgciSO7DXpSA7OqnZ9tski+FGerFBQm5jidxsUgmKHTsgCvN92qPJjuR+B
kxTKjef3VHTOoqmC88smrdT1u8gQDdwZfpWvH2AwiI2cz+Onj4gZFlAGnMmzl9Xa
bLr9WpUaY5qdvKyRnw9kyq/vodslhn4rLNNBr4/WdIIoc8y6vD7ZEtFYF6GTHdzp
i7Es0J0GlNDodLDocqhzsSBJPHU9HcE3L1tIgMOUBYLP1+M5qZPOJVaFk2OSgfS0
99tmJeMhaFd69jKrDGvVnb6FEsyUeTbSv6FGaCPcQACI8DmqSpIQmgiqXSSs6Khk
Nhrhdb7BvcWEknJebWiqHXLDBnoF3jxm6/LxWqpytx5Y9JmaHBTrDLnml7TJ+pxS
jqPba1IJE4tKiIZ+45wI4AOP79OfFT3YOP3Z/H2I+3lHC95rZhIF5gtr4fUmllL3
vWkzsG4vUYIzXTZ0QY13i6jNQUphhSMgOAjJjnRHgmMC/jOOvqWXlUq0WP6LDdSf
ek+0Iox160SgySj+tP61VvuAculRvR4NgFkkFvreNff1k9nKZSVopnxmF8EkvaOl
4vbC/EO6ElXXA1R3oT05CM2hSG9fm8B0C9MBCJXW6C6UR9UyAE8qPUFmQoblcaDT
QVkC3C9eAxvW08CMx2VVMHEiFGABID4knKLc5EEnWZjv0360EOuXvJpyP6Xu3uJM
Tupruo7zPAATf8jwMSz/YTCMByd5j852prYldW5ujLLBHDHrp5dYco8BTsjd64sY
OlIai3abyIyiSoPfHK5a/SipBBGwwal5LlJFksIxcNx1/nZIE3vwNXrZ4Mb0jUrz
W4oxY84dciSgaIQ83sQ60Yd0Jt2cJnjhKsaMAhLlr3zhkXiO87lmVIJ0YGJJNitv
PvFtPz8cHu9KbaJp/IXWRj0mZQ1uT6LhrOjmioDaOs7fQfOyxHJUYCCabU69haHR
rTxn5/aN0FyrIlE3X31bBCqEv4aCOmwOPBOhNg5l7zTfG85/KjVim/AtUkdU5WDa
fafpuDT/9w+Xwiona3EMANUc8LVR2SiQRI4DwUapjVVssiEbBmdDNtI/B7FlPpvm
mEhqEFURVVlJ8Aze5lqTW4plwIsA18h1LyBJFUfIvygD8f3v1rNwbUTI6mE6Oqi4
Zw4uDXMAaGj0TfOH9oU3ktKosIyRTpxvJezlbwRRCMHLeJah6QezkNQLvIRezB22
td3dV4QF7uwRD+aaONNIrUhGgPg/uKjHU3AT3StQpDgwoKgJUMsg/7L/ZbPcr8gS
94iO+Y1Ta8Ka3udwWE3a6kwTjAOEEnw/IlXnqVXE0ImgYXnd3S9wUngl3rV5iypS
kJe5AlUrJiANMbSQMggbmfKHCLSM3wHv0ffw6IgjyRHr9qCiiYcRDAw2CnS907MG
y0im9qUu/LQdjvbsJY2eQTumc1n+JMD7woGgn1YErb75Hwk6XyP8mNCbqNUOwAiP
tR0zDSuE7yhn0bYZ4qnBaUBnnsCKjznybZpfEgEsX6gBCyhLTgUbpcEX1Hmj2zRX
WV74LFt6eVE6OYlBj8w7ckGP3dWVX/RjI/K9LS/x9yJ2lkjqY9w3x5wqPEqQjM+7
0ZDzI9rqNeDIf/ahC/TbIWmVaNcNZqbcqBBCYpLQaZpI5Wa5d6ll93r7MJRh425c
GvW830Dbfkr/6aVQCSpfZOV9TLqddWpbGubTWfYDQxiPpQ1P7HGoIuxlAvq3Tj+Q
zfSfvGaBXWGLAfuyxmebw/S8QIY9hHGMIy7BA2j5R24rc7S/UOLtiPfoSCVqHY38
7lXTVN19MuS52ZxqXqn9JJ7gxkVKvPZRGBOYLlK1CM42wUmR1LXrsBB0hhghW+Mf
ACCiWWpa+RuGzLYOqwEe2kgsQ2OTwOhT12bNTlCj14w+qXRT3GXL0127VSTWfw/z
IbYMupX8U7wiGRpI2phR51X37vsrYmDtn9BWGC83bUhbxDNr1ID5nzDItFCGDMyb
3NKmu88zMWNtQyBenKB80LnN5k9yGZH8HUY8KqMN6INbqmk/EhODISQ/aaMHQDH7
Zhq6WvBLnlVClvx64C05mu0u8lT89vdNCrbtdps6R/XF7hud/+r4Vm1zylhpUsO7
9cvEUSDZpvKj08Egs/h2sNDEIWFoZzI4/QnRjjb+l0xjhCtNzYrSDjazZLpSaL28
JKKuzHINwLNg0qxg4XuYKqLL10FvJ/Hc6Xixeo7+tR5whvc8uK0bmlBW1xu9adMR
ich8IYoZolcH0MIkArfvY9u28sEfw9Oz+gnCTTdX5Aoz1B5k5m8EkSCUPSqAemxa
SgawyK8CVRG4f5MS/HIgq+r4oso03EZa2nLuxDkHVw3bZ+gUI2rO2RKr+fLCB8Jj
tmHSufkQL0bFOOUTM5F54pL/1w9eKPbWziN2KWWBXScrsy5xTwiSRjsl5t8MLiYl
74Vtyl/uVxs4DvVHGs0LWCLPGd8jJqXFbOSF+mG+JFPiieAFsYfcvzgebAgKuZBV
L5dEt9zkDzAjPbHw3orEfE2yGmbCLXMTroiQ5n0V+2MJGM9QeBEXciHnccEhOiO1
3f6kAjQ0POf3PhVeZBm+K6hAFFP8d7gqtusZkUfKC0WEYalSsvG6/hDczxwJ8z7J
RMwmdwprgKKsti3PUHXlENYK8bi/sVmfzXAxL22sbgXUxL+q85nlHJuUDB1nphwB
/1Y06w6E2d0ocvGuxyayXttNm3cU8iRJPqAmtBPAh4uwOC0+MedvU1KgW0MQDuoJ
dw3/2IEuVPp95xrBxffXiRS6CeL0ktC8GnyJMaqeXxeFx9LpijGGUqDutNja2Syp
+Qn1yg+ERtTbQ7w37l1q3btjqep3wbNw5j37ZyA806AY7FCKMT9uSyrbflhWfwrS
S5X+h9Dt3pMfiN03ZziU6lbIITGGLtj7OMKsggXcYT7c9/YFCgxV6UW0EKqW6qdj
dnFofpT3IYPdbQ8o0gc95iCaiTjLLcT2yg1mwnlR8Z9hwFTJ7IgW0jE1OqPwBr0X
qTWJtM2b7HmfPHFVnFRfhbtaQe8G3w+iU2Ioo8Mkmq34IokBR3tR6HqPGnPPbGhz
ElnXN83xLYLIS3hRmRmLK0PugVUIFzs0mOrzuxjiYEPrmnbQE3PaTD4kZmVBn8th
/pbWegSQsgUGWZv6HDbN2VQx+KzweyLqDJYvinL/4gKg6YOIVIaPd9IPiIE0HLgM
4rQi6U6MkpIsFpc2vlo2iuy1m7srg+OCK9G4yILBDWw+c/hLzcEvedm5v5Uq4fxV
Teybk9aBwAz8HE2UB41B21th+6jmf0QL/jBqItxswtqR+eK9i2BHTOxZ6z6Q6hpi
r1e2Udy4lT6QhOlgO2qjFo7yknEin1jeK+L28mzCF/OPkdLgeXBRZzN52bLZtcdB
qbhQWVwS2uKcAJkU6m/MQj6k0VrN6+mUMZpsjV4qOYIkholIMfS5+e2k6/8g+Zo9
JSi4HuNx0sWC+CD2fOW046eFPX2Z/Fljh77mYznijTCwd6KIsgT3gC/Mzuui/R3P
yDmpuYx0c6oRQsU0+Tc4XNw6HlyfTrUfc4/FQtqvXuSXNBh2jrTVBonkitFm6baE
AhzMjPjO0G8CGZbJ1+y4GJ6/RGx2Qic5yjENC+qircdUW5F137I4MLefneigWeBY
+4exAYmyjknnLLa7iBGxzpOWvi5g6znckdrMJ5dK6jmFc2+mp6zpajgv2I78URBY
UCLHdEXX/U3+jVskdeUsveEJnDqTcfAP7Bn/E7g5L3UyUzPqmeTGw8bHBYu92Kvu
BLJDDHGdhaKM1BH8jRIIQfn1YLBePeK2deoMm+ajxxb/zL81//SArUUqRieE58oN
bMjFu5/2JEZAxXEKKTAZAe7ujFgstTGFs0Xpjik73E+DCxrYSFGnJrGusmiZdLB/
Ks1PUfHxu/39PARdaiDx5bpKfC9lgmc0+Mxi2wZekhrLRws5lnud4oSXB1SIKTrY
ve0gpNyICUIa6VWESwzZnp0dnqZlRPrlwUR2gAwL7AH8nC1fsSPF5lyGwgGAKt0x
RPizSGM5s6YONNcArf6p8Mb9rpYe0aoc3AYYwtBSJjKTUmMg/h7myj1SViFvaVQj
2onzYyfngKOfLPdleqaFjVkX7T04LwZB8hCJf/LV9KY496HX0lGLwxIOyuq7WbmX
7n975JntNa5NpkMlKK8JxO15rfZsrccIkkI9NJx3SFWTonD+PbUMTB7193XyisAu
2Vd9kl2r0TbSGRFg1Ay0RVQ09sBCsopPiLygDScy4IOXyQgRhTbLRKhz52R6d/2E
SEuxicRvdVc9QoETrCD6NsT3g2Vk6IfZviShEE4I5KcR7+4x1Z8OWUro7JZekmuY
tJP1Opec/Wa9LtOLniRLLuS556jDj3pbnpuVQ9FTBNf0YWXbB17Y3559ClfnjOy+
H8Qq58zPNCKAID1R8Ixn++6T7a08ZqhTcM0qsx7YU+bQtrSEWoC60S5W4tdD0bn9
YUopY5SZcbQVMTDcPoSHIHATvZRsxu/0qsrUxeGeFhQFfJKPciFnFDtNhfM6IlhU
FQEqV8mSXeqby2zZQviFWDiUoi+YlJcRh8Z08y2vl9vRomTFTOvYfdt5gB4Opx4Y
GnLC0uBJrB7mJNplkANGyULQo1u1N0z1vrXq5chVGym9h6Cb/9NvrHRhj1hP8TM2
Dc+j+386ABYUAzEIAlHRkt3sGqUGADL0gbfUIns9WY8t94ujGsVvu6zMCj8eiNaA
kNDHsejOAIS85IwDewlF/eCEoUANxQEECLDqfVeTmZM0xeZXxsIgnz6rd8rV26tF
cWeunmamt5XpBth307FLAQ/lsw7BxPmK5gcaL+xwJgVqKJYfRIVBVM/BWJcMopd2
js5UaDdcTUxc3hV3iFgNHy8IJEp/8rvW077USMdoHx5Qs2/rLsC4KeJnrnPamaWR
AvF4j27PnaoEloDceQncR/boQ6MDckCSeFEWPr9eWw1DyeuLVPpMalUUp/0PoiSh
zLhpNx7GUrFwpVIkEHGBhdUJuqQB6Kl+gx74K5AllB1Gh7l7gC5rUlLs4NYOsDuk
bSILF427tKY4vMqwy9ncUhN3xwqLtFOtkKK0sV5v02XENpsLkNfIpWq996a1Br60
U7jnD7XNsTU61hb5nMWGwPc+ls6lq7jgE8h1Vqr7dJ0LGp+XvZWDU1GYicDOASN8
zUXKhFhgjmsO99Aa6OV4V0P0vaoTWV+dz7gX2PL1G0G1b5oBcl/cd/FP06KQvEO2
wlDeo9+bjHPz58K2wy1rZj3SSmeAUI83T5Ve5eTCbIqVAcEDJII2hpM08GVih14k
hzY3oPPKlqomAFjS/uoJB0Lf7SHw+2z2//lgLPSpMH9Aci1JSkhP0J2FimFWbNP/
2uKio7rf0Hh3auU0kbp9W4N8QWrBDLCzNdAOFjlph5kOqlbZe0nZEfOVUgymV+Ck
E0B0q9fG9fR30AGjyMzUf2rWkR/7VpCnk6tL5DiibRXX8NzRMJ2vQvJRDADuqHFH
2eS1MdQcBuf+kiChf3GWFeBQSlhx1jz5MIZyyozzsIpDMgtPQE7WUIJzpJO1JL7I
COPlP7GCtUSRok2f5SpsY+6vhhg6MAFyS2T/kUwhdLTn+isn1XAp5vV4v0nuveoc
Op5KkgZvqxbXg8UHr/H7lLBJRNTr5Vhxea3VpW9tzfsxF0LLBS6O0qFTO1zLAz6Y
wCEnV5ksdZhZbXJFwarhBzVNZJwdCUuUbghVlP69M27orfOFVJdyucvuAxzNrn25
xd+zuWPpOujHZypU+1mDm6qylXD2TOcpnKEDXTZXOeDJPNAngQQLUlNKIQ/zVgfT
xbUR1xYsxnhfqVilWcKnY368J1hi+lnuq/7uVlIcS25cBsS2MPlG2Plp34BhzZyP
wabe31bhGrefszygrZ82V+K8PYQbd9G5ZrMC0cJ3CzvOeDRazZq6JpbWYXBQ69zd
P2rSSgOV1oX8d/EuIFh/3iDAHmNFqoD40KhKQ6T7oWzZlPq7HF+UaFTG140NoZ+M
PuCDXzii3l/h+17vHIzUHqsAfHeG3oHa0lj0ahY8yLMXWsHpPSXSMpRoHNmrvgwV
yG+TD+76xK6lXobIzk7kRsm694Lb2GWXd+aT5ABJRkz05Vdcdprr534nuu7+Kh+B
023d+O+lVwUBijxYnYGQMhGe0PSWd3mKEC+T/sxE4AVRgaS8MRPdHkPq6Vri6RWl
yh23d3J6dnn7n2isvgswnMRbXzjjtYXVoOk/iP1pqshSaYHWKUUFzNnCCxxN0Zqf
BCy6EvIJWW6oJ+QrdaFtH1g7VqLHIWPVSbLlVa2vZq0dLAnwSk20Pb04+ya4n58H
uefFe7ol/+LxhWw/x9oFOjZGGWULi4hfdEp615fmW0aUEUSVOh+/9aESYaXXBmSP
/KLRzzTMadKFnFRvYJE2RqkZqbvpYxOqtPhxCpxM2Xginv37UYLPu6o8lE8DWLyd
xi21PQEtkWVA4m5+BQqaeYKG4qosi97fE8xuR+jNQF74K/KS92Lkqga+Jo0revv1
ly9/2yxeGyqG501SyBLYx1jFxTF2WUSbFGtyou7eLTUj+f05KDH3ASxt/SQSVEx/
sF9Wl/ityxSjxkHog2uY0Yl+0wCieX4XnKd4jcz1mZlnSZz47nu0L+4pxGp4uvpR
2efJkLxaqQpgwC4rUmfbu1b2O8nyoHcGX1KVV87YLB5Pi7/JtKdsvzxAnIxnL0iK
tTnL6jA8XsktEbYLOtZNkOy+gk/jMlX+6CzKcoaokv9+ULHzUhvLq8R4tDZcvDjQ
7uORzvJamazvQVjRl2UyOXWrb30So3MQp5qdOVz24aHw1MnDJogD29yYS/D3OYST
aXD5m+sT17au2/Apw53pipa/LHGTjIzrzVOcLy4QeGnfRwy3RaGXDGk2sobidJLw
+zFI1FD4I1oldSqcbXFNAZ7Y3jh85W1Lqw6mAWGX+lyvmwpXvdAAGe6YkDdpp7U0
WSSeKMqrJYMV8qpHkV3lGV/jdma2cxVKSD2uD3oU/tPrfP9ZCOqreyNU00hLT8qI
GPKOsIO31b9zl82cdvVUHJBTwne0JGz3Ic1Y+++nqLMNVHHrRDB3MGlK0NW02Goo
RirgfPG0br9D7DKhdT2V3yisFq7mV+UF9ySFV1z3iaolPw/Y/GOVb5latJmwJDAJ
paYgk+8dyHluyfdBCXlAqwaveuY0CHCoJ48uRmqxo02RLPfH/EGFa0YF4lpbEFq7
7JtjB9r3tGsLWtLyiSWWF6Eoy4fHcrR19YBooVUPsKeHiYzMEeM6XlTgXzP+UQ4C
qUOuIolkRWfy2wQfLYMXNCSxqL9A9iOXmOMy4IwZoTxUPkkvo5N/YmzvcT/emO0D
Xi+tYOCOV+g2RRF0xlkbBQeQhLdrVkcjyPT14HvRo2VT/LXiHCOqhoripeEkPc3g
rf0ACwwhZTKatAaKyIK4vGeBC7LEn0EdZh9m+foex8qWLOnAkR4vgbKqxPfEcFTl
sLE+oMrVmeoPf0t4HDeMKGCw5G6Cg7wjpJKv8M0ysoLw+nvBH8wRhypvNnYeIW91
0tlB56BwF23ms4ahq7/iiGgy6okH7TYwzrb7scdBSrjclPOfTfdvA8sJ+uyXVCfk
em0m2jVN55R+8GUut2uZO1G73T20rU67VU67mFQtb6CPa8H79gCeGhQbf6T5N2zD
k8qgN+8NMwb/rseWFXNRA7NVElaz7DQnAXNHJXOZ8/+/XoF7rwQAOeKjEIwdVfl0
xx7r61OLysGvC5u1XQl9A0nS4bMCYi9VYnPewDe7nbirMTc01tfjH2LJIiffQmgr
V2F0dmYQruAVErYiYjLAJ4tL4XHaaMlKST07Nh9K2I6egKkQfY3hCWIB9bXR1zkk
jZNSkSbM37Ls4cugdmyuVQ7ouRf6ALw68f4rdIxulSRSlogSfMhujl9YRCPcc2JJ
FUqCv2CMr4znWJPH7uzliRtoCPnBDoAFzGyJZ+dESuMAGiKabWIZnb3g+1e8vy9V
wi63zDPbFJhDbJovGU8rSxnodY53pDiBE1MwIca/cniPl6zJeO2BRcgnWuu6G8ha
gDBek2Iy2ers4TtZZWxYE3RG1lzru4MmOrSazNx0NqYTwW66JRoDCAqnJPgHQrrl
Oj3Jm0C5n8ZFsnpampiViUB+VHKho7JR1DsmCZDvS7Wnyrl5cs+a9AWJso6tmWNN
xW7bQqg5SYXKwGDRm9vaUl7Ym3FzshnXsKADhfL8VY6bQ8tAwQSI1tzC6tcLaUHt
jK0Ypyxf15986M8Q4N+of8+ceTWbKeQ6WtdnYA9qRuCySURkTj1BIPugXk+9goYp
Pe65J4T4nrss3hBxMmMgqIFi/3HiJmdHDCzLqkQGoaM2YA2ZYAo0u2AUckbJslln
JdkzwGfr9A/giRyn+99r+iBr2nRmu+aRislgB1FOlNVpxurNUCS6EKsmKr+rCyE0
SWbTeqwQoiW6luhHjtivODeYSxGSEthqlMRs41emO2c02/UWhE7Zw4QYLkq6azUG
35NtbjNM/muYZ0w3+WSyQeWyX4tczmtenSTT3S2lGv9/dgzX2WYnqaUyyaw3VttC
8lKmhompkcreQXUvEvlPqgqW+yg/ptNEKpE5hSZkiDJN3N5VKsvV/o5wrJtDTnYi
7bm2TXboliXatzyXrdYxpHHlzoJXRkeQunPNm71BRmZgafjUjKlcgYfreJ8Eb7wx
6EOqBf9YE+BQLlc33iVWXnTyDepwWKcHBBDYi5LX1xOGVaoXHUjwGuNmnL8v/TkR
aCVuXnpYHmE9rtg7pqvQ2WHrEc4Ge1e8EImLqM361lNzF78Zn+a74uJktLdf2jQW
U/kptctBdiBYdF92B1Kp5GkNsTgglfQdZTKQPbCkeYC7mNUqJv5Vt1SlgWEXhhAb
Ngpnvsd1Q0HNFoWxBLyozolGRCknQdiSGQdc9mLHHUMDzR5njTo9fQsrc0SwSh0z
IWPa0aIe19o0La1S6jRRWrHWkVq8ArTU2Escd3i86ki4tpr1SKJfrLofitRtpaa4
sipADSdheb/pGCZTdhfPMgUYOyi1eZ+I+VZ2Cwc7nhQQdn//m2LY50CZ5pnxqKUk
CgeUEQJts8HThm2OXN+XG/VlhWVWiHT9FZrPGtWzstMbVp56lrf1m4GfJ4F6YamF
mvmjsweu1F+GVg3X5N/P/3IuaXJk0AwgzeKu19gcUytRobImhNDyY1ijAPELE1KJ
WKcfn86ihcGBkV68tcJPByvzHzDNs7MqMrrGFHfwe4u64+Hn6IP/GoMkReR6ZHAI
kGlTDkjvvyGwRMzJDR/b4POr+8HAbnm6jQx/YZ/HdLdbfr2pPzsh1stOkQtHcJcL
iAl/oQynW11r1dY90Na7cHLTY0E57p7TRJB74ALwIHszd1ou7MVRMCZPQBwTPTLk
gyJ6HYBRm35GZnz2+DzPfG+MQQjuEklwSquBZFQAzLSvBMACRkX3fw6DkEoB3vwY
8+Jcuo6Y/b8sXMHX/gHucZkMPHaFV9W5xkUxfuYjT98Qys4zaIk01bQxvU8oQFhB
XAjxkypleTn7dpo/3BK4Kedxo2SKDmawfsS55igfexLP+nJLhguwCsLKf/w16zm7
BlkC4gqwffdgL1UKlATkT+ocFD44tpzMHIq0OJBBkseOR1VuRFKOfCyVr9JUW9Rf
0+tKy/hHB4DeJ1ZdNn+/D79csIf/fggTDPH+Ou5cZgC+fMB5CXTrNM/oVK1fDV1N
ePEpxxfjo0DuT6NMG+E+dpFEDA69MDPSGINwULRrUYdtPzCLlHEcB6TA1TzUtQpb
qe3cKI1CxZIRNXWsITrhSsxi/miXzVuSJ0M05Ocri8spAy293aHhVLtcIVEd/a6+
zP8OJvgEdOQ43NlvQmD3YWqFAE5G/dQqQZJC1V3ZwXVFczrea7eJZWv0MWUbgEj9
pUMW8BdtJzpg21o2AaKKkIks/CDiIejJI6WguV7huK8UqnC10N4CfbmjAKPGKJ0A
V2wfikSi7INeepC+4Ba0yYhnaxc/WCtPjBB5WhU6/QWC7nsgHNd1CKpExXz0ZxCa
iMWUlUtGS5YHzM9gwf6aOQ4fwXWRR/4s9grtr4pp+vMQS/2PSKHZCe4V8A3mQhfi
iS7l+gunslk3jE1RIkgQ9PN7qmVhOWyE8NbRyB799k8CNLfM+szIyOn8Q5UbMTH7
nuYfkPPi50rP1IIMDWuDRkaoS+rFktf6qF+1kI1dsuLL8tTjkMc4UIK6DoA2ciUG
87Pomv4qTUh0emIQrV8MQ2ZpVCZm8069iFikrPr29xQnKdVvMTiQMK81CwLTYQJz
M4Qunyny/v6Ii8b2j+uAILGTKWIsmpcdSuLVNGIaPpkMWDkUpdBynrp0LD/R7nwf
medC/4si2rLhrdYwv62j4Q62f4t9xIxyuVWXsG1hirwmnu0u9R/ZAmqwTAvX0oQq
RpMAND/i/M6d9TX6myUJSe4DjmGX024siacUVvAZgktAFDDuKs+hz2hT8XcixhC+
U3E+2SOsiS3BJDT5BjUOkBlS3sQ3nCpm06J5lPgz1q20TDNSMKn09r26q+wQ/tui
XklXsiANE28puVrzekMeUxT6IxAVFbPomoS1Ak8kCOnuDx5sqU2V9xZRmjASwgSq
VCY3eunNLUfyiFhX1u2XwsFXjgKtGew9yuBmhQ2mHEQoWWRi5LpJ3Vlz2Z8/0NLK
LrmzE0UZwigkF43OxcWdBfY9MV/gUv2qsvESYwS85eI1l9o7mAIfLoq5TH9c/mbK
nPm6kRI+xNTvzKtSYa3UjB0wUFgdBArgKYwRjNYg4QKtYxuMoT/qmgRSFn4ZAcfX
jepQiGbDrK0VxQnAnn0W1GKKf5Is+8D8qdxZH2EE+iz09p77w2Yd9Iv5BIOXgnbT
kkk4ORD0M7bPdZ0Uf5GAnL6Exkd+EZmqp1m0KkroQt6/KwhLRYb0czOhoEbXam6C
YhbHrB8NZcsVbCxO3xDzqe3S7q2jEakwP1GZLu/5+SEGfNLfe1QZdRg5KqiHKbhF
OkBV6MKl8ls4UeRM4kQcim/u9M3vAYY6S0c4n64GjuUZZi4OH5xkkLUeY0JOwOh1
8fYRSNpUy3HhEJEHEjInpsNsBpbglldv6pu4JkVKOmrcbDNth4vPBTAWaGGgNgQz
vmqQQSLHqPMCkhNCu+4UI3HHDw9fFaN1xHvtSeefGj9uZhiuedpbVPL2/JduqSFa
lTZjxoJ9JSOct4WjgvlDo0Iw3IMAyL02lT81mdk/sBxys5bXBpLHK3oA1hrAkc2F
RAYYPHRnERU9Ff53yn49bNbLQQ3LMlglF8HNe6Tk56gJy9xu55bR27YfNVfVPuEr
/7Z+dBabwNmyEuS7TU9WUx1ZSx72dH0TDpwlOAgGRM6V0CZd3c/XKxoS1PT6kyXP
GD58I04nT5d9/H8gSmpUzRT5J+5GgfRuAWeShQpa0/DB3BBkWuvKMD2i8vCHqrKE
Bpq1hZesL7LY17pYYS79ewU6Y51dg2BIdHvcBCbbwlgSNi7AubDlyyFik9L0U/PW
0VUARm+Eehca0blc/pqNIBNfkcq9SxA9kzUA4LHVHl64y35vYvhiG07M2Gl/yhJ2
9RNyOgiu5Q3DIQviWsfrvQc2y800FThajHrCuFsi8Snl+05TQ5QmGSqzBif4mZdG
Lf+54dPNZwvf9hvest45AUfrLiBfrCw+307Vhi0GZyOUfH/UVvam+/pH+FCDWBat
m1jPYW/izWi4oGXgpWFfNpL0XFWI37xYMKA++GHuYsVgdnvxbyM6z9sC2f7nyMhx
iTZaMq5t1muRLzsCAxxYoLqlF4LQzfzdZrDKO8OIMHjtzDJs6ZUQ9S5NJKdtyxRg
QV/3b7DNpYsia38mdyMMSA2q01WxLoEyPit7r/7l5Zmrnir4NGIMs4/2/Qr0VNr1
AcVoB/ViK8kIbEAPa1GyqFB+g4awYBHUFZZQAPr8DCxye2b24HDmyKmUXeGQDif7
IWHYNDJiwktM+P1Et+w5hvfu39I0IS/mEWhFZudDddj1OvbA2Rx0wZg1KitBmkzM
dxQfay9nhD8+lWsliWMDYTtJ4HXcqPh2gx/9bdjhY/hNwNoPWl8pSpLzSxhKoHgv
NGlzTGFGOw3M6nRwUfnhEDUHKbzZaA65nBr4amjZw0SJUF0XpJKDKH7k6eom44jl
9DtFLZkYE1GHURTlSM0ZBdi+G8V1bf5w4PGIKa5xT6mrpgrPMXQkxlo1VOOwtdpF
70/bH3ZRd+KQSc4N/3xcqbIZwiZwQtG5qW7JyHjgxUvHdGKSQTzP8hWY3cYQDUkm
JZZWFkAdc88OQ/qC7Ma3PraYeWCftlERMvtNGq9Ok0Ri6PslKlyb3sTZcMN3yT5R
fiYW0CnZOq6bTEHlmMvzfydPpnz6kMdFXNBQAvPDuyatwdkFpcjX5DxtAjM/jMVn
0cY6por8fJZC5P/I8uNyun0v0BzSYyMMnZRXXtm8GMRru4DnCrn1KEBVauAddkuA
URGcwD3pLqFMT+RUQk7FQZqQaOqbws0d7ZOOk7yVFOlDwZCPUUGr2eugKtGVARfA
t3aKSR7iC2TK1NtKeKQVIXL7FBh0suTKPpfX745PQKutfNn4woFan4sSliDjVLwN
C1AdHBUOZclFuFk/M5ncxKOeN9szvgSS4tbyoPRj5uSAgyBahnOoTCWvj8jZDcyx
9UA/b+2uh9xHWncgumoHfIpc88kOLJ+HyCSSNhRxv0FU8JQyJU5zB3KTS7LHg1gk
/pRR4wOBil5cLJ2BJLXWCeQWVPLoDnGEndpA/tJMe86wyNLheiYD7ICLn7YJzXKn
k8AuiTozqZ4U2saf7dz1jJy0f3r7dGeltEaO5+5E9Jqy8mQocFleM8ymygZUxj78
zAf03ds0nrgQOho6KTTE+lLngbhtIDKqvmo4ZDM9kuzH8mmNsPaERO95TCdrhEsq
q5DMLo/PTxw6SSrHxRWAxf+R//WabWfDqcwBYaq66Bv679c2jp9/Onjo2ZNkPwZ7
q1tCKWh26o4B8+ug5K0Uj2FgDGV7c7FgUtkWPLz86Cr4vi/jfO3AlsWL58uDRR5o
iejDUjibOauDXWGrSSiItXUyNTC6FTa2pTob89W+vpLV/17CdSesNbdrL39wAeNM
D6fA2RKtd4vilSTjZtKaC2XSRumCtIcK2WfNG5jYU3BTWD6+kBJS9JX7uBO74ots
SaMyHHNHESAKJypm856+t8odepkrbQ5GIMuU18uL+zjOgowLUqNFjxRzn4YX5Scf
POLBUDT+/CLoe2g4CWu2nfJ6CarhpUVtFcQBKY+uAJ/bkZGZLiEjL4zqV5NFyx2M
7KmIttIPuT87VEze4ZgbAsWKvt+KTWM69LJao5mskgT5+IGevMxydtBqiRI1xZZ/
emSPmLg8iDJGh/p5J0ERl5FKLsge3FFidXEzXyZghdnuTt/twbxpHpSK65O22UEw
f1e0O/IizNbORmTIFKw7vQJav90Y3T3iuhyfk523FhnwHgLECD6CcVH6vtdnbIjJ
1f6+rTwZphDW/SQqXNop4tbpAdxABM1C9yxG0CjHZ4flQ0T9hpu+ieabStGLdVV8
BB0iLduGz91ChjoZmVNFj9zrEzVXtXHKcDmTXmV43gJwSI+3fy01B7WUyRBIXUeW
14njRu1q5lHMZ2ZvaAshZuDCJI6fxq2c5UFcENiXNN4eO4bqUtPqPLeXTDC/LumE
uOo5kUGpJpgdFUgALZ188DTLewwcmlySgs1Pkrpryw8WUJOCnqG2rhBIjWpIZWiP
yn807JQVPqg5GtdhFqVY0FhVapu4MasVTbjohPK+TfpNAYF2K8M+FPEv3S7TmDZd
nvmceyzPiw1CKrOe72IBEYPRnUFzDBHNsMFetRyklqlQzjSGYzxUEuczhY+VBALn
6NmtceO7pAN1Sk+C0ujbLjjPSHtUqWlRrh7VAZgt9FNut1UPMPx5RUWnpDowYK/p
06/9P/TrgLy7ZUBnwswB4wbLhFYq4uN8DufgIJGm/EyffvK5cRZJHIqzQktLaNo9
wdoUgnPwb3BRdlku03yxYAgCU/sa8CYix/8S7HsLDFDtbENvHstTtsoUmsANUqWi
yGFvPlq0wBYzGnifNxsUnI+dpfIh5WAhFJNhG2dTQBdHVbl6tV85c2zxm8qEOejL
N33OjLvs0KtT4kZ+SQ2fv+rIzKIbHKkgPAExpFyzry9YtTN5QCFbEcRyj+Vnk4Yv
IfQC/MrE6eAQMiGo1I753rQYpDT2wZPwGDknY6pWpsI5zGV4+PJ8r8yLR0kJD8r1
cv+xnwRQjysqKh9B01pRDhuGtKCgZw26nDE608QZ3i1isj4KwNsxlBFyvcLN/TyM
kDn/gSREG7TvXI+CkVtG+sNcmLdCnEN+dfq8Tis2zHjs80wXsp+w9BFaoro50342
DBcFddyQ+DW2XWyXDjp3xeQ2GCxSjaG9fDN/smWzJJgdbxuKTUgwtRz0niEI+Qsx
YBml9MX/IOc76QVcH3Jckn88UTKJjVrc8Ijlu36347Iz19n5gnpE8REvAZjbfi0y
+Jb9PmkuXN4C8/16y2aa7r+zbl30BkzOVta58pZjdhei5YWvqHrvUafXCJspxH8Q
nA3YfFJGfvILJOkilgWZzjYjYmy7PILiCxyHsNuBOnIRzdlWoYXJegBlc5+rbSPm
o6eIyhRNiMc1Jtc97MbedOvDgWC0AJOrMuDuyGWaPxjjqnPUuJaG+fL1ag1zZQSC
Yx16O0bcy++jhyImJJdmpcAUNQuQbtaQX8kLVMmk8FsYq+AMkrfpMr5qv2AWBKKl
gaMiqcKyj28BZxaaOBek73ZN7lmWG+kW5ggBwJAgb8r/O1aTDTOMn/LY1DHW8Dgi
+y67QmIvvSykWqoO35pM+il+3db8111dvJ4V7BLvXpkl3wHtF2XmMIxEolGYJrdE
wXQvaosap3C4WYVN7IjinImKgt9Vozk+e1qzXxX0+Z23gqyK0EwtizEQwV85zVwD
Dtxp/PMBmzaAV1L5VlvCy6g0ZFqUsDJigA8yEmRwmCTHmVWiZp4kJsuxLzcvMuea
kjcpg7qwIhQEfpXGniVXxVkWDYlusws902YvIoJ/ql953Il3Kwo4Bk1XUaHDv66T
N1Bs4sSdU2ELIFaBZs5Rlc8eMHBjygq5N3Mcld9VWOtjn9PqyIXdgywjPPiO1+6u
MtSRVgSDFs+2iDg833V+nw/qPk8Kt2uZpW0gOsqFZQFvOjn7aaidBvZzvBUpYSUV
6iNLkd66Gve200QyB6AqXK2hs3Y++sHkVMVSRhhWN/Gk6ZDkib41FjsG88YZaUWU
29ZhtQ1SclZnawO5rUnTkXZ+DBJOXtO/ypPUpNjntKL8mPcDTxjPY4k7NcAywLho
gpIpz1lKG2WC3CR8DQ+agsXyVh7lRW7rkuvwUYv6deD6qOZ6V/+cpgfqBXSxJ7t1
UUmEm/V3KYJDPugYYemhL8c4mmKdPPMbcZPyhUVwMyADStcbzt1ulHQR5VLAbG5/
KOBZQ/1KnppHehaMafcAvNb2b3GQ2x8PjmbUUivcjfJ2BjjN9DisTm2hETMyxMCr
CHdKM/lc2jWjcJl/hG33/RX4b4ae+1iJ3kUT8bDihgfRQxpSCPWGVlEjbuCk9ZTt
q4BH70d/EGy0KUjrX2vVxD534W8tsCYBYk8TKz2ullr0wcVs/f+km3OXTqGITJA9
JBakucva//z7BCbzKFBiA1DFzD2d+U5YlIvuzmveThty26o1EykEIFJCIw13imDl
hdYrElHa1I4nUrYEaExwZX1mkwcaHhV996AhT01Kf0EMAM6rJD1HFjykV9MXR9kd
FyVkTaOci3590jucSQ89foaL+q6nCzf4lOsAz94hvBDpqlCuwJU/nR+9s/Pvh+pN
G3qL7ibXjOMfiJKQ5cdvfJotagVJMQa47shprzOBe4QRZr/3EuWD7aZb/8Krukkk
fA/SesbTbQ5dJyFcRq2h5xQxm13U2j8LOI14OHhb2CkQ+lpfAExquIxLusMz9CQy
kzt6wCxbmH4IbCEf70gs9v8C/81uc30vbYr38MDUye5rYAKcDEPuxznfEvLz0vFc
PKnt1loonqFYLFR2hzCCQl1fsGfHOqZC9VhyTxNSStQw1ySJgFkcBlMVsqu4qm52
b7eUi4VdVG8jtZq097yILg0Wl0v52xx4AI7HZCWnRCRGJ6oiANdo3dcxdOrvUMx8
/5Lu/0G3rp4hePsqzaYJ084GSS3fDIK08NswREO0opA4k9BPMDJX8liIz0aVoxfU
WquPrNGxpGNRe/Doj7/3S9y32zZvmGVsT8ExQpRrAFcuAEhZV6KNMBbeY/0oD1JL
Xbl8YwKC7c64ox/wKsbAcdS24AePuG5us7TOIEE2e5/1+tkRuDN7EjZmUNUzhg85
Dla26QTXLypOi27w64OQF76UgULeP4emZRchydKPy6BESuLaUzzwH/hvP4HsAMsk
rfNSpxO/ojatBCpNl5vzuoLvK1jWwy4JMR8qxKXiYoTLo4zqlwFpmEW+80J3Qdae
bftQBLemYGbFoTqHAd6SglfIFh1E2bTbkot4/t2JxPcHePs7dtdZCWKo941Bd3Wq
sGEnpZhDBoJEu8qIyCdSgCynxzmQzRsQLM/GjedEFtgBcutP7QdXKkhPirdWpAmr
/pRj5Z8wuediB8LUASJO4NigWEL0M2wQYJUnAFd1F/Eo3bj+DVxbXrTuPxEMwUWi
80wdC3wPgiDFzlCHr8VPIcAWtuCQ33TyBz7Ppl5n9iQdRJs/P+Bp7BIuYVpCTD1g
sPQarary/M70bSIUwn6Q1apgP/URzykwp2kRZ+AV/C/F9owgFjB6kdCGsyvJ7mwI
/dj+hDrIil0snco0yVeG3HnLXe7p7OF7Xp5j+hl8ARRMF76x1i8U+Qn/JtqWo62D
yrNZJchbPTa3kjo14wcXZoBWim8+XcuhnVtvtuXLimfgVCzvIdfC/lD0Re/KLBwz
5oFA1tkflon9owSybm/su+xpJ9N/ZbCZwC/hqwyLtuxSfwNfDGrWmoVx0YvquQhh
i7ztHCN5diZdzTK+SxxJETiiBALqCw4ZZ6uE0c3f3WarJ0/HS2LvY5HImVXkqs4Z
exf8nofSaUvwY4tOCEx2fm7tv5A6NIAAEuKTLZuauHXH2sZcK2l7rLa9aJFCA2MX
lt0//+DGl5ePVychM8FMOljFB/CC53oVKCm/Q9Pp+RpikHXKQ/6BguVmPhqsruAe
S+K2iAjvh9uGOgvOLfw47hBjbE38CtFutDAVVugGce3q39lACXHso8uXpTQoHo/3
8ornO+HG8qoxNGlw2nt+rRQ1u9dVGdHOwAmrhEzSBdzLUmeEnB3/BmCxrGGuNnCF
YJdRm0f+k0JzUdDbYqrLHsEIym5gz/KE1hZaazvjKK5pDlg3p4OaZGGVhq+K6xFT
BiXaRQs28JkJCYCP+qB6tTHlUJ4dire2BsAGPwMqyyCh1GLfGLVuZUGo5+06mkiD
9jjDoOBsWd19ozk0rWIuKkZ27BeTwdwp4c6cUd8EIUX8IedmfrBnfdqu/U7rRZ/w
d2HHenCHKIEQ3O4CC6/Z1uC1VHrE+TGIcCcz7Qsdeqz/JOQkkp8CEofz9FA8LF1V
voh9s6xUlRTvUHlHoxfUgkbKmmX2ukBOPp/l25g5zg9zzoVQbeAGY6CWv04vIzqP
FCWywNqe9JhwtMzbXpLhkG7nSU62zy/sJvk6YvA2LFIWf0TGT31Z2pL0148O9Pfe
HWRBYlpJPBzRwKiD8I+2e0xG7+bqupa07M/5y7G89Iqd4dIvJQAcSqTVfBKcaZAg
AGKb2C8XZiSisJ2fJ7mmV0OMDP1ock/Ko000z8YSZmg6HR5F8eVuX/DWoVMoOMon
g+yjfEUOsC1vTLdw8ttjfXmVtg/llG8gdZC2rKkvR3OFtdPFiBC4N6mE6yfyE/NA
GXYRn8oqJelk2cahwe1TtW7vDFoi2il08QK17h/xJwQfezHNZIsnojAOCooqEV2g
e4ia0qHW7BjH0YxzeDqWNK3OyZELLvAQLaGZOr2Gge1b6Ng2487BeULHHTyHrLLQ
lyGlfTzRrTUAalhYSxY4FUGWom8JsyoXnvlp8g2GNyaJutuGa8qOL/ifezdWZTL2
toigKNCtnoMpxtHr0+O3KFNLPUzJwQpKzHjZbWzOqRv/H+vg3rqKgjtiKvdj+MCV
0oQzOspZ1pU1syLvBYSFJgflIObJpmhM+FyQb46w/gV6Q/uCfMvEPJHq76iKrofA
XD4x03K2zZ1T+JLrSf6KXszRTHuWRjFouIHpm8nsS19VbZnm20Vfs32JeUunzgkE
NXV/zt52bPe8YZuHHxlnn7OJwnoUDEhKJbKmHLKOJHOV6V51eGqyR3yuZNchxvB2
/GsoVbU8u2DkZfZouwVshLdSQnSo8NyKOOyHxDDc2Gfiq+4gzxY362rTKn+J8xJv
+8taPZk5rL2IzhRU3x3SUYItpvluzSfK615qY0Pvhb9qFbSlhkavpBtjCtB9Th2T
0spPNR4lmNzpKAlrpTn+yScBcLCm0mtNujhkppl1lVRmOyP/py9tme3uNcq5M85o
rzUIpz+TWnNxL2bYaR44grTuQFrmgwqPFx2nTjRHfocT2sYPsaIrMDahIwuyja7Y
TTELsus58tZtE3zKib0jLc02xcpcAjOT4CGmCuZbW8A28wwUk0poSHKMR68RKFAQ
4jEh2+ET+Hv4GU16eB8lgi20hVYviQHl0BsnqGsXnzPCt/KkdWv3s15c4vDIQVTu
gQMi3782K/OTtfMtFYDvDuwW+K16hTZ2xPt994bHMiDVpmRK68jhx/G96S1XmURG
uRbKbV+qIxcgCj+eKFcl2ersd2OV7t7FkBpvHYK/y0Sv5uH5qDLVuooSov4MtkFV
opS9cTSDLeK83Crx0cojHrTs7mPyD6T2oKiuEwiNiDyLrJ7VEcnyhzHdYYsNx8sG
lssIZa7uIoKnjtp7mClyacqNWRklZu9cpthHCJtBsJhiy5I9eaNXCf5/Jgva1gEG
mrghdaPjb/a+OBMdX4BfQ4QTKOdiQvZ1I5Xw72XVf6h6eyjnFvWZVuZHbXT6B8qp
99zb0Ua1gVaqsUcSzpIPCzfaP4vTxlw46Qzg76IeCtUa6cV0Rr7FAO4tI4yzHSaY
T8RXGBwfTEsox0X65+GoAD3HTuc5F3aIUmO0ixyQp1Zki5XJ+pLUUOcIFYBftwaE
moc4tiDFL86xU9rq9FVBJbFR1yezlhYVACbP6iuAvUxls3VIsngCqwqRkloPVPXM
qCirrppjzCbKu7iKiE443JzXIj3noCpWS/b8uMgSKg0m+z2mapEJPjZcy3lJunAC
HttlnYXUGxu9PYOxTuvUqbDiF7KnayQkszx958fzKN2VOPupOIOUWfeafi/DeDuV
MdpPU+RuhWmczI4QK8ZMrtN4M36mxj713ek3GMqBuC3dTTuHLb8s/LNNvNv3zvnx
AED0qAtbs/mDv2hxR4JNVf3aGJ/FPLD6dQF9jOt55dZspN43NwMpy7TzCir69qg2
ATw3oq4WTz1xwJyG4qNEhP28KZWTOJuLgFou8FMOjf8EztEJvB1WfBvMYiQzfiiE
vNS7J2yD2RvnXmz8arsujgzHfR1O8Q5BmJlpZs/dQ2TJyqhg2SUcecZ2DAFcyAxm
o0gfLk8PIJs07U5bmOQtFsQEuNn4JjoPRiSdBcUEmy16z8XC8GuZ/nGnt0si0Slr
+8zd4AM6dif5C4zvT/OHCqzroxfLvY4XLBi7oy+A42+sap/r0N32hSLZFkoTkrLO
4Iqdy/bQUi/0WdqIXVPDENhqQSbatrXsD/cKJKtWCvAkxEKAKgdccU+6gFZ1VbBv
xeyTOYLOTK4S64udzmCiSDUgG8/9sTB6k2ql5MaiuTZZ6jNIUdrBptqeha1nKabb
5ei5DjtO94eyP9GroB+lRScGJVYqO+oPI7z1yBtGIulnjC+Kb3Dej7IxyV3jwLBu
8hbta3yFbkwbqM/GN2zQKHdDy2PahfKCdi3PCvsEsKrA1Dx24b/Fz1PG6dwyPO+U
7RkKAtoQ3A+oHsN21oNaQ3xO37HZZxRq+gQ/Nb+0pJO6nyaoxfuHPC1EKv/prKeo
qeLmKTKeS8djM0gOlPUM1aAFtYN6hIFL+UJjgcI9SGhtHvL2M0mYjRl3XQ4IvzTq
NyGpKdFibBsZTRWfu6CyXabDEINPREiMs0JC3XXzYPOMslIwC5kCQrsAszvBYEQK
LzvvApv1jil135SsiJkbOfwhJPCS4wOedGuKunOoe8nnswRwZS/T0YUZ3Inl9Hcp
fqZt0Xi+g6d4QLa5NlsjKz9zrLczeuQ+QDhb9e1ht3g5nO8no0mt6peOZv0bNWuV
8xr4wvvT0VIMoqj+uIuaBmqMRgekdvV/fy3rVeo/TRzxHUzfDey0AC2m12EGdoQ5
vTHIFQsrZXaQOSPURUFbKcKf4bF0n7L+2WWsW+0XpDg7il4ZxNbbKOkK8VYZwRrs
9OHwYs1MznU3VNcJiysuJNZTAJTqmyAley045Wuzg+YgF6d6tdT1oNh3IEH3O+Fi
dLZp11hU36Ov1rPhehFT7MjglI+dDpRj8DscSAWv5lSiOutQXbwM9ngBFiEk6URP
Z5BJP3WxCVBUwApkMuJHKsX0mPmEYkMvB2bPXr4bsSsK75Fo3hjx21RUyq5CQt7j
WEtUdaks+wcMi5hymqfGicL+KUv0HJwOy8O7bcXBbsj63Xpd970RG/8ROoYaKYsM
28zsyixjDXuUos0oQZMT6P6d2ZxGwE/fo8yKaOhNzsh1vGfFE/qeAKhoDtICW9uz
03T4PgRIWNxuqIhR6260tU97YlWe0o1DcFVQAi8KkIZ2oVhzlHkeQUEY+0UoxZwN
38ig0Adf25UXTze6Wgh8xA5/mRAyzGS/EGwdOBtBs+P41wodSY2zemy0M7Zpl/HW
xrE1cgVrDn8+s9c+b7ZlvU3hOTEtvSaVvlyLbFqRpXMYeDywmQ4yxw7wS6+55djB
Zrgh+sCxja+T3PpOpx+AocBiv8CRaz/eMEoXsiWW3kooTM1rbS9/NHWPb8qp88kR
G4aSp01J/z60eFV8DFbmwepWTYShYo0V2iWwtKhHe1Og44mkTjG9uqsEZBO+uafM
qUX8AiVddMKgiIEt47PuTvnIgs45RFBwLHe2AWWptsLFETn4ewU7l+R73fOdn+cZ
GH+hDOanANWY0sZcWNnVu9xYdC+F3uFVxSg23edzqkMgsdOiKbAnuh6/Ch9xDyq7
Ka27X0+Xfpa39c5Ujhn4uNA93DNSiv98pyIyEAhECL/vJL6IJZam9xUSGYPIw5yP
RrEnHelF1TQDgar1zj3wqNwtOW/oigHlf/d3Tx0CcZdUMt+xOHzzv3FbcWv69vNr
/Ba5V7vRk9xyJn1cl4zhLEk+owKYJh04jjnwZ1pxms4H2uux+Pz2DnZFnZiQ1Tu4
aSEqJASWsajrZU7+cTbcmTOFC999Mc/P+yr92CeExJ69mA4S+Ian2UiTFynnILW0
aJY08d1OpE8OFOgBB/YwXLGzIOmwVl/qT810fLTPGDunrWujfHMipYYBhj+63tuo
esqrfau/497oSuy32PmgvI7USYGxFNS0JoobGvgbCcS0LiM2UN+vsecd8ILcF4cq
XL5Ctnu9G7f8rqkfa1f5ywcxDQJjJffxCRs99j6nB7Wbmhl7PaUzsqRBxWudCPSR
OOPkAtK0zx6OnpHFOLSmLH90aR1PvayCULHYBJ1fjY49ll99HosoTTlQnWNruofY
XlXBbcs6iH3wFHFxCASyPppHZJGKnj78LdX8VJqpxKh6WsHDeRtL0FyWUCe59TFC
matfSaG8ULafO53IDjd3rEvL2vyjOWs2sWfXcwnK7Sc3/04jYUZCQgdNTWURT+GU
weCcWEKaUXNPYjtLr8oKYWoZEh0hg2v3Tu2rn5SgqPqJG+mm+Ce2/sGJJzREgBPJ
WbyUYkwOkaYHO2yJLhuuFNF2MDo7iRahGeGBuT452lTocusAJ4yw86XpcaNNQq12
GHYLlhfYsdzeU1fCA+9HvaA4ZJMdi/52uZUw7CBMx7APAEAx9v3QQJXd+dUbygCx
bYLMmbFkizovIKmPPuX8b9UutrdsQvekN1WzzEmtmd4lQIkt9neg5sCYSU7gF49I
Ue4oiV6O7yg2vYbRgBeMRClfaZhrlKYic4JBbqHRuGsBw+7iEns6RXk0ILKhPiLC
JVrVm3m9Om8MYiyXN1PMWvwB6mL2II+vHDepspIVPd2me6Ql5lv1z1DLYCoOIzUZ
CKNyWloQjvkyMbNsnxW6x09dHOy5sG1a7QQ1GN9YoPMR+DcwDON++S/ImOXMXc8+
jD6H6xmocWLe0KtrErP5bWvqApUetcqA4bAqf8ZptU/L7q9dZ6lr7imXMvxAK+ks
qVKo/ARz7Bt1DsK1kA3vyKOpnwmQlux1IrVCSIn8kXVoG0bFiT0aBh0BYF7glGHp
Hvlbl7moNIVqxkgHFV7YGNlMwvgU7fhTchaJuH/VgFMwi4r4zk0L5eoArk0YfMUa
eEZ5tTWxBNnNP3GxJVSamNbGx1zKHOCUxlNDpvIzERldVHjd4fcXE7dk+FYXdMu5
Za/yMz7N4iYmkPZIzO4w6e1A2RgW6Ad0FBgzKeoupq0khi/B+AB3Zi6ZgBeriWHo
rpyMDUqiT7BMFWxEfvHPe2GMcVdW0gUTV9qxZTIXTqUkEOUox++IftouBHJPzTqy
FAOnbj+6guOuz3JbQR6tzyuWzkB24d3mu0cWl1dkoMThB1gnUgZkDLzDb2N/YFlH
q1GjoMJYR+BsA8zT8QTogBJeVpTjcCEXQl8theoF4g3P7VnVafrnR6CcbMxDzFhJ
P0J0b74vgJzDOwFtw4pNBd8icjM5JN6Iiq9mpxkImQ9hXgclLxU182PG6qqNsMxU
kZBsZ5G9aWjbsQ09xE1BTgCZNAWZNyhWkLPQpRU0BTSm2pMCAPSHRmOjrapuDHZH
hn3W17cvd9+GH3EmDcAYMXiyN1QRsLMzqvpUZ77jIjKRXvbdZH+kLFRgeatmNISI
acMU1xaYWjYHBZ4Dkow+bJ8xqFFt4VLh+DXm3gNfUOqX9AvFbtz/Q+ADh8Safoyg
GcU15m6i/eNo9WcJS+2MEC3MZjIPB/dRfsR6mZI3uh5BNFQEowjcIzQl/4/3nCzN
nX7rzuD8Gx0syWGcTGW/vb3++VdF51E9IfzrWbAgxUABN46sCUGhB/E6bchZro53
PsO2OuHIzOSPey1WYyfF2PNgyj3jiC+mPkThbJUBQx2goABAfUly7DHl8mzWxSo5
FnfBNDFvIxQ8o4oWfg78GeZnYYTTmfkAtmHG6REAf0AK2UZjOJk7f8ULbcDgpOdJ
/RU7n9vVimUuVa50Bz5yTv39A5PW4DWhvhlGXzVdWBUWoKzfTuWzenmmE/ndkX1D
YVVCn4CC7OSjcYKGQNXUaq6mwpenms+pC5WBW5iTOgoSLd4rI2nhN7rSBZlkU7Q4
FonmaNdDXBLeaaulIpE3moDUwkNuWvdkMVZodoaxt5unEm4cqfD61dJp9xKr7nHc
I+/zXfhcg7xWeJ9PAaYHzKjptLTY4DcDP/A4BBB8H/nBrVwmucdXqpE+lZtwlX+7
y6BGYT4VRxNQXIhaFWBwEjIJN5674AQFYkMy3sxl0Wg/IZ3Okf2XjhqDdX4Cll84
grKknWTeCJhe+eXNVeX28mj4xCezS0IrPzJ80Wd3e3jrOrQZlNpbkSSrSig5N+Yv
Up9LVS14c+PS7nWG0jXGq4wBhajHJ7rmx2UZ5r/5JoTD6/sMSceARBmvjK6c3BR3
m+yBZBIUSvP3oAPQuMpcH0GSJX+mT0dcnLEvUEgx6uOXlYFqLB7aCyVlcEutlYb6
lOHP2WYi46nZpatdYXcW8/sMj+i8iHq13o3iuRYRWxkOX0UewS54kcjdPHSxLw4a
6u0jwmv1gHSQc40OpbgGPRqH/NHOENKOvrvAI5zge+aVcoO/cLFH8gTadPze/hEm
loLqIBJ+eqDaLfBBcVHJTvae0HdMipf9TiFr4gS8ppcPU5DlN37gkDC94xJ0Ghb3
s4y2oVus1knBCsG2c2b5qR1RrEaMJbyXxefh3tonn5C3eMR2b+8NiW60AabzYn1J
ohZEvUroryabESZqgymKyQVpfUMJHoRvvYLvjweAKHgYoZ0MhawMgJHyw+EX5cAQ
FIcMYVhbw1W97P+Easznk5B6B3KGo9eYat96v6uQ/JuLv+o1ZAPUX3w/fU2zzj38
mqu1RscCqTPEChJuDf2Z3zs/iPJN9im8TDYoRUABEsMedtbL3LJe6gg2CTFHJGAQ
0aPSh8fPSwU+wIpVcROudchVZCOO6gs70Ea9+Br06CyjCxNzy0CSep7dw7VGSxe4
9ninNp4OIQXZcp0WZzoPRUIblvnHlZl8sgnfN/YCygl/YZLKYEym6oImzI88EBvS
4RvfvhTJxhB0b/sIrQIa0imHH/gR+N/uSE/1V7zwc0YKJxaxMrVc5BE189b5VqV6
Cd4jCkOznaatyLPQyGx4y22RFasN6pu7m15fDkW+kKlb+dqCRnCi1oESoPg5Vy6l
4jYC9cSeAYynULyKFK+sevDIuvu3F9EUgPqODVysCEqbfwHM6sHOcWTOGZLpXFa7
BHYZity6vSYKuHwn1hmhU70jRIO7Z6U0sQ+U0B0ig5GBGtDygJEp3wI1n/IfYTGc
zMU+vSR2Mm77HXGmUgfDtwEaUtRkRh+Ra1GXsFnkf+2FDcSRzrLtZrc9eJYkd5W2
rixWtOG2FBxoKuNvId1oMGG7m6QiWwGRhyZhIXXXEIK6Dzk7ETDXVYeiPGrgGcYo
o12A2KvpGJTo1R89ao1hrGezkQqv18CMh0I5ImJVHHMmW4EqFJ45xzKFemiJVgNL
D6FstedoQa60hIh+zkBcFt8HwtUpAsl53X6zdz/h5wUUxl9t4VUqwpBELri0Ezog
OMCQBlGYoINE1LsTlBy/d5Vev+eXXYd1Gh6vC2pFhvEWvp9/F9CAzvHhWFqdnT0S
n7XKBmMZQMHtnOfOs2of1IFVE99l+dplz/3pcAkxsjLS4wcPFA0/oEkeok84Guo6
BYPvLhbjelKzrKCRFiWSf98HFPnxqPXLhfNpD2ZEn0LKPBeHBu39gyIWbYXdSRbf
j65yFihD9fsDsgOpnPoXMbCKoft4dBQtvUZZAoeUCdiwMBppCbtKhE670cmNKcx3
UHCuS9Q5fM8fK0M/dhLcqx5POW7KGFLGjP0syLq0zIKycd/c1OLbvftfgpVhrSPY
JUDJelq8N4nLPcsYgfOcx8XL8rzmTjwWl83Cnm8qqkQy4fOmd8Fg2/8pXBY2H8b4
fuDhNa5wGggta/yacUGPULH4kUtwt11OVsTPtad8dPOno425wLqzPXZMAW7pUj8I
a+qlTmvz8TdJv7nluojql0sH33VoDiloSMKk0ydiKewIo3Fb9i2//CM+GxckpGY1
EBXOBsxyC+MORYUYRkt30oBwlV8w4PKPS60s1HtHvUseficTbFigpPmIboAiEZqv
mKoA4BmZ+3aILPrAviph+GTtE9AWH9P+6nI+kqi9urijJpZg3omBuCMqfoXpJc/y
FhuZzF1Bh4vZClbGvSzojPAAQxrvtF3s/WjIzp+bSpC8bduDP1bOymEEgShbfXhV
7gVCap5W53Ju/ak3QtQIHSrmlsShNOmwXg/c4AqRVAt9P/kMm4zS6eurbP6rZew7
RPpXYwY1vR6pZK9VQL9LAbq1V7XjzIrjpJDXFcB/Nmdux2C1RTvvtR/GCHkdaBS5
QZHMtJcKFRcwLriAVvx4+hSt5AZztEgb7gRTXXQsAb98ph5XRM64mOQ6n1VKfTG5
ZOSBBg3PSzJkBE2enhzfeeAFEEvOVIZasuGnN6/HTCGUNjeYq+3DdlWJsCXDfXme
O9GsJqMnDCXrwmwE/gsxb6Wvqri30XXCBExLuYFMRCrIQVMDgDVt7QCsHoKzbLm+
gv0E712UIhQSj24wdEMPizH1vcQ1SXhMg87BZBtzfr5FokHjDE8fR9YgLaI31WLh
CvjD4i2V4rgMnkLIxeMeBNpeJo60347ve3eSfH7mvJcmtxbBHvocPY2hY7as8aR2
pa9Crehxla4Ikp1WCHiDM6Pjuh2qWJLEoFcv5+WFrz76V6l0LtfCzRMhFEOMHEg9
3mQOetp7AtbwzwJjpZMUUjghZuSyJUK2VBlPYSO67XdB8AQTOFY5rEhfMymtHxNH
GF7DluzH7BGdPLSB37MIR3UeiFp+L+THxTzDRq9P+xuMId7s41QE/W5Rd+An4FEp
s10wU1mRf6xLWhUYnYQWgGLnaNkOtfvgnvi41h5GGAOynF8cNzLgdNyKuUdJlano
+5b2ZsQcKHs4w9Ui/DcuZacRl+NPldMEaVk+HWMsaHLwplPAfJTEma82hNbXDDs7
IYl1/iLz5g0MiB/wo42kzS8N4FQdqHRbW/wQR/SftW+v40pg+T6yI97QMcsM30nU
ZmGePCbkiCp1a5LkovYOhRBDKvJpV+DeSuHJsxECjxT/ktKA5l95DQJ2yZgxe7lK
xRXV47JGMSmw/eCbh2UOEU+GFiBReBmVm16wq+mmZLooil69MgEwXuUQqNquPX0F
WKTSD+Iz7aBzwEiRlEx/kimVgTGTsie0RdoVMnaesqC8bKr6OXtm6IyUO0W/M2j9
Hnv7/Gv3o9dVFowCxVNzsteFStv19sDNeNG4+931xmvqeFiE7FdUIcZgcXmcF0mn
8rOfrIhKcd8q/Ia2mW8+yp/cYRbmuZbJE3yhvh077ZoIh+BXf/JF+b49ff3n0c1d
y+ymOJiUDs/mRW+LEdLqVcJzORi+PxMz1X+Jfi39YlkEYIPZmaF4bTr9z12+6lLT
7QNH4QA1X3gKdsvh6nOmvDoccZb+4dztEsafP2vzumkyGbDbpXXXvoEye/hifx9T
sdP81dBE98c1fFXhh4y4BZhj8jcwjNjDzKruKFuT7TLsqvz7h/EMpXd95S+BQHwK
SfcaCSBOdOFb7HIpffzIL18quCaGHeKIRychyAj5/ahigjG2u/FiPobZ3NIA5zxv
l9wR2lqoeR1Xlq7CEt8ulSS1MVUPhvu55P1AT180u0tWmZu2FIUjbUhmKxc1K5TJ
EBI6MXxQI+DnU0zo7BsHrPeY+RRLEu8BdJn76ZKgfQ8QoQYh8JvTUWi31bALtgMH
lGhSYeYH0TBRDIvg+XXxlosx6xRFcma7JGGvzDD+HWPDnHE80rBuDX3kadCIOFOf
6fOzPDrswJj/CGzB+3w5JWzytdqh/+/MMzfcKK2lv8P+H3pTLX94vDASV1LR9GsQ
NDgnRxe8/TLXPI/K55FdiepvhE10kjM3QQzpL2pK+iImPaFs75WiE1JBauE3blKP
oFFAR4R7yalFOFa12+0L4UCD8ZAIi107KGo3vViErrL0XDZVpdUa/ZnivdG4d9QJ
2blqjd+huHEBxOWz9FRTMfgqhfw2UcB2YlTlOWO7dAdAsPMdm+JBr6LKsb1bXyB/
B9ZEHhS0H6wGixWEmcd9IEjJ6KFnLF6pk/JIyAsaUQ0wjM/YLKAMdzD8db5DyyXj
JPQCaBoAOm8Nt4OkRk4gte5ihevdhL1MryO1JECScy0t7zU5rOXY514E/YfQiSxh
vHLVUC+y7U77+62RprDvozWkeDmLOQrindhVDBKw0bSR1AWzQqRZs4ls2JjmtdtW
H8t36Lio/XNhG5wErN3hOGbREevhcioH+QwcDXCE83fh6bbb8ACzddhPDh0CyNiS
KNJADNZadGYA6WMBArkqNYNFvpBXP4hi4BjkbSqRIWZrIbTEANC1Sgy98dQqg2wV
dPDFPu1w0vMuxx9XUfqibVd8g5dPGsgmW+2zvTvZwQQa6lXZSXvKiMt/vXvRbkdT
M2BAIOR7w8vkiqIsv8RWWB39+BS52wtRcNjHAoXX5VFze+Wi41ot+eOOKM+Ud7qa
0f2se/yjzFRrt0a3k6beT70fh93zYdaT29df1t59ajV22yKMcI7W0b+rtj7zhTX3
OWkA1w3RSCqoB8gfuci+k/qAcdWjE+p6w81A45q9QzEGU7J6JBUsHRTOlL1NlBTi
AqFG1J0OCU/B3mZihGuhMRBnU2isFTObt6rD0mL5O5VOpU+JNrYdDVnWCx/9Gql6
pzFEcS9RNIaSNnNY8CgUnj8jS6/b6fjdvN9pBx2pl7iC7JHt8VfnyL5Jysn6RFMb
Gc3Mw3o9eBJ2jEVgiCEFNLleXwMkRDefV3G8aMcCUSIQVRVknpUWeQ2THVselTZ7
ivu1IaeqEtXLQnCtR0+sMwNF7liX455kKe5Iw64dk86Cc2sg7mKYTtire9Q4KI4k
TxAtcjAjQLgVbSS62WBRBHOBwq8dOQhm194Yqv/bFW2CCAQVPrw+H2jA4BObtNtv
Q1iy2RSdmLZUj2SMf+INgQUfmfZ4OYU/HVSTTjEyEt8Q44/yLwmwAi6n0yEl2Qce
7YpoJge5LHIxiJezyyjejkkjYjPU9W6H9WLbrEb7iYsr/yym4kKJLBpOKLMYcQX7
ipNw0qB3FwKiie5/eukFIfO/rFNO8XcIz6GZg0w56hIXpKDuZQxfqR99ywIqWkhk
fVbt05CSjUh7Ov4CX18ZpC4e8JuACDxpLBTE+wdg3IuQOOFdMP0dYhn2M5LkHQbm
sD5Fx53nGCCLD00IWX9g8Z4WnN6JTnCWnnr55BMdy2+OKkXtmFyHMJhNeh7oF2RA
AYsTZI8ofIW/c4DYuIgoCau488C+391nlyFAqYNaaJ5FrGVX6HHthcZYfBjROwV2
IrrT4mIFgQS6c+YWWgEklTshWwpi2LVdhB8YMp4YbNADyzuDi4liBiUnsNIoZLRU
Oabqppd+nsfNXtMgQi/mzzRLwesL/MmBQ5NqTZWYTa0AdSe6Flvj4yQNNqySsTfc
DRsU+ktH8ddlFlEjEHjpouixsebdyk7MNvAV0sBqFp83fCvdRIN5oaYkZJlWvJX+
Kf20mptnl5glo6LLA2tJzfS0pTHwe7+6jd4YpRkG5WglhSrs679sjkfGA5ZVwjfe
XAgPiZuHUzO6yWByRDgZUZCvoWAU3/+u4fqmDakvoFU7jhqUN93JJ+AQcOtHiWkS
sUOnMU8mxUfcJ+1mpjh+tyj0JkJJCaf7yQE1Zr+BoUUmlWEI55iLgyEeaqimx1E3
0FPa14xMaM/M+OSVIMvgc+AbypAWKXb/F9dS/9s0Cn5wCsjKKQwCts4Xwy6pDCEY
ZXd8uJ3sumDg3V2YwqikI5fH9oeFkRubv9o6dXrdkxCUnw9BbqCDa0pOlDV4xvah
bj3fN/LOh3nXtu6q4o1j/kaHQ1/VrJvL69/wdISUafriEUA/ajJpzwRGjkJfp/WL
2+41haIthqaJJfVs3VqY+Qf9Q2SMpCmHrC+cVTzsJKy8U6e3lOeejsarETBeHDQE
ZpAFZArJufKBuv5XTwZEkjfSfl7S4Vuw8FOQMavHoJP4MRzLhv43A6/xneKnIaWc
t6pBuBm4FOyLYJBGOY6aj6A7Glr683n79vjY3NKf41TpnGo8y/sdDBKBgsAg1fHk
eI22sUdrF6ASCklK1xMUA9ffF2prvR4CFDnh89FiQb0b59FnFMxoNnKzGRqvCfZT
5TuHyYTSTEmYGNucrRSeAMWEfI3TyUnt5oy7h14LCcYTRzBT+89FYjwzcJ7dRyFB
OtIgi9rDgQNDMHT/21IO1mZI6kIoSCR+/6cSa0KyS8jCt3QlZw02FW9FE7sMDGCm
Ral5GD323N8SNASPh9DFVwea8JFZX+6srNv14ksEtuI0x36lRe4Qjz/2d9m9TYIL
EGs3nu9c6OF9bU02UF/ScEFB8IiM5fUkDvbOCdzTmj0b4P1pzS93VxmuEUFHQILP
vITvzwfhs70bqS8Hl0qWqml66olvSbg7GpTUw7RNHw3cSbcfKHkzfEZt8R3vY+CY
uXzFOghU2Rv2A2nLzNe3Xa3lcEWGQmgL1wrQau1IwDuSGxjZhjC5350rBSohMwiQ
KAMaMjYIl7u0+ntdHy6XUiBXoFe129byt91G2VlkcE5TP8TRqrkDxm5xFZe9tIDM
JCg3YRlTThIlNb2VMKMTY8Jd7RQCcinykc1xUKPFjDZ0LgPzm3WkooG+4fz4Y4WX
s+3SfXWxh37pvdQVreV6E5LGEhZslR1480BJsaoA0agWRsSSSB6rMaEEcww2kPuD
1IvGvpe8Qw9is0B8WwkB260ehL+oe+Lchb1ITh54c1xfYrBuxVLeFIP1eCkBtuAi
dni49wY75MVtOQ9Y5r/pSGUDBHMJg6oAC0J9w4LLd++B82uzkxpXIZ8Jm5gdKZca
nlUzXzyBmmlvET3VOYL+IYBbc7HGDOErOa19frUK93i1ansCbIHHJl1b0kdt6b7r
/kWh38r6C3UqNZHvPZMeeC6uaYYx6pj7pCHzw1o68efDIt3ajl1x52kQbh7hqtMB
K9zdcYKhi6GEq+Suw06WEr66Wzro2NVv/K4YdJndCXahCmsJ5tkTfe0IlwtsS1fF
ZGfCfahgHn7/xryHcyWZj7tOPiOYXppRmfQcGWIPCIu63ssnBBwJRy2yv/q91j0u
fwcIFYOPggIedxDm7S/M+IiF5L67gC/ONF1yVjMtXpjESMk0IZ8rRtanzesJn2kq
mhM6fIbVPjVAd3X4AXIJAO75d6yXNTS6md2mOIC53tqMJ5kDZktH/bRNJVbjpMC/
XHF3/RcHAEndYkv8JIUWcYwtgwtEI8vhhg9l4oWD8L4d5PAA79HjnRMjumBKYhgO
HIZr8y+eHGT6BbGI6koIxMLFoNZwHV1P/l9vBPx4pr7DnmB+D602cZMvVKxW/vLu
rTFKQ5iHVYAOhQA3k4HxkULn7Ag3HVQd8AGWDjonVc2ZsAU8hEljJ1cuViRaa7Np
RS47q01n63OtQPjCmz41KLV69BDzIztInGXFI78POKw8rLmB0N23aZdaLN74KRRc
bi1NACUMJHrbcorx+Q773dWVip8zoLdogXrTfjWbvn+azeNfEyCylBIBW4RAhlqA
dixX6NxRUtwBWwPad5qc+SurvG5+FbVoTL9NfgLWzZDV6JGIXQks+drQXc3K3xei
s/WtpLIGMWDhQrTd/i6ZbxSgmpsTPpUXvPfKvdN4n4k4QIfljBHtpmQN+8OpPzRt
+iTRPbmoYbBNSWOXHBppI3/geHGZB55ObIfRwUE10ulVWjyhdTMgrrmJUXmzOvYS
Ku+pe1CPQlSrQ5LWFhd9lUz7uRwchG8P/yyzoDhATpBiEeNQoN926VX8TnUbEEgQ
S1cmeWlaxQJjmeEV9qn67jQR0s7ihN4OPsmcfpJvEW/LR6q1t5m0I8KNO21uNB2Y
kMJhW+sHt/ULwMtuoqp2MwNCxYEyFuXwFcnq4mKKe6Z62Ph5k4TUKSzs9ge9qca+
bipNwHqQ7puu87/UnVvfE8bHPLdju/qTy4/nQa48rdWlxOVSh1fIPUzkoFufAHrF
Yk63ciUue7ECeg04TWR5vzvcLx5/N8+Sji9gv3Jvt1JsWzVEQUgkvjNrbsrP/raz
k9xV7U45SfudnIVPGen9tFwZRA8Yp+kmkPna7kGhx0vkZhCjIX1JSaRljOvO13bT
h4YCqvZzPoy+TPFA7q3k9omxJB/hWfvRqmPBhgHA+hvN88r3cd0fgxaWPW0AUHNM
XQwlpKHXCn50+3BCccBXq046aowTbJFticfO2HTdwONjEC+0jN45Wr3eCMnBtRHL
zpX2tGMPWckl+WBsNj6pRJAUFZiqLQPXwOAEd+qK/JD3i/Yf0MJ8c4j6hAt2C7Gk
5CZ7AcXSNww4AymZrBIBmuVa57aXJ52/3FC02YrK4ODKMfYJB+E7kUrNPRLtXVMm
HVM7eVg98hq7Ac6Oue5PAWcZ5lUChe3R3MUuH54oXi9EcfYqxa8ZkqBj3pqFvYgL
jHg+ISm9kQ+p8tIgrupjVjwMOfQl0jhUVM854NffbQ5lETFlfrfM7pee6G/xkZCG
5zeXd4PVM0qgcNzVciCqS9TDdn2gXjOHvMp0I2hNeJWbFSoluaTWYayS5dJspjfs
DQwuYh850jJfsrbPZHwfcZ7b9+MpujJfqy60sJMaPvDU4TfM+PsoEltN9ufWEV+d
edY36Qh0YoKNNMsPJA+8ARAbz2zK+RykTOjyIPV9ssI6+f5VVdNXkR6mfxHGWD8P
MEyuMVCLuHZZuzb1LmChvoujRp6Xc0abATmq54zEgwn4BrQ4HLETUnF4AyfYWtCj
7JjnX/67Orxs1XDpXT8HdS27kI8Se1jrHJmZPbRN81tPQq8HQcv8yjuptFzqbtwp
qQ55MI633SY27M6ZiNZvyM1fpcHmUU9JxTBHHl75/o65H+bxIV2q1SAd/hF11LOA
Z3uwcwTNZ5mgr3SBqufvrtkCLGKdbiLCYkUdw3QJiPJLngSDm5uRxv2CRaymrJDq
qOlR4dKztKTP0t2P+wIFNNGa3X6OXeTd/QSU3mq/42HpwZEWR8qDyv0SwrvyBp0T
HljNkr4GQncz/ymknG1BID5oHpo8k8gCLHwnecJCaIYu25GLz+Sv5/4zXCzjn/Ib
h7/kxRCaJpVMpkVTVZ44sLhOL0sUQmesjohFKHM2lAizVx+NWW6vbLk990FSAS+H
ncBY7lfOVHH2pYi/zsMxtBTk0Nlpe96v5YG7BxyYK8W2upVV1mUYcwVipDtd9G9m
seBq8jGqe3Y6liwwJ/9L1jqdw4LVfaHVih25OilyYpaJuz6WoJYA2prVo2wJVyBB
3Ag5DgeFkQkvln3k5maBSlW/BWDiv+Kec+1686osRuMr8JL5slfdMsoaXUPJ2Llr
0qfoRBtvWl7zCP0FojF/tCTaD3SfBdCWAugZKmisQOf6Kcy0iX17vxRiOl7RSKIo
8DYMewn54kHbkLH3PRSrWCj5VN+CkWbHRhQMYSppv7+sJ0WgAnOGHy7lvfVs3iVw
nbtKOuDhJtW7JA7FdP52zatQw9NHwzv+v1cvisebJ7nm9lgzHkZshSc/nnPdNDbm
xWosRnlBA7ohSRlAenUAO9dLszvMkZUWODLwrJ1TgZLnk9kylrprj+Z05WX/BpyJ
MWt5mmFVcoPQc0//GnuPWQ0/kLhlLsVi46UJopY3QM6QVwiU3MLZIel7m7CAZ5DQ
6SkINbFpHboQ41skV3mQBQCOtZSKDpWuWYzjJuesLaCXnlr7L2rgE82uOb0tZ7vh
o//DxSow4DBnQRWzrXWh0e5DQm8q5BKaz01iidKga7LInHg3PWNIKA9HtcrT2d0A
/nPXJudr3WEruJVINTDzZpjRwLh8n/WFZjJYnUuYgGDuvBQs15oZRC2cwM7R+o6X
KZygFnY8VOWSI9M4u47TsfAdlaQN17qGzyHYwHw8XsiTUNSGED/gLew5vY7V3FU/
XgvTGO8G6qNY1f7F45xhFwzgd8iVGVjJWFU1tYDEBcVeMfgp6Mibv5IyYVGXnQl8
rKrQwphGSIxBuiWPOyX3Ut8Vyl4L30VZYd9leeEQCIhkz7YhyQ1l6hx+AwkykuT5
x7GNQuB8Z+Q46dsyJO7GfH053B4F2p9NicmQJ1faMhyLzEXjX9/3RsyLNBC6saqV
zvQK0lqmD/YweucqtitofjEMRBJSixq1SbBkDMXwx1Tg3EuJBxz6CvHKY05bJgvU
j7bmd3EGDCCJva/gZSkdq9/fh14qpjBy2l2rbh6CL8ZQA6JTZVZxpDNXGDh5hW0H
nDFxuwUpscmUZ2qK0zdCHyqd13r+rleGeyFwEnDfossG/3NZjui6MEb5mXlHVYs/
oaImV4ex5QWpYthvt/1x2wU0vZ+K/XMsH/J0zEzpwNnCNvqzz+b2UbCx7/lZQTeH
KfFZ7STzG72eQ9aB94QZ/PM0ln0QGIAA6HgcZCqsompxXmw9PESZdmQS5rwcpBwj
lRSQDeKYs8GmLQYcCrotuDhOfgtIDJLAkDsGtM49//ksI128aWw9q2VqgJOFVFHH
KaTXne84y9BHy8Uq+kW9UzhSKJuDWf9KJZAiHCP+SFmEZckdcsX0j8Qm3kHmN0I+
lUt9yYM3E5MbIvSXKJ+G6aDq+/cM63gkyuChY/ANoe0HuMnclYuNc6AyblO0mjok
+jtssuErAL/qtD91VF8Xe3Bji94QWPNiPkY4DjnGJNzdrn1Q3l4A0KV/hDoRHQ9F
bqY7hYXcmthj4LjjRLsYxd1ESkFwU04+YlJgQaSSCYs/F8Vzl/JJqRwC9CYtDpSF
alys4l1MZEAbWl81Fg2woRaJ5GKoPshIzo5BebknMr1ttH2M+bXgN2/EgaILtqgR
17dMmk8gdY5FGDmq3ICQGm2hgFf3AAVKjA9Dq6F5pYIAAi/pJLDyHwRdUe2AT5ic
j7HxcD3tqA5TO83/5oniGhQcfCbJWe2n6PuRmu7nuc+pADjwj47ZFAjpfQow0Cwy
1hBx/M9r8YKGGDyms9yUt2PfLRA5gTv3wAecqj+L0+uq3n+hmcg60SEapD7S/Qg9
odKJqOYl3QZQdE1q2eYLA/0ylMBISCxhp30btKuqYFF2MfY+PODdKZo3QfN2nh7f
mtSPTPMDXOy4pW1wA6Uf5RBoCHKEhgiJS0Pv0viCtU6DJLXWdBqwwb+KHZKCEHCF
ZgRyEiSU2jLryEOfqvgZZAWo1Qkh8MiNNAp1YJT5WofmvPLT7i5Cmo9l1mQ/xbAc
NV+nL0FkVxktTA2VQZG6vvvMmGfXo7wqY3OBzsJE41aj4r0GD4/lTeHuxB54exXX
7tf8tV+G7zm5GHgnpWi3RTzpCKMqsxAzJk6IsHdR1XKinvOK/ha6xQKhvgA8+Ta6
hYfXifcdZguH8tIG7xPLTMAk6p6q2ADMSETNfklJbg9SIOd8ZU/C+Jlf8VVQeM3Z
jYFzhCrIzj2z53WtF5vEeEvBgcPKvRjnZdjbzqe/EddddQkpjJrwySAup3U53Rq/
Wxu2yoPAWWzbSHLjM0qekSlqkf+4LpHFbA3w3APsNZxJs/YjvERQHfKkkQZSB+94
ybfPLCIXKjecUxPtCDP92TZRsrUqU43fV7HHtdTDvO0g6aXdfgoMsxpnwDhHywFv
qUsWR2zj3BEOgmB3kHuCYESuTpPAZD8S8i0+S8ITjHRdSmFJgJ0fOMAa7zh5zGuS
hfzZo7/7Fyxxeo0fMPojpvPGcEX+cg6MqyPV+4ugD4kAo9SFHgcm0/MnVAybhI4r
+4VrynwfY4KIBVckcZ89/ApWoE5i+MG8BXUsbXIEAmDh/oM2/dyTcrdj+XRut0Po
Od2YuB+b7lob/cRl3r9tp7IEnNCxvbIXlzi1H9LRy5MAPYTltnYzUIcXxgFyR7cA
VNzR8952DDXgc8MzacSOs5glQdj48qYoQAeha2EitCiIgu3Q69Ex65kp34K9WFsP
Hqi5lD7NpZA4xSIywRrRPC7f+uphPfsm26okfSRSwWbYB7uE+dfdCuh2HlFk3orY
GLSqJUYgb42+bfnPuJaTGhvS6Ww1Ai0bhdxaGZCmXVq9CRHqIextqCEsXtIETKLf
LzxpYXDJMJfcmsh3o7FQBM+V+vL00w91/mNUYh3u0qTQ4ducUDN77iVEkl+V84zP
aWzPhMpZ8BamyeR12s0Q7rc0tj8aqxGtVOg0lIFQutcK1imbOPUVJBUlES9IaR5r
tK67b9QwncN/5brcmfxZI6Sn6d/hTATSEAufXmxvQeETtW7Xj+1GykWrrQiRREbV
XTQMLuLrgNcrkURHfRuOwu8mAJ2oMcm3EViS136WkaKNLyViZRbq5VXLY0vN4c98
xehkROcugc5lzzSfsoPHAsJpsz6Kb5+giFs3hBhBX9bS6I5K2LIe0f7V6C9E/txe
4AzWPiAegIMeXIATgU6qACqemhXSlCxIiKUxGA4tpJnZzxgwkA3yyNUNwTP673mO
HNcb1rBG2oJV+qulCbmwTEjZeoMQIlYQC7u7FfdSwRnMeArUFFf4aPs8031G+nSZ
eVosdUBINfMX06mE5v+bERVk14PZN+JLkOLJt9241XHGXooQxsr4lla5DbhEMr6B
Nk3iDszD/DKaRnwVQcIBmqLSLelYT4AmsLTGSMaBGGDN/CDWoHi1acAm8n9U5ePu
WaiXwMQE5jUare6R1K2fDHy7+wmqmyc1mbTkSA7TfVyCdi1zFv2sFPGOFQ94blpV
Ir17/DGyb+BAMSwzlkCPkaJAxtE5z+rTjDrnjzY6CGNUvWdMi1y5ajzymxXPX/7k
1sH3d2YVzVsYN5R7XbxVQOeyfgltPKEw458vU0mySnUBzkL0MEqLAF8g1IsSwbWY
cL1XHMi1ewfSi2+VFP6iLSV6CQ0HGId5FLF9CuSdvWSj+yOv00VQMkYn6QLhtwqN
UZa/5/ecXXhiOyMEbsR8dl+fd4/YYRNTxQCX86sDTOJEHybXzcP5MZgFida/8/Jz
kEqi7YiEGl9RZmF/fTHnJlZLFxAnUGPnh0zJdsb4S77ZbmqpZcLrK12mq17d9lfX
9qi0zM2ybilWdv5Gm3V/33eUVSb1uHNafVyPtWPbXR74auGop9WHWrB0XTNwOGeQ
A1+pUWcbAbPr1UYTDFdgmwZ5HneV5G2aLxunwqDlVehluwQ+Hf1FflGuEYsb5rY+
M4soYDkng6DU0hJC93XSNRn4y6qTDMiiA1HBADQ47sNkwOyZKhQBNVvhWak3xERO
GeL0PP7+vOQVRSGzBz/ZHcX6gCdDrfZkdu1e6gflL6lUK5Vxv5QsUEZziig4duTA
y6iVG9WZrb04Xa+fZpW51tGUTAfJHGK9Dcony+vRm4CoZ6+qOSrgBaDLQuChTAcv
rEL2vclCdUvjTlc7sNFOdIrH/g3HWfhatHYC2X6cpChk15KD4LOm3tZ2fZ2JyEzN
S8Nvnfou4Gxg1f+y1RLITm52UbwPNWP06bgA6x9m+0Lg/FasIO2X4KTkMD0XVnD+
49SRCxbtDDToz+foYJUOu/mu+saGkZArJmMXtP6gA5COqajxvc3OVDSHiZo7kAHY
AGCHVkfsRVVwsuJLYhe32+uA47ZrV1BzZ6HqPu5JDXQ+UY0/+3EOIVNq9jHDHHdq
MzlEd8OK5+WcgaIMG4Ny76Tav4AJStHLU/8PC4IXPhvxbOVgSOO2PONjdQiN/6dz
Fmpz4xWDF+t8Bgt5SL8oc3WmxqEoL6ORYOOFmtwZJrd5jtKyhb3eaD8RS3WE8R2Q
KbEbBeAq6qbJW/cdZKI9guhetOYCF7e0SU4Mn5sDRLqsFN5g5jUg6FjQnMDxLujq
/0qkQNfEmUrmWCQWuLaTubvqBkegdJ/g9/gu5z62rGyn0KOOHQVzbNUYOp0ikH2S
Zg7QUoUnWi9mnrsZmxYqut1hbRGJpTY/52NwKwrLky1qm0hFYhYM6UZGndUspWSO
thvKBhHqzzt+2Yz14o/L6Rs2aTbKDHIdHdX18yBHcxPQcWsddZ/czFU4wmd/jgNZ
fnbwH3zo7YrVr4A0RCHrPHAtwiDqx45tLrivYY3OsOBdUbP5CH8WaNzun0J+g6Ln
umLhu+VggMVC2I08RPncZ9e7aEnFziB1+OMx8ylxWu6YZXK2LBSsIDLd+lRDUeej
W/t5moUdEvCpkpRRE4VgOsz4AsMs4K8FGeGEgvcUAZomM2XppCCXzfwK1LsiGzBK
tLjekpMHa6qVDalm4rybDUGgyGGtTA4RRZH5ld8XaVupgBnevG9p/tzGlYNChZFP
7ArblS7KgHW3CTi/mh+tOw0vyRNUM7PBJoJyZvdHm10fmaf7xVz3fO5npjjdRXhM
tu4l8tHo8lVentfpaT+FNO30icOSHu5++I9qUspIYZTrLRmpe2k6jl1Bw+EDys6s
0c6dTyL4+ZZfij4JfybB5zn3E2dceA0Q8OKq5v6eQISs/6H7M6KV65dsQiqKt3kd
WZ+nihblXzkDIs/ELAOeCMuvq8t6hRIKSdsgoGHE0w7JmN0ztDIFy6/FpGsSIeew
EXkzL10kM5E2lrXs/CYFayME/E0e7ovi48ckdttYckjPbCFlwXzMtgr31kuA6Y3n
lel68lQUp8IlDEUEAC8VdvEHajXakkcMibBw0EAKHSM2ty9lMeFZS32Zl6IzUJnD
xsm3+g1prOibGZ/0d9oJ4szJcS2z8iBOtAmdm2wDo43gfDhdyyXKWhsANtuLRn50
h68wzJcIghdJLmEYw1fnWN4RygsBr+xflJRzTM7fazwBdZOZWMe365MbcLX7QB/7
rPAzZrcvVbC8nlrynFBiULKMExzwU0b9SCEFTaYfJ8KHTGw5PCSseRJVcQeVqooK
69G4cxZ60zre6l4C1Z9LFrUf+4A4FedNiTMXJnUGJakUm3F4MD7iI4u5JqC3COA9
16nbWxfOs7l5rmhzKW6PGU0xURvSjV9b42J1uhEm+eYShfjGEHLWbUoRXnJ9IOR9
sCjqjmRqI8M6WlxE6ns5RJp2iG7eC77TbQQI9GiE2AXy/DRKYrjY+IwXYX0Qs3jD
9XLkmU1fk1PgQBLZDMms/zgOZgWWcwkupLoQcFfDXyW+yIjm7lL2xe5cOh/z96A1
+qypH60bt3kMbl3QEhfAGgtycey1e74qVf6GFE8AkOEXw9viv3g9R438B0g4mIbD
zM5TMSUwPtqKd6vlrFfuhkFlT8g7VK/oG7356TB+vVizXx4csS5QyfUl7rax28fO
o4AimSeurChaoJSsqaTDlUQmU8xpSPA/mcmPlu2LMeAFe6ji3HSWexOB95IMa/vZ
SDq9ATliYZI/7yz7QR5YZpLdCOvSOcdnV/COZM+h4bgKs4+hJgYBoK7zSnctwVXX
tZdhlC3UaNh37Nq7EKD2JbjsnDaifz520VuyoZvo5Kmu23ntRYe1Yiw+P1+0fhW/
zG0DIl3EWXOP/+fLw/rjGNf9nNr6wwzqg2dos+qwDC52HBg1lodf/Mjs7st0g1ZV
tgSnmQRvxzpctXP2rtyX3A1WCTI4QzYLN5Eje/GnwKEsq07OpMxnkkonc1yTDQXO
XS1A01FCUHeSEwk5jgfcOIJhfVbMTT/NvN+p5VrfGEXvwdDv2OzDJs6IuCCepQcw
T3yqTHlEU0HSbmuvAWJg5KkeCa6alLrhyxwjqdM5anfmTK32ID8NWrjRu4NRf/Qi
WgAYUqqwWtVBmk19r2GoDqetR3pnDr1orDuWjpdQl1nmhxZUMZLmhyGFby+rAGYo
h0hj0MNxcOqGwcJrE1Jnglw1KTond5YWBmsK965oRRKBASU660VGLiptXy169+5N
ncy7enCoLiQ4ZZfJFrxXYRvVK8G3fJ58PVRZIWWC4ULZFKecXMrzyGX1YderD1zT
wlltEt0GvAiWQXX2rhCDZan9vPDsOushfLG2LLvMr/PkJkcE1VavP2EEDtgHdllh
mf4y+5jK6oQerAf8u52RL3CQWx0lEbAawxR7KTAxUht9JRCQvV6uz1F6ha2uI9iB
WUyAxWD+ljYWLDNWfYdqUUkgrh7SigPObb14DP/ZAoRsoRGwJOCqVLUkK0FOSlOb
414xN7+2zqpzRYuiUrconyQQDazupbd3+mQVG5xSVi40rFi8Vbb9zqbgVWpDU2WL
WPJXQUSEnEHjcOWlHDWzcbncYINmLQD1PB7vovltS0rYlh6a06MujwrPV1/5xL1q
uTxm8GvcmqPPGyp4ZfLaYwSM/ekMMgbSrsgtM9nne8HrLQd2+QR7WpquiOhddX6T
OSHUNXHpRhI4aqVlyu9pz30BrmU+TufqPOBCGk77MbbfCHk0wdNiGMg5SHeaIncL
FadYU+9pB4vcFxFLbP0NdWD54As3dPs7XgF4TexFM6YV2IC5ijiFOraug26vdNuu
C9mFeWruwXtZXMRUUxVbl+jCY4w/mRQxsRJ131jursVsWGRaEKkd5Rc4W3mRLrgR
ecweHV/JHB7zKOI/ucIn+cpbQfzXmUMD107s0Ll8yXdBBHm4qW+6LN+Evk/vfXgK
pGU8qxbNHYmchEEfowFlQ2v90rdew5OhXj4CCev/pFnvlHbh2xcHYLUb6lrKagKM
t+r7l/7qJqiBvWMXbvTqMYu1wrXK3l3+uaviaUI/qoaeNCCzBnoTu3HtQ/25B/zN
3rbrYVKhEdsm2cfuXozQR3Vc4X3Tsns1TzpLptlj2UfQqW7ksiwbA83FVp9WdhP4
lMwd76LAe9bnJqzV+mJX2cZltzZfnJC5X//HZZWYACtFyGrgbvncyQ4ksPh0LEe1
sBudXNuikgBAzLegHZqKIxOTP4uIn2QUip+CsOcGEid/GC+8yTClanROo8RQ5/pi
L3aYicEeNr94GlKSTQakyH/oJHf0wdYt4GsWSmoynWaZIsFFy1Ltim+w13cip7eO
sV072E89XHoORDpBpGMIWKTR+ULJBU8g7FV2KF1ym/b1TDoQA8uAO0B/F5MvngAv
U+qbjjuB/PPeI5sCWSAxJ2jnc5s8q6gce9DS7q072c673nCyznpmA7P11OyZD3gV
4G9qE8X0yR2UH36G1Gg171+LEVYDY0z6GawZ/7ORDLyGWkowGoSr30ZGggg3ESdr
qV08zWECoGY2CU433D49RTGQs84SOrGsqf6mJupfkmue9tc8Lx1r1CBwloQiZWPK
Chd9YRvAHMz4svdjgMfQnscnjLtcWxftyKmjJqKT7XpYThUjrHvEdQXKaHswKWj9
Ac4Jxk5wDceo4npgpsVS3pRZE7lRKiwi9vQSbC3TttPBKRGjpbrjy+DrjBIluLLU
WkxlM7WAm3r9ZhVsKnG5wT1OPxLXqOKowdi2xFUEOFhd/rbmxa3V19qUQhtFvmX0
zzjubGYjIw6YBUaohem9N4v9dvG94C2qE/kiV5DVrB76DFU4TahQRKPBOYFjqgVs
WSnWL3lwzi+x4IjJFB8Zonx4c6HL/N4iqb0kCSmSwHZPzxR8yOafTAkYwPUL67hX
n6aq3c0peTa56GXLa+FzB/eJb1m6M3YqJwnCAbeHF3mrYqnSzzLFSOs7CCM/S0Vm
Os20ph967uKd+ehC+bh7Z4ZUeqHPbRI86LRIfN5jB4gvpSucCvHkhStDkzO9zUeG
60pw2kl4ty9wpORlpgG2DsL+jZUpO5it2d6E9g6h4NrboOlb3zmyu2IqgdiY0RBT
4bqNOmv+4H12M3lJg2EDqwUmBFuDkx1sx7fB+H5OyeTbsZ4pW9gCT4KQcURPVQJc
NVvO7Eod0b+blE+OxayR5hwLkRrFtQoDZNpDKBbfDTdPswyDfLRVcggYMpDFct8P
qdyW1uD0OWuE8AMv33/unM1CbZMPeN5bbZb8anFc55bbHmmx1XR6tqdGs6eIISNC
ELrhMd1rzjPPQIhAzUMFy2C3O8YqQOaGc6muZakWqcpNJNtc5kixX/Qqt6iZSWNW
6kJPyFIG2X+IzNFKu87QzfoP0iCgSzsSD8KJM+HZfCG/MDlfQ34nfTs5unczrpl5
vIAO+Z2SYcO/gz4GDXz3fyOT1hxOy6R8NpX2NXpuZlf1qFgYvSaxNp68ylkb7WxX
eWxHytJRdVx+FiZC+UKVsHnTQEpYHiHl95/1FQnK8J4Q1CEQ2GfYsHLE4pbBbGwk
fYqSr2Qn8+/20yCwebajwokzK51viFT+ag+Ls8ubSwcOOtP0d0R+y6FjqAcu7gER
QYVRUSpKbG1MPYoIkFh4jDLKMP6FBxxmlqlIcJQpqjA8Bx+CDLPJKOKIw/zOdH+K
XIZvvEIOuVLATzqKWF2+rRlOm6yISBfj4jxgbaKC+5jLeNTLFX2r7zfKg4WWTOrU
sklyG1eU+8Un5+Zf0svQa5AHcOuzsk9DttKV3acsUXHU0Nb+FgVpZcU8rkm80pZI
WCXplU3IMv6QhwWpHQ5CDHro9P9vFkvBPtVP5Cf7rS2cVFVZVT0+8P6mPYZ3NBV7
njAO0qBgOrFFCITH1BvE3YaAQVjGtswiTnQaD+rQBoNaV0t63E7xf9hftnST62Nj
IPMSD4RtkbBqq4PO+cQZ0u++8y36FwW0ULrHsBONiYg5kh3oKehapR0sFz9FFmSD
hrsdr2/qPjW2SMHf/sP2AwxPJ+Avg0zwwTAWa9FxaJ2XcOvILxRiJzIi/BcDkpqT
epAGap0EdLefUWGOc2kg9qk1R2gBjLAUk7fgHxiLQ72cJzhRZC7+FXRXkilrUfwS
B6D4OxueBj7QsYxxQV67KibGgzX3NvGVHVpaxWDe0qMPBPMatSxlsmYVTUz7Roax
ifpiMujJkmA4ypEy6kSF0xjRF5oxFnWEYkwIqUGCaJlVdZpsuAIWS/JFu39bttzF
liYpqtwd+I4mmLeGZQFyarMoyhWMRl66DdL/z5CJp73sVlHrVms9LZfRuwQHHncW
1dSBoy0EZ7G/F6trteC47zwjbO7mrEcL0qLspvgdmtajM05VE9cS4GFCrG3M08/P
Q/h/1ZZQr+lqwAzSqRdZrDcu8SQ6eoFzqMlfWZK6gFPmmjRhtMEOIod3Tlx7LD/H
lTUpRvyfdSBGG0ktSfF5KHANASVmKfvEkArPAVpAOYW3WsfeeGmzYOSH8talUDRa
RUPg2ZMUwkYrJaVZgMcUrJJ5lH6z2lj8gVnwutvUT0brHpAow87lvsRuMSoeBbr6
oETulP0Pa05TU8PQ//m+s/ndi4uKHZW/LZq3MWncX9QHJ6Fg5OXKonxBktNOfLWa
0+3BYXxJ2QlNVrYm3sNPDGaoaEUhbDf2tV8mZD22pMLSHdS0v5d+oFzclJ99+U4h
eXPoBJVX5eV+sia1XB8UOpDx3bzjYi2cWrEFp6f3sawCnNynaQf3f5oUjKyhyoyP
uxn8KEE9si9AX8hQ3ky9HFbGcH5oXGqqJCS6AbbbFOTMK4vmHfWoaSf9iRWNtIzs
coVtnozw3RRL3+d4rpT7PRHvC/tNoRSB3avYxaKPpfl9mZ7ACXvs8PnSFpHoXdCs
Q4A3GzseMF1/rtgo/Psk8Z8BItTS8++Wq8nFVrAfyew3JOyPz2kuqYzA3UjiTPc/
IJ+33iFnw3Y5Jx1vxHksmmzdt7MjI5WTmPzV5tMBoRNRp+V1XRPS71JD1mXBXclZ
KI60HgL33vXYM5U62rM85vkta48w/GdpqOnySf3A/Uy3N8pjezVIExZuyQTYIc7R
RahROGj+JCP+NPH2Slo6ZbWWs2ATb95LcKlkCZ4asniWLxAgWUxWUGo2ATE51sH+
3YasHAiOD11Kv1XsJdG9JKjAaaZAvmP49BSjWDUsxpNRMDRDOCTpCGHV+2FZGgr4
usXqfenkZESOZoKNMxXzIzWIAicxND7xBd7r/M4++Mid4ml1MgUY8x+nO3iCCYN2
1FJQsZVChBM0uEjsKJm2IdwRucPbE/A80R+w2uxdM170ItEVqj3OJUistuleNdKM
bEeITB3EzYeKGRT26l+EZKL0wd7p24iim6qGJcSkTktRqToZ0g5zGNS+0BoN8fG2
/LDFaNpx/sbIEFESz8zgQHd23GlF65pcssfSLKHXw3AUd5/xqQQ59bEMZxk8nsQg
zc7OgLPpfCwQDpCBw6HVUFG+PpHETNSX/4FS6oBrNo/N/0O6exf7SCdllwtKFj5L
cV36y/QXKZElJ3rX7JxnYyQrbHYyGqnpWbc/aNDOLIe1+ax0or9n2hmExsgPrSRC
8e+KRhs4/pQ9QqH3uixyYF9wMstSqUE5b5GecPzaZiSzJEt3axK1roIOlpn9Zxk0
iMRDblEuyJCkqV6KwoBj8u3zQbEkSJo+OUrj5noQLVIUAqUKAZnEztH1y9bS2OmU
Oo3wsCCmW0e10BrT7ueDkxH8/k9OnwV2KcD4PcEJtnNGfV8tUv5HhnNE+pHpf2Qt
ctaCrAM6EdgzXqZFpEA/ZlYEvP9rU2qhL8KBxiOMhVF2AX+EIH2Gg9Myeg8wOZ5X
NdNXZU0dwrXQljPAQPWu7mGiAVkqF3G2DMCmycHPLINERWv3f0tTNHQ1kiFHK0wK
pUgbY2mk7eEyK6rY/420TQTGupq7jv8g/5Xuv3173zr/i0+jRIHAgUzNcDszSnek
50N4wWbuqg1yGaZZV5wLFYacPQespRxUIrqWtAQ8nuAtNShCRfCkOCpPeFoR5AtC
E29w6/MtQTVGcASd2WKLajZDXaEokUSt0C2KcgnUrAT5Cb3J3Ll84tv3hLw09rix
C2BzoW1EZBM/PunwS33dvA9ljg7ZY4gDpCv1KQLIbPvdvsDAesZYJvZCbGtTCIXz
v8kU3fKIeMeHzd7aJVxiOCmp0JK6W/3q5oUrBySDMVFjxFty73l6F8GBTah1z4j0
x6Hkd9S2E6NO6AEHrNugEx6MuWtWQ+szCWojUep0DFwaF7m2exTvs6BcmnnhfG5j
B3yjlaqkZ8Aqgx5l2iBRfyAzmfUCmSeqfOaBRzfJzCsIyD2ydAvCSq5R5tWAnA9q
E+KMBPb4Udd8totLARyNsU7rstbX4GHKtFXkDZTUT7CH1KRUnkAoRjIdsRcTOmcH
SnX1GlVq5gji6eZvyDMVxUMkQmWlwi128nxIUsOWXLlscz6TJliNWvVSxnjfy2nb
i9d79PqEjUlzwQ2tLw6xKAvlc5VsOaNl5lO3oruEsPlo3egMb+tMZMigl7dj5BYn
H+KeO2PtH34N/vE14WLZhVlq5w48dAfRxLngxuNixEtMhRBc8oT+fhOrNwBWEA1I
nRgsuPkCYPdXDemPnnuzO7UxeQsblgH4WzbCkKmRTrp3hvDgKfldg30vdkMT1Aqh
hhxqwfSxKK/zKG5p89/GNUgOS0RaIkaCeSwqZKzLiyzESoZMFb+nu+oEk5KDz9V1
UtIENfDHTNtu64I9lWT23ZtuVIL5nc0BlJBUlxBxUN2IKe8yU0O0B2fPAhHs2usf
k3sg6lUpSD7u3+bnonwPHIz2R8qVUGo2dolBQMpHA7kndx4eQPfuErU/VVM2NBSR
oQZs3+3hgI49EB/j7YYKPS1Xi8tX0ML0k+bmtD12yRhctqj6CZrcy0IK+JcxTQH/
UWEU9hKU5NV0BW/eccEEf+jLS6PzQPt4sZeyxphH1goDWHZ8WfECaw2NsA45YUIu
M5ypFXUplsn7Mc4CA2+u9GPSjBdl6GUxpQOhPw9j9P1A59z7KJapgwbF5tHxnSnL
1dmhVe2jtNn6uoU4o+9cGKAy4dhbtvLfQWN1+a3By4pbBcIQWKFSvAoAZx7RJ6EG
CekbISpMJaCjeSDdkmaOa1HdzR80XAj0KQqNFHans33uvXhwHl5jI7ehcSHJkzij
qnYwDAszg8yLirRLxl58+tzCwIk36Q+StIukf2VCaMnGzsHv1CNtmwV7hzitFfIm
QmdphYIG6eAi+xwJkXUgN36+AFP5LIsy0Vdqc4d2jtwKBhRrRFCpW4W7ISXx3NiG
uDBaaFOVoz0n0P+bbno/cuSqxUlpSbelKeNCErSSop72+7rLx5qzQTkZYMMEEiag
PZUT7qO6juEcWEIXw513pA2k6/2oUQOxseqfT+5IkvGhY476kMqLZF3jmB5huNGI
qfalQolbz1fmOr4GCMIsKXLkGc6IpIGHy4y3gHGmPdZs7RFQxUh9+dV9meekG+Eo
pW2ayy/tI2iMohjtAtH1PgnIdOWwkSBd2OUasUQniclvT0kMZib25jhKpajh3AWL
fgZAU8W2U/RfuHd+l2T7YE2LqhpU9yEwU8I9IbU8UZiwLW0PZX5j4Sh5R6yTWgM+
4qRDlHZNKzyQC4lm37iRngaxvCeLrRlaXUwPeCcWH/IbMZrAWYKk3n/bJ7jFWwOk
ekSgVDlGku7GN+pEUaXOllWNu6PyAVLqyPH67KJCJ1/EL2Uw0+HVUZckFjn526pP
wLUFAwU7eYnuMmYcCaYSQeDn3SVmFm2oU8ys9FBuMM+y/ld8b+poofC5lI9Ktnwn
VDHvqqm1V6G4Hjkkm5moy/G+cQTDjp4VersZQdebrKGs55Gw7/OAr0CUuc3QbtNB
n8Hp8HtQ5LeWtwr2U2EJ37+Aydr2icWPKsZZpBew2mKBwJPULBIHJ5rMrojZaXZr
YlSvXEfW+dV9lGsq+mNPMhCzABOTE8x3ZjTC595W1pAVRvQUxu1FUUjnXWlRvhM5
9aUP8dEtQ221/TXy/w4bbhl+1SDcUJPpzKN/LWmzLICr2OI61VSS01nyZnGXk23h
jJOZ1zDQpMq5QhbP/BgQmyrLD9CGhtsV4nFLsXg7lZ3uXgPywppo9epT+t0Nw3Q/
D63mzXztzLo/AEkMn2NHoR86f+pKoo/6YNZrm8pShsz4SCk/DIj9pkV5I4Xwe8f4
TdgEG4EA3istJSHwZY1iQKbGp7b6uvDHZNwKNzntFdbjKcrDoJX2lyD6H2YFVCW4
pVjy8/hNLbMqv2Q944kNF6vEumNTYjvhoCPezQPU4uYPmO8H3lABmX6GTT7qDuWA
RhuwZOCarmTz3ABKd4DIxAGduBOyyHsEdsTHj8liIyRkJzqpxTWgdIkxzXCYWfL7
doticEYxnNON1A1j0ulP2alF/kGYMESqyxv3EAD4fR7T0tP1zVMLAyqMiPQMueBj
Q1cFLLQQmx3mos2qKprL9DZJmUAzlkC/HjbCuuKoSa1QTHFQ6VN3xlQQMfZZMK8J
mqhWUiDkCBPTbM0YOzJzTBaavZmZ4BS1GqvEEBGu0kP1oJj1kPfAw/qBPODN3BoR
w7lJDrYvzizYy/ue7hPduTzFiKvdp88/9Y3eCR6++EtLw7GqS4a/0fkSVdFrrk6E
L+RjrkuHZXs5TXjgah7zXiOU3AWKw6bBx0l1Xb2IC99l55mNBkKWQX5+6tYOAzIu
oyUwJ7guDflaIi6U54qxRRmPrtEjGOYDXxbBkwPgrhERAHZeoUva2UXtYa1axzUq
MsIiWZ6UyZtC/zxWBrYH4f1L0I5Vw4nqqzJ1ayH+m+02P0Fm6ojfcVbEQR2WCqpZ
g8gPPNNL/42VebUZsu5e8kFukQhn9QkpEDXZVMIgi5K/c4fngqoTjdfllRvWHDG4
moLiSl0GgM+mEUe94fJXszu6PBWJRwSAlPXzh4xqwBq8B+qdx0dDIZXH9kf8CjfE
14I+ZhY1jFhKG8H0lcznIqGJh0dnSNLRbeM68VLj6FXqOm6EL255bzpkZlib2qYU
nboXv6hEP5HMpQiTZrpGzWqgbSzlS+BRalKee7tubti0K4sgErVJq4bDccxt0am8
+oRY8o7pgcXUpXk65OcLnFkhopv2J9t1xL9PwIdWEybmLLOT1sr4vlj/kgPU6aG+
cILN84EP6CP4Xrpw3OoQrOShYZqgQEF1fVSsrypyEXKRsy3LeW83GdVkcoyb/i0N
SCRKNFgZd76f5xlg4mj3f6K0G/aTOtr4HMyI9/SbbQ3zZpR9yoiYsGWe6jdLPILx
pjS8tb4L7rTybO8dz50OiAGMCpJ9t02mfrBhUqJyxAWr3s3ekDGyzbGXB4WN5+jn
1zwBLEla+P9NM701WQEmwoiC3q64L+yVev08ALQFeWZBkQI2+bERBvyrZwMkuSpK
KgI3M8Oy+LWtjLYOg3snBmm0Vy2XPqJcJvh9brWQioeK+G50XKqtfxFIxrqvxjdx
ksOaDslBdioCS+NT0JTcsdUmf/SfIzd6qAzhBf+5v+GatHPcAxVSM/OwJh3IhVNj
iLBZGpRQNVF/pD998aR/807yk2AJJTuycKxUXEGt4raB5UNVmClxDO1bNVndnIZ3
yqhqMR0X42zS/GaUKgPAcVbMzUqKTfPJ9mhNa1Oe+ykcv98nqrei41Fsn2aWBHxu
xTTesx3j/lRUfr7y1StuyuKrxCztHRQJV8jz/AmUcTaVydDyKZsh5PWG1RRFSD07
OcVMzOjSzCqu55oQG7EZITgVW87SXu69Vk3EnjNMi/KqMz6iUjUkGQqc5lkxkKL0
ZU+owrHAgppvHLID3e5IzsuTbrj4sNg4MY9wOjj1r9RhIdpSVCA5FRrk17Fuj9th
76rLwJSol7C0QkYygAkDYiYIxwSF8PKWO4Lx/X9aBGx7J7X9VT/nIgeCKqI4GSNf
FGQLL5Y79n2rS1cFzDZx8Mo0S679fBG2cInQH8b1dKwl3ts6ieahk36Lc/J3gOSU
9r/HykSSLpTuUWXYHkmcdcOCRyUh/4M2A+/pNa38qx/QiUc7ih2m+DIbk604rRRN
W0REKTbkgGrFB1IWFhC47uaIJhBbHLnXvJC0ftY6aqqRWwS8aHvOdflW1em3N/7S
NTng85gVSqwv4V9rZiovVCJkRRBfVborOLNlWrcaD/GC6ph+8XpMeKsbiBqfYGBg
j4Rh++fMa7a5qvX5FtiYJhZL+5VdLCpbV4uc+AfWA4fhog59E0mxYUQm7OWvpX53
PeVlKIN5vngdx4bpqVxdZyewynG9JgWlvx5ayW2si+KPGt+GuMTUvb8IB0trRBSb
VOQ6ST50ML+nB9CoeOc2A+szfAT7PKsNJYhQH8CsKaj6xPLJoeJD0vZDk1OsRQr8
A+KtCcDD8t1zDv/XK/a1kb4kH8xXj2QFTkbJ6JxRQXfNcaI98gMW9USjP7S4a1ap
q3sk4WT9P4JCHgpjGVDf+swilz9R08TkO6G3382rorgGVq0z7XAZrhkLWYQqMocn
EQoPBngE+VbVZQ/w33GytScsZ7EQYWJJ3Fn3O0HGG7DIIqARzgOVdtpIFSH4myFv
W+Q9vDVJ5miElIgm7+HxGZ6/oSXz1dCpTNUKkW7Mtfkj0uLcaBZbRzl2wGQe5IeH
lIDr9ge25VLM+lSvLFM29Avkp/s8LJOI2lXFOVSqMSdEycSEdP9M5nYqP3Dh3Ecw
Ln9wH+l5ZQGq144srb3lvAlWtRaLx1pxZII37QRFeGO97m2S6cDN6YFvUL7Wb5GL
vDSQKu/fuAFvTKkye4vyc4Dh1JEwxr8pCbgCdXf3YRhXSa0n4q4FVTpaa3mmDFNX
9tcRRTZahBd1dI7yhcvnfR+qinlfNsvItsLl5vYbqKhAC+1RprCgvFyaln+uBqtl
I/Pk0a/N3HdHksLaF1Nepk2kS4oqpo8QhRrEyYejFXzo8O3AgrPnX4iS3I50WIYT
7ahgjXnUlvtPlOZ4GijDUk0wGLtQlQGfOSyeDzEJrn/3XB+FN0rxZPHW1F2CR9LK
9TmG64/kPI1sCglBTaiFJDMoiP07+wAmSzvGjbgK9QhkLL3fEP5Cys/XhqHkBQjb
AERaB9P1h6rB4GYTUFHuX0aIbB9UxwYIiAJe+DqEYPydiBqdiyR+VejHfxVARvek
EEEJNFYAZREMO6kRqePPDtcrHt7Z8jDdDUeDx58rYSAC+e01eq5q95DUnolOoH0P
qWUj+K3nQ6VJD3NLy3ke9+QT17vku3XIiMmEm0EXuNktseCR25AaZ6skfABS74fj
zXMp0AMMjyOZAyEevwNRxsvIYuwB8xDVOLDDM+lDDzVoYqt3r++Xods5hafusXAJ
jKpyjosIBf5Th/BTRGsJuD1XMp1b7p4UbsK8qaO+w53d1eqDmzWRE9gqL9ciY3lK
wpHUWShHQmgnuu6ljHMOsDwiFWrhryAb/w1ZXx9S8n2VFatBxqVYPNJSpboh829f
lDGCjzNR/MKCC1jmoni0ZVOhdFsC/bwoi7tzFNi9AUnmDqzq4JTzE2xXFaPNsgZC
Esc2hq1+4F4gZBPpgXrOnyH6GMln7QSQ3i+eWhDILxRBG5kYw6G37fZKxDDl4+/U
bByPTYfTS0VbcIxNqhBDYLnNweFmjDxAeuBw38OgL6sXd3fvgJSUkU6ZxMgzD6m+
/5UWM3jIsxl6cnZlJR57FAAfTRrnELofs7LNdAkxG9/IKCmx7p8nWP37rjcgrrNA
Cif/6lZoMPMf13v05BSOOiromQ9IHw3+UlE4Sy35X9IbJHHxHAe+taFmnY8c3Pyl
mPhFdo5O0ZGmiod32FlplCSdDTd2gheLmjfvCeveeF00PsowdrIl4PDNpf9MuexO
AyVq46GmFSyb0uOeUCOwe878KYd1IqRX+2K2U5MAQ29a8TDt70LLDmvc8KKQ59j+
GUILgIs+zDAB3XkDn/uSBE9BxDh1s3LvPbk2nCcO4mIkRz8lzA/UE0EVKPvLeljE
ji/nG+00x2V0IhWOZpiF7iAdIX9rrEW5bV/gM/6OfXFMRkv1/+CibQpa9MhvaFDq
8JOtJ/Q2ujsCQeZkp9rL0UgFWrxHg14Hce1eez5xVouwZoPX/C1NMzlstYKvjq5N
vmjfmmWgYv6ROm7qAV7uqyJqA09h9axE4I+WxYuQmJ9YBWRGgNSKzhUketzN1pfZ
NIwWkhm0Bc0HQK8/m95GQt/SM6D1/C9wIFnmJKmcNupVIejqiaYpRXU9YMkz3lDa
bkKECMc9FL6rX5FJDGx3oWyHQiH3zn2yAI63E+S6DtU1PleAG+3Nu+AlrcV9ol9R
PCYMTJE/Bao9X+TLbhkwV2UEqhrdAjGTeUOJ/dunLGcnbQRlsSjAK3WZlI/XdWtx
6zIDkdxUCmV6GwL2JCPrJ4UHBY77VdXw9+ffApyG0wPEt1AU4DKbDHrfvtjAi5Gu
cxQd7P5hvdVKIMGAsDynncDG2RUCvNr9SQfx8JbQco1Qm2DMIdup3H3VW0bCLsQO
+RCGdNLb8IueoKmhQPBv+rmnm9ygA8Y7oJgjbr2rYdaMNhrLWdfzeQk7nIhgEb0n
P5QHwcM/cQvXllRIZSU/rpAj9ms2Ii7czEIXd0I9sqwJPzIRJZUVwwAlUntsUOIa
7wSXQOi+Tmbi9sWZOTj/wm5w5xMTApP0Ilj/jgn5fDJAiSVbfLgB5yrXJhCVZSk6
5Y7FKj/ToZat/7ZzY8AbqKAwtrf9R0fNj9JtrFggWG6+lLVq/RreVpMT6ly+B/Co
m83Pvws+ZH3NQCxhGg416e4pUfbl8H9+oNijwvU8tJY4NAFYxcHKwswaYAyDIJaS
nNYudxK/RnVn/3i2zCi2JLJgCWg9WIvh3BFF97y9U470TEpRybYPz5jEAiqmeoLy
YCkIUIs7XJziXPHDOXHIuSwUleR3PeCrarvoTkGg8kS7v8mO6jWBLZrz0qN881o+
aEqPG4ksmEv+AfTqUYrqVbNo3HR+W8QPDMbz3GnaTM74SRkgmh+5NKIYAGRxbb0J
OHkxAeEg44brF0ltC6s7WRCHp7ily1yzg2w3OqCP0swIHMI06XgoPtG9DhHjhvS7
HsgkkDTENUNZp+AD3PQ9YZGt1WFckdY8XVs1Ym5t9LpZKn2b1GzA9zlFk3RLKlA+
iV2nwPetFO0nVDAgS5da6xbHNq7wxl4DUu6Ji4GVxMjJayCuj04gJ057p6IdMNMN
5VEYyyCGAKL+/o+Tb0oNeSRotlHAyvjhdwtZpwkrde6bG92TFiS0qUqmlMJSUiPk
vJSb/UHHCcNaIPCUrag6mmf0h5/rbmtE9fAUfBI5VpNQhwtpZAMHG2eHyWnFYO4a
m1F0yXPFHzPcNYk+ovzBOBnzx/eivxuI7Oh8h+r5LZjcWHVtIdB6UbOMD9RwqFhO
wFccbeMig47V5yO/7NtpBD8wHPtEZkGjUP8+I3SEuexlE7580k3C3BfOEWIBV69B
k7ISVbM6kVcZgRonnhOZr9BHugEM6vga0cd20TyfTCeetC9dTSaVBFRrnU9O0ulM
bxdE7PzxENv9m+Im+vV+Y1kyVNlV8LUxgFhkYTrqFFDk0Inbq9F5lMIGNRdo7sQn
IHRTg0fFoccSNW2Tv7zI9oTf7u0dewgcYv3a9ieECGCvKzGqhezIrrYCeGptpjPn
0+0fXlnSFsMAoalBuZF2KB1tWyj9rhCMJm5+rE78jaQ3y0Y4DOAG3Dy1JogyOk1d
z65xPVwKcpt51MiQMTmpXCobvSU7D9uCSYtge90L8q/t6JfNx0JK0Ei8B8hAWGGB
UNvjK/ynRlOEHB7EDb6YYq0TrL09JFwvHE28EwF7vKfAdtRmgp6NOoBiT2I32Q9R
O/0l6FyDV+8/rT0dY/6BUzgz92Y67qX+Kb0WGWT88tQYZebQWLdmTGqC3J98OLtD
Wj0XZ6wJDUW4IOnk9eq5di/aWmWACxGEQPtprULsJUJDz/AReRdE5qyoFY+OJqVn
78zYWTnq9VHOpFri0bN4IYQri0S6tkOFBoore9/1uc+EBLjtzXwyXKhUvaWUviM2
69L8zftw5fufUC8YofPp1nmyyf7QK/rWP7B5RjsEXpGgXSKFL75X3kwoQ8YExjGD
Lqp9ks8mByP4z+3uKQXtPTJttrTX49O2buV6Aw/Fa6eBJMF7lKnLQJed6WerSJuA
ywWgUlkGoCuE32KSzBM017NiVVaohjWe1xy17T7HtA7rdV5XZx1W6aRJN9rCyMQH
Rj3/iGtiEJZrsW0sazdhWF7EqX0/BmEmi3dbWdQBgLnA4XGu3oBWBw0j5bUnDvOx
1q8djIhI6VCNcDZAm+qP07LY972PJiRu5KdfEUvYyWSm1VtilFjosA3L2UMMPtNV
P0rg+silDZmJ1STaUOn/iYMCekgoozWtFSgUoDLPvG+agf3W420hGUPIcmYMLt3Y
FP3LFIBcHIQyfVtNHhfs1rNPwMvLPcFHdM7C1+lW9dEOzIYU1MTuzeThZTrvg11K
vImQZxm2g92abkkdGg19C4RpIq54DQb4ecgYdZpxlxnVovNiUuX2+ncZDEnCY585
Xh6Zl5wdLLLx6BnUbL3VE7VmtXX0kQs4mtiMm3e4H4oXem9E/aKJ9RyJ5jQc68B8
omSFxz91kq61LhX4su3kvIv1ufmeEOKNUU9WOhXzDyjk6gFY2yBBS2FXC7jwu979
ORo4O6uaNseba9S0VYYnknRXd92U+TKlIzYms8Ukg8UCljxJT1gHWALMC9Uyt7M8
fB/I/ZlrrMMuERw/2TrVZp+EF0hEgr5SU8rxRBcBjzJtZWhqVzb++PtyaBvHOJi0
r3Kpz6dreZDT+aV1VONEzD4rjoDKB6qx+voxktJ1AQ07J/0vK0ka+fltkYIx5pzT
espFMgnCsTDF3PoaJT+q1MkmEPTtIpBz13/PFZ3rHvz5ZDQvp+dDguq99BefnaDQ
RLJr/0hPxjsxGUE1cb7klDxPS7e89m60CkT2BBzS3zSYGr74fj8BzLkuvRY57iUQ
6Unbb30pNLBNw9N2gLznEB8he1DjRg4hQB4xrJY6y5b7DuzgPWLiMZ46WfqTQARs
DmZRTz+1H5I0+W7qOxg0RUPi2aMP/yNjJYGjzjEQpTdYdSR61xZHHsJ4z2DpFVX/
E+owRi4caugF+RPr6dxo68ivA9g/LqFPwhW2nVpxj8V5zhDGZgQ+EnY2n8GS59s4
bf04cHqYYGGZqiW2dNSNhaFCD0UF4nGDxxNwmux+PfQ04GWwrHcm8efhUg78CDFD
Zm8KBqsLSjVaa7S3hDqCMPxexiqLSetfFS9hha0UcBGW5MjzH4NccTgniFIngA+s
HnygDLpLEvmhRkv2RSeXUJ/4930l+lECBK6VPeWOKWKdbJ9vIYuG62qkSkhBbjkG
F1mN8gvBEBmz9m+ViqC4g63Wge615cBQJtQ06j/c+7rJxOJHkxcieuoU9zXKuqTO
ctKC2mM7ih+iLVHbYONv3L8uECnm0PTkhyBRT5YQE1QseGzwwWWKRvtvTlu8j+O2
Uq/7B4FuYyhpkjxDUolEmKyI6+dG5tvtW+pWOrBLWzNS9e1s/EJ1ZTUK3dpVjizv
MS4KOBv7FfRpltLREXsAmsxsySRyrfxkAHS/6m0gegepEXHuvZNcBL4XiUF4c/DH
XSJo0yvvyTHkP/bMgYSyYKruxg791kGedlsAqrmHsl47zs00x/feBbe5sGLLaGh7
TTpKxm4Dr4/dpmiF4vFzOo9h8HUpSh1dmL4CGD5ek973AVjZvp05JvayRAPAD0NP
tqqMO6dRZ38G2qsbxV2aWMt2cUdiaT8YogDjq423KXKLcBJlvuGYri5wGZ+z/1pG
/yldlo3O/2abdb7C6/vP7YE3LVoHza/o4iVn7Y3iVg4k85ius+MXuccQA7kK8FHj
EGPEv+rZP0wRzd235rqnX/4OueIZZuA1B58WvcNkGwythjGJuogINp+hMRUVPnLy
94qJmYqPoxmejoT0Zu2vfBAglxjeeQTgI0nsxmIahQIUBL04tMsGp+3uu53LOvcq
apKbz3GOg7UPdPfjzsTyQs2BTQsC7XyXWw54JiugWfNgfJrg0IELc64nGF8uYN4/
NFq9eC2zuzMY1Hpi6SVaz4ewak2pcB6MJm8zpnzcMW3L31nrtm8F9j7iB4ZRhBpo
rJNxyN1ltQmnd6kfIuTLiYhavsKwSF5UHYtDb91LERpSlT/1ruMVo4sjXOgUoexP
MK/FIa17cHtaRwqdO22F2O0aus+ftpii6gXPLRG/XCMvNi+69YhwZgdATP25yrMq
vS0PCXKplXKi6R4rMjZPXjKL2gLXstGf6cB/JnAtBiF67zd84E3lH5Xo4Dx8RvLl
pRUkY4yznPpJMJu6vsZa33EOIdZmWVKlNQZ30Bg3q82XaIl3Avlv1otSqOa0S64t
bk+zXhFVuypuLiMDDeQ1Yw0skQ508/JnEHRy6ELdKX0W0Q/DpQzlbcV39cbEe+0s
r/T9OwyBYIQrtE4UFehqhhOavXgKLpba6RUwJOvhOLNrWwNPYQ8SZej3YpSsFb6Z
hwpI5sooL5RG3XMkR3O9bc769QYyA3QcjZFRq9rvloe6sFmoILtl/WHzbFrxcQv0
5b0leMJFXibY2K50BtYPaHdZr9DrnRU6DpfMT6IMzkl+i0koXVL992wfZaLhHLSu
sus+S3Gr50Q4LoafEBr1bzZaZoMqexGShinguRLRs19iaAfdKNMoLexGm10KaVEr
rdviRLdw7VcSDytWXzzm9g5Ijf4Is2/O9gC7NTcJ9X5pC3wZxJ1uLNCpbgJTde+1
b6Y4V30yjCV9hBbhqMemDdbNuoPFHTCbacvAY8PCtveWoGnQh4ZMsOK3ar/dqZqQ
h966XNBw7Yd0DnhE2EWV0e6pR7xEegFQAksSXv6IlGIfOnvV10V2Jcea1TGdwaTD
Q/tyFQseFz5wUQrWAoQT9gegRn1JDCB/CD4SeAabdNKjl7ynSx4WUls82Gn7GbuX
BhCcQu5CUtJld6oarkTN8ghf7pwCMOaJtpY4C+rfkY6zmT/64qwM2Zv7X+NKQDZp
/AyMEp7C2rbY0E2GSk4XezrcZMfJ/Qv9+RcxJxYGdfGw7xKuPToyMwF2Khm5p2EL
vyw1/dYV0eLnuAdp0CKtvVRhe3nodfBIfbnSfKxWuCOgH++Sjc70saUO4V9DX1BD
H49qnzFB4u/b/Bm3GAn7yF6zwNtjle8+0xQTLQJQDqKZ/lBzMuamSXXJlGqCIFHj
Dtp6ag8KYfvjtJeNF4htMNSHv7FrNwqhIqBWfdq6hRoPaIYQHZydfRDXRdWqNRPJ
nwATJ/LtoCGU2sMKyO6Uu3bZ2lIqBLhoMurMSOevGDq8vxJqWKSkJ161iksLvEIP
fwo3wjOTcgDNVbjUtxi8qHTOaW5bQBs41g10ftSHYG0ekYhoMrg5iryV8uFQ41XH
uVudXk6hWQCbHc5D+g+01o0UH+i0N3QJTRYI+7LDRY5K30adI+farAPGX/+FhOSQ
MK32LEOyXHgQ2H16hi5CgDRp/K7/aPHa1l6eD5weq9mx/awbp1mgs5Gb0YbmXLeO
2cZoVWZ4sSqVx/nz+cxgNjiYdqpSLOPkE+LOkEWggw7GihqOesm5liEyk98GQnTC
Q+rAcCdn/IujUj9CFI6MAUjn7IQquBhJGiAwsfGrqDPd1a/JXG55+6S7MYNTPmYR
NPPvzB8+vYKQGWMtBPNr8lDWs79SMV3Dgb7wXWNEIaB6GhZqdaFb2iU/SG4gfF+k
ZCAxs78uOxZnb5QDYa8/7pb4yE/Z1pEbjDe7L6qX2i/Uy7jRDgo38QGbrKuIPFSq
zFkni88fCPeM9NubSVOruDlR/dLKQV6bvKHyYDwseek71up4RJadaMQaGO97S/cZ
dIL/oCVHuyOzt9YMZeVN2lsw/6Rn1KHQY3KYfDnH/+/G19FAC5s6378E9Vqvo2NY
YVy0maQko8TprGA3HCH5yoX1jglSfubxS8JP6Deyk2sFNsAgOSn3I7ZFD49h+rfV
vwzl/WfzjNXXALx7IXA90qeqb59TV88udNA5reurK/1d4TCiuWq/WxfHJ2gFB5u/
d0dEGXfX6ThDim9DpJSa3iY8fzIZuIPZddqOkqu/Oiv/byjOgjnzLCIeYrqYsKSR
RcvCs64tKegU/Emyp/qAdOEiv2+Chh38tyhlP3s8nHYZzi7pxm7pY35odXFdIvLU
ceis3A/6eoRUWNjKkfnS+c5ghI23Xhck/20IlhHz86TP2N0z8Jo4Gh2TFAygmsx0
Z9vNY7PdPSo883xmxjflf9Zims7RJkTYYQe5BaT1IJ6RgMzcH9CuC1/wi1J6+wOP
IC+8hlhlv6tzvrOPqZe6GrAc+NrpLCiNEJ88ivonf7s6hCtcWoCzvMn/yyOGLIMo
rQekQ4szJy+GIhkBP80lj1NAASDLHP+M9oFJnSpe0uVVbouE1jWzgLjF7hopdFQO
xKsLCQL0aAbd+It52XKZOH3cH2qutO/Yb8OR6ew6oveeEX5cxUPwn00Pmmo9gl2N
o1eKU9ANg8Ej9FEx9wxJRUa6nQynmjFFYu/Sc2C9ASA36SurL079GxIPTzrqG8my
jM97IML7tr/Rfe+VApPxjI3xDP0e+ap0W+YMecsFbT1QZpFBPvBo0QJ4rJvLI/BB
FmFsIB5+VzawJyEYtmo7q4ei1pucc26MPZZ4f+CpGzfI7noyKzX6B3dO+eyRiaym
OfCpMT2Im5OuMY7NUQk0Pa/357B4tr4xnMz+2e6O/TtH3PqgnB9OG2DU1qEtA0ex
z7rsi60aYsZfQ6I87jXNzwAkj1bbrbuOe49TZMWuR9hfJkIIP0oaI11XOHWya3C8
hQYlqAXWgWNKDCwcWMiwmEiYoNHt8/qm79+N764T0biTlfGzJXRoTN55OqfZLCSW
466Hs1Pi97wnTpAJXMYZ8yTKI2oLtKRJI+2efq++YPNLP7YJrycdYa/OxLnt/wKr
kdNhohBAJXPJ972p2/2IOU6S4oUa+oGyX/1xZW8XBN6jYpTn0z6Egl5ZKvVDo5Yh
uLxWCmkBLsVy6DM7I5jPZrl7tQ/JTx12QX1BMzz6Deo72f/XQxeLD6DZkXWkP8qa
a3rJ3mFQ8cTyxD9rlQpAeOw12XtlpqmKSl4lLhfk1sBs5ZAypZ1znqsM8Z/AI5ze
sJ+Bg9zh283j5XyOwNHBt11p9rcKoFVmE8Ds3/qUwMLDyE8sE1UDB8vwjJ6ugr2D
4ueYC5vDxN4Ha85RNKgRHj2Hy8hyWwptbjZ4zoKB9rn7gH7elVUQOVC8T67rXi0J
n2t5HhOFSu7gC46Sbp8jAE4+GbiLMoLrVMt01IVD4vyQ9277Vf3PTF3+JkJxZNKl
Phk0pTLlqxuoUUBavp0Z1CVZCYSbtd/VhX7sC435dfskUu13Hw7seotzH+Rx9gCM
kmBgwwApx+sp+3HzP+VS7dBgYoyQ6GT9T9H/9p03sADmstBwCrb1Y8Qdrq9lFTsB
zdB37OoXp7xgRCkCMPuZuZ3XPDylrl9VO5lkBeUXXxRzojlX9LeqjwWAUokJPU3+
DnpDbJ2a1N5FXcGYgAM5cl8p7qF1aRzkw19b2uqQUR6pwZ/+D0ufeAW9IknEzMrX
hns5nOIr1+HNyxn2t75kXLfISTujmVPVVNzdUM/PK3LcItrotw12dUjz6NbuY5Pv
y/OC8o6ZSQcgolCfyxAKxf5UD7VDiyXNB+P40YAMiMqUZTAEmHyJN7wIHNLj48Sx
Vkgm7Sr9gQe6a39dYiOUrLWQZfD/GhlaVFf5ok0ylLuo4rBF9YX1oy6jLJern8jy
k2KB87pAJhWebS6KLPKaSiQVEHop/1PyQ2pT7y0OGVQuIyBWwNxisJ/ekGYvYwrF
b8pZDDNKdD8Rny1yQ810ry/XffyL9E/gAElWX2aLmYrOd6WEn5mtJXtuB/oAIEPm
9naiPZJA5tZE1xG1Sy1kVJQPH3rethbaCQ8byav6gxSG0GDhLOMtX2sm4AF+0Lj+
a6BO+AoklPkwIuLEWQX4Go/w6fqVNhcZzBoW5fO0voWZHi6PMV1EKB58u8QFN3Bo
of4EK6/9VvDunQIs78ab9Oau+015p+mOv7E0Ou3Lekn4HftJLTLHuJVJdN7h3/gz
8H/vC4um+0ss6y0GM1ZBVxNcdDYm9v+ZiguNU2la6z95SuNxYM9z3RSgQ7SIQ5Kl
15hCthMh3nMbNvA3qpaKQvgweGioBrF/bu3I4wIFRoCxkg8774F3Ux0PnO9L93cD
30zJQzR9T5jRHi40fuozpoLJHmNsVhdGUHn+J9BYvJCrY4vTZO3oiDY6n6lSf6Qr
dravSMSTnov7H3U9FzBqyRM3pAwToU9f+9cQxEfrQTrAqcwhFo1MzBBqxptPswUC
L8wR2Z+wsejEuWXPxyhA7AK0GaRsuBabiZ3f7NPXlTDvngab17MJsG07IWQMcQhR
icOflXy32gDmsgQ/W7d3YXYeqloFcAvqlBHk1UJ0naT7Vvsi7alHMRKgQVfIiyzB
cTP7WRONUM3aq+HeXM0xA4WXnOQ5ZTLOCiimlk4bfi2HhYsLoVJdgyVDcOgZpXlS
MnFXSDWmDF7Is/2eg+3joJitDoBEhPPCrt8OvDzR9LV0g4cC1hrvajtHT9CPgn6a
g4PgipEXXvVpVzU/BEWXzb1Ozi75lnQnQgii8q8C5ZnEMcCe8ZzRQcuKviGpRern
AkA+Q5OiXFE5To1ARYamET7QksiKkZ2xTbkGTCXqNZKu9e08/MZnqpmum1YY8wt2
8o/74mbuSXjL4AS2k6u/K3vWZiWpl4Stm483bVwjwG0gknnkWNCWqyotONh80NBi
HNncAcaT0O/96DxI9EAogiI8VxwEfDtQXPUKzngRnf1fKEuC2iVwlX4qlopWHwLJ
r3PI13cD42ZRV8DYFKPhVCngKN6bWU97kz9s2jmyzV9w59LnIjHqvmKY2+T2usMq
RADUTj0tTBJjeBtg96ostMp7qWdnTMQOCHn6DxxzMFaHlpeBiynYfFF7gXiC/u8B
d70EAAXy/QCxKgsByCI+p7lBEtAQ8rMgOU86uW2SWe9zTjvNh7gnB5XZQ7s5FiT0
WMK364PIHuotK+Z5BxDFjbJATARpFhpnH5o/Koj4lT9JU0fV50fgpVdbUaF0sR7p
+IfBHpWcYgH/jqfyEdMWCrBHk50QOZcStSQqkFAABQ/c8hI0+2uPQQrVesK7tqQB
Ucf0RPcl897YmEFMv4KPGQKYfHQip8AOcB2sOGBzP32n6H9TvxGW/yYwouV2oHqc
046uWJSthggiHLy5YezYK7EsU4+4wFdhffNWT990yY2zoeuFqRpDDRXIozvfW5SY
0HC8rNf42Xe/Qj4kKbv0tu/9VPXrjoVgZ/LzjmbKwgEVIO4uOzuvMeQy6b9+mwLG
B8i2aASNrpLn8jKl3eMbhavZ5+A01uuWO8KJLprzSOvEsbR9EP85PLWg5RDwkYwP
tsDl6DF3jB4DfaVCXVVBfNYwd9SZUvN5r0MV7nAunNEMcS8QiK0G2c6nT6Px9LgD
eAZbdSLbQAdqN0G+MHDyc05Sh+FGxmWzrANGlprpVAXdGepz5VtjYKbY4foTlYjs
DFVXnWe4/SwdPxOuzlKLi9DEx5gmFdIJ2vufZT2h306XGyJMlUsq2yF7xMUO4Wy2
HNKeouTJxdr41Y/N8ylyBN8PkQOSYExgW9q0ONhwUGJLU93dpsz7jZgRlVSKxVQJ
tU4RIzIU0u6DFo9HC5YHhUIlQQWhPVbBrTSA4K653ylglXX1I0T4cWlKKX5cBWNQ
yjb2DjY5od2q1CldIsfMMI8w9BHsV7nYgkIklvPtMI6qIAKdUL9PxQz6v1lFPGG8
BGkt9GY8oJNMxE6/HmfLHQsBUWRDo5dCwACQP58n97tzvG7e+/EAlXwChNZYgVME
Yyn16VzgMHKCewqUBP3cvuzN266gdz84foL0C2B12Gh/oewK5v/m9NbMRKxXM6aK
QQbTkJ5SLxQcepBsV2NmDY4OcEMSsqZx9WGqQTyA+/hIHmZ6koiUBSV01OFi8d1R
n/SAuLa17cMcVSU4Jp/dpvJInKS4hkG79zx7m1HDrK/qlLAEIWyHGyOFoc2VBsaW
4wceJh1IbQkhmUqCjYNsM1Um7oMIv+IvbEuQsQVsMNdMgAAifZGrC9H/nUe5BCu0
OyfmV+rz7E9tOmJxl8Z+zGCF8GNzqes7Ojd51jozRyeK4ifIS3oR/oF0pVe04DGb
69glq+FVlVhbf064Xdx6v67aSlrpYqnPmdwMeS1UYfUMOWzBkfYm4UZ0IzUiGSdx
gJTr16UMn+nSbsDLA5Z0/02ITrr3JhfJfGd3U1RqyHqNh5E/Rx933Xi36UYYw96a
5uAcY8nL4OkxheXnoUBTIaizsqmt6Iq4jhRVugt/DOohwdwXGIQ8/iIeYJMluHpu
/Bk6o9bfcE2NasNpMhKGKS7k95UyTnVgQCasfU7vwN5xVAaRiAwCLiUebZj3Npvt
h+h957LcZ7YWGweSbSG0iWy7Xj8TD6jzd+CV3fqiw/FKoKbZ6evWzhLM98R50cVc
KpAnrF/q3KzqpdHAs+nAl+ok3zdG2Ea6DaPFnyhazRwpLOWBqciug9VukNYLoUll
6AP0mcQZ4cpSWvCq3j9sf0zU4ZsSDdyvC9DCh6pp+MO+da+snIKQv1bO9z2S9pW1
zMGdd1brVDnM3MTeiLt7cWmEAKUxk1i8zv901EUS7S+BvuoFNQxyaO2zyGHutjao
Z6c+4AOmDlajqMJDr0EFuxu7XVMCuy6oGI0QZRqBpiZ2iP/UCH5NXjTothRheaGf
c6Pcoderz0bb3RB6CwBL2CCTbZlftk768ZcgV/4cfOfR+5SwPT1BtKl2AG0LbfIw
Nen+4wRydNQ9xvlYxBwSqY/nXUoTyiJXY+tXSESAUPFJoZNDdtC1q9YkyuwZNRwf
w9QlGAq4WR0ZoDcLBLrw6jje3UJZ9OGyZzpWYN6BRfY1R/CyXWbu8UGpoOR4cdSD
xoZHVnSG1CIRyYI4/gDVg9HHvipoK+QtudqRqI1QDQIqmufjUkk6UvYOsYEX8bSG
AcILMmNhS1szsUi3xl20wooqVhuxauN1KP9ZKxH3kqdNlWYDNwF+ObMA1dHLsmGx
EoC0b7/z6FrOdu/zXMeEWbZVJRyZPd3e3kxiqVzVI7Hv6OQ9IXU3uzFTM9ojx02d
RXLZZ53qW6NzjmxlsUB9rs5pNnHhEg8MzdC3NiFHvKI/3LDXVQCuJeEqOm5S/wV2
vW5/zz3soEBET6qgM7391gxJuynotJxltz/QkglrDjwpYnnuSw/l92I9RYl9UJSl
NbWFgvnpFHyws+u/B1HCuPfTC8CQ899M6XTGuvGccCw7pshivSv8V049WBgD2s3f
f7Re/kszbBZtOs/EKmzPZsr97G9mrCoakEUWvUgQLbcuylctU6iGps113HqqKW0Y
kMHuK3/NVsvxqSQDjnKVsdmbbWMYCaQcUtVU9AKRiffVbbS41n3WQCZmh2mBpN2d
xlc2kdKenow42AgkMF1CSJwgId4jMFy5F2xBkbfy/in/NW0Pwqh15ctY/bUH0CWM
DWNgljpYZJd+CCvy6xUK/GZKYFh2BSF53fClyE87kB0mxSG6ypFwn1+kq85stw+L
KMpz6lupyKGaVttkeq1ZuC/SWYRGPRjifSOW4MeGCuZpxG5fOpKdfKiKsNQxDcbo
NADo4L596lBXiqL3z+rmiI0ohEJv2KSnMV14t8a24S6+QjuboO5QvG+h/qrV221Z
v5pcmwdMVEReDYCu74rnpo+uCeKwq228yMkKpSTcPWfS1Urx/oLat+zGpL5rrfTp
7DEISohUXwBFw5YIwjhyllVI9KXzdgeI5zx1CovM6RBDi8NRnKuM/80sPwVKrs+a
g3F0/E6EkCRhYhQLJQl1zsXv9T6V4I2Fexv8DI14G8VJDSU/ZKPGOcwYK38QHLkX
WI1F6amt3lFJxOKoZsq2CSwCwIf7IRHJc/UlagskMBH7ciP70IGUT8edGhFSbVWA
RhKJSa6EfiuAz7RoKt0teMKkH0xD9yAHRqOAe7KjQ/Vt7DUYNDQQoULkWT+ixpNd
icP8zY5I4sB4+3Of0U6s8p60zsYB1VSis+0MT/az2cQjvfI8P6iXcVCutqKWo7La
82ppBb14ONaiHzRqCqc6SXjKr6XA2bGfIduChudzA9cH2eAN3nO+0RBkYOyMwDzZ
+3JkKSGAyCUn8wCI23DBj9AK91kNzHYxVacDKEmuCUzoSHe513rSY0EIiOix8bqu
sTxxwHe7dw2dpbS2SXf28Q99/5lX/UUKBMB/8+MpDHWiLtxKU1axrTB6+Iv309qX
eQDh7ruWN5du7DhJMtXwCXCh/DJ6TqT6pqNB5rVN+xGQxXDV8M7MuYaZZuC+RjBS
QDMvWWyExFVWgkPgufWvJv0lrbbEUU9ejFZsq7JTjCjiB08POAiHY5Ryt6k/0NnI
JdGzYQBuI5wDQU2vD3oGbQuhzow6mWJ2nG/GEjCD2X/B0ff2OvhM62M4m2TcKEQ7
oZAcPujaHcVcdExGIYaNMUu/vHSljGh0aFGTh8uQNtxkKZ+KG3XwnJ2LnpfkpYCV
Mox06O+2noOsq/TsWFgXZDI5niJ+332CdmkVDD9Ah2ulGXGI1rL3zKL5LVgmwfin
lA/a2OT12xmDLaXo4M6Go4Kc+zknbS+3btDnGx7kaboKW/aXF2EPYJSNwcfib1dV
1ZkW/Vc8fmz5f43srIXH5G+5UaMD45Txz+Spl9YuSBdvVdH6d1zDFFHCif1v0fVS
/NEEDQWUVAdZFefCyavnUlk23yqN2277kvWrJZH1+Ea/eFleOKX6PlbUxFbWiGOA
/C1yIWCoJZsaENsab7fsRCNCltmK0QnuCoJo3qOot2I7SE3qIIuwpUhHyu/24ZBj
Nkpe/O6CbYxPxYnTYeWuvnZthzGs6tud+C6n3opTORBC4yxKrdHLy5INv8TCyjh7
UQCnbV3XXi/YYzJt+IV5OqO/EBBTKndBUV17eANKUpsJBcyiA8nrc2xFUeRnjgG+
HId8QsDPSv/MSAG+t+QRsqqIE1117TMaA1Wb6UpJxsMuz9OQuBSmqU2Qkg7MuUo5
wxdTTpX3yjE5LNATQV4SAI5rSTq8zQd/U4rIymmEOytJ5tbge3KfbKx44S2qJ2WO
APlhNkCR0vUuwBxVS+YcNJOBtfIkEErnbPnlvdGsadnTApWePAbGqp0NGmhkWMtI
hivWYsXqaWDT34Wh3fOUQ7uFWErXYVbGRX1/VGasn4fNiVIxQEetSRtMB6CqrYLc
0qska71qJJwOdMKOsrJlianxz1211T3oKBtNpUosL63C2gxsWvX8BSdjbvwwGkk6
GIM0R7NECTQGuJElhDSTyAzaHoRHtv1nTo16Dselrhp/T2QhRpAzf6jsN6XIWQVH
cvoidXiMBk+QSsrBIAIl22J3l5CJmQeIcbpXgUKyhP9z3NKQsF7uimrmJ0A8J0xF
b214DYXm53dcxSqgWF6ApLtRuEyj7Tu+Qrr7z4du1qL6HVtveouHdt7s3Bqf+xg4
u960gO/boA3CkU/N28KA4yeU6m8FERBHBtiO+CJ5Q/T8Qm+tMVNee1Hz5dCwZIXQ
lmuivevQgtfnSV58DjkmYuVRZ5pe6NJWKr1J/eVKGAl9zFEHv9K9J14L9cTnoru6
pKZI0iPvoAThfsYb8avWzH4CMeUW6Ofud+gK/q6ZF7RVMl3GU5tv1sPVerpDdIVE
oKWY9pvhUMWyGeiX7wOwzZGtzKCip3Zzonv15NUONUxzK+ar8o+wVzyQl2SHVtIA
zMXfmaQ6cwQ4hKHUCcXlC2b25FjJ9NUwlaA+0bVSfD00xECe1gVvYt1T012H6jBb
vSddzwrxc37Nzj8y+hL3ad5td2sxqYgGF68EgT957BnfzATSQ1uoPOl10LUo+VKP
jNhuq/7i+7HAKP6Tsaf0KvUrUAnec++F+tqBdjqveJV6DTLR7aqfDgfi1ubTU/5g
imgEM7MUR5zVf8O41PCBeinuqj/zErjl4SwaxuKRCNQDRKQL4Yw+m//UxUUlEE62
B4W1/appgbOz36/BIFOr//8TG6Nu/176PnQeOq4k+XR6lDgKAouNoHxcGLiuodrK
3NnxrR9YL7JJFAq+xgPd4m0GnMVn58o5vmbgZ9mIa/eFIaV9Dz+DMQMzq4pt8KOa
Rxq7UFRMbZFAllnYDfwSNjsLqA1mzrjepdafnizobVXZr688RiMa65cZuTHImSUC
f1EwPn+ljF/XskYE2IcBRG7MElANO4X3lTIODZTTxRfdexY+iiyNgw6eFDvL+tQU
kPFuJwh1xwZZO8JVmi7JYNInOLKQuNOElOOotS1QWrwPNf7NKqW4fLYMyIElnpNA
q3pCyApluodt9Yhmyyb7VmPWenQ82Pg/+rXhENle2A0t4ZNip/UdUqIeA+pcOB+V
HRYGZgICbOHJPQK/vvwZtHPBDvnsw1uYdQDX1k6bUPta5h4R6HnPgdv9ByB4OF/8
AqqYBJsZ5VJgK0LMfrFbz0i0t8TTLWJ8MsgABxwmOtZ/Dyo4FDCqXt3QU8yVP/fh
EthJYbcDMxpQWV/pix6FwFIEooIhQ5/vE4ZZXsV+rXYYUuBO1ESN7TRi/e3C1nrZ
CugNm6mo6PJPkmatLv7TvzXQvStl+322TCxEL5kNRSuDFuEY02ysD2iTvvHFdVzh
bPz3zMPwAkl+RSFD0xgwBDZNdIkRU78BrEk9WtSacIGWmMm1aqyr8KNDkI7XSQOr
6tvfnPjPcUJzcdwO5Cta+LDVzaZmIP2X5r1ODcnUiHCc8eIC3iZ7uGCCFFPthhxl
Dq7N1hIj3gLX/Mva5v1WGDpvGKiQLFn/2/YHdeUYCmn8jnlCwjohhmm67EAFxzO4
TJSqQRZjZb2mrdH81g6UuBAYWO3vttOeiHL6K1i7dcvdfj/LnhgiH8j+0IL2UexA
BIUG9LInphhX4UJX2I40TteZhyxoFmJljN1rV/8bbwFJEab2xyXiateHtqEoiPbO
mNo2SKhcYKNsMv4dgujj5aA0PrdW0XXKG8tN+56HKC1dJqzpWlPGyUhgZulgt2Rk
Wknugn+OhTjuaqEv7DXngiNAPTp9BQ65vcMKX1LL6MO3pvUL0LC3VPKu4tWqm0t+
+xGE5Xo9mYq4VlKxfmg+R+f3kfmgK7D78stijtQ6U37WYGKQOiqY52QoJpQftw/Z
WW9D6JYrIRmh6TNT8szCRsBgGbT6gdg60voPlg0JGs72Z548zcUxTckwuHQYuTW4
/65EJCTtbEhEG2A/xxWbEWZ2ioYjHWcuZpFqaoxBoluBSRu1CzHgNkfH+2CjTZFQ
gogUztBqhzmb071SLFvgxVKSmivD495uMAMGrsNkz8Jq10zxwK4Wi+OUshOBVYCv
eMffVvNmc5EdNjcTkQAY3HHMxPUwXy5P3mQTJJ3xhKIOAwnu0N2M481Rz3HDVGJC
1eVjX8svUbthkELRcwsPuMnNSh7Dg4otRp/lUz/l3EQX4Tw3o8wqlr+5TZT5xsIA
cH/TFy7mxKntjrqN/lXXCD74GPSvunZZvhM9Kk4bCzgjB0lHRh3VuTp8713fgto7
BcwJ/TAFYnx7nwjXdaNYJtyJm0CsW/3m4eclfv70iULwtjbOQJglRH6+QMN/ZZS7
D/DSed+mwEtt+mzGVnWF5ax3DqysImumcHn+V64oPc1Jl1az8t/i0HJos4iKZhtJ
UCcAAk9oZMYxe71s9lYE3aELfosxav2Cgkewqscu3v4pPvgjGZS9se9FDJUSLA/d
HUtQI68zGKxlxcSZP+6yhL00qZMH+wbsP0DiffO95XdvFsPoFZDZHvBy7EAJOpeU
WLyghmZYbmKbLb5qrv9g7YmCiYvgPANzeTGStMKOGG2QJHQ7MHZP5njPhiPEk39K
B8cIqv3h/iZGIwIsiboNUqyiCk9dOKMZEQzw7KUKDd/QnDOXyT3NHyLiNlpOtfvQ
xEP81VCT2pAD+lutUCaNOza9QAtcY1YkCsLIPCGJDjewx+0eDsRpc9XWTVqFLQiS
EK3OtjZqSltnes2NAVAkRvWpIrj1LVY0tseFFFzd5t9XwCz4QJ8v4EF1nYFOjkej
82QfBT9KuKQOyIdHar++WKD4lYS2bWZ8KNlbxhaeJg2WlN8tdAui7fS7nrFcGAag
57pcf7ixjISACbQDKf+vjwoIjYGhgHDhWN5hlDOWgMId17uXmHXgXF3qKl67nSCq
Y+48b4cLG7DTZDZFlNcmRjtwt10fPQYkZgfifLOG17osbRLdyiwnLapt5Hd0MjK7
TlgYR0BuoICgwlQUup63biy2b1oV3Rc6dX2AzBakqrg9ryNKqHco03YsseByh6J6
rc+yhz4jSVw8mk4Ab6ve690DJk7zVVAXu3yULVJywy7+xfiVxUtljp2PTCIwlRUP
irvI8mnFPmc4maoIhBFnSNUuiGC+HHa8v/Pw+9u9Q6QJyA7FwEbCuc96f2KgGyRd
vSLEllKxK3puP2cp2bWNdALqHv6DiJpP50alAsrLIOZkm6E4FnX/sgkUBjkO7hzK
ksjj/gzz+nu9K/aoA8BHlNwjSnce3KfNJ2cUwpHYCefAjsytcZo+eoCyDXKjBJRU
aD3NMth6eAhahThNwjqNB4zT6SvYAfVR+FwrwUZ6jQ4MSuNmdLzno0QyGwPfuX+0
a44bQq94P6JNxBIx7+kYudlLxtFLlDS2K/zy8Gp8FniynZyHfkLFUoq7rpfLu/mP
rBsqjuSB++bdDVfrf+yLDgY/mxSWdK8F8R8TmhCgi1hdtJX/W3gIecHM80Tv+MZ7
b6dx+zKrjVCSMm9jFVTT6FBM+8FDpcyTKwbUUOIS8VLCCqXmwrGiJsi4oRmb/16M
jbvzEyRzukhyw2taGjTwyR8va1IJEs7fTqGRCC58XH0M7dlYYPxAVLBL4yK9jpxg
yqtwiJlCf5UNibKn2zOMZ0kRKE0TCSc/0O1mwZQa1rGwB1VgrOblAOAaQletG2Z4
8/ZRWMeXYt88WqUO33Uj653JjN69xjt7d21rctYxvYycmqnL2QJWwgjtpAiIQiDQ
5KrK/szbyHy+XseBjgrdFAdVnFU1WFzes4Y71DVdBPbK6RQ3eH/6bpKiuh+OI/Pd
Nn8W7nAn7AzOZzg/ze4EGhZb8Or2IpJL/J10clAfUIg/EJlsLeC7jD9CWmTXMN+v
F6Th7iosPxDWMCO2DGo15+dED2PasAQ+N5jyApbMXWNxxPODdlBvDHI+Yd2ubAJA
b3/F9Qw49q9xRjnplmxt01jVJv1icAB2WBVQ3DG7Q3KsRuy5TXaoy+8dUZtLz1Wr
c735OgZhF/CGuYDhKBY/dasNqdSlpwa2qTI6+Plm7yL1gwuL9EGzZi+z9Yp+v/e9
4VQVXduRYqUw+SXEh5FA/SXDFwFWYNlrUnZML9yFCXaldIOrIsMAxPULTP0f/uYg
AB2uBw0Cgb+pX0Y12Z4yQol9spt7xyJvDS1miOc3hjunvKE/dg+tv8NQrPU/Btrw
wrsDzVO8MD2zsoGOLW8OXuOS/7hk/YlUv2VmwCQTzIOWZsrsJJuZYwsnrrcG/0jI
DU7ZmZFKHIxpNFFz7+zqI5YcHo3pzuvrp657FvfFi5mSpjA5pcRH2knGjGBJPyZb
j6L5QzmVrwnn6uLJqQRbjrppueUWCJ44vQAVpCNsR5j/bFWAK209kc+/3o1R135K
uo83bzt9DEp19H3CMuuVSFE6K+F135DjtSK5AmZ8gCW/wZ/bjjah/5qiwZiGluk9
Vc7xhzs/tOyi47db5n6wRr/pSlvK8EYOZW8hCRehtTN5zNcszmh5t1iMzYGV91Af
2WI81iJeOpfqZYY2i4jqe0nmj5z0Lt0KQ+UHThfzHsm3xzNHGwQhJiGETpMPfwVE
JnAMUY8CYvFNMud1JWOoIYLC5j7WByhgkZZI7/h8G/noiefa4v0mCnIvYNhRAqD2
nKMR3R5O0eGtzjBQaJ2brQ3C4LekRtHtTNzH6RAyQfIoulikb19rnJX0vbJMbqYv
FvHO50LPp+yRNVqMMIiM+tOqyTAKg0K7EowGN9NApTBv5ZbAKfxohAQYzSGNcquV
sdXasD04OHOBaokTPW6yt6yb4XGL4xy3XH5N/VI9lOt57977GnEKmzfKmVy5v7Vs
/tHHOE1kVTZfVl4D43QX3MixMRjsiC6FU4GM/Nc8al7m68fbE55pXaT4+kdsqUyB
jpvNWlbISN0aoEK4uZ5nt5Fyyo6rks5QP5uVBjm+KqttzSy/RhE2GBdsbh5HnWGw
o4Hw1I1e4N2Yt3Uq9P5hLrU5Zw7z5nkA/YeUm4Q0yRvrTtPBduzZKUKJb6Xb7Wex
lV0+v3ebAyJcvyrCtrI3bP2B/97hVGuERhe0uJfZ79I2l7g3GhSFstTtHVEZMt3Q
uqm4WzT1pj+xbkVjhMVnEixKjU/Wjj5kG14TnlVtCObgugRkLbf6P1fzMeVlXMpn
11jFgm5TJAMN/7MjpAGa2Aywcw5qY2f0zcjm3aZ7rEHFLJI4XpXC3fb/7TJsVGDi
Ii5KOPi27Vfy9alzU08J9RGD3o/Zr3CkGXsa+fXht3ej6w0UQeXuy+zS97klUtMA
nHWRodpYzbQIQ9LocCQpsSZ1E0t1q4Zg9bZG+nzLNORNS3T0tkrFU14p5TqO1oJR
ni/mDJTDYBDxOm5i2LKwFResSikTwXXdcpiHkFxSxmtxm9zoP8MvZIUR1JJb3Zui
CoiF/V9HqE58rgoFCeM0Z0slF+RxnhVl//H8s8UUurxVpYajVVqgasEQwZx7GRay
ipk91mh6Xij1X7MxEFLLXMVf2JWq+EwTeTy8pH2LxtwTr7QfpH+1ridA7Aey81PS
CwUuojl0xok8rSy1kX+C841H/53Y9lOyTAvklISlfEgWJAOFzgkuXurjf+Nurme/
CVWtXvtD39dLHIYdqy6txqTujCOHRrHrK/mlIOymM84Nr/1aUJv1pP40N44Lc1gW
WrURRFH/js0OjeaQiVIPh3+Je9bcZHuWDBgYZPp/SSdN3zhgOHF8lPlqCs8gAy2m
tQMjNOyuzF7Z0uxtbP43rMo23ryiJderool5DBG+R1LIk9nV+A47YuMTCgQqzW5w
jLt8+R9maNKkwGO/ZQ6ESbdnbqmIU68s0/isrkQoutJUfpMUVn8gRAUliB3chn2o
X1usUQ+Uu0ofWSX3gzB6WKWzIUDtzNcay24ccyVXqR7hOnbM/L61O18rBlHm4jsF
t1gNk/cg+sCLAiLywDjdSwWpkeL84qBh7z+7BR7R/LzfM1ff7OmXwttN03BrYD0r
bJucjbeykUivvacWhVAz6Z54BjpAk2lnxniDpQh+XLMriNaw1i9V8aPdw+7WmvI3
5s4B0yjgdbti22gTXU4H9FxROFxjNg/piCO+CN9NU1OPqGGQkstiefFXrYcfqjPl
DpEsxh2BwXUzD6FPEJRXDEwD/ALuSL2JsHuOZe0SUTdjZ4fWs5iR4sZtwS013dpx
hA6hFdnOfh6ukui1ae3omsglWlISFEUf7zrqCjqerR2z5ZbOqU0gGxmGMr+piSSv
IBSOV/bmCfk2cnt0aKXb4FGaqbdz/HOaZ+IxssL0W0FIbBwEUrfwGAs531gzxXv0
ol+yX0gSCC0R00Z3kah3jdgUepgLglWdydCJF0eV1DGOrXtDVKwcVUR89Mf/VBfo
6FB5KpBoL9ItCQYyhWWWG4pIy5jYo3dYtLNT+qJ0pmBo+sE0XH/S7dA8YtpUrf9G
2VBqBBO/GQjCbv4WMrJlNXRUy5BTX0R28vIw2bz47kakgYdOOGUKLcYAtiwuLDp0
b4So7/XLbgOD0r7GrxY3OgQdUpyyM4l4g5TyQrCMXl6X+pakdn7JmEyuVoWG1n/4
NFQYC4r8dZOvoF6aENaIUFIzqf+lgV74Q5425M0+5Zb9iXHkDYT7U8BHMnWSM3Rd
Rz4tt5MpbQJhdv5241zv2wI0v/MH4XFLdnTCv6EmKPDXikq26o44KvlhYer3rhV+
W2W7ne05qtq1uXHQkhrEBDK5nBjCCqvdxlMCi5uW6MM2GGRncLb8cpjpWoPOaqL/
Calr7H4GRIChjtyiiJjgQPaSiIkNaAHI7S8VA1EacwiHQN1i35tKaOXCUrRudCYw
cQR8CbBMvqjpmLmlw4QOO1G9NY+2IdOMQtIXfSVoYHlFpUK6QNNJgN+bQyhKajOG
MSOzd8OSQ17RUUdkB8nsDw59qVbdMPXQ2FngXfUzJO2i0Wlvb4/u3uR/FYKdxyQ1
9rusDAYiUEk0gCtsjsBvEPPI8bHYMDpGAAmcr+/w4qKPVWXhJmLC2waxFb0VfLZk
tJvfXRtv6uqJS3waJQglpEa9PshktFDHmyqBDTGu4UBBv5WkES4egX7VjPdZSPG4
8cEOUVgTCLeexBuN1nIqJud83ze6K8zHVNb+N/f+LSdL/iJ1m1He+9xhr31csUVh
ONijTCmKGIYrTUcDeWt5gnEJVF05iYLGW4ZFuuTjRPD3syRHgO71JnuRSlu3m0R4
PBO52dut4XImuybnjKZqjF4fkH0n6prERzjV+gBWAPOI2MBuItQ1GEoCdNGtfBpG
BUDf+w12RF9/tIfBUIieqaH2KaZAMVtSdmR+GUWPcWFJ/awXpx6gdpGE4W0T7rhN
2XCs6U2dOaw7Mn7S3WbIaXUxusuubVC4DSXRZTl6xExOq5Myb/STCBZabPlA+fAK
H8rJC+aWluyrrfPvk7+O+JBlIrTFtbbPJRUugiQ53TMrG6LLGe4qWuwYqFBx0yxp
B9IUytgoupWb+lut5EQVXW0whIU6O7I/79NJRpsxooSiol/SApP3085lnwfoPLG8
u/snhtIGPi5j0rCfo/5mSfU3wGyI6o2ztDSkp6jqiK1N6jiq7hHdaQO415tpOCPb
1Ni5fh0tblaOJMUq3djOMd/A6TThPccDDcdOQI4i7GsM0m5dFWAx/Q4rOjji09kf
wLv7KJRDZYc6gloM/nibBLKa5xaoAqQE1iKzdgcTm/425ZqLDW52SwHW7mkjOGtK
cj/fUAJ1DrV8zY7jr+sdrdGGeXxD9XukRJD7hBneuuisiovyDG0hb6r/ccSpcz3y
P0WoCoi+NSRuwiSkZaeoGxjEkrSfLrlO7svlIXNbo81RmCrAg5sNkSvjkLePUb25
TbkPzyzKTM3N2u6+j/l3zwRltPjNN4MSMfBYqOWB9HdjzrbqqjV8CeVXJ/MH/WMU
9ae1VNVviiqi9VbYpHatA4cjR0DsjKPNdKseg2LqkmNv3dMAamxFZYTL65OMIoL3
pbPXKFYzfFmjzmuL0w/cWpBh+i1tgqw6rISyuMbxLwaC2bBPjVsMNIWXU3lNR8AC
ohZJudBoMEqMcz+qNh/n7dZtLFP9w3GiBparr/A6l13P+9toN7K6oMg9/YTVfhH/
Wcvukb+udMOMKVXeDyjDjdlJZVvyB3zB8BjsepSjLo/TQjkPy6RsvohHATiz31Pt
K8/de1VfCDXNOMg0OAaD6zLUTVIZ/S8hTpJhK8rNs/wZMv0BijkLglIa/JXe5Q7J
DqqwSb0ExztR9KlvRpk35I7PuEB1iidKuKkjrrD9v7v7ceQoHN1ZbOwgq+CC9Bjv
J10w+nsVWAb56DEbvYKXJIToSSJ+oKZ64gG0jqVWGBz1txXEw9MxZ0bKUa8JJ07V
6RrRbcvOFT0yKc83ALlLplQsWK3a/CK0P8bRBloj1Yhm2nyzshaQJBJSaa7a1mGf
wf4W1PwGhsZtkU8sOzluJ2v5yFROuOLBupQ5vii2VId1mIWE89CrdOvs3kUQ3csJ
J84GzetihDuQOAGyW006s+OdtDhdxj1KjCI8wPVeYSze85Cbatdsw42/Q+uEoltU
nZVzH0kqFRoqR1mnkQNA7imYDxpiSRhhmdpToeNLVPsPlBgR7UdMpZsLnHHGh09s
C08xlojUsn/91Gs+9TfH5BOjVKCVOyljsA000kwIf0Ouplqp2Fiy66+ZXBmYztNo
QyMDR+uu7zTfWKGxd7stmkWTAFZYQHPDhkfVkyug5kFuVAd5FQZeTk+dA4lKA9q8
cBq7FWfaewTUTXuX1H+FkDw5dOoBdauIlvgtn4y6YzNnNpBdECuoImgLLGhFVO05
4HYMj20XI8D2qqB5y5EgHhPB5W9MHr7swlmDzmtRNwUcTnv/OY7Y0RFBmNcZXzkF
G1T6RA2CAOmcPceg665zA15A20TJoRKJGkxrVCKCIAi6PQO7ZSpTUElM8pB/kp/F
Fd5TMj1OEvfTWtq8J4QxUrqPaPlroG68tkqji/mSH56TAyduTYLXQbbLzbpOJonL
MTDg88XUiDTBHB5v51nR2o5xh0YKUJkFbZhfbLtjK9d3GQId7pias0ADwuWyB/hQ
MEZzhyVt6t/aUY0vXn16gAMLwpTsY1PhK54LC86IPRDTFlgtEEqjdBu8uUeyOPkX
WJ3xA4JpvXQ4PBaAOF6GzdGCuEhc3ArykPy+ryOsgE/dtfN4ll8uul9l1SjeX/oq
QLsmIuUqyFZGyF/iBPL8Qvr6pdmQGctWnbMhuji/pT6upnVdOg8NVQHVaY3LvWV5
rTyiDRr4XKr7tQm5DYuGqW4iW49yCjIRQ5CNVoxmosd0kvF8CfUSmiGN0F9p7q3e
TUTPiKXLiKFfBKd7lhNIqr/vZKleRVBRddFniJauNeTzjiDjiIPih7pWerHvXDzh
ae3lhju0yHWuYie6UzAM0s+tWWiNHayGgNlzQXnoLAedE/USBNwJpjG1b3thjbYE
UFQp1p3jw5hTjGIS+w79Id1YahCkEjiTWDuufOq23uQdBdAYZuMYq2D2aJDSiBK7
08qu87U6KJj4ywp73RhUbBmq/cz2N+08newx1d1rRL0P//Jckro2Q2SBi31uzFkd
fQ1RfumU06zSr2Nygx8ntu+ysvWHU+YfNDUvNls8HwHgtJK1RfTfnhHN4/wscwik
ssECtvCkKbB+Fy36nBbONA2OA0JQRKyYON4PNb5x3GllJ964tQ4epJwnVYW39ZtU
b4CKFFiKtKJMGneV23MwPm4cmE1oIb3VJ4Zf/etecafxt3GY3DEv1XlGTOCzgUZC
lDY1PYm0DvJ+waVkiv+NCyT7LoahymX16nrs9JXNFFlcc+uy2fPvq91AQdjV4sfp
1h6HoxpK73cuNNSWrzTx/WBmaPkinUITox3THkn+t/VkykX2BzdoBpW1PYDtbF4k
Ou3sr9BqtakEh4A7QBQ//eDYXmVfjMrke+W2B4e+6DXcWVauem9fgU8t4Vo4d1MJ
HgCOnPKkovwhL8uKET0fpH4y4Se657R1oPYWl6fcbGDmKFNhFrWV8YueDPk7sOZK
dPpnu5IpvXIQpeHdmT3mvNMGJ0TwB4GX2tjTWTeJBJOz982JKcx690iJ037uN4u5
2v6Nz4KAFoYhhGfmwlIpy5gcticu3re9E8zSSTCzFj3GaxDCEqQnHTqJHrLhhb/C
e7NbGdj7EnfY3VStVEM06srIYQXSOUhd1DU1mZUfwXDH0wCcdmyJ1lnjBqypDPlL
3yZaCaISALRPm+m9xQh8tBjd6hqAQGZsVjulWzz6+f4GlnQWlINZLjDW/lRwIERz
RZDcRfLeRRqU4uC/LVyQu4Mz/7eJgDnAoOVSTkHqXtxEi+5I359la4aUf06vxmJB
s1dZCsqtH8PZ/ZM/x9smNcMXXynI2mbElcOjHIVnTMcuOLlmIA/65YXlHtCpxRgH
gyzc2iRYUz+MnvWZgMqW79d8cF5VKuddA4lKQmNbnb/yqtuuswCjNfPah0zHwtLH
HEcLK0WgtteaZyN34AaQ7ixHY0ICDWHwmnGKfPV5nfbSMREffcAkOxJDhkaAU3uh
sSkCZRiQF7CubhvpyMMZaI3n7MlpNwRJGsHctEjmBJ9iIWr9GVYFKsmC1OFY1q13
EdNgjjLGicUNp3sd3/cpHPukcu5xZzJpLqw0dVdBAKybMsllUmRQhg0FiP949COY
Gm5zKif/85vHOJrxWqCb9jo74PhWQSyI9zQBN+BCfZ9tnedPFu157HO9Xr1dyDA1
/OvMTpTUMf+9Y5GXJMlMTT0SJyxuf9o70/EmyTuzOBHD8T1y3LfXhWS/C0Y2kzAN
YCgkAh0vYRX2QZP2BDGx6YIL08NK5t1H+ZD4HS7m/MW71XhMpmU6EmtIuJY8cuzF
luR46ksKZ0wlAKqvO5DHvZkPRls19fdD+14M25+5abxGMn76KxNmQKgzSJBJmmuM
LpK70YF6tzyX0ytGwtZ1maob7jTA6TC0ce5Bk5IsN95SElTRc/lUCsIMHCXIHIQ9
t6+7ULg69RMQwPH0WHDD/bPyFIaPIuDp2tAzTeQe1cCamPmTSzcCYB+BRpcbO+Jj
Ja4q/cUCFiCPyl/9enCTTrCY4Xd72UK4l3xeutvNWU/IPcCtUPmkTyya0HW/4Ucd
baQ9Guy4/GihyYQYdx8Y/9cff1G+GHAhi0gNyJ21RBdZcTlVrrtvu9ZDUSa7Vr0w
N5YaLc+ZjOVWMACMLkuseDi4uBzJhn9WNL9a+/5/p/Zr2XMke/petingfkj901yP
1WYVJBelvFL/KSKeCzMThacdy8hTYj2zw1Nd7QMCPYNDRpPwH35DriInXJSV5s6M
uwEPDCnnhE2LVAaxqiWaaW9nlV7os+azcemnhR4tsURptBw/AjXXAXvWcOVFFERy
YUlLBf/sUinTvQC8o9smZrS79NYzpJnr3V44PWgdxWYsUKBNOsM8wEg7lI5eECdr
4VBugl2ARgeEbQuzJ06BzHhJFHijYwayLLuBsyV4BdA1JlLJ3QGOP3fwcVwdkzmy
sHmAEjbe1rzkcvys/v0aL6usDYJbs2ESoK1GO7c2izSvwJ9yetevIxjsJnwiqlNP
2gnBgMHEIEiSYnIO05XZxBRRFwlWS8YAO0coQoapPxoWIYyLYjgG9XpVGziYQcij
xj37sw9soGRBuNN1hRwjY1LWQ+Hy3569wYS5nCu9/TzYk8gUaHOVgeJxJna6uQyD
fEDyBlyWKvrnNkmyTbSzO0To0UNm57RcyDuSVsgoIOzImqUKPPmFmOtLRKwqTVr2
8v0TC5eBcvU1IuWNTPgzSugwptoXsOSn6RG7AqWXGMcUqNMyHYmnv4sclnsAFFgK
mZwgF4hTphpqgae8Jmuc12rlkRkAF7RV3gdeLrkQ8Rgzx/FQdn8w5zym3NHIJmrj
aT20f/leMP7lGsBKYw1X0Fj5DCKXywElg23fLPc2ZR72OUSOy3BP0I8jnltoOObR
yr2Kq0ugOLCJ71U8fWA1xIGYsF1I0YTCz/VBAbv9jdvVq8nKopSsNQO8ZpNxzQ1T
DBbRDapxqDkvIR1Cg9UsuIxhGVE4yq6rg3pGeKVzBi/uUAuba4ZGm7U2AZUTustz
hEzs/OwwEBnL8ftbe7D8XMYOePXB+cTNDo8SLCjkEAaWLwf+FoUQFUio4WeFJXZX
eNJ1PlTUgjhMSS0OVquesrNFB5HVM0BI23TO5NIcJHNTbH66ZxLsvsV2Uvra/XgJ
p1hSEfoD9KIoU5WB0HfZKyseykUxL4gpdFH8LbUQZ+hdQEy6F7yelzHvd66bWyTs
ctcffCI2o67f+WXAoAKSOrazJ/HKC1xeWo7EFAtQuT8NU5qyreVnuD079Eq/l5gH
XlOd+av19BS+9OjDjiYlosZC7HwhycpYkMN1EU6Igu1L1Rj/pCSlJgWWsYqkv+L1
XOqjxCj1YxDZV5Ve1OdBAQR39hdCLRCSiBaOCA/IPKmzup/N2OGKb9b76YBJ/tPJ
jwRZazSGfaCCbG8h7jFKyQwuwhTJhtTrjazgBTzC17MI7Ky8MTHH+rjgVe9ubQRj
5+B73R2n3WUXbvtmt/6Qfkj8wtySYFT/9KCjYsg9OcaropdSa6pHsKWxgPrpZwJ5
Sj8wbeIBUQJhMvq/Kz4pzAeDfkVKWgTgiNm02CnsLjivuyI8lV/o62+R+8WufsMw
YZJOWBKP2iwR3SFUUlAAh2qXAKEq1/OAkW/QTfTuo1eaixjQi3x3BJoj01jCZsI4
g1yUbBnPjTf5o2iW+d743nC81nxbDojjZacjaFFsFTBXeK4hT684sKedoa8jehIX
pB3LGQDVYW+10OB9HODypFAUV+UIyDB9Mux4iLaR/rsJph9fA3xwP8BqiT4ECgDS
sKZUFzFvZtK6TeNxtsMjlcoHSGSxSVlkrLhd4ocux/pV/Jowhm6BptZC0c7+iS10
ELMBDVaezFBEiHIndgxGfXQkMV4qqiufMsAxUDxSJpW9a4nFCJ6XYc+8/Dzu572s
3tvL2WJ5IW0mxQL1hutrqZlt5JmesqQ91puh9H8UnHNgPKn/0hoxd0YtkEUi5k8N
yFnvFFLNRZU/tOIpRGqCyPLMPwoQYEZsU7AkeK79Fr88XmQ5Ji0cHAWuDOt7Sd1P
exyKHryGTXx9SSTnlZtc2JboajzL+4+4sv11abYXxWlNMyfIYeG5FYeEmd653AGj
q5IfA1eiLbRUBRjPHIlwWpZQZ4CEiKoQIDScr9TIdJjzmqFTzaAmk2O4OIpwk1tl
0LcF6oQMHnKZYuJpzuGwRlDB1mcg8ucy6YUey/IKCsCoAVsqaQlZekAF8EgWO8Tx
YbeYlDCasimxu/bDWGihwnebBtHeJMR9W6xx1UQle2TtqkwgOXz9R/AeRyx1v6lz
V42w9lWXJICVy/Q8+nv4rnEaZZgMi+38LN9pMlSFp7ysNC/dtWvkeFBpYrgR4Dbt
y/ejWliq8zqTpQ44HlKoiotIHXTJFcJtCW+Aoc9UmvswKOUQUq+NSbw5IIWxKs7w
+Zvw4evFxlBApxmrfd3TpvV9Ox/YAJwQCJ2c4yEGL8+nz3x/z6eJFu51izIaaUPi
ApTi/oZTvTaZ71gexAt7zYjh8ncX8MczeYKSouClPwalxw81xpLeifm9vBsHu1na
9Gcve7I30n+pzBVVMjZcZrIWP6Hl0nuaGH0vw6s8aXvtNHgsjcAKVY12sQVjRg1Y
FWu6NBW2qtuFQAFh8lxo4uToBbRdUHRJOpAln6usxUnXOdLiR/EsiAuMjFdVeJGw
Spm3HI1N6EpLZ5R3B+NnilyrDF2MRuIdKGXDFj4XHu0T90II7QhnXadnlvcX1xoY
k9xfZ7dXa8kJ3wo7fzRpoUCwWrEsvXwhHv2cosA5k1W52KIY3nsSF2DFqmBDHAC8
yrzKFOnic5aKiIO7jOA0BSBYf3vY7hNm9nIdDNLNgrPkfDH4KXfNl7SqzlnFcfV4
K76X1ZipqNXl/3oSg6Ypuh9ro9M3MoNLf7+br0yVailDyQzfMdWgnvZkxMebmlDI
5aUzgp9A8HgG9+fC5D1YvwuPtOB5slR29ZEULLVIaL1kYzHbHNuhHSCyZsDPuvYL
2CuzFqdbi3uTe3GLqJspIX+i19PFAE2lsEQDW/IlTU5H+ItGnaEcN6xZVUU9tRsJ
n0bhSHBydF9JK9HauaIPqhq1mzDc2Emb0W3DnACIsipH3GP27J4iFUba8dM5swf0
3b6adPQbYNTUGJqYH64qojxlYjPuf5DXX6aD5GVmOWIUJvyfWePyHtN7FB5iseg0
iUJcL6SxNwt3a1vcvmpSmCu93byPnBUge6MZCEhrcQvLct/CHrFH+SzDr+zlu9x7
TQQEFKrxLVBrI3RsXkuQ8KVr2T79CgEtOTvh8o/tmNJasmPe9USO+m70oE3nz2UQ
KZVHqOoxjEr0K1v8bgFg08H+dCzZU/nkX+rMomwCuRIwHofkfFr+oLWsbd1bGRH7
uJXeKDeULnFu4kNrd7mehIKqE5aQgoINySdusecFVbdiL37XDcwScHWUPbGuTqWr
WLkaVOcPQFYkS+083Pa3mMCDq1uGZtQFNVp6IVsKLqmVRYolleCjtoA2en+aGhx5
YOfLNMqaItnw2MiDUG1wASeBqg4YxjZLRJLtautEsjkz3UQVGZqjbEmTTf3hUsmn
fRq0B/BF1MZBhZ/tN22dv5e68kBAAWNvdvrBQlkiFwT32QkU17r2x1JtrrH7zpTR
7SEB38dz1PBgWSOKX3BK7Q2fXiPJRwgVrpXB6M2J1SqXT+D+mNyrvAYu1U4LOnnr
jOenoIhBgFCZPyuk7zuCEVo4G7HyWgXSSUKYIeMww3k6M7OpRQhaGCwFs9ZY6nZG
ThjoC08CQK/uu/Hae2SVG9RYhh5ws2NvfNT1xqXfCCued3ZuBG2oSUuE7mKAHZXb
LwCpFi0+qlBh2JqvKiSOFhjC2+FSvlxF9ZmgomLqXpDR1jq5MMKIlrlFXwNqYXLK
Wc1RNPmuc0nUoywW6VFEja+ghtpj8OQz+7zhdFtsPGu/Hi0IQy8iIddDzHAj/U7a
y+WKBfVE7keyGek/slgyVfV1dIl4csFSyRZVXdVdfZtUrqZLjdLxsSOcxMQkKaNe
Z+TEBMj2y4odCLMiMumu0v/HjiaYhzMyQKrQrlvZ9gHJHU+z3q22JcqH4Wx/8ANH
AHoxnRsIHMMbF7g7QvAzMCKpoU2e7C2nwSu3mth5Zc7J2z2icijzT/YJM+2bbMOA
5OpaqJ2454aReKRW99oT2y46XfZQQxRUjnN+ocm8vIhHi6wUystyEe1A926WTyiM
jElLhetyPnWF4KQiOVYqohE4p18DdeKAgFt4mkk6UAYjs/W3IdeswpWUtVb3XbC0
Ri4PTR9qaoJc7UIObIARtEuqhxPmMpIsQ0XaEqEP+5pcjBX75GK1U044MnvZp8/D
+nrimERPlHacxte2cKxBhvXUYmKhkCYvCjFBFX4hAVGBhCH2Ba8HvoHU+KlDEeCC
2Nd8NqVt42cmgQdKjbS85VjPrZtuG2zVTjAnW/fkzmlN7Mz0ltO87dWEZk3UHjZV
Zt/c+vBar8mTjTQ82HPIMiQfGqURXBX3/GcW2We16iBPxgDN0TALSaLhfKD5CqII
eDMTnZz5pOoweQQa8K2UKOJjpENPcDvN6xF8sB9rzNGIWnuj7RK/T3mudEj0mp2B
y8+OF62AW5mXs9trxIbIJmXKP6qtQUTGeiLmTilB1Al6a1Dd1PSY6W74zix1vNTZ
BUNsBdGOzibC0Od4KsFQFsae5j4/QaPZgNkfBGm4xtDNTL8e2qEvvENBoUxifDyh
mLUMSS9j/nCR4JHjgRPovvYlpe7DAJUlPsnOhGs/vF7jJ6yVIGwzhog25UGjW9sU
kW/OdtipfDj+CNQfx0IHh2khYB4dB1A6qiJ+VoY5tZ78sSD2BZSfUEcovE2glVwN
yyv4rR3GGtf6WB7GK0/u3E2/BYNi6s15rlPM9f2/PTGRRC53al0+AfKgVFpRkbUd
BVAgEM6TJmQQAOvlHzG+c9Ak1vgTpiJCsTKfBGw103Zz8kcq6S93XFoGuXjFzamu
5R2ZUilZPSfbqLgbbhk7+qsvC4FMw8bWhjVpdM38EcPBP07k5DvSy8Ty5Cb7dcW6
adsvrqMU7iQQ2JzG83WfmqF4XvxaZpdGu3jSZS8CdVuQOqkDyoZy+Kv7/qICQcM2
Ta6cPdXqbgF96U7fMPPEw8Cmq7LiJX0BriaZ5U7s2wmymwDC8QGQmuPYQNYp8dqp
Oi+nr3AAZBPBsd5wQxrC791QURQys5n4rh9KX6wtQgtQIdoF9UkrVALdrImC9kuj
ZM+vhnopAsnz4msnxp1NCIL9talczJNX2pEyxlB+3m+VduQmlOmpapOEono8usdL
jWePSNhFy4LjePZlZ840iHUaVtsP62OZU6nV3Vsq94Q+1ONkJJGPdfP+RfnFpoj7
7W5hyQyt1MJC1vpOgx26RbWx1NN5aAhcSqmsJQarUf3YguXV65DkKtOPukg1aJQl
cVIupFkDRJsvXLGj0ABNASu+aloLKKmYPhgpRvEBtyNz6ye1yxFnEN6hSawTu08e
Jpiu9C+lmHnQQ5oAzpB6NpY901vpOw/0dAQzfJ/VRbmZwLHv+9MaZKdIvnpE8edR
X4d6IlLZfx/cLBPNrZvzedB3VeuT7iCevyr84rdijtMvGaXtEDB+jISdr7X6AfGf
nCvv81p+Nn2V2MzVxWSHv1pjoA2LyJIIP9IHE/k0XnerZWqtzJ6FTFLksZWATjBy
n346In10FN2SKturTQTQ3YARO0ms41Vx0wp1KkiYCwUUlDyNVP3fDZaXJbW1blrP
ccNiVTpnKqpTABqZbsGZWhYIt3Bhq045fYgMN1xKMlXQkpj2IJYQ86AsFXqIQxuA
TNcdRgqIobsJVZZghZDLkrPq6fyDCXPtjZjxuZkG11HVGvPI7F8esiFy9cFHrqx5
/WL2Ny2H1gf9CJ0qcazqjw+0vqIMDHIYoucQebOq8M5SqdDQkXboYgPm1QTaWdzD
gE7OAKZKPqjWCa6XYVaHVX+Gj7wK/NsKVgQ+4gd2pAs29lnCrwmokgQrGkgu1fLM
VveYH2vMRruLhc3XqdHbpOg98+KuFKBvvHJHyE3+/KuiGUyiyVAoZu1yfTCwjXgh
r3w802LR7PClSt6wFBp0LrOUIwZgj1TAO54VzdNzyo3wzSpjl/HPeIbGM57CrPRT
BFKC9HxfCxGL43FH7KPjmQPvDrs4JpXS8fO7zOcbker4IQ72EtCoWhyPn9Lz+Yc8
DSl8CKVvBi/RJBadkFGK2HiAqeDO07zV7spLTgB8vWR1cJ1ipVsaXkn95O+hZteB
NcmRCRcY0oKbwCEpJGtBQyReqGh45TfsiN7oEd67UMttSw3K/ZRw/0KswH1H9jmU
VqnWt4FF2o6a68VInNZPtmW5oVOrwYYqU63StLAFmHqbpW8jRAZAJhG3gkbm9VwU
/xbmnwjqrx0E9Fvqu/eHsZShJA6TqkB6xCDK16fxyCwUrkhShbREcjixwpXCXeJI
wygARs7gvV1bMYINg34S7jo2HDmXgatofbWMHLAlN9FHy83vU/EpIn+KV5/qsCqu
qBiyN4ppxhkWbbCof/INaCNOv5YtJl5dXqgkoIjpQxutCXFBA2wFsCkDoCOvMAqw
e4IjPNPr5++AHCeXmsQP890qPLxEtvalQH9c/7YffxIrXjuxEO6hUivgl8jbWCR6
F3hsojGfYp4ud1xCDKyaW5NaFShel/We+xd/oLguVHwmsv2/JSXWPvQ653nMGFZw
SOGaFZ7dvEV67h9vUVlue1JEWQk08NOQkjm3i+baq4EXuq54a6JUOoiNPo+Fnx1J
+yzIWe1RTZ2PvbG+/54kC4WXoTNA/V/rI7NDtkvi8IbI2kanuEGSChd6VHAb7F+w
mruc2MbNRLmys5IsOfJwUm4h5Lk5BH6++/WLNNVJpCXQ5FEa0j6fdgQBisSoSm0u
yVp507FhCGVZBXuqBfvu1MMN3bn9f0g8DFHyZSx3WWMSdnDoIXyZUEG3/BgJvsOW
SUymh7zEbFPByU0ZKVk/vYy/wo9CcbFxxih9BQObaGXKhWsvZMh3tui1WbnQ1dJ5
9J2q0OMVsPyYLKkKmFx7wQBNxPETjsx9P8seO20pONQmc4WLZiEta06Km77yU/7x
dyhC0JBIBSW88Jtx30rOvAD13aGpblJcnvS6Gs3cLqIRpsqBEvd6JhV8Giz16MvB
m6ZdKZyxBYlOC8L5laazg6sHx2jjsZGCT1mWIaxsriAvxOTN48p29AVzSud3XwSU
tWJ+1JTPWq/OH+suMwdkcWBSVJArXqZlCHRUI6o9989m/w92JS2xtth5btni3V20
Ue09nX68pndbmYzs8r9Aa9gqXzGUbXfsdqcn6OM2C8BaiFiGQ2cNxNZCMz5v0sHl
Zhqfesyv4nZnNY0pZH9kFZsWAA0roRGeYEvmOLd0jTNAg94y1/srs8bnsDEolk0c
7TFpwQXfrETqypVa7rb9SdxAEvXmru95/VWP+pTRBY8zoyR69hMLODT5XTZTA6os
utYOxKfmVnCWhraCnRJz5SaSIKzh/AZLTqCrw07/qVvFmeB5vG09lEi8KeOYgeF7
7vn5UeUlF4xSXWfqwFwurn00aVbGS3cbIz/CvGdkU4k+pIl3d1Y3XQq25y2pIsZd
troYidgr8dzYVkRLKlqBVVKVvSELd1ymUAoEnTujf7BbMxOSGdLfKsOsx3SC3KM0
GOqufMECskSGJ35IejZbqr2/L4t3ptK8KBEhxq3yn1bsE+O8AuyV54lZ1zEf9z7B
/nZ4CcszDssxFPjeIdSTNGN3q5J6VQYULjd8W5NfDuc3vyAkqbwRIZbqQxS+E3UB
MxEF3fl9lPfm0y63sBuHVDsNr88PL3yeB32kAONoUcnzLHA/pP4ToQXXZXK4y5gE
cyUQrcKr5c4MjVUMld4vhR9hl0Dtf/Vn4u276sQBZgjduscci34d6hKVCSbrF6bf
xz/TOgHKMF/xDeG3crOLjPtU41h58A1rfz66C3aOLbtI3Vap9ns1cpoPgGsVi6Zp
z2jcWZ8FGxzOeYM745CU6STKnmexmu2fr+cEdN1Tcxl1IV+f3AOBoCdHAgaAaLGA
8kvxZIG7bI9ekudxsVc64yHBHqpTyVu28D94CYfma1jA1TgjjFGaWgRKfFvIfwQx
MN1r/yJgFe3N9+pEfJhE+15ebU2r0n0+T1H141tp/pa5eDa6uVyR4iahJH+kdCQE
SIJMa6oMFYvls+/APLsY7HXDpI03L0MjeaTc9/84gmXpPHJga0qjnudeLagPWb6L
RTCQCv92sSwq5dCkDRaBHdZmYaethKaKPVkwbvgqOZi//9Z85twcDq9YZAWSjiXW
p5AeZbcV/7uxdGEOEpOjNMjjHzMjP1xpVflvWuiR5SCn15/4KRfyURdaKJ8lLxNK
a1x+FaFk7EDwDpFtD7WDB4mwJjpEtVidfvkWa3B7ShxH/zETZLRMlGd0fu2BWDrw
UGb+kb/GxvIBGz5xS2peY09hjS2Sj0dx4tNXl7ZJw+FAD0W9yhRjM34JVp3jsf0O
RMh8PT2n6PNnFFNYu+XmbPf/gUM3629nWy3Iv9Na6jI0CcWV5SiGkJ5nnNBQLqfm
mClGKu9F61cEpS3s9VCdnAImCs3hFt1IIKsooodPBJMfeLoSFdcXMzThr9brjZrI
aZZuNW2T24gqjXloBGBp7VeaJBsPV1koJE6u+b60D7DjDh74WuQPQX4/jkbQajHh
1tBHyAgPtH3OoUu5yMylp5wPTr66IQm7KhM9C3Q6caKq8PRBAt8QjT9AaWNP+FgS
+BKtqexmp6snZyySdcaDx4XH3SXDgnZRfsGT/MbaUoRed7z6TqBn+cqqEZ6eoKZX
dwG8i9MbyVzXERBBvVdeeWaIqScCFCBjJkHehJJ6XNFjhTFEQqTZLA4nE04fObCF
bdfvLDG2iZEny/PotYeqZiraBw1EKEIvVFXIPOr4XHBWt7eYek3g1hQNs9AQazZU
PCzEZDAUv+tciGSBzfR02K7RX/5u1R+3fwVYXl+ThTZhym9XxFaXVB8Z/CQHTbRF
yeW8ZRaXKz94GNuDzjvXRYWN0ZYhm/bgzY/FzZAPJ3CvvWCy4bWdc7CKTy7NvpBa
Yvu9ymlvbPulimH4P0EbyLyOyzKdSzoqK7/JHDGzAn8UjzMudCaZHfmE668rw3Ly
3MU+4Zc96s13wSoew9nVm0lISq7Pz4FZ9rWtkePZqxf0f2wBG0DxXNHOo5svrXjk
Izsytfiu/eHPiMtGzSCZt+XQO5vNTlUMMnTqHqSWxi3jDP3MT0i8OHe4aTaojyS5
qt8oAbZlGWrH4rcWDwOzGEQmhxVpUgr4QuCV+4V2oIuzdNl0qBJPrDjLmxoKHr0u
tP7vbJQDuz5RTOTxn/MloZ6t6IKSnGgBVwQ5/iJrTQFC901LQTP+USnc76ii0xdz
EhzUPKI3zK5kbsNaeIFF9hwF2jhn9rq4DL/jMcGtpY0IkpE/PXybt/PkXS7MYA9M
AeGSUA8uwxwa59H5wdGbB5JFNkqXXPCbFIvs7vbiWG1v99Fy7cdv5m+S2W+zNIZ5
UNC7fY8J/fwpIDvEdL8QXzskb9AOOfECNb5hfbLJLvEWXchOzgMnY6AMvM8cYOCZ
Yl5Ymi9rO8Lt4R3ZfYkfMbe7sNtuljAZ23vXzBmCtrnu7Afg+ItlYw1Cs2LoVaXE
zprc5psWKDMVCGlUd3EVpaadIeoxH86ZyZuVbgOvBjKuSpaxY3WoCUU6CFfhu1TA
Qrax72qy4wiCqd+pmfiEYiz1FNM2sn0cWq2Iuq4/0Hkt225KCYlMgY4Vz/gR/b2q
7zw24/bq9CdtcgPCbcuKEanczmgcKTMiOKEWlFcGUtqcDnA6a0/owsb+8baMasmL
Ss3BeIjBCOw/p4Lc8QgstVqdQye9tW9nw+6DgluPyUb5I+MDohfoHy1hOIHnTkrK
/6QyZF36Gt478iMaSCIjIjxHxb6CTDbp4Qw0srznPaEKIU+rD3AnJ9D9k1aBXdQY
yJyQDDyggnhacH0LOKKAJ2zYfarHUhj0CihLugubY97uWCZw0trdKjiQisjBjama
++i+8uZybBiLK7WDLmCju+n0zrc8+8wxWKunlowKJIVALY+3A9IvlQFyHsB8TjEF
mwUjzHVQEhiMacRk7an2TZeI0qbr/LWM0E0y7VAyB1GQ+sigpZh+ktAQRykWz3za
f87feELF1UMfKQDyQ955vq6ftMqxSoDqgklxb/oMnrf6TlGaelZc/MJsLFTyXMQH
76VFJ7InQISXcDr9iKiEG8dbHFhvoVOxISZXn2nEk1v1/hp1l6AuPAXuCQ2fZEZp
IVD8Q44qGOx5r/WK+uW/qylnTWEaJ53QfwUrLG2f3CIFc4NbDql3zc/ubwzX1SWo
bcQjK22LgNuZ3xCkfo2wKgE0TsZv18pvSbISa8H+3kGWZUYX3Cidc984inZdPLQ8
+OEMD28ZMfcntdDtjr8LQ0ZqYS+QhGOdaGCTiXsHcD0+UECWZiJ2QLbshnEshHtZ
YEO4y/rLfgK7Gwo/MZMKi1SumRrxAYCXdF5PYx2pA7j9a4pvkBquiN1VA8cR5R/M
4k+Ejgt5SEbT4VIjha3S9UI5KJIK52eGVKroThzvg2NGEQ/1dxENxJD9a5N7SgrA
+RUIiJE3wAqX5v7BeeAdG2fpCqlMbuQmyTksIsGFrb+BSnBG01Ol/rZh0TLHI5z6
Ukfl8PnDVIj+n59xV/jQ8Dwyv0TeVvvqWxql9MBcn85LQJHMKp2dPS29HtTuuAFb
V1KFN9liNDPTVM4N9X4bA4qTSJeQTo0ThsA7zr+sMWJt5Qv4mOWWmTFEvJSHpEEM
kI1cqyJjwtae5NUiTX2lu4XPhKGzSxpMgDIhof7+4+Kf3SXIBZwOVbiqF8yMy920
DPD0n/iHHjzMCQKPacXKd31ms7xpfMBP3wSLzFopbfmGp2cdkewdlkYl6UMUlLZK
X5UeelY3vBNvVbZo42DMds5PfKzU1Rjb/n6/s+lFAu0AGkNr/yHAdYXA1ZxPGg9S
vr9DujaQmHzyip/tI4hkRcreSw/U8FlZin18b2THq/+IPlh0zk9yY6Nu99yogY0D
i53iOgUStWoReGrEBa2nDgDB3BEdXZh20QcRFO7WD3SXc98+HuWW60XKYZdZWpJ4
QSNtvOSnzvQt7MDmumRvV6HBPJV1j6SmUH5ztXCP6JcEMQVPZFEyocWHEbbta4T2
aa+wNi/S9V1pAoGdV9nneyDqO0GaeamKP6Irw74BtNIKEkFhSjSo2T+ppM2EhrEJ
0wzDKX1+we+woj8m5XUJSRqR2JXaHtl0h8WLW1IEs8JTi1n5y3LrP2mCgfhK8WDV
6tvdzLiXfAIhpBB3xcgoQPZRIpiubROBuzdArZWLuvcd36sl1P2pkqnNBYfg9u3v
/tLsC6y8rQ4O+5F29i2DcpFVxxa+Lv3QL8OQRHCt0T6gFQavfObHF5oe265DZIMJ
DPq7ehgP1vH3C9j9pebWmf/EPZfen37+1l9MS1TWWzho/CP7o7xPjDGgO1GpBpLd
pgMLedeJD7H6b8iSA2tO4LJrDQ4OGW/RGute3rTh5H9korU3WrW5vkMNpmZ64bXj
i3pLnh1+/2RAJo6C/PK0I+1tuFd6Lx1BaWRlwP3AMnuJab8R19w0naOuJwonrMvL
MHHA2mFN5BLuwwYOeBO6B7KnY/PGnu+EfjnEqwG9CLEMqasyvXx7xQRHe34+kxe/
znkGlu+1o9PB7FUtIiWYZdgmFa9juQnWaONA9+CVYQtSH+apag7MGnRqHFlEV2el
/2xcjEEI5uPyefiU/UzSclFfmL815GkFflzEdQEku2fJHot1k6OWhQ16BZvX9OA0
lT4wOz0tQO1KtKkkL9LBYvAK3gUg3eEz48MEx7muP6TiHADC48Nv2G8M2HQNiBV+
Nrqpdj/C0WNNPWIlu2x9uHIVuswtOr6A/vDRfJBMQUoGz8F8HzEf270offMzoXJt
ukBfMqgx7J3ZSXmBy5C1EITvmK+//2HhRGL1drCA1k2pBnCFwbOd95I+xORR8Qo5
GzZGYhP5Ad7Vmrn+NohIVJbh5kGpqeRGZFFahpPR+DkmVXdQuKOSwbhEd1SYVmpk
RF1Mf50RQ1OzzqOS4Jy7tYPwCKz4su4iDva5XnHkbKXavc3402xs8z4bBzErVGp9
lvF5vctXsSzvFq6yHDpV2j82h2fNqbxMhQ11zpZ5gat5TvEz6W5IbygJb121ZJd7
445QyLBqEoOc9ce7GuRhklnL8JePMK6IsFlXl9O8oXOrmbKKlX/FYOIj4XbCG1s4
ST4cbm+nhY5+Dfk6HqqT61/+WJE4JwHeKWh5W+m2JatDtN2JB4xVkq0yW2go8UHu
aQloNxo0q3suN0l3JE9PYtiLwe2uYCM5GAWtWSoBpraS4H+Y/A0ulX8Z0+I4Y/Wv
e22ziSchhhJ7A4O1yYvsgTR1VihTYD4BikE+xW2DdBtIF7oXtJcBLjGIXXxoNr6B
SE3klTKft4CW/wz8TRuYtsAF0yvOV26n9nmID0pMYL1j29ImFUlmAfzUKZTtCxo4
JVUGr4XmgTTpn8j4FMgpZwXl7bTJ3ljI78PPVV2eYH5tpXJBch+015s8CZuZ4KcQ
pyHrSXjs0NVLPMufSzDTaxWKq+Q1n1RrNIS2dsAsIZ7NINPhH7A+i2CsDNMhYuT3
u9007ZGKmkHioMIszWTUBQSe31IP2OV2Ew3V2qleI4LQYvc+bD6//fWbhnjrIGAg
VCnwQWIMHV6kaiTR54AVZEZSPcSpjC90CHKnr4Qeb3DFlhypCL3xJ5EHXjBC4Py1
M8K7VvYtF92G5HJpOUoxrqQxsvfVFCfZDpt63jyolp8RC/XKaIOXX2UUIwOxjFpH
aCxDlG5gXiP9GmENFhcjFME8FFJeB6OW8P/K3hn7F1qVrMHrGuWnb8CxtlYlto/H
1Xr+3p+MDUVYPTtX2Ax4LsVzA8pAzuvZBhW3/OGTumMWsnh9T/R+c0JW90F63ZSA
BKvTPTjsNlYs4PXfWxnktvJf8aMsvvrxG74lTEXZY54bzV4M/oIgBwfE55GeuJjw
aR5KxGWoESFW+JSiWu8EFx1mqa9Me3+Q5mZKOXZrybjIx6zHGrPsaERBYtJWN52r
AfPxxo7XOdOLNpSZS+J/WOracSwMPdRcDyjRmLr2P/LYeSfAAGUinjPhhE88OvWF
Gd6/mNJ6JHKyflIQfU9EXCsuPD3ToNroDNm1XSpOQzwabs897ehVda4zToTUjHdK
ymC/ge2PuXyqSEkkLle6JzKzX7E8Epsbo69sCrNwtAKWNDi+PpiYSb4Xqal/jKmS
FeOQJf2yTGlb1ezlp0srvp+p7g1yuXeM2eFXevODnu+jVan8l29meqK4ieolWLMo
9ozSk2j1bXPoWN7hQb/91mAUtx7Sxu3kIfEnoHwLmhdCSgiLH33HPQc01of/y4te
iUqbRzkN8nRb3fiC9p8n0wX8YRU+K5QF/NCQ70jQDGwe6+8ccaosPIlAE/di1hIv
4rmUQzLEZHMppzgSENpEJ6AFUfVNTRITyvCtJIj02verJfzRJpMS4Thy9OPw56Xf
vM7d3LyCmENJ7UmC4tId7fV7Lz4qZbugOzhMbRtaD+tGAl303B9zin6fJ1BTuENH
+dnRZtaq4bYyzgum6fFSk7lzigiqG+LNuXfoU5aX9P6iHjAXnKwwwaj/Lrjldu0b
EF1mt3Y+2N83Et8cR645b5gEKe+6J9mIEh3TcmcEktMQggo7ExKMBUYj0eW5hhAj
8e8YzVbcxKGn4fCkG+y+MuliMhv45/RzPfrVjtfAxGMecYSohk4eBX3X3YfUdqzg
MAq4SmVECopHILBzWdaXLUuEhhivLruCeHrD9RdYf/KvjC3zfX6fWHzS0YWoLSNb
RDoX16C8SjcAsrRhffEWu/Fdj+eb0/4pfmB3JVUpF+Ko1CXrIaNSkPlUZpAFWrzz
CuKr4XB/8ndXhSDnP3jHmtAiNQBG6zO0HiD5OW+xYMs2TWco2rb7mfUUg4xt03C7
Ny0uw6XEgcBC6eiRh3VR4FZBcXMjdPJtCAlOAjf4jWe6rsW1Kftub4v86Oma3C3l
tRDyKPq1x0NvSiPDH1A5xk3tvJDMkI8oSiBel4jhPKi1u74+u/5D23sGVJ4z3fHL
p3ELmVvJ75RzpPq7NyqPiW2NcApayhAzOsYYv89OInkZhFr/LXJXccMBZWfZH/BQ
LGBWWw5WKYwMdOz1ypof29CPBkKm17vrX81NJnRodx90JL7h8HSMYotagQyB//U8
STEA2c0503vFfEUDTyTvt3pClxnd/9qmPt/sFVIlTgtBIcOUs+K2M3uRWFqOOOOf
lS2MW73Ggfxg8H8ot9ReEsGpGlQqKhPiHrTuBhOheSDfxUlZn+Lw8xuNIFFtfW7D
kHGV39wrlLN7GsdLcX1uXYQdzJA9x6zDcwmMNsP3jZDvCJMu7s9GSo1amrTea0s3
Q70Qu2p2d0QDqYxaPYmNIcA5fX9c1OgF8gQIF1Q+7Q8pt/G/WaXuGO3d4Z4ymYUk
dyGe9q2mfIgj2IzOrCTX+tiQVp/gHxRp26VQZr/3ynUjYh5nrwaNKjpIKeGa1976
ofiDvlIhgrcc0ShPKUcsh+QcnKqD4gOczQR150qNx4FIOkzQcTe8iWjc9mycTxwL
O4SMZlDQxLK6awHM9sV2FG3FiAR6wdry9rsiu1CLl3nvnJ5dC2DAYPXlwodbKSb1
CpJGnk3tFqavwr8xDSQNhv/1ugO2pAqSBukisKbnBI/y0/1+a9jHkJSm9wRV6uom
pBi6AEcBT09BbgW3jEbzhaqwg2LPayIEvpE3L+PIVLyPdIWEyayUcoRAyGxHGFCy
I5a8hNQRTBTyzeBZo2WQaHApRvdZO6ygXqtFnbVM1YhDb7i8SMfVbG//byzhclDO
rFxVX8AjrjwZMaSr4/6apeqsFu4yahXrNNguV6z1/m9CIfcIf7NmsznCbTs+EtaH
lGddftmFI1t2gODMdY4yks2m69hntXAZSXKDkJ4FxIZrKWEIzuQSFltnk7SygjXB
JeUKIaR3QoQ4bdWQ48RMGqWul5/6mmjkdzMgjflp7PKZ7av2Uoc/x/wmpc3X8Rwf
t41nu0SxFTXQeDf+tjwJ9nsEpXtJ7fQvnZCR1InPoVarnQsWO5zFLkQTLcLS26ZM
ebt5pt9jAjkkoZEI/pxzi5x2Ke09QeI5brM41cCRRFpwIkmk8aZJQXbhnPF2mK34
vFO9IwIFFKe3SdqeRDdGMhSM7erAklUcXkYgqRTMhh3g8eqZPTViG24l2X7p1Unb
ZgyTx8d0osqxeI13uct0Ob7NhE933bV3VqJupYH1BcBXp5Yu7v0j8jNfQmmHINLl
OMJ1zU2w3VfAfWVKErK3MPC+NLKw2UNljK1pQecSGiT5ksptMqY2h5xZ5pjfTRNU
u74YNwtt1uEqJ2c1L3A4Ocx5d+6dfcmqeHHr0E5DeB20GCZU3AiqY/ZpyPKi+biJ
y5KcA/ZKD29I0FZIu61PWOQc5iFEIPriH4HGSL9ahrKmTF6S6F3+FcaHOoYuJECY
fzbIc2oGL5XYUXPKyphmCT8PS2V0Zn15JMKijk4yPsFKmPwp9Fr3kKh0Up1Ml2TE
nw4LZD8ZZiSozkFonkB2ga2lRpHc8XdS7IdtHd4RqZ4ik7u/fSkUGqmR7YNxVc7F
z9NNn/VCil0APXrMdSJuSGsTEqyxZ7D6PHiONy6DYiyYuiId9TodcT4w5uy77ygX
IxyXDJMKGUq+oyp9rizqMyRDeqCnpxQuaZaShurVQXQ7FzURi8zitPvfdQJ+tGCn
M9RuzAKYPsUIjzypLev+cBf8usnWfUa0/cx4SeR4UX2EJuWJADrTtC6MsqhgiZ9M
D7YIS9+C6xe8he/LfkitncrNOe+cRK36se+WhOn5BX0WzEshk1CG21QOLQSV+b8G
YbB3kAYkdEtZaQEZwGzWMrnfTNPKqBRq0aFJ9ipbJA5MRXKyR0EDXEqw3cIBtqxh
QgLnNrEaeecpruTx1ViHo4EbrFeDxmo/ZjYZ/6brM4YHV6RMTG5iYNg73f/BuSLO
Q1aLosEVoSU75nYK7WpgpGH5MsiD3oFothuLzU1SGtAOm6APpzWSfFKfjwQh9fWV
vtLKQNhEf+3T4OgJ7KT726eKbXt/N8+TqGnLUL2RrzoIxGRr63knxbqTCECXoHES
SGWztrxzDsw2naaQCnHtLPHe+8WVqnXJ0bvspOgYlNxC3Ny6tDo98sK7414csgOT
2bsVR38A9+0Tjjvv/HJFg66s3T7uEdtMJpDWcVGcK1ODX8v9LyT9tRU0IT0AbKob
XtYTtwT3sYz/Ge9codOclDHVRpLlcxIN3+bH3jJZA9bJ00s96bl4C9MSl2x//RcU
+YA/jba1+s9C3P4h3EbQOJKCfdYE84Je1WS1Cc49bohDPSeylphohN6YNpeFaiJQ
eqmIpqLH8o78ycNfi1uf1kt6nOmXoodJSCiqO6cI5jSfhHYPT9lSG9PPS8FrO19p
aojhyIe9U64MlzIKfOvz+olQVg/XPpgxMYCfRjJax6FA6TYEXOBH+6q7rVDIqXJ6
utMcWcPkX+/VNFjXDLgRG0DLqGAho4S4RpnXOanrhaXCAAwRDWcTah0tBOBTSewk
H4UEDaNJAwsohc83FtQzxrJhVMan9BJ0ZRmGCgIQ6wNBNHGCx69e5jCa0ER2LR4Y
GTg7XKxI/Ipa1wL+/v4JclQZyxVIzM3+12WG9O5TnKvvO8me0nEkdIHOyk34B7oB
LFteuTbndELKrNoOc+D9jOLvSu9MOtC2ONyKlGuU9lForC3hlNEiAF45qbKhK9yx
U3ontBUH/FEJMmiRYkDPnC+jCzTaqRLRiLhkUSGzIzKUhV0VL9HSFbBGOIbnIbl5
3APlasIfP6F5Tnsoa8OWlzwE1bSo57zN+6mvCilrfooK3/BanHiOAKnBYHk7lz2z
H+39POvH9KZJ1QdmFgHLqmBlPmsHeq/SzGm8EtH9LM4eRGpdY0/JApp462G6U3Se
Iyg36i8qGWUSemMjivixqfwSh3Mp16eAoY6e/0LsfqbGAx1OE7piWc67tMQn7Vkk
az8YMzwfLq0sp4b2T8ofAjT4CuWWYX10zUifDoaxRIKEt3knBJWR140nl1ajM90G
BLwJhNGUnGYnyMu+9U8vRmNXt/BOerkTGkSaUkRpK545Hi4GoMG9V1hbBImKZ6BZ
vnD3/DBEBPRsnvrBBKTb2eYyf1/D3uhyMQR2ucoNJc7CLpXRVN65yyMKaywduczN
jLAHNOt9UenXsrINajLy+Vpkk8K0uSKoBaArdl8wA/SRQ3yPfYLV1X7ZMAG7wg/M
5uP1hoF5ZUwK4AVLdtEN6IgKJP+Mgh9948szP9KxP/enPiqJNjcMI1pccux1pOfk
Plfe0CpOomAHYKkopJqqc9KA22FcjlnpomICNqwkpIUlvdJmgXLgBy6MFkzIaviV
0atXTi44YgNDSqdS/e+GDfTlnlA7JTH6CqiRyRInZGOyeEvnPU31e3Bf+7M4H42/
/0Ck83hDKz1bKjIpB6Q8yL9x9m1DzNZJv/RZ7VOGRlXNUTTlh8vcWdXoQzK+CtnJ
o0ZcjXtDzGwOI0R83362hwdccGFuGEBfA/1kkhCbZ1eb4q5XALHaC2LXM8yxYjX/
j24wuflrmJyIPq1X7B0Znn7N432sZXEHMp4hM0wBs4XZsJlp2sRq+ttluBkFaRsT
47xPWoNFv+ZeQnakWu6KsXDzWo2osT9Sm7PKdG1WVcjafompNRc6XddUL7WHSgFv
UVQ422z03MyBcrCbQc+suNMPNhymWm1uIq8lq9x54NcaH3thY1BiboJhZLFQ+gVm
BkZkQqNGxY8Fq1GjmsD6ik/fyquNKkvcwHvgdX/2uGOyYA/s+2dzcchBkJmRfQ2f
n8BiarMLR1R+oLCxtY9EA5XoypeablEmSDDxF2s+JyDTXO8TH2h2HSlVlqnJBnQf
6XV9kAdKSTxhhVZTYClpj4RmjF8P/YB/g1hmrIReK1rtKLmSa3n7B/ejwE+DXNQa
ldP57WZf57LMAog0GxbhXDsSM6fPZz1lgM27NdfJ5V4GtKNV/rNIhTIc60vkie36
EeySoUOovsE6K77wZJ7FBAguGr47cFZTobmB3w4UqzkJ8M0ELHfHJt5kjGQ+2tVN
qX624mYQ2tESltbzbISbUudm4aYCsZHsg7ete1qbAN+gzIOpCWV0j3SkxWEyKpz6
N91Ia1G56xJHIK7LcFHjrwQAKAVeug73Y5wgTWn2ja+J+nXqo4s4g4mAaDIgyspU
tCajQBfPDG2OeMRUrPjUSUTJE2MqCirg2YLtAhqyhw5kqn+vpLMpE4KP2DK717sj
if30WOiqjxOnxlxjdiJ98kiHXoWeoPOMTXgcQhn1WMkrvsTh/l7ie2UxUAqjEE61
WRlalqavj2Ou9VZQWHGe7py1tECBCCS+0Ld6LLuTGBcjwgApZJR7v0nm9jpwbfwX
c5ZejyTsgPnLrCgQ38neeX1OPxf6TzZx00VxLpQhis8SRsb/6zQ3WwWloEqnoI6n
qMn+NSESe+1Q/z7wjQR+oHVylS+O3PF57K8xP4GdeLkRMoH9XqfnLMhqkLeAy3Xo
gp1I+CgNw2po0hIDCIdiur9PIZlrsQcrB0yHwihqJscu4QOVeW0O7v28auZtpchU
bUxr0tP8tVe0qSYwNPvczn41u2J4KJlgt2vY5GZ0ggOXjYY+GPlvXExrz6yPtTMF
gjFrEQMNChitU42xOkwFmh6whC1fdZunAZ7lUf9dICn7mslKLj1ingh3H3l5Nkeu
KqHN909JfyLjlMCMjkTyiAjiq2YNUcYqzZI0Cxt8O+5JHMAfxFE9q/6rVjl+hI/C
YITaLk4o6pfS1pGZPuqucYP3oGWGYVsw7VkK9wSbOlWGxfFE61ohCkJI+x8368z0
UoQ8RyUJZYpwHQWPITEJGbpt0tSqUzYTdlNBwbQbQfBLWetyKpA5iajCPzfz+7Yt
9GotM37nF7w+I5jVnoDWjKsPTeDkFF7ce79Id+LTPzTr+GtWqK0hLyqMZS1CL4ed
3NRCI8cEsp/P1fGmR/lVioSKykDHM+4YveGyniwHXWvXoJmFiQgG5FW6aIeSomMJ
2bNcqbvE1qPmJJ42/VYiCIMtkDH6W8/gIFYbRdtjD+h65l5jtEZmi8KV5TzCp/b8
xRUHti5i3AjUlHByFEd/xyHX4nWZukMSbFINHJHpusfHJCgaxTrlQn2YiKG8op+H
wD2kdpJ0PG5H+L909Armb8T7t2ILZMNW12FsD74p2Ll0hgWehcg6O0rb3fEHfwzd
nbVDHMumRWFeYlCKCXF46/Luh9QLcN4qGEYOowtN6vsdza1lHKYLSppkh0w8fNYl
NeauNDvOs1XfEImCFl4aNGVg/kqk9JdOfLcjXYX16gcqUy9d2LyF4VGewUguI4ev
XFDd0SrHORiphytV1Q3iS89pDAm/OF3UkMteeCBQ7bSZzwDqIivLCVO5DHT7F63X
xHigqGchReEHB2sqowPfP1CUgghEmqVGfs0mFwlQsWWZEH4+5GazTnlS/pB1XUrW
PnGC6i76v1YjMNmYsJD7AlxiRMP7jENZCNWA98coek6YFD34mNVYrw2LHA12WVcB
mkORv6PM1O10lsvGFgvzx6v3A2ly/4RXiEzfmVOZJfhuIzhVkKpkp4LUQHAV7lOB
+WUfyyyPPWKHA8RedHB0kYWYrTtiLmRGBYXtEtEaIwUcZ6bw+5ZnYpCQwhyjgvRX
/Xlj/XTBdhRts8e0yzGxTUZHxzQkKjnq+SzkO01AVNawFnehIMJDt7AU6/ifFF0s
ovusyt5FZHTFn9QJeyh7Eht5z3243zXOUEAhULksigDjIpfpZRRokWTwPpEJPUJE
VakMQyDOgCItHXeF5LeREwgT/arAIgGZPukful5AJYd+KXftrvvrSgruNs6C44bb
E0A+6o9wCAAs95ORr54tHsUDJ2L1OqmXKrv+dlkbnx6OWvH+bs+2meryOGPm2CdV
V08d12znUFksR5FQEnXl+cZI1UgDJ06L0Fv8qWkkNKUjvww9Qjg6Buiv0WwA0S+j
2t74Z65iFKiDHupIwFSxfMtNP3LUvECGGz54tA0hxfuueX+OAzALWaFvh93Okey6
yHHSL2oGUuRvryZg1ItaklJ4KOXCN63dvkUCqcJq67ozKyHHbZWXIR6dydnGqlLH
gl/f92COXVPFe+w2tQx+aZzS9wQu2Zr37VMHPOHgcF6ooV1KVLXEB0FpCkwOIpAU
RYpcet1CkVqaXkGhhJMZITEaEr8JFehqWWjjyBsuc04DtLsuNqSTAAblTx1lDaXm
FIE/LjP5/4EW2g1eUZwpqYJ7TwxRRzaRlShHxFlLEsy5jIJEO7L7gWFBY+C2JnhY
Kkry1qfrJbwQmTpGJfEaUgnQmsqPHAfdMZg7b0KNfWqZI0rrWKy1Dwga2jVOMCaT
gUKDeJ5Q6Xn0a/rWFcKMqZJv6f8iHiRKx/Lde1AAs78awBvalVUG1bIKtxdqfUpK
tSfphkcE22Tphiz+4oSD6lnvhyL54GxZ80kuMuvKdK+PGqU7LuuevjrLqDVRGQRI
jrPdnymCwbWMxTlrnH3fzP9OOFAulIZOiO7BwNJM89zAuCW/j1bXZzg4Z7dPObPh
8Am9HCwUkdpIoO2DF2Jlo1y24UOaAE0/P+T987mZvKdQyMd7TXAER6xqroYrH/1v
YG1+YH7EvxnNNzdmmfN7PrDf8Fp2xFx8Dcl47HeKLSyXXRirOF99LAjTylT6puzW
6k4yM1lG287yiQz/ihrlzwhffZX5tBOknr2xgleA5FKDowleimSgUWNpnUNrHAlf
uRTvvGDQUmC4pYcWWQD52PKtD1LWeukmHcTFnrrpFPMwzP40tpKxvMqfKqNRNs2M
uoKknc4JwW6PB63litPI6iJfjA5Q4zGKYj0pAb0QZY+2s/tpl40w/dnognegTrdB
fvNam2x58m/Nu97axLvhxx17gCoNhALfWZpc3IC6zBLZHgePma9NBZvjuDhZ41bD
0Hwk3hbYno99eTe/EFQRktwnjAdnNWyAItjq4rLfWPnxziZFN0dU7JLB3OA94eRp
7NjKuS1ipnmwdPDEAyd+Tr6UIZI3R0CJmChkn9Vo9QsNJ9c1q6n1t77eQ/sGberb
J2IQr8NbgbvqT2nx/uptOUVs3vA8FQ+GacEauSner7rqvepEi8xQlcjzZH7lNbgo
r9sSCkQ4W4cZnWSAfYy/PqdleKcbCowajVsm7dwuTN6CA/jQccZsUyY45ihBestm
uadZWqKRzapygk7E+ovLNbD+DFlPLBkR9Xsc0elMYvCK8bpXg76/NmgnEabAY7/2
02h9ebR3aDRIqOTzOvMWtGirlD9iQf4bcXs1rFDYlntdlZwhPkI1exOGfNnrESlW
1/UllKvmwAa2CzYBmW4AmfnfMhGypT1Ivd95NT319++SK0ZQS1J84T4ebkEQIkVm
LX6VxJA2wuIPS9R9kKqLG2n+7UYbszzge3LWMFgPPSJ5EwneIzfleTL4wvdF/4nO
PdPW/cN67FcO0l1joUipWXZmlq+Q1SaGnWyVHnEOSh00xsCZ+9ZYaat+YyUUW7bR
kiKAcERcgSlbUUe9FOONY3+vuDDC13NzE0wUGkt+wlXgYIy9PwB1IEanPJmwqrzU
ixQiQKLZmxC4To8VKAyvUSjVfKj2s4edZF6KCf2KEfDSKafuqkF5UT9iwuu2MdfK
g1rYx29sgVF7Yg5MApj3FMrl32yUxcgasI4xCSEWM99a79fWVou2ClW3FsoNMILs
zh5X37trWgKL1oMLc6INujJ45M9k1LEFQoFczD5iqKVy4ITy5euCmKII9IySrgA+
QHTM5fzv5BUR01nuywJNXQ3kFwY/MM5aKNGmzxDN2W1FnyPmP/NfQPZHRRTo8vaO
NU37dT+6bxAFyJHFm0ykxZWS/r/N42h+WUSqyafF5J0rWP0V+w9htKlnbpbXsABb
G/Vx45ri0RPYhSp4oco8dZlhhzb9PL76snmu/kqTmeNapMHWrNbkd+wbgjKEaOBX
7wofTeMJFRRAajF/1RAAIYd9FsuYR2wBL5bLYGEedb0j2P/EDo44Cs2ZDopWcu+J
mqVg8f/6j+5cITnNKIh6jlnfMPAvltKfy/8S95YhVha+blMgxGJesRx7QfIB+KQg
2Uf5CqhOp+YT6OFTulKzyk6aK+lksm0/QSyAEmCXKPyuB8I47E6kO4N5U1A7iW+3
H5XBh6WY9H+J+ur5FXYPLlantbUl3hX4OAwjG1EEzHSIIiP/Ms4J1hbmx/b9vwnG
ShR2/kqOnqgOAP2cpYd4zn/sGLKyro5WaUyG2doqjB2K7OnEtnkTHl6KyYhh/EWS
AvkhEZ/RpgOUEQ86U97PR2E3F4wn+EEYiBFbuTa6alDBfHzJzFGscSbeDp324Igh
mOQhBMOTjdTH/tg6aB1kkieTWlSCiP/bOq/LXv9XAuqycGJRV1MPZlqSuMJNrvXP
D+ydWoHJdJ3b0Sij6f4I7YhJipjiBDi4NkYHQGW+KW0/pSaCxhe7i4gN6vAW6xv/
KU9H5oMbh7+EoeKk8ikEe7wGDkL15W69AS8lxLaTbZw0zCocCfDB0sfzIYnz5vtW
z8J1cW7nnLTnF9jRWDhKWgM6hsiag3sDSFmdiP/4jEm7/16fC9rs0OvSBuRzlxx7
mUY32pX0i+6MuP4yDUlUzJeJ3O+34IL8NEW2SPuIGZXbT3a+tJv6ONmmCumXRX5u
MjK0UqbyWn/SW3HMKwBOdvqJkRu79YqowZq6Gn5+HqihzNF7n1rHSTgvtlmcLWnw
lmKAan+GLUVmQai6j13rBBcLccKwZZkt3wI7StK0Z/hArc7AgddNWyUZqEFuTVgK
Hy7yDSunLaKam9LPGd9T870sTRedBpy/o4uLkzj0e8j4zSMDBwVONXvfqgvTVkst
3/Bj3X+oOiPceJJgbP8mYPv3qkmesupH22mmYfFzx4lvsGfmPcX1iSyi9V+7QgP1
XktmfL5N1s40jJCH5Ik0da5rERqNd0U1F3IPocpcl+pHkPcnF/VvXG9GeNQRll6N
4oJLooBAFCbF6pDOJf/idRGVmMWOdKXqNM93RCnkti6ixfxdT8U9YbGfu+jzxHlv
7tEubTN9KtpwDV2kNFnrwl3+SrpzK4U9vtZPzVMZtjdNDYNBuboa6sPaE/pEF9sW
ks37BJqzTWXJqQYh9uPUqVGABweNL4XngksYikX4svXAo6tDD0WRvgk4Z2EZJOQF
l7E0yuwWHy+QE3UTnVymtwUH7xxZGlUf5QnWa6LhvXG2LlRBF+b5zU+xUvXZ+oSu
lgKG8on7AtbZAUcqrb2ryL9pI9/ML8HoFONqsIpy+rGaI3j+e1AiBPoikakSNk80
aU1Pdew/1Vg/SMR4M+ZepcZFvnlojtGdED4pyhUVON8bgM2hcvMeRSDDAWAqdLUn
QN4T+xPcyqrd7n1PWmhkB24VmF3ZMq+rNpV7fDdXCVtyeOoJlwiXNEXx0zczZCUe
aWlNhDCba6uKU3lhoAGsIhUrUMxuavMPQfxQAo56tELvwNIDdGoyGnDCnebiw4uK
mhliTKVo6ioBmSwgR+2pDp8Ebl5LzE6fzi1UOqVkiYDnCo0xIGOXFOWOG8hBCKXK
h7LFUNaKJiF1nabDBGnDonrCkbr+MJONy0kH8OcM9Q/lsDkhtFAdQD45LfFiGw/z
aK+P2vJW1yoG2wCQ0pR8gWjMjcYVNeCTkhsHOnZ5ELYlYYx8NR9liMhmHeXt1YC0
nHsR3BL4RXyyRd3HLiXzmoGrBSoPv4gxeeVJPatCZ0QOrZICEkDwLe1FyI5MyE6L
2EyayyUsQdG+twPBNhSR7doQJgqrisS7ecYbXVbSJN5JF6VpfS0tO0I3tsL5jMig
v37JNNx71RYRLSlvkZdalVge5DSAVtf/4gso29oIgXPRKgc8TfLUfoaV4czDUsde
8GdtMXtDiqvjoaoPF/7KLYZ2gGT0TQZn3ItU4L0AfSDTtjNQPg9pUdURqjsd1Ns4
iBuAGQPqKff6dMb3ra76WhEYYY+YicqgV0FsnNqe3VTAH7cerz7xbhp+kPUpB0bQ
Hio2XzkTTzSBMjynNBa9vP89+yg/7dWG+q6ltPXfre08r9ZubLF+5+ypjC5I5jy2
aijR96jXTzpWDZjWLhD2foHvo9xtYPC+OXYmuIeJjENRMfyGVbeIz2YnfJy2BIMq
uo8nLD304+iU3Sv1S4eZcNVErS4FOdvsQdQ/wlYRRQJ3UgJvidCtTTiSWJpnsMY0
qbpcSsBncW6hSrz2ol8UisZbUqK2GL6SoOY6LzV2VIcHJpYcLNwJzlNyqcof77tm
Syif+nAV/COqDu2q9naSxEOlketGbnYT1A/26XbEWS+U712bgurWACg2ZlurMk6X
d30/NsUodvLrHR8gt8M23yVzGSIhwgR8r8ciYwTWhqUxhIjbCjkLzdP5ew2D5XkW
Qoc0HkPcMwFtmjweOgEQOzBklrTJ8H0gH6nrp3v27UrE7glB+UHHqscnZMoeXaM/
pDXAAr9JaBAoXm5Bx1YebsuADkGhhW439Dr8YgiSDUTpD3p2WBbJx0hi2tIm/rHE
Gmt/AE+IGlC2yPUu+BR+YlBLLUbxrIHrxWycFgt0QcDSjDUyO9H4NKm9GC0MUmxF
C/BHIn/7HTDQNMi7vF2z5K5q8j3Z+ObzBVqaOmq1AlIOH8/CtmT1SoptuxnWeHlt
pM25e5ZiRCFKD8Kd1TL5acQctnnUqVl1o1wWbImWnKQQkUxJ+qGQ+I6BY5RtKbpF
uVhdvQV0VQfDy0D+fOC6FK9UR5lsJ3YibNYGsiuLMNf7BlJtaQwaHIh8MG1n9xlH
u8XWr2D5uY6A3JdIYgSathnT8h2CRe9xFzgDNJ+/Vx0Y4im/XgFlAFDNeM2ZNjXf
oH3kRt/xn+emUZJiK2IOdOuC7TocC1dwTsTPKSYqsU83DASJdrI3n8A0eVaZgRG9
/P2DKmFBerTlwH0ZVQr8KEgXSXrawNNQrn4lft990l/1ioIRbqYGI3yf8e5qDmek
yQ3jcH3fdlyP7OvTwI6aByQtSTpxGJBqGtejHkjTpSel/Mjd32vKzlcm5tkRTLSN
xFPcWZ6RfG5kojCDkeoibqnDPqSf3yTDCOV8Y0+0ySXcJTlox/CFtOGyO1TnzWw7
hXtXYFEPJVSW5y0W8iWc3Imwbb6cXdtT7mEee0VA4ridd5Ecvh0aoWMMBZVv2/hL
sw6DTqHjo+GEmN0c/agvX4WCV5QkNzA5KOCvMiUoDBVnHUjfJRzyUKuWwLk53bNP
2IeN9vEjIy3eqg6UBQIRtBGPQoZDkC6UD0lfs6o5SD1daMZGFoXmPD7OSxXbGjlJ
6OxugLU0uKoUCFw1YSP9rQvVpp7h79fnlYXvcRKD72uHZw1PTeTthbPciEaHcsPj
IPzGq9XeKQYtd166sBvC6Txqq+c2/zH5O7OlpfRSl8gYISuTXKjqJBWuzXMDia+8
Cx9ggeA2SGv8pT3Bbt/9YawcCZO6znJSYZNKUy1C5l8Nea1tPmn6qa2AEaHXVhNF
4toFFrhmqqE3lnID+6luukd7X8A7iaKR3TNp2JVTyfqJjphEnbCXuUncALG/XlG2
1zIRfkdszk0FSrqfAFPk5jgHn/EsukYZIKXO5DN49Q6JUroGJhsSpnhJqJnSMxA6
mB56x6LC90Ef2QWuR6iK9WloR+ITPlKBAX+aNF8Q5ieJz9jeH/fHasLe0m3iGkgL
zOTaM+xRa6IIqkkZokFP0bvNhKcHZ+8KZ0hxhE6tTO1KlkMINnXn0XH/l7rKQtlv
++FRo5NfdBDfovM0k8/mZce/kO16Zl//Vm1A43Qhk8QcG5XUZQlRM9Npsl2PGA6X
YfT05SOe6tQnQSnXHLEHs655AVfbeHrnMldIHLnHxq5JyWA2qez3z3DSEd4BTgc0
rQM/sgB8wA0W5gwwo0BUBH0u8OXeluO5kqgFEwICs/s6IWRagpsBCsSHpUfvL7k9
y57LKgbKt5JPMNrGgjRtv0nfgL6AonP7Zm6MSrsOX8I97W9eoeXqfD28EXN8p5IV
bn6bxT1UZy0RlQuA9fOAeF13nxDLeym3VrzeZS64wNvCey9LUjmGxvZ2vMtAnAbu
R+Bx/uFL9XOdrMGEjM8HyYSsbNZazC94OJ0YIgKFzb0jx7rVpDTLdJTrKGtNoVSQ
vh/u2TVDOnwd19owV9O6SGoWSA6n0IYeDPGqzI7pZ23ZALcdmkaN/TKyOooRoHJ7
8Mxu296x7X63MNDJjcGOa+J55XIgeVmDXfgDmXdVdmeeB0TY+9GCy+/JPK0BtJA1
sneZpjWdWXHjnNkFP6+y3aYP8zUmHlThx7ftwofRMup6cG7quW7f7S7hJK+6TVJ0
UBGo/9Q3a+PV6qUA7LDv+KR++DLMTgmq0nZsJWv/XHjkxQ5LEX2VooRPesNmk8s5
RIktZP82DDWPZm8WX9taBdL0tM86gmhHKAjTl9W7faPxwDVACXnwiyc6xAs5HpXD
bf7FJ5HisZ7t8szBvp6XT256zOJz4rVhcbQGPDJ89qmCynr4edlW9jHFBKo++8eq
JOK2hYLJzZp6VJw7J+qkF5Ej64v68DwNBxhIL14UEeC/3B+fkoWcjp8CVPKqXh7o
mXBlp1kqsTfdMnUlkQGNcShueamQY249MqOVNfWbKtLA3S5V1dQ9R2xsc/BXoQ0o
rAM6fBjQV/LqBGtTgtfinU9bDoLr6ltrxBLCX/jyoJi1uH7BKtuMV2hUJmjmALWk
bPObyuBj3DILHY0FICW+0WYwvUSA23Hbl5NB4BCqDgNgkl9iOF+r3Y8+LRKSk8og
GHuoJj7ca7CFQSuP6wrAJUzUpOSVGtK3dTzSuF97b8WoHB5pXpDp3mpu4NCi1rzm
A2Cix3ILcCb8pCm8eaizZxKXYUJl9wqkZFIvG/Y9e/pb0+YPqKY4XhrpoFA/AW3F
cGMofFcFm2QrrXFzOW108fRBsPK6jwgn3ycVB/Jh6XKVU9hECfXyUt0YPfHSJBb+
PFEwv/FGa6KVQMSL/q+870LxqwSbj8xuzwDT0TWBX4Tp85JFTU2VhZPBDVp231Kw
tAKxIByHvS+WAS72+aMoNg7CJjXGEz2Cc44EFkXD0AY89kaw1KD4/nAUOn5sPVOj
9slsK10Brbhw8RgzOuScJYGZbxs12+l9rEImspw7acOSoLz/2lrQwVxDv3Ban9BC
IR/T1J+pZjIWbe04yg44xannk/cEpdEPM398fde5njNQu0glarlIOUNu8bz8Yew6
skxTgrp/b1xu2bsUJIm7QZGDW0waWDfunEyGi/+y1Z+3Uf5S9jUaQRO/kV63YtDz
i3giB0A9l/3TTlPdWdJyr2OkdRqLnHJx02ZK30G+Onu1E2EYhsU6RN+NLCsl2Cbz
jSA+mDwTXRTAtr+9tG3kbRUXwuJwfF945nClPwBJe20plAhGBL+P1Bsh1DCdgEdw
Q9V2hxQ2D05mDNT/2vicTHmsiYa84u78dsv4nqLoZVJDk3zzKfwj6ak+ZbFZ/jfP
CWozOSUEjqVBtpKmjHN5hqHSrr0T4LOPJ5hmcfvzMP75Ytg3QGxYhuV2erYeVUhN
RMlEA2OGpYMX9m19zqDlQz6vMWfSbHBFjOvGGkOApRUJUp7NwSOq1Mj4c3+Y0h58
YH93z0tMuQeyu+wwI/yTAbwQfpGuURPz2j8E9UBQvsFX+2JuJaDx5hEW/C+m0Gz6
XK29KlEXVcVUFo0WFR/npgcbyvfGv5/PUG89paUCNj66gscwUA6c0vJCk74KewU5
Os4TTG+YKmStAr4Lm0DKVWlV6GmGKh+ljmA3Yv97E1wJ5DCVxcNIuUDRHHA7U0i9
zuEcQtXGJ5MJh657cbH4t5JQ98MnkOYSm0aCvwsVvaQnP48rWiFQC2mTiFTq+DIu
aGBNhLuz8m8XgUNuiIp/MLzcmA6x1lV1bKNJpyEubPbpS9k9EjsouV1qriazfAEL
d11u9sIbaBVUIHp7ForoV4zpeMISG1aDltC6BlkhN2vABsaqCf8w99NIrjEPx0lN
M9YF2wBMfZNuhpmEPX8M6G2AVc6U64lS7AVn5iv1h4p+etw3dbS1UZ5qeIfhr27Y
0Xpk3IusohDG6qfc135xNRR5xOUN/ikYDNGO/VKegreGfMvfBHvxFxbYhT1xCICp
+MpD1rSxnHWAmzNrBcWVDwkzf9fUPgbjWcY5Yk6vF8PMinMWJEKgQLU1AXjE1GtU
iRJZ7jvKxceRr6/E2m1Gf5nFt9rjmvOEIC9GnSlVfRj8gBzOkqd0/nZsBrtmoDLA
Oxge3T93WeSOSFtG5+mYpDXHA7WbB3JR3vydrlu88t6H45xXdGNpZ+PsfqHOvr/U
O0sw85pkRFgeiJuWOmWVW7iO8SngTxLCBQC3yVCDKMCDh0xhbVQT46JZVmHFwxEF
yi4ryv0Q1li6IRC0zcrGn7igSjmUMJxI/DFQ3bQ9eFNE4zQzJ4NB0OveBXFgUmPk
HcE564lgAVaOjQoequacS2axL99fUXVftdAjwRYL8XC9x6CKoXSfk3Q+VRN0GT8r
64lGDm/2A0mE/yldBRKo5Fch2lNvFtxEn898LccF+iTgM0t1Ww3unbqZuAc8vtXy
WP9ie3q8jQUbz06r1jxUTtZ6IrH5VxZrK1KB26SNHOlbpf5raCOr+s+wkuvyL/s6
6doWxZEHZwz+gesjxoMdYOIlFUQmm2z04P0ifx60cfehH4N+vl5f5WNH6iWHZTev
wv4GNuxgwdxxtG/nCaZMXFjor8JWSexir2PobUkOsyKYjrNNPTBS8i7mvNFXYRAc
Wo69UK9xdpbCY0aPUGNPIgsBJP6pAd0WGFgBmnUosARlfqvKNWPtuAvGI+1sjJIC
Kahve7yhwlrLJMia0R23mg1JV5p5ODTNe/LRS+RjheAn5r3qJQYQ4supw03HeBKD
b7pRLBS/smMG5UHLBJOO0QNKU4C/TbTSCaH87ShxAPoT12RwQyWXOj5cbKrmePjm
PAjGOMd59B4EyhXz9Tbl18LiNMtVdrg1/2LE0kSb/sn5wfagJqP1sBWimV3O4Wrc
sFJqF0wvauYao7ZfvmOflVR4pJRDdPw2QPnYgNxmKiB6QE57zaAZz84UUakfhTv9
U+EgLX++xsc9gWj9yH6JaF3yLqOWcLk8t+BHeUAr5vCeecV/0tmPdwRKjC8Ildrl
PRinbvlzNEc8x3zyNvojWPFP5HKh8qp/LOMpAR/82Aof6ZeO+mOZnPElYC/evl/Y
LGgeM7aybg+wXOcB+rSZD/kF3RWVBmbLikmr7Y5KrdwK1WwMi8VXPbOauXtk+Lhu
oQS0H9n4KjZj3E2O0IXlH2x6erhokTkBqwsghIPkmdoasFH7kYBjBLSDaVjqPmKI
MuaXKZivhKYpdlb6r0hGEzz0TCppUuGVmSjWFJJl9oBN8TcWqGQ4donRuBP0elWB
sg+YH6FRPw8iopuCW0QuNvU7cygcnjrzqIc2Gaw51htu+ieNbcpo2nb9BYqdt6iX
3NtCD42En0ci9v8eMg79ZIXC+wzTqaJgj1/k615Rj/+bMfD5GZqWYx+yy5VRw55/
No/6YRHM24ych0oMtCnmIYXAhc1rPbwviUr//4IcJD9NLFPNxpsv9UpKManDfK5/
+BD84emyDsPsvFL7JXbh/LxS6R6jUDZai0B1xIwXVxbg+0mET5F/LDYp/IsLF3hB
lXXi9ASii10A7W0wI5KdQIqiw1OfepwsDD2A+Tm56ef0dlo1p41MJEAuqb/mYpeE
REK9XOR/4bVbavZ2COCNtLhba3B3UsjL1G1nl2FkrwTjIWuEZzCrROegfqgIMeKW
WRcThWXYse3682ioPLeJDOshzGignHmWd2WZ13lIimrHF6+hFx0pinIQnjUa0ljC
1zhkitsGU+cuCbOP8BfefBy2S/gHY6r8W6ErGb6NmwD28kSia7vSwJ+RYhbC3Dgn
hXri+2uMDALD6qAd1cPRTvrPXgc3pVXkAazkiS6CYceXixe1iMQtsghO0EjsVS/+
4LDLwlj5YJzvF3DVYZi2oBW00QcXTdNzSC5ZBHyMlz2g0jMlQeiaGOKI3IyCpESy
9S6CQhMwj8osrtmiUGq3RvhBjdnqfezQLZNkLHLVEy84DVaVHRRhkfgWLGVai9Ky
FRtIslpyoE8XzDVUHdOvmAw+ZPwmx2OWJyVcZryPPZRN3FdXJdhn+vHVbf2p95e5
AsBKGoRD1KID0yPpbgmse1gB4nQbnkuuTsVELvVqncObc4qGLlOBUarEa71eT4QN
nW/1ssjduGtMwMFrWFyoP7UjNskZUNk2DK7FD6v+8qv3+SbOaMAdTkK0RrK/LbXj
5PuacepEapwzBFvBpU+GrVUq+jSQ8WRyY0988puzrS48MjjskpCbzdZq2DJI279m
Jwvc0XrymAqqETJWYUB9n0HlHF24QyrTNu1R08CzmMO5vw+zWztSgdZ7RlSMmbbE
/DStcM/BGFYAResisWQS/mUqElfT7HdoG8WcrtrWL0iAPA8a6xsN+rRcBsjsDnBU
8p/saq/hsZtKbjI5OSCvhLHXqb3HqgRLh+bKXkPfWka+E9b3GbUz90dgjDUV8dAE
Xq/quv3v+kY1k9gKqPenXoC+oKCHKt+ucPVEH0H7pz+YpQbJfFDDUi4MGQ7TfVNs
1O8toQANj3Sh7EHFT8lAWrMfXnBfmbe1h3OSNvM3s863/I2r3ipGDZRP/JVwHF13
fxTsAdo4xgDmWH+YhXmMbrDF3GKAT7nlpTSBUXh5IO5cO8aVJynntCD6nvXAAi+C
HQEgSFo/sKHDXitNnAm8OBckf/H/dYr7PjWOz211dVN9o3zLun4PWdEQMHdWjRW3
QnAS0pw/VRx/wMX6AfyiviUCnuPZ4UisHK72p8pLfxfXQZP1T1S1ZcuEa6cT+zrN
hsT8udC+52OsAZ/xaEE+nyhpc3NBktD4B6wzTC752J1CbygrNAgkHItqM531QzWK
O/KvReWemSM1oZvWxt417uFNejdH4sXG8A6293aUActYhPBxg+tRcJx34VK0beIP
bjDxNNTmOAP/arA7DCSiRkvGT6yZ+xNofDzeJN0Y7TcD6sFp2DiujDucxneehNyw
IZInZzAD58g29xCqBVAVeg1cV5TP6Ltm4rWLXGpC6qjNRXmYCi0Wfhj05uGSJECr
2kSPuXvGzQMTdN84cO7wpTLRHUegPcX4/bYZWJDrTe5t54kXUPLxNigSUSieK/3J
PTVGcz7sxNFn02BWjbms4Xoy69CiaBeg8A1BOGEICgb6SE+e6usv+nkaFACPntZ4
KKlBsqted3p3edV38Hcsjbz00uwhUCNkFJNEGEhrFuA9L468TayiOP9z3PtWuv1a
HXkUAc8n4fgSkrZ+4fsdZeSDh71wn0g+a5Rsljvw3b+ddFBxutTLq+vcAD2mizL1
vuCA1+TgpFyqRl9izdwz5n4iS1Qtbb2qNnEAu2vwgBj00T6GaAadz4oV8TRv3b7h
XHpp0tqauuZ4qWn9Ll/f92QGHETqqDhq9pTf+Q3imCdI3yMLMKzz+pOTT+d/kOer
8Up04nIImfo6OrpuQkQohpFMBmutCmoz8Nvw21VowydhyEwWNLdbpUOR8cZjjyFo
U2FIxJpS+VhIagqqvTi5Dh3G9LDP4seR0vP6tEjPiDFDNqmuCc3Gge3fUsqp17tL
juCtUpbJ5TyMTQr9d+Ns3gcKbDFQQ2eluFDXnllIgpw379XhwyDAQjvf3wk/Jjgr
v9gsgxQaW7m9C369nVIzYdGdfr9+7a5gRfJkAXngwD0vkRAkkh0EKFTahe4Z1jqv
W0WmMBVAkQmsExGCQxLZ3674lIuBIVOkfvcJRKNDdua4+ExpPzym0BoTcdRd2B4c
vTuHXDbLsU4wpGrDcv2Q/1M0IDcHRnbM66SmZrL8wggo9nOzkFzRS7/yJnn4oxpu
wfBgFFKZP3HqITswKqt3xAVQ87MllFA/if0CK+robRg6IPZmW3wpZGWad7EJzjo/
6HHao5M4N+orJVqBilxdWlYfD/9U5XBnwICPt9LVcvM9V2H71J1gzTdTj1hebZU6
jY9gKShUP1e+zMvheWefdw8tyBr8iMC0J10tHSwYSk0h8NY2hRcTOgE9XdJSGJeC
1RqtNPpk0iueb5XeQCuQQMpzR7mQfwiQ5RYbXJu6kIakv1P+JImfFcVCCv8TXJsy
upl36qTyJeUDugfccBiu5ov7fH1blSP8YC4cRSBHHxrrWRazhEK79ayB8anv+tAc
nLzmuwTRXXzXGyeFdC1Ak1MUYpYrExby4Nin4ymOVdkDVnAJJqEZFItJcNvaKGbK
TpOpwhdnCYBesc7UYFSOQBM6JC0Lhmeo9jXJnAgKjPK+t6bzn0Wm4alJ3OPwJ+9C
Ri/kpfFLqN9hCisgR8EydgknAezKz5kFftqAsTOxSiwDqeXkWJ+j2+s+lpIvScmA
TDi7tNNmVL0rDcgimnfNty0Dutff9DTRaOPwZUvlr5dLdGzKNaY+cKRE7mNjoBM1
MEKILy6iOhbz1WJXzZxHi+/kHZ62g8YfR+iCrJT3edoC9lHUihCTLSKSfnsTyK1p
XYJZZnIfyVnOCVp7pupXMPtsSdhE5QJAqDxqC0Anio2/1cxxibIWSVaongnhG2Cl
RYwSSNiKKtX5A+P3qFxX4nMg4oHgp1cKcIzLSjxo6XzbyBHFPuFbY+NeJq1NV7Dt
DCmz+6vfyxZQTwD1ChxqwVshuaClIZdfwtj/daLJqWf0N+8rvAgw5D6cOOENGxhy
X/rX/ImX4l4KiiCP0lidw2k2Fcutmbqtx7x6g/prLzdwAOnqiDu53moU10zuIvmz
CnW2tR9tvkLvVktTkhVRLWir3+wWyt7CO3xutu+AAlyr5WhBMEMNRXBUFMd8YWZj
7kAXg0IVbIZhd8Z7pQ23voZJvpY4IQ3wtW1mBTarJPNV2QD3LRyQBpWCmkIsJai2
ZlSgGMJ/8iBvqV0LXtd4sKng+U9YLOyRxWFPRsddoMhULyh7bFDhhva9SwtE7ovp
IQMf0ZKCsyxLA9zMgtOnjwLJICj7jIv8MRt+FtL1bKByNzGXPNAEt3GL9WqoMEyH
XdQguo3WQiLT/NmD2FI045Z8x+7d2bs2MDnHMh+oSP34M0Fvzacb0qyhWSsB9ZMK
0UazReNKNObWqQygthCPaziHmVEJEZ/GnTlBU54a9QaFNGFI3V2htyCCTom/FYOe
FS2r7FTaabY5q0HksZIYMTThLlx2KjKf5IbXo8N4BBUMLFekIlhKXGBsE2FkLlfw
9C8vwGfbcIJCmIrUVEjmGcS/+aolk1T/1MrjbJ8heX5dzX13hllr+K0HlCMmB5n8
FlpJ0claFd2AH/Jh1Cfh5DCZI2O3o2M05S5EwDqCkAfwtMyG8bzCaiQUiPMa9Gxd
e3FHBX96zFCC+CDBnDCU/VmmfBDHojIturED6JBzSkixPZxMChhBuC8nE070IzJy
qWRNxpyl1loSm198BO4f91XPddtytVz3VHSRO4bc4wAbQ8XrpnPE4Oh+PxWOvVJW
C/yCHVkJ1vRLe3EmMFr1jzw3yiIKB6TL2hHcPDIP7llsrGVMrJUa8GfNKX54GFrj
AWl7jRxHzpvcuhQf69xClBtbj04KMLk6oFKgfL2EB7tQQbsv2J8z7oIGmrnzypA0
9ohprMoNYL8k32Gy9wl+B0Mo68mMZbZJViWhGwEPnTpJzJj3R+ckd77wHRaII4v2
Sj2RqYT0Be49kX0sJuJSHX8EiFAHh7e8MnpnB4OsUmexI9v1JLw7kKLMG5yoSwJF
rLKzsAuseO5JC1iKFAWIA2DXcm5pr8pPFYdrlR5z3VZckWNY2UUFLml6wywpm9O5
9hqsbYZiCjr0u0Aq48pawaeKbZg3WeounbznFzra3uu4G81DHsYazekAZtWw4dHV
cRAOts2C4CcU0VRKhtBj5D2NOMoVrqrrG6Tpq/GEFcFRc1nEwG45nRzBbKCT7Ty1
rHokLfWL91AYT9I+a0a7UlKK+YcvKNBFSvDEwI45yiXov2ZFw9JUOjYVJKDBANWB
4yCFH/SWu2r6uXDGf0xM+fOmLA/8NeTYWfZCc4lCORSGmko9VRxbwAPk8y0j3Kbf
K/eEAuCbExLJ/yw+jX5tov/z8ajVzGEJ/MbgydBlDxKwMYHR7f61tWwXdxZNqQkL
NIIsPIlK7x9uS3vG5tUbD10M2mx4YDm7tWteNJWWeBk+qsUc6+YaYKRIgUuPc9lF
lTC64lNn/9/CNw3CZRTr/lmaE/H8xol/3oujX4smFTpHpIyRrPTGpfnpkAkonstc
oxmjWdtEEhb0j0bSBhGI9rVElhFRo1OGfHT+iMcNTsxrkj/QJNseGD7gU/1PCHSC
ADhpPnTdR/DRYeJEXQhAcqRyK7RDndO8dgZW73VHpg59LqAJ8+GBOR4UUBWrmntZ
DaQplBHRHEAkXAjEJ/1gX0R0LAcIId/CgMjSMQQlR/4+RITsY6YKDdabyArWKVrb
zP4fcLo+ijbpVI6LprwdHHxT/frW+Fv9pGohlKTlisTamoco2uYFMEKi28/IvelN
Tr5iUXSIZXa6WH+1aeW6s540rFxIHqNK4Qu8a19RP04qo9lkDI3jximknB7Gi072
1lZ6NBHirkDsJU3jpy463Widn4qNpYYXGkDDNOPMQl4a/KXQwr4Y7lKiPvXrGTN6
MxfRAoFRRYYmrDCsDWijPE0lCE75W/YGVvKrbjM32+5NJc65kCUQmQsMg0IrmWxY
Hq78pGJujsC1AXx3xaja9mtcTkRiBnHNVPHC0X4pLX7jF8mC54vdYExP93uwgjUj
yDKFu8OoaZBv5O4J5dFvskDIRiZNWUnhbGkFiZc3j6r9zvkfMywHwQd8C0V6YOJC
+7reZvh5PUG272CKMt3JZQz1dRZLEqpGknYeidMBuhdY4/j9iHcdbgP9LrO2yjEk
AoUMyXHILIJbB2ZTlAZNQZvToL8pcde7n/idMFZHpbx/jeXUmDKjffbxmnDID0Kv
9nJKLWjkBbXB05bdMBs6jbVpD95nP0/tV5tzRc4wnZ/WemIpeubbPHzgM2n6EzxP
Negm8wY9P4gY5iDwiQwdU2PixuUnIkEsBayhHL4Gokj+d7ViSRVp4xfIqeegLEVM
lJfCh2Qx/6RWg8MY2tWgJmMlb6Oe2hdoYZ+MUu8+liatVbqMFbtqICNDBNb+z/n+
QJWaiRQscoEGlDlOXMGBFi+hpEnL8YTmrDd0KHo/J5A/0oVabl2aMapJv7NX0vaD
QOLV85voUo4wXYGtSQIfU/vLDhPzzlYtg5spgRC/wbyFESdAi0a+jzFWeUNnp0vL
P/RehPlzgCUZ1IoGW/vsB4zxAlhwC+qVE2dT4grerT6NzgUcZtWUA5jcHFjCKGo1
BeYh7IS0QuRSRmYhIUMYExILJadwSXJ3qcgqG6wQU9O4j9i4tj6NnFvqaQWY+slY
2IiVCz1WqFzn4WSGQU8NbktuaggoM3k8gZZYZtTJjQaHSZnA8VD8E2Ql8ShV295z
uHOT3DohPmGo9+vsWhqAlrqV7XXRFZEVzyc46fGq8E3E+E01/GbQPqadvl+CkhC3
T04cehjMNooYgPm1QrGP2kaLYakirYdVq9Y6cgH74zTqHAUX+i/UFsmgNb3+iAG2
8aCpXtjx3+qCkcCCp+JiWaQMYJy6bwA42Moj3Hq405UnyUH7cfmLX1aSRwS4YC8A
FgpT/G5IZYVCd0IjhhdQIlnLtG5Uy0yQcr0xJ5FohAN+Hpt0uaLDKVeke52mViwZ
5ekeqqpgyTAK66wRImHsSVEWFEUI5p8/Lhg2NdjCAnm79ah8liZy+6qs/8Huyne4
5u/ZJc6LjE7MxFXaRElGzVZPQmAseHSW197rBPrq0FLgmedZ9KF0mZQXn4AeyvMj
PYfetYtmgsuMMtoUOWae0REFAiOeiTzT7Alcbed6imfdMZg6LaCez2GPu0fVHLh2
EiuvYN0DyRhodIXJ3zlEWrNAexPs+bDmC9IF8rJuS/cc23upPBRPeqTso8FMcHcU
f1drdWRIWQVoAhV5YBUQ6Um5aZnoyJ6fsZ/yz9UmT/yPgtmyu4VQ3U8yzIm0Jo3m
gnADRm1IlguqS4R/HiuvXH1PVW8wXYbE++t02zq2s76lJi6G9vR44MuDx+PjJqwF
xXBzhKnCvjP6E6rgDr8FRZkRE8hcTRMY2TtHcMTVzUowAduEoNLY7JlTZ2ktu8AC
mVbi1I5dmIC2bW1JWGVoGVtRWBXM8vVCPrHX7BaNaNlTL6vk9X4SuOSiH1uMhjsY
eVa+yqykHhxJAH0dQiCh3YnL6inCiMqx55bKWISuu6TmASB/+ubaBN+mzqUiNucU
kOti0eOnGdX0/Z28ChDnRNxofXs5brkxe/J2Bj5NjqvuBh62l/jauNJ2KNzYcBiO
GYRRRE9AtaH8LE423ygAUt7wJwtGSco4RXpWAHvYSKecdFAohS98IoY1HjaMYGVj
N5rqsx6/BKM/vIit4NyfQZQZ8XIM9et5iolLV4IGl/TkbIGXij8nPY6IjaS340Pg
hsGBnY1rhMLxLeqikQhxmh3UZIX29vsWN5QNlxNt4DHAo9ROd96BABiPs/UwhDWW
Z1pbrRZG6Rv0CEIWn0cIEvX6Z+UcJgj2tmzYif3YbuG/Cj/Wm2CenXZf9i9ewQDa
FKcmbtr1N1ujYfu1h86gPc1kEgutKli8Ryu/uoIQtny8zyfvuTOwKQQOI04ybs00
klv+fqPft4NEhNZV++7RQ1prKZ8noDXFamdYyMWPk6RlbXFCQKzN5nGoBibdvyOf
o+c+2anYG5d02VAI4k2XQjrY1LzuibFx/2zj2LiR6q9h2ZUPWbzFoIqJIdCnAzhq
MBrXh3TPcUOSrZyqkjJa8WE+VpVWnpGGeOZfe4gPCeFy/Vqmp5ILImbXWB5ziL+5
Pc5u2wroESrVlwz6pBKQDHy3F1yXrgw7iZ6nBHIJbzMqRiXWOgxwm4NWeSGc3lVP
tSTffyqo8daqVJG/89hXAzlXY+UK/gPoT2B1YhiCOqfx1u5tsk/9dOCTL/4aeBf+
41UKDhoOGMTI3xlmXC7NrKYAcu8lAW7NGz5xDuF6ZnG50J2fZnulcQ2SA/GWoH+l
q1Xlg8dpToDxePV04ZEHqYYNW26VPmRz6FChp89zGUzrZY/8bYo0jA4gRlubb6Ve
zeMM497ZQcC9BgRuHEmcf8ZSKCfK/10p2FPoOnrKHrC9tbPCnu8qv3JS8/Inh5aI
U2WcSZb+33K74Cf95DEHD0URzGnxKXgVyUvFZ/14HAdmGVSr7KURvPJ13G7RN1sa
hQB9/TR869E1pUVe4Ru1eGDrJnepclkOGsD/j2gm4yh4bIeYA9cmbEtoeP3r6Myl
+2DZoPXto35mpcr4NPPxUi9QK/DIIyCKwbzxsM/MI7mDeurgPZLBVz3zYjXx6cW3
zwFZ8HvYrwHizh6u5M8+fjAJGmx8xp7B3gWhyxNfYe3Qwg0qgbPfLd0rOIfE+Ts1
2ceXX/SQT+HD6Fht3yKmSaaMVfjU3qk6Jsq0++31HfceLE+4TeiXLHZ/X5NlaMo6
9XOlmObOgIN5rvLi8cEAlfQ0L9JrwqMDsgI/baEzcRkfvlZkxaBWum0uIWd55xmF
CP9HUqYsQ6lskacIeL5RmmIqOgZwNMxufv811ZxId2KzahhqS7GSzd7sS1rNQ+oT
FQM5iXxwxMPOgv29rBu4WcYcRbORRyXP76usez6Qx1UmOg4kxNIkZayVGwEFooWP
cO1UnrHR3Ds2hL84q4PTAnlKQGjc3119EDjGUtl9Wfgf5czyA3uFygRPZGyf7Hr0
lip4CGvElUqUlKxYG2yHyHxE7mBX1y2uSdNKAy8/OYNT1sKAdMpYjhvf79kceyRo
+T8NFeVK4SBc916Jgy62yA7Bab2COvXVbwEva0q4Nt44/8X56jOb0r+aYL19fN2Q
w2n8MKnL+hcxhfUENGjEYLwGbCDOtpNAmuJTrp/7925UsGAOCzz9DwKqVqmQC0nl
HuCSmGIhcCDSyCHqV5Oq9Z7ujX8n1TklLUyQmqQPqNH1WJTndyLupdQO5XUuRXn0
wy9EytHu5lTBTUQEPkFpJdB3yilKxy4KlxkISxTTwjcH9augv3HEkEAYX8b0hLGQ
lA8FHacc+hr6yqAMlt7Z4NyQlsUSRaQXA91SxFlO7WY/Sz9MmiHUGobjLkai6iPA
ueYgWJiLdWn5xLg0OGF4nGhxFmGwu7x0V6myB1nY0Dw2Q42kUZ5HkmVGcYtGcwJE
yNI4nLFP1h4YFxnXmr0nSrQBf0Y1AoF1JCo1PgrEtyGS5yvRsFqIYYF+Clsrypgb
eEbB7UafaWi+dzilff7ES7HAytdNC8QvFDPrCyC7XeS8o1waaXEOHeNzTb3osMA0
CxX9WrLLvSmej/ZGvjXSxKtXC1iGMjeNoaO8E/huiBSVeUTQnQrzLwEqVbOygY3B
AJYQH+Mf+33WFmfoZVC+g4hNm7QVrd8hmI7AF8OaSOzAlZJ65OmmjzWoPvR0XEs9
IfCBVhe5+zY1ZAvvTyrbSn7HglTFE32fk63jG2S0XD54EKMSG3fz1NQY5ckUFcWZ
nOOn2ROSM5rxES83iwMa7qHo3A06vuH4TbFIt7DJcuOunvJVqmr12pL0ROj3hz5C
Ra9Ggn+qOwt9YZFSr+ENn6PNpnukle21hWj1ar35sIJKfq8FNaaGfLSrooYfZCGa
6uuYTjaf/vsGZqiJ9W86PDR15OYYykmSL+F4Cqb/IJfjYD+wshv4SZt2tw/adlqu
NFp2+I/cEjriYmPe/jk32eL2knqHhwRI4QyT3UYqpbtNXYsHKZ5Z/i9JzlRbuHYk
18iccoiObFD5NPZmyV6yIfnkBYyxN0lZ6qFSJAbVegS9M7LYU8Ge6FgXZ5Hcl7Pi
HnMp61TVSlMNKtlglUN8wIjAc+nbvnDVQLIzicG5rFaEB4TVOK/i0Gd3+mUXG2w9
TprYldefh2svxzVjifNpee7jC4CVLKmHg2AHLm3h/iBYHp8Q8SEWPBipvZD0vEVk
tNMoaUvKAUtR0auffgpfx6oPVATYeM5N6+CPtSK8AXJQ3DM5ErxtZ4KJVdshz2pF
FW/Wcm6YCMdTEBG5O4j6Fc4le3ukk/RQ8Us4d6ZBIdDmfVsa4nmrdlG1nm+GJ2p+
isw9aecf/4xESnyIRzYjKExFOUBBntiqojaetoYk5gTibnXWuoSh3DPx8EioeCjC
+mIhchL6qjPIuirm5gabfwnusYfo3ni96Rv5jIXfAPQljxZDA12znhFjmAnIL1du
8j50Nlm39F6Rt6yH9dO/wsq0yUapQg3H/BDi27IZLUikv4VKMtIEnkUzRV8qXLnb
GpAyxKI3EoSIgat+hzeMd2+Fy91eg8476lz/1doilt8ukpctnNd6Ax7jdtFdcT05
Hog4V5Rf6GQrjo0q8PCShloLpTURV3H/xDlZTTkxbHlUmh/8N7rIC6wsCNpWnChT
XRuvZgBjro4rYxmFHHFK64MOBi8HityV4+e6Al+bD9B55BoTvFBG+aJOEf7hd8Gi
/fiTJlp4mCXveHkYquK8crC18MR5DNk/5j5iB0I5vtbg05B0mzMAEw7D/okBBE3+
odzydhip3nn+XZbKatnFujGe13tu2ggZZC3YCWoFxEv2nnI8U9kWiB6TLeWTzKUY
4k+b1kO0a4GUS2FP9T29MzFJeCSVXSGYtwsK4stfX5wi027C0+6JoX9xd5YlDxip
OVk0hZbISE+fRgS04Ay/XVASnG8rwO2WvtdAfndLg0WU0sYYd6HumZClMdDGmXz6
Ib5MOdSHUNZqF00RVVqvRnx/ApHwQqd0nuLJXKXc2JnW+hD9DubDCnufH7iw2Wxi
IwR6YK8LVp1BsD/K0u5PPu0LYQf4rHdfjn8+ZEOnCPZbaWIpd78WeyWcZ+ehZ3dW
gFNjTrjzju0KzslFIsuf4DtkUjfFFSLiJIcIOKNZufcrwfn8vMJTtADGC0U7cLAK
UKdODhUJZklDb2SnAAmF0PDcF/35Wc0m8tVCmBPH65MgN+FDqOxp4NAZ+9JgX9Ch
ieCaWZyhu4W57+x5yGukZDaiGdGlpTItbr7hABFj9cqNKbDw9dzXNgcjnlAaKhMF
EdeYBt3aFdM7cluxJ58rDPIpluvJ9yDGmzH0zKD6QPVp/97lPUaZ0SK9qMWQoE0d
4s1y+jRvLz9bNowL5/Z8Av1XHAU4tOlcseUfqkJ/OMtGCAvfF3/8OtMQNafEqFUB
btGocgsnOhjFWVaIGb1gOpjHcLYpK07dI70v0P5S/QXRSJ3sYRpNMnoA8kbnq5tL
kuCTZWBplyLBdf8k/Nvc6SI1q4I5qdYfnXtlzMK+wFB7jnR74PHk0zeGzFnod+sM
B8D7TjmR/3a7BL0TU/OLL654qcYZDYrbClGuWyEbFdoIS2tRWgCmWyGsSQwcJei+
yPSOvQ+mwNO+30k51aTcFI2TaYmABmrkPMAcwBWTl12uk3EaLFqWJyy1thxIMXSA
edjTiodIXfDuH7BEK8W14ZPoMLDy9T0qfuSW6B80Neg4hv6oEy2VMDB6PE9Xij6H
kwFcswtK5bmaRq/tHKTlLj+wNzalsutZ6YxVBoxkTxZ/HrXzNf/T1gfWaWmsocWu
1PUS2rfs7H5M+Lyt0xelzwJiEO3J893CrjL7I19SMZ4+B3WdDz7prnbz+kSs0idb
7wLSKu/j0w0U9CIY9rm++18EnbBEvbN19wBwTcwRrMdiAYbt5ccBFCKEW3UX21bz
RnrRcIgQqIIW8Hb0dT3d26iijHvbP2ucQA3Iz5L2FwovHV/LyKfYB1iKKRCsmqBR
xWJYuy/9yQCv0B6dSUOQ0QYUhPgJ1Om1WqWnIiKupPzWNXKAo+8Ah8zwdpQ46Ps7
ehkSihKNNuH+qN5BhxKjJafvq+zSCSisWOg3903HQH3r24Xtz0tOvQ6z8Ek22EDu
ISnfDMaRWED5/zCRQwSrvxCB/LllRYP+ldKOhqLWqpfDdyyuTsPo/DCljIKXvBWl
y8/WW9cjPuJlqBCTXqarbIO1siYVOtbGsiGS8KGbQbbeRp/uC5rAR/yaBm9Y648J
98jqIGOzehE4v9F/Rxvc74lIJQZq+lmQP77MM3z0+cWDwxtClJkqcWa75X3unaC/
N/AgAOBUHzJPeiPXEv7vxNfDkPOtJjBfNaa4NCt3KYdtIqGMNo0UPE+1N5UrvYU2
sOpTzGBPrs3QQGZ9i/S/w7+2Q8A6PIvIrpRb9f4OOIPjjVvxFAVBEvbwX0zcypbX
WiCsrm8Pn54HtFWSRNXi8Fp/CtB2u2/Qg+ZdGrxTvjOcQHsjfIX5uLPlWws5irhu
4sDOeKbrIC7fn8lDS3EX6iNDvfZuERK6AG+PyBR8Ct0Qn3DfMRmPaHusMdo4xTOi
AmqbWrS0k2lkDXg29RDz4a6jC0lCRItZBP60wyDfF7EvogLHuu0+Ynl15UQvz4Wz
k9hI8CNtW46jnuwowYp9TySpBt77rrrhXmobOm2vuxGscJVso35cHJ5kCcLAtCcR
BGOm5Av8d+IvH0h3y/tVAT6D3R9z6HFfzEjxVS5HJ373RsniLiYdciz3es5cgvmT
Nst00eP8aKliSJlOmiItu//dQsClZm9ApR9/keuSeTvJaSfOZGMJXZgKZfEpBxjk
R9ip3rCoUFCDsWQcc7HYfdzxbwI1phigbilj2tRN5wJHsG7K2a5aILkz77S7QaoC
mwi/FPOq85nl2nSc4AndFjp5NR912mfu19JO1+BTh/f7e7NfqMn/4ofKOjRAVawk
pOnB2XDi3ajfB9U9dCOEUPB8p0zT9x4fPuDxZHmmFZinNIOLac+QCs/WJy2VTiAH
ufzx2cxlczhnQcNDTvIwZ4Yptmd+n6EYQDU5DxvQ7sf6pk6nKwMzkoLb16havZiJ
MHUMBnuVa11sOwpmOGpNS6ljKUkiLlfkroHvd+OZS6WZRHGo83PCQedp/wBhDyf0
533OnOcgXybnjfclaM4J3KyrLWPsO5cgatROR29/ZZT4FRdfJIOOtlTch0JoWwTC
b+C35TAkU79bfR2RQTqL6dwtbKBSbjyy5XzfOeK8qwj1S4sQf+3zAyMZtCZOoqbY
OwdwAVlrPBaSRZQbtuZjOQSSippwmQ+9q94gCAfiJQdgW+LIvCvhAHZnld1TNMhg
clNRQySVCNebud1vJLgKz9T7ebvgO2agw07fgGRL5Ol8ZYZUIHhVVFtgqZlVo7ke
kTxWo0urfIAMYRKqhgceyO6virRSE3NYGCDk1jDBEzoVdI+zEBvcZuXMAztudjyK
XKo7C4aTW5+hIyyM0e8UfWQ4m6wWuPFq3H4o7ffdxMrYDKLNaXgjHfAlkTd2Ih37
iWDavTgjrievd555mAQ0hQe0DlA1Z+47//RIWiiKhyNJ2ND5iRJj17UJZYRVTBjY
cdiongYj6GOm+bu58vzbIR0dNry9mcpTDdBxpKt6LGQBONrIW25/NWfw4e8QF2xG
soNS+oT4k06uF3Huo/gJNHaAuJoCSs9BNkR1X2vy9e2jvhDB0vwssxlrcD9gYVin
JKdf4b3tTvIr2Sa4v1xsUptkOW5WvHMgHRNFVT7ZeAMX+34R/NpvguYBCrd7moit
ModsBcGBZMMX4yoAap1ZN/VavZ4P5pyVABEsFtwtYsczkESyDaUUjs0gklcGxtMB
s1jw+SyRMZaLBwxwk6DUTQg4Mc1FH6YctoGxz07QWtSaT64zo34IIwKh9ALpRZVe
tCy0pN4DYRydDrOvCQHGRHF7otihbp5FH0fOBcpM8AJtBAhnJwq0fpRmeolJTXdW
YOSFZaR9Wmm3LFZd1h5C0rToJRqVePN335IpLcbZgpatVQxRwDOt62IOJGOGlXvS
AXpQ+TWcME6Lj6usDSVINxZ30zY9BE+1hNgSS9C80hKjJMmqFNzsWBnKPEO6/noW
TIx5ZEv2WiJkWAe6ZdBgFbErWjpws0jtw2O30XgqL/JJNExBHr1OnXyuzjKMli07
dbsLsSo1tsoR9jEJw+tj02kQxyNzGk7FHhW7LUt/ACGqfQiF48iyXXqAJyIE5XNC
clmYboTDbNciHw1M7K21QoieGtQtTutoa+rHQNEmyagNCHd8xMDEKgrY1kMdpodw
eTpZRh5d/Z+FG1oAZn0Dd3QUialwKUOn+6CHbQHN1f70KJalrArjXnK8zPV3qVMx
PVxpCmsCnUAXZ21F5ranyUnhECU2n0dSeRWz56e0YrlfW1F4LjLmU2UbPkEuvI2O
vUIMc/LSqCk+o+jIK5s4fUskQQMsx6MVb1vjdYwlt1Kyg9Qj+rambPKCSVByrSYR
alHqBb73TyK3Wsg58FKTueHOQjxBbdxJf6LhjEyCZn9wkjmMwr/Y8kLFmwgnhgOl
BusbFttVKYoHVRCt9pXW30VAhf/E5Ff/cC7qc/7Sn+Kzsunh2euPUHGYsyevrNxt
iuiLm7lVifEgmFbBhaXKgg97l+SebVXgE6imlTQmdlfeQ0WofcZ5FCgYI6ycEOJu
LsDOhqaT9QwqqoVLvgdpA4ZltSA/PVAZ72gls4bVhv+1PypQr8KVtK6N/zd3kbrr
tecfCpvQDnHqQqfQhwyWoMcO+LgS9ZD0dOUJ04UueuQx+gGpn6HSkJ6Dy7PZa9MN
0r2wGTwdvdQRwul+VKrpsz4AUJXsiQevZD24+5Fc9c33RE8i6rBrA58upbVNBXv5
YMAiAYIhyoMIPFsAN31C1e+IkuFmXOoBKYRgFAPP/6JYJuOgyMa5LR80xyYay7r2
Gz+YWtYulyMHpuALUUmanbDjEm7cxdgoseF/8tz8x5zDG4EuHsPZYA1q7Zpj5/BS
1qahdB+lwkLPtJZf2zLWGKwdl4sdFVq1ZuRW4BbqOo71h8cT8k9vrlBmQSeVMWPk
Dq6Teky5+/1wftx/ex1BR6EHiwYnaI3bqe93AsapQLTqiyJ/kHrHdXLqUa2f2Y6w
MFkFrFxE3egLaJ7xxtwveMWyt2RPB1KXYJUrQ2mvxIHyPukekm3qrICRKfwJFRBR
4903taB+XrCMjErp8tQR/jDMBDAAd5VHUTHY9f9/j4v9IOiHr4I9/mxxgYzZ2sr1
G7+8tHhJ9qhjBfOugYaEbR87CiW0hJ8B2GQRrI8+95FS1nSbm2NulaoMkEiWPwDX
0yhYYqUJoERiJGzaDTAAfmJdg9AMNHCx6Anaxdbx44bG+N4LKH67Hiz4v/WtnRWW
IPzcuP0GX9koSrfzEvrtj4SqNAXbNp4bVZ25mm9brFcuF/lT8Va/ZHMLnkdljPUG
1am3LTQIjtmHKXKMnupXHb565CP8N6mrn4X1/Uw4BKkB5W+YnEpwg9FU5OuNHQnI
hfq3sSBi6FyiyyAPvJDHovAiXmKmkg3cR2elzH/V/sT1jwNg14bpUg701ukYElMm
IqoAD4oTJ8bg16gfmYltOE2rrJKENRuOVLi1xDfzUM6hOuRfJ2RBAz5UMtBvZxOe
AGoRujPtcQJabn759ml1PxveXX0bOMGMvuz1ry3POvMLjELKjuf4DTsbT0Aguvi+
TCU6hfUU2J1h9TebDKksicjmHg7zgeuQhyYj0zsm8KHN0m2W0dcyziLzAS8pvJKe
xk9/bYGEllinlOTTpPEiWtJaoFMGgr3S+wRJ0sLUGUq806s8S4SxJgiyzIMrON2d
UKDjaJ7/vAe1vAyMtME+cvYqGScf4mFDgDpVD/ruGvQNQLn2zBPiNlBHInYhAvjE
t3I8eYptrMR95d/0JTWyVqHy2j7R6kAbddKyXaQN+VgpHKxr8sM+14H8yOBSw3L/
So+uNDnIZH64uXHQnCwJHuY0D0uHx0kOBHIoID7CtTAzr0GBsh9Kdlff9n0I7QZv
ohPfwimLZCo2uEHy6yvScw+gRLxSFgPptLyctF6tVECrrs6rpBejoMykkD+cqLZ9
kgb9ufTA6uE8qQwNKvZ4pZPMV3Q1g9nUvbjQr5x0qat0E9NiuuQ8jEDPHEt8xM03
q+0TRM74U0qSmBqqUYW7V7Yayi7RV6FyqhaYyxfpcBkW9dzJR5Ssb8JClrBcxw8G
HI4G9vfdu4VEDpmgVdOxlmeYo8D5hgrRd5Ykk676QcwTtnZDsP0tQv8ZnOjVzmBW
6T1Yt5rSyyAko+yPDFilJB/O+lj0Yw6C71tXB8pq4q6q5Y9KA5DxVGG0qpnCh6/O
KnrkTkLdDo5WLjVYlNRKL0v3VHKevMPHVXpmvT1xcozduM+MW/4NvSWlNvLDm9tL
029zmZzs051ts8AfIdcMC3ICHXO6XZjuxOKX/52ccNNt44nkOa28wJ5SL91S2HgY
rWvaCtLvOOBEnTqA8IN74V82kyhEO5G5T1Ev0ptUD7212ssbsmguy0a694kCrukK
YZKjabX2CbKoPS/P0OPQ7DgruqA/g+heGKuNL1bY+GjA4EREFO5q3E66s4YAfzxu
UjaQT6AWWgFcRz3RibBPDFK68oGswo8a3JxKYnD1M+ykvkP8E6MeMf4IXucASsLm
8toqqATCGrgpXTG+M9vzQ1GKIRbCaAXgAFx/EQ3af4ql0eNzq6IqQtn8jzMdnaTe
+fIRSQZ/X2MVlVRC0krpEFT5/CHMIzOobCL1I//BZYzzmpnx4A1ixfzRpVEE0+To
QR+MGCPGdNUoCDTbXdvDNzI7OdIX9XveGzo21GrvZ7qJzhE0RBK+eCZG3nFcPEGm
zW7o/71d61/m9oQGl2iKYR2KPW/v9Y1CQ85bAHm0e+yL+mw7wqNVGqtCqDIlKNhV
Y8ZPbB1d6U+APs4M1KNkbmnkkDSu1dh2osC8VusbPL8FMuKpwHirbNLCMctW5PqH
afVO3FOC+OVf7rGuaEdLLTZX8vVkNuTXa15KJGbVAK2kUdWvFOu/c5O2o4k+Str5
azreeL0U04Ar8MS5aQIhDIwdHH485JRdyq806PO0S148nWJtIMNVOCRajy3SZoty
GO0VN3d7i31HRyfKgRAaFw7qeQ/YyyMJcWgARnPf8STHcNPR8c1wv5lwAbtY5y14
L0wZbeGeLpoxGSArcNWLhGni9nLZeZrBe8dL/WS55eJAtWPW8Q2IOeC+SwQSXWoW
T7BGXz4wmG1/lggG3bSjnRWoxxWArFiC4bu8aDmm+SsCuxwrpsewMAYrVKCHpHEy
CLPGMjdfqpLST6/q4FaIIjsUHsmBcsFVgvDqA7xEWVzS/EHR9a47cjLHM8M2x1Dd
LY8j/IstGKB6fMc/1//9yf08ZQ4C9nubRFSTc8saCKHgD+Cu5+1PCrwSDfu5o4dq
xrjg92RmwcQTOBpxToSgl3y4KbS4UOvT4fW2UTcvhG0Ry3Li9mlqav9tCBGzmne1
GXmjsK0cmcHIAXeuaS8FDNlzC0rMok5A/+2gkhdLx7fMtlTlkEAif1/m8FxJ76my
G38g2eZcCGrjlG3lEbAXfHfwhi0ABbFwrudiDqD/YioMjZ9sLm3K85HQ6jOPUjzH
4REl3zCfU00aCzvoKiySomCE40uU7d0jlU2NI+FT41WXVGxQY4hJqQnX8I8t9Ij1
+/Sxg4JQfjkox9cKOlH9f1j2TXvjMUdg5KOa0/ODCZWbCMW2ZC0tavGoi/oS5+k7
ZYHElVShskMe6AJqXEAwx08d0E+zY0g4WHss9MBdnU4u6vKw0wTww0Fu962fM2SI
bNZQvsTl6ap7VKm/f+yNMEBa5YMtAh4BbUho8CIpLUtgIGm/WXcKEZv/ubDRFzkD
lcG92LUFXXlFxCOwJuRGBi+kwkxw/PkIJ1YSdAqRS57wBv3PWavLbJyxB/xrO0S8
UtysO1IDlwWxNQZPhnk4MNj3AiJ3sTSTkk8UIuWBYgjps+/4BaW+ikSIq28oH5Ps
l3Ul2WLLDNmkfK18VVsBF+8B44jrKuateE0jI4LfTWkpv0q56Hit2M+IZ6UPGxrN
K85vpVwSMUizkm+2xlwblKW8q+9M7V1qHu3ZF4brv11WkzD7q7tmwb3gn6ypls8k
lIaBGsIwS8I06OLThpm1Ukwb0zx33qTXdMSPOk5Q2ZEYZzXvtk1wpTq9H+6NnzA3
0trB+zSjkvZlsnmh9hr5XsSdsP66HGlvyAG5mhqKYpu/tv9iNcJy77E++ZXPiwKK
AWmvR0dZfFqkjHs1ODKnUSNGwPLkdK+rKGYB2lhqOBCqXor2xLVSz146qOkxSxIW
XIrASkw6pUn4QtAgvPv8MoyEdjGOYsrMso3I65MzUEyRYtMrmqgIoaMRgOWPFOy1
9fGp7zdc3v6cOrv1/2SxsaYPLK5SdGWhHXC+cgNy/3C4ZASLSLIiKeyp8CgqA/QT
o5AzRh9AV3fP2HkVvzDWMG2Y4rC8n5JA1A1dHG2xA+aABFqXOZhq7mcMTHpp9CNb
s34dpRnAq4AxJEWqpKzt0kyS61gLsYOStatReI+akI0BDV8AnJpTuuxvJX3ML2KP
9Laoo90cCPtUOotWCdO9DeuWvXMV9ZK69HbVixNqTV43R3Lsz7v/5Ee/2FEz/SQE
xJevlXLrCMFdzKyuilEbKgh1JQ3u2LNKjOFTWyvKA0E1709YjOIQ7bFoBDN6HKt+
MLlID4wCcD4RqrtHgApcmdFEizcm2pN7Z5BAOUNDxobo1CB+agLxMvEj6LWbfFeg
5F7OBv9ZIBIJ+q/J/to4SK5amqb28S9/NCACefkMSVXQE6FCFUYl550nKL+7SmSg
iVsTMf0T77UhpBre6XvfXhW4DrpYQeqQQGB3zi37fNkX3Fia5UI9cXXa9QYpH36H
mJiO/73lE0UvxSxQPA2b9gv+e+u7OwZYQwZWHf1KyzuR28LPU88d9DxjlMcSFsI6
Nn7+vkD7obwCLWiYFuoI7PJ/T8a817WhtT7hhEVLGzB7613YOF7U88s7gfjlFXg8
TPtHAJjAAV3+D9BxlJV3IOERDMxZHwzxXBzLRr/M/J3ZyxsvATNBfH1Y7jCaGUQY
sHTSAh70jopPWuxl1di3+P2PY5NUqqaVY5TXax7UmeCR1VD20pFSPygjEWzKLYU8
pMMj4yL3n3xpvj9txn1rFBSAEkRKVttaUHzUt38zD5AcGZOeGkm/7C8AAbCGnClp
Ms4DgrHhGr0X1vok4pXvSf2GU7ElkoULGPgxdHUtH+Zebz0fjf1nqDeVsFm3XsLc
G1gY9mxSJeLCbwmn9rfD58v2DYRKaIG9oe7DPRRjbDaAzaTbp89nouJEsMdZgOpD
FVPC0pzV1PcImFK5gFrLdHSfgIlwWlSrueffV70VOrJqqu61quymsUIepB37bYPa
RN9UeVJor18SMDxID1SoMFAC/iys0q+1Yk6q8kVJhIbOVwItOM8LJTXxerlqKt6w
hPcXhY+WvJNyDxJ9ptcXid0GluKhbgTmDgQU2eBCmq+Bxa+KmzzjOSnO6szwl1zU
nGmYRu/DqMth2zXsInTMk5bByl3XxF8DcJBgh+Osp1ZbSuxUN0TyGv6jl8TRVC0b
AOenWqMrSsDhOVF5ofFH5a9QpW9rPQJQ/kIK0akeCCDkRrSvQO0hUhcUsXo7OJeL
7E75bQ4CSHjpYCxruH7kwMPY3R/N+Ji6UyNauijDfsxvydRLgllHgEe7DO8AMrdd
edqvKtMgfDRnculYSfFe6TYuG8D2XQIP6/uqfJyCtSPEZFPrsKSVYGo2mokLW9bu
giV53v6y9nncB/7Pvzym0bie9lP4s+iCxAMno5Z54XmeM2TQH0EtxBvHPghZkpiS
4qwaGCHhdDURfNml0AReoY9tlBWxaIFUwF2kdQYUZBJYExAluAuglpnIGp8pPDcy
xbzbHEZHN2i0kI9IHx3JnkXjVQpOX+LcPiCOj6NaDGbz7G9PQ+aa22weEzjmLS7F
3YkbEsb4Vajzbs2IGRKqaNjf+tTZAO/1BAjkSaW4bAEzV2czbGghh7qHq8hckHHY
BYjI8RQ3VWEpXNZTWKYUzEe6nMbBEvNFnVvhzsO+jDhkFp9lu8zvCjiBCFh1YDj+
TTglbKkiUlseSVfwm4ZkWVyjHyq4F0T1D9HaREs2oMeCBkFe/Z+XON/VZWw8b+Dn
AQqpQ9reYDL1viOHjrfivnpQO8KIui1GMFW6cdR/hkXE2ZaPCPGXsuuc8ECpSW1M
oSfQKNP4zoM3tz/ztI7iP0LrLCT0FJ/TIJ0/THN2/H5BYe78fPOY19ZdVVK6FIRa
HOC1RJwL+eLXuSTIeT1uk88/VZYPeJPocbCGvjdK3AW0NRNQu5RnSMFAjPF98+2/
AFtsg0dh3UQHlUTlrm+SA921pyDv4w40zJZdMnrmcU2IBU1U10Pi8OqilPRGOVvj
LXmcInCFzHU5uplc350mEDKdFzjxbLFQKqx3GBvD8eU6TmOqF7O+jSXpQXdzVtvc
wjzjvhJtYRNGo145jDgXgmRgDAwflxXO8RJ8VMguZiCe2LV81WBxO2mKCMgeUsRA
lbJzgCQHkh+tfWW6XdCGJSiXlDOcFe12EHTE6o18gcgkBoDmB5hDgofSpqKFhjG9
A0pQuvC7+cdBZNdKX56wiPRTyF9UEp0KuxQVsTWbu66EDeqsKz5bE8nkCsY/jm04
GeblGWxmx6JurzmzuI4vn10s+F3JE8bvqTbjaFDjCS9U49bkDvTnj1s4qs+36BDc
zuf/IYz2Kj+AnRF2lXmoEq/BN78YGBVjv3oTiXY1vHZ+tNBTGpM0Ti9QF/TpMrzw
2xP+wWoyk0Ngxo9sGzoN3pRx7K4kDFojgtZzW8zuE37QylXBETd7ijU/+IrXyUv6
MAgsF4DZaiLht3CvkVEfbBBb5lcV3VBNGRMll/KXkCYRzBXQ7E6GuIrVzVQYrKW9
+BZQeNYuJMwGlgYS+gI4uQ7LI4xKL0tPFSqFDgCldk0cj8dhytRyqk7rIj2IgyMD
arYqNWQNcQdeFIpM+11q6Pm8M1kWh7EQpMJFK0OrGN0GiMEpbNWskbnRhxpPftVH
sFC0P3j7Mw8lLaWoojT5ymzHoI50an2XwkV0j1LcftXsDzObsJgYtiCiMFJoQt+Y
SnntfeINh0Khc5u9P5UbTG/WT05tM2PtuJ2YhTKes+P+eltcKl1IRgiNRNqwPm1m
MsdDIktw6TG59StUZ2Rbt4NZQPe4nF6q7q+E7ZfYuz7sQdtXSmLb/4NfdZupJf0G
g9bIlUzBB5x3kr3xv1ZaEguYWCXTW9e5VYW3ENA1PYwHzdnNGmIL1CWTqK7oIU2n
Loa+e1O8WeTiTfWAgqraFhbMOBJNiQRfQeeLMJeF6qLJd+H/1rTO9uArQUqbVoWo
dAYf0Ga6LeNOa0DgWbhSQ+c61orE0Nl71phI6nxZX9wNRN9az9WO3WX5KTVZ/MOq
r8BzD0D4FJ5hXl6IoA0IuY7THHJBjOHQbQUZFFopgvAjzlFxCA/hsjja7wFdclgn
tClSM2WO9UIiWErA9fquVcOl/mORbLwG9NJNp2c72rQz+ID2NgCetEPuV+VnmUg2
nLs3Qb+7+NhY0iuBss4UAayS4rsqTJzhh21xgstUWpHHvi2mmvmvmg/IkDB11O09
+cFjQP1cFFAtjvyayhzI0iyIj20yMyocre/D5rmBTghCvxBdJrSL+szTQm+4iXiJ
Z1qk6dWsPnM8CEb3gqJHthc/KmXrSSauh70SHC8EG/j3tbTuSINZGo1jUHXIAVVj
+MlHTt3YFzLbqYjqAaaQNh/5WU0AKlvlt+gH2LW2uGcd5d3LRT7mOh0tq0tYkrTV
58monAdw3VzC4OpNCTtDkpdqqx+j8hwcOurggS6nUX15L0D3XrJ8XPuDgyt3Hbc8
IycaAaagDn5kdzKBRBqNcsVprOpwmiPoCZsw8Rop65v1Q13cvb5hiVU4fGX9GM0q
YoEavM9m1w18bxVBEnj+HiD0ynkA8EOO1pZLuGYZrcsEp7S9GTWXM75ipTT7+C8q
Pldmf5ClfCwQr1IYeIYns99txbOfb0xyXkqlHRyA4pdGaCuQaRn1u/eYm9EfExmG
xRcJiwMLAgn+oT1b2irhG2I+/5Qktvbp8Ss1k5RVo9SwM3SbqT7NDSjNin1mJXxI
9PN1wJ8FvzxdZJ9K+mNVqpHsTH1LT9C/H63ml4pufDU/Lk7UHBps1hJgD+Zh+eTQ
pQuRTluhGa8f6wVBbxAkrgrD98oZWvSGuEEINZ/dj9HAXxp9R6ooXoAbQdVksUiZ
tDk1E8jiWdON1sgyQPZrUPWuN31ELn3EdIPgxg4ZE/oqmQM69i0eQt0S5+56wORo
4bGdhExMZsYIT9luoc3DUsxlAqkoGGBWjqP+VK1Z5f9O5QcyktW2tfcHAc4+yaxR
yF22pOUsIH0GSgr1GcK9C+7bcJhhZJkkzcQ089HFn01Xcjvs63D+chX8KVS4uRSD
Bc0rJaldfUdF5mfo5HwLf18xH5ei233V2HsnBDe+EOrWgZw9c8BGrio4zyHdhWyW
EVyWGrr75rthqNcERYnZPzFsqRmhAf6c+kZRvf7+OGtIWkybyQwgepWE5FXNxjcC
cmqgbpf9qo1IdZXk2z+I5cZIPSjx2chSVRgyHVPLrsACUdoVRFFObK7MXvY0R5Mt
HPHb0Y5gXurQnRZi3k6HkIX9lmPJiBcAj2KoTYPQSGfy6bvlC7RAOxiB9/A/d2mj
kCk+sYNofKusLuokt07KTCwpvbniYO6XM7Jrt4cxxlzdt/V9WbAg+SSiYfskji/O
2KDe7w5VRxCe7p0kJTnZdBx/w7bfVfEg2pOxCJ2+kyo0NEt2nA9G4ru/y/SqNfFC
HszlAyzLYofpqZJYcSwpnyli7DjyuyS16S7lEowfzWmSK1IDUhetDwiYZuWXoHFR
BGSld1FStG9PiNnQf0FCOOH/0mHNO/3FhCr/vzvjT8mBw62+eHPGVHiE+diA7gpE
7UhEbbCOtcVsUSW/RtAN+cKSFRxn0DKpufb4Xa8MOQQ7HcJLDSWSlbw8YV9Ut1c8
tBJ3cUOQ/WtnledpuxYa87Gw3Rg1gFVTUQ5XycVAYMUN4TykyXD/3tft4Eeyub95
PDsFVq8VrydexV1uaWOHHIh5YiKNLuAJIojoDVw3Jd1PtsEV6/akucWp7BKSDjMG
UsmOHlk3amrA1168mRpPqwvJgZow1e+ki5540T2YbvwhMIDs0Yhc4xpUy21PWDp4
+DAmh89V2DjrQQ+WOboMO1bUVz2yIoKzdM3qmns8mkfc822ZQW/mu+RAe2+X7C66
VFnE6cYIrIL6QyeMbUrfwak50eeexfbsqkbq2bZ2bdJzlmoJyRGNwfFHlaONO1wj
Wg0z4foCbB4ARh0r+wqnQ22kPDD4OQn/azrtVFMJvUHYx/D3uJByRdn95qOSL5Mi
z00pJFP2EBMQdk9jaJEn/uOAGP7YEzBpad96+MaFpbU9V4cp0h70J75IEDe+nZrS
KNBRa8deMwheZrfGwL58ZXrdWftrF4DHT5R1NxvSgRqshl1xOslJsNIAhlo159/j
PR8wQT404aIQbCu4oMDh5eoNOOh6VbzyEEowZX7MeHPByiAt4rVMulkJXe5TmAby
RHL+QRaR/iKji527jpLPZvOJOKt15Cr85TuT979jJEkiNLI0qBphNDhTArMu72PX
+t5to2P979RYZDaVhccy4+Oehixe+ZVjfRdAx6Tlf13QkblnL4uQoh2HwJmLfwm+
hCBu9EIkH3H/YF2vcvErA3mnyu8RAhGxLkNGtCG3HsGdSaeinxBaQQjndsnVa+0G
Q6cwSF2g2JftJT5kY9FtPOBJiCVci2gxqvch3TEro5ZBFmCtd7mY4Uv5PvpUNlp7
SpcrPGyOC69x7qf3bJ/sKD0jzCOodsolghCbxBz13ZLy4ier+K1WRTSIP9jC0ilE
AC24Rw2NXMy1qPYxYlHCAAd00E0A/Vqu7N2V2IUxk5xVmdnGXI8PermoW3rnqQzv
V8aVbDpm2bIIBqMrME14ZWe+SYEnCn5UYuaYAj3FEHBkFamJ9NJyN9Ln3TjDEpK8
Wlb/WGTo0ISx7luyBFgNnJpUW0lHG2W18rYQaE5So7rIDuoXls/qrUmrrrFN3nbP
WQQCe6yhg25Ez12NgXg6oXH7v6fhkCRBPBDYHvumEVxabkIcZn47CpVe7CaHW+pm
0Wa2nL7q3OeLKFb3CoQ1j23ZoNbp2oQ5as7TBhiJNAlwf8hw/5lmuATD/ba8jt0H
Js95IQd0MG7ICAYe9KErbnw8hSOS7/E3ujXRdlZqsZ7N0BnQ7VyAKG/Ngz+l8cFt
o0X7clsL8XDL1cV9d2NoJgHuhxE/IZ1sAdn4eC9P/PC0ABz3d54U1NWLgPg02QZO
vU9yBEL6PE/B5quxwVeQ3l9ucZEIuVwmV+zUKwmCFcz3wcoxqUf/e4JcP1e49B/s
xdpWQAnovyy/wTep5yeLhRA0sz/9NszuZHDp6Ev3/qr1CIXy7tpJYXM+Y9SEA/VD
lWq9lyIGPKUVy27cGEWp6VCbdWOfVePNdesokuug2S71hrKt9RMfcfd56AnKTu7Z
CXdqiKCe0FGAMe+8zO89Z6ezzRWdQFgbTdLv7JgujqsaHgDQu6gFwxLMiaeIB68U
Qzbi7qTi2kfAfo8kwZanW6CgoRGZBHy8TfZ52tEMyfW6W49+Xz7e/dgnCryFcj5E
6ckiFP4k5QHV/xL2pVblnIY8xMQJFcfFd7HpTFhR2qMnTWkChUbDbzq2ttf60sa/
W3ekbc4wift/9xB8KLrjuYzqdWatmmaY1qNtHHF25kfBNAo2mqTBYX7AVQyOLi0c
T0zAlLKkHQPtjWHfv7Dyd4pgPto2D9MkX6kUY1DqiMdbTCtZevdxhSSvJH8CuSDk
UbymZl18K5eVZZXEiZPjZOhkrPHEhFi+wxJ59rLXeAq31A7R08p8DpUw5Kb7Gu8E
G/4LtKrlDbHDDmPUJCX49HiU2the6bGNh1hEAc3swKwPr+1JN9rwOeucR0BMs9gM
LbQXLpf8gODW8bFHMgvXZYJfd2R7Q7ADl4OxBJu3+hKcKCLevl5nQNt2KaAX2JBP
TdRfoL+2OSkXwkCuKj0zDKFY7WcnQAlpALuys8rQvk9M6Jy1P6I6KjcRx7oj2uH2
+V1bOsnkyhYRA9rLOIptD0uJRBs3YMIfIkv7F2bCm6Q5U3MGOPtSF5WwtsvIvQmS
dNKr+JfnXCQXoSK7oOfvxVf8vhalJhWpeL2qKZ2bg/NvktbLrDShAnYvRxHBKXYQ
wsRYQEavtWg9q7F4x5FxrSlkqj5YUa6cldfhsXZ+5CjVnbq6vkgBCYx0t6Y6f6p/
pYSx4+iUF2/3MOkM8XyhWG8AvWfT2taTDzNQ7Cvl1ozLHKKBFN+UKwAniaDROZNo
vGpuc6z7S/n/z6BLhweOmw/Ju9OC0BaRfPGddq7ULmm4dMtzj0FyzG2SjGSG7O5B
n9Piu3ydJsJmBHwZoP1lzMQDKr9zY2wik0PH4tc/SXOiIXNRZ67HKJDB3afIMIAu
bEGarA0JwfzWldotwXmz8O2qWBeRvs1Y5yqEUsAaB4NBp8x//4ulhaEiyY43Knc8
Y5sEHpXYAkBeWnLeMnsUgYgUVEg0YvXaeSEEFIN6gypRZMtFElOH4jFjkksF/iSy
+LkNjFwMu5ZXtX+zPkXXQjwGTqsbcFzwTdsm38YckT7sY32ZgIISB8M2bEV1mRlt
u1H/HuRYyVSZC5YhidgET9i+HGqkdseIsPuGf7p1EYH2uR3/5veebkGLauiJVMR5
FFrdk9paHW5E0kOnq9X6ZdPkISgFKeFc0ftiJ2UXEWgKKsFd87hHUCrnhxqlIVUY
F2/TMjUAH9y/53eciy3mTAMa2FdE/xFVoKenmMF6rY2+nRgs8Deg05aMT//VNW9u
AoSvPTY1i5nPTzHY+EYyAh1GCWMSVkhoMSIIiCj3nYYtU/YUD0ogQGp2Up0+U3eL
IWbSM4Em/DAI0Jy+TXzyDnnyL1QmtjG8hTf4LBOEHiNsUxhc8p0IOt2RlW/l8zJn
9bTyRaFjTLefxR9JC/MNbw/SbfzlJwq7rlZTldjsm6qd81Q6pW8oMgvXaNLAwKoU
00HgC1VyDP1QCYjiY0ZXYbpRhKkhngDTBX87pnUDnBGPS9uMaBNt01Pz8+hyJrvD
dIWbExSQnekh8iGxjNViaWjf1naobcreafp5c5eul08RMaQNjF5DSDQGx++kfxmx
kWTvJkuTzlytSovyOss8WlM7XHPE7QCsmXIqqfssxAVtP2PljcizCH2XDcCmSHEY
vn7i7f9I3yH7KCawlgzTSTbm8g40DDNsDqoPuqB2EWCdYMK+bYyJjWMk6cG8yNlD
6OrHQO22eX3TwoHOAGJiekpZKNG3nx9wm8Cr4rouUAHQdTHBc4uuR6m+rVL7EiM/
4Blrc2VFwztH8ztb4Q65CGSBJtv5OStD/3Zm9ghRhA85cuBmbT+KLL83kea4NDn6
Q1Os0y0L7GRFZkVTatx/wJAlEc0WkfjqqnvA+Mc0lWDM1CqqWVhGBrJq7HGLtSAC
LOH3NujeCB2zWqHcMhPnxRtwNaxecqAJiSeDJIMabQ4M/yaNokL6etWsCckiCYP9
U8rywX2D/D6tcGtVs48zH/YKbX6w+tq+ywFkAwe+1ZvPGhfY1F5uuqPY5HIYzRN7
w4wPIr5cmcTm86tZ1XwTcMBd2YoutuZ42HtY4/l+oOAigBk1sM0R9DmZbRJpYRbz
Y/PIPJgMoT5rl7cUk3bv3U0/VTMyyzns6zHKBnCypWJm828V5Uo1yK+uv2/+COj9
Oq3ZlWB6AHyTfGjWnCIsWOFKpZLphpa2J1PLoAXa8FuOtAoZhpYV1stE9Rhzq4IW
Nr5Z34zgOmtpiec03jYnSAQSrZo4CVVVNbmd/6u47brvI+SJ8a2sYIbvPotR+bgB
I+PZJUoGTv74j5V1bw7OclhfmdaBG58KsMvaoRu8VslExovxo7jy1FAd4Y606v4u
Rhpd5fG6gPsSwrnFipYfV6p7RflS2YE5++DWEsWyTR2JTmp076XKVst3ANg29NgW
fxO2C5zAlw1OVCUuePdqibZXoBXnoM8FBhqGnrC0Y9PBHLZueazdTVFWBXD6qViy
OGG7jN3NXmUayJaMcV0JtHdPYDc8+qmhrK0Gyx4z3B+c8cNUn4272vsClFikjdgP
UlB07Bf1TfAEEwk0RZEshlp95WQBSLmYeG1yCjL4bxfHe22ro/nu9Dkyd0kyKsV+
nwjn66ll7Ppb8xuckZA1XKD9ZqWuN/w6Qm8TpNB8KHuFweZnP12ZwCK9FQDszTAK
AfOh2kbHkb4UYEI5OHSn+2KBgDnZh6Pb0rkzx1bgxFnu6Hc9Kptq8vGhFjVeNy65
cyWiYXkaQVJsG8HD07nAilvpqf47ECQ9dYuuutEzFRK9jbbUtFl8YcLgI6A1XsuP
Vfl+wUdu1G77StR+AqNTbNNtjLPy6oJYuWUpt2wOrEgo6eE3OTk8GKsabDcfDlDG
2YVaa8pCs0OUKWv1iy6cMeV7LOdRGLNYqWHKfA2eJuiy3dyUEkKbHtnYvkld/leI
cBXqQJ3ZbXc/CWqgb2dYurRSY7PBLTYz2bByJFRr0JSHlcntHlgzrF3WH616lDB1
f8K2e3JzEwiu1cUoxiyGnQHWd3yiHD8n9PzcLzT4FwKx29GgllL+jEZvT/D7PSLH
eGw2qjHUq2rhSTu5OA+yxILU0SmytLDkLo8vvyMYzOcoamGOK/3+1zMn+xoIC21n
o2OQEdWwGey+QIC3D2BWLOc8qIP164HbX8S1GJY2VdkHr4s2RXobXtN5ygDGZMWX
mrdGjhvNVYcQC+KVi+mTtgO9qLKk5JlNXwiQVr0CL3Nxioldf6LWyYC+msLs2UFZ
Y9urHTkpCpCrWyeyJj+afREWc3jPQPsDsMyxQrWTP/La5LZHbBywlZcB7jJWRoS4
fW1kU7aj2roHeChD4XvUOcs0DKpRd27IWV8nEaRLNiZE0YAGPXuy+BvFR0Owl7vc
kTN9tenyyvZSLnvd8GmEPDCrPMpVTkR0zYCZ1KCese0+gQaR7hIntFDY1QyNJWoq
qtVPRmEq3h97JGWJKJ72+cT2+Rtxs1JSn5smf8O3j+o1OyfOtctFLJ4ndrq9CPna
2zkUDWosgJDui5Th2fjwAc4vtiTZOLpTDRYS4Jvumvul917dJu12kbTwdbjBeOer
+U9si6yhNxoCc1TrkrHJA0WqHJTawNed02nO2183ckqiytSKDkQNWfXuJK6RwjxX
UhNvJRxCfFBzwzZg7S6NpfnBrVASXSj+DcqGDAmnFaID818m0quxPtey05Zlwjyx
ax9h2bX9vsKzoQViJiX8Co4ULQnxtOj2+AMlDNUydfWbscgHjZMeY0Td/PE5gypi
6vY93UpqxQo5KOTEls75Ns2inGLk/cPcjqYwENccp3dS/gqgltQzdoAq3LugGE15
ePCUp0aLYHbuVuPV64QHThTyzqc9N40pKZBdH7ZaJ5Oy45qOmBWsvnMySfgcecIu
WpL2fEEq01Ar8eDUN6dr/c81DKUilWT9iYGU9/QXWz4HX3YytAcCePA4FYtUJ89t
Wktx91KpoVQKu1Xml38j+yLgFtHLzOTQ17M7/ja8TxmZ9JLRv1MiSKlL7m2qxe0G
0yLVLufvTrNJhu8owJYIG25dZQvNO6j0v149T27jmOQY85+USRv4oYgH3Uxq8dw0
oS7hRTzqwf5wc00lrg8Wo+jx9zCWZ0OcIzUBWKfALjzkbkG+Usmqk5cxpMsqvDEn
q4mxzvDUdWgHFCKehPDsShn1cPoUu06LKCGDbZBGiT5kj+jeNy6L3JtbtonU4R3S
RVoZE1lIOTvhNnxrmf7T8xYOOc5PCchFob8VLsvG98/Lwb96E5wtp0SsQDD92iT9
0KxlDgqU5K2mYePRkl5ChZvr8TwY47bO08oS20FVYiV4iiYE+LUo94JDyO31PtsW
nH1uVZDdJHgOuqQdjKnH/Yl+RwTlCeCKBp16LpdBRfA6B7TOEtPua9Uyjgb+lnhE
+dyuoYagZh0aL1CG9av5+c8CFqemRri57ZfkuT7s609rlhU/0Cg3EIa855k00IKf
CdD/DuTZElk8sNOmlcD9TNVPdmoPzVEjTwzVhALrrss0Vx2aHIDxGyQaCDdPoIG+
HVrH1AjFgQhy3pk37paYmBN+u+m5COOXLOtSDQyWnR5EFYVFT8Jn35Z9os5G5nPf
n3A+fJAMKwc1vfHO2aHvYm3ULRvrzAINJtb+4Ju97aHRUhMYZt20p/BU2ral2FEN
Y0h84Sfp/YzvR8JsfK+V0xIGuR27Q4dkdXDwOygznO9cMXIsgxwKI5h2NqsxS7RU
2eRSjQKqo2nXPFKRNQkaqU2VN9LWjJby5x9MJjM/ggPrDTqVMpzkGmpAaZ+54M1p
nIRiVRC06bL6zAbkq4gnbYHhuelIUw4z1rURnFHgl6hWXHT/3RkNhucPNTGPwS9d
ox1lFO8RV3kuqrKimnGW4A0iexDkiOvSJTweJUWApi2VO6qvNLxZVLbiavy/453C
AIqWo6H8pfGYN4rQ0vfCU8llHpHzpPXPRUHd6CsblCmcbkX0TfnPJta7DC2ix3b5
rb4FajweHblQoDp2JrEFompLjG0+A7R1vhVwbkH/Vomw/anFHqmTMDzZOK+EK4MZ
End4vXw1LkydJ1mRnfNV+x2IH2t3m0+3/wRfep8yDafhHPCEmpNfpdHXq35AeBKw
FdkU7/7/6VUBujIgSkvhLCnRl7DQCYepqDYr4EuMO/IpHo130sxIR+gR6I1nLKKX
3q+cNMJXe4eCYQeJqAyxS4x0IMjfUd10p5CkNk/KUlIlt7z2owaVyHRHSwGAOT0Q
jLWgJIzxEw/WCi6wXlO1agCHPpGzrQDF/0kyDl2RUhzBw4Hr0xoT/0fYdzdJG3cj
49AKU/GSu0pHLCdA69FB/EpkkB/tqrL5GrjnLgRlh8hAaoP8EKqumK9YlSPlZlf7
D7C4rgZWoMy3uYfYH1rSxx4Uqz8h48d7ZjT6Lo/Hb2lifYT/TrS8IH5EyUAmMr4L
LRvL4NppfJ7P/tMBg6Bv3xuI9iff6LFld7+i27DBRAd0YTM7/281+/rUAHrE+aqV
qzk76JCHzsF0E+Rhiq59siY20C2n5ePZpd45Z6WAVUgmE4ta/Y9o+N5/zvkjbIJn
95ykzwsdypuV4reAVACxAw3fM+eyXPA0VN9ezSY4xD/kaCVFNLUzd/uog72fgKee
/IVA5J+tghj/fWLvMHZwRf5Nncp6PBFESX/53xr87LwmnhrKQjfXBqFZpVkSP173
hz00xtZwZnP0Z2PN+pgarothml+Uj5fm3kZ4wBxNJvgge/HcBr0dfi6C9tcFs6qm
qyfb786PwS3kx/xW6L8TJlwoPiUHKeycMKBIQ6kydPtmSjZpPrVpadksre8HaXJl
DclrhJ7oMx3lUaKnwGvrJOHnINIAOkmhJMzp9tO1jV6y43+z68T+yIOwr5z9vsal
atzvaUQXXpNg2adVHtgHlAlg5t4vhtTagyxD2R3QNkreTiqc17sgrpsU6fWECo9K
XYTGyiiLb+1yWtNa0yqTIGwvsuOfmdG9RK3t3/CJ/tDGwnr8gJewhLSg9k5ycb7c
qpGHar/XepFge3GyfTTpRnTcRj0Hrnfd8PHnZOCAI7T4Yyqf0UXCGS4rjZtvBrF2
bYc9M/gcpt4ugxt2Glf6E0hsdu7WcU0AMe3Cx+t0Jb/cU1Al9JlBM7bB0OWZj+iK
bb9zLlGCGZOaAn8fVLPzSMVn6omnTM5V23X0k4hjB9N+VOvBwUXwDjz8QbWEcrd5
8Rt9v8ClJTxAzgYSADdamSlK0bPTZsKAEHpNpA59BCzUCFVkIrl4YsaTC4a96Q2Y
ZORuDaN/XmVMQ99SseqpRNZ363dDi7w0nvaBm2jE73JqqEOx/Q01VZcB3a/rrq9C
6v29UFCx4AIBF0g3lTutfZqTLDkQ5eDjojloJ5yc0iqsyFtxsqhQsdFBFhEg/UQj
cqB5dlBDz1/Jz/IOtcOv39V/OFhjlVJiv9zF/k4ogI5aTMni1VWusx91TyOkHm/z
/bO87mymwnKEhhKI/QYy/Xtv1pwUc40fAUYVHy3t8BJ9gOwXoX9pD/xIvw+DjfLt
v6sWs72GLr+hoFM2xXHByV3tvVq1TfewOosPSCAX8lxeYJ4mWA9ujDc0ll6H42Qg
YCebyFvbfX4Cd4pRRO88jUpNkvfpoq/GjWzxYjYNlkpW5/Bkqg/WW8QeRPBjTue1
huotO0c/Q+SgRArxmbttGzNrzuuv+q9FBue/il1wZEOwObXrZPH/vAOc//WMbDWZ
6pfdloUqSTj5gQLddG3KQR++s6sKSprZiV055ZYHOe3VEeps3HRhmxArjeuDYn2c
dh7BqwSE6vVJuHtBQgHU4vjirLblXMso96i+B9LKAYbVl+k9Lj2F/IOVglDEDbup
ytoalBqpzBXDSuxq8frYa1JGn1U+ytTWFAB3RqQ1/ftunoeB0Ch1KTiRS+L33P63
K69/gbH1g7MaCizpinxTn91mo1LW3Ai/cAspxoBEUT018oPJ9nSSEgvXlqITKbdT
jwFoE2KTGFeF3cYqSo+B6xKmyMH3DF6MM3HMnI2PFVP4gcKj9tULSm5ThTu4C0nd
L/ZJJSvU7knw8pQ3uB99h9m3/G0cTHwhz2PVdxoKmbhVDiuwmdqmco7B9tWIgQeq
bLkImRbRFqnhLcG6I2JnZT29frcNG31zv2H+gLTWLKhn//JK2R3arkg2H0BwBR3i
xAL3s+adC5WufJvxxUdYW985NJJusilrV+3Uk7PMNRtzrlp2kKT7KJT4lJgo7pMY
nXyqfvysJocKUOCQO2T5xTDt9mjALaz4qsiLwz898Jh3Q67EecuS14KN8UTUol76
jYHceb9XJVgpr0oAKdZVAcSREmZYn0xw8L9mHhYpuUv9K9ttdMOQfRZmzGzsXtFU
fN+oUWDSiVH72O4wzCN1nyKGd0IlZSg5Xf09j2KZMAehh4EWgafG8wjbZACY6TG6
N1zce4l3xIJwNphCw4TrjF99yz4IG1+lS92FAoGGrRKau35l3tAImUih71O2MMlg
57JjkSVn5XOd91Wl19c4zLWd12w0gUNf+Y3wA0rlJiFspYjThKbslE+uUYqyEaQ2
sYqtsA8Xc26E0K5FdL3vJ9qe9HwECLMzvm4CnL4DRSo6styjcHkiNkvNz2ZX/zX4
zG9ibcbo6PPi1T/HcjqzY5Z5jDpdAGWKR6jJpD21ZNoQCbtR9t4en0bF4YFutAxL
9unpkgi1g/TQw/EytwHIoUHggdTTtNJKz2BavQvtkDwnf2hMb94LMUOENvF492F/
ZEJuSU4FX/itZiCqGN3Oxjh0kpfo5lvKCs5JSACs5lCvNkCJxLaHt9tIcyOqK0+w
mSO7NoSfnMItv1bjwVbA1AZ+kumTkamt9VMJIpHTgr6qPjIsSiEecCzTYdvlJbXD
/U1L7xveTLcXgWwIa1+/Ha0dsvfC9I2BQrjavrcjv3Wzv7vloKXYfTvLVqpQwLfl
jl+uEjs+n2D8grWmsxVoRMtpHgQKG7difKkc+d3EnbQqgzigkFBFb4kWUI45CCAk
8dqD2OvFmsjC3eDNR2ETn+MO39aslXerXBon0wycEIgUDNgevo1QhWh3CuhShKvv
V6otIX4BMwuENxGnTBbLO6wOmxDqtniW4wQmV+6nPiTAnT8kgboSRKmKRs3wTrzN
I04HjmrguoldppPZ8ngg8qXiFsgyxFf+eB7w8M3iim3YqK4i3ltBmCwg1uTFMQBC
wMWfEPRgQqkM74+l7mmsl5j0f/euBhSmET5TX0Tn9IWbkoxxCSIpS1LqYFynVYyS
2s2FP9XI/uKbrUI/JhUDzQgW0akWE3p65nTccS01j0UfUHrdBIxP8O+tellyg2zc
dA19NR5HMH9PADx+0zRpaZrVi+5piYId4Pa1XguU3gxa+lhPZ+Z+/9bBgeRK9Fe9
n5qYuqGN/mrVbmlZyRPldKPsgUCuLBQeJ+rl1febaXOA3IP3KTvaEgKzwumBY87j
72l0lTU2QowAah2Jl6I2fU4+DJ9txgHWkfEG4pu5ftnm7nR+3JGod6E6zu4vb8dz
NMiXgkPDwDPQpQein/G++gtO3q6VqaJ1PKQfmcO1kaaxIKs163c01SLB6ElHYJni
N5msr++7AM6H6XA6ESVXJa4LYkq01BhypOY2c4cEXHxLyeHiJtyi+UAYVdm3NDi9
+a1j8g8uHy8jx2VsZU21D3Yf1qeb4tERUn+H+DcCm/baZh4mG6sLIxiTB3B3ytwg
BXLUVxl4gdbFhkiX66QRucwlGpVXS/YFtMPQ0xKoEyYRKpPlAWjmHOtOTRpdBoGK
r/V+eR3sI4rAavofeB2zIKOEnzXABJKCXvDIDaG46zYjQ64GcQkyUw8CcCiKW0tp
LEmuQWpUZNk3JY9rVlunG9/j2bOmiQ6VJ01H9KLGRpB8wLA/G9zDM1RkEkbtoTAt
mEOp/DtXIOxkhKwVExm4YsBFA70fr4qdVpSEYf4UeIwW4UqhDVjYLQkx76K+6hSz
wcv0UWnR9yaylzdejHwbsUZRF9c5XesZKD5/m6MwUUF+KVafiKNoU2iCLOPsnoDl
+b7ZlZ80g8xTYalHckkrOEY09j21FDduc1Pfz0eHdqFd1Ik/MdTCcj8bxyFcljzO
57Yx2q/irZC899n2UuvoaJz8XIz0gYTulg+EvUf1YRlp22FCa1BbJvIatJYdgEEz
sN77YJ2O3mt2CfQcByNhoEqWDG23SN2Hl3+LVh5aaJd6ooMnPYSMXbcVN0Ms0hOY
NW5YGpoQch6DlLvfmDjmqCDqvmxg6BCWYTtUDtux0wIKmKKZp7cWZwFKBiZn8bTu
TWy80tQZ8PPmdZSKx311nJuKBfR4O4itlxbeAsV+CKNABGUzouubDJ/+bEXhDNcv
wKEYbg6xn74bc9F8MwvSTE9JvXYbVUFjFrrbTKeWP8DzdhON6SRqnBBQA1S87yXW
OE2vesoep8EzxRYVA5Ehxe+YP0wFwXkjQ0Oc/h6kEwUnN2KIl7Hva0AiFNBGXhOE
YLvTKf2RslQ5vwc6J1GpZ2qUtqz0ZesZrd5cBWNuCJ/MxzMImVm+y+uo9+mIVPf6
F2joNuCbVLjxZ9hL7ZsMg1r/hebddX7yRmpD3waA3lDPHND1+fmUYZCieouMkvH9
dYL//AbNGqZ+gkfm2PCnUNdo+OnurkQs/VHAJUnBtCiw5bYO0flZw3/RJyf8Ze4X
9DLZ6hu+GFhM/MoT2dbs1VRR6jrGzDIuAdPE98cXQKdNrRATQPtc/PqzRniafvq9
IgrC3LdMZWpMVxqP3gG1vDrWTbVCZi6JnefThixKC7W3F2ELG2vfid4c1wDRvwS4
jpcStxWAvY41Cz/uuUcudjhxdtC7S+1wQsHD3wk5hIeTMttI/PXjikp4HyVaLWMb
wvBvas20oLy2kq5vGmXlVKtVUazvqSwhml2KRCR+u7RsGxARwn/pgnJ2KS6LZAsA
VnYNm3nqi3EYw2KiKwj3JkGEy3Y2pT5Nj7fweyV4hsxfqEDO4IwlEk3HDzoWeGNA
E/S2HxFzWSG0Si9CTpXfb4kShiw3U0AL+vG8eDwKV3YCrzZn3EVPXAPBJm9CPYRd
/MeZkOuWyW8SpZe7Le8wfyXZXzqcEyXyh/pZlusnGdrPskCXjC8yMWsEFlTvEf2l
hLLlK/26WMVArU4zCnufTYMKEHUGkqARBYjNV0Upbcz71oYaeU0IPvfCFMVLc0Rv
wDrME3ae/p9djY2ajXXLoO0BboyqEcPAzZXZDAuV3J36HmP38mCJnYygWR4olrCm
MvKR8GN9rh4j9dsiMLv08gnlh0cy52N7rlIjy/spbDQ5kl+0/Co4BgPw1+91mxLt
MgYiUheKR8B5PPvLGjqP8K5SRpFidapnxoaISTKWMHDn0L1lz/kFfXnwxgXxPPzh
SRTVoS3Lg8zaJqzXxVBg04oBBd1GmqanxKdknBWNqm8iHhAOp91LxUFZUE5mb6fq
vEWn2y9hNtkxYy4zAx1zIMfJFZoMACnUbRUZMo3w+GGAVMkx01qfboPmbaTuUM4S
P+gKsWZ9sqEsG5rxsQi5ccl8KD/8p2lIKXrdF19wfk48S2OqdvjS1qqL44zkTKY1
xzqFnq1W141DN+H05bsylrr0w8Vjcr9ZbFlsZFezlPSV4Ef6bX3WLaGRr9chZ692
MJYkxCp7fMePK6ZnbszGmNLO29T36FTNFkv5DYuQPRV6TZqsajDtqs2wPbyymIc/
tZ8s16kvW/qPs56BMPf/a3W55695Wo8kgHJgLlbHg/PRY7KPvMQSzJoQ0rhi8TcJ
0N2zzwuPyFM14hpw6QmdpXGfbydhN9X1TBEqVLuiTbA3kS5JlyK/ZwtYN5tfCn5/
t3rCIH4NWYp80308A7nb3Vlnp5/tW30yYztjbgYdpkfrG7ptUN1SnBCitEOx6EGF
mLUicFK08Qy2ZSjNwX13hrojXldSmyhI/B5YXYy/AX/k0lF3UxYsv8aSL30Paw6y
qL9rgetPjcknYxgWwzeV6NWxHgZdh2x5s5G7XFgz1Juk6doRMFh+sjnNKt75uuEG
rINaIldzjKm8fAESog6pjDeZhUQZxT1NhFlk1AVBiw7CzX6E4G6GL+9cKEN2yHy2
Wi4+gz9KtVSxwrFpD5VWom6yKRKPY4UenH2bfHb/ffEhgPNIV5Jf07zgLLG7vTHv
MSjBy6L86j36dVGmDgV87K10ggBZSXtBaVUAO16ALVPAa4vYEu5L5vpDSozQ2xzo
pioT1py2bWFTdlu2L9QJEdgpuSfl+yKtwjEAxzNmT9e5KHW50i+tnROdo0xvGePj
LcA4IGGOt65Gs/2Nxb/PpR3qrvd8VCRdL38+Nc8ZNBpbgx8dCQXbuxlxcaxEsoNP
jBTEVOJYL3fGGMlmwAwG8+qkML0kSxHsMNHY69Mhx3aNBb6UBGeNSDgbtJyR8dbw
0W5ceZHxY0UhlhllSTVpP1oNEBExTCcDZZCXwPFJfaJq/W9qxFpoeYE6s3zzdsou
8r/NQA6pzCPRK+/COFjPfaDBxwaCA5yzTgFXSaUZ/82vvv4Y0XjIiLsiu/MYrb2X
7/ozU5FIGpDrutURhp/iy1JRSt3TG3qF/3Gj0GMMjEuNNfJne7phtnlmMNQHX7GP
l/ZKFMvgTkH7d8owIfeJi0ann62Kez+lM/FhX5CSeCwvY0ZGc1n2CddHHmif5DmQ
tHA0IYlnIQ68ELx4tcUW7oTEW7kpaIsDvMJYkBtepNk2qxK3vp8GCrOsgbKOBCVi
7quUGhUOe+L2oj5iAXDB9eu1EqTU1I5MYTEvpgaQWwM+oBUmC0ezshZjBSmZkJ3W
0fnFk8iWBNJFlzf/GnRmLEwjmzc/2lwTMd4b0TmNpjGi6wwRFGVK+bKMP6pRSLTZ
kFYLqkkC/S0iNpGwdNr5WqfH7czMpD5of7VvgaDGUIgFwzkC8N4B+2MWGKleHVVg
7o82Dmtiek+XYIrGe+AtuIOhrkbdZj7wy8w3BVseL+HoS1CD9psfPcH8fLawxq1a
scSCZK4phb9Jnuoj82TzVyFgN3TeANvxQL5Wu0Ui62/wVneEAMQNzJNInh1qAI3w
VTyh/32pwNL8S/xCo6jj8ylinnN+vvn7Cm2m/fFdgC4kKklHXyfM0Obj2zPAUtwh
5lTiYnvvCNyoDt9eIy4RwZ/zy7r9lFH5IsdE9Z1m9gj6khKlCl3Fh671OMH0Bm4w
Toc3VJBBnHynpNhCS35N+U2fal3R3YLzrqZbjyL9kW472HIlSNMw8A0Z2+52OduF
3nXg51jsF0nZQpxTUXrxPawRaoh/Ub0iLrj9CrOPuagpdvT5OgwaZrg4QtsjWf59
VdplBuDyz6Lt2wEgFpqtMAYOqoKj4dIlghpzEnirM88tAzvtMjyUk3/dzkZ1YN2l
ogbpdxnc4ocINRZkE9EjA50WhJ8mAZFRw9t78d4jGNapAU6rTjoKRv77nEvAZaZ6
G+fhIgjKPpfeKuGy65ZlGLSaMZvmp5jyE7rnWVXpN1AEYpcBpza9a8RUtPYXWYnC
OWApgCcPou4evX3p6cGvJao+LWuKtigKUvujPMMsTT4QWF5HJPG1JUm/QE0IqE/e
KGozC9XXi9iiXQU1Nc+7szfoM5cydE3hruz50sCvnwga0IvgNkX/srODSP887+FE
+bjdRiLAqdavAQLvOtc5jQN7f8w6fwIPXMnIx5/HSXn/BGo5GQncyAUnzZV7KnUw
fg/wRbW3AQXI567B6rRYfSxHRcFCi87rPaZG37xpDqa/AxDtYzoJ94MIJDTMOg4z
IJ78tFCoHM3Fh8ftkkjLSTs+OlwWTzDfeYFaiKpx35Rl9rfQF3s2FDQUrImq1f52
qiEOvXySjh7RgkK0uuavOA628PREYf+ObaHbfUfbsdjg8mhgQsdcJdTKmZghbAyR
4sfu0xsGNCCqNWANfoirQcbIC9gMWwqu/DLWutfFl5OBtHz9JphmWfgpA0alRx2F
Cra5M5nK4axJF9UGsJa1WltH07eWbdGO4DfMSGums8UgGZL8rUY8AIt3xoSbn0iM
3BGx6X8kVYtnlXSx95EGSTLEfA80RUNWshAT0aW5q2wGcdT3U1v2J8FyYuiQTby5
X1bEbp7/nfVAeNLaIixXaTCFgWXagtbDwRXzGZwpOU4mzC4lUsg2R7M2sk4Z3hwL
/tQ+swnjN3ZKJiAlqxoi1v3J/YvEJzPEUuHJMTNiUuCmchCHoKN6IoiYRtR57lYG
14mK3z6UJ1MZxCgguj4D9NIjIzE/Jo6Vdp6fSgdygpe6htGeXHJueP3gbeb9QZfB
FcTYZ3DcZeGeqyRClEjYfV3H51aOFuRinZyHzZq6frUMoQpadrCSlmbcS2iEZCSR
++FPU2wPX5ynH5jheQ/w7s0n+kRmfI2sst0V+YLV9hNmmqXE+a0C4xGxzAU8lfrx
HpUd13AStuU66D69gJSXRj4IRx6cZJby8UIWcYCuwXwgJ8foKtYZkTli5llrSTnc
B6DkqE/x4qycHCjQ9ykh05ix1CChSfYMcvI2ibUVnDGUisGl4V8x+5/1AebrfOBD
cVrmY0y7GF0hQXNkfNzYc22s36u0ctLXs0DISzmd5+XCXQTzVbsikouPcDfMli8d
3xQqINsMuJ4RUSvFWwNzAQQl8Pjcl6J0y+duuTNOzk7vPCzNthK8mWHR/M1TnQHU
fDyyz4Ohofs7PuYi1409iVZer+8E33IaJzx469I2dn0S2CcOxoDXT+atj7MWddQ7
UbF08/7OgeuCHrun5ej/SYTRfrGe/3YNeETdER5DwSgAQfpJg/bp7USZShMYUcUO
AoqD5iNFacnXnIss5HDoUlbzVAOJlV98JpRC2kZRMMFCQ6cBP6OPe5wm4DVz9bvJ
38WDr643i3OAXdi3euBn0oMVK4ZOpb0YLCDTPb/j0ApyrN9cBdejEQYP/XIE8XNK
+XlubVlTW+0qWznGl1kVkXQWktGF5wj4oY1coay5qc1Goe9vqUoP+qviof/xTOEG
+nIsQd8unoXn+VfeKu1wZhQKmS/SmqhdgiC0p3nS9ErKUO5HfjjtjTO0CJ8Fg7X8
SJFV02WX9BRyJFv6DLUtFJPNLI9dy0YbZ+jiRqRGKTNGmHYgso8luNssNVU6QIZd
H9a7g4Abz+GkzNwHXcfQN7Q7IFq/2xPKP8/3wM3syPx14Iz1vuZF/CJKxWux6nCF
e7p1YOxW3/az1MSJBne4FeWGuFHwUTxdl2l+bmivTy5bOhmf+NdFOQAvgHReoOUE
o0PkAE8L7w+kKtCvxa/+I2wEo2IG+GmOIUfIHog61RFta02S5hV2HDY54OraHp+j
OdZtrfyfY+dbK1T2Ie271z2aZ0t1do4rHc+BYOaZB5eyvoFRuO99p3F7ZGJpHWJd
NWu4ZCPypSAsYG7Q8O5dyuspup2x5nTHdDqj9zZOP1F57RWJV+NYi+CT4uYvIH9V
aMbsv9jfsia0k/hR2SQnanm6AbR5xSVBOjkQ1Z6ymBMIiR921iD6hrLH3I+XYLDS
9T5CV+0C1WQDJl6An0kg7AzA+QwQi4N2YMhPmXAcKmFBIBki247CQc8vzat5XCBO
fXqfYVBRUqTUGMYOhtzV+CgWV1tM178A1ab9hvWghKNjp4ZSGkJdgzChZPzHpJaw
1Y1o3Z7gvXMwiBU2Q93VaiLrLOoU2lO5RNLDoEUVjOCkNP4C9u9CsZ8QDBSIxAnV
zLBCDzxAbM99u1ucjXocZaH2sMIBSoBayG0SRg4bZByNxJnBXd/57u1AZPsB+fmz
yRG6+RgCyZtAMusEBgsG81fd4B7zmoDDCPUR8HMwMMwI1gZyED7EcWH56RHwiBN8
YLKns7ZyOzwP29u+1gHZDsjyNgvNdznHfsX45sGhywvLPRu6PWFCJOcI/IakDAv2
ee7ezBpwFl1tLGbh9d7axgHvVg2i5lpCeDrd+jvfvy4yl/E3WzaDeUfIwXVnen0c
v3BjX6HB53w0NNJHTlDTlQxmDVJOJHEq5j8OIiyv9+iqVrBMYlZMpoj1FnShZek2
kc1EtfnNvtnGU8ExvHn+DFJzhLIVdApRLBqG3Dcx2dIIKPjj6Q/ioL7KWikXYXzw
UBhbrjIYAp9HBkpg8LHR8Je2vcmFXb/PuaQ2pf9KbpoJBUlfKmqZX0X4wK+DxR/c
OkcCJELd0kEvp1MAUSo6dvSpcmysN3ipwFFQwkzdraTZgQizA+Rx6BF/ZKK88GFX
NvndsVJaJW8qM4rkJzkr4WjF/nm3714rAkFvN0eAD0mzzUmZNgLDN/KaOFwl4TjJ
73qQ9/0pa1116afr7GVtd6oNS3ffRlSg/Zcc7cTatDPWoQm0jaq5aKZ4aJ8jjxmD
BdO13B3F5mmHUqGNDXOnXEh9qggpp5/WhzDks0JfSwh9jBdmX4naeh9P4zbBPBai
++SzII/p3aEBeUYhnJOuH1y315m9Dtb33i85X+/2O0F0HDhas+8Vs5kRcVZ0Qtmz
3dATVb5Yg5vbrPvCb0e7/Vf2MGA1pTaYAMSNARRBgmRuD2dkUNwBpT3quRhIsQTJ
CloAE3bX2DR9BDB/Nq6v+DtopwFFLkjALZPCb/S4kDZ291XApgogvLTDIaO6xUD+
8FLzsXEmAAnvXcpJSnGFnqCK4fph/2u745ECQo86GR/1gVjdwjbAnPBgtFex/X6T
RXROh94pzfSMTaKJowa5qfcBznbM0KVFbA8SnBbzQw9qqUH2zvU329Qlzzv+iQO2
Q4214S4PztpWw/dsChKAlhrZLlsxsAjOq9vCsjCaBh8/uYtOGNB7eduEhj5JF1Sh
lwIPpVnJaSuxlPIPd70EJSNfQ4dbTAjGNFqloAWtsnXbCfZDuv4XS4am/A1dS+tz
bvHI0SS5HDTOWMHmw9NiArTo1+nJ+IlKkdDM++foLy09P59ZsiHWNi6/9099rRjq
fYHKZuDPkuJ5BuclEvDzQ6sAa3pjDzPazVXPXIyTDKTDb6+wiodow3mjBc3uQsXd
pvwfvO7wdqw/6XkkkpnyKTdjV+POxlcXNKkQEMbBx/I+gWxXZWp6yIw2BKxagmjI
zZaiNiTjcdEukzkgrN6AjPApB5qn1uhNEAA/gHC0efAsohXWexrz6LG+QLyYVKEn
gTtHxg/dluL69r1efwhDyT9o+mtkpySmq6nczWWoh7bY94QwiPDV0zNz/EQewjjO
tQXRMUaha5qp5AK+SbJyyYKI/O6rzhXgDY1ZtnBYY9nCm9pQgiQCNaNGzy5IUHiF
02V61AlLTQnAT3ms8hJVl9n0n8+22hqYrYOxUnmxaJvSCY43uWYvNxbjI2l3rsez
aIUF3zNrYpoi9xXw1xugBSXLyIsTLvzWcsOrVuqeHONVQ13ns/KM4GtKdYnXOXjJ
64JI8X8Er8SShBk1zx8HgjMMcdYO0TPfshZVNC6OX5Pq/WW+SJquNM4A+e6AwsUv
RELr2xwCoTZmh1ozc1VR2sRhp7BTAGsJzMOQeniXZ9MyZF/zuI2xaYqvVAHIKzMT
s5AqEgViyiH2Ka5scrY0cRpI9EL92IUStYueRR+GxXtk9Mxt1KcQoa1A9w2A+k25
gX3M/L5cfBf215nD3JJ3W3Arg45D5p95TlWuikhWXDHmbT9akucSX08VsmmPgQ1K
2iveNGZNnhMEub7Dniofn4QQ2wvpbWJ2059JKHa9ZOQW6KJm8Fm7854fUlT4r8gA
+n7RZ00gdA1BDTADC6Z4rLdxAuIHIDOcpxZi3aU0yM47MQn5fgcZYOXndxojHSeE
CeMYpve6hF1vROcJ1K5xZDTvAWNeaXbiFMufn11zTVc/H4jW9lbpncKmbfR7Wyr0
M6Iu9iWtVJaFgXNbS9rY6YdrNHz5hJCJOkWL568DOrNADwgR6XjnoYeho0aeA8X1
XKA0OzO92E934p3NEQbzdoW0Ko2uSR9rIsaoGMclsCaYntf4Px+nb26r/BDZ2xiQ
GTYeGqk9vPs/ERNgoqr/fEKotOsvdWqLVQUNOutSI2vpT/qgtoMBQDmeV0iMdqNL
91pS2fMEd3JGrh3a7mk7KYztLBh3PyjwYn8S+GdPz3HHJiDQD+bFLT2CpKQ/INUn
YUi1ZiK7MB/YnJIdJU5b+EvcNZb2vSKe+SZb7bPuN9pj0LaSUUX2KjRnaHQmsTRW
Z7vcR30SBYiMRTP+GBIe8cafCbAo6sVbuAXkVhxzErIoG2OxL+jFEXMIPNr6Rcqv
Rc94BtfZnK8lSLy4S8SuNVFmRyw6iVzReLnwaIVzYz2wj4N17SBXpFmv4Fhjtmjw
rS2jp9ml30fRJ8q4qprwuRAxI+nA3L1GaINVXqmgk+GGYk0xo+kVc4PI+M4+TiK3
PvbF8FWsnsN0QEHP4MB+FkWa/po3JdTIeCOLmP2ls1gM6WLpHe5v/c5HpyHpuqQ/
l2qTBQzFX1ZCthyTJTopdjSylKFuJTuL/9patiQyyjlC6AWm3oYqHx9rTKFzMuWm
1kD1AhfraqFROhRM/YigL7GIFmlb4mmGj9NxMVqJOvx9GreXwvyMF7222fdUFGcc
3fm7tzI//byBAt/DXj/nDnYOrHPh+YO9as9zg2mR/lpmVHnl7u0SpZVj/b3IyILE
Bx/aug5UB5bT7+3XNHj7hl8galSUGJrgI6uiWOHq9NsQ+y0CjXsDMOyI5V+BF5D/
MeHfOW46bFN38pn8oftQ4eFcXTQYPaUyGG45DwfhiFYIIxEMTf9nhqFIoiAe/QUI
LcAmEmpfI6D1vLFfx36anD2rLSMfvjUc8H1fqD9Aj0LuQFTtnAw0ClyKrIee4U5K
iN7XsmnWVOMTBobrfEQAkizzi2qe0379dd8JLs4oV6JvZyEXLfKi9ThFxXhsPFXB
EnK0jbfwP+wjKFnrboYYK5W537yaHu4eOvQ/q6RG6ElMjOb1so4vw51jsVv9IzVo
VKgXmCgCf12tthGXV+2YpVI5si66gJA9jpwi3e4Uolrrsrn/L6EQ9j4mP3gZjIYl
kdoH/HUU3IRyQhwHqvfBCApPhXY3y1T51riW0L+fDp5dkOse76cqTnn/4uV498rU
ooYZKhaWBXUvAmeeoykGXFx87NBf1DGsJZLJHVjqXEP1kEBp4R88H721qxqdHONv
D6ASiS8EMAEPxz9tzRhkKi0GPpZUFjX9iL6eUVqdnnlxTu2rgn9eFnMQvv//19PF
0OPLH3LOwcVK0OmkQEouwSvS56Lu33/r1oLnvC8MKMBR4yRRE61odrmkw+L4xun6
wa/2naO09oHhMJpTcbQ6Z859dzmYRPI7Ys2aEUttuojkJ/XGIALFeNp8NDtuqaDY
9A0u/hEvXwdUdsUzu7OV8MzX9HAGFyQ/k1ornbMSIlBuUTqEaxROxxsTc7kW92OM
IeMKTbNxjQ0mGRXAdFFvbf4dnOMN2brkYjiW1Hvc5Y+BAQ69JVAzq3GOGWZI0sQE
WfBZvBtdfY5vnqmt2rdSQluUyHSKulCgJDDcEb8Jlbzxgn6yr825mi7Wkals+YMl
5CfQLKtKmZD7XF6cJE/8Dv8h3GRk6I85XUNUPpagWM+hjNYA2cSHl+LsAxEpb1Bv
XvZSfdlIHe92OHzeylMit/gp9ix+ec1f8j0pb2Tg+UdbzEVIQ7EY8cBLQiQCWUMP
NnyRGsJP95bCfY3V15mgtC7G+oT7aQpdgTTIKwJK19u5YhgqZAaOeFjqzKRJvF4A
72GZqxLZJrCpc+KXF13TsCVBTuVCE/XcXy0kI/jeZnb4LVPZVQfeYdlM/Bi5q/Qq
gFZ+UQDTJSrlAUDszzJm2XPqxQ5BNWL6VpImX/0OCGQNh9OSbldBySWaOelu1/o8
vqJy5TmWZAQpJ4Qg06ED61tpdJWBdYcy86eZ62jqYAHWGMtVYSdJRrMAFWZqwmGp
s0hC+6fxELscMwmSlvH3PxZxmml8Dn42xQkC+q/01Pi41WnABgocdfUhXyX0hjbv
WjIWzo+KP3lHgf7idkUU3C9VcG7jPwJm7YVD1xVNa7X4Dtcb7tqX7SSaUe4pbQq1
iVCp/VAMjmAYG1temEZe933OlPAgnKNJJIwW5CLOHzwTSEzZ0rf3hyhKqIwAqY1U
i6g8t5wun8iy7377Ayagu/cMsTnx8QkmG9UB4oin1MaYSAdsrdN/MBxTiVn6+TtT
sdnpSr5CU4/5F8n3HiSMWEYiVDQCLbV9RbwnrXWvOIociQ9Jb7GLHtmAfqUQmQ0m
3RtHr50kpfuphthRBbAYsNBEnp7PiKH1SKTRmTg4z1P/euIbuqcQ1yCBCVQkRML9
vqjMpkuDi+JCH4fssg1b/u+/ivdSPTxSDMDh0iJV1o9Ti3mr03xpuiQEV9OSub1h
wHN8S8Xq/tPRLA0Wc4cINHzGdXXQCBvATtX7s+wF+nG222c+fwgHKK/Z6hSjoXzs
BnAz9/SxH8y7UJQdc86YvvigxiFHmhb/rrZ95m29OuqdWHQudIN6yygKDJgUzs3Y
0DfAseo/HjMcKN9dlCB8CvkUKX4kyH7+iYw7lUlQ0o/QZw9tuCZ35g6t45Prv6Im
QQfh8k4OiOi9R9f0KGlq1P9iN13h/LCaAjBh9fC9Hjifgw02O2olSW1vP7Re5tTp
whQjl89h5SUK9bmqeNromUefXdchAKn1dQzh4CGTlpCIrzHPPS5EA1hBc0Mesfg0
f5J8KAOSuuNoYsegSOF35VPejJJcChA8or3K2/PgmN59BXkaJwRkvKLGV+lZ4S3Y
bc9SDtCmDjMkK7zCrSKoLQ84ysRMUrY5RjlVf5zBhR9I51+KA9EGdMn01tRYlSrw
opuyxpzPOn6ZzTjt7TI6UbumRgHfsAmcul7w8QPKK4LST+Dk1CYX/5pGRQ/wbHZc
rvd1E6QxTtJpSEJJrU+Pa9HySrClBJO09PpXnXFo8SRd3zB1dm1BaryQOwvYxoRs
sKZWMM3vZw1QUBP5jmnSLNJzVG3r2U+cfZhrbxETZlhEAEUsygKzt7W774d4mL2x
g3d7XepCveew4pTcP8NOjAB7fzbOZ6SoCtDjnDn19qmA4MS65TgoIRVILCNwkIab
TMa2gYqwXzoe5fheyKTbc2Ya63zF6szFCjiTQLAHnU2BpBt4FWI+om6YvYENxk7/
NWDWEI1PvU06rEnjqqbTJyVsPvGED0IN0b+eiB1v695bJO0/o9x8pD48PAzW607H
89dc9YZ9RqXl6dvgHLBC29lzQTvFJH3p6h0nihINVjiBKaAQkt3c2T7M0KJkjBf5
BLEXHKzs6RWLHCpiy+rm6VvqGjLM+eiSZzUpY/4IRyajvMRU8PHWFYUZKiWtFCUE
HEA4cviekYPxg9Y20DUhBTlnwCWGCIYvBI1WJ96pQzCbXI4lHV7nWcYGsc26vHqk
FmdteSQYFl0s2CguwhkPlh2bM9UTXsASs4t0UV7Ln5aXVKQoRgZRGBcdXV4CTCfn
ip3aFZfcyWsf4mdBahvMXYXqAc0HcLWo7Zbi/BqD4LB+JbD3rASGa7I0zSPbR8B6
tvwCMN+DkVnRaCO92KTyUDGtpuxlHEXV4dckIqa4o14015oTyQe/KY7AToadw1mz
vUHclecdSjatz+f8iK3hSakaL0+3Jqz2tmrO2Q1KUC24Wj5arq4cl3Zb6uMg6BEA
941DX/zSDEk0Y+TO8PjAIMv/IhyQ2RFqgvz+7jd5lU1Qe1u6W6a6TdoRMwKtw9EG
zP5G0QkN7T8tDRkfRKqxhoTFbnq8IWWtI1INC/qXIZQJPxph3bLNFVNlnwkGpogo
z3EaJbV6lw6Suajno0OG2GUWeYAl3AMSMcCpbus6AAu9EODXZhFNlL3Z84HTkPAG
cGTQq3ecORA3QGtQQYXtda3RX9hdumrTaV4P5vbsST5Dt/E4AFltclZJQPO7T5/u
zfTQltB9PBaLvruPyzMMZY24qOlxbE7uti6mO9Mo7HtvdMGOqd7Yt+oD+DeFBM1P
UgQ2C50RwT1jt+8PN88WJA9Sg7zgqk89YXDleS5Re2WeYHcA9TAKUKiEqgv7oQY9
eh7PtEJRQ5+OaHEAldu9NTmauPsOSYox0OGprOZy0lpIJRwanS1mpZf0VECXooGH
cX60/Hz9JywIufrmbtQow3plV2XUZxqUflBu5cAxawa7wJCfwgwTxna/CwQKBpaX
qbs8T0lkopdQL3tKNu94mK6BL734S/qoE5fVzkReK8U8+5RV/b1swKQqq66tyEUe
6NGObI6osDxF4WSEfSexVKAknuDsSTfykjP18HD9jbPkuncCPBhbWDrmPYexSjPu
Iyan5/VSUmJ8SVpd7y89PRtU0jv7l7xzLisVlklZuB3yVARGJdbbyB/DFPZusx2L
+6o0G+qp2vhZS8TPZFCz4R6Wuj7Fl3gtjh73bmB14YHfZTGGHHhWxg5IXSTKr15L
PdtKuyfXEdDbnYkVYfgl9IGEUobtLl6Fm4VXXb/yS0PPJC3OEGx1dxFYnGETWTAF
7eqHeBY7/CgdUfIh/mjwsS1mg06jAMDTTiy82JmWiKz67KzhOO56ZqvsxL2ODshX
YUmMpauZkNyW79SaBBYCD6U45MW4IOEKvPqXyWo3+QvTN6xJ5K0d0CN29ZsvvLdQ
/v3evQaSvlzetyQtpHpwDDlHs9PWXIQ+BGGQJ+MPXIWwnrDbBni1VMbTbi8JQfJA
0ENFXZq9MIYvm4EtcJQaEyD7d0sHb35igoPVYUm+SLNxO0MSYfd4niVxTX2t74Td
XPDEmC/QRVerSlHgol/L+HrS19UhlvNJuGZMcNc3ahYH2QRI/cW0FbmrWemtYV0A
wHf+7yn8kd2RZdv6WPWCxlf8alWrgPPCvTTL93fF08NxCDwgnoAMd2ePHv72703b
KidFvZHEX/tw9C/IfWUWDOQsJy98f6a524MYhK3z/Bu3beQErS1I32+DPL8AHWn3
HvbB4ADZQvQS7gLbsYZL6AlI3yUOKBNIlV7G4BMWrqOZutbmA2t1E8YspQkv8chw
s+3pPFOS8gXFU3ZkpqzZH6ZEkfKeG6NDBz/J0gLoSoDXArom2CzGgTSo7hkh0fTs
NqeXXNJ7rbe78bCwefahkzoO5GQ7716jOwhHXV5DEQ/qkQHF116MnWhgOhgORYzI
k4SK4Np3FSv8aKeKB5ZxEmjLq26vKpdbsQEn57GznRo06rlkAF4ZwlVAQUZ26nNe
6zT0g15mdrnLBSxLI3IadPbFmG+Lr8ww9sBVnOGAOyfBUrI8hsPxm4qFaLjVptRd
TXsvpi3r4BXkigQwOiRvVA+wROklYm/72XFrUjieVj2H6J7wFJJ8l/Cj1CIqA89O
ZHwdZdJAnZLv8FpfIwDFqee4DIgKbOH34QeNAAnegd48KbJW4axdNsivm5LxSrLY
YCcQKUkvR2HP+ntGZgPV/yU6nvywGBxOCmDq4xgcOu0RGXyvj7Gfaq9Vw8xF6BEv
oED+Y6tEBhWnaxCQTH3xLqGOUGIXbm+KDwzGpU3B06Aa34zY55SDQCtC8gU9GqP9
zOqUVnjWEAm8XFAeQ1rICaWPphKSBlPYbXELVS6nc7UCOwDbokdejNB32iKfsewD
UlkYO+U87rYP+tLVhjy6HWKIKHd2/cvEAKUufeKYZFx1D3RqlcOB7Z/AE6PoF3M+
9BRwBZIaoN0G6ZGyvRZ/AvOVE1vfc0YYm7FYgj7UfuzXpVD8BTe1IAnVwVpu2H5S
JCSUPicYOvOdE/Fc5s6bzGglpsITBsq1s2SDFKlCwxlHzdG9SmC3JnXLXxQGl+4d
menvvn0+E85Slrto2x698AtvhsHxFqWoM7NnkJw0864oKL/b300f6+C5S7O2JYZm
RG+DehtRx2ccMOjPzP8+7fr+bkv4j48N5zxKVXZuVUhykt00l30HA5kzPhYSCPTA
yo/Ulzhde9cYeL2RAAO7oUK36bZlux7zHAccZ+/y5fU+V4UQrefTMBXrc8/cjy5y
XUN9cgx3XWxVxV/oWCVnWosiT3abkM3sKkzDRaRd3t5UMcs6PhBuA5DCZDNX0Drb
2T62XZdPHsGbXWlfXu5g16P1eUafZ4fzmXTgyOO/TcwbsDcvVR788jlnfw3cWd0W
z96Iz0Ykpr5Ukv7NAjxd+fepQUWoTE/v8GZz3upi0Ov4maoiJZCf6+KOy8fKy1/Y
dckU/WVtR++YsXFDNCrGPe/zsh/m4zdhePkKB/SU1P3McCcDR6WVN7WqQzd/OEmV
eFo2itufQZc7RqJlfF0FU9i/4nK1CAuyOAJeL6/lxczFFbFKTN9+rbTkfW/bQ1lI
erp9DVBl0iJVh/iI++Jf5d/dcKVssGKMdQNWd1yOPblTlKQhbvBLUVI3Fr+PChHu
3Ux4apRr6knoXqtIHmpuTi2Ot2xs+mbal0NltQday/jQdZJKnSMiJ3jmsISB6Miu
x80dsHnL1WykZvJoM5tb6i8Lx7Crs2JphnrfCkW9TVjvwIZ1ujqaJs/i0bwivZpA
UkucKXTPsEpFxq6d/gn4M6JpczmdOKb37sPHNPA9dqpBM9encQ7gIvYktJwhcbip
mraJpmpJxOSSbsOpy3TUvLsMebYnCU7ZOHvQZSdM/HjJDX9tSMAT5F2ZlFRqYghG
e+2+Xhpd7XFb+dB6Y//Ev5yYKUtG4nPYlAksyt662HgCZSVcRdsRmbONwQSzTUIR
kObgceZmB+guXEq9eZkt0V3cLwD3/QQD0WhD+7bckouBVaoQ9LMFr4Zjx2IqUxxY
KjoYJ1MstayO4stx11U7x3zvZz6GEVrsnEq0a/8XsNsl1b4RurCYNgwV6T92gM8N
4t6my91S98X9TLTejQ68FrI8CfNfWJyBy4eZ40NJqHwZGoym/fP81iq6WCTrnXkD
msRPqa8nLdOE3xCbDcO9YGp0dN+IWkLbpY013VvihoTUc4vPLazNOvkZ99kG/JyK
ARf/gES2ePTH3f0mEh0u02WIFi2zpXbhvN4U+I2xWLp9b9oN785/TULT5IWFjh71
RYxu7oF0THTz9G/SsroY9D30LHI4LVY5OT3nHhJIXcNfYAG77c7ZKBFcP379sNFU
9ZJWKoPqAo5AcOmol8xN2GU3ryVXaW2BL9iYcz1j/ZH0wPgMrm4S3QKEPQfeE8rd
iOXno9Ap2ShNbyS0xeQbUQSiK0UZ3NZRfbK8iNeYS1GyBzchTj8789INEUDgK7Zh
8W767WVxxsCnr7KDLmUJBJjRaPfF5O19m5k3it+TrGDXVAWwT17mw/IgVn6zu4Au
sGjqGqEWEwNoOETgMk+Y/HU6Du0b622ZOJR2z2S8cIG/n0YEOg772bSuzmvT3buO
9i3TOTfn67QumgDq6z3noCm75ha5EHxc5uYQ+BTzczr3iH5h0lhccBZnYmD7Iixw
uCNbiHA/g04ytJLBDOe1mTT1cng3bt8777Relgynmbf92T7HdzqlvFaxDRJjWgJ1
27RTr3D1fn9p8L4pceUTlvUziK3vtQmkmMGRUh1asjswQidunVM0AVdl0dYniMOM
uI/jLgSw9TkgNwFBwR2mkkXtyY/nv56jsls/XofDkZj6xGoFrelW6XaRd6qB2onx
2nsJtOhqfx7dPZ4nZjW9Ag5AnlLp/TqQzSn2V/tw51X91KvVdBZEJpJKvq9kxQWK
T50biRwswUeaJFc/SKggjnhj66xdXJ25Q02lZZCqHBfLaG4TeuhgQXXoozSrAZmD
CKSzMT2SIKYuoOuRcBD44UNHCGTeNOxksBQ9JJuaXHLXdMKTF4H9Jmesw0PmwSh6
8UCoHH2zApgHc9ZCHpewi3FFEV9xzQW+yloSHirxqMypfPiPBHHoGZkwzNUdJaQ6
P1WUZlsGpXxlczUZzQwdcn2JOhHskBersBv+rt9Q9kYw+BPy1Im70l2+kx784nJ7
vhj0bdT2Daoi1Ry8Cut6UxfrqdbYhWEoNsaoFxImjl6JyzkjQ24sSAELgMvI1NV9
bjAtnifnBYpxPvHs3WVLcLHoVjkRidYOiuIq29l5H3dQt+pTiK2SbSh5q/a3sNro
IKQaSXP+AO9FW3Q1ul/b7NTK9aft5haOoiOrdPmYL6Ek/MB/su1KIVsc6ed/IKlU
vmBsBgXI/BuOo14rj9PIF2az4Sfum/L2ekvvhdBo6WFQQzAfEZdL1D5uG+6TVXH9
PnZMrBWqGLrqLG5REFhzJChnWSbW0mSqX19zEAkQJv55RecWDFApjm5Mnpw/taEJ
2lzGLghsvLJy0n2F8a78PLKyxSZ51toxvyWU4n4G2kqXr73hEkZslEpAdXc43iPH
DuTrtepxia2rcqG4fPvQ/NOFPaII3nV7rDHknKmwBi0Oh7GorYYkWwg7+vUUPILo
d57LtLW+J9Ajfxy+kQZpyPVT6ugYILnfxKcBI345FNt5nOVWtRLN8AFgSWmGlQKG
VyXtaiRLiqKwABm33M8/57W+ktKREIVimNYARRVIzprkPNv1Pr1Tzy4904h8rsZA
mhUF7KI8dZh2rT2HUFTtA9NLR8KF6g/7F2Fbj0PAVCHKp0H6ZDPi4u/qx7iJMY41
DygOm10AVLhJ4Pc7KIv9H6xCPs0xsCSjWSsOCLJmzaBP3xZfLyGswlHhdtEkwU2W
vdnXD0tbdmGwXr+O2QGHiVSv2YJh679juE9pd+7Ty5Na3TklQKdgD5XfQPvD8Mux
j2HDsq5NNsZVz1We4qKJuePjFesDyR/+RqAbuzg84jQbcpMfhzzWiAiWsE6bXWXJ
4FqPVEBnOn9k8mDJLmEohrLlfLKjw9AWV4B1zE0jDi35fw/vCd/67e/9QJFx5I8O
sevXL0DjXMw8rTEQDFZ7oMb3ylYENELl62/HwOTRTtw8DpP2inBsZN/Q7+E1olLd
ba3jr6q5idtGNj2MwjOGQaeFVNlkM/TlguXEBhDNYivPNtgIZLkb2HLm7nC4ziRC
jP6ghf98a1LAzNKPpVjoywwwNd7bniWCd8nV9/Xqf3qhVn5BcoO7XblujvUeY223
RwvtqoFnA6o3wZlKxKz8vCwWgsPy4r+6PoTmysyiCZ7Vccwy36hAIO//fjiJpjwF
P12Vv8keugZzjHjjwlVN8V97XO7KfeNFj8Mfku+QmUJ+79pHPGGZzTidqziyAj1j
CczDhIh233nGB4ia1fkSGWf4gCyzKETYFewLgRmQUP4newx4Zi0+RcwKkCm7blzQ
lnDwMFALWsSkp/W6ljTJKqv6zjNQyOij3bzhjcKCpc1M9KLc/8NTntBN83IlZYid
r0cgNxjdli2PF72Ldqatm6aYF9jpj4wZp14gClLYZyeVho/Y5L1GVKIwcSTpFbyB
fITBrgCn+vAXnQ+49G2W7EjdiHb38OZ5cr5dAn7ua6ZlJ31IRc5qWViKTNRJd9c/
ONDpCI9O6WBdJ23FJiNg0s8V3kMaDwosNNm+064oAYmH4O+7E2644qrFYO97IXC9
+z+TdLX06sikm22DkQ6SNq71VSeRmZV3JOWyZJcs0RTzzHbb8ZqETJ4iHBZLocif
MtlPSlrOFFcYb7amsqgP6lzyybhwnp7juNofJDA85EBjWifPxWK2SDvxjx9wZKID
f5gd+rmTkPLSYKu6VYmerBi0FMHChHH8kpPSE567uSpsrRMrzT3ynz12OGrZ0ph2
1hmO3xGdMvTgelv1wC03QGpTr4O6qY1YcI5k84TDCBOJnq2hB3EXxKwF85yDhyAz
mQNZxRP3RBu1H9xB0uVjtRh1ZykyrgyVYmB4Xkm12DF1Zw0jrJL9RAGZSPHaNtWH
67xC3NFTdFD/HBs0TtMF1oF5h78DEn5ANr1I2521mdHpS45x7ArDAi9ne0IwcVb8
veGF9ac9UH58olOJUa31mOPVuxu+QJ0XDya3T8qLiHdePvT7HRQR0D59tRN8nsUo
HiisKYYdqWKcJaFMkdzcLk8SPsZNKsobEgpzCMDqV3Fom1CQ3xI509EMhvNWulWi
HDtcRsiJZIYW3DKctO2iy2CEbHOEYy91hRxsUe1H1/RP46pSygmsBsOMpGyO9ehv
CHlhFVLYEYeShkcxfxWQgtkVX+KOmVLm4gQSLPSbX5z6G2EGD9Fwvx1Q3fOuaV9E
U6jwiHugbXbC87J2pthVO8cMjz0Lv6M8aQ1dLywwqOtfAfgmcIDfYdDQaqzcPCLg
6pkSC9aDOw1ldHf8KsSS9VTolWFzzM8ksZ3hVxuE3nd8K1ZLG0nmplibDCEbEqyW
zXTBP6I9XKWetrQ2yBzvlueX4t0RWfWVUHUtorRLxG5QjhXoCuWmebyNa2g57mBd
PCdW4/nQT9mcDmLLZOGqF9wW054GH2UgrGhxyTTLZKe7xLLyEWGGd8gg3EQ+NfL7
kFNhHcALcMksgS+gC0+zesHSf+L66jPPII8SN2BIs3f8cl78HV2cmLYMEOnEBijK
M6er/LutIXgpF/MDkdK/TBv0YzgZpGVSLP8Q91TTogi6tvdRvqR4HmCYl9SnaodR
+OGqQuU1n8PMIu4V+SkpUIdRoS+QOjHuK4KBzbl79gVLfJ/1pBzX44uewWYjvFih
uQLP/YKIXHuR8o0qNlGjV2wOEeepDAJJgykKg/5T4iPUAaQdC+1vItXuCq/yxaKR
Yvoexb5+Hwx6VCScZrtOlFPgRefhn7yLWViJf8/OTcChhM1HnDP90f5YXZsNwyOg
WOICFvrrJ8YS4y5Pw7FKIY//YdbXHqlZ/7BsYBIEwQ6gu3svd2mlPbOI0JsfFaqO
hR2A50PVlYSnVsWLXb7Q4n/wJjku/gfMjjJoSPRebhm8eA7aU3YoONg1/fig808x
vJQ6TbwXR2SPldiT7i7AEpWBBCfBzZtmLrHRP/GEAK+53jGFJfNxMliNtnfI6u+U
aB18kYc47sDRv7gX9Ki+PiRKh9/1J9hu7IVMNvsdZ2ldVB1hP1KGLjWvXdElRvju
foX6X5THBysYIOk+8n2/cR4o+XfMOGXNOFYF/vCJhPSZGe3RZ60q7T65Omxhfsz+
SxcwO8uE3ZsZBGG+UNibTEmAXTsAlaiJbcIzBvz2Dseeb2DPE4Yrd/9IJUSW368S
9S2Zf0ddybaw6mHs8L/pcpkhVEsnMjC3iMVYb3tOesb0qt4dJ75hjtMmzIAMqhe+
IgA6+N4mqiGhGI7ZNMxNq0VmoIdoyefh6bx6HB8xp9t5pRGyMt7jCp6HFE1DOOZo
81C09/zJsxWKbO82z3/yjTkcS5xnIOPtdZ5b6geBfTPEZC0VTGLYvbvClthsTvbj
etM9HXwWivBJ/CMYJ9sk5SFoJTwvaHYYQThITGTxkQcg8raoKY3bkSCv2fgIljXB
qa/RciHHHfjoNkW/xsOaQOlBUMN+eozH07uk0EPzUdgCcLodoBPalv4ajYQg3cZd
RjepdbHkVNOc8SfjoUEDXmABSa0qgU32j49AiCg50KccA/7u2CjtQ7uJ+NqciHzu
3J+hw0W4wMrjfMGnJjMErfxHhGjjUJqvi6O7y4b13yF3JmHrB3a0L7DxcXx3E1+s
nIZ9XrRvBnvlDiQV7e9zlduwBuBTBuKKWbj2x74khDMQdQf3AS/8Kcg5WBRtMdPb
kwB4gIiRDagClzKpuR+esGWWDRYRG8yJTrK4gBGRvxspzL5AuRYZue9OqIjGTTZi
iUVq2yoAsH9R9FHTuxWCk6nfibBdOdWm5NNuF+b/2EKbGF4A/i/gU+nQ3Nyg/9K4
aGEV0APxByqwfwX52wqiCGySecWqMjQTU9Ki1IARr/Q0kyLRceOMvxHKsFVNM+2e
2dFP7XRcDnuwnsfw3DOWiU4hnMky/GCd82/is+VSY+VDKtniJ1L6DhjFc3dDE00l
LLnoyQRbT119fSS9pWPcY3M6PNvYKaBCskp8DOudrE2WvMkt5D9l3oIipExgXJAM
VHSbVwwUYZLTlpRx45feafKog3ZPIeTIBToTYxKO43SMR57djoOB4muYLpENdZSo
7c+0GOYqYIa8YX1tEwhi/vvSgrelfNkPDz1SHWx9l6cFMiz6Pq5hGPOvuVctG+ie
wMZmBSROmbUgySIiglSFxM8EGD7o5jZBNcIksyR+MpaWBdLT5R8F69s7kQEUADfl
Q0q/kBjEmgghe71TgbFG7ZtI7N/icygWJXo+l0/NdnIErcjHXdZVaIgcohbm6MxV
qZ/3OdUoC/4C3avOwescamsq/i7xHxo/dsZ7rEMTb0g8n1yCJZE8CZDD1XOfnaIF
pqYMMUhpQ9z4pIhEDlvMwodOm5+elKf7YRsFkU6Uq3VDSxBHehbvqhFqFtuZiTQm
z8QEKU5xCYwK5BoJCxEvzRLcSc8dD4PEIlNFn1Uhi25Xs7RZjdvk0duZkayjgFoG
NZy3fB3GixDxGaYg5tL6nLCXo8fxZxU+pE3gCBF93T6ujjrS56zwyWyEFphIT7Rm
gSGNftTRRqJZA9usEMdaoxDMb3uEqNEgztb4OcFpPXCKhssSZpNFMb0RN3oc2N+l
BncLWDiOiAN1bbMeb4oZzTQvoi7bwkg9xRvYn+Vey0QzxQ9Olp7epmrTzyx4WjQY
u66fvXTekTb2l9OojAtGG7rq5LQT9AehAT/73YP0fXR1GzsgYaq0vrdGdnaWllCj
MIx3ymsO7LQpyqEvMIhOxgnNHcc+/i6scWznQGq5VmH/nVECy1vYEU+kU83p+DUt
1YexEtcgW3XzBunVoNk4ZnpRWSzUssV35WIOsp0gz5DU/D/eSq1C6WwHkQhT2OEh
qDI8cccn0ACMqztQL43RdoogNrDCs1VeYIfs8wYSp/ffsYeb9xdrwWrjHvelrIIe
uDxE5iqoZOLC09XtEGhpAhhH3ruqIqGwlKiolDQaEITpzNyC9yV2YBwF/f3tXPfa
G3dhe930n5j/asiimq2eDpzwgHCl9X/RGmgY/9G1/5XeLo+so2GeZvfKTqNeSumA
4onWdP6oOzma1pshWg5NOt5uvL//XlJxgzXRRRwpYsjmJK5nkGRGhMIt3IhvGAPp
XezIR5cg1vtGaJCeeWnzyRy1nyaL+TBjSzWQ2lHFt41tBF+OCmtJAwv1RcXq/6y9
i18B4y2wA1d7RGouH8c+hoYepo8T7Vx8+ndY6wdD1YrTQ+DP7i3VtlUumBsXWE0z
EPvH7YesZo6iSUjvNRdOM2Oh2RMICrRoxAolE7q1rBnfJiaRSVBK6p+TEmCGpZH7
dimxJ9DgltLx1uXC1aucbQxPE9QpAWyaBOY8yVf96K4pNGyYH4f9nsquzz0EAACM
dxKUYD5RFv5eSVsougcfnIrOT7trXggeum6wSagaaZ8tepN1jD3SS0fxkpwvL3bE
z37tsETwWIZs65iJ+ZEpN5tBk7l1DWiMZf/xRazAH/9YsS7mB3dhUc7qSVAKy87+
QkTjDi6xguXkwhwHBNhQkjv8zvicpbB/bhTHGVGGcjJJ4v341BgmZbb5SLv1jq/D
3YbmuSOPewg5VVCPpHxT6olRJB/ayT9yHVyklt12yxtzXu7pAz/7o4oXeEFu5M+s
vja2sWpFkLQEw/mpB2TCpyl0GXRWeDavN+3iATd+CSITfbtSHqCqvap0MfEHYu/g
uIHd27TkafqgJt6ASka/4dagZFpk81n7yM0hetHaCKTtOyDLAwizyMegjcEXGMDm
aOWwK19yYRy1l70gjWjNrvYi4fzubRh6EMwYZnok8Yl+Du/gSQF0Xt88cjsK2B2W
AehyFcNyLkRdfaRxcndk4PYEb4Zvhz4xEeYx/VSMHXwuMi7MP06qmgLywPTHqw/c
nHVc0vv7aMjGYpPhJbK8Sd4Pzw4s6bU/VjWXmS1ty7iD5WOfEo9+YjHA8RpfVlJR
IiOCl73BhN0hSX+iPX/q/LgczexHC3p0oD00Wgzy9Q8OG/0HhioYGNAsiHmC5j95
aGk/7oCdMizOL2buCOP/yVY0RlYJjSuU3kBpnXLqa+IjP3tidzzRj8s37TWu9sVL
m6TQoYgjqPcW4rj+qWjQ5GXq74DljHaOlcYbaG0MIn4ZN5cG8x58P+0PVmxx6Iaa
kCU9aM0eexO69Fd2UVChorAjkCw7Pf8MjeLkE6QnRO7a4UUZjerVtUxTX9khnKl/
ZFuc811GFkEJTCPlNsJdfmkVE0VlsdsTS4164XaSbSg9i1u5dgAzQRUp64tRa5J7
9PL/8izXIOYgiS0mOyUHaCY7x8TukRaGwFdQVki1ECeMjIHlqsiozqNTQG8fuuwz
+9CuSfTz3OFr4550e+Slmihzmgx5BQMwyf8Lr9zVjy6s1m6+75R43Dr9A/5vL6OD
d8oDvdc2QAKDK3RpZzooXZw6oeBKRPi0nyNo6AgzJMqnwndV4CfRHlMvzJF0m+9P
LhlpsoS7lQNh0fRiiAewzJIlHkAdp0lhBRyohdwr8PIrtnLC8qixswFKTwh40keg
t5ZA3KfNNtHIPDn2qYUC2g/DSnTzvSsK9pmXqB+sd3u1mnrVS85In4Zxz0tOfy6V
6pX4rF9pBr2fA0IxptLE2x/UP+5JkuaZQ5geHp3HDJzTw2Iq5tn4qkgwuBs2AEaA
ysqE/BzAZn+GPqF8UmEMjisHdiJtWBNbLLzVb1jIf+56C6MsHhZL1K+s+jKYHjd5
PbWRSTgDzGBVtFTE8hTS6znaDrQywR6u8c0i0nbJvkX2WJeMugaWgxnWU/uoqwLC
cwuHLDMzFpKzjLa9ICGXNXkuT+44tjg/bjj9rm4ttxUFcvB3vt/bwewoITy6h3ZD
bNtT1WaNkRXLhMWmemH0yCwROSzFhNyUtdMqwHOWHd1yiEQRVmUm+X2z3kmAEr2u
SoZFfxB3ef8VXfxmyWFW95Cbo5U+y45dRi8lSL2WFzyy07LLF0wEBeeV9ZjS3/r5
Y30NglFbX9J81olHY2e9/L7Kg5Q7JF9WmT56QVoMC8Za1ptkOytbHND0VGhNE7w+
Z18j9lNj7qB3l5RTL4HpRY8fkAcprza/VRCl87gaEMApFESF4bcETmqbQnopHkoH
M9Tzx37cGj4D4OJGUP/C/nfZIJrF2GyQedEdC6GLJoTN1Egdyo+z2nBb5LCldXy0
TMQt8pqpWKOBGMvzx84ZfxdXpNbr2xQ1kP+gIkwIIll2wmbxSa512YRRRXEkoGH2
TBAoTtqOypp68s7b5z9SYIGwDZG4zKFpVmVoOpCWDgQkFsKA0lShf8myR5UGSGNH
WLKNXDaoEyNdZ/APnS0JRtvfoT0SWQpO4OfLpPe/heeXcDyagNu3zoTzo/XQdk+f
GY1q/H/sTytU6U8h8Qn9fpgljn7rOpnhqvvD3NayDo8BgDCJlW3l+dr2Jo2eIkda
ox1ZJH8gG8jXgdXPwLUswJlV5Wixoo6MpjtvbPbgPHy0xlEY5RXOlBZNgSRu+Tcj
+E0M0otWTAbUxZiANlU5FOXYaFSYhk6JDxCyesni10nN2JgfSeoAYS7Hqq9/Zyz8
3Bcj1556w32OAa8cW51HjXB4VemjHX21bBbe7z++K0J14m5JZWMWbmpJVv9RLzmX
uIZ6X0NgMNPwShBg1bvZ+ks4FIT6r1A7wKxsMJHetldnHpyGAZvfxtaoA0t75eBd
yrOetLDiFc31Z37tsfY1d/m0A+DZnu+A+psoZX74iy9udHuZPtN9Kmj1XBbjx7mz
C+eErE3iPi4T5CTz6gyAASAe6lzqCJBnckgQiAf+u+Fl+bBQuQlwmMof3hITAdAy
uOGZeTBk2qL3Fs9q8SbRrP3ONvpVr9Y5ZBPFAvWACo13CcXN5n6iGNT0G+GvaLnf
5h2rUSX+mdBoqjF6oBtyLUsVkka4MHHf+ND1MMJESmd1x5LlSMzazXIER45AAW6H
c8qdh3Z0BSsKdNMdSAaGuEw9b/n60puCnQqkMimA2/T3GPV/1Hxn3COV4uG9jxRg
H0ySkMTTXQ8yAf4QKWNN+pxnV5YnZH5BikPOiCoi1jBCH99yeS9svucstdsymBf2
34HvOPlUPb1vf10/6ziixggmgp4aZ+LR9VOoc9Wpa5WRCzpCP7/dGXaq5ZASzDL6
SzIXHZYeGePTKzGgZ2ZWQI3NqthOnZaFuOb5oq4lUJhEfy4h42ugO/NyCNfl7cgt
kEE9R0yvoxps+gDQkegCiHuvm+aHKr1tYUexVNMwK87hx1o20ussPkhjgBDIFbju
pUV2PhftKy4aL0V6E17JsrcEGDmQOetynG8tzNR1fcehVRiNNnU0JVy5HAFZl7pG
wtLWCBN4CYNzb66f4nnP4eKnBtabU+bDoomOSixAi7kXFWw05gcQ0XBwj2CG2T/h
eZP/oCXZfKeZfRiQusBV28kdSDLjCGT0NRrb0i9fpbrxyoXbmqSVmSp2Kz4OD0XK
RgdVrDLtzfhHhaizgyTsaO2SDp5YvRM0VRAuUCENWqWvxOwry/CHBAHZ5XNMUAgH
vkvWIz3KnRmkJA3cCGFTMOwlR45QzlDXRAnp5Kg3D5slE8uTdP3TuGzWkcxLJfHb
yPOuVHQp/2e9hL8mP7E7BbpB3cjGPhkUgMtaJPEU2dsSUu0YhY8LnEisMXnyaNDH
xxZ1nbIEXAwAk6Eq8vKJTCWpEOZ+IBzd0KHoqInMKnDbHyBkfpgTIIO83z+Xsisw
9WagWDt4T59W5dCfljEw2NM9VYD9jd1pObAtBr1FT58xGhMG+NCDv8VMwpCge0Af
BBlXnZehbYxziIqgQixcEbU/S7L6VahLyOlICBeogU+qwi6Fd142EftntIiT9Wsj
VHVlQhnxtXUOGZDif4kM7x9R87gVcuZhFDqNsDS8+svCcfrRdyDmXqsQ+uuXBvib
0pK+1rxA47fzrr4AjFpbI73xMpCWHE58VFl5epAn17L/ko43QluQlr+uT7ZmLZwR
xCj9NLPrxOp2E1q44xgBcp2tUm/Lp2v6i5w/KBYJdHeVscTsmJIN5lsjbvsLNRBX
jiOUtjOonwMVZ2qTCUo3v/fMUje64ipZysU2PyXZtKfGOXsag82q1izcxBGuDkZV
u3Zq3DvKp3RCCZ7/PmGKGpWHKldHkjbnXmynyYbhLHv3tTtX636fdRpehUPAb7qz
ruO3+Or+ko22XT0Tv0vjoF4pu4yHnmoYzdzjYnPuwwh2FdTkInD3D5hhG2h1XvWw
aNcAL5nDXq3un4oeU6I9084rNaZh7H7Au9KY84nYvmUZAOZ5GXHIsTI1lBL/BfbU
qNP3Z3JpfGpXHTw+WhtainjmkwGCLaVBk+TsytiV4LweypKdO1ZMcOSjurPnDUHV
q6CFvhe4q6O1tWIkx/Rf5/AB8ZR3sFB0xvOUhodjRYeVtS+vshFxwN88v5xXwxFa
KY24fmjQAlKINgGv4L3PzGvuCIZXgRGlaNySM+fNdQqgFVugrVontnw3QulVTvnO
uB/jBRE9j+lzfUlsHc+qFw1yYNQeD3EM8gY4OxgjCPSN6cNTOzzqzrXVPDVzFO4M
gcklEAx7S7ExBLWuvwBwF2y8dnBCjveDqwkQHVY3+hvPG+y1Bv6ow2w8chI8kgCu
k8oyd1MS8lY1UyfnkT8BwkjsVWn2Bk+encsJfiEqoYvnOE2qzBGFytLooqSx7AYu
prAhUHAxx8S/yqaFWCNrPHPDVBlFl7dbgjLRYU21ZWpUKg4ytnh1EPLO1rFZ0aBc
dc09mId1lQjQpA0eufAsU1uFeKw77fuBSsCsnWH9OSR05K0KIwacoihDSqt3kky9
CuD3tdvRMehZnRZWmyibxMCoyPcRd1mPgPenuFSr/pgFolacabdtvbhZTc5icdJk
Z6GLt5spBSyb3O1qmlzm188Xv9qHkg/YvgjzdqsbFYLfxPt/sNdicauWupFmrM2y
CUmE5i/f8eGxdOKcodtnuw+GwLK99wyoTm5KHiMRnuNE9lHdDEWcmeaVNymgMdmF
wq5ebETXenhTkoC5xN5BEaT9A6k7wrTI9vqrUK/b6YfLoimnEORiyTks2S3FAQke
KWpOmQFOgsyivH6A3Ac0byjFmDIazzc9a6hTNa6VIZ54g77KbYB0fxIQkwKv+aF9
Vpt8GEE+/Yt96hMRMyUhHlyVUZiRjrzKh6eOGd1HIZP85Uh+oHnQZ8AGAuixwUcw
SgnuGPkiVRUWEi4o/2+3sczTTO9efPjkIMQdbb+3zjLnAm0Nuq+2PtpbMpuLGIzz
j/C5Nn2OrhXt1IR0A4VG1Ya8lUUtHhbXwxeanIEAm6dwpMsIU3Q8CnjsFsWxVuFf
z7BI4rWCEJie67pKHKZAx2QhzxYn8DP6i8Pd4kUaEYk2dS5cDgVAcKlfIB4vKG+z
6EwQCxMn3jTLZVdixSS+TrH5P81nOcDWiYhDcwXcrVeFe66HknX2LBjH3/k1lyjh
GF4q5j2QIJP0NlOFJ3B7jchKt22wsGPDdkYuJuoH+2i2y3HmGiguXK3VCl2+Qi23
SDdF4K5wTB1hwDamGHuu/C8y6h3NajvUob+GiXbFob0vF6xXnB7RpFsXD6j0VH6j
mWR6IPp1HGyRGMc1Ce0o4qxjpylaXmwZ7XigDvvZ7dWOpwJOqI0xz9RE57g6eIBn
kp13QWVjoLP8EteRHU41N5vyBzY36Sl66o87E3Z1ie/Ql2UPEBpziqnpd3hrcBTz
PP1XEwY4Di49kulFNLIZ7PjAAUqktgA/U8mpryiyoEQme28c9qTuqlse9NMoBRHT
e5CTnrBRttguyy14TRwujwyhiuNY2puPkEhFdTzlubwvBMRj/WDNhDUcY9tdOzoQ
eGvzW93I/f8ZQ8CONDkOp/CA9gcKk46+dYVcpUGg+rX2VgpAIgiC9xhS09olFcXV
glOas53h6mmIVqTr/giNmSRUw8NHibJBmxdUEKdevKPUmVXF1hSiNBtoWsTLsASL
V2E+UybaT0z0ISz/8TqBiCQ0X1sfcJ26++pIsaDOTCU3FOfC0in+ERgk6/LXSTws
qaEvpgd1WCudSSDDoNjG0iKkCt5BGRfr7IvOdfkN8nea/YCPNW2M6eMKvTUvoFDH
PqoSEKMcxTk/b6jL44EGePk8SnEII7Vhr2PM3y2Xz/IvC4pHd6mvRTrC3p1OG6ch
DqxYHTlMjaTlGOUkHJmShEmYVSoB5MJKs8ofCRYB6QTdEZOvJ54v2IZJqn3BzbUj
Yj3D0BLXnpeZ2+JJhN1UAmr0J4kfeNrFrtL+44HOYYfC7nPsTE8CXNee+tprNqo1
tt9N7ivMuuI/hrVVgm/I6ELFRorNBkFiforqFOrbfWTVuR6YUUEkvgqDsZ6/owVr
miSUuJHEYSKmNPBfI7mIQZ/KXVnJuk5vwstkeMW2G5SUlS6wg4/aA+RiCaUZzCfG
dHplA4YFuHq92JmSVvMnIBJEU7HLloszLZAP2KRuM2+7Zk0vshGObLLcgRQwAC3o
kucsUIBC7be03QLzUSepZeTvpQ4yHC/cshqsAo00SOfoEEsEeRoK44g/WIyIFZKh
Q5kYHKzUmuhbI2LGMOgZ+w/O39D4/o83A6IAtADoCHMWWo2v9/E4Goeytytzm6Lo
1LILRC0CoFIAC1C9AGDbBo1KbvWwx/QvWLyOU/KAvTTREIyVVE2DNeMXumNQs1T4
qJCm9ALWKSsmWVjZpjUoVIz1lGuVlZpuw3y3D5ihRlhez8dpkbkQ2jHJDucM+MGN
wFqKRmOGgYzwhRZ3DbeG+FQPdZVS2+XOQI8WPZkZED9NlLbfU8xC1re7ZNNLiP0r
YZ84h/mNMo+E3DoEqpIJ3IoF62kPTZw25VB4/nQSety7KUlcjIiMMDoh7YO7zzLQ
SSeZTnDVFt5ojdevx9AnVS866WuosUnzwAGH0eR8x2qb4lRSi2W6CBvG/dJHiAtg
FZOMfta6OHYxEu+JCADZQ7eFtxvy1kcbyjPQ5dsnVNhiGEoJuH/NZkSrnAOwmFz/
1gJgcbFvhLquTdGaablTLryUrBoreNpAcDwuixsXA8vdZZr+hIWuzzaVyiLEApnD
V+8otNyHUM0niisIMGRFwSgy+OtHNEbDBli7XkHqkweJtTsxOdkmNRNAFEYZ6MNs
OYalFsfRVqr/UPcyyV+tHwayBY8FdJve+SL/tZ9ApzzmSqFdY3aGa3TqCqhLA5bJ
fj0fBg0d08DfjghgUstFXKMRoYQg1QrBQV4F9HWS2tSx7QZ/qH4EOOS9Ezp3H2sM
sgInrnYn+tjvxpjFJiu/0pzrc1hY7ZdLFMGNOJUDV/vpqLJmoXAYy7oGqj+LsPK7
p1K5jWbU/S8ofWFCDZK3XoGZUti+YibGGXXneMeeOdG9x18ggRVz/y1vOsF2FwxN
/Oa2x/en28VNFWg+VOHh3sqsOn4skCRD0XshRaEFyeZ70Y2sZLUbHzTawdSpG3ME
k430+7zOZFLD87wjMm8K2wmSKiE1V1Y6UUBDssVgy8/z60ZCz91/Jr1OCaRSgxJg
SQmR18I5yqvGzuAr/XJfTpaBZaxl+gJPZ39GU+9fOBvBYXRBh/NvPI13KsD3gvu7
K0t6PQdJh7Xf8gpj9SPnh5Kc1E2tucteALI5gZ7BjFsoSizb0BEeiOTFKTo9I7lT
2TVg7FooE4Ag///p2khKOHzHEsLlu2yqTwBhllY1WxNh8Q86utPTcOLMvXuGEejP
OmooMwr431YDLPEtSo9qkqwngukTmquT+NahUaOU3BEaLcONZyrBa2m84zsGALSP
WD+WJ18HsBTJh+LVt2F4JrmdwJI+VDin91hTD2N7JEzOPZmO4JdfhjlFNzC048KQ
6r5AqnYGyxTylZ2yyRtaY4KXJMviSmXlDph6PvbJqDqnF671ErXprpWxiO/J6wZ2
ybUF6wPW2hYPond0nvxHEbT0lkfaPW/Uk+/nURAHmf3pdrDhv8HZbOrQYR7hVook
ss72UhhH/wbqKVTKCoULsGalVz9hNt7zzaJrEa3FA5S76Pg8P/yWimY+nhjPUagE
qis6Qq5mY84NxFB5eMvdlzlVSKizr4GaPLuujvbD6MJ5Zqp7+aiEFVqLMQtluDZi
WIxbr2LpQe+si6EmlNJ/6x0syYXXl/8lV28//KbjYInj5mlSO3eSCnWXrIjFuIk+
zLazCgX8Uo6/qWUiQk7/OItW1lDp8n1fF3nude79cKMtQCapGFnTAknihweUJWt4
TuwZ66GwTvRVhHXOFz1YGUY7wgwipVHO7dRKVziuzqRZq0pmGOPpVhECYPnbXt1L
XuyWaLVc4h9X5911M8e8QMa5BMZGux4rOgPaKC5hLdN2TUQAkErnaWazryd2LhXs
q6lzwMvHgKIpBw3V/3ZxFvkebkl9BIiYjA5/T+XtTiTWwuhQeWj61ZwCs+MNcXe+
Kls55TKWRdreYNlESCP9U4pV55QeCZgx+Lgvs1hMdZP7/QGRvn2qowv112TU9+Ew
0hrruZm2iQgRuu5wPkUrAdhgqSO9/vXDGo5HgLRE1ItmFEeZKJmHqIi2kpq8xyJw
CPacZ5tL9SzdgLhOt5GovShEqtJJ+ukO+F7IR3Hh0nrb6xq1uXp6dZuY3dVGogDQ
3AelFzypCa5MYxOJ2g7PVD+jkuMR/k3cACM9ey6VvbHDpVZNFAhcCNZIM/0lE3Lj
09Tjy6gZqhx6z5sj2xJcfECtOIP9b6zvx0oWd0qhdwuPSH55S+sUttcy05SB6j6s
QiRNrpeyjrq7drWygvjzoTnC3R7O6nvCsJ4uVYTy6wSW+uv8V2zMqAXLgQpBvNp5
RDNMDzzaIGySzRfcp13sTMhCXKUC0q9uRGPAESwi8sjfFtIC2R0nTlDpAW1k6LoD
gy+iyqyZ6N4gWOr3Fn+xQ5IqNQjhVdtJqqiahcLV+GVwCZ2r+8LlOd1Z7Spnqorg
VCC/gZjVHmvQr97Rnb5KcIGMsICudfOx0lZXiwZFQ0jQTDTGK1VURnXxm5bWPKur
hYmXKEmXaeHDofrojjWHa8VGk0uD3xLtTXU/FXcGjbNxrFb/GNfGfsBOEVmH3lpQ
B67q2AyJ7+8Y//z0rM4bnREFOWXYfz/HlU0lW8vhfxznSf8a/E+sknZoCuYwQQzq
1rxn9Ifk6kX7em4FIvTCsbmZQiJ+icIWS1AvbFHFxs1sUStFQyaSXxxodRAf/4ut
NTiLFJ7KftmzMy7wKUjHnu5/hHj9VumpHwq3A5pjZoPmHrAMZwGET6AmDocQaZek
kR7wbvkgGvl5sWowgrF66yyOSKOyBIrkouF5ngoLDMhU9lpIdIgGU4od4binpKir
NRDM2QcLXfxg9hmtBHA67ekmhK41+l85myJ1VwwxncimoEBzmx6CYrLaDd+plaom
VcY5uYi1ZKUy5Scgt2+wUL75PvqDSQfs9Yv209eJU3BRUvPJ0i31zBqeBcOyCCqA
QcHuSFVuowh6aasDAL04npgd3R/jaG+HQJXjqTHWBm6qeO+VHpS3qrn8/zLmu20d
XLGsA8GTf17UrbcPbV9zJRJHwhS9/FOcRjvbywhAuKGpGz/VuoXdpPyjOit4lHuG
mjR48i6boz/rYJsSf8h+MWVdTN7t8ZQQXDIi2WwpO+26+K9rheyBLY1DelxeEonr
SVHSnUP3Gu8sPCzj64QyGwVGIthREDlIAS05cAwU2q5slmi3uC7/Wasqd+j9KnJl
DF6XxY7BGlUl+yFSG+pzzaPQLkyPqfadd2c+q377QEK8f4Dxf5ia9W7kjkeWF4lR
h8j/6zTtpHcmqV/6Ravln+TPaIqOPh5KxrLY5XQ66dLyp93de2sAcgsP7aM2EOiJ
AZxlQ78ynlPvqJ5qUlctPRr5rX/08fq4hl9nmsHvb2o8P9y0FL8GPKOY2wz582+h
aewgriT4paLiLAbgu62KAwyCTKHQ8Lvwy785CzIL9R9bQuv+g6KiqPRb/dHEo490
4ODnKHiG1MiUSt8tXZCjiAak0Ksy478AqND9B4XZYK+KgThB7tsgwZqseZ0VEXPR
byv2E70RJueroQbVp+pG2/TblTBk4HZe/zm4xffcuCTfoH/YCwakECY140px+Kp/
mNob51j81uhRMtuZnYu7CtBfcOd2jhN0JUuVMrcrl58h19NpraRbghYPKC4I32yP
+XiOfyHUIbkLwH25rQRbiQq4yp3K0oXyDaLj78RsGA4yOe9F2lozsTzogHVqU5Xs
xGQWaM1DruJr/4F29JzOC6a7+lG8aqj+ZaJv2hw6h4skBBtZS1hyWwLzW7taGDJD
V3a7Y7k5eNVqaFG5dc04M1FZHntlOlTDYo7+1u3tNJp1r1SLQvYvEXlYgJHD8PtQ
+Jc/l3OFymoY1IT2IImDbksROqqOYwk8CFKLO3g3Myq88V2E9ssFIxes8gMEtRVU
EdxpjN/nlnddy1/sMWc2LTp2xgt1g6/2PMc1WxFikBzu/FOVCtFa7EydZLXyu8LL
C+ZMD3++xnH9SFK28NbsemEVIytVmJdMJsfthgYwBQtOELUyn36Ickg9GMAS+l1E
fkws6Yzh7JtJzqjX7FisGZ/S5Hwo4O2/qQHAqchZy45MlxoERFTl6h8oj6Vma28g
I0Y1AhGAy2/81PD/ia5f1ZObS8YB3hZbBw2aFWnoZh4znz2Y8jXufCj+W+WQXs1B
Lqsp16ea2OarkZc06oi4Qcs04PHDfFlkoaBEn3D1Awcx5duDiH2rvgkwuaCzc6nI
Wx5B5AlhKhhZY0gbBodI1RBY1XYVI0STJSTDz73Eot3SEwFHctuXNRa837MJm0iM
i4AUKk0tQ8A47qjpnU0LugMNiWb/371T+9iGXpe4StCzlQwF8LSnMJUaNoAB+5xy
Pzsh51eKuAvBBv4YfnSTbfdCPc6vAaBoOcjrj7XExtnPRKYJIca+J1OuEX+gY/Rq
bdH9gZZNyxqOC097QlkTZj9Q8Bv6YyDCQyp0FLy34bxG10IagDxOVh4SJ/IZ9koD
VC/o9l1xliiADcqAX4pt/tslWoc6XH6fbTFncufJcTKEgt9PR6Ta/uMK644Z5sFG
ahsrdMyCLJ2BJjwEq5rfmY5u8FysW1/JfDkXLiPtHJtXc+K+AJIKGV8Y4tToFNcz
1qnyuhFuHF4cohpP3Vpbj8xEgW9M1nAIUhWir7HnUk1HQO5qO4vDddwBAthIpwXv
i0/0nsQ7MnwvHSKiZlqMcjDuEzbKHovSOzaGIZAQg9i92+LZ59NfwGYe646rScb/
val1huFS266ccT8HRBtYWjtwV+G1Xioioa3SIbGPl6t+nMO39KTjnjcVS1hcqumI
nOUete654HLkfk7vWUEMGGCfu26V74AsKN3kPAoT1ev24sQlxA7t1Y6OQVPJRUnz
4dozihpFwgTbQmFEXWr7H6XiNoMpuwmohFhmtLUru4fBixs+a+2jTjhtuRt7H63e
cew0IjfKUeGmzwojZfTQ39mOadVOmc9otnJqZBekeCAo0D2jv5MhM9QLC981czJe
W4RWJyNEGl8qwO7+02rHJu6cMpScAUl0TOXrd+WHRSm/v3eDibhlDpEzaNoOClf3
AXOa5SUyWXqHUfScyvhumbi5w2JgLLucN3O7oQdWqwci3e4O/t4tRj9OVkOSsTfQ
h7MXznpeCcUbrScQI+RKZesybZeDsc+ktS+voCAbJvnxWPICtqsyxj60v7cjo0g+
+FGP4KP/Y/rw4CSqz4pOnz14bGOzc1J3b4VaneF1RDth5RGNjoO+ZtZMgOkyMftu
SRzzzClKjcyAVueAIfT7f2S9ZQyMTxbM6pWmBkSjE3L/PSr/DhtwOROcYhMxAR+F
QWl3j1AGeEm7WMHuX2XP4OK7/o9va8z6N0rW+UfhZP3DeVg+bEu8+WTr2mnx4bpR
YbDR2+7f5UQQ0GBI/Bd8jMRvoA0kgvm5P3ZirEdui1rLFLcin9q5v44EKYHKbc0i
98grw7XwahHQI36GrZ+3jNxoP61K3dNot8vJLIWj+pIgwjgTxMkN9IlHQTnJHuQd
PhgVfz20oTa+Hz0+A6Rf0xoMBC2BY0kiz1nyRT3QrnFEhczz8YIkLs7yHgpcDd4e
te80sMA6Wat70BD/mvoRVuGCykfFncXe7h0yY2R7a9upchaeDfm+OEGIKAMuo1AV
I5NhX0zIbgJoBq4HrUMAeFXM4r0cJCMoo5blg/CEPQXIFJ9N0Zv3XDFjjaIGd0Oy
eSTuh1ycibM3raJWjDen2h5xEwmamqvIJ6W5rUX6LLUvfvWpDgWXHEGWXOEo0D45
f6TW19PTUh2U3j9y8KdoL5txJ0sRKGIjyhV24Tjz557ybzgOWgfcgNNDJnYRpN5R
3naXEIi60L7NNnaVJe3vt7EbO6gvHkw27fd2tL34m0NmX1mKKh0K8Y+uuxtOcWt5
uMVMw9OMOyiz9MpJVHy+TsAW47zCdAU/HyxLw/u+xnVB85XmVxjy2T8UGuQPH7OH
gzNO7TSXemw/cSmLLP55Wi3H4vpT7IUNeBZjVmotobtXA9nrdJgWCE+bpAaY4Pgq
gTuQZmUbCY4iVloFBOZYOk8eCeZ2wnIAvojzWE52q58W6nFLatC2qXQ/I+iDPh0q
QgnbSCCKFm8eAesaRuxSaPN9htnPoVARZkkm55dwuWaR2cstw4WiTs+LaG4N6XKL
Worpr9qGyq4fSahLC7TSb4Tak06WDND/mXOc7wYL6Kq6g/bPeg/QehNT9rjwhybs
s6pdrO6tkk1oaKJYS6nD8iBP8kpY+sp0gtMdK3UDxyQss7n3Q+ZK7oALIfbRIwR3
LFbGWC9m0pvbqzC80C/oACFeTSlnGku2ta/+cTjkhfbEmOMgn3YxM9GazX0B7qFD
SC7K9gGObRafK+vascJD3DWOx0T7CREu2qhAh3xAZyQ+y6JWJDq966Zc2od5KRek
1TEODYLyUhxvAA2/gtmlggAlJXGWy/EkXVNc/xENeAZCLhxubQdtIntT9nNUsBe3
AupU4z81ae4TJDng734eLINXjOMo8umakCe9JhivTvCXi0sjvhWX2Bbc5kgDv+AC
3B7hmHNcfKZivqNcfQG0xBvL1yX5E0pRCelAs0MeiOASXs/oi5CB36S7O5SBm1f8
+4/gcyFLlB+N+PSNhFqbctevU0KboVoBfXeydRbhGEcLZkyo1vrZe/HbPSG79BD5
uQiXN3WGZ3txMx4ulZyxzgYF0X9hYkRbRGlqNpGE4gSzoxZkmzYtluc4KcRsty8j
GfZGqB3lg9q6Jd/YOM47x4bLb+Mi1tEI4TClyWpKWsAXssIlImjam1RXqCD1cLPy
9g6MCtuaMYHYnCmM6YMG04c6QWxONb5G5cKenTyundTv85KXTjijpkXziADubXU1
uGQMV/DdsRALNqoMPR75CRop49D16qh7jmDd3bfBDPbg2E2W5i7D5C538/3U6cct
xPuwv6fjR2teynTVr+hkjM/y8CHKAIMkGtC6sq24Bq2AXAKJ7HXXLZ7yM19lxkVE
KCmN8eF4kQVibEnNJRumJhy5UgsOwicJC2xm223U0N4xZLmFyc6wbP0aUrGBvC1G
Ok/N1iw5Vrm+wd7goOYvmoH4BoDpZK/fcEBkrLQW475ufnWOu8zdgvgMviFLEtUX
ITV/rMQOZ5ZFPaWxDtyHowCip7iPPVUk7k80BazEDv9IN2VFNoizDylLE5pRG0PH
CeiexY5nE+89LsXc0fY5K6o/hqyVb+7hut6Yv9uhv2g1ue2cIGsKeEyZTyePgNk/
i8uROZNB8CMP8rTXqH4Ko/3upTrSURaJ2Ui586thK1Fqc7SqmOM0Eu6XTeY/bxuJ
h+Kt2595yHaToAm4TMYMOL7xhCAfakW8M6Gsurfg1Lur2BJka5YfyHj8IMFCeXlQ
bqQcJKvseAENWWnHIXE4j3mtzu9a9fZ+JhGvPEalAnPWJ8nCfqGGwgUITh4ytTxz
o7cfpK244RibROyv1s8Mpvwa0AwivOtKcMQYex0Z0aosJnBSIh4bwhX9z2Lm9YUE
RH3VDVxC36id7O5//c/BXxyKMULdtamwQl5l0iVMH/XsrvYk4pZqycsgCHel9YVr
Bd4pMeQghtS+xCzNSrwqM5yw03cDVM3VNHOUwBe0noitzhgI0SP1pwCbuxU9mL8c
JKu3Lufg8w4so1YmOQIzRbt9PVH9wFFUf7EGR2geeh5hdsRbztit4ezaPOpSJ4Zh
/H2Fp43jqcSRgQ4xIMztpIMo5EzQB+Mdzn6+hiXhrziRs8hJEg3fyTMEInxOOZvQ
iKAcTV8fo8PCReSqNk33jwn4CxhovnF8u4hYD/lCPxbkf3FM6eFgoO0lRq3DAH5Y
x1MYzpbsd0A7aL1ue5jen441gytgazDczsA5YjronrbnqpAy7FXuRAHgePSgU1D9
+7fC7UpqldUU3hmYq4rzmtSMW0M4yM7K7jyRlbqLkHePfuSEq6imFWKKjto+P4A0
13KvBZrTMH/VzB+nhAqD7FdVGbPgLO5/aTKGVPr5MjrU798+nhDOb17Q5mkULUGt
IelcC7UzvIreSa+qZAkdSOSjUsqziaWcFGG/vN9crF2Rd9ik2QlLitPdq71FIYVD
Vf5/G3d1EuPHMOhZhSkb2+TSVnnRexpwx+IA99olY3oKPlHjGndcL6PEjup2l+w7
0s1L17EzHKqbPu4h2ncniYBxLhOuZ2n5vICsZ7irUdVU5FRd4aHzlJVUfSpYeSHx
QGFvySa9RPcSN4utisI/l/ScIFkXyR3YCMSLbNHDJdl+MQ0RKoPYsRH1V2Z09MDR
LrYvwI0Zkth7lvHU5m33S6voZkFYSRAlg3qf6bMjF6YY6UIs3ggT2ZvhsuJp3Rh+
+JvDqOX95Kh0yROagYcHTAdFdAyCD49nZrH3WojchxgPN8/PGsssnW2jSYXsNWQb
8p57gMzSSM4BH1nazQ9vZZadc5JqgrETG4zDNKq8rChLzjdKuqC34YMyK2H3hyjE
XoCbH59B0JoYWGn5gStlOrhxEJli3SBfn7Ou9Cs9l+ARvRuHvQmrO0FJvho1TYpJ
4OJM0tW4V/iTxEum109S9ARw1Lr7UWKjXONA2VZwFGFDQIe0XqqecMy2UOciUpDt
4PsOrf/PckH7JDnVBGTMgXIHmgy7rORnwGCJhFkUAR0IZ04y2QC6nZpZScAMOG1o
8a8gECgdbG+kJYUqqvN367ZcNcMGtU/0YSjQ92Py1ZO01Z8eLCddvYcWFtYAXhAw
sX/vBas+vGLvH4QEn7qfea97/W3Zk7EmeVhDOmLrcqUkX/AjPC8YGzip7vOGlyMj
gxdLLChswI8ZaAUkmBfh0Out2EyweA6V1b1djUsfiDQTHV2KHrOJEDy8Rckcwnhl
/HGcuEMTu2hfpAyj1xS72ts/r0IqwPq7cs7jvR1xaCfkHeaGTKsIAu3rjuEbOuMY
kRliiUY57aBMdCtskFNGi0wQC5JIkHZo9U3HRvsgCABdC9nfMD0pTvYlae45tTMX
oAl467kGIIIScQYWwL7o4FqfbNwoIM4d0IcLjdoDt662ooHBqvXHq5w2HH8CzYhJ
qR+gZbQDgBOWowMdIYr4AZp9RBcNYP8iDqW21wY2Zck2xe9axgkmpcT7dQ53jWjl
oIUnyQhWBy55LykU2xKJpISrgheuiKsfSB/JqH9VKjC3ukLcf8msExPBjHsX5VBG
WwVXW4q+EDxc1euIwFtecanh76NGV0puqk0pvbfIoIfxyFCrhXDSKRYr9qa5xm8Y
f0q4YmTdg+BRV6Yz14OJ/2+rumFKU7HbM0m9CcCYl0F29OgVk8W1nQ05gdYYZCVo
iJ7dftLmdxenk8UqRW/ZYy9PmVAfO/y+D6SKpOuwid2PLFgyAGdFd6t0CHyyFJSz
u5tTd9BOmnWqq6wGYEYnJvRBCOU5o7jNc0HL99fUvoEf5iIdz0TCVLyg2VGni1R7
IR94Q5MSO9U8muZjnAfDHV67Bp4gu9N/CyS8Lpm21tbnWAY5GGRU9x/NYiUhdqQk
i5gu6H1ZuLvay/+UaJ0mIUOIftL32CQ27hOFpcF4IkT+QMRPsxcfVGUmGGhbICdf
muc/8EpUQ1pfAEJiFwz6/RDtXaxgaqIcc3QtxM0bc335bbKHAmeYO8NdNci5urr4
y8biOG7f+vqDD21fFKG2dyVMtFFlE5vwX5H59f661AR6OQsdiu9rNgpnAw/UAQBW
OlM9RQlYiqaRRmgvcohJNSgw3T3SautD4CwCcpFSKdgSDdnu4k87AIt0LQNGW5vs
0+ot+kOtmnQV67Hy7/fXZoNp4XchG9Gkzq0RhP3eDG8IVWCv/jhdNcQeSXRUWnJD
jvxqg3zDXNeTgk7VP7m9Pw+eM7dGwDTtBsDRTY2Y64V3CBIqKsPlq4ZPiiQpUYh3
mvoyMdScVpgPUWB0+z14FFpwdCcx0ixf1QOifAqpDKgEBqB/xkHXbuhAWzJjnPqo
FJuEFYNQkK1xyWUssDrQtGxVlllvNnEboZoIihMi6pQqnMAB/gw9SdboeZU36VXK
EconbtwlE31RTwcmkWCvaXkI+Tc7pmVbPVoZsN50tiAahGK8hXmaVLA0NErEb8B6
JG4Hd2Glko23nXr5ZAC7o7WE3jFBukJQumfB6OM0e73ncGlllckDfnxCVSaYCL9p
fbv1aBxtlahlw/6RQQ8BOL0z01BwYyC+Wan/pskf0ol4gap9QHkqUatMxCp68yig
DrMYQf32w1fAoXg90zKR4bTGC65b53WnzFF19uuX2JNV1v5oxCiJaCXDQWAlTN1z
N3syaguQ038DZjLihLU7QEiJG4F4GPE2xqxNQGgpPa5VROUiYaR47NG8L/SXSMNY
SxVUWY9E+Tn8YXJBVv3IYFuq637aSta6B2FXkrLXl7OlnTWVCS/O84oQX3U2qpiL
53Gy2p4sGZMt5m93EGk+51z+vIzvj2Tk//kYL3X171+X3Z/AVrU70vLu91NfMAKT
058wRxiIKAlX5ttG60r7Zcp/huNPlRWZr4EgiL+W/UWuvHL2me8cFncOQdqcH7Ho
k7XJBYDsNCvAxXb0ColEZ8g41u+xqP/Hy3kE1ubaiRelYuKi0S2iTiRyXb1wa0nN
PrQraQfr9aSCn08YyWtI6TvZEhzbEOBvleXC07mRmwJhLVpDkhth7hFWz+UWfQ52
eZqeLb3YQCDYPBsUqxzn6CGRvbbfSbpyPaxOKFHPBxCos+FCzVfANJKbhebDXBvn
9R0XFMqNt41inM3s4fMTfE30gU900pe+ibx3CY3gnyFjHFLW1IM57X1+rGO6N2Ot
AdqEWvrzy9qgBufZ9KkU5ieKwglWOigDshOWbtmpKDHoPJ/iGGwOCX2bOaLWQew9
UcWKsbD2EH5WKiPUhrsJB/boJvaTJaZesbe9spVai/CPxx2cq1x0KvfQYoOHot1t
apC9HERw38+lZcPKxw525x6jBdgt4TfsxlCJjYVEvPe8lSFl2u6bvmzGCKk83m4s
wLhPJcshMSgx/xpQAWE/DLb7P0MbIdZnPEezW9zl4yPtZbw5dyscpGvnDihFXtq0
f3/iRHVHJ8kgltZmaNX+B+kWJ6iqcO6hX3RVNlMDnRwYtxcX1bXOD055WupDnqdU
dqm7NP90XOmTSkzV+ccB+mKMyDVDu5q+loUNTEBAh9SbutkBbVB9gYZcQN+cqJ+C
tv3Q3b1hg4Zq7AX3c/b4sULHfLqEBYuHG4QDO9pnQshDOsl5qZIy77t/HnfBZn2x
IY0EhbC6poaR5STU+nJG3bb+9b3ZnHzrwkKniVHlGk3EgCJ9wVAdO2BK5Q85EsFp
6Gd5hSd+7e9wZtkDdNaGiW1IGEl00e0h1pUBkhn7SbSPVJ7WaLoH52HSB0Flv90o
jp0qzSH+mjpRclClwug8s7+nWV9/8a3fM9oB22cPfKLIe5sZDcgUsgId8DWwplXO
ozVYA6du34iqSnuNEAkLf/IBX5KSjY14RFcYWo1Do2iKJUe98PzMmdPfLiVPTCKU
BF4Y66rP63bDAdnB320boYaJWLIncc527yHyFbL2sEVG7hmCt6ZogJno4mKYxZXx
JDMQvaS08DbzYiFCw3sAQzSfplFFtTSmyHF1ykC9xvdTo+QDftSZiMib8yeHZYfT
TDHgZzgjbhh9xkNFM2OR1c6IEPi6Vee19RG+zwvVMyax0EQl8mSMgrbTWooSeQRD
NRB5yVNsr1I3NkRXgyz8r2Mfph/Ri5Iq7xTnnUjqtQolw4nwqR2Zi1ZkKP7jpykP
fI0kZCSyfYO2Pbop81XkWF2KDst/li4Ou3+20Qre4t/2xPU7pTmw5lJf3pIRC/oj
gxTa59A2MluFFql60MkhAG9h8wQOUTMulvPG6HVzHKBGhh7cPjFBqoA91oN6PJ/H
0ZAxDPrCbpJ+mCkAVNbNcRgKdYxlcuVofzAFz+rNcZOCLoFRJ5fYaUWPx04wpoPP
nsMtjvYA5moBuwt90vAkTU7KuoFpxO0BQCKE4beWNKqbINpVhMWKHSIPUx/K1z8r
tDLGxODW5B/5bVAqV2Dbgc1EiWhYpF0oA6lFuhKRezWpF7ZsGYFtAdYNpK0M5iuG
AxZCxApokKu2zNDpLMv+QPQIPbJEw3umBPErLavH4xbc/803QCbz+kvZY7vCLBc6
mJpVN/2EptvKZTY9ZXRPvbVuNHE+05HwOdBBevRNhDRDGngKkh+UZLdU2pwFxo+u
8CvaooiT7Qp6bArNDPPDe6dG0S7PXeZOzCq7ABBSdRVd3sOkG5jzC4h6xwagJC4e
UA18czASHTaizcW70oxd5k0+l36MJqBH2pvG6onWaFR1N1Zhuwk1O78zdmrpGr1p
Y1mRvpUMU+9sCQGbQhQeMn1Eu0rqiIQy4kDIkgDaH1vHfC7UA6QeoJsv6+Gc1EBr
6l97Ax4+nTVQMmsdWA2UywSm9bb8YIqWNh9aiP03gW1e3/uOIbUQfUWt/1lEeSXd
WWevi/8HkLVJZMYNn8mZTjUW+3M7sChdGnhmv+z5N7UFCS3FBKZ9SWhSLQ/pmG9a
cM2W+z2lT5bzkAbL2wNLQWiLBHSpZKqjBj9RndalxvLt5fvecUN8UIv2/KfZQ4JT
XGdZxnnBBqkAUkXZH7ktGUqQUsx0FoW2rXe2eQ5I8RNrG7/FQrDs9wjeWYstYUY4
Pf1WtIQiFHw1SyUPaASh8w6wkGxfrudF05i50cLQjTqkm+NXXqGYA36y2D7ajefN
BxSFGGDYQh7ckN3A3dtwIuU1qOOelWVtZUG9amuDxav/liQmrE3PZYbMl6l9JM2U
C7KfxF0Iq/HxxWWkFMYyyZqPdExFRLuT1a/Kku1FoEfM0uuQnxh6d7X0vIvcMvFr
eLOHnkIXnL0DehRXyO2yF9sR8uhJ1TZor95ydDu9NyY6olX9D3BkmvW1kGVgQYlC
4vUjlvedB10PTgVLXpK+No1aRO7x4LXNV8LdH1OYKkPs8dCneWQQNiXFV5pTxx11
/r2cBUssVzADGmuLoC2PdF10Pb4GysWnDReL6ZfFIfUE4MHSttKy5bsb8EVdgc5q
gGtRr+vO33WaWGLdYwmKoEZ0pg93gE5HJpDb4816szlz05zXwe5Ugs1epl9LiEjc
O2XtI+d+3cpaFwKyVcV0CetRyZxbOFwrWVPFFTDNY32HUs5wmhHnWZmpeWeLlUA0
othtMLdVeitaQj4+4xJjlbySa+4mcpyBgTxzbN86SHUWKmVquK8vsqpYv5EOwfgP
z7iIzINAjdoUdMiQimpXyWYAqNLOPwzZcTZU42AZcYpsvB+UfURqZm7/FuL03eYQ
ullkky+bJAf07EZhy7GuRu+Ys34kUr58OaWmqo28kFLGBdLxn86dt278m7ZggQSQ
XrNV4KNbAss9ki1qQGCvfm8IrTQdItjiWcMPVm90VdQpbmIZvXFVeDC25bVFNUn0
01IOm1Ofsva5P+d8CFpS66vvLjMRWpAKCG0hkrVXxvCF7NTqyIA+vdClNYsckW7M
VpxPZS4OVmsKYFRxEjw4UujDnfRBRbLc2F1PWEkkkRHFMjFgbPHQQTXVW7VNDJHt
hADo0Eyw9lnp4v3yQlk9b+gsJwOS5tAMSOZsp9Pu9IFUNYS2OWJ+50fpI8PVYlcH
ruPUZP18+Jkbo/iHstZFVUAGP00BPNbqvmryjvKlJ0Z+GYjTr5JZ4nw7tX8RbWiN
HszZ06FHu0o3ddkGdGlKT4z+dTzQ3OjHFx5uB1vLvVvr3Jf0kTr0Fi8FpiDCGDxn
N/GlGHjphMuX8H/2mPPLjSsJHqbCwkjO2Dj0rIfIgRZ27drjcy82rarxO3Cy73GN
SBZhP9NSsPeo6hZ523DSaFMiLCR8YC+EcjbDd2Vp0ENc7/n6rN/s+CvYIGCkZbOC
pXgEXOkONRP+finJpsv8VVzE06PhflN2zehn/ukATv38msc4Q8TosQa7ZxaGWim+
Tcvw/omRWzU/x8ZVdQbW55UhfqPszxbsiLjMV5ULs+z27KQCJMIgR2AFVHzDeSp7
KI7LyYK4qXBifyWxEHCoZi+Otw+8DVavXamZuk30sRWn9IDOrX0IoLMkyDCi1MRK
OvONlaP6WJwPDAlefZ+VAWMFcYp27f8vGPUELTjfEQsh9lzEvRCPkmhjxNmwCghP
N0XZ57qHrd8oHRMxfxRtHNafOOkUIkhCggCnJt0zzqANe2ZNvF4+LNBXpHNFkw5E
A+exmOtqyykI3E7vXEhOJ0n7Ehi3/z/ecDE6gUs9i3BJaW9mqV52jBY/sky5VmNn
OXzQCznMvBFkeEZNAaHx/wFh20uWl0s3epxuVwUWH/v+mel9dD7Gaed0w9Qmfyne
6HGcSe+4zRG/dZAz2jgQeci/vHz7GOAEoQsdY+Le6PxCqsmz4qVM/U/y6dcf1oA5
wmECNqavz5iyKwTFY85THLn/XkitTxcmBnuefDfqFCjWy4MjfFwEMXMM59oWvgn/
EGRbgpc4Yf5Gl0H0egWQ1QFCtGx6GzAG1DoWW7VP7Vzh46EYBJTMCWSJ2V0Bhoko
ERCQy1FGroZuT3r6qlGMElyUcYOPHvvQGm5x9zlPuh623JOjUcC2lMWnDqrIpvW/
nQMIXbASm4NlMLV7o5ZL6XebIp5qDBsFlFd2gEDQat4UERueUDAUE/lNK8Qw6erP
Z1eBB31DNXUIab9rJkAbyXbbigEC6+GDA/+54u7Bjd59HU1aTGIMpX+QQvBjUUi3
E5X6CGyZPovaGIQMunQSKX3A86plivskqIDDhCuRhZgcLcdT+aYzpSTboG4ncf+o
p9HPUO9oSi0D/9yuHWmsHFO3JFqg27P/Blq8O9RAlWcNanQW9YLkQeMOKwbRlV9g
HT8m/afJCPvIb9lQd4QtJtr/PzbG7lB2in1OJYbJ2llDvmX4fXJVNqfFUwQLsPGD
lLwOovivrNYi6eII6PPxCbT5qHtxOmPxwSQwENO98A6edEYp2L/DQtwYtlkr+GW1
QbFkt94Uki4kTcdm1rUvVTahjEvz9otbUgQ3yy6aP7LZDfG66yqkJ3Y+ZOlMhUTn
uC91jZBfWaBIuk6WzCPI1tI15JSphhI9k4aLUw9kbGSwHiQ9LXiDqW6j+I7RnCeI
D14WcN6Cofc8/kdyxMthYK0ukLBxNuqLHISuwgkJ9fqFfETfNoCFkE1pwh1Rd7mS
tXh+HJUO2kkiqX+3kJnHK5Lf1HRk3z90la5yIVVuq+eM5Fk3wesxURaSJAZEXBus
jTcMmdxvDYEspkA1/6uZZJacOEIDF+H4g4UdtKdKoRBogXob3+9S7A+vHzLVFYc4
ts0swVsIjLEuUmW57ZiM63eVmMdevN9DBp3X/p/vCdf29+yai/TaVQcBYKZrRczY
d8PerAbIbmRtmNBPB2h9pcMhcF1L0VyjV3hU8fz+ha4LFSv2PqUHCXTkxtQ9XLP4
AvbvE2rpBUi8tvYWzeMkuLLClRuXHMp+Mftsa6MuPTyEnUoIZAi/uduJ+N9CImvn
4E9uA5+YwYA5+foiEeIeAuBduerhzphwpii17js0ZOOGt6zrqE367dWE0uLCDTCd
GEXgqNjzYyEMdxVPW9wbib7asLKNOjMwGOObdVp2zgk51NNDoITiHtdletpNqwC5
zelt7VJSEBBObnwkg9zndJSdJZx8KHJCs2R9OBheBB6KcWJh2NVRv6J1Nb67MFhb
/bvYty6lJbeDI7YGAnj7ZQsp4dQayrt8blCOSClyJ/3j3bPLgMpPcnog0/bUXoh7
GBt7I/RpqekiLIeV6dN7k/F4i1zq3KhLqoIRZ2Pz8F1wDQ+ji13XBXVjRxh3dAeZ
YjR9iZtHpidm0i2PYgJDGn8VS4CU56cu2ExzlCBtfKIUjFKQkuTVGnHY/x48K67d
w9NcPsWZ1J7gYce8Fw1ACGnmdDAGJwnge8qvuVJAj4lDP+MDFBHMsvEAAPZK1NGR
15brIvS00VBpIKPrGECHDaRy7yXI4XgANpj3pOrfhbKZVSzTUoigkPb9NGbJGnvC
2XA+pdUZuVQSRe6Z08+uBW343uwGvfkaZu8qHyNSYvoUK5nrN5z4KynIW+50isrS
zPOnOa00bfhj7vBpeySmtYXqWsrYNsKv5u5R+UY9MWc2BicOcrvQJ2y+XyKkizhQ
Igs1ONkIMmnl5k2Od0kemfnzWBJ2Ewo6sxc7SiOvPWKxzJl3waM/ATr6qMvuZveO
U0p9Sjj/rdGpAztQJ0JVCBUM6EVh+Aao+VXIa5I7GMO/KbeH/kmoFekLeDKWHzIh
gU/ABfV4wfpZScC8DZQh7Ea2g9MShClS/Q5OqZjrnXQg7h0oNyafNB+DJD4qRRSC
EUvnmAsufAWZeuW8YqV2Xxvl2wjvzwHC+kxpHCwUqJmuDiih3RJ58A4oMaHBOXZq
jS2j7L/PKjdx4oe8O9KKeDo7MheSI0XgldQoqTd6SZEAnRU6l4jMYJHT/8vQW3fA
i9IQfJqG4H7fSYK5MvIe/rGbZ1qQv/4xBAAwHou6s40L9WY8Ub1usjUAyGtr7cP6
honnbStJPh0M5p4WQZuRbm36UBrImsakKzi+K3rNbXO7dJkKdxXPyuYZo9VzSTHk
tOAlCYNk+l0rX2ewl0Eq1em2JYfiahtIetHzCp1AkClpLZcdPnjTioRItB388F5T
JUUFrNmQVqz6IsGsseuMf6xgqYhaN7dHK/ZQbel9SmN9C8mOjPhQOlMj4R+R7Fmj
d9K8XDRTpscQT18fWBPHDdkTc9YY5tAK24WpRNsCl4IgjlTSdPUE8WEduidOGR5e
THJNgtMG2078tCgMq9+n91S+9YmT+3wSA+pS3UlQWe+f4pwNl1VfN1jZnx9geLRi
WMzgNnZJzlcxIEzlkeGU29pBvnvqvE81FVyM/zHGmWW7Kf18w+ahhUuYJfMH1DIJ
vjqM2fgWGPOh3cxr/Gyg+xIj5dQxT+zias8gBtrDbjmYHkIBIU+Pnrp68Zq8YqpH
XHPYkI88n6QKQSah4DylMLySUKFjpEW9suE7HRmZzLV2tnUCPdVGVl+zM291E54o
2pY/Twee7RWCU9JzM645B6KuuPvv808ffmdgExEulG3N0vLcPgMfgyRPB6S72vDl
385ZmWX5523Y7jS77Md849UdzgkavoCRNnH3dWrGr9ouX36NHWpWZpuVJlQnvCUQ
hkA/Vpr7uIucBwlu7qrUdJL+d87tm/XEQbtLSgypRQzdx4O2PlwSdQ4JPXz9bnP/
pBW+P/GwoEqtds6PKzMW0ZNbCmxbGdP1Ef1v1W1jlbuolQxW5egKQpXwhuYh7nSw
weNpgYM+asBgXY6HFAimCm7CwjKKBOgldBjFzLbeIzZsAgoAOscLhMB+K8dOYdtf
TIXXSbu3E0akaOHqMM4qgPrlN4xMVTMkPMtwvwkgPJ6A7rDA3MP49IcY65w99TdT
lRwBy2aoF8TsjAgAUPcuzK5IGAwaQqOoVC44lRFPMRq63i3oDFX8jyB6pZP0Xz7A
vXc6KbEs0nDbMWIlcKXcUC5iVtt01onTfRshiAjcNYfZuZz9QkpF0zEz/9rPZgCo
KGbpQujQQXB9KaQP/evT1QkRoo+x2IagsvhOfTxcsU77YL120F23MEd7L+vYSG/c
pISEomDSHyMDvwXrbDHjrvJyILSsPPOROvRVcZeXjwJmweKqiuhGTtEWYHWhS9aK
v3EYZoWzKZ70+VPhmB9pZQC3MfWOTyD/LeC5fqUWG6yp99KlIpPpl2yvp6OZhMA2
rGko9QxbA/se1N0MiKaAhZ8YIuIfE/WQWqkVXzBaNwmTHimoW6jNJZp8C8lQKFiI
niCanHLT8eYv9FOu+2f/IK/oo2MZY8aLiaRoWDcfd6UhZa8skSwhEEqhm7gknkYD
1Ifi7BCnVlZ5/SrwgwOA1Oi8/aJ4hZYDCDbsGOEOofKErWKtNIG6dJfre5wRUOYH
sZAOZD2mO+hfD1JWZ8JVY7lKKxuQxH0XKxhzjC+m9hmogWDRr7S8X2v4pOMM1YE+
5kRpNbt3dUOdUOk1bBs0y+xdNGRF+hGpqCU1VnLVEEFvld7nPD+sHaD3UChfgqd8
ibA3LzueQdEEUnBE89EPPgMACBzZqR/DBZ9Qr83+DH5ZaTF0WfOCnmNKMGtKwIIR
Nqmd9gzH0K/KpdRxxuP32hvH3y1VJkZUtW4BVUWg/OXsamWCZpW/MXhVVwvl/rnn
BNtN04dpGadNGgy5YwnDXBOYAtOiOIx4GYsaTQFSB0oaNEx3rLT9ukJb4HRIB/tP
EQm9V09h0IjP1smZ3Ss4sxhAstjQFik6ixYsO2eAp3RJMgCw76IgAJ1CEaIZU+lO
sj0bhtiOyJrkm1VarJf0gDujQkVFMzaT5c9PqSxbORkTBBrHo2DBBA1oYUqlaIL8
ypCKeFB1sHwPQ1xfKEldM69b03XVCwzrlGkjH/oQXNliO9nMnbm0NhhB8JICenoN
I3vx3nqOGcb7aDx20+oS2f/y3O0au3ysTdcDCaF8m/TDP+I7Pagp3BGRMfJ+WMCL
CFprZ0Ijy5zNy9fKDcjX1M9YpvpRc2L7LGrfyah8oK67DnQ+k/gqS7k1+irALSWU
Hz7z9p5AfzUFvx02gtHbstvBxDY8FtGyMps8NF+X8a1iWKAMWlVdq1n6tEBgnRd7
JeukV/PrqJWojoILp9g+qlSv5P2A/FSN3WmiKaucfaiQEPHA5ASNnXxFCu8dqlbe
79DHPYUQgWEmk1c1PvreuRk9kjEC/myKmgdURxQUfB2Rm9O7UycCqBI3uaB5EQsj
HCQeWkEz2f/pD/Uat0a4ZLYWqKPJnQS9EBdKYk8+ycWEw5NOonpUDHLyrAarWWzP
6aHoZwGGMHFOxD7k9iUYflBbiLUYkZE0Cm2wowf3VDlB2nQY5e5+0ptAd1artrVG
ngLMYt9/PBZ76QlLsxgYgqLGJ9Z+JpSEy07fn2pYHtNl3mvyNAeraKxr5B60vtr2
PGdnoEQaCbJ7PGoAluCuxmVYQakXzbgTBNxcG1dvfNzm+2WC1RdWCyMk7RkpCyrd
m3vb/szR/RT3mzv7O5qKQzeVW+5gemwGTyUjYWxsv5oX4cEcBvvrtaaraKNvaM/P
EkHxo4JPj47aKRjvBd4vSGjaFK9bUxUMebz3hPMV+uIlM8ata3X3TUHfQhj9KtKb
ul9cWi36GPOw/i5uq2X902ItAxnlyUjYOzxohGeWgnM9oTsos1QkuXNRXpssw6ZB
B852dVdw8xuvLUTjkZuzkXcOruTy/gJGNA86VR9m8d5w5j/n0hhdJHZKgkwFC7HL
8e332Jq5OQ5Vxtn1Ti1MTWKWs8RLMxcK7lKD7wmkcpwSlRT0ud883rWEll4bq+uz
iwbsrnTQqTCd7tEcW3zKWhbyGoI9vUzjllf2Y0f3Mo0budqQGoysRpEVwPNFIEA1
37G2Xli2liGw65MK9AxXdDT1XcAHLCFlSSwW7+/lydLm8b4zt0rZAK52VdFFzauy
ADzvuXHvFrezj3OqzZ+5Y2NVkZ57m1PsN5IaabW9XEQ2vcsAKtQ8ZBrRN3TvYeJL
h3EOosJAn7wzkBUV/vZ2Vm0Q9DstbfeoMz1SvamjeX4SWiuZbxtUtrMb9fzWbieM
11iYot5autPQQSUKDyRYrKPUe8Ngw5AsoVrz6vn1PyQWTAJOxQ6Sf9E92iCXe+8y
ITz7I5vNpxdFMh5sLBNMgCPDHiaXy6soEMu2Po3+rFZYMf7TranolH72rT5OADWu
Dr3jgBtsyxGj/AKE4w57Z2BmzuftpC3Gw5XPzWV3LR+JjMZytgHjEXweLGXygq54
Omh5XTyDukPRZhjfewpwyN+GMJVyQmaLjiJaBXYKCxiD94ceSr5VFPIH8O+To+zB
BCo4sl8eqRLNeoNCyi027G37m/p+k8O+rYar4xDHOF9o946v82yy9KFVROtl9nkT
N612dARHFdFI3/oeVSCRwuYYlOfEI0Xt5CzYBZ9IBioqedJz+z+PLCNCmV8MvIx5
JZSzPXlkYzPkE2Ah68FZ9Dgo5PojBsW3v0YWnXZpwzSc+OkMrCmcZIvxZZPpL6Pg
jJeqoX0FLTHSJ+9A8GpsZNt7CWHtCBffvXv7kKrg2O9YD3m0DkMTZGsX4VCkdssK
9IZ+PkMvKYPiyKLFn+7i1bHE7g9WCEi30nDWDt/Ax8BjG/82D9Fan0yIh28MG94N
IWh1qkmwaV78ZnOO0NKyssY8su4SxdJ2LDkmuMnu2/PLEUPyoH2hRXd/ieyWmVg3
NewRt0JcuVO/AbQtOPjxFG5QYEGTYZTz7B6SsBDybFW7XihH4rTPGWiAaP7401uX
qOJR3D0OFhPzfsFuP1QRfy+60/ltINVgN2rUax9yEhrTDtQ2O1+tPsjRLnzMcYcG
vAYOdK6N8sAF1Nrn/NsA/kueGTQbOrBe/PSIXd2+TGQdHN7RJ5LSRbrGjIM441vc
MZEmauzAhMH0YFSNhyf3abkPQG+HWKCzrmSipZN+e6tsdE2i5rt1OOJcm6/SQaQe
5ymSdZAKyY74dXpWxw9Q+OrXHEe5LdOGP+wSt+me9+SF2eDzRhi5Bjo0GKFZLb6J
FKoYODm1l5B/hJ/wsmPFwczJzVAvd1MZR5bY9axd9iEMZVy0hpdEYFzmv+XURGWQ
qzBABXic0StlvuPRQ0KvnnGjQuban/Jv8CMF8Fd8RJ/J+w2YQAqlTHOLgtE8FU6Q
SBx4egKjUvtIQJcwf9vHxPioHZNy1DWXxuE1XanToKeU/AsrIjQv7eI0Rh8b+Adg
2PlALbXS1njHWiDnSbx8PVxbSywZ+RR7LRvsbV2Edf32V5WJ8Wfn7RWtqmszLFxN
fQR+zAmz3R3Hiy97RAqWErROeXNuca8sBItNZ4l7ADULXmqwEQokRi7Cpa6Ez6Gk
QjlNbU/AmrbkLqghwNkeRjgIekZWJ3svQ7oUtIJWvsP2CyG2Xqz3e0gKKf8kZbcS
FPhuFELslQXnTWB3ZtNATugjoJhEN+YMWcVmTv5SJFr8ZgN/TMnULR2xBsvLabvA
Y5Vgk05rsMMdTTvwszCBYA/Bx+iXtjxp+PYIt6VeFTB7u7OPOL9c1bxpifVW5B7H
g7oJYEDJFlqyJgBsnNtuho1oMdasHcgah0A5a3gRJRYvERESFAok0v64OoPEq3j+
fhnI9nFGyj+3uw9Uz82OmkzS96D/WKnvFH4ls9ZATL6UZ4vAx0SQtjKfIwvMqa7q
qWvaEL0CKZvRjVmU5wDijuhCtMgSYMCYujJa1P01r9KqwsgDLaRTLUZuHcYM1cnM
b84EPxecBa7n3C9Wpiyo0yOpFDMVmPz1+CdfZOCEAe957tZRsF5AcfA33pY1Bcxy
NzU3G5ISGEoU1pKRW4g74CkGoUDaAjlIAQfu6cTqha0T9e3t/ua1axqDIOZwPV3p
eGiBls3zlpdsUIfY8C24fGcnZrwGhdqQt91kBz6KliG7OZewTRScWk1rO8MlXXoY
voCpSLlDEL3oCzcBQJmVn5BD8s5EfXncfJELr4pxn/DdnAbd02VEVvwEStuD+aJd
Kud/DnfwlrxeRwd3FNML92/O7gHJ6pUV5vRWs1p3RK8JBlMMLZjgDgdTzTAQRemK
FN8VmnNRjPwlFv0zwG6x+cOryVqAWXHHSTXlXCeQ2Dm85dA5KWyqzkGASSbh1ZRW
5S0JaZwyv6deNSGNYoof+isi1hYdFUseL+okqK1TP5j0lnhpHOuJNbfEyYmzj+wN
MnqgZpDT4FXtkasFcU0iVaR85YoT0tZSTZ8Nok4mzuEF18QtVrIO9Fx9kDM+n0B0
NZMP7lK4pno97fDJuc+v5wjuS+LWlaAAqVmJiF6PbXxXMY5bz7ZDweInX9ydmmnC
tDepbeKvjxKpCHlkvbOH/Djt4ZzM7RyCsd4UheZ/zhNaITGZScavMYYfvUpw9rPT
iH98GSiaUdvn8iKBFthWiu3Jg5bLHLw6zQw+7laO+Rss2M2oHBxzpGTd00b5ipcO
RcW7Gb17tF9aKTnS/dtVz3C88PLc0aNujprgcAsmdunmCSMosIDEQL67cq0Vb5JS
Qgg7k7hhZTjDN3zkpr4Y9q7YWmD2sCONTzS1CdgFJTwAEztZtQyatzovIxmhUdTW
9667l5xwEDpYMDboruQIHraaTuuUsnnuwxrN5jT5z9gNlYfmNTNSbZapCCfJLnyh
oA0quzR32MC/NPoxBG9aUX7t23jjBpp3CEMA5EJsULFDQfE75f9pQbdUVCs5QDwd
v0TqbhlN4f5feTOw4umvbw05iU0KTjVg0j+dKdS3dmmqJD7+3csR7Ue73FwnCI/N
u3qgVEDBLlwx7+8xLIVeeyXF+qtpbwdjO5wqUZ+75N7QPY64jIaSzq1acE/uuvs3
l6z4WH9Em9qWrfniLYo7cuzHeWr8Bie8juvqvj8Llr0J8JbV8pAZjm8ivczy7vbG
m/G5WZJYtu+qf2BhEljL5c4arAZQyGB8uNGstRJs2pWDLpq8UUohZWbo0zJ1TouP
SSzwp371EVqrd2Sr5mTgUXdzhujeRwSzQg1cVXzE0pPUNaE9PHD82MpdRxdWDt3m
6Y9uOwzLmp3x0p/YhuHtnYIXsDXSJH1CqupsVRe9PBUkrefMAItv3I1y+GRTawGV
9Vt9COvCel+ISNxWbJSdGU/vXUZosJqGcRihWDDVfNQqck4vZlqrOqroZdVYNAGe
V1sAj2wwKRsDVUPrLlp9hzY+93YU4OcXyIjF5bHQl+KZ46Z6raLu7m0CMgMpX/Oc
7Vjn5yyjB8+sItdBhrJSdWWjsrzl/aw8Y4Z3f+PTkzOZMFYEcZWmrmk1inrpFLZD
UlFCB/ewKlmX8myBMVw1aBaN/gWLCwOSEry3qKzYLlJSld3D2e+3N79uGWvVKg10
80ztWUI5ZnDlhyT/Ma0NAjH+Pio+9zbLJMwWXAgz/paJzcPJxDCFgM9FFq3nqdQz
VHRFwa5echzAUNHawjz2mJCYGxa16enuoXaWo1HcMM3otsGtHrlZaMFLnmtD3eXZ
281Q8+RNrs117OqVnmVcpRS5nj4ghtsJ3V7RV0wfzT5iiybqKttnkE7U15NOUyeU
KDe6zjqmPloFTg3/85jogHsuwfe4Km+NiqFt5buAdD2+uED+chD/1r2imFJoE4Jf
dYz6XMH4fKMtaRkb4HxFqBSJZb45tTDFuOwu1MLXOLNheWVk8g4N5iJ1emZl7E56
vmISNlxnKzhA3tmiIk1WC6hXIeEftmyS190QMDdZr31jy4pIIylheeEqy2ol771d
zDT5GYREsw3YmVgbJzYmRU8lAM/wGaK87K5biL7x2U1isrzQINTkrx3XyhHUS7R7
2y8mtG9WpxChH9aqMdy9H/Bj1rRnKoiO26IOpx3Gob9c+bk+CUjnPZOkD1st4UyS
BRz+Q7OjAhZx9yIUSvdccc0E0VX2wA+dPUQzYCh6uuUTycP3bOtrnEoaXZGeXUNB
742d9IlW6N3wunTNLyAcPvfWIq6WnxwZm9fGzidIYUnbPW8zZrpVNjQiAKlWrxsP
576ulpuBB+6G0z1jQCwjvxayFP1IRf+FU3u5TRwIaiMC2V6H01evpzszCFredp5U
uwcccAG3Ai308C4C+d62U5674TUt0jKUYMgMyq037DwVIbiolI8WxmGeEeJcD/LV
5pMWTwdevkotDwDxAR0ZzRXgygC9dX0JQRFjig7sd9uHpbJ++BGVFNfamIgU5xQB
K7fNqe+/QnPcz5Db8/C7nq2J6MdFiKBXIlkg1dEkNWwG80Y68NrcHJVjTFOzEEQ0
G/P7BS6a33AKdoA8una1WvAtp3SWyUQyjKCt0J/q/zvE4ol/Q8sOWkJAwdGp3anL
+dapP0oqn3kuPII3Gx0c6LKOxMbHTd+LzeQJKG2Uoe7AUlKuHnoM7jFUvnwzoWNy
XNHbaIf3uu9GlosTgmJ+y+kWZCQprvRf4ydLP/Ql/t+UNkym5Y09XB8OToymgAvM
Mu2pmf5SSXY2BJvIE8QV6+BoLHZavS/8bzlgFLhxtXFIGA9SXuJAdefPYPmOQzVv
Bwche/jIL8paeBEzZsoPGBz+gSzFIMh1EPdXYZGMoHPs6Y1LQ4p1OfPwCTyZzrh/
AvLvxoKXGDA8GDqYur5nmVApuLCR2KFW60eLjc9XgeVFj/0lS0XMLjiLDuHW7T4k
5f02YujoayPEyLqRIvnpAqL8+mR0MtZmYU1heOZ2VgBHygmFwk+WqSNxlmkWfjGQ
7P8ETwjoYd4CDdWHTXdACk0JSrlPz5RRArlT+wtjJ7FGYrAbvZgGh0U+VZqUVEJZ
UXxu0xbCK/crr7ZlMReyKtbHVTLakDYFbBD4C1He17b/nmqQYuQXTmiJmZ8ERCNY
fv7ufZVkIPwEp5eZW8+NSSJTT+mqVz00OeZlBGtq9n3NmvhKhrtdCtBue8lemeV4
85xJXObWP42qvl3GrFJsEthW2snUb0c0kPt6MEyJyjnJjrA1lRcFSlbZ/883GWYI
8xn8cCTsCVRa8eIuoxdgbXNiAX/NHKYneT2r82VEvo7jSt5u11WdhQ5SnsIMyAPV
H5WNbQx6ngEtERSexYsBYIPCr/D10Y+c7Va4Q2P/Zc9kfWH7FPNpsO2LvL2zFfG+
6OOX0ROp1Ko1po+6tpKq9qjn5phyaZOXFEnCHtWqvMcQ/Tunsr0fjKi/iZTVFolX
J+9Xhus5/4AU66TPMi7fMRrwlV0t47b2WTs6QheeU3HRX8YJ5IrJSoJEzSDjUwzO
p2dZfBB5t+5/IxWPSb6hPaPN8kurFMq5T467qS0KHpYePMooMOfU4MM+lGbA521b
iJVfGWqSaL0z0iiculy9kP8IGZu3IkOsusPCBHvfYawXACnvfpCjCnJKZaMfnRhl
eTC3bi99cDSeoejFJxTYFNH3xdC0MdW0+AexL8ulG5+8Gj6vK+parxgZIK0B+dXJ
DEtbWhra5ehduLu795v7MaigGOrTR3kshijeoBzCDeqn9enVxBX6fwCsKNr5wi11
g60Kl1fETxH/1UuZbeiC4cG1eQE0+GLq1nR3sx6zdGTIo8YVfKYwdOkG5CnrAsbK
OmpctF6qwLNONFFPbDyCmgCU17aGpTAYCYKn/T+q1dSB2ahBx6o9BsbAFEreNRgE
5FprCe4H2NOvhJky/jHJSJrWTfoRMNp8xZyuTs36Td7S2rud7xVJcVJBmugPA5Hq
tAz+d74KL7HIOFOeBjhBys2vDBubP0fh9RaaZxOHfkhKhbGd4hBH+8lKnFjrraxX
9imZ+zxLtwDjg+AmZLXnHgIHLGvWGKfq7zXyQJTZMYNzSgDaMnF9mEKJ5ArZaQ5v
pQtxJ2KuaPv9t7vQ4eD5Yq8x0A3BDPH4sWnGwUlkWgUxLOXfGFPJPw34oZugR5De
soAA82bSql0TyJqHNN1ryvaAga9zZhvNDFynNuBGL7RU8pryM8JgexOTweUTEZhM
AZCHTvFnjwesPPfcbQBY+2QELm+iqxPG5MD96XfS2wAE/HDdGkgWS/gGoj4kWB9f
TrtpS7pqEKyXatCC1+MoxJ5TMXg2extv6jcysQLbU2L3/yx9vFGXyMoK+1Epx0SX
P0pzDoQQi34cnml6/ID8pcUNvZizrLWLa7ehp+RV1BE/DSLG0X/7TG+DRwc+MIX7
2VQikM/v7Bw2vgTFlMFTEwn/m3DN/SNvZTo+wvvAfBwrvYvJg0v1uvI3Kbbi97qS
kpTMvkGUR+zXogomf149E5IeNYI2h33M2+8bJEwlmEHg1zWfz/xAvg7ifFYA8VO+
hCEuYeTo4sPtMei9Q+1XZ4a5sHDEEwMXo/CXtCX8jVINt+kA7TdUx4Nq/fJNBCjL
rfauKfT504G3/C6b9OeJyrHeoBwGB8QSaY8UgH1UGOwuSKEkqiMxGHi5UOqzsgN7
uQyRvf6enGPgfmSIgDBFd0nIx20l6f7qBivpJzKxGEVYmutDWCycsDeo/4nlV7kI
SVA+bNEK6BAmlUlVAfMiRMBBQCtr3Qq9sVdXKhyowQuTrwr/lO4q0keJe3ect1vN
5STwboR+HcsyfbJJnO82LnCPerBzIzc4sxzwTY2e1SVN8w6Hiu6rYMVkEV6uKUVs
OfyfqSiwJQmWXsirQOYYO0bYcHeSDpXqVOxLgeVuftTv1JJeMTu2igTeMma7SkNm
/MIJIQT8eKI0pVhCO1AmOvcK2DGckJ61SgAachyKzyt3FXfvigBOKWcdNPcXdp3I
41UfsOAQ7D9oym3Y7kdj+iiHe4ZwiMZ/BBFD1RTCoe1QAdNOYXFB3d8LfQW62lDf
qt7KJjqZFsu0C033bcYbZanBn6SXOpYxomthFD0T+EGghbMi+kpKN5FLxhzoOD3a
xRflwdmBjfsp39B3IlXyc9RV4vPCx+w3uwF9X2bVs6TElMQxEL51zPV20puANt0T
Yjpqp5AunpZfhMsFkM3efpGPnl+sbnDxbeXnd6/F6xCVy71zb8ZLKjlbbgbz1cd/
OxkamuIk+cJa1izs8lEmrsz52aBOrLSLbLiK1fa4uvkkCPCO0n8Rw4q6b0kcT4uj
mqhJNDIqTcWG1KckrIVPLa/Uf6JgTJuvQUyA+c8WBSrLpvx3alvMn60vllI0IOuY
86eWsTlmtVsZ5qLn0KIgI7/ms/VzgjkYt0JOSxsqMwbrSKaRkKvrCSQeT1fH7YaY
eJkuKz06JZcApCk2dMKB15DBVVenttixplbJv35CeYSHpG001TJuW4a2lEapjg+K
39IPMPRG6RQhmvRP3AQFPXNv6lKxsin6tGFxV2R5CbKTUfMMB+1oZMSFrYhGZySB
3naDKhBN5EGl0AENDwVdo3x21fvpzEboGWVcZdS36yaLOMabkGEUMGbxvsAeWzad
D5531JwFVPUiaKknQJF0YNkH5c9LuzlLuiO+rC6+C1aeF8PKmkZvig0aAtHCuPjS
IqfB6JQ1tb+62uIBPsuKgceupP7ziit9thOIMxjBdQ7Nl6cnQKXhhHHfi6OSq9tu
F6RLQB7YJiTBgYy9wnSSfhbHb2vYtaiZ0CuwdxgaG9j4/Re6KA30d4QENMYYlip8
htQ9psnfYYPn414gh8MSPibNIFUdXBVAyMcoaiqpIIrClajYF4JJ8tklYReAePc0
bzoUSMV9qDCOgqMF4KIEVo/kqJJa5xJAFbrORxQr7PwE5EE9GC1Ll7PZ+5HUDzSa
MyhiRosPsCDFC+BI/kSiKLZlJrR5NbgswSUjm8CClBpDVUBjiflZrfzv7pxda121
RgngxR7RsrnxqCmwM9hcxz5N+rdl5X8dovjrTqcfv7mXslPPEcpL4TSTL7R9P7O4
R8pvGmDuKHFVT/XRPxxulSN13d+LUUcITxOWex4YiVj0z1VL1g2WB6ZWthKYg+2c
K8exeTQUY7tQI1DqFOt6KiRN07mWruf4Lw1ZjdY4/41o4eXlWq2axFqDbCO6gi1d
6V6ZMzIWqkFTppbuT48gWunpeKEcxaiCkbE2iO7HYVlvzyy6lzC1lRuT9s/6Jt9v
xHc8qXXTaOnLfa1BpUrE+GF0Y6g7pFe7q4Z7uTNAMzNTTHBlwhQglBEVIBc0NR+e
5SHjbHxGvntpLtKYrYBODVMQo5t8xiDkxmCIr8n1DEADymJDaJqyouSmweP39ZvY
eNQV0RkLQehkf4Q41pxHw1UmcTjuEL4fBi4629NqX8qhIh0ujrGOWbHtYglU9rc7
SprNJL2Jn57v99ZSnHebWzCz03j5D17uVCMAr+4asP9lFkJFJZ9qt0/I1xD/viPi
Y/zUaT6EwPdDwtPgwfd5N0F9c2x7TSwS3EemisrXhLTISQmU9lDzONNWHG+fq4RL
U5L6XNTQE/kV3tmjp3vn/Q/VuvcQQnUHovQXnHEfB4a+dF7tkA8ksSR/ApDXfejT
kEDirXVOfSxVIN9A7SlklIw5zDpfw8aTHplR1uMuoXeGFMdEgzfdztdvFKEch2qi
3JeAIR0LFDBCUW8aX0TEAfYXKnwl/8XSse7ub9e3q8VTZDUHosRGCLLx0pr5NAYt
fufQG5rtq+Oaoh6x788Q+Q1aHwY1/LePmZ/+DkN2nUlqKY+Mlw4JSS0nQu8x/cp+
1G6BElWgiLkNkvwXjiwHzbOz9hN4OBcVXS3OC2x3gQea+Oo1QaIv7gmkA/z7Ib8f
8LX57/KfjG5wUDruZBuWSrolIeUvPZB0phovwpaOx9DXpt6aM7DjZxPIbSy++LQ1
j0YwKCTbzN/c3y50k4hUBDCmhVErze1QOWTyYXtlG5q/b1zFDzJHUnk27bl+2yuB
KQDQdG//rK+NeMV70KVjgDaPgz3sI+eSBLk8eRKZnu98LKQWT0wNhk9zMIZZoyN+
FWqc610YDAFwKfKEVRIzGNq04A6IPsPjDL0+G2Yhf33qjEV54OXvYX4TW3DL/Ec5
XA4YwQiiRZnYoLRJZTg0UPmtiha+JmlFAoOCVod1WJQ1TPXUx+NVmAXxFJD+I/6u
rFQBpI8tKx2YamW1txiCe4V+ZH/jMr5kZ8dwlJBJmlUyVCHGM4abpaVht4rE0t4b
pvASdCea//FXuc5QzXp5Ie4o5O6zWWzF0fnA/2FNRcsmjZeHUrxvlvnNqEVyY05/
/e/GejEpT5d8SI4FT/Hgovh4Yx8VaY8WpUuFZvhsoMPDDS8ofFRDQ+RNVop5UxUp
7+RwSamxEdG11xdzD0VtkrgIwX01DuxijFoq5xk+cZBRBoYwKsFrSfXdNMjIdk9M
JqTEqGhPHz+X1Xuhk4A5Zf+GDuyPDcNoPGj1coCWaa0lv6HnN+H4zfXwa2u/URgo
zUAo8KT0R1L9iMPDJmR5wUK1/v0ell0czOPvZy7JdQKrZ5hej7CQnOtio9gVVrHz
bcLtt5eUguUcvkCCfVLhTIzqREd4AxCWztGRgYSWRHEUvpIElp9qezIJYSKaPGwb
5ZTKgnp385kx/yy5tvRjjkyeueF5luZ1cSVuI0V4Wx+g0XhP12G6aabrGIaMMydQ
m+CjQb6+SjoLcPfEm3ovKCAylK0CUalQwyBGNigMLCsUKr6pMneMczJ/i1zIof0z
B6jiz96SYld3FNYiDgiMCsMqrYNvK4LPNw//unIFRGOGNQJxzAvDQNPSE9l7woxk
/wfGSFeQAmUVmaUI0QAzLOFywoxTqd+D8MEnB6FTTxop3dEgza3xHpOPjIdu4iB6
ky84Curj8ccQ+H/VwH04gUEU5jTjQTk2OQ3JF/G5ur0tAUbL+bcgGFAR0fU8W24b
btI57hplGvbLOGk0bwzGG7fGdW+pMfkA1rucJAHgLZBaUxgWdji3NKJHP97xW5fB
ugb3sJmfHTEPtDc5h+L+mBdNtMTtC4HitwALE0I0hNTExDzCZZ6b3j1TTX7gL9an
hlJEAykB6IjncLLopg5h9UVpHXNYZYaXpoaj6cXhPmBiNHmnjdE+VWyg1KCcdQlj
dLeBk4+iQswXMEEE5j3go2lvNxJOX70lD6uxWW2ogmpXKiC7QFd+IAQdERoNlJ7h
sxJKEFfhX9krwcSFTw0HcuOT4YMKl7pzMpfxxYttQKnfDZol1kXzDvNDJmNZ0GYu
kVke/ahov2MFaWUG2Xp0qpvbyBDEMPVklcwgHmvFHyNvS5D8LMvqaAnZ3mztqQtW
E3Ob++n06C2ujIjApPaukL2zdUxchJ1NjCRg/67T5eFT7rcXQGB6PwZph7pHWTRo
mRyMZXFC6G9wuLvpoV7NHL8pZNFRTinOznpJcDAFopVo2nVTaZtmJmOI9fIDQW0Y
8pxwHg/7jTG3yDXMus7y0WCTMxg7X0a8LDQzUeZiZjVxV8C/VdGCaT4YoSYBAO2L
A/9KFdBAIRFlbIZakrkxtGm7DWTv0vBXMm0pI9sDAhnx3YiymEKQvdGPuQqhDSHb
fiQvitO/XiTCcZKy9CapY0N8WlXn8tfuqsWW044gNHWUYycm1LtTgn7EybGEv3Wt
exi68DXKtJYV2KGgPr/BUBuBK9wNsFed3XUNoxysakpqC/NVM/4f8KR65h68AQSx
ZfiDlFX8UudxjSqLwjYgXhjujqBzZ0nPV/NVyUKk9uHSM8OozlLxdO7H/6mtY3Kb
b9n9nzN9fbyYfp7aV8reeHOz+N3KlwbFMR2jGwRrBtERtuUHwbxHz7agFIONp9CP
mYgi5YRpVWL7GHaSDpjCraDNRmkk6dTPjYOJjye6WFIzRr8BuDTF8mV7+aJG2NFN
9mcmwetX2e5nm5CCuM/m5XTgT9N1cDzSnOVEVe6WAEn5Tx49cYSDzeeOL1KyF2Rd
eXUjeW1RzLXtC6KVuZAZxTMgNVQ+63+ZcHvm2oXbek+TvK8CuF7jlp4K/5QdEkkV
Z8x5rQR/jN9BCyDNkocRIuGkV9Rx14Mzw3Orii5YYE/oUvv+0Zs2aoadg4Lhswau
9Q9Be6oRsXt3xQ25o9aUF10qdGKpTVq7snp87vvc72i5sTBS6Gy1nXmqMrtT/sxJ
jEcvNttOhdXZIhBVjG+bsedQhk44eLLJLgxO+VoXhaWW2JTqkAeYky78OdYtJimR
T2b7F/QZnONZk0nGo3yMV6uOzYumryOMZTq5aUsYl3rzkeoUmoYKfBWZKyajdskk
oYBQnDg02Aq+wDousaJsI0KdlNGklNBRsIwbhARVfh1CH8hN06CiT1bZ13cJGi89
u3B9IbvqMRLuTJR20K1hJKF3gSprL73YF82b+An4vGokrb50anKYVUdEownfOzeM
ac5xgIw9uDJMG4ihxIzNybOZgwf36UhdKCeUXPjZ/oUCmf+v6JaNLVge2rf0zziN
KvNPvCziAkziV6QZ4R4vSNMCsEqnL7l72NHR2R2JltW7t+1uyU0KmHB33DE8hFS7
R9b0lwQO41xq88GzLK03DI7RLHVVum1Ex9jvQNm71mzjKKIw08Rjfg4DJgNhysi3
cvgrcDpVwLKH9Q7uRmYFH0x70oFgrLvLHo+OI6G/+HDUKopm3/Syt2Z+hhQUAWoW
LfSqtkm0npdz7nbMj9fbLe8UVw7R12H0S+w0XDJCoxGSJvpatOSHQ3aNPMiKgVkB
tLBUOJWacxZFfRxJxNgwXmkpugEpY4zEZcVxCUPZUbBMs9KBaUqHntqEhVhvnv/G
wEpVBkXGpQdYLw4CrqSMClnnivG2NqLvM41SbJEh5CUcytIuIZuG5lxznQJdEcqm
R6rvJX2L2nt6tm+cyLDuyZR0CBKdehODgJRyd066vn2A3x0GWA74cXoMc3m1mpTq
BpehtVm31+IwaWS3VeZ4EvLzMVPvkQY01L0gQZkVMp+gPFZXAXXgil3VnahJ7D/X
lPm+zVOJIg99AM4YZsvptgtJKuEh6UgLO1SXcrsoG8CsCKUpINN7u8tFHSfXBMfC
9mdLi6KJsz7j+KO9yAol3H2ZWdiXbSb9fMh0Kfn3LhHfFyDmTJiUEU2bHCawoghh
FGjJTczHMegB6LlPjtuBVoo1fWOCerOWTqmOKe8g3FDROngXIjgDLWYW+qRmwwrK
TQ8GVU7CsQh1HXMRDzKOKJdP8YhpnJZ6XKsy+RQK++lDs971lvDNVYNJaf5aqflS
SZed7oV9vfXPufzG9DiCERmxSDQbIsRLuV64qHpoRh2zwDZzKLxqNNkPbcKh4khA
45U/53QemtdQm3Xn82ZRoxF8ek1qn02kQidIYBaMtVVlSQ8qfWooQPAHTORtcQ9o
BB5mXwQ5n1Yt/Wk8++6yAzlpGSO727x9U+MD+gKjyBHCb88kBJK1wHQpRpfZT1pX
ndhhbSqvHl0vATCYPogmGBgNR22hkp8Rd3jgdla1skGyR9qoZ0AGEYtgppw3FEyt
qgFb9ATf2Qin5ldyLeBRwal4+XFygH08QW76ZmCMMY3gfmLwgC+767OdfNFX8vof
UYFpEbVk8w6EHoA8BHi48yvW64tuOSmo2ae+hI+tAiElQSbOj/cVZdacYzVzJCSR
Mmrlexg3TFQtnP0vCyYxeG3sX6fQnbjnOEt9vbYFh0MXBdo3a5afPmJxdTIeszPA
bRHfqbJCsbNbCr/AzGU6lwMWhYUqKsWuB4PAk6jNT8Bxai3h7ur+5Gkw37R1Rw5s
UCByqLFRjeSn/eQk8/7mYGkZSAAbDWUZ+bUA1FGY2wQZ+gTKMwwBCLgiuWBHYNUI
GwKDo6Q4i+LQ8kQCqYJGEI88OlRT91clAxyvDd+IKXJkNPAkd0Vz6H22tHAoSz8P
jS48MmOI4AX14U++JXDQT3t7ABtyZT/ESt/bzOXcA4Yn0y2d59XxfUBzL+n1PNbm
f9T/OmPp4K5BKYvO5a9EXdrC9/E2BGZHkKrixJFlMCFrYQzqSxRkx7CcBllItlP2
UbBEDIickJjhop/xQJrdEmXPStBAjvuorNZFYkqUZl8RkUrGA7WYzt8bNqPoPC0R
yfatosNyIDcEdRoTQHAdv19/SnAwU1O7GAVfg06WLUyx5InDPGK36bdGPEDVSgaO
cPgPxWanjm+kEf3y8FQ5uCKhvLhvOqjBZVf6bcVGb8Qq31HzEqRxXcG79guBGzFn
4F9VbwIqQfcV5kuYZUPXE6cJuyNOGZMiQshDcajj4gfW+plmVeKepspL2x7enH9d
1ScOtGSRyG7PycmtmxukfAUFUq8i1FkWK/IXyS6My7AuTIoKaCvJ51L9s0c6G2Sp
mdl1k54Doq5z/FT3A6HMXfIWb/89tomF2NI7S2NHqc1mLFm3rwVGyTKlpIIaoW1X
aCFplfcGfm+PEQ5j/VZGa8YHxxccMXLEBWRm+7Amv6w1T9PVKcHeVwFxCw4roklA
BknMVwHFF8kTjqACMooDTnzKjsqM+AckXgAyWHkoSYTHDbNaIv8pjJu6eZp0+E0W
ttWP5V7cmQfKjW1dg31DQDtPfPHrulHYdwiuhDjJhnWxgy0DHTR3IOuFpqzl2GCD
RKJ5b1o1XwhJzYX8ovCStG6gbFmcg1py0K25PjCyiE27xYrMtwoT/wdFtxrHUiT2
Dbk3ekYy/hoSYehza17GnCLSq9D9OSMITWB2wpeIlsTtbzrfQfkcXNoMIUicbMN1
4XTvL2I7gyZl1+mJ8BBuLKruOkKXXQIAU6BcuMxmtgCowI4yXVpJYZ52gNvhWkgg
Bq+pwiyy8B1xA2xekDX10CbVdb8erl6UDU71/YNPHhO8r1d2kKBsS+2ZUrNcfD5q
S30B/E4HRJHlQIW9aYrg8ooaxHe4cl4vmMkshoKK+PnBnuI9rYJODfL+OBwrZSCo
st0Z1hSOP30/ybHoY8fVjD/v89H2wZfJPP2u4ao3pWdbjZOKtPcnvThDWsV8qcka
14BT9CaiiNcs1loAKNUujU+2sDVMzWW4lNpGbMVOnfKxlWDdH+gCDIS2YrZ63F0q
BrTcdGqNLodM9rNw4zv2WQ1/PvEe5zCVEdWn/9wmwVXBSufqmgjVdvy1GKBhIiUJ
XJnfVACsF+7foUmtgMOHC+kqBpNiWj5NIkt51vqciML4lH1CtedV3UrgaTtFwEg+
ugzvT3XIDxNDikkvPYeJziT1ByH1EwJif0eKvOjC8cPTj0grgYOEJVSxdtE/oXgU
sP7KymV4QanBULSns1oeqUR4SddTUYUqUNxADKHUSWxgLwLPXf+VMzL1AtV7sZk5
GLmYnhtlGxHEbBkEFb90qfva/C4n2EmIg3W11rw8EzNXIDwNWIu8jbFZIydCDEMz
CFFyP32u5oun+RUIefNk6PrkxPP/bnn7iANASX/RnufOy0rITJ3NCYvjqVv4UpJ9
9em+WbdpOYq0JzSxjphfwXw1hZoMUyvGECNUMaAJx4oXukL9wJels1tWgQ4JvfX7
mAlfDUWTy2kk/jzzXJMliB7uGfyHxahR+9dBhN1NxFeoQK98sNchkFgxpUiE2zGU
wtbKo0b1M4oAVEWxr+VOcCTj6SDzwJBiIIcUL5sOhuOSW2QaDBGhCxtoaOo7r63Z
xq8liOU+oFGt3Cfj8c+7msBgr+aK9O8+iyyQyFPGwK3NzQczBbcCwh1iJJYSSOQs
0RU1A+dTrchd9tU+BmjVca6wXdgx/PPHHc8tgbXxEK6oKPpBueL3b8lQGvA/kVlM
cukHkSZ+m28nW9PlCPUVCJOjYiOKziEGvqdI9oOjcvUTC+KGVrDnCUTSeTei1Z8A
vXnb2Yy/yc7QxXVc7/5I0xnqYhRSH9gvVaDeiapx2LsksOtjxt2l+7H/FJZvSU8Y
GcPykGQwc8NLn3AtzStmHYBuQYhRfYJl3jRY6Z55g5EEW4rmEAoFNgL6UeNoLJFh
m4EYvLIa53YZiCF44MVQx0u9nJcxXYeOyckVm6Wf8whFqxfzougJK6gLbk7Pq8cX
y+D1IP5ZXlmgmw6m+B2nvEhYf5GzR6bleA/uKecgLWFnTRJG3kx5wORKRKo5VxM8
Tgetu+pNyJ5QK2lAD7W1KuBZCACL4PcRllBzQxceKj8FfbCpe1fFdj5BwGZ42tcl
UcRClk0IBv/hCo4Ep5B3Bmdd1y+mVzRbUv/7+VaRJTXSRh7IVV7Mgfg0Nl1JLm6f
e8fyBC55tf3ftbARYkc8+hDPYeVmafikdfYASXvsSUb9hu/uQfGDpuau6LE7dWfl
tndF0GNattQKLNLsWs/Tb4jn2ITEjYhcZKTDDrmJhe60FjLF3KiGkbKeAwqfnhEj
pYMd4jSDNATJSfVTMR4Cg6FSVrrYIagQ9geDpOopROXxJ/M0QlAZcbP2kCBU8+2F
gpL22zg7wZrxlmfw8r7SjhD7CP3aFQoDbchKXExTIfigy76ZKmEI/VHdKyWq6ZrA
T+9gjtGrrYyTCanLU9uDKAnzRc2OnFQr0MReU5VE95COfcTPcCGAmzWuFzOHJOlJ
NBCVTrMR30eHbENgDuRpQgY/0QNIGtoZfTDd8lclGhtaBB3BZgEhnZU3ee8aicWJ
cu/qAWC89FAhC3dps8mA5MhovzEWKBVK269H087NB346PQ8REGOVQgxWQMGgs4w3
Up8Of0zmCpNWbrYCuZFGQeEJ/XMsDVdDpGy2Twqb9zjXSR8fybGF7FJBwRuI9xrZ
kulToAXk0LctmDJwElyeoVxKiytAhGcXYBeZC2hOQUmPSWFSinbT4eq+KnKavLr0
Ku2snqgy58vmhUFmO4bgfuy9dlxXgp9wNqQbFZtp6ZLYSbHfyp973ZOfo40nuolm
cNkNq7DKiUmSgdi4flrN+ktkBkdO0g5vYVdpv7t5oLdElEiwAwk95iGLv4k6Dzg5
7Br7l5VLIcZrCOBAejdsXvY9BsFal7W//JV1/mMfcrOWJAYbXSEsSmzSsgun8hWc
gUuWiySrWyQGAOlyp/YJhlWL0UpWDzbhMlM7taZeQCjsKZ16L18DexQ/vtMzFD7V
zdjDqQTP6d95ZZyRl2TQ4z2+w4egRkMgO3JCffEWXWvuJcBSi+cxp1fI7Jjj7SX7
H6zTdz/zIwl6Sc3zDFxlxAmG4NxFwJhIM+OBvbFQ4Z2EcDd+qq6UyxY3Wyz0KnbW
lMvuDEfZ6YOV5uPNg8MrR0lFQV6V0BXZSyXCKAwDQtxl8Z1u1pQJ917P/tuEATZa
9Q60mZrXDm5fdOVKF3P9QCnL1mRAc06YjT6wBtdNnMlbrrKwWBK/7r2kJPluqvtA
dyDtsErjqxu3IPHKJaRk1AFHF3IH9b3Y3KRji3J+VbZkfEnOa16BXNHgpVmudZ8f
Oflv2IbmBRU/DQV2Yj7PISx6Zx530w56Vtt+Ugie2e4nIk/zqb5OpvBaqsILcWXs
mfrWlYleQlJi7VQfgsJUpUNMb8uJDVfCKyKVjge+iyrVvSO7LvZSjFh04U8hPy16
NBREIbafwY1Hz3b6Mdt3Q9c18zfuuVRv6kuUyoA/ad+ClUJmnJR+HQzDwcRplalP
kkeNGaPlihAmJvCuU5QOM5EVWXL9iBQvwhgYj3FUMgjptBwl1fJ3HB8MgS98vGBf
YOZjCpAfO/ZhNctMkyr+X76SpSWrZl4M0w5ajkacxOYmVDTOehp7rL5GIs3tPYbl
b6jLHlmx3YzcbTNgFkJKggKEr9gpimHV6LTprcUPvGHLLGx6LC+vMl4cnG45ihPD
RPVFxyqsVeay5jzk2sjVwLDAW26sMv0LnqTanjgV72JQXgpdNndFETgwJHKQm9/3
lk4nkjXJXXrESgRxM0TH1EkCgQK28rzm0GTCgzC66/XohNsqGz8SV1IJzx19oV/v
66atwG0/A8tJz04yvI60JNnFR+quarxnQV3lOelxB5/G19xXHs9lrojQYVIBC45T
mTsykLAvP4gutmVy5YgoFCzsHZ3lU1PNs5k66ekOPZdLzIJCyu9cXoqXH/2/G5fE
giaZNs6zXz8lc4vBt3lYlIWrj2HgGvusP2cN4TEZuBGop40bMHaMuf6NxQpA/vEd
y5TG7HLfOlReHnA9/0BDSA3YJd+xnUN9QIhxz8976rJ9vzTduVCdp9ycu4KZy4Au
IAm+bGSGNtkDOsGy2YhOLuM/L7pDRP56HyXs0ir6goDL26li5hPfOLo8myUsQ+Lf
SDpBFz/DCapzmp96XzE1l2vYrau6x+uWjrhVxy+Ed0+eDoRlw/5IWKmsow/21FUD
Iu4nSmQ6Z4NpvMYfHNDcuu8Jcug1IkZVxByhmRcx6bNS4CV40EtlsO22BHBRb67y
LVnPLNOQITyJ7CzJX5NEFRoUfchzU3GEaWS2Qe9qv5lDoASgk4bMglonHsdE0rCy
AsJjnqAmGxyM4d8YRYkHR96/b7ZaTg7ol+EGoxRLbP1OFpQXNhNtB0BeP+lnCXzl
cFdEW5SzLEYnKl6Xd4aznvv/kr/PrBEyI+ELlUb78/z2DafNUS3DUua3L58XlO7u
9U5xc7eqdWwzwk8rIZlkcTcLSzNO3xjsnDxlXOt+Zw71/sgPibQYvPO9ybV7u2ii
5Ax4/Rwxp5U3nsLjGoK+nCCoo8x6B35rtentwt+oFpeQnPwz7RFE723Q8oO3W7n7
rbL8XmBxG/riBG2ykjCqidDVWLaNhvINu2Rsjfd3HRX40YCYL7JrZw0J8SdUawpj
eBjvzHmJuzxDzyHVsEPJhA8bhv/n7oKdj/lnLPqWKqTUnI5B8NLdBqSdMzADW8jm
KMD0CE7Vm6X9s5/aNSmfgWj1iJPHoPpR3SP2clMyCBtlJW7CIx8+I1pHuOlNtTXV
8tHSeK6QbS+MYDfhvYL6DLv8JR9wYsgLNWUnQB8NgJPSw/wzffdNuXAK81iAI5nH
ILa180HyeInNCubTyrc4vKJWENFXAHWvlixKWUDIuxPvzKz4VLyOI6p6fC62ZwRZ
W01exS4GHLg0Nfaqa3PA5TGLgK6WT7jfD13awxVoCoOfSk9Pt+7Or38ZhTBVLDXA
xM29ES7OYmVrliutnpWxHFWuPOfpSOe5n6vsDWI5RjcFIrWLHY9mho+xaVN3aJ1M
RE3i1mwglyaseM/CtSHy3Z8p+4RDU9hbFoifxQc0vE55XqG981YQLz/HSz2Q3oBb
aq6V2jxq16sfmTyBosN93gGaRXsX5HPFFCn+Ws/+SlC17GAW2TrXMkMaVsG1Yi+N
QjVh2IfjQ/bJRovWuGdCvWZd/S85la1/cT7QgXzL2iw7JR1h8c/DytUa4W6881rx
N8CKUk3llbUbPkryOn2EL3Nco9Qy9pPpD84+RjO+Fz6SZpRYq3ys57hRx8ATno6H
UON/ZcShhN5su6WNixO8+MBUWpyV1ievO0KjL1ut37Bj/2H/+NTXWuQ++0cO1Bx8
fa3DRzvYykDm/JldfwhC0RnaQvZFkqPZ3iBj9HU8OTLO5BgB576C5JUn4AGmg3Vu
ifmC82qiSBHg3qtFr0oi3nRZ1oqfLkK6wri9ulXWpPwFeJZVc2KoRztDOD3HGnd4
M/PLZvdG2k9LCNNARorcU4HsjpDWthBBHUE4+yCY6soTS5X03uWKyh5uyZ06uB0y
Z1T6qmNS5lwW72xp8Anl5Lra1ZVy7ajQ6OMjO3C/WD4nJKiizNb2qTp1CqavxcoH
/rjx2Tu7nj1R8wJBqYpic7Wqw956/SGbCn9YCfgHOaumk7Iqa96wFd0obEQ/HywW
yEZCgfTWaaRGXEzjPVjI0Gafe2NSwG61phGE666ynoxXPywHuKjTnSWdG72Oklns
fcVoHuYDiEv5S4TrOVjnCWNDpfFGQtttoO9nJbuUHd4iSN+H5fC/d4CE44F5qZb8
dwbnEnV4VOKM29kS76/VMcs9oQ7YvXj2DRnbtH6oxsyD8Ki5JkHwxZEAe4xc/Oi0
kU/HgpjIXtcTA5yZdzdPfHx9nvJNiX1pDoE4Qj0AgjW478KcurtMb7yQZgjpEElr
Ez/rFWvk2JHHhJzhSPkmRYcynu+5pRJcc5nQsJ3Lbvn6I03fE5MFJEEkbIE/buvm
PnuBnV/Q8Z+dSiVnT50vWQqrVXhVVlhXrBXuIS0tvI/4t4Cw2fSSYL+Zi7XIxZNT
7paDZ4mBfxWkX0te1Yk3YL79R9INMNrKNYNIds+sC1HPCLuZX3TbtTmizWW7m5v5
SceVMCO29mADj0nDAtdAMSrpBL9fHidEh5ayiOd3u/ED3hxhOWs5lTJLX8d4GUjt
5ImPe/aeceBn0BuY6JAnYDDrEXLDW6dfXRXcrTT5CiurKFX78dpKtCoe8FyfL7yV
9vTr3bbarsJfl6yNYZIpCbyn6kD0+EeVNu/uPzLeRFoyq7FgXJK0CBoUFuRXzXeP
PZ9p5oTyke/AZt1rwk+zoNtePSEYhQxcxzK83LtnTsrikRCWWI8xgBGdXnYmDV1x
+RDCET4TtXeVhCfZkfI/BDwvqc9dOEG2m8wH5LfE3izFcBwUkFybjilIxaQGCW3j
tPsPy91AEDqzaD7JD1CyVIc9REmAeZVqxXOLoZOKhFZjkt5TMXv+iToDr+hd5VR0
0c6KzdGfxRTI4msbgDMbiHrzRVbfIEGuuMgRrLIZ6ELcEmIpQqvA31XFapNyWWBu
cYoo0/GgogqzGO7eFtHK6H/KcqaOnkvQZkzDkHwQ4i7jNawhZcFiMQjfnuzg6W1I
L42n1/tC8D5AgdP0Ew8UWhqOoUe1Amkf4ny6FtwYNykw2glRHEQjdXSpLkO/XGgV
crG1fHajewMqVkG/oevQHWmk+CNKqWp5EhzqaJcwBflPhD1aoLSsJ2TyztM1Kd3J
t3fdb72rH+qSL9nsCnR6diAGQ6J6smpepVTRtIoZUgiOTLV829pA5ND973XdwaQn
JrfdvOprxnFWIpY2fa48Q982Bwd2ru0jbbyoFocEmhb5ltJQctOOjZqKScToHuJd
NgTPDH6kL0VsBhJ0Ag7wHHx5p/aE500GOl0ad1IUxszMuBoEVuZ38kfPFNdHF4/b
y1m7N6kpqkph7CQr6Ta/dQO1XsYXymJ/NLz/EyTs4nvf6FHZOw71/6df3Q4JRB20
ueDu3En7h+LvXFtyW3fqDAvOStHr4wTSNp+jvFJPJsad3zZRNMYVZiLnBV4Fl426
M7dYYkvXX59gjab4AwbskYCXhs9DxE+9ZfX/zQkFxSS2ej6NLgpqn5Z8arpJ9Tdt
T8X89UyZ2/hNF8LbXvzrRCO/qpQ+vEcFAHRtjQKGyZko1SjsWxTskmEEXKW790qR
k3BZpe5yIRI9nnUUDbrvummddIQomXTjEDAXN1Z+n6kPsmdtWnNdXKyyF1FS6r9r
jQIaTrnXlevutgGNumMVvDCESlO96hl8UANJ2xb5eZYybapf6dsCADTDEsSCPHkS
ch8UgUNZLVPr3FPWitg1TJcIKbKANhknL/TRJW22k803lVxvNWNUZcccreLDwz/J
seAEymU0QGP+h6TYFxNmOVl/DGEYeguMpNc0Nfxhdw917lWPeL+AyavAfTngYLo8
3+8WrgXzC+wOoa3kUW8cnihZegj9/e8MJTEgE+Yz9AEOexeBJkWObdByCMMaOYCN
kCzzfPb0vaCXX8a/1aSocQ87gYOuOT4X7DvkooN5UVB74MwRAMtSzRGtCq4/WKij
b5jD93unHDbECv9MQZtG36QrE1JDBfr6zMlxFczIzEs5y7VT3YFJr7kK6gDWG5DL
332olLvrXWBy74jbt1EARvYD7hPy791YohNuHhepMIdmDKZqmPyIWjcehcNm7zbK
Tss5NfYxPwxAMiH15CumKVHiQ9RBRyj1PAifdPx7A6tsjuYNv4FQExxsv41Xl7dT
/YxQ1MEzzVL09rKNLB7LEYLcBFFLwKchQPNQj5QIZqIAts8s0VysrFn18pou9uI7
8oquY4zDaXZD0VkxRmRKAt2D4FoIE4kVjlhMZKVOV68X0/a6pvKMY71HnlHDDniz
BToDqPhUcjE/sY7tlocogrqZW4zh72qmWGqgl6CNeim8gwRBpeEsKiH66PXd3JeK
UF/W9vPKkm92ngAVrLIg2UteGxFR2Lz61NXNK6EqMgBB50HA0e7UujDL7U2EPRVJ
B4422M6pekBklp2BBQKZ3DCgSNSyNUiudm7zurthMdophuYhu8Q/My0SlabqPatj
quEMJvg7vRPYsIIDI1k9sWYHCK+OgnNPvAt6pKL9jr20c/hxyMTPcwEnfQgriqaY
0jI0g4ipi01nfgRBZyAuytl6dePnYEPZoSp+qPH/cuhQwJLZbhc/NDGDpJlplekc
8NZ4WvfY3Jq+iMvA/E4i0V6SoAbaQYFLRcWPIh2lQjJH917uynGOrtba7IChvIco
f7muz+pM0nEvgfQoUJV8hc6l35z11H+hy+9lBnWK2lZh1kRrBG0iN9mOKPkCDfEI
K8A+R/pF9Q6phBRYvJAKlR4jx7L23KRnB2+WmRRp3ESZGses18fkgnB+rdOzh1E2
81VGb5Dx4ZbGwrWkzNVvhNZJtGRX5M5xT1q3BKBtlC7NOv08rGrqjqz9Pgdc9INJ
JH4qFXKNm3JKtw4nUnre0rXfHNo/o+ThRoyJlSp+IwLOUTp3+V9hsiiki3fzYRrt
ovrTKVwFn+3BlJfA2eBuiiELRKixs2VxXytTD0tjlexoZhQiCGXZ43i95/nf4COS
Qj/M+gAUKQ90E341ZKDXORgHW5IOF+CHdqaiIj06ASCJ8V88OHjZMH9dlzeX5uGZ
3iQ2xdNdiyGNjkEUhAdWLtgK51uXiGW8GUGo6JHFBW62k9MPjWyXZ7PNXRhqceVK
k/TL6KOo3LmOCQlmtKJXuVrf2jnfs25xXDXlgr/C0ShqIsr7BjxbqONuyGEdDtan
VrunqGukDmwFU6aa11Vm69zZ/OLU9ml7t+ruaIF3cPxA8GjnQ2NfiNAEJNzaPQnP
k+SHo2Lit1LZ4gQHJ0j+5PJ3NLEzzlEukxfcSJTaHC4o8Cn9TPogupIMVD8HjnRJ
DLBEAT6IxlzracRh41HtwFHboayWq4bCmmaXl7kLvImFcfqW4RTtDvR99r6dcDok
c74HIChdbET7gzI7wUi7TNrtDRks/FozWbOn0gcW6NvuDjJ+BLpijo7v+xIa0yFe
BIUfqY1x2YIH54qDPQtKmMr+jXDeKoMwRfo4nnH9h9gAiw7vJchnZHa9HA9/WTHs
L7iD7spF+lBNEjx03haSa9EMY5XL6eeT37qlFBB/A99zb9oS2qyeeankMFTU1iqM
9ggcOUYbZxC5uBw9uIm4FesZaVEfB39ypSoyoAf+e1T2vCQfMa2yYtouhGfa2zCb
OjJD904OX5MVWosNulS9VWyUu2N3KsGTc+5h68amT9PKroA2uAmHSOPQ8ZRwaNy7
c8gLWDMP6RlmaZB0xHv6q8CYykzbJ5BNaAIN89wnvIV+N6NCweBGL6QDmlRMoI6H
aKWkGuya8DP0cMK+M88GaSV2ABYkFfsEpzmtP6O5sB4+pIcxE6HkDesV+YIryDjL
wUo2tqW4wr72RAvJ5atonAq84QAXxOcI8TPu9jG9d3A/KlyNaIHoxYBNp2XW08sM
JhGTUwXLHUv8EbXokUnhkT+AquISn13DR98M3tr2LP9bhZlryAFp9QJFerr7d5Sh
jbpIri4mxlYcp2/qXiS8fudRFXA8HAmAfg6hJgolYbdceaxy5YTqQQ9YkyyjX8ba
4Nqm9eO0+hw4PcRpkiYuVhCPW9f42ZYrr/aHCV3GOyRr1zypvmxxKDvNJ5n52RJR
cV/YC8dlWa4uFxnZzhlh8VTiXe7kaX9Vmbb93THcjhMMZ9DRSgavhCeLzBcv1nv6
gmOmSJfFsRw+/yUzqCNa8/aaKb/AeT377l/TP9h9VtdNdTHGoU1LI60JFxPZ/DFM
jfysD7nAyEorPJJuv5olBxnfht5Qxi+9GRoDtqMebqVd8Gvlg0dS3NsxfCMArjMw
siZVonMrc6lbjcv9vrlgf4iSrnBRxaUyhyz35Sm5SdSXGG6TRKmcJQVBKxb/tCP5
Sqv36c4QHTq+4emrCDtEkBX9sLSwOwFknecMtB85s6/KoPvkZ5yyd5IlbIb/RolA
+iOEdk5m8W6RgS7vdos1tPMqqD2kV5+xsNi2d9S9Tl0yqKVs8khPl8MBJ/c9Ynxd
GHTXqzbhsPLtun82UdovGRBzqJPrsLNaoOYJnN3AugltEA6mchK8YKctgVmJfBkC
kDARBqWjwwXFyKBJd00R+lxsgwTTKTQZyhXIb+4iV6tLPUBPJL+LuN7a8le7JmxA
EHUNRVJ4kWLb8F1F+TlXBa/qlJbwVhDHnKShY9zks+mcKPh/TpxxKI89sFUKfL20
jyjxM3oloHdnNr3yMpgUfpB30XhsZPqfeTAGNHaY+0KRdTVPGa2Q1k9SOZEo4QN8
JlZxiS2+40NO1D2uac/LkDoQRv5jz0tpljqs5aRzvrI1zNKvn1F6MRzm3iXMN7mM
rHJSbhrIFWnSwY0C1AYed6IT7bcthVmwCuK1iCYuq+sFyA0sO9pgDt7o5Z7leUUH
N2MTr/R/CcozaSGopQGsSbf/VdyvUyXK408Bk4ABYNh1JsHZUmu9B7UxN4Q2jPAT
q0Qp15x9zmVdZ3BnTJFJjRAVD9HFPbszQkiJ+tt1BnS54/B6vjudhV/4sI0hwV+M
cmCAC5QcHnvFAua4hFKqrkYFg4oLgOxtObNNBiADlY4XuAptpoWDZvCI+8hYc6Tt
Twa72tsk+oFuNPnHGE+geMnTreVU9HdUO5/TG537qcMti0/z39O1AV0E3Gh8Cw9c
EHPp7eu0jkgh1ttpa0X/A3Q6urIHxnWwRBAmkBCbMhEuPeNrSVzvSNbepo//5f32
tHS37GQli+jDDml6oPH37rVjX4Mos/ECmWQPcw+TuQ81OTP/si4iSp8j2qs+0Ymi
NDja1Lq2Uk78BWkMYKEiYV5ZBXnZZj+A/CveU0qNXrq1uwPiV5/gdymQN6OVeTAF
AzV9zoxE44AFf9Ineo32u17vfjNX+VLbxJtfd4CXb8L0fKQmq5uoqgCxjDRCp3sr
9W+Y6VqBIM6T3DgJKuCODEIOjjInFn44Lr413xMKl7pFy+zZLTZ6PHxQorotqfzJ
uPWF4tmyGi6gz3hh4hj4bS/E3UbvU5Q8KQiY2ywrKlB8glfj364I8DiJVYym+Lkd
12faXAdY1H/P39oWa3vAWmM0B0obApcMw2gsfmgXqL551I/Jgtce87ZvNSmC4IO4
vW5qdlla1y7f6IMvbYsg7Qz8bLsktiC5orkX9XUGbBQOr1kL95zAv2Q/Xk6csvhD
PskFVEaU0/V4cKeDPG7WGGZP6qTqXoouVPc8971lWXtKtB/ROq4YIWysgm7padMU
XFHNnWhTHW8EQqqYD1aMWT3heaztifVTG+N7Ilz76jvlKZiDJ4jVbyOOkTtrJBUM
R7bcYWfYYseMAp2hPBI5srAb0qz910aFrRn7GQQIo00kQrABSRUVTee23E/am0bO
c63/rrYYG6/054vTJnL2M+F7tuoAGfJxm85bERzxkC7a6sAf1eg3OUySpRpOyPZw
yv92sCbjOWepmbASqq4W5G8vtxPtSjZdiFrbPist+GTJ9304MLdh2t8XP++UAFLb
gCzBmc8X218ir0vdSA8Gh7jqop8/XTRjnRqYL9d3SescbwbWS1E85U+ElXiDl5dl
yJkL4O/0nHtg3ZpqCCYY13QnsTplD32qIyBUARIHvXBY8Ra5ERBRpESMVua+r34u
iqwJLk6SSovAejocT3UWbqNumzHBl3oOpXyS4zT2w/qS629Bxgz5T8NCKeusF3yQ
masxNNXN6Ibj9LpZrGohM6bMNucQHDhSmeIlRMm6Q0Sn7yntje91oDjosiSTP0xo
/7JpKB4on0JCCjSF+fVyZofucT2O8Ru8b7wY6p+n+nIkA62xhhuRF+Sens1qr3UA
MK5wHrE+V77rHBVGwAfvdCRXtJSwTooCjEkMQrkD2RgoNK+y55t5rBrCoQZv1n7K
nMs85yV6sRgdvVulB7SBNOM5MuacDoF4acSb7ErHEPwCvGhS+l2wR3uQ9zozbqBb
DcvyhE+kirKhpcSRj0fSeH4HT2wv1LjNW1pYV3oQCHvg0HNts4ZxhL+Rvd2ZkOBw
xOIpIUUmBb/KlQ52V6RhtzINfEHNNhBv8/przYSpHN4lbbGpq5hpvvpWvQgU99t/
+Phn9nfEit/R5kHKTEkbgKh+VXM6jBMVnEpPNy3+unbTf75FGQjvdFO8zlGHc3k0
U9np0ug2IPYddVmcLEhr7uehHlTHbG1AS5LGcrf383jYK2wYrkLE3Bo5zwdRXkxC
K3JDVI2PkJObQHPqHFb0anJc6g8lr5RXX3Bs+DN4oj6WuUh1KhS4pgiUADnL0/au
mXAunl3vtRQvLpY/ApUZ0jbWpicxdIcR34U4pWWMDQ/u6653JDzmEttU3+00gulV
rrbIjpsB8H0Zmfz3MDMVOqJMZgwYN66aE7riMHPC025VE1MyDIMhxbowDr6oYygY
ZT0O5BBUXEnUhCnIriRnJMRugbbG6H0Jmhq+kWtidqR6to0/uil5JoFMX7hNUwWH
ez/0ZRaRI4l8hcpopjpQtHdKJhyYuua4Q90VukAXX+yqyMePYV3r4Y7TBauvhoAG
YLP/VuggYv6XL6+AHBKjJGBpTiZsf+bzCxIZ9iUCxr9Wpv39PnxKv40DlMKfzSu7
L4MiPeFCsr+4GTNmxeAifLRF1j7F3nUz9gEhzFu68OVm8fqwH4D6CRyAF2JlDd/D
+u/jD5hFuFr4Fd+ZFYs/s/ATwyeyiFPw3eyDGTSOEt5I1drMkifv78gi5qrGy7p1
4NqPTshTawDVQZxO7l/M+NEmI0DzGHxUJLMu54X+g7qZfkY0LVHYFQDFWm4pzd59
iuvWMInzkvcWiT088CkgFMu5ufaa6ZO2c+pVmXHl3VdA6yEjtU6GI2sb2CetHX5f
puv+vIB2FKI6jX44DAasFbeGeMQVzCE+Xvx4rXVDDi2/5mHMQn/oqwuKR3CEvEPJ
kIGOudg8H4h8uyQi3JuPkEEr4Pyb4LRkvi+KKDdZzWusATI26aQV4QBgFXz6EDYI
OeGpmdpzZOFf4a1wbKxitIFCdMubcrVYiIYDo5VvD4va2HdSj6IChIA7JiN+wS5Y
fN3gKcHRh4Tloif3opJU3WaXtie+nM00uqISaDObh+e8JZV/ZKGa5APQeDmfWt7I
pgmzt3brfwRngAEHC28LO5BwLOFwSRgijZY/m5Cxx01qE7Q4ywW9sp1ciL+aS6dJ
sNZk95bCk3I3IFgGPhXRHSZkVmKnr3SKyb2PhexoKcEEgQVhlncGEceS3gU4eAcn
HHgWzv33Ta8Dv5QFuA0sVcQdcXgP+kabV3y01BKT2fDHTNhZotRvAMqMCm0qnTDU
4EeBNbsn3jFN0Cmw/zkIyz7V8XbJu+3a18qznZUA7Ex/6k61Sh6KsCABbpktstyJ
vpoP1U21UNCD4eMXHuCMHpTn8YBNIKfBamzJud3yfDlNnbdX5qB/F5ivHTp1T1Hq
AJX4NkZwUrNPZIFf4hZgNwwdPKg3/2H6KJFsVnoVFOHZI8eNaKIQEedMcaTeQ8z1
YC/YhmrwfY1uOsyOFzHnUL1hO7A35pYeYUnBYAE4ABR7hx6fgPzVsJH8BvB8PfnR
dlO9qZRTuqAgrv2Zrw9ZpAQGHLUVd+GyTZN3bFawHhT1CfPSkVkPScS0ekz/Ecco
5MX0d8Z7R/6qCA5Gqd33dU3tHGruN2EPJZ7TE7HYo/JJJHoAdUtVympb8lUA9AN0
5cP/OuWnsFAoiDywEBcQnYYIS0kW9/lmCDSm9ILt/j5mtCJbTEGmXV7gAMMwMkdt
XnryP0djJxeQM1oUl5MW1Vx+FOJi1gmx3Hg7tySKauAmlN8VUiMN+TCnitFkvxLU
AO4OynWPWy/y/l7cCfNgMlBvHX/HDDvjAroVD6ixgHf20PN40YZmr96xpxuN3FWe
f3HS+7GJkB7Dam6JvxlN/+CFXcqlC1C8Ghze9Tu62dDL2QOMXRogleMqteCRMjBg
jUJa6HLUUEPGyk5EO/wEILjlgHvqn/8IVVXNBVl5hP6/vd0hvTZrXzbIRqjruJwC
Y864B/eI4/Nn7zw9q6QEXjzLzLjyUPLOt/5RT/0WuRFsCHWiuSLf1g3J3h1/dB67
PSHlgKLUfEOQAKl+fdttGmPueR/9kH9ICMa7XOrcCEFGTk9FO4MSzPrsUrnSCugF
cxVz+CQyy9eZyJ8EyGm36TK8EsG1rblkfRB2vS5lB2fcJB8HPCVX/uJykEQ2bDN4
ymITPnORF2psOHqDWDHZXvOs+JId7rygBgGpm3tvWDcwJ+LvaoUJM6kowYdHg2+1
z3wOeUaCXImBGOuqUVS2N0NyO/HCu6vxEQjMHL03cwkeWaXOwdPneHxhhXJ+Hz6O
l37w33DEV1CJ2Ob45vIYI7gA2i7GhOW39Hr5KJfdGCsdsp8YKGb69Gwx+E02jV6D
vRQ6JnkkRytPNt52t/KXZVmFxfxeoZ+/RnRdOKmF8wzSc7sDvxG/n5rG0sj8kJEM
35s9k5NDuwTGsPajvEsRu3g8PsayhTOWxylxUWAI11TFrgbydMxrk1bzpbwDYPbR
f+iG/oP9ZaN1n2BsFDIPFFGJdmRHbFjNASfcTu5rEV19dMp/ZYxXqwr8ItIjOs4m
Iq4svfRW/l8Sr0XzsP0oD9YDANbUSx48R7U9EgdGoTSqQdyVBmQTEw4ydv2MJoc6
UdtEmFaOIapoxstMZM30MkDJl+V0YLABwgP/3IKkmc7ViQh8qahRyKF3eaPWdKuK
+50u+8MhAkSxsV0cEiMNVsHm5xQPuKeFm/1TwFJsjMk0XBEyAV75w6kW2Ggm7tMt
gANitz+KkzDpyJdOlvYehE+piwcEsjDy8h7jVb0iHLhEtXtQS4c6dvsfTEWHA0/7
swhDvi9NmmxHzMRc7v18JUT+HoWGJ3U3fokiFkoTQhysbthhWUQRZTcKEHQFiYet
aX1VS6HdhA/AD4i+nuDBs/aQjWb7KzACiN+6K5amRiwiILpcwdUAMpekFEY2YDCm
uGjRhZ9WG0Ke5QHkXy6mR1oK3RyvjuAd9sGnyfTEw31eTX5QJfKtbfKHvQR+KWgV
2JH8N7d51Av2S7umrziJyxdLppUVhqpyZIbXAhkTpKPAOMmeInrn5p1Sllbxs7m3
guAJJ39f4czBvBNv69SGpS905L5KQkDCpeU8eifmHoNRlZcePIVFL2G8T7WsFScQ
ClpxRFDjznGaNXHm7jBmhCYL3EG4JpdKqZkICNyanuWv4ljbaJVbuu6ppF937ff7
mSReWS1ezAKuZCz6YQgFuvnBVnHmJiZh0wBdNmKISBz+nbypF6wv4TMTHy2p0l0k
OHzWFaiK3AZ0KNTgJErv9WifyOInG2Bh64BSqPjqLxHSDeYeSgrXTZOzVT+Su3Pg
WgbwFPCqX8AL7fj7FljozlRYVTjcXwYY5DBWCalhzIBbTjvnnykf33Q8/iAZ1r1/
jY7LiJuvt+VKLA3fEJAQWX8+kWM2LZ/CUvDDJ3uR/Ycdp3kooWMbd9wgtvVnp+vW
2Ip2VhsYu+FE3e/SoeH0oUlecRaeo/Em0tJmCtoiZeJiQ4oZrGV2DeDG1PRji3D5
hmfSEAmEbEo8EWp3ooLPKlftYGirVKbtWg00wK9QNi6e1fYXJPd/imXBq8CAbZNZ
BzK6p5/p0OZKkFe6zLqoLMyx9MiMWPxrbkhNA7QBsxvIiIYkG5qQkkyO4vznbE4B
dY04+UUaGMTi9PFMvywZ4U1M8BzUk2Jyd0TNI6RibeHzFwWAYiU4ydgX4MXVPLI+
q5fohh8Li/Il9dMIuaVlpJdfv5itQgL4OU25O4A1N4tKxQmE8d8vInAF59gmr3zK
zR7J6lG65GxCDGSuPZvCMgbn1/KxRXmPIRa/MnuhCl/EbAYKOZWkapPzBvE9EpSD
Y4fj/+uCX2tISOXU1lTWTBZ78LX8PHwHBOiJjDBjmwZkn4ZcJy7WCXzkGOPo0Gr0
Oduqf5cuyQTchKs48xx0pNhfZPmkNFAV4t4Ox61QBGM0R9Bdn890OZKxTh4UQYAJ
WV7FlA+RZK5xcqLpcG/Kk9s1JXjgpS+4Ti6NvC2IfG+wOVswlzcPVJnMiDFrnjpj
Mk3y6YJ8tl3Aen8XmBq0msNW/58zt9wm6u5HfblNnzFq5MX1RRAqyirNGiB/lKlo
V4BmZ9YOn67mktEsEIsP451xbz7k/EsDucRqxGjsHDJBqlUzENyiXu5hkiZP8Vc+
Cn836JZOJI/KLBPudncOSG29hxf+vI2CHx8r821gtb/hGR2K5gdi1JleevLSKmYh
kygTUXFmhB1ZD41FGLOB5BDC2MlfOzUoKWSwY2W7mDZwLbXgWKQWTcPqCK+7yTbF
rLNl5wW1wy86GaolUamWmhm7LxiuY6krCP8Bq9pvcYGLJuj+REm27lxNgcxDbzoJ
3LOX0kPDIOsGxXTljuHNEDft66yoApb3Z3fwbsV8GohMpkmjfcXGnyh0Tn/YSFtw
ZgQMuRb3evpxk+JOjie4OuDDluF5hhjLeGga3QXY4RZ/FkdzCwjrDx8PB+r7bYdk
Bx7LdBrUImr345RSj3Lgg3tm5DsEt/t1RfvhECjmpXfb8QMWZUJ4x/3slBiR+Bwt
tCJJgyJuv9URV+8Uoz0lZzcM+dEkQXgwE3ERjT0aqCJVcUxQhik5NG8aLAvzDPEI
gdB7y+AzE35BgR3VAcDUqbMdRVvHQrnWkoz3pffXkrIFLUN0+Xa7vlYLLOet4NXe
9Bu3q3/Logdh+dNr6gVNjHSIsiIyhfkGe05RNFMbMC+9nrth0hHNq3gFUic/JBFi
yiv8k9xhT3FWNgPv0qG6PFWmNOXJlI5vhN8d1WLOjYGj71yxuP8Q1IRFDgaM9oOY
yDCxc41d4F80GNelgAC0x8EY49WXWVSoL3KP0u5uPqjPo6/j4xqKvHkw7UL2Dsb/
T7wQyQaIXSzlEPMIpqqRIv7ngewbg3Qu6GD7kXai6uIOJF6s1uWRN0zD6G0dn3Gc
p8T7kzIaheWyMEZw2JJEBFtWhOmkINTSmwSrbWt6g5u7FGii586EC8EIc0Xqj0X6
abQNnqey7JaL+ii9kKj8W3cJp6aDcIQRNI3nS16ufgi1N7qTtJh7ml/djW1+VCUk
ppDxiOvMd/gZNlvpTCR2VBtUTA+cwkdL2SK2S/QVsav7q/61HoTH1HYFdQHkC94Y
jk9UrJPXpHoqtIUk5VhMvagqSgrMaXpEGnOLVkYI/Zhv6UGn02JNqpEoO8TBRUPW
P122FNg4djh/NomHNRgdohnowj2ruIJ2Ml+acL9V4lZCX5pgd4IefdOvtYq2uQTT
dk3h2kOfa//uX8+iTXoCvRViCc167Z9zvmNa8ghO68Y8zCzn6n/E1HGADpP/opeZ
dlN+iXHdlNFwK3snenrrj99s+UFRoh1fk0h/Sx6SB5yg/1aA6Q7o1XTx5C1LmSy9
KCxzdH6QG80zNFeWMdJKRqaN2NXFLbAcMnW79G6dhTaPQJbJzx8VVfhOAf029esf
/PKNvs9SJS8PSOvZabxAvVbDzRBOiCJBg1hAK9sbtLsjFee1LsfUpomNRCR7sF0X
kw9Uu5+0VxlyVQ+5tGi3+30PK/NELYjD2qp9I28lFBBnB0gTHhSZaKs1c4BQzZ34
XtWq3AwktvVMVRYD6/VX1Seo0iPkanAqzGLZGwa0m+zHT4fuo7QgEKTRvvYePFc+
bEZkBN+0qDC9HEQ+Z9FZbYpbEPeRraKuBCEl27qFDmKCq9dggwtsHpvjLGyHao6a
YVgUTk4Dc267k5gKz7prsuJtWTmRqLbfVnlpbjxp/yGKfZYprbM1LZlNo477eNRk
u8IKpl8y/N2Na/W6icQd0maY/serGP1HttYQTM880NAy4ojHUjufxMUJu6mPuE0Q
4ALU4FzenXNFjsLA09pvgFqVqA+34EV1cNH1hqeTmrQi6HTxYwyS1WMnhSDfF1PU
OAkqMfIIdVapc67oJ/1iVxMMEoODFycaAn0Qb9loB0bJ0EYFgH627/J1MnZdQV1R
rKprb9sRKZK/xfSISBmoyIHchDcpiY80oD4a0whYJnC14WiLLoYhV7KNmZwCaWV4
UbbX+3RU5p0yOp1p1THY517sw3D/nWxrMCqx7Ck13Kom5RQ3Jd9Xvjijiqr7FY8S
GN5Ln89qbgCWf/F2dSbpm1gZ9HBFypRaklty5AnncNpbLRab4OA9yKnJL9O32Fzx
7UvKD6W+3Qlkj+OAxI2rPtBAn1V7BeanGZDtOgRdwp4jXl+F4HqAywxHQjp5lpaB
9n83biJP7CFTm6eK/PMUE89QpFtUAqCFfk1mKeoI37/wWP355Z+zjOsMq7aR+/IB
UHohcqG7rksl28C9l/W+s5oEfcHTgd4wfgW/76jgCQUpw4MzxsYU6z5wKR9KMKRm
ef5KxT2Y+lpY8zoEx3Bl05owsAqaEtsgLF5NEIGgZvtGGdYp5NvkEjcPhKlTFuz3
kdRJOQCR0xUczC87K+V/1UwVcUzCxlyQtMRzKGDEH4XQQIu0QSsF/3WTjePcldpe
KgJ5tzPk4sSgMV971R0Nupy2ym+Vu3Z6LSy17lkW8wt59nfzDKB/4rxXMlJ4dSrs
CgJABR43/besId16Bo6hvYTe6AYRz1g8XQwYs/6KFSCT3lm3Yt3GFwDeY8XJvjBU
ALzIobai/Oz9psDIf/c5cd1PsZEwyG/glQs/66yYSCNPrPp8D3rTE7/6AbMDAxow
+Es59DGDnTLZujoE2htpt8EWR05GmB3DbiNhlR0W2ijsdglnrDB5BWM+yKhqqSwR
sxzofJbBpZIO4a5k/SDRI4v8uhHZOPkKpWjmsJ/EUew5046R92gJg2tfYWHZBJep
gvxt3dP/Fg7fFirw0sHTlL4+c2GSauhE1mbqfsbHYiKStmfenueAqbpU+QTln7y0
Q+rLXHMWUgB4yttCEXvBnia8yktRGGF1DnK5YcaAGoLgD8oEiWox4CxiPKvkjLUi
F1XnPwEcTMhiEBzGEURYLFfanoJaK4O/hDutt5Y7k6oupm8p4YxArPzKagCsqXTG
6VHM4f4/uDTbAQ6W12Sd9pRnSPFGHIWPbwqLMSwiNvsIrtdvlJnTKYAKkU5arY/T
swOAHcKhGXb46or3geeHXDoTA2C6hv1f1f/Y04jmc0xMk/G7yTUvVwelyeaJlmcF
ciyz03anE5+heVj/x8HnG6NazXtRSZ2WmG4hQjT7RwhAh5YkfSf2auL6qUy9utDH
iXysP7yLnsd9q7ShQLXjb7qlnOGwzYaX2vqhE0CqarYY8eFB/vdUCvhkzWqQnd+0
Us+8tg8LILirL11/UVtX1EAMIpfkQGR0qKugq+/TKR+h3fkWz4udvMN5JnZ0PWFu
qfbJvEnK9Lt9Aislsbpd1T8IsvsjmKgwuJA5wMXVOdq0QD1AdvtSKKIokPET5GHe
+tsejh2rZgG6V8JvatRxNKZpGX9VfR/25J94XSV2gxTXeKdx8eeWOXEdDp2niIHQ
BhKLcNPldmmZIhDbuVHlCpDbu9L3CEpOB00nyR2cdWF8NVQwCUuiKCbP8W7J8pc1
CROUz40ZxRSgUo2FKa2PiyQAjjV3OfbdtrLzaY6DvXxLMEm2+X1ooWmXiv1hjQGS
ROcyPg4Ogtjb8o4PxmjssBngy+IW6IlZo32BI7ejY+r2b6Nne8/z048waxp6sTs3
IppllkHKgfZWNEOcrAfzlJezJUN82PmrslhYczyWTqoYqDuJObkoLLuX6LDkkAGX
Bb/g7UC6Z35CUrhLg2lVGvVFjLhjp7O9XkPN2InCUSNK3mlBoA/1hMBVzOjc5/dG
ZSJgEQyU/N1+J8Ig3yx39an69+tIKhF/AZVaDy8/7/XfaR4jeYKxC+r/q5EEHnhm
t+lh+gYi6zKFCRiC4ey5CJD68ZRuMinuF64XDX5NIIxj5EpKEj02wl+3kgO4c775
oDx9/IlO/gdyhrsodTnWlTB3vq+M577IT+vLGHP/VHyZ7fOdbJL0QPqphEhkF6UB
qVvaboO3v5bhG5SYT/GynIy9Manw9qyPD9c+U3WSqzshxcLcHhqljxXh3ZgFDjTu
m/VjPG1TRtYmEQYwnCk1OnWTLVgicTFrtzs/xKCFXYmJKZr11f5vC5tFQV7RZGTg
HJ1lxOl+hwZQWs+C6DfOUxDCVkv8I0e+oeIiWU1ocpjid0QNKlIIet13KjTNt79s
vPL6DSWA1PuEs/sUT3+XWI5uoWRoOl1qk1a+gOoDfmpeh8tNWyv7nq1gObZPgqRE
yUIYwEk6LijWRVxhF9s0PUUM/10xxow3ZWLcmgcKww3TDuNwBDVlPLL/RwGL4C0j
HwdY/b0nTbtPdeRbNF/RjV3HUqmkzoHg9nFAkNefBlYA78DeS3ua1YBPVIbju+C9
TiNT2nqD/emDnKaIOV+hvwO74wVGDeXg/vXwE459B8MG13dRHRI/OdVAAhCdlPWp
gtmZAYXtQdf2BKqsvSptaZg2neXgmq8WkeIT+IhJWg0vV6h0PFq7o7WFuDSIOOt5
juXintI432kFqLRVUMv1oStgiG0wTYz6HfLDCczyDpolz8JS3LKGbvmKFygNTv0m
hPWo6pNaYIhrj2zAHGDtWyhJxew/Oo50oiC0aaGqIyvl3IvaXS7E2vSGb7wCdhxJ
Nppzjzq4TE4KRDGRUEAQtkwGFk4ALSa2jbN7cjdhAANy7yAQ7qBkKW/Ir12CFZJq
y7HkvN3u7FoxbWXFB+hoSFZzGHVWoJrET7+psCxeI8GhhJ7A3J6xLsj7U5PErXd2
9QLoyozCgoW8wrczWRhuE3ukyDMgKjMzRhsYQHx/qbYmZlbkG48DbJHwZ4OgYupE
inweMKzKBG/ahbghwzeHwwDsO0PifX5U0zKf9hSvcO3fu341jGmtGRdow7NMkppA
S9Dyb5xtXhJySWNvHeojQyFipId9hKRfKUNSGXc5kRxtz5tBopbHIuBR/XQsoUk6
h/J0tlYSPj5Fu25fthqHLOYVlOy2bpiP8G/vvRJJBblBT/7AWwGBi+3bZbl3/zoK
9ogS2fgJDza8F6iDxNmL7N9YPhQZ7HG//TbfD2BCsqQC2b6Dl2FL2Eedk27876RP
by7qNmezoGsXJOj84fxF+lIkfzJh94pPypx2z/CiNFsIrKDHhaOLZcxow4ke9vV9
7IoC/7UubVePB1jnT4eVpLTmoOUzWt7/x6nIjXp/+ttPIKcMk+fbYDuJwhjDdGUV
hRxuH3Iy7en6ujLc1k0ppysLwMNrQ8uTeBYSM9DN+mckS0LQfgYxLxy6P0nxuUXj
fVMDqLfJl/XoFuzfVF85wXXHeEZzxo35G8V1I9+vKLApLJq9w7OrrFmWNDes8W/O
q6LE+jyb383w7fYAYjVxVJfPXRz5d1tz9lbHCgHUNBdyiP4v7KWlUhcVFD/rggOa
ws2Si7dX9RyCL+FuRnoS9lu5sxGsLU4r1BvanxGrBceCYoW6hZlzH1TEbWI7M6s9
ttDfT1ID67K8haMesOQSlK9muvuuIj7XrT0fwz4XnKKz077JbSiGsjoph8ypNWkZ
FhMazkTyAwjHhBZqLS/+Q1xuCZXYKiMV0A+HY0lkul2g6qeDBU84G8l2cSqaGAwp
lc1q3a+5r7FHTk8ExFFyYZj+O2JOP8wVvq5AD5wg9ZT12l6vEoO06cby8VQMsuZp
zkeDHOVYkgsGx/hw9on/q7kwMHHZM2Ys0OQBpA5PW/nd6MWiiOwUbOXIM6XzAhey
1pWWMcvb/lfoYkPuuUtjc2nzYveItWt3zvHIApqNOAQVF1/Cr2KCJOInFSoRaw2N
qWjJNysjWeiAzQa2uhYNfTLxcNbBowxufDwljvLv9RAN7iXKwyLwjmG1MvNqJIpQ
f4RxAtvQMVPvi3NzaNwNUzzs+SDN2QWYHH/l6n/gbiwn3nXe7kbe+vYQGGmxOo2T
Xa+D/mKlUO/m4vlSZ1Op9qni3BaaM9mexZFDtd52TZf3ZFUDq6d7/Xt/QegAA8W8
pPjDeL72bZBSESNReAjdNxOjGlUFVvSu4uX4pbi0E4shgqCDy/d4vCiVkvW9lNwk
9llSBO+kpeAtAkMgz1lMPMB/Lr1so4y9VmqkF3LHQxDPwIcIc1a++VRWlQA4Fi6K
FszvaQt9uSdbCoJ0PODW13xy0RGCuZwRdEZhYq6ScQs1suXShfnt37E3y70F0arU
jLKTlcPfFJ1OCZy5eKxfkZW52aJF+b2x28C2c9ojsgrIuk8DcMsjYBTdpy3/7yZw
BAbvb2zGKf+iiRbokIXDEz+wyua7gRnajpHiWWpb9Kmzh5p64Jfaw9baoy26s7gk
nLTUs8NyV3UEafJXY2VsSS3CMpN7BxzwxXARjS/utu7u9UqqJCw3Qeqps9zr4lG8
BycqRt0/WbOcqoyZCa5ebECvfoj6EG+KrNKifMhYPZTQ3CF1+rIUauLjPtwXXfco
HD7JTCFZGeTpvNa2TzYVASyFCV/Rw/BLypTdf9IfNRWXzQohrYEi10oehcWquNnc
5thoDytyQQ8daIBPwUijFRqaGxtpQtNVNpEybHPHkaZUTQzRPOfuGrU8p/jx44Lt
FESl3y1VE9IlAJfHAOSk9T47mnr6tLOjYuPFLlZRrpJ/n4zibhWc6BB9z4RLCkvi
H5p5XllZsY61Z1QsKcI6m56JlCmGCzDP8f2yiT65gJhJYNKOeTYUe+dmxHfygIM7
LOYGUaRO9N2XvklmYS9lbzwhNF5SN4jDTWVF45im2fC8khbaD4QDeLmY+1WX0eVw
vkjUyCB3f/mKrE1F8MwkBlYRI2wnlLBzwRJ4YtyXaWdxdBlqsRqLuRhLdwvXy/+d
Ot49FvdpxeeHbp5tO7+XPcOQ2Mf/kmAfKJo2teFLWqtHerGg4sRhGw+Df1d5ARXx
Ym4rSXgxkUqFb/F5rVC4wXbg27HfbPyT4H5DEXBcu8mdse3fohhkMTgol27AZzIO
McnDVycEFu+AeUNAJFtXRiKYGeLklYHuVuUbOICuHqFZBrMotj+M2lupipyHp8yf
tQMZVLaMo6ur0uzZz+qGAJHzBA3Oru9RKau7tCNrRYHwclCcp0QwLS+COsc1Du2B
FyPZ8Vyn4tfZlnIW9MujCycq3GUTLc+n/HRbILRHlu6cu5lZ4Q6SKa1JvJFi0f0C
0Ycwh8FDvEkXMvkEQUu583Ls8ETxz5zyorU4/i+AUgksv0g+duQmMa6SAt8s1SIA
Jv7goDgI/84RkEwWI2ULiGx4SKX8m8cAvAmSB8UVpOtYMBGSAEriHude1z11wgjW
rMDBM75IrkB/YQ4SAJtUuT9lY5X3qSWcNnmRsXSSY2rfUyG7I5FshQBhwr81rQr2
1fxZS20oZtkDM8bdZSdHxeH3HEb5SXfcz+Awqt/k1OD1PNI2jV3bKmwCcaJPX8ZF
cTe1WPCZK+FHF9SJ0DPStkbDXi/kh2gunAn2Bv7Z6apkaC+PwL/nv768Jpr/Etlc
gd6elejkJ2uLHHXxA/hWj4ZgzfhEG7WFbfxK42mcIBW12xG4jtdBHBuiXp7dGbVx
/iVXVPLRF180P59TdF04Dr19VwLjMyRXbKMEpe4Xvo3Xt/oz+jRRRrLsEgv1JYUF
8CFDLX1cPV+dCsTRrTCdYZMBFE4IQXzZlBwzXftle1Oon3TGYGq0s0Lck5LHmQeo
ZDa7OjahfO3Kyt6aEr3zs+zTiTsWGakGNrYBiJcmWeB4kfMuIy3ztjtYTGaGt0EQ
qGNm5/rw+fImwnNfQ5p5UGwMy5IQyHIDwHt5mzJqIQ7egP+C/dBawMo1XeRl5zAj
g2/XazovSUO7rUePLu7KuvBILcnMtb88+m9Uh9sMgQ6hNSfp1ajIsC6MuSq2T4yC
7kxekkwI8rJGH3sGzk6+HGIhLZyKLBIvKYo5gKuayxQA/py0ReEhg6feiFyPYXQp
jAchyqk1tD6YmNYulxe5CaGDFJ8keVvlZB6AxWFryyPd8BEFxiS6yl/eoOgvMN+X
xLAYCeQ6B7CO42zp3bvl4bv6QqtQ2ea2zfbwJ0AaRH39VkHx9pO+NmQzSK5Vz88T
pLpLQz5/+d8eHUeVOAOqknILQbbKUrf8BYOIDtbvfQlvR7eH+Og8cvQqgicpsPBg
4fvSqASmdMoJfddT5xks8kAJlBgs5j+AFfJp+s8QnX9680sHD4IotFmbwhceIM+z
gmzN93FaPvC9BLF2C0sCIHOzLULJQHB/KzghgOfpcCz7c9HQ2kBRPW629j8NNyA7
jRDRDAECCOBZskuaRuPiLW8aEAf2vqeDVICfAeDXmiQNcF0S9rPqI1t0FOC939fw
EE5UEPtq7UOkYB85/7AJqmwR7z0aKYqe5vMaLPGekKqiua9buReiXwT7oyxCd1iH
dzoV25qIV10H/QXo4tGTumUNuf0XrxpCcZNbRMdtBaqGfodymk0hFlqthqq04RgG
v58VzR5SeJDZaGFXOYL0Ykyfg2QNOqu5bSMN7ioQOsZziqvWtBdf4dPbOLARxtyc
bbW7hJJ2U+0LBKImds05dACLNVoUVXp4vHQmmwq+hMWOn9gvl1jygwK8/+QP+jvG
ZKcQtvzL/Ygr9lyAlKK3IPhYtp8v+oK403oPhDaoaEb62VqND8xpmUeM/HxSRqJW
1RumYQNylw7iROOdyd9l7SVbSA4Tar/vXuBQe+AGdj6AQCqzzzvCAJMUfdGAu7Mx
w1x0K+ozGpkdaU3lOVjKySPgcS0MH7i2etwn9/p1ZVunN7045U4OY6S/y2PFdANq
T1JkDLIXFsmiz0+rb0Fej2jsGWrjTJrfbLqeO1Lht53fTYbTxSz8Q1Q2oW945M49
H8XTJv/K2G+KMt5CHc/RotqmiCdAEE64xNBgA4e0G4m/7yHb4ovpcpwmTj7IP+ad
MsjFUolvRX0NR/m1NSFf0jXp78qbsmx4Gt0FgDKcghzRO9lf24h1WVytfpFbgzaU
wTnskfMpJaydZNO+fzNXXCv4+j98eHP8oHPJ3VsPpwMloMbZ6wWMqjqfu2iY3bpu
3jm2qFQNeCmtIf86rfLha4c+9Qr+bDlT6xxMpqBqMEuZvCjTHWT5rhl6AiWxLbsx
9M3L7wg98sxkvxfGwrlxqlfl5Mhv4aaq1/PC8yV6qbVGCV8ULOSGvlJFGv5F9sxC
tZc7D05AyOlmJiUwDjmNWqulQw3ufNZGQuej58F01oxVl7LegewwKK/jtXx3H2Ve
Qqu2YzvIwIx1z2pynn7GbOn2GRAx7DYQHg7EKEDX5B3yyKQOqhpMdDYja4HRfa7J
8TefsGpmBv3F8mKi7AftwgBhh5oB8SELVYOyiQgGrg3x/JQd7RGw5af/ixgnsvoT
atXx026+/4iJ7kH1CVP4W1CzylHGBGT1pt922BdfdZT809ygfrrWaUCiKr7yl8qN
VJMqa2wW85+AvTTk4VAdFOGsTxwvIViQhJ6YbGGHFTUG1hSPm7qWoqC0MOONVHSw
3lCxKy7C7oAulD+VaIqpXdDnzCC/pIIIJ1tjxtO2rODVs0y0QybLQFjUNSzMi40+
9pNUPqlEuOoRgx/BEUzpdzKltEEJpgsZGgXh0MDTtalH0N3BMMcOm17aMwzQUKNF
brLo7Nh4zr2qBvAZa2AaTpkkBpfBGf0JGT6p4UmGzqEZEuuO8IBK9/+CUf5/sYWI
rseZ7NnsPWEkjEBVr4PfaTth9ZgaJugeEnK9ZVmdUTxACLPIQ5XRLPo5shtnzefw
h9IFhkhfkukYfKUkDb6IC9LAgiR7lyd6HQmb2hx1awILDolfdXO+gMUatbyoe0zX
if0ahW3jzmwzwIOiJ/BKSmXXsYN6HiSpGotz+v9R+1IOWKQsAqOnhLrYxyQ3m7lc
+PW6xkz+kOhd3PvnpXHGRWaHpv8xLF6uZs1qVJVnZflvil6LvH6qEt43sU+jq2Lw
NXdHLW8St12Y3sXsdKi1jB0mQNC6nG9roUuI3j/bg0z4uxHzF3sqYPbRTSd9M33Q
TGwkIwtmuh1gE4lMRTrB4N1ysbNMHxDAtxPvXidh7EKNQy7EeMJlCTDIOA+//ZzB
cop8SVOqh0ABYIoJQxXsgVl8ju7/jxVvnv0Q+aruSAOBlW3kQ81DY1LwNwnhZ7Eh
feoFVxLvh+GffGPF9FVlZd233ZS0cvds3xF8C0X9mVjpQWrznyM8o2JTTqlVq+3H
rsM98f6YuE3re4dEo3t4JeV6wdbPRVYWIFQAZhHIuOFaUD4oABX+fZ66PhuTIfzo
ntKD6BnvpearD1qT+AbegY/pEPUt7a6xUr+VLDjj0G+54bVR03s3dnmlzBihI2Cv
9HTkQoZJlbH93T6ASpZElLqc0GKmwcEJ6h5yWILBdCNYTRzx1IO6vfqKEOi0wzSy
f3RgMIojtnzboP6uURsSpolVbLD4hWhRlKKhF7I+Q7JCZ8eaB69rxL+Un8NuA+4M
PPZtx7/mnRnuaG1eup6+4C0nwPXmsx6sG5Smbq4Jnpv5TRR9tN9HBYLPW3m8Rp2q
KSKl5YTODD5Ooh1cW6yru6cIgpW3YctxJCo9cf4sHs9GFamwzeNL9y4b21TFw7Ak
zyna5jZPZT2imuvsFsbK2dxFvVrrhbR7BP0BKV9lBw8eeepjgRh+wEINM4UybZnD
IHVO22yt1xfoInNJqI55P9Ieicux75XoVwUVXT5IgBP/3pYQxGiQnO01qIflzJ0U
pFFhIorgp+muNRlde3d5Pt76cwFO4kgVwY2oI0wQ8YPo5WESR+VaBNBWzY+LAJjs
ctv6/h+DOIiAQ24pA7UkZWObxFs+JDwRIJg3cGLnpO6WZq1rLiEuCgt8XjvUwG47
breFJDvRBTBNS9toGZK+P96biMp/A/bXKnBGMGI1YE99aggBwZKukQKjMvIRnmbV
bFyiNYpi3QQ//NdiXfsoHQhWhrd/d/QFqtj2EThdOlK3VlNMqLO3FFqXCJHq9Sgf
GABGQZFBl+QScwstS5i5FGGhJqQvU/vJiV7wdNtDPXQ2bO5oyU/UyrQT1yX76BC9
zQEgxxoDgKSYY0mywivNzFzmcCJQya6tPUaJ/4JVM5HeFsa1a8q778Ma9cQqhbKX
tKiAhyx9/e2c+c0FL+X2bOttr7Gavl4NCiZ5A0cUnQHXKaCw4HsA/otXE6HClugb
SiSSj4Gh6SPIwKlof4lkwy38qZNPa6gI1TrWoItB4wvHponwK7K/D+qgSiSZf8D3
y8aKdYAlJ1z5JWSxLiYaYVGdo6G8sSuHZ74FzWuqd0CzOKFno4lBxkvb9KYMeObz
qe5xvJVlVIzq5OEl/kJHwPkizXVH+1O+tz98YRmiVNsyPqOyrBPkX4kLaTm5n9s+
ngcUuFEI1s6mJc5JTt0awz4IbSXxkug3cfx4jF2fQfIE3Yh4hGRSAvDcZo/UIx+7
BPtg1Bg+ovjGeyOTHUtmOkIQPjNQzyEXKcUlgwAkhIPDSfBx/pqoSvfI+4Tc7tOn
Q19ICySx/jmJnT5nKGlNukdZ/XORAZ4npgI8cAuET0ElvHazLzK0ez1HX5J7XF/6
bBojtqDGrSKVpIHTi9ZJ5vx20h2SEmxfATdCsTtbVHYmq8AZQTz9a6o67UIHXRV2
nIKhkriv+9dJPhSvdG+iSmOL9muREJ1VpBQuv4dYMhX3nfnZvWEo49hgQ258zPoi
zbeRSx/5GyFMACNRjHxhWHOBp7NKR2MFx+bpoUcpz+dAUbVsY+4VZqHrBn7fBQ3X
CXLUYWEE9VuujVQXBmYWxg0QHf1wSXG3ofpv5q6pDQ0Ok+rL2mhPgoC1/C+STBAz
M52Le3xGSMlV2/8zN2n5+3mkKATvJvkUw1Vi6lHL5cGoBcMT5DU3l7vYKJ8D2GlX
CZLQMkJbNf6Uy99J/gffIUAfcCoAzP3uJ84HECDi4a7DrEqigmXvnQRFpIuTaE7L
h4ru0so8UAdW9adsJ4FV/UerpjQjRNROn9P7PxWZXbtOo5ZqsGO8ba8j31dxB4ku
1mow5Aw2Zfd9Nnv1rzkIzElMw8ro7S5Lo9WEAE6lDdX5YB8lHoynlNAWRYkAYsi/
DC+1qocbYjTkyRp/JD73cNefZattpm4BdYezs3i5BdPOABYCuKtmLx+OfLIKvPp9
STKDRH4oZti9x5w4z5DBcp4zfoDPa/y8Bq+zoGDZZN7yPJBwTZkwXqsn1nrkPu5w
9eOK6E8cgFPxo6SQSNC9zZYde4btMCLB/JC70y09h1arj5De3PB2pDv9yw/AjkZb
vmTCnm+BbDM/XJy5ZJqc9kttOPmNtGuK/zLWpPVoXxIc9mVfieQi8WcXfmXveb5X
rhd7Y1xjSLXHYlbL6fc1tsmxySKuM2vN5lgK1bNIHwcha4xAVhl6CltWrb2Qy3kN
5eNxj70bhJblUDSUXcqJx3xmPokQTpLRaD/piTpFTBWjMtVx44NAHHV9XcttDu78
lU2ybGe6PCpZwYUIefEMR5wkTXvZ8UQwPX4QoBRHzpbUAj1rKTT0WrFovb2Qc/E2
zePnA3srKWs4KYqLgrPsiwFQRH1/VDlIbmDruPIrVUwuRlhnmh4B+9x9/d2ufUOE
wN6ulw1IUjVcqZdE3htFg+FebfB2+WaaoqSjA0+bSNz4hStqpMRAYUck8LhmdISl
Rhk/fPKKO4wPUW5kTtpiFqLNDY9GWlFyS2s2V8QjxIBUz5MXkrRgWQtdev3x9e/e
4NI8C51VwwkFuv+cyDGD+1coVXfN1XtHCa98y11GI2fa7NX3nt11F7CDC98kK92a
ifjdlhx/62qBx7PIv1BO6vUvSICepxOkfapl8MVdLFWfpOtrFcUTk1B/52i1j7UI
xiw8Yjkz6NxxnxfypD7h8eYKYC8dDk2AEXhGqrJ+nuEmtz46ndhVmFC7tvcsf3n1
zy7G582X0YY3mGweApsbG9fPk/wmH2RwlGNrhuowKRKaXZrUZ7ieUSVKXr+dPYU1
AHp4yZ0norNlcSvUjdYrchN5BAjOZEHS1U5C5IsmZSppnlc9wowIa7LTm2pAdarm
vs7obCrGTbWiRr6XQBszT93LKMj/LaQs5yTdjIgdVSKdFM5pBEeoZe4qdqkvKXz9
fbFIaWojwmuv7wWGLzVRNC3IdF4M6Foy41g6Ibp9l7ybP7VvrN1t5KAsUreUf342
0S6/Xih/Q9+MZtV6/LnpXgoAOyT4a016wfFte0qfkUTxfAUHvHk3rvvKk3KhrYQW
roVXzAvWIbjee5Vj+OgmLY6TChIX5tJQ7GrS/IoRwl2SIgOFfM44uq4zVgdzhl8O
bGDWTdU47sYRtsC53EMAQtaKQktbmNW9PyBrRDGajFWM/1uNRT2NFmlfOgmkDkGq
9iJPFBChE54vnkU1qg9n5NVxuIAh75M9cVX7TZV7h8eiNfuuYDO3npZz4DTUwa1d
QNpqx8hx/fBc6BrrA5yM4OfFhv0y7NFDM9AZNmLhrZ+HBR4bUq8b30MrZ0jr2eXg
uAfvxtKI43EKJTyj8TMrRhXYm1TG+KOAxmdY2nlwv5p7Xub4imm/ZPdH4ovfKfRP
ymCS8on1CjtmwxyFev2ZIfdbN//r9+vv4ggC2njhco8EITofsoVbb7lUPQYrDwPA
7/w7AK5rs644yV6qf87AoMRuXpiAuxvY36TjuJZ2xfjhro3tDCbXEjmMo6lU1jbd
LDb3ikVyEWFqISSUnx5dyU/o34iSLNZmONbr4fdqiP6DOPuMmJyCncplthFP7nXT
szEtiYWBhXPekrTCQCXIT3ev/u6cI72xvv7JOwLnrxKVYjZYALGtH/69jRcz0vQk
fyoSETSWI8WP+zwYaHTi/KI/P1Mevozi43M+SPJdJ/lu6PpRLIGUXrjBYNPhvIsp
n6ha91fejYCtrc/z2x+DDtO4vtkvxJvy/rgjV98z8WwkPuJ0FYjPfZaCAJCo2/iB
yppzaV44LfIueJecLwOBSmvz6Yrz+2s8z62gQbfQFXVjNfXeQ80lSMfl8Ra8Y594
w1YIG94Y2b9apFiSvFm3m3Q1lI6dZOBrCOvHtREfTwM0PlLNVb7GeTH94yGEzW0d
t68grkiLlvc+est6V/L6mCsI0ZDqDlzOjL0aTSglXF/xVlNu+P/JIwjViBj4V9Qm
4a9m7Iq5DDg6WaUGNy5DoqBNhngUpxrtLja9aFFLLUM/nhXMv0uAgYLJzNR6JXlA
ARQ/rNXAPb7JjlYKqcvREr6NALZsO+7e8F/d1omwh8Djbm5GNHs34Vuu72IXH5EA
KpENe6iHq39JXED+JpC8fn+EUOkgJu3qV3/uD6rAzLqO/Vy7EjmAneE+cN1qeuLU
/ZoY5k30dmZrG8da3T8V5zq7Cw0qRB6UIw8tDv2+rYCLWOcfIFIXEPStvrXf4Zso
F2KAnNDx1MCjfkPzjXEKkZdzTHcBv1YeZKy0Z7YjfelQWaVD1omHXZJQXHSPOnhq
SMcGZoPaOlJ3HUkocTVfI0ouv+3bW0bOJllHU8Pe0Mnse7L3uKP/tDyMTYuCB5rn
Q5qOmFgXn5NKCgnq/x55qgYgdqrXuu0Z362F9tZ2/5YCxjnfEQm+ch4NqVnbSKOv
+5Kn3JfnZ3QNTvanJKPRruX61zX4qR8HXFhBgaKnhAIG3FQCxIi9SS3ATwmtbcWI
QOgto4+UG5C1/WLs8N2z0ofAyYdU5KwetvW0d7s0/63FzN6slSwfabbATRVLs3U4
iuBg+LSH0ShBjrGs+NpmwMuVYgVMo/AvOTmwfKD12+bW8URaiByNwr1VOGnjOXmi
2VVEqIL9hTHznviMy2iTAEr54/6vTKBlxKXh3MCdjEq8ZHiOmOwdoL5iV4wOGGqA
hETWDoLfqJXXO0NB362mZybnt8X22Nub5jd2eIBECDyHXfdfDtmPgQJ6/Dxp3y7x
WRcaKkQCB/57yUSqIaHGd6ObVJc1udRgGiCGtPKqlQi5g/KDK4c8vq6sq0liMBCS
Ljj1lTpEnuqcu6SJRlydwzF7zVdY+tqa8ffz+z5UeayeGV/N2ZG8U8IXf5eVIRfj
HLunSVFRRDX5RA6li+vvQ8FwY5CNRyftjzmotXlhnUMV7kRNl1weT9TFp5Q2pMKo
rfOPU5JtVDVLd6g7NDWxTlcxctAZr6uDzwHGO1HEohfvBCFssdiBT2PT1kSYCAkT
i1uREOw7TxRJeZM3D8ZLROJ1MsZeJLMWBwArYYktp9q1i2upzYLn7RBnKAwpzHz9
vQb6g1kgBgxJYCWzkAhAuXaBnmEaeuhd3keODvRH/TLLH6cD8TGh9/288aT3lX1K
W4DayDjD4X4w655d+oNYA0x4DqShaLk4y2I8R+c/JuNovWmkXjZ7GdzZArJkAdeX
sbikOhSiCwEU4lqzSmIkyapQJtsCV/ODO/TsDwHPEQJZI63qzxdu8rDN9wh6OuWe
HaJKqYuWFhodfdnfBVMU4drZIgXbR9AHt2/Fei3IbclsLB6rHXcj3lRc4WxXgsLT
Kehbs3FnGc3sgN8ROeuUWOjVKoS2fqneUR6c7+EC20iQr8AbdZeUQONm0sNo6Ig+
wpnP4TYM/jXyKbFOqbn9NITHr45Tki/NliZ1GduR0Kkyq0uv3Aq88cyGv1CaV64x
C8cQQgUvsk6yo8W3DeqbXWl14rBRMR9fE0EJInVRfCARzjHLP5fcgHCaOnRb96TK
0Yn+5wPf4UEJboef2JIrGa3yFLCnZFZYPmPi7v817jLQVu+p2dcRU/lmTPAaV6vm
XMEU5SzKuGP48cuhmOx35oa8WzXVcLsBgx8pfhInOr2U1PjOFt7ygH3TC3DF1NiV
3l2U19b4RLNnC8curntVfT3AjH7FmWyg1GTzYD/r8IyA1gAdXANW7EQ3XqD4JqEl
6erpM4HNeGK5XRfnjDNNRla2F1RqhCNBDmH1+yNlJN1XtGEWT+Y8J+b1bNhGId42
my3LW7E+FsPcqUPx2iigdlbkxmrRqWht2JYf23wJU9zm7Fm0i35QhUFR/Bbf0qMN
j6x20glef6oaux72yjwKN1NiuwJ6qzOmMJ4qvbEdHgQIL5bhyKmIRZoY2ToWKTKH
cQlqX2YgcYh49B1MSXLmpW0a3Lag9OmGX6nVbVXbngbe3tMyfNXidendMZOoHJMA
3TIMmN2wQuEMDFwtVsNxsfQX6Gs4VPteZfkNf4HMLoElDkzIjYqibSBk2TjgXZ5F
sRS2SRsJdTMpkBKbOnB0jGYkxMCRkt7pg7y0IyTPGUUEoZM68HQIWL/l087ZR5UY
8zgxG+DTFZGG2Shj2bkdnk5izncqscycFcjoyq21ZIbcnFnwtn8pRIQRklcWHiPA
pjDXeSGxwKO6AyU0iCSJdUTCNZuDQIMadsAoM+6g8CGUd2xaALoqEUMY+lhnwMYf
IFKC9Uh2i6ABFdS7aByDKZHnTW+o7f1Eb4LXcg9efWXpnLxtpn/EeRPfcKh5xf4t
jE0brnj0HINWlB8IZJoH/Ia8xcq2SBr/rshUB52zklSJ8wzpUrgQ3xUG1YTaxFJ9
JbdhujNeCqDJHlSLo0JYxlV6ex5sUk5dhNfQ+gVzbcHt/PYOpcyn7gcbzGD9yeBD
VoIHNue7/ZAokKZohzQSzuZWNHVb5gyzRISnZZtm9Za1kraN5LZZHioLPXbAVX0W
h/uGG2IadFau4bVikVMBkj4E5TBDS3ZRCMEBZONik7KYz1VpKUxC1mo14nda+r/D
xJ4Fa1iE1sbsXvJMSRKcU9wdgkPsnoy+OUso4WltBqM5Voei6lI2Xa+IHxFNbvqu
Nf9mO/roWqBBPpxlDijusct97WKteFtcnIm2RPnfVGmiiY4wVPfQmWgsR3ROHBJb
xGpLfnhuPljjgdQYsEDjCu/ZtDXONwMPmWphieg2gvxHO5L+vBkrubza5G3t0Axy
8vuKiVKlcDPD6oTKT7qPV/Kg35Ps/DFcviJzZPy+J1ZVevGXPc4Gk4yua5VpfMSY
t4caFY11Stn+sQ/cm/9/rGN/zM8Kln+JySbs4VSTmVL4XvtXJvEntNaK/Qo3Jv6S
VzpNc3YCqHzTH5igwLeZokhsxkotEyn5wFW84cs9DJDxO6DgRolfc6ml+Xrc1LIz
1DA6p/y36BHg6BiNLB1kS79VWrzhGSaCw0zGbaC0YrcdN9J2odSTshTwWJl4mWxx
/zz+A3UGKRWD6AJh5uegiVnyZvNhQ5fIIyE6109/4/jdBaRYkSynplliMMeImgOQ
OC+QNXNot6MAT8bWCv7lswQE2eCOE5M0djDywMeyuiPD3z6cMO5UPgaadinJqJgc
roWB93s7d9k2wrGb9k/cFhbi0+D5oLQJnCW+FPFpyA/TWoPBmILUNYMM9vsZQViO
NSNB+5SiB9KtWpwm3fIg3UJbQIOIUKluD5mZfZ3R1TiysAl8DNKSoVuuCF9iUbQG
bNqZPGAzXu2FH5je6qkqB/NsBdgri3DE/ivlG40OWCv4QMP5vD0SrzVVBrOGKbsh
L0cAvzaEOJdAz7U6s+xjVntspz9BZHb/hDn3TQwV612vGLgRv02Roy8fzMauWZiS
jOMSshWiqKbdClKIG4F9c9lpeinhwk0404Z4UL3X2RjNq/oZJCzj4mw7HIcwtckc
5Ty1xvctSe9BeW2sj8c0EXh5sz3mURTu9orLHdEpYfJfkzzGY+UJO83QJualUzdG
j05BT/penynuRjNRBtZzNUeh5Kkmc8u8WQ2Q70DXMM7SET82PFnGI4CYBJC87+4D
yP+29LdK8WubuPVKkPvguyZTbXRSFI6wlgcP3H0JVIOFmrAWMJO9WHQ/+FIZ/uKK
Yce8ni0rgld9j2H4Nv2JQZdQlJC+eVe4zissxFBHfvLEJwaSwNNtVmPRE3f9++9G
e1DNOr6MtEJSRR3kx/z7fhMweTbXkfI7dtfFDXJAX3b8M5QqnpZcg8tuIdprVcww
YSn5SwmsiQkY5fBoGTOIF+XiRuDwEWv5xB0gAOJJEqN9ssHBd1oIXInB1McvGWXU
amzPfyAE3A/A/3ltKohyGFREq39dvL1t0Pw4gpIkqGhe6C6jq8VnBKZw2hcSjy4R
1kxayE04zdBnPdFi0djSmNF8nfTReVzgDXMTyf9tiznbA58HQN/anVk3t2xqJS5E
Fjm4AGb11+3AqF6NPsmSkZUsWhNJ6elvvdNfPaQuSJjW+5whYj7echbPuYP+lIMD
6/IsFeC4tvvURIb220i/OYwqXh1evGn7/8G62+dtieICzgoa6uAk1+tRDBo39DBR
rlH7meI3a7RP7ybHVpFI2wQr2gEVjRdOZfg4zMLiD85y3vyC9rAsD7dv+kAiJJyz
N5sqxA32wGk3yUJibxaDxsa3nci36OioxjHdqrjLopKqGfNY3R0/f+bnMPtG1Exq
l+hPw0VcflnRnABRVLYC+q7cH8lyw2pNNyB8pN92jQtjfkPYrjecmI0gEVjSxqWe
Ys0q8DAzv66d7EVUjkb0A4EdN9PSVkY3o7cfOTaaijIBIQMsW9TJFnECbRxjnxwQ
9pF6tFmCIsy3Z+jSUjgCxNYF2ch1a9RLi0ezBi9j5bRI4StfrFaZqXSHPO5429LM
jUdzYb7S00+n/8Kb3K0T/2/bJVzSsWpagjnnipQDUPHIBtnTVr5slXrSG5BiPANG
vQYXO18wewHeH2+msYyKtlgHXjyd+Jgs0tCQmFm86gu6CltIazDZ/ZziCar859Gj
lb0N2UO9TZSVzquab6Be0Wto5UZAebUnxEtYzxO3qJYQc67yWvE5HivRvMHkteAo
oj395K8QfOPERnp29/OqtfDCMP8BI9M/3VKtMyireo2yviDXDZcy/szWgmduLqCC
ustLBYeoFmuh+r6tAasnmCP20ze6qCyE2nRVVLbFZdKulNTaFdGNsS0Sgr6KPrCL
tmcKb4zkk88djbuMreX6qw2xPt23fwIkEbpH7FF0D3eqrBuOA1J/D+e3ZbAnYt1z
O7l3Tv7BFGjAGu1m7u/Wfd0Gp2PtaaXHUzBVFxh7UbNa6e/gwaPkdEwtpRzwLyX9
Buimg7gdIMwqCMYWxkPNY7eDeQbOkQu/8HkW32Bw5lWtJGZ6VIelN7dI2YCGrKp4
2+QhiKzzcGZ/Uk9pWj2IX9LFLbDJFWeNXeNENb7HKmFbzvIuo39xdnOniY5VPTjs
UoGsyFnafxFSLvGwcpN8VyB/0g0rYkDghRD2C013Y1RhXy8/m3+kZZak1nXGebyS
8qcyEERsKmBpVzPWivh1KsJiTdwKqJMgTK3doyPNCCpRgTz3mZQFGfVbHgFd2UJG
G2azKrHUvQnPXFY7yUBYIDGY4+4lPWXGPu/15mYBq7ocM8LBJ02lDYaxyw/akR4o
9I2bBPNFCg4w6qUZphpsmqmMFsWfO8QGbJ496l9H0d+AhbhSOBPyaWPjJ8h8abIr
WA5M67Jlbp9yeODAvS+vUnxx+YBS7LKwwYGQ8qrRh/8mc+sijbuEfMPspJl6Yh/0
a7a3LBFtJEGxX5QP1PhQp1AS/Sjz2Hu3f5j4Tf1dNQ3ec3OY+lsIVM7wTl89xbIr
Zw4OtfL6MlIQUhuFj3SR6vJtP5wN5Er+gsUWftVCvKM0BBiE76DtSJXuQKKDAZrY
3XQoarKw39k/okYD2yeY6BX5dEhqdhUYDDBECMrD4ME4jhqusZY2hPEwaUlQVuA8
FJQ+W/GU1j9/QuBnF3tjQREYIqWjFc3i2yZMPtZWbPoc2kna1Ayg1vcpGIUbh0Lu
qRcUslZ2wpekQtsE2MMbVYnEyMeBu0yTluSrQ2n4DgCjmnvD2icIOP0ddTT5CJ+h
fgGNbMBLo5HSlrqc6kLN5YKnHP3VwP3scD2nalESkaub9StvZkojNoIsvgG9KQrD
LRG28Hx0o/3wZ6NAxQK7LrRkDgpdLoCQROz9k9Gw4GODJ21BLoDjAlmck3xQzymA
OruOmdPgOXcemsxM+Mg0mSZkrIQzTLYSBPt3jfXQCbsKgU3u2ynaVxKpb7vGewh4
wV6snzUjd3aBS3vY7/2/pO25WuCzwPwNXwXgzA9pF/tykAps3nPJKR3G2Ym5dF2U
dI//h5cnhEfL/hdHNkaF+M1vlKR94ggFofA/2SScv30cnMME2LoBsk1sV3Mo3zRq
LWN8qMZ2ae90B5b5LxYqOBgLnovMe8Eyhkc7FdRuwpGCpgznkhKS2oXbfaGzHOCG
iO4/y8TX3IDccn6ryWCj4OmmqSE6HX9YGZwCCL0JSdAlTj/A/MHKlY53jtd4LpWm
/R5xxiBmadJw3sSK0dv3FuQ9pdpW2w0y+fJ60/4iIZIkPL7dmin31i4kZe2EF1QW
OP5H26R+8St63JjEtLTosLBfyda6T+9Tcc9NqBbIRExjUx/QL3yBIE7O0t9c4+gj
tPLAEzvfm8/2XZlT4p/DUvMmGeZ82cIdPb03IS+r3qnuXo8lnG8OfKGyz4QZMNeM
TiGLaIQYxtD5x8DjNZNjAm8Y2eEpqti36T8EHLu8PjpXdcgHYBFn1NKJ5oo9yChI
eUJh5lEfQCsOGcxjAwUvwscGJoU0zI9Xo+C1o0+IGsiiSeZFbLNw8RNNwXbFMq+j
dZdg5uJDmoGEtPikeJR723mHs3Z7selDexTpNhpaKXw9lw4aXQ+v2ZJgVgFxzsNC
BHzArIRvXtXy6iMSUfmGudsmyZGzqQmMXo7kiLe1EBPOhp5x7IToMib+v7jk150M
PxwKnxvloWk2oYnNIkNvZ6Xffv4secNCnErMOiDCH1zEMO96V/UjyJFM++Nbtppk
T4OCAbUlAzyy64745sVlZleAxsy1PWuVYKM6/RuZpXQ+z9gHf3XRjYnaBNKgeRkw
8QdPsu7JWHqcIQhJbGiSgHf6tqfVm+8pnC9u2zm4tf18g3yK0rH781x8mO3XsbxP
8v1wvKiovvfqbPz81kOoyfrituFAOCksETGYA9eVrEU/Fkzu8FDhcVV0JSCZpscF
KJFMyEigYq3MDBh/7YTZkmr4LfyL8IQwQDmG+kq0e3xcvzeqKVe3sZX1GHvmp+Az
p6YF37FhqJQl0hEwq/cP0I3ee20jhhN4qVHM3TA0nJNcyBFnOVbtnxhTtVlVcTWU
j5rIn2Ghl8+aVmyeGtrx6IRwPOrCGVIemm/EliIN/kKaC4YW72GkeNbX0njehGoh
64vemHdvLNeE0fTsPjQh8o2eUoVd9QE/pZwAweXzBDoAKvih+1NFYf0kWha8PUAh
j17chAB8JR15SZ53KDhSNdEDImC8v9lJtg7TuUywl9wwNoLDfv0hSsSZYlzZ156V
Mh3kYwZBndnwQhKL/QlDTNei1KV/+EcTMjkSp5vu0hQMWZCYRqBU5635ZqR5ubgs
XndUPHSvr7I3lXGzx86DG+lDFADKqZPxUBJVj9u9PSFEzsMn0VNmPxO5iqv1qYFS
ww9gbG1By0lIku9jJwCn8HOt2E+CCSrAtJ080gzj7B9AXY+NokpqkRCNVOov2kY+
5SvUEmswDFaqtCsgZtH9EgXQIv1V4ajh9iqEO5dAwl99p2YUq8uIFFIFEChUIriD
o6WkGeyvIfnqBLxcW6HGehI1fboOzTd1gX/1U/jCNfdNq6ObwITCmo+IkqlsTIBp
c+zRdR72fMIJZPjRGL5BoRMysycG8f/Ghxu+pzGohaB2Xm+W3jgHCGwfchEaj7M1
p8euNdCaMeJ5EHG/gwRKyC3/C/MwESPQ6DQvVbYAz5vpNc84UDRGZt3x8N4kp0xU
+gkqotbBasUaYEg5jxYQdCc7p6KVu1YmgHUz14H2ZnreTtNSVq7p4R/WToXDMElG
K4MNm+ks8h4MppDupzmV6ehiPinHEvFwlOuu46/R2czyfK6Ke0/oePEWcjwsCmRi
amc0P8x0HjG3OjCBWJafvlfSzAz9XPRPQLzWceo8VXIVD+iAqG5P3Oi0u3sJOSav
6AtMg5id2H7DP9df8T/NOFInhX6pcqPmLQUKaEQ4p5GBPfgRBGGInTfFE85m+x30
FdA5n5mdaPDjogwtPCuGXEk+FcPZyf2qDNvwfzgOu7IZcGdbcmLdAT4cUf5N6W2h
f+GHJZu3+zdy2mX2cCPNmGxX5Mf7fIxtcTe6Vb6VziCFPbf7A9KZIqHT/W/0LZ1M
CF7FKgDd5FKrbJhvObpeoihHphNp4Kp8ER7waot4bAK5I3I6wN3zUIxPP3n1SnKR
r/cf3yrTaabAqbdDbDts3uu2qnCx+UElHMglUPNXgyQRsDZPC3sC7DcaXbLvcvnJ
+AYPV3sPfG1J9anjLRjprFgRKC315oNYdUw7fxRmz1LzEt3B53Xxq2p8sf9cE6hM
TE2zYCwTg5w4ko5wJBMeLIvBUGhw0lThhc+XjpPJ4y09rvDN9V8/k92J6xaukaGQ
h7sHO46lXnIjAY4KZCM0u/QRrGeBYGc00Np1vr8X3apZNYNzpZ5I8idp3+0bzx6q
1ccIMlbH1MEc/O2I5nT1J8p9LTOcBXiX36iBtYqVEdpQhy2Ffib1+8JyVVCRCKYi
Mw4RxONjE5T0W74J5lwqiQ8gXb+Seo5EG4YKo9gk/k8dZjtfe+tvkmiihnbxz7RM
07Nzksl6anOWOZQ12Nl5190+K+7yWf5m/z8f8YO0AJEkTR0p2lo818CpzYmFtrOg
sw5LZKLLMYF0uHPXVIihoJJTMfCnVMHD1abcpHKEWd5fAoZuQE3298fcwkXkKS2k
dkUoz6wsvvNo/cYecXn5Ye4QBkfX9m6h0ZvRYawyEvkHIUCguL0RyQtsNkvonHot
eckd2GCwSSqnxz32mOlv7R8TVTGRVGln/mOpH03b5cSchx9sfKWHeriALbhItTI8
NS/Pqlh2gmieDvXApn/zbAs+PlDOmL9kGiNPDXnH2HJG+/otqXKAbklDEh7w7D8b
QHk4+35Vaqwno0lbsXCEbOQS8tdocWFe9bCC5nHl2FUlYFiSWfU1QH0c7edSlmE/
0b/ANZfflW7wTBMwbeqhqfmnooD9Ardj9Ko4VkOCPt6ZEZQy9RkFmE+Xjv77PP4n
Njeic8CouGlmk8ihLrpaUYtswa6UsZNVyxjmZPX9V48gSpBi08Z5lICTux0Dcewv
Y7AMHw6B1lyC6lcMv3A8xh5UDMyAG+u4pbQjlzZ1yS5ilZ2COU0d3il7OPqJgjTg
3eeN2UDryZBr0aBnXkwha1hwAzVNZmvsn29btP2gMYmQBGFZh2rOW8UwEM7jiibo
AQATU65fDvhVv3f2jDL2F3nzYRJX3x1pudDpIswoVJ5KTO96yrX6ER4pWk1T0cnK
pzLr3XMzA761i2R8O1T+nuWEvpH+N7qEf5dftn4v6z0RV6TrSS5egQc0WXL4nFPm
ioju/rBqnfwVwCT3RzE995wjeIwmTL9chg7caKhqo1V8UO2Rk8XS4fi2rEV5tkQ/
x2r9m5nFcMnfVHFWHKfNhMTujm/RF5CdfESCYnrMO9zCozQxV4XS7pISvsHIcfFS
7j85lWcg6PB5K+abvFsFmtCkd4HViHcGdH3mlY3/zfdsudsdRIyjL94WQdIa80Bz
V7p0Zpx/inJGFc2sEsBUNSsUxbNdpjEM0xm7vE83XVXOoflEJhUy/WBWhhStzqY1
1CjJa1FXj0VTsKnw4OAo9wVQANjBBDrYo0JPjZUShRmhTEC4DeaHcHSdj1NqKC0F
jRm4Pd8NodGU2FmjEYL+lXgDxWe9snSHQkQ/gTyA5MvKZWaNcM/+qHFzzY+hiP7f
17FmducHxImCmI4exO3w2NPAwly9ZKyB2+NWRoBveuIYsx7AEmKy3qJvfFz8uYL4
bbXTE1mNO9BWbOtlUcXHYEhp7JcJ1jzA2e/Cy90dLESd9Dt2Jbz8heXzDS70iqXH
DCh7SOLrI+YjjRP0fxM2BaEIibeu54w90er40B6bxLwb2iKjmThUQU9AVr6ASlNe
4XKvlHQyn2le9TquAR8Zu4chyHSXvcjreotisVtv+xhaR5TUO0eZbzfdVTe0KR9H
T25KPJ3qFdWQLzXRceHTz3oy8LL6fVPAKox9sstc4T1hqzhUwuWMoi2W3m7J9joT
HsYJeOncMKpqgFVWt5idnqpZoYs+a7ziIfyf9pG2JONcHUR9dKXy+Quhl3GsZJNK
NbqOsWZ7wMgII/XsfUt8urRvCYT8+ELfo8cM+a/CYfk/aysI4eNI+29pLRennLzr
qHX7qHymU4F8s208ZTHZshmF2zdYvt7nshcGuPT+gd77Jtw6CXZnkVxoStvsGBMv
meZqHSk8zogPk/bx/DBRiQfU1lmHfPZsw9hfOrT+k75Qly8gT9Wd6wONXtZKRjG+
LFbsYiuCKl/5IlNRsr53sO26DzMh17KCgbuHPf6NAMBQTNtrIFdBUjLwfClGSnMe
jvqUd/O+wBQbf6UvR2MOGY/69RZdQpz27D8Emic/I3oW0rlnfGBbyMaRJj33Mz3X
YK7WgGBXcrm/tDcYyDJXKsb3CPAgztNtee+9hMz7Jb0k2iFBvJ5Goh5vx4FIt9Vo
UUMCe/DiOv7Bss0jJX1aQYHtdQqWtrzSnVGjhUG2JtYpSQfb5rfZvqyPK/6ZTxBC
Wok2SwRSQUxKlOrcIq1F8BzSBtg2xCe92zayjADXb9P8ga3+OiiYRX6ELUI68VmO
WvptJUbo9/pWYqJtFJ9w5+sfWU0zZkmOflCfiTOXyfERYDwfs/2GQtUK65SfkUmm
GnVeUWKVOuaCi4I2JMZvIiy8oStSXTp9rcQflFcBk1GIQFJ6rClGCrJRlURY5aRf
oLI48nXKahgSxxMmJX9eAjP2M7mnhb6f9Je66FxY5Ytb9Hy9F3s6t5q3Mue4IJd/
K6u2yK/HaM8zfRpZM6JAn5LvjUgSD2LVBCBupH7DFBDXg4zzHBy76IwGyQkqg58O
AqSl92q+FM46lk5ZlCLCnYozN84sM7s8eskeMuZY5cC8e3eQGYC8VZPsvN+zkU77
hjpPzEJOZUTCK0dM3rKQo5U96OQWBu9oojTzSFcaUkiFoHmCVcxO3T/tZCJzB2fe
Icvz1yg97qprjvRuYi2bkSWINwAM9J8iF/BGusrFB+bPehPvRCZyapUDseBcwWrv
ICpeMYx1PKlNwqKTU1RbYKmhMBRrM42YidONwzECFeXPBboxFRC+pFbV6uG2XOzJ
5h01yGntjCbUpsT1ZHG4MXKMwkctnbADeXqm8jQmq7cJkeX/BHGOZt0eDdJko05C
St1dw/uhNwYG3Yklf1QABLmNtj+d7CMnGUsH1UtuLrtXuIlDrSMA/OEJVqHFD7/r
eSAO1W6nFRlX8pkqSOsufJxSOM9cZogOkh/U/m1TqbkKn4nZVpVWiCX+OliMabQH
jz4vDUuBkpYNO9olOcr6vRs/vA7ajqdgSAwTB2COk3m61retj8x/qd3UDc5q5AND
mc5HpZfVyZnmC66KUnyHpaz17eYg73RskMh8lsN5+iuxuvKabI3AMvEaBcUwDlNL
twtbpgIo7H+sbea+vnV5V5v4iIFRRM71gWqytNgWjIJCx2oVWEtb69qxkncjHWUe
BX+YWG6A2z7e53JpMcJwCLYvHEp5W7Pt5Lg9+cuSv7tJOM7lQhLPBJGtgOA/Lkbh
+NSLqWQACNoQ4frH/oW61MGNDKUjga68CSEPXmu/dbqvjZlDpKIIWpPYRaol4jcU
PW62x2Gxk1x7hr0/YKxmhsm9A6615ykkE3ICnQyPIapmt/FhMFluo3LIudbEsDbw
5fj8/UG5T1bf9K4e5mwBg4w0vM1NGKwuJIjIhpxQQKusSpwohAQZVHHhPoWlELnY
/SX9T6IxR1pKV1C6aYXm0/yjFRXJi/81itUuAAoMXXF/FOk/DUFtPYi3FJB33X0G
zbF0fyfRaJsT5DzHQ3Kx5N5srmzpCwD4qNIjempLZV5X3DGz50FmXaomSJrO1cgP
y5sr9wxWrT4tDTaR8OO4UA4Br745yjKHafvveFn6kVw5fqiozTxVhtB9bsrtZfWs
xAhJzO3QOmKo3jKM2wLWH6EFjUgQvOelct9pEgzzgGBMzOIF8xyo+Nphqcbzy7wg
KY0x+FXS1Akxv0wW4o0wUsdhgOj6LG4HfwCqOJ00p9nN6XgppgsaBhJepw2GZeMW
yN8jHWtQETVkEaoms3h/I2OjTVjBXeMmSFahSnaxMowK3QaQ3qBV0ZqlCFxfYXiF
nlAkhKy5KEMe3WnXMHcqceheKj/+toi9AExDe9qYLryocmxjafekwQm5jx7NpBY1
fUXz8qz93OCMx2NZ7+3T2Q96He0YsnkYkM0YKaFlT9um6rGHntvh8vdG2oll9jNA
uiahF5aZ7wbMqQxs5yka2AMYBF3ppF11PprYSlSqB0QAFLTJCqs5kCGfknDd8ZjH
LgaQgQLgWh3fMET0OARsp0EfBpmnuMBKJ7xRTF2ZNjkU2x/HbHEQEBMSqDTUM2oQ
vqANUYeDakJcBndyxpXE84yFqc12VPFf+05R/FxSzQSGBFhUJdjPUhbW71LXPYSO
5cnCcI1VxoaKuF1m/gGPKlUrqq29Z8xthUtPcQA5nL0aOgP82doQjw9bz3vKrqrI
jikM0ukJr3zOUGEZQ/1HDrSr3B6+RGYW66lToqKagVS3NUASgZJrhcldrbBc8BzK
GBkDlvoowRzNx9A4b8fha/IlgVgwc4vVIgzUqjTWy4RBEaQjIhoS5J8r8WhFzGTE
DpONa5A8nCjYBqRbYTuN4jOUS8vOXrIGSvLWA5XmZ86XIcvvcyWAR76IJm2wUT56
zXHf1ZpVEiNpSq163GAuKDLihY1PRoabDYBpfx8/yK/vK3iPyYlh5ZtVQ7QpuGni
kKgjj0LRHaKmfOckGKK8D/o9ETC9bwt4JibHaIfBkbyi4gVW5+CNeoX2aSCRxMT1
VMhLN1qt+V7FEgalJxjELOEwOrn1V+cqH+RR69vzyyxr1KasZvAHiSt1ZLogeKe0
QkOeC2FdoouGWY7SXmdUmPa29037Ubtn65PVq5ZZrOdw9YEfa7f2KSauJiOT3kwB
VcjrQlDu/oT9M5G97EbP+W120zaUm1/8vDikGVZG6FVY1kp1fF0flHjbHTCdJVcC
55uZ2rRSPVD6gTTcS2ypuJ/S0HIGpPYmfOc9aaOAqWwFxhlfZ1DF3En92G8zPzWM
ZQcwyI+fR2Jt6mMw2dx22zvbS7JLO3uYYdWipN+8OkFpeWnTpelWIyAbsE/ncKZP
B18L5LHkleZNBHd/5eWdhM4hU0Yhaz3IBhjfg4+bOwliyEu9W3t4P9t9tr2T22Ws
30eg5JgLKeSemiRRkuZ0h2ArVVC1d+F7Kj5M8+eiWmdv3hJlXPOD8juLH+dNPma1
ko5VeJ339yj6IRGhbcza2NjQh5QnldG50sBhRYs9fqYlZfX/4vLg9f2nnt5YS6+r
tu88QI2iAvn60eZpn6ZBtxytOUC3mUm9bDTUExMSS7CkAvTl1OqHHhzKl7OAVaYD
AirMKtHRG8d1ntUqj6qD4fNXzN/92RA8z5MVIbax2J9rixhr9RxgQFu4N2ktakHH
prI7ufOMD32ouEHthP7VQlT+oa02Iwh6PDlg6WvZoMHIsRgRZ5KopRS3ENjwhBP8
KqaxoLdJFr5/rLzPdmS+Akx23Adu+/VEUl2hNRydwMLAWBfWOdQm3GRWoRhy+/vP
vhneEtTqpKyLyKKRNEP7WYWxKc0ea6DIwt5yBSAHEocqam47vMpUfqz/ff4t3b/e
HM0W7SulEBNJov41HMEPJvqQodpDRdtZaNLgEJIgysTZldhK71vf1lVSag9qz/bB
cJJDVTczxIYIXsmjT9pv16BAp58Yc2Y7JK8gviL4Wa5yOwbMVMSAmqi1szN5zAnf
e6VXGthsTTE/Kv9ZDpz0WmfUBZLF2EWHMWfZucFl4w6N8HdGRA+5yyNxQbOlKDUf
nDmwVQgFh60vItRu3ehdFXs+drXshHz9f6aPvb0tuqIALEDiBR2UL6LvcVJlVu98
Z8xY22ODSFhGBUwTGi9qUnYAkPGtFbIi+BAEZi84KQN8KGVOnHGsWzhDUwgKp/i1
8CXgkBhKmhucKiOC/GN/o005eWcqYne6qgswnCqkDq65c6aZqXYc739kiISyMdJG
76bymuHcCBOSzh6HY/IuI8iYZO3h+sSvK3JuRisQALEpSNc8IL9B8jWAGK5D3RNK
R2vcXG4iuCuCukQhxFMlLkoEyLxIB2Kcva10h6jlB5Nor1RHWIHl0IRDbk2RfiEc
RBTtcCrdhhp8/b3HiGiTthO6lwCGFwPmz0Xk/95R5rbRLWb5y+VrDTEoLjcXdsEB
3sxJFNAt52nnN8nrWB4yR9UQRCPDXOU8U5edAKUFIeyUUPCDLs7aP5IiJGb/YF/C
DAEMdtKZM5pl3vqPEeK/MG+uUp1ErbgmLNxuHh8BXYVsOCa7Y2KTis5evcQggvdN
MrI+dx9A8y/VFHsicXNH2sKSDLp4XrZWtLAu074xsQwJN+s+nrt7mGyKkyGLH4ul
IzBma46WerikUihTbp0/iJmYwFQpptEpHqZmxbTr7qxTTFWRYbFd3eZNVhkfJd0B
3eoVb4L2ws+IagtFYnFaFF5BvixwK27RhhuqON2kLNENs4PPGcam3ruZa+8eof9z
LJ7G9VBUDP2Mr42n6Ko6tSOWqnXaDfjLEieYoirqU+FAQUFxkwXoqiSfF9Ia5+XU
Lif55Slckj38lGB2MfGOSOw3o2SOnBUC+ppJrjcWRgc1vmgG5qiMAiCRSe8E5ZK5
xcbgR1lUsrLkfum8pWQX/pn+AAQo8pjFt88OvHDzhhUxOeJ6zj1ogyJPCJLD0Oh7
ebFA1OT3M4lpDhHu+5ACgqCMiMtAGbmNyUIsEl5TMs9teWQWJ4vQ9K9czMOZv2/Z
3GVAUwSr2KDrLGDzZus5+FkTRP4+F3G0URE+k+Vuu0d8q97exyT6a9A/fP6dpxyg
UpZQE6wWVg5bDoDYDFjhZB6GCzLkj0wbURS5WhJZkt0p6udBRguVNNbzNYYYXynI
P7msV24tBFBQeapUugNuTT0fMxqEFOftnrrHxPtHEPJgoFxVHW6Fmt2CZFgIlcpt
IYb51swL/IABk+HK18/JFB/hXyCatptx+xYiv8xEQIJIQmplYXHbKba9QT8Bp+QK
Z/IoaN06ggZK/PO8LUrqgHMMeUUOryBDZxASJLLw3co+yqN0j7W0qe3awZP/CWij
QjTScEjeZeBQxFTeJveSqscvjWwDH7JKsPWrke4MyUcbnejH0x5aKQ7eHy2YKROw
/tMOCHqNSLhDweneYYGGGdp34rRWK2nQsB7DwSy3g102b1yay8Rb3Qe2DUQ31ZuC
I+SVYII/qbxovhUSzjJ4Unze65yEvoLakF/8KhkIUZDepYOGWYmQlf8ZqTPkg3ZI
DvA17km5FQZ2/B76wF3LHZmK1SY+kGGaWPWl/49a0AAbCtcURWXScVyw4IYi+D7y
jOBWE40witMW/GLrHialZdQHTbOdlo9eRJmQgQ33X8WG7sUgod5tkFTgDizgk0dy
oD7KASjtB+D8GYhZC3tw4mz+jUTpM0i4JSxLtpHhVzAYmNAgxwH6G1nalnyL5QMC
4NSgrLW7Zf9jWkVKbPK2CGEPJSSc5k6MzaFG+Nxc9131B0/p/M8Iq1FfxFKaw32T
UEfkcsf8XcfEt6QSBsdijZZhc+v7js48y1mmeitD33K3hMGEheGwj80pwQnaxHOq
i9TnzV/a6+ZPkHLrkYdce3QAbgspus0fOCtrIMiKZ7G9w5rbc1HJigoHsDG4UoNJ
gUTHbdWjSJN+A1a4rWtp4gBCDLwu35BG1Dv6lZvAGoj1+NvHJw4aaNxdcAmAWHmz
4LuV7/vJXWMWf8VIZci8aKMvMDgzAQcGMF8Teohs3pkHYn7/Ah76+LHxBYZ4EgYo
NSW3P/Lv8tprQ45uPHS+ostKVh2w+DUBmHJeoHPSFFxRi33TR1ri6lzZ9B4f8pWO
4PmLJYQt/XELAa0UJjmYVc/yyDs8KQWpfHmEDDGsNd4Wq20aRyslauJNwnhODdyE
v3ySSyINOIR9w5sCt9yGDc875sqju0I5icT3GueSKxQD1NvpuRQCChXafXJ0n0qV
C0olb0vdqVE2j0JWcZ59qn4ftVWI1MTg2OnTu8fwg5zw3XhMChuVaMhqpDW/yG78
beMNCZXr/IeuUeEq+RuuSwcSUquOkX3IQwibB0L4ojCnmQBkkU8yi83AaPtGR5aO
TXDcII5iRLGhyBHI3hxTJZa4hGNPT7LAmMa5ZLvjoElnf08olOykRAi00ne/K0Bs
r/FXgXFnllojqjOy89LVnq336S7MkBqqd9ZayKkk2xBzjZuGYWE9AMqFeTeH/IBT
m21PnaqPtfp0dBDtzkoilnARleyiXh+1838HMY04hWnhVSZg65jAC2Fj4XMz2nPq
zpOxgJVZv3b6FRCpsDtQTg2FQa8eiDwK0lm1QTIEbDfO8sLMI8UL4ghMfqBfZ2Dn
hD4iWYL7Yyj5IfkVF6hPDmCbdL66gXPKgOdD5I5r/gXnHpn90VD5dvjJeATgcYoO
ieEvGCFM9Np+GLnLNlBvuoWmJRy7YlJwr4Ki7XrcccLUGRFoGc58lrmInS0pDJEt
G5cI6Ydfy2Wmo4k5AxnOU4NWwuIBfOTVjqrwRP/GCIsqSMXZJ2vneqDw15exFhrm
mIGL65LBPkcHTAMzP65s1JS/CnHIv/y2g81j2oj5XnG2ezFh0gMWIK2jiZP9JysY
9NOtm+uH4KnlvGuE68fmC+tR8TIG7zxxZE6uGM4JIPxuXejQlTe9BRU3Oxt6szMk
IevZ04hpIjCSy0OvG1RJPkvsi8krch63S0/PVQWKU15ErSMfxVG1yG5gChqT/UTr
o5HiASwG/h/8b2MXKRf2LYz0tA6ZnOnIG0PASal5EQ0jZTzYBd8w65J9Caz7Xtb/
GCTfmb/Ts4tMldh/imAlZ07FWQxYQ8EmnE7bdTH2uhJVKp8OOfRsfD9VH1kfXYPB
0JxibZtVQEhpKzDmZTXxutA+QlPDHi5VABDyVtSDVTe8+oxk/7mokkvZhI23gzVs
UfO6MSWLh5t2zDq83qokfo9usj9qpY2Ffr+N1dc++rx0wBnddGq0VufitOsPFq8c
1TWAhZdqRM+bwTclvW0royRGc851cUiWNOyfC9UZne37DSdYrDH0AiJOz/ZqcRYP
4SXzp0ryBxHDu3oPhOj1zDzMdDro363JQtnYUQ6p/CApUA8k8uX5K3kLDtiCZLYE
GOV3Pufo5gU29soVIy54vzIK+ekWRjrXWMIcdyugNoWiaJG0Tm4HMiv4GNgI/kpn
ZdWn9Num8CmlQRChh1P0HJpkbJcFQ0d5fUFx8ArjhRzpGjiAWVRNJpSPLaBk6wup
2Ae71R6KgAzqkP5CPhPaDXjqsj7iu+D7s11XD4yKTuB2cpDc7vnYRDqLMJEnNFzi
D0dWYp4wx/zudZepclSAV8AtVxqgnoHrZyAse2/S26P1u1HYevLxURoC9IvNqRsL
A7xkpE7b1k683nEdb9ivCoV7XFZaZ0MirOvqctPFKDmDMcgI5ZNwXZEMA6AYVzYg
cHtdn7SeBF6VFBCfFy2u4xkM3cQi1obl8YXCcrn3THsOZP14nSDJvOHa1pvbF3ul
1cpRVutemeu+kZFXQTQa7VzEjihbxSHYKaDLOpPjf7B3LXpA/ySZc7rMfisyvP/K
CGHea5D+gS8zY5SsUc2CkQS5CCdIrJDy8ACohiCOwb6/GbtkbPuininfCZ56Yz7B
wTzBDmsHtOymzFGOzvSDJFh83tKhJQmq4YxVLDno8jHc5XKblrgllY3ysa2ve/sx
lrjoJNW6l19za1F6zg4lX+1GKzcKFLhzC6zXPB9C22v0IhpJcVUfzH+jxvk+KQal
O1xQKdi2tYflINIQxmCaLxTs2caT5HZbSDeEBIM4c3YyfxJhz2T7/ydYnEVOyoFs
EYkgqEw8zAezl+iw3+kDr/oQh3ufsnbuZu+1ysvlV+9Zc7fZGAKD59u5gOfgxGGo
dX6yuE1b/NcA8qp2R2CwjK0gnO2aXjts8JwJ/eJTajrDlCwGYwonLIyQ4miCNzOA
pmi+4LON9vI7heREJ9UbpJOn3AhQVJ7PvcM7a16HCh4FPZGEIrMOQjaJtLzHPeSi
Boxukv6+/mPVZd1QajrufxfY/XlJQHYu06eeZEG+PqWM9Sb094pBv9FlVFDR7M/4
MOeCoPjLiFO7cdtnmfUAZvqNcPbDZ3WEiYl1rqxtnwWcZJ6Evpu15IYuGZZkXHc2
xizGooCGZELbNRItxaK5P3HOG5zUrHJTX4gqee/sRXKCTJ/Rvsg0U8freT/R78Dp
KWmY5JyjT/VAlEJYqmQVHfkRPotLclCdCFuvXWxTcA7m6iz9SXx26LTtQFmlBaOg
QWltoqdWk1dWaKCGjEKJeei1wHtRvKclaFY0HrAn/ppgO5EHZYbgso3zS/GYlsLn
bdhwmx2gufuxFefS8L2EaM46408U8faGYI9INBDTmztBhCpwn3rPCqR5MP3Vuzbq
AUiE3T++ube//OWkxUQy5qhZFw47Z8SKMISKiQ/iq/OTar66rpIWSa1oYNY6PMej
wJ/rmzp7+um4NceE1iC/bt+IRXjqUjhyZB4kE129QUqKPmb8hmnZRdbkJexb4W/1
DEjRBe3vwN/OIQeq3squT8Yl7KWTKqQbUWpJ9M9IejyGKcvcjF1BiZVd+20scq/o
NMx0x/FNgAzCHnIw7bEMomtjHnEPZBMOORby28hFpZf+n71yeYaUtAzkHw7XQn4M
hMBi7YmMjx34BkvCXoV5+y8TZux16+A/G1S6Zwe+06UWb0tb6RijK8vkPiD2FR+a
PSVKI1XsBb87erHzqEAermX02tzol467FJ2VGVIvN7X/L5vXJUZag2//NCJv+4Li
VhuMozTOYQTvVDxneCDIVlo+TKVBquYotS3XiVmWN5u4W9qyHNa8OLgy8ZTmSE6W
oGhsACQqPePSY6u3UyVoToxmQzV1zCPMTovb8f3RUqA1rwXrmfK6YCkQHgJeA1SE
nhM88+A/DprHd97ba0UHvmzVvK7/z5BYb3wY3Ak8fsOmm12RPAQcQj2w3hww2RU0
rwe4GYbmsJ/maUi9y+qWFYJTFGeinVyyzq+5sSd+Uf4NWUmnmAe9C/QO5IySEDNO
rgOi7e/QmebGL3hkohJ8pDH2ilGaZkAD0g2rUMD7Ps/VKJRWinmhb2UtDVynZ44l
TlCz01xL2OdmNeTT+2qQ71k3NHeCoUpCGct++aacWWOHUD1di7bBhxff+BgxnF+m
w1qUX6fCB1b8rqYV/Yrvbxtd7kQWMMDz3hfycqiBLSgLaD7EXWjmdcGroWjtjPHK
CtrIYmOUKJtlG/nTpZYRFgXX49lYQu7ze3OXOM0T68Ie5tSlaRUiDfOPM8eekReH
91nyq+8xxpN5bR+ZUD1Of3huScaA4Ui/Ne+iIWAiK8qvoUv3sXqoWLMxmVt3LArJ
BXTMkS3AmvxaQoIrUFd74gyJ0GMuB5yQ1wXtIvFBiP5buRnLqNax3UGIWLWcOqWA
Z2LD0Qh6s4IGya+G3eqO8n8lKZW8D2aSpkHZhaCFdvMNxXjtIbFrKW0M5WQff1We
expycdpty2qn10rZpY8wnD13EvFdXz320yWksxosrNxf+xWIBgtdsvH2NwW70TZ0
wGK5vKs+BjrUuQ3sEcDFhTCgmzdE6EaZBdWLpaC/8y1lm5fbZNWzCshZF4O3Dw61
ioELo0iHhOm3G36PA3eaODdQtO65Zmv1nctIyzNKhjxzrVCbefv/ptIhpoOsnpHl
gk4t6SzMSy0lA3maM+kUziEt24dd0ApsAUJSh/d4F7Dq9L4cXGBvJZWayUDTZiB+
PMyORpjoBEB9TgZ5LKspjSI6iiRQVDgWgJjbW7N0S/w98ZgZiHhjMp/oNANmV7hU
TrCDOqQQvMZYtnSgvr7zGfPpIcHFq7yEndEByNZg9tdzuIbQBj508FfMHUVFkS+a
xX219WUFxnJeTydCjkocVqtpk11tWsfw86YUaZMJ2yjREnUuDON0hsDpgvXwPub+
lfNEUUGWo3FozaUPHkW1yz3OvVNKjXZi7uAVWr65AbZpbyka1rGrZ2k/adn6jHlE
06gVEBM08Qa3ukp1qgASkxf6Czcu2tL+7SjLQJgwjT7Y7kChOu6k4FiFRq5sf9C1
djlwvS7PbV5zLn+bMGJeU03c8GkPoQjbm8RV2B/YLj0j0JQ0Zaje1KPJAdmInY9n
myWQafZAIkOpqfwStlMO6Tmjn4Rr0afzsP7oljlYUDWjYJvxH8g/3NrcOoZeLhg2
7QzT6stGjEjs/oUzfLV+ilLCMNjt7GY7m1yJi83GEnp+GNXPTaH/z37r259o4Btj
/RvJ0OqOzA9kaNTpoVOhCfek+ysFhn2uwsMS1Gkp7elojltkiggkRyTVE1irHdtg
4yL8oQPwcM4+TN2kuavGjOEH7NInfz72E3ViEC9NvyldG5VzuHGndof+bEK2HaAc
OcnI1uRNkUCOcEewhc2BsPC0dvnXlFDiRZMddPGDgeSd+59Y86GSXbsIHI7XRUHH
d8cX3uxL0K0pgq4UdagKZaEDFp0wschGT7FIcxeHluZ952w2hZA82tc7RZenFjf3
ffrWktxrHBR7Kq+IJKReW6y4r2nlJf9pq3lQWr1zSp68CwJZWZAbNl3SBCyTuozH
ZGNTTbYZc59ofl5NV5d0NhwwIEsp1cEjB3fZGTgeWS3uCYvzlw/2yca48ME2/0wb
ROw2Ktf2rHhuruzoajlBb0i69nlzs1e0XxnYLv1XWJo7J8h9vlKRXRsVBcVQKJko
VpmNol4nebONdKOts/3H2H+4YoqZn641tDX4F+uleLs5vFJ5/cYDF183PlXGiyRQ
TvPoOF1E9I6xoArc6pXj4CFW+rQOfV0GzZfXZ4a+u1C32Ydg0pj6Dt3SyzsyUhwj
omjf1opEhHwENeKjsI+rjDVPMdW3+i7RziLg71RBoy0Czs3Ykz+QlPYT5U5+tqtt
9PWMEOMn9sCUabdCcJahuJP3f8Cw0lSL/jFwdUwgfzrQvt0Ux7Y0PJ77lBCzagnz
G4LtH9quBwM+pIDb1U9PX6TwVIkK9OagmFqadpO6si36exkpsLJYJFLtnQ6dZufV
y9jp1z3Z9FUlUVDkGucj5CDYbtIeLVJczzpWmyr1exgZtNxlfRGTzQ7/cqcB5iD0
EC3ptbs4T1AH2LNEsURyHnP3vdGXlWLHYlcpqNqmDfiR/rZYfnyec3ZEuUz6aNzw
qz2euptO10vbpzcfyrASS8z1T+SL881/J0JyZ5PMzuNjQlrpBvJJl2AYbu9OKX+Z
IXDlWHyJse6eEHUrh525SvaJaTWYPR2xc7xuIPfvZYYAKwfyeVJ7QPw0FBaV3sDP
apTsYZv0Y9naNpktfEc+vrLWGdBAp1dK9xWY/12AJPpshHZNhbE3njM1ETjql68m
q/7S9PXkjpiizzqmCeTStT58zEJovV7xnhQCrjYfvFGpjnGsbMBpXaULlm1Iolna
wgT+q0iTzTk7uraLyuBhOuYNq88hGPhP26ej36nJ6j4RTAz0/iK5OoAqGzWRXhGl
JA+eTiWX/DM3hUUIkgg8/awKtpGeKy8nWRkkMGwN0w8DY8ZlyEVnpO4qIgHTtNrG
h7Qc4GNpr+khFQJMjYz8kxBrJa5MwaicYmAXA8bS37wSB0WYGSaDMu2UJi0AUl6i
LEorWLBxHqFcLb7QU+VXsR8ecm5HV8Kfc4DUu/GJfKK6pEA4mFR82jvYUFXU1I4Q
IkR2he+I40GjV4ubPhVdACjEaWSUmyRxkui2c13chUvi7ZF9+sJZIbvHaOiSQUBK
5tImw9xh2IPG/g6W8bO9S6Mbw0+sPmNealvh64ki8WSQQz7+iNAN9x8aVUIb+aMn
yIpk6re+lrKKoU0rrL4g/aRPS0OmJmoECpkJbBSZpIMzP5ClzfNsiRm81kEE7ngE
cbarX7pDwtxt7gl5t/LJ1vhjWSU8NxO9x3UpL001Ch5fAotOUlT2HgxeS7gO4499
hnOx03R1fCMCzJ87+T5n89ZEzPNQwxcSGMoqoL0iVdZ4BzxXKl2DyUvGDrKJsaCE
xPWFF3v5RezKDms0eKsCeMFeks+mzVy0Vm6sLgtv/g80HShN6iAWj5F0jOD/i7DD
+7RphyaIyQJxWisi+MM/BcwFE8J6oy4fGZE1mwe84QWvHpHEn0dPrVkEQXdTjaW6
qgYh4zUj85SIqtm3+aWJKTiFonhP2q7tiUu+mtUZEs6q3LNY+D97iqIeDw9TXGuL
+xVUbXRUs/CQZVzQaR8u2ZsHcNV5rAIk5YhOPJL9WGD81SeMPetGIv9qFSNADNyU
OM3Btqq8ZMD/xBQgceQcEi0wzuN7B6alg0a1wDJj5O6GIeZ/NAUvu1AhGSTL/7Up
rOqsZeQftu+UteHra8ecWVXStB2SnNRI7boqQpRLq+lHANyYQkWJ6VVbgXTOPfgp
RdvoLh2sRFrg7EsH/Gs1/q0pdRxLFyftEyjZ1+dz0Pdip8n0cYP6e72Z+B/CdDK4
ZK+No4TjXFe2O45IzEHmvJ6ANDFk9IpAj9XOUvgxkDw7Xe6Ob5sgphoIpottqhQ4
XSuIEkMhVuPzjXMAvNTKxP3rYGjQx3aXFzsS9Q5CeJ1rwr1abiZQy8IAsdY1RSDF
gU4oUAqETrlNaoUrUtYNJoNp8M0fcd0XZJiT8saTWhBz206U/KJesN6i8VdqGwJL
MQ99Fo+Lf7FDGbnXvfGPY50PnCWlztKeOpv05aBSMTmQWfb5KlSt8Cm5TzIPiAzl
yp3LTXeSAta33Sj/yRjVL7IojopDsX4D3mw1JqP4sgiG5W00zvmI2fSTaeUQPdt0
0XdccTnljMMAPobTp6opDW++AD3lb9Ewt0aifS1Iftafa/T644bJDR7LDz/sxY7G
NVc27hlJ8/wxH6S6KZgVQa0Tno0ROQRJAvvK2RWrZ3chLzQUIp3yH1xp1iteo0Y8
FMxScocI6MpHfJ2NdukH/7G3yx0COa4mtZT0bJuxDraUHhF/VpXNDTJ4lQQNbnCS
+XBWPTtqZ6dH8xZhV0jYwa1oEWNj8T+nC3tjBqeKraZX0jRYPq302YixTtXd17IS
nF9DRV6KylxQ8oaOIqtzfUDE5OV4s+SffOdIJIn8cGXdq0W3C2XITFQbfVEyUe7G
Rxr6yhBZtd8R4GeVYmJzI6CJ8FfCxrDR6o/4+NczQ/iRzkD3gMnMMC+hsgey3eM2
SOEpvA5bI1S6vCDNUuEBYwKptR0P4tQ0q6iQ41agG29HsyeJLgJzUCeHlwTM3dBT
AX+wxoA4hZ483dwas6hgnNF4BJTk/oflB4W5zyk3/Dt5gbzdRLGV8cmV1QNYw5A2
gVXeKh4d7aEsrsh6P11aMIe6Zaow5kEHYtWiWwkNVl/E9m5KpBOk5kJHzTjisB0z
DWab2gA0tP4JJLZ7GT919hwbGe+e++eSCgRVaJ6Ehsd/fStWnJJqLT+746ZBjOgG
P4N9YrBODFOqG2si5aKAcyQhxWHTM5f5zpIWPBBX6XZNIriO72vSUm7zcyGPvpOt
c7hx/d0zeDUnLteqqdXJLUcM5XPbdHtauO76TR787z8uxRak9QoEqqaCBXfPGq1d
kJAKTHle8q9pqSW/Ip8md75IvHYaAvoj8lpho9KL/tef8dhTdaCEJzSv43ZFcZlT
O0Q5pgMg552yejgeTXNQHqBSfP1vJ6N0cTjwu9Za8S+fFQ/nrXDfGvQRcMfpQLtV
XW2ufhYBVxz5uDUpKFNFJp416B+Nvb/OQy2fbiyNoJ3Sojt9Lr4hYvd6SdCK4516
FdRrKSAs7Fe9lE3Fwfzdjj8keEu7YVCAexSiaCdDcK7FfXeXlbsIJJaHNR9fPE02
6am7xLRQyYmUz1VcEY0bWQT9xnh+HHFDxfXtbF9urjb0cn0Wrr2Tv4ynXj1c3DM0
veZtbiURsOxnUo8k4pROVNE5Xv545ov55WwpQ2xGxzbhIadPUOChmFyNxYsQHsGJ
CF6WizW6+cOEfoGFn7/jeWXeeESKyVxcO/gKfJ/G+o3BRsGxgT3Xfalgqwbt9PCS
Ho6tdu3u3GoW6VX8LfhxCTd0+KyOWvsm6ikctHApNydF6FtH6wcqoVIaFngmxF/o
cEfckHChbuHVj6t8xkIMZ3PdBmsg9xBi+GhftzJnvuTYOh2dWJ+AO9qBcvcIaj4x
4Vh3hufxaAgZ7T+5ZdDKLDhXogMysWNaHjjTui48dboehNkKa+uTaN7RE5ZME4ua
8bCaMRSNW7cTYFYkj/RSY1v1r7dLFfnSoVoj3rH0jzipN/oW6kqpJeWS3JNMgmN5
6tSX2u0qz9rw+x4QTsrZVP1otZplnKczWLnhnLbniQyhmcJLAkT5Zj5RXA3FIyr5
gzYijOfjSZYDR5JBfm1TgMrMt4kyqUQ9OJ+goe/EP35JLMyaGrd9E3AvgjLgRbLA
+HgrSbIXWqn0Er3VMMrL3t6ZHw6x5BlAtwjdp3Or4IMGZHnEeYgHkbp6it8Q/UC6
dyekM8ekk1vTSOrq169yeJ+RKk7iX9qeuSGRE1Sb7GxH8hVuGRIvMcz1ECEOHM88
VrxCNHNfGKBgPiquDp5mRj7t6e1nykh7zT5dHly+Hn0HagMaYoKSdPFdO5qAQ8zk
xVXhCwrsw5hd/ZFzSwMCMbkrbtAyble1a5XP5m4z/KNKyYtIChyLyNdct1l30Vja
/1NyFGdFgxpxiKme6FUnHWeJmxnpctdjs4kO+kanTkcW/biuirKrwlVXfIB1VHlS
x8JTdnLfPPjVmNOzJ48T/Q1dRK1QZtLkcSf+rQQiQLmtk+Yd7FhTeLrF2Tl+fD5m
x56qZnApa0LcB33ltLOcPSV/Ii6s7WrvZRCItBxw3LIffobxe1oUrXZE5rWD1JTX
Z7v0bTfcKDnkwPPNq1NNWXBzlpCbjiNBTWUGkBXhHYgrBt8tRlE6489mrHgb+Vbo
OTtF0Zciiwhe8hd1mGver6Pd4vQFFtcKdQepy/9BhWbPrB7m9i7/D/z7n6Jb30Ka
3OYdscZYg0KK+46zQniDfF1SImt7y+Yoe/tMIRTVa4c1VWZTDd0WOCtgjJ5XPRB0
7Dwj90AqSNH5qRrMZ4Lo0KD5tdF/o3epVnnnSxlYb9FykeK9o1xn1Lal55i/pBL1
XaiCZaUc062iZ/E0UKz6FEnPOguQLdG2F1/AshqXIewXKBW0YAZGJst5C4H+53n1
YrQ1CnnUOGWDHRvR0fMVOhOxDTR4d+WWFXdexNQCqqldAVOmD4YRFtx6OG4p8rKj
oVO00n9ra1wt2g+0dVnU4fhoMl83eh3aejQq04iGmDaJ6YcDjj8Y/dRhWVAxogni
71MHVu8TaFFY+XjrXym1F/VnZbblwjWtKcrVMLG6BIPP/viJfGvHYQ+ujKQXXSr6
3e0bhRUyg5r4jZNwGglokloL8fQSDYd444yGybYEiMExzohHCyKLgLfjD1Vrntu/
a3nu0oiyWg9VUX+fBXU/nEzvcNXdYAlepJHwXGLIpC21wNk6J0TRsMqi+a1vT2Jk
sYYv1Gt9+rcOBIziR39hNpRpqNh8R7x0GrYLHXCvW0JL+xMLTocJYksRmqR67sK4
LSJviHNH3mVULo8NMjM9tK+IJ72/jv2Y9OdY2oZQfQdoKb8fne0BuAaxZ8eWawsW
rqf6FIHgHC/Nbrx7Npr4ORtfSPsqVh5o0SwwJzl99n9TJC9kon6aWO4NdVASihke
iBiJRy7T1DiTqFOqF5ruW7naqGafrIsuVB/1caECGVzFCDrUe3RVbQkh99B7+icD
GfRiqNcoIIB5dTtxiK2JOKKkBEjeUl8MPDf59DxYUVOs7o2bSbpiTxp+iaif+IWC
E3wMibKeLexIgElWqurGcKh7TDp1WTYIfKlmsQNChBu19Fg1hai6AufdylypmvCk
GkLzUZMj2uNNrAKomS6FzM9XsgGM0wLtcHR84B0eL7WlEHv6FB3c1EZY6G6cfn/Q
96louAEYfAxKa6seVNAzdsvPKA/IWfGygU5EU/0BUAylSci6ncYrIZWJjlanxs6W
JCMTCBvCHONoJevEKovoV0IhKYQ7po3LkqQKVFOJmw9wL/0tDADN/cEMMQyoH/4b
9fL+HvL/zwCCTmoUAnO3SB1F9KkU4eDMpkqyfG5zG3McpblXPkBVMpOHJP91NtRf
SoojDSeN86A1ianngJtlYFwOQ3lzIHUxLo2xeVQkTFgmPuYdr+qmSJj1xFHxElGl
V54KAom2PDEt138KM0SKauCdkkJxVZYKAyf6bZt75d4Mjv0zltHOTF7e97TMTurM
FRX84SY55MsCBTdIi6NfC0yseG3FPoyqPd2NMhrzxticwcZ2ctzkGhFbyQvhfYI6
H77rCuA1ejbdLgVuOFWICJZX0SQt1mLifUUrn7DqhML9goWroP05spujDN3DCqMf
4oEHuojN6IjfmrSdWE2aQjlhq62dTGWcfdxYCzZAgYgPfnej6askGGXq1m9gOk2Q
kqCb6Hrdc8JQchRSLozbE3HKhtaRUfBasNqNvFr+s7AvWxOIDkOYnIzZJ/IDVW+4
PCC4yNLju0CoaSLWqDlyBlDyh05hXEwvYW7oWGQPjncfLAocmxIyAZzI8caiUCNt
9Kce6lrXllfW26D5ZM+TK50zydUmt+9memN1YPN4NZMP0Hnu0NvL2YV/PFgF4xlI
FL4fOh6WvvPsE/qVTAj/rrPuDrUoQ3CHiQpRKzQMWy1M0TvHApwHi6jl8KaZOoQV
o+9WAioe9eWdnW6NREGzSrQeTor3fGLB7t7FrLFTQ02fZDxDG/8bK33o2HfVoab0
Qv7oZd0FJ31caoX/jqx1tu5Bcved6IsvUiEpnXno3dW/ADI14DWDE/XPGQmxrOAe
Szro1UvRnvL703AAJ+fKelvD7HuI46X/QMdxX7tKC1K0eR6E+5Tv3J2wZjzl1bYb
SaephLJiPxESy9IF4JipQ221VXSq2GbwXvQ2ysHBaxOFe8o48/sUmnb5foLFVmpV
A/pTeRIIoUSHd890ZcWQd1+Wgd53dKNqp7cipeDMLiuwVQZP/UgU7QetzV5Ok2Kv
83w4JurqbJtUrSO1xvZ1iE2p0PhiNYi70KdSqWv3PA+BXy4PL+X7HCYwaFJ/+xlC
UJi7FdMpKS9YUXyT0pSfKD4LFL0UGn/EwSotuyVf52VcuuYNOYFqjrBC6UEJFadN
LZes1C0KLB8V68tZWBEif98IElkiNyvfoesjM2TGLzylak8pQJPbttzL/FTLpe2L
8bblJo10cQZa5Y5VRXn8nDnJrhd2arINXr2KobO/KFkIOWQaQ/7KgrXAqqLYOJq8
c4ZV4vlfSDICO4zs5/l+rVzudpKklbRuMcFzJKyySJkTofOM/qvbhRPZ+KumAlCj
gDkjReiMmeVQHnZEdvqGLObH8t6Gc8JaBuVHFbuRBzvzUfw4M3gB2UHFFXYYD1mA
OnozGvZCdHoZdGxayJT267x89nszNkQR6fzhKE7c0fXaSDF5lNQzcuD23avEIiMA
M1RgNdDMGoPtxeyrHKImGIx9xsdL8I+b8XlVd2Z1Z9FJL9fffB3dM0DCCLdvJUr8
WgMrwVJIGvikC6eU2qk7QYJ8k6bFAVuJL9S/5pfo3yRpSC8hxI061gIPZpe0b/P6
oJVtb7EJE31jfTiBoYxESjZ95llRhAYXjRgwYGFGjqZ0RCrBARKtJI3075yPR+Y/
a3SjewWlfyKdLi5CaTHh4q+Bws2vRtiTM1zMd+ycPG3W1Lj8ywXLqg9d7zUKseGC
Exgqkh4o8TxlJ2Zz5rVJ/OOo5QC4bzYg9Mejyd2AORh9wBAkgdSAZJycUXqezYvG
iaocZwXAzySYojVd6T98Nx4GSiqWtNxrZkF3fMOiL6VwiL3eKctpk8PMkAoOW8G/
qRdQd9MgPOsmaEZN7ttElMdek97JDJ7BG/N6+ndE3b83oZW3zQQpVnaNQVrvmeDs
i0bNO/em6Xg8uZh8zq7dGkmSMEm4Hhd4TuCOSY+Uadyy/wDXT5Btq5ul9T5JBYrJ
Gjy4DLbrGagFIwn9WkDV7osq2Hy6P775/ok7Cpt7MLojbyQM+qpzDukqeoiVlHlh
bCDVYewHozwJke8Q6xAMV8IFn0CnPKTho7x6vUFxleGqN2VhhAy+zt8A3vAW++aP
PkG+YdOCz1ZP9gZPv2iCNksfi2HcUxJh0HD+bllNd60TwQsN5brz1egF0t7oTnIp
veswkDay5lQ70lt8T4yFy9hW+jnXrBx8NBdxYL0CFqCwdfiOVCilnhzwnMzs8SKG
6bvaCL3sWb6IVGdZtd/9w/kiJNvEC+g415w8EGnS5cg+KQe07UgrK9+GzQszuAdR
19E+KFx3hpMF3sHutmh2YDQXy50LYOZVoIYWlUf0GyhEUTzWK2a6/SRsSBf2GVqs
33Uq8EqXMJD8KrU0m3YxJ4j5oOVrs9p75pzuej5xJ1qZ4Vdaxn0woyXr3YhxDogM
SN4j5NTAKuzC3gGzpwBB3c/BBzcx4f00KlevFfKy6b21fIiL7d+Veuj/WXnWUzjo
5MP3PbINoxq7ICMWTN49UHW2ADi2CrhnT9OWzF0ZcGeMnhZZ6DLxEi9o3vkB3e0V
QpXiIO12aEb3S4jd3uxSox/ImPDjJ0K7Q/O+r7SZ7KHrMUr/3Cir03WV+0MIfi95
yhIl8evzESXdvnBrDnZDKUzLK8mL0YzWouAPikny36jWgJuoR1HZ/bdixupjMCMq
CBXXVX+PzeJezvhhBV2B97EW9J8WdNrv3vOzmkrKn3nvYg6LJOc9Gi5Q5+ey5koE
afy7IUfV/de5Nd5Ji9tANe46eWZ9bisEPClRntgdIWopyTvbpnRzet1LRYLIp4IQ
mRlbANhmR1y+3n7SgzHWYPFIcuYaB7ZuC1a21GjLfKDJvhIPXADFAoBi68IRQwHy
CrZguyeGR0s3eqfvSNX70AdcNAZmPqq1hWuuciRYWyPrvIxnSm/ccw3GKZM7dUeL
flH2VC1Kf192t/QxpnFL/CR/7NwCQFCrhzPr17LErGZICiTtY64XHmlgWixE3+0/
Tx37yfIXQhSIZMlNEkmwSmyfqIEUznZE48ts3oCki2cu0TzUivS4zb1S/3Cy1Xs+
0vsMvayM5X67RJ3Py1VHo2uUn4MFCN7iugrO0S1Jej/DR5jREv5kM5+9TWjLluhS
KGlsmT6SXOnI2g3pX4KsGG5qNKrq+UUxr1KBxTtp8Cizrz6kaID6yDQ/5w4/Ddo3
Fk77+JdZ2DFsMQD4U/mlFDAnLEEp0XH50gsceG/ygjEqQHoS/4Is3XX45wAuQZiq
iPd5m4oFSdEqBW631QtEVANZKAG5R66T0GiQwsEHKFoWP3Oju4vTy+vkVkEhDY9n
sROmLgNti5inbUpNj4s6vD2XH0qjxD1fGV64KZCTJvoIDacfIcrSmbm/Ic/xD8Cw
1zhlv7NOgnDLQsAErm3l7UTP+vqTaL6YC2sxakMUn8I7gnXXPWNw3xHqW11kcOwV
+i+6D8aHC8k1uz1zN62fVQxU8NmJGjROb3oJ3ar7uAVjw50NBnEV1ftHiF7HX/6e
hmNbzi34Nb3G1nqvPmB7lA7eBDpfdazccvRdktbUXWdwDQFNbbhdJsXoCBM8fiqI
s6dXxXo2BUkCbNIp7InUYpc9jwBFjenN6wo+76j0IdcyHRanwZGfJrXizPbNwqg+
sxwdpPPHTGGl8etc9K9ZQz7yH031BS7A2vQ8a2Dxq03/Q0zHcMhv1p9UyLZnVYNu
lg9MErB+Eb+vC5G9dzx35uskEl/Aq+Nm7Yh1zQ+UwOoarQ0EogTdIfQwxd9tqnSL
Exwcyc49g1Id49eqmkiwTpWJ9P9nP7N6rDShci5QRHAVvO2PxvvxY0M3AcTvWprN
ksF/ZBskkN81PLclPKNyEl1invBfb7TgHiJV0J93sv9tkoKNPu9cUT5Mb8GMBGce
hB8LcO1iyMYTYtnyJDDT30Nb/u5cmLF8uTNR5wenk8YEThXvgWS2+xZVRkNyogNg
Dq9ZdJKw+rKlBDKDYX2tfIjWUXcU0udMFFwUjB6gHItIS9r2Q3sTTizll0FhjG9r
5Qos8YyKVaMbMRfT3+wkyC5MT2hgWlOOx7D1k541r0c/1KB5/Ce+8q6JbiGTEP4C
kjNMOssBCXuxZ0DqJIsx1bP+gN/No1zdH9+wLDtgz7phCMJvxSfz47zIFN7oYWFm
S6LVHlr4TFSIB7RTGQN3d34oMjIQAS5fequfeJHm9PdIl3zi2WqSxm64JPmrFFso
CXoAWrKj6R5q8nj7+SOUZ82tOa2+KP70ZKkaN47Nf0ire+skoqDf/5+PSO6bhEX+
ZUYIiFBB8wzfnzbEUT3HKkc9RFOUIKwNYYWuzuNpYIbmN2+RkaykU27QyAINwg9T
j+xEeMTn94SHexBNsfqDcfL6sSlBD1LxfFtIvGHJn7domPaN9HThYepqDTrGMIAx
RYtya8NVfwSqyCELJOOG/FLbg7EUvXCh7b44Ig6KjxV3DZ3eR70ZrkQCiIBNg7+d
rrP/LY1Qo2J1ksU/b+s5o6HG0w5Ts5JC31nQIa1j1aQpsqTd1AhQA5/u7H9Xyy5J
QDoZuu+LUZeI9lbHraCaZ5pd5F+19j866dN+arlWU8eupeRK1Sq//Os3IZnxO1KT
6lldmjd/ErZ4M4om+5OFzl0b20yM8F/LezztqvHSK7vN1k8PybG9cpa5C9JFNTwQ
eMpqOYWOXp+0/zmNnkxglJS9EfFTre7xAysTx3GLrstvVh5ias7UQyfr4PdCCdXc
5oBMJXkQowpeYhCVtQrKFTb8K+INbkMlBwYNPO5nmkeI5GyR+eIIQDBtiSdpKsSV
s5tC6pzbkqGIt/hNVb1Qre3y+PipN7hAx8xlwDX3x9fNqMfEa2wDsNpCY1FmyLJV
ED0ET2pOMGgiJREQx/MZtkngGOAYzLaW3RpemfwVazfMa3z+LWw8yAUh6L+xD02+
a8qfLYHlinExAIsM03Z/vUCZ8O0hBJPwSEnqooAu5cSDFkDeF0bkNoAxkDOgGMU8
5NaGmTGBARItk6MQ7IHwfdzUbb5/6+wxjhf2CuK1V+P1MZpvqMbr/Tq5MEXrUOT7
pgc67tDpQRUQkcdf5Lf+sdcojTzpX2coBLE4+bWuUwlFT06Xf+e9wHdSeULWIInT
XunRar1TURnmfrQfZfmgQlOBewsn/+KqccRlznRXj/x1Qs0iLxivXIwaQxkDsl7d
G0twvQuwfwo6sg5ekcAz3wm/tRAi52d6IALRzB21xL92Khsk3keaUF221NY7lsrf
Eg55BkiHGiczqkjEnhXA0ErRZWc15t3u5EPeNbXwo6fQKCDMZEbtsajBNrg7fU/p
sdXZHou7dblDVOEFgH/0kBr5sdJon1Tq1KnoHXWyUr22Cf2PLciuiUz6e5hsvGaB
LtF0lvSIkEl7gd06nwFkVDr+EL+MfRCcgfj0KogvejYgA/f8dFhrnP0eq8+9J6JC
jskz8hvFzGQeSMkll51Wf4IJrIWTNgkbDt40omiCnriEosPTWLv67z/kXIQ4QYa+
cQI8uq/wlIj00Cxalz7+5PJggHY9z63eMm9jM3pAuHNYZf28KnOBy90PqNWTKEaY
ElYfBIGAPbGaPo3iRGdBrsuihULCWggESPWhvTn6Y1Lv9zeKJ7ZfZJ3b9ZhGwrps
rB44ELptB5OyMYZ04RtWBnB6/hxNpPAZ9rPOuluokkHZGimK97pu0nbiP0vXCjWZ
iXQGJzfhrtTVnoQTlerAmBJqLDJZJsMbLBnRVXl2J/6CYvqoaeHwEwI0jlkP5COA
K/QrzLqCOTZ4YCrPZs+t72Je9vIJFV3+VfPzeuibTfSw3zMB9ldMjpffFfH77Lrb
n99NR4WKwR5KkrCr37sUI60Kz0DM129syNJrea+D5QIXm6QKfNn0k8ddKuOfU+Dz
aqEBq6zatn/AKN3a/jLEXSUXiGkJ7tgdgPVk3rMZNuP9G+6Y/Gw6+EPteExzO/3L
o1xE6z4G7ovLtXR1hLjTYqYc+QTyZtV0fErL2oGlFvfEEI4Fyn9hU/W93R41bRmy
42fXla2iRx8j3X1QL/9+5mGiAky6isUPB9HxyA8wcN5sA5b5W3627fZdDOeM1EEy
oipzITiCREfs487UZov4VZmY/4ZztCToCS+e/2A84gNEzefIzGqIjO7US16hOuwY
NlBWfn9zOo1lsbgZsdnRQtE45dmM/F8r5sAvAZOMoAJQopmQU77O97GOJfx69z/j
/NuZdOnZCMdHNGxj4ljrw7o0zUemavI8e2q4uCf3jdN7YtKaZeMc0XuBsWrhNLUA
S2bKMCvEj2jlyZW5p5A8n+YXB7L+dl+qbuBm8QCASdOG06ryKJhITyfzzjyN2AH6
LramKH5NcXIUGikY2Lrmx8LfXCpCtVyQ0yqCBZsUPnGSuA+Fp3CAKZ9HRziXMabX
BUe/FHPi/gpU2RAMvAmia5IEstUgE+Wv76NhLiCrt3u0jWxxUg7N6acKAC8+T/JQ
f2uwZLLtc/QGUR7BKhEb3Z4tCg6jsNSTcFFvqZVk9P2+QzUKORrT2P2fSzWhKvin
VZ3R+Fnj1+kGepX9dX12rRAgOkcEVGmW0FZYw1PJrJyD48mfjNC/cItP1lW+/llK
cS4JK5rEl7Jw19hY//e2wLtANmRMyJROanppi3SR9T7qYzHodgZNG8DhIe9gFNa/
k9BlX9lQm90y/QJ/JWZUGYtgNGQdBWXXpG4J84M2BM5Cf+3mhwSl9CC02jeaCwjx
NzKzv2JCP6HhTmd2a/WoK03plT2p3/Ig7PqVsB7yRqeAnKtK/dkldfQFt499WE4T
vvQWeuA2cM1xiyL58m37cY7vp9m4Jj6j7VMsv7B3gxybi51WCwlnCIEfD0JL8oZv
mM6/hgdCL6hpgpGA7ZhIcBjScMDZKcyrtJG4oaO1yeDq/2CTNIKSJe4TPeSsZM//
/cn2qE7I90QqZZTuQiCHa4IHzvyA5PhncxWr0hvF+pB95k9ZzmZddsH4LK2F6rjH
YyMgcSd6DEilsdjDvVMru5ZHuk6x6yis4JcpZjPf9e71MZChDWYUI99bJZmmFqck
nkjALW1WVNR+VcADPt+pVaLwqlHwslqSFx06wX0TVnT9vO2FI1+pNKw+KwD+TyXu
By2OLM27dIH8VVKvogpZF0bsfAuz+LmWef3Dya2MYEiuExdlaNwO2dQw62UxL8KR
tSdjHEv4xF2hRkNr+k6+wkIKS9q9t9wHH2LkfTv/gvlHwzZwWZOBYTgRIRbCtnaH
JCL7Nz5gdzMrL4ddmxSr3H2JuVJzyjdmVq2sQBVE+quFfL7Q+C2MUxSdDjhGO1K1
OVThm8jee8Qg/KGuG+ZqzmsQjdu4v/ZOqJDGtXfgIh4YKKxUSdspXANHFAuw7qmu
2UZnM2akmtzh2CCKQQLeY4Cuq6woZc7Xy1c2clz/QIFA8r7TVoC1NBHOAtyRHAmi
X4+mDMOX9zc1+2Eh3PSd/irMm3taI8gqzFZdwHkn61TgT0cpsayAWCQck6DG0BIs
dPo5tElzzh/5FS7qaIJQp7pIz5piDn+6Wn3bdQFluabs43UGQgIGTiPggK2v8asx
qJQmkCHVcBc6RmshE87z+UNhb38mD5ZCH9JblfPogcLUPunnfoTFCXzeVaEgji3r
O9BhYP27xhh6sqM24wBAlARYNrQ8GRjWEQj9PPDEM0nsejXFK5+KG8oEFyZCDneO
NNAw7ILdqcQu6sWG5U5olT3ZAoqjEGHy/3mXL20s9AbL2yMGTgwWlx0Ah/n+wL8t
ORGr2ZuFhfCcDe4FSMozpC9U79gc50v6sDvDXz4Ho/+eJ1Od9GZbgFBVR/+MXzqZ
GDzCqmwlKm5iR9e8kA+OgI3dZKWO2NPR1TtEJVzVjVXBcHpfWEc8n1w4z8zkNjXb
jLcjZ6MwJxtiZ0tOgGMsthEl6JudHYrqWaSvYsnhxyxjqPfIvUhG/7SosbYdAFro
Mj66CElCxtNyjQOr5FXNxlPNkhi22q/JuGgLm38N1V0RJ9XYzaPFoYSRPHNlTFq3
iSp9WJzq1MLDyvSec0ChudpW0qOkUpRdWHf7nHABsN1YZnFUKVAYMhLPnyixDb85
zYqmWSiiRDNFcVHp1hxyzkb/iMVqYtzIxzs1ZdnEECbc4QIyk29INnDFzw/mquna
aSFTRtw0qRg7aumnbhd3QB5MUK0EjWKLTRQ2EyVYCZ0V9kVzSuNwKKMSk0ycgsZK
WetA9FfRfUbfd0vtAdTAtpRBS8qKSWfJPfmm9BwUN7EazFtC7KQG+9XXp/l7kXl6
2f2+Gljoy10vSm4rfAYrTyj/H5Z/5Ry8wcKObBTj2QfiPiIKCdy7Emt5YYXpMYg1
liuA7PUaGd82YJNXNw6WVvXRPv5Ujk07/tht2u2agx5oZ5uI/6W66/F/o6GlAfl0
bLhBnyGSo4lMDhShciu88s9m8IdpruQXyVtD/Nl9eYAvDZSVBMsQl/xQiMUMdssP
qAxO4tS/1Y0j7vXrmUyKCphnPA6lvMPe0py5+yA81W7RUt4e8bxvS0D2OrlEc/kM
sVJ2b8gVHZfe4nt7SiLJG5JTkSrIVBFhTLhV2uCG3g5OIPW2FyVsZypJDvVFWluk
gdnhDPmXMqruPg+MHFfoSZmnkMK2shtLqHRwnkEsGZ0XB5zF6C7E+HcyIhXlbDpr
OOqQ9QaeUxVOY9ej3aLIx/hiEwKRqKpG/hdHxaqqdHSTUBSc9RILw92QQg7mSaos
1SeRJWnj5YuCPmx5WbVpRbS8SfBtTnYumypRevvGoasZ7bmalExhWPOrL8wPE/+F
Mc2s1wVbB9WUhOvI77YA9khvLsv+YMjzlz6mu/S+2PSjRZj3KM6/kZ+gUu3gKiAx
FJtKVNGJBkAebQ9vwkaOFE8nwljsN48boLnLQPCP/rwsAWO2v3X3RkdTFF+mRFy1
/rMyytpSHoah16oeYc6kYb5/o4UuvfWhENCJu/UgeADMtAjj8e6+sbksuqROlxwQ
Zo+IeqeLzP5KgIczteRktoE39JZVhmgh1es91xZZoDhVBV+f8kP/ldaV71YuCUhd
Bhzel6ezgeDkXtsEbR7aVso9PnZXM3hvQrHtRJHVLizlSchk8SCAgFIoxtoEu5p/
40Ps9+LGpZyCfAkWKoY+N8i+JJrapTQKaHPLPFBD30vwAtckmnWiQl8OZHNvMURr
x6ozb4HCstlBx9w7B3F6/phfZpHep6ZxCySVMLHcgzEBffsarwSvcxhk9JYGVudn
BOu/jJlJHB2gPbzvQ77POIZy8HBt/m+jsBpifPC4wyCOiXq9WX7CS1KvttKmuXaF
dx/wK0BibLU9WTtTmMM7rWl5ERkqbc1zYyPgnEec5N0KvPanMGwa8sfeaI/A1wTm
rzkRvbJ2oXm7vMj1ry/QIxxACuuvteel/VNTdzArbPeDtH4FRIyKkOSQRs68f0bG
jni3LkvkkJ767c3kzzvuGNytCNpVR2zZPgiUyXYmjx1AQmr+qJgByDMOx1cyybdA
QYiNE5HMqhgiaD+6/5IeDA1/2rfmxikvB6Z3sPGHaYEl133S0P9CwOv2zr4pLb7t
QcIf3/3NHfh8/hR8PRcDk24bnzK6UVyH02LcZ2RoDpPdCU3ihFAehOWepZ7Zcxqj
v4knF3RC1DCVFq4oFVdCMtl+UEGVItPXu4atUNYaJUhdgqlzWhjR2sw9Xj9fX4Wu
u4pR5IpEOISVgGSA+eC7FWoJIHm7MF5N/B4CPa+cY19o6DSkL+iz9O8RHqGc63U3
vUZz1PpWuiogAGEkWNPWDl3eKagKExPEeCvwcin5HXdHpoTktcTQOCo3D/8018ac
Jw5ZwiQwNjLWrnW9vygzCHtAe0p68KtueMpWo7uOvfLs7Fs+N98bwwYYw6z3cpVv
O77JvW/iyhAOOUzVfUWQfoe3Fn0zJgBEr1I2wRXc+Facflzb/z7H2sPwIyj1mjW7
z0ONEVD7faCRY6k3NqyZdpgJxcJgwIRX5XDEfExZO04JpsBFMQ8s1V4r1QF8t66J
E68xKtepG/LwkJ6DNSBwvYnpJWUgWwNPz6rqudYIhZiaDHqu8mRnaN6NBfuBAAYf
Jt+S5IBAGjzSzDuaSYpZ09i9cA9zQct38OXaWH4RDVBQ1yTqJL5Svxz6py5h4zxf
BpmFmYFajdP/R+O/RyddvvHbm8dOis0MSI0+AlWci98Qhl2e5zMadTgY3XW9p5vv
TOmtkEMRFhRxs8KnUccUew5or2b8kAFiPSgjSYC7DLOOPBp7g5rjj4CuqHijO6eJ
xy8NGOOymWfOQ7td9A+HApwOswbVVv5JytWyKj/q0QoK+Tp015wtOYakAoiNM6zT
nLJvCzzmwl1riYXbvsz2jL6ASLHK2QTcKxmc2eKPqZvZAlsLrHa02d6jDxO+427b
Zh43LBq9b8DbfB9r8wt/mvRlFVnce3DmcZ2L3ZAMehdi64TVESRh4pyrbhjFInUM
08QrdSfjfa9NPlwtPNNP3LvCMit8Y2L8y+6QULDDaV7qdNd4dmJcWuN0FXAyKCdM
8qMoP1W40a1lmCJpMiwJ5NhX49t75Hfsg8O0BHTvRxRYK90ZQnsW/PqlYcefykD+
em1TQ6KlkDwFAGeH8a+I10V+nqbv7RLEPIMF2Lq7p/7atEE0BxQmHAe564LkncgA
uwD7hJ1zymY6fRfy9HEpN5dWCO69Bittb6El+x+vjQOJywynGHDnUirfcU1Bi+Ki
IMcFDFGK6V74gaM7hs7DrfAqlKvMxWwgyBSqg9ooDlvxrhRDpFCNGB8H3n391GVN
siMR4mU4yfcTgd9E/3ALQviEaVBfQpD8+uVKw6OsqKwSvuYybtIEW4sfWkE6u8pr
EUkL7wKifA8d8wHlU40xSHijjshFRAXVMPC994QveWiWLV8EO/ObOUf1yv3ymeV8
U9Fy6IgseggmuTjKOuqSFwzGZjBs31K2N8fPMnVw86pbKV8k5TmAWviVkgxWYyYa
djSVJVlp+k7xGVj9/gMNB/7qT/W79PhgLro8PSVTaM4SnZDBnHZVeqtUzm5SbOww
SjTimTjJjUA6I6Mpcl2xhPd8ME2Wlc7PhMJS/K+bWz2zVi9prLECbDiMwt9yh8pd
p7PPGEJeiopxxj6RZCNnFIMaNjddBSsvD+YWVdW6nyCbY+dbOA038q7pCtHwCRMB
ZNSLzhjaXq3lwYZNMyI6JKxTIluP0vhAJV1U+NaWLlG/yBYopGYdIm8alj196eni
fNJk88+dqqdPjU9q0q3LDhCipujSAbXwo4bMp+7gqkaxxphrVeRCXdk9MofZk38m
xWywWO9WOUbn0xsc3y3NX0qTWHX5MvfhhYif5Z5d2z2QY7YkzKMGRUTOcqy8lzCu
KYsLf/SFEFKKegIxLqUJbEct/H3Ahp9TG9oogYvXjmVPf8Lh1n2JtpL1WG5jyQSX
mTevIlLxD5BfiWdVmCUzX9j9SP4p7fgZaezrH+sVbS7NcOv5M5O+zn7sG8cRjkbO
ScOHTIRHzhJZEz2J9NCmoFjUWZ8t14N4VXe75LXPWiSMzySK7lvEipKUgfPUeF06
xWrEsg4hErsHlfFI8/Tx4peFHkV66cF+DvEFKqQSMXfdx2a39uXt9LovbYjpiqLa
oKA71NytXASXd/qxPqPNBFN/K2I+h2bvL2vrj7LVzMNVnfdBxfG0n3XVeBqhzMHB
u4uSbnD5UjiUAWBDBG3X6Bv3MXPa1IUzwWG/SFXHBvTLAmTtot0iictamhcbSWnF
PmxTXQEe3nJ5TTwyXTbf78P6bqZm/B5Kv0LxUeo5MJUcmzXX9AxxU25n7U2G/2Ss
dxadf2TM1I67yprn3xgreXhbfdm890oiLM5K9aS4f5/WdpF97KPNpw6T61I9uJXD
0ktMtehe5MVu/JsCxCSUPnYE9i9diyORYejA2AgPW0yeithKmy9so66TqDKDkknE
y4gE4KdaZT5aaURypH+16dRBWeRkuA6wBS4x6kPy2KT+0m/oTpTsFgFTkn7WKwMP
gBTrDhXjTuuGV6Cuy2XGzO4p5bZ1ZWZwFt+7bOFtVBg9HrLUqn4JGxuPCMI6Jknn
/9PbkCoXBBBZr0yoWGrJGCH2vqQebACenJMFiS0jCvUxgQN/H2vIB7l0QtddT8sq
bqz5VTGBctLv3jSFrH4kELOBqL8SrRRVgCPA27QXr+Bb0HEcQalIW/xwDhE15k3q
UjqsGPMI1PTe/Ljb/Jj9pkOQl7acXR+5Hk+iaJKUFh6aXU7RmSP0gbvLyJcD4SDL
ylML7eEz2ozbLxYPNE/FfPB4TNebJWOZLGS/Tmzt127sfTg1fHGn3WamzcqOIqnX
EQGb72xV/RyVaVvhbIrI+EKVVRnr/Dh3ra1FMuWhrUspmex3f6x9pUTS1+ousBgr
Hds71WbM1ijh3dPRTyaKpH8Ud8HmUTioQQ3TRDuKMLrOohXwoOmf9wsa0TpUPuss
tbiT4Y1nx0+AiNj/K+vT8j14caRuVPb+d7SR6mK3k+fJf8ieSW6AiIqDl6QqUvXr
zIUKQpV+2oONAtfLGaA3hi8iXJX/cTu9o3351h+B5Mc8vu2JxqTWac8ZGZ8uY0fZ
5QDgStFYZqmG+pOO2JOm466vcX8Q4edIyVxON6ncR/oeg1SRGYijYwgF6J18dQQK
7CZ0R/qbRxuRNM/BgNk8lbRFfJnNkg6MtqZ0tty6If3SPSwrUsgsymaGgjS+sQM7
7YmSTrSAIl3eRVtn6csDdwssbyqLywdtOn5myXkzDmJb06wgYPkMxLQjtICH7a5a
E3q32gwsQgQu33Ip10q0Z7bbNkFrFEjQfcmPz08zuFJrrGADYuus7KOpNGqt/M+N
g3fOoJozbQebvheqnKkkUlfVZExLlAGfCeTVdiLf66/2C+ERS7mfmmXQ1Ds8TMHF
Q8hwWu98kbAFmMooIGGt8Yx/3qmhGTpNvmrZJ2edv+lj+25DNLNiCJGHIwvk46w3
mO4vLnUt9LhkiuBR0n17SckffRB9ALmrb5W2/KuupLDUQI/IaoTp41VBNIRfkoAB
I8fRSwn94BE8ETh4XdiWM0QvnY1XoS12KxGVgMmgsXNmJ3vVx9cr7Sqby41RfBzb
O39vTZk5bhVyjFBNO68Wgb0QQz8HbuP+NOuTBki/JSWDyd5OCUIGuLrJzeeCDSPb
CHJPhGN718xbZHySBwviAPWjYh1TxXv+6KZwDN9pCYcbvB3Iwk49evfrryPUDoXS
mIGROoM0+3duvlU/AzfXLRFZWFu70/qjlm651SXFFbMS0BkekltPyO2cuOnTSJX1
vCoZjmBUXgPKuTC14fCBB0JRYl7wv23ymsvozFzVqgB98Gifu56uLEhmfDoqamvp
jTMbJ7C/K/+qYgoMnVQxqSQzlT+vxpEMpE30ozaQHrd4IOS6NsT1PT6ZS+B82h6R
J/bVdgPIFkZRswWU6bUJJMdG1XaGbVyDHIeq6ZT/mn3GqQVX6wB9ULE1Z/UDoSlt
u2o1F1QPULVt6yoOLqg4a5HOffTsGSmPdNwSKnEOTFWN2PiVl4Q07P5kJZ2BZ/1G
8OvRmunUuUeYu3CypQcmqvl9+25x8/t2BWvvpSfUNWTvfY+O7XvqmGyNaBRSdAOF
KrS7usoy4k0tp94qCFtAcxYKP8HGF7JN+Euq6/mKd7sOUUMPE/ReGW2rgSUdKJwa
DVN4liT9XvnHJt6Bqc9J4gSxFXxVAscHdY648b73veiab3jrybvZCfrPc1VGIqlV
gjvkJJImAJ03hPfQuNfFpNxBIBKIjsSfiTUohAiZ9jyPxsLl4p4hQwiVYQruu1zW
JXf4WzY49aagBYsfYi6j2ezfmzSicrm2Gn+5SGbe2APoORCFs/E6wbWOyD0O8mvt
R3uy8znQ75pvXVdHR+G/u/rrPHy4sVd6hK/dwsoXjWijgTH7WfuhtrNwqx+Ogaap
+b1AtrHAb5tbIABSPQeuOD6eHwqTtQNrNQVuUw/JR+wK3qmsBAspDQWYDsK5vtDv
DPKWtsS9KMqCCEopyAC6hTObgi+sov8hJcQBf6EotDg1zcntgiw5GLML05UNz53s
xbaaZaHIlvxC93HM/aLW7aEo8calZqh5i6Fh/6sf7RtXpeDGbA4obGa64cWaDUaY
cyeuMDId4w+7thEMx6+ZOn7XtaIgjHQUqxctiZsVrZfFhavSd76Rk1Lvt6fr1rZ2
+Jv72xJi0c4/W2ChNArzw1iFX7Z2q+d4tx7PvjyxXg4tkXJ8OrgLXfcnp8PrSqVQ
w2scIxdluve4u5oSeg2CDC6+h+aEvHYacj5ry+5Fr1XE3t7GnKkLR1JO3a1gQF4H
wiJ+v7osgfxvzuHmzsgB/j66CgT/NAhwBRInOxuRMKBabYfdcZN6ZnboLn/1a+1I
WWJ8vr2QT0/+SjuokLXglsVwK5FKCLBc6tXMBLB/tcxOQiiPpK5rEBtf4/IMeo0v
HDCaGvtwTecDqiiOIVrR2t7nIP0Jeg0/9QNCHxHTc5Oq0OgG9v8f1ddj+6PCK86z
pxVnTcT5AzYLu6ep4uezEUtUpQzRZ/0IM1qhdoCcb8dtOs2FHtxs5gfZFfpXqCvP
74OjR9aYLOosBFHTRzwbv5zKmRZj8VZcXa6WK0v5swSs4+4+RaumDrRWZDnrBa6p
M0BSecn5cpWZ1bbNPXBg9USLGxnHO9jlldZHhkEOYe+i2ME7E8DVT48O7ccweHvB
vSbztbXGHnEEnZ5kwH5rvonzsWfO6YAMV5DpM0bok3/v0VyulAPG9hGfmLgGFDvF
To03a0A6UWe9Ln9sdwukohMT5VL31cbZBs1jotevKRxE88+SoYF/8beHzBeuReAQ
zTsqwYWLN8A++OpGDBGqMsLn3psq3NMew9sDRk0LIeiHfyFKeEZKokYo4RNWcJR5
ZoleLqt4Mbq2I0tP6Sl00vX6SOfuvXt4+eA2B7zwEjCTUI1qyszuODawDeaQPQ14
9Oxnuql2VRF5rMHu/dlyEKN+KlL2j1T1ifw24CTmiqiMCwAGL9TTznvtX1KB8gW+
8ejGvPFmN+FUT6nTNzqBbeGEKP72P2NVm/x5qhVkWo51Da2JHrlT4/Fi3WLNRi+o
aOkSooGfnnbUbju9a18oq9atnNWyiuEOs+yN7QicRJ9zuGf53297iGcpa+jUhAmY
L4W8ISjtXYDr4LXTlmQpNhK0kwTeKYwjMwlU5dzIpC10fX/Nqxd6FxU2b7cUqgBc
9cKM4SYERrZUNIrUq5JH15zndc+pBEcsXx41a4sDUfyThGhNgUO2oQgyKET+L84+
l3zvYEnI3ma2627CSLvShV1ViYb7HygjFTICCkxRp6jh5kmhqBxdKIdgglvCu4v6
uOf0RXx4aMSqoOmOAoeCJPJckYV30/TF1xYg7tLLhGzqiiJoemQYlOp0tzphdpsH
oqoyO+tnfNto6ZokdTPp5TjOXlZrbhyJg/qBdilNbYwnSkqwkhnoo8s7XRC7QpKk
LYHs4iEZszWtUMCoU14dVkz0z83EZwEzN7NnKWgFAbCLDZbdd6y70bRrteLnGaN5
d7QJSEkPIFftalgGf7jHw2kyNgXRu8Ht5GERKIaH/MO4LYvzp/Tw6FlUgX3dS1pi
3RLMO0Lzs/UXTsBVhcAPPiVDmQ8i4kLDeOWJNF7/3adzepiuNigYxMT2xU600DLd
ovyg/5Ie+kWum1GqRBYz6y/r3MfvTh4X4AsjzcVSIhTEWFtC9cj8IF7t6As4aROG
p89MiPfIgwMepO6y0dkheD8HvwyHEX2rb/LqwEcQYpP3p0Qt8GhKqwGSTqu+1Hbr
UDY6UVgXcuXILsemPozbZewd2e2SdFhF+wUgFRKJr6m0m4CGuBlzwMWU7d5h6Frz
GLKrHtFcXPUlHXIg/ohIpx3g8Sjl1KBWv0GamCPWCW89S/9Zld8BY8kToOMEdwNv
+9o9S4a71vU9mOBL36czhFIvTr6GfuworIiPas/zigyOvlVxHALZXoSknHGt+HTR
00/3z+pN6fiIiFQughjzlZYc12+GLix1OgYXp0gng333MGRjaypNH8BjQ9+RlNbG
ZtQTOhfTSsfOom5K/1eq1anlSacu9RQhuFy3NK6J/qoSJwFR9WMjTaqXyWXzSIDX
dqbOGLz466N55dPzluwK6M+jn//qyA9hXLLtOEKzao7fGPfPH4EAnofiNNCFK/XF
xbq85UQwNDajAJpvItslXjxgjhXYB0n0hQMfgSczMGopRjhsJOJBx4/wWal2oYaL
FwcrU1b1Mt4BxfP+yxngqDZjlDuXPFkBKlyrG7AmdloCDAPh2sLXoddgMnYvHEvb
1+Le5KCalIRQL9nbcRuOduEfatSr362JJAZCm+0U4roPdcxK+CnWsGdfic30NQ6L
H3Owd64+ZTO3uW+dTDdeLpd/RGsskieIobioWGNi+gbXWo2kM2PeIjypEW5dZvfV
Vn8TJm8V4bjilf5e+ygrJg14iP9qLNvopbyiE7/vxxcPLCxY86JiAaWIPX0OR+iq
d/YaP5jp9hd9l9LiuH1s6tS5vnk4sLdBbM+NzoI9xVeVoMm8EsjIdcYyzFtlBQHX
fJ7hkFdqhZ4gYSErNAQWrCT8BQsNpOmyQ9o8j6JmxgN8rQDApykuVVzgqW9cej5b
s03JbaGk9rXOcbnm+uwDGiQ6iqxJUci9mSu/7Id0fz8mrHjSuR6cnN0yb/NlDf/L
1cB0Ovs2MXB8xqkS2wvimAjW7QWrBs+LSMi8UDiuZwXGyZ4+7W69gvD8wvTmdd/m
ig3iz79f+K1/F6Ggx0NHCORKgOKdqX6sD0p+3mKxChlW/KQuPYVFj5l4NYtrVgHQ
3bgNEbr8B3TEt5gc9oUA1O8PiarwuuVZ3/yWzNS+CZWiAIcbXzpl4z4DP35FsRx1
q52HqC2ACJQmmP6dxnP3upC3iomzdmfVuwc5Db2BLAOmd7Z0Emi0pcNqJr8pNZZF
O07Lgbdx5OYIL3OKpA6wIpYVyqas9wrcOzqxGZKU6m8O5xGHVr00VIv/hGYqn9TV
A5Qq7C2xMxljp808WWBQo8xZkSeBmvtmKOM/VLERGsRHqMfE/VCQKIDZcM8+qyOV
qWPiLJ2QX1rWUtBQ/cBL2N1r4trth4i4izvbiyUAG3VvCCLgsqwuQcDcNDTmtRG/
RKktkspcV/NqOuNZWMQAJPsN8EzkJIrZGa8cyusdg+uxL+1dRWsPi+XwjcMMKm1P
IKODzhmNYz0SVr3gv2LbSbGgSeymuwb22MZ7PjJys9NPZ7QSDREdk2dt8vkw+nDi
cAzF246YBCKx7U+D2sgS8lxQm+cbUC97bsf8X78Gpz9BzFw6xsaGVTWKdK8BR+m5
fjgoimN14XZ8BWrkRtoBMlmHxohLAmmgOsmiXiBph8xMA+Hf2wes+vhhncFh9VP3
o2OVFOy4xkCXjx8ky2huvFH9Nv+NcoSAYd+pU4YRafDHSvnvXkFFRBykssoBueyj
QGDJETgzf+qsA39QdtdymkaDBiEd5RYGdj11I/7Hyiu4D7qvz+ylLnyaveP2Qmke
lGcQypjLNwAe/ifONLqWx3JrNqC530hn0/MNXCGtGOx0l5sI4v5r7/D6++uracVG
71mmod7HBDZOyXS4Z0FKPhnJjgy587xjPnaaXq7dl20ulCj+Ni/eh7FQvQkhnrY2
ER8c6qofIHRKSZ7/qTdrzikZDVjNOGYzODVk289Vzat8c9MPwOj7njXAiaN4gOl8
5GJA1VB6IjSGtQDofMi7a+zSIkt6jgwIIma2WyIHHxgnWn0A88vAx5FA4srEYVDt
BTD340s1d+bFOEyscP8j3n7pmigfFQy0OG4APAAHU4was5Vcg8LCV+Wido2CpDCs
pBOhaT4LRctktfpxDYRvx+mTOlpMynMtXLroXA0mDJPPWUm9uqaPHymwZruphT20
sAVpIycjas55fwU8v1Jr7RZBY9ZhuBwPZnuwPuFosCZRDBMirz/M5ceHcRXqk0LQ
FYSc6DGf9OH+MYV88QVWdDS2h27X9RLHlDlAylraFPVwOf1eBaHbCEprqZlJPOxz
oBateqzzSZVkirrPwcDDsrc4o++eMHx6TUUOIyqUnVFHNsLf+bv0Udqtkxc58Xoj
trrXqWyrX5puWluplgTNXjZCNky8TndLmmDauTr22k7QV2b/ANOpz5q1/I1/8vvN
N1+7ynwcE2TkoJ9A6gbaFv0PHy97X1bRbpski5Zb4IfJ1nsqKzWmeDBPS+Rr4b+K
A2Jdz31+itWPVBOO94YdPHUiPeRwK1MdnbscAbaDa6/zyxRWbTuZB52e2S7JA7IJ
ZE8yhFrzdT8V6sxID5kazymnWJdpOPaIi6fjysJlk4/l1cbabnJGFyI8hH7ubxKc
55lbG1UxX/WnR3/tHz1L8l4dmPWOIiq1c2psb2/2JkweJaa2q6M7zSKq2i2jX15b
8IYVL6A9XLNDAGmMicj9NW1iEOoag0vF9omrSL0Ytzloqu0RAeOQ8OzwP4ju/Rhi
XUMm4ncNwnWWAEoqkea+8oU0UBzwZZ5SquBCJAwA7p0jznMbdXhQ++BdVc4uL/V2
5QVKPAHjmR+SUw95JF8VTmqMoQ7b3F8IbTuAboYs9ydgMaFJEahhX168zr3FCf5S
pz1LntuMqi2ilL4+ndMK96rTOr/CuHvTepnSHyo5P5TdP+rrb/KKcAcKv6ORkIBD
d/zQ70EovUWw3gRwo76EfOAIC6EGeBn0Pn5wxiSMUEeTP/TkH3aOd+YWiHl3utSW
GUxkxgLwfdOTwSwBfhjqLNBDtC7sC4rDcne4HMXcpia7v4aFcXeLYg52uTWYGLwq
jY3cgvz/pBNZtVU2Mi8+Z2OK+GzhsHXF7ZdXMPw9R/anEmI9IkZtSHsNmzf+DJct
RYRBzf2VrkOd2PJ7TNDOu3nHLAK8EAmUxQp02EQZK3scXE+nlqzAgx1kXvLGWCET
uBI8u3nphHo4w7oYQjcWD1wmFO2+oISTih/jGePG/jNQGoyAsqRSgLpnahc/063p
QjKRgfOtZTN8GuJg/mzsjkITg/ZTaItOrML3KiL4tcra+Pc9Ndis1tbdiDqrZPe/
+cnUOuQm2kxPtOX2cTPdI0GXMJylAjuwYKqnlAOjTgC7trg5FvgsDLq6adRT+3iP
47T3CyeAgKAPceZ0ikHKJuVipqGgXYyA/22bVrnt+Ab2KlMbTtdf54FxI2xYygLw
3K/rXiWyFxcpQWudqkieLYS+Qr1dUWsLPfqB9E0bosOU4iUr9Uj73VQ8Y1zc57Dw
tPjDl9Dp3YBBcbecKhEQteqxZgdfENV3cYHVnddCLiy6zg1bj8A3l9Fk+paWKAd2
JxYZzsYfI2lG1fIiXtcC1YWmtvhogEZtNt7AOMNRj7LxQ9EKzOUc1D9bt/w6PQv7
kNmrE3GRlsZGTccoAK+dUR40rtjJ5jH8TOwXF4BaYkbmm4tYkEAgg9gptzuC5AiY
jB1Me31tieBt9nz6MOS8aZS1f25BEMLiF0191DtRtUYFaRjWNkKGAxWZ/Q4Uig7t
iy6zQdzJFt2e2mf/o05tv0wH78guBFrZOR7uTkeUVYRoXZb5H3WnOEYGLkmKXwWJ
tULZv+JvO5ZZ8Talzb2QCKBOhdZOQT5JpBxop2alSc9PdFrlhsf16Z46EZZrAglb
RKHJrUVnLzrJh7qFJI6c6+G1GPoowsfYLA5cZNSIVY0P+5k9Y/OcsAkugaUuxA3I
pCCjgu+nVjK0cEYdsLtnCwVrYhlPBTmEfvLESthYTuokBQ2U8FmIkWUrCAPFVxY1
nB4kOUNwhO9i9B7P0t4cmht/LMb4g1u2inkCUpnjIDegQ9s0ZX0egHxujeJzI6Ro
jKnOYL+tys8ACpIUN9RBLu6DxBPdREEVbECwmsooBOoNKZyWuJTs3tLRX34Ce4Ln
dfeoJcdeitxOa2eJoQfM9XaJDg6gmFTWbk5TZSHOxPDRn7wVs8MfZ39FQbDoR2OA
CRzz67i/nol5VtZb4aRrHkbnYZKh+kn6kOAI63DxKyILM0KtLeU4c5WqlfjhDCaY
9QKgQBfLX/n4n2jsAyoJjNlvnWnEpkDh1QrZkHSpJxnbtMJXfuj+eIWF/BIVmwKN
8paSvebXnxvtdItaazgLexFROPbDFZx7hLGPNMasBYCA1oxUqec4z+i4SOwXjlZn
llpbpqjHK4Ep1fZJgq6wF0s3IbO/mvRloc4ty6U8sY24d0jCXx4Cr3csILlzRWbL
DvJ37VcdPtwRhZR/Ub3cWfuddKXZwkyUgbxvOxXxuIQ8JKnJKo40uQ+PFq6608Bd
VnJk7/xZhDceN1ciAbdwHyUcKTa/7XLc+/tDx5YU/OLk6V+81NrPfIHUhpnRWtAi
Twznmh256ACV2tBZngXsugjRuWXEuP6WqphSoijdH+cR7+v/DsiptQ/2n19d8kUy
09XoXekjCMhVp8ijtZHFDGUnQKjhZnhSH9FngEktUlTRJQ/iMY1o7uoOuVVct0O4
1mlidgKnlqqzb3tvq3EgyDwOU5kLuPoC6+NMXUSFUc7zZ1ubAE5KAKxY6cysJZyC
wwrvyN0BsL49Q3Fisoaj+Xs089cVuAt4kKfDIzTTnawGeto5pMDke18TauY3MMcI
lZv1snuwzbhNyqVDvY71d+cvXQnevthfGaLV7SU1xsvZ/g9CEzpVC03FXy5viWxP
4ysq2HvLze5ldG2VmVZXSCRpuhiAhheYWh9PYvuCZ3CMbV6J9gxll4VEcs+Uj5f+
TMbHKqDM80C9vj5fR0d6NYbARzGnvPW7grwM5J5+ptfIazR5Ysg989aIO/iNd3kS
LBapcUrxnTaXOhidV2LM/IeqGHCwqs346rqFt5dT0PnJXIHh2cixw7v2azEiUS+e
prB8QR2fGU0HylJR8kwmYESZIpB8HIQKNnlAyA8RPMyUUP6LBa4EAGJc4AfaSkc0
z4g81qouL0dpMhhLhDsV84YkgJipfiLiv6hbqjODj4cShDhvkRpYYaRfEeItaJyi
MZxU1K5R1g8M57DOgA3x6GerusUCHO/DcenGy16/CnydI+Y6M68zwjdBMWEZ7QK6
Vx6KZzrstFzth5Oc6GJXCXDILOHjKwoQlF1C5nLJBdGLZQqlMRXQGFhdFpjSD2Ai
H+WynJ60ey7dW7SqC+4JqaGK9i3obprOJHuu/7boSfjXqtfsWa8NXZUwuh78Oy2s
fRAYunDriccn0KMEsTo4L0HKHQZchbc+4kPODUBqscjlU+SR3+91BiBUZ4Nw/GHj
JovMhy0r1RYTYczgKZKAd70mGg9sW6Gj7h+cYlCmpOoMpzrf3mUptRgYDcpDNnMM
Vf79M54rGTfQJi45R0KGAXPX+3xoVfF/019zf9qQQnXY99Cm3avjjpfVpB5iTR+K
d97+wbZS/XdwvhAYuGU3pgEnIjE4WL9hfClTfpggypdduHigICyZg/Rhk9jdKhcp
4YlrBHrvZYmmuJV1YVQ9T3w+GEKlnGA7X/6ghWe7jhBfgneCla8SVjo3ucKEOX9s
Hwd2W1IdOxYBqJ/lOkLXzltwQW0vRxLo2h3+H1cUXrWXmz1b+kxGPX1o+5GZZ4E6
/Nians6qgwkibzxe/CxKQqChboWHGcoA4b2lmXaNXSr5Gky2TWvm+CqrvZSV+5K+
LWLduyxj8PlXYh1PnP3H/3AbtvXSvLui4cXOSYiwuptNcWafGLfB9H6au5CM/+PQ
883ZtdQw/Uq2GSRoA1KP+hAzi2WT6qyqXI99xAywkpFrBXmTTAXaZ4865HPm3NlL
Yc1AkHXIIhc/O/PTtrjVmTksE7/MnihjklQgcj3eVmFUJ/0YXV2M1UFoBZ3maqln
RM/WBHFQYliIA+F3MO/pZJuVes/mRvCHEZHe4qw1yqzJ04OL8nldIt+sM4Nx5dhW
pcUGqac4QQ/7fhB2JzHV5LfVyp/kHinFb1676JIglb+bu/WcuujES+J/1jtMEt6h
DqZOp+hps3HzootXbweDiCttRjlGSdM3GtgvOo0ePOpEJgY2yg/GaxIAPWbJPZLB
RNN9rkZsJBJuds8ib/D5JXhz6pAu4Dj9LPqKX3wBi4V61RpQeIDcrQRklyI+dsw0
tlSmGOR1TlmliHPBefDfi9Ir2EC6pBq6cv2uZPbbPMZcx5/AglrzRb5pJsIjug7f
gDM312QvSLRNh2Lh+VgONgpUyT7c2KZRNePzcTL7T95rYmIF4R8AGfxsPGgB6aY0
Q+4fztJjTtKGNA79BP9dYK56LPb0S6scu9oXKUDMxixvzyX7nDGQJMRNIYpoyNI1
ORVZnObA4OQAQwfpGVQlyJ2AhNR8EPP1dYsaW5uExGLlITY5OiMtyieqK3GUwatL
lNXekpQDeztGPxuweZ7YGURbUky3gRFVvqy0BejycBBBbjmMLyUz7qwOSUqD+PUN
Po2GKwJGzktOzc59PK2baOmsFVlp7fQQhPal/tSr8YraS3kB4nTPNuCgGkq3u2Gj
gfKK/p4+dBrBPTlJlKN4+BRGAiCloUW2WDdmhI/cWJHFCwI8P2mXKKc+GYbKsboC
WVHxX3YId9JEVxyO7jshFzDmvBfWkIEcP/OKOKrmu6fU3TB6/2Bfh4bFExfzWnBs
csiaDeAt6y2BbGR/uWVn0l/P78HdAD0yvN8vhh52c+fSrERUNDwXqmxYpNmWM43V
Rqc7CahSw+jiSn3S1OnG1dMz79O1CqwhGcie3hNBxeWxZXZguNGlD5HMw89Kda/N
NOq7KBqfD3lsaEv7F1AF8jyUXtZR8Q+l+5zGZTQLK5gah2xay6kqFBZkvoNP+WCF
LTUXfo2dOP3rEOHxaeV8VcVbnPnSae4M6f11kThIA1QvfAwMBZeSPzqBmLY/CznB
8JkiQzghsiTikcd1qmMZGaYtp/eA4aqcuGIm8pWzhyNUODokBwh+YBaQkhGCt0+x
RMmjKiK8iGhgx4Ytpqq0CGRmPUnBCvNfQAW4DZn3nRipT1dLXhdCPX+iSZ3mKD2U
l92l8mJGlmAEIMfJUmxkTghDF3cFtj7ahH7KfDmKFEa0VJZ5YcUKhppoeZzYQ2cU
Zv5J2XIgvAr6TEfJV2gRgWGh9lP5iGA3gu1hRCj3ilpN4bwddyl0vQNp9/xuhKgE
8Pzf8vi/JANH9Lfc1/mVmOHNE+0QxX/+RWnKC3+I11JV4B83VyMcE+pVasdXOU6M
fA3KIryZ9jGhDUQ4EBYCBGFrI9fdBB3UBj8XZc4vdfhyJhCzmsOmOa27F2A1mFh9
LZzksR8OYXacU/xIwwG0ah1+QLNbDOexhtRkNlrvqUzeJ5/BbKZQexC6VqwD2X4G
s2y8fy9dy82zPDhZLClQALsQKaLn11HZpTFO4EbwYK9m64Z17LwKFj3/F1Di3nHU
MMnglCqdNxxxu+V8RAyIfkzQd3QVdSW+ebWXE0SjRY6yIMbfzR16+mTK3JiROdik
V9WxzW3QX3CXEHlaBb26v2kicNfJnUevWAlEG0FdHrx4LZLf5NYlN5KdiZXr8aZ9
IQt1bNwEOyY3YcYqzIY/y4sN22qAG0Vck33cE85kNUBfg5ZtBTpSskiCYRTKRr6j
OyTOgZYGkZuMJNMnQR42GgXftp6Y7rkapxEvGNbFoxBPRpEk2DmumBeIEh4vhl/B
/bdnXrApwsWlxB361zyHhyo3rsQ1cvIyMdkb5jDQoeg9JP44BHkH2LC0A4t5Y6FJ
LUjzTnq2iIqf8rXcRyteevBXjEVlRS6xuBCctXXrlVeEPmxTCOMlU5H8tQC2ROni
nMyGg9dqaGpjOOMqNyh1ZOpYn/F69DZ0l5Eq1VUQXmWpI3jZyyVuDBMhjIxAOWB7
DhZejb+JIa9xZjsdLTL5btnDqKEye4y4anZV8tfqa2MSADZn4pRkyCJedR5upUTK
9wv/GE+oRih+hXBSUm+VozVbdYYSk9rNgvDwvKOLwCdy568SxUASKpBEZ/0sj/Ef
F8CUeJldkwRlnLHAVB6u8z6+ATrg9I50pVoE6yolQQV6+s67zxNXV6L6PXpciGth
Ymq8C9sabWaNCMHhIubaVI9oVf7x42GAF65CtNPQ5eJ9Vq8iX1AuKH1DQG1obSNO
Mc5P+IqsZXpVn5punLfr4Pyz4AegUolUqEFeNppezxll+/2kMs/fOn+UPs6gwaCh
RdVgtAN9TcwDqjjp3LkeT6t3qlwpHDtbJWpcCqApcmkOCeLL6s/PYHCVw+qG5YJs
9dvBE0JmPBsunnoBuH5L5vBAH0mZ8cIeDCu0QOuho4ISBpHf3YUicJ1TsoXhJmAU
py/4gzfnBFX64AhDXA2pEJOJsBR/hhI9ikmuA7BEm+tkRHyHtwmCFGWfxV96+dSz
+y4dQA4anMc8CoqoIq8XW8QBaSwokFksvB9fL8CA6iRDJeLmrJynna5svHTULucP
S1j9EeKPaewbTquYbMBhD7wlAxlc2fKMLDQcfm/Fgp7tFowokTt1OXITS1O4ADng
v9VdMDhziG5MwnOHWstRRfJOHyL0VjVrFz8+nxFenzhEWLivPGY2umpPImv/VbWO
gFshDRJGWIayqv6JgfQD1cVzRh2zex5Xh/kr7B4baBfkn/7sY0FUShbv5WGXU6xj
1oInJJ11CByfpEU2nChKSPflUl4bOcSgmwpdIucGhzXEUhpz1TPl/kBUyizKMwDs
I9fWwS3dwZc4FskiriHTHnSFsQI6h6hG1WFbSWOKYXaTIZuMVlan3PKEXSP6ICQD
3Wa7tuCGo0+g4B/w6Bw6khgTtEB6KHP8d6xHHCB9Zeo6BSBZ1ckBn9P8TAMvZZaT
V0J1VS+vNcUbHVdyDr+2TvZSNDOupcK2Mb3mveRL0WLT1GOzLpvumFzA1LNxhKpP
BT7BSKKC18H8DAkE8S4AzVAEppxuuLJcYCqHc7CpdiCDWfuxt77DNAwOUnUp+jAu
g8agwogBbMHH9gFNgewIm1rKwShpQzZtLc1Cstkj4ydRiu1y11R/SGD/GewpI8gd
1vlYoeWySU+Qrkk3ZJyako+JkcZ/3SWKB8ADssd+gnOZlbAY/f64WD21nzmMf0V4
MKh6pVvcUxygGSFlf+Hly1oacJhfVeUJsIV3j1W+t3FxRjiKTftfWv0vxqhpt33x
LH5XLbwvzs+8nJazEAb41/0jKrDEOzAjpc3g1OmSaL9TCIAwhzi9vjfdrLcGDRV9
V0ActG2FVp/A6OehQnaeTqOHHTJ5+T16otIFruOr5hWSrKC7CUY3l7e7PYoU5D61
XMn6VzBLfBJevIYyveO793VntUzByLGKYEZwn5EoQdTZz5yvyCfyhEn76FjNUVuL
Ck3H6gtNn5oGeWiSp+Ji621cW+tyo/4WPNEmaFA1t15eDoCX7+q6zVYhXAk76Vuy
stLs28qogygFqclwDo6ngbWJgEeuHe2JGcW7uhXyFoeEUiPW+skMpigVvbMxn1Kt
UpqkVnJPEjDD+9zwLd+Un799klZvd7muPJE3pRcPniVoSS8SG8nCsCbXnH7UeTSp
XmAdkk7K6NedpYAxbY+S2PnLfcOM7u56Jcwwu9B8djTEvIi0r12ZcD4n6DDd93Q2
C+ED+4Qn1/8mMz3qiX1XrJiKcfRp2ewccczrRSp8SbbDdkpqm2jmVb+rwYVLsL62
xewAUaihcjWi9D1UDRhK3xCGDsAP4jPvXFLkTtml1gLRSEAObUgoNlXi997P3Ml4
u0beVQ8wFTc9VsPLz9JNQLpoGUHwlHmo1SCdG29FtSLyQ8yETxtKMQa01ZJNDfCG
uTMdraeneBZH2sN3gRbYaFhQq26JirZYabR4Jc67Q6q3BYdrPGlnt27h6v3x969Q
GT+2E4js3EnP8N+Sy1No7g4GlvsvfGuFjZmYHaP87bIWJc5EJ09HqReZAqb3WVoJ
2yBlAtjboaMeHPI2bV1AQ8aVzqPRXK7Jr5u2cGFygsl0tZ3lE4DmsyileQ0MxM81
hLGi3Kh3HUITuJlgnidMZaF70jJWotbNVKNA/A4c/wat1YPCp/UrWrAE0aFQv5p2
a9mkOJJY4BWlwkjO5NWZv2GERD+Vgwa61RicFfUg4a7o3KwFhZsHRhWMK1BrYo2F
T9+s5kBkFmmhx+tiqmUjYBC+JocW/h0ZmudG15Nuvc8Gr40Lk0R3jpa4U8uOfj25
xwgldJD9B4+YhN8ZEw4BlWHnxY+e0I0YT0CLwSag2cUsVsHVfYsNKpe98S4pGF0a
+cYfPZJrihLobJMet9mWOEKQsvpnz5Lb5sRWAwxKMgSAP3CgG6tRPDtTFQoWUpmj
NkBluhXZ1KJ2gSL9hFnVESTFafRxhjhjzZVsrxOuEJeiPNpZ4N3Sh6dXkui2YlfC
wOR2PLB+GpA+nVysEOTFmhrES2p2DNtRhjVcjHuzl9giQGxew3uyQ+wkUX983P/I
ab1ySy56uMsd09Yt71+hNA7Ro8f/2NubObcHpkwqkwCWXE6wLLZOVsfT9pC5SWkD
K5y2lSRqL3fZxYej0951/8RudBf63KEfkekejsh1r3jcjfqLgL24edRQTZUkj1dt
D0D4EaaSoZUGApgL88r1TLyez2smvGIVEJSUaBh/lga3bxehZTHfKRcrs+rbF/53
yYHsB1M+DzqCL885jAr2Jgbb1JZxDEI50lHpHhJE7abkBtUn6bdMG5/HkoTfG+bi
2+TqIbl4JCNrKFx11fUrI8RH3N0BenQDhbNW6oWLxFENRG2Ql3M6s6SiE6VuY+we
/S3ptIADUid34tETEr6o39944Z2SSPTSwOMJrUPqnCKHAZmdIy14C0RR9QaA/XK1
nE5ocGQOV2Eo77R1Y4YvVOZWbNj3fANfmXTNClEDEDvZzgl+UTmeNEVtXm0NfGSS
kts5q2uWJscpLZZAiiXi5W7uXXUWNFqCXqjRur3dKo3ukTbCaZ7EvIV0YX71sRbK
SkvIJl/jrxz5NS9JV0fsbayU4nVKNtBhonja5NMauDKyYisrXf+y+vjUJNcea8YT
4Q7DSOKqwUYmCqhGAgq8uBQcn1+IO/D/ERuPnyP9R9j4JyDgSW4Gp1XntJElmdaO
5aoJ5f5AUOc6VBpI51/DsdAAa23T5ac/+m4lePiSI2tjeGDntNnZRiDu/yZy88ji
Xe9BpDohjzUsir0cWNJ4SDpeSwZdFWFC+OXCsA1aAxew0cI3NzPkSI/t4/wz+fvG
5tGMwFiBNSzaogecuVOJMzoDjirJCPd5keb1KYDM5waafSPtC2zQtGMb2gHkX3BU
a+3lR8e9l92uJ7Zfq1fuJO7sC2fcJFmeXAa1xoo/RxsBpi92lskWHorzTytorSdU
WcMJNLDwTZsq6va2dNZN7lrjYxWSKdTnySb6vI23PbTT2gGRo4R6EylzwwO22yd8
FdIuxI42boxGE6/AYj+zJAAQ96nI7gEkZxMLlZpLx7FoBq9c5zjPej4KJcqbMhYp
dRAXl7bR6HRhDEyyWtP7NywjYfXipaETPg1xlDsF8GZVHyzZg1oHt5xWCgV4/dZG
H9GDDbZNmeI2tnK7n4okgBnzAHu6RteUF9nikq1d23gMJNDxNB2QEBoPsN2SV61A
JWD6gRXMMMFXlGRTTQkuhRCR9nvIHEESW+uhfjuFOpp3L4yNCc8An1Yd5KrvE3rx
sE6rvXF3Go+6QIph/lanUM/MuW+7EbNnpfWAoZca0xkQ0kfK9IziBUJgwawQ8QVn
CLlkK9Q5lXpqOEfybJDmlG/ALffBAYVTbdsgWqamFO0ntFCWjbZDneIM6Lwfhz4D
ykTJTreJbfTvhSCCHgyMVOPPa/aNbFi4R3Ik6hFZHAHa3yC+9tDTFa/xYui9cnLa
T6ZfF7sqjnDlib8kwwUK/3pHl9+QSaV0qh1YMiT80DhGC21e+2E+t7JLWj3+C1Ma
UV41IwE2KHoxakMeYxMViyncKnCo4dv3zI2v8OHkbLXOMAGsYywI0tjltbzdSGEa
GJImSNijfDj1yYU7oZLvlZIVBmkJQyRsTeg4LJyOx4cX586rAsVUEFW1JuDEXnL6
27P3yQH/gcpBLZT0mbgJJ1T8AneI4WWpcgKDGzXcHMTI0jrAsnUNWoj6HwrIELTx
PGhLf08KXs+oelC44pRHsEhguHuVfGSzS90PZnZi0y2ppDFZwvESl8a5HynVNSIO
mf3/o49djdSFPZ5z1klfGksdkKu2QhGlpvrwoyv/sfNMufJ12LLxujSwB/Q+1mTs
QkCuyuoKfrgRKGv+tcxY5kO/85Au2ksGEJuSlg+iBVnH4ECQoghAEFGSrh/m8KhE
0WuVMwsbL2210f6shD33+lE8ODWvBOoznAthLFyS/C69rL7UfCJJ9iAtjkc9V608
DdEqNyfiErqs1BFJEtY7Op6eW/Bj9kwaGo14FOV63c1qXiL+ZX2OCvwHO+Udvk2J
0+r5bOMiFm3Qdz+kgRGu92ETMCacVxJAu7CIT5+xmIRlY/ID0ydup+WUudXao1RW
nXwng1UyDtkCt/N/m/6IhIMxwB7XWvnr5q+KRt9z2I28QROuTRBdj/ofFAfilwGf
XLbdRXA8ogGWJwYqDXz9e29ddoHz1Jj7DdZyMp6Wf0EG/FtNF80xxo9HXgLIe8Bt
lHCIahJMdxUCeKpZ0uMtP7PMVZeht9xPH0GeCJX2xhKXUavF+rPE2V/vHcTKVmdp
enpy4OZH+v4dZNjuvg59648WX6b/hrneRlKZzLFwfMUql9G4m/F7cWj88/0cr0IV
5rpV6GH0Dzauw53JRPfM1/Fq6AQ1y61pIAMgDsxh5Jvf9gmkJIetT40kTqD0lIO3
snrCbnPx/qLEqYG0R7DWppVVr5Kbf86DNJxNu6R9k3v7T3bYrZ7JGhfiE7Ig36IX
J8Ez1YRgeM/ZP7pftKMz9xlRIG71RpD3A/T5otoOJYZc/reTahwDZ/4mav7r6izl
nMalB6PFQmKxmnzDRMYi2nXaF2YdfWcXLI9r0DyicO2VlPqvkaTFb+Tzcd0lSAwa
CNlm3615H8knDlMuEXi+KzmjMQONn3tVnYWzN6co11aqdBa0sQtYRAUhiU/STJ13
W6bRRJy0lAxphM9Zm7GWmTOod5/HBorsH0jTr9DMJWTIUMw+5b1dvdkapRh9aEMC
4akQh2hDv3VkhpEbmbnZvJ1gGhxLrT1BukPm9nqIzqvsmG2em8Fvk4hoRiKpFUw1
MlusKVDpMUtF6JIXpfyHC3LhdyXOgKAtVi/TsDJ4zzNr7aWGmjuxLxnZ1kDfnXdY
co4qa8AYb1tuwTPgq3AbkL7QOyqYAusL1ruX/YVLsTGhjocPB9W0eA7Ac5mHSxrt
mGmmiZjOhh+AHB+NDp9uW7S57OX/4bym0wMs1WAWBc+CGwsuw5aw7/jcWJDDUSBt
vjGTWGWUXlF18jhMmsSL4n74jMBW1VcuYtKr9HPF0GAvQ+BBLN7D7ed6msEiWhjG
RWaM13DH3ve1HO1e/nozkKKoagvZXBQSj4Je0oiZiLMtY9+mMTtfmuRB4aS/LPcN
xd/Afzt8q9sV54yzVRmz6q1evtPnWD3DlXfe6iuFlkrDv46pBL7BqiOGtzrqXL5T
lPwuUpi8wvBlC4iJTaY05ZDhXurfGF8L+yyQXEmpKuMFkmwz5ahqFXhMbi2OoV2G
WFTMzPbB3MBqv5R7aOlY7qPOwGQJX8H+u6BUP0YWIJbsqF88dwM3ll9AYf4QCmdu
s67tNRZLlKDdSGOig0GMg7hO4bSlRRKymbBz+/VfsYM2E+7YOT1iwGGpVuVyPKJ0
IQQ7YhjljsVcD/3WpMSS14E4niw2lnYBqMZ+eEKJaBDbyrFRY+Ztf+Vjnoci4iMf
KMo7DJ3P8PCPBeOTT1r+5CucMYcXLIMhAF4IrtsGsdNGet9Na/bTEHS3KOABMQhr
yQjvfdPVBp4prJLMtUoMQJwvISf/yBO9mAD0Vy8OUV3hDuS667CVUoW4f/GE7EOH
pOrcxyBhXdi/cyyuCMUE1yfkfse0+db/iOUdGArwpLpSzFNqMJ+vRP5P1Twn5TrD
dcyRKXV0BP70G9J8C8YNq/ViCRySnVm9XR4oM2ebD4lW6U7xQlDP3k8QG9FnA+tn
XkNx9MTzXhk7tjwCxMxZZ/2LUgyC26mvmT4eIxKEZJIccXEcX1GSLr1dPoARqA7B
MA6oX6y+D5t/wdjBsf+4Cj1JQJIioTno9U0hrFVFqgX7HPPfn5CuVJKkj87pWIbm
8o9fitmopF8wl+hQSDHupNX0O9BQL/LrWEKI3SMMbmY1eHuZmnw80LPPWiyek69W
VZ1GsdWvdyX7NAxnGOKhoLRBsdG8B10YXHsK9i8RKQ2q9CNfVo2JRS2kyAT/sAxc
cnThsRWLGT9xcCySfGE7LtzfZ9CkIsA/2oUBLDh8a6xRIVMD8YVgINV0qAWS30o3
CbBJgrmdK1hobK8AMPywbtI1SSpYtPAnflIFLFS4VuEZaDRytlo2uIP8Dh0e6lvD
5qMQ8j2rTJ/f7GjyT2PLZSGq9cgIaGh0lYCw0MTGWrTnLmeQxTK7gKpqNCLUfr9J
XnED59uLuwnTnREbwCyKr0vSrVk/EPzQm/w1uenefOzHdRXwmnZl2Sd+WrYRLcHI
opo1VRJR+KRZ9jYVabTSurIduV26onJXo6vGcHMfMevqwoxNCT5nSyj7r/rHqFex
BzL6UKGsR2EfxMIr+ir1Rhe1yABXhU0t0kWhJ8dsRzQAK19Inwsj0IyxI9pzAZ/B
xepfqG5IjOt3v/G4du9Js/OmNEpirEDugepdXZc67LWo4tEBosK4qzDXOA94NuXV
RiAFBgqfPaV59lGeP8J4je0vif6LZz2NJkRexYhdlZBbon0XIfq8+XeCePFOGeu3
IdLQ15HMmbFMmkZruTxRBSnHzTeoRPg9fsAn7L46ipQ5uuasyKVd/XX7uZ7o0iAV
I8AXibP/Fdm5gxQNjTogQPmq3/WwFtOSGBk/VTNy55Clgta6EhJ+1mSfDtSmBbrS
BT4c7pm1PcGMwNXi7Tk/BP6RoXyrf0byfWmJQ36gKDSwu56QBf2OwOeDouihimdy
vN/Hbz0PTE6RM4PoaSxLVH+u5R/qRCQnefYlXjkqFEHCBhc6TJP/9lFe96Tv/zWa
1CXkkNlvuTxzQnhx1IQzqTC4nHjPVmnxnVhFf0tpE7Kcf8vK4exJyl2OUlLIpG+5
iSLoh8dIjVh4aYvUHsLRD1iZ+ZCKrfye5JAZNZ9VBj9qkp8loR3sUxZVYQdcjoWC
AjftAZU/B49St8bahnYYlSsoQp/IP5bNtlVHiooWqcua1sdnc6Nsrc9qdc76Rrwe
pX6SWzHnH0w93+EE6xU5YB3fC+GEq556tznBr6O7JS4qugJK00wZP1tVWHck0WfJ
O//lCvQJ808ZhYIYFB61toHYB4mMTyv9M7RXDdExMUsUxuPckM9g0SwI/rfTMPkQ
ZhDhc8wmApe0OXZCiOn6qqGSD05qPvLZIUNs5Ua67PULQOgxTG+DQgzDEbnuqD4k
8AJKsbVHAat7gNRkOBnB50lFTeVbslLYhXxN+OHFujdnzJY1T0W46MpeMza/fbK7
Z3A0pt8bAI0WQSUVK9TFzocGFUoyOJAdnYGW0mvuxKYGsFo2O4L6hu9uvetki+9H
MlVQ6BOjPLseqgHbYjE8dS58drDO+kANReC9VoHwDOWi6fYRLXIk08/CLqC6SBr/
6K+Qke4m7aw4vOJrc+2+axa16Vw/oFWKo+UylBZbYZ08g32wO7VK2HzezAU2Xl2k
2n7s/L6+6e5N+J/D31pY2wsHY232rUX8n4KkgOlsZx3WgE4kS9TWxfLh855oTGJl
YcAjTuY995QmR1/wsPFJSrLyLIIwvV2iynow6n1glK1XeArI2XSRVSkD6JvfE/Mi
gI203oXXXzcxltDO8uPaPhP4gz+Hj5KwStDzA8GPWz+GuDAfaBcRwXozQFkKyZFK
QiNxnw6ql4SjCps45cd5+nSv2cuIR6tZ0Erhqt7p8e9cTUspeMOLAaqw6aLN64fS
H7My7J6LkFi8RQeIdXZuMtsVt3yiUDRQiPvXTGdhu8QXI6E+SygRTcwGz2Hq50uj
Nx6E07SJ5nMW4rAawuNvK4Z1tMGlj/vWBGcD7Ry0tqbiojCv+Ndx5Kl52fXaq4sZ
dmf4C64+evPxAq8fsziZEODTWhi6ieoB4fwLQwrRngd1jdJMhcb5M3mww3PftX9r
D7XMC3QQgleVQq30KVw2oG98OJSd8Erhl1eYRoTvi06amaJ+JjccFoYx0P51nbkT
BxLTUMv48TJghLsU8QF5hIBRYzGu5700m6zOkDqTULfVrMTGfobLVdRuscJPniKm
IUBFCzyUQiX2p5UYWrTLT8pIYEMrB44KajqTSqUhRQMeGU14A8xRx8hiG35E2e7C
KXQQolpc+E6Vc2sz68CF8tG5kSkn36L0p+ITuEJxn8d7atKNWNAZzW+qfBX0K43N
bCfUYR+Rkg26UMmrlwvxIgVR6ZYW4i8fA5N2KzaHG9JCI7tkwLPrCntRKam9VFk3
kZpimHarDUcdGfe1TyjhKMQsdWOtq3kad6kiKo7SqdT8YY/NQZXvxJtVAUYzvbr/
9MoqF0UqHub05JdxfDyAGpW5EwE3NdnAoPeBl7O64Ur48Z/+XMjHo0OvUaor5PhA
NFvyk33Z+oA9WnizN7r46WkLKK+YCyR2vhA+D1MHvPTpog3fEq4otb6ttRo0S+ud
ezRMiZ+qn6h2iwcUYp1x2QO2kTJoGdtSThtGuayaq4DfM7NY4XhAmyFa2IadUY6R
0LO57HfvLjkTZ2mBrLsldvrTb2kUKP6jTxohNxs25Y0CqCgPbrwmNdu4efHTFflw
DU8u0ylUyjYAYslt+Opry+SKdk5+yy9fZs0SU70vXW8mTxMScyKmrfPIRLdPZurc
ex0Rgc50KVOvbTg/zitkCO3MYj68IdsaAkNZdAIgcm2SW/sqJf2ZhjPasGTwDN3y
8HHJkjoAuBM3W2KJfHcS/JwOAOdoPkX1vgfws5MqA+lM6+SjZDNYIoINDRvP3ksN
4ktfZ1/f8DnVuBkOyXmBLdGqgNaglhbkPF6ly/ydE6w3eF3mpiXSGbBAcbWOQirD
eWS/f/IaOB9L2cZU4ceRPWBamCrD9jg4cpf+yZXCBW7qTyvvZI7i4U6i6EA9a5Yp
A74XHpxF6862teOiB4HyL21Ykbl/+Tv5/mmtcvIWWjOrsYebl2C9W7jLgKIXcz8n
UOx72CCVBI5VvZaAROOlSRExQP+JueThZdjdXJ9U+VRqmWIWwGiS45xAmEl/0xXk
s/uyKUHkaZkgG8MG3jbnxMX3nomLs0HksN6gUbxkB36K8yRC1E0O+v7jq3HoxE1C
VJt/A4zLj8+t2ZFxII44GuW5bhygj4XNQjQ/BtgkvbiXnA1PmhPwVGPQ2RJ8ZSEs
VvUrwGy3HycRVKRKXYmzJ4ZBxj7sXbgdpKjnQg/Sm64By1EosIFmRHawgzwrGYIz
pRcrK+IHxr5F76G+pZOJfsFUvPAm8sIexSNcEsCQzfLLW+CFHg8iqM8ITZ05ruUC
f3zOVMzXZ7eaZnHf9DOqKUlPAfL8PODnEmpc6xoC4Fy35CrVxsD3Mnx4uejTosCU
UVH9NreaxBSvjphclOgKc9LeoH4TNCQZclII6ehuSSa6+i1jEQ13r1RNJ6+RCC6W
sCUptbNXQkYSyVxBhTaIBV7Mkq6hcqiUgsCui4ZF73lMV2JdYa+KKB+/9+1+4PYr
9IkiePbGFqhs/TxbcTupUhsrO7YJm3XQyjdwSXdsww9kHwYMVUT2D+1OgBe1ca2O
GeOFhQa/sVJi8l3Kuh033uENUWqC+xlOjZ42Q0bSNg76TubWXSaYFrEDGEUMXmFx
KcGQTDsbr4MSJGdDX3IWKfe0gxWK/3zgASv74aulmBgPYqwa5+xBg4VDUDtwn9ft
pYqw7cxnAIeaIMpuWYKRJnuQU8E1+fneaLCDqKRbCmcOTOZcHbq7HPBdfYb5lxro
VHv0yq+hosEdbbmb6RXp4hm4iv9VBULQQAzWOTsR2VR/+ZoZkscoCOVd5dIfQrVi
8h37g+daevq48qZC30b0PniNeKg04CB3QfvP9TxxWlmZchV6+UZALAaMwoAp1Ww1
lopVWJSNwbIT8BS23kragKSISNUmenEVR1/Mm4y43eA8/p6FeHMT3SfcCyGLHO8G
HM9OatQ3A0UbrzJy8cb23fmfQR7YQszVZAPGoxwPclm8Ns4rtORMqC+s9fIeyXrG
uGOjXYGQpYvy5uT725w20xrYH8d9nVudR1+2CG5ZOTUUA7Idi2Nph3nsnNVp2e66
dBsnDK5rlhzXu1UogqIttmAqgpGkT+EQmY+6BnZZfrsu+/VLXzuv++1uW80O1cRG
LW6bxbBcN2BFji22BJX52X4Nsx4gCfmuym4yczvl4k1Hg30sg7fCRChI0za5su2l
Rdi25EiV/cu0LVfH4a346rhSb6pELmgaBI79XfAhUfM7VxDAdOuC6hp4PDQUwkxj
TH7dO51loNXHsFQT+26PO0AHZzQxwYOYHP+UjKyjXkLksSjvi6xz92TBEY9odFas
gkfQumvO+JF5qTMOidfrPe3dPocThaocGATOR962sYxHgbbvQjLay2RPbGcggx0b
QQvk2NiJ9vukUFJ1frqMdEw6tdsRR9DZrISkxoPuJx3anbfWs4XhC9i586Vna5Tz
02bW4YtDAof6g1+iVQUsts8xSIml4vXVBU/qeuYfiPOeosUueJ4G1NRxiGNM4XHx
5q71T545xkKRCyKkwawAau8khbZ+2mjwtqsPrkAfyU+QUUDKozuXqQnIERCE7RGn
Ur1yaRgLlFQsWqaBCPmZhVAJPlN407ggY2h23V6TWwiv+XZgIvSRKc8FQHN56/NJ
LPofAioMkm31khhMOMkIV7bjsNthHKra1bpeipSIyvokoWmJNIL1SAF62THmuSpq
jvvgKqtCQQxiEkJj9NH50ts4G2O8FHR3o7a5fgfHLEbbvvIEtzup7/umiUutB2Zr
5R7bjLojeKGHXemca/9pVPCXBMZXf9Wcpz1MnWlh0/w+fX+D/bsdF7Mf9aSbaJ7B
q/bRYJF6kyYFx+pASWKecC3VrAWV4k8jR/RVXmiPSoLYx6arO3s4fda91ygp8hwl
s1875Zm9ilghdArL5OK9wrot/eNC5QsJ1+/stZdrqsNz1CyNo4GpBc7SvFWxCD+g
PH8LIDQtm7uRujUg5CQ5GfZFnwxOGegY/YuwjNOrNNQSFGBtjm2I+hs1e/ma/T33
0W/T/YYV4lZ3OYPlmm/MZurIR19IzqSJTdQ5nLsFTNSuZ6PGBDm1Fv6bC1B16FKL
+k9jR/b+LHRNsfQQFdVha59hbUCt32iMDarc7ZOctDpar/o1Ee7v+6r6JMOGWsVf
jg99XrHHi08TRAsy/UQVW0ilJyS6G/WeOscJSBxp7bQxkzXYBVXjneIT14rlSD14
eYNXvo2dNjQzv+QCQ3etS5BqeecRDfOtYETXq3QaXw4tDrx38TSfo/ChOyvrJLGd
IL03wLi0AVP06UsLlkyPjGW3I6MJC2SdwmQoBcrS4okrnHWz2Tit9wKo7FGZocKO
W87NHOLmm/5MnVToyUdyZxZ+mJMXlsU3qli8DiPGtMA0Z7cnfSl79vMoBE365lJn
iwzAwXbaV0e/RYyQikv5cRTfKKy7XvJWG/wzMq6iz3iE22OfFdAMGx9aztM3wg0b
eOgm3B65HpiK1etp6+4wz88PmqvKUE9OgKKIIjuM72nj9MC06X0PYsFgiO1Zn0NN
81bocMuX/BLzy4TYFHFeBj2C4cqH481dleCaRgFzUz54SQE5+du4fLpKA/uf4dGk
jcNL712u+WbyBEY47L3mPY1lHVQ9AjN3vkCFVkB4/V1CMO3HzQUierVUdG5Dc1wi
KgCqMiBseANX505fSTkKWN6OHQv1KqRlFCgEzVgxCQsKEMU1ZUauqanqvLZzysZW
B1G0eM6+g+bxCB9OLLIGft98dbGQSebvVdzfJa1pJpTrG7zrW4ec61J9LSX3N01B
1/ItAD1pcMArIzRW62zsrhrBub5lwIuIYvQcTOVqXWL6tixNSj1/3tAMMUdq8fYa
dV9kQamjBUVaXA22UxCvAn7YItaX1z7hf9br1UyzqEWoUsaOWItNkoZ46HePXDnf
GI28huqbovUGUQ21xgXwdhjzBMZ4SY/E5EyvDBSD29fjZ2+pkf+35yKFGutVudhz
r6d5LUiV4eaeCAkFk1OajKwD9N83Pq1N6R2yCHCsHOdfwNopnKYzspL8t8v+Yuxi
EHrIzpMtXTO1CvQerGRnbcNFl45zR58ny9kX3PqbZlvZv3BkMKnLvIIesoo3G+iN
Zmsfmux70UMNJ2TMKRpJzGxAB3qpXJNAJfxQVAh0N2Lpdg3VldL1VKNkpH4EiUxm
itkb538L0mVuer3YH6zfvqPzMkhcKmq/5Mvox6ARR214/YeoFvOLkUMl+mZFT8xy
e518Kym2Mud/lX/lXedklMGfovgmCVrO2ex9b5lrGS3iF2xq/iO+/Mk5b5RgyXFb
hnYozq3XQVDM0USbupLaGqYDAjKrBWNXtxA9y5N1fnBQ4eJd7OU44CjUKnwF3hKP
dESMql+hBVI/bj3tgtk7/G2owcuyrCii/7Z5kyMue7Z5ak1I8jqu7FVzNQq4S5Ku
LYxuxzoJXjq/4B0JFVXKT4sbadFgpRslwsatuhrruk5axPmmqDJSHiwObesmUphH
SWzk1/uy/PJOkaJvMwkOi7LplFwR+28CL/3fcPMQosT1VxukRa8alqXv+EGMejX/
w021RJdO64h6HFGYmd9j7Blrn2jT4a+UnQFiZumir6MvPMMT975B0llTdNSuZy92
HqMdoTmgidrjR1LhePNTo6k61EG4J3bnubZ06zfey67uAADU84BruYFARMsbGKDv
SGMbgzpAdGf8UGPjUuKEkfBb6qfxN+SDdcL4+iBS/+CLA6KKyAJ003cvd/GMBYoy
0avFowlliRDvzwhJ30HT9hBGRpnMxalw4sIZtiML++f6oQqanxin6vMevenbVqSq
issTtROmypTcJbCnwEnpzTrLy4ZsWSaN0H2y8MZIYXnTBgXUyvUA6YDpDk6xiGWu
zy7KvqrqwNIF2QCb4ysQVe8i3XOEeGzV90AfgUHyUXDIYGX5acyhcvTUW2o9ZVVV
Wx+OTgcLCbMQTLqjO5yXHju/LsjxdSioZ68LZUUGJZsbjkZoKjU+9s2a9aJf0U5d
PLVOSr7Zho27CCbVOoTef0r3/MAWBarYu/28ng7+LCD9SWGkrOmo7VBa6JbQMT7e
B0Yq+uE9vsF4+TvK9o0idZs6h1uooAAPSuVSFfsimAo5w5O8reBjHfimlPOBS4Sx
zeAoKcYELTFDvP4qHw9wuFav8G2jCL0D/L8X6NeAKt6goqPyAWXDGb8IUkPWNIbI
zrTqdiD6E9NY8TxxlKNCrijXmqvrOg8AbYhCWCGjUn/SQ363catlisILkfZwwjO+
fUE2dJjcrmUtW8Csy99fSbaW+H/z9Z/MY0+dh2U0igMiOa31dNNw2hnrDrGfxkWK
dfzLwp+BwyE9H5bEmhpC/VsbhyPs+kQvjKm1jqCFKGpEinRt4GlWqxafRXUXcQkp
nKH3JwWeog62+jZjaWObaVDR3y1FJVt8UuWysZzoXzzA5PMRXIx7FEuaUnjkKiq3
31fg2IKb8OhzIdCyR0OwFLM9ZndXxil86e53mhXCzsi/TDtqnmUDBUL6E0K+U+W9
UcUWdXYuTLCu3nGC1VLiPfCEYFqBIBHz4HpLzNu0GMrk/RUeFPtAjUUZTMQomuuU
dS54IYTQOgSeLLqlI+FKnP5nb1rDW9Wg04a8h165CPuhuPXnz5bEnDAXDsed91gf
lMR5qjdEc1Qzx97Q2rD9y/veWrFmn/uaEpkYqbfYQoZ3RxqIwiQXWJFmbL6qFbrL
FRO2ZfXqh8HOGAqfQ/Ufe5npk/ihPsRplrBz2fqM5/44mX4/x78aEu4mrYl+ZVKv
l/x0CjdIYKFR7aGXrk7m0JPRKS2HNbwn3EC9Sj3K+Me4phWE28uk0fdxK9Qi7zr2
Lor7CY1vAnpjAQ7pKE8/eSezFijZdySqX4Ff4wXUe60wHOcPQ2jEvsJ0JBNkcEsk
cOXW7Cru7PkYU2p1o8xE2ppUXQZKZ5H3gXotsn1Z5zEyc52l0Fz601f0J20PvRKo
yP01EnTvtLPY+SGcTUP9SqUq8dxjQzR1gULgZKV5ITF28mHpAlwtuLWrzYWf3K6h
9xqrvK/R0/mK2qQjm8aK4Lj8/EhOUr8m3H3KK4rAh/HkbbI/u0rILE7cgIj9NbIs
MkkdRU8V5jsqmTbuLFnIS7q6z2dTCDJw84LY2/omEY3yKsofbnSrlWU0Sfcn7lTt
XqCRQqfm1GlvpHQJ+Pwk/yrcpxOKH7u6NWJC3OSe8lRlq0htPWmUhpVVOVE3MVWB
8KqeacfdI+hR1WEzTuPgo4OwAF2SwNVIGS9K4WW/CHAU5GGITPpvrHG2ZHzAtNTf
JtiKGoqALcnD0T4eDL2cyhi7Sop5EQ5nZcybIv06euwAwWWDQNtIvgLthGcjz201
Ur0wTkNllG17tsgokP0Ho2uuXqiVkkWmKgP2rGAR5BQ1pAlBD9OMy99NcxK40UV+
qfbTks+UBJQMHIPWajcssd7mEKJUnN3DP6imDkCDWMDF2xnMn1MJMD4PGcd493gl
HHKU1D0SVhoyBGJwCvraz49QbT4hcvp++YyjRYxaf1D93KiZLnugZQB3hgMzIRaf
z22RFzRbVkjkvgiCCtL8xNwdmKZp9dLeBVo78cARvsZaKpI+4lvRphclQ79P7C48
DAgSYkjTRD7ewXGSUSSP5vaiflJCLlfafq32k0ku8z3PvPAPDkIBcPH+q95/KmqI
XfJjk5vkXAHnqvFGwd2bpnZ/2vwgdsl6toxW7Dc18L8wFFcJYAK0CXpS8ZHlr81A
r9KR/03DBm33qoDIA97/65bYCu5vD+kkhQ366HNWGbRwneRVuAhye1q3BSS4oUn4
r8NG+7JchYzrTxNzphTKj7LzKGmB0r/RO/hIAW7Ry6/gO7tLvespedshSuz/1EFj
Z/ni3ASAOMWinTRDZRQoRJHiwWvNk8RKYdIF5XB02g+Uqg4FJnjOfwHL2edXd4YN
mJnpY8tqqbosveDQoentXYpdlBhWit0rW9O6rNhuT6XPSI+bU95R/DJlz0mwd89D
73fcqmG8Gh8LNb+56EHk8ETd1C+1aKozxg9Suq112dJrU206fkB0ecgQlZ8bE8DB
fvEYP7nEjgC97DFc0ii6MEdDKuFzoItB02jSHfsPg4dw2orJLrtVse7wDyL9KhHq
oo2zBndtmu+Q/0T8RhoDDc2egvW9WhC7uRURjJv6vfwPDZsb4Ldu3CSjT63d6A1Y
S5L+YfMSNLDZKSQvui6hXkcotJg6Fu20usL6+D+CAwcl0MqQhF81U5RCSrzW3bNq
+rWhtykvwJ2AqT5j1buC/SHlTCPjwIb+fuJ04L4p5oQ0sGG8sgTJKcvNGx9oBM5B
TetRScgeb7AmYOuKHUu2MMS1Yg7W4AAvjE4JxCamz7pD/Cp1/HcheMa8NHsIxn2W
IyVpy1r428F1151g5hVnQsb+JuvqhNNufLst1cfit4wJF8nssbjdM5Bh0PT6ILIA
n0LgnqBED2UylfntLCcaINnpBSGpd4mP5HSc3vPB0Q+TisILQaEgIoq4+LpIyW91
rjR/1O5LsIl/jLI7PsCWsJwZOpp+UCOkw9nisQtNEF+RyBwTNG5Km+bv3Wm7OVUg
IuTQ/wIRh/s5jbJRyDJGRMJR71FjwSPQ53gcv+L1dlVIi7scyPL/us109D6Gn2IF
Ym5Ob16Rlo2i1hmYqRB/BvEClR3mydTObX7v6PS6hCYFpJjjqARglj2FJAyrYrbI
cs7JFT2eneiYylRrNQuwVaopfssWoyoVViQnjWbBP4IhBpKb+3aSLWN1L59GyUJE
WalMntKJfaQSK3k0fXw9jKYe1Cj1iYF0G6V5kAzrK6BqjyXtekqVmuaMlNPjXlhS
+OcT/ZZg2Q9pVVoFHRQiS/73rV4/bI+o201qk3uLx5X4S2vnFaWe+2UYdP7SgB5z
RMklgZWF2Ivjp6dThdTIIQk+R3QS8r2MkVH2vsNhkIVrOVXHuAJqXFfXX+OHEe45
ays2QZU5jY5c4fHG9V+Ta3IGzBWsHR/077qoDXuMkwY+tgB5qL8rHBVhVGe/67vq
lVbqBZb/IukJCWcnEJ4XjO/RwIEXgqHYt0a9LWOaeK6zR8US8zposoyLiO50wwFE
nUT15GZUxJr8myCFgGOx/9shjZXFDCiHo0a1LJDRYijRCYrtUiQdSRP4ZFf1koX6
mp1/BpN5UJn6iYDghWfTlqtUVwPGaP2CxbNSRSp5TpVI3sEaL6WVNn5x+mvIVrHX
sWCTPGielGPwlJAPFrJmjv3eHdHPb+m2ZuibugEdXPUvKPkNZu7NQvwjhFH4fA0W
V8KF1UGPZLq+m1MuFHCBi+6chIdQrmq5GGPue0s+I9cVoSETDQyXW+88dWZF6Sc8
ZA+8IVa4UdMZdqYwSdhAFN/KwQqhpCgEOU7g/mO1XnXIvfnWH3Ms3mEHP2EaexZA
AeWioWJzg0Wewc64xKjDd+SB/yWK7ycqhYNDedTfpW1lY/Bb8Hi6okxjAYTuue6b
e7WTcq/O7TAYXKJHPFlHe+KUOZccv71RZKu291E1wREqHPchBI1lzywx8wkTJ2nq
qd5JhKK/nkN8vq3zSRLnh7Srkv9ih99a/8/6LGrGob7/kbTfFrFEohEB6WBLYcBK
h0HjwfPNdy//ezE9duchc3LfSUzhGOj+Ec9GmZf1m18EEcrIs3/GEFkOHKibdtCT
bsM2mClrwbIov1jkL4xPTLsnLl4vIwjvXPkQSMgI7UwUmP/Ncn39v9Zks6NHmFff
rCTktaK3to0h6FvnFpeMbaVLsHJ/i5MuVuR6wZ8JyrHLxyZ4oqyy5QG9STpbVBip
p5+GXbkpDvlX9LP0mvX3EhCYnqdTflPrJNoX6dk2i9hk+zaPu9vf+Unou/xRAu7B
X3F8UBMLJ9aVasR6Ze60FatDANhFcRsWXOwnwy6yImJXicBSZ0Iyu+FPgnFyu+4s
Lri7AzO1z4A9HoEZ11q2fdIxXVDwwlEMYDMVwtoUe9u6GG0vw9g+M2D9VTK3pO32
dWkXENIA9FqDQ7RTNfCIqbr0OVwmOn7x7Xv5ItYxPuqictMv7S9PSmAdi2cN2n3B
9uX3gbr/ohkwjCMK0W8r5JzpgWrAug8qfmnTByw+FcFlzetaJW0s45Ngye6WVD8D
LAScf9UMK7xcHMv5wO/A32d1n9JfyujqXgkqc9luh1z7EDMSYp243FE+E2eJRqA4
BRyGpUdfI+gh05Sfj1RlFe2g/Ha2kW4NDmNK8OZeH/8E/y6aa6KUzqAHHp6U1vkA
KBvehDLPHAZW45U76jZmKd+9y1VhaNtIgvows61xbos6D0mcNoPbI3LS0t1A3C7B
XQo+Rs7+VhaFGjUZa6ogY8Ub9ADbe/eJ84cS/OD8h8MSPMS8Mq0OrZbYVAdEPO+2
ecvqMuBNZtCOic5jzQWy6V+xeq+0lGRPnfrOnC5zPR/tG/hTvaXt9w0Vx7kAwG2R
7r7lLOlATeQZZ5w5TCQp4OCJY2N1E1Uz0DF8GUdtMiZpAtdujmFslyDUBJFB8ogI
avfkMMC85uMTFH7LiGCx4qBgxpHlxnucxel4FfbECDfZTQmiBY/Gj8IdfirJg1WS
XdOkqY1V/h6Fqx6ejIdouNxfwwDmjfdKYWArnjn9hlA604/8+moWKNC29aiK1AEY
e8dTxmQ0FFA+IGBzoTvToXCTNHfun35BgKw63mIDwQUGO47z2Dd/k5K57M84CN9J
zS//iztIvFyUqPskjNVYDtXm0KSZ5w/XDo9DkVAS212feByZgGYENkbQbb7qE2te
6tgVP6r2k4PSWRBRWYvUnHCFZgNmsQCn2CLfGrKNUiDdKdQ7gEwb+1yS6WdDk5k2
tlZry0ozk/49GU3pCKH07nig8DaAjA/DjotpAcJwl2G6k5fLODy5KOF99Shxr+7N
WQPm5ZcO/kIgbzJ5j+4KE3d57lWB570JYV5GOPkC2loJwE3viFLhYaN1mRkfY2Zn
q42n0QUvNnLUgwbqsjGfXsSXZ42e6dngRyefCS73IWSAJ4xiHK/jBqmLq0O2nOTJ
zZ6beWmObVOVHliMA5jp/n/FkFPCGzyRi2SfLoA/RDT93D5mNWHel1AihlMc23o7
xkWGBm5X6+NLXKJB8OwOvu7quGnkZ6dH16bkubvEjElKMo1/7IKuTOK5lmNkVRNw
kYABOSiIMVHBQoh4xcOr+2tR/nYovaHtjdTZ08HlyYszVZ4yCFwplO7CdtkmYYcv
Yz7witcEBpfku96K2rNshGwVa4HL1dHqUOmVET32/zvTBKi/gKnnm+o83RycyV8u
8o3zDrmYwQ9z95XzO6nn0OvR7CUU481wDUokebHc5Kj50j3/p4zNc2E1Z97DGHOP
8nHGNfrxzQ0vDWW8kzpfgNn41GKOpZpGOhhUybzBgaCTOPMH49jkfkFZ2rd5SNhT
yK75+w+PpXGujC+YA9DbJL9YOd5Jyy0Y7DIX5bpRzZ+S6A68LZ9ovoh2tJbUeI0C
IwXgCfWnkRWcA67M6oQxVRIGS29Ym/ZlJJnjXSY/Ox9b9PQidME9HisSQccVhDHU
uCqBossEFDRLVHXPcqNw6fUhIRQEEP0PF09D3RDKVyMigJrf9fQ8nvvDFpkB6a9o
mB22SrWJ6QJzUEZsLplf2J9Ki5wKqZy+X6JmnilI4D5yD0sGDWDRvetFtRK8+X6N
cqOK+poR8Vk3Cg7nWXw2KzfO3GXsI27i0rtkxGWMVVo07KnZpohjdjHU+jtdqnSl
IIIGeaYySSLJrreLvMG2k92Q8eMtdcq4UxX+haiPIfg9FOg1vJY7VCryDG1GViVh
1NXeftvhM/tF47T8u9HL1kwAXpjFYaf87XiyR885tRc8lD5tSPuhgohzNZw0V0KC
4N7wi1VL7EPqoB8+pvRUqeX7w/55kc9dIxwqoowzQygMl4ZPAB2TFc/d2ffSmdFO
trvy8WLo1avOEYz//4ANWPHVdUBylVz3G//odrrqiJ0QBUZw22fJp2SEhsbqP5jP
DcoQ25i9fhCZYKaQkOgKtRWR1hRrjYS9HYotU8K9im8f01DAJjSZuTLRyB3RbOxH
CZdAoouBTEUoLHd0+BTmhSuj35GvOBGlsdhfAFxLtyguN76oaoehFiMIUlyXCcAY
UQDsnml+zHxltdtS9MivEwsbnrJbeNy7jB4FRWtg6mzEuQi9ONkWW5NFH9oKjSEE
5NNIStpp9oH6If8OFBWEC1AWsLO5mcYcYHY4dUIy3oNXOYVTtbW0acML3CIN8+Fh
VyuaxWaTOX1wbJLygS1dVm9xpjqpouw/MzToRutPsLC5pB8cgTgBMwfd6DiHRZUm
lOj2iyPXKJLipM2RA+XtGK5yFP7SebzsjA8lD9NsAfn2mKYuc44jJ05y55X0Mjvp
KKsgObBhFyQ+TbOyWXOPAkIkkbVXp9G1H/tAIeN6ondyZqrVyQU4Gq7bXaa8Sxh+
7X+wtH9HFJq5DdZ6wTLNYd1wG+yeZqek4P4TmyAnEhNQdo1x7aqqVMbbZV+vu9MI
XJtHrsElkpbNOfTJi3QW52129kTRoPSbvOrSTJIw+/r71+kLDATK1fIsYp4T6m5k
ymTeL/TDYqmK/G8bybiOA3kjIeB/vTlbQkolLhQui+zg9dj05tcGH2NraqSzQsbn
lfz+04NEXRoBiEJTfl1dkapVqSCkkujjuKFUlWMYS5pc5igqDpw/dC1bpnsQA7jB
KHARnSt1ajgwJgU3gmQmsDq/St+TnUksRktG7tZXEHGTxAklWVihldRFsH8QIi1p
5pNUGfpawV22LtLtMYA6VFcIXk9sYQVjauei+pAYaaHzAJJZHAP6r99K6pf+iGgk
tIhPW76aWvINbo1R6Hrw2geH9gzMY48+kjKFcddrEEfn8pqHZQfuey4eW735/Qx1
mdlAbOQIYJ/7D4sjpefUrC5nunDQEIRgC8h/RcqxlQ68aAXkkE+1s9u3u9cSiUpZ
YPAyFvDo+w5Ap1pacbmHhpeHoOx1I0nKn21mNOAkVYHzx26u/3t7vCt6CxH/ug6d
MP0XSXZhAc+3ZZA+yhdy090QmomtGmh1JRJaXtDI1S7iGX1CODdvCWmpu3aNoOBH
H0w51nRrxxhcKwxIB0Jf/zFzVVrQEynS3NeclbNSV1u7TapzxStIkkOO8YHeFJKk
Q2DfWiVrc2McuVAJ1kRmfZjXzMa0p8LcWRa63dHL2B7s9smiZF9tHUVqz4BB2FJS
fhPK1ynjAB1QFvrcObDJmpw9Shl/YjgfoBh7WdXBfvn0Tb2JadGw1Lw5A0TJ9fAP
W+nXZG95fo1rPh3/OrhvnDWp0xmm18p99BU8SDpLEiuA38EK5DWM0nIZscqIZWIJ
ERaLwgQUZZNzF4ZM7/yOmJjaf7JuYglxxa7oWV0pga1gpQqkMlhds/s3tuiDwfRR
ouMQNqVZxWMLjwSE9s/DHByCH0cSrHno6fKUptTYTJcpwhXm2nqpNPLMyNnKtKd7
zgg0UIyvDqxkTDxXbgIn+S0QEZ+1xHr0AuinEktTFFFcaYszP5SOQmpEZyI3/em0
hC95hCHNmC/g/YqnMmk6QG5RC8VMNiByihYr7ehGYnfS1fmW4NWllLpfcSaLhKE1
uldUBdrhytXqsMYcw9zwSRCQY/RmZDjpqldY2qG/eQBokpB5iHp7Zt9u78HUtvvp
Bm3rdEQtzHrNa7VbV3odSMOjSSh81m96IK1XAc/+Q7/XxAwhI+W/4Bdkkyjw8495
MUnrwFLvauXUVnOXrDS+7xwsL0RxAXgi52yx0suINTu7uRx3huWfpJfgcKAqgEMt
Q4uPBjVT6jg1NFxGrol6R+VmQj3ZWAXBwG+DtfYosRDiJHE6LErNupedW9f/FWOr
HsQ9tSQiiFcMBfBepXEXwg3/gEkKuOPAutlFeyap7gutRfPJHq3h0nbEVDrCGeoM
N+e/nJjBF068PU+t0zGLRwHAG4lOdnsIM4QKfAxEYAUc0BNRR4EvPQpEwa+R7hbf
VV2eShr2ZfW3rCTWuOKkObZpZgIOIbOFhAIR5xsiBdf9V9zMWM1teiinwVGzHh3K
3xk8S7rTnNrpWFAd0Fe2QnLU2QE6x76pPAE1r/uGBXimFHc/v0CxxCYc/+CZ0oen
0Ye+r27fK6U3tDN3Wky9E2KgnbQ8sEMhWEcmoOeHMQhsjb7Y10LxDqCo8v/NW+Ok
oHUUBJcEHec/EofQj9qIEzzF0cTLWBfmJAc2X0WHHQvlo39Y6X2nSmiNojtkWpwx
VHfukcGM+TpsRSi3eDm3J/514hly6+YlrtvamTRyQAI07q260bKY01fhp3L/e1Gb
3kX3bdn5WVrNKeRlaZfme287BoJAfTDDkBirlc2esw8cG/20VluxIYJbWNlOCXd8
qNwh6bkO7cCpYAk6B0XCnlBERc2O436jvZSRjXSyLDhqNu2MfA1RKRdP3C06FAJ2
mldXhF0HiV50uAeSZDG9StVZVN+AmjDwbDs48Cs1iAfUObTwYsrgCpVNpfHvSlfY
WoKQSmpQJi/jefw3eqVv9hJPda8Gb1oRCzEm9wbHTVi/PCXBrkIE+jzr+4Byzgvd
XKEuuBTtNEDPGegOl0Ah2Y+uZnscrdomme71HYbdOK7znp44xm3be9OUnWI6jTXk
1st3RRwpJX5dmi3YOjN4tPTxK9qSZvFLzI1b1s2hNN7ZQSkjXKwzSXOLjFe3zwXX
knfQXtkW93JiBzVCHv08AGTeZI/keARsiM3XTRQLNIweldkDH4Pr7G38TOE1fwUm
sWvp5h60TzAyc4X4vMK0yyEEW0AqAWCuVrvIXtpTRBATAZ1HbEfiKzWHhPf8Xp36
9KhTFuvyvv9I4HclaCKcnvyrL2YcLUTOvOaWncgO9CK3PcLGz6sF8+zLTSsqW8vT
kTSi6loacULO/6B2npCWvaXTKApPJW4DGP2TepKjLoq3ex5D/a/CluXocPVsSNO7
TZqJjsZPo/ksxA5iwKTij/YNIrShz95UpeCo4fyBs7p54jHAmm4Z9PahnO3RdlkF
qpVQAC8BLBIQG8WowJix35yOG72brryWnI0Ue3h2Q9gJxm2Hh83u10DaGIPqFwKd
TUuA5wDpqjObpMNgq3A2MXj1yHyWw2F6+dX/AhfJleVdEsOhUETYzEAr49ayOiHb
PRg6YX0DmlCjl6uB0TcPp4Tx+SE5f1Wke2M+h9Kk8vjEA3cN67cXoT8Sdr3R/duu
Z+oIgkO8zOeUNiRokY5ewiTaM8h4HprsLiaarklh3GCaPW7hbU5EdBTegkDLzRUD
URfBeAoj4VfSsYpV652DMOq/QKGirzyBpRGdpytcMy5DMAdrQD+UisDWxOGHPXN7
4Nlf3CQFR2TU+qIoKoBdTWRewN4hALTWY+kYviTd/uAyo9b3zGjecw6s8ddbPMIa
3bwX46jV32G9QSfOWgll5sK/uuXkjjlaY6fujxIy8oYbiPxQxHQ/xjrqE9iXZdVE
7RjMRd5z/zYhfnauhnH1ec+AJnLhAklfFdR1wirT4ybdz6JUWp1uILxf4UREyDgD
/YL3RJAC9wcSCwRajC0rF+ylQjX2ISFAcsqrCpo6v0hctDsjXkPc8YOfospT2Tl5
yUlW6WWf9u//Y3W3kad5RaG0K0bC7KPpWLTAsPGTEhnF37HO1Nw5QWU6gRPmZDmI
/Q5yFPag0vhopplWCz+amHU+fJ1e5l/+rrWCjXVGk5oDMNwChZe4/1ktrrO7+IgA
CMmVei3FabJtHJ9hrQZqyVh8LylUFcbRwCJBk4SNODwtFIk4KPDZOEMLMFKV8PE3
z8+nkAdpkmGXqvYRdFRaP7iEp/1FKOutYCmbhejIySBKOo4JPpnlxDngJZo9fmIg
G6autc+AjSn1WWkPeZrUlrBNYNCKABGtlvUil0FpIZnTaQlBAsEMLqzSdPUc61GT
OKW836UgdHKeej3it4d+cyt29huB9G79LTcJ1X3+5FfxjOkL9Ydb3QjDrtBAdPJ4
p2hfMGYKheA2YKJz3Q67+dqprrXdxBy/tAIndRpsFgjQMIbbAGZ4WNL4zHZkxu7v
JZlfbnFvZBfOdXYSmhG86SLm1/6doTKFLB69sq/sDIFPs3jw74ielA4oZOk4s88Z
yaIqB9tIR+6aniKeE3jP75KWUZ3GRsTmKhFQnfAhaM1J1tsPPyQ8aTcV80elf7cJ
Xv6PqsZgEadLazjHMMH2PvBFm/8Ep33icKvFfyqWFpHNBD2unSShWGcj7ctDrpXr
9pFEVjeOdQkJFVD8LWsw6Lte/nMDxyUfpNFzHC1xpiqcfr7K1RfUDmHjFDo6TROB
0UA58e9HzGjlf0tgWCQ0kEJjpKnmX4pTB0jprKNwsp0KosGEyHGOjtnzM+ZWqCmr
zoqAX9kKu/YkGsb/2HqY6q3fok1YApIEn60zlzJnKvYqlRSAxv0L34YuuVtyoBtN
bvKfwcQPztQvo1glUdrl0b0aJ+v/TEQgv6ZP+JBA/Ex69YVeAYU15RICDOoSMPDb
QzFvJVPof0EqtjO/yCuOnYgtCX8QSbp/tYoR7fkB/bNMmBNIhwbVLgkmj17N4xz8
vj3CA4rkj0TZMEuIf2738+RRxIX09bwqcCFagvXCfY9cuMchM/r0ATDoMsY4e02t
pjUZVWTpkDKbpkBl0PGYcZKiuaeKIWK5CeieOffmqUAUSTwP94G4FYzgJpAumb/H
cO9UcEH2vYXzrIIy0wf5/O4OgRuF9rlroL0YO3Dyq5JQ5zr/uiHwHqI8ZTBrBCeS
XlzHAsdz7W38GaLpZcF/RtzTsL9t2tLERTtDQUj1ut/57pdAKSV3SMnw1NsfMQhu
meb86BL6IzB1Tc5KpUplGojKnSLuRBXrZ6fg6i5G/5/UjU2cF0luovUMwOAXfz1/
skKB2jLDiFJ02uBv4/OuUlXl8tduAbu8GUzMsEPt/MwlAcpU1E6J4YUFDj7lfpbb
GO/iBfJTdYwbin2LldYBYNht46x8yladzO2+uBtjKDBUYZ48/OxTsUPi6mXNGszi
0sR39vpyt0uRjs/uUfheD7lti5Uh2+gfYd/+3S4phGmrx3hswXCEm3ch+dfKowWj
TrCu85RNVTDnKvfLwJCczYBWWzccl+iItJEj2a5Jz3IVp8bv/Hl8UPvGlo0NJg9l
qCYdGDxatiaNlYswDT2xkXIjhTbA4/hLRGIlomu13oWee3GG1YSqza6C+KgyppCD
rbTaavjQQAdn5MMKYJzaKvEFD/SNSpuaU4SOfcbVHWYZC/wTfGYy2E4/5uoN4K8W
M3PNnLE/F3DPwM46GOL80w/iEETUrSkHUpjVsrTgpP13XO5suv2abmeEA6e7R8yq
eN5c7vAa/yudHO4QoKhFJ2P99q1kHSzI+RtpC8rXWsJY/Rg2sAc/gYvUscgNlyLC
ecv7x5X3L2UvuCsMrOa9GVNMidGXKYFR5mGCX2jVbOiEoA43nZTxpMhGeEcgS88C
ijwuF6rogTBeIN3hwdJqeLXv++y3LVSJoCFphG/z7AMGYQvT/b5PRZ4yKG2TSKDI
nPm+ZC90sfJwGfmq2pkFF74RizsNF2bRE/pOxMeGIbxITJirnwe82oyXDyDA8qvU
AMAMnAnCsnoi5OMQd4geJIExYsQjx9F0jTjdpRYJYFArfaJSVmJdVhdO5RWJ7Ed7
97z3W3UA5xekqqAa5lkzxoPksZ1Z8D7+SAhDhaVZDHGKLbXisIrROTkqaQiNCpOP
bdgtbMxaNxk3hEsLYoDyA4XcKAlCvO04MiNBUm4awhtACE6R4z3/BGtYmtOdX6No
Yd1B05Rc1pywhDe/VcmwSO9Z21CiekV6lhSFFJ62HWUS8FIEtfGtWfEUfO0bAvjJ
PKg+QOmZ6/MOhOxkSke4zME7Wqzt43gVHs+56BqFemIU90fJX1JGJ/UppR6yRxZe
RhaIEXXDYe6gvO1D3tOEgPpo08UzaghejKrfrpL3+I/xPTk/RQtFbSZi6D4eImFS
X5DkeAhugD8ttJy/vlvPy302QB8CRdebU0H3cH8hFyTJ0OJnWdZO34vasJ8GSLhz
tjPHrBDax9WoUq3ezQ6CDf4XqDh9AJdVfz1r1XBKFSw7S9wPCfdlsJ7KQJT3xler
sEMlgML21mJfC3EOhfnyFOImd5TKfu4bYzdcaKHtahFoFydfIkAvXbtNvud9H3an
uhBCuN8ZA+I9uH7jmaae7Y+5+2obftg0IrYcZKmIP5LGcc7O/X4Mbid2wn6NcN8q
OkAv7qqhCRvwfyxHMDaTSLp18jkCpylqBbWI6kNij3MJGqRyQxljiE49lFa+Rl6d
mHpoIh+MEvXPO7Z/xSoiyThJO7ZHl1Z9Bvxs86AZNyOBSX9FCbqK2xCvsvAB49X+
oQIzdcy33TvV/5j4wa6N53KnWrToTejIVPeuKODBGLvImyJ+pAhrvzLGb/dF+YYB
ZH4+nIFwMn+nneRAUDs/+6Qb/gHn2xSeo4+G8j7oYA9YPF2aMTADdQJUdNcZE/6+
uSJ/ijDFpMOZL1G2qp88nGn8jdphTMJhQNe84hEIM/gJQyE4JV0uwhK2kpWluM58
1ytkBJZKQmcns0VX6spiaeKDwB2U30G3YHvE0pcWP7dezyvqVs1vFTKvo1pVCscl
/cuthjpnkr6tYtnRfc+OUjsBwLUCnAFHy7866snjOKnut9HbDI15klHQ3l2CXhYt
UlhCbQzCKiNWAYMmUtYabEi0K8/rxFc3lvtJ67JydHZ6YqWPGPEAWhprfN1OcEL/
+wWwtwXmX1BjGWBM4xaoEi4BKY/AW7X4eGB9FYXmVzp12Nt+em/s+cZ9JeYf3mdI
Nl0d7qcqNfiCQcd3lB/yTiUMDtawtYU0DUqT83emgogYNIwSpLPvufkmpPV7RfbS
TtaPT4HF0tSiLQUp5W5MhcOR5ydBsCh7m5MAloM88/32uoI7NQNcWLJSg2DvwKBq
cGzLcM+n2B+vz8kGQ24oD4OEEM51P39pJemNOWlfPMR9PnCR3apLOxFSKku0Kt6p
fNxRJ6RyQP2YTEjojILBH0kyTp7d71s/cKRX2701WSNTaUSTU1VkmjZ4zxJ6Tk0I
OShVRcmS8GCx20GloXRy0nerU1pEHP2SSGm8vzLii1PtYdBELxUvnGgAA6mjS31k
z/TT2Ij1tf1wOtz4XZtMWtW/63hXa5gBGqrfE1H2VfdkN6QcV8xPypheUKB1cFgJ
Cz0sh7W1DgrTVGJNk9amtNGrwe8n2VEYh8WthDzSkx0h5rU4AX5G2OJRlNuYZevK
cgUEJV05vjB1SfEblAd7zG0m+6X2h9W9sjFNukFmCpFUdRLSjKmTV2s4ze5XaVp4
ik5+V/KgtqRL3QX1uCI8I412Pwpb89NiYN/UO6GeTOCKrhyHS1TZtaLbKruKJ7zl
ZL6iZeMr2HixlxtCT7HICo303EbkHH/Se83C09l7Lt9lbMjZzLIjjDoeDKGQ9Boe
PC0jA4T7VV6QPOUC7smNWk5/DpDwM5WxQcFB2C9o9gOgSOXH3at0yO0EgvmZg5xY
EOdp1ov7t0D362R04AYYiXingM2wCfj4JKPucSJ3KHT0BFxVN5VAOjPPlcDa0XMM
kw9glYQDgcGzF4Gza9fpl8bniun9Jd0uHMs3YjNzmMPZ9v35h9KxMykOsYhZzdGn
4mSMa25lx1LE7WVItg+1l+pY8/XhBi/BbY9fPx2O40H6P/n2wgN9hBGcfnOb0HNI
9s+3gh8Su5ppxH9sI5IJpNn9VhVv3Z6docJLVfj3uLVh4b89b7+T+rpzlmRqPyJh
nJerafipsmN6t72aDhl807ab3yTjeX4gVQBsS76tUe4pTi7u/M32g3/kQfJ09qlJ
NCoXjBYFS5NyraBKbAXl5zRIQJZE9V6KFJ7a5wxV8h3CYpFsZE/u5rvdCIkQP5Zc
1sa7y4/dltUivph08MBO1QK6UKbMxs6aOiNpN8TBDFKsL9zCQQbl7FMwNoQs79HI
ObNtr4IDKN5QEwimAQfgRlLB5iwBWLUjcyBV/LSKpx+ikG6G1+vcG0MKBSgGOY/D
vwNVT7xOwtGh/tne9fTaXzHUpJ9v2z6VBDA1g1qJIgD+N40tcmr0HgDToZvs4wZb
jHzb/+O348is+z98SHXzsBjFJZz/tSjLNhQbVpjrQ+3qzbKXJ3kmJQ6Q1yc9eOG6
9rx/Lg5ATEG3LgcyBLZEcv9KQPBk1MrEDB+XWnMyti8AatK4lteththq70pyfB8b
QJSErz0Eazlwr0Jk9TbMC/DiUdspP9b5a1uZKeozla8pRA0a3CwhTTEWRGYI7QP6
O8Y7PsKy2UlMYcnmmsjYOqqsXHTkqLlqHMTQdZ9jKfh+rBRNv3pujSNNMYhmZGiy
G+UCwTA6wOIqJkP+Ix46NIz6gEYW22hPLq81YlyfPqyqTz7jK1+2LEf4T/VbBwPc
XchyJjc0GL2fePAlFjU8jnPmEmC747X1KCiMq5Pyw3oZCZHL1RJEvyBAXrzYMIXB
fx+9tfMU/H1XDM0VX9fCpCU6etc+YTuMAszUBnfIdpFQqEq0sBhoxGkAmH1ODNPJ
gW0HQMeQrWxvcXeaHXOtzSouGO+g1nQowxY8H1B+P9b0/iFqOKQhdbFDhc1SENGc
c+TKO6W7NWvyVWwlYZSIQI3dB5Zt+qHSd2r1eTB/L/bTScS5egWWF8oWPEWlVStg
+tNS791D5+0dvxnsjgqsWnx84UU9497GUG6kL4dKV/NhwRNa23NL9jBYaU7q8bJB
SBzprYSm64ncNYp5uMz2lQjkCrvrNmMT4a5hgbbrKGK7Pz9wkYoC4pqf9tgu04al
xjKuUbBkDYv2SkK1xa4G985Q2j7xIt0SSQ+Tpd20FMvVvXNt1UoQNqSZx+nTcJAt
CmTY8TcugWMqY7KlEmDBJQ1CqvUI/M7yh7zUQXpw/WXiHhLWk+PS1LikcjUqCA5J
cOXesrixdREJYdKwvBq+9T+pqM4OM5q4/F8Yoq56VBOaw6Bbut4kpoOBUferfvIk
1h65kKwsZk4rD20d4TbfC9uFLRQdTbdpQpxssmoaOOTL9ZyR5ZWCL5HWiepa2VYb
xCcDqNQx5sUbSycQVY0LYDJDcsGUK02NaWDAXyMAP0OqbsC8ghZyV5SgM0grVC/9
ZDjudgXdKJHjen2dXpaXhAKAjxW6tjbaDx8n2O3ixR0XtP2ABspwS0RifXmwe+g/
PwcauT0kqXRlyjY6MBhfP0tBpKdUN3xTGnnQ5rw5pwCA32jhx8hAPoSPFN0Bo7eD
iPS3Tv0yrMBhfiJUoX/f4Wq3MB/KNbtxGJ5qBeH1tjzC/Q0ecK/euUdijoHJ8Cb2
Mxhtk/QmJuG4nmWYJbjXMGrNeJzRNr2LbvnlzPXREGb969HF9moI5E09p4BCInIc
ihIEiuoRpXZrj3S+nLAvVUd9XruPje9A787TOieqncfY7NsAG+65d0RHbUfplyI4
Ey4PNub8MQ1bIUtwJon4VvWvU4HfhlSgc3nrhC3YHx2dTYMoXxsvFG1QU5TcG7Uy
B7xbsstm5CsDVE9b+CFRmYjxS9j+Vu1P0B4sipyxIMuNgEPlWWO8AtwXq3m4MHl8
CGdE7YqCFOoXL4xrdCAP9erW+4EZPXxLLJbvV7DYsLlMviuNfZ+vDzta8KAdT2Dz
5LJjwfwjTAq/QSR5rLJeNoW5/9mWGmvtLSWwGEHHYTbv1csyetYOtzcptndUUG/1
IaXqLGdlJ7LvZ1Hf8cwnTEplk5fGPe3RgW7AygDE64FUkKExB7p42eyeOfJqYsl7
eLQZodPwww27VRYT2M+67QtU4DDNdEHX4vlLrjNeJ537+zQCVCWNFAbVbytvWWhd
eUxUun+x6jW322DQXVpcV+zvkz+XDnS457V9rMdCnnTeDFVLd0ZeSY9DhssH2URI
bg1l1LlPuY1jiM2vM49xFUAQ7RpgnF6o9NDPLABP+GdFjy4fRhYQCPp1XEev171g
DJJKT9stYz1yN+wotOPgs7a+4LF9UsmqKDjXjwKEI6FUTTlwx3fnArLI4nza6DtH
IcIFgFmVjic2RqRGc2Y/zRGMK4OORS0JsBeWexE//FNAoZJFuVzQ5pmEXzK3mlwh
xYzbEgMkgTlgNOocN2RpdgBSLtIOejPsgb71yEjJ/XqzARblvLt/r/DfKG4Vb37V
fw+m+vJ9dpYQO2ONL85+fuQSAy8nsdWb67jL5bY7zM+wUzGDk651mYEKS8lXgdKX
cP7taEZsADk9Y/aBYWoJDLfpDkazqeKAL/cDkQPzsbnnoLAvU648NDEU/0NAGbhp
ASAspLk2xK3TSHvbXGZM/63dbRx7FtXmWbibvzzTgHr0NVjsKNA74G0MTdT1HKwC
z3dDLv4L4V07bQTtiME6Vj2N27uNUts+d/YdxICxJZ31MxX84l4UBx/oa9V15GWd
msr2pPbOFoudPOcSroFeQ17OyEh6qlE+OVJ2AuZYrbcvSeuNV26a9HV05AiIKGHw
YWFzZVeVUyPQpR6FuTitBcT5/592fg9RioqmdPXxvg7RSoLA/PJYBcSzMeFnvey0
n7r1jN2EwZX9o4jVZH9OBr+zUWgRdSrPkSPwjkX4R02uH/LP/SpvAS/B1JklY3Ms
S6idwjdv59gL/d5MsP3eB/BNlG9ANioTHR9+BHuKAoVKtyFvMMsEQuCnGADtWZEp
UHGRwCGmSUKhsB+xdD8F9bvwoLHWpi25fOYO1x8S7jKC09vB9+vIqw1e7bmQLbEm
V7vITzlV4tC1lS9LoyZndUSgGLqGlKKG4YK6JRixw4PJdHB0mk71rEbMM7piR13E
Tb98gu+JkU1uSsc0GoMSRFvjpK2DTQhNBjcyhOiS+AKuBZ7PeqKy91AHXtnH0I2p
M0/zhH8++fVknAA/GRaZxqZdMiuZoMBuhnp9DRnlSh1uqxDMs8StdyNprsORhRIx
gRQqZBxpFIvVtmMQwErJ2mJ3IpqfR0fZcWy5TmU5rcuOl20IciVPGmSjDOX0bpUI
7GONZBdbQ30BbcCMSUCSanrhOepmOHFn2puX8JyrKSCBdhfymAt5Dfri6x1HxPck
d8/RF2sxZHIwfhYdzSt+cUhGWyNNNLsrD3eoOQ9Vswm46TyQnS+H9ntR24amyqB9
ZJo4tSHSk6rINtJvaT1KkWeXYgfY5lHFdULU7EUNcbL5SKvBNjlwc5sVgtzACTjB
YFp6g2hD+41wzriQiKdZy2EO5Hn42PlR5ZndzO3lK7Pn/wqbxH/xHuGuk6a05W1W
wyi2I3S0FV9UfkrpuKotC0BGeAQQjmbYcNx2PR0F5ZOlpt8hAQne4uuPo9KP2lCd
fVQYpn7NWr7KXzkSsEu036Iisq3kC3N60I6KbXEKTyy6wyhH32mPJ6spo0FSUS1V
yl7NfDHHMDePCCCEwv+H0y9lOF88xygIjA6Xgg2GGTzEmoluRBe8FMeO5ptqwxkz
/RY8P0Lnc92Do9CuoESMECoaW9tXDDI19DshFxR30Oivt7t4VxzZOKiSVVdBVlGL
J1bRzPSMJBr9CWEbvOG3Z8T6VFItKE8xEdF1aJg4Rsgjr+34oqNbqsZ2JUO550F7
Y39wUdq28f8iscILtj03/Pnb+eXNmKlI8RE7Zj7f9QbL3b5KupY5NipxFm0Yl9h4
dsHpevkTiVbj0gN/WpBHNMRkhO7tFQSnesjlxVTVixlhgnRdfI55N+jk5BBwUQJ9
42AwT9gGkPLelnqGz3/3EL4exDG2nLMkyGkA8yg5PY3Sfs8/KT9VCHwcBAHdPP/m
zi2WFHrvw8Qqklo1bIUoPO08xPT3YSTVSfz2a+ukhscW6i+/3C4Fk71LH/Utp8aK
wp6uq3DFCxXdoyt7SVFjPSgizSKecGQxAmYOCmRIEdbyqVSvvPctopuHTQsemFcm
bG87OmjlWzCdJs2zXj8ascee+ipfl7R+26OIdlHSZW8hMx/tvfi4246rtdSNo0tG
8hceIp1+vSL6vRBX1zUck8Z4ogEgOd67hLPNrol4A+b1ZAui2dG8RyQWpdCkGaQF
vuThMYFZQggfRqyg6ug5vlYG87KQlK89AKKxJp9bXIMvLhi9HmFEyw5VFtP5luph
TNSEf1I6IVFnVuOz+9avR7RKB3gkByjCy3/C9vgXCPqC6Jl+dTaFlsourNXlsbXK
XLSul4ShZ2YfyFFxn4ya5STRO9vQxth1g7TlV5bpvy4Smm4Hlm9JVDotZT5rGAgh
lU01jEBNO3NzhIa+GjdlAF1c7XFiwjqehu3bBc71kpjJQGxk/NLlWYlOL9KCdg7G
4vUKDQ7JCHuSZWLdMjlOVkfPPc36aaxBZ3kS2WqzulSfq2Y2yYvwMdT4Tz0wqA+U
y0L7t7ZVgFp3KVTEL6/BR+AQVd2aHwDp/eWoH+f4s4NH9OOldcZbilvErlUbHO44
p8qygt1IuIH1gQDFpTSjc5a6KQ507KkXNF+wK/8wedNbrTZVdRuQeXOfRVXyp+6o
zYFisaKy4OGrsaG6J1qQG+7k2G9pVC410/VSCRXVXZr/c8cpvgj+ffCfO9gVxXAu
zho9hNQZmbVk/iKjlIws0BVTYpGCY1Z5mEUdoI4Dp/LTwt3k09l9MAVF+j//+Xsf
ZHN1JK5cibBWBGI8+j5kPu0fZmZDVOxh2xb99i3s1eKREg68dWAFU3QVtwhJpsjT
PGnYSw3HYiOTGGF8PwYBQjXNgw1SOPUfJ4ZAxzK75nCVM7swZXJbxgKooW3WVurw
BBayFhwCRrBRqgfGQG1iE/651itgxUvFnbPzxwQIG+GFmFUAuJ3ZGwCwz+uL73JF
ViduEQodgE1gIohirHPL7KfU/vDPIuI56prWGR+XebpNfxd95gMO2qagyB5AyXUT
Y1ahXT+KlHDpUqCMoedUii+y021mOldAPDApPiF4hsWCbDLG6FYyZyPFNCH1NDL8
lzwkYAMbu3BY6HArgrMfQ14+xLOCFtvbO41OWO0Pms1ymHR2S0Bl29RyIwYzFk8E
T2++Ip3zt7u60BAFGg6NE5EPA2qxHFcyn+Rrnm4YM6exgeWuoEJeaOoQSeRhvNF0
oFwLxrmPgJkB59s6U9oW0tR5wQz8ZsgM1TvTjgEDH4qs3U+EV4B/DQzRpQ3inilR
NHg5dCyWRtMphccOqZZynYHl/KYSPx2h4aBAq5mxsS+eH99mFrayivSPWFa/piUu
kNYjc3WB7wjfRlAzoq5PmVZh89mduhnHcuprJaQkhUq6o1nQfDjvfCxQyiFVRR5z
Kq2xKRqLeyjNhGz5soLSqhoOe2pAkwYpqaT3N4x2M8XNsJT6BdSQqfnYwHf4JFJb
BqCWjW6cXAFs8mucIse+K09ha7OIYkdyxqftATY5XYousf3lE2w53HDh8UpA/n72
kRZRT4oiYJGvaloNqq0iWeQA0IRt2yhP0p/iGoxyOW5uIAB7nhHyz6uRUI1xVMsa
8ESEalr60Kpf6lBkj9xVvnWl66dKpGRzQQGZVu+VQjqi9ARJKMUzzj5PR6+Wz3Rg
r2BR7q0skMzUjZi+yj2ULI6YLJScYwQ7A9Ocj0Pvf5JUOnUcO16Af5fybGuxuFs7
QndayxDVkmgY6ZIDvl3cum3DBRHauxgVWl9agQ+f6W8AKeZms7amNmwllDqSP7Zm
8F81pcTbjndNkXEkPrfcnRbpDHpcrFus4uyxxJdyfeWcIS5pkQxC4ShWX7ad+q1v
gdyN3ST8rKazKzMMSyGEwuqiuu8X0J0OU2Ee/ccO+OoElnxjNJlSmij48J+483pM
/J8jPFAcVpc5IUrBgE+2GBRq7SYffvQgwJrjBiTEvuzbThJUh0J9rLnD4iSY/Jqh
h1i6a5aiyX9i7mkQCd05VsucgeWpsT4BVz0E+HLKUQKKFAhuxwIVJFGa+ae8QzOu
QucoxGVCL9p4RBFD6V4Lo/xWoT0GvrpEaeOgWg40MfNJg7duGFgxcjO/qvOsnTRT
ngiMtjjFsYM2WxaF47t98Rsfi3GhvEgiLn030AwJD5sll9JwX719hp8XBeD1EO1z
DLad1ju93a/diWqp4RViUQMAWJSx7KaDvigLNj0YmN/otDdlAcT1Y7vaVnSmQ0Lv
Qv5AUsWjFQv9x9UjBtD00tNhfvpbhQyHM+L+LIPUEoQE3CqiKuGGRGHnBAtziU3z
eyUCRG8rs5TtFfdtaIF8dkl06368RapkW2vIOjZP5/iCXxhQwDJcXJVWBwuuZ43/
XI/JGFixzHascW1CQZRDEunduyiSXLarcifmYP+CD300mRkxUYJYR87Yv84Mhs94
z1c6/BtO9NvLo6OzoqzDoh5Mc3u3WToN9FPxhWb4wJSs8/33CEatN81nTKm78o2P
8lBXBOvSWjdTxtKe1hz8qxmtRMbpBMjRhKcE9rwg3LedEjVi+t2G8PzaD2IUMJD+
1WySmyKWIQCXv/Iy0EZoDsuQ0AYodlaum3rAiZQ8nf19n/7DrcXVD6s8XwSZe0e4
ofaw37GOPpM1FNmv1S196BsoPOUk/bo8MAU9SLAVFE1sgleQJhpDxflfZmRdtwaS
+eb6OvkU720N5hufc9lLYFdPvgfclGpuJYI3IBQlJSkvoCgYg01V0Drpq6DLOk8H
Sl9xudWB1KcVNVFRUWTqbD3xdORUuEVIiZrfOkSeky3TVNJa+En2oESi4dCCeqov
jwit5LUPZMOkcw2BqWGDn76a9F8qbRrD/bppKeZtjn/oX75EXk0Okes8sN88O5wc
4OjMDanBGREJJMoSS6ROaWVNh6bcq1z9c2gvQHjauW0J5tghiWnEFduj/2aav4ro
CZf+mgXz9gV+NLmMnbvXgOcKnaeLr4bBE+6N7yBz0MfTEx0SOy50xybWO7+MtrPi
3FDqbvjJzVSP/hwu4F2gK8aeB4l/YvZliQ6OmDN/R2wOzDaDiMOcMvrBbLXwa8fX
HjdPqTopqjBgwVj0RJLQ6LqYgt59JVRlwtRbMQe9wc87uwKphIDfz8QoonwNyCux
EJ+L+ibMvIo1oUWkPG3Yd9ICPW8bRB7AgavB8qwvUTGQ+4kami7VfN7bJySwL8N3
iLWS++UOA3Z8NF3+D4wwYGBLGuSxj0ij0aV6YELqiu8SYww9nDFcYI/F7YryaUaE
UVdifQtpXJejJQVotFzP8GBMXK9FrE5BBvWk9qIVQZaqakgYUmrdaR/Uo69oDAiF
t29Blkv7vWYWtEa6mt4xtB7fxjwwnivFKwRBlNF07o8nXe0RwWaonm1H1MFF7B6+
WHlKG7eg4tnCLcVVK1B7VSZXuHwmGFqz/qxFM3LvdX3+gHPXm2XeEBjyrh3VtUZe
ZBPY9N9Jcjr2rQ2QmuWbdFbsYdiKHvkhUdsmdaMeC4LawEo3FbTuIFbqixaSL78b
MeQejo1aqdDTcUv0S3SxaczuNR0V0snc22XaQfNLDQ/p9N6PfMmP2+H/NAHbGgZi
3aAUz1ofHRnhdW3AzzTEKWkgWCs7JBa62yd2BiH8bzqENtKx7E93M2AbvzE1N8V1
P4Y2d0XkNZXD5hBaiHhomXiiaJ2MxOZov43ARCFTmu8QuS4StUYTzk19GE8PsQxv
lAlA2EHSVmHuWgTewLju1uwfvtI4mbdJQdIOCUyjNBZm86XrPZXyzyO3zTLG1Grm
cr+hGuj+KELLJHYZKpJd04oH8w71hJ3FN0Ty6zziSO7Wuhd6A4a6vEJRYe/NMENG
mqiXTNHeYdHyLr+zVPpYVtpe4PYCgQVvAiR58+jn9KVEt5KRWeP8R76N+xjnK/Nk
mQjvvLtl12lw2nVa4e1u2EBCljUymf0Gm0YfFqpsSyR8Dpx07Uq3Quqg+E6Q+t7q
sVvNuwmO15g0Za1B6t6mA0Lgl57+/WfigK4UwnZlNdprwO767ThYsQ1y5qTZzPhd
8bORjbih1I0jawtNl6ffaYgv4ZQRW8hq7EHD/aI3bav2/qgI1BVGiFOKi5KLb3Dl
w1rO/NzveW+ZamQv10LbOMdFHSOCFdn0mJjYmyQVu47OUTVfeeXj6CDJGNrC0B0W
GRPzxEvgYGce3mkJUhFTUQn0gzbbU0VjOW7e9wUjnBq07ETLbLuGF0PgOZ4SdV0P
UBIxRNtipPGYAJqgDCIo/t+KhgGhUakYiwitp8UqTWaum6guL3XNcOF270jlmNad
yvM2PoabRrMh8EgY61qVm5a+YzwMd8I93auCeDzL0wrW0xxfqfc6Cu5eiLdPFpK4
DU1t5OxtzbCkZLrh6nx7LEb9qQCZYHaIt2gjxId+gnQ2aBydy7GdRM+T1QknA+xI
5SnWt1F6TjT5w+E/ureWC+O6PYBfb/QQoJlHqoDq5eTpblZKEsHNtrPZdOeOOlZ2
XIAo3bYyW3eUVDFGHNmE/QR4A84LTWZC6pq6Ow3gOsUHqHqeVuy+xDspWYPuMZY4
kF323fuVsmdoUtyOj64xF7Qfv2BJ4Hvs7lFyCowQZs43OhlqZ/DL+qk6EpWT49W4
du9NuFII3sPMszqRHAsYdCfSj758h/vz9+mwnSGMmtATWD6VQo22oCbT7a415O2Z
IKxPKkBR6b7tq3oFq6YGR772DWSW1N4kArLXQt7qtIOWVP6gOmAXaFAEb5PR4VbA
BhHCuTOhqJHd62/QvsAXJATvwitNz4s1dC3dtKcJCZVZdzvx2mq8Znc5PAq+j8Fv
FmZs7vhuq/WorLwrIvmq6psYhz3N2/UAU/j7BON9heeNTDDgTpz9wI4dIYTPo08q
ZW/DEtIM4ntw5JeUp7hJIt/S9AKcXf4W7bQqDgfL92wreiSo1mzHqXunshAYORIx
57zPPBqSQhEjHbVVtj3R97fNkwYbmw1iTLdqLNJrT2awmBP8h7zUFg9VwWRB/20Y
jTOoGLnUQWrHJrekgbH2zJxv7rdccRLHHOXEijic0ATIfgtBaDjaY/KM1fVumXeA
oNvVzc7ibKeIQ3p2X97mVtYPlJoZl6414vNqMK/vVB+ffHUQPDVbQGwIUSTUpFri
3f7h4TPGQarCgDg5vcMcvQVTpnXj06wudbaNRpn79FLCQuJbsKXdKWfB9yGhFtTA
gG0SKlRwb/xiW8vZ5W6plweFnYOAXIj/vdvG2Psom94DZhCS48bRH48t/mLqiNQW
vU4tOLlBLxn/Vjaw4rZPrcaioia5fYmF9YWe1g2zOkc4JaotLBV/D+VW3d61FpLX
OTs5Rv8hiKvnd6SVTndgEQ/pfHDxZljNe3plYfkWUnRYiauKumyT8aQ7QxeFikHs
qM4iCVOMphPtKMrx42hzy2AmbWmAayeqCRwiTlk+Oa37+K0ZgJ1p3GuWyRZdooBh
mQQ2ZEWvr0hPA6U31mwNb8vIDnMDXcI9OWl1UhicRiz8vFkcsgn3xDpZ8G7MLQSJ
DTVGJRAPHU2KoXj4CJmxaej9/1MxyKp4YJTy9qR/e/gwHb5vtUTl6HrbjVHGjplr
tsASENighTmL18LZKXJHQDNifENrZpdKvzcbOLq44ErFK2haG+xMJ9FnxhEuOFBo
jcV7SjZoWOlg5DZ2jpvVnCM13dLjoZdMcqnDWXt5Sq4iAW4Q5wv2pzL5ugpt6Vnb
CktiWyerfF9K1CUjct+/DMHFlBafVYAM+/i+hNIQky5JNCxN8W8gxD2jk05FjrUI
1eiRJDJy/Z8/rc9cEDdHHBRDaneSPenPvMnyc0SPxDehffcMQk8O8GnMy29m9WAQ
dFu7zcfkTBfWZBjUCkFGCqJWkkqTrBK/lu77NYE4pYh1rDvNb/qoARN1fJJNRdjY
rxZXETiYwJQRqxWiXkliVesaJ6haLAbI1OoIwXRDxcp5C/H0VrFtNY/P0qloILbX
Z8kK8QDXWMiA4GVY7M5Cl1UKR98bYk35SnGtdRc6ynQfgXnco0Kajug+5w7EPCY8
7LpzfTUK3Dtb8JMbhkqONhTGfYVvz6aqIJ6yFybz9cHQ7nku+f9QLvu9hKt2hXdv
kbiRQPdFzgn0OPZRv8Qe4dYR9ZJZeu2u23MGmcmyFc+JVgtmZQi3hk8/jezKQqW3
oMyO2lwaR4Ci9C4AAge852hQU2kPmuBc307n8i2k8S6XpGPVVJw2HOqe1DoxEQ8Q
F/2xyOxBCiQ9G+wwcLU8JiBJiu/ATfAYGZ366NrwZXpSIOU2wjQheZTOfsosHmgY
u4v8KPz7j7sg8y0N8+X2hlkq85mwMtkmBRkKJg7cHIYSOGjYIS4pUw+2D2bIDDD1
AAz7WhG5FRfW/8j9CjjL9Tn2LE/VH4zMMRsNKZtlozr6Wpxt88fB83L22RdVFBOc
1Cykauftdh3BL0cE6oFF+Y9B8U2OpC9bdT1nJj9l+63COswQ8G2wntYPVmre3yZ0
G84xMlAovKK/ibpFwmNZ3ZwAF44Ila9PnxRMtgvF0/f6Ff33EggRLfW55Eaez/F8
/Ckg5Bfafb48H+cWpOhis3y62tembQk4/FgQfp6QRUi3SVLgCOoNjMEqT5swkXTe
74fAsggS+dMckB269/27wOOmo95A/EXljiINN3jVECnXdG5tsWhgGWg8zqQeeS+9
F0ts4Hons9Qx3JRXoXu/pQvqsUbsGDxOvQUiI0k8ntVJyllmu8tz4bP7llNSvDLF
hAvuNd1FwBibie27rKM6E8bPGcgtvTsCYtSh6dJhBhtID1JbvtVHFOYXrm2imeWo
glMriQwRAcFhffcmmdXBG0fHdZbj0vv4jwHA9Lv7HHL4JHdWUPQ+eU+XMJKZuyoV
jgYsiicLB2jXVwbhoZ0l8mChHCG0FSCdmpJhDX5T33PHDnL+ovIlNyx0wRXip91G
dqB/rU3uDbt4pR5751b0299gne7hR2IJCIHafcABlfk78EyRVN433DywcZEfE+qa
TbWH83Kqd1XHxNj98Uh6qOux0UANd1hMk7dAeRdPo+LPZvzWEaGzzYAtOHT0fDa4
orGbrQxYF2jyiDulwrpYRlhwmtfStJ/M/zRx6ktQxVX90lBM6MruDYvuktZP8sGU
LI6bir+cO6dxRm6JjmCsQnWSRc1DXFtg1v4P4Z9dvQCVLP1r3F37yVBBEgtducs3
Mh8K6gzX0DsfLL5mmPG8XN7Ap0wUqkDzSIBHxCp8ACAgdgR02XEAwQNN4UpTxTrq
Z7yD8DwFxm5A0Hw3mupyqD8AcWbFKQIoW4oWGdM2LFV0iGNo0Z3Phi/k/E2ny1jD
ewezwyb8d575Vply6JDJdssOXj9r1/WWgljkA4DVQ1iiGckGbdfDpjCJOaBUW1dA
WNPjPxvZxm9w4bNeARUPu+G5umrtF0Av5ups0wT18dvujN1g/Oe4B/4lnou4uqyY
pORJIBD8/4hEb6iV+Vhdb5wcRZw+vwDC9dLmxIqbFaK5j6EEMdz5nj0Rh/seWUSU
dziZgJER2HjCovOeaV119jZ4ExWg870iRhq+J9z+flIbWXoXQiRYoMWGa75HGOcZ
qQD4ew10e69KLIsyajXZcoq3ibh9Af2H/T67VLxAdycY485AARCya3cO5IEIRZuv
xlc5/EXnCZCVO5LpmF8mDNA2czGlA3qnGHDbW8lzAPV5v1HDuGWqBty7VLBLGk2Z
SGsQYGEO0eaCTIw08Tbz82kNEyUhNCl4KonuSyLhtGxqZyvDPBGvbAdG0S6bi5IL
9yrlimpCrxd7eRFrMU369AIOF7sKFKMvcj3wEKOaiINoNr3L8sQK33Eq9Uttcc6t
x+jlfHC8UZxjqT7meI25ryRIEBORlydJoIfRBeLEZVCqltBU/+4qdp+8+Kq5zwR4
E77tZ5JuuZqhMPweVB5OHlaCG8XA/V29qB8qBcDTRT5mWS41+5OsSi7Uy2LE7qrI
tJSTH8L9nZ8oOj2I/5KLuPvBPKh51cTF2W2NwBlv7jNfBGThn9b2uhDyB0u7/3Ty
bRTHU+p1dN4/qubbxr6TaPoICT2cwaUenlQim9AMqtdjDubhuiESsgAGhJK67c75
DyHn938yxru/u7q31SmLK7SM4AD7s7upvTOBEVvA4irWXDSnRMjYkU+bVXGZUMDl
Lqf/XTDhAKjQZ9CNWxei20crjf3Qfa4M1X4UN98qZD0PFZ/h6UBXVGaHsTFPbN8H
Z19jtk9bmiDG5V0A9f1HAXSUAaaeOV5HVPlnZ1lNUZDnRH0C0r9iP4+ezZ065FD6
oc7o04MKDfkCuGuRDA5Sf97q0Ffeap6IYaRSS4VGs5PNbWhfVNh0YqRFmFVpCRLs
x4eMbj+rq9priszO36iv4dZ7TzMRpK3OWnhnCJoKtaX0mynWtqt5MwePk1UoQBDs
6R2WZsWzKJcYY3TBwX9Rt4M91Eq1JwbQ4qCNmjSbH097EK4yRLIUavhnXjyuo1Yo
SjgJeu2fo9ku+zIKRK2QSU4V+fCqulDByeLoMv3wUdGcUza4TXAkq1iJKgPu9+6H
lJuePcslwBOHoEHdebiY/+Pi/acr1x3aKQM7EgLwpjUmtQJ6aXoDBP9VvE9vPQY+
jljqFcsT3zWO+yFHJyFrEsrBcpIO7r0y9rQ7Flisfnvk+ZPRmfgNmVRMZhoGhkaA
GV0I1Fb/+6V4heBc6WpE9OxhYqaU5RE7qN0WDV1mHoGKKw8GY2sobvAMkMaFW1RK
WUrahiwlsqXofyfzA5LNFb4xsUhbt+wC/fTIqTEPPuBK7mBAXCiQ+lRwDiQnv6n9
0ajx8LyAS8wV2UW5EJ6l/Cs4vNV90/GezO5pjIkRDcJFPqyIwmuYpn/sIv+ToCQm
V1JZ/gjuuSSNEdbSw6YFOyKQEFi5wa1OvdjXj3rPI/51mDx7R6Jw2HXNPvy6Zq/y
EsYRaVFs48yfZT0UttaFSwAJRfpPXZmoPeib+o8ir0l0uffwlzppkII2IqeESmQy
Xi5L+8Tq/fsnvI5e6dnT/OHOVddNd6GuCcOArkLrre1T59dR8vmwXsdmtZMEYt4y
Pa6D2KKlk89VGunw7YqvrJMjaee8wP3Kho8NcrZiuvYk3ZQCe3sqexyh5L0mhe8f
2Q7tLTTPRS+eE+dTe+XDyt2wTGQVs3RIElTi29ztbhX9GfLHgg8fAwvWYwEgyIxM
SJ44fBBu6ZW/vkLK9GN5qU47FFmx4RoBEhYFcev1FwDJlyh6eW4AAiUJP6vcq/uL
SIjkKM3EeO4IU7Zd1M7gezfH2yMLfA0P0zirE7Z0nTzAi2qt3O24tMT0QkqupgXq
F14Dc/kECPdh1Ysa7mUHIX8XzS0A0M6Gsi7hieao165YdTahxLCP7Fpyk+8E8WxA
KJ9yMZSc7NQnEgNjSvHUYQM1gierwDbAWDAQ8jdVC/8q+Hm76PotOwPpb+vohLfg
5ZmZAw89qoOMqiy+qdFbcX3XTXv7zqJuNqO9p8Fvb7UGZN3Im9Idl5abxeSC4No8
9bZUz8UWRf/qs8GYg3ULfwcvUMxD2+Zs8wVAugc6x0awKv0dT6k53j1uHRgo0xKx
JvBrX8LdACK/IQaUJZZ6sCicNwHSIHmNL0tLGm37KZIhee7M7PlYclHHdfH6vTjG
5Ondh84MreoFu9IQ5qweSySceirBBtNCR8JFlw6NSuyjOeK3Afh79/pFA5Eiloxv
hiGD1oCIuw9CwxCWknqdHVe62N5TNzuk2xu0YDvMwNzjFsPi2muDlj56Liq7xjxt
q2zyfgEhzCUDJSmGjvjKnrXk8KW9ULWuzmqdB39ipmXH0URKjJd5xnrYPW4SSrrH
KVGKnZLpFF18PhuJMs66l9KFD6+S421Le/8aqJIY/bEMUBh90WUUXBKSP7hOn+Mx
L20LpRGMvLMz05Xkjez8Rsaul0urvHDQvpgu7IX8Z81kodfjYNvhNPcCc7wAN8mv
KOti/goZuk3QNSXM2tuonE9PS5dROAldzsJJyKMLg+NZ7Ls/cRzoI/EOLMr0Vpfc
+z//PrkE01NIt6jHr6bEOQ1QsYIlqTFUL1oaDYcyWJP4Yj2OJLSL6lghCezNHIvi
TbwY4zfOsCMitXbUl/mg4qXlBCs90JqAcctFkixpWuv2/RkW52YQMMOfJg1Fq6lw
f5WhwVAvaGCdQacGGkkftlmtSG/F6sUP1k0q7EcPXQbeBEJPmpMqKkT89M0zhz3X
XOaTAzUKGgT/BcCYUu6Q2n3C2NrZDD/jZNIzzPEYAtZNUDDZZG3wKdQP8Ymy7fP3
Cyccl9PZ22o2+3I/4M+THwICeWo/zlNZOkrfpwjEDTniuEoqStYMzCV2Pm+lRIgH
C/Chrhxr2KACHx1whu/CBF+RuBZ64vqHXLzzfs5TX8DRxo2dBOVuWHOpO3u6NCUt
oicgz+Ab2HrwwV3VJFyKWxf30IilvTzNT6DHUyPEMMdBvATaWxkqAtsKj5kXGDYE
9IU7aBjjAH9y1IATKvw697u2+goB09KgiJpANjE9J6/Zv9O/7H5peuNk7Y/+cv2e
tbnxnv6S/eYYbmfLB/r/SPmub4gjObndUpKrUMCOwflxlZtcKF/i5n5el6NQ09VQ
EdHX4YtK/XhcX4JIk3Vp/RJUj+ScjW4oNiktPyLurHS7bHC4wqLOZ1OUt7XnqUKX
aZyhZxHGk59q0+5zEmvrZh0ON2pPMYJV1sXBPuDHM+FdJLnr4gGP6K6fxuxljTUW
ovN8FZMyli8j4LHHAIu+/LvA8Crx1oBFvzJtB2hQrYM5gDlgN9hLxhcjDojMFoMZ
PJy/P2ebyJzCvAnt57pP5A+XIiAdZnzuYtJ8OqRmsWaAAE+gVpFwkUmslvazR0IJ
elAwedIkIlXFPfhzEAj1ZVx3+DXihWL11n5ZqKfQjuEBNrwPfjSP2+HpjIqOjYcX
j20tUKCyowrJ5ni7iXRtVmFZesd1/0TYSolb0YXfvX7NsZHvSD11t5JZSHv3BRi2
4nbBabHfj3RqiHVOhf7AHZXcrKijH8Viz1oeG9Yhl21lJjbcDct1EcMmss51nbu1
nuyLk0vyortZuUG4bgcbKNJL2TXRZNBLy2JEe96pEY7bsHh7mtXI7Q44v6EiPg3i
ZXjPyJKyAbJmbAObN1MGzS+sIHoxuYchMLtdL/ageWucnjN0JsKSvs0Jm8wPEitD
mcqZUX+q1dGGPkiSXbBjDxnuPHrG4ltXmQFA8rDhwKcddjGYkit12SjLqc2Yp8R/
u5BLeeto9nCpA6BcEJEcNULbFiFWu1p5yR41ETJkz7EmlnT/3OEXwmw7lJiN/WXo
lI1WdjwXOQxvB10lQhu4pS9VCEllvDpdPZJTxnK9LYHiOghDq7dSTCChQjesI4BK
7rqabDLSK4PCUF+QJ38+yKdjCS0g6H5pW9sHqxENs+jEjPrR7Zh/yYEBixK+WnoW
tvPiwCRsPihLSMvypdY5Fjk2QdxBza2KPxZY+/xVRoItrO/yJNUSpxl0mj1hKvkq
J72FjBdGtR5WrvuY5u+AO3v41YW77UKWOloBklb6ZbCflWJmdXt1HGxeMUGDI2jB
52A9M9T1wUF6lCzRQYvEfFFlLG1csfeHK6lOFdr+Op0AvcL90i04eQkq/xGjZ0eu
ObOO/jceOszwa+2ECoSMtsZh5idYnIjNKpZ9CKZ/NFA7hhcIZu7Lz24MSAx66NCq
ugKRXiBKje+/PqvMX71UBaaJzgXiJORE4btcNqVjX1HXIAodLJ2QudP4B1jpoBV6
BEhzSkQWUTFzj0P0vsUOVf6T/sHBD0ReWp5IRPoVco9F/IdJNV7RedsyMtIBEC7j
GQfKGRce+58DGeI4xo+hhFmnH5wZfFNAWi3EP9VShvKkaG5iV1wb5o21ndAc+IuD
TM6jI52osf1Fd+kAS1veI4EDd2f/UbQ18tZPIgxUZ4icxgaElwKnuZ7A3IhPdtmG
GtS8JuKytqSbml/Fdx8l8mQ+qCbfH4A1mMjep7w4EqzsXw8usc1kXYMZF1Z4iGpQ
6DJuWf8jm9hfv0b3iTiC64cZMpLge8LHolPqQhCPjBHFPuK50vQYZKtg9O0Fp7SH
PluLHWDQpmVB5Osd8zK5zSTJmmJeCfO1Bqb2sUJnix8h3ha+YmsVwrbwiMyCpAgE
oI8s9BcSko4aDLgO+lXEk5IJGOiEKrRG+hFcoYp4jpyGzREryte6tn7/RCT3tV6V
5zMM3Akut3J+QIXHhx9qdWkEkokvOQpcHilmxRsRJZdIoGCUPxBHqxmgaxE1xHrI
zX08UoQAGbH31cW8MeBlF0RrkcZtCpzGmMT7v+l978WrJbaQoTeyF0bli4b+GjeV
Tb7rblMQjqNVWUo/M7kjpwgPZx8QlnLWNzd9VaLWK1nJQB6oFl0EQlvscF308On3
Fxwte3QsNcw0CPQHkJ4+5AZsFjP4k5VZazQ/AEtAkAgIu4T1vGaxTy/sbEoHJxFv
mDWRm654LBUVwiDtAG0sLImwYey8Auv+PB314BmC0vO0W5DVVPDRMXHWg8+iQyVQ
5Hx2dgSZ2aMUPYtHG+5uTJAnG/xgbVbWONZsCgX73Cm4LJkNvP5e9g7H+1G1niJm
jmsZeXvL8gSDiP7GXiZPoZQw3Kza03b/kSjSMMNK93rS5ahRE8nSrFVEKLJFMlNU
iHrsne92afj90NYYklV9aZOYX8rtVPMi9aV9SjaR8vPoVZVcXfZTkt+mQkZMvmhj
0A9HFnHgakPSVcSXzwfuUoV/hEbgz1lBi5kb9I4fGCL/v5Ec5B9aTUchjYMeinTU
SC5PqDDU+LcsIZIu6XdwGC7RAxAr7QueBmHulYY9twOUUYXkluo2lvp/1DghpOwS
RAAnfAoD1AMMpOJbAYS7KmnXuZsgZWVYKU+2X3ID/o3GvAWWcuiQ6qS+xB5omz+D
7S/Q1B59nMPk3d6AS+NqY6SIu5L/GWwROQOKjHl8frIAPh/HvWUmXp8MGw8bSrmn
iFJlUYaWul+rEDjrSbmXxZ9+TlKYO4+oPADRBxHNEwfTEFrcyEBCnfW9IbA0u5LT
H3mKbrZh6xaOxL8FdhLnitxbUD3FzBNSRlRGb3XIOt6rfh3aHAeKMVY/ynDyLd0F
bth23XueYkefOl3X/NfcoQhMxDC012En4hKZmTp7zQFFE/xoa63Ray8BF3tqUMdr
ByiHm1Vqnn4Ps253P6R7z/CNHpOjvkLL2u7SfqLFREcPyxp2iissE882fFjAFDnY
pLi9SiftzXtTkOlMcllhhrvakYM63mnHsreKc6DHj7Q3EaDZ+vlg8U45Zt0v3+4I
OynZQfPQxZoLheP5lNrExZBm9jkrRmSESrOMyMvrXuSiA6bO3WH84p2F8EgEijVf
i/y2Bkb1dVKpaPRnmKaOdku0zmKJ0hUZsUy3z3TfOMmlyWZYuoqo4AzIdQNS270r
foVAxHmPOeuEtYvpCQMYgJm2f8idYUiln7bZO/2vuKueQ2jHJYmM1Vd9gqLOhrOD
LDxfkOxHruRqogLDV5fdSTWdj34iVIiMLP4mxQ7TRJMGnOjtnIZaoQ1Ghtoo9A9t
LreL8J5h58tCspz6J/sar0qWNTz9bpElF33N3q8xgtESFxzvcV56FjO8xN84C4WD
DfOmX83TWuBNIqKUrnAXRypdGkHVMZVsBSqLPPDdXpqLVpzssJh3LaE2CriQZ3hP
BXEemfq0o+gCd/GKUNSu+dI0KccbcDDA1ajQxCKDPCuNvEh/wF5HXqPMNASM2RU2
KOQ0P3bbl7fL+7yQwW+x7ayX8NOMqTOvpf0xLhOUdDRhJVcVq2TMNchZpkAe+u7I
04PxASNoVJLGd4V7uHTRKsyBU7WKwEN1qA2FqP1nGCr71jZvtRDN21wpso+UUoGi
owMBVGrWIFWO5McNMGTYjHVHsBTudPy/lybnWW235xN21Ors4rZL96SYE87e1pHM
1azdNY9yetj72AzWLACFxU03XBMvXzcoTBEFFmWTp2+jbC4YUZEI0mfATQnri6uz
5ujlFeBNLhmKpCf7Jx/oXlvU6+TGIyofPGie0WvYrnP57aWVv819gBwlEdjnpNRf
8P6VBWhvWqXGMhehNL+Dvppxnvef+l2sGCBhbi7GXsQzz5d5Z6MLPBOs37KjbcrD
a+eyIW7IPYHcccdz4FkJyxwSbyl5JXyXpktu0Sm49ho2fM8wYnfToybzdTk+APsl
VGkDY+49s6cR7exEXB7WBKt8TQL63tN7JmtkybYLWbb7VDQ797e2Q5JpW2/qDa5s
zHZhGBCuj+/uEluDZuH68KZ3AF6zFF2t5dwbiItAdzDjJ+CHKXctr7Zcpw3p5v5P
hkM23eKuu0ceuwGdhECZTz8+s6DH08s42ZQhlJLxuwqdVu35IBdMlQk1vXwn3pSD
dixQTccapJpi8KHxf9tjgFRLlHJRGmrL1kWvXAKnfeW4AiGJhNXFqaeaZRMbs1bb
fDEFdF/xNZpaqosWehZPOS0V0kPkMep43T9tRDQOQLgU80OU1M1J3Fl41aXf6Hz1
HUzcnYvL00gh5vQptwFe2Jjdv5Ew6l/DZiHKh7R12JQ5RVIQzS5qSi7kuckHq1bp
kebM+XaAydm3m07u5tjyCqKI1HeQXuleW+sF8HaQaOUWwO+DWfS02QTKgfAnxtQy
JyAThDa64tvKlPdGVjGCk6ugzrXGX7G6xLWnoDHmsIX+yiwzFdU4V+J0iaNLTAx1
yYvSZdrDfDAgSV1caCC1OKZRPnA4mDV3uR9FV3+KQQOYom0wk/1s0zMtlB9LeS3A
UrtZlHAkky6U33/6Ql5rXox9nkdOidRxsWE73VWr0pE+ZL793ZLNMTcTPThj9rR8
TYRNnE5+RnVz8XBGNDgFnyeVxwfTRPR/y7yzne2Mc7q86CEyiiwP1SPq5yjnPAjx
V5UB6xuIB0nFJ3QD/cWVYOG/+ap/MRQnFoINTNIdOHg79L1isgxbeQNwobYNxfZf
SqP3Zzdev1jVxU/Q4Mdb4GRhM+l9RNuMRglDMLppNoAMr1hcUuhKoPBB7sLNI/YU
ojexm3T3ak0goAxqyALQ/yH7x80WygeR2nQdEBPJnsILXfjNA+Rq6a/cSjrsc4wf
6dGbQfP0VM9DCFk+tncSFuy+5PGqFeSWPAn0PJ+77W8COQBa37CW1GiLR8ewia/Z
HeRnRrT1qMbjnZzCwgA3NhgN6fjowbW3lnrk2zY8So92oMioAIwGQMUvidHek3t1
cVDStP8vD60+01JvkxOlYqaDBpP7qQ0k0dSYMDY8KrnJV8HA/Ts5O6aAn2Esa57X
azB3CJx6I3R0ip/4YqXqMtVEbfxSTfhfokQMQTuQAySFoMr7hUURHFeowk548JUM
VqR95LAGxsA/gmhFjQ5kcxM5tJYXPocS3zZHjjbUmrBkK4l75IU2bwdJnA0ADnnh
FwGsA5P2p30SbMrfHhnhUqABPj2BfGZf9gG9rp9Sp2NgeKOUX7fyY81eYeYH6bkk
1Avv/ik1Dy0wdV7+EYsCYvISHm12mxRfjIXh51+RU7P4nL9PAidMgH6F1RzRkQn+
PYDGBolGwcSGWd6pUnrhxlscAPCwIj5Q4fkVSYw/FXbZc8P7wUmuWmy0LraCCJan
VynNfMjNJ0ZD2TUFm2uquZtSCUQh3e2CiLfJFWvEYSf44dTeGEmL9AjtB14zV9hY
x7sedCIlnL3o6EbOjTa1JAQL3pwF63AdcpJOXrpRntYqiss+PnZGgvOXvD/q6EvG
Cyk4XIPbA8HR5cTzYi/KkU6zwK7XwTbOY7aosaK9bXUV0+qYOpBkLm4FGzw6g5Z3
jKlI3trrI9ZGFAWmX+EHyfG4k+nsUbKLu7Y08+TzQdGrKypaLBLdMAuALTKZ5VcE
E6hD7oI8UMO32uTBiR+94naAf4eXHQ+WUBEZw1WF/TBUFfePVfaoVJa2LWukY1NY
03ehi7n5Ae9t0E9c7mVG7DB46r/DQEn39HOV6gycFuNHbPn4J2MwKQWtKgQ1DPoj
oN6hs0MMsdaAmDHz3mRBBjCqXFKieY6xyHYfZhp7bL0l3hp9dvGP3Artc95idf3H
dZnyh76skrfFAViB7uW9ORpvNeFzOzN41FPpCerVRARdivD4HCNhu1J7W9FIt6pG
xDSh8pqRzVj0VjOACM2aaIECTJv8x8YK6+wcu8df6SlVK0ZDR40HF9wItYLzrxQw
zykHMjrxeeF05fs6Yhdzg7pEOAbNCBi812ZZ5lrgRVDYXk+1m82dvhKI6WrIA1xm
T8NZ4JSgPGi+glZoYr2+V8RCLZ8Beg+eWtI9UsjskKaFd+JjtuZW5wX7A3xrZ/VP
RsMOOZN17M9zvlqcc+qjqgAW+DwIhwVPzpVuyYg30o1W+fbdWZMZaMVYGDP8ZVbK
W6X68/U8R4xQ6te6iXc4/zdq5vaD0dZMg89pjl2I5OIdRnSG8lucIUAhaqOxXAeW
SsASosmJXo7TV5hvLqwR+DqaZ072cr46o2UrpjWhKoh+eGuBGXB1mLQ2jkvQzhlX
3Fiuo5+5tu8rHIcSMK6Q6dqQ4NN0q37EBI7jO3OSAI7ecNbDgbPN/qUaVJGc00el
HAvjET26wd16LCqbvNp+jX0XyzRz0wzeDzyL6jq2hKcYl8TOpq/im4gQixDvd9+m
ZQSEg4vBe66UrVwu/4xjvhIYHLFcgP5UfsdWX/07iEyxpWOACd4xpxs77AcKPSLb
7dFoaBwZI4e4V3hfKjAhZxjjTTokfQeUoR6sh8ATbpOOiZTABrOr3QI99vk6o+gJ
855kQpyUYs3IOsJYi8zPH9gVV41goJ8mb7PSJsDo8DUaD8kOq0MA65mPmfdYp8Vs
i+YEm+EbwZob3RGGil6AnB3PCSLDypeKUvxwHR5+LJW6P7biHmNgVTFVCM3fJWkn
dutaMx5Fz1XBpcgL4wCKGsWrKN5wL5PDSOes52pnpaluw4BvOXUV68KxXOAdyeCB
WPu3JJ53ufV3IWNSFNmAYQGLFHcT/kuQFOtg6u712TnWVq2DBZxkyzNhdUnQwZWX
3bA65hOKGMPe7wYLjHfc84KQVpWL67S/9QJEWQS7KnXYZ/5b+5DFJvhauo2vQSOy
KlP4RP0Bxmn2mwsydr3ToRVbZFByT9Xae6STJiym7F9USC8XChr6vGD9Ad1X3fX3
kgeCXiqmIZ3iRaBe0FQlMApHD4CuG2VeDiPkJ3RvbBhGGIxtI8xRsWYakU5VCVA+
nnq+7C3Cq3kvUyzlr9RllNTyips69r/5WpaR/P/8zjNcI8viHfG4NqXi9pAEZkrY
wIclh45MQA5lzx4inDXfslcdmJqNl7G077Qjg+rfhYNKtM6Y0eTlGHNfYhcqyFcl
TtLb6zUJH0zds+DThSLWAp3VwshsrZwqkutkpKL+tnRphVxLrK0V/HoEdwY2rtD+
++DUtRlABti352OixhJ4/rYnrnce3dDnZOvSbGxXmzSRWTKY3zSRFc/L+DyOFORC
FQ6k52goNsK/kRNJrUtdqW5ftYoadBtIyjbjDhOvgqUGNNb77G6hI2rZsULHuWrL
Rh652SnJ/7oI4NeE9ZtHYBVq1waVLJKDa+6svEaNMUXzlrS9YtRlaUE4WpmV6gNx
l0DOmueeqBLzjZ/mSnKVxKtu80Op6H20olKFXecIWvIFI01KuZh0imtmDxMJD1Ef
tZuApY2/FoL6j31x/Nd3YAmAqtLVyiHLLtHk4+URX1GNDPjeafEIQWlgkpJ9jghS
y/ak6FkxgN4S7ic5L/xARg1IWysejNI8qGYE9WVsmp/SjS5E4Ma/q2cidcG73F7P
zHE+PiM7ox8nxKcsu0Uv6UcmY7uw8F23BZBtBoRoStKU+YzShtvyXEstozs2xpIi
C5BWwcuiNhgXeNvUOzLh3eFmPeKcpsU4XAa9yVzCVDaV5OOtT1ShW8honhj9v8+q
NSuup7Q3CdLkoa2pZIOVWKSvBb5D9rSQ5JUfrC1BITHUjalpgVpetdpdjidHa6SR
NbkvI+Y+YJwh5PPGD3itaBofjoV263vzYZ8s5x2Qvi3i5OTwKNgWdDxh5nNRcZFF
02Ygk5ctgRQU/dHA49/+x90+ISvHvBj8GquPrCirkeooNyvtvEY8egA+zPRFqWwj
xvD5oqC28rj4poIlgsRDbNarc2HFVA6CtzCJgKuRnd2Dm3RgbwiTqBcC/WlnFVGM
QUahWeox1yNpDqLCncDMkyHEnUT0smdC6HlGXpqQEi68KqlNhYzGw/HRoMMHSok5
kI18TCtCaUasPL9m8DzV/aTKtQIJlw/0nCe2am6RiawkD/lnGBE1vQ0FbdggWnYg
diLuyA/BA2aro+d0u+RAgr4muLdsangpWV+bDNQYOxS+61rp0OxXTqOOQKqvxYqT
DLPXsVqRhfCcECeKGit1zhvhYerr+7EvpCmMZF/Yk7os/hdlVsIeKaSPsycqkZTO
g0GJIvI8QlxikUu/MkEynYxQQQfeLbMjU6ZI3n5j+y5fdxiQ9HQtWafJ6S6KnjsG
cZ/g29OzddkTAlbwFP4+65yKAF+E2cxx7h42rZy3uA/Pbjq8BOiDM3gdSEdWVZIC
KMcur3tXcYSjexDcobXwI5SH/7VRTlxRmCqM8Gfpkla/Tz6NhpRgD3tIdMPp/RWG
oIgafz8aM2INuMI17Nw3cxBHO2rwOtTiktWhtmEdlUfn/12FNJm5BJOi0+m/sVBZ
qBBUbLonTJOS1mmWSLtLyg28ui7bawWikkUUWSDFuYCkmL3OoIOEySBBPj9lZSzm
QR4GygPnTgBM8sOPkAZvSPKiCI+03t5v+26EZ9xt2hV0uoXrIlD30/wruZgpEvfY
curDjlld+Y6/S0/UyLnoZpbpD8CFsQOriZyuYzq8Ke33youDnVwTpYoI1dxoXXKT
lBOE3/dYxzx7iULkY5mR729N54p+dmridIrIva129Re4UVH9knNj/fEnGX8ZnEWm
Jin0yaNf5hanPThcxgLZZgmB9sh51ET95WOX+q1diEuUPTdRmixtk8efROfPbo8E
WBlzaPuzHkuGeeP5JJpnedR0kt9DtIRQG4qSRc/peuQnPJI08tLluxP0/7VGBgHo
+zw74Z5fV6DnOp2dcO9Qs4LsfFvdFTFIC02VHigoFzrG7feS+U2+deuf9OPjQYKP
1HUjyLJYx1n04YhrwGBw/aYoa9oeQ9L72WMJuJWtaBDIp2qfVB4IeJ06/UBgfRLP
oGUQ1J7bD2otBWmSlgQ2KUXpWdv2pZn7g72bEA4fZYVDgUhuLeAompHyJHhbAVY9
9rfihk6YvWrI4OJi5wwitbUNEhNnk/2ZHJYs6U1Wz0dbMi3S4YM9rOv2qNZLhosk
9Vn6vQbkZglpszYoP4NAB2lfh5YNKwKtJpIfvXtSInH/Q606c08OuaVz/1Tb+FCh
8RY/A9poqu+1eDGOUFQPUkFrS+tvt5E2BDmvTDpXzmjWHAtUfohEICrBqcFsUaWm
VBr5RcKMFprLCQTgLJoUzRsIyBZ0/qyrC2q/P8Y+x4adhOusuR9Z7HRXz6IbgpuS
u514wOluSnUO3YuLobQQtbMPh83jcGV8JUuNEIHIFbuhPSY2HeMyY2qURhWHftOr
bAMZ+3jQY3D8uj19sobn8MnioWdgcnrey567VbPaUG5YusiZ9LUWEj9VmgTQwQzn
Q3S/qUOJ7dyI0LBFuWaAPjHGne1Yw4fjtMMPA/Od+bqqi2Ro7zRJsD+kLpchxpvb
ozOZdY9qOtZZYs0imu6HjSB3BXzvv8xMlNNrJ7FoqwA6cVOwlvVA/MIR3exNcFTc
G5dJnhigGGpoRppOjz/dQ19Yewsuer5tC8/C3pLnffeG62TEeadiGlcKmkDR20/2
RVSNZZ/42ICzGh2HOt9WqJCdZqgMyXKIv4vuTG2o8lxrg7CWMOlQSRT4Da0v3RLR
rUrm8qJIkHIw/077qy1Jv1C3my2/3SVdk+VULwwMQvWwXYfhW60vFkgxeod9KmBK
YOQPormDtENdjcWTm47qhLWu6F013bTfqedtloQ1rCVv12P8Onf/A1Nj9eeIkwD4
teMzljteSrbN38vA5rHD/QDL+pd8Bem2lpV4JmJqhDPaW9464atv0r1uAcAs6tCa
Q3wi8PuHwNHF+5h60W7csyJM/PIdb0uHbaRfD8iPLhpH+axd9IJYp/dpufHqAkW8
yo9tVNCKD6BpQe5aTCgqCANNQuIc66jJG+YnYmg5gpBMqzM/fW6BQXF7DsYC96F/
XWRLziT9HnbPm3uTIEMj2xtQrfmLz/RLN+2E5pNm/wZu/s2AMCp23/GpnA8pqF5v
miBZ6SqAloz7FfGgYBlP4rcQ88jJe/TFFl3DDMOZKtih3CenvNSFBHoOm5kJ7uk9
7pQbxuRMWr0/byf79JmE16wAMCRZxJn97Ls3QRAK62muQfu3jDRpAvjHT5y2/2Rz
Q6w+w0eFYsURsgCOc1rh+so7ucDN2rAY4DYmO9Ln5xHW72LujZoGj8tOFVX0cdrl
yauyPzVMsA6HkpUY2Di0L3OSDm7J7xgYzyhxAF4cbP3n3nQNzRoLSEbzlgrquDyD
Xm580iALjs050GLDt60lZUYsNWztSOTYqpTF66x3IY7iEPdVjl12Qm/yZpbFuid0
yJk7xdCisEWR4SlMEUg1HamHkttv0QKGZZIZzFMZOcLjAWmh93MpxJfOb/Akcg2A
4XFPjIC9BC8kHgs0Tr6p/VFZpt6lcTRd9TU/zVBpoMko6OJc1UcXWWB0NZcBFFA7
MllrPLESt1i0EWB+D8s6kPxEwHipeJScPZe9tgZfqKQkvaAvXBfEibke40QAnEYh
FMSRRSpnsY24bXFcwqbDneCKpCSGC1PVcIH+SsB6mnIQcDkqOxgrOdWOhXZ8wzcx
6eUPZo1GUWs14GbN5mtgqIOxpoTwpHED+Va5AgCV+RkVydQICwskQxIH5gpuBUCF
HAw5V1HSEEVk0CQL1L5zQ2qxxxHN3Tu3frEAXdkBvmTYVGWnhxq19CJYRKX66t0L
mMqCSQDqQLAFHHEMooXteB3/HbfOgvdXUWbjdpi+BgL+IBxHTUViYhT4EEJWH0LF
O3NcsOkHXtL27pdp5ALSK6+GZwk23c/NBmLuRsbafurOP6X6hUUuE0HXWJQ39j1b
MMYpJL3afmFaD88bktmh2jgxcIKrf7gIRUFpsSsQmGoFwaJ6dC0C+XJBpunQQNLh
bxhzn2hWQRdDeb6ZBZa7tH7l+a+EIbKIYeDqF+49xHTdvveTtS26XBAjvsFO9Mgi
PMFk6ZsEoP0dkJqgkNDxOJQ4xLYzLsobPDlxvwSEXzxtAhIDHWYayc4KT1Sp2uzr
CS1v+QmTM6KCBebxu95cI00zL1bwq5g8hnam5gk3F72QpdzRvNk7XvpntHbHjax5
Ysnf+EMYYuN0qocvST/UYYoEEQe/EvmYraZuYs7lrH4FONGFAG7JzSWxrLenQGF6
iixBzyP6it7FcvC6s38OvqJ26Cy+nYKTej2Y0FO6TWByluSQT/dbqLx1hr5hq2iO
Rmmj3sl4rneqFNebAeGNw2TQnNKvjIZC9n2GRP8MsVRtbBoQhkRAfmzMicqQR6eG
a08L9/ahzZYrZFAm8+S/VeVhchIN6SeZ5wd6EV4n6uX6Zl6l0adWWH0FNqHFihNu
skSBqyTqYUKfSJ0XKPOj/ajW42iIGmFlRV4Pklz6rwMSxhnJAkalMsVrA8ce4Lgr
waztj2s4fs2VuuK75Ex04x95Lia9m3jMx8sf4Udwaw2mtG5uVuPS1gdW40+6zz0z
VEQ01jNi4252zC7b89AtikAqe73zkalRLfIfEKaHod116qJHz2prmKyD9osFHAZn
xs1BnWyApG8qdR9tmnh4UdDx29LoyKf2DlGriIa1VtqJj1zlCelQE6E1i+cTW68y
NLm5MA/TUKM6G2pDWvPd3l2zwjWaZHmE5H3HFC9wsbmy9jw0mmKs1Ex2jFXiHK+K
9L5OArdu91dPd/J6+cdXqu/6qOIbnZWU7XfCwG91212vJDVzLKnjCFF8IVW5LD3X
HKyNDc1ce6mExoiBNiNzyx0/a6vaM4v59wCCKdATeOTs/8hZ/TOJL3DYcK/644Px
s4XCRvs9laMeLZgP0Kuf+3XNZXlQOVZ1gmVdyMBQDdO3XwmPu0MUhHbyh+oVW1cz
8sw59ak2LUteUHGr7mq2a4cT6muV4O4/aO/Jg4hG/0V19ovdPYR/MCrAzUuyzOzs
oHRCDSMAqn6nSiMopt47k588E8SJT2vcePtXN+cpp2h6XeiJO7LRNnbqdBeuIRw1
sj3bFhSZd5lbNDyjUII9fXdlvC5uCuRemEb9o9oEWqbl3mYKd9L1fr7jJOU0xKf2
H9xWHp2I0wDaT8BTsAC7Mjb+brEzV3tUPgiLQdP19W+F3z3pYFHIV4foIVaxr5p1
FGQqoqx1GIo8tHX8/eDx9h4xvjNl31iUKrexAH83MssbXNhgLXym2vPymqTx2x6M
XlgkrmCTPhnXJtO0x1pF4YnXSSmNfz7BKIpkyWLV5hnxxrFyjut0PB/0nCHpuSUm
nGKlJla6qU+A7eIHuMsxne3KRleXgBXTyUsPnDO/1DcLVwHzV9Y6jERu/MH3Di5z
guNY7svOI6xlF4zNiJUeTTMU+pJN9EzCx3LJpoLcvgQ4SmStSc4C80db1Z1x0x41
ewnFmEYOHDSKID6fhOsu6fFRhYbY+68TNowY7uCshge46VqdtsGGf8291QtSsIxJ
alou3ZrOWSnlSQDjuNHE5p8jijq1WBS2DS8dXyq/xZbB28wRnHxHsaCKGcJlI8j2
1QfEiPfF/fDLAfKsg6uLOHWaK85bwCWRires6PFq+iRm1E8UuTUj5nv7ahtMt0rJ
HrWAhg8T3FEFRLx4ptxFLPwtL3eJWqtd2UQNwdcR7fDWaP5txcL1S0WcnRX8/Ajf
EA1kPpBoy+325eezrggweYI8ZC2qxbMUkDoQ23q3dSdmX8EUzRVqg6PX0/MQVOTt
JNB4H2ZhDnrP1zt+i62uyiPA4Uk0X2namGbLCAQjVsQQONKt4oYrwIy8IRlGq755
TCdex8ft9psQQyQtR1ZB79jcWDabJmK2qEwY1Piw2wpKO4wZMxiJxmdHCKOvrB4e
Jl5DZfhspDbSCwg0+00z/bxJpksvC1KOY7IqI/6tT+Y5xC77v3p+3n9d9FagSbn7
SR8f9JaoWuk8qby0oAMj7sO5/BPdzXZwVb0wXWZ/Zg42MXaGtGtHzB1xy5MVCjxm
GVzbO3e7ioP7rS9a3KtMPISVGRWaL/+nSaYI+xsbrlnJ0lcQrsabjsh4OE+klN18
YOWUFMskjRF/2TGK7j9W+GtyFlRiKzYUlqio2IicuD4CgMELXMZn4iMxLmxqQcEH
4KDWUAjBO1NER1f9AnlkqxsrCEC8+dU+anEeD+iF2vAGUeXLDpQNh5BphghSdbNY
+tZKTYzQsOqjy+QLFbCE17P+XakoKAXFpCcC011qWh3yRNuYrkXJ78YouLMpIkNr
6FbOzdiVd8lvJenoKjZNcCS2PwOhhgqTDdzBfESik7VBXTZFw78cApSrT0D1RKdv
HBWV+9mMuFCMUWCtIfU9JRfx19vH8WZsM9WGnbug1aYOWY0pT+KksV+6ZU7Q1WsC
EQGeFGHBNSagXleBeRb+exmnoJH7/CdvMYt7Bgxw/6ESu/1cwxMUfZKXPylGubCS
b+GBRBmKRl4/9cN/7xzboIE1pP5zFJQ6EpwyNg/upykOHV7HyMnYWGAonsrQF6RD
xKtYB7AHuQMmlX6AxYq465GBkt7+L3+w0k+Mm7OQZ2gxflxksU2M5Q/lHs/1Qif5
WzSvUJ0gO1Pb4uzYwpdhQLQuWa+5j0HJvW9bm1Z/RvflU8D7rsOWFNkbkzwqUJIO
Vz0qu11OA7GlmZ6xv80LYXl/9zEWORdlSy4xj7dITOybhNfLkdDineBQbt+BrTMq
NmYEo+6KzRDGBIq5ud9z/pFOrwX3OSeyjF993cN84tghgyrLQMFrp68gwBhlXmv1
jSLSDMjnKNkGmN1oLtg3IT2DIoWYqykmnkULFxzNH5oR2WXwnVzE3VyYiHDxl+m/
GRAg6P2Ub0MHJdfFXdyAtYrQ8QKCCrjYFiy+jUuhjwbgLXO1nSpEgp7oc9VmItQQ
1Ff9ktLFWXwwF4dHomBJXC+nOpGGBC13uPavciAXfn6fTmN+pj220sPpiJrJRish
eAhA2sb1eTkjJuFyM+Qpmn+AlSNxGukCBaR6yGA5SsOMUDOV2eiuL9Wn4r59GOA+
Em1hbmVNfyKtUdIOjTXq2Vr8j1x5wLiZag5RjPwBbkWQJKI63yRrdNvNrArT1ccu
hJgL1KYtqLH8FaQtZxHXZf0Z7/a0ja9DzKcneOpWQKWTCwZ4Kqp6K8zaSWe7AK4T
SQonI/bpnZHLxYmt5aCPOwN3qgWeYFsOuH1LrlWtJctKLC7L8BqvxvcWh9ZdBKid
54s3GwXzcgbfM7b9cdeKp/WuQlXQg8iyOTwSws9L2xScEcfqkjUOPM852yjvFNJK
91t9uUC/symLsM3mgWofEQgYtr6vJoJuk+Tu9wHzWbdL8Tr9jBnQMl5Ei2/NxYC8
8wrkXcZkKe4iZ8GcE9dbMOEDnniz74YOMUYNyX6+aRpdyD2DBBXPfZi9ZVpPFgvh
gyWWlpF1KzpQ0cJ36ZX7owmyR4ePP2t8ImVOOZRsattipwAFtUN8wUohlCjcJSBo
KgMR394oJrXYQB2J928ML2grja+irnPngn0oQ/wrJeDRgstrXHmLtuNsXW93L70I
nsMi7t132s2UEVL77KDRS2XO/J26kJ7vEhqZp/ikZMuqOEueGrXULaEwTffm/ufk
ROe5XnZC1oNyeL838Pdk3wZ8XGTQdwdARjEg7q6rHlRVK7L1ISTGSeHK/efI2fNo
rmPkxF+BEHdEnTCGuMkCH0R24/l0pp345PtcFcB1gizOf3alvn0DGqjIZFXWFu1r
DQjLfMddVjGVX80yvGtg1t9d3AsQWaIKQIew6vDA4f8DmfophQEhFWkfbKP0pamy
fKHlhXssGx96CflXRLtbw2aR4IDQVwIRANQSU7NlvKo1T9ng6WVJI4o4PWLJ1r/5
H1lUcf29m1KuXPur1dxYFvA3BwzQ4xSpgfx1m+3va2E6KizYkxYlC+F5FEhCux/y
OaRMBw4ArPw0o+MYC0giTylNFw9pDr+uySlIFE2EyUqxqBQjN5qr2ka9umJBGN3I
dRNts9ZO+VBE3aw0w7C2sJg2zM9tVyXe7CMJRFe3I87W3cGnGrUFA4yTMmehCUTO
7ENSvP79N44QnqdJ2ebfKqFpjJL7Tu++gwKBVprxvclGUekeyMV4RdHpaJwa+QJ/
x1xrj1A2SPNez3EpkKschv+FjVQlPyCYewddJUu2KXtaiE/Op/4gf4Ta5KQpiPgi
wCcwnws49jlcGwfDzJmjN3b18syeZuuOAuIczpIsQ+H/TB9C4DrySL5c2xEP9thu
28egRP/QvONQPoB9G/Ssw8p5MUsNQrRIUZFCeVfU3noWyTrV9EDyOltb6z8GIEPV
JajFHNgJ/9tns8qbe2X7Y4xNDd3JQGt05j5dRqTYlCUIzFpP4QnHJl3rB+ZphA87
iWxGJWn9E/tRe/SvEuV+kQJPQmy8dv/SC7yeQ+mGsww2Fj6Z5qg778eWRURVZ8zh
/c8Et6B5GfGT/e2iv8iOcnfC3YNVmsYa96cCq1rK0b2znMGHQY2TYl78oH9u8o47
/FJlZWxRHJdoaiuHo+2QOXtIBEJnYrBWO8Os8ua+E30ddQyFO6Hxfo5pwKxGfEjC
WkRk6u6NuvKTz9yLFysbU7kP/XOEXIXay7pG+xzpEwxv/Voyjmt9rN3qYdu871d4
2m2reVyz7U6j70IPaNvD0gdjUrs9BFKKLi7Ds2FjDft8kmHftMTzLywoo4kUBcvn
dgU4JBJSI8+2N9LW2VqNkzXukkSVRH+HS3eQH8quc6TjjkD5raCd/UW4uFXcDgyK
Y5Dt1Kjcu4bBQ1JsebyQyxcBV2zU6AjxG3TBNTJWWyLrB4HzakxHCIxnSdcgvnyX
oEbUVMkVohOQLuj8U6t5FHMxlkRiKTLJrNeSwXuHws8g8DhETyyL8KnXLxQeI5uh
1EUJorsCQqF6L27+2umguNlUa0eR1or0TJhjDrRnl+nQ5fbc5C4Dpwi/RgQr/Xup
jxpo+ajLqorKNw+CYCuwsenbesk14K+KMuCmTGZpWTpbKGm0i4iAa5T8G6r1XjT6
rCyZjmWJXZFGCYaknvJoThTxv0lMGuzDuLll14BJZD5moT/nJeToxunGgTwvrITA
U7wgpPhiuEiSdSv+i8zqm4kefXX3Qd2WsKGDFbIgKZJ/gw4wmqTAX7RZEZT2m8dd
GKmFg8Tinz2ipO57WEngab6OrmoPGSMigbUPhAzghvy8fH4ln0H10IXrRigJTbTS
S9mPyQxi+iDgLXaWp3Jk9WLvMMyKa0Jto4JtTL/06xliJQF9UOYxl3SDsVJQESJO
5byokbU1HneLewbTEFYjcshWQHfYBc3gr+urpVcbCF/3EI5ysyyS7iVxfyzMcmJa
Itj62000MyRRWh0DE/gGjcqq66CJw225CiY6blHDF7p7LQLgqI1lojop2u9GxWpa
KEJ0IdMl3CXx4u6BUhlOeZAHZObnl8gBs/evJLf6Ika6KGLKcGgjMfmsChF3Ff1D
oNYsOwDsdB2YoloozZI2U/APnwpEz8eYz8/YE+IRQrVeYwaALHo7+xePd2nj+m5t
3AAW0GwIYaBXMsJ0h9c7LMTHpwDvwxuekccC3GFwSRwz9G2NMwXpWAfN8VOzpqJV
HE0Av+kSQ0+XiPs6iczSVuEyoDI6u6zKqpQAhcGjn6HRcgLV+PykkyP5IXo4g8UX
V28M6rSJRP4KvKCGRmryCCbThbZRfnI9UDb2hciahmcl+Ixx4jHWQJS+QtxdF1Uh
rHER8RqSTcu/WFloSQ5dlu526leGXRdrWYBBwdbGShVMlM2/wo9UgeWHxFezJYVW
PNdqxPTFuwEG0AEMopyes2LzliJWPGe9JQY6KIwu/uVvGyJG1vMc/1E/Aa1w/G8h
ib1hft7FanYK26PviBhe/SQi6afdh6xTdldmMWTnghb0tGNa6WvZiZeGL7kMkTgz
dEcPp7uvVdtSZw/y+fLCF+bG1a+K3DltwImGlLAWHCg1Rum7K3hMUzGQ3hl0fyZi
tSTLBepqKnAegcyeM/40amFpq+GwRg9l/SN/cU6mb4Ca8U6NRHP+ppfcf65NS9Ug
NAEQAajsfn7Sbzh1qsGiPYO0zpJ8mLjCKXI8Uwz4usfQcnL5yOR5aMOEyOnov2ba
b9tefCkheGdu/DAxNbiJEtWAQoEql+NrZDl6aEcyDEcHZsxDbJ8wH7rZ5SHkLJLe
nwuQOIJHmIGCSmIa49hAWvbglZkL5aLZzQOds42cD/PgatfGjiXFE2xVlOAQdEaq
lmI+75ThdkMVi5vMQKY1TknHUmHSU57t8DdOs42IpXqFTN/Pp5q/Msctde2AblrI
W95oU4IDCiOoou02AvDc9agO9QL3szWwbRtj4DPgoK6vU1iZeB29KkfXF7X6nsui
rthMkBe0w39nK/B/r1cLf+yeVBor+Wncz3Jwxgz9gRrHXboUFlmpoXxopjR1jcoR
l5f15l1+Wk9p7Tff4SPNqigJYhFxZCqEwoG1b1UmXpHCMw1beDciPV10Ta6uZNEf
RbebfCcBomeUl3XBcXEpSQG7LvaeS+HlNTOESk+XMda5VMS4hmNjKwAOKib+o+FO
9OJ15fo6AxEepDaZtjWNa2fakqOweI5MRPxff/jR2ZN/a64jxvjBDdEP+sjkVEQk
Px/An2ihgGh1jZgC54UMrf2WeUhJguQ6EuFC3NygwqYKAvy2ezwp83qNxKQTZVb5
n0y2yMMUi84Xf1zzcNrnZb2CjGE77Lr0Pk4D713g62FZ0WY8i7O38wv6lKHn37uV
MTLY3zujCtQT4QF4JBF2dZ1EbelnRgWXnMq7lL6oIOxQVvvprASuQ4lRVFa7E9cj
IlgwR94ZkRkPX1OxzUSwSRbstp30t37DslbVksLxtql/ndvWmiTwOof7zWfwjgo7
QmnLtM/DbKxM6oMgLoCJVCHeew6KZBh3zIRa936+d/W4ZQfZXkBFOqo5YCGzBSW0
RARW5TAemTwX5BnXtzzt1d68Thje4E+YZSrgUTCWNtIFF+VupJyBAwK1rBDQCOhC
19I+xIuXmi04RAAlEwTHZYIdMRBZlzLzAscdVL+fTFljFVhQPvS1/5UcqklaP3ME
641qxHDzXXbkqNlyMW5FCtUkgAWCJJi4nw4+plJ/wpOrol3SgRF/bUUtiJ9i1rhX
pTGAxyZm2xW4n1FUJ1VbUmviNurL8iy+El6f/bmf9mSumffn3yHwyGUOpGbDynDa
OlycYP/6ORxaKv5CGn45+tz5YQ7uI3ybytINWpKzgzuBd/w5sj1Gm1wh9jOkO0Y4
/QORH6NoEQk4vQifwPttHJ8LjsdeQHcTL4BddpJ9aS3yd8nZju3BwHHlB780MyBO
ppJrykJdrx+H0fC+SktIMLtGuSN0Gf0k/gbPaArsIUaYyAd7GnTBj83qGm/80VUo
B1VX5mcXlvxFuOnC/tmKfgBI83lfg4WyeG824bJLSorBjeaF/4K8uxbHQQVe7TTB
oF+Nq4TG98xixIpLHf/E4Zct0dP38dmLsxcUQ1zf1rMDAqvsPIdJFnd95sOnA1L5
8nOVHmY/VV+m50+Pc6Yx1Rjtt4wKWb5EkEoq5oCTKrvqvedWHk0ZmQlTpf122h3S
hYK5YdYOBHND9doozr9hRmhZchcclsjfze0Wjzf13d0mZnnL5Mub4haLyoCmd24e
GdyGai5o0XeTVV+KqamQn1fsjPnO3gySn7XoPtwvxAhr48gpdYI85K6wTvZ9YL70
0ScmXN6OwTmkybwdpNza+L/G8WDsGuFNcMWDtATuOqqyoy90n1kCnxzbKWq06jzU
SRrw4UD/soxY5RR0EaiW1bZQri9yJqUoqWs757EY7wp+nk0UzTLNG1CBo5QfpHXb
K6PCK+6ZTwF9Pj7Y1CT61MP1xgFP9vmvwZ1AnsFae42E9UXPpHNliIXEjET0AbVQ
4QEAiXZjqbyxRMDCaDREWLK4H3lFWff6+/OjLHXrwcoOI3eS+jt76NDaoD/Vakoq
ESGKhnZUQ9KA688HYXgbIv22RZWiIjFcyjSMLC7CSjBY78o3xgnlLWVmd5cRePFw
fKUbQIY3Be9mxqTvC0TwRLpKwZAD8vqAzBjIdWgadY/zU6/+tHdEpSeF+f1Mjm/P
bfTaFOK9oElRNXU6eJ4ciW2kML8TWE/hYtUN4gEOfbCRPxsoDCWkgd54h8VtoQLR
AFJ56jBCNsPp8i4jEeP5BJiF7cEQVJ3qyEG4HvRNJg/EZFf1zBrFP+7nnXOavrN/
CKpSq6kw13NM0CGMnK6ECqOr6UJ9BD193S0YU3HD9NQOIjJy0Ucf2U7Iq/vIaB7Y
I8dYuaJ9tMXDI6PhLA8Zzyhzu1eSur+MbqDA1SLCDLaIpGifVxe4sfuHx9bOCSk1
zYAjYbbFE14hdcM4odTR+M4KyllhzWzCAzMnkoyKTzkPnjx/etnMGTXXrraPlhj5
KKCGdlqEp5CaX844in3Pn8QVDOMhxg+/LtD3gWJ70bMajYoHq8kQjp61I8Wvdjjl
8ieS0Ue05VET9gDBRI6zhB5QvjdbHQQbe+1kmSGW9NsDZt5WDtfD7yzkQUnnIsdk
vxN1X7nkX1MYClq8++nmdfq4HT9mN8gstsMF2YZ71/s5JaLpqiFezdX8Q8iBc/eC
oPGmyxzTFC97DJKNZe9qhztiTwswoX4qaisCRJkAPq/8ajxPoiZ+Yztk2N+bRayJ
3V+sG6szG0r/+g3i22/7k4XnsTlyqT+KQJqBL0bavx1kolnEAHJ0yFR7Nh61Cwyw
1iohTKunHOmGVCyc7l7ZhlhqpZV5mpjldSsmQ7sSJat0SE9ztZNaPH1qHnLil3Fq
hG5HqKqnog6fkiSh7j7uQSj+xt0kuncNEnLOvDUrlWGk4a1NhyhSXPU+Fz+YGkuX
UsSaMNi7NXcQ8eNbzwHY8m8WL4785tKQCzI+0iWKh99LtGI/bYXQdstbnORSh53/
ufo0VUbGIetiZ5AMonzDIYOX6cn+xOOji2RWO9MKxH8XY0rsVtRs1KTsLWa6ZEnq
x2lZmfL7TK2hdSGYmQrR9pAJmJkasj6Ewjy/Lj7eYIJW/ciD5NMApDRoW9rwS8e/
Kee9RQyIbPh4adRYzi3rgqaG7VOslBkSNsH2AkDxBmJpUy7A80/xaik0BrrYZDRD
Gl6qYqbjl7rbX1df5Ae1XKvZ2AcLIvwni+fgFhcRL/Lmc82ccTe4/Y6dINBSqDIs
k1Esx2WcrjHP1j7CAbtRcI8fE2gc6dTdKpyrebUn/lBzqKrzubnZ+9MQm/uZhBEu
I2EKUT35DDa4HyK/5rkFMKVszf2AtnWoFJ3ZuBn6RRcYHeCHLfN2YOQ4MpzRWlWZ
cO1+rvCgWmYETNlBHSwBVLkhTl8L+n5ZTLSL++EnwrUE5rWUdwsV61nPX7xqsTOT
63nDZvwqOlVgiabPTXmTTbO4E0IzTp4bEJGsr9baPx/yEdb/PGIDUmRU8NavcI2h
v8BCjxjGguFE9EYNjEJXjsa93yH5LpfxtWYZE2kUczeiw5phUMKZK3mEPsT5U0/7
VPwFzbYD2m7VlOcL7xrjHLj43fEGuseQdpQQ3GCyzfNpR3gnN39ggiS1ScKWmgxc
jQ0qL0Ep7A/x68zXGnx1TW+1c6XFOjP7vEpsXAnFwqDUKZUnGNmKxfKG6WmBh1nk
TUU7oiDHnHlmjJrTDKXiENjMDHbRLE/SJ1eiaOeLUbTmutTfmrww2KKOHhdnKHBO
nVS9ILCpNxuovEiYyHiFwqokfjnlqNup4A3AYcY5YUUVlPj3lj2kyfNNdDs/pZH0
8Sk3Y18Ue/9DsmYmQ3EOQZ6u1nYw5fctXpvh3xYCF7RcqFvl65BItMgZhQ9bw7U5
1eWR5GuVGuxalCsuVioHOAyMVS1VdYx/kYWg8OjySePkeqGpYGMWX5ER+uVl2DTv
H5S4ME77ayMC/qlP2Jp0VBg/2otHHy+RZk8EbHZnjiPI55kedTZzovt0ADCpG1Vy
S9EBUIwqXS3NsPZqaCmw/SJZ9RGmfdQrTVXMRJ51hN9B3Y3aZigKJQH/wSAh+5xv
EgKg159mkOxuTIy2QwiylDmxN2irTkKPyXZrnwCs9EPWX4HnmxfT2yF0vwJCV4Nd
hmLWyn7U9ZQ7AeDmN/y8G1U9dRkjkEj9DTJ5NLS4eRi30nkQcgt5TTsmLrH/AQb0
poD+3SpciRcehHll5LIr8zIYYIZQTkdCG/HaexPz/sDkMg98oaTLnG1nXDHHwFu7
j0KgqJOsknuIUz2tANfR7ubI43C728PSoELswBV1IvfiTdTGBJOnqOqk+eMkMXcg
5ht2yWaeRNBtR4LbVVjJoSaVIJ+ElkuJkfFH5RJyhRk6AfRMmzZ8yxMBcBXPigUC
/Vp/RWxVWiZvySd06UzC8HFT/HBSwD/Xop9zkeVkvCYmaIjyYpcnkqJOHdussG7g
TnOCk2z7bpfih8XG1W0xr0Isv4E2YI8Mgtp4AIoxv4ZpebrI6cXFims4w977lWZz
NnoXGAB3z4M8aMeLEAlPza0BIIo/nCaB9hfeLSOm9XN6R7Go+6s4a6nBe/yPT0GG
G4PTYioj9+Vu0noBAQNKX/lSNjd+obzL5Ek8sKR1JQR9F7yDHxmrSyYtbS13j1jB
EyqUf+CBaQUI+ffFMkuMr3LCVatJyb17zZYjD6jDRAKu3JiX/9lU4Optwgs6cX+V
Mx6D3NnYnLBwmbwzz9FLxJywxgy0tOFXhVYfpSSf+zhnXtXcjBMyNBEZSqxDBPSt
+0PKLNrjKyiO2Fi8x/bvLOnyDXe1t3EstSpteGOSQ8GGOGK0a0VAkTjJq22rkZd6
oMH52AWgKnJzIv12cPyTU24pL6ZDNDJaB5wWtG5YlTVR6HwEpwNY+w7+A5xYT8tl
P47prr4/We1uVLXKxNq5YlpOq9YBKeCP6d1aQAmXA2Jr3Fg+FNTP5L8fUaUNOU4S
Ti1Ob2D9MYx1D6G2c/xjWl/LVoBb9WZZ/861dHhpC7+hoWnZWB5lhnt7yXkPHW0e
Hmw1XqPOevWI7/FKzlx5X1ydt3mCpIpwawx3WzCf8WKOMbNjfK8OaeOM6Iyf3dzd
6HqYsT39KWnS9S+Pt6eFZgvsmAd0rEO33XeUDKJGSLiZsXjUm1Rnl1Rc59VwR5eb
fLV4PFnGUJqMJSzIXKJE5Tv2DyJvTVTW1IQ+lo0D3klw5WthlHrJ7+DU/1FYkHuf
e7D4ZFAGF61bpvvEB804QtQxMziw88fkGl2vpjLbQfBXE5fdYXb4yDCuFBW84xKd
P3Nu76Qy3/oxfIcKvMJt0fh6A5p1z25vRkhxHrabX4V73SUbeDy8gsnc8L5/NqxV
YfwK7TjGsb1Kg+8LNNAPYB/93EO9YjlgHmDAZZQy0ia3wsr0wByHLRYufmWe5h5v
zEQ74EQb0iKeiPgDcge0hbLznXE50gA6l4Au3I+oKNl9bdW+g3aRWiK88FGOMCfQ
gx5WkVlcq2Giqj3uqSCo5A98RAm3xonQ+RbaZNmp2XrULGAhd/mRAQtojRX4dbLd
AcIfUT4X0YdBIFJWRi7v1LxNyRuX/EmhIgUJrnUBz7tXNwei4z8X/KyJ5TH7Po3f
mBzjyX+3R+q3hxypyFzJN5CvFlHXyzMAm6g91g6IsSxPcw67smkv6ZVtZjKTKPyE
zQrRD0U/DMefVY1w/J+lh8HwKqoEaevPTWp60s9QX/QC2IsvA43kIZoSJqs87wQB
3/VKLg/BydK1T9ElNooGj2rJLmgPqZfnfo0dOsNL2FKCpQjpFku7i8FODHVtavuy
O3SS/XrEyLlA6M3kaxjve+dqfwm0YQ7Dq9wuCO+0oeVfM2NlTEW1vuKHRJHsSXsf
jcB7lzxE/NXolvKAwFE2NyY48byZm1CLsQTmTs1FYLEnVoY1K2JJtD3m5Ng1y9Kc
TKiNYqXMpGudyp9sXep6QXRjI1n7PROCqwauf887PVoLuUrfDwDGNOOc8uK1Zd81
yvxeqQnAAlENCCqW9Cqa+oUbroXSU9jfQWnRbbt3H6q+d6pgHUg1EIxTTSbBjkkF
Iu1c5fQUy3XFzqGvx4YOLgg27fMrcjuZd0xLcj8bgdrFx3khxfBwKGdZ6hg/rb6y
ZaZtgI4Wuf/gxY5YCEDOKLE0c5EOezVqz4rlbwN6L/oZvxp1w4AM9rZEb3SJduyp
cQ0koUml4K3yCOXUwtBdC/bY1HGFoVSwdWMQ37tgPwsQtjpV0v623h2Ciap42HSv
3+rTghQvV9vnc6qW8x2EpHh3AuCeiAYb7A9NOHC8sGCW86PGfA9YRTncfpqdcxHS
15dcY438Zvw00bQV3mZhKk/BB90sN+8OWev/SVUZ/9Zx/n1euw+oH/fvS0OzIbCE
sm5o1NFC4MRo8lo7Yf749Pio6Q4tx63s+HBovIxrGyHKCz13Wax8dDgIGGHafrI3
+yQqR8HqRC4jU2ALpnMjop2Obx8MthlnwimdDTB0v5pKNEqSX63HmwtS+S2/TGNF
FsiAE9/jyfxF8/AVasPMtnhMitDJAaSII5tsMOduP02lk16KyJvKc6TVyXbgF6ym
B8uf/TiO9fMylF9h0jpainj2FpOBfqFFNqfsAad7ZHpwsII//iinG8jE5A2xcDqB
JkI6MQOU+4QUZyxXyk7GZDOSFMDVsFIWe7n0jg80XYAP/8midSP5u3QReNWlCVtq
5BlBuF8o8TvDnXr0lMT0SoFiy6JlL2PZEMolWWI+ETDa2lz4dNflq5czRuJjK1sE
9ZWDf2kRuNZ2heb0jjHLOqKWlUWTnf7JeO9uQUw3tmYfTiIY/E1qILZwdC8e5Jtc
nZw+ZrdIOKRWrFuHRi++o31z0rYONuN/zzrXKXj3ACq8Z0km3E1r8TDTIoS3wDqo
OP+yt1xlHJ+sUD7bRsil/eKrATY8h+WEVxiisIaoOeL8ngoYbJE4/2OECyen1kLO
SmFQPUtL+NPIIk2vciiBFIUy+1lF8nvtYBbaoqIgbpaMBmkWNzh9m9poGIRHnDm1
Tl6xVuLWZ5XlIrIJuE+cXsrPa6PeCBi1uXZKYx691SCAgxUpWtBsGin9HWqI69oY
SCp4+mjiyd+vjYpaa9HW1nDk4LQpxe5WjD00EfrsoKwmbyBIgSeMP+u2VDPbNGfI
PPz9SuVQb+A3MEqxVVkl18PdWlB5siM0CW4vFF+vzuSoUvmeC5Nws2PMg6HkCCsk
H3j4PtzyG5BrAyZ+tVCzh0p/tiIh1Dyb8Jetm8MD1Kh914Y3/eiAXpWKlr/YlVk+
thsrpajLUf4P7Yji6vryUsXxH4Fzv4m1FdSdtJ8L/8x3hisuqd+Xf6y1HtvJWLpA
8BwCpQyYhZ+Ybs7mL1LAW7y/id5LvkD4CJHj3Ah8W49KPl1Yz/Qu7WRmuhuDVz4E
693u2+angC9uWqKbmUzR43I/eDpRZepzesjXVwpIpxxOND2Kw0Fwz9Pc4N2eh8kI
E3qGsYkv7ZxLtezkLqa4ZnT5nRtoCSVc2jHGHPNdAu6VHW5dS2xhG5IhW6PN/kyE
vzUnD8Q9KPolghV3tSEQzlPGZY9JWddI1qDd5jkHSYrDeUwhjlywUejqgRzATDZr
Fg2W4iCZnmOxIVhlLQrpQxJv58kgMoHy+Hl2ThPc3kAoq16V1jYdKzeT+wbo5Rzh
uHTfULZ5ro+h/6RbvrHnhxYa4LUaxFmanRnaiqB/tBbp3DN1NnE9ykhig8BCVsrA
3E49V+XtbjTcSXpGNUQzbL5TRccc0LRM3Qr0SJyQHAFHS0WT1svKw16lKP9sTwoW
ytZCbxgKotKvcnbUsgYa4WqOITpALRaEOGKLGRq64WzaeMLxUnsx+wc85uubDMAJ
Sx2TA+faRlL8G1EP04bnqhPL4mUZ+Vzv7fIHFjE4o3a2S1GbizbGOlW7KcGhEYCn
YLSAO3APiyEN252KI78I/IEV2rocUlgD47knmmwfUIWO3lPHumxMORPp043Q4jzE
2Y5VfdFZ/Z3YtNeX+VXD4MxUSjU0XA8WgYui7ZM/rTU5ldRwvGI3b/22O71gDrOd
nggBNct2YBiRojrM1C7eKYc0Ae1fv4acHW7EkO9BF5Fg42N/JxhK0m8IGRri56dE
VF+hT5RuVKhrrjxOymmsVjg/AR6ZMu3H/8FUFDsd3VqQIEVj36YZqE0fpHOLXcjp
TuZCe3dACKUwKEtyRBuT+5lrelXUDyeYr0R12x3K8UrPUORaWdfrevXHyhST+UgC
VLyYWNkwM3MqcsDDBwHPBk/Gxx0UQ7aTDXUAFObgSZNVJtEhond89Icp6/64gikv
kbXayFOcqfytG+dBPyV8/x7ZTr5bmuaGfgTrtaQ+F/nRKJOrBOf+jJRjPPjnshE5
GS4673/rlqr+Regm6YDzI/bSS+mMFEDJGCWw5jwS03EU96q4WoqRoDvG2G3RRQ8j
fvvNH28kZ3eyLFcNtJh7FtuTsKPKc2HA6iruyWknqvsgyqcGglWVb1rIsKSz701j
mtOEcxeicARUCbcjzAmeG7KtGPgTkwR5V2BgPkBXkZeqTF9luaTz5OLIV4Isl9nz
69xZWuD2TcrkBuYnXiQpeMor7U7H5pfRWz+KIcCioaS36qDGgXAgyLHQBMs6nh5b
c49TStXUc1CXDcfL8dbcr55woDPNYgfnIDBCNwmTlwunO/UayA2yzHr0bw04M5Hr
cFDgrCmmKSqEbWUlGukyP43aUNQOZ9ww6lQAn8Bh83faRCa0+qns6JpDO9c2K/+Q
JH5GBMm3xN57psh4fjxjw57/OlUDkTRzNk5a/nA8sksCqCHGTygh+z0JgPvwIn2A
iIvi87NwlTmzWskR4SRGOmfhZsiMF5sDsTJS9RiqvVZ/HQBTySW0faZLdZYeEuAp
SK5O4aX8KkgX71fxKGg1oSlu8SbgRrPVzY1uwaJc7LqxWk3lid9wv7/GZJMAilUP
V/d0xB7U4kMauVfkl2UOMSw5t65AxSUdJEeCkMbkOGhT52/pZvkn8AyX1Eg/ZXyA
muhD8Y+jczdqwCwTJZB3+o227ee2FJFi6km4hMlShfAKajwq3Y9vUu9UpOOMBBQZ
2bYAcLul2V5+zDnok6hq+k43klTyNw+fGULJA6o5kkNWn3uVmJfXtYeihyB7Slv6
n07f/hX0zYR4EG5fRQw7CUnKvZPpfAPyJRQwzjW8mYfZVlfvT5y6pw/eBRLJ4qkP
CtAOMcPJs+TXNKz+CrsqV66oj+hbl7PL6cV5sNMDjEvJoK++uMuxVvRrIEVOaGrR
Tg7bjBmLdkd9jHSjSg8Qk0FVinfOphHcJuA+sLFHOBlsyHfbdBAdpJ+a+JwbYLdr
mAcCk8Uey/dHZ+KipHHfHYSDnzPyetSj37eX271am0V7aQV+5n/REnqkuVqXjbbS
eVNtMXxM4des5FkoHDfw4OEUIfURIHi9qMmDiKrUFX6pHfezMYZpDUswTHVOCIDE
Jw/l9109m9wdJsgsYgClSBrUrlITbqOG4Zg6aQqf6JszkuGjZEyqMA0V26AXfkhd
+ThBv4uXXmH8wEkuO5ZvXGPrGdeTXhGf4qmwYS4PSPTsz1BfbwRe/EDqO/HOqktb
xRFFu25BQGB05bsjUJ2olZJg6jDs8ojRMPYYVrlK+xS7FNnatnheGMCSi2x22kYz
rAf2q4gVsp3wnVDpg5g59ns/hKdmdWJeqizTD9fStoY2ta5E22EAP4QUAr4ZRNVp
GA4OMPH7krV3GAs99E/qsXOiL5epA2pQbYFkvrOGvEGDrfL2Of+hQGNzMNPcubl6
RyOYu+JwQl6oyT7Y6XWbD6i44t0UZhX76VJd2jQKn+Cz28whrCKFFMNlr3y8HaZW
KacQZ0jqPfkujR5klFJc1omC7pWJoyiBWkEF9taJhF+oEGx9RaE7jFMARhsz4e/t
vNTNhpAhIeeMO7tXeTRN5fSgMaU0zZo1grJ3WKiGRDNBW7qdwzK0X0v8BhJhvy6Z
U+TScWv1LaedUIp/J/VgIe4YkckCUJJMsBEp7LfhLpceBjfg+G3DkNNoDi+A9CT6
hzanbrahunNeqb/nJfSrwC2OBYEezYNeURWG9O1Y2GxxRgywUjxdnLV9pFGv46jy
r+8GWhrjcZRNZjd/jAmsRubvzZQQca7d+JePYsBfVRGXWt8Vaf1KuUT9ua0hTGDh
ALByHTm8Rl85Z1j5Cyk2sun6EUcIRia85+ap8oDBfc9LXqbWgDohCoghZtj60Fe+
tRmwmj1K+M+/ziRJM6kIugJoJyW77BSDhAtUTA83MIYy/5nFoErngenMewEDsSIg
hwlR7CjIvh57sSMWtjSWrLk/DMxemNJRWneBe0f8X9nSnib/5HST0tN/mHntXm9T
YYgpFZrZpdbgi7DOEymV5LGNqp7EWxdjQQuwJIWFRXoi7h7MId33czJGP3VVb2Ir
IjRGmaCpeZHrCjZ864DA1vkPAveTFxYqDg4Ts8D/NesEAVMvKGYzHdD80WME7VWQ
NeqCubMqVnrDBhD35CPL5PH1hdrCNVQelNiTx+ikmVYHXXOXO+0JDB3Ad729MH+I
SaBj16PV5q64bALEHZBdBqgKcFHU1w0K+BkChEwg++NJR+O0aTBwWrNU1Qhl9o+r
Slr2B6ItS5XidCA09UqGrJHPYJJ8xdJLnlgaQZ0Ox6YNgDOPjmLo13VkgL7djK4V
JDvm0k3A4u9fuEo4L1sg/KrKqlfWekuE9sEetPowjm228QlAQ9dBDSKr8HA2ev/C
8Hgg+6MF1gfWvP/B5X/AI2hya+Nc731tRV9cVHyb04HomogGJNOmNJwoCZX8ygPp
vjf3Wc1O7A8Zq1AhLRcoSKWlOBW/KrLdOGboA1Z79JGuLGH4DLrDJ3bvoyaOMMU6
WF271skRmij8U9h1tVm+oE1qSDkxlfjhwggxzhREcuyl1Gb9pFr0E4+2Gn3+6OOS
ra4ILlfHFy/pdNa572NUhf8KZ6BSKL8j+kwLuOoNfA88UShpKmJNQwJogO6yQKTT
VonCxbOY90jGioq4+FP8Qx8HY66lwMaWZ4CwQ7yrpTdTRFwHHqYn+fn8ky1RfXmo
0B//cJrtWC5zVdr/FG/ohj0hrbfSsRXLOzYt88MiQVBORev3lM5gR5Yp82qHZYlV
snMcIzwyybPb53MkP+7a+IAoGcjAG9Ygb1nFUxvDfXr9f8VTZTvu//8a6aa2UVnA
Lbbfd5lpNQTvB7BZLXzNN68U621CMw777aRnyoXrwsGzHb7RVk8lRjR+PY+B1GWT
aVTEQQS2FuRaWan8qNI20Q+lM097AK5pDSIQr8wv1P5j+fwRy/rlT9eFKfhS2LvI
RJBjSAngrmiQirBBH1cOYD29XfYHcJUL5dx1098O+hUogyB2+ZB77v/BL8zd2oU5
eLkpKkmAMUkyPwGr0VA6FITN0isyJtbzLoV0/h2xqdLZmPy+QojgKTBDp0aKrUVH
tItr58fonb3JqHIxjD/VyT9tPM0/cURlOqlKKRV4Nw+twbdWtbJJNgTwIaLGqPhj
VZ8LFSGYtFevzMeMELVCCNCtY/gjXtA9IlKrb7omAGPK8y4cCYEfl3vIRkCjl9vS
2LnMcxn2bdG9nr3s4RykzQInbMAfjSE42+KGF3PWudH+KJ5KBJp2gjMzTpbpH+PU
pz2Ov0yCzdQZ1wq0CYtKEtYPlyGyFH7fDwNCNiJVMisAAz9C9imyeDlJJsb5KIpZ
AJFi3Rsv+leMFnbNT6d+vd1OG84vMUoDhv/lDQhhTnUSzCPjgbnz+eI6inqbmlR9
hIoDEO6lG606d3CEpI71Eyf4DzivNjhACTNCA+an/oAWdEozypDbLsGkOcpOy1ej
FG9RqKTfAebGRnR8FrzvunOOrmqGykOL6+Oq6KM8C3KBDv8eciit+i4mRCRfMfm7
S779fIei+EKp/fHRYqN13ebcuBVtjACg6aSpVL90NRYPX9O0n6aR3ukDfvu8IDWu
tnAtx2x6l0GGqyY5opLm4C86iSCSTVsGZMq48HE72xh4g+c37dKSG5P4/Rn92b1m
meqx7XIIgLI7s7dsV8BTrUiN78pyY+1gslqy7BWlXOlY4QY5IcORsHkToCbb3F+7
Fmh/lioMS6XWWqNJv3ZlyhPBkgcIXRVBwVLedso8fykHZ4VO0+6a0GUFA+vxveXF
haFb8+wyd47mJpu/okZBOakE1ftrHGL5LMGcJRT/3zmqNsxkZEbquDT3KqdeIBmG
mhI2hg6cQDcJRsVWDEeOeB7I9Wg3/ucrfxCmfnN4LDpKQsaIgiYzvXP+q+Kxp/x4
35GzveilS8A1GAvegwb7N2Xt5VFR6tWq9P+xYPT68KmzV2LcvwT4rNrLu1DGHNBC
ovaXU4g09HEflfWzgOkpT+NE+O6YXq60YVI+oshLWZ0M3zzx0I+JkCzS6Gnakr4L
mMMciqZLY+/ktEE4ERXdgfJvsbyaqL8sk2gthgW6aPgdxDy5+uIvB39+sH73y4Rn
cVE0xQH1z4QVp5z3kLd91VO6LsUu8XpdRMZ2Gxd1hGcdYWSXaAH54LzalNdoMy8R
wUQ8YY8wW7E8+/ItC5lHg0hZy/XpPtaVX//ZrpjkY9JqSRsZ9qwfh+ILrQlsB2Kx
6YopS+UlwYv+wpPrkxmfhPVW+zFO1QzkzWFQTFqj7yZaJYFjaYXaMxhZdZUAAr0F
37Lj/eK3OtsSjRw3xQ7xK3txe7hIICY3UDD0eVp1NE42vtrxShB8OcperWyfVMll
ij87wmn9V7Mg/otXKsT9Jji0/8uWGsJxvlrkaAmvPpUpcVkDZ2vcwnJJY3d3tjc0
gQsNTSuOyAPWb/AXvhj0At7qEsU0j2rcNzel+N2TtvGIWnO/zN7vfT3JRDPAY7ED
I3k31PiM3/48jo0gSKlAVSK91npTMJYTsrUADRkzSb4yn/fe0ANrVulFaY2lXhX9
2Umt1hGl98xwQ52mKNMyarvZevbfWEZrXkdpjr04+R6El5//FP5iSIxFG7ZqXNWG
r5LdJbY2KRw8Q+TQ3yE19jZ6Gt/GD/VHT6Zl3khCMAKdFUnU7iFXwJu5vwYCUh3F
qlpfdAyAp/ne1BPXAkG2E369/g6Gxngak8tbSjqmAv246UrBZAYfgx5/eEIGRZh4
VJ3Q4QLEPQfS81tor5D5NIhUlf0v2kWrSaE3QXPjnQPlKxQuthGuUvGyNNOpxj63
+U+6jOTkNQVlXEP9fkNh4QWzLdnkZDtpuqBpuOw9wbM60CrPHSB5KpyAtSI5LXgb
sa7iiRpxlwXSWvtovXaJiz8epirI98L9twWtjFA0IcdbgSMpIBa8DxBugqMsHCYQ
lEd2Q2Pd7OhzNb3ta7AKsQIX1JSSrAJLSkWuqGHidrFgUZqwWSyY2WzEfYF2934u
phRtoxwWxCQTVS0Y1g0JQQTeo5z2PLzOO7asWxP8afdvqqydszp59fU21+JcVHRO
8ebOEAwtxCp+AcyuggLatepEueYzdrBUlogGf1dcAbRWK+jgkRQUNKnXpJ19OOI2
DEIJedt6V8xl8AD2KSNh9YkRqUL3FJMvgM+2Qnu+lWAg91M4hap68FyFMFsgkIrh
WIkSlAOTstwxcKQmvu+K57LE7lt6atKyq8hwr53hddLlMrdGXz5WtiVx2pkTeA8U
KBiNMvP6UrD/mUrgl8S8RD5BGVKzZC6HnLgh6WA4+f8FcY0TFV4IMDudideoFXXW
Ugha5NjkiIt4ug0IznTbq2p34PAGSaxgTndDnJrQ6dQ28nzOKhw0/muzHmRxFXNj
EF7cKtf5f793OaxonxPDGHLOEARohTJXrK7PlM4SezFJWCalUF5QbigMSxA7ex+/
FbR3euscTE7wnOxiY+IceXS43BchVGRmwDP9aC9C6JkloLpw594jXlnFmO2YMy0O
piQBl0jsfeFVs7J5v4HSq3x0+p79+vVRVKNX73+yxw09TMl60wNK+0aOwCEwOkJc
KcYbfbHiRULSaQ5TfZBxSCDij0wvGve/EVBgNQPErvw7UecVhpbt/YdItqH+S17h
oM0FOF0b2GI83vN6gsOoc+uLYsO7yYu0ERTlYuEE7V82iG3IyKSNgxyQJNx8N1WK
138AU0UvvAO8ftEGpMfjF+F6ulD7/bbXWzI7Wnj+Azj4Xqn31sa8Jp9hhMOXNpV5
4pVFxO9Zzn89wY2kzO8GV2OnSsTWXTnVY/Svvk/YsddOMJNxlZwjYHDdW1wEXnmb
2NDZ3UIA2dhD10juaeoti7Y5fmDsThuGEhAk4KxrpAzCdj0ACx6tWpjTY2vNaOMq
5vWLsw7PMfW3b/0x5bnC/VU+7amNm7XV38YeOdB2nYVKg6CpmtUd4H1Pc3HbkgbH
HngftbU+hIk22dfT6kERJXc62BTuvp2M5Y2LaR2FU50OHw4TUmq6/y4kzmr+8Rch
ObOyWXAD+Z0SeOnb0t834kNt/EL6yMDYXULO9QLsyq0WlT6IS8zYfimtesR37jiB
+uPMYuvXJw90E1Hc0kMcJtcmkbA7hVvIFj6hA1w7JXHis+7/Ewzo3y1ScjuQkzi0
AH+F7NYSSi90vfln6UfdhGRg2o+zutKVKUIibvxJFIdhY6s9K5CAHTxBm3tzQ+7D
qEKtPRMuVLNJTaVAiUxwoFh7iHZ1E8EITSw+wTen/NXL2K26FEM7AAYl1iRkycJp
L4mqJKk5taEaYOoevC8D6nBNJFI5uWVEssV7vyWc0uU+0O16MrgHfdktql8f/HST
UnDLqPwe0TUrpgtRxzcKe6FROeu369nB8tBiM5dJcnMx7nMQSsUAH1OE8Cy6Fdtq
73WD/kptCr8WP/hI/JQbmqfuGYHmO4Aqu0FWF2y4aqHv0XM+nJbBiNvXdp5RjOAa
lQZp2DBP50KICNJPuTM//scm05aelDy98DG7CxJ8UUVm/H2qqKoWmEntgr4uO8M6
jcWS+0oXy3yoQX132966GdAjwc4VHC3e752E1m4Q/mivF+lTzjPCIe/1kYcpBHLZ
tkQrNEXaQxsiKVY9YrkM0g1YRxCX3nH9QFz1u1Ft1i2J9bKSMZatwFMkrqSPsVzz
xjq+a5Am5JwwlNEkDw6sDLzpxEfKZ20GsRKSw0kU8aw2Sbhbox3LT7GpA21AS2OE
r0vVNaY9axXXuecSitIu+ELhkze6irDb1p7si/Kl92SO9YBZPgSupUmFKDezC5ZW
oij5ob3xbmxo5erqMAiuc1LH5YmxVQNqhRTNcLHAhkYdVXCCjDg4vCOkaEFkXuWv
/ilxmGlInreeuyt9UfQiXWIumZKPJ7WcJFZxldtQZwoZUDL7clX/w27MH39lD2RJ
NH7EAaSGdGM5kmT6O2h9PWHu8AUqWYnSHW2rebDE6s4Q8hgLgxG4WJbBZAFhVxKN
LKY2y+FJiI7l1sHgF2CkXW6+0TGsV6bM5J6MJFhYBHbm4SjCJGO9CJkQ/Qh8tZsF
3fDFNJUOt55CAclnqyMjAzSly9Z6TzHWNR/MxcnSOXNFVkHNsh6Vt2uKFGCufaHO
xI3vmDYLmaTbBlXtW4SW8W8cTU1nMHq3iNlXIiaFIZ59h80HZHZXoxVd4ZiaQYVg
TK/JUU9trdwt5mKtiIE6sP12lp6u7lQpTq51i0r47HcaDjKdM1rWMvdmdhNT2WLG
tCljP4l2O4OhA128a5AJfNmJqb1JL16PtxzwVAhbo4LmwQ96D5jd43nLNtdQXCtL
zD/mdCErwLPdQdCsUXh+Aa8k5kqlCUpLPQZ1vpIcFqejKAvfl0GjR3Q+TD3A8QHK
NsZDSdgDuV0sPvO1IR0gG7GpnMEv7XeS3ll38qB/zPvIgra+8zbj7Maug2va1kWS
bR7F+Zua1MCejs0dG1dK8mpJviqa1Rb6Cwu0ZlgRZwyha7AngNlCtmgxtRgQfx6V
Do5Nlh41MLn1yFicEnUt2jrWoTbDv3fPBxCESXKYGJyWj2GPIS0GzlKQtCK48p3f
OsaOYNxUL+6OOLMCcxz3nt31HqrXmZDDdr9/EvYs/ed13dt61wnX07uHXw4rp28H
+4T0eaS5gsrY2+Z/AWPDrIDzEmSppPLca491HjSV0G8doJuoyhrdY4qHg7R4CwgV
YBBaMptuROAkMBnkWB84cklctGRu/msWdB59MT+Ty/h3FqJNK+6DwGF0QJGIc8t4
6RgJnFesmWRNTp3Z82HnI65UimJg/VYyu66PsWKlX+4N8vE8+FbX3DkV+6cdZveG
aP2RbybmagShwxGtRDSOzW/q8ALbF+6nDdo02LSoBeiVQndjXm+5AvPI1uGtQZQa
KAtlQ+SBR1Hi/hJ3DGcxhsdjXsBjqRvsLuRd+WjmLbSSuvtAag7W+YYJGsM3xYY8
pwIlNQe6o2nRXCRJ3i2z5sr8wG+TK0wz4F8PiNcc4AxfZFpgn/DRJ2usV58PFxvm
0U7vBpt6lsagsz7S9gVpe6ZJFQ7VCeOvgdhELd/XIsgCmeglSaObKYjpcMmfF5Xf
6HnvAaawNlg+Cwby07Et7FHRJFM2Xs9tumrnFe9ZB6cVBh3Pesmn5UNb1198ih4a
eSLpZGKDHfbCxCBMCxHaVgjltJ5xj/uQp61ZqKqYrU8lGFCzIhME4wQH0lRSg9dx
HA/lvmLa/YFSw14aMuGGoRoSG8El2BKncWelij/tvSP0gDdOSRrflal02LCO/j02
5avvsplQZ1WTO8xx6BAhsMBGuTbetR41wSFjWwu2xHoMHfJyMzlUSQWRKWWh6BDv
U/YKQhXlnCcLl9PnX/ldQVlSUEjI8L5d9x5ptDgtDkVHwT8yTC0NMJFt49TKYcGB
FNp6v5+12RdJOLuceWMuQAfK9nWZoGZjpO97l/r3U1Ojzg9X00C0BEDaB+8WMEdE
j6WwVNo7v210ZQSxL9qwzEv+J/PB/33BN4xDvYT0kI16eWrY/vMEhV7zmZn6Cn3O
c4WjQjR1lTCYx0aLeOvrnhFQIcJY1ap56qUdrjRYdQHr1zpIMPIW4sQ8JEq7Eydg
lbNn/1BPXIJ6VPSmjYhbT68PD5UvsscUZlZjVK0cydyS+1p2FsX/7q9iTVuEjnSu
009cZ3/XYH/aImrdjXTIvXmWOQA8L1FYYdtK2KxAMNHvMUmIHh9PjmGDRBAjZhI6
G/t2qdZqe9Zsqf4bCDzeigQJhTxJ8vmshUOVlWwbb/iVyHbnGQQIIAQpG7UVFqzW
DfBzBpAn/zMnxClBg7CF51RvONn/d3IlyyN3aPo8uSqzOlaCQk7DsjDUhztygVLx
SKpNU9Vl/DEB25GdBfM6e/f5SZopdgQl5s7NIaECiShlTuyZkt7E/nuQlzq503iz
t01knmYLQKNfPkGi3wQfEB1Zx5OrpjKCikDAxg2/ZWnein0EaP/uEnc6AUJF4xb9
x9DFm9gS1D70DCdqKtiIyQfCxfYbLZmJFPyfgWp0nTCxomT5SncXRgr7DouOdN+F
dAEYfcV3TE4gBmz3dfdjyVvbVAvhbgzOF3vjtvC1H96faMyzmC2NO5uYuUzIAj1B
NykayzB+l7CdKwkAgghzT/JKehPqSJvcAxsckCtH00NwvSguw5Y6kAplam6Gu/qe
vy8DekGijk5JdQvR+9jAYaCk0+BNfTaoxfYilu/6f0cLP1/WpUHuFCbqyXB9z4Rv
kcTxz7OVAF4Mf9VnccjHrpH6OOpyGN27n/2TNNNEQk0icm5tbe8XVdm2BuA/C46W
2yzVeWk1eclRH+elN8BiNM5NB+MuD6KT74ujFzTe6fYgnrMQAEnuumFOLQTqovJL
+braSO3DA1mqdW5G8+k3oXwTJDXfqUUHWKYugOtcMcMv77PmqtNm0OXA/ShQ7E3Q
n6CtWUwUFKe3aM615i48/Wb6KjFkbMA2qXdjhONTvSOboBT+en9wJgvs06yj5jbP
/YrvYKs7CeYlblQZjC6OTO3/R4f3Su63F+NcB4bjOnBj23z2pwgCF1xhaKvNwv7B
V3bRIY7H9sUEM68b66ic28U+MRaeCzbC4SbrhVO4NmQhfDhv2XhggdT1IdYcsEEK
Ixos7OOEg1x1IEMh9jRbIoXqRHRTU/Brd9lKj0nVAMgP+Jjsx6Z2imzijZWDnhp7
T9rBzyX0hxxPn3VcE6jpTfW151jF5DXTOBWpMXx83vS/SUJmF8gYSaiIPLe4farI
BkzDlQ2E+u4SPl8Z8+di/U3VvPo4hER9R3BRkUmComczN7I3JUyJrE8YRwm42tl8
celfrbJYKVW7zRp+GvpIvtTu0VD5GUCp05heD3uUNjJEx3mHQKPgzHiaXBE66M20
VMM8BC54qChKKuQ7kUZY2Sjo6YkwzgTjARH+egqXm4IiKV3GcavkgnurCz2zxRN6
u3xZp9MbUU0xlmyEFrrCOWo8D+EGF/s870qEe27wnSTCgKBWeOBArE8jMWe6XTTC
hvPcXuSDaX/mux3xb3jlstXYsq+mmOaoZ24vz4o9UGwDICUYzi9vUP2OidrX3uns
IO/y8sgDPLNTcVPJPQL0UzvusSk/Xx1wqr2I2BqN4smQ+jAw1zG0JC/gS+Uv1g8V
KJNDb2Ra4kNDKi7FioSy+IUnDQzqwvSK3tllN+pC75+uos6jiH0IB1iliEv1UdE4
8bKgp3OxPdWAeg79LwD5MDHT5dH1s9oC+IKIGja0FTvOPh9wxVG1wndPICUA4xNS
FrBImtRhBFiOB2J/2JTNh6pIaG/0fY7qvA6fyvJUkJKIvakHxbBAN3+0vtscsAoL
m2AiNqiB9NPHKABRozzpyTd13CBdVBVrhdEMccAp6m1ER9JKzcN5c47JtGT4vOTC
0qnN4hNYXgZJ4QqyyHsOtq+RdmXnYGd7D408RAVZ+ytKVngyoSASr82P2b8FA6ND
e7MuqVXstTXLcupKYkxExi1h/Qm26l4oXa2P3dHyCJ5f//GtyUkV5JZ6SHB7zeYr
cE6q27ZjI8mofoNG7tqDQKi91NTH0zmt2FlvJ5bFP1xMHSOorfT3U0YfaXIE7zrm
qUkGd30oqpP5gwcAkP+O9l/IOM9P5CzqOx5Ie0klv3XUbmulqs6+GgXls25JELgI
kz06vRbgZ9vyJlU6DSrax8rHr4eoq3z/iH3G1R030WcNfsDgLVea/knLFM5N95sn
5RUMT3b+QHBlYVeULENqqo8OoDtmBtEiNHpB7gL2zWJ+6bESsl1EZD74guyDk8Fm
rQVkHBt+knWPPYcKXETycWM0mLvwCv1n7HaVRE/swGyFW9p+Kp20oVI3IfuF27eX
9fEX09/W4yP4DoBXAk6Da2Mfz+2HvvyfbpVI0/lmncP8ofzznkUIu5Oq1POrwFfM
cRw/N7EOQUhMzgiDzHQULPgvbRVwFCs5eNrv9JNcTJotPN6SAbN4BoL3wI4/1g7H
eAcUGKOgtchHgZWDcucC4TwF3scl72Pnb/yEtwAb/UC239zOn56RKTSGMVSdCGlm
4FFE+m2vzZ3XsLBlyt39s5dWxqhguQR9iWirdE9BA3GEEgoFjLAfsL1dyP4S6uPn
86h/wKoVzZxpZmkAxQJMWMITERMhnBCivOje7zAV2sudAYNmzB12PQH9QEzIZ76l
exjPSaRMmP/mqFUwlhQa2QGlpeoTXPa5ryFV/kHGLvMJ5ssTUIofL6nrd7nfK1pm
RvMoo/4+fdhk3AFl3ch/7y5i/fSAy4WMno990EPnsHc1DEdIwE9yy/wgSepLhvAq
2HTNRpdKBSIxVfD8lIz/OphAvOr2ei+vHxrvW+2qy/i76SvpBOPYqo9xGro/GxwW
AsYUktuPjkicy/2R+q6/ZGwmaJ3+sIWZpQNqEt5gOxMac6BzsaNxBLPkE1DLl8Ks
4YLUOfiPH6cdvksvDuX7MCj+8lb5bVtFbfs1LiOqk5UjcdFjf3dBN6/Hvgjy9ZGV
p2Fai2j5oPpnESFHWDEsPrj7T/ym5i5FyC0B3WAmCEWCj55SWBNedwT1UOozBfx3
BmpI5QR5fq2uyNyuW1mjthpxGPLva0bkjhUagdlOLBxsAEcDkKnnDYuZr2mreOPO
5CQc/tDLyEGetn7paQO6g/erItgxk+8aix03VBVPa3t2ibuszfZqp+bbR9bUZljR
LPfGD8zYvSrGh8RQZx91GTUJXXddXUSrK7jt9bssozKBFqffMgn4vyCUxwR8UAwY
XtO5Df65/mJoLkbslS7/mIbyvL4piK2bRw0ctKIhuzHojieo6AG9St9Px70AkhHf
nlT5KIUZdSIcYCmWK/YsrntEOFeUAuzuPAf7bHCbpOB1LMGT/NSnLN5qsnBBh+/n
s2o3ancG4jvpqdFDfxw8r57qESMozs75wX6Jvw/ct5eO5cqfAWRq1R/UTEEVjeDk
QEJseNA4spn1Yo6sB82r3ZH/Rz5nMKllOvTALzeAwibA2A1wz8LiIj9LqjGL+H7v
7WlIX0JegcVqIR4eYzp0BvPhRgz1RXPovnxEK7ivd+XOa1cI1mpqemezL9vphFgg
+K+v8WROkzZbwvgi6QFKJBue6cx9lv5gNEIsFU6u1i4WSE7O1cdGoE7PhywW61EW
JAZemEoF6TLIh0aOQX56vD8xi9XO5OMZvJHG6OEUTuEEMMGG724UBYwUTPnhqc3q
4NSFQqgpd6vUlm1EODsKKuTVNxNmMJ9O3tELiWWWs4SLBF/MUuIpGorHxl2YSAim
56tZV2JV/hh80Wf7KeFxeUXMbiXy3oqwer7tdSITosWNiA/fXtqyimjOzG/OP1nG
HBKpi030MAaLk7aCl+sasTucWLxSUn+bQZw3SA1VhcvN25UmxV7ZpfYY0nEVI+fD
2rsMXTHL/hmpuZFKDBIOrwz62MdSR+UOnkCtsf14sFxBZ/cOXPo+SDenDKMbWxt2
8Ru3AfBziZv+v6JrrryIz1FaA9q3I9qF99LTpewypo0aKj0xjHrm3xv2AUZrXUY7
MBxvHKGKbWXyZVt4Elw76NdMlLEXQWMcFDQOKLog+COuZ7oXjYKaIg59dEvNtuFB
O6myy/kmYSgmMBnozs8he559HSvFcAEio1i8OCwaMGed68xtbSF/Cqcpc+TmvfpU
UPilD6O/Qw7Pinja/ejS3FW2L6+06euA1jHpmaTYCZrzPpjkluv4gsHU8r6t5PM/
BbranxiLYFf7NOjay0jyORLiD+bwiUyDf3QYa1D+jy6Hj5gJtqknGbTaDE+jlhR5
0l3T591BQcigSlJ6e+RDbAiY75JhCfgdcZrXnl0zjs9F3CGWXJTC/+TfQq0xvFlv
Um7qg8aaHrblobKjJxq/T1BaJ4cgfUitvKJ60GZ8WpI0fsSQF+2WYSuU+tSOl4Ch
RmRbuaXdeZljs5u+LTxMkZn0QbFtOMI73/SRmXzXWLQtXYtVwt9P4gXyJKbkG1BE
rYfvvtlO1HaLpnlDgGVlZ+/KOJjTKjj80OPTecOGFbmOdbG1EYpLQUoVqSC55CFw
SLX7j0Gv/DMixMuumdJa1IQBKT1WLWui9vJY3H3bYDPr8IIMYlIkg2B9KVv3X8Yk
2jNGUjoYOu1swnoHYzowIg2kOqcT6jK+PVJo4hmFSpLuqMH/afaV3/0LM0qVi6V3
17KVBb5lgQ4gt1i9PIM3c6XhxBPrn56HD/L9kBZ+mZIESA5hmos2YlE/otDt0kbx
POnfG9xsPBMGeFqVJa2Se2APcs26lySaMT/8086yhARTglePhqVyDi8nSCk4s2j3
g2Cr8Ybi3y4E4Jt23Is4HdHJuU5nmoHUV/IaIKRioivs44fkLES6gseIEBkqAnLV
bQpL1bDiVo6LDTLaU0793x6uLstUlV1VtkwIu1VfgrmCCONycjv9viWZmzFSQNH6
EU3iAI3IiCt9t5GX+Ff1bp3hfn0rpWkkJ9heysSS6NJvoa4rFCOopm3Cbn99ix0u
jodKfVPSQFEHVe7DUupfzRWmjoU6oyxsk5ScWycoMb7D5YRQRo+geYzSmCUKLh3q
Zdnmg7x+JNOOg5yKjCQYs4d/x3Ia6bjpsrOP1DDKvmOL/Fn3Y6ZA1ZETW7U+Umq/
X5yYXZVHJliTvzk9iR/MwT3/bSkwPMRTRXwYG+66OmEYVu7DdBIc+BKCkSNHLhzM
PTqKg8avOjt4eQX18R8p5R5C7Lwy57LRKDYy2hcM2XEJqrkf235TjuE/ymS2FK2l
g/J7LIDtgoHfFevs41a791r/dN1EnVaNG9htbJU10MrNiwVeHf9a5GNeX7cQvmvC
VBnjzecR4Dx6E4cRkfwnL2lTup6YRjt3XALPx4yQHcp8+UY/qf66q2+LyxysbzVm
6mKa4FMUWVGPPoQrmeqAUDSMJX9EAGxhfZe51Qis6xBy3ah7b8gsXABzdLVlGfdD
S1V/FzUxXZXOKsSqYZp72wmr3BYrJg5mtrjKqt7vFpi34ChlI339CEBxqwxOSYzO
JkyYmJCoLpS31AjldNVRh/z4hiyvGajsvE359Q+heigbMCpLSRTyEPTPelWB7PUS
Yh4gkAb4RjiAjggVeJohD6iRtP3JeG4noX3E23nNEZk0yI+wI3d5OycEvl0qsbI/
H8+Mau3PYBE0UPb1Us5+9QIQIofzVe/Q9Q/pLZrtiy7Af1LG320c9gEnIL61K39f
hVSaogKKzvZt7Lr1NsLDDjSxETN7fClccWNtQRAd+g1BPhYfOpMnnXdkuV9PYRnG
VCFRkEot7bYx7gccyX0w0/5x1Bwp4N8beSLbSJtiEkh3fA7Wbx8DvXaFQbLcc3jO
V9sUlifXND8+viz/UmrSeO4SSrnvQxNxOA8PsTFxBQQjky3T3REzw9DLiEDOtJ5y
Zht624mmFe3F8OciiykQ4fzjAf4risW7Dld3YLEIGv07CMM72INgmf/TCLRp6aJm
KMAzqC9PzCBQ2CSfm+gVTN1BsBscAU0IV1kdn605l1km7HVXvgBBF8l9J/DkYFtd
YCgwaLqNuqIfQEez4xmhRz4VsC6F30TIcVzPf74K2o09sbl8FPljsrZT7maLcVmW
3plD/+bXB76nW2Wmy1cXBHdCaLzvu5eDPGSkxch0tDFvo4VHWS4kYmv7Huul5REW
OtCmp47GMxb9Rll/lkHsNRh011ohVhwqSU4GvZaZBd4Ix/8Kiuc1hlORubjFgnR1
v8TibIqy50g8VEIzOtcgsZYpo1UhCTlnaJRJofHESKyGy9hTSSMd7Tp7dpDQ2Hw1
q6beIXxNMbo2mwZ/NIbBaOpbvydawKvWuvaWTmGepAStZdatsbZ8VmX9pqelId4y
In+Rxf2c3Kj0aYUBcviJKrlv9lPoCbZ5ZQBsEoaXP6WGE4QxwMqU3HTgIYmi5sFq
MIwjOfvVIsEVPormlB+LdEuQKAJUM0w8fSykRETPQnDQMAv0Q45M7DauOeezoAnq
OfTy/1Dy9BqlfYqqglHpb/fNH6PNFuJmsLkmGpehrFHPmJX3KcB7m7qlczq7Ez69
vTInTkppETGxiFe+THtVUu21V22k3CmZ687QgvykFwsD8ix2RasWdUyfCv/GK1Yo
VgtdCPEMOE1+cRv5yghqQYhqNHxrkI7quylAOwR4wZGB9YTfPskwstLsQfhH3htd
mkerplQaKKW8aen5Z3k3bBpFK8xd6bPsfuA3+u/UsJEJhsH3ZEfBG2v2HB847/0Y
PKXg42CDhilAiKNWck7lz2diskcOBoObdLgyocli74brMLIVIsEuYfaJMsTqUycr
oOsRQpt+ROc5JNXH/FAqPwrdrT3YzLYmmwo3OvE/ZlMPPKeNeF8bpHLNFCC6nT0a
ulr61mKMHV5jWIpsEGIuEO9WCodP1MoXbtKVaSqR/AI/tfEdXypfEby0qp+Q+/3E
jpkvAJsrOuaOBzgyApEp8//7cSAocuJJCmHAQjD4fzEBhYgwovxd6NZ+mcyMWdXu
hvFJtBuoOA3YEFj+0SqACYE0Hit74flsyUvKGrcQLqL2tKntoqOYhFHByLAEpSx0
eEGNIwCCVoM9pq8PFkIa058IFqrhH/wYpLOvP1CySSiaq7/vpTZ8xSsnYfJTvi2O
2gsFcMu2rdFJkS5b/9SmvqUZ1iIYMyeFustnUECvTniP3wo7DAtqTjosGdZhVAQu
OipI6vlHxqKoDyMN8Bcb5C8IHFvcV80AfVOYlqNktAlT+LpdIl3qVZjqDuW1LYr9
EYv7zhpFrNPswYATzS6R2J7wBKOQu1a7FQaheRSG1WyeGYOjsxAlPzIZ9J83HV+G
Xqyb4aVslSoR0JmXy9yskHnQEraCRxATGcUgJpjuZBr7jtpPeiuhxEBt8KOukAyf
1Y5iyS9ciKPU/pNlSOa2JOhPDgeJUCwAsB4a7exXs0ZY07LNW+WpEpERz+/VZ3EP
32oAlFneopnsUOnZoLaT5Hv10ZDvkshQXDdaMFzvBwkynJ4/EyZK/e5dY3ubXy9e
C38sITugjCU1BPIq+8HdrOwUgjNh0hxzZhXVqpWzfwTh34RVZY3ivTLs9W/0w/5S
NulSi26AbIFC7UasGMprNh7phvrgAMJzeiv9uJ0mxAhLgEztTQfHynqkKxSnlRgz
gODb7BamxNyQQ3MxRPM3IGLXeTy6E+tDTxCaO1mhjHZ/gFdJwmO7uTEpvnBAdm/o
yWEBTWtK6g5cAqke0ff6WrC8q5Grjs4sFVUP3Ycqu7dlpUDs4NzycrGfReLWDK/D
n8sCXmvsrTN+us2iNaAaTy3QbR7LzObiB0wlUVlTZ8mLrdsPHQ+DZMALUGpndLd7
vhJSd07BkKzVrppScwLYaR9nqm1uvh4qxWwesv4Vj3xx8idHZ8t7SqR7mdXPfBhb
jiEerE/dXncTDkP4Q3/R+Nly5gWQKhnwnlEDaArFFuo94UxqKwu3p6724ZDN3uH/
PiBm7mauwamRhgv/YTK2vHQ5X5TR7Mbb4NEJ+GQa6mz0CwbW5Ivo8BHjUQXhU1hd
9VC8UGzuxUln/1n/BzwXI2wO1eZJtXwVxoQDm921Y2YMmfx66+JeidoiabQ3zKVA
70q5IiqOjSB1xsKMhuvvWeVDzY+cv8TPkxgePWc/J4cvBW06u9hAcbbY+U2XPjKT
zcHNLbJ8IiyBYjM/qwYNoWrNrcd9CcHWm4cHNz9C84XHqvlSZyPvLjuWwRUWoSxg
CDMP/k0epT8N5S0g2NoEgcHvqa6rYKkNNVgM6mvFjhhOfhs+8le7d5VRCi5hVh4I
pPuTDFC+4OjAW5vw01eqt3852P+HHi5wz6TcINJv3Wguo7DZCnUWrwVjelLzVjul
JnlnLevPUlzggerTGxIbuBnDwQUHFZ2K/NvIC1BYT55uRJpKrHFT39lnIzIHEPJt
HgqDj8N/9n4SK/sFvwxcgqePFR7KTXKA56iMFmeSfFNcqC/Hemzi5UQUior6zWEC
X1cR6rA8SIDtRBzqhwNO6iIg4RKdJ/14FmuhNvkULETaW+wU2oszFGGrNu/bPvEB
Qvbxnmr+gBickmc2k0YpoZAOUAr+SNxFTCRG5ufRoqMQQAMuzdOEoqE6w4OaMqsi
Gg+xR/9YWXbUlExUq0TfNxc8KgFttZ9MIOI9PJtGXSpRa66DbnPS9b9c64JKbi35
lKMDl967SnoAm9xrYZibRIE6c/NqbLJx2fD95slza41QRovV91iYMMqqCAMlNluj
UCTkjsdnQHUQzkuGF+uNqOM+w86RXxtch6dFudAC1gcyRR1EBDmytKz7PP1DkpLs
sCmnTuL6wT1vfgi6W9lQ20kZLwMTIMgx6CclMu6gBhCaL+klizFg4E5QANMI+fwg
vHhL1TjHWCrJ+Q0ee6JiSg95KVOiYt/Tkz4p46hon2BDDPaLroXeRnpsmqDD5Npe
bocxIef0LbVK5bQ4l+Ebw3QFpIYLnhNSgD6+l52z4XV64rBFimYGYTzKmTFUN/Uc
dv+IEpqtWpFm+uFSyFqPgz6Qx/DHOr0SOP3Y6vUHjDgcpZZ3BQDl7qnsS8W8zKD6
Tsz1MJKlvwutVi209w5Fk4uxfzmm8yGt1JI6hY2mh76chrrW+9S+8z2UJUBKs3Zi
7X67OQViJxRnbStAzwdqFVreWt1xJS/0TdIUQ287GPXkMsOJsxDpXWHyRGya4yP8
22SBH90QvTvLkl8OaMF/no3n+SVIrBNDql5UJy43hM2tdQdrI+pIkPU3n1u0FWaN
I4h8HNUf1GxRfEso6U0i1lpVXUYdwvgUHmQy9RAl5MPq7FwEcPwHH+R7S8KQKpIW
vm2vIntl4YrdMubiF3zrqWxoaQ2MQiPkXuaA6aBkVs8NxBRWbdaBXWoUtGpIaLiv
mynZxpNXTmxSnw/mSmwD/oKb4zElxNLeSXAThHqZ2Fi/ycrRcRGJ2tbJLSr1lBL2
rP7TNs62MkR2CeuHqyjuz96Z7Pp3Oe//hXGt/s76Q/3tJSjJHEvtpDX6cRJJWFGW
jXZsNYKPUqx7C6xwsRYPfFJS5QnZkVVsd1ULRP/A6XTQNvvjj5smlXsKZk38IUwh
muagRmiocOU/m41HDr2rle5vsJMJ8SJQsLcG6oL04iDhKS49+zOcIDdQB9BdKW3r
gu7HIrijdwS9LzSnMkzlfHNTjz6g223tgEm9rm3PYABoI3+MMb/pFl86yvA2n/2N
BFud9BveZvlZqFQbp2RvSoBhMX1EKCIXk4VUwCV4blNBgWA+FyA78anOavSEV+9Q
hYZJddJfJAhJcXSvv2Mm2C54Hddxh2oZmxYM7IQITbfOix9IRY41JbdlJQwx5rBX
u4tQqwqopG9k70kyVJsCOfkdurBDb1vi40/vxRNOJTHl2xbumzgaSljA+Z7EHlCa
gsf368w7szcWFn2A3089w7+Xd3yTkFBaSqguM72aXhkhf61RtAlFev2iwfhIMgJR
IF+j/mMfB/1tfgVFpIPFpWstwx/5O+MWy3WaEOTi/y3orrf39gigFU8ImqnxJeqr
P0CWz0KIHE+L7zuhBER77RIBF6T4ipkrkaajcdqtqwhO0a+7DXItqnFG66wDYENb
KiyJ47Qqm9TMNd3IXJ5da9RdWuEE1CGoLLqE06827veVwj9StcK3uDdhrcCJCtyR
yOOewlkm9l/cU27iNXJ82UTuoDOtjFvnfCAfWpEDVrjlZvLLVtg+xbXtrLibRUX+
n5Fn9GPvSdxycFKPOe0POvnA4R32nVRJr+6LjUhjuI1iJSymfQsN0rFPOXo5Nbdh
iOu7GRVJUFgRBRacTczmGFoMftxtSmVy4OycXaI3ricviSsBChjVsmY4IMDjxqHs
N+4zoMsnRrraWoIlCASNhRMgSZpdy0toziBvxpUq5CWKzBJTTch/80W9nAQV9GRA
1I9Ef9Xxtml2vCacvKryaK/Tn/RQlCic5PuxRlosJcL+HtsaYxLEifBS/coTnB4P
4j1rP2hg6oOIls6cZaPPFxzGAZm3N20bDv7StSQiaJQO0H5nzl6yWohLmoKEpmJW
4eD0rXj8qZGyR/WA+xby6ADKurMSJZP5viu5r/EYteVY9VAMUeKsUPav+PLXmCdf
vEyrmKKFGnUt/UasehTY343/n5ZC1oyzeU1XTkWXPUvJy0tDpj/CJxxRmsPxKWhO
NhclIIAc0VzdnzSgdbubqGs8d+TRt2l0BQsxl6CNo819fxtKVZC9aVK/ZyqxCzy4
PYnAGWnCwyayQNzEHSs09KmpJSXhahURi8fRD3gJ48/uCzOq9maxakHfIeKzrCru
Lav7JgQsiMKX7NK2PpkUUL0ip9dbS0Tfxl09e3+lfn33XzhmKFpUnFp+laILj/3V
BOJxdZHNrOyZIcBJWtwfpNxKrVDKnuAjG9j846BtMzMgCfnR4/77GhHoQmGL7DEk
hNhFyOe7DsGm/TGl7oe7vcRmhmpU22WGK8JnEUqqNhICHvGnSgMXm13YV2zj4xpM
J10lcwyNABrD38JV+098uYoTEbsjC26TtjUD+jShRJpIZldl1BNi30lfB4orUkP9
CrbxgDtKJAtPmG/myUZ8mPKUz7LB3xzsKNdP09GXliXS1mcEg8eAkyx95nqbrn9F
Xst6nkoVGxCxiScHM6Fg24HD0MZjKWC6nsIG6n4MZV3feXVfd6kqarmAwcFyoo0D
DdmNa41M8WlAZUJiHf6H/dtl5DJ9tDK6KhQZoXNYoRaoax/qc+IcUEd7WQgfWUuw
lyZ97sREQMO/9vP6fonFajvaZ+NEPYQt3ukpKOQdMwZjKIWk85+kHvln1xnZgujX
xfnWIgmmoMbEILM4bg2Qy1h/AbJ/H5+ELg/WLhM6O1jnCvDUPLyaz5U1jnZRxpBp
e7ZhNcrX7LfkIt/58AoVtIcQ40jkoQoc/UIK7ZlxAM5j+5qrfRx8gU4nFVISJDah
0j4iD225/4ZD0CjrRYiTk2tzkr415eqsBj9voCTwIyFZziphiCgI6CzxTGuUog32
a4trRsIynmBdYONfjWrYIrWnlAwo4phQFoRMlYQKT86sp5UH7uRTXmibi/9UUQ1e
+4kz/++PDItgIPIW7gw4HYEtQ4/ZXpkoa1tpz9cEosWr/nNA4Jx5Bj7R8Na/OuXb
9LFfG4VRb81e6blus3+aXplf85owlefxTEz3Vp9bVgmfmAs9YXRpMzM5e8fjPnne
OrOnCpHmMe0Fjo+8TXsNnjOs1mRnVMR0VpCeVqR5oRrFN/8tTfjC0LYuDGuWDm88
FfBb57jEyNVZO7bVkgk9prD4meDsn8b++D6YW2KhxjYrBci1+Sby8TByhZObO7FA
i1VTZQ76hE2PTOYftzxJxkloqyuZaaq9rE+3RYuuq6WaDBCRJ7j0NmfaJTOMyK58
jd0lAhZXO3/BU0SGfzAAgPgU7Llx2MLcA+PIZZdROz7uyKa0RSvG1QqMTw63jP7G
BGTFeT1ccmPrQBHKJjuFSGSwkmqOlCv3whyU18yYIWyoUsAyVO3Hb86TOvdUGVno
srmbLG0DeDhMyzPywHpkZ/1TTawvut+h4P4/Bepz9E67Ii8cIZfBOm7CRX2/dOdK
eSyXHx4u/kBDKRMgViOnL0jnVhBMcwVPbVCvopsJFeyq8+arH10P1M8OxR9y1L2y
J31oTpkOr9LGzM8X+XRHrjf2hwfKE84JH17+05y2CTeeGpN1AsVwmvrxiNhO7UFL
o9ljYIFnbvkJ4ttBtHuiw7a7JF7+WGmvYb+k/TVmC1I2jEgfbOXHLTITzlRUIY9i
0pQQonRtxuJVsP5zbPozTt2Jqnt0+hz5zvXXGLaEMEtpUeJ9b4hTRh8FrJzXmY3H
BBEZ/UmHeAhdfMt+iOowRJCVKmdY9qIZPoLMzL/rWPMsOtJyRmLb/eveF5eM9LTQ
mtUluk9/sZfP79dAY/0UC88lQVws9WvQUNwsiotH5PrQhS6E+NxkkuIqX1BexseT
vmiB8FEzoHsr8eb8LLaKrFhiFmus+oiw9/vrGixDdZVBU/Idu/h//Wwx374BBxVw
bT3jI6iDqvQDZMU7nYGOwkLy65GUbc5a5nVl/avTFe5Kc42maXb+lweVsmMdzDlh
uPLE+l0ba6Iu8EQ5R+DwGQfvZuzZhop/gqp05vSPhuIdfvsTCimGi85aqGpXCv58
8zFtEiQV3AXHn2wbVxZC3E6wjoa7rtrcLhjJ3JNU3zYCoENTZuJEC3c+CDrJCodh
bBEiBzpXy2l6p78vbQdiKviCiB5gz/M+I6ntu/CuaAud02Tlg33axFuvHG1jupVr
sYhx5PpD8UnTB5biuZeF4x/a5FUqw6izn2y3D3MXaLDd63GaVlMHZqwvD+ZeaDNe
t8W2pJsbPRfzH4VjPBlxEtMWmSujpdcD/05GBMHVFYc5a/oIP3zICwK1QczUChsR
e+x2CYQk506gNnu2N9FHP57gCTRFoldXlcG6zTw/zvsKa2a/AEClNIgiwxZOIFjT
rYcFNRyqVTcGmH37C8JeEnsdUM8k7aPK16qXxxAKz7eRgaU8CWmrdiIulXsQ5YNF
DMlrLKvegCnzEKcQ0k5WZvqWS6Evp76j1gS6lyREnqSLPGxZuzr5+68v4PsqPusC
OEqTT9l2otlW6L9a6SuLcfiafACTHw507y+3EUQzgfVDi3qk4Hx1hMWoW7mddmd/
sEhelnkX48byaXSKxQ6wiBok81oCe+nblSy5z1d7RSD//bq4wEeKxNteiCApAu0p
GzjH/4Xpwhg0GvUoFNe8vzlQ125tC86zxEEBCDp2fR5y/PoTtS3p88gR090gHNib
6aNvAsMQ9KHMBjSY5QymziFC+E0wgQC7lMKe41JtCwP96yQOg5UV/VOQytBfaw+Q
H5/5bU2b8poqdz96ykbJRFKhXzGWoUekZovrRNtu3GDmmNCOXuI8O3aIXe4IbE04
HknFYCX2HihMBcudHd/T2kL/Q5lCMn/84jHENJkq3E2iA8YWnjGg/mrtinGShmYH
Y0VwPcXUf2p9DncgIljYheiahPRs2DPc0q8HuZXZGVXQOhYU9mu4KSIJcElTWEIA
UERO8bR2XIXvI9PTMoX3CF/G0m16dJUXTzM3pfDiBOFFLEEYYdaCs+eTk6TrJofF
Z9zY4n0+l2ZN8lWvlwolxziXMUDSm3VuCT1knqDmw7lbXG+VjQ0i8+Qm02ThUQC+
7nEpmet3MoWP/R+BxbQw84HJM5mgg+860/R3dRbXMRQWCoTPR1NCerEdzd5daak+
nI2WU2gQSulg0Ddl90rd/onjy5BbwuukIYM8qfuNXwEh7cfFMJRDcrd3F7lfav6j
6lLoQUL+wimL8OkwgLDEeXYVkjNc0jmkOPDTrd/4GU/tNzQwq69C07HKFcQwCBGy
43mK16jIchvaZJhtiEi1adZ0gmKxxjAQeESvuQWMmJ1mcLi7zbF1rurQXbdMVnuZ
niUrZ9mg0Qb/lYnYmG3e3wgYNGOLMD0U5RyGIrDYQvW2cB+8AX8oamtvb/5dqTR0
PX76Brxhb+N1m5QP+/zaKLi+zAL2X5RWMvAUosj8Jg+NI2Kra8MfuvNBb9YsN1+/
OWWeq4rz4+p5EHfatOjMWhIvuvTST+QLCQyA7CRqbfuA32cosOiUUZ4/ikdUwyBG
pFXStW6wVwELVdbiD2hhafsGQvSCzKJeX34REte4d9PzsIr5yelo91LAPgZmHr8t
h6saa1uEzK1ITlqJF1za3UOED9NCvd9MukytpG1PabkOJj7UlJhAHFN8vdhnn9du
6pUzOwOnzqFUXmBbD5rwbWsj8lWEcNAg+QS+Ua70qwRGixqepkggImtoCU2qfm3/
Kk2FDnH2AhYoTl+vSWFUnKepCv7fU6MWkZc5YswgSjKNQNTk44w6nL0a9VbwD0WG
JBmlU9Q+iweBcov+zuTM3YVrre7vE9thf8fH5N5xuDvkEgc4fE0eJJzqKhtpHqkR
lSHp+LG1yqkp4pbTVnE9KTjPGtL9QkKuqL+M2X73Z6sdUeVb6BLy6M2cQ3ZMJl/f
aKeMOBGQLrCkoXGwNeTNPgWtY0IYiJGf7n1fO16tIq3kGVAPOyVQQQYu5AKitQMD
PHgWjnoIaOlmER7JAxGBU1gAg/LQKXrYNhHU/Nverh7Pv7T7lwiiw0bEeffSPO+e
q/xDO83RIE4QovTWFZ1nVhM7E0ZuqOshEorD+XUOoEPhMWWKVCyzYNfUx/ljYCbU
+w6PqiupNDwSuIfJeLplaw+BExW/HSl0HqGIv76Pr8SUDRRKZ72rcLIhwk06Lh67
+3rkIG3CcsK+bcZ8aTLDO5ndUS/Qe3QV+J3xl7bLHtuVBHzW4oZHNRQPmtzfo7XH
0Q1PaEQm2WihwVZA/quNtwsRDlfQl0IRSGUJkXHwjr8GnFtryaMYjwSckI4Mmcsy
HRYAGmnTHk1Om2qwYzXi3fgATQGB1unX7BXmunMnOgaECT1AKmvbzeRmnrvB/+c6
2nJV6vdIEvqrBm0996CJXeljJzydQzCPpWymauLAYcXRc+83u1NhB0pPo1iZqMtG
zJixkGDmVlXMnFDr91t76MhSbgWb3CvkEPKz9cWr6y1gwymk3IpZdtH6FlqbGB/O
x166jYLsIuB10Blkzjc/jDmtiwaK8/ol5ykjD7eR2ldqjXekLKL2TZd//QtLbc5h
P3dv1QrAYn2koWEPBSMOkJOW33zrX3BgFEJYItlo3f0y0uj53o+tg/9+6kWIN7kg
0nYCh1wJXfgNCkSRm/nidvQLTqcRMQlB+owqPDqczEKyF13ugx6/0LM0XEh2cD3I
xMhdi/S6SGWMpT4iJbEoQuzdh8EKfQ66xnxQOaCEfjqVW+wddXxRgBzojhgnZNeq
KNb06y6O3iFpr32ibH3OU0oIBCjhXQ5fOH0NGhXpIBEG21EaZ9cjvVbBGhHiuRaA
uJNbj35XlhIVKF/stJ7NSln6+yBoQbKS5xiW0sH1ttKSexJjSx+zM09HPJKWZVVk
MXu9SE8ulJeSc8J5ALldcOl1MJyQbWuPO/H1Ncsn4OQwTugxHCvG5brOjhPYTnJ2
6PNp2bSzT6ausYlYxdmJ+hcB6XgCVCPiiSSX7rdxJ9hm8+wVSk/roSIxWrK4v4sb
IyxRUYzl6gU0QArQODBmjHmbeXtWtDLdNow6fKcpbBmzoq1zS4Bh9eD7PLpX1nAy
XZAF4AAMYqMxmD+y9d0FzSoXBPMUECYNNaP5gY4Cxs17ZMj5/4RZb+YhTH7CaNSc
1o+XVFYZqtJ3gbaR906Br3Fc8/twt7dl6A3DsGxaBruzyKGMVHmwQfT3qB/XDtsL
ZctiNxBouxcalJlPK9xRFVrho9JA/yZNIF9CQFRM3dlF/ZJCZGqrP4n/jnlUzN4r
w3Iena6mT207WMFbDBcvGZN9VGKfb1tgTnaRP6R5C3oJbJKkuh6I/JdjJBkvxvqF
VP1acFFg4dhjFR0XHzHAQvn0/FG31tpKQXyJv++WxXdfUB1wPI3XyJxOBpLxjIyS
UM1zKJKxhD7qDBOwimd1FUbYjAvljg8s0cYCds1XXotzzowKfFITC2XZSGtPDv6P
prEAP5yind3ggP7CXId5O7IIVwrV471Ejo2N79HKStlf+IbwrIg4dgb6YnkQd6+A
OoaBI0Fuk3A+Nco1PqHXgDA0HwMePvN3nl4ZoW1R7t1UXHpMIIYLg1Z4rYm4Dq5B
jfM2US2VvHyltkba4OsPig8cRxQqfBsqZSfzznVDegRtltmYTNEm6DqmLXnGTPBD
nTfixn7YvQGeCr6TfpWMBY15U6WRH69ViVQRPT52oqVNjzhokOQImXE5FeOS737c
Gc3cM/icFD0xa6qkMM8IvbQ5J5M88KRhp6Dh7wPPE5Be0Ov9aHs5o7aSB+aL16x3
udiaxztS47+4k3BLxIm8d3f8bHEcuKlNPInZ9rj4an9blZ592S4phWhPbjwC8CVz
eYoNsWUz+lZaScvxv4YX/TQ3Syjyx40HErmFydSKZVPXjnW84QAinTboEAwrSbw7
d0gcgei71SM3fGJXAkA0biI5Si7la5TgCpxgnjOJwhM/tuO/hBEiKsA3pVTlgcW0
iBQUWFxb6VNMwERpSb8e5ayTTPs2BNpdss3wrXWfh4barEgDrmbDhvc16JA9iF6V
N6LOvBjQIkakqgD+D7npGkpU4MyOf8c7JhpJBzOt07PT4GnJUBOKPCvcRTyrW+fw
yBYewe3GEX8HjQ2/qvtxxrufG9VOpOCVIacpa0iWhjdHLq1MAqpKwssvs/tZDwv5
dQU8P4xefr2xvpOCIFbAC82LwLBfmiavChZskdbEFS33oA90rjuQSu5gfO7HiatM
ok9ojjj1K19mHZhcPOPrSu5BFgD5lLTAcQZvB/Ye+oxzwTnofjHal8UmvOlI3TVt
OQFqYe6LKdJ0zNBREmsiFhxzXRnhleCU06AeSJ1x/nO7atjb7GSWRUn0kupmwiFK
mMi29aQIhTTCxJ6AMKeD5GWEyCM0jHjnepeiiVaYSfMPgpvwZbT3i3AkfmdjnILe
Zpc6VU9EUeMBvhUAk3ISeC7H82/3wDyNkJDWiOJVHOPmcgjWgVwKRz6cUBP+Kfh4
lWWXMogTBECm9H1SnaC5OuKCGnK9mgVFRRIk4YAF/y7LZ5qymF1CtuKbAYeFdPc2
uhnZFfSkXxhCfBvCFZ81wFf0bypB1BoLsfqKSsua4jP0cLJOXndXmdDvfbSrazQO
MaxhdmGoZv23v3eWCwDBIXcbE+7Ud2+PB67gwvwBfzAZriAFqz1tnMK6QgNLJbRp
rvbTSS/Ya62CSS2dZVEYsHo3wKXDMBd/WOYYgUZbZsTZmgT83OlExVxJ72hHC3sp
qy2YrJqRG4/6/XKZJwnh9mfQZFM2Xh8Fv1NBhF23wAvnbQ3du/pAztgb47y0UPga
z76xZUrI5iOuIq2nhaQf+YoODjH0ad3CrRNc8O07OmK3TCOf9vRBv4x4DTHCkaLp
jBcOCqAp7md5AU940mGFati/29dyNxeEOSpoNo+4A3WKC3wTFNKzO+xs3mjA08up
dKD7QpyJs+QX6CRKZvvjVWGmTLVvOKX4jJCgJYoUCz5Gvavmvzg+O1oLtplw4BU/
VKuGPdNj5zEoIKk61pcX6KCn05/3pVmTukpdwqGQQL5cKLjXQbMGPllXBrcLAKe6
f8BWKa2V0iPb9xQMu+9+qxs3dbDeOF9S+AIbAbVscUInTG+K/XXqi083uw4MMsvU
ytnuF+ecVErizHeQt/B8yrj/tK3M3c2iYqQVeen7I/+r77dhC+MVk734XJ0boR4I
qKND4uVFA4YtYfliqa9bmu0BBnHmQ5uYpHN+9fmza6eSZ7RuRTWBcDb/Xy97ykJC
SdT3LVuzq+6VTO5ARNzwQbQQzaVwMM3JpMNNPs3wHJWn8xdQmnATuu9WYKGhJjxj
HqzzJeAQ9Mmxl9q23zNxP3gOblcZIqD9pkJfT8cb8WabHT1Hn4g4ssBH5kBClYMq
0CnauQxnIu2175yVm53xL3Vx7qV9UTIDI+EyGOmMHVIhDObAKZlJqq+2SDiLpb/9
9jOPWr37FzfG9WE0HrKpkhG5legqi0rzvkZDIMw0Ucz8ZNcH/sdpFKIQNj64El+0
K3STz7lZrJXd96qCn9jSeWAr85+pX9tDg1EXNU6UFAwV/AynyS2wUNKDourHQW5n
g/ay/Jx1MvclRCV3OXkWY/+tFVAoCyDLlW15xiVXlnkzqW0J3+VbxMbaBdBiIAZg
qdpafFWAn/KELlm4j3mYs6qcFuP/B2ah8vg5J0bTP5JELiVmNJdxDD2KiFvdnQE1
f7S5H76D78go0LA4nIElgPXR27EKvJ3c/pcxxNVuL2UTYqDNacQMkEsFPF+0xFAS
PupXef6RAMm7jfPTwq6EHwNSiRzjViCjowkG9T/Zn3c9UNf58hlRyJtrLxq7E+Ax
VXjk172WZEsl+rzlbzLwrzGHRe3PDlvv0PAdVleF/xUGRAwRFY58mTJlIj2S3I+7
SWOYqOZr6gDoAQZ7AdPj6QT7x8tm+0YG+WrB0uyWNrdSIi1bUVUxc1a78vUJ5D1K
U78iQ2woEs9PNk9drRVpAGTgdgeM+aXeRyiIeK1DBqyZJ6iIx65q1asstZhvaTDo
RU5kV8Eqe9OtuP4MDgEyEXf5bCOU7oH3kIW3bff69Jvbn8aWXbYsrt/gK6lrd7Xf
qKliXtsYw/Cf+4V04gY9/Ylhm394B8P/iuc1tImK34HjBz3DohDe1Fzb2ki7YPGC
Xn1VXJpRMI+SPkxNM3mUGa7S7+EEpl2P9ckfjbWDdMTpNwEasamrAcPrC+ziQEJV
NlyhKcMl1+W4mqbVNs5JocD03BS5o5LrdCMs5orkmYSBqWxlGEQAfS3QT6C67vWu
7Io4JpvcdpM1caUPhn6mkC1Fal/pJR/Jx9I4mPI3z/jSducEIZSkDVBnP1Spd/p2
nwpOp9RdgqAgstcJKgtVjtYi815CusRXY6hYBCadqGpilS8flVMQE/RrtglK6UAK
HE8b5USF31Qbc4hV6rfze21n++xG4Rk577YG4Gt45l2lDZnpGZb2XqOyt6aO59PR
v2QuxZACtlbdEXNIpy+hFwkjYU7tS43d9io8LE598nRLsMZQtlwiGFEnfxuuORWV
CgoKtPFEtD4upVqSCDi89a9+WvE5sBnlo1gz6ddFvY+nGabWwvpbSrtponWHd76h
IUbDJhkyyoV7qmnZiRYmaFo5cjU7LBWOJzGl3b3FQnEXYeLNqETusf6J84LfNqAA
b+ChO2ba+BRsqt8kiXturTFA5JxhMGpcRZlrlpEFevW7RHQ3IyhdGo3WuZCnoSEw
oYHoLb3thgAU3mkrjg+M4RJhqbVmupmBZXIYbacGYtX9JLGOylE/iKrDGKDAXUnt
SRXVTagt2GQMPqTuIX1yrcY7UbXN7Hbg6ZxhdRbGY6U8RMEEhEjzt0YkwynhRW6O
76qUMaMZCgZMz7lChAil1UrW3cwAL/2M1rkIT1fHx8e42pqlTEX7FUZ1u6QLWS/c
H6pj+gq+GilWpPMh4VdSFZ2sFPuu9IgC0yDQcilY7537FHHOzocRDkebgEY0SHWr
3TA8zXKmDN+2RDfWbdXGmVUxckVS+DxcKph4MctBRwQo7A1YTtLPRxK7Zas1Mt3t
WL8WChBQeCVhgVF6axuayAn4qUy84DyCeN8vlCIjqcxer87VJjDKSMjUQHbPQC/P
qbih8ANKtt9ckJcURKwDLNwIvJPU7/f0yXCD2XzHeYJLkrwp5P+No79iRlLIniU1
jslDuzmB/zZZdXXY0B0u4KHyZfbF6u/S6gvLare5WD5ujqQal29o4YY4TeFMOehl
SdPgskjzlOePtD+wZ6f9aO0AeRqvbwQqGE66fI0FrVEgRzQA+h2Xa7QEUoZlEFge
i70r+A0voMXsqBx+OfHEq/oGyU7cqvzASN/72KfhSp54EZUZXmESCyeMOU/3hZ5o
7xVJJodT+p5pNnSsT+AoCHBv5SKFwOZSLXpNOZVGjWzSMh8m9UZV5fWEiRiKvzXM
nSXNrrQG+LOuKp4Zc/yVQFMRo2JtDnBB20SoKsddf6JGRAM5TBDkYAasnjpk6yea
ki1D35Tf6gyCxam1xRQLWUwIwyLszf/dL4gMRohQ5y5ulFNr+r53rZEoDd7751Jf
+PdDQgWmykL//L9y9F6L29++4X3H9MNdrN2BzmU0ZmhCOb6cC6qMWJPqS0TqETLO
Gp9XGMTT91dRf9Nva6vHW6rlajIDijdj3l4B+1VEe8oLKmJlB/Mq/MdFq5X6Rmih
7QBL9kPfEV4DQo+mSCybZjXMp6oRLMEsXn3vXxICmBNEycU7Mg5wAIZbh4+FHkvV
vYdp4YfrKJkFIPIdhrxy1yJ5xHcXvZVYk+tsj2Ez+26FXBnV3YzE1dE8e0IxgMK5
18nC3CHCWbYZLHS2dNRTffpd6cK3u6Dw3aUTcUEyUIe90scTNCbGOgn2HBjuzGNX
Zkt+m29Cv9UM6gtZO/mOL8YjAegD1CzZfRzxHvID7KSk0D2j3WFByM6CBFIPX7tF
SIB9QFcbEmqGY27rBh9sbRR8eyxB1WR/LX15KaQiuC5wJghEdipqMdDx09Ertzri
0HrK4KxcqY3nlgkD34O+mXJzOz3zPsSSLwT08DOisBWA2wXREnC7UYrI3hK61YzU
Cm+1W3MqLsONoMvB+w+nXaTzqM7nJa27YZZQ1Yyu18qH9FwxvTL9n1u4nx2NDmH0
FUGppul/kgDQuQogfJnZNzS874y4l43NCpcAtSaHVa4eKxu2ShMB3tzdJ5LQAOSj
Adfz2LVlFInE46ykqXm4DTWCVIVLmIZfPFHKoOrn798KrI/ThchPqoGtZdZqwuR4
klz6hTCFC1+Yo81XKO0gdvUHVTUJiYULopnJX6jmjpC449dPd82gWrpJwTQnxU+B
oTpTGv3KSuT2/gGjMZC8RMh8djhsJl+e/A9Z4x17CiKSOKfMnqKvD0jVUd7MS/s4
UI32ImZ2/Jxw9iw1IyoVM6tH51iVBcT7p5CBIteye6Y1Z1laxLsGDYuQc3HD5jSp
p4aXCurTU7yRseXuddGssc6ubH2Tj5tW0UEz2Aul/vSGIe5Thfg++XHuUqctUTOs
FZaAAvMMDhNHQv6n0m1pnCUWxFQ/Ob456esfGnkhYPAChxfTnDv12gtOBb6MdIS5
tNrd5hGF6OQgrujcm2vGhcaOWMqD6UkU50wh7IldUxf8v04tRPZTWNMdtEODATLf
wpKNm43aP9cEinvKGx4Ziw7XDblwCshT8RXRM9pW8g6M+ltmEg2X8KrlLEbKIMvo
a6xPNUlSlJXyVKCcF3YvuP1bEA7YotEG4JpkUlFf0lfvo4BAJ68vS0bjhXPBe7wL
vspzRGbedmboC2dim5JY7WUciLtT+3SVKIGhfOTCbxijpTGrunlhEpzkt5xlUW29
BFwv85Jtu2J9VM0aegsEl92QrBzTS4CGV2XCJKP+FWcdQtBAzT64kZW8i1VbbuR4
ch+hvkJp40lG3w+J59SuiYdNbDmDsZbp29fVafB3keC4k1ZMg8VyGiAQi0OzSBDI
ft21aALkwo1UJt9HqTYLg0qkiKwKQ9SKWn6noolbJsMtSH4MxdgZpEg+9fiJ5bbw
qRV9pE8/ZucH8DF5k6hroZFUyTLMeKSGqLDkGJ9lMmihU9PHmBF2xjUZ1QaiQ5KT
OWNaq7SquX394i38a/TltY/9QDSIxJxm9uJlkI1WxJo7oyO0tXGgrGE15pMmtfsz
4NMmFGbR7delkHyLypIF2SqzyyKCbhDs3d1PyuV17xx37kjGRaNyewWrG1WaBHs/
mSs93ZDK2bFuNpknahXPdu2fWZ28O6rmVqtMBo98Y75d1Ng0X2cdjUwvg9/dylMh
/o3bbawHMTgAM3JTB6HtYTDOwXGoURj1FXyZtmJQSELSwgfnIcjfYUzqN/ot7dnP
onsXmXq6JkEYxtUBKMZCjo4hgAvMP5Vh04+MlgU/fQasCyRJD/33Ff1H+QT/VSzj
xUPvpWkAOBL5pLN+ityP2o7LsawiIEI/oatlPUP6wEwAsvQTxLzXvdbyH3il2Gtl
grmWQA2Io/1a+SWe8M0izKHDTcPXNzyM9wDvy5uC5Gj09La6NiL3pJakibINrpZt
7wWhERIwpkRWforecRxiNj2HbQ8d38/uRwMdJKFhcrJwaWTjmLzJMbvNhsEOadvO
q/6Y/Q+S0oSn/FcutlQtMRPBBXZjdzxq11qPSjW1FCJfDjMkDe1lYaHI7XHVGgU2
1ZlI2RyaxKDoCJ71dMtIwUvCka1hiGySNOUFeux13xuG/K6jwtx8bdU/aw5qMzmo
VRRsxk3i0foCWmlA8r3LOvOOk//yK8EpJB1NIDIOmG3LKEa/je02xd0zu3g7V2mB
169X1NA9htgO4fS/HJVIal1sYgINyQ26yYZmZLvJeRHjPpG6RahCj63ld0PQJU1A
cnl9XuFkg1/qU/s8LtJ7I8tc7zTjNDeHH6pbNGoALMFnjhpvfIruc+6auxPBtFIH
5+Ms+5fG6rtlnzrLSMb/DnuA+BR2Lyi5u78pNbxTkl1AyM47RHhYLabZ1GDyhhoo
gGZgVlowae8p/AgYw7fniL8H10Ubi/qAOF0gEiln32tKvG27kv7MS03EzY023nzO
dairLn5Rklgt4DlT/cruizaLf57T4WFw3Gtwn4gvoOlOMuG9iqiyP1zPZ72wfJbd
2vn3x0lVWb4wJs5lalwk1MpBhr2jWv9suHqJcNEJ6QlzQF+EXYzQL08NgJ7ebmWR
pt5Gs8lKeVDbUcteQ1MIvQ0BisV56LLMNMH/ZtyUjLm8im0+9leFDl8abP3yipkJ
GU6jjBkzjTaBFDzmBJkH0bXbkPV9TqcTf9XoTuO4TbdccQay7dwLmaM8rJxKhqdz
Mqc/HPO1oOpiDO+CwoEW4T4nfsNF5qrxz/+7fi9bP7zKZENIPs7NiTLV6qcZ9o7J
yks3RlbB28VFuTLild2WD5in9uRv9H5MhvjdD0JYDZD5v1XpZ8Bf/QH5/1/gzk1f
SjweEHiTM+0MYFz/d3xJyXp5RaqqBRuLi98mpHe559aqeh3F5+UyACqQj6AV0/7X
IW+UdLVGoKAnXU9yrn5g/YrbOO+EVzg6wQjuh8KUGjxGshb1Aa3SrBvHOzb5EWFq
3Tuee0Bu13p240LMEEFbDrsEMc1Z/ESX5XDaiYRBKcMo37c+RyrsKvd7zsiryaOd
e57aL8CJbNjEq136MBuH9+iwY1oX1RNJSAVM0wVSjjjh1bANNErFrka4SJs5p06k
n3yz1qaUaA8sPvWjxF8wnDLW1JwmblKzxkIHrGJmGzU+4YCrSOYG42tWugtlrzu8
SLmW5RBr9FtSDSgG7RIWNu6/GtQD30BX+LWI8VeMwG58ElU0FEW9RazyrwnuwYm4
YtYFzG5n3qoCGRcJfoenVKytI1D6TXPTRYGFp+R2sFYMA3QxEJ7U/WI1DbPg0kV1
7vVOxxyA8Gp5KncqsrCuA1Nc8C3J6+SSu98WksnijN4TgOPwL98zRYpRuX8Vtefm
h5HanlqdAYnWawsR57em41IygkQAjb9j1o8E8uSeujw82AlGkGT0GlhX7Qif6bqr
Kt4701KTvfNw4Q8wPKvHbOmV7NFIQBh/V4b/aTtCbDy4KMaB/CfXt3xBxiHI+0RU
zlPwSnMpXqJRKBQziVkqikjWwv3qOKvOmo2OJ8IHzjcecwvr5mTsEWnDgUl4eLw8
GM/LL/7+ZYzfZ66tL1hIIsiGXmTl6JCHusRWtonQGTtLLjQEMlz6WrBS5FEfxdEI
03PzBcXkc0tUCRgo7KgLHFx6HAj9gGwBUsdJpd+U96JiQGWMExdD20jK7O1LugoU
UlRjXnLWJVV0akbstT7DI748aQkMvTZPsW2mMdaO0db6Gk4vLJjhyIx0NjF4iEeA
lcLjbxPW25mjTRnXAgQFckWUOhkCtwBCTWu8J5t+gXp7szAr+pyMX2oml76lBh9z
3q+KTzznb6Aj8mZh7qUEBgYWp76cxb3WAVxQExvt3V7CZ3q6SkpCdljsXvhWGWjz
RECJcwyD1/Kl5BAYDbnv1722IpwNvVaOO/7VYeA9gyuzpYuwGCzgjSnePLO9BNIg
ZbE33rc359UTPOTLMSUzZbO6pBVdX+MZY7eV5EcGY22MEcJzQvOLL4O+XqqBKUtF
GJVSVNXLfbGRxW5ByhIxsB2khTuMF2ktVONvmbZf/cSIBzc4CpIuDPh6u+Nfe99r
Bkd6kNK+DTnfltgjDzdNLRGIMfHZf8m9phohDGQZEC6uUNb97ts96T+jiS/3bDJ7
1Cj6iD6A38GGnH7Q9F48al4m4DtQMWUa5OcDoqoc2fbwfDBEAdeq8HWyFMojmZEl
ZYJaza3tATrz6bTlSNUpwRaZ9O7Wn0KuIgfWZnO957rGElo63gKwnNU3DFdHrSRk
6mEuxMdhQxducDbj3HgEffDWTmPC/m4YfwYjIRLpgIsSo3B3Dl+16WtWUmqNbynY
K3SI5ehLe5dpxPQnLgIIm/7Kz11Ox8hb4da2uarX461DiKdsVXQq6aGScezWPAsM
wVFo2Uz+eMi4kaWbC8em6yHBG+Ep1DUkWFEL8VqpV029TB7i4aMq9RLhrlyfQs4/
mFr99efWv9sukNEVshUwNnU4DV4uFhzo3e2T4koGezkAeeqJvHoPDR3+mllhXExL
t8LXL6oRDLZNEkJgXtfgrZGCr4cpUgJW+1++3dVpvNIdpyvHCf1RCxQP4OGd+8tB
oH9674l3yZLMuWy1e9Y5Lk5RMqkYKEvRVagviKQD/MpYpga7Wg/LAxIxC88kwf7B
4SdahiGlKHINDZ+YC0YxpE1soWN/V3VmtVFJ547e3gQmxTlqFhZO6yHceMXUl6Bs
mKiBlMPf2TSqADtIAr/g/NCMrEs+D4tQhq1DeSKJqqHNmOREsd+phB86K3TUhvlZ
hSAQZJ8tRKFe4oGc/trmyNEatYDvnh2MyCWsO2z5txFioqFugg7edCAD5KnOZt/L
lp+v7I7T2Js3l+3NFvhFlFR1DEpEAEH1qvJ67T2KZl+a+ruCMfPUm1hzdGGXHRVS
iJ4slClBv23lcGtkfIwPQyLgSCC2nhcg0+dCyY3GnoB3TWJbM7cSP66d6HpTw5Sn
F9Qo4UhAWX9q2uiBos0Sf7fQH58wTOWoc9g2quZQwspXDDEH4A5gIOeXgSp5bwDu
SwlTYsLW7sXBw6cDEweJVgrVZwFMkQqcPUuLV5WAkXPg54SDHYOor5QM4PMtBhdo
6Cz5I8Df57LUIBrDC6jVlf97u7gPMJ6kJR7MSILxsJ1AdjfJ6XhAwcADczqHLWUe
9qp2e4k9c7SE9aKdEJelbXGk8V4tt2HpxZYiphPGpwWmPoh07spiO7duUXP95Qng
o0ngrTARx0jXxsx7cn0fjbEnJPaRlBiet5/1ktSGqXV5fu3c4Wq7Qmn49B4v2GPr
ghTGNgBEU0BAr2IEBYemworyXJUA5JcaEJoH7Xasu/G17ikdRvbTZilYMcZ3KfPO
DTWO9S7ch3y+ZTfB3AJtq5BXEe2kemgz/aGH5YrdmP61dCmjQpAj05uOzVv8B77A
+NS3E0zFI5XiIomcRrb5o5+hm56pYifnMy3aGbfZN0YsCoO35immJCCFCvtt8J6j
cN03y2aBO7EJiOGY/X+lhyzf7jg80DK36Yj8XxuszhYsgusk8pTqdWm2ABdKMfJT
TtfhJkURIXjA5tRR/qLk39r31RLXmHBvd7/FKFm+5aYhgdtCj3G+iaKSiBVL/FL1
FupML/McV8S5tP57vXfJMKzBD7Lha9fRPQwQ+8fePKXNMEBT49V8ewB6zcTUka8z
ZgTcwmajYGOKCUJpwGapEFK3pVTStKKYT0MWDYuMrUwk/wb9Uj1qVtOW/9oAD/UA
6HGAGoAGgRpRY7lKR7wpApWWweWw8iI2YZaKNHaAdaS1+EAS9O+hG2BF8ircnHoI
zGVe4srvYhqJ8wkUfiVB6OteuMqTYgNpiAOrADoZArxemhMsup+MN817ygv2Dkrb
ehHx3+cs9ro6RcvDKWkznB/HIRILBxb+TdjuM4Dsu1RxOIpp18cktx7G7q+D+19K
ncQQQF3E7BQmSIRUcMR4ItGVzPZtjzXVGXgfmC4omIBCnRDU75XIzNdOXTOIoM1a
liBhh+KmoG3t4ID/amYxvbzLpm9OExYFwXfl1Xe9MNKQ6240GafqHHEWfgeYOFE/
Ru5d9r62OpDwrKJMleNpNMZBXa1bBBbNqd1UXBRb+BL+dPVIhSoxbIbQwXO70jrb
NRT0X4EiIIuhdNI1L15bLTWS5I+6/EeW7dMchkFodJDSquvamX/RYA/C6g0LutYj
e3yMj/XLMjx0b3jjy9kWqfwbrWEIlbd5t2Fx8dr+nwHs8C7TCfVKf1XU0bPZfETZ
iu6OPpw4dZEQlpPhmVd4rTEQuTu5OV6uZMfhC1Ak2BQ3BJHjuGsuS3jfEPbWMrnU
IGVaANajwZ1LNKKkoCTFFm8wCirIRjyZTsbEXSlKDe1QFavuxmLvxdQocChZCrkh
ScH6ee+kkayi4ZMYh2XL7EPsM2mYcCrgeZAV9x1HM9MPI8oBNDmNsSekZlIxfWag
wSA66Wkt59sQjJ62JRsFirRltUAf5FNDCsCORytsrBXCxTOF29+Wu0bexHItBQOB
mkJ5gpfApeqhaVuDrnIwZ/y3r5e56Gdz4yLQLaqj24Xq+yggJgr0dzLrwX/wTP2V
InFW9vIeXMW+LwVPLgJMTcz/ncEk52kuD5pmEJfQb+iJT+ausZvxID/KSqsGXE00
eVNNbUat95eYzxvAKFx2Vah1FLyG8UvUbF4Jtj0yoDATiN6fBsaT1xVkosoUyOnR
OorOpA/TTpN8NwllWIrGcY43vTV+uG3HFKShPCo1W9e+79+jnF7HhJrZ43wd+qoB
7szZb82CLdTVwOK9YKF6yzYaSmAZTkDn7ni6/+Gjr3TssL95hzwjzSYO9XdVZOA0
qvcaRBw86nS/IVkD2gfVPEhYbiBQaWvjZi9B4wR/RFhl+xLmvZ/HzXZTZJGXRIZa
8/88aUnv0YURs0ieBzBJGghSbqTwKzyBQdR1Ab47ocqE8jw5zvfP600FVpzjEB7P
qpNfxEWQw8D7PrvyeILKL3f1IYJSTkkX44Dzk+LWhC8uUipblQd8yjGuahlq5tov
Y3jWH1xtO5nlpDrOx3ySVLxrPfLgAEToc4R0rzHmLPyN9gqMvIF8oPIIeZ66gCwU
Qr0oQOigP3Jr2RgWrCMl3+wisqGmWwdhMZ2glmwYkgMMqeZtczVot6x84SVG5b/k
Num4Ap9Ya6WzP8LcOWCFC5j56ICtnQhqM++Ln8FXl3+Dt5ZPl6ai9/edOSC5/3Uo
D9LnfjOuzx5CvBso1FEgYhDbMM9xwbcPBO8tZ7QyqBguUSCPph/fVxVKGhMW0ytd
aKJDyVp49g+7fZmr0ugRtcqyOkQhO17kBGWbzFQFTlDCP4V4f8wTJFx39TDuCLf1
YFgVfxD2CTVTCmsEkDoNRCzHWkGgtjG55TtuFYDvnwCxw9ZNVuxXFQmCojix0GtY
+OQdmGwrT5+vpMMHjF6YISAo7KQoO1zNC0dxV6DbgP7uFYN22MRHdsAxCf2ElTdQ
wvjuSm/VS4ZRZvs1eBCCBobca7xy8XqPfSkOJT8WgxWXI7wNVbkj94L5gjVX5lfa
sFrrrkIQmoe9ugdncOhW/cfQ6PmKMdIiylBf3WN3qg73vhc3e/Wq0OkRsKr7PVuo
aKxLr8HaLLFaZ5NecwTqDDQhRDNNdoJUnpSKXwIOQMoHJgKA4jcuWL5P5wUiFbzP
K2XlXHLVM4x/6Ya488742vsX23h9z00KOToJWmL6ysWAsju6BoUZqSqPmyIqrvBe
i/X1hY+8PWPCcAj4wIi2vEO8lP+eGVx4BOtkx710fsrv+CLLGG0XtpFmStJtn3Da
d4sR+ViRY+XvgWWn0O8kVWiDcFDWy1wpoW7fEum07r14ewM3Ekfj6TljCUJYAQQC
05w+8L+65dl5p2Q9uDuIaYtzQ6cx9UQlBfyaxSxA8C5KnNzrX82kJVj/FL00SFbA
9KxgbhbXTYoRmtY04/kw7VsV3QnpucsGSAt1qJOgScggD0zoDzvG4G7+vA+dXjw2
EWTwe6GBHBWDhsmlsThORT9h0xXipWf3ESS1tvm/ZUkNkIWiHTowMzRx54DCuiUb
5s9SLgu1OQ2F4Iat+J6phoXmWcEuXydPECga6DtzDHNOZIjYZnxFCfalBbydcVxT
6cThl+ZS5bQRjsN64Np+46LEEqjfmK5Rh52aA4ALXJUw9TjBAwIY+JKlfBgs8czE
CciTZB5WFL0tZb0CndHJXL69iRXI++JQneelPGmdDt2BuOphMKZiF+6ZQR0rw0La
2zNH/dfggKreIXeXiVNmiYEleS0zypRSGMLiQ1eNB8+ze2KGhfcKuSWRQXNHN0BH
bwXDMp3aiz7NPVqdvDc2eP8zvMhNtLNJeZ/6fHkdbNna00ghjdyUJHC7UOfaPsnQ
q55h3OYifjc8AIU5G2y49StOSabPU7vcFwjl9LDDme70yc4Gs7kzXn0mSFR5wG3t
vWlQnNTEQEDhK8XzFhT8ku9t9Mjw2rI73fhcwc9CZbrb+g0TLzyHe8Ko6QPWk0az
WsY8z7MOKwtVjCvrB3rxrnMxBvLDGonaPGcOFTQ5wARXb/dmbRwRhBu8sCQJ0PAA
6MYy4yhC9fRGhPmvH8jAm1GQCBEKPh5gxgcLL3uHsVOHaAkacZImAyBqymlAVzAv
EVhlIAGelHI1X/n/iJiHES5egvQiQYws//FmuFmQFhvAykQl92cRm0qy48Awirua
mvImabni/YSxlC9cg1hXCYLS/etF1eoDir09V0aQathzgjILwgwIYik1h2PTwlsP
gJ6sF9OgWIQ9Ybp0+SIri6bPHABBcMASSl7okbCGRs9Mvx84pYV0rk2yXU3B9ADm
PDzN1n8D9OOsiOU+AJCe/TwYwq8+jfcBl8dNVaPqqehdcCgYyJGxoDgPLTUoOfmw
lX/jmICQ3YFgiN9Tmw82cXCuZKWOIfJyL68+hSJ5xhoEi0+6cEdWen4HCzh77yoV
GfosCiNL+rRCrjLEWq6VxhBRFSztume/GRVnsHjYYKCnzjBKd+QnJMkWJVNp366S
I9IC3Aajs55wrYvdmVoZhpeczEdtVDVaxo0piS44qaedkEX8FDu3AZfT3AI2Fe8R
wC/augftBjDP0uZJ33DzH9rdSjrfQnphRB9BQCaYtPv2jyNWXCNEk19ZkLpyHawh
S+m/V5pksBYZX4Vc2qDtK/4eWoCmnsVcjg6VHPSq+YRq5tz6aYNQ2Js9g5pXF4lo
E7ou61OV1YmK9eU05TM0CPRisHpc5Ragxq4T1cGLJpOL1TFPgTRTdqHDjzOsomdF
IjRtfXvLAtYcJ7TOuUUUiTYRSBrvdwqRb7TPf2GSc+jHwX4yMXfrs2XglgGA1Px7
IrsRZU17ZMwqWokCqBcRWBQPNmf5hItUoWeIK8m7E6WpGN0T4mNaDiF27jki1AzR
rV4z5ww33L6wG8CqXoqApQ6RrDrq9I7Pv1Apfn7f+X6tpSLWGXWkscVjK9v0xylF
NJZhX4JZyobuu7AfKcs+aHxRHUzLkV7MTRc2iFOqugZrRxMJIn9BGZLskky+Bzax
ixSysNKxBGG31YtreCwwx4gM78NkCT/Be2VDN9BSAwGGFEUGTN0nfo+qEBR44YL1
nJ+oVUiHF0psYSNDoxbsPaGaWs3UpZrVYLxr+H+7u9bLDD9L6I5V6MMjXH4wLkKd
h3aYdpLKare8J0ml7Q03lSE4PcpJo48n/ogjJfYEcb3im01kSoWSb9lV2Rc5dL+g
uQAMJQENpeQg8LvKftCTuKIohd4s71DYWh5TCS4x8deFsxhgoxyD2EFwHt2NBZhp
ptxVJ9AsRDA264rseXP8F9baep+a9sm8lYZfY/qdY5CT+VSQyNQhSxQsf8PUFIYF
IzobfU6MBTgKZFpEPGVdS/KcDmYz3/WR+YPPYjMZttdoTNFS361uIsUvX9UoxzY9
zJk9GBzkQ2/Yujnpw3bYIVYyCF5ww4mXWBpe3szKhzmznsGEsPou/rgzN7K9S0iP
WGsLDh24ZbYHG4mYzjtcs3svzLuMmXYPH8SJQgasFuAm8SJPNuQodXMuLvZeEAJK
1xfeUABZekM78PlKF1yPvm6efG7obbhcp7ELCmfFcIcoGH0hjgQg1gtH8XrMB997
wCVKRZm5T4IIehDCU1yZvI9lCjjfA8NkbOqFFi7fB19Aix356TdLKQOfp/iMJQYz
fEj1Dq9tz6/sS8sRwjliQGcEAOYDPlgerFiTC3P03ZI70xoPy3WFITQSekIa9FU7
fdq2FMj7ue3GBDSYptZL5+Z+vNL60VsqTDSe6jAvUq3kFLoys7jHO5e4y73bgzMX
5LAN1cI1KPmA3gkUhN2SOvx9+cUev7HIvFxtBhRYDaWDjXBcRZ5pail+sd0VpnEf
xkGRis4IrWihHFy+wc4XCaNo2783UOqqZI+pkWfFkp7XXbN+HRWq+INjVeQICIsw
XJzj3YhSkdS++jWG8eZaLMtIT6N5SvPvNShCv5OI8ik5wiaNunGQ/l2t86+JniLs
b/QdXGMP6HmRLP+9xet3xfTOExicOUkZKgiOUZYjmbTt5rN7JB2ESyrXzQfIJ3h7
LeQ3Qkf88rOZYcLNZQfDXsVIGQIim9A0tqaxWapL9Mrg8k8+uBD5DTqgp1K42tvk
K90zwAZ/Z/yFGZU0FR5PJEEDTC6yjrCC+HCeXclMANhE+62Vu3g9KhJ9nFzf3tnu
GYPp6z3qHtXULG35cqry/fVPzyCJBbZnmw4delPTEMSRBtxm0BFNtZxBqL0JgxYb
bLhcN3f0B0yXmIQ8mKcjalqMbpdqBvtiUPa0hZKHLZSkoTfsrnGaHh+2xvvONhqV
HLj7cNyyooUimifmligtKaHmoE1Kb8KdLoxR8vvXUNuJxVBt8Ubv21g++lXK3h7w
1IduU2i5qcumvbsroRoDUZAClwGF2W/Ku35TXssEbj4+k5P/4HJ5wsv3k15IW2UP
QqdpFc7SYWZ3NAY34yMJ4mXn3Z9+HlI0Lmkk2dVc3cxGmtUBk1ayxcj7Y9MdwjT4
rJlSnghBsHO0kOi3ww8Sn2h7EZlfun63YzfK3CervkOFd+bwq2oHpuU1HOpefRkL
R2ZWAxaPtHhJoKtc5HGrcBV1Y5nQ6BUGHbJXIlRCIKS9yhRVNcg/KLwlfmATyOY/
Zxwm2bi9z5EeKUWvmhUaO1ClWDiZ2pLhy3hM+cd+Cyv5H9dicWOFXvDbhbYUmSSf
y+BF5LUw3PSwgYNxObbgvoYfMY5lUyPMkRHJPNryRrWpZq4DdR949CrrUgv6zQ/W
7YTtQNKGqrGO+FfwWoGr//Xkq4bK5D9EjNWPANjo2w3AxzRKdQeXbnzLCDXRbLXB
k9iiz3u6CVyCL/dy6cAa9cgSaMkO+WvnZCy74QawVYakck/5k6Tt3NWTyynj5JbL
w8/daRSDfmvmMiUGg9Z28R+N1Xd3OsN6YI3kN03PjAkDjf5/NO3ny53Rzt8gwjX/
tAuqrYeCA/Ym1Rwf7N828/JXJHpv6pKa8c6zUYLStmW1qhU9nJGHvdYBnbXYG5sS
5+X2njphVwfyCaIbZd6fLEa0NCXZqgSrMyykuwqA87JZTw6wkeLayTSOy+aKYVvY
RCZ/TqlAyqYrUomRtf3M5V9IrOSDOHOIctw2uz24dz7jI0pqbLKQ061SsQNOtMJ3
PtrWEyOAss1IZ8z2jC05+xScUH42CskS76tsm54/5h83w394Tmb87F1gTfxw6+db
QSk1H/oUZkLIumpxBCS3SWk7DlyrttpnjKD9OGaULmLEZNrTv+SOngTSUneeIMl6
hWZtQALuQ82QKzhCUe29AM+b93e3KXM3GWKZ3CUe8gUSSbeT1Xfc2P/LSJbpqgW5
AlSOKXQsYrhWo5/lBszBZfmuZlKMfFOe0tyZCXL4kSDnueJ8zYOO+Ca+zPzm/DuM
G3t2lRcgp+pOcUxspRgY0B6KByA4Op/dawrppFaClCTnyo8hdD502pbBxCarP6mp
GcP2JYb5YplGHi/YSyJ+jhE9LpZIf5DTJIEuGpNYiEYCNqqqZIQkCkTk3Cx6HIuj
oHeXTZgK30goCRbLW+PpT7lQNYcmgyUdaWf/81eN5xzrx25i+hGdf0eoNWejLC60
ydJoyoowVpigKgzTvYpUbWJj8KJbAXFKLd6qJOWU6MXszqTnxd15Cxw2vbRMtNmb
+7HRvvrD5Ah7SKlVq1WCgK06qb6xMruiZti+sehSAwKIVAjCsEU1889S+H3VM52y
TT/C65Ju+WXUabWRK3Jg13RtwTeqFwkgu5mSVhSJQ6ogWC/VZp49cx1WlcYAGueQ
cyY2V5HY8NDjvUzJ3FU9rMfZ/Hb00pkABoQ2OwYBTZRWrcm38b24vd9chP3AjJCN
o+rpUSmG9ccwQAG2lBXfu8VA1CGyP2J9WMoc+h6aIfIIHpQqTvU8II2jinSRQJUa
pxfP+eCADL0BTypvxoIuAnNj8H/syQooKblRXoP5c0j6QVaNbbk/mt0N+tkzZBpL
UzkIbD9lcdp+touOZbS6yaZWn/A4XxcVt2QFhHfIAxfpNWAauePNU8OEqK6I9zbL
xFh2w9fMyRQWRw6VZm/UUp0JELyJvzzdROk8F96+DYq7iNXXRIBwqLeWGnicJ/xO
U2Bs35eIXvqZtdACuS6NKWOWM2XZwwsLAG3LeMnLLQIvRRydVI2p9pd0Q1nF31EV
ukpKukBVocqW7EQP0Scz2LwmXxwKbNfUDCQ9UGL/8j+uheMmHvEtyEWKA7Gvvk6/
2Whcgzc6Fcml3mwh371SsoX7AQDxSrz0p9AnaUmuU+kqtSX6RnQT8YHCC15KNj+x
pgLEL8ITlYLiU/W8K2hoFtvuedyMNh4JJQ+PRxknKXxm2OlvXxwsP5mC8qDiwG8r
BNa3kF1xieWZ5q7rDUFPjbArkjuQSmbyjGqaNZNHUMvriwQIGU7I27zksv4ZntTP
7kXip8L3vnCZPnjVlUQ9OC80L5D4S8qMh/yXzFyeqFUM3+ZlqCOxcYf6sYJwUN3y
nZpKQwaumzio4KOMz37t4qkGeohlhtWyj+PPF58u5FC4tlgI5glelkZa5OqrWc68
orT2Gy0K+V60sctEa/MkkRCz7NrJ6G0CY6ZKlUGg6qR5FQnaJBpiWmYyo2jRPzv6
GK+a7TjVO3ZW/M3jO42syh4MUb1D6ol7tMY/U7aD96GMcsrgAKH9YGwZ87WM1S9F
isO+iLWVv+axSJUe7qbg/NDfgyUoO/DRpvZng1OK8AhwYqRNnlBp+F8geICoGLJw
/E/eXTJxITfwZgAvFGrneoVtUYmjjFl88Qcc8jNOY6aBbkMyzomiZAjvTKlOgMK7
s1VvNbLOIGvmDxOSXkuuQgjw93GaM0M7s2A5ezueeqb7+EowwUAAP1/CMoo/+yeN
sZYQzD7GhWflN9Klt5Vboaawd0unZmQK4bp+yBWyC9SsxtFLuGRX9IP4Ej/HqioW
0iNz/Ap/BqNSIzOBGmZS7FJ7T20tYs6cgTPk+LD6WfwHSRQI2SzSWjael5qwNY6X
QpKFa6lTv3/iaRzSDSUsEiVtcY8nvD9ROyPsJm4lIpEiGJPDUHQm+IuTTvxuMDqG
sHn0HJP468rjoHx9pyvx0oXP8xcz7C2mrDgD9PDpotD+AbJFuDUBLwiOA9biI3jh
YQ4ci5n5gz6M6aOGhPm6hqxlwHGFT0Ocz4lHDJtFMj+w0Q7buTZNHV9aL/C7cx+T
MaRfIYU8603xTauIqhkYEHdV05EssdQ9VgDDVzHKx+7zeeKqsod189eaMBh1ydjv
mXTZBJvAEG1LpHuG1bXiUz/k51Q7mnQBEkhQdWSwwJ6Lv5nMuYFLHpI3oOsyHbdh
NtLm1xRjxsCjFndRNZ4jKx72kxDhaCZg7VSDtdVjkeqU4qE48PGQO5FPAyPrJ3bZ
kPUMqJ6sTNiwzA2xokRHtFovhl51QOhR+soogFiM2TlXgHc0p23koQhVPodh8ZfL
K7SOCCyPMgOrTvOZhslv72uJhP3MAQirHnhJ7p8wf95alpx4pPK+pl1JMr6OgJcm
iQ4p/mDDIWw6bjTDNTlNjnz7XGivxry4bSE+ZHuWmjkRfuVPbye8F+lRFd3AxQXH
2syBsYzZ/l1nY6ZeIXkVMLnO75gm5ydSsIrevho99UtR1c4viu9mNAC++FQWMSVq
vuM76elI6DExx8BDw3G/7fzh2/tOtSOTqJmBSvANnnLxsPF81XCLtiBk/53RdDNL
ySkQuv9IXTJ5gsCwu7GGgx7QXIDL7wY7y9HjMbNo4b5VM0TCn8tR/WA09Pq7NoHC
biih034viVM+v1Cnw/ILOC/p8lbEmTdYtLCZFHv0HyuRv78Lug6h/0R5bhNRxs54
xz+Rd5a7U4d6yUqk/fLyEtlDzMsQwgNUON47I5R/ErxL3NrnlsFGuPJVQVK4Ic9J
pdt8nfRf5WSIiE14xF6EyeahJWrgcgPftdNtzccEfta8gjZ9ZRc++TW7W9IBv8S+
BPi7S1gMKipOC5x8uQGGQaMFWIR8+rsQThIWpb1SSsQVCmFTtaYLEmLbHzP1pMP/
w8W6Yg0+qPClnGgSQxyso9ED3R6AOMfbxJi6U45j6rnzjX/jQojXv3eIIQJaiAzC
C3ojNSeKeoNcyInGkmME5h3d3tUJ03+oG6IHpF51vgmu5EfXKgCjGV4aC8Usoicr
IbyWS/ZpyfZaKSnF3jpdiSCorE5HBIPEpdcV1uHBvgFLBjkCJdKJOiHgz8ONjnYR
PHy2NaogzIhKVX8/tOSHZ0pM8r7Rz/OUTkgyv0h94PHgM5fOJZ2d6Dg8Muvt7fwo
N4qQYmNl9Zc6HWcQM2AeufGXmSwp3XDU9EmhsOQMs5CsBtNWWZ7ubNdi6gwe7tp/
IDwtfKwd2ng7hubi0H8XzdxbNR26ea0VgirWIiQwDlRRJa6zvqMhHE3JWDUZeADc
T86IWw1VE40veYdfDPs6aSBFs2vVSIS9DSexra4ltQOK0bsxRH0N9TuVahE97J59
KyYMdt9eXqBDX/8etRa6TA0nmWBt4kHZZbdKaEr2XdywQDeWl8DnIl4Yle9HYH3V
vJBobp/n8FI7hkGBERBWx/64TPXIix+hRw96r6N5DAcoMRvfgjlJNY10VsHh4U4g
65Nzxk5mKUJQWr/nHosyyAH4cxXzg2IRHYw8bH0TkvCZSJd5zzTFfxfiixVIKveA
JnMD7xB1r1KajAGO5kJg0LeToZBHnQRGuTM1DyiZ08oBvV2Il8wPG/WBEZpcEfeK
vaIidzPg+w4fl3sZbEEZnAldh4TZyQYtv8IuJB3DomxzfE/TBV7rLfYIRQtsZMTD
HFl7xw/EEE2GO6Ekqictr/Qk80450e95mdw5flwc5pk5fhTGSDDERlQ/oF8m0fQs
OuRLycuaHEK758LBYJsLhUHEANzigeqFIdeJPQEpMcGlX1fwh/0UROeo5UB0FXAW
CHheedUF2WSLo9zRg4sXKwk28uTXuSMED0P7Y1T55i8+E7kn1vHZCCDOOsdiTv1u
JLkzxuGEKSByTA/MFzb79N97CLH0rbl4VdcSjE1kPdfp12AF4ukXYT6/5VAClp+1
G92Dh6b/l4qy05A7sz0p/INU4/Rn2YZtEXOE2x3Ar+IvC9IC83ktzWEKcw2BQ9w1
wfyinnO5bN+z1aySWWIMD7VxCEQT2FNrBfDvKR7lcyyfHUi2TZ89rsGTbG4hCCcf
/20wcVzPqTtD21dpF0AhBjvy0m1f7E2rlii8f10dC5I+I7Xb2Q392gI2pR+qlJ0z
vM/WPKdd2qMBuvv8qhZA8dmMdT0NE30qSz/02LxtkA/DnNE/kIijMwnpX0pc/Z3D
oqasr5x/u4Pp+eowIoXnY8QgV84hCg9VyVGCU24htA1QC19++i7jWP0JnLFavzHK
8WOW2zCPw/72Wpk7wR/m7MoYxfoXKR1Ejb3lQ+7H1iKbplOa19PWIaxhdhLURJKm
04S62+7IJw8/f+mubSChv59Qp1AC4pgsPlX2Rsuay6ui6sz93mlsT4LGD/su1EoF
XB8pM17V9pp24dcGNuMLqv0StWChtR65Q8CMqTBahIOsa7H179KanlhhOdvcyNgF
AHhbZQLp6LIB0DC6AOXi7gdTDYHFIYlHpc9SAmb6rZhwz758yWIaEFjtP5SMNhP4
Ogk5sbqGhYSqJRfvxb/C70iupvWpxHesVgTV9+t3gg2Tn9Z088pPugV15doczmKr
b2iSHK/83KbScVAexMs2W/vRgMT11/KPgU8ccrifSyIoFFipL2TPVImtPtJvGH9Q
YMOQu5Ck35tr91AkO7qIAnfPaR2EAlkIkrMnIOwRuRIEE1nWGAaG5CLLbzFnIsO0
iklh2QkoMuS6gho22FtCtbunFks9AW3zTdfrNs5KfVrdsjalB0dSbq+Fhsr5M45g
gH7+j2w+Akt/ZPqVbd7k0NkXYR3SjzjXWWpEMKtFpO44zX6oD4pWtjNNc5PfQPMZ
NFFgpjvRn5oSZqZ93rEAfFMeNULzjylTy7a05ADiSLOnMWibDXkVu5zDFrtMw6VX
o/efd4Xv6d4xFkZqv3JJGBr01wMqpnqpPtO8sHbKFDACDR8TI/MqypQFV8F4sujr
BYVNwdjVLN0kRvKm62a8K91nHJJkMwihVhdS6tOgZgkz4rrAjbfwGuY1IKngnq/A
KN4e9/tp0qq1jgHO8HUf0YhScyms1sLbViSJ2/J3AmK2MIJZqcAotf4Axt9kkF1r
+og8I1pXX2F6KwW9pXv1+8ekyYRvNwmVu3B29lQs3xuN1CjL8EvJay3AIuM3snjB
tY+oqSfmLFXfhxtvC8c113ZLmHaK6XHtmNPYdZOYmXEoOIvBDKEkZnsBnvk8FcJ1
urPqmAGdo4uPD2r8wF352AaAT4xjYTkm1uePj6VNm6gt+wWNaUcuLIJfywj0COZw
SpCCQSp8yXzLcE+FwM1iwtF0QFg1Se/mU7/+YY7mUBJ33wtwan6KkmcIoneOZ6i9
DIEbHOsASixIajYBJeXNz5qeYk9X2vJH46PI6Jin+zhQccjUHmisIE6MEcXB6bGk
VPOIhs+eYKbeuTVebFKeqqEJFigoJQRBxZk1oq6KhBw0dO8iltHs6rHb+mkTY6TQ
ifwV/bP8ymks5hADPceonpH2dleZXI3pjEkULzBaMV/Mv0VliFgXLYXCeYqWhnr7
ItU4HpIr0QgetAJMw6qQLtlfzC5JChFCINuuXmqt7zIZxUj+gJHKW6l1+RTWkT95
nA/EGqjZbB4PbO9nA9ObWyLP0goDjppBpCtsHp75SnNtnlWtTQgeikbhiVhH6Vdn
8GSac4UDyLsLIqCptWfEQXDXUTYNsAL4rI3Gi8oAvqinp6JVXJFidVmynn/wnWj5
nkVXcvLLCaSyqbdFxZvJj9+vcxEbAjdwwKffjYMG8dft1XlOLk4iLhyelB+/ewgK
awLI/79VxxFuar1pkm+kZCXEy7LyiFJB5I1nHcKjfb0tkvB9s7eGPSCenx8gRqbC
C1FF7PP8Ur53rj9gJewAgNlEO4BE5epJdEivPEB0DHxYXU7Nm4DWfn00lQz6FqLW
ecC1UhWP/ZZhU/iAFGfJCv4MyVRntEHV4lZaYOX+Mc3UTNoaTTEKnOamoUWRMB2S
q6WX50waz+hHnBi1zX0u8tvLW2O6U95jGRibqsSNSN92IuX5GMKqxGgzalSuLQnG
KO6HRKEFcUEjbb7B6/EYwNPcm4BDrbobrEL2DX3vMbCLtLdJCQ7+s7AyVb7vwfjS
EC6olwFOu6anvsLBWgKsy7cOQAJqMOUH61k/LdeR6zS77WoTXcYR6T7Y0ZWs/dlv
1furg5gW5oA6mnJD4nbFZzeazWD3EMcz78rfmkrrbYJ40YZAwvH/UyTDRq540Crm
I89MP7w8dXLJtSdZOfdWcZyd2mALJY/PVTLaGgw3R8j0ExxvvFNz9oM1ENMMxFz3
Z4GkFDUChZo0mKiQz7WBD8KbzgaEeXTXLp9ELrIgCgX0/IMYco3b5NAUeFQN4tkr
EmKTHIVPEZo/0FJDADuNkjph24jqshafO8MDNR1zezbfp3u3+/P1Bh3qRmOLs/Ik
8vR4uu1vGF2VhVUxHfb3tyN+VQh+s/OcO9bydca3NWKMOJ7iqtbn/U/58WwmCgtj
ZNESnCCMaJsyXOL+3Zrb0Er5RffpvJ5eS+tZg6IyhoYtTrj135pZhj68v2pJcGKp
QxHQ/2W0fzDe327xbQkLlQdaPIlZrUgec0187icAF3Shutbf99SiuhpJj5yNanvN
V2GS2CujcxMno58Kkf6XJNhTBWh1SVY0NL67lRPyvc314omu6Y+gpd6LZkhxmZn6
rVYo7E8+R3P4/jVDNK22gZOJEmYT4T2ctnTuOJ4dxAt3p+dAe6XJwiQ9l1r4k+cK
QL73ysJnI5/Z6rFAr/brkrieGeQrOUmUnMGs6ckWS9I2Wt4TFMFgbZKwCrOt3ZOh
Z3Y7rGpD8JboPrvSyca1SrxDDD0gjcbVksgE0DQCoK9eFhx+XCsY5vcV7HvdInP3
A7+1Iuavoudbws9K5tNzItWD48fPcUWySkWyp6Pf1aloWSP6S+O21V2F/7lfB2yS
MG+gsCiKaY11kIiWLj+ySXQVf9Z1HTvw9JPy0RQSrU3Ci8XsPhmLMs/z5JEmzYDL
qFKuc4FbM2iiqg5x3si5p76eO3UxG8rSY666Rvixvbvpu/2BNrCoEeGktYSvuc7m
0E0faXKgc4RyvaMnJemiwgF4Iim7a8L9MpziUflft/Yg1WYGYEVzUGuEFP2Csgby
zWo5FrrUqeRt2KvkzxQ6UAYTnhV7ZCoUyo9AUxqsHfdKq/pymIMszN9Y/V07PFPV
Dk5tg+RlvBNIjoqxom+mxPnX3icA3Upj4pdEypmXeutVymaTuBN7GOrg8GVarG4t
ywtD14jUZYI161ZyD75T4RIhUqCZ5iZnKqwpD/NrMI9eURF/r8PCv2hitxPf1VIk
/fLb23qaVNup7L3jc5SjUoiHYolZ4ASIxinRicrN29ltjk4hHASHgnpQ3eJzK3D5
eTbhU7+s2g9zd5plQUrMXlEtjVBP6EqPAny4yy1WASTHj48xi6oawZJ/mvGZXPZv
jlYwAd0g+NS4daC873zvndPXcb720yAh/N1p8bhRKVyVwunppsI6aDBtHSsCClfN
JrRgFWPGbn/c0rMDMscBJNU97EBr84P4Dg2hh6j3yF1/U6Qdhdrhn+Ijc2RUs45k
vfA27dNj3XGbCjx8autBVluuFwhyC95VvGQQRlaCp9EYek5HcTrDZjesj80HXj3G
K82N+JR5TAvLzVUji/FTvFm3eSjFeU+l6hDLbc00VzT5kpe5QUU4ivt73IQb6lUz
6l3wuLsI/zHqmGcLGG7V/RrHc/YE/jVqdXiV4+2chPWlgtf4rlKw0nuo5vFW47VY
+xY1Kk5hxve8pAjokKpGUMHxMz0faJCPhy0CTWR5ZK5XNYMCZs/4PZTy17b9gPKk
OUFwxvP4JS0pmR86z7TIHxMakGCbhE4sCfwCDa9fkUjp4wm3/59/toH1ORsOnC5s
u7EcfY8+L13GwCWVWEYt7RXNxYAiQt3pnOoP6tKAtOwul7Eyc5wNQy3p0kunkNue
S051YfUSCHLqC2EBmqm18C88My0ly1pfRbj/pIPMGPykRveLeSygHnVQD4jsedxP
+dqW/jaZb2Vcq9YxTK75YQCr5ea/yNe3AB15yX6XxA6HSa3MgYteUnjTKOhCoTnc
Ui//Dq0VWeCdJpcSNSTFYeL4ItmAVFi9aODGQJwB6zIJmb95QQy6VtF2T/Efe3UU
D3xgZ6ZV3F1+HjCtbZT6wElgflWNRofe9dUl1/UU17Xc+r846i0ggBK50S0aAlZm
DrJ96d9pYA0FCr9eBb+lmkQrQ0yJ7P7indra5xA5GR+YPFz8bfJbsF/cfVB2TrE4
msH8GOcJObXNS9mUlsK868usQTbc9kTNky0ucBbImqhH3nvJIuOfEnD+yrHHpJNW
gj24bxtROLnTD1VWwHvAluZGPht9MBbvzFLsjIA+Yp0ZLkSRqdu91vMujEAU5kEZ
ABkx7pQwO1opSJ/dXlb36Ww+91FnUR+xkdDNpAFQUnY0X5cP5zXxKR1MvOGZIhfa
Vbvt/muECHjkg4MOe2LM6n7ny9anDJvbfJLaE1GampKqtyuI9p+ILJYtDvBk2ZWZ
rasFDV0GCLLJYy9JgMSvVI1c39T0sC8LXpDuRgEG+3Q3nyGa1WrJYWJW+a7u0lpQ
KlZ8FJuqM5e2dhMzBgUG8jguTlilEVbC8qgc/jBCdGeCZ+SG5u2lMTujWzlJynD8
6RgUi71lJswmTM5pzGdweEmVo4Vr399FMCXemEcW/Hykh9hIILybsmfn6TycVNSo
7nwpRx3tKb6FhP6HDXBZVMzDCPkNOaY7xeOO12M4zs3JgqOPEzvoAE5gs/NF5DLr
pGNhvFDOlNV27Jn7WzmChzNx2A+rEPI2bt1ZIGlknWU/xQ3IyU6rykzBZeMC4ymD
+H/rXB3o6oUyFM93SvxZBtbCybLHIAQbc6/pKvONJxyeX9gWvQahFczxIJTY/e9W
+vptobs2POD8HKeHY+S+rK3mAQ1M+zmJM/zzjobDbNlR3MASSvzbm9BKUu2br99z
mf6vlpscQ9cFJc9ghXvAJW9rFFDEyAW1niVvbn6BU75FVHwRYvn+4aCbLNm3nZqN
rhI2UuXzJxLLTdMx/1EQznSTzJrDdrsvxfDJcst0rH0NiQGk7ZDyGIjAi0/GTRND
ih1PVgCB045ZF7GLeLGHgOOlXk1jdVbWEaV25GGVLWwoo+fMI+hmD7381sFcui0s
Yh4ZFe839Gu9a9HvZ2ipqEOExRJUxctnntvThbnjepdr0zbDppMkMigJZ8sGijNT
Dg5+lHlD02hgGApkds2/JBcvjEUS4oz4+6fdXK+eUBNJScrqQ+GE8uugFE2WVSYO
beG6GS26/xXE3twnJ+WnMonOv9QxofgFztF76WSsQ204KPYh7dKYAfzUXPibsk8d
a6lnjZ0JtFSaM4vvZjMxW4jJ7ziXj9JcCdYr2ZrtoIF79h2Xey2U9aWwTGGCzize
t9EXIP1xFcrV/jF2mnZSKm9XjBGm7rH2vdhHvSCpFkwsP7Vp8BNf+L4Vrv8rC/Ds
9qcOGsqhPxmihmnLLjWbt3kfrttT0kHjT1kwh8wOTGI9QJvELhwWiyGUGG8qdx1m
51Je/ntn4cpcocURHoVwmpdADauSGvB0L1agdNyDgy+hk/M9fLZcso91GIrh4NjU
W9kt1wjXBJffVbz4ZFUQuaWoo7ldNxIg0oA+8wymyPs5pLdcp+GIQEzOLXd3RZrI
FGZI4cNTyTcRD8FfHhEQevRnsoidWTSsXqPB9bQ8Ip/vEukKbcpDECd+KbT4zjR0
FWLd1BjQVZanzE635NDX7seJTECHmXqWtcJLanCtdDhxts0yjPAJc5MvUoGJTKub
0xI3cxpdaBokOe968NRvqgJSMzLhlbis7KJAU4UsuCQC9ry/rlLuAV1R9+gSjHjX
L+abNj8WCPpaLwpkjgv8UhRFH1W8HWx1KaPzsvi/p2BAPFgJ08JvcAmhzjYiCxTx
UOEzQVHml+oQOAiTdaWrLrVmJTnxxt00G0jqV+rIGC0EWqm4fjDNSc4ly43KPtb5
ZLuu8m9XcEl7wdh+JYdTBM5vnIk20OmouyMYcz+aA2vrqJFxtgA1D5FLXoLjp+6S
soH2ssAOwb46jqYuSPZD9TuOD2b/8G3Aiz1D4EGd7c2bwiupG7z6QkbtymF6V/G/
QFQGeEZfZkTJKZ7FzuQp7LUCwFMsT98eRUABtI2fNqkdpF5D2fTatiP70AV/vR8g
KtMDr08R/BYwMBqBxkcxN7/Q4Lz4QsXffCOHWloHGhqBLio7uwqztmLi7yJakA6b
xLw8nrDIMZ3dsaEU6ma8ff1Y+Cpq3wAkZP9bb70pVwXh5LdhqG2/EZ3dZkGkIvJP
zt6ckv8VvtjEGOPpSl2Qiy/IavS7lS4NoU6RFQ5lty2q4QvyxD2GHusMblPJ/gtr
l/noVkUrOpXYcqEO64Q7cMfXvPbM9KLV7eq2/kbqwa3CguM75Ij67Boi0+6gtf5l
DQmmiU/1HGjzhVdKLV/HLQZ3giGCRJiGFRlzbBT48WZJDyBtIVHsvnbSfOuN0Q9C
E2fXP0xD+ymQ8ZYltba/d4zcJwVucnDPS08rZQDT7CzqLcY5dj1q6iS5NRj6in67
mk/B7Ps9g1Ms+oZMormGmqW2mGWFXBQU5F24o2co55Iz1YMnlR69IdzAuLHdY9bt
UAG8Pg/NhvAStoDAjm4WeCpvqovp918F12FDLl4EF2hjJOizmGk+I2HQJ24yCuCG
75yoZg8FfkfdqroNq/J13E34xL/FnsgznvCaxQ2H+z1ANkF0A8ZPXpFQlUHDqIvA
Upp+wsXkCcOmbmXb1iyQExodRY+akQqDbtwkv5KMFDacIQWrz9vu2voOiGGFrUAt
YD2S98eT8RpRvyRyyEBDRobN6Mnm7uaEmnZ862tGdw0SE2JmuHwDcMSXD4HucC+K
bAwF05a01pc97iT93Vgi/sIxy360TjrybaYdqItLraEEM20Tm84juCq58vRNtkJI
NcONurSZ5f7uFO2dQO1QQUZYBGt55AsUgqy41nbvmg+PmWXX0U+K4en+NqaykVqR
+S2sPOU363xTUOe260LgQLw59tkEZPc3vyadnICyzrAICBsQX39IZp0lXdKcCs9H
2w0w9ks3jcOuZcEkxn3IcE2B3aAYgzGpIURIlo122TSP3mRZThGWWuGa2oeXCF2y
LC2syl8qbv8RZVNZ2WyjRW2eBxYuwbBqNwFt9sTCelBKjVZE2lsbU8+m1nG7LC8h
t942FAa3CLoquFD9EU1KQANx1bHWVb4NP4VlExTJTjgsGBmp7aS/D4V//N63ED6L
Z6agjmd0QS2Bj8dV143mRj3UVo6xscEd/7RW1XSM/try4JT0Idfbi8gjZPq+4LBm
uB0DV752R5uc3eINZq57g28cpcPJ9It9kw74MwGphm5H/8ALwRWQolSv0zZCM1QR
u6WSv0KcSFEODzu1whS39Am18dNf5o0s43GkJDbe5WSp4vpZ+gsMYb7VKGiTvDNM
PaZvp+OpkdJ1fobrzGbT+GSUhQPCpp9O14Spu0Vth1uPGIING47xwfUa+UGoFaCs
MoKwne0seJ/6hduFG47mdEugh5m9BrLQRy/rMfVWKQt2O3rkRd6cfG59/DOBwTAA
y4gi1+S1f6kJEWSb5YVkCpUACfuG2VtVXPfeWdaJ8YC7AVmjm3Sk8wBhd01cHqbz
i6megVE94+qZWvY/NgR1Uw2b/xON4MEVHFPi7Jumeh91pMLLwIuLTagdNvMiRJiS
mkBXz140LBbbj6eG8V56i91SzAXpQDNJdr7KFPTraJMLPWaBAJLNbdVR3BnUjcPg
0nIh9nsGPLPvDHnB8glfc713Lb/8VaJ2k+nLE1XTMn03gyeLWNRrH6fbR4Xl/Mor
MGmIe7qM4uwL9Y7bRPD9qXcmrCiDyie5h1UmvPsh5aVjYriMVW0YioLTBpCG3H55
hQZEvnK8bhtDKDp0p9QnhqUG5KfzQtjHla/pmDH31r2Te1eXzHNEpkl9Esy7nU9e
zs61TwZURRPQqRxxWmVnfka4OghC0aH6F4JLjvlrRAv/XD+7t6FhNKgP/3w4j5fe
XZtJ35hFGyewWzAR5CWSXH4t9aVacUcXG8Xxo5NCUskEKTNRacscKbKn7tZY30dS
IEDgwj6BObBk0k+kYoKFGYaD25zBzWGCTZ+TlN96zkyCTtbIOj6QQJ0opagB4cSY
P7xwB5O2xbYXbHWJX16JLEyMWeOdb2QdHJuqn1TIr7pKlqu0f+FVs5HG5kceExhq
zE6G13sictF/E5jrz1tuktmKr9yAnlcm7Fyh15p8OEsYfMQw8pnvmfPK2OYex/Yv
ni1KGiNN8Bpt3lNQ9aYtVREsBWgHMMBfKXY28rxBMNGYfdjDv0Aj+dYVbO1YPL7R
1JIUW034sJjZ4518+dLLhXs7297aAZXooNtB9+VuuA6IZl3iE1WR618z2dFqwCp2
rYofYToTkKljM0cayRHmOv3KEG4vT/d/QK91YEAOSdzA5EW9QAVm2k4YkZbuqGLQ
i933BWflr1NVdRyQLQ4Wvu75p4lYEFdOxHjlcr666uXG21aNgY9apFZuWAiFxYfd
PreDpNY2DxpFXTi7acGPStf1ZDTTNYyea6qim1CxCIJ9x2/mR+NT1OXW2DdIWEqm
uOUyNvFsF20Nbr2eTruURPQP8DUDqd7rj0pzvxiNZIcuNKsM6UISKUXCBVagj0Qp
7T8f6Ma0JbFRbB0+Rlf24urV2MDOhsCir4Jt/Fubrl5TOLgN6h0ZZ4fkDyvgobk9
18yB76Azn/AV1Y/utg/9yDwBfCRPKFQGXwZtz98WLOcU7feuNr2MK3yCYcuqRd7b
wOthTkTw7I9Q93FiK+rqoOAKUWUo1bf4DWYO1PiwHRrPWaFdwZCkqGcTS+fakknR
2utsYx4DhV/it6vrf2x4jdvet6uj+yUulifIR7Qw/cMCeXv/x998LwQplc+18oem
BpOZSEswxCBiE25FgsSae0e7WbRoaxXKF3DOKkg1zA6jv/Zy+bnWWgXKyJtGWs4i
nx2qe1yc3xp2ZJz44SbKQL4Z4oAe5D+hWfMHjwk96K5y6NiHxanAaIwoSWrIJfUW
8YeukXvfXTE1BKvAmgakgpLpvZybU3huy2L2MRjh412hIhvFwdApy1cagS4uJGmu
FwWzJor/R5/EcDu1tv0o+gbWDaC284xo/bqwkFAtk4WygPe5rwsr5e1TofLM0Zwd
VXHunvbjYNMhq7yCfIZGWdIOjuN52v/lE2XNMoBLuujla7+3/pTPZLh9g7Bq5fW7
ASqP9Gac32vMT4o/xyVNKBwXFdO2qvdJOZ9lrNmhkTcBdZvUucqdzU8jD0OEaW1+
TUW7kwV8Fimtin2EEOGT3ctPFFe/o4UitPP7TaBwEjo5YnE4JF/vgsnkRf96WILy
guoL6nwTb2fFCn/UscO8Gg2udCpoL0gqIW1RFjRt5Iq0+eWrDNrtbokCcZceyTWI
aak3warjc1iO0O0pLcUJOD+uq7+0Mkv1u9dexd3h9O4V73sfOPYqsulKuOxmMmSL
wdvvyPEnP0VSPwskPbzVWAzvp0GlGrCJbfmM7p0pkUlT3bnJgd7UX1XF1F9Jq+S1
+qvMLJeM+gsAjF8OF/WUQosWJuRTD6bT5OCq5c58gw22vp2xe3xzu10V7WFVyB3b
GH0+Gmar+bNUXz8nqPq5P/n6JN1hhxzejNiZnA83IOo35vdHpv+xa8pIohT2EMPA
q4lX9V9pouoxjnA0wgMN0AsWA00yC1rl21fQgk10UHWQY9n5qErLL69Pe/5lkl/P
QZIZMiNAhQZZtkjnw/YvG1XRPnMjFRDBH9WWpOjGWs9HxiB9WWLOIx2ODpwC5EUi
gSkFXolZ+H0YbXKNrS7r8bhC2S/z0qYJfZe4Tp8HTqXtgnm9x8uozSsm37qhanwT
gaY/HiemQPGI9lCbzVquu1cGhahKZLT7vHNydfDgQ5jlTPp1QqGPWJ4UpbMnSneT
kip2TKerNsM/zP0PkIUDPvsoXVoveyy3Q3Pz2He2qTzeoWTMAL0l8gZgTn3wqgHR
hfiu0aVcprydtx/11oB/f5QrFjtKaeg8bY1GGWpUzyBLLQROkLlZG+VZeswGOM4J
uHjx2hQ9Cdtt1LJzPZ/SMfMF8xLj6AacTBFwuynAr9lz8o3rc4bZmc2lb7vhiA0n
C3TgseYLRb2UXm34/qPSXwbcr9FUiq4SNMIPCU8GGNiXk0HD7h1uL/VuzU/lx7AQ
ZmBopAuWn4FvIsaO6XIh7iautK5uuOOKseE5Ukq9WZVqYEgY0IEyTwMXH2zXa0b0
E7NQF3cRCzEDStr9AU2uf8GgxfFKJLSNoqRMWRzgcMkBvzpHlqoA1FBtIw2jzxvg
5kVM3BS+sG0/7fG8KzU1/eZqrm2D+NNrkFKJA1jQaU4h7UnxlStVY2md5qjg2U+h
CB5M3sBH45lzjTN2BNejKDzJPp2v0p1TDa2U6/HdxTsOVMjGZ0lKAQHXAllRsRoM
2JExg2GfqlK46i69BB5SHNbAoTu5nVfkfip8W7hp5bc2SOEw1osrG/94mHZ/Rkyq
0ZGbNx4m3Box15aV93S0Sm9WlIZfzM5QOSxCvgZBujvuju790/WYFUyQHriJ4BgV
dYEzeB04/3Gs2Ug68ScNkH0+8pIw8Mu3peCNVDrPwwYFVAgDHlaRNK6rx4njk7YL
yAW6ON3Gjq7nypIYkorIncV7K0hraGeLEzj/12Jp/e7GOBCrNjA5ADsK0YvNMX74
HjZXw7K7SSaVrPEcMj+W31rbm466m32duEbVb0w8BNW0wsJFDV7xjHp4TeNEd8wx
oDGitd07bEn0/s0UgQ2nUIgQXe06l5riIgvnLUA7AUe+TG76D823KVPX/xrCOFkk
DKlTNRvtkdM/Jy8pzco2Wm7qHZ0LzV4dd2Cw6dHswYryODAraK1w1QadeD5sRf3Q
xcmcJJz36W7r0PuezKMUXJhOpqQH/LD8R/3vSuHSFllEjiuys975HNioQsRnLlLE
ujkousKq18zm6+g4eUGFwrHwrzhr8hORSmfpZqwyFzYocWUqLVg9BK2t5k5e0wbJ
Vg7WiT4OV9yj1NbD/DaXOYBK84knvyAOViqSYeAi+0DtBsqedK5L9a39/l7iovFe
ekIZ1tpcu1vnh+wBT5UTZfBLiiSF7IJ2Gn843d3bwYUFJETzVQBgy/eAoBTdjNjb
lveHahdc88RgD0ccYi6sYCRmgX5mfv/zAWLNtWomH/wmhaxGdZvFc3zuEJF8fuCX
NxCOy6KRLiPgli6rjKL9eWLv+lZd1iRYb73ELgqN32ngEwgEAScYSIYAoZOauPY0
2edd/IBVKwr4oS/Xfi08p632o81M0AFk+a91qBvqkYHFsN3WU3vEmppLbpWGguQH
qAS59ycMzFGxpDhmzd3MqTQzTaHt0YqMcNF/mBG3ndXNQHY/y2p2JiK54iVoc24K
szcAihvk1sxtwQJuOKFJT5cLrIC1adr9rznXsUzZ1E06PZxBvtWgEpd6eX2pp5Us
aRs0dsi0wQJzh6V82m4EghbXFMY2yNBRnu11A1mqPwGtXkEj3O+6HeVG8CO982Em
7qveBh/2B627TzmeLsXAdknR03w6ka6t6kN5RGr6lCCt1ZH4R+xMZsBDHaCvU7iG
aIqcuz2Bx2sSvyoN5Qa5sT4qCZ+0pnTOPbjQqc34PPEXFkdCoHRRNtDuRB057sal
kN3br8P8xa/o07nK3A22N7jC10y56a3t4xsPZgO7D71VCjd5LK6Hi1bKvqQfnZOl
rBHf8WYz+tNXr08rgK+eflldZ1lAp4XwIqLs2VAut3jqK00Nyr6VmeGCGG2cPxUM
Awv2+eGxAtfF4tw8JWOwV9EkPOIa6LNL5TTOp86s4iY5/3DU9K6RZaA75Bk9nVlL
PXI9g6mArLc67XVyzBD3dX4mZ1lY5jtvFyKZjWgqmat5jd9xPlnhEO2qFSsaUZZn
tZkvzZ3Y1ot6tkrlIGTZIIcnGI4Bc0c9MkMIbY8PrM7GQhJyRHE4cyDGw3gBHaOF
S7S8kpwEFwOLjk9iHwIK2H3vldUVYI1wN0aun+gunoSgu3fskX/zqqGWTQuNr72E
OHyJlzeYtk7P81jzZI/N5fDv1/s3xUXZQLveMWhxrt2KTtKZk9xuu4pQgA64M1Rg
iVrXhiS5hi9AxEiJeqzKRxg5ooL5owx0J21co6El9YNe2YqVER8rlr/EETfTD83a
DSGtiekPiXWsCClH8kOXEUAb3mX6RuELaONUTWzxnVJKxP3sLtgN06fCzeW8BJjz
DljjVQ/0+j47Ft0NrUd/cu5YWnWWrKctYc+PQBU+q8h8di5AnRz73FoYHrcHf0dt
hpp+YETmLmNI8EJYY2WJunqGBtQfvpCvalJ2/0LBInsYu52byLJYMKAGsn4P8U1l
YMR+0OF5Z9hfeyVijr53iEB9EaTiEw1TDsXIYYJflsrrV/VonoHdregZcCAeuYJo
MvKqrP0BvlUOccDfZgXs+3s1pI5lrGWzlBLZ69vienBlK1IJopnckG11oywzJXNH
B/uHSAlfP5TnvbwbDZKtSZo8GxGAVUi7m6Ou+nowFaFj9N5aainjUir38bBOeyb4
j83qqAYy/A6oIoY5AMXmyf0ZaRPzuMFFwOdCZ1IJOzKWeFvhcym1r3N/X/KlhMpj
xnKyj23oBwC1kBxtvQFnCv1GB0yDSEh8uaFTvDEaXZcEcsrRzgF5Z8ngJdiiCPN5
MMsRCEAQTFKe81kExPyGPFv2Rn4B+wE9FjtKbKL7ub+Wra5ShTAJh1OjnEm+RkS7
qHAF4vsXHxYIt7+KkPx1lhugmY0kdsom0WO+2E4x711yrpMBRTsdIig9przamEfs
nDXR/LFqVYyKaMW4tBFulcwIcROzIzP1r+UkGEZKog38N1Qg+9NTnaTQn/m5Mcsd
QK9jy4rcvsqOD7+Ko7gPAkMi4jwOs6sy9ggEX1xNijA1+3AZ6OlsrtqgvFyys8Ey
4EByIfr/F8wMgsfu6CV9AlWS7CeFfsQqzm67sY0K3pX7Yo7y3l+AkbuFw94CuozT
EAyA5heNeXSGEMcY3i5DqZaRlnjHMLPtmqTNOXw2hcxFtg0ifyRH1qpCgkrtwUwp
NFEmhhUiYjPhA/6NlT62s5p/skA+DiG7Ge4XV3sPxgG6EkjvVfUYWsNi1hWDht7l
Y460iCFwjVqd4hQ0nr7lKRnSD6fsEIo/00385xtdz+pc2xnpTmitH8/64GuqVpJE
8pnHwzPX00JoTEwSam6F8WBNjaM41NsAjQ/NU6D59t1nmvQ9Xvvwp1gk7WZbtRRc
kyQ6GB1Fm8jG20q9caeytDM1hWlJITlkkTQlLktBn9QHqkP2AWFFbcGVMdeKSMHa
ktY/xp8yt6H16ZrY0itJYKbjbJYrRdqVaaxCjJMkTFAyNcHJZ6rMSgcdENuQK4VE
jRTMg3USowOiLKYTwd4Zw/dVpQYr5PbH6V3LzUFkmq72lQuLBzdZkhayaDOXRqnd
R4EnC73ccF3qNQAsfUZbYiXbVJW/rZrqLCUgmWZxnGNGuU114WeTV5JqugBvMRYJ
3jpJrpO7dhYoS/qM1FS7SyYUu18mvvSBGHA1Dlio6EZflnHh18WebOw+lUibwzP+
r8YuC3v0QlsSgqAdSAVteiV2mV66mVgLC5OzeVPjwOj/OvCoL95RuU7A82xU9CbJ
hMwBR0IDu3UEsJxKl9Ifot/tAsuRBa6SFnJeZcsG86ivAfEeDcfK339r9Daj788M
ihg1hba8V6zF8IvOlOzRtDADPbsldQvnUT1Exip5tV+M9byaIOJwTXMbY77fpKvu
cOPNDffsspDenLSH+mocHGT7fAv4dVUBLtiieCfwcCoRir8CameatSuZXUGDJ+CW
waMVQP+goQny5l1dSKNKvL5XfA4Tclxw3TQMqIobOl0xZQpHV1c2Oo1yeAXoWFyj
iXqlluIXOKAgg36lYvC8zFQ0UAOUBkhttiXT+CvcZJR8LeKVz/oa1XaYiCHqy6sg
soIMUAWYzBKLEU3NHnXp6/c6vUE7KmVfKz7i9BZkJY4kyXb41DEbFkUJWhAiUsTa
AcBQ3mK2ENqnMJIs5xfLYX2wZ/nzLEt1sDEZWFX1o0pQrY2vy9IoKd0ruYT3GHmi
6k8GGPyQxj0AmPmdxev2YwUS8U+3Tcdd6vozCRWawljKHg8Piraisplbw685//vw
UQadV/UTJ9pyu+GPUZ2/UzMBEsvZmp6Sv6M4665t1RfgbWmcBEJzT/X3d7uUb9WR
7fbTLQyCo3jCEWF7tTNrTdQ8ihkfVjkkJEFwVTry2r0/tXp2Y9cs3Wg7mOT6o0K1
D1lSQmxm0NG/QJK3bp5VniqGWrDquirUlMInmugUw2ovUVFQYIZXgNX4eBSWsi3o
hf+6Ia2DMlc+8/Kssd29K3usg5Pklr4B8L69Nw92bVPy4X2NVM3uQRW34zYrtN2a
P5QIXTr3Xv4pSkyK2x5QZoXj+hT/HimVUxe3zp8BIUwfsGrRP6M6pkPi7+QxQvjb
2IprT4BeagQQUPB9OvSr9bYOdl2fPhf03xAyasN2laYQ/dgkmRIWUvDsMwmXkpLq
Rr9H43nhr9LzuiXmFK/YGIzhdAA6xeXnzGv2omAXde2gDHc2A8T5/JVfVuC9evNS
91RXcOJf65xDAyxfOYxil+rLjMs+2acUtk61/7Gq7IKR5Mm7zpCB7viuZqlCqQSW
Cf4pbABOUwuT2SDcNeCZ8iNODxRhsQ4HTK/dWhJPkHcIxajDHZIQ+adnpat4UzR9
wuc2rJvfnz6bbMiZ8eE+Gz1zUF8THOPNrS9b55mNNLe1abOgVlYtQr92hBDxbVGw
+kL3TFSgrNPaNlJSMmaTaLy33gL2jdg2UWXLrMde2fLcQliPr/LE2zsszrQfK/Pp
ciEqjZgodmb3tCuwZ4Z47Dk1iHbLXbhF8PUgmOGtiO6t2F07+J1wwg+oj7qhsBFg
GqCgjHIXKWBsn4jaUhhH1U6AUj+0VNAh4ZasMwkgE9Bfm0ofUCKIIpbjf/sADReW
laHIGabD8zPcKQ7mWpbxHdzGlTJDAwuEhwf0R1bJCWHJS+RC4Q9mIJt4uqN2o6Lw
qVOIFXxaIpkdq0Z1vvfH33Nwl82CIR4YS4J+R1MQrLQJ9TvpcNI7DSt47gZ5Skzo
3NT1O+z/4mtKva2Zfonveq5QF8voFF1Nn7iXVNdhA6l7LV4gN9g2j1A07OM7LjgO
YiuaAuttsBW6gU//tlD2AFeorUryZcguX1oVhaf7y7lDwWevZOrY51s7sfZyXKfg
pdN9vo/PHIEuESk54f/oIH8M772J3DSXN4oB8fdRtr6fDAY71A97/eJZBVXwCtah
yZpcxw6Op+sJrzLW+pZBlNQjMQlxyEo+05UAAkcUo83t8IehEg0UKXLCPI1SPjBS
Inq3ewxnJDPqEpDaRh8Ouzk8i6Tq5F4cmOIMzISdnQbPqJzoMKvo1sps2cPBLt8M
0Z/BFkqaJKzs66Bbumpxf9tRWeOfAG8DEugmwhsNQWogd0QhLOJPY8l8aki1vdUE
qv9lazezU8rXkvISqm05tRj1DOnz7Nzin+M+zpift1UrfGYq9aQJqOkKgSHOYrSx
urvbauCs09VViuS1fnZNSppuQARZZ0fIJRaQzetGbVOFDCvlSSXD2Q8dTns9zWxc
99Vo2rYpLgEDhnpsqOjMhB46Wjp/luAMn6TBypHWJBTrBuRR1sfRpGxKISKZGrre
4iK9+d2I3KKqeUdq5vu18YQSon77gBjBMZlpJiSmmzsL7VhXbAvgNGQLsFvNbusw
AU5doUsePxIo8XqwJS8vupXWO6k86cTjh8BZvlKe+ajIg4VhCXMH8pGQD/HN5cyZ
XTPX5n0wEafcQmuvx5o2uQEpZqm5glT5BfeZFZtZZKBjck/49l0r9s2e/a0A7yuM
ad2TMLQOXsnFyMEbOJNjAHx9NGZpcW8kKrHFAQ6ZmU1dntXXobQaumdtlwqtburS
MazpsOnYxL6d+RrBbDFR92QFnUsEFMchrpxVcqdm2gFAWSbaNKL2hTN+zU1ylNMx
EtwMkGBI5uZHMq+HpINMPBxSs78UDktXAP32Nqjh5NN3fmCngSvorU0LxsTbhVWe
J6jb+OzJGDt6EXz3EixWQnf7fjY9zzCQ3NUaZ2SMy8B+j2AfeFnF4NzgmzRmsUvi
bkRBMKgYfRqWiLyAKZTf8s0f0JWJIiXIKVlVSSqK/Ub30+iJgC1Tq9jPxLccGnx2
z+ZQMiIUX6riZFH+k+RcYRH42hQpyCb8IVfCQ2Du8ylNdiou6xHPy4JwecETZjYW
W9FW3ft8vjORvI2eb89Gr/hl2rxJGwsIHir91TMOYBQ29fNTanPlrZx+1ePVSF0X
swzWd8/6sfDrRzJe4Jhi8kyn/owQ7VMVg29QJbnjC5xPLovUhiS52p3Ha5cmG1fj
J41CVEWf0qUFJ+a1XvygQ9/jErmA7PvOK1ajSGua0otQGKeXDlHgCIgVps+q9+Ti
dlPGBvEgXLx4nCXWl7uB7tPm3trR1H1r4R6YKFX2JzX7ECMvNweqJdAFQJpM5e4X
SRjXyrGhy6ZcxrQCwVHKjBzgheE5omw/xytM3odEWFpaDdDsyCQLsWGmP2y6m47D
pXsaLw/y5Ab9m6nyAsnBEA0fPUoOwHnDbBZfnZLDriQ0u4ssYqrzwUbZE4zlcFtJ
7pqbkWbBmeKyJ2iu5YYIX2w5zWgmG1VW1cjQm/E0Y7Mh3KGPDkP491fVOCfUEAS8
b4sm50UU65NpXLrJPFkA/bRIQ1NDLfbV64eRpQahTT6bJ1SoBZK8cYDrF/zMCKut
Z02OWXiPtj/FC7HUs3MZC3B7qqmPfdSBQFPoKtkEgH7mFjCE1hvRNiAEohEaFpK+
5T/ROjVQYboM2smpRbOmEsGimcA0xyX7/uZGy7Cep2Q/4EKlKJp4HmZsnOSO6+e1
qCQmZkseNwCnNbhO2cUfglVLcawPaeDZXHfF86Q19skwXJqCX7bTO7P6IsBZvcD3
meRP/uoSp41d7RNRZELOeeqVAPHWCzSqaDS8m92agBbDOg3jo3kZ09nrir3416Ir
kaoNN8/+5KkIs9aZlY5bu2Oc2roI8u2ulk5iOA+cZqkoF4jh8UkuTIUMJ9fot4dI
azdeZgKzcb3WnWH5HhBf5lIpeF50Dx+jgEs2z6y63PgUuaerPwzDK7IQT/uiYgQW
Fg6hUJXDDxTTYlyzh2PWIFqLlx0o4A5dfhPyde65rwOFaGUdRlhrGq6zA8DBQueu
eLpSgLCkcrCbKP0iUGsE7Esllk2SdyKL6hBQBWOx6iCXcyZYQ2gYAUUNA0Obc9mi
5HFeMbQHnq254AGo4ZUnBj4pwlnS5lb23sFp3bDGauIFWYmwB38nm0SLNgbxkXlG
PyzB85nGcrY/EUcSRWs37g9ecmwsGKdOxqGGS+hppV2e8FJWRq7LRDHjwIWKHG3t
rzQ/PxPG+7tQd3B+QjQjz8QMxEkS2cCIsysFG94zOOwYfO6ctPNOI+kIDBD6j1XG
D0CAlAFIwmUYYzNHUAHvzMIXAPOLbDO4eRQIsQCRQ0uC/9FkuCEhw+1zyL8odBmN
fIiFw3dy6TZDLmP27y7tkMWLhlHKe1BaG8YgU5s+R/ypfA9KGF6OC0IwVZggK89W
o+oVFTA5NNQT1gEBRybOYJ5i79s0pSwRnu5oQnm3YA+XRkkRm7zk0h7D72QNs7Nr
ZUPN4W2nY4yJ/YmufUlCJUdcp3zkgMOI2NvMXfXs6J63t4Q5HRaam0tOnoFYsunc
KItvMlprawXmdrev3Lb7RoEtJdKqUP0O3QgyCzftDO7xUiOwZkiGgT+C4cjuyzpe
xB2msbn/CAKbBU5//ge/X16qiyF3mTnkE2wKjp2Pj+JLXUa2k4dheYbA0pe6p22w
qqgSvWiPe5QDJPdPpiEQRAfhNSGyie989dqYQ8Q63XZp80pzE4RwDdWNRRcPo0xg
oYrdKcvYkFdyXMNdHckDT9IJbkWrcz4ZxDZGLvtXFxdqer6OuSISQ89ub8cJWxfX
XRM2hWy+Rt0e2/VUzwyMmKgZvPGuyf0JnLQqhKaA1gpJDPNNin6fDbvB+dTjUGDl
Yw/NEdVxJ0fgVUs4LdhglYHFbiZ97u4G5PhSayStdl2K+1yriL3OLhVc0ukBTHnD
RvXUGBToKu8ixOTTzdRiD5WaCkTe2I3IFfeWjFYNnJo7LH3tVHPpD/yZWtu3p74U
95KaWaqhMy0onjz3E7jnAnjoo+tXcdXZj4DvYSYdxDl8NvsRgkd5Q79W5mFSoLLd
xLFZBkcuo31KD4G1QaK3areJ+OVuv4pr28mq0jugqioieZU12Nbi/iL41mwoDqQZ
FDzBcwjEJWp3bOw1nvwK1V+139TCACCWM5JwCK2xf5MeqNbRuVbEnQ09vWzeqXtc
EKoTHS4B7obdJMCN4XGylIblG6vVdYn08q8vkQqLt7pyxm3/JJcd7stY7tBe5OWn
VvXeoGZV4/PJxXo8xEqAYbPnUjM6iMP9Bp8zk9WzN9teNKTixV1tWAJ7wWfmXKTb
SyaELZhxeXzXgdWP2fSbxLG42cujGId3FxIUgWmnWG6jymgMU6+svSDR0OumL11d
iTYhSnrwEJsVZ91ytyn4Gr4pTEnZwKtdgl3JAB/05+vZ7gH4KnDqLZQCNQXYmvFS
9l/XZQDl7QJ3fJGPPUMqsqaFF2QmbhmKqpG+5h7pAfXRmqUJLzultHcyBrtQSEfW
1lxgkA5e4wXRsu76hX+otkv0BSm7CjYenHy7GQtzj+FJRpHT1KcKMfGPCWoIVkb1
u6Hwv9p+sqfEmUJbBq9K51TdQsZfO/PGHDtIw1qrthfboSP13tcS0hexZ2AEggxf
2e9FEeltct+iJ0D0OQLAjCHfv71/X5DGSOmIsHMpSh7oo5JNGL4R9PimDv3akCzO
/ZZizMhMz2VaLpy+U+DNHeHlmoHUG9Q8Wsgcdm3a4691Est83BEh8pMgRrEW9Z5S
V5CnlT7U1lNaN9W5sSfEiFFeJgshSimzDAD4d71BU/k3fM3nI71hkYrjh9kDPebA
wvuBb91dYFpyQYAZBl6CcOj5OLV39rqyfa8KmX9ZUqY6foMvj98x6siz0a0PFx3S
MfhAVCd3vQGgMEyCz8lB5NE9QRrbN0SHRuzlBwI6wZ6vfiwkme9GFcC0MI3jRG+O
jWgjrgsKsdEofQqwkzyvjol62ej9SCwjsL3mNabtW5HhaWRejO6T5T35hBNOA+Uj
z3FTcbLnmKF8PmOJQOosi6A3g/a8dbOrIIbg8R+KE2n4qaKmYaywioes2IANwels
oAZtjbDJ6lFVdSi8/OM/GqESmCPIUv/tQl9vHVyOhzlkQFkgHQlriVzaNODIy3J3
xYq2+rTtgMRNehghKbTbJEGkONX1RHfY+ytYqtRzGbJYjw1DJTpmDXiqadx+vBI2
GTqQlJpq2Qk8xglJJwK6gOZbzkO9T2ZrKO5op5tJ3H3TKQfr6Hdhpo9DPWo1cnt/
mAyNqDn3qQSYahxRJyC5x1w2iN4779VV/XwYSCB+T4hBEt0/ernP6vdf1jzHPksP
wOCUKtcflGSgB16MA5YhCVCSD3+WE0rMUQJe3g2f2mYMkNwpGci3InsQuRdqY0n8
yYgUNZ1SW8skAoqSVCYSS/+6XsW7REDw/+WEgKl7uLJaDh+oGY8HSIjp776OSbwX
uCTnWrOYHm/Zgb3qxWdEEDS3/DvKav4erBN0Hzm/EcgxlGpGaB1wcrl7kCZLAFwI
3dMu2RAXz0nl4xD+lVhQCPsAKhZ9WspZlyiSF8ewxJtiZuRsSYnUb7HEILCpPKd2
7dWQOmOcAlF5zste6Nxa1DAyeKSB9r9iXHkqI2UmdZiihFl2jo9UzzCOJ5rh9iNf
dRzHSJkNBudnjO2B9WvmVX0KtosjlhcCU0PT0tN2pqdsfNtC/FjYFS6o6s4kQ4aW
zoJDCpupFtLsa1n1etApNgOdLEIi1soPCOsPqAW/NhpOYqgidBchdJWcIRYIoBv9
TP71EU07rY9rDY6RGjKs0tF4WdWeLHmxvCUFCXWUOrMmf5szEhYar4FesYLcqUro
8Sg/V4Dt9aQZZ/COqCHmzw7zWcWSuDPIdClW93eOUVzfalHak+Iht3HPrWvSJnV5
o/ugkMAZBRe2dOKcjreyLfyhrIVPMriNdg2qPPp7Ud3Wf6vEja921h3JCgoBrBBF
ThndVihx8SIk305+ejinZEQwplGnDlb4s8lM3KTMpr1GrlLQyG0bUqag1jdoHsax
IDgrl48qGwvWFP6kTzUADmXo34Ja9MQsPN5rGGRXT2LBoxwZajfNbJyxQZUQeOVf
rlEX4Urf5QuzU/1yF2YQjL4aBtbakZFa3TxiwvvUm/brV1uvNLO8K2MQLopaBAHX
oXAqFw/XArTI1LK2E4e5UiHQgOiPXpb55GoHUEagpKLC3pJN5ztI0TrEDTBmRZvY
TjQnZ6u7Weq4sKdVpQ9T7LOBuw+hZ0Jh1LdhB6xICn/vp++CXmB6j/fUGoiiWuj1
8fyj558YgtTfpMGyW7UdNq9Z7KAhWCHGWM6vWmHjA97x2QL62zqw/i1+++C6R0V1
+RM5bEwnMQ4SR9H9JSVMl4fOTtxTgA720lspMG3YHaBVLyIboiGIcBPKD8AKDfjN
d2oGlMhvpFzpLAfQWmhCf5kV8R1IkXIe6QvZuzgk9i6I+hnTtxz5ipfKiD95xjj7
8gSTmRrhOmbZTt4Utp3KQ1N8fxF7RkKD2080rSEEQ4eEcmrq/wMPPFxnW6pgN61A
Qbk7ZgnwVTdAE8A75spzgp3K9t49iL1b0zEJWgyvqC5o8v9amK11qqaCQvxz0EF+
SdvH+Ymf7Go/c1SqdbG+5fwQ2zbMKfLEasgfQNHYcSIrYV6f/nguszI0pZKZj272
7WtXuAxE41QxPavjGxllNO8Q2Iwqjyq38pLtKJ4a0gnuynw555/0+Wo8E3L/k7zo
i8GijVG9QiKZY5IOfuVdT8h93SuPCEexBn6H57zO4ZNTcYrF8vvfQs3qKQ7NOJnX
MSt1MaCcAt7l4wQxE+CZQYYx6GZ0qSa+r0agJngGbRvZgoag/LUs5tOWS7X995Mj
ChIDWM5189oQzgSK3//YtoRhb2sskASbvJKP5E8I2N+ST9goeYQD/winqZT4VfdF
7nlFuTurg2w7My3KKuiqj8zZhGnGrPynj8vQdthR8c0r8TZid+9jiM57cJLKVMx5
Yj6X83lsVGLh8srLsOR0IsdZm5wtR6wftad+2u19VF6gWRto0dT+oD0Uxj3bfPgF
EalaYUwedp31JY2oc4zhasGgvGAp7wDYaow36uexxS0=
`pragma protect end_protected

// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
rqjcad237Dy1hsniRz4u27PQiMiJ8I8tyR0snzY8j4NTdrDdFIoEJPJL5puxPJCLGOGDLTtRu5wk
vgYdVw26tVycqRA44ddawjmzTuOggeg8a7jtFtorBIaCEy+4nTK1f6qvMlwLeZfEwJtP9+0JiNjM
MUttYvBGh3flPFH6WAUXbL/cBf5jC0yAXdcCRjcFTnGXHmCjOnh5poG4vcLVnTjwgtoyRXPbiGgW
wb3k7SpuuZyna7ucrCxq3blXjsXQCFOvov+TCWc9TqvBE1Y6w9JrBilNq7msNUHh6k0zX+vDo0vq
bMaUs87l6gJbCz0MkIwupKKaN/RaJxvl5GI9Cg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 36912)
RUCx9QfH0gGO/ZTFFs03TTT7cFTVJcnjhDC5uB86k2m4HDM6ks0z5tepRMIGKIp1a1a+zcjhUM4r
2I89zydT14L9pELtTmVU4QK3K9A+kL6oTEwGf4/uZPR/r6UQ6Hwfj3/7PdnEdl8VTkbyE1X51u6i
L7sagaqIZs19XcWt9j08nJnQXtza1I4oOw+qbShUhvhqLwVPBemhVOVraOjo04sjTQhD+ed3UJ9n
6RA/cwhIRuNuURLPd3Rn7J9/kF8TtWuzc8o90ZaQSVBKEtXj2jgVk9EfD3qogcEQegdJ001qLumQ
MDqqpSt+ujGtOvtO4V/a3jHLRoWzWQi2jpjLHIZR+95Y1qqBClk6hFTbP1SH/JNc/w+G3H6LdWw8
b5bxzten0UBBqUXnwvgAv6xIn/PaBo9GuQn60Aru8P3XODJjevQQFaJtYCh7F0b4ILhrAiCMzaK9
EGMgusF+AWu8pRD8DHCRzpQ6MYKqcN3O+apeulkBCq1WlxQBHn0daSKmGu/+F1f9q8KU44NpygZk
izmKJshXUuHldDp86khT0W4lraa0n442JFnf+x0evwtllQozvleNVR0lKQoKrEw3LpuC2yR1cYPx
Qb21Gb/nprgGR6bgQbGlKaEDYnr0cWFCxJb/8gVUlw5ubCTe5Ob/WP7wsRpaODQ2McB8LGeJCYh4
wCOMEKtV5hMJhV4sfXZQuBCPbvU7tdnuIAXroqHnxESrnEEjikrOE4AMeb+hnjp+nNw43mTp0KWk
RbFdD2Z3SNmfF8eeeM8jgbk4Py2iXOAnr6eOVnAv8TJ/D/QDCG3OXCeroy/owXu6/2pl5V/LEHpt
ILdW3ant5FAHnknyMOe2TzqAVtMOYCASOMqHpy0MUusRzruqeK57dJWL6BytAZZKI0XVTsDeX1Hs
LE1FdHc5eFjqivb3TtW0glhe8S+g55Q7HYlUgRaAGOVcwn/V4ID4SFER33KFDwQNG1xprJboeRaE
VSSJtYfql8fii+njDl8LpQpV/Md63Nx+5pl9aXs45A1rjVQsA0fN49ME9PGQHGa28mBQGtLxcyij
q4GyfIf3M2mxU9ovcBSPOZMVOdt9koSy4HXV0Dx2Wql85pdGULa+qECSL0vMKrYrmuS4wfXCnpCs
sYCfgKQmO16aoT4YMx49d1t+DOitLzothPHF+HKukk/Xt31fGFLMHm/ranRuk8/9C9AmY9bLOeWh
LZRCVHf/46a2LQ5j1pX/q0tFLoIYRL+24/ZgaxEBEQg6+HmGu/hXLcNtSAU7SaqTzONtjFgnN1bp
0ERfa+7edIZ8WIX9E8k/DARMyyiWpleFVRhaBmaKedpcnFhz+nrRvtOXMW45aqyU2mLNjiu//e6P
zcLg5uVD2AZiqHU1yIhC2lKrAax7B5IyDNvkalVp+3TRar7eYb87wIQ4WXQou3vvkUkRGoX8mq0Y
PPXC/0Gn3/Sb5ndXA0V8ZycRA3YXysXQzUBfnjBkLiypgCaT2l4khuAlPmqb7eOxlGmJdFhpzAed
klEmCvSCJPs6ijQ4YE4mZiG+nUHWHtTL3QZqrHOEwK+LY37lDUs1qEaKkW2whm2W4dTmzqxsslzM
Vmq9wwmi0LzBhWZrxPErEeGE7ddI2oMbg5nuJHxKuq8WcUK5WV/jUpEvkKmdK+4p1oJV0cekm6DU
tj9FT5OtWWH/MdjXzYD+DzDICCfrN3udddORq0Pcmr63mOV3fQSzJYKLuEOrc56pTqsJzqcDQIvX
p6m7R064WY556TKIMPoBvbp3n6w+9S77qG1fF8uzn5tb83SxWKiVL0e69zPvFXwX5/YWDYV1EtTH
2u6JhnmwnDBO7G/UQdLmTDkPVnQYV1eJvfjXeCX2QlX6FizjeP0eX6LmeXICeaMDLumlCnVWIgEw
ijX+IDMijBXH9sJUngvhCXJULPvtrnJCe4qmjtQnXWHxkPyXYOMha6MhpGwWdx6JU8CvTgciHQth
7Xz2PS3eSU64DinAUXzs0Yp+i1JZ7lDNZXXZsRLPjDD0UWMa9osXbfQdhKSMmPPXLHxomPhQrEuc
mi0makMwhRMpgIozu6eshtRCVSTxmDFX1NvJkyhDFUkZN5azeKupq+fLnTiroyeGGnPgm8Ex8MYP
3kTxXMMmCaDAzzygHExajNjdLNUjdJ9gBcQFhLPJNR4qKFlbvaL0ovgX2R1XE5giDtTVejW9eKT2
Lxj77yYPOricKszURWHlHN96IdD+CY78szRH0VV9zsBXmzuYR4/wFnpA34o9c/hT+IWYmygae4T6
iLfmRNa7wH/1b1BWAwYS9j6+C1zoAfeSPFjJNpzy2ExbxRLMNbmaDVinqzvlSHb3zNIWQ1FH8Mee
lOY9vfcbsLK1p4hbK3N27SJrNd2nrqtpVBvZd6ORwr0xZQ85fHRXf24ocDrlRRKvT/NKz/EtHD/z
FpzLVdAC+s4O3CuAn3tgvKg1vc1DhstE2Z8XMDt6HExAsJ1pKZYJwh/RrzwBzFpq+3FtJSoFahl6
A4e6GrS1wJExKjnN+gb+omPTsGmrkbWkNyFPeRUaIJNHKbwj+Ev1M35+wq7ECLuxJOLSpCkh0ROA
s4MZDzBBdTdxWodY9TWPvxKkPVidSIlbp6lzP220dxrzLtbsgyCcZHVwNC/imbNeKU742lsw11Yd
pjeu+1E32VuM7hXy8ECqrqxltqtpLjRMl872Mkk1zEB91opfReWjcdQDSDKB+N5doOW2yz+hq/VH
1vYoyETaTRKAX4EvPwXuvGfkHz0pASTs+cHCCiCdTCltU5f7kc0CN+5Sohr/IVj6q6HxvtA9P9XK
CFx5gg3kLOpSAozPH+JKVEFaa/Xdx5xFPpv+kVTtGDOiQvwN9Xlw0x9oSYDOFv+X6ShXtIF+XdgA
TLOWeKp3J9yIJLkMEgOFQWxGOm6CO5H/hKsZ+uezIjaly4wkRsk69oEMH74u9yMjAGhUyAcYJpkq
HilTbxhfK/lsiGcdfB7BiShIv0WjLcWv0bMzEKa5aTJbt5Do0IvosKiebRYeRUeWhbdxCFqeSfxG
PHLS/Y3A5GfD6ZPDTUB5JCGBEOijk94rfrmfFzeaO6VtwbAVqm4KVeITqM7PX+zwH8WyRnjrUUbY
UA8kgDYO3sYrD3EHRwYd/oi6gc7EWwyCSKuDtaux3bu3Z+tzzPL2igWbELpDIW66gubhKOgZqjPf
fHGh78aRUrr1xa2rRwG6ALDi9GQmj4gMVBwjS8gU94cEnDGezqYHFyiaRTiSuZxNH43TWajBy/Ex
n74kMaX5DgjhtgtpKpTnokjWSPcGlq7GuKcMwKgoYdV5KqYHZ9/Jn0nY3IgZ/L4iMIJNzBL3uaiE
2Ci2GPiSYGuTL6iQXFdwfwj0W1HS8tiO6W58tZR/IGeOMkFo4WGFcHJL5J7fQEnNCTbn4f/FtwMu
J7APdWlICKlGzdbDJLoZzb5ZEO8jzJiTccAtMJqmp9SM6F46999H5JtlftyWBEjVSLWepPunsjTt
AZYDf2d6zHlWfndqIt4B4C3nobU6GLV0LF8sMSV1y2HMv3hRVZ4BsRRtoVF0Bn8tqgkV744ng2lJ
0/x1NDClygwt3ru2EaCsXIx7IfQwIS0FPjgAcRAGQKhVyCii6m9b4JT/7vc88PiNJxFtTlcaL3ga
AyjJI9y1Dt363BGcRtdjlhLUsc9t0PLivi+c+EX3FoHBSvPujnHkyMx7r2S7gDWS3J7X7l1Wi0V+
fbZ5OvWwkBVkHUkVu4mQJQNacOGUj8rGzz9tPzICoo0dhD8cnnNZx72sZjOd3COE5FSURbQhAxRy
hp+4iwbmwjbtxMiG/S2R48TYlyEfO4v7PMG931VxnZuZsuOrDsCScJlGjtfJqs/AVsk8+BR+CzLp
oiyCj4EldDLUmPzMHEvF1a6G7k3yqzYwX97VU6nHxTSna62FNnXXFl8HtYzBU5/il7z8fVwV0Pa4
TzeA0LcaMiG2q/3C4+RJ8bKyHWfq/SpkOw69TkOSe5wBscCc6M8If+cuq3FQYk4b88DK3dqQ71/F
0LG/LQX41veZ6DCKHKezncQJmSbjv/gLDtPFHor5PFkwWKJRSiVwjKi5GwRjFAXVsXNFSckn+6t0
0qQKFjzi13hSe0KCkJBxF8q+YxmrS4P0hxD75BYHlLrVXLGVhZXpGYJHfIrfDXnIFJJ0lKUbPzq3
+/XgJWfQejT7RqWqGju4PnxPhgS8dkANLoHd2itKuZZ9iwqobOHlJGTkPP3Uc/VXKaD/gXp9/svK
cj5C5AyIOEZywPnR5g7/eoBV+Jnyd/HRfb7eqRnzmMC/wifXtTogCdVCURfJKrNFJhfT/886+Zha
bXemXwkR4FzFCZo865sfkuRPbCkQ0Vl8S88KpbeI1iyP8H91Vz3feMaig1Ewaf1WztccI1yR8Ane
iNj9V1BCIptdJ+FTxA4D0BBE0uoKqwfl1567yQdrfHHV47Y8MxiJqAONFYkNUpXhpxYcnUkHdnmi
7+39Tofb7pzWfA3d7audzFgIXjyqwHwION2KVn1VzriWpMcKgmXo6pIxXHoooy+hLzzS1kiTB1cH
vyGNMknE5F6JTJ0w+Vo7OSq1ydkyHzeytlsbnzNTNvYIZWxEgD3MIyAKGcKSwl1GzK+xIRWAEbe1
ET+gZsKhV9AVcn9OzQEirEuYGtMKrKosiGlwO9nDniQUopwGM8q02GZvuv0x9uHoOHHCHGwBqQZx
W6VXQTosQhVHWTnqqoGgqbfntbKBD7B7bTjPITqFuHXMQ4PIyO1ReJaPHXjTjDF/Ly5lJCgZQepu
zOZf/ry5QaFYbqF/JowuiZns9pOU9np7KuLsqz4h37/Tp6+8GBc2p2uCqrOCEAGLJIlgcazEn2mh
OTF6Qwb5yykpSe2mdCv7MDFU3zHrB3In1XJ9nIkMR2B9z5KKrftABmdg28IR5bIGLV70Ps3euDqV
29miO+avLMD2l59ZqyJdkrhCDvWaGWI/fW/o2yrhLliUqQohfSEKQllUVpRoCEpmSE2aMh21eNtV
o4TXpYpkpWWHeyKk6lWUcsbftYk7Ey+mVhZG/O+xm3H9WNR5fU73CltGwagPngaO6eAqiTlUF881
XPNTcED5hLhCytKf+/khliuBMoIMMOiFO9nxDZXQTkb4gyPTRPnvxNWTMsA7MJKaiMPkiU2nerHU
VC8q5L/en9ojpcUPjCDzeHNbj+xn4G/tBh3S1jd3XBMibF1nNPkLGfn7AEEC4cto+a1h06q1iitB
cCTTk1FWSuNknFgy3dg2btJfb+jy19unRApSRC0HIOFqkrWer7bONLDSNqJAS2+0k2mpxRjE/1Yw
Y3KOYkZ2Ff8RpmTFBlbrwKen5YJZ17uVRIpQeA5jIZwsXXIDQF19zhLxbpj9eifoRXEIM2H02fCI
fCrOvTm5LzjyxZgk1TlSlMLvNFEbCm8q3+nr7c6YLwJr0337r7okjnVEQRFwqQrAFeVJmcQktu+1
dOcKXta172Nydp07jrgLvfel0vvvqzKuDCREZ3RG3kOtbQeiKaK/p//Vyoy9RzgyMNgWKzgdjrfE
h/RTdBBufU5Y9jkPv/it0ron3Oo4fFo8K0N915ZXVe3S3iroT5nb+lRqupYwSnOehUz+nYn6bIUj
rqW8FOq86i4SBhsK6EobPeWutHIoxQSYV1dEfXl+b+u7dp9763fbT6ssT+0Vb42zCTGiafupItpx
IjChyFevK0UzPKR9fEeo8GDqoXrHNWc43lGjooQc2Q1sXLn7J9fLg+5TG/U9jiJze6ELON0EzZTG
KuNnvt1n4LwnkBqVeunK92K3SmuPmz0V3SYXpFFIQN8EnX0lytTtcWiu8y4ijg3wBMPOdh1N094w
yP08I8kjWmaQ9EPJznNg1vGNOSzyK1QA3FglRv/pDH3k6K/H25UH280xruF9iph2+uY0Y/Gvclbi
jH8kTJWZyrhCgnHrHPdmcrG84g/zuCeIcsgJLRbnXR4Ia8tXcBwkKOIt0zaFFsrH6k/DkqEpAjHR
wThOT4+2feVxT6M/t4dOydq2JijbfiLFDJ6wfwH1EJ4du6xRFPOdXk1syT6WXnKE0GUAXnTKAf2i
H24nSCniHV7OwCOiU+iaY0mP0JrGmWwtQzuTsJ1Jg8Ed3/VyIvq/8jKi/5L7brluOCuoDNdB3Cwn
en7sK+pkeqKcykZDB8cjnO5o6ezllnUWlawB3wT4686FqNdw+dBdWjH9b/XqrJbB1TE+8jE/RDdv
i7lgAX9fiypKHbrGL6wc7pJlksXF4cVZWkMlQ3PwSL5qM508cP0Gt4hAZuIiO9v40K0l28zHD8sS
JQxBAwfZsNFov/U6eeMXMp+oo+E2TAO/ABnYVigF6+oTeijwkKH2t6I7387t7Q2OvSQv2aOjuHAP
pPc05hKbzgZ0r16eXfNr9VSMJtttiFyyungU+MeX08VrwwUE93wpzOrimu6b8g4pP9nJYBFmo4+F
y/pK+uS+lINNOcH8Ybqk+g8sVEO7BI3ZTJyzSsc/NuMNlkaI8KWuIyyTri9HY2Xxzhp2QhSDAG+Q
ehQ2ZzBXHCGMMRqBeQxPa4Qm7x6YzMAQEJbe8yZcqMK3V13QMkwpPPpwn0i/I38jtaiaruvb16uv
4X8fgpe0JAlwCUX50EEusvBAXEKON7nBydRIGG/a6AOzig0ZZdoiFtInycTu94QzWOh5feNUa0E2
1FkPZI3pRyNxsghaHQVZtd8rmSFvYqc8N77BJFJnkt85gDAOZ4BIbRUpoCNqCzUJzde7ahtL/SNs
V2g6BOiiJwoYkQQvCcBpU1O0FTUxCDftJJJmwXq3vwxAdlhTvMjdiftS8KdnrkV7LthAkzDoanGF
PmhEAS1FLpw1g3uglV1yu2WuneqP3H6K5PCPPrSwlEhgV9WM2QGxaaxbgUlNIF8Gbxw+NnQreLlj
YHTo51xsJk11OUe3wyGXtONVDZ1ftJo/WIWwVDUJNEDOw07QANsEpgvIfQelo9gRMo8hBVw5NQ0E
nw6DkqN+JUFNYkuPVEfWsfJb94GHD7kpr75+FRsKMMGznj8Wn00uilBxa1Ff8Dtaaog+6cC/agTM
oIep7cvLrJq8JttJBVH+tBkAb+EhihCUyt9s8un/MM+K8S+aGvqZl0WZ6zOBMJX0sMdRYXHepTZE
tSkJi2g698fRHq+hEInQZioN1UWCuvqdaIn334xEVdXG4oLlbn049UmoEdfLOxL9wMoqB9ELjoif
jPVMMiWubP8Wy99TFqFIpegfHofxOiwBeiDtTQmKmbyaBOGavFBOBQvMAT/+SniNDisl8zE+5hcn
ksZHilM9w9zqwnyaCVN51bP0J7/e6+QNFyMncz3AjfcaeC9rdn/lkmlNA+ZqNATy0MQUujzNB29W
JG3rHzeJ07PNR0Ala/e5/0Ee+9e403viHYBVX5a7LoQWqfpfDv2SO5tlwb4x+rU/w5N6MB5RR97q
u+SHQtcY8YBwnFH1y5i/49SOIMngyopIsczvtp9LXeU2AFiLJymJDb+Rs3oY4pSmvPr4ZJSuPcs4
FpqNnbMYrUB5VxIdCeDFpUKNWaz6lw1GzDtQ06EpHViDZjdmh01EMHR5O4jYo7UiDLZgSXbeY22n
u8ebhpEVdbqfTtnjAGZJuGBmvhpIv5AJ7vifg+3LcbstMq4E6hhbQ49rkYs8xae2i4ntEN/Vlfql
yIP5asPQVmB/inMpNsLgIjdXV9QNQVYSiLcCnx3NYfzlqwj1IFd64o6VvqFmz0TkCx2g2T7C/2VF
ltWpv/f8RJRKsPi5CwO4fKSpTWCD4UUhvu3uYj2ozGbDKTN7EgqgkqhzlUXFXkx6qxIQPv3pCNJe
VgXy3Bwp0Z+NeFphKyjP9Tcqk99RO7OJC/j7CAcgO93y5P3FYjCBwUr8inK/IVxJ8Z27puuWJ7xJ
6FMo2gEHYUXBITIgaLFwT3ZdaU+jfhPHC0m2kLQ8gXVJknFyIwwFGMeqVQXov3b+AomvNzhcyWga
2M7IotyoTlKXey4t2/Sw0EWkG+txBb1crxnYOchsXxxUWBmRcSEvUmU42j8ppcbsUp+f1R+mJCic
3dyq9G9VIa3ptZuh4harRtvfr4KbzcMXpAMi6uis5usLaSKs21gVDdir90fl5Sxgoh85Ppj4IkGl
++/3aIecD3fNmRDcTiBU+rRt/tK9qvEAzzxdyK5HO05hFtRON4RAP6qr2IK9YNL4E+eRl7hHxwgz
Bpww+ePeIqp3CrCH+CSnLWB85qJzMKbGHf2fci63eCpdBtcTv2H+E/UJP4nCKe2H2jXh2e69WSL8
QvNqXjh5jmaDV+qf1ZPnlcFGR3CGVPf+zqdqM/LAwaGtZf7tmf2LZ9AfrZd24YGV9VQEHiv6Gbqw
9AMmL1Xary6TPrUErtIZyoYrQ3XDfcxsQdsrjf/cJzjqzo+YwQNkxQ134oPHd4BXZuS0GlWaxjFg
xfYwyCPwhOUqUN6XKO3ofF9rwlxerfQhZw5CKXVZ8sFB4Ng7sh6jqRM7XxQF+qNu9WqkG9t2/q/Z
/qioZHVcMPxygdxmtMzqt6XoAXdECCaIPTLMLOLwI27rTI63mX180CjYf9BMuOuOZa8HNf/WbLVI
odt1NRCs/iw+R82zVarqCAx+EvF2Fjk6qPVdd7LOQaKFgJVlbt4ONlOC68vwd2dk6EmYeXuJNNWM
uPDAHPzOEXEUabrk49YtS1c/Cjy4f23zhNJZuXNT2glws+zAmKvwUvh4uHftwOOf39F2nM5ZleaQ
ieq7D4J9yhVDtummuTtMb0xqlcZ1j2zc9kDyMnI/hpXocRxmoLDyHg7f2+eDOU4HFZwwsdZY31bA
n7G+hUj+6Ki1aL0b9kMo7u7sVP+YB8yzE30lWyR42rEqEDVsZt1dyeFqDkkpatmKLgK1aIaVCdql
jJMUULeAfFynEUasBDlklNpKTwau26x6cIEOuJ7ld7iJRJhsxnnC+oCRH1Lx17L5RktYTgSafKQx
pKFG2nBGemcwcH6HAQzNrEVM09sAeFNlL7WwiOv+CftWoRoNEz/Dk4vpxwFkFuwHP43f7f0Gk8Nf
6Z5kooefdtL2NuXZ6JvLh8iIZ3A42JT1Zw+2d0mWc9Qie50MqCeZ81GZ45RzdN9i8UzP+QjeSLPS
fEW6Qtql3eYCxdtLm+ydbUZxqe+K7xxuCe3kf5lwjGqEBTQNRqpPAOKgp8OgPY6o3/OZCeFtXZNF
+I7wUslNdBsXjwUptgMaLGT7Fj7LYWVbqEdvnAyvu2w3ZNlsrPLly0y7YQMDvtRha4uGCRs69sEi
inXJWyBPzAGZISzFXaZtfsYa9saWtuDQPLEYzo+6dcvGI/ONHym1gkpABjVI/b26bpKcumS+wG2r
WCZZqNVHqvkgbJoLYanu3VisPoT/JSXHGspDAI1NqSzx2yjHmF2rrgfxgMLRfX1mymX2zHBKvbxt
lsOcp6ZQ0qtzo5tXDEfxYd3a7oRnrjU9bouPnHSntfhkaajERlzAiQoPwl7altMk7F1MUML1unlA
CVmI1syOJKrKW+4FZ9b+wxtT6FHmb0uuwbB5W62ziGwuw7UuMJZc0M9K8mB/IwZvElvAqRPljvIR
6oO26cAsMAstC3ZXqUIR32MNnpQKgn3suK7VWM3tIVJz023XkCRSWZIn0NGilldCtwu2mM1OE+zM
SrLeVj01ORiAEuvZS2C7O6+6y0A8ZMN45S5z8zoV8YkoLasaO6inKipwvVS/6DWIfSwFHrhs18/n
OvxCe09JOs+eA3Dgi0kL24qof18W7O2W6lDECNyKdreqtknCY4q0CRufl2vLKVG9QoOcJcIyKQ1p
iAVcWYQgIFWdJj/7EBJtoafD458lJnsFKvD6YeD6OMzQP6GlSS8qTMcKZoDVJuecZoFLbxjlferm
WhxGJkHdPbvaRtJM/lsncV1AsPUJnne8po48uN5SkU6NfSDLBbQEVrSq9wQGS4JKWwUlODkAOXbf
GEbMjeDL8UUfmMxDa8RQ4aN/tQ5wfez0MdceLqtF/QEcJ07EQ7tfbktbHm30v5cwqiUqzJUYb2kS
uIKGcwboJkwUxebg16KZfEf0X1zfWuvKxrnSZpGR8j1UH5XCOV2rfykiwTen+xXdYoyZYzyl80Wi
ja/NqDt69TbT1VvuKl2diFZoDnZXvhkkEHea7ZkXjXJOcN3GPRtX+24RHp220CAyuhB9vQYR90Gr
H+ZNbTeobvQP9M5r1iqjvMUHrC/OQ8Y8DBkXs/pcjfXnGey22SlMpj1f1PvnHvGXINNv80kVrv5D
uHjyMLaeM0RadJk37hfreiCqfTy3lu+XCNiBCWOqYns/WdOn5VckW6udkF/feGLZiiR8jd1zhCso
jp2znPnb47EeEZTo31q58o/KbKi7kO8YZJu9Z6TWHAlj4l5+n6FwEVLTt8pQhWaxvUOqmC2duAAk
GWquZzNZJ7kaCo8GXyqF1b7kY3a6Xh1WqNhgsxShWFwL2lK098KWEUD+Ryy3Sd6Xlwpo1UhXDizW
02NHtYSFTGnF7MnnxU89p8aK+KkLCmPlMIPml/kqUvDULPqKotzn4P+1BwJ8HaPd3fNs25kl2MUq
UsczBc52ri+2nxn+SU1Lzq8GWReotkRyV45Ves7VqHCs6ImUOBpv4iXQsHa42w72NoTiaTgQBqm1
G/4TVcl2NGnrCyx/Hii1Fj9HFTNth8UDGCaiBN/o8xPBuXRz1af6qRJpOZUu6XmWZZwkOt4GzMm0
wskFa74ubKE8P/uS3QW/QGWon0GhyxcjNELMYuxREdueTSRcfG38xSqHiVQpXxVtbYOv7+izOIJE
SZnMpC9ojDZkfHCh1Z/HsBBreG0VS8rGojh5iZEx66FSJ8DsbG5TvgIq8Go4n730oyUI5i1zfEIB
xpOlv6UcLRRVywks05B2yp6f2bWskY4fknymDHA846kr1zc85C0DXtxC1Q8yo4TVXdG2W918vxz2
aOdDPZ/d1tDLEuir0NZZa+uDuA/EssTCDBwSqDrq979x4AJRq4CoL+TnLimdIQvWBcRB1yiS2HF0
OJz4eFBC63LbxS24Q9tLTvPWwUdognSqGvpQAI41ll4AMXvsxB5A9eKqPXexxxjOmCpz0Ri/YcWv
5k01PO73Ndo0prWoXKI3LB1eA+bgql2nFBNDn+DniwmmLTgXZkZVb61fktOVfjXlWmXsyO44RgUp
4CnrhObm4QIymizgbJqbbUKHnhIq2XZq6Tby1AbVgGba/BBS4lPxPXYRhfKjUwF76EytXph5m9d0
LbTdf0g7gx5LoUW+eQl5oW45xz06KkWzA6DchWjAvvEzoV5xOtrxi7Jm6EOiumW0rSD4HsXUJv5H
MrhnZFUlr+aT1t3iaQWLScV3WMiDrxN1f+PwybDaw5sS5fambdIBmicSivJnNi92W7BFvIayEkZz
Q7YTaGHCkv3esTw3ALvxOBZ3eA1WJ0YGbQUJFOLpQbEzHzzm0DYM4HE5924MZniibup9gpfApthA
3P2+MIJFx9KUxCHXygudO3n16nL92B0h6bVb9vmR18/whCNXK8WDlmg+XlnG4CakUigUCHlQ1/Je
Wlev9Xl/Korb1aeMhz/M/csN4NtBqGNuOcDfG4ojlfZnmKYtKFeXqBBGwMJL8zuittdcpyCFzGIK
5IwP7Ig0AJ/rSDx8xHgaXuFE070X/amEWWzgS6uans03CK6UnMS5i7iOyMY2qU/IAlPNGjuS9G0c
asKMXt1MtfJMCduw+glQjNO5kNi9rKvZAJ2focYOvWszbXfDt8xcxAYBphq3/XNjRD1TmF70VBNX
i/sqzaQNgAw/V5j7qteRk2JblPTKk+qsPJDwnyRW80OBDnuHb4reve0JIosnROYot9bWsWjbRqpR
Bjw2nSmyu6MrngqTlTfdZ+cUwJ0sc/lWb56e0H9MKXOpQhJ/a8XtRVuNgPCwhXzkYVCHMRBWxsZ7
cNUmqdXwvunE0KFtUsO6kFSf/WdaD8HKXAgK64rxq+zd4Qts2si89OuIs6dPoug8TiJsuX4ocBHr
9dGidsLBsETlaKdYzHNTyo6IIwnenmGa39rcVOddiZfSaVUmK+4AHDeW0IIoyBtW7sVWM6oNAHlR
Qv/Rlvke4fVHH1kGTTaAOuzJCt9YIqvK5MeYAoCTSoGKJxOvQfB2oTUEo8yJqR0n6y3k70fcobDf
SI+dxjpEE595lUF1h52VmnwNFoLhmGjw/pUluLUeIUPqUsOXYMYot+8ERw+CmwDYQktBDdRZkVkW
wS/R/Eqkp8sEtxAHrjTSObQSulw6TBD5D3ZIQgCIo0BSGpzo+0V1S2BiubpwglrfZYRZMbHmiIFC
Tsm+FR4ni/QJA99UzKrTHwxCkEMgStLgQDrKj5yAZCmRl9QKbsSE37sLixAoQk8IGvY/lJ+BDqs9
DaX7Nki+hwkazuWHcjTDhqbfitBBlykg12g8W5p1Bpms06YoBRnkNV+3h8gEZY4Vj175GiEofyT2
W6v1nXBYXnFOLTSxWRXLiNKNbZ8z7/ZfpagWXm8u4/4b57R1b+siA9RDLvGaJhfDdWpNePaX6hwa
JzOI1WXLmvjcfzIINmTABYbbEiUAlLGRo6KeYYQ0wlJidlZch8ow+Fr/YoFRylUlBAPglv+knicP
no2eXuHEEZzdr1+6BgseSWf4kg9FHM7m8XH+LAprnc+tS01w2duZXzV0FXG80ujc/pt0/jxYnCwz
FUSz3px6j+ii7WIbK2mtIfUP1JzXXvImdlQVRxMmnLsZvo7uOIyj0EhDS+hyHuSCjLFb26DjXxGp
qYlp7BQuxP78HidAmvYIiC5L10G6DtGpOh1v9V5K5ttyGBnBxzuKxXwfdDs+SBS4DYJjKlNzctRp
zLzMdCeXMHcaJWr9uFgbOde+yzQIuEQCZ8OgQyibM642odJJcVRYo+LdiSjLcs3mb42WW4dROtYj
SbT1dZ3Z3R+ZWjFup9l1dWQfWypGqdlos3CT4FMGp+G+OYh6MgxchFJ10lxCvOoUuQyuxVtVsmGo
78BMsR/5uS6eCL4MLxvExDsXSU1Nywa4hqCj9if4LGmnxZHFUOGgvXsswUv7ot7DBSBx2IB37p3B
2mT3IOkbSWjsJGukpl+Nl1oyccka2k82Wi76j3szFUIptwDAS+BWFOXNv96i6BQYDCmxK2h6L5XB
8it7ywgb2fdA6otF6r5ErN7Kd4GcpYhJJK+fMcj80EU7qUlClY+WxVa9byZuRqTgDM+ySDcNhPWv
MN5Ba2TtwzYHa0v8XnGm3QDyfZjs1B26u3s+TxbrGUQHAjZhMzP/Z2r+Cd8yCZFq5EV+aigBoOMK
1bY4Kz2yG5uIHQhrLuxEb7TxoSciS2rCl3Vu3PGPYvW3MvcFiVca4oj2R+TBqAbBnsYUFdrlLWHX
XQmOuJ7jpSKLEQbp22pg28fri7T8Cwqn5QZlsq01rXz7GPGdALeqiLEEiwBOy9CM8QjnQM9cHpwC
9VHS/fns0h/vDCkgZr20e5YFVFNr1gghs2IqQyZeLLma34137c/lsFWhTC8UVdbBO3qIYh5cBC7w
u/8+pjEqLLUS7muUBeGZm0Xy4sIMQS7B/+om4cz03JIYbhk9pczaf6gcYNciqwxQAcTIrYEQBDPb
TBfx6ZA9Ub/ZPlQFyACS1uCBH4qEmQUEVGimHpiFCZhLJJ1tTaJwfNq2fjCc7IzfgOPyGY1fgxPW
4v9mr5Z1bW5RKYwZIEbMycx4C1Oapa9x06JLDkeiqLmC8KGRUUDFVy6176QszKObfCG+Zl8q0jzg
kpFo9N1myoWYY4iDJ1oE0pcXBWtRStVArg0lq4oCnKKdh2RSiH1QlDwJSqKRHdO9NrAexhsDYf/I
TcdRQmwE6/LHJ7yDS1SQLoD1L+IxwkooFaVXMYKz4c1mVGiU4116saNo15ZVMwtovlp4IbI6h15j
Fh5L6v3oRQ0RU0G+sysZX2j8VfUlDf6LpZ6WbFPiOR/5QsCeqePDiesOT90gyi3NYUuUblc092Tc
H34HDVd48y0e6O4Q6Pfh48qyTzFami2vKl+227/hGtPH34/mV/lJNv14tN7x3Fx8acavTTiNvM7d
sGnb/XlW/qlukRgHqTHU/Q24by4uWMNl83FqWDVP3bClAAk6ocFwzf64Nhy+wsnb71kEErCfgEEX
cfWYKBVuEizPWwb4lmFvBMpw/mg+l3QH1EgJgi5aUUWMwuUBmzLt0+GZk05vhoVqdvCZVIt52RA7
iVm+pgEJ//Uxy6R49nl2XEO946gAtpDogyORa0eCtqQmHMqbWyPDWwBTynU4spYTA9mVXbA6MO49
QbBY+xyQ9XOrlSeGf+u61Rr3HJb9fgpFa8gyuK+B+xCYrY9KhyEAN08Gl+JYFTqoAuf3VhurIQz7
P9pLnyNjgg5BLebnKZAAB79p0e0x39/1w37pltnvqPmJn8MlTSb8Djmsi2oCa1Bz+JDt2iJG4ZsN
3cxdgLk9Q5T/qyJLlRYZP/aTvUA7DLzEbkwIjh1sYXzaD0fc5qgXADtLAsu+1AF3PP8Tuz3HFRk2
wY50GmnxQf40wkDEX+FMJYgEH4vvjvSjumh//yfzqmyMhNhCIPl5+//JqPoiJ9T6NSAIKEDkUbp/
/0qw82nyoFjVFvmvuc5RPC2H8ySqJ8/uA4kEQo/2JrjmDY9idJYgk17N2dVHkCAUFmu3Q/x7TOeG
MCPlfqFndsJGj1xPnaXYKp95vNf2/ryDb0CLFv46EpyMnoErxzx+c3U0g6uGH4x1fYeXxdupyJVy
Z85bxCr+tuy6Ww4NqNmgCyfozBy6E0jpEc8NpQStiFdPGkFVGzG/LGzs6YIUl/pcDJCllndsXCnW
DtuyhrH5n/iZHnYg3RYm9DizkfRwvU8G+WHFWFYg4s9R6P+S27cS8VGhjGHF5QcS7DgirrLQ43ve
o1bSK/D/J29NIFvyHb34+eqY0EvT3gOJhmbER7w65b6FYsfHTrovy9eeGYm/6580xklwmYFpN+k3
pVUjDwBLhNRduHvjc9Pqih0Ulg3pKy3lqyZdnMyeHLxocXzgBbihEIXXWij/GXz/YbbdwwjELBN6
i1iBZQnNBiWHZMLPAtwVtGammVbv4L5A01l52Xrt0oZXVqXQjyAOON4+J994ddZ6QrenA8XUMiZ6
/9s5CIfaFXuIeWvhDJCqDO8cQoZATKBvVvm4YcWXPkyidtJZkXEgxDs7uS12XNcowUIiy2hdqJ0X
8eM5I9QzT1BJ2Qa7QLTmhmNMhs//ad60QUv83rSsEMh42cZVOQ/OeUYl1LrSMCwvFK+Wblqy9pZQ
ln77s+6qcVkqwRta3nHbFR3Aw8ChiRyVM7gVlNTucniu2HhMWSkzePtgaww4jGvR9CkI1oytRYnA
kpjRhywNeCriu7+vDDmVpP/2kdGoylGu95VNd1WLoQdaQCCe2e5se8JwdfgiKbABMJi5uvr793jK
q+E+2bzfDwylKn8Coqqryn/t01l1BGb0PtUaPaQNvFuLWWBy0gkFugiv4K9kqwDodeMhMPsDlb4S
bR45debXUvwcJZBQHR4PSHJ1z7Udvnr1u+S4QXTpoENXi6sanHnVeHLCiiKsaPRN+4Wb2upJSUl9
Dpwx0vdDsvqKE+Fj+DhyVTPg/+XL6xbZwGxAOI8dl/WQ18zemzyk/eNOZzEmFQpiIfYyMmuSmHRP
yVpGZ5jeZNCz13wRjtbeAk9aShgkgcSWUhhLOBe2RNGV1Ze7n2FB5mlyGjawdss03a8LZKU0vkhD
jb7KvvzoASp7Mn0gcD3VvUhi3kYujRrxtviDbxXg/pLKm8eSKDhEOvkNICPmpP97UrKwfqvpABYV
qE7nJXwPUpj4LzB/9rFgS4YxxHE1ZUqTmzxMEoFDA1G5+7udkAV2uIMi2D/Flunn7AGB/7VkIKkN
t0HvC1kXsdZChSF7vTis/wpEeji/A7E7AV7CP/qvgsai3o0gUJ0T50C09A2U9v2xIxAzjcCFBNlN
ZmhrE8EDlwk2UwDMTTfw2R+AmoxZ6d9xpd4RJCpOmEJs+NCBvk2elAxP92MSLyxr+D2iIsUCrrMF
Vj+d+eXQPCDQ13yJhwmUpev4hpeIfchvCI4o2F3BcpLbElz/6wurHJP4wQokFKBXUVMv0tvsvW+8
LfB4bY07rxrqPWXy1pNBNlDvdjnYhQQaGjd9s6RZr3YrbogXC9lK8S0pXCdzgtAV8aWI7Z/bfvdB
8/99rNmuL5oCmaHMOG52eo0QwF/htwgweic9G6A/jTe++H20J0P1Ky4D066f6EwcPJvbOUdmA1cI
FU6FxjXpIZCbTmq9caPO0bEuFiGcV2QBiZqoY5VLWccLGbgXiKrjGSnyYnRYEcZ60HNJSEQvX0JX
v7R2lk5/VdGL5C0HckjB0yIAeRIoy4sdJHtR2P3pJspyWQK+MqAfI0rRNZfjC/+T1R5GpLDF1nfH
ZjKyk1hFZQOWESUVuIzNDlJu7xnDGa4xKwv14ZUECFr1wtj9R13VqSEct3C9r6qiQ7CEKkHOdYWy
ulfXlX2E+TmbEG2tbV3Kxy7bqU8B+mwWLPhYwcAShYfrS9CG+BbZolx3rvgwkhxp7oUFgz9i883h
5lQUuwx81Ti0BcVS16X5yaA9BJ4PevAdW8nguffSLMz/1vkaIOVzJbnlZYmBRh75LIBMTk5HEEyL
zrN3E486QnCanzEEwn2q13WPZGUs5xamD+TVglR6zNyY6f76s0MKNYk2Q6rhQhwQNRHj951eTZFi
l8Ajyd1R9RzSA/9oqKlylFDyQXxL/H2Jz6WhblhB/yrBT/BZqVj6Z1vlxfDP2LsWmxRHP0A5RTRk
9SlmmRx4f52jrUTJVFS957zOnGrqwQb3jag9XNCtwAoC6krdB1Ael2cuMgVUoUHA+87gmPnqZoUg
Y+tE0oqeyaL2/+r9CawlrMw5N4NXevW6QTzACNNxuDS4hrJVbCNWh3hzt0pFmf98n2wN4j9mSJ7y
lHIRwhyp0LesjDAM8F1vw6X55DsYJY+DcHGsnunyw5fYio1WjZ0YDmuxbBSwBqYFhmO7XgjR37UO
+pdl0SBYWmvnEg/PjX0mxZNR1/N71gaKtU821NGFJqDFuyk/s6geS6S4z6VU1/tcZxJqVcHGQHON
qDLagA9F5q/hFGb9eNTv2X1QoUM8V7vXqXKG+Yy9KO+d0jCOSqAkV8/r1hjseRMArbokjUkYDMdI
w33RIekLFtkcXLHeIjdCdBresScus/tIptDXKzM95/gjw9edG82hGtND7a3n4/tCxY+BdQSDb0h/
gVRGI/+q+CWyB15r5jxcacOs/I4p/RDUohbuvt4lSMEprgK7pWvQwB0U67cey8NJksOd51LZeua8
kKeEUVx25bK8dGgM9qx/KAa5guGH3cksLeTXxwYBOVqzHauDTe4mI6cJ7yMxctLDKEnlmi/KhZpm
3QmxLSRCNZVjquJPERGA6CtpjijIJ8kNnkvKjZ9b46xFZyMAaqKkcsHmdzmP53FBjC0wG2lAMPl0
5M46C1ljdBCdL3bTO+DHNNAeLMJwZdlMvbUkB9GHIk2XPmhzQRYF7KtfAXsYQkS/MLK+JEjdSmrN
5YKcS/Wrp0MYe4NcDyKNUowRkMdtkgTpDmqynR/U4eigifUuoiV6maZNeBl+oXwPQjhlldGjuj8c
9NTdYZgYut/vGS84IheeHvNG5bTir7oBQmMbeN4FYI09cprIpWI3NftYaIjtUHKEiQMDdPTKNDhm
z+bV9JxCd3n1inTV/nrMYFFLk+eAqMJQgyCaoEKkMZE/kXn+dDp7ssFhCwPLDRWnnJEeIUf565++
dg3+68T5ikngDWgWp5iPx/iuxS6gPyGLsdmYLjeiKiaaSLVKM8/oM+K63pMBWSh9HxvRifgdzDnG
s7l3/C2axte4hVLXOCNBIzrsuZKZyKg9rAc9yFoFn8VEct8x3ME3i70/8emmJTthZToKbemMfGY/
nzrIcAW8DK6LwvDaTfwH4//sd7t8jilED4qIr6Tuy0ehafHtulQKt8HNDRrcCfg21Tv0ToO7m2KF
L4g1FCb+gjitUFNqrSfTx6qIkhqR6YsK1R0K5CVpLiJkV/RRT9PQJWfrPH6gSoGwPFmq5jyBfkrG
CbIgT3AMi213rBVgQjG2ZHCTLZYxsIXGBV72bNmiv6gnXjD4rHZ4lBSGdbl+eI+ClO/L04nx/CaW
2BrtxMF7PDmqopDqYtOFDQGFWE3cvxYD37HFV0Q4TWlM0rjxe3ZNH0+wWtQFWgQBDaJBP6aCLOCI
mI+Ylnh8LFlh47OfDBLtSTQKfYimveSKejWeTwrZcX7WvbW3mEfWsgm2JoOLHp3i41+CP1cmHmp0
59IxE06mgdfh7P03XVEZw596ak9oS0AFJFjJX4ZtjyTbBLc4rIfDdYSH2fU8/GLPSYNBNaOoKDCA
dMemmHjw39qUeXHYPzYhz5v7mM4LJg8kMWuL9ZOHYCFmtgPNAQ3DxhN996Njuwj8ubb1GSChOZkT
blTzrwYtKDuVuk2pbJuiTavGxpY8fROOIVyIXnxgwQbK7svp105Po+CGEVNdnBj5lChuDcPO7dlH
g8nFQ6dQXV0NizTWrIPtsRjXVEPge4UinNvSRn9B2SBjw+sPZ2xGYOzdHfR35AXOkPxr6piLNGsV
uZvjB3cNd14dZ5SB7hnxQ4wsWuERv/HcEpuQ777T0Uw+lo1jJoQVa2+aJ+5ogV0IV7ezxiB1L90m
Dl5K48E2NZISLvgTycYqCz4Gj0h1OcR1MUVkaRu4FlbLMZ3/Jmf8Uf5qfiRoq5esNRjq59tAYzZ1
gh2nGJ2M+5/RjEsYyvNT6mIPnNTbgASDcmbyXuyI71pwugJlwaQXIfGT6r9sKT3MU4Kytzn2uhgX
UATsZZTbJpU1FJqxgNblUIKLX/jYihbPpGcUk1D3gsOE5+AEqiuNK1mjT2PZ+O92cYnd/riS7lHO
LQ0UJaKNvnPbubozjgZPbGPCo9zixTa7KkkiZudLXAMT+F8QpHN5Cuf1zJGp8ZKaIvL1u8cvjmoK
krjJCyA53mGGDzwICbiYVq9aDUJPrZ7AZn2gmvazRLJcljdap6+fuxTFe00oCbpyS8i7Dn72w1vl
ie0cX6+qsdoI654zplXVcK78QJrmPAxFbrySreqCPaEkUR13Zafk0wfJ6jnOzmzIDPWR2sJngJ4Z
6WdXk269GAUQXQSpiXZdXW4fq04lB/cTa8WIftJDc16R7vk6roevur9ynWvj8w4hDOrxFw9zGj0b
73sk21//3t06hMmyzRJfVgDD2D7bpQwiTTYH3FBYlvgjsczbgC3ou/j4ytgDhpYGf1n2UJ84/wHu
Qb66WT2rrP616pSFli1JBnyXQnrZ6MyCRB1DT8hEiKJfbuSyP8rg0uH1RXGRhIC8+Sr/FD8gUfKp
ASoFNdLyfTWwMgweNUDv6Qc0Oe6oc4tdvaNb+RkI+W8WpXt6RFA22fuAgytUnRsW989lUb7qbE8K
iUA+vzNNt27m8sXLTURZ0Kvw82AkLwL/rHJ9afDAClG5cAS6cLkrnlueBYxSDHBJG4D3BL2MFDBu
nIOOtJmoK+aMI3okTh1ffjQPNMyDORIU8/ktAI8v+KgOkwSryp4NzjBMkeeZH0psSTTsJOKyLcJJ
x7gOMKfXvPPL9i9pZcnAQtfLZEfM2VNWjIpp7QD7B22WrRjEWu01kgHE7GvFf/KaGReKBZCImdfc
NEw7tKzyjI0omHfpULBxFI1rLQ6QcDmfxwk45rc4f2ARED2DJU9vSW8ckKkC+egt/96nUFDZlD6y
qy8ijegm0+9JBJlYKRmhf7uGI+7j6KhO4cb0I8LOzalsOHdSdVI/o9/7ZjkAEzonLGd1rtE3P/dx
JF1ycXGcFw4mt4A/kWppDJBklsIaseEYWybmdNuRiNhGTuhk0ARBwrUkVK/TBLyFuBH28zbCEC2u
TkjHb9ZtBrgjp7VBD0FigD1CvnvONqhReEW5Js9twre4Th+3v4M7oU2K6aOZ4HVdeha01bkfssqi
vs7qCfAP266d3Ev8TrPNQQ3vO/d23qOnfEPtbvEbRdqtm1AgrVdocXWDLvH5gAODscn5L4JtP5lu
THDnaYXMhdyYSOcbJ8pICxFYvnh7qKot/wp/k9xasABc9A8lt4FR9dMYAt/0z3W15Bb1aQheDJTw
4OrYJ3nMm5MdF2KmFntK+nqnnZBnkFa0s+/oZ3XDkUQ8UAcIokAtdiaiBwMiTrw/HGrvi7zjjioN
SkKAP/+8Tjwhox+gZRlXFxNnxdYjtBv2nb0hdm2iebpYh2bhbFpn68NnLhgWJttkGZ6PLUJ7wY1q
g9Q3yEa64qQb2AfLLn8+0Yk6006c1TxBhf1z6W964FoQl1o2y58oAVEwxd4VQ25BO5QKZrtKO4cr
KPWhWqrxk4USJf6adS85dHtIRVXelVOGHgbT3SMVjwuzfnX8QLs158TQWPKKkDCRH6RigSPBZgIJ
a1/XmNbxE1ehQo6de9xwQ/lzOLHxvCxe8nIn+QYc7eqSzMmyQWMHxO0dR3xnR8xXAAkiyqjA82yr
hrylCtLHuxryu4spj06m189yMSI6r5a1kty4VhNa7uHTqOtmI4ywc4Psfwm0uj+Pxb78+fUiaxtX
pu9x74E+kEvnxf8GxjJdOsaqDvRTHrtYQoEIElj4ctxRo2kNkppTLWkvv3VQpaWGyO1b//puHIUe
r03c/sHGnOGOeG8ck9WAOpmYuFt4nvBixypM+Z/EHN34e3yvCkNFueEdvNbXf+ER5bdiGCkZC196
QrJPITeWvixW4xg2ukT4r6pBxfjKglswEnJyqZynIIEMwp7/9/3KWub3CgMQ84CpUX8IQ4LQoXql
qrgqawBC5glvTouu+7HNHDjrvidh1no1W1JnYwcQ+HOwmzav7nL5nlHbzWqbV+VzTazCzDOuo+d6
R3U97L+8EK4zTiyx9A+qi0ERW5YiMhNsLfr92meTg9NGfozMdYS0u1wzToKqt7rBkwgkDQM+5iQk
tsAqwCqjIkx1/PmIxDkO4TEdu5rRcH0J3KgQaGIED61hNVo81cOESMiNy3V1ZDU6tKbEEbCv9X9k
dph9S0XqY2uXeC+DHj53CefRlQk7aQHd9cf9j163FtnBs4QdnPLoQaGLOyiV+7NPAoMzDmTsE0hw
02rBaqU/ssLVWZZKXe1cRcB4YhUsCYVLA4zQ6AHkiJchq1sluhEshO4+0ciJVUM4dNUTGB0rVwHa
HaxQeBM8yQcCaoE3UOVgsHUOYNy5I2FYm6EQjes3nXrcepf9Qdz0jNZDZfyshyYWRsdLclwoll/n
95xUcRSgAkwuTRVcmq4/4JOHwrzOLywC7fxHX2eaU28+UE1ZM7KG0LcjzqTb6XWfKEPGMe02+Bp8
6WY/bF+mbcjirO/se57lGFmGgkM1na7vuLvMjxJdjvcXRbWAcRiequPy/zbpOhpOLzab2NcGGpAD
JFOJ6DTITCogMg84zYYZAIpQJ/d3vw7LlzbiKzDQNXOQDSQygjK0BzrIx6bSCPLrsD6XnQCflJZa
6gaOlbP/fh1OnCY3dcNA4npAVhGgweqEKlfPS3ndsDKEcbRx+forrwJmS/0YgaowpFU3QM1dHegk
r3zB+mURneOTWrOARQmNT+xIeW3RR5eFLCAvHLueMgM44dAX5GmipzwANyS1Nlp/I73pXOgmHVm9
BVr/hoPNyAKb+aeEXeGzgkH8I++K4c0bODRcqqu2yrSBjWxxEh8IlmRSiP6y9km0BsuaGvxWD3pQ
mzAbBTXjUotUtR9FOcePy20PaP6Jg7Jupb+gROza3O/Mb7Dgux+Skkq8njxevXO3MFLcfi3C1sEY
V1vy+6UlmHpHM3IzPWeW2jID3N9+XQc29ms9J2bxrt9/FFMdkWhg+Hk4ScBKicOMCr66MCSJQdLI
EFgXUDreHvzpyz0vUH25Vllrk5TyRwslFidgD03h0OrGOccJeJ+2Nk8shV6NcgS2hWaJWI0RcwMj
hdw2cwLztdswiMoZH7Les5jW9utBauz2OsvPODkVKETqc4Wuj9ju2wj9fZi7DamRadKU3erdO3Et
PN3rWOwr9Eb/jWAEofudWZEygHPFcmYN+52b+AHTz1M9Fe7aQDS6ZqnAUEJ0CKtBD3Cu8FfEk2+t
COFi9pag+gXconXveDTlzb9mhZKpoVf7DgI43NWrkiRHOWPM1Rm2CJCOfasXHNHYW+GsCMECHExp
7lEbBX9RBc/Ufv5xUfZI0KD2l6DUjvYt4reim+Ykke/ucJV/vdpW+BjRO7LZlwqjdjw610KW+YwD
Qvy3xkF7fO2zlzaYS1G8qrxVVtXZ20kZKXd83fhk6fd0PnkZCocbJkf0UrBUkR3/APDdwTiEFO6P
ijaQBdcqLi8neHU5VzN3sKi3gVo72SeT0WEVaul4/X4ewd8V16vc3Z35Wu1kw0Q6mfm0KfYga1wp
c2hHIKE7jCcUC4NZ/n/l1o/7pkwZN/Ah8XXfJQjs6RPXPmxLCG0Rk4nker0n3hYJIq9pksGSRkhI
A2GXDuIBujEvwtxlUgY9LMOX/qDCSrZ4ObHGvuoLk/x030DKXk415bURnpPfUfA/WJwBtgsqzGGl
+YrtSXD/VqrZ1kDkEGPuwidHwr4W6ASvxg/VxOxD9S7hjTSEeZGaDTKQ8Tj6/IGbsn6cOGidOmbz
5EECbEArMUEAC5zyZqIXqNVL/zxXdFJL8glm7E+uUaUn3wuYoah57Ou6czdQaopd8gTCU1BWsT23
Xj7XIfEaAdAxPKcQLvUDkbFnHTqWf76FegyOfXq4WCU+AkZH3/FbMVN4Bvv6/D73RyxSlkZfBrzz
h2LS+3cBFmwZPqAmo4t2/vweNN5FV2iBDfotO/ZOmTAok1iEuTKCB7wIqcG5XpSDrIDemLmtGqnq
731HnrX3efu5RdYihEO8tPTi8oc7a675KDiNjmVj4mGqijsEGwmgFFshG2LaJkyM8BSuyNcPD7gF
/UHEhGfnia4BYR2qmnIw6010ZFRto2mZotuVh/QPBj1CVuVX1ehWYw49LfquDRC39alL4Fr4JE0c
eXE1yqUiLo8JW3jTJuFXEWa8MTtsnXcQe+9chTmWVk/2K92W3Pjzq2m+tXXoTctQuETDsKmGkN3x
+JjomTl2+Sge66cLURjKcZWwB8gUrs4LY9jmVJpI2nk5hjXFE3WN+5Dp6m3aTw4FvbuXMOvWLXy+
6v7yK7+SxtwaGaFCpIOaycIVQVrETN72PwzEXdgsMhTO2BPsWEjC4XzngswrDXcr8Kzmodst7IhJ
CUjqpkbcNI5BZJfoPYJx1aDTBMV5JBwVc5zDD1LcG6Bq1byuGNIrQs0AD3Lh7nlbTawD/S6dyvsb
TBl3JDamd24XuRgXijMwLTC10wlxhY4xTuWIrEQ3966Unf6IIKHLQZxRr7iazMRcBK3Dum3MLont
xBk74G5kb6dezPsLoZ+yh8ePmddU16QOGp8dFEkdqjsK4Ll+g0+yHzxX6XUrWwg2wOQ6RC9Xv4Y5
PWxUMghk7m/mfrZ3xYKEwQf5zcnu9XddymwPs8VNxYPw6zlMhlbOsqx7HszMtb4sMqV1Fdhj/8Hk
ylrb4b0Nj3gvsoJV28z4RZ8e0b5vGt/OqpTtDusRPI3QdnAVCVswIEHMvnpzaxYa8gPbDXH1Ukdr
CgAfAf01Yn4jVrpKo0+bsVnmHuypa/5RLuYiyru4I23xU/wBJ+ssjjsq+yJNAuKU04b7Xsct6TTm
Wg1OKIy8nhSLxRe1xez2uJHwUFFRaiWOPlcGdLFEgdiMiwsTXBfEWg2JUzB2bgWKaTtzkXXsMM+x
ivbGdKSf9Py0XmWEBduD5foCz+troC/0pdSpxDpNyml5DjvDR1KoQZdflZRP26QzyWgg8PRegosi
w34Wss8P/MIhykV/UZzNSnChyBLHr86mBJtfn1FyUfSWgEbM3kV/ji4Bv1uKVYQZKw/7B0wgStYA
so+UJ9zlyqMpPKiofQyReWpLTOE1/uTEwTETi2q64sgXfUVxK/2VQZSFzw8gPXH6ZqYWxsOMw04C
UNd3XYPJuEwVZZuiAlmUDrbN/UeGEBvZJpjEmB+xnNGOl3k7TtssTiPqRYOQraI4tKH0+SDbvmds
5c2lyc5hjtYWheqwp+K11cwnc5v4Mefqg6dwS5gXwmD2SekJ2c3RqVRkfnNEF18GDMcOZOCIVHNd
NIynNo3H/zfjgVs0XpvnkK/pNjceHZoFo34MBrx/zbEqXommX4U47vuSOmBIj1PX44wxbhyNMcTt
B7QOHJt9ukBU7qfVafd6OYQZbA62d0MEmQEMhwb3Q+OQLSiUvEeZzEJ67cafMs37FOsi6CmR5YXR
1aCpBqyZeiRgo8hYRcMihqx99podpG8PeszOoVfxsyR7QItOV4ptAxf4p3VLvJ6PxtP26K7lidbP
z2bJrE75MpnI9P11bzD99NWv9/Zap4krLLbNwh4TmJsAv09MaYh0T5LSo4XQU19iRUtYwUKaTaln
/spQVtCiCbkedy1gtSKh3Nxzf0nYZ57Rvk+fXbD60hzBVbpIr1s2g3xK2+fmwZ1l6PLH49P/lHY1
3HK5CvhU5EQjy7194AgwTZHf5YCdhJ3pCvEfWmuKb/kFcYeZRJ2jrMo/XT56OgapYfU4qe8uvqTI
fOvN95sTuzEzYFIn+JYHUsGkBMTztDE74NUyIH2rh30TYsivCo4O/hGdoODgnlxrt6R/O06SK5T2
EhTCpBdJAkfv3hKiDcLsQPJhamQP6edxgXMWEjK7W0+TqagOPZHQE2ABNhZ21q70BvnRWrFpmyRT
xCAAM1DxYZbKLRhA9YWnS99+0HeN8p5zi+5HIrFBOqizgvjUF+edARYj2YWb1/hhffnTGftqYNBN
qAJY0KYlEOvBMe9MuG3x0Eg16aB2NeQRf1DYC9p7U2jfOT5eP0L4DsHt04hWaO6XjPHWV3ahXusv
Sjx4l9phGANwvwEKXnbwzMjq2Tf5u+D/+amXJobxBqCQICLe1zC2FcX2scpjV8Qc4Dh0wmbq0ux6
2xtDq0YBwKOIzKwxE7wTHc09zGHzF3ph9AkGv+yLtZDQpasl7IODcvUpDsbhB1L0oMVzlSjSmde1
zovq9d8RXYrNLBMTjscZzpFsl0kEpmKYsEu8Qxm01jw39QTCvjVKnf4z+p5b+jg74D36flCwl5HG
DyR7Tn8/7zRyWRxDIdMraC1uQDfMRniHT+BtggRO9i7YMGRQwuhGCvZ1ZKpQ8HydfR0s2bOnWyFV
C0IT6qiyTA4D4r7V2AbTdudPtM+OB6GLlB8olgNd2+T7btvF68B1Xccmb+wWyRNeWh7meZZ+kYFz
iwHpQpRmGJ/lwQ+qszaqZ3dypPuBRoc90Nxm7GuiLm8cm6BMbLjZmqpWQQU/cmAHQHQ5woZa4c2r
BlcNqsUBLci/blVRdUiYkBL/RV/dDqtyBoGGw5B+UIlWoOLm3OsQxwDDmCqwIa+8cg1K/mHIOY9U
XwXpSRrxMh10Iyi/21EncC/uqBrx+38Dq4ywZfhsNi2fTOEg0FZ380Z+CUCacQtR3HmhObk66Z7M
7XNdLa3x1rRm7chHPxsM752sa6/yHuZnqY96MnO0+TFGcLClpxiy95aSfWIKmaOBYtWZeSrQh2t8
ofiNwCU0Xf8AdxQdy2cYlYdVF14GLeWGjv8Wnt3MnFcWuF+wMLNn0bWDaI+cx3Azn/Ntd/Z2sVL3
cQR02kyOOroxOXM+s3Yo8TO+Ht3HZcfZhIlmOvGr1GT9iikZjzFfjsJUMJW6ll6AQBJqLuzidoO/
eaOQHHUuXehr47LlHo6yboGVp8WKrytMQdTvCOI9WMbuWn5VecmGaggD/jQMtg1xmUWqdILCA2Ra
aKW4oWw+gbx3zroEexIXxMvEWq1dnTMXW6EsrYrGbs6Eo35cIBSYzykXJ0HMsKQTC65benCS0Ny0
M0Egrh4Q3UGBqztrVp6vkmkGv9P4K1Jqgstd31Ev45NDO29IbrfjSh/cQQb+cNpmladdoxNYxFIt
705q0QypUoNZnY6lSMX80sav5CLmSNFsB4sbMFjY7Ld3ydtHORizoQybhxow5y4o0tyXhnIr5wWt
ljbp9K86/lX4AYjcUMm+MpFvtzIx5wzIOwIZwqFh/D5IqvJZgjeQxtVTemUifbK5DumeZnMcQqE5
/JwhQe/K4/EGJTaAAWdpHIHk2qRnsIM7gDd7INxs6Z/bpVxmWPkbsW+hTv2cU3tb80nf5/ZMqbkl
8VgPtaJhmBOek0sUdXBMqKLDWSEhPQC0d7Pds+7StdUF17JAh3VnYczZyDVbAtIqg34/GVicQi1y
ht5NWHTObZ9p0Ggx3cyR66B8CooHunTVno9mC1CoOtKcQgVaQ0ToxfNiT03wDEwCG3VW4q25p/cS
qMDF0N16nNzToYfRisAqlQaqQ62vkUEzOT7NqxW7nWoTHuE3oHawPeQ/M5ysKVjk2GUVjvb2CfER
ZfYqS2+pzGLaMX+flXs8v8wAGPmDnvRrOHukdG+QSNCQTbAS3F3O0vrJFt3YL06JWloCmWfWaSFb
A32C12RdnUrk7VDUWPtW+e1BYZzHqsBmiSW5TUxBAxPYn2H33A8ZZ0PZFmpTzQfVe6KqTmmuuU+L
t+6tF7AdxPvarZ2F6q0JbnYr98RKAZ+l9AAHOROKzRpkgbe1qNMtgsHijzdPbgQLLTsQXOBXRWwF
00HIYagv9hkdsbQbrAwwXFkLQGt1o0+WHKhd6KZG6qazD26s0MAenBJDXTt5H77ZFVw8060Aa8KJ
g7SZFJLo2+QiRMSIx9h/lLvc4xinUnbLSlo13tinHzcPbtYuKsNWrkmvdv5qHcvJ5Q/+4sllc6F0
y5rCPMpCxm7IO/X68uebfeUku+mOXSx00aXG/1ScmRFm40OAbf4W7YX++7rX0pb+/TtzoiH6J1Py
u6peNFx9V/zJoni9sCETxnt8Q2qoUuDZKUyrdFXznB6t1NNQ4D3E05c6QaIQoJHobfHp7immR5AH
rG7ZCII2eD3awnMVOhmCQvTWdCTODC9YgavjZylWY1CtGEyh0jtGG9Ya6/T++keFQ/Gysnkb5ekZ
8tyPRF3ey7LS+JBYCyjX9KWeAlWLpfRjM6UvmWLbhdAM9dLW6CUvRbDbSeHgfA2AmrCbDPSLGOrI
pnHcPho2kM00G5EDiA6gqO8TacQatmfVRBpNT+JWLpoJlKDeevet0leQdfY6+uuJX0g0Nm3dezXF
rkInYiw5V+uzPSZyKIwsb1bZJjWFptz0fZl7ebgS5dnAmDlWGSzSFyDyWqdx1bJEQyLpE3hLwxFz
4ZmBK2E7M5N1lUzYS74BhR81JH4jcx7A+y4P7B5UvcmVEkjgzCv2ExpNGW5nD4mXgFlyXI8kSn9D
JQrTrisbds2TX+xAvsbNsZf76tNikpfOb5YLcD9eEbo95jFnxgk6hux5jb1FzHVKF0+nTGfpqmjb
imqXNUBiQ3q6cY6UHHSqHdDuWr4P6P8yqjnjeLo1L2M0YETYIkmIEfdMCd6l62cULiFHDzCrLeuQ
Fh6AF/rgeuX9nlUUCkGJY/tgygDFJoDZ+19++vbYajDoeBUKPf3P5ilicbQzMvz7Ezui7HNNthv7
Etn6iIHgCVXVIjCyRVb71wUoIS4j/K17SquUNa+PUbMrRzxLCxAXlOz822kjye36Vgkt9NwtvNsj
2wiK33UzK6YQlkrIWpd+AqnqccJDxoIEkIJo9gxx4O2MGp04FwcLImvp66At07OA74ZVhZQTSQyw
PF30NFer3aTM26zCefZXxMcQ/MjeNHeMyiCu0zgq+JH2y/MmgYG4F54FbDeVIZydaN2wECt2R8Ri
Y2eVYmlz78SDN2noKUd8dPspf9cvlRPcwCp3sJ8pPtFNKx24rxIsv/uh8WeWfuoyHntSKDZT3aPC
OOZMpsv9+Or6V/NEZXnfbkevrtFOXK1vMm5f4cQVnxeJRl1/6R1h9SzLo7i82FhK8pCmIAIoe060
j8Z8NixaAa0q6qcBLUhNz7ZbcYp65EboQvnGPEB/Hf9hL1mwxtNx3t9g1Yx489hUA3A+nxzIRuHi
OVIVcbqbQCiGCvdnQcrpP5nztXnyL56fkcUNSGA0bC2jqnHJj2Y04Dqnm5p3Cp1D3QIaKbx1Yxjo
5Ocymz+TDvpZKCZ8H3LlAkHxSFONC1fB/WKL2k5ehzl6e6P2VSeYaykdcgg0mhL7NB92VrnWEa8q
FKrPO4TKIuttYqF1iIZcNvkhyhs768X4HnS+0sf1yEw/M/8zG2Fy1aG+5DQVTrK6aplBaOMSzUQ8
q33Ffq19FrLljagKmvYtAx25dMX2VO48mKPP7twBCAxxJuHJNHs7sagDbaOR/DRjz4dZKvTJxcCH
jE2QdlyRY+FvrlhFWm7yUZ1/U3jGKfaXsEhRbL3S/oEvyKAhBG+PRhrF/fCyWLYa+7V1z4eQOYGs
TQKtBLR7MlTVJSjwIHkWgXALOcbayKnwhyz98H4wA90AojCICLwAYa0p5WRJ3GqEupGvhJBHu/4s
MMGdQJ8KzU3kPDxb90S/hfnxp9C/HBJ52IrJ/pZICM/GSBHJgFfbrzNPNHMKXkdxea5QCcFG011b
ZGdFZAC8iUE8cXn2ygIIG1gVCkyCqOD9K+W/o+QCPXAX6oml1RZvyTLLu0CJqamNT8VG/ejXq7o8
dnRo30n/zjiNQ+CgnsYMcavXHRotmCbUPYA7TpCsJt3I72ZfNkqhG5JUrcTvQv//VpMsRaJVpThO
a/m9RBI5kozJo9PIuR9XLA+egDmBAwGLhYH/gnlYMQOLQKS1YpExNOpNXGdDVg7Tw9tMi2BfCm45
3QQLfB6MPXeCcKWXPA4crneZzqTYz2HGbnr6EpqrskBGIaJzjJlCDiO8rk5kiiHEP4BV+Oc7VmHy
7VRG6zpWsafR55jCCqgGKagX2FwExv+kqgNgSLcIOQHmCZK4PRwJAPvg73In956VIEp03WuvLkrv
EclEYBWe18eguKPy7r7WswZfIsZkEu2XBRvaVCmO+FmABeBf6Tr8VGl1IHTQUOvCAcsdQUFQNjfH
oULx9TKtftEPnJ4Xk97nGEGxmtdjUDdGd6IXX5yW7bfNY2APxUGDFeQGSNTlwfcwRAxjT+FiIyLa
OWNZQsWnPNs3mvp78NhIOmMV7ZMbFVp4kCis0C5BHZ6s7lhmoUE4jdvp/2fRSEo00rSaY0g+7UXi
W3TlRS+Ote2cKu7ZGxHBKj70ivoiIn1pQsKhKClXNsOAgGuI63De8Y4PndzoE5+i/QEL6U73w4pG
BmDyJa9I8aVbPmpRhKNsIvCHe8/Ui6Gr9aKdAMdDFg31qU0m8GCHoKWPlwtj1zuja9zZbAd6EPVb
9TABJsVWFM7GehvradCl51NBmgLpb/ebj5ykOR7cOyr06ZWDK5/LlPVHRYob9flYVe8HvSjR9CdV
q1OTb6urD5deCMwqAJ9OCjoJ7y6gpj8VZI046mjtP5+10OTd6EEWJVSpKdqYMgbjeMpNY7zIb9m9
FkMUfOdsVUvbISnxM1vtpCL44W/GpUfg2aa7oLLUr1ILUfZz4nWEHQGQMKMIQKpkeoYaXDJd2jxL
RiNWQESQb3doHJKcXggXBBxdOCPfaHKr5pIu/GHha1bSmGQ1KpiHrPF/KR/wzp/27tabbzzDQcBq
G+0p3SEYuxD68LFBSTVan5NUy7vhY5tqLDbNZKEX/BCFy2eVxWWgycs/90uW5+E9glRNPvS8G7xm
AaqU81thnCJYksPkMMLSxUETq194HcGOsi/Fu72XnM6XjlsaePNuyloHebHKqNvsEnMQC5AZY09w
o/ErqkspwPGcOqADi1FmgQRAuTb/AqTR7B5opxtbywS4zbutsQ3nQnudVCq75XbQou6W9B0q5jRJ
sagd0QUzliRqvNvXrkjlCrzOsMQ9sB+zOJGWARMog69F1RirqK+Kr67aMbc7E7EzZFt1aQr5C/5l
UYAP1Ac7+dE78uEAgg1V9ZeK49J9wGL0F9Ictn7bYcuZbWbiIZBmcFdNLS9K0WwYSTg3Jr0u0eVA
+fNJqe339mO4jPKpJ+0PgJDlyc9LBzkyvguOr5kWJ8597OMiQlrpcU03OyFRzUOkHBr6qcOkMxMj
KzZYrM2HoLGu3tbNQHMGynQcikv++Kf5YapsARf4NqZt2ctxnVXrUv93CssV9LQgb25m9o/Y/6y5
o4/MWbNasU5PQYKU6xVLwInKryEZb7AbnaCmb8y1ptvAD6zOrqj9OPuryabEHXMZcoXZ3aR/KlBl
u1eTr0jaf5dR01IPhJGkf+0vhM2P0BZ/H1XWNiepAhWAhF701URnonGtZJpK0S+go0nSLu0t3YWo
/7/HuaVHO8MmH/EpOH1AwmLJkCrqU+6O2L40zRq8nbnCH/SKGokDObyHJ72hza4CEoM0IIUBf8En
y1NjfTNtI3CGPrgJzt4ZOEqsj4REgqr4pyglQetk9dd6B9X6olvx1QZgfViw07FJv38xDQ+nPu1S
T+kyD7j2Bfn6lXxMyNPNxVk120cKQOTAXihGcPNC3RWMW93DuTApnX/4CXv6b7J22glSDcZHC6LJ
9O++AzD2kTXStpwCNoF2eMxjttJQRe5m4ZBHoo8nWVHZnlZN9MSw2DtzONV8tjE9fadzY7LSGiE8
UZ0njCBhPJ7YbI7uO1R4U9A5qJrFyJ99ilBp0Cwn6W6Bk8b0CKCKCUj8OkeP0DQEbKBzpvXLeJkJ
LKQ2w9pd0EaM5nX+hpy+Ls/zTVsj2NLWjlXTjPDX8T3MFqtqdCRl+Z+GTTSQMwaVivSIfzfUWjdd
OvHYvbuUJHgoTYYJjgSRTGHoZeh/6AsS/9YsRhqz6EmCoQRSRv7l1mzOfDBnz/nYx7taHyR5CUxq
W/aGS15wBcd9ouN7hAJH9be/A/qLRCy+MC8f6V7WtXsPvAwaGihwH1TF7AmFfKAMQkR/RukIJBZP
tQ/LWi3qMum22A7LYhP+ZyZ1/IOcTDW1QC3un5mr2VHrkSkgy+Oy5XmwUUdjTwkqsgUlOUpHCf6x
8rF5sCcXptr5MWKzalmmEkYHdbjQ/xppb59gKUIQo7tvL2xrmojxJwX6xF3gUi17tq6Ekppb9T4M
rYUQFLlkRxjegPMGUtwb4VjNpAlZ0F07EinP82MNN8fWcea0+OS2b9mBBGddmSpiMcQSjOSP5NCR
axFYmjQrdc/skcRPY17lSq17clt0A/iSoal7eapgxgpoZeAe3lsUyRjHKVm/5c/fUohsEq+K5TQc
8dz92gKnGd1cg2nO5toBFITm1LMf+yP692Z18Vq0Blc6H7qWSiP3YMIkDqxac55hQH2kaFfQsgK8
ogZ12h8wzirAFNO+5AOXTKKOhECEtLO/7VMQ9yPVzS8xnBD2sW1ZjXN5j3aRg9iWvzni4a2zP5Wr
6v27ZsFbltTkqpXa0+50Tncy8dZjshu1UNDcHGIeFwZlxcGtVeIuXYlK9FYJ3AlAs/doNXLl/B5D
xwb2nZEbFg/aXzNnObaQZ3sphsqUrHhKDkAjKi6n9PzD0BxrsH1Hn30MOe8l0bN9+Jjwdi1dAYuE
uJXskO5jgF8Plqe+wbhFcAqFpbms5SnLJugKTaHLUUyD5+iU0sXjmZuugV1zsAbZ/JVj1BXyjl0y
3BHzvba/dCQksLDE5pjeeZ2lSZD97GDJlHySNbl60nbXO5bCPu2nUFBWGAv/zVXA8EobhnmhHQsv
23WoT7Yo/K02D7p9Z3G1vEjsDcGOfsFlztjqjQ35y8HLY+/JOIGyX7nbTQKuIVLorgK8/hUi858p
NdN+QqI9ZjA13jDtRnyCEyLVvTjojgqXxMikquTn+4Q5UKDbT8mQyMTXN9SqA0dU2ZvjvC4I+Z6f
Hfx7iOKXopaqc0zBIxGKZOZU+c+TuWBhVOQJo8MRKlzbpBL2fnaBpzi561xqBizUlYCW8PgYfJoc
4UxrcjDlfxbPk+qUENcdw8SvQvDu8LV4AmkAvScvo34iMqKQKKLU+Te5gcJuHcoZg4MZFOyiWVLM
GL6yXpwbAXCQSyuJNUBpiL0yQrU9xT7bIqNr8c3Ndql+AdpbgCIhmPXz2MkghuwPcLk+Y2W8g1k7
riOB+JfJf3tTLhzrnC6CGXN0WZDKRROI2pQGC6Ci7GzNqh1QHYluWZzkpl6UXUIPYFDPFyUfk/sQ
qKzZmlqTrK2vbTYxrucOf9x+w247bB3fZTIyiA/LaCROQSAvqvNthcGV/wbLMbXPYy+FSiaT6IAw
8G/jBehgIohr7quDZCMIEVXMlBl5WSQlnZJBhi3H44L7+su+n0TAR/X48VQ4GU0591kCl7/lLYbX
7ge4VvI6DGyMLy5GEybUwKYLhwasO7KiNeiIG7QwaezztVSEz/q+qBUZF4UbA3JoovI49jUSF0t+
bZ760WmMbC41HvVG4EzexfwHldY6nW1LYoUXFMbjv2p17Fv0B2X5scsJuty91tgpT1uEIt7pKfEa
rg0nMa4gIr8wvxdU2n8aErFfb5jOkX6B5HqNdBlRvnyAbUHQZ5+i92b+Ed+jjHt+fkQ6LvQ9qCOW
wyrFXVtyrnf4qjBRR9+UxQ42ZuMBGS7OOvD/QLQJ1tIuCcwzxEmb1mz3xBS0tUaFcS+zgZDIuVBg
dFe2ohw7OJUTy+CzZnWYMw9W0oyYNu8Dbx8pHieY1hUq33IPFngTB7V0hLZ8VjeNC9en1Eiz7to7
j/RaM075y35JFjlMzd/dCNLEUOqgJGE8+bp9SZKzsf+Qp68ja33dGo1NozZoeQb0he8Q8lITLSqC
c2CFZ9ivI/dHLi6jtcBcIgvCyhlilY37reHvEbr8/hkfITcpibFxQC96JgTNe0QlSUCp0mAyHht3
p/v0wQ9HMF/PfhB/DCHp9jZDslVCLaw8fdQLqVi9PY3Vk7/wtI69rY8DnqVaoFU0z0YvSLV/ktS0
fVUs9ddm5N1x7he6NYf4tbpkDv1/i3L19fr2asW2rQSl6Hs3wxjtJSQsZcmy/H6KX9gYfFWs6LfC
QPKX517hEVawHzrs4Xg37ONqp0SetwTC5LHyAS/TMwrSu3VQFpvt3xNgQCdf68Vy+Dde4vIv1HM0
G0Xdamf5W8MVTPIXHXLNbGM/3xbkZ3iML5BPS0WK6SHmXV9BdF21B1XMXUIGrgdg4tGheOlMkrpi
fWxUxnCzjII0Tn3lXcu3Gfd1upOUYgilCQvgvR848zpANyLzbFXcYkNciaMOpv+7Yo5vLhn3+mdw
4ihAJQWxfHI/2IUa1RG5Y7OsTnK6oIqAfSJt6M345t1EQ7XVv+SnUQxCXtXLaMlGvg5JIx4jQqkZ
wHUyC3YAt6uhxjDAw4jGtvik2naLMlpp8N4wq1N5TBIE2VtA9dkoLSP8XbZ2rXPc5o1QH4cbNcTZ
ZQP0ZTpdc6pum5+21lekzT+aBY5+K7GvKPuNNczZPORWMdfXoBTyhP51YbjrufIXYRoUpJ66Naz2
7FKlfobRZUO26MTEh3IMQhW/uvadI7ycekDmEbe9I3TR6NZynI2GpjuZlmWfRZcY3h/kvJ8aPput
wZNFnXPp/pb5EPmibuEMaPtVniPH09PofXwZfnVx43Fm3ip88HndRRb1Y0WCdou3e68+HhFvXGWK
gCdFK54Hkai00E5Cr528Dz0R57V4Ip393cdxojmw2h2kejvh91jdelkojFdBryDx4ty0obDFxv8G
g3uxw8toUREza0ckYoGWHTXxqnBu0aVu1cspJOkuolNAnx0yDdw+Xjsm8KMuqCJTrkSNof2SjnvP
kqcFO12O5jCegiLq8xUM9kdHtp27WK+3ZRTkufGqQQj/N/KUjC4+wdHQ5lfCYd6L6ILaLCd9ST8I
gpuoC1USD8Xrcidq2rVh51mVkekQa6o27ckSX6WbjPpCb8cblGMVRo24A71N16KNnyC+12ZfTo4u
I9G8xKDccIxjCvTtvutnua0tbC9O2jjlnm1pawvq3CywZgGfTuPRBbb6h54PTzTk9RWb6uvQt541
9iNacOO2lR7QzlqBKt4oHZQ+maVc7NDK3LO6ZhKDCB8Ct7+3G9LJyg32IhTuO62t2RasAWc5V86M
lfEg3r5JIbIDablV49O4fEUOC0qc6+zpTOBkKNiPH/6XSEDDdw/NBUVxUWpN5vgS1mAik4DuSHJJ
rEAhf47cJXgWocbC8bxs5iiDyBTSwFl3ufY2Dj9Pw7jmgynJAwlJVVM4bMsvl8w51ZnWrTvq2k3p
IHGGv/Zr8CRvGE+cSSWyycXM59cg2jzCN0BBBZtAgZQewAkEmYXCXschHQRTqe5HaxM6XfTV2VX6
CY1edKpyQU1EA6HQZQuIn46BwBggl35R+BEGP1FbEPU9jVoOm++KX2uJYf5XIcyeztcVtd4vaXU8
zdTaaQfBKm9wqYau/ztHwoWwdHLn1OIUo3WvMIh+eUD4bp+vIfTkkJL8xadr53ZkqAGtbhF4yrWf
l+1UzEE28X2XvspGgvEbTaMhX6FD3LzELLLzgcQUv//YQoFZTdlUQdFDHLA80pc2KIZi76peCbvz
gjbwTCx7NTAG6waXlH46JzlvJ4OFJfy5Yle3/Wntbdre0Afsz2oNn4TRttKJdm8GvjxbaERjSqIL
9x00+HPoboRIVuRhQA8ReRULYX0pb9cv9AuS6/wblQfGBrhXpiZXySfe4bnE44iDrjiiPI9b5Fam
RQPfW7pVsovOYnuO4vEF2kkSSH/kjfVcSs5uhG8EX23iMJ7HyBX/DuoLHU96zCH44pDYxU25M45g
is5cwNeK6X2VmUazp4Jhk5GB1zWmQ2Zz/bEaD8gBxidnyXTC65jTSCVZKm2hFzyRkJF+HAX0i4On
ozdwZBv/LYL+nOrgVZ99MlXwHKSqRhWikBv6/BKWaWGvR9cyEstgX+EpJeEHzaftCMXh/bwfuAwJ
WwkiJcoW37xZTOSqPkY7xScPMgpMIzic802MWcfDbVEln5leErkY+4B4GHdGAwkdqtKV5sginuuF
1fomgNYff4ZccgrfzhwAoCnL20VEN925Mg7E/gpJhnvRAzRPMHwX87FfaA1cY+W1hqSCH564dNO7
4yKaQqN2eTEG31gBUnEeyDcpJje1ws/5MPyB3tUGoJydYGFNGj3jAnZdFTE2t2Fb0MBhv+a3XbbR
GnwrmfvyyHeAOugfPXhZ61NBBbfqGomZIdXM3yxW47fjEhRhjioYMxmY3Gr4xpmTeDVfyUYKJUeP
nJSJ9otbsvd3cKCd5K3l4l6xIfUylWqqBunfyxUZSYlcBhdOe3iBI6tC6mB05q3uhWOOtxrGO4dg
2h4L/zGeqsZL6f7RKjoHPzLlhJhPUfYLasNkg1c7KD54InaMDsiqBA4ZxvmtD/gXq8VFiz8xHqQn
j15hLMIKgqFZDQN9M4+h4mBkFCQUpC8ZUnB3aXgoXal3Sdgf+m5Z/VFIkIOTmBc3H3tJAYQW8x/V
zQEKro9E03u5cIiOza2bDO83HLz5wN7/6fqgU29WHAA5Vk4tkYa8J6kraABrEFHf8VSEYBF3Cqkc
0vCziYUrnQiIWDAYifGCZxkL9eMCpOKZdr1j7qNjdzFuv2RJb9dfwOwn49qlEtllWh1DoiCI5Bja
P1+oYMNfzI1/sx9pHxuuKmO5HTF9t/+eriGZvAJgnfpOT8fte/XYamdLPl8ItmIbCK75ViTCeKXr
2fwbe61dlgkzrsDbBkG2vseGk67Y6kI0WGZFlEHRwHOimr1DdkOK+cs5TdvBaaLL+wPE6YGssOgI
7CQJJXvL6EflNmqdgJSJ8ltebA+OMvNYoQ5NLLRQaVbdqDDcApOOMXPKT//W03bACsHKVdUokxVK
Vh3rE4EXlmyryZ/79tn1F0Y1X8e9+TpX+bnIm9Sw2AZuTEx7H4qnf9yOO9Ym3sy0jL6fZRZXr4ZD
MnE77mL0hL2fl2PXwo0R59X1ZV5OrorlvwJhAuVopx+zB+ulCqcRJKnc+9iCY8vv5Q5VcO3rjEO9
fDk1ET9FSSFbecXFdnEmMB2cndPnnHW/UFahcHE2hZpRuHW0r7jf5Tor0uvDiJURk2uHd/9HU0Lb
btg4NIP2AZ4kca0kBWpYOvuagGX6e7mozxYmx+aCcOJ39mCOPYcbkBJl+YzuLQLUSn+B8joDafbp
KMqQaCXIMb1O+o6PPmqD07XTDIMbf7ge54Ft9Zcp5l4xEJDxqQmwqCPIMVXItx8S4njSjakUIUIQ
e9lI7mlrDhPIoUUAgr6KQ5I8AXkI5/BErpw+jQP+weInlINP/HlVDG6NFSJXACWa7/VTdNZVFMRr
YNojDy4NUYAXbB3SR8Ulz6JnIPQrL8bO9CTrgGCvHFzViYAUdyt2fAO3creAChAwNy5CVoUCjCM9
tvsMcNRkFy3gf/F7MVyQ4ZaNV5tpPbVg2dZYyNP2VNDuSzzuNnxdvyGrY9cLBa9tJCOdrHCRW8xp
BU3yWmbKuumA8UgISzwX+yyk+DOqDWn9w7G9p8g1g/uvdfQL8KO4rGcMiaBCCWgiZqwVZoq8+hQm
gWWyn5zPKKhWzQb+RROvpXW8alTYN1+TKDbId0ylUyugvPT2V2JbFw58kcnElNE8HCeGsHY7ER1g
5/VZqei3Imb7J3dP+ySV39BOExQZyd+DA7DWimvkL7n/GBl7Qh/A+6FI36BAfW52XwJ9qzCzxBlz
WxW02UTWUICUGR18lGOMrLoUVTai3HEdisE3gyPNaXfmmyOR6x3VGr3qdTinmTx0D+ommfuykuta
ko440Lf+hVIhuHNIN83TaZoZJBXEOMvK+RFV2LbIYmoxt70hC/jejgyWfJvMOKwnYGorfcNeC6nc
OQ7SqNmmWJQM9JaiRtHrrkW2jZtVlJ/tNHzDvCPyUO1ZhzIUTyvjVWC/CBfvKfczc5uKb/T/bunL
snFQEHF4F59crwNnkbfZn23c2yoZJp8cKxN20fscriab3fURprDCIEyFJzN5g+kZym5coOncW317
9UAzb5amaQU5Gglhha1I7MHZwlw3p5cM5BAo4nD+qmGkAgas4jM/IVkbrBn51jojtHdnPxfP0INN
/1m27L5jCMbsV/oYV2TVKpiHpf/T3O/zcAp/Rt/507Bzb6HnwscQqkQ105SGd7DnOe74jb40WiNs
lF1Jp2dpbl+f5jnWMYXyFPgYCRHJA8c4ZcodOMwtMSlJJOd7RZFkVGZgYTSyEKIHBHTBZW+Jmh2o
lXJ1+wmC9+7/1nw+oeqJiNfQ9uL6VDVK5J5eQVKBQdiwLocffebOJfxZCPhCLeWHw/EuGrzYXwIZ
hZcn5SR6Zh12mis2bOiuveygEC3wFM3qzsmUl3rs/rmSMgofcpcyiQG7gmkSEInEgLaKU0f4wdkP
sL6jMNRkvh2WOOcjpd70pcT7lE1PeffI0PW4qLdQLksO7kKCmSWj2N/d63Ogfxb1tFR3/o2iflb9
OyJ29+kIwiM/92m5yGSs8OvcMRmB+uIxPmBt4buu+X9xSiMNsLQ6vmv2VSPiCTzaVlcak2NQKDol
ZoIP7tkT3G8PbQkhoqMgTSfCQo9vdwBdGZXu+CEJOfkuRTiRcBcawaCN/mTFOrGIL1jAI51XQEgO
6e3/FOnrKEMoR7VknV0rUW7lteuu1VIoAB9P7pO7y/vg7G45ghcnMg9Vsd6c14tOlUIpCuGKqT8N
RH51eu8R6vqCEQ2D6/m/h/mL8POngW7ol8embxvQgO6e85idMYgOLH1bL5zeQZhNQCLkqUaaU+B1
Ib4MUuuM4eFiPH3BrpPrVinuIomoA4j2Qq/Q6mkzrOeo3Htz6uYKPfVvg5tZU30FNcS++Y0bvCna
LwX9zBbU4c4LUgQYsJvHIYQm3rgNOy0F6178cgp7ou1YMmjAojA3tHBLHwUaKkg8B40m9T6cDh7+
cT0p41vGAaPjWKJDJz5FRq512zWR9H9dV3limRHz1Fk0XW0h4MlGM5ewLKthqnlYDGBOseIsDi6j
MxOr9YqF8j0Z7Ff18gzsuMMXMhPvuwe2UAnJ4RAD9uTa1wRdzKYeJ+7kmnojQvFP34q4DCJqDo6C
oVLIwR+Uy6boGY8FicW9iujUMGeOX1P6QP0wt1HwIr5V8giJ1F77DgPe53qUYq9HuroxlTVyrbWQ
GVxlegl1wGMYtlTwOLzVF7+6kI0LiIxlAlmL3vz6KmOV8NE4s0kbrho/8euL7Roi5j2BZtRfHe+i
TYBjWAZrmHnJApYi4ZTEa97Etcc480zPbgfqBOrlzoJ969pbva6lAlxbEivgmxDjghYMKI4B5zQC
Ibu0+Tn91yoXvL9ke1SfW6WJjBgflVWnxTnuiKMvHU441J3Cs4BmIhcvXqmBa7y6fiA8jKhszraU
aYOGo/Z+3m5oit9lHaAUUbA5K4fPqQV1SocWYo5JAEDnWk7Q0TZHiHDQGJq7aTO/8HAKPUFEJZD4
nYihS1hkUM0rYOGdQh/P/UxrSJg3JxP0VwZx8Gj4hoyNKEtEkQPs1rp+Ote1xSSmGYjoyrPdOVqp
s6qhctfKP63QmRk/46W2Xho13p+wlrcmaIfvgQEKiq/+A68433zZLY2JL9BwJZ8P+NUGNECgFtfy
6U6jeKWESEnkf2Kgo6JHg/T/yky1aqAmh+lqI5fDUSuqQ00AS9bIb80Uy6Q6iayhCBV77xN0auyR
sILSdlDs4ZlPcFVk/xLT36WGL3PpeMZjydFy/JRwTLyE7YgvzVLh14+91BIXvP+c6LvlYPDne3Tn
xN7pBpiVq/Cs8k1uBA7+JuumXD8tXvRbLi9QqW/oE1X8waLEH+68Lc50HOG6DcZ+3J8sFCw4IobL
bsy2MypARcx0zzURITS3iqzHzW4iqP+iAKaqD5U8vspVFgexu0YKbGjgvUZD+g8NqxJuI5dxPjIB
81bl4X1VDi/ZY8ytgZhLPPS+JrponMetGXP7Bp8dvxwl50D+hJN5bW1L/4KqnqwrmY/jQn/wXTtC
nNsRedkIoppYl3jbnBaml1HAJo6kAXZ5KSI36NtTnx6stxIoVsgIAq2QNIxop1dqH5xU/kKPsMsu
9niq3rUXyXajJdRWe2vVjrF1NobKyM/cDGKopyi0h6ocER2ycTfjdTdwuTbbvYeeEhTtgHPT0zUn
bqY+jL0WoAMUEdrt4m3uMRIdGSRdcCW4WRcApZOE+DQtxury1/u1UOxL1tOtcw+Qe2nOJpg2IQnH
Ql3YxVMVBfzPBu/WxRkpTFU+3m1NsHfV4JyGJ9MjszDzsK5jqokcFsjoK+tR6tRa2Y9rcbgO0rRN
FNbB5c3k835cUcAA8LjTtPlNxNcQdkDy1fBAaacrcg5TES0Y9GoXrG2UrXLuVLeuy0YZcpbDi/0c
w2jzro0EvcitYL8eiA2EfFJI61l+9LohT09TrbCGP0b6/9tns2Pj8Lf4mkEsaIAW7+uaSGowsp0U
4+nWg5BY1AG+o/8hzyFwdLGtDsqZMTGleBjuZGghtSoAq/kt3JS1J3KYRFmuGeOwGHs3vXx0EEnV
2iq7l9gGbuD3spR/iiieTTA25oaKcg+lVBI+ce5w0lEHarX9vKDiUMB3pTT9Z3dPc4sGvB61NfC0
1KX5kzdSpIxhCrTiC0Sr3/6Q4qJecHIZZ6btbmfYubUDBD8Md9kNpi8y6J8bnv6QXaJAUEh6O8qP
ksRAaohNFViNemig0sTZEIek/ClK26UKqLgWOP9N4NgRRrGBpUboB5/zTNgKGgY3sN6mwiOJjzv0
SBdsu6dnbtritXPO22tVCsy7Ub/a0Yeu12pR4fSdnWIthwL3wXSIg/G2m5TymcHP6gtgz0OqsnLd
UddIIpX5sPfUcUGX+a6tkuljHyQivpSbfNMp/5w87MoZVsb8hKqvIcYO4OMTVAGQNFKKA6u7RsQr
dMI7zD0eSoYauslyZ6ny7cVKYZ6Fn9ZOBSLCOxzyJrc7Wf0hMCiuFkVCCMzcKTUgfvBU9haXFyHP
dMUYMkxqaQf44Ej7QOe/SyyQNYB2dwtQz/UumgqoHHDqcRtz3ybHPjZZvwjHpHdD/IeG9PaSa1Es
fIlexi92tNsPju44eaiTzdk8QZSgYWA6S4I7PMrL1LVylZt+pD3u07FigZrxc1iCcD4ci4rkIbsP
i+aoSBfqumm23cWnrxpE4MNaXxUCyfUshxdpo8Hnl6DR083VUgzDMqQBKZzYDeZNgl+ygP+HoPG2
bjOIXVY1iCZBGhXpWjXFqop+i+xWRWR3bFvC+VRhJC1oGbctmloGf9bt6rAb+FpF6bEKgknSpMUk
BZYNXApv0X8mikICuVGmorF5f77mKcQsc15RMfK7HZRcKqjhhgztZNHZDv8OmXX8JlhGcr5inqTP
QPbZ0vpIH3jqpWZLzOUKXr9CI6eyeN16zKvRNmYYjDV6Astf3+IEfqDY2csMoTEu9QdAGamxyWAM
hTth8KOqZ3VwtvcwyoRfRmlhyCHwN3IqHxxijZMi3O1X14L88RqDejSEHF0SJf2IkngN0pO6dvH1
OumoKbVgGsIL1Q+0+PfCBbsIn7v+dDjqkEtGq0PtsjNOLVGJbCaO3Aw/Eyy1zvtA0n1E3RmYioKk
HQQURfn7iHT7l2rBOIhku9BJpDsurE7HVvQHupOeIcGJWfB6AV10flA9QWVPj9GsMFcffG6PeVRH
7FK53QwKDWnIBeDR6oLJUfwGirGVVofjj055iZQjLqqRXSSiClqapYcmEwFzIoq7o/WbttpypCQs
E9B5gsmFCEs3GrqUAn6EhqdcdUW8xWFE12ZyNAkqva+vA2K6gGNzjdimUKD6psNrKjo0X5c/QbPF
rnuLzSE+iW4sy1wDo2PGrPWLiRsND9s0tPsVkVxJtavzy3xWAvVFUIhvAK2HyCNJUQgPA6PpN8n+
1Vd+MQEBiIFjdg11Bcfk4rJbMJJMR3zZNgZipNBACgK/CAAWUcic5+AqI3rZs5Xy+skiFNQX2ncw
PRcJsZVX0wnAaa/Vkq1mZSvrF9ngLvjiGg+mkV1b1SubrhVkrJpVFP/GjtZiAO8k8WilRUTWyNZx
XXxTmeRdG1tKMQOCLKJcBtBob8w2pOP3QXHzFzGFFGI0IGMsqFIgukcNmKqoWxTzWa7gft0OsJuX
ri81t24DSXvFOOTpYG9AmXzl+PDIEcnVcctiNFcjTy+2R9oaMDRnt8+iR7qNa088OcP/N0WBbkIc
5uNuwcZ/dftbznO80WS25gK1r7g9NW3BwRHyCzSDf37gQ81asvGj0AxULp9oIj10R3+AYPDU0Iuz
4RRUUkraBQ4/1e5mTvc7HKgvHnHBf8V3OlUK47h6wwOnGPPt2jBZQrqtljk0ofPQeSt3V+I2Pv38
BMxddAnM/qWj7M9ryreKuorRjUa/+2rpVV9SoGWrIKTjbQ93rkp4eeZIarK7pElCZxvR8DQKh3Ga
nBofFj5c1WT4fiLWXWyrfMkiNBCQ2DKsxk2dLEU9zeXB2BgrOXEwfXuS5JUJ66+IiEFxd+Cuyp32
+CsV5/7mKdU5aI6v9MaSHsCC+vfdpgM5SkqMFQSgIVjOjdajhO9U+SaVuMp2RJwlRt3/QHLwW2F3
ypqhr1niP8J9G9CNZE72jihGVNGNq0B5/HpOww3vio1uM33MjMhFJFmCoBQuypOlOnnMpzldFymD
kKq9kcxDu3Kb8pmDtN47GpqEMUPCs54Hhe2OxX/6q1r2gjjlq+1SFqKmdNpLEeiOn8M942icSvpB
aYBIopOEC9Lq8YWJA5evD68AUWQ8z4xdzKRQ2pSY3miVqLzEAN30c0VkGnmoJskrdCjjvUtr1TU5
2i/mq5bNdh5tbhKJFS/BjVhiZjK0vyE1P+MGaezVa7YGF4YcfviaClH2YtxZQscgESqZVT+5SKYU
4N42DZddR7AYBS7esFPF4mwJZKRR86K4pa86m8J5M+sQWgEeuZTu7BuZU/T9bqimOTuHlVD8rqC9
nFGh6V4mHTiDuvErYgZXKYN1UaSlBTYZhsggSwfIlJYBGjYZjnn1ni7nLJESr/l8Mu9u9pROip8D
0uEp1tW6Ak+Fda1PtTMuudYI81sJUMkK4jYMQFyaiVgW9loD66FGp7REtqh3f7i1LYyZ/1xyxEEY
kKJYRQ5xLyoZQRLNS9Ck8ooxpDyHimZNrzUyoO+P5I0hzfw9NIWwRlOzSg/XPSDpDQEQkkwpdiTQ
ibfNvzAj/gClNp9lw/3YMiSvxNpfb+KdbnCD9EEZXhnZSn0yiuvJvF7XlcJBRlP22UxuhKHeY+u8
dT0Yop0l1hYN8YKV8pg/RW4IBPzvn+pTclZis341i7j2c/pKFOG+67bta+D97G2UtYbrAvFUXoLc
+Et0zUkdygUqy8GR/nhxL7iBYsQnN7RSKWDTxv1bWzMXPSMZ3W0AwPb2K6pBtszM+GlrbFssc7Am
G+/O147MAhmz8etoxvvDwy9Csgbai+HIq2qDYpV/WFzpnGfPZd8lpUlmsV2ccV+IaOQ6Ap+z7VrN
U+U64Vkr6D8fUwuRIMHX5yOhuRDhjRox5vfLnPWyBtsZqNZZbKB3NiF2YXdppSKyKR3VcIa2cKK2
whtKJyl+TvHCH6hBG5c4g9IjVBWAJt0SOdnGk0AoIFaEZ1ptI8zf6xrtIx0KKYhfRgZAEjUzqAIi
D5MGcKeGDxIDSNaJwAgBuU+ub8ndMMP9SIwj7Duan3QGsGs2EEKHk23e811P9GVsumpv2x7Ibhd2
HyzaoTybcerPE7UiwIVd0ZhDSNGK0EcUTNXg+x5+orThbHd+vKj1toHn7VvC2/j+nVDoxOSo40fM
MGqzQGImu8HWnoSXoJbzwMCmXPkiSE94C1S1fbpqf3fDsJOjLuJ8u3AwXVWyvKn3aTmQK23aoZsI
2CdvmjreZvo3U/Lrx/SlU1bWTrdhMFm28206Ugekc1EgoeL5q2is8Je0shO8/75InT7T2OWBGBjs
JUxIpmkBCff+6ZJQ9vJUiLlTuSE1IfBKXI0uOF+icZ83zpWSj6IajPAWSrF1gsaJ1C62IVpbulVS
iXitrjew8UBG/K1RtZRM5SeOOl3O0bLVr69+PhP5enn74X0y3QsHht8b9fT8FFXF14grUUjSLJTN
wMZ0NS4iOYUkWY/LrCAXbW1fn9X30MnSJdZXMVog2deAoQeNrJd7W7vpOE1L4sZuUNwYfQabKVXx
oAibbLztgtunsBcI7QDU8HpBZ6jPjD0n3NklR1BvhsOE5VH5LtaxSckX8v30uOo5xUApTDKFLYTg
FnlEwDKmhXaV9ri2sorOYfQgPKYK3sA4dTHhSFNwyHhpc9xuVGRp5sts4XD0l06ZdT/qoabzj4tl
GiGe/rUb1A1x7xDn0z2JSIGq2BaMz2hhoQJ9pFACzyk8YeQhmGqHj2eQzqMHTBtSFIdn0286nERi
jaYzGnXnBsbB7/tzU42GOdEYqsWtymF66WsVMhFdXpKbX/s6hxuOPjku/IU0wvRd3iauhN/BnjtV
nBEV9Xt35Be/WhIQbVgvv7x0ciMkvy6p6Z7mf5RpbH3wMLK6Xtltcghtn4eP5VJV3vUOF8loJhnJ
jZNdoKbU/JcVeG/5If6fdMWq1uN0lBt7K9go6cUnuwU01a5oB0liM0C8m7hZ6lQHvs4x1uTruWsc
UUUwgIodFCwKajOOubTfsZLY7f5is1dV0xNbt5CsIVe1UJrHshu79NJfX2NzESWCsnNf9n/9e31M
mRrs37sD8pslPwuh5WUnfbiHn3vhD+SpttbwJr39Emt18g04/0v7byIlwJmZsRebJwENVMg9rGE3
NLFQ7iLE8GcNQxec6GW2idQCnjKLVA8XiuCYEKMdauA410phkVmgUeisjtmiXlrOTssNNlsJ5gGe
kQlvPVDBvKkgh/6HxSudjmczChym9tEsCju9rg8DAclIld4L1tNaECmSS82bhED+BYQ28v885hSr
PnY5DkEfIqENImFA/lOzIA7bNZ0X2Y5B91tO1YMFL0TSIQJPUzMrVYBSDOedCrBRTj06l24ptUdV
WFJg91/eNl6aoKX1OX+8hI9qqK1jvTul32kCT+hpssj+RyyZqGQEIKNp3jLZ9ueyx8OUbk6RMBFe
+eJCQz8eURx8So3PJG+KohEqFKEftDUVL+TG/CqC9SolMQGR5lDj9wp/ubc+5LivwIhlUqmw0iZj
laW3pwwlLIpDy5FL8pKXJeznVtTb6XdZ/2eL1c1raU0XUG9jvwhZtmzJ+Fow03hwAoVCAKil+P5u
XbGBk4BfV3LObVtVfR8NINbqZER4XGTDhSjvIRAvc4aEX0Oy/Auo26RD655H08L4hKLwW7B6lLtN
tXbRvJ3vd8lYtks5jeYVJeXjguAkcGudzSff6KEUeCU+9mGLsiMMH/KaAs+4BgDj4mSCzx/n6OU9
1oluVtIEkhN/4Onxi3irtJcCxctPDeDfgYmLyFocB386yPCmv+SySo4EtsR7SmBwQJ6tx2ULS2Ld
RZ9aJiIThMjOCPy4xVOGsMm04c272XTpP+JTEVwgzaD6VPZ5chwDVdGKG1dNTG6RsYQLh8vCmDin
xRabCKdQH91FeoAvAFih9BdqSEBgpjqJcRgxv/+ZhP2nXZ8qt51v/0mek51OiHfU7OMt37jfV/bG
nJz+G+wHud5A6A8tJ+IyK9Sg4QaHPmDZyZUuwbyLEopVGxFBwI2qHRujU7r4bB/OikdCjb/Q4iGv
L5GcWgQpzHiGY+6IOPDgF2C1wKIsVpEX5ZRPeluNyi3yyEXhXm7D1D4BEsfXJLzs//Tc2i+uTJ/S
MHkmGeXQKNvvyCAc6bXwPt9qzTLnX8t9+x52mY7UvwCmfLILAE0QAGaA4AblNNBh7s4dFcdcUD0X
hs3EnLEFu1pI/5WtaiX3x0t6676YeCsgHjMPk58AuwfdqMXNDq/PB0pz3esdmIg843Hb0li2EugM
NpV1EZdNuPcc4/ieFoPQbLjl7dLtj0+Yp4UHJA8gzqQo1Pz21oipg6Nbf7O6fgz0OHsnTRXES/QS
ob1suOgizx7c9uOUd3kHUtnd6qgHefTm3KjUtMqFDNJ5Pq3KhrxUsm9q2lsjxOgO6p93+5w1ij7t
U9TBfgCT0G3i721SYHwm6WT/fCRSLKPb7TKk6W/VcCbwWwkccHRvbkNDuwOg4LORTkKKj9Tt6D/z
L78Hwq9M9dG31rovHpqPKYB0owYcGME/IQFJ73MID94GxsSQFA/bV1r3NAdTbGJqugdhW5RhfOD1
ppzasAY7bulzmI8zWUF9QDa03jbYRP3aCPM8IzhR5f/mgpF3O/RMWK5FvSTXOWbfogOjKHJeR3M9
T6Cvko7uDrtAP4lHmvVywze9q7IjKzWNSH4CnN4rBU+TQ1Ijl9Tls+//+e/D//ve0cEOm9/Y5lnp
/MtCVqLkBlSlPD3a0lbnJoecUO9d0/0kQCWnS7aSRG88/5QWYPV0WDuqbqAeiz0GfDJcgWxo6I3/
xaiXJZZXofWgktAhlIpMzMbSQtg+mV4MGQeFJMwWeqT0koOWc+BNkJc/5NbdPBSjWJq0vbIT+Mb9
Z4mZGrN2WAcFakjNPoewXPTAbwBJtaMBR+6tvIslGSoRW4UqUyW+rwKqw8/8xYd4IwRHYH7a9Ooz
VX4jy/EDJ97d8cW3sb9aoG8HalXr2DC6tahrXqgaWUIBbiZ4+DMazd2CzR1QSg9Mb6ZUuySrGgDk
PUbV6UOb6iuftbcnyDGMXREOEbHUvTHSU8JjKmoj1qX7skl0D0trqiOtkZPwpSgXHxLEK7JxKvOe
GA2Xg15vv/cUvkm/62RE1eTHpBAUlaR/zbmmOu9nX0teSpo8zw1pLjACEzNDies232K4v0erG8to
1APjCa80bnZ8xkO4Wj70M42CFUYOXGjEIxxOHixG1UE9gIC8TCBVhWYR/ImI1Txx7OQnR4kAezjZ
bdirhY9SAqYleLUVQ6oMo2U+Y7hMDbgSWhkgnW2t2TdUdwJdI0RBPvDo8kKbQKU3LNGGhOc1uQ+a
QCuENk3cbB6TsNuIVsKvjJEh2V30sblTzp69rwRL5JpDBWGlNMSMI/dIokf/80pjk9Bf4Vpv0slz
58PrfMYhRJI5YmGe8wKKdQPJoBJKHkE+grsh7MKFcz9lhdMd4UIfBiTIH7v2tOBrKPEHTw83/ynb
EqsNCzv/XcPj+Mvqo+3wcv7DPjKMNUnyo/JT+/MRd5fRdYboGWqIIuhx7wXMfYdjAuibXCYeam3o
UaWNEwqtyqbwy8ohxg9B/KTLscsm9k5xm/g3A7FQyIYRUB1UuVLh3EsWj2fx20KHAa+VOSFOUvLd
Z5h1NNzsmmak4LA+GIpHOxH4mU1BJp+e9mAwMcnd9qvBo6Pg1y5I+jTowsnI1mVGuvmzFl0zdlMA
lkb5htIdC/FsMaOQ+cZmUfx/bVL9dB0TT3YnviJJLxjUZ7uhkACFALGr7+HPsB1WRneZ0SLj2BUK
Kci0JWpLU7KfBYjpUNiVdItgIbbKqsfZpgeDsuNMVQqXuigougDLjHIkP6XnyazNdqpG/9BfOWU3
St4DDZvOfayXxIBPIaKaI5CS7DV2/MiYa1be616Rj6OzdJEmSh7yNXBRBYIjJwdfXTQvz38drRSz
h2H9SArvfqMN0YyYviGHLY1WnwV7ujIODv4z5/sHj82+k4fzh/v065mWyWSlCKpbQcCUEKiGxJhh
7PFrWjvGodkGSPEg0ouZmVElYwQ4blT3NnCrbMaX5GhY/blao24wWby7jDs9KhNt/i1bkLz2PITP
tcSy7dYf5sfuRalsqtmtxPmoa4TO02boVU8rxFULPBoZlwes+3oK3aJc6R5nUGjV16ACa0fbT3K3
SN1hsGzYQs26cqUMJDTinlPjKAJmnJJQ6k3L0HoaoiY5drB0XnoIE2VVsA8J8h8ELpQO2bOQj3N5
PhyGE9yUE7okxtXt96oPcssrgqXeTvcXfPqZyvBa6k+0HR9++YKYSthyfD9BRQ3WhPDBYosXsKIE
BfHdHeI89i9+JZ1V3xuOjJt6ybNpNNTwLT/P9HIrCkewgrhvo9zQmzgTwQqYQLWDN7g7SyiMzdq6
8xDBL6Rm05Qmt2xKYBoskTikWJdygM6jDxQBZA9v/yUc84+mmb9M1Da/RiVRppL2Ieg6gNOYP9RF
e6mEbJD9xEycvvMuHesCgq1JIpQ0Qw4/7QJg2ZsoP12syXjf5Q8gaqw03EZDXoME/1IkV6uMY7fI
mPo3zTLoa+sEuceM8QfGfqdGTqMp92Q/kTKhTzf5OlDCb4JTtu/vlXslOxHDQGW7TsgzwpLFiBXS
KK6LoqAL1pBMC99nl9VHCvpNN8i8F9qUdBegI4sjrEGnd1Ap9lQUVwKc36JeV8XN2xl2nYzMbGCH
ucBAq/coKTO7q3VHJ7Amy9doBVmdCVlDwxHku/0kfrI4rfdqLn+475pPk1ufxAnA5JMgbHax5sL1
KSY2CIMtryBon5V9YtpFSEgWx7KkiHMGtRV6da3iDPaKW3v4ZNbElfT/unU0bRB31jSzKEFJrJUb
+xR5vJahTQfmNCI7m8UlkzO8VGHKoQfGtPelWePcGPxZ8VlO0zvg1chxTY4HaV1tvyGJ9dE9Nls9
ZGLbwz9NfxMNdNLYdLdm1PXeyhSZdVSmMn2/nirlMOi3Qy+13wMvK0oAu8SZM+l6erGehOx99THb
yxdnn/uhc5Z0CdRYpLnM6FnRtQ281wA02IrSzUvTbiwLzk5dnrpkIBkTRwIhcHb/qAAg8AiANf1U
avelw7/O+hYamwqnOcDWCKgRel7qwlidtbtrIotkMF+SjdFh++rxfe96slzsDxPRTxXpQZoAPQMF
FsOYtbvmpWDY8Rxd9Jm8m6SgIEgnf7qNkz2FvLiS0Za0QDpErfIhG4LPdbiw4Cse4GJFAAsbHjs4
6VgPIHlX7vEMrZTdefIhtzowHloeb03Czs2xcpJN1QaF/Vu3ld7XQkN1G7OdU35HBF7G16jYS/3j
vhcG+/THFrSD3ap+yR2khU8DSvOfn/qCiGgA77Jz2Qoq2e2Maj5hmhcFXwDfUP7rrmReHSxRV89h
vVyV9a0lDiBsrcSrMeSFUMbhAokSGpOY7Oy6IWDCPqeVXhcHVU2u9zWvJLcTEmLTYIDxIcLx+VZ1
/QIHzmSKxg80wRGMCPwcIcaVCI3lZHY0U8PkdJlFP/7jkok28XmnfxGSZzjs9YrCGvAWaWA6g3Eb
cu3HzmCDOttsGJvqTiGrJACur5fPjYYtg3bIp0ZQjWTgqok71kMHoVqi1jdc4zfaWKl+OvWjtgu2
QkIYyOvNCjdbY0R6XEoLHA2HYrdO/aY2r8b7OLdXG7pnN1/e577/DNAKq8sMxJmIrZsLIb8IwOZI
eIAhyjRXaddQRjMOHcXEv+MFYTo4oAJYYdD+XpOcOVDdkQa5Sd74r6Shw9PqURNXFEJhuMSV1/ai
gnukkv6iPOoi8inJ/DZAdaktvAnUguri8wdk3uvCL24+11i52iyuQeFnffj/r1lVLiF1O0VgesR6
9kSZIfGk9Jr3lUWsq3bkJyFg0XpJNXSdpwVeFdlkvfgCT7GGc2tup7Ig4SbFm7Isxt2nca40ZvBd
oSsuCSnjkmY/L8PvPoWqFYFzOCx4ypa7InEIwSHKAaGZOsIE8SnuiwgwVO+Ix1wLOMzoy0OYGBLx
7BbWXKQ0jGLgX86NBAI+PS0Oz2v1MMbHp33kkirCQID/EbLrKjd0oC8BgKLbMe4g3jvrGwTI9mJ7
teg+UU0skN4UYIWJWCQLUgPVTs32zkPHteJs6rHBX6J++Q7Fq+62oKHzD15ZGfOr2Je+b5B3DA+W
ss8758bVgXF9pl1R+8kD6ABWeKMr69Wa7IczFop8+4wjjMZ0+98LgUgxJ4b8OSnekgct1IoAFncz
ELmnTmPY2GvhK5uRdHDOCpUFlIMQ4qiCNeJZbqTYRvegX4Jg7Bvt6GhdeMoHkYRfRPwzF/kILvbl
kO+yRWCvtBLt8zhN8j2Q8aE/3qJVdAm5SVdhIZblCEbU7R5r6UveYzSmVHoozNDG4G58HK1SAlrw
bcRhv2n4+ZJn89GxmgY7qpkihTlQMgW28gtIQ/B4bXxRbef0n/ff40uX0errgJMd08r6NQMLOR4T
dGn8kLqwq3ys4gJ4f2B8Qv+h5h56rlW4XP0ad2AKBmsXvW+vRAtpkShD+Ve+dJRWazOvu/E3ClBc
Ys3yrCXKOLyq6iK8GAvvLU41VVGDUj1QXN3qSThK3Jz0n9ICHygN1cu2dJNnPT6q0+jUcoaJT6TK
cwJVcM6CC3xSr3cISppinH0wsItWcpcZm8I/Dtd/QJk+
`pragma protect end_protected

// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
O+O8vOKH9DFUyFL3t5YImMdgIdhydwL3/V7iLO4U0E4Eq9OLaewlVVoL0WIr8kis6kM5RlIkyYae
jdtJkdVch3u2lSJmmxbYBO7K7pwzGGZPXAkMQ30i4H3C/j54LXK3wXSWvCO1oCR/XFI2wCSY5eRl
O1Eh7QpVXFrVZ+AJFLaxX0sZHM+RWcSOA4DKiLfxgYaRLqNSqFPKqCRSJsyOLjonYr0tIZP8dJ/u
isG42KfKOEoeKa7Cys4vBx75vKuEtPMKNAXkaTovmbLI4MFVCfqdXnOF30GihWbfhDJ9iPW6fR+f
FCFiYTkEL/Q0qLh87affiX3rbA6f5Mg/TdY4SA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 9008)
j4OnVGCse79ZlB0YgMr9pDsf2r5q7bgFijUvuZ7e6EFp05hPdr8TvWKZwUYhquPiQBbWL9Fg4jcx
93uEYm6ecEPuALO1gXJ0ir2dtL5Y151Y7tRB7mEv7UaERa28ViKo8NdFoJUG5jB7WcMHebN8JZ4t
DDAyLjDLGD7wsZJK8BYgxPW64aTprIaS0/zoGFmdOuy0lOoYqpiru8LN7HPcC9ARf5+NJAtFCRp5
dh0Uix1HwrJRoinbSJjAKpGE015CmBTN1vD/PkPekSkrVsXBSqOI3iCBE0iLYgk7jwZHYZwXTwmk
U9TkOtZrKAoIjN+wRHHNafLZHSq6psXP5n2HGSAt0yKruqYPy99Xl4puGQKcF0EddAgiuTZqqbyO
G9h2UvHhUx/yIZP8QIET+qyzwc8N2gzcXfl2X8PDxTgPRcv0bvQn31dK9qzV7jHQFi/hqBOZv53+
P+XbkwzPlmoQkeFlmDiJB/maNn6RpfP0CMAhO1rSRQZWGChbKzH4pd+noeKbRytK/2/Y9sywm4dc
QR1rxnG5CwRB0kgGg1x3JAPmLsJVOMk0zo1ItJMIceXRRCsuo9MSw5kscE5OAGINyQQG3F43egus
yE3qqDDlSfCQQmF6LjUoLcvlsQ569Slavn8vq4X6CZjJ+nvcMZb/xPU0WR4OwT6G/jjbeOX17L7j
G3dP0lXMVDZXai0rSGVEfxYiHio1GxW/C0VOhQuL7iPWdTt8ugyZvniUA43gzhmP2iLJNydARLN4
UdMu7bl+Z6vnJkph8ic4cxM4K5aX76/XYXFwyQDY6Q3TyVSpl32q5AiZZyw7p9lOc2g1ohD8CvDq
fS7qIERiEfFugjDp+9nrtrlMsr3BVnS9g6uJQa+zhZNx9dmmJRUZSBMQm400ugNQLghUwJimO+VW
h45MbteCfzOnVxSRBbmj78nvxlbDwzJuMXZ+FPF1EkB3/q4FxMrW1F2//1JSp47tBKV9rcNmqzNg
gOu9S+zggKQR07AnsJLfE8AimwnslhiKBecKhKBKBZw8cZNeJnfg3GwEtQ81RvXYEgThpp3tTLJK
8IgM24Rmkv+HKAF4VeUjmExl6xoCxZ5ZjX3Mu9QvXTo3yPiFVRiVB89uYraysrUcg3Y9yBiRKbp1
6zzYfwDj/fQGkndWHDY7fOqugMaqc/w+tH0YYyNAi9RseutSNuW5Bpd6E2uY6BOSQUy4uoid6bgI
xiPx/uGq2vaZJ8wMt2gGyadWEftJrb0S6PnceBkW6QOlDEQH4tsReI4MKfA1MeFT/IrLM5YOb/Sd
Iv7DHqiZojC7+/7Fhr4IkYDZeloaLwYOT4musONL5SWHm6KSGA8s46Rd5Qx4GUgDR4mEMniXDOiU
419tU3OoKeh480epFAZNO4BA30uDkJeN4J0JEncbAe/wX7AxbTzwKl/nvGZkB1tPt5jNXa87rJOL
A5NtLIEMxUWh5Cz9ZHL6Fz4/shnA7OksITlkoZGopSQZ+CmjjPkWCX5tq1yDSxojxSzajNjTgN3g
zxazmWRt9qqBCYQdjaWotB++eDYWWqldi9l8gq3RUcZoyyYS3181c74kyigqOrtQmHJ5gjsu/bKH
qJ+hrda65ekGwdDJaxgPzJCSUu/XoP5wLRrcRZ5cpPc65nXPR5ZBZNl+NWl89Vvg8bF3OcWTyZvg
avzV90kLPuTXEWY9wXJ68zPalP+zTwwyQgJ80+M4Jv1H2yG570xUs94NisAJ5LR/BFq971uNfOf7
X73YItsWHPrb5DY59/NbslNyDuwFoGa6stOo+QDFQv3AbcuNONuMniM7QsdidEfWO5clRszSODHU
nf/RRuAmhEdVIOG06eqhKOZXcNKDlkK2a452luU2u1AMsz7DAX/p4rkUUV2taELeMPZMbJK+uSvV
A0LIFvwWK/io+iq4GEMK/NKMPb3fq9MGT+6SR0GxCW3o9fuHCLcWPIstFdLIVmB9cw8i10Z2YnYc
Mz/wbIo02idZP2CuIqobdNJOOCHZkuF5EaiPq+kx7veL9zE280gakHU0N0ofpcjbGoEI/Gx+j8Jy
njfRG+A39dFDkwwiV6pktx7ciHob8x1IMV/YHIHmsWsoB6uTbfFYyM4rzHEa90SxFcP3oHzmeCSK
Ou2306eLOrb1iCXQEt3WoObk6h0jWsJk87iTUAzo+LO5DTrlNjq/OpbLLjNhP+I78IbZ6DFNnsUB
emaPNbPpFH04S/wS0uxFJQZkO2ZC/XmySBzz/OwRSHtBVvyVj4MfKQ1D5u8AdaA4Dgi5s/VnObkw
QDUh9B4RLiqgnSpAA7RX8GNt9Ny8dSVrHc9sw+Pay4t2V3qf5LolgtUDBi9OWwJ3G6O6lhkHIBUs
YhRBb12d4wnHOg66kc3MTi8MvVgPR6yjq8LdemWZxQ7jDB8uzsWKgIUQDpBtiLax7nIGkeq9W+Yb
rqnMSGCdIcF6pNN/NMpx/4aPxUvwUm8XeJ86BQ+Qg0ht8t30ZzfGYEMFmVWbyV7umMbZLF73mB38
jR5EnDxhtKFANqzQ0frpmlKRdFlv0zj2rKtEICXj3fmCxEVVmg7HvSjngv4QjMNBdyK+NPQGokx4
C01yqFDWIjd4sXrDDewYDSJsZZv7UxQjdML3GVJ14pMrU8z7vf7qW7wWUNaktJapyIJ6SQMyiya2
yvVwylN2o9YPugPTiNr/gUCTZZUaKKeLSVSWmGLsvS7M8W3zYxIHbY73cd9cXRqRVfPEC+0sQrD5
HMfr/exYVDCglM69MLjYoEJ/RQd5dbCfCgUZoF5ntCyD0ERZwOCvP5bfILvkBy2zjDlVdLzqpteA
evYRwH3yqHFHSB45CX6QpgypOP7AfG3m8LG6may7+ResHkJDHlSBqCC2h+qAJp8RoG6ClWrBmop5
5rnl4J4gktWYbnDm2gv5CQp0wYT2YekHN8eQuU6JRXaSPQIr5SUrDlueSCyVsColDXT9bFYEh+fa
l0mKQjjeDOeRuQUfBwhwFqz2NEwA3onu2bOKgGuL8HxWgiQ6oMqn//i+ftHd9DlK5LUSPcYKDtMK
02y/re6krRSvEz9Lun5FS+YoP8hsVbOeJygWUV6YbzANCR37qY2+eTP0ppFk+lsG+TKPMHdTIwCm
81P53f330YCQ9mbi0Scmf7z5c0/8vcKJEc9RZawgKluP52Z9RYplk+D4bqJRpU353ItWEa3ea17/
WzVx41HxhoYjpiJAOFS5eV/4ZBpaBsSq/3wZeC5zNASak/UNeKAwDmEy8Q0fcfxgV0nNRJf5fSFB
98yDfPuTw3FctBagh+nR4R4NDGzTkhXU4e89dc3+H9q36tvnDYR7BzGBEny/WkOXPvFWDPuLlHwk
DeSjcYL0bRWe93J59qyjGD+wfM4oYdUH04RMcwzEg/Vm4v+RFVP63IB5h+22PstowY/Fyirh1Frx
7CLLx65Dh4ZbYcWs/nJbuybGtUvuLR/SwtV6bQBi3fSOdwA/YUCEUT6j7NeTHPUfXfJ/RtkpqMeg
zE/xyrnj3qja6qoQR8Gl4ZLu//uc/PGXndsNl/zIry9hRDzRST9LHnCiFyOc5tHf6Jnj+M1BkO9z
rNgCGQJPOoU7xUzLYEiomxuilerBsWzAh6Z1xgQiCnRrZ8WSe4Fh2wfMbIt21vqoSTpmFR8PkHft
8XoYTrXgOKXQj5HPAy9+Y5Bj3BaEMLOHQF1AiI3W4J5b4eNq+JN6LRJZ1NL1WrEeiimHNhkMaXX0
qCrf7hthXa58jWMjqnkxYERoJ2muGg/+3J9QcueMah84kkLmhydChl6/wJbB1m/PAMp9R/B2RdpZ
E4yXPbJk7JqX14nlza3MfyFUAvQ4pc13ilxiQSYVKcGNDbU7fGwUKBle8fnIh7QxtrlsS8cTYbRE
xVxYGsUqmpfjW466lQ934A0c3mFLKGNvPNkN2b5g4UdyFTiMLkuYQPDxoCzPM5Ya9uIgf1p4ePI/
lpMXVXzzIhDaJl/r6IYoiUSKKAKEoiOnm20nCiOPkXaHu2uXfHI1Hks93BvEuJGiTPSglImDE0Cs
pn7YFNethO2G4FIGG3vxLhOAPL45ynrgKRRDnmidlmbsDFnRyLQ5aeqbTMmWJu4GoEkJ0GNU2Ma7
vx8d2u//ImXIE5FEYcpUBE55aNSGMI6mmH+IO1Hf3hO+t/Im2zCV4eaWgr/BX4deQ25ShLeYKt4a
Z7gh/Dr4TPRuZdp8uGE+id+O3PsjfuSr/cdCEp5MsxsFr6pOufkBjMpWrPb09jp2FyJMbeWqmqny
++NsJvyV0HvrYdQT8zI0DY86qFFCwoaOmsxXPaayyn3bZU2hmh44sdE6RDW/FdL6lsIad7UlbgGf
4N3waJgScfvEUOJuYjjhkqzz2au3vx+CgkX3TdcqV1UcY9Ak0nvsgE6AUG7QazVsou91CTl5e0AF
lLzWNTQkuPn2A/vbPqnJ5TW1A2zHbCMvyjDtY2gu6/8wLsc6ZUf/k8ztrSXmXd3AIXVItdy9xO3B
ZWWXlz6V122peqeLPaW7bKSU0GmC4ZI0R603J+UM51xYeWsaPrpjMFXQxgYt9Ojv3BKDMfhUQzhj
xYfOcfDY5lrTzMSR/cnzjVMPfuqeGXTSClE+ZvzReQMXUM6gZ78HbHu6c1TvpYFKjEHfQR62U/ZI
w1u3R68mfel7mu6YBj6ve3yzZsnOGQWJZBW08xJNz4uSOImP3xySoE0Im9ndi0ak/yprym0FoDkq
PyKyDDL99FhcmOvdfgpLDhbPABfus9URa1GvDwVE0EveR93K/kwQfQJXrnY8Y3RG63UNAOiXsl6Y
fl9/ewZkDLZDxJtTQ5gG10Q3h5MS6m88AcKpaao77xXoyZk0Ufu3VAQSrXcDb7sI7YgHc98Aqr6N
tt2CuLjKxOdoYd5WrwpC3+qZALfkw5k2YvhzRCU7fgwZ/svGF6cbRZTZZpkYCKWFwoomVoEQsX3k
CwfJ/lsr16vTX7CxlVkFabnqOh8KEYejkllU/Shj7nIMp/M+gZ6hm6VJpVcTqH/R5ScmcwdOcZKg
or8nLPpGjv3C45qpgbnCvFOuUQpXwv6hAFNaQp8qkLh2kPLPgt4BL3oYT4zcMuiLymPiaMJbAW1G
0OPcZve1U7fb/TLJ4qluRXy/OptD8rGEXhVVfW9n/L3y4L88NM3t1rWXEot8gdJsIF1+w8lLEnfd
CK5yDfduOSj+vmeOHc5arKaimp/XYFGuaHd8yBjKPWOK60IROfjtFumGi2/784H89l0HqPkrzaXQ
9zqb0vBC0dCcV5h8CpzNe3/bIjHV1r3d5XHtf9lH+q90MJMV07YhlTijbf2nBrfOZZgO7fxn86KN
Mw1eZ56KxgN4PlP31DcVWQ/ER/KLvXg8nI+0aNrllEnNNz7+vrg3GmOSdLkKJSMvG8vwghDyVx0J
SljANgJrZM65mG8WQt9wqx2guPtyf+MEdXQl7/Rbg63nb46zkIOG83anNXCq8jRv4b3wMxfj/g4O
svasMoEB66KZLwLPq9TXsr5379yRZI3h/hM/3TxLI7qZP3hINAfR0JdywOq0PnbmKg9H/Jzmnt8s
Jq+3eB0jO2DrG0KLRdtVgXnBt64+Jh3wTLubtiTwyrAdfBp4/3zbnEoq50W2zMBF96uL87peF7TR
4owJauT2iEsUQ81AWjWi9bsSy+3EI0h/J0ixnlsNtUpUh/9JOdtoAd3UJEXln4vAasETb1lCCEjU
oMHzR5qgaGCtq3sCHnN1J8MzjskBIo0CuQFfUlaTnGJEZN7c0CQjDILQEcEyUZIfPWmf2djk0Xfn
F31v2p8aw840a8uIPqHMvfp8kMkbjEICT/JvgIwWEbeg2DxwXSILiTztn4RxNgBl31yxvElmUItG
3YtLIH9NdJhCYebpXdhqBEI1sFgwuIx7SJExHXsaWSENZNDwZ7DOA7+Tyo5QKl6q1DI0BQ+yz8Dm
JOFKR8gQr8riHEY1St1JeJS4NNT44KnPV8xZFFs6oJ5LGKazF+QGQ7fzKVa+UwjbL7gi2k0t1VXj
svl/3hyOCDVmH8YF68ko6PIxWuyp+CIYU+oPBOJvlJJ3bRSD875qRLk/nH+Amw2+wEsDGNxer8nn
BBDduVD/9eFfpngWdJqzpTvOs1OyzAI+Po0U/I3c879LnhLOK+WH0XmUzHfR8bHmzAzqB2N6RmWQ
2/pZBjd/4/miF/0+dE2qrpR45PGqJJaLZ8UqIa3tUSdDXz6NXcPeazV+dxJorIoIoi0Ni/Mt24Z/
RhMPh05BRxHkZYR3xNNR8TS7rJOPEqHew7KyXi55H7bbvUdd/alRiWnRxHR6x+R/dcqyrS/Srax9
TliSiXpR28jdDrC0Ewk3KR+ra0wCXK7QwH6PbXcwAj5CIBQ9vG0G1U7XmlNkHEy0MbvecuBLRZP5
aivjfyUtGnmOpuNQG5YhtGr3+94AP9f/J2gLWHxXo8U1Ng/ToJ4PO/ajQpb/IE7fC0Zm9s055uYw
fT7/N2q0NleQ+it8DJauXw2+H2mg7u8s35s2h5TPvQRsPeIQ6DpKBGc65y6CG9n/grqeO6v9IW9K
+b/b+m+hIDCiS/spcYn08VUoNYMQ9cIZ3NPqNFtJoXtv9LPJl9Wr0g6U2W9ZdgEnaXzwa4vL/Vgy
VFjRM6+8HUuhsOfAiSeWAHAsqWOSzz7mgEMtgpoKxlviiZsna9aUMhqUpd5Bc4WRJ6PIYbmJvisY
HJN7Rzbki8oNKp9nBkxM8U4eIQ0IEyjJE1qhFarqL/PMxgRlBz/ld37xLkN08AGD0tpEjP1yANMQ
0f+CxaWfpsv+XRQ9ouxopkH0BhBwtfYkIbqJVOfLuAjuEs4Ri99nnFclDivaxSburLup5j+3M0n4
x6JwArOQ/K4mIxL/LKfMuamm+hASTFTt3nJcxDP64Zx62RRLAcapopcRM81JoHXucsjqrJbK7gqb
D1CWmgs19gayEGWVaRFEIZl4sdStoc/VZIp2zdTwV6DmMz4AlG4sFdyqoZTC3EW43LaALVs1MET+
7yHBMmRFT221KYsr7WjvlPljW+RQx6TmG/C6W0AsHI0h1xD3q/mvYhuOsrrD5IIRqSFax7xSZX14
znhsw/MuuQ1oS4BF/dEUHnayqJ8zLacphbh1v2xbYqQvZuK0thXPC69VFbDmfhkeFdwY6uJc9otU
gapQ23FUOv7sebx8IHRGQj2e0WR3qWWcO4ANXHoZKoP+9l0LixcNNu8EpFAcWl9NKRgZvgux6/nm
Z6ab3S1403PXGHX5u6sRiv8jJWRfDhkq+tSasi+yiA+/kC1ChR7Nbu+aAk7jMDBVO2greuHe6Q96
e8Tu56Sby7DJKtDkctI9uwH6ThFcxKXr7SXDQyHnjqdykgqUEI3WFLbYjBhCG31KjMfDhYqdLWV8
GpxkZ0BI5NyT0puzR7R7Zgadgt5i+CHJI2Avk0ryheLIVprdsPmmVp9sgdRGpDUFOBuN38MdQ+xA
Z+XFxTc5mdZ0bA4DcoShLEJDbKzMVdRxEzPzo7BpV9fjJtJbZuiF1i0DuakLpWCZFPU3Od2yYC+2
/S+sxri82ECHb/qcqIUskHwLPI+D5vqz0CwQeqLKnzYY+V9zqZN8NZKZN5fWTRP7VztVngzArGsA
QZigQEOjmjZ/XcJBqyQjgRJnkvWUSqNyoaZTJrwaQm0qfCC8s6GaZfmONMY/vZkrV+7NQXNlO7bD
Gwk4SkBnl0P5pTChFJvJTMgfXgvU+igJ+SecpB0vSbZ7JgdxXlU9atfXcujCkIuG0i2PcaKuz6gu
K/94UHP49pffWtJG3ZfiaoCz9h+GPu5OFZ6hD3rvTaA22aAidPuaaB1CCy7CoulUAZB9QLJhQcNQ
qpvxtfRUjusfZ/zaA5FEpqo4upm7FEibxgYAxz4Yirm8EXBxV01i6WjkLq4qjbLw8i38IVKvZByo
xki6e0iyXhetva9QAE92nv6m4fE/sDZqMNtSPQlLbWj4GuuYEPXq6k7fuoXeUoESPKNjDs/slEP6
jZ2uMAnGfXlokmZAaZ+VldQo4ofEZfnv9DzWD0VEcnq+dzgcFdhYAc9ocXxx6wUScVJQmO4I6+HR
iF1SlUnBEe9YFwz4kGdeiZ1lcJhykfp0wW5/03KvbFA6/KRMtiYcLkWcc1lLNKN9tgaklsW1QJTi
+ZzWmDJU15nkYYkXSFh15NbKQX8Kij749rVdWRFvlJyEPl2JhOzdBs8djB1qe/V7egsEkxzTGc+V
ryu53F/eD9waJ11cJU09l4J6nj9QPwptSK9Oh1YAOtShqPCh+VhJBlz0MIwn65M+1IuyTHMX7d9p
L/ByVOfuLNMUEab8ElCq1aYDMB432DoLeQVNiBNP8e+m8e4p6SHb+QE6DUcN1sKhB8MCvVor4I7O
DrFXJ5mbvIIdrAF6OEV4Go7B6BIGvvPt9abcaYZf/hXjx0PjtjFyhrsqNx3LRlaHrmQIYalGvQmv
ZKRRE90QdRayGNqbsKqw/LlDmBiomoujl8WZVjNPc88m9P3gSzYmnKsEAAeLU0OSNM9nRXoopBm1
TxODqntzZRC0ROMCyZV3byvlO/+ScCbJ7VlD6y9vkKO/mYoGKMJjm809oeiKzp285pGdJBinBlDn
BU5O1ldDQYR1puvfK5C63VJoWj5G1yWiZ/nj/rZyFFCnMwJ14ZqQvCvSyUIF/MOf/IWahqWypWnZ
lticiJ3A3gOjJzNy/V3qTk2VSUHoJt0lYC7S1Lc9T1BV9h0+h//M3deR3oZ2P8zk2L013UgnBTgw
qSI/aX/AGV+A8w7uhQNU0Ck+ZQHBQ9iGmcHx+3SJLpWAmkgUNWQWm38wDxuSqijvpkHrGwst2ymU
+CteRSHfI10lKhgsoU2il+rSZV/QGor7GqiRpc7gQZBZ3rc17VE6DUDekqzhBP8ogAAOWsEqHIWm
66W4b8q+o/nXJG7KGTY/5sIuc3W+EPkhehzQmIHa7+BYPJNKXstOG8SvzEcFK7GxUQbk4Lf/XnTY
SbKmj1wpH14vgOFWdnzDgllq9FEhcAyPbwhxj/hm8rO5kemG8M10Pt1nSEyfgl6kZPr9oGtwEjiA
Bxq4xmiRPGjze/vX6/eG74SUJPMNyWhy43b9BkK4E4KFH3m+qtDu4iYpkf2yIoF3Tied/W4hDopk
qzo4+NyoOAXavFEQUi898zWMnkHsqDhYePjI0IPryBciq/FkKYw2DZ1vHL6bVgTcMlZUUD6nV++n
h++b/57nw0lYMCMju1SFlHEhJWfxZEiFD0M/k8wAG5iGpUwpJqV0DiC/dqS0ZS0Dk3yZLa7meP5d
CBMROC4c+pkUTw54FGbMR+gFYEBxFXwrnbpWqXg6azRdg7N4kIj7TZNN8zc3tzdhl5FzweXZ4A2B
fTEDA/JCMotIkgSM+zrceUtOq9m2hilZmg+kglxAy6kf6wUM1a09ECEMCeadH7pUvmlGal+QoZE1
Ung7DhudH55AZCJRxtci+hVKkLlh9VZS+fG0fT0qI1Canc4cEAHkJ7Wq+eDysxz6KA+Wt6xPcRVE
ExFYCJBHjM8R9B2Cv9taNrYH8uXjQjiOGx6kAUehDDTBhSRmLhyv2fja/BfbcX6p/fb17JahFQZp
Forf4ECXr2l5UPCZ5Hw2vUzs/D9EX0uvBt2Ddzn6KTLZrrRVp5GQCOexZVFTk1bp2447NNnsJt8s
GTlhG6rs6elntlidTB4GUTiPbcGuXoUCMu8CwEZGliuJ4apRzLj+MAPwHXwjA+xu/pGZopMr4Muk
E5qL3LNSACR0SccYFRae8+yyk4fQTeB8XYBHGT95D7I/s++NUujGdNqqwC2MuckUYyA49N8PBCRz
u6poMK6eW6e04137jc2LbDym7+LBcOnmg+ueQo+N4OFG3NG+gU1BJq12WLsdkNxwkQu10Ax8CVug
EZ3+CYUZA92PPejaqgmsi7GdZRzMK4QuvR88gY4yV3baiBvwXyseNE8knj5SQtYMbaD48c1pjbTQ
FPTXZCJRyk/OOT+B8KYuo5DbstFuzk9HejiJ4QkpbVAtK0FNYO8Xr6EBFfyUbu46TbrLTIpWKwEH
gqFvc+2X2vNIZcvHvYMjUz0UbZs1i4sw6xPyI7MfC911r8xg0HEcT6UdLFavGi+MTsx72oIpw74J
ISNoidP94ywtUB/ALRxF7YOpEUer2EH/F2EE3kDiDYn8v6EpLuB6MTXob3dyJv1blju9qKzCHm5x
rElbDykzUWew7ZjC3J5zOZq0vkX8oZlsUy8gEftUDBWPU8smNDKBBr9T1TriJ98ff1HDAUBoxWhj
7ihsejxJAHYT/hqpwgk6E+Gp6bwff0Hgchi/rrpYGU/CkXb72zATcAGD4iysiJ0GGfDWCiN7x+nr
i3HKNmtTfBGrcsdTm7Mg7C4F59NcAko5UV15SbTIEV7NuzUZZZjxb2YFdDu3cjeNPgpq/ZuekNCz
N/YF5FgDhHE8KWnINo0izMbVb+RGFOUY4Z47GSk7BkwXqsdigG/yc4nt6k2zrEnrcbU4RoBL+LTm
YHoTyjvXKm771HH3AE9nVYoM7FkZMzoDriPuNu3gBLJTbQedEPlGz22GVHTl5c3Bj8rfWdYFhEos
oEt58YSWRkElVCTXKt9CK4EiIHa4NjtMZfxrHu2cWOgOE/+8DwZi4n6bUqZ0X1xZ8pyPGTPMukxw
/+CrsJve2O9hjv3Pt/d+YLOWGFGbDGhOeGR7F5cZokcFf8HBxVzrDl9I5aks1sP5weLHyJa9CE5b
40mxpCFQWH7I69K2RuoCYV1pBBLRgs3UCFWwObSmoUqZdo0L8EccJqX7mGe4vZpUr76zI8sv40zQ
a4W88kL6H9wgVC6JZcyZ08JcwTxuhu+vPe1wPY8YxdgvMyyaw0K14Q9Sh+Cww9eypru0CINFVEb0
RKuHRPWieJWNNYqWfJGM+w4MVNqeNWPDNuPDecodP8j5U51SuQO/tJbpQTor1cW8T+BFaMMGOQyQ
L0GobLX//dfHc5LinJipH/zfaVrVmdDj+AuMLqAQ7vhLjW48Dga155opdtfSOssvnmLfg6fUxoZw
moETdOBZ7gMZMJArira3l8OPkaE9qSkYBZVT+19OUExAgjw/xDaY7ExXRAG3EbvtqX9JRRAe71BC
tok6/P3ibhI+ZSckZVf9AIPEkA6bovjlOaKJiAgs0W+fY1yqr1e+/mZ86vrMWSOxB5rv0dfAaVcT
1groWSLemvWOXd2hsosFsOHHdgAKtOy4q2vyJm4UoGU+ad1Qf1tVRWmokyb4rV90u32OHKbVQLHP
TpQlVMtElo7PCgEfb3eeLG852vl3c/SFjzC4hWTCP2aTEQXBFJ86axQ7Pz2EG+W9gnpdF6n68vF7
wpDGbCvarS+S721aaJuNw68lBKG1g/61MPn+JRoPexFOq6V8cs4XhlkkXX3JfO5UIfbaDmwij5OF
YSJbPk4fXSgVZl/1lDZGTv0pNVogXIffceN2sj95ibpvpQBKdF25j1/Ev9rZd72vH+jFUqER6+Hh
HX7CkFYZyoe6KNsUB7ebRU1P928OvFniZO83i8s9lttn1/PKjPtIYfacbiijyqfiwrvvhR2/bHgh
Si5tfVsiaBKhNtLXOCVhGmOCKhfyLuEVnhfma+kzdL1Yr9CiXxEiV6AGs0yMedNLy4bl5N3rVulb
6WovsacWLWfNGu5xJea8EML9y1k2ts1QWO9PQHTXHpWj5SuIcobDcqPxBgZEt9JGRDtgVjZoi2av
Dppown4LIuFCvZkjomWjq3ks8np8AxxaHrSs+jUn2JqU8H5/nPJ+u1ty1Y+LQ8tNcgf6bVPKaExW
ChOjJxqOmHNX0v0AG1WvgQSrhR8BbaRdZSX4aSn0ZL5leWRVFm+Y66A66/Uw/IyO3c0EI6th1re/
k1b6HiRPM4Z7unLjBwue9NWRfm+49SD5uhHumYfqiEHou29Ikw2jtSOARJHCBTactMgfcZN95G1P
Mlf81RkPPeYIUOrFfXNXU0VK21vQNgPL0kncXaAIQIQho7PZv7RRbm5uMvzS5RohLbVUTHjhSG8u
psc=
`pragma protect end_protected

// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
K+BWFWfBrBXLZRqrjFXzUDtjSyZA3EPRMD8EvRi0Z72an1SXuEBfqJq10dVOZCGs679TkYy+Rlrd
HzFcYe5nR4xKxFAp63kow7L/3sFX3fLDkdm+QlIgAN4pDF/yIIC/MwGKyzvRMUdpxNew/IPgbauo
hxD3lLhmG9a1PiDTv7StXLJVVhfupLrIRVM6TJ8nbMeD4VJIZKrqqgf5CBSkJ+09v7qBvXAoNH/b
0ntS8iSQjLeccISIpCnoBueZvYBxX5hkPARLkaykKigREkub7WVfZxisQHVJjW5b5cw56/WUfVH7
gPiahMf0K3K3k/L64WLEaBEpNHUzsuTHjc9l+w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 91072)
gRk7j8la6Xn27gBubHJx/jjzABob2FaUyrVBCjiiKI4NkHLwBUnnMo6srdSffcECytcJax0JK+3b
Kx85FisiwYj28qP42uuso9G9+6azzfDq67IpGjstgYgTZ49zOpe/Jn0xgWy6iOMa8FrKSNOi0nUO
/TC3j0tlTX+OV346JEzZtpr33UacGepYT3GtOfmF3Rd9tyuf0AqQgpDvcxijxPr38O2Al8fQznnZ
1oTCS2koaXEo040qFP483wsl9mG8b3Ht8gSFPYwuKk0/XuzWBIRXaMdjUBaWH2UaTUoL2XMXCj/E
izD3dCaYUVi0uWiaDJSlmJ0IVAlYKH7RhagT69fPDX94v8HYqt9os3OvwEzjxb3ZuyDH5i8Jyoye
A5HQZezpcGuMnjop2fwZOmoxx+yxbuOfgVfpnD1S+9Ifz7QHrrKXBtGe1Zzn1veaulC/MDaZu16U
yWu3UWayQuUloDXMkDjv59xDqWouKf77GucazThtgb7U+pBs+m4JisGmvc/trPVMnuNjCD2Fs//Z
txlEdeq0YsIRAvBEDT/rhcaDrrLlUx2aPg/21bKNoJfQiSliPvKnaQO0F9uAKVElGS6ILn33U7Fd
Pjlup12smGXkuEkNQnVeSyfpGjG0k5yemD4Zl9IT5s1Fkl/KLJZHi/j9H+SBwGuCJ0fFFSZ0uauI
4Ob5hyWBje8Qyf0X/HdeaoHUfuGbW4ZSklRX3qXQnV8dk/A8qbvOSM9ZEaxjqHkYquNLXY69PSmc
8cmRYPeTSeFaV1jiAP2//rpTFIukZc2ITZ3wlG9YvKiJgVTq8/u3gyMDN83ZyGDza2W4aqMJUsq4
ue0NImdR8h2llGyCKuQE/f4a4nXK9Eaoy19mAMj/7c3goDdxcZEeK6qap4oNGrzdTWBzuQtIy6TS
hSwoup2r0PqTWQ33RaPlJ17jHm1WfX/TzuKZMaesprpFyQ3qwd02r6Ub/jba493WkPJujh1mDCQF
oAMcd9eC1FtzJU8P+3Rii69xpfxIEme1Zf+PVaYRufhEEinyzw65GE39J6jw0jqCKXbNGamnHMKh
5To4Es5Mz6ysMjXylAf+NuCzk+q0fMKbAuPj+UDzr8+ZDEwHdtiUo3fsSYBl3DG9qxFilrjq0liX
eM7dG0VVapGxviTW0C6fzbE18Y3JrBGINsW7LaEmS/JKtF8CoIrwayzqXwd8BiXbxanBcwR9hgV5
2nEv5Fj6y6hWI05eh9y0eXmUbP3MITYUta6qiSbXfdIshCDi0mmuI2AUK2BG2nD8Xg6Lu70l3hWi
A2drjrxHhBTdkxGKTSEE6tqS0+OEeKCcTgtgxO2XxUO4aHowa25atbk+nHjwRkzyTF6GeT/oqTpX
yQMAqJG1TlBUXRxeQgpxeLaFfz8YAXnNFZwllPK6Os7unW9ViegmTQA01VJcGXR2XcbPitV9rjZX
uSNzX8bZ4jRRq6ZCAIHzWqntVoW6mrg815jIQlke85fLxIdxUnldqBd9lzaB3+KPoKKqbdbcS9cH
jN4/eZf9Wf63qiyBLwybWVKzfjfQkdpedxf/GR1G+hoky1DDcuZ0A/pIacIx1jTzm/kGzWoTUK1p
yG0iJxIBi2Bco3DPHBR9ZcUX97ZQ+59OW66lXkPSHMAmS4MIfwm7YeT+NoOVmvn/2AXRSBpMY73T
4Zc54YICrcg3x8HZTVOD4P4mmED9LTdGrC7r5JU8NteXqkcIeuMTsuunGkMb7MyLLs6q7oRU1vAg
WRV/i0N87sXPnGjdjiD5JWg1GR8Jmq0Xc4dSp8NaS7CV4CuuHu2xRaemzxM/2Risgl+hQob6ipqU
FPETGC1/WTn1nwJfMNOt6WDdZS+BudGRWlsvEr27HLBd/8ic6+h+DR5Xh8cd+5v+1/Qsr7+onNWK
HR8JquCHstQSJC7KX/6j9NlgjTdxa5iOIW6P71d1hIWcHPYfxYrP51GfH8N5yixzcsIIFAKHRB1t
bV1F8iCUvZmq3WoI4GcLjV9HqLr14/0wFmU9LLarH1bzxHGFLdyypVKaxOpz5Mdxo98Plpwmpwk0
eWFQbK+jtE41lM+20aUmD27gVLS+ndjOVnpW/8lw1COgohpSZPD2HSwCKqfHOKgzDQD30pxZrGx5
QfIsaEjfFRcIQfh0zGI4HyvhF297PsDoZavQMWrl59aVXZxRsNOvkMgRBz3aSmTT3klm3yDuL+ar
aggfcWxCz9jM2BDB4n80TxbEA07ANL6S5vZGXQq+M/FzzzZy05uor8SoOK6UN7k099EyW9Sbt9h6
cqmef+Or9cNZORggr3yBKRjl0FHf05hsTIfI2BTia5iYaHvGu6oQ4t6xEx2kdtdj+2lc6Ql/v3aU
OLq2iwkSk810qkIXqmYVGOvqTKSZSDs5FMK6HCnSibNzV7wVIaFGULh5UCM87883T0eUg29oaZ+l
mAsUKbp7FIwBH3lhmDa7R8AnUqygC11HGcYxnyy+J2K2UUlkNYVqSRKVN3ymQQdzAlcEJJWAsN7k
22p7JoyyAiCeJ62kE87ZO4LeMY1HW2IcI8RtsQO4InBfYJZSIibEQnxAfCUrTuZeDV3Hu6lB1QSw
D2PGmh2cPetqQT4loK7sf8xNnMUC5Fe39EXfHfzUn3ebdaDu7DdtlXurqJG9uyuPVNmwuLY4vMNc
jwOFY7ePMF1IGy8fPmyE9kt2MnhFBbOvWdn7Jv8UMCFcK4eJa4bb0uAOBUIuRWrqFOfzpFvwSBSs
cWVDnfTOgES7Wpv159gIWcOi9ReHQlVL9or66klC5m7QOiF5UGqYtdUPZPx13+uiDyR0mdNqBApj
X76ZX88O+kr+MU/qup+kryw8AD0c3l/UtPlYISjdeF+PVUlHW4W8oRBqsTglsQYLIzySQmetMI4A
8nAsx8YYqd77uJ7L5oNFSSjpcJ47R/sYTlSq95QmcgXSZWd9u4iEsBIE/jyhKEa1x+hivKpwhoew
KQXRi0fKa7gde6dioz6SNaXCWsdMus3XIO0Lc+0EbAgarTTa+CMyMO1LLYVKXWNEmXypX2KVs836
vyywzUkysqtW693l5ZiUb/yFx9NpvCeRt3FIQUYImHqLl7Xk/PueD0TPWURlKwAA9NypjEeHalLy
lT31jsLtFlopzDBMfndqwcNdjQRQrh12VzrB/BirJ0LbPUwYqNv4Wq8yNhVAyeniYqe5YmbKx0aR
LPEbMNEJ0yuV44iaEIcxsCBUMY11XQuuRQ4Kv1Sp2rTqkpmJpnvH8QoqWKrrKpMnIrvHGKMapWqt
0rqVxXUQaDWEVCFwsNqnUGnGrUWBqVW2LBptTESq3jp91LMSBNEhzE07yaT8GCmC5pywbMwX4KSh
W+QpJ0JDBOnZT+3R4Xf5iZH+fuKWOg8lU3ZcmuCEcUW5zatgbOfRAlLEI4qZgG8hXdRlwl9GP18J
UcR/c58M4qqAoQJMAIDiFPg9npwYVRoIYSJia+pAgPZJmS233gHKddHfx5QAYfRP9QRyZKVhbZQk
a+uwb1GDeXmD6bN/XCe8fZxkeQnDm8TeuVShaSkAcar22ZlLrS4AmRZ/61NniyIsvUuQISzyMoXv
hs2gkBnoOATzM21gIzyYpsvvR3bXbM4HRwTpFUiEV+0F9RzVMvnmZ1zDcapUev/doBqYc8dnehST
a9nF1d46vVmsnom8kgXkJrkfZKfBVc7fygSJvRDMA3Sqgl9D6Oy0zX9viItSKKogBrSovwkwHJvy
pHYdt2hmuTc2MHSQRp7BqioKl9wp8paSiYWp321DZbZRW+uO++8jH10W6yIhGpMJhkM8M0IQMxd/
v8fKsJOya6oqYEtiyfCkbZ0l/gZox3hFTpQ2rkkC5+Cl7JwkXEho7ihydNm7GCeuhX+TbPn75yad
2rBXnMH2rptSZkoUoIvUrUQW0pdrjD63DCFNbOr72hRV6MBGGIvbOorS4DtDdFH03pA8y8tLYJlk
HJo5GJXgAf3zXC/EG/Ngg5paj8Voy5EHuZ9S9X75KZBrLe74j54dMV388tMsNBwVIVgOHaiA13IL
x4rAYWV8VbmR+OxO6WIAZ6K6xUgUCyD5C/dwQvQq8hVyMRDUFTRCLpSrZ6WD0+wSYPk98gRYVk1k
HJwGrG0v2qyap7F5taKrmFf/JEuSAR+YO+Huqp3dRX1HzwWQa+gaxHkdWpOQ68HmOHrKcANo1hkr
odsOLEoLM8YcoGkE6LmCBKQlT5tdtm/DUmvP8R3326V1BWVZG7ZRZsciP5Dp7W9+/BX7glBjmtF4
yL1a3N3xndz34dVh7WDwAUV5hceTk/CUUyhk2SJrdcalXdGQRLu/LDjIMf/JxrlPDyoDEH2VcLkn
463TAXZZx0qQ6xNzoJKRBvL6YzICklV/tHaX4ObbXL1X4pLcZ7bcGFhG8XrGEgc1bwNG6LKJZPJs
Oq6mTVbFGwxEHmTePtJD4TBMX5WuOoXtGwqjIr8sKV8CL+5Miu1M6+YDuTIlLdOeIC4DLcxEY78C
UEN6nlRdX01cY2SPbvciaOnRBLi4GVbf4yrkFjip4aVJ9swE9fOfOHbQtKZmy5sq7124oZP0d5lr
NGvqN9jpc2PNOu6ml7HPOdmtMRmj4aPGYqF3e61LxZj5kV8HeBtUJitgC4FwqoA7NTO3LU0uoneh
JlbGCVDLXFVGJiGGRrCr+hA9O6QjWmDmMq+oRiLbohFTkb4cTcVZz8VF1x5/S1vXScqkiAkfugWk
im1h4AKF5bZsxHH7ZRerAHObcTpjbjqRtIx5YrkBVqcHwqtQR7f8KCMx0kZBvOm2aYZwVd9Q/bHu
y1vr2VXa7CGJPy9s7gCgUB/K59xonkbL4OYN4TwWbFdsrLVpVXyPPpiao5QbP7LPQH7iSG87UwQF
uq/Co27xWCQ2pt+/YzkRoLmrxk+wcrePfZ6tE98DUvLUE97FSb25ndiUKHgkjYN8FiruTN5GgPoz
4MnrO1vtfyLssIOSLr9nkSJWLiBLdRQS0e529ww4oPHABf5t2j+CrFswueWAISiCRGrJSIYAhEKq
QpJk0/HPqbCmwV+s8Mko6j3EJszhd4PrP/IGu4iSQ7UqguYGRM4LpDiDL+mILUZC+oTCSWsHnur1
nAKUt9OaclUDw+eDB/6oo2GrXiTUg7JJCbXnBZuEK9//VVcswlL84St6mujqOmixVrmFIDz/m0ih
iY3S4kJhqx/FGRgwcZBEyk3f5rJ4qiiwOOxmY04TDtZufyrvwzSHHt2H5R0EOTBTzGzV2PFlsCBT
s5Im4xbJ3FyS401aLk44TGsYFH0OyZvprp1S32XDBE2Z89eQKGMy0Gxb/XVMAcRtZR2h6h0Xh1fn
RakIjkBijsAfKHRdP6N8KNJQaxNeN2anq6A/i/jRjtoNWvGGDEI9LqttMZFoSyT4qwFb3kCmmJhZ
4ktz+eL31YChnWwDu5z9bDKe5jpMYXR6HW9aAxRM2GiQ+8qRP9wGnQ4PafA6JPIQjmrHy0A8JR9R
YIVCXD/LvjVnyxpEE0Fv3+Q0hovFtmQMOxhOW3D6j5k7zjgdTPBZOmHTdZaIaqX6mrQ0nn5wTEsQ
tfJWRWfWi8El0ocsT/e2Ap/DLg6wbNvag9A2dmOQvi79xIjLJf46EtMmTG/izlQhtOeJ8HMdIbtU
gS3nET891hElqVM+FAji2gPSDEhS5pAngokEqz0D8XNSMVnVfPdbJHjJdhWfrKBsOqtG5p16AH1b
HZ0xo89j+JXBnEnA9pv/KpAKnEvDNcf99/HIaIOCusSRJkY0XUT13Z83BkOSYzds1Ao3v2J2D/iN
gMA3lOJvecf/6A3EucZSTl6Kvj/ya5eWxgdzXaA/avQMWEDmcWPoeeIoziMGSzyphAdWhBo2q+af
VdhNNRhuk9iASX2Skh6nSLTSlhariixgUUlRjpgLeQTLvol+GP98ODwVW5IN2wERoPkvklQoBEOn
gaWrQSYp5T2ivND/EoA0C2o735HhqUJ/leERY90sbNZJBf7YFw7/DREcy7YjDvkPaY1/TISYhq6f
X7w/WQf7BWjSKhE4Y/dbZZgNslGSs7UXuQfVmV22od0WCfQbZriiktXa92bIsG5qri1zel4NZe4S
NUlr4yRZs3nz5K30Gz6JnjbpZNtoDBMt/NoVMqXhlvYOF8mm6iYfyOrzAR84CFnyB+k2+mQ69mk+
ydg/lASawEC/5vK1WkpxjkAaKuA+WazEe1iRWf3nBlD4IWW2Pi1aR4P7VbF72lA1/4lg3qJap2+y
TgpoOhVEVd1w79CMCZKdknN4HhHB6C0enR62NBRFcgEG2Fj+kXdEvLmMoLYqoN+9t0sxdRCk+zhq
Cfl7GhTB6xNQeqo/4ij7LKkujxEgMy0/MR/XPBeoQlVIQGhLQj5naLtFvl+Ww98oziX9cc0FB3Lc
cAmmQhSsrHCKHUJewKTj7VJFGTla+Hi6XHbT/8IUNWhKP7lOj2CdRFgo3Bg4YYuF3halDA1a7gN/
AsbuCUOk6IR90TLw5MK1J1kQQ3sIXHOhD5uJ0WehuRfAsViaoSQYteHYKpqu7or+G83Xd9iUqF7P
i76rZSIRK2DYz/Nd5C4O0VqzuLJw3njJ48vVAlSz51jqOPeSuSFWI/MS8KgFFoxLbabmybOVwY0a
kAvMRM67WkIh3Vr9ZEtc3Lr/q3lgtnJHp/vM3uIPDJ46wc4d8t9QJyUwdWitYR5246b0SWZMyoO7
VVh4RwS15rpgJ6l7AQcOy7bLhC+ayKtQTeM84zi7MLcomhHpe1TiJLsdLEFLzeCEEbzwKxk26Ws2
bD9v+QKeZTVKASUITUe1kAd4PL1076QisMTfmaii+3cfk3OyT8zBTDFnrjZmNcgN54CBmaVK3Cll
2eg0HB6AWL7c18m8HFICNOgnerBpo5SCVCPYWSK4P+KhXfSOHURh06R6cHCT0h06IOfYAWxm5Bba
a3JW4Ca/TG5ylyPf5AAT/vgnZk+NthlXjd2gvFYqS0ksj6ciNv2Ku3upKcs2m0pDNVmpCKv4E0Uv
JL+dJAqGkS/42qI+lauJQ0qRqzlSPofLCmPugnqsAhYHtS99s3wni3oLTYWt9cQc5utKpPLQU6WQ
HnJuvTQDk0dS/ZqdFyaGXrsPWSLFImY1oQOuvN7Qsgxpj0bc1rJcQsvFuW97aT8o4KYHZarOWLR2
gYS701hyOXz+8WQqYUm6rFmsEritZOF1FBuRsaM01Pf2MP4qoYEAx0GJ1NFQy32nSqKvTxPAM6bR
AvhPJuWaDbF6LJF+E54LKE+uG9jhmmN3H5JExXwzMYfTvF0wG4c0D2dm87+uHZfhwHxe4K+DfT9j
qvYnv4pxsk+Osq1auIvGhSAwSB5WMgJ+R99fv7Ey8JRr4yGvnvoR+Ll6R1y5cuG6j3w+62RZV/JU
n81QYHDwRSOZUqS5YUe37X+Xx1uBQCLFHxonVT9kyjQZN9QKEKp7mhSr84BvWKFFHqgJB/xNwbpq
8NFtS4AxmwWcTpNRGPQXOX3wspxQeVoOxTjZv7sw4gYchPLE0f4eWcvwrhiU/przn2vn9e2sB/Cm
sWfQkBjzBAJ9CN2kEH6tUC7J9r4rIqIsJCM+bsxhGYmNKAwvSH9jcEGe/6RIkbXSb5zgfyRwaeYF
LNh4ow23NbZ9svVtdQaTGbTF9Z0a4LBOZvzULtNCMc/fLFY8nwc36KKc6rk/ijf5iR9fBl/8+W+M
iAY3BoGG+Xky60F7O9+DIcYbe1GT/MDWAxpxGK6liXFpCrvWJyNJHO5GwFvMN1Wj2T3U0TZI9gx8
ZiPz+p3HFiOuiABIz65JjAWCLUw+rzVRmkJpGt2Oh+7gKbsWPekmY2UkLCKrTfoMSTWjtGmk7wPX
zCAs77dmS3wVjDVjvksucEThf8SBRBOIcmsefFh1GhnrHuteqkELNbPeSO8P2ultb/4UmOc7Uhal
Qp37YZtpUP0XTjpvtc7uIc+780l+Xgi7g/2ZM1yr1lLlbS/bmIqBET8zZl9rpXCtQbt9WCu1ZGQW
ukgeau8aOx+lR1MjH6CTScvjA8pLTMHOBXwmTnhGT8UnBHdpjNj/yJoYItDwZrzQtBJopN+Ym2ZE
zke5DKM1YDGlq3Z4GLIo7q19B0C1BuG1MDrmaSwkim+kPKcH7IExr2cIk5eiT+H1xcf8CgwioHX/
jazWJEcIDO+65tyrMvMXeB8N2vHUKBE+4993O93P1oxCDtWX8kVOAizktvpFHbm+aRyre2fromeJ
v4iO6LPCWXXlj0d6jQ86KyVSDynXl2IJKjp1O+58c6X6P3chYB7rENImE128XhOnyePJdXgvasPL
Hvv+Q+M3729YvNT++aHx7Ic8a68bCzezmL7qEOKr4RShvsRyukpEtegDYfZihZHHhl1g6JgZ2/th
gUq2YywtoF1li4X72OfBi523x6Wfe01S85E8rDBAsixcggdtedCB9xte4AldCkNz7/Y62VzZFATj
VwEXS/zYBpz8ly28DLTVIEOpvIArn/JRdXe+WsOfKVRDfU0NTyfq4h+TK0XUzkvHTSr9xF7+JZzZ
5CEz9/bZBxmhAUjH3qht5XZ7U98gQjA+Lno6Fj0KK5o5WRG5vWv/mLP9M//oWIDlfacS+k6TzbFb
UAm8vbFkSOcXUZl5im+AtgvQSs7d9fYu0yShXYlCSK2TtRXoO2CsdG6nudHntTjmdL5DU0RGByaP
Plzw+vhIX/a4316fHVJa1Vz+Rb5wledoFBlJL7QCwo4WEVTkc2ZOgeUtKI+XBdcpchBgsT9PwLds
qFOWslUaYCZN/Ek1s2MLJWy25XnFxK+rSGkxgrv9fu32y0ULRidZl91U3QuO1flSpxYIrARPKdUH
tqGZAnpRaGAFDuQu2R0ZNSKcZ5DVPs4M+csCQMexvZpvuZMUHrbmdjc2onYondN+2zuHMAZyuYOj
nUdtf03AS+4Zzoy4UTNe2g7TChGGnKf5fd/h24ifuE6UVY8/ok74X4JJZWAAOWMJ0G+UgrAw/1Th
5yflpFHrTr4zqd89VWw+ZDDPv4A+vnmUuSHUTMHE76V9l6ogyXmo91pWrlDqFsG9/Y8pHv7Ap5p3
4U4Ki8mKOQAemVwV1CfgPFg/eaS09YeJNJ4hjIJTEpREYH3C+L3RaDkIUemwm2mNK73o23ll1Uv3
Hs0LgIgceovOFHJMV8lwARk5ZT/jK+W3yx65Mf8daYeNfsRzE95M9eXmdNrOl2ZILs83hLTUywPE
94MVc+AgZGcr6pandYcTMO2eUIkplY7MkbzEEJC9gjkM9gEZqU93jX/V3AGGX+SL/Co0BYJYaLTa
CXA3RT2ZTA/dCkRpULkx2MpoU8Qb/sYoSxfmXNBxGCI9c0nlrn3aRAiWXaBaDyzC31jtW6vpDDzd
y9eDJ0Hi7N+H6F3L4ARK9dCzJ7nigiH6ZnvSg++QmogjxLsDiTJo9KDVDy5RuX640Rts5soOagww
6pmz/ErpZxUjOf10FfuHSwWzQf5HnpEU8zPL2jwhXqNFI2bmY18n6TIfzldPrU7jqEbrNkWHdEKn
Bwyoz8w4D8Q3jPN/9kt/dhCofPyZICoXuS1GhklEAGHrK6n6onfFwDLTSq9grqbTmzFS7f129kd1
SUZtUy7RxFHANoYRkUDiI6VcsHa3jc/M/ZxB/fGRnVllIh7Ae1Gm8klC9AGL97V/riGmlNs00jjM
IDhpffmKmLzVrtPkGFXeD9U6SkxXhWhzs46JzPdC7TkMKXsmWo6YQXkjWMuzNcYPeTciua1TZRKK
oGZR5xvjCt93lG7UY1+EVt4X2Xu57wLh+fqC2w2QXQ7wBV9NxdAgWxRPoGwVmXIpwIPfa7ly0DEh
v2UhiTZUf4h5vPRcL4ViQC0O6Wgi+cfViNZ1xTuVmjJpzHY3TvgkNBaRTsrOYrBLx/l6h/fre0KG
PkDOysEPGbR8XvnQcrLQu+rg+uVWdiLN16uocsS6dpkFoi8gWyrejbe8IKYSpne1VHqIO5WkD4fX
w7LpTeQFmj6KYH3bTPC4eWdHOup4G4+mkGpUm/0RlBJuUtiBKvphLRIOJ52N5LKc6skb2VxjB2Wc
ZcY//H5EY/vcHNTYyAGXUieGKlNv9VcaAZD+LCE8OJs9taeWsKbzGVfpSxBU9MBmZ19/l7TWQRR7
tK0ppj8oYVZhZeF1QYz8GdXa9sYp0lpqlUTGuT5AWGxI7nbMI0qL7ifm/Q4sGAT/Rsdf4RHamDhs
mAMpXdj2D0/D61jqgdmw11qCAXZWJMyLFYjsKJ1HfnYj2+lRe5mWLYaVRYxUh89i8gpN8Ei5/0j/
aaFLhXx+JceSCylgKGpi/L7EG6gAZANjcG+NWyDNT+sd/4zG8KaQztRMJszF5NjYb/aaZOlE4L5o
4kyXUwFWW4I31ZGB0oatFEsSFddQZupviVw7EOKJ/ps8JbhcQrgbRQTJ3qPOdUNPbBwlwN3iFx7e
MdRS8pwWxV9a/fCqOSQj4U/Y5AepBZPA+5+HDfwzwu02awAITCSXhzy1DMfKwwcrnvE5WFb/Kl7m
9vk5/wBJ9hNHdavQmjE9y0JnodFJUDogU5HcQmn7I6Kgolh08LxxSlKWLq+8bNs/ecdABXR5z4uO
CN17oyL0wQK9EopH5YAr0oir+pihuA9BF7u9gpNGm4w/jLSMwp3zcIy9LZRa9tq/nPnNRqmPFlHb
B9BkGet1qT5Z79dbg6VvrPtFh1IbQTACQ0hyF6tIZp8l6mvrAIxMf8VHOuYHQsi6d492etjQrU5A
G8SYO3S6jlIOPY2KSkekB7echIpnNeBHm8EiWWgBoBujgcD60OzxU12rySWDLyacli9FzVcWLC6l
jXZ1UI48mFqzFImQi5NswuhmL4AGYPvERsBKyBYaMUzga44aHKVhHslPLKTX6wI0VZ4jo02XO6dP
Ud5LxbCO3EpT87AkimbobfLc2ShGPHDFPFPv6DMRvgekRqkHP/4VL3cYrArb8tHwlRFc6jNeIL2B
F3TrmHn5hTHT5AyBbc7217im6ohvP/qWy3NuOdrHAkh+KFzNoQ+7UN7evd9hZVi3uyV9lhGgeD2S
3c6eJqlRUpKZO6TeH2cKJY/T0ybPnsemm/rMfcQaiPYfDp+W2RKJ9IZveGr2S5+yToShw36HWEfN
9bS8hg0+IdyDQfcmEKOL6WLZPAbBEZatRGzp48HF0EXBNqewc7EGaJrSCgSGldYQYQNYYrt421Us
F8pBiAtDI+RKoyBB2MusSxdI1fPN3eAYROjA2NGxYhUp5kkGXyDSPF5g4fag4Uf/aoVSS48NoPhG
i+s6Ytuw3zz4rV5LeUflei0Qik6/AJBTR1TyBsDGL2/JrqMtbZ1qtR2Chnd6PR1bp6AR7VL4llOs
SHWkYWMi9lr2f6IKy9fLBSZC5SVV+yPZhhzHpk5mid518/7ZfNdsS3IJ9hcavjeEhyoMED6sXXS3
zBfjc6Ds91qUEbPbLaL86doQWk5CtWvwPTKsDNU20PwnQAdl1Rtd8jhOuxZzGPyLtthKHmLBG85n
ATYvjKgmQBN1kAJhNyJIzZgt/yfpnb5hdYXWBQMkWILbnfCVjlxHX6rtdBViWAezxtQUCbs9M3Tq
mi2iZ2SSXC8GHD2tpAevqHwa/6G590QPEfIrIsq1FeA+AXE33gNJvJgjE6dR/1m8JaaJEBWSSef1
KUWJi1M16YPp1yi1MFWoF6wl694eUoAl5kQtx0g8pgjrGdu+nQfCVbaKzPW6opzJDsKq+Ch3eBoH
72Lub6wdfNZl/uSHoBM0VTwqwYVoY2fWW75O7c5jyUeqjHDuooChhESXyHu2Tt698Vn5tynOZP22
8+ziDLoLm5t9CS6mjjYTZ4bjE3Zb7XlG9ose9czJxjjoWasEj4KteAzuCrKQj/WY8m6KW7R8iyUi
bFcM3R72b1GiGpbePA9ZG4zdgYNhIlWu5v5gFGyz51euzNh5ckVZgAGFeUUuv6BnQJ3rM20KkMZF
V0AVILogCbkWpilbzYfGHV0b5tOvk7gF3ZBpZTf/XVMq15dLu87ZO+fbEKso//LIpCRKqu9pOkiJ
wWtPa9ym/jSky6/sVlePE2ioWJfWaSgg/4XL6BlKHI18wkosHv+6TV0MzO69s5L789juRMK6KWJP
nVyLtHZ/HSjygYKk9krw5Rbwg1G8v4xyHnZMo8YPzXiBSVF03EwNQC1uzuToUSrA5g9gb2ZoNVaH
FHsIa2gKar8ad/6CJp9JVhKmgl9zdpfxQOsjAxPAHoiWuvdVAWk4/q8EUwxummudTqHKI1upgAxI
Tvk4pOW3hgT9cX1tyZNxQ/4fR5beo9lRttOYTyfOuwxtY5HjUtQ9RvRTG4XuiE9/AdHGKiJOz90w
RBW7xYhTZSPIi6jEclAqYHs48YJAmj86oP31RHmy6ymaQqgLaCJwyJjq+4PO3ki+305jlDEZfLZy
xWqfq4QwwLEBrrn628WeQFKfYaLABNaovw7UWfo/v5X70yhPDhEJK6lVxa7I8Hy041qQkSFwca0Z
gwb2xEC4LTLXxZp9Fa+JQc8b8zXkhr7ptYCrTpCxkQsdSBBufPEzpI4QVtOGgxEVhtA2MIv0SVAt
WSjDYEr/ZwjjY1PAXCr0k3ze7XsUEGoArQJjv6/ynvjCk7oyBSg+BITAZymvQLq1QZSdgmljLVqC
eASGJp71gSq+dmY1vm2n8U6N+t38nubT7fOln2WX1ZUk1SSHuo3VbfYZeixyE1tVzepNneT6gbng
bC/5/z8J9lD37bqjjC4t35cA0iNxqntzUMUJSNpeinndRg6H2/mIWJF6dsm796e4tQUppYEbXA30
6NXQsV51oLUbAkz4i1rF61CHF3SXtJ0TT9enAvikzDi2lxJLwqres9IXqnfRs5KFxJaVhBNNhM5m
dRjRk3gj0qwRT/K3ey7AjsXc7HXK+25Lq1SgHri5HPyimqbTHGDsNYTKR/5eZVxlP3x3ySndXlOg
hoSp/AnW5s8DOGcCd909aVuTls1UYe7qEU9hLFQgici6KGVeXAFh+TNs3lsRqREljgtZpguYeDFO
TiUEuFMa+ZjJ2cVo3Sui1fcVEJhovJKjCiwxfYStlVJGEW0bZAbkPAS6bden0GGUW9l4X+iOsv29
WADXNyraqhXUWOWvEmfEi83ztESY7PoB8nIyK7X8BPk58lD66R0+LTptqf44zjmXB+gTkrCzDZHE
9ml0OjL+s5MJSHy3V7dFgIpVeaT0uNqzYs6hVn0AmUMZ7RGd6r+Xgb62S6YJaTqfVgBpt0j4SJJq
3ypahZHYRbaATPkYj/2ygrM19KrrYA+XKBHa+AOj6E6YSWJLh2LOPBV9D60jkF5t+sg8Y9JSsrnN
xVP5EIYzdrZBnFyBrLYTP3mEE9qfQv17XcnkPXnVxzDJ48qpfhBPENnIjWEuFVbPhiWfpb/up+qB
Od8+jgXu9RrrLe+dtZr1HbW3A+cj+sgzE5s99I569zrmKZ56eBjf8Yo1aC3ro5t9m2pPI8Rfs6l1
y/JcG/VVKjHBflulAFvD49qEiBjbQrsfEwVQTg73J4d9cQ/iwudg1vlGc1X5TtsVzK8rr0ghzlqy
IEYrPknLEBfwIuAQCZw9+hwGAJ713bEAcYhqRdLJMWMaioS1daZd3As3QtnxY8iF0zCCM/IgdZbS
SmxQ/rn45/OPtb6tka7V+TrEDyabU6Q2BMDDmKSfX+oTavUj+MGS/Y3jPQnKeh36OIPpD+dXHMjn
mXfn+p4JD8nl21veYbe530atzFpRcGj1ROBqrqshq0aO+5zdflA1xS+GwMFTbT7LGhhE25z3qjJA
OcB7TKR9DvOfu66h7FeHvaTsUXLe1VDfgcwFWypLCI8Mc35n13zFMPJfXB2QJBbXR55PezS4ZyxH
33y4gIXoso4OYIsQdxdJnTGtJCLmrBHsfN5iw6e/jC+DrRS22uqINSaHeZ9Aa42Zb8c4HcyowyVk
VB9zRM4DIIVIt8SsPpsXgP+5znoAPD5ae4LRZ4TUsc+n/HmiKbR8ZucoGoVeWaYUL8cWHvtJWUqF
b/0AnbIEWvVZq9G4adELGyP02cPAqK6JxEA0zDPsTxCU3t07OJBQknpGHgha2PBjZ+0vovdfaRWq
tZHTKExmE/mxs/2QQ3UAeH1BfBY+57MZ6Ae+ziun9Krrt11+9SMJaEhyEEkxZbVxu8qCTmll42OZ
RuTGyNg4nyCX4jDVF3NcS25R9tr/hDXkdvUwVF3CKhp1gVlV5tqMAUQAWv74bNQWeixmS4bg7VXQ
fsb1uyXa7EoC5JrVcAocnJEJlDQETJgzBAojYJs8e7V9nFZtOWlnYMXbJCXPm786LCGS+i5dVJZ5
LZGw48wTl4kV12EgW8tlb3KM3kbSVpdpxDJt4uzRcVCL7bOj0Fb+d6qHU3SZwxvlAJEGsOfN9twD
rQE/DQFK9YUqGcuXgzgb9fevoB40d+KxFq1h2GsowQQw8Yu/q5qNBaaLwpktEqzBOjaP0v9W32tS
pryup5o+8k+UsOlUSdCmazwQbTBwt7bH4eq3D8vilfCxh+XakZYYN3bmAYdG3xefoF9eHwISF4Ol
cbfQzmsRbFURt6zjSTbHv7rRCPedf/CQ9kv8FZp4T/1Rued+E+sW3mzva5qIaASdkDMrJEzwSfy5
ds+RCIFVmb/xNs4+XjGJsDUiJBi7+y3J1rditgXmGd0B4Fgr96YartZ2T5qeSl4O+vln2Y+rXdNb
Haa12Z7bZCcnqUHPjyy1XYsAVIKH1czbWln9KBL5+rAiNXd6ehe5YZfR78ctYX/tlRI5gSklf+3f
RoWtQmqmjBSZR5VSIHy1AGRe5ihMr+RzyNZKhlhn32leuUtBPAiSL7XFch7XGX/NQkX/3gqD5Bkh
OnSQs1x0ajxoz8UKxmFWkhvf8oPslZO+b7hwqPh5IE1ad3tUjilkgmiSH1TP/wYGlygZ2LeEkpGO
u0PEJ7RslRZFWe6N41doFCmtQF6TGCuKua51rlK/vV8VFH7yp+jOJRHViStvkLyQIKwBN+fSysyp
7VNQWG54UzSBzsj8ifr2JoLMVNnMIM6j3h0RWzPAptkjgLQNsA66yBC5UkkVqjXyfnG53IhpRCg8
NWEu5oYmK18Z+TUKoYqgUmhVoirsQnQygQ62zZ2lVAqjV2HhSDVF9dxgPeT8EMx9UJRR4c+bYGnk
79xsQm4396QyjPwoy5yKC1sz2HCXpnJmMHhnEuHV+WJi872X5QPp7BYNJo5ioJcVqm+8GjWINgx0
WMp1XmJJDr5co7+XVNXFNOdUu4Roim65N28E5V8Cag56FWI5GDuwRCtA+s7M7FcChJABOHZCdgtv
/rsAp8gdEdmAcwgPYu+GuJ70UUs8tlBx4j1yLAQHcRV0AijxDShBF2NqLbIk2oYmnwLbf6fUEnXl
mb6JJbJSgtihPUWnWLpZ24Sfy3F/wDNau2y9CiI+WlWKEK+GJugAlTroIrSOUphnSeZoKx7ENsAJ
GuojwKXMbpSIxkHvtjicNNvRg2qU6YWvW9NMO7CZ8KBg3fA5PEl6Joht4Ow/JNjvDXK6hRUgqAX5
4vyMFl8g5Dq0SnYaz59Oxc1DbPsEnyAmiOWD7WDDR+rY9C9X8jRKG8zxcuWsmwVqbQZogyWoAXzm
WJGc/Ro/1cihjmiBiQxfFgWwl0v3zv7IBiRmOUQvxdyjKy5TCmG4uNpAIjlVpFHIt1NJvQrWQR50
g98g0bjljKTQUqtlO790rudtQzlxbktMft4JdCkc5OCNhHybRH6iOh7Omwacy2fJnwPUkxq7DzSj
wUZ/A5WG7tz6+gR8s7PzH0AhVw5A9UnjVUrC+rrPW109+o+JVaoGOyzpHTnUcBl/xrCs9099jOiw
EKbkPxNUMNBVBAXSeOCRYFypQkEEgsneKLNYjewtgRAm6gqvQkE/aaLRYB1RyBYI+b9shv48+9eu
yqC9C6NLdbKhqkxkOotbi+lYqAp05r2An5PZyk7EF3PKrY2j/SeNEvqcDxM5MqMnShM+sOe0EYK0
9U5IssMWEqGzLA9RTmM6FumU6LSJT5IxuPbwIc69R4y2EBY9eH+JS/jM600/VaKlUht5DfbmWgMF
OybzaxbCQ1c+zWZ1Il+RB+yJoqZloH8DQ7bJ9O5R/c7ukilc2O7Hq/JRKw/Nc5Gdboe07+qM0K5l
oMDBEh7++TX8e7p/xXO9egAWqUy8CVV4EwHeiDBG5ZzIRJhedNmMMiA2W1jSbD2kifnbtgQrE+yP
BBuvys/+8bgvvfRX7rRuDYKv0E2VM3omO6LhyBOce7hn9YOSw+rQRLwZrdPH/RdIc9/9TnCwuotD
H5JBGbs+xRkiv9UvPChKSNvu9GsV7be1LZ5DgEiwcrmgGjE/NgI9rwbuMDz9QoaCMeiZI2Ckj4EP
62xBzIdcNXPJJ8rr861V+inQupGSiKEQUUTyliq4OrKjpg0RiTlezPqXu5QuQXLFcRBhQPMyvikU
klfJXMKhsjxZbqmgWlGkiZGrV4+ECpkhshzXROlYE4qLz91t+hQ1ZRoncrkAL2lEUiUHb6MbSQb/
tjPveD8UzXn02KizX33ThnE4u/nIzSREgMcOUIuoEkyoPNRK2vqZ0559VK9cokPh5/evVzimVmRM
dJc0h1l+CH8pTJPqdN5QZmQ28Un/Otgntf4RJOV8jcB3UZ7zRFOcphbZmCYAQ0iWb4+hm/TjdTRQ
3riuFKDUKE+tRHmcmGJLpeFRZ/wDbYyvpqt95d3LIsnAE17bo4FlnCxuyOTuHDYuOT0sY8mqf71w
91NY2Fc2RfzYSTEY+buyXcTu3PkOq8TIR/53DcCNJPgLKg4EWndKLXxrSREoUuhiMsLm3Jwp9XTj
ON1h8z2ep5Yq7uEOnuV8DLKRWevey/i6efcjF2oVb3Je0aOnXpgCSNgqeTBUHlHRoIbsDeKS8rWu
qbLRYspVvgB7QV76ea5Xhm7sqizibErNkU3iDyAj45LxRVkF83uhaT1XKApYT2MTXJADTjohxMFI
xNuvoahmtu6oTWXBp7V3B8HCUUkGRwBdd6wXPRZmTFx0ErI2QCB/L/v3eBtYRADUeIeDzUrOWj+V
4kkK6HzB4XVY9zlFV3OG5X7pVKmLgxNvAG7CyaeeNMXQ6O92GX36snvhSVjI8Wu/DEvYrI8jVZR4
vQQNIjzP393coRu4iAAga4lRix1pYEfreg3N1Isl+d/pz4r+8CnvrHMNPAJ4TC/HdM1uhjqhOehK
xkzDiwNuP9Wgvwq3yCi8xPLlabBnkW9P94lzHqCWCUeL5rA8aZsC2yFgThlNFR9PGsIQiKu7Jede
ZrNVm4dHTtRN+0ntay7x6qapEKKY/LFla+97Kg2Y05VoarVRnbW4+XKVv26mixihibdW2/3Ce1UV
E2IH/gntVcQr655XpAV/2gNP8gqXIUXNbV/OIch5yj46LZFm1hm+5Y3QlmUf5N/flUsSZoO1T/cL
dLBxuhXsuyAFtKtO7WTECeZ3c6PgGgccKiF7Xu+XIe1Iwl5BAElRZq+IBQ8aJG0fu+adHsFm1cM2
ZAQtbM/pKK3fU8bMLeNcmaVjhZKGFaoi8vSIiSJIZSyYB1cIXI4LXlunIU3xpMsz8MreaiXWqpsU
LMsy4q8lDgd/hJn0zIDO3FQGM6aigQvixOqi9FHwf71IpO/lj9DwZRBHcPOcIccyg0NssVqN7ZAC
JjCQ2G1wrcoh43vZqRy5LXBY7NGnrDKxE+akGQ5q2of2R0mxSGE3mIH155OrIieNa92FcjalwQWV
MCNAZYGGM6/rxcm7qayJe/tK8/vPwaJwo5W4nQaOSYostXyyceh1Nc39B3W8I07VuY6WZ9iRE6s6
IajdG3im9SNuEbWpQMtubqfMyvWQrtFhZHJEFWyOGviuRdzVOb/Tyu8Vc75k8TEBPoHUH/sxGJ99
CrQB3stNMej+tWEun4UVoabAe4uA9o+D13E7d/pWudfp9zxLqOhfTDPCitqObNIcjb5PwYmigKB+
BltRG+iLzLTtf2odqKmgOD8d8d4noyawUBBmw/kdKXdlG3FoqVsBXpvJORZw50f++qjxyzfY5vc5
KRBgAubMR9FQdYBQH/K70VlLH39VQd80yfPrQh/xkctRLSth9hfOwdcjeNOLKNxYMzplOXuNg17z
lbhXi9wZTqYBqP7p6b+4DIkuAJnScob+JAV5AGEKDxKmI0J0Z8EBZGt3qbnNL/DhtPl+rXgrPPWD
9dZhjeAJ2zZZyxJyPfxhmf9wK5ZNfTL/sGlks+oAUiowHN4ACstUB3AYZswqnnvXbSJEpigdJNbG
GR51cQaE5MeqAV5feIZRuP+S8cpKrDSOxviyuefmrxLsuPb8gkv+hqFgPr3yMqR1J+kumwuKhaiV
q7jtSaJLGDUoGuHm5m7Es3lG4cwO5hS1Tzo64zvp34vFtAWhz1HYi+V/KbDNOtH/HUiD1qtPeH6m
UDyFb73x42TR4uqWThjWu88OCZebSZnVtLqvUXhdOy5j8wN9DpdDAEpzJpvjYtmrpsDrJrWPbdYi
4boAr55waDL8pyte0FNWOtT8FaG6ARn89eN132zG+zz7cV3S54iem8WOwsPpKOl1q9yTv7Rt5r1a
cu2ikA6XvHrcCS6MdOfYeJUqwofSFvIExGlHYvIpjaXN3xDVhTU6QvDUEtrsxhySeFTpRvoRq39V
BtaFG/5l3IRXEbw8YGUodS2z3WKPlQSrNM0Hjz46sHYUNuce0tHw6rMAFVk7Pha+xQ8AO1FyhXAO
jWufk8VZpXrur3NmGnyt3oCYJyCLpyg9SVnkQz/9CblH+2gst0L8nSPg3fMfC86AybGojudbywXu
BiPUP1rJI2tUkd0izHcPAb1RSHl8K4aVYMwxbOZ6W/uhtrEnPATyN5clBi8cf8pBst5lPd++aKAW
THECyqwWEOhFHFwF2HRi0rtA5ufxpOR+qYoLmJo/0rvnnGrfvpbespz8kMm3IzaX8tDXAJ2UVXE9
UyZYreON28pwFdblFWhr/EtLJDitE5V8FsIbXFkFSCBcBquSIlfkALhZHzSIe9di8atX10VMfU++
xlKz4vb3tI+61a5ToLWLt1LcnN7pGlHXwBvfQdsGxNb7e1omm+2CyDYFPlJP8rqqqbTYxUDbz9N9
5Ap7UXxCY4v530y8/0SfYdueJWMh8eyf1+fSMs+GH0AJqWaXwSdE/b8g5Ope+TDAZzr6gqHUI7wK
rtfzY08PcLiPP/AjGKTic0qW6CoX7JLnnIHF2QcPvkGa/mjHuQjA2Bj12GNq70f0EP6U8eFCQkcZ
BT4cK+y8eDdVTEOixczvo6JtQUymjZeutsqZn4BY/zwY0QBWegn4MZeiIvNxG8zAdPsw0ATkXHVl
CSiUcIgEFFqKU/F9XgCU9BufW+wYWqkTg6xtL0VqCVx/0eelTeJ/muPYTNTEpbCdDBF9yg1/3Due
98Q1PE86EqAytT784c9kMfgHGXshT9owTVKrp+nf6DmRmQ6QLIYwOOzFztnD6CltvjVaBgjLOUgV
1oNf9w3B81rslSHfd3BtM4VxVOjVCBvebh2T/WYdyWQz2JN/uC1Foe3duDEmlx3IBgtjcCGR0o/g
su+vwriVa460qmt5gOfKPi6KKQ5VbaozGoVD41jcwez0ET/UTO/rcSuez0QkrslF7kPUcXkbLfdS
6qMzClc5uf6bXZ7kOe8aKz/h/nhfaBZzNvYodxLdlbb6uOt05IA5aJDeuryxlTVu6RQA2ggWWSdw
1nsfV5m3KK3fW2CHAH1QhHALzKTZGp2Jl37cfK5WSRdlbgfv+ai7y8Vfuz3frsY/HBp0rMrfyQ01
Mfx8dQk8RMndNU3XwzGDmkAxUfuv+YboXv2TWMjr6TMMXg4DsnWGoKQiDctHUPmYgmWU52nhgIW0
nG8XS5NOVHmYO+mzeJucnIf59OHpjgZJtG82QSXdr6d5038YBERD5m8t5B0q3yTBp/L8nr/NFz2W
Pr9H9S6NnOtrA3LUD2RvtaDjhSJ3xxVypgly/jyr8HbifkuxuhfklE1o8wuJEp/njzCRib4ZdnkT
qivqFfJ4PqgdSCP1+0GRz8dxepBWuIQZIMLMNTQzsGT4+5q4vvjFrM4GlZ3PctR/+pKLKWbAzmw4
+KHmHRSYBK8Mp/kzcHbOtdfQaeCG2zxFoawNLqjkdgNCxoeK7edRdwDdpsS2k7vQhfHlTpY91dWS
ayFMwOsvIdBysRaBotAymMBtesOI4/XQN8T71HmHtBKCuqMNH2jCZTxyVsKentcwpN2s6QO9EWII
B9b4D8Y+mbaTU8y6Vp/mN5BzbdNv2E73Q6cqK1YgRgHmuUEOfYUCny/sPKD+F/vvz4z83mC/PLgc
yK0v475HM9SXrUPiKBQievSuxe6FoQE3dhU0/e6BZQ5w5ufIUqO08grXGlq/+rVxKmiDJNS1TUAJ
bU4RbBHNqtybe4ZdJ51xcTTR2EXWXy6SQrNgK7jPveDl+xxg1MJGTdCHp2Yg+EBzJZcLVZVufnL/
t7nBedeyy+68j8b/j5fMyzMxHOMf60gCghrBiA0QB12wFMp0UUraBrC6zN1DnzPL9Ri/4iZ+eZuq
1xjaN0WqydFGVWdPlGPjmHE0kExDwSy33pkuP7UJzX+ak9FfAR+SvgNqnYwwb5ntiOTXmkeiQXOt
tGccA4YPVgBAuwamlT9vuhAmVUpxKXOGumC/9mG+TAxdnOuJsYOXn9h8OWA/U3t6DiOsNVhPRCdj
suRAGpZygwyPCdo89eCuSHUKEARm6txZZYw9xRyV8BRWkxe/f4yfCHXGkq92sORiUoA2vYMj2x6B
gEZRruHHESX4k2+PRBvc60XlZddV0JSNEAlX1806NOD0ftfYb/AvFnIJSYsHZc131+FDis0709ji
mNQky1k1ZCFS2ENymntKzXhxBd6v3Fy07VeiZWIBYIj1WvpodfJfVtyEsIvlDgN/QpYlrXhW1KrL
vLWmj7w3WA0qMtse2pJojYNmAZVRYDYe0Em+hfIiInyafjnh+ctIFUBP5yKkcY6FYwmKreGJFS0S
O3oif3qWLgX8nxGdauJcn1UiUKpsKISTF6fOaaCDcLZ3evV0QfLZDkkgoxormYy5WoFjOBpD5P07
7Y4m50v6sJDwuoXJdjJhNorQonkfgO8MKyv7WqCaoCUwe2CfGeE2hDpbRgM6OIEfFw3+AlrQm+dL
x2/sK9q3IruvZ6x0/V5sOaOB5dWl+quCzR4heGNmYTdWTOOAD+HlUWJFjLsg2fogKTpne6nH532l
36pVXS8tUrUcclg0oye8sps/7EpaLW3ua5c9YXklMxbSnCH5kFKphT5oIZun+oAu1yPMD8OLq00c
y4xM2EkXq4HX+IzrXARGEVHDqv8XShEw83LVgN1HRSw1838iuZ51jWHxzvS5np91/r8JuSJj0uo9
5myp2oABpgXjuX7ApRvUW/5m5l0+csqb83bzS6222S90ge/42ngum1QFriRZ7jKIMOdwpzuWdNTB
XrNUh8VDjT/YK7Skm9rxoA26AK5Sf9BNbwbfaXVqaMnaS0EjxAIlsG2r1Vcbk8DJSuoUY2cqtWXr
geDOnrzXGo+wzf0s1O5+dCLMGqXUOf6yLMldrn8J5hMn94H8/UV8d3fjeZyK0GmZiKwj+FvoKlt1
3aItZZUphBfdAGoMdMtO7ELkNQDZ4Rssc1rC/UWb9MZK62aWGpdZAmflXd5f2pu3ruBFXwfUTQbp
dvnKrlrJWhiz6+w2jTFPYKZBfZcLSA6BUECNZlEH5SHJMGaACTEzIpQRon0oZU44H1HrKNEqgcrF
ySZ4W1RXO50fcDrWQ3kCCTMTHjnc9Ait2z7gxZIqYMdYim8ygSbsE8aLNe0C90fNxsBqDZz5zXko
LkQCUkcQZ2Ogo2zGswls+qcEI03V9cmt5sq+ndf+8i0Pa6ddvfxon2wney42rl56j3lxiNL4Zbdx
7RzQoukAx80UVXqX8GU2jIQH0lrkSSQLJiF23cpb/lV0UjO7zps1Ckopnsh4FhH4VAgS8dG6R8we
sF13jIWEmG+VKR3XeQDwHe9LhdydBytnVgKlvNcMhLgS3vIKizWMJZlQi3sBTwR4FE6FrCWcoSVF
QXWVdmccwGkNd35m2sklVSuM/d6tK3jd1giFcJ/yP1gom1srtA+xC2atLT4cB8bs/xGDyUi7E5CV
itrYPVRqoxZw/73QZFzWeRyZM7lH7x9o6Nkkx2+BkapeiVdP8OnttsMFctOu4Z4lyMlJQemm6S4a
TofW72oO9su/hl0Cm5yEd600Ax3M0Z8Xz2m/PlN5BAFUjsNrBKp9Wo1m0hPlvvW57MIRPShlDfBI
U7oy08LMzXtG4X+uAgSEkNTImk3K6TKkPwV8gMv8fcAbHbbZ/NgCzU5HlgI4a0Ws4Rn9/8zEAikK
3zXSS6mLdk0bQADuDAeatrttZW6OnYjtMFvrvgmR3hy1SwQ1Zfqoj9eyOgRtGp6VTHFYejnPRiVN
kUJox4hTUjw7b8r6P/NwjCq9KTZIk1i6owPr29xXYiER/GtIPFLPA84Hbg6oPZz3SHwp7jUgB4ON
vEruZRZHHn+F3p8ELl47wJcy4BYY5KsM4Cl0CwRSZNPSkWndLygacQYYjeULQxofp+u6PF860Q0K
oUflU9uC8DQBW43autlDEx+cZfUJ9LAL0OaP4LBJx3JZVFyYwA9RCpw0RftNo8zXZSyiWWcwmxwp
VOw+gIDH18QQYZx02NqBpX96q8VDi8oDnOqoGV6nCf1PDIAfQGB3YxDnnTaKIDal5xUDdkBAGLdo
vTtNip7XErCTxLExUKKVzv8O2qxB3EIWAecYLBgkt/wCl5vEYRgJXNWjYPpzgHWkAxB12PfyfqpL
qqFhrZtRRxN24MgJJiQ3rAmbeD4qMLa5NVBCX0uqqBLhktdqO1WBLvEBfYUwqzQFJSJRsGMmaGLw
kkmGQRQ0aVgRyZkOhjL7NpV3bLU2PoZftIQ1DYHzYy87niqpuHw9J5nn29QZM+Trt3K39/KOAPWV
CJb0CgqRGF9G4by3h/KRlZG5F0lfWPhdi3GG6T9WL0iWRSW39rQ1bLbCFmKtZyYcGbM9b8ZrmX/F
caAMuy/Vwx6hPds5B1mRH09eGsNR7L1UravquPw7gSPjDpgrWK87J/5NhDK95DIZD+luVL0Ua4Q0
gOZ03Jkj2uM3MvQPQQu2Az/PqpfR9wdjUUg0bELi9R04HQKpmzh1UbEkrw7LcEuW11Z7jHpgKvdf
WcS/DXuXINwdgmtZJ0VT6/fjojKMvyOnzQkHvm6fExOPng+K5yzlI17rbvuEs1DCpHzlbBW9maNb
sjYHYFCyKTg2A8Zn11yiiZjxr7CKHgSn4DmvEJ+Q5h9Q3eVWoNrs73AIllU+/cO0HFdM0B6lGkHe
haT4bNY2MXQsGTfCskJNUmWpkRIxIkXRy8q1c0LxzC4xCqwyoqNR2/7l3ylyaoXGCbT96gIzJqFX
bExi58viVyI9g9ELuA0lTzm6sf0CbwDRYeCpCJF2vpv7PsZiSLPoLIkPJrHyC9MAXqsGgo7BN/qj
IOpP3rzuLH+gsTeglDV6Y8hiSJgT928DHxpbl1ohgVcsx63wQPj2THlNLRtB8xO0r+f9sDD+kY1x
tbfti8TFOwgL8SAVHZkssCRxQeZVqkXGhr34eFxa3GE30gsgtPIReNvp09v6bR6k861Mz/sFDor3
2pHSsBdpA/scrLNC0uzg2sqjnVS3efV0pq5nT5+k+IeuZVvgHTR+AhlgJh6JvUkMG4PLrDajMEXS
mT+qxAzQ0tPWYH14+icuHR6n9Yw4v9t+TBfoVNI/fugIWb9NGVMAGwTHqOcS3+mNzCnL+DPDQTAW
4IgC1m2FpoG9EEUVNSI11P6AIzPKipLdFZpKV4hI7UOc1VCHXAWuu4+cLm+9+VGLOFgShiA8WmeG
/UV8w3Pxm1v1r0cijrVk5evALKfHhMI5awcDKyK+hQgV5cDo2mCZxbV3JZMSU8M+DJ91I1bpkmTg
Kko3xSVrUV6/uZrIJaOBwvLpnDkb2q9ZH6TSmXY5yevb5BeiUzr89owPGKMpz+FwRNkrfqiMqPSV
QXXWpzuICT/E2z8QFp+wACw4EN6uEDKNBhRKzkWAGaXXgg7tThrvbdrCnYrzUdhS+73Jt/VoMI6U
TW2fT/VZQMUd/aXuTOYMZ+6sWDaS1ygbe6gH8gb4dLKVkJsB64yer1SMtbwg3NtHlnbdbLu1jg+4
l+BbLtyCqFHL2dIKyAZmTexbo3dxpnxMcDPqGMqt0hzqioAwzvh7I4bAg/JVlFR2Sblms2su6fbG
9AuUI1oMCtVeTeMFU8mm8UScNzrfePI0Vd8aM3v01Z03/imQClbA95cVC0LkKwMWHRP5BT/TQEfs
9uIM/+AeJ6gtF/BOOdFc5IQvuA7eMQ+r3fZ7v80IJH+mHthMNBgdJQNpj9TOz43+hJIFPvLb2YqW
VYfAAgeBhRRIHONl/xQ0orCaln2ZxqnrnuRueTGjXrKXneWHD6nEGNz2D7k5hTgZftdxFiuCZe6U
djx1CxOuOJezT6S3BOdu0md3E2yB/CAvmUE4NRV92RBbRL+1anTbQCpMbxJx1Y+8S94JaYLu5Mi5
8Lvlmtz5SKDEIQNNghv93Lxxm3EYGKJxWISw/hMsgIF1SSIQ1ghMIekJI8J6FdzwhVH02zK/sVoE
AxK+cla5MieorhlCzKoo5gZpCXVaJ/E2NFubiZLFfco5tFHlDWP1PW9cndDe/QDe0JFuZmtwO9/G
NkbF8ECpglZ5Y//Rki8WQ3IEc6Ve0M63lXx9Yk4hBIJRmFjXxuUTYVeFf7NvXVqiPdt8WFiEfMqH
b26FWrBh5vAR/SJ1UQX5qEkcqRi5pnTPnCht9zJLk9PGFVspPwHpUXi7jbqP1roM4QnjP7M+zPOk
lm7STI5+zixTZI41NCu+Yv+NkaboB7ld+xi7xQZQ7xGf3nrt/H+Ych542jZxF7B12lJ7mlX6KtM2
VMV2VZOxpRQJjUR6FkqaF7rDRfd4NFgF67fq+6U2f7hOF/YO8QB4hxRXeChG88UeXe69Hb5C1bdJ
aM5IQfBiNeFtPyUqW5r7SfhiWokdfB+AB5lNsni/7OvN8toQKpdAW31hzmdjQE2gWDrKHgOimGh9
HLQCmVrf2G1Qd4q40iLbpR/6aRPm0daXPOAt0I6jD9FO9+mES4ZZ0iT2rAwllf+6UQllsew3yGI7
s0QEq05biJxQr+vEx47IN48VIbLlh2lcYA0mGblmnVPm/U2Vkr2YVPoQbyo0R2Yw49XVqInbqMw1
YAU9rGjhDlddJzDtNElD9ZSelReA2TS4j5qLWi2QJ2/ha+lXn7lNJF8Ovy6GxJMH85FbEKp3GQCk
h/MlAY7s0h3GX3D2hqukMvWEE3Zno9M2JWVSuVZI1xGHAfk0VEcu6FjDldoGGGiXIDxUU6ExdHtl
WTVzr6dBTYNAnGHESVjUzShefHnE0blUKW0whWU/x+njeQBbjUK0PpxsP1Ka7WuKOeZO3YFW1uQq
GW5EwjPTj4WLMVF2aTmoXQgWhZ6QptizNvnzsTsh4WRAqigqSVNIwX47ycOBxpMlespJ0j5eJ3cP
AYsUy5FmvHustK6Yr0eFFi1no+SGdxanvb8DtUQT14fMpQbh4iLEzi0mSiIwcG3WwXq0sxTh3lXS
D/9Od1/QLa8giolyWwPpbfETqf1DXCTNVpZRgzIK4p/tfiNbixGx/es9mwqtLTOMpht0Z6unnhzB
J67N/32dpw9ANCGdWYgEp5JPEgfQqHhpTA224Wqcw+tHZf+0ZlY6462tP1WlpJpt9AiLg+TX83Yk
IbkCHSmiR56vBzHvxyqXnZ1SdeMJED78YV1MdblWW8TgEfDgnMJeKdr6JkPdCaefgpzhae0RoIwz
TgMjwRJxKrWcBLBMKxYVzxQuVIQzOZGOI6jadLLpSNwrm2SEHRWUwYRW7dx5b0UOTNBriwq/MNYx
AM4kXcfRDVErb4pzZTPjipcdQBlYoU8JKe0TbBduEfWlS5pdkJejSDjyOO60lqkml6obCPc093Yg
wLLAQzSLYtCYYGZTeWjHhwd/hBiFt4NX1EjJjuoirz0gSFlVc5xjUDskS7yzO4dXhrIau+C54dc0
AXuOu+nrGt/ytpt81+PAYmgPbojDoM3g06p3d9BFNLovprQ/bu2YXoqLukV9BcsqsJgqyxT2rIZ4
Cm+8L2rhtSOw7DjsB+ZcgAqtfsxjo8HmbtkOCM/EwMVGSkC+SwX6TeLlPo3dY+0Fa46mtz26XDpd
SARLbgwuzCPlxZmIn5VwF7hMzuaF1C+5Kt5/Ywa1IHtahTzOeAs0tGdTdLXoFoNyajd6WuSUA4u0
B2Zi/lts2ZUZd0Ybuw/o67pqHXYjXZPozNMDCdaaMKptsi3ANp+WT/cincY5I8Uls+/VBdgJyHoD
JE818BhWpEDWLVulej4bz8sYKEvMjIFhRaLKk7c74OAULrcH/zO7L+AxU5/5oB7toRKA/LSynHjD
5udQ1GjzhhkA5u47j6PLTBQzfHKXv9ACc7fVKjCoeLARqysZCIAW27qOVArNY4qTK35h4nv2T4Yc
/TuIaxE2n0Kg465no5d8oipJBk/hv/xu7pzpYRNzMgvMzDkuGkmYbXlZexERlcWMQcrcP3LeZouO
HYoxJsboyNbFpRIU5yNHZReDIE5ol7sJzD8fx9pcB4y635Zmf9fyvB2m7guKhZJ/PJC/updoGH2J
oZ+9U89b+u3MJwhJ64exEarv8n7H9KczQGQvPejHsm0SC6DW65TMy7xl+2DfZB1L3a/g23qxUTaS
tT7EV7+m0OG+g1vz9Qjik43A+15oZYnxgY/yieefUVerlwq/KB3BCiVfkbqOlEhn9itbKOiBw3lb
fcWgXmFyh/jkm3NeeZIPpS3okjbwYVJK44QTnKmaGhfTMdXC7ZQgdXrceAj19QABElKJL3NbUmYG
K1GROm7yx/F4ObEfFRba/jJUdE6MQcRkaCd8Xddof+TK3Zn+YduXWr+2+CA0yyiYktWTKjCP/6vW
TQ43R3cMzFKXe+h4Gp6/JL1792r4cgbzqGql0iDWztdwYbntH8FD959HCCK9YYUegkmA9XUOa6N2
BjbwD3isTDJzmQkqLDXMwt9iTIuFga5XWNTVbGiZ2YCW0mhztRRiraEJngHKkTDA0a4gguW7FvxF
8tdCdnArLh4bNSTG3RRiT94HlpKWRvdd64uiFbnwrboL5zGOgo2QU7yDR0QwKss52fMLzfaiZKCh
DPeX5rB4Oz9MEpTxZmYsZKgH+EINw4Vj8lcY+8MkOgQNvNFOwuNh3A9d3BYjQIIhyuBbLxuHzZPS
wX3wHPQAqDA2A4V17kLSqrKv3CKj/h/tntzSANo9ufYvV7m7bFXZjTsMxLTtMAfsQIthB98UDCNz
3R7iJHEIPr+ICNP7uTFuL7pEEobYYY3vXUzOQya8Ll3S00MFJufSAkh3ISokg3TzmBLrb4trHIj0
m6+gOU0lTTLUfOoBj6yU86pyzb4zGPojvIBhun9vwFF5cVxAmNsFnY6l0wFWEccb8kneTrdsRqdP
c26ojznucGx9D0iQDJ5Rey1XYmOOwBbBMpOFcB9InKU2D3Qv0CzOWjdqc/b1001MFsgktvLY9imb
sEIbdOnHyGaY2ljIfG+NEnThX0m/VPYrSOiIH6CtNIWpK4ChwVgdSi2ME7Xtcxise8vISqTqr0J5
qVSxlQVOB+lyht9UKw7pWVBAeVgG0uxhzXDOKuWaIORiH9Vqev+y1/m7XjH4b1Yn9Gt1uKMN7QXS
6UyzVhGxEMp1bL9TkZzVfpdH2XdNNLEMfaadpeaotwPzKxxkvEpoWzgE03hIY16+YCsOkkOsir/0
ko/uL1WPI4AxdQtjjQSjrUJbOU1oaylWiFHlc5HG5bBzua4R6CqBlNmbFFRYeDgBSK3mm9nHpraD
LsNszB+SgiqcdQ8nKp7MWC3VoZU+SNNU+Q6CXYzDNvr32q0EuGbT93o0gz/6dj66L96ah+esR6GY
+bglwc5z96m6dD9bgUCrGA3fpFKnz3PODL4EhWj08KJj6CjG7EvQPKWD81pLYJF+azlZBMGSgOjL
J37/WdIM+tezBzRKGy7xTuwAAtyLlpuqI+LUIBLsI96EfRIAeK2kPT4JcaNbVnkpIItWR+6nR88C
n0XeEGkI11egYEyXl6zxZwbn7RpKSNnuirltweXSs98SWUzrvKsr7N4+rStznFtnY8JzmAifm+Sf
RvawKvI6jGCbgaDnwsfGUljGzJjvP15CqSM58mYGRKO4+tcf+jSOdftXXOchwKmSCgM+roHDrHSL
HuWfZKsqva/TsHVTb1EX2skwqfS+at8OHCOAz+ZY7xe5cpPEBD8NCzVMbldYEi3eidFBE+qjynQJ
aVQkJahQHA0IliiAwpTE0+CTyNlxCKJU7MslG8cKj3TgDla63P6+f+PRD8VKpU36KTATaDs9f5TR
yarM4FQRvIHlE+eanQcq8avGQdKgmJp1JR7WOtYdjklAv8cMsU+TsT4MiLvSe29i1ibjazTTRx+7
OpzgK7NFUOXhMRGxzfMpfA2gFjty6Y118UjYGtVoJxak4kzzwT5n0L/9yBzqAB8VxLjrLAFzhJY1
y6VBkNQSXodmFQkPyequ/OUBeQzmUvVrOEacFbbU9QK3262Slv+gLF7poskeRb7wQVuok+Fdb7HQ
qzhKu6nYEe6+W9b/4gWiIKMGPe7bNcvXXp8N2ulMiHHN84m92XoVpwpgTG8+A6NU+wcBUWxrPum1
x/ISPsX8U/PBGMziicgQ57fU4k8pJ3iJ2M9eFrLJ9Id5Po7kwW3p9hNStdp5OUzgeTuv0SXnDWiS
MxHu2GRl6PDXdfl7W8sAvx1CUjzmcGS4KjgY5trzDJQPXwGE4YJDL5oduNabUUbFdbposUBYagSC
pKywRwqn4Ks23t2vx+8ytaDAALp0tbT0AXwzaVhoaNzSz3TU3mgefVT5IRwQnqNKhV5MoyIqd0Fv
3Ad6S+YZT/OwxjNhKpECZZjAaHtVwc1TuYsJaNKQRhChdM9KgIuYZ3lhNwrYA0MxFmBFJnXgHi7u
l7VtAUMHPHbokPW6KpxhhMbHt7BAB0hkulb2AMbiMxrY48hmuVjqvE3V1QGeDy9k7dhMK5vCq3sx
ezQhMrtCXRLVcwzuKaHvckiNxIVFROjrtyYKxEvgZaBRFHZ2LT3QcC2GbCN9QO36NuCOeQC+nuo3
3NE29deb9qRdkJRIUgGJad/xDb9HbJjaym3wLzyHMRaWMgZB/cOLOhUjZKlEiTrPC4jrr8wumoew
t1aeONNOYN74XnWfR04pLOQC+ChyYKkR1gmv65IwVU9vKmGleVZU8EZSEYrmNPZrnVRNQzoTIRXq
UXuNm+6vgk+9rB8F3pCFDXRA+zAn8kZeSdKVQQTF0FUXkEtMqh5qH3KPDKaTUfML7JAcItbqULnL
9JwR4oXpL3tpCkrjxqy+mt9M4ArQDYIY63n84iIHze11bFjaQ7deEzinWTJFuTjXbOYXyCdmj55p
bQD8PND39xkfK5kskCG1roSd6d4Ol+OnDh6UXeX4sLnI6MJgJasDyev1FLty0NdnFE7JeKAzG1yA
nHhVRjNFQGJvxcvDWa1j9x0UPLPZ1+Eak2CiTYcQ2UoywApulKLE7Wr9yoqPA5lKs2Ilrs1YTdLZ
h8ZBBSBCoYgdSHx7uz2zFaISWQPivxM+TGlmjfX+6BKEEXuGZTGFh/SSkom1u0/4Mi7tFg8n1wcP
+d69pqfVPD+c7lnO4FbKoxh3xdUAG7k3TqHKwhtsY3jLjKqm48049FPG8jpgLx4Zbh0sG1qswBCH
ZACeN1T4D2D6g2yBd8vEJRslLStEz+whsO0yxfuji/0CJp9jCcFruxmyOP/L7gH1he7LsaobHFBW
pc4Zx89P6E7qobO2JSrCN7pq+/uYrehSjDa1Lozy81j947M53EydGY6xKEcHPtxwWQ7CVr9Kc7ni
waLALQv1HGFEiMCNpJkGXSkxCuti5DY91tkIoXbjsGZkleE6kaw6I6E6nI7AV64+98s1J6HKsJLP
VXfcdMrMigQtpzSxfGz1EbywmPT2IvY9LiaYbKluqqVKozKj2Xvkr9C7bPOJGwuJrsr8jyfO0yuJ
ekxwXmpfoTlNImhqfZNb+l8F1Xe1B0QN1NX5SOh++61ylQ+lAln42asfBwTRUGTu75XpI/7fI/t8
ybKMHbNserQjLuaV7JjX7b/CNs3lSmbUiBE2LkBjZtaa7vamr9kW2mWv6Id0EGFVNO7amW6nwfqL
0SActVQCzzbhBeCIkb4+P89bAX22ta/UlWI60tb0Rt59H4ql+95l4MAFF0A49OQuBVoo8fnlyz7I
c7WL2EtfeZCeqIAVVhmZ0XcJ4/kB1kZKtO6qdLe4UB8QRth9rIdGmqUDTb9XjMolvh0Pdhkw+hQD
PVfbX1hhN9wJM4zMBvcUZ4XW9BEPSFnDGhvFfr9LPt/74j0dkysSYP/TZ+lOrLJ58YwKDumeHTl1
U0Tc74CzGVOU392OrRq5hClKvyOQgAg5SdC54KNtQaK+cUnlVnpp2swP1wR5L19j5LypL3T14BAZ
YXP9LAFu0UFg5wLqoRXY9HgP+Isng9Q9zM0xU7Gd7HOb9SDwx58xszwyKAYrzWt4IkpT/Lsad1PD
6becGR5Q/zYlwgUacyvQlHulsZmAqkXJCFXuLbU7VcssjDRw+A3oX7B8JRZtiKlhUaZc8hjUYET6
eb7lbut6s22FynUjS1GqMWKI93l3/nhXSFM8WQkQFAI/cu4W5hBEadeNEDwsGpPh1WbzCzivXdXU
5uMZV/bguTrXaib3JqnsGnMtQEzOB7N/+iuR2SGxf0O3yrAq0P+u3UU4indmivNcWsXaaey7yZZx
jihYAE4y234WHBJQhuu/cceuj5zY5Ju4A8Ifc2C4EZN6BOtWDauUflBGANMMCbHLMx4GCIIV15Fq
/8982ZmpMTfPjuFOO82HLhEeJaDp17Dhvi5iaTs6FA8saT7FagqRfIKWW8u93aSyNwBKt+Pa3C+8
JECPsCSBN752usClkne7jibQ4xxRKzxToKNoCHkuzyQXutf8i0uewKixyII/rgYFRpEM4SCCCXUX
BKnIZ8kFYMmqcdQpdZrWs8DwIaO3rV6d7esXOohszs76D6avY12orZSdXlitDxCfjNsyfGrAyAeu
yXU0yH44Ipp6t5QZf7PTMTfaWOEmiQfMKvsOM321ft59apqE2TUvqsjkmf4eWQErlOTP2yfetWFa
HkY/4kFBaR7qknuTZwD/Wuz0G3SaC+cWuZpR6wA+twHTU35WTA91IFxvGkyFePgULyUWrjdb9ZqH
vwHyNUaU1Pp0pCRvB0fHcgKNVf9Ke8LUH3HeC9ZQbljruLCH8E54HsNbr1XpxupXqj9wEVxV8ja9
W3fIIfN+zfg7uwf0NH6xSlNhIcZeYeAMB2XWVggImwgFluaoeSVTwgdISnNjTokJrFJkpCDDxzlJ
pa3xOKDyHITlCmQ/ZforcXuwiVQSbh0xjGYPAiV42bDMsoryB+0q/SB6RCKOTBz57Xzh4OQEy0o0
M+v9BXuGE5tIu6caxj1TEZ2sgVRaJ1tU0ikLMfyh63pQ1lK3iE4cK85E+n9xlUY96fspneDaDY/+
cest+Md/R3EQtsl9iUEaoSKqV/2ubDyDhhEIhbNRQTRZYzztORWdkGuWcdtAGMdFErpeqIMCfiA3
fSwtU+u4BkeD6RrVV9kaxfXcnSZp5tNI9kBJeIaVX1Qv1YGXaIJMO69Ic86RZ28qXQ6ffkvCtReF
6x7QBwkvtMuoPNg2fec6fwp9SdC+G1CG0qvNQDx9ZmEgw89z3AqZEanQ9VhIGxtQZ1PtnBY0dfqj
koKgBCnhnZ06X0kaK0V/vfoGj5mD2RuRcRa6j3dP8FKAJWV657LQgwzS+c6suuuYMd30wWiBDxE3
LgJAH95liR3abTAhBZGlWrAVTtp6TBaTV5KOWRBjbu9Si9d1SJ/Mx8EXWIakaOoweskGtK1E25NY
AyCMeTdjfL/1HpIBsrwSA060JJfJFzjQMeB1S/GcckstXWAGX8t/swAHjJNO99qSManFR7T3zKwy
v5mgvub2ktl8e+TI2NDyfkCk5FfufEtQA7JqIvBEadj0C1hj7xqxZI+hFrjEWxAV6iEog9iI9Rc2
CL1dPCG/3oz1sKqnoVnCwbo8BZMm3JSUd9jntV+z3Y5e9ObBvNzVpc6TrrAAyVkLjk4vA6X8Aeq9
M270eMYV5xjTstcATiLp7k3i+4go+QTf2KWhmnqWE4F+ZNXIbtAzb7i76b6sawBmcQvds1jKce9O
MvUMxR9M54D7lw5ZDk902sWYtpuroHXuR+fnFwdLA0rJTj7IVze+V3lhO7wIufVyVmm0O1LrLcuJ
nXmt6iFdFlcNuYyI3WqXqIN5M83Z7LwaEYFMcFYNPeWrw8DZBsSjW5/gVULM2C+Ur+M+zL98xnOL
qSW17SICAYww9FJ9Lwe9k3/qm59omGdIYKrtehZpW6UnQZg76x1U4EEftrrW8GmBdu1YjK8YR/UO
uW7hiRXnqPQa21iHtJW+tezPngaeQsuuifYBiQevJkEOkhAq/g4XSZ8DDVd9F5xnozHZZgN//Ybs
KnQ5oc98cCB6KDvxGDNUpccEFxij2bXUspCuNXO9GIDFhJvvOAc8y2Gs9MN2XAi24F+5jwMtKrGh
YUrtTmr4xf8u1DYNFFr+NuoPaBrNxRX5Wiwz9arT2K2mN9YS/5kPmWFY+S+hBXpWSqJuY3O38pl5
/8sUwNxsajmHcbjQquDpCDUSqcDQ8NxHj0GZkgP9B50JKySCaw1+RqjQYFtZKQYOCAWrbW10S6Am
MHezwoVEDUNSX3u0sfrc2rRj8F9nN5wt/FkPJJPyt4IumJEeQ/oUhMGrzJ8H0QB1tLTgf0yL2Dzb
aaInvCCgL0BC1E1+lksfAIPDWsWg8BpMqUd4b8m2KMcFNvtF3MdztTvXTifWCDJTFj8vwtMJwW1/
EK9rZqXX84dXXtBX0Ii927oPdfHltbOkDiZrbw1P+KqPiXinWsDx4Vx9OmbWqjpJxpPKwOttfqt7
ooMuRooYrmgFBOFlk2X+VvHZd58INWzjUYRNxkMBkmskSIqZCTAefFlqiP8l3r9xGqz8AHwMJ2Kb
ibwUoJtanaTjkWwy56a0MAuDeiYJ426WTjkn3v/vrxdwXKjjUJlNzGb5+lUcM9W1Hp7LIIjaA2GV
64Ofdc5GJkWarWKasrufOHj1HIq7T2WAz7O1VOHT17UPR3LkQagjdu+HCCEBmKnIG/ZSBdDTb9iC
r2EFJ+RfLeqdC0djtStZRvMplAwhFNp4HsjaeiU651yk5HeyD0tjOiaF6S7uD8os/T97Ui9hFtno
InIJtJSjTaq8JF+qocT/gM3UqzxCP568Ii1r7Q8Sbtd8CTSuqNYIku6s4oVUGl+aqxvfxZGE4Ut6
9Qham3uOxHktH0V93HNS/KVi8mKtu9c/CQGab7QkaT6ayr7wzXSaGYTmVEA0+utN6l0dny2S5wYb
4mNK4aAwcXdv5F1sZWEI9cQq00h1uoWwBmDxb82zJI6qD7O29UfgAJz/00LnPtYltBVeJQj0gBAB
1aATFVh6AFNGCL9C3z2mH39tpV3Ad47PYVmHjkVH8lLWH9F3UHgnkT9esnhAJBnLgUaRQxVyhQTp
kHHuVmJLAo2R3iuNBiP6moSHBhVvsoFdxONqrnrQpHD7uys5i6TkSwQTVuItEdhooJzSnFHaaEi/
sVnllXbxmzJ8V2Morbet0N+4dly6fqwxRFcCi+0Fd7bgtE22fu6OWi4EI6JH0wMp6zBKd6rqoLM7
WPfcOQ8VG5x2QpOgS2UtdZngDGY2iqPNmNDYO0VUtf2ilOJwXnMwCjTK20J/6uQq3h7jAu10YqIb
JAAEH1+8rcO0llygNoVfcCah6NGHjpB0Hv+AxW1E9cnDWO4mjG7qW24vXSB75ADvEvpDtBrD4ffL
UcqzSCBLMhG2akY4ZksPzgGhUSXGVcVccpSSbLm1puO4VkS0uIdHpEVbYXFy5GSWMXKtF0JMcLkL
VS962+MqccHk/J1vjqvW1nHsz9NmgC3SNJD8FttoZzeRAuc9wkpFzMF82PKfeTW9+xZTMHFLXRai
4gs6x16dAGmmAdp8Y38kYSfP5VKKwt0rfJ5HJ7gUMARH/ZR+GWy0KywiR+Lwge9puESvCCVlCHQp
wrmzlJUCm3UEJZc1XyFebflPat9HvmqPGsqsSWBVhBt6Nmd88nR+0G4JP6km1FZY3bqAlbI2VPZE
Lhf9o4KW4gTGvVRQqqONnqb4AHfhG30bxpkFKy2hz5IgkPprVxxC2w/buh2v6sQVXYifrkkY/6Ig
F4yP4p2VlbZB0Pdhk1X+e+xqlubfWyTWpkY/sdt9sPf1dfsq1K2LNvINT9vqcImUswul60YKbisu
SsYYc8dYeCSRZkkdGhFlDzvXqbPzzPgEV1sQ9+/DzjBkfyC3J6FR2ExtsjKUYy1FSl/l7GIp2zi6
5qP6laRdDxArRDZc7weJ3ssWyVZnzcMvat6iCrqRc1JVlIe4FRambtEBY2mR98c6FynRocAQt0JP
VSNTM0QvED3ekVA2kEy4zH+97mg/LQhRDqJiyR4Xt+rPi9fphH3XjYvLBuxyJj3LwkW/GkiU6CbI
Zc01n4+6AAsasOhIe0zmlGa6H6iUbonluyvYGEJt3pNwARIIcxxYNJNVgQgmXtRsVfsPHWO6iNx6
T7nNJM2hpoQcXM+MW5FX/8pWDMWbLqDMQW9JChyBLQz7Svn1JHW7Hpqj7QO0r/6WZ8uqCaRip/Dl
+MkUHEYCwwDZkoncc4ux3M1R+dMmptBevGdpQUy10adhAkNLplMKgm1xMGAK9pBrjFOwAkGTJoxl
MtNQVlrgammq4AR3gCrJ7yrpLbNYW+qgDCl57eJ9weewHeZdpiMvuRpgZa0YF7b6nM93t9d9tojq
WNvtBdOy55+ImLms7xo5yjsYDwZ0SHqhwVaUerA6mkLeXZcJnNlmPnMi6msrGTGLTSMAuLQRRoNM
fPmNaM51vVmAKzNvjJVXP9erAWgKMP2+rJlMyODB4rZUVy2hM9INW0XVBZdiKoDtphrZYywLikVc
T2FNC8mAePFQnuJidFlECI0HGh2Ko9Ud8CO68ET+M5kkBB3ALwWzUfPcC6OlqCylnWG1BotsCald
WmjJLsUKC3b0cCPYAlOObnhZrvmR9TFF80nomgfyN0gxeSpBz3PC0IMQtMtP0kTmVj1zcjXCW/5m
elrHXm/0D04yJXy+op6bPVDf1Mo/USbDT6La30k7xewFjtfwmqrPRzm0RIPq+UMkctKbiGJJTsiC
KEueAneb0VrhkuvR0YF2CavW3R59LXHMOXJ92gfKmmlRviu8DT0Uza3wXRzSIcXaNlgBPIamXGfw
QnlSBUYFTVzqHJrFQKQOKh+Uv5nXubpBI/jwf8UtLvs8KtdoXPDWNr8CRg2ZWW2BcBokT+K/erUx
Mb5VFLysOlLhlLVdU9zpBg1KPzV0PhKTQrrXwz3WGm3vouHo67E6d/dAiH/ApBA6yVTHS2ycungs
MYUR2JGksF6uJv23cymuQ9CiWE0e4VaAdnFp8EuY+zFTgaZsMtvDTdP0Fbu26dToGuwgpVkkcEL6
mBdFv565f9LJGfWiYSyTtns5pfHseGaSOAQQlEMcvla4W64IMvo7/JRkeCfIHlWFMLFZkZ75e3Nf
3Qmp6TG+lVD+MRmsAJvFjHPwv+vbxGBKnVMdrZ4Iq7m7m9kgYzHtrJwbLyCtq1XmdkFU+/+u3RYa
DtG1KlMpQYphcKcLzLdaYwA6A32NFBSzAz6kc8/+W5+SiKQHWjDzwnJIi+5I1xKgGDVu3Ba5MXC6
Oy2DVZnLrHoehOatAVYdaz7dXGzrHIOEdscGQIkuFyrvQBuLgqlvivszyXaNiA2DdfIGId+NHlv7
F7D12gUf/FlmuChpXlLxcQNieeqbZpqf18k4tGT6iWx/YAsIN8jgiIjbOL54K+l5nGsIGo4XmioE
KunA1CAUPbJVw9eq5aOLu6CPDMpKJEhrtjRz4q4L0UhgVP1XHTIDkiUloITS6gmlCTOJCK7Twx0a
LipIexHXk29gpA4/K1A5z96QuK3Icto8a4VZB5gg0XJo8OOyvom6qRhnsAfCP0nnguuQA9v88Zpt
x+j+/zz7J7eIQRiL/AbPQIpMuRSLC5G5w5DMzYiVgqtH0Yiemt+1IfgmMrTUgJg8kK0gT3ZlgAYa
9iHHJt09apjqh3xBxcRxLUW7PmUANfenHlXqEJQTGcoo+sKoNjSelGNJT7X2/ala3mmWS4JSWw10
ntb8LDntcnCVkaJdbyMTyVAjJQviia8AWQID53ZiAMB89pNe67PS264fIhHhBAczGVRmily2pE/t
gEeg70V8W+MVfs9WKuc605Fk1femQBds00yzgfzsXQVjhw3NMBNmQGES/AOPYPLbU6l9iKvdlXbC
ofMNyt9b5Hbczw9Bosle3Tunm/EclqO//vEmfwPDjI5fKcesVwrtpEuxqmnT5ESrY+Pmg7g8sYPj
d1grWQRnwLBzCeCs6fbP/Br4gd5U35pmZs/trU7Mys3YSS709HZ7cGe8DW9gZvzId1LlJ8WXMKP7
qYHPfuGkQPhqylAowZYSvGkZagXRI8DGLC4p4StOHq4F4oP4x8nV8WaT2J1M2Fo1/5VCQX+YaXCF
7Mg16+wuKSrjbT5/DfPeq8Tgd+qfoP8mSVDMOnBMqmsZVRsBiVfdbACdMhoPR00tp7q1+05ESh9o
LAQZQe22r7kNCCNf9KW8S1bgY7MqFBlcXG9Gclwhh/TgdOluRnTjUWeoyFTHgHld9DRhE2rmam+g
kZmmxZOQETp9wHVQgEFC67m4krFyf8Oep6PnYIyBX1cyNFa1OUPKNLoOrMs5qt6YSJ3lQooM5n+3
ZJqoj/vw6hsCuGvD/fJRzjkMlQu4oLrIyOOjXC7qaGbIJZGFjjhNBq7mzBRJ/JCtHSSj/Tps53ii
P6f/z7Og2kukkos6kU5PiYYSzCmcvf5jsBnhjNLtVkdte1hS2b6nVxawr4eQdoCLnCPjaO+aBbqf
QdIbxafmKn7q/k23Arwocd7vuag7hIBEd4QoNoW06yDilZRjC615ZE74Y5yY0vGDjmqJRrrC/fOi
iBZk+hK30Swf3eJbX4pBNkPvPNZ87Ey7g+4yU98OLAGh1FnbQcYMWYT+cCv40FT6HT4CrcUVI5wj
jmcGyH8EwC1Bd4BgqU4lk3TOZR+1Fen+Q7edc0Y673DQAzdxaWYemHXwYf/4a8KGGB9sK7fvwo31
CET9sUgYgrIuOC8EZ9uZhB0HvIeGw7H0KJXphkkSkAR1FoRhvAlDMNOdnSTzHTYtIS0EM95Z3ANp
3E/2B4mr9zGTIEo4KRUYylF8vLTRIMmd9N6YOVHoqfL6vs4VA/MQNiMuzszEsJQ8tNPkl3Uja6Sg
jZBDnQc3v3MJ/HfT03tK5kN2FCJ3Kkv0b9CurwvNYX/EKqx2lySRs8keeSqr5HKUXYjocqozMKOJ
Ly4tZzooJ810zfcCjCG6jh/qpVamzxqUHyOfyV+bysWlmoVTE30zC52h1rA4FMRqBemJux3mEqmC
Xo11sFTt8AHbS7hxb+P6a4+llyOJhPu6k6Rx4KoATpYeYy8eoxjzQfvG9/LFJ4Qmcd54tpQyDyvO
I50Esvww0MyTDem/k+biUJix6zLgfXAPnfPZsNR+7sSMVpR7CLrqt/k1/wXU4jEBBC7RgIsKV0gu
cAY3pwrAau5CXBNzlBIWlgByQxG2yLlws9usrC8etUatIjMZMrWV7VdztKm0AEnUG0KYycUv7qyA
Y7Pv+ChXVFl3YTmvym703FJPHvJp9soBNJWRA/qBVUAtZduwOvLjXoZemWdmCmBXe2Z1BknmiDYG
pAUgvvyAKmhIbMHf/8M9HPNEyjvnTXuByL7xUVpTDbQdHJqO4qjCoRnUj5PrisCfFyqgZ9Z3RMG6
oO4xuZD2IcgMdvLsaCEnPRt25aiyxVepz1pQ/0HA+7TxAfeMTdqz7TJ5eaSV6N31mvv7yAPbH1/D
t6YxlVlv63D9hy/qRisSU9WCN46djb1GLRJC83GUm9uHj4RPy6bGhQbbgl6qoAeY194p1g8Pl9Cs
EFEoIxRkeJT5aT+iSiYl/Q67w09/Wn/sKtR5Zo9w+XUlKCc15kDWe3/LkaCPGlP0cwyVoBPIH66j
SaL8BIHS+Kub3p0NJvPiY3Ek8Jx0S2JWoxdeGP/hoFbf/8PTN5D5QsoxPUQKQxyz11cB+KzDZ2YU
xa2boD2M/oS19WgtUlX5PMBaXsi18eX1uZ3shEpdzA0BP0/2OAB7o5t8AKGDsl2ZhbOQlUSw5eYS
toWnenNqJJz9kYoJaa0TyvzLNkq55UAsiFilq6uJo38RBB7pY7igfo6b0U//ggMXhMoetYcClJom
uV19QuonJFa68ga+cJcEkZ+nslCLtv3/PQgrwhK/tss6qvaJFLhp53rRNMOkYqHm6hnxtDZPI8cU
7AUyiI+iZ7klvE+zJJFlclXzJH6ZEzGWIKOvxqo4Fe36wWuFBFUziWcFXSLa9RtAXCZQnyZWHmwN
vWLcp7a0zWwSDU++ojcNk2QKqNVYKD3xnj6ww0IDdMa+pneQJCB8A7LjoFdMk5Q2HFnVW0mD1zn8
4PPZxIS1L38aYqMCcOM42xFdn/TVmt0Z6sstWEyUbz8nSzzZo9fOboqNBL5CCWLXJaVZ1Ez34AeD
aOI53FR18YwoDffocoENmtFMfnrDnbxTu69aYjSHeiI19gZFxW3unvvQCP76y8ynxGlvZzl1FJEL
chpyHEr7O/diLjKuvea1pRblrGn5v7q8paWBfJ4qR6V4PFdwVFB0vVjihXafPWIwQpabDJS9R5/J
GiKzsT2MWuo6N1Ucs8wT0TEim4UjspT7JkI+2xRA5Bh06BrPo8kz72CHJkhoG9IWbL2dvqV82W5/
L87Mr/ySmouPilaZyw+ioCXRgnqapGUwCG8eG7aTGdAt0FF6FxbaYhA9qe3wkiAD1Vp06AfnwcBu
rXCNgotAZAE8I9lo7xXOE2t2NIB/elFtU+DXHHXj+hukjFcCFB7O1LLuVFfis4Ulum7C4rx3Lg50
yeVhKH1j0ut9k1XOtF5CbJfLfHeiVZxbCMVNm7fIfAaJtll35rZq3ci+jH1EVzECSofnhMRevC+Z
4FTKxCMKr1sXqPGF1z0wt/84jl8NUjD8vx0iyYk35ri4fiO4L+15OO+PKYfQyhdXSvcypVoGJ3VP
NuwrCm3ypNkdu87tgn/IFEMasVj4G+wuvQzPH+m5ozmkwxG6mop/vnog5OLoQeZk1RbZbwp2XC/V
V/HtRTXfTRdmxSLXioCb/nGFY9EPGFAlkWSGOT23+rPMuIS/S2X2qGJ2UK7s4Q6owvUQfI7xxxhl
6bRcNmehxCrCG6HQ8P2XXLU/eN/O0s0+81RP7jlzNzMWnRiEl1Pv4MHvpFX7Zqo1AwaBisiJaOmO
kU+IBzgdHZq+iw2/6TUQ9Jne4GYP3pI8Du5QVu0Ry8o4Nj/LYS/8HrKBGCqjjP3RNGOMIroZc3hl
egJQ3Zz9pgIYKUoa8MPhBvOcXzpBYJowuj/DJQoHsNsdKLJAg2KT0bpYbXbZjWZ6hkINBDnRwtVK
qSBZgJIEXqN5MXz3/7aabbDsFa728xszaKU8+cgRijttXE85M27IiLRGx7iJz3NsvORMa9qDRY+C
6SgiV2YG6d4WkJHGX5R1ECFfIyJEY7+qWRfIwHu3FILrMpq4gemEENNaUVmI0fwQa1Kz73/5daS2
k7kJB3Jxo2DSWCBNzKZNutkQylEfDsGOnV+syCTRuVfgeLDQdM4cwJDEaaLRNky5LLn5qu/zCOlE
gorDm1Lfaj/3b2dUQEkfCmijO2Uusgp85fLYNADMAYhtMOwUxhGdZITMhqJVbjpbRl1KNWAbUjd8
IoZw92wGLbLfkF545qYCHPwjxE2SDtRo9Xjmjyv6mibU6XuJfeT/LNz2P4RiEbq70vWumb5UVkCN
QFRagOFY7VXB+Del8Zl+rXWRTf4NzmCQ12FGSz6qGeSsPUJJkwXqhkKxaUcbP/znVt6pV85Ybex9
L7PeoE4lzCleiD0P5zFKPi0KNy1G+3/Y3FMXekLpa7a1gooSb/KjBtJFeuqGXLSVrCNrytU1fYKU
lVetC/yBJUJovB4r+nWkcXCpERlcfyfREpPyry+FpVbJLL2oLQ52ruI76oovIsVxb7zry9buoqeD
DUOoBX2NHRBXX77Dm3d83v6y7zQZYBgpz+iqR+4Ra5WQSGA6BeAgTOwCaHmhwd/FlbD8Z0yL53AD
Xto25zVrInn9VjP/6QJt1BoxmjqSZA+LQ0VrZnzxxmV/lsMgWv1GSsFw7SdTEoAlDFkHoo1fjCjm
nWUFvDEhV9p+J1z9jcYCyAqtPoeq+n/DO9SUzM4fS672chw0RrZe12uZq0+fSwx155n2E2ZBsEn0
gZT2mTiwUFzK+epaImPhXVbqeAmd9KQ1B4zXo+WhDnDzDeB0jEUh3Y8fb0gi9fyhQlauUC/fCpaL
k5v8SJDYSFX7ref4+lf7SBmXKSU4oDicTTQt2qIAS1GwSJrBlHLyxIRMCSuuHQTLxCV+zsa4NXWe
t9s4CEmr4oRFXwq0Tlna3F5NLVZtB84ieF2xFUaG+rbFoFobeBVz7vjxOw2OnQJXkzOz21PjiX1s
gwirw9DnrAuiA1i2mTygG4mryd3+1+xziPJLaifuW0s5oj52Mjbg0IEAiAhbeGANiWrXEomJkfo8
WtplXEY18x/jAeXLvPruX6R07oajtT7iDTd3X6taWoQ11w2coHmAuFrqtOXCKhf0sJZkT6GfnR4k
aeYgDFi5XHQulVe0zK54uMMK6c4EmRfnpAYYWlUThoGDKowTIoanMTYSCpbcbTVIqmJKv7zl5/eA
9cfgSUKkQYZa3HVPjkg2cFf6ahsGmIXytorWboFh7NvPQZmeY83/e57qdd0dXw1MkS1NDSxOXr3V
kTlOzg7tTnqTPlltZC+pvLs+rnNs+ok4hCfeHbUgF5rjnhuN7/1y9nauyhb5Sr0+n3kSjdv895SR
L/p7yTsFZXxP25eyrmrpE/laKXf76s2fm5LDtG62lfumx8Uz+XVZ5uAc82aNwnvGiMy1ODkOEviO
disHe+Xxmzr88Qbj3nG7wcGd/HRU8mxu8muU9jECjWQTbHpU3d4PAaOzwfK5ObGsYzuEDW5xVCtO
YeqCfXDUsxlIyUjx0Q4HLNCQ9JcUFEArVIsLK4n+guKYZBCqrcIFthXZHp0QIkwxkNkYrLG0kup6
0btesxvAweoWoSsI54lDa+qinjDZysGyOdFkf69SXaRncSs2drJuF33QYBzak7gtNkQZmrwcgZPF
y9LwmkFscNtke07QBjCT7yhgiW+KTc2wQccXgE0+BXbmuvF7zFUktQR9Z1WlVB1cPE8G6y7h6zfE
TkSwf+UMHy11ioSVmLVq9t1ge10WdfuJiouh0GywjIPvSvseUMpGPaToERa+HDYu0cLi8kUJ6N9t
K/cbX7i94IZZibK5+sHQjet+Hq00sAbatJfSH9gZroo1FahSV2Av7pOBGcpaZhSM6h08LdmDprWh
4e1HZITzlmFWItntR2Oy2z9KL1Hfq99v+EvVABgQ3O23GLlTn4GartXzf3HIyL9PBkBEAC0icXIi
qiTG2XI7dOOkeWVc12qdglEuMyIShzt5wPpdf2ArkFdGzKssaXHYaJzxBAcyUwKSTT8swGt6t/1N
xeu3c1y5rNnA7EGEFxRT1OQkisqH5qFX77teUqc1p7RtZTNtoujZ2biWCbqCtKz84QLsA3smTvVu
hFT0HvGQo3TXY/iIOwLsyzNTTRLxKv/pui9eo5uunInRFdEAUhgjDC7gqjnOWVGL/wzN6BBFCoND
JMZLuKwAmXIgEaDYHFJflCdLNMz192fOqO78zbBlo6v+2A1+Wvf13UkT1R1Ji4q8t/u9uPPaesgD
3dyER0lUfF1GjSiL91pP97CubVjekAJvckRd6Wz+LlSjM6me1a45Jkf1h8kf9ps/4CtlUXQMgfbe
1KZKql1EXsTLoopjsCI0GvNUFQp55AZMURPDeCOzPOzvLUu91eZJ2hZMBbLcEuHP7xxtAI+6UYPe
LaRDefBYuqXMJCy6uOfWEiOre7YhXrHx6L5uDUz7rNMzeiIJaUuSA7juNNQ6m1kmFwE7z4v/9Kjb
Sp/4YXakNd3dnlMVTmuvemeILThUaU6uSpfI2px2qjOqM+bJ+DUQnCc6IfDWpgGnT0jvXWJxMKhc
SIDFRjPhgYZgvP1ItWxWLVChiTP/rk/aL4D9QbR1UxiN5q+GgBUgE9WA6UxV6mG0sHOEe/lb9zJ0
Pfb/zaB4itExADw4zLaY9g0/cJk2MIRG/PTlsAr0pU0BNy4NGIiqOX0Nz+5VUVGjlY96Dlw7s1NF
bFUOHluX8Gpqowt2DQRgt449Ja+WRW0t3J4Q6+5Wnt0KDP0UrtlGQcXGt2s21wLPFEPJE4UZ8JBI
g1/pi691R5UzgYQZa9SfPPbEO8adv+gDvz6QQbmwMeJG+gt1HTB0Qxacz2uZpSBz8RmwXUyccAHg
BGGewOiRuyvN7SP9Useu7Nufxe/MhltQdlVd0ExgPXWvWEYVZ264XvdpMmwxk6X3GLvBO3EBXW0T
XMetCyxH7zMMKlRs/j3raVLLGwBC1C1K74jjd3ZKt/5BhYP19AzzIir16TGhZycSuP/e45g6ZGoJ
uSXaq/UUAcgPwyk4FauvuFAQgIwSvPykCMQHp19aGGSrqrWrCg9mNYsUrk8LkUtQ+ZUdXMdW8Mf6
dtWsBt42t1W5uxQTjQJnnc8kl6x7L6w28EogXEbvoAiGPxB9HsuvufLCHsoKzRsv490a3OLMMFqT
gnLRF7jZE2FcA1GAoAg71cmsM1OTNhJoiZVhgDqAGfDOZ0+LiQFQC7E/GbSjX0vUXPTDWhRNXzgo
XYkCoBb44/dip10Eq1P56eJckmCdNScRbAWHLBMjfaRDDVXMULbeGMeIOwJ1Cl9TsfuYldb1qmj4
7Ai93Mmv7EkPr3cecVcuPfzYAYri72t33AYX6ckJ7XaC506Z12mdG8kH2cUC39UG6N5WGyvn4oXX
bFCQBBv3lONq5kA3UAVIPfdZjdSQZiUdMsRN7TYQizydwkvmzrwIWX/qkDCaf9gsxDXz7fWWZleN
752cyUSTlpEBG8UizfAdfrc5dkLynvfUGMvNSDyY80TD9KuZfMRu57juSsADcseE+jnfRWiP4LPv
0IEC04lU7pmz/X5PjSt3mavNPO+vjTFi7A2gy1fc+E8gepxbOKcxK/XTcccQlSGb589K4RoJfdza
TVPodr7M8uvthPQU5uN24VcfKdFjbnss0vZ+u3Zn1nqyaOLDkEzlVxOy1nNJOdv60uY8M5r9ZAN4
jF9FUn41sjZqhgAA/uFWaokJ8yTuFdD5qKFhZBdy7EM0LeNh4pDprxlXbO8uET73Wojn0/ilvOVj
QDEpITzMkkwPp0MVFYnYFKdTdgtffHWm16ulpefX7NG23yeExdTaIPTQ7RllTMBNm6UfWBAks+Zp
pnXg1m80mx/25jhQxNg6E53qFkGWjcKPBzo26gIbATpJgHZXVe7ZZIZpTCGNKJkjil0wqPHKsK27
sptjYIWB4fD2ZAQjjTEX3kbfC1CpyMhVgZYnQWV7HgQBY/cGFj3cI5sCVLED0RyvfLeDKTH+/s1q
ycHR/5hjhNLWEkic0gE/IcJC3aDOJllH0lCiAY3mWs/Ijk9YOhYetFgA2+5d1Mxgeyx9YLzcgtYm
Hm4l9+eaN2XmEppXF3alw4Sh77albTiLL0AC7byjrt2RZNebPo578C5I2zF4XGDoLacR0ui8pLqp
ugasjMMCEcnlG6S3MRvvpYd3aNV3dp9KHpJ92tuTnKn5GM7oVdl85PLIULFXt2WHS0ceZqqlGxGR
vC6z6FYyUVj5/sfvVWKsmkKh1C3Lkm8GE0o81GOKj5YjYM1/nnfdmd3BUdEoAHDQxV3pcsQ3XcGs
sw8I08ANe+dBiem0j+omsdGCWN8dkoZomyHQWRHveKSPAQGpjByue8zyitFiJLaDT3paE2bvGzDh
JGIRO9OHJikzNlfuGauzgkQO+f5fjJ71fmSwmEGYPMTfCnIMhJQYY032J1Fw/S/d63daHqcy0ZEp
eAV/LB9v/4BxNET+sZ2/+JR0lqhIwgQyF6Vee8s8EUrbbNBnZc2U0/irxkkuEJslUoxIGhaJghur
35ieId3JxcvMQfSxDC4sWrzXGEYvNslVuAXWGX55t8xzLwJuX6jStGigbia7zqJweTBmaIPCyqFK
cAjkzQzSkY/cvnutD+v0QXLcuASvcQkAA82pYAq47EdEs8QwQYpCLkCz7BdZO9MZJNcAHDkUYjPg
iT+5ElS3RCjuuhGXBQFNnk4RfHmESyU6afxMi42gNlDVqa5zfNj3AIJCuGnRw/2hGdlyd6zKrNjF
S0a+nIplgTDRilyNDO0wX6o+s9oqYTBQYWRClNXEHHAdKn+FbLEKONrU6JLrSHo8ytiZqg45ve94
Zs3XyNIiFsNTdzuxgPPp7hkapDmo1ZUwpXP5ZfBECdwnFnJlazvSKrImbx8QfbVuZTui4HjnIrQc
egSi9m6spla5PbCbXRI7MxqYQ3ETwiyZy2hq10z6BKUg4SCrHAezCk3Cbj3Y0If5mGPvAnnZewpC
X0eS7gDIg/FkzrfIUn4vNYT0yfhkEqy+72J4M5twkFlB3JHCgQdQDnp8I2JLXH/5l2yY9LFJLmo8
9wdJOIAnG4SeoP1o+W/FeEkSGn4FJA35Nv2z+y8kRDlySsR4XUYbP3gOWT8jm1UUSSi4E/KZ3CJF
ssWw8ZllJasisQh0I85iwFuVl2PclMJ7NWVxvGZuc/s2LcdjDUTdUP/W6wrIHSfvQByMwwuE3nvL
HEK6Uqsa1f58TVuQYTnNnq5k23lr1LeF89zjh9ScRl8NfHTYTbj1PLsq5u8ciYyeTDCHDIJ6vaHs
G8T4FSwTXzzBROLXey8NY1+eK3yLDhMlBFYz0i9xiFBOh/A3SvK8hm9sga5lU1o6d6GaA6zmwY0A
Jzc2Jh7pQtuUnievxdCyACPw+QwFgxjk6yRVHCgjUFY4mGwPkCavRMW3Anef0MQaUBacoO3IhRZC
RdgK81t7pSxRRF4Ue/A5frMxrWF1pz6KecOwcO1SVr7YB91Yfz9mi6XTdQEvYVzUXOmPdCrDHzpX
C06VeG8albLmLagnSiLPFAgCkqfByY60ijdEtFpeDyYF/WNJTsyHMT5kRDS/ZLJstJzcMkkM9GYp
ahrkTXSjZxZWc8n6uv+LZ2anx9QtgeBgB2+vnf3XciqRfIvRfyVsShGxNdywSn/YofRLMmmJNe4K
q5uI/V7DMfAsXoGturbvRwBWLCAdfWfkG3TdYAuP7ansn0cw2TowRzmiq4jVrYf65mwx2A62YNuq
ldYps7aS1GK9+xiF3UyWehOWS8gQHDOZm49a3bMcYwC11ceLeyDDutUubUlELnBKHvMcL0osa4pr
LA4rMpdwvmfoWuY43h5vyeSWfzaCTkL77NUPaGduBrrmIm6x42ak9weWXdxOSHH6fadH8nSeNcku
IUF7gbfqAsUCu+kKRucNLh1OTrWNaRdruoia1al4iS+SoBSSzT8rRePcL0Gmf7ueDjvUke61puKE
uV7cfI5HuVDLe5dSi1TQPhwlr4c4h3MemCHArsjlltKa8rE/LrG6X0w26wzRz2WSfbbG7vSJcwd4
iraDKxGatJsyrG7vhno0KUe9oCK5LgUjMC+j4Jw6byxN1TWerKXnuGLOqmZC+viUzDAbbBbbp/or
nXz677i9d/lCQXy98CjRfKlLvqmT1sHMGK16n8CcojwUyrqx4urdC7Qmy083aKGc2PUEUSbX6igC
ArViNdQhGOiumm+IZs2D1uAhclkKhYVNpSCMq8KUNSgx36Kkx7lPu/2+6vCheMRPF94kf9qcds74
VyqWekwX40K72JlKxROgXOmivgXmfR7cq96nCX5e/NEO06HzblD3BmqfFQY7ODMizPyQtRGgb/4p
YjTQ9B3ZJ+iZfdfYieSTqJNqAZmM83FBgwmlartUvcufbEGT6LAsnwhGGbm4SFlYKC8GVw3e/QoP
xeRwb9qcQuk2xoAZLJoSnUHSgtP4vvwN1v8ZgXiGfuFI7lUgLYYmft5VD7IAn7Aq/zYKF4V2c98A
eeITV1Q7i92g5YRmXG2dyEOG3d1ua/XFuIHjs330UnOrJTJUbLR+uprSVMniMtKC/jaDUr1eG7m4
wvKtR/G9WbqXSI3rOIn4j09jE5bTOT5gRnAkaPdYa/cG22MfFxo2ixTwkW61UbwVJ9K2S38hnfdp
fRJ/7nyDVOziSCah71AwVN1hKcPyD0zM2QyLo54/7QNo/HtLKcjzg0cfYb0yBPADdTPqCn7Mcabs
TRP3ESgh/pR9YlQjjHlxRYUOJHv/V4/b7eTvp52azvGMR/UoLom1iu+6EarTcPFQaGx8JhLZJZyA
FWvUdSl125DpLIZnXe/mow/d0nfkH4XUpLp4kZk+eaPzcKtwo/SleNjE5IxjO33ycatYcbHnxXPV
etbU203eyzDa8xMieQZSgYB9vKuEzjSOtE4KE5Zcgy4+e+64jMm9k6/q+giqzvOdX48B6LJUrqQd
e6ukOYBH6VYy5SEZD43rlLj03PxHG+30926oNYR7jCiIk+M1afIWCjZ7w/diJinwYsz5cFeu+Tzy
hzTDL8D1SCjtlorhdZxPGtWlk3uAIM6JFc2kHu154fUcINxW73yZfCl57penvJCvLWo7xZVQ3rqU
4DCZd2/eHC9L21f28nMmOpnHqw07qX0ZFMv/jedkcEx+0qqKO1mr/kKuuRq8tccn992YesWWV+cM
QVi2ayyapyfzsRVQVMNV+ubteOU6NMc3pm5H9gOu6icgD8K/N2uelw/b5A9OhqOdA47V85NGJA4K
ozTd721bjdL4FloS/VMXLbc+8DEc/HKeSC+e4o+OwwPbhOaE7qDoNltUSgmNrMthcDN1psm6j0Mf
+Mvc4X5QtFWJp5TVZbLk81Uedb93GBeo9nkW4qeexWIWj0R+I2sfC/TgFDkupJwTH42vDpjkznVx
J8QwJ6cp7ZyGESlyG/gppkcIm8LyAmhrMbme8odaI6Eve0zv3PqDLMfHcA3wa/CS9zY2rznAh3Sv
SPubbQBshJidveu1F8bNV9JyaYmDKV1JGwmZkYtPq0anejmbHllZHoLvEytv2X7Sh/YoKOEmmFon
bVi3ON944wopLPS09Lxq5vJ/ubJCj8wZEBS/X0WPo+2EqkrU5hwXi6BoYmyAj2rFGbeUD3s6CGW1
JqcdcejnIyw+TT1UWla9M7pFAvE2+BnLthsM0eCvoAJrGILUyFH804v5tc6HmqX+4TEXWzy0nzu7
9fzttMuLDD98IzVN0G/DrCp7RM03KUA15D3q/4L911xiXq5ojRI0IjLvM8eI7xWpz1qFCYg4sVpd
aHx1LYddujYqgiik2ZJqsh1YXVya3jUWvACuEDHEt/uu7bUFddwGyEFKqdvgxizc54atTyKK3q5T
zT1Ud+Hd6zztqBrhRsPZcFj8J7oGSZMl5vii820kpK00aU1kty75TaMth0kSVMnygOshwM/opnc2
R6gbCZftKA6P2UurzmZyq/eMSUl0IlsUSUQw20mcrxmZ7Foo4qEOy+VViff0GvhUAD8Yr7f5coba
AuxuadmsHv84wAMn9HL98czcGpBtbRE6tH0P9JsZQZg/3BX+jpyLSukyXUzyZQVF/XcamOiRKym6
lJ8z11K7P31vn2x+RL6fFS8NG5wiSkk3WzB+q07mpS/D0SjgP9bwawDSPmdDqN2knwRSD+G+9AMQ
C3C3j5aGLhfm0rWY54ZEVGReKSCgx8Cwxy5m/Tvuo8iXCpjbJXwIEd0eep1boh8B1Gu5toxHvqmc
JBqK8XFYz5heeQX5zcDTXq0SoWw/e1poFaY8xsef9dRiqzo8LKYhr8VmrPSqNU+XCSULR+e19HeJ
Ayc4wNvDgh7L3Jfi3cs7DfWLIFV0tA63ti4G+ZrczjcThSJUMzEzStFygpd3fYY9T4XFVfjXGR1p
7nz6Gv3lU/YhtJFTvMG4SioR40Kgj7GGMGm45eosk6KicfRNvIIIDnhKAyLT5alR5ZUM2vc9B7Uv
hHZtk4VslXuuvJtE2gdK6i6oiS5U95H0sA3omQQfqeDPLcPdVvVmZPCb/D31COVjefoArAbkGaJV
uMoThcdtRozTqfsTtvymMyUdI6cHtbTHEesvbiIS4oyEaCKZ46PjFRG7mUZljo+ORpoaqtXTD05O
i1h3LYS/KeQKUuEKa5jRfyfKhC5eo3n9NbELGwKjooxbETGf2KDIHFQ1YsmTAEd3ayGtBLyzp6hS
ekOIMwpgdSlibwppb6L7R0F586CpkpBV/4UKWy/oHIC9SnYDT9nNaiO6if+6DiP18S/D7riAuCie
E9oiLWRmEwUTbuY34LhTnMQT6ZmbgirB6J7mHbCUSXGC95mehn+X3x+f9dqTzDGuz+0SVaBIJtp6
9eCrOTGx17c5Pj83+mffnetW+mCw28lLAOkRonlfx7qu610RO9Q7LWw+sV08/Dnp0g+5wtQZ3y25
65Iid6SVKJE+gQ2Qe5hc6yh4YW47rgiCbT2WLX55MeCUcGOgvhi8ZrR+8SwFr9xsb5alv0KQq969
O7cZYojKYvEuwdTgpN3WhVrsOxETcPP9A49+F6np+fX6dl53RKeKawk301C/5djR/UvGa9EMjy1K
uhaeDNNdKf8YQn4FrjMbf1tDMyTVmQV4Mibp6P2NM7R7G89VM+lOpeiN8lt9ddp9lAyikmWtQRq8
a4Q58eJr5nakGCTqAFkXZKcN/QMddFVeIuDpth3fBeIVaoxjw+0n6SpfUt2YvSgKorjljVwA5Kkz
lTSPqIWljxP8VUnVpzuaRy5xQms9E0i3CEtMPj9koJXcWQ4MfsJneqBOg262Af2sr4hqnfUtZtNL
uSoLtHzBHHeIwgi4CCJZuDLy0GfvuoCeUKuI+kTXe19Z3oPndJK8dvlDY6CIbh5EStFTkScPuCLM
ovtKqEaArcoipLs5bvZs4Aw5qtBmLClUN6fL85+zfJoXJJjfswed7v84taXS2+cefAgeBhl0wW7Q
u+gfb87QZeym2hKgxOl9fUn30nxPDSF+koyxx1OzXMLWYzHn3eDUr0yUKG0SeNJTCa1ZYTBKt7T2
uGzbisqDbiRZAfRwOUf0+oUINoTFo6ycTRNkeTOE5AT7xOyaxWfQcOCWkLU2g+p6oPdzylyKNLGW
6sDW6FoMoTVfB5Fy+MssYAMbZpgfS6qR9bWUBIXAP5rUvj+yWGhtegYwYj8duYiNG3sxKEs1Z5Mm
WIolgRAysALaNKNHtn/vkdN//XEn+H0sTOOj17qctDGK2HaAjfoVtmZf6Ry+k1OqPDffsLtvEY9n
eTzSJ7Wwis6A+lJEL/hUXAPs7Z+9mPXZtDY4iIc3+eLwzHO7r1Ra/xHoOfy/9v/NvSONvaTRV5DV
QOGdBGwrJgjMctooZ57C32VZCKKKb4XzbAXeQN5IT0Vq/mDn8w4SuJQzad3QTcmRLGTKGS8flRJb
SCmpK+o5x7Yn3VLLT+lmjMrALPxere4MMbevwgiz3U58+4c6SW4A3wRAi9+6mwzn2i7t0ggYfS/h
kSQSig6gTHHTDLmu4xue99HduLLg5ktc8ZP+pWF48qTBEyqreauXFa5fLAlf3KgD47qjFtbwCQdf
TaO7hVbPogtvd2RnWAJdzAS+BhzJfgqiJieUMLQUvIVE8w2di8uwkyqHFy0zHYfVgTYMF62JD7/w
dnpYtlm3pBG8NhWhXwCTuPtrvbcZEH9UTWh2JCENalQ+0UphoHvpMt0J3iQZ7rXvrvqVcjoQyszm
FJknKkZxCgK/sagHJeleJCISANklVt9+uqW7ZkCqOFxjnq0lMpgL+V5kKAnESi/9z2EbYo5kCQ39
xp1aP+i6f+3nHOREJkc9yhJ4PDTfJ+PVzcBdhF9vTlZcs/fxS7eUvPhxGjDZQV8dWJGHK/8i+9cS
A6wKC45u9xH3jFnOBgayl35vq3SGXS2fH/n1m3AuiCe/TY4Di50ITf8UZVd2KWKPNSnYErhkIAem
3L9yahC34zurVfTdW7wfHeWfLBhbscbrJh/qOUQmkp+YVs7c/UTi7e91LjvSh8Zha7K9Z95SiEnK
6+QeOnk6LqbGevRwW8u6QWLEfbfBDS9UFVRh9NabnlEXCfNGkHWSIX3Kt9Hi2+4arUT3ymf0svMZ
bAAkkcRzBn6OtUg2DdRDd81koPLEmy4YP7THqzn1IPgt7Iyb714jrJmyAHXYREF0GMknd+9ifqqj
H3eK6hliO7XSFM43VzCPKhz+VJQMdROSxa4nN1xLWQDLP+E/+BkEcPNl/GvkZtAlrYjOyRVEJkbF
aeohey6CZ5BNTlpfsz2gOJIX2p+QBQG346Ot6F5N3jkqExi6onBx1wBkQeGfWGpTnfDiO0LOc+V8
5+mrKPdWnOilWI73jXl9BLJbM+bJU+7qtzkdPsYZyT69//BC7oClro4Xi3YzNbabsYQTNuJiduMO
WZLwiK3PupnIG5IA/ps8p0NWkw/uBid+ToAUb9/0Tl/c5K6UsA/tgu0uRMCfWypeMaT8O2nHRr94
u6j14uLULFTTCmhLk7aU8Pij+uv5EruZHOn0RkTyWxwNwWt7/XHZa5oLIka6iYMuB1R4Ky38uM02
4ABlbQPcOV6aiqolxitPrUk+QCYOYpnBUNRvcJds668d9ojRkJuWrnaL7ks1CMr3PgX0mpkyxV63
zv7tOqbPzZYzvStp3F+Q8P6gRm1INAefZiJhdfgZaJ+wySWj1wJCDWsw6HF7qCbrOGUtuDol271g
PrMSAXynDkyTD2VhtjpORjU9+Q1kXcRFyekvEm9b6SjNuplcTjFwi2WkW4eJGKHyxOJeoodv5Voz
a13SOInd/7PjcMK60m4di4uymm70FoGnbdPBLFWfZQnbgZ57Fmb0i7cELk5/1IS6zMtLl6fH0sAK
D1e96qtPsfFdp8pQJ8gDeK7T+owezToJJJ5VaO93x4Qlujv4C5AXGG9bHaM0IVsSw+rB05Yi8bps
QYUKJH/aWhBEszPBS5aya+imEdx8V6p6dhpI0gFSbiGQwsJ/dQT5SiVL1UYtVIteHcqKuNx6VKrj
rqCgAMQIPswqP5/mytEk7Mp/lSOwzxUhOUqhTNWsYT5CRRsMZZz96slDZwzbj2ElCuL5TO7Tajcs
Hmwr0WF+VCVp/bownz88YDGDzCEUX0d6lHVHez1YQoiWgRQVtCMufna9nJICE/t1+VqcY3SlWk+g
dVsL5P3SC25SjDYe9C6jpyGq5kR0ke1SFxfpjlVsS8y7ETutIK7G78o1AemOI6ESWGxXxRRaJmFt
RbdAlhsTq7pOU4ftO5lsyBRo9UbH9Qo/5h3gGgji91i7dctlwx43HJvri8G3OESI8j1tVbd4vsOG
MApBzucRwMT8HvUFGcZmPgf+Fva1uuTHDwq1pWo1W5KF1XCcVJpl+b2Hv0yNmgyVikbu0v9iqCiW
SCfk8aJFHIuTq8H+nWGfSaV+XlYIrI9FY3YeF0BIm1qbys67b0kfA52pBHXomtsbrA2pAG6NC5cD
Fl8Yt165QTsV66rbRk78BlCf4CnfAcrM+9nCprz2uHGZPTYy9lUbthyDloJmeJApOnyBUuMOt/TB
C/P9iD3eoO6xiDC6SymefNA2byE3ApV9F/0x5sIOfO3ZAN3BL45iFMAVSiOF1L2JzpQSvSVB93Ri
hEeBwnXOd6RnbSlL/tmFE9E2HtRmS69rIpNKOWNQGJGU7aftuUIJJ+gb0wog/It5nBedF9hx/aMj
msZ2O6LziHq5NyYKBg3ARDWuhoI8yS0tXKzAv19Zcd0XqG8i6ESR5Ox+Q2bFl0yHY/BOkdRdmhz5
ihgpwIPAOcCGHboJFl3WvA2bMl7mhj/qfQCv+to//49T3EFQD/btKF/dYnOOgmSjarXITpGhSmAj
alcuov2SXOPrRK9532+MfZfcpKoO/uRLVc7MSIr3FubUC5UuQHDCawGETi9GGPAgFzGrkixVRksb
HMZldn24a1o6BAk08HnfKXJwCZLecuYdkmsJ0gwM/vdGYNYRz/qC6PpMme5oMM6e3Bk71r9quZU+
QhnxZ73qH7VWqUNBsY+cKPGgKBPCCyjoyqYEbqmsGxR96kA3Y25HaWuj8bxYHcddM8uL/IzaxWuP
SblccC0ko6+dcad1uYp7m+uqFVUW+gIkufje68PQHOtMPdKS28TeaKNpN/3NDff/UC7iex8NoVMO
d4x81ca9Ycl4BuhHZdvHQ7L6zBHR2hOSCgHXuAeIYa3jTGeMIdpQ2fq+F5rKRmKiY3Nq0H8IGjdm
AADeAc4gp6tXGjfeHkhHInwM9IO+mWkdzNShQdfIFZSTw/V3/uWOrwz+ZKFaUlE2lZaei5YNwHKY
KHv8ffFvU5+eny9uXncB+b61uCSevG67iT3QZjjksEkopDYEOSe+rFczxdzZIqV2QmH7oFZk3ST0
w0jfZBJkhFqF4xam7AdWw//MKyYuPmwx4BZ/AvjmrAoGKQp2Cabqk7lJcIpMDrGzPw74FAzGDRb5
4tQumQelcePm2LRimHwnZ97zUzgmwPTXIyZU4aCXjq3718jYmpqXgNPdG0EQ7sLNJy/IE7D1Nz3J
/NSy0OpGuiV7CR/hk66EvNdLyd7uB8ERqCspNh2V8e83RCKUlHr6urZNt/uGXB1G5f17jvXcChB2
Sty1XA82IDX1jzupefwx7w1XkRlYa1J4Hlhyk/gfzKj31bMxEP9CtoN5vO/vv0AompYclseKZrEq
p99eo7nXW9QXthqNe6eYtnPcRB6Aj/WtOEwW7S0tWzMTg3891cuq8dueyEENobBNDR4si3ayRmLj
tIT6pEwEf23xBWCkkrITOzcC0AjDOEI3mo/88H9qxOSdCiVo8uTk0/0kG23wUfCu8I6i2vdllB3s
13IjITSA+JjOIHg3qigzUc4F8Ss4YYKu4dkxp6Nszwmu6nlB+Uo/WDW2Gwea/G5sQr6QFjoTJSUv
4wGagUV4lliBK2AUrFPkfCFk6YfRwJrnQCzt3mf5DEH3EZZFy0iJEweIhmTwMkjgKjW8198FJvBh
FQA9IoSSZDpO+JlE0lNS4eJ25rDJWUxS8pAFvfZya+RU9AQbAU9h2Upq75IFneG++2WqcghPDoOT
RGbIIk5SoNRohtbOB7CrYGbLFqWnGm392p1Z/HfefyqXoDLQIxhLt1/Jd4v5Y8T6bLPYamH6oszQ
YqIRPCVqJe9FRstJlgzeHHChKSKOaisBXNn6lSLwUD9FGYZ+XP1YpyLfrMXTsILP5zhdYXpobTW8
AfOjOzzhCyz5W4MP5u69hJS5GiagegMN/pU1w9120ZuqHUuIxdRMjkEXAnUECpQ1pvrszwT9XS0W
CFl9eqVYalDOIlYj1Z4nfDBP1pnssRkqLDM6C6dmmeCzrmsgulM8nmp4kjmTmSn4578KFt1XUAkp
AHOh9G44RSwTeX8IXxt38BdZlTTmNgn8t7Wz/cj1CJ7Vg5PnYxSxyfMoMAR8k3MvF3XgMUdFBzdQ
+BZD8DIt9A12m34Z08AxfeV8I7KRZzMHublxQEpTU3Ux3lI4waomNgXdmutZj5bchuw2+AVLORGJ
PQI7OUzXun1iFRrYxY2xeFRyE1rarPen3It1TO9u2V5dwVdeqcLhDdrP8KCfsQ5RWZdTUXizjWS/
ARsvazGKNyjcKYh8njMFmkvhkGjMfYcKc1Kq/cFPZopqc+WKt6i8axWxbOlRMdGSCAMRBz1lHex3
+mVM9fO5LfZFudtU8PcrtmGL3quxP4n4LToJx0JKQAn35LWSEpaqZCKXDXnnTuX0f789uF75uwZO
LN7kQSzJtO+YsQ/1KqMmHzt5aZU5HL18qun7+2onVdWrRjC1iGGojUPr1339uBO+GiZzoUQ8zTWN
V8jgXHIDc62p1ShlaSMqaLepAcrtUVCwN7tX0GW/jJinyjOkMiWjXxsjwUXS+mm1U8Kqp/Jkb4Rb
/Rbmvj5fiVrH5J/roFBHnjZAr/o9LBKaq2xvd9rvmPrYs4c+nzcOtz5dkPJXzBjNJKCwOpLbOk4K
Z+ygy/ZHqijjm/6MuCJp/hdOKgBYlXApYjjQLxNhk4JYRex4CvSJ7ZyuhfJWyqKpnkkBK9uldUx0
nTt7/6BySD5jgiLrZ/B6+JMut0auLUn16vGMUmmc722t+wy8WSOAXNSJSTCekExtQE53xtfRZ0NI
+tqw2QEt/CUPfaaHyyzjysIkyQAHpw/XVHUe7P82ZPpkqMc7wLhLqIT9HozZZ7/J4a8MQ4iR0lh4
SsSWD1UEueML0dm0ElG1dWxXy3/VWyqaME60DRl9UhKZ80gd0sUAxqAdN9ZOGRNxKCiwxT7QhQbz
Wvfsi8jAfpnYal1Sy21wdfc5KUDeMNplGkI0wq2nd+oux4FjkCYe8QiaiPC+UGIUq2m9MTFsixWE
dNnAZvudaw2dCatel8n40Drw4qbUCEo4MbeZcxgwRtqz5WahBGKVIlgAsnQjU8MJ4PROpAPnkA2n
B8ppgnG+/+JfuRMYFYt+vSMkZf6altRz5SjYQQ6otPZizp+C/1B9+6M77YQyOTzRpMp80/gXFPPK
FzITSFXIbKOqQeLMbt4lTjKYQ25r+jhGuI9VW+SluhquvULPF24ZSIyHIkmr9zsZWhF3POhXrLza
NXy7S9wMYYFvwYQ4I2PLr9qIp9S6+VJQim5TZwuMYODwDra6NX18Gu2Lo77PevoAOJ9son2h2Znt
D4P84HD2tbsnnGgMS9yGWvCEsS9YnuVpHWrXAMPNWGMuCmbs9pSXCadmblSPP8HwnptFinpUu8Ib
P/pCrYk4dtu70ZU3FFxzGhITBD0I53oTW0jke8jiJhen+3itpSeBdLBEPTPPKV5ML90wkyv7MEvu
lVyQQIILC+QOenJ69iU1sMeDdgOUMVX0DjcOFNdklY07astxkDfKV2V9iy11/Wdr1q8ZzbhV718L
sVOYWU6nkRxc+cnI/QI7DjJL4BawZLqgfXh473+rYlH2niZH8oMVb2s06ESMRWia9pHX3gXJPPEW
fEoy4wl8lOvVrcn9kqcRAV6SbBIQl0PM4vrkvWTMronUBUfCbnksLxp9PRY5N6jw5UYJZfGLPGUK
4TpIfvtyZMfrnKiE4Ncq4alg0ffGLThK1NXc1rk+u+Aw4uWcCQ3M4yxR5q6U10gqMdQ6MoV2869M
K8f/gselgNtfV4h2lOGutckNYdll9TUNn079YYsXMhZKe0I5dtbh6vIbkus+B73rNTugOaZ8jYzj
+kw0kRO7dQioG4byThFrt8xdUfb1+rkUG2bwB3wnD7FEUaPuIINth2UL49e81uX+Kd4/ZuBQfF0P
vFSvquGYUvmx4COV5oADiEHM1Rk3jE+R84pSEbFdraaQTEUQEVKiA6L0ZJYZojbyscqhi7KIl1Aj
4TZ/g2eeoo6Tg+x1zRwy70nx5PgBFScKQLculYY98vAmKFIU95xBHTwd9bKbhpuLt8eqnXHDx30V
ejor8ZLq40QUvcUviCZtWALVphsE99Ck0OM2+5rLEgY/ctKvPOfeGIEiXj9uUxnVgbYn2AdhNCq1
Ous2mnJL3uLSJvxA68Ex/Zd9f5VONeAcLVqfCfAdg0ptXmR9t3F4kyUMknPA4P9rfyazTuysdglR
AF6KSykrvjrEeX8RE70jqLoQ/3w+OTtmIQ66RY2GTl6Q9kmkGtI8iAbX8Q49fqfK/WBBmWav6by9
4+SL3DL5/6LKj3zqPzu0vidP2p6uyJsCzqDXuRuxomiwEEPwLn5rYi54TonAOiELWq1GeiWsM0R9
QJ464MGcFr/1quec6Xlo6LGE/TBV2+KsevzJQUZIWaL9PQcvq7cU142dLEQewErdd2GicFhm6Cjk
Xg8uFPWapcrWpNbKn7XIMJdlh4nNHKyzPmQoDYf1GZZpcYuKGZPtBDHQYg9f4digS8ndFyzxhp2f
CTIQJ6G3RVIsMrayGwDQFV5ShuoNP+u5/HjKyu57jqJe052JfApvRXap0+dlW3gKCT4Yw8rZQPNB
X9Vx3wxtXuxFaNpPusGYU463LTCozpGzgP3AJV19BqVB4pAYXVaAG95pDYCa9MpkGItwvfC9k83v
T6qdebM9KO78GveYpRGSBAEuFi84xsIvy1IVW/QC39sBUy8P/dQx+m5B/jGvjJSpzHY2jDIGUfuw
xrN3xwnlnUF4qbjsnpoSM9/KM+O4Zt+luJKKalOMb9UkksXDGhpwliOb7VhaZFL9+iKGJE52b4RS
kVvFhYNTzAAWBaInV36/QKq3/DyijjOWE43MIsUK4wlgHF7gEdeR9MvmV3ByaBC14ttGMDR2l2Ze
nFXOuREhDy83jW/mBDyTiYsFLSb7WMOfv/EfNdv75jdEwfUd6ncMZOCgi5VpZuno3/0yxKAqtx+f
vBQCY5LheM8Vool8MgmgXSSMKKGxqe2BGMf0NgajJURyhY5Ewtv44i9CYwAU6UlmOzQQkAumX8BR
8Nbm7wa9e4dJdQmrVOA9j4muym/D/nTema2Im9r0SyyXDYRzzDCvpnSDwkqFcDJdmCK5zwECa2Xc
s33w249OpeQX0RUlfquVq0+0D6syTs6v5qRwDK4mmkHE+ZDp77cWH/3ilEyRgRKKzap+vcVGl+ze
45ThJir0d9qvvXffUCSo7fdszXdWWx5Jefki2RxvIvA0my1SY24z+oX8WCSrkANY0d8FP3tMUZDS
FvjRv3FzXV/RTiKrhYbQnGRDR5XqNgqZDfFmWVb5i36j6LfzapFBUehflzTMWAj5QC1i8f3Z9xzm
TAlv1AA4b9ypfReZWAriL5UU/SvsCDn++tjpf0jRjUT8Hfq7N0e+37dgEzrd+jObaXHBRVqmijOL
P/7bi7a1wchkbWp6H0wTkVBshXAp3RQ2wGRM9uoXjT6EY6vFIWjR0mmdkb4snAFCFW+vSMy719cq
zuGuQz7oRtwbKvPOwoYCZDVMG5DvST3KCEYTKcOL41dE03Plg09m8O+zB1UsVOq+DbQv/qE0PM8v
LdUxbnOxyiysKr+d+qWVw6YXTp6CxgZ63PVWAflLnpR+7SbTkB7e6qI9cK40C2a27kb0E3591p5y
KXhK5YIRy6klvjtNs1M8vm78ZmXKCpz9QC+ifFdgx02DclgoY2977uvrK5eXB02Q4nR1682DuOhz
XaKo5WpY8hlrg04+Bw7W3kfwOWR+6AWtrFvUpGf2RkFM0SqxyKdHC+Gb4M/GB+J/UxhM02/kxidc
BE+S75Sr+RAlkSUh7irY6WM4WWkiP8OamXwAMMPcGwWHWjFqNRy1N83+VZjAYVpnQcL+uGqAeEKo
I7wl6sTTomaPO5SWryXgbgIwHgm9ziXQRb/wxmS0fSUbcQfA8FzTvU6ddt94D2g0t++Rmm/uOfBm
Vv1l/QqndyzXO6P7i/Z5xwPhuVE7rpj3qeVqvrNBY49+808W2EaZbZpPYd7F0AvaGd5R7jyYOUju
9scbKAoHTGlJ4CFvFbGv0dglvqRYMWBDfBIjABD/XIl04Cj9xAMh9mait+Z3w+dZeGEv/6u/KRpb
wmHjAqvRr3hajlHpV2/V5ChMpxKGGWl9aNesB1oOikyVqucKR/2YQQnHF989jUIvTbeZRwXtaE76
NQ6mq44T1Atn/g9BitDKJTW4jh1EUN5WsH/+Zqi8CNs10pukAHmoGcUVxny0fqFgX+MaHIDSShZo
SamPhEGOffLKXMNHTTZ7WaS1o7tbVOKgNfk5ZwfWkQDtfjhMnhOVkrDbyymN7ftlLGULi02g44J6
QXh/2u/gSfnz+k2xoEq7QOZhKic0/cM6AU3pcQBdoBdkhofPCTj6yhfG+euT0PFXekgPkLRjmM1x
7gvyQnEsczbG8sB+n5Z7wt9MS8L/qhKZ8a+fXWFfd4GYOdW7EJ04vtjZsJBSBPXpj5jF05pq5nhw
Q7a+UEHyLRQA/iUp7fLtOGRqM1vVYjFiqEpOcHBGY3mbMUy6fN6TzXMvSmAQ9HJBnaCfySxfCImQ
juS9l28nqrJ88n6QmS0yUHt2wWxsMaAt9F4J8XhRJ0HMxjhTaQO/38C/HrkP8iJb4xFNTd88fufl
/485xZ196rAGyvYuSoYaBIDWAylZiVmWzLfT8wUlHN0L6aDXmh6shEq0yNRfk+FS9M8M177WCPe5
C4VFfIw/wcJKX0YvSOJ4Cisq5JDvm1E/oAlhD1fvcy4EJoxS7DKjs5VFtSknoL+j877KRjf47Pie
Dqr6sZER/Pp0G0yjENrPv9a0PLn999l734GoO1kYfxPHg0nRdk6AyqTzvkF574Zy7iV7IuR6rXFo
IT48dj1WCbcPu9tu4emvwWcsie1tIO6m5dSaTMfn0k4jx2JxU9dfapaignOI8+FfbDMKfpx2Kbyc
KopIm9hs0yIVVP788HHAGZx9x6nr/4vaXK8LbN3i/ddWIkdQu1u0uQHC40ny399gUP+FwIM9XMLZ
f6MYht5p4GVv4WpfyjNQSvbO1H0byIT515AOY/qe/4ekAuA38Vu5mEpF/po1TqMq085CeZ0jNzSf
HwFtg/4jU0umM9I0UFFdFy3DEJ0DM7imBSdbQU81weTKFs7UPWErV9TtNXEM+A0suZyUIGR4nLVJ
1N8QajEovEddW4OFbIGwN6WH9IHHVbglT6a2TFS75nT8i0R6XmmcBE25PtGmn5gqCBPu5eCTUbiM
aO3uDcQO72fJHMMDLc6EtLho/gDvidSIpZ/v3YpahJ8l3SIVkojYovdvb2tY0nLW0OVnU1pyh08Q
j9LXu4eTqLiXok5/h77ziaQv//nyWkHNDLXzHROY1PJjWV8kTYxp22Zy21FK2VomdIIJLk2hFXKp
UbPG/HNkYWFgtVkUdCLzQD6MWVSIAMYCOYOwsIQ9LUKwV0F/rH1sZXKYotxmH+Do0qdgYXJE6cSg
CwY2ZoZXPKMKwUfa8of143ulDxYcYTaFdD84oiyhZgFI8jZr70cuuL8VAl98oS6Ed2lQaD1htqCj
DzGKwScXTTEas0jQLCYx33HbOA54CVZx7P2+92zKrCRBt0LD6N3oaRXXejiAqjZEwh8iBK0uyJWk
cg7F5BL8ydyMO4eu7sF9TKbjHLFHxsAzZz/E+MQDaFi2n3YAq4Q9o1j+w+Epyc7SIxqqEhQtXcQ/
jTQUmrZMbYXuEXmVvB4EGlV0vAGiCKUjiR1nd1FPNoPtr9tL6WWpKpAdApumG2EVFi625FJLfCa+
KI9iQC092fHhIFkvUUHnIdwioKEf7GzBgAdqzme4xw683TXLTwSPKZCQ1jQYE8rXV0oJiJcRnNry
EuLxSHJVqIjDKXQ8qlHQ1Z8TGuEAJLJ4cx0t2m0RBNRRWO+gVGMl16PyI2fCsLtrLga1in1J8oJs
86ExA0MZuz3e7CzVd+SIpJoZw6q+vFd4C5fzsyI0DqBcXFnzPU8pmAhYUhRcgT5SfP7+xBdVaiAW
IG1yAxseHSgZv5TEHf6FcxToX1lpECuDYR1MgER5CqNDsLkQL49CThgvc+Ey/wtQHXR03fMZBPkD
wkgKaA73E/45Xbdg9Zk6Iw2ibiYxfaGDs4qUengLjU6WfJpNuzdRDYQdChH+HMOX6CQDejp2qipQ
p959LzPpqiwrnav7t7OnfaSb7XgJc3HgByBHHVe2ixh2qpYyG0PQsXIKCGNNy3AlvqY29W2clHVi
WZC7j7+1tkfUX+fSEpZuTkPLc52tRyLBmZDISgdUbcKLYcduD2w+IGs/g5K2F/hscFGyvdEsWnH1
oiX14Ha2urD0gD2D8b/AXpnYwzSo5E8OrAT1Kq5Z1Lll+MMvVpoPyklsHp5KpiB3FreKyErJzJfx
ctcNqT1Oeei4RZ92wEBMqxL4LKX0L6r8yk54Uay26SF10JdPQIYwCUYC/kcdpSjHo7BzY3zZmczr
V0dU379+jpVLZQuGdsPExyB5TBAAe/nFgTse6I3PBRkaNwoAlIbjKvxFPasghOL9qh29AniWvgV3
j7VBdkXE5Vz04OgrE1vrGc4rqvTSRJh4tsSrqd2P9e8Db3nel/ccvBl3qSNp/+0vci7r/P4eSQdr
7SHtJ8IAMYvIc8fWFh0PWBHon+xxXD0Nfm0ht5ZpV//nyxG53Y1JoytMz0MkA/EN0KuDmX/HG5In
UwFi/nBXlwRdnfAfZaKCkgIZrIZL4BMOGlELp73rMT7hhSU7+7VCPirbNzaVobnTIA+IvZjX3vCv
/tcHESUxq4dF9BchceM+WZqhX9oorepS+4oVh3iTnqAVBA2evcv5JTYX3xg5hYiuFsSiSM1ls7NH
/m6R4d8/ga120b194JboN4qXwCQS/fbUwMDrjcbemMB+BczWEwKbv2wufceXt4gycnPjW/U0XhY5
xisebqoEWcbFXoDX2cTmepzEfMLfDlMC2gnJAkRsVwPx8qAgcNe/qmv37K01cw86r8vPC8qEG9b6
VY92+V6eQ+remkJ4oma2KQTNgkkC2y9qafq8KItBetjGfNjpLXd9ODlQatzVxgD4vcAOD4eMPsjs
m9uuBf3Wxi6Kb+/87DmdwdpseCriKgDd6hr1ii8fWxyqpK66ctN1xpCbn6lA7XMIaqWgODAm+MG7
0Vt1wtGp5MK0MH9JjFriJSll3w5UOPztYdT5rFfXhFbsPBk7ZSaZWVzbP57A2qk2AaZo8Xz0wiGf
xs8pGlFEDSLa6S9HFgom5YBxGIzx/W40pKn0bqtzp9x4xRzPCykKHq2Pn0g72R5/zl/7CmBKko70
2l6FcwpAv/AnvL0iZQSBZPSNSPSOg5LeHsTZMZx+zj5JTqZhFFUNoFZ8BELzNqU1P9rgqQxx/OEi
s+ZSDzlxOuPAc1yS+5C1eUhgTzgFWO3MamunSZLQyt1K8AO766Pcou3/96H7eoxTn5BuiI7ToQ7y
AxusvQHy8Vwfd5tv1ls4/1Kk1BHvpKxMARDp6yEZtaSdJHFYCtzNUPHzaS/YL/edfuYE9GIs4glz
p6gtQz8T0FcNtpqElZiwjETwzaBDM9Hwj9vpINw3N/j37IhpdG+UVP8i0k2gvC/NpOlX42PZwP6C
W5uyrNtJyiPQXtPWKSm7HuDdDzV7Fz8XgG11PbSK9P+TRboKWqh36E3xsbTNsJnsHRQMBY+DfUMn
Yp/xHT/EcnzqePCy2VDO1n/ggZallMlYVvvov+N/maImbLPj0cLrrY/zHBFEuSSlHxLe8nr82Xhh
glP7WuDSULGg6QOdUrsrkkc/c7aPOpMKewB/h7ledGuxyXDsBwvUkrAPou+5DkMs/Zqc1A3Jk3Qj
cifgQX/t9bTg7EY9wSLVtjp6YTxVi2eRfphrHwh6Sikz3Nqo1x9dLwPob7+nMyXMkLlyfM1G1TQo
n+UqD0gJRxBDd2JNpJTsRR0V7Nw4lgt/2Na94X7UBQFqM6UnWAUbvd1vjcki9jVALpH72Mi9c0oR
fB/FHYi9wnrnTWM6Rd43SklKcXFhvk8soVgmaUQ2zLgMoDYpTnMLEa8dvYow0apeZ8WughQMy8C3
ufr7TDmN/R/4xuIuzzXDS9KJM6HKRf64mFBKvmZ29kQopInr/pn/nsg4MQd6+Z9du30WfRBQjGXJ
PwDnE6ea64ryaqvnhNbT8uZ+nC1VgUzZnTBNPCvz1F1veAd7epnnWQomSjvM1Sc33Cqx/9dtE/SP
RXiQXKIwSIXfncq0zU2nCel9y4qtzYy20eUABDIVV5wMvSCYAnni/w++w0VzKO7p+8y+bsYcDIPz
Fie2Bmt89eS+wFTMfgyMqNaPkPaFW+vVABZdOqrVXkyT696YHHACWyGHBZRmfMZ0yWeIlfSqopdP
dJ9PVt+3kiTv7UkZNOu+bXe6ivIbf/mb6nfaVDzkKCFGabnSS4+wtr+xj/sZ1TALnCjWkmMz7cu6
g8cHtVeLNORg3nnLpRdGzeEcTBG1e9vvVvJZxnrKSU1j2p9kTXw+e531H6lgM+NwmbImjtzKfDxY
nAaZD+6W5qo8pXirkDkPwL08v8F4EoxyItks0W2mno9meJxglbFjX62IQaw5bHirDubh6lLqcRuY
yA9oMfMyzfHvy61fuvawwkTt4F4hOVvCRHYAQDyn6rpIuv7T4wKz7p7Rxr6RLyfusjQbTDB3hwwL
AsbJfR8x1Ebp2hMJxZr+Dwbrbz/YFoNU2OZ9Tb0AxJ4v8+Q7G81GzVcWIhIq/3NcGgU6hHhDyAQT
1A/YLU5bK76+PNvz+Cw0Mtq1esYFSUQWnq9GAOmeL0rt6qcaA79ub93Tf1GpXBXApcwRIIUwUH7y
K34JB73rLBcYPTysfgXOhRkWcqBxOSwiAXNVmrH23iWM/K+w9qxNt8aY7g2XjmuXBwfQ0gXNXIyg
q4raX9bplJLS3tioZOEwnIMB+cAlYWuVVtSwvfYUxuDXWAWsjXdHXpQMnoZoN6ckS7nVtwsr1m9B
u7GkG9jIqC4q998zcz8ATUQjxsEEsji+L8ExxQMP6yKHwIO7gqwi0Cb/i+R1oWGRitMc7AYNO47s
XVvffIZ7QfYSWkgl5boRBmS2k9jnv8oneqIhDFTHCU2vyzcIAybpE/IGDhvZ8HwfJjqVqP8MLcOi
Ci6bRYF4fswBvLm4guUb9L0xnpiT7fstc9GxOuzUuBu4NU10FhXAh8Pmm4XuuoE+SnNWK83gyxm7
qj1WTMuPAMq/c0rFrq8Eu1oKShY95pSU6oohSvuGmAYyJIgS2LxLOYK0CGPsBlp14pt3NzdzXtDz
BIN3Wp7Fi07hDkieYHynPTpd/9LfPSk3FhYVdeKm/uWhteg3xCIsTwLuDu1xCkFwWhhGesddmSSE
A5doB6WvESZNDw1yuAifoN24La/m/7/4tzUosSnuuB/GkMjvyatFEgoRUUVuQ+G5ErBFIrVAAsdg
ffnt0Jy3vvI7fIU+WK1gQrCq0rwMI8NCElK1Jin4XnLSeUJblkpnrK3wgocZK+AcgtOkhk0Cnvz2
79kQ0UGEpuXuipbYjDCFK36QdPFMUcmCBfy2i8VyZhAe2E6M+fb/SSAwGjZoO2nvy1jfToYuOWW5
Dmu9wuAhVCDajiAyhWIrAXcZRdcw6BIiBFoe/3YJ6iH/tXWb3i7WtMxS/sdHF9jozRlGP7wJ+r88
qq6aFiakFX9O/gKZslQ5Tob9c2mJBkVkJ9j4FJ3lwrGPTYUfPg79pQ/roLN1ABCE7DEWgrGn0BeX
0bmTzu4SM2O56hMZ2j3Y534yEzOWZO2UUwDbpkcDM7OZ3OwpEuA8rYY25g5WTfD2oK2YkhZirsiV
C5IlQm2RmRSRMVCXQXvlPyt4ah5Zgn734SMCpazf81wFDD93u02n9M22r8aB39LDb5SxF4Vw2xla
KgAVMIobcpuGoE08++lhClS1ehGABoSENUeJmfGQu2xosQlfKqRVUu6DRIkkNGpwQtZkwiwECwmg
ykpJz7TlNvYiBLUVOvgZQIlrO59AJW+vpb/WLcz3zBOlQ+3P+RrQFYD012RPU7SBrY1bEkOuxNPP
0lt7oFxUqqFzc83geTGGjkK3rwr676o4GU5A9r6AaZtxgZh+cocIFxEI4OC/cn3wRUhmIisHIX+K
1tbVxLxJHr98aWA9/ihaKGOjAY29pOpBc5Bo1GsSLxgApKh5Iz7dj+2hd0Pq6rYwBzwKTC+nlzzM
uFWzUMaT3JxCIvViB7nhUrxbU6dQk0VshOR0H/fmNGp7y7RuhP+VBY3K/eqK+3ZqKwt9tFowxS9c
/rUYQV61Vyh2g5ru3rhDWvTPF4exI7i1wVRqTM/z2zGdKK7InZmigg85nKcmvcWN4XrSmsNWQZGJ
YnRNEsi/tx9NIcbWBdDPyZrMcIaR090eDi1KWHHfhH706z7vJE7/9OEKD0YEdPrQk18Oe3csEdEy
GLCzqyMlFWNjVxy3sUYVeEmSqUA0KCLhCBUmR21XM5C2Ppfc2jiUrRaoaLZE3u6BTe5lCasrPVEB
nNUM1FploC7ShL7Nb51+VzbEKUHuow4GLXifGH6ujHEVKy0uvI2EHNe6xSNcOJ4byZo/zpvHx3cS
4l6V8AbOdg/h/SLAB1L4SZ0Sdx+sH+RiDO/PIGh3DYcAcjvJ4717/bacGvUM6eHG/0zzaT0djUb3
cly4bWllOfrSMCIPQadC+KLZ/U99ltsEIvne/nSUUcQyg1zKyW6IHAPyeDf0LxE7URGCCdxip8ur
u6s7FQUCBER1FQ17WAjsEc1hy8p8oZY4UNhXYsZqcQIJSii78A6hf+FgVDuuiHOC4R9x3Nj5kqwv
YLl6fbqqxQ7ULaxqUtQbWw7c9GwH1NPIgSGQ3o/XND3dbocR6A9/YEz5eqjOtjH1HWQUbwiKF5d8
kIw3Yqf7XQ6pTTwZtVkv9mV0OgqdT4EidFDUHuxvuRaFqba510/MyunJTuzw8nktHbgiouRkLD5v
cHrn4EwDBA5qTB0L1S8bvKCGFVZZy0PZCspGm59RwhIy8kqNNYBhu6HUQPmB22GqR314fySGPjXB
+Q9Yk8/KUoPo/0QJKZA5z3E4BM0UMgcX6HUEweVdMxFUUtwW1XzDEOL++Q0J21FI6LLhoxmzP9WP
pOt4XYVukCFzCa9UoHaInwXguSUzAZNzOtX/OJwJOwnHpZTQr4UwsxW4Hb4LdHooS59Ns+IRlDy8
x0imjt3JuDKDibXFYP/lkjUEGjFZa3dM8puL79xlbp+CDndp9dSX8bN4fjUXiJ9FAG+aMmqsVwcK
9QohANYg/c+lZ1CYn+tu3uRGff6H0gTIYXNZKZypLKYMh+9ULUbBWP5VewYBqhAHGs5D6brdiyF+
zM/d4vFqscC2ZbZ5acjmkI8e9dTFL8LTQpiKq8SWD19Sxu6To2RL8DdhMJEf04scDRkhzo69D2f9
UospHvv9ykAasjw3B5Od7H8FgDCKzoT6+nQ0M1gvRBq1jB/q/kxOZWUBtd68bUc2kJlzMjp0iuuK
SnmLhI6JlFMABV3olFg/IjCZ7XUdcrwmEYW+gO6bIFn9oUYcz/aKtmJSbjm6L88ropdselu2U8rw
Jw4Bsg+ESKFR5DnHZxgJnx/eu5vsWF0yEnE5v8uNO+0DoAhZbHE7KjfgwucjU760X8xhUxTEahK7
Ecvzaogz+TnyokAtL7tW/mCb5oYKFGjlBMR2RiwXrV7OBV8nN0HU1+EFkJ7uFoK8DDQh+uzTLrZI
kUbcAzi0LMdzqPZdl0aptdKjHAFzhcIzhh60FrgSnqOaDZ3mwIpeaioeO/ZthWY8OKL/vn93wu6J
gXiTEtpFudK5A7XqvLGeYdusNAQ9/9BGDXCB8SXPOvxtn/20adNPPW4L8OF0UlTq6UXX9oHU5aKw
o04Dwp2Vm3OBvEk2SZ90JlOW+Vze3PxoK5e2mz9qj1yQUfSIo1Ah9Ix5QD0ALSPMoriizWHNLVn6
QqADbmjoQbypdzQ6lbtOazBWos39GXUqDakwy4XM7pcvqZo26E36RL2d08cQ8JIaFFKB1b+IPcZ2
lNi0dNlr4RFNi+ffUhUPYhXOhChxH1J1wkEwgbx0YrUHI8+WBABthLFWQU4ushcuq+qzADmPrYWj
zW6d5A+HKKXlL4v0SF5Jj37OT+Kp8qE6GIyD5TA1qCCUg2/Tas9Rxy6mIM5u4S0S+S0wiwiEi+v9
aJN66PUcmgL+1CyCUdv9VJU/+8gQvZI5Ln3tv8Tq1kanPad6JXO3yWm/LeVmu5lTCSKEX1q5B34R
E/CFrC+GLXnoe2/CQBJkceoexaTszJY2Om0K6WQVuB/sx/dX0w6wyFanAHuLXuNp54G/SSQOFN1A
VghcajbNr8Qxmk0jD7UhVR1HsM7NDqh1+tFPaVD8VZf/IzCzEjrUl/fLYTmV0m7O9edM3tmDyy1K
C9mh/+7UGJ8nwuvfIyKIe42SSFj8Zs4VwNuwzEbNrsOnfCOE2aEBsJKlLNmtVd9cp1S8N7z0nmXd
kDr0aSzBaUmYpszKXWkNPJbO8pdxOD/NFFyK5N967VLA8kbGSAdAVZyap6hykaATISSLZ/UvjXkn
1kNXLdyKgRJ0XpAnEoLaU5yxxVjSEyGBD3V55N3YBkry/MgpX4pJE0h2Hz6drVOcqSIqfbYUsRDK
6FsFf3j7wWxYSJPjAgw1ePnL6nqIlxpFsifhlzPoIc7jQqxn9Bc96FZw+LvYCvd10llJU0P9mREh
Ng7Pv58A3xB4vaUz589JxP6vN5FFjyx2/v994cQOsIaoHD+0gu1BGNJIM6wIIWmB6UFdMkfsfBe0
JHlDVnBb59hZhoC12J0sxrYJ3eBNJj7xLBTWFCG6751NaDiSjDh34WQJ6Ivs/3bEdvzf21LTYl8I
tI3+X4cPUnZJi4TuDSjTbQIh0CdkgUyV+0rV7w8CvZNx4+dgOZ5P0j30AkxXvPAMREpU9JEqqkpr
OVJYG8kqz3RhxczfZCdlhKClxwNaA/X7Cz8bbeou78olRU/8qZ9rx6S8Ti3TJtDcCR3w+I62NPM3
mvXHe0aOQeUtdPe1HUKVHRPQaIPmv9JNMlrLYAOqPNKJ5/1yciVKtSNK7FLhhoEyqcZx0YZB8Wsk
rAKVMqO78dXldDC2/SU8FHDTPNaotLZQK3izW0srvdX/GhPD9wjXQgrHtycScNyhH1UO+BDLpk7b
Ld4D44YNXor12BmkXDhs0OCL13H6dbEX1VtHWrsVL0RFdqUu5xzPPWZzcCRERBQV7aEcUxb084o4
D5Tm3/kHEZej7CcE5xtETF1llPCYD2HkAD4p7KXkfnk7Fo6t9gdL47muUcFDR1HsJfAh4GPj0OT/
YVGaWEP9b3nSgs+kYAro115s6THi3JMe9kNPOn10xhA2mUih20Bpd6mN9bRigsR60WY4JvTc+AUA
l0hA1/YQjwnIhCXBys6wwMxtitAf4AALa0f9ZcTflo/fgjvwdjHBDw/0wxp0Co35LwKI5gOwtk93
rpag8I11rgz2ts6+iR21AvzcnUDm3FjJ6956tUZBxwnx7y3L5UywGW45p21IodPHPJNJ6BbmJWPr
/pQ4+xbEwT7aqHkffZP7XpcMA8hqyc4sO7E/uaXHI4Ab5/a5gSt0PnAKP7iVqr7MQubOO5PG01V4
7sA22nIQtFqZsi1mErgeit/Uix4zlGvr0BYYBX71rAES5Arhr5ZJA6vtAugoXHqZ6m95wZlVhZPj
ybRh6xhzn2j8AdMb2e74T2B5ARCvgPjQ4W38woddTka/CdqvAyxwckeV+mECV7lheofVWnZX+QGX
uKSTh1A394v9g0nwS9jJ2bhXdFsP+AQuMvXWwNLYMGnSpf/2+FYeZhVh3DeEJK+XC+r/+KaS3jdE
lUYkiX/mWUt56xH3wdR1Erf9H6UfxpLrVAu89oP9S9Ob6P6vtp2OBGdPKnEMNSyLJQC7dckdJido
oNKX0PJJaykWw2b5W5Kb8iK3mL5IIk8OlHz+Nx3W3Tar6+TtmexHAh9W4Yox8/+49Trb4xRqCAxS
x9+gW6vc3hUFwMruDn/UAsvTtgUV0Cnh6FuYikd6C64Kf2NxaVfU0zWCdeogPvwSEJ7iEb/ds2Au
z9F43iIJs+VnEvnKhxDm8LDcDWzaQFwdB7PIL6VFI9vuFHdev7xeXpo8RfJ0L8C8PfACxddWFUib
1jSy7TXSx4S6JXSuwLRaoRIfUdOETGtOi+MFA94BEEEUZ9eEdDlzWt/GvfFmrjJyTQfh4Y5rcbp+
gN5YP/fhiddGjGOidiyV+pCUBqy9ku2MKMnTeVDdBZcvKXxwiIYiya08kWBrQV8TZNtWhx3W37LJ
FHmDBSX+dqmDHXpYT1ejH36W6ojsyRnzIMtHyzBk0ltcADXSnuOhZe1i13ZZQ6PEMIOX2B3FewAZ
NI9WNciJofJRNnnlBWpFjSd6L/3IxJydCJ6MLtt+zmR7+slvtr39w0E1PPDGwCI7fJYLW4FHOAKK
DffAleKc97WUrpgc+VyRxhwmtdpLJKdUoq9tLbnAJkWkX93ra0eVGysfToluakE3S5oZqD6MV1kC
25/twiyjrHccMhcJBk8krYM9MbyLqDcRZ00PTg2SMpBOHaf/kG1Js+UYtPE9LE0f+2F+oNbyZR79
dkiJv2okMcmVKygRMZ+7yF/KEsYuRC5r2g5vee7VGEtK2+9KuaAHMW1V+JAWAPAly9RXlIEDsFfs
1UhFqzTaOuiPyTeHEwIVi1K9vPVeiA3g6Vbn3892KyO68d+yrphrFm3wTGmdRW7ZJT2t8BAYfK9c
K4/zNy9F1c2NhUcBnIlYRQ3aBTfusRieC6u0HRN8I0tEZw6W06gyE2C4/9GpcsiVamzkvI37guQc
Qiu7gT8ILMsybuD8uGvlnml1g6eSklEAwBfp+mhcyW+aWCKM1OTa5eO82bqWrb+rVPAC72a+IxfD
CapNahldA8lyqT1f49SdBTXF9nuxZY9b/zGUV09FURmGi/tbtPYZ26hy6cF6NLh3JVDCw5sBTiuE
FpHy6SFt/LizhVKXT0A7iwVTyviIMjDvI+hLDzPcZp7tqSrxmjNgqEnjEi6oqcChpSElAgsb2Dsd
HXoI/+KSlFQnkKLt9+7ddlajXVZVekfxnMmIuSWAyaz4qPdCgN4VoLU3TujxUQd1c27BW900X6An
dAprd6AjV3e8q2FW4aDusf191/qGNCIoNq+w8/lRhnR+LWc+pm6o8AVlRasN/Nsq4+ATKRJpU+qN
Kvbr82gGKBBaZO69LoDei/Nlmeud1e4za1FikN/Q/i9vUeQTAQYauG3wjKgRv+4uTmnOlb52tP4a
E3ZRfyT9TK6TPGgUY4rK1eqFz86nZ0KvmwxFMKhGzTNWhwsL5wUHOVa/WoIsco0vF1wPo7AojnUM
NO4dUEyLz9wr/cl2KUXGi+pqFPerTlk22EJrewMKAXZjluMQuzUicSg+ZP9X3cUJUwTV6IFUYB91
H7FdLKgT+Tuc8n2Cp6gZbDxfEfStqYpy8OS/fzHGMTUmBr4kEEAy7bWdTP7lAR7kmVDEjWpN3DNE
HID5p02SbWLGHKDBJVLIwPEZHrffuluoVMXNW2bfmrAahFTNLSlXpcKaXrakLQFua/LcIxnBipEg
EDQkWGtTp66kte65ghJS7gK5E9AsI+mGjlF9A2dSZRGq8kKL/8qCPbYaW6hbc/AO8YnhR+i/xbqc
Zod5Sm4Obr9AVjWdr2SxW/OPZ9r0mFqzVNqWj6hsClcKppU/J/oJ4YnqsQD4RKYrG4zxLmk8YVRY
O7P04gog+AxTNhhPG1RI61N1z7vONSV9q7UYUc+9X7XGwil3VZkFvXgfWbwEP4T5GlGlX2BJ9mQH
YjHmAr/ogqnGbXXCbXzSuzS/WiFLEeZIuK0pnw2ZKSPprs6bjV9oHVtgRBsJNyA9LaERRf+/LK1X
EasC7MjhwQfE/AdCjOE6V2pqMkRgW9YXQQ7zp3dWIsdZQq5PCyYrZ3A63dtVulHEN0mwVDQr5DYV
oeHwS1mNSwpJxkB3rAZrD4Ngs51WtgmXPkAF8Wdzqxg3OZmug7sk/VTUJaKra+o0Uoj7USJb/to4
EJJU4J2HERWxdpJojmhqgAq7pb/EXGp3rR0Q8BJDrX/u6aPdKl/WhJ+QaECSZtvYS5aAr46eOHqA
nJnd0kj+5HeTetYHwz6Y8OWHZZ6oggnVbY38SbKJVxiotP8JPfoHiK0QzzFk8ZYSfPRA4EIms7xk
Fdmh7j020lqeRq6yH0zz2lwknEZRBsY/7SIdHIOpE9+kaRj+r2JPz7Bj78GJ8JbIk1dwGg0Ilk1H
7dnwapENbBDla+psTYNAbRgBFMFwqulQYuZD/a48N2Pz/vkpkeO134R8RIaOChZ08aiV24yhZSR8
uggsCbwI+QcKFW0ObW+tdxX2PT2mPstypj1m9jBMhnnqnHjQ41rZIHV1nipuwr/QM6Qunt8gsoWS
NZF1e6miyUvMC8vdfu60MEskUHc4IuHtRhzmdO82EBqjDC9zYFrPE3jlxm7miQMRnIvd+YXCDtFd
v47WT+Ncq61ha92AYk/fK+C/ErkJ5j9HYeE5SGHQp/pP+PrF279ehZk4v0hKkIS6gjgRITfR2Gzy
+bwi8soqavhpE0O4DQdO7tn2wTE1AOjgVXp8Xn9j2qQkPXDlR6KZ3ihHRkbwpYsLeTH6KwtY0XOp
zO7mwqKL2K7Wf/rVBrTdCHMsoOGKXBUguufMpEIYUXndUQIK6Vttg+o6lbjVetF9fP+ClrOFPU9f
11RXExGurWJVdkk1KUJSNJVdmZw3IUXqskdin4O98adL6sKoW06O8oZpNtA0lh/h4zg12xbKokEo
mkr2t6dL/TpUFsKIpLcIe5R9fHZ7eupyYiq1Hl8WxlBCUdV1Vd51C7HLGjMS2hTtIVvpf48hJYT0
Tu9QYQWGKThn3dClWGABPSyMeFUtPoqRutdB+I/Fp/rzQB+EKoAIx8JNsTL4bQG6oP63pnb62yky
NDrJnwfzrXw8IzVMeb2ll+wNZW1JIElElC5y4hThQQYcoyaSfyQV3HdL01Z+YmhMT0bwwKA7jEVT
MOq7h2/ulqupPof5KWHsi86vjUCTu3M5bnJ6cVi+mftzKFwgG0z2e+wPJBxfERABA4aoCLCuSsgX
+hV/iU6SElzHlFyDdQk7ThuC/aip5VdUcja3vTs5mKLTtL8o5BnvXVB8Q9JRr4HrkeicadQHcVW9
nbxdXMw5sHBDGLX/k55WSMq8tGwN/L1DmxD/1hvNVHGPLYEWzCoARyaKtHF9jiIl4ersfsbVaKup
zzH0OiHfic3eszGglfgHHG4Xqn0qM6PZ56aW3Sk+qjnXEScHfghgs5n6JcfaW0ajh9mUnnVgH77V
B3BDv3S9d7AA/s40RXo9F+vpH18hDKlvAWNOIn4A6KLP1prWrTN+pjG2GXO+pPHCtJcZM9R+nvDu
sEk91iDLgn2wOnaXmYlIYx4c/fChJBbmMbhAIARLazAs/MaM7yS8i8d/+S2+H7xCgZY2T6vm5WU+
ZCor/GpflQEOwo6B4co2AfvmQKqdC0li2rUZX3evRPvHgFZMb/J0gSvwFdeg4+OdIqUoAbUPrp4d
pZohq5T9GCB3tcQbcA+Gf2jhkYtLdXWF72GD8XmolASB9SUsG9WkUC0VI00jrVD5AuTIqFtHfiy1
FDmqJ24NFR28f2YO8ZZMGjX/nit5Jy+OsQ/UGtGRHXayk0KSoxy3/jcabquLTDAEobh7VxbjkFMs
r8IanIwfgBrI4TFpGfwBsvuNBGgOSZM39gze57a2Lni7YYEL4i5v+Yv8XBpU+f+jRSZkPwdn5/hu
QGiPwKxrlZQAg20xZUDNhErsiKXztpARfqbZqyjvm+Gu5Lok1QLLC7xl0IXHNov5f513y53aqqFI
saPGF9HNuN6hVUu4S7DP8J+ha7MAXEIt1MeafrgHXA8z88Vzq2iYSY6jHhYqtsXeUv+znus8Mtl4
/6RkELZ6qjeoZ8BpDLejGO9upv5isI084BbHIaZLxR6D90srh4jgKJqxhAkRIQWe7rd7zRDnrcLE
J26SWCjdQlTG4h6sQQiex5VkCsyvVErTQz9fgJwwsa3DKyoZ/swrIhIHD4UYwXKqhgXgbHCrOED6
UCWpgvtLwLaExZpux+TWEUO5lB1MVo6BT7e6I7gQ0YHtCOJth6h4D9yV/BcqIbTuBqY2/0G1jCjT
GCWitmdbz8i0Qcgg23eZHDfxMcFs8FeW/y9MIfUe/XSeoq0j4qo8P9bbiu8yAWcJcxj5I1iqleg0
eOXroEKdh4AcL+btujwOncZQbkLRtzWD+Uu+feaPZo5TAnXHkjF6Lx8nCcYm8vRj1eqO48iVFGIc
CpmWBivm13uTj9XwVxRvAIciIYbQDMtQ22sRx1LEFN7MDqD5JqeuWUMHnRlMjSyDRvhnsdGo5lM7
5HAoB1DoGO597DlkM8I1IaXI7TSPwBFwd+mImRLfxV7YZq4FemA8ylgApdJXN3DFigjakAAtmEYd
W5bHG3LJtCkLT6lneQlbbtrfqw4qfjFc/fVkp4+JjMupaGivoUEomNPxD/t4uC7qkYKeZMEj6UCk
q4VdEQJJquhsOAnwFNy0IowVt2cH0uIYcMjIxa7e6Y3yOAM67FvXydCcqSvhMkhZadIHnQVVtb2w
FNYlHS+LZjh0vcVGT0Qk0IQ0AWs+gAkfwLkTw7G9UeN8Nls4gnTvIV+ZzOU70qZ/cVXNnzoi92gu
xiip9QcFYRq+DnsOF3rj/4y1tM7ccfFptLDoidG2lN01rEh6nHoGib0qhVSoB3+mbVoUKbgGLS5X
tGGTHcPMThB2plGlAPq7aUjTrx+nAzyMYbJhsjLiyAseGz3JkDQHqAdt/TgjRDKan5s0V8bT+BcC
Ji9K5cznpyoIVzsAbp1BlfsgMep9KX29cPb09bbt46H6rjLEfCvLYLyVGVXD4V3qpR+ZqQ6IVoXJ
ov12yjfQ8XMuQbibW1D2ag7WynEa2tRwKLagJGhrySiCGZAQ7H3yjQqK+aFy2ydtiyzvZC1ayBhw
ztUlUTPT5e4oHj368vK8mvhTaPFCPgsIRBj8snte+oSLK7uAf0inTM8ij4sGcmwdmO92K0QhIlvA
aznhWJS9kqTc1sROftEKOi6irt+0/MlseomFy9HZrxck6X9U6T4l8KwC3QAQ5RcfKnxfd+ed8jfC
wV3Y0UZy3Kz4VRhR+PKnbTlTL0fCvDWPjoddqvKUH80BVn7a/I1IxC+4xo8AOVuA7YEWJ4CqJIUw
rOpo6MLwSTK4BYIKGHn4q1jMyROq3Gjw2HnBN/YFFfnw+yFjnSBWjIheGWu+m89OL88sQSMNEQmi
pxLcvhbzeI1eeY85w5LgBtq1Ab5DpVUPAZpwI47dpW4Hkaq7W5PCCju0t96LtFUqQEEyo7EnAPY4
OC6qUhH1DO+ujGyND1o0ob3DcnnORS5o1EbVX+Qparob5qu7eRdjubg5//TVz60ZPy0gVy4478SV
gQEj1Zz5f8N+OQIyas9sL0Ie1adjgjNQfjYy8O4A7ek+KmEfCAw77CG6upm2aD4sA8AlMov1fE3y
MyXAiqp5y43ORsBSxujrx1C8nQYodTjzfSFg7MUYc6YqNXN1vopnw4aZx14JZgRIFieF48kxaNcv
R4FL+9CgMMxKHC8howcqqTpyhKljMI9J4hgAqT8+/MEEAgQR1XBVah2wnCm4SZziow41r9YoPjDi
/YF3cCh4RXXN+WZWuGhl6q5VUnXtp2owtr+1gHQuJbi7V68zDUXVwMz15rPoIuRyWOGg6+/A8R02
lmrSdYhMwsk9urH2zuokwHARaHc6nI0M+FOg06istfMZOc2YzaXZ/DKRKMcK7mDykc4ed3CccPDZ
/sZYozMMp0bpdG7Bxwy9D95ztYzhm2ARunfSNH1jWcDrhoRmfV3l7UbDVzm3scI8f7WvzSTTJ3yo
0vqwvXqdPBh0FJk6AwB1sp/rV3CSE3wJt6s+DL/MGh3M1tyYdHJNoQ/aotLPqhvY9wXemD9366Ve
Ouf0W5JB0aTGhy1vk0CD5QLFc5JK3OxU16CWDWUqNFN1ehaZK1OdomiOrhRSy9V4tNl/ep4JeJom
T4dbbhPdDnuClvvtRo23+rFUgVjHQ9z99IxYQsGrRthX5FCqtBVvwKNWrsqyyHtBe/hkctzPb3FJ
0rUrZJetuAcNCVHhv39cpwr5fk5dDHQlrwiMXCkpAx4J6ngZC7IYJoDijitw0Br/VRf3Q+19hMtU
iy8Mltp7AshZyBAifitPqYZBpez9R4B0oX6yuDzjwiC9cGe+ENFpaKOxttH1RB7PQIcKzgE5NvUJ
0VKUDCoVqOrjgh25G6YmHwHYCteJ5FJKUuYkI6NAx5KgRits4Q3S29at4ppxrdTb9UMFTJEjmydy
2SZu4bbh6kt6yln1IAw3o/vYvO6vpkuKVHlhErnKwlbZXwztbf/+i4P0tGWK0dWqETccHNOjM3MI
ecf9TZ0Bc1SVMfxzjBaT/f5j7r8exxzeohofEkQTp4sn0A4bm+cG/RYO5Shszck2ERjbjeZDOsAO
psctKwFToJxzo8XO8yLWLKR201BS/0mPSVTdg/4tm4gUlpVC1mNNw/IC4mrOojbKcfDIGsdxRZGQ
GfBXFbz0s7W+z6vL4/MkZTy2wpSeMIKsl67RYIHCS2lu6fdf8vUP4dvtHbGwmDirGaRbmses98v4
AoTjpR5POH1YSHFDBKmTpl83iyzKGlWo0Wu3Xar8zoD/KQnnYLNmLq4yFhaDR/Kro7IPb+NXXhOF
ujySLV0ThWodYaUV6Mn8K3JpzKTIy2rn/lWq+vOaM3OxTg5l4OncLeRInt5N6ALMF/CDZuQN/VLX
XZohHkPGYrvN4DCWA3p24iJqYmUXKjYLqdgVf8TATiSIdpV9BNFNAxQi9tet8Us0VzcbmvIGsk6Y
WHwYe9cWj/sU66O7NBrZ7NAmPetTbqooY+sTTlKiZaoJDF1pQg5tgTm8jVdII3If+PB1JaoCaC1G
4UFPtNdrZA5ixRnCuwgSz9ajkoTYFQRSEHwYh6/UDQ6PYnwhpDD12sKPbo1YypSvEm+PufGYGM9w
O2GPO6t19/nDnc/qhFEiTCK6Epdfzd6jCmUG0DETRT17fAQvF5B/ppWv8tQXccGo36+LdXHQYlpP
acPxmhsKfsTjyUHAheXW6WYnRwQzeznYy2yLoEzp36rgRFOYtKQ0laduJdYRSi8z6yH2zaVZxCYj
U9YL003hxF6TP+Fdfx1pjgrLymSVxJP8HbdwyFsHdxnXX013TQZmbAQtuuyBa7AAma+JMSRqc4yu
OCxa7o7VRm5v2lf/tqH62ceW4319qEqYUsL5lIZj2uj9au+WmkvdJ1a3jOg4d0HLtRStBefBS3Yn
17b0vGHKTA+WmJjixX0Vlal3SQsAfT7W+64gesuN26BOz+D6j9n76P9FZofj+dqssxw8x88BAQk6
qxz4CvRdUNVv3ph+Y7igd89Aow/kXJSGNDnF1xLtaV8hJNS4OAjbuFpKA85JxQVfrVHYSZe5xykN
gVHz5TP32VyGBZjhA4ecAOVALg2jPBp2xPOFxewgme4GqUaS5HabGZdLziLsTtl4Gyn/fItPuHcT
qd93Ip/BCgQfs2h3BCgxHLcJqZLYdl42k0izYM2SQtpHgWhd/0W6hDD3Dgd2aPEQo28/Y8VLc/5E
niVWzK7aO2e9AQr4KM5GKHAPHMamrt8OKdsqPFYTU/HU0FOmXCZfJcNgvgdUSB2WluL/tyKvoBO1
o7rh4AfYFnMoqRVGuPOk+lk9iLdIlrF7It3uMR010j3b/k6h7CWLGxwhi1NxgIudsIG8pt4p4Crt
rTfoOGxUtdk5lrgR1DMa/xy0Tr4c5Tw02goP5ETR3TBMP7rk1yr6hTXVUtvqoqPY8k2/dn+PO2TW
9mG2czIRTfjDcGhmmtMIuEpQlqQehXvWKziJX/jaczuUio3CJjt8xLsqoCxXMzwnZWasuATZrIhj
LGFSzGQf0mHTEmayV/qtjawlbTKjOhtOhhY9swBxONNiCmdyT//WSKmp3/J9itQ3lE5pOhvFUg6a
34Ria5ckKP71xOQ0APvBi6i1tcaxtFN3TtmTMA0oq1/2fQxfTkRrEE+6VL3YdPprMvuTZzqSoaoD
qQKgeoI825RYMQXj1jTEAFHdl56UwDBwQQcbigB6UW2ocswFwLZhrQ+4iguyiy8iZZKctQtPuys+
N1bMQPL6C/xKcq1wHGNW5ZGKcXmHyNquQ4LEIZt05CHfilhZ9kd3W1IGYCixdnHV5BTSse1S3NNl
J+Io4PeFfmH+qi2HuqaJ5+NweC757Ixjbb0jvtK5NVWJl2WW/P+JFjltcfdukvG80vx/McZptjjq
EK4jncQlOEInDeOalFpfhaAzILUvbW6fvFSe+LZ9yltNx+DmQDV41HB0KSfXjpcjq2HCzcdwSt/b
49se2JFwQwYO1nSbS4RsMclyfDGVtYOWgZq8vgo5/i0w2vXwguKnD8Qk7m9dY1XXYj1/lzmVU/Qy
dMGFbtbbkqDPhffFpLQc4n7cdYS2mDwyA8sc6AUzCvPOMmrirvHPE6wg4oHwEz3fOVxcQUZgUX/c
MZJbzxtV0pY23zhPdbOP2+3ikGc5XAlu0gfbrqRxgYqu0iU0SYCPlKE2tMZkQ3aD7waZme9TMmJM
Oi/z4w7Nmw30vgB0vps5KodXJidPruBXETAqtkzltS8C6D0RS60O8jpJPgMv6NrMgf/YdYVMUckO
EPhHt86K5QWYBZwdit0K7GWB3a7c15ctdC9yGrU834QBme/2O+7eig0Ubcd0dHN47ajYM9RjWqfL
84p1yXhOk19YAV2aClyPkReoVFcXOIgSJaY6wN2JEps8Qsw7hF+wxntmSK30gI2EWTfGwatEcixG
whv//rIKtW1rKPXaMi0Xk0exaFoATTbY0QONjWYLDGPO6p3o5Elu7ywH/Auty822RxJpP59v391/
AQgDS5f4KABwO1A1tJY6TfzU6I0IQxKjCz0s5a+xmcvIUIUdcZ5G5bfNT4xU+s7O2DQeM9xZ2tjL
nj8o9JIRYF5NB3CMi/kfhgVM+zmwMN+ECtW8E4SujJzJrvTT9Yys2ANsgN9iMDz1MIGuStQHbAn4
Vh+07JTLNzzrT84dJ1k29jBTY8y4m7JH9Nx/Xnh4lh5/GFbHphFlny9VTjqb+Pkl7VlZOt6G2Q5x
mKM8bPZubYJ5VVsy5PQJmep8W4yjToDrB3EFSjMtFTFu8rmZ9vlR9orVwpltnYtOKCZXrBJTm5Ds
EH1B7/cGQVxTzgBxvJK8hlrY/5dn7IF0Pu6hBqFa7uukYZafasegwapXHYf8BLoluMDiSEElfhVo
5j0otOggiK6FA6KDVir2B9tdBtL3YQBj+xQI4y9Dd+RMQkbBrGDHiK87XSr20pjzihgYxXtCo1zL
sMc4hlmpxhttsQmBOFHsDX20vEPWFExXzVGarkSKDAAnOLf2Hhq2CAhfruCG0ucV6y/CxWxbVVa/
bynJRT/5XrFz1viQZkAQOKE4UnpiTT6S+NvA1HlUsLiCPknfc8TFG7dQ26CV9s3UqquWSOweyRk7
EzBkLadD+4zYxjcFGNXXs7BHZn8S8gcuZ/0MEGhMdlEDuqEwD6GvPY1PH4GsBxFzjJSoxqlg5M5r
JJE4SOIAu0HyRr0D8clhJylBrN9DUMR9qh2fDyHSUYgTUnS06OgqeOzvpG34FqbIVlrNCB0Vt3Xx
v85S1632pa8IMZf6WiTW9lOBu7LE4IjqngsNyXdSLzt50nMv4mdkwnWMBVbw20UZSU1KWmKSA2qf
+H9rydCIMCfScdir9zP4peVEvJY0vdaCWgHDY0w4ENKIHwFu++0E/ufKYyBhlsBy1sgnuon/QUwv
GEjdZdg3QW2D4cf7lik+6nkm05+f/L77E0363Yn3unV3eOd0waceZLYeXIXEdix8PsV01jihPf1o
wVXVdCto5ceccXbl1dgh+szzSKTvYRptrxLWBiAffU6nusvrbB3CAP9TS3ttkkuCZMivqF0bFgi0
M1bIihdjTPutXudQYu+B5LGMkardjwx/oAQBHeaKfeDSqNsL/yTJ/dTXflTlPUrwqWVA7imPkZkK
hy5IURenW+Tu+vbZee9Gk7CwtN55xySy25pbNpJx6kzq/CNugIn6LWrwKOm1ORqjH2pvv8Ho8LTE
cZ4zyb+zmBmkU1Mr0Qk/qO5c4Yl0T/w3Lx4FdxsQ9pVQhSZfAfTmIUepB5oAdhitwGwJY34icucz
+MHie7WUzavfQTVlVBlxtjlfZbUKGwy8ziosD/K6ekW4Xw4Rg26TRqK3mEdBDHqzFGHkZbqNd1UB
DsWJiMA+iyuU2Cr7l0cVXD/sP8lzgX/X88lFWaf2z5yplaZzHDaeoG8sATgP/pKJyTkgFY7H72tm
iZqyloUoja/GJ66btzapHe6WMfYLUTSltGJM9t4yXo3fs3coMvGgRN2pt5WQLe0injfM2BaHDILs
fascxJLUhmp8cE2FaV8mRU+MuhImSChVC82vCOq+a0dfOFN/iQbXR2Rti+oU/J02SNneTZmwytAN
vbEHZcyst1Ez82gymdf3vTT+DYM5v5BqLYAEBbM/gjMe9KCr//M0sU8o3/fC0QA9QloVJYWRytUR
2GOSPMG9H+KAStm+eBbEa9Pru8DXumet1hgf5sGcVbGf3+2OFDMcNi4t9UNu82hk+RDDr1XCWgeJ
3CJRZPgyrNggjfwBGQb8IuXw61lOq8pQy6ReAl4O0lIq924vUGiE5prKEP4Iga03kSRwG2GeJy7m
seLn2cADgvy/Ycvu8t0MWW1+zXd29sy9p/QYfNEUVfhXNp5UzXqJt8SIPEsdaR1GaDVvYC3TfH5s
QEkfkZByC5n1v+UdmvqTOnydQV2WIxGgW9QgEJzfb8woNrl3+Wy3VTePNy/tMbPEwjyqDPXfn37U
CVm0HDZ+nYjWVR72RQPc818G5UcvH0o2klBP1saDf4ELvnQeM2jMhX0J5ZeMVrbtfIvSDtWjFM/4
tfkYG05P0vUW6TYsr+7UTzlgUOFHqdyohO3fLHbNBqBaD6uJ7bwucu1cljbw57x5H3ng9HYR01VK
wWqujPRCvxAkXDZ25Y9rPkIU2WMttWEqzAqXX8Mw11zUJJbn6qaqcUNS0MVaglvWY3dkuZfMz7f/
h4+a+KyimWHDLtJwmGFdxWNRjO5juwIbKV5TuE1f5vZFnhq0T7aA5TBh/QWZDFBztBlsqzcBXgmg
GixybJAz/53apa+/0htvOvBrTmBttk4vBh69bYKbJeGIgTLEV6vqruAdnDPte7KZ+OMFZLBjgiu2
NFVGqhiCDJpWjs1yt/qK0IXkYQWVHocqtYQQYvBs0w4uWc1Pjxq/8cApvOsJSOGaZQQg0k7vWJfV
N5PlJcf95d/UN7W1q1UuwYNftR8vlPzr+Z2FjbaaDGYFE4+QcC+uIyrtgDeY0ViCEnODNuXm44Mb
U9AiNCiK/7PJ3wJ4Eqj5cpEmm0il2NIVPCGPlcNkfxn2XDRDgcMsZ2Pp32V4NdEU3Ww30Uap+qNH
eI/HLoN4jIPcOHOpJOaz5IzH0Wnvy5xz3AJX/zitt0PzpTD1+2j8/Iery8B7nDyEbFjVSqKN9UC+
CLUgcoa1H5tvI1tAqdxzQ0iC/TP++YO+SIdFl9r7aYh32vB4+0B50yy2g8iJksGUKidMEuoYpPgg
TAcENyVr053IGTtU2fy+BKNMBBcl78tUYZQF6F9EJFycbyYYM7DK1F+AcV6UBIEm0NmkfzE9oCQJ
VyGZQTOOYXyNu2D7iDhaYo3d/z4+ltno1+5cn48WjzKLP3NprlcSANuOWACSERmDNs9ITRRry4r0
Dq6H2+l43bQ/031uk7W5QHWw+dXG8GgpGHH3+Hx5L0xDdlDjPVq8UnlIJMZ8H9c18On3n87VZK8P
6uRKv162Qpyu/B+7njbFC5KZO6QOSPuHC58g9NltBrgBL5ATqN+9YcfC8axhOJlZjSPFLLl0dq49
5zjBSBd5nnG5aQnxMMQJ5Il1he7c3GHmQvGbtsWoFC42j2+ZULk0bSSrBSbrJLWfx/u01fY3HAB/
HMtHbaKU0wU0xs+gnG3yziawLa8WP/6G50g44EB8x9O8FnlYejFoK6KR85aFqa9FbmCefNR3EIoB
4tsqYRFT3CJjq6oQyxNEPK0Q6vO625+3jOqOJ1TtsrblC1os+otblaiWQYxpsYmwX4ub/lI5AzaA
HVRM0WZlwWL6SpDEIARUKo3M9m9tnUGh03JBY73G60xJ+j9vfX6he5+l+AcuaKBbgr3VlgZvVJr3
9HoZPiNaj0UMWLOYHDGvhA3PDNknupFhqD+KEx04FHFeS7WvUq5nD22lRdYrSCLHveXCgB5KjOzz
pSTTmIBeuxcAVbLOqqTnu0Lbq4+m3Ihs1iowd47HhXx5ssS/SzNqeELCoeNArOPQAxIW/2u0GuYl
RzIUGrrHp9bmABiHoeUtVLWZGgmonBrax3n0rG8EkdcaYhIxfB6ujNQAQZ2QZQuPQbi/v7n5qZT8
QFA2WIdC4JfLXVVAOdmm8zQPq9jaWSz0xZQAHQbr07obyrJXn4jqvPObYIKMaRrqmFixzqcF11Yi
mHTD6HNN46UfUY+9cFb4rkN+DwDr/Q1ZqNqCcgI7FTjIMbes17akf6ZI1uNgLycT6QlJfKclW5xZ
yum8khN+xYq87KJtfAy+q7CiwdmVIazvM67C6qZaDi11R/iW2zD6WTODSZHg/onMd4kuUVbi7Eov
noqvMDwImeMEl8ffjJxQihil8PXCaCuQO7HqGVZZBByszOKFJ9rYSIRLJFi3lHsbGah4+E2FPrG3
UNw3KZdmvcEK3VpHtyYxfGWy20ixr7Cp1faF3c2U1I4qUSKm9LLADWhkpVrqt2cBFG+0v6h9Cks3
B464kBDszYZXdlH4GlbdGujWWuZg7Nf5zisZsnnCUKTVLD3RpF43f7Y0Ww9L0cB9YEMsye1y2HyU
HIa6Y8TZNXXfcxtfOBQj/coWULNkmJOeRqBN3IO9tUNvn/T7+gFeMK1uB24D0ChPIWhtmNBYWWBn
tkJpYKeAGOMpBuOpN425vV8oE9zzJHwZ+qmzuZWtQADwTyqRfVdQh6GFruf9swi+WmT8OcWgTmTD
J3ZsL66cEts7DVmchgjefqBhnL+/Mf3X0xBzBFeZeHP0lbhS7La4/a5iukcsp1GRkUwDdnwnc3hd
i1z78vEUnrdik78ueJR/Pr0pFdzR7q5YeZNU7ZVIjQn3APbgv0dgHbEsMQoDael7Bg1Rm7Y6E1N5
VsVD8yLimFIHfuiOX8F60nSy8YUBUGLO4oDNhYZLPJqiGJQH+LUf7fpmlWCBy589R7sExn6zPGuS
KJjXlsRuq2SUOOusgp4+OPRd1QKaqHZ06HIvhNG5RbFa0g6+Rw4TcUZs0u4tjdp4M1g7WTGiMfe1
AQ+bZiZjeQ4aXo+O+/H4ZktG7yFZEjspkTmgMXnEvbVA3HkoB/4BYFGO5laXIS1UgW5IQdtoCvHo
gOL6Qpjyd64T7EzHKlPbHd8l9CSdb1uKSJTu7BV+ocLlUgyfNfR1tWDgQCIL+zAttEijtN3Pduq5
RqEEFoKRetPQt3cx0cENzWLwhZHNE8mPMic0KU6O5xdlLmve2p0TdDqWLHuR7kwiCbrFgC+p7j7F
n+3siUX0g/Q6ygBWqfVTfF5FstvlXffEI1je7StV4AUTyt06wxnC51T6DOYhZ13vyoIW0oNgFB6Y
BQxFMTXwCjHZjYbm5AgIH1C5qBLwkUY6P1b72iBno/qMYjJ+zl+hF9G7x8hu7k4ZUKrn+20JWC2D
hiCnciNe8yZY8v4RF94YqWRIqMJQ0Oj9EQuzen52tiWoTLf4NDoZbfwZlQKtVc5DcPq9CwyIS96a
HdCsHQAAx5xZ+AtaeQlxA72mpggsR553gF0QBKEJx7CigV8JwrFhgtmQLAMPndt07JOXowXafmoH
O86+mtabnbEvtRkCAbCnnnSzuZGwA0abQNY/oCq6/1gmpbohq7C6t5bw5Iw/9mmeltxSQ/F2/r66
gTmoJAaPlpAV1QYrsn0X8dvC+3fD6wdSBg0YAmOK1KgothXW/9gZeDsGVSobGOCfd1Or4CY91J7l
3pDt+ZyD4odwqkye4sP83cX4gmc3CDHFFIzjkiUQy2N0a3QCjebQsw82mUbNCULHz+HX3ooEZqBF
W47gmao7nMuzGlQqbUOxg9qS2ST+Yrjl/5Vx3GPdlHklizD6SngCFngEQUcVUI3Xv/QiLdhbwxgo
CyAWQybdWTplg0jAy3wvYWumxy8r1ixMKvPZcB+RNgDJy4KZHPqYuznI/vNdFaJbG/shDs+oIUy6
7f9hAO9kuvfeV8EMg+Z1Klz3AAAlCtE4/lL7+uaoziJnJ9MDwaOQ3nIhpvauyXjIdXqCd8lp/+aj
AfBR3WO1aAaq1aoyOkAWeNO0Ig26F/zaLKpwDtck6hRbfjJSMgnrQuV45AoGnheVDR9FqLea+RBM
SGCUWXmQz2te7Amz+753QuzxzT+CuV92tDPN2wpAgNWAK7NvG+yI6wQ16if+sCy8uiQD3lmiTkOm
rSGD92Qrq1zX7TgXCSQgEIwhqGOR1tyV2DuSuPyFcRgIbZrKHdMiGNWswDLIeobkEwYMKRCszA0O
xbXIdGNB998AG0j84ZxOobVspKfho05cpZZOgQHyq8io58YWSkvrr2mjhgKeGCJa1vTwKDDSgcOd
GHyMFgChXj5TqOEevw5qEWOZlPtI9Ma232AeD3df3rYnW92xy4/bWK2Whrj/0yNhqlbxzwXhlKTl
3ZqT3ptuDtgAAGMRBU7+SCCkpguOcncWHgzlja5y3vJXxfvaBYphpiNXrGnGrm48VD64btRf71FS
2xGGsfkKWQBzylsPkmVcScbp+aGHkx98v744AKnXZdEWgoEj7y47OaAcGPUi+oLBQi+XbeG/Kj07
xthKwarmUL9zFAibds+TOZ7tqKCP8PinejG3omBoZxqgy6Dffx/7z8hfSP8AsKvL7JFcuo5m397S
hjRLT80E7u3+cfoMBdyVhog47tfkiSzeBdXallaBn3wtHWJvcDIBbP98zPKhbhWwitcc5zQDQIWO
dzsf+a0jp9S9AhdnVHS9N3Lx49YpLxwmAOorR59YrB1DG+Hl7mdmlXZVdM2PTnCp95OUmn8GKwkq
6mS4d+3Q2dtm07be1FeMlV9DwAZclq10XINRbVpsTpKxO+uzwx6ky4bVIGvcFkPKr7L7c0sNHGDg
Gv+0r9dzNvGYsmsxxk9pcNxPinirV1bHgCITzJyInpgA0r1Azbar5SymXt6WfayI911ZcwiJdY6i
5HOZVNrSRoWhymwYgNWhzWvnQ8J9tntLSwLATBvIfXoBFtzh+GkXdog80NIY+atI7OlqFt8sfV5o
ciEZE2086ES97sTHT91oEMdhBgizwy2ZZ+OdlLbYS6qIHcGUOPBzUaD4UNL4TkhJfb0uIgmBLTe5
UmV/tqC5d6YDMuNjapflrGuVtBa8Ob53AHun7wbygSFhHzYy4M2Pz89L6I7nzjKDTSZ5+FiA5nwo
Cq0NCS0PSKHePrs+YYsGE2zpZjExxSM5x7pheS7NAX5cv9f9UOTNY88YwdkAO45FfRKD6X5SZpCO
sm667yFHJMKkKDJ5erUCYm+wxEb39At6IHsaK8tL71czfXuDb6ukG1npx91snW+6+RQhN6YnsjLQ
MNmTiEfdYnX6bqirUJTucbp+S1M4wKVuieOhbRs1aJiY9F0hrGFmCqv4Swn4jJ+Ym67oYkA7sATk
lvn3+zWhJSv0Wrm8MPMDmODuPPigXIeH+zgLmlvYz4dt6qOH7HFGus/clCLf/epeMje9eZjc1box
4btKZIx8FSK7V60I2kEK/aFnQ+9pkPh66tZIbvwBzXgSKsuP0jVEoc9IbtHJtgNb2LkcTnfpEcTV
XFGU3lkuVGeg2qzYhy6574OwYitQsZ3HYRh468pgpHOxR64E+mZC9xjqFeOAAxThflAgEMti51T3
DiqE//8Mp/o1AfNkxd5LayjJFPrZvJVr4Vo3r4ZNgDI44w+2X7hVC9ZyJxj9fIDX4cx9y1bdJTHQ
Bc6g7SBfbdCd7waHnI0i4GwS8A+tWtOygkLDIh1BE2nBj2kLqqS4L5rx+UIxeLJvgu7hbqdUwErB
HFo/UG+MuRpL+NGNTnY/XeiCQTHzVJNllIJ3gZ1SET3GROwVIMXDOpHbLjbI9rnd7zFEFoxpqWUo
n5ROkwGb19PJz1uEk2NBrKtugOKSiSmr9ck1W728aA8Im1USSNYtBoH5UDMnWIe8/wx0omPThNgk
Rl72wEhkp9SEH8xFwquToJt60q0P1BzBn00qWNRnu3PHe5otz2OXpJqq9kv2jwVrpaP78T1UB2Uc
rMDNCT0nTeGAgpzWBEsCod6MSeBiPariivqXQ/5//yGi7iDfuB78fWfxQH3hGlM3BFvI39Kjax8N
qYOTmY5IVlGSZyNeard8gBRzJPSENJkp3fuh06OHwPJ5W+PN7KmTM9kAUuqb0fxzWril2peu5gpZ
IJEbVeEzFoNWakk+zxZbUkFsBKdUU9H/KBtq09eA9Npu23V2dfXwblkeOl0VqvIVY54q4twjQ9fc
UFIUOHmKgB/hGR0FcZ11v55EVKfvK09H1tGP1QpdJKBUFYR4EEoQyP7lW9zHm9q4VB0ST8q9yYvn
LiB2+028RxODsOQcvJQ0W+TsRGIbUrc6po+USmP4em5aEljiPUS+wcqIkKHVmbb92fuajoKI6oiW
bFZIFezwOK6Hd29XFByH2CRix8Cutx+q6Lqaw2eJno4TJmjKA+2lnZsuH7hnG/BjfusrBeXO00y4
1hHPaSfF8wWDyLg3OAJ9+RYlkO8fM4qkJtTdywWGmGHcl9iPoVIqZpm0s3cwWTM8WMqvqf8WdYqb
CYXZ6pTezoBYUuIf9uYheOd/qDG8WJtYn7oF+MjukRtwwFp7RMFFCZlPKJR7ceeMjJyW9D0NulTI
StGRlaN/sDKS6x+6qO9EN5Ok9j5nvh2excx1HUc/WP1H8Bnz2GrSzS8xQE9ilVzxth0kQAWHXxYB
2ISNlEjjzPsI3CVErm0K7UKQOdeQK5zQeMffThlLxWgLdqzDqnd+W1G/1eeEOb6/am1KDb+T0qZ4
VQL+T3rR7k0zf7+IOIGPi+kYcUepilsHU0fYlzKYIvQ2kuvnyfq2kXLIA7hdS+jGRkH7lDLq0PdV
aJMFZMIM53Nh2w1jow6NCDwbP2HYNKKQByZX4fBAb4AEVsq819LPX0IVijtm8dQuy1SOlUlFDT2U
HuhFKzuabyEXW9FCt01HTyyJGv9+nzd+CCQsuMJJR1HeNEfvTrnQkurGiFKVkV/fKzq7m2ipWLwO
eoA01FUBPe3n6s//rs3C9HPFn9o6PGFaCOpJ5E7oxGi4Yt6axwZAMli66W7aoWsWjGR+GH7JPua1
CZcbZFnWLOHJiaGRK6yPNBB7Td+tUuKUooudzsWPHMwQU6VD+nWZGmaGVcC+1Dgu0aiY1Idln1Jg
dYpLm6QNiWpVNONueFrS849F19944rPklvOIqLhgJ/ZYH2aoHx95szhKe0UuA3TqIQwFPp7Vn95M
1DFkxHWUCmKoU7sqNgThiQavx2AwcVLMeHWB/z7fDayOzgEmkpcSIUN8FA/P1kC0UaxC269iuELI
dz/xZFiCNoYI18smE8ND3c8NDvNpKA+prBSnmstmwyazwjH+rxYz3eLvh0Fa5Y8AJ+MDNIIJ5srW
2Tn6WH5d9xGiL4wTf+3ReY+yhsW4RCZsg3uvdKoQUHMUlcuunQ4Xx4EDwsiQFPZkoKYlX4mwJNpT
JmTQs1amDz5hBtsEAawe2j8slmrwtp3eKm51ucSGstkepPkDiUQH52hZcCPVB2v1WT8t55LKXz4/
bJkesrz2IIWIXGd4mxMP6AYgQxmSVLzsUuG2JliAGe827P2RV3YmkhlFzVK/q8NSF6WA3ReSrmtS
HhF/xBZN3X/Sz9rGiEkbICRqow4Ud+h/AGR6gIyr1TeZmyweADvZojfzxhE4J45Linn6opl+iiwF
kjJgyikcw8p3oFH/81NeKRkc+fSpSqMoWv2Ddd00mF5Xb5gtuaNqF0lQ6JUQ31Kqkq3WUfIQaIsM
R3xRFcY8kwjTj8kK+V1jzXIYaVc1t9yv4QlVoIS/AchzQ5ZG12Dnx/ZvSKXPxNzmDY0QYZ5PDbnU
xAhqOscYX9BIHpzQQMayPqeOL0sSVNI4AAoh2Xrc5jOPkw9FuAseY2evUcKSwB/+7TMLYhb3wGNZ
YZTcY0tVlTQ7h0EyG2AXMeBEekpRCeBHkRNWf6QF4tvKujSN547brDv25NyeElhzSqFjmODftdFM
0S6e42fBMXXojmWr1SzhZUZ5Q7rsyzlYEaLYZdxMMRgD1VJ4zj8v0jZbQ+HM4diONKGq2q8sv/y5
ucY+zZ01spfAKN9/MsgwDn/gpqofgbzdT/teGD23ElrEdsDAwjXNVgZx6Ak20kGOVOFBr6HP6c27
FCsc+IrmuydmTA5afutuAD06CZCr/SmBNHBLmNIoXKfOG02ypFb9pA33746EMMwn/7SI6cWHN3Qs
Nyt2q4uL+J1bksV7KgQNcywCDWe58JiHe9cPLt39FnyaP+0iKSqPveh1tMz/QvIAqnHgykHW9+Ot
i4dh4Uqpty+6txdLkKmWF0vSBsqNI+pKCVM9ZKXUU1NhmcMaH/q+6QGGQNFCeK61dvapgREbWy+u
trSuvuSW8dR3WQrrYv8XMJ0pvCuPNylEPRiBCID6duGtdVmiuUlhzotIXajc6JOcpzSsYVeEAcMx
EXCLHaswSftAxUxLNj1rJpCx6fc8/zTFpg+kZ0tWWRP1Joej6QE5L+QehgMu3A7/n2eErwQIRor8
DwkUZZDiYyPCTx2SoyvmQ6i7lMIAWF7GykH+cgrozeFknOfyQtP/kD7wloOaA0+dUHgP9GfVUmml
mJXCZM1BPtQCcDsp6yszM8aLXO1FB+rjWhpIqOXxeZcC6/dngIwlqWtP4CUaRF2DljwK8rqYAOFP
cEdr2ELIOkLo2srk7bw7NzxtHxt1rBM0NkcYLphgFTejQRIqOv71swDpdV8WKNnm09q94i72Obm8
0MyPtBPedbNrtM557IMz7lo4yu/PwUKA8bKI3fuBAzWzhoFVUSOXTpNUnL12lk7GKVGl+oAEXpJi
rXcRLYtnD6bWq+T3skDYTs/kJQp9ApxKwt+2eVNgn5XVQ1CtfSd9njgpZWrKSor4SRUrwv4Dk06f
ltsY6302PLHUbVhpOm5l/cPKERhqUVSs/0tmvxSLr8wDHGyuqoUvjXH5CMcMeuIn2VvE1h5iUEoa
ulmURTEr8EE6wSxJ6cgFqqw46DBEQ8Of1Tt5zu9KYSUXkddJ1eQlyjUTbu/Hw7YsTD7qfbGgdc2/
OQBdiMHtmLG6ZNv/g4cnsn2TXKIlX/GeUK6dyt1u8VGKGhIZXMxv40gmi6xZlgN4/JPf1jbknd4E
9XiwTqeRgRoZcMz2vqiv3xGt2LtDE/hWB1uQVH9xYaWL7jHsopwdDVI0kK9nBpievoRX6qiSWgtX
lEZDSlrx9D9fBe4dKiI9acZxyxjSxsPikbrXSv+mqHPSM+4mJ6ZsNjo/gzPu2S/648H6WaHcnh6N
0l21V0ZH/Pi5jT3iQaKwi+1+V9eTRkXq5h0ylkTnKHrn2E2zC2mdGbrTPFnkRvyEb2RWoNy9zjSV
iH34Xwu0XKve8me9CYwL1UdrIrUM2C0RmKe6jEREyU7VSbKYKVc3UJJN7fECXGKJTt7xsk67Rwej
f/hWlQr4EaAlW7E5iPKTd3Gxm453wpdsZ5/HzbFKqaVFbgVmE5bHb5lqJB8uFKG2yYtXKTKpW2yr
MCoaJ8bIFjmTS1+UU8vI5x4LkRFfpXby8U5AnA6eWCK1fBPPsVpf0KLZrVvcvdjFPg8MbYuj1icQ
fv06EGzhdS0fIl12yAnr/4D5QJuIYg2fVgaUdhxhuWtJhAm/NNnlcJzmXACHhg4RFOLMxs84ULxv
TdsrgDTtLDPmC/OIdObZluDT/hAG1VdJATyM++cv3C7JvTespW3dALnx1fZLWEQxQdULhriTAUBi
HbRFGVFw1NuS5kfmczdTVXkCLSYJ+R4mJbC6yVC7iI4PfNa44rPWxM/2+MaG/Qw13xi+IpxFdVq6
2W2GUeloXJb9fLelP2zfsQUApnbjq/CtvNyrLaNIjcXk5GB+lD9Izya60MhmLI0Zla5RO1E8e+E8
3k0KiZT338abu2xV1U4nCU7oZ9C+8w9OyzZUF55HPhc+oC9YxrDUM83s0rbt5YH3fT0hCOCo03mw
jqGeE4B8de+0YGHsNAhBftlxFwvWCcCdlXyJHdx9K6QsjgCQPfcve2eqvkTB2fi1YIOjwzJHj/JR
eD/tmShEi2IEKzYj7q8vXGWJ64ZnepnDuqaZvZgc3a0+8aGJnNtg7ca1wHmTEPW6nrNspRvJrVU+
9thfva6hM4q+bTf1vsuY2S7YTjqqGuIz2xdMSmko3m4yovA4Xygv/PTPv1V+hTw5jNZOZQtIZw+s
wuyAPkqXDxTGTIUyF2zpE3aza4GoS9+RMi8CKSE7GH9KgaHNIsDJTxOUFSa2gpVzbSIWpsjVR+GZ
T7JcQ/iJlYtySCE+TSGn+R+3pTTPGbg3hlcDim7MIklweF+W5pJpkJjgIJpzvS6SH9GFmbo0rHE+
SVm0HwZP9g92avclsk6gJUV4Bh0vzn2dSF6P105QnkltvaAj/yR0wmRzyyVrRDVkiUkpbbzc9D6J
3PWYkZlJgEzlDRWXqErz9c6WO8p7NlRkcnQ9zhndqacUc5+r98zlMvuJDi2LClp9S2YtQ95u9iln
poII38/d8/4ECVWoiFSTkUYIU+bFzvwmc2JZVmyYrG5jij1WIaryEcbvv7hAO4o0g+ftqJAy7+Ve
+HLuPYipwXjRpXOkSOpwXoQNAdik/3kdfYZBrzzwViwg98aX18XkglMGe5Bme2qCKlhr0avAjimp
5suosh9/41JgeaKQmaK7xrBmA3xec+du1rmqyEtzSJJYjCYF0IMWW5kEsUmD230CAK91nF19JFo5
1X0AmQix6dxWVfEHQdsGjnXBKnwWB/O1n6oFyTpUWi3ocvUnHuio5oo88O0PFQVF8uQWvk4IHgCO
cWL79f152slbB6tifwRxerCgC/BuU+JC7VWC90RihrjryN/KzaeYagjzbPL/3jFcrKQ5wA68IbAd
47v2hRWWZN3aZ4S+Jk85FwtLv0oM7IXwQKSYSyyICaviI/tB6/cGJeuT2sj6SBMzjBcJoA5NrZNB
gDi/Ose2OI8bdEOMaHwasimexu8sTxp5NR2uYEHU4mjViFwRZo93isd0/Il1kcSiXNFvNzM0zyxy
qNtFur/Hk1RQOSH4LZlOKDNABoNbbbQxE/DXVj9QiB2PF/3FNe6ckRk+2dxtV6SM/lb4BYd8SNex
cVnJC0rH6HC4JhnnpCdtsorj2LZPN1dQUCWbWDwCC5dzYR3ffACGUVYzKb+CtQ+TV0RN0vYaf1OX
tk/gSCD7Ig5TAyVEFmvdzeX1MDf1VWhCkHfTG4JZZxS62M7T5fQO3y69IQi6RzcgbHDDcPXgBLVI
ruWHi0+V4XJnlp27HTEvmCfraKrAJ5dB/RFARuRUKTX1eVtxFteJtx5o8eB1wWMnGJ+5tO8DSNLq
NVwDk9Sh8BGUgqVm4mV5acrwzLO0lXzEtJhu3fSHqP3I1jZvae+CaXMmpHcFvop4sU/L77vr3fe1
ZSCDf8+vAiYrcge/d+1bU7LUr/RoYclXndYB3huJ4yToVtFt8P9Nshu+ff14cPO4Gigco4zVWjjZ
DuCqtN1Ctvk9TmSxF2uFX2ZHY48hNL+7KQr8YMolxQN/jJbpk/l/MO1MVjg4Hbo3LPZTrs/38JYh
MmqtC6SU+pBeXjRkDFDUnUi0JsTVHvGEUdj9LPFEcea7eFdHJba70p3JTxfLX3NxJc44Lv2E3Yre
upe58rIKe5jiJU/doZ4/PF2d2sZ5oQdJbJ1vH8yEuVa00fWIE5aV8830BMPMzj4Xm1nh3EwBh+Ya
oW8RnrSWIAdHNcmfb5POHjrxl80ldmpcaEiEBwP4zrqSUeQovo8uMzyGeJ1ivLi73zNpRfUtdW8Q
u7mGksA35jEyO4Q5s6SlQeEhz4hEz2YHni6zRN0dEo1TJvUy6DztmJ4CRJLLSJ/VugDSKHv8yFEN
ayKbMwP+UM1oq/co5gjE776HJ1lHTnMcS93RJlflxzOppSU4BRhV+G3xnV3XMcZF+w5z9FGTVf4e
GRZu1NtuH6sltuHbJZEEoJPUCFkkwSgR0gBsSh6v3cGMsD1rodM/4Cwt8o8Nz7Mz0ovCVnZCl/xd
56x4C41KVfK+mZkBEN5zkrIvQjryt2y9hrQQ4HV3oeUFDXR+4R0gTw4xRtjIDgzF2Hbogr6roApA
WN0sB8x2BwjTKZP9Z6wB/h6SrpS2IIWFI69z4l4bwEjc5yZm6Z6ZISqGfZmliQ4xtHfz9mNG/6yA
4oOXmeYKqAI8v0anjS1gyGTfevV7lG86k8nCpo/+i1q3heUNJy4nO8lqfl8kscB0vdqW8OW4D7ta
T9Cg2o6OxMpcH0eVxX6czgsT4JT0wZ8Z1AJ7dp2asY0FGF26IbqNIddYpFMJlowvbu+DxXb53QFO
V5Ce6L17foq1ESpJOj6pN6dSiVoPtHFa5N+cHMkNb6nD8/rfeXu81aF7+vNYokalZiTMsFaoUYyt
SeUkrfQLzdOuqKD/A7nt884tA6DZTykyTqwPyg8lYrdwI7f2rFrLDROS35lUBy2eLXwTyAwdPNdw
Tk8kwyLf5o6oZuE/IjqBkDbHg5yLfdK9mgjEnfSjdSD7Be9nuwxM8YHNN/0zvjwDVuZfA1EznKpM
ZtarpYyDi2eaI8HuHtk7Z3Dur3w+6Pgimr040juzmP1XqgRo2vVrQNte8F/BNumKfka7K99fhFyC
3p2PLRzI1xEyDmTAu/hXIWSPWIreISyqOkQwlaD/zAXfcc/B9azeBAU9TnBnfJ35LQvsyYEf4UCP
NiN+el6L8IDU7HUkiD0UE2l0nmzgoau1WGwX3/4OTriMWIVETURTCiolrCnf7tXfaKvqOIRJ+ZGq
kAqHlYLF2llI7R98+ddCMvAJjmmv1tiRbhEeJz8A1Wt2YXBUEJTo+oj8LZXEZ9L71nYNSvalGRs5
M+j9VFfaY2eux/7FUk64YJ+uKF0Z2E26QqiUSVcaOdk6OrnWetAsQXlbULIpVSbeRMJ4fxu2Y1ds
zrOYj7Sp6WRfHbLvwGNq06orfG6U4ZEHJqinyG246Gy2zNdjT0lmZfcnr6tlT1zbxKcZ5VaMi419
e2cQWUj5VN1PpSfQ2fiqmi3iMsq1bDM0iA1CNHPnHA5eEQNNukvY3T0eRNHwtup5X0Rs5oqMXaXE
jIwyi1yURG75rnec9AavLZBzWFS03kaeAQlIJk8gOnTgd98MlFFiTf8Tez8vennkzCHcLocbLsZU
ClvzzTLxvTNnje5ZduHJLJX3wR4HhA81OqoNTxLCFxmZVEFhCDNceM1SjfZh1rxWYioZxAv5oUrc
oHCGuIFSW++LPBrYEh/pZ64YfD2fFjRONVzzVyE/pC6IiIlsFYMQD86xCjPBcfcW1D3+Gxu8oz31
JwLqapyUAfQKVw1voVGYKNfe29HiXrMfA+vo3NBEVa/d5D/doKJ0qvz8oNEePA0wCsKhD1oJwn1s
r4kEb22NBHVuJ+O+BL2DuNXq98p8YiQOjU7/MaXiM3IyuenaCR42JWKa6A+nhKTem58KL38nyk5v
kKJu8krLW5u5C64plFI9EsfccJCzvswrA4ZZiHW4pv6yaNaczQINz99+VEbPbKJ/1JKZQdiT012l
xQoSNOJv8WMwHWrAJQubIb1F+kSsU+PSdr6FsMbbwj6oU4lpwsoZI4Y1tHjQEII824iAPxdNHs5e
rMjc3/pDWnViFcvomosHAW5LaYaRMClnHnI97XP+XUarJyvFT3REdNqON/hGsB+EsWmAQT2Vkj5s
m5ZUOMOSjFMj7+TfzP5YIIPNExb39Kwf2QNUamtAm4LF1ZTcBfyCEGoRS2tl8I9oOb3+yCQGxrOW
oWEBrs0N95kYhrv9nWPtGdD/t5UoBm5xHn0ux0LOfPPEjAwLjIXgRnmMSG7DyRXKzdGFUIBle0HP
UYxjPwfxXzYkkLGq7ac7zMQnOroOdBdtTA0Vr7KtI3OG3hhoGUhv8hcI4ET6J3NdLiQWSlLiR1mU
AJBTRYs7yRvxDpcwWNXXJkRVXIKbahBi9skTaH7YUwFlp8t7pNAlr/Pxo2jKZ8qOy03BrJKJJ4Wg
9BLIs41Lsq48s9Gpsuh4Tv0NDlqSvnPLwmUot9RdYmvpAoVgXl1Zt35Zu3pmaAhbIUZRCMX4/7/J
7ZoteldEIclUNKeW2rYwk+TVJ2RhsqPAevTfyhW7tsTncYnewMiriO5Hs9I7PiETWujdntKJlzBX
fHTZmQoouotKVZSrd1+owoe435ViEuwSn0jiE76W6/+d21J4pFCIPe43qgFDWVmvqOUxeIHVl03w
5VAAcLr3k7zzhDBwOWxCIbIZmZsnz0Rtxisti/AO7kWNpTdUX49L1cc4t1ihkNE9JqAoeIO0tYFv
htVNSViFwSqPL6xVyAqAuAHqezm+x8FT6YDa+JsSZEGd9e6Nnp3fBxxJ+xd15pQo23SPWUpk1DDA
7cNlKUTgXx+JI8I7uszNzpMcWFlrMV87yktUb7I2SQhCfBNAkaWn+CVyFq7QLAoLyPMI7NeZPvaX
nLxM82Ma2UIHw7gQ7LJzZ8o8tPDr58svmECmgNALV3P4bU8nLXZMzJc5efrUFMfBjXg/kRnelhpD
ySsZXUdjn+pEivWjImZSeY5oLdohUnboOAvfwwJwyQuKgBm94OEZEpMCi1JTm0dt5io6/JTgAHGm
kCKHMyBX5Z9JNr7EUgOmyvp9WuWuHMNTtP/VeqUdq1Jqb44wT7++I9EAU90Yf82LIuhPb999flS9
4sCUTi1u3Mj1AMdW6Pg0xPlKY7H07YC19d2k+dmdfaHHEwM2M6DivmczlZn0dWDyETwPOm3/r7WC
18FQZaz6DGWCaibLKQ4fj3vAdkZdM5QBfWlZ1rmWMsjycxGiX475NyO1fO/Qmg+yQLgIgDtZ3UOT
PEh+g2AiTsH3p76d1u0008VCFez9l6nX02z4m0wz900dg2YwVPEIi7XWf9wLfojAREyTyGxFxMfX
EL0YQkd/UIjEZKNwDmWzH0TqAo2QmLq3JAJKTpdxov+t22MWuYVFMdwN0UmO0aP42rzqbMKA8mn8
KrftLXY4061tWTetuXjyQlGQSNuuMdOgOGQf9rIH0sDZ2uad6m94jFN6CPEvFzaDlb1BGJ9K3Fy3
6Jm+I6+C+cTrffqjtEZ8l1HtOVXKfD5yxdJehTQXfx0/1VlG/Mseh+QxVGyes5KpUR1JvK05ul1k
D+rmPDXukD9tMhyUueOc84x+unczEbmTkZ6Oh0wTlE73kjIwaWdy9WnPy7b6nSCjxz0Nw66wvfA7
l2IiqK6Mwm3o4DEca52RioelgClyaGqJx1fHOETIb+F5aBnHEeyF2P+pxqkAIw+1Uv5b/eHJ7HTB
OarZbd+nuvEsQLZFq0e+KEla4qf6F/3p44HBpK2mkvKqUINsIoY0q1Tb3W0Nn5Zbsom8TFl3jJx/
+yX8FRpTd5EuFtfq+ZvdmS5AZ4pqOCov8s8gUOZVujY59Fk9nCNgKAORJJUIRLJgRbahIYQe/chW
FYYO7AbBL6V7rnp8TL0CJ/4TDokWOo+RiGk471AvpIgHPRHtQsiuQaX6pQl1tRB14YEN+/gGYmYr
3CwCMJQ+As5m/A5xerMOk8ekXXN16R7CVRWqTCK2PP61h01DKN3Bztb4yb64BFUFOWBdFQPO8FzE
LY5zEPXWkFx3hw4g/RTKzpiwtk7unyAdCiaq1fSD3SPDDfN8kFiEnGkQ5bGIUEpwn5l4e6stLLbn
v2+0I1iKojed/hLgpZpv83k9gQZ+jQnd7nD0z+N7JKuxgDSBFaX0M+DfPv/zNHzdKzZlp9aAGoXZ
MhJOXz34IhGByNXnfCxuuklvz7j5tCtLhB3pgqyLgwTh2RrNbS4A5Yso7D6vq2ZK6tx54gZ1hUcZ
LYvVIGxghm4d+B9svF/pUs0EZ0QKOp4vqd+tPI+AJ+Yq0cqlGglNpapzV3UxH9GZGQv5xPxQHc6a
eNkcRjPwanZTWioxOxZP7d7C5+BHGw1jPw4Ub4ls0XfvM5VwCgFuDOD6fIJKxkIZTL5p3TZBJMRj
PIdGLA8bDplwv6winvqOls+MWzib31XvSevV3AA7UoEoV3sNCMaJMPQxxRPRB6lwijqH6jv6cSKl
XdDEcS/eDe01wu6DehC3wmuBvxvHYEpuYZAox2Y+zQs6P64wAkyrXu9kvov0l5+38WJtjvhYW0cD
QvYoEvJfDdTPvA/7nBDEdYdC0ksYJpHOm/zcQXjPKYUWU/IB2VJ7J3tpz3bDmuUhDqWjwi6P3656
/+cKvD/RB7GW/0jryXvz4YurPDgNhGyN3lQEYvp359gWjLg7dJPEvpmyLBP33+ihAKbKWEJtlAFd
FCrpaNX5NVeBQF+bRMiwbOykAS9HW1rR8lOz9XQ7QBHNPSpaRmZUh9yBHBxazY8A4rDC5n9TRUt3
RixJx7WPU5xooXDi1QBUGtoFSV1xYZD9Iz4CRTxw5zEjbrPfgtWl2uYDgZZqn54u7E3/6qh+X4Z7
M7uK2UMXy7iEJlOQ+VPSmCat6SnEwgS8leuvZyVhgwnmMv7RsaRrYofSI4iIOmYU1FCHScijyk1+
VBShylrZJ4VwOAASt0YN/X32W31CYeFbDLKadJwQo6YkM0RIGuI2M6ZpF843mIOXj8YoY/zJWTJT
A4FyXNM5x4whAqYIbZQFTUfZ994bOdJ5BwfMlyTwcjvGl1MutahUs2Ahi3FQXMApOL4DDgyWxAoh
GM6H9QTlzzCscCqeZ6DS8DiU7ZeoyIA96KQnT14WQ+Jrb3RaWDTmiDOq2rx2hdWvIFsS4C+QLUSO
jJr052ACo5YM3ScLw7stRRZhQ2hntUCFqPfYtO7CoBAjHzkM4WM9+Snfkq2AaF9rb3kop8kaoVXU
5cypOyxK70vE0WirUO4yXWWQpUloiNUekwDJ3+RlJa+Q6x9tf93sn+N2X7elBDSI1XijnK2VbzFU
jMAcMQkQziXxFsCPd5lIUUxnY0XQVWsrCWji361zyQBKmAso4YhyVWsfCNmKEPfNafpAhcm+HsKn
nCflUhizRY4jqcQCCBzPIcGxIraeR6T7AJE7HIJe2a5R7f6p+V1b5eEXf3msX9SnvxtGXPfHqMpt
zwc6+k3zYUglKSXkMwg0dPbJrVU8vhDgHdu3qHaWclaoEJf0in2az2N8x88BfVaoKxoe2kqt6dBM
jp/iz5IkOe2RJAXQKY5t0jMGXqtwvY09WOfIR/Jc1NxKp218avMqVP8KwxuBY+Gx91dSBNVjPp+I
Z2jW7JbF64Y3BHWgpogJbEJNtJdBVe4U6IeeSNaMpY3ME3DtYnogqASenEF81lfu40eZgsFl18u4
A39x3gdYlA0PpZboqATEF/jKCDue3cqobd9sEpsfD+dKfGzXIBUasqLXLzddpoyrq4WHlOlongc5
FRmeVXm7NOIp+LmUxSZxk4eMakjuTnkxZZv5QVKkhxWu5JJOojWxNZpNOnMv72v0yUoJ0lpgriKp
cTRot6Zn/ivSCgaeWd6h7qGg64VqDiHX+FQOPX/4mNe3jGfV5u1XPgtI1NoOpKumT7zBxd96FCVb
Gao37JWf6DTrkRSEz/gA58Dn6JV86Hkhm1h5Vvv6SvsqQyLzpqz8hDFKQomEnQBRxWJluexsPl0K
eW5v2zl5qKiuOqLzW2qHwzTiFKl/00x4dGO6Qebktt3FweCdENXh+kgpWPZHSoQ8hZx/k3QeIqPQ
cR/PKogOLZ7mwzpvYkrJt1xs1grPYYYWVQP8FA1O/8PD7thHezODVgFPwSIKEfPwq2vUBNHcZgB1
i15ZC9V/ttV2ao8pNE4CIfb2GRsySRvQ435F8nVhWv4hMX3KhJLpxeEzh2scP9fOucLHMxqytlqv
sPmV+bw0gRH9ibBhckhlIOnq/dv25pvZFs8+yl5ovc5TNGGJXWvQHZnmsUtCKVzi24mw40fA2Cyp
/OdCqi0U4qqVY1oTCGioLLdM53tztvCB+T2RpXLiwYtHJiAp5fMPUWy62JYhxkAgqEUP44TP5r/P
CH0agqqyuch8XyHI3iikw8GZKsDoAPC0csypxthBq7gHm1O2g7Glrf23VERgnNEeeb3ibi7la5lK
gLjqMRijuG51DHy9fEHAWhPb21pmNH+Ha9/MC4/qH0NHOE0yEYUP+zYrDiHCrXHRoBkUVDzq0MjW
3qvEe9IzG6JZeFLpxWE9NEMfZBcu3vYHbivfK1uwGTbiPyFA43wbj2LFsDAyj/dOGDwozsoDpEiO
chH7NK5fMDIijy+nHpZtS/E6/KYNa9NNS5Y/ts8ocbiKy+uIPebasgD7P+8HjA70R3wVVBC/x/wR
wAsAWFLrOLRZMGo0f+yiRZ0HGv9AaLqTYJkx/lN52XjkBNgBSwnPoYkBcMJ+7OLsLT2iouYenPjK
WF4yStdom1DKTOvEP9rETyB4J8xEB/d7Vi3HPQPONb+PldImF8GtTkPjR7kgavJxOCIlv78u/yJp
Ayuz4O0O2JrpSZ1X92KxpNdS+DwGq9KedPIpPG+I1U4nZV661qA7dTv3pxeg2tpUkRGcXxallVUL
8UCXrZwpDz29Vv4WMowYhEwUdfxCxQCwVb5aZ7ZWO7BUk+1l03u6/zwp3K1XVq+NtjSOae3Oo27r
RTJPKRJx3K2SuKtq18BJndcaRpJNbp6JFe/DRAZUWuTLmOe6VDlXERozonRR2wcybB62el03plr7
ezm54pqSRON77GAqoAAl/MzoY6y9kE/K+1xrOhrSCnbLlEFtTWEk7efmBc880aSaVHatg4bssrwd
sh0/wWjKp5KbjQGL2QSRjhRC675cHB91AWXZ/krrbqJCFPWT0uyXKaHUCaE2pHYR9NwgZnwnrLaP
6CdIYs9BRgZXYfM6NjhetX0TXXgDVhK6txzufSprVhjg2/7tLK63fk2n+NLPR9EXqti52kFwiPTC
I5Gw2cPt4SrvYOuUdVC+tYBaf4tmfSIxvYsfPM23quT2KJ961iu/YsR408fztHDjgV8JuIThTYUB
xdq7HTrAbuiCD8j1hv7pEKATsgQUetWsBMeahI2iv6h/NE6KfRUCDiiXYMEXvYrEoB7lLU5zri4S
tyxQkQPTFydMmfXS+rgBjmY/xGpu7pFoEiC9OxRo9TA+bSa6WRcmv7lRs1tFIYwRhoLlPwFosJ9d
hig/Q42XX6M9IJ402p12BtxdWsCf/+q8Rg4ySJCpCfq/P95qYaI62HU2hvwPhdOLBexgmoE8PT/h
5G1VopUYbXKbexknLkqo2F6h/awpBl5MwiSc+7UaxBBhoP4hxmfnl0c1sBagQu7YhWmj/OEu4Yoh
dnhKviKOlGmTzitM3qWn73oG45ALPyQ5e813fIC/9m3orDyea89qOJcZ/E951lzAoJA3VGZDEQyN
yoKPHkcptwv4vv42lHAdmIfKAHWZmxvWz0nbl4xHPSvC4TTXTJb44jIU9xImovoeZUKvKuNyVk2K
l9a/pbCfWSfFHnzqYs1WJwZflQN0qUZ2WAq1WHdLxQs90VGPBLrdH6q2EMKMXKnVE5huNVBonJ4U
Uxp0Z1XIsKtZXBPE2roBk//dxft9rDk8+FNdRUxpfAP0s52ZCv8K8OBK/aWj5Q0Il5CIznH21H8+
0gXTqWIrTLto8e6guvcpfyxJqhdhxzHZ5ZhghILMehF216sa/EF0dR285Wp/VPd+efqvTJAWVE6I
HJIpHJZ3D/olouZznVTTFHhviXe1wjUDRj2YZOAODIMfmKhAjZyjCZWpTbtEOBL4vwNUkqNn/IEe
KLUmHHSmmlpDOEjO9U98kr3HK6+2tfhlyFtaGxWkPDh4xnUDY8oPxTEvTlkT/0iCur93B72KzVqg
tLEteHEcHK8ynkpQCbCZ3rZWs8m1+POhjasSJAXKsl7kLUWrZf4cbZNDeZekmBaZ1c6ip6EBseJa
2rls3GHrz41dugit6qiyOvNKRuR7w8loqMwpXHPWyT6OKfa+XY9f3LVYjahpvTk3E7HNrL4XfamD
+rV77tLHO04a7ggD6HxuppummzrQPUx/m64wS6qUUfEDkL2gPYAmxl3ol5MgnxQ27oSdmEewnJyX
lxcBebZUg3s6ZKvDQDh9VVZEZs3//vjeaZo9R3II+/8ZlJTiHHo6YjgYnjO+Jes/bxarimn9zeTu
Jgcx1kx6k+7OpyrpCs3m+7/kpGmdVJsJNpBfV+pr8OeRDNNpn0vT3s7t+JDg9cWcDeoW2HfJLSkc
u8MGWOoSRw0deYS14R54HVrmTspfOglh1euQkavwNom+F1Ka4MNYod7981xxNJiGwtloCOWTpS3j
ywDw3rHPG958lj9GNb97+qbbXKAapL9Vwgm0s5iDspuxfa9X6iBfHR/0b4ZvlDkU4tGlsR3RbL5R
0hnXLaJBAcTW3BdESy9HQxgmn5Cra9yXDrgj9wshBaD7DfKZCbzn6WugLwZt/4HNl4sh11YVWXFA
bFfW+J+ZQvAors7HJa1XpCVgrROeKyfraNtxPmBtPS8NscMJ4Bx2su595/Mnuvdo5PcZRkw1L7Zm
ZomjaMCY274iabE/nxutr4yz60WVaAM9o57P3h1M+4q4y8Rpt6b0RAe9pXLf696JxEondzMBDwHm
Ew9+JyFJn2cw9b1UEzUp0Op77EMdHblV4zol9wtx65lBhmttAMlaAO6WrKr44AxpyxSMcL2LJ+Iu
0f0wc14Tu+LZWmYs8QVJ8BFrDHf7ndoPVFl2B5zC/8rJ+oYJASZwVyy2WoOpIHPuEdjTp2UfWiPl
aCoaEsenKGHVU2uR3BDOB43rfJOxTwwje1X8RsAvEmIa9VSiemhHLw/vjR0G/cjva51cQMH86Dvw
TNHv+hkFM+bEwQK1mrbGI30JHoMu37cYdabFuPEksJR7G+cV2s8AFlPrY8WBuL9xGSYVw+l+hD7k
WuMdm0GuYhAEnTJjtyma+3j/40tbGqJImA4IOho3YUjrsCLlfbqjIO1jeIqO47Jw9nXzpj0drmcB
FXDlZbaNzdBP0fv4vo9cZup97cifRJ9210bMICN8wTXv+TSallDycZjRBkntAmNybOaei21ndtr5
ccYDfTYr4d5R3dm2Zsa1mgqZ0tq3TCZbbWtaim6g09CF/C5RB1ISWOJVrt5rfnwP5jzFfWL4dG3u
I95SyxAhvhp51rMxESlUskV/d2pfjQykaKit5dN7g3LCPsG9UdvYRjmTHlFan8+b8MHHWdnhB8fU
XbKu+0YdhAT13Gz/i2p+/IM6B403Mp3+VpXaLbjvOc+OwjbO8WApLhk365rE1dmC3nMO4z+zRXGd
sUrWELUw/0Q2frW2fYFVjzFBGPZMVGMTUutazPFR2kfZSwPkwZIfbcOuPm9tXY8zgP6HzEEsbZme
HYaeo05KuWVSsRrYi4V74qXowS/Wvf+ASB1q8BLuyeVJhl3gckvbBLMLPsFdZly0s7rh2O1gLphD
vU+AxbyFa55QvAtK7WeM7XNwrW7vFhz9ZzVhCpSLKunMrm2SpXBRfkDtIIgqWXoDH/vlM8Sh2D2Z
YCqC+99fAMfrafNNvS+BAE6U4NNI9V5A+N/Sjab9gl09jBhB9/QnNbZvz6rWtHCME99ZC2dvRPoX
Ouukl09J211FuYYGfpahqcmtuSSWehCyz2SnVRWnnWXoJSnaIa0HdGXG05oY7iF4Xa0sdo9KhfJM
0Q18CSED6Pa6bjS5xGKKksDKCZkHJ2aNZgpDm5nVap3r5Z+twuuwAqc39NRJaqsNg9V3qhxmJFvc
GnRQKqD24FRqD2e1R7HUFn3IGo1YVa+M9ZgBDM3M5R3ktkmsNAu7s+6MiN0hUHVnXaCLPq1MPGxN
5Efgoy7DmKYYYQ47QLmw2Ul/WgAmxtsrkdf/N3ba7IdvXdGQyosRNIWcPfAjBmjiqm6AUQQ/3rOl
gKlvmLEyiqd+6zYSweYqs2elayrFIJeAfB/mU3X9QVk9zFeSgxfE+aQj5NuJIIMvBe8NVxjpQL5A
lXr4fv14y5yr4Cv5FdvCfNnnVwcioyiHLFrVG9MqsmcwBa1mb5xpDor847vUeeqKT5500/HMQV+r
lAWhPzkcub59gCx+6S9egYDw3p2JrRmWfyJeMHZAdWDtAkq8hkC9i9ioALg0M/on4eOIhR3dOcDi
bJk3n3kTrWmpMl5QHWutXa7M6lHI3yPWSQTEqYfnR8xio+qnZmvl99kZn9nXgRI2he+eAFYfwtna
QhE/SV68QA3scnSf5r7A0oVpsYKpwKh2Pjkwe211yLb16UG1KxbLxzZLts16JFqszjXzq3Y0Z8Uo
TWMwO1S+U18YJ6HYEF3rEMfmWunpbxVj4ulz3pUdiHfYKeKezlG7yj3KQ1K6nJpZHkUzFc1e4VxW
qnV2zx5a6uqLaEK+hKN9s/hSN5x3T3dRwMatd7owi5TcLQeie2z+q0IWvdeNqjnvL5ea8L0xQqPf
T6aXaziVXSX6cYR0OHbxRpYxjtPgR5/A+yueSzMbYd5HB+mL87EQtlzSVO590bRO096lAdE44AyL
orC+ExnjhlM+7sVwr5VFFXAjae5NbTzb8ma2eTi4aR2TCGJCJBCCoqFlu9pE6gujSm26jUJLtcl+
AsHBP1OulNoGEDWXprobOMmihyGeo79mKv/JD1wlSA72AzEQ+7mDuYVjzd9AhOyP8LR9bZiPu2kJ
ycLv915n8k7LuR92kpuz/KzP1UKqqOgVPOBb/aZiWaeBayctCyj8mxl1DthGa3w1UEH1VJWHt3fe
Wsd6YiqSQQlPOBPm+vFXVWUyOWozq9IOtzPqj6pds+qpIFtQRns9TiKuLzR5GJZln+Gf3t/8Ga+j
tmcTpE85MW77rmHfkn4RPBuvSUSDLTfPPezN6PtcwzezsxM06GXiokTz+f6UgZYGEfGsuFDSq+3e
fJVm3JXGEcJV++2rxIfDlqMg5sHHhqGDIzyo87Lgy4S36td+fqwJSTjIBh8/poYSb33tT10mmqnK
QdQxOxtxyLDsvvbko8jg109lFtWgw0Hl2aiKx9ArkVb8HEOK9qPUe/sJoxH9gwcLR7RJws+NAl0S
M6rDtUBMJGeQJ8+pDjIcs7JrIoN6sCcdxB6tdVeapEzE4LnLySk9jSFHxkMFrVrZbuBWCoMp/b3j
ANNTqWXJxJ8IRr8wnq4hS1XHirJaIM24HOoOkmIeJIJJZbMqPJx1US4WUIy2OMRZHmrexwwbTteK
qBJKBofhq8Bm/vWbHpe7KQ/shfkCq3yF++BchedP1uUTZR158Jva25Tq/IHwTdcD2FRi3RJJEvU7
SqTZyO0+8n2k1Vg8LG26y7YPWXNVESo/rCTT5xdYHwY4U//eeD3svmhqUQQ9DkXpv3ZebdyxyqEP
Pka2O9rA2kjqbXKj7cBvCNc8YJmAUgJDImcg42FHYxKJgTnTz1LVpqcpaj0cDeqOPZrZrDqq+Scv
nlqVA0FHUcSzRk7954kLfyOxtUPPkrqGmvpOoVYOqUj32vjHsHVdgiEfAqyiRw7FcFOA7fGUOP3q
M3BYk03T6+QUef1iAcoO8HjG1ovu8YS/lQsbjLfAHH8+IatF2tUCLc43Vg0Ksq9mv5wYUNiZ6Ydq
RZd7BkCjdEuJP91QV8/Y7I3V2zjLgLPwKazDj31RqIF3JWzDMVu7DUIQHcQuFxEH+VypKPlmDqYN
pX2e1J9t/I6fgeR2B0NfdR4loEvDsEQg4lwdnsOaGj4aPYzmYo5rdNU3zBO4Hdr1o2MMw0tfRM/f
SDsXv+CNXBne7QYOjPDIIFDIJfB/sHI37LbfTJm+bqf12PUbpqgor3cLRiiJxGCOIe7Hi8/Nx1OT
tRbisPHzSdckwjDtJTA1qcbikqmhO1Rk2WKOfO6jT3NNWhyEy6G2zfnMwjUpEWMEsdDEjknaJ0Vn
ntDJMnS1vvJI0f+LzPlGsXtA5NTODNeXYI1Je5TIfWt28n3n4Ne2bkld5nXMAgChgxw2dXQI7zQN
2K2udM9GSonSWU9hhy5abr+rRpciBPvxBMEa+oeiTALF1fVFv9DpP9xWG6dk3TXWDBgB2fXCFJAF
qybpTQ3C+xexhvXTVlaUuuwMDuERcyd0s/u2Ak51UYiEvOWsptgkcFLH8FRZ39UycpKJXXMz39ES
6q7iUXtLvIJ+zoyEigrYhXpOeRmPoebxWFKpvsKGGEK54ffH8H2SBZ3ooOjSUft1Qhfoec5LriQK
Qa+EXWqHGvvgY4KPuCXVmpi9RG8p3JidQUK5PFoViTOwKDecbDVWQnH75MeJg/S+KzCI1FBo4w6G
eVE+KbtsZ1V4V2+/nyCqypFXTW5CjUUlxt2d8DQY2HcZvnsPkRsonoadOPrlevwUmByYYoVr8Js4
pgTpQCSkxnGR6TwmD/chXUpOJsqDsGK46p/pUd9CczvrpRbSgkWNZDvhzTj6yHAtioJMrT/dVb8x
0mZYOfRQF/MbW47TNfRt1fddZRL8F9Wh0hI7CyfLi3wTfmYkvKPpA91axfNP5BQL052Oxx71vShL
xtmt/5ztahP6pq2oBN+pTgqv/nHMDAFf7vGPL3wMxqpWPDnSq7l0o1eu5u9ABuzCf3RzGcWcHABm
Av9v2oLXvTHceFoBlOr51z+9pC5w6kjxtSJVjukhZoOycggLsYUaX9gvkxlCoGn3nPy273MzQQRK
CEMZcz14GEdPXh8rBED2z3KJTvU0BUDyv22OJH5Ddp8XAcSt7e8DBp5MTR/G6h40NsmtRQcmmUZO
ygIGB24LWqYw/qW/lqBp5Z4qSJHoeiYw/FmXyAu1DBGgv3SH9cI3JiZXpNT4fQzQcBRu8pvnyrSv
L8Uz0RUIZjXq+4Y3tFJj2Gl4rq6XCDkfea+GF63Rl4bBS2Xyf3KK/ydzV5gshVMbMzALZVIfA1Cy
SM3t4X/IbPjzj3+YS4QxBaDzUiSyRH2fZAD4TdBO2biYl81Zg4G9KFZeAJo3yOlFiUPcbGHywCsf
NrGVsil6VHk7gyLHW00udtKudKJvhELM11enxogWpgmAykOxrSdRlES4NNTrraITI0INFSdiQktY
IC0XHtPuMvJrPtFtJD59tzJ03+5Fk8ELzA7B56tDSTNMCnYZyXNNxDW1suUhS/ialq/VgOr91v2E
57apvkGM6TtpXxAbhLhF62s1FCBEGqxNjIfArqQ4xGalCtugJtvH1mzw2o5xsakjzEh13J8Kfa/5
B6EELKri/go41UZoujQsGGfm7aTiBZ4eNE2a5/AQKPqcNtYE4R/mla+oWfpbWMV8F3Z8+WiL01mn
QOkMc9S9Tf9kdx1sJpEAUsg7/GptgkQPgQCscTZnw+Ta77+fZKk41/Z/1jR/0/Bn20k+gtBJ74y2
8X2/zUmpeFeyJKK+XF3z+7xpp6RimOukU9kXLeyl+8Y47AFCMeFUmuT69BZ+OIWwWHrvFWqIurfc
iBsON4pvg998NKIMBHQEyzFaxl1ITq3B952flKl5UXjS45Jx9bQXry1R7Tn6qeRHbW06Xd5EYNMS
kHdOpLJzE836WxndiimbTZnVCqN69agnNUrm5M459HLgA7x0bJBKtf0hrIjmgsUoYYBvZ8cezjRX
oicx6TL4r6uvRZmXAzmjbhDUXEdIc7MJkf53UX1fSByPGjBDnJzOkzXIibDJd+CMj9ZzWqDPJNTK
Dy9Rl4Q490uywGkzDWo8tq8AshQSlkebdyTwhD84EaRic4SBvOZIUdE6kLVBaYFbx7kzOxwj5klX
i6fxllV1ha0yEFW94uaq5yuXvEWJtN0NKEaNZEaE+2nbfnZOWKCcG6TOeMF+h6wlNNghKJuSS1un
fT6uMrsyNIO847pwx4nBFvUL7BjNc02R2TB/YOPk8yBQ2diAk/fNli9sDz+28JhbOQa10NfxOOeQ
UHGWe7hB6bw9y8T3gtBfw0sSfROG33hc9pJJCRgPtPMB7gKQ/dPo7xp2Iif4f/Of9v/e+NeZ8umm
niisn6yz1oFf3wpsjiSjYUF78/90xRQmzDKZrIZvioTKYkZCiX8P3uD0iwxNIGXyTqg2yPkFL2iD
/Whi7DD42tIuRj51HLTOgntn8WqJAdJkoRB6Cf8EM9eUZe02O9LYQOYHUls0Aa8w6WyFFi8PZsTE
ogNlfpGlD/57Sd1h8LGMAA1Q0abtXBvkevqd2D6SAfad5UQhuMo2GoodMwXEKe0CyEzhp9E5sKqq
CsyY4GN1hUWyBKB006GqOq56NNxHmJNGCLlg09tDavWvGUCOrbcP4OesYGvKsSwRNuxi8VlGtz3l
jE7KXgG4EraG5g2+owbOzHSB7rTqWIO/BshIFf1R0sC5ct1oIOnkifKEDKYAK6NAD5swbeS+PfHH
U2bkjPffTdMnOoiEOjOp5840HJT1T4u3vQtOVbxPB84IJ0v8vMAZorxaZCNnUD5ZzQXNpaSHA7Ww
Mek/kNB7rczNFst681R7YDkickkXGP9SQ04L9pP+Up5mWa841Lqj0OvfhQq0Ovd6vK2atcQ+I1qG
gWbICjzvQcKuh1fq+zKMLOVNF5quxe3NYxleiGuFu14k+fo4Ow9heWMy4cfL7s9hjVSz0PhySFT2
/z98M02PIixCaae4OtwSiIz5Ife4Qz91OkHytYKxSN+Opcun3UVtk0CcWH/lKi7iM3jVhlmE6WjG
gUc/rZez8dRw1suvGYUoMEN5p5PEMvXg5cJvyH9hccikXF2PeL3gnrxjYUZWYNDVDcF6S3Z7/m/o
0Qt55DwDZK+zWzngYLY/6ENbgS5QDUyPiwJHSOul2SJpjpAyWDtPXebqaaAZJ9tDVIUuEtJFXYnX
WYX8nvdKfDcxCXHJusvI1UvbXa3HI8rrAMwGuA2rLZbRz7yifrhZO+t7KtHYhn2J8dW4JAb8CFNE
hehzD3eV/UCpHHy1bWv67YloTK3Muf6CmHn3XsLTZglT0ogWIWh/3H1hDBUbHKm3uOmQGe8c3ddi
Ws/tiQ+H965HNZ6zLcxd07xVxQJdcJtWErCU1gMHfpOTDbFrCYnwwk+lyFlbBqbPw+X1XBKu9vJi
lojMXBB2RM6VfJopVVOMf/A/xzl7tACt1jXtfcmy+2UQqZCQk00sQsNL/h4IAxE/LIx+vf9hPIJi
Ww/tYIB84jtp9jsbxrHfB/Ozi/khyrPphXtCvLbnJl54kcUQwY6InaYfIMOOhM/ep9EmaTrAwiLg
qgH2aNQaGyChCh2LSfrJd7IgVDf/TO7SrDUImLH01usoq5kQD1aq7X0lJG2sZGfKEhyHHNemO/P/
VSpuMJYrHJEzJLtKe5OPnzH5QciDUJL6DSB+7ZdIAA1oJvP2BSuy5x2loPFkxpqh2/Vw73w2t2l2
F2lhDhGj5MhrcyN4rF7i6kveqCltoQeYhXMqfQ+7553ztoM9crZ7uXu7KVGtk6wcfzfRKbF3OXb8
BtnTLpJMFq0YkYyN1miaJ//9PNlPGXYSgvRWQq/CHBiRd/9Nn0gaT3hPtKtRfqAQjzy/7BR+z7yU
oWJpOTAkp0TIGqv4IDmKegsu7RDsSmCFMIhpB+wWMk1jASL9e3AmDD4l2XNrZCZa6eiwbIqz6/6Q
KVWDa/YfLyuwCKqBFu/3iAmouCibxUQd80xHkHcJouwkUIlgVPVC5rT2/5bzMjuqmnmLSMdvLE70
OFeRKGu/PjZnxoUJcmSif1dt3MfOaK+sl56GhBBrrTd0L3NJbLwEcNwa+hvmy/yKbTQ5LfXudZHG
wjw4SsqycMS4auZ17gEPI2qU54G/yaoDdjHQ9yejr25vtE+ioIm3eCg2FrvjNPPK9CqTgjSoIK9g
WdN8LIvoww7HrGQNtsL86PAxvdsiZ3FinboEdKpQ3Sb4hOtBYuXzREgBBI9m3YC3ySTgKfMPg81r
CMMNngKlt0NgEMiKKWb5YA09MQ60a0hrU8lRbWG7KlZiOE2KXSVAQaBv1eZdAMjrFRQweIoJOFS7
uU8vBSc1kQS0JSGX8f1g//xiKCT93gr6YlU7dP1efj0NBT6GBdBVkElH0pcUPDIPX+X81kR0IhdF
n+KSyFMRkssE2WsSZUOLnlyk4hJHi8plnl212Vd27lNGUBHYKlYatW5Jz7MZdompU6MWpwJ/USpo
8XhRw6X0OGo8EdoKl4keqICkTqIRAgt+wdO39yauCU+pHLxKbc65QFU0mthqOELXf1PjLwsjlsek
uRWrbG3IqNQoD2FxX0GtI4EQph/IkDNRw2Bkr+ie0EwzUNrxQ1kQT0aXNVfaAFiCsB6mrXTSzAH4
DEDyWXOEIoEhm0e6HZdztUUKmuTfUYtlR4Kj7EPqDxd0xqSBEnEWKNMYc7MsIdSkFZZw3Jmr5xXG
mPHliFrqjCFie/2Cuawr8n+Tq/CbSzJPB+NEzQ15C9ls0EaWvyY0QCu3bAwvhEnltgPNWXRDI7Ll
KZjkr6yvJHo9HkxT1kliVRHkLEJVhbzNK3/CS3GFaqrPTlW54lra9t8I2gwC9eXgsqdMOUUsauHr
JBoEsUt6NGPhrsw9FUIT5yVzy7w0HWtI8H8vIuZ/X/ArVhl9S/lRrZ8sCfh0M4JdiMBsYUCYSXaD
w7i69VNcSXfKnYcgccnzp1de2kIOk/C9auydswPtDowjGzWJ2Ha3vzOm6OQzHWtoyrNFyZ6ITL3E
4K1mvZPEqzHgv9KTBAPERinVz6hEvmn7jacf8f43NgcxKj9KzG2p4eQd9HH0Dkp/uZPlFBNuTThx
7EAgU6L4fKa5ffISRmVvhfshL18Nvn+spdhLGfMHrmTE4wnudw9hc3dIKXTCR3WniuCsnBsOz+Nh
TzJhGdxUMGI4HuATqK70xAe3cBk+d0O6+peyDAmF7bstH/+tMC7fyJa3Qlsnl66z2p1kFYWUEThj
gVs4UiTX+6vxxvN0A3gY7rmN0Dswb6/k38nDk/9IZe6FffcI4tSGeEfQSXy/XiHoD5O5Rnk8Dk8r
XNOykJQmk5p/4Oh31+cjo5AD1Eb2YBoq5m6hDM4snJJj/N0gV0YYEtfxVleDu/0hMV27yp34vL67
Mn7VRJJxvLDDlWacyg4cRoxtxXxUK4Y2cwEhqxpa6z/qMYk79zNk99d7ZMz3Q8/qMuh2yFAw31uN
So0QUIpnI0pexeTja1y7ttvzO2D0Y+YezhG21oKRrv87hFO0DlTEE5I5sOWZyYWBMpKYL10MZkd+
rY6jDfE1IUp1lSASXgexN0v67ocEn4a8Mf8E/6DngyBSKzl1p3YBlPMDko1MAMlHVWnH6skhfdwk
+zsocFLx57RCqvzBTqZfqXqvPfI+m5VkLmnfNVRQe7O2+bnRI0NyFaqANjWGeX5Xn6EyrBMxbFHX
ZYv6MQ16EOYhRVgYswuVk9kkL9fUXmjWnaQOsv85DF6WDSWcVjBSjVKFLlbxzHJrdbz6hmn3IH0q
zTzDXRbhLtIa3d4G4B1J6h0H/9Z1xjR67Z/IW9xNH7+flTVVV+52A5m6Da3AzHRVMi7skXvKupau
x/uto72/I/0nilQvCivzGgthMjKEj8a1/laMzR6Ra/w1niH/j95thjy7Y0mxEU5f7/tyOSRc21oO
bANaqAS6A1MnaQy3KM0cEMQX2hfYlNbO/Y5iFWZDFBUJb27/eWZLlJUGFujmZHubLU8ITwQvGEte
GIvIpG3bQ+Y9srK79aqpE8mqnRpAsBhtt9cKexnEOiFMDSPBatwWZqAECs6L0fbFTEArx4Wjz2Ee
s0JdMaoR/HP4XLdQUmetQuIeaD7umi4yak5smv9riv/CKRw+8abeENumpgmUwYuxlfPdItynMs1i
W2wxajuMXK0+PR2/K1UWcwQjQenpwPBuxEta6S8zxv2+8K/QlkgC5FP50RwWwi8SOsuScTxO7eJQ
6l9ziR8CVkgTorb6f/voB3v3C7gVY47TnxbM6FquQ3gfBEk/FAbrwielAuaOApF3CweuoqlQIRQh
3u4HEWqQXWp3W0PP8tkKYzp6Pvnq+J/2G8NDQx7asBX+dRqXA8NwDPCLSm1N5v0MYgx/T4HvfpD6
TczTmwjvggpYgDO/LMNUgqNlg32r26z32Q19Vb3SeRo/fzIRtPUtBlMofPiYHTipwvN3LnRKBE0+
msBnHShhtDAIeL3fE8twn+vAYQYuX7uPYGwOv262AJMgaETt4DAKiqQhZW8vtuV8KlqYqeiv9y5M
Dw1q8wvI120VhvEMcAB76WEP7Dn7/XXkdpk8diEu2YOQ2+xoAjcw0DTcM88wiv3vqGBQkU3L9sbF
0LCp5FEipkQmQ79xSkPkdpulmS9neO+0iqUcpRRtB37RFaaM90APGRRR8hSj4qSpZTzNBV9H9P5m
cMyU3MGi4SQUWa/h9Ion7lpaRlEZOlZbYU+x87uWMhMQegy06ji61l6LNWKy8xkO1KCo6Mab7O5U
v4IAoh/34OBNkemKkz144B6KaLdK90D0QdjctoovbotHR3CBTygwTV7F+Glzx+gOeeox3AHpDCFX
APKg9AmJbfGhWgWzHFIWdZaCWqCWIYXUSncmYdlMBrlosvLDXQ1w3RMZ122NbzNhWwlDF61AkXUh
qRuhhB1nClN/rBlNVI++XtnDNEoq8T9ulcdL7ETZTQRfIy8Ozid4WDW213ANrFvHFYCvJ5bnImHE
YW6q75tn/9jJPgrhjM4ZXnKc2NxbI2p1o79TpxvX4cm4X07gMcKp0Fhhs8ybpByIKiyei3MQ5MaI
+VXIQvglyQeCeTJeWxCmSV1Bt8ura+PTqmdu+f4vNooqauGl7bWk/JgpzClBPBFiB+bU3hDOEkLY
TVuyFX5aVM/Bx6b22l+aWhu8GeP0N6JUMr9sMuX9c5JUNppK1Jl1+ceoRTpdcaDq5+TgSBzyCZYM
0rEWNos9dQcOjhgU1F1lFfUssHerHSxpstt4sM9cDuDFCSNI20kDgFkyhcsKJJwlam4KCioFGy50
7TCHwPtqMF5ZfZrNq0O3v2irTngs6u2JQOwXm9hoO/DkuOvbG4Tia3/pme9/np9/Heqh+Q3xULPc
ILK7Im2MZc/sgsF0+mB2NcRvMFxaDI23f4kRJ/VTuXG2IyRkYXmJlDYCOl4ww6+yVQq4hLQK8Flf
QnSlynjz+Nw8PP1jgbaQpShGeoaDKKQpCwsv1Agd9teUi3OB/0UG7CEyL/d4M94vejZJNN7AGi/H
8HS33U4QKxLSVxl2RALZ+rIQcTN+sda4HlIuqxGsZF/oFcCk+7RR3PU46NtbIerIlfQy1lO5VUiu
eWkIMdDESc4Ljo4dw0onsoGDFqKPt782ZEaHpcDUdeL5KIV8X17ZWQqiXXGWiqFeZ8G1veolb4aW
6NZDz5cHZKnAmirdSON2Tqwn4WJ1xY8UKxMrAJeNuGSQxAaBRgLUxykA+CZq/asoyw9rT4e2SThw
xE476O5JAvZaqaP3mAZKqPZ3jGQlM+Rzaw05K1whMTsiP7odUn2gSM7AhCgDWXcQ7QkcyrSrXfHd
36pRy061UKD3I6ENvpKZKMJ6aVbLl84vosb53eQKKwt6znTHX0uKJDaSdhd+iXE/i6zKvQjyXivC
/WaKQIv6rN1Afxr+ijhxik0cTgN6pNeaNlXVIJMo2K6jZv755lBwv1L4HHx3CLr4HIPA+NO9ZSlk
3+wLLpJ/muSTiw7oM1Y0xyjEwjuBqn3Kc8CdheefwNpRV9QwUDwQuvoUNdnr4ZpVNb9CH0A9mNjp
PHRa+C7lnNmm3fPGHPguMdMfBQ+1mB2bY+uxdtDwPpdWLvrp5pndl3YBGp4ZrjemmDLUBzGE0NSU
SAgegykU1ER05lE00xN7unEKsxSDwkQ1xLrDq8a/KVvyU7EWtkBqqbbjNwZk353oOoI9bbnzjCOe
RQHyBTdeiGpt9LUyDMesnB0szc8t61FaoLm30tAgtTus2jqujxPvAdROPiPeRPQmHIPJgviHDPOg
+PYbScf7nbsi1MTK/xTPD5Y5a99ySAIDDhRMm5Pya31ObEiieV3HpEf8asIC3ANYZaEXMHHaX5cp
EU7R8ZAuv55T3KElyXloD8EmC7Pys7aY4upJqqcaMHpVQlwN3odnF7JbP1m3SamLZlsd5UhCD+Wm
HTF7UQE/9ybOz95R0vIaOKq0LxoOxzlZaEsFJ+RASec5bLOD5KI+roIl327UQfPN5Baq/WW+0nvu
jOTyzkSjK2QQnnI1Uyyao9LVM8Iy/4ycLyjXlwsUtXEPz+tAQ/Rxg0EChvn1tKkx53u7J3ec0wGW
JEKUbVpcZoWVi2HedZWgZo1OUztbn24jPdxt0YoQ7wmD/SjuMS5V7sEwlwwVhzYhJw5Nf0/sqdot
1qoLhHHzljP0RlJ9r5OteadV3LkiqlL+N+pY28Zrn/eKTqpIN5CZLODRYKryXXu5zqIaaHt9h8Tm
Hc4dn5skhdFbBHKTB4Ty0GXwZg9JErJ1h56Fq/K2D+A27luHgAjkLMJBSlGBYfx2UR7Ns9IMlav3
sZkgLn3S1JPvSPMeC8xQEkDFoe0gtD8NBf9W7mq9ayuIlcWnmjIoyE51zDw4+KZ5lmqYGSDBLMn+
VJ98mBAeHEXL+ks8Thq+t2NTIXnHNDrhODygYNYclgUXnWAwGnca0rvx2NWJL8WQFXNFqjGx58qM
uEUjUEOJ9k8OjvrEJzPk2sHjvFForlSlQ0vSldXfT7JiEj9fIJD+c8Ds+HDiu7opc84CMN7ADMEP
6KOb4Aysa33MRz9KdwHxi0femqurhHjvkSk4MQuo0Oa/Hs1ecyWtoT7DHdWM2R8Um1W3qT87LyMq
r8Nbdi408AuRK+lk5z0z3bmKRaJ0AxlJ7p0vvc921ARDfX10W+mfE2I58MFz4IfTh0qbYH6pcYtw
RgZORjSlavyxOks451Toiq66TEG/1ogKdJhdW41fCrRHcLXVg7xHJXvBl4VS+ANfdyjebhq1HtQe
QuqtVf1+MycefLCP+xRWdEHApgRSL7gZejrhqxrl96ZfwEAPzTHxgZh9LIbsa2fS7j+iPVTk4NAB
iqhld7eL165HFC2M4xTW1013zSMgSEjhONcO4G24X55ZFEavWV/GoKUTx/ZzTimpNgz90imY/nql
kHIen5z7qCsV+wQ9yM9ldqi7S9dnNQfu9Qfs0CRKTQ1WJf5ZUQeYTayH0qTe5Yfv7bGDthWWEOfr
TqjW6gizvKVNJCrqSBE97ZoLc8JZSYzhG2uY3FJ8s7kW1rgjRioqhr2xJk/Jj2U2lOZ0p2eo6QTR
ahGTwO18WUhkrW8CYKqkLqLQiZzlqo+YlwnI+OvSjpld+LKgobrpCA1dYrcNMwTRE8OQdAvH+Gpw
Y73JKGqyNyEzRNY30mqqFMaLyeISLsS9A167arOHkb5Ug0jQUVYrehabIlI16HnxC7wf/zcnbRJv
jfjDutCu2k6zeXEdDPWtXvdhjIQ6DDunlo2r+Z0RfLoQ5CoqN6rBFthyh+GaR7bWRcXtQujq/j6R
KLhXN4KQtbwduq4E+xAFRW7ZDMpvjApMbsh/bilBB2jUppPbzYeBeZncF1UYw05OjJVgs8cMKmCn
AV4N4rtt0/hQSSzaE4KcAqibOKF97+FxA1VyYY2Aj8pKEK/2cMpgoZD9C1y6wQJmTvRVMx8vZAuU
2VYDiIs7ylFo8w3VB0QUtomb+GXpoOy+jPS9HQb6/rb33Q3IBXTeH3gq4n71KcTJ0y+AYQ/CAv6+
I2YrVx2IRZdVoO0SbSIWJF9Kg8hCQ/gkyduPypnH0n+tszolNKDMNpXIAX/7eLD2wfAxy+U++GNV
iopv7MseqPHvfY9DpAxLV/Oy/WtoVw+50WM+sJu40kedg4G81o1llGw5r3l1uUc6W+vitEPAPR1s
+2ZSaH1RIjDMM/FpN7cDkGbhZpMD/iOa95yPwwO2r9CeyJORdVb/vJVUFW29MAAC3HCTHbq7xE5o
4gUiBw8GjJnIdyc61gD0XFpz0/UM6eYDtpfpAqZfG5YW8NTjRqjj0m5/9+Gvp59bMaAAD24cCxPZ
EH8WEzUzl0WGQSgkaM0JgkSWNi3L4W/Ih7rGOuMPJPCi1Td784+1cBF6L2zBNYXBKji3vwoe9cd+
mTOL05SDKx3jnOpP0BYt5bhLhMAl+uSxi6E+YO1NLgV1WAjmxtuu60ocn0m798IWc1U3KemsKjqE
6C1ym18BjrPpaxEGQL1zQtyKC+ZM3yj/z/RLeZeBdF7C4gq92+Qg271WtVum+GmLZqCf6N+QdzuJ
OlUunltbR1BHqvq24/M6tERvyft5imL3nRls0w8kVL5o3yl5afwS2BSY8WsogkuKTCkQbcuQEIvz
ViIBkEv+QnLUUI5zOortpIXa+JPBq/LM3LpT6Ll3GOmuiMZAkfA7gZuAaoPSOPZh2tyD87uLdeuU
JXUPETBHTaud+g1XYl/9/rBa/A19Qc/dMKSXZwcbQVF9tAtsL1DfGbf47U/HWJF5P/fe1rxuSZjn
+tVQ9+24zBID71xtK3iCySldNWcOG113oL/F1wmy1RXlqROe1tm0HmjUZqGxMyV7UKJG23Nc83q0
/1CiBeaXnu4QXxSW6QEgzcyX2HYxiLFqoFlm5CKrET+8S7sFeq+PD1VngAFNC8oVMUHdiCEOdmCH
IphC2+R3TIP8gM4237bHkpeLi6jSb6VCCosvfQpAVtFlVBdUTOQRboncNOhEqsdwO4KH09m5YM50
5e/62Mo0lHYb+oFdD41B8O8XKDZ6thJeVnE8ESQpc79e177G1NxbRhd3F5viYdD9g7K0aN7tNwRv
nOA+hKwvWylBR9Psc4QVE6IWNYZK3FWESjNV4E9CJ0RSech/yEEn9j+L+Q+nMYUc25S8nJ+HOLor
qAZarXiGiDCpO2XjH6py/x6gLLsDhF6bI+J7sDUxzgDsbJnifkc1p5IQTEdXPiB5mz4RfKQQt4bk
y9GntKmB4HTlfeGlKVH7XOSdhG1G/+CtkYWIiNQCO+8lN391b+UeghXYyR/T52UrCoaRXOsYUPg5
Ij8wExSIG7P0Nt11HBO0rG0bfrAWTeNed0gYKVqkD+sYe71jsqBoWWjYzVru6CvT/n/oJwgd/y/K
rrze3mM4pzMoTAySmmxBXjhhY+DQ2LtV4oCR1fPz9IYZuPBB3b/KSIumcM9y5/mANTn0pttUK/qZ
GyYr2mFINNUqBIpXb8FNFW/F9vfN9eIq07P6K3vI09URjvVbOYl1uIRBegpx0T9pRYqse91THPkw
hnkCowJ6Rm7E4ItjjPGLR3ANgY1WMkdOTtcafwCIgWnt7LJ+44qt8lR/wYgFfJ09g7YR7fGJnLwp
rr1GmY8X9iqsg6iae7aTpx2YsZ+3V/knU0w5uIVjb5C5/16Mf9odAOKkhzUgTBM9N9AAWs8wLcC1
+Z3qtcaqrdMW0FbNCg+qKSPAx9LecVAe8BQW2A2O7ZTpQUfakdrD/ib5i8yoc/ywoEfUaT0P9OdZ
r9tLJOZc/jK2FD5vnKxs2tWPtIem6KBdLVzw7HdCt17widxkijmFbl6vwZdl7PMVXGUvf6n7zUP+
aI0R4tRFvsOwRyQrZ1dmiG2pQZVKivDFQLvW0WcLO9rinKn42CHuGACUb2m+alK2ItpSgzOXFIeZ
tx2qSfpLrLW1SPe62SPJ6ZMBd0Zq0dJgV1pwfRVRyQTM3wwE3Z/sh9tQjhVPxzZdQ+PgFc4VkGKN
SDLpczMjQFDtoxcfndzCP870doIxjETLQ9LmwdJbwSqiLkDh/ayRjJMhVoBaBnOOR7RL+/z/m6wA
RanHK7vH+Z1hTORHinv75883kIkNf5UxqE4f5oq9ghQSgNi2k/koBMONJcbe/YDEaYN7ljcCe9hl
nFA+m2R4P6fyvSODSwoHuLLs5cR0j1a6TQxdEbhYy8gC2U7SxPiSDpJg4ZcFaJTHUo+nmehXcDqZ
dxABt2Adl90JHoAJ8/DhQ6uMutkLFeiqRGfWvifCdC7LXN3b8q54MMlcP3wr1V7XMPSlD7mFRbIq
pnmce1wb4CaM+TjcjYYE1qMxjKUEI4G81uvjL/4HOdx2jbTvzWq8RFKOoD8DlpVQePolrwHOLzpg
0oDLR+UQ2NN1/Zia8m5+Ooc+vkmU9Px6bpweygMAHyQG6yH2lh6XdbYAV6/4IsTKhLV3Qf/UmBY3
Nm9e4QXM3ha9R9volSZFEybQVX0fZtRXEYxBqaEaK0akGYT5j0SIdGTl6goGb6XOmjmlb41yIwda
7AxJwrTgAulojipIDCs+2PQ0ne46EtRmUYmUl/O7ApuLb7w5027vOcfNZWx7233/p1LVe1JtI7Qw
CU/5OKbGzj5w4VH3Hc0Q+TGXBYntk6ULeZ3/Vfq5jAfESOq5NiQCg5p0bZWj3J4Qpf8Xu4iPYTfr
xq+YIUBSt78FVHbONK1S41Y0ewdj7gjtauUg2ghWFcfnbGcSe9YuRgREW0E02qTSCJdjN8hlT5AL
sWMBz4DShehYN5hs/LLaxsI1ip4RMrER2r71zXlys8n/XNuriaWrfXNPoYmzw47u4N31G5D6aFvw
z2SjaDQIHCv+G0JqFS4FozUqtJVxrtGL3DJS5vy7ub6K1Eviv+MqfQswx9HmVlhjP66p019fCtTC
vUxP0L4SfTNJtTds/Ed/91pG+pbHjdVjNW1GqG7niRoOV3o/bVMLPs+1xjFEaakD3QEhxmYzzEjH
nP60tzyKvn2Qqz84AiplxipPZ6tidi2YYXMM4yqJmocYH+XD89bKohCvNgRXrzWeF3N0GsUk4Lol
Y/2JTArwuJZMuRtrDzyYfppyh+gNAFoHB92cKlOzQTAohGWq769Mzm4t+Kp3kDihZtizzEmK7vRK
0fxiEvGg57IA4vAjK5+H5WiZz3Y0l7qbLDFtASzb9ycuKr7A8GikEiU2ZwDKlzUFzcHz4waJ25qp
o3JCoaQeGoKg6grb1WQMeZBeXfLvfPKRBYt8wnHxtwmT7eubF5jk/3iTc//rJAaCll1Kwa7J7IhI
s84autx1GDubtKAindABT1GDVPk+I4wA4Sy7fOP1ZC8I4Ti6OpNf4JFRMYV9nSLIH1tS6J2EVbky
AoQ1Ve55uR7hbNq/ISs2nJo8fVZtEETs6D4pSVbfZFkvsg6FgqdUmqhheoV0TmMnGVrccMIEB0tF
DR1/AxieZJPwIFAjLKd6jeoHU7kWGW36rKMS824/ZBoCRn5T33nb+NsBgzhgRoUxd6M4nqw4p8GL
jGkNKGpLrCAPC0+Y2X/y9qsikeJkuPSlupfuox+JcdfZVrR78oM0fcG2JRXmG/ZKEvqFNLumg/vJ
jE+r6dBrxGef/0k2clBAExDdB0yu6+I9MDax3J3LEuMedvzGpjIfNwzXDU1NdRXXEUHR6z7MRp24
kauvrcNLlp89mex7ZGyD/Z6786II4kT/z6ofSS1+o6dN78v5yE0om5H1QAl4MQNBwurKUgChcsF4
yLN+cwv8Q2MpGBSt0t3q0eeFmJ3OXDMuwFZbAi11fG5dOJeuYvfmNitfGqTLrpV2DDgY4VHosXmP
t1Y83DBDVIKOsL2uCw+EoT2euI31IONY3cZE9MYL1jcmU+cPXwty6JXxcfliqT0lWY2oUUbqLhzr
Q4+LIogyBbWlpnRrf9srAt9sfSHln7H6w76M6zQDDFVDZfmgIfx+WCCyLiVcZgNqvfgjZ4LFc5+E
cr5BaoiSP/NivFSKG50WE2l85SFihP73UfIaqpeK/mfftZtMMUcbG0zQe4qB9OU+nTsac0wkYk/J
Po7ioNQrM97pxiTvZYmEQPqDCxEEyO0nNSSnzqwcEOCsuhzuKRfNr+goFJS48/5XD1/Q7ctmOdRE
8xOM9y/1GKpdhvdGMsQLCWqtTHw1HHWR9ma+6bF5utBPYZ2Rkx2q6ODnLc+nEWP/CSf6ShJfv8sc
xSSSk9V/OVm6zyk6mpw1olqFwSq+8r82TMBttqN5QiLTyotBb9IlCdIVvRFnCt4wDljy3rDLp0+H
Aa4clSabab8kbCScRWcLpEnl94jBdL1qAAbeh8JgFyLp06EwDrP5D3Oji51YQLTQlFRbRn5ghuSc
gjWXX76YzeqR97uGVQI7EgIiDhvV6i/3p0Sz1pKEq2Ef5bGgf3eaSLXyrv6HXvNH8RxY1Cbqyd6W
zhMOSdMkfEYgbk/ZaK3R+oSyaPQjbIET8dev/JiDyrEo9C6zHddVmpr4SOAI9yBMJchMU+mY47RL
LU5Y81vWRgaXfb2C0Djz21ZrpNRqwOa2voh+4eaIDEKnt3rFlum8ZPfzH53ikBxWsua0gCsA06q6
CG8etRaQyPVBAYpASGWT2+6K/P6fyR0klYahGNmwSF57KwmLHe5xayeomvG0RaS8puLzsE0t7AhC
JqTCfyrNbWCiJA3GU88PerDFiBTlyJFCa7LkLEnO5kxS28vHGHTJJrHgy8SHvVyFjF9KmbfoKrVN
XfvK/jbfftjpq1xS1I2VLJKrKkbJp5Xy0t9uBRdbnIxNRt0n7YlJeFe4kO496LicfwOY0hvqv+Wn
CoICiFRfVctf92xw9AqwZv+mrVrlu0jFAL/llPOqqYYX5hmXArdsjp9UHp0aPJFv8llNf0df9Brs
6FMYPrPBZKkdkDGJWBTuozThzn6pgAGslCOCelStkjssmtTLFdbN+tkdVubC14PR3/Xiu4rrMdgT
u8Q5FGG7z95fMeVqh9QrnpRjn/ES7oBj2nlrBUdl8fsZyQRQ3QxhaMe55g3XmwpYkaHd3qalnYpw
E4Lx9cUJGJ2lOQmO55FIwUIlGi5uxrWBH/d9dwYGeJvjx1GBLawbGxUiiSOWufSWpnuGIhqfs1ZN
3p53UWe4bSCqYaydJpuazGemq+D3br3qnHaotF4Kp3PnINUvC/BsTnW6OAiiM18fOLHQ7bUE/7Dc
VA50hGZGWnYtIVbOD2ec8w+CM6y3Y6evxLXl5tKNuVQJEk0Ad03gNonrmzJviTOZDqm9AeQDMmNF
v/WKAaFR9E6irRAoAR1TZmeVeDLtOp/9SyYnMgaV01S1nyhUIYg9iNR0mAoPJR69prsvuJzuV3kT
cboin8H304d8MZrOkf32ZOQ1Bk2/+eGxgQgwBGNfvygkdOMPdu+lEbNMeDRKtpDYJ2nfhda9GMPn
A93CPeUi1rvSzU+sB8MSOPr8KPCOFN6yl8rd9SjkdOpkT+QbWAn9ALthEKRKxqVcUl4QXbWo2WBo
QrprJeXzeHNn6EfZGElhzYJpQIMQRnPe64x+epUq1cZCUaF1itgNiyNMwkVxWsb66Hg8HckE51Mp
CVq77OprSbMcvSbftQXwt74hDySURFhNQCTs4PxavfskhnPsM+M/wKFu85FLQE1vA+/ycueRTty0
BFFvh3/egi5yvcoWhee/CY659bWokLUY2vdZvkZwWLAfeKeGmNlPn9Lu/QcnFGEICTlqr2bUGqu5
9PR5OV+fKB3AAqFV/QLBZ2asuAXLg2BmYi3/cO1MYlKQM1X2obkbC4gEk6eD3bVW+KLlvumcBD2n
aPkgNL6P6x20e6X54qDFOd5LMOZgJXC1tUcc49Z49bWIkUaF7sOliImsK7RLNEySqp0cYwz2Ksbp
MUUACyl/ihyhFDpV0RbhWzWLvw5C9SdlJUb3iFiJzRBJmGkVpk9zRlzXCYMlT2uAc5BpQXjx0YLc
7i6Ct0R+oX5ZIuCcjZfNZXi5Jn/3aXtjzfbbp7jnp7RYvwPUwFkwvJTV50Q4JkiHS3zJYUJLRu48
POZD0TPOQx39hXetsd/A96Cxzzg7PfaJRw8uQlWIlJYjtlbIxzw7yW/8HQ8Cnb70Tdf8k9FcXCGd
yQ70QTWAJJYmqLojXlR/8NZMHkNtbE2oIJPj3XmI+UBPzGMvCKo9Nuk8B2EOAJ+RDNtmht4hWVDW
LfccJxyB+7sGkzXhvQotm3VXKMnNAzV/mfEpzYbC6KcudI1o0+fHGrf9WF6Ikf42W07o9DGvVV1f
U9pNsV8yVG4OgD2kn3GSM2RfMd80+ooCQOvXQGCd9hREKVVJUPGx6NF5U+eRMTe5nOSzqR2TqTsA
uBQsn1sbGjuTBchrpEYYLTq3OkFthUMstdfXWaRXZxicqhL1y3mKmy7kx+PrDIUe+K0ovPCRh5V2
29ofnWXBSr4T91E4PtYKVZan1g9CoWLW+yXDyAmjBpVG5iHwMEROBUBxKSJ7dJdVuj09OK+Kye0A
g47s3jHPcojfSWF6A6XFqSkyU+wXhbb0DO4ZyZ1pep6ZwV+wN+cJTA7M8SPxWzaTRm3FN51Ffbe6
rIWZRVpSnLJKSn+PGV2243n7M2gosMP+EF0qlsEidWPZ6Oo2sqMzBhJAmDdwQrPmd9sGZ2a7VCeQ
MvZLfuGIgdEYoQnZZOax5w0GhmLswgCvZ688BIlwQPannccS/XjBoBEwrwSnr54ulbmn15dMnBkv
Ksnkf+v89EupFZEGS7FmKuCo7jGzv4wptH9HJBrhNfDa9I4G84q/G6N9UgPXF4KoRjRsTEGGzoAq
T6Xoc3Ev2WnDJArrtcyH1zVUYD3aA0EfdV1+GUx+TkuDFaE/weHYlNfMEt8mgOo+0REk2RFfNqRj
UBGNzei9F63NB55MFnEBVNEW1Nc1ri5pUh9jYcqdY46usOTcyBHE6oHIHdw69kybik3BAYrKMp3I
VC+lo/tfM21dC3s2WAxuxVtPfL1FiBv+h8qPqs0fiyktRqPOuN21hTu/OyLHFAIatLgGm7pybHXW
QAKUlhCeQXnGVNZUMDVYr5VUzF1qk2Qz2he839JaXZB+qjPQSL4y08FRK7b+plWrN6pYlVqXyeKF
mb4y5qVWvVuqCy7B+mNokvsNWLiY520K/O+Ox1iPHwkyQkPqBjphb4mtSUzPAZZ9flH3aRL7HS5N
5LIU1ghZlh043VcCSsoAcuVeoD2BzP8G+PAbRjJK8JYi4YzbV1Ryme0Nbd3MJDfWkunNOg1QLWBM
Ci6RW7/lFfWiNC5qCC5lBNO5wX4xC2OZnFAfi9iwRWcWSS/rtCDOc2sH2tmK6N9MOUe5q8oVrjaF
vcMkzM+xlYoSWLTint7AWh4A1QXW7mGQPTkzOyeW4NGUU19ti8n90gVPkaMxyezH2bJC2TMSgMqn
yHhOs+Xx9hbBsrfPdRNX2qafx6r7ITrWpQPxfonMx57Pc0iTSaPYBVcmBnZhI168y+kE+uqVBWxx
nOXQs0WVYKYxrh45mwm/dHkQa96DH3ZaiAkTakCh7y0Dqd/LsOF4B5OXFTZJVmV+iubVjQDGQIuy
7bmyNNsjTHDSyOhoJ22Ots8WGHM1BBEeoDRzzt2k+QoEyQJ9Ey6J7T4nzZBpE5m15Z5IxoBIwoN6
Jp/FwAUJx1Mt7VZlgXhJCUvCGlPqEalekZvRVh3DPsHLh2L6r8CuUFiLVkPJ1c+iu48oFQrPR5aX
ysRVoAZ086+AH/nariAzatyi8Mvc4qRli//BlbQmWdkkxYMB4iIMSHoe7gY0Njza83RwhT1WICyA
F1TyaBbJnMje+qVE+jIZEk8VyZG4zyLeE4HUOhqYZPbl+1FXAYUY4/xoqbuLZC4xNGU2tyE7TWxM
dUrntWQBnJLYM4NwAra8TQ0zAh4gOGPNy5KTTR1k1XhKIbaJiHxmHIZ9hwBpsq03QRAK6ML8CmAs
ZHv5pc7Fp8srWyHXt6urQ4/KWk1IXNC3Xgr4kwY9A94lo6Mkl0CYMMFvuv0t7RyKYzT0uxOsFChB
DCKqlCrPHwEdEqsMvgMrpm5AYbHQyDWx9oUvMjOIJ/HyT2zqay0aELnwoFhv9o3ivE2/KCKyF1BJ
E1emf7BE7QFyWJD5EEfpSM7h/UBZ1Er9/5z3aBi4KF8FYLS9A6bmWcfp4NutqRi8O6IX7CXX2o+g
1xUC49Vgfb6eSZoBW/a8rUzGy+Cbpu0F5VZM73EQIljdTBVUSIbnwbeOiTzLUHpAlECbFygk+331
QU3iAwGN3Rfc2cscWmPT9y++XmwmfJlgJexZdCmZayFAWcUaOLXn5UAc5DsduCuEVj/yf8A1zoAU
B9Q6Rq7Bx75PmnAVvW9YlNj9FeoqStmJ4U2rfH6+hh6FmMCZ74QOO4aKWNONSv97Rc2PrVaO9P+b
8YYvVyubm7rAByqNoKvh8FwwElGVnHOMnFImV0zN3rGw+mMTVwmuFf2uCos0IZGRjr3chIa3rMcX
ESR8iNdDnp6aAT/F03aFKxdAYdo85NEdGpM1R2ckd/qw8hUF/DUf/4ldsM1w0qhPlZY6LTVpHO8G
faaMturlLfIcVer4Lc6iMewDdRcdX4Mzu83j0t25nP47fUCnw44/MDITQX3uyS0vnPwFKA1rtWlp
P4FafRNeXILLcWGH2852ZkF7MbajgwfFVRw6kk8jOSUnZqbdRNHYnOr97RvaZYFAoFkhc7Q6LBGH
U/sZGLiFY3CYErfevw+sZAkHymmlq0dR8XqdGSORvWvsmAWQh2U/cYKgvIk0i9uJoErh4Ww7P5Aj
zaegnxNceXO+2UUYo2bNqNc/VjyxWOZV1uetmpSKFZ3E1lA3sHesvRUAqPborUnmJJ1hCuiFs/V6
iVy0uVm6Z52E4nNbm2TJAqDwHOmqmAr/HR2NtgTcl9BwjepeQdzXdKN4/xQBH6tIHMMCY6xkg/nr
Uw2mL2mHovfRRyxKLFUxLDBk48CL6ZaCIDyRTch0HNrnAytFrA6nbqFfGzNm95h9VG2x7uqgEprj
AxIpgSpwMnMKIF/N+bv+CSWnPUdHqHWqMk0atduUK8ukPHRF1X/Pz5xejc3E6Gryhvix/S7Lhufj
m6Wk+0/FKacwnrCJMEDGzf5CyeLxT7gMWVqd7999xov4ZJrzf5J2uHohVv1sK1NbmDOPIapaS5sH
gNiA+YkV5JM0bVT/TGE/xnAo//yuSIUFlLWXmLi7p1EvK86e6/MFMcigjQAgFNKWYUtKwrfAZlW+
BbRUX0FQ1Oeqx3Y7YcvHeChGAHmKSCQvQ1Ztl2wM2PhVLtq28p4VAeEwYCBrF1HV3jcA63byeiPJ
AOsKaOsFi+ZzAwxYzsA3liFkZf9ojSg2dSoKP+hyi4AGtbk4r0in+s6ZDMeMmFNYf3QzWaGfTyU5
jMqGzLIGgPN6d897PoMHuRXL/cgdbHpjBjB7n1o1vX2lRKhatzWNiGW9T9XnLiA+B0U+hH9FDgB2
t4yZvWKOUzBo98fdIaxyk91tNSz/HA8nbO1VfRZP/63HTlDZt5jLtbLo4tPYRqQx1yYQkKVYR+uA
GMgmJ65cKA/S9/orS+L51snebo0SDDJ8aKU0HHcnYnHSmCeOOIiYi4TWRU3tywIuKd3NOoYr0Uei
97QyumCPZ/qXJNUgu42QdfTqiq8xo9I/pSy4K0mTvu0yKdmJb0M3CXuEFAUTJaiOKt+VpTOmsB6l
LG5Xn4nngRMIVrot8BpzKV+J/ixNM3S9+K0FM4mdsYSO7lU+R3g9xp0pqUN/eBuTN2HYEVRJDTHc
+IBLtf283s7CmZI7hhk4we54pM7MmSqV3h2GRCcOu6MOFgM2PcHsTaZck92um+S3pFLTigAW5FWq
hqAI8A8YMUxBkHwag5QtaqXN4aAAZGVNqD7Trc1S3Y3diAMPPaguOfOPIQ==
`pragma protect end_protected

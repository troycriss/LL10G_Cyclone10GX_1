// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
Bkb2cu7YbdFmDQjUYIO9+yYBJyP0sMRezjWXxkO+VVlOr1ktDiFj6O3D//rm89NAehRBzeY64rQw
AZlU+YWeN1ad+g4hPkvlqH+thRzymA4ugpBdcLg4juoJyzN3cVn6yuavPfJQWwFqDhJ0P3jFQKX5
fHFf7xRY31zCDu+ob4wpdoHodZDlRKueArQ9mOGNFTQrk7dqjEMvLmKiwHP7XcHRmmgd4ElUmXaQ
kxMDaGBRRBS1AYqsqenLXLAHyA0jrsSOw8gcXYehEfOU6H96hf6AyHGdEsuuHTPr3/hU3XNBWkVY
W05Uwv3yh2GnRAxdgOU2ChPwEyxb0tXxxYsIWA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 11456)
9BQJvTN8vkgtBHiKKtk40uwcP64WrjCGFs9BpwbhiemwNpkrw963E/M9SOZkOjkpgn+yCcBHmTQ4
Asj2TlLBfAuLyQL2z/Md5XCt24m90thd8mYOWHQLjkQzF2YDlJTQ9M8xnU5DWShDAIUGZP6rhCN/
S1J0yOL4H3tV8otwaACOlBIgQUuh4mdxoQFvNyBiANU7lXA0D4f8aF+fNhnD0C8/rG6Ap6TC30hp
aYcd7QmZQPr6THv9fP5yoSgzV2VTqAomdPzk5ZElzgbwe9Yt2PW4Xcmx/D8yOL/athSOFnHhd6Ph
HYd5CrmViwkLF3MUy3rv5LrHjsWASVb6AYl5rUL/HwS5Zv6nMgqmTeblqIE3AaBPaIZPS1yGs/Ws
jYS8eIm4QNZSdL6WDYpS+ru9OVE9BqgAnCZk8A1ZW8kpzREjbOmxLvYw9pjhjgkmXwg1VfKwSgZS
F6Q3WuLdCJM8Uyf4NuyRLVkElAP0JfLwonvJgZyiEgv3XSXPXy/w5UdcXddmg/dJOfiGG9KItiCm
J6T0RuD+NDaZnwKIVxfBvKAhbWDUzivVDtxUXDBDs3pLbeB5hLNg7Fk9Ghye6iTaqT3h/Lez54av
um10RQFXTwFRm1HjYiSQ2yzg6G8N+C8Mko9w6qu0kY/GHZaft0Yd0GZImWLNSMTy1Nkygksy9uk3
gS8j1jZv/Emf9JHkyfWYjPpkh0EPh9r9Yh5F3iW9MxJqYkn4qffihmF6EOlnwcatAgUlbU55a63S
0rSg2l3NXwpVqZUQySGklb/Rh9sKzsJS1RyOBSPAP0nk2adznfCX8rvmNyFjKyaYGURL2zxtvCJU
99w5gMMo2PipbyFr4ZgotE5GxTs9qtBg7CR1zRXFVBxIFcEp/AcS9mR1IQ//zOdeA1YMnadaoLKn
w6pEaz+qRKlCcaunKH/pHKUZVhVYOJ5CF+oSefMUZoEJLT7AWY7a9BKKex4BjHA/smlnd4pYdtr7
mIDfSQFGKizru6gaYFfGr5NHxSvv8lhD5L1dLswb7tm6JoBgaQ4tB4Clo+5I5pYD5cf0sN3lVGR2
NtbrrTtnpaizrH4aoJymu+HkAC2x8HaNzCdJtGj/MWdUiJWt7Tjb06PV7WSDvZ52rb1G3DOGy8JQ
HBMGRQrQ2fE8IRHruZ/KMQxQWpA1tdlhMOvx5wjXfZWc2/9Pr23ql2IbjfKGte/7mzHH8IIdI9Gz
gHRi4gHmhtxfYFWu3ZsFZ0grb3fgqLqTLIcrtvqZUJHwpnk0hT9Nx2PDMrFA0uxChxhBakIvvnt+
dRYkPk0RnZYFISLbnVVhF71fIy/Z5d8kjS0D3hUUq+oLlRQ3nsANOAmyuacM1lBqi9f5AJXO3+cA
Wy+w0GXv1zWHrVPWllfOsCZVwwM/DzdLC74xZS+GWGj0uEU8/NXanRuXL/bDwu6ZP4K2FbNgZs1y
nFv3xnFln04lVfEQdJ7M2wqc7jUhXbEWZQ5/2bTHJJrdk/G79reLBDAsj/eBNu4qRVHs4akVN3C5
RBv7dt8HkWmjnzi5OpiIYHxWq/G7ocVhbxRiYHxwUJ1U51417Zzdwj9bhHaIdlO8nKa0PuLbAj0b
2YCwAsO07yJ6hwJZyDO9syulVb0IYEAQpYZBW6CFObNSuy7WkxTKSBVET9FpNpSGtyS5fJY5tnHi
Wx+xeTP9I5W8l9LY6RxIgkeAL63POyy9p3oMu1pHGcSUshV8y8W4VR56oOgTUe+sBHCExCg48bGs
c6tQjwLPUoVesT7UEVdH+wqnxFqFyEieIP3DfE0QX/XVti3Yj6Jo1/46ea3KW+KMOu1ng9/sgK23
0UOjRq7lWKcyIQXsrPYkhMudIZsMAKY9W8b+9lu6Gl0jIyyevLfPd2huegQCHO1gdpykJHjKke9d
JSZxoCPLlY8LSZOJwOdMLft4lBA30/kG1lNz5xfznRmnFVl9xEkgSb7nXwhifciPp9u17A8BVwes
NilMlh8LPbUk8Dxk2dbIxTxQzoCyCWGVB2Arr8hnWNKcF/Ton8PSlZbmlkZR4rhJBpqYTm+bqBE5
YDVBTSPrC70VcNga2Yz/xd3UZTjA/rQ6U72EKbeRmDB9Q1OULN/eyFJoi8QSIT+5PWCvEHAUCfXq
j/Qq7jvUpqtBDBkrWjjuETvpz5f7ecIeftLrUAXyVO59j9j8dwxg6ecIS+TS9aTZ/tCYomcpxAR6
9rEleHXbnB8T+50xg/ihaXNaQ8SL1yBn8kWmfT0+CEBgxDvcPqymrYhjzqLGZ8JVW5CyYMyxQFuo
BUaYIlwvBMXFfwxzgudwCBMS10L3079RA6uHjNr7XDBJawSOXgfQOAitXQjrzjsU+khILWYKpeie
9s25DTAwfeK4u67XBR7KZlLI7bjbaQ7WZmyC05PVKWvfICW7PMH93oQE5LmTNxrSaghSxozam9Zl
Tq0WYhlwxmKcF/KC3/1O+f/w4xOrqjlJf7d6sUv9y9w1h+QWopuN7dfIH8d0Zb46x4o+/44ojEiA
E70OZFQhcuWmMC5vn3oK2H9qf4HmyOMMDS7WNhTDTLFL+FK39mVVDy/gzKFGhaVITx1vKHq2sLVL
s/3GDz/6ivLGeQCB2e7K295SnvVVWiTL+YwgtKj5kYqVpFEljgaZAbLAyV82LmF5fEw7BygDjLrs
9dEg80syehFhioZf24uu8qhZtExgZSl/0Wog6DtjdptWbb254fKpRwpfpFjeZEdZkage4voZKqXv
+WLZy9iTXBNr+51tMJnN94LGnGpvM/ccBHlaVKDNuq+RKNwJ4srJJJ+wVulRX7s+y2hf+BSpy12e
v3glbAn5+rcTIoelZ40GMHNSysE+rzbYNL0FED3unuBLQkocDvE//CN7A8eWGKUfp8fdAJNfAYhQ
l5k4rVVpvp379jzuWAQCbCU2x4nLFmQgZqcZ3nMtNx4uwVJ48iqSKvON/dMW4IB9DKgIPWaJ08a9
pMZ7oUSFj+yipXbrxfOECZiQ1BOHNnXDa7MWtulmtuPamj2827Hs1PUzBh8RE7zBlr6OTPTugJb/
dPrkXjDygwKVebA5vsqlJpoNC7nsICU5KRsUrZsfZdWVtsPBw35XLnk9XA9fbTWx1HY/JVDtIk0D
Jk69OyEYYveAfML+cHyMW2V2LiuxYIMCkMCROrgJRHxOeoGJcADqWnj4h1p19BhRjuDLFshMh8hn
t54Pk1cZhGbTC1NN26WjPHKeay9FyHgOv7GeqglcrdAUITrTQDpOkdhk7L8KgwO06ait7sWhYIZ2
+7P73zE3DyT3tzDxQK4m0A8e5ivJnpp78nWXe4krn7aEI+29Kw5kwtrhIGCJk1nO5SRDaI1uB2pY
HAGHAu/qBYmEDOuavI/6wymvMYeER3CF4fRH1g6tx4d1F1klti7YkiyQQZ3gcUHIgl9U1ZcDdxnV
1SmSj/H+ROFfiJ8z6+JI15y3U630in8wa8+ei+Rbnzyi1lj+ZBaz1s78YlMIQD8/sfr5cRh6EvWj
slyM4qeVXciME5nZhxG2Zlzuqlj9FUy9UiwsGoPgZIgz3fcUWVxkryMY7eyWthThuEfeBLAsT8JJ
Z42ViXT4zL9wFC9Z0dko++bhgaN6Xn+Sb7j9SCq4+BN0T0bA/E6C6KXHQoUfoq8aSSfRH981n9gJ
hmhPYi0f9ruK8obiu4w3xfZ8iTs9WNCSPAvH9r+mVvnwVtSjuFQRjFmVWg+3UtcGqnGjoKfwKYTz
xutey35TmbCW6J0uH7hRoC9ScZOglqOim7rZrjFmw20CH9VC0tIYIClHcJcBehxHsZETQsnpxBLx
pul8LASEh4BKpU1Wzu+aCBo+mAD+bttmb2m+4I6jfBqS+IkMFw6tcRMTANGV7SB7RHVLE21/NIaF
rbwjTQMsrQgTPNrpaYMuxcTcTLAYWUp3kPXXyBZ0/1VvR54NSgIdHdpZswRuvCK11sveIuyh9NcK
5lVlUDZmmfyeBXSosDzkbl6PKrvqt1HN+05rxFWFO/6nGNCOjymIV7wM+JPWbRkP4uDe9smJZbTN
e4+IKVuXFBr7edZGz2AIzgWS58+UidY4qHmA+PpSLNHVMxf+Yub43Zxbbie1rrexiCUlSIsapH/B
VCH9Ls/ZS46PU7wiN0a6o8haC8j0uikhN7kz4xoCsGGorLekE4m6ErSfAf/K1xjy3DMNpa3T2TWP
BNmdfo3aH6XgrQ7nmXul1bi/axozPDkKtlS07L71ZbE9bC8evAbgeiORX3nHK6SdT+Yf5C21Ug9x
ioyU3OdRncQqMCmY+PCq6ABs/dgf2/ztts/raojp4BwhMBr2QngGTDWv+DAVdf2qKEt6lToUW5FK
sjnFPzgRpK/N+SV+XApTqc3t3K/2U5p6gY56Y8kWQJxYhroOihQU+Sq4+BuR4Jbl3Alf2396Y2DR
e1mzTrQi6a5dIHv+uSmkvtDo+ygIHfYeMQGj9pxt8ImZXIM8tVg4OBkMZb1LcXT/962AxLBcdchy
D+CZioCqjTCgzoWGTHFoxG2Z5zoSap84VBUjkFkNLYZDCxb7cPisa3Tkk5mI4kpUvFuoBra3N13X
qbN1WBXfGiLvo7++vPKvZ+4vTcUPmF8TByBst+kWTHBbIuo+PStUuXNO1FxOVJp+fSL7ogxa3fgo
t2cU6cHZI21J6Dn+K789PO6vjrzFRaXfVM9hsWk4bqUDemS9hOa5UlbEI0TyH2HGuRYA5Coyiqlm
MG4BxpjuFq+lBtVK8jraEo3/uOqkpE+87z3m2IJTg3qc6FpwXyWjSxGa7xN+siDmCZmU0Da/YaLR
zCUq6yB/M9oQ1iAk8QIQajUN9qCNbSwE7V9TNkNVJW9DKV2XHz/yQzJnhWe8vFW6rrcHtLZQgNIC
6OkexJnmfNBKZp/TxgmPImtFvgCTpW6HcPyMs/QVTKEPL1QfUNfUZYJsoWQnkptMeE9GSG9SfW6M
NXyyGt08wlqVpqkwjJHWDqttHBIyLJTreM8/SnnfIlE/6zBGO3OID9smKQMAkhypcmznQHBTma/M
K9GSSH+hMdw7A58k1DIVMEnFndqIUcx65Wrf44+xwqZU2p9sitJg/TVLl22JmKqCrUr4bUl8d5p8
/aCP+Cmk/Ol9aFQMh0ZJB8AnHcLQYrg62dWJdpawkJxBrk8pt+AuuHVHUFfnas69NuYxkdM2L4EQ
1O72W34U3jU0Hov0kwztGjOuoJuTG1Gi3UCVfVJxTR43uFjtedPa4081DnTQMvm/SAuEM8XUXJ+e
i+nQ5rJVC269nrVmh+952wNu7PALCi/8U6U2gKeJceuOGSqSBC/2vEYvOivn4eJ0ENxnWf1EPNpY
GTROsSB0kE3f6j8mXD0gG+NulcUuRLK6373uaUIhkfAjuEJWF7gVnTLsNznszjmLyYTMnnb+Cob2
GLRwAM8fkSUf8w9C3XBtAd9bzpx2BOn36dMFQ1/6TRLwk1oiQ3Hgg5vJRiASYrqpufZ4P8L79XfR
LPGFzUWTUD7FZcPIkhPln3X/yMayQT6/0ORnnM+lQXkn34640wVdEOfKnOf42rxwwEjTRBrS03g5
U2lyx22cjpAxBUjQTCuoPds67UIU0GUBMwPiY2pAVFPcexZjIi2//XOgZYE3usG2ZPRMDtHXtFln
Dx5ljK5iZE4BlkNTPoKOgbpxHgoUNtqrLoJf9R5GZ0e1JOPfi2ZMJm9MtCsIaZTvbFIk5oyQPnsf
dQ566hP01w4IshnvpeJjjGA06Nn9x5KasYoPJYNumqx8PoR4PlAM3od3APllVRxWen7Bxap7qORt
IMtbr3TGAcyxn4w1TYsP1XZuEqe5/0MDzNzglL2KVO2CsG+bYyqWOhmjyHDskiOP4sBqNoRuLVx4
dImRDqluIWkAZIpT1PZ46CKDLHsqXP6QsSs24YX9OyqlQM37zOvLgPtX/TA8FuScsKBZ226vIA1Y
GfCBsWnBYOBqbYiuDIKpSjiD4iuIzDOHDG/N0xQpw52T7YUhG2i0dLdvKl1ST6op9V5m/PdhFi9T
g4Aku50e5WKZ38HxgO/LvdzOfIpXk5MDa7/ge8v6PR6tK01PL5TeZVw8xReasknUpyOngI0PNOlL
KRZuEIcLXF/BYTUkgqTfcWzNmd3SphZ93ZZpUt5kZIWiWF9jWRkNE0HbXuyej52kDIOPys0H/L4d
19BZHD89rTwYw51hdMtBv2pSDmDp3yTlCnpGt4mqW08OAoVLK9l3BkihqztdjAh1Trz1+/KoidS4
JbrDNJv9/vr4hICj/wTzUlGuxkOglIFX9StAqVnpVtpDrHDn6jtMYclTa+fkdulL86xCo/M0YubO
6uN2mwuHu1qws7kBnHUtLKIyhdVevYQJctJTGTzvX87qrDlU0zyrvqCo0hxCdjWbvIVQXdGxSgc3
M7ZayO3Q61VDs2b4HBy/dl9RYQQFXocTHMM5NIcbl7GTjaaRkc0UtMcv9q+j28Xv0luEOemwY43M
wwp2y3fw62jdx1HoLT0q3eFv41ZTygUZaLCLne7MToZAWUZc9yLBfKVKJpkZISgRPtXyYuRg7Aqy
wHP0uyNdzysGvsEJTg+va8O6yy+M5g7XKTJASKQDdbretfRANKcYhQeGAIOyisro6jhPomtTGT2W
m1wbg+vVRATvjuIcF5nV9u41hxciDM57wPVIhy9RinSTHHMiKgeP7jFFL5T7QLgBCTy7HSktH7Y6
Ej9bADzag6/f4STt/nIKa5nJzC4/Nj0yIfZWZEMUsSQVv8MdumuGK9lyssFhW/+rtUvrLctk1tz1
5jp4PV7RzTOSkHHSPp4nXgEMTLL/aZHCw/CiQbO3twEmsRg0AyrvwdEEnFsHoFJt+zFD6qTJCe7u
/k0eH+6RefrAylR5ZmGGsRiL/CNeLwR6vmxa3RUzPOXOmSTFiQKtqJBe7mOKylujftMBOg1dOlDT
p9Br2pV18HqUQIbKU+yLKy1HxwRfOQd3eKSxwvTo36C1YThiYN2ioBM/VCojsNqYYK/r/Q0Hnqfy
URqAYSAVSi44qP1BarsauFdrwkH3RMw9N+LNVSMPdVLCMDK1qGTSA1mPRAIwm4tgdN3bsMU3uOQd
Rz+CbtaXFZYADgtbWaA2gPzeMhB6q87BF/yUWPBNnY8ZMaOBAw328607+CrX4qnP6DtRs3CwxC21
Dh5NVhosGcqcNCD2iXuSx8VVxn4F6LU7fMwRPKk93EQ6lsABFKim8Up+xbfCpPa9WY3PvGu3vEJS
8cKU8cpVMAaMVj552T1AzMES02OCqjWWw+2jkbrTm9ocWjsQpZKecLc6ECwY/rTy/dgTcd1N7CFP
HWKZBODrdBFe52/W22/7Jy6/w1HVQYGbz9xkUffudTHdt9ADrrIqy+fKdw/3p3TZPrdcqKrO6nOu
x/sa6SgKNiLrmEEJbqm5R8OjwNpwM3BP4r8S94E79IQtC6efqiLHsBDroTSAiCBNN69ofnF7Dl8Y
G57LvyX4GcaV25oFEinKlG9Ojw0aLzvDMR88mOSMI4MPQPLR3YgUafgRDClV5j3ncqdaIAwiWQ/2
PfpqhpZ6MXJoowmToODLx15xJ5NLDSPQcWdc207RvhJqx57MWAuMwlXbpyDeWfnMnXNVKJSFnsk2
fzPpu5G0HBxaXm2MvxUqwTU5cgWFe9/WI2ugaaFmPKMh7LDCviO0nGz6NnH/LciLNjInpDD1WHYE
aKPfmqVMpmZrYVM2LQq5M2HD45Tuwis+SPp1H7618TlCHqsLd5Zz4UuBdIRFp56HKoqr0NT+R8DP
BRFszZMqvMleB9UQDoeHL9RdyppwsLUYkgJQSo/fWOk1vqRzkdh3tG4i+NANQf8ZpcZcuRvJyFmM
Dmyy9IgWY9Edfy39Gl9qCB1HMsh8SKGZUF5QLaM4RLyMsSsGMimv+MUWZo6S0KxirhhoF6hYf4pM
oduyVMQTaTIQycHiUX3AefqKk8Umwq1Y3G8o7ckf8ysxje3FNwgYggHQctHw86+Kxz9eoIX/QdBt
aTv3cMsHaG4VTXG8ouOX3Q+7j0eeouMqaTZQMtJqjrFdv+hUJvBZ9zDY9LpL1D00EklXqEnCiK9R
B7TUoen3BkBwDaCZ6GFGCu6PkvvADI7A03tvOB26U3TAlSskrPrEHzqB9RFrSjkROvOJmmOcDtAf
tPiyQEiBosVeAHZFJisTjNcNqJTKf7w1o9wnxKeBSZ2Fe0PhSO4PhUhrBSlEjP3xPnhhE7vLODV4
TfQE+dk9q5Mfi9fFGFTrkxn/XnQuAPFZtI12rOZF3ab3DM6Whpk6qyoEFYBJAbff0E9oEfkxREnc
l/pXsY1XiKt5L0lVq0Q2LlOxTYil6pSoICDnCuu2tbe3IeAjeDo8vuDPl7EXjLStwGmMWZOfGNlG
+Po3WbepkOquW6sQ3HxQCbmS/6x+bt0fhXcmwMrzhWFiC6fqyTzY2qBw4bk/oVxsmvRjo18/pIbH
cOoaPFtu/gr1xTqpf0Eyn8V/ut24u+yRp6r1gxtWEFhc0tCP0GHai8VLs6YNRW7tkGN1bS7SZ1gO
3ly1itD+andlhUT1a/joCnCgXqeIhfBkoZ2BxvqtpcU40UlTUDXmnakWplls/7e7MhDvPLeQDo0W
NnlYVd7gqT9AYR7OL3F9i7/C2rZ63a25pteH/IvDv9VJFU8o8xL468XDROCsQNC+YUDPMf8zx42m
+IeH4hOezROF13CXBi+5oJ1f/CGYgsDAUL0j0ND4M89jdgGifwRq1bb6FYDG+TtdAdHCHbMz/38b
9QAGs8UDjc/4FG6k0fYcQrz663Pnj4FiCZHtmGUU5mzcVedsNAan6ZRu0/gy6Ilyu/kssG+WfJXo
8j78sePgXfc9Wqu+NY2Aq67TePXt7TB/ejAxdn2rC4cwptfCY4KGyjwub1AU2u3857jrtDW98Dfb
LMWgkolM9ldE9b2klu0+thG9meXHRAMggGOdsOEy0xsQCRfMsqDD65CnOozleO0CfzDbLGYRXASh
mxJWfEwf1FJdeKoyWtorugIbKCci2/Y8AFgdy5T45zXb+2ffYpzpjZqX9ZJqftYRff/W7EWfPBbi
kEj3J7jL1Xs3DeWxlfVvmgqsTd+7kMw7Q+XV7AtmBZtsi3tjifw6tLO+F3DRYHVGMu2XQkmdLnr3
mTr+w9z1g1s/FcwIT7XbW1S7GvP9pXM2mo2K+Fh599HHVhVkwW6SJf9gRW5ZDOOba3Bx8h1LjMQC
FNJ4gRI5gSiW8NaQ0nrw3GeDozVjhj1juNetv6ZscgRzrT3J4XxU2YLWxqqzyYrodhyODVb7EsWv
KVLMVjrPpQvRBVcfDj6Q51VQFRk+jxaDtDGOTwT0zdI18On5ANB3ZoNxG7RS6BO+IVtyhasRLAl6
UUeRfpNmh1/vqYzfEC2mYgTqhAva6AMZdqUtbDfPTxeUy06eFEOeaTXyaU+s3mMaR8wY9DABko5a
RDy5vObhCtod956t/iGTKz93t4AUlk4A0rhSLurlUtOfaGoHEom2qnfVE1upW1k4neDEAmgP/x43
OglT+CpCLXkmhBsogiahVqqtU5rJfiuaFyR8ZXk9HQKthr7JcYqFosxz9VCDavkEW6W1k/lkBw2V
zAxjr9hQL8QiYnJOZ6OP8MOM4NhTTGB4xXNvTj+dEIaRqcyU8D7V4RqafsK9N9fwWFr6lW3I6e6v
kkFvXjpldfMdRR9yV5zQI12drpCY2y6Byb92+rsW9BDbryBVCR0lPwu2lqqKiSgGrPlQeZ2PMqtr
RTms3YkqMFXPdAuRf9CLKM9dDqnJ5Gh7kU809ctv5pIoHJZFG95N7lYg+4Bv2HBvEnX4Crc6Nkbe
ghfm8ITAogTxfSqTyAcGaisfzay5uZsDG+7OX6j++qrrdQ4wTWqTrUy3XBOwsHKcb1/IoydQyas9
VAIHH4z1uPZUUMY7iKEJEWTJqFy5nNiULPdje2odTnghKr6iZ8Gvah4cyegC+Kw38MghAmDqtMcF
UlCOJ6yd/KQ8/wcPOgaIEAWZ015UcRqxb4PAjytqyM1rcGItO+v6mCssq7teOW/dPlE4rzdMXOEm
aIV9A2awHWfrGeDMdxsk+asfLjrbNzqYQKtWyMYTOwSBgYu6QRjf9lrtVG9rm4jO/wjK096A13um
EMtkqarxdMB/oAk0PBNpZPo7QJvQELeLHGRXZdoi14L9xpmV31olI1RA+tWkm4G0RqyfSnHorc+l
dgJET/WFSJ0OzPrDvv6pgsT9siDZmzrsSjOWkbO//1unSVVun0YNDZyVvIovZcAW9reQssfMvf86
EMTsCxDPsWfhHPJbJT9qxrN+CFbnjyTOZiubC9HWtcFdlH2cjPvpK84qv+BWUOJpN/YBlFpgApGl
rE1yN+Nhqqgby/SD3xZtQLPdxYJvSA8BVMgSCYwi8aKtJtQuNoeok0jWqJFB71zsXaNDwf8yJa7X
ZbN9vG5MreXNbzZN6sj77Kv+XfffJt5/tCpWxPpjjbKC4my/C2G/Gtw7xagmKmUlzu1IfaDfrurX
bWoRfMPIqWOU222AmkyXd5PbkjaAoV5sNtcn2760HPoAnA+CCdOyQex31vxCtHrWFcdHeq/ABrP1
kuU44Hfk22jnpxnq7Yj1qUeI0QtGSmeo/Dz+lr4+tpMUClwKgfJCDG8TZY6MrdFvtvyKmwE4qQ+q
q6VOliyh1oIhN5NjHS2zACS5c8wXBOekkm1HHBLUEw2cYNE7yfghblpwOM77ghfGDYRmsGyix4CG
9JVSFjPtb7aVYSokn6Ambyiih1jIQ2JdcYBbXfFTwFEAdClmmmLse9QEoN68QzA24MU/t31xUL0w
Lj8gGBdlwT+iEp/n75O4jW+zZx42Pxz9VInmTcj5TSA1DBS1nFmKg7CG3t7dqtNsEnsfLtiSj/Dz
HYC9Ak+NIFUTITl9Mnt/yqTXCMQ0Ke/kYAVRZ8nPMvegybm0ciA5HcPKmdi5+PoO1LDQfTbM0Dog
MeUqWMi/9KVQM15KeW3p8Y2TTApE1+eo7iKY/mpKiEYM9zDIybPmMrkCID1DOh/8ErLu5c/YdYyK
GpHrOI/dttMeCW1dZrTB5Td2UUQv/1Upeup/gbTRFxluq9kZD/zBDr0D5+b/J56/vQgdiLZY/Z2+
0KDxHEcQKhSSlX/IAn49uHgBsaRnRr0AM9J8SFIh7Zt+RT7M4Ro9aK8lWkr5qNmQpnrKPg/02hD8
rEEQgx4vYYP3x7RRcBFJ+pkxw8TUZHXiJOftv6Mk2sLaRxgvCyHsIvTUWmVNVvr051k8drJMFzoH
meoVcDfJsianK6MpneqHDQ2ACw+E3KgPpAW5I3E07FK4ea+ik7IXHbH/2xZOV2wGQ7nAs8rghO1v
/1PErfZI9QHQ7L8cN9ZAfP131o005+NCA9M1r7WrXO0lZIzHsYCl3bZs4hN1kygVeMNPHd6ACDIv
0wR5GV50zngcigc3UsgwUsT6K5m1YvpI8mzH5e/3m8x6ez/Z2ehCtmOa/u/UsAo4npVYh3Fimwhi
RlnUQsJ+/+EXQ8nS5rN6ng3o7icFs1EcdRGnlaDU8pOMWxAPcixS4bt/65bnUZD3Vi9BmDK56VOJ
9NhuvZFUeGI97NyYKHt8GVzZkl3DCBH/o3b4msV/r9wpRoLr9h0OxHT/SPPS277d/d2Yiaa5MBrf
36z67rDAEjSoqaNlMOQ2Yxwaghn0sPt3/4l3kpZNf/5sT9AUX/Iqt25rm6uNlAPOqhVHn3qpFwre
l+6AvFPIpEVUdOK6NgUOhnrCLYvPvefQqDYCI4iEec5Gv/E/Xc/PukamlvNzd8nUxzEtTZxGGCIW
2H/X+0M8iZOa4Z5cp2BtaNvJYPZQ7Mlh0YAj6aCwMaRH9hS511Ai10E0fBXRFmxlKfbpjWdFi4EP
s60adIFZpVMOKqba2zzS/yMqtyDy/FoK+Kzn3q5W/P+ftxoeod/N+Fw5dwn8O4P6nGrjt3v09zYg
3mCobybzaw909WjOM7dIe3TPkjTOI79Kbit7VCu0cMGB/g/axtYCsz1WCKgV4eLQVoCzaTNIyzjj
XTIRT0Ptjkbc7Q51jw12AtMEq+3iBqcwpFqqMU5qlrZjgyJtZ+SMxbWES12RkiQwY2AeGBga8qRu
S4abdKCcnaCebmKc1VpY8iO4N7psCAq1eLPO5C2mJRNeuD3msUJPyckBh6P1g8vjKtxxU6avhfXR
MK0SkBQOuoQ6XZqWjNs5QS5IGmpLWISK5GeEqT4OSxkulJblP6xcZAujUWg8K270E75c0L+hsHv2
r94M0NYB5P4sVL/lHKibF9B5mpWdsexTRyrTEEXUrwmWQQlTEYY7GZaaXLe15M8jr+vjHhhCaene
rmSJKZHo7IibaoIQRTzXoM6fbr5iMFm5uyNa0KvgVAzybrnBmzVut8cVzZB2/ITsNhSwFV3oYLOF
HVquqL/RpE+GAl5R8y2bQ8rY2eaWu0ZCUXixzLd1bXdDs4+UlqntMADrZ3yLty7ViWH9fxm0nwlD
aoi1cd2IgBw9ftrmqYqltSXl4XSPVwy2clUCIFYTiCb+X48B0rU7vZw3QELc7BUefqsD6IdWygdZ
e5H8Ppzls+XM3VckyMu3tNR8xPM6gghgCLr2XCEN5aJ4zXm0IAK1qMUvRxxbF++4gnTJd4rrcsZV
r+xpO8TeoKbYWXgsonwW9l7ZlKDCQfmGLKpASS/jAstch7p+PvBGJjnqXlJh8phuHEfowOO2AMKQ
l4bECptdY4qnJuE0WMawiv+4y3rE/GN3Mc7+ajaiRlzqV647ke9f2Pnt6vL0hw2dE1Ld3gpK4Wak
Ll6o5dQaIirpMCFGcIs86nSUHDUM+/Wi6yzLK5Qxlo6Xp2K+5Sb2KPhgAw/0wd4R60/sBZ+OxXvp
gXSLT+vPjQo5Ewqq0tZjvQlCDCoT32gJzvn/Jb0pTmhJ8r3J3XX2+z9ujvOvbWwVL//Fe4NLq0vD
FEL1iWIet2HnAiCxwZXa/VG2D3Bxa9fL3W1e4SNCPRVCY3Nx/kBQ6v5zzOQaKBYkFqO4SpUt3Kjw
I2TSv57zBSgvJ6eQiPVItqhVQvYTE1jM9DA3xccvK7FlSbccQ9LY3PodgxdxWqOkxI6u+rwPvHDX
wdLVTLnYHpWgAKM+K/uQIQXD21bXlwLNWDk7n+3wunc+rZ7qJOVdrSVC4b4opZfREHyFW29SVqZ+
rN6CO213130GFe6+fCbfRKnsK5AEiawsmAozKRV5o5Z/U1QHafPP2/ZqQ5gawi7lzpimnD/XKquU
FXJhEehh77wqjGy8Q08m72vdMsdSTikR+mdd2fKP8KrnQexUKHrflWCGQPPZPRYoIt2cKZy1TEJN
+/lULMvI/WiG1ywHophpjovP7h3O78EvxpXK2tvQBhvuHxzG+LvNu1UiTjroik1wyJW9+yrf3QZ7
EkQiki2ggeNM2abM2XcGiozw/Dsx5zrQSeUuYo/0cegW6rKTOyNN9sCFothqKBYPUPlUFKQ05eRT
miZO1eDPViLSiJ67LHkVP6AELxZCVKzjgsUXXkCuO2dEM90gcM/nwdS3jnBPf8GkMMFE+23H3hF0
0sJtZzvkF9kYXMC9x9M3cAqeNiNzrXRdCF3cj5pZZE2GxylzO0QlHutmkhbZzIucF5m/O26i1tcW
3v/u3DJJ9ShWAphiymwLQMBzZS2caYE4ZPKKZFA4EKF23OFdheyJ7UOEGV+EKObhUBmuNAdyUiie
35Wsa5XrkXZXJI7ac/d8CdBmj6HNoQjPUbneyK5rPZJvxcRApeJY3cFH4Ruc+ldLAhT+mYatBpRx
iMmKEg1uZyO+RNr85N+P9LI4cQ+QewpzRCFgCXPwcG1JMenBMzMiqwBoobEpcL8q7gkVc91JzYAh
V3vMUTDG1vo41XzbYdsVFgWDRst8+OolWnrObaxbMWy8GSebmE0Eqcj8N+KXyrK4tKygZwuDjzRf
hawnF+CnyIlAj40MbCoeWdD9uvzXzZ0h3MMIocYI5PBgstuOAJNazJJyNTcgCtujOPhyOSj2m8rt
m94chwBfzYPvCd99kdaDBR37pqo5u5cbgi3TEt/C/qtqYX3GdsfwevBh0muaCmrKFEPvkW3UOM6r
OtjtTwRv4Nm4AGbXkfj5SxxQ3detkcSG7UCIDol+HdpYbaadt9M4gCDGS299Wl56AUYmKMC9c7Ee
DXnAMtZFqIf/DCwyHDUGi02kEcTGyw7yDLhMwtbILWkssc0TKydMU9sH8DolJoWbCvtmc6LBrHPA
P8kIUctGKthq2+DXb6YOUVIVlXVWy1lQhJnMJwqejXLdVyl7damuDPK6HYko+xRNWt5Gu4XwmSTZ
o+Z+0htFiHwMux5S5LyNZOcncaV3iNMfzIOKE+AiurbvL8Zxg0h+SnoVaScMIZ9ti6T+cWbibgyR
gg7x1aCe6BJPbIUj3T1GSbqBdAsrRrztT2xAjRaR3+14jCeXnTEopf9N3o/QK/k8csnjwgKju3W5
XS1FVmVNSDLcWVGmCZ8W2oD34PaBlyFyDyyj+8J+Oy7JZF2rKM6PH05OljDFEnUhQXASVlFXsWSb
3/MPWlZM0uKPXjotivWlN2DfDDaV8Nh0crh0xmwILUzSsOUOLTC5ThyXgXvqBFeJlYsXsm8pfWOq
XtxDCokkjNFHDlW/lVtFtK5hnXJxbrENw8HYwX0xOPA+A3I4kBe2SHVpVCsPNh8Fg38WpBYE9KcF
cSAstx0sw1msJisKgU+k5YgyHOF8sLmYv+Y7XEb4LE+eIiIYtZMM4+ykMbkOx3AAvGwIOmCsOPvQ
lKtYhXccjm7wq4G6JlVr5JWXJyb5VVSgK3UA2IV5ZYqr+emVkUVasU2o3i13R8Ji0UNXvDmo22UC
XpRVJAWvpqM9mix0QztWxXfLZAk3vzGzXAuLor70Bw+mwKVh+s1jWngEz6FkZKf9amZ/05Gtwbbm
cufDlELz5Uhqxsbvd6JIU2RySVAB8g/bZt5QUl3EBc6P3bU7FFgYKQSgvsAZDO8qLHF4XR3FhtLI
HfVlZpFSNiCSqPhN8xMlQ1nZUYQFhlNH98ewS3eb1ksvLjWq0/eOsD+PPjHb5uAqPh+Dl7MhzC+1
FGCixW8yPxHzOxKbtjKoO6gU+e4+zJ0HGFYloE8Y621l4SUg/Mr8dfb/0+Fa0o0D7al2TK6PNlfF
LC1NSanS4B2k97RPDbmSokJqxKLqGNH+zIW5QgnBSOLj3QAP3ikkjEIBkG5yF/3h7xj+vUq6qlJh
lIiMGnYBr4t5YbKqXAN1ad2+camWii8jfL1Zz9qVEG7tCG9z8mq1DnjcvT4m5fo8zIJN3JdF5Lc=
`pragma protect end_protected

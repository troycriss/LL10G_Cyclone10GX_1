`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
KSqrVcVEOZegiWUTBPsbfeEU8A/bP3klE7Z0i3wPrCKevyAtAYj+eLsBdd9GTQxF
N3mS7fJK90yzPKnOmjzgc+ZCOSRYonM/dOpRkGgU2NDdPvD6XDKt3Ib6Qr5T+6dk
VcK1hS6I6mvLlYKDHb/sErKvZl0s2rfUoVere7mOfGE=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 19328), data_block
QYTSyXiRDUJFwpuJHHP40mVV2iPnpcesgia1GEg9Wlp6O+88JzOEs/K9nQ5ivfI2
07rcb0hquFADFiAvBGOIfxMYJrgmTB5UpdDmt5nDBXGm0Ar5yD7o8Ikgc10lHPA1
5Kz0PvjPW6eZKe3WPmXqRsBeYhecMzszNuf5pgitvjysaALTKL9nlAIf2cOPLTxd
tlW3Ttk4ZSB+fItCQ4RGMLrWy3I5qTH5XKTi5MjxMrU9kvq3QNoAcpfK31aQ7dAj
lJu6oN3aZgVeUphjz/Iz/8xcKWXItM21hmfEd+oU7PncN7G+PtI7zhYqpjSSxLLo
2mqLhzL9V/VNjItY22Rgiy80fRATttbW3XBl3dy2ovJlnBpDrucX9mcL2evPLU5W
MMBNpuamhuoCPLVago6YH9a4JzG5K2wqVAVmY/T2bSpVsYP4tQOb4UeaAcXBrtG2
0kCDwvnEJvvMtVI/3+tVubUdOt1xgw4LIs/RrBQvLTUWMUxQsSs7BlB0ASSX35yx
rZZumHb5eIfwWI9V2qveg/ks/VYnnYh2CaC0ZevqgVlSsroinn2DInS1mOzjapO+
DKKfsysSEBNYkYcw4xryt8mqdxGsogROFkKgE89gSxnvIUiMQk7/G7jD7xLZYavc
rYn9E4Hi4DWo09SNiux+iU1KgCqvDSUs5ydyDKttkFP2uKYVXe5YVoduUYvg6bkV
ANVbKGbyZWG5ej4IkgW4s6R4LnPbKKS4aBher2qTsbsm1eEWh3MzLuTB7NekqRbN
u+Ssi27PhVvLESAx6lP56OPfIJRWNyiSxjQRi1qPawKUQ3QTw0F7m5S4HIyw7Zk1
CgFtLX+e1ucGZ3/A1ge45/hrG6WC2R154TwnsaOuN7XqSMlamvyRWO/3cih+zfwe
WmyGUQe4iZYJH+VTBunSVfemX1HCzKUk2cNSwZPlL74SHCe/ZRe00xNLJ8EQdLNw
Vo3YGdLKxHFJUVRwuhs9WE3lGZEcW6GNfZsRLkaySaS3T8pMbkuF8a7G0BrvA1l0
synGlLbqmmPxezML+nEyzBOcIUgibHnXWJQif3jIyFw7aCRyKbDClWc6lxr4zkV9
jxl7Se4Ik3opcbqhvSK24X6Zjtjiyflh9qPGyOSu2WMfzCZvBbEEf59AHuJyH0aZ
wnOWx2y0ipTcXt6WYt6Jy2DSG+Bsk96+dIpn+irZXXuXr2qmuTWpAFr6+qxzZOHv
Wkm3e+xiE4neOxidmwHEuNkuDYP09RKGC3h01Gp2eoraCkhm5zSAmNhfodbNdpTg
Zjw46ZIqwPMz3Eu6/hIIo6lf+9MUMKlE+ed7zUJPA07Cg1rx6pzLb300ZM0Ny5XR
8QFFzNoX1nOcx2JX11Nb38NRwr7SfOiSGM1vjCKvUhIPvLPN+HMHJVDn+A/hXO7r
VG3ieGXtOwQ6xXi7N6l8CifFJ5ePZDUIPxys8TVEr+D/aKRypofawnqxagq5a4CZ
tdXUgP7KtQY5hGZn+RO/wR1f1XrZSk2nBgcRkGN7p55ncRUCDZSdB2mANqn804Gj
BQ9goGlicGLGGzGTwA2/fM9a/l+h/+4JjzX8X0z8ChUvbRK8F3HUUbbErToFvGkL
I1/dMrmmkuSKB7PMpsAJLlSy1DIiBFDOztqOtFlmVLwd0sISyDPcTyWk5jlIUFjI
rRe+teU3IfjgUsaDQSzqFHYK7Lc7/9nkxSVJhMcA12mpjODEZMPOXPEMrumkn+3x
bDyg+a1AE81NIi16VLwCuQAky28Z7GywPRSltSt5a/OJiKRKYomiuw25NNwXCkM7
CQnydkQGc+4Xme0xMBU9FMY4LRwVvkp4ITGB3k++eMi0yAHaBEmXy/z4C3ZiOnL2
rOHZ4PKr2LxtUzHYjiJpinnlLXt9U3fYfMudUmkwzWBNtmmpyfxdd5LGxw4aIcdy
JWaIkwDuBy+8gpe6vNWAypvXFhQqoGtNBk42PuD+Dw4PkF9CkBfN9oF5Ibr5kupF
ZW8FtTKZ8nPAid74YXH0rgFLO2Go6P9ngO/AQaqM++B57ibNiCzKPX6jcPHm4rJ9
G2fuPVdPjRT6WACkfHzBiSboDt352+4VS96+t5jxAQtVC/7N1KAxA0iuFkGOAbe0
4GAjQIZDs/0o65ug/W0YTqT+UPrTj1Ko7sTyOrqzLxwdIEZ2m1bbJeqdib2uZE6a
hm7EgS5zGte3uMaD94RIGnmeXZW35CmGJem7493r49JqE5KpzlFl2qxaLAUKkPjs
ULC/rex3OmwKG0qyRRcMSxVmY4HAbqQzeJXLvjRACqjUdt7O3fEzuDj5mUvaTg8T
VieU9N+PfbwUlRLIWtQm9g8WW7jUXsTPloUycuszwmUA75ZD0aucXVKpDsZeIM5O
uqQUMPO/EHzhMFzlaPouel0PphKl9H78pGpkOLiWuOx7WAx0PXwSXRCqSyKEhAiw
8ysC7CYI/ZdzvXk2JVoRuDPDG1V706DgYHBy1skDImf1yYCmPNNoyUP8zKqelUFU
kSAhKokZnrV+NibSQE9cihIq/CBoZPywQLEjf2dJnya5h1dqxFw6tldfOcRtb+7Z
uQeee5rvfe1gxW/wSjKHeNcHz3FZH84FVgVCXlbwt6ynWlmD/Kc7XtSQA27Kb6zO
WOjB2UrHWpz91DbsHtlnHzE8kmDRxu5Ks437XeyZm9o5Cp09cZhbEPXeB88VTnAY
hwBO0bhNneB7FtaKZw2RJ1Emya04xuc6Aqw/z3627jSfcBmS4vNi5GBT0JLzuv/n
kYPoGYqUQU5ScwvkKlMPsXegedivxiEKggn5KwyBSA4gGj2O8wsK+o31eJNAT8Tt
4cdV6bTctvZeeBve8WNJAQIzGWe/EsNrR2nIOLvsgC3z0svXhT+/0uZk/NzsFqh5
8+0EYOEdLKNnqCR9u9A6yKw8mxvtMCYeF36egKYL3//UldlpEHjfJai8U/bYrMad
vSDgliUB3skB3N1+nbfclYiOSAVTdbp1csPNCYC4/ve93PgqNZg97Zi0sRiPoNGG
100pP0dLF39ur3vzYhvS2jZk6HiJqlVOlzSo3r8CmfgE1o1hYAG7cZ+Du9O0QpEg
c4pmUkf17Yu4n8vzYW1IGXtolMl7Kck1W//oqt6iBu10m9olzzDOGp7DBmTmgH+f
KW4o8SSl0DXrnJ3ZMAiCGHatl6HZjeqd2mxsYCKQRpglsqDi3t0oav1C9SkQDuRA
jZdlxoMDU+dlPgOrs1Rh+2L0tPvnILQVW0obcZeXgmfbzHKiLVdyMxpKTxVRVb/J
Y7jB9z9f5pf3fhKs6cSSMni6mgXKZXWINaPOeeYmd5zv27pJDx6T/nJZ7uMWgFix
yZ3iKpb6j5KaoTLM5py83Tg0F4Qv6/OleHXhcXD3IbJRGj9riEuN8uGFSYEQ5beC
RsWVTXjhChYiDmW+txDhTEj9ArDIOpduZDk0PcLqNlZrywRL0Ez9PPwFBRkNdgi3
E+7LRK69dPyt0MCEdNKhKPO7QaWmbfMllYrFvieBAl0WV4dT5C3T2RWrVttf3UEZ
dhCYIXghJmtBdZCOR45Nk7Qo7mPRWW1d9jdQh0KRD4MeEtgSmTHaRe9vclntWjbD
QfKYFRdrm5+lCb+haDsLbFWQPzrzZvdDhdMYBf6BVSOPsbXVKuGEe1dN7d5yDMDe
etTUMbP+YlmMItn2GkuN02BaLpaiJltsEOmbtuimculnMR8mH87OS1WsfCD1UEPu
4qRt6+6vCP3SzIRnlmzXwNQi1HqmnN+lA7E1GEcMqhMQKMVKfce7pMi0kqO1xyoN
N1b66x3JMAdK1bEEMGtFUdKWJm3zrNbg0ptNioAQm/GYA/qzqTt7+AA6OoU7gh9r
7azxqpDfHiRnyFaA6SfwNHYYgNkY9ZxvzwRpcvK1vYCQeD3GzizRNdcjj75yxmO4
8al+1iiRia7gYMM96t4FV8cR6GJGG8diobIa4KtGQOpp9DOzrN/SHqYGD7TjN31w
9q87oFWk1MR+j2IjUD2rj/6aspPPdT0GqdxmrIm8WCHaSLqeSsrnm8Si8SpLqVII
4to2ocMcmDYpK/r9gOGwB0sV+GOp+wBt8W9hePpTGqCp02o9izjndweEF7QaWRGa
nfGmc4e3+T+mN/0H7Exqds7Ezk9hzjDif01zkkPskhKRyNBiokrJSnA3iwsKPjwR
taPDoooU/4ciD4HLnd592YM7tvOnCATWuMAKbC83dej3Ru7AJ4fVm7AWojDuM8ZT
9aLauUdJHcsl3ZclDvgPfIyRSsW0WytEa8VxRgjNHAD8bV5bPFIPidMjGkHAiWHk
B3jU6wCIrMXdTYLjP7BdjTidP6UCY1c/tZW5YPTHvjK4tepXn8BgPefDGPSTRhAi
idx6+Vjkd+uWZANozfJ+d01Ro2GJNaT1PbKaZFFwVZoTsCR7QeECjS9yTc7bRXlB
Fgg1eRRThb40fga0lVnXinq+RIo5jkHr8Z12WAcPOOUMOE2ISVGDiCiobCG1bvHa
FSYJ7/I7W6aQmFAHs+PKWAcs1tsWOlu7Uw10DctYKzJVcWFn+ffh0HGnxKcPv4AX
2p2LzpjupHskbF2KxoDpMvfrZrDzdcjIKPYkKodQ6lycpBIlWTVR6vFzdnnLV5xi
vBMkbAzDpbY7AgpJ/CEacc4pyTjYo3+qSCfo1PoZ/sRmCLduQEUS7gIzWnNecymE
pk4JHaHPskN/OZpFup+XRWQI3geN/DUXIRffRvSXY3zYwWf62hdTtmYGh27uLKKX
khAO80dBcMaAq6sYjW8B5vglvbHcFlCKIKpisqZTdzY0HfrgqTt0irOp7gMvx36d
krCpyW+mhWTBh0zdj8Qp9ylpHg4qWRtE1bUT6ELC6k9q3hs4SfIfkMXsM/5K9QnU
E8J5wQAnUWIUUSsDHJ/LNN+3l9MTXNPm65a2allpNP8I5m/TUT/bTrHzyzm6QcuG
VwfBkEPZvw+VxV52dmUVuZc849GGTT4C/vRcIegjbsCp6xyHPT3PS0aOTAbj1H+d
H/p6hKAr6q90QzGcDe8u6jGH/2ReFz6RHCtqmdhp2f3d14oh6U9CmyDr63DZybEb
kVznjrojdtcQRNBKQgpKoC3tE0bSPrzCIq56c642MKDIH+q8y3BRhG3KnqQrxcuQ
SiOGloDPW+zirWN/QALks6cg132slmGX/DkitTR0X2i+HdLaxbolG+9+CB5HLidH
LtQ1DHXtOUxrAo6rvKaHLNtufxQ/NZawRrYXWbGMJVSBzq/UL0/bNz+YUDIg2TLg
/8SJ7L17djEqbCkg7MZOhX2Ya9dlDPFtlHtYoPi9cDpbOuec1G9G4RLxOdJNKTSm
IZjr0Jxn3z2MdBj3HPHfYjUOdj2ODKXWaxB9mrj4fBAEXGNAV80nQbFUlSS097mY
RqSkTOkcD+XFEQc3zBb/Wcfsv6kitfV+MV41GEm25kZ0BK6lKZDWy4z8X0qTla7E
BoO4NTSR3UxTrnDdB+PWXKf/R4W+OZrOPXqVIoPx5ATSUhpn15BpZaClAe/D75y1
CHxXLa3hcM5bbhBg0OWl3qHoID3mrFp4S3AIFVf9wb4QoWZhMmnTii5N8YGGwE33
TsjGNoMwDUJVvJCAoum+kv7gOS2FJTd3B9NY+pnvGrT7HjAvfL8BBaA8vNf7Sx1r
pek9ujyHU4MAfIfBJ34WjFzvP/ftW58JdUOgCybwwzCcSfoe9vbOKDPZ7qq8qwqk
tiLDQq1rNCUl7hAR+TXHa1A9B5X4T+rEu6L4K1fa3uthE2CIl67bpIo49zF3Ktki
WwxhOYHof3Mj1VKyAMVEwUJm736mp1H3VqvLmdIFm/8H3JweRlKXOAp9WM+4QM7R
P5uTCyIuBYcFbXgwd+DDWtoVlpJrDEJAtpQtvK9CBBZYj15nsEBWkOkvmsg2Tr/Z
M8mgI/MTFvxwEnn2QIj+Va/Sgt9PzfrKt1+wZrpK7I4+AINrjXcOEwldeAJ0AH2L
D+Ix6cE9xSIq4LKxsklxO+bJskUrL4q66k65brRpYhh79JcwN41aZJV4om7hG76B
v2lUXv/SYLOVeJEHAYI1w2MzEHlJF8Mb5FQDWPHdCU/w2KiGhc2svbqwMIPDqM36
COSKQ3hR4vUXD82U3kCf05F1Vod25uK9TIyJnaJ9RGGKYwDXpYI2lRS31Fhi8Bf/
GmGj5rdxdtwqAJol0n01mjihPe0WKhXc2qWHvWHsLWFBPhCof2YDsivPz3hORv1a
JR/I24fQEuXFdIPQRZwEQxLCqWbtY4qdam0IKzZx1Miq53AxfnogbgcxLaIjuY5y
KYKNZN/Hlz26U/gWWssg/PhrPDHp8vYrVFqyEWDnGpdzPwuIp47XJRVal1v6cCDA
cMK2brUZMDlCWjJYBMnCBEMBjjsf0CG5oS85EJx5DXiUpzKm9uURSVRSU8sZDFp7
l76qoqUq7xenXUAxA1WxQfdrgYwqq8wQqysapfuyKJxg4m1kgmsiEfPEcncYCBkG
OhRpRzGaxFmmRlTRdrDEh4czouuU218gdkgi7dgdcdmEgzZdcH32NFaExlacUfjV
mannvCB7fcBNGznVOuUeWQehtAJ/I/w8i5n5/2FtdHy+bEcaxXAe/tPwbQdWkzNj
UctJ9HlHov2hDdXnWoZWVayCtXCO79t52joJuVAIpV2X6KG2ZapxqIvIOMgcjUds
dp+Ujj6Y+YQ4PCmlkbUHMKUkea3XdiDqvgHXfY/hI4dWqlNsA+2vsCaA9l1FdhHM
yBIdiDxfFx/VovjazSkgwdZ5YaRok+60Ff8BSbE/tAOPCRsLu9I8D6vA9JhPhXTJ
nfJaHMRWXjxzSQd8Jx+0OWXui3ruVcOPD879eJ6ZeUGFKyOlcAWjfqwQkC06rx7C
HiOcUq8uzaBzd4O99UIwPrZNZTuCUZ8K9ozmz2Mo96UO1kmMC9H+PExraW53Ggub
nT6MrB5VcMARc1nlP4N0XYyXbwcvTFJ4jsrG94Jg6TvChVAgoTwSb7qKId+55pAw
VFpZYJYkDXsvQ4b2qj6m61C0MZyQSOqp3EG2J3EWDF+0xR5CKpxrvnPrnQxlPE+p
644v6gr+t3xTio1cpNMlB6MqXtYzugBUGlq+7p3r6GN8v4c0DEpZAz5quf1Cy/QZ
sugj1cJ0EPeB4q1ONuhxuWkhLEyrmffIz9G+D15+SFyz9KYcjTIRi182CaQvFFWQ
PPYpziJMvjqjzclzqAae2EuniBrmGeqbGcrHCXrJw3tz+Fimr8E2qiVkWq0tnpV3
YMkgFMWWH1qVhOWPnRB4JuHo0tfw3YlrBFmtOIhlm8EnTnhkXf5hlIpE+7ZubACT
LlJaiWRBSE5EjKxLTVE2jS1ALZA2zSQmXgBPvRndhSlrzlHnfk1yaiccuZuxMDjf
x293HzVcLHsD82On9pVaKZClKfjVWnWumIQf71GBQo3AO366EkjUP6sntFNMnTEv
swk1ado8NIUxxammARq9F4L2cGt4KwKy+hxi3sIwRg5iN5KWdfE8HljdP7myXqM7
DUBToXa+mFtnLZs2TpunsQLgl1sq6PiPVnntAP7Tyc3h7pYFAsRCHINxZdpfct3x
XdYmsejzuiIEL5CImkHxZbrHeSPxzdETHzNglwGwhVLfW5mBt23LEpdHJdk7omW1
weX/0mW0q/4cXzJfj9mZchb4URLuSSCq8YFloi2/59wWo+RN/3kk8jf+PqL99AKg
FtCkVSJm17VEetnucLpzLJDfx/InGpVdNZKz7oF4NJp5dfXp5S0nPQXDXVahLb3z
D1noIvD4OedNhs/2R2rUGHPyUiBn8HgICxs/yl5yrVFMlXwJlX4du/N6sydd68O3
4gQ7QuwuZy45v0Mcaq6HiESnEYGZqunBhk02LIi5e1ak3ifjaVMAteXdUtQDOJfY
w7SPUNF16qOhZIFtxMAsstJGi3M7g6vo6UCqcR2smGnstsVw1hZecT7PnP4Q6PBv
sHxgS27yj+tEjBpH/mL1bpW//q3CExNB+N7tP6ABCH8KDMLVsUof30gp6Zl9FDQ5
3uDrVDedajp3pj1I+GG5NhzWmFegENjYXL9R7YHWNP7KSzztWU/XyylSYjq9djxw
6eYwP6Jj3DHfdimlD37Lx/YjkMPOKyBoy/1isEmW2m0vMam9So8HqVJ5DQf7qYjA
nf2GQMrF3a6VVXI9i1a4TAHsf87y1F/ksFkUNSHiWe3aKfPBoUxxT1Sp+JZFQoBI
Q9+7LYenQTNfYyWXI+Ih8vPvKaYkbvUKVdCZQEGORkLS6oPng1NlUX4zGJaJAiVw
uHWPPEoPA4Ep+JSo1RM4L9QHqfdeVzBVyL3xPFjMAaLvZ7QrYqZsmdEGNJIwwLNm
nCTnZ20R+f/Gki2WflwvwvRttTbQlj0Zet9bc8/62axu1WBk85ji2Ew9D+NmMF5A
Zvur6o3iLM8lbPyYnEO09F3XdMe/U1dHMCDTdtFdi1DYoi01tzaq8hnu7nFywzIa
MY8PZQx1ZC8yIm+lNMy8UoGO2hnbM8lrNxvyrgB85OzdBIBcGutUof2UgjFcRGtG
ErbwHjt1yn/Ziqw27t+gZJqzzb2ubUT2iHUf9kCKqmnB5Tzrw3QYfzw9DtALbaqd
5WJx8Tu4ltYwgQSkYaLofNMPQL2xzZdD9+doLFNoabs1iUzSLLOmY0kGRAb0dyKW
iyiey4GMw/WDaH1If1R1qIV42BwSDbHx3r1Q84tm7TXGWTYsea2cj5l2315DPM4Y
zZ5BSp3O0d9J4H804XRx5KHw7+YC2dDlUjnuAn60A5S9MBH0q7F9JhPiWHlGTnyr
u+WFb4II9KdLpP4kuMD+LigEn4o4yzQSaztHICahSo4nwYtw46qB7/0l3fFr28RD
9iBFVVAkSCSdUwRe6lOuuliKjQWE4qDIgaobyNNEaGp2aV8pnvxNB6oe+NerEMZA
vR8jkFhUtw2gO++FY3bxuQ4nMFgUYhgvhBVl34WHO/hDiFPvWE901jijZf+shQF3
T8+d9mAKnLKKdEm/NvtsxQONkR+uMCMoy3iJdIoWjfg+0K6i6tiZSP8kYwOSzUm8
sKN5TTho/Gmfle8zrv95btm+0PHFstynNir8PYCxd85k++FTb5cdb+/Vlb0Kd/nH
gPmgHGl6iMhMwMyR2AK6TP8TMABpPvbnFnms93/va+gRM3cZUOgY6gP8QYYbWJj9
zXIVKkBOn6FJ+wk3h6nr79QDW6FqQDZTX53JnWtYgmtV3vejUtgh06p7XQXapcpk
ng/p61ZbUN9y6YUxThrDz9Kfs9//nwxegjBtI15MpDIyfGmxK1Nyyj6kgfkQ8RtZ
pgeJT8WRYBVtSw1+4pv9dZ0cVTe1wtWt2gjJmRf9lrmDh5ajuWLf/90z5oZ6AIGu
Qf77XFr/ySdCQAYCMe2wPsDOq4rHMeqiF+Cmobb2bCGUyVAd7PMBIsgZecHmWtur
8NgyQRMmgC0C/TByfaeQLTRxBZLXtUvkWwft42YDuOWav/0YEiDFC+XpYlOe6Hi6
sEb/niXluRNLZttLyiIDtlIZm4FBcBEaYe1S4WS6zHODE4o5aD02KhavLnXr/EpC
7KFZh/Fo8gqUhVaeQr12HP5OokJ6XZJ2QaFkwSswPlgwQ/ILg7sqXtm3oStYNQdP
qirh7ML36UXVO2HKlrBYTfQmPlrkJjBlHiwiTEMcNNDSBrFBzh7hXLy8HJAG+0vO
Srfq/ohHOmPCpRHiwUMcNczDVXU+3Wq1p2Sn9XfTIpIDZLXoTpS11tgzL9nHyVkm
ZBqnPcRciBqepr5M1EQiZHradMLnJDGoaDVzSy0QVq1pHNzixjdpK7cBiIu7OGk5
94QVxWaP6g3kFF/UGIKE9dqK7VlwTlUu/+I/ZuPp7GGFAZvyRHUuOeYjZQzY7lDo
UJps511vJpe4skEJLFfugHYZ4j6HEAfQ7ZahY6pdTazz2LGZNUE1zcFCyYBTvJa3
lYYHqhblmhec+QaSd1nVa3AhEDRU24iNiRLSxTa23Kj4LwVU4xjMMygEEPYcqQKm
nrTcNayysNWkSskOpEk12aXbWV9vnqjhTQR+pKasee1Xp9/oqCpH+BGFZq7h7OqX
SEN0YdJrWcM3Heo/YhkFDXuecfCfzemsSE+YWou50OF+P3UIKvDKZAXAdqIL23dg
g9xiNoNE0C0msMefORYlOQMDt3R57OtGzH0gDac+ymeCVmots4RjdnSZ1LK9Dekp
/kNNUeH4fwPncOVUIZQJU+8awppd7jUW+g4S7wvjHzpAQ6oWG/kzBKcdsu3g5JZW
szSeBGCQx+IPJCS+4ZqhdsdY5WJbI4zx4XmS2d0w1wPYxD4S/ibKWswGF+TOuqZk
n7ceN+Xghoi8Iss4C2pDVHjW0FJ8JYAEJ8YY81g9CdPzxZgzVOdn6ufq6tMlV7Jo
SozF4u5CIJtgkpEYiPimgAV040wXmPuMYXJyjTpfoMvNuA1vDnN6AX+aP4OBpuol
r6jv19BhPD1emrmy/EjjgxfPxMhN2szeTGTk16VDt5C/kF22yAv0HuIgKQaxeEj7
X7Jzdv54HLsmlErL7JmqOF3b1DDzma8Gm6bJSi0WffoUgjWDj2GgIVEijPW+TZCz
y7EWH2RXQkxjmAskexzJsXuLWNq1qST9/8DfDWQKN3PQAVR5f+8i1XS5n3QH0bFZ
P1gZQljI337FbR+Vhe2BFFzir8+r/5+m2G8aKbStHdt38pqBjm//gYF/quJmz/qA
u94DiY/tdZ9Sy6M42edPqKKqrImWPtV4/QLm/nj7omkG5Oh0S0YWFRR/sBKaJ8fh
+VaJ3r1dXzT97fld4vYNHvilj7UI6GSpihW/jpJhnzTgn2XSXgZf6hCjmTdgFrwl
73Vg4w3DPuRw8HhMV6d+ezC4Qezdf92687JZqYJefdkoE+PAuMo1miqaoDktj4S2
5nf9XoeRPNfccikqpGoStaL/JfuM9tK0Xjm+xekQ7vYXFXAs/8Xgbz/WFhoNCX1I
xpK92pPLk7U8HRTzDjwTVyOIXKznTbi1AcFio5zD90p91Q75V2u4/O4aWFPFMsLT
WBnWo9y9j/xA4ljlAPibgNbCNJHMruuM4lTf7WYkGkryLt/U3tnFY4ZrNnViYRDc
EvEK/P2+PfzcGZa7KD2Yc1KIaj7HFYDVlOmHqxZHvN8uK1kq9t9Z7Jzflnevejye
3WIuE2RrwEH8wqx5L9HfoSvs2dgYSigzSxwz6LghVnD1R9GL/tFPGMt5GTtosThg
RpK9Ov2GcAA30J4/jcZVozLJwyerdaQ5gOm5mlzJmpbqr6+HuSO2SjoPJEQE/cdK
v7O6Ika39xn8IcQKBTWdoyPWQrAnsD/tiv3bz7VSwJk7OIwihaOXmho3WF8qz131
9+KFAKKqe9uC/RqNFmkynKFsnAlYh3Wxv71qy1peE6kLNcs2KsHmmLcxOcdKY2av
pECvBV0cQDnSDRStmysvGFqD69b5J7KzzZjkN0yIiv7Ft4QDIKbCTsLjbRArkCJf
QC61jFs+8C/94cVyeBxtP4LlCaeb1Z874tAOPCAe5YfHJgKwDdLSZ/hQ6JaoCOYz
sW58Drocy32FGamuJHdghH3zZ3wJOEEvr1KzJlPjOpMFLki8sAcT56yoUM7CdUXI
ZyxxKP6SqS+Bma3iDHw+3pukBSpRgACAeJGNhn6r/psnmh7lQxnJKOe3cTVjs99Z
c7UfQGDZphf38suLy51Us5x9prI0L/R7cElUIxPzJ6sCvcL4qWU+IVzNYctenQ2n
KQtLVJsURQo0Ad5ETI+dpF/EHrnwmNM5ZrlFpwpw6glG/2d2XWnuCDKPgziLJWkD
urYlVB9zk2ak6y7cmIMUEKD34WKcLtQ0Cd+JqPPkLQeDHq2H9Uam53kxrIhokeT5
ikzNDagoXZIUMnS4PsTVlpFTrerlGG7+JLabiioFS4KUP/mbTWcihxRtmRpYEJyT
k8gIadd6ONDGQc8YSOmU+vgj5IkddVQjYCfFK09gqxjzcrzoE706qRbPt9+TCT+R
Mr+XbjkZg05KmgT+uJmHTnvjIaRweeCMHfwEa5CgPdVrK/wpqvMl9QtfNCf39ph5
sATLdE84N0OzFGKkW41GK+qCSDq7rA37LXOtCMELGoG06dkQ9p2gkw0Kc3e1Xay/
ertErx8rSQ+9e1y5eYQY2LxAnbiQeygLkW4idqJgYlHo3HUcFCTlL86e35DP+rKI
uWNc1XgTh4daB7/nPCLlPEVc4RG9W7Ug1aJm1Zu0ptsbiWth38Sb2bwkmd4XBuCm
8y2YaJomTASQFr0P/Syy49zRT8GOAPRLC0BWxhXvm5BNfh46ycWe/7AXZCMa/Iti
zOiX5pymFNAyG4AUYELPxMJ8vWrRja1cx9fCfpC2fDPZOID/7xQQTJUXqJ/5Htzy
ulgPvGGm/DPcW3diciFhL6oXEQXwXEkBiN6jhmfQs9DTyiwNXnVLVK030f3N+7R+
rehe+S1sjpRo0kjL6wyuEEZNvIDIyUTOluDuWgscu/F0WywzOVwe3fql+4z4fLau
iaax+XDgDGOpheSUqiUtBR9BIAmmAEoYg/zY67CL1h92sf46C+MpviHYg44wphOP
cCm7TYnP7TAiA6SZYIbP3sNcOtug6Hak1nUEOsIVf/AIEJHTwe/d47KDLBM32M26
PIb5YzRArE1JRmdfPmXD+ITfPuXHu4PZcCRMImkV/l13cujRc5TBnhRnCciSxfrN
nFxcK1Ub22RHLpea5JEDIIihMMDctwZIfG+rN0mP9PA8WutDkyR0K9LJzxFsDgQe
GesYJTuUBSNuTiYftj7AS8yBSd/LEF0FW5POXGvv94diu80aYVrSei65y4PcP/D/
7ReEFW/+xzhpDWAsY+3WqrDwvDNCYajzQOQ7Dn/IC01nEQXc1n1StjdElWVvyAMX
OJuMy0S0P9w3I2ImlauYrFnsS751qEw4EGo1enrOVsY9NWtTMgI4DzBjvXLZCaY7
CeI6TVk9/GYGESfQzQKAizNWvzZTrqCSRlXYZ82T7SrgiAJpoWkhyrASMpKbCN6f
YMRqEJHnErQZ9+RFVjfe38Phvcr1nyxxwIH0Q9fvYSs5diM7qH1GLbbx/j4KWfXk
EGvCqmUtd1hnQkDYdiwvN2hMepSKKi+IzS7Rlm4WIuKk+Mh50ybfD4HKPljiVOec
UgpMDnBRDBDLgVffmt/aXLnoHwUzl/IA7Fg18DsFfozdhs2FYDeS6JCTvHyFWaPS
wZXMC21hor2i+1EQEyaJKHt4KjPa+Hgr+bwM6kehOaOGL9aqFQZ5qpjg6gu994eO
4vyHENz9UhUwFBUToBVt/p3lqQnVhiU5612vfNfoqH2pLXlUZpfkAM3R+tr7W+Pu
1mcNK+Ii7GpP5e0q0UqYZi/KrQ2vpOpEOo3i0NzHLc6go3ztSSoWd8y6WkQb0Rhs
m+Z5SIqdmPxdi07VgCwh+vIl4IdVd8rEKhjCds5nXO0OXGKuB5uuoWW8lhIWBbZp
gg5IC57sZOv5Z9CVVeorgWcWQUv1jBaxOyRMrJ7qhEzs7ycstY4IZt4w605mkYhv
UtJWZOEDTPDzzRr0UZF3RgOf0Gq0mhlKB3KonsCckuZfgYt7XAAoNRyiiv0zOFpm
BIi3KUnmtNuZeVZpItzKHKkgIdEKE/kyLJGktZOy2zb5NlWB2KbBV6z70KmLqHT2
yzZwcnugSJ8CKdozvApBs3h8CjnWRrW5Xdtv60/Lb5omGO5VIEIotzd89c2eqDin
o3xp/LQnFzDc6/XAVMHCdx9zp1OjIowY6Q7CoXgS8hOt0kkjmwOF7+bkSXG4Ivx1
CELa+dSBCrJ308PI/2FyxC2GBavytQaoEdotku48vzcah3inDU3wprVQFqJ77XHh
zVVBAi+tCztGzzdrAhVHvshjdCTDm8fYrXo1aZjRiWQVnQJ5h469wt20S3cHd1WA
tnUir5Ci8K6UubzE04912UsX/viPKmYvQ/JQXuSBuhWT0SgjK/0dPi63zBhd2xgv
vualhvm/Ysbk6f6zQNhFhMjMJ9AMB2HVTZyM0+k2PlxZN15Pz8OYQcF5BGU/ESJn
Oozrrx2IWLyUXBy701BYbnz8RQ2IzcLToVJI2OScxGuQGXMFk/e7aJiJwg56gXZK
Hjqt/JvFhkyPEJNlw1y6nskXIaFD91RDSk+8HXVO2Q8+fSVnbBv8heB2wQYlpvbx
odiLYhFAUKQ7Ho6vfxT3wxbOMIs/G/Cqy+qHYSldwwTsbjFtzmLxq1hxO6RBQauv
Os3vGnZxkgpuoT/2qXH18j1q5pPmc2TYL4G3xdibcHzGEvJipfm3vrHUDLdTctt7
kQuFHE1HX8woWoAWsY4/S8G5bb8L3eQUMwifzpPg2JN2D2R6XhIcRi2amyO6Riq/
0VdZIHt+hWAIDbLPS7A11MlYx6KJTllpNAIAZQKunSx9uqi6TDxgkl3OqXiKINxN
B5rxk6DaOtbq+8S6ZwZyX1OwjXou9MOGoFURAD7YQIZDiBgcivdvxhljd+cLaeDY
zmBMDAx4lOTeRvW1RNVYfZug2sMmXfQN3f1XCRrBu21SgQYtB1PZoIgQ0MLHMznE
EzFOcGrcAiimy8RCGx95EWlJ19K8Z5R17mNWZx0XXznNGGCZv3F90HsvZISdXGsX
Iux7JRbhL3qNF1wwUjy9r8qfehxOPGbDOzNSxAEEgwYCPDkGVrECcYY8EfYHjs7b
pneTwzBWWt8hCTS0tz7GSUtUTovANctnOFJf10n4LL59B+3OzQvOtLY4e46I7kPl
tVxxEUjvjhN+a7L7C+yJQSB6YVHjBHqp6Pw2552ZFygyCdPVL7cX25NiiWlnFIqF
YE9LJixocr/i2bhYdfV+FEmIl6nSPHP8sRd5G3y3X5dg/ft3kjydOStcvlQV99GW
Ltiqc+UD+oZ2BA3I+aQLAVgf3jgn+kN79fZEBqZWl3ATS6gDD0ntJzUTXlwzscya
KdeIM9L3jKrtEx83OKIqt4YqZNaUxfbspxC68QZ7o3DomDTyhDpIlBTrQV5mn7L0
/TVvjUJIkr2fqpd6IOqKFnAjTXXWm6XlhfWNcq+eVfgN41WrY7Z8aVDiRNw+mofh
RtteULtuuZF0L8GOqOgZ6DbqD0NI6qfKuaQhUerdDRUz1zGsEcfd6jhEqCz+fPMO
dLqDnq2q1bYxLNjpxEl+g56h3YXhpK+Kp9KIz6v2JE7Pxmz7dK6fjc2XwvehCLnV
slgVvwxtxXbsyE20JxlkVl3z5MeMd/1Q+MCP8szwjA0k1EF8yHjw47uQcJPJC0jZ
b3P0/y+0vKI4v8dC7rL+3mVE0KFHUqJlMpxwaRXDmbIoTnFnUbxMQWzwShvAt6Aq
delH9rJnWvueqCr7yF/HqR2AfDL6AugfQvQd2sgulvmJJczLgUmG5V1JhyRMS6RY
X8OSrKXbQKy4OPaM5F7AFs3jN0P2lccnkaaI91FUngdwsqqR0wHtz9DxYBZRHVsZ
bePjkdWvQJwWhqtvq1T/oSROKpkcc7tghTWb5M3U6JAc5u6IhO8DfevecLtxYvDJ
ab2GUrnr4oCgoN/tHorNAOz6MdBjsAlxw+jyQ1wn6QJ60fQ4SOlLqED6WY0E773Q
qvTvg9q2s+AYbaV3xHrBRz7voDBI94aKxjnqWYiTHKTh2mSJ8bj5LOQO5L7ROAhZ
tXs7u9jVI9P3ZDmPKWWV2VItz9KHQAuF1ED2OwrfwYqkhtgzyOojB9bhCZjRR7QQ
Z0odWwhkyEA9VAxDZoY6/x+F8XJm5wrlBozRhqfqlHv1qf5bakyLVmtzB/zrtCE3
fK0u7+R02Syq5T/3fvKDKUuhefTG+fImB8+OgsvjZafWXnqpYoptvSTz5wSGzTLz
C8b8l/x8QIAJQ1gmJLXoOVHlcJgIRpqNHoW/SSr/Veh76g7j2zmttGGDpFbyiMhV
4ZDF545iF+8iY4e5e5wv7bbbydiLNJ3C3yqc4tdsI9jbmOn2Gd8eg1NsWDktW4Aa
t5TfQ1+QVQIRmbJ42hvWWXjUNFKEpIa+SNHuTDZ6r5eENtLYF6U65EHgjIcXT7FK
JjuusLQjObkO86WZikb+r+zYX4COGwLdCW3JAUhE4QnhSMEwzP3bF25zTP2yQbcJ
jICPdbgb5A5Uqq59tq4JPqXhTlJXtZqn3rRPMRHEaW+DQL7bZIifIU7Ub+GLZ9su
r+3AknX/hehdR8AoipHx5f2F/Rqu6DBS7aIYLMIs9iAiwp8B6+jAjsJFQLoAl2nF
D8OiDZJlS+7/g9xNM0gQQQK8stvnsm8mstqgaLGxCkxWB9eSpQ4ic1rAwWRaokCd
AlR3Ze9dMlinc6ThIsaAMixj4Pz9PWgaiP3g/79zbI0KymGQRDkMe414Tlzl8WoX
fJ8LgB6oZ34O7gRLN1NgAMKkXrdtH+WBo+N8UjRNG/6C1Xwo+V7jUOc+JaibSPGr
QH9k6Kv5n5KGL6CmLouZwimV3v+4ZiUjS3IrumZT5QOA0+YiD1q3JQosbZiPjzGQ
4BxoTnQ43R5SuQufRqGwphYUcVXAl3S+vGlWLj4kJL1UxcK2k2aZU9/ON52brTCB
zvdugzgbKos+xM/RvmMqkdrtrc93OKO8PA/s87mpVp2acud8UyoKLfZOMP0iz7Yj
xgeOhI28dHZmfFAyXvSJNcCUPiIJW/vaRTyDM4Hmc0pBGeM+6p0+sXgkOaHWplN3
ww/tqYsawLQ5yiakFKYfylKgEXPEEPYKmDqHKGkluzbTnI+KejyLuOGom1A+vHdt
KON4o3m2KEuYNlSd1Q7/GFSFiS5dKScxgfPv7WLv53O3vE7fvVB8hyFKx0cu2r2M
fk6CYkyauzkKFbm0r3gKfsQ37arAwfDNesd2z21fMQ0rr8GFL+fAVpGKVubzbu3U
qn68IWqTDOn0V06ZrPU9+kTas1V2GQNkdlzptmmcd04jMI8uua+//gy7XQ52wNQA
mfoHuQcaL1ezoP/e7RoL9mTsAthJBArAJeCTmuZ4Gc0izX8DFwXw4tXkr0NBZYQf
7/WbaFgbdERWno75OJxjxVi+cC209NVXgE/iB0AZifM+fFbTbAKxdRDtFWmWmXXC
oU1jZK2E5vi9L1zowA+dT5Dn6YvYCmHTvXPT5z+mPDogMffRurpZ+0UbBK5g3ir0
8IJEBnjY7+cAZbhH+OH+IlxHGQ/QXX3wnDNvC6MvBbIQvKvR0PDlI3kqxlIsWQIJ
zQAoJ6trpcoEoNpfk5vLlfN95IFQo/wfz32u/3JZr0H4GZtJVIqqAnqycEIBs4rb
v+QCe3FLiuUxap0M6dlxVr6vM7U4vKNJkZCb3LAlGfK5Z33x/ogNml2FNIjSEgVC
+fZc05v+Wx209m78UsIeTzH/WgdlC9Xa/+y/3mhqaPyN3im1asKZT2gHG33olGkE
Z6Bp4vMDHMmoLVVsGSWfDfzlDB+5PLe1CYzSAyT3HSTvPYR91OzcTkuTa+yKfL+F
lDOLeWN3A6GXBGyDIhedzlXSnq3RPAln43sKIbm7JusKB9A/fV/D0f4UdZsfom8I
JQHULDmv4pJFEN0exGC6TgtNzDMvjfR6pDF9pS2etTAH4McX3ZI/n3+jYP7DlVRB
P8JkVBe8Qs/fdCrP1GeAZbTEP/Yg2NJm4u7UseZLlt0AX/9htfhYh8wcy4kzx1KN
+WnKyzCO3UPqLvnhdhqnNou8SZ1OAisoJ8g15jC/DY0sLu2cBMCJd9ovRkQW15Ye
f3fQm/PujqL656bdlY1GKJ8dlRGgEhDb5tg84ivMnQw9xsYqMXZt/LTYvzvqSSvv
iPufDTUkI/wpifhvYiepSRHd73vXOkojXFhTMMce7drHPJQjlaQX0w/B/dfUN29Y
4zCldb8hY3+zIbOjTkdWO7OhFh+jAQJkjVUtGVCmuMTliGVsLd1gqsZKSpPOJWT9
QHs47mv44vURqAcqqUMFEK9zQQzYLdzTlkOLy5C5Ev1LtOZdtsGZoLc+adxr6Izd
UV6YgFpeEZrTHOmvNR6oWjzDfMbNWzs+HggfEji85kqVdrGACnn6v8Eh+kwm2rU/
4YmNC9CuRsjJeAYwC+DU5tF717d+xPjbT8CExbU1bqFbxHfml3tH8EFo98/ZSkOn
fuPhnsNmj+n9GzymdUOdH6ur/fvCoLWLUuZymJQN2TJ8itV9IaL6gmKEjn2QqUeC
NZ4qXyyX5H+qT14MqT2XaqQ4FJUZDQmwn0+e1RM6cYflLfMzW33upfFBNMq4nlF4
i1JtKnzxpV+XjYYuQkrj4Xa0BhSLk9+xjDxZ5soYPO3LESF4Cmq/XJfSzgEa0bzM
4ZFijcKI3g8bM02MpLhUqkmeJH52f01nXF4pjovoDXvQ9iDz6cB70ONJpeysLWWr
s11v3JG5Pg189s5Xbv6nqXswSQkRJ8OEzwJfmi9+43Y6y7mQlJaqWeXk6k21wm0C
HQAno1deNX9+J4ECy635VxM8K84q4gVOcDxNrgbE8NO5r4ix281bfDbs8TaZQx71
dGSYC9pecJevDpWniHBO126i/eRiKq1+w1o/IZ7aNNoOaGczDhJGcZwQwh/uRLWh
gBuvTg3yuYWBXB8ni/mwrhDggKZ0evYACD84Auy/Dq8kRGqab9s4kR5v/2hz8YZP
yfDgLhus7Z1EJd+Y/ImMo3gJF2OPh31/HXotADQs81H+S61WGKKLUJn4+E4RCmPl
A7CRJX33sLijxG/wviv7YPU4opdOEbUqwoMFvmIBz759whnYx/CWnW0+Y9XdmBgS
qio1y4XViaiG5fql3UV8wHYJmyKztafzX6PEyN45MMNfYJbPCsriPaOVzdZKCepd
DA1Er/N6zBgYVLVKZhhIRDiMs/jHDkiYgLJxa0Z4gDeXMuWwx0yhV04zB2P/+F7Z
whIcOPBaE8A541f4rKm5B3w9XwPFauaDOrZ7fFVCMJ9dYloA7w8MzU60Lep5cm82
vFad/QN4rWoSYMwxgZKGgdTbjjrdRlUsR1D5a+IB0ckaicKAN7R1DpkcjttIyhwW
vELBEQZBUx4pGwHSNKS+MFfaR0y2iv/I2Zlcg87EhfyLqVUTS7sGeTMs9Sq3fMEH
FmFlZfN2L0pIbXelQ1XruEjGUhTSCF1DA2bfoX1jpnCSK0GJPJugAfAcJTTRDDkE
n9zV2EowHr4H/ER/YMMisRn6qZGNotvjRfrOjsJwPB61Ii/bf6gXWVaZsHD5bfnc
9XN1Rne3Kgbnj4dDitM8nvOnhKV4GtaaSaRrwWb6zQ8JjcDQZCrJAf3YRW0DwNUM
fiow4svAN505CcPrfiHfXB1cKBhHsW4Rs8UB2+aD6nwYjlfByFRKYTt10fGcv2Lg
9T581JRHF/rE7jxgRFXRbZ0UEpO3FJFr6vsiQ/naSJlnJQg+XDIOe6KJNlWvBC5N
2D4TpMLUgG7v5DfsP17zuEIiSUXSwxCtmMVLbdBdHF7OKOOt8ybowrbyp9tcD+8H
xXBhnG88lZLf0zTrFYicH+WZAmi8/n8JIPeiURbT8ZYu9g0YyKiO8WXWHyXFcSiC
lwzDLMpui4i2DcNmMpCMsFwR20OSwEUW9Vwffk0ieeYViHO7aEZrjyjdPfJZnCqp
l1amKIdiDyaoi6CHwf5BoCXOel8QCAOHysGnAdKtBN1JGduO7MyH0EQWuBEXaU/a
Li4kwXxg6nBk8htz3OH3u/QU6oeuu6GPlE6plRNZGR/tScW6ZrmWQ27yAsasvDg4
Utfp29m/jO2yRBA3HkePBltiv9lDowb6GdmzQVLDfR8f7gZi8G/wSccilALRLvOQ
HFSfefj1wo69+5XHZ9KQfkevT/0h/mHVsSRmE5JdVYnBA1rpwpIKPCbtsUuOlqdW
5fnutDx3zzNNIr9Cs9vtKfTKVmAgfmGeo4kSX5pB7I7uBMCLJhlfDUREuGtpRhdt
rC0tgJtT30QJMnmQRFmCd4jPZRpYZGhoVrYo58CjExa4nnw/NmxowWBfqqFH2Kmh
iZCXNCRJ/7XdvQsOqM8IRULCEMTGoeVjp8be95QSbYXOEFkSz9dKjmDDetzv8sB8
SLaYD22tjcoWhWH1J/zNyQMiIX+XMqS5hrmRKXbaYkOMo7VGCWv3ImlhYOWAWw5B
ud/G0zGvOyjpjNbbMMyOWHhgIYdV6ZUSj2Q/K0cPOiMxlyH34zN/HZpHnp8gB5l1
x2B+ycYgt4UAsc1k1zso4yPeOgs1j1qk3Wjk9/ADyiZ+yjmwLDwNnlcJ77szuKF9
s3WN6itX5Ixg1WnTdw9od6+ZFKjHiGvfSMF6RAEKzY+uSGYKtUlJVSRUO3sMg5QO
K/9DpK+S7Ni+I0NKCsUgylGIdFDYXEtN8nqcgkRYe5/Vd0HnWb7cYahvUaic19nP
GAPSFsJAsoov20jzyRYA7lCWGuMt905OvSlyr4CMUKHKmgirN4/wSLd8oyhwNA6O
XqmEqMEE1bqGA2Z8P87zzlWST1lkhWOlx+icno+XmXxS35MzfPo5Eip/ohz+Y8+P
73zPcEF8V234cK5QgbACgn5Ez5/W2m7ylkU2MlQt6aJXodQhJUnzelwLwGKEFI9Y
CSxboT75+Llujy7mWQtn0A38umI4GX67DjeiiDX+YejOxJcQxC349Yi7TcGIFcOr
tat9MbGri47OiijtYbPcHisto83d40A9hPciQd291TnU3QriOVGMJfE9JALM/lLz
HJgPsAQLtPmAAU702CaPeIeH1TPsMiU81enLE/sbPzczGYGEN47b1mIjoWd4nFXI
UpkGyUZ051F8X7GOhm/ps4tCQfJ9UP0pZkAgueEV7JcNt/54Oq1zv/CsWBS6GJO5
gOGwfgZ55IiAj+eIIsOq6fiRi4Pj1PG0NEJIPhHsCKsrsd2tlGw5qGf8kZORr8xm
VwL8B5+xDn/tcAazOlZKhZEyTBXKIJAq//vAfAFjY5KwZReo/Bcf/R/YbUCdJVfm
ufT/ulItM7UrDM4EIwZMUWQjX6tme/qcDkEOGTMNeNmjGF0ZOD+7mbQtYg+6myui
maP5IEQ369zg8JyJQclxWm8FyJET0VldL/L+C8ZOqXXXBZLDgFXgwlU5hsLDzFIC
MgS1SqCwi+uomlDcDPcBNwqRoqiRvEWVNS2ekt8FTCKcl2xqmCJL56SyiXyfrFo3
3ErWA+7Xhbce90TFFBROqOg4arVn+DZl5Pp6Ye828xjhb7Zn4A+kS94l3NEtA9Xx
TF/yoGIR/WUsOnBZmak2Dr8FAHnDRxr39A6BBusqM7e0ACMmIMWzkWUjzOs+3xyM
LmsT4D+23ycCWT5mEasQIyBD4zG5umOhIqY7AxHzClP7J8W98Km7fziZuiNdIDPz
J2+hofb2NIYFwrjxv5pj0NyNEX+bxoOlO6u2RRQa+6mlH6to5plnhZoMH07mfQ+D
P4PvTd1T9gcR8KrPh0MAJf/H8lL8Kn50iQA7qn6EKCqrkjAZiMB9lFnoH/g5uOZm
MQNhywbBEBhFntaSqNOQRuymC2RdlpcpdVID1UaXHocBNIFrrWvFGFGdJGRKrrks
a/tAKSFbK4q76PECXtZsWRjmTcLS51fC0KGhpkQgAsbKG8LulZtYAgVIYp5gJmlb
XhNPrk5n1WqnTXMuQ3jHv9m3t6WidEF6UEJvkDsc9NZUtHH7KVi2PD5elTo426CT
N41spve8ZZ/zL/eREoO8Jd2uKQh9kb9iTvNHsRw5QRxjI0ZHyZQPfL8fibBs76Yc
BTmt+Y4faAYL/ba+jFwvUqVdv8+IP/NoupNFRGdhjcOjWpfXID5PLmu5C9YoJMsc
qUTeNuT9QdTjEENWjMw5bmfYlRv+r2EfgtVhwwVZHHPW/eyBW8XLuKSfNwgt2syE
9UGXwfiM8tsw5CnZ2QnJwpnKx6u2Ge2r84TQ8gnjUEPF2xjX9rgwM58JyR7zT+i0
MbxVxvj8AWZi4uahiuRkB/BGfS0qopLsG6SZM4Zcl7a0b5543sYsdkM6/BktmN1Z
6S9D4vtaREQwnJ8vkMrOet2bkNIhvxXNMnirBZR2vNf68tOrzuMVkqOljMBODXJd
DtP9IMtyt4Fm7aspRpM9jQO5Gi1uDPKP1D49ufGqTMAXABnUGs5+cZNCu5565OEk
FgPKcxn93s0sWJ436hqbG9W44Kij3KBYgmbrLjRfwOwfAm/ouEVprxXHFIHBxEFt
KYnSJDkW70uyWAp52qO8fWre2KV7euGsIsG15o+6JN42kbY6G3imCYkj7Uu3PuXI
z3FMVNnoayg3NjYwWidfzlacmLt6LZAckjAkQCAJVxYAKkr2oP4lTfFPBDiEwt0n
xIHqqlpz3BHaoEk3h+eUles2PtopRnYVp8qxCjSdJ3fFWPmZYlp7A4IOKmH23MUE
UhBslaYjCOeaWWzyOHu3FbZgr5XPNQiT5Sao5S9boI7LmtcmRMoJW2X7xxyB+IfI
TYBNWKV22VKRXsO+WKATSQVOI/UKPeELVa4UL6IpzonlyFkvG9wggM+QJt+oP1cO
ppU1jkRQN9PyBexuNdpvsPGXtcsUbeTPIFraTp4cK4JXjYb7YIyg/ab1+lD9XrLb
fIYnYX+WQknYX2roL57u1+48hV73fciVxcHGznHoEwpu6vgdbz9NY1a5voT/KWgD
+sQgREuBZoH3rOC9FLwWyvM9VF8LCjWsMFSsA5Fv7cbOZJQeWMKtVlHDr2g7TYSt
0zy6KH/KqVNVh23mNhTozSePZy8CD8KQ0dZ2bdWT8Q94hr2sxxp8wRC/YvPDGNrM
ERypLiFH0juEJYvKeqJ4JfrkTS1K73iGqV2Ksm0gX/QGj+Ti9SuLJ4IP+fptQOG4
lHaJyW2OV3c/K/R9zGuyAERLUKeFL1YSjue5LS3uf6UjWS8Rm3E8/GmzdQxibx1D
M/S3avVO0frSHT/qfPBJCy+jraEU2s8K/BBFdThhASMEJYTma86ByR54Eeh90HcK
vFLjnOEETTS2T5BrcRPqCl/obG001LQnW3bi4ZWo7n6pWqJD3YoFpgu/fPBeQ+fN
3r0e5Y+SkotCQazecFwPjFNBueetcH9TctrTVp1ouX5VgTZL1ivaALtg6waEzsUT
9Td3b5EGcYITIzFg+8Zxg0FDRk6sIrxKGHfth61BoesOzNoDK+qG5DUwM5venzsb
WFeqbisyIuzP8OiFC4rtUra4ArI06mkw0L6ijrINqXSeFFtdnAo8ZWPVHZfxngHx
xhhbwH49Jsy9KavFxXRqHCEyAXULQg5uJHNM1A+reniGVwzfH+8W9QdujW6Opnn4
HAoVYkWsCXY/8r6zL7c9y8tSw5onFhb84OV05SJae9ZuyBMY/0kkFICTvklN/dwr
RzUxY63rK23P5WaK+/xKzlgvu15c8IEnykfWF1RMlHDuO7RvjEIDmgLpG8zDGVEo
TxkI4zA/Y59RajhifGbaiO2EruwOVcdIhFKLWd5F4kwea9HlwdmKP2lwLIFZI03Y
03+zjaaPnOl7lGiHoh1NHeKXZio9WKsLdID5pRQJdcrOB+EKv3fYu1F+n9e6NtEg
+j5mdi9AyCvyJ/uU0hnmwyh2Io+/smtaYwufKy6I8uQV05S56UtX8iTV50nuq4Sk
Q927W64+CzG4GzmtfS8/0jg0jeNPfoC/OEqs2UZGNqG513cXwZlvhu5jXQW8xNld
8cK07PfdDXAJozg2Xti94QLcGxEh4TVdBpg/5aefIvPxbqVOjzjo0MhmccnkGQSR
Dt2n69KC0ARaOd7qrinE+WCdeQA+ia/Quc7hW48eCkcoZQdX+THjTcm40N8z1vwA
Ydbolr0YTqpckhlvbGDxHMUdtoJJAciUKruUczYkY9d5DeJ8MNp5NVwU01eJGVhQ
7Upkl467CrIDRWPAk6PAUr7rt/QWS7HRm/ArwrC5CiJDf5dt63JYR6KAg9QXPS9p
7AYnEEpyXYIMZCiSsD6Twbwiy59g7/yNjDbOYYfAtM0cat5Z4o8it7uduBVHArrj
VOaiGfxYbX+rlbXtDh8q8pqUK3YmcOLqwyXcrgsW9dXE+pnIgy9aUeLbTh/BeSdl
XBtxSiTxZ46lkpXZJSfRQcJtWsghjoYYGotAGaBwPIZdIwWyApHuZ7HBFxe22hSF
2h3AUWwFxbolpEUyTA5K+MuDEyCqvSbPE20xyS0FMbpMszPZt9FwDUFEeHmMOJwL
X+LnErSU8zYcJbHYGE+gQqkc/Yxin4p2ug87yQBDS+9UOjjlKas3hpjFBkNPkITa
SgJBwUYOcM/8aK2JHbkYEAIfFp4oDmD+NC0Wx5t8x6xKzrcfApcoeUYwcC8njC1+
PSzbZok1FMnm70qC8waPNdFI5mfj2wMmw4v/z+e0xPEBeA4QVXtjKjq4+KruEUUz
TOQU6hRo7+IROzopeT9QE6vQkSyv7FbYdfLtSo5EQUKLCosqQhA88qpteuZBr5fS
v8yryDvXnqGRGANydSIAuYcJC3gd+aZaod74FzQI8MOOaA3JfXrUOzqAkWJRTCjB
GHsx2KJG8E3yA8VJEV1ZkbXogoyGfeDS7bIqsWxHl6FNg6+FSSX7DtoX4NtZY7MP
Xq/rxnRrf+M7wOC2MZI3+EvB93XCPpz/UTCciNj+qEtYKhHKMDQS14HG1JBbfjRU
X/gAVYC4EnvjZj5Ysw4R0wunVgcpHNw+sbEsxVUsx9PATD3Yj4dQocxqHJWl7vzJ
hW5WVKPWQGfKIhgr6no+Z7l7pBXH9ZiTO7ih0oVAifqoPKKEJ0N9Tl/LH9e1r/W7
xeCINcgoFLOb9030n2AzNwREKb5/Ur39IpazZlKf6eD20GwaGxLKukqdwisc1hA/
wltFi2a3WmtZDHDthBX/x+vLTKxg/qIFm5OkYwQQKZIeHY9nkCILgl+Ilr7tySii
bP8khcrDbD/BtoLem5ajtugPFJOqufeBkrRjXf8hcjJF1HkvA/AiHuqUHESJFBgt
7vdUfivR0EdNSL0SCvNTzQMaCgP1AxipJKHZdrk0OxSpXRJGBqkeY2CVVavSuiRg
q0TZQfiuSeB2yuWGoX177Sz5pVw1ClBltDne6GDYd64zJDseyAbQYBg3cZX8HFYi
7vRbdCiDz6Bevx7gNvVSzDvc5n4vkBWEbVwm21pjJ08IhiCpnkA51+gcwhTI9i21
u5b9WnL99nv71OhOKAmXFYfsm63K6f95Iio/I37vKFGsRmSTQQ9gl0XZ2mH3ecIO
RRld8ye9HPB8IzNAOBU2kN3LLxECEc4fkHGBkGoSnfuF6QHDRYu5zJ++ecPOrEo5
GwIUFrPM3KjZDpzQYuJ847S2+mP+847jSGMM0Xbe7Gcq4gtRqOxubYT1IfXJayIj
yvPNDUBLHtybzk/PVM7h2BYsdjxMTFqrXLquNSTIuuIvfTFds3bDH5mnOqOIRCsB
vTDyTf3+jED+OR6i/bp5IAbxQt0DNjQqV7bVtCuMhiwIREmd5nGRT0X6Qd75k105
I6Rf+K1E3xMTpZqkqXTmpGLMxKlOBKmxxETcMCP6YwLRRh/9Kj8c3AXAhE7xit7+
cIWMYsmU2B5oGP6LO5ZPpBeL9QUO4nowORQKbUcX7lh0eF/nxDWcPieLUiA0Idtu
G3+nG/KOSRbHO1ZwLJvaJu0IT9+ARAS9SHKl3NpDDZSsnC/jjIGjKzfIRRAQ7qnV
XZfEPzkQHVsRQLJkvKZVTkoNLZazR1o4ZXuwgX80vvNPBBBJZWELA+FlGfYd/pGf
XWbtd6bR+Y4dC63JbZ1ZT+Wb6TzWzaVb8Jw1PtJezgu7RMtOzsH1S0mBFLhiNj74
7OdaMZKDhdeoj6PpDv6DRwg9oAVFbz3O5xjysOKbKoGIneyDeMnFvACZVmMbmhiJ
wHcE6IoR1xZXjuE2vevIA1+KKumQviNJTq5skLGPQcw=
`pragma protect end_protected

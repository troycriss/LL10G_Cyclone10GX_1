`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
Z2SNCVOMs+ZvYrPgwPYOevC2rZxEp3ny2kY/Au4X4DYaqTfKHqSHaj595DCwefas
8uInh0Y+cCdREUoPrzf1jou4D7FAvrZjED/gFWvJaFFCZeezAVh8u63cBO8Gfw20
QMaYa4u9g3nx5G1kg1eM50BBK3uA1GbRJJ42hqYaIh0=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 2475584), data_block
7lSFOQ7vwAC4DjG+sng9VlgPmXcRKga2MY2+XAd00r3HG47rV3yRdhJOQI6WGIJF
1Q5KjSWYcC1+KIdG0UpzuZ24zNxHBCKTPyu6so7QboViYQn8KnLuCtTsrSsBapm9
ZFMlS+yT57+eY8tbvWXfkgbAu+rnJjaPzFpkY11msWiKbN9Fg1UkKoJ3a4Kh0DsN
9H0AlhbAeMvvf7kkzCn8HvrbW5kfy8mSNtqW78eiEmwF7zqNaoPgwqLyVSyEf8MB
Ad5jn19zyq2kAl81hsj1e6OLl36iYu1vwzNnvieQOrSOE7ePePvYyh8gckRb1jOd
3Dur3nwj3jZUUuTbu8Yi7Q6HuCJlet6g2D+0sO7VsQ7samqxGYD0Q++44KbxDIWs
sdts6y2GYqNLEW2FUJ2LhEXETR6xGz/3Uga6hjPbwmfXbwz21Vys0/TFUj4TeHoI
Px3hF5k4KgZ/f5y2ofBjuLAa9RVyIEj+S5bwa8s0lEa+Z79265QRvCouXnFxVQe6
AHGcqTbTqAgOrSV6+Y2lXigy/nlCbgYuhWtLUgFrK4xyFCrNlZHJytiyJoy3GA4Y
4zh4VOnGB2IFcqD8/aT/AY9gizxK8pX7w0L38EZpGBZ1OKR0UaNg9AR36ZMsBwpB
xf8GVMd0FkQcWrSZF39owwCbSaY+93MoszlDLvtKtRLuhA2mxDgFvGh+ou88QUue
tFIHbrO+SVH8poBpu0TWPnEJ+M3CkwQxn0Tx4Nn3h9Dhod+Rd3UHy0WacWvwMEBY
U3LAwQCbZD4SAw2IJRBJiuHrbif/G+TOnzFEn+oes6HXWmhXSMvjb7RJlhPDEo0x
buQuzIcvchKLUDK8lb3iZi3JpEybKfDzLDlf6YF5LNCApmTRAObGwQ2umtLBbIHG
Nibl57WelmMMirQsZsdT5f+wTpb+3KJNospn83n5tQL/2kDQ8le5n5+J5OnWU5Sv
hVEHIxlPSGovSEhAlLyDSAs8NMHGdmW+416SPhYLgpF2n8rW9TqBu4f7Q1zv5I6R
Zm7qq9KkGwCSWHfOekYCFrUUEs71lD3L0Fvc3TpUnHnlZ1t3jzYchKsB+2ylQ8P3
pwvrJMLnXQnC41zPk0Xi91NNv55eFrsfzKooDQkUH2PuG15AgccZE8XAqmth1oSp
G/6V3bk5BasVhpzv3gurOQwKRFT8iEEFZiC7XBrMTjIS88AWaOoBWZKOGhO4e7lO
oHz90pUw92DFwcyh+B9ils8RtEiePbtzZ77t84bZ69KEfujeMIgCTk3cpU1mkee4
Q7xWBuowA79UzvnyqafbYUMr5RnnDmpckrnDqg6I/dqbreR8Up/CSA6fMWsLsTQ7
UPNgrdlDakthX/DCYoolfjRKDlZkalem7nJdUNKPI9RbhNhca6ZslmjiviETuziV
ro2E2Vr1gJ/ZIlG/FcdbVYpQ+sf2o0llcYjqAk5ANA1qCJe/3Hl57sDQbzxPWXjH
4+GTCRF24pq2pNfXW/zSUcHFZb9jfnbgZq0zHIQzDdgJc7I635gyWBud4wk6w8o9
QaqPcGvYaj37/pRbL6otjsTzt7SSYbMNQWKAraeptWA4xMrbs/8fPKc/VUt291zG
kibQjj3ZHwkj3k3YO3Xg+8zLcHjGaMFSkBZhAV0hFOdELydC6dMIqIerqbjh5czT
eJln9aZBbMB4if0sWr7Dj8HlzU55HbuAxRWNx3rM84Oxha3fe5ju7D+ExV2J4kGT
Sm+2o+cMqfKj8LxEAMx6DmHE3+BF5yybDEbp2E8YDmjVQmIlx5s0htv9NCpjzJG9
gZDdKOEDWSbatbL/f2tIj0/bo3IxRWBfSYTlGlhWccblPkyNU6V7SIqtDWvfEFSw
/zfiZkdvWq0UlTFTpuLKeEs/6xbNXGjavsM2dqpFwroZiYsak9iQNQnHDLKQFCKe
g4rzLQW4yIU8u6Me2LGUYTfnJcQ+fl6uY44nNtvZLch7aGKihhm4rvhgOSrzOkQU
j6BxpQSfdjfxgBiUIxJqv3T/7iucU+E1pbxyp32KpIuT25FABgt2PXI2+fyfRHGR
+PrBZEJg8Qo+Xy8hYlSHeADaObfy9J1zfEQI8p3FA2tE7AtGPH8z341uSRQdKfQu
hagI26PUQwSqL976VfVJK1udoEi/8vjuQpp26ng79bQJ62NjYv9ABPAh8SZcrqLs
DMcfhr0CyM22smq6Cpii128bytnTsta5vxDQPX9mAWvEkCtMSOIDMCYc/SYEUmHF
4Axs6Hv6h7YaNJryaOgYI06qvap5E5HjEUAj5pvPwcfbDF2lTGSQWZo1mxPaTO8r
fjk9/BWZNpj+IBcfZUSSMfSSq9MlNNBEL0wjz22JqyqLMjRT5Ox3rsb2GmRivfLq
ZVRJMVIwYNVMD/x0zf+feWc3dmyhwNeoGYZbWzpVVzuKS49YiVwu5Fz9LASLagtK
yz1JGHgvzfOOTidVCg6EZIg8ynvSWwj469J8YSEVFVLwAjEua3KUUr4Xy2Xln1bM
tHVD1Th7Cg2SDcPqct1oXc5Qpx2592lqF05VdPpaLkKyxO7nPYqjwM1P0likyB0U
PBricSC657pA6yFrITss3m6ECBBHO7mLYHjL71T9zpqFhNBsLYYBPCpHvm3SkhdY
Ah0hpJsw8icAsJHGuYAfTdDxAApxksA0hC3XNvBNcpvPXpxrpTLieDtHVB0LCaaL
kFkEDyo2kXSPjD9e3Ml+UK6PfvzO4hPO8nJUUnpJESCVJda/T7U0s9wfSnuUyWlQ
qp2AKivPqMWdxpT5DBjd6I7V5fJ6VmZA53Xq/zTmF7xf8IFargRryqzx04hf36jd
3sa841+x8O3hZ/h6K2J3bw6YRn7O0WWzB806BEk4nUGuJU91448Hm+VxYWRMTg0n
IVUKsTL1/GupivhuRt+2s6smla8vSfbwqaJ8M/ZWfwQzEMVPkvtwb6tVSlNb5Vxm
EiSPR6Pp1SnpTYvLWseT3O5JT+vpEfI8nb7jEjTwv39Fp4PHMqHrY8/Ld+03aTPn
15aPyVdBnxT+mwW9YNdIq73mMmBVNRHz6hpGXw1PJI6gTptBxvituSGf/fefrtrl
oPwEbZAhKYhtv6PsoSardXHUYHqLRHJ1yONZOYbu7Q+qNcK7jo1qT80LL5CJeJ58
8NO7F//lOXiFg0jtfracf0fyjIuFitbzU6QGtZcJ2Lo94pJZemHchWctfF6+w0M2
7lk8xsigij0CpaBbAU88t0cNukIqMDG1/w8uORLzY0pg7WMpFC4RUbJzryHA+OSd
/UMHpRAt/vnNADCAgtMUO/ucClTHXogcTWZfbSNIonky42b+iqQ5aYnUwBO4ZHiS
Se6mkfN3KELgJjkHCy8Cffenb2MgEUpID8K6v8yVEwBppEaJETSjdY+tWhPrT+gD
ByOGRw1FPh65eaoG1sd/FbHghf+xNRrk3FT1R2rrHVl7zcc37i6stAH6HwR+FgBq
kZqcuOhTfILmU7QQFPYbYtWMS/LuFe9BtJevaFvqUPV8pO0IIjqIVv4YnCRX2Sjo
RA+kXmB6MRs3mIX7jq8PlkZSsrpkhpTvx1H8EU3wRk8n55fa+FX0hyOqvw8rK1ue
e5xYbbAGS41eLBBVoQiXLazPRyR+FcPnQPyNHci+K7LL1lK0Px/yh36iWHabquqw
DoVsMA0k/rXjENqfOmeV9RK4v2d9Z/meP26ei2huFbRTFlF2gVqv0Xua40x80lSQ
dW0D4YU8i+NhKAbSHVT0hwBAr5JFAeWvd8tv0scnGX7FRyPrlgbCVONV0cw3UUnP
fO1ni5eWqWV0s5/cP5Yld3r4HDpuJwTW+z6Cr1DYmRWg4Rs3y28dbJQfwnNg7n4T
qQD7Qjug/vFf8VBGxuT2PZoltA9dPogru5/WyukXV06f62T91TJtOc33WNZt4cKe
zA0y5D1YjFvfd2DluyO8w8phHA168JPEuaFDp+q8AOgb1tKdgBvglVkgwMYerzzc
nH5+C8qXurmMMq4DZR5TqJicusaCIv27lDegG5jfyJy9zVEGdnNGXmDGNTD7AfK6
suWvNO4uoV5HZCPWwcchUOVVyIbOBwtyt5fyBfNFOb+HaomLjcDVwuiL/SBsauc7
S/nW4lI+RKq30XNQtMYhObW/ITrZC/4XjxyMZzgTSv4Qgyo3bevAJyA0qgB+bjCB
hqB6EDjuS8btUcGbYFrQk3qWJRHxOGnqvnYlhxOZNXTePy8i9KlJqqbxF7CtpslA
Kw5DJfCJDxir0N9nH2s7GYPuTDCbUuRqciZNF+A2JQ1WHkJP8gDNwJnTwuBT2OAM
3bYtlFQe79BXhfF6AaDxNjvRxHwWXdGijm2wuEM3Rr5BAHs7aL1qDhw5rGnuWXB5
gDFv1RKFeW9O+tiOLLrtaKHTp2AMegN2c6Hxmykxg7IcM2I3rsIMna/YYXLBpxzE
QogPIOCbsP3YgzFhubzhD6aIB17vbtLDq9vSaaGPsParEnpi1N8H4TGqHWJpz+nB
gfFdD2sLFZe5b/I311lmMXbq6WrxnZaiPHsaoIkkejPFT6vJqW7Tvhr/oW15O7YB
GTYOv7HsCXZvag1aFPGuGoGJWys7Mz3z546P5jC7sBNUcqO/9S8V7Zvrq+S7dsRI
ZTfZVSTTnntGZ8wM5ITNAGhCq/YKiKaM7UBkowz59UZ33Dr0a2Yn2HuMcgC4C03N
ot2jxhjwd18Ah22y+JYnNzUr/tSgCuDBpmLgnCFfWL8d1OYA4gg0HH/dNPMj5IOX
g6VQKamzGiTHcR/DYg8awFKcKNmfeakcnwMBCo5dvsZHParOJs/xuJOTr67zFwLP
8Z3dqhFzBfMHTn64nETO152UNgJxbYXCLriLr5aJjPaBSzEf6xWGCiVWXTffPBZQ
IizUzxmf0Sc5pVB1nvJUIFJLDPYeGSx2ctiQLnG72xOO+rkwQhv6LvDyqa6bY5VY
dBjksp31xDLAfXE4iUNGP+wZwY+uM9gVxJkIseG21Ry2FtDS0yNGS1w/+A3rpHyC
oM3W1PgSEFV3L0w0iu0J94s1zypJT0Tn+HupkPK0Ea4s+hA3qu0ckN+vZ1+QPX+z
mUBBcyow8+J+AG+49+aJtjzPvyH/Vjpf74LFC6TTeClOTBLvnj+ifLVrCslaLxma
k3owiNPr7nTIkz1JVGt7Bq9+DNZ7RwM2k8aMggq4JECmuBN4YPXAqbvMJ2TuwNaO
y2LR6Ay35CaqtMmiKkeyvzDtbL9KWR2pXX1r9wcKvq3ZnSGV8XFA0XfYgbQK2aZT
L0lzdlOsuESsIFd5XSYaZiDz6FWzSvztp1+SM+fEEM1KNFWQS53EvBK/GPBtih78
1YFWpj3oFGeblQYOPQwAJqwPQc8Qt3exUwPFis6UGsWsh2pcP9XniEXKmJjk0rFY
RYWTTkM0SnRIJoA4GciDayWkz2t77s+B5Ccfo5OFujjKtpikwYb+cVD64KBLY5cW
IibovmjXfwfJ1AhZz9bRIORsqKKJzMn9OQ+JfyxV0g0hgfErbVlvFvWVQefrC/TV
CHiMB01Mco0/2x5KT2qnToR8784pSmpJ7eIh5hmCAKYDVNbeIA0eMP9hSa+1EVrC
UUx2neK8UJUjW2W8iNLUEVEPMdnsTyn1OcIybSg002mxECqPSkCRs9iOhy2scBTi
AMWR7wgk5QJ94AM5Vjjcnp7xDHP5ATJY/e7mBMsqp1z/0zJEY/wA6g5J/CWh5BPU
oE0JOisN9osLfaGrte42f3pvm+9/lbOkhCY+Z+3xZ0YUicK9bJjokkNgAkmWPnwR
ES4oKoBfvluFt0zPJdiG1wu/H+eLW9BgoH5ahOydWV/l0w2TSYCsw9fhaKfHRCKw
t+HSRt77liVC1VK7NdmtGRWn+zMY79XHmLlglzoHYeC/nvR/iSNFkfPT+kzay/Mn
f0f5wkmXDzFwQk8p6ebb47YSfmfFiqj0+3zoRZwQC+o1m7AK/0wZENxf415RV03h
JPHd54hN6d+EE02g62qcMKytHljR0wuVHeqJWLWW/EDiKhk3+jCvwdoX3vaB+xfP
sA+BbjrHz0dSuVrXaGPXkPZojyUuhbjQpPjIbpkryD4D37bMHrAZhPed3KQarJbA
Ogr39/GwcNFugEdm2rkCuGoygo1sWzd/NuHttamLG0GuGNrohNkSg+IGg7WRuHy2
IOw4oMVPF2TmUk58IFZbvi7OIWVRX3iNyDHw3aTWnEOzFyXE/Ujej/TY3ToPWZQB
DzRWt/wQO55MSSgDLT+5iVpAuqFJmHxn8hBkNIttP4RiiD6DSyvB3Dhk13lEW8W7
JaPTEIz8H5gfDucYLRHytLljt3f/WczUckXqEBdqeNlcReUPWDwcEnHF7ZdMfbhL
aCAcZsBVVz1eaL9YMuRFLhd0phCChTtA8sum+JZKwBWGvzLKpLgWdI6TyzHaPlgI
hwqSpxG+3OIPcCeOpxNB+5QMc4LyLHnBiJKTSIzNBoZM0hxy6HyI3ESN3Ir5s573
d2K3c9OFHjoZ9TcOz6PXXd+tjJ1Jaafr77GgvDx1rpwXYAebeDjjKZpn4ywfgu3y
QpU0TTDGQCTjNCkfVD2g5XY4Blxa9U4oozx5KTYMIv0FafFWaws34v4g5TcngF64
xKYPOBuyablV5IXqL208FNzehqAG/CToDkJJgDzG2Jx5GpW0mmbSsCsFXSCXmZ/u
IcMOPPkCMTxGV7TuaQs4JgQUYvlaMWp9Q6WLSAcwda4CetWmWH1cHOQbTFs4KP8Y
0f3yWS/5+RiPVJtVICvSirrTLuvRwo5OHaLY8GH9Xnmx6mZsqrDKywE7XPEu9mKb
1G/FzR9bKnWl2hyZ3mPFs/ebXbyxavceedlmqjHbRKNFSWVM4CzCn3QaYf5vQr+8
PdoC3JT0+MhWcSmuZgSvMmAQ/rAYfita/AA8KKuJrq0dqC6wqmv8oUvvULu9kR3n
xoBef6RtsG11Rg589k3b3+cOn5zkvaUQGQVY/Y2HiSDLxoqtp9aea+jf/+oiriQp
Upt8GSTCdylGc+nwjRSqUfoLTf6PkjIMOARkuyYfRISWpcHTPhd9IHD8EjcI+H3y
AS4pmmt0V677IlXf2n0+VaUckk6KZitxU1FfU/19y3RFofrH1jluzc26IkGpGn8h
tTck96AvN11hq3VhtRHX0xFqOfiHEvvTQT4d4AfqxQqrXeHbqfYzLYIWctMrdAVz
sLyCfP9bQxwJU5tepjoBXDo+Vce2yLQ6Ff2S/igfX92fXNT5ZZf1ko4dWzKjKRY5
+zppIU+P7EBzy1Ei9nnoCgv/rCV9bp3oVh8AR/lYjauBn9nLifB0dD6yWto0Db1t
qam36cq58tREdDrIjGD5fjgNp9g6hhFCVbRgAQ/l1v5a9TVjJeTLsheBolyqJu1i
mzvoIUS2bcUCzplX1Czj6MMkmggnDw7o+z1Nk98pFwLIV5n1pq7gCWYXGdcnAyOb
P8shNvnZWpdCbGjd2sE78blA4cwOiaWZteKDQENIxStiVCwx0ECbXZEDJA5yc+DQ
TRl+DlnPMPLdn3AKO0Bpyzwj4TxIalty8MEbcuxjY7p3bspvoKH8WkeKp6ZIJBeU
D+jk2/93AzTVN7uhO5TT9kvZvpI+cjFIAotn6hS00MlKS/x0jSz6I2mM0tQCcXL6
bAwYrqUuNQwbi+V/nedbiIZNQ3xsEG5eCbBjwcB3P8/27l1zjcxsSLrC1/2hYdJG
n2/VIjEFOl6b8pVKNkOnJtLILvPnzktQCaZgnb3y27jOJg1wKsQQGvYQTOhH+qfM
g05MG1zigxENvaEhA1ELGtDxvrKLHhs/Lgib/tL/TOgYpK7h5rU5qvoHxuaYp3hQ
HpRr5LCmPjRLUUdu0XspgtFUVEIi9PFANj1BrBcpoMj1RgPxQ+Pj+tp/Lr+IqlAZ
FUe4Fgo/2UODI2RidsNazGknNA3USX5afPN4yt8zD0H+j2LvNIziuU8SfemKhqVw
E9mGZ9oYYxXFc+qYOpPm+SiGP/8TviEQj7Xn9qsnB1IpAgDbKZCg2m3jOlpVA5Al
wTX25G/cyciWmouh1GNHCIzblyMw8G4U9Wr85xd2WIDGz//ndk+ckhz2DNi6YENl
heIvZlhgmw4hzjtdbb07I57q4VwpUl6LNJAtMEhI9D+C/yl/9SFVFZWDd6PL4R+0
5wgS4AEx19JgFPzlyD/bLQsBEL4+R7dzGr7nZndv+0Q2WnBkx5T8spcpyREB27Rc
sxpEulPqlMpk+GfrzP0KoAjqPmgDjVw3+hQjEZAyqMLSyrZ4B00R7VEk+BDdKx8d
WYA2KGDsrgW6q29Jk+R7xXE2qQUQbB2J6BvTFxYStvscSuS6t78vmJIMWKZXWPHm
y39/Y/PKbsxAA3LnM9Q4FbQ0O3GknkoIqIeRgO91Dkq3yrDdm7IgS6q1xaw7iry7
JAe2tK2+QoZg0ji1nv1tHICteBbbhDbep4RLH/H5lTGtkIko++6uj1yWSjIKVynG
VkKmQcoIsx3K0+vNMFWCl1pmGWjRATGgM0hC7uu1rvzIDmxJorsbrsMbkPK7OIku
gLJsYW7ABipUyuk1Q5cwPSF+Afs61w8N4nnwkNH6y/rzC72RQcwdAopZygoK1MqG
nXVn5vSwTuWEITVu3CXfOO7hU9H3deMoLdV6rCbVG8sPvrZsdflCY11nBC5lA68F
aLxe1KDQ4wRIyl6Wy9C84wMrusdZdqD4ekLFQIiTzmB9jEXvSoO0UGA7lNh8dxFz
wXY7fT58sZLFf5HZWIZTpAylzmf2izF+u0xI7x8eP6q9iihRL/VMlQi1yBg7/NEU
LWBE+LylZhFn3eKlpDRtZX08QtlgjshRJLbzZyEfHF5MinSVQLNlUe1aMpaXeJRi
WzGjuIbzHI4grnYboYOAk5McDsspCx7c0OpVk3YWc8/crrlJDiSmJXj/ZjZ9YoEu
9ogmCyVjBVOENUUrtmZXyKFp0yvuuxgy8GbdQhre63ETiY6Sdwy0bqmYleKPfoin
vA1b4Aablc+//hLJHbmzfqOfUgMO843OOayXQ0Xj2IkmL5pSv0L64AA2Iv/QZCIZ
EpT2yZ46oOIJ84y5NZF9C+FqiRcvzya2wetJ/1WiHHgtg2WgGLAy4kU3XcWuDLsd
+ZqxQ+GjB8ASBWzb+36YFDM4h+l0ooQOmYuEs+0GmKrmmqblNp5yK7sSHrAZVu2T
oGBTzn76qd1kfS3tKpGbyA9YvEezJY/6/luGCuWUgZqvKbVARkcZm3T5dGNFAwyD
eoqUGoU5zjmIeDk6kkbz9jcbK/OAdISZWbtuG/RURaRaVYmKGPUMHMnofNtZpaCc
Pu1y7q/0ZO3lccpgXHR8D2VvKdL35RJGe0GP6WYp3YCveJEBfaZ8dnZnP9PZiP2i
FF9HTw3gsR1bkqaBCeqWmaRH3pSk4/0atRoOSGx/tYQUl7DaKdC0xl7g71EsvzBz
F7QX6JEQbiK51uKFkjiG+pEBrUjmRH5aN8EQsYW58Tr4EIMVBGIZKh742ZxGtBzi
r5E4tnQrZRClfiGMUWPnDQklIMbPWo8Vul/RByRnC6FQh3lMyfupbobFjIxeitwo
9KQHalF84HeKCJVaMyIIdzQB1Rgk8H73MYQbIWDjJJ6x3qBB22FjUSOBQRgYLAkC
MkQOw/UvxB2CnXJzievuPNPwVtAseIaO5kDWwus83KdxZv/2Chi/1fEDmRC9D2kn
uJnqLN/wmdEj3uEebCoNoKqTb/c8KhM+mmXDZH1U04pxnJo4GEpaDcx3Xs3nig5s
nUekm+IG9tPJdrBONo5jA3voSyGmcd5vgJW6DCPCexQ5zha6utn0WQEH44fIQcCX
OmJgguEmYZkVwSho/e99dRH2VyHeSrCtflse2zRLA8h9UxDRCRxhQhjqlloTMWa/
DVhcV5T1FnHuTEo4e40CRc6QrJPtXNQ9+dq+FD5BNcfFp5ujtPHN+kkGNWVp59BR
YgdTeMi7hWCa3Gigc8urzXC1VsIfpwKCu3OIfWexvBpcDeAPCAG6Ukt6ewXSOaFg
gUTMMmTZQMPOuf78IDggHpCWfcz3/2Ep9oXP7fzIJ7GYWZOqC+vDIeiiNWoEh8mu
qo/t7cvluk8VGunmkEKcT9Isk+7teKEjs1Ayw9Bik2x1RXgogLCH8KwwqzfGjmAx
14bJE7/a4svplT1EpK3AmM911oQzTQ8X3+6HthCDKajrDO44EOAqbx6EF5/NctiN
1DXgRdQfAUKvClpl/Wl6lVspErS4bViShVCNxC5K8ShamBclPgtJOzaOyDIitZJG
CrGhZ467IqKOHpYy8Itu0gP6sAGVSvXytmQO12ifbb7y2hlN1AEhUMSYA5rlpzS9
Pem5XoDlKiO1zqAyOwpPkDpvTvXmTQivMhBc6eIeHxmdiNnX4qMTy5UNQuXtUriQ
a+ikgyWTL8NFpRuvURCx2ktUL26ztLSIBBsppQtPsG3hc2TPCTiSRj0SASCgrT4A
n/4zVobfR5Vc8tmtGLk7y+QGrdpCpPJ07GKbDcDF4bJdDk7obKYvw6fel8GMC0f9
Y46LP24p/gq/KYF+EHfXWmv0AAxbkiUo2O+9Oy6AeUsOP6AnB1rq1ftZ8J94l0WL
nesOuKiEU/FZ/w6ufeTbEjqaxVL4Pxap1IMr8o5FtiOaImbl8wSdlEg9V9LmoQpn
IGyEMhsQr+mZHZGsrSStWNQ2PKIGm4llaeOIomv5cKjaF6G1zXdcgEWUPSHNcomh
nrWThazo0pDxlAbS3Cmha1O2n1jwUrS0ME36Eph/WuisV7XVTLHZmTbjbXTpXB1U
gCFqoqtRD0cmxA3CXSsFcrEFqpDpdFyVqwp4bIMdnlbQj+XO8lBBelQ+gZ7dMV3X
xcWPQp24Pq4i6br1sNcObDsH+lXchGRGUkVjUZvYJN4rK8pygAHlKnLLfgMZGwj/
1Rh7k/p9KpvcXCwnqh1hjHHnTw/j/hCmhW5zzvlgxiGVnDWmokFpbPMCbpFgL12C
7cmq4bUE5MNOKn3Vbr9mnCQfMrFJpi3MwOBGwxWN/7RnGQgXX8XUSj+no3ecnUfV
fatkKQ0fd4BnM7IFqVna3zz1jh0GfsUPW0SJiYP7aeGSHrhF2pmVdG7ui311I+3c
x2FegCZOozN859GSGgyoNBLI9+CbTKkqPrazZ94kOp4H+VCmP5UadLTOgGKIyNex
15S42G4waqjSifpp/BqVKbtVP7rf6HD4MeaBFk+6zS5lCjztJbMbQLeBbdyT7SeM
ZG2kQNxEYFYGXt07yCV/eh8EkZDh3o/6YLN4stSWGTIrSIZxtNRGcclizVi9IbhN
gdKtBHJUO3vOBjTG1dXCQXMyOXydhT2JKYBpuLvDKdgpAvPutut5SKDnONvFw1ho
SpdtYHAxATgzEt6We6QvM8JbWFxocOyGvF7O2ckUMhzEnL7XAVUidMxjyjG8LDkJ
BD4EnzKVhS9uxkdmcupfTUxQcb2XQyLHojfMNRpPqGySWOPkSYyqPUKiUHxZLeKe
F9HkHuFk/yuCFwQa+dPPfxwCCfoxfHNA8SsO1rf4GzcdfvaD8v6zp82Xd+mxseEg
UJpWwl5doQ+/4VrZSWJVwn+suK7TRoVXdqfLj727g/xy6oTseBvASBle9aSa9MR9
Fhwwma5vB40D58i8dHc0SelxgWaa+K6DG9Zgqy+KM9wQfCQuSc4xcX7sXlTL1tDx
4FQqycBSX+xJO+SirVp1qqFNw5NBTSY9O5OiDxbBNozxMy0l6GnCt6nyuP2NtZt4
AkCYVUWyDMGkaMCVooX1Ur95DareV3wj1Uf/quZFg5vGOOwPtNEKeWqEhKUZj0V1
3blVllgpv00ZJyWzgRqkihDGTHThmLHWN7bxgzrVp7q5LL/gC/ZtnRqfGWcnNpGF
yeTxkbQzeFRAyN3QCU5vm889LuVG+WDGOapmv3ZbpihaabYykuqANKHwj9j0NwFy
lbxCoqPjQzRNrl7NGCzbYnWO3FBoqxbWEd0Z7l16mntjlNkFdTVTB0E/oVZp6grq
RMfiH1YMSKPpf4Jj6klsNAG81SlMaFFem5wTLCpC9O1GIpHwPLq1+9pQN63wL+Gt
4radNl53Qk1xsZC/KBNEoGAOHOGR+1jKo02pGSW615Art0NNM/F8MKb2EEFpukGm
mn1ldEJ5KNYmn9KxPPdakE4lIYkRzKmKhW4kYB7IUn7uxB8wnyELsP78oUaVctD/
RIw5cDxCpAk8iqMKps9oxVGO/FKqf/eZ1xBXmj4AG6ZPD53Lyz1rSHINLxjocTga
RJxQEFtnPHf2aU0stN618Mp1NzOPYDhE+iNDKd6JkE7sGF1lOQKhaLZSePdI10fB
NuiaCc6CPQQR4oqd70szc/36uceEuRKNH4bkurd3rgjXoIrk14K6A6sM0EvBHoPC
FmYwXgMuM7v++3KhT4WIIhZ1FtUVu4/3rx6cuxbr/GCXQQ0pcdnOdo/a88HREnur
SxwA+Lx2IJBWZ8RF83Ca/1/2YQS/nzY8zXfMRNXFomuLaWbkqExda20RpiVJINj7
N64lcphohGhQJw/su+T+WBYQgUlQ+ggJeWV1YARGPvSAh4bL9sY6g8R5vcF2uVRx
+BeGlE2ZXv1nR4Cz7KyN1iM0Dh2ne2e2DClI7PlMdrINDeBZajHHl2V9fXkVCLKR
a5vMpPwKp7zByCcew7JQR0n/kvO+tuv/T0WFA9pW1NZ4iw6+hO/jC4fg19suDzQd
XA8ONZtjqdPaNW4P9ieuPegR3Cw3YgVMRmJc1NpO9T42guyKUlcYeP71gF1ogElM
7PoDolzVvvKPfDRaGooLzfVBMKsGd+58/N7WMYM7FHjOEUn+voS+H1seVtXwpDe9
17h6MylG2I0Z7wks31yhtsxzcyARg0Cix78saWHlHbnnHNRr2arFtZwgYDE0NGNP
tH76UPS6pFcZvKr72Namm1hS4ZKW+iyqHuLRZYB4ca0h9CyxWRe9YckgCBSetZiU
77HrIi7uBkdGH/PXjG//6Sla0rVI6o+dwrj5wcdbqNUvUTKcA3zzst0DZKtjeQpt
fD/Py3tkFABVcQfXl+bAyx91RPvr9UX0sCEOxeJp9CN3Wen9o1jTJyvMhgHG6GYZ
9IOHAVLgAeoRdIpRTqtVd1HCe+wk+vCl1BYJLiGsEZtjK6nDFZ8NT0yBwOPwHOeK
aOlVKUYUGCd2YmVr+aIYG/hD9k9HqGtWlvbMvCPHiG0HvOgKGPNBkg1djWI28iqV
Z0c4ZB/XV1bIdsxNCZz4nnjcsRj1LiLv4P3SxbGd16dG0Z2PeH2kHMdcKKg/7pjP
2/0u8AXtx1qV4czg/qLcr77agRUrnse0KtgADCE8HFua/HropITgaDGxGl77MAzO
JQyQcYdqP0N8nsPo6vq+lsy7/nnJRI41mcWrlx2pP7a0SypROw0zdV7QyypVr6+W
cnUcCWEhDgq8/4S6ERQwfHalwHomFVF15UZm66Xpbp+MiXuDd/hXLkKXi4AaXCqa
+Du/kL7EOZVL1UaPc77d/VXUYJItKJO3RRerHBfSAKffoUU5BNQk2fqN1N4KtSvZ
DkOqrZa2Ae4Uqgip3kvZfAvE4+xNs4Uao+0VApaFGZJGfVlcXhLkOWlxpVHkPd1M
ER1y9xq6ehEjFNryHgRU41vv021CuiJ0zSyW6BeazOYoTueS1agdts4JtiG0MfAL
0N9Ibham9gVTpWaFBO09DoYY9lqKRIdrM25ZB2qGf6nkpWIpApHY+4baBXke6NBY
k5UmX4kmi/LYDG71CEra2RVpU9q5sRowfuBauDAAWtbG3un/+mqFVTl39rXyt6da
PYm8BON85lMSKCWZ42aMBi19NSGVDo4/DZZqupKcMtr5zplMD4qPhpSbXY2CTafb
S+RPEkZ1JIS/NXnub8lgq2DS561YCmMW8aPcYfbSpornxo22JwmrdptEblDUH0nl
/uL8xZavgi+YpxFSwogNgCFMQJz7cBQghc2RbYruqJ85JY6VkN4ZVtukr4byeAUN
CofSJ5Q+AHBVPo5MpBHIRw9Md6rmKOafpJZq0uTA6LPLXRRP2R+LDzzJrRyL7nni
NYlvoQf7rgNBcp2nUo+3NPNCiqYfrt1Eeq9v3ujyKS//r2/loZ2TKuJkSFDMrY1I
kpwJr2RZYLLxWb3VGW5iDQS42xjp50tq2RCzmdNBOOAsHRsG9eVzAoz3nR+WnMRx
7omp15+UtARPglkokdzMDBzTAZvgUpoZ3bnNqNjhvWynq6K0zoQtdIcG+EqjszZ/
ONVwG31vvkChOQ+nfRqKGhknEogc16HB8ocTXy+g66ncze+7HrI5ImywmZ0sMGQ/
ErKFT6PjcA/p+Z/VQ1f5/8E8Ad7OuXjhT8ZMPfObXtyAVnDo9v10qIXnoUfXQZjy
yQhl6W4fcaUnJxqi6h/yuIP6Hcj2KatN8FJSFIGqkEEDdQhEuTAgiq1V2AjnGAcY
xVGh5fSt8QWlNnwl7FiXcCPtjs0Kl7gNuKerKEL2OhQAJul+tSAZYJy082mXQJ4J
aYFU7EkUkoYFfjNRlVx/VYX1vOmLWf9q9W8+4D3N98dAHNXGimVDEiK+LzfT9J78
lcbd1j41eqRfBteGCqepv4GwHgmNXzYH+lcci402xktp9oOpOSoGunbHEVB3wWie
FST2ubg/xVrM+qy0Ot19MCUUPbq13C9DCWu4xsocyaQR5fTR+UQIois6WrIuRiRq
Z8xbc6QRyaWVm/8D2oBloMN4meeY1S+jLnz0mgvlz6ml10a+rHbyIlAvE+P3dbSK
BjtPeBdYRySd7AzkxgFeqh2z3Z2I9Et9vH243CMs7wqZubRT0/+lCQ7Em9sij8Kx
tUHmSwsjC7Atoj3UklG0ZwbcvVoWfIhTrvG3/s3LypBQNHxaZFKQxoUtcuIpAo2F
cXkq5LO2DkOyfd3IvACXsv9FZDn7McUpdRolSWbUnIpbVPz2RgDHRCu2CcqdSQ+k
fZ8D5RIcekT/pOJBMJUVd92C1AffctkT9JpjYak70T97920eJsfNUIfrkdJILjtR
INWg7K8pNJs35YWaPD5b3XIZgUyTye8tkv0r+YgR7ozOxaeIWl+OohMnAkyJHWFf
ArB9M9ax/wgD5W/Aal6X/OOESw2Fo/3jCwR9qbR8lIIvUqUrzGC04EJgE1FzwwAJ
+TbFlCrPV97SPjPaRJgHhmHxDxjFYGdg+U4HKKvbhgtUmnP8k2AJRVdvg8jVCNAO
McdYLXjL7eqmTESOmXC9jLio9ueL0wfU2Jd12GaLBb52bbHr8Qi6wHo6KIIrAJ4V
5fZN0Vb4/sRFPQ7da5m37MzddpAR68bjFfNgecmwDLY8WiL2aEQa7c5qCTOSqR7i
2vOrQ1vTZuLLYzWb5QU/DX6cEpXmjZAcQbT6LNYTA9WgvplxujsqlBpMzjUjLDPn
GWMxUMPpieo8QAvR+qGpGeILdazLNgqWMpqmUcX8fulBxsixsIRCVEJtCggoGgVn
wnMQIOhcs5yzn+4w+bh6NnpBnXp5ZxbOu08tlbaGhVtedPTPsaXgdbbjxwV6guYR
RWrCD8kOWTLWERlkUO55GsNR1/z3CYm+w+nAhxtiKpBTBSzgmdo3P1bXfedje/mN
VTz8tK5Ov5yRHkOWaOS3wOmXURBMdy3MLy1quQNuOuKXAx0zIq55LTNrif1U71sy
v/tnkhCNDYl9qXyhMmXvFTFK4edkUBMj85GLtIYzeDRezr84IK/8k8CHPR44mpP1
tolRxZOfi4sLA2lv9tLNdvk1ILfJRZvmWmiQYsFlep5Fw4f+yWaiK2EUP9E7e7K1
HE4mRe+tnEHGEFYkFjtxVCyLfszSS9iX+ga8QJUnJb4GcLgi/u2H/39Pamni2kn7
ZGxm/3+x79yCcrWuYFEeuXNOrYKHXR2ogkctrrg+DW407qDchkZTxLWAbcixiKL8
i6zc4k9mClCqmSxKG7Uyu2Gxc2H0Jv6kgQLVYd/pctJCr/j7IL6VAZUyC2q68Xvs
nty3RqyzKUNZFlaZUUxIXO38Mkq5hSfxqg8mZ3o7v+GLn/RF9gqP+bZa3D//+2dK
cp1x732oWdD64nhgYXNkWPqaR28Q0pFdD/fuEHAghv6hFfPOtfLbtuGsH9PGUSKo
+d/bGpHFc+zV/plv26RAya+DFYs3iOwK4Uu2KNTclHB2DWxKh+FShup3QHCnWjmN
wnKv0kwNI0dtV0sSaFiWJMs1LanoxQEH9H2O/T35nlINpxCheeaBAwTGF/OclX6u
0OPztgL7hlDM3HwlPm01CDdIQE4JbmxpJaM3g6vIgrQp1zJMAyDG4jnkYcrKzbUz
GozDHInUyHzUJ2v/wRM/s11eDsVCiMPIAW+ZYHYoFkn6w7pDBsBNly4Da/L9zKgA
bE8i23wIjmA4QfrEHHJPPCQ52tTBjVIapJtV5iqnwl+P1Y9kYNzZDnSn8lJ3U8oX
BRb9mD4isils201Fuvyks/WlWv/YidyaCLZ6geb7D99gYljYccxgcTDYDs+b12ay
BR8St9yKUKg8A8DpNyAZ93t5/jRvVn7a4iRXOig6+dmaxDlKbocqkTW33ww5pi54
pQDl9vJ9h641WkxT9iLRdbaleQKK5fDsBAlWMFjz8FO1vORci72nGWl8tr7WpUGK
5mS4RKgE7F3XBVa9vvlZO7733/YetX0g0Eudg7cCtrMms2ALP9N9KP5M+BcXje63
6NgfUdrrIeHicNfxFUEhfs0dBl1OyFHWKA8OJ/d4lJjcSwtZ8gI7ERVUuuuwP9CR
xe52h+BL/t/FgzYQAp5kiW8knKQWdK0P4StnGNUSXgYyAVKPrIPM6md3VmLFmUV/
Y39sGxYcPLwEkwn0H2PI3kaP7Mi1i7EtiChZHgdiP2YFHugd+aq3UTXhNH36OnH+
UhHUdnfaPbgq37gV+cgmdbt1NM5J78KjfTZD67ijU75hkS9K+SA76fh7DwhiIB1H
KXWByduyYfs9zMFX1jhrp0tXKk/4ZdW2ASljnOEmxXVPaifXFn8t5UHqWyvvczBt
wQrs37FdAdECHDwNUrCMXaNALNBcBw+Jg5xTF6fsSZpy4zUFzSSYyhtFpkyNiYHQ
RyC98DIyF5KHtIUATGXySH/FZC6uMZDpUU+T3AJZk7LQgAqwKYqh3ur0jP7MRRge
vQk8nZNUz6s9clkHIqEaNP6peoWSXRIJ1mGlxvHFC8q7xCputOlJHGTWm/fZ+ALP
5BTPOwfzvEToK0PU9fh+EkpopY1cZSvWnrXI5+PFUNBNZ2YxLdocCBiGmavN2R0l
vpsvc4RTc5gLbxSVsimEeEmQ7uC/3Y2O67m6NJg8wKkczVP5pnASgLypG/p1L/AH
0xIkS7ZMEec0UwsRhor4T/xA9HqZKlo6P7Tlo09mo61XWSRJ9nrglty7wEO/Du2a
pUs3QLL/TB2jBG8jVWX7OMGC6P6EXcYK8qBSs7HMaNO71I/SHPOS68UjniLHQLj2
89TM/7w/Qr8cCGLt4r1erXR7ZU/mabFm8A/yeiFJoWpXKizW6mE8BKw1Fv5SirrQ
vwD8SurCYLN3VVgc+fi74QjMLy5eLzXYvp0PmK+RevKHIpCM8nN/oQdtWL71Wrg5
M2Zz2LHMCyHaWfviRPeOlc36A3DAlD4ssrwWhH9TZJ8dHeicdBhXt+y2i8Vsl3Bf
Uo58MrX+EEAFzVX+JIA2WP5HL4SspsOUWUVmYl/4PwgGkEdtU8nlmKhSBVlb0g6C
631UQKsEXRVoH9Mx0xcH5/XAhxAaQEoht2VCMD+XSCSJuYyQnymDG7sbKw2Lme3N
Llao5LSLzKnSbBff5YtV0u6P9lUtxen9rm5jB0gy4zeFEnyPNN7ypXccNasMHNzb
tCythEDqzykyMKBML/rUtKdAA4gHykgrSuOUlg5lmEgb6s7El5NDuTKrHvUE56BK
fGpY1q0ALyGF3H5MDR8p5GU1yhsQyVj7sF1+4gmhjw3gebRQ3iyTRSeRuDmsIMFP
FH1BQgK283oFBrCjxUE+wgdrFfnxvwemP4++x3mCBGfeNfZS6HNr9VvH5ZDITlm/
yDZoHCxwW/izfpf6ZKxRe2v9PrIRcCfP9C5u3/fPUBFPJlstYCzPD+pEW/8CgNln
00wyAruNifcZ2SDP/84QpKdzY1dYuk33oMuP2OTuMl8UbFvARNvpJzexBEZqXguT
3mA6vGfQ5gYP6OllD/8BJUeuAzKHlAgtJhmz4+/pd+LE1GXtERKQqYPP3W63Cpgb
/CkIZoVWtTg2DLQV/CqNOczr6DgqL9PvzEo54rkmNvwCMcVSwOImCwpyMc+JZEQ+
oyCxPR6QfK3FwXENTN7NAGtrSa8+Fl9l2rc6BU2gr8AiBYk+Zt4Pv7EtnIdi5Zt8
v5iDil0pHeCnDGWT0hNRdO98RRN25e6e6Mqh+aieIiUKKYTIWDAOAGR9BNZg6jN/
eYh2P/hYtsui0PyXAMOOJ/ePZ+mn9+KCVEQnV6Xw+Hq/kOr5MQ1XMfQSCg1uMhd3
KFaTD9XZEBMVlsNh1HmG5Zzef2NhFnoEKYEfgkdq5pjSxtD5xfllM6z2gNzJpByA
YQA9ErmnFYolM9tighmo6QJZHjefstEskA2IGdQlgA63Q+ZY3Im4+mkis8Zeci+b
ZoyEAQQkFkWuX3plh6+LzipEC7/HLL8eJByepHGndrDSSqV/muOFiET6XOAYBhzd
7EPEQ5SgC729uUh9+f5B3W7lDjaG/DQxVxrQDf2y3UNyPor+zyLeGojgXpzV06h1
0swnpn60OjFuC8F07+PxkBmR7tON6v5i1T0IGvsdske7YAkFBbWoa145d5iDG/9X
zzIsyZpvfFJWYtONFeX6PX2KnxQ+tmztPNMOPkdPhq3feZr8qTUiDxDslllF71qM
Lf6aC8rqsz4+ZspvyD00f0t/2BaynICT3zNJU4tcuu42ytWcmA+h2mzv/qKH1W9Z
1bIpsJsjqXo0naeg8mfh2c4eR5EzoRH7kveS9OirlmodAmVEwrtQQwKjr43SCg/A
tDBgHhIt7u2x5ZMSMCTsKgmW2mO0PmP9Cpwi2Kvk98LXfH+SYWJqzdj+HU1tnXd0
Q6h7GfDG7y5XHNFBr1f7ADLn5BmkFK6TaXsU5R9n4d9xM7j+qNZntMngJdz876xv
/CSS3345wPPIfigBza5x2G311ML+HN5BrP/4vwxSBAh/3hv6TzC3xRYLBefkTSXd
9KcRUzDfjxGJWB+5h7wVqHIssVrDylJq2lTAUd5ILiFTTjjFJGL3WGODcRMbjba5
a1Ws4++YuBrJVInKRvqA3jihj4cPtrQkNWVZTkZIdfjxnKhyoCR36FQpAsx0JTs0
waBC+UPmgnae9vNLdCemUSggefKJfSa2L9JASiXtodWA57kDOI9cVRMbdjkFDhC/
SGs/Ffv5qdvPqutFWLjIIhAntaxnFkXQI2n1n257oVRPMHuFv0DCF7TP34p8n/qI
1PmTTMQTtGsWW9WkzLiHgbIQx4KQXOe2ubAvwXhVHZx8PESMZaXXH571jk9lV/4x
54JmktKYbxPE4DNRETwwh5lTgy3WmZ7NDQFNOKzJNtizYHQePlmBr3wzKg2ASOr+
0P0Y4FMtARJy7B8QHYw+GwOwOWIR3UEVJBGVqJ8K7MeTd7u2s9NJw/K6dwJ2K+EG
rhz1PkZMfEE+99Lgeo5AQbCZJs2yYfDLZ2GbK2IuFWG+NPVw8S//px/sy598aLRs
6/cI1RRx7tpaH0h8/mHUb5ng31EBarrRYCVq2+TFgvvUN7CmFC/0bn0doawt7FVD
B6brUpZToru7T7o1CH06J8aYrCxEecBW+Eh69eNJlsINwjsZ7bCq6ecktIzZbf71
5nJjhXaXBSRIyESUeFfXRKLxZmbmhaJEBc0bZX8Sz1pFifzBrdj7RS2gpiz35O2E
HvCsQtKqQn19GACYlE+erKkAChe8CPEsotmwJb9qb+Vbcwf5cV0zFFU5NE8LSPi0
KGttcGxVvQZH6LT1tZHthW2YLwQIrfyz3vGbqYH3tQyo4iNDB71Y7WCXIav1iBjE
Az66VWg0BILarbGgHFtzbWNW6Knea2a/pEd+q7ZRlO7MTB7MzFI6ESL8jgqcZ/jc
kxcdeoK05hxNOmkWfY07sRgHIuQTT/qKtZjh1klIBjkj5nktmpAXMRv4CTywbsBW
MmNZv8itSXwHCbxo6LmffraC8GS2jrzd29uoGrdgcElCyIScZbiPgFjwCN8cOh/a
FboQXpIGJgUFfiCFrBaE9vz6jJ0XNLZ2+tYJ0t/SxMyCgVa4meDaGlHo+adGmVw7
ac4mw/lI7a+T3wVHUvSOhTl5F1uyNDe5ETwGpDRieGAv72m7kNKpYkkKgaruQrPn
h3Hh5Qcdj7tDyn2BxnC+7N3p3WiTS8cW6cpvJEQSHb1E+mSgi+l2FPXvlPk6leJZ
MIpkyIQWqsQHJ3m4gw/cQnnbJ4uNNFffYThfP/B5aqjCskivPFaeOxxin6WmChBo
lvWTQ5XwYSYMMX4KnBH4iakJw8nqfrioaU/t55/C4Md6rvkXCbk4y434zzVzBTy9
un9K8fmVAlOOpZgXBWZYENjE5q48lDzvqxUoIhdvlpwemRGH6pznZRd41kwIUrpG
Y+oNzM7huN5W7TMODK9Q9+hbIyG9sjy694ql5Yl5KGqpNQDHWci0S4SNGB8UzduE
tNOzAswa/nzp77rtce40G4N7aanWJOwfShAfEXyAtwBmOrbiJJiUyDS1O8h3WS+2
PlVDzYRYo2QCP68tzsrwM7tqLnROm/T7f+1h66/f/ebBwplgX6yPqQB5PBFFc2dq
1r7jL/7QFioWtHQb84/7fB4M/6H3478A9I45jMW2de3/jSB784akhRErJDBtPP4Q
ICKkAeykcI8gd/NAzDQ/Hv2lfyuWP+EtKCA8iMgS7NRIWquE2hRIenMwYKWIAeST
GO4HOcpQOpLuVg1L6v0SU0cPG1lUIegliMwobD0JzIpJLzlAc4NTaBwOzzDu+5SU
xCu0A7GiEwk0EgDgx74P687MZYfhLccV9UHYQwgk+0IeK10xEGc80Rymt/U4giv+
CRRSOPnqhnYE7Dxfe2CWSpfJctyAU72cP+K/q9rqgcNlkAgH0BJ4pA/ZIX5ex/WC
yBbZud/rFavwJdbZ60ZxG4Dm1oVfbo2CFmDWCsFn6eF4gfFm7/+R0GI+Fgoc1KaI
Sb0jbzW4EGe/R5fVIFf92wTICVjRywYMubDBC3//SG2xYfjs+VxoHJw9oPDr2Wrq
QVJo0NeEtcgPqgmHkVY+mvTOpbJECS6P9gsr/St4xmgPeWbipQ+np0CL5ZTCUB61
esGaeEsl7abtxi32BETM9K4rOhG+gokFNYJsV2JZ3ExRy8Wov1Yp24wqi/uwOULi
T/zIQj/3+3oD4ReZi1L7bXbUeqakSwY760GliWTo2GjJNwu+K09LjWdeyAXuivmQ
Z9kfR2fPw1FHSImvsymFD7xhQAtIUsUb9FvU2PXthn4UztPN5hdAFiTjPOWMSIZ2
EiQxlo1x4ye6tvyG/wlZVepg7Nerx7FoTYXFzdM+3Qs25kdZ7+M9LncOY6jOTZzF
EXQarBSNWPcOUK+ioPrKh6f9vjz8kn6aSTjcxz6yUV4Tvw5KGiDznCBLqzBylXmH
ckKjYXLzgxMXTYUIGzvxcfZPNoH5OpqpgK419kL/fWqyEr0pwV29Z/e7/8I/dASL
n3PGxg2mQrrO1MUGt9sIM+Jlw8bKvyYMpbaYi7SZ0LgRzKNO8UkpKgXIKSlnMj8c
A/mWbSSq5CSzzOpaAngIzPqQFNpVzClEogjhPzIBuRc8JWWQaM4HvcMsvx0SCw57
I/i+tENp3bQYM8VAOC1drM1QnMdvYWx4bUC0SbMJ4lmcw50i99IfbQ71eOtyBcdB
SvYb/fJx1FL9+ovnbyuafmkARIcdeSrnufnBGC9LwwsdtgABnf1SO1yOuoXqqhlp
Vz1ievpdiobR0RxFkI+kdZnmnJNhd0ZYXqRnBMNUZG2HWk9qcN5hk575Hse1cCAv
ZyyY78IgXoJBUlnxSs33fCRLHmaZ/MhwMgnqryGKRwBFYS1C8rs6mcS+K1VpJUC3
PXS6gLvIyXxHPPRCSwnhKblyd9z+vuY7YJ0HNzeOeexGSDyFVLCqs428Rf2jXFm4
46+eAUzYyJ46xK6WWdecnmaqroE6Y/XTd/EX/D1trRdDvbPUQ9hFON3TOU7twcY6
LgmMA5rR1uYNw2PK8OIFSGdj/jTVQ1RaInuVS3lY9aV7exvU2fGgyixk2oMobSgm
phsq+roh/HbxzbzplqoWUjSvQGAiAdcV7r5IjEK4BuclgYbe4G8xPAmKK5mEsEzH
E/mUzDVw8qCI0dgo37tuYtHobXuyTojOovm357DIvj7uxZ0DpSoLhERarz4tc2Hg
ahAwnztwwwQCfTDr/HWsMCFGGsu2ZFqolLwgbPE4KKhFiYGSlhLbwmBTdv23AwtP
iq4ANM5fdbFL+pJTiHgfRLy8YOJIWJ8jxDBv+Jf0DUZJhp/TGJpdkaKoEs7Btdu0
3YYiXUxl/OImlaBSiQ6frwCLb7se1CCG9SKzyq8uxxpWNHfjFyaA6TfKkQn0bOfG
m73Zh6ZTVpki5GrsuoHnvNS/GIhUnAjCMujtlhERN9CuahrsJqskSgsjt501tnge
UsQJQEQpT0o59uTl86BP92lFgavtyZxWZMNvUhlUab7E7E476ptBJjN/kJquyr1Z
1itPBzClXvSXLVW92fUtowSegwOjLvCiU+VWA72vFqjXRbzjWgJsSZg/7vL5dy51
t9a6SHlVGajYVR6mCoJlSEPxOXHCpu9ht46GVGBESnC8XIHQAOhjqzqZ7LVyPHgI
2nKdnKtz3e7gE4vbumuGemHWzbY0Vm1pfaNEdhxcRQz+/9yZGrsLJA4eN7mwTR+8
LFYyHKl/8lAk1xBtGmaT9laqx4XcBUH49dSgeEQJ330/Wphj6hoNCzWEc0I4hQaw
mYMO/bscHxogV3KimoRqqQpVj+X5AJ8YDlQ6f3T+RzATrQgUkkPI/0tfCpyWB09Y
AggKtr6QRHPYpKBOhFKwjH7Hmw4Oz4LwfWbZv9QzeW9plFZRXlWQQdMsZZDTB/Fk
zNMIgHNcDIieodxLAfhji0qDbamEiByPZGwZ/Jx9MVcAyOIuOQRfdQFmubhKTwWL
p0xmYhv9tK2E2zmHdPyrtp6bvvTj55PNZIhC3wThpstuRhD1Qf21d2jBeyD7RiZW
i8UXVT/NUJvRcWs1pvk05bKLpXErBafmYzyiGBwMLbV3HjlWsWyj4Cv/W82u1vK5
gZsSctiUW+U4VRdBhU9Cd4WsTIoeks3POvAyvXRYthuAxui6O2DZTYuy9mF6T7vz
cWXllbb5T+TDT7ERiGgZdiQov05fF3G9PU/VYTuRRZ8kPcurJMrahaeAmC/+O5Ce
eUOkFCnS+9kCCfMxhGFGOkjFRs37ubGDC3WvJ4GdpWITvgywpnCQ6d5DXngYq4dM
FKEnYoLjwj+UjhcMj4ZkC5yRDH2FMziXG7SWh/Sil5koH3h7A3cLR1mtWFiR7iIF
Aaukggtud5TAFca3fD0gLtleJaJdoE9fsGtXcEUOdenHaczu7IpnGQTHHkqCKqDD
hYU2qNan9hLcnlRMaDyU0NN35qe5UxXk1EYfketKd4q/JHGSliMGncNF17kPOYF9
GYkESGtQV922pSlBetza7VWhx9q4qYSr7N56C9mrGxSmX/kNaqlirgDwZCawJyjp
8qsLXXI310emoiIxnLyfWWOdlgs4Dy69ajv0tjVSRftt5Xxz1SJykv8n7gb3eGn/
1JmW/daqAlEo/9ouVRs1sVK/uv8Jr752OUW7yNXSn28NgB6fWHyhFJmVWRY/bELn
QCyV3/1BeHRu3BFzXxPNWRTNqPdJAMyzTKNIeOcnw2hclFpBqN3p89vXuUq7Q4IS
M+NRy4l1+igK1XejAk5IX3WQkkHxxjfFpZm8TEGdOSzfefDYl4SoQ/7WBYeiVgSd
4gSex3GDQMetTOVgrQrpJdVcLQcmx3VZMcc4Z7V9TiEvlmbkvO+5d2Baf2V4iK1z
dd2iux8hbZ+qBJ9B20pkzJlwHqOSNo7Ecse4GOjyUK8nrfBDk/u0wNw5orkqDNQS
87f7i9/k90CfI1CLcuvgAsBJaCYaY0nZAoPjB3nUF6VFacIdBTlhg3o2nOrrhywJ
mcUI16E/FqppB7/ZXZNyhD2XIb3IjHdoYnCmLuuNlti/yDv/xLSqvqHy23Bz/Ucp
fuq8jblJ3ZPxV1tCr5kUao2i/si/Zd4LCjUxlYWkuoL64zcjtWtd+7y3bhKmN0gE
+HLQ9w0pJ5IsEexgmu4kZgxKUeVF8DMMQkJyHE0BCAoEuDl8MFsFkdcLmxe4WQSb
hzPaK8XW5fkDtBQn953y0x7vR6NvwjaRdz6Oqv4R34Vwlc121z3jZt49N9Hi8i8g
JWjhL2aKfznxAZpkxtJLu0wd2qWRrSHKzvD0s8/tD57euV2INdBb7y8f0+A4uIpR
uVVeFpoaHxiuyeVn7R8gVf+oJP2OR5M2n+bmxY+oKQD4x87s5fY3OTp0qOpG2a3R
tv9fnJj0BDRiT5V9Ip8NNJ6UhgRh0sHxWilkw4Un0a8AaYjtqojEu4wAoVFG1eC7
fXlJw9PzFnUNcQZCd54WVI6MAxVyD9Le/uimIU+3IK1M7SunPW1DlB5RcidkGSRa
T3U7rIolE/NAAOyXWyJYgMhF481ZCCpnMnlTj/974Az5iVJOX2kp77+DybrQ01vu
bUMlDBBKARtZdeQ+T+ug8OgWsGJn0SV1XPVbfdTQO1RVpc/pvvTuR8FyYIXg63r3
71FTxJZuWNpSRHTfIDCZnzWOBQm0WpD5pMZDeO9lstaDPNjvQZYq3fSuDLcr/PMK
ku9IkVdb5eW0HknUj+BoYHj8oK/7ns0bjJumGVkjOSRLIdsRW6V3snSqgfOB06/Q
9ximQ4MzUPxB1G2hV70aVI1fXQqEufj9c/WwyzQq1dPS+5T1vJMdVMLoG2eyKb7h
/ot5dSDWP7yldIgTb9dWxxXuxVtvzuRKaBXKxG5dS1k/e0CMxwfq79j3jkeSSzoK
QRJ4Tkqy3GSD74FV3I3+UJ27wzTnK1waKa9tJm/r7TXXKp53axPsH/ziifZ3Y7AG
rrCYBqBlOJOwBu1BRi70qlm5UGQFiKN2MkOtp6N50ghxqwC+rUj10XmOkHpptyO6
mRjH19p5LICwb4FMGkqhKQ6thAJhO7yrWDSVRK6hDX4ehhuN1fdXtjWPJjgBSX3V
Miunh1NhdPnC7naeDdjK5G0EMXM4dSAM/Rs7x7wnCjj3rX36oo8JsYBVlVyXFp7b
WqgGLxTg8oaotc7Rt8Et9mVLJRFG8gt4GDWobEEChrq78XSm16mUHwwM6flKqcxQ
S4qNhnALR88q5UKPO5vMGB/T6IcOWEbu6gjFS+Zjj67aO3UACJHf29vuryYdIsVA
Cg50JPmxNUJu3RA28O31Tl+pD+alYH+4lIJkw7W/wC2TaydQzgBxDhBND5E8qX2H
jyJRIw2xKKUdPvX7ZJBMllb5021HvgAPSVblj6j5+tJkk95K19BuBl1VOXcgYvDU
LqCCc7SpOSr/KeQ4NcLxTECtH8aZverj46ZCeaXCfGfskULKlkqfYLPqOE3txgaW
3B06Uhb2m3rmloG0deJX9E528q3dNhz/O73w3Jf4rH9kiO5ZOzWxyJAr5byZ62ce
Jka6TBDxWWmaIXfoJccbJ1hQ0BNnTdOL8zaZWg0E8t4kH4g3vMkcQlDS3SZqTuw8
sdXBX1zzH/uRq57NuwemRjBITFtzjbz2qWkDI+x4464HgQUSLZ+CZbNBa7Kwo1sn
a+kQTmH6l7UcOsM4g2TPmRwkipke+pOp+kTK3wGjKNOUZVDA8XycwgoaBtFYAmdz
I/bkr0+C01jnKNPhjhTnR0sryNVbk09QTi0Dcb0fkdXVAGxuD9e/g8zmwi53TrYO
RLjZVZX3+pV07l54CbY4UyiFKirE50/bUYfGwkZTXC1XYKZQmzr97bQcYIMPOghK
Wqy/I4HYjaR4EMhwQA54WxIsENqCSkWDhixb328oQ+P8kgI7FztyayPT/LnhmsnL
+eCXCayBUgsanToGzc04yWKweL+RiiBw1ETQ5Lz7DEqZuD/Emw5GUXS5+6O2Csxj
E5khKSeUQNV37iiP6EaCCP6lxbdc0HUBFCcFD1pcU05HFZY9T8Dzgwd8jUYKRpUy
YNbnjU3hqnNmkIFgWkW/qj0BUO4c/ZviZwCtInkybg1BaDviavO10fTad9C2q8/r
i++4fDdfE355edBj3NuV7acqmRQgBsJIpb+Ge16qBIu+h2uUVbsexYP0Qijhu/M2
aNCXdLBtMDJyBj/7QKob3TinFCcL9ICSpY1p9r/tEBYMDPf66YLgF4GuTztOCYSh
SOdniINWBjtctrmzZ+ODGkiUqSvLp3nzlumnZmHvbgnGnMwjai7I6ajRm/VZDSt2
qXrhr+lQU4U3AD7InMDTGVNpadZgM3+eC+d23Z8nWH48g+Tz1BuO+4of5hu/PBFd
9B5ZIfYtMO0gyGsa++ia3Z+um8FjuZboovL4mFaJY+2dcEllXvcuxC6uFwkx0Gcv
Aq3fiqkN3nIjmvzuyOBgw9t44wdoucdQoIWlEx17gDEnhn2lvTR9qGjLtLvRYUh2
vOiJ/gBg/zFrsx/8zL35581Nd/BKK6SW4X8p+eJ57zTWc/BlvW/QN1zg92kACd57
fhrvyisg6EgLV6HvTQusie8bG0or+ipIdi+QKKQXksBfp5G+BTTPKMv5HGzCM4PS
c2zJVUvF3JgqavZHWmeNf/KuRE4m5Llb9fkcjp5CUJTzn9DlP8i1xQV4yyw5IuMR
MtZ6vDhO309trAayH8RCWZzhN89sHCj+5aTAdqDZrph28najD0UKxnlu5gloCuEC
NzsujF0llL3gKxlcgRIamROoZSCfMnlTmTCY7tjx6kQFRlj9wbYxlbm45gDq6bV6
nAe1Zh2dtihvlrNhgmVLy8uaCe/9sELJjKPj04lElB0bEN17+Fl8O9C5+XL1Ajf2
OkdOku9m8HhOrRh5e1pqXKVEQz8/uKkZ0L5zEjeUSreM9ai2+z9cvFPiWnxw3ruu
Fyu9xqQ2dBj7Gj5qxE1UTlOEcDO6DmN1vLIE/fKvYQpl9Spzsgrw337sK++TNsYx
zemD5/0GshjL7FVmeImEY72Fdx6hpSAwnehP22xFMtoC6UZRKlPT1xcnGo6DEFT3
8ZG+RXepr3G5HlEOkf92Pyq4docfG7Ml5eDXN5rYcFgGh3hdByImYtE8xdPPyULg
BiNNorujfnnHKKEgrd2YoBJHwyHJOhDtB69SN168Cm1CXuUha0URYuLeoRY+/EP5
H223sQbYu6v6jEbpiwyZpMvqVhyhS7VM+UrnQtkLkpzZHGCVzUBzMIzBKErBeJ+f
A6j0eadDmma14vReD7alEfFyaT8KJAU2qYBxkIK3Dp5HN1E4y0xttta792X+ruo9
RSvpwOUsNi4FLRJwf0qM3zcM4ELg2ZGUdg0WLpb9nRlRav5cGghDa0GCp1BqA86j
+We09la8f6cVNPoxOeZJQe3qCxGoBPg1liKTrk8G1JhB+RftaoNuZRxiboUv43LO
wl2ehp17JIp0n5BfsSRF3peuSDKFIShZySYSoybrKhNtXUhPiutzJeAhjXd6it3U
HrYOc+hSwe3fpw5b7fdvK9ID+fs+fJNs8ZWrKNfb3pdswiESdVcVBiJVUxwIAKd6
AenZjsnzxDQGK1CTkefSvT4Yd0MRkfsDq5Ss39Zok+kikacBVPiN5HmFE8d+K75Q
NU2tRmm6qENPy1yq+WMT/Gt3LaJAcCfoIpLt+mp+bW6yNtMZnst7rfhPAMloCNcG
GlHS2NpG3G0dnUj3PxSoNotCgigp8OxB31incaySdvQV59mzp3QN+bq2K5ZaOSZ9
frqwhGaPPbZro1uzbHyIN8WdOTR6ntbAoatxYr/h4ibIxqEc4bD8Ox0uOGzQoQZy
JnAR8qcpD4KibfcV80axmsUCZkE2vu+e3AVFLbML9rSSpn9OTVumYhuzTzaNIvnK
z0ESL7nX/wYN9cZ90dtb+LV2yOuPlzCoIm4exDlmDOHSGpMgLg+Bp6ipQpLGVfA2
wwwE2KEkb6bI4q6gSrdwQZP/HyFw/bHWy+tOZq/NRrbLcOr68ZcUeGW/7cdQt3nC
hPcrnc6Kxoil4ymFjDKYfo1cPi5uD+aEmSyqSAoEIekGe6Eq5Sm8YFdMAOlyLfTr
vz1KC3Y60dWv3QM1xlqVrZCijmjusD+oNZ8lRFiN/a/PNePAvO9VrMjU+p7odkV2
aVHbKlkpL9q4Y7evUxatREbbTa9pDC2rq4h+jpsM6A4wSU3oYK/kZmlysAmu+DwT
ZyUexutjC6/VkDj0M8VTkKlCwKRhL4LKOLCcCVG2pxajHgsBDfWmgOFgG+3dKnQ3
tVoFa3vX3ccwfw+loQB5C0dZvwGmqeBUpBE6O2R+OV7trQa8U+o6Cb/KDHa/1mT8
MuwrqyqMYhBxNJe7u0glt0eovItXZpzKBDiCVXl5WdIc67E2I68UigW90yEkCB/U
WBqoUhxEya3tuxNhnxM51z17qRKyHFUPeZTqsp6hesr3x4cBlDDlLAEYfQZBm1zD
f1apqGV/5B1fkyhakjB0HMD3FiFpBA9gRwFrqlnAPtgv+BkXe6JoziqyU5NsddAK
1r8fgU72UlIZB2zwYNUAU+JS+Z00ip7DUyzkCCg9QNNWd0tD8ibUaDD684Ra6XEe
T7Dkv6nD/1HPMt4KW4u3E8JnvrnOxjkWqx2J2+y6u7R5TFgMLqhzGlgbo6EwkCqS
f64iq84O2czJMTb8C73YEyo2Bp/DFJDCOiTlUkqMvPnCnl6+zmTwyve5g90dX/OY
9UPODRW/v+o/fzFii6BF5W/Pr2za1s90n3IvOc52Sar6w1cyJWSOIgCDC/N90xmh
QfukFJ++1lUlY4q8Lk2Lozzm97QT3owY3kcmlrCfNZGo0ur6JSgiK/lBmWLz/6iz
deeWsDzvyB1QJqdNtxdUIY7f8jQ9uvP5ra3+QWFzKsv50872thc4ZdD/9sJHwhzP
HgbwbT20aapdiRtxPYa4giGl+caeaqAu+XKKOniLvUBY2OcEe6p/Mv5Agx8/v9F2
Gki6T1/HQfFR3wpjyL5CCAVHXEYbUijLWcbt0OPB0jv3XHT/F/97jWDlGWquVOsT
rF9+pg4P1WZnOtlQlJhw5rcMCI+bClNO3zoSuEiepw3tPcPCqOJEPhmZNx8wxmKG
8VJzRJSYEappicJ0rwVKkL1xF32a2jYoRykdLxVb30l+K0M5qpCac/skygnzqWqc
5zmH9QV+kSWUjgOnjDXwP3bRvlPs8IaYo/b86RuszFD7BZJ6HTJskKaV3KESGMbT
J8QlWBds3n5W4iVFGbJm2EqA451m6z1c1kZoPlAcJ7RCxPLYgGFcBeROkL2H7e/s
SzNAW23ycy33tr2gPUURCYTs6sOZwNFnQR/qqiC/BJ8sFn7ixD+s0ejFbVd9ySgA
1PstaoHy89bFLgkxoJlFpMUI/IV8rSJrJb2kAF9zCTvFgXo07P5gmKogygi7sVtp
ESDS/sovEUOL31z/tiOMs6QGVFInpnEzIFWnrAtHSPQOJ7wirEGcuDYpPclaYkso
kMPCg29D9pzsjh5ruSeontKZ8mXDyanBHWllvfxZSj2pDRj9ITBbu7vTXC2RON4z
jZIXdkwQDlzPsnOgzCBZ3ISLWSatJo/mR28G4j87OlRQ+rsx4ocLOGei4xhZfkQp
9ggS9tJcik4oWAGkPGY49LOcpgS5z1OEsdLcmOK4e73DMPaUDJY9jkbakx34Bc90
O+cohzOwXJ78A2mVkQeinHO6CYYkultFsSrF9F6L2fIaRELvZKjLJOt+w36Z5F8K
4YR1K/mpckhSuv+Ga/X0MWR4jMtXoXvOORSYZV9Wp4mRNl+3qzYt7oPDIjltm5Yp
X+dxLPLdbzjaIPsogCsFiDCrZalI3bG6wFg4JJ7tfxlE9fBvGtNXrJ5LgecqzOvJ
dvDIRtmZxWrITxKmC/lUhUZ0FpUzhpZ31BcU3vK6AjphOgaglrXs+ZWbJRp7ymzO
Sr03PZ9QhJx0WV6FB5qKLsu6YFZRD7dg4TpbVBuvkbGL+4L1cK3Bw4uTlZ3QFkB/
LO4tHs8uMhs9nXFiU6GatVBlYVs+nZIU/7RJY0JCJp8q/jhFGIsJHBjwCeL27zOV
FQ2r6l1Wlj18uqIFIDK+pntBjlVyx08/UX90vBHiO2w0oXLAwfskLnlrOLTu40k7
2oHpbzxTuWdH+3+NOIUhxAu+IeGsc8AbKocNgpLte4jgIB7VUZ2Cq+HSuJGEtN4w
imLyDxDE8UkdQ87De3zMKJjGTVRZ8iJtIHTYBUPnQsLsV8tqSiJPMdy31RL+Wf8E
Lg2pO88n9lQ9UBP/pA1lWpdJ2/BZjjmEDarbY6MwnHnIWyEAEVJsIRInNVTN8l2U
g3ixWeFUudWQMgRWeKlsTS7UnKenzazFhXWkEgC1BE0wmM4TzzH1eZTmSR052Y/h
QvdKquz488Dw8ioY9oicw9FdRNvDr2LtT4LJTwooh4rWLI2hdU5KhJ1UUzYrnihJ
pALTQ91IMruScMldy8je4DHQBPOvdpriC5LvYcY/2jj3+KsxOhig3HhWLs5eSGKK
WU8gNfzyy89wtjXS2swhFZi8v9deNMu5HQS2+wbjiWMK4MChtgwEr26oZevEmCXV
Fo6GRETW2QB4P6SJj1qI+3vhZczFggqemvgSvG540lJnvTYsdxRGT2k9biLRXavz
iFTj+7ncHWnMZoXWiAtGw/UxbxLJEXGFn+Ce1EzlmnYFjQUecVDhavwApgN2yLYs
XhkzJahQUzYL2NiBx+PpzNxN9nwoyJMJ0MNfxDChmPfAd24WwfK8bF/yYoOKjB4n
AXOGQY0ETDAzSOkasnnbrsDVVxtgf/SSVxZkhogKOTXzOBctyldkjFXyuySW4qcE
B+vAnitlojsHOOBp8OIPYp+Y0jSDRswcoAMUpE72bAMgBceOY3QJK2h9/HhW7J+W
p7EqHf6GUktDhoG0ttCQxt6RydsUfLrb75Cav4ErpahPXQXk2+Oc5J96j28MIwZy
XwuQ6ACilklOkY3ecH91pTh7iPK+Mp/MxpHE7n+bftOJiiZKMyFCcZ0nZR9YZ36b
f47uTM3lQb+vQowy5qEErFSJotCIQLCmSocp9ms1creaRHnZrwNXN7TOYJQ3cUJW
rkhQSrmD/yl/dZRBZmx8cqCMtp7FCpNiR/6zoJYkmsBsQoRmP4PYbP/gepcnhr6H
oNPDs3Tgw46e9yt7BhLXMpzX/blBDW45ZmsHW2AAXVFFyEg5rD/+En23irs/de8S
xSHMKUSWD4YwTtXC+zFPGTZrM47SVTYbKPW6ylQsWvw4XCYkPkEfY5q5FJeaDzZu
mlVv1EWe7835vfDTBb8wNPxSMmBxUM3yC8vJEXobNylz+VW50YjvDtPjdPk5Knar
YrOCtHTCadLsDVWSZxYUU/3bmncGW3uJXRxnYfG7AiGqeXIbFze2cD4IuL+FcQ+g
tHZMGR9zrp8zvWTuYhnRaj7ko4P8hST1MVfnZFbNXW7VebWG3CKHl+J32nwRBlun
HifEzIvFU1fQ4kSlyOMcjHo96jZvUbw/fhYhOqNRIFQwZ5LV9hGTGRH9hOsMx8zq
Oe1A8/U0h5K3/IwUkH9uDPq8CDFQ8ZRWMSdU5ZMswctNmCZwOa96MXr43XTut053
271uPkv1KDSsMez4o+MtNnRczuNmPulOk/APlJN6KIHRC7RwzV9K2TVhYo8FckkS
LF8D1a3a11mHyJ2xJ1gwp7pFGdwYK/8KLKtV32CoitvABOfGPGARvBj7OdaBhQrm
57l9yRhyUnIJxX3hFVjq/3Cy0lwlMWny+3Qj/g14Oxrjimer3ZYZ0+j447FeXS5i
Fh/jR0fb6JWAo3eAYMDAn8lvS+xUUfI77iYZVf1ehvFFXqfRFtvuY9Nd+6qxSErO
36c1+cmyxGqL5JfnsMf0l8fjwOVdO7QOmuDncqwjnviv6wlll+QN82B9tyfARe/Y
I0JYYMI6OO+kNEIl5Cj6YXOSL1iTTjo7KJo/2Zd5ZYEhH4d7Agw9yXEB1Utfo6zN
Nwp43OWRmCu/aiy8RCZshqvjXcYrKEtAPvhIdEGQwLj9JHqQJrSYEmSveKNX4qfz
m+C4vFF/Sk9ym3FS7/54U/ow6UREO7tr9HJebqxHRMFhhOFAGF6B2YttHvnWelzl
tUl4NusLNc6sv6o/WN5rutVPpMh958j0yS+CErazwiHdMSRfpHv+RhVoj8ZgXMDo
8x51/b3Bm8P/Qyf6IRL+PcLsv60ntixU83UxDvkUmdxTz4rvDA63XZ7X84dRrxup
wrskWhG2yMwcV3I33eDiYEFoEKBtevV/oc70Sc1kPOMAo+5NH+gLpbSi2K4bMvkQ
aXyqXiVxj8VkKQtWMRXnNS+zCboB3hMauQWOHlSXTZbavI/MYIknohdW3T+wIKn/
fdoAHE8OTqla3BArvg+Cop2pyUJF4dCu3J+1ohZyBcRIuLHLSWKQxeWcnzeoFdYQ
mwVa2dbX4lu4zE2P0vp8NklNuylNLgobICBFNm8bKCoiM+9f2vtJbiMVHfTn60Y/
WJ/DRdZCySUTRqnqth6HSvyF5YrtXTFnpmHz7Oh4Nd0vsHrZTuOBB37OVEI84Cp0
D/qLIE1Wq0i+gCGX9GGW2VESPy+/6ZOntZoCIvKvuOjSvlw12+7fCxv3W4mj3g9B
ndYK6K02eBoBAev2a3jKoLD/QgFHdiAp8oJygW5qNVeqocGVW4CKMCKxR5zlUhZ4
SNMj/ZWr+yQN0tZxxGWuokkwyl4rAVM5muvhfetS2t7wqkfSRY6RgILp6hUWsmU3
s/ya6zFvj9FcccAxyQbALWQNQoKsmE3iHIjIh8jQRUk5T1oYV1up0gmYZg58TDis
LK/bXFGdJCmELis/9xxd9vPFGY/Al1HZXW7d1nvfKmJRsyVCUgYBdmyZsD32czyu
y6Z7mivjiDrS9pk42o2duROuiWZVSEpVwenOsXxzjCU4s7cB/g9SZsJBZQnaBxa0
7X2Wdg9sIjdDAkBYz0PwowkRp/I1wUChPqrxvOdUlsa4H9qs/nw3fI1TZCRTL/KS
PyzcsvvUEkrlkjOowN1r86Rij7ktl7tXDMIZyCHzv23xEEz9T71lTVo/Nq3TXYM6
hDvX6+cSvjkFv2FXVTMa90GBDhVkMHgWR7Ccd2Q+8jKS7TNn5Oje3lrOYnH1gj8I
QgT0++EFX1uK1q2qncq1JPVdcP8QWNuaai2jvvB3WnHt+Q5/JPxMgB9hI6C9XgJ7
O4+7FR9xu6qgUiyALaq4z/gWR7PWF3mgWhVuSqrY2qMhJEQz0v1UR9NcyRrCLU+E
qFz/Obzy7E+E4vC9rK4XEBpfqz0NGYq5Ox/BxTto37RHaPkfjqYsBMzMsUVy9w+K
NfkUxZ0suJdzLjGfZ5meT8rMLsLpU2aBHHnaI1XeFQC3aczQgfWyIcuCfXsKzKVO
kwe/0c4Id7x0tkbjWx3lrHeLzQFSxKXj4xWDLgyodWbqk0AxTkmMsy1xNvmkdcbz
SrDCL57Fcofh1IN8gnFvgzSaYuz/B1XEYRJCrruvt2SGnGIOVJKFq758q8halJWN
9wMBCH1fdp1Hm+Uyuhhryokcyt9hbw7JjI1aNo0lNRmxYe2XqIREAcCsrsgJRrbE
lUn4AS98r9IM71SR/ino9U9+DhPjsuETO79BM4ud88Zprt+btKg8tagPFlMZ4cri
wjgCnUzlIMGhKaai8Q1zcKw2BYjN0nsA57+KT32n6WqJP8HU6Ciz9q1zlxqJfZEp
3nz7m+wDvMBXqHsYlYbRE1hI5fe4Nm8vYOOJ07NKH/JVT5s9txonOIuBRgR4iiMH
WQO7Ye9mO9IbiQu0Xy7Ak1HifxDwbVhwF9PwoH7reecrkswQJbdTvIZjhaR79N+R
HFxQzLyxvUH3Gaf8FBPtnEYj1CEtgd79FOsPF6Zit78OZsg10XlVMv31JHa2O8NW
KGhoWgG8fD2pAWdZHZ92PD51bWtLNA24soHhWVV7vD4O7xwbq8GRsYASFsRBEK1X
7tFvEenaHnV3J0Bl+S1cL155zaPGBOqRf12hRnrAXt+41TvWg1xXDXOGzQhVmehN
Rpf2MlSUzyoNaEGrGdNAC73WLuSkV04Gs1bo9xOStdzK7BM1qmqa5RsAWxccIAUf
RcpFDdSiqUav2LtepfW5Ahut7eJLHbKx6IrCXvBaabxVK5vFWIJ5zlgxtZX9zQ22
4t+V32trQ01+0riSYXRZaUoVG3s8fUVYR0B329NMekuPnVlaEqac8+u1E8S9wPgK
Xl1wBOojRKUFQ4v9b4tF4HwGvfL1Zhe9PfHWCgEriOoMgstN/AxdaFwlScBYOy9y
5zfPD2Vj39hfdDid4HiN01Kjhvknv78PBPCaWwCJbXQg+dspjoR5p0KkScooMjuI
vK5PXr/yixZCmq5C2dht+rAbz2C/ZRAdmO6lk0G5f90FXrLdk0KuIT+vMKAS39Ob
SenxEcQ8mvoW9ZtOeDbGNYWWIDtAAyN+dyaNNxA5hvJjo2GH2Q4B9iglSdAUse41
IEsEjema01wyrF5UhsmPx1Ia85eHBbry3aidVT2QYiqpxTkjeskoXtDzRvd/HDiQ
MUxFkf9I+b1qOP8jke+7+0Rwpg1eVmXQlZwBEbLrgCDU+JWzwniWI6KIiH01UjoP
OBmNLqZ7nIAlM9wLh22SAXfhMWFxT/NzXJ4oRk9Fz9YAdtV8wB64Mwtdx2RIXVFs
PWGa7MePtD4jR6eyohzj2uT8E3C9DnH+n+MAdrcf0Pu14uBjXCcC5MaHIILPkpHt
ybf6aVt3a6duYybs/41MgrJwFUSVvHZl7iEEM65A6qOD7s0NIn5DByEgH0bSz42S
MkbswvlYhz3f+F+UwqO7ymtDVDYqQYVng+BHbaqPWuJDb6rMz+Afb0INwZtyAaaW
Qs6JwjCBmpTYAdUKNdV0WPGoATC48LEqxzNJgO96FZFaBqkhYiTkxNtAqw+Hwctp
AyXMmTn9UA9yZdv10rS4jhreHrfAovtG+O4KolSZnyA73JcpmuxLyxDvvQgo+4Y2
JKMYAEyaG7ZhSMwrILIGT8IeRykSc3o9fpf66u0ImcgrahlOIj6+Yreib3drj2XG
djDU3UXirFtTZ1URwiDcKp/oAHNQapy7L+qiuGQzjedJgl3X/8bpOF/AsIHsIOus
fHemJeHCSFD6kMvp1osbfXEw6P5LXPHIYGA88dMLZD4Aev0ihnJS181NB/qX47/e
QJwWzNh2n7edTBgNumRddUpEYHWzZTXTScwjKt7EfWmntawmeAyMJFTN9ax9dSXf
1sI/LBweEvkMvDqUfzmXgJrrNZyxx8ilEkUSnYwVs+LOqg88+rAcyGcAqUYkK7+m
WhXrMKcPoTrVcQ5UI1AMDkuHHUz09eW+NGgaut9n/NR08bJTIFRAzAqrTGkiHDvT
QNive2slklxowE+6BBAt/8Pg4Ii4tOa+rZCBvRXPIXYElNEVXF4HxcA6JDS627NM
KXwkHtv+cVB3cCsjkhc81nty+PYYGXqy+7QyxEzFb1NJTEZwcuy75FSU5VGM1JcR
Rz5oMsOvUabWud46SMekS1fibVr/KIxORgaMKwpyDTW2DSO+uY4yO2ZahtuxvIms
xB5xewdI2EuZ+ARmleRAZKuy11H60HvsYe7as9ZCMLWa6BiRrhrmG2yTv3TXecZJ
U6nacHNnTPOhsg25R/+Hm99dZ0VuKXGMKgm5sbpTnjhApftzRkd7/N3rXnFRRAnP
3RnCbDYj7Zcl0z2f0qPV7PF93cmo3dkM5P3GF32WFLP5q/oSGW27G0+DHjDpF9KU
TrhpsSfGOqzlyFZtheXgDVNuW/hIpofAmcY2py7hdie01R+N8Ojve+9xXLmUqfyN
cCD2AoPjPXSa6QBHZ0b0Dp+newEa5UErjARdXWdsH0KoJRNYhYZ4CaUeLZX20854
FAB5oEYsZxL4VRZW2UhKy0XJnT0MilCXT8H2CJKsnRbuQze73v79lMWNw51EmVQ9
CIeSNGO0UrXbEpgC4vyFRzQwPmWdkBscAYMD6Vxg0qjLU5NWqE4ilGN6ZC567BlY
2em4Tkigmj2XdX8wAKU/M8WjZoa9KYvV007QOLvfb60ii1eRgI9Zoni1n+KpKxSe
AZ0BvPRLo8QZb6kBmRxIDuavdYWS8keAYYQgbaFeppkm+xDPm3VHpwHuGsJm7diu
xWn53bHeeN5UtgQW9gs7SeO5ls7GdJauoLDLz72WUzxNqdrVmhu/R9g2mmBvXD4I
9SYe7oCQFJWbyFMqnzD6L4Qz7udoTwTrg98DikgIYZPUHJ+ZM2Vme7VV4EC0UkQr
MuBoroFx7FE7Lg5xh//pJX0JeS+K5h34I7uSTDdXOl4LURk4bZ/3CNQQsJW1jbZj
53SI3/U9XgnjhzLvWf6EYe4Csa1t71Y9Fprwy51m+PzrbSu5ARGtk1dRfEjhyqU1
VTga6kegQcTku7loAOeEjNWkS+LdQc3V4qTGw7Mz3cWMvtT/qxgtjiSWSajIFIrH
RyHjCIMyzX3+ElPuG/klUh3jgS0Ncw4waZQ4N7QILA8zfodzOX1FKVxSX/Bi20rL
AkA7hc0BKxoOQxrqacdv61ScILfwRHvU7QZMC9J1Nf/E4ruKyzJgV6/11xlQvNyj
nQJS+1Y5JOxQETPyKI4MxamP9ErtBHv/wFhCCYpbClDqzKDe/+n2FOsXAyZ54KoZ
mCAwA9z7XRKruTRsWRnvtHU0Li/mybe+gHTiqySZcqUVVdOVNpcUbcA6SYWHmmLJ
yiNqWg17eAvB54h3Nd8IJ3pWDf32A6F0jYtYo8bOuv8NewQY+Hjb15RpCWmA92fu
YPMSayeMdyiiGdlVCvcumFXIn/u2YPezAxXrhlEAWY0sVrQfE2mDcSJQ94zqDgU9
PVrO8DUf01uKkXnz3UkD40cDxqmEjRJitMV/M/0+rldJ+DKZqejmZsGFhnkyHxw8
kHLn+4tRfHJCgg1TtkCPuZVwLSLoUmf5ClRIVES2IT3vYdC/LbHKhXYFhCoq+8WN
TjDrUptQbLkwZ32sf9+AbVuNfugGuCj0lO2t0UAlVqiuerhE8vop6KF/9eQH9AFp
FzCy6Qouabfe6Sn5nkQWptJ16t6TaytaPt4/YmLZZ84kzVJC9kUSxkurrWZRp3qg
N9DZUDVrM5r5IFC14OLX1OkcA7yZHR5Sq+QZH36sl3TDusxtLM99qxKI6FfHMQg4
Q7lfsN3lr9LelGbA88Ad1M0cmexp6jh71axQqxwIT8E1lYZ/EoXnGAFjN5CNiWEl
Me1fQ2c/ggYLPpu/vWWPqvYY73QRusPlCkALdGIuc73nXc9+uRXD8Bzo7f1kcB8i
00woNvcSCYS96Ceutw8fe4CoFFrSAnoMutYH04PoIMQvu+MbCz9MI6WGjNCcEad2
hu+kGAk4sN2vAhhEKrLMJFCFtD9HZf8r1TkDw0S1f+u6fh2hzKRFTjIAiX9tkHpI
0lwv6zD2pLbXPqpeSJMJbWC8TrZdGv+d/O3p8Zun2DPrgNSzNfNdVYCzH1LHhPmt
Lc2jyXUl0WOLNiPJCZzA0qxt7fJizxiu+x+e0VhvKIFxU5qnNPgV9F/KNsmeJPlV
+dZN0Ft5ehTUDaEDanfrPSvrszGZ4UM6YDRZdbTY3o8mlABReVQxTa29I5C+FZ7X
JUqeOujzjcdKPZ7Yv8ogj/fjLOWJydebneR4hXqzTD/xeaVNR//TBLwHQkTXGa8e
EIsmT/T+CmT8G9jMoM2BwdyneQfT15yCnOqHANcx1HJ4O/SBAHfEv4NnSv4n1Bf8
5D5wpzO0Yfa+l0X8Arpn1+jS9zEujs2ZQdZSTHl145j0msmGbPletXpFoWfIs4YF
uKYBMF8v24SwgAMM1AAW3FCU+QOeocsy/XNts2qoZakJHRvGCjtCdeabWMuRBkII
1Mb/Fmal8/8trIIRI+fusl1JOCSbyAoz5pV2ZO5M2UQabhiWv6CR9PoNWZrxrjW3
QjTU0rzbQpMRYbYxKHR6Q7gR3Ab0CCMGNjlr1EBtXbfpigm8jXSRMX1UDBANH6PX
0Rm07Hog3GSYti+1+imQGTV5m8VzCm8+Ts3B8TBraFhkeiToCx+HYfQX9ckqa/ma
vciYpPqlUHkHrQBUnLMr0rdtJvP3ihcHXnfhh4xck9zHF9fIOzJXyNLGJWSJ/IjF
/mxSBRU5VpeaTnobXXs5m5kEpfkaK7wMUAVLlfBk/BhAMI5SgCqeahDG3SXg67UI
Y8zFjG1qpU2cHTiJYSe0TWsHvAADTEaPN74Y9gBHqzFIQtr/ecKSZZBKR8tlvaqQ
DojpRTTtlZxrvTltoA9OqPIRfpq3KFH3vyvFu2euw4r835dEHuXGXpw8zu/LLJN9
KIamN8DL1hzNaoH3gctkkTD4FllZQ5CFJKd5Q4MR8uvNFYg4mUcG1KM2LmDYEJGL
M8GacRQYn+74r3JPIvzUhQuDiiFZr+ZUrF7AI3RibV2+hvvvRC2KKLDkG13WOkD1
GX93+brA3jcaZHF0ISxA2Mlzv5ZRbKhEby+HNer0SpHEcmEz4sGNqrtcLOamq79e
hUHh5K4LvAv9NxBf4Nk1Z7etgBivekpUdFCba3kaazKEB8LljLCiNE7ebj1a7I/b
mNSwVt1Fo3IL5cA3EGRp6+Iw9wcmEBbvNpyAC4shaQEBQs9GACixXlwDKaqKFSPp
hp/th+KXhlCCo/C41/uvIelGNGTel+ifAFZXU8/cIYEycX0RtFNwKJcwdcUjHRSX
cC3tTltLMFooCrNtUVJd0h9rEv+/V5Dut4uiaN7FZQAp6sLyMfOiBJVGqUPTqy2p
7SuJjfx4BvgNRtvl9P2FIdq4Igi08SzZjr+9aW6AuDMqDs9/CwwMF6+dTn6TheKv
VYzcxH7rdhUW9gqCaCOIaXP1Ho7Ewx0nNzqUbgtb79L9SF8+reuJdnsCNH1MqJUA
Y3sCuuW4EY8D54r46K36D5nyIgpaAn+n8oAhv1XTPyWuG5plMOSWnKUh4fN2ti+5
8PRBxz8liu2hs/z8PlM2i47He+JGvT2NPrhqrb13AZfijAjqh3+4MuMqQ6koDtq1
AJ5z/NlvYQQMfWWNn+GS952N4Eko+z0ngqXewTM47tmXO7XMPJzcBb9VZoCejlVI
cSW9yo7QLmaKjct19NvgP6nxCU3MmsbZmL5Zc+JEgyBFRO3PMZCcbeQdFJ2FJNZ6
3SnqI7+WZFoJt5ify4bpx7nf/oiWcPrIu/ymwLYGkHwsHrO07xNSggKDHWSi0MZS
wQ8cKKGuAM21bcF7DsrQK8+y+pOgborQJbIi9QfsqgqgxtJtHcrBbF4tENMelvts
JBybhg1SYzgnmqgsNbN9Lxl5ULOvfIp3GpeRy22J4zUXvM6rSxVO9/3sBEzyg6FK
7pNAGLTJc0m+BaqDb4XXLt3oe9/Ss8u3Idk6/h2sIyC46ZV85pYrfGpTbFZnNry1
aipdswyGQY0DxNr5F0Eeb4J8KNUGVxwVaTujBjfssUhmuB5822WZEhLrRlCtK+iK
so6w8i4WNePmqQ6yLskUM5mXje6SjTARcrw+BkUA8VkvGRWsWgA7KyVa/Nw0iObH
5gVcP5EnG9/pWsnKgg4f3Kk2rZD35kv8cwaqItNwHlvmYA47zrdc8xRJJ+0IfK/5
+UkiukOQpOsXpFLjpQ68ZRo5MN8O6835j4FlmkWsJC0Pvul8cxILKkwdsIXjkklL
/JMwiZ1FO/XmX3LZhaiPSMHPmYRkMVQMDrvmwp62an0Cdp4L5rzb26+00QMMJp9z
iVWyhDbFskl15/2uFn2m3wjlSeaHpYHSOXUDzCogaFrp9+ECYrwI7dWqow1WCXdS
Kol/UF4GQOyp+t2rPEtWEVc23TcfsVVXCYGCSOc7MTRkwJ1l3mTkFHf7tCcCVtth
xNfaXnJtK9LgKPwFAsp3ixzj/jiOhL08SiTuhNh11K52Al0YxDBelOTkyWx2r2x4
XjCXCvnq/6w5b1KYtMICFyI5e80PBWJnhnFlkIN55ToZ2ARmpjExdbK7aVM+JTe7
BWQAndxQ2kolDFLWT9P3Nyr5T5hhqqEb+K8mYdWpS7SieDXxcMvhwE4UHzEovb2g
XtHtzQouOw6EzTT50nQRAbtXaDRY2dPeTsZL/idinW8CgKnDkWWdbTWQICIy3sl3
V4LMy/BmXIacXubqXQjxrNwhd77fZKtzFtBLI8QRoBRybhWazjiGZylj2zcM9rBO
OwS6urt1y+2MaZB/KZ9xIZyjVAr+Y8+sCJJn7bf34Wupy5TJ6Hg5Jtq99GECqJ1t
HyEQjE9i0egdehegW1mxKHTA+KHKXVpUjRfGb97EaPzVN8uI6Y+zG7NJuaX1EYpK
I7SLOx0SyXA+eosbtGWsglTCjwMCi1osNipluss85NVYexfzdnOQBpEHTCzN6wLF
eq3ph4HPeSU+ka79nYoaWrgZEHmRMs3gqpnPVT0nlYXLlJviXlE58z6YVYPn+z/m
NJWQYK7xoIjlYJo1ziCYlnimy4uKRa0JU0GZimoPjei/QXG36TUykjWal7e6O2Zg
Y5q67IXkIkUs7QB3yxDzqfUJmHvSDmufvND/AQ6tCeXZNbY1MxdDnYlT7sjUi3FF
umj+ryOBN+s789+tmkV8dRAcV71qGFSNFLm2z3paJtPevhGQjAwG59erwHvX8ozI
haDsMf88BckaP4r8JL8AcySVuczzWSBrAHNlRgaINGlBq2D1t32M2pcSHXh+a6MP
ZKsJzwVa3mO7VDo2D4NPtJH5pF+kL5+0fAJ9jIEnuD4zjze/5XKOYW220VlBiKRG
WIW2CdBrWH7SSsEgsnjaWfdz8du27T+IC2W9+IqAkdBPmQeHNH0M+2NrUM4HudKn
mMxOUTv2eYYUAdXvUqwyZxq9IycQFOeerNwrN9oHd7L6X7YHBVkEGlqREUKZ8NXR
vyG1MyVIZpkaESk1YLIr+7eixAPGNMNrDC5yJwzAU3Vg8yxL6AhYeR7mk3yl56VD
CbOFzkmQakF6bn5kxz3M55HthrL7OfgTmKvdUCaDvRxENhwOF0djwuYNmNJuK1+s
DYEQ7k7u4fYUKglz1csCGcRwG9rTPXQp7JFecmSDRlc55/Mw1nyQzKSVStECVJb0
vlJs4Nd8ZHQMq6NKccheJFyTcg1IUDj+F41Voj+6zYQrZJ/Q7QFd3ULdVAcmCLiQ
whN/W33CcNhhCTjdBTXATqI7wBMQDDqMLNck9i1ziUr3ud6s+CdXg1R8cnEeaPFg
pZB1z9eFelIZ/8DXB3oG5ycEImgXveyS8GYnX+PoyITCxrEnqBvnzx12zkX+r5Pq
9ab2np4KhU6fdEvwKepuPz2EbSgVIzgNGFg+8Tef8Xzgkzexiiun24DpHCTzTEyc
UtqHSw/ke2ABhWD77YbeIEoet8nydo3mkRniwV/l3iRSCc3RGTMmZIzZF56rHG48
JIfg6u1QqLzni6I9VY5STLM5MYhkV0cuFeRiAS3/7msK/yTWCKB+LJ6PetzS7JG8
yG4N3Dud6JKawMdUOzAePukorqlJGFZ44y+WQ79TKE+uj3UVMM7hcDU9CVquu50S
LCVzFbFDakr1hgaz3Q/YDMJXBSzmTszelBnIPqD75ZSl9cPz+JX8xjtrd5vRq8V4
/cdcZ9xL1Mcs4NyEIUbiehO9revccHDRiqWna0vdBDq0G4OQSH9Ode0rCtOc2Mmw
68J7dRsiXQHwK0bRpGGv7+/PSMvEXSjTHdUHg9+XZvANXsAcfc2qjnRlYxM5TBEY
RK8w1ia+1PESizuizg0/phZMH2pplqe8kRDbYxiVqhZpNmVAjqRq/JAZabsYTvW/
uvFt2w9HZElyZXHKVi23lkYBGEWnNVJIaTaO2Ms9xa+PQkw1pBrJD0M30EQfLJwc
8YwCufTVTCBP17tTJsz93ORQBYD76j/2/hITRK4+Mrw6yWLMd1ByNQXzhjERxoTD
O/8ZEF7gJol+2Z8Lr3qVTtL48ekndoHqZUS0Yn0uR+dOkGdHHk9ieltahd0wWnd2
iu+qc2ZGMmSuPVSYo69AqQ6xEa/nVouA+/3NDTfiLNPvHqX3RCh7Sg+cr0mTc0sy
Xcv5g7Pr8gsDJZVKcpbuZgyx2e8WwRJuUs944O/SeXhekay2fr+sfnfQ7l55pwVk
f+l1nbrPNTY4zLblVStAnslfxbU45cT/6ailKsfxnqcMHC9BsK9vqHMgZBPEUHdT
dYyc5z4uGDMBSmW6P5a7RIyLWkUYuH3l2c1MQifssUuuMJuX9Sz6F74Tpm1ddxok
h2mq0ylTmLWWEbP8QG39AzZGQWSzwwkb1jwyntd/WE+7N7lf2uMX/gg2YwPraASr
g8D/pqlcO5FBukjTxOd13f9WROCn2VJOS3a2yBj2AIJCedhdFyxfN/0F3bXmKCfu
HYv8XUfjmkmHbg63gckvtwC/V4VtTkk0u6VAXlfgwWp5NGmGTPLw8xgkCTAl3ev7
14E9oOowuLE9EO3hNfrWFgzULWtL2497l8n8DwQDhVpGM6mpG+mcCFJHtWn5xBPz
XUB66oA4WpIo0Qg8V7zdeWBBYLOz8wz3rdGQ1ixPN5WMeCyPcQlhc2JK9RyoeZMz
XJ+z9a5UUtXiVKGhHySNN4jnc4WZnzfWmtaJp7tnJJZGe+gLzhWfFvKWZZsKXojC
2JK1ALnFt7tSsJf9hqtFqxjXTtMBsCNTeeIzt7oTzENzIU3aVa3k4z2GI2F4RPbD
PZRCu35qxCGtyVzrY0PnyFCSmVqarNmw70c6f5Rlgewxodj/L9JXaZApfwULBHKD
p99ttQ1bSkuRW/6jwdvRX9oBOr15OFNWNCZd1oYe8posOccQpT+8OUq3ATrvb2EW
yaqW2TZK4bz5S3yZlJ2NA0tDVOvsHYSz8TzYnrUpXST9h/6M+7cNw4v6MzgYgpDW
uK1WIgkhgIuLEM6yke42jOTo9APuN2TihlHLzsxURpEKbDkZBOgp/jxEUSWT0VtA
Zr9QftI5znwXp9wY7R0uAYwVpBIlb5IMgMaJdrtj7eio+RcK0C+6HRHGBbwdKjUc
atsfdk8ZwJxGlkUbwpBLfcwx76VMHai1B2Le2sDdbrO7px6BK4HqJLKABe0Q0DI8
IjyCX1CWR8+GBEN96nsXnNQVRA62x0N+gAxB3G3HPM9pxzqI7/dQob9HV4P5hvLq
GQ5A4TnyGUq3/yXsOO5STQyEEVW+UUVxZVInLBXnyDJLTGicDOrWmG6nYburAFox
SUhH41pdPy5nhAGTY/QfJOymLsHYCGP2jwb/xJpW5yePElzkPgrroheLT2W7io2j
PY1E10uQvLG7o1Vz0pTkBlHxgcbj4WPBVQQ8JeB5kHzHw61vKkNuoAFxA/N8WZ6Q
YZr6r+7574PXHZYGAU131tFDqhW5HMClb5viRraHNvYPRf4ENlFt+Y9ZtgIgOiv0
Q3CxJ+KWoO0zzYZ7jMOAhmB4+jCGQ1N/tX63/cFaAIxsELlb/NmeMuCTx+7Iz3S+
6TGsrL2W1V0r7nDQyYYhVLXc649TMlbMFHDPqWRaswr05c75ay3IpX8Lra53gAmK
S4YwRHIe0ORnPvO4EcnhOI4CSWIdRTvgGPROx02S0XhPt3HmboMR8vI6JsTgEjHa
rj9XZer1cWafIlyJox/RtEIaegrtAmhPG1GJPBl4JR4eFDr9LKAqUC1xustYspwC
bfbROY64hfs5NkUlsaQ0fWArBVO0loNzPLu1TR2rB8KGGpbTJCgyy3VecVcZKnEa
qgjaJN1zvf6HflvGsmaUWrsw5KVUIEqjbMr52ecqPVp/7FJoqAYWedUSWVp6wqst
KSJcU7h5rgSnDuDXVl2ODafmWUS+zdLarlG4qK83JeqiEtegSqpKTVmxnnUFLkC1
1eU20c76Zj4g7u1XKwNYcDG+omZeMeASFf51WGt9vXVWohRtVl0GQVNhZ2D2vnHX
mI3u+L5M5CTcZP4xpc4a7DyTf6DtvefYZVJ65QYih6TzUg65a6imjlUpUwSij+mP
sHKq8+GttOPfFLVzzTcx0yQBiOSe+12lOGDOu6NY8RMULlugmjBucor4rPCWheZ0
dsmgyn4pGP4f4JTu/Rk/DTozAceABH5hXgRZD+56Ssj7NpvzxVjAn7aaXpnJ5FIW
6kRBWuO2UXt7Rz4i+wL+DXokw79DWfsYgvG70eySnEULg5LdFm2wVxiXCjhea6pX
Ht0uU+55hP3lZlBZnSwrDuP2c70KPyPGncGZqlmRCxboc1GdhtfMIX0856wNeBua
9inp2a9Pu8lJJqJRBg7QmPwwMIVVJFNsCdWj1bfwTDw3bPFog1gcywCrAQ5491b4
y67TEhnYmxJuaAqiNEavPHtCF2gGt++yxfr0AFwLosBFlMAVdLnXbNMkPPpQVUOE
/IbSPzsQhWQnhQa/CQ1Yxdq7nrDUiGu88ydfvUgdpzneOh168oYLovJn3DPSLrUz
cT6ecq9crahYXg3DTLvNByW/z8prY9MqCB0Hbg1Xb0HahWXRjgq3Z0ZWVOb/Zhak
FuI9iJpl1LaGTQu9QsfLHUm4L1EB0g86zrSJFXXopfqGgL6pNvpv2kcXZESuKhzf
5Nqe4B5f/gLV5/gxCtZt9Ped4W6WbxgQrHGVK66wfh5aQZTvkyuCmPYX1cHVopE8
TbKt/n3kTkIUbMQVq0RBJZ6yj83QxmJ/Dv9jHOinONipgACI0fW2NkOuP3sP2eqA
/JsCrnWHx2Yd284BLpCJaLmZyMv4jOuDYd90ph813v3HvO1hBtgX+ImcOC0wVacp
6Ouo0OXxU7nN5yPNsqER1j1zOMad+yYc/WLcgPVp8RDMKVH/eA9LU8pkPZSl86y3
nJB5Uu6VUs4VSs3cqmUqFQQScMxxHj9XYnjnhjoiQ/+6OhYTMlJr9fI4UPoWQL6m
ZTY4ewKzy4QdAUo4uok0JeUH4FJnFor1s9N4rDRPWAW58aaIeXQ1bJ633iBxXQzW
EVKLiu7s0cEYcb3ch8ygRIEGeAFLzDegP2SfPPaJScwG07a4z023SixmFoQT85mL
bmcwadgoZECYMp2MTpGMqLgBJIi9yx9aVTE6AIMJoTrMxrZUz4+u03Jd7pogdDX1
DmJyDIMtFC6JonUhmnFwcnrTsuxLE9AA7b7bUVrUfPxW6JIkmangO/yglZW3tbZW
ZIo8kS8DP9SvO28ZhTJJoNS2BWkY2hltZKGTHlRu2Lwsx33qZZIJrMPRoRKt6rh/
QBBjP6zOE83h4q5q/8DIqNvtO9vJJhupfY8VjnBThuwOV8choqwxHJaM/1fMkoQu
hzF42bpsw+nW1J2qZG2CUNwPO7KhdE3bSBVrl86h7KwkmT8uitCpG967TaMW2vEs
RiZAODf8G7N+GPBFXZTuMoxm7yE/Vg+LTAN/O7NJE0/YcFB82OMN1NUsoB0lsDeG
BinC77mDYWHRUsC+4vPl49c/GvD3HqxSaopZyzhZPqA/K1V/T5iy141ao5hkmSbU
N/Rbh+16Basp/s24lrnWNxYeP6JGfaFnzsGBAMK/150MccjNmZTmuO6IHSs6aSpv
xwt6CL6sNyLjF6Kmg58+sj8OOXGN8RvfwjYKllE34Ich3fh7C2Rlo9JjW0qGlao1
ZvMf9XGuQ+oNrRE6NiqUQN5FWQJZvhcFrJ133cYhV0w0cicuV6o/Qhw8JRl+ED1e
wmdtCm5N7PlbMH5huu25GfEO4uUUesrl9yGoo79VObO5kkVVV8FT4RX6z2FEPZfW
5pTCaDk59eTOizVRW6Oj/c0KcIZljZVlT03GNeiigiIBLnK+nlphSfvpVsKm8DRH
0I4aaW97f5rFm1Tcifc6POxSjIVh7aQkg9Qi1gSn1ifjVzsXTY6kOqZOaQlEtyCs
/+HGeF023TnmOg+skJDKt/NB/seVsTONo3FmZi5b0OgFvboStEpTZxEWxenPVW40
vQyflazW9Od+uq+BxZ0CNvZLzRygk8JF2DM8Rjq7ePBQJxzUp/aRI2Rq9fObTziv
92hyzrd+wkDEj7/KFlRsqa3D1uO8GKLhkc6Cmwrf/6FmiWFBmR6/UIPD6BJsX3R+
jzczvQSNLugIUIbHp5oowyPCt8kx4/zXDpE/6MU1W+pUlsVzQ7mdJkUGba0xOGiY
RmZvdJRkRIoQEGfPmB2h8SZu84ONcetKXCJKFw14DTNxN4zKg5MP77NlRxOctvl2
WMwGUATOvo/U/+tDuHUNWPOcEj0otfO1gpKhkShSkjuBzwODbB7L2Hz+1xt/Aonh
x5lCzllRRW8aSaOCJcDCXIqvhHgX+2pgD4Z6GcdM7n7QoNN9DXw/y7wOnyGsXvOJ
gSQsoWmewjAxmLVhTYlkMcdRJSQA90sLS/saD2mnF4neCXK2HLtzLyyfd/yvrMDm
OJuCfxWQ+tVeFU8iBF582OayVS2YFnuNZSTQwaBpa+zF9/6d7UCmnWmKo0arCLNZ
gmLUGz3GL0SAByrc7jOYpQMfitnx0ufG3X6XlW1F269qobDTZiuXbSsKR5Nk2nUT
Q5rBFTwcwOOJ4nSP5EdM7ky30XCj7ugPFKKmHNSQBIYNs8l1mWot8RQrHT6Sb27Q
8dvhSirt9FtoT26FgdkfZfeewFAcjokSpWp671UtCSinUeFLMM7aG4yMyUwkLYGM
BGU9nKWlRnUr6l3tZ3D6qUgCPdBulXydc9Ju/kDvx72W778SiWVAg+1+3l/0PxwF
UJkrd/EETKnhwjbzwcCW2OGspzL7Z+S1Ti1INHjMxCeB0bLgBCMIfK5EBCn/sQi8
onkxbPn6PAlBFoRzaP/nq7FMhD2YO9AZ/ZKAH6l42NP5zZdHNZ3cvOzjib26AecF
l9Nm604NP1g8fXfXQH/MWiKaJELWI4dYgYcAUomsZrb4g4XY7E0hcE6EIWn290Wr
d3gbxxAAUDkyx2nLW3h67kjpxz2z26dUxANrgZA5JAtZCkMzZoYJgfkjhAOgK8OZ
UrYxAP9JsgWb4z0H8J1XpC860A2XbFSPUbPWXpO/u7hIfsN+FWp3k049JTWIwmoe
HwQ3k6eibk9zpCG3UDOJNFJxP1i76Co8errAd1l7IcaGv8+D/tAgX4G4gS/zFAqI
EHk6ZmwTndkVhi3bq4I1aDnNp+AA0d56rznejDeGdsLlKBco0D/uEweJMwbZaLrP
Rt4UnZoweWU7Fgn3nsjMBorZy/L4O+uWkJ7IRkk1yqd+JLkKOcW7nknTxY3n0x7k
SP8MfBEsYV5Z4+v7g8izgP4kSIkqUiC62Ri+UaMTwDg0MaD/etRihlLDIZHdq3/J
pSSws+WMTbMaxKvEUUv4cSooqjHHL8w/j50nL26WqOWT0GHp3ECOJFnetesDgXI7
Oxooo2hfsZ1X1+4N6KTfmLu3DPx+JWiGRGBv2t5Chyd8ZMIK/gJwb3KIAIytPzTi
9ct3pstw16WKivF7xagVtDwhHmHT8vdKvwTTqA8OMnpLz/a1X2eHE7qJfgRt+gfv
RmeQvYo1i69qc6jTvcNWVKWFahHr/xGsTJUxBeUNGcavD+PmAivKfI2r/22hVnmM
ZCL6Xx6ZjT6EoEeMQ9GsqSOyZR5quuKQLeYRLN0Y3ZmNZFHE2wqSQaTNB/deDWlq
+WKYbwAn1DVTRV2SxEvXgG8kfZKWAPoX+Ibtg7qZ6L76TK0x5i5BwIMCZwNutkJi
Bwpa7DOkIYFSJz6TO6Vrogx5SWqRRkbL6roftwgweg14fpouuSym6hIU7SCJ2iBO
MpNVceNn7+U7an07w5NLMhuzvBPM5u6WOkv7bnUSnE0JUfv67v5HaUeAXr8noNuy
bRa8kHAeE01sgG9xJVABGFL/ybmYP0/WrTdDxKBzRp4nLqRYiKNcfh2LyYjHo5Z5
ZdXvnfFLt1wJIOGu7KNq+wX/nfQZAI7Mn4ZEcfZ9e+I5enTQ6f2mDVgDP0r4asyn
SwlM8e7GGXczFM6f0Dcuq0mCI6iISJk3VKBBbA0jLYSTQ/GQeDl+Vtq6W7XKZJiF
TLo/y1bUEozaGGwfkuMO16+fbWl87mwfiGJbjFvANEmsirVQC1O2ZdBLTjRHSheG
j+4M8XO7vrtS6ef5SmB7CemvhwNkI1iSxH42Qqym+m3bzUUDJbPDNj1ZRwfm+4EO
Y+XS3SpP5cDoBLyREOrmjjsk4kh78eaVkfsrfcH2O6cEAYFXM2e4bqW+LJPqa9Ez
vSqhd6Aa0p/FVDlBMhA9kE5oIYOhoJ1e/79lnzk+2FWthHb9Kxy9H/LjHvIFZ3i1
pi2a4KRRjpr9WfoVNYIpu0DVM3lvRNQBCUQ2Cmo1LaBafVX/OJnpt9QKJkbnQ2mh
zUP1EZfrzXN6CNikFyd4+VSnP0YCq3UNQ30bIEV48e1iBGjiHRFn9SGrzKN3jRo7
x6CsEROvOgnttp6PT1vj06virhQ65Is4X9Yk06n/2gxjkgKhdl8oIT4ts6peg0xU
4Fcs3MTaB1KMVd6RK/tDWW7ZGVWDBrdEA6x8bCM+5Hq0GwSQY+QzF+k9C43nYHI/
pM35//LbJ+t/gDoan6TVbfAC6LgUlwQYvm2zlM84VDy7PRPRaO/CbVgKh3gBlO85
uTTB3ZYTMmRpK/QMw1d4v8lV/LsIixWz+TUrMU19NiwTMUBDaXSiYFXdKaOj556j
dHxbOXJwTI2vipDeVb3+xDFMl5BGzNvLRLEi9k4TCMXR0+tdpa+vPwiyEnQPmIBP
51bIglSnKMPB23a/GgNYfH1MRKi2XFnDF5wP3ZGq9yj8uYm4mTMBU2UeXfoStWrg
1p/GIaZbl8NjOpNhPqWQQMdjMHMl9m36RebVjIvVqLkvXdkPMyUw95pfndPxHehy
kAaY6D+mZqYfVfoTwEy0D4ux5BonzA+RqZ7CxV7vcSiY87BmM4PxGR1Q0WRSkPiW
QFM0qtqWzjnzOVyd9G++woOeo5EjyKTGfU5eOvC3duyie3HNjFWyA/dmK6Yr8pJF
te1v2bHELzR8Pczk572eXu2YdSTFXHhD2C4WbyDJsFwAOR4h7i+NluEW1MdlDrE8
ORKrGKI/u3/KzfyGPGzq6XVQiuUfiu4cazTYoA8Uoq9ZRsuW+eEnt8gnC6u1myhL
NUW7C8untPzksAC4Ff6+bL72zY5Ljwy3+kHdmaX+lGBHtlC8hlh8Jmi9kqluaiFx
Wi0te0dPk1wO184PyBBQTd1ZyN2lCgZopO1rJOuH35IVT/zDL1T8Tm0Sqmm9OfIK
IMpBy/jiTrci7nDlXscdknl87MPaAvkePpSNNTYh1tZeCYAAKqO/dEPcGt2tjoiv
v6MZrSXMGnHkSQ681PiA0Beg1B3FCPmsivchCJ/46X6PBC0dmyYj8iSYNBgasL2c
EzpEovt2gysvfvOO1jRK5SI7vu6vMV56c1anLRQMqh29wKl3hS5diQFLOUnHNB3/
SLtOPVmJ+mjCUhQ2KrtRkPzzQ0+cG763+Lvn0XvuD9Aq/2bJW9M7Fp/7BOTQNQwG
5X+/LZ2/MVQ9z0aUSqppwxPP3sWwzWAajIztPHexeiac2zJF1eGwf4kCHBGFbH6A
3fqnKNXWstlnibhT9AmmN/uKPv+qylbXBV6p+IlvnGNEzXxzmmrGHdnff4q33BCw
EhbvtwXRilb1Qu/x83ctbpohPgAOBCcfDvtHJ5IhBqSw5LKFSpJSXUl8Ui6VbaOM
AilHmpwVFcjmFHrcox64u+iTcyapXc5gAyMJkFRvBfj0zYIj6vn206XUqNky9caN
ZmHm4/23mTJb15a1SpYhHYDr9rLMY6baUOfHPFM2ZcS02cWEsWP5K3VHE09RQmgl
NHAuEcJyUgq/trbv5ATN+wvqpEpYqwpmGvt65In5L+8+MFuTiNg6BlbBPUsyML9N
PXUqj7FiT6M6c7Hp7TKhMzgJ7ZqT1wTFC13+1OoY7UtujMpKWDQWCu6iaJ5nXXbw
etWsiu6OYEb+LWzBo3VgInDBUAruOJgdLS3vyhE9fMrTT9rPIFI9p7cjH4l/lzFR
jLGMy5Zx+apB4iWU/vKglr6RovXDMnhh7uT1Ci3PquoAd2JkDscnhOApUUieGuwA
t4vJTRbkYUmqsE0AF6krnwlKYuSIeA0sUd2T3XMogA7LgFt/J9vpt+uQMdFEe5/n
8UEBARICwSSgAbJcOl0Fi9iBHNz4c49Tz5MF5Wh+IAQWXfJM+Vla5/9QhSaKfb48
4In+NvaSPNynFjdhDEsiX2wT8cLWvXUSl1tr/8G9kUx4pHEGs91zUCXMNY9Fm1K3
ZIZCEQJe9fMaoan+92QuWAWUZa0fNfOMhi2aY4gGPIMZFrhntmBj7Z+jvPmxu6EU
NPTPkgLHn1Lz/syRQEEtjmSG0bK5RdsjX7PpbbK14Ylkwp77V3UBp9v0/Fpcazz/
oKyRJRKYnplUMxd1zdPaBJiQ/HIcxSAqAivsXx5Vas0okEyTjRhYZUMhgvDXR9+7
cUck5juN16rfJjB7WispdgUCOnPoSWRC8UTV418N5ekW6fWWnP4r93ZnnLruevFK
Mlro9gTTejoT0n+bs9L0Szf0HoLknCjUSfxI7xylLXfkTWesEnHbEMixgJlYV5ub
YMGXRnP0gDbk/bU3tedPcWEUHhCuMaNiBKSqKe8mXd0OfhvbT2KGBaC/I0HqDZ2b
pukuQ7LGK92igKxP5nsIJK+fJ8ONYx+Qe5WtHe2PrL1vkH6y25VNAQSgRIwiUxxm
quQjnv7k9WZgji7Maxq0D8oWZzcO2+tWa8nSpxowGUL5FYHiDob5ilSE/OEPjEbY
t/iJVSYCccIXahf/axmLkiZLZ2PgWysrOBVOQE9z/JU6xr3EUZdo00JPNl8Y3lqT
qMrlO3k64GgfoGQEGoKPrlc3iw4h5nfiiosQ/LHPAdcaWkUfZCrS/CopKy16ORKB
spqVfimISd3aPxGKMGFx+AxXH1LzIJXP/FYhwNWAquurhSb6cZAcWaN8zevaQwj6
LAC06EXLri6HfRxJNhlLJFjbtxegyfBhiCu3IeYxY6hy+BRzYL4oA//W2L8Uz7bC
dY8lbCr19y3BaHC+NCyi/Go8BHSJpSRtWVNJcRrb7SUj56jU5hfW6vcUOcdppfBG
ujPG0ZiIHeqKPsLFqlpidCMGA8AWzs1VTG5bVLFALtynELcRtiH6VK50DYYficd1
MfouQpsB+w22vLTepUaj+OtI4nYQxvD5Ioj3N+RkKZAVaDPSFyuFdad1Kb9V9qIe
+eiqmtzIKb5648BU66Uh77mQRK88F5znkt9LP3GGYM+n8inqq+pBvHT8XNJY4Pi0
xUj317UpFoxSJyWS+yloowccqVxMta69hJJ5j+ZPiZRARxa3WAt0wt+raiHUycEI
yFycY0bbuhhHaYbFGrf8ZNczILJqrgGRdC3O6mHNIR5C3mcE0lRY/MxIU7hHNXZW
Vg6kpMVuBRpMj/ZZS3KKkc6uuNNPMWqVcf3aP8ecq7lkvvtepeCac/rZFtbe/evZ
WT1BUYlMn392GYdgWaQmhvHPgggHsUoQayQmsi9ndlsMfqgGcTz9wuF48tNWyi+B
v/7LaE6nhAAGIgF2/Wj1xlqWKIPZ5Fy7wO+FBa4jJQskjTuvfaSFcwvI8stxjNRP
RgY2d813PLLyPY7z/2hOJAat9sBhr36fmRQEsAh9XbvXM9wmECZC0c4p0p/wO6LW
uenefsEmbTRBauKd76/S0/zzvy8/FhxqarluiLFBB2g5Zz4I7Pi9JYFzhT0zuxRQ
YBseEdgCTovLZmYVNYdMYZ+vGd+O9fX6MUTAZbKV+55kFAD3H0hAsYy8phP5wewr
7NI/CgYUisVbbWzjy7w73pQmJ+d+6GGpYQNWbKS2ds2h++9uCkCRsV7l2YKi2bjQ
JYnafsu6qyu8ilvTuAWE5ZEeL5C4+r+VFwnL+gFWZm/2nq3uTK2hOC0FzFg+XMhH
IGQcN4yBa2I8c+yOFtC23u19Do+8f9FnssYTAVJQFC6tHaUsgFxJ9Lmwtei0Gi/E
X0d62gjgIhFu/fc91jtnam69qWgQqMKq3eYxFUxY6JKB0/2Swea3z+ENgtrdfdK3
Xf/MtYYOc1z3UEiks3oVatnlw71nxmw8bCN1DqKReRTcozevv21wQVYo9rx5M9yO
h5DNNA+lihCbpkCwgq4YZ458haubYlIcV7BugiTt7pp0cxm0U8f6SDgvfO2shoE9
i2+yosigwWtvBG8Wbyp7LPuMQ42r8js1HWfestSETMP5q7Qmz4B0An5W0DAsNm5M
pm0/NT9mf9jffHRUqCY7zbMzYmmwOCxJZRevOA/m/xZjkSVivaQ5FaROsVQVn7Vd
shoD5R9Y1TzKXFDdljwSTaVizCHivtsQka8BdI3ZZ9QFUnz7TXfYfSL56QFAB5+y
TsvVs/EDPBGA47mw4wvh9zaR4hTMF8xLhDuq/3Iw7mKDKMvFP84wPoVKOIXY6XdW
0jgcx8pKrB4TzOZk3kF+9nRdTAlu4z27Or3QK4o/peDt6CGoNJpSgnjfWkvdHXON
UIF8+9heKAxCtIFLOa1t0pP0drfmz4UCbfvmWcOu/jYK/OHa6vZznkt2tOPAJZTS
h70DGAXkbSSlRJG1pObINJXr63m95tJMmjmZdaTLZwtKW7zdYE5VGHhPJI75z208
gZjRzTeWNKhRh3CmS1YKVbbXCiiWKR1hDdN9SYDdzgrScTIwDFt7TNeJAuGdliCS
jzgTPI0sL9JdlKj8eEpNpuytRLMm9auh5KDJWCGXOdBVSCydPX+VsJ7xkZKd3LPT
tO+EnJZaSIzbhsGSGRPcx/ac55/+kb3FfEOPEc2g4cR4wFKWA84efsmk30d/sqRi
fLpMZgKvDoO9FQdKeNgPTop66n4HIG3CoJ/9FDDAoUf52C8Nr0F5qs7+SLxVe5Fa
k6YeK/GP6v9utxj6YNytbuWYZc+IIfPDvhDHwP7tDyicS/6XsBx86z49wLqBc4WT
OLcNO9uqnBMQ1oLsL/EmX2rTN/QQ3F7YKkfzfklFIughWe4DLEyA3s+uYM5KoGHb
pBrKj2qk6og5SnABm22n03AyzaU26W9gOxHuFbZoViJd7q//rUxM2caNmKKcHZPT
i9+8eYaeXVoZvSANjikxnq/RRMke9mUKsO8BwF5IPhXtopRQ2UnaUgeN0BWpg4wn
p/SnyvvMExBnMYhTC7zWxS9JPnKwb+tA7fGWADZLjR4TPXn6iGGUj8MsZ6BYRuSE
VpHXa3dflnEIa3LZLLqvCgKPdYlOxTPY1C+3f87WtjGJogylVyCDWrKAlL+1mcbL
JgVpsCW5W8/V382zqhl0HNLQw2DXXf4GOiUrlclfj0YdkW+I/YyKABGVUCiMSsYV
6Vootpnaq2Rdc/abVhB3d9HhM3gTrtsorWMDWOfho00oMhJqYTbINKUT9HSi1qj/
wZJWyTHaFnJfqJ4NFGjFbLUk3lez2VfVjEnou0HRhtsQpdlLaPgis9NUACYMrH8M
mu3kyka8f4K5xTdn+tNpmcahkxMq5+y4Ek1Ewn8bChMfgAUus/BUmrxqXWV5qO4g
b/2I63Ql4CAWd8RN9x+ABQjSWiD5Z/Av7qyg+8j8SoTpvRZImk2KivEwup6mcXaX
RVMLTCPu16Asd1Suu36VAdbMiHRLoMhqE2iQKJ1hUPhynbLhFrKBV5yzC66x7KwS
CV6saZC0BIgZRbEYMD9fIFXfnnXq2cKYqPSkrOmCMYbyLnSSPSt+Ay7scCW8cLSo
PGQUmn4rnJVqPhv0N5uGTsvdXSgZkgCqlegd/AKsvJMCY3K088fmSX1WUIuTuIen
BWe7RHekJ0luExN+FbC5FE9TXVmiZmtLf1QQZXWLKWZ3IthqMalvrrJK9MJfbeSK
FHMef2bbbdBnfpQFz13eJDuvmDFbo4lrcP/OurUbm50hFTp8s/M/MKgP4ei8lPO+
F+6YM/LOdotZ/+7uTmLPGNn2QKGupz2t1MpqoXkgaJqEtGKfXtiZt/IEPIOY+cAz
Z809jl8cn7pu2C3aetkFBUpmJI4RCSk2+kOL7Pnhy5+0m3jBnoNqNS/J/Ms+KNLT
mje4fCjku8F++YQLcMNdMqdnlHMuQso+ubs63jqZNmfNoCn5kudx/SEwp0me6J/I
DMMZDHch132ki6eWLu0+Md2teANsWjtSBQYQ88YMifz4kBF3X07hgy3W+aFrSXSE
H974YIU9oGAaNEIrJnftIUl2c4uPCuguw91+XrWToebHSYR+nRRJwhITjdmnSv09
s3juiuhb8fK7zmzQr0jmxBVq5VkDNN4Bgn054xtKqXxm3vfnPNzbZXg/OGIvyfs8
9woCAhRbF84y4D59Od3cQxROcCd0aI3gkpyockBcN4eaM35ljFn6MgtQSf9+12QT
1Nd7prWULasiga9yTgB++bUqMGZLF9tF42N9Thj15sXL4l9LipgBoEJnQ4vmGExr
ZNRjIGrOhclyLrDSGQIU95lMarWJN9I1jMlCi1wByhClak5UmPrZhOo0kefkyzSE
X5VglY3Ud004bCHdr+Ujx7ruGN0cawENLxvK97UEtApNlD7zOAqOLPdyrIZ5VQhl
Qe51gheFfPSoYJtwfaDfP+ht3z+mgE+C5kCPS7TPTHF8QSz36j/yY6jtbB4ObAPC
odlOxtdD6/Hqt1V/+acgOlF8ei8+FpUXpe6Xni8oDODo2asCFXE+XGNQtDvpQZyO
0ZHNdxp9MGNG/D3jUbxtkLRmRXNmcTgcnVXqWXImU1lbc2ALaHmBpJheFSXdEjWT
28ZAAxLtqs/W8sYGgeoBqHH0vTJIcd5HG/7DXthBeVIQAzmP0e15iINGF0eUSWzn
kDbuXvlowzU9TMjB7tmx8SoSiAfQxXkffaZpRsjXspKdIQvXPcxtKdNxNTM1fLcY
ZTXGTA/Bv1/l2Eq0NZ+sWD62EMxkK4h9aaTOVL6jIPtnRvzg2bIRi4IXtOv12TL5
+ibUApcA80Yh9hT00Wq0z22H734GgXq+ZV1xHM8l7U5LEnUQfY9eZ5uqZDoatFEi
O9wqO7hst7jynfAk9xRxtU92AeIILYjOwLVac1gHSqppMNObl7Rn0c+4XeCu8jsu
oBAWyN98wf0QZOcR8oylb9Amx7gzQsBw8cz6zcL7BP9mGGWv/Oy4p9WqyWP9sXL6
YYlyN7A0w10IkqmaI/iSOUhaNSww0Qw9ih4x8p0Nfsz4TeORp3ohMY6sRZopfJyj
pKdb0rziIAAyvKP0YCF7apqmxHZHWOdIfV5dvfFQpu2rpQqn0ziiaGH6/VP521tL
SOTMhXd2WEiuzwUWT67t/KRtrw+Cd/a/0e2DMoXxloN3DFyVIP0Nzl+zyVB6DnzG
ESDSRApgDS2eQluWSfMTr65G9+SPlA6PWbDcxB1H/3tg7hMw8cnUxI139IVU4cFm
FWL5q/oR4EfhqXMUye9m6uxO32br1Ed2qvoyOlRZ904Nqk444ebzQ/n5lFQvUiPd
QxBjyT+90m3XjbO93L81IfzCpwQpCw9bUW4qYXhX06Tn8j2oJlPMFouLXLYxsmHs
yZG9creaLXPBjn7TgzDcU2ldfm+yq6+WPXq9HBWCDBh5pMLkPskFywAN6y16eXa9
eP4T846SrEeKR8WAJtHNe3gmF5sjtcPEoZPiDoGFV5r7ZLqAboCtjokoa4f3sIFM
mkjaSDA33kjLLwNIHoop2CcBWKq17abSxSICVlM8RkVUcNcZy/n2xvG9KsdPB+KO
GTsroXApSTsK1xUMGBsqABFQMX9s0uKYEA6EQZBkbdnL4FKgDgNglYf0SROiIZwW
RjmBCxqbf5K5m7VHdhRGWtEKGNMdv92aObzgDKmJOGdDvn78mlO7tYi39hiig/bB
IOIVUwvDmoBZ9j1IqQNxsxYgZVFxx4BRilr6yLssxY75xFtnN6sZzMg1afB/2Xle
aMmRK25z/6gAmhZ5zU9Xh25vgNer37EdDI1/WZDCsNNek0+u/lrQ2klm982Cw40C
2IEnsv8t8kmzWsZyjxrdQkda5kUcnrE2oIgSNPBlbZaVC8LKQ+kZUbh9iqSQ9AuD
+mWyctqthLrBQ90xzgxPVeGQI9Uj3OFR3MNKpcLG3U0O4FmFLdu51ja8egkhuHE0
b24feEf8u3uLN0tXJn6rdYrdxtMt5MhJZyEaHJlATqd8BUKb0KAhbujFg7QCjf0q
ZnLaabrrfQnq9ls3vuGx6CgYgNJP5qkGgz4+bW37OdXoOvYhjDrAOWRGN9rlpuGj
7MA/YMvvjryQHOltvNxgX2yJ0+Y4y0UlfADP2kPvnanNa6t6hcj7mPKb9AJ9BwPq
MGLWKEI4V+1WeEnRRzu2G2en3Rl4pVpLYf4hVCa+OFQ/x+TDQmZSa48bhhpYerh/
LNPhGRrUu2cNbbD3s1mjTTES3fsLjDvuHRk8HZsSvZ6qvZR1Rv84nyjOtvLTLCdl
I3XkxNsOp9FhVUl0mT3KOT6b57S8+izjAxsaF7A6nWr9JEqnUtVFNJJtfHdOUD4P
UTuVKPshKzW+tSIAv0xRVIVxxzN+i+H0rA2w406F0U3m7/0o61JnkN6rA5ht4YMJ
jwIEJMWCuTgLKuFlAdWGBNUmlba9aPjJrGiMSLqXyQjBWj5GzZamQg5j79zpPGYp
ze6bVQDKLzuf9YCTc5TNQrvegAVZE0DUaiWktn4lmYN2pTuLCo3jNzjuJTAeynKQ
F0ediRPLJTAmEjoRYI1iXR9ZZngfgFqMp6CysPAlZsgBNMLsNnVBd+vxjQ/RPA5H
L0x12abu3fSHSRrJ3/18VjuIPBq/We6c5wTUGP+PFObsySQubueiUJhjlyIKcy9j
0mF21uS12LGngvt+5xMS8Cr5X4sPYJ91V902MlT0LiXUcG20whJKeyEBCIoWFxHv
IOnDJWYUDh/FG4i1pCRmAp8RfOg2YXrGj70xTT/T0DUNiSFHK/TvGyxGHv4OPP3+
3tR92TKfBaJOgZLeNS8MwVjlWfaOgeZnafjRmyFs5ETVamUjnVuhFQlVo1CJta0N
RE+h/TXPSIL3W5uxhBQ9DiZZpye0UpfbPBTdHfhxmnAGpXLmt9O00pFASJMObJbu
fayOvy8VW/Ki/Bw7NqfL3EJDvBt47r0KPWeMp/CcbPcHB+FxHW43Y9EnBN8wQRz5
OSd4pFTebRe8yeXRo5EIwzgU8XwMUcLv7aS6qMUlky0qNbMJNpRw7LsewJBfwvGF
Dl2pcet4GrPzfA1R2/nIAhUobqnOdJHbzG33/4VCXkbs99aSBpwDt4lBh6U+EsLO
264Ef0zWEthv4GPQEUDb7t3noONSikrHNVJ0vqECxUMhQ3Tcp3L+A+KZFW3Ic4WE
aiQd64jPC0vFDzI7T5uy0gUp8zOyxsRqWjcUZ1RURQCFYEvVHMEVX6csPG2IdkNJ
MN4tkui21jY+9voyFhtH4nKBPMCWbCcnBQtHPckhg2ELg/BDmSglPXyUflVG7dg9
coZEuFNMxhZTAqfhC79Q+LaljuvRRZS2R06ord/jWYAJISZuQunNoWKMSd09VASX
SeYqxPNh+jsJk6exHdx3gIR5HI6RCkW8aMB9LewiXK39a+m4djYjo4DYG4Hdiy4k
7Q6faIuplDGFjz/EfcnSPxgR2v4RWbdTI3wSD+XWfJUGoIWjyhE63lS7XhYhlEvU
XsL76ZNDH0JxP7LLoqUKLw674M/I7TpofSsHD5n8V9nficQCwQGHHUPwunVNI+GK
TTlh/AnfN8xDlLElckwmYwXofQFrhLv4SgRW4DJDGKfkjEVTMVk2Oo6gmRQBmNdg
wZLeHpliiEll7rGLV8ww7QLgTxBpwMpG2O71oxXA6khGXOpij7RMeSm7CtHjdUSo
6LzhZUy4Av2vPWzOlhLLrIDS135/+nkiTP3IwGAmGqJzk7HFDYnEEVDOcwAywUmU
PrSEdXVVzE6VHV4jV2fIXzYdHyQ8pNQHqeTVcIQ4LM48r3QODD9xPr2znJTBxNet
s8Hb8CLfDOifYDE+COvGVZSF4JMcep65eaaa9M/Q94/lc0aVvzC1cEqqUwqNsTD3
ORkpjPEs8eGggp8ZU+sQ46Gc8hyqkojuNYpCRctDx/FVlltdnywqUIG8MEeWyMEs
d1XkME4ImW2OmOJMEh2Sul0zj681Qe9C1DxNnss3G7C0jV62/W/HHbWbvrw2gCoz
IbpTnioMIkGB2Kp9L25DQDgDXvTsW/8EW1r8XjXwDp4gIxJr4frQFEfHiWJc709e
Oj4zV8+uyiia8BxTHfgQ1Z5ZUADJhsrnjCsALNai52bNJrpP3m8wpXSBSz7nymmG
cdlmAAWacmfZ9gvFlLPmk+BUAErCXADRQ0Nm/KTfIlhdNTbwnBZxnYmXDD0tPovd
8rLysrYTV4TdxWP9dm2ex2OC/w3FyiDd5mCd6sp2gQ7WuszGdR3Fj8xhk+1xouZ6
HqPNLjF1xR98Y1eIJRpjSA1j4L/rXoNXRnC0qR6Gc68HS6wFLc5ZZRzz/2b+jLNK
7wJiHT1Fmmblp2siSngdDj6oxMz0IBybtWVcPPfqcm+UfjU+QlEv2jwQ/1X8kbIO
AUfm/q3N1BtJFav5uwen0EBFIezjPIN96K+hH60KzO1cr3k3WGiwGUFW9iAuvoPy
8hVM3//5Px+XgaT6AP619fQMoAuIckDCCwgA/Jg4Buiawhij+XCyg9sNR8Hk7AdG
PbQZvFDAFCKUZTGcrdOjgp4cjPVcBbluj/s0J16oGddpL1CTFU0AjIyWVL9cS0MC
yY2MDl4+m86Dtu2q6j766Ljli37mpBamaeesOumFiu6YWHWFGLOlLrtHiocihRCv
dy5T15CMoQCkhQC9JKbL+P/S+V0lzH/7gXTcDlZYlkttNcc+mnninJ5osB6LlTow
PcsAENDUpgvuKLITB3vcvPk78XoXzuQ/eUooaoU/W/6cCFqM2cpnx+xZjaYFdhFq
f7NlkmuPFeYXrrJOP0ssT/WDuvohiUTABGvezgg8gTNk1M47hbMEFoOkxjGoRdAs
k03C5PUoAHNbjiCdbs5i7buyKtIeaXD9z553MRnjqaJPH8GGtj7WtYOSewSZDcrL
ErX44aifMqMaGRTPQwJOBIcIWNA3TOSd+b1NX32UrV/yXebyki09xV/O/cXwEQzm
Lt3/PtqEP0OW++a04OQyeJFCIArLJs7DfAK6TnlSAxNZaY5bIsMVx3xiU3EfmPgE
/8F3zEFguWtCghOlx/LzjW4xLK6jnGo58RXQbWvoSJCyQvn+0ral6rGHV3LTUzGh
GzDGZLRwWQsvu+77kC1ZWCOiQGiVZC5AZikqe/bJnXjkM0FE1JgxDdxZiKs4MyVH
Lyq9sPrt+cU481E8r6nXzihCaTc73GAKJSdN+rLmnrqO+otDXSwcS22EyXbByvnC
+EbN9Ryrj4aU5GMkiVQd0qCqPro7pEFJ8hVBzZvewOg9GIcdEb1MU6KKmna18HPo
MnNyKAR1wIvmpzgQWuGY8Q7kjzkZeabRH94NsqsYVPKX3UnuvGBdYIsUE5l6C6vV
Eg1KZ9W9wawfpWzzUok/VFKtnuBc5SJo5OxiBl/jjW+MfNPeTfW3UtyxKIV5XlEP
GgBEebdu7lHZqdoNiUIZgNo6xFvW4R38c3roDqdDbi1WuVVMCb8wbEDxUtwlRNHA
F8sA0Q0vGkktzzs1NDjNHIr014Yo5clIWUkudnBEnR/la0QGUG9HsIeM/yOCcdCY
o2cWuf73ivaJ5C98Yhr1D5M9pR2k4z2rNzXEAJTvDrxiNGG62PFiRtMNGxRDc9Tm
ME2WHr94CSUIxFcDQYndhZOzkZpXPDEs6zkwjEXpc1QB747ElTnaU9RfIW7dJMuk
orN/ul3r2TvWcZlmO+qxeCjCeDmQDbJNw7L7OdSMpgpLVU/0oSahu8LqKG/06Wyt
FzTUUtBUNL1vpuaIzkFI5g5DDV9pwH2Sp9fxzfMtu6RY1JddBqMv6qXXPwY0c2PY
rkLCcH+9WYBW8RnTg3jY04WMi4Zcj6q0HH6ScEsiVq6+aPscDbcfuIp0Er9/Pyrd
hg0u5VchKTtZ90s6EJdUm/zzEkDFhIuyqBr6EBnujQlWOO/NR8jz/EyBkOqlWtYc
RysYu5Q0OCDWN9bRyFH+XIvhvISkibj9nxKaPDgChcdnwEz9cr08TjcsmRo4TVS+
9OC13ruNF3LM1KdsyQRFsZoSglcMZokrGHs5lfyco19eu2jhPG27r5vMgGg5PWYC
6g2aIYjgzjBwFkaRVdGyU7M8INe4xZmuRunr79I/q4EiQNAmp3mAE33d8yD1BmpP
+NR71lyHPMSH97kMbETc3UuTv8bNC7kw6YJFCLMi7NBEgMKAP+3xY5Nc/2I0vgII
cgX7wBr+9ywxHx+3E/4KLUfWYVI7fyp85k/blS20sdoEkucbHEQPjA3KT1pIRwyz
QC8vzuDeYIHWieUQY9jG/RI7FE16KWJww3czCu2jURPhA6Fys5unLrkudyBsHj6I
aWIElZloZGoyWpYtz5qBGvX/HiRW13c/SLhlbztVHlI7/SD0k+wRJiHP1ZDEHRQX
ScJH2B7gE8hVo1Gxau4E04n1wO+C3eggkzktclTDyZdmNjZHzpPudVcJgOQyNV9O
g0dxFx+URCDR17eZQVkqqt0JOhHMKdMh24eHMUK8Ne980NCz3bGKAFGLKv5IJaoG
7JaR6I0PYYegFZM5a5xfebl18VEPFdeVYj/NmCL3DMEMYfCqlXsqhKxxquekT2cH
FNdSrNgZRj7MRp6QaVV2Q5ZMzuexbnTUO5UD3V3kKwdpjACylEg/jsPZE3XAbYH2
3gp7O7M40qY+5IyZsc7zz2N8P95QWNE2NGmAgnL1CBKc+GFAY/rT0qARRk5kS4Do
vXEgTBtJ1tzifB58/qv9A/9z2DeAqCwNhZXHjc7ejqP5Yj0a/yxDq+z3PobZNh+5
dxSgcXZ8VWAC9P2wg0hKKe7h14Qam76JcUoz/z9ZoxsVYZcCRZmriVHLYQ3pE6m6
0m8grKpaw91acU56UtzStLIRi272Ipiwm48idnm1uHyFrAdqXuifQqv7TkGJz565
Wip7dK7+2PVegfq3UkLOirC7jDuAIJPwZahcKxF6xxEkDQEcbj4g2gvLVk8MZbVT
3ssT4cTQf44ElSt65IGHQkx/W5uLZmBOcVQvOkosueAbXxyWYSEj9x8aoe55SuWt
hwAiufkEqmQAF/pqRyaOXq9lBZpYUb6VzbRaNOMgys3IPsXQQscHs2S1B6J+KaBL
Llx3Uf5USD3+RZgKYEK+TRqbGYQ08lohV4dFR2JfHiwUHlwS5rZJemgz0z3zf2i4
iWR00/z2HsCeuznKs8zW9OxvjDINw3hwKaOXIr2qmU7IK3Ea8AueHOt6vxLFr1xv
6zZ8kqrlvePxJvbTE/BrknadxWSCNcYprOwPmGjh0JM/w2ysZUf5oNFYJ/opXoza
k/cAHxCak7tJRUS7JUm0jTsJXiwmrfProQgJCRLqe1wWAnoiX0h7aW1UTe1ycNsn
q1wbkohR01arynAzAThBrOAdBd0LX/YQYek/+KTCEO5FfsUTXig53tahaXqp0vdd
SxnVRXud53RGi3sJlzmAN7FecCm8RSGPFOUqBFsZ8ANSe/+tEtvXm5MgvvXiH9ri
C+9vzia/XrITRTZB5nYpLt7gemujUq7YpspS/hkllcqV65UEQYCzUMrLRL32z8e3
+LJMhGtm55vN7GSuZkWLIfUyKOYHict4sPDK1q3k+1URfipVtbWhQ5zLa4eDCJh/
1F1SqUq5bwqC+IutCbtDta165vFYHjvvBnu6thhj0SwZgud8XWNQv7Sjkq92WO5V
hYs89xdU3wvaCQDyTorr8FPOMk0GDmGLgsSooTqZgY61awC8wSRcsxeebGAjbL7v
G8tI06AyJ7DGuR5zXfgkai2jWke2mJ6Mp9E5cK/ddVQI0qV+rGF6PIcXG5SJDGXV
NnY/upzEysPEfSSmoLGQS8kd8vOEfTFglXFMnMy3vihZGYOHgD3oLNpH+oue1YMZ
dwd7GX0Sdj6Yl9i15tLZ5LFjlI/Lmb+g8guyRwHKGhTB1c3HOMWfhujVsUIUS0oP
FaoUr5YRkSSxxa+NytAfTL3VMpZFmUh03v9q0UxaY7I3zwyNa7hvF3gAra9Ob9VF
z87ZZbMjazYjoCLgiyPPfgjKSytejJdLf25a8gY0kh3yfpoiW84NEIQq6VZxInSE
V7ErcXmNFoDYveeArcyGhYhDzfhhtpPXiqMQ48bkLkT7RwQayICeMfWCJ6f6mPD0
6E28FjGw2O3tztcPdXdSENiKXNTXwQUJDiL/kf0IPbo/X9GBPmWQeR0Ahf4jfYrs
9kTLSyVGBJomuj+HA+bSqjrfngCjZk+v8oXVfUxpwgHyd3JCQFP6JqOQhumDDZ6U
hhWe+ncXTAFrCkomQCUdXWRKXxDdXnUEmUHMv1Rir78FkwGpgdkJ8+yGZi5pLZQH
P3xRzZgJgH0MFUqNWMExOaVyOaY+eC/fQf2G6Ju5VxSNsrAu5qu/uSuKdvIBdwbm
mgjFJCCzmJg+SoWi1yPne3otenP0NARqDetR0EKQGJHSWD/7Mb4bj9wnuOLVSrdv
bsPdLPgg5nBMxHzCM7xB6sr2KGluk6i3Hgc88+7WPabzfQ8pfTZrTFrVCtQZB+Lc
I1ffw+Y3oWO/OBISNLBDiCUwqVCaD9fxCukPO08Sr/C1w8zfOZKMaKB6f5nqfiDE
tkD0wFLuyl7Y90tKPRobB4+9dweD5AVGfL0NwLMALLcWKwnIFlxZQumzNipRDd0h
QueK/R4RibLSLuS7QY9DhS6/uxOkGtYGKww2oMk4Oh6I4jgaHY3AnesNavmw1zIl
z0VjB8vOuJBBPSyFNREMnbdgYGK9WtzF5KTEm1qiLprDYb9L228e0sY0LWtwlTIA
Cec/JyJeHtIIEoWb/KpHNDltMqHXEIqLw1EwiV5FS+FOiT6hymOsk02va5sdJfzs
H5SePKHgzB/ROm/+jQOZ26M2b7fXT+8hNlXXwbkXqbedqAIsk45pU+j/ESjJnYL4
JQH/3CfdFgMm5L4fyjgrMVMZ1RuWRBXjdbzj7wNayKpaaYWdwDfUjOoE2KNo+xVw
8+/JuLnN9x+QmfKi2neH+As0ZFfuj5jvj0xn04ozqDkdcbnYeGgqdG12ebWRNcWW
dxjRtzeq3Ep2R6rJGF77oqU9Q8je9P5u4psoUwhGEm40n80Qw0S6nwVgwOzCtY8G
RkQodL8JRbz1OM7LtSHBnIqGIP30w2DaalbHIDyW2uJdD3N4VoW0isgMdZB/CFDR
fr2y9qcEvI9Ek6DBehJiieJj/l9KyrX31scjI5h9FluWFqQGjYubVTT8hj61bIyd
jCrz2KcXsqkDtaSRX+5BfHPxOiBgXyNqdxBe2Zmuygv559wRjlCrKZf0vGXjhZJA
ffWRxqshGMpDXwSatQj63SUOSyCS7zB50Y4FOxQx3d6KCWJ6J6dqfTsR2PdBrkVR
rTQIv3ZVUO03J9Y6JnZhVDNHZC/cQOeLLXjsnU00ArOuPruD3j56Kquo457elmfk
qnrEXahuzeLE8OnECkR0iPn3RJHD0hR7Q026E0Aa0w53OLFpLic5KLHSjcDzzCjb
T87SG3be3i63jpwBGveQ879deW1wO7+VXPllyoydZRZTy/nGQq0IL3kllmjD8KIr
XUrpHdSEtBBMniySWpbFyIiGKZYpZ+5s0vBxe41BGEs5+qTu9r6o/pg2kQ5upoNZ
69OtWTzFJ8fd21OYGO/vAcQyFXPVooeGtY/jh8rgUGL4mO057e7mQDTcOpV80AcQ
Qq5qqFT3CBHfVsa+iVf6RjlAnP/O80KE/P2JgQC0t74RnKxAouGUgfyi8r1R/Iq3
K26gTtPnjPMcXciAI7Z0hsmQJonKAgFnelSVDWzixE7DnVZihx7QWZEjgMdO8LYr
uuQCtwQq2tEbK/B+F3pdG+kponDtOs4phGrba0vH3RDUk+AllooG1+ydliN4Z1EY
GoKgPvjmca/xdV+eEOV1cimepMOWYLoFyNgunwhTZtU1Xcd7NYHoOPWsHVro6BZv
+jDYZaunS2hj2WAB/4/UBOGcEHhxdSU6y3/LQfxwd9PjEkUfQuDcXTXD9VKlSdho
jwf5May9AG4U7ivDTD5/mU6mrf576U83qfk9bZz4p798aKI94ytLLpYYWTYhD+p+
MjS5ByaE5egV8PEAgwHXVt2E8rCiMW0tY4vzcIHQ1TpKX5QETArOdcesnGOovbPB
ULUxh/V0smz93bTSVh76e+Xjao1weqR3T1e78M+lE9oVWSpLlhYxDZ2NDygs3uaZ
X0QDo2ty//JQUK7asV/U2xfZiYV6sp1LJv2bFz4JU4gxfNLk3u1ECPd0qz7lNzxL
z5J879tiLMJ5rLCNjXvcMLcpUwmkdtYfMwzmpQSoB5uNnij85WWRzW+rSe1hLtam
Zu1EpqMMkTs51DLq62E5/CaYsTP2otYJKlDYsmfBteFIEXUA3iBRUheaJdTPiXN0
HqYP4jTNj4IWDahSgIG4BxNKISJGJpqeqJVkuwuHKRWoiabwqNWChD0QjsslHRcD
Nj9tn4diDdZHAqkC5hCfwYRgEXZ2QWINDykfQsU4/HnWpMtcrljF6nQ72Tor4Dg4
CigxDh1deL3jtHIHnfLOBWNpwM+wDA3yIptSZste9pQNJd7/U2jU+18bDYWiOstd
NQhZ45n4mViXKe9d7Qxud48VVpnpF/oA4GdMpMKc2KqgFlhAj/COtY3rTwuZu3jx
rq4WXLSVsf8144/3HypLJt0hJ/4J8LeJDfAaTuW2Jo7tPCnxTANaY30CYLA6K5GJ
Ift+ObsgGcyHgHJ/oH33eQghoFDMlEbBaZADyQ9NzwfzvnUbBtnPKIe4V+saXKQi
gvoOhRFQDZ/7msbZYfC+q6rGEZ6LChbpCGqS4BcTiy+0E+mqFKF+4bibvv3/GZs8
7v29nmxFj/Awqb855uRxoogVhG3QZRWhsy7awmiIydWIu0aY+f6dzwC++v5ctrdf
KTZ99tr+dGZOA+QqhjfKXC7RtFHwNCJxezactTJE8FYhR1hBIQh6I3Z7BBcLTiBa
bdKN4jIfsm/1nEVgveNr1rBtLgk8fXHyEHQywIH7n2t1lXvTvkggeP6V9e/nZGw8
gcyujLpGNSWtEG8Pk63fkoTZISsxd5EpsVEGXDFS46dDFrxXZFmX0LMjng9mrg5L
NBHKPBClNiKIIQiPcGpksgSCFNULkrkuZEYAT/jzqTpdd+8oEpSbHcfSY6kQeBpV
92Xte9NTvDQG5uigckvOXHVsTpL7KyFgbv39SXeWscemGtdr4QqvBG9vx/ncbeoW
kxabi8vGHso7ooRH8+rXW7sakL1NveqQVm+7T8VxvBiOhUb85CzvA+FZFQembbBO
yfPYNQe+9XA6kaU0Uiwega0XdtC0JxaGsC3ZalIcL9e8MxCoFCApD0DgebIGKuJb
uOtvGr4+oqIJIXunuizD6NR491NBciRpGOeL39AIGU9P6A/FpUtTDInes2LSm7t2
Eq/MoNwSekqtQB8A7jj/x6Gbt7Ny6SBQ+2WvRZ0IlVtZ81GJtb9D3l56SNxI3tNW
4Xf52Z0Pr6Bj8Ye805U8MQ5MKDnVA+61Z0I9RvbqwMsASZ/l7tFmihEJ4UWMknbA
2RWafdYoJDrSeF+h5guNfXH9ydQ6JKAP5E+ryT1e/kWngUKkPb9UglhGPBATUwbp
kJq2FQOxQI9eI53lpnLyINhu2sCZVeTkXnndtEUtmcAPyREvmI/ibS9BW23R20DC
Nl1eCRUGHgQnE2NENmWRFK2oFP3O38hlf2BsYz8hozgkPOu5OaheK82FI8jCA3PS
eN2Sb1HfT57akG2lroLqh3HPDuW37BREBo4iE/MBmn3UtwWCL/x3qhyxPcUOTUBG
2m5F+QVUs7cHM1YED3S8tBXq67K6qgYG9CEqnEs2gRjZnZb7s2ZdrFCmgcUtk2DX
0fJ+FYjd2eNP3teNY4NagozbQfMAfz4YO9HbWfhks3ynmEhFCbPBOjtGtfbzGEuw
gHM4Ztf5m/yrDsdowr7Ifhjh2P2pbi+mazhO6S13yr58JK8pLii5dNynI0L5Zqo6
dORlem8Fqpqb3FImpSmhZB3qacE3kVQ7Yr1RIhft0YjkiyfpmSczG8VqExJLqgiD
SVUCcvWUHxH0quNONLk1jTRqvpgjSLteroptCkpqEVXQV0ydw7fG/1BbhYZXVkCD
a/k9kzOf+aVYl9TkYyjOIhSbtY9w7DzVKbeA9pzYclBERhfqA1efv8DA+SQC/F8a
UKotNr+6u8wR8YXFgIAzrMtQM88I5nXhzvoaZv/IgNxXHcI0iRVwVtoWxEwJYDoG
+ayGuG0JJB8OI8C1wm3VclpC0P3uyz83JFDPoJLckg2HUL4sQA2MygBYWmbjTNiN
zty23KSmEvetJVSEtPmcAiG1qk/Y+n62IGjA/F3MEMpmnebULlrI2qcz5yMv84CY
HUQ6MHjGBKvKbK80v9+0PZXZ17BlDMFQR7Ozp+4iMpqMGcd8fb0SMTtmXF6KSUwr
cnFHsu6xpuCDqBnZBO1lKUcutmgaW8dIfeKMb83I8AV4NPexM+hYPtrr/yJn5lqh
MJ/7p8+z0eKAayKbKs99JzTUbEx6Yf7Juq3/KupwMoUd+sH3Xh0Bg7ZY7DKtahIM
XvpUy9cU/zUxj7JtJEjvHmpVuHjFIUAAoIThBAnz30coSQpNjJLXAqkvXeJ2ocuA
FEy8L+EteS3CfeMpc13OByixi8AM3sTAjasmzi21QBvAxqwbmJyfyHh1PEOK6RUP
0wkZtXIjUbYfk1BAp3/x0E3SDdf2ORQa9ZmcaKPHfmGTcueKr1rFL5BA34CEZNhb
6hL5Curfen+tw9siwefwICzrd1vWp8LPDVrq/kAeZnruUAbRSl9v/NRtmsBZEBDm
FVj2tZUgE842/QMRdgx2dxT37jerxoNKJOVsJWhhR4aDkVW/tp/qN1dEiJw1TdEt
gqPOP2uWMTiSQx8wdi+vv4H0xWkXvPb1KkRC+WGFCw6qwZt7qZZqFMmZSnrTW91f
5Z2KSFVmv07RlhruBQfmwmukoSRfZx/N7Kw0wxT2DQfJtLxcvMHlUJ4PCDOYGf6h
/Rsl96IcLw9M0Kg66zLPn6o304M3srzTGybVCLFrsrMN/04LqUi0cViyRpgZiYxt
MAK16u0wE0j9dRYoXqNnijEGWdXX32YZ//HgXU46LfuXyYw1HAB0cfzaqyj6FL6u
Tgq4OaB9x/KeknRBhlE8Wc4KJ4xSp6nFXdNZHRlfqs6dV69HeEK+U/Wm4hyMIvYA
i6GdYt5hEJz5KHMHF0TnP1KLONqhcLlvsaUe3BHbJynRvaLwz/nzuCMNT4Y1e4XG
7VBM8tpfVyMve6zesGyHZeu4CBSdvLibnWgbAv1uILXAMirlWXNUVypRH/fCdh34
nctRaQNgzb7gduHqJStiL/EknSe+Lv34oAWlfa/xHHTQrnCd4k9+rufwW7xnDexi
broqZ/AFBYthhe+wgjRDeIJ6a9Bsfs4F/dXDKEqAiOV4pYR47l84MWreWmvQKgl/
noueTMP8p3dKJr1EB1M9FdJFWuhTgQh1R1DAAoVDOvDWUFzy5sGokTuecuuuwcpH
Xz8zSXUw98ZxR51BxxwFJNQeSlStnsvNpEeCTOUi0Ce9paDLc1DB5hpnQdYVzIsv
C4JCCDhu7Ql+3JEibKjypwJ05DQ486FIe6r+BzV/eGUILDrI3QeVB5GYs4GAhmQZ
QkVrf9pvoIQgGs/4dvOM7F2oXPDgM2g5FEozS5KD9LZ7ZjfxUzGE6SRiVj2nR7IZ
Ww/6dL1Mkb+XUL5UQ5qYViFCprI3ySwxXNfaGAL2iV+iYji/R5jpMeNwmxYrw7hc
le+tT1JUmD5tw4ZbUNWnMR68ATbCuEVDk1ks3LGMw6M0cKOM9Om/Sa9pRUP/ffTC
HAas9QOAZ3BPXm9iMAilDvYqoCK0ny3bvDSoFdmWtsKc3gLA7beKtrk8YPyj1dic
dWZz/HUfBIwCfpPfPfG3EwS3dNI1NV35XNMqIkuJB1lZglEb759+qoyUCUeGSCAs
6A+8yYfyG4G5BBoesusG0dOMuyvzID5odAXTRYDfa65qLTOubQCOOxwNIEWfE+qk
UK5wLGPC7qFqcXyPbnC+mLCHAtB6uFtz9yVDP3hJxCOe0WczUSMr0bwIx6iw+nWE
rgvwoa9wmSmCrwVQ0bhvGNXkibG6plhoawyRKM6MrfaksCm/yW/xR77XbFZCGTN7
ARnf6N2yLWdnsJet4Hdry/iJ7w4voW0/KtlWNhZ/DhlTJ9CpZ3wvz0OmSAW51L0X
zGFlLF4kZvjTenvKJGjV3BHilN1hTSJo7dUfLc5jrgrODe4LipOzUoPQdrQyQS3V
pLT+/GgBvEZbGzgmAxl/yYg8q7/49tLzjNcIstjJUQC86r8T+4/kSNwdMD3nrFW9
kJsQvkYXjWA4wdHt1qkzu8ux13pDpgIPyJ8jlGMc6yqu4ckxb0qRPuPQk1Z6Ck7b
fhqHuv29/+V8QNKP3dnF+ShkeXX4MwL5cvNO5YlGlgFCFihr+59UzWk+ww2BCCWE
eSSlizNcakcm6iepihZuTRqMJI8nr3ZKldE/5ALe6gcPeO8JgGuXVH5jgBLVCtRm
DIw8JZkNqowxYV1bMg2Ho0hSbkcql3mo8EMOQ6y+hSoCPGwx9cywZYUYuW+7J52i
wkFgaI6hNiph3unTGXjjUTNOX9iQVFPPkOM9ANpj1irxFwImpujU5S3gUqM0UJR6
jYosJNaSqRJL0ackq/MvRZyEUYwdjZNqjoxPrlkKhrUvU7I+VJXve7HVXpIn0HsT
F0fnJNOTfcIGTRNU8bjzfMe5ApkE1yEgAULQ3BmlecZ+d70DExTYgNIC9gPfZjWH
MHlk6erT8Ti9O8Ms3K2cu7yqiY0oWH08HYn7nhN5r1PkUH6njjYktcsfXyNuwZqY
UZr53KiVGfxRcFjBzQ3bcVOiJnNndUAwop7VvnLLTcZdPnL+fLu2robLPI96e9/e
fRbBQJA5eunEcG5/ylYO+necGdC37MsrqH+y4CBOWMxUiUdb8NFUxnEqVMC0cuNG
g8wbauLqm1F1BR8S5Q19OyD0YsetGrTJ5Est5cGS8UkSCR0yxKHjzALYoSMfrSnS
hN2Kd5dOf4SsVQLdh08n3NSfQ6LKeqnnnua/pFqB65dYS6v/vr48mtBD4aN6wcfR
jmzWOm2r7FMBz6ChoZclkUYjkfdGH23Nofk5h81/A9vAR5heCiklOlwCIVyT4Dxe
oGLqlBUrOkxy+IQGI3NaYjSGnIgYuZkzFUiYBCC7s1pjee4HUQRwlR7UCkHV76w8
euzndIm0iNKlGu2JdDcT2XUj/8jd6R/ixysjnItSzNErLF5Aziw3n35aTMDFAF6I
SxPWEeLbqy3JNPrINypbrqrzxA8q8cIYswk3nhmYvIbTaTN4kPozml9PeINVZrka
4tbcQa5QclzTpZC7kSyyFoJtKagCPHUU+FqjlRwC2di83rEkvl8BfSylwsFnvwKK
7yAGa0cx+EO2c15vtacHSCXONEaLy8n7s/50bFUmwtwPDd0/52lF2k9Fy4cwtF72
S1OHduRDuwms6PvpXUcLMCeD6kxLra9eqHih5Yu6Fbee5cfKiJFdmKUJq4eIu4HK
SgpjwQPRTVH1GclBQ5OSy8aKu3i0b2e9Tt8QgcJhYfE69Ldadp9Qo8GLpdk2DXd2
PKitqy9ScLm4SwrufXD4n3vnplLA5JpLQawZ38mcOmha85SXlqIB/yDRIwotS6+0
VO8GrOBluUjClHZArTPVXg1HWuIHJQtl2YqPA8OmAs5osuOzuX0HzeV0RCRoa33t
agwIY4VLe+EqeGCZhKr0pDwflthGx4zMg6uTrtRy2xrc9C4Js8KnvCVr6I+KZnni
05uK146MVZr3swzdGg4HFTwF54LPoYcz/D0yZNR18ghoPRGlOyjFGDVzTFBS+et+
w7/5I5Ek8ZYhc7J8H832TXo3mfkQqA/IBwObkb2goiK3BMQj7A1qXhnG4SW8wolK
CIquOTlh4jd6lKWJDGSk5TuSo/IBnbiySVI2PMpO846eQhs26PX78G04xm5aKBMX
3OQrBUroJQyZZWNJbO/vGhgKw/s/TNxFhyXT1A2f9tUn2Emv5x0pkjvKi2guQQ4E
wrGEyv7RkDAKNoXzu8WyD39Lrcujseg1NouJBnQ5B/uvSuu9ajHsCLgDjgTHg4jd
pqPGAJYNXr0En9dqIe3HydG96cWwRV1kdH0xkoUDbUnn7dLd8DNg9qJDXIKVoJkx
m9ZH89/SCpiDXfMN/wRa4Gu0lMIPawko+SDakwa4U0zQvx8b51jOz+hCKR6np/2C
ajVTbSGokUgD5oS52O28/9MwA3CWacvAhEseRviRGKYtuJ18GX/nU8tGVk6MmB/2
yzpw0VlgXtnBshfwtRinAM+8e5oDsbVrk7AoznrTrlHoNvJ7E1Sppr7GCkmplaur
IG26qL6rUUmaTkBefNGUYSaNaOC5br/ZXZ4H6cOGwKBghEq5awli5UhCwipHfDdv
/eAupZWmM1dMDA0C4IyP0j6DVbS9eoaRwCP0nO9ZWhLgiQNJyGBK5KQ/Gki9ZVKp
uciNy+mUrDeiM+KBHf17KUyUQ3CTLNlGHiIfjU6z+Y3umNVfYMrB1Y+gCbXyhpNc
5vONyqu4tm6GR0v4JV0nihxiC4ZjqYrLnI3vObk7VWlXdHO/E2KTaN+394kaeKV8
rAcg1/SWTJ+8wMDUf7pHM9jI6qTomFaq2NGa2XdJRECFxUvM6poWwxRZ29Uj858u
B2bz+V6gKc7yqCMDWzm105dH5bmjc0URbNB/Qp5RAWYgo/8xdfhkteFMAM3JmFxo
XcjZ3pCYIhxrbp2n1DoZIgUjG2bItThDSJcgbUylweOTY2AXKuRk5sIOVDBYvRIj
NX154h+uK6U7kcLMkvxNH+6VcW7tfx2Srvhq+z/Q1KK7/Yvcy8PsXYuKL9WIMHDD
hCL6p7U0Arx+HYAGLX1GhTuS7Y4txiM/9lAE5AwuLpRatmOJrfY76kx2rdatuVGZ
mJLgfsO4tPsTM117zrXTkG/XtlSvKgT+j/9HboUKepAK6R+TOhlTT6LxGSGAjdDL
PN2NninhnkFSEySrTJhb7IKqD3GybRjVUwCAn943LNvSUi6zq836Bn+mROoFab3m
DQ6+85S0akyr36ZUtWCZEainVURK14tcGnSRYJ4JyFqx0seEGGJN8ynRJpVgzgLm
mSg1BGzJ0m6tU1ZLLadaRZTCPIYtUXhY2ichw9vJJbDTkphOSEYnhavtxo42T8Sj
lhOJiRQCotUHgT7/92+XVwEZlR/pPeRZM+dz3MEp7v9oGMSXBuEss6v5eG3M9ed/
vM/KwxvpzowJb45G94ftonInYvzE+6DhafmgHilxcaDlq5JkqeKPA/5LXuyy8D0i
iHQ7pZK5p2ChsNssUnm/dj05HERoccEXtXGOTEDfYaPKrkvKOV0SJVA2VRYgDNly
xkX/t/+fA1uFMCq9UdYrt3VgE9wpcjL0mK3G36muFG1VzXHmZRCbiiioivWWObiO
YBEt550b0rFgzEADo7yeQOOFMe/EoMg2pj4qyHjrO24aRSmDk4uBU5xAcoGJUQuy
TY1lPk1Fu7Nlr9PJADQH9EwgNUVFYCEv2sZavPUXng0QN89fB/wPqmJCpkG6u1wq
pvOAh+zaWCvxlbhMg5mI8KkrQggsO4qNv1YYB+WxV3Rr82hV63HjRr+Cb30Zbko6
0LnBQBEl2PeXUcmt4gVLL7T/9KEI6jaOXB3aXM9rrd0dmXm288bN9ppn8kUp0x3h
GxC/NacNGFe1TjttBV+AeYriP7XL1TyuZmJWTsoZ5IvCx+/x3kcG3HAm5aGhZVLv
Ox/WFqlLBN/zfvyMvpi7Gy9mwurcrm9EqRM7ySUld7y5SGc/s9ysLn9hpUP5QJWK
J5aLd9SzEQGojlov69aLCxDM+ulXMcMyzF5NGEJYFvzzfPsSU5j/lG5LSqsN33XE
Q5PT4VxygCStWTVGzXD02oDzWD3Xj8f4Ne7EsEZnMyYfXwmKQYMp22hQSpRpwKPz
yuaLzOXeeUTNqgFy7u8ATkH+beDBYNzhAZbZeDhiFZVyDRv4jhKC2GPc6PXt3oZt
I+uikykjYdETttXXr4QE65YqevMEMMVew0FnEwwQmZ9Cq/4hT0H0AOyyiBYGMtVe
ObA0I9nhu+65NzKpZmM1QvcGRA4aQ/Qabl9BogMLWu8q9k+hNbPGaWIZMphP4IGC
crBlroD/t0F2lGNcG19XaKOXnI78cPZfRupJy+xjhnn+wZC7//dEt0Ue1mG8hccs
WmbjHpyFfMt/kAY8BubMB86aw+rPCGVr3MIBtI0eW763KyKad4HbqfrfqXT82UGs
GF0vA/fKG+PJnZbuM9kzBVUpTqGut6oRUb6cPjzQ0xouX6UsOhF36dRAVv3m/CNK
z6MKSNRQfJwtt6Gr/WfDAoJRQil7A2Zmi1iBCYauDGsRCEccSJCRujr79pyimwZ6
cRCCH8qqqU39PDqjsrc1o7ZCazO4D25G65y34czZSWZS5VOhP5/RHR2CNhdX43V1
YfzIrnSmIsZgLGYJ5eANOEdjmBpzu3pq1VxHy184w2FaDCbi8QjdyZqU+iisHCpd
suNQHo9gdqwEpd2RpwiO2MiSRGUFpbOZdw3rhsTVo88PmuvEuzevEhcA2KU/7uEa
9Q7dGSg33F0x4okXo/F7Wn9WREEfB6o+aO4A7rfg+42W/NfiMg7VyEfDk392PNkA
IMi7DfcLr8tmgPtz/npgdCIZ3/ksv3EhVVvJw7cVEd/0jnp2G4VWinIKpUvTGxF8
DDhaiH/T94snwlEgRIikpRx4zHEs3j/VfhuocpMlWxf1p0c7luOj1aRsVT+obrc2
Fu8huclDtvwmP2mvFophp5c6txGOt/StSpf4E4FsQzMn22jQ+IN8PLPT0eAI6Nsg
MrBj6TQKvzqEWUkM5Cr5qvfauPom2BmeTk5YSUXHEQYfLDiEqDJvXcV/MfYAU32Z
rnuIMhL8axgKY5tTUrgg94P89eB3M3jonq8Jk7iHVa9hRLrAa+KDn9uAw7sgImOu
sPvATn4xTkayCPwu8+wLkW+vbkVuy7QI9XQ741rGIipNaYQYiBrCGgr4voLoQOBm
p7JUDBelkxFrYfWuGwBnJmujpQfhvwbbh/MygAuUzRcj7M1zJLEc7Z5uYXT4nj6s
tFZ4P5ElFooxUoYrRcQQWGo3VfPvlc5QqzWecIXDtb6KbCyV4d8nd8OMAPD3e3hs
96CjNm8I+1JSOxNfRtKxmQXhIO0Y+wvwqB1gSMrxVyiXh7w0uF3zd/KlHVMVoXHh
/IQqRP14K6ETSy+xFZfExO7zky1CIPMqpwZQ/UmhB+uR9rY9eb3b+hMfbb3dkYDT
T5ZsKfjs+++D0vJ9Zsd0BxOctu4KBmCwatSs3OJoUFBtS+T6zdBsyX529rYRHuvk
XbNxPavpdJHwZEQEZTS+bxADS+Wqsk5NQWt1T8j5Gxsr8ZIzM1km0HnVS+Bv2bE9
kGKGaCqmLcMyKRkV4m4+YfPVybuOatlWotKGEfmCJEcDfl7f2jCbQTLEcJ2wpcCz
YgS98VWZwJE3ErH+UT7NqN8VhNmkKa5+WY9s4eufREDMR9e9D4/26F5tlLc2fjLG
CpdrcMEjOSHHj43OMYIBf9ELU7OYUMXxEopsgkmUvGl0pKBeFNdRXIpgifGwV8iZ
YyUlRrcw4JU+SyQrVJA1L47Aj2LRS14hi29PRohKTm9RJ+Wo4lMO1v4COZr38f3o
lPop4dCH4Bep8tLEvydEHPRpRvbYzZw+30cAICkWTStlBIlfAHLeNJo21mA95h2T
ULEmL40iI8tMYOuG6tNwJaqGZqBGUh0wPlPizhGv7p6h+1FNYBBITXg9mqCKH3O0
B5adpdhTBYgEzoHO2+LnY+TXR+9C5+lg//+Jrk4nCdk6NEEcwZbBBQSIj1BOGVzW
Bw1CHIk4J70fL5dGVzjFIsZVZUik3zslE6yxa6iC5bG9b/22B1UBzDnnlR9k68Yx
FRIseyWxATvtZ0m3WS8ptYn0+Vkah70wnMAHRfmDe6LksX7o4YqfJcXKDkIMwfQM
d+mqZQ6hsOveAtLYRcFnjcEMy0WAi48Gl+3TEl5Ea6fgg9qJ2BGPrnh/CVZPww6Q
rldrloOBUrov/fCiF+HJtm5RWKFSDKGRyfdJGJ/jR6+YBsiP3EnRx3vMhb3pGArS
oI7/OELjNx5MF75PyxQB/KW8h731JgXvERWy2c50MfYuUfcrvnHQUwT5HIY6brFi
gsYghvN/zYyxqXfoehFKICBkrssVVceM55YJBdvOHYQffqNv+EooL0rvUVGuY9ry
XRRJ+xTL6u5rYEe5X22zIgf0fE9ZSGc87aGnMm1SgFp8rLpKbc2IQlvNLXETBMxb
8iULRb/F4j+DUAvlO7mPpVBCKJ0JJIetCUb6VeIcmWnN/pNh/RuTE9HTbfOzuQCO
hnnaJYf+o7vqsYLnOk4sjb9V6XjnSj0yYu5qcrBvaaaSOivkrpdZBrykOV1lYH1T
W6Hc3rmm9cGmou9sUk4H7LFYEMisFo7FuuhhaRhUHRgbNxMDCnhNPwNkhNDY79eK
nFgXiKixUcetUfM/R4vMQBAZz5ZzZkVQfzR7cHya7pt1JA3yZ4qwvVk1na8++amJ
vuY/J5qqLO4pbZDRy/84l4tg22Twe1QJcceFslVzbluw8eaFl9DRwIfjQN7l+qeS
Fyf9da323FYV/GRlsEOA83xHPIdzkFx/SMl10fAMQ2xF+NU8aSkbFu8ZV2clPV9G
mcPfLp8xflDWqB54O1bM5el6hoppKVH/dTjsPn/ZBkSViSkxW/c0018rqC2ErL4F
ZURnNJ8GiHjsjiHgzb3djFj8EJmECCuHXollTC64+E1k5UwijHRIB+JzKjJvz5rE
If1sFmlL11eBK9KZMxG1Xy0ies539kV/abywh95ghc+AEcx3ZVWutnEpP/Hjody5
s1H1m1LlPOhBEGsqtW7Tcn4rKUdXIHEMuhP+cXBjnOqPb1TwxoxtvdeYigUxtnSA
XzRDX7O3x3CC/W6nndGMJRgueCxTsUA5U5CBuEj/6L415OOUYWgv2dG4gM8eVLvy
YadqjA7W8KZ2r5wCuzGrH9rE4XBrAZ6PzWa8Panl61iw0GDaZAedr/z744ocHpR6
RyH2Xaxkc2hyJPxqpYNWNybDwTWCE+U3YOQVqKp476aZUvtR6hsyWhpx8qLO93pI
HWffWFFBoEtnfUDjyRhvBezjyl2chBD5SwGQHhVlmo1In3eYmbAy5CtOM8ZKtQND
P8TT1Cl9ekQcotocgqbvaVH3bTsHxLqNVcMdHberIrCoEKZvosg75CpC3+PQLVxu
VWa6ME/HT4JbW7D5Wp/HVSsPHqHDwon/zaTcLPza3sMUmShNqWsJXxKlPoFOIUcb
sXr/wG4hASlO9Iw7sxXLlE/xoDehogRLjDjjesOZQgYD5/hhybVnsFDLZTTjlEkU
RGhM7MqmHFNEhfbxUFEFkd89DULEBzCGpdswgO/a5ipos8HWgCqwcX8Sd3iKfCfN
3xxn14WnvFeOTyEbq8kkgYKOPNLw/XY75+2niOqkavSdCqIMRpqcK2GkbTDvqDTw
Q8d2jrOji5wXBxE8miH6M7Z0Ns0rstF7Ox3QuWwDtNL1AHPL2LpXKGblFpz4G8et
BIZg5KW2FuMKopQnKFxzqUh93hfll03b1daKgSr/5a24ChKiLpCvkK2GNOyhTzfS
KbscCYhAeFK2I/oP4i9b6quO85Q14dfoDVk1oK0bd7DR8v4A1SfiWTtxoPOdAnJC
AgZArJ1zPJm2dqvtD88MOXy4qqpcqWeKvjADesZWRNP3NJh0c6l9D+w3RnZLsHzR
FfLu2n517I3UkkCkYa6WCYUtekMUi5nacOizB3IPa7u5qpEwX8RT+QMdXCUor+0V
BsFmOZ4/yvGyjKi7FL598XF8NvyTlmb6rYgiyv5GYTGxQX0lOO2Moj0ZZddJC78P
beymnUYPQgmC/mzrsgmxPFffd8kSQxBqJHMoSkNgUAA2tht9ZmCHzNIkb0lQjajx
iYGa4TtNmXK1StQrCwBFwQ9fdiC6u3VSC1MZzhHItp3akmFa31+OX2S1Qk68KHY+
Uozj+L/WcDLW1T6gXglmyCEBV8WaYRXOIZM/9h75FquBHNBikSZXgpuOH6vzDunt
BeMGKmI+510cwHVTpJqhNcjL3jV3SrZvp/HR2/jmJ0bg91HyzIudkf7Dc/Y53EM5
1XJSwplO1cMXdnxTStD1UxYtgxf3TKf4FiSCdE/bNifsfsaXr50cywmzsxJCRdYq
lr/8WL8PQhr7rP2Sj2/EFp8d11LceKICwTgD773zSUNEKd2+dYlN7wKsVIL3dwcD
j7gBrbfXY9+ifKiYktFd+DeU/sg7keO8gHxIESisU+8GadLQ4OpKIjoJdbgbLuTr
py8cKtje4MaJxlCi6lL/IVsqnyYPsGnES0mBvTH+OnimtBT6KscmH23klJPlnxKK
gZZ1iPOQNKV5T53WBQqTWFs00lUgYYGrruRqoxm79orn2yKAxGDI03DV8dr2qwPU
Cu1IFkuOR1zfBK/4SD3YXBJR8RezyUsjlao0MdNzgKqynzhiTNuhyuIBBjmSnmdq
1M/0YkRwIuNNrvClp4Bzoam6J1bvZ2G8g+8ompdMkkbEKMFQyYF/AHaNNcI2APQz
Gfnl4qey9s9gRp8yhVW06359nVa1SMy/BpspP7MbKtxqZUV7THqjY8yQuLHlsW3a
MDoYZkwXYPt8cO20qna7bjTyQYtm13jU7g+8CiizRjlHRxYORntOgy05CNyfB9Mi
mdXJvw1m0ocfiizfP4QDQDHsi51tzGA8I2ghpRx8NrhUw7LmxXmr8TnkAAuPhFD5
TiD/C8Ca8ItC1vg/cUX8cVYVsvtmMx8fKfmlQpZSNR9a64Gn3xalTtJFcn8ffZZB
5ozSGn4Tg+NMj4cENHSfZ0guD6hdGEQPQ4Gj6RKzoJ5pM+igM4N+l++nu4H9hpWV
s+5BYZs4f6pZpYPJm5eWNHwNPBa+B6eECZ89EyNVtnaO6pU6gqHBmOlJsgt5VGFM
kb7dU2w/cNiPcxrGz/6r4Zyo47v8eibBii2Q0WTnNqq2i9BaoZbsJnIEG+oLdmZi
4iKg5w2oC0B5kmHjWN6vGh8gOwgsNKXDfIH6MJkevds2rVJh+MAdmdLdnD5ZvII+
0DHZAYAH1HfiyJ9sIfod+LWjqFcYRv3BWq3n2Fyn+ANqvCwbg9hyUXHCLrMuQVph
ih13edcLpBKEkyL+n/xP7V5xx7kq0KoejEuTEqp3iVLPL1C5VzWuSCSP2PGIGUiz
gdh//+fVGq1GFuhJJ5Qsm47R8QpCR6Dtq6aVNyGoxJ1L+avfP9ww+NIW/BCXy9Ka
RBWa3epoW1CYNEf/ZphpaybFoCN33w40EkJD6YMO/CUw7f7zXd2b85maZnS39z2e
rsunuhqeopvvbujPzIeinvB8s5TOiq0E6iMHlGzCvbmMehe2LVmEuXYimAU1AAKe
X5+zyB4r/qpkoBDkg7brD2sgw9ojozsh2JcAvbFM74loUWeRgb6psMczbARDXdVk
PVfhe5P7wQEE/hmG054j5U80K3G6zh9ZCPpZr+WLXc4oeU9GSIgQWdWQiID1D5Ns
DUCNhzuf3ICcnJ07cgNPZhqfpaQRlC2ADeN/byiwXOV5k5q4O6kskXVDLlH70hC7
rFoztwjfJwq6Y9/3/Eo4iMuvT3CG87efakpkdR1zrs+Tr/BPsifEfeAn5ZWUWdvY
RYnwBv4P10O4EZdTRK+3txo3d80dfbp32jaMdcPshRH94zppfONk2Abq/H+wAoBj
UOmqJOA3FNeIPeuGXVj1dO+f/YCKcUx3/r6MRQEluPDYvLEH9AsX4vyZY/a4yI74
mrTQdCW0s0pwOcjAM7xnMibBi3FZlM6hX3me6mKPUk3VQzDlVdg3zxsFMxCa86Lj
YqQsAOQj3LQ44hoXRkKAri6bDUtBXTNvqe7aOKHyQHbp5CxeIFF1PaY8nf0/aUA6
hENngQBNJ+ovsvKeBjQZolp1ckRI2NXtGjTk6IEJnRrTlAx+IfGOoRTligDTVJjV
RsajvYnqcvpDY2VFCW8dnf1FI5smaCRH5n9gCQIdyNZOmpGMK95b9ULGSbcY/7MW
HLHtpdCZKkb/IpxOCP/zYKjBWEAFCp+GusO1W8ipC/kjimRxykyqbpowCjQtmvps
Ro1d8XdA2WzGLisB7bnFcEbjZCYOdjUcCyID1nP2dp+jRqTDJmALCSwtimBhPWSO
1mcv4ObWi+orXGGuHDy1OYlAt2JkWBpbdt7I6UXE1jHj8pymj9gP3HnX7+4NrfPP
mb5oPb4QObplBXETUxJVEuKkDe1Ug7WlzVLNM9ouvVMiRewIb3ug9yjcj1Vfu8vc
cbFH1kLfezH+/I0vbqopQ+oODY+SHuK8VRk9Oq8uFYHJHfJ2rSDU6gNI2ryJYkhi
wJvAbDz58Kgziafyu0+gKiDAuujQcMx0XlaAZHyfBjeYrgV2XL0vnnsGx9vXiE7L
zg1hVsBZpmR2TCvpTsZejJfCaQVU2dkt+2Rxxm+XrvWWXjNZwLZqKCiK3gS+8yfT
OLRn0GoFwJI6QVcjuIj4PDxRigJht4MtJ0dvGLXK9KBLxIfIsdnj4/ReDo+rXWN9
T35s56J9l3fyhTQCHP3gM2Qj3tGbIoeUYpzgMiRTK3wO6DFRC1AGUGdR+WrPf9TH
hxzhPwFeF4RhYGH8mHLWiMQwjC1yN1Uu30tMemoxwSnXwoaSIUoorq+7+LVHF8Eh
3sL5h7YfWvnQFKDiCHHIKQ4NfrucH8w/A9KCWA5zIDpYEU/OTFb8NRSsu7tMldAr
qTgSLcBh/ltk3bMniBOlhf74DEunDCv0BLCNyEHeR44irKHmc7z+UVefICn9MaHT
rT9+mp024mAP1pE2Hc0D079uTPkAx0Bme3BKoCtM5uSB+9YVStkyNjYiOKw9Q26g
2NZJQm4e6tDu0hx1lXJVmEE2Yjur8W8Qqdd08bEijnQLsUV5aVOpg7+XZtF681Y8
TuE/JTEpfIORcnzyBkIN4k6tOjN4avhoQ3zcolqzb+HAi5j3CetvlOO1WVuUSFp+
hiuSRdUMQhLEM2/jO6eSguig1xcRQisMrHshlfZDdP5H+L1S9IHTpb4D68pP27UZ
PyKVQFkyAQRNUH622vZknnEGKUuFG2o2vqBjrsX3GwLhDDeYYz3UXPCAgCLOwVO5
RXnaBYSW5Opy0vI2gdabTXVJW2ewUpUUcBYJHRLpgDTgQRRmWy3yCRcFdmIQFIXP
LzW191jzu14xZwsd1DXtFMbSW2/GytjX1Q3RKeUJ/wzPMtbdDc8B/pONfehDvDC3
qFqnhdv0LlwM2GKTZE0thIEN1B91MPT+SXtXfXbHntaJHjqmOlM/ZcFepF6IWhb0
bncIiMMdN61HKlXK/QdIEmliHKo7FaHWzmLA5/xFq8DOyAmbyk0AhDPw2XkLbg7e
ejWwX0p8WohhOiO9/HE0QNd9B7ndvk8M8LDJK3D9Ki5XKK22h/4YHW7WaeUoC1Ya
dxr9jzv2OpcRBQeNGGq7Erzx5LOcjcMNBLi07zSEkcia1jcT4dLX8rq+0Q33Movx
InqvqdaScE+VcR74JdrVM9jvrgCjouu7HiqSv48b8p9o7Y/yFGeVVqnLEEn6I5sc
jVaEvhUbGGhMV8QT2w5xWhS2+0jIjO/vFRGZBdcWXkXIpTUv7v0/ghtz/y5HzKOn
K2NpqwGKKmSLQ2kOXBYxeXIm7nOzUl9YqQfijaIfqlYQljzhz3K0uvPFz4CiTUQb
+qLyPYEanZd7EpEli3L2iyUPfZDsQ+pPPB9QxZMirytUl1PaQwMsEJUqguYAnsKk
v/dOiksSntpKW3HkZzzlKJdVTG7HF089zRmVr54u4iqfJcphRHaqHt3trnQPd/Gh
qHIdi3CDaCfzjwWSmDlyt8ugfZnoTN3VVQGR7uoKYB1jcKv+/TvrTqo2pL24ZTku
O0ebK8Rn+STht6heTN6k0lm92UauYuj+kXHp0JQHyBrpCTNQiw6VwhbmOXeAGeE5
nyno1yCHCz2GCS2VmnSSaMnhhwuCh4wALz1kbk/pU1Y1t4RlDB98MZEXlrXVoQA0
hRZFHHhefeAlg+gy+TrD8Ti9yH371gfw2AQ6tdKLofrM2Rov4dM8XgcwHU3MX2Kk
ar19h4pMZcVieVjM74cKFWCXQ16cobAjTq58tLEhWvSoEsNYs0A7+lAB6D6GAXgW
+f8y/Q+QbNM0Rr4FA9Cf9oD7TJsT9Qv9xqFXw/jHmXvprAAS3YAwhR1mUvyPJ4Ea
EI4/1auFFe/I562SS+GPhvljoYEkCUJfZtHsJG1rNo1MgW+rh/HSMKK/LTn/a5t4
VeASDogRBk2fi4mtl3RlIEZJhE4W6vYC5UPIwo1keP5AFyzJGbVrs4w7zC+Vz8GF
TKz/80lYzjG9hZxQcXNOBgt1nMy4nsanCxcz/kZg5ejRpA7a3Cc5lr9Oc5SBN4Wd
X2eBhDERgl81IchbJw821B6xcgsB0RLO6Le0z916FndCWjb/9SUJLhgOFmAgVc6c
s5WxAKY106rdwVAbtjSrp0z9//MoIiiF7Ocx6cinDHQrhhXP5FfmJjRd/+ywtQtc
z87iEkJj5XRVYI6dTEqjVDwfzu07V15gkx+MFqK3t4EIYSUjeTVbR5hcBMDBTYjr
ZPRf6eiuNBn5plOmm6RyEr+5GYe0IJ4sIfybM/vuAw10cv2kk23ypOwEimr5RQXO
vKotklI1hnRbEs9JmoGpRr4EX49iNWIDsV5zo20XkyoyhCsh2k1ew/paapsJXST2
jOJu2jKx/ltRINjrWANA/B2oMJAIl3THx8ihazzHtUYSEZTAFJbAXLF2NKE8uNhz
yBYF4YUeAqfXfrPCtBNDIFWj/eOVDiE5M30TzyAPqoonszty+C14mE3xFJsXJsbs
O0wjN3t7WfzVuMJGAz7MHPOQHZt7nfjQe26pMm6fh3GXzV4zPuM+LJYQIAPpv/uw
Kun8n3EF1Khuou3ef5yN2uxTtgqbweDcujIop69++lQ6Ej5qtnRJM8LeyFESd+nn
Efw6J934vLvy3lGgYCcFNT27aYTPQq5HzR5J18LnosciOQKRjA+pyk2HN7u7loHz
FOI6Wludq8fVkYn6ShhbeTUOIBBgZP6noGh0BtkR6CIYld+AthD6nKQ4jWp4sEt2
u/EUty2J37SSNKEqgwFY3k4wEfK73vsWzfrUjrIXH0Y/mKqxmEqvL2xsKgMMjDg1
3Fyd+Sdp31G3H3eJ5gMIDqHwcq/VINjWh95JjKij55NxfSQ4a9UCFILqQ1I4gxrz
pXulIvJdVq3OhBWiKoLNrM0GgcsU05vcYq+gubqJRqcwNEPy9Jn9ZhVDR5HTRLn8
t4IYKHOYCPcgzwCcySPf53Rg2KhKzd+d2aF1Lc/IBhZbUhMr3W80vl3AQqRs1x25
DIr3j/YhE6Bc3Ywi6d7cZ7KtoK00V1lDTMjgJGz3KTQ86IabZbfKKwn/chYIEghS
426MoifiG0gxGfYr/+T3jYj0wqAn6/0/AM/LLGjyvIdDwO5GB2Hk0wkwzib5OiX+
WhOGSiGyF6z7sLlbp38qQ84GUXD3E1cCHYCg1ErYXOZLYVritMYAzRCfQmsdkFum
gY3toH6SHwydu2IMiEM1OFc0KkWlY8NGRAlWTJi4XPiNJiSjiB4/+bthMA7RqF/H
dt8CKBn6KvB1FeS9ndyFLhF8W6PDRJ03O6jRLLV6zn6n47krH8km47AD15VjAujQ
dOlC1iEwpRUIzqokC2foMN1lLlycdsUR0uRWDAuX26rUEUzzrETlljPFtCSRdtUL
kSK2H+RYl4YrLoIpChRBiAfLLBKWE6Obq35GbBSDrl6ELoO2Hf5scCIZn4EDAxU5
B4AG5yXfX/BTEvoK8fWN/UrHCDyLW5p9GZp7U69cXH+ny3/ylx/Zyn9wC/mXovZs
SAY0OuIXjIxHvuCayk0w3FBjxpMiRaA0SjlFrz51BR7USQn2Cgp9h/1Wn1k3ah2e
pfJgHMB1KscvaYNc8BVVWI9mtZBqd15Z0W55DlKNkTK0PdIgUshW6sBKJiKmbk1r
SBoh3HK+wiyLEdaXZmLdku1IGrWELwPiFVYF1wW3QiBAspRdhrvaGzfnC9RC8Jpp
C2I2WJGpveV6itMe21f5ClfMEZyIVF69iq5NN4PZb0jGCwguXuqqdU6k9qPweCKy
cRuTIq8L9YwAjLeoRg06Es0CVX7XQmEEU/rKxXU3Pf6OjDBotkiT56d6YbjPPy6q
HM1HohC1G1jI7DqHtC/F6VpStj+Xg6W+qAVG3JGQPmXha5yuFg7q8sDXjQVjDg5w
wo6gK+dpEwUTJhOxx8QlT2Xk4joN/a7mSe8Us384iVrKQoo4lpDVUm9e94Et/JWe
2sm11H3PDrQrSBqEFzUb8RVDJ7/rGJo2Bz9aNXCw9/MSXmWyIZxqYrrhjHJy0y6m
lc4wgQTDCQm8v3O/T4dfxnrV6qV5aSI4FExqkSlWNNOHUjc+C3Gz1ZIeoZ2zR922
LBtCoCm6AbslUARLOymOr+5WIwHEP51f2lebsmXIik1WNwVcxxQqU2IIykT4yDDO
2pG5jK7hLWkwNwJUxeL1tZ6iED8l8ps4MS0JvszVqkDcgb78E4uZ4jLjabVNm5TM
dMIWAbvqmxvwBrPUaRNV5JUk4USbIhCAYt0XFmt9QGY9KWX/hoO7swstvCzP1VVp
h3M407rZOq9ZnwAtY6kXFs5+sfqGLhfyxU6do2Is7h2YzaPRqF+0YgFcT9361X7U
YWMdusnMYuu7jZkS2hubcxUWupcAES2qeCCGS4+cw5EZKK/ulUWIxYw9BKhYG7YV
ERIEzyYWho3Esuu3H4mIFYTn23jYmiZTjoBnYxEAc3wrl300GJxfOVKky/ics5k7
aBY8tk/lPHZd3uxKtwMKehnZ0ziXR1FBIjeMbdbht4pRXgXI7hArw0UcdDZbgpht
uvPwE0zfkCikXAGknBm8XbDKmpydXg8W9dWaI0zm023pAfyhobXBtCrIbPfMSNWt
ZIlCjx53UsO7h3XZacNox/iR7osF55We+FEhWnvNtQTs7twl/bLWnG3N18Y+AOkA
Y76uiNF4+gBxxDtuwf7Y3p/Mc+R5fcvEYdZxgxf0CKUkitbTGpoLMFvcAV4gvD8i
WNgCPOm9fcWj7O6QQ1FpTIGVObb4oaQok1BxZHQAiuliW35cw1MUekdk5oMhtBYc
alDW7mKaUhO+H7Zit2Y5ei4YjSm0sKqdcJBcv5BQb/OUScFbPlTMQFyfA6prmYmc
0wRgDYEvr8LlTBGqDtqq9NC2PJeRqL3GbBBksjXHb8ZSjtl8Z4A+b47fpiUHgNN/
QXq2M8mZy8fU55lu+LN52HDaybPMjGpOaxtGoGumUBstsexaP8b4arBzGc4N9XVB
2v9TatzodUgwPtKFO7Ktd68BY4XYmV7xbp2IEtwUG3MtXDhs3Gmq3kweYQvgiKzp
QpiDzYsuLCQEZYFaK/0EWfx+O4XK66g+7CdfRBic1umy3L1axDO6+9iELs4UgvZZ
RYS4V2dxpQ48LhEbIow0zrnXkV6YKb1fQKHkoBloXyc6B4o7I6IOgpvLENEp6bWw
o/x5OcnB2yMH8N3ma6jxZFgz+onwsZTUWlt5WculR5bqWXQ04WF0Q58dr69KpLpx
/S98MBG4LuMCBJGPgmEtNe+sdWL73uGhb9nOjhTLxpIM+Y0I5A25SycqMGxbMyCo
6zO/bq4i3NwTBG/Ft6tAxMtORLETWdj6r6RGS2wYRxRdH9y1AG/tc78wdsR1UaiS
f/yIjzr+4ixdwFkCDpEYpwiZTpPNMQOjSizOvFS0WdKQIs8MO9OaHtPMvnFu4XBO
0QAs/tmhbow0+6T3d93NlXUHJvlkOoldkegUP12NZe/UPur+Y6Xk7wQK7RoCB9+u
zllsWxPy1di3ddUuFnrLYfmgL4FNmi3msYAkSrDrOXhAUEfb+QwcKT+TZTShBqMb
WiRJJVvJXbUS23CnaIehzYQAJqHyuAkCK9aHkA/1gdRT+ySkSQvTsBCx/jyq82o7
jh2w8z70D/HQR7Cxo4be47Y5uoGzKcXm6Ux1ktQk2Dp7c2tM+7Q2Y+HqJlb/Prt1
Z5yMVLpg2D3zVmtRp2bUg8/Lc6OhcAd2GSYAr1KhNVvWzFWuf9SKkpZrYC7PxfE3
NKbyK56/tcZax0xcghMkMHGq4j+oKq6EWqZgXG8StBPrLuSzDtPfGbE6LRFFQcCB
iSy528dpS8WvnTmhv5A7e/7etzOItRvmxecH1ZAUZVR6VCsrFSDPB2NyX3YIC28L
inRN8o6Q5Xq9cq9DX1A9cwrekZnHquZEL5fT70bEDVNoOgWyxUwryff7Y56fC4lC
K26PmjB5asrS0MHpy3KyFYJJ7S8ej95uz7YaGaZyUEX2Hsfx8SaB0B/+osK/rpvW
HtO0MaxrSJ2g02nIUZ0yIoXDRBwCbistRBcbOmsWVhUTvxdlXlFNpSL3ruXMzlxz
oFADfbODIsCcEt9Vl7rlhsRqZ9udGIkmSaQsxEgqh9tgC8Da5v2sNHFiQ2kjpkkP
9y0qUbV40TkbtxSZG2DKQizgFF78DLCfDWNKcjyQX3REma91ChPjFdlMCanr9TU5
K3u6bKHNlY2+kMloMfi1gc+MIKjUoBZADqiWF4Z1U1logMF1LGayh9sgndOR21/K
/qK8ZFC0uE/zYjdedZyfVKY6ON+NLqbS2VWO2EXlG9+3Q8FUfF4TVW0zMVHr3vq/
0UIXHI0Sbovgz0kEu1euTIitNAuS3hagniZXwclZDiXouUkT9dhNVrPNUjnhROVS
IQukQ7WN9DWGVNP9aWir1fO8hvZVBosj2cL5XQems/Jf7Op8nT7Vfh4tfGUClasV
wBoDLaJVB1crBSIuUF4+v6kmshtPF8AsqNE0nKoJ2T6UEXOdCkMt71bAwtjcBYeY
+4w694S7qxq8IhdU2M65nhlCi38DW4HEQBszqxKjvi0FidwdTNK3Dae5M0dcLMct
/hZ+4rbN3/ztnrnWD+DdchVyY4Abx4gbxGN0p4C5Me2fIDSo72ize0VxKSP4qFdC
PN1GFVqk7P9xLqR3V+44VfCMIIYF6Mj8grOrG0taL42ODjvyFsSHJIA68Q3/DB9p
OhjQcVWRg66WRrUlPPCjDwWvWMeT6XvOXYcTBI2LwY4DqvTSFPzdwR12RcTCR3Qg
iGkETGykDWg4zgLLqRlt1D5DlpPjc++Nm5MV8NN2m7PyN7+vwPWTgTAlDe56a0D+
SM6MnB1kaJqUBFlE/kxRNN9IY8uzlrs1AiQ3QvTcoAC8gdpn35QPmQlJW9rUzYe5
+VK0dQGRYcovUZlEAWgA7NeD8ING0CcZ2/MLa5ePhaor4Eac4Lw+sAW86Vi34TFR
ZtrIeg2Ty5/7AV+G1C6r7RrPTaSqlGx879ef1naOFK1DIKiYxAGkG4nT4MUFiz/E
30Re8NQMNO7abfqPJniUz1nzKrBIH0kJ9UCcMrNccVMKSFx3ABIVVTeReu7iacUf
M2i280MEdPIK9tNDM2jFAvTswxILUY+treDzvS2tsNOJqDQPj4BOXWqRc5pb3jLH
BLiQomxLNNQPl1f9C7PJQXJw2cOGftlj/Pj/I043G1dHhF6LyKbaO+qlxv5gTG/H
TkmkS8JVKWQzENsh2Xw5CwVlZY+re3RnebotJeHt6jckYcd+cx52nG8DbBVNmh8C
hjgGriibS1ap3XCTAFUAM6UCz/8dSCvCOAXGmM5Bzjm3kX6M83KLqNPzdSi4bDu1
CHDyGNIdj9QjeGu6M/VS4KG23M/oeqJgk5xvPbnqfDyj9pUUFxm5T8ESCJ7Zk1al
QdqwJJCjDH9UbdW02k+/oA3OgK5Jmtlb1inTjkyg9aoJjLK/dtrNMWaBUzXWiNm4
K28gcCPztC1N0AwsYU2D7C0g+zOVLZInDy1S0f9yErLgXkzNpPI+ZTScFrn3MOhU
pLyatjsJ9Mnzk0dBCg91l6jMte+V4gUuY8XgxhCDixD4qvGolcujyQLWf+8z0xPr
6dit+ruy3GI+UPKnnWBpMEXp3VP5NstFpRNqsTRHyvfCS6fYHo24uMH/8FgRVKno
Jqwo1c7Apgzjg86VFGEyXluhyjru3mfgNZGZmWpZapbKg6KU68TFnBy+yr3yD09A
jJyy1MdlKqooz4vWN77tQfLs3KDcNpyW8s+fjg6pKbYnUyn2AmZI0kcGPzWx5NfO
yznWZLRTeVzCSlO1dUAMFWw/aY8195e7HimTDYopTriFY+wM/TJIH/37FKWwrnHo
W13/QaXdw9dSmGOuCYCak9piMUVYkotqAvyQpbwULq16qNBk8GOUqXvx+MmIcWP5
kxj0WBuAyaxGv5Ep6jJ3g8x03pSiJd1Ux0c/QpHDqzkbGzzzIWrncXYoDic/30QN
cW2HnHn9Oz1OtwKJmCMoTOLVFdOLrHZXx7iugzZU80kT8UydWjdjIO8MAZCHZTvl
GvS3ofu8rBJGrAwTOHmtke3/MZt8IPlQdJ+I8HDwDksUhI0wWjBSu3jXYCus2Hvs
v47enbmx1Xyu+4aOcjqVlWnDO+LWT5LyXpZ9iRQqhRnoLtK4mVUbxf6PLcGN5yH0
54qx0qUDut9IEEpCUImwIxDj4okjvaqJzx8cj5P+3jwgTaw0P+KmsqVLJ02Lh7he
HsqhDRKgshijuDMfFoWNLUnzCU4b/W6mMbjKik73nOHYCZIvwiUyeMAbz3QTt9rL
nSlMzaNzE3TuEF/98sK07n2RJFQOOhC7VGIce3D6zJz1voYl1rmGCG3y4kGBbaaM
/MSXOW1ixwlJwdiLusulMboNRbjvX5IQlM9sKInxSpaArVVxwkYDapmwIBS4YuCp
4BmD/ZuijJSHuHuNCmy/SojOu55/UFaWdEHmOJ0bFSfN2rm/tK30SslOccG7mls5
LQLGZ3io55dzhSlMFPbQob0wkIgyIVYrCVob3HJN7gqQYQmx2sPIvr5L1G7ZrHPZ
onMUXh1zeGvBrf0tF/2j5PVZel8bnrx9gtirEt713ZH4jPV0+5m+IaffN35/e4vy
FwmjFHmBQq+HY/zl+pztdAnYTp3Scgth0vwEq7bWOBnPw7UEkl5jLcdEcxlD/VFf
yk5uW6qnF9cAzLDg2Ixtn1dlwUivrzejmwbZUzmSd7fyxGzBnmJ0awOOA66b8sOF
SJs3yUshbmZ5GN99xaWwwBUJwa5Ao2fYJlAixypOc8VEp9rkeG6L5q7DS2vapn+E
vhNu1l81vPxzidmf+HidoTpk3DqQfjkHc2UJBBnih0yuCZ0f2PFbUQHciXuZfCA1
RsnHgwQaxXi4t1DbBNfDcweDm5BU+OSbm/h/U2sSsYWe2Ava/Zpx3FVBZiC0UV+C
sGIKQQJ+jySahKvhZsj55Cm3xEoX0f6gGysThV6BY+h+c1JS1xHbifplD5wB16tE
Oij40P76obZ6ycviYBk5PpenKV9RTcSd7OVLbYP2ZTe3vcWuMG4VaQp7/7t87+8W
3dfLrq1QL+LAGWErcsM4Jh5zIs5nMGOPdT/7jq/IIP3t3eWpEGVjpR6e8udyhSDh
eSFy6dBLu3M6EMmmx46AKxyP5I+wJEQvCkdDMO5AZx/9TVub064NU+VY/srCO0i2
elvQuil5c3iT2m8/2Op+H6dtUphn9hUlHeMycbltzbfSnpCyTw8ziXT+nsxDJz1w
kpiNF3ILHJURiqWF7MdIYVQXoYd1lY7zZdRlK2vZVwv6sYDqfZub9xZtVnxIGI+0
66dDRVHAC/flwpJ5deJ7H0JHInEygpig8Lk0qRKkRFEPYXhi0hnnTLXXvaOgA7FN
G9UpRxdlg4M49RmMznkC59p6zSmNaVAH0Am/FA0AbrlnCYKKjAS4D06NnFmtKYk1
16CuYeVLOjiIjCwjj52H5zu09ye9FCGB6v9o2mUV7JIrvxs25ZUC14IxApS3cpJv
YcdZPU8BwJcRrZFjEx439JRzvLTDwXTcB4i4akJmHTHTieHlyzLF+JsL97oujtuL
Xms4Vy74UsFB3R2y5I+8AALM6gh8DeG+ndizf2wXVEpHlGTkx0MHEmcOG1Fb/xvC
3sYvoR8bqPFLbXBUgNiphHFW4vojUFfdsYxlAonm9aHTH5DMgNVl2Y8EIzRw+Saw
ZwZIHaL3u0M1MwfKR1ZPr3lJv1qES4ES11x5QSiOfBebCUAyN1wlkzQWplc7fuIm
hXnaJ4eXSnq1WHqcXI2IP2OVtPGiRYGYmFX0PgR0M/vnkRCc+twlL6j5a7da7nu7
GAZ+z1MdGcFOV3QXEoYKmroV+mbTId9AH4Bx53bLs+/3nZjHnSqFQMvStGSjGGNg
z0T81dPFsQidotzjAa1hviGja2VAMw9N92/SDPMYAEpXFLtLxJqYcXNIY9RpeQTh
U2UCBlwkfcmWEQ2lXRUAxWh3uQeBYVjx4CyEZOvpS5pa2+7oQ9oDaWr2SFj/woDj
XRmFaYgH86QYdGNz61SWUCKiomJB0CVgPQMG8HZWUb6xXkwsXkXheT1F/9HkBa7C
l7im26Tk3We8837OW+fHbynflHI2LzykTHy5QDJTgj5I2LgyWVNFsFZTTEzuDwdu
dHo97zv33T+LKlfeZgN1GnsfM5PBkJ8bIeHm7ttWq+HacPmE6vENJiOik/cUwNow
uE/0BQCmPFEFg8qeOIpWG4b6Jag2WKcoYfZyIH/zA1pPofgoOAMmkDwxvR/WtKxn
tmCkwo1l2iHNP/gEwAMUFLuR4B10cmQGPcuJwux8FitcB3rdwILxqBc/KBzC0iZ6
SfnBAmZffJ5I4Bg8Te889Lf877gzr6WCNjl35CEi51WgxN+nrtwuLSmLKqAcYiqp
uZk6LtnBt7iOgwzGaQXzkS/YwWyNmiUqP9QFb0ulMWLYJ99uitJv38JoEJ+WrCvD
+yQg/28+4M9SyhAAaSrj6wGjurcdtP1C1xprEHCj/vYOr7EePgurMzzqMy22Ywiw
vMOMdHWG+ffBaRtR8ZtGqeK9470spAqwPmEmzusvwkRpzDvwemRxE5pI4EScskH9
gzQAMuuq3tfqZyJYrcdw8QpZ2skKHktrmyFBJCBSKTeX5gIGpaa2/wl5ZCqXQ0g2
jw+hfwmj68xZn1JLee5YXZXOHaGTCFhYfV6e9awWU6w9OaNN6ZCINnUGZa91RmV/
W0V/03b3Zke0ANzDDUohtKB+BG50kh+Hs5KGKFcQYuCEF/CtRQrSHfNOepkYLa3m
oSkZNvi4gry0Y85XFYqRkzxGecRClnrWF3zTfpVa4aBbnFJCI01GbDNZ9vfpsLV4
/7k9U70qDsd1VaFE4+gjSK2L9lhbekMBl8pYsqxgMkUU1i/KAW65g5MAuA+NAMPK
W+YMn/roAnozpcrgZPeHLrPBfV1YcDBqKYezBsTDpPy0kE7Jhr6ToufWHckIS69A
uVkuxpfA9YPhYarp2MrhAxCvcl+TOeZeoZwL8V7X3RxGUFrNgY92GLkOt/gUkp8n
v4+3wE9057JeUJHZbOxWZylAeBdVzLQN/2yqmEFSSDkvFo74TXap3EmqPkJxoSD/
Nwk/Gs+kLJvmZPX/t90JMKR2/hYs0rFylvdpJSNcJ/Lb/UlMXVtUAPgQep79gM1p
tfIo/NdgloOJim8snwF72cqW8MZ1Yohrm0e5WI/5oEvMIUm7hbAANASbwlbYKQco
Ok9dge1Nf4ssjse21fjr9ldtRJyWQLg6pmmx/17CaYrm3hrx5hTvcJMJbvEYnHo+
Z7hPh0w/QpNrYqe7KWEs8MUfJ7wJQfcY1m8V0SyXBPv0DNNtZQ8gKYH6Ph7JVbAF
KhvAI3XWAf2VF+Ni64jmhb4AaF1yxNPoUDRA/Zcf+vPH//1r1T/Iqhq26N/ivZcL
keytKuNgK5DWI0CdtjcUGf7BjdlBdduCYt8q2EACfEh5azw6LBSav7053VKoDX1B
FGWxuJatSQRNgDe6ajH3b76b71iqryzRQfW9FkOOlUrN5emTMdkYMFiWkD+lfe4O
/wvjG9xX5aHfW/TMujw5H9RGiDEhIevB5TWhxkeOzVZaluQofkLUvO8x76n4VRkn
rFRaw11bBzcwhbIHRqU8NfB//hTyeyrlVSd3YjM4UDKsT6/RuBybVPQm/1XoQNOt
v8jUVhzeER4gXUtGkKxyix4uTtqfjb3Cin79RrLJ2U4mdV1/EyQxKuRtRSiREbUl
nW3EFYI8sjvqLEdHIq1AddzZNqfQk8GpJluptyGfYGoAcPzH2LgcgbIhL00nrdcM
vKWVO8pGStU8P2bCpwL78zHo5HwZoDR91gN2unsDjac+Y+WRlNLnmwJYsa10TXVJ
L5v1BcVWhGyqksbEp1JAzAXro1mcikDEuOqFzni8ogy5f8vOogv6ZHZ7vqjZyjPb
7kkEKC1OvaJXgMpjXLrdhwYQZwozCpBGqwQKIrlKlYkCvxyxb0AyQB60BQIyARpq
ed0QYsdg9avsBeXmSY8ll8hm9hHgUrij3UWKZ5NbRQ8FCa5iS76Ae+8axCxmO6sJ
4uALXhtHKwRZyJ/RhdDRr192TIElbdxFBjg7FrRxelzfkDSj00ldSXuzLlqlNWtO
9J+5lT2KZKq70yf18mP4ay6V+ar9L1I1jZ2LzrGF2yvMKZNmynH9ZzBpPM8BFxqL
GbsMloYSLHzYehuNmiiasrW9CoSKfTQykbTn9F5W0PVyGfvXvRsxoKdExSDAUU82
6ZSpUIMMg/vK+V2ZDH3OdtxiOe+4nk86XR49E4gKDwoBJVP0gr0RRUXoEvakr4yb
OUnxnZ6FYqq0YcxT42RFV+YC/qv9rGsfknLiZ6cxHRzlth9t8dIfrGRqvbaO0ony
scAs3LbGZxy6DC8iS0v7c4QJKI/3JEYqo6CJJczC7SWqHNNZct95xnWhGbCpAMix
X96Tr+aPzTOKxKGpGtfAIqbCOz5N5lGWe3zoofpu7o4uQoxmUnEhlGgk0WpCd+MB
NyoaR0IvfEnO96j5GIdKLlxYLW6Xn+qvucBtuRDN6Z7so1nnKMa3tKhzrQvQiD9R
v5oqhzn1qMSEYidxtGgyM66srHF1UmMJ49e1/FdIgxfXS5J6zQcBIpTrtEafC11a
3Qw3cWNzE2SqQiBx/Rbz9AkYvhuAj0vMeRIG+b13ssFkViHWDA39xZ3fHLKQjrGa
PMoidj2Nl8bEFf+p5LCKiHDfnlf1043wrbeVWgcU3nfiqC++U4puwKAQ5564Es5X
WByEQ7MdCx015w0DYejHfqo3cwbKhrbOZtOB+bd0tvF4d0TVjxKsnpRXm3DGHpoc
okpO9zYjC6h1sYUOwssCSs9Z1JYZ29/iS5tVtQwF3AmT/U2XomvM4CdatBFXBioI
me1tBj1e8tvzgsMVOHP1r+e2zx8ZRDxsWaDxTPEp1yJMdjbC8U3FnjSfrhxOcZQ/
YdWPu/XrWYOItc2jGO2D3l16gqt1AtRTN3G8uT9HTwtM5xsOqN50m0emPpUpdS1S
kv1jEtpeFle9mZdMx2zdpTZp/xhPc2SnWYpbrxxXsk+mpirwYqVg6hZpRnLRf4QV
kfK/Uj9jzYISwh0VBJx9iqKodrN8D+05Bvr+7LHzm+jlQ9yQtfKpYqb2VbCvpbr9
WlzZRWBNld9snMlD8nk1tY0zxSRtiC1DfRxaAKIKLPrK7l7Fwe8GfKZaY6VmEfo3
MwGlaDS5S543Lgn1DG7W2tb9Cosu9BhTuMZiyLTVEynLwzk1+yDHvD1W5XaMuugk
WvPXGJ01Quza75qk2lXNxj+dhN7NXIHy5ZH94J7WjnKw2OoOofrSEgYEj4Bm7qw+
8qIshklxfOru/E8bqQUv2eJTaHQSJkbcltn+5VcmO9quykErnnbacjMHHfTtZ9aC
IBBvR02FnDvNwZsZayhgnDZoXNG8JeZD4/ZqrFqXdipjhEBODoGwBS3xTkLjlJcZ
8SYfn4Ccd70QS2xbVNjAmS2xa6g2bWOyJTLCyDURCK+R07riB37fIUskR6C3sNnh
VsDs3gEgV2yxtPXrL7myOtY7Yjob4l5uLh5ffE76zTBS6zrHVU8XsXAGFcHpAxum
MUuhQVIoOvFKzIFLchCZdTESzoDbVm4BJZ4Su1rnowoA6glcnnyiV1GfohfOC89F
ZAhbMcJ6u5hbtkpkCLUPFRjp0sh4NM22xmnFrIz4QUcs4qfnCA9/eAR+Q47MqvQS
p5fjEZpDgrFeya2kP8vUCLWeFLXEnkSv3kyJJZpJ1IXOoAmSojZir1WBQQp/xVef
izGq3Yb8ekyXWEgZ4/4bWZBgAJQmGyDAHp484DAzaR+zSYF0pyZuURiC6wJTb061
ZKh7CkviK0bOt0qaGXFGzqKvSkAcvTVEZF+3aFKc+u+qyjlpcwy1g3M3wj/D5g68
QYAEvAbjXUIZYrODXHnZCiOtvk5KlXx5oquARN35q0Xj99SQZBNkBzS7WV29YRnb
2l5GDtHTUvDm337cDXy+peS++Rf8na5K2vlJovQUvcujnaFYGm8pyR9hE6tQl3kO
DVlXqyuHhJnhG0ag4LN+erVcz8AbT/IfgckjjxahXIfDZKNOk+srbdWmEIPQ+042
+4hdI1GBMIE7eMsEJJ7NrvKNd8sGdMYk3uVKqSK2mkM4n2gzJSh03xaZIEz8mDa9
9gpU1bGchVgzX7/rvHO/J9i/TA4dY0CGCRdGuXqJQyjGgMsJQCKhOF9PDSkGWomf
9g8nS3upOH+bjQYYN2wo6sh1kapr0WJOmn2uTUgt1/o5S/pIQl46Age1KVP4aSl7
bItMfo4uF8b5CyVpAQ0wTS+sU8GsPd00ykzBbuNvNuXBaQIBpJrzdKNVK69AAYxI
R7M8IjlY7ZT07a2+2BrCQfnOIxhspQrUUV1ZVZjzlni2ipg/ddXhVmBd3VxBav93
x6KHCdCGKa66Y5cw96kgm6uHQ4mL/PIoi4jzWyFOK7HQMwqcBy7HsTWUu1mCmuQD
NlFgzZaYFqqvZUknlDBeXHyS5ter7UEB4gNs6+OhmAIF6UZWso0GBN8btNOqbodP
i+HUPy8zsQtVCBOKylIrDbFEzA3mQXESNAD0KaWB/OlDNxPtZJ+Fc42aURoIRTId
IFkMphQi/tL5+qv5bGvunUGLLVd416t8TCP2Quu98a80VyeeCnCSPY7cMK/vUyG5
gLQjEb/TiF1/G9EHjaDB9AI+b2xqK3ad1tUQZat5ObZUm7WF+79pblBYj0gtGMZA
nPrOFj8yqqegILHHBvs1XWfdO6S7MPi1D9IJmv4xqsT3zh9FEBj/aCn0eEFiEwpP
WHNenTTdL8YI8VQ7NNmms83j+c7sPANtvzK7KQhWDPuaM373TBFvqiENNiCMbRcc
YGnLVwL2WtvT1NpWhkyg+MqccEAPEGpMBADnHJDhl7hncz9cIQm3unl4wXJnf8Xq
Oa460XLOy4bh5H0fyfsBS0UD0xd86197h3gjqQVYPLJz/tGTeREnd3cs4DnSV9Dj
S7foSHPHcha3ZT63f6xn90JeCa2hYuwFhpazwMWfK39+gkO/4kDGggKjl77EwyxT
ZQM+OvY0X08hDLVGv7NkHDjHtHxpbRYwZYN9Pllk2Jku/qLApa31QwgCwLETdCep
nyH035JuZXcEEwfzmi+J0daviIMwRZovAnAtTSGSCTOFZm4wHDulqWTcU2lwb9XR
TJbytCTmUoyxtuUe73Yx82sXoibsi548oS9LzsT3XiaCsQv2ntQcJ+aiZ4wr4I0o
rdJ36lmpj5ZQEvxquYevmPBk4VPJK7im2wNHHKBneG9R+lIZToN4uAhXFbpHsxXk
FrSn3cJ6CM3lAzy6r40VjbbVDS1al3ele6dbdLg3Qjecs1NaiP7tUa2Hj88n4GYc
vmg8Hd75C2iMPfu36PH9Hi/Z4jz3oz5iNG8O1dtx6nGIp65ofSe705HAy9Z0XeZC
WTz1LTegRXPExvGUR11jk38MBavAQJ+C1rxtjh08TLuukDWVXOhnKQ2HapvorDGT
5KCf+mRRjEqEm4JSb8/2YRCT6RKlc1+mrbmXv0Xcb4fHz0zBQU9MoFlexPG5azyJ
ueXAjhEUgUDWHmuEetvfQmEqan1OExEVCzuuSNU9O/GvGxk0Ahim9tfxvyJ82h8R
BqpUjgLxgWy8Ip8iFntGMh89/Ben499BGozDuXXrJUvmJDzwc/b1165zfCg2RPez
+3W59KS1RjfRxXsOJZE6a+5t7uzVuzmide4ajKa7J4cdTPPhdPOYc0mFzttQIXrG
XXXEyhtEJ6rli/bxeQ5OjSWquN2VqmPShhDEy+ZW5Ju2Hi479oZ3oeQt6WGiDQP9
ix4AvqSoFz+K/3bP3il57fQGoank70WYimk7sx+gXRvpAkL0yAmwZDLwaacyOEyh
dRcLNwcvQHNWlZti/PHU5wIt+1FC/y3DZjy3hxxh1EI+tT5fMt0gNslGIoOAMEND
gVysYskEgfY1sT8tLwYTtygnjMpI0RLXOG4w/Fc5jGq+R88NaCH/NanKPFCcGAYB
nrKpqsKJTTTfPYPLEsfVCnZ1d2Cd0vLzvaL+aOgBdCuPhnXojr9xr8zNdOFRQpO3
XadLWIQl1q991jnIHg7URIfr/ry+aQVprl9xT21dfqh4zbWpxWzTYGTCdPI4hDZp
bPZP64DtO7wZ9Xaj1B8RkpDq1+MmYop8Y9fuM65T9k426YZ8oZrT51R+4s+y8ZFx
sFtVYd3OcJAAnDID299xd89wCSR8r8Vc3RW7VmXBH0hu+tNACxtqNfqEuacwHy0D
eU9ewSdhtfGXkT2PLzAau/x4FGa+EFI6GiWfMWQLHFtUAVRy6PFWuQ1FbxK5NyME
ptSz9yjirgEMynVRk03eMRxjoQ1gAtIXzc8WGKFy+8tmQ/uCRBOPooDQrMDeUeSF
ySthzVcGrIgDgiJdR9f2Eynd+UcnTRzTwXJfkKNXGKRKlBQfx9+EnTCPdVJxIgXV
Ks5zqMH42rjrIJqZRCRMEue11cAcrXH2nc0/n3w/oGEZ6vZjxLSPblI3iDgH4WCb
wjLWNH9OVhx32RzA7sAsvxABetUHteG3ZcksLVPTvbz4q8RdJ/x/xt6d8BqBcxKd
xZkab2YASAu15GF//xbGEBC4oIQd5NWf3vBzCtbNHVrcVzrH3GJw889wnQchGbV8
/ba19nObFnAtFopVYZ1DkaQy7KG6tc8cFDUeIveC6yygGVAhsKv47vdlC9uM0IGI
gooDQkW9zCEdCxMmt8HkaF2Hu3UVJXmswORYWauFfdCNNR11yW2Z3LHKfH2thgPV
Gic+0WEiMmBciT8jMzZjI7v8kqlkux3SO1BQv7Oi2Ig6JgG7WprPTAWwGVFtCh7q
D7IsHqxNKcB4jbuIs1kyx74IeWvJS/+lcMdHY2EGUBT1RwYOA4C5uGd8ZeHyPtWx
T2xRi2OZTuu2sUx35lvAIwIO6q/Ysfpg/cePIEi+0dZYuU1trbGM0/PR74myrdEF
n1Xn/oSnKtiLTYxzTHEF+xOdITjtQG9OK7x8nkVkzNAl8jvls6gvU7sasK4SMH58
sZr1gkxAd9Rdjsp0JzopOdX9kKoMCNbOxNBtnZJEAdN6Rnt6W+bgLJbU4IWeBYUw
8XNYEftRnM546kry4nDzd97nQuOpoXwayY3ttujMie063r+FHc0Q+gkdgc0ehmIE
ISgQCCBXjpF9I4USZZ/dsGMhvCvfE1TCfDke+TEg0e98dxP1dF9FXklZg5Om9nU/
bQvYUz8dHNB3Ej+T9MHbsJbPhV+4ELRarOkgtgeoAZAxZoV9iyP3rNbQEB0Q+kvj
A49kwewHAwx0R+fEwEwDw/v5fIk5haqfSTVqHI/N+6PeGdCTobAL94Jj0yXTu3G/
CI40gkA16iG8yKHN4KdotvhpjVtBWmLWHzx7m86XvTCmQGu0XbAUgD0ihgY4Rgr/
FKYKkCp+/qSy3taJCbvQWR/IXpZs22welPwwmLoLVBwzCpBZ8XJX5jUQbHKUfopB
UGACch/sykfQKfjPly78xpKvvWNek9qiJk86zU5g9Sf8VJ42mKFlOcMLk/+ZMBkC
cLFXYOhP729pKNXBP6UrjDKg+QABTOOT+nUzF7TfQiDBfwfobs6rhND/pT3uqkxF
btJQQve/iHM6XGUyH0MPwgbssOKR7kLfkt7VP8WfciY4FYfViGMcJHp9smT3UOxH
8pNMjSs8+qskD5CdJVDtEkJb6ztrmJsI7ATy7i4sCBHbvR1C1EnJXkLSrwnDRCRS
AW3EInvJkUpcPWofuwbkIS1ZbDmIm+dK9NfWjGyqVs7ZAazq1i6a3WQVcA5UMDZX
HQs8jN5gbTmg+uGummMwcUlQOorNWqI7c5R0FDde3bKuOqxYxO1QxjfZPG49KOj8
sV8NJ9erjMzIeOZ3+Tgy2OdpMz2wOe66nJbgjq4gVEEJNG6Wft20JtOOS05v6zry
ZVU0u95SYGVkNo/cWZtk3pfmVa5470cj0l18Jyr1en+kuWnZBOMZkd8eYwOBU/P6
Spkf/uL60OVT97ieK+rnhwMHiOmOSXKLuTIS3sA1xVjCjSzzUUpfLMbSOTHNLrr3
7T37+O0vLsYzycFfShNh+6D7Jz4g7461HMvutlQRr8ZO5BrySOJ9ivkJZq3dYXH4
G7Dzm/sEPVy8A4ZW679HrbjBY17PP3CIY29r8ORB6AZ39exFxGCKv8plsRnQLrQn
zm0EMTg5zHmmjffoukQHDL6KBBwJA9f9XwQ92RnWP1AHV9+BrWOh4gRwXC8Z4f3I
mfDv6ign7qO55XrfbWSx0okyIvR5VhW/eBm6xBsh3Qd6N8U6wibgYZk7jcEz6WWp
GaaoCRaj9BBFAelSSAKJy4YwwByEQL0UaUj1zwExN2LJusLdpCbGOQnhx3NT+/Vu
TslxRer1mqj9Tih2eXVTAFfcfWoLL14D/U31NgYa/QlY1u/IK56/oDezNhP5fLlK
gGYFlg5LUUFS9/Rbo2IWmiJaHSX0406QQSoyl++IvubSkSQ5MRadlG5X5Za8eQwG
J6qH+z+Isl0CHkoqoZkqaAMLtBB6jEDG7Fze59A/ZG86teUGwl1cgGG9SlD0dHym
UQbUnBfMWPTlkfUQLD5ijoJdQRegT0MTheq/qD6bi/m0JugqY3xFt7mZ4ITfA+Y9
H3dtUeQblGwWLMakepgDdjj9qcuyvQ40y+m9r1Y9lYVHCApLDQqW2PFZQ5APYt+C
P67wGAKnSZCGC15U7RFs7MJ2FaxWf9PmtaxX5BBEVQqasc07NNLHwMOg0kOSHw3v
/yChcREx7o0I3CzHiD8xWEFzFZ2ZmgTGbJqYfoeq9PCGLggn8qgmlptfwztUiuBp
krUP0MwJxQKyAe7km/IpbY6VCJxIdaRwIJBBG8TWrzJx47n1HinVkyrK3YJBv4v1
5E6SOWbtIzaU19K2eQFPot67FCOMroKQxhPPmIYnyuWQeL7HIrqlNpcQ8rCkWk2A
GOrUQ/Trp/ZoAq0oGaFWw0gptOz2U+u8uwzTOJQMlqyuFbDqgICbqo5izBmM/IyU
4TzycEWLgJyUchaqKS6T0z4Lt0MEbqVYCCcZCkKf2c9yaDJ0N+dr1EARoivgMV8e
evUb94LFC6p5XLrkxs/J8wYPeR0tVVIr2qR91aXtN9gF3xcgGVCKmkg/fNIF2OfC
TllPc4fVBPNuxTpbA+K2N5B60r6EmDz7R5vr22KsH14i9Mc7xsZYZiJORxcfW1Ex
2x++eX2C+7Q+GeZvUF5kXnq3oQf27qZty5DxqyXkbDsr/jcXqqWoC/1hogrwWfxn
v4Hh05kGx9L0WlkBshXujKNtUYsS85h+vHtdWXWg0xCepRiG2P1CNkBImIsrnyvx
gfm1kYnDaxQCJ7CbCiP0vYejc9pv/I3wGQ2HXWkEjG+4Q6X80u0DOj6Bzupo26Te
W8DymXia8symzNMWouthMLX2dJaYH8eRUaNGPm/lLzHI06RKjzIcVgU5I0lPMkJc
Qu/WHwZo6KdVl7jFNoHWLKnlTP6eIisPQTRETm6qlm2W8LjdiY5gVAPpL5whcEOs
W6ogxlxaDGXFMGut/84IIEcQzhZYzPAQuxLTcRtPZYj01ki+FHOwp8M3d+azfj4d
IGjd7o9P6PDR4LEE0zby2ugh8rAk+pX6A4RrWMEjQyLOE6zuw3VLWUqZhHLk/07N
rO2tK3kb4Qgl6a99yxYuh1d02dGv9icIZFXtEnXLEOA3W8O+nzJd53SLCb/FFxpa
ZGMjKCsANvLOYj/7pcdVhfSl3IAewaIKTfIlWA/gr2ZDkhcYqzJ75ILnvbwIx0jm
dEYssAWHZYAYEmjRd39Qrq+ersNldVt6DAvV4vpAVTX8U9h8FpTBMBbX40WPaywx
cfdV/PV6NQresylhDS2JWXc6Si+zuEi/lo02s54uchD74GhmNtAK3Rr+p+hV1HDO
8U5ej6FQL7w281T7mebryBE5j5pWPsyYs4miZrU63+42OErjlT1LWnd8NqRoUcce
QgMk9qhAvVm9aLaxpZHimvBw9xgcN2UgG/9xkRm1TSXagJ2rg4Wnw+RXEoL6lPdA
JT877v9GwfNGPEtvw9JWpLOyGfv+JsAD4oTvcAq8sd3VbseI/eA21qXmtflMonku
puMFfQnFccceU3VADHGiAFx4Ah6fPxnSgRG8vkPjhQUn20OhEEOm4YQIL5ZMMbrX
/YJADxIu3eY2NXj1fgujqHri8kKu2pPMorNbiNjkWyOAMSQ61DsEfZXYFtmCN26E
BNGwgVv47w0Rw7f0GKHEiaIz4HYkCdbTWqZ2CknvQc2ONcT7klULIpMw6U7MHIr8
0BlPkq60l8oRwscitS6OakD+nxxJ6qmRSvB4I2EhehMoOdyazs5QnRmvXd02sFnA
y6g0/i8LqqqvjJGL+lr18iGc1D/kNvek+/8z9IYCg1qEAG3vXS5Ryj5JtHXrI4AW
i6j7FHfRRM0Rxl3qLiw6Rjc9s5Dp2ojq+nE84g2y0XmL5vtun8mrjLs5Q3O0I8/T
JUoUJIm3i2EQHOYWXe5pttTFWl6uZgILcLwgm7OEOPqtKfTQYU9frIgmmPL4PpTi
s3B4RQGOefHghPDJKOapAoJkfi73OvK2svw+SsJhVkDRYfPVbb3tI409eanSCSGe
lsxjPiOvFlc3ITyxMaxhENNb4PYFBP6nZrhcgYYRVOqrA3bvDQTkbx2pAG81pVGR
yR4qIZNNn2GEANYWS7TpFOzzM+9m5pCwNbemIuw3+A5ble8pFL/ho7WsJzKlr/tW
JdswzEoyUuWrItIPG3BYKgeSh1/oJnDMoHPCR8S36uiAwME/jWHP6iOeBZoUNNRY
++zFx85rkuV3oxzTTliSoVE06FA0sBHaOVTZS5LKhZbm4yKgGr0lEdHpSh39GH8g
iH8eVC0HIwexG+bPVWnPNYjs3a/ykig7Bremvy5Curt5BVKUXqk3A95HEQUQjiNi
VAeNND1dp3XHljrtyoOC7ONiCeUVDFhTXU/Nh3BeOi+jOkamrTRajksodOCq7xSv
kRMxba7nE9w/Wkgdt39McapCpvYX1g/fL+M4Gj2Pcnqyur+58CKrbzBVzclRvMXO
g6iXclqdKbVb+f605RPNuS2S9OVv/geuCvx9l4RunF/fIyCDhoIby3xJ7NcAJUUw
1c9qYf+pAVqXbOVs/MaDii78YmyN6uS5JmF/zXw9aP6i3Gcc3ux5oiUTnRbx/Pvb
PLs+/K0fVJ3En6AhWPr6D6TlasslkqYKlzvb2PjJmik1Xlos9twU4lCmEkj1EbVi
F3gePEFK1/CByf+4a1tnvQ5CEjqS0Dco+nqnbhpVFw3YuMBd5v+VtvnuNCNumFNG
s/0wQp58nEPaP3qJZ5uUw4BNjrvnNAl4HosjuqlubQ4G/4JXb4hlCXVnqCkrrZtF
4Q/M55y+u8XluJWFF6IOTLak6IjoYv/9tAhiZPeeWh7n7301RucBYxrAWALqyNSZ
qDdcHUiHk3tBisaFWrgbNilHMBFEtXiqsRbUxia9C5WGv7tDuXdJ9KM6gGJoyrkX
LBX3PIG+YfzEEDC/KP/MBA9/PyVqrar/8jcEYg+JqmtyyJt82MoFq4JeQHy9jw3S
Y2tcXMoqebCqtMyTqvghTNWFuDZ/pdzMeYL0KE54304W0psJZqYNhUJQt7R9UMlu
HcDhn9ErpEZN9951DgcwAX8JNGzFVAmnpHDy3zBIcO2LYEjuzpWT1UWVXqsKYLhY
qUk8B+OvzENd+efp38rwWMX7t3FhV3SIr+feVl6v3TitRLs+nLCYUqIO2wkIY/Sy
Sz+mDLMrXjkld0YDvZEeDFCBoWIGttDd2W/qcmv48wJ7oCjh9jEJUj8f4BFkC17g
CWSNfWmzKFf/dtwggTqTgDMGjn7GAXrZ2sMZCsmlzYb8XwwDy3q2DxTmYCLj5/vX
BzcMQVvx88w542hbJxx50YPxd9NpQDMmjl89xPXHV7vf5xg8TiYZWLlO+b1miOFS
EXCQszbErsohUz9SeKI3+3CfbojZf+yQUSiE2L6MZZvgYWKPjSD4nNP4iJgg2B5w
130GZWNjRFbKx/UMUEdCvEMlylXX8VcL+Yj+w1eM32r486Jpk1Woq0PVFPNzS9wi
xd0EzObc3P/v+SLKouT/9dOnPzWm04XYNqzYx2MRf6pOcugGSWjE099yRRzu8mnQ
Mwt8AkoTj3asGhg+lmRLIMcsvPOINSPvp0yfFgnst9eit4KUC0adR6FXXMdFrWZQ
Ac91RPEs4EfHW7pFJ6ORh2oFD6euPVXHPtlQx8OAT2bNCSVG3YsZmmXe0vVL2Tr4
PQbGDHA9ya/khUsAGMLizhxlqIcJnl0yg/ljqa1pJssmc6iQOqABJ1Pi/w30ZCRD
eBTDqvocUMN4z//yfCJhOI2zd89lI6AwINYPBnmEtfrnjN0Jp0rYe4UHVfUxTeue
EeI2Kx20V9O7bLiwMAeBhLAbmXvk6SrH2CGf76E4onWoxJQEu8/YDBfR8eJ5m6Jk
myURxlgyPAKa8wc5P9xPL1+SQcaIzNgmd88ag3/TIljzO9Z+eI4DNcqX9KKjE4Of
dTlj0jmDO30dKm/kc9FcTEHZSowAdvuCuI6z5QDWMGC8ggcFS3zWdo/qXto95CJd
6rH6Yu+3hVVd6NkHAlsCPkAtTDjAbFrNDibb0TVzPqfEihRT1gpdtyTh6/yR6Izj
j6Gl/YXyiLAH727T/DTuIRAjWmIX9lbMR/7tgo18WWDC0hA66KljouMd7zXzfE2Y
kDgnLXe4XNQ9XIgod78B6KrpcTbAAhQNp50PFg6hPoqePSHNPFd41nfeluI4bRcV
mBYkHZkM7vC+kXpUMfAr41iooE1Ed9KNJMXRE9I9FV6FRD0PCw4p5afpw/v87XG9
WVEJz06U7fr+cftO2HSasREXKTISJJTHRhKaO26xum1Z3ws6UhKJwizw8cv5X9p1
CdXgyKvuO20W3CQm5jX+TVtVJlFrMAl0k9HIXBCZ579O/+zKj9Va7w1q7V8HLnrJ
ZD2UXM2lYSWUUQ2cOvOXGEEmqphZzbW4ZuSo/AGUUbZWcYdMsa+7DoEk9dAD33Ey
Av/2+mF4q5LLWMxfNcZPsS2rjwv79yer+38rXwrR6pYGD9rYzAffmjpQnkcKUbj0
BZKvfs7IbrjDQ+VQZ69KdoCVMBnEJvfFzkpMVoLZhf6HePF7b6xYK6BljzVDdiRh
idgzU+FS0HHuIimp6nzGpjqmrsH6GBl5VHrFnmcTyX/XpriGjjEiGzD1JgGRAD8T
UPLcSbkHziRUZxvNt0X06hI1q7YCsIKh1XzvqmgAPbvB3e3rXN/cTkKS+Tyd9Nms
OpaFcScPdRgbVpZe9dmfogAwpGzILUR3KFJ1bdO+FnmoXPZj9WywyQvUpTCNFwmS
saI3P7e8XM9ceee0uDYEZAYMuxvpIOJDNV1ZGEk7vWVujG4+JFMxrhTT6Du1ozcj
5Pci2pfeuOD7djFUlpGrq7ou8vAi1K43VbGjc2KCpt4yKmH5s5YOqGH65L0ulA92
UHCoOp3gZ7ZktPY2fDnU/NsUuiNVCxsmITRAJvbLIlh8g7LFQSA/ZKtUoZAD9u1+
wTVc6b2tx4PSnzPrGNVuWnvJrC3ulj31lwhYCYkw8NvnjBLeKZNI7dYiUuuPYxWc
/YgX8etorWDhBWr7hBzEgN1UdLZjeaHjInq6rfL6JorOBl7r/mCYYkG/qUghdGy6
lLsT+W+by/QHIjypxgCKoOE3YsY+5zPnwGwCjmnHefpfPZIA+pZ4WxV+tNcL+T3j
iJp8ehtH69wRqdXEMEnpK+dPR9pxPThOMWn49Nai5SIXe7ya+At+mbijk+YAqG+6
RJKJTi5xr/KPxSVm9GIBE2BhNzvC6d8bwoJVrFJXIyvRx9FNiAy5sAWeq2zSHSr7
Nz1X22163X7dqJOrrGLbxkwDhNcYS9+OFe4AFg6PDIFzZH/8ZH5c99tONYfuip1+
ZJUDU/nmF/qn7v233QT6v5b/Y0BC8kjDOEWE213iNm3WyXBDqzP2TE5Al5BfWo9r
exF4ZgGvtWgsiHRD4MIHBRQcH86mYZcCZvlnwx7Zulnf10Drh4qsUQCYbZGUMaD5
kmXEDFQ3Khs2NPWNAL8rPnU5JFgr+NugYKncYS0Gm2D/As2CfxKSc94G94JV3Gx+
BfaGNoZ0mEqJ751ZbWK06XQzaH23y6yYUFzmFpOzD0mGsRR33pvdAYT3H8GqxHcL
KVpprx3fNhXFyTTxL95jqxrvrNAvWJ3m8JdxrGT4vij6zdlqShJs1VhTmJ4QB2N9
a/RERnOPWGbx8HyNg3/Nx85yoIGur8YhGsAatNdBRL8G+Ow7G4mUuhgmOAkQhMDx
eW7OS5xiXGNyBjZlLjTH5QL37YNjiSvEo7tHxCiQICB1SSoT/gVd4Wur2aeXZeZw
OIFLtLFWlNbMZEiA2a7+CWabVJjVnIqMTv/aaHA2rnoD6QxENkw4tBs3Q5xPnexZ
WvXWfFckRE2ehdrgyAM0t4tnaqcJzzTv3P/PnlaEL1McQOo+niPtOQ6I+PZQj5As
aSKOHKn+Hqd9lmEhObM0Ikk881MBGJeKmSlo/PZ8/SFOKBYty0+9Nod6R7ZRIB6o
TnNg1/AzkFY6NyVJ8Qy9ZNDZRl2djUkuIsRHYxNz++XxWZSm+MGQ7e3v4Nfpwy1L
rF8fzYu8+yDCm8pTrlIckd4UyOm0SeuYqALC4HjwUQ8OlNNLK7vTiXwh3Nt7sRKU
m35G02fUCQjM6mlV5kodAMH/dEMWBhh8uT9i+NFD2cPBsc30HUyKJ6r8OJJkJKrK
nv6d75dktsL8Pir8SAoEW+7odGWaA+5e6YDWVX+7FA/SJxuiY8barqxE2advU9NF
xTFpMcr2r74cufBGu5OeREPcGrxKiOYFR7qDxpW3hz5SRX1biw3C6mPUsPSHNo/f
OIXP01SuhWABeY/k0zSrY0U7ahDYYbVyqk6kSR6yiasZNumYbL2hkF8Sz/9lsPba
ZtrBLrrpyjGykd2LjbmvNIl06KMcuBAUr1H+UhPT7myGYyBHy0viIHKVkzizItn0
vSdOuhbQ5lXBr2rQh0Vh2HTEiE8B+iO0TH/i64XRmnsxbbLJ+hYXGerVGIDAlvDf
eWvt5k2RiklcrbFmTvgNknoieYxqaONBWN5a+uSkB0rOtmLnS1VYIWgeTwg6L/ko
8jRcrwelx6R/6AzLPpHG2UeIwvw1ht8fpAURgRGK65CL/Zw3xPiXg+TTDufdbc9u
/lD6sF9wYys7wCCxS+LatLIjBPxutOKKSg83Vu8OaXUh4g8YWXSXNGLqKEOnwrNH
hi1IZ3k/feGpmVfGh/rmPhoYOnP8Ui6MpZuLu83R7o4jt/V9iTo3nBLjLW9NNyem
23IcFifW08l6tVFTyqaPjch6BdcNxAtJqHpjg0kXVk7GyPRQja/kmMR6JFu8MB32
C/1bj0sAVM7znQjaE+7Vso8P0XiQRmIt3R2y+q95MYB0u7lGj6BBrxtwqJ2VeBsr
a6aREl0x4JWhQtAB8wRCU+XpryieIQmDujzG0k16xwzUVpkzHUogfLKJMmziqJT0
6sBz+ziMd3BULmVqsCbdh4ufsPmUfksPucJYUUtfsFsJ2Lb5DZbsB7IWqd2/tf8l
Q/6L9eAXvdZqZEjLt0H21Tp4z1obltpzd7W983jBqKE1n3nl5TAvr2J4kQL1c2tY
/OAXR81o9GMAj6aidRcUUEATuErf/6an6Av2akxPmKJURbQS70wNp6HItq+usQDZ
VG/ACM4BtSw4L0c1M4sPCCQHxd1lu9EYPREbZBqkYW3sC3k78kwIOp25j6lgl+Pt
fsIlaOPSFqW5Q4rmN6VYjFWAV61Cfm6z6OMYf1PPD+wAXfPJ3mVouxUWlB/54e20
Z4pRrBtGnHszbRenzfpD5/7tHwwg02nPSVA45+nd5SXvhH6Nz5FOqBdLVTuNtA0I
wGmu79/u9cZG7zZid6e2ABI0qZ0ckF/DhkS6ags1Fhnu6Rirk+D4iAiK6UbMuGAK
AOeWAH594bMjFDpD/MXPOV/d1WOen+YDB7WBrpAOM7fjR+f9dmpcHorM0mZPWS0R
slOL2oR7ZOq6zDLdzXHrp+DoGRHPQjY3I3+FYUUJArQw0vCPJbfT9yjWWriG1M1n
2GMcqtsQ8JE9F2w7WBQYHJq/mjutkXZSgzzysPsHlDfXJa1e930JGQPZN3G7UpEb
n845Ys4988TZZnQ22mFqGaLNsX07BFydlWRNEHskUdzh5O7GtkiAHA5x413D8FCb
rLo8Q+ZGalsSM9Ktlg0pvWru23nHjBFXhUQwm7TGEzjk2UBtdbfM/i+dEDR3fs13
FefahbLvl2Del0UVU4ydQn6XSiYIudIsE6+Om55ws1oXYOVQn7zisvqJefMzOQmQ
SLx8f6oVpF95BsglnW1ADkeZdBBbCzgZgfQrGcOQcx3ptucfu5KSf6pN1+XCv72T
Y5cwtG/Fnr+WwjQVwW16GH6RKqrLWlHBFxe6ClHg6mGCRyh//rnodEKyqxLwgMjr
68+6xvFY49gFg66icD4yXjU9L0GHEaFOhONAe0KP+cpqapnToUYEXmpJruZpxMFt
3l4In6YKzCZ8GH4pbgpv0PW+RQBLubu6QsneD8SLljlGrwCtRp+LeEARQZqvXMJQ
ym5xMy4XBlODrWZ5LMYE+esaSYyQ/Rfkqq4J5vSnebrsxLXXAZGBNwur7JCIJm6Q
deV1h1gEQyO3enZK3Is/CIzn8HMNUGmvsVVGsjQSZkxJJUqoqFwlhfup5QfCchNW
XMqkIR4uOrKJxBH1u3PR7W9pqyqukKyTY88gxcr7GFhX+J+ZL6i18xXzhYWJdrHS
0tcyKFj8QcN6MmxgoJ/DKYN5Fi7UF4ubDxBv5efqdazrnJQ4hubS39qY0iTujjoH
oA57aN5ggqyX63ehZWS3l9oKPA72zDbkS8khTLil299EA1ujdTIeYj1bBykmGi6x
8vSpgLFqD8aMk6z0vmtOylMMQt3V7ybgkrgd5PLo1iy5+7wOSu+EYeDk1xNhP75v
QQ3hd677caq3Dj4ypMwiQEoGAhtqbsrmy/HpYl2h3CnXedrBOjky1qbQxUfEL2ro
5bD6lFXKm4c8z3a7H8Z1GsT8WfJ4wbImPKq1Tnu+pctCz6zg8pEvjiqbjvmxhoMg
7gBmrso3/sMEegDdStqmEtVpUCnMDfFqxhYGWZX2mZA46j6gtbHMbffMxCIMnwOm
ag5DLM/Qn8Jy4j7wv37Je2WZCpWt9ZJJrZrvACDTXsfhZkuQKyl0ceSa9WzPJf3p
I8DptlBdRttYp3hAzrGZo+lqfroLyEiFRbYJyRJmFJsydcb8nzMwroFsfpTleXHy
E/otcnkx7IPO6Yv2UyaRiZPxifMROzuMLDCpWUSW+xkIRW5gH5LcD8A1QnP/JJpT
yaOa/V5ZyPAsV6BZIL1KN+Z8Zm6Di9HuKKskTdNv7+w7a+/792idAYbFSBUBUJYP
yfsuJKsAbDvhWF+z0TICs+78RnEXY/YE12MXDaXx++ttshZLFpOyB+1aOL4yjAXi
2WG72gOfZuw18FgDkVydVEfimwPHI7YUoftuILbv94qMuwfNJdE7s5mQdUUSNzuu
731euB/QktDDSZBZcFpgTIO3v6riF26QbBakM7ELJ5pCUwTLEXau7oY/oxtPqqHQ
/qtDsATPhjQD3Ek5R/7xKFp9H/sF7AzJmjnLY2nzIkpT5CFthzMHl0VhkmUlA8SC
F532byvqoOItRddIX2BSjCSXMqazpVqUhEuwZae04OTyTunc+eL3R4uw8GQmSWmA
VExnIe1nLTxw8R3t6z7BHDggIZrjHMYVRuFBGEoNaUYTbj17v4fpwoY1o5tnYT0u
TnK95I387UgwsLbmI+qVtkCP1axC2Roav/0qPa+nj8BMaHuR/baXcN1ExXEwzZ0Q
tIzdWP4wSfxLLkCoNllLf6kJx7dRAAxzvPZiv1WsabQxmO1yA5Ozb1FAo/qnzeIi
5bttZakKMtWgC/sx5/pGHkWy00KLnbNM7Vf9xyR0fsyYYOg/qNBeZC0T0ioi8Bq/
K9pCz2uZXpFSYAUHEvvpWD34gMMGN4dFtuiPMx73cIe2njZHh34v9dwlgVApDgWg
pp6YrQZGf0kJykzzFCR5BV+KDpSmRmNN21kG49YlscV6Ju/DKhQfccVPmdavHPeK
qC62KmZ2MsH/xkcQ5GIJSQH+F59by9GXl/RX5RHQFwr8o87Yd8vTwHmtfG2X6uJg
lBZtCBf5/XuCH+JLR5snvBYpelqBHMNxMl7OMeYLr/PPhW+oNjSVTX1cyEs6jwc1
HRu6NJukMP+GQG/EYRsSXpoYmSfkDqUL7oBxPt/QI6Pl8q4a1eF5E6M1RKS1f2In
ulbHgMFu5CBZIaRTKwOddG1e+gwVsCLF83lz7HAd4xtz5YAAEdHKPzvexZB3I9Yi
AxLGFv8y0o0LBGkgHXlu1OpDqcLHgjZ8BvBbyHpG5t6TGev443lUTN/vOhGgufqc
kltcXVFT4N7M/YUAB/e9rAUmthO/NgkX72GxmBtBhJzX8JWts9FU/1mdrNr+Kyqp
XzOSLnmYe4zZYJK3iUuohFvGJVXpvGxCZHjH3Wj1LfbyoAbUzt+GHw1rr6DX3YuU
rK52ofm6PTG1ajXp2/X45Prar7Efb5SaT2zcX78DTAgC1gOibVWBWHsJLB+MxPMS
FwDE34M90m6BuV3e2d7qVFFzs3evGwgackGsND8Q1LN6wXEGZMGh9fXpmz5vs/Ca
ubPDzKtuUfWiUQf2XOpPIgj0lWo5NNJCjEIj3LVmgR1qIyqxIVIzfJL2DFjTov9e
Zy5qK4/b5CabEpfl3InGB/GMP4iOkX0XkZXh7/Rd/aHCMzWPKt8HA2+/BNHuLx7B
Dj9d6vl0JZgb/TTngMRwDoQZh3JMCYfHi5NyKaa9GhGBU4GobJjtj8X0ayPOf07d
3+m5xVRSgL2Tt0Hhhyx9jOqAyefk+PcNwyIayavRwszN7rjHOo/95L0CRv2+eaag
cgfUYKh7PZ3h7DhojqhkDbMbGsh+E6hK5gZHUR7Ip3zpBkH/IATzd5t+fRPH5YBF
ZygxOZolVeqGwIPO7ivE/uabP0r4IuOE81kwCRQZCWpPJYbQbSsVAXDwBbTRtiNy
BpNl5BbBzOZcGtKE+/XVJLnwxvio5sVx1qA709S0s7Ol/zL6KGN4a77fz6eyrLt7
iomFSih6HbZV2vxZbIWTauDuj5jtz6WTyKX3Jt96lHrkWSbyzcuwSxq1HC1vSnyg
WF4kRElEmEvYGPlp9qQpXgC9UnTb6JiF0id7oud8Ufw2FXOgt0oiUGACW8XwqeSQ
D4R1r2+wah6HXYCAFsJ41QrdRgNBlS0AQU11kIMm2X5fJxYV2lwdSl1qf7iih6Cq
rw3GVCVEFqscmqKXJ6Ch5vb4l/7Niy7vs+ak1J7pwXzFEQMr/1FYiRoOcoGx7P/z
PJjNftoHCVNWmoiGA+ZMhz5fOoHZi8Zu9os0HYhMgU5URFu8qByOXVOLVFoecIgC
X6nh9DlcBRqyYGfVso4/sodSSZ6YjegFZvqYFJobU7+UR/6gHeqUypcHRUpAuXJe
Lm13wvp01B/E1NNWtijYJ4Q0hGNJo95/PJmK3lsIVfhqrteq77aw6pWiImStgmRU
A8u0ARvT/7+r5ns3x8EdUmGbx+jRKi1Pj61RI2GEIwX9B3WqiWt1ePiy42KYQ6Q2
Viwi5PYK8xcinqPLrpSdk5xFxuVWbranwyDpAk9mSD599Ih4TYQU5uCDg1nL8b7Q
57kZb9ausab1cV81xcqkd1SLhfOXn50gwdQ+/Zu3aJt+kvOiM+8UipH8o3bQs5EV
B3HxleclBrJM7dNmpGOk761HbuqprSTKfAjmsQyha/S8Q6gQYIon3j5g2E9R4zmA
lwbC68fJB+FOsmwEb/5lERcLjYPGOklqWrulEo55PD5x3w7Xt7zXI8iOAhi77s2q
T1wo2+BICic1Y3QEsRzBzXVLzbjUiXn1INzu5liVWuLjWcQgVuhBRDI48YWpsv2m
wSJiBKvHgSgTHFH2fqL0A/s+6G5k0/MCc7SIJMfiCnGU9U/vfvL6Fv8phdN/tmea
tg3wGwIWubZ8aWj56FAO5KTInYMzmPq7JuiGzfYO4PYfwlQR5qU8uI8z/I582FBQ
ZApUQmGVl3BNbAgoOgVenEW8emtZd8JuiqjiqdHcM/rWCH9omOpH+0lXl9jLz6hz
N++vs2HpjGz26X9DQPFV31H7Ex2LiAAeaAE014BrnCHG+unOlyiRlyGLfS2lk0VZ
C+a667BB8vL2I/8AdTaftW8QXHqyE9Bd1xaJDMZbxHdYk8PHfiXaB44mdb1sjZdR
CE/6YPqZpwECWj8XnicJsNZvtxVysKlIUhTaf2gs3MuKwUhQMbYMPEN2FuJp5GU+
ptwNsD/J2NzWKgpLu0GdV2SKNQRB8vnHgI21nAdwdFAUBDbf/eeupBcoALZUBdoM
A7uL8wzA483Bom+TG7SHPZ2ZofHSl3IwZ1E4W8WfRWcWtoKsDsnZEQlgpRJmFUFT
sU+BByZ0RWb/Uok6WwCzNuL0AI2pOb8mQnjCxj6yaXw5JhDFseF2zJj1Rby4cCzK
dOsa0SDdREr3Vba3O0S7RpN1lqLuP9vLYeUYLnJan86/bOT9iYrZQOVq5yccegKK
yM0y1Avq9a+QdMBJ4ypddrAFTYZwTNQdqvf3WipYN8ieq3ww7KMln1fYZhQE8fyO
mQsMPYnh1gOWTj+U6hR6N4Ep64JLLZBL7kgvfcGA/SVi9UkT/6tqOeFcJJBBMw6Q
v7XJrOk/MojduurMrQbfKPqslFU8smY/+wtPXctEeWOdm7hW3/XhFq+qpDAlFQwn
4e0HlTYhQd5HDM8KdbuHjkLE7DAk9kdYswq0AmY/NEaRNnDnmlxM7Harsq6f7LYP
+dDCxc11T03VJoEdCTYHWQ7O6oCn7mDyvDrsD0eJeR7lGJsYHyvsz1FCJvuExXRj
lkqmr4KeA9SVFFZ66Gp4Vaf0dg94qbbvJesSJjzdklDsHVZyjdak5N19Zm/KBiB4
biJWiYUEnn+wPM1JKczU2XBEWcElb9I8XqB0OpNKSy1B5Ga/IQ03OwnV6VAWFkPK
b9IGIme6EOVIpBxhzykBVvmwNnGxmBU7qHSOXjYzBh6fDCTLBf6NZAAktXzvdPh4
j59Y9WCemLy4ZLxVXfFnOFL4RkdPoRaTtq+0c915J6cO7gqqTkOmNgVZD77YaMlS
NYx328fLK6pxIW1fxDTQfkbwQhxcZwOTmDx4Top6czZmxz7GOIx7wGyLOD4N3IDa
JxYppTO0i977B/tJVLz4ZHU+JfLCXP3vDhOZK5zMF4YYd8hMfWxfoejvSl2dpGG0
iQ0AaEW2M/W4NMohx4KwF/IS84FZpo962nn6fyVNFH3wmSereJtV8m3qIwu0JxaK
Yc5mv8l8BSsX5w5O0d7Gp0Dyx4MiALJu5zHeqsomW7ESl5LtHOCHUxFCQOK32Q/m
gSKJ0TteYdaPDkt4AXLVOCwDv4/IRLrdaNhuOuFuJqMUG64QkwmkpOClrA5Azkm+
HN2y7bP9hIhLH5aYv29xztfqzvOQ0jQ6xuDJ8ueMFOA3unCGrQVJe3peYdlZAqJI
HwIEopokHLysMSejT1nq3YT7bMy87g0/cZmqVFNdQ/jHfQtEOOSUwfAi0LGJZujP
tsQ8UyHcUBAXDWv2vzBhegVITTxJ98vbxE9oV2npbFkXgEjGUIaQt2PG1Yx95yt+
TrcEHHVA7do5eJ8Lrlt6CcrqqP0722OJNVk7qVWJdmXWR31QLxN4Vye8Wi7/IHyl
+GP2QYgJJjeFvpVduSAxej1ee8mMH2q5ZoWIxx/42rgTNg/FWuMYiclguogW1/G+
nTf9CzfqHJguqgsogMr9txOiGpK8mc6jBmQJ5/4PS36ylgkbifk/n6yRVPGEO4xk
4x3R5XgNrnQjE8i36qdwZg7GZAOvTg1zUtuQTi90VuIrnVRziHFZk4O1Yzd2WnUr
iyfkhANNFc+mMAdCbH9gGrI3+9/cKn3RzvU0/6HXKghFA7pcYQSw6W3eYWhZw2l5
RMtp+INicpLI54P4cIms6GPkUhVFcHmx4Su0+iz4mbY8IvBO65fuQNJkH/mdG2wB
PwnEG5FTzj/l5cBrHeDLj6/m3cu0BLut+J7xrQCrzokRG3roNhRjm+uO1Ppjfeui
Jrqn15ukK/R6XTi1qRij3eAk0gJ2s99nacRHePOOs9T16nPK8izoULN3CFUJ0Oqk
mq5lBHuNOKxKEyREppPklGfG3enLqNv6/C8jYn5G4EX1GBq7VVdAZIavm09yxZCp
gKXsANtkGPIPAYhpP0x9BHC1UOrZxJdPQMiLbBMkWDItgJrdSjQajcV75lB27SXv
OoHXAVDhLy2ToQepcWEV40lhWF8+6lO7W7FUAKOMbuvmHe1yNJbwlAYUSW7wT/2t
MIX3yvR5VURfVhsRpo/iXvGWm02bBaRO3zmG4G9V4/JHPhJUCn1VU8L2XMQhlEKR
FCvr6U0W8ieSTbtGaJm8noNREqL5h/hEJwLk+nFLkZicTeoPXAWkrIlLjDYsgf2N
ZVMjSo1fEWMDu/fNmoUA69BZZc79PprpJmfrHwypMgmqxgnvyNJ7rC4pvWGhk0Na
msLSvAI4MVpgk+EjsxAWlRPfM7vdEpcJkCzIcENRHSyDkkr+3dhOyIDsG6XTAQEB
oJtukoAUN0eBojVDTJZ5OkBU6JE5N6wFSKCwMfgoi6a4ULDft+2n7ADfmCk0GHXq
IlUOxm156Bdue7JdYTX0SlpF4OLyttlDgdh4/2sC+CysNrPmAnVcQs7ZavQHT/D7
cYAZrDnmzT7M48zm6t68NgHTihmdKzdurepWrDb4nyIPPwq173zL/gfK5E9JBP+f
LltQ9K04Y3wwXxvH9Gm2XuVMtE//72fqzuIo8g1akrVLe19E0VzzhEf3vLaqnKi4
l8JnbSTyemT6US4to2izHP40gOfJT76FCVtFPYVwrmNQN4SufpAcwPTMQNy0my6g
uY+dDb+4iYTOcv+EE99GyEDv7erMC1v9gNEIXU+QR/Dg2up2lSGAlwttR+JALnDF
Xl02QzjMjd7IcKVTDcNgkD+o5ZXevTClFJcgf73SjXCPGgDM9Y4YCmSiuD3szNeu
UQADI0rpkDFij48VsE87U6IivStHI7tlZBdpPTpaXl202Nsy+9n7TbpsTkDzVh9t
PV8diEOCttGxhbMAuxMOMsYo5CLbAvdON2/Qyvq7y/+O4y7S4W5QzSC0xd6CQ/38
BJkqXEwreo1lV1s9ZY3wy1kxVmlXt068Sb2STHwx0XvbCo6ddt3+QJI97a5SBSqj
+Z/Rhob9T25G32mNHMIQ/tY3+TTKE9++uvNP/3kwtW6iGg+F4FpkfTk9OtyziYPT
4NOBRm/n7lEWmUNqLq1qtvE12XPUeFjYobW0k/bg4wIjRV0myK+jopYaK9MCviiC
sArLjy/umZfinvLhROZLy3IQ1y9IiUwSBDO/WC33XVLo6BHZHXS398Dcd+iC9CQL
H+5bMw7Hs5wAgksh48xh+dHVKZSTaZg/mmvkw9C+a1DffKqOoXolfVnhxNU0Xmg8
5be+Ol+YPgTLFaI57hdFNBcSvd54L8lNH22yJ7plFXwChm+KutSLyqgWncLbMJgD
c94lpClLbdC4pJRZN/3B+REHj3IJfHgdMZ2w5PF5dLxkmUook+zr0DTNDWPJdVeP
Os96Xgpnh+CMqUYsYvZbNPwyUb2UzB6RaGZTEazGHJuY2Aeus9kngsqHmkhDKXd3
kh5oKHQADHcsa0eJaJE0AyVBjcXLPkgJPuMfpfkA9wU9S9DLO+V1S/m7h4qSiltZ
S1DkOVmogslabrtWyZpPyiP0Ket9I9DPU2lS6o0Qqziq4w9DW/k9XWdMbWjzIymp
D2oegDzqLcrGaz0TP4YcOr73yg1KIM659agtZRfMpwz/LOtRlqhojNJWda0R3ubP
TK3h7/SIU5J+EXGK3GUlidX2qM6heXCWZRopJojXYn5esauZ48PvBnecrDbsw6Hl
Z/JbN++ABDtLsM/oh73brQUhtax1dOx01cbMhJG/eogTIXLNzPtkOb5Ljjcl+i6k
i8eLOIJIl6L68RXFMCkBNPK4fY+3Ob+clW13pEDD3krjJBRArxzbUU+dwcLC+UGz
YFrBJeTBCgmmBxCZCPY+pgqCUnpnFUbydBfAk5J88uXVcoj3tdfNe6xzmnoQk5xv
LdWmj1qXr2kA9wbdJS9JCmFZNHr8rZXAgWr7WeDEedRXDI3pTdSY+gLbzDSCJKnY
dflSQQSgui+8VDwPujDgiPIBho7v/XPyQkIvhajgRgeqe8BykFMCfm1g4UKLLctw
Gv0B3rdILVXj8Wd3Mlsf3EFkj6SI7mZPHoGgplIweFsq46iB58wGI3/frVgsZZFe
547mOAoY05Z8Wuk94rJeNB6UH8oo8nNQLWe0wd693NZHBG5pftyupPF5nToR1Rn7
3F0X3VojPzO29F9COFH3dTqzuCNcI1QTh0FUcP3fMWX1aFywJYCPIYtVIzniZy46
FxAZ22DV2iNV4jXdm6nOaGJTRg8yN5IA1cDy6Dm1RH9m0JTg6zcMGxpR+3FYVxT+
agCKrV+sfphzhzZVAIpHDds1SM77oMSCEzH+lk0pXdQe+6OUlhUh4HBFis5z3Uez
Jwr8tUp/VbfwsAYy4dE5v1McXt6Vq6h1yIRlBCa69S6DiCWL+RHiyjwhYdy3+ete
8GaFIAiYFT1XX8zEC0cOGrjl0Y7G6CtjTUAsjHrRN1wWTylTjrDgtp4i90cKxO02
w2a8eJ7OB//LR1OAvGgpKqrTMZlaenYzjFSqEeg+YoitaZhSQmy5YQX1QpBVXwrm
nwEaWW9X2dBrIlIWEa6JtxfVH6glt8ZfslVTwlUQM4zS5/hQSqSt9FBrwZ0rTtaI
aQ1sf5bhW+V1LNO5SJsWu2VAUDOy269piUDXV99wDdT57gaULIsMZUOAWr2TyHhr
/ftwztzP3zb9dSFt0YJJJyU4pLQT3YV+PHln7XzCjI1yV6eID7fSkiuCJy8AioPf
/YUifx6+uDlD5apJ6KUJniBTvRArfuhTZA83eOQ0E5Ny/2OtoQoQQsSoGRvuzqvZ
wj5rDhSmtJixNT7TTw8ibLYPknYRY1LkkCE7wGfD5uifJkRUl1WO8bffD6JVxihW
kOaBDD8X5KlonyVeG0IPFWg+TLgfXqv4npKD3oLgx7FHTYzDKXNhcPh1tyV36TCa
e1uIcTB3DsXf2zFrciLW9QVNTZrABLiG2CqRKXHhzlQdovmZUf+imlFuqRZsoo0n
4wWvg8oHfQ7wi0g2oGzS/tOje4tuo4byYaVVwtkwPNISgPJQY4CZlZw5YTeKjhWT
dpHdd8q2yFikcOHZ/AAHKCQtsaVhlihDDYbG6juNzcXQGUCDfIN5n5TbCLUlia93
fvCnmY0IczQ/tAp/DCqkr4G/zO8ctUTSr8nzIB/CPtu/niXWwQlrIzc5OzDBdWLG
6qZeqir8klAm909CmSTHW5wF5OwndKHq41mJqghsZlAULmnaKBPIAawBNcQM3oWU
IYZcD/imMnG3xew5QiSS+heoGKwlX0gg0W+zr3r5rQEe9C7/12jDqar/WxSoVMB6
oMbx+ffVI5Dp4lpPE3nkfY7/up/wYCJn293UbX7WyJI1ussUguiiqnVkALQoVTtM
CerV4nX7nrBIiKKWamQjxn4Tj48n/LZURP9nZZKVUOOyy+oU3IUTeCwJUGpMSb/i
riI+oedjSQhIV3gWZZQeadtQBR5A2adwLBL3WpUiEvFPmM9OhwRXajyCoO4o8tUL
mM5CF6EP9yzj0u3dvubkbVERDtVoSBTNdZpzpAP3P+FwuP/dpE8Xom/wzzdpHDYi
cen3SluuR/I5G4hGgO0Rts1ZmLzM+zQTo2+lK0gyC6Pex+CJd5Av5MniQKqN01wB
UzwZLtfSzW8haRK08n/ecIlvpgv/cVDQ9w7i2qtVTib3o/CtnRjsfHtC/eqL085g
01tk0KLiRu/P5s9RazT7FvijUCQvkPOGIgJc9mMkzgwWiMo+bQmZfHVR/VNy6wHA
pX2SL/8SNQozl8CLI/VZRvr1ZTjlbdtB1rqFyT/frO6cxCGRnkgiLdR8v83ZnlNX
PHWkYujDL0TOpfMn8iy/gQzFwnx0M/qUXEoE4u5QOuy+E1GOastzQRtkr7yk2SR2
2NhbgI3Im7dAxDg5d7UrYSmSMmK+Xe7VfPOgG5gJk0GPZwpUSTDNMJqcrym4N16N
iT1iZzfZELxG7Dl/+rW5H0F/K4xk4x6m5VNy632DUohlbFXsI1qBm5ewxZ66yPbX
RaB9WAZnXi8Zt+QEDE3Kp/+nTuKn8TdzRm/NbW7G3+u485kLSXgpkDTKoMRbGJ0l
DWD8iOxA3XLvPIvbMmOr3Ybvu7grZhU7EqGstAguxm5qfuhGizTTkh0WLhwde0od
Mwsv2KZY/2Zaq31c4NBaeGIjLpb3pCgjzig6ue0aIRyMdhdDVMVFk8cHxjtzN9mG
xJEvkg3jU9ugn6omqMkD4eR6E3RDWAPz0hSowmRiy5F5ojtvcSMALT5J7BP/28gs
46sTavPOo6/Lsth5bAgTC1iREylYSmigiy4Xb/ePS5JaNb4VGo76W+YcpnmJ/ha+
jKl7wse5t2aMS1y/t+D9F93SMqsy2o9PI2Qyp8gzpDVvz5LnaZzvNEHv2YY1Lj93
gE9tiEivdhqWFhwfNHMvRGfW7Bk98FmOe6DEi/T+urGAoEoTmnTF9OWLBWgyuZ9B
C6AHJCb4Q2d16y5U0ARFOEd82/6S/n7jEqJy75qF6sW+agKQ/4d2JNyMT5TQaXN8
OGg27gGwrx+fnMobh+G7jclAJR/ioBC4DNejlVfHEIvwV3+stvKqA7oWaF8eJbyd
VdsC7OQoRAmQzpiRpxcbTKndtYAA1NfeJiQnlJ2rXhM9AXruI0mKam/XWkqa/fzr
lbFxhnVN8ycl0r1mXD0KViGLsq6LJfJzJGe6aWDpdFcEmcpHvTH/Nlto0ulKIpbL
6yFnv5WR+LlB7o2nh0IcqrvpBkT5PfKApw/vqomSGRGfwbpN233amgbsLiApYLys
Kk8lMKl/Esb6E35sqOtA4zB3XwikZ+TQFCsF90EgpMSMN+POJoDvzgOpcaudjJmt
jqNpFCgTGSdPBn5L2IZ+4+EmT3OTXDa0kHMSqjlyRR+Uc4wOTt3Ii5K7L4SKJ9sl
tPDX9E5/v2RF2JwQ1/fX6QwnfIB2NQH9QM5iqABa9A3zScmsdxA+bvcGK7ydp0Gz
fGnGckCnlT58RfMirPo+aWHzaPjW1E2UI+aUTYqXcfK7f6N2RbMtBJsPmR3e/+NL
KTziISw4cYJqvg7CElcvZWlt972qwlXBA1mqU1cwAhWz6HA5+nULfwZTL8y8LzFO
qhIwU9CQEeZgEg+YKLAb2F7CxCu0e3KAus8CIVjaN1Rd+A/VplCJ4o51Qqy0BdLp
tcCyYL3md83hWRwheU/gDV8lkWsw5mhDR+O3/S9NhSCmirQZryIg613uBxpFm/u6
EcaXBHidqp1FuP0/VP0uRnVAsceDyyrgeFKwt/mdVo16abcYJGFr8j14ZW2bqtIW
tbaZZVaKc7kYUG4UE8C/fX58KGWrviGp0UUbBtXX6yq+iZiuN/d4mKqaJ4mXHdBx
qCoasHRsK7m6d5G0exncLk1iCgnapj1kO8Z2CKIRIhSHWyDcCVV0l9aOMVa04yL0
pXImTjloBN6VE5yYOc2binji3LVXxOYKBxG9OzTo7pBzmfk1f1NCTEJ/QAQfqRnb
k8isjp5/q0NJUqz2mWLk4I4i2kthDswMTpoA7fJJnLs11hPYI9JgjfdOHgMXtD5T
f8SUASmWK02/gD5PfFeS9imWa9nAEdbtEoiUjuJ9T1iNWDo8+73zJ5LvS5tlJovp
qSUToRtwWK+L0B4p/z/fTpksF+CxKhC0DX+3ZfK+WacnNUoRucuc29yOBQftmtKJ
eJX0GMKHQGRNDQw4lP/Q1p0f33JE3IHMrJc6AT08OTPrUD81U5Qq/6ShHXIsR3pj
D0r5axeV7nkKJ8z0983BjO+ZI1GrFXNgEZUzcDJM973CyMZEtS7IfX6kn4pQWafL
QmlG1VWYvbrelkFn1iBnt2lNvnm6ZlDO4iDGr45THBL10XTVla/UC7dHhgAl3O07
lXCbgxafaJzxg18elhhScIUuNNKM4fawDCBkSpqxyPs7Lsu7l8xXc50gjCAo3lBm
RfsisQ71BSuBJ5x044c/+fatiNsc/KPPzun6a7wTDZrnuWKeZjvwA0/zVw/HUbVX
ARl3RxUJSQokXWOxiX1xx8I3eqyOxts+qXRpyn3clyeD7fMW8cESWe8GJcCRJR5f
cnoi844J5Ocq2omlkFpzXiacY6KI4KdZXQV3lGaeXjLwdqPTGkw4pXALTgZmOW7f
qt7ScQQUA75/TCum3BzEPI3ha15BDBnW8DOY+AN+yu1Tlro6ERmw1Be+318d7IFo
wZnEJmdhoU4Zu67QlXL+f00QRmfdDS3+55iPrAHNwlzCfIeRQmz+PI0MqlIdNOW7
TrnupZzykiKI0lxESBP96Duj1nAPaCjjWg6Tx5DpENvj6l9gZ9SrwfkyFT+0R4tx
KU/X8R0ZHh9gJu/MYnomsLVOFv3R9nTEScnqxFGNe3bMd/PKoLynp2OrBPvmudyZ
KfJwP1kqAqh4MNoL3aM+uGAQHsVYNEvm0PbGLRg/85DgiLdC0e4if2gIWUvusMHm
UOYwUHCgaT0VsgYdQFGhhK4PeLPQJ3EEUR2l+vDPfTN6Q9q8XufnB77i3cvM0nXT
W+MTnm3zJ2guP57q2yrPMpo+NnAwVIL6YuHuCHPNgqYWF+HtV9PapRjd8WMJ14R3
AlSjkoXHNXGWPU1Q1L2Z4DRlBZ76rvjEA9nNlOq8TXjkhMKGmm8CeaEWfV0KAGvm
7tiMYZl3m0AsQkj39zs7vCnAVJKbrqgzUAZbVCAw1LTliM1nPgLHzoD9VM7TWTBZ
ZEsOqoFSiRn6HP5aD7lTKLX2IQQ7f5dgVRHLme8sCy371EW9yFdT4+zga8gWO+Ua
kWusHD815B22lQYmNCud2DMzb+yBsn2XDW4YYve2oQfVpnbXga7GSRV8PDz18g/3
CVUwGBAuyPvZeTG8IGrAQGztiPFDgSkFHUv6nHXDBTZAunmpUuy1FR8N/f9gGl7f
6CfLQUobzA0WiB7zY2HajzM3mhCMcormDo60dcfaW7BlL7fdIJdh/RU80VvkC6Yf
QgfK4m52rUS0G74mfbueWJhceG0KEWZfVF1twJWFD3yqMQpbOW+c06/e+kluSUC9
+lYQXpObZgc83xlkfIb7rNSdfEana9gLeVqN3SHmqzQrmIv+p4tnTVoers7CmSB0
QutaoHCl8QFYW3c+3k2qZ+NlGOIKCFq4EfSm0iKN0YfJoYi3Mu/g6soF0XrCklTP
VASn8BNr/HHzxMCGMkJ9ePZKOQQjl8oGCOsoDufTFL4m62NsldnnEIbWGN9of6/9
ux3iqSFP3uLdFRVBOkhyxgWe8Rh2MTl5lBJ6zQ5B6gKnVB+vzHMA2A8no2drbwrs
rVAU/UM1qRlyG+nUidwoFzETDquLEm8kXXK0kKPFTVvzqn9TatNtRwam1cA/7jBe
AqjAJQJsoWEhNVD9qByyLsmFhgPIHiYCzBFw+jm4vWrmyik60C6gLqSGeW6XIpG3
3Dob/azT6d6p3z4XsCOFYs1GG+IC796c7e2wCJ/+Tr8XjvEzNHUXVBF62Vufv8IH
8mryMryryfcCrsMSIBa1Xyd1LqQ4iBLuqnk/bify3mRq3CSP1J9JOdEDQ6otIJ3k
C0MJoRx/eLDXkPcmBuIb+lX+SYhQtAb4/z+tyxu6oX7JYwIq8mWvNdpH8ZsKILri
V3BNCO3WTjoNwyVTIkgagW0BDPiQFA3wtNUayyXeH5qCEY4RCnxMTvuRC+w8M5YA
T/P7p3euMiSgN3vaBOhYkd+D+R3arKxQTW20P3KCky4N4PlLnIAYg+v9dy/Nm+OC
BqN3bTZq62s86NR+mDwAvuNySKdpZ5ajSolrz/ONXrspoQhwbrZUhdyS2sQrshYp
fym0uQ4ypuXtiRuGdMWhiNa0qJ/l9A3n58DBgEa14XLQxpz5tlvjsYzNL/1IFh5z
fgJIsNXtJx6gW6hd+qs1bp3NAwZWs1dzqYkiyFCLyoMNL7VONJkneCadMbF70/rr
KtbhTOMETpttvzSPlbw8jqYpF9gVQOOPPrGXuAWRbKiOqiZKFWHOZbB/z4GZ7DyD
0ZhEDLI9JpLhB7STKcfIfXwRNZ/CU0xRwNqYnO87liAo7MFDVJMroLTbMD9mRBkV
bbbwFKmpSH0nD7th0KL4EI8qbJ9qM1uGItZEo81QmcXQzTWCWapDt1wKxrEVZ5gP
z9vzjsgdMHpySkUrt9x8tiUzC3VTw+B7YTj+xMuI6XOlNsHOCRG4+tpY9sB2xuVO
P+JZdbNDBJvZhWa7joNFJE42KiDQL1/KA4VIBmJGSr1X4uJNBJlNeyUNPon/4dGA
bil4StEQl/SZQVRoWKrOuFhtFAxWozIIc9CVrvOvcwu701RomBjaY0F7WlRYxW4m
qiRjziuyxnRlW6iRV6JgmnPVFO9wXI28nDIt1wJ7lHdg9fqMoYtiVFk/j4dZkeWB
CmaUWwhpvVUoeDCNNFIda956VfhsZTrlPYdjQ5jTm6XdnUbG/xcwH4N2in6fSea0
zSwJNufScr0J9BSK2r9QM86sefiWXNlFkMBEgk6kWgJiAItoICEiKD2l//94rnRV
NvMbv7COqU+g1DqiNK7rSsuvdG+kBouyxGpD5qp/qIEypRpvrNEEdIWVfTkdBaF0
ix2ggsy0cqSfk1tGgyQJqiEGvBZnksnMEjFy1QBqFmHgV+z8flPH3L8/qdQX6DLq
paazwahVbhyUcVSz76Y+dmLHha6smPQwPfr4UoW7uwdWUxSNcmGc0K7s3dUqRCBf
GBF9/l23DU6zjT+QqdK9PfffK66RwojxbR4ANRMHLf/hPxQh4U6S8uV1Za38Irwd
0tOwUgPuTXCXq86PwvTFVKT8bKO1zpz3emjUzyA/XFhNaDmLAM41PkrZoQFsQ5f9
Api/qqbyn7gs0wYFAzTBVKegvXeGeM40dw5bKvAsjZ9w6/1/OKH43eXjAU6NfASn
GmcaGyU+OP5CWC2uI378YqXKLXePm5UwG3GBaCqj6AH+1FRPSo4kANigTBVcERvR
l3DRLkT8ILNTUnwLVOsH3J/yB1fJzw/rsNemCNQYLMGB5/frN2ZAcsIQYgvm9ymP
1XsyjJ4oeX5qmA58pkle90KY+ZZRkcogHCTxsMhYfUjdE6C2vySFqaT5NnHajYfY
ybsIiEEbNCmoIrFVvXBseGX4hM8u1KeH7PrcVeptLeADS4aaZe3hVRpJtztbuCjK
6agL+QiOUFGwZT8m2WmmIVHVQJY1i3WuGPg5IuLgnKyU08h5wY4HH95/NSl7fcx8
RWmADUSEliMuB5lVPHS9SkJwjC4kvwMh0dC6J4PCx/C6PeppwLC0TQSrDn8k4zgh
ZCFklme3PSOQmVEK4ORMS/t00a2qih4Sjq07DuK3oMO6u36jh5ccM+iC0KJ5F8Y1
mzgrDVfQ+wOEuMHxOJuBKtVdo2HAZy6EFieLzMiJ8p3TkuuCiQATb8WsnjHhI8ET
h2mHv2iqY4fQW0B//657J/dDmyN0brsxdWCOTsq7QO8CnWkgMEi7tgo13z8HTXpG
Cuph6xOyxIog0JQXN+d7hyHIuZbKpvzekDIRrtmyoSCw4wYrQCg22abcmrGyRqHx
zmRCIFaUoSLC4D6FfjzLjIovLb0hs/CK5d62HwdpTKH88H6j7Dc/L74ylTl+/0Hg
rVO4ADL3dJCOIQPtbh9A9fJzH1RUHAJ+Bl+4dMxhu1RTgAUniVgEOKDqDKp1+UEF
9YBarYMZu7RRedhYGyqO98WK6VM+l/4bm/lUpl+/pcm4uSZWQL7wJpQ6pbT+LvW6
EpxicezqqQuTig9Kkx58U6HsJ5wi1lgTgg84nFVtu6FyXu6oz+eLcjh1kjwrTjj2
pFlk02GfWsjQ8wcywS+sKFfW1jSV5ePM3bA49KiMVoM2aqGVSKER/KZfyl7U6uYK
yAsmAOmoJYSaynthHMQ0XE8i+x+qZ+ceofJydVkRHzaw2797I05VsH4lCDcDdJQT
+Sgqjxhkjq7p5NRCg6ageTsOsQ3p9MndahDBgUdwL/9ui7BTjZrqHchpCFxkdCWJ
He6ICxVerRDEO2rCh/MYvtJtWTUA8H5rIg8t3axofzgNJ/k056rp9aOS/JCzzSkW
YEMtMEDXWFpln7WJcqiJgYYLShb+uLo5+eoFIWFCDzrQ0ivatydm22PeLge2q3dj
HuS+XxaEAHLnz/262+Vxo9XW+sZuNzffeWJfxoTKXlZKbYZHTm1QMqkqwZhmLIn6
JKzPw0fQq5qUtzAQIYwZKNTX0VoRcHtnXxxMzgKnQYXHOEyQGDGeifxk3u3RlY93
A2XY6ygRdklvcD/6yyo3qpsxsi8w4+gcPr8HbEoISbROph0Q6OhQkgTO8rKflXoa
yydaG4f63aBCaXjXR/r79LDM06rYDkrt7ighvly5URxRyzUKLQuu3fqas77KSKWG
89mA0JdktmBk4Hu5LTqDaK2khkF/7TOwXbrHfDpq5U3t9jaXvHMRT/7ln3ebMIQj
hTBK9i0yLde7BoH128s0+PO4S0WWWAdAPeDg72fDCPBjSrcCq2QWFhry/s8wkzU+
Sb2bryaEW6xzPqY+XvM7xQ3SGG0rWT4Kwo7G9Z/lOrymMogUcl720jdVcTIoBS74
Gfeqxt0EaEADAcDRVhcFeIf0TXGXgafMNXQ+Sr/JOBGiR2w/koAwcEVm2NII/ayO
t+X7wP+JmldxJU82epY2kfi6FEXkdvlFVrecSiwxG3z4JctMhx2ynVrB+BHpxgtr
FiKDtrrOpi6p+QvDsGQXT+TWdniflY1ehvPmAof8sgju0vwCR6+2q6wg9bc7tP31
dEdhA6uYQ+pGqU2swZVNUAYfNJMYhVDgOKQvrv4fhjPuwBlww4kkvmoUpCDXF6+a
Xxniu0YeQwHnfOaVDfX/iADTDycV2ZrvC55XhzdOBo+4DVJqyGjHe1N9gPoN65Pf
Yt8Un/UfEPAY/6lJQ0S79XbeoUGSfJiL8QHiz1GuujSXKUgvvXiNKaZ7ILfMzqVH
gBEJPpa4KmDeCzTLDpF48rMMvMrQOUQ/Jev87o88HMedckXoaCU0Qt8ro3Jbo7rQ
7FwRroizV2a3BzVAagt6tCl+gMRpLZdKTgKOqAZLHGswrBYTMA2vgyhFmdM6wrmt
bfUCqpSCZCEjKmNXVIl7v+EQUE4kFk4c5E8Mba9+UA2a5brwV2ba0mnL3OV/uCM6
UoCi15D7j997QXGB757jjRTUP0Ql+6fHDkGGap3PKmOsACGbVHCRGt8SOisdjJEQ
CqyxFyP+5YmVEs0meGXsGetvugdlw32r+Shntnug2EnKanRnYtnbpq2pRdzo83NU
XYYuO81JrzPKDpaI1tqj5yighMZetrEq7EZI6mUXaU4dwQaXy1QaDZfvQEnjRxoq
0SZ6/2/qvUdL4J6elBDI/KkTNcpKhhSEKXjgk9BGkjIGepH8seZgxMvLiDERzowK
UcuNchZv8pMRe+u0LUn25G2yCMuph1Lqo/oI71fgcPHgzLFKZsYsvNYWCDXzD7RT
W/UCnztFs8Ssv+2kzxxONWqZdfTVLZYTQI6eYdoyBIG3Rq7a+702Xm0wH/5c1Ari
s4C4qFMeTIYwvh1VPu+qYYdbY0ZvT7SOFV+RSf70f9ky7/YGzfUXbgZQmk3aftKu
U+ueOZQWEKOuKS1+oCeR7tB2OSfkNBrSqlEt3DP/IsjMCIpqg+iwlC9r/8sWDo9q
G6I/48T9cAZqM4syv4IxsTwfUqMIf2r4bk6pHNgP4sC7YhHeYzSIvOVmBNg3LgWe
EX7deSm99q4cQiNsrPszmwq00NHy7xTfuYew34+AHB9M63aqRvtrNVmxhIeXhFjb
jZOwUTQ+gOF/9N5b59ej63IM6LykXgzPOvUkUSTViEhBPprMaWmeum5vuSdxBoRg
E2FtkHaTxeuzbi5rIGYYW4uhbwHMOjPWxzr2/bkurhY+/L0ri2HW6kh79nVQOVZ7
qWHy1KNOUrRmokSWlXfW5HxzBpwcd3Ey0oyaAjI5I/2hw+wnJ2IOd8bzCBtNs/Rv
WNW/txtr8j4Vrc3vnlae6VjkP6AG8jYg40lrX4tAkgONJ13e7BnkHleSypeWWgP8
mzQZd/3SBfnH7s+I8IESj3K4wO0KsNeTmKrE8NyPQ2kjpAQ7sObALvmXtzxrBXjx
BQHJoz+tflzeLh+g8UsyC64AfzJ94DcfVl0YDbCNiLXqFdioT6f9jx2vr50TYEyo
C/9wXfj6rLboKMK8vs69VBbTN9tOPv0Kp6M8crImVvMkncgxqH4PKBJhCUJFFAPh
ee07pMP1McKynI9r9ekOSMechcmskWUTYfo/GJsLolIoEZ3HEAoI5hdbpG8KoWeZ
mBrlTs7MzmQbHucUer9tlrGQbCGgRYxPDMwstmM6NLT09rf6GG1LbYdVNNkN3B5z
BStOABAI2cFyNpxSLvPo7+elqQr1MD5cOyMK/rdTXXfvdhgHpqS1ZEGtG//JdhHr
5C3k/pHip+ra7Y0tfoo4LS5AEO33hx9/Nz6exWxKjcWPWScZ2HwWNtGqNykz+Tu7
qSjoLdQQAtKN/tw3YCmkNkphPERvD7Qo36QZi49qAHGgNB4vDp/LhnkIbl45VLYK
1C7YAbXR6IHKfCYTr+xOuBrTvFLa5aEJD2pRqf+FK0wuzNLJvNXdvvy6TlxkIFag
0d8joOjP9o2SguR7O/Boooektj3re2q/pW1J42li4MNmQqatpYPDCNdpzTgQYdHV
Pd1ZsMZcM5RlD2gE0V2qeG9TKV/gYHoDYwxu7Q/UyP4jVSyCh3HNgCkB/7EZ6EnL
1n5NeI+SppKB8jKhmjZmnFJavdsixrvdy2oa6L++N1H6K6/ezOkYMDncHj7tdB1X
+R7iM83gwOeHuJJrT/b2WL4xtEYqVVraXzFPiXEuJn/QmrDpGXi8uMXsLGZA4fdn
jlJH+pb1GScv4i9MBDbspHF5gEO9QuWEGIj7lRYAy6CFjtkuolbkcxM7iNoy/IE9
cEX1pL6FUkSgiOxHzyaSvL6HNaxdWG1H5pisC40qtAw4QQt2kz5MXyKRIRtAcnhq
0nhSuzE/cIZ5O8YA6xMERmzmm5uALmcPX/BQhV1PI17AY04COGcUHUIUVl8nRtAL
0LGkJbsVDi12e9YSqegxW9efXwmjCurcFDe1DYWez8bgPMGpxSqrvhonVq7WhAOW
+YcNAIi4ZJfFyHi6KJBFnpIUt45Ggw7DmFAgIVz+aRLEuTXkApGQd/uaUnkymMPf
4b3fZkT1WoQ9zQfiGFahz3B55wTPHxKVjhGMJlA7CM1UlyoGo+i1+mh0aqwgM+8j
b6Mnfc5XhN/86CI8Yd+QKV46QfCl3xraKqoM+kDApsYtt2wqi6411TvZbsTs9mDn
7dgd2+YqVWXVC3iZdbaqaP8A91ox324vtUSETLRYw/yTxP8UUpHDnETBJgdyc9AE
REBMKfLE5JeDv3nl6SUCtVJrl7jvJQu+3ocUNwixx4XBDJ3dqpgkRdzEMr4ueBn2
jU2IOY0ePmsil0IYu1GoR5oqJzgTqx2p1SedOTlkMpkEGxqfQblecflJ4rmb2mZK
Es3xeKnHZ5emacD0NPE4cJwI5DsQBJrFnZyEBOLBpwx5p5GgxJv9cqfPQImMVzy4
JzayuEFcBSE22oUZYbQM90ypZpxxTet/l+dycJF+vE/1q9U0D4xyuoS3IvB7T+Yr
H1F/2QdbBE7XyBabcublmFPZe+uW/RKmZBpKNa2E2As7liMKj6ZlGbu/+eSeY4X7
UG88cks24GhXSkeC05uX0mC2JODKJjUjOOURLMM8+zr9CjQcFS5aTAGnqF71l9gm
lVdrpWE2aFLjVbODjD28lhuTRQfDBSYsgTqqnZgk2cosRpUJLc7Z93ozCW2gNaSr
EUMQTZML6FfjRUrI1VE0iFcue+HYMepgDVYPrdlsSNT/HRrY6uFspudd8QL24idX
TzrSUvIT/7OUuPepYkPKDYwyIaUt6uj8RerTLIx8e1JyuWpYOfUqF/yV3fzxHx7H
bU7fYvQrx10NK3Yat4b8W1PH3xhCi7i+y98D7NGLFI20vjwpd3CClx+3ux5924w8
7D7Ge57EGvgdW1vYmv4Lu5G35LCoaPxqVNC+CRyfC8z71RD3gm6+m/li1PjGUb41
co1r7hWlxA4UIRdgfMHpvrUP1SJBTSTr1CX00xSgScX0rfP5ti9+0/PBJGTL0Noi
B02FDJ1ZwAYdz7kYpkjyBP8AhXv48iQQam76gwOAI78bcfcW7VNRTZQHBvKpg5Ql
95woFYmtUx4wsXUGWkmTDfcB0k+KSByYKQLeGJLlo/DJpAP7ZoD7qduOMU4fRuuF
cb64F6uoZAfMUBSbvtAqZcoFdzLq9zNS6KkipkMgHDT3pBsh3D70FyxYs3r84nSu
dtfJU/Ij+zGM4RiOstTFFkJj0MhwVu/CVFnGSFBaYIVcmT0dCGfNWwPNHxGFaMbk
u4OB1D8dUgEz7cLF5XxEHt0JmYkOzHp0+T2O58wef2w3xvm6Pz0PPqvy9ZtI2jE+
wkJbb4uH0os0TPvYwATA6TvermaSQTkt4qsl/aO1pQVk9Wl2h3Sk2EvIfb6tH8gH
As9vXzQlZbUGopFY6iPUWe/CK/LAOLMvS9y6Pf57qEqvNFyfcDyC9py2uudqFTvF
gryhsd/IfnDNYu0ZqKKY32i+8aIERVcgxxBSTLIndYW4DAeiTEDN9dEeyrfoPDY0
FUCjFaGYIO7VDmfAjypkufJl+1DfxhnOyXaW+ZjqWvQxumD01PT+cKlZrnb/y1f8
6clpbyP/6T1+l6oC8tTZ3UQ8vlu5Q2XZcg4PulZFXRzfq6vIkm9SEkskq0XpbfED
cMXf3MhOnguNzOnVCLA9LvwDiK3N/hcTopFAdjkWEXNjB1HIwMxrmN8XW1eKVGoh
A+PwxXH2GZCF6/8qMu/CgbNKu2j44p/IXxcPkHoyYskFfnB6CuzRyc0ZtBG61jS7
Xr9/78BFoLAm7j/0tfkK5t8fVjVz9/rjso8fgnJSPI03lT7iDVfNUwGdrYJPwfzX
EKBC2EFZR7mVyMKgnDoLdBujljFNN/L+jf9tze0bZYDQJQT34KM/rre5x+b4XgKg
LvIbUpUDo5qM3GHXQt2WpcCCNnR3at88pktOsRYFOM8sE7MT2Mri9oWO2Qn69urF
X5/5oDZ8MxMxe5HZ3hXYN5Vtjl5PO0x+H1qhoGR2w9bq/8pDqasQWUMjsL15GGl6
sDHr6fyr7YlYDCkyavyUbaAwQWCO4TsYbxwJRkmLcZ7hHsrUAEQ6N+ZOCfEqtJ5O
vLDStnTMvW3LoceY7aw5nsFrAU11vJiS0wjVu24Wg6B25nspkR0/iWEqcLHesqud
5GAIkqz/UBgB7wBUbWupu5jHm5Ni0dtA/xbEH2VPhYw5oI58IsY0TxkS9cvA8svW
2Xh6SK6MUHdjtmIZHLkXVI9s8sUevX0P+6sNMRUnBpeR82bezNd3w+QDvwva5aO5
hPqfOMFJmtKri9q4XyQPsmN8mYwMRkb2JfGBKXUQO8bdPOkg4ptu8gbv6tkt2OsT
3PZL+PVDfJpZb4qq93UgD+6O3dtO+3Tqg29wo+39JBgxGk0pfqIEjufj2D7/dtWK
DXAKk5jBI1+MQ6hdpWiql5wrfUHB6xClmIHGcRdqd8Hhu+du1z0cjXadSFpdXWqr
ejVKuZwOEwIze/Qd22jsFBG+gDWV3ADtUTpWuKsZf8Gr1YbVjctpFkILu+QtOzCg
iNZBJtvyRKQZFxuQgdtnGHs2k5QWNjBPVW06lAcYtt7M933DYmzM9q+XNYLqnefp
c+XDTYNWUse32VUZ3nqncXVt1Iz2W4h/wqB/dtk2n1rG7WKfTTj00bNm/Wj6uK0M
eR3M4qdoikRbqVDWSSdFlAeziION69UJB8SKxl1DDMljKY+8w3Zk/vsiiVfT6pTR
FrmcQEotRX1ZHw6RXxaJFCdoBveRcSx8oElPTKbDPKUioIvT+aPEOoQU7zrVxfnk
ISZn5AFjr6iWp0TwUWkD2mHcKNMtROYf0cNpaaRaUofFr9jPuvbdMzz4QDrk3kv9
Yl0iuZdRK9jFXS6yTzQTuoiprmXCws+lEP6rhlSgx+TS2DldVR5Lg995knHDHclQ
w1M8tqtc+qjSWa4VV6lr/vo6nw3txXPpMf99pz9lw1bG9icaLEDbaj6Ho9aKH4dF
+j0UQU/QTlX5tlSyrq9XKqnKvFwJX9orwmj0mXRWFTbwGLybDETtpK4+kIvz1A7K
tyfe9r79vKkWNcquXhG/iB0/4DYThT2PEYzXoHlFGszb5NzAnJhWPGJNZ5B3UYwv
cdc9YjhSzzxM5c1O9zSL53boLVIKjopVoNEye6cTx0Vwvny7wfRRvjiHmpR/VvgQ
+alCnwevF+iMBS7jeF0ZB8U17qZ55xzIqetmFfIXiu2JqcATjqYOZFvw8gPHDvYc
EouvcaGjWmKwFCRQFAd4YAWUctaVBUb1LZjAyjy/UGny5VWKAloRVY+hIBfoOTxf
V6+9tzBnT5rdM+tQ1XTyP/+keTuFCnpYAuVnj0r2zvyXtRYs9DWyluE84CgtCSwZ
Yoy9c2T7uagPKlCAVu+b2LpbZyM1VQtd3VKIQyP9Zqn3I6C1QrP+UXRE8z1uKF39
XwUK6IANJOT0crLUFO45Qn66S1y7AZlKVopYr6mmibtEn1h4QiG47AuwroFlYe04
oEkeMKMm3UCskiOfESo/6kRfvAqFLrnFuMzBSXrfqZAzQK0j9jHbYT549SsJcZnv
Rba3ToaO7oSTDYpXMC3KcqeaUxH+QN1iN9BZR4URgF+Er8uLStsp6sKuCA/X89S2
TW/P4cFiEhiEDpQwdp1tl17tY3cdb0D6FfIVLFQ6nNY5pZIx3N0B/Hxqn8bI+Y+8
6FFxHUXwOFzj126bXRmS2Br1iqPgd2y2VWKPUX335G2iLaMs6Fzp7Sn7UGYXiayS
bqz61W9HB5kik6nZP/i6SG0Qv0UbDukmYcOYrKDDtHWOl3oNqy7liiSIULFRR+/B
2dKPyxuWcRiCrSAVVHgjCUiM8KqOjWdqXFg1t4dWBa2P7v2n6kzkygFI81XLOjlE
voc60fxCBRJgBBmQ2rLWoOWoA+gRwQmEfGFK9PvYoll/L4JNCiNsILaXzojeKpnV
ZctUiYbhwb8T1KS2LmW+oys/1BZwSTzYbiYVcG99JqZ47tjoJkNUp3MIdsM81flm
EH2mVn+QG1xmitiksMHL/ffa6vsvtIeWUT7rOKfrwzggjgG+/+gtJFWRdO/6eCIE
yZVjDx8ntc7S3e5/sRNXwdZOrtYGcR2b00KE9+3KLE8KXiIiyeTF7ArALW9w9o0L
p8GkWiBol3RCAlxsNX9/gbV63GmhbghN6xNbxQolxcvga8IICBpmZTSloUVonQ0G
J4UPqY3J2RMzMxwGNXG00V/1LqVMKPlzQy5ifHfzi0dOcse0IFYLfVGlLLjXsgsp
bNY8VjI+M48yrlPylU1WpKEJuav9TU6rV429zAO2+gYy0rmO9DuywTCOFFyL6vu1
fuCcvMOoam2uvtycx6jkI/PQTNB1hyXQcTsJxKZxyDXjLkJqEaL9GRQrcEzSsqR2
yNbITkoMa3f/BxRJb3x1Bt424Ed3qoUAfdsNJ3Y8LA7xbsMxx1r596gddi4FeJ5g
UwZ4OlXZpSkLs42oROpGhtgII/ZgTDv7xN0E2fimg5KIe1EoPdCgg3+mkKKyxtEt
wkFE5YDsLuVoC6mJ0dGewakhZU9etjh7IJYtfm6NyRKH2JoAoF/YNOIfKxNFVbjl
jZ4jnKQBmK94gdSOr72d92gJdOlbgiyJPPHm2qBXY3hpivfQZBlHzOxo69Oh4WaJ
Nq4y467FbKZl+/1Qp/bg6hZe6Wj6zD/AsqYU4DAD174TDOz7QO7zfXzga9zAvwue
f64hIxYgu4cKAEFhG8IpzAjaBI/adjE7B9Vpe4om0dg+peNZZoywYhuyRbR23sq2
z3YysFcS/Ii55Tv3RBUnp7kZ20FotUlzX4UEPpBjpDFKY3gVMYcZ/XeCmvJDc6jl
DxNO3CybfIXeIz5xGAseJ0rCBo4al/hNC0mBc2d7Von0trZf03mVog5wqiqKzL7k
0/0nyCwMHQwGvmasoZtbomYsDOIgTQb2dWuJzq1NmofB0iY+veMizK3hG2R6c6QM
frUWN613rRpDPCKDFIknC8s2Nt0zid4RvTdFEvoFNbKvAxb4ecf4LgNQJHG1k9VQ
FjTUr4xoS7WA6Y8lxojHkZHjmtKom1S28xZoxT4T+ASwBSg0qBbGYCSI596olNN4
f0jB18DRQnNbO+mJCRjBtTElTKY1xVtKzo7rq6dvpHbVpN/bpwFvesKx7VAAM6Er
d1+ZFBPT6fJDeRRAyS50HSpqGI4TOswJ8Emyi/Y+AKslL3sEM4U9Xr58lZ+XU622
LGr0Jbo2UjXp0DoeFWB55AQcc/FXUwPXIMxOJzJ+vmP66I3fMS4sfa5sn4sxYCww
diC9tZbbR7926/LfY2Egtt8sYgtivO2MuhiBNK0UYYK3pLXSXYmjZ9FnkcQBk3Ko
umZ62MUmYzvmkfn5sLnTuU5pld0BcypCf5LOVJ0MnD2qfYzfawYtlew6bgxVjGQQ
7zjgFXXTX/zHAjrj7JPrDuDVDafiOM7Ew5l0WQasMyqkM0kci0U3T2v9K6VqZIKL
7mvAO2SGbAwSYU0Qy7YcsG1zjpqopxHTDoClhiP8NrAWklxkeO0xmJuRMsUdD+Ua
c54koDeJnwh9jgMJgy45+OpAFQ6JFNJbrnl3K4VkMXMOPg+9Wv/lLUq6f4bN2cRe
xOpnXYhcxanwh4i7/tdCTproGwIwIB34NBjs6F2Geso0fcGk5YVNXmrw03hdD/cK
nJuxbqYlJ0ATxdB2zfjJLXm93TMcSUTvllnvmrThiLFZyGxmpe6O6mMarnD2RvQN
RDVMjFlIOhnryzwVNmYLW2yDNJt9HJY7RYASf4Tk0Ju5dzuTRcNBEPcWCUS6TlXU
V6qi73ykrgEvHd88fTU5dZUOyUQLYozSwfTtdkFB2HKLPT5ogeVjScr2i+DLvYNY
/mEeoN430q8ibJ4gJc5RPKGl8eg+AYMokGJPGPFJ6BYLZT2G/HlJVQf4HfRW8/5p
NtR4jHVFlTei+9rNdPM8UF0d/bFXzRDLCoBQFU9V0NX8yem0ml276vCWuxIOZ29D
7dREV+kVFnpp5HVMDjAZjSlQLbtlwfGRDe7EhzFHHWcUZRo9xC6+WvvQLTdiWDSg
w8oVrUN7j36s2mlqrZPe2UzMjNPrBCeF5cXssZrsLMIOuHcT3KDwh09tBKZGWgBr
Zmwyi1Kles/fVda3GC4u91UVQjxMsZyKGuOWRebiwOoDHlz9/fVtIt2B/mzCAdWJ
aK25JDZnt4ewKHUQuJ81lB9DL+3VYPt/Bep7LfXNjEfry9I7wCIAeOYah6jShmb3
vNHNJN6P4qaEjxq5D/jg3SB9/P2+L2yRuL9hNkjmFnc/YqXOFTjiZzCpwzZGqqnT
o9Rm0kN5v3WqNWMIT0Tuh1ug/cCH6UzA7hSGU+WzPpBtDmY8jd/HQDtDK1Ah7lNC
6vAm9ENBrW2qFtzafUZeKTqZEQONmROjZpS6BQ/H0HvAoszgdfVKRa1aQIKhXmoY
nRmOCMPj0zcnEL977Q/8JADjYdE3e+ia58be2MIwqn9ejE8Ay/fvT7DOvyOGbVZ2
Bm5cm6B/dAOMxLKv7kr4sYGMnV/JU4GLv4789iRtO3gsUjYCd1BIaxKB3Nww20F0
O5a3M0QxxmW0mY1kBzedRhJrrzgt4C7YN0nY0ZeLYBMl/2ju/nJ+f6qg628eE7Jk
m0ScsIeZGwwTr2LHT9SUvPPvSUtcgxrDXOabFxPL32vKXpncclWS1doXDDty9MiY
xxv/Ts4RkFBid+PcUfN6iLNxLxxWUXHyDy5jrm2+UM+lwhC9JwV4PXQzZpmlz9CP
u1brAerDVtVMmqayW5XYZ5IDqLLtSGVqeAjtsl8VO4SxL8yRp5YJh5TwrS+fiRJn
hFc6AvtXROTDvh9/1D+vuD0rlCQRbbIiZQsr+RceKmcHIQ8+4kDImizqFWvSKFCI
GgeLORLXjmt5+Nta8puKzf6xTBszYPWF4gVEZOL61z4cN45vfDVUM89ap//wpk2h
9H/hIW1SD2DpPLvxXefbYzQ0ttEpt2Xdzqs5aivuoP8LB15E6jUmGg5gZfZFLgS2
COJ0KAYU6CukMibI79nXVq2XF+px+vPJpHCzw2RhasgLwRgb8v9O2hZmCUWrXyhz
VCWKKiR/j/SrYoz8ErXJOONzX0CgsMeCvJg6uOjHJzfKnSEzMEkKroGkSVm0di+A
7NP66KNEaM4KaRdRBHyPsU3Q79qdxRDnH60zYLxXlRlg8D6BaAf7Q4fQWjgba0zB
OxEci1tHb9pckedLQP1z7+qhR6OFy46tLpR26lJTrleWCjx10wy6xEHJlf9K+/kP
+k+PHAEVcXumwQtQGZdAT+UONAURxQSPJzf+dAChF3nJe+C8JU/XD+LNMa1uyW+1
kopJBCsM82hc8zQNqQ2XI8XqZ6vVuM9rFI4t7kgM+SHmMTA67R7pSDtO0EbiijZU
rx3Q4JQ7ADC1qMx4lBQ1VqXhN/+4OhgNa3VWJTXABTaVQldxQjV96cTUz8Rake1M
N9f/YXSl8tTnfqGRjC7RHiuUQhvpRgcVuycQhWikMwSzucAE/NgfvnkeNcBJTP3/
SmMB4+jir6ZOKsSBE1QrAn8SRwLUNeEjwMbZZIdEgWy1fPYXHzHgXfOND9bIu+5S
S5lc9NFtRQ7wGohIxmKbuFJRVj+j1V7AMo3wnHAg7KuG+3Hs3oyESy/QtD8vUQS0
YfPmOKR6xeBbwNupELQYIg2WTZ6RqTodW5xPlH0Al+4I/zG23n5734/TtMTnP6Cd
UhXEtoHNWbY20jxAwXb3PeGyoOmhUO8ow9QCwR2Hi3ffInvBRRkr5YSkDBqhLGu5
Cq5FoUeMZXbwAxw9VPlkDkyexhAsMM1JpJbR2qJ+r4v1wx64GgjwME7/8eCQL0hE
ZY5pdIp/Gw5NGnbo/IpwcAlHdgSF4ovDq1/08nYiAPvVmZNmxNMDIjrVsiT6fYS+
7z0ocmc3/qkLtJWxrXkIPrB08IBvfmzAG0XDPvwS6OrmWPZDIFRJa1kYZLH2yuIF
zXcp8r7MTumtZDT+0wTS+/v/Qy8xWprDnZE4piFq1AMwSEuI/78zNxrySC4RUimO
MaDAM5tbPAdFHPk51q4KTXZ0gsjkaAqMDJFNQF5UqRirRbwTD4fpCQ4wje71PKkw
B7kVX4gt6jY3DAC2J8dTgWzDOb/TxGUxAYWg2bdax+whgMXO85sQuG3lNvk0PGFt
dxqwtTrt3oeQcvDVfragEQf99CbkfR9m7yZBlkxxw4g/uCEKrek2nKKXIf24TcMO
N+jCvui4C41YvTrMct3nYR3tF5Uk9w/UbU4ZFswTe0VaisM8m22MPzOYeW/6UYR7
fmDRGX/nV5obngoxr6JCEC+cz37qlV9LYPzyWdIu1s9gdSU5UX2h5L6POe+wFFoH
xpwPQ114oaa2Mq4CRwxn0aYUfN+QJxxG9ojCtETKeU+vSv8snyAtkLNQyExxIH9J
YxN4Is+fZRy45U1De+2KWk2mGHrrqho1QJj2UqfWkr2l4qCL4a6mHVzz0g9+7jb/
ymqdvigcyoA/4Dcwgx1W26Z5ksr8g3jRGTg7cGvmdKfPjPnVdssvOy55vbzj2ZKo
RHj3zSglNKpe3RDBDsDnCxTF2qcPq004Novq8/1WISoKoe28JICE9/x2u+M79kBs
cO3ZjbR/v470IzBeclsSSjnhCzHB4jD/a2wNqLR8k+zE7mUHMiT/1fHKccQMxcA0
EV4+rwyevV2T8VucG0o+QCJ8NnaI+YxvLILiidwgwuVhVRbYg75B+F+PhXEzOvF4
SFwCTsGQRu4B43uZHEHhEerEHt/9yYDYG7RQgVqf25hurDYVwDALGPXntNo9LBzq
BS04oF318fV/XREv8/z+jlFFq1xKOSlt7yU4ClCx3H+mwQ0UXruAB7mVo4xZTW6Z
YgLi/hEFWGYNhzYRI2H48ipUEEjrA6OKMUMNGEqi009H0RzQ+EtJ1ZCUf/Az9Xdq
OkmdanEpIiNgm3i1WPPNrjfsFdrLZ+S6sctui3+YuGml8qO/EkLomM8xUTijzUdH
iOpFAQKHooUzcMHu6ZU/NC1pp9l+9qfzouQB7plBtOS8PnQ/tDNtTVoTpBnPQmmY
YorH/bB9iZfBUvexg1bjYzb4mTS6k8/ayHm9yufTh3PJHKjo26CltARSUpX3CcMr
SMs2V6saFSo3KS1oeFC7HDPKeyWM1mPjCQw3d1S4mlov3gMcdnZtC2hjHcgF8lXb
ZfjSaAYWhi2S00Bi0bHQCXoyEj0IdXu11CPXAw2/znN73A8ImGrei9BlyMsPdUt2
RJcebGm9cee6u5mlzDPXn1jbwnSdRCabYHtZLxpqWnPTv9SSqbNmXJeCEjFBGWhF
bOaz91lroBoD2l2rbMFiF4EhZGalcfxb/Faed/smdgLi3RF4deh97ZGSDGBG4VbI
kEixITdOnwv/RISQ/u0FXQR3Q2RiF5d0xhwQZhIh5VuRQphtMXfuNa/oUYwWrwOX
5WMErOtdrXLrA4vTwyrd5cgj2IIsPvdTgneLNJExCiX2dTxjYt47e7zyOugmsLio
JKJoyA1x4Gw3NuCHJk9LPDLocy7U9fViXHD6jAMWoF6M5yIxaBBrQRw7ossH+idh
MN4ING45m4HLMewwZEKw4QETFY6SGwbTMH7kM6PLeRM1KVSwcUXmV8voYYiqguJ+
7B3p/takJKb1hbIjMal/dJPngw48jBm2ZEIAX8C1PJUnruRq+tBhvcdDq4XO3Jbe
5zvVzO/A2m2Nz+oX6nceV026PTrP006fEDPdM5LYn93F36J+vXkVqnFiC+sZJjmE
YHXHAwP4XtJZvDHlMxRpHPatGIrn322W6tbHM+QtANuF43Cfvqwt3VD7w81sf5mz
DSWiIuAYJgGFJdAs8Bx4mIFlnTigkphYLKAd36DDz4hv8by6TYxsCK0zm/+x5GHo
R2SYmftNSOUj3PkS51eobVu2g9SY3/pZzAiZQHpZZ0IoENO1p1Ru23rZHyB2DwE5
KTJR3pRl/wI9749Wgvvyu9jmQ5M3ZqnE9z9PuCoQmr2sq6flg0gHIlgA2WqrdYvF
Dy3f/lJ7OjHbavks9U5IRkmpHcCbggobWY48xnv1+Jr1w0yzhzoj3WQnzpWW/OXs
tUUoihmwSUgzovNznYdiHQdqjDjihtx6i5S+DUw2Anj/48CqyTz8MiJfjRY17zfV
/8eV0/oUT1yPJ0mlCz5ukuRBsOWeqFMrV/KHBk/HM4ZQkIXENt1bK1LWJ9VjxCK0
4iK/H44lYVHtw/1k5WRGyuXqxQQlyfEXMJfT2DiUlQVdMN17Q+b9lvpcICUUDMgK
W9ft8PISzIDUzPj0r2mPRUN9Ynyu4/lFbCWS3CD9zvwNYQ/mPUnzxKA4LbaY39CX
+XmZjU+g7zcY0zvJsYbGH+h27LHbRkFfv3+017kDonj1bM3TxBX/U8MO2ZD/VKN9
LZQBjlvf44Vj+Uie7cUbLZXGUDf4JZyYvFz7A82Xih2wjqs61WzS/JogvWcTmU+u
m3dpDR2712M/3ohYjPRHvbk9kiadxkxVMNmnQj69flJByUR4HYpiXfAIV2E7kJ7Z
jaL405CiJ3FPDm6pqWyJTlD26Kv1cbpLoxvPzSAijSFOdyhnRVviBKK5KSDbOYh8
dtd9VT/MDOyCnko9dGktAZMG7syxPN3bLMA77BlBPhQx9fnebUV7z+1/AMhlRSLU
TooRQ3vOXfYJSMcg4y1eL7fuZ9skgpmtB4NgSeViW+8JnrBrwsEQ7AtZtgnxLB69
PLNOtQMKEFt8+6CsuavXGAIVSX0Z2G6eFQ7LBx0hx/fDGUNi4St4Z/qvwdJBz8j6
nMR0srdCasYxHYAlCdO5t2bl+QuCyd/NfPCuJOyEH4hJtUzhFYOgUIDEWltOhj2m
ZbZW8nEyxEYZpfcMdUtiy5VROg7r/JqF/zgR/QWO+/to7ePEm3jmgqvIgkQ/IQEN
vxAzhK0EEI4qAUWY/o55T4Bhpi2x8qqSPfcsxDYdRcYK61eX121Zdo4K3b4VXsQR
i824eelK8Cj/rvlENyOQUbVvZcmxYgGUHNp12tTG31HdVu2C2UJxVqc87gDrkF9f
2WJfiTNj5Wxo8b8OVc2aPjfzMe4nF928TWvLz3vl66+ng1eSwj3aI/aTZn0cVXaj
nf+e6K5HxA2hHPueEnBgNMDebRbNRPxiVvpRC4bQCq7k/eLqtujRUA28+GW3suBY
js8ypuXipSIlc8mXqL7vaKWg0zlwLSnrdcXML2kG0wLutX01rM8J3qzbKfxfG4NI
jka5Mprsmjo/OSOArkPCufqfEwqww77toVQ7cLu69nGDiMlkrhOsfb8EBetaFlez
3Jc3c7tTVLtl7YUw7YB1odRP+riA+mjTdgdI1Eg4VGnPZHWvHuCKwtoFN117dhXg
PPq8Lrv5vbZZbOYgqH9EX4Azrv8XRs/tMsDwBtRAb6qaOpZM00oTUWTsxOIo7Al5
g350O7c7ulEwGD+yHxGS4SCBTI280wQlUQ6nblOjrvESckfsdJHGdT1sCLXVfUPw
rrdr7cwye+Oee0QO54sSfTbn/DNsmKp3Qy8QnasZLUwn7tcb5fpK8ERgDbCd3RsT
H4TWZcPcFnEPIIJiEccl6x6gzQIoHSwyWdKs3nSpor/CJOjuueSogWYxBsgb3dk8
3vxNIh2qyjVM9AKoONcHlZ2IekXW+/4Et16hFDtc96NU7ptnedUUZSprO9cg9VTW
rfK1bZN3QZTtiscg2rk1Mwfs/0CI+8Qc+QgdJCWbwdk6cS7JbONq28izzGL5FhKV
APhYXqf5SjjM69mSYcxnSc2AYCZ4PxChG7wJGG4+pdMZUAE2IQNf3jHThYQxdOhj
CUii9iWy7JEQw0QQ/XSwFp4QPQrXTf/TmPDWiEswm/E4jpcFBat4LEjhPHHqsSZH
1AMYUyMjVctyU7B792zdTNovvT7xJzsJ35/37Z1WCqVlG2SSt0DoK6/xnG1E0NpI
6wz7A5A1XyqiY1f6/uUi/XT+Q9uYA9SiTylrgCci6QHN8+0XxZLq6uaB/U8oVogQ
qEOfh8VqjSTYzq5gPMI2AjM7GGoz6FSvkQIKj5FxEU6690NIenv5mjgIpFum9qK7
cs0pCIFYc4REDHYnSRMoRll12ISDve6v2IklPsAJ7/aFpkQLLo8eGkWP9VLeTdx6
/GGS2ExXT0w3aJUUzRFnV3g48W5TFX2p+XJDXIIygd+NtN/grRuzPnZ6vjLcDlcD
J+bTJDQwDXrH5ld4XYIWVOv2cfGIOWygpLcFJktUwca+SwRNsK4TbyPzFirn7BUv
8q8hzfuzfsGF/eCVXfZ9tvrwHuqy9670Xj+6dtJeM8V3itIclqT2q/sqYdkQCTsU
n8MBXUSorACSahUvb7Q++0j4Gwxm2LoW2ljewYr2bkkSLPFe0u/sFyffU/d8SOz8
C2pPs3SStyo3QvOvqsvQDyXttQz/K2/SHXU+bpZHBjOijyq/8b04tgdWaOHt/KMG
WQ3k9jy6sOmXKJDU3xxHX+yudRf5GeQD3qK0pANmznRFQZF8LAFm8/MVN+r3ezkt
xLL9IWrde/skwKh0JjS6rdAkuHmdDqCCPWsDy5ueWsNd4YmufVhQ1y1Xun0ta8W7
AAmPpeQgCbVvtZJkxmmqzRqU4v0NjQZH1DF/1opgWFG+xQ3l/NNdxt6sn7x/1MX6
REajXPu/rqnu+sbJMfI36WqLf6GPicypm1DVMUPh4ac88c5ldoaPiqX3dR3WKBv2
gcfvnCsUQNarJAZQnbbVABqgDNjX+2MdqQq1BGoA0NHTEvAS+giKA3v8Eo3EnYPN
uqxZNSQSsvCXmSAoTV+AUsYXwvvmwFjWPxvUcQtH5NP+tTp5e393FDlLeIo3SK2t
s70tVYU2AmnVFJnYyinsVUXl4PgIsbHKFJ7/OzSQjBXQhLKCqEBDVqLbgs5+WQEJ
cy5Y1yX48CsPTWVO8gDlIuv+9869QI/07BP9BOGphZodOjz0u7e5/cgiUZi/nYW7
NWjhgTFdA/kZqmzIqY6Y35lXjHjr0JNKHnHgZiNvdHBMiUh7SoJiYNPxXqRSeOUf
FO7KKUtQCaDJt6+XzzqZu+Hhg82j+S5X77QrLZvpNH4Dt2nWheVYW0EoLcK9WiPJ
Ec2AdPsNNZcqx7KFsWaIqFVk5knjBBIixLnZfGtstrC0a7EMMxRYrbSDcAlTS0hB
2bShxpsfraroslSFZ3Sf9Zv8vyk23t51NGSUvfH+2gk+8Zv6B4K5GyEtAVkXwPAj
9Pm2E9hpLEL4tfJgq16wIbMk3i+HracnRH5DEVPSE2FhAwzm7ccKi3fzOsgWTZf3
mdxUedpovg2TZMP9toNsFO9YoaY5t44d+GJP/pIHcXxrZ0/B5+p23SnsWIRwTlES
KGLz1wuTUPgZ279OfOfeMrLQ+r0e6ntI68UxMEz3JcIHBfmfuX1VLNKsGhLNo/sD
LD10YrCvA2uv+Y7yeE60CO9QHkucVI3jwMhzrS0nzG0TTgPUthPFxUKWqJm3E3Vn
f+DBFoppGuxAu05PIPB8lr/9nw6z57Pu/XKJAoAlMjpbgajFDsbngAugY+7cklpO
fhPEj8LHCArk9wUK24lf+aaxZWYVMxCf83koXPT2aYUUPGcpaRU4rlm33ydutuys
hYWAoC0etQk0aGopFJXKM4bRfs5r6jkh0Xl3biqLc2mXfHGxvk9R5mupTtJffJyt
tWV+mEV5zPLcmLcHYA+u7MtwcIngtgr3PLigC2PjtalUWWROksVEa127CckiFQ71
sDwu9EdniXwEuCG2qHj2Ux9UVYPJ1Vns56zsSJiE7+NzxsmvLP7oWaJ/5pz9kosE
AF9tPTpsMsBxID0b4gs1zaM2yl1s58TBqdjiVgQ9WLDzWMyDKmWVRKHzSmRaMlpM
c8C4E3XsnpdgHD1/d9ZGrgIYemxJIyIyKOJGPaIyYn/Q+Fw3wg6qvjYpqicifOBv
Lg/OJkz+R9CiLd0B4MfsLrAgZHqsPEae66MCtDtfbzwVu0ni3sjgugYfTQJEvq99
G7Y1v3NvSLN43X9zVcTF+1uTYWEPwxZwT4XBT7mceZd213Z9uDHLTY35xHlJxFwt
ChsP8Pb477vfNqKM9Qw3KfsLUFDCjaMuzL5ncAZFNespxVMOQmxQx4DJnuzsxsWM
AX7ZzF5GwYqc/CbPPhZEIBy/644poa8pheQROhGANYYakL41tQz6Y9cem9ECsQwD
RBsLfZjINF9l6iSajYYeFCC3jdR9meZy3XcWtFPwPmhGelWdrEYE2xhFPRAsOgci
X77XM71dK7Zf2/VsNQGF1OEywnH8meJJb/VBMG3KMm/ZytUoF9EgM0rQ3+uVIzCf
Hz+jU/wrENfVLvAqMjjCFrqfg0u+LFkW2CALKh34eQWp1YNVc31q/4AL3caIOzv0
xzGwh2XX5XaCJyIKfQH5CvX0udJQzUsLnxjxmZR6fva+qiQ/PwoWc76CnDhsIAK3
075wifuSPK+PGATQm3tmvL+Yh/ywHEeCDoqFCgmqGw24toOsm3fXuvzhpIgkxLRf
m9q5jls7znzmwPMBRBliOmv9gcAoFrCP0y1+Wcq9Xmjxo2+lhOvYKYxiIwYDP+1u
aaTSTxjOtltaYuCRDCGgFP7B2sZGwi9GWBfWM4vKhj+V/WB4cw6ymiuC3Zu1g2tE
ZUoIsNswiuVuG9o/phd2mhVcHeexS3aA4VqZM0AeLrmhtoFCZtTvN0P9ORHXn9BO
uDHreG4qHKQUTnz8k/j+7U2lGBkbg52KQMP4gHBk1fcHxQ6s3cDuQZMd5hVASVjd
cyI/eOhPBoeTptDYuKRySS+jaDQ+L29G6TzBoltGZNEnKo9rJH5r6i8K06lTfFn1
5gfXvaWzzPWCYOY/NCRXLxcOqJNxOeSjl+sAfm5prAD5IAdrVq/QVXkHkLHElBdI
TeSipKdBSv/LdDzoFv7q9G0T1KENEhWfZm16/qhGSOL0/zS0IWqsGs4CoF3IGvdl
WrEt9O2xDwAJdyKO4dmB6Wngf8Qk5P/D0pK0hTAwqJ+d5OcIr6o2DYSTVFkmBSGA
kLeppN82MCh/0Yev/anc3t+4b7qJ2Fgzqmo7I4Xrh0P+1K2quma5z/VHafh3seRQ
enCp98s75oRKxZjYJfBtHJ13CWGvZm8NW49Pz+Q1ae61Y7tIlgzVpz7rkxa7DXHt
Dsmr+a0d9qul0Cob0ksv00gI1XGOvHrO2Wr5L3/AHUx1ESlU9etZ8TXLOIQ1Gv3B
aLy0odTAt1N7s0sjHoKxIGVKi3g7PPslnqWMMrz2FJKTtoUTYdciPnRgYnSYCon/
ZgzEMT8n3HxE25vn8GWiVnZkChizd6saD2zf437G1lSeUOoMeaTvckbLYT+NPx6+
w+DM8CLQPATxj1oSN8SzyggfYK0yZgNtcduKUx42jiTYk98BUJEYiTiiiy9oJz1Z
HBGwNKUXuXp1Hn2GWTFgqQwNBKXR9GUnAcdis19amCqX4PrOL30MN7oLZgmjNRFO
RsYEoG5iCwsPKKN9d5/ca4NEe3LZZq23sDRMPG/blKmYEHOr60G+q8b2p5vVLi92
ChsM+qXcbAh/FWZlNgSShE0zsFaIT/RCd2A4rZqh95RIoz5his9hKscTvWukLcVn
bEH726osIhVYCKjM2lNVSZ8+ZmmkNXhJpJxyQf5CATAAt7YdpIa7XQGHVcjcLLgp
NNLSAszcjMiAySNWcLBykUUByuvmD5QKPgHArle3xD/lpxZm9U/tkTTF/oHhJZSm
qKQ9cnIf/hLHYFikAh536B0m1x68TRqqa7FyKSC+ipIGw895YIstf6fDc/ViDOOb
W5XvbfXuM6IZVCjOOFp8b86yLELBl1OfGgkSV3rkr0NyhA7+ctZUM/hgDiSGeCu2
dnnLg57CmGTETgbVL3CJ7T7si6ecA2zC26MdPtVWPsoVAc7sD9iNy8fmKOaswqsE
21E9S8dRHfPP5SESVRruYM8AQr1tyQ0Lt29I4zGXkQLkrwbm8t74N0fTJOhm0itX
2ZeBZ4/rfctEqfi3CaeR4Y+K/bQgzNfMTZdfNC1imMhZRs5x2/Vifydz4us/iHYv
GMILqR4/DnbgsZWNxt+3HXnAvLY1XEPPa+yGQFq8P8ladmwA+XOmNzFVyTuPBgqz
MfQrJzVbRPTLAc5T7gcjTkOoleSFTiVeXrNagBp1oyXQ6yivugeLMJTp/GjiAK9g
S/gMjAfEEg7wkQga7zQevYGfyiGaVZpmoqknSi2v6dceQ3xfSP2tPy0ThbKE+Ecj
fJyr1ysXlf7W4u1UUQAA3ipEsSr8pEUKYUJnoJJ2sQFVYqQaqptZn7yPG/QPDF0s
9UynUkt4sT0C5go8G2JhmcxW8fkpQOsy2Kdad0AIeO1qPtR5varCNTbLn0RvNPe/
GBC9c31WesJHGo+DiEX9ZrG1s6TkF9Iw4558TjB1PjbH7SKC076CtT6RPbTeN+jb
640JA3fZR3l1yGfVNH3ZMT6/FhS+cW1M+SGLnRKoGm5MeRO8qJvGYQVjdRWDUIr/
GhenmokYfi8cK1L9VBUPlZx719HSjGgkr1Rwosoto+2c5QFPPm4vP7yJdi1e1uy6
AxM63UnLCZD9b2hk9Gdhq5Ift0y+lkXQ1zU8LUXx4nIUzaO5SD0nZ9mjQLcOi3uv
EzMwReEGw3e/x85napz8JyD4W1Uxy3GgeolBoUCtkq30+wQC0lf3tUBrmDd3Sqhd
aPXOdMG2mFWkQDKbvJ387TunttSpdhuHsB1+Qp+8JsrdLOV797kFS7cvmU/szdwT
Yi3bSd626bT46ReoDXLYn0YhV10I4hBerNEhIHkaNyiH79KOvVJI8jt2mNF2l3Ol
udSi4nsQXBx+vWWgoFMzTc6TXPIbTaU3oHIY9+cBRW2I4quLykfxVhM9XdvAZJ+j
GW9ZVVL/oWZ4S0cZ76ZT4BYqOhcPeZMiU+gC4IChxwXW6PYMJKbR2py5ZygqViKR
GosJhAqzLU9ss3nSK8bTK8Io34pZh6HMz82gwvivK1x+9dv/ZuEV7XHNSjEghv27
L/GH6eosOYC2h8vI+yzi1otdEND+x9KpRDpOs8CG3wOBIqNoE1MnAocXgsO1k4Yk
35/JSOq7u7gXeFN6DNslsYjwbIGTpktxmikL/usCgdsO8v7mfdAj555KLxLbKtmO
X9ymAtPPMU9O7CUR2Y5e0ynuLN4XBCvma0cPLDycQZMGLWhrPb3NuKF3uvp3wZdw
JeEsENNkHMGrgpVpfPVgcDniubYuQc+vbZlNrIYBLjXaqtQHF8A5m43O7ZhCfnyO
/BUdJEhhbhuYKKFgwD+9Hi+aRgQtLUaqlJlwKctqWu+7Gn41f3thF9qSsHIdzZIY
2MCrWx1VdYZPOTQHMuu6D7stQeLEe2F/ctB37bfc/ZvwtM4shImPtkqu5QFMiZP5
rhDsttIuowEijo5QO2rjtWeIC3UC2eMfnEb9fKlmZ63eM2fiIGzcTm1qASYii0rU
neNnKgQ82A84sZfkO/xj7dofkRvQ1MkUEcKV5WIp9bzoXQSbMlx7SgoMh3Eu3lF5
aVvu3LwppuQH5fcqWa7TxdX2pQQzjnz4eKKkLScUnK5Q0CiaTZd3UBRhBOwQpLC6
3+q2jBs2ojvXcywl0lvM+Y7tuMghfatUY5Oox4W9xbzHgGHq9CSSqKgG3XkCMu5o
s+KsNjZk5eqHf4mN9dLHGJZq3ehW1YyGiPSW09WUvW4xa0cOZOGWKSqRQioZnRxd
mJSOTAziuPG+xoyq0Oo0MxFdZSJP/PCB3NdHrjn7beeCilc2tgVN2Dg/vRKv1vNm
2pgnb4z5v48XIbsWnVNupcxoGy47yAbBp5Nl2UtdjyYtjZR/3vN1EbQXeyi0O+QV
aQx7acuokWgrTrvwvOiicVtMdsHtQsYo03IU0zI46a0egjAjLTjh4I57EJty0ogk
iQim3957qsqTKj+NVX/gYsWXRzNZrC3tfzx3nk82uAcT23/Csga9cum2SzV+XZPW
tnEdImVR2gq9wMo0fGer2mGwJg4zPsBw1oWiRhff2Fk4e5jcccTAxEJUmfWPubXX
9vY55h0YUCEF+S3IjyKN2Mw1LqV8R+ps1jkTW2yEMrwhnkdkF1NJ6MZpFyURk7r7
59C0fk+oGB8JO5JiLh2UbjCR39F0j+BY6gZli3dnnmY4WHCv1wPn94AN18nJVxN7
ZTUOXlw5Oyldr/tpOhaJVRaneaSEhxwpHJH0E1g9+WuXHr8Myx1KSdOJcjGuA7st
EM1xDc33PZSPKxU+QXb8mw+BC/y+Gq6mClq2dfWzPyZReuPzNxVu1tQwSMOe67ky
VVq/ETcXLFy2p972RnlM11afpcQEJgV2SYF+ekIRLw8WfZDdSihScDpaPiZvZLFJ
KfBHv2uQJfWj/DqN6PHmlyC/Vej6DZtnjHe/t4Z+7BvDCw8D+tBtbvgtB/HRRe3y
IbXka8GBb8KzonMfHkiUQXBw7WAa9MR+yaCeA3dgVOqVcRYdbu7gadhhK+Vvuhvd
XdrlCSezC578oQumUg2Uc4R6LY27xML6OxJ+THx4heQdVjccYVaE3f+A4Ijr7vN0
WPdaPXVeH05qtQkLf3DVISahWE6fcGYCcm9wAbIIqPdwpcqukEdOok9Yg9+Z7qzi
B2tuGgy5ciXsz7eTofAu2A1mVdsrjW51WPq2iNBGwAb6B23MfaOqXfLcaAjxmGG5
x1vUQHt2oZod1Cf9Jlx4DOxQUoE+kk7kT0cZVR6taoHwcLM/LQSF6zXXq7LFdhXa
8CaSznUYwD957/COlN9+HAXxmyBuVjGhRbhFSa/UMbpbcS8MIvUhR4KhfLwWY7zI
0x7JESpSNjCHz6ffuze4orV72PTEPTdNXrCFn2S9Plpj0uAuhcQlbcAZKNbfXvZt
Sh4YuCcHMD+Z2TgXJO4Z/1or8ShuEHzaXCixPUUq8ApjmQurkNZ+BZZ4/lKxCwFE
hHbuLKJjpZrDBdBNTN0uGJbCbGWc6f5AUmKGAhLI8GhwJAEnYKPy8LuKwlmd+d6L
l17RA+taPgbMHyQZQdcbIOvGV9g6sBBziI9BdXr6SICVraucv6jTGWs3h+6C3p8v
gUioOE0Pzb1itf25rxwn00vVfdT5n0SQnX4AfyRyL4azjutlvMlbfYg2CkzyW/2l
IVD3QuUaCjxkvJAHugif+cJnqAiRfxmmwobhnz4c7MzekE72zzf801cAJVGCcatD
kco3pIvmYD164vo9Q538g9DZV90RjRgO/rglp8tX7Cotua0xVYu0Nkt3mMUltry8
AXOzJmcyj7siZvNFlPrywQAeC3RpyGhrLl3083yF2oRHXotE/ySf5547X662QQNw
2rwwynrkwQV1xCTAkDvZ8VDZtR/cGAjWAfzmg++jUIp0GGD+QghyICw10gJC73di
1C4KvXtkqehvTNajijVi4fBL5DkjTZDy6Uq0/8AtgC9Qh7KRRveFVFsl8z/GUB3i
R8euEA6TPzqSKe+uZFdeAwwoXqQwwJh/+FiLFhOZemYrqMSYGNqpINexic3sSlW2
FFO4MV7vG6PO++Hy842s0cNFfAswpE3V3CWRYZDkhCDTydNpcTnZd6MMUKtEuujo
FCtjma2v2A2OlwQePaGhjgszlp2olz1FizY/8xjsEQJ8FWvqbPGKanhcQfYk6X3g
S19V7soTEn4e49I6yQ3Ux9eqqoANndsGpr3pXHUdgkXCY9gEFnvwGQ3L6LojXxcp
y4CAnCeLAM/HInq0PX+QRywkAXVulop5mWN7r9a1062KekGUd1XHPMceqbKkkpm4
wOpTO2xq8G9KjK2MpuhnjqKiRyNGltCOKUQDU8kz4fwlL7Z6klesSbMfjRgolGqd
FzgieBMMTjMYXC9OZa8SHNOIVJN0tKFmGoQa6Vm3VQXElMN8AjtL2qQ7VXhCnFdm
MOV+k9l/u77y/XgY+ib7vy7EBxJTuzSw6XA143QkQR/+5Vfa4tKS4PsB90Qsf+te
h9qQx6vFEsyhmnsC3o4SZf3uMSPnIyARTST42BsQqyXtvyvk7ekxuBOXl2w/MzXY
tmI/5WaZCTpqFaf5fycbTxsMCRz1OYTI6Z4xG9nM0cVgft/mY5riclHiqoZnT7LO
d01HOSkhiliCB8VqHBCuOQJ4/RN3yF2s6g9WUlj5/UNuuG1E4cVzHDLrE7OSJv1u
XAc+PFDiZ3lNgU87UZM/jl3kgHO+rpE11tvUR8HCEUskJ2SE/3XL9k1q/oaLkb5H
JzXyevI2AGxeHd8U6IYzQwKbdpTdkA37tsvNEfadA8x2gfrzXDHymtc5OK8VGTnv
byG5wCnUwpht7lGhb2zF9yTyPQGx9h6lMgW5BIgwtqnWqzR/mR04X15X/LRRz0Ll
ZJLMukFzlYp1EpN6O2xaUWrXPmMmDvlQd6LABsHXcXepUVIQ9NmIhebQZ4+ep/8M
hGRAqU4x6tSlrmGDy8PFuDvYMg6cq3hPMaeGsFW9bL/UU8B6kKR4SNTKIQh8uNo7
k+nG+xoDyqPEPRnCF6kfZTYyG+70SOompbcvmE+I9TQzaijyyP89Eq3nBWq4nLvr
UKx29PSh3LddqR4BQP/mZIR3IViYKsgpq6OyS8dQDT1in7PcUHXxARL9BxjIJCiO
6XRz7uaGbOobYs6coKoqjQReTGAUv80/2n93RNyVlz+MwrphzKCx5dGyQn+UNMOZ
CNcx8p9mCWrBQpixsWnGogW6TWKCz/Pfb05n+e85QTnsC+3y8Air6Ap3zPzxlNdX
fSMO/zmUcApsyU7txZLKXDds7f0W0OPq3eCpfwr3BuhEfOWCALcsia0X5FZOQv+J
wNyYZId5iSxuqaqC3F9WfmKnGj+aEUj1M7UlkFqHO4NHxFXFUaol+L3GtVDOfLkk
EQgbZK0Zmc4reuU94x428jMYzIwNcvlALylDj9zsUHeG40AhTjVKqf0XVqbXTEgp
a+IuxykMiRc/RxB2rxzvLNeETzx5k7JK0R9vEnLHFReXNqj8EVIo6W3yCDIerltL
GBNmqbtbbtJU9HSpzBg/9dm1XnN8aOeoQEToJlGwKK6vivJtsxn+WLBm/yS04cIs
0Ki5YrirLHYxW3xojvgsitoD7GpAzQWi42cnzZRwa5o95/19na5p6VSdBZVD/SGl
s2TBulltB2Ra37aR7Yg48IETBQk3mxZei+n1bMgdRSEhROsktXKRN+M8E6EjgmhM
k8WLRwt5ptArs6hKW+WvfgU1wb7Gtv+KouOojZjX3lCQFZWa/XgXlWYg5LLorxTw
bnyrgs7NyT3/skG0LAatHGfOkJzfiOT66tcd+a9kzwHiSNPnFYd3Ut2ryDiCUruN
tlp1t+o/s9iuA9BPRYhvdn8W/JHoxc+ELC9znnNq0SIg79VOpD1GUmdTDPtsdf8s
NEp8zrcWNokyW3ZjJi+7dQv0vejk2L1ae1usZUpJRZJYUvM0RqutC9AZWjNQgFL8
qKtjik3fM5ciyfMogCOOIHdFbEWVS/pfLg5xVuPCYash4VUE8qhskzHiy77lsmoF
/Lk+C9gECL0c6CswOp4jBK7Z7zQy2DAlhN7MmYKBfcazA4KA+342lHXmkWAT+AIk
SLHqePAa3hzAR3SGwXFTbgtEW+jdwnLHoyYivI4htRwOuoDfoeCVR1SaGCbOprQK
t4SrM143NMIOobo5k0gsWVcgxyGpzALjQVU7u8nWL22MH89mtTLT5E0MfG1wux3z
NeKDYerrh1fOU3EZEW8oIMrZ9GdPgJqdxeKxp3HUap2Q6yvodAKpt2/VjHOxoZKh
NVgzCYUoFVgGESkljETH8U+PMHJC226621SduFn3urixtTfABqDBwZhrRqhAeO/a
kA3hg2qJfXj2v4/oqFgTsgKq2gLKP2Y6ykaCpm7aOd0RxL64IIMXrnDLWroGX8d/
68LL0t3gfRT5o6w07Tmr7P8Nhu6cTYdSbw6hryQVnyI+d4r7KLkmVjV0IRNlVu2s
nxZ3AA5R0xdMjCJg+PNMIBqNNJ6b+JwYTGQE8+Az8bBa/nv4ktVU0f+4DlA28m7v
iNHGNrf/DaiHBkXAJBCA651iv58MJfQYUBu8tp8Z2Iy0LlobPCf8dmQupRxzgz5v
0sJcgVkrfwqV7QeWB/unzj6oTvSghlMO82CpbONXfJ++ZwD1BBzSWukCG8MVlQhS
TTEwjd/EWxpNmatcErSiPSt+pfyNhGUMsUjtPSn3evpOwVbws7CTrkMAxYsHdDwN
SdFY/A2Tdubk0mVjgD4v4HPgnMgEkTloiEgky3xPldR8Kbdt9IkzykvxaOjaCrC8
jqphOkCdHobbaFLcBQVujxjxmCnlDEwwKdfbxi+deLbW/SqaCVefPy9NJ/CZXhL6
zclYKbOPf6MC/qEMwayCSV8k5vTEEwp+NRvhdEB5cOPKWI+8GJoQnGxH/qddZr/s
XsnpKds9JRev4TNpMB4uBaOITjYf996izsK31qgol+UNCuLYaP7LSNemRCXUzczL
s9jIgHA/RitEC3SKTxa0O/ywMgQvGgVElZ1ojAMB2kwIxvniIxS2NgaCwG0YH/JA
XNbfcae2FMLYjrwM8COIpZBzPV58lk79+s4EgqbS4+qnEJTklZugPjsDPjZ2O39N
Ubs9h2SId80XCVh/2PO++tJCY/b11eQZhXoTHlV4+4EnIinSjAGiukpFPiYTtoW8
5XRJV3CZUAuFkx1ddf6WWhIToZSADceDKDouOBwQgGaxBdvx3UWLw662VlEQ9pLw
+mDEFfEoLsNJLXE0gMzGQFoSODtmMzQpnpD9cnuFiLYSFw7coOSF6QGrPY04D7mx
5sVZuxDvf3Qa3yI9pUqTR2uqnP42YqgfhdwTINQ1S6oBE3k9oMOohPCWQUHGNvYs
iy+jNB8/2kXykqX5rcn0tvIt9EfE3jOvGzZH1Us4JGu0GdB+uLoy8NQq0OmW0N/n
IDIRstoKjQ/3bZcvuPhdgHw+Eva0LU+1ytJxKjr02yyRy29qO0DjCHXRjO2/C/32
05oEXnua6wvNnFof7NzwbJioy596ghKYRQZRcTjUnz00ew+ZhzhuufBXB6g50LRI
IxeO3+DlrhJoA6jtcEuESvrFuKnF9Ac14K5ZaXOwpmvhhLZzkRvWlM6hIhVfiNLq
bMRESpTTz8obliiz44HL8FcXGG4r3qCYU5zmlj5OOYweneQVkvLMj5exE4OxcfEF
+QSPdp6O1kHzO/w7VtUXLaB39T9rkFct7ZYZe6NJFQKDWp4pJ0XM/4bu04Oaj7UO
FVVs81hnrRst/J5nIOuelzGbjBJ3IiRUJJGiow1nJzUMIwSodP5BScfq4VL9h7d4
eWD4mDCHyLq6rMOoIY1FV3NUOTtU2D/9LF5fqDBx2o4b3upW5wNywa6WpDjmnsba
kc0uYsnewPLuJcPO81v0tvWmgoHZckPT2gvwkCufhtCsbfAn0r8PX3DrSN2/Y8rb
BE8Asfx9Tp85x26O4mfZkBs6UalCaazGXZN/fEg3JVyd69FWVcqhxEKJ+uOSV1us
m7OpmkSkbgVX5FtjRJiUdyGcYRC3Guw68/s9J8NTCayxT7nfz2mIAgrtqUkOF/zI
jMQRLqXRX20KzjNZLbp1BWLlPvW8PBi1Pw57rNEAG1aPysVGFCKboZXmMQ5UImGO
UKL2D49Bim979UK8RS8Ua174QIKhC4DfssC2IUp9lxIIHsz/EGZrZQrfJ53gAkLS
M7HGOWgwm+3iaM1EtjLCsLt66uDr7Jj+K4bM3K4XVoAg/mP5b2lgXE1d9rfySzCS
x6xNec4AWOsk1EB3uXRRF6ptrUdLhe1rO7pR6VYwPd06GkSv+L1tKnufnlqTLBaM
FYzj0pTv0KKcwmS7sqAazeYYnmbrfkwp41VzG11SZ+0zNOVQXP50GxedXyNIwqll
1T9b4Nw7ExB2SSLuFlDd2DikmqIQcfrf0xJaCCS1sRXniSb3yy7yY33xcsuLdgD/
DCGmk6j1GiA4P03psU+QsjTCTOygZUcTMB10sW4IPyJ/ytKtSM9aFam9RJXR11lb
nLLa7/hwT0Lz1fILLE0sxaMmMOk7x7Lem+NiQtHGSiBbag/aP2bj89taeRh82A7K
0LwaozhqzfIOrV+3pnp1KavCwAxgLqwMkUIDq4NKkuevVM/zGWZ6EGMgTPXz6ekX
3585yDOB5WdCul0hMAluY6ZQUP0ZVlllCCyb7EMPE6lHpCbVq76wSF3GX4O0j0EY
FkmeZF5hq7HPsOxeD79R6yAaKTWAxC7bDzeVRULQvzK3lVh2uXrEkgDrNeNsQ4qY
GnGQtXJqRbrSc3qJAQTW+W1G3IGWliKTQ0y0QB5z6GNUBqtTwizCx067ihlhs67j
aAh060nRUdl8fNITrfI/M+3xvWsj33pXGtY8H0XRgA4FtzXSNvlQtkO3BY3q/GWH
KLvvKBl+drJE8q2H6kYsAbd091sLTLvp0mn05RonqUPA2VAC4GojcHnxZezoIr/S
1kkYXqgifZRx0nnWkqxenfYjOyyZ6U9QzYd1ywvaPFwBZSy+bNRJIm2cS1q1J7+W
HoIbGuKJlxUoEF5dhjJeuM1DZ4gmy8oBxgMtnqGJ5Oz8Gt6TIlkswot+GMNWZ5a6
it1UN13W5dGQ25BakK1ap7Clo7w4PLn7DbUgP76y8grfFgcZ3R+6uXAsepnaiH2O
lDxC/K8FqCHP+wf5KVNzDARGysmZ0TNg50ISjRzYGy90LIWAvyuyv1xJp21ETyfL
w4bkLsSxCvA9rBfKFlJDPRUspETg0BK9wzxACv8gNtO8gxRY9NJz+nZ/f2uENv/I
ZyDQyf69lZdsALUR+a0iaTcED0iq0Gv2fBn6RBmaUzjlwrmQqsbUGY+c9FrnuK7R
C3RQFpdcmJRzKCvuFP63NYPniQAZ8mThFAV1Fj/UAWLwrlVG5gHuUBLR1xKvxav6
rUB4veDRAlN3xUDf3/ClhUsFBjMBF3kGZPPh2uZdByv65B30GILj08/6j0kFagh1
LmNtqH6fEbddJRZFSm3JWyKWcabuS8pByzrU/aId9zU47hh9PweiD2Znd2mLw3tP
3+/kz3Xmw+Bfi2AuNHnVSlZ8z1Tq6612AR7ofcd5ovm+sSKID3KSGu8nfl/AB4Yx
H+95bg61fEokNz6XUXg4SF9964n/wqhOz6IM2DDCOgLMa3CGIhyyzF9xk8xZ49nx
bWFyXfbdgDefoHymc1945TVjK1xlMd6GWd6cmY8Cn59vFkKhHLmo+Tny2kX0vbli
M6gzB185EqhH3z3at5HrO0sCvTLdTWwbHqvYCu25QoafdOWOm9lBGIJ7YNXerCFf
GAZA14Y5KCAp0N7yFIAIiiX60ru+/fPnyp4vwWysX02fuD/dlYBEe+3Rg31BepOV
tP4FTZla8OBtvyYVd8gIeVlu3xeWhemoYVNb4cQThRSRoSgi+8Pfm+am/jTxF/9y
O9XclWeNxargDGgpQBhtGucCkPk7vIWR00TE0fSIb6lahvfgnYRdnPI9CDe72cGP
ICwDYVdiYtJZut7PlUMqhu0E3+5zCyOvAu9IvPjhn6Xe5tmBRwvCqtWR9GxoG86d
FXLCzhHwdr7kFG/s4Q1yn8fncozrUtLRcaQdXcUt7VonW/NdvQsY4QzFmxT7XsdM
S1ynTtZsuyLZFa9xZ4nf1DrT9jseSJwzTgw1g4ql92LTc7SsF6OIGakClO3bzamU
wJpUxB5kheDS8GwmvdcfBv95wmGonuUkf1GeDfgnTimjn16YrrJEiZ/xYlISeaxB
vcUUwGc1Ot5cblJ0kLefAiDcNPB06XDxSQHESoq+Taf8v2q6JWHV/xpqVbL8rJaj
nRuFNxApLVqNLOz7e0s3JhZDEx4htobkFwtZIE20W3hm28LWtBRXBcyH8z1ktJaW
EwF2XJPEvUXsIShoKVif6+YfZFlCI75ZQmROge8B+BzpSlAbZgoJXvo4NciOvFNu
BDmbc4mErRr7OUtNmSqbIRZ1DDXQBTIvu3FasYhoheQoHaX3tXD28KfLKGPGxfO5
Rq3qdSK72HLtrrWRPHEGigcwcHR2QfFflKtSweh6xddjJzNxlZzsMo9ytM2FlF9e
MVVHSoaS/3ogCZ39X5ustrf7HXzcHYyWrIOy6tHlRMGseAuEU+6HrvM77Z3zrMjA
33lStOMX+GU+MsQUwtW0URvFSsDDGfhvSYTYp8msaerQWTV2nLn5bak64doLgVWz
NPNSuEEg66SoBWUNhZpy/vzw8SVJ3BVUnjyaqivFpwW+yW3MwzAOkHMx2AhhtThC
ODXYZImndChtEmBy1PHO0S+sG/l0XvLJogus2xt7Oqk8TbeqD6Dl69Hd6fAAsRjS
KPrwLWL2SlzsN+1o7II3ClHPZzpxlhTTrgTCLGHmNj+tHNwO0/s5LvsvKVC+KPwq
M6RmT8XsHZFpSCG5LyA1VnnHEwNvyve/NnuV9/0VQIAbZtbbiX21vfWdjjJLZY0m
RpMYN9zfwdM5WGRROMVZ/znGvyEkJPdKd/pfvEZ758R/UdBT/cigOUycPFHw+CNa
092JN4IlMlFULS84zRDUmlElioZ4m4Vh1+8Xo6iRe7wJAVSL/JTmnDIHiIjdTs/n
ftgYZO3onpLwnlglAmjgs7wzc5OIf/iopLbZeSWiST4VB4+Vwi8UXwjLcLwyesss
wwaQ4cAbgbURQuUAi8kjj/l1pa4eGCG0wQrz6waNigvIjUa4AkTZvX/h7dipxoxL
CYtNfAs1hOLr7jygpN1dtj2zHxXaEFr6bTG9c+Q7v5Lodk8cW+uFF3XP/M5NCUTp
uMN7g8MPfroQoT8R56zYp7p7oTQQw3cdw6+6aH6yE3GJl8HgDfsGl7r6E9HvYnzo
Ob6Z18pSkEb1Ly5zhCoR8Jt2BC1ZefwtfTiR6W5q/EeFecv7rdDzAoXjuroJhTEp
GuFkRYRSDUjCEDpS0+wWZc8YxhrJqViqjwOFuS6m6Bu5WHvBPfTjStV2Fqg5L4+f
UB/AedAYXTb3Ej34LCbKcMndRPDa82cUMf2536uq0qgp6OuBROWjjtyzfbZgnQk4
8h0A87BYBBBomZWGGgbvhM2kEMFVoEbwXDnl/IUGeMbcZ91CY8Ld4lmpEV6+SyJ1
YzjIXzxIYx07lVQ1eBHRLsp8xDuoea8EsXds50Goh0usXbBMbg9p+EY4LQ/q95tg
QLjwkFNa0zipFNzXsC7EkNtpGVyF14UjqZyjm6JLFxyQldv9xpikJn0v1gxXe7R1
5HyHBXfNCkdBKEhVI5Au6AbS1kqCryc84oEQUKi1M0C+n0cmdadKrpCWZhFDWx0k
ohE6ISmbX7YJya4izJTazmZRY44iTbRBgIcqKcJ5KA9G4/5h36xcXygsGBspWMXw
DOWAwrT8AI2MwlHxWMZalnDv20M86xtZx31sJ1ZoJey1rtgcyFquc3HSHfiwWOsx
Yqstc0+lnXPq/VNzBG1/++crKSsn8+5vPWULUXCXIEPAelT/Tob2hSJfN7IM34QT
FHaGXf0a7/Gk1WacQkS8EHgj0R+XN/XxBA/r/nSzLpf9NwcyOAkUEd3f0V+BGqHi
NfOsurIdXcmFBVP77GUckC2VcY9Hyxo/Mh7uGYyiPLHLUkLwUTz8l+ddM/qRyY4n
tu/fhjSosaSfe2b1MCrB82k8hRI6IPchLcVdb2yZy6lvkFtwrh+wUKjPp4K3s2AU
HwsBlVfGfDNasx5xGaTKtTqGVuFb3iTa68Xz8Ulp1BxLda8DlhQ9Q/4aQEX7Mssl
NCd+y7FWIdiKE/tx/LEbMpRHhk7AEH8Q1wwDIzoAa1gfabin8+rp5B0Mo0vw34sh
0tN+geUzQQN2M4PuN3UlhLJrRO/eazVIS4pM7gUddYcx3XV3nbRIJdRjf9Ce+ZvW
HYOj4LD7xuPKXxoChySM1oNcujANOJ1nxG/fxDZy61fVtVBvDSBSAdO2W9pBsZEM
JrzmKQo4Npf8Lf2pmFXCWDY9X+edYwYp+4sI93TwMXJAqdoYrEHayd45AnsiuPVz
gEQIHfRpDqo0Xi1ZhBJMBx0T1754ITZqPgh+WtyqmqB/36tMpus2R8ZN/C2IbF60
wVMbZsSlZw5anrQlM6I1OwfFzPVMJMXZZVC417Lc3bbPlhW7fg7m2mYVbDOIMZV0
+ZBZq5yVKxG+GWvNlsgZJXu1+okY+Y0/kBuxXjQCOSX6jOO0XAjoiRzrBwNbehYa
XuupSMqDq3wkFaIRBX2wphKr2RgjD7Eb1h7tpMeDIgFbJlcrP8LrGXmDjP4FtLhQ
4hJuVvrY63pDAuVtNzAHnY0GYIdL/44RroecXoltJ5yQZqoMn1SxWEG7Ci2h2QkU
nHANp/3L7WmoAgbt8ILikBVup3CRgABZQcoHsTSye+J0Umsbe8HQMk85WSF4MyGc
HP7eg/kzykMCxykoi9gZQ+JHRWvfVlBhfUm826s2lvwwo5SM7GVaR/lc4kAhHHgY
7tZFFgZOqG/Qv8+06lUVu0GqzC4/OV0mwcxU9Qx/c5iUGFdiaGALEgALzNu5Yei7
DnbRY87pVpoDD57b7zYHoV3wzH79byyG8HFuHYdSPfvXAjI3oljJwhyVIRnB9sel
0wGs4vsqwtaNwgdv/hePeZitvo2wv4ANoXFwEabaF4V4kz2URPUETTPl1r4GwY8+
Be8D+N7N59LqxKohaTZQzo8ol9VbEFFPXSCJ/YJnJOpYMBOSiJ4frYx3Yh76LSHN
2ARgvjF+snFaM/Ih9Vzrj/V6pdwu3kWC/aqYgRmGJqDAVTn3+5jnZK8mcqw24Db5
M883Rz2U3wONCYszaVu7kwO1XHNeluCzcjKpxUQZifTgvz5lajx6zNbx0iCnvaW9
ce5V2mvNaMsJWffnJU+IjYjaoVwPSS18V+lI430fnmryY2B08k6QhsZ0NZD8gmWF
hfQ8FsWKPIGGCi8AJpBnJ4M6MC5dsMUBpwHM/QZ59SvBJZ5IeRZJLnZBvAmpWmgG
8iO6OvkZ8s9W7dzrgt1zthi4n5JOqS3Ebas2hKUxfmJwL8Nza3NzQttpBS4o6ASS
YmqV9yV/opxqCAtfhv4Z6KGjvmp2ekIiWB+KIKAJhTGZjxwK0uJWHuxdsVBb3tMD
55/1Wdgv0uoMurQmZxNPG2dadv57pPixu8tGxQFMzebsLGbPuTxp13+neSIwVaA9
yOdjw6R/Q41ZIfrV2xBVfN0+FO8HuvGIXEpGZK+mA834Jp8txfcftJcA8s/7GICa
l/KgDZ06tfMrn/ZcVdZQjMg/dO3F+N7WdWBR5VlNOkMipaNs3PufacIEcVcSKbpe
/aXg4L52ygufpIlqnmZIe0wgo9I+ApsReFwRrHEksGYggye7kW4jmTGJrAjS8RGB
W2t9/TR1FxVHVL3obWMly6FwpcFBk7eDbThrc1Zav+KS6XIaaihRlYOq1qBRjVcy
j+A/eyZ7Thtt0nFzGg1GKtZBwwiikIxVoD6aFpyaGTOIDKOuF7MCwURuLwSFM+Ay
7qEesmPkr+yii0nxmpxL7iPItNKlwf+3mU1eClNr2j5aV+ikaz788R75lgjY+qET
G271HNNCpoA/o2STH3dBmgukl9sUR5nDnXagjybNJ5epWy15lZBvcibHvYpE3IaU
sjAxJxKnYXNalksFDPTA9AWsbuo2vz6sJ8uAgmBKFCkffstXIp7OhufTbrVH9MvF
IHDn013l2gyaKsPM/sb6SWFXXIumEOVw2pm3/yYfCgcPdLBsSkYsG2yT10kDsoik
sqqifP7Wina0Bu4/H9dgO27XR2Mv3wLnpnnMBpCQ8ISRVnjr+9oVicOxz84LW9tK
GqeONlwdwXXrGvMvX+IO3I9K2gho4KTl4XfC3PwHRIIsAJtDpcRVZFtMKSo/5OA/
JNZaZJQGJYKztmHXmiS3wYZM97CtKTSRRrgyjeM1WGY9SiwDzQ2EM8o0SpAYPiKs
wAgUU1O3It0aB87nCLn+hhFrD+5VMBBTBe/dg7VVeioKHnrrJKyWSlyAec/ZaN7v
sABJQUDyeC/kBtgT31SpZ+xMmCbkHR1Hfm2PGr9Hp94tDED3KvyZfB2x9GpRDsHe
dCCQXdd0CQ8jym8oQkQv9VrZqhkEViTaqOb8mkonXkE7jZ3t0UWYGZuunIQwu++u
jnx/Ns49Vfhm+vT+eun2rbl/WQcf+xaDLoeN/1eVObfHMmzzo9bCzBIW9AKp/wJ8
x4aLl0gNH91xGtIarQ00ztOM4p/g+0il2lmMy35vNj4Hx41NaZh87PaVFq9j+CTC
3P34PRBZkZFajH1Za3UBEwl06Mn6uPliitERI9LnK58DSI9Aasfo63E1aEJrQHZ7
3sm3+NRAF/bZYm6pfVEgK3Fs2CQu0cNxWN1w+wLEvCctScUR4oeBH2Adqy9UmDee
sDNWIWLgmkUrnR7DTLuY4c0GX0yb9Cx8cfLv7kR5jQGIhYqbQLGX7ibCyLNgr7OY
maqpYVXPLmGvhcFiP0WDyY1DC8L8qgfkqa54JBKSE/9mH9BWwmYO6/wCaES4eu8X
wLCO4c/WnkKBuxSy5l/j3E3oefgOkHTOikXL/uCgybkt6yGU1DkSoodtvI00CwMI
sY+L4awhFz4GBhIcobamTtPr0j6Tot/n9CiGwY1COQJVZv6/O5i2n+SreBCjvx0G
h6Uk2HvStixfwjBC6zeDVdggtEi4Ef0Xwz4HZFaJ5AwbxIdX106vYdgQnPnRFh2+
xgNnxoL3KZSTrTxxpDWOFSlGu8zcasRUphVTazUF3K/llf6l8vV9TTRmuBldOseT
XeYYbUf0BcP5UrdzT82IfAA3eEHIGCo3Hgk7PWhtUgocSpLQmX2Zc51XuQKsong6
7DdP4BeF8Sq5O4IVa5260AvpBe3+j5WUox6Ry/2kWWCePGG+H1to52u/NQ+dGDwX
hj/woOvEtfp1jqq1jnTKduUtcZgXkd3XkC9aJ1AJ2WEZ6EfbWmvv5Ods767zEfpm
qLNQ/5f3XghRqThGeblM6e8a1DGF1bMHa42T08WIgxclYaJerOtNi5OZKzQ0x5GC
P4TnqTsQ82IOjROv7zb+ImJnqu2wikxmH8YxUpPeoPKBXwMImYOOdG3KjU16ooSg
zwwGEQu6hxMd8gB+i/+dAuVkoqIfTYP2V7m5HjPtOrWtsAwwb6AX8Nv45AM+v0P3
BP3goUYF1prOpiEPzEVSxFI3PSWUyeE0drls/4hdoMHkD1xEu9yA/D4v0srkybN3
pXmPSReisem+CQsQiooXqLCVSAWSf7yDkuAcAzCyTw99z9EDD2uWfx2gWB5tSy2X
NNc6a3nsEbVk2E7l4oF75Q0YV/c/5e4fmha8sDST75jGWZhywxehbu/KTh4lhy9a
/CwIa81e2R6dERvvrGUrIAR+sPLHM2y14dGlX8tK9l36d+6dMWXDpcZ+F8dV3CwS
m5cV0R4RQW0gku6kq6BbOEF+2N7IaEqqiHnKwgLDoGkZTNqdCzwlDOHpYtwwykK3
6CQYUC+iCOilXRNHh0e2G4s7PX90bO+iH4anemqVNsYuicom5CTTT0tp12c4fx8H
djf9OjFORBu9vBHb0M0efL/ff3aqSrzzpNBcqsZqWs69cgzrsmh+iz3PocIAlY0E
lcdxkQfHvZqv6RnBl1GbJoTzOTI4RvRtSOpZVWKZv3wqu24x6mPGUhqgpKtoMrGQ
CVproXrQjZXvvP45MP4q5hdSjllw10Vf6u5MR1qNusU25fctGOJTmArZvOxjqn9M
Xt0h249ZYij0i6JSB1VqB8agjnMy6nEe+Yw+JXENCrAH4BMmiz7CHNLCZwRqHFvY
SXpSD+z10x3B8bsc1JiubMDcXNB0VeS2xRbf1l1zBxbgHEcLuPXm+tVEiF3HLAql
VnhXsjk9u2Ch6zBASY2lanyud0wIytSVjtmus6FEJ84dT3UKtCCKBRGWpbR/IWdW
rUeIx6D7Nzg1qMjgSokrFzEaGA9DiGGU4AXo2dI4fnYMOXFmt8ZZZhh2shXlrMLJ
Fe7y1dhGrrh6gWfPEVU4yymigBc/gpGQUZWsOsMCiXLy4711vVCTsE5S5Hmas6ml
lpsuFEiZe2VHO4MvZYoz0Hc2fEYNG8lKJ19X5wG9Zbe6VFd1/IdtgvidHIKK+yAa
FXHAm0Y0WSa0ks5ALWnkFbqaLLtjAw9h2tS0Q6QLShf60vtKzT4hm5ompRI0tnsC
IVgCiu6X+q8A7aHf1Dsa8ExzZThozGG1Ze7DFczsCcwcakbEMKBXuCJmTkXUX9D7
QGVQQcpEzaPIr2cb3JmMJnh2Xj/CNtb6NL+k44qpkfSwAa6UViBGUxiez/BoOilb
7W5iJyQFAJYC/ZH77zKQZT1DikykKvJjUxnSQryDFIH9Gs4ciIQ15hJ0tZ8AKgay
L3zZTAXDtZSiFNaKYuanB/vG0nnR67GNsOGV9Re7tNKHV4+zKOsTQ/U5PSYHnJCM
3gRwHgxotpZ2iSdXc3iUe6N2nIZeU8pnVRccuQ9dLKHbVNefVkdkNmrK0/1K3iws
2ROK1FaVI7r15417+2zsoyEIjMBRZQc0epcQd5PqKj+ExQTLe6sVysZCKn7cjDFJ
Kg7K+G0aEYxhUhXfKYMnshJAIdOcMf7WcBICgcksTXGEm51hheKqeuYX4eSOAV4e
oLPHHBD84stFyA5nXLfnE+D/+flxki+f5rYd1dBBQb/GS5rmvvq557mPV5I7p9Ap
irL0+iTY/0uwYQuuxdp9RXTRY1vnSN4OgYnETFy3Tc23xMcPu2t4KjGNvU6DjOpv
aFrIZ2S1kZjGD3yPnnWAHhFjZsCW0gHkkbmRg4qg3nwa4SXIeJPgp61y5TjOpI3f
sA9mCplToeodaoEfOMRVLxfXiuun61yuOGWZf5F4ju+epCtNHmAVbmxrKalpGhXS
1lALqnXZoel5BN8zhDGhmZq7rHTDpxCNhnwjL64iBq97Rm1tyibImZxxWNBRM2nW
JcbKOo5UssS+vWF4OBPWzdE0AL1q6gUqkUi6Ina4cAUAAWQmgMBXcLLDBMdDK1on
mUnI9gREJ3vRaKRCzJFTTvEcmTZC72+CxvFUeoUCSu8R3jfHDS8PAv7Qi1gsyY6W
THEZmDS7q3k9O914LLNDeSzs0GBSvle59922VM/+5DsXvK9h04AQIILVIyx8157N
jL4uWnp42VdoEKRLIdiD7mjgLjucMPZa8EKnmLw+vx4WZ5D/ggELz9xW0FMkt4nn
/eIHpQfMvBAqD7QMm2a6pUn5kJeSTF5qHg5jswTk1vQY9poWRnPemSAZ0Az4lDyI
Z+95lWqIGLAvE9vE1eDekQFsLZWQ+YUALAXQA/10paja8uJiMEhL0ZR+/zwU+Dv+
Fc1dA35yIiJctCw3u3JTlSyAgcDStv5YoqllfcwcfsMtAq+e1HRZm0YUYHkoOsrj
eGiv9ZAolZ7+J9PmO/j0I+3yEaqzvfh4+gxxvcumnSFW+Nz3c59VyOD7OQK5sYJs
iLDv2E+cuLSpsnE6Sa+ffCsUM4bHHxoGAqwksuaAVflIlIw3mqFaNoBLKUQV+x1E
S+RATlIe64JvejKFBuav9crzVs1lDR1vq2jIJTBAmba/9NTrCra5o4a6MNWiH/RS
Gg3UQv94/eVbD9ekjIcJpn0TgaP2Q54j27nCTyD0jGKABXTnvuI//qq4JWpafN6O
9JtMJsmJP/bPsY4KSIFq3D1DlSYoX0LoS71eBL77IvAY4LLv16lpW1xgsmzpoEsx
+mb48E5wFCeF6zJs+vuKCJh+kE6Ajlabl+VjsEvr+A5O5wSPmRHEHsMhc3pm45SN
MU4UorMxl5/NXH73Xxtjj1e0mVdQbL8OSqTuuRMJVYa6UjNasva3lS4VSje1zM15
OIijt4Q7y8RC6BEEbXaocZO/Ujl+rwHdrEw9vfIGBK1wnwn2mla3krSzciUrP5p6
pkPIZlgb9ZsBRdd+xh/pgGJm9k9EjIgn+RnSbSnrCiDOgqWC1OzoBaOf+1fG9Q/M
yjQF5xxZTvinhoG1A4ZJENy+hXtW1tqvM7oJNC76GF5HiubEhLPmioUN8sgcUHcL
fL8GPOdBMYwFBGF0MzEgGTzisAHX7RyQReE8m2WcWkvTQp6oTr6yqik7hVL1axwx
QMP9ibt8Ncn0iBkMDqkDtcPEidLPhX/Ct6F+NQYzUxcV2NDsvkaGiII40zGtrHbV
dHUGnWWeHbQFi3SCKqBFdJfZdnPGR5ZRx/etCTQ9qU4JgjTarbCY7aJ8A2hQ6YNv
lILfYXmB8GbRO4Cw721ev1as1GUQJI42CNLsdU4Xj5KaSLCtHEuXTtbZDohJO2x7
7q9eeME3ETyuRrmUkGVCH+4sLxVqlxdqyiLbPVJFnf9cn+xQqfFzm8KjvSdfTNDC
ZoMfOf2TFxI5Att4gqUczzlbQLfz9KmQ6H/UeWiLBkAUwWkQfyP0UvZDpq7lLTJN
/ISZ797yv9NPbejFDdgOvoRdJ5nHUQRHNQzI0NyKzvdH5AQoRFIG3u/Th+41pYC9
UEK+1wuEvuMiF8sYZt7xKESLB9PIlkhtQE4yQ2wv41LsRCQPDDNmI+gFMihiLzEd
fv11Ya3wUaCljoNZ8m20BBSiZOwUA6AKiWv4Dw6wDA2tw2LHwprba4ZhXOk58kbv
fH2sotPP1Vm46k6qXjD1rv6wLRB4eQcaPznpPGK9M74HCAHoBmunYOilB27Zs/53
Bgc22ltqEn2J8Ie1QuY+RoYTmHc8DD/NDHgZpNoE6QvD4OiEeQDnrGBLQR2cHWn+
gdt0YReR64YpghddH8ddJr8iaPVlAKVTKj1QLaHWFO/lkgE0/uYNIWocYb8z2aM7
QcDWz7XbAgs8pK3X+oyNoKoCB4EBE5oUtzulS/0Gvz0O7QGnShV7MvDVeX87lxvw
ZFOyzb0SPEVJ647K21F8LRaiZEQtuiJhq55mrD2yDpuqq8+jOxD+HtYeJ6y5u8uf
e+/eRLON72Js2+nNJP8uuHIBt/RjKlEXqA9+kKQzIUVmHYl7Ez2y1e2JxUZWEf6E
iTIq6jm27DUW7YcO4BELgftkYezXbD6EqK2TtPPl5/osiDyqpw9QMNIBLF9xYVnq
qOKxpi3+971cbf5G0cxLSMYZhesmnb/9IjvWywZWldJsJfIyGBwFfFQVsIdllbs6
HVI1xpgxxGf4ssaAEynHpSG+P1aRND94r0ZZj4kW0Ty53totLXEwVooCtaa7Hzq/
+4Aw6POrz+wKbB6QNFbUWyDPTW8pEEaKmE3vnGW1G1u4D6rEV3TOKXKEZ5M44Kep
a6oRj0P5uV6IY0XZOefF+hrdibqFi0XO0P3qphMBu4rjoy1AR5oNiaHGKH1vnhHf
XITnlGVnJiZr7Iu134IOOO3Ghl2vTu5oarJ4HWQZho0lVRbo21xw7hZrCc3GcoLJ
kBWIWXLJpT8RAgPPhDbjZT1FjUWBcuOYNm0t0FusEEeCSoBHH9qhV+2iScCwxpJf
eSB+lGcAu1Aq/UU5uh+0YFRfSGHq5K3Lrl3HU52h1E2FU9QEe/W9Ll0fBr3pznRR
NhYLsJEEPbHIVi9SxuERVXxrUzXJeTdxOBKVoXxBrgiFw5RSWeg2KRLHPau06BvT
hEykYfKl3ZOIBmRPKw6v0wmIMoyhcVR0CBlgxaKXCPTL7/hJ1JNz4gkh0kXH7SUp
CFSkgRsJ+iYqVm7Nd/c40PKxluyKeLw93/M//STAvpwmNJ7ffUoVxubhLdBNoLsi
hsePRA8D8nP7DpaBYKLk4lyv0SJ3tW7gHZM3YPar717MfUFDrB+CV2xGnXFgmY/m
IKOX0xQT4FQ1/1v3P0JwcaEFT+1yYBTcSrknWXBKkBfooDGAL/N7I9VQTXl2L/qW
REja4gBa+MckSXERUDZC9ijCFhEhN7j0/ef/mbESXXZuSld76zncJqG5y8mrslqb
q7LkSPc2TH1L2CV8PkfOquO0ZS2AzKoPkuemk9zzgp+pUVSd/GMEOSlb/w+nLAzr
50ufTfTOIfrXVQAuFJu0wGjY3l97mGpAu3NTyKgiD9436equnnxsDAh5wEkZo8PS
VqZ3Ea27M7PE4/t3ZS3X9Pv52m+AlzbPObpDfiaamkDd457iYNLffLL/zut2DMYN
zQdTUPQJOFkc2rC1OF43ersG2R/h0O6OXPSQ82AEs/Lg/TylyS0POZmXdWQ4d9/S
zp/8PLxH/CJ/l8TD9Rbq0EIPcwGFsVWiJtu+b/YiG2VAsnjx97tz4qLsdAEFPAdm
UKhA2+tjNjf6d1wFMhtb3Qxzh7Iwj7YHSd4krb43wkIqdZUyTNR7FdKK9BHIL1qR
Wh/gyco0BUempQVhvzl6AR3kckyvW3my/iXiVotOeAUyQ/odGerPCvw3NOqnLsQM
Xi4FFYgD/ugsvhopjRpQOkmXhFQDZ2DkFGmLOEM/EzHU3zMSBMSUZIUDsZL9iHVc
s/8k77gmGM6s9pvU1aeuk+N4S1T9/9+kdfAgZ2neLyizvELaQFNScuusaUczNSwl
0co0wkkUansMTRqtwa6q6CtSrv/j8HygB9DoTAdjn+fPqclftfkwQo6MWpH4/JhH
wFbCAQ7K+dFILxp5USZ7LRbOvEpB8fc4wn/Lz9fIkATh5oZXoMh3LG2FJEhskT1v
HRfsCkNnBzTNPfsQG1gtUe7d2v3Mgsb3J5qpGhdgrSGj/Kf+QBop7PeCq0wfFrfn
mKgRQiMTaBocaLd6qQPm2IGyHyi6zNBirghg1Ttob9tUx7sjWetKkv3r305s5yOr
c/vAx0EkEfjm9B8AGg3yo+ZqJLY1S8QDD3IlO43Ubtda76s+3vEezOOwTvvKmdDO
0Gyn/0m+HAIJy9vJqpHcmcg++d41bwr1Msi3VW6LpCR5/3bMx2cF2pFd9SoKKUEL
DcphA0R+yUtjDUCM2BAR063M0YQ+7rTYyO02tZ3DiWbxmfkVq3JvTBsO4gVAMO0D
QAZM0YMMrGAeT8x/nqaWHywMu14WkiMUDAt4vnqcdK/jF/1HlFdbdKI4cnkcBnt+
aiHx310V8LB22MxLQeObZ7Y2W+ziz8OqvIZC0wcg1i5kGFotwjatcHogV2YgqUNd
ja2O16QC2dwT9Czd/rc/u0c+VheVq4R97A0VFyARkRDD2IR3WCKMM2mY6zQxN0MB
rwP3czB4C99PIuK4Xkglyj0dLL4Ash4Rv35hUmsggHK4S3z7GJfhjnYK1+zUNYsc
T59SLRyfX5MyWEnbBgfFmbsF7K97J6LmGCWHZwtRO/RxJtGQ3o/PwuNO/SvedtV4
XokJo7oxb1P457gsJgq35/yixRcQvBP1q5vGTXizs25KoNvntABN4+ExAepkmU7Z
cktPXRhXKaW59cJ52DwmymYpq5DwMHRf5+Ye7/3UwfwC2Ccbrwvai5OC5FCpw1Tn
TAOoHDSFzWoC/XRIY0h+hUbA1SOK/kRurWnxgK9hsU/rv9SWcENXOW8sL526+xu3
3M92hy9Cb/ZgG+o7WGBghvHB8+qUZXQVpURR/R6IIsx9wnOqpelIUlZotTZlazZS
v5zpvlnsHVQ609xwqMx4L/Xcx5UtTznuulagxvThx4C092sN700OaEpIhNkeIGtD
m2EiAi3FxpSMR7czSYF1+5H5wkMPcszht2ksU0DlZhHQdzixBlwn4j46lINt86Ij
1ROIdlOkEwPdAnQHHqskCAhEF7bhsU3ox9GgWO5WbWP+EHMhV1xZMcRlyzce6ubL
/wZ2Wv6Mb5PluVDrT80drmC5hKClwqj9soyQeX88PiMf+RimE0Eh0etUDsNaFUfr
84WMeC++7FE2Ja5Au49b4RvdHz7SvQPCPbKN6m3lZvUPtUlfpKJfDsVZIgP7rssq
d2rC9NH+wn1/TxOdR2HU7srZGjfaoBPGO31fViRkHSP3zF1TW4fdOurq5Y8aBYIU
kLoCttk56kzMiOt/+03Uc6UZpdO7PAllY5v3v898d+cmea/9AoQJ7USaZIA+W779
VZAZNxuZlA6NE+4rn4BDF7nZopiAL1GY64rIcwmNiYj7CBa7gTvx5qwYZZSFBMs2
6xWr+hFi5D4ol/tckJ5TS0N/1r9Dem/ubOJyemNYWTx1UOnMKzrpaMaHVQpOq97L
M6j9QIvPUwns+QSraVmOnf65/pLAGicka29KQTzonqIBRlYWmVZXIM2MKxj2Fh4n
OmeQNf8kVWZ6elMmxmOfgaBrHINHITSFiUcTJ28rfO55z4Z8DGXzb+4xh3NOvF90
qUpH4teqIbZmdFGl/W8NG/1V/7/Cam5cg0Vq++UC9O71hhoKEL+dOeuU4PO8beh/
0aAyZJ453dZHl5iRkGTgLfPgPZK5VaI7L0A93n5YScMarhXN88ULaMgZBB3vrwjH
vZl5uXKAYsp90nSGMICTx0wYOflYUBroNjrI3eEgLjkp1x/n327ZdM5CDSrBAXr1
pdu1OjVlMR3spPofsuriLPy8odIgq7Aie+tMeK4R5VJpicokX2w9cGDkNXMVG7bR
wMFG8eYC/GaudCC61tnIEsFpIu79PhQncWjs2mRaY6E2WKd48JZk8vL9eCt3rQvM
/C69WhRdLSGt3tx3eqcFCvXkfy+Ly69j+24n28dMtyG3EbFx3T8+EcASXOGEV5xq
VO51qmJp3d/uhAKyetNx31kBYOfBtrNdfJIksutD8Wzyktp5Cw0mRb7xzNT+hXdC
J9OdC92VKKWSoLe/+CVtCZDeO+JlLMPUnznVdLbaPk20+jhzNSEcp/sOsBORfG4c
OvCitKAkQLlzgyd413An6K/1VGs3rDd9jjMGLr+BJhUOfCmLblAZDgXg8i43CxkH
T1d18rEBz/Fy0muhRn/sfi3q4bdmJnaQnAJjTBOshQjWb2IYPDmP+ypIQC92yYzG
QJBguD/1W83/zNhM3cawNMSnf+GbB12nqYMHZdnrvdoGXhCPjLFbBaqP1w4bANMW
18zbKllcAbc5/w0O3FfB/WmC7Ndf3JupTVSb1kmgXaAQH8b9jrJ83au9WsI6ADgd
uy/wJ/qnZphDXIxnT5T/6HkFI/BRLMx81FKTF9mbTM7GlSIkYQTNnc8zCBkFg4vi
sMVfBxgvU1na6xxiaJEOaEG3x//4bllbdNBHtrDfdClZmx3ON0Wd6+Cvlqc5sHtK
zTPkc6uXbPlgo2R+xY8kuP8f17rvHJAM9YcjQdzEzvMJzvrK2CDbtIgOJ7G/Yh6x
dXGijYMwknFl9yIFYi1Gh3O4dDSi4V264Qo8G6+itVXrQt25ANn7vAgOKqLBXUGv
JQKquLmQi//8Rt2k+xRMra2GTmXQDF6eBAWGYk0i8xNsevJ2cmaYQJ4I7hDSDq+V
7t3iXr2IAKBDpQhLwk+HbUVvFZ4PwHF+72HbCrjt6VS+6ox9JxNaUmacH9gh/XSo
uupTQExrijk8r4y7den/YkPKUYhh1AWlkwtovz6ygeCwONq8oTxGAn+hdIGO1tuV
MMPd3kOe/kDpiMnS8NNHfPVbnzy49Ds/wF/6zg5jbA9LfpadG4jQwbGYwTOWGxfm
uL5XTNQk3rKtC1GcsqA9grWJScNkxP9Tb9h9mTmfgV8hTZVUPKTOK/vv4CMTzFC+
MMC8O3VpWamUpi5h/avG2JACjbePP4XB5ATCvVNtqhwIq5ECZwkKbWPurGNAzYrY
kmj/qW29rpYqbR6+Zhx37Sky/GI0cujP65tSkyQgnkgky9imRwXSWXe9nnCOf19T
ToIRKRYm45+NTJFO24ZPfXtKzM69y/N/47L6WBM/g2iYu5c+qFZ9BfzW5vXljnc8
0MtYLWit3L7sa6gWcwDiWu2veE/IOI+EVHQ9PRrQgmyZFiEduObKxOdHmIzlcLG7
rP176q4EVXEto8Rp99/1QG8N9o4UidoJjDeh0uNenswuimOPU6V286KrOkspo78o
nrcOPqXNmZ6E9wWBGfHFkfJyZlLvE6n5UXttT0xTGe8bQ7ej8NNqscTmLDvPLcYm
JYOqM+UPE4ekEMhuskE+4VGETF1uMmNlFg2N5tGcyQ5h9aVxXupgFwqySUUrdN6J
jyzfF9iNBPttY5Q486Yjb2ZRmp6Ws32uLuxKBGg+51ySWvHWWiy2WUQj7QVV1/bN
A73jWtRn3n8Z5orMWxo3l07XSkAGvbK6DFq+WlR37ol/ZFMw0s5xyr/95C9T6SdW
gLQ3zLKXIbQjEKTgf3VZj/hIg83mu4tuBU/mI8psT0lXe0gq1iFkSCDwCYjw0xTN
nJHYB+fXolakno3b4uVuJq/9iU42YF9SQ6jvKE4muKLRni47JC1UNNQAXoEgONQb
B/6J/R6jQY7kxS5+LJcNOs7G4uvrERJQzMMX0OZKJRhZL+xJIgdJ5/u4KnF4PSrH
x2W/fLPmQaWGpjY4Gn4s+SYEs9hWJaMbbxbBJCGNrLAd/K4UMq6VP/7OUKbsGWW4
V9xfrJdAILTXGLU5xFfkD6qPzAUZYhBPBEkjynOEdBCnpKR0d2QHf08QwSt33NVE
vJTwcWB8e3Nw8vQt+0njutG0TRyGHL1bl4Aqq4PiMHy678NEammX5/4t1XpHb63X
a9jHsBA6FWD2ftGEqLUXSuzsZrb58HnHmdBA32B9/uROQSN4mOW9WQVLQ7v5L1lB
xjYIV/3DTWxwBCR4BQI5/ywUo+Nah+J0g4sjbnT4Tbmbd6dWTDAc25xIsULgN8oG
8T3JlVsTi/vrg8P2/rHJuyGU9yDiPTzuR1PYXBKYU0I78/byLjO3DFmjuVwPh/QQ
X851DJzY5+L5u7cs0Y1wqyAxfTbkl+c6aVyS7O2T+LFNjXtNf+h8fxvmbgKUdmBb
tEbY2X9VXA/VJMzTOj8EQtZPk84cq2Chv6rK0B0sejJhNerXvpcNnvJm7r29X+fH
IgVaeFu+4lubeQeLFnHZHeOvStmk5QI7qF3fhN0zt1xrcU6iHETvts09v+2W2apa
nm2Nv2etVe2UVcBhj6hSy4SlngcV6MbHWwvSMag4uHzXnsX5zXhkc+Kz1J2nwVuv
vdO9GKQLq2dBiHrI8kBM9OC232LE+AkP1f2DjkBCe1xGQ49Fc4oFAGfqdjql74r9
fdbyxYe/OKZ4fvFFL21X6QNFcPbJlHE9M0BzUsh7zkTqBEz5rt144Tt7ESDxzDch
y9hrUSm0BVU4n2TquTEczIiFlUFJZ/Bi5RooslZGdXkl71od0LWsU1WrJv7XSapf
i4nBGse3pCgMUNd/HlMCZd+K3anAiJsELcI9Fwfn1HU9wgSvCqLBK4ZunFPL4Gt6
6tYweWVEmHHTJgsMi+at+dM4p+1k2uFwl2c1F4OJkSoGKw60Wy7lVCFLqdErcw1W
Zo34blmjCawD0TE4j07ISUaJY8KxxvQHOkxJpx8Bxqp7Ew9o4MwMB2y9sWjqmQSM
VjUu8D9xAWVDBZtzToUKQULs2sUIbK3Nq/eheFOCpAzgueIYVhQECQCjKZKqGfXr
aWL8xq8iJZqLQuI+qjDy5hQafGv2si/nIXxptov8fd1SAV09a2UoFmob+8NFoOJZ
jNiKNVCLf9rQjsqWkJcEG7sF8iQ1ZYPbfjjAWyALJgYfTZIsBInWKN8rRSByb3d4
RZOWin5+gzHscfu8vFze4k70O4Nz2LyGXnYYgaZwWitsBp9miXThcFfdafvXsQW7
yWEL/orFdTCnVupQx5SmC9+JD2KTJ6Htw1mJxdCzwzdfelNsoLdnUhAqnO5Tn+uY
LQmN0wRINJjUES3mT3eBDhlSUAzyNhoUHkFv+iKsdtP6qBfSDhaw6Bmv68psEJbD
9Z9qPHuHL1tm5oyNVxRAdmnqzMsqwzB9rhVjxZFEyktH5YkIMAqaIghxjEuPinyU
EaVsPHyDjEdWjo0LL1YGaiZ5WrLfqV+kes+e2fHYKvOgXbQHfLXHBOpdD6/NEPgd
qeRYIw8ggVs17qzZqrKCe6fcSW2kfbNqb+5IsiDGquV6jx16JHUMkYrmwfoeIcqV
gbj3y3kgc2aimiyC8qSSnftwLXe42wzdX2sHC1HRfJ1bi11i6Swr0SNWOkIfim1j
vgYSOi5T0kQF/tbTdfcIiIEHY5fFz2mBAWTgYiE3Wehd4F7/EM4A84rjuLErD3m3
WCrxf6i1drBlsuKS7WaWbogUaCcQdljrymV+aDnmQs+Yh+QedQMCykq+zH7MJSnt
aieyquUFsU6lmMfNrZIa0lv8tpRGXjcCjrJFOOXJiVAUcObYv7zTZaQCNkcH0baS
Ly1JJ9oG3otLxs0zo07rewcUXF04j1GkmOaaD55iWrMZrHBZBq4LYIkW+maBvnA6
uJvAbF3W4qZDgpqL8f8GPgVXxZGUr1BmqF/EGTUkpefHsjZmzI2t4SCsGOnjPmgu
kLY3Ijz0E9+f7PysZOlhsvCjQPP6RRnmCWc/zueOWL2N0rnDTdeUHto3dJLkbwsk
4Lrx9jvaQGuUISfkq9x/5xkTwk5Ml+mCWrFJaFuqrL9ROpzgyJZf/RIyPfBgrd1l
QmjNdjNVpQkeb15WD5LsjsdMws3z2NGY/UdegKO0LKH2fOuhJ2fSlxd7Hy0gr7BZ
+7QxErzZRbRcVk/ZMvYC6KqISyg/DgQ2C8wCM6W6H/6XzEzqjMjM8A3IOAC/FqWH
PFW0NI0nb7AEQxNv+mUC+MLGXo8xxuWNGRs9nOllJSbm4WWWg+ICW5FHBHEKPQUK
nixahpgdYVAycB0f+zfV167Uj0ZhBOZ3ufqdNTGe4SmUzL3bcSSDZLG0EuNw0M1v
ACKcAhU7niVga2annC8gKWx1R9Brt4CtWDvRS7xAF7qRzPmKj0TDuYBGHWP2LKz0
R994i/89M9fIINE7WQ+O4iclDRamB3hzhmY8M85Y2IGTuU/PSHGDGnNh13i2GWlP
+r8FTwAr1va6lGE3RLESFTDs2Foo6kc6HpRiVLEaMgbDEdJ+7tufEguXmka1LSDw
YS4ViazTVKqfJkuJynyZRHCrmJ5oreVgMCDeWsnsh/qQHZRooweNzQdujBQqoYrv
PGhIJsWUwPC1iY1/UtHjM21sQFQ5o8u5McjS2QMKaCvpvGmVvnI0qnTiQl5CzdqX
hm6qJAxCrglOVRQ7QE2ucMx11k3RVnGTj5ltD9VHmCApqd0bzbYOJD3wuqX5xks5
FfyDcX8aycIu/bCuQNhf80qnXUT28um1QYhWZRUO0PU4WS9+UfzTjy2xveoYwGJc
EKjmMtIfC7Rp9k3ynGO3/ZRP/dkdPemfimoA+w+DzU4q1dutV/ouP8r9iIpX7od1
dRjk8FVAlucQpvFg3uUugnnRBUbVylpyXKbpEaEjPD4Ky7J0HTqVfR8bS3gBmla3
Lmx3Up6YfWqDfFWSoFM3A4RlxW3JQ+lQ48TY1G783zuLHZh9WmokrLTy5652JYFo
HTVGZiMmJ7FC6OzISG1fT8MWVsLxkSRLmmz5k/aKVFO/JhEaWFAD5ZuECJ5ZbQrq
Jqs4apQPDziYSMWTTjQv0oNJqa1rsU3YSYZsFqbJzS6UUCxOzigI8hDtaPn+89dr
tSubf4uYKeAqlcQJwbUzgKK7suIyuukuuQRKKuFPaHX1V8O0NZwu8w7dG9/ApXK/
39OdmBft2Paun+FihcZ4/MlbNQh/510Edv6MKo80LMfMT7sg4WJvh1GJgSV3Oyn6
q+D2G7xdl0DorOLPf+W88K4j3Li3bibfDnhQgMjcw7BUzO5F/ml2UZ2pMVo7Xs/C
VxkqIdqUE5/0g1F7K97r4OmPVe5QGNOO6YhBrFmvvL3DuhGn03iGVsOHfBm4sNjM
kAw8UoDYGW570BkgAMndPkOaP69stDXNYF9DwB7fwh/O6Z90oZCJCQ5Q5vifAqPO
+AWSdQeukUpK8PvCuD7ApD3vuuUIc+nX5eKNn7iZPQ3+t77SQl67msDM/yOu9ASI
TM3Daa3hA0MArQCKS2oa5ew073+oI27gWvogMvd35g+1hd6zbkquAMVpCf/LvSMp
W6Xf/3TNjgojZRaJyyO06OjvMCQU9Rrmst6ecynwGHWtCStg73Uf/LCcQXUnx4NV
C+MoLpWAovwyqfjksp8MsQXBonlaE5tckf5g4vxfXXw6xehuyvMSCM0xu8RboNoW
bpPmOcw84Dc8+z3YfMIBK9+tviNqhbMVIukZMJHP/oVTFFkKCkRCWyLgsWvm0wTL
BDYCwHp+0p+SZ78J9+VlkcC5Wv9c62a6gYnmZGria8rD6y4lt8lnEMOfNvL8YxLI
8MHBN/D5jQaMkNxxZTZPkjKTXdX0FNA5aoOcLsWUJ4dW8ELJV8R3LmGwoFLGOyws
DiaZuMAO8G6jdqabxNi+BsVBajo7VI4JkN6zdIzoKbmOsnAdDjYh8dILPmEiKGDD
57OGRnWkhYo44W8P92QNY8h1TDypAT+DksuM5Db23BeWAbVJwhRsiN4mkJ9jL+1b
WHLE3sG+CF3Ynb6mE87mr0lg808NLEl6vvbhFzMVDlJQIiOifX/e4WEy8Jdrcnir
5A59+Jx2nV8WYG/hl9yVvT+9AYPBUv5vO4eXmEox0By5hln7Xbog+1QRAqgoNt8P
VeeRc16xqYkVyQeYjFdhKKPKUmu/nyYk3+FdsFJK4LgqzMzNxPGJtTyvtzTtzv9I
QohfD4ExDdBvsmzU9g+x5fh9ZfMJTknR1N6E8+3jlPnzRaIzMsmRatF/twNS2QRy
7Sc2HXdyt0cEDdSZOlfzIjHIZ3IqQ7vZ9fVb72QHELro/V61h8AovRedIuKdE2ax
R7VVlExUaxFjRfUFjEx/SSc3ZsP1PWL9093ZGY2N9UJPKKG+fFnwa9ktDbuU2MfG
gqf1Ck8h8P08cm1kmQgLRatV70bVD5nfRHM0bxRUFZ7Dpztj336mwchb5bQUxV6j
MBprkwT8sJUFVMTzfbUA969VCnTl1JdOe56X84Xde53dGdaMMuonm/3gNvSiwy30
l+iwRmdWnMMHPUk9rysPCPjTP0XQysbeeOFnPEYN/IvXAc4iPb/wsegj/u+r+0cL
8eJzYAfahbISl4Yp7GOQy51eIz+JLfLdb+tPRkRfMyF2pWbtgcAm2ukdxlB+gN2X
9KkJipdHUL08dCbDQ+68mFULEDrAQxZ4LVYElHhI5F5SCU3Ug1h8TomPJln+uKxW
eXoYifA2c5tpGPgPpOsDnyKU5Xg1539icFVSbQLUBMSJkdDgP+RKeC0He81ko0ga
dlohYnhGWg5ebgSXhCAvNx69JooEGXG4MeS0UEEjn73YSrJ1gafQyiwHKRFpEfXl
tUzf+l1qkKi8idA29842U174ortK4yCi1J3mLVvCmGNo21JfCH5gg7U38YVP7j9K
wTbBZfi8ZMkLQSbC1UIKNMWK5qylV6nto23VUAlhqE4o0bXhvkrDxYljBfZ5gZ8b
HmLORfy0aQhQBo6xYEy5gLOGCoaF6VCt9Y8xjPS9yV49kFUHSTZuvfK9HwV1HeVi
SdU7iZwnMDjgp5fxUUSD2OzrlWGBfKdKlEgXIBbKWHu9VIfVpolScu/JxYzl0SVV
tc85VI109CYrsVftSlqDFq1lvUM+z6+wmSrMAXlkczEY/hH4+C/Cx9h12eRBt41Z
2aXGvhZz7p5gE/CiHcrMR4I1nI0bDzhlUk4G5pCXhIuL9oS0lIU7iXt1lM6BfhXm
2bO5MggPPVQmiy8/3K9I7O4evmH7RaiiTLypfJBcGXEd3xoagp0fk31V8oPQ0I3Z
TZ/jeWZ+hT6a8Y5m0fJJI8JA+GgebUqepvkf8EQgwc9JH31ArKz/Oqv60NTUGFbk
MDYSpa5E/YY9ZxIJY2Teye+n7fq9u3nBg8H7tPAm/r1rifZtJrXgVhh4nFcJEeGu
wICeGqns5Fy/FvUuX5dPktugFuMeXVTlkJfP9zdXNoMGUexPHMLEuVLbM9sghdTP
q6QdAVaAD7c24jaC86YbVL6yTv64E197GsLKy0txJHG62F7GBs16b7aUU4UlCPrl
UkD1wXDChZkrfbgUU0HwWv+hK9mmBnY1c8kD1AIK0W7WGLqcDgiReLWE/pMmtWG5
eo8jAPoROTYalQ6jDFVKc8kMHO0zYp3CoIVUmRA0nRojI0N/6u3QSVpHIjxUxCyh
7uizEVLJsXzXncEYL8/t1Cv0PhdbiKYhfyt7PApMND+oMYGleaCIPxB3ZqjrrSdZ
yWJBXxSbbYGpJGHhvnDzBrZI6meJsZo1rR7rw+ouB7O1Gu7K49TmkjDd3IaOIaV/
Rci0/aZFZOd1Z61Tijkdt0vwH5IRYAq+9fFZMozWBpyV2ay1qVqBJfm62wT0dJmb
R26KRXT9bgUOw3EBCBb8PB7N9di9T42FEyxXn9Fu6TyBUALaps+QKfBjapFDiNIM
ap1Oa12e2L7MNMmiRp4L+L2R1jG2jj6+XOUvFdsNwYhC5MxBw5IEOEdoCJMXItZG
GRQN/ncgc3s+IFJT13oHnZxJgWJPDNnzge1Y+FSIKHQo/GXaTgp/EKM68VpZ46di
abWus9dNxDw6A3IgeP2HF6xRqIyWvWsuSuO4Ok5Fpd1+4YH4Ff3bGfGq8ssjY/zH
JEnMfQgYp1VaRU3XEOuzv+GbVlybThxry1jVaHv6k9xWPJh0suu61rLjnd7fCG+4
Z9Vnoli6NeWQY97YAX7rDpFjI1TEj58rAPb2ZYviFVgX1l20U66A1Qn2T4OEzZIl
NHGAxU8TOTyq9NwYZJvr8O3QEfHfwRxMKHqT6CxTf1R7DDG3CPpLrsBdHtl6shuT
PCwHTZ/s4Tc4jCaMS/+FxnCeyqevqixWgNnsRxxEJXhR1ax6A1DxfXuC/YgJjtXi
0TZ7ZiiNMXrxo4cZVBcFEhYVhD7VXXnnY0U8OVZktViu4tWAwqWEF/DthbKBr26Y
sbfJX/8kVl/+qkUvYvRomimP9gA5g32n632ysNAUjKYiAWaQdwOUHrens/tfcC9d
VbEZgDi6l67D0hmwYxCBRNNYrGW/G49iuZ6R9M1xyFV5hKJlPQ9LvUdBIKUVU6ds
cpZLBfItwOuCeVMIPYejLERXvDUPc9hZzPlmlo9ppDV8XHK2MErhJi+LRZnE9hQQ
zUnfWM72X3XYOJWPi1WygvlzRny5RyPyWbJALItFKO59gOjFA527GRX9dit5d+2+
lDjaoHQs2HJKBBqDi/TaBnJMW79K/ftdOSB5qVObdliH47bYkrungvrIpcbUdMe5
3WikbURvBFVb+8vp0puEXIY3uDpoU44a2pU2OutDP/QrhtgSHIBpBm1zE9PP/Y+d
i/eT3zPDFB+GPy3G9KtOIYXHjcGUADb11PXt/bKysRMRJHCutR4FSw2mQOomDU4h
d7vyXPxI0kkHnNiBjUrcf1IKfvklFE23dTCRtaXMoMLEpWGccJFJM+1IJLv7YcpF
ygum0WiabK/CFd2iCiwZcIDJ5RzU4Iw5hY6EQpzKr4y4iHfU4eVlmvBgvITmdkDc
UD2JIhBCT1Vi2PBv1+ZgNrfYCaV8f9MeO+Y8q9PkPHThKvO6yKkxrX56EpNFzqdt
ICCxV5XV9g7KlW1uLNVJS5nszNfrSPWmvG1zVLVIhos1ie76YFM4g3Ki9+KCxUIr
sTe3AR9qW/Jv7UBPgbDaIkbOPyAH/07aqq+eAQEprJSGKAOAm25FCmfVAOTitUOb
38dy5TC5Jcm3zcop9rzBTy4z3r2ao4/Nl+jL8OArwkR72Q/bbWGK+Ws22qWLtIoQ
MqM+7U5kRKH/BRYQu/tZjMDrWuGjvUyVS+LmtSMxfXiF9v+Bhl7o/AyFs/ZGu9Ki
Zmz9W4RDmelQVz9qZDqC4oPshLmwnwkZtWVzaI4OSDdEAjMwyEGFCP005YAetRyD
wT4MxLYchZDvzykLQKS4q+Ws2YBAjdBb9r9Vw+o/4INSWvrAzTTczMiyCUEj6wTQ
QcxGPX6J8OXsQiP7yp1wGXBSYOaz/iSWm9l77ra2svIq8JVjXs8k6EStXtnq94Z6
1T5UrzxSmu/w7SO2M018cua+e0sCOMEtzN/RH0iqDgpIMFvKgPAcT9wACRTL5DLz
UkB4dGGTCOr/YePDT2Y1cVVXah9UEcTrsECTbBG3UoAavRv9Hrbf4lf8Czonm0Zn
UuvH3boRiG5GunzNJSQxV4KMghqq8yUeSv2QHBHXSCYcJ8wyy/SV7Ezo/jgdrThQ
OarzQl/9aXqjaP7ylQchGGcK1nabSrIils2M9tzYgHtXdR9idgm2Y+CUuSZgSaOT
cuFVgscDeHgydJvkFXigNrDJLXXCWQKRIx0abvNYOxpslUaIuz7fFGrMHO9c+o5U
ro+1WTxUM4vyRigpLvrbG4g7bdBCvILE+tCQwRK95e43XgLxt5yTzs/ry5ebdglO
dXaHlYkTROo1/jzucOCrQpvNPtGJU2B6rFH6DVd8ZOh3H47qRzcEzEZ9ux37/zP4
0VulHhib/9rHuNDqIgDsMol7vDoptN1rIct3eES/VqMs6w3tO/zyNoei1Q5j3A8p
Q/r6Ku4fABC0eJGkTyy8xhdFdWNyE+pP6g+VOsew+gK4/+kY1HcwKhV04/otrsb6
suGo5fEThoRLJrSYVvP632FoGZ3IjSvD8xSFLDZDxgFR4sZ93lXkFweC8MTjfzh/
Cy/LKhzaDsm1sRbmBxZjrTtrDFtHaahYSwClQCmSK6JlkV3CEQKt5A4aP0emp4lj
rxSv2GQ0utTMgDkJbY0IxF41N8C4nDQ8MSGJf+Zp2Q+iJ1GmH7m7vP7txhz7lYLI
tvJs53TFUzBjCyvPDyrHH4VFD+4l+8JVrUjIrMz3iKdvOv2Qr2yU/9pMDSrxiKIx
Q15Ad87FggFVYIkQja8RIz62bvmIhhDuuGW9Z6zsEZwmp6ys4VH1MOJT4fr86cDK
D4k2SEO6Hha2XbVqOLTbwshfuWTT5iBH4vOdBls29wAp4CeMatJ/fOE42K9/KCYU
Q3hT45h6LudO5o1fdmC05Alx80np7b3s7cM4m8owfIKlG1dLMU4fvCCCRqx18aVd
bqKGak3XkkuLH+lSMtQ6k7LNCjZ3WPzQBauzndWQdDpVkAAj4JN2gZUsXfvP+bYS
w2XyQZt84Og5upBuZD2syORNSDmayjaWlzTgDHIwsfwUyWpROwJC3TEniDy91v8l
794m+Ss+Wh8fro7kpqHfp6iwv4S3Yra40+5TjuYARlAnOXaoWtadEe3MnzXXmM3U
p32nZZN3F3L7AkDGQBvBUvJWIv3zvLAQcemlynUcrEPu7fOiRR9vg/Cz6vA/Eme+
Jp2wOebLvXtiPegG6Uy02/0G2kVyVe8i/UXbpyWLeKDe3ou7ljYlDgw3kGSKS9rD
Wd1I6wm0fAaLDYecSLMJPGpvU9wIIkmm5dT/SK8Ob2zxZRxPsLrrP8G3yr9ZWE2+
kqOwRVfMaKpNhwzj3G+5Y9k0UsnO3MYEzjfIjIxGGPqhLnEJ0Prg7bgUQYuqLska
0d0h3EE0I1gzys1NL+AtgD2tCVzrxRtOh/1ARDGtgCeL+MC62t/qR2W7JxNkmKTb
Tjt/Qq3NXAkM0xHBzwfmtLcY2orskGL6tl0q8ZIRuO69fp4oHovrCQTYuUOTXDaO
AJCBXNlrDAJR8ifJNoGFh/Go0wWp51WnjHLkXBFSpU2kSxh+DJlc6yCddVF56D1r
DwSj/TyV0EtWQPCgv1t+NrfYylULFJwzX8nS959FKOV+6SD9f5u3PQ7GkS3bNRbO
Ibh+xAdg+GdT0UlmCLkWc8CYZvGJEm7+2cMRcwGdPqqdCF9rgkSmkP9NEKw7lQ8p
lsxjY6gNSgpAtIpG+ZW/xQgsK3j97FtABEpoO/0WOebpcFO82So1pTay24NzypQr
Bm6gC6uhT/W1c7JZPBaQpYquOd5XXBFWevoLQQbLTXBMeRwdWVe8JJBG3BaAr9+N
mdQyhXSj1K/X+MKsdcJvRASBbd32pyBm+/Loh9P85ashqkwVKaU4uicJ22WqTuw+
rmS5mvtfYQDHxkGRWIhNWKl6mfpRyZg10EtoRodYOSgMkT6smpQzhqk1OZ/DxwHy
l3ave72MANf1RcUlRPkxNl0WAfXVzLTWnCkDrqNR7XCiAhYLRF5YhzCVIkgzzDng
YrsiWavDNT4USMyfwzFdxbPzoSi6nYTClH3rSIzjL79WBLGmS8df0Ai0NY3PaUo/
V0EFrBFDgIqF9eudQ+fi2KbJhdNMRxvSFA3J1YYAIQ04YUhUd19tMyRDst0ISNUs
0ih0fNHoVnAk0K41iGLXpnlKpQPZRwfiiACEerbR4jBQ+b46+vIkDQh4CYw1E9MZ
aeSs/MWt9+McE8rQ99VKRp5FKtFktgLzVi1H4pwNrcq/Nfj/yU4sgwqMuK0nrB28
2sC20J/Awaw6mUuNGEBtV6P8UQCGw1S8veJ1aS0LhQrMTjuWFpYEP2ea+McPdvT3
y4G1ClYEjJcK3XW7luHuZ7M7TGpCE1cTGhZ4d4qiMH76wMkIiN0wxN3RojKkfYjv
b3mnNy+IJc/bmMjX8CjLb1qKWoKtMsmdIHH5CmNM6qeoChYnaYP812ZWkVDQ57o2
0IHPasFXz6QVyioABuzMZmR/eDaeDvUrraxNY56VRMRU007K4exgPvkTTc+Yv3QR
/vklA7UVz6pIS4OXsaqoownpXvL99JxIhJUnWFUawkbtPij1Ux0P4g+KI4y1ZG7w
rR5iJdtkRNK1tmSt4g8iBZhayXw9DsOAUI2/qFRjEmGnBi01CW/sB8PxTKyTM/JB
zFgIJ037IkctgF9WF/+296xhJY7Gfks//oTlRkyZTUohg7qyg3Z1SSTD2PgtN/dd
+HS/Z/BEFR10h+Wg2oHW1Tlu4Mt407S7NIi8O93WJoeXruOOLwJd5psjAiluvka6
gEULhFUyTAQhpSNse1UxdPVbbEnG/j94W6DYafAn9PRmv8cEYt2W8XtPxXzE7f/B
Fa69KqaQrw/GX4rIdigM5LbZQImU0N+8uxeEPuUYtI9pBEItE0ngx6qw109eTzQR
26o2iGriPiBKAb9bD5FJeX0QtRlHm20Tmfa7pJzRvCRLT7mx24b2zbgqOsegbKbZ
ziFY7FZuirVOJfHpBTAl7CwSDGaok3teG1NXoyqS7C7zWF68VCKZpptt0mi+dZbO
4lc7OJPQp67VDFmbiJ8jRN87RFWEXFE+2bwrmsa2qeSfoaU9GvGUe8wEHOUFKSiX
Mi5Ff1D8TYZhyu8xvxnycexc3r7/GnGkiVfthzZDlOY+YgQD9Q+ALEK8UzN12SeW
Qnz0fAqHiN2HS+lWqImELsp3sf+az4RGhsHfVJ6PEAebHJ9J4F1Pz0ZXFFY2MNTO
aiHZs3AF5evcMrkTTG/cPmOTx9xInrRQ+jZ2bLk3LFeiUknpDc4V6+HucTjk5Uk+
ZoSxYCTe1WxzMs/s8Uw0EN/I0+Kq+K8Bubq8kc2Qm2yByzqHGvZpEkKI0rnitMqz
OPja1chorgFkXzN2TyE+53nA/jt+Ddh1CIJszr2pwHm/0HJxYJ1+cqqz23DnM8XN
84XV/PSvG+aMDaJa3/FdgNmuU4mtxKN5lSOx1KonGjrwYQYdzz20qHGmv8zh3AOP
IDlBsA6P6fSBgqqARIingeWtQ72p5SpWHpnKGYCMzcIvC/y1BnvHYAiOZFVPHCN5
Iytb8H6CBOH9w5xXrRM7Q633Pljy/L5vPdN8B6ETzEgXuT2hlXjzGSQgz7X92que
vwcFikkL2n5ROWrtmRtk8Q32dLK91fADmhNZubYBZFtAVecKeIgtWbTovJBhzC76
DfXRIMvdlI1pEH9LcwBccrrXDXAlL0b80tX2Mp1sK1WdTDFW2W5Won1uZgdxShKv
OrfkfwNr9eV07e6xRmKttrJyUi3SVPfZ3McSMqI4H/yxyJfHeBJze/T8NtGJbF8r
BjB/8SAbbmOI4pEB3hOLbKd14ubgoXKn1ghM3QObQUHWrv9XF4cYCximtYwH0So2
J6imqsdCEEFPAZHc36SZiXPdHOaX66bkUO/ZSwlyigSGVoh6DyZCOOJqBcwbTheh
wd0Uq53sLTDXfgfPfbP4YKnxeVD3olvu0INAFegTDJbdYXaZ8vukTeb839YtyACK
k6CU4KKCh90ZHSWngBQQ/6r6AZXY3Ld+voH/tkBrCjwSY09td4CyIqPqk9urxDQx
ydwzyDn5gP9/TTChpD3z+wmKoM92ppXFzeWQd7RcK29YsQMu+oN0ACJJ7xQRI/s0
e+1v/vfmbB3UbxT9KUOnl0v/C9I24P3kesUBoJ6c0sEa96c0Y1zPd36Eb67GyYsg
AbthnWzdBPsrZHbs7mZS1tPdrg3mMJTYnHJBHFE+CfIDbRU2Z+dsrku/PYMeJSs8
XnA+JkdCQ+9WAuGZB6FgLqKb49wixP4jOw1XFfhQOs8X+rd1lrbKhJYoGSyxdqNC
vps6c+HbaGadRgzmPqBirp/BVjHIyNfO7q7vB+SPaxC+H5cZiEheLD4MVSVGSbD8
P+6s/TYcbNFEEJuWk46ytoUkR4NHMc19V5ID8SbOZyaerlD29ZE7BPe46nuGMqfy
O/gLddWdOY1nPpXPxW+5KYKXk5YmhNvYcfv7AwP2QATlI/iwyAGU53CjgT1Vvq79
sP8menqDrDsd7NBvD3C1beqF8YW3PI5mC1uv9dec0jxdA8RKaXZWDhkSP4Yh0szY
F5zM04TVDiPSkItGluFwbiZ6l7o0YUq2l33/CwNs6UbsJOY28qMgzZuQCf1yvGR1
GTHezY0/tqH7IztC+29PYbqCZ4buqci2XgHFgZoeKHSJKMy4nPxnuKf68DSo1yQb
PbWwE2F5uuRylZKrrVXSYnGbsBoiLsY8AlyBlJMmR/KlSQUlr90IfgjT1LWJaQa/
quo3hP6hk3+uE4zB8yMyV8HAxkkdWn181+ND1oFnA+BMNURMsl/4rlkp08Blo9VO
HOKGe+Pk8KsD+0fSFcepnZirVH7kD/+GGfUYl+HKy/9OQIz4w90mZ09MLeSMcyMp
lk3XEN2+Tar+inNjOPo1bbTfLg04qXjDWgEMkquo/GVqhA2XIvwRVmUJ3rvIYcSk
kuWogivqdftKjCAxSX3DIvQobxlSL1J83JGxTPYzQ3sMjjM9A9a6+OUuKvd8sLHk
PH7uQ0YQBD5YI2S2hPBk1MhM2GY6AGZW3+PfzR9eKBxkfCNJFXFHnfYPdVix7Vx5
C1LczAksWAtA1bSXDxxx1luaXCnPsRU3uWn41pAAAZnpDI837eQtm/ypVK+6Z8oK
CxR2bwo7mlHuFmd9wzDJx9JpSS6o1IPh8qsldNtCZMwzgwfJMAlZnL2PA7O27xdn
Ds7BUqFGbbDrvyqrm07ULbDrlpGIem0wyBIGHxZ4r4JBA1LO6Hjwpxmr/Ng5NLLC
rWL0NYtpq+anfP56aTqqD+A3xJdy44f7lkIGuFgIZwVTTnkldKcZ0p4/bsxzXCA7
wQIDU8fXChvtbzyn2qTKRUpCp280rLzf07nD7h+LXQJZNr7p5hQXrM3l1U8Bws/u
Aaa9zj0xkH3jzOQ42ISwWkeKk2XwO8Eq6LnBzeupxpOenz6hmD6PT4267b0IuRRd
y5vAJ1Eq7gzInqELNCKeQrElECkuL+1bNa6X/NPidjrjT9szygAaPcdJVUR4qyVW
Qt2z4hQe+BFyiBVf043LhFw6B6Q6elDGd4ezPPXFnG6yGzObBqmVCBVOCZ3Z+MYw
/XntmBpG4+avcv2qSXL9k43BdX/YVE3ay65UrMLQhdfbpoN17rIRlBzFDkv2kvw1
Pe1GF0yUu+mE+/d0MbZxomjebxkTzSA6yaEZhv3hPUZ2DCM4E+OOKhY290+C4/qT
pGT2N4nx1q80HERqvQ6BTqrD5u/P67qQa44f4ETGtskuVI4NdhObM0GcJmMVn9aj
CXUlAijVmjV5Kii/13YnmAcTDUqBiKXZS1Ff9/DWz5wVR8kbzuxYcG1e/DsGnSAQ
FzVLfGus9E/aTsxnCcNEvaCGhabA8B7DeXxFrjdWAXfTvHCHub4kiUs6ZaXhNtkP
G/TUjJ2BwtHROUbHO3aTsfHfiqVxcm0CCX+zPayO+IWcSlcqlZzZipzz+jrH7kpk
vUMhR9NOeciy8mJZO0HFR1wNWASzoe+mdOoCB43o32sHM8j8wRQ2QIWleVhzZ1tj
crkz3CuWQoUX//Ex12Xo6vbwiPw9pzRzsIBVtaqiK0PO5YWynVe2LOc7y8BvcKKM
ycHwJb1cOgtnOk27YeQqXz9HejtHmDE7bDXvPaQKNeAwjFB+mO918cA89QUVLkCL
NuBQnWY+nDCPAiRy0pM/U86HMeU67Vf6PyqZ8MF03WgbfVi3h3PHIejzJtwW2mCo
DW7YzJ0LqiBBHArUtn8aHMTvOHmqPkLXYEB42mXKPqixF90sObLjJRsNKBg8Ll7h
9LDqL8CYa8Fxy7P7b8TgdCWvHsr5yHwO6oy8jtQHYdt5K8hZ0Xvos1p1mTLDpa9c
np+VhYlKXbAxcyZiOJ7w+iSBAwLT9UwQZ7LMF9Qquy2hquXGKtBohQ7q3NCF17SF
M8trkvnFMmZ19QknHatAAsSCXAw4fdObl4BVxHybgdQxatweKIdcl6iQ7qRAJVCO
NE2tBOez+ppriyHQwPuNLKTrm4chzkxi9+wdt8vbabySFHzcYQXeGlMXCQBWBtd7
PmhEP1bJEmI70KU+8kDgDhdw5gXKDxgzZlT5nQEuYCCsCwZ2bbssX2AfdJ9POv0T
fw0HbzuduXDxesb2Jrxgb72RGbL3688YmuuFYU5u1omqrrv9e/X2jbHgYhGVx1+3
aOJmtkZSSwNzvJgFv4y9a6XxAzvSC2KFAMVrfq8DVDJJ7bp5eCsBJw/kYFj/C5FO
IWqWawddUkvjkhavIjxLI0g7JNngbQn9MugU3MExfhxkNWSC9LzdJICjb5I+yAAs
jaDmFY9IXFzCUeJyF46EcNE4eEnIXTh+QvfRXT5yDi3WqlXhH30AaB+XjA676D96
+97ST3++VCv1M0cKvYMqje9/JEv9LyyCppcHw8DKW/iu2BYaF2k6adZ8joeUc9wb
W8v7vLW73nbgJ+LNnsA25+RRDNZueD0aR4tGB1GBbSixlAC9SzvYG49iAdGHu3Xy
s5FnMbth86x0ZwQfor/VmQt3IzRQlfl1uks8Fu1cU5MIQLkz4ltsbZlR65rAjAIW
SCW7ji6B38qhiiLBVpytjeLICWx7MVSKGvFgY5VdaPdOLQMKSYGboYA/eEmhjWx5
NYleiMQ4vUoJkMvNBKSkhFpz2YmNfm+9Cyv54ewAPZD/o04H+vsRWlFBQ6UgLHQN
EsxjD/S/T3APj+khP95xdRYOzvGjvaLJfVFfWCHaZZCJwsCDBYUxm74eejeoeFWs
ZAujTFPM9ujMB5nb82xEUurwCk/9qPESBrWcDG2vuFPrRvzuj+zC68I/37NxllkY
JtKnAcBW3dfFRKmi0QnY9wiktKABg5fJWSJEcWFn8U5JOJ6oH4cIRu4zfXFxkdkh
L1JzHoIE34huOeojADUAwHhNAKJ94c0zcYVWDm5ynTvgf3HnqcMsI/CXyoic0ZDo
aNDoOfhZzbZRk5uJ70X7BH23Y20jOnlAPYMct3tbvdk4z2gy6uXSAumHQJGt+pUc
nw94qumQeUKT+c2uENP6ZpRQEGiQIFPgYy9/kPqjxsSCxHlx99/g+0vPBcfML1W6
8dEfxQw+OIN2ZQGbGE0cmsyqr43R9bmPKHWiobCXzorBbbF9lAj2vLM0R93w4vNK
GSL/yzHfTsuTnsL7b8XcyKdvNNfJb2WZg7Hs/4W+k3igs2AOPq8vcu4qneqb8DCH
Yyui39FSfsC/dPZgSuL+kiexdcR1P+7kjN+1gAyLTboH5kLLtG4DoZkHSj0yz1LD
N8i0MiO1v6sfiCFpIB6rAMU+RtbvZ0Jd2FL/X7KCIuPK6pTvJcVFrP1ArqGrESlO
gvr28QKmIdhkN/uy0xHLZEKzCU/FNySR7KozCL5sYT/1otIBiiLFbsA+mbMlTOXu
MW0fmIAZP2sU/T2fdOZZZu6KUOvH0pG2Q4RiazD4geSN0OdrZT9VBKLrdDaUgYh4
J8apWQl01qCaGqcIlaJCr/IWt4NcUoB8JOs5JPgz2Kn1J9pHbiczoy1cuEV4yGs4
Hic7MXP+7Jcftc9aKP4CSmvUVvTLeQ8Jv54hwGYb7G0Kb8RgTmi0nty6Yec1ctWx
Okq+CmRORY/+nBSpM1FQoUlGvvOOkdPPqupWSzBJKViz57Qlil/84UCArfffZbrb
hN7auIysEagYdhytpJChFzRmOmiUrfpHru9irJNwzJx2zaw/lFsLQcdqyyu17GAr
NEcBMNlHbB5heMJhdY077lbrKfqMXQ8Z5SV3Q1xP6jMjnuUBmgfqwSoF2KBy706F
0sBZCHD2Uf+JCyVORAndJFn8Kbzxr39Mz8FA/8oTBFAjez6IOc0S9uAvcbjQhugd
e0j21nD99Th08so74e71Ny+0fh5Qj28Ummh+eibBPnmWhSLJyBKIkmVxNZyDOw5M
f2cFDORYq7IZaDrW1CbN2taQVCI6MrMRgoAihUGrVtiHPtmHyB0J/uN/gpDRi2lN
D0Pg5e4eS+Rm8y0GKXYFdlylGQgABK1rQyKre8fiHBf6dDzDbhaorj5lAY9DKrXN
eQ69a5dTuWkTGZvMpo+6nNRQdN9qsgvZTsZQ4yi+VeJf9QWEXbGjZr6kdG0N0ymL
DmcNgvNCrtd4v/2BcI4h3FbUmirz+tT/1AZ8w7ltVJ6GuBg4c0AyCajPzFj2EIh6
109W8i+gnW6YqWr5nhyKQ9cMv4kqwwpq79QkNmAcI6Jps9Sji7ue2py3CKuJzFaJ
aWyDys+0daUUYJZTW/7XALYtBqB83tSKY1lt1vD7nQwg5uE1J1TCEk3iAkfmVULt
cL/zr723/G1mU5GTB2HIWc8ITBaM2yZYrR907+49Os8k9mRBrTAu/T8Dq0cTORd5
v3v7JyYv9D2J6vZP+OKP8CwNQ1sAmzC56r/HTcGC66Ppt+IfNFqhH/3Qi47B+rAT
yYmZOIxYs/UhzNRgiDaWZiZt6g0eWprsqchX6vK8S9SY07VuVq6Wv4LOO62R9tSt
KhyzuSQRm8Nl9s9bW2OBqCobqpdLyc+9BQmYvtG4MF7zF3wIaimKbB5sevaiKZSv
BV1Crk45QbD8G+Aig8+Vsm6ENILHNbykaoOSbqnCYposT2wKpzSr2d6oHVFwBqOV
NAKlLPQZVY9Th0ToOOSk6ryHScvo8i2DDt9yoixK9kXgK9+OOWKoxhgeD7BTiKhd
Rvys8b6WR8eAXgb4adfLVbhdx+qnsgwwHJ7Bb/WWmak12xbiMgXoJPVZTi/a1Xn+
XWOGTsJaZJSkY1JZvamFH8R6R8hp4kdtKmS5ujlYy4RY14+W5jxUP0uSbo840YZr
r1L9HPrcSD/hRNZgPCBeL/39EJAXqBKgpdqdVfC7RbHccCOqQB4IpCvL1RHhioln
5+MnnTUJ98bsx5tc/P5cOyfSKLhMOvVOCps3+Ij2146jIETxyNhT3rLMasY2Z8jp
tPQBbywOY9QgXenPcsk2M62m3d4cIczT+mdkRBXpP4g1ceB9DuzsK5lsnDQBBgfh
jQyw/JVdugk4SOpWllum8r/W8pSjHMtSTbhaKXssEYQB0M0zU5pNIPdId0iv+a4f
UY+E/UEyVuBV5o+gIiNgkQMRFVmjSDXDG/MHgb8/bsDI69ZSJFokDDPr2q4acuAg
KLqLzVYl2uHjztRQsw9BYrJUvtXTr4cuIsoMoOd0E4vC9dBUrExGhUtmkpTpr2/e
lzSM/YUU39MNzgqhcCO3JbVw8v5ZAuJxX1cuQjc87V4Yuw145MdQbdM8BDExmX7j
lt0VK4eOKVz7sqnghoFw49ybM5a+e6Iq9g2MvGDPC6UNssNbPNRKNGZCxJMug0dO
WjYsa6MlaemniNfIfB7I3JFbd2XVMeQXbygqW4mkwuNn1O52jl4YEBXArTlhjv8I
/sHl3Gc95dkK29u2JF9I5ScBilgNYbpW4yz3MSLiGzsuDsO1zcdSD9KPgABsr+c1
6pa0Q+S3bU65mMhRuPcr97mBxfztaHxjoG/Xn7IRiqHxPhu8IFwGGGoA6cZ3nH0W
wSpi/loBky2PFbBrPV6Et2s8vWg2YIa518dbKs7KmRw4qiyMkBIHI2hZp7jZoyxl
2szqiFqHVWlgRd5+hCiuBW+hxOnNYGQBTyjNXLT4KArJr1c7o124a1L+JGRmia3i
hVdicHO99Tb58BKjnOtKUhlcJRw/XVwd1NXGaQMNxoQYYBPrt+o6FQSO4o/jmq6c
gNy3kz/Qf2Np6/l9xs979DcGRWe0RWMAlYilpsHTsevuHzWq2heIfkKkvHZK84Em
pkW7/q84P22kRvnPAETkYEauwEiAFlr0HDdggrSDTJyn020OZq8jusPRsvh2lp5p
vsLAFxgkGs5c70Wh8MYOnpVjjLMjPGg6WTHJsmyhiqDdu+yjIBUEw39Pc2BOwoiD
1CU2bJlra8PJhX/Zb+2qy/HGnfyC63ySptJL0gaMii/RaCOmSQe8B3vJSXwPytNU
vVHfC8gcg+W4OLsYJiZr3p0gwuKNwkr0hcYvn+bMePE0GfNqC1Jh+9/L3rga0BAg
fGkKEeyxCz88wSxUT9q0hnm1DLQ/nVC7zcvr4nuFJqIwy+5JVAo20I5td77pG7JO
6JZYBELakt9q9kM5rCqA2ShGbECbPOhJk8wkQG60OwZA/z7snu3Fwv6I4xTEb24Z
fsNuf6i1eCZdoukaavmmWOgiPyBDWWoyLPJuj2IGCrVNlXR8JFueQhC3Xn80xAoT
kX1O7E/O9Ia5wndhBMQyUTkntytz3iLTAlkxZAzT7dEFD24j2ZqHygXntw8BZGea
i+QWr/GmUTLcnO/J3/kTKsunAnmkxAJIjgoPttu7j6qNhzZ9hZShq2ovFcbs2tW6
qyPx7J2NlXunFkaCFSuJ14UsgZ0FfU3Xf97I968o/+miGwE9WxvkQYNKDQl3uGfx
f0Wqzw7V5ztNUib0KW9+PPtfWc08HLSxMSY2KB/gfw3mtCVqSe/N0ie0tONi9nRN
Ax6Rd+biL869OgrmutES3WwMFn6+DuK2cgCnDIhohnoSwW16q04eLPtAwW6vcD/w
O3wF/M10CdoqGTizuMMbi43RgYeum/5eneixFZupnjiM6qsiVylwAbLAkcgWvwV1
iIlI5sF60q9gPlpqMeGawVjTpWDmF24vwyxknfgdVxQibk9n3xdIBRbuU2CoZmaK
k/ObC7r6VM+/IKMGAZJLtKcIODidi0fHIouZI+DbfGiv5if6EyphlpgOgpjEPfw8
JCK4REZ2HAjkXkfpxTceMoG62GpuaIT6rh38c02C3fi6ob856FSvBWnQwIDzS1II
SzpD6SHb06SWSBrLDD+tO+h5YccvIq89bQ082Xh74MC7hXAeQBj6sq/niTc04W6A
yl1oaf+Yl/jJRR4w4R8cyjiCxJpeWfI9Tmhu4M0Qn8Sfh//+Uz7AZvXtRIlnmZBl
9NkeG8xgKR5B/Mf30SoBmS91TgIe07NvUTORBXY6PkNbmxUOTzgDWMO6zOCY39a8
KmLEFd+92amV//pqXwyibV6K9lWg7YOcu+BWUp5AF70lm05dp6cBqi+3Wm5dngLx
9kz9NKh8Tc6A+rMsWbN/c23FFFpl9awTTiJENmI+S+pRHg+MRctuQoBvhee8uKWF
qtOI7UF8lloNkbWg2EMbghyBWRpIh3rf00/WCKznxRCfsTWxFqY76trSxtqFN2wk
B75SooFtS7UPIaRpF1b9Bk+bX4CjYrPBdreG+KZT4z3wNBg0Ps6R5/goeHthRewN
EhZGY/QTASEQCI44vTZDHBe/KazV9fLrCAHRvSlEml7vdb7xCTZWF+qKPErzW5iX
siF1qf6+CVKMQNIoBQWmdglFQ2/A/cvyEcXsUQVHU0P//N5zsgZ36BhLJX8Zl9Yg
PA594eyr8zA2zbDF68XDH0KqIWC0w5PGz5o8K8096e7ZQPEGGu94OoLwCpLBzXUO
8k3zpDwHnRhT4qU1gcOosszh+hmt4Px14ExrD3uPm4XjuJR00RCdmlgB2/OzE1gu
rZHXK7qPhUCuLBH1dEUFIUKg8hvEaBpAFWjA7SdN/3+b1fbvbRMhNk6kB9SASQXH
p6y0bTeDKtbQZNxIwKeOYSF/0CEbpEmWOBRvG57fBnFKyioek+zKs4MMo9qgEc4h
zeWvxiem6eRcNfsRFZs6o9Fa6t+KXeR0r7lXghuyWw7YxYV00aRhKBywNLHZpgND
z/Zf4ZpfCpon8qQ97vNs13xBoIoD3CtuVoJNHBa6kwmCqrNCTo9BTvsNPOl9NmRT
JRzzeTnsgpnhqttpGKYNMng299KMuPQzScrEIqAGydpQyCWkpbSwAgsuxYUaDONj
xXLjfsdzXp1URQcbrKOPCaq47dGvUi6WANuYwt2PW8CyXJmJ6zOuUC2Q2XzMQCn2
9+zPvS9PvYowe/Gxou5RulF+iOLlqfZIntyB0G/KFg55hDXEduKUcmVf+jP1KUKH
ddXFdZNkHfSoii04xqhkw9XZpfgjAJTvCaqebNz4iPwUjI2kjsQbR39nQa+F8Z5d
FQ6sBOdcAU7j8dm86dAMwwLxeSWVqwxWcrV9KWf1GtNIltCJt8QEoytNtt+ngisJ
S/iKfgL2FdhEqPEJmmIj/lv4WsQM1mWVAGwP8nW4olCB2b/4PbM4BGI1h6WHWTkY
P3FoZ+qVtRuZMBt0saj2SQvotSlVNjPbB62zwZrBldAna7ILODHWZXpDY9p7nQ+7
VFGp8HzSv4DebVvqSqV9QvsB+DZX+02mQZ3aiAkV5m2NgOpBOKxmaglp0uqMep1f
RbPvAfpcNKxShu2D8t0pPIsmR0u5ldgTEiz0aj6iI14+63xa3iF31G5iAXAZ+jg0
leTNmFIliBCSUhzN55KYP4b29hzvprAshMz2ueZPT128TZMw2tPQ+IulMToDG2mv
5wBllKKpieIzYa36q6/HRJ5YS6ml3DFch7wb4V+9NweMsNsuM8Q2s1w/gfTy7QKG
FndGvAB57sDSaoZNktGPF/1VcpxYaiXK130MenStYUZi9XPxhFlfuENHJzpHCYAe
NALURH+d/NKgp9bO39s2ye4mUH+TlfRkMefPXl7BR/xIs99/C6auUysHrGzT7jND
DXML1YyKZqJsZhWJreb2lUU/zB69Xk2HWedMy6VmMTCXTo5L6cZeHn55K/ifh1uW
NUF32dqnBHfa2st8cWIxhMjcGzw9W4uitiwObc4N2VV527O1IU8predav+YFecGB
jWDr7CJ/8IffB5qiqF6jaMPboniBT7a+2qWjNPS/VG2m5S6hgX26FncKC4FmJDkE
h6/1HGxc0K66ZTFztE4yS5x0Ks4iN7oRDO1mohCQXvv8pnGg3j8u1Tfbct9esDSX
YCaLuBGPxG4aNYCMfJPF1o1pyxocwrclJtXuyngAtroE88QRQR1HLbdPAevL9B6Y
x2F7aUYjxsZO+GNcwDmdPuY1kyrcW3R1Vn1DEZaZDWNFy8g1O/eB1kNmeYGehz2e
1KhHipHZCMhJCIrQxa+QGCHBRVytIBWg3nA37GxemqX4P1CYIve6vbs0+Ah+E5eV
yMNQPqoDaqi44lbc/YXb6VhSq3v/U1iccR6pWPGE6SdQh/sNiavwN6kkDyWAsUX8
xXVODwiR5aFlZIpA1eVxcpyOBf6tQf9OFWYJyUKDRf1jbHrJS5oiQ4aRQ3HX4JmI
ZJL1nNIZp7kifHW88wxmKFNK+aImA+vjfXKbl8+yPDtu8WQGij67PXOVevju65VE
96U7QKPZssuuCUcgJ/rKizxQ1I89Zxwkm74iLaWhOrEEV0U5VvyQqQ+bdcHUw8Ru
W6/dsmK6Viad3wY9Ba9Lnzjm5DhBMB16RCvp9TZZUZTAO6e0hAIgqRRTRsGwnmlD
ln7GfKVQktaoH7Ul7sgvlfY138gV5zJZhE3uocBCBO1JVLBQ2cAoJwSvwE0+1Qy1
LQc3Cm641j+eP0Ofvf0fqyGStq77X2e8AbkZVquAvqS56Ki6YWbFR2Xs7Rc1F4y1
qPk/4o7bgVZLb67bu85C8LaOZEokF/me0g4BwGq56eTfuEJaJycz0CvTix2eUko6
PE7i44Y2kGWL3cp5ak5OOoqbEFwdPl9a2d8OnpK572fMtod9RUrlaaGuiLWnGUOu
sQzrpNjHWvEA16OqVTMPiVMx69bOQIru2bcD19kx5urcD6ZAWsnmEnPphodqHy5t
nVaBwW30wATgZBli88Mq2AfLewhWKXZNj5Buv7iIHFhYnottzMKI56710w9xq0QW
fNFSMCenFMAr6rGaf+PAin7enmUvmVz5nY7xkAcVJBFzV3YwsloeoWVz1OBVYC1L
EBM0iqyKGizugZxPbv2Sd2DhC+wjY7kYw1LZ6+8kb7PYPsKamQjcXh5OUV3MZEZh
LzmzbmFJWA30u6OiWT4InzzavS2X6r9EtGyO2GwUcNfAhKLYbQEnKjiBjSl+p1x5
M5+gLV8CSawoLKT4pah/4oCLpTb+ugap4u6wxz/993d/l0xJklePSbPOtWiml+Qx
wutT4PfynA7xCK4b9L57q33hIhUJerr/jA9ZXfeBILQSKSt1kU60/5NoF7F8Ow3n
plVQiB4jSTCI4Qz1zSJQ8D/n0VyeAksL3bFmBXeOhmHmpdv0CLF6xrTZcQvVi6Yk
gWoYYSj6weooyUpRgOXDJf5pbnCPb/GMoQMWJqsjfVqSOJxUsxiK+pcNUHmWNa2a
gSnK8hH9gVh6bL2f7sPMoUyjeY2SgBlfPDts+j796uKf6yp6VRd3SFgrlLnucHK0
qbFrBnK7CkXMmBTZ0x2MELVy50VXpyQf79MR+0EUFJiZ7aUAsnhlO8fPl+qM1uXT
hdrmD0eCFywHRAr+sdPdAIlKTG9pq83x4zihIYx5NWjHnyf7szKE5iEzRRJBzQG5
hcSlnqSFR1UwLssaSPOJPJB0bGYaaF2O5deYIVEkEGZ2HI8U66m/NzNbzD2ga8q0
P2I0QhnWOXQsaj25VN3axHBlzyhpAECn6oYdZGSlo234yQD3m3Sfx0Tn0pkJm2dJ
GJhMiGfxt6foJx5iEy/VlrtHzd4GugYWta4OQw9arYfFDPnyJL23HwLwbVIFrGxU
iXVdSq4pfyOc3RpjTvTKDv4yjBl/YgYoSTHZMqkAu/pAoHGfihx+s9yBVZNynrpb
WR1K9BnEMAPA2bdR7EfbwMcBSHvrjGEcfimzKAe9eKqCT+rpyax7Gzr7TKIIDYEy
OEcS68hbc6S+2sC88lqLw8fMeX5LZhX6SYtpC9OgUp4C+Na69EmDHMAhBGGWgn1a
TjjPyWTbtcIvnFfKrGQ7kc4GEzkU1KehjWlFYXTe5uwmmja86yJb9ER9d9L/tz+G
pAU80Dvoh4uR9kgvl2N+tEcIu7x4++vZ95F6mH4XMuew8FP42P5F0goa5i5doYXl
3h+fXzqm9c1m184nIkjySHLg9QxWQKDg284SC5zAy459+F6UOfCiynfUjBv10XEL
H3+3W33LFjtK/iynThX+0f/LeakN4Svcw8PCR3nKh/hIFHedujaLcGGbmOxQIWWd
SIKeyUrJ2GC+l/HeMYlxj3D8VOXwo5GCXrv9TFE+Vb9xhtxhOegg67Dcejp6/Khk
Ekm0oW9ITbFQn6v5gOqgi+VBgoslrtFUy8Y10RILQ7NXkF5DEiKySD9UbPn7gsMS
pNO3JZb6dHSSmV0xKFd9TjQj+IiF/YPSVFSTLSmh0OvMtZD02KR246rGt2W/KJMl
SN2XUxkUrEXUSWmQkv1xHQeUwt/H+V75hHU1q/N72UQE41xAhc1YGROdY+MD0RVc
CfWRJT0YmS+j4+wSMdkOcqQdO/sOFO4xgXTaS7HDRdR8w9HS9D6Hj/bbVBie1z0M
EpllesLrW7VbOXLruHBfxHGz9zWxQFjEcga4a6k6lNOEcbwYAcR7mo+/Q/yQ4TTa
rwFYtOuhkz59QQ/7SHPw8qPCyzc+SDSbMU+Tsm1FlQgYBIgJ+91mU79fpyHqHUcP
YXB1WhTdkMjkTVuNLrSbuAeU47qy5n7RFGM5ol7VyADboZ+OYrpaldIa1oEv1rBC
AybRxWyPgBRrxayC8RPBGBOeJU9UzmN4iO3M8hDE6i7nGypSSkZaBxTsfWzYlLuo
/BN2BHkJDCHBPqC3QSo4gxAB+LmjNBcUpSzxeHYSncXjZFBfGkfrfj+iMvggHEid
xsyvPx+nETJ5VPBWvKxQTjrlAcA+jXEzQ8tvVTSuPOAV14QNgCuT47G16ytA/11F
B1/uU7Sj2qCGjcONuMFMNNVjPX/VnAE9Sdi0QNVtvRKRuu46xrBaaWU6NpWZf9fr
iB0vazzbP3TNf2xBY+lBXP7Vugg316NYz6eEmQgSC8TiZXRNB2S6hlYs+cv0bVxH
vk56HEwkqL9+yhKOzjQZukjtEoiczKoiOcv7RQSNvuDJE0p4mqorx1M2u33kFnUf
j1bO8M+EjOLDN5CkWzwlS+D7fs0KsJpRPgb95f1AEdx/0+fDqr8Z6bxOdRPnabX/
vRt/cxNWfk6AASOAyTMYGOxpnNi0bNSVBWQb+W6z28F58NnQwx9iHLabnyA1xH2k
zAdhLQWHTGCcKfDKfgYtlF5GLwbwfHj+qKJfB5eXTDal52Yzf9/N3o3y+U2hgUWv
Jr55doGbkt/lTEmJyg4EheLHj0zgD2Uw/sqZKWwEWvaMMkYNIr0LSoJFuJ+KIfRG
vffme7foJOsdNn7/E3cYeNIWnbKkikSU7fDviM8IBTuhKNh5bDMpZyRynUXpPOrD
+XDHR9hXC2fFp8AzWT+3KfFJmhLZMeYE49HLIGKXF044WDKkDodHhbiSsHqlFLqR
fuJl1JFSqjXivy9Vln2qvclHrqtSF4ovN0h1On7IAjXuaFOdwo8BRII2J+1q4/8Y
hJbTXDrTbncCJpg7fpD4mvxq8umJDw8vC2ZtHNOys5psJX3wQ+9tPgM9QjjdT7nG
Ju3mWQPTstKnfHglsQDIWJkWbPu/ZRGz7jBXNiHJp4DP062I5AfRPqxSnLU1OEOJ
sinj/e41UuzzC6jjw0AG+SQIWDoH/tHyBHxoGRMWCIdWUYNFn/MBqh53jCzXkuFc
9KR3tIV7Lu622c2tHERrK6tH4Vz992hSKiKn0PgYX4cK9oaVvGVAvs8xE1dExdxQ
Jr7Dkceg0FwlxY5JNbgYSb/408cDZctngn4FNtPRPtIwA9JjdZK1YDIhkVU0i+4b
6w8XAMv5M1sNcfd38QgMPlJd3YW9disr+ZX7rxIpl8G2CjPtmJgQibE+ReA2FcZA
WNQr+na6hYC+SiQGDQHAQZV7EYPwAaFKQ0J02pflu3WPhipUL1QZquEvVDowhJrA
6B3QujIYbijStZrM2xBTx2DDJpNPxtdPQ0MZ+01FUzrg60H9GTPjGhg8AMD+HSYo
ZsThYEEO6yPG82DSDeuAVkAiGZ3juwymjYt23DQdqV/e/i0E8Xc1WwjcUTlicSqY
meX1raSCKpjutzbdemu8sQD+Ssx5Bv+sYtfG01mXXqZxL6Cj0EYzn6WMDFac2SrV
uDW+nVPeVuB2cq6h4lVMcMS82TGasTphmdoqFAIUf1Ln9w6Upn7mXyslxmJVmpLE
r1k2P0xBpQwPpuHCVeCdupPGeNaxyws3/DTfpmGOlYvsmC7TODk8g3BFKuxrr4vX
u/2WK7ijXXchsWK6S+xDtrg8Mk7Myoufw+RPU0IqxmEohpFFXcWKsPEEU6Dt9SEJ
u8lODlLJdnQ9kkrgls5kUSXJ4aMOtJrh7FI6NK2qWDvdI2HUw4EQ+75mnyOTCz2e
UUusVhSh/9coAl3sh+zozlAVuE58zGW3/71zTCGQOP9AZ18UqGiJ947JSQb7oqi7
huCcnwMPrbtESTYOqZ+awTVfm2LGDobQLuV6y4UgQATQ90YnIYek2oNfIPSGDT1N
Fvgt5KVvkuRcXaGR+xwvHqWLuzdsKwk6V4bE7J8xSkuYZOd3DTVslDqzRcnGeKja
kIXDu82KqxFCueUr+lsnnpRWfJklPZY9jMDF4YrBF96wsDroKuwkxG5WTO4el5EB
48GBOlomLhodCsGgtZusAThJwbRJzT8cHCvyt1J1CbHfnPgj6NdYfdlMcbY/9EDl
g+zIRu/g0SEefAC4yf8lihGpUzL7dMqLJ1ypNlwCP4cuiSuPskuZE9iLhWEAWji4
TXNu3oBjJMKCQo9a9OioOq/wVSS8V9GLc8RE0OALkj1SEJ+Xquo1ACvPUTIAnY2w
S1/laTFxdXANR66S7B6p1VzJrzpiG4fUIMt/vwcapPXdgRxLDFSkOsPhubJJkBfa
IVHclhzlJH1M9GzNogl5v4/PCwikcbyZcY/dwdcbGlnDpaE2d2ZlQhT3lKQyfWPq
zRwakT0D6YeEkHE/yKgSl9UKsQxtMLiEUFiFzQVF3od26ZOyqE0IIVANBA+gMB5s
LMmG9sIjAI8wBwbTQQP1ZBLozK8RFna4Vy6HNr90YsL+BPUXsxcg5Ibp7Hflt3fR
I9an1+deKP+zdeY0RwbE2covqBbcOnfnr4cIJ1in9ORMVqaNWgU3gR1MFHYB82Np
IvvtijaOOfluZyXjpMFYHl4mBmo0Lez+aPCZhu7HkCR7M1Db89pX/zlZJ8ybVI35
Njce53VjBWyAcz0MfEV4PnXg5wcz2wV4m45a41GRugB3BtJsw/ZcaZjC76KGBrCO
GKlva8Ze1jlZ1G/mDYB5frsWep8CZaFAoR7HjGmI74AGsVzQMlQFl2CZd2IU+aqD
Z279oShiknBaNpwR0mY6favABUXnyIuMCVBwNXP5E/2mrULYxJhb7IRwSyRiVa72
VEjRPOCgpr7o3G+bFj/fSoyEMhs04wYDvUK2bGFnnLv7g46BsTVzKfkoCN3sS+XG
U70Gl+NiwWIbygqDbgCaMRAxMbvpeP/CyyXAuEy6F7pcnwWiJG128+xt7+9cqhcb
jn2g/5ycJajb6yfaHqYd+My7XAdsMbFCCHmgY7Jq3TTMG2kkjEdYqZ4F1uomXl5D
oqzjo+e0h9y6fgNeGJKCI1WWx0FwoTZmbmOipSyMYjvc1jPRROYDpcc4iU4y+yhp
hg7QW4KenlheGT8yX20CMt+mJqIRHfxhdc6EBwzRUqB5S8p1XU2YBGNVd0JvqzCb
BIqQE7lwcw3LKFLhMGVVbt5NNpZtM9VlPLllo5WzmH0jrnW9B6TWoPZCrVl45/Dp
lkKk15vFb2Dq24gcUSkAkkpSoCTLYu3M8Hzgy7fVcUqK0Trx6SNtAcYJSVoW7cXH
75tbdSTmVZIXO6OAkpCn60ocLsK882dmDrov/LkCCr519lOeViQI+i91yqWVFtkb
CyDFsHo6ijSW/7gX/GFbj6FI0lKNLekgtfJNGs/hHYMtpXU9Q81xBCQk/Tvr815+
Rl03jAps4hIeadeOA5GkPlGKJ1tTZjnFbBtdbg5x9iO2HWuqJAqg/dmyD1JVDPCd
CUnoz/C/inMbu5nHxGmBPTVqsPGbEbgwts3c9Rsaws8hgbrAnJ0d/fL15qqczHop
dHtXkwrYw/QAXY03QrUXzkdGg6Tg1LeXYmEX8BG8LK/pEveRT6nmZ0kZbQgVfAi2
wOSvyAElsabJ0OzrVoYxglUatOxBm66BEpLrG/Fy0LvE85SKs6DttqqRTi4pRiCB
NmpS3JLW4mfTjYRMOYmh9FW1aTsSH86szMGoy/ue/TvNzLDOKCehIQoapBpn1cy3
NJv8F463lWBKJDasHxwBXMVjN/qS/StlguFESIs3rGh7p2Bqkrg2QY+2Rn5xrXdA
IMTKCPCX2VtU3tZh7cMjNe6li/i/RJ+aFGvjr1Q0lGTk5+D/3GJfHfhCQBue7Nio
K9Xdw8Iuh5W4sO0Llx+qmbi8bdlZS+P++xxKWDt97sUx+v8mQifX1oEvaqpZ7jQn
NpgK1zll3ZyA4YzYV99X+3I7V+BvOXbeJqgpiAlQCHVa4Bdf/cKgBoE0FAgmwrIo
pzJrIKMY+VT7UDbiP3bu2Pq7e4sjjme6jOMdqEiRsyRcohugY3wUD+KRSo/uLje8
BZMN2ucJew3lMv6vanYCLnic93P3LDNQpAku1SnJcpybHcdS9HWwTfQ6iKXQan+w
87OLYN6sCSRLvKXCoMdphuqW1Mk0eembMQKCwBO3GyjFb//s90k5fGtTu5A6j3hV
fBL9lQwLlouv+uvf7gr4SxIHA17lKCO6Trm6Bk/+n4lWqAThhyTXhAXyFuqDdhr1
FAIpjhfoOWoFVxHsxaOLHY1faIOaTZlLitUhLwZEVk6NJJnukZl0QbPsQNEQO4tu
QkeGEB3K3+Osi4rveT0ze5CnvQvoeO314Yq+yMPxwfHpJfG0QJNYl53DLugZm+vX
4e0F2dx76QQD7n87cBo/fwpxOC4Y1UdSRwQXwXFCcsQ5qtEFsuALg8e+GsUGmY00
zdbPi1LW7uJKmC3ydhSBXE2gdwlXlAu9IQ0Dt2dpVDsPH/vDunhuTvHdz+W1L3E2
3GHwX+h4e4DXZUZLM5eHuU3J3aZpD11/apDEtV1B7EUhGB7+2tW959qncn42zvPh
AMzmbiIbOx2OcR+Xf9jM8wviHtoUYcw/GvtyJLZovgnXzoGPBXwh5v20R6AGpXsn
EqJPyk6KyT3pUT5GZ9Kv1bTxmWuTTV2aSzVfvHWZdNdvz7bB5BLaZe5EiKivB58s
AxjD0VPTPLUa+SU7Ao9pYOnTJYg7eaAogtBXicU6sDOlwMxUSW3KyxLl/0e+ExQJ
2JnWruoMbJ8J0aH+ku9YknyiezhBi8mvmZxU4ax0ST6LpkltN02cdQxUzN8qKK0p
UJA1oG8is8RafQzGjEB4WcOxFNYrcfyLUrIBad1AySZPirhoXfLvNXp7W3iWZwZI
2dBO5aePsqSMtiStLAeNQ+bDDp0Te3mYF+l3lVOAr7mkSel5zMIypkn60uchGANk
jvch53uscNq1irO4aQVA+pN5nMummUB8QkevibAVw3yeubKYehkzUXTqJu5Aj6ib
S3n4plhw2HL/Vdq+hm9sO586jMBcyzXshbX0VvguayroqODKjUYAatWjaFITjWGw
dTVedcpz0qaUfwawgAVbOftzATyJJEglsQDtuo/8lTum8LpaWukux6pIxD8zw9dM
jZ2tSJOooD2aa2Wk/9Aqdb3hRq3cf8EJwFc3ID4MVQhUi/fTuDpdnsg39khwnUcN
rE07Lgsv3QpSowrWz34dAWXAknGBFjH0S4M1/1ysM9siZYyis3wfvyyW8eH/kh+L
oR96I8XED4KURTJgJtxrnvsKKywg7Elg4uWVMgDVRGvkbtCr2j4J2isMdb3FUBQL
8VQVihoUtNE6sx3dvsgpdAp0xaVdOiFqzMaDOvAVswOY6G1T8VBXDx/+nDLDjnza
KfKTEFXnrigQIGp+4fgqUldcF793uZmwldXpE49SAkabPprpm1+qJIoiUH3dk3tc
vq4m7eI8UnGEz8z1/GNqr3GRwQ9Fl9gDuzYbKmlq7w4Hae5W1hct4b+22PExOOZ9
ve/UhgtbplURkCm/nHZUueKYMDH7l7+uLTgolzg+j//+DJTAc9+CTr5U5ab5PZsX
rvLJqVZ7jrdqXlHAg4uC+Oq3tppwmwJJqDu7VhZh0DnDeDZymTX+zrXbEqUGblsU
ZoWR/RCDE4Ew/tYj3whMLUmg07Xu5zYhpk06ihi4LerKcn0QRaxgpxdca7fsvyyB
usdDVsu8Abh+nmOP2aYCmYe2LoSjKAP+Fbt3/0JaK58VMD+gA9nEuY19QmddqJtu
jrFMekPHNUxquGXFxFkuxR6qJvw5TPT9bY7r36o61nplPzaHLjWuXWBJsmnSTJfl
p/r7MvItm77j4KjHNuSXmxEZgMmqMyxA3ArUJIsStxJcn19Ndy2TWlOX9G9dzQNZ
g3gJUtzeYFKTmeBMhajTX++j2RcqHdvKZIg76EQAbp6Y5pK+wfG+sumK/ewtFx6x
4bVTxhFz/wv5EVQ6n8ZHa0ejqd/xFMXKyr2B9H9Rq6B/x3nf7UPmcOMshXQzIAb4
Pyb0J2RZLkVubvbcwu1p8qYRFPM7KyLJI50jJJKux6w9yhFCELu8xwZU6sdodt/Y
Ovz349DDY7N1HJZy1Lr966ZW48nGvPjgFqqoJ9BehOQTf4wohhedx4lzgj0qSEIX
XMqom4DEzRSiCUQorEuQuENxZsTtIjjVIrcrS8VJyvcyI19htkYrDv+nhVeGnmzT
Q04VUBug2LapUqTzwzDcsIDK6qQP6L1VzQAZEVjh7HKNsxuKcvewWMUgYxe8s9PW
rUPosrWFRdNecLcvfUO5E7iF9dU9OBNtwkUGoUua5CKqOJfRh4WC7vTu0Yb/pKxv
820lfmJDKEOB2EEXahk0YD7Or2HKkgoc7pofcSfC1TWt+qM43QjynoX/TWJamtgZ
v6uafBxQvS4LQ4tiw2Q0hK6jWKqlat+eaWaKARJP/3oeVfZTnDSMGNVLrAxyt8Uu
Z7lv+ZYSypUfShuw+9VSfZtb2AK+dc8r25EX9Ets0Q8bkWTDcC4V9MAWhNyQbfyY
0BzpAkOs5INAOji/bVSsyLzhtFXbSbe+jbtOFwQaAIRtiKS3+KG1mhOcbshJf1B+
BcmR+q/VnUYRixsCDcdjJ8eySAdKbVyhoBhpEGdNXZOiej2qJoGcpSaQ/xqiOUhj
nXL4ZF75XRiMIE/AyzmJYVwMSAghhI0iTtlPuzEK3cbuCqkKu9/Y2QQICrH4OofV
pz2SLDiTpyW9G8+vG6UMHuAzgIC5rVed1H5Vd1jVq3a7luGOkcyPv196ayF+F1sj
mm2G7TNhgHPFd/Kfgc3Naglrr7SZ95f5mIRKOhl5Gs/2rPNwgzF622ecNFVpdxRB
SNdFZXIbonbaYJXxC6SGbvKu2vIHbWQbprKFE/S3RxC6WlPgqLoZr3GOeRiS3O/I
eufwaUaidj/MwI/BhZt4DeKYkOAJyEs9sT7OLOsecsym4EAhSaowBX5NQCHYT73Z
XjQmMQwdCMNUMVlYszwSP62XzZLvFuKbBk3tOCouc5k0B0qfddV2rb4P2AtsuWCd
QkwFokV3jlVdVrMevEaaoUfHkSBVX3CWayeCIBBJOCVHoUWzT/6uggtV01rYuuYf
JXg8woz6Aadq5DYCI7S6RQoFkOL1gaWcx2tCaul5Bo0szqoiQxGE9Y3T+5nN+phP
PYlbYip/TU7oRmQrjH8aNqGZCKMunrYvVeksCadHQeIai++IIFziW7BC6xUwUxag
+JHYSm2i2C7HUFgrAvGe4+dTLz3KyZfgPTl2QwvGnG6503EQilvXXpPb40axJs2p
KSD3leQtonDT8Ozj8DTzVUgYmN3psxF35MaNdo8tWkhub91WhPUUpUJtVwXH2MnV
3cR4vlyI5/ciymi0HbCbA8Qb0nd8xikfK9pei7lv0HqVsbzVHPHZmEqW4HoTQzDZ
Dry+bgnzxDLRwO4aqpdaCkWLiO7pFiIRFRoge9OOeJ6cgdwLLNNHcPgltzC6AYjw
DgMfsuOs50pYeRxKRzm/0e7CRFyKwqWnyjHVzrduDGGB91hCzBrr6JdUkDAOM8C1
HrV+tYZmKXkuklRpBjrTTfGb7nA+N0rJMQug/+7LA84YfuKX0wGrX0eCZy4IY/M9
qvxcO3M02ptLZwFaowZGRw8Kse/aBaY6nMcPkH8qZ9itey65+OrQG50haq6o4ygo
ZILmldLNwRcWIvAmtmdxlp/PDOzXsK6Op8kyBS1SZToGuXRf2X7q5e/opazjg71Z
3WTxiY/z5mhHefl/su/T7jGWobihaG0+tha438txL0HyU6Fa8dDocSHreD3DzhZ4
epNAWTeSZQYBcBz20JcxWQUuDaBEJV66P8JaXCK5zsWFeb3JUREZXvoFtXD2s7aR
cwk2uYi7PexZD3pnMxPraTph8PaoPS5NNovIWV7xB9BbUns/H8oRMxYgN+MaX2GG
w1QntuetRR+lPkgrSQaZcgmRKQbmcY16uw72WGe2X5mNP5PH9GX4p6c7dGoBP8Bj
L3qODTRCtqlJ/9aTbsIoJHvj79XYGwz3mvLQp0rM7bKuUoaa6GxDZawXwkiMwW5p
Pgov9i/tMTYr4AVskgoNYxIDdvhH4Vpf1bz0WbhLhDNjkcZaAnsflG90JkUNbtsh
qHcepr4MQKt8crONCZEIxClWXec8xW+EOYgUGwUkgSESZkTKbRrTq9J9p/pwhzZC
I2SiivzbkYg01fTOx2PU5hMW3KFaZM3LcKdrr+jN7b4TPiHQgouA3bt02+nm1yQV
I8/eoZd3Q9n9iLi0c1dLEO/lu/tYHuAIFTs5QqBe6PkhVj8YXzPWUc7dPi8iv0wu
eDBo/x0jfmiMwGFHmtn8JLjQDQ2xYJBvpd2neje4aQyamCBvV31m+4603xNkE21T
ykkqZnJAyQmq2lmFkCZC+hF0jKeJLGIrLezmbSntHWplapixcT0sO5tPNJlqx2Sp
nEnnWu8ZVLppffCeV137Kaa5UhDII8SCdHkUbfyrVw4d23iDG9SW972VQnnFx1M3
3+cB8UtsS6/qig8LYxAsTR6Wk+5lfsLnU185GMkCHDxX0lq5j0rOb/VfprKAMvS5
4W6g7CiWs4rJBi8eb9arC64oJp74cDH4D0vt2DrX1A/dzjms3p+ThVR++XqUJPlq
pBEfREKEAnYSeZi75mzElT82Rjs0ku5doeX4iNr375XH73kinTuos0+cihJsIvJh
qJ5VXtbCkkVRPaWlILHS6EITod2Ji4X6RDzFwFADp7li/cBoPujtRAInbIX57Luq
EGJGXGzvy57KcetMJfPSAuGd3Td4ilEO4cUf53Q0A0lzaDIRkExguw9SuYb2nkPd
WQttt2jNVJFl2I/AyR8dCwJaOTBo2vlv+KV/IoAwxwBBzt9ZC+/0cQySD3C5RiCU
JNFwVQqFIAbnZsfmWoozRDLx0sNyH70ZV+mjYOVBq+Bc1QmFFUSMCPIJkNnysmbT
yHXLbJGahFrYgjz4joNfxd5z72KRNTEThTVUorhpzUEaotHszyYGg09/b3uSwkgQ
/aLtB9xtE1VpFt1OmLAetteW8GWKmrvnwSJTucNCOmQKr+7oRY88NCg/WUAp7X0j
hUXqJwUUaitUJg29apkahEJWjH1u6LmVeBLt64m24ss2Jg5LD4x0VLnIQAMQtIsV
aaWxysFhn6r4U4xb3lmvPz7dHQ4X31yTf6Ovh+zlPcXwjXSV24C9FrrX78rSaec9
mqFVGETXNxaMmbnx7KbVxa9xbPo6OeSrzBBRIpTWcd2xR2WrstSNtZHnQIzyd6aR
QIGayU4+TVJAnCC6xaNt8HLQ+07BY0CBBw4+CHTBSK1S84+OpAs89jRXsq+Ab4YM
EUTXOfRbWCNX0Ckif1XWxzORFygvb+WuNyT49LovT0UfLRiVACOEFJS64oeQo/qm
S+r0xa6BcPWFS5BCds0je/ql24rV18z/TbG9RS/zbdiospvk/cg0TBkf/1UlwQ8P
R+JtsbzX4/8/qbKZWMUo9wVlY5V+uwJ08mOdx5Pj/KPKLD5g3BGlu+Rec6YXusdW
Hvr7H3HlHHSiSKr720XsicbydG3jhj4BzIs1e8PN1BxPRT3shubxTNLGZDLtYYO9
FE1Wnsaus2pI0DCEbY2FDvEk3IEehAxf1vrwBfLBnreQiuTmdoRnDyu6lRSrw1pb
TcwkOGolrp4PjEACbTwWE1UqJJ9R2APGQk5NUtLlyUsOZP9L2yPTF7+Hu8Y4qkeA
vtjS1TKD5JZ+qtCmXDSMrY2ILeLeAh3aEVQnQeuHppEa6JrIqkOwvP8FEmvIPIVs
dwCl4lBCY0iS6yYY4UZIeSw4JE5eeppM1GWjFks2U3JTeI5C9xYErtVGGZQBCVkZ
0SCUpCyOOAfEYL6s5YUIKIeu1LH6R3I8BiGdPl8bLe8o0jJz5rbuGCohM0AYkLCV
1/CS0Uaf81zOOlTEAimzv3NzOZ2bEzJNGiHsVJlCdvioMTZXY5Ye9at0/eXlnTFv
h2wT8RvNGWw6Zm0cGo/eudIyfJYK/DpxnLi7BVCT55uLVMYPKo0HKtWAKfwQBPFs
UzlAslNomT0AK23f9dP2+FLptswRdKJ6s7uKi9ABStAtHmFcx0iCm0i3o7RIFHrS
/6Zgd5o0pDvOGC96WsOuPGjvu3mw6P9tBr+jn2WoSqON7L8RxLI+Y1SZxTEzAUgI
TLnVYg7QCCXjR8/8BnuyQM/irGy4WAo41TH+VA+CAxgSV2VBQdUj4Lsl8YZ1/8P3
NO+Tr9JoJ8ImMtBnSyjb4ELZREXEjdzpGg7Ew/KnOdx6k2CPqqohBEz6OnNHsVU9
hyd2gQPoBppLrNfQlEXgiHD9ZnSIWwG0HbwHFqgG9rsXdceAXy8B/n7n/UPSsEUI
Q2V7ubLximbkuxjgGwZAB9BRvKBpWhE0n/OefpN4ifOH5UT3INa3oNgB9nKjkC6g
8Sokk6dH3hU2RqD8yYxcFFUTnZpxRPevPWDiprqikidX2738se6mkqZWFctG3DO0
qn3C7XwfMu0lpdzPLLQylL9KSc7xhEyVLj2nGb4E07amSaec39pDNF+qk9/3YPNX
TTNpSjOgylqCRNpj2Y4XhZOLgEBF3zTG+UmSFY1r9h2kt4kUD/oa2hvcLD1huF1e
J/frV7tYO7X/vYpBJsHn+h3Y3qhDcJcUxfPXzc1YGf9kR9hNiEHVRdlmo1FENHhs
Qvb/b82dLy8wtWYNC1K9W7SW0+fvtHIWUeMYpCy5fV2B/Dv8zVUTINnPs5Rp2eHa
ifFdFxrs9UEpFsv5nH3P/Qymc0udKFPnUpRONI/OjfjnipPHU2d+sxL4ic/oOnWc
bzvqiLqy+jsUOUHJXke+fzY+3Qbb06nvFkIxCVJh2yYsFlvnEpk0nAEwkacBej1m
aB1PNhgZPwNQFKOAw2elNBa63Jz8+HM2sksB1XtAJFeUDR/8lLUlC/PD7ImePR+T
m+tUxaXihd+VweyB8pa9XQMhNlI989Wcv9aChdWWjZyQ2EvOlbJiJWe8L1eD+pZB
TCnPKJmPDLIFyNjxX/ntuyNugsOG2c2MsbMSJ15IJnkrRP5aj+Bb7HwCvbEbx8Zk
avaTckkD/7pqOzLOKZTBHIaxWMkNEGrUuCt1aQlhVerj9LfxVyJmDQwp8Ml7h1HF
JvzscKvDyjE/G2ulyh2K/tgvjZ/rJ+q6LqK+BhWkX3yadZJlgPLYvykQf4wBpo0t
c/E+TCYofy12h/AlPpWJk/IdOnwF4R9uzPtWKtkE+vnZ50whl52tqt/8tNv8+fo0
vFejO80B72g8f6Ttml4YbUCzZLAspoFCS1v5SLOTU5c6PQvE67lf6F7JqinvqS3x
KUJMxioDWBliNLwplirMfco7Ck/Ech/0EkkW7TjbZe6KcpjxjP3bMy3lMpzAB0+l
x4TraIqg6O74u4ICcqC9wWTYF+aefvDweT8NZfl+/ZtUdi8+SmRJbtQ8DtSzWne1
Vs2VL3aZLesQ16j0F3s2WAnalabuC52ieQc7FDLHOpxH1m5bG14IAjhimJXqIFkd
Kk0VWbRRuxK+y/s9os/4A4UgtiQzqyBGH08qHvCFs4PsPFRF8NbWBtbtaeZhJOxS
6krfcJj8CMgTqctDW1Zs9HXMk9p3BBon75XQ9z2Tj6615ZPLDiGnYnbsgh8teY2v
Jb6MlM34VBcen5Yl7UEGrGv+2PPybdoj6CC3TPMPhcaeNqdrsizk0Q2uz7AUKGKP
g41/sxoaltmo4ihP/k6tL3y6+/KizyW5JyJPRdSN5WGGTGCz16/536Ow0xUH0yLL
QX3Ffi/C4VTVF0pOv1w8zQb9UzZfzIs3c8OaTt/fEhszGw+sC2BPsVeRyf6Fev0o
jiWxyW6pSJvWCdphXJPSWmhADA3bqB0Yn5VsbcGbtBkZ+h4R3razJislZxURkOUB
o1+ba/62ojJ3t8AibRnI4PHyUXYlj4hz9xhVVPjYV56yjFIeD8N3SEf6SahDrT57
9TdcR+aBrJonuA96eiLvA3En+/5aEhrcptQ16Genwl351N0/lzlC+/eu2/tZYdBT
ZquRjmNIjtOxBeTeQ2GEWM40rarZL2Qxx94lhp+AEfFg1fjUXq4Bi2WanHLUK9xm
4DrJ59foxLd1RRziF1MBqGrQLKG5OPgS5NHLnx2I4R5W/fif3GTktF18egwFf75b
cKZQ01SgtbiDdLiw0eC0PG3JPr4FIxCp8eqGOql4UVC+A8svB5t4I2E+g9hYCTi6
o9JMyOIvCkNSkNGWyFNC68o/7povJeYFV+tBjbJlyc77FL0rWvDL4dwlUJe1Ewrv
f/l3prG4IOjsrckEWygJ3tG6Sgk6iQhPWld5zlLESUEXEmjki4yFfCP1waSm2JrS
oS2BkGeOwCyrIc3Wg7N4K3dbzQM4W4cL4kFhaJE6WRo7lqxZVk4rVBbAA45yWD5W
ybs5jDrZfc4Y9XY8ikmvInqal/0xvNqkp6TxAztlnF2oVR12ejaNnvvs34keQbCM
4uTF3hX84IWZE94+AKG/QrjLILZsqBDCBbu57i6SxQvoWt5mPIxVxql85cIqyGBL
fYTkRx5OxD7xhst0aJjtcZG8SXEHCGVc44zTiltiFWE7qqrxe6z6i6hMYV6rcY4D
+VbsmyDtUGUqQjogHWs6a5fikfDbJ3nRFqupRxW6uz8y/fosxtO4mAdyYsUv261O
5X9+2xiBdb62bsZ8PTOmtz6CjNqiPKqSsbFMdfLSkSUMaajttpV2FHAS9LBHLysK
YGfIXPMeF8HsZ1zuWSzh9wwIsVSYlCAz6HTXLugWoWg+xpeXe3s6XGaxCzuXU4/R
eZjgXLmvE8VaSWJf5LhmnecTFnPhQyDYUyiu0IjK37WLd0gw5MOZVwYAog5ztRWu
mXAdIKDMxUbJWJoyWAsleCRg9SvnqnMEdDGZ328ddaYRz6iafRidE2ie/OYNw5fP
G7tlJXvl2U6QqxgL5Nvnq0qP7bmwyJcDTKcKitCbcq/ftlO9on4G7J4NS9muoU39
GEEPXmzvgMdzCQQYrSVAIYKmP4v4KFg8oPPYfPaTQ3cOMEDgTbPEyL5yu3dZRSzc
eNGuOF6S174DGsRXmBD7VDmHkqVA76U6UQHEGSdFl++3tRLc5n8e92hE499yh4vF
SZFGStRvuUUr5UO/fZIcOYlEko36m0+aNMEHXacThr0eV4Ba65Wg2YxoafheV+kN
jmWE5LnWHh/uCF0UKHb+URHrDnCUQ7deDSxXC/vnC30tgeH/YVUxcu1767OkvQo2
aTxGqA7SGfpTtId6xUS/SYQS2afUe15/VcaVi18kRCc9GXqa3Jh1O0THaB/Ziq0o
qvfocM4/UaFRHT4ClZtlcTBW86aedTxic7dSwWwBMplJFmciOebzFq3xNLLHPCKN
tng0QEvvro5KPfOG6M1vFt3P1uBxgMy/3LDj2ArI+V6i38QyEDbzR4bD0TmyV6HU
dIHmJfNZJL+3WP4UeSG44zgvFE46MqCtrjKRd35fT2CrSAAXR2RyCN/F+JztvXNd
Ih0kQygnBC4jDuTGb5nx9/sOEiAjFeYoAeUiP0MoiXyZJsULOURUHT9zQf2af73m
tLNdp6cwjZ08+52s5QVAmF8qGVGjSBupXpN3kzaaEH4nMWqNKHbWWWodGQR42yQN
dkvxXacyyVD5YhotUYfyB4S+IhMfjQZUUf4AiM2GF2pKRVfRoM6Py3DqIz7e/qhc
RwrvBh90hCwH2e4HN352HMEWnHnJ3prvTWyri/9J3stgFLYq1g5vXfQROw8toxRv
LLqX0g6EUlBNpnuY43jZ2oSNXNlAAlHLRT5QvVIriCS3rAJ8jCexc/L7+ZD4MAzz
gYj1NOQxyHHn1UtuNz6WyXkTcILHlmyKgRtWZForkYwZIqSKDCTNVdGD2fTz1aPV
X5+nixDd9xl0xT2YUvPvXYPrmM0jwpz0yhnGhHcROK863ViAjE5vT6zHrGHnIF8G
Y4uYAEcf/7zH27vXeijPKvd5NZ1dOETPDl5HKTWQ6Hf7caPo65MZYrT3S2Y1hp+o
Y+1Da9YGCTeneLTIdL9NxW/g9JMCVjMWyQmuDPbkp7OTNwgvwOKF0nd829+0DgjR
lS+aUN8rFur4SZ+tjrwBCrMVh/7osfroNvXlBXMNhxOCYY9wnnoRF4/HMALGxqcU
UsNf1TQxRM4bFGsrQwjKodGtcb4c0bQ6mA1OigLBiRMRtnPGroRleb83s9dAOe2t
pLpWKggnbEPDC9jXIZjhWH1bzBgQwSa6/O0ivccxn7bHi+E82X/dqfB/XQGR0vx3
8j4sc9eYVYDr40Zj2KrSUtv2RXkPjdMP4+Q/VA2sl9Y4vhk4FwAMmEaupxDUcz47
BG5oj5GKCXh3eBKasJNEK/mOa5t9T+bkFGCblAAnpIFDPppEE+CBFizxYbyKySy5
AHgHqGfGpFKfSu51GWK3BDb3PkA+t/9zAf0ouX2nN0qg4UWcxa5ZLpJleli2iJHZ
08Vh9LU/NeNzWE06zQuoaNSKTSjXTlN0+YFtWnTTZen4xOrW1P6JtVX7Cd8gIcMz
K1rtPNSDIMkzZ0eKgZsVvb1DJvrrcfiE9TaIw8/SwYpHW9k04kYpOEd0mHs6ktZQ
59BLBKqxlProJyZ5g0uOEj2q/g1dItA4xrZ1s677SCSbk6AMBkyMeg6HvI2rtVBh
k2TqDfSeaYj6P9virrlOUovaof+llxZWvs2RM6zq5Y7KNgoyAjXztDMn7OYatgOs
Dhaxk8F4fHQ8XX6zNuoN8twSA5aRu2zhn0ax9iIUOFe/YjyZCjHDrv5OivfwAsQu
gESuWpLM9wZpUWFhX3sOXYIKL1/9Lob4utmRWUSYWxtSksGS3L54vMxcCDM4gXmq
hfppTy6rRQw0Hw9WSyVNL6/qXfNFKWqP3YKsA4JK4fasBh6NtH/Oy1OlcRNWS9h5
7EcHS7UeQgQxgu15sMpy5oQ/QlcyGZQBGPUhQ51zm4hVC2Wp0OAetjg6mN7hRVN6
jecv41oulZpe/bcMp51U7c7dwZCfRT2Olb/uE22Iet1PGGqjq8m1TiSgC35kl9/v
XIkcypv3kWXp4czeyhj/RvfFfBOSRrpij12nF9R2s1VTJegxQ/UWWh4H1TBHldOI
kA4xkI6Pwh7zHXVBo2oMHEqOmYN5PpBR+er00Ds9uI7qj/sQRqsZmnIx+KMh0Ixr
VINvmBYwolzO+Fv98XOtb2GRyk5S5AgNuiYzZrZFsOhM9AbAYE88tZGXDoxNjFjy
VkRizTxYPiIgv8blTFHSj3cRhaWz5kCFAC0AXIm9czCclJW+XxqFRi6eRxDKey62
4NiFaHVeWBu+vUkU/KCIDlMuHQ7ISrFSYjH8G5f8gQp0Pdx5w1xa7XbyYGcT1cp7
bbnH3UlObpR1VVs7Y8ZW+vO7EuK4F/t4xTYcKD9Qrxtvp9CEpGT1t5pAcE1JjgdP
EKb6Ssw57RQ/w/1LDtPnGT7a6xxEtEteX0r8ifrhsDA/pTcbb7/Zi9RgAdk94zDE
QJhCn519frXUNLJyohkre5xlcSWEVBBY+AB5P5xaxVBnen8kwwzQ47phJDYSzvDX
wBjTI8/slinEKsiu10U9JEh1fi1s029GPiHxM2VgXMSVcJio9vKGSEhC2D02JaTD
qeBXM2AgPdtWT6rATLSvLNOGBPEgPlfhdv69mh4ocSKrxBoNez4evkV8Nt41LOTZ
6xwqmqqONZ+naucsFIpqCuvZS6TqRaQg2enYlFNs6L8mvOu194rpWasTyc7RHKhM
WaXNSnH9/NxJTtjW7kwWj8HJHknvP9oRhhuaW1hpFYcRgyNWp4oEGHyEpXI/Fpqy
ttdAqhCPkF1YXGtxXFvyTL7jSKaQwv4QfxTKHPzUw7PKZRpMHDzJIiWBH/qITms7
T7ods0VC0uaorp6JTW6tm9QEl11+UDZi3aQ9fNaydKEra8l2FNQuTwdPTY4MM6S7
CdPZSXJeN1ze/xDpuGr8rSJ8dKhA68Kv7qRWCWMRtjHc8RGHWgmshNkekv9BqWJl
VX9h1I+xZVqOn06ozCHDBjIvqsCM+3euZeuy7WnHbX/Y11nymcLOn7gIqN3uzfRR
C9g0Yc3auKqpBjYAdt6yzE1D/5kWc+kxGPgNGpp/5fDCZcQNXYC8MTT2p9V4K5Kr
gDR+sFcWLLqQ8994DcFwwNlYaCY9F1SZouazXuXvW554ownDT3hwkKQdV2gZ8wo2
tSKJ16BFAwP1c3dxrQWQJy3TIW/TgXZYAWEgsXByKbifCXMZQ+PMjdtffedHg5FS
PaluijGxbxd/4VzAFQpB3/C50LyjhdL3fnddTTLoZzMXboQKiD9yzDoAcBrsdpeH
9CgSaB7n+fVex+6+Squ+1nALwecK41PsEKhQ6zeYKyFLrKpmgK1SEzFeuirSxqh9
F2OWBjcZM+XjpLVbH+AfzKYLEGLAUkuElYjtrR3I9g4nWzSJ3EKKMPFJ0fgDWJ97
MJ3XAsNVFzM7gRLfJMS1fldVNNBNI+Dd/hoAgQ8b6A9oKqXs0gX23lFMhS/LCDwp
1nZ/f7I2O88kFMMJfaGUwuR5JjTt1dGOYvYYuIoyYG79ePQ4TySIZVnVZFCZcVcE
15GxWe2UbaKgqVlnCrgLy7bGr8sJFyrJI7T2chvYHmGzbWZge6IdK9ps3+HmgxYQ
cfmsO51iqnaXW4zcHubOvXbqNqDfEE0R5j1seTXqEldNJnnT4agHm8KgbkbRPfrd
Z1+Mwiw3FRnt1KNBlQcni/jXySHTydeR8X3d49wN33oesuFVDN2PK74Wb6DBc+bN
S0+XC1ZORX2Hi6fKkINFj/GSDNpCnVmi5PfEUVvEDZ1BbXxfXZ6KgsWrL5SHE3O1
ABXh3gD0Qbi4W13Bz0cHBgXNMz+FBfr5Lth9o6KLb0JvUN7eF/xl5LzmnA5UqpI0
bQ8TMbo9RRPUpEp2jh8oDnLIdVBsRmh3qUVsbNpup8BRq3HgCzEqidU87DkRYEm3
y2lgHCFYAyH/C+7C25eSZszqFkLazD1lX8K9743xuQc6XB2AtzQ02Eq4zgrGOsD1
bDt5Lm12OABhpMMnv9e1uGQwefsk3H3K6aQ3SWdEgNUN8YcjEGvtiYMqyHwg+7sm
ZxvSdkclKGQi4xgBYqIcilyBLAhSd+fIk5m8vOExhAyJCYoU5nV6fT6DI8UUZbE5
fg+1FopQAUszUiaZPRFUMyEq0i5yoGsNUk2fsj4XUdT3VFVG+VrlBmRQALEY5Dnh
tKmv6ox0rqoKrm0cQ0V+i/LssgN/LflzLsDQFGNfp/sQWjmU4op/Mtm0+Eyi/+N+
LCGAkTMX00qDWkWuAzzBdgDVcY21Rmk4oHzQZAv9O5VxSED+VvirOFyuEHmlwHuV
DGcjQbGehdz72MIF4yauiPStjJ+IshgT6UQCIm08L7NenpyviCTixg5vx6IzJIBN
G+Frv7pK49XsifNCr4VQfRhby9sreNk95rNmSf4NWP+X7NrwaKVwwyLKlhKlB370
c+1K2rmW0ezTcMB94t3INbONd9lCtHeGl9cUtmW8p09f0DJJEaCtxhDluETJQU8T
wB/hwHwcvEygVFqrVtO58v9RxV+zAd1ZEJVvvxdiFtNOs8YhN6nMytRdhg55lhDy
gcU4+7UwFCvGdVoN2ucmWKIm665ZsGEthcQREXMyb8+auo6DuZherpnnmKXKGF0w
CzLqVyxxl4wXLmHZFY3fYkST+9MKk8/+3++k4phffWJ8WW39/YVm37mrFb944RTy
rlMXqrty60EeZQd8oIk4V477q0ywqBKjes0qgB98BYddmrgogTC+c3exziwE/1zE
ZDh9JoZP8iwDRFPZroSRw9tU4LRLtes2Bsm46kQkH5tPDifsVrAeUKnaWs08BkFZ
2YIm/WQrL4tceOpciu8QQIRon7fHq5n5H+0sIlb0J+z1s4gvJz0Bh8lpNP4SZxST
9DSXTiAPnYOuyay5n8HMYK+vJ0ET6BHB3P8aLmxz5Fjito8iSwYQpvsJQztEZlju
ZNUgUfrtmf4OQeI7wRmZaU2qpkZG2SZOGP23rO6Sqas/8u2IFyGrJMOtGhBUwPHH
i4nmjEAwklbivh/S/zsAJl9z6GzRNSC3XEyyya1TOnZX3Ow5ACeIN+y4tR2/JlMk
CvTfZuWM31CqgUbC8cJtxbfdwtZSoXgugxJVxAOA+1C/jt221yhIlEyEtEZlc07g
m/kfLnT5f41fSfJBFSODOdxfrudVxB7TKbuFbfMk3an869Gg2jaQg3DvmFpjzRJ2
KOhiNhKPf9XNQZm255HZtnNGvS7FN73SueE3QTjMnxffEGfUKDv3UgKuaLr5ka4k
sB0JvMeIsHwIddEPixoFhO3RsMAyhyQroMEKY95S0byMt7Ho3yUKLjS/HoOMkdvc
T3eMw8rSeG56WXdDgYEfpte6kxPLnee2yBgD3hcpwFTZJV2QkFfx2dusD2XjMNup
6Zj7uTNdNB5JHbfuNT5dk3XPznuaOkThVvA5ULTsAXRlpwZmOSQVAIAULCWgMFjE
xy3Dw5Mz76o7/6b4giL5ASj3JLQz/7CWsBZJ/BCxLtPJXYxnr13UfzmoEcAQAcmc
+f8a1WHCO0L0w6HqF9TU1oP6UUOZ1qe8WpfWY2BgF3y3rs3yRIiCF5yBlqAWs/H0
m1Td1iVmEi7MJD5vRKWizeZcdhKOC/e7hykQ8iw14kxLVy8f6FeUSSIHfpGfdDgB
l6+X2r0rlH+VjF8xO8JtwpTr0r+tJZAyzPYwLZzyi3U8Cj6lB63uSHe/+wwl6+SL
niCkJyI5LtG/oCYwayXxkGeJVuOJzk/pu3aGMmqFf7lYA0PN2lsg++es7+1g85iX
yPdwDggGmAXpUSgfegl/vdQi5Ytq0crvnpV/+XlYAVvLmfmDFSy1xQpYogZjMbF/
8a6C4kLa6UMnc/9ua2qKpE3mt/UZqQNau4JZzlJba21mywgNnX8SEjiw49CFu/eX
Es7QeW9lY9fn5Q3ki7YQAiFl44cEBoN2NAJ/tb/twfU8XVU7vRetpB6eEWYn2pZ2
HXf//NoSwgOnGLFeqk2UMJN8ZBz5VT75/EaPjhg55vqWre8XBzCK8F+onXeij04R
gdx4MnP9PtgyFTNu3RvXi41PqvuK6aM4tSe+XPnSEFNZjkELH6v0hcAFomRh2Au0
aR1sZ4EPsdhZ6FOEI7w1x67USqa8whByrjerU4QYJ9IjeXNUkzoVayHXoZw7hQ9G
+0ZBE0sBaJQ03Rsol5237C7CI2RnqAD6FkHHAkz4teCZm7pbvVs3Sl62qd99HUsK
wrxK4PUTbhifrOCLvD67vAGQ5X8JO3ok1gb/hkUuVMJ2vTyf/MYnTu9GrYYubjJX
tz9oiaD1jODtWscoI9QOsouvSILO43jQFogufQ9nIXjEO0Gc+xfTWeDoY1UJBLlA
9fl0KSZK31RY11a4IiBYjRgFBReVhUt+nz/MPlCDc2iJxENadMWAil//WB8M50f2
oFJ5SXBtjIPIKC26lH2hEnwHLNsfCaoEHdvsFH60jDRdxM+SUGHvB8Mn145nr4qm
ZhmkSju0oHTsLb7SSuKAkoGLSTycykK9sExJz0qjR+pHyEnTdaYpKnPh4oG/ca8Z
fM9GHqlD1Qx1+9RLhzKeB1YE20E1iyTZv7Gi6DD1WUK/3roRbjg6DJ48F0Hyc9At
GpXQHSTJuVJGggnHbo5yATXbY02oSCNalO/Qw2PE/7omjotvhru0au/GpLoPcQOA
nsZvLBDswRiLtZg+sIYr2j730c9exRGRWFFAW8/yKZXiPwTfqn8CSmOnf5bSciMV
8Pu4jV0/L3PbBIMS58TOkoBsBZPex9MGh3kUIRBSLOLLPjUUxO+bq7M2WvW3m78n
E+YmesN5pNmnJ4IpyMPstU8vsZJ/79lcgbA9my6Q8ymO1GRCGYQZHE/pRRvgbEDm
uFUS9P1aTbd9gKghWEt8H1lIgebOEFDWedvSoE2e8eN+vNsRjVxBuVEs13OYIijV
9rWv0PNv2vmTYBFH6FUpu+8xu9WQfdKXHKIuKRZOpDVdQ+TjsC6IoaxdQWrIeACa
wxtHFixx9nCzMa1rgxQJTvb2bEzBsNzZOvsFQ2QClPTZ/i/7A+iV6egzb3uELN/N
OtmwgGuRIAwcSUYW2C65JXQIxkJeX5nZN8+U+ia3FJoGTFm/5tU4kHUvqB1bRIbn
xhsqv4AM+4/A2qY7kye5ruW+h9pu+7GGtdSJ7bGNXm8+DnSYlgn/6dfovKLNkSZH
UaxrXYjBwsMo0LWJ2SOVl+UgENhdvXgh5/khiCjXwdyoNZRQIdh8Qc/Y3d10mhP4
CfWXRydIrLoiwDAvDJ6n+pLbn89WyD9PsyxOlNXWvX1N4xjZDRCR5UuPD8CnzX/f
r2N+JPbuVbdPSMTqYjhpYMlHd9VY9HyU8s8A1TfrT8yLmguTq5Jl4Ao14natbdB+
cuw0vDD4gq4Zh74zijcqqx/QL3seNLkoOKInfDzCh46+ZQ1uiwJ5WyZDXqYNdxo1
hQtsSn+N4nJzS4q3S7SU342+xk2mhGMWJqrnhSSIo9GMD+2GXeEc4N7ZuM5jOcNf
UUEyHEsw2xiHLH0XWIZFSZFK7qVCAUFEm8lRFhaVMMeiZLyumTwC5q2bj1rUIT3s
5JaD9iH5I7Ir4wulPLDUxthDfslkF5/2257y1YCl/gVhpj87gYX9MfLcL4g/QD3H
cFwCB/nTdFHf+uYemlMbdoJgeqM4iNVnOgtEeRTLO86VAbWgzcJFdmTCq+94KJxe
QEzURfbeATmC47LZ2UhtJQH6H+bakfJBdqukdfrF1wuwkS1rk8/JTRBn1PhRxV/D
jb5mlPSn/mZZYWY3IcTTc2Bay9U9uQ7prZrLmCy11YC1i3hw5UyTHvFEKT2WaThX
u7Q0yXHtF+NEU0PG1/GFyNeRs76bvRm+4fCG2qls//x5/DM4dPLPR4cA/4CZyRkR
pCbVRcTYnTEHPpd2tti/gE7Af84bP6ns0B7r5oLzqlPzRqEKMjU1yseWIwiS3Rxx
QahKNB+F9iQlKHw1S0Sv28tZ/hVIeajE0Pu+tQO08uqZaFHDV+nw07F7rlNcl1ea
cvxYOaZYDW/ilbh4BhQ4fhoxs/F0IGgrafgDRymD01RtUmdQOWSJhX+rq2BEg22z
YxzSlWkD7kafckn/BVfGTfRGsL18NWuotAFl7wvxdGVY8fIkPYzLtrvxE6L+VqR6
iDdb3WSJGjX6Hl1v+Mh5u6yEM/6O0EQmb4Z0fzQPm0j7mU20fPUEhB44IHq4Ht56
zGamZYDF/g+KzZU/TA1i0/+qPVw/QhAiEM5RBKm4Rhjt7abRu1RJCqXjAV81kuas
RrOFfS9Ceu2/S5g9NoBxFIO8bOpenClt2hWyl+YFW9jLMOHFHdw1GYnRKm0yRy/2
yrJqmoxs3CQIvbo6pvVmMGuLH6zI3XXUoQ583Jt8TQVBQzsfTudo2nu3WmvwAt8G
BS/bC+4I0fXmxQ03qi6d51OIGLdOFsmzZut1XJN8dtQRVtzArIfldbKUdSD3oUXK
LSRffraicDPpdhle0euihL+fBHf6GRU7P4jEIPAtvAaWV0efhlbWfLAa3/0z0R2R
7I4f8JwVWTswHFbW2iUsPddYZIqlNGzCmCMGM5yhlh5X02kpztfWAaRw9+LV86d3
TvQIyAE3m1bcm3p1RFelMxtoCnrT+ZcMYZvRH6RoDP6MMaC489Cm9MiuIYzImP8d
+y94bX4mVPW2qlGr/WeHJWlZ/y39lG9xbSkaqB+ilZLbW6bj23R2JaotNPBB+un9
KE32NqCpE+qHsSrG7Jjd8kZ9EgjhlJ5ngMjGRXWbGSFvhqNeitZxx5HI/MQURo9j
+I9UP9xz0RrA3B5Ub/SiqEWFTS5JPFii5/X56IetSwVeGmxs04Zyn0tiZWEZqQ+c
2MjABri4YEv0cWpZUB/uLpa1zxR9eIdMA2A6Cg3AHhr6lTAVL++qY1vYoqTgFkDM
QgbkZF3jc6l43pPhh0mWrf3X1aKSZAmQlxexn+TU4LirDCOCQFHR0nbVqeihCk33
4YzQz46x6alQWljRmLwrwaHLl4yJS6j7tft1gf8J16Kj7R4iASEbN0yXQ6bMDyMO
unKXIxoH8aCZs95gZK0Hg1YuoYDwP5FJIK5r5/xlgYyVchv1p5m0pl/u4/FvPpsa
ra4bO4YwVJjCRu9tExvL2ZDZCUUX09+sJxnugmPcsYihhFH0uj3XtdOKexUWqMRu
2L9Jjbto98Rx8GAXkogSEIaUEt5HPKLbl8NPJfSyk9UL2i3k/lwSC5nn4sjb2yaG
qS5jxW95TS222nCzjTYy0G03k7mXffXVEIRP3iqznumzVY5kxOec2AkeaSLvD3Oh
m4gFTC4p8NjSZE2b95OteCrL/i3nMHDoaLMOCq7PRt7eh2xmn/MjgcJegk2s3Lrm
FXKBPWWI47Ds3qA64NArs6/i9K9fEXjVxipNGa1zONGN7rZs8VioqxFN8b70Gwv5
Fh2FMj7RCBHfI9WJ1VHsCnFjkV1yBhXSqVRJ4LJ4+tlZWJbWLvNiSqw7L98lBPNh
KvvXHuXIyk4y3uoOM8l21CR2nhVvK00ZU2lCqeNWgXwiusDPPc10tgpFdq3DVB9N
uAwQGag88rLDHZ2KAB+DGpewTSWaOYFbAwMaTHSkZMxP3QrRHJEsKcAcEKlGvfHA
IZxhqqiMWYmWcCBo4fm4ut1VUYJY0v9mFGR0ECoolMEYQ4emWoDXZpekOx4Q/0h1
pnoXjPWht5Cn3DiVXYZ2+M9GkfTUH6ZkRTY4DtJWcsWph78/UBNldnz4tLPPsoMG
oZPYhE6OxYmVeGCZzDsL+NoTIt756/HAt2OFMQS/iwqFEU69RW08YuBHAaOKoMdM
YeCC4uhb2CWaGZqwBK6Bs+ixNKN/y/OpYCf0XeP/ivEUwgIJ6WtZsv5NLPYuDLFo
r7VBeDDQ5MYJRttDLrKu5K5ofiEnoIXEmA2MczaUWt3kB4+9g6fhre01zq3z3XmD
JfW0RI7Tb3xKthIx0hnOlbQ+v2STksAv0fH7sP1Kp4i6a/DR5totCCg/LMxtPh7g
hG5GAOqY8awatzzNOt7epUwb3FB89mglVLzBqiX2R3h2Dt2WVoSA3VCNBdnCjisX
/ktDhLvMFbfQIF6n/InyTn0bbsNvlhAcer1cKUkTZBnc6YQ3hSrecqLbeD1Os1Ij
UJPZJR4tcsgDzuPfTbKThaW2QIgVQSle1JYODWQjw0zWu1DL9VO3tcIZafLv42QZ
LRW1Xsla9Gs5kXLMzM8w0kb2/kYfXV77r0ryilrA2cHIUWrlgXt1q5l/R1HFfH6T
ES37Ge7TOQWYabfTqy0qFn8Fjhik8R0Nra1KGmgDTSynCWCG0iN9ZhbHUxyX/TMm
ryEypskLk9jMM0dlwtOil/W3boD1Vf1X2V2W7eHpr5aS0B+4HkMNLlAfxijtJwi3
ujygNA0PZb1WlgiL5IkjoOp3HBdQSS6eIgph2ruYwwD5/XYWNw+XUnSnsm/Ekq8M
pptAO2cYJrc8Cqr+lJ/XoNVRgN/l5YtBV7G13Ta/bRDSUXSXJ3IS2yb7/1J8pBNL
YjTKozz8mBVjB/JAZ9ZYE0g6gmDcNhzDdUBmgkhuxuz2H/+UWd7PgKvfKCCFh8Pz
16BSyRitxH1qyWsv/jjChimgVreouYiQ398ne+iCS3CSCSnpoCkzuLSpHJyDmRnG
78CyzR9GAI2lam/QQwNdnwM8RcxVnYktrHcGr95saFHlpsJm8Nvq2dqWJsV8I28A
xs8WoNZiIl1UgFHF76ZnAbC0SBuv3gZ1x2V+PLvPHj8vJTRrIulgtZ6MeFOxZdxF
wnvU2qCpJUAUM1NXDj72ZbzLbcqa7GysZks8Ju/bGK9LY4Y5ivmMIdlAwbEnhGZt
tm7GPHg82VZT/+qkKKrUfhIuLmB6wtIRfbtndPav4Ei7DEdrUUJTwTeECoEBF6sQ
oxLmICWZ+SsJsu0OADtSfIkDNP7H5FfAd2fAIQe34EHi2xi6HjbOy05kRMagQ94T
tvdPnAowFDhfovstMDdS+clkjKaadwAC5ES0ee4hg2bE1owzMggEecG90CJpFign
Q+w2IBEtL+z0qMiTI4aUum5xAUsOEWU4oaiF+W+XKC+7DbHgX6+HiaA7EtGUNLoc
0U54+rUPQQB36GhKR5XO4JpgAwZx7kQoT858ExKyeM4iXHOqGaz9n9ikNnuB/Gn6
nBabR5TlQm1BFBdx4KnezkyC+LvcP5tIy4gvISrk5HYr2wa1qTeliuOwPwWZhADL
FLV8pLaQPfz5iyYghZwgJkrTGvy98f6mXWKWfANXX2eSXPBgQ7kNoQO8KREyzYs/
LDw2yjJoqFoImeTyi4EjPRzdsP31PCe/NL0F8FIVR09hUt7IUmBX1/0/aiJGswG9
bWdAN+yGhKqV/JQBmnNeweY4Hr1KITZHFBU4KjzmNIwA02wKWr27oVoUwB8XjDqQ
5g9oLAwa6+0wISGyNvANPm0As5KIK9ZFO063t6DnoRYPT/R+4HJeJfLiHuJnem9b
4ZsOaY89OPH55zHkfK/jKNoWg3IdYmTqK/zzfci4lmGSS2HcPLyxz9Q6wui4o2H9
U4RM6jozzeF/yVesiyCSSdpJxmW+TlzqZaUhPQj4bLi6BeZutFNxtU8pyVX8Pr7F
+Ux/cq+PfWSXqE0J2RAQbmRlYXhpQzK4MJOpppg/yXeieSXC7LXZVeOib1vo275O
DKu+kkcRFnz+ax5Hc1M+t9UK/pEKXClXOq9FRs7E1Nyzx9lCXFKVYhJefV3/b8d1
Zzjtv4jnehIG1cftF54KODp4hO2rb0hoO7eND8M1T4ruoN0zxF2+sVLE1W5BL753
aSobfB0JGbQFgMvcaMv0eqayrgbNK1qKaPS99jhyFvUo5U0IG5a5hPRhU8CxMHBK
aAXGWujUqzrFTIBxw6SWl0HIoWVAK7UOJhzZ+/M+OJyFA7QoRlgOf+0XYBJTXsev
50KqZqxSp9jhMgggrT8hFNC87FSyrnBaEm4aGP+B1Yh/q9mnD/83BgRK8UptC3yV
eWUYdqB5F01G9sPvQLVA3zyyQiHPM9ScdJzWKPVNlMraOIv+rPiQSLqqIs+kXuQY
qPr5gRK5bcfSE5kcv4VjcU5/DV+oMFzhhJvOqTz7jtNZ8nJtyT+vLfsexvbXXH90
hS1SI5yqRxpjGz6JGrR4HaOvZuhC1mg5uexBxgiaUat8xqEXq2nyPdwRynSQeytE
cOVJ78U+PpgOPZOBPAvF+8kpxO737Ae8VJhFj0l6t/usHsAIncG/CCdHoPIDdLO0
eXR24WkdS6GdPsLWqG3HWrZq6RftxM38Ea8FJShU8fSTA/DNjws5XdSOWw4EqLB8
3HM6bjU8J5LukS2ASji6d2EAZ8gg9fPg6/HpzGO9sMMLnYidEaR/AMAwp2UtNInU
pd5szOC3gcpTAq7FONI0h5RAe+Er88sMSOwsiFJV4BqCWefXUnF2HzeHt4SuQ0te
TTet5ak0cK12uG02AneoXC7eNmI/9pKxTu+LskaI5oYlXhNAdgvVEZawEn8Xh5zS
Nz2sQhKg6YdBW1mNp43wAz+BPiuoE1r5Kvy/aBxEe26ifFGCO3CWdMdP7AEBffVx
q29J9pmDInM2nbawoBAOrGtFWkCLtvaxLMsNcHSKzNbWMRfskowq+EirQUplyaO/
eD8lfHsvThH2Qf5O2dRNYrkmxFTb71KOhAlo/CvsK3DkmBKMgFoCuf1g2DD54R1v
yjLuyHGVPGqTBQIJBe/TCOikopj/Y6F//pSun/yCq6FWSPEbZkF2+K34RN+oIw9N
ul2WFg+e2NGn0nX9d3ZNZ2sMeSGgbM8Zaz1mWgtGrzPXdcaoYHWzLr2ZDRQmxJdI
r4c+Th0cJaS10DHpf1pUUm3WstctGiKwMd9DAnWCERN7lVGcG6Deri+Jn1TBMxL4
kCvKu5cmi7g0gVqRLig9mkpc6LqSCXGpMgVDiFJdYW22Y7P9NlOsDZ0VrH6svarM
0QIm952XKPCUsPBPTjlNZB2+7ydMhEzT8R5YOVxKBn6AJ64JLq74n6mV8y8ip7k2
S0nTJvThEfqnlyG8UGSNbs4lHG1EXaneivVKDJ31/1BjAL+3Ykidker9lN0FYlKf
s6W4ewmHVsAysBaNWQyG1ggJv2jfzUNcYANz26Glyn35697ECJIdyIKK5nsy0Ccl
Baz4K0sNsEamRp137HhV2+HZqTf4gWUQsVwXWp02Ev++0zLcmZDZ+lIsyKq2i3LV
DtTjyy9G3RyNv3mTAv5BsAkZqW46O5iFlOQCMHIRiZsW8ExGCvGxaI4zAMDGi4Je
2gVwFAIi/SmceEAO6UQ2Ua2kgFq6+dUGW8fMmOAoxbEKDt9QdarMtzRBZk79U+Y3
M0t7e/oivGwIbrjANz3ZHxHmUwXR+DrZ6pUjmu14+VHKk7coLOCQZT6A/c2RpYGv
iemXG30O1h6N7FWlp36EvUi39WWy4JcWQFOVOWE5+aQCIwDdHpWR1TEw8pnzkpSz
0hs6aoeNDgo3GKACRVYs+X9dKgvNugiQXF15deMC5tu8pKoG0tvLQDvST51JYM1+
tjL7GkSHC0pGsVnFt78Y+gSBlbCSdLRGaCrmROqOPgyweAt1CwEj6j1izdA4W0FH
m5GpsO7+72k0Pw4rI1hyLEhf6phiTwwYK58zFlO1rLeDUSq0JrBkM2MzNCPzeTMv
1arKh73+kx+KNR2mminPyO4Ccw/pVhuerfD5yiAkbffSmfGWdjqDZE8X5EaLVxZx
gDf4HZvy1Vde/iaCkQ+bUuLPQ7Y3g6QCmXtPOcp/35wiNe+1X/hjkZG3mPblX/yA
mzP7Q+zJTW2x6p8A9mHszLlAWG+Gz5DklYB/9tUkiPEpvdsztQSOzpd/l+X3rks+
s2Iqn2I6wJ1LBPEAWSU+9PE7LEmp37Fexj1+cUjUemg9qDeMLjxDOJJTy5SgBI6F
lXc2nl64KomoCycuw3whQD4H1TuSsvG4dHKB0eCZCmsihcjc4hoGNIJ+Z+Ogt/bo
Dz4hoE2hRBCzYSTTl6QhZDc3ltSBk7EH5BXUOid7ufI4lm0JiCprW2GlaNB0n9Gh
wIOL3u5KufKIfsEYYaG+gZM83dL0TtqTTYmi/slYLtI9edhKGw1h+7p8zJIWaI8z
/QpqOlRzdGlzcVGvwJ2bSD/TzfZGwbS1ux3oyb//4+H0EruFFbiw2SwrbDateL1u
BOFPpx3Xha4nQj1iHivcFpLYQdvC5cWG3cM3M92RFRp6XScbtonaCF+Itla7R9jy
IYR457rpxZHPsLFEa42V91olr/eeNVeDJserxU3XOn1A6wuKffKzk+zif65TF1HL
yolrQMn0wmZPszGX4/xO3fQaALTlf4BkvSn0f42/Sm2EGztHiK9VUHJJGIzHlR+E
HoJDn4HGR2x62baXX5/hP60nTRK3nUH3fa1F7qUwOrtlZK8pTbDZmIwSVo2lm0pF
I1ZUr2BfBgsXBhsfS4cYQgW/sJF5XErauE9H8Wuyzywh+ETRpm9hlhSrWmLmVypj
dwuysLTloT+qLTQUfLXe7HFZLWwZaPxATWqisuvGl0QWNMf5bDeaSEg+iutJrQ2Y
rVDPcX9BT+Ix0Js7gA2WNqiiwwEi0bfRjVLFiaEUxVIU3fsaQrZco7x4QZTpMQ5+
kkEHHjGv6Xmj/YbdpozHxVCt7MwY9+DIeYq+BRrkbayVOgTY6UBHlZF4ouWA46qv
KNuuqnr5ItczxzFkfTz0oJljVzEIbBAr3pCjEFdH+Ky7ViIop0kdpPMe/gga4DoX
C+9uxi/QrZIbYLvzmW9NMhCIOALvYqgpX0hZam4fJmKQllyIUb/n8FKjLrXiznFE
EJopacar0rmTFNGpbahOxMeyC78VfNBMfhZhBA4OETDGffCqaoqPaGmg5udai32L
HAhYLUv8jLpIfyxAdMw0DXwEcGwZu2bF1h/U8Zm+YXR6x1CNHd3lgQyKqGGs0cdC
582Zw9xFD9c/BD8+KsnXZGZ79gjWbnVokFiK559uaJfMV6VuxJmJzrSha+/qDRxE
3mH1z5ccSf5sdpC/Agw5Bmp9AAj2DyhkGDDMyZB4ZiGA4lAWBZKarjI8Wy93fLXZ
KIxxy/By4opHjNyR4G/VXR7rG95a3H2ues10eKKgSFb+oHqS8PIMcvjhYG6DPXz9
O0Bj2F9dbxxUrNTzLktbZZT1gsy644iGkcAtTVG5RGXwaS35AhImePptlaVVLPkw
aqA+VVHBjF2eT3kOh4DZI750YO6S1ZPXt32W/GHOzg8WwQ0URMiJXI1POQGGKDqD
Jt1VnqckIACFncWh221tvQIjX5lBmu3MG7XxrJ+J3V34hxF2NICe7uw6sBbEtXIh
4moTEb1253F7dkOlMcbUP0f8uM/6Vn/GmEGDgEBdAeG/oSnJ48qw71yc0suq6hDP
iicrxt8J2i4IDiotSlIacXVvkmO+vTKIGjagWaddTdaxTFKBbO4883LYKNWFtVy1
zt0UD9t6IK/X0PeFcwrXwn0UWQ8rdkfEUTZqZ0Sl5ZeSVIjZz8I1ldntdNKOlqEn
CH5oA2tx44eF8FFR/8hazJp+WqJ4YR9FClT+4874YJ2rOr6e9Lr7b2SQ9rNVXbxf
wGWt2aD4/rylBpg5C5QyzBCYjwxBVnxojpfvjb2h8dGZlZv8takQ4Plh7uGNWr3w
otzKt117dv2HwHLOn1l6b3ozPEH22INB/pw2pMcKRfwLQ5skVyc0jCZIFwkF1ULb
uLRCbrEljs6W+WW/yX1ANC83EF++6vr3bFYI3DQBy6KT0qT0mNwwv3smDMUPcopB
BvkxVvNIRHNRP84PMKUugdI3TF+OcDz8MOQeQaINSxjIafg4UjgKFdCmv8BptRtL
s10161AzxFwn3ftVSyj6aUb1aZmf5lN5QCP4vnKHjKfw7b7ZL8UuAgAk7IuJJHFn
ENlFk0z4DTk+zqnx/vJP5svw/0gajc3yYn10fcmh50iWt9AmaTLWMVRsbniLIlrB
Zr1gjSzSmafcxyUKtdTnnMyFHtChlX4ZJ2pWnYXumAL4qyUFk1LGupqvXrO8koeK
6fun8ds1hyNVTlet7NiNr9xcfDFjCgcG1fVR9eLKoa5GL3v8iRQzlFozyOhEYWTO
ABx2juoXRSxESOOhdjLKspvzWfFS6wBWKmUmrzm1bvzCHsCmn3DSv3hqijGrx9GK
7ZntYp32LRcBVicmblsh+NJNBJ3IP8G+7PVrcfaK2H5Ed5hssQ5Ku7pmWGjyF3cw
1M5SFIW3NhwWDvF1SaF8e/9ilvebuL1nrAD/F7/2XqTh7qMBHdy3udtLkqcPkKYl
Vj+cb75RE3hC9M+T2ltj6N+2k9kRlJFpXdNwd6D55QgHwxOgZfYoBkMgHo/aceN/
0AZvv7Lh61Hvah0oLe5HjaiEoTBRwmtxq+wuBwd82UJu0I74E7Ji7/AWfA+Y5/mk
7uuqC+OraGZEJVNsZg/QdH3rb5bK6E4FrMAWhZtff2WJ45kuO9twltvMmkiE5POn
DC8EVgCliWJEiTIxM9Tg3H0LLNe6uG71eTrl14kFGx8sOzW3hTPLk5BGkRBRrMK0
s1Cd6LeR5Qc208ZL16263aF8qPPpa3eotF2UcyV4m5GZdohxlr22z2zKcZ11pwt4
q9hGwWMJjygDYoLK/qNj98hrMuNjcQOQ5VAXi4hbpkcEfnudoyyrjj7ZwigHy4/s
gF8bNH9R8P0kUSSY1C8QNkNmEJ5l43MQIchSWmiWLz6bzCEXpxmgJq3zvZuSNobd
Bd+HOBLJPMM3RGyTUsEhCjGQPK+vptZCZcPkZFzLWkZ1JZG8uymlay6lFzNDU7bu
V4qWhfO/WK6hkl9fDCWLeFO+/9AkNzZe9V7iqg3EF7pmlqLPLgHgYHZ2WfQHBGpW
2VSl506npPHfVHdL1ych3ruBUfXyCaxy/izMfI4/FUMBBOPFK1TBfIzU4Lnp85U2
3jEVP+MIfCgrHxPnj6kulbxQclhKKYt7Nt55jbzDBv7ocKAfX5PNrlQd2wixhocr
ZkV4YLWLuUevIEikcL7/IJS+z7c3uVIC82maDh26mtfumJPYToGjoof+131Dxngi
oDcf9CclaB4PRWIE52HQCHx9T+JcPtXYzGu0hFmokXX3tw0i5sPdkGByrWT7KZqt
z91Ih/iHzhjTHKDilJrxbXdRpsEq9X59toabgY+yQvG8SUVDqzbiL02rKErYqHAT
eaBG/dMEhOUsLsradYhiBocAJuBgEIHdTYScMeapDiK1CH9J/sV+SUC+VKPetA/Q
uCyFJ+3cN6qhUz83W4/7KB3wFRqqO3q/ciRtckUs87ub9GxgPhzmso00ZSyuabos
mR1kC9DQk98q7JIWOF5R4bgAN+bAi/0ZTrr85wDrwrinF6KLgSn6q6lcuWGIjh9+
P600ZE+WD9az0BLrzw24rDiuTh8hrl6hoBeAc5tH881Cwv98AsMdsgsB4JmeKL2o
gQKfKmifbnYquuv04LcnqOYtHzRYQ54Ms/SlNbKfW5mSKkzVcoNFIaSFvCka8DwO
K0glKcFL7vp5SgbWB8OG6twqUBEYrZNskktDPnrzcQTzYXFJAvfD8Be2uyUA6Kjv
B6U61DED2UJ3Ld63y+TlC/1m1jiyThwY7CLW50Y/0BzsVr9CON6HPGUxZifv0cKt
F0rEG3QJXGyRvrRfzHZlmOvVoNa1vZgnNUYzO9ebW7yDkwHXcIRuJSvRe3RFe7ne
AlEAdqzrkOTxIScc+NBrmXA7bBU5bcax+m1g/hNjK44UkMLHWa5SLzrcXHSNM0hq
9Nvwh9xOn6grKb8h5D1tJMyjE73l4rYb4nSwIpUyf7Nv7MJ5gNHbPcziZxHu6NYP
wBzRbVAZKDbwnT8Y0H1NpFZMllTeBCvnn8BkuUxsqU5CNSF8g0MDZ2PH9WfTDWEK
YL7vRaaI/a2+p6BZKl5KKZDNvhnnz0RzVMC/7Ym275YXyHVpiInB17b85mPyRJj4
/aX6pzb17wqfKfVkJMiVP/IzKMqVMEAdch1Pnl/zzmXPz+tqliQtZzp4hK1cL35P
9uWfJKbWQGXAejK7WEYZhFPwYO9iElmsWqyCpwiXyarXV45kUzKbkT01TlEvnknH
gdGqs4NZ9sIDARnNPBYY7ZqlIxJIGzviaeKelh+dOqUwzCdhA7cBkrnqgrfBnFju
rsoDLTFFI7b/i1k2DXmgMT/pRU6D12fEBC2ImPhC0GTS4Z8dvjNqzt9WFclmwq1k
LHZ37HYJ2vxRWzVaRBAuAlygc5/X/to2x4/6A/m2UaARijzrFhyI7a4deq1kr17z
yURHLb0nKPEo/j9sN1+kcfupMj0MM9dlpmA7RgdfSaHffA35FOFR8XDkTGSegchZ
X5Ai2RI/TOpoLfeePASydHCzGsRvmCmcII7BiixQJ2COpsnkG6JB3Z2CJDa4Cmfc
M7Xu1HWJef4Q/y/agoCVa0NEOu56EyKlNzfQxbl1/3xT4cqr5HwP6CXzoUFGX28Q
OQ39Fj9gc9eaIOlhM8yoMvR9C0PsUToiydfLusldFEsAWPbehdJ+c7hia+bpcA54
MvMqu80GreEBm2Xbtz9BNV3ohDvPOWYeoogzZe/mXzABRskuptOHzO8rP6oQjxw0
Ua2+cdpxnJa8tt3nbqgy0L6ZFNi+zqo11ogAxCmYfC7OItpSENbQcPhTdPLj2f0v
8qrfx0p7+l76I4NOgiHgV9vGjRR6UvW8R7Q0sxM9fnZPP/8Z4fEL0Zd1A/toVhNE
DPgRGaP07BFXJBkAt7AM+G70NdFqe+rSJj7tYoy7nNPkJFWQ9aaRke7U+w7qR24L
8lzWBoE9qjS/rUkGaywSwu2b5sWiNpO4Zv22dhSwxXHplWQFDS5h0Jj29D8fwMsC
T5/FoIKNDXz+N9t7dn9g49dJBoM3+on+1j6Uj7LLSAbIgivOeehglBBIdSvZBMFf
lo8J26P55QUhApoWbt/QjQ9GJk2Ek0fSPA73XcfgM0Zdc2p7icAAQsMqnLxIbetA
MSYvaLHFRky7T2tgrnTiPB4zJaKCT569ZYi7n/xbv+bnOpvhifMhy45oktIlIVtF
Y2G5539ZQNAt11NGPRqFUNePyWoY3CE0tY03UCL6B/00Au8diENTJ1lSi9leJT3M
dq6SaM4nTmBmpRSiDUNpWJm6OhXGSqWtG7SVQG6YhEly4Un6g8EFEQZLEQnIQkSB
NQdGq1q11+uOIAQ/+JXYOZWcVus8Z+iYIIQHq3Yowl+XuKaAF2KDAv9lB4pxT6bd
zZPK+08frOnWx4fs2hGGSjnBACxZN4Y5BaBStwP7wFdWB0mw0bXcOH7mEK7WEg59
StEa6RTHSJSVX1uFW7ZranZwudVE7rLxfacYFDXg5oEIqg+uV24p6QPHQdZZldvO
AP+H/3har1OGX9EG9DnCtOMmL9PgMMUomFZAvBV8n/qgBk0Riwv4cgOPXrLTyBQf
xoWVwa6LJAlUFm/WJJA7SGaN6WJj9vl28U7w0sEE++tuaOkHrEROit+XNAqiimxt
C94CW3WXHfH35y1+5t9nGCOVvrCx3ecAmSevGxMKwjMXkrv4nfdhEwT+DM5TjKBW
03j0kE3j7p0CC8d6EsVbwcWOU4gjcmstvkW1/mQq7HIDpduA2dGGTdMtWxCv0WLE
P1j3kO30uE+w6N/EoxmFQm8ctgKqQNsjE5f/4kTy5Bn7PPV+3+1jZ4iJyyFPtE4s
ca1umc/kDxLJsk6GaCTYnguyzAEaoPJVQ6H7ivmT2szRoVCg+DFWJmG4CPJCJH0C
SzTO/0Lj2f8VgP3Q/illDmquXnu9S/uHkBKrBiZQocFJOqHye/RlL7rMqrwUnVrY
LsItbNicHd7742vXaHh0lQB4NeMqyplbTgh/pS+Xl+TCZVzXKPbEvLTGyekelPli
I3EQvKgmNWaly/tFXGeYMW95hXpGxvtzR7rTde1KN1/ajfwN3gYXikVjTnSahq/6
aLwH1sFMqPQ1cSkjyC4xk19D5HGRW7S0o1Zhv96dVaXF5KdGvzBaaf/9L2e5INWN
8TjMx40NdDb7xOcVZ6Qp+feqh6bs+Ik2G0CVbrLdpbNeIkpzeYjHeKpT9ZshbaED
3tBle/YJBeHQsZdKTv0K/5HtYpQLJr/bBCGqzrrbjNcjJCZFsjQpRpBQW2kppA4C
HIbDbm1pRPz2NplBz8VTcmMXHGuG878Fg59TDGgemVfmz6h7cBn2Cb2HazTmMbzO
RqxJEcFKtMsCHLfvDGSL0yRUVaONIJBoGEfflocTvmnY7lazcpwMlmVMN8VBACkG
KKRV+xA3G99vBHaQMFYA746dQtqBDuK9brPnM6gYd80EyDKeNGaUO0vb1qN+4jx6
N2iIouvAFwdGDWkwTpdlkGBygZQTMwQF/ocP61Ow81L8+AEPOMMCF6LdTtYKfOyw
2NIdbguGrYgnsY/8umaa3ZYf23W1UsES2SCr0CJGSwHBFPAt2ghA8CQmBso18XWJ
AUVdbY3lChPTUFdd6Kl/lkG/0d0wIR8OMg/I7hOu6HxnLdMooetMsBCkoBqPLAFF
B0Sa/A2FzU0EcXVBUVwIFmdEKsxJl3OV4VCRmZE+X4SHfPNftwwareBETFgYV1+0
bdSDV8Bbch7iOJ1QF7bEM8QmJ7vmvxETaFpky4RSJHjHUSKs1SvIDR0eHrx8Ft2v
GdAfcDglulTIz62oZx+sppkkx6Jx9OpMtuedxk6N9SHQ9Qm/8wiOQQhkWn6oNU1q
3uaMbe5kKCY9ACtmMiwSh2i0vmYONVq1awkgWPBALaOjUrYy26SnyhFAR+OQakc9
BDq7qItOyJ9ZVDzwdJbBsUBwPP+avkDqbas5+aC/loteydCDUY//nd/tVbZ5mOD5
K4N6l7WxXP6f2mvv94dDwLgeJ1TT9w+KqqvrKRJ9WbTtUkffQetL2x8ktSsDFz4J
DcunToomzl528v8yLc9kv9o2umhlf+k8zStFg1eb9FnCXH60OnM2bNDvN1cFZaIJ
bicUUzzzUKgBeCYZIKJidJvF9T0fcODO/9hDZnMNdmfaF8vVwGCl4CJo1P4vGunm
PKUu/sFSY5IzjgD/iILr/b8NMABwCsWgOqiVyBsSaInCtT5aGhUIqIKgJ/8lQw9J
Xe9wlEgADr3/Ba9tDk1Pn+oj0rW5TX7beeMDSTZakiZ45lelaALzqR/kBbaZD9e2
1dPLGx5068au8+y6rvpNXm2z2YYR1EtOm7CVEjlQhkM6CkEbkO6JBmqFOANTpbXL
I/g2d+la2VPQcUpZnNemBEaBIlboTCuImrRVqlRBB56X/UwddO6oq6+OxskTjoRB
AHy+xUsrP1Ph0bB8rXgeU5yVNY9KzniVV2k3i90A9eK4+5aUCIILlTgnmw49cLH8
KlmGP8jIxVJmdAMErgdG8qJSoSelwyROcwn7HMZZxEOiKBWYVtDnVqIT3X+Xdc6z
FyR0eWSYTqJrNsFPa6cMWq4Joj4pkmPTi8beN70x/QMQpBgCMnVlv2NirV6CVURA
X94Cl0LyOzjSitIh07oBPmHVA6gcPmaiXxN0uMZ1vQbNnaY92Gn8Roz6FJeTrkmA
lIrMlyWLG1Zdi8Y2PhYST0nJPPiO3ZzA0ELzIP4QyGLYVMndqRlaHecbs6LppH+D
PMl07gZyzK7b/rAhn0CKo/fwx32QwTdQIAIS5SwFDo+W+SiMcEnQTxs3a2ItZoCq
dSJ9EY6pbN8ZfOaDx/QNktt7MtVOnpRpIJy3wcQVJMikeET299Rbim8BmDpo2De+
V3gRSk4guDJi2WBLZNOT03a/wI2gIFOSlUeulSBs4x34qW4gMB0TrigNi73JnE7O
2PHiSWGedVCytAHufO5thasK0iXIoTwK3pOlVou2j5G96oV8HCZKhg0Dc6fWj3r2
P4MQ+In0CIQCyy7kFhqTv2z4ZfESJ/bu+ro1SwfscBIULEdFhFZ+BsjtTPXmrw11
g3XcEE9xMP9ZEQAtVF7HoJhTfa8PiobSfXFMYhTLBrdY5QJZSSv0k7ioIkr0hz1c
7fcwmrYpUEzm/ZukzHbwMchwHdDRJi0MVAtGHrxaW3LnaVKYY8CsKqC7swA6S5WK
gUDlsYP7yZ6eyTFol5KkVlssLt9bzjI0ZhUEDXyB89pN9xzRMLiTUHW7HMSi+e+Q
dRDst7vC0ASkq9Xtm7oI6+qk5UfPI8YNKSiKHW50NvgQVV2L10zn+dVJa55Ira94
mtQWATSN/nztlp/UNHs2EV3nbAzb2rzUXgvt/B7MIrOtKO702c6ylwQwtmqEfqnq
ibrrc41R/Q91T5JPyNCXaX27B7Zo34VP66eRPWjV6/7xUhUinRTq3RSVLQe0emZl
WmdBAJO5iBqlxRmsj8PP7+TwrUORCcqjjYyBSXxWtQ/SYoqViy4fznP0l+n7GUQ+
YuR+i2OC+FG5tTZ4CFuTTd/Nk3eSM05hnM64UYUAti1dzkBPzl62vCsKkMjSHu+B
XMVzQ0IFgf5FB61henYwmTXpoTFb4RStQ4n6o5DeLQEC9ox5zM6GwJwbM+HgVLSk
w4xL+QOHiNiajZfgxUJftJfjiViBapaw8tC8qhPn6KZtiRRmQPfea70+RX+32URg
Xn/KPk3j59slfaBY5h/y7v63w9r4xG0pqoqc3nXSOB4dcpruYrxnfbkTUwPI79gr
ODK/CyasdU6wIaEyWn84ngeEgMz/NY2iA3ggq73em54KN0RgZNwKaN/ZnRItc0Et
FAMSRBmNB2QzUQqHjG+2gnl/7YI8JDcQfhvDtfEO4t20F7m4//WJPdaZED5l0P8y
uqApAHL0AAMnX3y2a/4MO1KBFZx2vgCXm+NfxXt4D5C0+aZbrnADjypBpr3eTvnC
Y8q4XjecqW62tXboFthaInvpYHnSQHjzuwkI7FfTQFQclQMkFX3CMx6YhlTV1Qs6
0oo3eS5CZrTFJ9cEP/+4kzEm+Kwnlyd9sd/AbDwAs0KUBzhfsKEuYbxmXbnq8Q6N
jGBoW0yG8pElbfXq0tcHqxwH6l+bvNZMXJhXFoJlDrX0D2uHELqh8seA5Y52Mfl3
3FfdYcSLp01ua7S/2+ke+ykDvA2caRqXDEsJktZxV2V63BIraNGOyDmKQxM/ijCK
EeYQQcuPOIvmXIDPbI3Hu1evPglnNkJ7XLOSRLJx1Gwx+/8GJtpjBzdyXaEHfyNz
s15AshNCzJGY2hT+z7a8J6BwMxg4+gJXtPLeH4v5h2dSAYzrI3OrvPx1HRhj1Syv
SFKPgc2QcPhpId/NuydtCEcZchtXil6SgA/V3fFbqqjb0+8hR5IKgHB8pjjruk3U
n8e4RVUCcDlpuWooYfLHHM18XyHM3XmS6xlvCd9QlJok8xm3io3zIywhYEAU9qtU
sL8cKP9rTpJwE9iSP42lEuPxLQfZhMntEubs1DFEhhaXfxSOI9lD1isM0yGbpsCB
CGaVRJJ14MdM2s4BrjWL1wHmWvH7ttWw7TQS+fOyZ4Ln2daUnaALY6MvTOIOJQRW
IwdMzjksW3wvkSmbkRTbXn08pjWqZS+PzW5ukSOTyNHrWdRxHN7iuX7y1a+xTzq2
p96Vzm7eiLQrUGwo2xGoZ8T5D2+rRSunaOdpFBQEjAARJy0jeJM524MLCjQb51M7
D0kfBSVwXdMlgneYynGyfE0I0Z3OD7lb63k9SDEXP3qfUl+tKA2P0+tbvZr//SZP
5GS4rktYfqu/eoUjb4B2kX3fFKCxfd5p2PnQpLotnzl/XzydD0v/wKRyUPY3SI1w
8mOS4WGA+vUM6Wf+RywG9jE3fXlxAo2k0xe9OsB2CnOIRg+rsI/5onq2kLT6bDZ2
naaeZL66RLplEAiPKLH6Jxmzr/82bavhiuusllheU1AD+RPXEAxqPywZ94uReSl/
fgSHXrwnauSLp0pdFzleA75m3YIyyTOZZmNygM3Xwe77egW1V7hk9hUE/FpUn3+I
taoX0ilW76jS8vPCVBsDflNo8704pwklfgaAaaubFDZhwjw54gBEhNMY26UtPjq/
3i2CIqoEoIZsLSEZqdzEfIGjnJD8YYg+S7+kbjhXRTJqEoX0xoIgqPuvwFXnYdX4
milpH0hplkEY0G1HeXvhKXIu1W/fnBNBkBKuXwh5qstSVSQMUA61Ya1/YOHHiG4b
JcSUlrb4C0CKsEsUqinBmHpogPSo3ptaUQuSAg49R/6g1pB5DzBJgkyDmUx9X0Rc
PWAXfTgAO6vZfys9+aJJ2vTRiIXIRZlfupg9XlZ2GCSBCD+r078PxQAnHRc8R4bN
BKO6f4QdNtx9Qo3dge8WGdkQfiEz5Al8n1Py3/Ef4TbS9j8e6MQkGNPqrcwNM2kq
GVd2VZqEYopXlSwgKWtC6ZtvvkOo4d8DuBucQsuLE8n+s8p2lWZ70WWwEwh0ejoU
GVTJz2e75k6G2et2KCGQyHQDaCS11Q7RJm75sHwqEOtSsumG7vzWcX7umPjyqTjl
wFOpjy/pthUxSTfciBxMulA4JY3XOk+4M84PnRLj2Bgl0ddGdZIAvKJWrMIzWBdH
qmc4XbHt+XpMj/YZPg/k1SrRk2haxzojogSivIcHp8Q2/gKnAC2vNEY8H04e3GoH
4j0gtepOXFdBNvS78y9cqOYVhkTU+sNUWfO4b3nUtM14RueEbhzRXY41977TFExL
R62flQyJMgu2fu2t8is+O2Rgj4JQITv8Qy9WJAjZ8Qm7BJxTZw1IypDAp7J9czWh
nx838erzdEEK2IZoIN/CXGe3NvDKFJo3MCB2ynfc/6IPp4di752PdqDHHL+pFY2a
hsiGQbaEsVI47xpQcBKSmAuWjQBbPiOAj+8jAjp8Hucx2mjcTHgUV8Fl/CUGYn1m
Cz4l0D3wqwcBbURSPs8qR3UsL4KMlMlwJkC0gBC/JT3FUURZMWVX6QwDjSU3d+Os
5M1ZD3DRVzUEBbXONq3SarzmWI0tOOe4+YTcXeZeZy3CwT+tZQRrExqonKG706eT
4+S54fnU4xzgORgPR37LGpL7O6TIA1hV1Oq5eTGR2nVDAv9YYsu/vrhrvLJVH1EV
qJOEPPArQSDTlYLMkJDTMgb40kNRWwMNB6C5rzKyw2mQLt2LCBtGT8Wb3JPStbJV
4xDX1QuOA/1xypAvtPfbcuOkPwJTOv+xp8zwoRbdZNAwFjWOtYM555Th/QYlhVOR
9hw2U1HZutdiWWtaubzsgokqYS/6ECh63eJQ/O0Wr+rduEUTCq2v8brHijm5Lmqa
vFilZDREMXetjKJDF/6OL9QIJfWafdzyCHfSBBMWtZA0vz4knwYuHndCZktV8X5l
MSgV7wsbi7Mh2UGLgHiRX2rBDiGijgh50QJEjbZvCceodnIBACSEFi2dPQRKj0da
uyKurxUlj+okpDteL5ERWePqyhnNNfffp9cFT6+Eii0hVAwiep1q7jWWmhFlvmGb
YhzoeK3VMHtsvKOZFOiHJHTYvNPfZDKcth1HmYTooKQkRjBZg8aVpspKWAqj1ZGl
xJmmyku4jfBFzHGCi9tf/YDmuBEF9IShUvRBpLQXfuKTNrP/PMtJObN/ss7G0T6M
4jcgcPABPXkO2OOgL2LVGvkwnfuRvg9GTg2tDUbm/66NViUKB33MfbPlBynvwP9E
QRMMYdv5JL1bO0Fis1br7HR3JVGF4q3vfldFYOgbk3vHDcpdeYPnoRWPQKwQ7ezq
QEyqLC5qfxyf2PDWOXM8tZijpAnKUIrY1mnpaDkyO+CpBiGw3t+mWPy/1riaBHs+
SflfOh0D+A2/RSBisfxGw/mcUXHVX7Dqv0JeichcO6MEmCiF6hOZwHUwRzn9fnF9
bWnv9VgXF+iMhNzOLpUasltQf5aL2tc2OP1/kkCmVEz5y/zac5liTK8Snp/uDgk4
eH4IgkZgrqWFWSjAE1nf2fwItEBWXRJQoucRjuzOLql0ki8tN9tOoJ77ZwUvE+oJ
PoI55nTUyKYWerGuPSHGRepmeYC4vNa7rY2oP1t6DtEADapK+8BxCOjzZZXoYrcY
6rJtxKmgO9bOCgInASDQbdxoPcSzW+9Oa6NMzmyYXwu9YZBMmRu1f8ioOCDMXEk4
CoKNV0zJRzSp9rTHsgL1EyhAovReWST3PrTku/DlRox3BK93vLb6WSin7vATeJjC
trdqp/nfpQK24iesFLPp1u0PJUuwMQhbHm+QG/KjbtWMNYIxVwKXB7+8T1LpdW+H
ZCwv6Mbw6d6hWrHenzhiDT7W679Hx2M9cQgS0wT3c9WKA87btoNstP+M1Ks9W5R/
VsErPCsmgG3ywjuoHSemdZ0CI7cpS31JlUvjBFL/JeRt0K4pzRN3rioHVu6zuGX0
0lrwcAyW/LcRC2JPV2m3c0ZoSF3oi0wZh1K4UTDmw5dHu2LB6WWUgDnu1YqGhRS2
O8Ieerhn1KzESNnhMzWhUqtFODhCDNxMmAC4kcq/lwslska5lVFn0Buj7Mr+arA+
hu4s1pdtpvW2YZC4zuKHdYt4pXAcpnCVAuDzOWxU0dHLssOpmpXtzcgMl/fYY+FO
OvWYqMPTtky2TzEMZphqjEEUnzesUkpw2iqKKgo3hxaAuBiV2gLFTtETzPvKXMr3
7JlrjLU2/zFG0V49DP+1FqipKkpDCC8lyAWB+/5I1hP7LCrEVxsv5otreYuFgPY9
310ao1ByGtDpM/8LIkJVR+uVJoUpoMRKYpNBS/k8+2E1gLqvlCT15YqGP9lBQmaw
5WyItMLBfBOzKZD0EvwptgO096YiRufPh74h7DjVy6oz0GZFBCHjDmfqxG/ed3Kb
Q+6QNga9rQWCC3o2Bw03gI4LqZ1wtCKAza13FM6N/BwwEyOX1nn/SusoYXVw6bpt
BFQaDHKVcvhxIy6Fjm5IVImqwoEY1rt5Em6mToXrOHkaqz5EPTcPzG0mRmkQv6s2
B/s+d1tCss4hvQUW36e5RavgvPxrdmtihQLorBbV9QP35fbpO2tmKRZsc7dWVHVu
oQOy0yqJKfXcK5KsZwDVGzjmFJ0sK9yfG6bL5838olk2e46tFfuP1u02/oZwlH6Y
c6h1BkTuvUj8U8SiieS3m1P7jcCrToY9eY4hlhZ9sxObeRg1Ky5096tqoJ4BHgC3
foZor6tOQLNNbp1JMwwFhgbWjn+goNfBRpBxLJF9jQ/iBNfZ3m9+IkSay9xEyauC
hSKLO9Tq2cIwQEHhOZeqZpBL6LPj8x01hunLGIlnDOpJ7cu2QLu4Cvk/gGiZy/Se
tSqWl2VdT2NJrlR5u0wepH+4E2yqeSwxxRYX2KFlQ6KeNn0sDbnMgl2AVf5KDELx
fApGta54VY07vK2LQcRMi1cvhMC+8ter77vakNxbFGV65HvS6onSDuf7G0lxY4h+
e4LCd5Uf4RVakwW6lgcgdUQ2IUQvP87A3hq28UVZByjjnrmwD5YSvxWoABFzMwLA
en28n9c7zVURvNHhnG2XTjknnQiHGi00tBJkG9pdVh9vHcIq0bB7inrUe1yGB3eC
lz+qCx/HVYHzlBQGDz0mHi4P9UGGzGcYY7DBnWA7jDCRNa7bhVroM0FdUQervPXB
+2Ahg4s50YLKSVqGWVM1QeQx49SpBg/+zeCeeeN8PYYw1epbiC4zMWqJ/7SWgzni
BCQ/hnUkNwDuo1JxX+3CNvp2NqpqJrIDKBFGQ2psYC+1xTbzcmpMpfd7O17QPfpf
N11OI9M6ck1eCDy28HEDhnOznoQopT4ob/ZhGP1L8hsNBAFoSRtcTv/NpOFIOYx7
M9feBOg/PB78ifW/kpL238VXVYv6gwcrScNdafC64sER9hjgjTlS9YXwfgDVzDUw
AS2HGthxbGQ2qmmHtXEIEFlOLjJL7Zx5MJHRvRz2v9X+RHt7taeHPHrzMgM0xaQE
/+AEjRtUagIIZOVdSwOYmwb3vYq87kaGlI5dV2Y6ZnvozZhtvfY2dP8ohPG8L+X0
BBX+fK4OlhTLHX4v6rMLw/CXk35qLqvZKPAWM6B+IMH0I73MP4zy4Z1nmbFMX/HN
EJ/mKjDWOtZLWH01l6DpU9BMyh04pDFqIv9zP4stZmoBxC53e5shIn2nQ0kLac7H
+kmu2/8SAEw2C9BKlWcD1YhwuD5TeUmUG+ZwFMwovcUF4Yk0BJlOuy4zzEoZT4KW
9NtPi2pmhRq1pQnWWVPI9IpKKc25oKYblBcU7Ph6nvP8quxpXxOhgwlLFzO+fnP5
q8Jl5dt6hAgaSlujLDxY4EMLWcRclFZme+u8XvdTdU+/37FOH1zswhszQROSFoZw
pV68RZiU/B1oIpMFv8CS6Q//DaDg10IyPIS+XTRh9wqPj1COefywdYvkk2+FGJ72
UZTY+gPFk3FZfx30gYULJL6MI7U0S3+lV3qoC9IFA5AuhxP7CicmYUVIT9ZKjBr0
komyZNykK2UY0wm1BQg/3oEvRszSrvUIdS9SR4Dx6L5CsdzwGwJQxAlwuhgHc9Jp
DVuvabPOHO+ldlcfrjSAd0y2oa2rJMR4R0GEQ3wlepGysx8vw/lkztBLjVfTW8Z6
t73r7HqqM+1OHw67iI57zm+cI2L1uUUl2cUt57g5nZJ0ax9MvaEQbjRUfU1NVN9U
yQL+hNkMpXvxfwmAmleN2eOuXDpObp1Wqv8tZqFBLw5SvRhxRm8iOoC2qxx01nOd
tmnqNWDlKbuZboIRNqgNVECAK3AW/RXUNPtuleOYrr9dHSPFYIRQN8R1ZKAGz6eg
+6hDAZxrlkLWPyMMPyTrnqwqoYmyqRfgZR1yRLdOrKVK9hEmAlxv4i6Nyc3I2Orm
iXt2OyhyyfB5khnTONGMH+VoSxJoBZHLo8LZwo2nm/OsOxsPDq59zaOdl45x3V/c
yA1PrwKxkpRbluunVfkITTTn3p0Sj/jmLd2x+lZJnlgKf97NzMZDdTgDwAGeC/VE
xxKX/XVPoYe5BIJjquUGAxCSiK6UNdGQL5fp/cJQX8VNiN5sNVQdaFwwbf7othhD
rnRomBEg2zfrI8KVxBpDFG9CD/k8AdNpRtyQdDliORHgO5hw6a+Essq2mSJLZynG
Tn3DsUNEcsOQEUJtqUsneI8kjaoTapdHfR0u0L84og/EHqnmORiJ4pbUZIDpB5ZP
2q9QArofWjH+Fw4cmcYMUy7NnFMGMsSUDkHmSBqCOOJrJDJhHNeDJ4VZLmauV/ly
g1Q5/F91LP6fzmW729CGObDayvGQNgiTMdnzWc4ICDIYxRSMI38ievC3+OKUz0rx
h/HtvwUkPn2LfXdI07VnIWQJo99B1ACktLyUqUH7K6KUPvbDj6NbTObeqlTJpQu/
qcj3hYgdYO6sUPpZmpRmgJL+YsTCrkU2BUB21TN/cDeSBt5reJyNaGagv9YpLtEc
1Ici49a5RoW93s1kZXo2663yr/hLOfR9imtLXIz1KJ7QzBPFkYhd4Iu8zCxFNEjl
xT02/bsqTGb7A0IHeBQ1ZP3U5Hi0GsAYHW0fpq3n0bjUNXj9pbt5KmL8GVr1w5BB
ZHaDxRu1klTlsrEBuyOmONNp4oXH8v+9PTnY/Xi4kn8Ur7qhcdnZUq9Cj+umBByE
kcitnTN5ejV7h5ntPP1w5G9NtBspFX+ufJb2+YGjEBNPd01oHCTGD882r7T2/cTJ
JgZRmYUP3btSSLhLBKmcmMZn6zaJ4QKPecpqz9F0bfgacdZ4rhu/sCdUfGLjcmaS
gjgMV1gz+ORsCc9Y9gL/9dczzbuNugAfa9gUtGqHcYe+75Lr+9aXYsKXtTkGdRA+
GInmUqslDc/xXZv4v6QWnrMV6ZhmafUCXgqlYu9sGYQJKNj6HHQOiTlpBiNW1SPy
XlsOCj5Ii0FhpwaAWMQQrsprJp//HoyvvUsCHh9fjwwrX3U8QiIR+8M3yc5JcGvB
WZSDeBFRykJOEmtd/4WOR75zCprPzFFtHUF+KRrbkMuJb/OLs4FJR5nZ0y/Orfjr
nrlArkUn0GlKuWwALVx0BQNtz7Od3qt89cqA/LqosLm+QJqi7Hx3e/i5ATTQYcF6
AF6TvXHBrlWvOPHp+686kW4paVgw5AIW8mG6VKv2tYfXqEPrxqLCT7V7IyRKfjuR
DUQXYMFh0V7vdarU7+i7rVv8yy+rAEsLDzQ3BX7aO+pxhRpsejf+tb676cPfPI4y
4NJyafPDjccaFzX5zKD3wPASOQvhO71YXDIAePmzkVDiamFRn4tAbarvE+UAXNaf
98PZI3unnDKi6uKtldOgsqC+QyZv13EtkRFVnd8vSE8nmUSwtfn1mjqFQQD0Mwma
d8sDgV5ARKaFvX9JQltoVk1jUUR45ZMxgT9wsQgqXGVLBG6Ty8Ffljlzo9GPh9gK
KpSJ4keBcFnMDliZkgMs7qlC62Oij+3yfDiUY4qenuk4CQ0/Wf8GI94iHqdk8xSb
TdHAQT84VMG971N7+IWGabKGgl+FMyeF26l60mdPOTFzaEd4QkT/sSWAdHov5fWh
8mj8CU4lbuzfwRobPsshb5IBMVyTG3STHzg4oejyXe69Vl0CA4CWWlkCsLEYcauV
HzHNx0EuYrCABSVTY7vh8SCaUQTyS6L4g8ROup+B8wQBTbMU/rG/KjfaTBNxfYwt
Bk/3XpggdkVjonE7VMEzq9TIw5yi6bBX9+VfZIhg23gTrHhG54uCMHi9ZlU0uR9F
pgy9zzaqegDoEuGYXk/jzbMTHeDO8ZnbkBoBvawj4JhcIy6XVyM8z4fiu7LuJLT0
y1NaprGz6RNaZIook3thoRsLhq5KrVeMC3uVbVEUc+kilY2LbcaWzEIp4aniPGN8
tAVIVqU/QhVUqK+nwz5lzLjF/wntrM9IvBMYbm8xdJpAb23hpDHUDmmv7EkoepGB
EATBNUEpA0WwQy1NQemARmnY6VUoRkyq+XKTy+3iH+zyZAFLht+HNo5PfXsbErnE
yKp3mUY+7D5CD2rYt2zZhlfdMkOhOK5n6re1q0SvNd+9w6Rj6e3mh55guWgejIE2
fRwddmALw1gM7ELq6P+nVf9B8u1193P1ciwlJR0Y9Af6Xcnxb7/W3tt8OS8FsWiQ
a3Us7jtjRQ/ZGN3lZmT4iCJNgXL4heqR280+6QcXni9+B3j6AuHF6u9GwS11HYom
kG9wGBVbzpW7SpRm+Zc69IyjeDxmkl/g5xniqK6NyWrPvaxNE0m4hieyGPlRQ7xl
I6cp1cJ/Y5z23tl4JfVjLfAibaufqGetnZamIYeIW4hGUkW5GP7t8BqcSaIxWM0B
j8ZIuU0hfO5xXg9FijMejnUTkGEoiqPHlW3gqMyBQTzs14TZkCzqgLVRgqhw6xp1
WlSUnN4hDADeQdPQ4GJMzMkFdrjUeeaqooUBkqwg1j+kgS2U3pQ49X14zmFkQgbY
D2ecKScWRp0y9YpytD1PHnrTNKSZCP0tirY9ow5TuJr6Iay8YJ7nxhJ+Fh1xo5P2
9+DtNgC6MQzWmlzs1h5FQhuGIyDtIHy20d89LkKKmFMd2zfs2r7VQNyrlNJ9sIz9
moYw4BaZE1khPLg8e8wRyolfdsX4+K9KNeHziicomoHFh0wEvEoDvnhlPJ7qmGNp
7t9orskg3YptfO9P7yk5/sRBs1z8sM3dptNK0u2W05WDKJ3mtk0LFBu4CYdzT4oz
2xeelU6FW6imJ4Hr5OEJI503QgNXujTNKK8uplAgFeYtoS/KZuxKy9ZZdMlipBfA
mnXJ9/9q8U9qUK10aDPGc4t8eYPlzys/kc4UKnPJuO+5/REgt1O6zoc4F5+slwR4
opqQuG7J8z/ny/+Ip7KCUUeXEdToGuXwkcjjQ4Y9zTVxTND0nPzq1EJQWSLZRtXO
92iFB8gdXrLde3SSqIBapVwuzQkaBI/7YD0wNPoR06HjD9SYT5UtHm+DZKsmkjD8
o/DLzR2Wd7SLq9TJLR7PTnHaEIFjVmBkcHmAvlApLSgeUa6aKyAS/eu16Q3icVee
4BfGToDndXhMjN4ANgZt9gQjNlFKYFC4nzCDXE8sSIlZy4fsRa/IqszxELZMgbA3
MxqmR+z70Fowy8YSSJQx1dMIc+HZgcCuF7d5CncBAFmYrSPUUQnF/37RnVf7xOAS
zj59AKpoDHgENLpYOZkCCkXq2Sfq+3MH0ztPAHj7X+6z4YzDBiJB1z6mkzc3n7lT
dpWTw/5VEaMzQGdErNTvx/oG06FAmomDipeod4ymx869KRbHSWgeUJ0EgDrMxG4Y
WvTcM0VZVhUJRzZs2nxwn0omnjXAUkmgMG/qtrjzRwdC2vXO1gFoj6H88dpAZieR
LdnufTtp0OaxtaizMpYV59eZ1xnschO7+yH9hS43REQS5trtnSWYm4tbsjazm9NX
usRWgcdSXF+UkQQKN87zE1t15TqtA3/yN5zIPOZHOHh7R61zwWFd+LlsxMhix/XN
xBNRdTN+e6SBS4Rue8wxwWEOPEfKAA6C2iny1vD7TwyAE5dTYVJNBWB55Fcljfph
j9UPGJFzMEiJ/pAMSA5iYYGobulyFg3VLJPnMUpZBoeXbDZSwsKSnmWFFPPS9zcq
bi2e0EtpkTXriop/u8Wf3sjN62B4GxcwIKi+aPbjbu/7A9ZRY8c9uPYHvP46u83f
DVy/L9IGqM926J+tLoVx9AxTos8xJG+6swJpbNGvH9cLLDgdZPyhsYc0bnB4oeYH
plXi5c9+AOmfAq5dvtCWIm/KEOmljeLxx13Pk217ZuFavVEaD0J0e/evzHnt3vsA
/BIzHZ24eF5iUFXWtj7jeuJOrK3/CkStc/pc94PkJVRYmPEyTjQixCPRvRpfKG7T
l0MWxwHKT/qk3gSENRZDJQTmnWxhjhTEHukTBa/s+o1BPjFHJ3QW0Y4P9y8uxlNB
VrFxkfeHl3WiH/UHPf9oz6SaXSQ0H2BPxovlMcFe4vtxZUGjwIHqrjmfWpjIlp0d
TrP08YzY53O0doQxGUtCJsjR9PoRrGM46T+RgIg5liAm63JmasbFoILxHuwW25Ze
BtBieGcQS/MC0jhXHdgDSKGVWqJiuFE07AUZc7zBCZwuramGR5DuzrcI+89CNfnv
xc8nHOSG47zVG7bbq6rN56qZoMnTvmC6RIHCK98n7M0j2mcpC708b9KC3m8/lt60
0VdHwKdDm5i2B++HfKBNNYxlF7ZcyPrR4ex5Cn6hcaI8/cOxS+iob1wya50CUtpA
y+mEuQoJx7ybbwjht5mWTliI189+TnDolfbgBTmUWHh4wman/DcYGkrmgChrKi88
WkpDdIjaRmC14MLAqpGWn9QF+3bSgW8aWCG4aQFJPWNqW4emQ+73RlEP2OIkXkDp
UqnDSQdfZhEBhXGSbB9tEsBiUnj4RR7uPbFoaGhlteMql6qQAfCfIXWtTz/fjT3t
IqcgcQp9PoFIkNWQx3BeAcpZP7MOAVqjmcvfFctepPlRzcB6SBYrdGVtL15rIa9A
3XB3WFpgv/FFViFC1EPWcLjKw4l54zuW0CAdDtt1hN4ZwTfxAM9YIYxEMFlotbxh
zpBAHWG794IpN/ELzdbLTo6mOege5Hjk/m8CLdAIP6T9EXrgZ1rJ5gEINKSRTldU
GrP8bPuGdEH0/IbMW8+lkLh30E3jKnpAT6gsK955j2DdW5r/N/wG6aZIYwXRnGUC
/fuakWftPvfJr7owzIAGaJ1KebcP9S6+btgYeyb3/49hqt/7YDP7VEvEXsgiRkxR
V9Q7PbAAfeFf9uyB2Nd/f1XerCvELVWJZIQll3Kaa1B3vD3fJN3Nyj91KEdJjGgP
74TyvAehOrXW+HT4FHhQIiIwD9tjoMdi0rSYYmuQRRYBVJhaizZPQOf7FF7fn2BW
lLmx5X131Nxf1+IZYGAoXmOh1oSm+UfgxtoQWJVR5aVuOMhEE0ic4SAW6yC72R03
k3U8nUnnVA/niT92vvxkzAqwivRY9TzzZaTA6T/kRR9FSXjpFioCXwjDLb9RulyB
EqTNHWE95RsqM/KE4nT01sNP2XryaScA+xUUnx/RgCZc9WbGGV0qXx4kwrY9aoPg
puXE2EeIhKnouJvAt6YrYgc8W2gU/kzfBgl9QZljuGaWX6dEcQdE8pVfAqfwY9Zm
sr7tCyM99GYSD+19wbmVQ/+9GqKXVm24j18823Y4PftDHHLnXVezsx31CSTRuJ4D
dY1sYZSAFIsvu+tGFt3Q3WLFQ+yrHYMFnledRiPMQOQGrHka9aYVtsVxTdGOuq9W
7uvzqin1ZyspuUb7pzfp29UZbmCeZ0ZwZzTEZ3dlgB64ipZrKvu+JOm6wgV+v2Y3
i6WZjvQFll6TX3I8U/qLI1AlWw4EFrYcurq5FdYSD62VGif6ck/GmhjufpL5gZev
cZRfnuWoyU3zTrxhLYcUyYWmdGKN4Xox5dCpHasQ75QJf3YmHsb5f2/nMDnUaA4S
XT5Y0E+JeqPl0DTdW+Y5ybD+Po0UlNSE3OI43eCY4alCTHKyuTIb45GdFPAQpuQD
+lpVXRxGTUkxWcJeD2hxk45VzZ9Ch3VekCN/nHDT8e0H7byCXTfjpqQSj0PEnOnI
MgYEw5a6yE+YxV3OsA7D/Ysn2wx1s8r+QkvC86od7tRU7sUKPdmsETXEPOZ26HqB
OKub/c9AzJaUps6Z3mlhOMW6Qrqz+nTbfhml/Dg+FQHrxWoflI7on91c2+rZNdrT
28uwxdoiYrq01C4pLvgx3RxwWWO1+ku+RzW69HEFN4ySd6unum9IJoyyR+qR89hW
A0eQ6sy+7sWJKDKoPnC1wmbD2cBPT7unN9myazzbJMt/yKAsROSiK+QSN3diT0iO
dk0YF13JFqfK9w0Jv8SfjQgKjIUFmEkSp32IhFlRBNk8kRyrIWaTrem348kMWoz8
6vQt18FdI+zhLhGIiL5fuWzdUq54o4w5tSf0QMPb1JCGhpXeUMtBjNvo5qF5xLUO
cXbWSLkG/3uDX6zwuzO/ZLl962jeZuZEKz6z2sfDZHuGdpmGW7RqMnQoiBib2ykn
KJeO4OyQQ9Rq2I5KpPVBo23415Pd5u48aBjsCx1KnvWnPYcswWgCA5fz8Sa6CeCc
tEz4iagnyr6waHCgq0bnTyHz9Cl8VmZwNtUnbXNrUSc95fbvrweY5367f4ddwx4H
oaLIk960waLPNq1VQwmmKaZBgEqPTAFJTjGdTOfhgw/aZy4PYsR+kXXSeFueAmeL
XyXiLN51Q0SnehCliZ4WvF1eO8xJ6TR2I7mo/MX5wS95Wpp2CLENZJahJ1X6yQ9U
VvTBNHwrbabZ3gZ/acnO4iAVaUP/4m8wS9DfDCtfeoVGE0DUX4bisU/gQY2dPayx
nr8KmFXCNVgUOLeE25fwN51LWWIULl/YYRiYE6tHP41UzDNQxztT3FUfgGCdQa1r
lSnB3UHtmhDNRH8t9y5kYIB4BSDBr9A74KQpsHfYQe3ZhUeVRCQ/FQJKK+30pZa2
RMVC+mc4XjqIVM6Owz1dLKQJiS0Fa5W4zoS0Sp0PQEsUVY7OfZwhpyCJh61wxBcR
mJLmOwm8j/1lqbjqPjUsOFLD4kFuPOki5W0BwdJT9Fr+9A4X9Pt9BeogZO2IVLBZ
hHDsR2NS+choyiShOka3cIS6eAaENTyCAwlutfxp0Cmbc1MpvkrQMzZUhpo8Oo3h
eTuBxQpub8uzvY6YZc7XLaugGDlJh4ml469a7q9cjDQpxwFfCPQqt9gVOKZKtGAC
CIdVlPuCgzDK/VWr300lIsxdWnIJJuWIK0bvRWBfzF8DzQKnL69MlAkZ1hWa1k+4
xqmQJtaKXYoGpu+BPEhuyF38KV58Ckuxw4eDP7SxpyXruG6GQ4KvLp7VxaW+bhoY
lh9hotv7zjaQ8i0fMl22exg7eVkgV9stWWl/Q4o4QcoJjFPUsabN75PGolvKNgaZ
Ce3wuYCK30za7LbgnVEAqX1JpdYh3KSW5NDjrHY+6OXwHraOsGHNXvTzikdZ0Vbt
aoBZfaWiOgp0Kv8Hkz+mRlrsLVbOG5vqioBOyQxpP/Pl2K8uqcaFmUCCJzTAoqj4
8UJqWW9eEECSuEBiX6rngciI0pzuqTbcVYAxmC98/LVgR3M8Miy1bG2JNm+GFoEs
3iZ5HgBXRx/a5DZom02gwHqb1mJ0tCB86TPY+jBJvxKrlNFz/nGDlen8uI4Mqas/
zcoEghV9QkO41NJJko/VmGIwtZrPQUML/eo65gigQmIBnuG1rIFkdn8WaT37XBuP
HO/HU34J+/i6BtkCb53BHhQoQdqCRO/dsWIcR5zz8zGXa6BUBrbYpK/vQPMwpzSX
8s0EDIpBgzMtGaN5bd3vi+73auYhfgRAhjOrAgnFf7O9O/Nxk1f9Zz/oMknJ0hiS
D3Pl3PrPvHJ3DNDHANo+z8sw/n2nR4bAw7xz1dUIosko1KOvQXIjiU5zYB68gkj/
N+gqXKa6OeM1EFxG0a8Vit/p75XBK1O/Au9YSG05SZOACWtKZPcBb/pejGwv+uj2
lMJInyJmn7cxoh+RolzJybrPvjQ7ZfwU5wvxgGq2kBsLt8LM1zExD/099FrYYP3A
DK5tGYnN6evA1dya1d0ROxRyr7d2DJ1SvAfflJhB1CGBhtImC7XazkmNHDxdZvOW
S9B7ZArkQECcvDpqKXRxFvSdy0k+0Chk4sHykyRhfw6WPp8DG5kZMMF7ORcAwKKU
VptAv96Oi6KmBaavNG1ic4SRNgpAF1LEfQeMVSrcggo1JxBt4PIcLQIghtqhJPWJ
GDUyXeMbrZnTu/kywh9OqOeovtSx1vuIFBn/9pl1NEtq23xSiO4h8xANoILYwZlw
luGwdey/4og+MoDbxSjTkmbbTmhadOSXHSmn5ovyTIhZq9KzfcUmYyWSzOsMQBd9
xZrEYrkOhlrfX5IrQjq4Dj72Y6VHMcIqSDyElzH6gqCLHuKx1OOXi4sgpGHCJqij
kERkm4Z6ru2dVW2HWdlQ/H8fRQUzhNUC2Rs/f3xE/XfkWH4MmvvXceR0Q65qnf67
2i3tray4heagpH0trVimsgPKxLaMflW4zovPmIQCNDQJs0T6qR6CeLgk/00WmwId
VWFto+mgkbJ5vSuI5ZhnNe20FZPyvnchQD1G/E/gBCHUEo5aCEchgP+bkmQIYHoY
PoZKUbS6Yl/8KBz9srGy+t7+rXycFn8i/WkRmZY4+2s4lRralKM/ziA1iDAsksB0
t5MFqLGNzaDJaNNLLkGYw1bEHVkMriptsjrA843HFm2+W9PW7QCDR+mlRF85hSPO
tFrBhrnbHQd6khJngnAhN5eOocYRtGTEYBAcSwvKoZUxZWpBsEU6HeQbtsxxMp97
D/wIPR6KKSctunXvyXwnlwWPlhc01ssUVHu0QHMjRo7MeDfmwELGC7jUNFgmEs5H
LDxcqJXeW9coXMEF68Rizk0JKBp09Py698z5WV95b+0PfzG3vKGu2d3AWwJjtyvI
oDsdqHzZ5bRRW7HfEVPbGpR4NW5Cuej0A8ExVJK7e4fa4RoTq5Yop5j1hXH8nhOG
V6xGequ/ye3LBa2ssV+Ne/ZV4GEGRtyB3Hrk52AwP1PSPwQXm8KK0FuGKGT/DJVc
7Dhq9JldqZJ/PiBPYZhl0ADPeFydnZA0vu2gk4PSXoKwt32xb1QUr+7hXa4Up2/O
g78FgA9/Qn2ce4XkFr4I9cMg7eDz051rTIq6+jUVw8JJjxxbAwKYVYmu/d/IWU0C
jDDmz2mn4Dd+qGyhxVS5bBOMHIYBbOnQij8y99ICIveTbfJBM5WI7NQ2rdn8tTsg
FIPq63bsj7ma7amfnRMckC0bLI5sm1HbOLMJ8BHBjt9XMIZrfDZqoLT5sQs9g7mD
UDk8x2uj0JZxyDwVq42239+XvM37SZiaP7rKjvSI+kwFcB07ug8u1E18gik79Of4
a0qsKPJ2+wCRl4YNc8fgR7rsRFyx4iiq0AwQsc4Y5hLuqkgqvkKiLZqpKfwztegC
FGoKUQCtBcunRHg5MRKqwlZUrA+z7oS9cTq55OKoG3YvsInB6AUq2opK5WKIYsZo
YpYWFHGfszAL0HZlRqCBiF5astta1L6l9o+zie64q86VWMN5w8y67lMJxKKi5KhC
EGDyoeR4+JDT7XzgbmLySUJGPljcx1bfXdWw4naA6+A2STLvbhFtOI9Evuh8nQiL
j4Kze8Os2f+jABsroNRaDO9M4PsV2P3O+0gNPeBsLd8stntw1iNRZKnbjODtp3Fp
wxtd/sqndPIwjwfhvNNYKDHMu1utopit9ySa7MD4SvrvFU/jyFLI4oSKMP8MlxMi
28g6NAgTqMVRgjY5/FlXQQa4cJghkx73UU7E87j9hVWyiTTT60OAEZRjw778TGO9
ll3VuR4mAFAzX5Bu37WruQQDg1MvjP47L0aE+bytejDzxVAYp3QE5IVXOsdlX7Fl
5KfI2VRXZU1u/EAnf65ttgEisfXhc3+OKSF1VWRLprHX1NW2e9UpQniGg25IplM4
+ryYX1WdeydK2WaxdtyFuUuz/bqZuQPmfkvw5LuxJiTGQtl+PuoSP1hRjLIB0/w3
pkMkVpzumAaqajTKkfQqFNCtH1y5xurZ6ARnW0iY9Gb9qlcEzDeOt1FpF6XRFDd7
FMYdy0bz+i2Hk5ll0l1mQ0yHNC8yzAY5MsROJ9Q2QPmmv2GyuOick47aq56jMJne
a0E/eLNNw+NP5avztYOq8GvI2VKZjb0/azx7ZXoBpF8hbIXzBW/0yzBFvipkK8JH
0xVuBLmMYsb1EbjrfTEDsgYQtnzQkts3k/w+DTbVgwQTXto9sK08cFBFtvXqdkzp
/G/noR4u1qjo+5BRRLlVhdZY1REkfBJGHhNd49dQQVzXjkKCAa5AV+KSq6dwTsOo
Tcm9fiHCXRO9wcDH63jhXfG0mai1gmkwP0wNZr0BML2i+Qbg2cdnmUVHZjtGDE8E
mzWfAYRF5XRrr6+G2akn+F+6/2ZajB8jXC/bR9hsLM30b+UWAcbcKu7XeImnMFM7
ki+3u9D0r1zB5MbvC+9sY5M4/mI/qxRKNRwUH0Gu82Frx/d+ueTDGaOmAqZUpfOt
eCExlVauSaH9GFRcstt3T+TL04TWiDMyU2vUhFRKS0E22sR0O4TdDVX11Mkp/kUw
JS+ar3DLwCGXsiOjVAfJGb571JfHygUe2rPalYkYwQB+/M24v8eqQswU/ctpfKsu
TyKANfoBjy9XPzwZkHciY+0HTdkzfz45mFmkrUVLIPUWn9XB8lUYWx9IkkbJMxD9
KScFJHdC+GR3vzCze8ChruHhZcLUD0tYf7MlEZ90ONh0Pju0BoMf0ENv8nhIDgG+
Gvz+B3XYOf15lbvtrtFUrGygJMwzw0c+3uw9C4pW3iGFvI5pJMAKjw3piKPaX7P0
Ql5HLUtTV4LMR8qY8HA36xXbKIbfcAa/2F6y5l2ibfTV3SpqEUy2QWmAJ+yg7YZy
yAyJ6LBvsVit4j3OLl+WYbaoZs4kgfeI5O3ETZj2N8U5cFOzukPurUAeGIDTvJCW
pxYk1iV0DELtGGY3woE4f2QJaVKnSgT3Lcc/8HPSIIWo6xcz1P+nRZWXUDaad3kY
b+x60frCVJGgXS517MyPGUho0bceCyIyL9qPpxNOk3M4Efq8uN2bx/HSZ6T0r+62
8YWUig9Pj09uH1/8hn3VWeUSZDd5N4O68XochPPQIMtlC68rGGedjE5J91B5salz
nRAa3XLuZvP4GoHEZD1n7glqt3bxOz1odcmJFk14YXq/z/EtMPB7U0P4F4dJPdDk
vLJ7+bwTtT03rshMaeroOFnALJWVu5H0Hk8EBP3rfd8B+4g0UTg/pVV7pmzfDy+L
b2rGAX2bu99WsumdXerQNM4BhmT6cwUJCt18ojqBJMKzeMzIG1DSbV4NzuqTpk7M
d9IbfPTJv22gU6qDzrX+2Z7Y1w9jUfWV8h9beCSLF51MDwSECmzwuZ6cSQFKAfCI
8bLkhaUaHyUxeIYWqZDQBQtevsB9x3cxTH28kV+TneWSpNWiuXfRCmlJCZ2Y6Ld1
IL5tkgvyVsC/2v+eoG3VU73z6c2PWh5H4v9km4lLOr3MZRme7wCi6Ziz1ULtYoay
dEKvV6wo3B6V+e0F4XzEmS4SN66CtkmTCnfq1OpZ9CPFXyD0M28emh4CL/aSPlpT
jiO3m0N1SMAeMgEeGrGP7zwKSextogs2IUirLZrQj9Z6nqNalShiWV1l3X2gA19D
gg4+NmRCnCVZquCTK8MsSk9j3nLepLAgrU0CiSNeis+dbVLGfs9tWwo/NEzJQIKM
Uu2FphPzlb9pYkQ93CXISKRua5rUUF68HltsScq3h+k1rB+0CNIP+wdLjv+dMW+R
jalRnkPUlEJ+OAjHj8kGvvNJYbBlgAtXfqf/+h5X3CotE3qE4YByvIS9LLLgfPJe
47Edu/Qq+cIE3sf3xI5PUU29e5WZMNeDkMvOOqmm2bMDLbM8xDJorG6f1bEeRt6h
kRI0uS66t6Wqhyrv0Ddca+X3+Ls3cBQbHq/PgPtYgwsun91030VWx6r5gvuletR8
IvedJcXO+FHODMXHouau/GnPsIYQtTuv6KDgi6mLvhSvBp3OW5TAiGkQsVKcztET
m92DYBdPf2RA5boBAHK6mhAFcCuT9vwOR+XK7eT4mepjhgUmev0u3RGVbtyksVGL
8Av9VUX5BV1DssiSaUv9JZqL6o0Q/Nykr6NzDX7Xhvb2/cDFc1YeKTsa6gkuo+kN
NloFiS0PSRK2dc1qSV3fddak5oAmj74nLCAroxwSJFa0+i1PmCvlPdOeXYBi7Cyp
gXG8OuoBSxmSVGjeaAvzQatfuNiQPq2XDcKJ1zFR8K0n81Qce5OE+54lStKACOnC
LXJ63Dvbk9XzC5D1o0aY0fJiQBP5ELG+Fn7Mnd/58NG9cWMFhgiDRdc7CBKFS9jc
/Tw0hl/e2dkxMBOEvWnuCxSURRUlc4R82lGnz4fTiPwxdnCRS1ENSeGChf/SoZqo
IhqMqzD4nMNrwKC+WeSnlZkxmGLcKsRDmIn3giN6BgmS38GsZNOcRmmRpw4xCzol
zfS4vCUy8Yhnl52TtPiWd+rzdsr0c72E15Q5o4Z8oATkskXXEt2PO91zWtvgh4ri
nA6Vq3eBjbU3DZBh72FXB09QcEJiJO8wLcodI/rYm29jLKw8v6tPgMqa17X2ZXr9
LdxCn7onnguV/JGM62BsfbRX4lla61kzwwBOzUiH0GppR3LE1+jtl2x9S8or+x/i
On0K8REwGdBtgqsqw4ihD/qxzOYj8pZrE+lE2GioGMTQLPtCLD1ORppcsTuc6wwV
8QgNX4br1KtoOhCmpioTvmMnQr9UaxQEPm7Of94toUzFMgZf1zJVc9Mi+wBLYOMo
WkPd861a/wTC8hLDxwifn3JRkEMOtuRWeGmx5GdsPmRj3tf9KHNhFofKU/5Oom57
qxiaZ8WCFfg3wtcye8wc40qr/E/Nt2cOeo1ExwND0k/fQni5FC0BHganivhELG1S
DTKrYTuzUxOCyr/lkPUjwIO3+TqVXNl7dlpuR/c2fCszzeKF1kVV1o62NukyHYtP
TE0eqN56a2GpDYe0SlAEaabYYb3HwcTY/NqgrXUcKCmmRssbBWR68eafDzJ+NKBT
xLkUDD922bJKDaBjMD8RpxnxQDG+PAy3DO6dngUEPhYWjjZbJr5g6/rmrdJweLxW
It3ctoVYXy4jU1diHBP6uY8R539UR0fkJnawYrkXk2IHm3jUPKFCSkpQuItKdHbE
WiU26MniQ5KVkLCl3DRBCv+9dyqdn41bKQgnmUFY2rODfaeL67C1l8BKqMZvbiFJ
JApwpiE137J8erMCEgeaJjGdJRY17CMZFZmuGjPqUtZiFtZFAWBtX8jepCRsH1Dv
iWLcIIDjp++LvM5KJRRF2w9qRsYUymRFWujbMZY8N/IKm9idugi5rIv4OeRrpQFS
4tefCX/1x5txGHtr0wtGiWzcEJuzHsz1hDmDy4IhvtXIM5W+Xf4/O08+QWYm8ACr
0e3CU0kiUN9hJTbL0ACrBoWlmmMlCGMNWqpRU4Ls9CO/6ZlNIAZNiSJmwdNs+krC
PB3ZzPQgci6JaRcyY/7lqj3AsdsodMpZG1S4Kw76pT4J3hVxLrNRPmwynWcYLX0p
dN6we1Q9R9Kg2CpQKMG+PfKNQ2viAenIOJYJxQa0zB4CIh9dTxeLEfpaLAKe50LP
d6BI34gykZliX4mrKOJLrcgBFRkO06dpDMZ5tbMVNESxWCOhja+EK75TyMgfbcHd
gjoUONf6BVjZy0lO+UrPJNABryx0Drhe9wnIYIfCQer7lV7YZuK9oZFMfCXwfw46
/sjEGZTEPuYnjey9og5KGDPwVz+VwE6hXzc0FxQtUs8hCSGVrkrAowOlttCKy5c3
0T52rdxAm5IIEj5QHwHtPgwcWyugbSp8+gulx9TpdaJNf0J/dwOP1r5T6h6NH1gD
c3O4xlxwCUAT6hCdlwi4dCCFj4MhL1BN/+j1UWSLYmtdeOc/BgSGhZ/DRRONhtZb
XW87C9KghfMGmF96zNZLVLojyBc0rbTdq97OP7d0vv9AXp/khSdmzujlcb9UpLe6
LBWEJXLSFMYUxWJCaDYtuChn5win0ZkpFKw5ekSq0Jd7gioXBjG4rr24oGCIadHx
lYhbVASc3pTpyM2LOdo8g2qPuGE7Sj8eGmjNZEadBlLTV9c+CnrGUpuj05ussza1
q3OVlaBhi42OtLyaS69a5us/o6J0F1hq3/jULixBIJrSkDgE8IWXj5p4fCYauASc
ksQMvNIedCvVV/qGgLrm4al8E5KJJxGGHalfsMu9gJkP4jbmAG49pM/9XgbPg3G1
VZFf+SzTM7ojNtGXtIoZb+4K2NyVwkQP3RfWHIUguQK/prLRE+vk1xhtfhhLGPpC
+rRn57t3h9+iROaVKlw2bzTVi19KNxOrdDJeKjEEuzHDXyd4xbclJGLqeaN04gKq
Z2FGVVGaHYy4QvmlSxIO//1/2FiIDR3aGLmYE0DBvjdC27hn375pRccv6Cs6QpfW
g7Soky+ToMQ/fjWnDpi0vwr/tOI9wdMMtBNAbQFoejGsRkw1YQhyaeXptUHkPiL1
lZbDJUndqadpkRMM4i2RTJ/qmI63H5Y0VYhwKgZRvUZu7j/er3e84O5VC0/prfhx
NpOQv5yV1e4AadZq19JQipHiR0RQUp82MirMCF2PG4Thvd2E9WTqW9bshJOzuwJu
aNyHRgqCDAlaF9Wy1F+k8fZQ2HtrHPqK8AlVy4fgSyHChYGJZW0318c0kKasNhp/
fEpTV57WVIr2FNwwowunlxGqLnlzKA8b4c2OUI++SJWK8payezYSmdxKIXiKr1W7
IdWJsF1EobXdUH9Aagq8FPgB8cKa+GAxCNDwOj6Gt95fNHEwyk3BdVU+lQ3D2qEj
0X2nx+mS5qmCFPXFHZV7ziKTC+v6jiuBpCFvj4xYf6XZnEGqZr6Gd/CObjaAPL/Q
I3bFXpIyda+uGG5UJvM7WqaYHRDZf+mnul9uaHmOeWea2lfXyaifzPOhikwUQ9Yp
YtrT+eGCAhjIrYJgHNw3Kf7NdE98eL7DeVn8tqDqd6KJuIXWE/U54/w47/2YbHQW
AlE6kmwVwCdgBQeqyGnsqlYhAzQQ6blDqfxhGDFPczsGdYXXyM2Kb4o9ZlV0R+Qg
0FYLIz+u4zPqshtqGEf8XGjOUTSmwOvaolkds7b9nz73nwLk3NfvaBFB39zyHFWQ
jOjg1loEwJTWwN5ikKWv+k4ctzN0P3vHo7z36fefnVbZqwWC+QWCLOfmZzfM7dh0
kNCHXbUw3tL3+FiRax51sO4XwBO/cyuPj83bboeTw5AWL16H8Wn6VWx7kMbn9r1k
xIVvdeOMfvQG91bXpOgSb8yQiIYSQjDh1CKi0xcdANUeWz85+QKmDuBw2gchvhpU
9ZSGQ5muzekHrxTND/QQnWKqgenKm34BiMNRKuuzK3bdKIUluz2eVxk7DqNcqAN7
cYSZ9oAZ7hLxhy7hM5GOQo6BcnVXOa8VJiTslOcN+E9aP8k7Tut6iTKNQwu+Sstt
3jAxUVfD4dbyJPoZK2UbHlzjjEtvUjiwhDquM//pTNK/7wDjqi0kUQOgulpjRRTf
1TbPTQZEHlJqTvyIrhF0cTymL+JoANffncTiVAFmmCvajESwaT+S5PPh30DIzlGl
ZBhOGsTA60zG0E07xxm7n9VXfc/tuzeKaJGyKBftI+2QSA07CmtfdfxxMjmrxvfp
G3oqzFvzWnUkqRufVbanNf0UfgXLSOWuC/Pi1y0n2/io4wOG7HK7voRgOGYh3K8F
1nWHev+NgAHKnLaXh+XMc0tDaUlShXF+WskUHYCCOItEi3ocO5tU8WIv4TzgjZLm
YcPnVZ2ACwwB+X6mVJ0EyB3yAtZlwaVRsspfrePqSIuwRwskABaUclSt5JH/nGCk
OpdprtgplVmh7RqIljSbHwEU5YV+Yc0wS616hSTnunOCpLWoNU10MtMMlVlzLjrM
9dCCWiG/wsDYkfBT5im5CksqdN7mUPkSeL5hXVgObf+NIcB9x42Xp5VxL5AemPh7
b0lBvH49OU1mnGKScRvEtkNZrbysLw9DhUx1Qv15PW7XGGLPrXUV5Xcv7lypC/UO
Psor3R33t7aAmVq3bWUb0n7bnTw7hUE9yU0QWzK3azqQWk6I+/LJXeVNeBPQCmAa
x/2uR/AAidkmi2vXvHcJc+eMAfbihCH8Ks7qjmPRoi23Jr7YN5tbruGc0oF7qFT8
qd00oRD13/ho/luCX4itDM/heLVbsLKoHz6Sw1LNfDr5rj0kXCJNbVwMr6q2aOfM
yoJTR4BmWJzUE1/6q1BiBqbxPZVMCu77YuxNOWP4zziSpEFsfOQfXi5Orw9SGj8u
Ltjr97imO4i2LS8A1QWPVjoW5VerfnA/9B8r9+SQzUp4fGcYvgfkpDhbiyz0kHcN
oTA9omg+Ypbdu6WxfEw/bSxG3RFjYku/yHYqHchwwNb/gWbUfK/rePW3CG4FKeWB
ULX3Pq4z19We1/p9AXRTFBACea4Bo2ELpT90Q+sPIZu0DUfpUHXbmCgvm1SKCYgf
4nQg5PaD6CJJ4EDGPhTjlQeqxaSf9svKydDIFhkFZ1eo7xGmGHXkUrnpeRsIG3iy
lofSvDN+VwKmATDKGitnRx4J/nXEghMO2OXx8KWQ0Pt4XkutR1CzdSII2yYk5hqj
gZ2YlEIKgoyNv4E4E6lEjU1rNspLZbuemzOzEVnO7SpHMzzRaOcNdYh8umHIoQNv
4EGRRu9nwERCMlNtuI0G+4o1Tm1JnelXaA9f6dYADAYhOuuiZLfgeUR3F/igIq+H
yDJe1X0LtRKwakdOL4Hu3eU2M1pr8SkB598TJWm2emuaq7g3a/iY0pka00W/0aBv
s5D095vw04Jc12QCDvEmtZ/h9bZ9HGqmOJ1nm3eINEhHAIdpDe7oOGJwvmUveVSb
x6UFzq+IkfRyuh6wrrJ+PbIqBaMdQBdAzpowGt/rYNnzU88Y0h/MtyWDBfA0mCU1
91fGOGXRqMhKfoTnpKko2QyV7+om03ZPXF+E2bccIcBLhiRrMQCcVVaRCJHYMOVt
PAAulBjHby+qAwQSAO9JvbhrDgB0KPZrwg/0+jnxjFOhwJWILU1kUEYd9GCVz7t3
b8XfcXXEKDmAnaEMJPjRIvROpIPbGYUn8pzYnyeQQF4Z0FCtZ7NioipceBIQ70ue
T9cH5bAiED9QtMGhDTGl6csi7/yW45cV0SrDTSUOa4vIYF85f/uAAHOVXkBEPrWc
m/py1aOxy9tkQAe7QPDDQ7N0BVaSu2RmH+Xp0paeENwW9IEXVLGqucuhB/25lhJy
Xml1SPYEz2ziP4QVtXVEdENcn4d4qu31hx8Ms0YlaouzrW7Be/Z8SpgXMy0Jv5Oi
X8IZppF9y6Gc/2zj1VUbsvtXEFiWxAgPxsASKA2p1dYASXhJghyesq189kQCN9He
Au9F4KQEJuQbU5FJgNtoNBjqPeMlha2klaT+lNQZP01PzQjfmjqEYEGIGozFxGJa
TF8ufO+CQ6JYx/pLIaBULuFECSLx/GMeCwvTDgWPkiB6VPyEckTgHNQXX2AEXNvL
uhwJ4DsjD1002AogbqPVyf3bore2aqj3emLqMjKgaiclr8g53tddXrRF+ogxzbFU
iXcVdCtD/Mm9D7bfbioULIBIZY4cWxI0nUEQ2TjitCl8lAYACHYeCg5+xubqi015
btXjSWxg04008uxo/rZqu8dGMpq0T0376Vq4OjW4N6C5Ofn66AUXWw4ORjGLk0vH
55t6mjqueurbJQQnk0NUbMZXKp6KWnPX5tmOKCCKhqnwm35CPVHCA9/2yXsfcT6K
1MEUHRjNOvlsVzUU75eZ9EzWnytVzQ27U+6HGk3l7xML0SCmLVvN2eYMRezxN6mu
Yb4F5hrhgwafJ6JWX758n4lkNbvg+FBndwCKGHPwsWYNP6lMvtamMGr5RRzH/omO
PMEUWiU2eXiCF1yoMy2P+0WgTSNEvbeWq9D7ofZ+xTRksKKdAq9dQWdf3mn0ik4K
9DxP0hznJrCNm6TCZLFcVbDcHLPAr2TskCfeQVn9q9LLj4ga0UN/H5qEEURYyyLs
32wLp5Y2gV7QqiBf40Pxb0B1g0teFMgOgPFp0jkozkdFjGMiYU3cUAxBKblhsrxM
hn7jrUTLnZElhld3lJ70EGwdSw4uyEnOzgRrz4jUCzWQU+XgdvukM3IRccgXdL3e
nvsU8ql0WMXP8HLV0U6KYbeGSh0ghHX7IjvSCqm/L96g5wuyjyRKvO6gojhIGjUr
JJyy3BEU+hd30L5rdybu52ysn0R+9BUoo+2Xsr3gNxMzcuUQ77/UUABlFTvE+APu
H3HdlBk5eK5fSfME8CiIRNtGDFE7pndYH5olasggCpQGIpLrCDIq1BQA+a3zJ4W5
8k3hWVpnrRgXuDpNQWmwl5KD/r9FRZy7y9Xl74zvmpIPE9sFhuEyZaYeL2rhQDsN
/QNR6jq7DXj6ZRwUwcD+BsuJ2hhgeLPLlfd5X0W60XWyFGce2ci2KkeN1RJrT/20
qRrHUNTcgQlWhSsTgD15ClpHnjDpxo/LkldIurf45snRbtom7RZllFhlm5dfc4/b
qUrTgUFrx8lwJPrKlg2xhTLssqqy2DwvatE3pORNyg2TQtcFGDAMBa5/7y+SgGUO
huJZ/IGMgTWRI6OUbaKXt+c3+yDGacrkauO+st4+G77kQn/Wej9mvIcUea7xyVIw
WRn5xNN/tPgnOsJXmPAE51AA6wH5WsVNmUb8dHlrCRidaROXIYFyug8ZrTBquvse
JgNIS0RBghZbXnkEVruiLp3gSN19Vt8yIOUh1zLfvsLF8ca/GpzO6e8aecQRPs9z
/FavCnk+AtobwxO/LWm3cewdn0i6wiYJctKqBx31pNmtH9XcRZvK3y2bLe8i6N3e
YcJVo2W73Pv7YONFKlw3fgpBy/A/T4Bk+Q7kaFWTppJ8yg0Z/bBuXCYSTDQm1HKP
AXV+q+2Q/V0nzKA6O+j3y3TWSPxUlVc6nR+F5Ks+fa8dfpEZJVR5E7axp2XfcjD3
qvVh6KBhEPgbtUVmfZGO7Ybape8nT4xJN5uQzmClwr8CdQ4L5QcCC8oGmG2zf+7j
zS6ET3H7YpzsHECogqNBC3f6TxW7umDe6Z/ozD/NZUPfVRVDxA3UKqtL5lLmWK2n
5dkZOhWPi2NAhr1jastaaaX4IA7M3/oWaSngYfrgCYJ+z92Woaywv69MuynafsIS
LLA1cxy5jX97E3NLbP+2VCfxlNWhzfHTD3Z2HOpbEuzJyrgoab6JWmKsU5qsfI9B
dk9u9TIM1bJaUh0YIJ1bQKUD4REpz0AahO8eZlalxUZAK/pfvlSJaD2uTo7ilJSI
2zyLSn46lhkK1mA/+oSKG8eRVnjCzHQ5Kad7yI4wxulA2Vgi3rRKNZfcXXEyCwbp
DfmI6kvVVS35OROxAFS2vGrDbh68oxcgXlyRNWjpMakj8Q2CH85sg0VyBJATsro0
n9BqzKNFDWO9/j3i4aFWXTP9IohDw6J7Od75PvPhIBdwwkMIC1Y+LqMpU0HYMbyE
1C/DUxNqHid/VaZjtsE+kjTWvClJlBmhWQaslyxZxME9bxzcVsHOtGTRUeodsNWn
6ypWWkTzozI3Tc56BR3CKZG2vSGMj6qVw3HyR5TVFLKbHEbPka3KHwij0I175wYi
5xHiRyouNGmDT71xa/VaDSvPJiIxo/yGgp15UI/Q8c/vKF4XQFQTf8GB/BwAf4Wx
oPK4Zt+em5ptZnSRSfFblWfxlQyHbqAvfXRMo608tVSMLWotESPeOItIBZ6nfcLS
8OoUTXzAaYFo6bHDrYvlfhgRwqRr9ERACW9LajYI4Nl0vc03FJDe++VdP4AwYvbq
XAx63jPqEEhhowCEiIL8JR6+locXojWsA8Evbh5j+w4TZl27WK44eEZHwCD6GKFc
B068Zig+/GZEs1OUZTPnktY48icsv0pQbXtCgxGpVQjvBbmQn0os/7/nPfG14Zfy
zYrtvzrsXh72rpYswYAmUXISO6v+UA0onIQ1fkp/6LyvJZapUjVLN4Au5A1g6+JM
8+Dwh0PcCbeIlPu38LdaIp3KrNiC4AdmIR71mrbHAX2+v0ibsP2S7UwseLaMm0JZ
3dcB7L6zUCWFRn8MZ834Ex65aH1em7w902qnSJx6ZrAtsbJrYWx6tWynyZa3w2Cc
JlycI7RK7IB6zv7zamfEnz0scAoTy4LO8cA5SoGZ5JEBFa9Hx3OfPQVAN6yN1X3R
TgzhyS5A+SGk84K8GMfpwW4/f+KE77nsghoN6OyfZ/P0HfjUcZaX36cP4KSOaOQ7
U/vLF8WKJ7rKgZHy8JQgANUcH9BHRovPZA5KRm1c0ZMtz4OrMwap0wkFwAAGgRNC
ZQAz9vU0GeYJoudIMtWI+uzDFxyZPupUH73DUkdYS78hVD6bg2/TwOcuZrUJowTx
mWso0cVkSMAkqnEDHpZTNclSaUYTTW9ggiTz1dsVWTOhHEM6JDPlzs4Kb2IFc+hF
ADwKgiogF4WpAcGUME5CA4yiv24FsB9GfKQiTq1tbXYxQ59MdcRsgNOsk7RKf1/c
J9g8tOoF/bXQ3+sVVfmZpMMcOd6RdEAoPibMjpZ0y3adwapYOhALKC5EIuH2gNsq
rpPxdHgJTu9i2CLOior2QWEN6eSyZzv48cNWhhdA+JlLVk+AtQKVweNBxTwV0I0G
4XtMNxy3q9q4lL/J/toML4AuR6X0Rp6gsBlzhVQ98SzVMWfwlLZeRPqWxdca00jz
vqYtYgJ7yFpknuqrJNc6/fmuTrS180DcWgxslqH+OHHQpMaofCMbKj0vPU6Wq4YV
mUfUQae5QzxfY2PCZj3tIrljPvJ/SiPHm/beEiT3IJGFjC410gzftxDB0z5c/AWf
GoxLYeQfubMR1+Ja6peaCt50cP3l0/KWPXNyDjWl+I8EfRd2JBxjH5Sl+wvu+VGM
L06/hoWoGbOTPubM7tnT2YUO+0LaV0vjtRbL+m1Uy7+0IZFAs0Xmu5ZCLoCkon+Y
6CcvMkER+SthqhtIf5hF5QBWsyBIOkg6YbULQM0SBoyO0w0xxlCIyXPNvsITLbtL
+YRqzuMfHCL0BIWhcAF4YKJKpoF2PzMqVWGrgrx07EKniPydPs+X5VHZflGSdiJP
9U8YUV12VMNTYUUHKoCcsrSJCoWe+oWNi1Iq/5vk9+U72U+dYd5JvQIkfPNm40c3
BS/tCp5HfwaN/3uW+fN0BAVg/NS09EAxhTwsPVbqa9ujVCMQSlRRdVCZzOJsK/6b
TSeOfjgVrVbHbbzKSo1/xTeI0a4CPYAzwrKesY4AGaq0SAzQXS2WfXNdzhpzWjmZ
sPz3mHXTmbI1SDsXdCwUmft7oCPCVMfEN5Z8Po9z1U/+lgb67B1A5GCtbibKYNlm
OgfO/oqSoq88GcmOAIFFVuEjzDv0gWnlManNYHahcO6EOoqsTP5vDGRhfarFQPFe
0CAF8RpgbtknsHpQmeV8NF0efa1ib0dyWRRTtfv/dWrwxZ8hcgZW41AR5g/5zWXy
6w0zvequ5xUznzA0W5BeMayb+Ghc+0NW4z9yaTM04A5h6tlhk6DquJzt8f4DltOq
S7O7kpaIlneTj4LCLKq3k3Mh60j0KtWO22SFz7qItGgnaK2XHSvTH4m0Kq4B372B
PUDYM2lK2uLX4Iu8lkmbYF0sQRkkh7op8vulr8MQJzDgD3200MVmQEHjnjVliZBx
8eLYWkiK5EGj74kq4flYkD70f6Wk/0LFEHiwe2T3Xe433nnLmOecYvWM5kjwuNYY
5MCrMt3zdFkNaGeScBn1yxx0zPAbG9GQTjrT/YKi946nimzDHe+cpefpl4xfyaEG
OX1T+uDyVLiYj44ZTJwcBoBablyQMs9Ntzvade/BQFMjbKP0jykj/LkYvrLE2u+K
pL+AE7VwLnAAVlOBaaU0Cn7Yuy8JxAmMHPPGXIkI7TmcuQlzjBqvsdJTlxL8vSW1
pPjFDysuyTZUKLfcnVc7kf2RiuNQ6dxFacMn+SFyWE+JCFiKDKjgEh1+M4L3eH8b
2WwW7RG+OVD7nQ7SwWr99SkAzsfWX+oUSbJmfLpgHDPNj4NHSZvpmbIInqgRDTMg
+Re6pCm8ELgbrkRi0nvCmCU/T1Jc1hvYUJjVbGU8mQd60m3vsxD29murfj0mmrxZ
FDJm0da4m38HhlTIfdl9MRZCkNUbkctE6GH2JIyrsURtzCyoa9ozJrVFA/pb0IdY
JK5Zm7aAWeTEYvBBypFmUUPjcviy9/OsZUONTENSwpOQ45Cf790tBQym0J3/nZJr
fDuOaGNNezFS6qV++ab44XfxjNXssISAfs9x7HUHxaVbQPweqFO5vx1RfaU1oNf2
m5fcjmTby/hqxntF4r58E9cWF2v+I2IF4TDXR2h2dd+EQoR2P++PLvXFzjWz6a5R
QeHc/rVkJZlhUt0/QKKTczC8n74+wGTTg45MfXDZtxlOhUGgdB/SEJgI7Z9M4VwB
dbkOr6s0RmpKcBN2r7GIsrgj2/q1GMVqT68eGOnW+vMAFkjD7qAk8uXmB56cjW40
PE3kZQVmxJ7g6O4HrzD7+3RVS11BabO3DxHKGqjO2T3brAYDs/9ZONUa7J8bW+zU
hqrZxvu0qj/46BHshHWD9tyrE72LfGs76N59Ja8/uf0GtcgCnHa2gpYCXs2B/+qs
pW8cS0alI81mUMWylwujGVg0PM41dPXxobeZ9K1qjigt+/wNXhfO5ZoEYvj1thoY
uHj0rSoLjoPzS8TiJxlkxG5PV9Io9E2g6axvpq242a574xpsRn243wl+8uDPlqdg
091FP4Q+ipAC3qqZcWQCH1ZlTXbgNwuOhyIpFG9h8TS8KeyAe/dLw6CAQguwd3mN
OV3IrzO6+qwykvejxeZIwYgnbWcnpR+6KAMV7cm1mYlF4nR38U7HD59EBvd4+9hm
xOvaXJa8wLck0Qs4sNbLxx86zFPwmVGpL7Zs96BnP2WDgSif9PyWqTR8+kZtW3ui
DYuQxA8TpX/ls+Oy5JjKPdJiwiEZguuNjbmNCUDpoEWovaFY35mZbtCnaFokQlRA
IbzJGPeJR+Ca7F0L9y8Yreo7w7tccqQr32SNE+836G6qHMlU3uMxxhgi8lztDoXt
KBNf1VByie2Af4sigbDFODomyx67xcTGBlaYkIdqjf7rEtdxXELZFIrUP4MlUPK2
oqtqxG9oYCK5f8rv3rHsv7HMNThyoyL1bJvQLAEM6sSvH8V4A8nsaScaHuA5AAPZ
eOpeFGmh+TDI6ptd2gdT7PPMguubDnrEUV9VFNedkunnKGPF49NAzE1VNodSW5Dd
y0ybMOmYXCUbMYLFfFkcLXf8ncdhqCqYohmybwKAYLGnUULiDkw4odGOIpvz4Tqm
RpMo+hPXUaUNeHvlEZYYlcPs+/TpF0MfTbVNOvWVWtrArlx5/WvnDYULsAEHp7Xq
MWVbsWHrZxY2A//5ZwWkVi9ruv4kCHAW2EfyIptn513w3Grl36ebXquqPvO4JDaj
nF9cee/SYv0ZmpiYvWnioYI7y0r8euKZEUdzCKMxzybae6UWQXEvC+TUIK1mLYyb
YEJr2v0o3Z7RTYZq/hSlvrb2A4tzCqjQeIWJu2f59qiP8m2IewlWPWYbl2vItMKC
b/Y5tb6krtHEBfBUX43RB1BYO3jPJ0wF9ckGbUMpsVXh4M4z6CHiKWVZAVsDsu3o
AGuZeBroLeUIJWM35WN1Cs5mn3b/xRZF3yBmXemO6ur657odtS38VIJHcKcr3w6s
9Y5ScCXZkXtbOiSkUWGXznUFUAm0Li65u/Bbjx55OQpL1gkagnRhvE4Msqej51q4
JffxyXIeC0q7zLAqLnU3Zu+OPqBTNj847jtypqj4Go8kIwIn5neNsMCZwyCJi5tU
OxfuQD5HfYwgIyU9c+vm1+lwhjaWlyiUtaqyq1hv2pwqbW0XSwDOqJa6AATyurWp
Iw68cgYEje2EpZ94nsOzNNJsVkiemc2cW1MO898mps6C57QLF/3drNXiw2Ydc3SX
/+4PDeg7Z0vy4KO6z7qnYOqERDRBOuT9b53tIExetAmgWrnWzPx6eWqncTT1/mms
78zx9VIoP6+Bvp9qwN5fhKaUgYzODkY/3DciU1Ol+km8eWAPcS1ufcpjqLQwNWZz
MLrYXhCUub+rnxlpidkj4Q08iBysLlOK7Ve2ztmz9/VoEnA1ss/LZDxvBb5OHPd7
H+3kfRFHvyxiCvDyjxEXAV6XdSauF+UWhpTlR5FFsdhXDcaRnUUYc1s+Kr9nVs3H
XAR1Kw1O4d3IMMZVxJo8IsqJPUhKhVyV8twePnXAsJcO9EO/4tNytIuaJXNvVbIo
4shuqiV1oBwbYBe4gAzftDaLhUKoT+c2F0OFZiLNA7T5XZlrOgVMxq3d6kU6W9dA
LOxDf+L6kCH0UieWHNEOOpy8YprKJO1jN6eeUex2m5bicIl9ikvgEAQB0PSbvMgU
jnSqEuau+QJkcmxn2/2KPkwNV9wh8UamLv7ZIgNJZzGYD14LOi7uuCp8edBAm3BG
BxEgW1FscTYMh3cFFlY6MJelzk7ommYeeAf+vu38oQzMrhKaa2xNYJX/c7jo//9R
I5Nc+92uufxiMi0xZ8tVRO93ub/VbOYH6H7+ZecuALWS6RtPYMtr28PC7ZSlO03J
fMsqxkRqxShG9iGh6Ib7vJK3tmuOgsrrdwU5g6XeAF89NtmJEWI/PFppXkjAIIzT
R+ihHIyfBQQiaK3pWcedp6KFMCPgfD/5okjwUl4dkmQG63Dna3sHk3rQVBihHpLh
2TTo4BH8gEeTY5dOFjQ3aZ5nAPszRqDBdlY+prEIf2qY8GgRrOxum4LGCHs5fOOI
kgr5hY1PWeted0m/4i1O/Usn7ra52hKZhp/ENQZrmxFqz28dAhJKZHhav5QGDqdm
UITvj3cp89NQlGXFIFrqsAMtBHhoAB9HCgxlT/HH7ieiGdgQtR8+QO1qVtOWk/6z
Hb9J2xTpbQ1+k2btxnRsLN7O/NGafvKeVPZYqV8tTEEG0NjayGcjA1YLKbny0WsY
/2IAmFTWISlCswAjYczBTmiSYskfOYCwouU16dikQ/NtGbpPs1lqPAkC+VNylPtu
oaT1xNEhWIldcdJWoPeYy4TAEOMJj20w9wm9Ghl+Rfy0PuYRh0O7n08nK9ZALKaV
3ECD2AcfjEHH/vf8mOVilWuZ2ayb8HDos5NZtgqO8kaCnwKkZDK9NGgq3/ZYeAWK
Lqqr+zFSuh511DPnnK2T0RTUSvA5n8gNONKGvWPuyJzFFla9XvA2enqK9yFnyG55
wPJHQaYQPhw12WlWoYgddTT4u26G2ZC1CD1v9ACy/6agV3EI7n+hDJJJiQNwx18E
qWFjbs3NnVcxnkpL5a2W2RaMltdwmiZRAwXNWJCdKNKzHyqjueBPotGh0afiFWHh
wDPuZ9EXUQlt0t3b72cFw+Si5SigMetphfhFCwE8EXkQ6HqeZBteUWGR5neP1vvL
X1HgB0lpZJpuGZxK3E/0wzcN6hcZD5ucGeAKE2nd76yHidJ/YeYLn/uX4E1rQTs1
r90C7DAcJ192d/QqOqA+zvTdjM6YPaR3ar59NBrYbG5PEZiaaFkJEoe6nnRtXa9+
/zdS0SeZSbKtghhF1W+J6TLuDfA3/YENkp8WEgRCuhdzByiOyXJ4aykCcjTPCS3P
Flz33t6MqX9NpUfIT6qfgiLYr16gTh8zK2e/hOmzkpafUVI2EbsTPa6QGYPjhdTE
WFZa6hkeuFCUAOgFAtw2JVeA/5gsgzT6PF30bWWb94IRMkOVqvS7gKeDr1OElV66
DhXWni0ZN1Ivc53BotJxwue7zXqYynd9A5uOPD4n9jyavajkTzQ7AIbnYanHnzQt
I/7HJPhCaEsda20emBQLdrB/NKDbYhbsrx5EO/WLrvwFdC2Mkmb9OWsA7VgBKypj
TUYNfoJmMXHxxEDdz7Uiu65+PJ+nEHZMjXG6qWKI3/qGryPQ3se7RG+qr8/3+jB3
JTsccnU1Yr8HTs4tqj24wRdLgt+SV/DK9tSuMgai/QK8QSTWx2NwuejTCfSe4JDo
bTdibOKCtUuUb6SaPgd/YxVERsoIHUE4gOugDyUTuTMUAN7CpgLmF949t9sTRdcr
X5kdBlvkewklKp6FeIPe/VkT610wCIWdTfft8IgRhg7HKqqMs/3scgay3ZNhhxM+
G0SyGJ0Fn2K5QJHLdV1zK4U5znzhI9RrQ9/yugm4FLnRl1mvMxxqu1g3jda6Af6h
zv6BTWCNSuFsWFX4n2WDUuVMWUTDvNobem40WaGaLhKJ2M2esVmFpkjDiDjwaZAp
kHFpY5L1YEanlJVYQLVmGYSE9P2emVWe8Lt/T0RIlNp0mlXZmVTzX9ORMU21On6d
TW8aCGfVS+dIcLlL24pSFil1wmYVqzgdJ0oLPtzmE5WjLt6fuoQwIZT+ZYqwxh0/
MLlC0Gac5ozli2pJALBNBE5x2HydHB8qrBOPnAFk51xcft9Uo7a6eYsVFFXrXLYU
9r+UtdFjuWx1K7h9IzLVoyaCnsN7NJVvFuwx7GOWR2eWZ7YetfziHziPClDaDtN3
/4G/9hCXat+5X2tD6KQckwoR9S6/J4kBFUBodyHDQWE8MCrK2cvj7ljZJd8IOTHG
p46DheTKT4QL+g+/jR+S6I/61Tj2o3/GQFFVCAJxDb78q6hjzg/Z1jIWtVFIdZOi
34h+zR1YgNJDUVG+QQYZ9og9OqFGbDQPTLRyCAPNQFXyuoHbAS8ZIlDvmvnpq65q
o6H+cLjkfeonugCauMXEiyMY2Hz+011uehFd9IO2WBJEVj4x4QF8quSa6g6OEto6
6xBkzWdm79TOSB8LsylgpW6m5cjb8qg/Z/kpQB7fSdkhIYbXxDqNnaqoK5vMpiy/
ZrfQiMfngOLWE+IngP1qd2LsK67n0NFFCWbQ7hjlJWdcDVDT4M6XA9/TcsXI/aWB
xZcYPxn/ZkK6Al1p9YGwCTTe8k2JxeASMXzsz3rL5PaX+TUDj8iFDGMuFmF3UEGk
In8CveO7viH+eeIcr4Ew5RSk3qMQKMM8B/Whw2JmXfi/HaK3o+VDR69oyC/w3ECu
eOGhP8cXHU/rDwXPUcr82+YBPthoAHa+Fe7hzRuhT80juMUYcmDiLRrjSTwOxfJy
bjcGw1e7dsL9qm33/Yvz0aHtpR001NUdU5ma/4En5upNcfWkAASI2Jl+vFBLe5DO
tux4+Mlgdt/qaYDkCaCk3iUxsJSIoKLkgc16EMO/ZCxLdxIbAZBDVi468lla1gZd
wq26SjXu9BdxTiff8OOXL3ntM47FA/Flyowed5qSIHrcQKdSTyJZlbV3Mf0WOTZA
B5OcPtapC399nWxflFPGUeLTMEI4vRRiGxblwh1hzSc0FRiroghvsQ3/Q5x0CiO8
RdQMZiA1EwyD6K7mx1iF7ugjCq+Y7Un7GsV5q1cOfEBnJU8YT2qo5w/j3H082OCf
DNl18yZHKqmCqrvTFsrijyB60AvMryRIB4ozyZ/aHqpl29/3mPVTgccD5BqHdRpX
a0QX3M6LTcDDKCeQzOXYQOG8caLsTiYz7PxEn1dtLuI2NnKSiyo53BQiVUQC1/mS
ksefi/RcmDjE+hEKgyfky2oH6MFaHZlN3e2buPOM5VSXwM0TnrNxc6aKae1D5WNa
snbnlKfcJ88XCBf5FxKXp4ZGkrtGsMFUr4WV4R8SnQR35M+9qMIJybj7+PXOiCk1
DJeGe96rt9YjQetVlosvgGWxMPny4oOKy+hdEjjzoAv5t6xNy9V2OHNShQQewQ5t
3AAlzkXsSZ0u54zbMWjvlsXftKGyJFNeNiLZilJ0he99nGS1J0/j+A1pzwwfN3Yt
V7KtzXKBtmfqLX0CjWAtiEZQvykqqn/JII8Qjwq2cmwzzQ5u1iXdbdtiDr3LUMeJ
F6+ogi70O9FmcpBCfJMimH+lyTYlZocdGORrkSLsTNF3pVR3LLEKP6vdf7gihbmB
Ct1V0fY0LCAyjmWBpNLIU9QQt9+vhJzzGS9Pw31eEJjAGXXg8IMUQoU0dc508FOg
toq8DQ+sMGzzypd8t2ldWqOioKG4xC7668H+GGt2uWnuB9BaHr9zzBTWs164sA5H
n88DlQaJrxd7S0wpynNnj617WVvyNdc2+Tod2U3vcumCCk/4HJu7TaudmG4VOJBJ
eBmwygZPaD5uPMF//gIH2zcBa0baM9fPiBu8GmKmXVUUPbKFHzAQ7iL13asMmEJL
auXxxh585AQMqzv2kMqxaDf1dwZ8gyTB1emOPtFBcYSLu3zYpG46rRk2lLnYMrCu
MzDszwKqQUGdkJYcst79Y7ygTQo2qfG+UVq1G0r2QY9ReOOKtjIqe1JYEOTqhgr7
QIZ7W6V1O5gwftCi2fza7eEe/SMAS5BoKhObs/O3RFjxAMg7dfXNNrsw00GR6ox+
8+zw7nKoL+MQ3NadWPei8JyilOw4RcTwLqeeaC6DsFba61QZ8+4pUmapRBfTz43h
sZkC0ilpwgZ/NJ0faSq+XIkAnXg1S0ndjWm/5fOt/PVm5OwC7+inxcocPZyhCl6+
swymZFXwXzOzIOGOB+bqj0Ibxe5iUwt/UIOlAwDM6MdCQ7i4YmynSIBr99GQmeqO
SlStxTP5mSqH8KUIPMhLmgermMmgienD+K4CT8ZNiL6xB97mcDyKr/dPE6uBgqCa
Sth78ltUhcXEIRN0HDP+fxKa7OwnTDEPzFZsRT9O1kD9DVZQL6Ev3Yd9uS8RlA7W
1U6ypWM/OpriejFRJajH/ekf2yGP3dBjcjlzNhm/uq/yBqVVLq4TRUbV8Vx7Xs1N
r10rHaeM/dHVYTYSLvbVYfNIqhl5GkeJkO0OsSYRjshNnfeSZTtKiHjimXT/VU6q
pjBT8TUs1a2BLXxHw/ZQdOgRDmTN5GILXwy4nvIldsJAbch6eAfMB5cj6Xb4cmkF
akQxEH6dz8uZ79YfwHEXOhfEiG+4pVzMSEbV5PE0urfPjw+gqR/XAuH4DMDJvoRv
unN9TYcR+XFVfypltI21JiirQIH+6o0XzLa4ITjxMILfcfzusi8zBd3CfoUY5bJX
0SpxkGt+3OAsKBhw3ZBvvIjVve4ovVTODow6B3TCD43W5bwY7AZUPkPuKAeMeaM4
IY6wIjBQFcXLIV6Fe0MTOiu23/M9DbcAZxQuXcZ9AK6bwVSBgSmO2zKCVEOHggqN
+Laflb5GsHGbKW1sUW6ps3LFjJzHLwwl+I7p086C4xKn5qewb8Jp/cHE1m1muIfV
39vhUjLJnDm/FKPoHO6RX0NOi35VUmj4Au/RNBGUVJKL+gWjwCuMnQORQKUyoqAO
XEFg9f25klJ6SAt9nZOZ8EA0nVx32rdDQVRyt98IvK7RxMrsIV+MEdgJ8vdttvRC
nLgaQYHlYi/TVnCQ8TPLKsiLaaGrAYX1dbTax860LYSlGs99F+ON3cH4TF1wafCn
UGumv1JV7e2dsaBMo1GMuyCowhXZpDJlj/lzA0lCJLR4sAs/NxUiBklmapJajI4j
ZwZeXV6SFEnCsNLe7gHC2Ryb8jUewJRk0juQgvV/KRwYbT5lAuIcvlYG1fZIAh48
1wdb2Im9dwSzIGpEYlX+XIm+6U40jAusmNFbHbR64zZMiOrast+i931Rj78GjLCC
NTkXpf1KdKrDho5OpwQSFw3mw6GqZ65xZbbgz/hkfjAj9w5TMnwEXVTh0IhjzkU1
HS+4/wXOc+bN1xIQ58sG5Gnwmj2vMSBdMvmWSMetGP1FSZf6RH5O9DOUGzHpE6vU
g9k5IwkCiJ0z71trOcegbVi/e6ZTOv0eDrDKTy/oxvMJY3Ql5t6L0yR7LTJPU2v3
R6WZnf8R2QWZy2MUkr8scPh1Eg5fZwCEveQzbI5RMIOeoKb5bT1w4FQKCmfTlP2T
EwTMhzqz6JqXg4Qoogc4pI9xWA4yvqkH4QORuExkfjXqag9d6uDC8YAj//KP7mCp
8iR/zxZNgYKhdTbUxv3O90YD9iFaCFh61BcPpilKV6g9Er2ne0x9AgofmoM+1glO
4EoOMgTJWR6WDP9zWn7SNXeRCRcP3h9e9RPqy21W75/1M2oj87Hey4WMXHvkokYk
wzv5zaix4Am0uFCq/AzvyjwSC8Me2ArmjhdA2mDsi1GesrG79lFEd2XjSyGQ+7Q1
NeZU5N/Ja2NzRwKBqhjpsByqAh+CqrDWgrsZbdxJC802TTVPBjW0d2Q2bThTheMO
CXZuOOVhLOHR3O2jUEV8pW7gS/kdBRStcftoY4RXj8pvor7uFfJ1uTlNUIRnhzVJ
pK8JwDGuBhe7+ZFmpIwIFecvR0wXmPlaM6dAK0cA2BLPDQaF0kBZFmOQpz+gpjhF
6Nimyj5nKIYdR/9qc2jJ/S1Dna4xR87nBv9PJP3LQTd0rWN4/gFjf37/hsObBXwN
nFR5Kl11vNpBHcLh8RqBoWxcCgaS7hsBF9kNy8I97Ukf1I33k3WR8wXP2BEFyteA
tTP3iv77A+9QSqmkE9we7iAIVDLTgLhyqIKWK1gkMC1Gs07gJavus35BEA9/9MHs
PKyO0sitp1fu59+8uepyCkRkrhUOPbYeYzJvQ1/7WlX6WwQresQPjka4VsbVCGoF
TTnLDxJE6LbcEzXcRIG/98jbJS3ViYiaN72Yl+0DC6oregEwcqLIL9cW4hZpABS/
72bOrhqMDxan3WNQl0JWD52AZK5Myg2v6ozFaHLV1GiovCoPpHGvd4FDth7tbm3E
3Rcb++F5KNlhHn6LeXoyMwywilplOZ66t4TLh0+BYwl0s2NQSFdTXo7OT/tldTZw
/ACGvLOeqE/T4H01mbh2ENAMIqmU8U8ab4vsWn0bZ7b+nPGf29TbQCPrfiEHs+hH
dPTl8KOu8C1KpzDshUVchM9xfUWcEUByKyDhzipRK0nYXgLfy99zJRzqK4qhaOTc
6z2df4qJWNBF3Z26lyG8T2S5Qpictq+wviWexE/iSFq36+yCGZK0WETht94y1SI8
IWCnfxO8dCfYhh35KeYLIEtCcTJKspbYLSmrZXJM+uFqU1wsIvo6yla5qypI6Vaq
7x6TZD0N/LIEaidbRYR6xEvYO9FcfmqH5scAyAKFCTcCcU4mTddPvAPm0VChnjdW
S0g/5OeqCmTGOBV5u7PgNkt0xBBmB9TdMjb1eoclOb3aY3tXSx2JaJoewEanSbCT
Al3I776R9OzhVF5uZoodOVDPJWhCfXl1NKlRt6IyKdtxKygeonjnzgJfW36jP8EK
kZwiHcVGbiz0cseCESZK8uERS0tkBdBBS66cf11oWzAHo6Mg54ZATNItlFphCsWK
VKaTEWEmYDkz9AFD05IwBh+iRiVYfZs1enJq2k+5syeb7iloGaYAAUuAlZVL0crl
8zolV5UCHfUARoRu6FoNNris2+35supM6XX/M/Qyq8QZuxGWhhpceiDCfij/p2+J
N9zfcIJm8lMZVL7c14sL+PJEKeEtvZeGoM+bF87qZi0taHrvmCkfG//wT9E8YEgJ
V4VK/lfTGtGLQeY5OkLObQMByj8jYoO6iG91Ihl2tSHYWslEvHjnPxwSKPg5z6g/
9iT/GWR+M5jYTldwYxsVj+lxQOa6qefbqXjgZ40z7QKKuYOprLxjS+gSgfkV10VT
OsXtSTRg22UB3/rlGVsXQCseTPrUdPvDZsFXAAePQLtgXG8Nzmt6NX/4SPhkwrHk
RAFk+rcvRSwRBACPwN5wOl5Tk+j0xp8XsKRIU0W8FOeqiOPSekcMyvkEc5XNe3tY
K0y2qkU6bKVYCTUEI3iWNemLf2Z5rWusjR+m1xWTmMvNhGoN0JkSJ4BlaMU/HJx7
KLuKK1xW9Nk/mlPWKoQoM0xQv0Ea4H+lGGRrOHEVTT7IgNfc+DwCdHPvbQIqIuel
mbdBaHlQwAJ0thgDo4DqAGy1pj85wj2VGbumd2cna+HnPEEJj1VfpYpM2+R+LWkD
fn9+aKOYiSTkbTdqZlzhXqD1g5y9w1HnGA4dcaPboQ+MZCs22+QNLj81UNgKgkwA
i/kB5DZ8d9h+KqpRz4JsgBfpg2RbEpNGnxbBn83Kr07lH9MgI4hTJdqgrsBt3hiB
Bg/CJgzso8iZzemtDj39NSvQEvcyxeQ42mcD/4pGkcglT/9/gtlu5fkeoBrsYQ+N
Unhbojpvk7r8BwQwmpBSw7JE/38kHiS3+WNhUAefFUkTer7zkO1GXwtHO4ioKKK1
xEPNh0QURgYdYQyGkubbkbm71/4fjnO1/48lSBnhXAzwFbzhe0eL426bMkGada7z
mY2AuFyj+1unQOXPH6m9A5ESH0DyZ1ry3q34Eh6ma2OtC41xqOuQTHBw1dGG4UDg
qIiMMpCY2gI39ngjWAlkG/KU/iaC/nzZne98PeaAd2agrisAybFXYHtw7FuMnGIm
xLCq91hKiCT+/jp+Y9BCCCq6zZFGHOfyLu4BVMm3XaBGzQyUtqOZGobCqoOcBUhl
oLW4ZUBOTjd4YPEIJxn4AxkEVFonXczKEaEdVjiNKUGlOk5aCr/DelD5YnRHtxkH
RFaF/J2wBdYgo29fKJkoZ2cO60O6/oY1tvaVyltgEfAZV6YGsQzU0d3uh7vfZs6b
zsP8OG8EIEAUxbjwJM8OoUDDQ4lqUQQRRhSr0g0Xbu9ivg1NImdS35uB9Jo5Keqq
FNFLWWx4I5+BKertmUclaeEK0VPnwE05ZyXYU+eWlRAndPg7UuOWpQG7TMEG2SRI
LGa9h37StLJ56EqBfE5EdefeyWZPDVCd8rXjOFMaLy6LkEZK3Dl2CFLh14VDindM
Fyx2NHWdio8CWCgoUM9pD74SxKRUUKO5lUWz1uNVu2EDjNkc2QmtCs0qJwGhoG2E
27uZVcUe2a6Tde7G1IAOoleC3ZE+4yYhut5OU0sx4C8dXPJrhvlrQZYmCX+jxqhi
6e744jPLBNwb5r3H4ohj2lTGDwBcKk8Stox5oqV2yZG5H1ulD05Or4T/gq24t/XO
89GLoeJvxpWxbPg/4uQHzK8hTKOetQyDyjmUno9w6QQlc2Ow/nXMQYiN9MeK2PJQ
Rm+lRis1yFvmsCNKFPEznEr+JTw8BXks7PtzTNiU6x52XzVrX9de7GpT3oaSojq2
A+u/YU2yEEwIZBItzC1s+rdQe4eEs8o3kIeWzmPglwnxGyJVbfH8D5OUDREus3n3
VXqtxKKV7eFaRnyuBr++AeYwNoEHOgqvBK6HRxWngSlK+GNdMM6/r48R3mbUtTbG
FuzQqEWRYjcKLAhrH7kCgxje4V/dCFbciDmCz8P8H4cT1irzfI2zkm01cvn2B8LV
1oSVi0Ycf79az8kcUKoFGoy54aemZbCOcEi4BxvlU+L6yAl1rlBe96XVg7n02Pah
Fy9RsKKCVPPUPSq6RF2+d4FZKSCVOt/HJ2LW/79pXyub0ppJlHThNc+pMqxCtHPU
FOy/48VwxKckrmDyAs8TGS3mNyNL5Czb/2f85u/Kqh4un+bnD7ONjXCU+9K7onSc
YytyM2nvsKAKz2ZR9L2dPlAlMAMii2J4JiG4g+1F3qg0w/JAKUxcfzW4JNAjuEyZ
iv7YH8+n/lgF3t/Tt3EZozrCjV7D3Fo5jON8DPGOEdJO1jBCX2QA64isWza9kC+L
w4CKRU2LRP+dODZg8OByrYgppDjG2YH0Zoii9sHowR0SnNo5tG6C4vG48Ws38C7G
bWvBvcXWx95pODvaelRtS+K6qJ70aXR/O0yOh7bee2M2fhFZBM7ahHQ4I5g46xhE
xcMEVQ8oVWb39Bfocv34YAr4PD+JJ7tQJA1YrEvk/sbW+1XxJoFL8U/aQ9GKUrv5
c9S5g6KrNSuO/8qL3QtX+lW5F8z8x4yAgIH9snvBLbbJ2Kaf1zKaRWi+NjLU/IyN
vIA/b0n12Gdo3kjNMtnfgnOTrqZIdHkGAkFiDVCjldaUaVWmytb4Nzv4M/Cocp1x
ErEco4JgNyntcIeRMmMZrRc1j2pDBCAmWCh56Vh4KlNW2lf2QXZOPvYlRfF3bDKA
P/bwa5Y9HA7KZ5A/4E4wfjNB6wTVi+JrZGWiaM8NDVO0Xokvs5wDThTG8gbDv+C3
GtgK+aZZ3He4ceyqzRvEXBs07ker7YLYJe4nxWtFvWXgO70GHBI2ZZZqB+zlVZIy
ObV3iDmdtYEoUMdd33OJ8s8VB0qhPDZ/0YKHNrETRdeY7qrsFlOPllylhCm8hVJR
J8okNFh9FdfvPPwQU3kLQ7pOdYrXV1xGUHohpSY7YXn4PUDk1/OjyGVeVAiJSheG
Qq7b2ajM9aZfNe0jX4t35H05vkOxiowR6aJP7raMgN1bEH1ogsLG2nCkW5XQ46QK
fQ1HFGwk41/VObNDVhKU1apMEdtIy8GhMhhDERX0rBdJrZU6ZCWSMX5F+LMTlLXJ
S1b1XGE3vfRNM4mR8KhV7i+0A0tJiKLS+6hkm73x+Wycr89gBed7z49ZRmeJeV5H
eO9xh9n1B47WlQnrEazyst8uOTwRx4LdgR1ZxE9Jnzbf4q3xMc1B5WEozzQvsat6
dZicZGbjZrxt4Rs+JsfagSIb/EtPYl1fsn9Ooj7wFKFOegZ38Qm8myjZQjIp3if1
ctE43NMJJpJD7MJYUUmHJJ+0NZcjsYfnOH7WDnkBylpIqzkPOLiV0idXkeH5rVNC
jANPEQ181KWPqMtOo3jfRrVXHZuQ85vpeZdU9twb0u+SuU1Gi5SHXvZuY6ABqLgk
Erb8cEA9akuRWdqbbVg3ATkbc9EELIzsrTnrBrTGk5VXeMdfbLTAXTacKP4XOLFk
oI5qRQm15CuQ2rArudYL2aP/HxDGLCSCCWekM+hLf9WlLO81GyPYE6eerkrM0irQ
H1kA3kpl5DQ8ptOywYwGZVz1L8onaBzABPd9/TTuLSM6iKLLDPTcQAeJj+ZmJGfE
PwDggppyO9l3YlUijA38XZ0fUkEDhmpqbbL7Uhz0eph0ZQt9iRFvxO+D6S0/GlUu
/nWzLYsfHE9laJM7nxxVgTCtVYSE8ViKxJFA4RJcirpgiuREmkaLg5/v1KoWHhAw
lGPm67A9vH51Kx13qKSDQaZ1F5ScHhu/ZJjgHZHAwPciMS6/+T4knPvPJPCdRERO
tBdj96GfcQ6/F5f74PCYxQ8TVs8qrqGOgztLrKfq40oeoox066vKdXx3kjQ80trp
mdkv8Hr7vzhqwlbLhyADn3qMwafWszJIdk2i2JR0qG/4AOAK9R2DGgStWacK0RyB
OBTlP5JH6qvlEse/wwShN9EIPRBekMHnavMJKYtku93tOFysbjlQlG0CLTmAnge6
yMA6x47eScvQ1LehMaVENk61Fj8yfxMbA4vE7rQ0FQ9jDJKUxXuY4C/n4ZeGw1K3
T9EaVVW7ydChle+2G3wIAwM+uc/aJeABvOdhr8sxAfp1Q6fVl5hV5BpTM+k9ykBF
OXV0uZmgK+2jYcwtI05W4ulf2wJ1WC6x5rrNT5OgABsrs3PT9XUCfMsAPvdWr0/c
ZBoL0xotM02RE4EmqZ54uUPSESTQDbRIEmm/KjE9rN2SWwG5Givv4HzLxOU97dMz
QS4pO2BenVBe0Ict7KZoCM9hqCn+COjLrhLxIcoQGr+QIek6XlvX5QhkKDXyzY7M
fd5Y21HVP5FmpW31pp9NHgv7eCi6uGc4l5pQstSLXpy47mUnfmDfn/66pkB0yVzl
XhY0dp1kB+iV5iz3c0FalfhnZXcYpEvEkuwKuCfzOeparSICHeNia5tGP0Ljs7mZ
lWES/FkE21E7TxpA070S4/8YntUsiAK/jyCMhL/OlMopWExa0Ru79IcXEKXdtbXO
WFe4as+KdLFCyOC0T7vbAx4IhMIV1Qo7rq/qipxSPh+UzExCMBKthWt0uUPEpfew
IF+eikMZCLYyxxHRB2wnExd24t9p+kRPo9HlFJhv14KVtpnE7SAWFLgG9StyjO0I
epraPW6gv8cEB6wD61yRoalh8JsZoTx7kQk8atsXpNdFShVFOL/M/jipNTIomBhX
l3EbamWI9zRRyLfP6XAJHIS9EDgRfYwi8lijA5c/rus6g4x0xEL5QIb+NpSo8Mb6
pI72wVAj97jStYXqShSf7ZyDDDMr94NJ2hNWrSkOKnY3W0gjh7kh2L/VOgSZIoBX
QVJlpfjOvB1cXruUI1+RLlf8ZVI1d7soCstB8+aULw02hr3eDqWQZCsR6oseCWBH
qiyk1BcHDeHpq+B97biE7wh44JDelmNslsBiFrmKlm8Dz4SNu3yhilx7u2bqNVZK
1y1ED+2EYf2ONnKplSALOzSMSBxxA0pw5vWgQesXLCTBEiPiMPrDKlNshgnkStXk
x8Treu74+oGeoCneSWWBqVrbeN7zi6+SPe7gipbcU6avYqu3AwgPtazJY510rFm4
XrxDWr3BZ6buAIa5nXB9jl9VFfcvVuc3YPST0LCnKsT+Ae5+CdBC9DpRvHoFJTzx
K0Q9K8tp3TnktrVs4jKJRG0qSQ8gSH4tQBfWsJc2uqfAeVQjHefr2ZXd4N6d/r77
5wvb/xsjpL8S+8nx7KrZI87XL0YE9TS5HoTsfUmUTYczoxWhXFbGUvNvs491E8Xh
taqpptHwQCmWHwiDwj4e4qD0OB0XaWQIo/HYKF8c4et95XHDzVhn9wNxYl8TbkOi
+2LwF3hW6higD8OG5WHOvszwUe6vN3vhyUf+0YYTtE2Ci7CawG8M4eNVuofYRZuV
QSsUK+nCWsFujncYKxn5eBRv3NsalcQoyqOVIt8FRq7PPJovIfSYRXcsEENdRREc
WlqQxNfcES9WcRyNZU+4ELB4OymMU0Bqu6iUDjlcBom24VY8UTRoNtSlQl9bNXXB
YXGKaurUzcihMx6RDj1Yh0GCV3dwJvjBY/vaYeRYxZPoDuBl/dpZZnZpusKRh0d9
wI+n+PO7a/EOIXr+4bvJNxyCyubeP/wqtlJxRzco35UfLukuoF0Wi61ayEo4Wkls
MgZRbCRugBGMx1BKhC0RmDdKcpZlxZYX5LrqW+XKDmONFkeN2lpCEv6YqQR7Re4x
cHDZQHoQyDxOQoIUDs5NzPsPMn7nuwEy+scMgfxrH+ldZCwnusZgdkjmcFROKVYv
pvK+P9srzLl2uSsDgDhXYTrxBNOwgw+Ci5iXkdLkzff55tmnHMWB5b2LntyzmZIw
Cl7fS9N2ZEtHCbzdwmmicNjwWKNfYGjzODIEYYP8Q95s1F/QD2dV4K5ygS3L3W9H
MtGLD4bQJoKY/Au8cDHKBDdB3RgEADhDJaTYPjUes00Ve1IoqhGrVkJ+3MXADkW3
j9V9CmojqOg3l4tYYwDpE0NSZE9igPTYqOgp+oNUFRKKopJrTgCBRUINFli9Cj1y
rvl+XPb5tXkhbYznyBRLPYL8Qv67CWRmQlKxhYCv1CcfSlKSGNXuRudsYLK9pqc1
qj8RvoD1N4Fr52JFhTk71QuEROZuT/TRjLxBXleq9nq+Rrcs1LFNvbw9RtxLHI8U
jEV8Axgv9ph3rNTrlndaVpqXiqMDJCNKjsSDHD7CQ0TJPoNNL8nHGMd1/0erhXmh
/z9ExuQJ/BGfXHc9qpsCeHHmCC1glgJQUYK5yhmIZgYBoKW9+2PgCYKSlE/l3gkc
td/ZPgjO3vMBW19nZKeeokGr96e5Yixs/cacEAFzspxMvFrZopsG8TrzYGqy6sXk
XRp4Uh/mW0Ik28IZfO5GhclrZ5wLdy5Fufd1n0c8k6F+q0dONqCCyYGsXLwmwBHu
xhNYBKQTJdA/aLHW6FKKd/2dkOzFSMgIwUD6V8j0LpLr0TlCwHqQla1Q0Wt1yveX
VXCHLFqrYuZJGz0xOU+xtTAkY1cTCYOd2pM6bvEdR6wiLuKhIomlz1bo8jpTzu/z
lqyFd5R0kqRpvk9Cp9XdE7OG7ouhG1dwx0Se/Pdmf7en9Y9Rgeq4J8tReF391LPo
c/JtFWNUPxwxTcJf1Wg/08LiJrXqABYhJp84W2obsBXyz/nVMn4Un6mX3zIFQReh
p49NpGBbQ/8r4F+bZtpcfeBL0deZHyy9ZdwUkn7BpGW6C4flbn6uXDkpD8vv4ZGl
AuibHIoqf2+cwxi9Ub02mNSEQh82K4HQ65RTKKI0gtAGYKsIKKtcJsWsG0pcCwLZ
6watSUFmBBS8NvL8oWF+rIycoI1cRc2CEM5tU98LtmakkBnhHFsFWWVFhAbmFCAe
cF8S1wc6K0+ji1IJjNx2pcTYb8bKO353ea5zfbT8XLk846GTpMCpJCxRnhM6Aq/q
3a1uVryZlKEPcFPrCaeqda18aUPo83juIwzf/bE8qEO9vR7x7g2ic70nOY4G49NW
Dah+89r1/qY70tU4Ok9yQhP7eXw0emY8HXGr+LqyGf0wERt3EU/nWYwCbppSK6vE
2CQgfHcrJyx78WJHoCjk01hpyNKARuJeN8ibg86SOHMZh4h+lCla1L0fHcgUw7Z8
p0DGlXy3ysQHyfnuBFP9HuCxGSh4FOdOkHci1gFfjq97NAVad5KW6eeJqO6nkgE5
QbnqTKL4KwduM1WGsykXECdQzEszjvhtecK7EssKm1BBtPcJbm+55JrhP0SY7cv+
gD3n7TECuXA39pI+Fk568T4Dowt+G1jIuiGAV9l5zPHrFtVhA/w7eC5Yv5oCsYb1
i9MY8xmcO3xeqV08+9wa5KN35Bslxn+yxEqBT6RnhvV5dBJEFydTpa583qE30YD6
5RziDKUAkt0y0PVRD/XZSPJw29AdTVn1aQD0k8xmMdx7qhN3DMOmqCNE8TmkHZOI
Z3F3KMP7uYP9DUf5CQjUEOtwbzttJwfl4Bnd3PGKLEU3tBapdy4zPMhfoE00vtGF
E1EQhAiI3gkNNiePxt3DRo5xlVQHMzrcN52vlRhIZen6SZM5YKJnV9wPsTnQ2Tkk
Ywxyt626OPtbeJ6AkdydF/Dm3BaGwO52fXT3I+UEoVSI0ULodHd0x2EsyjDlxCI+
KwrLfjia9eG2HYxeMD6r6EFTyXu8Ly7pWdyRIsG8fV6aTRxI0kAntfXIQaBRm2/g
EDMEB0NgGFN9hokvVZ09fxe/cYn2FfsNTpL+krVJTLUNdVFlnfxmlfgbQ/fFMQ4I
v314O7cCaj9PiOsDkIdkQoHik03wbsWwxECWtAWZAn1WyFl2TGEuHvynB+Rp/Xiy
zUa1CyWxVmdgWA01XgbRkLwGmSE/sqhLovEfatvk07CkTjnasyBdfNNNj6hswlJp
JUU58oCe5NI7V4LC5fbwyopA6bJbUEvjQhX4NpA+fyLt8cs/Bq3K89wId7+HbhlT
GORJnqvozqL0AEhBi2/986bMM2MQjKxS8gKpkMMkmwt+3WK3tWvE7RKVfqy4Tn0l
KllxpBfgDSRMsp1jfygtNGHCp9Yqw7K+KAeonoHPBkyzvrJ7LnrUC2hNCIB7MtPw
BXfi84Kj25ksSMjcBuKeQaEy/jQLQbtY5plDmQR086plB6VFDnuEIaRkiZRz2amR
Z92PN+ay7xUw+hZeg/IqKjGMz1DVen+994VN5SSDjfUrTChFAFGPAayd5bAhN2cn
5AQcqG83rvawBoJXVu/m1hYn7MWrz4Q+TSx2Tfgiy28HqHmKm1QNTKAPFA2rtmll
CgJeulnqiMOwWACdhqktUtrX1gP7TRrKVbdOLMJ9WZmIJZvJ83/QDh49Gl0MoOIa
qrN5by6zuLUEIUxZMrs5RMfzr/Z+Y5LtETkozExNpYr4tAjCbroZUvXaECWonIKp
DiPX/CygCv4esesxMXQFH+X6FtgAZ5K9USrPMThIrRg6VYSYFS5ZfWkyLjolKnhf
M/Wkgpz4nWrOmHQMcqHXTgCOB0u5K6isbHmQpH0ajsHhE7FtXuj8b7YAkdBu98rl
30kH/BZvGQKezpVMm0Am5T3liCWsYOvGqUphiJK3Q/0j/wpjVWyhtvX+otQ+TKY7
SkLO4UM6eD+V9RZtazAM8thPhmVu6hnFowPTYa6ol0IV/TrFplE0tr8iVJf7wbme
tYYIjFXiIm+wFi3mfNCk5UTs71gAeF9pq7qq0o5vZJKuPD9wgEKJZgp/3S8D560B
6e2SHnmerzJZwC8GVgkBIEneZr5o/RoTZtatYgUuidOI5KxyxclilFS7X48o/lVt
SJ0ioZuRRFAjn47ai0focZNof3+eGZCgSSK3hm0FRIQs0Nrx22g1n1zgiIKtdIwp
2nBWmfG9hk0tOKHKJDpqbiFPeRP/z8leTDVlfYvRDLqFq6FC6SnRVoRWHoutkPgI
KfWAGt5uzf8fLNcPkXdb4bR6Hfu0Ss7vuBZI12UHykMhl7j/zyl4t03sHKg0M5wW
Ptv+H2X6MmC8daVi1GzU3dz2GN7B2pQWne/CNBVLPYgcT8iktbfofh/5boLpXhzI
Y7M1214Fk8Cstc64Sp1kA5EfhT0SRNLOUqcE4diUhNiXl1wrz90eI/77XmOWX0Bu
jitEJfTT2Jp+WHpeasL/A6saCi3yqJRqzs9hElHOrDNxe+89yKDA5h3/qhFX5MiW
q8dbTpI1y7FiJ3QqW60gR7WcibG1j78G5XebSsNpMgkuQn+XDMP5/No4lDx52xN4
Nm3gXhywMm6mGQSg2mAR8imxp63/8lL1cirD/v9Yxx69ZaljrgeQsCGDRv31yTV5
fROcZH3/yqGaHjO8lvPrTWX0dpcn0jQ/0jNfUE2Cn6sH/DXu3HF3j4WRUSTtuDpk
mbCHZ3zbR0rMg1+J+SXUSIaMljvTo9X3WzU+wi5mThElzWJfasPTJzy2FiPkTfLd
eGdCSvFfW4DbLhqUUwDA/OD3ct0EaHADRgEUC1qWqriP+sjObQqXFDVU4vA9LAWD
le8mvkiLuE4/B1UDa8IG6Er0wxYYtg2Z8iSh0JLwZwPCKUhC1ePvbLUYp6ATirf+
4JD4HXh/ABx7DVU4m0oALFPfCh6BS1haQfpmxTM5Hixpa9VvpBOYbgxXy63xjD6R
IRrmttE7hlLjLa1NBeYXyzOo/zssUMlCE7T8lO+zdW3Rz8OuK/Ca8ML/wMa3xTTd
DBQFHzlel3KsQMMBgcxtHcfMjc9BgyKCsnwz1JOXawaNEIQKFMqaheTl5sNSHR57
ypKzRMIbqbOE4Kf2SuCwTF8I8dnX/rnjIRek7lpmkxbxeLUof5jfTpFKUYprEmjt
lzap730HgiVC/CgkmrBYvmxve6tZYdVVKFeldiVQueGn/uned47jvXske2srmw7R
FdMH3UUoHt63QxoYwgbWWdKs9r08o3ityOjNLA7i4W7dBtQ/5Z3eyOW3OBEBugjV
g+SJEkHji+3a1Gn4hCnR0SRJH27qbatMHbXbVYPa8ZHufvilPggj1lamf9DFZrRw
14ABqlPRJh1TywA7BM52Rcpj4EiJ6oBFqO6cY5qFbMqmfpEC2BgMwQWrCjpe+S4G
aKggws1z3Yj+clKrQszqr9nZWzoxN/gOP8ni5RjlLUftQWVppecnABwEifw4dW66
jhfTgXyd3nErl/IbzB54yrSmDUBHxGM5tpUo6W4rwqyhLvbi5rN++1cy5Ec2dcQ5
jSGilX2ovct5/jbIjD1akH2UAw1OlslCJfX/HvhXqiTUVkOo9McPG2XaiphMnNQr
7FTbzjBwq00cQxUCb7lJYvIZPxnIx3CCsyETpY3cvzh+SUhhenRnPitLg7/txU5B
bKY0OwyVhEtv6wEBmEqvIJqlumovW/QnCKRrPklRR1dCb+tCe6Sjfmk6/UgLzgzF
nH837cfwUJUeN7GNmF/2yPvyq3vW4nInp6HfNAquFusvCoyaehWx1pCXSpwn/dOX
RJ9c2u+gIQTEUHIfRFAkayh+H5MOAgZMFu9uWi0VS9pdU7QfndgbaaegOcQoxXQB
580MHhyVGPAm+OTyt1aIWUvQVzAnRl8u/gtNvXSG2g7VBLWPfVNDXWgh4J/GsQZZ
PmLmTTwG8wCffWVZzLnLbL+bCYESxM8CnPy6HsDvSzbbklyPWC8HSrzKu/bmVkq9
YDbwCX2UERaSwDKF4rYGT1bnLNR0vB9hUPuHF7vEOaJ+kGvVG3NKTXz2/ncRFdzo
cq0JZ9yZVPt1fB50+4F2omCb2oXlu9kTXyajfhAreOmRUJ6JVSzIr7/DcLXg/Bu2
MDVVdIvs1YcX6B6U08Iq6pAiK+jHg4JIP4f5VeLr2uKgIpUxo2XXuZ7ltGXeZJFt
awrJ0nT6u2ePJta3g6RgpTfMxHJ9CDGeNrAQxK1z5TA/0VdFium+pub5Ax0/2Ot5
4cmLC02GUYC44+BxvsJixn7OWPvi5FxjOyQ4llB03Nx6let0fq9t78wT0IF1paL5
0JUhs0XJj4kneQ5c8Ju48NvWU8+1t4Sg4nofIfH2hE8dooocoN4rTJiZSFrFM2I3
S3tOvoaMJm0U/spI2GWdAZ4kX/oUFpFbJm/thrZwXoQ1ffAGPwm3ZIZy2cm1U1P6
5B1GtE14fkUjdyHdD43MySLn7mClIzl9WN67lSNPTS3j8EgeYziUKwNggn49G+yQ
bORqHjG7ZfwP+mUG+3gnVZrgC3Sa1hER8+8LKAUYoxTMaHAyfFjJJNKAWzlcYawu
Bco/sQevaJLiE/2BgFrp2Xe19wiMXQn7N/podU2R9HSSbSl6gdsQe+2820I4mPoc
jvBLQEjaGGmUt6zC+KlchrSu1OlxaoVYCnTysMoe84Q7R5qf0lfCPvI9QQrpMb6k
sRbRTQJEkoP+w/LR6xqPrXTooZhvYDZhzeONfCR4lceJ1K39HE96EDuetMVA5nKD
eM3blstVHnOCcABCw5zJvoXrzxcQrAJ85st0fBx0BT6MjEX/mRUPIskbByXJc4wf
OjYI3mEGSyhQAfv+uca1ZsGmHBZUS5sMG1UdliqCwDxPW27wvUuO3bDNA1okwcvM
7m9H8BAjIFRozJPHwnC0L7zDF91ZgSLr6CkMdClePd0b1ELqTHMH8Z6KW3kP8nuU
+Da267FlEkI7R2tWyDyJharR+7XmtOvWNeWmTJ06fV4hAGTmXceZ7c4mvFudHN/J
nB9XJ7lRY2dEsqx2c61pR7baPc5ehfM8+yyrp5+zHVtvG0Ap/thqRCsoNDJR2MT3
48majwtUOt9SyZlDrqdsAqvp988KYrfTt3NRaY5ftmj/s5w+n4u98G2iH0p0h4Bg
NHPh+I4kVKa35O40qT92yk0kvaK/DQXQBHwoCJ/oultNrPmTKjOsdJoOWnyZSoui
srY7bc3JdkbOidGuyGSxCaf5HiIY6Dci+BiC6ClsAwF/e/7KIRTOXnZCf/KfZ6SG
a4QmnchAg5nQHYE1elQuLe80SgLsL116SQPMDpTrAEhusn4HlaxVG6L0m0Piemes
NDp9+oaM6p1XMFEGKJhEPlk+ow6UNqQVTs+HTE9WmiWYV+adTbtmScYwzrATO4gy
pEYcR63ZiRREwNOPpB+oI321mQsNadTNoMCr3+6pHx3LnR9aU3Nh4s7CRkDT4SEt
7znVeV8WWfzVRwHb74s8jWPCmrNQ9H/45ovacBMuwkh8Hen8ZJtgdITIqgMHTv3F
i4oMuS7t9b+lNJh7+RtNif0vXDNS+EG1PddWTv+3uRtaGYKGoaSjj9GdfPrav103
+k3jHCGtd4Kxzwj2eoCraJBXYMB6mLzHjpbgN/e05rbLP7g+PYK0rIMxN2wrBU4Z
RP0GsmzHBsJWerX2sQOToPWK1gj7XlerZcKQJ0KhrRg7dJ7GL5j25a7xcdPaUluo
KIoxfv8CaoSNq92zoZPqBAZxrBB569CPd5G4TtPV+jfTMlg9pase/aN53YUX0BWa
O1ccGtqeVlgCpYbLld/jG4+sqvMBivwmeRR8s2NJ3FxPQYPviPbAKbdVd4q81RSf
fwTDBQLJ1K4BCiaNnuXOpuXPhiwTFiVCLR/rP1EHPzF8ahRUQInbyn7nxNrg/M7z
GB3U2W5v/Tjb+hmAW3sL/GEpnBDyfeTky9qZaob/OT2p516Ty8vPs8b8T1BFkzAn
Va0w1kkTjBHkXm3NAhxqNQJyeYfX41/GbLyl13gKNZxyh5oUXjSeitswKFhqQn8U
ExIchSOv8KqsXLk/yDMl8CLj3BoTKCWuR6u7d3TEveLLFJx3wn9RTPkPHUlSbySL
DpwmKc+S38+e/sL8ICnHSgvYHZMAdZkX9bjauUh7dZSNSVqYMwZvjkcY9bN2svps
z1y9sbbj4sofXcOfb8U3d2PyhtPLmKEf+1TnJmQsGLnXLs6VmhhB+Y16+K9f/LU8
zQFY43wlBQww42xPQI3IN2LaYHr8oBeEXZFRonOKXqZle0U78bKNToZ0H2pl6C9x
Ijr/8psJ9YWTXhb6xJzymFJCex6t8EvaqMlHPN2sKv9y/S8PTiulmzPlgOgZLXVT
k4HSnfhEqcjR3OoTRqR0nt1X5LudlNlfT0WaCY0pBeC8pV9HLY4skAOBYacceZsX
gpML2723aVaJt0DhgjhW+WXxdPY00k1LzTQeYh8Xuqk7MitCqWNm3eDqAVfcEbgP
gENfAg7o+z2PZH7/vfRPbvHRGr2Jw76/VGXHaeVn/dsUQnfzaH2ImxN9EPn4719r
fbgvZvB7V4e9A7mUszQ3trSR1Q+6xCquDRhKyA1/xQlr7NyI42pwIl4OJ0dlCePm
DPVVPaWWzLEt6Mi3QvF9J4musGK9RIuMBU7t6RfMm/qfbm220GytuQ3x0UFqPbXh
A0piWktiV9bATghcVcNlBq9l+GDQIrZk3YWYx02WuNmtYKRysiinwm9ZckhGDfpR
GUPMX5F41W9RgdjnGw8RUA32rzmTdNbu3Zij5Isx8M34CPaWvDPxb/g0V1NKj0zS
DvgvStoDNu+S7o2ti/LFFnIx+bXocTguRwxJYmTtlm5rkKe+t67VVc0d1bZwb9pT
d6Hp3vfVDbMiOGn/mugby4QUnUu9yIgekX/feZ1CNdNzyoQTVmLPkLLlKp9yrje9
SoWTh2ZdOkQnU+AqFYEINTSx4bTblOTNd2agqKZ8PUKsaRlNx1w+edUnJhxzNhwx
sGFj0t5ftpDSwR068Q99kVCaM1vDPno9xPSkbe9ZFOy5huXnIZKw9xn1I04TuJ3H
FuMDHjdBjDXDx7uwEGVcfRoNpoMFXNJ8V6DY1mzgwDdQWSsLi9f0pVYjT+yjNNjz
Fs/cF2D0jlCE1leRTru/URcr3S2vD8XVsA2EAAZu+W7o6BhVv1sGz72TJy6QZuTz
JBWfrFD/Te3myxEIzPlCNFz67t4O+ZbNmAdf6H13pr5vA3xMNBe6/tRwXF9AGEgo
o3SXk1YMXDeVDwkSbFth6Y947IeFE+g3MaIgwLRNNEb2W4Df51MyJywRpmo2XbFk
+A5CxtF7s+JLzhlFJ+f9h5So0jdP0w7IIolRML2XTCdGxxtTh9SMY9FQUOvP3QMY
8w6TODQYddmzFvm0QJAiwnjT1928R74bFkm8bEe4a68c2EFswDMhyAERsiEavQpW
tU/7xn2t1b7UtdAqkMELKegYuFbhD+5O2HZ9hAmlo2d9okpr4Nzq3OiWeI3uU3+/
5oQYFRolEjtEP6LnUnGcHSS6qA9x/jroNgAf0p4jtdReokle9isyAM+pX2pnLA/1
xxC9/xgI3OUuZ6J3ajCu34txHYxXZkbtSFNShprz0GOJ+qOdpbpYRsHJSn2vjfJM
H96XoVL152NwGOP6q06LN+M3gyKsS3SWL39cwQ8mUZFy7uqZ8M+kMcp+/KZYDfiB
jeh5KTj097SkCdKk317eY/Pf8EENGjgbRSvH2rnwb/Ws5GGxqS0cLCPw5QWtsEK3
3J0+s9hNRyef3aoy3Q3DFaqwvEuC5Rv0NhXpEF6w+3IIJ8OCZZMgSMwncrM8Ck6R
/vfYLZI96hNKk6FF1eYgzMh1oAlxp4wzRk5hfxU40QgshzXaFwip+M54orEclJM5
qfq1/Ib6MJiRt/fBL0Ggl78FLZBC7YQmY1G5d3DNoou0pDYASRV9A6t4uHFNprmG
IqQr//9B4qNU6ynM4a8STEIR7PSw2oYM9xkIvwtLYoV30ueaRJoMr5qPbBtV1pRH
gGUD05C9PDh9Z7Tzm5cjgAexCDQdebEfm6VxB2ZIGdiXBe4Wx09Y3d2gAKhGGA6m
+l6uUtx4LeHMilzQ4RGfPn7HA3oi99iif/nySajfKlqxs6+PyHROvBGOsg79HAcj
8VR2rpaDRKlj3VaLhQMR24USPnNHOyxiusP8R+JCNB/9TgwLb7cxQtYgtxggzfDx
xZAoULtHsZlmwYpeF46h3q/eig4HuXqW1ML91A8ac/UEpnSpZgNvA0FWTtFgAMvN
bo8d8kpW1zNcYUtHKb3/oSBF/ovqw8QEmFbEAp6acIXPXmXcQu2OnROa37ioP/ro
8Q72wdAP1GoXgJptYc6875e6XdwC5JwqSPdYNgxP1oHQzgOEpd0MIdBAp4AGG1QH
sA68HFGzrqpqnAOdTYrCOpeobegd5PyTCYtEDv/ZA5dKnxUTN3wIAXAL5/wckEMM
SBARpYEXtcGXu97IIYxCSJVgb42UXjjFA0maN+uOLNynsC+xmdFNfzkVxrNJx/nD
S+uyDYvfmQAxvtq5zgP3Gc0ZFqxE6dpzwlxv0P6+zgGErt9BfsYmIP9Ejj6DW9Sg
1fFVWBcCvG+uIouOqVS9g+sow5RrY0UFJd8yu/7Qx1n458Z6X3Of9d6e/anmiIIv
j29eyn0SlkGWcCt3PK1PK295uZIQdbu+K0R4yw4ZWNZEPCKzrWYnGtpWd4HhTv6M
TsDqir4h9OtbIi8SmewwHW8mnJB7mk5jbH6EzhGeYbxJYmn/A7m5BpZtaEhPfTx3
madmrN2dCU707wYQ+cZkv8tgJsZ0X76P5tTaHwoV8qmi+ghRgckEdljLXNAprp0N
ITI4vFiw5410bFSKTzs7l7zM5rnYoUPGZgJ50v1qshYG87MGWu8gzx3ZousEf1CJ
Ay9kvAUFkA4hjUSbR/5E37HlbMY2n+z/tZoC2I0XH8xlEA2n8HmcTrce/gOy5X+s
EjhBG0ZM1i4eZBuDXSyKe7fCh1fNzUI00juKiqQ7FDNpYbRvaTm+J2QJ+mV1N71s
p7GK5BhjY4LEUgldfHFYc5p1PxebVB3ewp8Y8kWrzJmp6Nm83UhSZ4p47EpnE82I
+nlRsJ5KYKAlSfVSoIMflguCCOUyRfQpeZCVmPZAI+p4drmLPMOqO7hXvtsgWxVC
jwNvYGCGR4m123Clo2MbJHpLPcNmjzYXH3vWBhUczcvs7RthdqV9PZ9rwjV5wAu+
3ZJf/kLmSSVpPmdVqaxfgY74sOdxhnwLmWocRRyuDekRwxkHB+ufOB/W1a5jIcVW
XGlcB3dEgV7GZXdMghwLLhk5E+0zNHHbfy+KMcFwiiEQP3bH6QGlbXxtVgKg3KJm
ZkKr/7q5DRDy2TYWEvnbqX+7qt9faxZquY24Ma9AqpeX2aWz9IPytjtVqESGru4A
Y/TodJA1j0c1UhEo9aePmJtyT1bXAoB1WNCdZhj0NsYn7jMmGoZOy5vgR40+ACF7
LOgAP2Z0XoPuYsO5zJV91Pqz/m83ZkCx+mI30jyWJ6min7H9lkt7h6NkF69hKIbS
m4hG+J6grelkiO698CjR0dIShVPbpVdmC/yFFCR30SYTgGlyaxONcTOU3JYah4WX
IGN3qCYpddaFggj/4u7cSCAIBwtMwMOl8m3yX3FTM9HT5xG1tpcVw7Khi4BHJuJf
Zpn3hB94UfHrxzGWXCjKQqMsraAEVjlvqqi83vK6RpaBkIeemWHpHkDM+Kad3T41
d7GV/YyUH2FgkZ8wtcdbMKz3yOKE2O0R+xe8kRcJB8ws0T9y9KvrZCluLj3ShR/B
A+WVZQdCYovwqDIUegMWORzAa8pxxKbsIMo+Rm+rYYWNicy0gtIFV9i2RgYhM47E
2tO0CbymZC5vijUy07/gfITCpjojOKvVwhN3tJE3gdmXlfBV2PlxDm/lLwsDYp4S
Y9Yhnj92N35997YT5wQznPppxJebRY0dn2shNIKiMs+BQUNNEFDCOzy7hLNcLvbZ
wO3/SSAeEy5jHeuKkxUnIacJHlQzAQflqY8qZugh/iiIAKfRXWinQf4RZxUw/Idg
fE7XEsHpL/uys7Bpy2WriqvLU8Ny8eoYiMulF0yN2r8FObINt0cICkExTqOsoBdf
MHnFzdXMTULQ2Vrzcu1OBOae6zdu7W6EqL2tRBIalfB0VGTbU5sm/y7o0QGvl7to
REl0zjs13JVFPaXzrz+tqo+hP1AOPvA1FeN8aL5C575h+FTCI0z6yVe8tprM25d/
F4dBDNaJGFdYUf16DB8tEKAZGDoBYlfNKbwHYJ/9+WU78nSnkca/qrkFIN22YO/d
35Ov0alYm2MhYHVKnK19g99B1xMp6RM3XNk9C/eLd6+mnGyDuS979ly3HLnXr7oT
n7ypVMQBm349tngHIc2aaJQtdQt4l5hg1PK1nKkX2DOI40w/QNh+5l0pw9DMu3FI
Gp0gO35KvyYgqRfuI3rz6YVp9IE6au77kd9rmpaNqF1sSTCZtCPpLrgGitWRFEEc
LweNSK3p6x/CcvlQsmcbQLRHT0XjxIARKOUsz82gCA+2FFz/SdMrjrBhzCIwbhWz
Wovbf3R8gDPUKGw55aaQLUT/F2RSAMIe/jWSeKeQZt7QJgIJPNi+wbVCAwZK6aJ9
CDdyMrwWQ8NxKfZCMvXYa/o1lWhDqu13MyFXNE9gyXlRbncSUXi8SnvhV++kk9bs
YOLoOeOPesWFI4hbMw7RH2HOic3F0XckIn2r6zy8LO959f3Kg+Wtj2tByzrNM7gc
b7qfvBz7q/OFPnI3CvOVB2DL6Epp++42Uij0Brw5fns8CyskgZE1+OJgkfEI5UZ+
6JPchTCDcPYTFQuvCmcnX7Nf3J9dSFr8UxcgblZFUUtsWSiB1DFEZtBEznZE7XhI
D+o66mVTdaifhEemPmaG/cBbls5dU9YLz47DDTmksytLRq3+Ilzt0+KtageuxueS
BYoPMQFO998t7F8rk3AnjjLYLyi/QqYckfz8Xea9FQxxfFOqP3FBYDjlzVH19s0H
GJ3TjQ5JV4NuGeXlT1pToziACgTJl/iIA+b17EbDRIImC5UuMkYvuUIzhDjHamI3
9EoJ+qXfmtJeNgI1nUduVZV3l8K9xFrASgNL3f/9HEyEzzH1T80/xnaRWzcgAFAF
93wUEEylh1FBaYO/9LW1LyhIkWGnC3WQcfnIyrpRl7CthUljt79S7fZXkn0FIT+K
uIhFwxMdZaq7JHSkgRDgNVP4FvmMI3mP9mhSYzmLYVeZ2DB9e3QQP0OWwflhRo+g
4xgR9/kiH0+YutrtEh8PRw7jo8JRQ0puqNCpzWztmXBjArlXY2+NrPorAXMygWNZ
yBi1vNnT8b/ZrnwcNeNYdHpeM8Ru1XfNKXYKffHwvYAqaE5cbBEpQw9j65yteEK/
F86VURY8PFeaYq8gjJL6MlkiKsWcpgsCNbQhJ9l9NKgzniWUlPnl5nLdr5659KF8
7nNxtoIE1H4E+etJ3I7GKyQewlBuUQgSF4BFtyqZ9u+ucgmAd/QCdSlT4BYW3H2V
imyM9EH6hTF26U/rgQxZIHHyPgmAC7rolgeSV6wrtBPqBlQIau09z6ts5b+RSuZw
IGlP6ZIiwEV1wZ7dA2e2y7MyH9s6daFbk07QpqixhUFvey3yLaX+AsUrHEYvGU0C
N3MFiE/qLFTBjFeEjsfQGQt54/2W+bkrp8TCM1uN39u/SAWnFa/E6Kzfkr6o8FxG
G2nkZKvLIN+4PBo1v0MUpOIVOOpIWFbZ7YdYZYWjvWIA7qewvY3ZGQR81FInQgGr
oPkn37Agy2lBgCuSrTLdplP4rQCGHpV3bTWsLmABdsIbqul5bVsHfnHk+pfqxvKc
rGGsJBqGJ8y5XvXRvPGpVZ31qVbjGD91rI4vjQvUsYBpUJtfHapi0S4v24FgbCAJ
aHUeauhL8W+7ys7xaBt+OSU12eW1aXBOuonid0rCTKY6RD4zoVUQA3bAzVBZYVUB
wzaDqViXr2MyjZ07QDWN4pLeZn1u5n2lFOOpvEakib/qWwYL1tshVmkhiQFv7lmj
m9Xi6fJtrp5qf0Nnp5GqmxsrJNNCLJ4ueBjo6ZzqnEQu20q0D7UAVxVpT3zMOJ9v
PrSoge2kYM6davLl8KXoam4lejqLhJSq20qtcmOWKf81WTcZTH1JMWRovuROf+Im
UbYTkcbLUe2SWFrYf9epkiWFx5F+5+9K6zhoRQxIw13LN5KlE8jSxivp7mMp6YGZ
szbHHx6b+G9962/I5AWQLd+KhyT4BSpmvEXNutlZrEhvU3eCR4hulkaJY+UaMEnH
VFps8o7wsnhoO1YjT0A0Vv6SwETOtoKnxQ4VorXLpqvGIxxRT1GhjO17I6u/3Kr3
mysMcDUSoBxyNpAyIFIoMS3dbAbfx70XdbjBOQgTnhs4Z6bajIeo385g8+8v3ISh
9e6IHFzcFkLn7GVww/5xXS2ZBJL+HBptU/iQTv/y951p10juNIifYyTD1c9VaYZU
P/VDBjxDeFfohJMYijJRW3E7Prscws0385uWoAnf4yBZJZOZxC/wEsUDzmlSgojM
+hWBIJ55ZWlh1VAquHvpP4M0r0IL2meG3GG0RFrPLu2Lv3wdH1saGjyPI9ZjciCN
RFzZXefiuZjexjXpLIDDdOG+VKaIUaToZylP+Ts5h/Q3tHPiF793qb3S1b9kIox0
gvL1iyPfeg0JzW1DjRqJQ7U3bqhZo3gxaaoOFuQN1CNwoEyjLFCA+KIyG1RBRc2f
x/EZxt56R/DkfhSDaZ7GWUaaB7E80N1YVRphTUU3WiL719NZpJ4UmqviMznIsL+D
Rh76xDSB65O38zFGu9f3GvriG3TvdlIdRzsUNUacp8OoXhWv9YpSyUkrBAEbvzCm
nIwaxF5e/ATey/k3yEBqKHJdRhZ2OFR5R0QmkYFx5f823QpuRmNzGNSQyOf/5xy4
dnrgkDIna1GSh4CROK+MGp7C6rEK+pio4pIEFi0laZsVLppcvMsTxpmSKKjZTLYI
j9i7ICuNURjJj/xt6U5mtuSqA7nu7yX3BlyTqwkLB3gH/M1uRDHJ//gJ1xTTS2u1
i6kvMmbRBO2uK92EJgxqafiixCja8oRJPi3q3SDnVHwOXf7bSjppWPHtw4LlRuKb
ZtbDhQjdy5X4Hbnqs8nkn1MWM+LRaaNCjZ2EdzxLdBMaMyNvt8wWbURmIgiXhg7/
UXVFXqNmUbnzR9cwLt/rSFZoOP4fcVoszUokFLJXLhbgmct5yKpPVPiYvJVrYJIp
kC2ePPP333Mve9ntjS9VTY2dqAstXDLvD6pt1w0GjBCL7GOiIwcuzTlP+MRw2Uoc
SEsHhKFb+aRJc7R/I1YRb0lvXG50DqZCj5a1PMlkVDsxTrOGjRGdGOErfr8b9MaN
7KGghvm4Rtkm1PLiUVeirh+obDjnQLpRHFXk9Eh7oKqcpX/rtBCQf19Rv7C5Y6Uz
J7gvcR6LUKdG1eTNubb5kDtWKwet+ZVhne/KZiUpCeaI+S1P3u6CkVNDl/5xUjbM
tPj5KsVE/ALiaiF+L1HTHwV0EiF0GIiYAQjz+LevbmtopUruGMk/4ajafvsTmvCv
xprVODE2gJH/ZJaOlt8yab2ThAzV7VuBLtW9imhPBSCalCTd8h3vyM+qS5H0sPX5
DhM1P8GQp4h22nqdv+sfKhrKuKC3AfNSq6YglGCJtP5wsY7X4WaoXr/LhQZvEOlq
BFd0qF8/WxzUezXAwDz2B49C0m/VteW0o5Ig5xBie06Wtfc6CtUDlepW6ZQQSlKU
W8u/5HxXZx2kapgpHrwODrI0Iab4NKXrpMU/hqiIhn9y2vmSuiLE2vQQ9GuR+Snd
4S2ohgw2r0rl9y5wW7EekyZ4X2Nf8vfmR536FzxDnD+CufPNqJP2OspLDNoa9fuG
iMyhFEP1iK9/d4NgV/et6EPwHNL6NwWOaVwLvU58YRT+2GFqhhxd2Sl3hLwJ60iN
dUojpyApxJVjW7nzYqducE5Nq3HJ1BBWVn8oK3hVx0z7XBqVk2+vBJqU9ZO4eH+5
8SG60q0+B5Em+Pyv30gxtiUSjC4EHn22cFg2M8844mp0c9GxZz/bNRaWs7wuN8Wk
tJ9V21vdzGcB7tNuRx4M2HMha9z+hEMk0znD8d0poZ6RVfu9ODIp6bXQ8Z3FTtZN
O3oFrHidVF3W+EiXG//rLI73vp1ez8bL/01vLI00kEeL2NQUQPJRjytaQLbAqBeF
5yvVz1lCQJ744cOpjeMM10F+AajeTSCcIuHNgZLhUCuRQIqwmhNsdfTSnh21HpIn
cpRQ4NetKeRJdu/eK52eG/dvQ5LVyiHfxftUxH59pOmX0gyAsuAJcGC4UKu250ZB
qSfaKd29iuibE+ahnEYhQInVxcQY+CALE2hT2DNGu86JD22wwXLlZF/lIoI4HvNK
4KBo7fAUEadHXOw0cSiCHcgg1dbUklB5g8SZrPNlHF1bcgKnMmcvcdlBZoWV40al
UqDn12NBVaqMNGfeQULqLUTebIdB9ylxSSSkJ4tJV503APG2Wx5yZEF9zC5CT/zQ
Ix6wzGl2y5+3PHF4/ulxDvGj6iB2VNah8sH60/ATAPx84/Wdw8Vlt4Yhbh0L+5zB
HmFrvivRsjzmgNlI3VI/JL+lNaYJ7gLIi4QOZr0TjacrVf9Z+pWE/pwBJnXYDJb9
7xR9sNSImNXMvhEZwWSqKbHxICiTXdf80e4uNBnfAssah6Ge6dOK3E3yb29jFPiA
pOkkFNVcJ5+rShHQs7YerUEE3cv+eDfUHs8ZL0H2leBG0XCwUkVpR+8IQAjC3aA+
yzkeNbMtQbW04ebqBa/PxMKKfXNjU1tnDrZa7seYOB3O3x+QdVVKNqu7jwadvJ98
UCh4C1q9hKL9ir+e1WyiVgwYdVR4eMO1Ay6OBu/tgvFBlYC34EUGmnBY9GmLTTwP
HJWcrYCUNRgpZJjDfm1NiXCQjhVZ8RAHM0hlrYWGhRgmO4pwnPzfeLX0+m5DVD+n
4JV0/kyG3dk+6zFr1Yqn62cr4bEmNcVCjYfck23YtI9B4tEh1s7KW7cgAW3vfbGV
yATgcTN5WwhS82S+y8tN3+jpLiLd8ibLyQ6cbAl8MHStm7VxKgRbvFAKeGIsKe8r
uAztOJQ0F87GkTfXGSnB2I9RXvCn9zELO0EcPTP9k0PQUlIJ1BBB+xCea+SjlaXc
qjCfksVDpl1Dp512rirmid2k03CdHWkj7r5fsw2CViUI/buvPFxCOZKlN86RANhT
CAq/PxKQs+VzvPICeq73pxekTdFNqKKVY1dCOJHQ03utwbpttNe2Hw8rX+BWTdmv
azPJyoGOy0NlFecuFfM6YCM2waHQQTpINECr68zbA8j+Pfl7wUM/w/JNkqDgHwsr
jIUx6AEMafvvTrbARXQNCWTgkLIqgEn7XEYkZhsHwUfPg5ZCpp0KMwNwOwpmExxP
HzJjBFQiccwEmVZlz4YEMtyKG/jW5RYkK/PKqBqjPbbXpAplAxMLyBcOKm9FqjfF
W323LRVG+uIov+jA5ooCDTJuS1f33qma+IC3u47/TH8wPRgR7BiJAtnJU0CWZlCU
Id/xfzmwLlQGlsJ1gqGiObHL2WSuZyKi0ovqLNlqJ9Oac2bfzkv0Vf+R7j8j8gDZ
jzl8Z/u57ficGCQ1WHuFoVqZsekPEKrfKc28RCin5RAAhJkqPCETCzuE8ji7azwd
gs6Exk6q4J7EB0t+D7rjEX4/mKEgCe5l2t5DFGQl2kUfQVEnJs0O2GqkkJ5wIzvm
RYk50C9n0sQY09deE+uZ8J2qmfxqHdb4MxSH+rAZ4fsm1EGDRL3iv1JdZFIvk5Iz
WCybC8hFz1N4wvaV/xQIgfiTb1zv3HFZTnblzfS53wSmLGlsGXvi6XQv2T4EbpX3
/AFhHPsdlX4avSiy2YODC4KPwOX97HeSnKamQ1WSaN+l1M+L9ArUxhuI2SP84hjB
14e2RWn8yWP2+Lyq98f0fn/T8F7C0EWOBp3dP1s7DYeRO6PyNwM+HOs8AzRVeyGE
UT2i14mJshJIIA+FB/2ZcvkxQTSAPkGr2qT9gF9CBb29VfZJM03nW3/gTlkqXd1N
oK1dubnv1RJWbTqeSNHOuPK4BpfMYQnkDZVL3U8mEkRk3ndqm1s3ZupzjmccbHKt
Z3rWWgYpSwI8OWNtA8eZsSXjRR6tUJbF+WAO8pxbwFfEOVdrfjZPC/mhywRbvjUt
PWlMNt5vp2qb55c8zBLFCaEoUvwkKzUJydx4nhNj5m5EYc8P60fhcnvjdJE7Rb/4
DlBluds0ormob7F2n+kw9jnb3rWBpcX//j3Hst+9xQUWQl/IeJzuQ6jilGgy92qF
SNxFkBFFWyRnPYk/A5Xy0zhHYZ7+WbMRPYKaiyN0FSrTLpmdzhpo+xmhHr/GUuij
9nDypZj3RhPLmJs2cNCqnpcHI/ocxo/ZrPluKlGvxArRr+gLFGg5i/Z1E6cbYRp/
86+DikcmFenDq/gSc7iRqU54Kd2mMsnnRoP66DoABkVok95SoEIOEpMQ+5ExzqfY
zV9Mje+ov/mkmbH3mATfPjkSLWb9FFno0uKgG50ciJHnf41mUvqN6Itds1iVbenB
Vz9fsg7KK8Gx8vJj3+xpQxQQVTif3xCZUdqYm7d1zG8z/eB7uHvxSD78kKKssYXM
13SBiPot+zJwjP9cWB+Q0RC1vN8kkhPzv7RbJ8m8Q9woED/VxGn8Sdn0gaKo2BqJ
Y/6pBZ4ukTO7FhIWVKhYjeTJ3MX/z6egXqKa93cit+JS45fTkYQU0Zcz23coZoNr
QzuEvIcDFZ79FgvpGyOXOEnUNKKnLUh1TQLJOhFGteWIjiIz9lm/P2jGz0/C9ytA
pY9C0joXMMX9O0Oe6HKnFW9UxAhMn4l1f8Xy7zsHlE1CRK4gH15ykY050VhqDsrD
wzWnc9Zu8S31np9tyXRmcwyzOZaQdIxhtddLqOuI+ZSO/JXJqknHjVLgjIjhWIeD
sD9DkDf+OH5vRg0ISgZeRhtnTknDb63BKF0heks5epT8KELB5KFeNHfu8VoZsw0x
uHQkPQevw4uCoQav/CRsvMNpgzp4rJGePs3cSFkdCPtxGdQaUgpE24FLW6q+1f7n
m2kHKshuEMCY1RBZ7pSzXmf5yZORiYnookhDdcc2il0Bm9ElN0/UEoDGJQdk3vdl
xac4EONRGpH2+UTG2ugb8Y4UlXFh3xA1cGa8bwoGD/Xwrukh9VuMCHK46kIk907Z
ZIlheD1E5BnSAjnBxuSmMDHOQxgW7n5PJhfH/FRUi0zaJT6QEshcDHLbm1y4i3bE
+s80u4E0gzwZM8GiXMQbizOcguDN+WI4wYxqZYmGYd2DeiifibNVXqtBMHJD4gmY
0HfL/HcI1weEROJQBfAIfU9DblxiUYt8MynoNluyieJ12BYzky40MWa4otC0Zx1d
L4wZ1x5xHu2rUkVjq8GnApGfPOyJ8zFU9lOiFThmdiQR/diVcOZCbCt33xkrPbiu
HwnOcrI4QIF6RtmwdSaiiMgE/xNKchIp5Z++WEclcc/jyQAZiG5GuGw4p7AJNQ3e
h77aFPo4xfBXl/n6BP9rtpKqoju1/42JoVWHXE2kHm8/LzK8fBHPVG7vk0RXEUpK
X5YDPoPqezFkwkCTO6BpGy/13oZTxUxU+k6TaiLTaLJl4jJHWoS0m3KBgpDqYAG1
Cv5zpdDN3VYBviogI4CVF/+aqHSBkJWz1OCAzERqtag764c/kjKBxl9iyaycsz3S
ovBhEF2RbZ88ojTeG03hairb4TnbCqfSjtXrEDPkXVpss5BcnJPrjBjUxT+okBb4
R5XZfbRNIt7f87lDpaQG2u+9C5VbwRaSiWJe/ViyVNTipTvrMLDjvE+NIU4OP7qC
skYSvnb/EETWfY1W+U8hHLGWIh6r1Nt4X0aQERK0Qb36T2vS5BBmWueYrVTxf+HJ
Gjyo8d3iJdKIn6i/LPYkO5vHjHuv6OS+bFDx2z5YmcAUT7/jnmexhcqeTviUzsqO
KsfO8NUutQWR38gNBeNMbMCp/2fxhRqnHV6zz4MSyIuYv45b1ncymyABM8AbuLoq
jSn54lybj0tYw5y7JWkZandFGTBObXaICDzWZYiG15OBEMOYJBPaQh0sGpbAgNqT
Svj86xlgZBVnhw589M28Cmjcg5auHUx3SOhcCwwlIgiVqE7nd/+E27S7x4VPcpdc
Rp1WGTY5pmlRPeDH6qSZhqKM4tIqbIUeoSLlblpPGoHdJmuoyQkV25SADpyVgaOt
3i2vmZh0ZVrhAxGDOgfc0Vjss9+j7v5LIgadLGr5gym41j9Qk3tSmbuWf4sFtwQz
2vGu10Kju0GGkSX9o5Qfmz4EXVsXztk3ba3NSr5U7x+bxU8o/IcIF/OnbmdzjpFq
5yNVXx8zc23haVMa45f3s7Oeo9eJ6koNfxQm9gpy/mRC3R1pvXyMQbVuiF5yfg1D
E7xDdSI7MpboIs9d6Wx3MzpwPubWg+Kggp5SAU+6XKXvGu31mtSOmoEHt9rRFu9k
JrWD4vLa1wrbxsx0nSPXe/IRTsSnHG25aaTHldwe2I8uWSgO9G6EUFC1q89n0vTT
EdhhJPI+3P4Fh6ctHhxB+MmgieCI4A4BYqz2ncvm44B6WqpZLXpoooMhqn7E8eWk
pMXzTWkE+SmxL9lY9uQDhHtB3SDappDPryUenHZlKpGv48VaPw2Blmp4W6SMDppn
s5gKmvQUvx9vZOVUxHnJF1nm7ahD081QNp1CZMoKac8JBbYoB7VDCefLkGE6rh/i
tek6GUEw2CXHn73GmmbkflpAxKDyYbpSBvUg3Y03Nc4GdoCnrmteB4jk6Ixl2BFx
I98ffyJ2tqkEEZiKEH9BbXLk42KWlo8qsTxpLUjCNh74GHUaa7s4S7oc+nGZDJ62
NEdNzkglM5grQV5SNtIdqEmYEdDMbm/F2r1bCS5iIDu3zzFPPB7R7NDMytiLgLKC
MM3zjiolmAR3yFJqW9oPm8V3UjamnFXbISK9dDiYVl8/99KrTQGggTyng9PruliT
XRcOTu8IdNtwbvg2v57un+CiVud6AJ77fDWIsH/rJrPDFm/Ef4i0i7m+MaOjFcUR
XyMISUQ51zZbyk877mrKy1D2dkDqb5dkEPXdUmSJXOmgag7KvU3yHDlFrJ6XcyLd
5TszWK0EsfmYTDsp5jUxE52Qhi6Pb2xZdmuJDB+Xu6BuchO6mDszPVKlmEt1PUXW
PzFyDMZ2Jr4oBYUp0t9sHFKXzhkoPX6ix2jyoRizOG+bYK5DbunowaLmOrMgmvNi
ernnuRVTaIidiOto+nF8lDee8H1sb411Kdz3HPmGWv/auk8iHsfCTAgZW9jYdylK
1O9TAzLBDJDhKPdRUMo5gnlA89tY97Ztv9600p9DM/K3cxNCvaOocpXd5WywFL64
f98Da07Zq7Y/Gh9VU4B9p5lV0IG+v4z+OzIGzPQXYVOwo0aikIGu9KVRFFmj107+
GjBcpolb8tr2GOqHGnrM2WJOraaJXwjhc1iX32eV9CDBd1xkR3Sw6WgybwRebBdG
ngXKnLIrxgqbQN1SmwHYwLQPj/giSp0og9XK24r3OlPQABysI24bSnfaKEDgseKt
3rIeLXRNbewbIaqxsA+Qv5Ng3Jf4eP+64CneFs1BQgNKZJTAwQSsJb0S3diPCB1E
Qvfs5e9WwS0h/XF9C3vgYmrXy5kXWQ3A+Xa6kBXa+ACcW9T1xtzdh6Y8QqnK3NMh
ZaPNvJGtVdp3I482/XkcqqK5qrnrsiTao7ip0Aey2TZspoEXdE457U2Oe1CLnrhS
VPse92406qlaF7xz9m+6JJD1KJ2AbdBN3Ojd9gyge1BCitrHvJZVaELpbzM+9tvj
SelwHXD1HayLjbivIMf0YmniPFNJ+Qq3uht4BH5NwnY380HYE0yTh/suFBzs4TWa
4hwMVTzTB82IbPoQSPo3EUS3zAxIQXWgFLedkMslrHyyhV0iRpIhSlEzRIMnZZLf
9GzrLf+PzasGqfmD9/yirqSNEvngqhdFhgMJsOZ/ESPuvh1U5qdsmHaPpEp0EADE
3rYeKcCci7+cYvnIT1ENbfKI41HON99iQs11orWZvtp7XIMzzJkwi5tROY3sISer
cuyD2ExzqNzo2I74RUPZdYF2HU9B0DY5AFbmRWm+bFupqtho2RHGsYPKCDa0Q+ZZ
uBxqTwaUH1TC3kHoVJiGM7cNKakIiutyctFo+ZbQcVQYZXz0ftckNyyPd+Q7mq6n
Ikc9zuu58awV4Jrs6P58tYu03BD+Kmvj4/Y0HRSX9HFjvdeEwLZAp9/A+2oP4NxG
VIJtOW14mKcgVnSbptttKqNXcvvxt6N/xTQV05tFwv9bNs6n/ESwVPDdV3gzSz/p
YWaLJ3TN80I1HHTXzHT6mmbBa5r4O/nidmUGaobi0LCxPAry8i1s6hpe7QaF4Ef+
C3GkviDt8vilZeKtegxQnAPn3bFWOFawXe9zz0wEU4vag+GdC7Y1ODIY9YUQ+ZT9
vUbTyzVF9xyHWkXLP2iSEZUmsv55xJM+RWhOnOhrpLsr9WXobfurkWJ4ah72Ww9V
CodXGBH8lU+XMB5gGyPEaDg1d0pwcvdyt/wc/8spHwB7jXTxTDn9vN4hA6mkDLhm
0vehTC1IBqoXXF/olJXeennZeGKeCvXSJRNxBYifDugcFKe79R3qKCDjvo4WKveY
6N7r332ONZmYvhDXy3H2g6gHMqCgQixfaCTlhs3AM9aSwO8y/pHpxMFInmUDA00y
gnU/4W30rG6A/+uQXnOKG6gsupETHJVGgwZcz78Qx1h/Q5TCry/wVbVdyrM1bswn
lAtxt4QraI6bowimJMzxsq0VR3qQ45AlYwf2U49x+AOMVQRWGPPsQNsTyb+DARM2
BefO60VUkjF5ra2w2HdUtZf3EXY2O3ZIgFyKfpo4McJB0S+7X1/AFisc78jppEuv
prM8YGHWYRfQo79bRDeAq14iCivLyT+/FtiPavJklmxvBpC8zBvLBqTU9FMhdlz+
4UhTUuaD75niLO9bax34qk03pKnTvszeV1C6tk10p/JyTodzzI6eeWCqWLt3sREP
4OrqnmN84QkGz3B+YXo3Gy5RXlHqhuFPn21gP3lEUonmP5FqU7Qe24OspL+MRvkj
ukeOOoNAmSd3nnzytMz7TzW9XGyJeErS8/ffJpheenQcelsz7GLXTFKzaex+NcoH
/Ar40TN2DNCto7jEu1X5RGvLbJi8kL0zsxkI3bDRwWPWiy2wgLJhB5CSrkglUOmU
dWuOoIrXzP/d6O+K0PYnaVXlRC8b4AQIhm74FltnNWQi1PUSoNgKPVhoUsLzfvqU
caaqeskY1/LuR2GTPLn/YyO9CckCK5h5R/eyYdRCMpW2tjSmEpdbjBi6Y5bD244i
dWFhOWvl89NQaWCGpVVVl4kR6HAnIZX5YPLMRkVUhCafUFKUWmk+QMqzF+gWkBnz
nwrRnYs0DznP1wYOh6RIrosLOmCoLKcSL0XYRtG8wuS8R8bth7OaqXeJhFRx1isi
iiR+058yFhpv0Q6O/PnsL0BlI32XxbZW9lWOI+RNjkyD9Ekk+xzUFWmlf5qioe4D
ZzYwGZuic/j+5E1PLQJ6NUxdbxM+2F0csLQzVMVJhX+KzV4xIU4lwc89yYN8mfSt
fgYKm2dsTWePaKkNsRralmAnEbT8Bjkakrf5GJKuUz2S2cjHAhGDMyFToT0g2hGd
ubkCuFe4Go00REI1UIJo7pPMA7RQuq6uIxhTKOoqUEvH47D58mcIV35kyjt8jYeJ
wuD6bS+NDuKODV7QqJDXtsua1C/KZ1U5FBu4ZNKhNG4Dm9kczTr50KpmFBtC6qbJ
3wpDwKPNHGxlqFAysqoPKwS1J5mxXDblvfjNQHySv45Yx37phk3rGLmbvBx8oKBr
a10hvpOPRy5KIl7+Zied7xxntjHSPZUAfJOOpPOSN2T9pyhyPdyGkIf7hXGeR27N
0EKo8ZBK+OER5J0SyS94ZRGdGLF+yt4mZ3rbuVO70CI7nFBdJiqW++j1zwwsOEpY
u/z36SGMP4XoM2TYUKu+3YR3gRT+Zak4X3tFcdMaD5bHZnPt70fhRHoM0dIixl/y
/Tot0IMzLL/KgSKEPQ3IQTHVDI2NeNg8JsNCW31rTpztgOTQmN1cRZ+Lj1RIj/ue
KrlCYjxwui5iBEJLbVYTIw6CXx7j7ufKQ6jH1wEW1YGZurqv4LWlHYmfQz1jHFM6
bDzGUQOMzUEiPxag1g2ouQse2RO9qroDYut4DiFyq1UPboAPYS/G2lsjDmvdt7R0
K7dAZ+7gU+85jWAmomGsmGhyceN1a5hqLcfcqxapOEcZ7+NVlq8cRUgaBBD/BoT/
ZT19J67w9ehyBzwPZUvixidngyx7ECvUamcC9ERb2S0HCW0/mxJ8HEdQHXRT7wtM
7MMoNDQ3LvLcnB35jrS+yKc9/V62Tdq25/MKy8V56PF3sjt18ELIyneqSMCn/PJw
pN269t7TLUi0n39dmembZ/6XUa93FIMen3NaWJV1TMikVCFXCJAQys0WvoLbk/Pe
IsiAwUqHLAtz93Yr2KgNdwgYk8q2nFs3/ccMG+3sMhixnLKgrOYkEvwn0dB8Ctf0
PCGN2YHqwrRvDY1m8rFqcCE1vZG/e5MKONhCsu0ydsU8LTyVHP+Em2TL5bmwBkUp
8NwNuQUNzucs8IOsQhrB57yEwnpFDPBWvg6E6lQfIPTRA/BAmdA3a5P5fRn1jM8v
tJEtbD25F/JoBUQmDPTNqNA9mulD+O8ywGknil1nk+SIvO7Uvi0/jqnjf25mQv3A
ioBArY1VdPhAV3AQhTeKj/LbPoqiMfnMucGWkW5XuDIpldomrHh5BzOwkm4KF13J
lHkqfcwMyeO2AsLbbJ8CKa5i0E5TA4aJrHUIdEnWy/bfZ2Q8rxyTxiRF0/kFxkyx
ieDvq03dterc8Yj2dMpnXAeQioIriA5g3R6WbMmDL9WiiaYwz/2ZXgbWlLG0+pdd
i2zCQC122doNG/CqK6vUn9nipzCWJPq2vp147GEdd2UggQVbOYfxR6fRbKWqZzdj
1Flkaj7huK8jSybmfTBMOpRckn4JIM8Vt3GlIHvOqBJy0cp096Y6E/rg5s7ioIHS
/Vz9f/yd/ESqa5J+F9Vp/rWw4I3f+19Whc7WDkL/binXAvHiOVVKE/7RZgCW6ANr
ItDTWTCU5I0jQi+nJeqIs+bCQfMg4BoYpxGwIRTylpO/pdhFO/sKL9NXbhFj/x4q
l+RAiPMXnREHWL4jNbzltrbQkBaUUHneDj0erCa4nhEbIhWvdGYeUK45Hy+jioW4
BKLPKYN4hk1iz5HDWb45Gr2naT3V9ZtpdE97pOiF4Xk33ValuGgBmu/Pmz9njsUX
TAfmsFCOpR2WxtgyYQ5Md4tAYXZCjt47L7QKyQyy3yC6Ycrs/kNb71JDDHDzka++
6B1fE82LjbS/O1eI5WLgvzch3rnVavsGLLZmNWg/6A7KSvJlckkjA7mala3Orddp
Ppac3j/FgquclZXphQJagXpdemW06C1IeEgbgGCURSrhFEGoM+0ujUaxUQseZIDK
XboR3D3j8MbSQIxv1i4h4WX073bf5Zh9FgS+7WEnbMfWlSZO+e7PSdeknsaaMeS9
Ux64ULKdUiV+54HgJxx3faw+eshckDM8+hpg6P4P/Gtt/nIGI3Fc3ChvP3JJhIo/
MCsa6IrUQpUk7HW83m33QKvlQMueXcpmTakpyDBzQLDQKlCtcdKqQPBPxxWVokAD
jiz0t8zlqeHTM9vlwd2IaKd4OWO1+ywqkEwm1yAkKPCObRuqpj3kRczRfo/FIffB
wuBSoOkZA51KgZArpd2VtBCscW5wETPyYN0QqopjA9jEAly0zdq9/tDuOu8eHNnx
jLCHTTP80MfriTp7X4UwQwNWQvzMmsZEgcrBBc8HDNTgAu8owoD14TbIMzC/qsP+
K4oR4Z5FQXrTZ68uiPCBAefZaSZMiXY0UfgP3ZLvcpMrTA00VD22US7bK9DItOcV
1CxeS1ymOlCDXZBKQef4uJB/ILNTGGVPQ7a5Lg8zQe3mG5UoJ0qtb/l5HtPWD735
Y7VJvBkWx79gS7ceHVgmtb3ekMVnj3WrY2KkPqtd2peDfIQmOctHkKmO1bt++3ZN
ZaL+oxxKA60+FNXg1495b64J/0FB8KUUBwsfYE4F1B/3a4RxWT9NhX0ZGsfcOVJH
03rctXxd+TXcUty/1bwTecm5juX2O0ulKx4+g5vnMdDqLZHF8H/Tf+6AUQiuN2WZ
sBlPw2cIG3fxGOFFDttnABn+HPfduTjX4Jq5DnKDraokxOt42CRC/HtZ2FWucGwU
90ur+F7AvuwMiLw8L+UK9uvQE+2+qDlBgAdEL5Xwbl+HgLFJxcV6VWyED1K/WBJN
ay1/fDgHiNfucADtqA3Ra/phE5PQM+unPyDniL9cwudL5lvLIE/y3ksv/lsDDzai
O6/+5mPiF/TW6gTX9rH4LQDLaubrzQSr4hBPgZSP7yLqgc1G82QIXsw1ajc3zT5A
p01OjwyPiufBoM9qN5jxcZgY89xNIJ2w9nUGb+gT0N7Ezlh33rIssqFA0Kbe0Snj
mduOw75OnH8yZAYOF+gAFkn3s2D4e8prfdgVitValUYczj5uBLlcP9l7y/cVHbE+
+n0WV3mChSSvYowOCK8vEIQ4sFrqOgVkHSLX0uHHsDu2A2MksrYTD3sGKY4HXM1Y
wjVR4OVNUo5B0Bz6xGaCv3BJIxtiGUFH2Ys5twrPeIZnIgo5uFpm+Jm1HJS2RGx6
AvofLe+9HXRofgHfSMg3lB8DUoDNGXIXLzGlsGuKNbkuF2MmxGvDZaTnbfa5NiR7
5aps1gS96xeJcwsqjUdK5L7hRCWmJhOu1tbpsy3ii+Qjndq1bjjhedZfKG7oyDcX
uIQsPpWFHTfdEKmjgOdCSQlKvX5e3Rz+XoKu6ujwqgrm1Zs/TG0RRTvxoKTGLZrm
MLsRXjsddS7XdMR+EUY4vdHE6HLtgmfegSUPLMhn35qE4z6uuDhppEtig9Myp71b
waAQ5fy6P5i3ahZVmOe09yMkCCehpdVSfGVEBd1YSX3hkBy9KV/PsuPgg4ldvKvk
Dnj6slESli5FwVIZZ+HsDnMtRWg30xMLnhQb33PsgyhSBpfiGRJfzRg6H63u940Y
SmeugK9dB6964hDxVEHlAnt5tBm2/gKJ5Ug04Mj31UFQb45nQBanlmdtTtsmIWM6
vXfWvBCCLGv2IiTfKljc3TwDUkq1uriuytWvP2jtGPQ6MXQSpw2xvRcOUi0DrYiX
eVZoAZ1/56PjBs4wFC0B/Y6WHlJgKAkIWsKZ8vAQbitJY1/T05wQoiRKWtEwzm8j
9Ddg0FdrlNy6l+1CFgpH0E4uyt5P4fjx1xN5svCoPJ0SinL5/EgCiZ4I0BNTvuA8
qR195dZKZHyUD9/6G3TZc3oepFwnP7mYR5eziPnjCwdbWmdR1zeuQ7/4/uU0xDfp
keCtuDCYp84Ypm5ATSygR1tzCTUn5wAUs4Q/UtJ9SXVhzyLpw8bPVVxVNRnzm2qe
9xT1eeicjWh/NTq7SAuGFHSxuLUQq6UVoiIK/8SIYwaNYjtaBE8s2EKuZNa0yxm0
9cg5TcxFtxEdotY/OpXUXJSqFHvzRe1k5jLPm7F+Ykuaux2chHtXtY7evw+dBu2H
t58lB8+9lycBja6bO6+U7Hz4q7C0MSBMrqHilxLdgzay+3TCWg4O+p5NxBDK7cGy
7ul/xr/qCTbq8f6H8zA9VIgchVwWZL0+Fjd/5WOHILaOSSiomPz2MrGbEo1cxvKO
6A6SyryhddbvKWE+XZdmmm69p15Ns2eEcUdd/wNbCgnc2PvBB3K3Vsl+H6FPGl+2
3mem5vczz7rsoA/aDhne6AlXLcs4BJbXMtC8HsavBQJvuvZEj0o7wNwJijEKwMMX
kSuvl3RR5JjLFzjjwvnQR1AO2Vj++BSbidDrpKdw9xdBctXeOpAdKeLRYClHmkYo
v1yPsL/0A0lCclgR3UyQRFA5fRwmciOWCQ+9xOZoov7W9LLmVsanNu66OLc3gqLG
LyIOXCF3MxsuGyMQPWZlXtGWbNAyMu8BcoFEusv3vhNBp1SD55qsLNjYjscGgp3R
R0CY1MTdeVjSwKQQXwt8TF+lGuqRMiHu3cKKddqoLfxuSP51j7QBckKKNtasd2GO
uYWXrk3nh01UR3cDlitSB+S/2tG8a7PjdAOfAAhiTzgcGxYUMEcxpO4jHhu231M3
m4O+50z36c04zvAs7/ScXJJWaU/UyAaTR/M1HQPYQi7l/285Y9hi7fALvxwK1c0k
zZcGrK7sMLkzh4T2hukz9m5BS626gRtlAiYxJ6qAyCJF/cVauMb8KDhEsSf+RZXO
mVp8h6IngjrEGMPEx5xPEhA6Lxg26CedouMaGIjdwOLtUr6kBaSPascawcnUFarK
WQ0nYArHS1fBG3xwueomeyyZyI7PFkQF/zRABbBnnRflWL9vGryXzpmuC3KKODcw
gifWeDm8Rh4sa7Y2NaCTYZiEdMNFHm7m3QnTJsRusA2KxItZhze8PmPeTIT6edqv
jDlwKRR5GnOcC9upLiAMjlYyu+B0nsx5BqtbGXhgYMI+QvEqrgipZ+nc25JEN+hp
lHuGgXtgr8uaT+6NZHzdOrHgeRB5Q9Kd2cyb61Nblz6EYfaAWTAeU1PYSpWj19KH
jV7hQv9b4BbFzRA6irBtWhqG/hzXkyoTimizKvxwvampNG5lCZf7xO2vYacylNa8
opNz4VnNf8c6+bsVWBDAoL123KfT6eJf7JbXXE+tWhRaibbFQo/Z71c5QxyHa6yc
gqgecYcSKUefg5yCNkmytsiZXnMbUMcBZVwCBAKEKAmqkU59njGHcPK7u9EhaTZY
V3MLVT++W7hNiOqmFVcM1xRIdahH8yw20gnmLVJTDV6Un8ghoNzGv8YSDGABDZmv
zV8WuEwJtPaOYtCxTguxYClMhuvz6TH5g36NQkYdVTG8HSp/aP7e2/4ClyJEsCRK
pwELWKZQFZD7r1ZCy2RoXthyso1y7O1gA8pOkDa1EOpWgBLtaFswlSaXDgDRxnEv
i9/wsrvAbQxURSwq5DQ47/0mRcfEkwPTc9Zw/yy1Ua6v4byOZBDpijBLXS53gMyL
Y52rGNpW35M8b1zuClBOfRbyrP4DEVTRgdAPFsrz6DhfUcAhzWTDhxyIrHKEuWsy
5Yn5k6rqPyS9CH2nKCH0OhTvSXCuuiTu9dk6to5QBwStSuikmNXWAlAR6+yQa66W
0hBLHTVyMUlAZWIFPy2uD1KQf8XoDO16DPJYJpDvJySDfD12py/oXtqfkDCr2Me5
aLW/AiwFMpoNz7NMhfxCH5mbDJDOciHqzbVoYAT4YLMBxG1rgX20glCiCKUmEfXo
7j+qtBTmq3o8g8K1UmVgTa17sl4vZrvpc6SVtujG2HvrAVx3VE3qB38JZ+ZbMf1X
ODp6CMP0cgcb8wfn324cKgIjl97dNmZrH3WXlKZa8826O6uWOzCd0jfot9ZekEjz
rpyXmOngA74kVVuhP73w7gkrIS0Kayc4q7XCqL4qLEJZraotkIJGOdzQrTpHxqzo
F2O/25c27TowAp8dkMQJxHmq8RM34DJyNHcyireCeg/+R877rTnnsnfFxl4qU+C/
33Wevo7nSHrFZprpCD8gr4O4QgTWDhoXRI6beI37wL2jxtH9374RRkhbRDnfd9mr
lRDXRUj4jRnswHZAhlr/gnbR8DTlY0hHUV0GfLrKMDLH6lpRBIsV7sgIzFcSS6QS
znOaXVKgeSF8aHL4EQRJ1MXcbsbf2iaHdZiei8vio2wsVfegxQ0PBvgLJiQKZp3C
lVGqQp4XHR/GGNg6CpXpTKBvlmcPHTqDTdkeFuxjYbpR+yoa6R9nhgcgWV9/m6SY
PyMbyqMP9/qIl9RK9a2jLzJyxn9a8rY0WLgn7q+tSLz0jylrwuOpbyzY0XL4vMwd
UZMcBCz+mTq/DeamDFQLPH3qxp2vn5sohNVASyMGn5AKYURX8anGzOWxMEhjyFhe
/2NsiIXaXN9I+05NQbvWKfpbaP9/pbNApVF7bkv0xl+IvaJMomYMesVEpuEWf7EC
Wdd35Dii4Ln+0/XVi7VvoJiCT8yOUVXr3Tzpzp5RhyQaWKxu9Cq2T3He9ytyNg7H
m7ziPKRc6SAC6blirOzBbW1lyK4/5k/CapRD4bE96Il4MSy8lhivcA7AvGc20+Ky
gkSq6VhRdrfj6SY1BfSJ3/CRWzdNxH3G/8wLts2UnF2c2kVeRuLct9LcETrbPgbh
JX4gF4QDs7ppKdLQSdRPR7plzUGL41O1aq2apVMgtaQ6o6vIKhcrIWQa44zYUyu3
jJIhGaiUuM4xN+MDFwgo3l5ZYpsgZXZ3BOxMtk/mJ6gm29RuJk69bvORwgFy24Mu
eXZXLm9IQIG/whAFTwrf0qglI8Dv5zOwvQhzj7LjOb2CFjTcJV5l9Ye/7vfXYrjX
2aChEhjeVcxsGHDECrzmi1+3HiG/Z0o5+m7rgZA+GT4ThXjAbx0sfMTuY+4T076n
y+P3KTdQWVe9yKcz+sv3eZGpzytcTMZdu5WuAKU/2UdOeiBcNYa/sMZDk2wmND66
J7Ji4madgezzLM4KseNshGgRhzcKesxdsiHH49jckIL3qroEXq3xkVQXaBuyqMuj
Whf2JmXwXPFG4yTd3FZvMUu8Y48ijrofwkHi4qPQ2Zx8Q4dYAHQK/aS/H1Ee09Di
pdvKfb3FigDvQxVDrzVS02LTNn6tvXs9/0aB+jr+Xlny+c5/oGx3ZsaxtUxpcLtK
ta2RAKi/0XaZeb24Sm1alKCDARwrh0XMrVNg4SjqSi5JMTa9BIIPEQCVyqFWfr1L
OU5mjMyidZfdy559IzhocZSTYUk3968wn0Z0i9jNOXNld1VbP0+iweTUVrzWVs8z
rMr/NL6LtWxBp6Zxei7MWlYZ2GunXSaM421MzbpyMKeLwySghOQVJE/Z3DYKuIoV
WmHL+Fq658NkkRi676pJlhTDkVTaqDaxfTr/5LgsOYo9kCwG6MHIZkiDPBYvZ2Ye
qZ4asfnrfmvrb1ma1/Vkb7qnfnczuKH8B2scnKeGjd9rg7ZwlQmKBimVwiUKfUul
RDaxu8oqzeGv9TJ7yClbkg7bEqDIu9wDEuBcv+FpaaXLPXzs5EqwnDGINTih47Do
YaaL1IXEF5IV7MAGLtzNRYyggca58Fdc5rzLx256PY7P8fSMcUtb8fCxXYErafZi
P6GkOQPpXCIeqAT0eG62JTuUujGzeP62IpVfN/ACH0Wwo8qYAqkeGknkYha7k7YC
kcaesmJ7T7yBYckWm9XvTE/Rz4Gk1P5I/oNKkm546NNPHumF6/+oVOoStEbHyc7o
5ko74BWwo8uh7jVM1uLXhxU0E9fQzkUNC55WZGyT+36fP7RMbr0/gUpNjDemr6W4
aQN6h0481Lr0qaIWXHegnDzolJdK+65tNptcfWLOacRn1+SSArIGc3F2IMxx+448
2AAJRvPBbmlWaZJYsoidjhDzbdxov9St6mgKmXbRxpHxOE14UDQL3lhmK5vZENkG
eXxXJhnecKtPBdKsKAwqWqrVaR8XnqA8Cn6NwylOcqp/aXRCPSN14Xg6YJtfJYZw
F6Kz7jn3RdHjlL0sgilnO/h/sd0+QdR29YB2zMYuUNbZYI2xrmuCwAuE5SCFlWV8
+qTjHStKvBNq2nlbOgL2zKigXPJVWCCROMLSP88ODX1Y95tS/jYK/rwYYIh9yAg3
ZqERxqX4biFaxMEWQr7SRJEAVBAD/EaSyH4uagdPSVWPEXJZYmg82jbOn8kPAlIr
26f2EgZJoR6MlgGm+7lDqlnWFnQVKkGuZ6JY8sjvoF7KSwG/Q1XC8mQ0a16zS5vJ
vAfbM9HYmTEpV1V2/fGXweBdK1Fzal5ODWFTmIvVeyBvABNUuqnUGH5L/mwUpdMp
8J09xtGRRI6+91XfTFVUNFlCpkfaVD02jWYlVPqOsEFVQm4x6Rc+kBmL7DyuXwZ/
+S+2/0ZufFlipPmf9U0JgCw2n7SQb4qti411Ej4HFV2m+/X9slV59xWCIt4FWF5Q
oH6p3pQHQNePeNq6X4CD0lXpVy5CiQD3XGyvwnsdQaohCXKLlA+iH6dgeZ1oz+By
UZW22GDrIjfTUGiNHa+WpIbu4xKFCfXFQKFL21hQW4Fqs/Tu0OMs6nv7GBqiSuPU
AY3y/DzCMtgVc9bAnP8ddyvRazwvPu8+kIcWUCKde4HA145tkpfddBTFtcnxX/p7
h9mRpuSNr/npe6us58/4g1oQD9CX8DmvyizIcCvGux4C9u8INuMiAewAM+ld4hd0
zxn5obh2A1uwQPKqxnhfl8htTTi0JeHkel6zm7/mS+5NGKFzUs3oEWtM0jtoDgLI
cVqbthGL094bdI9sxgG/1ME5nRfLDhmj8rtx1A14gr8I3cxk5eAhrG5s9flUhkZs
4moeSAefBg2Yw7cWcNE44h4rWXxk0Z9kTJE9vovH3VcmzZqwDxSUj+yqgoD9IRRg
amWwg+eVC99xoWW0rhcST8lfLpjtyrventHUFTbi3HwbAzKQAqvY3L4MBHJeMGkh
Oc4g3pGDZvDT5jTb1uJMJohHQQVMRo2z8gWNipEFMTH04Z6E6UXd7owut5dcTfc1
uHqHI5B5n/PwKHHplX0uKgI4fho0MdCX2zBwuKPvK9N/kvbrxJ5g0oR/zBhTKvKl
w/zk0tNnkLv/Zd2VVhFw6V+C+YyJ5IvDOmJQfXinA8Wp6leB6v0S6V6to1LtDZbI
LPFw+cpSuRn2V75Zz+fC9+RcoaltjV97XmRIPPp5GVlZWJX17Gp5ohEgVeZHtGwd
B6Btc7aqcpGqSi/jvW2cvWF36cy8WejCTuj+Hh/T25qeMpCtN+6gP5j2Hjxz2XHp
L8/CeoN1Qc7n1mlWQbROmoN5p9Lcu4Z3XyXJreIxDhyfPDaZJZsx0YBnPCUnHOno
Wg/q0jWpUnW1+3aMc7ovgi0HgYmBGqDnuDihAWzvy34IKba+FUOAv2D99wlltH81
vKujxd8rnk+K759x7+fwEVNeTSzEaOrEUVFOgEzOm9ovZouSdagSFHFkoQHO3KHe
NduL72RJitqKkLYhq4vCAf30OmwIGuRw9weCVkdHy4d0Em91fYDIogvEzcd0BOUF
dqbHh9k4wnPj7h7ghKVHoptrHiD18LS+SuY8nagwh736CyD/wF6CVFWYnTOmrWMH
GgONvHYFrFCuc5rmqCJJd6DyZntQZkZfbRr0KAYhyCNSORSBHBJ26IHBdM9XFrKQ
p2Ek4iqSWRJ548maXnheqjTE4x1PYgGr/tX7vJpXuKByAybCz0ByCRwxeXLlT89D
hbgId9NtPr7x++MH/jnG+v1MKlc7YpQ9t4SzCRuuti55QsThxnyYb6riB3a4+NsC
CTZ7nd4NchrzXeJoZvFAUGI00YvMf5SUZwaqMG+nO0Bu8BwXTJ+GZTTYaxNS4Gvr
0e5QlVnFH2er2Ix53RlaRwPTqAUf80ObiZTvt0Q8INhGlLkFOeNDu9RizHgZU2U9
z5G3te/FLo5ms61GEuVaLXd4St/zSDH+jrEOsDeqtex0zEkrNODOFVm+/lAq4U/V
+4YKtiKkMsUZvWkRRAP9lRGnc3bDqqNkgpiJY1XopZXdQ1uWq+pwbLCTUQ8oATvw
fkfBE14yWZqiXAr+6borAaJbfHaMfEM5dsNgF39ksHyeRUIsNh9G15r/1od4YbmG
b8XiC+yzpoQxhFCOL8B/PSVW4kgRFtfehi5Th2dXqz0RLrDFE0aRVWK4DbneHf40
/Yt/FOJTlJ+krHrlOAZw+oln1zpfREviz8bpmTJ37mXEnfSvyrg/QaIaIoAa5zR4
oMKRoOPdcAv8Onxdw93e5TWHW008a/xdMpMHuYxlZwW1B5XhERYVQXuOLSfrNmnL
EvN9Swgno5+tG1GT3zPS2IqOwV1Be4JFAHCaeMiBOJY58HwtjjMpkKUzExveQmlm
G6yWfmrsieGprCkDXGtqvXrFTB5CjF8cyL7paqIFgkzbbNopwoEvCVEEH/W0Pndw
Znay8A+fwzeAkUq5Ayv9llbyi3jPJ81n9WyNBnsZwtWnomgQhDso04vDFmCuGsv+
9u5LCOkRRo6xFwZjAjG9JZYhJP3zPWINupCY9VbQht7gA0YxB7wLQW5MZJP07Ced
GbI8sOl7Lynaf/r1wdgpqBovutbsa8delWLfzMJp0WyYANGCEWvY7WAUT1/KAy6/
BTvY0aJHNw8VhVi8vdHngVlO7ofz/CAPBW1mPCz2zQYFxXZ+Hht2L4865XBP+cb+
ET+oaX1fSJ6MhDMTPBfKqKGSClCuBLK1R2GowJ4lTB+qXwugeYKXw55Ai0OG6bjn
/udl7oDTgWFRXCqNoTWi5JOMfwUXxzX9G7Xu4msx/67yqaoq7UdXl0HNVgSbkgrC
M72Wh5cOJNa8lo4AS40JUfwQDd9BAQ0OE8vghmAb7gyVzsnxaL32sEBowd/dMTHt
cgzQx1VpcPQGJ4Ny5iKttDzvP8+Zg8PZ1ZMCU94vL9224eNWCWe5WRv5IScoGrzd
d2L2vLivKsIzrvxuAILDpnNYbSICSgBT6cq0X6MXz0May3ELS/uIBlVg5Y1QsFnz
WZuMeXR8UVxskSLMhmXVMHfsSlIfRQ6+yem3/h8vFd5OlzWwqYAoYjpPljryLw1s
5tWzOjezCtESUC+9FOaSir5RF1wXoy9rgSLuA0GGVAwAbnrAuZs6Af18Ma+qO5Dh
2ACeceU+p0LZbXUrEazexqH2ZWOWdxA5nG0Ca9Zk75QC7Phedw76uD4heG9k69p8
cZUF3bG1vZ6aVQ/Morriy80aDotrbpEJF84yQSgDL2TstleigsV9qGJmlhAekNTD
ZpB4o/pHbdiTRIAe29xbPSxuGO9aEV+6uuRGpeMftbXU4gchjJZl5cDAuZ6hloAP
2utSJEtWdD6xHFEfmBlgjVEdE4/LLQSBCppk50iwXEI6HhVc4KBfz5iMpureAKNB
gPfi2olSot4uiS2ovpEtMWDoXwJcx6xYexaeflLYtgEc16T7Xl+7MUYnhsxhqpvb
zQkLE9nIElKdJVI7VXH14c4HXCA3uYUTI+jJ5wYyuSOGdnhWxRWCaElY9UjNsdHV
j197Wqngz8cnZNCFSScFNgbg+RCuNv2d50WSoC4wUjv+m9S0X/bsakD6cjJlJPIM
WocAR0Vp8hfKg2k9x6xeMYgwFc+7BXku+GRmQEUcqnzhSNLzsB49XgS21y/rxPn3
YqbgqM9Am/E9c4NsSQUKpJX6uGk08/jMEBqMsLaAOlGM769uC9EWVLkaX2WUfZeH
y/yGDOYydK99nllz5fej6pp6pgEXv3gVXf5zH5r/iUaN34oYTenYHA5zMrnPI7Yi
5JIzRl6NKiVPT8wQ7WExkeIQMbY6npXwF3Gir9X3wf745VT8gbQnRw8Ye9HM8Sof
vB8W+IWGrdaK0WO6alkKbvAtDtL2mhN5r9We9kFDggpkdZ2lK2vQn/R22RBSe5xF
ywmlF5cVvgEME/wi8ba2F2y2V1G2kg6PfwAwfj2shTTWTYHPWK9W/6z7eBt/SXrd
h/VY0shBlCjTLFEvZNLVL+idmJ1i19xrGC+qVfZbG+mSyOAruI7iklM3AlB34XSt
U48oLuYHLFf0ewqyxlSdHt7fy+Y9dqNa6kekTGshoHvBzIGZI8OJOxWgnP0fo4FF
VmxiInCXfJvfzhU3bgD/g6+7C0JhWmuKcEPdYpZTHBt717ou2RVvgwWTR+bRzqBd
yh51Jg6PTdIvax9jFPi4kuUpQyOjLHWcOQNYLKQopUeijJFCZzZMqLs1rig8AQVt
Zw03C2Tb7+lfUOunuLoKrhBE3FHgPTzSIeMNFyBPyDjJV6Ypg2RdU6ym925YqSaA
3PPXBu5gNO4YJuxYnDyw5p8B9xyeaZn03jDyCjjnVXeuqHq/oB7AC+dvJUtimYoY
4SfYwpzCwUaf5s1dXsmHTiadE/JHMItXxG0r2CXr7aZB2tdQKrzhnTgL3i4t+sdH
zJRw3wq33aqK+uguDyAk0Z4itHHTkKi/KurocckoJ4u1RdTnZvQDdNNkh+mSHRIe
s9l+qAHveldk61sGno2tjsj3Mf5llUr5WI9bYmpmRZQJJyefna4HYiIw7zEQK9wP
kDKqqI0kPp4OeUw1pxP1XSmps6qivymUmXQ5NiohUtte7vBsB12tSRaC9dG8SRmH
vLkaT+r6eab+FCBPDAuCokBBpzxYsJmfqzqYWOs3Jwz01IwJASn1ztO6dN+8FgBN
5P9EVbCZn0F2f5VxLgCBPLFwkuaq1sKqaUkm+fJTbKpTYqnVsEw9if9n5ePmT6m0
qgYTPWlFLjrRsDW8hUTaBQOkGZhzEEKe7O36Dnz3t1AOVf24hz5kiyxgP5MJOINx
GaSAjB2RzropnhlKHlT9DkXuVo2m9PTnqsOYj3j9jMCC19AMQKOdJVx2yoovbcA9
AwL2lsXZr71jW/ApM77bbMZDfWgNP5tszWoSqlD4HF2qI1DfWluuo0S/UyBCmC0G
ZIW/g5LYlOIVMg1mLU384ZPYVouherBkUKju5ANo7pXg5C2R8aqFQpGa34vwBaob
EN8+vkKedsX8N2ePyBab22Cf4goBfQ6ncCGkjPnXFe2DpK/I1icZNw2+LN6XN1qz
444TISq1/0xeDjHlVt0bG91b99QZ8VoS0F0FRFmto4H7IDYRv5eqnNvl9l+sIrHZ
ACdp0o/wBJ6YRHHLgwNcrr5N27oG/7ezEkT0jkq/8a3Bq7JtirTFTvN/xOr0DAd1
6ydR+YOARUB+iE1aPcPAO/6W8z6FRV63BBbA4RENv5YDolxgwaXF4ZSydrjMorQl
K+4xhdiSdaElkmsqRqAU/I8Mrjz7Jdj48LjaVH2lTjGe/19O0igBLGgg8HkU7d9Y
1G8s2YsOy/IFwYIh/i/obZS4rFtbpvYKr7kjTmlzMKhEy8Ge84N+wvvFuLtYVaxQ
UZTc3Du/npINIKx1Fl+tor27o3PKSU7NJvaBXt67fR8BSCSYqBgCQjrbcS9xTq4t
YzkUZlHODG6p4d5qub5aHzOEm3LbA0tMJwmZhWrkOGIxOFhcv8gw1V05M+Ue3JQ6
HiMoAa9L/uzWjeaQXueZMiNjJGILeJsQ+ffQppGbwhjYk+gKB4/OeX44QTSYzh6t
1ErmaaEwBA0MwfC7b/oMXwIaOiFVaDEXMwQy/ZAtBvtGJWIOkmaKbvP6brf7XBHj
cU0dm3ptwGBTSmtQSZEF62SKVXfo4Ik+cH6bumo1sXGpU0UIL3Q5omUmi1UV2NLA
jx6cD3/XQtazvttbqyZfj9JS9RnohWy1o4aHhh9daQFkWop6ZDO5Smh1ce45QIjP
DjbiYRgGkzjV1fN3+VFCTXeLPWnw+eELnWZzqu+kp+XTG8WabhvOnNxCEHo+3zFk
2mfQsCMVcklnmf2FssdLIJkwdL+Z+zIJVA1+NvU8IOdZwDa+ahWpliey/KsFRh4P
ekAQk9Je/dR9v/JcwDE/cX8viS5wwg6wWbG01co6rUeA9yF46i2GZfa7fiEC9X+6
kI3OXgcGdEFOoJQCvkmIxOgR9nCE2GTcc+idhubFpdgjUCG3juziVzcIo3NMObPL
3ZGYM48KiwAetkgWbxvXG/kfFfFOMnL5OcTLFyBCQ/I4+Ph27H7SswtGvEKmTRNg
F2rYIt8RCAMc1g/KrAXfQ/MKz9tHT6eIUgZpUp5rkkx95eF/dvaJT4KpxFntVj0w
jRz7JGUxbAh6y0UsBNQ4vSyEqOcB8QXZV+BWOyHR6tQb3pNhJzypvUikk+eYe7DY
DlZnftf4xRPfx4FFhN005IKlLVSt9xyXhbQZyGZL3Z05huGSWow2wsvjfcXq/6oh
iU3bjq9Qth3/N6hOGWxn5n0Jdm55fFDSG26hU0/IaB+U+x+E5l8ghANiKMTG0LAt
aP92C0pC5q0ZIqtQf/AbM5DZd8S/QJHeHQVpx/iyU885LfH1H+wX74X/QSKkVrDb
bNDAJW+60B36MpaTZr+sIDN5Y299PFmWrh8Feor+R6qfSmyXZ5T6g3sZ6LsNDQoI
GaycIvnMNl+A07qRuqSLpFIvGzuMRAi9dCIwbn095612Lez2eDmnDuTw6C/tHq8p
7hJomIBt65LIagdb+iF/CyOXO8aDjUKbJKlPcZySwb684I46e6dw0lGD7rUG66Ur
ZaxFXr93XJeFoi+fluYKp3BnA1pd6fR4HKRbG+vLvn/MQmefgtOv+UBR6WaZiExG
Fgniana+X1hVMYV8aCi8jnjYDs9O/6u9uCpSuaP8Pe9DUTaDNmxl5ssUN67u/XLe
lezgJUMzvkcRoF/8inxjjY15jexi69stmRFQb0mNfhxGZ89k23LYLItyONykLlYp
pj16yBykK/HaqyR0HyIGLc1Fw5AK5dKm79LuHmMKucpabq1R5GObdamDgr4xg+eX
wlqdYy5zd2J8NpIli63PUnU5q/0chPwPKMnV2+8GaCavFL6sBuXtAGFazxe/dPe6
07cnH8AkeS5wgxq7rJyPjv5R082K5w4c8H6oStDlCySVJ7g1FoI0IUI6yPMoRm2K
IkPjiI38NxK2esLCERQLr/E1fhiZRzRlFNlrWXsz5IA57RdhkO9PPd7qxE3dmcnD
n+cdQxj9vqCnZrcq0Sca8xiVxgHtrYSmClTmOe5Q0m6b7IssNV8CSg7u7xSIVHEN
7ZvHE8KSUM5Cap57fQ35dWateGJ+KeconPr/L257JWBeOfHnEbk72DdJ50h8CkJp
S88qftmi8irCo+M9sq162d/AWIn0sF2Hsb/MxvANXGA57/KCX5an3UN5lRDqej87
evlrb+IYJRokvP42y1Z4NnVifud2Ea7xwmA7+amXCYBRJbI3QKdJR6znZnlkeayI
DhPnHaV7huxG2lKj2tUFHTwlpdy/aClI43oKfsvZB+CpxOQI6L7bJkCyJ+5sjXyx
tBJ/qPwBdJ1SrIvGBMUeU9kvN6Mizvt1DS9MC1Ix63dizjIhwrKVZLlVGnSe18h/
B/hqrLiXP3XSk3aJXfH+fnJyFY1jnnyQL+fU7vkCD/dlHr755Ob9dCU0Hya2pcX6
QRI3wUjza0ri5RWORagNBOCgcVQWw9Ymc0xtwg7zg0j+EAKIpjmqdY5tA5Z/iIkz
D30OnfmkSUAARzOo50tx9albbRDaxa2rLWS9HC/sncAp7XyNO8LWe4WkglXG8jr1
0KeEyHUx8bOSdQEo1PVbD1U4IF2lrC9kiI8Ri8/y8XTJZf2Ruc9ZQFPwcQZFPhOk
zHx4MOpIvX/43/mKkry8D7pWnTVsUUeasRnrXjm/QPn599pq2kuYbGgohuGHmv/Y
Fgi6C3SgZQ+xTjjHwchJxIr+RmH4P4550cqk1HLm7R4xk8U81sCRWrftgz7tHHQS
kuldroyqDQSAzExW5wVy5zWt6y3Y34yqkBJCVx2TwIhwSR7CTvSQ61yQXZSjfhf3
WSIDPn41pFutDacWBRgMibx7OoCWgHdwXzvCqgEyj1dhFjzM7F09Dzq/f6sH3+qi
nFDmEZ4EZnjZs1cqIV0mHlGskvqK2SIbAt6ncZdj69qN89UG/2dT8+BMdAQeIXS1
qRskhH8nvAtvqCiNxaddr4dkKq9WnMmRx6u4fZxEFDlzNjsOJOoQNNlATUjHGTM+
HhSIg60Vw6+EDhnzKtCFUw8ZLp8mXYvJXk5swYHb3Jcy6vpXKyoMxQUKqkhmFGya
DZdRIPh2VKt0Lyw8C3VRv5huCfCvMQiqVAYu4i5L40xaIey0bllhYZ0SqqW28CnT
g4Dj9/r7sx3A8aGBpMi2+kfMwm7qbgW1PbKyz/ox5zUeHi4UHtUpzMD6HkIqNSYB
rW6PotiPmZ/8nUN/9FnbZ0aQobqDAZca1CTUjeAKkRmFJMw5Sg6RzW1ekHuRYYiO
wyrY4RvIxXtnt5tu9mqk9sisYRaGe4HJjVP/8pn366TPzmNy74Q4BrxgdO6QlpTS
SDLXyoap8hbwpQgm7DnnZaXEJW/YaANXwq5DzGsRRlqoB4u84eQ7TpqRYroSj8sX
JCgUMt/uMsFWIS2HipoZVI1WDIaXqysHbZoIl6n0CEu0cUsWccIF/vsgky8fqrZW
i1GZkiS6XKZLmj94wtrPsS6KxCXTpMA5eKyMeEXKpaLzCuC4T0/FhrjBHEfUu8vK
NvCHCJtQmEuAixoC8azLU1ankhvWENzbD5K7R4oIoxhL0iOMahkvaIY7TKX/AV2S
0fI2KDDfR9bnBXhjRKpSDA1ZXW30H/7Ums4N30OXEI2Z+Ef8qcPUcthfTHDb5Sd+
M5iRxhZ76y9YkveauelvMttPgG+Fh3Tmfnze/gE6+/HjAzgy4mTPmuHkhqXq7vhc
fkCXbnPxzeyWFbdaQxEQk6MxxjftF6Ko+aYebpTTUMkX2Do8Pg8aDKE+8YgCJEo3
ptgtOOUZ5JXrCPw1/vWv9+uwT2MzYQCQDNvm5a2QVevP9qnhn0m9z7MjeAi6YaMI
8gkf5G6NLGuFVNLoNLjKicgH+9ec8aEjF9J/6uVYaK13tBRMfVDB25bewUzPqEnB
xnmcHG9870xKDySTzEbE7Jowkxfoy2FWive9e+pD3uHi3IgmcDoYrOLuSoMq5vv6
bNXCaQ863KXlF3sQi1vg9qsifolqNkQM29DHv1kTq3PJe6M0cz9l2ZlvSnH+RZmq
F8RD6X8RCHHSw15OU8so1MMNJdQ1Hy3g/l4zT/VK6c3vLj3d72u+Z2Lenv0G10EY
Vy+lB8xMHp4jWGk6p7Bf4EUAn5aH6Btn6NAT8VM89VI3eYnewj9SUWca3b/e55cZ
/IemjS0wPu4iXG1kjLq9bxj4ZM36h+gQ7UVdCu+YzeRO7RqanJRmAtAegH4BRMCC
EJUNSveYZwJ2GBIjxXxszblcvEuRIjCNTaQz4hWPkyAF81uIyp+U7dulp4SCBENN
n3DD24cyB/7zyqEX+7uTr79GopL1oJXJtM8S3mewDeOGLUklfjMfWTllxAH3/HWt
vID8cBI0b5Ew+SFFAIrogxNU1p8H+Rgf6aTlEgoSb+SxKa56W7PVcbRDWhvIgBg/
Rkp1bxW4EAwbOfjmToQd6JIpIcHxTXQYlPELoqdHmrPkmPNB2dKgI6fQ141j/oo5
0Rk4pusU/A5ntlbuHtNi02cBlG6LxkrtHrOywAlzuRarzZEDgivsYlNqitIM9li5
y1fWM8v9jQk8zX2JZ8H/Nx/EyG9MvY7/5Rj7qTSWLKhzDfoJnPYP4gKgZHBIfZyX
mcFbnpB4BvKPY16okek6O1p8clhJ8wWwLEQmfwrVKU/sd2w20daM6QNqm7CaAdyp
ARxK0eHSfgzTDNOjaRpaVPhNQpE+58evT/DfBtMv7DNFz8z0AgtGGHFxWs6YF8PO
1uLkqtEHMHE8XG9kiIOS239OTxa8/eLjBx4TVvUFtxmQINSugIUfEGWsweUfxFhx
I/PbGhq/c9Ulxw6Q52adUQ9nwFrNCXZk1jv3+fzoEjodvCjPEHQJYhg/VkN0VIT2
yPHLa53e2MVfolQXgO3SwmOd/sB94jJypUO8QcfuydzS/5GPidEzLwdLjFFgr7Yy
Qk4ZohOq6sGKUH58MmPiebBtK3Mnmv37hjwYfN5l5Tdbyovuiaded2VHn/mEtYxj
IwaizjmlwiKwv+YbZ4z1uvXPtIqbeyiJBE2NU7TUiFLUbZy62B1qdzbbmDEE8Fkf
0kJPDeUDzNhskmSfsSMooO0VO4YrssDdkmvLogMlureVxMAnAQOaxJYuaTY31lNI
976pFv3I8isBnXE/Qtb7Y9af5oi/d5Xy9gx6xygI9pVrAxs3R68MgY7g677nCREi
cm9LtobN5dOaFZHfAWkLeMkMNFNak5+v9Up6bAmw3vxfElExkC0Z+5J5BIfOF30X
58apmQStc52y3b309w32B/rB0L5o1C+n6QidYYVlbr808EFwHfssz/NKh83xbexR
XiSkPW7Iz1W7hrm6lA2p69LlHJxLHq7/9GATLhB83oCxGIbbrJsaIUtazJWzf2CK
XHl8cQDQGKwZAz6hmxZRkbxnnMogsKe1jJZ9h03TLLm7TIFkpkQsE6XDOmegiPBr
+WaLJ1IV/TA8175R0DDWZrDwlZmM5jLZWOssjB+gSUZzjMvGkYU2EavLkB3EbbmL
0mxY/HeuSDb0XdGN0K4DR1wyLXw0EbWxlsj7jaWFU2LlWiqqgG6PuS11oTTTWXQo
USOA0QWpVHT4rdfv7+eiR5W4BeQf5bi7a23zb63/G8kUuhuzsqvz3eRY9wqypDfo
Xctw6wrvxIiP26bw04tFdwgI3qTQyXpVuGuvlaanXPVTv7hYjlZ4t6p23TGydAbZ
zIeLLZbXTTtih80EiltmDJAxBVZfc304YFceVO/SsqJErgkV16y77gZ6IQsiPc4e
RT9H6ssd+Dkz06oqQGUApsVPDu3OqxeAljj0Oqi79ID7nOPRG5WYc5wnP3Kb63Ip
DCGyG2ALySOd9iWUcfWXyldMo0WV8P4UODsoBlaMK40Gt05pKE7H/0XjLImbPjqb
5e2mEWhBCqddGh28A9Yo+/22PjzqFYNHnTexS3vuTPmvob/TbFnFUZj6CQRdNxEV
GEqvIBgOuL45jGartBnk428Z0frbWBP0C8iJqE+CsZf2XR5k4yS9X1tgODMzmz9Y
ii1b3D4aQtbYCLmt5fjMp+ox+9lODZ1DYuFF8Q4Tp6Q49GcnIJRUQKSyaRANB2MF
lIGZHrevzBDRWNpYo/1UAIQWNOg4jYdQIce3K1EvkD7V+GDSKZ7bILrSzFrM7Ggw
nZDMz34g8OR3xdlGuW8i/N1HPjMT8Nb386U1JU9hDzJu+eI/caXT5LemM1MeTi/l
pEa/fenFF84oJdXgYzK7ztgvjJLC1VgQrB21Ei59XzJTYHsfKLFz7l+EH3VLad2B
ka16q1J5XwsBiH5K36L5Vy1tukLZjmGGYTXToNak+uy/daNaqrgpFxgFrBm7fT6s
QnBEtQR0vjQY+9tPIb0rXjFL4zkO1+iQ8rueEpGcGcSQSdi0mPjx8m+JB2khtQxk
0yBfWVWRZGLCRikDhZy0l6HyAbydmTGvUnWdUPW9BRWAVmbp1TiqDy+2daqkqfd1
a0cq/O1qYO1mFdqaGb111UIpv1Qf1T681fvPpPM1in8KO4rO0lXsoVnzWr2utRci
hp3WnwIdel7pG0+aUMBsMBXP8D0H1LTrKtCYEsmsv00lCvI4hCmw8Mb7Jy8MXNeP
jRAFDq/ULRaHHAgUf0Mtu8kQBKf9WMX8rpoxGHA6iF0txDFR+jj3JtUYjOsPz89R
DpHgqnLRgvUQ4CBY2f8Y+NqHqC2nqSU15hkFJJArxUDjJEnmS4U1NBkWupdT/Z7q
v8n4jsALpfcJxQ8z5I3jD/rr5kFyfBgFddUGld80RbAUnkt+jw/gANOmOW+MvBBP
P2GyBLjPgFJ0AkQ7U4EtMpmF1rCyBdWjRjLsara+8CinBMJG/gj9Z3YApbRE/tEj
pPoY3KXIl90IKDpBSABX9hoeXaKrwR7ZnLZus0tU2OLmr+YqyEsn2LlL+3sGrB37
8K0a2AAOEWUnl1pCKbpD6IUtx6a/Pf3JGe/MU4Np0qp+u5Y3SVAlUHniW3KLTzSL
6nB8vabMrojZMn6TAJNHoC+/tzyuVSg7SUfqQKiKRXz2cKRjIowJysorSmt9Xy/q
BksxCZ5UBloo2qfOjiuWHn9AlSXlqx4eiK5RNUeyG26bcPiFDPaMT2r0luOpODGt
AA+TQGj4cV7guzWBB58XVNnnqur4LrOev+//AIf/vRz7RdOX7CFQJA2OVVYqUlaZ
t2p+nBlcXx2yNONWmMFsAJv/EgImc3yIlU2FkJZU5JJh5ZPTCGAT39oUftBjRk1h
fBTkTaliwjFmc9EawaWM6X/TOSAbwkpI5MgMbhVLCWShQnmt15wNl4532jGgtSP7
RJUQEhAs3uEQONlpTR5GTyhR+sVtamgGKA/T+92bZbIrj/T4ZJB+lXWbStl4iUZl
yy+em7CqZXdhNgqclTSifTNS0WdXf3aOA5jbvpXfEQBhAsbKn8zZPlX6uEFdfR1K
2gfxTRmgTgoP6btNu1fy274NJwBVSPZ/Lqv9cxlkF6smEM7yNLZQtWaetmZBcX9B
8IybR+wocQ3kT0P/r04RiIQzcwHqvwOziFvvoHSTvUSETrY3Fk6NRWlCThcfRfNF
DQqqvFDh21ogvmnEswerAIdMm4Cym46wF155BR91p9Ivg6BpOqqOsPF/up648Od4
UL3hnOfdsK2/PCBr5c0mf9xJ6OJoF7DP5j5if70/iC1T9opOT7nZyQzXAZSILP6l
NRefQklqZMmI2HRFp4mEMJhUo3A21tC3n8T8HPeZKjqOjiG1patV2Z/Rvb65Yrey
9tWGr5HhUwjafT5ZpkacGo/3+ZCTH/lOYus+IsCNaVM5D+yt/gfALDVwJvFs/y2v
hik4/IEM2H9FLc8cltw3g46w7PxTxsaSKvhA+PgSkWI1CnkGmg0joFkpWevBPQ1w
JqS4M7GVkgMcP2CYMou0qwgt3ySdpy8NQsK9Wwme5YD3eBJGCtex2NrvXEJIt1vj
cTejqfhxHIwjtG4IH/mUzIkmmApEESY+OI0vLmIApQjIMtqIpAgQbFz2Jm1h40Fi
4U5toryOICSllOTs1zl+4Jf67izTLFCDUzTLV6jfXijqC5P2XxqTqbet2LGNH8hV
wbCggg/eZ0SdvOjgBm9v/EZQ34IzV03zXYCBWECRWay9b01zDwaO/MGChZ2RsPIc
7dEMZXVEdcIFsB4zE0pJ/DNc/WKVT+krdT2CPxUDMhbkjbl6qKm9/m5OCvDHykoo
/2Hxps0K1/02Q3A+JhctYF/eEz+ooHj5d/V5olwo9AgCdzPlGgm4fNUAKUo4kDwr
3HsxXmC+/twwNwFZYRoH0YztTWdayqJ84jF4NdQfyl4Hd41/ClAPDhqlP2PfCc8R
mWuh1wte3JSQYHv3mjMAP4KukI43hs4cE+aQHkzT/weInDZ55i036d/crsfbz26E
Pp3+sjxBIfxwzVSKyl0rgG/mRIGWNVoVp0R1nuvSYTlpVN24kW0DdTJyNxFQm4LX
Obx/NXAmrgd3suEvvdidtsULk1gFj+PN7alMF4EKYSV8TABO6hDdbg4aSd7hMfw3
dMw48pbUN2k9aKLmxXYkGyk88TydFYK2pYcEGhB3KBkPfEk0sy9+mh3v66nIiK2g
kegzmBXxDF2qd8MsJ6Rd2HI91guMu8jQYVxX8AR2WB/FtGBTmTiFv2XLivjnUn46
7daVpB8knvYlGRNIF4CAVGIAPICKM102V5YMYaqIgybgf405p+RAfwP4VhDei13u
Ku0WnPo5+7cMOCkqjbzGxRdwe29xNc7nnVt48Kkq4OLbTWAOs23UXnTqY0brMGA1
AjX1VcC6bAK4oZrvbRMwtv8IWvXsUnCO7zTUbFLvl6BPuAiZXhpS8eWtsELMgZtr
DdyLN8Du9HYT7D18gDSmGsBeENPMGFn5DLV0WY4K30jUoUZFehV+NMl4qShR3hhB
esah0W0LNy2sUrrq5TLM6MyC1pAnmZHvzY+npFCrGtKv9sfdKRfCCaFacaQIvtcN
YFJhbXubonGhlwxpQ/qdnJnvoFAb7mDDE9WX4zA1AgqkaMSAaSncylwXggtRnnAl
E0L9uM4xXhGc/uI7ZHRUswsy8rUwqruirs+yFGgi70O7GcLuLscFIqXwMswF9W/d
igDb5g5igq6FrQCPdcbWs6LxIJbY9DYMpg9WZGNEnoJbhVBS9BVYYMDE73M0k9pc
EPHbyognH+24LIQXpKYWFRGgBWAn3RtlB+PVVBz0f0QWPj92zZCrnZLgxIX8fCpT
s/YXo1qGQmX/YoZewen/TadGRdwIMm85tn7c8Zz3z0Wqlj9jyGOLH//Ge48HNFRy
c+0OdMLDSBKW959aCfuSy4/66RVFg5YgGO33B9WPvNMs3ktNSJYHi80XUnWrshmt
fqd2bYcME5wBQpV8Ahjm2UQUGJt2FHe2ocCsl2Fxmz8HrBFbbb0lQYKEJP0kXc/1
rFA7WNryOax7mYvV1trAA3i7lhl+pcdeBp82Hr7skesfM/biL9m7BdR/lw5F49CV
ff+GnApOF05HRI/39ctiakD1wmhR3aUGaaYVJ2ocREPczhspJy/6HXf3/lzRC/1m
8La5UZyhExpJXTRdqzDBKBPJRTquAkWohLhL76rBSWJCOJo/xGm4Wn3knrjuFlr8
064LmhkdWa9zigKRclDLMzgKGxNrifll5FGrx2Leu2BUWSlTZFtB+0izJQJ8ImfT
LZ5r87r8yAfvYcBepjPPk2+SJOiV+GQ/6ResjVaFrvnLXluHJSb1BReaU9PI/NmI
8j7jMn+G48/uEiDQ12K8YlZPvOmDwwbvt/krABmwxVvER1P/ixU+wdn8PuRqHdQX
sHYl1MHOj3DDHT1a0vSFlQX+wLqfaJJp5CRIx4AZLMZA/4UQpG1xtoAMgtcHaTd1
bkw5KwqzxcMUOYDge0ATggP10YpLLoNtG0+qVmUYYrGgjpslfO9HeBLrAFa+34MK
L1mTd+9xn1tSB3xJnBABvnixrqquiYJ9rXUBAYlquhzeFF+KePonMakCaxOG2r0J
3q/O9s2wmPN97SGAcyEm49N2zVkg7HQdL92gk1lEJ+aNXe2NGcpZcVBCaxzQWQiY
+B13riJYJr4ke0dSAfohw5rY22TtmpAoOI1OOMz5gaeYiA+P8QUhi0TnXSLyvvSz
0CA/tySUGwInA6QDgickmIBGSVe0iAwpWJkM6h5AwMl2rRJvMZUqBhK0HnIbq4jk
oQClXHFjt4Dz6moR53TE5x0WD9i4ySi+5j+lpOkZTjQ69AZz77lG9yYktI2pvhUY
O5ReVm5UurQnF7/wYMjK21r9KYWHwmadCmEpV3UN6OH7j6SQQPEwWIhvJ69NZ4fJ
hq+dTKcd+cpRHfK5RWH1r+qTcIKUzIUNEtiKB7oqMfnrWr4gWkRBPPTS8WXvBnZF
EmZ/KCMYyfsDdfnG/h/2zVJyXYRxQuSnovMf7/W2gEhX/RNZ8bDMSwmJpV3XEZ7j
gxyMO4IX9sAf7YOVJU/GzYyEyxOiDA6iH5UVCmJUQQljW/SiB8GdoeGylAoa1tz/
y99V28pGYm578bKXEDc25h/9haq3k4BdyrYdxEuS+Ia+OH7xVOvrn8VFqbBjdJo/
L3pkWcNvGeyB2mYUhtGHOnL6wCJJOhPqktr2hExTBa5yavqHfQWdzU02/VsdXy6G
mGo9gchjrukkkmILcA83v3fsEsf0KDN2VGmzktvVwybo/Zf7totfcHmv/kBsrk2D
AfN+qTVdWFYlzbDEZVA/2tcRFzmzmeHyFNmpS5jdOnQZBFN7y/M274CguN6Gi75Z
6XtpMpIoqV8t1JBGUbRCFdQkBrg+Zfe8Hvz2bxEGQkAhGCWcdPji2uStrcAPbrW0
sFHgM/L+5ZYUgKDw+jo4+vf3hJihLEFd1powwIscuf5BnHcCPozURGaI70B4B5zX
E5lMGzYfAoUW6mXgr7rPQOSWR+g2XQjsbhbeyQY3IV1PepL9atG2SJNWauWnFMUT
xt59mbasT1lIH0ITd7XRbfgRiuTTEnCje5kNP39KXIWv7KOlPadQTdJwodmpuT7G
knqebsZFdnEF+VcohE3q8ERQyt7twSyfI+3Pc9wdZvMI6PC0OMwZHH7VZuDAd+Er
/BuR5DC0BOub2B5YF/XCy6sntAWKBQf59xiEKzGilKQLGHGgIwTwur+2YyE60TR8
ksw5n9uKpfsZ6zwrBmEBH8eJrPy4MjkzoZHUklyOB987WUFLklhyIpDDsXDcgxRw
vRDwFAvs28u220CGnCZvlkir1h3D8QV6yBbYPJSZe7yIqjGva1xSjAfCUBDzl0Xk
9khO0AQ0ibFdHl0QOK9CtNaL4uuzBQpdZ9uRcGLufnrGlvhyVEPi9SAW5CT+CzmX
CVoPe+M8VlK55iGjXKDhf1MGibXBRwSqS5qSL7nOh5q9f7YqHk2eAtbqbz0ISyZx
51qGhtMvEOE7yRRtslva6oDQpFeRiayJHLfbr7PTlFc3SkB3kSpKUKaiOd9lsW5G
mEs/78rw/MBhTXPeQIoorwvFRRGkJ57ae59M6XQN8bveQ7YvOJf+2ebPPsbbC+SS
eViFae68rnIK3NwCcj62+mxRZ++8Wge+X7H/UWfl72CqvX76qN5UwoBzkv7YkqA8
pYA4viCq32Es0nNIczzrlWzqhVCD0WUg80uPZjBiE03V3MPFbFfhhxv6Y+KMSQi8
jhcbiUOceqUyNkWwAXXJo8U1mQhV3mOZUxAhdDCoBnTs/f3FaNX4WprxU1VM79l1
R3SgThNi8/629VcoQ7p6fuRFFHaXKgT8ea1DEFDWaPEES9RyF8Ef75Sg+HID2eMc
ZYmDrKDpmkn9758DZNgouQoAHh2qzyIz5KTnEfBnoPX/MHSXXlt6bBidpYqyx95K
duJuBZPWASgrDelq2fvo6hagpZDIMME6Pk2LQq0Hoh1akv8+Cir8V3ND0svI2zrm
vqibcWvvi9pVWoVVD4vZdACWZqMja7msw/udvyHePtb+vGECOZtXc337rnMaBwak
Q5exu//bvSvP0oIvbxu9iNyUC1XewwRd8EHTY7KeQJpw4VigAUGICf1z4mTGHxJd
jihvLFV4nyep07bW1jPP4G2bk3yxNaoE9b7IHXJW7zxB9noNmPLcaKS9fo5dOscu
H8+MzYiRpmUeOt2KMs5nI1QweXHI6gAxrWQtCxAfJcLnkNqguTgboa6nVfQ703Ts
N/Je6KEBe56e1sAzMt0aZ5emdVnzkqfJ2f3pb0o+fwukgRKTrfNKKODh9/nN05rH
4mZ/ajyBDexqLUvWYrMErGw1FuaCJjNj5hAGZvcja3cuV9em1DlPZ0iK5vk43zo5
MejLdHV6dT/QsqdLWZwTGOOfFmaCphw8SZF41SJTBCSxdzn/9VWBHnm9MDE1fYvo
+M2k9ldCOkOGRtcPtKDJRSPOSf47z3KX+F+FZWqgKFZDKRx6Bv7gCzZE9Az1KICy
6V6q+0+4BxmXl1LHvp1M18nOKmv0+q0PG5ZUZVcoadtcnMvxE3+n1Z72glchvjt6
hYPdo7ydYwDCuX+v6ddlgor/ngSgacZti2VRuyhxbXgDwvSbkU56l9HQySpdvEBY
ytUpcsV4lFv5UrQc27gM40GuCRXUi1SCYFfXO8hjsBxZfjklB6J1QjiitKPcag/0
yrfEor8u7lgHl8wXfruoWMhxhO2nz9Jv+hrfUAdnlTkIwBWmWiRdm26BIqSY9nFi
lKa/cFsgFonZrH4Bgpb5Di7Y0rpP+LFinX7Q/+f2SH81s/PXo6AYNxzW9X3vbKKD
TF+aoHKUZLDsQxrF+MvfplrQhloscI9Gf4+a8JsiX2qYVQCOpT3XEMUy/DwQLUiD
EZ/gIFlWvwhHAqQyPAWLcuxwwJcAQeY1K6l/7QWmjVZ5HibsGExy1ahyBXWSsfdR
MQK3KJYFCA5brkLD9YmaeYxk6f3yI1QiHx/D+bP3UW6TrqyYPkG8a6F52mJxMX7J
rtVtj+wlIkHHl+nKlRajFQo/NEOSubRQyjlSq4BqXGjpZ9kIb6YmPQuRf6nMWOLX
99L9OPRg3HUabYd3ypxpWAyM23u/G5EvRLgDBOZaBtizIrfvc7FheLXwZnSwmy4m
pBjxEHN7nn5R1dSWa5Qa6FPBeBPdt92sWeMOE4ZSqYfF+z9yr8OrD5nYKJ1jm3p3
vsbqI7wfI5JH7W3XSH+NuUFLzn6Dk/Pkugjxn7Xm9qtYx5BBqles6lVWMqLjKL+r
q/g5tNLfwyHMN4GztJ4oH4epR1Vl/EbfUQW5bKEq/uPMFF5FiUczLeZzP1V5y5TJ
iqowORi3PvJEheXtJFEQRwl6wQ19BSRM8b8TNVlIZWL1W6kbI5H/pQWUS7V0VWZf
OsEah0JtuaTmKAqL7Vf2RfhfRihQ3dMeacTB+McKgiQy7uL4bDDHhTRovMbsmOuQ
FD0ZZ2z3YaeDU9+uYYT0+D96da9iHcRy9WLeLgp+XmFIaHk+uAd8AHARguf3BGVv
tt5rc7HFmiOv0HTf3k0dh3DSnJlVDf65wdIfuXmx6aWys6ZsJBUItS7N9cJGbh0E
eFOjwhWxjSlFcXmoXUWBQQqnHI4XZY4AeUTY3WXulBjvfEG6OTgMHcmIZDcbGojM
tfsjXuo+6hfBnYCmNS7XfP4qmaxdoXokyTG4JxjeWJe7oqzmXR0lEn6qR4LZ+Iz9
t8ViUPJrIwfSbmXQA9KiW6HzmSSz34EUO01+enjNFV6uqf+3n7ZCe56WSb6JqC3V
d3hRSM18XwbyFAj/DD1IlrDweKloWY69dR2D0gKVqnn9q+eoyaJcnvCRcFZ5cRu4
RvMwGAEmVSRXyYXRLPlkWKDFE7h1qh6afxIuEi6ese61wj6MEnsehIdiOk99K/nw
HV3UY3L4rZSRxVXNs62DCC3zwdv2FFan0yZq3T+T9AF91bGCjXHrPcYUbe66BztU
D6VKmxAoRP0FkDZqQpwveBkgsY6igUAVE41xaRnqKqyKu+Dz1i4rPjlfpaLbQnSJ
m1SmqKqZ8Hvp6g61t5D90JqROE6jgOAl5AI15U3m0eIm1bQy1aqZIPFK2IPeEFBf
NkinGz4wqWUnZTQ1tUihA5kpUZCj5kJORmp4d5i+z9Bm4d1f1QXduqZZHOvbn4fA
95bfh/8gP7KQRvdB3SBif//ZNeQpau2PEQmk1D5TEqWZGwAIn1l/J+zFa38LLLE7
DNLfwUQPNFBh0NmhMY67g/S5NXoq6fWrtrSAAqb2Fsg+xt49MZj1eXZ9ydNd1tId
0R3d08BooIFNT5xZGZ6hd7uQ1f6SY8w4fxYT1zyRzX9j7DdmJLhVJ0VK606YDWNt
pAr8/Sxk6L80XC4I67q8zC8zHv09rp/rZ/G+/YRX4EZD9ag8/hlZXeSxWeb440rY
kbyusPeQxIm6VTRFWBVuZXX7iNgK1dhVpGhgv87zVX2QdQ2bfCQbjXWVPJg1AJ19
Hnmuyds/5cZUYZUCrnFNC09ro7Xv3ctm5YdoRFTZ9+som3hfn3OJUq8SJMgRlqoX
CJrBcxFeBClVTp2OiNGywVaacOo33/8I8bIGg7y0Z/DV/xVanjQJHjXaCj7HL6zk
MiWs3OYJ/R63SV7QhUpFsgaILWYCgNIoXlYgei27BjQX+ZqmvACKPNTQEmHFQvB4
OqpLLtiTjbDoO6Yl5l04Hqyu5L4UQ1IwU0kmMgBR8Qx3wUcNl7KciN/yfEBpYKet
qlCMnKTlXv8KbQ1c43orHtlzv9dSFz2xNUzLeSDXVfdx/O3Oxon79aamOhHRYsOZ
yfHSzjlKIABWSa2fWFg0XJSq1xUiUplnu8p4REnfww1Ja9KO4OVWBnr7g/IQIEgC
7276zeCUuyP7sy1JeuJRPu4PwtEVprdFOFhnr1gd4F9hQAHjK77D+a+fLIRvot3Y
gbv5PUe2RbyhxFEVRU+93342kXkho8qEh10lCoOPONLFhuXmqkvpofW4653CVkr0
66/j+lrnT5iNzZOwl3kAbeka7ToO0Ceplov4t6O4jpSglEWyxChblIur2v7otJae
WKKUATxAMKJ7JuB0RJbs7LuUcLLixKJfz0V/QNBqunhOaGcxr1DmVEW8yzAnh7m8
ztcGD6/ECwltmONq0QyDt16DgGTXWwfAWVPlP18DN7Spmt4808BGqVLL1CHKO2Wa
u1+aSzMH7n4+zc1RER6FLbIsj5Blw2JMBGXVCxYgJMPibDeC5xPHn3FK1n6S8cRz
LqRBr5W1GJWQc3jckFhkbKcwB6Pf/GoP97/kMaaxnHxEcbmw9FiWh9l287Oj/JEP
V/SS1ykRdYBf3Pfeu9G9u2uCTo62bqL8uBwQLm0Vy0JGt3VQf56Cximj4xZqgXmW
4VaSlxy99Bd2ws+TU7IawYY6SS+EFBygoXEdrk8Ijo6mqXoUlsKQQ8AD3dE8Ox6t
QNR0mejtmRpshzyJIScs8ttZTYHxDzectDefcu8hl0VNojcTS7+PCW42jvMHfns9
9aolDyoh/XffPJTNp/dGPpXW+uebZfUvnuGoeTymfr+4Uau6gNGWV5Aq2ePs87ps
yxzW/6Ov3jWJLu0fVNZ7PFQPp0jBdFJKw1PWv+AAUcR2sAYn3lGaJ5tD8wK3TLzR
J+o5cwR0Vm0Iop4qhFX+QCY5a3VX9OVg4a6PGYxndVtXEkEZvKmYNKwafcz4VhnM
LDG4Pu44MjnGsk+ZBWjDe398TYVU1Rke/QKpFwDOp/swAKhVtXCm9pVWHjB1nf97
1Z6nmIM/+ziUjxCP6okfaroSBz7D2IOi3ilLo3WZqu94qw8l68ZLE0yXgZTMaOOZ
KSP7fxUZ+u8C0hXIPOyebjmedg5YogbSguEPFfkOrr+L3cxRmISqdqq8RcudPi1x
fgcopbZ6gf5zjPg0K2p4K1sM7PXCycFMnXqU+1eGV0MknOfnAqdwHRkowPyM92LN
Srzf+z7SUNEdePut2mKhFPQYHuGdp/IBN83ZM/Cy8Bx3ZdeqF3G1OS7MslsP9x5e
pjwGpED8G8OwqpgP8OWio0M71XSOmdpBp4Qlvqa3nGo5YDuLW/K1FbD2zY4fi9F8
fb7joxvZuvvsjMnWBPBnZODFQyXUKx/NIjCUPjUNZHtBU8NHpW56qSNfw5Tz7QFx
IpFtqRVSlh+IepBykjSFiASj1XKDHJGGol9ZeApplnHtUFZ4P9rJSwBZq7MnWDFm
UAAFzdT8c3mefx9CoU6b527jLOzK9SnkxL/mJ6MIVxZ6qPOQ+u8/otoZEBegX613
gsqzE1hSNKHAnivrksWa2Do2OCHL0qIAXfz8RqnO87p7qj3lENGGXv5N5xag3SYL
sLvLIRJpL6cVNJS4slhicrYK4dnKd/Y6qD2rPrPjccsYzebSK9lS85Oi2vUwcsWf
+z+PlV12k3wVhnhpDq+jFvn3diCvYpa6WyVqRnzkjzCaSG/Lp4osETnevK+3+drE
loq/E8azVCvIPbQm+jyYYnQxMk5EQ8eqOQftV/fu28EAm3RYdxM4ibJO5TfXEg/h
Vhgp1SDu0yR5kso80C/Kj0U4KtqX/sS3gnEvqg+g1gVwQgDpUVC4EE1Alx4KZenQ
xsaf8lwt5WsfAKBhJXM3aNgzuYq2CHl6+EhcbENhxgjgtKtjCsDMVGX2ee6y8HMR
G4J+Nd1zvbCqBXg7H9i9JS68rfpUfPlDx1BHgSf+fz/R7JraLzT3iqMJqe717Mpb
TVSvbC8f5cwoQh8IPUFr8g1B+BjwDKtUe5QRIVU3Wv0WY5aP+A8zfal3KZpoUb7d
Qchf57+O2vEd+HNmrVeP726KlG2vk5ACaomkDTuagZGrlwkEqb72B7fKVFPsxbD/
0yyY++ZNvPlsEZr5c6aJEe4lSEv04j7dmTy8TCc48DianMV7Tkr2QtHD8EWkjmnR
7mvhIGnlEVYPr5XXjR/28UBRcMZ+LhjIpKquPMduVeSHdxjoFru8Wz4TnfW96yVK
kn+xBIFmBKxZnQaPAkydsIuKCga6RONRVI4YN2tR3/+s2/qXsPiLDRjuI5I5rHj2
1D1MAN18ZuHqBoJxVxBVHYSyp9/xIpXjZ0qs/PQqdW+5pCFxmIYBP2L+h28nutxK
rWbe4OpVzOjlk7pz/NpvVvffvxPNdSfiR1O05SMgo/aO2Dh3KMe0a3QoWMfS2eom
BFUtHT4RXpoH1xWzV3DOOT+ZrLQ7ZPC5f4TaNSHyQ64rOtfb6jWWopURBvB4ZQEF
7QjrIyQ/0IpeyyNYaM3Yfd+nmOw27WMXaP6xzVxPQJ5IGjSAu/6wIDIsZvVrcZYd
ZHwElEnDN8JjfXepY7HnyH+H19aKlXYauiykBiioZPrploJiOjh/pum86NlG8okh
whKXfa/k8b+QPKwzwtR1mmLfRIBLBHYxLCWRFIcI9pa5H6A3+Dc5D80IXIq0ESBQ
bNlu/c4lD8UT34vhjFKIZQr0ZQnQ4U5Fvxs3QvBjoM+zkdkfT7PKdYQtEH/VtSW/
deESMB8joxagvS8I6RM5TECHgxjU6T1zVJTy2z/LKrjqre35EdyFRliRbIpnyRCx
PtuICrawl8KJCwsKEhDrSSGX6NOZq4pHgtZ83KoRiFUFYbF/uKJrAR0Pv50eoLiS
Q9SyAl+/U4ls7J9vOCDNDzcqaHEWJu/Jbb1AuTP0zCPj/EcqNA1NMLWUCArqSJJZ
DyhL3ZkvmnF7kJxUTCEr5WcCIMurqEMUawjzNKKIXrI7Dca5LduB5gfL+5/UUsvw
AqgcEVSBLHkCKugP0dcPqdg5sfbqEGGBGe7+17SjR/gq/nv/h1+sCRJWbcKT0e2d
otaibPnUvxw0NMoGvM4I7nvNn/HYUAN6dsSrTqNN0/XBLyXo5zkV7/3YKcnSGK/Z
Hwqf608ocstSrO/DzMRAbGprxky+kIrXy7QWb8Ijzyyx1iYfhPDKSLuvEXSj94xt
/fQZTaIMaTS9+Jd9NCPgE/7WUGA6fb+j6I6qhZbG8NrpuUNkSrpmdJZOR5DaKSDT
ACiHNZx/W5Edu2NScDM6tW+LqNA6dQfDRascBpONaHtgM+NZ+doDkwcQIQ6Z0BHp
xqnIpTA0X+d9mL9r9/+drGjLKnRbYsPijt4cnTNp7mEjbDemj2hi7D9hKBSn8dEv
fZuTdk8FGmlzgjtow4kyq9XCv9/UpmMUU56r7AeerM1ORSYzMlBQzoWAMruYxe4y
nYwP0yclPYC+irJlG7btpZaIhU9gu289l2tIDZBzczddy/m41cZ+V5anhoVgox4R
H8MT/zViGMDhNRv9jD/da+egpU2+JnBeerRFftl+Ki7q6no1YJYB4y/42yRQcMLR
H6vnL+9tDuPiAoHLhcmjavW5R5zM894CpQsR08wriPnb4Dzvbx4BXRHvgpEU3YC6
DFZ90x2pEM0ElBCEHLBx+wecxJZGGJuN60dJ2WrSgi2MhJCXaIgGg6jSl7Fu4C/h
4uF/6LDtq0RyycmnmZc0oj9MZdPB67ICRq0jbdMZ/Oh9s/8rcEhi53321Lmhtqcf
6sPe60WI9rCk1aZSY5US+j4VhDfVKHGV+G8ZdeHfzxhtiZBp6WCm4g2R4PTYoLub
AntnIGnBAE5fa184MXYpKptH62lu0j/2SqqrO61roALgJlTZGjZmLZTAFdXeKTcX
OoVQFej5qy2uW4SczsXOOqLg7gGq16I8GlUqaYNcKNOnL0KN/p9WOgcIlY3qbsHr
hpzscQuUylghVxJ0mGfkyP4NyZEXvZVh0mZDc1sp/+SXmklms1kyCZn+alW8HQ3S
btODCLNgDKephN14sxa+PSmu7gG2bFBLMZothjIKrrSOC5epe2+TfOZBtNkdv1Hx
m+Bpc3vfaV5z0lM2jdL4lj1LYXSDsbA7cT53BLZgWfPXLvECBT0a2xV83e1zYbmN
pZGgjLqPjwPWQ1MQHxlKF/ZEbdGXCAbjQkc3Hzfk5ryWxiGTxGlmn//Zro+jF0DK
8rrdIc4fYIGoY0s31eBMTln7qcfOp9hI+vk7YFVQ6nSZhpHNvsgRAImqf2eKw2Qz
jZpxsmYQOWH6ifVZXCoH0BACtPxmJbbFp23wBJ4iWjX4FQ0UMsTnUxoTBg4sVwdk
t14ge5T1cecXLrtgBAoJz/SVXWagvIOIEBnD0HcjEevxKGpXKSKtooUGC1CvAv8S
omTc0AflGP18sgPKcV4Cx0UfmAjxauJFXrdsfO1MQ6tFaDLXLVgoDmuONor9A53g
MAq7sfi2vwKB957/B46FRMmn9+CCB03SkWRkwOUwNhKEuZE7F94ZiDH2wk8KyWzP
spc5yVCXfuDpyQaLPz18ryBQZjiKdDw37o2GHDy++TZ6y0cOJbfT2/ou/XaXBLfX
a70juJbc2Sk59G6nwO5/AFDiIp0XS5/DoNQUr2TH/KmJ5Gq12BWzzbE81ijNrGZp
r6Lk6UbxXXCqoeOdeVzvYaVnnN58MctfBQvo4ty3PEKdWd58GNpzBU9yPUTH3gUT
kLDRHZHkwabnuvBn2E6Zf23O1gfaWR1x1AxA9vyrRlYFpq9Z31MRfsOjpcRU0ArR
XfLlhX83op32PzK9BiGEIYNn4tLAd5UjGFKj+NTj/Hlb26TVjTeBXl141ehnGG3n
2n92twv/SWHgYk7/6NW8vgkNqeyKu9toVQW59AL7s8hcWKgvkVlSPR4Hj3ryFs70
8fOVsxUQGZPLuX/+qGh9t+4txqps39969pjvZB/t2DL0HTvP+4HdpTA4XAe4MfdX
AmKk4WaXsrsOmsnhQJ1gTn/NXwrjXPm2VrKOxbdNIZS3S7LE9VlVCkGNfusde4OH
LBb6shunqpcugKlturialVfzLxUhi6d6cp0KwBCdxlhy1g4h8bGUmtX9t5AKz5fp
sL3nkB9gIKReIvgL+6Ore1R0m5DdYPvS/PVkIl9+RPpdykrAx0K4phL6XAscRa9i
qx1R2N7erbJ+M3sDQtMjUi5sBDmD2r+xgUapcG1vbDWN2fk7u0Tbhj9Ttv77GDQf
ac4tPLIZ257VkEejJxOB7R/AnnAx3acMFagD6YpT9wMcKD4uOqdY92qxIMdvBZAS
vrpfT0U1yhwgMem/6iHmTtuOJyoIFQ+FyCOw/rtnyHSsClJIqDtItFwWY/Y6wL2N
NA/qokh8FBbG649NtDo0WrNOeD2cSIGlDzmkyXhVTjuUDaRcm8/l8IqjVi+R/A4O
wJiiLtXA/MRNRO0VK1fv4BOFXvkpGu4r4X8mqRn36YrtwoBgERmaENvzCAcrxNXg
I3klKj85HA5A5QtwwpcP/rYAos762pTlddx8RHKSQlWWnvfNoc820Bo267VZqk3N
q3QvGa4YKPzuuVTY4kOEt3p9e0Hve4XwHoSBRLRSWLX8OZ0ERnhk8MoROFQjFEvs
9xdogGJPPAalTm2dPJ4OsU5MLnYb0kD9CPnz9SDyNPFV0ODIQdmIFOolOulSNhQK
Glv+A/Fao/JSh1CbmODU+RdCAbZeSjtT1UiosrmxQH3EUQ0DtDM8iW6eqVvD1t/1
LR0ZTFGAV9spQ5L7r5opCEdO/RumezOHisaU7+ki1tAEIcyKRyuiF3FP1pntAla9
VEaGusf+Ioork6ig5mUjP/pIRgQULiH30ZZOZOnqBDA6FxkL8+TtanEiMkI5xKyR
j0kF/XxG4y2IwSt2YAeeDAljFWDeB7gnyH+kh6resGWNqFUBQ0XB7lpL6s7X06bA
vAl8QoBRdR6mGu2nffAe6z9FVWZDkyV6lOzho5hCbEv5b19waJJ4uw0XBL4RHYnJ
RaIkt6fom5LdejMF4WDZq6rSD/NA5+qf4PjWhcBrti54zlyjI0Vk4GlSVCxo5Q4y
oSdIRu7TNM/FETtHWmRKcFNHvNh9kcJph8VHJzQDSnAm+MFsmS+Lrknn8w8llxjw
4Rnt7vhHuOn+QYOd2ec2hV8zjvBzd3gXOUui++ZAC4u7wr45DAJfaQ4bRU1M6BfN
YUK0P5bhA/KqE90VV/uzUOsSDMwbqStc+qj7rkVdxvmC11T+dwMY8kXllOiTV2pW
l6Q4ULfQSbiJ0GXVbH0ZVJIzUmUlvbXRL25HmN1jtCOPGOp+UhyfETo3JTUG5HXt
q+BePaf8o+Ntqiy7bLwmkoBWE8V5ZA8FZ1u511Po+KCvVXK5IhUrZnbhhqQVd+hA
P5ZWz7F1opiRXG8TmbA/Fh2qPBJzYCs+lUo5aOGkjAJDQip5N2gHvNQvJJGZErLE
1BHYXptE4kcP/epXDqgQ1xxWgst7ffCds2tKsyWDMMoZIebbfW0Osv3mlPEMBqdw
oqtKxSzPGadfab8Vn+d3Ah/WZ4ktozSuFx0xjgfrNW0d7E8xWMnLRMxfQKd//VSn
ZeyXsM2ySb4TlLHRWz5PxPGpWSCnjSAqL2jy+8Q/kOTfrjxettcEhUoQyZI3B3OQ
B0E3ivPYsD9D/rdCXkchQEAfh+AWCQtlG0/zmWyk9J+q9j/4821ZXPYzqsvo9Lcy
AnkHjiQVftfBGyypqjQw6grE9SF8aB0yzZx9hXi9Sp6RAqxys/gVDXFDa2FztKI0
T0AlvzgxraYc7My6BBhfylNUi+MCco2z7XGbdRK87cALBHkVWoO+1TZc5GnhOgLk
XMBJQAhva3GJsmbnb2m5YxMxzPS9J2wpjS1fReHeHogN+W0Eaj7nuFDRNTeEt98O
dssld3pJRmS/I74+1FTeskR4Dmi3cCI02IjpLfvWIwNVJUyWIVMT2ww9xajIHsV1
bXoOQako51dTCDXDv5Cyn71qNJmNE7xbsvCLY0dk+9ObrbiKjzMjQCD1+v0PxxF+
arpM4YRRFYwT/++nqqE5v2dYKVdzLXc9QyFmHkdq4DgadZJaJ2W9CXJdWzzrN00H
xIGinbYks0JsGLeNruwlwv5rtHdLApDLaPZDTtMtzHemWXZfAqHlN2E1wnxFbjsp
tVGEJieyrCVBSGGSgKt2oQAaHa5gSUDZHaYQbUsfYWpPBlJTonln2zvwvyG+c4lI
eQSBXUEJFi02gG1YRQF1wT2eNS5uYkZI+6g9KnmFZ3yljODzn2Grzv8mR0/klwoE
/sBnsEMYcj6/2p5lOSI5oPj9oCn0Mh3QmzMPGyQfmQ5YGaP8HZt8oR0QXMb1apGm
9nlkcr2YAZm+CHPitp9ujGrxxafO1V1IoAoHSYm0VGtlDYdCaV7V7AAu3JRBvOpE
PP48EdEgkk1IqPphE/2YDlWh4jPc2kGsUKDdjZqCLVMhx6rAP1zi+7NdS4PWYS5D
GQzNcyiIEdat3UwMevVrYgh/gwy4j1An/v9GAhvhzNn6uwKqNXU/qHaIF8Vedh/N
ASEPsnI9bM2ldA1QFKjWd2d9GPPuk22fV6JX5jWImFjyc282FW3dol/HzwS31qRh
PKZsQEJb+YyjRMXZMlj+dDvteAwHnC5PNwRZyntN45Dv4ZtAtdbFGPjv403Q9QEV
t/UsrnPDfy5W5QfABQ1u+PLKRIfrAWme4YiLp6hX36y8FCaQZdCT3Lch5YfE+pH5
BuI9CgkQhXxH8gvhth6mz4tCDNCahyH1b7xarMp+p8Gz2h/9mB8WBa9g2yKJF5jh
wZhDmbR3faWsiPLHN0unixwk9/i5AFpGNRT6Pd/2wT4FasU4RtJTcn/3C2QAIboP
ZtHwchRP41r78dn7+/PZSIGKIZogdH4OXspQhl0eKpMBN7lE0NZuV4U53nUNm1rD
082z2FodKfWgzlTZs6ioQkJ1lfpwVZ+hum82YYjcJIri0oPz4LtHXX4nxOiqRCqy
0TDqQmSV03TEoioWboaUKkA//GyCgtSPx0eXuRTshngeMngJdaMRoChvB7wG98FS
lPuZnx/Lgt1ANaO6yiEwK25KqigJYCzZoDirFWFCIhORQsUmVInINHR3Yzb6/tfc
FzdcfvCknw7DBDZbYE23aO8IXJ1E9heyCaoo+eW+RIXIyPUZP/pOqBpEINGHO6FG
gmroyev5ivPT93GeiJ9TbwdOnR2LV8QLVGim4Ept7pwzkQnekbPT7GgMsNTzfCe6
/uktLDthz9iUzZ5ckqR11ZQplZU1kaw9jqTcdG4UrhP5L/dGGk6t39BkgKeorIsT
P/rXzFg9+PBsNzL3omgXgifKi+N2lsEXgl+5oZ8GJ9TcuCvJN389PoaBWm2q8mrs
IjL00n0lVCsZv77Ds9NoKXZYPaEEIrjAuU/znJEjUGcKkDGbPaoUIdXhyKktdbZW
C8IWjDVthY6C4WVUjW284vsh7JLWZTdXouAdJNU1U0+jhEKdpgxvAe9vLhpc5ECX
qC9rN1fF9/Ojv0+/0I4Xc90O8Naw7SxJFPcOJbNZJyaBssOY4K8egIy7ORp5ImUA
tYpT54HZ97kXfohYWsl4H+vRwBysZxykrjOjVHBTI/bIhTBAZpqFpXACx7jZQjTj
hKrxfAs1GsgxD4AdMNpRGULh7MeDzBEeplq0RorJysuLmJMudUT4nXmF9ETKf7dP
BYOq552TvvFb7Hyh/gm6o3qaXT1z5Z1kkXk8JIwAJhKS9iNWueFALgKHk7YPOt8/
x+qmBPxh4bLpM5AE6PQTVrN+O+rbx6bcUzrDFlelcTwx76r4u3aw+rk7wzcCYChz
DJ9qZTsu0JAVMDuvkBm8uUUacQVKjkxop1uuypscmHL8Xt2h8AhbBIdqQN67qSEh
qqTTmO32IEArpi2Jf//dL64zjp1d78U7hFE9ZTPII81T7UotussoTCWGMR962CJM
U+nz5mBm7mNxY8PjWgSLCCe0XTfPB20aI5ct79n0KTCA0KcDT3fAZ8PPHFXoDDJ6
sjweFOHzPpPnMroo/NdJr5zM/Xl7+JIAxTLq63E1AuG+e2B02i2LodOqTv4gnng+
p3Rkm3nN9tMh2DuAkKGy/zh8MujuA8k2sJ1SrIPbK+zGtpiHqCBc02TrmEeNDSjY
cx4MhBEqWpMYIYwoY0WPAiEJB3RU1hmQ/5cIc+C+tqCefrKrqfY+KRE723XT94pB
p3bcPpJiPBNcgVDId0aIWTXvJvS+OmTC8tp/ntDIs3xN0jcdRBdjtJUpvx7cgHX8
McBYF7esOVjJVaLSblLt8gYeFPKiKp+4N9rIK7WPMykAV0i17FkaWUxWDOnRIU5i
zZ2DBltl37X2FiSEECJnFW9fL+8tu5QVLasbQ1kLsv7B1W+NlK14lzuYSQf5ULbd
xPw8f8c+Wi46BZSm3a9HX3UX1Uc8rkxnFV+2kv+hTqWXWdJV0ISp2DGrL7rzIDra
sop7uQ/S9GS81rvYLc6NPbfRijpVPwYFgpJ91O3Quhg0cgU1iWvpcz3dGtgzalIw
hJBbnqP5x2olL/B2MAMbwHRDagLW4qC5njurriQTebufzgWw1CsSmA5IN+jLyGZF
q0xWg8Dfefmko1MFF05iuFlPeMTJx96Vyw65TkwXTY/LAQqGAa9GNipOzC4mdkx4
guYeo+jzRvCNsMa3vj1vw4dVJwXSwG4YFpBdKR2avzcUmcDKvxQVvW+JjJu/uN0k
g5Cszyl2XYrR16/sz77HO8XQSY9pkK8Oa5xzdBjmGQ1bZxmdJ8rxG34NpnAC6Zqv
9R+/1CZ/CUE/4wWgHmpAJpNebZWEhCte5cKLnL3k56SInNKfG+zK6aKj/mJPMsIJ
jdVUib+VUzvdccrmP8sfMCHskhZTq/akMc/+F+PUqhi8uEUaQjq0G1IyMtYcM9US
XujC9FaWNaeg4wZZTcG+vmsjYO+8trx+3dhgTN2B224NDoHNPg7DuPsQI8YtoX8u
ySsCBKyzFWAeuTGWJVsO0ZVrBsT+RQNi8tU8i5Qgncb+ySLaO4gDRieG9vm92/jS
uxGsSStGAnpq2Fu/w7gwJTXBZQpa68EWtSxtkI1lnNjL3Dac0DX0fpj+Pm8iMrT9
uG7jd4Dh1QaehHwJFqqTyplGaN2gykLu90DqtmfuCVgyAQwcfCwK2njORPrNU5wy
k07pWDk6AiKuz7YQkuGl+iTuDZY2AiKESfgI2OlOE/WZ+H1YJVw1nEs2cq62enHC
8JGc4Cyr9vdhKi+K22a11QFy2MTN6yagAqovQaPR2WSBZnmUh3YxcUUtiP4GjNPe
bkfzhyVx8yt4xNpksxEWNRWKsGU+eVn+A/eRhT5p58zV8sAfSJGT4gV0crkBISIv
eeV2dJFCqdubX8JpSfc7fbw+UnUjmpvhFQKPRgJcE195IYfz85JU5yZTWnwaNtrc
ehWfSCpyaZCcJexfwyDwI4YIyFoGYemWV4GocZfL3cTc0V6CSTsYY4BLOHwU6BQq
MxihrurlmUeQ0/Ds9YKNa4Y74wJEglWqwJmWn7/x+EhjS4elbCg6ZdjOotz9gAuj
08smVZol+gHl69SR259C2y8wbckTbERRwsnpTVDKHet672D9fhNJcwceHfk9lQct
xoD0GdSY73AL+r4GTCKJKK2ntiFWml921rk0vzIoYpE5WRwn6hvYdNvw9uPl3thY
ujqjac/tEx2pLH49Doyv5YcEPpKpaNaC7rtqZSUGMovnjmPfjrwPPMBAFLyKOPN9
eT78O/KTXgaXurELS6yCCLKr/ikPg9jFNB8Tbs91eMIRHIuzAK00RwG8E9nh1T3h
7/ypriWV+v1FO9W+ugkX/1emaoZUzNE8KPNO8v3l1MWQu9zt4wy4jWYZPFKaj1RX
1dySkI+NhvrjSpe50MeNWhS9KkVzKAq9iJgOYS9hsXM9nnm1qbg672D4o/Bo4nOS
qqNh3sX85ZJErm5libNi9xZEbJ4XRWUuIrvVSIqnuKM38yEMdZhFL4AUSwz1jqwc
IvHttU1X3wKMi+n0hW5AfLHTnC8dmE07Kfovkt9EAv3JrUvliiNSXGtGjqOHsXGP
KQp1w2StyrRMGpwAIm4+JRy5D3YywC4TSKAQwzythmq5MHgyAJNkLRJaXWzD3uwC
VbfXr+wFW6FX9X/4LaS3AtguHJiVqxjnBNRZMdkuAvdF96fKP3Ei3gGSO1Q59vWv
tTueC9Xj6duuc/c2OXH4Ma+dqBeWK8lm7M/WwKcZRhlyXWVOMez9/g01v43M5grZ
rWS30Jq4Lsd8DOmdYFI5aUFMZCCkCZDCsVE5xpsK26X+29QOyVopBQ0I92Xdc5Sy
P/AWE4yq601FIJzoDinHemqL8imtDEXbmjWv3B0zNTUknMQbYd1Z1IbAmYT4i2MX
BY0xLpKO6t2c4pUOXDXu2zGf7Dp8GI+RXxODcDR0IE0QAYmJ8yAsQAnq2QHxVSG6
Ph4sCGT6INiU8Oqei81LXaEQREl5c8u1qC/IZ/yzZylm3abiAMhkywzPFIU4RMfV
jIUO8R0ZfeVZHep/t+oNtzbX84OUceO0ppkGkp8+3nhROv2lfFWb/zWur479NYpp
piFnJY4wN9N6VFNt8xlk57lTRVm1TrdD+OSV7ammN+GR4Ii0+HWGUONgrWSZRUOe
pyS+8nK6zVxW2JzMldMqW1CLKO0b00P/5lCxCZXoAv32Efv4D1B1awcTB2D1OT3b
ufK9fxgHJ9ijHFbydBnYOKWsXS4YShDcD9VFbcjCL4YxkzA1Q1GGCk5JS7xCzWDi
QUkthUi/D6L11q7FyprTTRfJAVUVVooiVgOTAuz1I7QEx450gRBtpwWxv5eHIbMe
RF74Ie8E0LIRBctNezTprsudKeg2g5ldbrJ/JBTDVfWBFiuj2VNQm2AVE246R+PD
jqNRaq/2/RVcinuxX1G9aej09VMaxT1LO0thq2rIP7Ayqkl6/5ZPqgaxrXW1ZCod
zFU1JuEOwhJRQGo64wu79UHVlaVuLtW5Wfa7x3grwWiTGPVGDFEFohBax9q+dEuj
zA8u11LDB7fHKZAiM/jwvYL3LwUkHCLBrI5u2F2AM8u9TeV0+U0j9nWNVoOcTTfj
1UNuPLHLslJH9Oc4cosZugLRefGC550HOaH4Juog1uyW1FmXFDYdF0Put7SA1cpS
B3LSe6SN1TTtWd3jfLGmOL3p9FpRStMnlDNvl+0Sy9UyUfVsT9xOGVRSXwGriGAy
u0BkD/m19xjgM8B9Htxd695UN4r+JUzLhm7sRJ0quOod6snXYVkFbCQZYaHIExwO
PzUgyMWjl6PfJe/Gk6DPiXIr7tE6ITZbX+y3lhFIHmQ2wkLolkub0ATVGx+mlvam
CI6dgYLPMktpw4zs61+AEczFYcm2wnd8I2KkARpRsCZnAPd5dbMiGJ2en7MbmrqA
sLqUvMJRKoX7t/ZrUVGOR+3bje6MjbcKG6mV2skrKucBhymMi97biaP8kHIaJmOB
lkIOH7EwjA6UGSTYN7eIL6OP5n2L5xp7RT4VHhJcZbF7lKyaYRTXAp+AnBxw3Gok
GPqqV66u4WqjkQ02DtdfmFFNoEHfJAqYELhbJH9REymctWOYLuYegZ6Ou6ycWoye
R24Igfclr9ehft1ueG4iv4bkJ3EiWszRPonuZwcQssRQY7Hycu/I3y945PfcCzGu
Rompr6b+AXaGjHtZ39xxN/yzW2HA29T35W+JWKLiY77wy9L+bsbD4Jjq8yMBm657
BpnZJid8oqYi4NguLj2MfIqclK2jMVyxPg5Bvz0gzNqb/e+sRcDBIf60e5mZvFhA
VvKJR+0pkOWB0MwTkz4C7kg+PSiU5AxI0EEwnR91XMClA0tU9PhInWhbT5w/CyCg
7LsaaYm+8NF2uLJJ6VZJ7iZfHcFtUvOE8zYxpF9Chsge1P47rM0TXKeHOWIEY352
27pwlbZ9mjky0iI9f5ATD8WsRsmkD9LC9U2jyOnmztRjDHnZQcJ36cNhBBgeGTwi
EnkCRJaIiDiQAeZm5hji+Xbs0rRcbwsHO6NhgjGUy8eMFLz2NzV1PJcPyGpnvM8W
kP6MbqMWV0wzfBjbTYR07C10UAYcwufF8aNGXKayHsyVTZ4rd44e9mbvYkJ2NgjG
/hQ8dd8xucEm3Fc6sSZEwDE0G3xIz5jBvjdKzr6BMklDmXGoU8HQd9Z346v7yxkS
wtCpPUEKnzUpUSlEOE196xD62CLHIdbIwpH00e0yNSJpYAOJh6c3cM49Wug8pTJ0
dQ2xAOfkwZiYBLt78XCWQOPR6UHD67SYjZCxPy/tVEgLvHv1hlxNhvVss4ko3X7f
YReJV5iLn+Rmv1+adxDnjWujjUgfMcYRv1a0egIl1mI04/pgKM8Y5gVdNVbm/Ngp
nzxjVt7+chQ2eLDol9csWjwM5iNS18C/ssc1FEjLN9KCcotLD/gLnzlgqLvKPgqf
cN+7FYZ39dqow/ZbM/wP1A/pLtWDEwT1SIR+nvA+eSiUDgdS994HkjFKaQPGk4M6
qHrD7tGGYRsEZFFpJCproLGeoJvud5VdPg6pOwUcszrglTCfDrgchQRpcf7OPmoP
dzhcCT/YCcU8ppWwdJy7qP+Ee0ujebGwRUd5xW1cuvUgVrwPx52ZZqc5Csx0N5yQ
QX4gpUOfMPIeAns1qiRSDI4iBvM4FuQCDwHnwKz5EMKXMo5m7QLFxI/KDRXjvHh/
8ZUapMxD+8c4kLFPaICqoW27cf7+toY7vhNNA7qjcaKYYayultp0TmLxuADsi3vk
MiDsvsxU1Q8hLgk9o6sPUXpRNY11euehvsD0lXTXs0FpyytLM6lBpgw4J1mv5jox
r17jpYSMRP2kSe+BfkZtrYBM5nQznMw8neXxoSOcYpwfc9sdl7N6HN/tf0j9tWg9
GdNQx0s2absQQRCO9hTsaC9IkN0gP0lcWZ13DznMKaVmDdSWGfDL/GSyK2K9x7uu
FWtLe71w+yZ71GdpLg/AwCrY3LJz6NulcDoTpmjn7OX6XaJEYsozFrFNnox/M/JF
Z75jWqnZHTGs8/rOliTRcigjmF/bm9oOG4pnZ3XQRI//VD1f8MtTzdAy1HqN73Tk
ZdZETFCA5XDUwdpZJybcfgRQb7f025FsOkYjOR4QAy3pE4w88t5iWlxzH4HUsGoq
nyzX8ajg1UtTIW7/r+L/E0fT2JxXi99ocSqOrpVw3XcU1c7Nb1iVShpBXt9WFxMD
9C8FPAtAoR15Jv4rjp7dUVl2RPTP5p/CqjzQzQceWC677nAeV5WzCedsnxjfWW8c
LwPGLtQpw9YTRC2T//ezc7pdb3V+oy07wsgVCWcfbnKqFa2iyksOV5lb801CK118
bPOSi9lWQuyy7xVjfVccc3zRZI+05wAHaCQTHdW74BbtRJ5l2naC9P5tuntCbXe9
yMqP+h5pHXLWSu8GsLa3k9Y/kb9HQRM0u2i2BGxz/9Jyewz0RlNR5ArgbOXwgYLr
XmiZGkBtx2z2PGJsDRXDXY90eBgf8UeqGvMgpeXBVI7tmMF+HugEH81jp6GOWr84
hmJ5XBszRSgIyDnBn6+o9uAnR1CHm2EuWi3e0FhycPZMwFgcaIUfVdg8dGOE4p2y
obUMSpSQDq/oAO7DWzdfE4HH2wT0Sn9DGpHPb41fnABcFYEA71rAfTvGQ/gSzsrL
JcaRqYPDdmx7+5m9kl7wiW9ctdPy/tbtuaLGvocxjXgb7+uIMEbzH2FbLL/uGIbo
zPPGfvGjUGpbi//7/hEJhcrkWZoCRZZoWTmqmx0wgNrsy4W7AfZTY1hzbnbdKuHT
9vegTJj0bJqAhzaezv5iOUQsSqKsXW++kFPBaEg3s/RlheNLWjtkXHqOcDtpCt0i
Z1V21Wxx047YiPBPqx7Y0WEPWI7LmRgebgD6T67WQGxmqrALlZGeX48CvCBNPwuh
oFPRqyQwz1wziknNpYcHFURj2yRqYxvj/+kbHpZzR+zzEjKTKsBFeqGaykxfeAQE
GX7zIi1TjRSGdCAVuUSHunk/kkuHq2PKAzrpYk1f1WeDfqSNYuks2CoL8w1kiwhE
n0P91933VQoUk2EE1iq5Wv/Cq4aQNQot7K7QcQiTQ57WMS1VetQ3aAhCDffHVen9
QMMo2Jsz6qfG6IQ8AhbhcKYhoK5e3Ey8IfrCk1jf8l9GahXgvb5OtN28PBwfCkQb
DOQ39swhz1s08Zzw41P5rs8KF4rXDRxHK6qvw1a/1hzOkruZrJUWfw3O8mlVWG4V
rorQYZmhdnLx3HEarTZ2qYe9jnr44wj633XbN0zwuOloImMrEiw8+raulj+KpBgh
cjlbx2lB9SMSnuL/1/hFeJmikKUQxO4eUNiiR4AFVGJ5U9N/IQ3ODsoHPRkRuxi8
tqImFnH2/ROtqzH2FZXvW6NuLwayI4SK9DwxxR7hkJ7Afug+CG4rHD4rMznVvnEE
sE/DBBVKDWCFfq6GhRn/wwr+dur3z21rSKVAIF/tEATDFKzM3u5q7QtSjw3qcuIe
AkuTVal0ZG5GO9miheOxT861wDNjMNP7V5ewBT8uu5LkCj9fmS5UvL9Y1ZnySiVg
D4qdL2CvHZmCcljBZXPCfWU/KwfMOzyJ45JID2lC6xcRwPiJYXogbAi9pipzPxoA
JbiZKgGsO7UZFJpff3yzIf0wLBmwZNGEiUTfnat8TLSCEirFYOkdxzZYdLlICqku
NE9+zvxeRsqn6DS0bcAl+lw+ijlyqUPIp0OgWjpCgWfMlHjhR5vdLkiLILUDhiN2
IetngQa1fXPTF8gVzY+rphWg+76zcsAIbWBVbhsjLaq3Zw81R/6CnjI7wbDXoFJH
0ehxlNiXXtVu3Z8x6kkKdhbL0fSJPXsL/MDXeTF8AxJh2LbqvuHfL9T78bLQf8lo
9Wl+rHsMEcrmROBQe/+2uDvLTaplx2vO61zqxQS/iDLNdjGhwsjr8eapdf9uZcr1
8vOaXkZI/X3EjTzHWCC2u03s8BA9kyY15CJVgeqHC3hzOAtlv/eDbBL66ChTG5p9
QECxDvkMNwsFMFn9yLwLt+WB3tacOiObAvf8Zrkk9naIVlNvL5vPW2eavSH9c+eK
k48xdwLl9JmtRHGVylg4a0rQpXW/eESTUlaD9NVwbrUe2phjCg5C/AUanTxfOc1j
/f9y5JORBSGcWVr8N/uxGOGtPjJrLvyq8ux0IpU6dGMvP4EQ6Lwy0qV0hUstJqQ7
3TWC3x9EaLVd7xxx1mjwY+XO7H+P/p4437LMcfr+K4deAfH63Z8T9XTsrThu2kl7
S77AgTQyb/ljar5UGkpY54E9a5zIh9VyNuQcpwXLj9FPc+IpM8yXpBNxDiTnSg2J
qQXP3XaTZcFXGnIiK8Gaw4OKYCQXP1O+2YARez8Kj7k+bNXMTaygNI7//z5rtpgV
t55oUs2lChR9XCy9vQOAhWjIJCrFNVUHHiWTj55Z0pdPiB3wEBQV6e96jSaFxL0d
EBjcd5fZj8scTFA4uirJTtpEV/IctZe0y0czYInu8yq1ReCcuOXDeGlnXC8yPuUf
+IYcZFMoF95mZKIeVGGZ1i7JWFA/1rguUumJspyplY5xuDjvDp/tYMiaOm1TcuVo
LST2UfcZQJNwZClZwUL3g0jbPx+7ZxRyVlbWPM8xfOD81OUXnRl/frLKy3JEKjPU
+xe7z3mmcjzpGXGA2xclIwzrt56eyZY5el2UkvZhyEdqLawkYsmG5HgYQ1qcxsKT
z5+1WGYauBXWQZWXmbT2yTcHkHSb2D6GxAsn4Ll1wuWnDyplvVfDOsGUAx9xDpBG
z+sHr63JSNHQDKkeKHVfPvfduvvEOc+vrnJ156+vyo9IkWEdz/GX3ilMVyvG0r5U
dXdnwmWY7lXbTLfuStonccgA5FyDT9bTzI+/HnXPNpl4KRf07fMRlUBAEp+1mtkz
3REw+a9OX85448VaCQ8Miq/B2gbXAnEVd3P92vRZKEEvfW8O0fZQRUaUCsK2LEgh
ZR9mF5rDyf0I2MRRp1+QWlLlXNHDtoUAdo7X8wGrfE5v9bPKsTIFdunBfbbXhIfk
jHFuweHq8qHBubNmmV8cAmurPfRVOETKdT/70MoLT5qkLd5+G3ee9KE4AUH81ktJ
WgdsfV1EIGSbSzRkH2Ptl4sIlzukhIRqY48u6gHhWBG2gYaciF7y/rn9XVY1IqZU
wguten85S4amvZLOZEuAuC9BTIO4odDjZq6UMuHCho/AxQkDKYG9lryqgSkWqmFU
4CtrNVrqg9DywwEi3wa6/t5QRagPEFARqIirj7yI7/UM0KZ/hwdXp+5BAF8QzOFJ
IEzseKSDJOb4DJSy67tYV2BLjp60/phwSnCwcHGo8I8SkGsLL2eYEK9eqTYPkQqA
ToZ1C7jw+eRWy2aK1QHyZGBN1P8vx/txhi74s09MH7CRr9Ey3Uk5Wd2Iligz1IbX
14kcyeBzN3rP31gIw7hiKmz2yzkc5lnsiYgECYmyd8ebb2tWI2SBSW9ua3M2ceBn
xd4TDsWiz9DLGtoulgaLiU7BluidC227SKH0RZfZdhK3eankgZuBJ829UD9OfHwl
UY0lh5ERCvcCywWErHoMhARo51NMuIRwzPAhd2mbRVwcqvp4siSvJWenUDfnSKIc
aLuI4JF0L6rY270ou6gks2IHIgZMmhwdT5Nw9de5mxx9VzrKLQTrCuA61puDuPWC
EYdDhgKz7HEkUCM8r/WKkmociCCyO08gf9XtNGDCtUQ3o7KJyvWsgyrJS8d49tuE
mphriXZsp0vqOOOyDBulrAXBRpLGNQMLLop2cwRcn33PniYgM1/JXH1jdURNO8mp
H0MnLDLw7u5UkuqiO1ISETnh+IIk3GL68qcIUWUxwuwhEODp4jKlGR7/Y/qYhr2X
5tBaJZQob3NKePD9H/w9QWVBZUGrX0/XoZ1ZfmqiQvwcout4YcwXEu3hVZRyQlrT
biEo+h4cUj29fP70ThkioWAgjzxvDWkxhTLjWjG0n2QTSOshoHR9jH7xDezRcBVJ
iuMDtktjfhj3Za3DZcygTWwS7Ntf5MN8AkdHoxPo1HoN2zmXTX7JNNkRZSe45nTf
u6t7l/A2LH8hOkBJR67zxzyX7oQ5zhWj84GeDjV8BhCVm33gL8pk6SeK0GvWTidY
Q6qtL5L1ljsFCcFS1vfID7A2eEoIzkqMODqMk7wAeZBm7E6y4Gx0daz6F6HXn/cC
Fn61VngTYoDxIXSMIwZ5pneDuzTOXgVVH/nB/dHLeucqb8ziJXDe/XLuh/aYvJIP
ukxmW5MvhI/0zBqqPfqDsR1gJBcJ/lbjBbbxKPzmGS6IhzXNRQfoEBfykWli7tPA
xKBwYlvurL+IU/FbyoWFj3PYQ4/KnwTmS7pG5m3rGdjFJtMEgJmecHlOqGMQME6e
azu2U9lcBwDTfxsGlmJso9gymtWVVD3cF62mBYSsh7Tx7t2hUpJOstNJwtk8lvbK
huzucaGaYkqVoGA2vVGIrZr6NKnv5VfvZ/lGOAMyHeEz6db1BanUrgnCGgg5VHUi
QzJO0T7uxrHiyrO+5zvicjqwAhXKDGL1FJJhQ5eC9uR8hIHCql0Opz8isNeaIPCx
qXYsoDDhGTaXZQXi6PgC1kG9bg9KB6OISFT2TYTQfLHIzwJC30QG5tXEAhvehiSs
YQkxnuk+F4jYZoOJu0TYxuMxT12yuunCbhk711IjyipnrSAs3aR6njCa35TIxrmJ
nMj58jMwZ8NxS0aGaZihI2CVD23UAp18xp1Lme2rRxKxMGkmSCwT8xUk2nWUzfbo
fQsxzkM8vOWWudUB9MW3joG/KLt/6opC/1FUEEz8r3PLEG2/1ZE+gEFvRQ50gDY0
tPVpv/VY6YaUl66GECK1i4MbL7pedikAcXRnVvRjyFblkH7S14AulionMbzilGd6
Bd0uBYBI9Y/k0+rEhsZBYXab5jAxOEsqxY2/es1Pb8u9a9dm2Kv5nXI4RaEyRlBX
x47RcBnPuwJalJS8j5Jl+Vh7vcEDUp9PAuZ8AzhR/gsUz5zMhtMA7xRuVhvA2Jks
hUmSBNJKP0w/CioRuAVcAvOZDwKpW2M5zxsvuuOZ3HXF9d0sI3UKbessGH7AyH3d
K1D3z43XpZOSlbK18/dvxpNwVM/8hBMW92AHRhU0gFAMOgYw8TAQr/Ik9pxt3CB5
2I/wBq5As8sDjCU0j05ofUBcRIfsnv38NXyksg/uaqdlE78pAr4CDMXfKuGx4aXM
icgDfVFUxUCnx9ce07n1Dtp5pb7XbjUlqsnOVQwqONsZtMTmmQ0rpvWsupvF2RlW
xxC7aw6Ieatu8BZarVQGcauZk0bSM88yDpbidAv8pVfcHMmlCglfzNOGKai++Yxg
wwbZdfB13jt2MRZc804+/IowXb3p7/dSz17Xt/zECm4egFv7ATzpFCDoPRtaRBz+
AGEqDIV09wwa/d+u99aXEVVwWlRwB9/H75z3ApFlNSkziJJNKOEAaKsUmgrwm4G6
u1ufPspdeKTh4s5re26lCaEHMjSadrWoyjhFtFAI8TqhWkmzFZsp5aHbTO8E+Esf
ts36Q+0aSSmj5EH/HpPnZR5x2jSL/onwiO50AK2045A5laazBih6TFQ4+9a0iV9G
dspspLVUVeFh9ETaelFGS3QGaeHFnOdv7yAjPh+ICf7Vgn/tdnoS5SaRIsEthnnQ
Uo4e4surgxPqGLsUkyAA0n3hGv/vOrJk2vf6+gzeZzJ70mE8EaRdcp8zPO8p2/u7
nUfoAEkxPCIsBbeMG5arutmpJ1ACdBt04I40JH+XWQX9rMeRhCTJn7NMpOWU4WVb
roMszLHJl/n3YeKrgdCDv4pxUmIvTcv9yGnexX2gccwLdwO4pYtdaSjAqj/EivTf
c0Y6WK/r5aXvECbvyBzf7J8a//XwF90mMw+dQ8QGZDTcZiEuOiTUtoXC6NM07Fhl
bJYEWCzN/YrMZt2FdT2jVnR9kkOLvm6rc+YnAfyeDCj216vCWh4128DEv0T9YavA
TGBOe43V50dfFomWs7/NMMbzQReYNyPnoOsTrn9gSK2HoBuzSvaIerFv38FxQ2fQ
PAdrtzmKyP2zu1SGcTxvpY+mkCpntWRDBqcfWMwkILxfpg83w+nD5ms/rb0aHJZy
zqSNaQt3EOJNwQByRFs9djNdKy6Vq0q8s0yLTfgciqanUXoWi3l/LpSp2seyvCMZ
AaVcgwQkAZnPBNvVKSqXeouDlTWkenmvu43ryVxQMTiL2IeFJtA89X++vXs/EuAc
vpnI31NSH7FxLEc8urGA//tQ695+zcf16lx3gjeRiOAqo2TPwj98bbhEM6rqjiph
uoZq7bNPvnaWX4LVaavwIH+Zqke0feRTmes6fV4C9yV3xYhr7KXOEv0aV8Eu0Jd2
EL//kh8vvwcPRHOCHuDWGEGiCBWsvxRA9FVSmINkrekJjM+NYaBhh3gmilex0cf1
i8YWCKrBL+E50nrcClYZuWtzqauelyu4+U+Bs7Sn96x6POQX0+EdV0t7pZZNKZ9U
YWF8omCIibm/tWCCvWBF9Htwwhfux4gILuA6IUHKoKh6PNeZdE9nwL1NDJpvErKl
QItBrSx4gi3JN8nL5HIM96v/WDpZw49ztvTGg+03NWBQY343cJA441L3VqGtKB4e
L0JKDsLUPnhMsCdnM8soVQD7b+RRfizwVVAzC7Is7BxtkdA0RasL4gJWBgfk+M0D
Bc+1xSvYI7+7vcFE+ha6aDIiGRF1QvRXkmxzZX3n8FcYXXpL64xvIhDrrm0k6nq0
wupixmquk4KXgVxBs2luvh/HWL0mQrWt4klSu5Hlb28MWGlugDizMbqD/PFbUfS3
dT/isN3uGpDn9e2uffoeX2H9xL+QLSrcPn4BZikqSGBUj2rVjw2Qvo5tj6ziD/8I
92rh0NXUugIlSkit8NKxmvw/MGrSwkO8kmaT05znIViEqJZOV8wuGDmZmsuGP6ju
1k0W1B0YmoIekuk2o1fhNW9PITO8GTRqPrrDSGHrH6hIhTLqZlcTpsJrolULyTmN
moR93fg8LN1uUKy6u2UYXUgIGqH8LKaqpFig1iJ8Gj5IMPsoh19VUmW1EyWKYU9v
zqO5pDDwxRcpX9JUyKuT+6gV+Sk8d7nC2QuhyaSQXjcRnupsVTZqE4PC+QGiro6O
7cqYDMal0Pa/VA9V/tP9b+aWwcRKgFF9DhiO3FUeYZ0w9pXOxVtcEVDdrUxByjyy
34PV2VBlWjmHNtuZcIoBuGRrorOcDaTkLLsji81bi2TN8QmuUVkGugQot9v35nJw
m0UQKDpYiff1Gu8xPwb/Whb/OPJXuwyewxwLDXLLTSditPsG85OnsLUWwwCL40TU
vL2zQx9o7JhSd4wecEwUzJILSuEHLzH7d1DMOO8mv1nHFC7cWmurj24mys+XGL2G
FOzozIXsI7PNTuqUQjwdGehO4zlyHXgfrZy7MJnpYTipGVzq5069MrVDk3+Jo5WF
0lFDaB3jbWSMuz3TFy6xkDMc2QTiNZKmvfPWYmYyi9ei8Xcnde6nQMPRpymHOSAU
XMjhX/4SEVRbY0+JjEDPrh70JV/0/LanK/AyGs1RDHZYag4ZZp2w1W05A3Hr03jq
w4TbKPJ2HWuSMHNfimFl8lzCfMjg2WcYycoa+KBkauy/Rk65RzFDic8gz4pwHtLh
d7TRWnEa4BBJLSCBtvUTnkl9gzazfCI7YIuCEgwKB/csrrku8y69GdJcosfptEPl
icrohBQtQeBo2q8zCCKQ0NqLA5olqB/0C52b6SMx8l41TNAB6CpachcXKJ6/EwTh
MkcCEjBKJwqgagw3iIyNcgZ1WoEJ4fBQOGZ6a9J0OcG+enKmhZy++qFCe8Q9hscL
8Lw29/AJ+XIoG3RLGqNmja6CSmTLglDteIgYSlEeeT4CFvticzUlZ1g3uOUj0LOe
ZaX3qO+bzvOQQSL48or4wYAf64uwSBXbV2iti6WbijcBuxkV4y9PeSOdCfbavkA/
3SZnPl0FNdbUIDNvmhMQBa9Q0nRIoYFLK90D1tHz8eDjO5EhySHvqnpmD8HT3Wxk
vHOsr3TB1hlMdxGFmmUd1MsdiM22eXc0jlFWN+QR8G743V+DM+mLVjcozdk9D4bd
crTVnskcARCBVTZM+Bj+fhzWGC+WXKUtvkzF6Kp5zlL3sA0y0Hf+s6Dc0iROV2vb
l5eu/FHqq0mwAf/xleQpqp2mbHrwWZeiw5PS5g7+NcWmhxW3JdLI06giURWiPUAq
T58hurk//qJucK6RfEevKng2VVknOQKNqbn5P2JQ2uxBE2a6jF2WFEnlAen0v+9E
DGZ8SA2GYRcJPZnzbDftSgPcqHpjmbQEgMySWiaAQrpKlyDDVjIwMC5mHXDwOguZ
9fdpCfnkndmsupDqNoloq2De3lL1rXJWJYbwO979NcdwR0TRETmoYI3k+M0TUlA0
AcS/VWjM5cYSLPu+N/k6/ndacSX5M+KDbEzUo4Gwlb6pH9j+v6kAoOFsZYJfpSMH
OGjHz9g2yaeLI/X9L8QfTgUbEAkUEU02uNpJYbS1gE/a6FzWmuDVHzJKh+rMpYuQ
xFlPMmxRGyjzo82U0pu+vMH4G3NJh62PJlOnuO044HNejDdNthJj/hA6sUL9/SJX
NOjDp5XcZRMcdBJKYQRpflVIYNVMAvPMmhRfqPMabbwEFOTIqpD+x46dzyQso0gS
p0N+GyWeb2cgBElOnoRLDhGQblSzuMlfjXyi4Np5+LNokJB/O6DaB+Bs1qLaRFs0
Eh/igW7NUSHUCqXEqHH/XDMy48eew1mQJnPiZ8PqDD2PHJM94+UQY5o1DT23TJa9
CLHzKc14KS0kPQGL1OlaRBZs0vJGx6RHdV9VC1Q1k1SnHjJ/hE6BuCli/Eze+URp
AeFcNoUm/myghXKPpsGer7ZMxOfxX4oW8TXGyDjCVMTwzs5uqsUcxhH5jAPZpY5Z
XFgcbqFpcjun6P47NsAMTXE/me4P24nTjmoLD0f/Ugf84DSNYSbIvXFuuph+xbFg
B8hIuWC3uLwVd9gnTh/DLp/UP9mefboVA3kraMaGIkAKDU+eav+o05wLpimaWfWI
2Vip+kxUGwT92GAWaVD9ithEikATt5xd4BcfJz3LtdJH4/xIFHY6nKdOfvRM0dod
Vbq7Imtl76g4eaT45smDcMKxOvkEJo0sGWvDb+SJ6BGKRTjWHsPabD2ugoCQU4S8
XWZwGj1kVYEowRldW7qBZQgpkHMq5t5ptOqPko19LvemLts30iNrULz+SEmDvdSS
z+P8VQQu4F9hnzlvrFe6Q+bbBQIfMmM0JRky8W/YednXxNZ0JjsmBYy0gZRQvqEJ
gj0Y033BsRo80eDVRz+IU/UdaMneEDGAseq6B5pmTSpe3TaS0bC79UXjuPI8piO+
0LT0oo1WuhDYwW+q2ccDBh17K7MUiT/P61CsLcvkaNGWmLM/lR+nHd+2i9TOhSgX
NRnotf0NGyEPVpsD553pOTy3WQ14f8q6KMVF31q639u1ib5eY3AZulTTmNq9v9Pw
tlhFZRzPkArBOufaidTkNo0Ut2dEqk0/cSlkZp7HNfFeCTpb0f4zb7SHDmhDLXhb
G0CN1EV9aEc95+v6flNr6edYCLhT+62WkTziY21GWHuCnB6wiqwCkpuPcI47T3fa
D3Ur9ZMiLaN4RHXpo+gx0k6p1jAx4lO8ApKPVKZmiT3ZePQfJPRrZThM7J5dCtlr
sEkJBRWfzi7wkfdV3/JMcPDoMY5tN1cBnGZl5UU8Bcz3TQdH68+DflhmStJoeA+/
MVgre5soG9FSIBlvCpx+QoP9JS45rXufn9YvDRf0CvXfxhOCZMXl4+x69Y7M0kmY
408kCw1ztnuvqya18HhE//y5qxvX6o+mdfFgnMdeuTiNUY/JIDURPutTu5B6TZpN
PqgnyaYZKUpk4CewBkxyyNS60/+gY2MMBO6AzutB0F14kQtYpQmetByz4ISduYDR
1J+pD/umCMm4l192dU8KeNnM26TpYV4s27rlBXP5ZW9f/HsLiwYhO9jd0TJL/6dx
c5+1hK/dPkhkPJn92qAFmZe9fR4SODvz4W1syl20zVbk6lTTmNKemGbeOoCTbcAf
c5/882HbSHtE8/lpeGKPQHTOsdRtdaEtTxKZ8oHG0TMN21wQrfm42Vwbqs3OqJd9
Sz5jB4pBVWaA4D+UFyTAlvD0yhiWv/fN6ejlDuQda/8IpMOZqD1DB0o1WSHYYNe1
wuHv65PUm0naR7Koe56AK3knmfl0veErbghK10sZagnEZAzlT3LnSqk+1wAhGUhu
WaUnG5pH2I3XK0+pAdTOJbxinySOv1/8A8+XBJyf+ry3A9rnH7rgnmAjuEr1gye2
xjstPwCjlWOCKcks1AUb44qDOy1h9e8wd+agqsn9cr3GRPI/rgsrBBcZiHNKRNLp
7agYUTM25FzLAgKf0yHZMjO5oWkjrQM5MELcpGEkYWsdj5uuINUJ6Ds635H0YL8j
DZHOuVHuZNR2tSWh7uQVn9ftjTbBQwoyZ08wZ/DIFJ8dkQP3XEIHwN1qlAN1oZoC
+7gfYKlgZb5UELCE7Ppiny54ONC7sN92rDSuYDpSxQRM8qv7+X6mrV84FfHDICFH
2C1OX99tTbbBCN496Dpe++ElymlhMbH/9eUAQw5SOpROkyfHxPBWESYgDPTbTeAq
oTttgg6dX506qEJd4tClz82rACwe3JpkMJnDWD1OvGVvSz06YnF1LxbcPJ7ZfEy9
rdzEXU5yD55L/sKb+xtCcDy7m/hHPsxIj9J0ikM0jsSgpkGWE15KF5m+epxKsi6o
uxvsdP4giiwS04b/Otoohx5jG74f3y063+ll9gnOkhyLCutkvUs2i6I/Kt9w7C9r
GcFxlBAyr3u00ta9gtDlwsrJsDlOFtTyjE7GGiCRvfTvXwq8fdvKWkboHw3Q1h33
p0KELYaaG/n/gcIMHazqYXncd1oDoKS2GsywXHUr1Ip5xdVABE0zaBO+D/nr8+51
4+UQO7mS779NN6QDLkXZ/8rw79EwL/MXnqjSAhDZZ2ylunMdGPV4m36vPvOqgDEE
hQ06bSKoXaH7U57oW95V5aVLLOedQt+nddCP0Xaa2NJ8y7pCxMbLzW5sF+ZZz5Hp
z93HgB0ceKuleTrC1xwrvmW+KBAYImoGr445XCzW2EpNJzNfdVIuqzTlMmcTVeK8
i9hoLiAxNKFcMtu7fxQsNwerKDSKgp75M8KZCjZYY2gPgK4y5og4XtcW9S/tlZcw
wW/Dre5++UIYhkBg/23QGM3M12wF0oKC7Cyk5KytSsXo4OiAm4me5QTZc8csmZpv
ZXw0PpmQYTJP7c2qAsCVXYhJvRv1WBzYZIkv83ef9wsThHN32SnpVD1BbPRdLJfP
dnRbe4YAgGrwkVwngNzOKYCxas5WsOiZxBO1cTxdRFCa8PfqOqNNr8dHjsBKeHbS
tugsKeXsFB3eLt2l+jvq36+tiipokMFKPA0TMswbF1tf1L/S/39FJ/84OPl3X3x5
StFYF7q9D4F7yyKODfGeUe5cG+uNFjJZ4/TPgP5HdeRCckW7dT4+dfRTdYdwXdH5
lE3D95Q0kT7ttO99G6OxNroRaQkit0NBqbFcl6+4Szt/QcXuHxbv+u9le8RKXpmU
hYJlNbtPO/sKDe/tWZqQYcAQKoPDmBk7633psdHYVB9cIN4SgATapH1xlY2EcEkC
dy3sgw3Fka/hSJLsvJb/9h9exdrNnHPadoZv3WGaHzk/EIYR86vWZAs+8edMMe2H
RM5n5JG1Edu3vcFpefprV7BRDgYbFk+7ZnUkoTcvYqqeN09PQaUikkJ/D1Ds4qzp
X2JHhCr8mFwL9M10CU7yduSV5upUzrlE2CNf4/6nxAAvgMyd1t/ncS4DeZj822gO
pLpZzFnMh+lKGfZeLLkRSwgMCpC2WE99KkN7nAjg8KM/ilWJ1PUvFq2g93DRhckp
rWbJ6/mWIy5vOOurSBKP0+pMp5c0fzSwEb6rAODzzTiSNI6I6Beql59ozYWQr94z
2ipShQ2FO644gd7AjWJg6nQodbRhFkSo5tLxlBORkBMIr25GvMBcafgjB4nSkwWj
XZxCwc2qGERfqQrTAWAM3WmviOP0HApet+mvZ3GKciO1ltGsr1/O0TKfOtfTI+PB
Hhe32BtptYVVPiWW1dopwtzM15rPeq5ybjpO1sY5ujxuBg1hOYXkC4UuGO9jD/Mf
tLsyt59m7WsObcS8ueMgNTOGb3a4jNESYTfBpoX5kBdvhvXVTKqgThgckTtgedf9
9cqBUsu4Tp9UqmnkvBGxBWjiL1wCP94tu0Q0PV7Gi7YhMi/EgyuZFFuhLs53Y7uv
CsBMKPia9JanNv7wm1yfYcYVH3Bb8pap9h5Wq8oMjHXHoTPSNlgxiq8rNLtuO/Q3
obVxxcV34VBgiQIBqrfJjJZfQExVzhDX5A3PVkxYPuRrfCCmF+tKwPD9pcqKkJZI
wjC6raWaiwD+UpAQ0J1kPlpxzsSO3Wdmi0GIKNCPKASSMsqDRt0zuKNplKMiKT8E
V46vNoWzfeURnjauNBtkEGxCVmRyMkji17vwBaXgGEjme+oJ42xq6BmmLoPCuRmj
pABdVnJTEADfmAfMwUUTAlK2e7Z9FSuzwEhZZlWsPGkBK52aNM3yKz8eiO+uP1KS
3pbutmk31/DsVjKoaTh1I52M4ugMRsFdYnDeqKjp+ndL98X1cOTb6wTUqBbkqduQ
z7EFEUqeFwM7lAGEfPAn7qh/PfEvardJiavBF8TFgr1EOIOofAUacSP1PjRRAEkH
UvfHE9tfyUihaBXszF5QwuHi15eLPBME3jQzQP3f+eODlxZURgLU5gT87KxZ3Fav
iAS9UIoDthDIfHs+L1FFZO20tnVSvuc1lsX1QRqMgXy4wbrYlDHG3P4vvHaRUO2A
pJfpMTj9raYBjSdLW2tntqPlKm6XB1HEXJihTTPIPzk24eJFLr95bZ0ar9YIehGd
p8sdgHlXOvKxKqlLXViPVFkP2xpAr5BVxCfQMCCVViUkoF8TVL/ULfWtHZ7yGYRj
5XA5NRKVmF1f++1NecbNDMI51lmPZvj/lRAcTYtggcSqP7xbCCcDo1npQ/mY95ha
Z4n940mv5HWGbEktiS/B2WNO6/peCrovqlURrKoI/Hc3PEgOLN7/S7tcwS1CfUZI
taz+St6CWV5Oixy8rnqsqyqs4HzJC4vzHca/HxgxQyCulhsaKOI7K71OEYc1TfU1
6YagPYg1L1ByO73UHep4WniJWHIGFjkJmoYlF6w/hQ1r75I46sv9tfnCNpUsNvfJ
niLx1tJWY+sAju3FDfbsRsBW4ZLLts+Ebn9Bn2nrB9zq6vq4z7x8qynbNdtPietE
zu4sM9ZJWkrzYxro24TW8KRyGC8Yb5AYmKapcHHdKeRp9C5OhA/UhQdkE/vbNi3T
QXTn6HEK1VcF/bTm4IZ5f9Zl2s9WerboOvy7M0jweqLS2SQY8ZrDIXalQJ2T6FWj
GaaFngRNlWE2YK95A6qw87yxGwd1M6C/vWsV2Z5Mx0d8t6ghRg0qkE5hB/YruaUz
oTRn8DQakz8VC0T5qgy3zIrcgsahIUp8uK+JITc3NoH6UHKYFwe5sIgBQnvDHtxJ
q0qm2S0fGxgmclLh7ANJyecUfLRcYoEdqFwp4XuHDaTo9uz/tIlYgQ5AYHVYSCxg
I9q21iVyGwYUzwqJwbBIuiCT2lBlJMVNGcDwyUXLP93l/mG6KFhxZIztGlW94Q3j
yZ/7JIbfhjFsC8BjZAqGfnjmrvcumu3x0zLwXafXD/ZuhfqjWm/AQKR6TSEKFzNt
/d5MTl1GX0AOKUL4ni/KSuN0Z0Ieiaa3Vt8RjEF4eG4ibNtPtbskBCC+cFHv/FQ2
50IeRDclqrBhk9AUB0dbfqioh5ovRLO1qNaR6xIvuf1wA7mXYcaEDym1RbFxS+CN
PXgu3ITbAvrMkA0J0EzEFhXIx4P5kg89Ptz8eGx6iDxcF5yjPJaAqpdiFCVHR6Od
IrO2xFAjF1MtqKqV2yKJZMEdUQqDLFs5N5vv+/1t0FtxPcQ19lICL4cxlk+aILAb
wtq76G4vL744YeokjUdGiIwZEXtpQeRaaRckBJdvZBGdbjeYZt2tk8y/ZddAG9ug
TuPrcPxzEwF0OTlPABYeAY0TkQ5aaMnONMUG4e2FJqmFLLg1TIo4c90p0v093hYG
s6KGvLrSBPgOdfozmLMreN8dB/PaGJ6Gpw9pNeOEbYDC1iAUHxUOfsvbsTaFXi0o
gpVV447D6ypPyjgKH7HX0VL9oDFzvET2AqSmmn5Ja+GG0PHFkV7wdW6bHOkcwDHg
Em39tCpOa33jPfllMRbCUlgWizvVD/NMBnVk5xFGUubdxv2foVD6+/G5vypI6M0N
tFS8KCJmvHfquPMvR2M8gdAovgzsRSztbJKgzJVeU+LF9ei4/Pnygs/ncIkg01xD
jTFB9gFU8qZQHw3+a26rvgYqDW7i+8zlqJs5qPXDmUt2M6XL8m3XbWNVh8hxYQgS
vKsZIF/BVWmFPNTBixLcQaA5fjbLwrnMzZLet8EpgJEw64vWnq9SipbxP66JFQ4O
punzo93O1Df34CJcuW4SNWprWPdv8r7xZ1dGnKoedlHZg4gqk0vPf9YhK3SJ5hH7
OTq1DutbiWCkeamBX1nfLDsr+o4BNCiEMwfkPzc7HprJ2TLSoSTpAo+Ywzn95Una
epFgEpIGXS2Uvk3Bcsi+hv6OBqHtmFwiUS8f+d6cz8zyBXEOpbzPalhzCgK4H7DI
JSAuyWmQJRp2Am/P9LjPk8/Rg7ZpMpWkoGn2Mh41Cn5dljJOO3S3ahaejYgsXo6U
49phdSdvGDW6PqN5gQujGExFxLH7MeVmuwi9jmbUtAFIkf074sg7Bav3UE7KJrHJ
RXe2iuEld2aSWEOtSW2I1V8noTWhwSRZQbVV6V+k40yzqzE5rEZjAFVm4hgDVPiM
JKXsHm4tWpPVo2oMqfsOUwF2b9GbiAQfOUk+glTw5JPZ4FIlJzRsip1VHb0cAdwJ
zIJc/651tlcBMFB5CS7a92wE1CcSeJmxv0uvuBq/nr5qILYYOMKe3bbwrBhcSRFC
HqtenFOYamXv9JE3JyuXOmu4hwMcKi4I3ZYDG87N5qHW17uhQjEUnxuMCnPTZvuT
xsZTT0Op+jz/b0gmSEU6hi6dhU2rKifekd6FLYXpPzKd7RKCDL8shzZg3XmRMDWg
7YA4iwcXeryuIdv0PMDsKiM6gnNAxN0BhZ5ryJFYfnfzTE52gXsgOTKBSYVwHAd/
dGjidFf/mNjP1PTkRWOecqrlwGaQkAhEGCf3rIzUv0nOrlF0JgwzaKsxgRuGM3SV
EA7GaaVkOq7ZIcbrWxkPkR73j73+PhS6C/7886bDHEE6h4bLBI5T83AQ+7wnKl1y
owdY0gL3Ywjy5IyW3IDf8Dfs8dATbjszV1hCerw2oDKnacJVd8WvGOA4u97xLTNu
QW8LKMi8GPCakcDzea1n4CqF3KoDqbsTg25n3F+dPQEfnZgwio60JLE8tDU1m+Cs
YxuQGnBQ7CfXUd78xL58fKBoTvKqgR9lhlDfWebXJSZBngDjiY376bOpwZtrXGwH
QTtUVfjEGwwveAX+UEEeFu9Q9+fkWE1h2AqCebgANBsAs77E9t8a6hobwaHW+qaW
9haFUBmCAzCsbZFfbmeoQFXIR8doB3/TqXBxRhGs73FpLk+MjsYEfY0NS3bQhf3O
nTMNzDlRebJg0H16YFuHi/+eHldj7d5/CIC4uQnEUVTtYUCr12Jls+QTW34dWfEy
h3SRqkREVT1TDL9lmickX/cjLrDm830T9ZXp5h88ZDGD7v85N+itNiU2UFrzKjsM
ewxFrg4KbiCN0LLxjee8XFthSaye5xlPTINEeirPx2Nt5J7vGzQqd/YPmw1I/p3x
eiCeibndB0O1ebqc4FUmLsnBBqGjRLrP9t5geHiVnwM+SG42oBKrlXSfZD+qQIXZ
G9VKe7ccSpOCnhC4jmPTygUahOqAzmSNvZ/zBzFckfvxZ42stijYEIGBUs32lVJd
22fM1T76V/QQY4BOuVKE+KXR9JOL8AJzvCKzBvnT+Vdopu1ckss7FSYVZL0LCt2Q
QN20H58n0i6sdttFkwZ3LF4YuStkbf0aa81ODq5J0H7dOUtCzuIYX3EontoLpzF7
8zHduusIM0GLPbNKJPMKTfOo/KgUqpsuywQs7+pqgrzxT1iFn93JVwpc1nGpgT1Q
CgQ32VeqIMMeCK8UssqNy0OPQwpa7J8IRfsUWNNQZtFkkzEsiLAsjN60/kwiD4O8
LOiGz3vPc0DSASYumGrhwiY3Ra0sOrB6iHAd6WY2RW9mG1jhvBXP90KYEej4srIg
LB5rZAFHqSgXPTN8X2hFITYUdXUglr3qDCtlVUoI3uzmg5hMFvrOKgFYvhD6CHZv
/V4xEqUA84/98ypbqpg4I2FIHdbI9d8OoRm1mxWsEHZeZiFgA8kcyPk8nTF7/EFJ
N7DrqPv7yyWzRBz5vZl/vToQ2+xrE6z/wJmjKbQKhZ3fdmCHHGhXQCJI7V8f1CYl
aLmHCFuiWxkP7qKGnmtlkhetSg51pU/eoHai0vlebb+MGTT/9if/LuLSlJ2CRueh
avRVYv5wb0x/Z6aclc1Owa2oZScV0tMjQZFjwXndfWseMwEI+7ihmujwSP+9ljPM
DDo5/KyaNTpNNeD3ufyYKDiCLljcktaaz/NaxKMfPLH6mPaboprKOTqyzufEolcj
zHVdjBAFGBXFXmLCREM3mS+PnGKVEyD98JTuOrUFS11Bp4rf9UbxR/qEIkcViIfn
47Rd+OsupW7BT9uFdMFWQeX2peA+yl6bJuB73VwkRe5BEYTg46KlPV1pBtZW5JYK
GhrP+gPwN/YVriloqWfzWRf9sRbazYAlEjdaLYoPH3CWmWj6pmmETwbrVDICcnpZ
RCezoYq5pV4kdXaZ4NV03EKZLmV5Ux3WNdqNjK39/3nKU3NQJVVC4snwKBSds8Zr
jJNDwQwSK82+QtkUDZIyfkFTv3m1lPOX9ackCup7Kc+rBgMeyWR2l21df3rt9TWm
8e6x4uLy2Z7Q1gt6WM1lB2TQp9o8sBMBW+JaTz0s0MRpYkp7eYvnGpSumLoInGFH
9pcoOGbmqoD1RsBQBjoUH65pojfUIplAAr12jkzLbcUFzO3J892dx+32ciqyVwjr
Y6nOMZow2rxwMaAxLmrZtwg+oTe0j8nlWSs4avFlDEX+nfjA4rSNJKbGOBVrs5u/
8PUstIqWtIokJkvd/oFNMxRG0WRQwWq7zP/MO+KVDk4asKa+Gt0InTlyeAeQ96dp
jxcdesc0MLThUkhNB6rXGBTPoq/Pya653iYOD3xEL4dHVSM63fd0xqtpKH27JzLh
cz1X3h//g4P5LCV+Da4P70bm6tV1BKv1Ima+bxKtT7mLORCYafSCSsR/cpweWY5V
z0tm9qameX+i7/AYPJqC2WTGDNESjF1VGxJJPNSYayuHhmNLpJnT4cVvB0AGtvMR
Gtw6KacyXuu0n1Ng2tT8skH4Z5rzfkRhjkGY57MIVARNU2BU9jJe33TtvWeDGWN/
kaaqJe0oUhFKC1XdyD0S6DUoExWfqfm+GDYUtZAjlRO9xUrTPJ1Af/DI0Ece7LFg
4DjJliNX6+Tv8Ylzu8H2le969EowjBbFknXbw0+x9GOYxvhHNlECBhYjC5+QJVWm
Y0pbhpqqStGV2/tIXTJlqum2dZRwuVwo6XPBfhpATLKpgitFpkeXg2b2qEsTxNu4
1dW4cDnvxT9+qoPuNkwwZdD4belL4ClsbYtejaL7d7nHGQF0IG+iIgDeeV+yw3U3
WQeQMpPDXiAFVjo8c4IYJzYZrc+coCtlgnulifslDpVEeRiBePmD8ZTus+oyHpKP
twyvpgXhxT9xlKoOeSB60Vn1r4ntYmWlMpqQdsJ5jN2ATsTSIqivo020nN6w3eFj
Fi0OF2yjC43qmaW7S6BKJgpts/LNAyj1D47RCl77FzGHGFoujn4G213T9j6Mpiv4
Xg9cUwsHMODPxne/8lUy0eZk9T2ztwkwT+TEWgmZ/SGHDRh5pZEWao3nYOMg/Hch
C2uJ70p0ZiGjxVX/ibfrxfA9wTPblEiRsPoqcXxaF9sPF8Mt/CgA6VAh9wgVlN1S
6lce+Y6Iys5PIzK7ovzeN/0u/JcR25yFIuTEagOETVzAzRjeDqkaDd/nkVMbVTuq
ZxJucUaH9JysJQtCPiAy+qctNMd//uxinzcxWreHF5e6OxuDp0DklNB+Qn8C2XDV
re4B5ZpHoXh5dn7x6ssXGJ9CreFQQ2qZLgplSmN2AZ6+Bi+U4rGC0QO4MNWe7TGN
rA8lHOA1kPiY+k1bh5vjef1S4gZjhzJcSNElcRGvxv7HjkmMdFxyfFQKFyzQiN0I
IYWqZWNRnRtxqJCNjVKC7Uj3yPALEIzNBNX8ZLt7KuE4CLNxHlAC6K2elhCvR1Pv
bfeHLcw1DnEgSPhM7wXUXlY8nQJxc09bUxG9xWNMD0WsUFq5GvAFdm3jFPaIIFWh
7tCCkCXu4FxiHmf3C/4otn66EVYEc5FXUXWwX/WmtkPZWzyVWCycEvDhLwwWVAXr
1Q5hCVpSvV9fWeCOh3BowrpZUL4FiGvgDsLVjavoD7H/pAQL+gMcVqCQi1ZrqtvF
8C2+ht0itoCazKQnU+8jVxUJf9q6CgaVy9qpWkl4aFGyMZYsNCNs8zC0LlMM2Kc9
E9XSUMzADYG2NOKhEpJal0I2CvNHcwPOfGSEtnZ+sTFdJsmWxMFLK83tlUr1ziDg
w5r6ubGOGo8uokKrbuPjEKCPsG56WRE0fJonvWUq4n/xJiZGxJULiM76jrioMuFb
dndYur/qkM49Cb1bMCD3Rx5K/mGlR7KcOzn0rhHB68k/BMA1k7ch7/j0Z9b3psT/
7p/3VSIA+gOcQXnlKYpr7DX9jBbmPfzeUVBpH4/1UItQJ+zZWWrlvQ/f1Z37d7cM
rKOz2pMUw0zJiTJkwNRdlW+O7+hhVvX4lOM2xTDJ1A8SSV2XRb8u7B7o+MazfE6j
Y9yzruBo2DnXfLhu5djIMqNeaR1OYabjK/m+QpJEvEqTKIQ1wmE3ow1j0G2N7SkP
Hi9OQJPyqk3GhXXvgkfxMvdmyX3igaGowk/TFYOy9ii48HV53lrkhwVPrDyJnyQE
yal3763t5HBQbc6FhpVL05lNKPUypNdrneZiW0CBvcAgJnrO5GdjZt9PDIbskMtD
ppExP+KP7GDrC1E7Wqp38XnfbQZs824YpIdFe7bwkYQeaoO/Fdm8HgtRqiBj7DZT
M4UaYjFLkdg/J8ZrOvV78J3btyO7c8pGTdFe63GFUHa/dzJPutyaR8rkBYY0ljiD
zk1o0JiUgtgB4Tk5dGrqe3IvhvZjTCG9ZKE1dNEHWLe6CvChEvmdT+NXiGBFsyh1
TrDvzs0M4/+hf2vlXg9OMXnaM3G7XL7HgFb1ugn6xsOmNO/5PK61l0HvC+jYRqzg
jY/mm3UFoKXHs7anjYgzZu1XHFHJPalO5mjybUyWJ7HjOrAw0d96yUDNzDBnd+h0
3leOiC2/II+ioElO9zAPFgAuQQv7hCW0aul18Q6QNwIPX0XmZBqMmJ8LMHGmPiBA
YiYX2WBdB9cmSSYmY8nZUSyfkpcHns6STU7MZ8orkDieqiWbDyqeu08fBZCDUHIx
QjI9eLELzMx9XD+N0KPN2XvCohLCp6g/uwDDX6V+sKreyPbjIjgazJ0yCjjJ237+
ohq67Dxm7kjhAY6EK76nm51e8YDvKDv7al4kZ0VShWXIccr2GYvFx4BiRRVh12Mg
mDX2G5JGo4lotN5LkcOrGvbZGKf5g/ac3jD9woEfHkLAjcMl6fRSRlfbBHTFsFAf
uKvpvngXrrcsGLtbb29OIkPSHg7b7oh2sHBC1e7ES5rJMBydeQN+BBYHDRiOVHw6
RiIwmJh9KevWLkKeJxn/S+PJfTnNhOgUTezzcldY84u2FBqkvK0m+X3NOPdpjQ1C
aMzydYB2DMx+OAFen8sdQjdnx6ThdKj8dcXcJ/hbDdoUwuFFltbCykbVq6EpVDjT
jt1Nk1e6DJ7AJ1iLNvN3/ZY+PmQHT1cO5giWMdKUQMIvfBcm4TpWVF//kbWFDUpK
34v9JooJ0fNv8KFZyaeouGqUBs0P5nhaj0HGkinwvm+ME3/A6URYWZ0zcKvkY1/J
c4BLhZyP5ZdbMwWeWPCjCFhlg2nHoZp9dpMsHbPR54ACFtu9Gx81cJh3koxRaPvZ
PAKCMCU4urlaLmejDyZ4FypyhON0CfsG2YUgrnL8Xi99OD1ZVZU9aBpILMQAUMJm
pgD8JfgkNiTlZb9jkpT96867U1DdK1uEqEs48XHWtm9flgaNwuxoFkefvRozzeJd
aXzjQTPwAWUVWkLYBs3jHfgck6wlwIKIhgRgX9lOfopBS4Cxnf2Kh/toAJ0fnSb6
2oJByWANMMxDWFyrVg0zV1tqqN8YG3XmAlZmz1HO/4TgF703BDataAGUy4T+j9HY
nBdccOzRqTlr9k7RCXCrUODxfUkosw0YSTP5mE1/D1XuvRF8CDEUVnWtoMazH6yD
Fd31ZvW7vLJ+B2oamLqqi75VPWjKZH6G1FpXlKaTSuhvrLdQXr5rs/tq0J69WjwL
nRDCpbxKn+ZO4mbLSaKEKi1inuN9vYOBavYn/rTDOBiy8vkCp+KxdJ8jx63xgFSu
kKwM7bDLX35xTlqyMRXzHIUO0wQnrst/KlV6QY2mSP3rmGtatKSQy4oNUvm9SSCf
e1GRTk9lmWfUTry+RYu4LzukuOHROEKayXayF/pPn3niH6yIt9O+QobTYwC+1QnF
Kc1qneRWaCga7geeeaUOLXeX/xMhwsNSW7OFTiqwJiX2vKo4bqIxY5Q6uHJdJ5qY
W0qoEcbi3iN3sy9opxJklC2TLDk7c09gxsszfT76I9ZMTWJi6WZx5M3OEDyuUCb+
lgzlPu0seoG7sW30i0s7ruxwkh164kxHIJvMt8m55DnXe4FumiqVLEq6SPlMESXZ
EVokyza4R77SlLcouHUlZoAaC8f2/wCwlFdmzFoTMhktiHEcRvhkLJ9Ce6xH8p2W
TicFh4Wa2pAarcDywNlDISSBDXnqbFFSDRudWlOyj7klU5TmEIzZv+qdHfNsrKB+
EgmnLTpG1cTBQqxJJndgfyImWIitQ75cDn/fruW59QVSImUGWk9C+Mu9kelwNVBJ
F9ajKuh1MZrGD9uIwhULFtbavlI0wkUsI//uP7+5pm24lNNhPJcM3FMXlooRWLhM
je/Z0I8za3SvFZbmN7ertnRK65wMfHHmR5sVbClc8hCjhv/r7fMOLD/bB7lvS334
0HRJOUF0XUhz8UsKFXBSW0kXnD6F/38Dc0xynPdf5eWRw7K6Xvy3lmeIykev4l7N
HQYpNfBvqMVN3iznRbs/2vPk9AjJ6q4YtrQNbFfP4axrK6W/2YEgQ5nnn+ZIr1QU
AnbH3NGWsZb4TfQpKKsbEIHMT8c6Pv+7RqBUZ+b6TV+C8kpmpwpfn+E7ztjmQYNb
9nOAUOe7Vl5d0Rxb/DABjIH3NfYR52R/92sYPyCld8INmB0luCNp/ZCaVRFDctbs
niF8LoOfRAOQipdN2NO+VXwpLA2upNtauuhRdCwDAWwsAKoofmhBekyQisJXTwDc
F+JtcU5WINJXH+0D9qfTPasjNgnlGc005kvWU4u/8kmtyFtzN2pdGtR5d7vMq6KE
uhpUeRLag4imRBbjSpqFiEZWh7eD5gg2P9jaIDBwUw9xE0929oQKKRk7S3wvNezT
ib+BU91UmyAR509Pwi/7JPrjC54H0EvItcSh1Hr73ToGM5y0z5ZZ+jIdM+UuzWKV
5hHveHwuU++bEDsXr6YyuSha4UQ+d87inTV6/ha1kzNQEX3/5CteH9Dgah50yE0k
CJdrxSbf8l78MY7vh7zk+VBiBekGsUOYcsSgqI9TTZ7jDDOvCeTRz97MgcxyW1GX
aOvcV/E4DtaOW2aXwPqyzE8Rk0hyVPL4sx2Y+5R98VEZU6H3tsRRXSF/6BpguU9/
Wm/O3zGAjMMJwFrX91PHeCWLMnQ08GLewM30zhaH4Rj45aozTWOTTf5i91bYiXeM
mElmmX8Rcc1YZQX+63oFjYRrL4aUkpkBAdGse9IMTn1Xwy3y+ANi7T8h/UNmJltZ
yKxLMD9ekfxEYECd2AaDfroaadSUFS1JGCL8uwAOP/Ncym8fiAkP4hI0AIdjgHJB
MRDpDrmUjs8e/xHm9nNHhbK4/1yP4Wq+YoiduifSNvvEhs/wJhGM5RYBcz+h/pQg
zFrgE9Rs1lRsVkTeg7ljxChvaHyarHhVtHdhmquqUnSac/s9lerarvch8Vj87fp9
J8PCiTv70VNgO0eilWxdD9wSUN/j88v8M0CSgSn6I7Ps2IhgAf5jmX+JJtt5gUl5
IaDIpAx9xn81rKKDx5CpA1wt04M357ifB6pv1uZdLsd1Lh8q681QjFYxrL/5Rko2
PFSrLbzTDghCMt+e7uOlvt/1hGYbdE5x8jEgM4VA9ARzQ+heRsaWMJkOXAcEFQay
eoXSLVD9y78H1zvHxNOXt4KSkb1L56SbAvP6S5oFY9pPfkpEToGkiC7YJCrj5Igp
cjDjPAdx/yyySoT9ETml25QARswD6LubtBFjgN+tfWrMX8Po5IO1z7LfmKlbeXhD
eRW+hExqAzWl/ORoSkek2YVP3VzEhZ06TfIpe/gqL6BijDJjgfd+Hty0gsWoQNU2
1UNmLj8l5Wox/qeR6tsuGmqMtrUL0HZWqJusZ49FJ/Ja8lxW/ylZNEQ8BwwbQhzX
sua3d1RlmyHF/4kjGi5baOgDZqyhtOuCxrDXu2JVf9FR/mCia4c/yx3AA2j18lLd
+1YYC3d+Vl4oHMfEiCMjoagIXLxUP4rELPy/1kS25tQ3a//lKidxR18ti2aIuidT
MM7NLt5lVzoGiWACS+k5FGSVuScPRKFBOygmEGuZjcdAUBGzG2jKc47o9LdUGWbl
kLzo7GorRJfH/LIuxd0tSFWkQorTHWQanhJ30T6L7kWM+GH3VHm17Bdvt6lEJBoC
grqw4HvO2tYtFZSNGWslldnF3A2W+ncobq0LFiOAM5iQE6ZuQgGhLszWxZn9Mn26
6Po06YFHnk3v5I290FkqbYqQY3Lqtbcs8PJTyrzY+rvUQiGmquV8E2H+boDKlgek
gITYIaU+TWz71PU4JduAlOaAQCFk2ovBZrs3/JQxpXnurOgoD7/lbDdtordeICqG
DYnFJU9OBybNFElol0ysW8uYPA3S5SsewiYVzvlU9eY2MTaL89sRJCJk2XV+zgff
ObMZUatk7GfPm0BySOpum03sy3Vm/KZDrHA28Dn2xJomdeUbbLByu0NwKaowOb0M
mVKwRLO0d387fDswzvpg4HhQ8WeJfIg4ob0MEuqiXonqt0DuSyCK/mDHFHn/wzsY
kHqhzVFgoBwzzLpyZCOQfCxIOM1xFw88HftnHz0I6777cPvEb1SSw8QC/J240/AW
ihOyFrmF/iHGjn7WhXCAt1HcVvqU5yO4IK78hqcztCsHvN3MkhP0Gfeixl+x03PK
KgfXnb63YPzrPZuwrAJVqtm7r46WJbG8eOZRdkvuVRWMX2HimVNixMSqmPCsgiui
c6xButyVc/5rPA9YFxK/gcvuN3NRyahaIBndY5op/8tpCoBBXRcx0b3Vd7lEMnV4
/QNllTLkR6w2/bOmHYfYdXSSqlYDFLtP2wd5ubn1+pCSIXkqsaG93aaACajbrs6n
3P0t/R2oymS2DFeOhyGYB61Z4Xx4joqdxxsRrwQnXApTKxDJfQUKVelHW/ZkIqGA
soo/celBr8kPkUfKFgeX9OGsM/WVlfCfNTF4hZilGe9X7Jf6Prz7Kqv86NcckXRx
kqy6OYSXwQ3gEoUZ9TB2xPLOBAyAyi4U8uFhsCdZnLGBRSdIW970xM1s+0SQ3Wdw
jjbpeBfIWVT+qNjD9VJ7vmhafq5XuGCCXq4vZudXc3LhBwHMFejvwNMAn+ooBte+
vckYHet9k8mn1SEV+nFnzVGiRdUi9DuW/WDlo/E2aszr1eQHlAf5wwTr4LHf3lP9
+r3jQj61d+6ihrd1VD/QOygl6mN+HEdGVqOxz+rLFDWGEzrN2NceU1ZMI75KgRf0
MEaImdO0y5iEBmoKeAXLv1scX9GpDnY8NUcy70c4Skf1AalSrQy3a8/EpqBN4zOY
iw8yTNflcAMFgaSJfgkFKSqZKeEEMe7TIJ32w/JBPz0hkujQHEJBJAe2is6MgL6E
438shzbeIHZ8mDbTvg8QWLBnP9+6qqyAPc3Bxkl3ls4cEAb1TtALPaI/qKSQ7gfl
+09/14NjOHuthKbxWBhOtIi5l8DJ+ztZSPgogx7u+DL0QR800Gx+sIOrsGCF8Fpm
49W9dMem/ALP5jix7rMwLdJHQd9J3m6zrG2n2R8d3Ba0Z7440PZwgFvdPR6/CQGf
pGSo/WKIg0s/AnwIwLStAyvi4hSrh0Vs8gSX0ABOXx2urT/DRrbaC3lLkds8GWS7
bYNyawBwGsJEHHrbmGRu8ORJmWPMyYyVk1w3ybPbvUDyLLf164PvBJXk3wQ+cLah
mF2QN+Grz8/0JZT16oqY2m1HJafwiaYwDzd7yO/3G2o0c6uQHBZhoRXBZxRYXuD+
4rEmKuZvDvf45YKFMx85Mc0X+FeJBz7o/7D6bCoIYsud/a7GJZ4Wx+nCbwQb4PBG
zlMO1k7o5d/e3+ZVHKm8mWe0QUP9XnPNFcj0teAy4N3iQTkuKN6zrU6RPg0mBzqU
VLmMKEh7Q3Uu6hF+qYpgZy+uE5PgKiNaH8kKg3m7cM4/QGvXTG9OfDDACavaDI/A
WF4Pcb4hSH2J6AmRKjxZ4R8Eng2bDmG8Vl+Ugj9rWbOgi8eGlrFJbAWETGqAOZYF
0hk5u6xGTvu1oh64sh+phsRIPYBIbZer2635r/0XZXNgu0opBJotzD4Fu6NmWVal
hyeeuuPijIxzIWDQYi6m5yEEmoBL6DUa3931oqToZS+7ck7Z9hriCaf+2v6vJ3xm
KhgjkXkWimKlF3TU8qJj0JU2hxnPybzwU1bg9AnsAx0dpop1bLvdZ/1SsnOBMPM0
o/VS8gThDdgXP4IPO2FT1+r6tpe9YLacIbeZYlOAE8FcRydYjS749PXq0+0zI7Q8
I3l56zaEYqBnRjJA/8QBnYttdalOOFoqcVZMgqhlMrJ0agObzL/yQVn+RkA0ngRf
myqTlI0qPJj5OHZmYuwbQMInvTpspjK7peZFjJuyLEyycLVVHQBIV2kVCfJLX3aW
ur7L5pdvpCSTARZSfXi7SVoCPjwra8ylTySrp0hKyqCMjRLuw0XNzBpZXoLRUYk9
Sv0k3Ym2gTyBVju80cuaYqdonrOxdxY1f3+f3enVeIXpro/zhHkg/vto0D1zBimR
zMA3df5VUtXvK0+Adt02Re2CihBhHU/S6e2gyAPiyrD86MDAyXEwpgmIVqgvTmTX
gqnegBnL9gJ71Kh+GNjnnTjeViKKnnVpwdq65KcnX5UpPLvr9Jyf4FuGAatXXL6o
C8VX76eGILmedOIPYvWnc4rfWU11+SKs5swrlULIkOQ7ufjWJjtwWlpN+8/P8rqe
GQtetmdBX32bS7gxHW8NWuut+dL/JgCsTp5s/NMwPU5ZVcYvJGBBZ3dUF1e1Pkqn
woHLK8zVI9X73o0WkCP3mG3OryNIcDOpuf2/Exumaa9lvP4trjnIA/Qu1EskzK+U
Kc6IhS1B7dJZWGAsTgpelUrRUDQcfyZkM9ILLaS3fmAJjmnflwhS1Z69Ff+ay37E
un13JAKAXMhi98J5Yw0vzSSjrZ4EQoui6euan0mPqBrVpxG9DXQWjaMG0ZPvAgdx
bf7pBdbQNwf6PptkICvcx3AJMjRg6Kr3YUiWbzoUybYdkW5pK/8fmPBb7sTU/ey2
WUc9BQJTl8HWL4J0q3YspFcGiVNz0fIzKC9NKHrfqUR5Zo8UO/MO7nKXKlxccZVb
oJJWuAYJi+J6tP4ap5Nq9UUqESskJ7ChI5Upbz1rYqCFFOf/sAQuQ3wM5v+jjfgF
Da4NwHGK6/RYIHiOlkiXdM3wOwe+a4bG+raWri+p35dBLEorDxRafiH75slz9STj
J6dL9dRwSQ5P7xxt3fg5duR+UBkAi7KBACW6BRNddj42c68uDOSbqijdt/NSkt4D
OG+Px0u1xG1yDt6CP47wiPYdT8FwydfEokKMmNu7KqrQ6RtDnQuMRV3Sj2vDYmWV
+Xdf2MTItsWEed9ZKo8f8c0fZNPzMqmf313uKMeN44L6PPT6+VNlyUeu0/ksNQyP
SQs/mA5qOfw//4Jfew0S3s5zeEhTlHHVII/qjy9O/V8Y/7A3AGgMcGPpbznTEBAW
jXBLEr0f6FkK4JNw6HiljoMcpLbrUezcGQo4mFkGyzcKpHnV4ZCE3YKVR9woZUhD
rmAKJUrGz8b1bfzQh59x6fcopNb//wSuN5r//wzgwyrgHiLzx3YpVB148mALyJFa
PSYqt0sKsovnH5a4QCch2aQrUCaQWNIv8lqLgV+gELnAfAVgTXWDEY5t3t7vKgCm
f/lrztR+56KeBV/p7wJ2jk13L9BkyqWCbQge/zQXQCzaes2JoibFbLdoeoPTapjy
5x6pI9S5l8UQ3Zg1s5pQuz0ek8C3alvNaDI8ge0Y6NfEuumvuQiMrZQvPavycOD5
dfLPXgDsPpMI93u683Phu2poqvBAAFlvZ9qFr7E0LKk8By6Wt26frypHpAy19T1h
G9Rmv/9dC/Ou6OWsbsgSdRq1beOuB4gVAaJlyOzN7xJ9JTnPuXiqdIc9RVUV25p9
2EOUb9ra6P9MI41AYDbT54tZWDVXpJOSKxwouq6+k2G4aihyfJeguseCpH1RL1ra
kAlaJmwvU6D7XdLJFdhNVvZf/WZAllsnzyP2Da6QUaJBHeERlsSvnUioyQdpLVqu
kNIfWldwD9yxeVUd0ieF1knsCvznqvwKYDC7DSt671n9pk+SahLFmAzyvnYFAX/p
N9nLh6+u2CEnag73RmeWtyj7ebUQ7UKSmaFI4E5NV0mpy3LQ40YxFpIzxvdEvgpT
wImcGDWs7aHryCXWlWJcBRprr2JZ807JD6YoV6VchMN6f2AMlSkxuzdUOpPD3e1w
nfbMS4AISoHWaWKePGLyUNniJ30/01YNW5a71ZhjoZiCeYRz2R2DElkS0hglBE9E
AYIyNWWlUAqg9KMop2C+7qK2qA3WzzCXuu++O2WKXfYo9GNlDcrcr2BzokSbNgTa
ODD2My38gsr5joEQCm+a0zjEc6ODWvJPchliJZakuGe8+sQpVyEa55AeZuxeEoqk
ei6Zfz9ZUea2PO7/5BTgVXo1enF2TSwCA1kuu17Lh5ROzAOOifiFIm0rhiENoE8D
CP/qgV5e5JKjoqatlvywoTDmiI8VeqF/GcXusnjP51CocYF52d9IODOhO1FruEUc
0OeiwRmVs5+iLWrYWdagEuHGdbEyDrqNb06cee+jritDMnmSdXXMFsKITMbFqHDT
af8Sp19D4CbMLSomHmWplGw1B1zfetyLG6b/NfupCE054WoVUnu9UNkF0i7cxkn+
RFKIoDdXN2esRdDch+hy5SAkAg6yZHbbZVcNmJibUI3XXyZxIge5PHJaGFOx2s5T
DNX4uXYhNUfk5UlIIXhE681T9/Td8QfL81mYT5GDBRJj9N2D52nIkbMWzwxN+iG4
duFQh3KOUWOC2rekMGSfGLUQlqONVzf/1HFeSKrD6KQEeEWcqzTNRs3PX4ZUqE4l
n3uv3uGrh5azUd+Ih87pXhNR0ESP2vpE51RaX9DsK7ycytDJl1SeEQnkQqAoN2mt
WBbbFkBGqLewFdtqVMfE4h4koqoFophU+vRKd6tbi+qMRhjOIWDTtRZcgl02JXkf
FtT5M+QWIPwjYrbuhv1RCk1UK07ABdmIiwD8qka6z9uBFvIgNOSmZaVrPEg+qjhB
SUtwhvcCT8lZp9qBymOphcQXfqg/hlekstzwhm/k1+t0EdB4PEZt+N/TLW5qbkP3
TrxjgE1Eu/2lAw2fAgRXYbe2nC6ZxjuunITfvznGjvK+D2S81XzuNEjoyFrnky7S
M4S7UVmeMSkz4xkbrTWB745x47css8KGpFwVIey1H16p+2nqjmB5GP1u3JV+nkTY
YKQcs25cQa2YScwaUXM+bEZnFOp9/IqYJlsLsfQHlQiac+RuG/uj3x5RK97Bh7ZK
lbTIT4NlUAO6fIPRlmqYGZDT2ffiX0zu9i6CQ9vrWH5FMrjYe8CYRgYnbAEVuVJI
1z/1aLHm594ZNKONRwVWe9AT6TjgSXx6T12sDu8ZlrQiaXf61asnzXeo4ekFUuq8
Pcu5tSuPoSBXtrPBFTnlAMMZVxX3VZpWRwSC8VIKBG8R82hXgOQPABSdSMCAHQ3C
StAyMC5sRMdIwSI9UbG8VTyhhNikZpt+xgrZMMrt2LpBHX4jgXgryo2i7ANL/0Yo
zgYIrOJUrxD4svcisZMeJ1AEuDTB691PjU162ja360vROxQiARJtvel41tL0YIUQ
Yh4DX0SuMmUod7Cn65OP4qV2j4L3DajCTub1sa6aTRJDBgxmU8+tl1/v/T6SfvPi
oHVMMLgS39cAFTaBtC2XofeMiVRseAXc3SfX6y96w0iPFqk6Lnqd43n+xsvtf0+H
wyv3c+x/6f14qip2LRDSL4NswyUxGrtfAX02E34Tt0DzIxBpH3eeovGBUuQmxwin
klOQlIt0LAHU4IzHNwjcPukFhA+XdWCpPWncjKh7RdXgsDZ33Xe/RvqqqXa93wAH
CjxFIUiLPV22McO2not0sJxSts+ZAdmJowl1tRj+LHQ1Xy6nm/qRf4BoGNs3XNFh
eyH136l1weNQHeP9sdkB9DzEv6DX6cCvX1FwIKQN8LRlAVlX2vd1En9/dx+eFVsH
OqaKEB3LUvqTBmf9CqVmBf2zaYvx24xn3vSMe5uLKyHC4k4CuJHrn8F0ty7NxfsQ
pa9df0wzlunKN82GgH3dE3utuPVhfRmGK3UMvutkdxRr4crRiFVoh+/93vG8kPUZ
YqC6xY2EmzqPOBD6vEzjp/E4fI8zvOWaFIKyf26fwBgh5pWZWxRYcvljs2/VysTS
l+jV5ij2Dz9CgosCJC5sbdFBcK9EiGmMAK0Kl4u4VYA+JrWMrMueSmLPYTmxfKy1
sZy17PWwNhCz6YWG8RCegi3xsGbEPIVFAyhdIw+CrKgOVI92iZXiaZuODFTzXH6R
zshmVqyqojOUQS2gFfuxKqt5ApWhB8SPWflqfJV7NhLxCPQOFCSIMqY9XO0vD6at
EkotY1hYbunzF+a+Ztc5RuK5exNuJRRunxfIjeVE+TS3nv58f55uQ5hvPO2KuOG6
Sg64erYGZZChB26D+dXGvTaHwa5XMBwLeU79/vAndLI+n7wf3MXmJkCMHz4LpmAN
wY9Brkubdn5wi190/pHVDG3EdVopn2Oi7427i+MDmRV9Bg3aboOsKuDJG3gcjjN6
9RmY7nKw2m/xDb970ogI1DgkVxKR6NHVSaon8lrs1VC9jBmVjyv48/0FitIjE9D3
sfur+fO/rOSHN7Dli/hK9U/H+EcQAIzqPSoWzXu7bgEHoIqd549Wa84LgUPu6gfs
vlhKfb7nRVJHvF6dXnCRAF9d9OT2P1JOzBs/uxpmeSCeUCX11+nWTg9wNx2E6Nj3
haW5fxt+ns2oe4ACUvft6StiqnUHpqxMQ1ASjKNsfCCvWHXaDw4Mqb45TX0qwYxY
6UrKFca8u2xB4BckR7ln3YB8ic1ZLIQQlJ8RY/DNAghhz0N1wzyf5kVgCdJAVX8+
e4eD4bARLMkdkFbiT3qiTsl60oxKVM8gykX5P4XYodSQPBJHSNzgqpDgQI9+5oG+
yespV7yEnkXqzfvukz6sK6YoXctbngxy6fOk8qAigkkZxeEOSY15aJ9+thKLcp9C
o5vifnhCuTbkDQg/gUw5i+J5JW/hLib6t+RggXIIFCWN3s8Z7OC5wZLLp5pKt3mN
05ux7tUuDZJmPuboG72MCUmiq56htVcqVE861abQZyxwZO2Yu2mhTK7+svRFVos2
6f6kjYGo6PAU38GHCdOS5X4f38qpvLT1ZdfL0BtMY+iol3Y4jvVi42da6NH3C+PR
HxOFr4jlRGUF+2LIUOFbs8nB9rhrwhmQFBpAMIfC6KWoUfiQY7NutHumM9BoHZmN
/f9qXeGAm64kCbDq6UwBlayUdlXREMDPw5XqYRw+/MzL/0suo7MVj3OezrSNzMau
WfkqqDvgZ+mdBsMBA6dgRqVGqu+P1Il84UTzjmmXQeXofmBaFhTd2CqPvKGSthvD
3RIAj2u9/CiwreNsr7FGqnV2hjywuL2X5Sw15K6FKwjMVId+AnzPRei4EgFd41Pm
PkQuLQ+SjM4FJcc3pKjIgNYdsxw98XvP2WnLcHSQbIhK4y7k3L8qESSZhoFliQ8G
G4CgPKPgpNIVr+uxNuF3VwNUjcjlgVm9jEIawiOcTtGGp6GvdDx9mcGUJersczbp
BTh3UO8+I3Dy5wILL2MyDcIGWlsaWVAV3fthWoCnE42hRKdejD1bg7pJ1oMf+pAj
7vVpBIbqyoyybdZTuuOsd/Y6AA97CDjx31p0rTzq1+Tpxj7VZ69Ir/eFRE1KGuvE
YsW2SJLBsxLeyLJPxLxxxXyNy4EF/LuIsKROZtU5SJXpFWpciB4P9t0Ufa7HhEe/
zLGB2iBI4PjFXw46o5urrkAO00nBfmPbsBDK+CY0rafZzqE1lqGNw+lPWvgjCzGR
jcsIhW0hudkkdiLOGmg16IqEDVSXrRm+Q45x60CynPpXNB5AMgZNmu9YqH+sz3lX
7MY1FY5UKzPMK5iM2wJk/zvnMVhLjR2x+9jM8nzzs5ivQqOmZX/AP0M7dKge/ZhD
vC4aLn8pqbYWLCLm0PO7NRVKdpflj36lTxzhL74pWbBOo4kTGLIC6quPNsBcaS5t
0u7ApQmVlxcj8SdM5vCKZ1o+UIuwczmEpTL9w8ZPRnIdMVfP5/BYjzyuuyyhrfGB
bISHNNWMXd3cdgFBMIHrkanUr9ZztmxG0cnUBIhFf5QSh5bAN7ogO1l16og/9OqQ
mvlFwAPA97FgUGNaSNcQJeG6hZAFAk0zfJ3sL43tL07eS19Jq6ngCij66gZlgLA9
eiJq2lJ0rYTc+uXJPAonVjqP+olh3IhCUulmUuuideCne9xxjhpI395QHdMEJWbH
43Pq29A+dtUwkyQaic6d8x2/LHr/Xb+tA5t7lkAn3np+42EXu1Cqsuzj2UJVEY4G
0VskRolKmsSFoVSh4zKxVtVORBburTXB/pC1WF22bVBFXApknSOGNb94I9ccL8lD
zkrWFq8gQEMpHsiHKtVp/xuM2Ip0VokxJTN45VZGVS4eY6tR6h/B/C59yAx1DV7J
ekyFUMjhRycvuSVtqGdXSVjjsJLepbm9/BI31V3c+fx0mjo0DUseFq2+2QyAyXxf
mfpITlQcuc7ISeKDeeTRSptS4qlYSq29jBrG2o8CzLRPqzG2VGJAu4w6MCssFisq
S0o1pAJQTUouaqwBV950HTSIJur9Czbjo/saRgoObbiOEOx8kyQlZTp++bB+HbpR
7iagIQM99FcVcsXQGQRjDSjbpB7cznMpbomL7ybf2qEXgfI7qzacGe1q7WR2Wk4A
0iweYVQI2OtMJHi+Eb39sLWcyILIx9MYA4AKqQ8OM+htQu6mm3fxKiYoGUpwOjBY
/fAoGB8EH2UNyHzOJ2hKzn6xcymN3+5tEvjwqY91jAGAizLU80RRyS7nRhXI539W
1cdg00y5v97pLTzTog0IBzMazM7BRGffIDDwq5fjayziC7WgmrRYA7iFwF8tqfzd
zRDHYiEVtRzErrSa1A/5Es4IuSdhRnSzqq8S8rn4VJJ46Hp/81r/jbVDaxHcTx3J
dWKiGVHimKxBi5VxbCmb0A5YhbMYVsVvr4y1+Dvtyfa0vCmKwohBfBJJ1vny+U31
QLUc4DHqJCQIy3Q8D4JTiARWUQw37QbV46yniBSO/FripYLRONv/DBCeT5mTnue2
TUMgADP5r5tQ9JLkLX/nfezwGn7BtKvrVDZOGzSivdbF0NR8X7WvEVbvLCyt6ELv
3jidhTdKqV8QZTPnw4hmcWElVJogD/M+p4SEp6B/eD5n1dld8wK8XhQWydbqBlob
4R/WvTjEBB/o0+Q2s2sPkNoEF/Ix+oTo4RQE/ZRcAPvMFbvXP8PQD2l3YCiq1/9K
zFktljmkLCpKuX4P+KvOJ/rpMQFynm6Jl6AOIvJCcKcQH/gBKfBL5EuIdEfQuENx
8Hgzvn2Asum4L4Cfnysvv4ANiX1ChihUQ6/hGZgz3e0K8b8VXuUiQjU8nqtdndyt
MAUZqdxnvunpj/is75vwAmrFRbSsIBfv0eg8Gq2y9pyiSzgM4Drr5TwpeeVQjJmF
FOAGnDfNSQ/I2OgKvml3WveYlq+XKgEiVAPPYNFLMDHRuktTXW07mVZ4dfozBHcD
4aNyLg2jbMEGG39cS2R5LEt5u44m8693jzAwkEKpyk++Zm4TjMh2tsXEzuvDDhV0
42H8r32RXjQ1I4gg51Q8MmQX29bwTiIGJORae5VMjgCXo17vbDIOEELoLE+GmZNW
AQRLZCj+m8Bt4CB3d1tEyyrQ6InQsaFqE0vBNfkAGSLbyD3MjJUNPioPdA391oyF
ryZ8N+O3RkH8E8UypMFAEgGV5jJiCmsiHdPhdv4ZIQnld+SDjXYoh8DSfUNbRqKe
BIrsJPSlqrEWvmVu6AA2hJ5cHGMWbx4ndMpvnpMzWCmAwcBN0km9ntf+3QnrcgVw
Diq8TmaxToTGdDhKQViXjgJ2aPItSUHFINItoMOK8xlfZu07vJbQRnTo5IXPKqGZ
dqoCMG4ms01iAEyXaNJ2cgKmw0zm3pFzzYKLH54YdeCZZAkSU1LcI94prBfXpTVe
9bdloyu8dxZcEhvNEa7PkLqbTJU1E3wMJIZDiTJXHBj3R+42o06PCDpjiEu4y8k6
wq1rr68XBBK8YIs6HGNe1m9OMRy87mAcerkOmsevkMHxNoPKWo6WsP/7uE/EjmIO
SF3YHkhXPQHB7WijTIfJZ6WYwTTJdnf/o2iS3jeIDILhrO15WoVsjMXVGRDewRXI
HVCk3NHY34j+WiT92cL6aNZEPz/1CaS3FIc6HXpH7dQkJ4NyzLgZQ0lAaZiwW1CW
FwjN7dZE+N9OXZJnuscTfEcjaOv7h8vkjklqSkHBozkg00bZsRRvUpg9KsTB5Nif
E0Iis+nG6b49t3F1GzQpxwNie4y2jHUpyA4QZUVrGbuyHWB5BW7nywVOjc8DC2Ax
Tc4SH0VOddF0Z4OhMT6AdMIh4NlwEwT3ixkaTkn/wmfP5IhoX7PqIsgfctsWeSKK
uB4v5Prv1AKyw6meiXek+cRzxDnVjgaTrezp/buAABogkLA+teu+plammGHw1fxe
lpHxvqj8Ah+guwDeK2lmveulJvE45yOxnHDY70KB5QNPQorxQrlR/3ggQGE90hNo
Q4BpmZDMDkzRa97bfFubQOq+28rakF+lBPOQue0X1skEuS1kW5KTP/kcrY4blek3
DohMZA10eCn74ZY+xk/N/LiCutt6N0CwUGFztFxhME8Voyon7XP/8QbwIgnkMbmk
v/n8OcLRlG6ND1cBNOXf5DAMX5j37UFvbhAVvXHE1XfDrr0iKGi+IcCZB35yPNu1
RwH7VH58MokGLZq/ltn30xmgiuW4B181/SsHQARU10tL/hN6LbCXApmPjFHktAaM
9tBArEKcqFqlKbe48k/AZchSOFtQsEpPge7hKDsuR9nGf19FDAYEr9oRdnxbtIAE
uRwhjJg2r+hlqE53TSzpG+xVCSO8VIuMdHzRNKh/Uls+cRp1Cz3WEVPtwN5KLIek
QVxrhHESCjTO+sUiLTkSGQLwGm0GhESYtsaCY1xZz5VHqWwLznlSNXm3xIglUenF
qiMmKEpqeZWlOnmyGXwCVrNZx+6/Kl5pn2XUfDnOX0OD3As4ggS2uU184Pryo2M+
gBLhgfhr6GWIov6MOb287sdw/HrMIWpIXPT5Q2mU85FELtJM7rKFUnqaAaObFhkW
ztkTO5UXRT7Q4vWkKEf55ygOWW42asfbo4kxYajjQVJSnt58jNdv8Qte9JL07rN5
qj113TVE5X+8oJZJjLMrZ2/r0+6AvkL8Gh9zsj55jLS+pTMZsJfZH1nr5OFFrRen
BmOBWtaSbiS/whKBg52KTmyL5McFcypmLkZ17ECY7n0573b0nh6B2cJ/c+rOif96
H0Em1lW5q9S7QrHgf3iEMsmpODs4cG2m4lpCoUXwNzP8D3A/R6miuZ+qiOOu2s8A
/J9PxtqaziwUKkwkSOGWfNdSV9qPJDdcANk72/emXolNMbbLrQknWiBu9jVAlB3R
ysMqisXdBl2/Y6GA2soAG29C2U2jwy7omQ/JcDlSjdYykcGdYH5RdRmJR8Vy9qg/
oHyNvWnlTnXo8ottF2KF7OkYuUN6KDxlA03iwbRNsOjWLvsPDOZPxU/OVfE0IRcl
lUf/tlFG93MbWt7CFKxt4vWOyWErHoXHV9jEGVZBPLRFSRJ7hpSpE9Pkv3XgnyH8
KvYDh78lRITpNtAewdYMdMVhlQMIx8ySy02S7+DZvOnp9UBk8Cp3m6JUrXiJ7wOz
K7HmWQHUhfD1eqyyUQJxmOwkgnKySsiAh5IIEoCcapj3nejtHlsI45bYOQmlt1j/
kvSqKOwOGKDsMBs2UHco/jYti6LprjLt+qpadTBuMXCFHxZ1z4Xb7/sHB845LFmd
/i1ffAQ4Hsh/PsBDoWg4j7gdv/wH1xFBeQ9ynQJsyG2nT4dXGzTY34aYBVdDW03g
DkZGmWTDcxxxFnU4sOD+ZKBtK/5/f6k/Te2e11bYkhTVGtj3/CHkqW9QZRSRg4RH
mTrod1Em0zHHsOMjF9Hjl9HTE0pnBZA5lH9XSTbQMOIo7Q/b5Nq+oSNrnrp1ZCs3
dkaEbxy70gdEkZgDD/GXEYVsLBC7X5nvg3XwJSGoE2DF2/XrtzG1sEmQChVVz2wF
DFDUhP2RwnTUuupmVW4Pdl6AGMN1iW2vIaUvHbVOjdZEecibyYnocrAKH8M/wZDd
dD5UZGTZsZlVAmL10ufMe5QK+k51H/lQ4b4WT9G2JZkElYesUm34qNV316dMVNkK
CiaDsbyXuNSOPAoD01d96w2C/Y7KuGD4d0CAelq2SMIzf2RBrdk+lgTOb56ejj/R
nvNXjNgtbXdhlNObBuBxkoAjrpEPyk9B+ZxOmLVY25Ojq56xytvIrZVd51fF7WuV
49xHMMiNzm+jXTElltl1aVH0qAp5d63qGNTqjJeIuxOk8fSr4qjgOnPF8kEV0cs5
hWKe70kDPhB53FtrYek19CQo/8iBxUkO37Ozr6u40L8br7grTXNrKq9ICPuDtSY9
r8zj2AB/HCFmfNcRC+rzx89WAA9kDECIZCgzGmYPoma2u9X+5Ne9jn/8mGj6sWy4
u3uwDMFnk3lAx/TJqromn066e/i7TWg3pMmlu7d4JYAcGcKlZNHrJ/837338rv9e
voLidlOAZ56r/IJehG8/JUvlRcxaLwRyv+qHpOkOtzNoq0RR+XDZiaWsQgx5e0F6
muDv2AcBkH7O5D2D6iCb3WhDlBoIgoSx6RbWCAkqo48usvfvRvMH825wuVFM7iJc
Lh3tpkUvRYMC5tWS7HhguHZ4ebk3CWuw6DCBiI6z8o29TitPTeMgczR2STcMswiN
2IKUIJIQ/lU+nqkt/MWqfLe7mXocZVEEYWTWEZrD3lETaXn4m+UJM0ZxpNsI4Mer
agm4nuaB+vFBPVs4t11q0SqrCsf6XNxJOwWpCXH1Kg9MhCH0J2Ar8ed8jv8/KJrN
e3UGQUKBZYV2yzTqvPz3WBeGWa0pP0bKYfXNA8dD2YqThdkaXwFdWUrHOIJiK5Oz
4bTqrqH/UNA2J52cGRgOgAg8CIKafap++v3w5TG1DYYsF2eb9M9RQqubWkcsPI1O
mbReS4KLGJhkeklDKAcHty/mQoXwc0pv35/a0PSEPcAOHOhTqt/8MBnW/NslMwqA
gpdF3LKvofWfO95Y3hcdp1CiQGehYz8s9Xkry/DNp1qaRs9dMt4pZUcf7kl1Tofb
xLfzqjR3gHrOymMlCl8Z9kwAFLR7j47K4eYvNjwctL7Xm93Sn4NOxswA5Uij+yo2
FeM1qey7GtxP8HieGhDBsdHEyHvxtyODrqizZ0B8CjoxG6Gb0kd9hWGRbnW67kg3
H3KTO1b6ZkSWLQuKZvkyharNpByaJBjA/yX0RlB6Dww1/g/pOgTA3UDdE21LO7At
pBS9JcpgbQghtYYMxsOk72el65mM8UTHrd53cfBQkUG8WkWqrmpxbkvaJ/Uvu7MW
lLU7tftGmmE5mZZj9rcbprPv34t0yBHKwsH2/E8jAND47gkXa09X6z31bhH9abXL
1TwgKjIv+VmZn4ucQ+4gCHiS6U1c7Pr/jEa6XN0rfCkl1sAu4GdHWBdOXDFoAU/A
mYPvaJ3GqwIYkgJrKYAJCMyEMiep/82kfoo3h8nrFGueLSTVTtBE3h2MUPSwJqlU
QacI4yi4yEcSvLL0CJbBLWfBWnSBjCZr2iXsOlrpXuPPUIyWFlSApmx5z5/rlcCS
X8qO7UF9vpFOh196Tnh1RtWwEtoaoHadk9ST5NYVb+BXbraJUfb/qtHZYiEE9oPa
tL1bmS0vF7Tbgrt+H7Oy90yhRc3SdA13vZSWlckh9bEaRCDWVDM6s81k1p7wSIUk
PwoGjRmnv7EWNjP+A3Q90MTmUAVRX4qbT8AZDKsqTTqstrX7dHeU3qGh8UjxAFiN
mcFOb2gfRo5OsKMP1ndTyjunmHa/SjRw5TvmOsuPYdMLiwwQeQKkFZwW8vi2/SEC
swP/ULcYMWuDpBqNV1zwylPG5QY0JUL5co14YVqo+PdMZHGWtHfeuJButc2sCbRL
7aNizPT3tHEoeCmn5rWwipblBZKm9FK7qLZw6Nr+8W+IpqK/9DIoAup9kaRmnBY8
4BKQGmCHsV9FBSJvYOo+Dk6NNHtXsUUyjjkYS+ZlDrwvfYpiNiYho1g2IxDDTYA4
FQ+Q0eMooTvNgY6xKnnNKLQWSuB/mMdsLuv42JNupMgDZccX2Qb9SmBU1KHY9Hke
1nOSMtbMI+fQJZJOA/G8O/+3Er2Opm4+ffeOGgyFJKIgSOpzSBq6HKXonJS4m9lU
aYDhsBODZMnSuwmcYGylZXZVNObV6xpvYoEzzqvww6Hwkjz17RaRXbfNjdYZMqyl
ChuI/rczHeEDFisJHS/F8emCvsaBdLgHZSb6o+ap69T7Hqkr9Yi6dgRHa946jZyo
dv34YPLm3PXfFdZk26bQuGbbaSgW0m7WKQNl6UpVnOqaQMmHfNKnjXJbnzzS/tAC
BJ52nfhxJysenRWgccnW7jeSxcGqGosTC9ms/yeOSuqqUjvQTP2C6PrO6qsCe1ig
ZKnd5A9QD/vtEO+pFdsbBnXS33ycD7XcTa3sDDrDOchVTmt++GiKLwi9auHXURcN
SYnVffXZERclauCz8YIbG16637UQin7iMnqWGx2vZiahNrIb03c+svLDFN/QXW/N
NogDI2eLFizUUQyvUwNcXBVWLUPG6SMF6HqZLikD5JoDX4iwLhyL7BdKMtaKw+uI
83SUQ+dzXwJG55jgsdXst2RklHMu3C0mJilR33nf8hLVui8BTz9H1gG96BRn5aoR
crj5AL1/djlFWyxKTPYGffktyjPjky8ITnVpHz+5EEgkTVFy8pDiY8H+qhR9Sk6I
ZQuGIj13wLIDH/vLn2IAVXiVhnIGqtc/vjb8v9xXF8MFig5kpiS6egwXddReQHU6
YJBY79bwk4uQkN7v4jWFDd9sJiMBcyxttbtyzqEbzP8G0TcvEn0Sth5swzK/AED7
b7FKITZXARjBp1G+qVspKGVdXr4xCI9k/JndowtF1TEq1FlUgUaPY09qAOAy2Ux6
5jVuYsdFlOnqQfEs4xHI0OYTYhFwOu3FYAjKcQqQnRHqCV3uPZwwMHPYbzlwmyPg
o6QSHwvsh8h9zEXHNA+Z9L8EwYW6DrcsrXV/n8kV8kLN9SGx9Z9CI/kBW6JMxEe5
aUdGmCBlY4EYxZnlC6YzNEGdxo6bMaLNXpO9tdExC2b73VetROb9Y0vnBRmOKeHI
RrFDalnrEm6W9iq23r8mZycQUFqdiyt7qySv9Y2oOdyyv5pYvp0ogUZrMXCuHy+W
l9VYlxKRneIPX8FOAfP8p3fi5bTOA9qErF/zUBiVTSY97YfOV/AF2yUfZaUbdCYB
5NLEUzHhfceGh8caM4qy4nDWjv+4IewHeEewkePwy3r899TKQchFTwaYr2uoRbYx
bUU+Sx/3lgKJOYy6I/Y73iEJJQG9M+R1fzbkeb7Updi5VYIS4UlVYiuWQY8PrP/U
P4q5QcHpBvHwH7iAffGPknViv9gL3kKiAeRWuF7BH7+J+s/QDM8k1SUf6ZYUPv7m
aWu8iGvAhSTsQuGVsIsFd34U9dhOdH3Tqi5G2lYttwp7IpXDkU0eD+Nr8OqhZ6Kb
WKatH9oO6n/6drqHo5zy+6WqroVQvvvMrZA7z44UF8ftp4COwoYvc1ONgCXjN3Cz
hl/zPmRm81A9fA6adLRIGX0Kwzd7RxsTiCOZBdeuhvLtoa2ggSuXrpK8CKrhhxTU
jlGb71BkvvP0wtMlJqHXHCUV+plcaJW0hkaBjJxu5ZkJfhjQiJkeBWZ7iyeCHIl1
DDAmW8x3J750DWyOdKuYr5w3OwZNS5hGK2Ngchx34tvs80aQpcOpR+ElluLxtG6v
8OLSvyprc2gicYlSe44kf7QgDTzf5LQ3MK4Xo5wKBC4GwtiSBDB2jxw+j/xTaybj
Tu4Zy2OaujhBwWtit6z7txTeuMzoCA+b+hqNTiwxcl0mayOtNofr5R4NlUoefGli
m3VtUXJdzR+OyLZBc6OCN57YqbWoc6sBD7qnJ52O5mr8N7iQ+dk0XV9hRD2n2jgR
dZPdOZQWUoIEgi7mvoh4Tcsw3RaLuujs1/ZpTqH1q/uaXzZeQK7W5AF+6yvgYK1a
1riNuYHFnFNqZLJCFCpSM10pSmLle9wwDp9G4W0oCpJEygoooGY26TkLuQXQSpzz
BKKUFMe4obpEXdjUeAMoAA+7Rbnm4nShRpl0zHbiuiE9zGcxl8jnPkWynPXk0VUI
INYt8E4BpQlGfdn91Y7FifHm4hylezHmV50Z3k9/YUDLglWA6omwG47U+eZ5A7eJ
TMWgvw7/CGifw4GS5/shWwlKJ7JnxY9v+1Zhl1GXpFF+fOhIdz3yPQP1LwAj3L4e
tX28a0zNmCYuy6GTaF0b9sru0zj93XBYhNkFA67BgXdhlanCGgcIe1EsyaYKIPJD
6x/eafC4aKYvo/J8/LimCbg7xYyofGI+SUb3CUS10aiWQTxH98qHhKvnLInhpuPL
wE0ON/f0vt/Ja4GwPuzGl5zsZHM0F6L9KwPiJJQQEshfTEGfJFzYcepfxjPfP3T7
zcLq6i+QYSR7oT8wltD08mWLv2cqgk0ilgQRmgREe9Mff6bnQwCjDJOEWuHRh5K2
WEBFRzQl+a5RmuHV8k+v3HiGahhgQ40n2Qf3PxnrKFuF7viE8jGQdUH4p4mmoGA7
4LRtdJEKKZM1t6a4LwapAbFlSa/0VB7OsxADaYhgLuCmv/wleIOZLgE0GJFE9mdg
2nHw1U9xHwSfbBNcu3oT9mBsGOijKMb8pTVcaM+UPQq+XQw9AnuMLMf6bjPcz80w
+An8m6xFxJIHSuLi/eK1swLjrxot3Qg0hMpRII9scBA5VBRDKgr8UxHOvxr5CTH8
Lj9IwBn5/P9VAjccwp1dVzStWZeZQ4ETitKjkkhXOKaqBMcq/hAHbPB2iEZejG0Q
Y2qoZrOsXiGbTA093xXsvPHKBwmdrQlKEYKFbc1DXPtYbW6IHLd8+b9droaUOL67
hURG7BBHmilG3qbjugp/11BRV4tw6qd5AjzGkkNCEjnGNDSPxHiie5unsRmca9+F
E6PGuVIR/YVLk5mbVz3fkHzCPl+cEXSmn1rtBDzMjDSH9JCx4xY5zEzNblTkI7hL
vsPwoWEJoNNB/rfnPJe2EwfiisDJmQ2BApfMYV1OIWQhTA6CzLMZOuBBbGFK6FHJ
bnOiGszMDy00LoPh8mGA3x/gS5A+7scU+dHieLw43/c+jL3QlGmlkRgcmZnF23nq
Wt+WBfQ9sNfD7q/PSYKOemvOjSQITCGhDNVrVwBRxQpcBhicqspzsE94pYQNQ4u+
dj4ora7xYIfutMwFA1FDy7NpYvGEsEiU3U2kM+RSufP1eF+xoFdTP4+U01/Pv+jn
gCHG7hIwgb9Rxubqn9ACbqygkGEx+hyV10FDz+mfkqUHr5qlC38Sy0QEKo9NPLbk
HzWvp4ifuIwN/Q0PFF7ro+pxcO7+i9zejkinOUcW7XSSbv5e2CwBR1bC5NBj2ImW
lOu4DG6t/2aO2qZnyq1xp7oLKjR3dY6N6RmEySHCVBzDxCIBTPnXAdRpR6teCfOE
NxgH28TUybbuRGIvrtmn8va0SZpxdUXzmvFNCAGZpvcsKkSloOobrdWhgdrcUT9T
+DhyJiPFIF6fU/tliZUhkJv7qlIeQWkRo9W32VKD8WpKb6En1zSD1FgOJdARUmuX
/Z+U7c3la9Yd60IydU6NNnSFASoXaLImG5tF8fq2jleUedxaiQBHNIGddlmzg099
gORAbcGf5WzI/f48MjBiz4kvsV4SeWyE6+PI7wqNAAp7Guzs009bMIPY1u7GA2th
RB97LdRU43bjd27YF1KpBS9dzF4qdU70txBcmkA4L8sQ4WbZdCwlmEufrgIs5L87
pipqMxQq3IBxPXthl7rraFaYephnPe6Tv4gJPnSlg8wAsibX6/AKupV4/up7C09M
DJ0MJ+ASb0tFu/S4BGNJEorpYVYkEtrL6OPYTVXaOjRxRBE/sFrwuWG4VgX3ASxf
8vG0t9PCEc5g/HxC9x9r6YY2VR4AFyue7aH7QrqHedP4U3yoQ+RtWm2qimEOHMj2
KasOPIMRRlcirxSgSTZ28b16wFSz/5U1J6dPb4OYKb1Yeu2eGrEtFNogIQqXqZJw
a7q0Ka1H82zT7197H8aN/ZQzNV1SuVoGBuzErsuIdXcZhG1Wec8em4thXimatUwF
RG0mPKEZC4YAgP46JZyLgYiR8dT1ucvYQ17CaycUNqf99/+XZHQNt6aPT4ngBMk9
7ihhHntqkhlebZApejDSaraVIeNlb+j1293VW+JvsTN1elQYXjKbgjEGJ/PTvO2N
wdXILwZyJv9hUKdMnExv6mjMNeqG3tVE/RO8XK4Wg1mrZBi+BHV1wOwneV0MC9tW
7CIvtydTE4ogHPFswx7O4wmQ0EyzPrEBwwTlJ9GpfqLkY4n8FkmhVvb5ZRbIMr1G
GViBiXTCtobihQdQpq+KhMajSl5uRRqL5s5ZKNR2tP0ougAsen/NOZL4+QSSnVCR
3fmyO9AA563vjMP5CkE+zm8kVi4oxAnk5J1dcRgWVvOsUlvftQHegVYG5jHILoky
4t3/UeNNhj+WFsd1sxM5TZeIEoUzwlaoVSzBBJoaFLSq4XWXf4k7HyZn3ORJdFb7
QjOyBFySl6qju1zza6lQ530OPr6AIYSg2Yc8qZpUJefyqIv9yjpCmHVzgafjds/s
iNhj2euFx2ZPcDj718X5qBeEtL89Lw35OKzWrsx4dadcJR4RNVKeOXhKKJTOHQcj
nA78W/RNzIFf/v0S9YlaHS7Lw7scfSzQAKc0MsUzdXyhuO9TuN/Q1RJQuMUcQF+W
HEQ3enaI+7dUYM/F6Cp0K7NbyRUFVn+KZiRwFj4esq9NgFAcplq3ZA45FY8rx9+3
hLMfYs/OBWlHo8xmHKSui6YHQCLxd+9WEWP3FFQy2EnzDblKgucpejPBCz71FnxK
YzGOYAJqaNf4xuq/fFhY569lVXX0yeDTMWgnWDiFNZ27EdBW/oM+n2BtGEt3ykXp
+rK2rxTqZ55wl8cYZs5RfKewTXhebCmnwiEXfnxpEm4ea+VZTwz8vE1aVTfxHZH2
GyBGnVy21khrClBEXgGdjjUyKGhaDbyIR5ZNlqX1MRAT37aZcxRx+uPyHRPHKRVY
9m5Dpd/TjC0T/f7WJST8BHw7GsZ3x6L9G0H9+XsM2Sgk1RVjOMqVuXDZAC/FpbRL
MChGE9nJBrDU4NsFTL3htyqkZ1LmGG/0gpgY3L12GJlqMm3oFOZBUjLzzC0Z8s7w
5h78OzzQjAz77ski7PaHffkrwPfafwteD8a7EFHUG9nWWyViLNvEr+kJyxa+dFWW
uhp+B6e1Y6pTDDbq7A9ntxJvWfWGql6j9pygs1JLRnpKLzBt0jJSFGteICPP/ri7
aPaq5qwS6dZfzVMbbCVMmMyz+JpNSZNKgKpRpmAfEK7NQBsZu4l4LxKjoNS/TBFA
BD04HGUNqdCLKukpohDNKss2IcxGdJht8JoCcdniupEMEv9/S9VtwOFhjeCmMeev
VcJf+k7A5fU9FduoyLwhA69rg5CJrg3qo0vjdhfGb+SfwYvuNBKNyYRxkPCwvQaC
KtcXYqoOw2ZJxr0rcGSkaWPnEISwA2lGu5RMTnz5lSM7T2jeSMQi9xJ8RUEF2zsa
Gxdf7gWhKcCQ8QLGKYUeNErx2i7UXldTN8L9nGe0Q8BiG331fg1wa/J/cEpy6s/U
FlWjdYE4G7u1XjwH1+NwmJqOk1JFTCg/30yy3gPAdxffzoXBAymRsxLQ8MvVj50w
exXXWAyTtPie41ZzS9imRU279TdzC4xjOzHJ6228lgIdTN9kuWj0xFW657pU7tHp
Ra+SxJez3uzit1jGV0PRPjMTJKN2wTVGe91QQzxfymWt1UrEx+AefQA9kSoeJot7
ZWoEmRoJRjRFq3QGtJ4/KKj7K4GBiipIluCVEi3VCcFB0RwbCreHFbJ6W62v8MwG
x3sCCYQTM4b6bz53Sqk/oNwmwdCp8/cy2U6Ojp+E+CA6E0y9dFQPUQzAryHFa1pv
7hb+3BRmfSKUgrX8ks7x14AXE/ZQY+/Ox7GKSkJP36xuSAbwROlh1+7RAN6lLY+m
gYceBnuorfBzhs4i3FRRJJ4XtalGQX7gfkqKV6Sfye/iJW/HHaLgK1UdM05BUEdz
Z+fUhhLB7bqh+nkWr4pyHPzczbZcuaJqb/rrRBQJBDBjqMLdHf/EH1WQE1+QqKEp
7KkuYXtsr3T9k8WIKZxdgsN/Rb9asjlgE2OoKzH5kJOSLDImmrcQjDtzebBX+RR8
/8nbsTpm8Nb1GjjXXTQ14B1+3VoifjwzmTDthTsLQ5ap4x6i7CLhH829VWgO1nvd
tS0nsZ+mRpJvM4yz5zZFuI1i4omDVQsVV6e7srzoke/t1uV1YUjG+vyBMguLbNTN
cF0WXwgw6d/MS9OwngIA78QMyB7hthlez5vOshZdIi1nJYTudKjHmsZ70a7Gkhfp
bmybRcvLYFN+NCfooIJqjgK+RXIJkEEU2THaYtx2pYbOeUeGrsIE47vJrlygDYhE
LVPnT6/r/GvEmMsFbAn0iarav2yVNbu9QTJTi6dTbBhGrkSbpmacCKpQ+K8IXJ4B
mkRevf4PQwl7yLE9ZDTCCLnbIZAApe6VTOzTmgBnnsFr1cT9blwoGLQLnGCwKBg/
Pulpv+wpRvNRFIr8sT9iq2EEK8DuaY1c1LPKz/PQBtDn8VsapPf9B+ssm9UbYpik
41mA78+FK+QnSu+UVpT1kRTuMP5slFiXy6KOzHzyc7uXNmNEr7vTf8MkM0fxMER2
ejMpkQ5GqkcYoJi/BzKXoAsboO52l1zV9s8hWQwMDNRJvyXfRuiZsPJUUtNgv1ZZ
9xcjaWTKo5u7zl/vAnRrrZcToccqCKdgXGUveN7LZBGhpAGOfJSas9DeqipsNtLm
BH11Q+6/0gDXUJaYcQxDNtmnILOA4yEz0lTjiOwGSgJyHwwkAWrRMqMawf8lStov
ytDrh2uiMq2jq/Qxbe6KIfOtn2qvdCgqCEmi+RPk6mrXXv4NfooEccOZ8QJa3QY8
a4UdTg9JwjGLbDiBw7c/hbxp7TWe6yceLWKcxHGQJWH2WPo8tLizjpN2mFMiW4nT
0bYB8rJmcMkMtAVzonM+uU+uts7c6vBudd4ZhbtbnAluPh+L6hLURRuM/IY0DORP
xQzOM8OHTtOcv7BRX/ZH02/XY+nO4F5bbhygr0Sw7rYQTuWVmemJAuUlCAizFeCq
SC5AUMXu74GtNzbEHyYddG0sTGuoGjesZzR+O5ZjTDMpVso+l+MNFa9nc/p2uMqi
Qco5wlG4q/q+QNaWgRweVmmKHZpG/+7wPAajqv3YEgFv/fNbRk8dMf+GL7B4W7hg
maFNFnRgHgf1K+N2vmt8/sYV8VT5bhnNzQSvmkhAxHaXJqAIQb16QXeeENnSf81v
cdWtmqHegG+Wp/c6P4570yMv1nbg9voFlXnesMzcMFhI6C+9CwHOi07fr+ZJFqLa
pixud96iY/uYkgQH6aPJP5OSzY+awoqTRCSj1nRowEwSNWV+nKgzTmN6KpHlynnM
jQM3O9S9eTv3fRqNLgznh69R0n9eByyuMlCG/W3bWykiYjkq/hsZNCrWd92zrgdL
Hy8pKu12JeqUWxdfhogtnAZXeKfWBTUl5v9mmJsU/iVJrxAgsImy8daIjCmDfEkm
pMixsMRVy/teuVZDjlrWgwarGhorq6kLxBNKT2X2aY45GAV+v7JvjaMbB/tXUyby
YDUaYOv5VkUAUMHMp7XRcdmbjS5cli7JOjJz+GNi1odO601DIRjGRuyPHM1rcWtD
XWMBVFtENSm2R/X0YIIPhsNVwAkDeeybZLCM6Rr/KE8nCwCV+Zbp1+Qoj9iurj7w
5xBtLjFUCb4RL0xvXymeqK9nHtFkbNtOZbOrghn+BD9JUgOcZYki0B6iXY3wAxzV
SDb/kRbqPjbXVWtBGYSnA5HOvhXqR6EHscoRxnq2n9b0IuM8+p8t0k6S2wRgzHaz
r8F6izo1DI9lgnXmL4YvcdmkM5TakCrYChkVhKdB66YQlrzH09rRpXfdDPQpvTpJ
DprVjfGKV/1ptwNahh1Lbw5vPXDdhRh48ISSE9zr5BmJVBY7alVt91a9Q/GduDTc
OqE5KGZhON424RCK+gj+IZJhE71WBVr4f7ajyKLWtMZikNpHhR8nvjQ29Dml4YOz
TBqVb8SPIpuzCIe9W+UnByP95VMHL92ENjT9CVI8xmQ44XCfK1bB1h/XMy+MDNKr
3nC7i6LPdZE/Y1CFBns2EDyHyIb0dxfg4zppcrKN+l/ILwENfPnyt1hRrHRirLzc
SUlkiIRRzZpSN7YysTIZj9GbFwV7vtl1d7eDtiyVlarEZow7u87oIQNRDDSJf+Gg
HiiHFylyxl+LQKSytoxxZ9mv4bskw9tVvH4Ixj+hzABBQUGzyUfx5XP+VqHkDQY+
46p4PQml2Ya1bcKk+LkNCjYVEtQJjm4wOUb6m3p3XBgkLmFVDodhmZc/22eniNGk
up/WExc2CQ3GRJt6kwVHOLP9mI1bkE93H+i+SJLMWtF01CNXaOCwgB1VgmhrqrKN
8Z/M5EjnFalfxuSl3empFc2H7kh30v7g3K14n6CFjfT0Dn0r4WzX0Mq/koHQafMf
Kjpbau9fv0+GC5LBaGwJgTYkxuAE3s8hw6x5MYdxUuEjQRSovrgwZ0dowQAnkSAT
leetuTBHjQ1mhDB5NPAUfThgJhoDFKTvhNQU1B9AyNdmFJ1bA8FpJB4q/Q9sDfyV
WbkorxnXi8/BjO5puOThmpA57w1oNQq8a4QfmfJmajvU9PcuX2XGvWgatQQOeQdq
edF3PvLQYQWfw8ID43XtuNeyjS3s/S8FB4sZMxPJagcwsbBBgBvt5hLgHfOBPz98
ouVBf8xDLPhSfQeOGzPKYrDiLiFrA/BKUteU7RiRvn4JRp1HA9QMGkExRU1xDxFB
4vEWfwTYlKv917IFAYZGpaZd39TebZj/U+1hgL9owQURBdaS26NK/o/iRUvoc72H
rDmktIqQgdxZ0u/P6BEdAmJXALFh7sWogd0XztgJkTkynuWWjljrALYx5uzRZiDy
ODFfI74yB6YYmQjJh9b4hyCwIaSb4cDpx7WkyScw3k1K8++lAcPpSK+NJ2QKj5xp
LATYm+XABY8pHYOsPqrTh2SiE9VwgAnb9gG76/21Xt/3vu+UjWTepk4LEDn/MaLN
CM1LAHm64/3mEwdDjqkghE6ICloqlkYX8gwiV+MNVqJ3WnY0mGDgsPenUlmLmxD6
0L7lavh8foBDDUtGEHFV0ONJSog75uEriN5QGi/l2a63ku9+ahE7eD0E/lJwdbqd
vDJoREc7zO+6VSE9O7w7sTN9AdHcr1Ns0ghJq37LLOB2/G6SUO95rSGsGaayRl7z
ndIb5bTBZSH9bhypTvqpMzLO+lmF23w38eIZK1f7XkjrchZsVKuoHe//ZsvTCJLR
0Yjrrtu/CVByQuL0pFOzIGsmXzk7SPWFLLXv4g6UHeliCtFMAOqYhcHiXh/474Kz
ANyTf6sXnPu9O5iYrvOOADiw66akdo3C3yzi78yKKvM/VGkygtS6zolfiZCrz7fC
+Vkz4o7AOjN6J6ggYYSoSkfOSJfByAaJjlCT0XFup5zcF5CBPSqW54t8AxQlkMny
ECbYfJ3abybTA4Lqfn8gzUag+ZNbN0Udp2jrNwe1GqDMKQwuFmYw4ezjJMheVPyL
sTsS1J/0a/4BdSzRU02ztDcas4chCb0SJKAoaMkDbCvhdglTHp0UHtjmjEpf3zTI
L6DHUZ+BgHxQDDHFdUIKFxA709CJr7NxvBrXQ2Mz7YGZ+yOfPzXQ+wSikzmyGGKO
6MFEB7HvUPdDQBMuXDNm7IuVXQhryxnRK7t+Z/hGchL0RhvwfSCl4CqWUTAfUc6l
0WYukyQfPPi0cx0IgxqeBRIgAvXqa8I0q+HYH+IUrWRoZnQ1VQrxTqJy+w2d8GRF
4Ht8Rj8XTTUXOi2OlrS9RV/VPNxVWrHA3wLGNMsEhVXcsvXIzvx+453DzrSra7Od
MZBg+T8cuNAVBPJAHdZ2qANVtYP7wMP2zB6ap8Nw2UFygibUtQwD0Rz8YkvbUSlQ
dOZrBHoOiwHNw2vKzwYPnr+utYqipvwW/a1IY76jeRPkQl557C55O1uyJRExGvv2
QqHlPa0F6+oOCSH+SkRUyrteBsh74icQp1QuQ8Z91F0awsYOKdcvBSMX3LQW35ZZ
bD7qSQY4rS3YX9c6DjqWrZGty9caqpKnm70hzMaqSwgErZwk/e7i8WYEqe48x79f
W+rLVrIp8ZnQDWEjKLgFNBWTkH3ePM4/8WjUyUq4begUlUcxfvJGWtY265FUaasu
JjntYZu8QAoApOuRo8CuW1DWVTGcMlvi3Ai1v6QhzgAVgRrGBW/AtgKQmzkuY6ix
zlMZVUN+XWt6Q5akIQ7nj+Z3nvD568wB2+rJb4W7FDpracj8c3r1tK1wJ80/Elrz
FqXMHMi4+nBN3T/rcpXByLDb0TVzYOXFzJ6AoP/oa2HV3OWaOqov3Jt8ot28NtVb
quScrZKoYFNaFRTIHmbb5kZzfZ2Tdzz8boZgbYxQpg/J/6o4G6IQn3gBp9gsAgH/
DYKQjacLGWy+EnhNDhZAcpf75IxjAPnSbIbwQNiKsVK4jiKfS5he9hEAJPggmWB8
h92OBoHREMV/kml62/fg1bCEr6DxiNJ9kBWreqryVFPWbQBWhYy7+SjVbd+HL5M8
2j03GAPex94rC6zV0k5C/SCmcQWUk6sTxhNSa8jRc4zWwRyNULf2SyQKEkby1s1+
QQHYM6aQf9TS6TU6KukKl6xDxGOt3GaTuCdAQHJ3D0WHLU3hr1y713kvpCeHgQ2j
k1IpcNbtVSd7gVI4Ni/Dg5G0aPYcz9HUIltnXmmwl9ukIF9tOwIDacTy6nh2Ifad
BySYWhiXMstce9tdihw0XbOxrjzp4XrOZow9C232N5rQdocswL9UXPDAonF6t9ok
2EJro/aj8UhvdNmtMaHDLjUlFpMgX6+tN6zGmUoFqIfFmLx7AMEakqXfixu8Im9s
gheoisKRXdyGrlueBl/5NB+lVPU3BXI5RV91LMY+jF/A8iGVDiWbdQgq9VoJPMlL
kk/0NYIudclelOih5ZEzLDwKnr+sQvsrKrt4Ear33cbyKxmAB6BKhmHczxQo3+mR
KErvrnRRVfvjFnpYTMl7XdEWE52pHBbZrpq36D6miXKXpQN4gJDWBrEzFBAr5suV
jCYIl0lvF/66M/goyllvgAF62N5i3aOBFRmk/QQVMxBpFFjTEqt99UdH87RQofxi
iUM8S9XgsT9qmDoWgKHAOgBft7VSsNReKwDPh4usMk/MYiUSMLMtoeyNc4voMzsC
3C31wAc+Jo3RN8XPCNTBZS8k5Yedbgrzmlv4NFW9OW3d3X9gjb1o+b0h/LJ1dFaL
szczZNA0c3nipg3w72hnvoq4pVPtc4dlaALZp/vypegczIkhIHM0OVtjB2Sdlpst
EXmOvxIc6dr4xHFEAYChHBy816Tvy3bJUcPe1vQt/q1PyMr0EnlC+PZQs6pOoUrc
CnNFB5qxbj82OIOOep2AQrFflE8ey8ry0Cy90KwtdnFpMbGCMth7EyFnc8jP0RCU
W4yx/0qE48EtOLzbbnYbGohXrG/N9b8cIDp9vtw+IrHDcsLt5d7FCnLqcjoyi3rh
cUnbJFgAaJndGJARmxD4KmMCJkBZYlkhIMAtje9X59QjigqTF3cbTro/yUIC7Brh
Uni1jmOzcs/fAL/dWhBpxYaj+TBzvpxgjWkUclHzA52mJU9x5gXJxZiIVzyjNkxW
IP0oCgu/6iDub1+ZdgVeKJgAG8xRbmt2sA+aqn8avNlc4lawyIB3YP1zjPJP7ulj
5NLLLYkIR5MxgIP87qKupgUDDMN6iDZhOGuNzlwJIwUiEqeuvmPg9QJlOaez9LBj
bmkFjaEZya3qgximOVfQGoYCf34SalNxPCpUbfQ+WctJrKIU65OJH8yDKE6haqke
EGWKpCTdZ7WZUtQAgv+X+5g7T9ALCizOR2nAx4aKFojfF3cXxw1Ju1AVrA72TioZ
f2OzkTXuyBEp8tFL/Qh65RpPJle9bqWF4FbhFskcbr+UATVHZa9GW90NEEpwo9Di
nalvsBY9A5tcpqWH7RVlUwqUHn+R+2MBTJLqeMH1F8T9HCUCP5KovhSaOnaQT97S
DqJ11VLlU4dA+LQX+TAwkDGRmyqzWuFLVwcVRsm7IsitOPj2CmdHIsXW0CWPdVnv
ibibIttJiETGGscqUnHiy/flz09IiXVRg4ABxkVXqQogtInoSovzjUCdTgEsJYcP
pHoNZZjMxBM69fSMtFyaDNkZEWMBHy25f4BWpRfQl8nzX/eP6InP2mldrO/MjEQ3
E78z7WcpLelvBCpEXcKYN2YM5SVRhvWoC8UVbOa1Zx+692ggLeEfbwroigJW9pUY
En1c3ioCJ30UpyyVSmPsNp+e/md47TSwg7YDaGy+fu8rxZdOmtAP6p6NE8U7aFzF
09oaJnQDSxj3tPtu61sO/F3VK20UD9RnXgHtOMy/Lsxky5UeNWbxdS7qlDN5Nbdj
sENtWM20wWiVsquF8yfwrYNQyZFJ6JzM45W1Nva0Hw9kdlZ1ApD6UOo+x16x/3SM
qBcwvqJceIpavgqMIEirEQHwXvGlR3BCFmxqIQFEczCcpiT+EpdvxQqRZ9vZFYA1
ehB841jCVrCwg73JxOgty5fIbMvwE3GLwZ9yrYu6Zc5hZMgEJ8WknqLr7d4W3cZw
EAmS89oT5wMeVcpA9f55444qMjqVMxxUnaCpG8XlbQKprsSy65ZjDz8AxKl6XT5j
DFlWr0hWItwyFXVehbeFbTJ3H5L6G9loqbasjWqKH4h7Wrjy2S82h4SiiNQLhcNo
nuuLIDnqyZWrE5dGFJ0v1H0iZMSvUtDVT2h0ubOvk9DXxA9k/p6Ffd7rn7s9JY8o
z4C8ky/4vSx/JPWSkm7hGYiyphrTaVxf8WFIQhz46X+IVTgqRQEfMbQy63Xwajb2
s3DnKBA8BOUeigUXPsyRxq8IH1VLYWQSBDoOd/wfbNNRHn9Gb6C3C47SrtFClWwF
cVAJy8FwqfzjHywRd46LtCSGe06gnrqQwhU6ZGQudfVcTNyCWtmRD3osCtODYWf/
FTatOcgEDsjbkZAdK73nMPpq8BS3oA37ljWiKyS8pqeU8utDHIn5e1/N6oxyMWlx
8NWga1jkZfXc6QoC+NIgSq/dzh4AimtaptunX5pvYkZyaUpgKVpJ2D+S8Kx64LXh
0lVfTTIEUgCvLWZN/4oF3KUXUZtV540Fx5hQInVPnm+bcnpSP+TmM6c73H38lQkg
TsNzbvcngoS0pj/+bTpPDbOCW3trTHcN9R/uiTsOUV3E+SFGouRrJ8Q7Je+8g8gI
OB+U2b5Z9EMBu4FF0MK7ut9o0vUf8FBrWB8DFE6V1DSwkRYZj1oGGT2meakZW6nq
NdSnHT+0Q9wWQ9BNGBByNNzNLGj4R2UU65apxpn66+HG4Ian5iKiC3zG47Bxoafd
0NWV++8k9J0yJTj5IyJGGKU0VK2BvD/iDUtpn1BYx6gf73xU2yUlN2JbraVFGDpU
oQ8mfOFXZubnQ8faiaIvX6a90ICCpnwQYM7Yw+CKhLKR7whQs2IiiP/HjpzCXAhc
F7ZmPMXmcVQWyLq667Cz7/irMhSMi1fFNaPSv3KpMR/w1AnxdiTvT7cxBVrnm5Wv
nJNisLOe1Oyc/mVgzGvC60gVPgjBke6FW/YOcYwDs0uEPL4u2lcdcfztgMmOW5aA
hx8awql3yGnWKQJ24FhndKZg97md7ZUfYX8gwh05VXZ8wo1RSzDmXeXH4ua44u18
MTOrb/eKMAK7MWHUhfUb8Jj5MFgeg9NPgosghODYNyIDqIapd6Vf3K0Wv9EM6QPl
tbQqHuxHsOb2RMYGjl/5maeLCx2hX8e7/5gOc1nDQ6iZbvb3GwMrE1i5veEkKyUD
ZlngVzRPNFOYqnTcmnDP5Z2bWtGXre7WBmZzz3fIXmQV5cZwj4C7CwNgL2qzKHRk
bmP68ICpuv0wnhlNgnZ0qCTEMASl2zLFHJlo5fmslZf2A3KI0dc2yW7JBONGqjhc
8QX81flNs8g6rNZih0gHw7zU8MWmqGMFRSDBTKlCyt1y01B4REUUmnMXOixjumWH
MTjdl6h9DoOsVmDPj2pDyrSKeuIWjIBX5bdNtRduqxwwUqgPQDxR5Lq6ADMrcbaM
6tpZCLiseJzbuMHycPia+NbDi1DnzsJ6B8fOXgYVWdCDk+25xpmwo+aD3rJa4Xja
gtRLcNMdfGGVry74LK+ZuEcl3At4QtCs4r78ftOLnxV/eu72NsPhG1Oa59JjQiRO
gf9gnnCfPMANYYIpGw61V2TyTy+pA99MiGf/fs5Eg3cwrF2KgL6inTQwKq4XsUxK
HzOlsrj09keaKZydCBCSWY6cHtU97fbrqWnSpwrvTfdaBWvYeVpMC1skAI66zZSJ
iBHK671vr+0MzQGqTXrvbSuSUJx4Q1EK9Zo4xPCIHZPFx3H/eV+2mq/GOHWntf7T
Jhf2eycqELzkn5hZ9e/upjJV4WRHLof5mk0igKXaOp0Z9ulkou31hgOUwQtkBsMS
QzD0LfEEmUvEquanSBsSm5ya+OwaBQccum8LTSckFeDoODnbru2zJNLYcbYEWz4D
veHlsINvqlBpuEAVgG04LMSnoBjqWlc07ViwJMyrFX0VvO+J6xqBS9nWxFcZbPYb
mUU1zbSRtKb1ZNslCqpE/oTBmzQrKY5FAmrx4Hr9cY4t+mTRZwfUVgsNQCVp+olT
OBLXr7L+JUKu9RPEpaq5nnsSkVT6rRfOVehAlVhJR1YUJNJCkzHET+qxpwqiRmKa
YUDljjLifEYNVWJjIp2ma9MZspguBFPk5gE+hj5Pn4Fiyq6cb2E/F37TcTtkYZCz
9ycK1TBhz+8wXcz4bnnnHkrv/itX7oQnQe6e1g+053CdzDyOnjKA8edm9r0StEUv
8RSfBjwp2MCd8UoWjfF5F3FW11RAwXbJdleEHMR/cDyVN/N/uGkumExIekccMLLk
sfQJVuZVCIB7CRvYgIwcaAZBmbNitEVFQWA2I1Y7twlVXxoOYNrCkBRt/plVYOxQ
DVPmGBzK2OqoeH13oNB5Q/XbqSagsX/WGhTVdSLE8Kike1HAe0JNuD3x//XUYXbZ
QlheIQRTFt4iv3NDpDoQ0ggk99u2maz0nvcVV4IvgRtiY8YVRYeFRM4YSDbqqG+v
jLijC+nZBclqqEXO8YkP+msMglhZj2YvXopm3L14T1IxogoWxhh6zuG5tJepx0ka
zkwNTyU/yRkH8vHLncL9jF5x14sIvAvkNf5b7qenBaZbRF50iU25rxXr5og1kOJk
yuJh83Idm0t4ehyidU1pmfxwlLz57I4WP2Qq5YXglwAVbypPo6AJI45O31oFDbqb
aNN3F0/uW6jeSjnXdxSWP7L8g0SZCypUlszTS2USK2OKfyWB78N63dnjB0DZonUp
QCOFLewE05XzK537kFrBzg365xq+FWpzDVyBvVawwW0AvAR3GfFjTi30Iq4dPwfT
TDLdp7NWF6syh92dYYZRxzGUqCDOSG5GKyx98XV2h2T3FoZQYho6J8Ddy5w8d+ZR
PYMXfwy7bvV0qg24l8uAKuC1HsVdmiZhD+rMSYjSRvDh+bZv1I+Upd8OZUOCT94d
/x+cQC7eXVe0bYD9neQpaJziVVrxItvR7+kCgNBB6taDZAvfs+jJ1fFRVvu1pX5f
LMhTVTEV/jehcbvD/GUcti7pma8px7DRDtEDe4EZAcFpb+hEvHJPnlqpX7u/mLXf
XWMCcBGSQY50xrRyEQwzmxUr4hc18UVSm56eFWnTYUEbh/Y3KGPfULqilBnf7THk
MdFqoukW9BhOFvT18BijYrDuWa5jcQXvqMK6K0o+4Dj/sOsVciRfVkljHhIQhCDd
cNCQlX9OONW56ElAk+GNGBJgRI1lQ9DhkNbv50L+zcRtAKY/jHRca/doXCHQFTdj
VMx+4y79sykm0dhdZxUDgf6CZoDi5cGi1aohk43MowPnyR+tz6fQOVJerbZB5+Io
hRcYhldaf2dIcTJ3EdUS2k6kUh+UmgVgKOm82GjjIo1JQU5b/BpB2sR4mutW7rlj
037fRTJA44HAPfeGyaagKuqZh28BExZOYb/c3dlraMyNhvdrxXc/UpyC6HRVx14a
mkavtK+ZPGPxMPsO2scwRLuIesFjheFncFynU7Q9ezA/P4C8RB766f29qeJsBBMw
7exHlYhITQTQ5Z3atWP8a6wtjQg1d+MTtDGJ7wDytSuludnix46wZ9Jafc4dAnFQ
mX5BYiqtaRTprjNXfqNFBDtC39iqwy7K0z/KGxTFw5WyIYxkCK+ZL5v0adJVTsRy
5yYc0Mg+Jo8pFdA+teZn5yJcab/uCEGmrPXfuPJ5AHhDlEmHeUSV/046A3Yy9gsw
Ny98gcIy5ZNHfZlJnYoCyHw7zyEij4BjGr4PA9VjSddPABiADuinGvy4+LieeZov
WG8xNGpP5nj+Z55DlrGpu18AfwGzgP4jYRpL3hgns79GHwHCin/tbQHcuP9IlVj7
Rxj3TcUBn0ng3LwNjYKOHSwMt+Jp3Yq6lneyw35OiAEaKezftF/9ADZf105mBuuH
k6Z2My53phEMv+Dd7MEA/qJ9dCCeXIuGAdd7K7fj6c8qSU7Xpx1bKoG1Juk9rjCt
3haKBwPCuSmI4hGTNgzhhl1ZxTxfJqnPWFvNQTvWNKpgu3Dtfti196TiyqT46eKe
0AZeEgxbqS9JWWq0etxIGyJjtMlYTlPcOthrRMe/Mu/geM//kiYmIctDyApDy+DG
L1+vlk8GMgJkPw9DT9eA0C2LpLZaH/EmDKsEuWnMRYpC0vVBo9wDyDNm3KR3rIKF
vmaNV78EvmpXcbbN++Pds2anGcJZNm1UA5DgjFuZfQi8jhkJ2Ax5tcyPie7ARm4v
LCgXwPmx4qMFq/Bnb6+3tW9oZ1Fb+JmHi+w/8vaitJY7LWh0Bb0vte7FkEUNLE40
4i/JynAwHcyGxDobgbXZd7UnE73Lzn/flko62tk3w93Wm3IduSfsDmEPSK3nf7rS
Wh/U88tsGU0pp+VdH8gWkq8b4cWFeAsdKVNYrk04Gy1p0mYe6SwTNWZc7PFu8EN3
+7ddh1eINMXSoYp655WrhsNRxy7wLgpxptgehbYsXFdQ8cd3QT+fn2taER1tBovT
18wPCKu/PjyQRf+2yiTKC1jiootvGqn0h4PW5Hu3VC2Qled5aYhRhmVCJX4ZfQTK
tGVQtDPYJakEmwSWH3oTYs1HFkT3b0qEPD8mHV92Oeu3MMirXRLKtBqwvVDZqERX
xdchQHYgaJfWYsM8dsLgsuKMjrxt1uzvJjM+kDNACOnR4u5qudxrDU18gSXBTra+
dY0oS4e5wnhsBs3V7Pe49AuQ5ptnFgF91c8GEisoGdw0/D1LZ9L3/ZVIcdb2Q10r
MWsJ59+5xsvTmMWeBFVVdoeQH5udxpZ5ui5dNs2zmdIEGP6UJhLZymVIWD6peHfy
7Hu0RqCytbTHI7upmxsEvqbu/tvv2MpPiU3F0NbjAYW2pVF6ZkscTd/CxJiPmT+0
yOIuV1PmrvIfh6LK1gVQWJlTjxBAzAAazTmWvAESGnX79Ml0zUXRdO5q3WhXRv9R
MXXbLeU9OIzzoPpyOAeNkrJ5O1Pxerv/Bk//e+PpTjs/4aUHJwiEHjjISEOZGJQx
CvN/SdVrALAdzQzYNAvtoiZ0t3kM3LKBgsLKs/XAFIQ7gtWqyPCv5WsN8y0veeAr
AaqeKoauimrwRwJWSVnythX3q2aVr6X1ZyZZZT3LVLND8RlCvw1TkyvoPqzls/WB
ud03XxC0wSfkyz7zQf4dyo6OUCojfoOsz2lt9SHsFn/lhjRM1U6VuYI+kec/0Yc5
uE/aNOm1X6/chyEYsJvdE84AjIXWpQ9i9HGVKhkMpXfi6EDjYOxec+qoZSphYqyn
+8aZhzg8XMHDr5VcNMnBX6aMvf9yy3MMS9+AkoVL7VR3lAULTvraDG9/criZLm4w
rH54EEqCZF8V5csxbkem7qG2TCS6dDjfEHfQFZpQRCCwFYM2iEAkQRa8Q2EUHJR0
024EJhkrFuvJ4rOOU+SB6hbdIMzvRDImdayndCoPSgUjlbAnIus1sQeB83u9opjR
/CqujggpKORhqG0RDN+TkR94SP8rI+jGwQbo3skasbPuub8TubTDaXIjSheWGfdm
s4/c9NkW3LSSLjK4t8TzoVtxKSbN7OojGqyqKHnYL1I/rXDAMRZYw4yZevD4aIeP
JQ2whHSdKokrK3yQDGQfUuBt2nO8NfOwAmXcB8yVtdq3ZCmX2W68+S53wGg0f0LZ
4PwIA3yBV0D7azus8LyZxByWoHtAT8IgQKxz5r8DsH3y2r6MhP6tnwGv9IAx9xMu
a8+rEoDK6fv69r7jWJ1/AS4ePMjtnoLaIsgwJ1nz0ckUKfMnurIvFLlvOStwDZML
3rGQqB+JBqPjldGoFKHF6js9Ii2lP89wQ9179HB4KJErp0o/MG/u2xqZlGT+ZCVZ
0DL2/VS5edCTbfB5Iv51qBq/AS/ubAV1zuOZIjNmYQHwBx3eWypwj4aRkh25FYRD
PKzpNhnFI+WRAryZg18TGWq38gFwYhlg8AeTcmBm3EI/T5+gCWLfMi0HxwtwpSGs
IF2qRqydw+7VT9St41T4yKCj0xxew+MfKIr6UiQG+qE2o7MjiXfe7MirTFKl+rDa
5C8+A2vGGT8amMobqB6znRrPzcUTAF+dvJLGfD4XqJvRESfd3CMk0xii6PUNAZKA
QQCKPxtUMyx8R/y7QRbCjYRyX8/k8UywG7lM+28rCjwMoZwMuv78g+w9mw9b1R0j
AkJNnTVlxHgS7Yvl04VvzEUDplwUAFcAf0hzfvRv5Mjow+JjKRW5A++nvM+Xrzgb
uRIaY7XiMenP5d0eeriEkji+Va7xUTSOBxDyoaOiZnde1m/9oLtepnlYGMmYSxyc
lAaiDX3aZbpk3rFwuGvYf399iy0DPYYeT9RSaZrS56PZI2AZeYPmGy1ZDyvlEjcI
8r9v+z+01CGOr+WckMgKaju7JpbSeilJTald13psCjkAiosxvOTbiGLFiNn2FZoa
/2Rh//5erRqyWvZgWi4UANx7NU6hgVN5OztwLVC3C97Fv+quZi430ZQVL3lYam1R
8isWIo94uneWN066MYo9NGYh8gZ+LzTKTxVmcsVLD3kNnxmuTifzs9OTCTMW91+M
YF8d4QzCkJMZVvMxnExXzj2zyLDLDpfIzwyA+6nCSdD4UwKPzXdDPVtKCbE5MT94
5PhJeWCcMP12SNjvg3eWcpr/5XkRY+WhWxPFaYIsBhse02Ez5nhIKNX90q3tohZn
tOj31W1NZFY8FqjPoTJ8as/LBQJ2c9a6gpx+wtxb9EY8J5H17o2ahfyS7NphCoAW
Lzteo1hXNKMcCZV+LcL7UXTbSg/qRHURp2tYR7rAG+PLb6Of3QA8QHh61MiTHtYZ
KSmd/VqBsg1/Hg9xAlVYjsEpc1N3NcKroykyenKknief3UJeKYS+IqN8GtR3PeJ7
DJPDnMUhJ54sm0bYPoxovmzvkrurbb72aOLmjpANpt1c25CV4rsLs0kHDjMwMoD9
HU7Za7L7LqG5CnT7rIDYNmSM2X1tq3iZjnu+8WRZP9GApTxlvCHEUJqIWT+sRBU/
8fA+38lR6YTgbDVPihLpXwsdrwHkxGS6ThmYuFbd2ONzv51kIEApvdjBlNVfpPFV
QRr+YEyEWi/GEyAvd4KSkvBfMeRzGzwrMS9G4Nz6jRHao7xxYYRRNCTXZDwcKKhD
00gh4KF5OVmnnJ6Af5l7okizzSNyALVaUw5g5DVeQSCe0DpIAuSr4EjRcRYK3un1
gInkKMOZoGsj9qgZvpR+BBveG5jk1CpwavEtxCb6l4BX1H2gxcnW5jlkqq80554m
QDE0b5UTo0ObOuDCShLi0V3AXRWz1gSkgAJHGvuPIAeDGivuDXZzrJ3z7uIEljlJ
DdgkR7g4qU9PdtR/qFYo1tQuFNsJzpuWLUHh4cehZygYV1WzQ8DeXLQ2e90JUgdn
y79ZK9im4s3jErDZpFaX6lfKDG0idkdeA4E0eyftgKyOPcF/cwR3aGa2FjzYgoIT
lMYu/eCzVhnwba4s/kp9f1ET6IJ2lbTAGKjhhNAVkfaUxLF2h7WlxR4BHkZrPelU
gv1twKyBWomuuQFzkxMI0QOoalz2QVcaR8C6tjyFY2dENJO0+1aVfSJtbCuLeeBk
53aKpn2qOkvT8Ysxi2bVLwtRXn70QVi+6N39wKLd+aw2bew4lGIYNzxSOgrNmhQ6
f0SGn+7x0vZ5j1cOhxTW4FjHRoZ1XNCugZ0u+Z/URoTmiMiMfhjVL4PyV4JXnI1M
FVzQgdOpquihBnO3If2VhD7Kp19G/m5kkt+CLSd6DyBtawHAKRCCaWx+1YHU2Bcz
hpPJpbbl4ieV3lrPky5EqEjWSq5r8A4TMseeKlgC4kP3du+0azCSmyK1Jh3KlfYh
D5evHumOsnr0D/r6h3Gu9pHcdBKZTJk3oWOf8wkFthqK9O0vbFtyU2qXiFb0qIC0
pIY7A+AEHyYJGp3RchOauyNcJ8IQG5NHSECdM0ZY65j0MNFm5R98xypsXEokOrrh
0l6Aijo0gZL0PmTOpp85xObThtN6N482//GP1ixXOiXXIeAat+oeOxIeLg5p90wP
REfBXSa5cMVtHCg2qosEHtzMVGjcmQ3rqCsFwDtNJb1Xup2TO5zLqxEYuN7aKJq5
7lnZGsng3iaQeGah80HCKI05YeEpYio0yC45DJcd4NTqVktvu6pHLi1dZTifKr2c
1FValzlr25J2ULQRVSrtKZwMGsvLBnEgQpYb1rci/yywJadzeMYErR8nANO1D5it
cqeL5R7jNG1opfTi2nz0Gl7PAB8n5oRK6LUPmTsv8pjci1iZz+QqtVrWUjazup5Y
AWSgZc7Wi42D2UtIIxMAdPNPOmnYVIrZ/FTHSBdG38odtLrIIDGv3LSSf5s0QGgS
grHsbMqlAzXZ8BSQM6iwZ7+XuVEIoh3hpYhrg1JHva1P1oIqYs1VRiwgnvcSESH/
miB+gDW9XecQPO+REmCZLwpe2apwtudQXaGD9ESrbIeY4ySBokGmk/HQu0xjgOX4
iMrqq5WXoGaNwMD+j82Q6EmqEBCuN2G2lJLM0cfZsA1+vC4QyqJnFVGa1NF0eikw
s01LY9DW7kWsVgv0CLaPVEcuAFUD7hXBojkGtW2NUmLsY2WsM7a6KNz5VGj2oLOV
PK2+CmZRetZFQqETN7gBirQTYgvdThxNpKHPvbDyA19yAGqY8W5XlS4sBVzQr5tT
jmbJMlThCKzFaoal6nhUij3rsetwD1gRkRiThJ8JzZso5a1S66VIwvrGc9UgOAAW
nLTy1x/E9iUYFahIRJmi25+mc7IcQyNqrWdIXaWSp6DMrjrx0WuCzLkYuNQZSz3P
AIY1keTQeRdr3CgDZasyUS7a8k/uwo1Mn0SG5djr+/URTY1l2F0/2dnVchW0Lq70
PnsiaZKu2Pw0WSSdrfKtrQ+1H0fmmnkmt7Oz3WHrEUwYT1I1ORNfTHos6Gvvfrv/
s0qYIOBMdjaYtKFtTJGSeJ9evtmuvdauWJFx4IUmt/M7cDOwl46roZgsJawmgv6b
lju1WvuixQBSH1osXJsEzE8cYabALvY+Dyq4W7EwBiqO56WipWO7m6Kof8j35Q3H
piH1zoTHuOlxcfT4wSD4B+hjadIbToi0cK5tOKWo46+tW0TCr8hzE7bh93GDTQeM
7Iykseac7nF5oW2kCFqU63bXHeKDy98Trytz0Ll0uLHId38V1BuY0G4ficlZgn1a
Lm5jPBSLADRaDeA5j/YgAsd7fFjwP2uKojj5RuRhMe1z/8yYM3fdAzgVQbHQD4qW
oEmvKbsfUIHSIMPbBRw2Sc3yY2MLidVFdbQ5PNbc0jOJD9WNYP9nSAYmFixStuMd
BKeyD7a4wGnA1gnEq80iEnmZWpDOZdcJBj1fPrmRwUPqe3QO4PWpfpRxwsNMQjlA
Pm6GIdQYfhdXPo/AUQ4H0xaI/+EhW+QJdv3nkjSZYtPdALwjQEFSjU5qTcYVUlY3
7f6yU2WyZuFlzgdq198UL2tTdb14vMtxGeCiqZXcRrxC5HTyFZQuuJIoIipofTws
Vorh3h/lPomRnuP/37IIwyJRvc89u5dECF8Z5+yDd2hl7K6cIt7jnOXe6WjlVW+O
ZVZwvgqqpyVscJO7aADLlLnphzhZ2i3E2MPAGWVHm3cOLety/6D08ERtWqqCOQyE
xysMwdMDhrhahDvAYXScPc3fVzA62ZJ6M8HkZY/skEVSYrofIoB31aLQt1rj+L29
ob9yvAMmW0B4rVtScuA8WVe9JREvNfa23S5R6JYyaXZ8ejFaV7rpdYqqSGoa49db
Ie7YWjZzIAv51zQCYUVyFSfRVkrHS1LscVDxiiAAiI/o/xlGchRL5I/zI8M4yFiJ
FqoIpUszO7XUcAM5XNA91R90SI/RYd2PNSD6Cn7tFDyA3G7OfQknGFOxfONzjbdW
AOr4YDvqLxxUlmh4sYovYEwoqG9x6h1MwcPTMg6sozaW1IefNODTXpQFoTG5xYhS
lydTEgV8FzXPZjl+U7VPqHOezvVX4FDtBKeNIQIu7PxbfG2zMm9DiT79BqGNI0aA
YpmQ2zjvSi/hCPVCylMQZdiiCN7s5yOW1ngZmezf9jtXFrEoEAt4fcnQeEPK1YAs
QBlASNVBYlUOVS2zHEQrzjBLAOPjFcFuL1W8fV15S7bH0unnDQcMHMYkoTK7YWqv
KxZz3ZgIYUQO9syxGpKxM+KpVaScFAq5Slsq+VtjbR1xG175KbRFkeGOmOPKOaCX
bHYoCsqljwNzk+Af7xS/YRi96zmyKhGrJlAJhu0WWkwjLcbW0hySDm/RWEPP4udX
ih2nf9DFX73HeEE73+m5G9du6f5TM/ZFYkq5VqqrHuGlMuFLglZbUk/s84rOKPsn
WUwRw9Jo/ZfgVzlajHdIfR78uHuCwFqC63+xM4bV5G3cv+K3/IvazS3KkvWysAt5
VLnrguo0ybvmhLuxpaQK6a09hTSaVf03VIJRvWERMrSg+yB3rryES6hXz8poa+V0
qbWGTewhPlgznpt1aywSI/xlBY0/i3gJOTr9UBHwDORy7T1mGBW1wGCotUyvLntn
TOmVIi6228fZ60dfCT2qdasfIv2GZVwoXaachzw2mU3xM5ftvnQJjXBbiW8iyym6
Zap6KgbKreBVpWmwrL92J6d/suXztpvLZaOqOjVvdbss3FmRHmG7BtFfN6Cp7f+A
4bvfKr9iM4T60AeuYbyS42FQq7rUDTmFLg1VogAAfIrnYdvA05RYaYqZnDr+AX0g
5s9gnPMK1GKn1zW5mL2V07DIvcYrpInMGLdVuidZ495W6ttqvXlMGLHtganltMut
JOt9QuQxgDZ8A6WHzNfa6R4TG4CamL4zzaoBy6ensXuLEFPwiUaeIU+YvCuvTFDc
7aoxlnnvwh3OK8wcl8gQ5zwE8v7/JuzzYd1QVfiN/f+TY1vVeZMohWNNwCOxnhaa
7AV1bzGaCDlpY3pkSzqRYFQsytb+s7cSAak5DiwKMHqtK9Lmyj8HlKiJhsBne+bE
z6IpuXQa/fH+SCsO+vhgQgwE1JcRxwrTwFBnEEq7Z+VwLQ6h5EASLj74LfveZlmJ
fEqCmTbWCsVOtG3Xx/IESU+hpq2soA6+i2UUS4LOaF4ly3EKHTK5gVWD/YqXcNEO
HHalzcdSNGA6ZsEdCUHjazlc6/PaafccInQn60+NQvdj8O13YUYrdQYDUWqVr+WQ
ukDA7+xNWZghbmm6xRf3npj68Wkez2rFwo/sq+cW+4t6RIXRi0vw5KwlrLNRpsLU
UDvBf/a34KdGnP9ZrNsUB5KRBdHqerjUdBEhguzK1Ad4bES905jd3X9fnxPs8o1Q
xPQIx9x3chjo0bH3qXTyhNiJLMHrVAf10eKFbJ6AhNuV9lF+LsaEKKF9KDaZa6/a
iJ8wewMbcsRzznQxIFV0zEPm82LZFAD1rd6XQx5ZY0L7s8m0M6CKnwwMwzAwAA9T
GIeuAU9MmtBbeJVxQyAIvgcErWHJK2UB/O7Frsb/4sTwcFP8Khccz33yicDcztNu
rLo7jxyzZtkVHXU/tEo1OX2Q14tEdyykwYUkiPooEsW5TxS/Di50HKVa+Eol5TFn
Si42pT+RDRvXO3enqjEcUc+cdIqiadWoojshD+Nfd4u2CtNCkHN6jxq2rkIKnSta
YrSG1943pX1+0LB1Wwa1DXMR+5tGGetav5gxw5dTXABLQzdfCHBna1bTbgdU1z9G
B/n07RIM0dosvdYeDOJJiF2jsCI/GNoPhF+o7xNqCJRlTXw5lmC8xDHH2xNnNMfq
Hc+oBRi++QKvjSh71jEd/f7KHSRH8f6R+E3hIPNVEO+sHkTwNIFjhGUIF2zBY5Mu
RgnSRcsrsSVQOycDN+POGn9P2CCtARpGjAhpxLHBsXSDXuV8dbdeYM4auOsFS0jM
f0xDEyh7PeCm+v1tJCr85k+xXVh4hNxLA9USoJQuXVKapi2cb09XRzieuqIkHgK+
6RwNxbyB8pu+FCRP8LV8GFKdOIe5B4/CJV6bBEoYIJcdKWK8QTdFjp9j8ii+QCRK
/fScyzCiMhKQFVH7pniCJorgiMJmnGkiBhzeONhaRjZzNctFWuGdBYR80zHzk1cl
/olrw5iutBID+yyO6mowVqr61/rJYJnrZ/shTrL4EVVDfRj6LWgurpa4LXSUBXP9
6OaD7ZpcInGmQE6GcyumIvAxkf2HfIEYuFJG1Tkyg0joZQSrES0htiddunBLNk2a
F/5u8/oeKfajGYSuAwmMiVWr7nDHYMnDD6vodOSii6x55+INaHaRD4bFeeejs2N6
F9L5mP/BVfh2M6UHQjS4b+zR91xzyTqBRzvb0TBZRCFYjZutR5Y/rZyeEU0xo3Is
C1s69GIrlBnRoMIFZDdeir1RevLGd0Tc8cgQiTE6McbzCRONKC46JBxVliSjn+QR
WUxGKDgSLnbC41zznDVHUuYlXnWYhpTliqICxxDWIfa3YyeddSz2t273gbuEsA1M
6UNqr6mNeV0P+r2dQdk8Z0gdz8z9MZjw1ojqTOP86QF/PwJlylVDgVCl/IxKtwhh
Skym7DYG6ItgJbNTUPi+ZcRvbU3kShm3FXC4neAs5XTjfaQm+q5QZNWO0knInNnD
yaQhZSpQ/pLyEtuK0HFm6VQ0F2cFL6c6s3o+QvIDTJF95uwDqUSy2TTcuV0nzap1
+5dBRkSNJsRTG+4BAvPnZhzYHz1gsngmEHEx7KvzpbfQgc/Cz1N7r1MsNHR0SCdD
WMe7TsJTOIiz7hyc2SwFu/bylcwXh/GLR5c8uGmIrOR9yfgnqB76CPaQpK6U724c
wsj6yp3Tan1VPzwqPtD3WLxS+OdeFpTitLV3THBzmwQhbXj2OGCF4FRK3As6HZm7
iJBT2rKUpn1jucFJaColyrd/9c9J2jjLdbfe3JgSmKoaZkTYFqKUowXJR8lIx49j
rNjdqPgFwvGyS5VgKQQqF0GarqmxpjSEmpW4tZfEYumQwtcE2GtsU/u+XksWr/rb
M8gsSDYa8aeDRNViS/qR4M62qQWB1MEYdP7qn9qJxfVZe3hT7Vj17q5apBUYJVlk
40v+gUuGsk/YXgLSaFodC7dwz+nTyFTjHIxMzmdA9WqmILFxmHXTgPwhkTb1DXoN
WBcY5Rr5HfRhZx09boL8Qp4BYvSyODE3VWgLMBO1Sq5U/b60b3An0zr/foRXN9l0
Jk5wTWwxfRZ8UbryoyaRvpImaJRiNJHT4WFIpBhOgFgnTeynb7u7FVvrkP+UXamJ
XJT5Gtzl68a2jsTIkgYDayVtnow1bsvZbxM8Ee2GtY0Q0JknaxXqG8O0QKx0Z2Ba
th/p5n5+ls2OPuyCwpwtutB1TNI9RPYITJYcwO1zHjKnVMu82yN9WzeO6P4UT+LM
k9+c8UKXp4pzdXub6S9b0eFN10S8DvirpS2IUc4BCeKE1kDztXXupcfTQ+yWhxDv
UMLYknhzwh/SnEYQsYsmQgcBAA9hFFVUYoawmQhAlDx/UyHUhkC83EVlt97xPpke
brH/R9NEmcRpfbl0QgBNdvJCYn0coN7vpjjq2wu5Ti5hh/ZiXQ2i1SvCfr1/rVEV
5H8mNZV0/PWc5LXA0yYIsHlaRpWku3nliYwkqA8p615cs0LrFxyuWOJNMBtTEMlR
fHunkY8nvFp5qZ4hyac/VaVHpb8K+/xBCcaOdrsIrmZXSP6aHkW8gQ+KnuGCcuWH
immbSZ/8Qxgugad4NNFmcifH9jOEXIg/fLs15z9Rf08YMxyA174D+2oPVKw8ZKw5
delbOG0oS2BFq9GMfyTkglsnAhWxSSEfqtETJHIs09lZVqNKf4zCohEBA+X8Ea1m
hf5rPi1oB+dPMM8iFtWqf50atrufmhciJUPP+3+gpHNeOFuXfEINqPF6xPDGW7J3
8+Cspu0+jiB7+eVpmGmgd3QHhJTkfYnu0SkEAd9qlkK0w8kpx4iuhsRszI6oY3fJ
mYnghawtCGT0kZymkEg8RgC0HOILDw3EkUPBbpA8rkYO8ehAmk6Lio0LG12vXDt8
t5pmOCj2sOHZBTsXtvK2eIgS/utAAPahclYZD3tT8eUuyQiCYffZNrN3wR+BYVgy
PCcPiXGAIGQCFFL6ZorcMqCasiWldZ2k9OQfUkMt1TtWtbvNVq3fOtgQ4SbE4Bqk
g7TH4gdfucQH3lBBKCYszI0z9hd2S7tnDCDuIuOKRZrhnXby2y7MmnCgE4kysxS+
w373mjKylTE7RTQfUqlEZHKLx5+sGRrbaCITcAHoOd/BqkLGuEXUV2QEvrkZnU1p
rPZM0HAFwP2EnwMIqYu8XScnzh6xhBjIbDDkmHzOXWcuweEQUTsKo2r4Y9At5m3J
kboHG7k5QkOonU34s2aV96AgQdwZcNv6iX23CdS1J+phYU6+hapanFI9JKWR9Hop
fvVq3Q6SPkdz89bcJHpjgvy0220pj/3pVChwhWsH0RWjvgwKhu8YbvOnX2NRmO+i
3JJJyxK/uKU85c4vcYvkiWrgsIsKcdI1exF/zzCg9zTC7kMkpdsNQZLwSPhIi3YG
AJyD1/onQ9QvqXTjk1IRaNZ3GrR94mQCbXkIkYaxiSS8803Q8/OD9p7tUXzW59gf
cX+lHEOfkjQBVvZsZYVEcxrdVpgRqBZv9wsZP0NEPrTEaIoasmFMmCx+1owb13Q6
7m+A6CoMcfYHjEDtNHNArogd3qC82l5pTXM19QGUp1vTQ45MY9CN8x7VcpBPJ9YZ
VdURPZNtRho67zR5eHJSJOpaGDxDxEROM3orSEoW+bXu1Xw8CMwmmVji7HuXgwhm
ekR2bh7N0255fH7ggQP4gfOlh2UtfR25kyycPJyI6UACx84kpBR5wrGKKtsKVpr+
wfoBivEUawEHEQKMBlGa45Kt+JVTDBmiZ2icKOM17TVppjkCk/z/UnJ25kQcfD0b
72MAUHTjhqUf1vbEQe+gByx+rPDESMiBtNY2Ek6zj1xzxsmeFs8P3BjaYD+zzfNm
31kJOhx1pCge+ks6iF7sFbK2uPRynbKzj02Nr0w0BbKcSUh+rfCj4p21Pgbch/qN
YmGNGCwxbMHYx0aE8SlSuykSQIFdIrEDlPQ1B2yWC61yN59oMy17S1wDUwA11UX6
IMCnpl9eIa+Q6knUEGSfdLb4vDTBr6UrvlPcPxdktxeIxdDNB2W0rNZ0QLq5hP7b
bejpswgzpU8+4kUxEmO2MVJttKrc5ZI6gjZUKItg6SsCth9plxDq9sCrC8/Tc72a
DhEQjcmfvSe3+93qjP1qbRSqn03UJGcVsy8jgkccVYn1bXZ3EdbV65VLscv5/tVK
6i+jTncRcm0moSbKIuCxN89li7rkleHnfVQHV/aVChTfKirdj6NdwTQqoZPRwNlc
WGXubeXIjt3K0D82nzZHT60IPmGuzRE+5G+8pu1OT/Gpt4X/4VkTvVBqKD5hMUuQ
jBVhxpEdRUU4qAhvyql8Refd8ZPMPX+XuxACRG+OI31wWQsgmpVFGrcN3Y7bhdmj
YsnIqXfhRYa1Pg8u/Fs8rCFWH2oOsCAeo4KkZahiAONew+RzdAZj9q29HmBQt2GF
TenQmUJd+Dt06DXp+fImz2iFTzl/HnEiV8/6xp32i/IdvHMSmwtLTWIfUeespY17
zlHcbCoD8ouIXzNxDEoA4pcjWvmSAjedzlz1wOb8I71c0kF6PLpr8qah2rLZDOZp
s/w5XOr9qzBKlQO2sCIAk2rAxWiO8ZknbFbkybgVfK/PN82juqCsEu1OPywMUj0/
WYg8CtR3wmrBpJj+oO2IVzuBsqPB2liM3SGpFklo1T5NsC8cBEWQhpZ5o1MgekSC
HA9RiEiL061qrtRHlWNn1KemXXxF3whCaGHDrUIx+lRM8vhhm8D6Ux/yWuO60eqE
rQVzH+T5QtRKR9Jr3drvFLQXR/vdfwdeR1Uvb0EqkYHRSph68siEuP/WbJ0c1Cui
/4hB9cPSV2kO41XbpiBoNzQKF3IF/4UC1AqsiKsGGV+FAFRofNo/M+yQLskSPLPx
2ONy4lDxeDJJXpS5lzvAxMFPWnBsxI23/PjbVDYeIccXaKceKHGNb+ZIEZg7bbL1
XX+Hr0LrNsmsNi6CgF+qIwhIKCgzny12rFnXhDDE+68Bjw80voQ8C6W7+qpR2+oI
oJweBQr8czEMcANGUvxJBfHamka51FILzHWVKDR5LYmDkUynlSEyc49JhfTKDW/1
CmoUT5/ea3cNZS85+My2f7jBfFBTyzYIsWHcRHnnRQ0ISu5WX/AjtMPDAvEW/7Zx
tE/uUYAHJI36CHBqe8VJ/5D9nJw9SjglOgwJecOte5SWvIEX++ygcl5bw29RKnrk
Mitvf3v3GIw3/M/bl8oBY92u2QERFoy7Lp0SpI4OPaaGLneQyHdFkfYm7+FkKqin
72j+fQ+zVLyviaA0ZyIFKm713C5m8GTHvLwcF3ltFGyM1/gi5Yp+UHXg8S9snk1x
8zmX5+HOYyO+WX9TFuqJSnSD3RDkmdAjVkjcRrYxxPfEcUf1s4Kz47txERHgV2nV
wfJuFRKBaIc7akPNkn0D1jYef6iNiBvM1tNBEQKK2JjqqTrGSKkbDEYVt+r5qExJ
GO1F0XhIQH5U476SU6vyz9U1Ir021WEvV42aDkD6uEBa6B8hacXx38gUKjYBWder
LELEUKY3E9ZmHBjl+z/OKtXDmj61BWpOtSaOgx+B9N26ZMvkXFbuQ2/8xyBXmB1m
+iuO9BwEJj1EmujiN77i8EGi4Yyk2/Gltzku9fuanqe3CNDsXXhoN1cyvyaIstPy
e7UdPKGuq9lvH1TU4K2/GBL9VnriBeq27vkv62chmn14VUs4JdK6C+kgEDcGaI/x
GvoRD0vN4Im+noFc5v4kzTJgHsWkMwUYxGMIS4KNj84uzXhBPt5CoTwQsCOM7hd8
ivsqA3rvv5v8lzSzfghvA8p71OO++JA+aaq/JZC7ogNZGedhUSCj1NwtjeMNv5Vx
MJJR5HSyxuZCt40qqVg2nNYwEWXzw4xNvByTxp1GFBg0YQsIaENvTNfj6aKAcEgw
FCtUc6X3k9CkqY690Pbm8oG/3gyD6mrdhJqpxR4Yw00Qzr/ZRQdPM18ptbsHiUun
eqcVYLXGbO4IPSoOFtm4+ujhhneCc8nynYss7FLWF7oJpjW41TXSMuyI1f9HcK7Z
xM+FI7sSrpSrSU3u3s5WOatCm3C9WS+NreXp13uzeNQo9/nnJl5fkyYPsd7KpFnL
Tp/Zm0qxYbSDuOJygDJi1G0e442pUH4kjpTnVMeNrda75zy0anCqHJWBxs3BGWKF
k31PimB3qPbVHVUgizXu7IppUA2g0udmORJb3x45lBtwhPtwMoyOPHV8/t6LNboy
nCRO+5dYH+EIWx8vPfDw3zh/3KMKVALGU0E0+24PCo9/ZYd//WYwCthCEA1piZk8
Lia/csAdVZEh+SW0LVXeQvbz+PzWHXq0HTKs9jb4Z+xmU1lXPkLa+YmC9hhCx68U
VGXwa+kx7n0NU8OSxfTNw4fJDZu+Hy+C0P33WgDKag3Zk5JNt+qrcw6x/buNeqO6
M7sXpdH0Pf1rOoIQ62iRvWXFFIpJh17ULtt1gGvDrFmZfRgryEQh/X05wZsEJqs8
HRZ+/FFIuRePIR6Rmmbi9QqqVvVbuTefld0GvS90cp1uC7ovcpJmScUKE2oDgOUg
CmhPGdulNx8J2orCRZ1mV0eKmzd5/wsaRj8mHY7P2dlRLAccrlkj+m+3xOAGtVW7
y7dVSCnS0h1qGaW0dEbi5dw4sl7hFKZosR5bKo4BFeiwFpaVaE8wcP/TtaDF7r25
2v/HmthepuqgqLHUCcNxYOpnpSp0WCcNTJJYsoVSVxVNSijTmXdajpp8so/0WtbX
hjS2ZwNsstOey02FTd+Hw+t1bjBOf4d03cauv6xWdc0NbUOuy3gPa5EfMXcaYzfs
TJIs5R/IsihekwcgkzU4hKczMfnn8p3l4qyz+1cZgl1nJ5eeBg1jDconsYsO/VkF
omqgEgHPlsAnbZNLeO8bVZKN0glNRG4WBuCd0LARM+GMKEer+uAoCqXKvZPEV9xR
/whByujZ73uMRSPaUUozMfsnc3jRV0Frj3GPx3eNjfcSVnNE2h25uNgVl+JXAnuI
Bf6xqfYczpHd7PZP+5O9UOfNdIzWVtb9N/Yi2t3WPGAX5IALUhTQGkVE0v6N1J4g
TbN+La7ZGvAgDbnNmfqxwORj4MoIuyzm2RmyJb3+uPgBirrRKt1MbbTJ7T8k/KU7
CxMIIWf+YnGbMBCHMIm7edCa4ccj4QvLxlhAZ6rPI+WYPNq8Gy8ARf0sRJlQqMwN
AwfWs6yRULiP8acYAkcKKyFif+idTWYgpcljagq9rIkQxzmcKDVzOC34DLTkKW93
WkGCcUwPQlPUw9jiZIwspiSp6cYU1mkWJz22kJTNEsqDbBoq8C6DTQGIQmh88DdW
tN6eAj6Os1qiVmk0ybJxnMz9vS02303IWfcfaXDK6IfMB4OMBtueIsCyZVkqwh9G
Naw5sLobcsghF2mNpPQbZUCIX9vLIL+kBGWvzzTCqtCqCk2vo/w2OV6R4V1ZDRcJ
llYZqPLmTxK7VweuFkD2EN1s9H2/bFKXQgUZeaEnyMRpO+7WoFrxNwDQzlbOSvNb
0CjFjcTGiHjNx538jUi8cVXJtOkMoeIn9lJw8bNZmgX0/j2xj/lV+t73DRCb1qLc
ehB5VaOFasapvTVxcHbj2DZS8X8g0+1DKyAyC8/sAuQVOV51Dy1nz1d/wpXN7S1U
nBA9gEEqfr1t3ajBh4cHjlM5fSiIut8ZMaJKcwobJ6YvuJCE818/8o+HipFBp1e/
zN+mjYcNxkdvDc7wIVfKKi6BtOZgFZQ5Ws9z0SDg0TmgjHUj0Sb/2cq0BHeQRc66
z17wAl94BYRW1W4PKTnxWjSJ/0mRshYNCUJgdFyU/WzfxPxTnQ3ERFaMdXyeNCXp
As0wzKic9PZ/R2sBPrxIO0P2t7JnA7Fghx2PoLKx/ShMDgA1CGk9PYY0KXpLCcCi
h9yTZH8l8qbjhjX1SNtPzXZhEgaEQRfwW8tNFLCWV35fjjGoT/3eO30c3tMB7h50
T4tq9SWPl9twT7O04rPa+6VGwmteYFqyayOfJ5w0V3+A4yLsy2mwLV2xBsYD0SJ1
O0z5VP9x/CsBA2OXDc7SJIcYPwfBKChKaWY5KRU3HcE5QsvfgS/9hYXTJFinNIsn
UAPynr2m4QsEdr6BEiMakjaO0Itw6YswFL85tOJ9hhCLeMhbNM5sJed8/e9rbRrG
o+6A4QfvCfb53AN6PF5mzvF829gLxwHCL9mvZ1kg4V7IDhEKxX5ahi/rU/FjRLbg
puSYN1AUsUPRC+de0jEt832tSzzk72VzvtSv3tnooIVVJqxvmWjaglasPoDuZQGT
3yWCR2dMsyCSum7fWpVxBNDocfmaWbqpnrwnkkyygHTxSgV+oFzRUA0bkGzIOvaW
A3LGSrZesZ8Z5UnJzTQN0LmjPt+C9X0+SdmESiTqSu3SiDUzsdXfWr4LGrkZtV/p
zsRy7crn6xDvPoVY2bpT4mwtuZMQsV+JpWq88Bbr9+ZO/qRAfcLfFfrP7SuUqIxO
7yA1AtihZd7KRsSL+TyFLwn1MDT+BGuUndeuVAYklTKSPNrBs4mGOW6DhzJyia2T
gY5F0dzblXtswkfGpUdTekiYUT21I54WxRmjp2Rn++xiBsyDJWzpzS4eBM/U/9jH
VNVS7yeLv74lEFQr1ZTxHK3Es6t5T3o1kxSQl9+I+cLVrYDa+/QnDydZIqTliRxY
e2wZFRpzz1sHKwIk3tO1nBZwqUOHRH8PWd1aW+BXOScn269nLF4If6w4aUSAe+rd
+lGPoun+t0hgccRUlonP1mBI669NA3pl2vBPOpt1dbu5lT9mUQvidbIGM+KRtDdt
YlIndY1o5Sm6RHsnRsnVMaZbiFmHPIVgpLrZjIeKqMvWkUB3FnOY2geYjpPlwCl4
ycF8+nU1ojLXWS3CTlwcJ+nElThLyPMY/f4XzptQg0YJ0LzkTH6O+W56fYmav5gd
+hUAZEKA3hz5GXael/0MfV+Uinlj5BxEs19HdyaG4XXbEeKYtkNtxnHtm8Se6ofe
Fc4madMCA6+fzlo/88A0dmsMx143AWbTEA9EQGPGoD92slftf79TV/0o/ta1HO0s
O8zXOrEYhYrQmfsb1Qwd89bLnuoVRXRAudJE6Fs45EN5n+04RWdbSZ7RuLUfyAF9
8Oltfu1yrGhK5xjlD3YyKI5V+8xlBNc2N7rB4lmxFTEa5TRPtUWscezwh0q29cd8
lld/MkTo3wcDAbq+U2DflUcXx5mcnD48LrSTRZAn+GJXUWk0aAFUo8D09+PcBLaN
duM5xlQTZ6slEnQzMn+f6NclicRCqnzoP6XKbLtiildLe/lDyeBz+E0e5LRUN7f8
Oc7Xs0SPG14lfGo3Lg5pOvSPlr7pxVd4pR8NDj3Pld5Z0yWlDIG0NcUUUoO7K8As
uLsZ6XRYT+wvZ6a5X00WPCR0OzHWXrzcP8+8HlH8TWQx+LIkrFcyx0lHwuh+Dk6T
RATyA7cWW6U/X7svERTZmsb9brthPejCYoczfILM3L64ZGrFX+0CoHSZ1Ytq13YF
nrBgCA16Nt0x9lGFR7AKoaiGWmmXIX5ASA0YkUW2HoqDGDKn1c5Tqt9X7NsXU643
iGoN6aPl7E32jH8ms2IZPfYROacmyZDEcBZklgQUbeeZxP9zZw6fNNUH8EQ2hV2c
6qi8OLCycelLKYlLq5A2HxdcKaoDiwyWHjkWB2fOT78IfPShxIGWit1RuTlI+yoL
b0HbtcZih9O4Wi/BXK6uMY8bujrgTCpJ6D21X9dK8aQNGvUdMRQKERc6Yi6gy02R
helj8j4UYA4bqZtXIkMZaZyh5lneN8m1/OqPbayLMsFhT24KNvRCuhZh8vI2sq3D
WBo46DHDsiCn6jPjf79LeNe4UnI1Ej7GYNEL1T2IOHDPimNnrmXdkuBn+TdBKUJG
c2x3+6fSsiSjrV8YDD6UrWtxlXL7tsbE/GzVwTk5uDkGFG6d+xpFsenTa+otE04J
iSSgNa2/Vj81DwPKRR8Ex8d4TFe8WeFqZdRXAp68EK5McpbQ5SxzPPGt7EsnhCk0
hsHTWjoTfMgbLcY9HGmo1kbJmjQ2p1N72fsoNrJtldkicdpu8sgJnYPiwUSsr4MQ
Htc9pokK9j/H+TyXNWBuwdnzJ7vf2snG1Bg8Ypx7X0DvcLWkAlu/KZS3jDZrzbSc
L0NE18ivBvgJXyXIneQFqhdibrNqMmf7bvzg57LxW0AkJKSdVH4kQ4cqGr7SLJUF
MtG3Y3Xp1IXJixYTbJtnVJiOdUcEF2rHTx6uJzph3N3e9momWlM23hhVAT5m6L2F
ti+VAMBnDfRphr34o7Ah/ZOFHCnX5BFLyiAMTAyUow5j0DHNh2XMO9+adPKWfeHm
dmKnvuCbnnuzLTz92YGUh/WtfnOc/g9g2SpTE1Nc2q3358kuKezLwE0Vtn3EbSXd
yrY2IFkGxDWKc/o5hsZe6fYrcgpXU2006qBVGXQCSJn9J1uERzvV5QVTbdf7xD+Z
w+8QvsRkNxJbAO8gKH/UZEVgbhZ0fphL2OZMpM4iGW0r+339r9Biw4KYCtq4fEJO
Eb9Rc+3O7riZQ8RS/mcKmy6RF/FSiPV24wRtESBjlmGA5OfDPAXgBZSOBvq3JIMK
C7CivIJTUOtY+ptxIeX9Y3iCNjsdF129qbvzI2aOSqeUdXx/HxnEXi4379s+DqU2
ssu4OVfP9r+we9Ryar0bSZJYha8m4yG/cSeIKc1BM2356H1aLyM4D442N0d0twew
OGAx/3W3ZT88sBCVk7NS5+mbjIYNaTD9rPa6JnhNG5Wt1GCnEaxc6a991NW5QP0C
BE4sm4WDpOc6yAHW8DvQr2KC7UvizKBerSEh+ZHLuyyg/VWHzps+SaTpvUN3Ksj4
sOraGOv0B2zLJ6jT1t9M+DAJ9JDAtLV5TC3AqFTVYVAbJn593G3YO1gXxaHkXoIJ
byazKLGGZIb20uOLudtBV2PEfv7pwKj8WrvLsKRjmeQXte8pdcTtvyWK+NGM739d
T2uRdoYZClJso9cxI/PJckNs+QR43li137RPQszxKMh+fqBq3nGXmzdjsJ0yDvFg
ydFqgB7zqI4M7ZnOihiW4baOjB5F8EMAvxpbM0yl+0bw2w6wDb86zARyMq/OfABw
EaMVXoaEvIRJcbHQFGDKNb7iTL0y4TtDRlax35KH2XhZD7ufYgkxewL8dRD0oKBn
GK7r448VftbMhZB9v0xGRGUMXMiF/kPQ4FB+GkyFaQ6hKmGdeEyGAmOzMVBuoTYw
RjZN821cKKuiXCHjWibOB5yWHpe9MhJgkFqiOPz/2PAnrKyFL0aH+BDKu6otHKV7
Ksb2RgGieYfWhbIK9bpylxipnq8bcNNZQGk8Lig2CUwQ2oDknI3wJrXZ3iuoJiKF
yRJJeySjSdyeXuY3wzf3Xu792iAno703BbzYMBRCEDezeB9U70+Eh/4jPk7COAF0
zQdc2FCwX06ep+TS5pE7AB6hPYu5oAcj6prJMKqX9ApgUlmzfxBUDidi90icv5a1
G1/5R5T4ApctlNaBQ59lBvUhg6r+0NX8MSL5YEXXjBZ07VUGLWjo6mqyIxdwOLMG
1nk9Wg2q1N8TBKfFU30oFjqXmBPKx9Qg8g1WCIih0Cx84Jv6Kin2e8p1bqF1u0Xz
74IYUfKPjI/pb511FVKjVsKe+aN21/x2oIXSqcr0jN2teGoV6H0HguIUaQWP7wk5
3xYaXEP6QxEbqt5Ei1zAmvTnGCHCk7eaCBt4R7SfOiOmqepZQe00ZZhrRsS1AMbR
xKOd9rv9RCy1HqTMuJ859zhSDwe656TBZ2yHX2VTwYNuZp0L+QHv4nsXiHB+/4Id
aY2je19iN4EkSnhlQtY8D9bRP1fKNgvYvAbCsyodi8Zb4uSKRdq3AvxwltPdYifN
P7KsxXDNJvqTU3wUmr1TdPgUsrC00YdMsHPYeOQRhipoTwJfxSR7+qPfaDHB6sl0
xsdR8aC7GGPEtsY/606ogu/8iStrK6Va17ZNPvB43nJweRvX+MGGcVXIXhbLRQTX
YVO/NSUp3tK/87VzMSe3oU6VFwJnpfBJKMzUZKoxyIuARfGgDfjnOMS4rgk0WwAz
vexSnK1dXKxFwhTc8NCulh6UEqmkLEODG39LfMawUqFn/EFDcZhbbXK5UhOKRtbC
iPq+ubacjUZC82BE0DnKTzJZmIBKn4MQjF5vhEGRSl9EFhyrN9sIS4ZTLCLcJNy8
JyLH2LdmRVXnW9Oqa60BqiauhmPHzL5oTE5+4knwh8yUcgZbHG4W6rWMCDSRNZDe
GWkK95SRSzA4SLfaMa5PDSHy+nK0NP8QZGA+rP2vjfoS/tKEBt3HhFUt1LCiHcnc
OjP6G21jG0DJ/7R6XU5tRVloGX6HqC35XLl92jVWNxAO76wIcPBzuVBujWCqPgK7
30ZuyoFUKl2QMuUte2NuIUKRLABmwtg9uKAsbUS6r2Nd+tBf4JoH7L3pstDkoggH
zoohn01pDPMhQvRWF8HItQCR+kMjnbKxvbECGCojPpS6yfgHiyuzn+CAZ80UCo2C
ADA9b9yYgDlSU+vjZSdxYk74xxZUClArtHcEUlhOzDLysyd2dhQgMLIogngvCUad
7tzjy7d361Usn5CvuldH2PbX6fo1cmxJ/hAL4kZJWqsmn8U5dTlJMJrkvDpnvI/q
/HscpH1wYcDyXwbPPOb0rRxcLeeCE0VaYAJhqP78qVA6kCaZ6uOgUh3f8uhCe4DJ
JoboPYnFLAHj4dkGG7TTK/xHSRQsA+JxbTEVU+B1CKAHe5z2lgKJ9A0ESpijkHup
jg7yLpidmYgGjM0bJvd/KLLxDHxWeOqqf+Y753Tksd0eaNWInY7ieorb4J2wK+Xb
Zd2OoUKK1lQKqWQi2eLc7kf5cXKeMxTKxiDsTkWyBf0wIFfJsrimUrRvFVDlrt/K
TLzVXk5CuhG4i0pbKrnJQwYVzJH21CxQTEd+JQcNy8Q8T/aP4bLTzkypUkc1Ee+6
Y/o4SRXOAHDiVMHwRs/G6Csr2hZreOplwtze/x+QjjPzdFYWq6YTkS1Nbb/thuk1
oVaTfITTsiuksSVZu6L2OELHyJNZRCX7Greaua8eP+2QvvcsKzy+ewOP6/3RNBBN
7ayqIpWPwRXW6nHwpQu/ORJ0k28ClBFyNhRtgHctvZkUAx70DfW4EsCykMI39pU2
Yqk6CyWkEREbZ8QGHgkPjCxatRBn7wOFlR1EreiTWBvRsoRhNoASHbDWuzBeWT8t
EEIybhQ39KblyH3/MKmmR8W2C31OvgMLh05nowD8QupqPm1H4D79t4HRPMNREEK9
mAprC8iwtcHPC6kw5uZ9LMxV8PAIZe+mBzDX3MAEVXegRObXXIF1J3/bBV+k2RBk
CnV1Khkwtpq/KbOa3Sa8e2dy8mSN368HYw43ZRrpa1G1j00Obr1TaKJ62CGFQBU/
ux5QC8ZB8ZO46ekGL0EKkY5APm5u7tMWPC2N/vfeg308+MIIOFbTk55B+fy7hKGf
cJiLwGZ3F2MmxXQEk0l8RWwHvII3oUuuL8uimGhjAVSKoOLvue10BTy+FcWAImKB
QEr9C/OVll2BNEoT/vSQHxEjBFphesWytFu6voKQfk9OteQqP0cwgoAe7necMmEd
PCVmVIpvBZ/RfOc9FInKh2lOIFaLV0I3v4Lhjsn1FSUax46rFyPYcXKbGo+Cv+In
o3XElK1rCfn+beTEc9czH8702MuWeG/IPSWP1zFHnqNuDEr6P5EXaBz4s18fVc3c
OVwFsFVBNPuLkjtue3nQWYDHzZu8d8Ir5/evOfjXWe016YkUOnDJay/9HWVmYHO5
VXynOWZNkLOkQjtw2eMHBJz6tADwcnUNpLTxaJe/gtRR5JCGWOKG0CDgVGG3smcX
3SqYj+QNkLys8mEYOCGG+ZK4HwQOe2qVqpxTzr1KbWPuEF7VB+bYeh8IdC5lkrdo
Gnn3ocOLG+gynLcLmekF60qJLaKrmJ2eb7f6tLnOoZecbTRhW3uMts45HAiw+FEt
Z86PNtUfyP2bOw+xc1c34LQRT2QCoFJ9Q3t3JnzSzLtrXNTqx2T9U6K1IRpj5SlY
5L3KhtsDPSfv3wPhaVrkx9mwnIfd8SbLECeLAHX4C001sKljUObaic/rg4Nj5b4R
kxU2Zir+1mh/Fv2p32AxtXyJOu0A2JyMqMf+eq9VYc/IrezNrM1CJ9LRm2vp5mE3
V4U/FznGU3rHGr6qXkTKCW/og0Rz+mnw9WAR1UWIJFZzdCmNkOXrWsHriG5CO2UV
6zemTqy+6TUefHNald7PVtYOA3i3aD5fyNnCfbaiY7UmzUI5yV3mEsVQjV9/KcLA
gigq1Fm0QPwvR7+KryTtiQZLZBNOnKuo4h5yLIlRyzV+OaUG1PIcsb7MNCOYCxjr
q44ON7oJqIqIFK2hW1Gt3uh6GBGtnDpFaZk34M68jMPqe7K6Q1QVT3vvtlkrcs3H
v8WTCO1eysV8Z1tB6amX2FnkPOmk95Qtjy3ktPELHBe5QXs6XczEcHuw8vc7C9EJ
RKzEqMUFWufLfBkZM3Fjv+grQeteqDL5S1TNXAdV5eut5xejhhpazrkGG2ZjWHmv
ICCiOA7iJRab8g93n0VWD5tdzVN/z+QaP2/vLg3GCiz7mb/MbVAI5Bnz4oraFaKv
1MsArevvsUgxE6u/2MLF2u5c9dkGrE9tcrVikslDwFdFZSgqjizL0VoL3DsT5Sk3
EoO6zcHLPmtB1RcDBMOK+GjMUUvRRK/x0yTIA4du6xaGBTP+XtjcBFkarMvalK5j
SJrnaw4Nu/Ok17HBY1Pgh41aDHQyrM27dpklBVrRGgeMywHiKNqOl5/oWOklR+3q
TOY8vUlSUseYFM3IaIV2uNx/43i4gKFAZB1S7skywbNyGeiv1ixS5I1kH9bLiDKT
E4isPDMS5dO82by5pPIO/UHZZ3WMex2JEZEDy+Rt9Fw+TsBQgL7zGWBna4KCoH1v
FvpTUPiQS42epYDonbZFbp4qM24xM7Xip2SKL7WurzWX16+tmhdbjKNJXHbuPWOA
wT9ieAx6jnodRoUDDMPAtMAJj9rBDKwgOxUppOOcoOEBKak9p/3tP5DZEgyuRbuu
vvbqJLdcjbJ8M7hlkwCXbkvUiRwfU7l0bjJB0ZFvq2n2d+S75un/gYaiKZezuDa1
xZp/+1ncBlppdRiPzpJ9ykVCWDmf73Vp7SHHzS3rDXxVwmLzLVpvMVQWT9IsWfVC
XlCrfwlMAzRzGlLgydFtvMuWs2/+LUEvlv+j2QkgdufKuoAna5QsH6cgmkKMQVQS
8/aEUusDNEmsmVVxddLu0Q2rAo9AvII9bvInsvkCmTCffVJUnPW6SJEJ5otUvRxy
7E8XsLYsF5hiceUMHHQhdatMlkkk42x+jbs6mxJapyeo2PgbCHCyPselkuWihDue
mwQ3juppzm7NXecnrY+CZsXfawZdjW1QdzyQ5kWXKo8IP/rGblZqee4V6fPoslwS
8l0LxroSDoJ4lBhezPMJTqmHFt1tZU5+73Nn0Is+a1SyNaXN1N6XPZ8Muois6OoY
n5ROzkJi5YlTFIoZyta04OeYsyvqifIEXGCobh2m5dNwG8taIFr+F4HQBvYNVa9Q
4IdSvCxryxNo8C4QMbrGK465x1LnscyLKTXIFxT7zUjfEboCSdeOML9yhkY8F6GC
R7wKG2K8ksYCyBaIpbmTEQPaJbfncJ+eWDFW6+XWz/EnpgbiYRcF+/3bFDQ42B07
XVOlJVXgFefTRD5ERmsvKjnuO29bgywQXjcLiBGCRfwuGlHE3pLL6yuyyGmhTtxP
JvGeSguJERg4aU/ecgCC9IlJoYlmNzeiLaLJKjxPvRJfYCYOxd+XXuVhj3OBRRL5
g9K4fGL8Qmk/dSBKsvd6cj/YkL0rZzJiIQWD/UmBUhDcaG74baKwd9eI6Zo4e8pw
WEvuMAqb93DEVibz9W4OUHL2v9BWX0Gaf3PWzM9TmyV5nokuJYt7P9zlenA0qzNs
lQOmgx63OVdecDPd9VCZu3LymWeKCnZz9S/uVC3FzVYqTP+XH4D3a1fHk8K6xwxR
c9/LAg5Yd+0skvgNFA6jlEaC/Kfw6IBAnDq5rKgzmTx56AzB/EEgf3OVMIcRDKZf
uP2RvOqhJ4tyRVkiximfxLTiqz0IAU1HQJhNeWwmoJb+NX5+/VQNjiwVP1VevX/T
Vp07dLSZod/S/Fy8DAiYfqopAV3dy6RfSFh1YKzhyyIlaEOC/TZ/BM6zk7AEetNV
270jHBEV6ZEN/ZymTPNVEDeZsB6EQTJwAV9k4006VqzPnkhRb6Q3MvD1keE6DSOz
6QNRwEGqZWDdTlEKVWFjuggOWEdTpvn4wS1PlFhhZvENF+I+vw42gbp2cqOZOYhM
IxBkK/rTYQnUSR6XJGyYiyPJCsswVr7XLgyH2jvr7QcZ6KTQklQtI3Tze7po73Ak
mrEFA/8H95wFBGP7NBrFkRFUqZMZJZE3W8ysS+xjRZbaWezRhkmBoUvmzmpSMxHh
0qFFlhLOwohmX+CtGuWuqNaqCsCr+3sbdjhxxXBeJp3DUJjy9/Xso/CnSL5FDD24
WrYl2RKgyLieqs8Et6ym0pe8UZX30fjlQLWHK9wKLrZ9b/Qszeg1ZRbbg4BRdXjx
4QEr1StNLokt7FhTah9Xtwqp382wOsoy64z/BINQP8CpiGQdUxm5QekOngQbawAk
sPRmIyddJaCqxjV1AdnAhUvM2ZpxpbLyP0nUC3pnV90lhsklus3ci/fAxRIfuSqV
17Ikc7MDXm8yhDSI5jrUeJJBM6uWGUsdHgsPMVxJQ1XEie6lwpKXtp4oysn8fD7u
0MEtHwb7brjaXKKzuxLovw2Wh4c3Z1Hy7YDB3P1W2LIrb06J3bdEyHbZG8JvEDcA
kEqvbstnCZxaPlwPwbCMeVRokLkpobcR/jmFw7t5acyTewea8cdAxDBEEy/kCUyd
03dZ+eqcZayEfRbU51W3iEQjsaXNmxJlamXrMLgULncD32GuHCNJ8efrN/X/nyWH
sl6ZA4L6yeuGfBPvuq7dr9UEkjBxBoXdQJk4fWuPhtotSlkssZ4DIsIiPyhTuTw+
l5+ocwrFXXGDcaSvnu2CckUZWpRGEsFgzZS8VLBU+P1MMc8vxDicPBk4pNta6N/q
gflcDuA9RE/JBOMnOOOJ+IYcUphek5MoIZTW9CcH3noLr2xgugf9LvIjzgx2n5+K
KPkmE/q/ptrJQG2154rqMRg/dUd9JqkH/EOq5dePKdz1aHloQfH1570ztQp0c6y0
WFydZWdHyIILbwXAA6TRj5UwzUzRiFQ5BPXfkO0rIM45b1E2KsfondajGe3vloFL
fmcZcebw43Ovon2+nd0duqNwJnYkIGcN7mFBQV6y/h3LHrhuGNRnye9aREG18VdD
S9GnRD2SidKnWoh0SIRftGdOthq5bYmyGUwU3btMdtbOBZmh74fPTOOLnn6oGjDa
2MdgCMsuO7cBaXX5+cDmGIJY7cSaM1xmk3v8mzWkUVEaL33z41dMri6I6+m67ZiA
dWp5Avk35cC6q/eUDb5fhkXLDqXqUp8fCQGGC+3/VGXtFS8fPb2cfaw76aieTPAQ
HBJ1U5X4CZ+lcJzaNjA+ARTvcFS+oQ+ORiu2OeTwB+sSY/DB4XhvdYcTHgSOguH2
/jHhg7PCeXI7ZptzF8QstNJRkpQT0Y1XQT1aV/pbsbEvBNArxBVzbOdfJ/sFmt2+
HRb0BYKlSDaDM6G512FTNJVt14brGCgwRS6EoFPVyOfjRNTqJzeDqcC/ArlBPQwd
h5jRpstkVU5FTEwBKjJTSoxeoisL3lTIsVDXGmwf5tjdfucBH7T/Ch1jxRGn1WkO
U1Pvdoj3EzbLgUGkWg+n37oTKIw19yoMgIM14GfjKgePeI13jAMo4ZiDcSWeZ48C
jOE+hBnAM3tqr2mPC/r7quZcjdUU6A5UiDauYJgAtke+p0K75pfN6ZqDcKJIVPzH
/JhSZGeONVKBE0SdPD8fDiFQpR1pS3lMs7hVHaPyDqHFih4EBGyAisugP0hQhuQ2
Hrw/6KlNpvoI4KF1gny+i3cH184+3tc4OhQ0BCduYWqHsEMW9FGnSx4xyUrpiEbP
6cUdYzgtPtDdTixxt+in0Yap84pk5jgIdI4Pr7LMZYVsKDpUUeexDHV+DZGeGEyy
U4FZpnlzJt3FbNh3tl9w2B+0omLfWERuzU19tQIZQRiLKL/b2gz4wkb8f/UWRFWu
OCivzQoTKdfcbOIqPFJvNQxuVlZIlxLlv5nQZxENG9/s9nmB1fDOo21vKREuoI+m
7Eq9Ma0JxnIK3nZViYTtYbj0Qh4FuVDaAGygckfzOZ+3C12JCHVGv0LFr87tOXDb
Ii0ZfQDSVt3RDZfjpErpxlhcD+KFxeX5N7BpU+Pi8N/UCjvfVeKNYkLXdbRuuSd1
dwRfs+Kv+Anrd+Rd6mSAUIGvP5cJMrOfL1g6eH2G12j7VInl7dFAl33t7a/Keitf
u14DVpBrk1QkG2tpxpXhrtWDPvbMZ04Sh2iTL0ux/v/X9/aUGaPhuba5SXB8YVSr
opyqEgwFNJVIaeWVdmE1SNZNSspqyo8kxeYerDTIj7zh3n8krBBmT3O4no/ip3Tm
1eTkz83UlmBUOo+7WWsf9+ZgFnG/5yOQGs+LZ36ROADeR6B2OOgxQDFDwifqGONk
t30bUekQ6OCzO3E3QSD9WE15TWDE2oqPbAAdgHlxsBR2XKgQbw1faA2/i2nX5LLl
kiZnCeoTxnCDL5Vu8MZF+1/BS+sVs1AxINkvpEWH+09KtAzzp1nxWZKyQLPELaXB
emoM7cDe8M4RLp6b8fA4QZ8eh2xnu0IvnPoPSsH2gg7g7S7RlvmWLjbVsGc9VoI4
JWkHEIzj/Aqs+BLOjKs6nzbOGDdMVt155tCdeR/SrIL0pohivJpJGbyVt8p9woRU
2mOUh/CfwkFuUO4KTGizkSOeBMuxvbxbw6R+P/WN1qFnqsSaJ3k0ePtwBvGIbKuU
qm6jRYQOwpl7xuuLcfdZEOVCgHj/xsqxA8E1v8r13WH8ZASLQzcN87DuoiEv5O4L
PKmvC0kKKHWMutmdQaf9vWgZZUdw5LSdkC20IYnMGWUgS+Bak3wnnMAJ35piQpBb
pOxlzK+KcHS4xLZvtXVxvcCm7dvQQF9imPM/vOlRroj/9DehIPoELEzwmHOt86zq
+yWyOx+/fThsyG/8WfH7jv5X9UU51YH45EncHg5ZrqkrxIMRes2pvLz3DeUYhbne
E4+kQhBu5xk7eOgRLFFRKlCzvh7qCmBjReNzezvIYr+UG8/1i60Cag775TB5Ncji
vNcINLvtOxucYqSmZWSc1qu+DZ6FcQE3bV6rjG3tU35MkrR4yvpz+A0IHsGEAaa1
HV57/Xrhy+ZOcAa9JISda6QA+3wJEyxI69Tu7aoTTinytlZRXBGGgLQQcv4kHmaZ
VpPbELmL4JqgWJylERbM8lWZfUXnEX1rgUS9A98t122U0nZpT1oZN2cGOGIZbpj3
Dm9JdanyC4ucVuEUjfirvPgHPsFxhstxerOU+AAbWKGSog3G4IRgO8pHl4vTKPPk
Z4Zv1ZumjCUrfSiGD6onFQP/U9X1OwWn+tYe5fXUUpcIIwQ67ivJQOMCcA7DBHGc
ISZNkjCSseUguTUFGc5SPdpXawu4906+Q8Qe2gxIUE96gKHzEKGPasj+n79dYCPr
wlbnnfgi1rLjwjaDH3kamg+8JZVyEW5lhqcKnLEYGLtV7JwOjpV8f2hHXeX3+PdO
2ASiQTJVV/T7DhlZ8C7swg93hYZnYrapAVVR3Tg5pGZVSKWynlBLvnol1AuiaFEV
ckZiVF9ecknhTB8l4/jZOwR56/lfuTlLsmtpWdRBp6kwNE4IxcCM5vYCYmQfPpgV
QG0GWCVwPpoJsVhKP9YrsPHSDZkD8gBkcpDJ9ZiiATLM+aW/tYi05x2kzvvaBWlq
syJviPRZoJGXNHqJobaW3C6BB/vPbXccAT+jPg/VFWsX0y3CIGS0oL46pAOf641K
H4DM4f4MFh+PLg9vaQ73xA/3a4Ztix8XTR+DcH4VIQ9gcN9rzbaWlFARz0BfZYFw
t70LYeHTdQFQ5FmmjpyvgtFsu+LYRZDAOKRpjAFxnVuEcXFXPWW3aEDj3JkFgkdh
AuY0SPC7liZBaodV/Z6bKvXKEAUZiuUxfTEUjRUD7KPmGZqnwyB/S0/mRHrv+RRV
GYbzFwF1l0fwYrhDrJmlZmQgs0kGRcmKhq8yQCiQWIyIdXyxCYWZq70cNatBLDfd
xSCOVEh6K2f8qdCD+7wyGN+MS78opxjqp/CmGMZZKmJlKYmc6vFrMFGvG/oJW1HG
2FuOtD3WbOkfekywmZ8z7IwyDPOKemiPHdqNhDt1eSHoZHj8A0pSV1trsN9+KByw
aszahtoHY6KU+5Q6821921+5Og/F3fB2vDTFXeli9iTjSVPTDTmgucqKRSSZJkna
q8Go6ysbUcn5dH2WrVEun2H0qpMFmlWAsXXXJOr2rCaOAWRiWxCo2qcqjt4Dks3W
qv2XZeTMJnenmv5+iMnq3Y+DV11lLuH89HWx9S08S5Bxc2zvCeI1DCy7BAzcz/QD
pJ2Up1j8pWkJWbWH175sgo0xSb4SMaRjsyTefuLa3948qiV+hZBhDvo2rXfcsoBn
1VCfxE3k7IFRuvhfMPznMXt1IzfgxNCHONx7e8qQlNkovqJy/Azh3cNWIy+tB10p
+8fcsyW8eCTux8CwmWVbv3Qe2N+PkXYW+kdzOYRrBROW3o3d8qQ7TAkC4cs261As
VCVKYeJun/3hbDvQCOhWqvv8J5PF0UZym25eeteQzoCTwUwDwE8k4O1bsUZpYSHZ
yr37B0qqLDl2Z8SZKDlKi/HwFyBhu6cIXbRWRibay5z+cjgZ66KtHLe6uKI/KT7a
CXXvIcLekAlaNjP7M0BL2i6iP4CZ3ZHkvYuQwNDL20/optxGk/2U+fseRkSLWVFM
nkbV6H9aakoTQKyc2S3T8FC3G36kQLbEztQIy+60LskHE8rOYocPDSxeQMWPO+6A
38lSO2tHdu9cTzLeUtS/fZjF3KzrRRWFccQiCdQj1ZTWG7e3dAYpglP+FLHQ8fsf
cu1l1SLlNtyKcvksOW7lIq8WFQR+Z0zQjCmu8If6rhFjlKtoLMqOFqgsTCEKFAhY
itYRj3dNCZmpw/4C+dFvRR3pZNVGR0Tg0QzQGzrXRbtjzPCiX0yQk8OgAsRsp5x2
Z1xoFZdWO0GR+E83EmL4amJbLS1Cv/CePyn6JKDwLx8mqvKPmHoHRwn44F8Qk5Hg
q+QRZ5nLmDg+TqoloBkTI3K9N8yB16ihaMrGupHfvcPjkwgJKxZA8Z9wI1lXaB+z
sPmJJ9aBk2Kl3+3CEkpqotQygKnnOP/hr7+BGHaWVtpVgGFGuam4l5/yo/5Q6J0c
XXwBuKyrUxARgj5D4K/1DmvGrRO3iAXlObyorB8vBDBDIeBsMBd1yA7aI329Zek+
3sEBOXIzATRl90hxwQKkyPqin2QLp77H5UyWOUzATk3/PIqncSO1MrVVRNGOqgF5
diqQsVxKyY8+W5vfrIGfzSzKtRJmyvo0IwrDpWND7siNfn8t3qq2RzANwNvbs4Tn
cfRs8RbOhGl3dgssFUsrMB2ANEYYLXE7H1HB7auzKjp9oJKVJYKsunVkJ2qtv3L/
qOqwgUwb1LSXHqoVCG8CCUUEGC/6Iim0c9VdTWZhkpirgBGjB4kJcgo3JgKmXdTV
jxKLRs6lrHbdGkIuD6WWc8ADN0U+YGcpX+pPmhSH6u4n22f2auHOCVv1XDRqk+4z
FpufV0bu6ASwKjccJtGmKgDp3/mmJ1uuicOOUsyKnBrBrdwJVQa3BmmVLKotIqmk
97b/8BIeLKlrabMVjMckznRqL3WaEHbHxkEIh9ycJlTZj7+quD6CSt4OThqmASZT
C68ztC4FgiyDZoQQlxfkkIEUzZbvCnXAYLEKrkzcSJkcxFxSDUPnzxKFldcWjD/M
Gv3w6awmzpTw8WGblWwkzlUAe7pl6j9n7KPzskRuxg7h1QgLcBNn3NB3Ngv89ri4
g1weONNTNgMejEbfsjLmCiiBTL5r4lyaNjznWkvMi7KA38oyIW+pum38NUrhbV41
0wrIO163+KzEskJA2qBI6pzOyI++OCWOcoOn5BkZCGAeDWYLCyLW4Vl/mHXbYGEI
f2y4s07BVhl9jPkmsl+7C7/XpoPBK69je31kvVz3pGZ90KxIqp/fXxr0Zhez9AxD
ieAfrIf8GN17ygPDSBrfQeXUEbh8Ppu5ds2kRELPU1nS9bJDgJ+Ayb/S7+RZ5/Kh
Sfj3d/NJdpgKyBH4AZWZRmfnipcsBSkWlMYBNpxCOJq5cDQty5RgR9h51MdQKOxf
pE7HTMZYBPB/g+8OL0FhYMo+km02mFdQXCsrdkWW7bYKh1PUyWOMbuMSmlXIRMFr
Nu/j3Q8Gt4Y7euNZDpiVoWtzA24Gtho2RCJ1UVMmEGdUtwvVdrnGqM23kJUEBQrc
HziqVg2+xjyKIIlTeZkY1DvgHwoyPwguRKZ7CjtQBI+c3PF0PJ6lDlMP3MijOWSy
2NfWXOUwiJARXMfERCbN7ksJKOMpukh46IsqskYdxUPihhZOFc16+4qyQ++cT8BV
o13ms/LjlMI7GBHY2lfLuu66Dkt77oapLHtyM/5aOsdwub85DQYuNzGK7qT8btn5
v7XyKtldgfOCMvfurREOQvcsl8G1HboIZAO6V0rwbtiBuY8qmK9rjxYjd8nHmTdl
H/yTfGxengCU8EOBD4qYheN7NDMlR5WUBS2t56P9L/zgFsfGw7bzrlyuZwGXarRR
4jxhT3+EinKfU4pyEgendJDZyT43pUGJv3OFycJz91lLbfCo458/S90Gx8TqKqj6
b8R3on0fA35RMplso14yhJDGg/0I7l5U5aayJTapXvmuW9BqIIUYDE028PWRT/oa
TJEsXNaXuKvy2JoG+sZk8aa697RgNq2V5kxjx71XAZqbADpBKiE5Cf2iZ5GbOGG0
Y/5IcWzj6szDbDfj9uUr/493o83VXDPgLJxOTNC/0e+FwFHWrGYSGrWw+BVkLlRY
zK8szA43STob8oxyvXslBGghM3HOAic85XIUagucO7LCxutTWrWd5gWngmttyY+K
D3WABsNskFQR1wkSYH0Cv+Aq5bYcTnIi4GrjHz0lV+nKcInOSyBx0efq26oWpY4q
cDOmUAzADurPge/BAH6yhHisxCU3BLbG49bW8Er/UQcrzlAJIN5kevmZUKS0Cg6D
IhILgRZsD9w2xwjz3EORG4hV+bmmC6zbVaCKJSZlIczoLTToM4rXvqvvJxvC/d+I
QWIN7WKyLn1SahcK11Y54PLrJs3YJikEvLii9VKfv/4gonZCrNlQPgCTQmY81ojZ
dDkqiulMUkkWCiTPpvwPlcX/h7Kkm/1p7sy8Tstcw5oJ5lfwXh9F9JiTWY1ZTrKf
Gll/rEXMNJXLtqjHJwOQXZkOZwoB4r121qBvrlFUBzRdVKz9Cm5BxPXGQKgso7no
BbJtrevsdBCvr0TpV0hxF/Fw1gHwf7vxHJuRD/JC0DS+Q1DFFu/qHoV0ev2Tm7GR
0zUQ5JnNEejHa/1Vmhh78b+76hsHIPeREWbqjPlj90WnjADdhjaHrB0lRM4W4U9g
dSwzNAff907YsaYquYDzN5C+yaTHQI31ZQ7LlOFgpeXiB/CzEoFb0yHHQBaiGXyR
JH/tVTg1+UdXe6BstpSR47SjgbtU2tqdg7+Mfc8kMLCmbXn+SEh+p7uGaJdtbHp+
oLaZW0vh0DiMJWAhpMqzgVRtydS/EcvWHI8pVjEnbxUm+sjKkwlL+d4HJEpEOlHL
BUmwRaIlldFBzFj2el54yjYCpYcCVT/8r2os4K1oHk9fU993p8sJRIPKlfA+8WZL
lF+qCg+UMw2J0cNgLU6TCXfKuE+Jrlgsm6oLI6hZSXiYxxzTRfq/UQ91SyXoJlce
98ROoFjOr/tTpL8BsOoBYb1P4ejLGrIS5w21JfeTXx8tFF+I/IIXDlOoKgSLtzom
BlYlIpn5reOxAh53Ki9yIo9q0uOTPiha8l2+2aiPgOUT+Aiiuq2F5eW/zR9p3+sw
3w1bntCRMSVoJ1UVyK6KlP80hl5WMKQkPmKmP32vJbEQCeFu0ymAGxM7wNJCCsfQ
nXdAiuV/1pTPptEmIIfVdyu16SVboLY71adk8oFmxXFJ+SuD0gjcgupf0g52bE3B
/W56J2QksaO/VZHEc19jnDAnXpkp+gC+TY1DxPBAdtOmhKdjTOhV6rj+Dr9iBNA7
UF2vzLPBpROitz0U9TU4gAHZa6bvcdIwAvBkdk/JeEjUxcRw3MZ+oO+SQJwsyCUe
OxbzgPAWPmBd/+Ss+WDRNjwVvu1M+JC8wT68jK3zhgpI/vg4Q1otI62q4lW66U4X
dC6bb+7yrWxGT/v7ZkpjovVBkVjr+bv3GPWuRCt+lwi6GB8PGH/3YbnOFR1O1C/l
jg8itEL2YLbVKwOPh37w02OR+aPxMEbmNKiEOXGFYyFFMRmSDekycuvNeFVLwlO/
GXTuL1k3uxv6G1mAr5kQSHOiPc/Tv34FkR8jyZbAWL6AuFDlM9N0UGVMFK5+Vjza
qAUFakHwufeqBkEROTlu0B6YNXYTd01AvB9UXvh4eo6mc6yQIrEIMD+qpLapZ4ln
q9+fCWzLDq9ikejIzjTJCFSUgg0dRjeuT3l+X1vJzjCR6eb7U3MyKW1dXUIvDZZO
7S0FldzS9h5RUkuu/7r7dkyq2DpzGdl5OLZEjg4nsFmY2cAWTPNr4+JNgNngcCPR
C8x30oxGQRAynqrND3bdKk8hyItw0pOJYoC/VqBKeZN6nuGxw4NjteeLTgKuDme3
L8vutVyuydFgjpEc06q2mnb5v7XO6i7trejysAynnWl57jMm/kanc8OWxtBB0I99
L7Jwem2TWq7uEit98Y59SrJp6ssW1RPzxHRIvJOP+YrdF3LMnp2E+fQNQUMqqlDM
b9FgBMWyQYLRPypZ46UFcfgL1kLtJRZHz176EQJ7XYAlJIYRApIyEvpUn00j/cAf
8VyxKjiBfddViEmqg5arxPhCQNPu9yRnMFHfLAcg2Ucxx/iadA90x3ZaUTVX8eK0
Pub/cVZEZRbKjmaVrefgu5m4QLkbKugAgrxqlYziRBjIPKL3w8sxi196Y/dHvGOH
HoHR5Asy4MO+NNEGpLCOkTO5tQeUrnKVRN86VBJJcpXMbvZV53BNFmBerYJDCmdU
bYG7flpOrRUynzUGMKKob03nfCZM1ZsQzOs76x5iEdfI671PMUv7P+q3S07uMtds
1FZd3eKZmMIxEicgiG7TLcQeJEzEextG3BCoYWFIKlAD2oOgWc6CbuETGzTSCMii
aQCAvM9571IbUIoLOCr6hZMwuRR/EbOubkdxm70Unvo8132I7VmPLXFaPGozlO8P
5D39wqkhhJ2Gp9csuNcwJZRLFPK1SbUwRjeLAF6od0q+YRVlrlkHVGFnfVOPx+S+
wJW5NJeirBD83eeUKHC/r5e0kYTJiJyj5b5Bf7oRayUy12ZmwJEXgieuKbDIAYk0
laCRSKtfgzZfhr8NcE+TS92DgkBqEbf8nMnwOZMlv2sIxpyFdLj7gYHjIYIE84lL
feD8Qv2GPvqtfR2n+St5JHHJO9uCN6vO+5l3QE+ck/jvJHXMWGNYpNYrKK6qHQjs
cVTa/+i269NO/wHv/LOdgQ+Pi/NDdbFG/sKNJt7zvhNcKvy36W0gKt+Hm54ojfqE
kI8wj8boTg9fGMswwvL5kpCmBJyVIIQnEvcUcBWV0GQuFaSZwcVkKsFqJHUMmrNX
x4C0Lsr/GQ6hyabahrOpmhvNNcAwvXbn2gVA2F5WhHT2V7KIVaGCiHCtdv1en+jV
BwrCna7PZQIooYXwCV3q7DaaBQ3kClvQ40KytBxrYbblS4KUvTaq/H72PHyZqMR3
tjm5uAa567FVRh5t5YdeE1wnxK8WiYgZPwcySMeaUuB7XUU+4/3LOMoDM3UfY5RH
oMN9sl8XjxglsFfxVecXQHi+UsASQe66OiPrR6Qe0Emiu0fRpLgko+SAA2XU47Hf
NoNWgIYtIKJOIX5feCavVe0fpmhjiJUbqaGnb7zeW0TYD7Rz1PMpjdv6VspfpNkm
R1Q+WLumVMTviKx74p0FHxRyocirlWQVezYr0QpJLtIBD7Ss7qmDBDANZBp7J0e2
31PJWLgpeLAYuSzjL9O4cRzYkyepXpEmJvpEHK53lmgRNjGFGshhBblOoYsF1d+E
bG7JPhwEcZO0UgnbMVTtXAWs0T14BepVpHHCL6VJnHNRLjm4vv73ZebdeaxflIZc
wRg3/2X0JJZK9sQWT2C6YyxI1il4d9sGa5LhYRrbNPBSAFpVzIABwujqrExytel7
aKy1YBePcS6fLNv+bQ81E9CKY5RD8zm+ubMRQ4KFnuxVD9KHeJRcmnHZVcQ3Uh/s
J+OZudj9CR8lZUJ6JfjyS9mWFEurPT4KPuDI914oBCLZKvpfoH1wpGH6/g0paJMK
obJ3nYR1f4JQtHMwTJPuviUS1EY4iexSmYGnBl9f81wZX316QhB+zvuuPQJffqbB
AGLT8N0J6ei79KZqHo4v+zvq0dYDKyIX3HIJlFr/mq0p5cgALYk7euB8HcWvzscb
xaE/y4as+BolUGPfMjRrwUw3jjEnqiWwSN58qcwhLHktWZBLO+lD+KB4M5jdCAa3
OhtlOBTR+SZhXuq41LS5SowTSvlRMUZNmw0LioF27iNciKgkbNd7hEuiDUeuzABl
GUjU7G8c0PWSC+aGE6ZevX2woPSu5PPl65tg8aLjoGwP1NFvy9n8x/jpPzC9Jld9
QMZN//A2Tjt2LJgdUviGpdUi3ksjqGmOGVfEgucAXoZlWV7umfH011kOzM4PBy+k
QSdn6vK9x4yt9h1ErPW60JhUfVh+a5Ten7N4zycL29FErkYYj/XD6kfMXUhU1WR2
5rC5Ge0nzmdnsTSlFGGezMr+x1sj2IDMY42/87VnNY6htbbU5Ng9Fxt83heSvmve
R5adlLGMBrC1S6LdsIDwZf9SShY7drzdyd/xf55IKBkWQAwl0SJOIWMDwW4jdtG5
2hrHobV0P0NDu/WQXn5yx+SPjdUpLkdWJvU8l7hs8qOv0hQDvifEAAfYGSv33mSk
E21GJeqlVbjg2wEo4dpsEt19Vbiwd7GMbAdaj6UCMFR01jhicnXqf8XH8lWRUXNE
iv8kGX7i2kq3yePW29K3QpjZBBui3M+y6xNu+0ZEZCKYrEx/i6hd+8f5WpGmmRuj
OOMYvmMKdxnD00tOBmgbZSMLVQvphs330ezEsedv/tljcdnDUXn0vTQJNJoTQWIr
kJQcZZ/UxHzvNzjZ6SkrcqDLrRLEZUzftA1zn1kTI2k+Rl1gCeDYi++a7WCZSLoB
1efO1VoWdp1APUnvn2LuwHzRhbLllxKX/Q+0rDg+6L/titr60WWLn3Hgh5rGi/JW
VJFTxHo4wT12lKPMvrYoN44OaQVZ/X6uAyLXQhXcW+yODm9UrFFZqgRie7eU2OH4
159sJEw/AU7dGmhdodorAIk7b3/OCrU2Wd5dEfDCqGcNHr7quzNcc/4jAsEQlXM5
rC5YDmlmTRad2Nnh1SNEhtQbaYyxk9FPwPJRC4luKqmzYyOXvqHRaRh9r5HjtqRc
d1k0RAu5rnJpT6ypCPPU8NBytEORUzJknF3NFkHMXFrmLCG6GNWIvJUcK9AWbDwb
Ac04wTStKSoN863dCZfSG4zm1PXynpI7zpGBpxI8D21F3CxwMg34IJ6iaIg+YDP7
8D0yeaEkIXIZ+CU2jUWp9hkTTO40ZguNDvqvn0IMyBBB2aBTdiQyfuvsqhL+0IZp
q4EQABVpzGIj6mdQ4oLZ/6Idjalu9kBehIjgjYRsI+HqHlkXa8jYz4XVSTS0UgPX
LpP5JVgMU7eDk3jJQ89C0Ey/H9wSagYZk4VE3o06EDM8Z7t82YbwFNWMlIjRkXoI
wNNjXrTRlgfOVE48aIwRgqVVn4li1GrytDgBeqzLDVKye1Q3JaD/Nd24f/YuaaBV
1RRernCwUMUIV/Rnqa6+8Hpj6DGDBDVKoYZ46KMVKuzqNJT49zOToLj0wfVZgz5p
2RcnJ3AIfpjeFY1xWyrHiLQcyGT0dlgMVlZ+EYpfFKiV5O/QIttI66fSBKtx1WdJ
ScDrA4V0FrEkVcOkMxRs+eUl53gEDgDlD4dqchl3FVhUdjQgg4PDeHWDtWhDUgRh
tyt2xTgzIknjIwYT0FuR8hkt/1jR4CLYW6wstCY+yRdDjkRq9fO/jGPpnMSy+SF0
wLGeAEhIAp2GtzOXgkabD5I/um69BLyqOaGO0FRm42/8c4ZARWRQqCjNwrQL009w
MmoUzdKy0SrZ83dCsQULvd0cxKE7QzxMsyZdFTi/X3L8UuNsVoaS9fAUSxlen1M1
KUVWMN7/T3qwg8Vq6PSaIkOx36QPUmA8nwcTosKiJzu1gyPMaPUDRycudahk2xBD
wCGo2E0KBkNqFtLfr5PW4jWMndXv018hE9ewHWkRgMZJU/nieQzzR8ekrodUtkHa
UiaXR84sL+LVz+EHp9XjP/q+XvHIs3Eiy3sv7HSB2QoQohrBEMIniwj0Bhl0wDp8
hxaB0op+QQ13ZfRMXceKDX3ZsDFpM/iWmwMwGA2pFKYANLPL8dkn8ZsTBKRlHbQ5
pbJT/jJWVt7OuNDyjiokOHNOluUE1zrWbASA8KGbCJkwam3TeNZcijOhFVZ+W2W9
yzDvMSLeGtiwFYgIaebpfjH4wgYg8NNe3Ucgc4HbsjQBYSmhcelCmZnHAS2VWXSw
LOmXGcewA5cs9LI6pACDFXHK0/F6n5Nz3T4M7m3d1m4UjOttpp75cvRRiCHp6UVT
vGZ70iqAZIajO2LoChhFNqrGx3W+qo4dy0+bTKxINLsdwyFChqJTiaQlP6TRw/tb
oEMtct87+uTRNX5thocRikHCzFcbwYTA9jPiU8fdSwcACpgitS6LHF7BcN6gzI9S
71gvD2hBr52zpoozqIr+zqQKE2IX0J+pcrvpaR7at8l5tA2VtDSwqrgKg4xlavCv
bELKODLACWnU0tz2F5gdkiB74gFii3g7lGS6P4L/dCO8uCpzdyGJFf+AC80Ycx6e
6bsHkXEDO7vwsPvFKaOeUL1LUUc6vCRYy1L83pHMWlHnyW4cZIyGwBMp4Kqc/lVR
m83hARgwQWOV3S9EIylglpu3lccf5EqOWwWdxOcmNjE3Ww1KNUttcQ2m7DgqztH3
0ENjTlfYeS3ZL5GAqAO3sxiufATS40rpzpDFqPVHDi2QBRDZRaORA78bQ/iiI58O
u+KqUmj/2sJ5WwnOImHxeJ+CdcoHuTYOsZOpen0aSmFdPlws1ZsKLJiRiQr06f9E
EzP/otvbp9OVfdZVUBzjEnHhwvrsLQNGmdJKUcvU8qK3Vv+fqBUvBc3+Yscj+9MB
SjXo4GgS6bLVb+ABJ3vQfu36IFYB1tD/SXZKbBHzDbybYPtBHUZNYxaJN0o7gSru
sJNtoGDUQJ5NNXonJ66fZiquIzVeprXNcJ1F6m1OWduLBadB9F8QfPcm2i1A5P9y
iFRRIByZlI3BCQhLg8fYkGYIUTlEi0PozVmEx9PH5OGc2rMcYbAK/2C6U4OeKXK4
g4sE/wlh0kGmtnPQD4Fwn8ZNjYC6IhNmvumLoZNLsuX1zre4QDn1M1stxOnP8YlC
0VW39f6KNSJw88jWpyQ4JE4RZtTMGYQLu+a0HPBAr3Ug7Gy2x9Op5I4v1E1mf2Gl
nyAhmagV0mPa447XkAGojbf0XyH/t1b5WD5m9z9D161aoddKd7Q4Svt6xIp3POzN
x1PTSV1B0olb8kkTsXMsuqBIRaHg8DNlaTl3HSpvIG2e50Tvip2IujR6oLMlsgTg
XTH+lFLeJ1pb2/c1b6XsV4EbhFZtgGoX3Ik2XDxAnO6Akrw0xI7bSkvqvv1vIYH2
gfITsbSZn4jsBJFk+aPdcdMpIlTYEhna9PpGCYCAu30gJZZej9ClosVoVK/5K51J
S6BXg04zHdV9e2+mTOpt04RDX1el2h8+H+A6YoQ5Dx9C0QFoQS5M7Jh7uPoHhPUh
TfQcszYZMoMFpmekN/tdgo9uXOQUaSD1MWBxj7ZX8jZ6gGBFhqsTaLBrlZKMvYY3
ldEBK6Q76Foc2AoqMzAUVXvmiFMNy9aONR/cXOMLCllig1LYZQ8gynRFd0TttJqF
h9shkDTYsmNh14xU6yIFZRpG9wnPZNIKgRu8tkDuqyz/gcncM9048YNaAs/VoJtF
tmXUKSCiSPHO80yZPIbEa4k2uLDd6gTf+ib0V/Y8M+nMucx6kJ6Eft8cQkpoZn9Z
z4c5wo5BbpEQm/rjJ1mBVvK4oRzzd9NXMI7a0zpw5GbxfVx8auV+JEjYhZk9pvZD
z6UJNU4NdnEIwOjzWp6J0rH3ir6Zv+h2Jededkdklw+bQl340JqeDM5SFuCOE+ab
yYbXqcVdvw8RmFNTMV9sBC/tqVNL2ZmpAZXuirPd89iAIe87YbX6JhnaUdSeVqBE
kz4WySFXdv7kNK+JaoMSgx2icGNb+zCxshHZIaT39lBcZDkZUHwUgarRIY0OcXtO
qohPlKGYtr71TwHefum994IrhHH2R3494kQBCYgy7wTlDME6smG8eCgJeDSp/qnm
0jP/ev1N+KHtuEM+L41p+AFsSASaD64skKxqLgqt5orebOirYCIJdcSPvGrC6VP4
uVeIYJTwuf0QnteNIO91SCtTmW4KR+wQ1I4QZmMuILyerC7AP4V4t+vFSQa+feJz
rKiaopkUltwU++0N2EnoeCNcxAwLEMlqZmDp7P6ohv+NuTyVyFNlAUf3M+7JabEb
IlsrzqLob15Yb+/wPHAlykMKteMxS/NzXM0Ea/JPBkV007s0meujHao1xBLpbqLX
daCzq7tWTAAEG8gJ/zFVlKr9qTpsVyCUGISnhup5alL6Sq6Mog9Gx2Ly8WaaZWRF
2wGuA8IEtllvcK6pd5Gc8ilCnhYsepuCLjy+W52zcN3pHtoTx8IWArbaielEzC0y
90bw/zd8P7HeXwUyDmyUOsP8J5szWO4YlpMm/fGSZb2zoJ/tkkLVo2VFphGefmjP
DT/dyYlmlQBMtdKTkqzSiMwqGfN9M7bUdskZyubwzMbpuJDTyc0LpvA/0PEJYFdp
vYPxAyXAd6DydzqKBY6rzhKy+zFGuajxq9syiAgQTaiO2OMjzjD817rjgr8T6FWq
r/1z2FEjh6dWw6ESVTBhFTTFvFXDo56Ix9iczCjrgXiHtinu43PbUfZXM9oddiqz
grOl5Y9MlUBhmyQTL3kRmzxx6r79Yum5ozB+eztout7AgYbQLqoD3ynZQdQbVRcn
CWximRbGME2lap+y4m5PDUTa7OUx5xudBOqGvb6CD4Q79bP9O/a11/Gu/Fb6Pnrm
rrlLWIm6YSlvH1AFChRAAgISFmDpPtgWYA6/xvpOKSquNI130iRHORND2jMLrz2e
MmvrhY0zBg0RmZGZ627dDjaNXYhEqhz2NoLZGd4aSWUNFmsv0XrcN2vfRlTnRsJS
3nuiZlBGfinPkofmV7T9FgeNL1Nh+kkQMQBbmpQY4ghjNDss3dHn+yNhEt9Hp7Jy
jIf3f8b8x6yKciumIw6is67azyR/e8RhczAzadQzUjm481+lyK1394bIhzT9B8TE
SqofTk2jBX3PaDduU4pnd4D9HElNtccaKWcZKkfYTc829x5Z8Xdu9yzKfqrL1lcD
KdYf4yep03meC3yEVIE128rOAx1ELEAhHN8AS1D/0qj5jLVGOzHIkBkCh6zj3Iyq
iO9UITJ9xiTAmdIA7ypaf8+m5GJOMA4FzG8SVS6N2/2u5Y99pFsEPElXu9YXrbEq
GXlctnpEHZZAE8WwQ2JbhUmGRvrfHt3F9lM09SJ5mcD90DJWVGHgNjRi4j9zdqsh
N1vY1htP8ZDClxFox+n8JcyJYKzDh79QxTfvoBm23cUj3mYtURPINoOxtyZWnC9H
AyhHUgvL/WK+VsAwaRepNTo04iZLnPANp9aqQZEuniRaAbev55kLfroQLZ4w7Kae
e04L1Iw/k4N5EBY3qcVLQar2KAIa6L1rZzzGM8SM9P/7AHeDWIC7GHPmF4D+qlC4
WE4A8NmAf+KqGD0y1WSQej7RommovckKSOyyf/VNJC5JizQIPUh/nDSY5K2NgRb3
SI9uB4vLR1pI5bZiBXV+UG0BWVthbtzL1BTnSIVrHlL0QhGP9sryvJ55lMbGzX0e
Kt+p/DhLW55G4CUIjqeKSiycEilkAjykTcIkfBeCCSb3Lnc4RpiaYz0TmIyWOhiM
7+N5rHylS8bimWC7DuyCSwMVJEps/ztye7ZDP0NiCI9N1GbJLLT0fikCf0hSW0CB
zCE0Ps5mcVZckHBBJcfao1zhPPAKx3LxEiNaJGdJJHPkJyfXMj2DOqVL0HH0MYFD
J04V3N531fPivOAaDwzgsdQGpWCa5kD96HmidS7lxrBhkHxe9Wpgty36dm6dUrKR
1/zqoEjgDZc3mnvF8yfxc1LuZDM245lqHk6R72uaFgyQsIzeEuayLKi7oW3wMaK1
5PIzJ5ggfDvw1d5t7krXNH2s2CXgwCv2c8ii5FkTZAHN7sPHkrgitI6zmbS7f8Vm
nmKefgKIjac+O9I0nDzXTswgFnaYKFcGmlFAPh54Amk8XlLb9uNY/LB29PGwMPx+
jo+Nscpm98nJTSTIPOTdGO4PHa+Bq3puAvFZ4wjcvTzh13vJxipahxZto4Roay8k
UQX7g+h0pLYAKEvutumy0ert0p/SyQX0aOIkjA0k5BDNTUSxgWiSKUq1qkIAPiBY
dhUO6pihJMtGN6ENHK6sqRRrf5+r1BqxQ5Z1OQ+1DZ90Ev63eJavfXgSsdBtJA1c
kKT1tOciJjap+7IQGoNJ1Udl8Hk6MQtZCF/f48/ZwjdsJ1wpbx0DJ25Ebg2febJn
Cdnr1akh2rCJ7Z8Kw1zmK4UskXk/XqhFeH3TE6fAs+Hto3nArH0x0FIgBRBhydsa
k8y4mdJCyEqGKpZVlc9QJBCcchKwrLKC1lTE5x7xzGJC5dCAno8yWZiv86WR1xmS
9XuYssKOnQJrQf6NmTYY4ns40kE9fMk3Txj4o47VWn5GmyqqS3zL3aP++riRgq60
jZdNkhRJ2RraZqOFAEp9/rpW5GlDV6xMrAwaU2HbLxHKGyQ6k2URC9gcnsj1QtL6
eTVhiXghrRHqeaKkghDbruxbERKF0jQm/d9MLX7BSOnSBZyPRh/4oBDo9afYU9bi
Jxtuqd+6d/UeOw15b0eqUNnmoQjJYq0KWu/ZB3Vf2NlbrwGGBCRFsvcQrcXlQb5z
mu7jCvwxyv4h0/EEhB7G6xrq8yKvP35/1gnBCUs5pPimPumxZ+/1nXUXHx9Ggw5T
PFHdPOiIxPfVIOMh+ort2mjOJKe3ovEhfIzE5Za2hH4blVzIRhlLKpAlSUpT8BR8
FMnIHlotG5HLalz9HG/Vm368gQUpqf/CDj2iOW8j6aGXfDwuGcY/zkvStK1OTUts
C8mI/4Vl9ZqpK8bSyV1bs163T8SjicyNNu18KaENp6uahH3PImEeSpjPYqNRH0HO
aAoVaoGNzxFwQke85g36ymfslqVuZVoqpeMdrN9qiLeyvItOz8mssmrILnfxtZwk
L5NlQM67WHQ/SvdWkBl6lOed8Kh1Vsyrc7WwMWdrByfXdby4hhjwQBpYJLVIVCEx
77b8yr0kvMF+T6Eq/JE9gm7rFaU1/Acb8Q+46Xy6hliH4ldCzKMh7DJMC8bambxh
STSveGgLTgILGejaInm3H0Mz+KgE6e5o/Fo8k2Mj26jlu3pnlH1+VHdIuQSWLdjj
8CnN+bezoOnSYdWzM0MkjPic+axhIfLT4yp3Wrws/3+BGz+3vEHMYMzFnobVmO5D
2EcXufKtMdP7+MWF7Mq47x7PvjMM0SxBlHQ/RJSGkCosAfs6S2u0TW6iYGym4RXP
Hpt+B5IJjgnG+/BJM3IkdVMNJfz+a5MQ4mJM9AFLmniiMsWkXF/gxLZCJavh7nUN
5dPhPvLrnNyggbQCYGyq7KAIE5D6lvifo4AiJXaOilTkkyxiVgvPbuUxTnXAmRNK
eHxLbpN5MwJkmfqmxP4L1+PVOAL+I+EgcaTHk0PzjecY3+M1IUfOi9AWJlGFbuy5
jZYkG+ckorqV+fMuWjbmXp3wmObIMqBKgZOcIaJfjnS1Szrx6BXUzD6UC6RVpyv9
I3cBSrNDw03hCAM7p396xqX0CCX3QIPsZx/D2j10jIL78HM6T1ZvUdXrQyGBZp5k
auqYfK1+m6AFjYoxoIugGQ5WqjJrR1nI0xsxKWxn7RWyvEuR4FhzrAGwxDmrLxu1
3YEXkWCPWG41pKTMfwFdVR7w2RdDSNgdY5vOViDRObC9Y7okZmZ5G++NeDhB2Vip
spsR8cgFqJMXrDPCD5YCwTAW6nE2YSdPmQxC6NK/zq6Dw62Q8QdxIKLeqxLpWgdH
nqWtsmkCM8QZtYRqZwdgIOhibWKD0R7StcclrvvFv1yEzicePoC93WtHPgv7Ou5B
RDipil09/Q1Ix4f0T8LpgD4SRTfcOpU0eyYGtiMNJhlzim1xer9PmUx1STfzFvRI
iZSw2YarfDRnq3bbFJNPQrxb8EPVs2Sc6eoxA69EPgLecCeJuOSpDh2qkEuxm++E
TwAV57r9psCIWLpk6/c4t5fng/R4j0H1XT/9qRv7c2poe80edWWNRH5C8sG2MUE2
ipUNQnVQCXyZHLr/BrYnTP0PqM1l+KIYSPimWKqTtNLQB8OnVzCgnvrYn464TgqL
6vFdSs+eHgo/Kx8ZB2VJ8xi+XWDm3dedTMIMs4EgUWXHJZN/qDLfoGM9Ruoc7vN+
25MU06VvhdK2jah/FI1D9ZNfZcQn2cszRY5A0mj5TKYHYFmimC2rzIuuM8CEifTo
RHKxZ1d2BYprD2XW3PtyeN8AWmJjpkk0yFsMRk4hJMAGZZ0tsZoJVZ14U74PpGwp
dFKozNMnJO+pdcFd1TW4QXP4i0bvEEnw9TFTz5yRenji5eAp9x43T/xiK1kRGQbN
PtqPc1oaPUMPEHK1J4Ar/Oy0F1UrrK6SgoXQ0GkTJYhz+SbR6Tcgzw1lSK4LVbM5
JDICuFfRdLwhUIG4kYoZSmC8iP+25jsh3g5wwKM0DA/1B0TlJgjTgSl4MtG/FyHG
r342jfJCeFyY5eExCUUhuCxXU+uPnmXeRTA0OO3zyZfBcbWDN2oz+W3FLZsmtiIi
234LOXRobE6QDsZyLyF8BNdrov6X/G/rvC90lBdXDq7PREy192qaYEpFSedAGNEB
2OPC+gsUVmcCoKgQTAOv1te3YbIzlzXTAONzSRuD3c+0LSj5HFNqkqpg5REdzAyq
YO/vTf2kt/LbBvSzPeXyjO0A29wzbXdgPr9VfSIWCn0Y/TFjRfFMLtoXmg7+RWyM
8i/vlmDVjKP9YosH3thuX+PxRSpstMKMBwgwL1Sqml/HILK6JzjklccGkyM1To4u
1KbKzUhESru4QlJlpxa1J3F3us1P1DEeLVwE0SNPLrXaI3yfSbdKPFYylR/qKdk0
PiUaOfGfIJcGndj8dL5Tx9Fu9bqMRgVoY5qoABsL6JFbDA895TTgZ815QIBc+i/g
4e6Ym4LWG7HoNT/KbRLNcsT+00yKfFjW9zI+Wc4/UCuOqrgxIqqeEqIMJBOQ4eF+
oLlHszDVtbY7TUhDOWMl/7Cmm47qeyaZ8A5fNadnbZghkMabWbl2WTGenbt3G6fv
J/7g9PI7qC7FnF3BG5LUtTL0zhpqqvgaNzcAHAvuLd6udZtvtfoVtB1MRgJ3Grhq
u5O6gHfFKD5tB1Ve3KjXRLjFZtY5IrofX/+T3iRRp2j+7N41J4OZPMmgbvgSBO82
fFV1y/+lGuye61oDiN6xPAmoCCXbzMqMmjWnssK5+h9NCOCimZS/mvQrdp+qh/yp
8TRivqztGKviKVYet9Gtn4UnAl+WsOqDGPJi+mliuaqo3xCpya5bHeU0Zjwiz26F
zrKOPAO4DQB1+0IHXf3gmBGbiXz4ALM2g3FZI8T81/BaqRFp2y8TAzI+dZsHQft5
HznRSPh1LxCG8Umo9GI7cUQ6XtZYtseFhRmLVI9WcALdACTxgy2vdBoW9y999Skn
QnAV6vh4HgNt+wDjPrEjmPITIS2P7q9VSigsMkTyUcn8JgwtKM/ILVJekpiyCNSi
7cSr67v3uSF4gcCOO8QP4Q0AvZM1Mv5GP/QXyh9Wa1E3rbHjkHSh950megu3oUGp
YsbjYORYGpK84Cp8HQxWJOSCAl2SS45gUJ+XlCOg7d5N7aRALHWwEm/U6NIWatQK
WEHgxJm70Xa0O5elFx2esj/EhxCRC4pV4C+e3aWVTIBlGuPeIjlP8JcE/Neoh/+I
ACUZ4sL4M7YMF7nUcjPOSdwf9mRvFWhOdTNc6F0ibsq1LhNP6zS90RHVO8xjfc2s
hz5DQdf6KVnQM6IFQyQCYDTcOAJI7vCoXWykipd03VABF7BD2W20Tioa8MA1mJiz
YHwbTWU955rmLrEtSxcGfc9YAgJUdrUJqjxyFcuJGRvc5PR76a1A8tnqCO1EAJGR
bxUGN1veHZWmR2F8+UvpCQtddYlogbgF4R9YzM+uEmCwgdNV4gpz0qjJZknOgoQm
mCT2SGU7zubeFGBAzfUlS+QOK8xly+QICq7qI0sRUUxEXkNXqCtdzbDkIW4rzrYJ
KsqgWGbU9ZjdIioLGE/d7i8B/6Twa485MxrAHdQOtE9crFxBXMzFWtDJ4xnd7gMW
B6g7YXvdi8LZEHl87y6Y5HOEhVxl9pFLozLmpZCO6L4t/l7yxbaIepaxxSw/QJkb
IzlK5hZZWkdBvAPNwnWy+OjgWRN749Ug9ns6x0UI9iVoqt0zqmByk+FZQaMJG620
ojNKKxAbuYrCopZd5yFJosa6ETsHb52Web+Ynm8RDtEnozn7EDK2Q135vWmfTW5f
lI/MgENzDMYZQUjrLY/UW/Xy4IQDo6THgdn3HbV4e+YGMoJ9FVMteLk0a7XvtfEN
JzLHM1Hitdf9s/1si9McXGp8iw/hi3IZ0R6zgo2UviMP/sSd7Mn94BHJ2APIZukk
qkfdMfiF+aydWbPbycHcsdu3/UnmUIshZGEEolbjhZjlpM+YwAcohklByNvN6My6
4oYKHkpWCQpMM5MaVa6SFyiiAW1/81dALdgKrXgBfFskiVNHSIE7hU/T8pRQXk+w
6TPoKYF11jys2uOINtr3i410b7NOiZXlS17lPENk/guJaLI/03DdbQP677F/MAFt
5w5sPugP8j8lvowxBhWSUiaBdCYH9CocKFFGGugzU+Rup9G8CL34OLMHnjoNtQ45
awonCi/013dihkD9wFUmhQQSE5aq1/LMSbez8Ikzp4wFs1tZWR5LyHNFmUqi2nqd
UFgV703/NCUDOJzC3O/cGu835j14uk0Mgy3CV6IvnuRfr6sLwtfeU2urDPn0m1lZ
BzJwl5Ksregr2aLQCvcu2uA7cwBA9vODzHhijFoZyF+cp8DSOfdhyLHJsa73cVJM
JdUu/Flg9I+qNq9M6bHbT7bGSouIwk37yCBCKR62efoZ9kgPchQhSJbEcOXy2Geu
5w2NcMomvoisDGv+vHKP6ExdLZPvwOmzmRdw4pGznMq/SsS6qk8m1J8on4xqBnOO
nXJS5rYgaU3tgeISTATP8R2nVcktxQzJ+/mC6HSDlpeREzGtemr00C3+az5cpW04
EOSgQWuP8xQTjZf3hsK1K9u2qP9rXV9CPTSkWXSX1jEkv1yQiUXxPboamHaBho0K
Y1g4thB7TPU+4SZ6hKy0C61hm7W1fUTWOdxLK6vOTJB4mar1pNPuWEJFzGJsOZst
Og0E41IQvwRGA/2UMuHGTlSq6ojO2NF7TqdjNptDv4KEvFXqP5T1Am3YgJkX4Snd
fzaJ8sgHZVRFiXe4oMSpCNkH9hUVh0gth9p5B5S/3YEvbkFnDXKlJbQu4QrBkFRj
Fun+OUpNfcap/obPXJBxxnryL51110Av/S6M54Pziix7BcuO+zw6Co2Qfbd1MAvP
yFo9njsuIND9gHDVtSoKWMZxhnAPnnOdx19iCVAsmgnNKXIC8ijPAq6yBIpy67sd
cVJXZQeTnl8NN8RpPp3HhRbxYHG95QkzM4UvxLf+SSajkLtoIw7J+HKSBDiYeCr8
V3uC0aHYBm+LLyMIJ+GJoNh5K0vt63WqWGWVP3MnqOKFADFAU00VgYw1Q6yF+3Lr
flytXALGFY1Mda6sdMMG2waRj710gl/4Kj2MHa5lxNLubb6QazapbRFUfeZ6EIkQ
2wAytieqYOfN2Be90MwmFbprfhaNTcAIWmVDgfJ51Gqf0IqhNYoVxdyXVoeYCEww
A9cJO4lSwUNlDkOuhMBNWyOEjWgNGLR89fQLaLTEmKbWzq049h4sZMbW5WmyKNAM
qeEGko8tIHLo6w72E8PwjzXyC4wfrH10EMrdLZqVOouQhQhpCFmvzIaEMdp/00ml
RMnq9Oy3dfgP0eo3y1REmIjzUplHK9PH2lGcR7tRXASHAEN3RlRJs+q953J1G6Q8
evpiRNroKpyFdU2OyCVWTGHImbk5yDS9ik7BamTsOzj2ZwfBAkzguq/MDILZSoaS
BL/aHEURm8wUjc++nWIdiL9uOUt/LEFfNvPx8HDYTYrK7p4nrewpMSl9lzPuFm9p
qBKriFGVQLOnRAma5BQ3/CQIIwP6ps6TcDbUWNDTbthIdWtFm9r6Ogs9VyHMwjyh
Yi9W+MDf4n3TccbM2FpewImzPaN7E4Mm6GLsINx08uMdb8iPIlU1liO1HLktnZyv
Qx0t5iysBIBDXNckKratgcVIFjqnbVR5P/aevZt2SskcjKPHlIEoEvFgnWXQbzfe
eAqT+Q1mVw34ClY0qN9FvD7tpx7oJEQG3A0HwKqEbTywL8aVel3qGaQMp/7zB+I4
YbK26fNhRNFPpfW4RXBzbW5CZctBikjB6xh8k3wzSvvOBuMwsRN5qEuYvTCQ42IZ
SC1tFFCi8jXb5Fmomg6/qtgVOQ8y9gL2i9YLgz2cCGSFcFpBDDe3kymQRFWkT+Mc
g5gz/OpuGVggqVZJDxsBfuJfiw+KmmAM+nkClmbrSMk4NAMaSXGg302AQ2IKNzIP
cWnypQ/W9Df2I/usI8E12wqu+NTfPxN5W5/JmPpPth8UinT4fy1v1tKquPFNvjOe
XNF32zu2LOLXIigFci+DkG1bUntiH1jh8btkFlntaxEDEJXsFc/MfL4fdmfRwCEL
b7bhqy3llA0JSMqBY33yfkP5VQLdVtLFCyHOs/lduCN3ZLEcARKg+6Q5Zgje3uZn
c5kZoGHPaFyPBfPPtQEOOwhiYksFKsfdls1vdWBQwmG3YJVbAcvfVt+bVFkKLGBt
1v2uvLj8i9Au0tJuIIiDkdY+usWOOW/v8zTvlBGtdp8JbwCN/HuhPOKaIo1qkra0
T0cpI1RGFoP3JosjKPJhCb/8CfNUbP2t7Rb+D3N9tlYxjeUjBspNunMYSgNxQm3E
8ap857rDtQ2KPXMwd4cAMQLM8KpYl0PtRzFyfcK3soy2FVFb++p4U4XCqwVun0n8
MHXkb+uBZU9n1ucxuODYzRlFSuQLy36b5jEo89qfm2s08wJmvoNE3jmIOGUqxszA
KUTy54JhgXBrMnmRSp0bQHl88eUVZKmVuLN+DLzjuad0k4+zFpvLbk2nYs8apZSg
K7uFpJVO7SSH0Xfg4Xsd+JDoqC+X+buydJF+H52+hTlL4uOQJppZwaBrfAv9dkWP
V2bPKKJnDA+iMMuoupvNnfQJxcyt8pZ0A1Ez5x45pwTYwDdrdWAxEBqpFOvaU2C9
DFicpgrTFQpi8HY7hdz2BOdrsOaI8Sv8FAl3HZCBSZYoHdG9f5Od3zz015SQ5xH2
i9qAodyOap6z6usppja9PYcRUThuQb8gjDj8Qi2BlNiSF3eh5bqYZ++i+bsazTeZ
ljmexil3ggxZTpEhS8cZz9mmswxBnAtzTp86CbRuuJFN4fn6lvrvrz310YpF0r2T
d8xloTJwFlYrH3Iu+C1qtwGU1wcM6u33ipNNZ3KY21wxlBUSLeikNfAw+WPo/1Nz
BL/XJcDdBFVeVPBXPHtLRShBrBXmUeX69YU1ugcFwhAZF/5lg27OX87lVqmXUFVK
NlZSbqtR6ygRw1JXYOIw8G+Mdn6wOZqawtSMtoP/q7bLLwt7CYOvKKuPni6CqnEM
tgMDBAk1tVdzWj52S/q1kMP6suM5jtbKbcQzH2e3X+6ZTjAwyMcdPiOpoPW9KfyA
Nv0mCQ13kDz21wTb4rGlqNlmvOXb0pswC7W1apzwOEvq7ryQ8Lyx8Wd9MF4bNWPW
tFiHD078hKrFfVHxU5p8mA2eGPHl5Z5zNtHOaCcza4BNVk20BVDtrQrsRG8CPBHw
8+nt5xIa+WtTDCIZpL06UNLJY/IgPz19bTpsCgWlboFEF7ahjRgd+K8LNHBl3q6T
qfTNtmqnF0YzWqm4EYYSPL8gD0FYAXFYneUuhyQvqiVf8EpXaO0RrS4cDV70PoBq
Yo0M6TbXgTu79mKewveeP0ZaLz7oPFayKQA9v2lSNIF65EGv+Om6RydWKBgXxnv9
NuOU7z4p9XzlXQGlj4oiGNH37ZSIfUeEmHAZGmJvK4vZhOdvHmezEodvayrptghq
pBjoI20FXgjthCJepmHKa7795Z2xBb1BnRwWCRvakkdzDreX0uFsJw6eoflbj+m+
VD4Cf0FA6xLjdcE0wxocdvP9bC6LfPSRJ3S0Z02+zd6bB9T0r0LNiABkzeHETScw
xtpNBl7AJG1eyS/Xivx/qxZONaGnTxF2xqqPvpraS9YVwGG2Zv8GOqf/jB1tOi9M
XYGjiydFtf/3O5VByq+xnipjK6lhKvcu74UyiIhAfpR6uMa67x7HnxSDTeyTmfhD
UVT1Yk7AFLJ5O6XAxNokCB06PM/c9MN6IsD/uDVcmfeymYnXiIVfE7mxl3R8siKN
Uj9kPM3oGjSSdAlZRTrHuJvTPuss7q4tzQZA6l+QvR/hst2YHZyKmDW0whbSmXvG
xlbWqe6FFaeSQqQj16zOwuUy73jlujIdIdqo77dIqbz5fb6/ahHx/66dt7FViQY/
0yJxSrzzwQ3VdGfhW1AudmV9se6KNJ5D5w3XJdaQGnXXhh3YgBd/qWWDykfp2uWw
KXuVfSWfO+ZGsZfYgAd6DSQ8yKtKk/sDnnNaVJczsWSz5BCf7c38iEZcpVoPQDEi
O4JRvoCaluyBfqnFt6KnliEDYIlfMU+tKKUlfmEwNvS7jj7HamQG7rsdCVCdezyy
iQBX7qXEw7aY5MvIkpMnDubvjZJdcWuXOXFSLjMUuK8m8XJazqNIEbIINte6PlnS
Mseb9naZkw+wp5UDanI509v2K7p022ubfrkQM/FP0GDPnjSvwaERTgmgGFufS6vP
JQSWz4+sljoQ2gEzW/XRDk0U6z5iJGP8YolY5CwcIxErK5xjx9xSjKg5BFSWyA+u
xnyWTqv7/GDGOYva5SiF0ukYFgEdQAmF75WEqvQ4315ydPKHH6hjU3yjXI0a9bUH
I+D1be/LrIqAVscziOhGUsEdAqobi8viGoQR5pX2PE5eV6lWRzcRxEqHkjRsN2dy
FeAmlIA91/uf3wUZsOEOA3kkd1P3TLxCUhwK76aFUIdjgYivCdHqFsV361NFQPX1
hPQnhkdcXy0DGZ875t6fUUS+n/cZVMRivuO8bA07CxVM14XF9ec24AQpKLwQhK++
9a9xFvkzVBwxNsAzWQeeJK7ftL4rNBRLOoKPRzl3loFviGYfKT0/3nLjI1i9vFD2
fAps6xMqmdk8kkaoG6B/O4SWrocJOmiC3zC1rejtu8zvdigaW3Pv5dzq/G7cS4rp
xmKVsUjH0yfEFs0Am2wewS0e7qKrFhWDhEooeqTyMBh4v5npIkBgN9cjwbmycnYA
wrEqd/hMgg3kaF7YtZB2fCO1Po5JYNzomA9Z2hz5+thGu47dDbZaW8Siy6OP3etB
JBFZYrzsPb4ubFgHvLOzhKRPZLlgkqcuPfRVDO9COYJeewGRDMhHRXCJjRjsby3x
WdKZ+iB51TBOWJypc6P3XiH2rxN5p8DqBy03Xh9BnHve3xR18nHhH1Fytxc1zAMg
GZ7Ivl/9ZfT3AZSv/s+AciIl0RHcpBNnX/9NY8bdJxb07vfzIsTb/Gqe1NaKJ04M
g8Y9Z0HiS2FNivcE71oLd0c5I4qKLxGPCyy9iRQGg4SpVIsGxzRghDlS02xq+fvP
o5+5qvMHsu/+M0znzLxcnyScnOgXzbcc6eZEmxxRaULUkxGGo5cI+ojBz+ec1dXE
UaKrIQu7Arpy8xYazNTsS3MtoHRGla7yx8Gxk4LSnuI6qlfCsLBZNBGo9M3ZAyoe
US3edhxqBLPToGQIcwLGvIquv62YZ9RvSx8QtXlnvMlKKi5oRFjKVmlcqAJae8Hw
ury+9yiFm6n834twXqZBkuBifzyFsG/J+rTBYC5nC/U97fHVO9G6+lR6KLImjqgf
aTYmgZa1gu+EHLBhNBOgpUMOfIfSK50QhM3PPw4rCArQLL7DAxKeh5R9DIMaftZ7
HN+rNAsDCHRcEzX7jVcTTzvWVrVRVtmVtkPsScojF0T321VMdVpA2D3D+L6nOhkg
8u8GMEQEJaMYOE4i5EHQoqV2ZY+HR723XxIVrFo1HLNLHEruLtI9QiZpYQORnveE
2SDKANwUIj6Dm2eTBELM6fNtTML98YcCsEuBUIywYWlZBEW2eVbiJZj6hIWhu/1P
OSDtiBp/yq3MeTRSyfkIRVkqWpAAvLZc4HxZ+AdKk3Be4ivPegSTG2QVfgZyA7E+
EFfy7NscDBU1wjhvd7PaST4+by+VAulFAbnQsi7aUQywZJAMOFfmQS4mhdeqvsLa
NVVc05OFgfKIhgjCvHAbWevdztZ80O3VVkRuoS1RFbfVWjjiJKcvvqfGXsa2p4rC
ItM53he8cpWQqVRvCzcMRjBRTNKeQt0WT/5pJyEB9Q2xB9f+bVzhm/NYZcfmfp0i
J9d+cZTgN33Lc+LIRClIbUCqooA6q0TsbJzaB0OfIXYm/gR/u/QpW2fKruxkyKjx
e3zU9VyAtd1d5bWqFunJg7P9hXf1leMC9lUsIuRHa/qAb+duC9SvlVbkzTdPC+gc
ISOFHhHCZ31OqXKzSU7lMxxOt/Twp/Kd2wb1HQXEpv3i7rUv0b0g2ftmL7ZdTUt8
/Ynne0jcn6U5t6M2MpWXqQD1b+JDKqGTJ9hQcCRIdfcdzFAITTQKf1Na+PGcm89C
UaXsSD+o8bc/u1lUfBjoex1Emifzij/VsY1uR2lnIGaZIVVUAS4+YodZhDdRX7FH
a2DAysD37yfZxSjpLkt7ZQtYC2xdca73XdBsMwVAuLMbl1Ogb8XP+hsFzH3e10QR
dgKP3Te/pa8fep9nszZUAvuT8js+Sz43MI/bPwrM3ZQnk4njOINBNbi0S2rXt/Z2
6X8dq0sn/mQGloZt6+plT1sj28LF857eV+aWufCqpKZD/Q86st3xUzrGYOK6w67/
9jQW7I0mtSuYjq+1PJXBiSWfFHVy6oed3VskV8FY8hkJ5Ic3YAwHvhAf59dC7vPq
SnGHS296q2boEBYqMvtak7IedbBppMNBBTqI9+EdUIZAzkuiv4LxzvNZXV0heH7Z
EcsW/ssDLkSjWjir2vsx+kJZl7Vkgypd41EGixLrQN9yK1Pjr68km73GvSADJYRV
dh64g8CXkstsk+ifDK0LqNiyXYtrcIb3H9itxz34jRfp6CUQ+anc3/ths1O55TLu
au83j7UAI62jdAo11O5QhkHTK7TDrzzeCNfHiEBvr2Hw7qj2/mI/bX+H2QoMEzRf
m7btApVRgpcPOh93xpBlg+hgXo3zoaPRKMMCNZsbKU53Gmoa5HtzixXxad59uGdV
pQ3rFm0wBCgPBAGl8AgAxW7AkX4Qf6M1psUWG9+R+6SnMAKFemzUjz4JAgQzA7Zk
Aho+lshAI4IGVJOhlUQ5ljQrx1ENgWKBSe4MKtEQXgiv1TJqcEGVuZK0cwxUoY47
UqpycyQ54rZ/YV+wogPOQlgZg4o9N1I8Xp6NXq13rKztH69jv9W3A4C4VKAPQ79Z
DAYUjV6qqfEytFOuqQV87+YGwCC+er0XiIDk0Mwt9Ezy4+9yH6448AYoNwDz/2QZ
O9qLVTjwfNEDvJNazgD0x8VXPzceyLp2yJuJhFqAkmNoa5WgT+E2smta5sSttAeu
jC+10Go7uMw7BcLKdyPbQreC+LShzYhc1gE8RKjoz4+SEKjZf3iOc4LMBjK8/yJz
2D6chZgRWbIy1n2sqd5r57uhn2cyGUrN7ZZuSwdcKlgBeVluLPxIbbXXlNirWVZQ
HyXDYeBLNKp2cBI4Z5gYXc4e9/hex5kbpTU1vcUB5AAe5P6c76VEOdbCLLBPG9t/
mVZz9LGfRY9QESq+1RRcDN5mk5LmRSFde4TZokvGntfIF6p7K0thDwXtT45jN1xY
PPYKpztiCBww5vKQnnqKmw2DHUf065uvr0i4nDpg1kI5eeYQT17ZFBJ4BIQwR2+I
HDy1RVyh73C3Be6+lL8dT4etc6XXJeneWPKvY6hyV57Tt2NfLWFUVwwQ2lsCltG+
fXPhEfoABfJ/nEpoc/LmcqJO3hVhWkcMWtWUfGDGl4WONMm7frLmc9iBLfQpoyvA
R7/YAU79IxQaEchupAb0B3xs5Bz7HbkqGUz1mn1rdBgb6cKcSIDDbuWCBf/8Ixvp
bmBlBDQHJz9QP5vsmS6gYe7C1ZZlf604+NySAaht05GS2G8/ABF8erOLR7ElcPaN
d469i6IkJF11EPcJk8KzsA9MhklZtjQ3aqGdZ6bYAY8Pe55cp8pDZpDsVSlR391J
VKcR0BhK4gidCHv4Y23oPox9uc0sk7KLogrfzVcavsXdN2DgPl4CyJl18HrYWrfq
3P8TOpQhLywOPyMEw77vhcI1KfOK6IP+BvUsFU63ahIQenbbOtZ0bgGets//kesw
1psLaOU6L75Zf9C2R7ABIe73FsT9nUQIAOH04B2SA32qhxHnYTqH+uuAzZ1W/CSk
S8DRkuG7gKo5EhzDViuiBQewIut/sWE9Gwub7tmRX2ECBAnrnFV0IffY812ZoW5p
9bRPt0zlWzMxb+V8x8o53L2g/fpORgN1EtjRYfQLcRisqfSPO+Usvn8kf5byScs0
O4dNKCctS7wYoW5Aufo6VAOJSQtFTTbcZEjQiVzE/gwdQG0R9jyLKFA4HAHxdahz
W43uxewMYb3HP7wiemUqNJsaoQ8ROt6IX5NEFTBCFOfOV3ZA+eHTmKDvaJZw0N2Q
wadGaeytTLDjVcwoayCi5YNf+QqWQihnHY/WBXWLEZwfZHejf4DLnoueDTAS/YSS
fvJPgTqvEkKVI2swiMZyo16G7reK0rGk2ECMCapsejzuDchy5r5+8K4Sxpr8YA2J
Ia8IwnjQE9EOdGMbl1eYOw5ud2U60fc7FCkcfnknVEvE2k5w1G2ImXGO4+nYxK1V
Eg7U6BQBc/OSJ3u8BQPEPdFZgm79WH8w7qtWVA2WrUeRSsYBnrGZvudFCI3ZC6HR
GnWqLmtZs7Cq1S5VTbosnGL+R2y1HwURLnSwUBT8iHweKjQnVJYQ2K5lzaAYCWDi
oDzk72pOIeiGes1NRC7YWJrZ7bzg2jkLzEBvqjQrEJemnb5B6RLgyu/d5NaakfDx
znAeo9rvscR5KtXGKUogUR1B2HTbDgo+zTp+9ni4iHvnMDnmopD42zMK1Nbc7mXR
Cj00CVXjNkebFSQwtB0g/FIEqP++f02YsWYtPofpcjrqBJXbC7CFy/2SDVTS2Hc+
z4twdee03jtQJXUuGCF1fCptWUjIqohF88TmgP+opTbqqTp4a7fuqtPXNtlLVRU/
p1+s/SgQcR8Vy9ocDdefktWl2k/L9m/5iWjfISfbhoNXDdhbm7Fb/CVv6VaIJ+1a
TpvglHc3zGhjmB6uoLC1v+jd5m1PkthD3AcFD93N550FASQvbYbO1VcVJaTwao1k
Ni0x1lscKdrwTqwfapp39NzW9n/D9DDQsf4ZuvVpy65Q4sbCr6u7T5feJjaJvSvm
5zgS9MCul5uPlSRMgPRP/DuJDnH6XuBkw1+OM0L1+KGWSTT9SVVo2A/NfHe0bPWQ
COeH6Fc+tDc6Kg8LOGb/JOATNHlqGa9B0mVWiUQE0WSTuY6CxYPpu/qm99DQbXVG
TrqNqCVTqe+rgv9/VOiYo0uMwKHkwd+zqVPGeo8cWRViEUDfSTWgLOfxU8p5u09q
+22LgbnGXiuWhZhuqzcLMripvIBAuU4/keVn+JM4JLk71vksAWXpMkoHoOtH74gb
MY1MGMU9EusnPAz0CvZJmW3otsn+0CxQAqzG9GkpmsRngo+ZVJO9dTr63lDR7Atp
AG+7KGIVqgVHN9y9lqja6ezWzFeR2xqz6lAOFDfph8wKsZYyGiWhOyvz/WNLUH/2
KwWNrgoLWmzoG1IMw5LARleevjVPE9V9JV3i2GukROYALZzbIyPSFx7GZ6C4J5dQ
nalxSu/OouLJSgbewLfjVJgzWJoSEs7lloJ/t8QJvqvMEoq2tiWmMOpjRvpbf0zs
XNFFOQVh/qgLZr7BibBehErjw7cnEBJUZ8RoHTFhOKzOKGc2mvwsh9btzsRTKanV
fWzPuCpU5q04ddLNXo63PeqfbnmOSr8oRz2lPgyZi/wkk8DUfyC2KyGD0abjxNfv
jrota5uDzsdhTZ4AZMllm/stt2mJoCAbozi7TtJYx7F77D//uBwD85dSIv/y6y0l
rsox4R5K84lYSc59iSegIlOhZbiM0Kbm2/2FPADVIqmq6/IYZbKjPUUzV7wtamSS
DLm2HEYAq0stXo76HYdsdJowZT8ehbzuaZqitgzAQH0VeWZLyQvroXptpYGwGDDl
EW+QhdDzhjdVaPaFlf61mCUX+7tlT+1H3Lc6eI57/OAwGsHRyNJUh9JebRTKykL1
KbjRSsqyvvurV9e7S/JIgk0bYi3pjT47DzqC2XIgFouqArfk4TDlvrXSdfbqUNPB
MZFNPVkJERXy+Xnkl1Gjs4fRbVkAcfVeT5oNL0U4Xnr9nMbaqPrBCTmwPM/RF9j7
PmDa/PdYDOACevXc+by5deGirod1a9CZQvojU3vzLw1HgvyqaPGfXJN/tOtNvM3O
uBgA4Hqmq4G/XC3/NN873TRC0hD3k2TQtjLuErv8xUjgew5UZvRc/zrwjIycgZ/L
yQM4njFMctVQrGA359FBJzqWYzn2UZPiXi3918EK9w2qX6yN3ikQ0IkLfieWz2ZQ
Y9G2uMdC1KeZ6sRcZt4PJpiQHhhOmkwRS/0iUpePD+Vcs0j71ysrtP8Z4q3oOqB4
qVUVRRbK74g620dbTVoKut2QAeyG/A/9yPy0PHEjhYk2xtdv02eulDwp6uveeaIe
KilD0LkCOKMgOMGfACtezW5orSGk5njYh/a0Qpm008VtuqF/Um7udt2Ta5bRz3MK
fMkbEB0Km17wpuOoe5reBuVPZMYJTEVL3XTWc6MSWl0dzsaFU18Z8+lVlcHnuYDj
zofMSXHhk9jUpAnh9ZirkQ5E4juaKHzTufKMoiLdrU3Hz6lvgFrjOS2eIVlaO33j
MkoDITGOac3NO9ea/2FlKpH7NYBA5UPNtLstvThyCMMngA65ErlYm6OtDb5qrbyY
8LYCWx1tgKCcyTbBN2gD8l/od435MRhBk+JMa8wf78eWkzyPMFIEIqR3UPis9GFo
YpxMmnalzVf4DVJ784CcMWv40NNDE3JJvQ0LOuhcDFOw0reGVcGz19kw16zaSd+p
TLYXSZ8bpfbDTlLAneGR2mYJWRgolCek3YtriPXSw0wEubX7Ux1nbps3yaLHTtGc
v5M1PluZgVYxhYxhfrwkNd/t4pUaFMO3SoWhZq7fX7vzPCuuTMZFgAY4IGZLjJsa
h/wPFNAvBVywIgDkkE6m6CdKlYXaEUrvhI/Gp/VzfPwEA7qiFPdF+2jRY/b6scch
I4bAecL8kdyFHGV0uvfvFvhIJXvWmKv9PbQDN1hCNiaHYo65nHrVTrYPObvibjtl
Rb7aBND1hZjOd2lrIl9VHCZx0wFlIo9IS++qv1xR4ri323VP4GtMv6XLU2AcCU7w
pEfHna24ByhRr4VloWXD2ALcUPm3HtTiWu9A2V8TaeGM8jYkO4usAMrNPEqP62lG
KQU4Jy6A4RFjyAE9Qj0gR55qlKLgiUTD/RLIkM9HAKcAFLHyhPj/CokkciJN2buk
lyco0gcCK+tICnlz/1gPKCPgHc/dhkkKChkZkzwbuBQL57ZsaUnqRR6xdSnllc1G
4ZGZR1e7W51YRTgFrPy+G9dekE1apJsfvoBLgX3SykhLSry3YW9kdC1H2tuVMil7
9C1nVsjHeYxvlMyzmLW6kC/tnZDdjicbiHSlqFErZpffgQ75U1FCNL17aMClF7cE
oseB6oz3anKi739uCEpXD2oXELIkUn8Z2k2nj4bJquGyIErojWpjXfhkOtXR1mYM
lPP741A5YAj8dYyTrCTr27G65acAAvPTSHiD6xxU7y4oe4T8ib99v+oNie7ZHscq
/FPxCibTALa/2B43EKsa/IOt45d0cBuG+H3VTf5PZg+b2DoKs6e9zMCX8P3t90/D
NLJRwrGzCXD76LOK9NCG9HHbAYghFseY3HyDcGqFIxgXPgiqB0SMTZoLiD++Ror6
0l9cB6lNO48US6qnvOw79fPh4Eo+pdKuR08nigS44c9s3zfuvKjIxyx1TRjKoDE0
r0723XHq8G34z5tbi29i6Hfc0Hr7eRz6Uk4Qs2bnZv5fqpbn4/Fa+d9f9VcpMUEB
RJBXGjBiBcRO3zBdDJLHNBOdOy7KnXZW9GmveQKiXs79DzA1ceVftLJOvetO7bGi
XCDet24Bv/XJmzL/ytnxhlc4AEHy5tixu9T8YnrGFdZ8F3FBsu8nfugEZNYRWXL/
OAvx9peu3DFgpkZGuswsQP5hnAvuhc/O78N0qP4B7GDhPkRw8fz5l6PKWS7LFlyw
xOviZcob6sWmm2nQG02yqd0gC2ugs0z8uH3kqVaZH3QayDXTDOQ0e9sP9Znqeano
re6kqIK3qaqRbjS+9onkMyF5u74lAn6fplHBPUiXKk2Kb3VIFngzbZTkVKdc6/cS
zYF8polsKIvJFRaytB48f2ct5G/pB4dcxzJlla5UH4u+0M60n8PhdLPGyoEGKWW7
TIAJgIVZpglkdBeF1xvjzQFUZkesc/ylDObU9pc1wqJslKhpH7A1Y/edMDv1aWy5
V8YEI4EJ3daplNd3FrxQ8DtZrwBhVOPm5Xi/Quvf9nf0YrwVMqFlQ2S3f7pHU4vF
ecMBlXpUNBNMV+aE/fg5DCT+cv0OFmMdkKCeNdAZf43x/CgoNavT/TDgXsGE0LXt
uF0j3d2gdpw5ZfjPQKnWiPX0K6HRcbxEYj31qyiBmFYZIbHkVjT/MU/KCcMRrhHY
8sM3mMTG9Z+mJSdX+Bq3sInxFcDQnV8Hz2m1QXUse50Pe68VBLA1oi41/afASRAb
5jMluURtWrEgfH2Ee+3VVBbHlX1q9TA9Yma84mvL3X920ZTdoNodufkhOIaWFgMB
3SkFkyFfLuzPLvZHdCu5oIw59hm2MrlM4lZzNEUlgIZafvJFuuQGYj9zRxbkue5F
oPQaxeEkV60vx/OiYL3FoyYR/u/6vEV7fk9Z0gQgfd9LX7B4u9N+fOjUG6yH3SkR
ppRp1pSeQRDfnMJJ1ksbwgol0I2O2HS2ORaUIVzk704XgczhqiwFK/stiF+6lHp/
2CboYeYB43FUcy2fc4Zyy1CLCWHqm8gCJdV6kZOh3FDexLi6cFAoTBXRn/wXig2Z
xxgW5YSNJVQrpqguF48Yprq0rtPbhZBieTgsUyOWxzlElPIw9XYOwcQL1h1MYTfG
lzlbu8nCcdum2kCP/RmlozLmJerWiiTqHk2lL9wdN9S5rMwU5kedq+uqNhyXnQHJ
werU6AwwgsMo6xLe3Mk5/BLAcUQKc5T7AnNhqFtNP935rXwHNfWY/liK1d9ZOdHK
OmO+np2KHfs/ZT4pnrwIw5rWIKI3rVFG1xpG21mvG5i5FOyeLrr9wb/Xt/dQjzEk
gIp/+c17bC37S8fSoaEYQlOyEHrpsf+WWr0D8Gr9uz2kRzNP1emHAFkhwJt2l7Ew
WcE2oEYsvqf/vXd5A93pMkrPJQCpLYpV1ThwaxQXp6hDd1KcjlQMsEuHEo7LhRGT
qfrw79A0wGFt3nVhR3ISOxg4KWG+v/+YKKNp9FOR4+jkupSYTopH7W1NjybSo1oy
EXYXJmMMI4aRQhVw+NRGK+69q50jOCsrmXz6bzMOfqyfM+tv+ua8VvBEsD4iaxlQ
M/HGrRPW5cZIAuIkuKZI4GupDpR1Bod8zPLbG+pAS26IYtb0ThXf9e5IN+drFjo2
SoFdTw1pPTEXpt+jtJHXv5EI8HhBhUhBSCHQxIOhNvM7dg6txozsAPLFaVoIrAzP
+0px2np9UiLWw1AigZ36pG+gEazHvnnaCbrMMMnJcNmknmp/q9m9TffWgBth+C+J
dVFJ0yNN/XKcmk2rqQYWk/Gedh3523zmtcX+6GX0N/x5H4fAXItg608N4QwFgTDF
G7SHKB1KoReLM6UFT71hi+7jSBynCDiMTBw2wgn4he9tGctDXo2Y708+9u7andga
CfpGshpm3oPuFCNj4f1tLOKYRLUe9Rhk3xLkKeHSoLq03S5V+53A6YOA+EpdzqiC
2fX5h2HIvU0ztX2VI02bLOL9CqtZ+XK3fIiJOkNHRbWCfVTcwejJPeTKKhbFdXSm
TkefZ3RbJni9EwM/NQ5knrRKK1zgd5qDcyWFstIQOz+QMx6TdwVgNu2B+3nR7tnh
/Ad7WJ/7I2PsyXwYCDP+R4hfcCZGtHJqZdiku6ruhhq8hF4xQjas/RYiqdJlVBHx
bc3l8HceJXqySmrkNq693f3xmngUEfo/b9GX/BWSxny2h/L3LH76UP01qtHUS9TS
d/Kf961vfaQu5oPFUV6S0fPy42iqXO9W7x658Jh8XDICDjRWEyPZVruF5j519RCr
zDTl4lvuzySPgI+c04HMr0Qxo96PCY3YPC6v+J6W8AioZpWHAySavFZL6Fqmk9+a
QWvSAAXBEGJVLQTGl7pMinA1CF5Ww4EpsNHR5mTrTdMJo7/AzMF3NNROpuDKX5en
onYmDZcTZDDXZF6s4iNU2/NsjQ57ZR9BfQ3DI3Kci00/COXwW4/aZINYjljAGzKf
SN1fqWofkTQ7ivqUrxFGc1oZNrHR5xmEcL/ndI2mJaz9qganu4L3akn7SSCqVOn9
Z3FjGFRM3yVlbr0I7Q+ztEkb/UfinTrlmmIRJhhRFN/iQdAlcWHobDLR8whcu3Cy
7O3HHrtwmnViocu2ogK+dMwYsxCMOLmnKGH2KpjR4qni+a/amKaDy5VCOve0J6T7
iFc2cdcJgRD92/rcr1lV552kkTcsBWIRZ4a5w6048rGK3bjZ0BovIcRMxpM2Pn2j
C3ORTtnUOXMnD3610CB3VzyRlJDkgDrVzEQX1IFIJMfNfCIYrI6uOzbZJ9qistO4
gVE1eu/HPy2rYdf19Sxhkp9zpR32XjcnOPGiGr05ajL8cWXfcOnBWwG9p4N0nvfJ
VEqVKSF2BbKz88inbQlw/ocwMQTXc4zdqBtG7mQHhOo6HFyv3IIDVoKdUY1c/E39
OsncCltmr9nwOgdKniul2g9wVR/cdJItgS9amRNQgPCtd+92NYhDnZCZqRCAc+ns
RLC6dF7UEjolh4JZDWTXPJdF65ftjVI03+w1d18lT95EVn7aQmEV+6pTmzoEF8Q6
yMGMaeoUZkX5lnAV9nPPk9I/2Xbsnplt2PWlcgTjJWCcjOjMBm2cZ6kexX2OvwKH
c4sWn7Er2D89RDzYwS5a2M9M/Zkffb6gt7dT4PKmfwvocQS25omtsWiojRKbRx0s
cqSIQJ8GsaGsfm09EaRUq9nYYqDm7A92Pxih+pP4YP6sOqoVpStmJPGczPHPK4O3
q8Th3zktP1G1vFsXFnHQByP3BbzV63Paof463aBDPUpqBPoQagHZp2irDJnr+yyL
UuHD2md3FaVJazJzAE9ZCv6TTjUour43ORS+gm7o/LXvWxA5Q6zhHddTGs+zrkTt
nCUV6jILIl3/Zl09cULnhMduUhp1+C+MVWWev/40SXjWNohOAdwETLRxF74HVmdp
ClYTGnCCPJckI1+IaZ5XbIe7/NEXVsL2psGFr3A8z+wYBLpORiZM8+aAuU2/XniI
yUSgXprwjpdHiO2Kyy93mSoUAyNnCHhcvGRGA7TG5M+CCPkgQhDCaY9/Dza/iOU8
YyPTXWALXu+114d8afb+3zsnXwJVF9LEC4g9RibP0sIuuZuTTbXTpTVduGZ91DxT
R0M4XVSugBSE1V0FdyMVBjCNye9+ZM5vXfKcjnjm3aDupxM5oaBb+QFwcxRUEebP
tJvX5gx/TJK+A794YufvSS62MSQ5OlApCq4SZPSZn8NxdxUhQaR91OVcdnozPm8p
xKElRxITpPuvnn52okayix2aG5XOKO+KwFXLDmd15e3wux+7GzZJxlmirGar2F2s
T9wTWa1eikkV1g7zyVzrrYMdXFh4RiHMLY1LMaeolijwuGn/hKC8LeoobL8JtJFE
eijgAsFLudml14h88rGxRNTVyDtdC4/AMHiAgdcGkt334W9mWdgHXdU3Y4w0LHQ5
UJNueFK0JXcr+Td+e+WHVtxY+xLr0eSF+Cnq+HKkDhHHbdnloDDaYbZLiLprFmXu
ZZRDQZ3ptX4rTMxFh72SM2qFy/XQhZKCS6CVrOt8MuDOLPuaw4+tiBFDOEte3Pn3
//cpKlW40uaCV5fTIgJP6SN4T86NM5sjrBfzA53vvGo7sGDhi9oJFdf2lvKfZD9C
qdIgunta1jLqRW6/71jjk5QIrO34iJbwREpBnOn5sHzGtlGWIjFOOxbGhsEG4j5h
UMcQaGaRNvruG85MTNR8b4NpoDytHgij/LJYJbKrSlEAOvA4uiyYfRvuE3Xj2Olz
X0EzfM50d3rpNsHF57GcMSZsA0Jn5BaqmFZFJ8bvP6wF2IQxdaMu/H1gVJzhBz1I
HTe1egccxkT3Ta4MJWoOBHgYl5ZiZQrid84qOlwVdYkl4d8WCH/4++T1pzQ0eRty
V/EzvEVpQxcD07DSZYpx7gFMAzV1P/O2SII8Fi44Y3nUzd5PD5qDGukzb3nSQyC6
Nfp3zDXfGP+sWSTBeypOWRKTbSpteN8rqSz3IfLvs4qRbqRA5FxMA0klOBqqHzOP
YEYAIH8A+F3WAf0oHX2v7otpeMnX+VRn3AIVO+vkvSgT5STJUXORMumc2fT+Yhmo
18ZOgogmHtyyYkLqBLu+otJ7TukDZ8s7QoRCWuayA/lcLzQGqzjw7Fo/Pg8jxByK
mGxxUGexUPTGaepNIUlJOWJP0xVdj76NdE596CZwkU3LKRDUdycDDn6ad0TbBD3+
O1kT4+TNdBP2dEHPC2FJ1D0uCHO5/qcrEwK2v9qBp4TAGg/BjQS/ZAU5uDjzkKZ9
YC7msa8LzWHqeksaIwVqbLXEzkbEvoJsN9C4hdDtcyacyfu9jr9Y5+h09RcltOoP
ac+Y414XTR4zzpIpopKyGHc84FqNKGo6c2eViq483xtIWNfy5tcE/xoePVo9k9Ca
MllYzeNm8/+BSpaGN2a5cf5xzfcSLjyHwgUvQy/1k9DQ9erGFTws+XD2B/mKN7JJ
v3LRb0bPdpiaxKepILx3Lm4C0F/+uuCcztwF+wpHjQmgddSmfuvDVy9x/ajxHS1z
Sr9mwwn0tYiHrvVrd75pZRteZ1ZTpmW2lvsHUQafhgNUaZmWx35JXUud+yPQiSNg
9qIhHRDWhtXYLXnvWFhRCmTa0kzMEWsNCwwqo6rjwSaHSbKjiQT+JoPFWrlehej+
1WABL/2T3HbFmSNqkYMoCOt5qO9UVSZCJdIfgPMauNEA3E4fsk4jAlfnQRZjJCfu
Lk0wqQyI7OgrUHHgqGY16pBbx3bqKzOMwsk54PLmhMvBFHotMP0BmukuDpsHtd3w
ZRIKVEtYE15/zJfHYPAnSOhEA4ah65PfMxaTzGQRKye4OVtwsF8KjB2NvGQyEaqb
il05bSaXX7Rf2IisI+j3mcVJXCbP9nf1DjQ8mIvdIej+IBqs2LX54febPf1aBazv
DlG8mJebFvXgz1E6BqCzFJ6XN7fpDUVf0oGrdlfyPB2FMmZxxwR/DW9S5VBzaVLZ
/d2Sboft/Sb5r0MNOmAMCZa3oIXM8SZCP2+ywAb+C/ZwFx3Z4NI7xoQgYCNSFJoL
zENJTcKt2r2/OcozTztx1P0Y7brLepnidLl7Vih9UKq5LgsptRfcmWn/a+nLeFYi
GTnX22ClNJ9DKSYCxtBHLx72eln+YcYon58p/yFGf8UQr1rKW7YJ+Iagz+JUshoo
eFiI10C2kVRayoNAtJCwFRjGDSZ5O9ws2qmDT+5XO6CbctJQSAgHVHvYh6B/o+M9
at9AcRwAI9WhZZDPV0WNqU/YEbq0GpGehe7r/ivaUgeCTKoHrXbtHaXSmNLyXsdU
yWrWNlI2sMW1VP1lBZo/qqp3COgn8bHu0drnIMLF7O7RD220+QOmPL40GE9Fexl0
zdH4sL/3Sf7yb3CKPUbPi0YEKTzPGDTc4Ta0xIzirbZ0Ejo4PynrOx3D+F1E4qFV
LSJav0yNHo/mrcpuYR/+T4c8sryZ40WFw9GUQtzsFUmYfUQMaNX51jL0+btyyEb3
62VtyEWdXrOL6VVNoJ8K7cEsxubj1pnz7/9HzzjUUANNxX2CJT2MVazmA2wqULTu
B2FPsyDraEzdksKUPWjDUkrMwIa/9HSeumh94T+Q4Rq15KIMkWcKXKTo/ydjeEHN
j1y6NHp7WbB3GsR4vfpYDUt3x/lF1OiyCXujUItQtjQjhP8KjTtn2RXuuTFMeUUL
bVImIGD8u91V/BJk4glIbvEwcvbywW7OM3mSAEonQrn3O1Nncun1CXOxi2ykDIxh
2trcMCEvZZEig1Rum2fI+CJzi9yy/a8MBebElr65T/5QZT4vlwyPS1w2jiTLp4TT
SQgTSV4NAvd4WPPz2wveb8dzAO4u/e7Rp+EvKL1BiC98YMJdiA7K6vPV1+2YIs3C
hovDejJ+J1bR6xxmh8b7JZg+EvAEO6Jwl4j6aO/AtS87E291YJu4XTrpT1WGF3GU
0bGyXA1TDOIo+esWnk7n7/7iBtTVc8w++VaR1RmcBPREUp2jlM60VzZGmgolSWui
KHWSok6eiXM0g4oEnWIsj5Cb8fqrYmdFe446gq/WyDBKvjHh0FOMpPqjpRcv9FFW
iBQgaxl/YkY7fXQYXMgDqnEDla8KOO6Am9XdLm1zfZAtJdI5pO1QHAeQom9+bwSL
gefBPD+h9g5H9XpJL0QO5dctDhhlxER/9stEidbmeWx8NQ04vy9L4zMBX2V/EFr2
wfP9G7P/p0CVGbqyEajWwnr1/HzCquPlfe6fx+/rz7/TmwKlg9CvdrpVClovjG/z
yNt38468UFgEQ4h8Vp8f9fIeW9S5wVpCHh6Wl+qhS1qsA5oaPNqrzAkO8u2eMsgW
KrA+Ae897qu95wtHmlpzNyK2pY0F/MRnky0LLnqRVOB34bQC70LEdO9P0v7IgiDS
8puYS0iRLUj1vSBiIuK5AQji+mUKK51ecV1RGxEi9woIFeB9jUuKZLA9LaIiP+NF
J8Vw3p8HA5hX/omrD8QMpy8HT6uKpEVYpKMQvfdJBBtuWaq6ujzqvkxc7GOSoZYG
+5SBmQtmYdHhTLJiqb69+xyMFn+U/vdLliSES61SX/D28XZVUubLe56GzIHHIl4x
aceOgA+ReBtZREU3TD7MJha1t2zpGhJ7nvdBNvlDhiJ+nZBuXrVB6Svufgx+NMTO
9Mwx8g7AdmthlqI5utALoN70f2t5vtxZ0Z7VXr+767TtNnlEWaWDj4+PgVJTHuAX
+/nKvYSaVWwHVX9bhcgu1vRztTuYeotA9uw7Q10MiHoz0i7XvKasB60uCPy96wWN
4hDiJ0tdnp79ZXfFJ/DgBz8tDvFQkt/EVOO3iDQcZzG4QHBfyVMLqHUbzCPc5b3l
Y7np8nD+5NkhmwqsM1SIwgY3db0z9qxc2BUJJkoeRhlMsEIQA8Ac+hEW4Ywz4u04
F92za8zni24Bge4acmyvRSmGk2+hvtEI85vEwffRjEieeU7VbEQSmUZrkcLGKcvG
0KeK7yEnpdi2XVF4DCp4FZSKm+BO4R1R1a0SUkSNB1pFHtM1oR1ui72/xu+7Sde+
jmEecNXohiyb5/OmfEiKmVwXaW4Kdp0VsWe/1X44SN+EmDK0Ivd7+U5U+O0BsBBd
G7e/pAtzh6mWdhGUx3J6aP2jbI/GEdWaSHEvJB2sOVcEvL1iPiD3BQWfoMfoiJzV
PUz2yVApmmUF9Z5dRvjSa7fSL0npNgIDAaZp7AZBuY/DLHZtfm+ReSK3IsJ05OvE
gC9m1tJ6AntebAi7mGfYCFy62a6zBmfx5txYaJegsMUmwBxP3bD4xzCHVHFHY0dP
eLo6alt8Jd2qM7IFFaea2yLgTk7ecnwki858Xh3ZE6mgAq5ifqjrU141ArVeuW+F
7y1EpvgvfnGent4bttjGqdJEEe/suBvIDBbDxul9vgGTtFzGGlC7cAwZ5SgEpOci
7GISVzLmx+X0mEDivQQ1r11Lwg7ByOOab1qlaL1nPheA+N0xG6UamSxpRCOEkm9M
wBqF3ObikE8Yr++KxiexqDwsbidjWvewauGSJKWYbK1zAhQdVCh2bX8jeirsm/zB
QdBemIGsFEXJqT4yrcxTW2cRBxNlGdgVdyK9pdqe2w286Ocaul2VdbyCFCx86vob
G52gR38E4VRlf3yoTw8jqMkpenslfajfg+R3al0WptNF6/nenXeRhD2/XgiUoiqo
lqsaii9s/FVl5Cpo0PhrP4Vq7n389iG6nb8NNTbBGDgXMK+3RrAZ0Z3d0RCvhchH
URMdZjLL6+QeI947rG2B0hhBRaXnP3xk+fxSAbSJyLKizBJDGeiQOEJzckcCymvu
vvcm2Xc95zCKiLSLVEEt+nrBObPoTYJvLjoacMlymWv2+UkFvFRtQJbayahCWHBm
3uyisTAntEHfg6t5iMR8p+qASTvFePP2JXJGNN/VCsEuWOppyluBpcdQcwEL4XdY
At2PDV1HJ2h3xo7gIh1DU4HCrFH3TdtMrcCWzKioJU3RXXzT0k77qy5Giw7y4mwd
pg9uVCTsM7iO47Rh8RaJ+3KYdy7lRkaumAY2PBMC+ciwZZ69/N1Sb467nkKLQYxg
akNUkWgQLcq6g5MUHBu91Jp0jvuGhZI64XRIiH/voArdCrCSOnOJ79Le+S2SGEAz
kd0l7vVkHrbpVwJa6u9mDfp3W7s3htatVMHIPHNAmO5U+8jJczWz8g4MxXGDWVKS
njJkwcJRhVVmITfroN2aovRe0N7VjnJbIb99O6JCYIFnj+dbHkrvIuV8t23ewNG/
3NcU9hGEpALQocnEuV5AdlBRBo+eRaqibkeF2Fk2mk4KaSW7nYB6L9LEeU5EXDl9
dNdJtbaQG2vQiQ6N57Ga48xS1p/LYMZpDp1xM9FnmglAATquVTE6/jTunnMwyFNA
y8x06cR8EE0cc1QZESnI/d9f2Mz09y2LLwRGkOEzqESC/n6fY+HtQcYpXYA81THO
JFSZt+FbB5lQHm8pGOZTHLeCrRRFaRK6TsJ54kaharhfzliXZpdVDf1YDgK5eswd
c7kdRqK7gV9R7tjkvegqYgRfhT73gRvBGQN5rgJk44CdVN93LY2/S7dewPPnAIHP
JOBrRTnCB4k0ALK1cM8ph4/7gKzV98ZrZVQIA6jsPqwpyF67j7F/1YL7QmWyVDkA
m/8jwL6X+vBK4jVmeAt0WjAkVlC+9e8RdX52Dcs7OpAJesZet6bpl4EJ3kZ0PQ+J
gbjjLWvYfnJ2/8qukwjYMdhPhC11+4k+UX8jwI2kmZq5BHj9+Xrlz46iPAdB0k5n
vUDP+8oeeeCoC8deaU/jzGqd9ReaPMnloenbwEeDpFyxIBTXpWatOiZPw9fP0/e5
VLGyiv943p3gsq7Y52QF2wRyYQzzuB96KYzp3iCB+1Nqsb4sGrFFM/jAgfzbykYM
Wc4arl/NuEzdQBXv3V6YyPipcFaNoJL86nUzkbK8tRNzwEnXCTr5kgi42mvyixYE
HNRgrSpRVRtU8LI83qIOxqK9lKamcJwuJ9cEPOMWhgyPWKNz/pNvgIRF6pvMWv+T
AOjnTUpLexoYl9r/+AePcZ9/GsX0gb1c0640rVc41823nzzxjp8XjmNk0CfRiVBj
1FQ3HyH5oCBX2TlC4i+sbFye663nUxT9smJ6iaoUQjzEsqc6Iz40T3Wf+sucnKGZ
8bG4cBBU/L1J+WIbwo84Xe7+SWVpZlppl+ar1HCh7ygOhlykLisAU8eqyk6umpo8
k2w92DCkjC5IsjkQLYfokzp7faIsGMMnpHKYelZUqws67DtpzxTpCJcvFCuu2pdi
sOu5MYJ0p3wEX2KLviQtSG3Iy+qZyQYYCSGRLi0RJlkldmrlxc769tajNnSYW4g5
n2l0Et0UPpYGPrWDafhkNwJYJwM91zT89aCF+TVnkLK/9jidVlgib21NbamGVrIl
92NrXMvCS2ERAhuqIHAYBKXW5idDSI/PjCom+eDhNEql9MIs+TGFYEuaATudwoXx
Z4UDcuoEaHG7l7GxBJL017Ri4DhLtG3BYARvtVMFXNn7hdsKJ+njpr7y3AMUhHgr
4FwIsioDA8Y3W66nRPGEdLtKOxIF53xvRI9nXr/1Hat3MVAzwGHTo3Gkd/ULnW7R
gnYWMvSmZv9dtsLv6ynkHY4vqO76MhMUxA5ACOpoKm9pMmlYlJOeXXWGd1ZGOXE2
1TXx9csa3nq1vUhjMZTSa5u3QdbqJwhewCMjDGb8SnzTtLGDGeVmDcCA93fMZe4b
ChOCFLk/0xj9hs4UJhuq+tdf64oNzC9EkrQ605VbClhm6OqcARTKbN2eI40vHVEl
nx8KlVJblO3Otkv3o0p0uS2+xGkPyKTWjviwyEEMqMRK+qUVEbiuo2I2PH1COQGV
4jn/hFJX4Asg1G3QcYB1PP4x3Oi/wnf0heQXoZcuzyQ81PH5QCYkd5X/ObBEgjPA
zt8pQSbTFDMUKm54uRgDoCbYqfaW2mH2wWQ2G4y1ebGUHulSCMbCVVe4OCFt2Cq0
Npxv2Lbp5CVU7OkmN5Zfia8KesLlrcPa5KyWOhlulbHcC4UAbYeG+iwNZylzPZLR
/Cwv76/WdC+giOrp0bejfo3bjVmuZ55GvFIxqeQm9mDSUlrAomvf48rcJOiuTsX5
eqwslAQ+A+//tDLPyagLlMknpZHpMCnA8AjTuxCBJYXfAHQzfSgqnQMPqzUz4qiW
gDc9VfxCrNoCbI9CRdKrJ1eit6UE6cKCEiMetZ+S84DM/7Pof4P5u3m6DYiYi6Xj
ywnY3KzwtrMxlG/UiIB9rrq6wJCQ2n2ZeTPMS7cw6YJk8Cl93yy8mr0UslQOIJ6B
uxAUrhorGXM1rDh7pCqU95PamUAq1j8ctfsjoqrZp5w6srjBXrnpJrjhYdsIzH5c
MNP7YArcWSxWq0rdfyrlxERVORV24WsPu4YuFN9cMJ19yIyggDeVWcNJHAOCuZvE
InaPwPI8GVv3u6m9boxruJ+JuVyTDKEZK4LLYI376zoGdAfED+3yN7kptrlxVtSt
3HfiVvW/fzHGnX9Aj27losHZyqi3sTqBSGlxKFGpF8ddxrP1wTV+ZkaQs+iCtWYT
YxGRQBvqGwtf5rnyYs8nzI3qir0WJG9OLAEIlEeHGb1sZ1eRQ2vbzcjhzIBNum/N
EbLxikSHlCal/F3Fee5KY9bW7g1L8u+LGBYdowsoYZpgd76cmULqfQjMYj/voOh2
halgSsuwKT1lCa5s2MGEAkLiyAfuD70blCJEzneo6yEv/rry/vb/BFxVkd8iKCOM
Y/Mnlq2h3nh5Zk8NtjL5Oc0MhLXbfQadHgoq8rxYzfmT7yF8vlcqAQQKi/hqpThy
aw6a72L7kkIvVPtXvEWdD0S3IEanTGsvvwfZ9RQT+fpUp5SAbwid/4EQZYP3wr7f
AyKWKjiHx09zjCTZ1PpVSEbtDcQootFTBhG8G8dUj+ujsqrVH7908ybKBU436HXc
bOvQC50dOadQs4LsKOUkviaoZb8S5we1rR+IHXqofYCIwcV7//EWGmk0tT8p1zVV
kZUl0MZt2OoqUf9VDEZc1IvP1sUzbBD8ouMxK4G7yTMlfLQ6BT0Z4XYbAVlhF519
GgFKO1eerwhZBFGcK5YnqHzEHUMxnnEgg41GKROhIwYWiuLEd8nsbTA1w5dZVOlH
PTQyJYtr9KEppCeRnPKXOf9vObx5DZEL+CTq2b+NJqo6NbQ/EdQtcOFmr0YsVxZx
vZB+h8kLRRLU9LmDkb6QKq66qgscRLoKNKHTm1VAWe8GlWmAUhssHOorb0Rn2alq
uYopHzA/Ae5SsgLRcHOWpfy+U4wkYbzCaiEGG6FTwEFw3sRFp5TgoQf0MIRv7oHT
BteWHx6mZFWWuT3BcKviDPYsV1Mvs6LSe2a8aPbi+NmoOjmyx0Ke1yvGiICx8fm8
hkiUGUw4PuG0iTh1lpvF3iHWbcD0fnmIR5JlaAXPWXegHo9DwJQ2mGCCprs8L2gi
9u9AZzeVtMzoOKn3gzq9Z+Aw41L3RUtoG6KYrPAOz10zL0jMd0bWOEH9uZ6cvgE3
IPwN7PYKCYirxZJ2OClG6d9xp3i9CRaWfUzpDbFU+v92z2NT7/5ALYOPKU4iln4W
6Ax3EPusIxEtiEIxjypY/oDzjz1YeSPYkYhf7yYVQe97Urtt38HrlUOSIimmUGbP
2mkd9mlYYtFP2qGx7zeW248g2gtdbEvdPIrpmANGK7nAh/gmkZgU20gIW64mbge3
PwjbCsahsL8d4RAU9MacX4pEFInwFQ/V3yEYrHmHGqQPwYSCdTmOJSDJ5uebxy3T
oInvZG3uXR7QPu6xYzKP1qxO2bog5h8k9knjAV4cNySSnYgVXyp+6lxTC09dC1lt
OM/4NHGMNm+f+dI8rYVKqNSZP4mOZJa2DZIE2V+PO9rlqIdenjujwmo1PEDQq8mm
AjJo2/qZ/s5WD1obx5UxzSux+IbHQ2v+YwCgGQSGhtkIMW9oWnWB+4k6F4QpjqEc
Lh7zUZdgLbY/F+8q4B5zGtPCo2rK78VNKXO2U81KT604u3Z0BlSl8tWelEXaQ9p7
MwDFPJx5+1wMdOTYWcEKk1xdk+VWHqtUSSc136mdvF1z76de4IxYmpwqlOywz70J
oDM/BieNfIjjrrJEI+sgEPnvK5rn1NBUzzAjvIMJ0sBBj/abt9RdDPIi8QoFKL/Y
/5CNed8H82obcGEUnxf31xX2d+PsQWMfjKb+80Xr7FbNmE+2gBjZ44w/4JMcV/nw
0/qoHpgcI5yJZflqnh8/qwwNkcOw+GL5+vvhZOe66aL0S0ZjtBswpOGNEMvkwAuJ
6n3lpG5MWS1e0W19vhYSo32Ksl4LQrVzZv1oVILhw2CeW2fZtoh3s2nUEYS6nIcS
HVHiFjLS98T1MXKpZBu4Utd8OY6vbxoJ7CgoTl0SX5YOL8UjGQUVERG/wK9yCT7c
0h4j1RbLsYdZSQaOemtM8QRlw0RjDo91UK1jpfaIQHCIRFsYUbtLg5MAqm1P6qFv
8qwhJkuEwrpV3Qznxu7+8GvF/o2YExlMXCu8laEUJpgZxgsHj1RkH0I92UoJnAMk
VNEyjXlN52lruxTutuMxkPGki7TkzKXXObGyPgTSp6VdL/v2i9zggm715QEhdlvM
KRCsvOuqzNeN3v5UcrdqOROOLgAtowLssSYdBuJNdJZhSrjPlmjYuo8lgEUjbO+I
RHa9L+4zRdWOZ7Gpa+q2S7sX7yyuFIxxxDlZyZQPt25S6nnhBh0b5xEjbkWi2f2I
VzIMblredp0FIcLWCrPxI4fGCU+fXZ80RoyuGIPvPlxdyWQ1dxdMk1an9hG23132
k5UbAFvxGmeLzMOU7lvMz9HVbIucd/35AWKcRDMty2aD36GJv5HxojhFDehZO9VK
a2+VDs1CEpNWAiLeVywGRkBpoHuzf5ipYYCs/xAAo6Vjaa8M1XfEP/+R9gZaazGF
zyWudzGuN/+eHxXD4Q2vWe8yWkW3jJM56KNYk9U1GxFxC8CdqLLa0J8UrGZSGCkj
bYkUCleZt0JcWF+6yR8Kfk7Nz9oA4uMrN1e9hweK0ZJNJnNj1U5Y0EmIq6EiwO6M
HMv9nE/lS/jTClM2AiSVo8QNeb8HbV7/ZbAdYfMyf6asD0+gDuDznN7scLSqOX3m
K4sJrdAPPM9Mr1OmN4VCC+QsaFzkuHllq0jWrnrrnzxtZf6rIR875VFlCrcOKmtS
qcpj4qnrA0KbqjFRattOYGCzMVylUtgGSK/YKsWDzGS1+yqtMVWMVfn/ynZnvxP3
kZj6Clq4jzyKgSi3vO9M0z41bScICaTDZrzlnogYivuaWCWQpvbO6ie3x13hqO/n
XKjc7/Gf4+WTDUXk9TYw279oGi+n5mifGNddoaW4LFutAd97159MDIL/17fg1b/t
T2bwlSX+89WUB4+WpC7zhaZ067kr3M1ZegoIW0dw+TojepWBBPNmhrAnjzK0vw/V
vGjs/iTbxcnwPeGTNx+/gx5AiMuF6zPhHdC76q7jT3Ge+vRsrXiKYfgjkSullrNv
z2vKs5MEbxAv7RD3w51xjvOPgkaiSz8gch92j4N+0KsBv+3ub5W2TF/ZFkjtz6wO
JiZeOjOriUTTiNGbXP2qJEyVYVaJGAMSC6Eb78J2bcLBrmV3tkzRqvEE+yatjPnR
cZO4h0JYY4V9djR1YVZyIAxFhvMC4rk/95UZnh6anfe1CNj8pE28BhuG6ATiBMI/
9ttFFig1ckkXK9QTNoZNPniBw8H7y+DyFipVSIp2SYL71tx69UTRxJjkSS9m+eEt
YhMraGPpcGOlxE1epyDYZk+WgJhE6Vc9Lwtw6ZR4IA/xxIjJBFUz1SDuW7TAhgok
ZxL2cnGLOvgDP7IcKTCRkgHCdzGyGC4bKl2/8Wt90IqPTVHEj/V4NrSd8WPCteOE
xBmlDKAIw3dj+SXggHHvnDlnSt+VUSer7ttVfXOXPCGuAV4an2+UI4qFFcXYd64z
u6tHWtgRM2UDpjYnX+mh64MYfqYwWR8NIswhhG7P9oZuSUALZpK6kMvzaDF7+LPY
Jr18faBSfubXAQGRWQK73fB83WXc7A5l5vDqs3L3m6mYx6yAwb39KSyaaf5fG2tV
puwjCAtuUGGHy2OhdqTv8oiYu3V+7BfCxANWWz0VauGOOT7JCEjoP+fSCb9MYiyn
L6Y1li+bf+/uuQPS6ya6Wl6wCzk3oqPfpNf2/CgjPcqXJk18336S/Xhd81QTKKwo
ZOG3zI2XvLEO6IX47l/9nql3l5bjmCQBPgeIXsftAnwJ/Wkw1qjtM0Zt3OCZStqx
VUglmW7L05bo2mGXtHmwVBAfqsanzS9poaeg6e2S2GCso+z5wYUcgdX3mJu/g37c
jBQpmpSmG287NNCocw6JDRtkparF4hGKQGUcSVHQAxjbQXxv+5GAXOa7Mtq3q4bg
vL0C+tTwDZU3Oa0S4wCZJgLVLeChTo1EzlGaf/YxW5ctRphntU8o46BEWoxrsKah
Kv29saPkwo8b1XJc6GVlrmrf5DcqSviwJQG9I2Gaw4/klcIvoJbbTI5XDswy4uyn
qBw7hDA5CswNkqgfmeP6Fx8L2X7Hgkh4kdUL0YDEVjFcNrMaVyptaC9dTaNaGesS
phxqBI3Pf8FrIO+IfWZo56LqvC6lDDX/QgLsJp9WqKia6n+x0yuERwRSpUcDewmt
JC5opml1mn2t8Iad1/n/qT7dwQwTSy5Zc4Vhs9eTu5W0m7tAFORihnyqGVW5DtO5
Fu2W0v3xVCJ8RufsvLeKxss0GeDEN1M88AYvGzdDE6zONoSgM9IqHD314SPeDvfm
EYVaQgJMuOoy+hFr5sLgjhpOKsIe+sXgE8uLj86QADBET9ThM6mJLtC8TgasGCXu
/8TcWwIjfRZuZD49aPi1OusRBDENPdOn20MKs22IXJ/d8CwSWLzr0RjjICAlkYFy
/YJKFO3Ywj+LfyL+yck8daiQe1ddbtcCAbhVv5b74+dhkGZuFyAE0bRwwtMIlKa6
yRYLLJAlHnIgt6ZTezuh7TiSQqggiYIDCKC6Sr27i6hse6M55KoC82f3NwTVVikN
bv/4T3cCAVezYjlnK3WG6+ycjL7eolaVWUhZTsyckIO0muRIziwu7tpZ9LyR/tuV
Opo8LFGYpJDMJplX7hrU8+9DmhpRgrXgQBliiRKHEJaGkzoARMgGROLxrDB8Qw6z
krI5gfQtKyxIyW3GqTqt5S69QTYEzWWtvjMIcAYihRAR8rrCoOymsiarnAd9u+Vu
rk9YFhFVU2do1MCwwkJ+tGXxtmNjyvBVpLrADpkzAcO2pzhBlA2Hd1I3To8B6ROw
Ft8s+zYUVsOmfCd4LKAx9E9egCGT2oiA1pEWSkuRWkVv+4W4d4zI2sBKCbvxwpnV
7LcJsjiEq7ChsDnA9eNzx2YzW2nWNJrBE50I2dF+ZOVnPMVGPM8ysguKYZJYO1bT
ThusqQ1zaKDg/qJ/qsiSQf7HYWRI9iEea9hgxLcSb57vReDrEZBThaRe/XIjFzJd
WfYk/LTTxGa1v5S4yYRSkoEBEiwYtqCEH32vSChOiEgUDegZuInu4Mbr+gBqQ2z+
X2GUnTCNNUXmQn6L7AG+XgERVehB8MD08yrMstHOlWyBt+lVI/FlgXvLUPDrKjB8
PPTrxs1/e4QYNe1k8FZZpdx27vl+sTkgeQPWnQ2qhlZpXAv+S5DahnrEJ/VNdcdM
kS6EYRQD6H9E9pXrFWRNCZ9fjE5XLz7E0qtbX9vFph9VTAS3KskG+oXzoOqg6lDn
4u0dUevGwlq+nqNxg8/UZifOLlTq1LqEthq6nqzFbn8i3g97dSh8mEgs6iIIzHkw
s38PhwOUBgNfaZGhAc1RW4/vchGdbAjGuTk4Ps56xNt/gfCdpMZ5FE1pOn6oexGi
JqjLOllDvNpwbo6bxIwk1XFZOLaYVRpKrgrUR1UXmQheE6ZTIc+DZEKnvDI9jyJg
i8DX62IhbP4TZV9n3BrkBygkwkhsd3qX7kiVYe6gSsQZz5gLOxdYf13nx0x5r73r
gLiIja4aXwx6YyST/hIoRXKqwgJhMBT2njpnUJ2doYI6ymsxeufEZSg6/96/sNL5
9wYIdUfzjAfem9hpplF7neT+XINe4ONCUzPApOSU8qQztaZVz5gSFb0QjJQ1vsfh
nfhGQ7zYCkXGKZEUGW2BGAid18u3+NL5X3kuGnmpP2UoiGaG9KrhWzwY5myMz37j
sTy5h/FCUnoMDva/OTdGr/0lbDdf03k3kHcq2AyEYdZ1nmv4YgKAQ3daXkMUA69c
wSv2vWgVk/O/rsK1/9C7qs0EvUbD8B1kF0T+TpTAjDDfr/4fjOvgSX9B4+ytt8I+
ULn8dhUuseWWkegmkRgAjyXJiZRSdT6EqoIxQv3GiO7osytuyxkL0CLja5QSaiaC
VjjqFUnj7ZCszBy5tud5q4ON0k8pTpYdWu9g0jtZC5TsXSF/yXB3Y7JRKJLlVEuA
V3tjq6JxIXG9jGNSCKGnpc/oFPZChLLRHFqhmd4D54URHXYT6HOX13DVRPAaXqU+
FakVrP8Nc4mTzOEEdqNBcpCz8UsjjTk7pJRWyAc3aGQj9eH3c61fNwI8g40YlqQG
eezekUNIiZHV0BJEzInk45u6MKxq5xNqavtnyfCeJim2zkSJLQfiOaCtd/lbS1+H
T36o+L036BuGX5l6uXqvnROn4KMA270meZXdc1mJ1cmT8gSfvvGDo4Msj1p2tuNv
y6AYjLCgsuLgjck0wBQ2S2dK79gDAVpJg1MovST0msE633G0pKZvFGrnJ2GZc1+/
k6PqAhSxwoL1pavOo0Q1Qg8QItVFbHXefv5fB8wBBxO0mNHRAoNyu23iXBcUtkp7
mvp/oi/+THIxtE2VBVxSf+knRy4PIARgDFw6tPCVaJbj64yrcKpcpu8ui8m+gDgJ
eBTspujQVSBHRq2jfhthvTb+rnUgov+svUcp1b/BGsOtsGP31plX4ssraKsJKqty
DemuUGUdCZorRMQudYqdJSCE1ZPTWdYgJxJKjzzmHuiekVqc2eGMIQRHHASTRobn
R4lJeIzuFqmASrjcQ2zQE+vJC3Jb39mHrZOEYOMoQtl5l8qsuQMjS41ooAdUCmW/
z72Es4aVfhyE2K8C6xQjGYczET6bVkNBEzzWEhFLLJoytt+BLP5jVT8s5134Zete
G3oJ4hEjqamPSwU5iAcFqZWZkPM3opWKaf3ol4XP5pcb+YMUzvaO7qN0aw22puYK
O6Tp45ZGiqfF+Nuj09sR7JbLiOTHGOUCyF6jI7Vy2+LoSLs8/XfE2/gM9aAjVImv
oi8y/n53W8I500y97d+I/4DLVzCMROLbq/cQHuophVScXBDlOclIXr9SpFS/N0v3
Yp5vu2ET9yoZgL56l4EoWdql47+loeusRmXSSADU1ZrQp5BhlK6EzNJGySf+tqoh
yNqehCIdq6g5H+kJ8NlMhKGyzLQkNsFx8liTlYSfC2xlD+RbwIhwv+XT8ZWb41rL
wwpaGNCEHPExFxXyY4kNjyH0tcOgRagQ91jJauYUQnPcKWw6pNCLQE/FMFkJPhUE
dDetv4FElOr3ezCWl/k5ygxvYTOciF4snyd9JyIteQBFRuDvkJ1NfHCWq6iO7rTC
pvDyn3THjyXrWHFiKTfiXxqn+lZOW69MUkO+JLPjG5GmqYCcYAOcBWZO4A9xSQYW
0cpTjDA17F6npkHI46GygCgASVfxJNYDOtoRI+yqGRFevsItsAAu7Vj/6rfKXNhG
bT7BBGfhAAu+Ux+FCE1FJCad6OXFLqgUiuAtbNY2ERtL0XEd/xVWKdUOThezlUnt
5lgr+zKzWr6rT6Jbbnp1fSrL/dcSygFRuyk6ZkS1ueagBopHQZ/O1to612iHSITh
acB7MD4aJP+hwGq3VsOowuo4nEyZGe4qPOid+bNo8Dy2SNnduGEqKbkpmvWKTA24
OZU/xWo1nOEb/wPXJ+ETbHXox9p/6YXnG0PgjdnBf1wsT4ErrbY0f2mPv3MueeUb
Rhbk4WlsmbuxwM627vd/pj2+ZjY+knKPfyelAPeb1nAMLdJvTBJylWUTIyELLfgw
IMoYwhouZjXcD232HyeHzBGqumk6k6dXIlhpAvi4u+gmwwwiMLTXms6LVvG9m2y7
BzOuze/veFxsSkuAbEu2G1xUIloksaLc8tp87pF6z1SIf3Y9Wge8AKjxVSX/C+x2
dKKcEC27ueZXPlmmqhfO+4LpwQkBp/p2OcUyoOs+17qGmXZbiiI2LVwleLArzvMW
vj2g/Y9wQqRu2lod1c2fUOYZmIE2tMkMPKbcRDUCXMXLVCCVo56wG5BdJ96Vunf6
cyHu2lLk6D6HwJMycquuOF+B67Zb/e9fKQ6gcu/L2jf+GSR1gCqsTU12+t9G9Xg/
/H+BkIkZ4VJZ4vDt1qy+OgEXKt0hBRE0cR9vo19qj1dlEHuYBk3JG5RszV1yGHdn
TbpcF8K2DGJOIfnLP43DlGVAUmudQ1LZK3kLrP5fnNzssYlh1Xo9TdmbuldMWOWd
OEBe4BrJlEhiKaq9rrA+j1FxZ2O9QQLvWM+7tJMXrKrcMG4rdsdfZ5kckrpV8CB9
rD4QvAazr2v3kPeUm3kLj29VM56X1F7PiOIqvgaH4LpOcEqKlPd7EQQB62sTT8ye
0GEqcHfHFckL4WXDXyyPC5tQiJQua2q5JPwk6M19ilyMREQ9PCfdleBGzsRLnM3k
686JywXtvgFVVoSFiN01FmfRF/iNPd1vUqqpdlZH27oGW0Tb7g4zSNyxQfqIepjS
ixaEYunFPFTQMoeMSBEHI5XIx328KTxD1fevMJjsil8RpbeT62jHYmfbGGRuywR0
kDW32lObm76ktKOrgvVc+3ePGeRW+3kSSthBGC4zOWkHpPgYSjw4arlstSZ6wNHh
6qFB4vTGG8pw7/CG17G7xkGYIlatpLIIdEQsk4YiYv05H1P8l+yj5XagX96UHVe5
w3MDP8zsejqRU26sp4H0PZBKkLbbJGhlRbNLUFj5Abahv01FNScsDCSHEcFAYXhv
L2Q0a2H7YMyg7s7pW08kCnsV64Q7M1nLYqTAoINNiIGlRcJ1oqntycdzgBsMz1OX
eOZ1A2fGWJYRfBGDvPfuayQWS1AMBxtyIs1yESKVA777hJ3u478epKn7vo7YqYVX
l2rVnqTrmzcOxplOE5aifo2xNWYepqP5cZqdBz7cNc6/V9BIeAX79f768YtTEq/m
5/gBmlQ9bjLB1GRgZ+jSeCHPQvs+bw7FXtRxChofsn2nJGlkeFq3u1qHjfYlBSus
yazjxG63lL4mdXbcD1YxKlG7d33n57ZS8kwV6tJXhJzM4Rf2ftXHCdjXPfR0YeqP
UG9L3rdp4uo2h1+eDQ0jdwdPf67lU5LTPe+Irebupf3HemBoT0vrSVskMdkOMuM/
21esk/sj2LhRsjZWwC4ileB5+KOgTwk5LCdPki8yp46REdU1VbBQ+00hAizL0VhZ
21sj4Ri/6vvD0gmlkE5EDZwq/iLrQ2eyhhjnnarv3s+h67bCjb8Y6Bm+vZawV5aI
9MA+fBpQhMpHmRtvFHM+cr2A/IgSeBWi9AQDUuvvklhSDn5HPDDXZ59V3RsuTjr2
5kak/OWpXqVMgSmBGAdLeXIHsA/4Oo74RUnaTfy3q9uzLrtRbZ47sPGTOPXAgqYC
IFwIVO5rXhseRPOK4jNKA55tzEWcIoAzJMwjapGXOHrX6zO5F4raijZLILMcHllM
x8WmxP+R0Yzew0q800bW+A96qbRlG3EfPkpy67RZ5B4v4xo5l925lCp1ZmnRfUr8
8pjKLZKsb/WmnUgANyb1ucP7lrYCKJBrMHmlyuZrp9IMwmznIpsTlMQUXbmNrMaa
gEnXZePci7qMr9uxn234XlLpUqWNO5RPDRqRJFVwlEWhDcDY7i5eA6QKUQdB1ZDU
1uL4/JPBTgLHVRYh+onb+FxGOAR8pganAuSjHq5IupKramMUi7n/KSjArXdG2c5+
z1kl6wOOunRUCQelF3yo7hFKndQZbmAmIDmvSTGh1W0dyV4O5ZSq3Qn5UsqOxNSA
LXW23eqFTEuA9YJr+lcHXfZk1gZCD3JR3Z2yh4u+GGcLLN2GDfj+MzKbZO9DnUXS
OckelaOzi0azN1uPaqRV7zBfVo27ib29IHt+b18iZ9sjXc1iPDl2ygJf9AAPiCf/
1WozrVJGVQRIlYwdUmqOCGv9HQZykMpRqGEByGmQc88SLrRCJdRoChjjj4lMKMIF
j/OjtIrky9OKSzB7JdFETXU4QQVmAG/aSwnN0X6OWephGqSCcr/N+yWoH490vS1y
PYMWoNtL+BT3en5FmnRO2JOsoOskuQEfgmVsvdeCqNYh/AXJScZjKpqED63YYpC8
mTeOaoFQHaAsgyRXZk3/ndE7h7uz8XjUW0Wq3hPHVeiWz3xTpZNXTkGad12agw9z
5kU9iw2TdO580C2WflS+vqghu4hO4YTpx9cyOJbdmrVVierK9GSaeJWNHBvPUCys
4nDhAbT7TAtGsvuzIUOZJwDlhPOcnEW9WQEWXkvLi/ScrgFqQZ6OMZyfPCklTFvo
UMHC9Vf4CjGn32HR5HBegyCogGI+mdJDl5IizI0fWf5t7zik7nVMGgrPsP+Qfew3
v7dXrTQMMrSDqwWQb8UTn6le8NQhy0HvzA53cuk3c/OIrR7EHp03eO1o1EOQaMr4
LfvBWibmvtMouV2oGAaaZXCqezSsu1LZ3u0mOoq+2fLfEITEiZlqbtmlJrl7+88E
Q8mz3LRF7ry+Xh40i8fzhnUS3EEONTTSJRfHLpFKkc5YpMIYfjUtB1KWvuJAU0f/
GxG/Tg6W56SVmvw/ZftB3NZUqc8n1bY/1/6tbvOTsczaTiQzPUuZcYJhRZC7t+LQ
CXm7vlWXrp7gKtdebgD8Em2wCjr5lkc9NyciEsZhd46gSPrRCBAPr3Mj7ddLkeGY
ivA6oHCA4osFVGadZN/lMq48QvFgmsASAGixqVz/UYJhw2y/Ty0tly9Is9/qXIM3
SpxMF6SZqRtqHi81DWYw9+6nxFK+3T2zf8pe0fk3fsTeBzJQgq0PxoPiVEYyP+T5
CVNoEmqiNAThnmqTWRDd2JJ4W8lqNqGgl3vv2Z3Ve+8+fwP2dt7YE1x4JHAliPOj
xwmH0bTXRD1FF2nAUj9V5CF2t7zeiuk3TxQiw4HY1muL1SDNyYhMT96P70VvodI6
zY4bPyM8hJS0u6GQy0QJe/D2AaEWuBytVMkVoajlsQrFDTtKHnZDembi2b73ZtcB
x8EXou5jmMyeDSIeE0voj/Cth7waNuH81GF0evu6ffqPB5haw9kFksxcTC6yGJo3
FglVxCt/J3uV6zBTwkHMv6oYehSW2vXEwS/a2o5Zr04apT6HGmQl+54xaZWLADZg
GJRAR+jSwpME/ZWNCmCSA8qC/AiumQ8YhAn3dr9LvnBLh/EtYf6wlOUzJqsFJUbF
3mmyu2vRhNM1xH6gQ7av/XJfxqpoVOj1sjWIRvOsG402VkQ4FX/z1odarRf+v8ko
061Mfptps/qsmGg9XXvMPsymdh/alSlho1iUV2/msrV6JLfwYdEAYVu8u6K5zgzy
O6ZTxDHEZMb/aSjolI/TecWcoNDS8X2lcKST1OiIWnTkoVIVPiVtgpQfxOw+1eHN
f4uyDX563dmRNJNrWsY1k9IYN3LT4VwTalE74ZO/UON4JE1jrMJ4HmcZq+dSIkN4
uH2rDqQhYPEX+CnVGbbE0Mn6Gh3rFNu9yN1+rlTaoMIZcZxmc8lz1eny6SutOsUH
ZXO1HSFDaImW2oH0tFt33hxSwKTiIjYhi9m9F6RW597bnzbUUMYpMOJ2vMM8i/UA
8RMBGXTq86nZZZcGN2zcF3XVcAFmkIXFP4YAC+8WxXEUh6iQ1L0wzV0g96F0WA74
BNWsrnnZiCb+ApLnef2Iu5uYbjEGqeMLzMvHDQBu8Boh5nLYikckoEoeX+BwXWRh
EcwI6+9W3XqH8Y/UVdxB8J8c89wDwpdaCoTBAKa3Q1tW0q6k9pa/B3PrHJIZ/+Zs
2NwEcbc2P5eo5ogdKn5kO6Z04GtQ5i4JpPfmcvyJIRLDTiW+5Tej2TFvVHu8JhZR
gGmK6kECa0AVgbwNaWu3GGkfm9c0xuj4bBsKrvNGKxRPdVtaTBO6UP4mSlYX36xf
+cCwY/4EkVhW4KXgRoRnGA5uX2L7ePd4EMtjWj/9w7c/WgtraySInuJ+GiH99W3n
C95WvJjE8kmfxEdsPGbnmGz6CXQv9lenMnDvMhFV9lGFNDCzAPA7DEdZQbiF0+0I
RjfcGocePp/+bj7MeaaaSTkbEYdQqeWle86VMrI+66n9+Q6GVCZ3g8BxBW2/OeOG
53D2egM9Ft4uBGt1opRtsD6cftznKIYC/L4nwG3yUs/EGXuZZ2EDwb9PYgCIDnJf
Be+cEcvWMMBCqh7gy9lj3/8712X7JSkA//cQJqCnNW9UZDHkHfZiIES/ZXhl/f66
DrHmbUuAYhlM+4CqZ0h2yGF5POETXpzFppJ0YDCKB2CCjMM1FB93DceqKJxyJqKE
2BOLyDcipK5y6/IXQooqqTrs3V3ylssuxE7Yv0nh1dEwDVzaBVsWugOMusX5dUjk
3FFVfX16sMIMja1T1kBzmRL/45PI9S2+41ZxhZKTqtkvLHM6h+q48BgUi4GxxYWk
XVnyF7vkGmlsxdeJ6jGwH7CrwBqeuVo65nVamRT8iPUhbgNVulFOvTAVq3pdq1zx
niCyJKqLQr0dFD3si8zanY0gfVLGLR9o3q8Gx6N8GW2niVF8rSKtTecRwIWlsxg3
/RSd3rfSRjyT3Nsqk2gSwnxJlYSJX14vPr/DOpJjMTsZNv5dLAUES1hqpb9IdEOM
dvPnH9T2/cyXCN+VRLL1U/W9xZxDSYUHnXiLRFWfq8Tr3UVnWsY7H7qqU7+8O4NW
UN8y43ZTfzgBRyxVP+ZXwktDjlPtOEOQhHLefGXVn1H+rBJLs9eMHlqgQiToH4ru
EsSFE5mXtllUISVbaRnitqIvrNUYCIN63rJELFr8hd6ao9Vmednv+HO07aA4bdg4
MYQei7zKhwDUPzrP4rNSAO2x5VHvwcl3Y/rlq+QC51wzCP+hJV8FPrYrVcb0jqKw
RdvG8da77ET+vidHFL3Wtb3BnJppGn6Q+SOj+hN8kE0STrIoj19EwObkYRKgbtD8
Z6Iw5rFia7ZqahmoJLN5HeBzjGjKuxg69oN7ldVhxZjCuGRx5K/t6R5GBhYLvgk+
trJNpDZmQnBwa4IjNEeGM/Khp5HDXKqy+ynYf0kosYZjJk2Ir+cMUmXyNZ+/OUmr
PbPu5WGwEWTFi5WXHTXdEFpSbt+a+foUmDMTUid/WwMXCQUroeUrwulzK2gDEQqs
tEGtzxBldk6p11npt9cSBRB4UyOKmRNMyVlciKFRmKxkCvB4rH77e1vZBtRUqJIJ
NjNyK64oDzPEUXYm4zkyFJPNDiDv2hdYUZi29vt3+JMRyqn6GcwxQ7Gf+4Z7Y6mb
/j//ZRlULz+deW+Y2c9V+yVnf3EGbTvfoGPGzXLcsnNSKIuvco5qJp2LywFROTim
rKOrxPn7kQeJw20RJ3NmBwDzEuNHyuM2eKdY7oPBKUn2ce9a4KqJhjP29YzFHROz
gKst0iVTdJ1+92H9ZKH17rRsiMt25beFCqYjDflpkQT32xDR6+SYg+R9znLXXbwZ
6a9YbpNGBFSW4WuEg05h36UlgFB0rfmhsEqCl4o9h6c3ux55sWG07yz0mCK7OZLW
blrr11kLsGc86Am34Eor/4P8D2O/0vTB8btOuW0V4/sV5zp2I7u00MxbWZQfUVbl
hd+AEEo7JxcKJY8L15JYR7GA1JzSfLSk1R3LQ3/vWt8nSf2b6jeoHAo0TgubHm9E
HU95R0TPa4xVyRPfgwPOAP4V9xKSJrF520gw74/Y8gFdQOy0MnIlfnk9k4FmiYLH
s8eabuSaI2v3MD/UKgCwmJDtZNvz+JoqcLjy6wt1VSW/rMKc8wumh1RsFBEwYhXY
ANGi61tXE5YWoIjrmwh7d+Jz7X1XISRiRVu97+iNycS2bJgm0exUi+VJzgqhhJql
tWTp0H9miTm8W+JAyWLAeM8n1zXpEvtZX9RnejB2z+zKv/LzMVphiHZMLK83JxNw
T4JSDEmoAdXfEmIUbDomG3qChu1MNYeBeo0Gtf6b6TPrc3DQ2k387+NVJCpaNyoT
mzifQL2L/dUj9R2Jxhr1PTWQ5aMokXV+F2+Szxk1x3DZdwLlzwAFZKhwDqB1MGCB
UZ5y/03EUqDhJqih+1z7nAbUNr8YFDX2V5c5sdWF5vSBV1aXr68dCKwTqgY6U4w2
asrJLsjHQsoZcvMeG83Dm6p8KsncT90Wk5X0upmAFhkI1sUvLa8diHxpfkpnkRrP
lan3FIrKT37udcfIrKrWK2MUVVvKyWHpgpyWxdDQ6M/0JBN8dz/gcv6W4X2JG2uM
nmFFkuMTgIud5pbH076oU9R6TNVxujJrIT9gag7yLZ/aX2PfuY3FhhXBsSZc25v8
8Chxlp0Ry38wmDUH9T6sCH3ouA7EuhjMTtVYDS0j0PBeWqc1gx328wR58qb0a8Sv
v/Nir454cta/O7jndI7DW/aRuu+lH1DmSuBnLRLtZSJnG/nIxmSTAzxkyHdJ0+/z
743X72Aa7HaBkwQy/fSnfYICTZTBpOnVgPDg7YL1BsEV9IufyY8Kylc5w69yZE6b
wHhK6EpE0DFhsQdMZRDUHQ3sAMdpht9uKKofdWzwKKu+dmDmzs1FkajmCRkB6KJw
SabUUxcFKpIRbGWyTZF2sE8n4ebeez9ANUONvB750yYTll87pltemixw4HBOiECY
ypYhgXblZb1mcBQ/54c1q3/sNB8vkb6XfDWcIBe0doN7F4PE1k4XAs+HXMT3uFUl
SmYeo99G4rOwcqorR/gjLdWR6msSaN/Sn7J8uDA0OUidfcziERtOBPxNSfGXjheb
4x1dcK7TxBUfoGq+WKWHU9j4J7Ooxyduxyl3CDWuWF9d18HO6S75a++yhxISPgTa
z2twG4ZCOcLCuWOwamDxMKS/C9i2G5kfdiMHv4F3dyKey+aXIjPJcomd6DykAzHv
VLpCElRVn30yVoxN7pwodJqd2iLsrabQzSBjmriWORdCR0GFJiW/lpVF+4KjQ4X8
y28F2zFqWvPgA09JGPPPcyx+h0i4MH/qt1fL91Np0hXziuEIvYwNTY7OmV41xP6H
aSNhu1td8GPWHKHpAneyod+RCG/5WVI18UJnilNbK6MKO36RsLPhOMuI/nkdBjGr
XyqHyF8kO8i5+APiCvrQI8z0h/ya9ArTp71r67Nu/CWeXR28s1auXDPj01+Cgrrd
lxRmV2Ebhknuw5VRLQc4Pyy5a3ZEx/hoEwa1u8g2zHuxlBGnvDwWWp0NFyOHinPR
NW8a1HLcWCTW5v4qIWA1KTC7tnIJ6WQxW+hZr6UrIpDWz5ExCjbuDDhm5UUJml5H
FbhfJ5EnfuWs7YzEjvOxsF0xzlGgIB6dNrEtec/nFc/qVI0aClv+Jdle5WRqsEj6
cnhiE9su2ikZEgKVOElE71kwJe26GS+H7WXA0qG/ZQFDwYDsTe8uJxBq7TFf06hK
ZKGdZbmy+eyNIKUFL4ttevljS2dg5F63DIBaFRFBGIJ34S+KYrtnx8+dBsWhOvB/
PpVPzCyFSIiEdE5QCDMOcgLTmSRMxkNx9A44eOySDIKlM0j02voTZyXDZwOVtCPm
FMHBKWXtpi64c5FnglGySOfT8vxizREF2f7f/5LBD6WSC+11+OgUFxN1cp1d81Nq
q8CncTRLg7hN80CSdfJzxALjoD7ch/hj6ISZfdUl5LN68XU2xbLP3kEy4ROriYv+
DjTR4oBnGinfCzlWahesvXtqG9UL1S9VFfuwqrtoSn/NmpHKciL2fzSF5pc5MDWC
AkLrd/abie20lKhFJ4+pN8ha+X9Fft5c224Jfh7Mny1YadoJwH6xbUK8gwNJjRgw
1Yvec2cxM0w+JeABNPLL8NqKSqVyfe1RQLLF6eCUbePgetNi17pd2nWrB5kNLaFv
4niY45viFJdoSH6VwUNNmK6vglGZmpe1by8o9InVPWPDyClSwAHpWVU8q1HRvCru
4p6P8G854gFrLnLxuLIXAoVpl2HWVJaiPg+jD5UemMGwJs4iqknRd+yUzGFV0Hap
LggQUmzihEC2tzRYABtfX9iY9g5r+Asp2kd26xEWnPwQb0SzTowgvuXuQjxm5VOi
rYQA4eMzgBt1KaRpnK1q/tOqnGlsg6LcGl/zeCTGEUYlHkVegQxPrbnlmDg0F6/B
7ZGV63kU6o/x5kbN1ytw16xpwuZiZuIi6a6NZC6X2hf7BOHuwKm29zBq6rR0Q267
mCMPZFb1OhZVFJ4zsm8mVTUs8rIHAgDXfbl1z7KmgziR6JN2sXijejyU0WJDoqj8
q7riHUnaNkRwcbQqiMvQ4cr2YYohSSHxmoKXwoe4fVprwP7Yt/SIaWPgYenBN71o
85sHmxCNfOphmzxRE0EyHAWiyVWDhhgjBoyu/lPCVBTyqw006ZZ77qlGkth4a11y
NW0F4WSgKLC2Dbcs5ZBJ3B/gLt4nE3EpDvo7JtFmDVdHL93MesyD6+9F3cytXp7p
2lUusfvAK0bVCaSvTkPgduknbtEVtdNqWiTuYw2p+40zwuDSSW9iw6v0HReFajGn
/Rqy9In1qpDMhu1xW/D/5NGNCbOC0TzCqcJGUjdDPeYlquAvwHOdODj9QzsWvbgU
b6DN4pX/DKK4ktm8naHNSOQWmlALThZyiYg372k4ZawoQOIGsFQGeL7Yxe+tLRVJ
B/VzM9S3KocP0n84e4nEIvnWVofDX51ln7c8b6tbNzPu68CecB7rzyk191c6UJID
1PP2itWLONd9fWg28csbzR1intSwsOMmEi0DQmolEX7Ql9ROBFwTJAd9BSrKbJHU
f6Iijx3iAiTPgwOP/WGdlUzxYZFu6rpc/PAAiPDDMg/oPhUfRKDNyGvjEplpweP+
an4tza1fAdleyFn0rC0YT2YV8oItDEcXjXYguWrwg7kIvrBoA0L53oNlb/bEln/H
rGfR1f/1priotyYuKcLjJZaLEJDQqPnUtcCqkjOQvpi3Z5113gPWHIZxaNHWW+2A
MvMIG6NDy0rCynxSRGgKmpPSGy6r9vzT/5OD9c8TNjUyHZF1DyaJIS9P1FU2DwVk
JhCpJGKwSsJE/pg7VJ1mr8YAT1l1J+KtaMZXk85fVooclxElemBHhBtzyUkRCN9K
LgdYo8mUeJ/iKQZ2mqw+02icYNVAxe3zJ0E6ECEV6dNTmn8IkL/BS8OwDWBLWzoW
matDWiM+ljc8ECF6ER9+g1/0zu8se/pZnwfSvLAU8rQTNF1NvAc5W/162ilh2eam
/LWhJlgQ1EgdOWflVD9UvR2w/zVD5r9SP0oAzQx2HXMfdL4RtWCQHS5VUT+Vc+rw
Pvit0i/Jjaf4Mun/dbp35fcEpL8Sq9J427dpqQDsTZRmGj1e5PpXiZSgT/pqWp4i
HCnXQa3SO7GNv54vkVKUDTqJjyNGgwQh7LKCeoICC/fld11WUDaYBm77/7w91NRu
k0rD1Vk5qaW5E6vo3tk+ZFGOdrrRYERwUnMg4FEwazYziikLW3tleGMH1JJChT74
krrVIkEu4k7e5mYSj+kjDyJl0tjm85oKQ43aeH9GQEHgVNGVbrw36hB9vMJy2HmL
7jt9Itfu2DPmjE5MxRbJj3JzSQhx3bwEDg6V8FgzXE3HIboKxWzQMQ6xlNeFwdaX
+CJutA6/TzzT9PDa5jVan0mB1SEwPJN+srQYAYZdjumgtbITQN7CsjsBXBbc1wNh
Q6CvXom+AHmzdU0cXCGX5DpudXRal8G5fjitCYdGhT2D0noHwyIvlcTpH+72m9L1
UMpzjC/wWpdInnaxAqXJj+DpY/YILoDHqRvGEp0J0rUGVVWUK8YOlXsC4BidVrGK
0rvBDS7II5VnaGGyUdM0gUqIA1A+2r7+ENe2JTPK/yP4kq3xPflNH6Z3angFlm8u
m6WhJKNUF6h7W1HZx0BEWLFD13C2dd2VTE/fbk6T2eF6wxB1Ip88Oq7bHDXiNDzJ
o0Dont+kw4e25fUHDwnfMDsH9jk61tD6x1KB6MfSsJ60aQvPpz0i0WogLN5t1eGL
m/VLBgSuOntgLNoByeU6jv9lTui3W9FnoJta28GF7a1+hTDQgmXQar/XD+UP2RfU
thTy6JVwz/kT/4nAtdAuMjQgkgbKA7WL1xXeDZdYL2u1QxS58S7HvAaDesbxZAKF
DSpDiuJnadfI7OtlZGHLtVuaI/eXlX2YvYBr86l8+MN0CCAEkk3iYpczpXBu3C7T
o2leW4CsDbOLltZtgotgRUKoUAkb8KFMgACanNgEikoz/VJwCILua+mleBrgVbwv
IqNhpr1rnYkHDUXVqMDiuWDgL3q7M6BNV4xKZ+VhoRaDxT99p9aOTrVNYb2kGf7w
r5SKYZszj95NLdAFnS3Xs+fmvLski/r7G67YGyJ+tBBLC8KBFBJYdXxjH3Nj97Oa
iGHnab04I7gSn8WWD8Ma6kM+rODtkWFNrGXvDheSpYT2pcbO4XXvj8S/ZGyTVsMK
l/Kwic3ROXs8xQE5By7oAbRs0LeyenDgmB67ZqFpWIaUxPZQgS4lvzuRXLduDjMY
C5H85H/5ijh9MZOfRqmkUZxcwYZUENdO4tLmpbfjdwOuakNtRxUCXGFxfr1Y4zUV
OwDhJh5urZUsQANVdUI2tltCtTJRvR1zhSBebyjHrWxtWF2Yewwi95XYP4MFpPCn
pI00KlpmcyGQ3qx0vUmTKi572qwmDgLhHfWKnYvv3ZwH5M7osZIpV4tCInIXvj61
z4XEvrvk2s9as1i+8sK0lZsmflgv327325GlYajqp/VUQFDvEOU/r+1DiFm1tKoz
EcIncM2Ry9CyLiLflcWnsrEQcYD8Kti5qXGceH9CE17xiRlTKx4VKLI05iW9KzYR
YB3yJ1VfkS8g4AfcgFscZDFABgtJADqf5vAS2UeSRwg4caNtDKk3EISvl/QV0Ygt
28UdI3YHH5/TEsT7EeRGjVsQhdMYxhtR0jO/grYuiINk94JSjO8eYqCSkhZpUAkb
C06ZclP8K+KS41E5A8Qg3dwymxrQkXudzqOdTY7bU7AgFTp51zR3yPeGMz5FE/4q
tzHRmuZCsVTQv3ZCyZRSsb4UtMeI29eaa/fd+26Fuv5qd80bRKEsGzg9l08Hiox8
Rm6g9Kb/4XB0j6Pc+wDIZ3bM1P1j7Zt6QFp5IaTUej29RRwdNwJu5bW9pFNonY08
qQUCk9RLUMEPnxnQYx5llWlzGJ/K8Q1bIEA0WGk/KYUMlJWbumt+LDVtIAg+Pezt
NPT0lx2XyQCCPYasjAiDjqtB1Du13CbkcYgEcuYzoFCB1ewM7uAQ1i2dNNeagWb9
LXkVA3eqxBx3KUUVrO/X8xhceMMhGYarbYvU2QIV+/CV3nvLvHd50J4WFi7Nboc0
22ejoaY7lYwsew6x1VSHzKMcpFy7dOnLr8uZq2K0KgbX0g9ujopy7vWOKtW8Usqa
fA/AoaqcN77PhAKqQiRgzEX4Lf7pRvNS94HWq5/tMTGLRf7V5rQ/Kyup5nhhDg4I
mdaBjNxE7u/xgQ9T+WuqWXohBOPgYoLAIK6WPE85wf0RXnAoJlARU6rQqcA86z2C
xeRCD2EOd9nnGQ/cCblhdk0ox3mYISIoCxzCk+XfIbtAvx1MR7rQ+yQvD6bHjj5N
Z9Xy4FYfwp0Cm2RcegQlCyC22gtAJEJFiE4hVvmLZXqc77TUOG6WifAMOi9MhLZk
ST1OGsrFeV7+k0VUfIXMp0a9654BcZ51U9qKUUGeXJNmUurlS3CCE6KgfanZUvCv
yA+ti5ere3yfbuqUj+Gpin1F9kIY3366O/dKhA+vuovGg1S3NmRKjlyX+chzBQgQ
Vi8ruR2SkapoBfSd2nRA6jXWgM7TPoYGQ0SrHkXuKLS4TadPrT/6oJ77wRG3GC1O
I/37wCaa2xI5aPFW2uqTDqP0KGtTd6zedpw5PoeTeX4VSzeH7zepusV05Yo32rlB
Zc1lcQ5CIfbTU5AMVuBupRkqVfQTBWAekB8o2ALKGTrBMxVgIJHBp7Sw6KXgw5bH
2ubKWXw78lyOouJXc2Il3edDoZJog5bU81MtMuLotQ9y4ggbgFR6nvR2RMdOuqTb
G+J95t3IbL0W3vO7fUvrFnQBYV5txO54xDelz+va833E7gw/cPgMW3rBAxTMW8NU
efmOa+aSthtdVB0b4XEqoFAtb0Q9rGpLRZ08ylEW60pcjeo+qSdbTs0MiDfxNSM9
h4n32OK73c3Qi66mIIz6Nyo/UMV+Daauk3CsuE+IqNKpHmTJVgvraEDcJpUhauZp
Rqx39F9PfaKXa89ow0YhehscQ9B4UVvu1g2W7QMewSt1K5Pekqma1RfMzJB4caQv
GnzkWU9XFBWq614zRS7S3T4qS6ncq+AnFIwNJEFJotU0mfU/TxeScnEX3ruTQzW9
XuCABIiKkFreWM+pvJ56/HYU8Zx4plBhbyDFoCJfqehEdspH2eXU4jnCXTcyt3yQ
yhfruasaHzZzx69zBstksK8zs7N2DeE+h6kpxAg0z+qlsljeQCpE7A04VXYZ+lGP
45wnnQlq1/aMde1x54VTP6JGKXALYHItTByoaYUh6Y7YkexOADTcLtiVt5voE+OY
ww9TrOOTZ5iJWy/xC1ZQ+Inj2Jm5SxGMOCykRz9n1GB22B2aieBDHc5xcBiyACm+
Ikh1r1qOVHbHMyv/u/zGL0uf7hFOhxcNNw80KL1G367Cv/TFo1dcOwih8YUC0AWu
5aVuzh40hIoB4Uh7yjQeL9cKqpLzjtR5/aS8827UYw8c+y0lhcl4lxt0mCypx+J6
neF5YM8KW92CCEjZuODgGExBJWDhSHWLJyDjaFnicfcSiXEI2d2y5q+OvDfCSGBW
wYjTwOMTeqM9/fDYgXss9/gohSYte8ZF7IMVDbPKuDGGi7w+nJRkX0xrDsZcS34k
A6/Z1dJRZFXldPyHy/lGc1tizSoySP+a2+kjX/ZjDj551HB2stUv19fdZDbwpD6/
kkVrtTpLM9jC3aKdZdJlQcJk7NLOhVvZkuuaqvVEdl5VcapnNh2+CClVl3cFwjh6
BNtBJfULyWVGX16z/vhVVo7O+UzOuTDs5NS7b2Ekr9mOQx+Uz5ii/X41ev4ArYTZ
1+ky/Efsx/NrGQ+kEsArr5dhplDUZf7IEQXSQoXORCmbvueZEfpTgQhWN67sn5iZ
+uDQ9CQG3B+ZsE/xqVAvYOlA5b1N9jZGAfiX61wYszEZv1FvJFGEG++9+J07vrre
Okug0WjQqMkkfeGTrNm0ySUNdINz2VMAJgkr9t7+MzPUl2yNl9ImNKDSzOjIhbII
JbFykzjYrTdTNxADVHXiTkCO01C6w2/0nOomdUN2XXW3p6eAXguFtC/qcnLGu8AO
MWCO9p6wOcOCitxalj5XmlTEB5NI125lctY8ZJ5VVLNjogWcghaJfCHT6aCM8OJs
+4iiboKqdsQgchhhCryBTdfObWxxc8dH7wpGfYnQ3jUK2emR/kzBK546wXz/yZcx
g94w7ezR74Tm+FcOdHwM7EMPOnyT6lOg0bGobgSfUu3tcy1q5qNw/lbOsV0fLlPM
4F+rTJuhW5isWzSuO48Z+OqzSBBSItnjlTAolB0RC9J9a8hDrmTQ2H/ybft36mGf
FUO80C5Tcs2lwS1vjHGg3NOfRFCZ2DqhB0XmJITqtWrRbAqezqC6mwOogj8S3m1r
RDZ+b9Or59OdYFwC6ZHipdG03JXTTOxWh8zmrisyxr6TtVs3yxp573bl3SdrINVj
LQf9YZ5KJUzSGiE7fY0NIQ2cX/AX1dJMHlatj2yoL02APns8YD5rsJpVX79KVLN3
HXK+q7qdvLTU/wQTf77yGWgzCcWmeDm/18PLGHVbTU0UxrQ3fn/ClDnQ48IYw7rK
fRPlZGy+W+jpBBKqWC61a5/G9MAxwgXmVenf5ydZQtX0Gx20nz8j86i0mrRu12kk
eM+JaWGmBjaGrlIaI97Al9LJPgDvvOnVm22hewhQmRqFYuTR++lmU/regBKnZMBZ
TTgS94qc4/UhQFcBwMweOY+W1J5SuSTJ8nds9jKxCGL4oXjbvhIAobycuSc8iMf1
53xnBJ1gqXnMc2SM8r282WBPdkJxtUTtg0dwGp5CxOwPBu5Gfja1PGQmDrqfvvUE
jmsyc+WsvUzWbkIlaF0EmbpuYSS1C6EA7T95gqgHvxNgqkMM2miTNH6u9ckUkW0y
t9v/iIFGE/7/ql5aF2Ng99LwZWfeE9Ta1O28Vnlbf/5+Clpdwgg78op1pZbdAzc5
bHWzClXugDy7UPlxVxHAkB9cA0e9c7WFk1KHO8dll107TYyfsYamhVGdCY5re1Ag
31hBAqSAR0KjCEMUoy27/5YQAP6YCKNKVWNqztqvoKp0r2XmemgJK1BryL0Vk++x
9E9VA0tTvSGpgqrE9b/JvMMe1D6TZ5Ya4SG+8D76udZ2P2ce7gYzwB3TZn8crqNj
kWdKDopEnlXR8/+y+fWW8N02NLniZz82EFB5dUqDGNafz+dgcQMRo5YpMAH8fFSW
QlKLObu4sgR/Ki1VRiM9dLWSKeiwYtNHFG5fVLKNASOhnULlnSwCyfgN5gKa8iAe
lXjMzDqq1YJ491WuNvdZS3fBEclJQFU5VvvZyVRcgSihN0ab00f9+vAbuP+hTC/O
VE5XRnYQddGJTc8WfZK3Lb7Z3104MBP1mzCC6nvyGjpmbxE3Da3ft1T0/fbIy6/Z
T6D0KOQ8Tu9BDAyBpVKUyrBKfoboDzYDqR1lcLSprrWAzA9A8HOmfYtj8nSf5Qym
2ke93hwb3ivqIsik8shqJijeRkQMHLP0y1A4oyuhQhFURWuQXX9cPXULdvKw18wJ
RJC8eBpVsVAvGRJpjT5EF/VAkW+i2WRNw+Z7m9FCYJLVdO/1gfsrnx1LiDP/NQ2l
/80WJPF7senFpXv0iT2gmLmLDPDDbahjjAOpUQZStqupkagGmGqiWF6pTyxZMsfG
9DKvMFJbF5QVJSvNcubRSYkftYdaiWDZ9VGA9cNE3jId/zc2LtomVyfALYAMl1HF
tTdWu1TxxqGwq2mdta/lAfaNWR12v6ziHWf8HLW2Nfzo4xtiieQQTT+/07EbHRPK
4d7y4XVxtH+SJl6RdowuxTAZaQDYNQoMLnxFAl+bqOPa0434IJiYTo+H7LQ8NYBk
1RHkybGfHZev4yt2m1Yv61UaLbMbZ9zo/5wD12G8QmP3QEommWNJo+TVr+0qj5hZ
fPNh/SsyF9y9YITBFOl4AzaybhJzqvRjwVupQyvDEiSxu++xYspBIvsIdctJx4RK
OOaMV6iglMx1Z6UW4ksSaK2qI5RPYS6RnNJoPyTslmRVQ1wcKPGwt7MUf4q+vilr
SBpjRGJmkDbFXd6d0YXDUw5hMgGvAYaT8MVT21LoY+Bkg+r4aRMLL+YxJVImTd2M
3lEJmdEuf7QkP+mVUSwhtOsEHgq2bQaqt9imA0gg81NYqWcJjTXD8tcnnKjsiP4G
GqbrtzNPwcs1DNbnh3fPe3qShrf8gb19xYeGH6pCAC84FTxStTMqLcTu94vcYvzS
UcbxLm0H/gKopACLa/zKus+ELvHlitcjmSMASzb3anKF298pWXFITWPkJfzO+KjD
pA/qa1an0CVIDMPwCsKZGy3H8hLv7dS0QxPaS5pAtNb4XUetYhblzOL55BLcvetc
bGyOo/9xFXrficOCg5tHXayYdePU989+aJSwOZH+XTg6vzmttKhBno3HldfTM4N0
zu/Dm4wnXKCEzkYr3c/ADrU/mUADtHr6OVcYhKED3crfeeOfUbNGVjzNiG4C/k40
5xh7EXGyfkCaG72eDm4kwMczd5WC95Ti9OihVlQ78s8LedXh26BJffXvIEzXP5zr
E0nRTgs9cZJ6cjhtdrnfmkUZgHgo85jAfcHy55055GdPNfNH7QKAeAMZcLFn03lC
0c3DaCZH/fSYYIppAYJ7GASjbW+S8yj/FTRizZPS/lP0TZrclQwzcjfqJwSrgnWc
rn/PV0CjCRc+/nnxdOSajzBjT+fC1BE+KhqXhkVGGlV8O/qfhBHgZ9RtdyCbLrg+
7xEmsc7KNXNBvQagokaGehCXUhlLTLlQgtojR1y0CXgSYnaFyub/YPmzLISAl551
6j7m5uPOtgrp9/6G8ewkXDCUvX1whj02beUY+lpCIpCh5/YdgC4lD+8xkXr6bsaR
u9kMZvikKDtpln4qIC5Hxf0Cu+r8ipSmWThIe4qDtNqw+/PW2YHmvw5Ax6VFzGQK
HKSrAkw+e6jiEI2t7toQcp/HqaV4vtThYRpWyXri8UJEjQ9+/V96QEqh67ailzuV
/jZBXsjPmGeThp19oYmNdVDoQxxRWeSZin/LBSvYeIacmesF5yTdoi1VANkVRf3N
JoIiCjKz9BJ5o2elaeo+YD//LF5m0G9d1DetCLpJ19alZCPhtRgkVxVLY0fNhDhD
qsT51BHI4a+FFPJ7dkLLuAnodcL+3UphIu3+BNJAVJ311Zkik/fQ+WV/BU/+gUnu
AY+1BOWcJNvuyQTDRFhkYvgYzhTvxsnTDXlkNDv43GgY5WxZbyZfokdVqiHZNhnt
zlE21zzSQ3KkZgbl+TMxXCRZONI6HUPoBOiXIOmd7KlhGj6seVZKDfKyDRmPfCPo
GO1yHPmtevt3IJUl5xLq/Mgv64lgaed4w+hmmZj4XKq3VI9Xcm8RVrDB0tMmv9O/
qKj41Cn46hA2LRrHR5LUAYmTjU3a3FuwdzeASDZ2jFDFas2XKQ62MHSTigIu5pMH
63sCOq6vUiAkLjUUPYcLxASYw2C7WlFjbmSssXpXbIWnbXuJKMkbW3bFqr0PPHu/
Q/V4iTXFmUIu3VpoPZR52oWrSr/LJm8g4by3INWAo+hTaH3NxTG/ASY+8TLkhjM8
qM/8xirS+ui0OUdtcrvrwo/fDP/YM+wwTRqU+8qkvg4nes091Y6N0GEJbTJNwH/H
2TQJcuHCFCrCzVaaKHPcCL+4CKBWXOGi9WNnZdrA6fDZF4hyvERFtTIP8b7XR0qA
Il7G+KrgqqcKmlmJFA4BzKkr/1qhGWCsYHG9EYaGswHkisBQP+X1krzFUK3UG9yh
rSbr5/ETI/vv48LsdhERi9qFLOdgfj1PPNjC+vUBRTGmxIkEF9LJrB+cSweqe4AJ
z8N9/J96JY11BYkZg+iVk50YNnx8nXmyFwd03ZcR+Y7aItHgoSbvedcGQBFlZiSo
OyfMG/05FGDC3awRmFQA6959+mGeivWItE/eoubcK9KUQpzfotFQqX+0DzED/EDF
ae1cIQ4NvklZJpWbszfdfNlAyNI+D5Z8l9qXhiQeqzpxmBI0ZcPWMZ2icp99rnqO
4zkCuyDyYpxJT3FzrI58ABYkcZ8BPe4NCSD5sq+H2qJKbOrdeeQihcjXYWqU6Los
jtWpDzUzWMAIdUs3KzQUuaaaMF2Za0JlOcx26r+6pnIfR8mL6QS3UhWfocSvb3+Y
nEWD6wEbh/1YL/E78R4G6LE68WMfHBD4eAURRWJFb1BAIyB+ahchwuYrY3/XkdLQ
PPPpydPwAJVPbZAuQvYhaIP51nYDrcJrfY1dfhKi7ELFW9mUqOeVR/Tx3gLm+IUu
0lqDR1EMHlRyevTxr0OnqjA6bKre9mxO2iv1ucLtDJFpO8YJLn5T4j614dxDTiB4
DHLfD5cOMjjRAKF5TeOl5clifX5n3LQrjxfZFZ2bXr0JTzsUL/1dfZRCpFGqavc9
Ri/AZPHOZyQ0ytf9HR2eRQMBFRK7dFMagfWEYKHxSQx0ErmpHuZvF74Ma+Gsaz9d
J1YdSqGGpGj9FW9vEjRTB5izfs6HHFunH2jtImeUI0gnKd0gu2N5Klnj5zCcn/r9
XTXbFso5EIMA63eytMpTubkxxSFjIzVjPMbD4raUEhOw3y/xrHXhtBY4Vy288bBm
KqwriieqqEKOFen80JG1c9kSD/ZZ/gPzjUem5RN7Sr7ILxtzX6XOooIq0B8AtaqU
Xdyh/r8iQzrNp4kmIcMNF3GIumNwziAHVp0YvzHPf5defTyC7EMWyLdfB1NNI72j
em8DpOxG1XZIKkOuQWC5lVhL0zwR9K1zpV/GD5hA0uy2R3MtFKTS3knrqwgTencZ
GXnlJXA1kNaQDsEpl+BrK1lMORzgSW5rdI+kWYyDRclNoLtn1nscxyg6yM8qUoTa
4JSF2my00fkTIQr069LHGguyTQcgqTG9n45rq2bjV1G6+xk6nRo9DEi/NnC7RiCr
pUgVe3uzYiARrKaaabQpYK4SleQQPCvCwjDb2bgFMqFfbhE1Z6wuaBpsphFAQZ6U
xyQvS50LrcfP4ZlQjJ30HBVB0YcGVhvSZIGyizea0zBnfzYwsvlR6CmWkZIQmVGB
wSB+WTmL7LhGj0/uzgI9Mb7nguBtf3A/4dUB7JDucHI82MVtmFGYXf8ZAXiNLEcS
zyT4sO8MQsAveYGI48Hx0Sc5YE2KWr4wcBxw6ct5EVmKjMDev8qk3T2DUH/y/1Ot
kVBOL7vL/Ncr+OKpK6xqgpE/bN+uRN1l8VDDwCSDQIaZKvJe6fUTl5bN93ArpiJg
th4pKS0xcFIttLEoSlRaIVDksj7JQaSa7eR1tGIc2AQxIrO8/hJB+sn7veB4qvQk
VUAbDXswG2XP4m695bX4nL2zEanis6ZUhs7/uA2XbY5GCYD2VE/aAb1i8P7Sgk1z
ZBQB03NRnevhe0FweWt57ZBxfpdrlh0RMInnAIN4953xKLMIJI6AjMpC+/TGFVsU
xa2Rf0mIaQR4OgXa5NHTKhmXbjykMwfpdugygpZHUTrv2Kxy2UnVrp+nZGBM65Hw
okRQNqstwhEog3r+wSX6bXM42HyhgPv3kTPThdHx9Ju42yeyeFQZ639u8l+CDdCy
UzRXCfYf9zFAwjxtogaY+cJsv8eyerbK4Qu9VpE0vUjssjI04djSeuSgGVA2Lp+V
giRboHIodf1yCUW5eMrGPq9uYgIg56W1+MN++Jfw/MwIIGOd1btbw8aVn3VtLJk+
+GDZkvd/X9Kiq5zfLFvHZ2bhKdE5JrCEAbvhlA/zqvCNB9gaXH/Yaa7K+JD/1l8B
9CN1lpARal9TtF2YQoODbrCwLP6iboo7QwEsOdMIcXkUzguJkk0ZFHcUTBqvVYEz
QpMkWcRHYW0PFku4WAAVaNquX0KeiWF0QI2L+FCafR2aflDSfhOo6ySbCc9qSwrl
P03+cJz/+GUOdpS15Pv56RC730/QPLPY33V+Tl8aPMwCVOz86EtM3w09sKaKvvf9
JdI12x9b74j0g2hXsdD6GevjjHjW2RBbFJrWXUjkmDMdyt+ExTvfDzBvsV/JLXBf
cDeFldPOmDJf1cAMpDGBiSa3xA+LaFqzBIGjbUwFoZfxmQ+fITrQRNcuQde+MgUn
xX8G6seXNX6vSEUYrRfqw2FWZaQ9TPd4mgpAf4owGQ0s9yVCE4U+v/o8655Kro18
+XMuDWAT4l7PovJf5Xbk4oBXZj4UXi6LIUFhTRPp+aB3pzgXzqGUpTJDiB5nS7Vm
wtV0ErcvP/q8SLs3E22NUnZyUQ/ON/aHUiHGZqY8Z3o0JOxcmXov9wiFR8ZYTDBL
3fQcSfw/aYMLn+wLba1K0RgrUdWwOPcj8HvNciVeCud492ARO6NGhpfE1TB6tqO6
eAMTUIDCZIB2fV957df+Yqolib2BuOAAtBF5xzxVYBR40Bvlg4tZ8FJdPIdhUrFq
+4GMEAhwkLiBIAlxKzD0LGPYasZNf+O+TancY85AEQsygs8FRldyN+//XFyt192f
DedazHVvrXvmryQd8k/dXBM1EHoxM9uAQcpC1YU3yrRH4ux/qUvhQgNvaznVZTz7
bZcY78VldMeEtNqeirxYvO+OAyoyS/PSB4OIUkcYQdoHnw8Eljg1E+0EeOrW2QYI
S3TiADJaspoNaSkszf+jgqIotvFfD8inas8mqaOjTgz8rDPkxiu9/B7b454AsFJ/
ZRMPVFMPRf8AvadOp67uaPSdMJddp/C0slle3wp2+Dpx0VxSBnIsS0qqcNQbswED
++oGpjnbD67cH4IHQ5ittVkkjUUMny87CLG6y2S41DKGtz9Rwrh/38DmSmu8oHdQ
QboH2SnkqWIl7Kpq5xgol1La0IKwJJqQaQs39wkiYbNvFRS6eB1xtDAIqAFpR2xe
POvlSUExk4GSxb5U+164MMLj4bnKFcgDCC9D0+f/NJR3amu6Bn4Vg+mJwXCH0vCL
NTRFJYwYT8L6IXRQWXsVdbomMAyDMV78/JC3exXuUFBSXU5sY25NO84iCj9SP8Js
8bpwL4gvsqQ8WcP+aEgQ5JS5fiVfoI/T7yxOpmA9dv64VOzonacBAQselZ2EWbuG
rtfLH2WdMEGzsIo+o/kY1KBB5tf/9zMGvNBJReDRxmNcs8jWiFs5dOOnQ3NiUuIT
Us/2CkdsVJHbTlzAvKl6iSG/+w5/3tTCrJkGVSjwwHUjN3jn2CGqJJO6VZziPrvR
l21gJUu0bpZc5IaEEN6pPW5MZrrnzTLItmG5k0vS2N85hRcZ5ixZzGojutNPEVuf
UM3j7SRKD6JVY/AlKj1BXul925eSUJJm7CLZphUEiizywNGYYuTNJVM0GqQG45r1
fOVCUHauDK4AaMhtppyTik36GqIW7LPZbTDM9uVBg3OyUZoxzo13a0vCiDiQXJoz
qSH28IBMtLhqloyrdiaEv/C/++l8YWXypDVJWTgx2W4P/HsV2iZV3FpiMaafKtiD
o7ZYcDluv2tChzw5QkkkcVNfO2NQXWN8lTsiVIUPhi1QwKLBsxr/HjuyfPzqYnYd
lb5311pfIYxmoaf9B35y3uuFtWxCRLKgGUw4Chsuy2yGORA4kxviBFVrNVg1TFCs
8Cds7FF6WojuXiN2b4kV/cB6Ta4qfm6MIVRJ0U6VVSYGjJdtC8Mi2e8OUdjS8I4I
3WZAI1ilFO3z5ZtqCXma175VEyzYj+vQx6VpJ4OazwrbL+7ZtujcpgAVLrpLd+zx
mJLBpl725H6+r/QrWRqz5uN6ZvxUAoG2TFTnw/GVy2gM6BLO1fxxGxu47kI8xDfH
RO8IVtxqNE5OC5Hl6rm0BjJjBfoG5PG2d1AN0aa+o16zM3tWKKap+mds66ruY7B9
zO4hnsGtu17VIQ9T6bSzk6AL1KtvIwvDKk/mYYuBAPGqx5WJzla6nzI+ORMtNf79
L79oM6WzuGCYnoke/DSjYPvofzY3FnLmYZh09eorLBLXaGaCxN2eq76LV0k/mF18
pQYhI/KP+FBI/pUtmRwfJ4D6NJLBJpslKHOX389LafCnujMdQRS/srkKkjgPe9Kb
tjFdHo0efMytJ7nVWKFpuxZnZ9/l+yOb/dLvjlURcmBUGnNTOJnEbzWbGGsL+gGy
yrsFtUecXqDLXghb5LjcJia/nr8Ds355rifDuv3w0M0n4YDKMaJpNy6TkUMpPrDQ
dikboFSZBLhhe4SxP0RtiXxitCzJXwa7ZIHWB+HSuhpqdSv7u8+VnNG5KWbfm4Ff
97AxjqJQiL0V2sx2cJzuz0toDv3eHqY1nKG7XOsKnubXuE5k7o9dbceq7mmeBPGN
rdoZzPtuC1nhADYqpjSmo+mRGScBezGJ6BfaKrzVIJ/PWQM1L6dbszerA5S2DUie
Oklc8CrHNtwZivEBzy+dKAOf+PHbfwRiHZcCxgrIYa3uIjmwLNNyl1BRDAE212F4
WgxDSgutZP0NvfE6MGmircrpuxC0yjgitJ0k/JiqKM925YTib5zvti+vdxbvqUxM
k8NPIKFYGyQuI5PXkDYhimFyf7vUWgcQwVSp0H2gutBSLq3kiGFNh120fWHIf+35
QoOGc+c4WHMoJ7KH4WluEBd0KsfM9u270ZWLZSl2R1j12gtGGKESH/KX8Defj7AJ
gLeHiqp1iiuOvpdYFhrLduIT1ATNZmIWj9onGRf7cfPNfLYdfj6uE21ak+xQBBk0
bsLdaMzCbIUMtPypo5a0AF7cjMnhIW+XQ3EOrUdeF+AGcI1LjMoycbaDSZxdLVFy
77SRDaPSKq2hDAWVjpIwkJNHhbS086z7JM/6KXSQqsCZ/BgtZ6QihAk8vbSuIqTu
ohECjwao0di9CXTu6rWQTH6mZ5f3Zf1RpshEICxIi/IHO837DmTqFX5dk13mazN/
/xalV88rjLqhx4FiO7OHepAnDLV0sXXtfsNLcrLXykqfjuGlTabmuDgAdRL2tnM3
8Vr1504Rn1Zd9nqbbs/C9ViHOUnichBbmZXk0lMFJ9QRRWdr4HunvMtSYLRNsFCq
sxc9XXnaBkWE7yz+UzXbV/E9t7HCp+GUsPYtdztODstwlNMdHTs1scLU2BS76lFK
vhkQ+TUOkj/HWkljHyiBE6KeD7sCTzE6aUAwWktJkXlpdELAUILQYJbKiGsr/uTr
NcA6BJHOi7V2RGyXYfDGKGqvwluZ15n/yAAgvyaTe+iAVHC4ajW/zyrcT54q2IpM
vU1N8eTuWezDn0hBSMy4iUqjKSXuKx1M6bcWtPB2LSTiqw2rQElqwWzP+LGg6bAm
vZuZpOn0WFahxRR+qpKkIMun2k7lCKvX0fM0nsiyTNj1P7HmXoAMJvUqKIBdYPZk
XMLskAo6QKaTW+cejEnfXzTXv98gSWRq560zjHoplE7IIgutWyzZGl7kR8BVTv7w
2/rnpobDN7WS3JDyGoLdwJ+lFxuVqPzPjKLMbQJdXwEX4sTF25CM7YerKwq/yRQ9
rIRmFNuPW3/jqSUdjF4v3rAdX+UBBB/sa/OR2qsBoqiB6DzC/Z5WpaiuKPKsrA0c
syM/eUA7/kb+99NqHtQhUohH3gRaomBCv/aevfTehVgkYbhwgIe7PRVzvaY5QKib
VGJ6A7q48BSHUIVo7LnjjR8v14e7t8ccxxn9wRH7wD29HQooRWnD+4i4varEuFMB
s8JKBS3G6OklzidQR0uome71xo7KFLx760W8T+8H7PlWd3ssunQmfeOnbUWbTgJQ
iiiBbnMNNUBGzzClls9erbo1IAJCp+u4fmG40FcDsNJm8X3k30LQlg/Pgsk84hxB
57iHU4xXUjwqDpmHx9r1GTyKjL8eLGmjn/EYo8IKkd1NVuNOyg/hDBd8w365S4bn
jJAyfCxEj7S2qB/oYqqrB89RYhlbbv8YRBkKyLuul/3K9vEyPWHJutGR0lpnnvuq
cyxkkYgkUH49TVo0DHIsFdhbY9y3Wkq9bKbY2walXaQneBVOxHiuWI2GcljMzcZ2
vQpHY9+UOWNCj3CTqjcVKX0Q6cdiIrlv58cs7UH/GpIcNOyDJfFer5X2O1p8s2Bk
AfcLY/lK3KDoL9+s+qrI/6Z57X1bKELMzkCRkiqghErezx1abzs7YKvV8+eHpsIK
Ax9MZb8HT8TMyCA+WtOEW5YIZreU3NjNcyEKe4sZZHESavjD3KgZGq/hN2zm0eKo
nKxWkbWjqbxb71870kXP4hNjFSKg/SyErSzQFt3+BOsNFkrPCQpqu+GA6kvayslW
hbam0TwbvEGcJdR+g7XewZANK63h+XGjK3rwoTFBhD21Sap9uvYOYJwN3KuObyCu
+BrYAgCum4UjdmlwyIYy/ZxyLuzACFhrZODZ25WxEX+YrN4G6MtgjggmfRlbQ6bN
ZoLYE2oJ34V9dLJh7cdlnKvtdrV7sCgDYC63DSAN3BXf6mGD6XGRM0K8OmpTaO/e
sHvU9TSePZ+NWbEHCtR6xjRO1eaNYzgC2OMZ/UJAcY0weIqfrPJtO6MaBuv83Lay
jXcfBT+IGRoUg65osMa8LLQ6jcAgnZYjBHB5ajO6LOvXiPwUsnzfzXUELRbYNVlq
sBJh7BmQWzM0YHMuvGganFGzB4KdjGgDiphSRUmqhRDhZ6H9qkRsLD2qz9B3/0hX
UWuuQM1ounZZxG3jJhANEMRD4aoMHyl0kOuzAf0iF3daraHqYGLsj6SS4BYUEQ1W
P6/eJB0jc3ETghIWR6537IsPNfgsfjDBN7WUQED3gMChTFs3U1o+m9/FIxdDZYBC
5PLUfk3BAk9hP6KEpp9y82Vy/33pJenH7+Y0FzGgqyTm/ljVMr7AipFvzetj4gIB
pp0wnm81y2rLupRYbQGDlXp35fy1629MQyN/1vOLPoykKsAEukIt7Y1nqDCrmSYt
8YM/JyhFtR9rSahyW3Xv572tTXVed6Wyubw4Y6rsoOhYfanyVTraVIKFqKUaBjb9
inqv2U7jYPQW50cYEjq+eiixpoke29mQ5rM4/+8AWdWwhKXQvI3yq1HmNMK82SBA
HezauiH0nuOfzUoUZYdN3/e/mM9SylifK+YPtodhxdMi1Eq2B/0jue1scpKxeID1
JwUE+2zbOJak2BHd6upg/gxmEfZAgiMlMgGsy/cspMAHh77q+GPU8zyoJSsB/Dzk
5CUmhNQFxF1fuiYplruFiHlvivBCaQpH7XINHXgsVEw4mAsXDwJxt3RWob+h3mFN
wnxudqAwP6cKPNmJNT54OVYVkzyJ9TkPbyazd+d3OBA5H8xKd6xyRgmT/+rPG9ir
AtRQzlyp/o/cgIQlJtGHriIfktiprldauxjw6FhNgGuO8b6rnOS1K1nwp95LxsXg
ASUPvDydr32pcvL/py3crCFEmqERkF1EWQdd/ecLSLw/kdLMAIOJwvyHM4ilFTzt
dt0EKxwMM00ZfV80yQKtv8tgG+VSDOHFRNSuLUyd/tvpWLOQfGVn/V3uAJn0fNuB
xf7klJaz85FxBhpxpIbRVqIyZjhzCw9+Mm8VGS+QlnQIZ2qrzqeyYvTLqiGKoxHt
J4kl+pIuOj/1Prox9L3KNnavo/jE2dG88Vp+KEFro9/2BBMjaOHZk/jbk1EAnfJM
q+/fvnu8ZRaRQVTWwUIbbWPyIQQRXsAhtWhYwowBa2S2l/Kh3f4HSnebYnZA+wOK
I34fLodSelvk2Yizb+UPviMKMzeFy4ywOivburGPkYzmfNLZr3aXTLXLPuYeVQBZ
n7vMPKuDRzcRU16hpb38HiXN33aXj38A1Qy9XjcYo5IikfmuLpIi1kpRxJqRe67V
z3s+WqXN+61dmZonurMB8kSoqeEgoogPWJqRJBBfzsYZX7iaW97uXmSiohcnWG79
SY7E/UNEO/nCKBwWYZMOhcv9PrWqK60Ng3JvXn2dk7gm9GwUU9fzYPswnGBjsWfH
1ksaEBoTJIcvqvIVXEkDqJaDVmS87UA5CGIFEvHEBFwYfwAqktxt6oFe+2G2IU9C
AAipDpnb+EZi1C2OEKU4wkw99ORD3MIKB7UTvRHB9RwsZVH8OY49AmlIbH9nTQIi
d7sK0G5BLanWQ+TXL+pTbh7EbtpBNsHuGwd5GuBRKoxiQO+ca2bvNT/6alOertqA
FDR3df239YKwzKcE/le2zwM2xHNMFmU4IdTOAJIQ1q+gfC57Ku4WkDXdPtl4qiX2
1H0yqN/XiOVQfS8X87qeNysoiLaZ9ka1LrNI7f4pLWeDGc8XYXZRv+/LhEctqheG
MC86oLA/jEkFAjakq/2OnRPLviVNmXXuOcxQvP48fgHGDrYZTP/klOFS8PQk6dIR
ITrxKs0eChD1z2cxAApNFnDGvC2PgxGJcQdXxJGA5LHaR3dQBe3xbo4ZauIc7eEC
6Q3jq3K5LQnyAR30YvcrLm6/Un3jFzLL1l3NGZl7QUaJlN+cmDY+1VMBXAGzvZpg
MHepnbG8e8R+xbqcD4QnceqFCa936x81Yw3iI/dVeb6bGNSxbazBPkw7MdwIfE3y
oQRQSYnV9glMsFBwTPW70bp4JOBTURzXyzPuAYmggrhpkXFrrTK11euiCZmvBIBu
jBDaYqw6w4v+dKWuiMZwPacF6aeaEXJtJsKlwmDJv44CbBUZAAOuuH2W6IUTC8ds
KMz8yKZE+kjxKgmaiAO5zA8n9LIi82MegoVSt2MgdutYcQ2BV6vvGKjFAg9UWjFd
RN4Nbcl+esK+PYeXnceC8NlfUov5M7oTi94zGHfpNZhlCXpiXoZuY1DSjBwMP8JI
m7PvfmDNjIxCmLdP7JeicRi1XAoBDVV08nH7kMsfxkm89Kjf4yoxHurQoFPSvlYu
WHsO0kWY4Rh1w7pkb2oCTcgi/WaMQDwRbJpa/ICI4CatLjCKv5cLD61K7u1ohQeG
PPgd+ImeeGQtNl2xEHwi2UFay9myioiFai3Ojtc+/RG1jJGiRDyuxIpYAGPRQbf6
qOCvIhnbVVtAIsinklh/W70RhFS4me6ObdVES4DxObjxy59jnGyLEm7UYwaYdg/0
LTWGDoX/FlupOC5mmI+l4d3d48+dGrLESWWkhyZrqPi5/lF4J+AVTVGfTLiDBrm7
4fEn7F+yw7OnDtU/xJXv/BLK9cfGmMRULb+E0XJdIZJGTFq5kr/9uZYxQOS0Lc86
ZHHSz14NevZ6GBP916xfRqz+6NmQt21BemAcL4wdwuX4XAjlUaG7oquCl03HSN84
fAL4cY8pIxTGjpxyV0LRUise900rmbRJ66dMKXEMcTS3VfqFIlKg0wTWDqeLJD9v
bvJpOjiI+MaYA621AIjfD4ffOlYbiSyitekZyaNQk9ZpeRwZU7WO07Oni8Yvh46A
I8PABTsi3eNkayocnQsFITIqfj/3KiwUmS+7UwVsziDDmfOp14dAS4bPgw+uX7a6
jl9WEl5yGqImytbiwk9Ctnokf/4yjaZow7ZKuNDXcO5pzQ18w50uL2cIL9S1aXKo
rlTj0WUxuAMvtvEZ+PgMxXGSk5ivpoYrucQQ3ow7ee+tY3skJSNbTip0Axi6tjes
opOTETU6fNhEZD3vz/Cp8tkDgSh9/q0pROAVJqJ3BVf2obg8596FVDREMXSsfrrL
rOsSKpye0hajVVpGADR/ynDV/o4V0vSKqePk7hnzQwwBG/Eb2aTQOcVTSkIAMAkH
Ucz3Ax/FdtxzM5gNtZPx5uPNNjj3KFkPuU3hNp9T0k8oJ6gjvwwNpr048xQEEZwf
R8uMEyItIuoFveAITBQx6PAcsO3m0xedPfh60d/pNd68CtTfr5M4Ie4DX4DOTniX
+TqqBB2riUAt/zDXLwBwN7sjn+n6Ico0BRCifoR1K/abLdNBH0alN7YjfX5LtHoM
gBsIH2OYxQIlxk14rxuVOTyMEYGKSYm603o9LPydmw+OpFdskwBPdM62CfFW9Q+Q
NWQ+YrOBbntWIkaT3L5DPPYFK3I/p2s4rTLd5atsHhBLtGBZydZZiajgSRNrogZ6
riptV7KunehcU0SX9U0EK6GvU4hwWvxmnMCtdN/PkK9NPHs6U0FIMAVDFp1CsAqv
p0iFQLmO9mkWqTogW4bldZnuDussSLbEPvKVCKh/5Wk9gD2JL1lE1CSRtMewOV6w
lUN8EaAZtLLykLjkWWtGXQ0TlExX6KELcPd/BNTrUF54ADVUyd1OImbxKtahfZTO
M5b5lgYsGm/hQmaNLU+Clt606nQFiY2O9rpe4bupW6uT6xJCqLSaLONs0dSshBnc
MhreoctaDEYOngeULNqn5anyO3EQ2f50oqQDqSmTp2W0esfkNhRpRxB2cpkTa/MN
BlGIG0kfg9+xznBYE3QrSb5LMWkHuALQIS4EroVITLYobev917Z4ktaZB+/kRUYr
vssYpXzk97Wkj4NbjL/6UXtk1o6J2xyTdYiZjZaWsGIelWYn7l4lTiRs0Xq5tSKy
jat4mSVXH72Cae3cDyB4PIjsscOZqmoyjTfBjXkxOYICpbK0yRBznnzvE+nYoQsR
tLnjgw0iX0d+5htvtVxjCYbur4sQpgAlgQmLkM/LQHQvX7dSYrQCcvcx5RIfWylw
2spOOI2OiekxXDBCGGWcC1cwibXLPRNK92/kcstGlKLoQ0PWsL0WuhtlJWARbg1q
BCuNUzNge3jcZCREd9/byaLcb0chad4QqhcxzAlg7XvgOZZYsthYJnKnvk69dhK4
5aBVxLc3t1Nj/3v9oHXwZ1UB7N/xfl7FWp4OG6eQxz75zqUK2JnYoTkgG5CQRAQ1
A+nl10KRkLJ//uh98PHFgqHOOqpQD1vWhTarVm/ArDGuZOVsBkc7uqk0RvFNtQRY
8S6WEAPyd/y42eWRMx+67K78/pZsVXk1VaqebQo6rL9IoZz0yHZ+EeG+5nIb0HTN
j8FbDr/EhJAFIGhX1a4IA0eUWfQQwV90VIL1O2BV5A8HRDdxAEZO75u9Z8VEPyy5
k+00ryWKrIwicnwaXUbmYSmMP6Ubdlv3BFexGBLVdO3d78WlAjhfeMsWuTUIt+/W
eSVODxmKRC6a0zh3MYcjU1xURbJZa+fBHb6LvOp4xf0IjWAYUd/2mzRXeIi6I0ln
bthmRO39OQ8mnk3OsJm1h2Lpm9T3w/WgoGbnVcy/HHeUx40jYKuy3IgAEmbviwGs
g45g2E3LNCdgZ7FFnJYpDR4+G7rdC0dZrlcDCqIbeeDsf+rZEIvWOmtNStbgsOdz
SmmuypfW3Awi70yLsnsWfRRMn6duPHytZjWXvnEzke1JzJYIal01RVhBn4il7OmU
RNQaVUhNXcrQC2+xYZ/2YBkY7qhT6URWI/+1xx24LAYxQ+pdyqLeyEaQBYEO1KvW
IcZCBU2KYD46vvoqun9Fbgt5pOXlm/8DKo67NdsDEmq5dk/Xi5CWL2ZGwvL+0iB6
ttEsxjTaokZqxqFT00vEN2SqpI5lwH026WbDw1l5Dw0RqLqSgFz+TTdsTS/UeLGG
C6JzT73Msdbhx10vtWegx041T8dr6Sml3YD1DqXEcmwawQEPRhvgBhnNbmDYgcvf
1PYnPutbz7u1qE2Gsnh299Pm+ErQu0xLJo32rMDqzuTbtCplbLMn3bokb3zEGIJf
U1iq7LpNADR2FM+KLIjwbZVF2Cim6DSZnJKVBM2lBDADz9LN62zJ9zH0VkTEj9rX
eUKDC54IV2BPseUi/Y3DyNuq7UmmNBkVFTM2UrOCP+sMeSbuZIdJ9tjO56uZzaBZ
yqlR5bRWMEM80PLHJ+4fj5YL4CpArucpQnngms6usZ3Ba9ZnvYPXEhXBhEZ3LKwu
z2P326f8x3LtqnJgqvpM+S1+3djLp1HLiaqmOabzlJjvTtnH0CNcFLUyC0u94K5r
6+S3NIkMbo2Zq6WTKhiYC60IUc+MvoTiUJu2ggArSwLzajXprJVLr3abeu+s9AM7
O64pDl8Jz5SIGCKtBf98sSLHFhfIoOhZpiLHkehG3jb/Z/Gjogf7tPY0g20f4Dro
vXoFnZrccFsN1x7j5n/CHms2D+OuLgTvsEqBzloSA5qd9W7yRn2UpC1MxZJsPmp+
btck1RqYzD8/oTz1DovIiuG/jocCAsoDES3i7Tt1t2Z7pP/N+h8aDDTNsWxn393L
VjhZeLzQoE+IQs26rUiKnDM4af/vukxZ1rGrgFTqIPhWPEVQ/fPai/O1KNy2zWTz
MkX6wASEK8lQyib9YGjbiAfyfhI9j/KymBu21hZbbslcW6NoLn8ZtSZtKntmh2RT
hdEJSQebABDppmChBD6TnIU2ff0UVhM3PZ3wGurcHl+PfaX9WetAdpOUQQmq4qz2
4XlgLVoq4lgIOm2sf7Fq4pVT8/QrCXlJjHHgdLtqz1fR+x6bV8C9ZdR1XF1278u2
no5DxoP5crhMPmnd3tL7Fz97wLO1thqNKV9c5ky20/lYLRc+AjMENn3dsvd9E8tL
c6zHsXCz1pLVut2jJD1jzPBT8YOeslVvGAKlG7fD+yB8jeXa/IDqRF42Xxmpv1F9
a7PFk5U6tI3zI5s4I9YOp+F4fFpAr13XHkZK+HZDG2QkH5hXv3EeW8izM3rd47dp
E9469TiV1PiSdsT2CdZqmQTvhTyIze2cukmFgvM4RVXNaDH+AUn1OUOxpJ6odLzN
96PQhZvTLgnBTkT8hXweVYzA0robneBulVpmZFhO1s7dKKnaQTWwLT2/FqRMIarq
covHV7c3BCH2h/hXkXCRwFuyzJ43tqwZS4aXhZ3HSdEUWGWf96EYxi2y95+sB301
4fx05KA5x3STdNCjNDEo86k5yj8kqGMWeLWmgxDolKigpPKd8droooPUURsNqGYl
9UZmrQMfGesp1W9p0BX/+PgH17IOuP2SlFXRo2cB5p3nBCk/7LnIbaXoD9L5QbEw
WZQrOcty6BvSSwlUynB8wtXZx8jiuUFgMRE63sYEF9gVgxvjoE1kDrjzAWW0rbnO
8yb+kJlba2yymsAzIfxanBkdbjspoJX/SOT5mWPUtukVTINnoMEJ51EXQ8HtI1nM
l84xdT8jZg6hlU8mj2vcNBov7rHyGcXQQMaP6TvmoPFKBWyb331Vz2D3ST72J01P
cj+YKbSSjKvWMw1ZJ5kiApgu1LrHY9u9iNo0PnFTMuvd/es8ISLX2DZ9R/wMBXwP
T7BIZIMu4zDbDw0GHz6IVqwX9k8RbG6Ua4v38LCVq3lamqA/XQfVtkWV4/+czjPy
s5BOUpRShc7ig7P42ZbE2jQ5QOE0OLRjtk4gujUg+/tEttI1z6mtcImB4c3EfDlC
4iBfGBPaNxjXxbo9Jud/4+R50xxmrZrwiPcouAv4ftyvAbWTgu3k7sL8nX4pb9Gj
Rg06Fxhzdihw3NDvtysu9OlkFOrL1y3yAmMuc4X/6hl+EwbZByTc3mFrqFosnkL0
EzuBnw7A6ZhptONdy/K8u30JkMT7lXlAg3bE2iBnU1aOOM5Wuxz6T/fD9Mz1m5b8
NfGz/7H6Vyq6W5Oz8AAVju8muGx9oRzwfniBesBElN5wUkvjSwWJ3vzqW1OCIrfI
CVsVvsAfPoz0RACsI2VnTCDQ9yVN6B3x52B0GtKjY5X+1ATTHg3lKyL70ZVuCITA
4wdRvgVrp6y+VVsEENZDHCkVlJ+cP+IPE5ITqCp0D3bnp41IbE3rEQIQxdx5sQzS
SY2MZW0M68LgbekDBmetrY7gUy7Sg53XHULyTGTfD0gUMylknKevJWJw+YevBw/W
mrD7BCYaHIq4NC3I9P9pP0P7+AcVSQHA9ZNVZSU9eFaKTB5yHpOsVpgi6Vs77VUk
JBnrKtnb3MseGREwiZxGN/knvUCSfsDqqv5pqhAeayZQe0TGiCQs1WIBkmUGU+OD
GT3o2BCZY5c04c2prHLU92I+uRFCrHDn23qDAMyOlFRb8BWAcGJ594anTXEgNjCb
qpygmUX5W7cUEU1GqoRJZc7Pljq20UlOjWQqnD1F4bc1je4MrMrTxQLYjSyDLnnp
PBzr6s9sN0QN/8kiKJZFFgoYRrV3gscm9RwjkzFfLlRfUmP1m+oan+v9p70X2D1O
2Jmx2sTAlW+3e5wiS0nBmTtFC4rCqdW+k071fHkJajgLRpUpeAp8qhkRMeGs8/nH
7k34IBv26axa65mjii6v45GW9XA8vgJq1rw8+zmGx9JHSY1pce+Sp1zS1AD45+tS
aqNay5VgHtb42XhimOE/jT/bLblZe+wFBs7e8n6xu5l/HfDbqA4dhqK3H3GdYQ1I
35Nyc53CSGgW61Or2hM31UvMJ6AjMPlfrZPR+NNUBe8H245Dz6c0SrEfTjzpnuY1
Obp9OhTkrVBAWtJ/X9dh3dIKbBSwqI610RhkwXdbogZESlkxKiC7TtrPtVCRaXbe
uTWUtSXZ933KRfvyN6HbnZKOShgVav90SM2SHo81ViNquGJxLW4KtRV2gnkAc/2s
6nc7fGZKaduCAdn53EMyvbPoQesFp+bzE1oTOvEGNtdXj7CUbVpw9KRKyRfYQk8z
8DhCL3HV0rDwrvIy0QR6BMEQfxMDp4KqDuFhDP2qB0M2dQ3U32NVQH23PhPBhgOS
IOwNZmwCV4ANA3GIp6smG2fy1tYaws4/KBL4/46CrX0wn8+cgHTq9K6S91s/t0q+
Sfdjtfb1CidyqHws5vhBqSIc4J0LPXUZb9xA4u6SjdQd3tPqeZmrozFydACXHD99
nPo3T2/fPdSQt9rptL9RQzayCnCBjDKsv2f38w+43LtV61BRPVRQ4itKQyuMwo3x
X8P682yTIww3IaqPlOkUXErSozIV1PkyRajN38n+dWXnR52pxRoI5Ixxpq+JXFS+
/3LecYg4ifi/RqS11QQ8a/RaCanHPWtE1gV7jQfetnmnBRTZLRNfST8R/0boB0cg
znKG/zk4NLno8gpPhCzzGTc6BkJj8jMWLZhZb3S+a3yFP2EdFJh3QsCkLoN7Rddw
1BbHuaT3W96r0GPDsd2SdLb+HvoP5YHKT1PqCRvRL7wBbiuOnRU+sCI7eAnl3/dP
alW2+ad873Qz1C8dZzdIR14/tE2ZTObdaeCXP1mjk5pBc1sV2bRPf9Cfpn6j7hKZ
QtdE5cW9TaOcjCEtAPUBgtVFiYs/4j25NIKUvs30kDgnbemOTyAaoe4r+w1Fipbc
Bbi0sYifaBpDJyKNiijq40skPkNjh+07EFppRQhagTlDoCln8Htp9V2ELnOXRBbs
GP1Eio8r9Ad7r+3es6XGUk9UtMd4Q17QoXEnnRjDirO9UBp3dFUrEgvkIMeJNPoF
Bmu3dJQtpXDfYzCIXPmC8WEMJBYBJWq933TcuMhxg++GSXW9nfelGoc+rrosdgBv
spvcNeH+RgCGDNId1tY7hQjowl80t9mQ9AWvuLSAbwaPDzrxScNd3eSWL4B2SV1v
tOyTIHZ/NVAxg14OJFTko6oL1louRq43bWOAqyWXB/Dys0Q7+KD45C03pGTryL+F
g0OyHWAZqkobs931OTWhY5iOgHViBFvbD5EF+X16gRdtS6AL/6rb85eb4ydZ8qQv
0LC6fZVx03r1Lk9FUl5bRpcYh6ktQzQ9nR5/+XeXFiq6rNoQsfm2FBdWsFlMVavm
f/zz9lKhcDMBVsSy4gGvOASu/cii7A1YsWEXUYEynmRtvfsf15HZvSYdzLYU+hE4
lgs2uGLgTiM+hV6Gaei2jfc4LFHiKbc5YdlROS8DZv8oJP9TE+waFKhqXzFUZ9nZ
Nk1ADybrm5D7r+LOd20Q+Z8opoePtKujFyEgbRpMU/uCNeDyFC7qYK4ES9GWJ48R
oSCY+d0HXkavAjnNRc8/jM82ZUWkM0o+9etaA2SFJkr1akFWeHM1wfVJYYxuM1SJ
xOcokNlKe5NWUNE+1cj2Si7poyQ1Pq2z+G+owe+sbwBuxdKKmVH5vLG0CaoJIWRu
yhA4j2vNWdLMCW8ueCzI4kwycMeD4P5LY/ijJV++ZefkZGu7f4OrTTyeIuYkFYvr
iFDzbTykLI8Ir6kwONe7XsWLjlx58AnOy+s8NxIN+1QBndY3RpoWXT/2KQk+7kEV
yepbyQYUsVq//svHF47pyrbfIyfGRjERf9R66WcOImERQbrE9D2RmOxklx+y6NQa
fIpumWDOvcK5qcITvKqYCxCnHnokwf48ZQUnTgwPXJWKqS/pj+nO7fcduL+YG3qP
QdXVcFdCkB30cDz1X1ogqgRTTgei2t7E6sA9IFryBLk3gDNk2dsupUsUzztYy0fG
0LlcQcF9bf7MEnxEdS+Ygtb3ED6KlG9ytZjRw4eZVrBmNrNOsA4vz+620V2ml2Sw
17eXwGzjubEUxNpQYbCmtsJmYOq/bDJM9PU0TI97N0b7FOAP1jqFtPV/G6ZRQzYk
qSxct/VHbv73KSQTxYEZbK99p3HbD/ZChzjyilOV+OLdVH6qGrMhhZ6ulpXbw5Lu
Ou393VLE7DjtVZcKViviovbzyfr+urHA/Rft7+Rr5RKHM7yo6uRCXyFzu/bDn7uY
N6kHiAUVHRLhw203oJqelNY3WL+QZt76BKMj3bal0/9ClIybM26i5w+GG0JW0eSx
jWbS+EGIas19sJQd7dQT4DDXROPRGM4W50HnmMpCMN2ZQ51OhmMp9b+FWxL88jIo
L4sIn0JXOlfJTU7E07thfa8dxAvP2/6rxUL41vxATR+NbRUyhOgytNMf/Db+FCcM
K1N5ILYLtOu4s1Tp/IJ98lGhHDAdMdeOwStiuLao337Cw5PZFYs5KTt/cPuP8tIN
3/oNhUOEovnBts1kaFaW01h/ad7sccf7igd9+FrvBWLl5LU0oviW+PEGKRHBfiUn
QoBbWs9Iz15AA9jbOG8XD0zL3wcqT6A2rWuDteDHkc2UjWOTIVzSm7o4w2ytOb8Y
C6bc6ZVNBD2Y+OUklDzYsODe4s3Q3b8ji76WqcZZiPxAedXH5QTnnwEHY+5uZS8m
5gQLC6HiLZ5gz01SwwCUazwcNJOx8RKo5zSqZPhcvoCYYZy9sURGOaYc9KeMV56N
ovVIKS5vd78k7S8dZ51KXaUtXDkAcbQsTyxzbKyRcI8kI52LxrZAQrOs81QdFYiz
kPLYleRfz4VDRfgifl7DxSd4AMvO5zBf2EgGRPCHvaDb/9jDjcKmgLBX5YjwAvCO
chQ9tvgOccX5owEyvnGAgQM4Oebg9pjC7p4gD5unvfE0CAOP0Ko/w9jipZkrt7BZ
81jz724uqK+dRcRTTCUUYW34Y2rehNxS4h7ZhiRODN6ad4a25RLbjt2gASlweogs
nwxWwobQeWat24KS2NZj3sQd+2LJOoGgo5O3yEJTWi7WoIE56eYxDknZnPe2sAqt
Ygmt6izRt5F9sjbbmcFXv9qWsi0Dpo0iysuDg2AO0jMZPhCq0B0JGPd/jhade7jT
90vY5QJNUQwjYR+vABtN2bU1cfBRVwcXFHqoD4cRCMPtWZ4+DgKZRFvKSVnhonbi
1oT8iw7gJvQhwNoiECoPnF0k5q7fBPrJHDZ/HE7NbrR/G80GLoQ0TygS9m+XSfQP
LU5Qmh10TYnI0gGFa9miiU+TkTGpD/L1e1+/Pe23+gOfLSUNrhlacSHQ3eVvi9hI
jPz2hkkQgV2iXHUMQPi1XP5z8z/oLPnFsjO7nhqVWEgZQF5XVxPuUxYH1EVE6n7r
dpJgOFL0Ys4Pmw4oxooYClyWFP/xDklsTCdRYfNBR5hoF8VA+4ZEl8MWnD0IrRaP
9AhptL+8U0BFgxyWqaVws0G94Q+ByM2t1wPY6bZonPBedmtdH219EPJY4jEGpxQK
Iw05fCMoJqL3yFDNH1rZBF29/n/vbUlOAiTaort8jA3mk8NOWym0I7SkoR1ldLgZ
00/HlUUf0oLbqveDqFDNBRG7g1ZyMJjo45MkUxjZ0FBqr3nDqNq4GagJ/6xc6uiG
kjTxlX97VdA5ylwl1rDrJzF4KHiYq0xB7KVP4P72O6CYWXcRclzJ+Hko9Y+6zcu0
a9JQ3AksMFlZskZt+s4nNnXRxlMM1njSrUrR6N4bAtmrdsJm76BoxhgNhA3qk3Cb
TplWnlLGYLwC7afpyP1rCOfeojHcd94CPNdVFgCmk8kUd6MQ8LiqCqvgknMa6UVx
rDTNYjpb9WYopMBI/LLGrb7XQw8GEZb1O1FlVCPX+KKGPV4onEhtGLP0kj8R6MWl
gU/Hf2/8nEXTvse0mAZxf6jvmdqF9kztxQr4aRffwzHHxkmMb7EocXCxxUvzGlan
hHLGUknQeLyhd1xnUPVe/lAOzokgnxLFgD2Qff/DOOHYXsBhfoeDHV9U1G9768wo
3qiecdvRJOiLEpKbc9qrBUk2RZi9mZPrZiFcDF4GuDXXoUcAy52oTnw9g1FtTeXo
jaxeyoeGeGXYHuBZDixOQUUKKUCK1awPer2Rp+jtOnpG2iU6PeuN2muJ3qt12NOY
9TP2lA8f18eh3CfyW7GGk6SrtYJu/3K4Y0HlKIFASRkrKDrouzpxxu2g7fKor54F
AqMUQN958e/K8Y1zsn0Z82Sdqt4NjQjhpTdLVnUW4Whsm2R6n1aW657yc9QxSr+I
HKVl8ZajuBfzeR4mMke/DugiDE/5JVORfEG32bir8HNHNsx0XZFu7eCp5uu5NVsR
7xB2esTS/AxojWbxV/wOxRwwZ9+ZmMfFvCAI33u4qNlbLlw7CYQzst2QYd0sELuG
hMDAj/h7ymSpHa1TT3jpo4zVoyM5ci+oGOvvyzf7CfNQw3XcxoLTO5Z+N9mUAI69
3hHPbEtsNgC4hI19x+PHKmYXDTkMgj/kMIiTEerkOtUg1vUmmreVYzUqlyCkOqB5
06kX/d/4fETiHNlBPKvY5w3XmUyEIFqoxvOiz+HMRYyM+HVuOf4nXf4nAmf3hUFd
zh/6rPh+IvQr8EczfwUqrBM4VfFFUeUJzZLFJxilzn6OHFqK2JxK6pWfH7p7pJsj
5+KuUtj07JyUqapDGhXlrtGwWkdFsCz6dpWXfYm5/rYU5OyOMJUl4cQAG++wRFX3
Ickt2q0Rd80qIRzpqo/sGibeZnhkjRHDrL1P38YMacJEDdVlwaMOEgpV3qTK/7Kc
9O9Z5Q0NaXs+MJeelKd1YNW5vDEXMo6UiCNVyTQjnZ0A0dL9hlB5s2Aof7u8t+D4
csuPXQCknQEnQQ3csh3BhH+cTB9OTkjhx/LWPH7p8mC9TWOaN7LmQc993wESfmvQ
27K7vfV8JlWbmPoBvp8OJjURUPGhKgXe9klNXODDKhLHMZJupj4p7z6AkPOMBUY4
tfEcUm06tQbmxo9NMlunSQ17jXtOuuirFkJ3E5mAM/AfiF/ie/z8Px/LhD8dYikl
ixCBekkTvOKc6J4eIP5PSDAeDSKSxV1oiWe1u0hxLHaMyyfpCBtuUvW00655Y+U5
nMqcq3engTWNXGvyayXBdUr1+EAaCEeVrNdY5h2nA7mf2fK/HlTCffWAJAesk5Wt
dfrMMS0gE/utpui9BBhIsXR6+XCESHrD5WleUKgM3ARRUMhG3QjEhmBL2ifuaKBg
1tVrPrlJoBHOzi8sH0NYBgc7/uGCQ7cONItLSbM/EjkITQlVnLJiioP/JD3skHoZ
Z/mOZd6kncWaTKSvp1xL/q0itkXsaSUkvWlHozTO/YpCVKll00jU8EupZbAsZ0Sv
gzvwpn/LLaAQtf3st4T1JEpry8y7ZdXcYZT4IoPLboaWKFBTDwYLOij/0Bis1/2X
kz/X2WVxpqPjUH/wuvFcIt5y0vJd251gEEF6qmCVan1S6tpWQl8QesDEbXmtsfH/
od0sxKV421o2XR4OtmC7OiOXHJp/cTIsjS4aq+tFNvRAa/vO335dRJQpnsMcTy1U
Rc7Yj/nBrDRsaJgf1AWS2Qguv3wGLmnYlU5ctfof5ZIdlJ6qPUwypTIKz0DzMkBl
LfMyXmbTYyLiH+lFuZf/YkrE94DVj2KCkuZ3lkoOyRCAfbVvIYpAFtmMJDrIfUjs
Y53+/ThxUQcqH8E+B45AbgLTxdhvAt0RuJBuB6dhpjpxN8v5tC4Eu90Nn5PmHa7U
lkCXklDn0z92ZVOcTKtPcLIDvBXsY7V1EOxUUXkoLU3dyRYk2qsVJOBCqE2EiX5E
P3eaBgc+MwjKD8gZMwLwAdQkkr2X36qJmBHiMUWSn5i1tw/9DDOaGGkx2PeAHbvZ
hrTg8ySjOHVh3ARnkDSZwDJq6E/khBxZSEnVlJfsyQCCIw1cTBbV5Izxo8zgjkGM
YINN11fXd4CT34IFtw3nhojsqmNg9sq7Or98VayufWDx1EGqyzTEWWclCVvNYeyr
aLG/T0vxAja7fpOG2HMJm2vuA48Ch3rU0GSnqhNxaiCZdnEOsa4FbQlFwr8Bihhu
LL7Ma+tFmGo1GrQIDEtCsrHbISGi7/1PnY7C9GXiBKn97kR8hwmq5Eo3ipdKO0sK
MmuOg4hqIXWji0BLXyUTML9iyKfOykYGzRnKi0VhG/borgdz9ai1XIhH5GYE1NuV
ykjS3bWbP9axVLrKaeROGN46lU5zlbv8rckvEu3YXf69IoSV4IZQgCceuCY8KuJ6
78UtuZ2UDGJIkODRviBP/U4jNQXsedSmR4u/9eEHzMZp+fXmApC0AMMEYM6/pv3S
ty8fXmc5TyvgqsLJ/8ff2xRwjV6nAQiGkFVK4yIXBeE6X/9FyRzYopknaOf+uqTT
7LkSCX1FjtOFZ1FLpDBOYAm39UFeh47eZDsHiAgDP/DjjfffAWfF9KDqzDv18yn9
fc0anOp+Adyg8Nj3XWVpTOJrpwYwI08VnlM5uOpBmC+hsRrj6YAjEOjv8u0Nqzdj
DnMymteVeXMb/qifAZesFgAPp9H8BlM/9Sb/cGSO4iJpl1A3GYIPIVgV3NoKFnrP
lJJbOhZNX8nI08/IyG6yNdjophHq0t5ldzBil03HM+9OBAKiFg+0kR8Z2+SFU7xZ
Kx2vQoccoxkgIRDPEr/GPSJQ8PqsQGNPfvgUI4fvLbAZTLMi9cyGo3kvWSUYAJBS
zvq4RYMJ9V/uuJ5Hd5tk3g3/7gzsLP3Elv0iUUerd5aLzrx11oXVo/gMptkSszH0
ofFf3En1Ib6Hsg98DhrmAm0IVptdiscDREtYQlzsq801lzaiCE4miTV+M7YyZbkS
qWmuRbVhl8MT1jjjaAAff+KQnNVWkqQxpM0Pg2tTuorBQkdgFYnUxPfYna023kcb
PBDbySmB5ceXyoiH3VnTK8wGJNg54kTkzJZbzhZdVpqVmXeRkNmrKitMUFA18kJ8
QVhkmiKE22/fjoojEZ+7LIq2LF52PBU66O/ekD5oUYeom34GbtOZ0k0HiK/MuGsH
pgOj+MDPNIQtBpOrwxc9ytK0Ys2K46BF65RgZ6y5W5ALkLmOqFXxmmbWLYwlNZ2i
UT1zqGSBRD5u0UPudqv1mFlerAK379ztQWdSTQWVfeOZ4ZSRuEAiUhGR5p0mg1SA
zLmnYDhDsG5eYzEQjW+NSBnSn5WfOjeW9YXGwfj+r/zbfaJ9r2473xe1NcVMooOv
+i+H63JMAG5Mz+4t4793mRcmZpxOKep50Oe0YLT/QyhMh7Fu8cB6sfxzjqPaNF2U
EYP3DY0AJwGyYTtwD0WmCXzoX+BvLKsohHLHepQyDg87l8kJd+bzsFpKPCx+3Jnd
yP6yxQ3LXuDj95cjkMuSj85t8HRMueDqkTHXXyh95SpAxCIpKLVOCTOPDcTxXJzb
RlFv/xAxoBHZaJZVTj62AJEIxqsRpmtjuzF3BWfZqbdqtAvfva4+tX06+92EuOaV
Rs4x3BJQ192jqIPsQ3oOxlZvq/YtHGEpmj73pMHpUB0d97mJ25iJG3kvO4/ks1yX
EK2uR9JCLsJvhnR1ao2scLA9eKp0wlaVBhlHGiDvkGlWfhjuEAnIjVbOgdHx9vj4
pJ4GvbR1js+dd4HlK/lMVgNX/zBECRAlbBlmqTyy2sUo1Duj+Q77tNtrK4rEZN6Z
WspmMuFe13Kiqae0iwi6I61hkEo0zSBONvbAGaHRY/QpD/Y7qxam+GMUYokTWVik
o1ZwZbaeFjMUcgAVEArgcPYCIYtBiv9fGhTZGt73IICn4RVLEBzB518AzAiTDg1x
Cvi7+6YTHW22bTm4o4yAJmS+MVjVCmdUavQsBypGlJOoVJPk1NoGDG2KN1v/uMwV
c91L1pSC86f4s61J0guTNrtoDxyBkzAfiFFIKXnZRJHidXtmImy41Il2G+Qm9OYg
5oZVQkGgF1sYea1YD4NBlSJ97X1HUDnVKGmHZtcNm8EdrOWFAhb5b9Va+UxlmRCz
YM4MkpS6ardFhigP5JTu/ctASoSGwd0KQQjLqMqjSybx2s5gR6dYVFPaN9aTXMhG
bYAz8lJoyk0kJAMimKAr6UpTVmMUwcVrcZC1Ti1qOcLAQFTKB9nDZOiImv0FY0uh
b6gAWwsWQHP8a+LbXlgRSnWcSqIS8x8xzluvLXF49/U6gCR+TQQMCBgPcO/b4UYT
kib2R55wZaXe2rfYL7gjReOwPBb8+E4fOf8y34HAJ6w6wEsN5BbDhfh4LXJHqDxe
hIfUpJHCZ7uEEqGripMO0Od9RZZGpSY+2vO2oNvkW4FmOarI4YwY/OEAO/XPTPRL
zU1NmItWnd9s02T922S4YCsOG0fKs/bxvvpHqylBnEpK4ekOW8D1Mw8cqRXIYfaD
NTMSHyBytvVyBRPGa04SQ3NkE9mDyo4tiffoerbk2Q+UiehH54yfBZHTdj8DRKLe
lDwRS7qb4xB0aTJSvAsFVGLw0M9kfR/sbU9V8x0rLGhR8LeOIZM0qWYTtyRu/wwO
bqWcTgXoIjSsAvVyqQ/Yz6qJGxwAOaIT++M2+4fU32H5jAn1gZNa43qlk7I8PqMY
nZ+xVQbhi7/ZOEIMlxVrW7c4wY9e/mzaDC0mlWvR96wu4hAQdJPs8vglVkCR91A+
8vXX8Ox9yb2FXHyBFarK+F2Qv83SAiseBFVElUi2g6+iGbdwtScMJ6lqh3j6ITx0
NI5t+R+kfmLPJmZAFp7HZONWewSgXSV4icRkKvsZQcpMVGvTSR2gUQj/CqzYSpnV
1BKs5V323Zic9+7AAJ4OKoXvYrWUXdcnXinrDjuqLarFwkBvuVrnapiXoUz+Wita
ntebFntrH3rI8GnGM8mEElTynX8yME/8iIpNT1ZLxJ5Fxr/jcAxb/xPrKCVFOYV/
BEwQr+SHVlbq/aozcHbUccLUR+1OLd8hFFMk7L7nrSYF7gO8n1JA0SDfXaC7Gl6p
n//X2MpnEM2OmFmtdyOuSuheISa6W/eJ7y90WTFDQuIh3fhTtggC5GAC2tNWhR1j
XjMUD46/KvKiwhNmoQe+O48gIMAqftksd5kwsXaHse82Aa2r8N+uIE6OOcU1mLoA
DRwX0LDalmKdnMOl0Wz5JMJhMgLreaD4xo+p/VzzpcZQ5mgb6mb9jl6ydsoxKQ2q
CTfhltzAdi3gFoZILOFjQuNA0SjeTWm3BC3oaxf0YftTpdzlLjCbW9I+mJPolI2C
HBThMpLN5u/CnwdBiquSblRUzWxkbTvX99QpAJvO7CC6ZBUIl4XQcwGlPJpK3vKk
C1oHUUo2pJ4GI1OEdAeobASmiAh6Ff6soAK3zBHgTVxH3E6QENcJsOVjNsPL3bQ6
1lJKDDHeoFYASOF0Bb9eGtf7TL4TuuWGWmSPcPx3IUKeUHflfkb15eTDP2C6AQ44
HDwtYCGlZO00DyamB/fuABdqvn0kQmYCgjGAMLG6u/TLDgqI2PhJ86G+4if11hn/
yByHylzIil0QucWFlJP6i2aJvFR+rG0Tm5NLeO9bxin+NXkVoaSoDjqD39J/nG0b
ao6ygHNXOEF5XHXOFNa//gc/iJSumPDCKEMPpzXMEzXkJFKlHDXPLB+FiP5Gq1cB
UNznIqrVFYHIGn8+Tb9NPUel1qoUBWkO426UAUqXJJhAzYCUqBtSHh75PVkEuUhs
e684EhUA9gsh4t4N/kHk5KeHxH9TvppIoiZqEIxxX7Rk29e1STNcQUdJ5TmVuKBG
VLHWBaDHBdlYcjSMo/Cw3uWoriA/MLoQTpXZbwNr/MtZoHUpY854RGAMoBCJGJ8c
MinbpvnMAvBgAv40Kq6QrGHvJf02OG/ubHnFTxo33oLJbsxay5fGaqHxVu0aX9oP
WNyeDo7Pvl8lS/rKeGbqEKMpfkzm0xGvxywnnhUDk7Q3Fd2gZbsUPjY7/SoMd7qV
uC4QL1sAYNeYiNCsaHganpv754qFnRyT6oj8OR/O+7HBRQpoyix00kqk2h3T3Gjw
dGy3PiscO5pvtk/0Xp1VePpHnYUH3GF1l7hRtWNnIa9VCc0Gi0nlZK/WlleAFQGk
ZCBB+GXn6wchTlFaxwzle8gFcIi8c+RkjX5XPuIXbT3QgrFjkeDi+MzglZyOwshm
5q8dxFajKgai/sgP9N/SWIUe8+8H2+dksF026nzJLHDSBckvci9kk41nQ6kF2Zth
m4251YTjDaMeTP0spKS00j8QZyH9APFwWrRd90h6Yi/QvMNqmLiN3NpCCyOWf0rc
J9K4JvT4MH9ggigQB5HuACua67ryvTrIpEbxjrvUJ6Bjo3qsCXPnFJ0guSBdL8uy
nbmIZ2Hwm3pEDEz9Lu8YTNndGdOTo0WnpVWOj7t8Getom/E+6Tl90rc0/+s9lZwa
atqWq7zx+WJ7w2qmsUtoiEwL2PemIKL8MVqWFYm1XxPpf32jsHt1i5YkN+AiEUEq
v8U7+RQEp19omHcja2QpjOP4z8D9EF8mIcMyqkC+7tBWOjvdl6WZrrSyXsozgSWP
laC1ju4jCh8aoMHG9Eu/NSKSC/Z1bmH5JM57LkwebG3TcAcobn4lZjzya/9qR7W/
h9Z+8uYPbKMHgF6qjXoBI6ldsRqkbVbUyGikX86CT6HUFp1uNIiJTkxWG5AEGXS+
YPywkpIxQenni5AcbSRPeAW/Qldh5HjYWhj3dqK5whhFbZzAQrj/jRemlXLp2L1+
q29Whs5vSUG+NPwIaDyfgBxAvZ2zW8igPKbhdvREdiRDMLcGTAGFFcb3M2X5I8Cv
21+KJ2lMCFT5AkmUdMu+Qwqny+er4V5l6pV+qnFjj4ZR/LRYDrETzpQsR0IVzpLZ
SkSJtz02h/ds9j+xmUe5v1SeSvjVXnDnc/HMF0QIvw6Ob3JDBfCKRXceU7AGgCRU
/Cqo9yAv4DYcERiZ8nG/RxqTtkrkWQvd+lVjtSja0hH1HidEhRI/WdUuprsh6SZh
FDGLSijSQIs7Xw9rJOzGFbgbhQYUGhMx7i1N015AUIUiuY8Wsg3GvcxHTCiCltF4
akJ1bYKrxItEtuAB6qVmvuBVUY9c1bMUeCBQFy5bfy/v3N9eq1VfKOUtympTI9fw
74ZxIZZEkZC1fXcUpmeiumN5YFOzRMqvUNCSliRY0UT1RqnkAo/vxuQ+zflXeDbW
+Tn6J25gwFODwSYtOcmr04lQhzttLm3cXB61CEZzuRxquHBVkMlfcJXIctawstw4
4EQAIz7lSGIbC0x59JXSGWq6l8pXmhyQBUhUD5ajnYqA+dqZeh5gLkLdZzYQIR7C
sw9BmR6SnOSkQjZllCAnF+Hm4ls7/aQkzBpuJsAtM+pj379mKK+LbrIFujXI966I
FhNR8A7NbkzSEa3g74TMP+PNSmZkzSAs1XxqemMOCwUMIcIWZ4V0pSkwaWuarEu3
1+WFvtDx3ZzZIBJcOPjaMPtMj97nixjh1JxBHr8jMMn7zpnJnxutnhfRAO35ErH/
5Z7IeCSNtPPgakWb0IIkZOQIyQrWJsPxgsnN2HY1CkC+2Jh7yWx6E22ZB7axT4/Y
90y1DNJbUVoOpXU9MIsskJgeBtWPS+r3xbXraNF2v0gaxFUP/L/xo7FJAea8jmh4
WW6tjsy8idQ/RCjY3eJItfysVG+FMn5sOHADcKj6Nmf6taZ0+rFYlZFPb00VZ/b6
7AlLw25UjSVL/Wc+JC6HmiWseGltjLRmQaTbwl5vUH1v6tqdlHxG/JU0J/VgtxGw
uLMnlijWrwyNFCz156znHakIBj0plPJ4HYxiPZIcvP6q2U0CSotsGWmoSN7WQtzl
1z7ncq4KrjPmN8+xhRm7MjJtPFDP2ByzZ2k6qNSJBmLvpa5r5zbx47Qa007lK1dy
9pJewdDm3po1SYivsWMkM3wQDxIacJpSYkf4AVH1P2UuK21j9lqSeFDyixXT9HNi
9P9p/Ehpr3kLSGPxjZALp8SDV6OtjW2JcIYQQCGt2GX/cjAAxMcpfxfekQ8E7/8n
AL3mJJUg9CLTNxprOVcVB4Ks3ha39kccPzm1oBMD6ZGHAJCoQnS8NIm80mripcp1
GYr6BenvfOWgh6uNemP0hXeAmo3EQzxIZRiCuCAjggBgWpm4w3fHl1KXpH8Pj+Dv
J1SojBlD7XoP3D+ALjOuR7sLUC0idiv2rIV+SObrqwhEslW2MUWK2Np6yKAslMVV
pAEQYBflZViIcmjIcM2j0ZFe0qc2P4Cr7cRMHYVtHO3l1ORUaDHK2XFsYkw2FbXe
+sBwEtl5ixIYQEwFqyjDC0HirY7sif1VRHTusIe+rP9yPilnOtizfjBEjVOAJLba
Htso190dgppITbMIYZRETIzs2Z9HpLULxbe4ZB9lnmxd5kWTdeQZ89TlcsrmdreR
l43dx+xkhER2mECQTX/ZGJnw3cno37dVGU7pO2luQLggOCHXGGzzYUR+vMlnBc/O
aRUJwou7wEmE3Nxi4vmZ4azsBDmPg6aothyac8tDPA+6VA75WHAQK1R539cTqYJh
9aiWCnThx/gmsazEOlGVO3rWVnjRPP+LLt4Ou8gobXD1evNyBzVGjEsW7xaroRK5
d3WHfQIavRqy8QB2NoHsW0n6+sG6oGDdaPis/6u5Jd5kddrHhB+V4hCW4DUBsRFH
JCq6pQE32cmWNAsdqo/9bMZZW/If523T+Yo+iT+noYsMVbtTC7t8BaDSEBHvgWgm
nVzgUamF80sTFZjr7uMZ0vh+h3EarmV/FdEK2zYR+dFLDUDulJd5O7yfjDUyLEcR
sCePJR+C5HAMi8RxWX7P3MpdAXjRcYp5SRJzRwGef6jB0uMtH8gowggPJeYwo65E
7lv2uFmfmeX/VgPnCXsteu3YYMBHP0EX23MnvVaeKxr2ueB/VYZ/CkZOIXjzHIL8
QxIDW1Cu5JUhk503FoA1h3b9s1Pl3SvJ/nujFjpvRPYqfIFyBxEo74csZ5Emf7Z6
Ckn4QdB+LBa6Y3noWEsDXTs+30tSQn35Y/HjjediQke6KKUL2wioTBk5OfrjLo/z
jflFpLGUh25SHoFVwhfmu80HewU9WtbHj6oUqfcQoFfC/gnpn+eVA4lFpy2+PSQr
zGLEQXT8hlVKKIKqTFvJXlQ90Q4h0mz7W5usv/tGGaNjK8fPj0lZADvxHOel9ucw
rLgY8ic6OBpbTl1Ll823xsZ5VBPFGj/kI+wK1f9CCQTo11/8pSU6b4pigbeevg7E
Hu9hsuIx43QMdUWThI1DYUoaFMnyLKz2bDZCkYfY5VSEU5ysHRewIol0TlbNI5JP
VmUyuNkDNV//a8L2e13czcsfymbPP9K+fDfLmc4Hssj+z3SZdlcf8rOrLmiFTdWK
MSTTNo7tjuq1R3dBW24jfj3teGIVc4L4FXv597CoFOZilg5OV3TycKqgCixIfE6G
BoulX/zm2iPJzCACnXbif/dsVlq3hvZe64j7yxkDtBal6gJGXaf/rO3lHwSon+ly
b+r7q2QHOM7TQK7GBfpnlWy9K8/JLBkFEYbwbulLhNTs21mHaB/DYhwPfLuhX6Ua
jc59JhplY1349FVuZQP0ZYTF84px+sWrdklDOWFrN3tQCRVMB34Id3BapPal3Gc1
ld+1HZ2lLYvWC5py9m5o3v/P7cm1ioAoatLqAz/Jna7yps/IMoBW7ETxu4TX1rfh
DPp0hgsNu2lH7W9hlazv9L9a3TIXDgwtN8WR3jTrnNpKLRtOZEZdFxNBgCRuoSEQ
DTo9lp+/Ky6XLjiC1n4y5vtHtkfIzWPVwfUnc2RPQMecirRik2+k77ui090fz535
oqbYtBKSnfovwR7TFYFpp3UkVcng3e0Y9g1fjBZNh2tlZ15TZFm5ah/fjQogfnQI
9OsUz9Abpdl07MpLzGbSgB5EGB/jATWX1LSODUtqUBH1+nTY26zYOjP3c4/yMGqX
NdHDEOIrMoLCzb3+PUKJjcXEtnL+lzOJRGR9gJZXW9DrgT0PFwBTo+Xu6SZW65BF
4MqS8NmywRE/95GDoxdVpGZD5l++CMGmHmpgD0XbzncxY2HIvFAfPblVtTyPIkNQ
TlG6ztWCaCCuVYU2dWrCuXEO8YsL5bdm0AHc3rtohsKlybQIHq/OCP4AK1zzBK2/
Z+jEaKARuQ33XLaCTP2MYPCtsYcloFdqGJzFH9KXJAZDeIkv6EJ+1UpHpE/BIMbr
WBIJAJZ+3CcF6oGFY4IbbyLvm8nBBGUZmZdchMlXnR6Zn3o1/4HpO3qqFaoCk9fO
nDcFFV/BHe84E7SbVfFnKtU2vCFbBOV3+C4N+thDFN+Wr2/USzvvvyxk3F1ZVkvg
GEc6BMxlWuRpHo+9/+8uve5Eq6WKWwQ3arYoS5ZgtEg3jzTARvJ2RonA1VXPG7/s
NhfJeQDdVIza262IxhutH2q9ckI2L9aIAZAESrv8/7MUF2K2wrFvGQnUx+aiIDSN
AUW1TZVfup+ImYF/cxx6OQJ6RgVd5fk+agqz2Xe28Jbf7Z8oHIScON5iM7fSrpA9
XTCEIY5gDwSi1hS4QPjH+fRhQvEkiX7ADwDbi5x6LZrs+uaoj0UUptzotFbmc9M+
jG0a3PrPkyA+gkLDivhPjP+qBfdrRE1m4cfb2YZz12Nql6Tloe2pG1KwqRaxLWFG
xXz3EdazffuFhq5NL/Ruv/msvk/osSQ1NZqWc1I6RbibWBTOC6pxwblrOBUE6+Kj
PSa8yQvam6grO34uSwEQ48EM4qTE7ckmxW2RiWPThzyGDgl3ddzUrERTp+WUtYu2
tmuffXADmMPnjE4PWlCbPni8m55WMJ6Gq+SSji1zvnsMBEjVKxT5WSvIA8q0+1d5
kBy5t6FngVhguQOmMU1dTb0tDFnkyWGyLVdGr1ZraF/LZAkQt0JJuKlRrq3pqSTo
ExmYVIa68Ns+eJSINB6lQrcmLrChQkwWhfGQXfNgoCIiX5sJ48RynQypBfjXi48g
jKOWCxfrXbqnWj3bttFdu+5r9st+qLO2dNhPdXSz+0c1JOmrKQLUFMC+rHy2gGZa
HOEhUaFAVmsS2dpB0CNO24yL+En755ptCTqcbha1ppTp62M7BPGEMQtnYih7E8A9
+VDCQs3ifLOJ+2ZzOVlNZz8CPRViCkxhCvnjHuSVwaOwcCiBRgplVDwgW3Ok7RoY
gGj67ISK/Ew8YuGy+iTIB1yxaY+HzJffHjZzVJGBaE3kY0DzqvGVCYDt5MvVLIic
N6/Jl5UV7o+Bgdmmovau4QwWrf+MBbUahiq8hdptPnX69E48JzuAsIZIP2SrTNJr
RkMW+waQzv3rkXMK/3f1AjcMB7CwvrbkComxOoZAAg4D1N3CJaszd/enGLlD358h
wluwitk7HoNG9hCWJDLxwXLiPr1NomlGFVliQ2pzUiAoT49qxrzQxupSA3QnrGi1
WjP4REuRN/wgXHpUJha10B0V+304fVnbcVjcCp3D9qoQSazc8IqDBx0lyXXEbBMg
/dM3V2qfoGDY104gizARyGNDTgtkKGpkHgitPq0GH7mMr28KhPp6uwJmqeQpv+Wz
NEtqU2LM7Z+RAEMoN8gkN0ll/pjdX7HXgEnd6ucEVksHRWTbfFxs0h+ARLzitAS3
Y+RHh/SkQEs7trDu8i68YrMi80aNuNj1jCkej5TeriZ0mfHzeF7Pr3ji4wLYz1ZY
S1UEoiX+EPgWR6hAvA3cQ2jN1CEXg0F2hLN9NNICEdCTqFvqU1/+XrmKrXwM0TZS
/l4xcP00hrR6tdb5CEoDd784rKAGoHOWxhdc885JRakAT7mJsum70D61gFCI0wcg
uGWYWId572G72Rk67OX6C4WNVhOulJ4TmHaOAsSu/9DK2MP+eM9KppW4R7U0Yz6g
JoHLwcgrn7KobX4/4+xylRNOqJqYPqqNyvE0bGsF2c7JPHCg9Sr7TOfzcyj/K6xh
6hF/++xqu727vmGlF4tlskiP0X2YODjk1PlwbKLZuJigzTnTxD5Yka+ZJdGzMu7x
V3iHMds/Qz0Snj1xZcQzcLYXAYLUDqOsfnMbUG5dsxz4DkRIJ2kB6bQC3cks6ZyX
gWBaJ2iZUxkwABXpTX9WxPoRayHSd0jWAhdRaeGuJjqG5MjrriDRaMuttOj4ZLcS
nQhO61e4ZTtfWx36TBmHUbTdzAdbJlE+xc1KrgxvuWCUkedSP40cNHuMGamw5Nsb
+Nc+NurO8vZ4vHe4ji2ErIWjAqTkrGuR1xMGi6aX6AsU/E3PSpKxuod1fuKQJ57F
vURdup6XsWvOi6osPmqyNt6p61lqluY4Wm/TW8dQl453ZAjR46i7OPDLANOIqcz0
8Lbf5MfL1zcLb5AyR0a5bkF7wAnOKCF/KipUkBH7m8+6IiDYNgQhsh8DK3Hl38B8
XYorp4+QE6XbW54RT4nRTZzuCmLrerFmErU9bU0S2iAeGoRi/RgWBJmKIXXprVN1
GPUbNIjvtwlsjhIcSCaTbrO3l0aZauzRT3rfUozQ3RYgZ10J6GlUcniNLXGi4u1B
6Kc0OwC7KguVqsopWgzPxNrzJPuo2KNme2dttyaQLlqwIcPKAkWlZgcMkGtILeBT
kQ8cO0MzZhMCAX9aQvhcDkvwr9WZSM5oIr8Qp6v5phjyc4YZJmERzH++0DcM2mrp
33wf++ocWebhm9tb3vbSOktjA6AJOsVX5C93f1eOuFfmXxzJSW63YuKhNqoBfNh7
51SgdJUFCJW3+Hers+lhlDN5AMtmT3OwdkoqY5RXg/FC60y15GMnNPd1NaW8Onqi
FebTGt3iiSzCkALfQMd3ZsL5byFhaucWIh8rrJtqCi40QBTuKoZXuI58d3R0xTk7
Gd8DSMoCbOu0qmCiLgiRSWNIy6d9d5FAOXMtDa9xoPrD6gjE7Y9hHxDwodtsDDPe
95FZF7qD77W1o1kI8lCFETkVrrFOcpUXWjY3mrxMG7AfTD4tsmyhHyq4cfJcYGMj
Ic7zwOhtjaoEqUoDX/Htm9hWP3xJjqC4vYNk0mwfYJAleCK9WAOiC0Ix4ccrTHuZ
Nya2Jw4EXl7pRJefjwsZoYZP9/iX9YsKr1uTYQSIIYWRq5jfXlM3DyfilqhOAqGS
4X5kbL9GoU/EJ39WHNhT1HvHHenMA2QBwWkGCBdEcKI4GbuH40OBn0nCrzROQwA6
LcrDI2G9tKQ5d84X9ePl/2EBJxykbF3lUV27GbyZY9vFaFvXTGfsZ8YKE85dJnmn
rtS+3MI6s6U2tA/8nvmn6DE0TFRJUKtFuBdp5YAzB0/JiO/nXDGn6s7CdSloPNAO
EWfHNQMUcLBs2hLI489aCZz4ZBzOcJneZEYCAqAcxOTSKasxU4Flc8rmQkzfPxB+
nLaW5C5sAugWsrZId42tNxsrH2bxBSxfBufXwxhf0UHd8P0tXZQ1YZrujKVQGNlv
oMFJksWevT97QXDhgl5BMhOE+ZZAxG/UZnk/KG/+gcztutbLof6tnPTx/40xYegW
0WD6bemxUSXOM6DpQU8EKHvxN1GgplCJyjiOYXujvWJ1UX9z4XHiMNscAZhv+VMB
A8zOm6DQ2tq7hZIsuSz7QRZvfildeQF6flQIDOD7d+WPfpuTfU2LU8dqpewL1zuC
eWCvhr2iXsyAfPf7QZdFDB1znQXPRVpQ690tMwRYZEME3JEH6i4afFVQatRQl4XI
atZEz/DWdsYD96mPe0Xt0wiOYEJWeDdCNoOCNEAX49ZBQaoOYRtmw/ld5Gf6STd7
L+S1B8vf1EjVpMfFby3FjepVm4eBdt3ky4kCXPtQy9Skdl4bORdEfjHZlA00xtm9
UJaPAUqJmw3yeKK6TTKwpNaAgyMYbtVtZ25BuW1+Y2moNbDvv82ouNwIePethqo/
7DfMsrf/QHasZE8oyLmSPtIL3E4TY2l1BFfWxLNeZ8woXHLcNrjYKgkPraj9j4Lj
JYwFbDiDisfhk3QaLAfofmC2Kw0rZifsNN49T5iIIlVPaBm0zFSfiEq8RlKBIPPn
roxvjXWtSMRuwJSGKTjmDgPJyfnDZEtQwhF7CJkcGucqv24MNHDlfbOYfayhN2Ky
zmnAk0pTuD7QZ0mA9+P6NXfXlQbSQ+vtER4R7jjDOd+SpT/Bd8MfC7EHB6quVKQP
/tOw9hntA4fokLdQ+JYUurYYDdqut4GMhT4WpuSWd0kK+pnATYW0PtMXk1TW2ayS
or4dA3HWlV+MbMRPtv4ckVkmNM7dCDHMtXPFQXZo//RkL/L5sxnx0fhvS1w3EGqr
iD686wvpipmla5lwMsUS2t/ACvxkvtSkObLorbZWb4vgHpiVsSRH+xi0hCXB+4yr
M/IC5baek+aaAssZwrsnn8wJkjwaHolgT/LEIRL11hqo5WsXrcvWcZZRlTgHwR88
+ave0rlHCTkq4MLpMTU70aCziq/MNnt959kawU9o6BpaXLR7or59t6sZSGbcEaKN
lptFMStnKMuegfuKySjXqgQZCu5iwVGm9UCnhTvf+6L/eQSzVm93ur0qMnZDdaXU
puyNLhd2o8EbfVtTgzXUb2RTe5YUEtHdg1+SCuZew4r1NHebiblibM3HHK2Bbr0Y
MBdIRfX4IYbNXCf/lALrx4wIPpTIabPQMJm8F34Zn9JwleDp8cAx1lxpILo2+2MV
rfXSQFbOrqV46uy/cNQfmdSaDvJ4Ae81cJZArpGPtAhrkFKGeA0VfB/AyoM1nHYh
dO+5VT1ZQw7D5Ycf5ZENNalHj8suoG9nQtlcu6v7uWYykalz1AcUOf3kMRDEQ8OV
rDahF1QPkc96bodtAHd5vogHwrJL2hZ/YoPXAQvYks1Y5Uvo5EzBW+xj3ofrEFTK
4egXwIewWEQ1+zuGuHDmiw9bBfKb2irJYRC0PVO64CuWwFw51bhNoujAed5lDYmE
UBad+CjusVgyBYeAmCYpKkhoNksrE/4S49DkFoq7e9NZ+EbUXxhAS2tbuCRgy3dC
lK6KbcgbgJL76pgasnqnQTDH86U7ox/dF/JL/4s9p7riOl9dt6O+HhIPPNQNczxY
HLLUu2inXDtjjD/kBvR+49+pffXH4B5+hUmY4WRaZWt94hgk5nAnekBv+Y+s/f8i
MpVXKQQvTxFI2IAqpMsgtR/Mu+m7lZwIMRkrlVu2iYZI6qIvB4GhFbemnEXLo2U4
X9F4BDlnoWmsVtEEBHKG/lM87BLFns7Yk8sONUnl76USCdycpmn/11ZmeJ+c6TRN
25s1/sk5WRoBMCsN4xvhuX+SqUwpp4ubt5pyWgmzVSz7B/WEjVum52LI5tGeTWin
MjaDyn9VpwcZYuCnrRI2Rs3oEKlK2IJIup1IQGj13etbAA7UfQpffW0NiGHNeH/x
bHvMkvOX/3PTtrW6lVEnP9LTakkWkajaJ0iF6s8hj4O6IZAJ2P8NlAVB6mHUGEhA
cHmKVdj+N406UxqqvWAAJHm+fmulS9qfZFSDH8erVzNC7h4k1aOzmgypkGGgHTSy
2pciVSe643cWnQjpd3J8Eb+xD9fSP3TyYLTBmMwJMTFOrjOavXrH/v32W7wo9l1E
nak9x21g9ncOEPofV3Q/WDLWwko4ojmWvKG7yMwz8/heXGsG9SwOaHU9aUYWyfhJ
C90iv9ULKjHG56GuZ4zqnMk76qEnhetJVUkmA21aTn9+T3UlMz42YfwkRM9EKEk1
wzP0tLBB+qOkTki1Agv9KfN0sJvZREMzH065s4FHg0mWGdLfndr/LatV5sFBNBmN
xZ2jQgfS/kTWiPC4pUdMTFcgauedpKb77ngDy9fYkf9OAzBUZJN6j94jfW0pYahi
7AYJqor2YEOJP4kk5e4mc+4SdR0OErmhccFdVC6N6075kr01IMo60z+GATxvugcl
WKwga31/3p3R7YNZwl/q0uyUjo3NpSLVrIgRX8U+DkD+bsgFQ9la2d5jnsqmzCpO
89bFMP0ZMNsdq7W2++fIwwOjbYGj4jFMku1TaQtiPeYCTv6hLZDA5hAB/8cD/O4y
BrBQH+tw6dAyzucsbhKZL64duNOcTLHnduX3KE8X2qzBnJ2JrUeg8NP20XneOwBa
fNbSfpJZ7oYb8sd23x7DtQ4vt2Lkbxv8HRSXsIdT3p96NFTAi4hIAuMqEGxm/LA9
30woHhjpv26arWCl+jtqKx1W4eCSfb5egIaFJbl66M0cjXYHqoosX2ew71XxF94K
EDOW/iJF3KcE8zzzYeolCuca1B5xj1j9KdDqN2kWTp2mWnns5RXpajX27jMsyGRY
B9WxPpBVVQQaCkHGCsnuya863XY8egkDyokH9M2ZmNAGGVPiAl/rADLCyU1TmzGg
sgZUiCnTsiRQeS4NE4jEsTXCc60dHW5RJbRYVreumGFuTWVIYX/49U/24XMEUDog
0M3zUOjd38aYzOjZ8gwjOFd9GQXsUUi9m9f8yWMZ8VrpQgpIUnDPrYKOqh0BjvIm
ef32p7wXryXwUSzW3ljv1INk7AKO2zZxBYB/tPnkLvjuGzGbTx+a+B5hR094T/3e
3GpjzCi4mTGONWXb/cAxbFnqaecJwzI6IHFYuTM1jg3gfdgoFTV+m75c7jxrrKC2
gfLoZigKrJg/AF4iwwuZutdiQDJcLQR+nd5g+NoIlFoTwOCBqVfSoMdJ4ra6Qi56
70NBtYtfMcbgKRDGC9UISE6Vn5qUAjiHPp17dDTB8LmDFijEgaRWKFkDphAgWRee
POKQ5nKlkSJ/DczKPMVUJzzG9aoMBAsXasdlVGeQU7krV7gChJczc2kayTrpczRP
Aw2Pw9R3KT9e3f6JRBvKrkx22s0JSm8OKRcD7Rp62R7wqcsvvyEpiFgEc/rAk2E0
3AdyLOrhmvU95aSUrK0f9MZheFwVw7nylB5mEAfjaMj2O75UpKNb5OcBpsENHdAx
OjnfceUlek/sc/q09sBxvFu0JFOAQapWN0WmBzQM6nXqBkvpGEK+9SXZyks/wZsm
TiIGBOk5faM/fl9Qn9jHZzo6c9HgRWLWQcmQZLwPSsDb+5HYPHUvP3ERh/dND/Fh
nkcrSzCG4CXKO6phBbBG988A3zIMMpVp9Lwkd1/w9H/d1LYem11K3BPukJsBE3T2
wdRvK7zyY4UrOPzz4IMmHQpkQ37rDL7lDHeLeRHyYCT1d9UR6bFzLsuU0HdMNxjm
b0aSPeeyacMGTR+ykXWoA9bCy/fV5ra5SyOo5BREJrQ5xtagtt6rRcur16oK5YjW
ebj3XVRt0OcOx2aZKz1EUXxAJio37wMTT4S0B0i+zpgLqCqmIqrxo7NnoRju9D4Z
pUEFnDOaiu3V4KgLwgbzOojArsVZqvjgMm0CVEMODty++7UuxCp2rkGqbtbZOYzd
d5i1YGjQnp/PX7Sf07OHQFm2/ebCfR1F7f4My0ETJIxJN9VQwWZeWWRlXOu2wxKO
ySFzbvUpf60drD6ZQ1lfABQg88cE+ZEjj27skY+klJb6r8fT0wkqZmesNCvlx8rs
GvrLAZsKgwMQwiP5MA/ORIGHRcCQ4WB7ST3KsCkZMrDHTN8QsIZjS1wZmaI2T52E
lo+z7QOV6YQdMjuWQXjl53gGBBZmeZJXpResa2ecaJdELXtxmqPUrDMFfUsd4EDi
FVFaIcwjF1IlJBgIbAvqMxZK0L0YSlGqs+RiKbzpq6C30vSaKtHvjyyrkJxtCQ7O
G7XF/YBKDNubLu6wd2shwH2kE9sBEAuzD635OmjZYU1XhLXmSrN5IscLGaeFpKDg
zRsQXMU1x0UP0jthQ9nYrgC/x0gBdv2cbh05KDGPMfp6wefOTzrJs/zGnP6HL0pU
hTKtF9gFlsrvlTGall3hU/00Tk8l95RGNmx5UCAHCuI8RtVxclJY1+HXtGXVJHYd
t4VWxpjyTLTrLGYksGfVP9+qIp7vevZpNvLzZi0aWtd1nag7kAsnGhEUF8hgHpsP
+GXCDJ6ECwC5i8m2w+9hqS0d5ot5/8/eZy2TqcX+b4koG4lXsGPxAQqC5JzHf/ZJ
bbyob5/Gjt5nRKtH0grPuneIyT2JwXjjVNK8+pLJUHaWFm7Acoc+UaRGO3xNaymf
f66vUUBymVIt7AAwP7F6rmJdL5wo3JVdy4LK5lXS4hslJFkyMaVoId4ydo+TmhB4
dGQOQyVF77635eQcIb0Vh1gGtEZTNDGMymfPeBCT7onEPNPaaki56ZIS/WDdO9Ej
vYRHMTbrzDqlxzSlkwdLKFyOCUpQFcDKDQASQ0Pmr+uq7qoCHW/kyvmvc4Syyp9j
aLoIt4z/oCGXwgw56fxO+sLxDWVnfY4TQQPk36G+Zj3J3zSsKZi0iDICIr9dS4Sl
Bk6iMGlI8zhgQFvyXpcWf9qeMIHxa4bwPe4siZFmTvggh9nE99ivylov+hpcNHPB
/GoZwTSDH8Slv+g/+BT05GyEvexlSX0Nwy5NV0V/GIydGKkZLEG+dTi2B+T6sP73
gaOnGZ++E4kfk4MxCZEVZeMRt7M3z6NE0Zwgi5ZaWbhUZXLpb00FxJlVq/oUYENB
ztrX/J5scK+US5X7y6JcJLRG6PmNUv/uqhWx8n10l056cP6OiL9JxDNTwIm8wwVY
zWJnBSKmsD+aIoTtaNuAwOM9Aw6y+8wEOnD/hO+O48KxLXDw3neSh79TDAhYtJ5p
tSsAtiuKrAueLCAsaeazou2tCCtF8klF1fIghxFlzg5BSPrVIhR0IMrDI2eq6ccc
5Jql88Eh2ygraKaWzR8u1JNpwLLTnQQqvt8FiVAQIrIu5e4ytUV5jDv053Wm7P7N
W9Qw9MozXgTu6hhCQEloaj2UZTHSA/WoDedbI/KAjM6plo/8WjJ2Z2XKEBwGBB66
37IUgRxISmyK46Nsoyk5fLTWYZ117e3GWeSMrPt143LjdF/hRB2PpeSyq7wpEZmv
hL+FTuX0z6r8isMVPGedXR1agdO4kvJHfpmByO9C+89vJTViep9NCU3gcODRE6LS
1vFk2FuUmL73EaXrFpoWFkWIG0GSFCVEJ+cMZSE1dIMQUJJwKFs2hphte4DfBE9A
uNIrAqQFxmZLS/VIcNK3TtGOIAlw6FbwKo78pYXOCsvdB0AfGgWE+fxpBTgzLHF+
rWGDkaVSfj1ktfCIXjFMqHh3O1LpIX6OpytUMh+By2SU6FtPYtg0qD19YDt6vri0
gW+QgYHuZF3fRO/If+ZiahAmM9yPWY+AySROfkfUXB16X6CIZUpsAh7VL8w9gpFm
3M9N10j8FxLPT2JPepjnk2AtqrPklPusGMt595GQocEVWsNrBB0VsTvPbuqCR+3x
xyzogs4ra6XD8u7QvLXwvGuoH+CnWxSwqZtFzZCUTqfdr7x8h0oumXAXnym3+zOI
k5cFQf/jSEfYvoENYcNtRhBGpf03ZEAI2HMBnpJAirBkx/5sC5wIzQL7WhYuewUW
y+B0fhiDripgaC4HIo4GZCKE5v1aqZWJLZcfSDrrF9ing80xn7lHvYDqc7oIgOji
UomeCzWRzpeDz3oo5uWQkVCYjL3sszgEoANrAGzKG+NyVgzYianDGsfg6qcs7N2o
c9GzkRvxWn49oBTYNB0Ynvjj+ZWeh12yrWBdvlzC9gognVbSFSDGaIzee89mtXyX
3InIWQBC3D0/MgWzKjdK0ZZREPxVRCy5c63iwu7JohqbOne9feJO5APE7Gv7Pjcd
xTeLPLuZxlRrmV79UJVwJQqfwVI9HRfTr3nSwfpXw8K21tYd41iuv6uo0mi237hn
ujck6pyJwh4ieCf9IEIvvJzXkX2u+JhKZrwQeqL4xeZF7pn4G+clTqEBxDirh2KG
zFz88XHvT+vqb5z9wAqZ83ZU9ENf2m99LmctyGDAC6uakSmpz3PsCh95zQarKxP+
wwY6T7paVsUsx9aGG2l+hQgCTmj5TiDSTD9HLuZYZYokvXuQgBUyXvjxgcdyw23q
Wed+IRt/xDi96Rt/5zvCF/xArejnrA9xU7DfACzRdwQX9Sn7nf6fRliF4RRWQ/IT
tUBPWwr3ErFJhj5ZwgLL0ilFDUXR//OzjQPcWpjErxxyK4EaomB1MOnhVqzwXMeo
nZVkEwhBiDLyjmxGP257kKfOLs8yQVx5NVATEcpI33vi94aiTh3WvAh2X1XMBMKi
Z/YwBZF0k+Hh2kCx+bAOWJB9mhEkOq0WLna0xQFpvuowSpOHV+6mMHHr6c1qWBcf
+0hKI1WlVQEzErlGq0njKMQAETcVwTXHObSZzxFDvN1AGvmnLyKDpyM+hWY1qFrX
YCXW1sBXpzT/m4sphbIf3ga2zHjl1QECBFK6Dmp+9dNxaJl7kE4XmkEPiLZVd7+v
jG/sbTVQNI2G3icd5SSVjvshoQ91NajkEA7hJxO52LRlJutYsolRMT6Ss7pZF94y
BeHy57RLMTEZrk/Fscjc02duXPmncCs1AceQzH6nwnSMhk2+ybfUrAobC5H4Cysh
+cqgsS5nHSPNvNNLwsYdH0ZZgB9uvF/A5CUCre3j8SyuTdO5FiFCZMM0A854m1Y0
z55VHEHltWjmlsSIrl8U5OxaxY8PMG1T6XdrZ+ps2rGSEA9LR1/LdSA9uez4H9fB
pW0aj8dh7dKJ0lY7t0umyvB6Gfq4XuAG1WrxPSi7du7F/XJNuo42LtwilVFxhl44
mvYdM1h1pxPy5ayAB/QZ+dyM3FOy0ETKtCvU6S/g/pWxEeFqG1KRv5WjJbRgwqnq
jZFPGy0Q9j/CeixTIgoIQWz4CHNipH8i2wBb3mvgzQVOtYCfnD2FDjPjI6+gjWIj
P/U8lUx3JaeiVjR0rWKs5NX37hygoJepxn2MuYzM3zujBxEqypM7Po0fW+fqkEjn
q03lJmCLVPwrWC5diMpIcnG3UdcSdQzCr2SDhhyVda6LSHm4XWbP1fSMPHQeKaP5
G8PYvdFVQhsYf5Nb1iM80og6DbT0g63QXe7uPNCUllk+PLQzdYGQBeiMRKtPpsN1
KEmW+AHj/Y9nov1QqEFi9DeC1wBtVnsDRzC68t5ByDXcf1XVt/3votFi0k7HucVL
4vQB1UKnWEA3HdzwL3fLfmi/Ly3izGkiafkxoBA/RSZf1/xhXowOCHcyt3wtdpyu
OtaNriUvYat6eXrIEZCY7mJEvLXsKW3WlXvnsd2xG/87+feowujtQiHY/DZpK1J1
CzcOH5jICTcJa7xchBjKueUZ52YY7dz1a82uX1VjZYw0k6pJBpN2NzeQ9QveO/jv
N/Hb539i6wK6karsQVqQUyw3W/z1Pdsg3MNmnD22X3NV4a/ZkkcAhETq/J+4ohHq
VJSqXOgmjqcfhlBlyURgd8VtTapLTjX5bkMR+LF2paRYJnn1Pe4CDy5JZzjCKVEF
2wxTfKxmE9/cn7jo2iyl/FtrlYzYEdCxkLCkFWiNE1Su5G7KVzgO3punRjcpv5p8
+OJ65OJZSFq8ufDvEmKE3eSxywOsdIuLsGGNGEpkr4u4/krfyBus5eGykY0gylIi
O6Sv9KQftnmkocvRIrw1UG31W0C9nQPzafX8kAwaeHthdeEC7EaINTrpBOoUiGQz
uYbVGP9yj01v0G56fCCVsXPum64VLL9wm5hblq4JFbWA7YGmo1YlEPESPnP2waXV
3UiePS6nmw0m5tuYuIMO1YvAO1Hc86P3P2pSmEPJeLdOj2LNz2daUDaYfs+RIeqR
GwSsrUww3/qi3PV/OTTEXSvEKeHMF5MQ4gjiAvzaVi+ha5l/kxFozXhMFSb0IUar
eFHFrKhDWpMhkhRrNqKL0FS7Q3+P+mSapk6xoS5AYPxmmqyi8fi56+mx5GA20+bo
aqsbdZFDKf14rmiru88/Mzr7t9lw3mBshoRc314nsi3PXxxiPknv/MCJZ7Yp3s0k
Z23XkH6bwKY/yJHWzRhdGzbJ2LCDSMQmSfwfQf9WQkAmAc+6audd8wzqqZMfsLr/
CpZXOs4WL75TYwlMPpw/D+Zxe1TnGUSf0q0+5fu5ZWA0MdedOxfqB0TPp/G74DlS
yfH0fGyLJzvNfEIEzp8Wnvx9M3dnV3m25HKKZJH29oN2mdyiC2GMgN3W6IJCi9bC
ojCK8ettDGZYQ1peSDp2/MHJDw1CF8fp1XO7qDicmgrxCsyJudEeGcmtpUxKhHQy
mCUjTJFGqXUuDWIaTHxuAj4TkDd+oF9FHW4pFjA+rTqJuX8w4/QEK7ieC6q/HnEj
fe6VeT/ykkumyDcAJAPLDnaEG/XsvUnHG1rydL73eFoQgk0HPLuiseMqAHrtNHpm
0hF0bMWRKp0Q1f2XnRrvC3B7lzH1toRpuozRoXuiEF7ESxMbg054b91rooauXCGm
rTnac/7ypgJf9sRd/C7Z+8dmQMZbFnCDDAjA2crZODxGaCp7pOJeWLDb8egCGfTv
5zx8VA5b96a0T/mopt3HV5VMBVmx/ieoVTRSCTxH7UtwFKT1OPm7mGdnqpmlUb3K
YtK+NgPSCw3tcr9qisobl3aLPwz17yMqf+9XsXhxtAyn9BHJbpzvrUgXXZZnKU4E
1agtojpTWIv/8Ngs6JWsUxRYBIMg+Ku62BySbAKUnXbHNzqkSlHrdOvBHnDeuZvq
fEhTyuiI7axTEJ/E6wKFItO8v6GV4UgRCNHT9VbN56iEulemUcmgVOxYbburSl1m
F1Wg5XdVBctpL8rG7X0G8ljhmtOtLMzkAY2B+2715i17KDgb3OnQ5i8myiRqhfFy
Np9xUQePrlQgoOaHnNHoHeRj/7f+lqd/mK5fQjeHZKX6BH56Go6+LYTi27uGnImA
+7EdFzeE6QHzUZmt6YVu5JqdEGsvm3EZHkI8tUxhpPf+5MskinEEsJJ5rpTmDIBy
jyUCb6jBqDybZ48RiWC/4wTIFL1qwu2AsLvRmH7X27XOCOBbDR2YU/FtmQhYmIuE
DGzCYKSnhoZuzTTt3FvKt+C1I0eg4Vea9iMb7KXj1wFm3r7XBpyYinwANQTUxP1S
T8+XkENyI1S619UrNK/zcbVjVhCKYzPW1E8ALZsgdi+RlCUptfQOPw+cI6dDoDm3
V1f2T5VSaeSDTZjdaIU9gcUzcNsLYVPAAxqrIGt6Hn3PZ5q+q4DmcFMAp+Xpz5l+
3PUKBsYB8DrOpXoO0vaInyVAJ4DKSnfvvrmhBBhTQ2GWXo6zu3FyJzYYnLhVZI5y
r3ptQcuU2mj8UAHQBbeHXAneEeD92dd1aBWShQIouOONKnU3l1C5N/NfMMiI3UcM
9f0ZuQ44HtNYtB1Wz7TQ/LYmaR91c8xb7r/Q+Zr40SK3BpY1VHdSwf3yEs6ORkBj
fHVAF3UDli5xykn/iWetD9YB62oAb8zrnW4S5M3SSNlVc123GE4bQsrUyxGo2zjQ
MKBHZZP/OqevLopxNacl0jM0JYagYaet9G7KB+VabS54rK1vsekvo9LFZqhEGNTG
V3gAeJuDkzCkH7ksy65lpZXxiEJOTxQnctyIY8xw0BUqJ3KEkA8IhOjkcw+eDVuL
r2xuQNdBDkDf6bqS0f1hXyam9V6HS0jowB1sDeJPfJeoaOxklXYhFVHZcomWeH9y
c46i3qwRHARZrDuACE8c7AeYV3BZcSNbaEjhJt1rlZFMtOkoCkRlgRWWxDPybhc3
+2uL2PBRio11udJuPMppF7S4pvC3MRVM6P9Ia2WtMc59Ot7JGV3CegkQykYhcsci
pNiHrQDOh3eSyaakseSWMiDIYimiJHqHKtkXbDNneRqgndZcloK+O3/Ee4xINqmQ
eVU77IcRK1F7XMNrSSIUxyX2O+IyMNDgBZIqDi5/53tzJuailHA1VxuxqnGzrKfl
U7dpPXJAf6SYuU/YXnb2gddefWaimNj4P3RcrFKby1iWfE+P8rC90y0co677bN57
YuOkTUD0qa3Hotu1sodtd/FXVat7ZDImgsDGb1NiD7XA1WG0yQVwpN/C0coRYvFO
9OFqwUpwLZyuy6EmzGARopujkUajZ+gqn0AwqMyKPPHc+keRgFDbR3uqchOc9EQH
KGe1oTKtOHpOClZrOIFN9espLdwlcADnXsjXK8YYBuLdx0Ri+tIZOLttgkaGL51f
06LVnwLcRnxp5LjoIuUHv3nhSkdUhveX6prfjYZS2yPsMZcCqXWvyBP2KSauqhXw
neS/pLUCAHJd5SuabYAxkqdzDz1ujwqaiQI+8sIAHsJv7XPydoUYFjaeiAuJQHIo
Z7uVtlfii5b4h7O/jZstSms2/4by3XtAAEKfcM+/CyzSbGfMPmTGeneBHC/KT1nc
RnLFdhv4iaZPjSAXzN7JLZK6Vqj+7J80Po46T74CJJ5MOE8Kr5o3VKYeJX8bZamW
lKZcZQJlLsWKgc+xVOVK9pxmZWkdXzXJemKYVjI1mjxVrAsImfnKYB32HuzncZNT
bAR+CPguQRQBJ9M1MCdMUF1YVn6bzM+c3qe62qL3agwfqlXI/JK6nYP7Zk1q/MDm
ZazHmmAGLfTa5rYejVU4YTFyFD2SODJFWp9r+pgfEnXvTwZ8oJ2rHmtSVGQZILrN
T6AEvUIA6FYSKTdDM13LK4n2IIBkcHudZDC06jquzIzSAc13nbjTIcDcbQnoBj5N
T01GZICvG8T6sRL07/cLnj8TNWnL/da2iuC6GdkEy/x/r5bfK+xj+g7CGwfb6bcR
jE6OOHrAG+P/YMG+SxmDqNwmnoPXs2MnvS6sHW7A6DLR2CdBw449/sfTKUmP9W4r
PfpcDeL0b9zRPTVFoPumy/jmDDs9yXqDH5n3sdh8/8xcmY8QBLwn7Htc689j1KwY
9dXpNRvKpioUbc2eTwt7msSp8Eg0Vg92sJSUug1+fo3c4UEtbTm+XbT0h1TC41dK
Zny8CWkEG6KemCZtJyu+8OjJMqC1RjFJDByAcwqVWckLYNKpoRjX+CnACDgRto1N
2eJ5/+AUyYjAauClWmZ+MXk3hfwl/sVtNPEjgUc+BKh6ZnLNM4J/1ivAtW+gh909
Fo6aY2l2saPSLJyg0YW+K9PX2dFERegnb7hRbbXAXkRYDMbhgWsqxKFVD9BA4cjB
72e64d/zPQRFnKRxa+DkFCC1FjlftI6JZ3X2O1B+xyT4wFO7uTpbcfGI8JjGBuQe
BMyGRbfwTAh7VmlYcevsq5zB3BNyPjpc71PTMfH+7+VKGbk+GmaEwbZB3gtmkr9b
8VwGxT/w4MidjuOkRF8mBHrCJ3N0jdKl5xZDiJFx/K74skIAhMi3DiZF5TxgOMWY
/QGKBA4UW1ldSeU7U/4kvcPLP3Rxh2le7YFUv4US6SY6ncyXFHNPySu6x908+FVN
kXdkmBTbWx+B6o2woMi61pmKJm2vhMX99ZjF8zFXDPvrpTsubOH3kkXFfWGjvn5d
rKaXyoQvtlmJnKJA+a4njRz9WdRy2A0feF4QFgMgv7yfuIHAVDfxrljw8yZlDdgm
2pEcVc2zY9gRP75YVTxO1/AP800ej1sZ8hpCjigOiriY8MmHu6Wbxj6yLgUGcKQ5
tb3p70rGP6KBOdTKOZnVpUJbp91v3VCYVSgJ182bS/ED54MWNac3mEoCXykYgPq6
2WnaZWBV9EcSw06sPt9vD3JaHu9K4aACbzC4RrIAXTCQX0pC3ZBcAm0N1C4MwaKl
KzZukfglDgQ8ursnFcEtA6q42GI0Y6WUm7CQ20D2RkQSqTknGjITKzYAjUqu0U4g
Y7SLSJim9HdiQ3GSsWvxww1/X5uJBdLqud3SVPb8druBEUVcjNeM0gi4v9i3owR7
IgOpf1MmByxlWJqFwsllxDxpu9X5Jq3f8Ue5RuAnpwqSs+FydsmKStRYCzDtBqx4
7VT4hCrIDMRIIruX2PhFaYlmNvvvQqdgWL08H33BGaQscp+xoExIrVHu7YSOQdG/
8goI2jkZublrR52xszK5gqwKx+e3Oh2rSgZx3znUk5O2f4nz9WeEbFphJ+4EypQI
woJZw5LoDGnB12WfIlXKuUExHcrO88ut6j2cRjlmXSUPE6gYxe+H2TU54u8pbk+I
SOF8qkXE3xhcBMwOCPI1w1z0B5Gp1yhie3XhSnLkhXxlOiEcc80jaJgO/n09TdHR
7Qs9nFsfHyVI6kd6mswfyz+P1xyDxn9L+aAAwSQsXGV7KR4bvLxyYhZ/n7187+h0
hfGiqbqvdF788KntYw0anguUwNQeaOKRwc8EvtpzAoaVWwx389+TC731f0J7wjMU
ZCjwDPm3yjaSEpGPvXNw1SVtIwuKtAmY/I38wQbH9iZXwk5z9k42JTeZUkDqWwiX
kPclVsieA4XUD+cDeULhpsBL2t4aafLHUQzcbQBcsuC7UF2uJRTlyMbyN6fX8gW6
6spgjDcW1O83Hhhh6W/K5oylldWFf6cUcNJyYzbUA2CFp0W2ShrQVypsWMnODCQk
Fv5rnpMR/DbzvMF/gpVqHgtfmsfYSDP2jKqJNToQfe24NrC7OIT7fHEntstkgWKC
fWcgE9wvSa9nvRu7PVaMoLcJ0Z8RuvWaHn+BYT15fcLYKxRG3P26ahJZcPIquV25
mU8O9TJe8t8jdKa65rjZRxjYNOVhb0oVhrKbVT2aMGfuMX8by57Ea9YAFJ0/oUcd
EjvWHwYO8Uo4083yIgE5FJ7FfjsbjHlvinWniB/Shc721qL936ZFyHaVc190wLe+
yZWggMvHwmI7A1xBkFt7RDWR2sK1HdqoRCnnZViZzn4UYEhr4s2Et45PZVvMDAmp
FpFpP2IyGEES6q78oTX9CcGhEDWS7SD7ENR1xIVczw9ams3aWFon/6qTz4SOrU0h
vLNL9C7oPvQXvtMqW8ctf5SOjTiFFPdVFWIQbzrJfvjV0W2shhsbzvv0eetZS1GE
KbWE4RlU+L9GpzosUJy1hSEU9XUjXB5tZWN6+dzNHg7RtlKlaBipOWEDg6w7yktV
/M1Bj9CjdXQJBzzh0TOJvV3hEaetlGkB97jEqXV7Ml0H4sbAXH0GOOnjK1Nz39jU
XW3NYQjhi/f2gdOQ3e8MNJX9/30xwneyvffP7DdrYdL2fxN0FwPG7LSm/3BOx3js
fGxpwfY32bss3Q6Zf7ecweAxTbijNbAcms7sTNwgp3RRePvP1g6rYiMBaTl0hxCJ
3qn49ylCOTiR6lR/fyaE1Bq8X7WzPEZdGYnIMV6eQK/6D8JxXHkDQkIY0FMQBBDc
BN+KVyoKzRrhlTTYKhpx1S4/jHZzRX7S+6cA1qYubkIUsOv0/trvfgBY2IbRrp1/
O3r4GKL1wjLFz134cVZE/Gsh/5VPzqehIvPbqhUwMY8UgCXY0FMpdDUKH02qBtaS
XibJk9axjUpYBUmcKxZTYq8QFzaLp3G7/LofVylr5Ym1RCLhSzhP3gbjbTQeEPkC
g5p32AXoSZ3lFNQdmVq9sI42/j6VCkUQlbOiX1RCfCWrAUquWROqcn6D5Wnwm/BX
4l+9o5fx++AZM5wpDMklnB3G384Fna+PShZZMqAc4yfI0IZivyXNmpBkq79JHg0k
mUfpquc3OXH9mERoZyN2ftaSzphSEXfcOsb1aMpy0S9C+AjszSLk1VatN2l+T0Ra
1pl0FvWDaBnsFf5rjFvFr61xkzbXUfT4IsNhBGFS7T0jvjvHRWU7qUu2qMW6gpcb
QCi+uYHR5Rnd9W3FCJXbQ5jTgVdKZ54z4Bvj3N/nWjQUK4BA9FD4EucbC1MmuvWl
1SicGtPtiyW7CF3tdC6tBuxkz3I+S74zBuOpSN6wMSPVD2H/BfhdbxHynIFtOEiu
GUeP8VHbPs5JtSHNtPHRbujOAl/0MWExtRK0L4+Ke0GXomIdfxkbP0A0ovKCxBGE
Vjxfdbw565KgtVmW3q+5SJjUY6pKiXHG27i0lq2LbMIREHPlFtlydPlRDNUFJFQP
RYrRuWDVorFSpr/w/E4Pa74IEc6W2AcSbpeTMYUjoPu8Mj7HXO3K9f6LgviIlXad
+brF5aTyN99TPjy6SuhiXDiswTgyMPKAIiIqunyJuSWaSISsuwFiGH8+2FLfijj7
dbN4BcByqT3QqVqUZxe6wnQIhWh+/3UJQigetueCFA/52n8n8AS6dfPw/SoqJYRq
x8PavoL9FOuVnF8IfNErAazvpyIb41DnHaTwGdf0ZBvXFFmlA6aUv0qx4Wm01yv4
RDXANHmNYoYLzYosSIZiMVB9155fK3niPO3kxPVCUk7ysWWWtqjqnApM13V48bs3
iV6Kd76F0zTw0Zburup4dVsWQ4jYw+UYI5TM1bBRsiJluh95bjqpTeMKoa8z7sF2
MqNWwRj62vPC7Y7tLuvnP8HPsshgA84YbV0zmpAK6zq/V3pr7bWSjAXL6OUnW4+M
Atm3HI9OiFO1CUw5teoql650Gw2nEct6fpH/VbHuum7slO3KClhQRXMIQromib1b
d+hDmmcf+Z9yH9ulnoWPjpo+e37h2E79v5ALO+viiIBYceJwCJdKO+MRyR5EZcSS
F5KFwMVKOn1IE5ZELEGvWR5J71QmZdwVHwK+SuyaS9J2ChBGRUGuyewHM/phlisa
kCUHEl/WWpFNgOKjmUNEx/Q7HNapM25LNYpeRJInEyzHPoEm5nO+hT9ctqetIes7
UjbBRV7MnZkrJma8tFbhAx9NWbldq9s5DJJeWpxhGv23vb35QXBWoHj1Qk8sW9pA
lHdpxgsWby7rfFb7G2OiiTl75RKEhebVo2RTTP62A0K27L9F8k/fZC6FmVt0tzaR
MRxIAw48qj1Jb0g1z8NJIWM7IENdNG2ielbMOA9Ma/Y20bTeVyTc/ea+4eXD2XBt
eQm2P6+kQ+OSf7u14D4oW39izVv46BqF5U2z7cYw+NXSuzH9ocxUzAG+7QbJywRX
ztvl2rBPlR4gMUWdROuA/yBcrzXjPDyqp5hFhn+VaLM8no/TT7K/8dpsAFlMg2hP
K6siTmd83EqGM78RC5HFS0Y3e+ZeXMgH6Z3bmG7XdF5gm4+eAx8/PmcCQ+mE/5Hd
zM51MBhsJIknm90mxaLEUNy9AwccepQNdt+XIELsYILP72xDniqJ83LPPYxvlFck
4JYyk4kg28eP/yJJdFwjdjDYbmbYKpv7XwvhVED7Y29dxJecQoeza5UnP5eG73+t
Wp1yeELs/o+FpIS37aQDXfcpFS+uNpHAZmbocjhgRuJJjp/oQA4xR/jWBshonFYP
UZPh+ECqigbWm9tRV6/TaJW24a25907VP7ZKcOSV5Smj44Qz55BSD7gw/jfcglXi
najRLajV90/ipgI2NT4FJgS6VDRZ4EBKiXHfbWm9mKZ0noiJOWJ7G6W198XI5WfX
GSi57qQkUbWkIRlKTZeUYywcVlTxfxxzN3Xs1KQI8D1r2Cl9pla2t7kSFd2Wap2w
N1LkirxLOBBPfp8QP8zPTMmgSvIw2hmTKZ86TyTvrnXHCOuCBBfU09x2RaAJp5dx
avvF0Me7Ia1yH57IOzaWgv/BCPDwmtQwXO0GBN7VMl5re8YoYchnSs6/3eGSXqw7
K1Soje+UGFwtcjXNZ/nglByieOrTryv5IwDMeyhDVkFx99kKcIC8DZQbV7a68Kt8
2CXWew9V47M0gA4jv2f2Y6YbLqbuPDuan87G/KLM8LPD9IDm8ScqDsB2QAzoewgC
o8fc4BExU/FFP/Imfa0siV3P0hgzndc68q4qK/d6S3B//ER63qrb9GhTgo1TdarI
MJQLm6daAHKQl6dU/PI7K3xhd0hwrF9htCRqRDr5wR+hcLJmeOfj2pOF5eHyBIOh
mxS0QVuqbt9/9rKAiPoY2/KZ8ASq2amwtxc8g4O9bVo6kDg+P8x7XY9U96oN17/M
x2NIDHDAwsrWkKwRo7+9UpNO+vECTJRhskg/D+CKuzYDb+eV2UYZfbe7fpSeA931
tuNZ86KoGPcv/2QwbImKZsJNWBV2UXNy4VmYqUESn7eHZV081Glg/XCtnAPBHOy/
05b0//kfhP8OukkxlGlyyF58PdegMLhi1dhDpwh8xaJ1HPyj9FlNVSevoTgkQKev
A3sWK2/ev3iiH9WvJh6ETBJwdOCPNO288jZ+AXCnsQUVpqWdCINFvHYic8bB+pi8
1TaDju+jne6fjDwfdd1s78VYrqMcv/taAUGJy5SMqqeEpKSUeHSphnjjACa9R2IH
FyQJxryCbq85VacX4/rH7kJs80b+qJMdWRZEh0yhD0eFLiwUjV3M671LUf4S6SJ6
RX9wKwTkOxzVM+ofzPlerbm+y/JYAZffYv697lL0igTDBaEle+GXShEZ09jeJNU8
XY+qzBqE9OVS1LUOVeP29P0ox9Y2N3kwHT+JYhlG55OQ1FRel7Y/JMXdATkSZIV0
IwyBlbtjwLza5766XH5jCAwWpUZir+9GKlWxd5Tm4tYegSO5lGM1Rd2grqc05/mb
4v1DacFcMgyMJ9j5QR2DpZUdkWNoxeg0w08yyYSvCZl8HLwVgqvMa35fwHYqyuB8
Y1Sep4Sbn9jAw+H648EDcbnGBXrnJ7W30m4jJkYnJqwMJqyRerF40wYgUD4xc2GE
zw6fz4dm+KK+wXKZBUqTkML+5n9iBNm3eHKMk2K8fTU2STY3vng7LelJ3w0Ryw6z
zz5/WP+cEEw1JnNkIergtgwJl2DCjOcXi3zIQRK/q1pbZi+pfiKyQBaWEgOXNAyx
UypHxeLE/OclFskdweiSw36FmYicGrj9tZwTuFX6z+uqLaqEaBDwrWsFDR1t4swi
pi+TN9q2PWyujC5qykE1VhdcnGo8eMPMpV00dazTVxGVktf7FbFfcXoXrJI1SBYl
ShqP5DVw+KfhpdkcjDoqBIetqUI4WKuZMOfk6rAUK32U2ZPaaZtIHeOZaxIC9lt5
4UTemk9BfnRoMFso2z89Duj/kjC8cOnsljwAUw22xI2vM9gjGHoFP1RCeMbXe194
TuDm2bNlNO3MYChXEBAw6BgtJ/itw3J0DiukkBSN+Mf/HePFMlHdwpd8iBbbSvUH
vlVgfZJcjnOJ8R2WpSnescaxacRcZX07YbOW4eSjh81gDANZndcMF4s5r2UgYKzG
Fwgzy98r+T1lXRHKKVGG0ziA4GQYfsRnEKwcc2FsbpXCkqh9jxuxXEW4XLp5+MwC
+EV8tk7fiO/kyf+/qiZx1N07hv3P+S1PlMydsvwsM5L4VZchDvXHpEXV5bx4ab43
LFewc2v121owvUm0X8XSDDvn0zlP+yF5Ae9nmoPFbWvWacDNckzBikq3HE7G7b/z
8ty7iErsOxU7uTPIV7Ze8DhHBwkAMqLn2tpzZDcfpPSETs6wTANoWaVq46dAeVg8
3/p2zNbmTnXlCM7ebBidMRhvkSX5rZa5xGPtzyziI9/SA2r2tgKJKwK1YDO4E+M6
fpbAihSbTcQQ1omECYHRdBUn5ISYLTR4aDESh1zxpgjX9Waj08ha5ddbHEddVajx
kQnqo+WTyaRSQRDdSs96VOHbSSBz/lif4OnYLJJtNlGfKGrnJwU/lert/5wHIJDV
LrFTyCPcaE0OKGJzV4kZCSRs7yv7EixOR+mZLp8bffPRmILXAh4S2x5p7nrPRGG8
7Rsh951jZiWE2dPmXcxGwq8qyGSgFRb/nNEKEK2eYIC8nviIU5zL44429UpJ3e+w
Fu0chyTtQBR22wbMQPF0vomC5qawB9J9MQPysmXdVmne5YVEzDXUIdZKdwZxLDTj
h65veiptrvouRox8qxhfFAu4oymWoGy3EpbU5KP9p74VQMtJm8RH1do9ZLNZkzmz
TJNk6Y4GJ6hPvKbFVzRl5iF8dC2D3UfFuDCr2NSb9Skhdtc8DyqIXMUZRhQt7Ox8
Hr+E4VZZes/lp4rniiSkR4eAP1OzZTGX0HYwhJeW0X0OrlVW6tk7K/oITJ9DdueP
KLK3ILawp8v4I2y0HW9Nki3LT+q1p6KIG/LHdRi96EztnLKDCnx7kNx9BM626A/F
YTqWuMmgn06VnA+vTor5U0E9pTjgJWsoBK9YwkzT8LuxEmTnGs+xpsH2UQFOvPsp
HGDDp0bAXFMlXTP3VgBaw9ojIi/Ln2rbCZawejOn5Y8dHWW2/fHSD+3vJrF6p2O7
R7YpEjyBSbedGEkaRsSPYO6X5iOG+3xruM+TDt5Xs1WevuSh9W/3D/L/UJN9U5S2
Z/gJd7KYaTBR9Rtdg3+/Wun1/ADdLGEm1O/3Uyf/Vc9ivYjgVuTizDZjfUSKGiNu
Slwnkval6gZZmPGNqu8vvmBQKZ7iI3dd2fr+FDb1/wJfJY1UHr77WOZ8l8rIp2V4
rVjFwMzyxkeUjd0IiIlBWjUZeDzhoK2m+2rr9XBIwuxG7qOIga1yP0b0fFU8euwf
kZRaNZex91trO2QpSZmgXhwegQdYazW0K9cDZtdEm2CyKhrVtqERLPM1+R93KbuQ
osXxM5CwFfQIQvi9hcwjaGdsLJVSyQVBOu0m1UaHuwAQut1B1NXMVKy2GKklT7+K
giQBkYVtzClVTsQX6xeQ7JAUTihXS+9oXIMccBQfmwYhpkGTzis2mWC6kqdqLSmg
xHIKa5NX8I5NnAdUdD+zN9QiJPdAX/TqA37Lh5i+LJwwx/Zksa/imCWRroUNAGTW
gOPoQ8B54FcocfJpkpe1ISfUpd5GKl9J0T1tHe6Oa1oU/QA1T4+ygZJE4acFXlXl
aK+mUXAbsNdcCi6/RREZVplQRJeVfqyukjqB3J6rL87l6hOyoTgM7Tzjx5QD4fAy
HngmwuMGtE84vTWQK3+FKzTaLasK0T6Vtax3xJzV4K/ut2xSy/mGWJNX0qfvUMFx
AI1vjx75u+LhNECLb6f92/jnB1wlf0wfhbgpulqQIC6E7dvXABt4gTx7AZKAPy0F
YoX/NuMVbmM9NRnW7x+qo8wCmAB4b3XS8ZUJDkOmnkZ1YR0l6iIfQ7jaIdaXhhBa
oLLD0uZ2rwMgVBMYacN1UbnZjXQDjT4YRTLSroxUsUUt5SFlAe8hFLYT+Djrjky9
yUa5AKBpCV1TuhVOXSu4A7670+ALyUcd0tzlen7KRszpX88mcvKiOEg1Xv9YRkyI
x+8sCSn3L8rsVskTsYJJY0bAQRdJgKf/Q/eNXXy6wJtpp69tfCBRUeYHFjqj9HHj
Ykt4LyfKXahMFceY7vdTWCtJE9LSyMgla29paNy4XwYuQlVO7lKSvfPj9oRGqcvH
gx8FEOqJj/3jtBKBCpOxgJt2FoIXomnbCNYcQbYV7bdfKukaIPLDy28uBrYWmnuJ
SfNqA0Cr1NwZvcG20fKfrIx1iisvTX2GgHJDSqpgeXHunZUrxUg9yYR8vEZJffXa
suJqVkpSKhlHC3S6qUArdcfHaedebqPgKYrtrNTXE7mX5CcTFNQcWTlecILxayWI
o1H/wn521t/ovkUJJp/igaKqK7ULWiGDpVjP+Lzk27p3ahsR+GN+9yIPeuoC/VSl
IPiRsoilxzqy21YiQy5FYeppwww2+yQcHgO2Bht34/iKVm5wpIcS+mPSQ+ePQJ8O
II3AT8q93CK5/ECjH4yNmjYkJtvLMZi5+7yNzapMN3Bh7x99/EheCS+JA8pSrDXP
mpNJYKKg42x6USM4Ef1qibmFXux6gGACr/SgFM5Nw/K0IaTS2yopm2+S6x/Zj7DL
GKalnbkUumsaNA1N/6TNZwZztjSvfyPv0KMg6+7zi4vHLIMe2LK4uvV+SPiZy4uO
vjUZsLKY1cZw9Q+0y7G4tnGHayrrPVN5hohfTSrYyTWL0ajIYQwzs6ihLA2mAXGW
YyDG7X9YyaJAYsZh86Htm4SEN2LodP5NLiax4gk3n21eh6ZCcZ8cIqy82EVdX/N/
OQ7j5FbZiNYpuBmE5AMYmgCOEaJRtkpUmKS68nDLROx4iJMOh0etPpFTswzRTB/K
++DjPPSSS8VOVS0dYeqG3anVzQaxd7QVyIb2xsM8jsex+PSPMxvRc1zI+6Kd0oUH
WMGTY5it4NUBbU1wBF0dKBZBWa44GFfZZioT9MILwDW3fa/BrbL07CFcBDMKo4qC
w5tYYnXCHFUtcU2AliyWBKynGtsUPwJX5RE0jKKiAgYxS8oI29qAZcMr01iu1mIH
Bzha0LXnUjExh0GytU2rLLwIaFBi7IRTzyJGDAd6SQKs7tMqFTmKSgfLUUlRiunj
YqDDode7FHgfAjOX86XigP5Br8ji+YPnLnxKwEuyLIKUvF4bZrFtXfdLLPByIsl9
Yx206XXUG6IPEkZVig7GUwyQLghoeK4xc85IzKMFRVfEdCQoX2tF5zzRlaVVRtYU
a/K56BCT0rZI5cMbOYHfdbU1hAviq0SI1C4keLVkCGnn/5QW1qf3n1mXmgiNopuG
fbqHkCpoZhKviKxeNcOxKHsqzJM8E1p1j1ktr5DQY/iT/sum7yeOlfIuN4xMi0KF
quCPA+l8rQQvUm4/EHutYUBVzigPJE9s0QlGt2Nv8ESkqwUfrcJ8V4Vfqmlk4+mR
dxnIt4A5KgS279ooUjRPD5yO1qaFyj89Oi6eZ6yobXAHQcy4ybJoWadnxxTBYomU
h/RthaaE7uBwxB3a+FlKUo5J0nMsTWZU23AUqQGFOk/nBf2QaSTDlxLM2YxGQs6R
w2df7GUmqCvC4xeGG3Gk9LbGGCSuXiGJy1Bs6gTb7t8BiWASP6WFOR40wqKrCFjZ
wcbj6srpT0jafQtJVRNUeJyXKFNeb57LyBss2jN0tocp57wZnMfDcLf1Q34QaF70
Y25/LQgmK93WuDFc9KHAhUdyfBXwvR/6/mIRYWAux3/ZaQC87K1UfOD4J3VKxNo6
KTFdejVHLEV6ekdvVsr2Vee8alng5lO0M3muJNq2dvkb10EcCvVgGB1g/eQlxBMR
bZkwyGI1ah7OHO2NUi42v9Yk22MHAJVD8iv1ZcCpDPDHTw+ebXM1BKSuur3pFTcH
+oiKdeUa1mz/l46wMLgcPDhu/Tbb3AjVI7gvriJK7ufMDVhQB5d6xeuZxjQLG9dS
86DBpHsBYjr2ZyppjSvxbAswUaAE5Ct3oXFt8/rNjbWN3dAsKS6JD8gXdUjPBA+x
H+YL5RJB5xZWHcz6pdE1do7eDMlumoxbVPUcCOZZwJcbmnMnMpUsTQb1Wm7GFHCV
KUoeWrjjLwfiZ4UgNMUWOTxHlJjAJfzdscZ6TebIyJDvHsvuq65yTfEVQjaXNDvV
t4sh3JTKEQY3bpSy/4AkCJjlD3eIfMLLmdFPyZo08LMj2z+/Q2ROZj2HDYgB7Qmb
VtRCzgT6ZO0lxTGCkx5lCnFx7GIt6NqNFYBst9WJ/LJNq8j4PG+OIP1C6r07y7C2
ZCh95oTwNpW5wZ6LkQn+9gbdwWP5IKIkjsYD4YkyrfzpRcLl+xruPrgwGJlZlqi/
AbgDW6VwdlEBN73hn1dcWE9aMx8KapGZGwF6bUHNKNwvbBYfvLW8jFDTr7Mg1MIi
1G/iWjXUtEiAg4xQ7drlBWY0h+eC1kVqsVb7cvrHKCW/m8wjU1i/yB3oL1LC9in2
+gHFRO3s3moMCNCrZqYQYDpN/XQhqY8fnsEhr4uXfrd14rsiYxPhsxKhaUpmbTLn
J1sLqujB1AT3Ll4zZ3btOy1QD6P8rtHgDhPmKPAnorNHx9YEl4WcP8VSF3T03ZYA
glyA1SBYhfZs1nSwg8dDUm8R75lyZaZaWK0jWzuop7b83iRt/HgoY+z21dIoCr99
afuQnhSuJkEpwe5K3+LnWiU0ehqiVMuHSFY477Fq6t3uxU1fYPO0Pnp8c59gWgtb
vo/PHeMYPdj+dQUaXbcJPOZHX7/QIBgDM7y/i6u4XKmWFJDvuKk52Zi346TQ8/Bn
vZ5CGT/73d/sgQoA3PmgTbyv4hKrAsZ3gW1AN41cIQc2u+qldUb0JQ8PSlRwogA6
ITAbtpwTEbbfHf6dEo8qYLBZ/8TL7E0JGaTHFYrekD7pf9Ru1HQr84S6SY+cQM9H
EWEiKbGRNNPZG9urYlZAOSxu3reiKDMSuZX2imh2JIEt7mMwW1oVtfDU91T2FZZN
2TC26yRArhU4KSeWX6ks7kRxupmFHSLLvRuj5wqeMSdvED8QTI/8ZGDIaOFUHa8m
5CcwcKV9p3w32MiTstNi/DYXBqt3qXZryZpQyWIIrtht9G4Y8pZz6PGBMKv0/cY3
42THnJ5ipXoyrU71D9hvcmIHF+DbtH3vMjq7WSCLf+Z4bK7xH7a1vLlWHGKPFrgX
PM1qh6KoqBgDhr7yNpfxEX2f4ebbBpzeRg09ucv+qVVBMedEMQioeypWOm1rqg7Z
macU7gxCtINXNL0u0NvsSAxMvggsHQERsYmuHXu2mICU+S+iV6WiLoimuUUb+K04
tY+g3cRap5RCZaj3XGT3DG7v3nyydfbli+bszqjzysnq7AjCiz0N0NzOSVwO47+P
nMxLpLHSfBtRgOsxMn347tRNsdm6XrGTS6LY444PjbBEi38bcT1mU+ZnH4N6yRUD
N3y9RRQvmg2HgJPu2gLs9CpWjUufAQDwODW3j9ordPYVobGEYcJoPum6kkpHt/7T
Zbcu9oyka3QzCptds+5Zun192X0hlhLCBX85MRtFH2yKyf8gNmEsyRw8tuX1lp8U
Nw16n0zJHnLtW57o00J9r7SdlKfmEw7hO6sD92rVV/ZG1Hr6Qk9qzkN+n1wJJ960
4mJNJTjmmSDVOKfRzocUIMzjRXB2WlBEiIfhw4aZwdjwtiE1/Xd0++RX2FsnOwjO
4EQ3yOyzIzOV08k4n8nItOkB4YTll7+ezQHoTB3uEkOV+OABHvtm/IS4KWqS+ff+
Qn5TEsc+jdMfhChU3+sNMrEV5HWPVAqLoTRrz6RFsWj+NEQYrmtyCUA6/iezYCWM
qRJyUxNmYc/jkztKcYBcVINT5UT5kCe45yjFTKgoUcJWYgltS33bZHqGsWpQ+ucZ
oJ3fl3ZbANz3W1UlVXhz+2tiFfarUCbfKHVGDLuSz/nVGg166Y46T5VaQgJia2Zr
dcjjccVH5ZI4CSM6NkfE59JDvsn4KZfQZmrkYfSza9plF3RDkE3wqlbvfgctRN3b
ZbPhXhz03oHfkJYjL0DfNzFyECScA6zcx+Mh5lmvtj6UBDA3IQavjQEODHJf/ZqG
PLmx0SDVrRRdPIvAWUyXoYMP53NO+bMkLAO2mCGhbBqlKkXdZHDmeRgNDJYLsURR
iYCVqJ+FHm0YId/U+n0TfpoFqONWbkU3f+SsblqzJNR/xsa0XVjQHh0tnbIRQC59
woNRGi/warLopE6yFxUyRuOFL6krhoJek66Iq/xzdlLBK8wKvmnjahDjzP4oOqbj
O3P5Z0oHa6q5QZ1SagbFY8aNSRaKWp1cbawBO/DdyPkDmfH3FUjrlqUiXeyjOQ29
VHAeuaRxOfHOnzScPdWdCAahLYw2H/rSBInUmSUqXn5VNVPR5K2/n29l3U6QQDbC
XtSAy2/EEJRWKytBBsx9jCwiFpV9/pqmQiyzsOPGeswM2lnEy9GHcDMlZqKSiE6t
aJ87aP1EktxSuMCrl/IkMZuoJgOVzNwlsnL/mBF4C3CSgGL5hpuTZDzkNFL6MVgI
mmC5AytY5TvIBt6xwn9OZ2bwhG4WKZJd+QRH4O02Axy/SYYIO50sbvhDAMxUbsW9
2TUNiiUe0hwSStiqWMpjt9Sb5T8DlMdBl05o6PWnOBLd+dKo5f82saZTSf+4JMlN
PAk5k5yW39NYqlGslaEuMczmy/qMwcGGAi0OTzO2S1kake5Ejvcp/GRE6x0sWvRO
RLNwc/yjFylhih4DTGa6JmEXs/r5xJ6sPPB1R1MdXOHReTYzKJoo6YCb2hNj9/B4
2Fqz+fBXkjJPT2IwVXSiuXdpWnB1OY+/s53t9X7i3jBEzPgkISp3b6EAUyXfF9oP
TTeC8Schfg3eQjlsULboMT7tnmSukEK6VtDVVxWR8kiFKGETZRXcdlnnE1ZQ3XBF
vFM41bNChYz7gp63V60VN+62J9eU8HiYcrJ/1oAfDTfmR5CnUKkSESb0o3s5iX9U
nzbyKukFTWP6wzzUE66uiiSSFQjQPwH/594QnycDMeCFht9jOKNQIyorO3HLkK8+
CnC9UxoWnBJzZci7iEZCjC4IawhhDvzYeOFkZxpoLQVLgF4ujhadFqmwYY7Q66NS
Y6odetlUCoyE/cIzeE37Ud0RPY5+ApBhgoRX79BWkn0LwjdfGBkxNYjc9Cekz7lE
16LhVH2lQ+12FzFwdasI6RL0LmuODGG+0Yd24oMKwzWmGZZ2SzEOBPMG9k0FiJKG
Wc1VsDW3SYtl/QudPtZdi6pu8z9YCQRBVds9pzCNHdcTh8+yeUv7q+s1v7AAvX76
YPTk4/G9qTxL2B6Y2M0hYdP+ZgkBfvyujt5sS+yuEOKNZr/++j+GAsw1j7KugfQl
L9bmteDl+9fgfoIxkCGv0bmWw/G7CY3nfe39guN67wdq7zO08CVPPEknfdmd26rb
iJ8NzvHZnLlTcWwYnyBDfq0dazlu4V258p4eFVf2/Or0NPaePRgLrPX3tOlbTS57
mu9oLATwfbw354cwqE7is7wNY75At8OWtaVX8NbUIqhPsmEe1iWtf7/e6SFZBqdo
NcjRxxl4ofheq58j+Zj/6TkCOQm2zHOCXkKfI4utZmfI+usBCGhGmDY2Woe37QeC
CMt8gCXtCf3XRId8LI0c+vu8e/Ij+zU5uXr7kmi+OISiHIrxVuqqpQQY5ChdXgVJ
4wwJgMVovGFEpl6wXIqb7DGgBSQepwj0I2lOSIIyOcOFJSPA2e3oq2VJx9lnc5cZ
QnB42fK/PlCjBcDe2IYGUdBaY0uYqexmQsxnGKFUPLUt75G5dBplyfZPUtxrj8X+
exnjl0SIpYL+nFsD6XxzrdsVkuX1IPyfZON9YnBbtzfNc0CCSDtNmzJvEU6WsBg6
93H5IOfkm6WGbABm0c6p4cGG49aOBNyUja7yr9rYRnLSRA7HGFs9PxcsoVK2b8S8
yVOO1zqiUGWClgc4bXaFz9w45bdDPfJyA2pZNGPrK2NMEB33MsIUQIq6U3kDh5Qd
QZoLU5rDS6h46EkHGXW0rauqdtDrp1aDSZGhi7+dyBlNrCw+NvcisBPsht/0fRzW
5v60uqar2BtuOFWkmLzs4Y0K39TBeyO+lc3st7Ly2JeEdRH/EGiuT68/Y9NhgkJg
gXVOkQGdvxcLxyF7PLQiiknFChU3J34SX1uaey5Ys39NsqEbjDdNgYsKaWsU2UpU
4pComW04RMU9JhoDXt0vCHHD714dXg41Q/l2daJiuPTErCQhhzuibmV/lXVJ+MOl
kdcCA3ZjJpB95tE3c1kz7mzdlKFTIhXMW8rZ6JmANPH0B4jKAOLuVJhVI1C64m6B
mNycT8LLXWyHy6wkbxdqC3KK9Og5yls3xliz1ow9xcDWOUIoPUGe70yONmXb2aMb
j7J+gSyY4KVMpmpAnGiK2R7MWFz8ru0XjJba70Sd2ZxCvgzjIrw4zWksyM5NjVBM
zO1wc9yVBWVb/xcXh6uvnE6491GInSfows9iUPtPunSkwDwPjQj7oycH299H8xkQ
rPzpXDwv1jBJxfIBqftm3741Ds1BR/i9W5bCuiATON3o2Z484AwfHqcSfbvQmGHx
BQFme/ymrAlntw2trrzXSzA2Y68iisCgFc7zbv/rq3xv7YeIT10cq5W9Y0XCqfWo
84usTFhO3TJnW9RFt1lZmtKOYPpwqwUR3skE8j3SwQX55dzIT1YBig05X4NeEGcP
+ZqpqlviSQHcod658WZD15a4LvcVsqW5gj3MahshUNzANxLfvPlM1ucD4/y53bR5
1W2VLeu0d0p4htLx1r7H5uGgEhNrlZ94H7jdnBldYOrJ4qNnrOvCstj3wstVZJuj
v2n1bn/FltS1UaNzkHJHnrZxJhKToP0Yfwo8DM9+s1ID7xbAlYH4GdJMZqfyo2Uw
t2U1hN52nwTVQ31YD8rEPk/oM51SlvGHDHfivjUuXSTok2V0c6FuHV9LIpjHO+18
lFK8drsLlvHZfnW6z/evBgl0W8uR8D7Fuf8MeJiuS9ag0cky0e5vnzyzOJxDDCjB
OU/kFHXDWN8M4gK4AYsOab90cK4ILm+1SgDZAnFjyUTpffSPhJWKGR7sp7Zdwtr7
8jHfCc51OpFELiC4JOAVltdWe/09AObit/bWnXoQVY4ktPcmo0qqEDx3/iTvTSI9
KfEEhu7T93rJ5fIeAEhiClgjZL0C0G6d7l3CGWHRZHVXRRD0muQFecg7elCw/P3P
hswmNE77Y4lz/bBdhBBvDGP00J96FM+9klzqkP9MMZ10j3NPmyNm4eUefHqJFylN
jLUG0ytqgagc76A5w9itcHyQ3XznFYxWxrKuaQPPt6W+POyeD2N1XzMX/DBx2e3P
4qzJkqqaTqKvYKsOdF5dRzcEP2q2XFwHSw5jIv+5h/0N8xy40i3P6jKThvO5M4AU
FgJuKHPqQre8LfCAYS148zB62xb+M+1E4NtO9Sqb9eAxyaDq0fymYSo5IHzECYzZ
nFPzlXuzOsaWN0ahHFEBDmbI36xkzlzLnkFEmiZazvgruQ1Q19K12MEzi38R5wot
InHQdBcjP3iaOtX0sx81j7ETHwzowJChcicPrWaoY9HvXKH68zUbK9RjNtST89WN
hnk+jzMkTTtmcJYsBWXFGJ5XK9L5vci89njt3gQa6YM3T7MRSLMorgVw01ZvzQka
lJ4MvVh21BP9ohVGXhzNbV2eMAil7YN7+M13dz9xq+fapbQGy8+3k8g0rG2eFEMX
vY/wfaF6b6Rmcmnv17yCtbttWQeQavIT7GMMmdUsNHHXOJ69QB2HlesFUVxv0tn+
+58QoRq1Xu5qPyEXyStIV0J7DUNV0Z/zCm3BanMPLp2BW28qjCAi39Y41MhNC1IL
LdQphpCWn7ubzzIfELyjkGXk36i8vMu/S2psGeZFsV8kD8/M7wNlj5phw8iK6PCS
Ro0OuyavLxhXUAPpc5CBB/zm5QnwhsHnHsoKYiaF1qqUR0S4cHLzzA5ZD5q9w+H+
i9JYoO4iaF9pgMtLAQ636mcLox9D7ZkktcQvNrFa1i1GAW6MST299gbYnl6ryt6v
53YSYbBhLkk+PS8eWMIhr7OliiaOGuNUlyKQ4Y56+4tfY0N2e6Js8vw7bhDEblTL
PvYdjgoP+OQCgZswAbs4X4W8kdqNaqP9SSPjdw0JyDPb1rvUQeWW3qKdudhT6/O6
oIytlLw+mLDeBNmNjV7/o7Mr0OW4ac9/rgavOzJGcQoHerEvqL4W4WPKzxpG7n6Z
s4160pU1BSWn6W1/rA5qKWEj0zBegjO4OP4g8knIGYD+hdNZPwWQHbMBg7Qd0Zh7
mCBKstQ8+BX8vjKEfzG5DZe7oBgHbOapteD0uVEE4f7lY02VQ8YwvfbqcrSGumQV
wIulNwuNeXmYV2v6G8MwpxYI+ev+ZnDk/oW72VIVSZ8tz2ZtaSdNQXmH5E+WD7wq
C5JsTcL2AGceSJBp2dG/A3u57eIff4r7ccHE9Qy9DttgGEfmIHDJzcJNwbmSp67e
k7JAkOkgwuEygJnE1R9yKpkLQrRIOg1qU2vxSOOKqa7RuU58JBNFYGeA/hu3GYS4
1Bbw24dkRrHgVoykC7dDKbP23o+PkFe6wSEpSYQ2sTMvm5CwZucenBH9/iSOvFih
61AJZtynFa3ara6IauJ55tU2wxkGHlnMo5nE7T+BeKoGMorfVl8QW2YJdRaNwEqb
rGLp2liW1rDCX8NcNO3zQAYL5cn6F0aSOqep1aK+kKuIpjDUrgQD0xknW31AYItR
0zDPeVDnAA75YBHXlmn633CF6BlOqViqpmsuY+iqYxG20WatnR4f+URQLtFSK4Ev
fFPYqQ6zES+4kIzlVtl91+GW5HEfyLM67WB4q6v/eWm1fp4jnvyB/EvavS4vOXee
RqJ9+fmQIaET+pHM2QKpSk0BXGVaqWu7BVZQLBCMriU/m3s6wWq5bAeLSqdbYZ3+
gKOTuis6v0G2dtab95XSR40Ji4lIGme7nEY0oNpEtsdHHN3TE7MvIDOUqiTrNjHt
l6rQSsAwKJ9Vqgemftnlv7pAqXdfsveSvNoAzPbPC9fVjh3H5kFqOfkGvU6qAefg
W4fBAf96FBDVm21B4ufxnsAhdQXOrW5tac40coOZ0XWTTo7pES4TFQECc3u/PEVZ
9uOUSsRDcGNdq+8IseZMqpZ8/sqt0SIn3hjuuFpC8iOpZpb7NMKQ6dYZuORkp2le
JEHYIG/yD0eU1Q7EsrkzeICtpJ6Hw+lQ20byByID3x52Xf4A6o8cGEXR18qFNAsd
FLuiVruiRWC0XyK0ak49a9ybBkSCtmujmQ+QZWOrFuuoSXOpcPfyDpkBrHph9i+b
eUccejs+JChj/iIrTew2jDykDIBGehgCen9SEEQEdH9SKoSAsP/SGhSBVRL2Oadz
og8Y80Lm4N3mJ+YteIMhL1HQuRxINRd53AGesgwK04N7owdqrYTYeo0pksV8xgyo
2fVo01n42/nOAxQrAYN19lyTbxtmJr+Hr6acUAjL2pwUioyqcL9k9QeTpcZl3mIX
oBfc6IpBys9yKxi53DRas64RX5sXrxfiqREO2oQKgYnUbzXL+P/ZfmUNWFhVoclG
nIsAUgpbuaOZZVGpCFqVwng8w78H+Ks/l2lRPZ6cBVE9/HDR/U8Bl5JTs4JTXEQb
Xp0JroCUJ10ptiCuodoyR1LLMQS2bT5N+oVLeLEdIX5HDpXvAKY/vi+rzE9Ow4ZR
xxfEMXGJylffDSKYlKF/hMao+TUvWRoMmcljUphixzWCTUozl+SG82cV1RjBb9H+
v/aoPuTg5EoQuvFibC2hO0/cUWx8/tOdnq0jy446kzi22vdX58vqXQwHLTFvS0Vt
Er0859Mk7SW9QQLR/WQoydiOy+L3IOwETafXykbO4IowKrM2mLPPnBsnwa482S6/
A/AQnLBoSs5hOGfrR+XkKEB9+3GLPv2XwNtqitrnuHtxUIlryLiSefpYkOMicU7i
WlzUgk0mVexlCXd5hfpDF9eXXCo8oBSZBpftQFRyQM7Yx+HZWR2DQ8mo05QHAq5i
kVBzzUSPpQjbXsUrUaRTy+Uw9QbBj0AFHlrvpxXLNtChSbpjdJNQSL31w5sukt76
rVPebsqGWOkG7DtgsSSZZDgFa1ooVgx6QLA6WJu4HlELIsg737IWufCHj+v9dFKT
PIgTE1oN0BiYy9Z9ukE5smpcxNJvxdSv46sWgeyu5Pk/DpXxGXV74UnO8PpsclqU
YCpLnJKErHXmK+a7yWqK2aErLuHl+wRyOeLZNZUdh21TWjzohsQKbJkA6BO0XL3G
G689WM4VU57560d1CpD5xaIqp5ZCEVgCmGVpEaMJMdyag362I7yehu6lKdeQCF6C
Z4sMlhXp0XnO73ZyQ9ILUvVWUXmsjfSePVgcQXU+Sw+NjM033vRtS+Pf/54QBlYd
Nk8OxCMhA3NNR2noPGy3pfI/flaY1LOkqe29JMvg8IOwi6Lta0iwzE9Flb3UrwOg
6GJAQQmf6Z9pb6/ZuTHAX6mU4qcAMhQ4BsWfQAySYlhjD+GgToehY9BwAKsFastK
ZQszGoEtSmH/IEWJNv0oEi8PnnKI9jxmswetNZSZBhBYurkxdusCn7tvb2UHLySY
RUa2Y7Lg4MoHxCqe5SDcUxNmLkeneOoA0CELqEhq3/eJjKd65nXkKulmalXVJywl
oHh1A2xOXd4hfo4x2/pmqJDt1cadooU5IaDerF4OfdWF1IK54Dfd/SGGSXzW8i+I
ZOFa3Q/LmsmkP0lZa7WOFJFoKec5tD9kq/uexQluRA+ENghT+RZXTTFKSD+2KvT9
hxQuZCMzxRFAlo8kCC8mq2D9nXEKhXLatVMSowdUnvQozLe2BFZqE/KhLoiH+EsR
et3YelJMM48rrAzBlIvUBYhCaWLaDmrkCrSVjmLp6o84h60mjFcNFSjgj8OHaiqD
CYJPmhCUo3qfO2nspjnYacY+hEpjrVG7iKTkeZ4eyHM6fh/bZBvzQD3I4LH5o1JJ
LZvrP2+Pfia2fbcY4OQXDV3FCP7+BeBJv9oE+JlK6AFfCZ/Sgf5TegBSDspHpGLI
3+9tGTcYHcG7azhEFcKjVdzES8UiuSjyWlpQdBcnXqxNUZgRuSF3HYcrdY3kd4sa
xlCe90j/fiPHQfqNvmYpR7dOJ9s7ROq74Yv45VbzBOQNJhR0997cTrTAMUsR+RKE
/dKOfmtkrzl4Hc+YiKc2RynajTCk2r/ldJkT1XUhpszoiqsLzXIWYFWTTddUCmsE
cAsI5dur7eTQRNWbcdXqtE4k777mDf7XxNCrbPsbkSu63UIKkAYPBw45UtOamRUd
KMlyIuSB0w77r6Ce6G9gilaYl4YZECsv72uYkF8PmiuWPEyIg3JD8e3Hin2r/CaX
DIA0Uj3sotv62S/9Un0vGGDZPcgXZFyu3J90Dabmrrp4bdbkIxvAiNGfmPuDTLUj
utEP1plNh3/ezUTZC9UtsQ2454sk1y1xw9OanSNDyZiFlrBzxHQ5uWI2HnbAJjgy
kMv71kDzGhZ2rKe0tC4d62Dw+kCdiTqdvwSl7o4eUGwrCCVdti7FYl2AyZCwYLZi
HPb7kiL8VgIjwdDh524IYr9zRnq/5m8s5mxilhnxD5PT7UdcxcLPI+6i8xv2aRR+
7PbqM5UY6K0uOICShYVWOcOjdAPSnlF37nk/eyTItwXe/WDmuUeNyJyLBFf2R4E6
2DtiNlMiX3yxzJhx8imAfhVuURmIGgKlNWyAHK+Bit8iScgIjTwDxvN31D7MxVTS
35OCFZH6+RkfagBBd7iDLzna05z0YWw1XgIGQ7t6xc/w3QRZ2poAuCoUzkcmkLrA
n/V2TBMT2ajnlkJP0EHE6copuavC8q1g0K5QIc7JUbwjRRCq2ttk6t5Sjill/9yl
5tz5QMYIgf9z/xgKWuF8LODIR4YWcRlN7jGHondARSTwH4bWCeV5Ij43sLnuSRlQ
508ZpYegdMzSC3wM4LBPMMQzVpxEXi+VY47Pvkd1A9JNDl0f542R0zvX6umDZPve
M4GywPO7AUa7XUHZptrmevNtEDpcivZHjZ6wW9tYk0jTCkjIWN8/IrPyO8Bete6E
fIkbljyrxFMO/BhfdwCgy5o2abxxBO318eGwvW6sSRq8nVhnK/5MRGk3Iu1t4xfe
WPZIVdOevpetRLHY8+stzq8g9ZJvnmM0z7TCax2pg52jRdTurkDaPoBSMIjJ165k
8al6ySoaFKwrCcU0KPxtdc42r2YA92881WyoDu0c66Ea9q7tgLoqVKoYPGnA2Kn6
cQOsiE7juyk2QzFjdsIjGzwAA3ZtLHLTUad/uyW2Ybiofqs8f/qxPbcs0pIQxuER
mDgddmrMx1Ch5Q0eq0uAg8/8heuhmWEmljrvwn2qVXcLx86gBFxsdoTneZBANFwE
52stM6Lr9j56uwC18Oci2TaD8Be8RHGiJcanG98hz6XeoUIXYqkyGF8wQuynVlRU
rNL2jw6TDihAARStZaq7F9+GeOAKmaA9XhB9rqJ7O12YebIudPYCqydOwKlKqMoX
rtgdvsyvWaboL1JkRseM1VDiAWlttekgD7hRVSS9jC4V6H7LnR8rK2Oe3ms7XceU
mg3Zek5deRXHbonLXJsTP7jkI9pum3bLPtuaN/ZMkeTxxEk+SO7G1Eg29/2MDqtK
J44dPqbHKogWnm/VOlJ0nYCEkX40fOW7vKfz2UJjh4spcXtDsZWufKuX5s7AiC+P
RAfizHyV6RPAVdDQtC19SVW1WBNif+e9ok6mwUIxjylNLR2X+RLoHb7CdsP5t955
pS8uzue2NPKd2weuGa4bhgVnJnKtY6wUAs5nTJ8ZNmdz3270DQY6IiLlFEfxOJA/
TFKo5pgrN5mlTQfA7OOUWuditfNOR/xuYzSsKM8NxwVS3ZbajdNRNAiCA+Lqmp4p
MemFu3UeQtNif2OfoA/Ie1zurdcqyZnrq1dU0Yy6UParJM/HMsLF5Th4U6v6AlMd
RoORwwSKwD/dR2f9IhQrZcoMRRfN6EfdKUejmBYGMkxYw73WlL1B1vvfZanDpkHT
ZHTpFrgWi09sWOUzrGGaJCRkEPIMEkYi4eIU3fW/M/4Z8o1vVRo5NWrtVNSR+8ac
WL5FlpvThdqXPv0qFbQmZWpecCufrPBorGSXh34Zj/hCFE5VG8rtytHvL3XWTPmi
qtIrZYAvKPBjYn2L+kYqXAs/Of7iFx39h9NVWmQtzX9UoPm7Jpwh6dm6EeSO6Nqd
sNPjOtV//X/k5kovpFnlaoPHbyrhykJKBvJ4WpZzAtL12ohAi2VucA+YYbT9g5/1
T/h0N4f5F7CXxNF5vVqbRwt9gUdNu9pxW2svtXLh403G9hPg2zT4/MRd2I/4tXsY
I7Eqv1I7qUQRjCuiWUb7DswCOWBocoHG+8b8WgLjOjyuzFGP6TkT8Ye1AXHUrLqJ
7ac8pQ/6Itm1y4grjJWZYWljNHMwVvnCHMTZg3H9qkyq6RYbBeiizNrTsKMbBRlR
vktVgVJAIgaKrB+SrTY++U7cNEDn/hi3vFNHjXSKk8fH22VKF5u0P42FgBR/5Eb3
K8VWWvmzU9VoBSctDm0smZkRx5OGYmrbmcXvuWZNXbr/9aR5gdgJEbgS12y4zIEc
bTZRDb+R5kcmzICoKYyeDai+R618AgK9/cP5fl6d+ig42wMWsOPpAOPDqfyt+q48
nWiMU3iXjKYHltoKHo4Vn8EnhVkWuK7UAT6pNn2L/ZXtuAssmbsbgyAJyJCO2uaj
RQKcdHCd3CvkfBAFEtd4LPbZe+Sf//lQaPoMO8O40EhMsIH/TwJwv7H0yfdkdo0M
yxY1NhADs/VkkKdv6pILHIfHdCIKn91wyaSf7BK7nbyQEjbZfTuojuVNghwatyNj
BClVn6FHhCXqfqzE+BRiradi8kA8q6Xdu+h/exxI2U/zcYOBy0bYc8YTg47+kdmw
d3MQ/31fjwZv+YgjHp6+tp4OknD1gJbRIec2XF2BVvOm4eLgWyXE035ItNmxgATi
rVCEEoIT/SyEz2dH91yoyZZ6QJa+M8s/EFDHcz0Oz//UbdVAqbaYPYWQR122jfQ0
LUdxCOFVzWhpAc5HM3gbmQcp2ghP4BOm8h2e53UWJ70VpfvYrQamFy/sMJcGg2X/
j422tOd4qivUl4fRZNpZNwp/NXyqNlOf5uUcoOQ4Ack6uGZfhQcLesT2PZcEuxzr
JY8chAmw+ffPazcjYPvcuzuOjevlRsKDpdh3slTpQqTqRjfYjZRGmrsKKgRbYPPL
isVoaH2kJN7kg7Vw6HXz9re5AHP41Ji2z5PnCTVzRaESxJcuREYeU6dfwXHQoeZP
G38cNkzHxCZwdas7WATHBIKCBXoHbHT7WrAwqxXlLLPpNV+mr2+2M3jy4bfLBb3P
UNFjrsH/7XuP9B6J5bQgPNc7WxZf18w7K7/jhX0cL/x3tZUpQnGzMv3pzG2G4uJT
Z4UlEayrc5U1VmTIlWPxrPhiVFOWvzMACddeMKP5FpQxI0rwt4+s9YwIdJesq+GJ
U0ewcllntHPtVSXMl3ozgREMjbC4TfYm6aLatwxu1ZjH3jYIV5i9W4gNKH/wQUgr
1aWHbS6bFutZGwSkVay+3A6cvG6IAlNuYdDw7jMGcxIxZthcajr+fBGXHy3S51z0
MnuXOM2Zayu5C1if0hw0evadbobbmyVqpQ8WUSj4IZAqyV3WVhcklLM/bGqBdtqc
psjlLJhzL2ZGfVWDFZAUxYcY+TGmwQXMoy71o5vSWLBB2j0cX9YbCGaH5FXoq4LY
8p/d9q27hvmWMTmMb3Pqrhkge6xIOaUi3GKD4IkVtbuh/pWqg3jYKZvVks3gbkKE
D5I1kp8WgVL7HVYLdE3Zhaex90KjFO5z764aKW0zX0DwFAPegC960krwsu9AwI+F
AePyDMc/tPyKx8k6+4YOE5/MP0VrbKEkJi4Ud1JgW7psR04DB5GkjPoInvW6m+wo
ETL111ARg+aE2QtwY5CWU9PbKP6NrMNIyV7Cg4L8PwYvZXmujuMfGyZecFTYDDKa
DdicRSs7uWuKu23OQxRbaP4qiIPnkSEjGpT05QGZs+IgFx+TVvtF2AaUvfXcQBsm
QM1Ulu2FRLprikw4nM9ow2V443uedGZJggmYUVKnKwziGu6DlV+/XHsSyPx6TH/0
QaegNDGjwgBNBWF03yI0r2O17TAHLXFKJTNNZHzIsC5vY04gG4wSPdPa7j9Qjm5c
3EPG8h8Pt2JQkfYQwllURS6Cjk27Aut+IF2XSf2QSl56wqCwJ9THB247018ADwDf
HVTNVMWvsu1ZRLqctPz1ZmHz0hzrdPya3NdzSQO2+02QjFAjN8bB4Nuw1rhYv4U9
pfHxg/aYm4R0zX/v5uHRJ/y7k9xBTgHCW4/9h+UrwOr1fsyBlgAuGAk1KJXGZYsR
buyfksAZ+CosDz9v/dGoPyJXIrsNsmBXRCbTwp4OGdicYlyNCxGjvYjgdYAvBQnR
Z9OjX5R6A1J6Ako6tHixIS0Xc5nX5lH3h5+xsBtPzDhHaCbzh2SEDPOja9Bd9flC
s2eY81QYmR1+wpp4gYzhHSkxs+XStnrLUq8zkMENf/ITAcsolxfVKNvQzMVgYDiR
5zmV4qBbn2jrDDu9qzVj134eR92vvcV1MmUJ/1Zf4+TOx4KAdd2TYmow4kEwS0fZ
v5NFrSA0qhOwgCMlGrS/cc7Vb3wJ2zqYAkDvo3api0G4+MMlBUbAJ7IFJV9ufj4b
5a0ipqqalomE+z5COvpR9lui9LggLUoI6xdMb0v7UWbT5x9aNTSZb10C+5qM6knM
2oxJjgk53TUFwrvXSFCS2kX/LE/f1hrVAKsZOOze7FhaE7XLI6zqEEDOBO5AuXoq
tZmou/u1SCEXIR2jue3sGgR9lR8EzOKHqupXNZTC978exrppTz/RKE9d0SU3iSgx
tYjkAoW2BtuZkAhvXXVFdpDWbd2QGubA8OG3pugwV3acEg8rTGi86JIA0wAea07e
0jxijPbquWz4tdTxSm5Unv1hco83JdZccgBWEYrWtWP74wFTwvclXbaJkAj6fjzL
9Z/j5+L6uT3JAT/P9P6lGQddkjvtMaqLqlgo76JlPUt7FrpgcWcFCmUlN7yA2THj
F97L7hhDUfOAaOu3fwpvU9zSa7qHEWZR2AuL1plXDrpqCgfDGlcBnmQ0iSGKOrWI
ejCzJs+rGVvmxckr8uQrE+YLP7/HFYSy1nm7AkmQ4fDUkhkforrVdF6yHp898uwG
ZjMfQZqSdz/tN7c+1aO1jZXa3MQe3LlpKvXvU1VOXztHSLBbUR4Hjei/rZj4AKP4
5zlfhEpDqyDmfBVe2ASp7sC3eCOjrKa6ExRN+Whnbnq1jOhySECm5lL9Q5Rvmrp4
Pj4ivNCpzEvTLyD9yibzP3Fz7U+ZOgYPDxIMrz/j6CGFgKzH75JZhQ6A6Ef5UXuN
hcaWvfh5B7+QHGfldBOnenZsztgVaT8kQzg/92jorze9GrVF590I7AeQTKkHOnrL
47kr0JUuMxahlTQ+XRAb41CW8ytGgBeeJeT6PgjzUQbjYgiq/4dswGfUPYvwST9I
Oo3OdTDv3norsS2tHCS2t78Tgo+xwkYqJngo8WHAtM1IIq7vx0MMx13f/ACr73/O
6CFOS1wE0sTUWY0ReDb2bAtAM+giMm3MjP0Hj5XihCPCZ++PPKt6/bNAQn8BoJ5I
+w/D3fGl0QY9pvre3a5eDwjWZi+Vd/WP9ILW6kUxNmatbsxrbi2CaLUaPOdkN6uI
UFwFaQVjo68Dc2uLL5+LAou2jd9KIrkoR2S3oPvgV7kxbWHApDVFMnXyQZC1/Q7m
TWU4FYc5k6z8PLq1ICAodEJ06IRohMzhykuqdosU0EdXfsGLSOLs+FO0AkncZJrO
AhECKpftwsfDGRep7ysQHlM84LfsivRVrFj/7h3pKmHB/IrGit21GhYNcsDZP0k/
24KVx1WJxpSiWsgG+xXaEsEV7F72NUsOpvRWuG9NY+quWqnXpl0w+Wg3pT5dzDug
Y8vlt54ILIXXeDRTPp+5qqXGt2twY1OO+2Uhc/uBdUJd7jTgjFXFM5qeCD4Vq2ui
9GKThnQJUIbol79ElVslHXicQWXkJg76C0mryA55k0d+SyRTp1noGHob8+rteNH6
NjTHuK2Yzfz1VR2BYQSaGq7m/WcoQHEwo9D7rngzBKyGAd1kmOi5raeIj34as2hi
3ODX8mvJzEEkkxypv+vlHGx0wnpch91pDAPU1RJOtTwFSkbXuqPzO7ultnPvghVy
fEdfD2zFZfooe5dBCIF5DIRQV5o4Cy11w1r6NeCiRQoV0GqS7S0gW9iIdWYpB6te
84IcMHdM1l3dC4IWWtNo3jP+3Sl5BYa2u3N2bvgbdtnOEx0J11DGL15XLWjPuoYs
iH1hlJZV+KpZebc/jCWxrNROT6q1OVME/8AFs5Wfi53jHl4EeQZqPIf/a09+f04/
TbbkSd5ZasUs65t9SdxRVWDaR1moqCl8wXwmwIhcCwfR0aoXZa5qlA+KZW0L4jEQ
GlnOACtMhT4iFFepddFJ8TKn77dLChdwwYr6V5uS1BOgCJD7v+Pb2xkHfDPlMrKY
mNxUjXDU8wnMf8htbnSUfncUaR53f02ZntEBxXkoLhGLl6vUSbvFqCneHwRI4Ruh
hFg/esdjJfqdcZ+JZFGmNq15GXjblacrWJsvYMpFe2Iyzz9p5lX8jewS8h12Sw0/
i07acOdfQZngJ7acKAqp0RUcgI9ydiDzanRI81qqtmrvLxzchO3miT0uw6r5VKD4
p3BywWp2h7JuqmQZrPmAk2/RL2vGv/+AyJuXo4f9vaqFpXvW925o+wDLGm1dTG7v
il/f5oXgrSHiJWsjttcyp+50C+fV+Wmftf3SN5jLS0+/rYrOLHno40X5A3RcaB9h
X4strdL/aB8ds8cTJ+LeKX/hiS+4J58C/WtrMRVhRw+8c8sbBFkcB2ll7T2pmXZu
g6JBPA3oYfgY0C+ChAfyqKjV0zM710zFHuY0Ai7V805F/uiMVQIGWov5a7PJJHDK
tvawBhdNlj3gyY7ouN12JYba4maHjddqjS/t59PbfkUfJhhT4UO15VeinSKcWPnj
Fe1g+T2no/z8PpdZBISXmroK9zPseGFSN8kvh5mIyETbTA+1+HyOTdM3bw+tLp3y
ejI9NrQZESrOfQ7lIIQloIK2539G5r/cBGVFK1Oza89Ly4JsMivmp4JW8pEXNJMK
QiLS9L4AFNJJKt9Nc92dazUiphZQMJ0giJkt8MwCPvyuEGL0LFVGpOhEOtaBqiX5
hR2A9l2jXSkeFqUx3Wq+3Asc3KcnCryhw2QREKPzeGNf+ymb5Kvx9JymVfYBI2Ha
fO7kqastdKH8cP1gxhx6n6m7977lppZVS9xzXnJerKlfweFz9wqf0TvOVy+LVWSR
J/zgsod6gWdNRImMB59PJ1YsMmQte8KA2bQyOKa36mFFvmbA4jECcJiQynUGX0Iy
47nr5PHJUY83foktC6YeLBnQPwOERsuVJWXnhus3J/839DtGfS2oaAjVE+vR92Bd
gzs8HGVBHK2qX9ambd26Hv7KYURLhHDjKrYZRSY0paBmbQ/3DBTmLznC29bPz2gZ
XvHm/xppl2ZFrv97ZTkuBQyzE73P771fuJCR0Fyv/BqV6w7W+MpSePlJT3eVNKna
57YPOPyh250f8Ng1eBI7nl2yaWHfNt9bOFGbH6bJ6Feg4OcEB9NXmDSBE9QYpCQV
Ns1Zoe8dEE8ewXCPKABM2LuRKXC4Ncxq9gGCcpWXEx2ZlNt3BSL6/FQ/6V4ZIhrp
v1fY005+eVA9e7228V8tDR6qIUZKoIm1vvwtYGzDbjbWPKn0kTEnD2We2gGZpbJ2
DnNgZY5LSbVmZW7JeBfA7QmaoQtu7kOIeOpiF3mm4shj+K5y/ru2D7NzvT1v9ahR
HqmSU2n2GJY3IBT/kQU6XXAUOggfAaQMGvjLHrSzXmBlJo1Rj8kgBcKvqsHYOd53
slvB1of1Bj2R3n0YcLa3t8rOFwFlN4jAhBzNSbNdBK+lZO2ujFwnNDv+lFdbRSQW
AaHv0N8gHqxNzWEx0Fq9yrgaKNJ80BUmNHViCDr24OHCbfiv8a0brkKPrG0WCsSZ
9VlXMC90puVmv6PK2vkxebntevrRGX7DucOFf6UJKEs9f9SAT0Wef5hGxYWKY38C
uhOZktaEI9XjoWhYCjvo9SKGf4GAPKp5coGWw4R2DBfMAnDqoQSRf6rvEkP+gt0k
0hirxdn6cycKYjfn7Cc2qEsZpwPaAEFjpmz3qCfVToBNifuMgQB0dTs810XMtlf8
3cbAl7ieMZoPvT6POw3ZX+VWttLUIlvAJj/3/LYT/4RreV4VRLGS6AJEqvlHd5KJ
Lfzr0Z5F41b+2ern82eOrqClHHir+aypcUJ4BPmxQXfb0jSMO4i0RphhpiTheuos
KqR8BdgQL1JpX0NLMFBQkV0PqyQEqXa6wdtNhSC7jWBgu6YVmYqxrjHaKbaWKxff
1xh/xWR/X7MkS9NDHfMjQGjVRZbr5YXeJ57RN/F1CV1hVzBxuoQObw3IYB/PyJ8U
Zim6aD5xTrMttPOd2mTrmFx00HOU11LOwdYFeV4NaAT2JFk2WCUhKRKchTu1p1MJ
I7UDNx4xSi+GSomS7zsECUmJeylIVKNq5RwUQKH02OF/cKlSZyz/Wfr0Oen7vLHR
6aiqv+bZoIgsstvFwRqY6rhKD8srVISnlD/t/TyS8Mle6wAVXgHapY4JrbaQmpEd
S0fneUhv6nXkfspz3BAcjXdohm1EgvSl2sR0b1SgtkBAGOHxhvEUOwpiNrUthNSt
5KKr2+giJmjDCT0rVvNy1NZwbwg85qLatCrxCTKA0JN1w5eQ3a4mekSTQDbnAcOf
bj5xvsJ5gP4YJGeNRRrvcmfs/xBZtONQXdLosrgon10/2+7UJBAVCOu3iLrTMfD2
9qbWBmUjRWjNaw2q4pwEHKRj37TOFTEHRzR/QRF6xMf0wZ1wxM12LrQah17pGg1X
iVb1Tt+c0k5MCqzNTCOiuP5Pfnt3AFTERL/OSUhZ/bqBDWVqEi+F6aRGq7aIxgnF
i5ZEhg/TxJPr+gpgOb2dNIejFp80tkjRBkeyqnmFIx/qPifKaiKORIgqiUhGx80k
CuNpqPmDta60lStn+O8mD1O3uU6Dndh+3giUXDL/HCZdpmFycMQn8uP9jF5Zkdwt
6IMrEzx22AqlfFNRu960dMiN4LyxHsKb36nzyRoYwQ4Zqn/bGoXx9+4RJWy9jJRn
CAeJfe8Hp6uJaZ+COctkUms2SHVzQEi+XUC8a3XM3O94qbuEiap01ZPzr4lUrkXu
LwTh9GuWHJOJn/ZqR3YM63gfDK28HgNwjCM2rEJaeIjqGbvf3NPgsz2OfDPkWHgE
1pXg9W6UDgZQeM9fmcaI9wpQengtsgaTawYVPSQf//j9EeQY1OGKQRrJVgVE21eO
9CFDwCG8yPgJAvYUjuZMVtBVVfv9Y6LOQAwnsqcuLla0ytHz4sn5IzFvB0r5DVHW
nT3RJtFO8StYVIttHgIsFbCmLOIA2Yd9sDGGQvPCGYc6J9QVbC3eW8wVO3rOZ5Sy
iccjEQfLimzaGaDakHT0ZUNNl8Jl56YIDwHBZPG75vpoUOByUemovdM19rsghJxp
aJ5fnfsQ1MvXU+u9sjt1wPifkjy2hIxR0kmiYix51KlffOCMj+uMehwdMvl2cI12
WXkYGp6PjSxC2ddzotEExhu7BmZxspc9oYfvQAMOAr7BvRilJMHYXuVliD1pS3Vc
DsFcG3wQc715PwauNGsAhRhv3es6jgBFAhFkeJkyrQMhtKQ2DbO1V+PjaGhAIhGD
JoUD4FOxC2gAixiLxQUoBk0PDMBcZ+DIzuSzLgVoQ+ruy2bagAzoMqEymoZbRQ39
RAtVKuMxzTv0eNJ/GbKLvP5wQWs/LoALDBcyIDrjETNFILx3D8/WMadL5Nwb6cXE
EDQo7InACWZbY7GtJBGnMx4CBrLApSaZ6tWIIZSGEe8FSS8VdAfeHXmu2Gm+sYRi
Ul2x+kj5soWnGW73+dl0G5F4rrtxexRor9Lsf8OAEvvqTCdmj3CXUzNPkrpreH8s
6mEkAC6yLpkuKGKi5mq/oRGCfkB+4nVxx0aKVDJSpno0MT+UkLzJ0l6wv9tp51yP
HFVcQrM3weMKrY3QPSkwhzejJJ4GK0js9jRXAHhkSCb+FxHSpidTxcx8PCT+Jef0
tO4KbHD3oW5zFnyYLBlfeR6KMyQ9i1MT8Bdj7mtDh+6ji5yE0OQ+nB/iohzLAFJL
rChnGyUD0hkEe3yL1IkypW/QFBe1MEccd0A91bwB9OhwH8buq4f26pWrlDz1Xi5S
T9StVR4fRL7R4EVzW/XcDycEt8RBZyb4sJB85Q+XLjyumRGX2Qj8fyR01/ed29Z/
lmvyEUpXRwnqqmmJee2cMULlELSlmeqcI7x5QBWAHrOiQkX4/doqo9ILZxvn5HmG
LASkXbNPJVixAxBs9mCq6jWZRn6kPeFVjN1EZbxGt9uj/Xpv9Z0QmGIPwwU9Pgt1
KIT9t60XZpD8F5ckX9pLJgVKgL5fxYdBkbF468fgpnBV7NeA0r8piZPyjDw1Nhfz
6vCGA3PIlLjDmBBz4jgeaMMFucHTn+BmZWq2+efIty4m7cC9EOrU5GfrIByEvcGv
2zmKoWP+U4KO82UTh1ML/9auBbLJCO4IbRMe223LH/OJFhCDrxTlNYoJfP/Uw/cC
oHVDM/k9XY77rVz9Zspf1KiYbOv1I9eqNp5VJSo98oXCiho5jYQ3FHh06ALaVwKs
1KbeT4QhZIKorzOsxSK5k5l6tbma/Bc24rnxpVdjDkquu6frzkFinyzqF5agkvhz
GAaVIDH48QCJZ82y6b7ZJlfH7vOpmbtCCG0zN1T5dUtt3YX1oFVoemDh1aYbzLgy
AA++mYwHfJUL3prgTMxcCnNjVWm1Q+d1XpN6OekbsPg05UCQ+a5zzzxAAIIaq4jx
EhGWAxNjcEQEJHtGGkj6FDqK+/ZeVJuroLv+lUyv/Yu4kz46g+HDlU51ivR30Z1T
d6CaF98kzr5ynSv2AqsvHFS8A4NBEVr0LOUwVmPFDtN7JfiFuOfa83rXh1PXgFDY
DFWz8bdpTmNwKcTeHmZ2qwTI4JdgHf7iSVgIpbS5fGEmoetnZ9MK8SdVVpyjzf79
Ha3ex1uLwKP31vbPpsskX+Ncvh6XyEG4OhWi6fIZOJK0nPpJB7mTm08zpxc4VCtf
12tCImiY4Glk+MqveTs6lYMrIT0P9VXCtZ7I9lEpNychta4hKmPIhCef7PIsNI0B
yCG2DgKSyhDCXdDhGHmZ3MDL24CGjyp5RSUzoTaJxsCTOSCwasRqpZlbLT+57KsS
zHRa81TMRjiB3kpGbyQkAi8S9r0fJmbLxplx5dUZlFmyz706b5ZrxNoS50COio61
msThotdhmlRpTF1Qcn9srNvH0tFtaDOlJslGLjKSOcY2vw7wgNYEta8nXsJAYGIc
0IUWyRVWgyFNDwZNcrZ4w2rgWYEurjSevCoxJqR3LZu/7HwbhS65ClOltmrg0Lli
KpSD+xdOVY/eueKW5UExe/5VnkGXZRyPD2paDlLFwkVzIjblUHoYhyVeEkus1GTk
5H1wDuCYnqr+Uebk9+gBRVD77AdNQpqmL+7chD5HuAn7Gkqyv9+bn0mm+3ZuvA6e
RMNgaaYBdAdK7mTtfYpsEAh7rd4ynOJvAT7fL0NEmPmIiQFwBiUXoJD/1zmfJreo
gAOXG6l5XcAzgcE3RT/B0aKYJaXD1dhgceh+etAYXWjcVrJTBuhNNnqFXuh5WEaP
f4IYSSAqtMmimosK4SDxq5kfEydRSEWcOsq+TZViZhOHeMcBLdXVTLtNP8HWKkT4
Wx9xO2Z4EXFYnhZBeYb/vFF0eV/lAopwlAENflZbwOCmtqNZ7gZ1c++KqTxaKgZ3
No/20HvMB0RdNmah62eVUUE2k2P1vGBXAsWH66I5JM80ipurd3h77m6Yuyipq5Zy
DeNnjy/Fbxlcd7BdtVrpyHvujElVY2joV8NcAaSahwd5+pKYJk+uEovCAOidLL27
6qacXwyYC1miizB/PoQL8hQiflcfD3hvDWlWcrJm8B6u64lF2Eg9P0bMx5o5kJaW
BXGf57P4W/Y6cgIPMyJkr0oEdflfNMZ1QOv0bUzbyeSxrKYhrX8bm4tYcewNMLbE
q5laEftS6mBHvJd18WfvX+VYtUGT0GTLdL+59Clz1Zw1mrL7l1r10zf9wiqwiFum
pMeOQ3GZio9YuyWFbOwChb95n6DDtY3U9p615JQ5uRm8RYODAfVPsfzSGCbmNLSM
kV9CKBQHHx/xMPNIz2vBcAl5NgosbrZGw3ynOEgq0JphyDDxubyBEmVYXYCWvgaw
Bp3VGxikDkfbznfOXx1wegnL0LwXzzf9Ym3Mb6v4anrKsNNp68Fy3DtJriLfn44r
Aw26Vpbdy+KC4DGMufJJmd8gPelBPIH0qBfWumE6/NExD3CMaEiOGfj7Ubces+Zs
j6NyNIPYRCbKjRQmbtr9ozO3mJrehZUQEL7iJuAsKdlg1L/A6y4j8MV56Mdty9wP
FKwCrp/My5SaiqaI/VHZr+s/QpGYn+Hf919j7nMLW3CQU8ZTlxa3jcs6hlxFbu/5
qCr6dATw2lDUxfi2eXUbREZWvxO97kHysi4/w6WD8yDmtqCrUtOfd7AguEeYzqjq
WeaBl5zjaUqhWTLephKAGupq89rFDY6/0uXAfKaFz3NlZZLxYEF80uE2Am/ov6HV
fvKq9OKRWoxjdirGG1O0yO8FdlAq1gxXMj87kiE0AIeEjsSr8BbZ2/tK/2EBGaEZ
HgDaQYKC8+7ArdkJrlWbBEYm65jWFsazJ8vOmlywHsnWd9kgfXzwFF/V5oB8FBwn
hOuOKwwy/1jx5zpCiTqG4mQxj6J3JgBjfFJX9m3Z1Z1yHvhQrpotPSoRlyefG8Ep
7n83EqLIXrxyOX3lyIdEwWP3RsmccQYyKA6fFcRkBnr/r8iPd94EXFvg/LTksz85
ZOawYPltdtAdjY+C191dRdS1TI3g2JHWVcvA1WfTC0mfKqKx2jO0g3x8dtt5PwiV
Fpt20Wz5Tf3dZQlWB2V95Dbun7HtBe2zTEMXPhf1zvj+sNN4p8empXwM2lNYNPW8
C3efNG+2n6OScbNk3XYuwB4b/gbyXphsW3FsNvRYNOYTnW06HVeaNtEVHqVmDJ4x
odM+bkjysmXiOk2hO3OBtCEOAb8TM/iRqN1D3ha3oezCQqavGsrMtjb4IRbyPovv
JfeHX+fYCNhKiwgc9AcupLoGUd2BhZ23eJcl4MSQBM9iPfnzgvUyeU0FVkcZ5vWA
Khwlojn6WxLxQ5EsOQIeRLtGgZY3mWMntOWOZN0W11j+rK7uIlsoPNgzJuGUONpc
iC2GrWZRUMXXkFgKepaUjuABf5A4pxsgw2bN0ls9e57YhyeaJjSDhzIX0sA0Vtrk
TO5z25dkXqL20V/vspzrpIClx3bTFS89WFKLkMcEU9a7bvFfLQ6BkzHFCe8URpnH
dNhRjMDgD0qVzvPXz8X/bDwBlXEj+XjaBZkylILsTuTxxxiWrHx8y7u0zJN3/XQG
WQ+fDdKcYApOeHJwpsHOcjzS9tOgLHIbR42tTzFeF9kHztKwTk5YaIP/626sDl4F
yQJGpn/3tRHfBpfoIEdwAUo3phD2/S9EF2+RMgsu7UB0LW448eBSJ+QhvNSQHmG6
ee7gSRvwYXB7AHSf/Zh0sdcAqOBS+yEWl2l1dM5jzcXQ908APGUrw/Y8+lbiJ5JT
NLuC4Tj6uHrJEwATsMaAYcpsqthZQ9a65rpppH4hon8oFP2ispPfFM4UFxMRgdjv
N6ZpybPcmwXBeSE8t0wxgdXPcgb30AqskrvmzdDYacNa5ZD8IjAq1P4lN5Ms0ZDz
R0XGFrf6h6YLrF6Oga9VU75nlXkFYmj46VtoSz8zcBKLjCAaXpiRz1nFmAYXvWjK
I4rYBfEepj+FO4s+lFTLzBQPSobwtQXf+H4Tp1tarbPtzD6xvue6Din89kTe57vv
n+mROz679dXqZg5meXH97QYvSfW4JqGqBW+qxEA0j58wJOJz98MPhIsPDvbW4G9N
JZgM7WpKme/TJ5kZTq11hDv/xFdygTKzvWAmKD474u5se6/3qEdF/bQC3E6pL4n0
Xn+6pTb6oyDrYwnqqIuJbg7MYXPuMigA9utO74mfcG57pdZGq1UI2f3d5BSEQcL3
S06XMI+JxNy5WStT0nT/9PM7xN+d3zs5xutNZspfLE1zJ/+W5kF6sHUXx+gcPrcD
373iP6X2pU+ZCjqSKLwNdaBFDuMPopXEr0qBcAN6+sJOjEQKW1iouYdbC9P4PRFN
hwvIgM0h+c8jsVVP19y9UJieGrIWujuodI3SWbb7pf/r/1CWVA5whb7HH6HBCd6Q
mMTAaIkgT4LT/OL5XjiTiAkKfsxRYyMxvJTX4R77Djd/7dNCuFROkrXj7/5EUg09
6WOHBfK4hgUXjVmHfpSV0gKXSvuOXkXf3zl5/q4HTVWk/8ZcxjgX3lCtucn3Xa1L
N2uBGBYZqw1M65KmaGorEGMjzh0po7CthOQN85EBkmjUX1HddS+p831QYnK+syuk
a59VDZ00Z7fRDPW04YOAKpsDE5jdPu1y+AIzgAX3PNg7qeSJbVX2KOkNvMK/mG/7
LOdgl0hNFP5La/Vuhz/6CSSV/prVKQE2FDGHOgVswqWbJpQkBkzCKSsyau24DyEy
bXoSpcJAKj5dXnD/PZOnakMB1oXJpT6Ou0QLnEQBDO6r7zSlWfoSlWJ/jDE5zjoC
i/AiP8E2xIj9yXS5tED/waQqPz9chqpBYk/pDzZEGtfqXVHpv4EgY6O0J3XpDr7X
gbq2SPp+eN+mj7JBN8hbE0uFCCWDQH2iwCbCzsR2SFSEX6MWbQnpzZcNHiZgIw91
1+DjerbuEZbb3S2GACa675ymTCkk4EOuQqMRXvYXNuLNmiusbgbH8mLmovNweY22
TNeVtIgyv8D0Ijz7g8EFswzEs1zMU20Acimen1fCRbZwO9rjmMoZ4FVA2dBV1ndj
/WGhPraA08n/d2okxXPZh/ElIbW1DAn26inxTHVLJjFDvf/8gB5h3f5cYeHcpF/l
qKNT2HpWxu9hGLTUJg83iB8eHTqzemBO8NinNkDz6OM748KuKhkA1nM8PtvjG0Ug
ZgDw7/Z+u06BmmNbcQCh0K2vemyqkrSiiqbtUmA7Xaj5Dcd4+RHzv3V20BYEnyQY
QQcQ/24HVVYoDG29OxZ5Th2NMQS0SbZ2mLiwtSS8OrPLnnm+Op5XB0QwaNPTUTk1
t9fHGBcxSDxIFc0ybiiik6ek2CHmj9V9DvnJ10Earl4zrGTU0jf6OEB1sRV+IshH
qETGToIYz+aKU/pEStB1h+JdTj2BglW/XmlYtBH3UTJYytVyZafw75JA8TMvUJke
sGMZZLmyTHtayu5PsrmCHL6XDW20x4Cowo7OwA+jQQPBP8mGkHokZARmJ+smb/R2
hGgY0jYdsaL/H6/1udSrr2l1VqZbxlOY1XkPoEkmV+cJrnDi9e9xr8IEp5p3zZ9M
10Ug9Xk3eBYAGxyssWgz9GfXROCSEZvOvb4LfQwRiZVLhllqEizaIvdRTBmSmefN
e33dAiJT0pzwWvp9uR7XhAIEzWmN7CP35iQcMjbYfszNy/hZ758mCAPgTcRXy5NH
fIDcrUxNO1AfUbpAk1iqEZHe176wD6EXw6EaKNrQA8jQPFYCPfNkWsWIBONcnffS
8OASMLZWCMCplbVXpbbkAuTsN1z41NONjJrK7AYgWSRaaQW1KIy88KlYIZbDEdIH
fm1PXWMN0UkQEwWZXnEhzkX0JFwEMcPTY46RYwUCtblLmL0SB2KHVsRWO6Mvm3El
yVSVIc9vWfXVSM/NbTJVlLM9ehMA9Ie1wtfS4gqs9IhmS66CJzGjhbf+Pz5uxtGN
9h/Git5yGeKu7kxGVSQ5dGpVaq5rAfw1c9F1ARxESkx2/l88qbK3PqJi/Nn0G0Dp
oH4T0NhbvHyzWR/yb8SMKWmCUMiU1Zi5JA36GMuH1lrATNPNy1d+Le1zf8laQ08N
pqbpSEzk6UAj6lc9//qfXG8XeyzGFdIFYpc1HQ9eAmqoN9mjU9yty0bNzPB5Zgp8
p8AS6qZgCecglWju6wkaz86fevre/Mm06dJ+fhCh5eOMK8gBMn7RHfb/pAOAVAyI
ByPHT3B5Pf7i4iDcmMR8731K8hF1R9s7FEoSjAE3ge9zLWkNSjWXZ6XKf9iu12JH
sdXnEzS/udD0KRojfznLPQ8XbrUV/i3c9/UxpMg2DOEeqDSwV5jYkC1H43CPNJCq
S41kF40n4vN3kgnIX9Zy0T+hrToevkqQMckRCyVjl8fI23BqJSsrT6hHbiOGuND2
fa7YaLFfCnEz73XjsiYo9koAF8nSpQCrjE3q/agLIbur1E2mt9RV4aRZvvF5/He5
KX4IPLSy3hqFLfFDcruR4vq87hxi65JXFPxhSS1Jjuqv520snB8BwdjTnyQjcVTb
6U0SxFJannsnvlWa8RBj3CeQjA4YJv+h6F+D1LX8ZFl8LOR9nU1aJX/zN6dVmjla
/kKjiRSeP0U/pz+S83qHfxJm6qCPMhnyX0jPJ09X14FLcQZSfXHgfHG+deLUORym
W1Ock3iTqgksKYHcG5YYqrNLcu7932o5TmsLcxJRxKS4q0w4tOiqA/rBPvWAwiwT
sY4kO46Iia7OjbV7S7sKgHDsyyo2FbTW+Vt3eMtaVzuQxDUZhkFdzplBN1QikvPf
hH5IeBaV/vCsvkrBsdLYVjVM43Zq2Rqwp54tFlrVXr4uTtXkt8NHONHpIcCWxBst
Q1s7/BoFw0nJ4aqRUAFOAdpGkZc31l44szG5tWTU2wsgZR8fMchjED53d28/VwnU
jVHr5Hm0w6CuMmz1AMyyHb1UbQGfsW6CYovJEUdjMN1EczbmuBxB/8scy+aGHIB5
UI2gs5RlWHmj+FRlt7i8RdmQ3utH5inFRFJ13eRFNi4KDLHRdbfNTJFq2pJeUFkn
jv5XgUSIUtNepfHU1cfAKHqpCRr+EMTMoThKMEm61vTy71KeO23YPRsNBEccJGVI
OmmISv3m8OsKuTDSyWA+Alqoq2Gx5O4zNsIhlGY9/zkb/VZ6arxVhUaaCEwZUdtA
ZqGnRVAhVcEWygTZ8f/0umcCsZtLCJyFAc2gWTk/8V3YkFX7mpcVZDwC+RnDApXX
LnP7TJA96EhfMaUZNsNOdpPvVNwribnTxckh+102GDffE7VDfaY7UESrvc+42vc0
5nkaepKVcWxrYWpHZwv7az/9sXVp9xisNimEa168rbg5gbxmkeleURkKtG8T5cn8
K3skA/nVOgiUqtQ9HCUUXyHdAOsQK/G0YOCWThzkHaq62JGsQQlwCj8/Z0889oAA
rVbiwBtEX9mRj7CGO+bccKlXViqmn3fdv45AQcbMXSHNiG0XnGyW65Md4KOzBlKd
8cDi/elDo4Phy/1gBy0csw6N5i6080BHbzu6o//7XM71xnTejrHV6z4ovgJbkWZg
Y0PyaFINrG/jFQoYlAJJT8UdgIbSWZqr2J7U4nRHpLDAl+YkWbaFCc/so/uY/01T
uhgBm61KQxqCc5nKMt1k/Z2o2zMGfgxDtQd1GsMrXci4dY0wvw0bC+00e6x0fT92
GRNT6J7foWHv5zE+z/kFX/M1+bFPy+B7fow60PHC5V569S/vEy17h+lryFIb0QvO
EE/AU5OiCZQEZpBLIRt7bLB51K5mVClNjzpq16sSgMDWzpbkHUs3tpxoQpJ6QSlc
aODnzc72DA1eUW/rMiFulID+UdYOML1s7DnVuvv5xlhN126sJH30aXuFDIqqiKlL
jGSPhxNEUCC25RfDGKcpjLOdl0B71wnfK5McnMagmSvhlpqoNYvq4bfGwertwNsQ
n3nz10t1jDvyAbMTLCmJLJPAW6LirdPFZZns3/DOY+zyG6pfgSBTVh5Ndtuosn/C
NGHS8A8zPGwUxhWqZPFHeAvkgDqmpTS2FaZp6nHC7nJsvquwe4TgsDWrSa4MJwp/
YDLilfjUwLu+Ddpn572FRS9G+V5ZQ4fM5C3SHYhd3pOY/i/r/CqvFHUlf6u75Z81
cVD9NeKJlH/Nw+3RfB2vBi1mXsTReHCfQFyPAPqeM9NB0TdNXqxvN73/6pQpU1Dc
IKv3/uJ3wj0rRwL4JRUUO1LpVajQn3u8zL8hapaHTyjeox5SLZRsjUQzpNPP+TlB
wFiUsFSMDLZ9CGBc3vLNfnJvZUeGB8/EsLG9Wt/rO+7Y4itXtaBuDfSKOenaK/yy
uwpcYB/QfCPRvuuQX4yxBVPsKDRB9FXjo1JdYB5abljsChxqUhnPxDzhspKDlltD
qNP0KIz/k3E3PWnzcYtRuHw1zYNyNcqOYCNL3nYakJrR/Ro74qyZ8oufwqadkS/E
zSnNCfZtKhzCBn9AYv9tkLQad0+0ChqUqWO7M7tjaAplT7v3tjNz7sSoyiN4q5du
4yMkZmAFLp7YTxqcJqFqcd1G4POXIHdi7+h3VFWWDJhFfYuZOnHQzqULKEXDHVzk
+TZ+f0Kd0NoL2lXI36/EyaTKoFxW66KbqgHJGfp5D3GuZLY2hTgTSAkds0YfTvMQ
On4gDk3DhwUQrrW3xtAJYzdkbgdsduBEC6p5KT9/ncXj1EqwtaVOVWXSwVIEnf69
bWCgOk1DYb87qap4kUht6im+KdZO72P5EraKraXWlrWGftsvfcI2IdY2h4bEzLHC
eEa28JcU23Zww61nyjSRj6az9wXRF42e+EoawzOR2GVn2aGH8o7uVeciA/wybjp9
/egu2S5OpYN/jdII+t0M/rEgBpjCwIukaHWz0YyQWLIyvvxhBsMkGds9xKeU5OO0
tBZYWBVGUUVNOFBmZnZTzB1uLdgYgeSofpbg5Vc9EuHeACxomJsg+UbiTnF6klvI
FGZLqn4RUCYqXJJMmajsEaKxDXwY7SnGg3EoqOpn84AZ1RDePHa1/aYNr07wtjE/
PbsJu7Hw3wmGdZCdPi8RwHnbEu7diBqButbYDqHlaAYSB+i/uTolHMk1FbI9cKGa
HkmX0/DztgkK1vPkBn4H2lXFY7cvA6Hiaau2UILzR6/cp1+IpmoboRIhmBcdwuYY
MKkx1G3iNzvtbKXgD7L6K+WVI41qwX4IouZK21PqlcByA7JRA9ffWRor/IC7HkDK
CUTw6YNhoYhKkAeqOq6nX8xhRVFM4oTkyJPhcWwS6ks740lkANvvVkkcsqMJmxKh
hNYE4ynpYoFuCPAMaw4REz2hk/beP6L9mdbMBEjqGfIrwReyTZ1aJSI3bKcITpII
0Z9QeBYpCXaKZUJMprKTJm0yDmaPjXMAW2ml2T/SeRUg5B2mnaYCDJMye9rqsHod
GPneUMsoJbPIT7FnNwBPK0rLU6TqeLmTcgwCZb9vFat1Afibqqk4oytkWlxC/cYf
p0H8XL/Afc2hfA9TI9ioXaDWpu0MNmi9AqlPZAWFBupFtpm/dDutJOUk5d0OYbIP
JpMMch9OJqhp8QjLtgWiOCmNF76YelTAFZhkc1J0jwNn5mnLbhhWoO5k3MEAqE2F
LxRzJ3Pi2/xT9UqzTK/WlPee89vfzea4u2WpRnp2npGIQa8vksPm0tp+FuQnNlCh
6FvWPMH9jdHsrCDKI1Z3X8AYsNBh7HWC3UCTQgVxqdV1tEWZOubJ80ywXqQO1tHe
yjYd7dl0J83WRNkQO1+TDj3oEvcKFWMcMytX40IQVjqzLwHoKER+tE/WKwhM7qqy
4L3GZ2uZKqZ2CoFOVuc+Bk9Heil705nSkg0y8qU4Q/olQh9d9huNb+rhsAh/cyg9
Lop9AJISmuYyUw2GyA7Jps64HUe3Ak142hAxFeO+yAyF5DrZ2hFmf3N+wUi5ksOG
Fvuvhi5HJq0AhJe26TONEXCSeX5RjJyrByWgya+A7rsUZx/3XMlvk1cPHnT0KQjQ
gkoO3xjlZetLkxJMBBZQm3JdFXObZpcPjEysXP6uA0A8Qfc8NoEHhGmrylvGQbHD
xYCLRSTFbX5+HWOh931HwHfEZmY/wAX9tRNSC496xSnqf18CpVkF4NPvm9lBSdQm
RunPxmpya+PdG4gIkUSGDQeue25w9jwH2ImSEMUK/eIa5VOoFB0bkjtiH0K65MJA
M7eXeRm5r6DOoIbBDyqcMmWlphg0ryNs9OHefa0C3b/GQv9w2Wuae950TDrUJ47Q
nccnw/QbEePBOnHPalNj9M+lyKVKXXWpiWf3+VKBC/I6lf/e6Xx7lklynW3PfjjK
iD4UkG3TD4b5kWfI7Lwl9uE9+S03qIcvf2wbS+HIGiwAne/6n7FC0VEO2k1po9sC
Bd9t5TnekoDisq6TAxOIL0MXS+4PK1h4MH5sIvOFFlBvW/9D9BE/qTk5u1RUuznP
yc4c488tYXcWF5SpSIhd5I32ldLu1rNSNbjHN8eYxSSmGx2gkH0ENpQWuzwLndzi
HoGmuKtgbq27iU+Ch23tMXfl1aKwlLmPWoIdhlNFI2Gm7uoMe6ZSfyra0UnbQed/
hvxYCLH7LVAIweaPN1xsOsYW6T/h9+xlPKeMTVpMUDJp1NgmbjCXxq3dKXPTUFfh
irSsuRhsLeeVs5J5Cg5jrjedDYAFFh7Q9zz6CdkqSsjpkr+LGoUOBaeW3yCptVrx
yFkGLyJiUumEh4nXARRB7CQDvzALvoB3uUn5m0dZco8o3kmDboXGpuYTbTzOuDgB
RlmyNAFsVReXTTHgBEER7O5lVT0smD+YRo+7JZwhYgXCS34tvi2yWYwFeO4eDaox
k7Zf1qpdhR4Jy3i8P+6oqg9lPFdFvEmX2BYbNkQHkQJCIZcm6uwD98h9zSEPgoLR
Wh9L3TkgY1Op6TlFESNdzZ2JIz1qVpsI997lSY0Fn+OP3y0D4TBQE45pzVOGibM6
1K9cSxGzHF8j/s7SAvq6vf25kRgIZ44k1uQW5qAsL2heteZOhXSR9uCdzhde3mi1
czRSy/6j+P5BvuKfS8FfaQI9p8t4odrqhPFvH0CsG2QFfZRrD8PjVduw3NTXj8nN
kMZp5cPsB+bkLo2p/Ia8wm89agZOS3q1yw9T98HpBOO3tWHpqAjCiV6AhaN/qtJg
HduMlGbGjEI/3uhlfgJZ3uKnyFgsBTPFk2YhaJFr4/ThZHUcVz10+4DMwgJK+q+B
eRV9D7DnDvN0gbH4HprzBIOnM3YImwnmTjmekkqjZ3/orGzMzadAP0lFyU5nwNyt
z8pKVeKti6KTzgIuoOS87W0mDCo680Mw1e3PTOYxEGC6tuHyMh/Jz5bNkyR6RLRJ
JOhA43ZujPNobYO4MawzG5dQ3V2zpQo9EawuwogO9Qx9n/5/PMGw5AUOiJrMlkul
Q9i9/GfDcUdc5Kj2H8EOvzVJgNccW4Z+rSZbuRgphn2mYHjPT0hYW3miAiGwcI/c
dTPbsWv8MwsVNHH1AwtQQkdM0gfxoODp35DX3QEu0k5AULSyLc2nsEEXarLo1KRP
ubMqXXkPT+lBuOpxrjtvGusPEtDZUXvDdS3i62tSGhnJUPfKYNsYOeqCXugoJcx/
W5BPordi/J4bgpOZQI4aVXmvMbV5sF+Z3K0Gz+Mi1b3ByLznZmgE+/oX9JVQCeG/
gu5uXLtu6PmddLHtOvDEpvYjxmthvcSbocBgzgInUwZYeD20fYPWbjHNWTwtOXlk
sQ5ESWx23yTwqq0NyyecPAQ13U2t0/5tdfqrBQrDsp0aj3dRx7xxA46e9vLybmP/
bOmxC4lVZOBz80enG+2ObL1fV7a0wtgMXd8YJ+vu7IiJqvRrXZ5leWY2udY0cB9t
+udyWTfvYUify/9uR5fVbNAm/bAStDA8sGNVHkS6lE9BwZ7Ib19xXSaZxFWcBIgi
QNO0lp4jBhpf1DMMf/YWYA/uaesb5saYXEB/rIjHHGtt6eiGxedCTEQHI9bIVEZC
+KWW+ALvNDQs3XoqeO8NMehx5J8Leioys9CXE/WUZQkP3/i46YljJRPUTDEARd1d
4MrdddVZnre/N6Fgf3FECGY9/8ejh6d+IbPazvsSPcRes8iXtqlcV3ih7bt5SNrs
+xM8pM255D1/Lba0ju2z60ev5xrrxoAQHMA+iTnh61FERHKLhXiuZlobno8rciyr
cxrl5VtvcgMt4tmZY+EmgKjFDPsQlJkoinb8AxiTVkO8B+55r+wqtJMqNSaEz+Li
3KwxeV6Hkl7sG/jM9iYeg1m1JMoifG9VATNP/NaSeGD3k6JPfkQhVdME5PKb9XNo
LX4QiYznWuhiSNU3yCO5H7xM/pShJMNqsEtJ84Io5X7aSRTDNlYv0pPEY91q1bxL
jT3c6lmqleDmvGAWxpXxuHSmIQ5ApVbHVEZZoYqJ5IgrigVkvW0ewjpzoXuQ5Pss
6O9XgvSNmNKcv89hRmKJvdSPASuRahgkHQfaoxRm/5ZasHYGNWVyKJh2XTk7yPAI
+nFUBECmqcF0vIdKI8Tqpj/G/ttQw7ALrN6bxC1YIC3SR+QWRREuJVsz4RGFmcXK
wzaBSGpchPitoyFOpsOoWP17S+T84FbdEa/8okdD7vBlfS585RR6/57uGHtS5gcW
F1lcKuwaP1UbpZ2d3AQrzBLeR5wvvjO1f7h7Dbg6cJcYoflrpndW7LcTeHko0+uJ
sh5Ru42z20+m8Lsx28cq0vsgKtssgAquFL9ZVZpN47Ur13/jKILQZzrwqRsx/gb/
NH5ObLDGuZ6ap87O7cK++Dr3J4GjE5onYdqdIUiOOOsgGpQEdtb+OjfNyn9dLN2l
P4hy6mfKinAy4sT/flIgYb/qmuq7mJ5VjaT13LgB5y4ggBwkomREP4b0hENuygwU
10xRSoICnbqegyVNiVzyr70XcS0Z2VR68BNXvCpJ+bu72nr3kXJXW6Yt61Fs0flh
r4Y/Xy0FDnjXf7+cpI4X/+UuqCPjt3P5MfS9SvQmZGLYu/4rSqebJHqypQ4Gj9im
Pyz3SR/atBkWt9Q7hx030n7n/J8NlYSZ4J5RRhU8ajesT2GE85yTvX460G9YPtkz
xD/AxJLsAmd5hvtRaRo5kgjPKJ+a1cFF2XO11jyfD2qGydaRGuS7ZPQLplvqdZKh
QGmpPXNoAUhIatMywSTeL6qAHC34qKWB2UpDIriVK6BOqTfALmjiNV9hm4K/azjw
q5L+qo5C+wehswnqLV8SsmGGDoS0g9azj7HwPcgTXNZQob/haEV1UX/KseTa3ytc
0jUNwvovr3o7BlXhv8m55U4ssid4DGfD6XhxYeeOw1wpDuI8WFL6CgcANMKc5WJP
6ASejGC0Ph57xXztKcyyGlRx8x6K2sfU32u+E55ZojqULfvMMGQqSosAT1x7Yqa2
GrIfM3Uqys/sUXV1UmMOo+E6I5/NIZ+QW2lOABFBo3KKduky1RQvRO/lNaqwddJu
m01McwgnIEcLAFhRuvoKLsjNTZb1x3FHBF07+pPDZx516HknlOCmJmoPjERMbicZ
0cajZ0ND8biItM7hBcbjn+9T8Y4sdZjyKh85u8r4JGe2maFThsn7Hq98J8L4SGdT
2cevE/JQXspve7JNKPPT8mhyt2N7KcZRqA/vneytSFhI+XKP+TEMchv3msGGZryD
A5YgCnGzxQPs0LlekWp5NYZPDrEtXUJe7A3sF49w4F+nvxg+l49mYeMB/RhPs9EZ
j8CQGOFoDU9ftALRO0ibO7pFU1Sjk9a2DX3r9R0BQbpEgs3Q2XwoH6XLRgRDt3Vj
ihGOQR7wTHnsUoGhdREG0BPLlAJwdrdpwrPPqgaktXrdTCVmp/YiZNoIEjQP0uWe
LxizrKgh/rxoE0802wjVDaqzdckDpHKv3D2gVPC65vTp9bMzUUEoZ/bb+1iGS1F2
iVhPIkBE+bBgCw7o6kCAnrxBW/kCSVvkcXmVEfswWrShyLQPb2f0LbHJOYBX3TZh
JlmRQ2OjjwOrFZNraGXYu11rPO7KZSxssG/vdG9a4yiKDr2vUMXWYDrkfoU061kg
f2eGPZ0efPMKy9OaEmnuYaV0/xlXsRZvnX9AsgJT6amzn0zZwJCIFPn5hjEsYqsg
xLV+pyFyZVja1fmTzty7PwkgtzEVOLZ+fZz7jWZjSmS2Wkfml7l3031734033lBe
j1b7anybiwzhlS1PnQD97PiHPgmgxjCPlyWGkXrhUHP2gyud/tvgOCrn+NerQT8L
KqI81FGr5flk0LJCDdc8u0ssjib3rFmKtvm+8FGCkH8EOQSExf0MZ+1BZHfb0g/P
4OrBoiVUiQMV2a44j7nFYieMtLGzC8VwRUz/USIZvBbGa1FNuJxSmanNgZvFdP6Y
vbdTxVpD/xZn7FwSYTTczNhGjbd7++a11nwKf1s9enqif6Hh91kqoYlhqMkYuDt7
1EAoAwz1vFdCtPbcBMKQvj8yucJrO/nGZrTkzkrsOySIm8Tdkgs5atmEQkThoIWe
8lBdaFRVYev/PpgdnXA6bg6yY5/9oKg4LavPZVo8p5pM3aD1pZQMO9mO/xrXNRdv
YcpbQr0Xk/UKWFL6Mn9mFsv5tPrXVmq1cDmZ0yf8vt3btyE4Z9f+P883fs4XN1hR
g8qcFjuB9JKfeliS3iK/+Gy8BEOPLd4XCJi2XEoRhIOUNMfSwpkv1T8yowDXbUN/
hnQL31ZROp1pKyA1ZFoclkcOdD2fqexGyUclgQ07gJyXm95MOoqXWSCzPzctkfSx
va3PXAZDZ3N2gd0a69Fp582KPonyDnIL7f9C/QijLiDfQf9+XpMkq6q+oOnen4Pt
/fQdlo8oYJFQv8oopXMBQJMFWNaHZ9cCOUCW6eFo+CorxhKkcF3w3BIRFgsEGohM
Ewb3wY8ctxPTW3dT6vXm/lkNoXxecXDG+tUMhl8ZEOw/la63CAbkSW5bFbqvn/xI
Jt7/loYs+JOSIlW9wF4HxQ9cH8SU5CO49sXs5g44mTk5pn9p/gVPv9fKcu+KF9Sh
C8i/TqCV5rOXtQ+gng0+ODpn3UK45j2YKAcwPyF+wPxxiVJT8oG7I6NCBV5iIEh9
F7R90XlqwTpNmP2TgB0eog8h1HQhZRRzqD2ws3L0m9ej7E31zCtdCMc78Z/1EE+l
Mb8mwuDRcO8rIXN7rf2UmUV15CVxI0h8FBpxaNshlY5/wyz3JH/kNs7GiMnIL9WG
GqP47PxtZiJG/M3an1/xrQK8PEFz3njcRdpop9CtfX5FvV29EGLNMIYK7a2yQhdz
4A10J87d99aW5X/2O5YCuAfCD07vnT2LYN+QfuKPEllOmd67X3qd1/Fnz/GugNRE
Abl+ArwJ+6n14Me3cVQKYgo2O+woCLYdeefTtibDL7FJkNOxD7FfrECuwzO4B1nR
1Ykm/kPkhS9ObflFO6n2B6iaZxB/B7QFxxgdHR5L0/rNFud7PaSiIrZN7mzH/WPV
wt54G3r1dx2O51AIBEpEC7Uynm+GMJbumJI8BwTlXv5rywcICT5M2SgF7WUk8s/M
NgOQfb9pt9m8VUW9g2/6u51c7VUcly8x/bI9dNFc3Sb6Gars1lnxDsN394xiNj87
0r/IZ1MuuWDljs/RvcGL/HymPjPfFDHZ+80sLl0SlM6NL1P9VonGNqcYGirWuW7m
YPLT4nTgc5UdpSGc09BlAite+CLwDJr69WFAeK7I+LnSObCS90yqYit9/0Vgm3Af
dnbFpY4pKfSa0zGkwm1DyZFTv97XZ1++JrqdZtXJEVE1SNNaIXB1knW5nCK64n9t
GQD2QUZZAmzJROfRNdqT3iNncIjII1JniSzDx9QC8g4+OXuDgcOYFQJ/153YkIuL
3CMt/S376AaGWeIdm9tMULlnbCFSX3A6YlY3lMYb7FNvQMnHD0geVyDagyWXBMP8
MXtacXRaZt8XJMbNc0GWr/IhqvZ2OR/XzEefdhyGzxt4EV+G/VSzg6D48rWYuLPh
jLc2MNRhCUzsPIkT9vVEZcGXl0qfjVck4+RuZi0TFK7trvMt0C54eOaDUS9pjkbJ
YkbpfSAemh6d4W/FEGXvVDbciNxzYuyPEXr53IUpsr5VZzxF7vxbl3kkDnyF/jVD
h8P0tiDZ6CWi5VRmUzyQyt5zUOdGX0HIqqFStiRKY/4jUN8SHL7veCuhhPNQt/Dg
wXONCYBk9IPyRiafTBtRHRINgV5pwT7yTab6WoES+Ac6vZy19fQlLZnOqbKr3iLf
9v03OKEJy2nDV4QdPESOzkb6NgxaD1920VKQ/kOoQhJDDd77tNg8cKhwEYjxr72k
4RNNvENdIWvRssGqaU9sHxIZ9RPg6BZkE9CQiLx/zK9WFXmg8jBAxDuQAwzkeYke
zCL6QJ2M7nSLGCQibpyoMsnzp2UuL08SOolr5kYgtKTuNGxK7kbu+pgHxYYUZrep
U8XQ7QDv6bK12JuEPbgmeIQ0BeVLp6wMotGqiIhlZXHlhl9ZMqstc/1YO0u79Z+j
Ne99fSACH9u+3dDUEAeQ2xxLM6S8r3X+itmLUP6dEcU4M/TtjKD1VYOoR4ghWlGS
kqxQXbwY5trze8He3on1dpuZ7+z/WWrSfuyynI+BAvjXRpVW1QJKcOdXonDTviSS
qV5moknA0YtvfVYTFjMMlJUOrmUQ/AkLKGNdiNXNA0RFseLheWRT8dUst/uzF7vg
Ile2JvV2ASgI61GuLwZTW/Ras5s+p+tObZveWqu+P456EmWfDWL+NNJN3QnrQXe6
jFpNdQ/VEG0tpuPoXHmZIZEZ1DMHDrY1nrmhdnBaLcl6a7l8whG2SbBd+EDMeI/E
aWynrWXep89x3VykhrBOxgk+Sg5shoWprmFn6f/7wL3P6lUxPyOJVJ9zVP0dxR9D
nc2fZ3B+jgU1fTKDIq+Nbq3gkkBvZeKr+lmfUeVEnxHH/FmCaV3kKJSCkn4RQ6+i
T8euQVMTf42WPxk1WsGGUcPaylzTGXIQkxjQKP/2jXUqKIqOLRf3NyOgyTg+jaML
eG67zHYzOmNtSsU4qEU3ETjI5huvBbZT7JDvaz5MUF9PqHdBaNhaMLNL/WxWTEOS
k2pMi9PPlIdq1MxHen6wJriRlIv2lzCHmgrVtcMK/VlJnh9JBGrINZEKh9Zs+byz
uMQQoPlt62wlz8QCII2sJ221D2Fw4iOV4sZNLpgSylKc15gaKRnzciYVQYEGSRf7
eKpu3sB3YVKJuUmkmIb7NS7bfGxNCweLuCwr4Ro2vfstfCkK+kfU3D1tjun/mPNV
8I0Xty8UQXAfGDmZF/UXqJg/dFL245OvpZTKmkGgov6fxvBLqPac5LYlzKfHjYvY
mnEoKbfqu19Nf3JOvqmHohu+rGvIoEI9wfZa5Ct6i42gxLS8YHhu1KV9t0dbxyUz
SksytF7moQimF34aEO/Ne1rpnVkpLDctK5U6ToVty2g30lDwSZw8XfgVlLhDHiP2
89qn33Kh1MxpWaC0+mVXGZ7XoPZZk+uukr1QSMKmJwPCu6V0s67lAmnDPMBzgsI9
B/qxz3jRDNFahpKuam9zfJl3Kb5U/atHO3faeESGuypwQwa00L3Y+et4ql1/z4/E
dj4E6gg4vw98t/j23uPQkst+SnZU1w9oVLsxAm7tkxKk3gZ0OzRA1+DbowE/qD/L
xosnxql31lu9xOx2fqrymnF9Tt6yYQXEL+7o2QxZRrvVDKzIktJuVM0hAGYcg6w/
9MYTk5I2xCosskbOnWbroU9+K0WA4llKr1VbghSBQUms8ZjMlysohr93dQ9yBYAX
QL7RcYWFYV78+BcK13f7EXbrOAvqioxejuXnZXczpezkp0ol1doPKFeQMQSAM3ZA
XfZ+zxWUD/HWfK1Lgd2v89vg1PkqHqTaIFl36jH8azEE5UyczfN7LnM4tEKjyVnQ
YGzfDrT9cPNcOSssvqUJg/40pE7tYRTZYCa9LSmKoRNeUZdh4viEwe9tz3b0LzUW
5eriMQIPKmshMhVlcRoFRgvZqqfA4dYPFj8AQAAuemOBxVuz674+KsPn8r7FUfni
8JCmatsrienTyOVfXI/UhETrQPNion7bMKi6aTaQBM9upv7ofijtNJ9OMjAJcZYQ
Rh/Wc9Y8/R1nm11CMq9BacZHnbHt5xVj9srCbKrVmAbPWuc7Q+iJ7TJHMyR7o+XV
JU58mPhVOzq1qLE8VIxeWBuITj9U/Eaiga/8Mn+VdJSyRauwdyc26JTm5TH0jg+Z
vXka8SAXqLg1Z7UzaDDrXBsLtRnEgVgCuEO3xBlS7u9djXWIHl2KEXhhcpBRQGDO
v5vnyiJ72MoeJPE2AA05ztG+S9JEewfcJNFGPrlK2JSIIx57lec89OMo2zt8dj8j
FIy16VpWsCxcHMQOgz6FgdxMJ6GPXf7jukfgSZ0xKFc0oV07DQwD5fj90kK7jyOh
fliHO8+B032SZ/y3V84r/fJLdpLimBdd2Abu7VM/Y5VpT9eHl5CPdUB7LWx/1Qtl
lXgQj93f6F8UpYDGy6EixVG1Wt4K/sor/4Zv9Q62PI4khP7NZTJArirWwxv1kA/M
hgf8LxpVnxab+O3k/TxZmUxIf0PDmeVOTZVjeYC4YH7jJB2jOUDEX1oiHR0aB6YA
yKHWKNjMNb+2sn9ePrX+rSwhwWPwoF4191sNkVdahsHHLIMelP8+xvU/4h4lqpl1
iTYF9SqM8H+qmV5xBEdLII/DM9ykl1yzhx2FlQvb2awYH/yVbH/xCCuf9XD6nOzZ
ubfjO1PrBXb5gGAvlcDszb+BqM82CCVTNawSu0EDiTU07cvr9E11NDN1sWIZ6GLQ
gxnkxDA0XbSEfD3fGDMaJXEZaCP01yaA3NVzs/ppzcMLlInSGAnHIj2EUYnPVUwT
3bwy6cJdFf8TTChmSBDvs6+6AoZYpMoWNPxkWuQfrOcoCCu3v0cz+T+sHbvst4ZT
nmNHQlKICHL43u0S4++eIDxdElBenVDjhKE3e8d0LOPTQfxOesZwG+tY9lFyVZAj
5FohE5PNrmva5TH4SRGVKwoUSYoFVUxa3HEvYZhWXvp/LrFt/B8a9+asNctIz0uW
xX8yjwAuFq9+N7Zemb1l49vfIJ1mn5FHQt0rq8wP4oO6LoZWb7wZZhfT+LRKNEUq
bA1ZBcRdGtVvBDYAgC2D44FtnBq05rpMoNjJyhH0yv/52i13xQdvDs5QTkk/514z
XaNtJTYTMvUZXk9XGQuF/EK4Brf2R0+t1CmrnOackwpLmU/OodIUzrafhEyDjzrh
PChH4hzMSlUNZpKqLwWiO6Vh1ONAEWbWd26oQ5nva/m9nkgMqFS8rSdfGp7JiLJi
2jz03Kwd2cLJ9EKdkBAw7emWjmBefRTo5JMBxLWW1N9a1joH18VH91hRYzR+Drhf
U8YBZRmSQfxUEt2h9T2N9C8BxpYwETETugYMvnbfQSbBcHpugw0efv4W/sqI2ElE
HYSM1h3P9cH2ot9GkbtEHOdmGaOOapwtz7dq/6xtyklhrCnzKe6udEWEuAqp4O/Y
EHp+Dz9Cp4TKI+DAeQNqZdN1kDHEeWaiFjUFOeMJzUzJ1QdmOkhaF6Ue8/E3IQjc
itzKOilVhp8v/gGVbMaKCGgapICfM33xiIEsxpF3FQYTFxb0eC0VbWqqkotSlpZl
oD00J6ZC7FE8JqjR1AOsoD4hooa7E2ebN2ySadnVVbLXSJLCLeTOnD8ZiHau12uE
GcNP7wMqr5IDvsEarYJiQgM3UP6JsfYdraOBCct3tXrdUxGEanPA4Fv1a+wL1AwX
IagdWMjRzSI6PWNGOoFWmzgeV7a9Lp+vRyWc3qoqcNtVvzNRfmjlYJnBFfg3L1DZ
G86vtNyx2RMv0NcxtxpHOAXbVJYVeqFlxB5EVyn1AEy+P3++pNZAiW/UZu3qcORI
rro+vsTBG4UZjk1juBvMnPrZv85o9rHcyUTu6anccvTw/wuPkqcQ0NV3cOyAYWDV
IeNoRkEWklmK+6jM3NN1a05T2fUZHMQ37Fr48uZoLlK7ynID0XVp69VZ1ORbKKfJ
6Ak2Rt9X5ApNBMWL88l1IiqCfwxwQfU8ChKYScSFmk9GRdAd565eRTVAfeI7VqMc
dYfGBe0VsXD73K7lD9Uge0W362racle0bk1gQbJ28tzOHe+nF9vlqsqJiTphmvOm
y9680mCYxk/MxA4THwkHVzau1mds5K+i86vLnVd8GXJlsZA8cwYZUDIISQdQyOU2
rFCVUpqTKjFHUGFuGKzIo9E1IkI+J0lhrsbfcw4VJx3M8qq2gUA8iTq7PFuPXQii
tWnYfbouzlE3Dv3lqThi7sTwv/P9OjtnQf2GazcNZOProOAjsvncVTLYY2ttfpel
0dsdAZ/CJgqFPqTUTXukA743ukQr1T/khRRmdmtcUm5n1s8IQFb8ZWkQ3Jxp2jbh
oe+QDTeJJd+CV1HpxqAFWqwN0+U2soZpOYuVFXk4AK1mMlxl8T5LsPIuJTAZL8fS
cqolHpO2qvQDoHwwP6W6M/6FrfZK+3XHUTux9nVKkj3arB/qeBmZmUKUrVbfdiY8
wmQEBL762KrkonuYuu9ED27Tya99XfmmG2EF9rLQU5xFKHnidxPH/cTRNHqLcdHA
53OhBQK+csxnPZoVZ6yQsuAgHpdGMjCO9Iogvx+pRZi8+ZOFSdtp+8Ot270NO8oL
bqWvsq+XLchk5fYHYCK/H7SeZafmo8yJZVdbQQDwAq7uLKSVDd2JAd4r2fITPgN3
IHT3I8mGz4QX9+REv+1mtB7/VuANdmSJHvd2zky3gls9ax65Q39FPZuCPmXwUuVx
gia1dXHVPgp2kI9oggZQ5BMXU0516ZLtDSnl6wZ3nyPwyXB7QZgBgN8SfYfNEYkM
lSMsFFRfwo/iftQjio+cjZb/7JKU2zis0KBSgJGlcRvVSAzy+LqSwRjiVO2JEAH8
8GyEkFKxoQ32AdGEXyFUHGrlTC9nRg7TQLksMVtS/fvpzJ5HJLuEMOsdSRmY1Vd4
jr80RXKCpBpsn8vRoTb5x4ynfCQOGgej8e6DVeNLOBR1kb1UFiIfVdeA94F7WKsm
bIoCNrBPcKU/dQS7OFY7jLS4uR4XZml/NA5Zc3DLkXd4ki/rEjF6BtcYpovRM66p
8pPoYiCBhte4a5GSemF3V229h0nbEB95/fxPWD2w+0tF2iGQki7fARixeqJ6bJAV
2l5DxKBhNZ0kEV6u9eOOgEN9dTP7sQtVX2ajVXZXmRQkNS0jgM/iJriOHvyvu0PA
2qTGV4ix9DVKKlYniWNm7BBFLXk/0yjejEE8MIt3WJSodN1U25NFnUwzumAe9ScB
YMi/mbTe3ahBNyk0sjGvRFQmUmezRtlZqMOAQo132cVaEBEIg5V/XWE6X8Kby32l
0f9YpTR+oh1xnGadNMqsWsPRY8yBEjZMdrOBn6N4qbe0C60TVAo3lSe4iA+Yni7L
06WruPq4xSGUZtlQchmfP++BE6dwLD8oIWfUq30GzNv2wYOpErRWT8/qvOPWEmTD
RIAb25rUUMAj/bx2m0dimf9JZ+KTk4PluSf0bGVYC87Yjb2MmJngC6kNQu2RlA3R
7nF/ivivy6C4ehOjFKFEzRN1J6QJYYJmlRPwvVJfr4BJh+kqU6rgO2UUPrRl1hoP
UqHxJrHL2smlfB13dfofrDK96lOQb0qGXOCKTPoYeJged45R7TLcw8yJpNYj3Yk1
Jo9Wfiwap89D8vuXa1dp0u5HC8BwWAgwROQ1Rv+KC+c3RbesysC5Nx8tTuyoPJJP
DThZwSCPU50FJNg6VBcuOX8AWgAg3KqmVd7Guas7EragS/Vlr7Dj7f0XY79zRFGg
LcGz/EcYq1XEYwH8a0wZz4RP0ZmrPGAb6HP9vRgxortPRl1tQDLeS7iD0LiAoQeQ
pbSFW6JwBRKNCK7B4khPda7CN46mbT3iqT96T9K9mfjuJ/jpqRTZrqazfoQMvsfB
xXO5ls3LBdX3oTJXjYPFwcbkawtXH+xwqkWT9FE44S4MOh7+DNzvV5E4gu2Thigq
k44Hw/9nRL9i7yj4hbgWT5HzPHJnaolam4YN7lCqP8rE1mX5Iq5UKjvLJdi/Ok2U
jajGdpmtHoOXZOsAdrSZUGe3V7Vu1+2Uo/iN4Wr4f4M8l0LewPilA0QQw5PgEhFN
jLZDqZYbg4LQkkRqu8beIj3+DvWhi42wl4U64HCaAO71Xq78JYFdQRJlXE+gmOR/
ft9uKjjz+2h8iwEacBQEIcRulj/QHATe9iO1+27I69Ok9uO/S0vMM4R31MQFH040
cJbliakRFCxdch8hrXgvVMe6WDa4BmHEHApt4BXsHWQC8eIf+Umd1NNYMrpgxuSI
Rb6QjQIQ8rwZi6icjLHis21usWv7iFylD3zHhQGp8Hm3+lnEOrrVkSDhupXZ+Pek
eAYbSpz0xG0X+nXXkkWgVh86v+YOkZ9+D/4wlZ1A123RNlSZEFfjT1R1uyP/eqqX
22gy/xl0ISh5WBBfBDdYZFKdjBMGa75gomcXoXHMIjmuwWr/xF4jF8Oj7L0LRPLV
yIoFSbLPgjUCKQjHtJpvKnOrijgTv6Yi3+bgzNuvRH1CUZ3LJMGbjD5rQjwp/qzm
ejztLX8sSCz34f5JFsWqRjjOgCvDIrej/O/ITr8+YZEhPu7Cd29B3P1Bdq4W9F+V
0OSwytTyAGnHWRaexg2wilmENFsda4xkZBxBD1jlAOiXBasPywxcecC8X0Q3jU54
QsxXwvPl9okBRKpIOPBgLlzegCg+T/seNjvDSn5a2d+0sNurxMFmPcDXWcDSF5z1
Es0nOxt2lIDdPUroG6s/kfaMxEbK6GgXXR94n9cUJzzYOxo9nTv0CzIEcgTQ/AOh
CaalRT0hh40WVrr93s+bo0CURF+gEed88C/8NSW7We2kSkZjSxKWQ0ZwjLuY+lf4
fzeE0kHXhH4OstXpKszxPT0NJOlMsc6pTlwCdFyhSpHrN50I9oyNuT2VBC/f0m+X
XBkpvl58iNHRIt4fYhrTZoBT7mJVXrMLL7eUrG8TJRKrU6RUA1T66bDLPqG+c8iR
VUn/4R/WXiJveGG3KYng2rJ3IOPGEebqKlI6XrRZmfA/j90XRi7jhbgSt9HkU0Wm
rOnKipx7TE9EKav8aJg3eC+CBA1o+cqRd8VHuWWJNmQznlz/x5FfPAGUqv905siN
i0MkZasLM6uM4oaffjcZ7Zj+pPG0n7WcMF8hpV8gZ/upFmEodBTohNLcMDtt/g0+
qZ6/RR7eBd/GZ3P8Fplzc4dxUrBHNi4G/DGWYiGn+rQAXTFxXhcUJcylg3oylSig
w7sfH7VZ3aSbAKRW+vDal/zlQgpbnhlkwFR6pcY7JGF1MxiUHvIiP4H/Kkkgx88h
DBJ4L9XK7mNv8IsPhgz/jmz6MXQ/UZWHRlBwec+yInDm+Cvvh1bTS44Az5X99zLb
OAUMfkWkDioYeJfc0QD7zbiZPYNRGgNx3Hv6SU1zXEJOc9k6oP2fXIH4Rjm6ARX7
B2+Wi+ZXlvIHZBPDb/zHFyZvL4TYTx9z0YkcTMu3zbn30fT97euAwqkd6XYlDzja
sZBWJyNmYfITxPcG02e2dkLBH4RxqFd6JtsUi9gjnNCjW3+xbYUKP0xm05hBKuXO
92oxoAfmNoE1qNFoYkJwGxlyy/5FKCnkMUS7BQVinCqoXVKSUXj9Br4LG1NAqAed
LTRhsOhoMnVRcavG9BrDVAoHIN6yqK9P2j0qyQqa8ReECq/K71l+sH2AIMa8yhWt
+GwvyyM7w3mLPDwl8F8k96VeiLZPi9FnPHpMYhBpg2xwHXJlJ5dpzTXBlgD2Husl
Whak+whd0O/tvTUA57nP8Wmx668N7N5ix8IKK7LFRKmdxgJXCRb701LKAwsEYZhT
Fg6PGYsTCRVPMhGFPhYZfoOHzC3V7HMQ/ioQQH9MvijVxMD395rvHYCqbhwp7o76
662vaKtJgLYe/3AO+qLGOTNZCDtU4HO7waUuFSGFZLb1PMZWE3LDDucNSq0GkS3w
GtjznCYoE//eiHItK2jo6bP1QV0M3BT5Yucw2FjruHBvoE62o7xmAJq0mFt/TFhn
r5a+ISVLgcdeffaaduXgN/fJBU0zF+DR+fsYGbi3D6DYT4lYsmVzXyMpM2CmZH3X
0CSjpqZLb1VSsX3A/MvV2AkJVLMst9j1G4y3qx84NYUVjT7tccDkgWuOjYoxzOBf
mby+hIzh2Mh9YFSsekMWLg0I1bXfGoIGds0HhpaMHucHPWUR9bA3Xui6ssXoTReM
+qyubCScSMzL6zdZNSgt5IaPbjGRHkGJ7kxM2VsjWh0aTigokHB1VgB3D6BfNeFr
A5NZqwwX6x2lWuZsDHk5LX6qwbfSSdPIid3gBWtqzRaGrOagDVeX9br4NZZRWFus
Z1jdfKj6U7cW/FT7XrsrZ++kosE968Qu3j9nE0oM/nrDOyD6JCVGh1ln8DBpqHqy
yOHWRHc1AfcJTmHgyyB0DJuMrw02RFFFpfGDmBDRXrpyhnHxQitnitxWQTIBQHJx
+3oCQB8cvRtEmUzzTIfYc0aoexDGeQy+O/KtPtwn72z6ltz3UkK6+FfABRDURHss
4oviEi1WbTTvIgTLwFTLNrrMOZ3L4aEwdQ6/467X+HJSuLJdZjOAfc3xsVcDzahZ
6PTca9NnAK49mocULOyDOHC33iuf0K7Nh4N2+YHTg/7qozbWN7sPNXAhhOG2s32v
h894rivM4LoD3CRGKyHVSrzshTTvtZy4aPNuLQ3nhwfXVbRQHE6sgi/pNjfciGXP
G75hLzvV5Vuour5YNR97bMXeB7KE58an1BL4LpLVpB2yn5wlBMDOrqISP76SRa9W
GLkqNL3V8HJk6+HYbKjbTUDALxNc2MwzzGL1EGkBuKjc6j+155iRG/KF/23vPMp0
LEJzYOqaTvRwGvCtd9J7LacqKzRZfVmoE3L/yS7g0bluizbnlEJOkwjxrLRb4D62
UM9zWNhRFS4YO2W1fBrGn0fSFmmQtwzj81oZ1a472KhYvHoHDZV7urwwnJXbnFUc
I9WgsiCb+DreZepMA0b0dbn8J2PdNDvodYAuctY808460dfq1z6yXWfJ/N6aEPXk
nMXO2j7LP67bYM7vBOzBivVZD0gqqzyBoKxn7rDYZSRAX6PYmNPphjGSuUUwYSy2
o6ldKu1E1Y5CRuyXQSuDSYo4jdTBZmXcacHJJq9aCaaoTWaVbEyfJwV7wHuyyhfw
GZJ1ydhLy5rfVnQZfGUrvDge/Tbh3a67j6aC9dbIYwA24Stzl3JbvSmMjr6wekv7
v5GErhXAU1uidBWIPDy/G0yFKR+HbQ9BD8CcRlY2jQkDKqcbaO//IG5qxHXMEGbC
mKR19qO7z5iIkpezSwLHwXCffJ36GOUGutqIW3b8MTLBsAM5GN176etsaGdt+EGb
6FX5H51ipyj9MmS4IhA3KYnHmWqR07VvPFyRBMN2jVUZW8P5QeHXo0ttOSujUZIw
Iovjqsd1Hvo6Syt4cpD00NEWZEOGohNbUjzNWqyGGFcxTTF0wF1gxkyC5DE4yuqX
X/yYQCCu1fWytfEbm+kyqx2U5OwrL4RWasiFSQ0pCRpMZHbDEkB8HG5tPYWL5Sqr
v9RxC8Smc6paKdn3MU9xGuw3pRZw6YSmlGDdVuwGKfkwR6URicl1yBsqlh/yFLRj
LYzfJV6RJV0iG56MiM35mMgYFGmK4ptD9NKSVr9d010W0N/hu+CqwUr66OALmUWk
5iShNdkeVC/crdOrD5J3AHoI6Lph8uMAVJzcCWarxfOIeuKfFCU0T5DStu10OFPF
MdzvJLEvizBT8FxTFh/H7VgBLxFoSJzqiIJmzo4RqdJq+88w+WnXTPMG/63wdfHC
r+7rPTmkdx+5DozX47GKF8s3BB8Zh8uam1r1+oP/J++rQN6IT7eprlDCFxeldXSc
MtwcqhdV9WcEtjREJFYBmQLOZLtAulQsG3xeyl6Pu5djFCx40qQKykf6XuGFpJiq
nnaV9NH2q2RhDBBVflkLh8pohJDMLTIaxvZ2xH9+uhHO7v+J7spk+P2SD40R4WU8
APLGBgVkgXS//EvJoA1Xcb0b583cqoupGxF4fTcRtYmbEjjNnOlV2hEVQIET6hMy
lFiekyURHDXh+4T4D3SZ3wSDASPTKmvMkdgyC06Xm7e5puhaeEVMue3dVbww/2ZZ
gnwKmvQ+jY1hhX0g+2qzxS4MSi5RluwL+u3cY0VX7zVLZx3dxrcxjYvzoXA/5y0s
2QHNfmkNVtVqtY6zVSV9pRpAc9IJ+UJ6m/HDIobOQPqcc6fb5D8P8BQ/YXPXo7YF
HHLZzzqHmpmZf+mwj9hkDLy8GoiQgcXMRSVioYh54MJAV6edzmT710LJZQmLqPV9
ujbc7h+534Tr70To1if5PZNbmddC938woHdOT7//xj8sE3WGX8kOR5YOzH9muIG9
CDjgu5PzYvomgYLGFyNiHlY8paDY3oyUWxoHs4IpEnrUspa0vBsmIrBFSlG9xVEu
OFglf5YAoNzsnt20W8l0IIQTYqb86KknKT6vFXaQbCegjFTIrZz3E7doMh9fdY6z
11h2VULw+3AWhLR/pZUbIJiDqxsGkM1ZjSRteuDrplkYyCk3Dcx9yi51DL6JeXTQ
crFuWBcqY0ZvGfmG7tXGw+IvLgElnMfpk0m5/6zp6+VjTaqK/uJm2fY7Hf20FyFX
XjKXSPwgC51b/2zNm3VbTxYc9DID09ozYHOY3dn0stNcS7Q0QUKmwM4J5TFGzmGq
+O3mZgY7D3XdtLRrcSMKX+X10jIji6Xx1/Fo1HT5XSBKL3ezVBKUBCWeCZw89hbM
goIeYpPJPQthRPuligMc0Li1r2HXUOV7vajwUBT7vJ5qkkvyR2lnQYqkw54wfreg
uHnUMP5M5x4N+vsSKrq2AnGPN5T0ZWtyh5qRmx7dqQI+LOw8A9l6Zx7Kwo7hr4Do
V169oyNH4+LNS8Gv7cwFQThg+DBQXq6qBpWooVbmLmomP/YuHBNpix/SRuhqhp3L
uC6H2F3yEh8gKArTKf40LAtZSkQoeShRdvLquJD7cp7zfMWf5nYWS6CFuqlzwIyW
fmH1xM0GOUtnKHkD7KLPAdwMehumxpMOgMfH9CAdgKwhbpuF/6buhcNu+4sxUJky
NK1JXFTTt0ErIK7jj5kqWeh/FqifsN73JUBFMDqTnoNC0nC6lkiI9g/CGnAeFOSy
gtg+xXeVnvQjRX3w4rsAfobpvVgUuUtHf/HFjgZg4sDD+Zwxgh/K+6MGcAYXHy++
xyBrB4dhHreT7EVkAO8O+LbhxPSkAUj6tfUwPIdJyd7fQvWF1IvhT10thYB8M6nB
ndLWQg1gRcHYlDsUBnIWrrOiq3nIJh7XMUS42BX4WhP+45BCiuNCtlEIkGITnmFp
X+S54zAaYkPlbnJsP5PWagLBhFogQ2KnUzeirEHCDH6YhuXQB2/URxo1916O+GQF
l5khx1YXhxP5tkObvYzuYizsLyrvw+FAI5UYxNevTjJ7oMTfgOQXB3nnjjOuFAIk
xk2j63hpuIcUxH+N/xAgO1ipwXYBjugXR9H5cNA8DkmJ3jewqkKE8l8GNrtj/IbG
89m4RRoo6YJZgczjQyZ0vEKY+49vYSsDbqP+4HsrYhZZ1zG2o1ik0zVPRp/PzwFK
sIovBUtc5Qn/qOobNB9EzEVERj9BHbVGZfJ1EvTtkdqX33h8eRi6E9e+LXBWh2DM
OoDSzSLRjVNmFC3vNM+cz4eknKNEUYG97gg4r7NbH/0G5ztjTdLz2FE3NvRQhtBt
PAK3wBBKcwfkww8QnidL8mNWNRSAdLMqqsKE+NPesSkCwrXKoBUokBxVrXlx2mdf
Fe+aO4FmuL0fMYb7OM+LpyLKwgqn6LNddVwadW78E6MXvFryGscmyeRiQFwx0Utg
TxiMFr2Eup1GxIWQ56Da1AqMvXLYlHmykQT9NONGTwDTi/UJZ0TRbv5TjebU9E5q
1pgMJcOsqJWPGk5H+6fDAqewLk/jqJP1rPw55mBky7WgYAt2kWFcDtQiMhwSO/WR
7c6YVNb5v76TEdGhVomYYpbkNAbo6T6NQwfioY9cKpZfTApt4geiOnuuV455t6YO
EKv/jYF8p1nG8PMYgdOaON8WTymOlE3/iN0rIM0T6mvKd+LVwAbKveXvJVwdfRO8
1kdnGCkAjoT+JSG6N8S9vaLUXTeVOIgWfKVHF6/etkePJ4O3Ja2A84T9AoGc85hm
TsGjx7FViBw38NxC9aBC6ZsNp49xpUaxyPir6jFZz9V+fxZg/pgce9mH7T+MQmIl
aDnrSn+vY8PlMuAMYz+RTwLVCAb7YzE2GQQlzYR1UNQn3MblSmDCoJONeNG78AkM
vG1QTH13Qb7ZmDeROhxhq+gHhaEEjeKNkN9A2eZHHsnScMs0SuAdQw3niZ753kez
aDOUQRhEw/lcUtYkdHsnGAbT5MQhgtPJT3+AgS4zzxp+230jVxlyqyPIiu8wRmDE
GuZTL5Z3uHKWD/by8V8NxKvWdwgIt3Za02pkWzDUOmp6vLXroA3mcXKOtRHrPfL9
F/kJdG8oEG6oX/lvLs0E7OLxQD3fcbOrd9C9NCuBi/lZNs/NZYSKxaRapnYKlx8X
SVxFwq+mWQZWH+QDowtQJWbn4VHsKKcQBkxN7Z8OUuGTZxQ3BJzZxoOR440JVqZ8
28GVm5Ktk74Gib8YvgVC2jdvjQTPoeJeoHK2Z3Ckjc1b+E7wH8JFbAZKfigtakcc
12G6Yj2kfZhPlUhlrFTh3I81/Gn77uJiEKHBZsgCZaTozl6n59IdX1q9J/AU7XJE
NOQfSAnpKEFMoI1PgciFmrRqJzF/ZU2LIwFUkTokDNDhlEaQsHefF5PfG+cSHrIp
aogZkOFAlED7tuEclRL9c5aguNl+DEDEoFAyPcYvYkLgpLb3njGu9oFH6o4ajOb+
yvRFi1Ua+U6FGU+erLmRNorFFrPasu5JpKqzT3cuDcvFEzYxDS9TTr1KdKQy4+Kh
WIohNOUvuZmU7LS0itV15fggBVV4sY0nNw4uvun45/1/uFNJd9FvqlmEeW0nnkn8
0/bhCq2wX6V3NZK+vxgfQ5eVU3L/+285psqMhLDvSK+C1rlCqrllQsAouEvv/b/s
t3hkoc1o2yLdKYUhH9hThSwBNjMh23BdpzdzGFD0mNd8sbs80ljaIMhaTl0b68V6
92i8LxjniiIV2pcJSdq3O24GE4B7rfIjTZ5H/I+owozmwPlioslHjcnIfyk9YqE4
ceEVaMuoh9T6fQj842CVLBjoH2YYWiv+Moi3WO05VvzJAEl7i3m1nnG3TdRnkcm6
JnRoxOVgJ8n6fLV5oVBxSEHogSc16iojvcDg1cPquQF8UU8a37MhZke6wNdZG0pc
c2YTCn3WDQAL8sPMeTxyKQ+SMuHBv07d4LZWTePnyOh+MQcfjyATfzRbUJTIGfnV
FWTZX2r599l7RxIW8fJPTVSryjq4EpiUCzdET1l+2JWPtjaWGVOTNePbCWyq0YkW
0RoKorBWPV+zSaS0MPYTYMGdR6VyIiGevLAxjPW06hqg2BsKturNP+IZOfA/36W8
ZMKsb14sjjEXqYBEg2ynLNgyBMp/KbzYiCqzn9wdJB3WEIH2BTM+Lfg944W5qqnM
PDzye/fOgxZSo9Pl+j/jkxIUDcPuHKzwyc0v0kUFG0ThiwFq5D+7YlF1myWzcGTg
5mjPEIOjtyzQiktao19CmlJsKFr6EXb7ch1PxQ1t6jR5aGi4ou7vSFQMXfiji2kM
p+2dvCYBSjnEAVJOp+8q2a9VuAsXOtlqNhxC+UdFtUfGhMIsosMOQHhnb/WC4xZM
tPRMXyhJmGlhBVWdV6F3IJN7HRiDxcwi8BWVR0vHaYjbMTwQFu4jvbKAH5epsSYO
zqq2fv3mDm1fTQ9/L7y2KX77Z8pv4d2EYAg1mnIx7+Ac0HxNS4wU8UQarQ1YDQlr
aGnHjejuXj+3I57X72B2dlc+0P8qIXTObIKnhlaZs6gqflJXZfC7NHRg6s1Qq9h3
iWn7XvBoDfH8R/X+ggAYACSDpMScuz4YjU/Y5f9bih0CwFZV1K1Uwymr5QFP4A7x
jjUxlQ2jvz++xg4ISVzd8U9S1bGrEjq57yxe0dHAMHDNjfyQkVjQcteN1vktHvs8
uJVvSm5os1jBd+G3AAuCihQ/m9dJkfK3GHIIMjFT294AbJEr844xr+PVedUOLu8V
DE3ugBvApHTcsenb3QycgvRr63N1fG97j7BH/FZv4270e//tSeArm8C5V9yFKKab
rlwafVmUMaRmGusEh501vMOcWD6fixGiwJOg2yGNo18slTwiiDk8e66FyQC6+Ukt
obZ6hdmUlfKiJqnikkC6yox5vhi83fylBY5hv+1jnTByAjYisk4inIvy/U12/ic1
7D/UjMcxr5YF2N8iWufsx4/3gMopRHLgFR3Cjvv8N8/EUlFFFW0NJwZNpkl7WDGV
9ARPg6+J5fQtGGbnHRkdyQZg7RpqF0RvLCRn1SIFF0CwBavWZuEPH7C+1HWzQbs3
sxPWDdb4u6snU5+WwGWl27QB+3c8pvq+fITSGGFeJSpuj/EJdo4NO1uZooouwmDe
rWiVrktJPqKpkxEBgG8sdsRwIgGW0nFLAvQKv9/BOoMVrPD8fVR5UbgvlbjCoP68
wT2oFiNeVwtj8E5Ig/YYbFPi//Id0lNSeXL+TBcPHqNIHdtWKNbcv2s/80qElYKO
aYkHsUjyPbLoUl7GDZaaJsROqgLi1CbxDUFAGIdg0N3Y2PUKuTeoV2+kUphKaKvY
e3XY1ugNcguvnVD3P0jAPtIH7aPBkNMKjK7AsR0POUisAGBCdz/as9h1wW7V4E3k
L517X9lOHc9GF59e72/1LnWaa63gsRYvXTNtO5OrGm50UbGZycKSXmR9F6675iz9
DkSSpKbLL9c1ee8fCD/c60mnmuZSz/6lrmi6ooMZdHro40U/8McPIIuSu9GYRscG
+haFLIquusVZ41ufa0Q/RcutELDtY1pPYCt9SPpcrZfQpbGd8ZG/bGeWhY4sGW5C
7Y12gbTs24huo7oZfB72wubuHzJe4ExThZ5Vohu3sevqMUFX5V2mQ45OunONstZm
jL23HM5FlyVyxzQRaVgQQpwpIJDjpOy7fDVUG2Lq8uTXBtgLH0tAYtQgvrVwiRPR
5XMMDdiYV1l9OpQtNNXLL+HH9pwb5Jmw8YV0nq8f5+SMTVbfnQuk0v/fDKhQqxCa
mqFrOL4w+ci36Hul/NQb9TuXt4BIJ43QThRCiNB3DBjOKnldOTlwj7lCIpgWxw17
LLV98choNsUn+ALjMPlz0094G0a3MIGPQEcxGZPWZBmyI5H+HHsuM2ICgCg8s7uc
ZwYpOrt6oiPgHq9dkXEptJhE0dSsP1jyEGPqlVLSXhCXf1/dlu0iVjrXSWlZm83E
a/wN6uMeodQpXV5BMFHnjp9hjZ2hEGWK5rpGntyfkg4zOPzGi+4VldQWl+cdIRck
JPVU/0b0YV+v1zJSW1Je+9FJvFPqcVABT9yuwDO50C5xTi+jd1yfNPYxz5TcrXfa
dQDRu8YA2lt68IGpMvtqLBDDFUXwnY+mKb4cpib2QRZ4mv9tDf8QlT7kdf78D08D
Nn+qRdE0+0RQPt0sqdF0BcxI9mZohdTSEEK1vwMlCOQAPu+cqGlGLuCRjmRJtj18
sl2sfzffA4p7aq0VQ/ngjMsr3Dme+SmspXF/rN1nj4FbXR6cc3nAmh8SRaSv8nJE
rQ/wyjEIAQdmD4uIk7K+JjQgETUGLPPOoOcmuea+4ARcX9zifmetoUQGrMtXbZ9l
MrBLRWEqp5dGhpSnDPiklxmfwcyfKvGgvslM3lEjH2AzzRJO59L7LDR6gSSEr1XV
8ISUn8/s5PiDJ3CHXrV6545W4Fvs4lA2BmQr5H2+qCX72FZbX7WYnTXTrL6O7vpb
xNdAnssWj43AkxVx6RjSLnICo1AAR/jLNQqhl7wOn29z8e/0nqk6nXfBda4um4//
ElmripSzgVk281XRRscjrc/DASNweGYsXXdnKLU4exYAqZctkHf2NSm7mdmvSXtj
CxK6dCDWROe/Rr75WCZcdP912qrRlQV70Qwy7TfRi9EZdXes0Xv/DJS94zpnCqVp
v0erNx6oYn9pZ/mi0QR4UcC4VJaw1UFU6R636KECkGC5VpK1U76bzYQ4bYVYw1R7
yTUWX73D7pVTmzbl06YMvUqKiYvahFwkwuw4bnESH6XAa62GbOcvuDMoLyjl0k2F
IivAsmk+lbm86H0AyjAoNjStdD9eVwyOeCcWUfNU8Ybz7xOAIYis3cGP8MC2+bfn
6UafUXWPvZ3RC0W24LJ23baJPgtEj6qqlQXFiCCsDhkqdnax3VHQJhzaumjWFVZl
kzzpyb/UrUVcg5O6GfJqTutyWOVyH7+iy73/ZJWKZ9mW25oCoyT/lo1hAkRMDDuh
jCrebGTFmt/3ldtnhGwUgyZLEGiYxDLPRlHiroQa+LsGhYnEwJORSO1tvBWiF+P2
wJvPpnMVs82YolrwGt0mucggPESsYGwYWFAA149NmZ+5ry0XAsWxjnYYH3Fw33H/
GqNLjBJGQnrSlzPsU+J8w00SaaTV+3VGJxqM5ZAeTPknyrmEbZvqgs+bvlMv2BkS
gc29BkkhOCOwlpjU98LmjwUamTT4G2KbmgyKlBRh1hgIk4ZIuXH40KdWbYMEKD6G
N+tXrx6FUpKci5rkBjCeDEeFhEKhVRMV3ab2EdFND51rMc2FyhrxWjPAs4hH/N76
bvIm0FUscH8vyInLyeN2udYnupxtNoVECtO1cD1WpfcZ0CUJ/OexTcDFO4HxI0vH
Neu32fVl4SaPhnqX+ZOKbhBQmtvY8+LbxpYQRlP1/Fyjpl5UECC9auRl+0oov5dE
LaG3oLr6xpvAi5GS6bTPXN9Go8D8Wx6brJ7KdMDKJ9qe6kG9kR9diyIgW14ijPi5
ZWpNLXwnS7/QPe/SjeSIYyqkfglqJmTH6xducGYHGe6dMsb5SJ3rgu6prppo3H/c
E60wOvpe9Al73YMiG5++hYxLYe3hxG5qdWyU6R4K9DyaY1tWbGzH4PdIkFETkNv7
YRqS7SzeD00ez+ftKsl4O0ykrtU9sRqpEHumGbz28HyXlPQxjFH2rZr3q9Tv7LxE
l/uyWZUod1c+N+xE67T/oioxYAy3TEZ1xXqvoOOR8Bq6u5lBEi6KaLip5ZbYjFro
9qEZCoYJu0/pOOpfVb2ZvaTi71r4+philCJCXTF11BaFm5M+ob911xmjnC6nvHNh
0lbyttiZXpZMKyu8eLJp0oCl1WMNGfvw01BdhTkoojvNMACMMp4T5NWDqYRdqq2r
veEh8ppjIYTw9yWd+9KXjJW8VgxTZXOzvBwQox08Qvye/BDWYF5ab8HhD27gCDIe
feWTbkbpq8lk7S8J/Wl6OYHE18rnrjQ2/I7D1K3LFqlBzLufgiUY9P/2ijXENVuK
w1jFj1XjnQJW+zfm7VSdqCx6bLK1GX0WtvlcUefrBOPaZVXMS34EosmH7wVAl6th
PSx5ezVkaV656hVUqpw+82X481CszXNsvg+dSVGHrUlxM7Mf75PzMsolc4U764jd
fF92J9i0ywziLymtGgrpU/GG33Es/1oE6CnI+ZHxDQwEqcP9xxgj13nPMHvgaotM
BUVSZ/kuJwYf5jtU+hLVCEPm6tfqgIZU177hnlkAhqtWx7ZevXMlOv2bMqyJRz2r
ANuSKdMqVPaiUvDFhLTe01Sczd7ZyLxqKjA9d6SnypgdbHrNt5u6ZDrY+jFAH+C6
mL9cUqNVwZJlxxbfbHKo5r4fXn0TaMVFf1toPz4nf6aEAI+11nqK5aVJoenAI2/t
J6HdRU4FYyhhGgqzJ1aujNhMCqw2x/ShHa4ZIgJJM12lq5m3JE2V4jXKSXDcbA61
Lm0NSqqMg0Z2s/f+7j9W5nHIxUgd1pvOXE/xX0J6lfZD2VkOv2O+4APcNHavTbqH
RzoUPWbxHQxH16K8tmCmZnX1XbLDUoCmhwTro2vor2u79wPOF3YGjga47T/jcuhM
5ly+QfcZPMKquhdxGMHfCQSGuR1JDa7AMD+lx4/vHOdCju5jVnJU80i2JkmYg+cb
cNvWh/t1K22YjxwIXOVEZF5rZEecAhIErzO4rI25bDdFo7WjUxMDs3ArEjcwHjY7
VsTijdkKa4BqvD10DTB1zxEc2SJ2ercG2KH0sJQrT8oINhJKbKirD8UMG2qGbC35
vWut5dCTjaBIuAlREsdmctX/E0Pu6eSEPplNK5RVb6y8K8QuvXqQssHURPGJbKTQ
4ct1QyOpbYskxieZNDzcC7QTuvqEyYsTx37AMbZ9lL4B1m7jwtNDwXHjLSO+RShe
s4tmkJ0pdadmpZZHvRulvO0X7c09gImU9n9Al/mDEVW16EXOFN5kfDtKJiAUi3Po
Rj4mGLTIrhHxqRM8qndSCGYPPxG2I1WxIW+En3ElmH/mDPqEhL6X8Eh8dhxKxnca
WHk5PbNgOCUP+bA8E7KI8EX8yoBJV/ROb1CzeB3NZxh5cNOPc763pSRvMo4mfD0D
jYxIGrk/4esJ1xqLVmC4wEDFrHd0cr4e6PwOoz1hl6U0yFIIhqmiP+7xni0ksq8B
8NQvZzAUyuPF4oVAz+FLcFD33mMEsLphH7Gbdzlqg9haDfDiut1GBWBu7sdLRA0/
mDICgixj4Ypukn8ujNI0PO289l0XsNNBcMk7YTbLuvb/mvSkpEz5JZ5W9NT7HbeG
GZvTGj0gmE+AP/A5xV2TlP1YSIaRN48mXnbMMzH4yPTrzWAI0YH5skeAhmWoLqIi
x/h4Zsyd7+2Rm5vBmyxfzQA+tmR7o31EUA9zr4iRHp4uUvLOgkL7i9bkAN2bj/aa
f30p5OfC4aExpPRniF0TFQJOY/TytaG64ifvUz21DEGd1Te1/qnMrcpypOAQA0mr
G4sO4hmotacIsqKOSPa+W2QM0e1dkMptw4qv6wu/wzqI6yHQ1uKCrxH/me6nlrRU
4Cesc52UMU9sclIeluJ9bFLUaxY8ktHmFHbAsWasQzEiFenUncbJUyj1HMpX5Aww
KYKns/xGcwlvnptYTbVGGEyUiQAM1UNh3z0MVQvll01OrzvTlCiCY7zg0omzjFzJ
hKRo+h7Pw3e3QURZAPuH4DHLz0YNkdSemyfOA5JyC9IMtIC+1jbOSySj4qFvCsBh
4FqmJ0Gc4iE5HKE1lSnvg9hJOCTA1ZKryPlf+aOlrQZAS1aoBu4D/8JCl/HlVMFn
YKms2g5rHTY9S3gR5nPAioD793WxWUHs3jpi6WjoWeSb0LFxbidvnWZeF6MKvhT3
rYSrL3ZnuxyNfaV2iXvzc3f+c2yhpTamNedP+1ebVavZxzNlrINSb3LjR9HlCsnw
C8qn1Rr5ddDLBf9kJBO8MP08gRkoSxAUzNNMQCGfwIltY0FX6Ef1BagbMd6fqTpy
tOV/gSWW0tvbCxxRE7oNgOZDH4wkH+jgrGMW67iHKDdRrTOhEou4eADy+tzX4sQ7
8YK4YDdDaduqEAPX5f2Zb6ILUg8qc/2aVYG6RmqBeNYirUrrigr+pk/vsofjaa3o
lHGq3O2zoZ44/f7pZZ0x9ROA3kEe87+mzkaXZ3xzO2YF8TzPSQRnlSddsampyU72
UrfipHqJ30UN9+dqGSFYeY8VDKzyeI3QSNoI8smt9ERdTpfxv5aVUrUYPwVR8rAU
UhPHTyw2KtjQ2uAHMhQLs7gCLkF/6BwnRqmRiPiy0K7xGGnbJfQABnhx6rGIdmLe
xO76pChqDiLlbAp6+C84K94Zx/tfFkk4Xt6Mwive0A+jeP1sQHS3XQ+Fss9Nn+8N
QHqa0x+ffFTeXKSWLI96hRVPfpL81A5DuYK0TBFenhac3HNVcgydoX+OCpPiPkvA
okwRcZXHmVfDCtK+JJ9L/Z+/IyBifAwBZ1vHKMzGFL5BL2u6/6yO3cCjIlXNwB+L
PBkcDQVcyljuRGRHuTQ3HeY0i3wW5qVJspfU1crG6cHi/Z+XKhdikIJh50tFUjwP
Ng5toISU6GOOoaW7jS1mSNuLKFSeGs4VFOB9c54YzExJPprSacnsdzNU09Zo2vXQ
TtrxvpPpga5fYkl6D9VupsHz0Oos5hEqZ8C9HO62S2UQnxwdPHd5C0LdXpWdtdI0
T2NSdyoYyRkffIpfe6xGuJ2pVAlesprtz2ur+09KkROTYFu05GPHFtcImkwqIPub
sY6Ifatxw75017UtHFideK/sX/pFoASz3/JSF744CCKbX69d3PuJ3VHa6nvoTCo9
X2YH6L0tSQiQY/0wI7wNFRldZiyAYfcJcRsbsZthdpShTYuJopYLGDicifEHVAqQ
wqaCHYMaDxFa9iuqZUYPpCwTpf5+VRXPnPywYq55AqSZFndpZ/KPXjKUREvzEANu
NHGMb+vuzeivoh5AV5736/YHjVFZ4RmVxBiKGVaG5h9tRtst7/oDH60hCcT6BGmt
7eEQzgQACQRcJL1YLRjJQ8BJ6CIXZS319ZpmfuV2XpR11sTUEfe0s8P38ZXkuAvV
8y6JHqdilJvtcqBwMyJOwtjx8a48l4/IiqxV+7384lJ8k6Uj45YCH5+NLVMDkdHC
WC4fCLAmQIjCirDhBY/RmugTslA8fz7//HX+bRMjPwu+a6GezPTRim+gpCcTEBbu
tqdAq/2G8CFq7juQnvBRtrkg3nYfWlaMTZJSFjgXDAz5a0nO6bJHJjKf1pnMZBeA
pI9pHJE7Upy/Pn3okwml5SizwUExJ/f27SV3yNkWefszoj514tpDSrpvlacdheNS
CXM/Pxqj0sxiafnE5kWhkOVJ0YjLVpdZs/ZR8pP/JavKSepzEKfQahVlkGZK/ROq
fP2lQwB5xY08GOzdDLPlX/zkWy1K6Z+zyQVX0XhTmBE6ob2svVQrgoKdZseNUSrI
lt1BNRzB1GJJf9Zv4KX2U9pQW6vIS42xax3pPkBhQpUPkpmCrvWTRCFJLyIrQlXf
5XjsIiZmfW7PBu+wAmxip2uYcfEsGhCUSa1ZA/em9u/5Ryey8Oo34tJSgjsfMdYE
XKbMZNW18jHpzFSlwauHvUiqp/JcwwCH7yWSv/hAgfJU+MFAaz+aqu2QUqBimtsg
6TlKyIWgFLhy1ZhhfKBqi9SG+8YO9kjKfSi+xSZp0Ozke3kYrqrIOMsKpngH1f6Q
HmhbT3NO67DgrFM9kBEH4sANJqtw4FzlLxiETfncXEyXxhxe47ZqUK2fVnB0l2iH
PCvb/OZMYrQx6TfBW4hEvpyXYpwclrMIh5Jy72eu1eMUPynynOGyixjWqXN/9iif
5CjSLYCyQ0zxmYxeJBQAcM2umY/6Qc9yJa83/PV4ck1OzqGhQwJmOp9xiaVd0r4Y
CfRXXDEkMPdX7Uy5qVmGWBMdHyjgHu9lzAKBFuO0gkLcGH7OLeWi6QnSUCjiC6za
nhuxQlK0BY9il+3QVDqq7LK/u+fMNyiTaRFTfcWNNEUcMYvTfe2XIpFj5qGGSFiH
z95j0Zifg8BGsxIt1WwpXrmNh25F3SMpIsld/5NrRQsPd6BPsb7r0BSYkZ2aPa9+
ICTW08UZP+GZsEqgbALtH3mNNO7E0ulVg/86UEky08WkXrd2gnJbnB6dcYs/5frl
natyIHvo8Wmj/X9XZgTIrif8i/dDyOtzNJ+JjRKdPuWthumx7toWHQ0WDqYm2Khu
etpOoKTiuw3t2fD0j6hv2xbSxwq6TZWbJzGVYMHu4+fbX8Y/u5Z70sqmRX6eRNCN
cJ6qMC9cuBrYEcV8led+d/YwV5nXuW24IXZINcbN8G1fU69mpPVYhmbZc015Fg+2
8wxnni3b7+5oavgO7b1YaWOu37pTNveb8mSWb9rTI4zn9RcW0nrdorDdQldcqU3V
IxCMMBpJ/eVPjpS62ktVC1w6e1fFoqJ7PNkXsMwVE02Q38xITM4BA5GSKnDYHvt9
2ypY+qvRj3yhnqlbFgYM+ZdeRoHAntMfXCJq2ubuxdZMWeRABVk6MK+vqV8bVLi8
F8ppcRuE/GCIRpTTXpGkYHyfqXPYrpD0CS27FPrUWCuysk8Ev5Dtkf9cMBSKfQJS
uzRGbrqMQycONlDBH9hZHe+cATIUL+/DwBfvbnfLk2H8N+zSIsxo5rY2iUyx1K12
qZaroix5rR4EqwyHYkibL4pAOlRE+pn7+cgttfzHPFlBRcucoNOgcrrhgWU8Um9w
CzwDbg/3TQzTruwclce1iDSWMQp1am9xttR03qbFa9p+ymGkSnUpSWD25qbCRm1A
B4krDK7s/S6H6LLjmFStQ4sycaMYs8QuEwYHCYhwGO6DkH9rG6jMuQGQ3y2658wF
B3FNwSO92nBq+w1GoN1ff5NcV8ZB5mZEnZ6n1lVaJAziXSMd30p3Wq9JTJsEkg1k
QAXcE9+2dLxdIQCssvjvWrBaF7w/5XWtX0BDQ8SElUeBiVC2B/z7wRuX9flWlAuT
u0uBsBgU+7vwWxOb/4vHG7E1MfRI3BBbnNGZNWUrIiFWz0lLAPvcVUBoRlOFYuzu
KtxSbEM080oiC6i9a7ZBi1gOwU9fOYXGhksGRLuX8FGSTpp9lKJvypwBVg1DGpsA
Ryxo7gKKBygFItjQ6Z98ZFHqsPDj7JgG7RLsDehTWZsd6NpsPIOc/rlar/PPIj8D
RDHBdrIGbtY2Ff8nSKo6ynGk4joDBTalgu6KFKawhgMdABlMujP0vFAOa5Sowji6
TWu7pdni1DSJ0lBkYCG3Ny0RkFfQurF6oU32PYQKgFCdE8EBXX4TJxnlPNsCg1vt
Gexxu+50oCrpwK1XeqLWOjLiBV9UWPmeE0/LfwiQd0I/nS7Fwen3JLEHe4eeSS4O
LhyrgAM4AsLlvfiM0CeJr+7jGdhbdqmW+Jxqs/eZWSxl3qcr8T/wnJ1N2Lmyw7+N
aRgxf+Ifvcc7L9H1beoJs2qG0KBICo6HUBX6H6f/x414FCjGDzLn0rMoUPP3SJ4Y
kSYv3+UIu0QeTI3tzbZoanXVYuL6huz8YYw7TR15O7qMy42HEYGkn2p5t65mYdyS
BRbXx4+pEnLRCErZX0lV801UqOuen44r9m6m0p2nyjjjJgLZzKPbIflkXiwWEuMK
mJeTS5mexGXU2zV0EuQtYRBzSaJCOxSGXb1qsiz9ZQTcmHIbAC/EOSsPfHtIxSgO
5RW9autTz3tHpysQZaWnUCTrAhhmZ0sxMNB7emwOcrsF5+X0UcJ8UHtqvPZEwGD8
KGuH+tCbJPMFFoNbG+mHEM/NgMXb9SytttPcP0RsW5CIogRt449tRh3i809NAzsI
qAAmcZ++J9Ekp7ERlJa9JCrb9B3T8wK0mkSTLZUT85ivqQr2BR+vnzJLUFo2ILZ9
hJlVrdpQijqFnWOj9uZcQFJ/cAQMn8RPH1KSvyoKL3OBzP/ecDDTUFq4jX81/sYK
B31+3qsdIs0aCES3NU+AdHgC2s2GU7xef3PUBAc7kECWNqEF1VLE1jG0wawwPN1I
m5UwhcZxG8piCVwX6rAT6yHRpL65YiBrb+Aud13NCIheEzzElSRmbZAB3/MZUTX7
UpmM3p+piwNC4Ede8hnppThQ6kpUYnE0VaZnwVWCHe/zzs5sRNfLAnMFj8QBF22i
I3npj3H6zfTQqBIyASyDMoUW9esXWnlp6kM4GqQFkdwRfGjLH/7yxq6UnMVO5iWd
b9mGRg1veC8cLRbWSCAthkejF+VRquyjLXNEaU5FrpSi6cGNblxbIMAgPRMdbg9i
yaK4xWXwS/7KD+QdbMVdZmPOzVaCAb1+/Z0L+8ms0ifkqWsHHMs2xECiYqYIU6sb
aDIXwNOKXeSJza68l5nEjW/lNF82TKOw03cbn/WjnVr24iEDJCXAxm2+Yg6hm3Yw
lrZFZtbVxok5oQOYaPx4SMbD6bKJCusV1BymNtN+/nefd8hB3V+bNz+Yj5j9vDSx
Nxae9tRznKyddG+taLmXFVGR1YogygslZufPEPFUONLm/J6OxF5PBavlLAhIgXK5
GNg65kvgZV0r3WCBdIsKcTPPyNL5mUnJ8L+zF+dvuho37BNnLTvVD2xHBwRmNIEu
zOwShkobxsgszIYsySaxhSkVCJiWZDKM7NJEgNJFjDkloEB9oqMSqt4BASUBOn/Y
+bNjA4oaPmKRa66bqCjONlBZCFLGsjqraa/k/41Sc3qE41+fzcNNMT9pxfW3K7LG
c8ew/sCvYgmBoaZHQIuFQr8ozMW/M106GReoXCBRzsC/n6TNxvt2xQLrvQfuM7FN
2dVjA1st5k8fp+gIlr0aSXin0UmIqbsaDQyaVPtyh4D73KqszahhWZ2t1l0bEYLz
QZX5itBf8qQ7+ZjmnP5MnyWmr5O+22/ld+w42Jy1zQdXaItZAAuA4GFRN4tHnh56
LVuq1Kgk6Q6Cy6t0pmncwPuwOA0ToWiAgjf/b30eCyNXqJmc+is3MlFwGdEhpkzm
nZMjqE40PjpvnD/HGNvBcuMEGtSwecfz1zWZ8FRaZiivNkAywR2mss29gNAhVpaN
ZabrDsitl8sAlDUEhT+P0S17xuLqgfva5s/OKbmhSUgbsVVjAwTPmAoZ6YfiDIpa
9taDjpQAcdYxrtsaeHYIaHLAW2rOaK+uHkPOXuyVeBnR2FnXPg/UwTqtVxAra8wY
35lQaxau+6h7gAKGwuWBev7HYotH31DxaCxyMxHLJH0Zwr2e2ZHVqw8u4sBEAvCP
+hip4ET/KPpVLd6blI6yfDjKx53Ij5xitMNDeUecee90QqzUy8KBcsYngJJWI2Tm
/ImKuUyG9biG2m8Rb9jQd6vQNg5Pk8LRxzE9RudSkAVNZp0RDacgdhjWrippdCkx
5NSFinM/Rs8N+4aDCnOV4m6SXJzjihdauOwXIZTw87hLUpEJ+Z8ZuiAy2QpblyZt
btrQZC3K0NCrJNmjzLJIiSzGnbG5soL3gqG73Tqos5Ig4fyaq4/SS81DVZ5E9kkX
cHKrFX1NN821dxPCkBztiFfeRhBNFzNVqozXx9ynhGVQHCJrdpXz+wcyb2hRknF5
wRSTqfq+FyOx7ftDaRJnrfp9ccv1o3Dsslh4hNDwpwZkAGzWQ4p1enoU3I7WhXUU
j5H26TXb1Y6qnHhEblRlkVTZoUGWadzC++ZtcZ1APJEf2+sr3ucfC0rfH55kL0Qb
oV8p2sHJ0RQMIyGJOn40rSVGVPvoUY/UzYJVgjCanEAUo0CMXKmC2G2qHf7i/47D
W8q35gsSEbm0QQqcty5/ssbVyC5D2pM4rEwrhE/GUHX22oD/y0x0Z/k4pyAbIFbr
5+saL2YLCy8jnN+bzNpRQqdtNShqJ25slaAuqdlKGDLJax59wRY7KtKb849va3il
JPi1dgnxdJgKoDpXdyVIU8Jt7ee2B74n4OJWFJCJqO3v8EHDiytDdd0aN69WPZ5N
YbX5uUfOqH3vDr8WEjD63FBtFBqvTprjW7ZYjakBG8V8RTa/Q9KMMOe0fR5Sxij+
McDmxtzu/tuaBp0c3Dt6qGHeehIz+g/urjSmRmT2AiOdmEh9hXILIkzubrQmbAt1
VkIQQWkBvqRI7WoQqvDN/UF6BHBpZw3dnJYsoryFUa0glz2Ty21fTH4wwPYQ3l4L
HGqZcbzJjS4kVOxFWGHm6BuBjmbe03NudKCMyiBAYdjuhpWdHzoOM0k0mM3hApya
aBtFVVb3iU2/LtFK1kjftvzDM3EwZRU0TCdDcZzFh5KyXILxhAK2gMX1+p/0SLBy
8q++pKWot3uS9hq+DhEAIsOsz3SW2i3BqhMReCimqwlsVR308Osi0weCtkQ4gPdU
9LiTDPtJ3pRxNlxYRIsr8ZL9IuUuHV8W8QoIleHjxOWut9oymShjdc9Y1eY5a3ny
fEkgUNlvrGHevXb3tpP/oSR/1juBnGa/Jt26UaBMJPglUlSGt7510Jyj/T3KUmx7
bcI+vyJroiLZlTHCw+bzJg2HhPGR4cNhMr7CIZvstqdBzmnERvC/QCv7gzFWiRV1
slnpq7mSjWL/7Pb8V/Fwj0YOmuGnhPkcI3kW6jr3GWHKIoS5D+ZaYS1+QJPRsoTA
en/KJmvQM+CzN+LKtFwSiUJudojdJ6EVoNc/6xoWTIolTW3u/3MmusU6EgqCTg2t
q1VUyDEDmLtqnlToQvDSqDpun5pb2GiJXP+AvK8uNvkl7IXn0REoAD+F2XkavLsh
bK896+styu++QM8HFEny+dZXzVh+sOUoR7+NdJliJjcvEunwCze6Azkv18TAp3yH
gEW5UtCsnDVRfjBrwOgiUJpfucAuZiWSXhuAEAPzsnqSvg/fxvP/LMXYRP1lRuRE
rKEwNgKeW2HfEyMSC3nQFeNQH97G+gwzpZ23rT6Na75ZM79Dnx9/0WXRsopNfCz2
5YE/Jgqe4ERL7/XKd9HKdfcbg/cOatMiGhE1RiN8Gu30b5s0XMyPr0/vRQrJeqiJ
vdTLye5YX+F47nZ7tyb99u4Dc90ERG/wUPzkS/IRUf7Nf8K5AnkDTVA9G+3Y03u5
9Iwar1yaQA8xdsbcAO8jb9g2E79nGHeLQ1jt3Ymt6S4nLbN7fuNem9oWWwIsi18N
GwhK5RzTI4d34KpOPvGdrJcXtpwqjaix8pIngEq3YEkNV1lpzT6dc9K9t49X0hHO
BZJZ023+H9IUyLV2fYcHhX0PQOsbHMG0eSLRZpHfjhDbX6ac5/ihEPb3FLGZtXDk
hAGwyBZNaSm4d/xWqRfyhrPJ5ole0d1fCL6zgMwK5TFzsa7DtEMjUOxgw4HUL7+5
PvIKvCEUZKR8DyrWBa/IT8m5+LMehduT4n2cIbTpuAaHqDWdvX9qG2JpwYkO5fm4
FcdrXOLibctXDgEh8GP2tR3S+HGbJMEKLbm0IaVx9ucez3Rveglsonlb2INTj5t9
Ld/cLCLWn3RKlCnrSEWw60D0xfhIqgmWFx+9MXEZLaYcONKDgYqqgMmK0tUVp2U5
WeG/Bx86/PHXsw9/dHYRLVmC3zSPu3Hv2sfyU/gzm6bJ2aL5KyyuNUKxs0e9M4KU
W6Keg3ka9cccWid159fNBOzJnfDRKHpZnJpN07gh4ZvTPbydu6xAOYvEhMJUA3NE
0kpIJfgkJP9Mc6F2RgduZvVJvuf1FpWXXyBXiHh/0ow7E/SJsOQwcc0BNsIcODRN
bdSzqOR2OgehAGxX0Bh3C1SRprkvWegl7R47+z9zMHpmJOgjyTSS3RukgMxCClqG
NQQKliKODv5VUhbMVd9+jvX+FtvXBcDOZ2x2ROCMJWHaexi0WyD9HQZ81QysBCg/
v4xanorYnhrA0aO3QVqxJMS7G9l1DfCtw9KiEsxz5fZEaBFC50GXJa2AZT26vANx
KibvN+fOJ5AkAdzQB2M90XS/6htv5KrqvVGOAXi603TJ7MyYDmSfdQP4PynNAafA
CHkDRDcRK1DGWSfBs/AVc4pmwYtJJ2jh7TCWmA3/9secYBoXHO4cgbJ9bmAtb4m+
Dgvt0BNRU0xLNQ7l5hFml2tbQ74+5Zt8buicuN7EXg8dFUb7eDG8q8MYOFsOl/wA
pMvfWrqv7k27M9ruga9jtbhwU0/CZXIS6eP6ytRqN/4piB2bp4egduS59/kZX+JK
o+G12WKVceZQilUwzWYza2JMdboqRiwIU3c9YyhpLTV++wZEJogj31OhFaCKQMS6
T8Jw0oQk7hholMUzAduucGESnXsumXIv/bksWenNH4PcuQOltM/SZN3NC4E76112
tXLWLPV/xHwj17nNDhipTSCrIhCFqrkJLIprDVSnt/sgITabSVJAXXbmtw5sHms2
5XE4MLOyxcsLvyeBMwjRQQ3l8DfBBQsr/6PP7ehUjCkZzB6GDzWUyEOuqoNwHWla
6w4JxDY6El7bViXjKV9hibhzvtr3lfBfRjgJg0VyhIgXimJug+jAaf1G8i182+Gq
oy5FqdZmp/8j8406wmBRaiWZHl4FTSbtmAT8vVgJYkhI4s0MxbW29vRLJ/RIwZg/
IGGxFOoX9ljgwYwWWgjQ2oYB7tTXcs2CW3EeNKJSCd70NZ6IDvizdvMBNAQ2HQjM
txmLZHE8MN4maqPH6FSrEXJoQNaGqkg0c0w2YciWZe0lybtXHHq3vddIA6Ans+Hu
Fy6bOZwDklM7I9HUCnx9L1f8GuxGGkyOVOfc8rSyh3Zwm4a7IC5lAFcvhvLcupR9
f4ZAJaUTH3vvBaYBiWv3bgBp6/Nv8XtDiuhKhzjVleLASVfN8sKfaSIMAcRKb0ch
BdhM926H1fMceyaIdP4LkDuDAeB4VZpqZFjvUyjiQhUJA92i9M4TbRDiownCZv6i
9VOQIQtVMv1lTpyqZg3jEj+gkLGYyvEOxhRhOZsS06DZYWldlu82mAU+iP0nc1ns
hpAnd9z9NzRHKujw+GVUMbTor1XogPaccPx2RUOFyeexuyXYNo208giB0bnjA/HL
JfO04HS3fUir4sCjp1Rgt8YEOEfp/EH8DG3ThrAvWi/LO/M1+QUEddtpKM7RjEaz
nApL9gblGKQ0qA1a9Sg5jdY3nARvaJItTOSXvPvaKUzb3av8iDKzKMywPvuSjkHW
GDOOGKiHiBswnUYDuj2C5UJX9iOd8SZa9y8T1B6sE+ciw1qXYTi0Zxz2Hx+e3Qca
5WHZJWmBvVCaoJAqlzi50jTQdt9GCgai04Sm6RadadN2pT9UjctBKFHQi/4a09zY
VP42Il0+nBBD/fNo+k+/igxkPHkwzhojmF3+uDsnWkxuMNJ9/WS1sArUCAtrCHGp
xxhdhfq0+om7ifwf/N6AGYiDgnBVfFqVoYeR1d6PwPhYF2kaPImfRIo+53UZ9wVP
sg7H7OJ3wWcr82KW67vX6oRl2xIX3Zy8SuZceyo2Y6HeVmDbbLlci8qNUCapPb56
3Q2Mdr3/018iXJeGOKVXrtrdd5VtKGtvVdGXQmt7rVD8IRPisjh9H2PRpurJOJHC
rrb9Xcf2ghejYWCxwJHe92PbJ1sEvw2JMssNEyyi15IDz6KlRZKt2d/AVHvKNEmp
FoYEolLMGqixGgwiVF9Z88fU3Uvc9GAhdqQDfa3D6W4g8mCDHcpKCG7gxhjPTln2
Rj/YOYff4agUn9qaG6YmYfn1+CAIa2gHaR3xMDWM0dpGz8Dt6+6iB5i8ylqkRj2p
bJDMSa5JKD8DPBJVfAfM01qLc1hObI1H4N0oADNZ0uftaHa/YQGkyRG0xQWlf7UP
bD1eoorXxQdeZQ5q72FCEGRhnvFf+NsmPXLz28Y/hWuL21bI/honLzw3bWUgkYAz
JUJkSjT/0gsU7H2UiT9W+Ul26+Nlnf74xQSY/qAGhhhRPn5W6QXXWATRZvtgi5gr
/7+dO5GZ0rxynJ4zk4oOJfyc3UNy1K5AgLkSmgRzj1v1tegTTJWSUzYvox7AfLf6
CAw9Kuq9VgDgDsEf1Cqe4iIdbxgXnRG28GWmYVmxN+xsLRdLW3caYVLAhKyZcbBo
Xy37my1M8fuSwN88LZw4KCSpEKyz5CpRvVYjZcNVDJBVe0PikDWfSwdsky+UEPzk
J7vd1rYPJz88vTUiUhljixTn/nWtLelwK+OveTuVJFr2WrTuHVbumvQCQDoULNep
PUK2ui1Fxs+cxCBpRx6dz+i3R5yGirgUc2py/Oa7ji99Tx47gIecmXlkahi9LrEC
ldHCHbNanXhLC3RpD0hc4ZuOi0gaVPlVxui9GiuXJyegzdoBH3OyugyzcwPDOPuY
Skarq5V57vh/ZrFP7bOSaLv+L6eKNYmtIAJXHdCNIRRZADBJr4qpjgLh6LvColTb
3/7ek5R47yCQwhrEUYLTbrcK1kjfmWj0YHLEePXFwTfxcJDpogL9nUFOqlHFS1zv
yMWvaJS/8cLryRhzxzAZufxaPcaMNcSlVtRKRKtOvUdcbBsD7J8V40UCwhILkeuk
vWWAmP50boS0LMMThGgPlKVI5icnD6ssOiYBetdIbIfag9yssLdzBbsRqyP2B5H7
MZoASXtrbEkxpq+ufrwgk2iutWO5GwmoH5urM5joY6VYt+HJBtBIlZMJ5NFrz7cq
OGBmcgZ85gwClIquXwZnZSmdkZs1KwGsrIYTF+IaquZzHvdc0JlU7jylxFh6wSsy
hpiOXhSbvbZvuETtJVHlxLq3PaQiPxs9MgGiHwmpdSX5ZMWbdxMag5HEsM95QR85
WO08ZkNPQ64tbwT1NNW91tjarMNcX22ANLcCVxDbAB05ZwwRoAjNgnR5Zx2ncRZJ
/4J7drEpHrZYpBwaXiy712PoPqrI/TZyzzz7LJBgR6tOhuOaWfpkvQMrDVoM2cig
iEocEm1NTIgjEgxgbNPG231sP4s6TJN06CK3Evg+Yvy7Pbkw76jm2OeGyfDtf2zc
x0Ofp5pI52AemSnXUPmynlkby9oDj8nevXlxDLhg53rmrGmhGL+b7pqSTiAgX++g
/rYwGUtmavWNjALh37eFlV/s1jcWBMrQtnZiVafz7EEA0I3AMp04G2lDwhzLZ3LE
0TFlBfjJCo+TAdzS6GxCMm5rEeS2FV9D2RexdvP/emmP+Z19pYzMUISBUR9kRlaC
/MkiVcCpNd/qs3+7l+xg0BGfXebX7fscBphk/h1ZFMX3e3vYy1sny5Li8t+b3Z99
A8/mgZoGhQQXN+JU6uSAR9kL8sb6HdvYZJvJCh4+x9Iv+J5NN8aa1r4DIxcd9yxe
4zsyv8HExnS+eLMDdFxffH3omKYuH5pl4dX5ov7YSMKsora9t2VK+GyjWTdl1DmU
BmB0UnWNY/zF+QD6x+OdE6Y0+DUbicYLD9CiGSM77akfrqxBXt+QjjS5rFFCaRth
Ja3OX921+8zIIx5NtdyxNdq8ivVJ83phOGM9dfgElzgWIm2QaktSvF5FNAe+OpDk
6V0cXDjB7qypENOwEKJbXQLScwakQFYnBSH8axzywuk5Ovjedj0XYpZkaXpvvAUl
hdd2Rv6HXU0DN1PyvctZSNh+fomgcFoa19/GbZk68yukss3C4zWI4ZdBmzzedRz7
UhuEhVoXJS+DkEc/3Mzn0JBmcgj/SEoa/3P7pjAGx2AmOI49tAESjkrpQ3UL0UzY
pawDb3pWYwMRnNUX6U5J7kuU1fhDntvSb2r+ooUR6+q6Cz7hVZVzFD9f2Ksm0ekJ
7OSrBxyGBCIsIsTJUjXsea/6VVVSWj4CfNOc13OTETem8rf5LsX4O5ylDPr3fI4V
A7StsTu0XJ6wkrXOltmwUEp73+5nKdhCqw0dZHT7czjas4hjmBzG0gidBiXY21as
5+6FA5zT4B9NCcPzE/9RXUlBz+TvGLnUrBIC1boFSdnbPayk0NyvXG0P/DMUQ7Lu
3RkQe5Or/5Jd2JVmDirM6VwaGwBJjhfRXHj2zGNL5Jn2oY9vJMaWWAZESpL65W6p
CmdZK1kXy2p0xnkny6whgPDRgtuODUwNSiRYf7dpviqUh7nQbfwl0DeA7Iokvy3e
nXm4tkrA1koSfEvxD4Uqc9/8z0REcoSFpO1AbtDXU6F4Wzqe6F4N7zXT82EzCh1m
7C499Y4xQgE6/I48uiuNowMPshPUwVGWVsQUJY3/Y9Bb6z63aQUmGlISFzfzbfeW
i54bFatHmGaOMXQh0gXjlECcIrbbygl/lk24RLheLf7mMO7eLTTLcUY2/VniK89v
CtHDInLlA2lk6o3onF3Eu22FJcUlpgGgzGFEV63SQhJsJVyOkQWatiuYKdnGQ7vn
cUt4fxDfBqM0zQEE+xB1xGvYM9oYV2GyjrGdbY4A00umLdFyKaZctNF5lWbdFx/P
2Ko8NMOQp8w3e8O9DuiXMfToB3EpUSPhT98s2WMVVO+1pUyl79Qo7KolvefElb8U
kUfjBE1tFARaaUSSTUL8AplJuZPoFVwsmRneYWFmsj2LJRKJ/yFepVpAFGmQPdaw
X19h0T2VJXMImeROB8KfCwgwxrsYItcw3hwDnL4Tvl2OtB2TGsDU7sg0B0ocyvIg
2EtQyZjYQqD3PFY+UMCOuhMnrrG0mvEOUdzbp74QxqvsM7kpISjKR8DTTsbwVRBD
nndyUAen5/FKS5YNzo+GIiTDHjLazeHo49/6zGuWB+WoKypk6Vzs9rYfVMT3/OM9
Y4gwutP3/IjMc6CmGUorDoKCBwj+1BwQznq93C1RWFrLcxna5idqR08+9n+D70e6
+5cmIBtLm4qRVZpH+21XXRViG12q/vjQEa1iyajLNTWisCPP1WKo/wqabgOJ1UHG
6XqiGHBq8Fb09GVcl1PyWJs/QddozVyhoOBF26vM/obk/j3yY+j8IPQy31PRo8ti
imwO75eptjimeLBwwwXm05Niz/b+3VQ/ny4ABa+QiSFpNEZfKvAmbaN1HdMpgEJ0
xw+R6r4fiVfcHXKl4xkopOnuljHkPp947pfmMbKqoHdwr+2/HasThRy0XuoVNiES
l2Ual3GSyk7KYrKdHnwlvZ7enjOmgjPJ9cbvbCdTKbpHoIfktESj6ENOODmlc2AI
0Ks8bjifZSAb9t5Lvo79ZTilUFTVDIdG/N0t1OTz1p4NA5j4KLo0jPryC1/yoA7L
QZZfpCYCnYBJVYklkoDG794RK6XlXfVPVawXtK2ZiXv6e9e2wI+xE66qHqAfGwOc
Zd3Dwoz1e9Iz21zjB7pV/28ISh/LofB+vmSHJtDJi0IZ2iiKQVpb5pkNgkQztvhk
16olHj9P6Rcu449X6gzOp8XnufKFu7nvF6xspffieH5I08hmAvFdS8HTOMtdvm5W
Hac/42OWuQpPeMCgwG6MBFldlUkP/h7kLLfeg1Xac0O8wHlo/MI6R3uSOmE4yq7k
Q/Wk1R9GtUKp4KH0eDEL4DU620cMGIJD4qBJcLgQCoO1u2XZ3gLXxx1w1ERycOnu
cS8mKf0a43eqQgVHEf5YX2p6Edj7kZa6QNopuaMZHQ+5R3U+PU5tojhYpk0CTTWV
CUfK3siWbptnHfi+Lp7psrpPD0GzIwltKA9lIvlGvrAqpv+f8fvrHH3DleJyHCrT
5i3aDGVq2ws+Nx3STNlYkfah/299ifT4WYr2WHK7zU/TEYW5lPsDCgeRaOnACiZI
WSg0b0ORGxx2lAbRuQrduQ96PDLG0pxgs/tzYQ6C4d+71PIzEYhZ71GPS259QkP4
Jrkt1nOyUTV2c4yPqTMP09PbO7VOrsEBpnBq21ZJIm8OrsUhFFPT9CNqAFkSh20A
HQpA8RMwfHiyR+CT6l0tyjyNXgRYX3KdxB4mFm3LkKY3TJx/UWLlnONFQwecc7eh
fjsTy84dTDiI0KoRZEop3d7UAPGE2IVmECwWXRTgw4bc0pH1pi5bm22OQ7MYXAiX
ZjpE6o624aIwEDhmbTpd8ozyy0/hjBAKyZY8jbvjMlHucsJd6aqMNQFvqglPHt58
84YS2ETuSFatHWUAryg0sVQGN+qAgxK9GWL4/ur30PauJ/0zfeJCoF4EvLLDFSHC
z8lpRF7KJIf9pf+WY4bQtlSJp5xEo94GnvZw8jj3Wlx0cVk84qvyi31JHFYMtQbF
gdInUyrfQSzTUhdC4YownAswYfeDSOMjD+SEssoazFlx4cWT7t6UFQ2mPSGX4eII
NcBlbL8dKjintKgfVY3Ofe+JckYY2z78/aCa5XPPIN+43GRA67yYDaGixjI+64zb
N+LufdUkpt8CDgmpyNtLlDs9aML9ztDU4OY4lD8KKRFeLdCkC+XKpanNbsQyHorS
l0Fe/HG42fz6jJ2U9rSvh2QuTSWuoYfK4KSDldUwrA62uHSIb0z62vpo6QB+JLPJ
I06X7YQgOItjj9eaU3jEDrlBYVy/CJzkRmmItvevjEsMaEuZ4Sp24YqW62r3AMJd
0tYdawZsV0/pX9Ksoq2HSrCaphSBgA/8mz12GuQapVpHiwbBmidJDsCQf8xInFz1
F+kIDrJnmnG66g2GNxfWyaCR7/kf7qVysSFANKkE1oGlocY8dwc4ffQopsKMZSNR
MYGoOfZObh5TxRRwKeUl9x9CtPmJNDIrJBkafd8WON3gn5X2uDHNkXJNSQq169fa
IvNWyXEFZeJUEnrFSvhEA7VgWIBk6vKXR7D4iSjaLmkNrImng1mlTWQEPccIvUGX
inSk4nS2SD9TPKJ/naaeTudf6yGfoclen90qiiXzS6svju2IbPyKnrk/biejGFri
k5CAPjS1WwTn2/ng49sqt9AQGtO2mvNHcUvUSrQW8UHynFjEYLX4G3A69Ueu1ILr
iownut69YIOK/p2yFK/elHo6MckE0vmJDb+7bgHloJMdOvsZRTuL8Nwo4D5ttwJp
oIpNsjjLxxNRd/8V83O1Il9eMOi1FsLrJnZGWX+PnkvrVaTRlxqtFGvMRTzlH43k
ZDT8YPng+MW731jFpBlXGama4bhrMU9SnHAbqoekhtuE4tfigB9umOejVK6Wfafr
nR+Mrl8PoMpxaSwjiieRLSselhzNCzntEKW3bRt6LTmFbXbfjacfO4zTwoqY4p1q
yzPpnYpfpQjZy71KlGrlnuQuMHmd6BrkgR3likTHtHX+V9b6IPXYiUD7z0lZVwcG
MecbDPd9XDn/DViKtSUXqHc15X7eVZ0PIUmXYVJlsYnqC+NBY+XmVwGVnno0phlm
s4PRAzuAW3a9FHNjGALoPJujpojTvIcjV9zmJq0juphy3xPnrGxhRaoBjUQdzRuL
awWLzaKvS1mspqNXAMEkPR2sAerQ/ULVo9SQbz7/fhUWitZqXWngaaN4/2g8uPel
C63WGNDsSLaIcwJzn7SnHlygJMlr29DT4AhW2Rui10O8+CKvjCAW79nWQznrwdSX
NWA4iP3NSJzvi8Eo+KyX+OKDbAafeVgWzLYoLkLFyxWBsPVD63+pXgxGcYlXyZJW
3WUHlciirJ1axNEzO2AHmuwbbXdN3pK6U8rJsTYnI/Gt/vv/t3+mMzPQY8QUnIfL
7psJYSBZQYkh+MvUyU9V4mIuoyPLOS3IBicgNGS5Q1FG9C/wa2nC+rJc0qs1GKj5
pGmp9dBSHRGlCeoIH/EYS/ToErK66kVqdty9usx0JFOty39YuO+BKSPdUm6dxWR4
4HZTHc5GwCzoa2gQrlzbvQAF+PBOCmztuyq/8CCxbXFq2qdCTHH+7Qd3QhSOL2vU
N5K52d9eWf0CXq1/viO5zZeR44gr7tNQenPEhBE6rbC9VCNt/EnGs814rsrboPbC
W7zm+dl0KcwOqqpwjgdE98kr0V4bLmP7gw69416tIb7A+IMQc9HytlEQLAn6BrUd
E5tP7p3p5Jm/O4wxOFUyXnCwX26Btf51ydIuCFRJsyOlclu1j1I0JUgTbRrvy2UH
hhINzMA3rtwR+Q0d1Fxk/0PFKnDa2DvkxG4ock/SkDE5vUwzPbsntraoONiHQ2GS
PVLSCkuOVJo93IZWbiTQ67dmFKEBjziV1gAUg1jJSrARj6oN1TTF5FokqdAtjn7u
tCPgmvXm1PSVFoDHyyA6uFC4FjWOGFjrygBLwZPfwikja2aP/OgYjkchu3vviPMp
RV4qCfwXKW3Bzn6ytrOjGbApvUsMYPIFIGpcDjHki09rfzmmioiKgzopbX5x/3pK
+QBK1H+Jp+TFMUapfsfKX7C2OKsZrh6l1DCDQ/T1HddOdpx3Nlp+LdvGApVtBmZe
qI2/sHD6YrY+RQp1CfNqv6DYxJ1HdtPKA87m2OorbYBQ66NLX42ZsVUPW8hevlBP
Oj2eLeWpx9hJ5xEAfy4jfzLgzkIFzBDBZQSLAS/MJxT1uBlgrUXRXIxa3QrtpwD7
WDSWxgtDqwQp5IesMTgnWGJlhPbYR8VV2hGNtgdsAT+0FdYYyzIZ6REgnXRHLWZg
m8Fuj4qR+agy3tJiYvmIJcorqGOk48EmNiNxgE3TrRuPTB6fAwSJgSFHbpJireul
laZ+jgsDKLea0t1pwX7fq3TyJcq2s7suzoa/7psnYXQ4L1gM51Hqz/P5bwk82xYQ
eKYYMwP+vY29wo33jKOv+3KlzIIzBnNT/zBuVfymvJtYI5tR/4nOnS1naKQXOB3p
FyBGI3nnnLJaKV47vWR78vYPpQ4GB0VPaM9llCnyWIGGcLsXcg5anIshDlfv4jtZ
axDrLG4vTV/zbYYT8C4nLf6m1cSUwKu62CE7QUB+F6sQhx4pruUBHkVVf8x1jUIO
eXgZJhJnb50uOdDvWcuhsR8oJwYSEDm16JiBA1Dg1g480vSSKrb094fBUUhQjLTj
rAENZZm7tzXy/esHq/Z9DLotVaGA+Dd0SoikugCG3oHGNiXbVd8hSfxg0Nia9iTO
S9kV9AO0z4makSzs4zNP/Bl1AS/Fh91444KXaaMRdR4XWJ1Tb4PNEAfVHE45lczR
AV3PBPZjkGiE0Dpn5jdinOjUMMlwF07iyVx5CUHvFOCabHrgyuC3SDikiVxt8fo+
yuv+csu/293e9tncDV7oXqqoQXD3e9YfCFUVGyXOy4w25yJS64dYOpltCPAF8rSo
eic35Bcz9jMmcgFHDLA56+tJwJvXpUc1tvMm0L6bBSyUOwKpmqQ+yfbtbc6h3tZZ
8dCptrl1NpLoRtjnKmJOFqgSrEwf0V3h/pY2gQk+9Ra53J4hdpI8ATJXXVB6jcys
wU5MDRI8OYdDmsPVy2me+QWBslhKaE3upht7Voyulobw1u80mKoGwPth5rfvT78k
ckHg2+GDVTxmdhgEn5PWqrjIo5zqgTKmgDqFzmcJjzxetbBbwGu7bQ6JJkZhJRx0
fVJayh/qVNHW4+UfpMqCT8FBNm3ZMOqTjR7epdMwGDlll7OtO2IzmjarUFB0LdWq
ed+kZ80c7pms+oZ9uPIfpgRtJnZYIZCFHX6CsaeNIJf1ExA9dn9fkVD5jXM2ree6
igMmqSGc5Ugs0LB0vkDJ/A8NNUVKNQ2lm7ELZI+WABFM87SnfKLEdjjv+v+LtFeD
/N3WSr+xyLAjdob5C0X2noJGbssBSMPacE0NYZ3xXVWRMLmWpTIJnv4F5VR6ou/i
xDFmgA4G+mbhWktI1pwphd1XbzESDiOsiVxzs3XF/1ZGTHpaCII4DzxzmR2mcTi8
59upoRYFWU60dQ97LY+QHgaQ4WCjVfg5gcdlBTRMtk29sckx0GaqPqsulF7nrFWT
13zpcHJTKdl21JfD5PSxmPLAF8xhwAqKNS/pOBbbiJXIbdMSJPncInmqIQ4wQvzA
abr19xRSoNNoHJ7jLTJiL6iLIUIM8ETcOR8wRDywwQW/yc/fnL2jOL7tuqBBLMxA
D4N1S3X0WPEL/NI8kpGAKzA9tEDBcy5dhbsHB4HjVLoLzji2WUb74KJAjxNLXkkQ
WrPsqQO4JfBa16tpvsI196Rd/y6piDfLRGLh5NdJOFaH+841hq5F5nw/EVsj8dnV
R/pMcsAY8MBb66qwHsVXgjfBF4GHrOge6OJPpa5jLJUAMU3WivgWNvqrPk2HZNlp
WBDeWe/oNwsDfjy9swtd4P6rbueqz2eBxL3oO+pjMLIYsiCkQUwq1Bu8NT+kWSZd
e9JT9R5zq9Ya96fLRs8DaNecoYBWeSsStUpkUIWpdgiQ1oREgtFL45jVuzZjSEkv
QmPwXVxeuAct+HPe7/1DvosYJIgFDilRia5y1AwjTjNhI5lewbdUWcMqxn7N5qXJ
UOCI4B2Em9GLDx/vV9XovsftnxMGoAVfG16f5ky0e48l+L/C1l/ST7pihXJb1jDY
HRMU0xileeObJNIJoIbZ4xUFgNXg50vX8bIuA90XretnvZvQdFFIhp1qhAx3CCW6
59Ng8Umycf5L8bRn7Ksgcq5E1PwLehqUt25mOLzR4WjBsfgn6v6U33x9Y/u7Fk8S
+whx9LmUS5tsoaaZ7XjjHcrDibYyLo5LfpweeOQQ2i2arQ5sisSvpuiwq5HlZ2Yc
AhrXt1ZqnMNDNKVhsonub5QfYrLTZcVDq8gBK1ZtKcfGheGbJ5dFZNhc8N5jMvTj
2/bVc8pGWg1lL/XpAUc+3KNsg+MOOPXOe4UvtJ2mAUYUL01UQlfrQQ7A3JO8+5qx
bUwKvp+9bVognIDLPicsfAgrcG6r42GCcg24sU7vixUr0tJ5YMMo/GZ1uphdo1Fn
IWiHMLykrolKjSBA/cbEV1Xj6WhjDjm7VfOnJJ/rvwXd8sqUzaR3IehQAEu71MMA
POH85SSHUx9QOcoruAFxBpvuqZXJIl1/UiN6SUGTbURNBBbIv07DYmVLf/iJRiXK
/gOAuyUH/mKnKJcFqqSopr91Hrf3cdUSVvv7dkBexfhOQK9jiRLKnnaTEqaRtEJC
/ejUzpBxRJYnEIRSqKJP6OX0h+3pM3UpMSoGRHjyxMHg5DepluCg+QZmKvSNunxw
sdwfsan2BWXoVzAV2KVplsxmMYzzfcAXik53atuH6dXfpM+ERvacX9YBH7BTTrf5
fNBaIbXK6+HGGatRKXvZ5Z0U3/645kkUyZlo43BkG1NEUOvkD0lSd9JsMWHxbBtj
9Az0h8lC175J7wrJuAU+q7FG8ieentfsH5lwWuTPATAhBNXR8Jvp+jYxEJqsqhjr
sC1SG9nhrbtPHyzGRvwenELV3f5z5seIorScaeQqYuM+n8S9yx4zeyGrpCft2Nnf
jwpB3X+fjEhwCp5SEgx18tPJVMhWg4UvDbPmWbiUa+GJI3uC+otvHKwQBV1i6Pax
5JGCacfFmS3cOyHDSRL0hNQP2ueaXS/0oTyTBBzZHbJUPZQqji96VKKOlwZ1Rz1y
GwvzncA/OWfytdaS5Jwxk9ETDch7HmPD0a915obx2QM4U0cmZz8xUsDfQ2WmJSX5
xJ341YqW2smk0LEbCuC8mMIDJ+fXRRcGFYOfWr2uyI6xbSZxv+o9k1dvDh4FD39C
yKkC5qGjXE6TX3Dpds6cZ5A9t1E9BgT2uHTxNbXoU/D86CyiMBCSGO7y/ECv2o+w
z2CcqSeII7z/URfSrWq5fvjozlndBwsk3Xk1mIV10cjXXd4A96dCBbmBV+uyfWs2
WWKs8NmWMST47CwzP6bdJwgIkeiPIGOFfqv2/w9LWRCj3+7MTkAWQLhnGQadLeE5
AJ/jXgmPPfZXQX/0D1ZIa+Vor7Qr0RlnJEBlMLlcQKbJUqxikCbtov8K1AxVDScn
OlS6UcQ5bFoYl4qNY/imdfXtlFga89shqLUtcSJCuafaPRS4F0lS+D+6vNrABzK5
1fXidUkVqccvgg9zX9UGgets+qPMpySrI4QiEVgmpQWm/Mfw8zmtTyFKDTTwEz+k
KTyZVIY7w2ex7IHn/KzGVKaovh3s9GMG1xLwQtwFx9mrF9TuaZy9vW5bWQsDCr/n
DyRRNVYbVIrDalVFDhQierKI97hMtptpWA6zYrpGd5xM8dYr0nRao+COMyrwwLMU
8qDgkSv4ekUCNyHHU5eS3SSUI3luHG6gNregbHOr8U0u3ynbZkvvhnxHXGa2YQup
HYE7qrzwWyg9Mm/rqxbT53icP7WrYqnLuB+noNUIZGVRzh84Iyfi65E5aXFViWhl
FJuj5YWrhzttxycy+af7yO/3OuM1qpvznYc6Tgs9EvhWAzMYfg4mtVFJe9el6LPj
SHo9Xgq20uiWBhLFkWHo5jWMIOIgMDDxa14VQzy35QcDVWg8up9Y2amL+myBnMAB
31js3+0CVLxtVaV8R26Y14E6rwC7hTFUL9aAkM5XhngImDVuvdXORw29yxB420oe
A6yS9WRRlgb+tuy+NLOz7fpKmJseDp4iM+eZ8fVl1Tq0AhbfE+t5Iffk1QaOepIT
/XNm9XbqTSVQpENLLwpDixWJi9bBu3JdfOerNfDmib04FK4wuV0j+rRNrwkMS3sd
tHWK4uiGX8Km8WFty6JY7zk3ApAHrTLNH8PFQT5AzOu3liMtmPxxrqxbe9Z/tNJd
hIBSz80nIH4TeyyVASxXus8FxSLigTks20rMjjwGuRFCrTkzVHrHCYNNaiusEZA0
OLohdeAea2+rV9koHRcKHBQDihCmx6Wi3WtVBe31jRtFLYmqOfM2cI+jZv8zwcZr
oQpBDJpsXkrE8uZPDkHIA7xm/2yUmBgQlynxiyt/cqG59Mzv3ObiBLHImG1jkHJM
9IGRml/OTwnZaZRrVkCwlG/leXAz8pZYB3eqJ91YYIeyTs6NayAHpPQw33dhHRxc
+/eTEkmh0V27tuAQp/Hf7l4xY1B6lFkfzo/2VZ7thMR2LhyVMurVDwVgPcLISYTG
7Q3mBmBmX2VMZhYxy6FcusTUmDnIFvdJveVt2BvLhQWny6+l/GmlZ/MlVLKPXtyo
Fh3WNx4fDJ/FaVpdioQ5OEHk3cTVSsKackkYaQSTj3kMZdSt34BgB6W+hWYbyS88
vJUj9s0bHBj8cWTRJ4xzwQ1HHOGTCGlLur1CiIJzp6v2hJVNmkFyEw0uyXkTBdlD
mmOCbgLEaiwAk+t3TrmTlNzO0a2smdXHLuc2DNLInc8DbtPbIiXKYNRVNP2BX7PV
SrwXyNoTIw5dc2S/T94mz6Zf1c0Y89wBdD9lYZu5U3LYyR+BobsahTs+MHnDCjAq
lLGgyiVt1y0icvOumfKcHug1kJB4KzaDBasi+x4zrPw+IE7d8EMtiGWxq7PhyZ7K
CPDhll8ToAtVizDoIDTG75UbQhF2kCYBGhQ35NupBWLNKFBp81Z8/caFoRGF1pt4
U6b37EIN5t8r33QjKZc14iwCWNaW4/CNe6ONczgcyxlWT2HSdoAlQCPJeYpOaYWh
g/5iQC49r/84HMY1aN1BqTmTsf9ItN2ZBKF+FQPK++n71wjJhOw3LrUycFOC0Tgl
lUuGBAFNp0GZOvXmIKJeZzShUw+1YL2iYX9Dk7KSOtLjj3PfzvTCwKxqJLNjX87h
h5DqP/pluTj2nWzKoz/qFqSV/G3IV3k8C3Snqy8fouYwjWsjcdqRAUcKCA9NvE/w
XPtNRZDUbuZNKcZ3eszQmthMkdxILFtTIJqYrLthYiun8hh3kx8bSrl+yqpUu1lV
Occ70h/HF0CZ5rOIwW6rQxkxkWA8T8tzp/pthajGUeVtnyUf521w3P3Trf0JcLik
VV7GmJ5NMa0A5jhKJzC/z2X2j2Wo89jTZMV6A/boUCL17Ag8hTeyHvjU+0PkXFUK
1em0Xj+LR1bAGgn150UorJ2cA9TQ9Ww6wQAsvNTs4BNyA8QA8DG4oPVhnb70LGnQ
RIILLucyokYGgY9YYwkU/eTwXOtGGi/xq3cSRhD/pPgfvm1WuhRNNTp6uU/qlUM6
wNs4+pFU1UcCc+Z5i2WKW8X0nMjb8JAYWfVvdNLjXwLz8nu55FIolcchSx6uV8aI
9EWImljR4wUlLmXSnwoqdawS9ZrOO4TLsfo7dXfGbY3FCxYjrvnP4DHvKKUHIOka
J0AMEqN6MQ8PGE985lbeNwEwV49qYWdAuxy6LBSAaEpcTq/tAOMH32AVeq3Yq9VJ
t5nMVq/maO7XBqO/r/0wC7Feio78NKzCemPeTZQoTnSD/xduKzMVlnzM96c3F3+1
woEZslZUNvdlca95B2vhoic43Hi67a/Oz2MJORnS/1treFiWfjS4vKIQq467PVmT
rvFYq88PU0KZNzPxznamOo6dPBRPNmicATHn7yi5LTfLcNUXE7zfpQcNr2nkwbiU
ysckViBoOtwkCmwKCxRTGeU4LiHl1evVWzSQDp7bQojQI8jF6IvCB992N5+GqRGa
TbOSqIgr26lNi5jgZ9cz7zehgBbz4unFCWNMTNUZleT6ljEnno3iRzQz2dKHSYVP
qxdG3G1vsuuKK3TaocuiFaEbqoqf8IusB5u6lNENRRqpkFf2NOmTZxRHu5XRPuPK
K5MS+jxNG3D68L/DUQGw9aHnWSO4Otwl8TtbH8emCaDC/E0O3Ykonlu2dgYnLk7o
s3kCnAxEDf+oY/okRPDcXsz32WxqARCEAP1W6Nz46rIULTynwlMcgC5A6QlAmtfA
pEvJQEbnBrTd+Bc+xWZO9c3i3q5nG3utfdneV0Hy1in4KvmbFXlnBsn7fMTnrw+N
QqV3zlItBRYOMy6ntqtYZquFUzfV80RgNHnfFiSpfyLYSIg18Pf6CEbWeymif1se
b2KmoWibF9RSCcskCB4D/o+yIo95qoTdIz7IWvAFry06PrW7cmpf6ZSq0koea3lz
9AFe5TbEJ+xrw9pLWKXfpsE+gQveUxZfHp6b8mk83ApCT95CXErkTPZ5rjMRNjfY
quZ8PNNdYPJBakM0F/70zWq+ymjUfdcoE9aYXmSKEPcToDTZtFuBQuX66GQfMHzP
6Se4Qs7fv93iCP5EJPLqn5HpMczNMbQMbmHj6XDut3F7so9rDWEekCDDmTpjfHo7
4VRWdO5sGzLYVwMHsOqSFr8QZzKDfjeCc1pz4xv14f5gO/uVqyefILA09UQSiny8
PNAIrGei3vArpJzEmo+YsOayAA7vYIoq0xA7hIydtIPaVLe3qxh3ijf0bgY/Dxgm
K3OB+Gz+k4kacWVbRUvBu6zZ8dXP0FTm8TjHnx6Uwa8FjvCunMUbLeaxdVod5yaz
1ZRzi4uMHVILHDl/0R6JVR4nCDK63zTiv7Ey7O+eu8arGFIa9fj+q0y8r32R2Erc
Xv8N7FdTVKrVEmKAtSmpV4AqLTMpIWSkatylT4AulEheoboVlKdemrlu8Hi/Eaup
p8xwF5nTs3wv49CFSL6QDn8URDM+w9S+QNh//wds5s+2LCq4JtPvE8r1TPHhBPdC
WEX7fhfxM5GzEz2pD7J8eqjfsGwa4lfnFasxvd5wN2sKdqY8yyZIvZ47Sfk6FHFY
98ectlGW4kaGz9ldeuWEzR0tHfAyCkJc+boowDValOJEKoi0n5lZmhuftZofIAGJ
aOujvPwjgoDF3w+5YUkY9IzXOZY4bbsBRjDXCRcvFtnKfPiJzF7mAC6SzxkURAmt
E0wCZV3FDLuoTVFL0WrO8X/RRN0kSw/DU/+E49OYPDaxL0a9xQtysVj3ihhgqi4a
Aq1ugaw73rsKztiI5V049h7lCg/JHPL6RhDaFmz0PnJ1sCYDUkkk2W89PiDSPvjP
aygQMdWEVZS+lH3MDvWcf5llzpFEV2fI+UjbmAzp9//6ZJJYVGDZKG9+gf1lb4QG
s7QZWbWdAM+E0ASuNdmJ5qvlOhd2FyTBcF2jQBxLjdIqrStFmMrupTJKM7yDwrOW
aI73xLSNGOcbpAGMnQQstiJnqcEozGV20POwNVcFGnIEhB7aqjWYiE6Vz62MXICw
hNCL8xAty/oOcn7Q9izDKgYQ6QaIQV5vaKiQAw7eo4BLYw2Exbz0YuSHQatuHh1x
+OHZjTOpHyMSLFb2wLHdDBzCqmS95FWbfWBLNqxDBuL29diCs1mbaEKwahee2r8m
ZG7azddhdq6gv9SwZlBLar/nMMjB1t2FmQzbPDeUgcthUONRPJ6GIX9hbgfKCam5
Wex+Sw08WRATNiF+SRx2BBjY3BcWULUArzVasfbb3lxHxdzrrhg/SkpBMvJe3/sm
9lhOf44E4gmyJDD+m6+DU265LGf8SadAwNOz7Hq9K2S3nXUVZak8FEM7f7DOiids
XPPO177TL70VGHLiId7RFbolKx6llExG6Y8gIXqDhJWfEtuPNt+f36SwPOl0/I3L
UOockkK+QwS2mJESjbXhwMVntZO0Oe8tVCWJizN5cSoQEfhKU3D3af0nJuoIHhpD
EGTfRqtN9YcmP9GM+iE+bMc0lvz6fPgy6j6KUKnzXhoClre7E/uCBsIMsltn3Q4/
0ykmFZixw+jZHzG5mx4SlxMuZ3xbT14gnuqD3vfE4/I+nv7K5gkCfxcX54gO9YSi
ur2GqV0xA7C0egI2g/zLdYYng/4+zVabJTinWWnIYzcc5qhlnmlA6kCOkXvVnYyC
CifjBoCV2H3EgyU2FRjv6Q1Xnzd66T5KO3VJu/q70PdI9CBKVLlSQ05Mulxkw/Kk
eNaxotdpkbS3b4rox7Jr3FmSRpVfNEi5bwmls+vYaJWtrUcrm5rhZSZsdrtiJkI6
jfA8tn08Cro0N7VAA8Ug66Efw1MRDqAgfTd9s4aujJuqP6V5HNBxVyaBL6a1JBQg
S9p0+4/CHTFY/lHi85c5uzG5UIxV7+Wf3IFFj7PTgP3iY2LFB91jY9UgrjOWzMUR
QdVlPcqkAAHzmdfgaZxUaDMchYp7g0A14H3dMKlRnhpgr5epWhdFWhMOAf6Mpqy/
81ROSle/8X+sYxOTwIYR4Cbqg/kIiuFENcwE06UdwhS8OkgQB7MXwOGgSs6rInhE
PUZHeHmS6Y7lGxeWOEcXB0Ru6WZOnDvWIK5aM16s+ZULAhqAL2i96y3Z1/x7WC1D
YTIqS9Z0UZSvYudBZPlaFkct6sBfqjCm90uBQrnowPmlQG34uKitzZwxiOoQ3fgT
QArjbaq/t64tj0GO3dabC6xafm40Gh02/38RO7OjyVXkKRss31Ncb4I37eFHde38
65fXs5rK7XFFnZYnJI4Z18wGsWyzsmAqdfGfozI13GAa6eWjNZ8bmudBpRbyXA1Z
o39Vac0N5vqDQERCmxlp/5PEM47+iWqoCYx7QsnA0yoKHDj9NuqtlWJK3WnxLjjD
M9/dUMNzbdey30YGLkWwVVaR9a7K0khZUs+RmRXpd32Ee3RciDT7nrwYBbAl+XLb
JIiLBzqTMhoQ9Qwo5iq5WCf6+tpdEHoud38eGUQM/zTeamyZTt911tIuTERBWgiv
2oY04tP3j40YZ83/ECSFQmalLdxqoDPtGtqlMwmwHObzOs3y3SflaqUuknaJOfpi
8EHjSISoQm5kZm68MID4HWJ1HGcp7nKsWZcx+bRSFfQxH5Cwme9ATtwiJEHA2ZCh
f+WJQHfFmrGb3GUNQ63TGz+K0vli4Mm5TWx1EO0fZVJl7KHMfs9v8h2uwP2wgfkS
YyKvC4LuCodMFLJmoOKDPg8reSEZ+cM8WnPwbvLwk9GjG7Y4RiGKMVqNmVN04jGA
cRD05lVog308EmWBga609js8CGbHecuOsAObGth7JEVvuZ4JZh2CJ94btwr6THQc
vbs7/GdJvTNM0OrdudjX/6uocS0IYhDqydOLsjmb2GKdSJXS7HO29Du9z/3qmKm8
j5ptf4LHEsEaEZEAAauwmY9WwRDCcoLl0gwimd6yvxFw5hlehaLvt3MdTov1WuJB
m+/jt0HcM1ajnlnUABeP8gUYCgbNlJqk/4ct/rfRmxaY5t3XsJgSvEkkzJWAXCUV
/poPv+W4kZvygD4v41tx2oT5PSqI26SXjPs1Hn5t8RFDNR5bpS32OSnhsST2fftT
1kNDQh91Oe4kudI20TBqFWrUZkLwCwNnFI6HIbyYXnhh2YbuJp5wRVUR8M52r1uK
X7AX8waB/8jsgVCN1IklXMPJHutZVJmxnxpih/u3ZPWUzeWoSCnkg9X1Nc3TVVH6
LbejSGv7fQjBG65lvpWgUng06Ax9XVznnciag8dFmphRqiHGK+GQLBbSKlXLuYp0
2uE+sHgdJ5bOVcmF0UWgxgEcNHzvOarkOciITUF1a/PDuhoKN6kJ/o2e52A9qEB0
MXixhe85zXDVf3QAFO6CtzBRoTHsDMAnzm8R8TD6lH1OuQTB8qduxfx94mzo9NE9
iUzjKed13f5Zdl5ZKDA81Gm66vL1lvotXqXXUuJ+qYA70OeZb3aOGiYLOtQSQQi3
y3ig5w3kAdVuxavdcI7gdWJvou/6F3eS/6izqC1g7EFmZyTmYIG0OQmY2c+MHFOs
HbQLybWJ1fiNqGmwfjToAH6Lw96wZFfozXvDzuimRhIgqp9E4/8XsijltCXwWwUs
zL5+NX4P5BX71c/3/1qJ0A+vJ1KkfcCfcB/HcW2XT57Ui5z6znSq3VAT9IRSfFA9
72W9VbKLl/oCtNtpY741M4LCGa1IJgyX2UbnfWYqONe1XAasiuF9zxmYQwd635nY
Znssn6u1K2WpNjV4moqqPTxRyxbWTwBFylJbPANVaXLimtjlGqAGw2pmgMnrIElR
utYrdvMaNEggIYhgO/bQSdWzzZ8XrqgaSnRsxMqU1t5CF4agkPKHGL2BbOiXfvEw
tzem30ZybBVd1OUa67Y6yCA6HBJheQhYM6Oryw0tlGVGQaoEz4ApkcBQWHLEsorN
gUhZhc49HfXAsTe9wYdiFHBSe9Xi5p/QuOl25pDJCGewlGsF6gTrzeG3pPoJqlq9
lDIOsShn+lSdVusNV6IIEoZMfJ/K/ytpRAZ+/OaT434Vnj2T00LuEQ8COlRjhUxS
zbsN0KZYX5y/qbjnPz2uMO9+fthENwv4lPq1X7vaunF4NVkv/oo2mSYbCvx8ZHtw
fhfmITq2eHj6z2JwKfTa7zkVUyLB265hC7xHly84p/j1j5br6FTbAAusNYCALVdR
/iskpu0Jd5kgIbiGHTA9D0ZyIjhXiOQV1jowSCurqtxRUeQ5TedCZCqCGtVO+vO9
peQqGIq1OnEIBwP5gDvSJV18kGpcur4CksKSmB1Yr0k8yFC9nMeHifJ7jCXWCfGJ
Xn6nx4IRAB5dY/S9HYWr7wA/upClZgA9uMflclM5H6KkTvGsGbwJPbPENc4jvyPk
Mc5X3MqDLPo3xMFcXZv0l7C6a2tVYaScnLEag+y5258scayAUGHJ/8U5KtyfmgZP
CjzQRm9/XTbt/z5vmnkVD4cMPpu2vsAqecV5U5Jpw1C971zoJ/eZT3rWowJQQF69
9icCXpFcnubsMwyNB8ZlD+ZbZxlJZyc16Fhcszmnb9diWoCD76FaYWXK7bqDFoaC
FrWfKi290au2qExZw2a7l1682Quj2lDi198e/xlxfxaVsN6vLDc0MNZsKA50Wgx6
jsqaHtOt6HteXxjguZ1Du3FaWgVCQ/3n8cFJxL2LDEgSa6fg8XgvzFb8h0j0lbO+
Igz8R+C3dbBWPTfM7hQDLCb98uWNT8gxJghGcmC7hPkDgcl1XaBjtzSE0ucaUkco
YG5gZQ29AREsWZw65RkxE+sF0ooOWwdubrsLBSi51Z4ZTGopNGGceXgyDi7YV2J3
rwV8UbWs09V/Hw9ZhnCHFQDHcVs7tFNgZvVTcgz54ory7DejHKDeeC8Z1JK+PORz
YQuJ/UEReDQp042El0j+ylXgvSK9NRQtDEFWht36RGwpsa8/1SdLNYocaRr5FHMx
65jSgSb3vIbnr2A/DQFU8X05Lpyhf9r36VhlqNYu9QSBKtlZs/ar6A5XTyu+Mu3B
4U5zOE6oGHEMZl4QinFCWs0Otddy69kjYFdL2Wu5gx/c+RelE+igbWhLfTMKVfI8
Qrx1g1/qqIhgNFvjGaQzQb2rkFNr0+r75D/BavOOiSO8Um7mpzkKRmkKjOQYnjnU
Axp+uf606wQ+VRgZZwpNEHXhCRbIXFmMqRM1ghx+UfkDhweG4mgQztI+QuDNL8Cj
y00pudsCVrlXuanxqOeE7+YkaCl9Prxn+6ui6EcA6C3+O/zOwrO6Ieen68uK5dV5
guOS/ye3s0tb01WE0eFNHn7ygPpt0bDPIYw5Zb7Ph9UfG9rvRu0DiI+26v91D7a0
SzDn/CYcNaa1rHTT25QjXzgAlbH8eWtq0+hEJhkBcjHOBQqCeReJc5Bu01/gTunr
7DtCL6RDQcn5NlxsqMFbFFJVuwgobmNjlt3ZyoFzZ8BEBx54jzoHHmqNaKT16+bC
Iiaqp9soRc+BgpabcgjQ6an7x+PQGQ5wPO3cGn30txZzcKd68j/BOowcuXforDs3
HqFvDzEqoyuvl6RRAxTxPPKdgE1b8zI1Vqo11tZOYMtTNJbq6Ga4K/ICSWzrHTJn
djb4hRnEJ5uF+PZBNg2TOydT8IsmrGz4JvUmKwbQvuBvq1mhZDppMBDP3WgPSwtf
dQBs1KvoUWjbZZ8xfHNr+uMN0ytxN4NxjKLC+wU3+SC2UWdg7Yty+Br6S98pYtKY
v1SSDbUKXyVSVwQq/5YN83knFTcitTaHatpXyZOIu9SjNo2xIeXcqEKJZdXtZzp2
2x4eT9Sx4X5k7jT09ehbxnt6K9sSHUfFY0v+L61p88A90XN+U5xJDUFE1x82QM7y
MEUHbLdft0yo8cS/bN1I2KQMVhf/dlehp3soSpXt5qjO3aZWFu4EmtqivRnZ3X+D
k9o1XNw2ST10CXDQ3+Q85jc22U6cjvxUsMZz2Mfxe+17+UexzBSivPHDSPcnHI22
EW/1fzJEvtwiNWFHB/zqkGGhxLBfYhBYo/eELZg0PtIN5O19fqjoMJuIUrgxf7J0
ymzC5NE3VtGoqEEtR7Kq4it36oxWdQBGNouctSrE6iFEcdryswyj9XokzxkKoMQf
ppmCyVMwporktG8KrwKyu11s7GPcbvJtoqtyjzYLBNpsprO04eTu5B1jJ4hplbFp
WiSTnubo15sSoqBLw9m7i+N24RsHFpcdHB3zcJwbhcEMOJWyUky/7d+9PPyhAO4O
TY5eP0WlBKW9K/qWptwCR5/h37QvdI/vaJhwKx85OH3jSLlJBs6jUq+gbPuOVSYu
sKv6qXSGMtAvEfNXAKh3l9nGW64G2CRw3ysIuAnz616P6EUvnYrob6vJkqU/Uezl
rIUmhEavQzULqyFIylir9owB+sSGE+T6iJzA4EDFW6B3NIYp+16Gqk80p6M/Trxt
qMRIdT1qOolWJz41jEbiek4uAv7nrPqlKJlAu3FMLpwfWQuLnB9ICJKYkzCIlAED
Fgj9Crv/NcP137ZWUF5pQY0p7SdH5j6IpAYTaU1J8Io84XlTYZptjz3LqDvDaEwD
KK2b5Ulkz3eROKCcoPncd04Uza9yqT8dbmtdb0wbkRgFpQbnm+bR9CtcA3DNRxi7
xTnDaSqsC2/9xJ4csTniq//ZsmgtnPnIIU9lZDlqGhQ3JF6r5S7DztKLNmVLb/7P
qr4P8AjMy+zmGjFAUScg2+xmscOQy4ibR/X681NKEgcaK4+St2VNmHH4VVfn5XXi
J+V3qCnAgBXuClmRwz/gB0kIl4a3l7F48kUYyE6j/7WyvO9CMUwR1nt7kbKL3wSH
yDE1Ex7PxgS9qv1EgKvU5pYJfP2phbnpRbYwByn6o4tZYAgaGRLzhspkw+VeutHP
cE7aSPeH0vQQpVJTZN4HEC2ienYLjQ8dE3uJUB1lpk8ub8lNFgsA06QpLBGxzB3X
uEIGHdu7pwERRN9Vo9vWMvdP+45NXI1Zlc+b6I98kqBIToM0MuA39Ngp1f0KaG5M
NlVzMwakJDHtmjUXzabUaj4KMKneVldPi9q1MioBghI0i39D+sZmz6fyQkyX7Dvp
njBuYFVD28HDdOEaXgTnmoJspJ+++MT8s06J9p8QuPUF/LHfIaBJbHg7I6as/V6n
8fu9jgMyT634FbDwZmWAH7X8GkatMjYsQcUdYzFds1bsT81+LsSnDQJoIf4JteuV
z1RozCWExZOPNiwiPimDQCLoaR7KtonfKxTNuHXiZxKcxG+h3Wacy2TfhvRe0p2j
9Y4joC+9fusxv2qzT+a+v0Cyr2+DFNXJbJ2X5dDuEgr5HFJXONKK4k7PgFZ++H0n
qHzM/63A7fxEd+hmVhpTm60GsYnc+zpPKqL+T7JVJgSlNIY+RWL46tmvJ9CXZe0I
FO6+NxypNDgamDkN4vyPXmgY2E/CQkLrZjIK8p72MhE3InNmZ9mTuwwn7/9mYHoR
y3HBr+lG1EbHE8lRScU935jhJ8oDYfZ8v+CYhCtZF0PdptTlu36LMxEAqdecppo7
+X5FkNmjtUc9aM0A24EC6LagHfioPKl43lgVKRrfa/8obbGXnz4YqwEJuV2Tcbfs
dIkZ1+/+MesLrwZmB9qib46oaGFS6tzlfx/yXMeYlToIhpIWg+If4FZn8gvjtdVM
6WhH/y6o+RZCL12PgZsN4/tpmnMkQHGLTDEoxCXR/EGTvkDeZ89K7mrqrtyK5F5v
cPh2K6UMvL8lA8BcwYt00MRSZTZLFf6Pb+eV5UBNJCOVB/Kr1utnkq+OQ4Hymi6L
/PvyX1lrX8ATtLruPV17+1bV0ojcsh5DNyrXpYf/XGQBHKFCNRk3Qcnx8YaBTs6o
NnAZyR6laqa4X5B4ylQ77uYmYwANtkV9v7gQZGWKCfFpZ+aeA8Uyf4Z4rlm6uLLf
Z4L3FPsvmyavrNxh4fiqjICPtgoskSyILuY4tnpfXxzbuj1vyNdWxHsAQ0WPTcSx
2TAcy9uY1HecbzbZwYtfk3SbMvZSzHK9zN0dVn5xai8RP5x2ybpircLnuE0PLACK
lniQD8Cw637Y2dWZzkOJ/MX6/ArW3lYHyDvXV1fkB0koKPBa/mKEyRvYhtXOKmvg
4wjiRJKoJ+HFKgP4YsAzZ4UuVuDGZbgegVC13j/s8c8l6SzEr9NmYCPkyQhliTiT
t8L/avFZ5+x0P2R6jXArNsiFlm8Im5IZ7AcessdPfbm5zMww6+wLAkqfbx5NYtey
XtOsjlcNOWHq1aKuYx7ZZUnpmNqkKSo6RtZBcxQ96sGDDeRbGYyZDbrSWZhW+Eg/
770nsHDhQSXjlyyczWyxBqINaIjHF7dV7XmwA3pIFpQQKOlJwpa3fKvOK6r06wF2
YI0rn2pOy1gmd3ibNYq2t7nNjGpqiScE66PEmNseVVRb8KD+di14LmbJfhgjbTHu
2qRNmyQEZyLL/wISAb64cPejbTLrsk7165faVQ8yuefBFIqxc9YkCYbY+blXanJ4
0JPuKT7I1vRRMbdqvC6yg41zATWpL8/qQeymwFUB+UuctI5HJcOuzmUK7e7DzLKW
OJTL+3dLcYcKo5us3S+u8bwUlDQSbPcbPc6iKTOXx2i79dhVGQ3onvkaWteD1sgM
msdE4IqRQW8+d5PVAxq6bpV1CnU5FUrGkcpL2j+Q0kMMfAW2iE5cqUP7kLMH0WXx
00P0PLZoOTCdGqDNUBHwC2yBjdu3YdacCwlJ4klE3CHqL/soKMrFj30/cO93/K2T
lDLstQ3rUVt9FAJ8P/QsSu8EEbMXD69VHFNIxG8LbndG9p9dwxcybqozg+WX8X8l
u4S3VTp7Et2u/oPRHo75/d/MS12XzTDKKoPFYnm/N1W+CEttU21XyrMfCJzU6bZY
6N+9XExgzbaWS4BWEc2K+KyBvJFV1RjbUp975ELIyQsmzLbZJ+Lmu0QW4gVSuihP
XAmHnA9JedKPg1CGRSRhHU6zdpFVULXm1MNvrVK/8x/BWUraHM0qEVT4AbxJjpia
P+0GvCx5tEGgsHC2qoC9gzn3s/LaiU5GbnMickarVsa8isHjJ9qd2/c/vfyus0MX
R1EO2OFJiGVEdPKVnHg9x5AY07nxNXu21JByXua8fSJog05/5Wx43LulwcF60ItJ
QZbJRKxrqjETDdsi1mk16iz/FgAnkHPIvfuzN0IPlpBv9m7K9S3NmjCtIWkOAZol
XuJtKbjxJ52tYk1V8PJc98SYzTK8K2IcwXWQ8Gw0+9c/htT3rseYrBm0cWvDhwQW
HfkNhp8+d+JC62NOpK5wiv7g/WFvxFpYJEy+lc9zq3mZ4GhF2h3KnnkzD1UH+sK9
6VjJXvJ6CnrQkdA+H7Va7J1y0g7rT0DTsNa8NHBPPrmOhkKUhKEC5tfIGOdPb1oE
YXy0NWysSlBk5zJnrx2wvA6D8kHXur8v0xUJb0tEySCFJDJPCxr9v5YUpFkrS5v8
w8AstZkA33Prw0me7cgzdMN/aW3viIpOmthTERCNaieE5ETPXONrK8lU7L5hSCwH
1t6nCciuutd5XEBFquLk8KGyOjNbQHTM4RJELiz6eZplv/oao0Cuhs7C2TyZvTlX
y6AFySLEWwU0rwqPV3jmPqjjeefgXqZMZf/ybX6sFVuUy/93EWgXBh03IRHHwCAo
fplDim8kCa4FaCu+Cb/5FxXHl6dz1E22NFV3a/eeghotRqUaL7OE+eA1NQYzoM5e
4hfDzd78Oy3gGB3r1WtMhIliOHQLvzL7vJ25M1i2rV9FwEb1d5bgyRt6T4m7qi/R
uI5g71S10bI8A54GqCyRISmjPW//TzLXSbMCVfw2emPNsAhBGuoKHno5FyGCpBIE
mffJfChwL0M4INXvS0kQPr6d6G5av9eGncJV8oE+b7dCQi+kNv1rKiqygfsVTzTu
ZTB9qoojg+iTJgc/P65LswHx5gKvRh7vtBHaXHKHAqqFevjl7Cm1lq+IONNQ6Lec
aXz/aP+CqtWf34XyA+f3sLpqdYGRxUD6s04RntNtVPQX8RVFQkhn2j8yo2MocmHR
Zg+PU0erqkfQ4K/TmIe/dGdWNJExghRsJUxjGgbUTtdOZ9upOj7GJJm4fCZojWft
8NcMzhik7iOwnYk9CDCQTrsQb+55C6usV5cB6kzB4Hn1l1PcA845vvtWmCsKp+kX
2zbJpIdUi53ETTzDbnGnKmobn0L7kBGCFTVqnczEIDbtjV/D3cIHBO14TaFyMLv5
6n0e6dBc3udJj7HfcC9kB2q/vxpAHP9mzlUNUdQFX4xwhpgsCBY7VCzFYEZpbtfZ
97XG/i30HimyicU2FbkNg3hIbb5/mflXE0vcgMruSGyHP5PrglYIxwRQlzjUYN97
4QxvgRID9jgIJ9/igs7mya9NFEFp4c4IKKyCXipceTluH/6I66pRMm7OpYi6Zxmh
dh2Cir3tiyGOvm5+sPNLxNTPCZrNrYUzeCJVp/R6B25nl40lE6S9dvxnfHbxl77h
7OLE9DfI71Y2xUY0DsekPDLFAuHFYqdrO0SP3Hz8KzP9cJMM3cLGVKEqu9c85MIx
JyRpt5KbWNvwTd7D1MEMq/dSKwMIyCINN2uIVJFhctPxsoZD5j27cAByd99a2Gl9
dNst3Rub3fC4wBEUC6qpm7ltN4kU4YTiRmIL2JDPgj5WypWpe008IrAv117QfqnY
rKNMpsNB28+xYUT/dKT2epIPzizai794GbsSZdV5lmfxMQ3xEU4vP1cCrBZNPJNm
hQo/jB/fsn0OSzgRsJ2jkf8H/qbSa3EMk23GmjtYlxd2w4tOWgLYDyCbirb4rVDk
THTNSDC44FpH7JLUeFZd5beaSesZ4qDcee0IHsCqDByMXZJWRkrjKIBthyblAUVe
cKM91PXsQd7G/kQowFSxmgP7HnR6eLhXYAMgWraJNIGi1kQ5WE0MJg0eVcPubowd
3rTgMQ20RuxUfmoLJcWsdYprHitTBrROQ7CKx2iut+LvTAO8N3Mb2wQKgc48itPU
Jvq19SVxUSQDEMNVg/WF6nU5TuKzSQGcTWcCj9EbDXQrYE+XF3W4p578fZ1MZSK6
cokJrpGaT/W0aNNrTmwECQAp7jB/oBZmngLgZM0AevCN2m29aC5v+JR/is6YXjCn
kYo+APLwc5UQAV6537+YIiK0lkjaW945SHoWeU6JDzTR1kywujzFyOxg2dG+AinP
7ruOjhqN4V6FXwvD47ghJh00SE+BkTEfcXWq2xfkKbx5jcS1m+mk1wNJBaviptLr
RExbpGGEqQ/ymtK08IEgudalikN67cNvZhx+nvLRtt4jzJYY3oaKEOyWNqTQ0Zh4
x2f5nzpQdzZHbJC+CKLnHoyUnU3SX4ADeF1ezGJca4YQvywsHBmtz3wZ4itfTw64
+O4OhbSRyUkbM8q3M7ZSDAOwuMoSdoh6+DHjHiRg/iCaCjLKo8brrM5ScvyOTMy8
GFiv2/kZI/fZmNk3Ewjmg3Jbes/IPELwl/T25cv3GRVuZ7B6RTyi5E92AakvKod+
KzxUeAuN/AbUSe7lmbKr0t6YKAGTjOEm8kMphdBUOKCiTrwaeGNn5HARu9z9rB5V
8bn+3QIfi+o+emGL3hcByGsB4Z2lYPvEr+1N/PNIS6MWx4gId2D7c/gR2Mm9aSfW
5HikmMMCkVmQzHh5bYLf1LwQlmQBbNGJRRipFThrp4tlNLrb/fTmLSW2fceo1URL
EGvE5Yv6g+gp91lUH9LgWsafYsw9/euUU28MzwSpPLuTj6gANU7d1D5+3UAu/Nkl
MEDhkrCrig32Jo4xZmpuj4HLGvhsYiw+1sR8KnGnloEyuDoIIziE6pdZ8rAbalLJ
T5oXlUy6J/4cLZSe8vpMtg1h8rivX38n2jvfZDoBcoth/C1lRc+tsEvJD703gPnI
EMDO35jbHMPap8KBb0cTHZ6JnKTAJUnF2ivnLLB8g4Md/bOVRxweLhg4dH40dBXR
MLaRD3jSJxV7IX5MGYDTHgVgp6rMh1ydAptcI6TeGkcEx1tgjd1OuT0Nr81o70i3
RUvpT/cGV6draR8eJKy0geE2aj76uwKG8A1kuF3zzfYMHMPCSURv3AwaFqFLeJ9q
17fzFFhk6z/262KFJHrMN6XE4gtFxqvqSilJeFAI0qRuGYNYV/VfiNZRe7IsHth9
cqDsza8g4Bt56MJVE2O9wwqVp2xFjFRvAW3P5J+h/OWxCKDN4FWHXqPjilMGrSAA
YMM8C625KFTk1aEqsjOrm5FyfI+J1yitMLKitOF0DbLFbof+XaXXTafWJpeJez/8
zHbB1Km7NkNJajKPIN2FgMKNBm2joS+CGd5Yxy8UhJsqeDn4U+KUF2h+PLqeLZK0
EkBOdKe367jCNVtwyk8jhH18/pFp54+Ja7scpXVy7+hTehIHNS1m3ZWeaN0337Kl
yvivXeqXN2zddnWsQTS8Rvdo93KO485vDE+xgjlaJPsL4MXdp5GIh+YFIC+L+s42
QT+soXNgSGnnlcXwyFjIB5jWiUyCF32MAwlgpf4hjroJGM7+9bQ8R7uVZ/lgQGiI
ZMq1QPKRMp7IaEEuqscqOmeDK8LGtrHn0iEYcbv4/qguo0YItUtAsZNDB3inVizH
QrrUJF+ZNMBmXOpQnb0LgpjvuDM4V5tGeq6IQ/KLRNtfB5YynqY99wJw1g5hxmFC
E1vmCBP70CP7YuBtbKtxMlIsSa2u+5zZUaaUkZjm+qDVi5z+j3ZaMKZIOPQeo6Rq
eE/ALFcjcX48VDuPDZ94ijBpXwdU8r4SXNDyw29XjmQXP4B7a8uZ1EVTAS0qCqxx
rdZm8YVSp7uj+71yT41+ltg0gCnBCLYq3nFSEVnmio30G546a6iiVikUeH8dKTnE
bloushUt67giAdIVkfrH/2LE1bu4SZcSKRWthpQU3bRFurK9MkfgJjgN8zTGK3/z
y6vwd7xAChqxB2LY5hA3TmxyWgU0ZOHkS+ndtKYYaNTo9g3SbRcwqSWZfS/iNS0g
CSPK6vRY+gMTgrFuxSdfhqk4kSRBhYPSGLJTAyIMPJO0PYu0lGFzEZcHl0J+d9iM
uLNj0UNMfArvB0M8lteXOrVVh2acNyn/J60WW4cPLgkVf5SISTSJTqtKUfPCz4sQ
BDwCJwYovaZsapxf+amIKVfaIQaJS70EfoSLaFFCSMCot5a7ytNB1UyecaPzgMf5
LRTRYeOATePSUyWpNcSw6klnEVOL6SYX1hHBop9lbifR9X4yAgqjDj1qFh+OxLcl
YKreuQ0MjVBdrLZ55snfEaKLjQZHb20dp34GPqBemJFGIo3ZJFn+sPUiJj0ixSK8
gwoVKittTjGjAMizfV+7xTCGGcy5KPD8ztjtxVbAZgMm+O/6kqsdmZllrH25zVh/
c4kR6RbtN1jQ2PFIwoM2FoXMWrCSm5/50ryYsJ2FhKnczNwQadOFjot7WemAbmhG
v6Syz+hqZ4Ov7wmKr/kek8qYPA78XMieUA5nWBk5N0OhGopEiUZTvqStBQuxmw0L
xPnFwHnpriBvzpRY7zY07+nQh66dmykWSvKlZR4uan2IHJuLtGsX49zthX2Dkptl
9tEYOw7xJcsEdxkyk69sSGrkwPgMsIiXlY8SceKNIe7I9eww1fuXAcRDVnuyfYsW
Q+f2m+Qi9JxeX35c/srijGj0n/sKqGz/bM3bfKOZzI6CQ/zXCA0LHR8/lHfPfcOc
hVAjdP/9GPeyVvKbILgiZvkrkpyt9maxymATe50gebKYqyULbjVN1zjEmrLcuMGH
h8ciodjc3AN/f43UVzjAuJ9x9mayav9dno8TQcUZ88L8SuVURf9lKQ0cG2bzHHNF
R6Q2+z7t2BH2BMOW8UvUvdOnbEzLJoqgdBcKpOB92tWMUulY/VEax52XQQsP7jQG
lsnHLVMXbD3D21tcwfH6PvFhdTDcDYOBU/B3Lm+LAFgYeetlDKE/u73il5IHOaoB
PCSm6Hq1UrnVPBxq+ouZvaMg6QSPXNKeCd2WHA+bsIGSkIfYyrW56uHRwsCy70fQ
WzfkwKFqOsR1kr1YlNyK8tt1zgBsSrAq34vBOgc1XjR7yLyUlHHp9jQkV8/NNKAv
juBZyaewGu1ejUpMNKrxamHTW7jr3YZ+vmG2PNMH5vdtNfRKg29zBrLUMm2xoiUK
CR9FI1qEEeP6vL+Fdg0fa93Qz2woHjAISUlFRKzpDD9HP0pXZ/hH8mfSVzqWEaOu
yJNQszYQzHZS+Qonr22B+7Ukmglzw5jLQ9MIDUSEo5P7on8b0ungNBDYc+BS+di0
85nVBeEI/Igz7UavwN23dFnjOn1gk8qOJfo4cb9Hwgo1GwY7baYLw2XwAlXoKw2K
CJYQrcxtux53rWRoUsd1/u1I9MbKDbZ9HZs8AADdFHe3IUwrsHJIe2X/QyjbVg7D
QMvnwDFH9jw5duy7C6IwiIzOtAcpmziMXhUf9zV39ELJbl0S9DnEvM1T2kKlNgm+
8qTue9FNO7HwrUkUPHii3uPAQg0mvB2N1DECn0VhiqcQmWkKJ5ZHnaDGer6CD+Z0
IAVB1ub7ToaOEAqCOPPL6KzC6BlnicP/FDpwP/4qJbhxp7kQL0/zJHw6fuqbbu0l
noehLUzKFTqfpurzpzDgin00BAW6N3ilWjMB6lyoqqzXH1Fw0FyXUs7dKiEgxkjw
J+I9L+f5nVDy4Y8vwb7QdM0ywFCxuvt0vHRB0kGnkgMKC1zH38ukOfmJ0Ceg1o7v
ZtH6LYlehhgcX2C8g0dTKhteVD48vE4Q6URO0piHQFsGKZx/+m7HpuKatM8yK3b1
MNmd03YVbUCCGw5wggFPs/V3L/wkaGudrTuVZe2CMpOVVlkfXIQ4ou7a+kXBhFOW
iuZXLQQDFeAAsHSJG6c/RJrFye3fi9cgo0WpoYp2HGvzVj3uxyeTygx3yIZ6GVvN
EyAmK20/qjBj0NJcqNqUy+pgEfe9oimYZGhODFcZz6oS6LZmFS+l+PkmPrmpfnf4
UHJXsK9LpeKdb7DOF0ygji7wz9/LWYyVdi2yTguKLVYtFkwzpIumKfC1DAlkejJ2
u9BrsmOOyHBavGGV3+eChTbnK2acd0MxbRKzarWX5bHpm8CInfsw7FhjIrrMNdSJ
AjK82SeJMBVhWQ3bZpvzt54wPYs07brUv0VUx1rrKxPAVs0bj0wHdxepzehweBvi
JIsn0v6YvzZQgrT7F/IaRFrt+F5punsQJ5NS951wp2c+EKjysf/jZdF6abzRS5pq
d9wRQkYvCaYtq6ZxfJGmoi+hMNanSTUGEV+eb7HZ2IijKf15HQRhf9fLx8ITCiRt
MxS68QQONFS7L+yLL0sMGixUatmAEsdy9+rN2gKKN2FpE4G6KIWGspz3ERsUQieZ
9/FMn/B09FvbWud2oRYhDeJPP5mS6fqUwRcL/71rUfAxNoJj1GR9yw8PPAWVfK+X
5KURbcoADy+C5PWuAul7Er+LnfTTDWDW+EveGkKT36Lm4MbpA6etYSIwh7QwVcC1
Ba55N1ZeVHkivTieEL1uUrD5rF8XgNvXE6Jdms8tLWKnpvln3U4lw3OLP2ED5Qwc
sbwBZuUAzyB5mBIsEmVGYFNnxCHp3hHZO6MJ1+GUzi5Y0zKjd+htWf3v1ma/Fnfk
GOahqTW9qaHt4MBdUYCXfw0vhxo2E53uuc3G4dfvaxHmBupS49oaG5UlIBbBzjMm
SCsQOa+GQ7NGRkkSGKYnSM2qmHjDa48OMRGZ8gy4yzt69MmmZ2X1Ib/My0solhNR
f0L+zIWf2JpOaeasz4MWwCVbm/uEpk0UiZvzox/4lVpfwuvop9kz3dOO8AqzZDVX
Emk2B3jQVkMYBB4Fss7TWxuUq+gGHcp+sW46SpfeITOvyDn+XUa3cJjOWF261mMa
cUVsUfxLMFf29d9geat2QvHi+tcJNc6eNpgtoa54UC4qsyAxgeK/cMnlOYlPIsjz
7XbxMm/cXP7s8yuUJeYhV2WP/v4fSVeeOAvMp5U/90Mqr88dhIhs7gpAG+Kj3PyX
K+29JjDW1CuGNqW2+uN4Y4jwuVZAgS72+2cS2fX2d3mz8IA/HeELUdI1cUUMfmgP
6N3ytNBjWQaWczY4RJKlTaFYrwBueMhYDJEkDWniXD3QkrfHjp7UoAHqpFvOCEdK
aK4XaceIQRakqomPB9+G2L7mvr/RaXWGhRLP400s+dGE1Thgf53yLsmIExZc67NA
hgvdV0w4QSC0Y2LNPOGy7ijb7n/y3cERcJDW/hwSb3UBaNHVZY2bSN+61fqlEVJE
GknS1+Mk129iurQ9pzQaVlhAFFcjQi0SQn8m6fSIlfFtJMCsjoOhE9gTqbyKdogl
XPW1Lwo1L1AwKp4cXiYUidirKo8OlTEdBIdYtSUQEFwpb+LXyqo1MWu4j5jvDb/k
XkwHP5WihWYvqz8nGTfNCDpUVmR8p0ONAr5Y2M/xYR5voTvxUdy5L81rlq/2sd7X
o+JHYbHw597+XpRO+qETS4eUfh8U9Yvvzp6sobnwmxY7XjYyyDZwpYlX1f8+2Ydk
DSBgQcf6yYt5z65CiRCDCsT+xJx+MH9C39ucCbkWpBRxbZCjC54FwfJHkMdUGKXY
UnHIaFgi2rT+5KYFRACPMjeDNqxOaWgyoavY75kxjwSAB9tJAk8NuzVPVK8sMYz7
6wr775sRwACtqftxK/qYdqm7LpZjypz1zhUDAu32JPpvKqKlgIDYra/1WwieBF2v
Y4lHcP4gwAZNLI/pQE12Z5m3EBWGXOJ0g+EiGzruCz2ZqseWp905HHfRnjdJKSZl
C3Dp7ixcMt3DY1MeHfU26CQOY06/ahGTOm+94vNg5uuDAvNE72N5p35pUh1ZTJIX
nzuSEZNxAsPl3IDuO8+NNzQLUj3tAqSQHL+lhD1Juqbi2RFWaD810p3ZLss7iLgn
tCq/elpiqv28+z/A0GZPWl9pVz1vqmH+lm7LZhZENxIDgpIYUkhthKMO//5Ul7SH
JuFoPwE2wXAc1XIv5o16bPTN4//3Ngi/fqAblGHRwJTNIKkjNntq8wwEGmUh3DNa
rlWDZnWHsyyVsBi6LzraXTDAvzIJP4lcqXXh6Mhov3U3JSmaSa50dVYY+Afcj0aS
gpfM+1BeRN3EhkqfwHinpMt9hgv8hVy4qVdL3hBLJMVe8LmyVO8asa7iQfD/B/KD
Tx6T4TPSUxYNVPL1o9+HU8j41ukPwhgvZtNRgn43wGZxHC9ey5iMVNMeN38fh0zW
sAbK+kZ5ihoFCoaBc+6M3KaMO4TEont7bz1BzazCLMDQe5tdcEESnqCfPuaJIMWS
hnKWjpm/eBinZWLGAae+I2K5PG4sRTXRaCOKov/56EfJQ4V1D5XP4P3fGavp532s
AMYShN6yo21rrXQbqVP3uAuajodPFeEVhe5a0Fqmdv727LHgTCrfYrlBjszuKXoG
eWZzRQ6T7G5771BC2H9fA6Zi16fggNmkI4weA0uZkxlqSOMHHSAcaoyLX8/hLMNe
/516Onb2c12OwrUQLtR1lkCNS4At38JUDZFqeBgUAOKerf1OqGIS+L8SooGyR5r7
6NkvaCErgPzzxwmAR2g7ig8AWCGmSWyZx/1En15heLxkICodJR5izfHpFcN2n72K
27MmoPGoFVaq/DrgPXq1qgR6XWzs9fJy0Y88tXddG7Xtxf74XatOBDHE2HZUTZts
yA3eGVQ9n9HTyPKvLmnIrbj/Bqg5lkXLLgwUf4IJmFnoreFau5EiIGt8rxJqbZPz
rPZ+soFbF3gLZeUWifgkxntd23b2xEWKzCQCU2wHJk4JcFx+x1oR7NV+SYZBhGA7
Qm6Gc691zPve815ct+D+xEdYi5xPoSk7t5saDJ+7qLnmlnIScbYZH5epLPfdKUhw
a2z+B3QgStd4fV4Qo3l0MYbaObP/nQvNU8rqX4uvLro2yLuOSLwmoI981Ll8QpjL
wqBhKVcvnM+594g3HGF6yrsQz3hvZ/JvAm9Cu1Yn9n/hzkGiV/P+1EeDs5UYjf0h
4rx2eGWVoN/X/Blm8ASAdn0Cv4Mtt2lHfHP8Y0uQQNoRQ3L7K5qpbvsz8B2a0UD7
0kmCI+5VmZpxF3bnzhs/9BFhnG6E3vr/IIfQ/tZrP8dfNejSKTG8RhwZzWQPhGp/
h/nYAn4iIHCJGBnfEgdQPrIsCzXoZ3+SNl2AiXrj7biGPSvgUPs8Q6Z3gvAZevef
fHKFPA/eR75m6djS1jkn+JNY5hkqsOsKAdossNLr2o4jDo5l2LBCXFIl1WksgLbh
383iopL+Blzcajbmc2V3blAfwN0AnxovdDXQzDu+naeCtiX6yPgxCeu5Yk9CDjDJ
k2gI/BURatFHFhCFP1eumcG2Qxhc8vuseCC0Fd2acbKUGTsuQvl6hSgdgecoupmG
FTP5St4Cbx6mTKVV/SJEqD26DtBis/bOM0abUCw9MNWz7DMckP/v2RcbWOb4OrOG
C8V0+wegR6uh4BylZJoRdr8FodbLlCfjxyTuBd7e1KkVHjNyAg7QMzTgBrQHFA8s
lX7Kh+6s7M+cZ3BToD21/CuYV+EaDHEG2FOme8Z7R15zYc0HfAUHSeHONqtt1orz
gbJi6a+D+9wQEGIVXYo3yvXJZz272xT8IO2qsLFWciV8eiCAiI3Ezt/hRbuuTi/6
X0qnidBuwvm3bl6ZxctrrVO+LGfmpfhdLkwESAMMH0nAKzx8gQqFRuN4unXX2P9e
ybI7t6wOUXFqqQreLdRu2xL54iYs/G/4RhAi+/0AVq22KF3RIPpLF6ofkz+II/Qj
FOkshndMnNTfNFvqBdzlXZj/+boz0ZZ+D8DnrPMQ2Ii6MvO3q6QaINODT3DraPfV
Q9wghGpW9uBFzFPQHoQZOdAvX/EPw8aPxR95HlS+so9ctYnpnB2qBQbzAbZwxhNH
pUSrby3EAjMgkimJDHtQyg36kqWOfxueHRtc+JcGaod4DVPtiyEvRgtCmtVi6lBk
27JZz9jQXk5txVM512PyXtamalW3hGZydkC8GmtNx3OY+51kE1/k21kFTo24NwYn
XvCGVNSVQOuJQXkDh6NYGbQ+hu0oTiY5jY2ZJsNmZudrxwfrGNpM/Z0oGF2GkCT4
G1lbltPerbkRt6aCxzPA0IIDK/KIQPqCNET4AV9PoOnx8P8KvkBenEn+ESVr04gv
ZNoPlpfN7U22QJWO2h4A/HzFBvGhR/KKS5NEVOkOqtL0u4CIKrbu7I8DYdmaVS0X
xHCUTSZOX2dWoJaUx4vyvRxqx5zbhQUOX8Ucf2ATlF8QKrkuVn/1fWgw4S9qGTis
kABR+QYCaoiCcnbVCvtaXvQWM99hDCfUvtBaFwSKKHbx777DVA1awh2G5W1LX3XF
2s7WkgMSltU4UvhmUXqSeYnFBzXkjdLtg0q9UW57IpXFPJjtU7/+Y5lVwEnF4Ead
lp5YZTVZdqvUZBb28locw5wdetI3ZrOlP05jZjl2ZyMMURKuuq0qYxgLNLmT9KN8
0wajHnabwgEVKaXmd9X433rBK1PnLP+NMEadqJAGSjq7i2gB9pSL75T1f+60HF1x
mg++vj3p0QdIkEQtHFDi6fNW2xSYYNgtdqcKyHeFOMfu+uIxmFiLkBhortL55ffo
2ajjEpf8l1FtqTqa2gpdMk4fjsQdtKLBJGp5cieITIf/87sulXDREziRyoZvIUWA
SpSCEYPbwj+PZl5Lxvss+FbTOgUQbWDTevRVcUHW5brpJQmZlnEMJ5zWtQmkwPU+
8gUDbKRar9oXKRrIpxjb83fggKbayYBfHY1GTf+XN02wEW8UPPT0jMn9ZH5AU99n
q0kWgz1eA36pH7HhWe597sNilsSSgCWJewTx279YIkgieN5LU2AvPEYrrcg6SuYF
Ai1/DzAVr68AsvGE7PMzORYuhFRsXpGcfeSeo0vfY1+ZWM5RXzO8P6GlbkkUlf7K
Y6rrEGomyv42jQCHYw/TclKD5cedFSEd/lA3la6VepaN5ggvePMyOw/PmtnGNGS0
WuJ0DPEnMRU9L4UTP0cDcpNH7q1kNuPsD4GxmTzozg48QhokB/BSQPVMt4TAmFbt
4bSpnsfS1oLj5HhtX/NF+llmmvql4TtbcvmuJ217IuvOVeoKNJZsfPbB0VqVdgdI
hupk1HaR2X/UAnHAimWyG312v5RWvYUrAlMV5ZSSnwfD55wrorw0qX6K1vafkxJF
yV5YkgttbMDM60leBiQLITr9Lz/0d/gQZz3bUf+nRuFH3SZIOAFlRcePMCHZTkf0
P9hm9HMt2I6OuJMX6YDxMmNXJ7J0fKXY+iW8/qDtUVF0mv9izmmooJbsJvKAqK7U
XiCor8XvK657gU7+eyue+JIt3ByyCQq8CfALjy0SXMjULyTtmYTshlmw+5QXBjol
azm/ntZSgt5p9uXgldEIX5ypaBpUTsyytNSTQHGpjB/+H79XtssNYjI2LpCj98XY
X4S7JZ7l+j6R8U87Ma82/ipC+evK9EOrGqkY6bQJFFBDmKgejAJJA+W3S2mM0j5m
59TE+fUTHaCHfeBoBg6OT+p43mYZr3Y/1wobGYXSEJ0DnuFml4lNFV6feP7HD++U
ozufGvClBazqsKcV5t6L6qON50DAlCrrLJzmVX9fxjNhZz1TAa1AJ/RZi1QcYHr/
symFMjJQl4Oqc3DYckrFShI4IDiTuh6OQIz+hl3co6stbTvBreLyPqYANIYLebAJ
SlEd7THCqKcv2w2awvmmf8gurXC/lrjvaZJ8+GQ6eUFHiC9x6pR+m6UDAaMjWVfH
gey4N0n3xZ6zfUIzlOoNs7pl8LrbSi3xF1w3SyuN+IexJCfkWOPV15tqfIplecfa
y4TUPPVyu9pbpWn/gLOlsMW+SCMz4A1AtpsysACfdJMgnEPHdXzUCdFmKM+KduQi
GqDmrCFtFWDFomVfnn3/IxQkf2ZxKh++xp7VLlBrYVQ0lGhbWyy00RgdZfxXIMwa
uOwuZxmYQempLMFnVdBE/BgMT4XADhm/V2wsizUVYQZjduJyL01y4R2uhDjYhXOW
g/sz0VvgFc8vte5tRO8zrVjidNhtfCENihYyFoQIzwsZbRJv/ClQ0bD8R7mglkFq
yNmuRFLThQGiyLlEWo08/iTqS1SqzOPhcW0MLPCsksScSeH9wq1P1TnOmJ1qT54k
K3AlpPRaSE38gjiiDbPzv/ZzZKyGqTjfqSnz3brSSRpzQGpL2nStiZNZcQ5ftrd4
Ei0EeaPAoSnJOJsr2K0J8OJI/XPLGeIrbf2m75VI4IWwxps11EvZNPbIr/Omnant
XYXJqJXrQKxsEZX0hG3KMApQ6YiNSTfWn6Y441/D1JvecLtftQCyifu5pwmumwGk
s5zegeVtF+ByHTqzWCdMEovG9lsMM5kAVA8mdtr08kkE4xpEC2NX+fyhfeyXVueV
YnO95gmotc3ppTQcWT1C+grG5bPHCWouBYpFiSNCIY9mX6Zb4nBO/CcNMKEpu3zd
NmqbvmYR4opKr3oStlTbRTBpxNSe5GSRA+PPECZNjc3sUpFUFfoPRFyoMHAsl1m3
4o18FcFdq/4sCFgLA9ivW9vjfzDd/W4CUqKyoLb5tXGrkGoWA0kndI4hQ5xonMZS
LCh4W1Z8GacwIZwwjz2OtTtCgYnh01rXByw7HdudnUkSBqwpbeiRLgovvExbiZc5
Iu2jkgFF+fRJJH+tOQzTPvzLMcfhhqrj0m/S56xz6bcUUBSgzx9Qgk2Dpj+3/+UT
kGjVZc5MVWC2Aby7sjiKak0OUCKXhEXlRhvynwNqVa4aL0+xU0wa8eiOftRKzRTP
qhMuseBROGpc1qbR3uHarYrEKgnX6Xnv8pPKfuGTzoGj5FgoBNg8/evXvaQstMXS
8pDgbx1Si0Wc1KvoEepemueGVnVfa4Y061f0gwscW0YjdPaOpZreplnYBwZsT7e6
vqxWMZy4ATyCUOINml713N5Th/LxdU/nTiL2/OmVnObr+/X32REoqRWoy5FzD5eM
F4gFiVFc2ZUmLDp0L8SUBsjqhPidRpDpPbRT/DO7HY3858EE/TbREKJqL15Mo6yk
GpILdULXWa3QKnBxw3N6YqUbfC3d56lzFtluz4TptYiv5Yv/ChgqI99yX622qWz9
3Huzwf7aEh2Zeg6y5HkMAYIRYPvy9QQ+MaebIzpcUajr/NaL7CnjUqbqmfcEhJah
Q0N2GXGfLQ6+hOiBioU3GMRBTHzXQKkd2/+ROpSj7Fjy4vu9Exz3ETtXPY5d/YnX
42LgPnrb0Aipjqru3WMFZj3IY+J2an8FUcdJCV99xBys95faxEH6O2KqstI8UZnS
HRxSjr+O5pyMGTxk39kWSD9kZYUK0hZfGO5nAbs9Ifv0OOQUOzy6z6o+luYkkPvZ
BnmPA5EXnMpipvBxQ0OknrH39z5n9EEgpPthwKIPh7xn4/MaUz+oQUaLeEZPmlVX
U/aGCJ+QLJS3L+oQR0DTEE9uJwrlbURWOe0pz5OnhizToX8p0FaUqvEjNpitbRD0
DY0MFnOYeqfbmR1SA+HlKv5huWb+JU0x3UwXLhBH0OsAJ/oo8mkHTLnag9ndkVFU
PAuqi0QI6EAWe7PQVnPAEH8bK951xwlpSj94PctffqZ1iIJtIElDYms3S1CZWRQw
5VpvoxjCIhcBiSnIZfKJB2dzvcYUT0aZF3CUxRd2pL/NXpJEmi6Xnr/K183yvxZS
4ol03pTPTNbjNQGRoqrYp7F1WKXH9T9MBb8xTlfAmwNei+svH1skYiy92teHWUsh
f54+rglxmeefjO9Zga5Zw10hda4Fxfi9aJkfzk0vnITU2YSCut8umE9GFUrYYMb/
i8gf409rQKGzA8prKZad4NjmAlGBsNDd3yjJ25CtX+gE0ye4hc9pIIEoj8yeEcDS
co+SFWu34cacsiI1Yzz/ejZszDlD6p3jP/oEVj5cRpIkAjupQyJRXjXRN42W+XPt
v1hmqkCK40gAla+hzhVJtgRp+JmWEfHx8n6bztDzUaAtgRj9I4kGfL5JehazO6K7
teEOtXgz2VSbIvpRAhfqrjoFJfFhMs0bQ0/AekgiyyUtI87i6lMZpmFU2F4F+ixh
LsQncgUiAw/BGN1xuzM2dU/XlWa0XDFqadoI2r4fHcsdxqaqFo7id5FFr/vmu4Hp
gCreaQv/Nx1Pfk67RgqO5gyIs+4o5JzsDDTb7rHgs7PVD+6pQ6nfdc/kucB4LdFH
Z3Z+PZhkOncnH/5CAFRVo5VsK8U/PfSvZK78YOdONJzQTjpWc+S7HKjOGfcMMrma
Ukx5Awv1kVpi8WrFDDORAjDjGovR/mt5YgZ43G8cOfskwBTbYsFHi+EBuJqTUihn
jOywvxtf6wJoFPnuN1mOZbo/uC48+JvWjmqYhuPB/wtthDRJOLksuVpA+3s1j25I
40f3FYQZffzjIU9cghzoW1xeJO1NJHW3JdbBPvXC2YG1y1h8A7Bs9n+8ob5s8Zmp
4+5itlHZU4Iig3vRceOF20z+p0G9mhNQmImTrE3fntujgGmPc2USa8l9M1LfaxBU
Uil1ndv6U7xLA4ljuk9cwlT+tbvDsphobbXIrEqXRetqInACCO0J1JRMOrfpHOp3
PhsD2TXMqM+G5X3ldshuv4a0mycofocz9P2orhiiGZQnrorSBIVM+iuXYj6gdcQd
3WboafYyQ0cTa6eY9OiHbHa2HSDLhyYLzNz5eEOompXmXev3cAgf9EeVCabov5tt
HZiGEhd4uLQW9P9fSGp6xm0HGltA7v0ysV+Pu5+VKfMn5InarQME+/obxJh8F86b
lSF8H+fjWYpD8YJtO+lGMxrNUtT6LW2m1fOjdrFX9d5OgOGwHH4amSXpS3tPi41D
X3hCv3y3L50jq0bdyerHNQzMXhML+QAnunCBnKVNKZNq0UYeAHNPR+Ow+AB4APn1
z0D6dPttiRsggDzrHkwVEFmUScTLE82MkQmFuGcurBz8/5FaFNG3TN+wCYObieFT
Ssi5kMMYT27/3J6O+mb20GgB2Gh/GfrnOkjezGZ78vrjs8804c8sCWbjITe96EJC
nOdgO1w4vO3HHmOh+RQJrR2HIXyoaqQtZSdY43in11HjPnyktav9Uzq8usYZpHGw
bjVyBT2GGNY6WORIosJyl6dsWtIjCU/HRWltJ489FVm6/Qcfc6zK2zbtRjr8GxhK
1ZepR0vmnXkS2+IOlUDZoRA+z6vy/kntzXCazLmroAZFtB34rc9J/n59Cnmju52E
sTuzBTCsU8qcgQGb033goqRDDP+FPdz0x1oAfg5TcAGXiGH0f44eUuMEJpeFvFKV
JBg4Y2krc7cNm0ST1jP6Ats7mqZA1vAZ2UuUQPtop0OZcGXlfa89vN+xuRaadw2+
EJn7tnidJt8N3Paldwnhf4AX5TUkaUu5QACr/ZFndTXebYm77+aGP3EcpXIUQtmr
123NpbNcR2fTAQ9VPdovSvS6fybN2LeEOyBNOhOwHfej6r1+hnP2HB8Hku32BxEh
D72Ea8P7dQg303LETh0Hm+h9O/g6WfzFrO8/8j0x3Tok4aB2aOJH3sNS962aVoe0
z8zVK3mDkfT7IXBb8e8uX+UQu2ZSIvpCPqmEadW7EgXSx0sS0QTK9L85GLuzFmGf
7WdJ2Zb7F+jypvPKajOovaNDjBfLPWyt+nTSN3uAZOta8cbCxyv+lsEYZ0chxDBT
hTfASNdnrJ5J7ej4vWZHqU/1tHaFPL6R7iLksayLPaNz6g5n4SF+IMHDO3NSsfPR
92GGZhGIchmbH5DCsIc4eO9KOj8nL1RivZlU3JQnvDetWeELgQrahtRgMkLdAYCy
SvdBF+vLVdNWwzqhQhk4x8SjcyDcuR1V5u2YdwxzFrXL5S+1vdCftSY7olREHFq/
YJ+gD7JLEObM+E5qvAfcWriDcRggNHMttH6YeNQ35GqN3KiU0GkedyqvCHXFNfEw
prdZOH8dxkclI3Zlavm6svRTHN0nJZaDBPyyPNR6ZtKdwikj9H7JBtsRCiCuuBPe
jwx7xPHA79QsM+0jcKXfYjhwBoXE5FFlrOf3xX6I59rKidX5IuTzIrpgRjxDeB+E
zqoCU+g4jLiObpd6jPWsybDCXXOtmDHZH8KpIAV1IvVw9xnvi0RJwJvSP7beGHPF
dK4uQ38jwvFeHxolZmJBmBXuf8eSZOYS8VU1PLwyR2Z6Z338gFcxlHI1nCUfOTSg
h+eMP0Hx3nbdsDjqzV1/FmK5H9tOQV3fOqGlDwLk/BoyJB+QGf0vXwh+nqJj14hs
JuiJGhkPC6CRrnhVw/cD+6LjXT5BbY+BGD/3z9dOt8Jpiu9bM9PjmlsREH+TtqYM
FarPrSYpPTgh2mvMXEiiwv7GVJX13VMnKwONNCxVX9WvAvK6Sw/lYyKVb1G6NM3v
uFWFVb6M0p5JjjhjMKPEthetgwsMXmiXMpoObuhtzD1xpfA/dsFXhsh9ycquwBKJ
imXA/apRe45NbKwrEgV6NZzTl3SV2H26fkhIjkheITV/CviVSnfaljZfEj0q5YRB
K34smhSSm5UROaQVi3Ppgk8X5QTOLs9KpdPoxWoO08FCR0Pv1vT49oBzyaesMJxb
fQAOUijoQGWQx85bhsGeM6l3wIYEhR2+PdV8sExjNI9hGbzJ2glkDUc5+4/XZYWC
+gJzYkYCSIulMmlFnWjSXxUCr8Aw8gFvwvGLmn7Juo1Z/J4wbyS8/K4wLS53oftv
ieKv1Vf0QEOL7ti5zrQrCaPTbZ406IRisI1Ukwor9LdlwRqD9Mfn+qQ0QK9jYMpV
x4ArAcOYa2JlO3HBvNnsnQJ125OqDzfEQzP2rXkyn7UD08pX8GdbPrQiOXO+2gW0
9xzfzeHE/fQ+JcHidBK3QRjf6lUsZPv5+rR2w3t3j4av+/lC1x4Yn/rHJ+Yh7EwM
nMzjDOx8U86LmrbTouUsxSKMzZ7nIRP4OluQh5Z8+6xyCBAjfnkgaJq6zR2mKexX
Q1dRVU1QJF9NNo5zs8oHHX3skxOd69rr9xySXR5cFVj46pMzC9//esONZLAM826C
sRrT3JaZThOHCbfckaNtRE6gGNnrnhGEgueBbReRi1t/uYBzXJxCtDyEGjWdhdAu
fGZwsxujR708bmTGiasj3i+9YhFvqsvLCh9XOILINdjaggARzgweye042ErEXSoD
rE257Hf1MWHfdbKEzTIzNYekqMAUKwjWHTzhSot+10inFqGAG9+kzSAea+8Qw3GH
ZMawUsf1aVQKsqcnqwrHVY3UrLpdMPDHCdtLlMVP8pjr+l70KgDGt5HI3TXZmtve
G/Q0PXiUp+cjICm5iUQZ2JfdQVAc2UU01fqYEqk5rCwGxCv+2QEXJau50+BA8y48
AEGV4OixIoWNQW5RK6o/Vc4I9cfbFkKiIpCsGCBUFBn9U83aug5g+FDHszbuUR4F
lAK3cpeS0PuCc4P5gC80gBiWtO9INgRm8bhpVsKGiqtqtV4ZIARYYnJZ66Xr5H1P
OiHpxg9DvFcPxuOZzV58Vz17zB30L9el9g0I9sWabUhiKax6kI4j5ZEeeiT7J5et
988bxfDeLg4GnnDDWgemFyHYWIUDRBesvUWvc8dlid6H2F0Nj5vyHgCEutLIMX+4
SuacU+2jTipERk+zWCc/KnaWT5nCCJ4pFcJLXxAoOxSqs0tii2AUGqSFZOlgpS0v
7raonD8vzBU7quXIAX4eIgMUNIanhbsTyxvufXcSxHmtTWIepuWGgqm3fa2lk0zF
fgPBIrZPSTFt2Ifm27kuwRwO1O6d47eEt8IOprsSQLr4Aw3XTbSTEtV78xjuYfFJ
YBXjliZE3CSHEa8swRlqgQybi3MC4Pqs19u53zzBJOAUesc0nXFuifidIa3rIFeu
Vna6s8OjRsB5KcLdp6ipSdBtBQUuYiNGvv3/06uhjGhDiG0KzNzCQTMV9xWi1NbP
DsmRZA4FxcU5LBg59JsSLhqhQ4STo1XAq22AUyLDyLK4CTZLyPfJJuCbfuVpRy5F
KvAfxaxC0njCIbRRcHM9NdbLG/MZ8wUlAo7EBaxCefjNyX+GQ12SDoMg6Ets5+we
4WOBoE76aKKqvfsund/65AthN4mL+OeJRqWKErw9JNo2DI3PD6yHS45n5y9sSfO2
wTucCG6sXcQlyGZvPOIufwmnvx7k7XvoQ1bHW1nHD3q5jGysNa8rJa3+AmA+e2+L
qg+yJ0Hk+k+nhDh9Rg8ZnUuXXeQZA5GECWse+wjYtrNZNvmj+wRMPrnXzSNW9mM5
jTDhC+A9luYEAB/kQtkqRIF5F2Fi4zvMNpALOsd4BagpVIDsAX3YuihcUObsV47h
jdUTVwC9bP0xmEsDoaRH1EimMVWueQpEpIGPfx5US5YrAS2dP10WHe5qqVq8icqL
bncyIGL8nTsZlrBkdwsNNL4k3NaDC8s1a48HuptsFU5IZCIDvPzXFikCzOTbcVjm
g6yRhwR2JLK2BfgP1ayhgOxyvr89Q10TOXpVcdcbcZzv5VzPD1YzTzXYdLFWyJZq
oL1CsD1iwR82wzB7rDvWdBZmY8SsBjiHDhElrB603MYEt+JJUYCifnYIMCFvzF4V
RlHhjX34zk3k2MXPvbGUWJztJfLBl3dVdAH1cz1etMBdOaQc23dTiaVwxhy5qHRo
a3HwlnGoTNmq+2K/K4gx9tN8548QcpnKv4F+ke2B2N+L5rc/8/PEkpxqpH3sf/Zt
xJ6Cqf9KSoyn2RbJHliUHmnCtOP1EqCx5BqVIn2F5lbDks9Fdy/5s/YtV6ILnwTe
nGmoIR7eLq+szpnsv+1LHe0Mafl9Bp83h9TFs/FD54H7VKhtmWFF8BW3jsitFIit
U9iUpeHhcM1zj1jt+tTe6o0kml0Xp58pFYU16LdvgGmGYfgvPw6or5Vmeenw1ZvA
OO1jVgYYgGsRGaUc0h0Mmixk9tSl98yUFh3xKIS7lTbThrfrkqST8+aTla55MM/A
OiV1v9UiKxrikpp4XMF4vDcREdJ5YD8ljqW1KTcwVNQo5BViVmrnJmx39trhr5Tb
msP/Zw61lzBaZdkPA2tWjMjnpaIROwJRAkZfvsFhxdzixjTBkat7/Nwy2yIG6ONe
QrwrQqcQwBk28Fe/eMtlzVh3vbDJAzSgCZwbOzWqQBzGSP3w00ERT39bwK4VroAz
KD502rRifwTLCwxsngF0b6E1EqprqMgB4sp07XiM770HJMrltEAKdByoFYnj915y
f+v4EfsUDPVlIaYYU1FviOp2XrtZLjxkzJAGyDAQmw6X0LhDfD7UD+QA5gLt/Fxj
eaf5qbYxjrfgjsrKlmENv4+qePZVYLT3X8WHlQunNNYUIR6kJUtr0Wxq68wAx0si
F2xU/GEymz2hnQ5k65IgvW55ShmnIqzO7+ZaKmV8GJj+6Jn/FkhVyPkcpBZvBlMT
BCfmctWPy02xyKr8sDzClrNCoMwryUn+i4YKPjZ5V/70tc7fobAkdWpMFpzTuXKz
j9mas9G1Yv2voPMhEas6/Sy53gnEQl+JiatAZ09HYKBbRCrJBP9LGHbmUjNceIby
bOF4Cssct6Lr7ez4tUAaGFtFAY5J2FvAB6h6c8zJS1pB+cBmWDw+Yb5wpNGCuial
laIv0yxurxAdcHNIrbUnEEqKne/pfMIBVIolRvkjHpvsY+T0ZQsYhvd+KrOYQBd5
igfpyR416RbEVdFINOsjUt7DtYhfefIBxYGO1d6EttwMQMQn0oR78fFZ8kIBoumv
GrrK7gkOqXk86xD8ELd2kcNVcJOdZEkLxDgcPtZqSAqsis/2YV3uT5nAtz3kw6u4
nnNnPjan7BO3nQ+fJREHCpyOiIJxXg9kD+/H0CZF0OVT5HjJ/tAnsepebJLVtPsP
CSTBZbJnsDJ3CeoUy/x94skR6aUqHOK/9iNhtG7AJX7LtPVE85vM7KQhkxJYzHJf
pQs9m2g8PlPXreBDOk6pprtk/tPFCmhwRfPXfX5Hwh+TXD/TCMkMTwfgKqkt7xLT
LILCRG9eTq0wnAdrb3YDsX4IObfKD/0xsXqe+9AI+mKBXV8h4oQKv09PHJW1YfOx
T8L2TEknBxpcTINydXt80w3hSECwreTMAuZt7uAAIi18gZHoLrXf6L0rN9C3IDhJ
6DcUFtb4EsNRwKFTMjFO+6DQ9EBuDJPOTZtIG/fWO5k2Tc1aELVeN9mfxHV5wDqm
RDQhGGQWdkDXc78ga9fEWdO709XBOhhl57h0hz+G2wcai79j7kjNocj6sotzvuIP
NwXwhyBOPfLoWGAYWXfSsTAsK2u4njHSxR149hAXwmKBlyoMENwMmsPRC8J6FJ9N
hgMndKXebZn6XIaMxdJP0VmSov5je00Amjo7Orw4hJdSTdxyMIRID9uAz9MEDCqC
wlKTaAwKHb3P/9Nw8ft2yFpqkSa9B8LFyvtLiMr6whqdJRFrX4WQ3+XFwdCDlQf/
WHqeDJJ3ox8kbqBlhnTWFL2jsSI1tMmjfWHpxcrS3aYK+5MPJGJsM3K98ZTQhjqD
8X4uBlJRy+4w+ajZ2ky4vOtttknfKWn380yc2byvL0nqZ7vb76Fm3vj3mJxOQj93
uAjV3/ZiM60iJyhOs9jw17e4DCw40zDhn9oR6B+woqNDOHbeuqUnTkkCLy62qMwM
txS424baTRqSU3tnybe96DUVhiXJSs7UzNcSIGqrJXX/cxwJCDaBNSwWDuR59jPK
YgyNwFDXMEX2EE5cE6AT/fCaQdM8Si1VU6/9YYb5+ce851JRAALm/AnMWPXWIDxy
sPa63ByesnfapXpo2U71QBO45b7qgBczv+dBWCKftpDy3WY+CwHs4PinvulrBdjV
accDPTtkX6bPMDDmS3ZBccmixVRj0fF9mrTNpepTG2E8eBjJCC90Z/iYKkC/d5tj
qJIJo+6aXUr+yUyP3bUPt7Vnp4DF1c3J8YF1HHyJCvv9JAi227BSmBua2cWouLhX
SfDe3Yj+4fZfILi1m3wAJzGwBVpMIEVn1Uj0E9knCwiMnwgbrlEE/Pv0hseXcHbx
TDF6TT44aGQmExk3qyVK3cIUgXjurJ/Ji6nB4HgD33g2QDQksbw2IObNrvmgVCvR
DnH+caEPHWJtQx0OP15NH7TL9DB+C3YYOGiWn+euzYFiYhNtu8anit6vNnrAXkNz
DUhOu/YRIVbkyFR3FDNJdim64CIAZblEm8lpOqKfcYVUfKHB/FG2XmI4V/EjOZlV
CBxTqPK3dnunN34UU+dQzjSoRnQNB9dFdEqCLcmdhoAm+oxlIw0AMF4tungPlrgo
q6p6OG+Fae3/3TUEtP3tgohdkh/CIWIdVVEc5Yb2AYpNJwW7Qy/78Wcdcd+TXNaK
Lde3UXnVkn9xNEXx2OqsmDFXcZ75cHnJILukCDg5VIcAjzA+HDMsAszs2p8fJ7vD
S8ZdDgh9TsmktBvdV3qQ+ZERuYfofH0iJX2Q/ju648TuCSAu6uJbXj7YzsBX6+iE
J4tvll9bYHt/I8trT/zVtUCpO+gd3iUtgR7lvlm9b89vSYc5nbHlnz/3Rx4obKvS
G0FBiyGCDDLTjXsdpG3jJxr/xtmemK7Bu5UhVrF2rP/9Lbs1Re10JsejlU33TlSu
WqAuyi2R2vQGCUrGMM3jF6843KaKBEo41y0tHcn+Ln5x4ZFySFd5Mh+vmKhsRR6W
YLFBVwGWaIr1/cUcRUPCVVlH5pP3wsGmZCW/9q8khj8tW+rj2UchyDOuxIilQOh/
/3RqXBJTzT22e2dsUatlQD44nBkzs/abS4922kjoDo+5+bOrfH3b7dax/jWxz3nK
PSt+1eDsS7Ght9otGQqBqNi9UUZk/SC0RX1emlVDSE+zdqIEF3vc/N1K5qYG6xpK
SY5JKlgGzVWyzzS5cHcv0uMIGlL2sk91bU9JwpREe3sYx99sQuW+qCeN21ZRkGnO
KONOG7p7I+pBhDqRQeu5qybMlwJqhVcwvInz+Y3H6rkclhBXD5ghDKEDLb1dv2yZ
5WdDCyARmhj7lLpa/BBWMxw1scZHOgo19r4yx25V9XjelFOptRHm5tp/8Yid40sH
mOM2M00TRWVFlBWRgB7OezV+QldHcxAYkPo3CQYAw0RPb41i5TPVW2pTM0/3rKDN
gVMDbr0rf8WUKoz/oStqyMMInQuy2zsYAwjOcLTRVFSmn61vYdpakjD+4ol9YraE
SphrQ78MzWEiZRH50txtnLzMuln+1vVI4VRBI9TGAGJMpuVRkE3bYBk6WbQA6O6h
aixHNdo3I2TboGKbsE7RAyi5Nw81K0NrJNC/Hm+fV5b/zvF8XNa/0141C1PQ0Kg0
wkjrV36ogqvqIUAvHKHsrRMr7DeM8eL+UljqWBp4UBgpy/HgKkvSq+1clVRKHt2X
lsPH+ITdScGQ/wPtw0wLIvmCeyaRlP57w3k0s1gfNw0uNmGTVYTt+RlXNPrA6gpK
WvXuMIklcz09PMLa3ALxcLrTzCGh6zOjECrzURGDRW7JI0n+rMLaY4epC0Wtp7WV
4xdoPFYTzpydwet9EEdVwKe50MD0B275RVKyjT+T2iM0+H8zQFVBW1WiwGCaLs9z
Z2qwNH/EczdxZWUXuw29NDupZHZTAoQeyjfFaZ1jgpM4T3qKt1k9TGjfBaWgkwN0
ijV3W47fisUI544jSJdGFb3D170r0PiOO78/ilUhsiz75ZVSHO4ODIvMRbrXfar7
KokRZf1H2jcMQR2ot8zcuOxc1v84FcyW3NjOS063H0DYzK+CMuSSd3w7V7JBWxHA
qQ6ZaYz4eTbYO5GCiqeB/PQT4n2XxbIPIR4DeqxIOOZsKqG1g0PBZ1C7Nq1nqhb9
qgxEgLbfp3e38JFNeL0QlUJQVKDX/xBwtsN5DU6JiaX/CBLvlJgsIGAeDUmONoo+
oBoFx2eW7S11LUTo9ef/2JAQxBxmCPgTof3G3zZRM+34YSNaCaiE9Ce2mrXV1a89
8BbfV5130yaxpRKrNi/7GD23sFGNVuF4uzyk/YgRAnXxUfppvT+XsnYQ89uRwnGr
7j3Pvg5xEkC6dg5hh9GmOyu6hXreFO2FhkFoVcg2LtMgXmLElhx1xGyhA/hJB20O
qh5RVvpEu7our5cD23JpAs1sIKbrwAiVxgbBw+J3V9zZH250MVx/MQcl2dpmOY6a
ghm8QiWx6IwpM+DcA19agdAHQDhC7XmN1fKFcY7OKDWR0eQ3nvRq/8L6O771sZtU
Hl4A791SNsZuHPxRIlIzcbUGxFdfVX+Ge45dVqjKC8t8JUzZLYc50xffeVrsa0of
ohjBg2B6zwNWGCUAABWaRmB1ZuqwhXXUJKEG24MH8u6VADrQOmprMwNTHq3PnDhS
+Wa3EtOwI2zTiX6eCVQ8ugQTrpfY0dbMLWk60PN8iSXVVy0UbaSj12HYVQntnALh
EJtG/g70RX/5XYP6igp6xZCtz1oTYpP0cVmred0fuRSKqUBkjGuhcTcBiAriB59R
K/hRIjA+mRHidOf8a+Q+jebhuw35jw1aQcrkQ51+OWjhjv8R+tkZ8ZR4jxOjFsQR
v3l+OA14G00pyAgMxL4chdP0pTgIr3RQNHnfqH9vpXzChkk4xRSPU5it2TUFh6pi
MavRsKzlE7w+ZERySnji6XFJxypgd3ztKaY1s4sXLt+fJ3cfY9kzVm+mEL+higr1
g9dL4NvDmdAJy5q3YiKdfagmsPOWFs2R1xrINGyVcg7OtoaH7oYNJKWtjTKKafyR
hiTsEiL/On9c9RsfgGUn2sCPIyccW/VKUv/srnkCc2A9KRdvCpTU2SeN8a6D6Bgu
3S8f45sVSkJiNGFUMVij/B3OZpPC3ayZaVq58T4sFK3vFmsnKlgqd0iLwBSG/7e5
K7i3iRNon/73RjThoOP7YoPx3Sh2DtkZl9ZUYuXiKIvJfOlRqaEPeXaKbwdWttzd
MLZeRDN8Raqe8Wq7J8A0/EjXkK09D1qtInbx+PYA9gPb3LuzAOZtSc5+UzCBrOaI
EnMjhATvieoharSMThH7aMC++aBLQp7q5+rcVJfnTfwhvLX1xiS5D1OG9QXVXsHD
oYDV6g8agbzyUdWvp5ANDCUQQpiwHQVZl/Nl2NQ96Te1Ku8z+BGkyk5BMUX09M7W
t6Afpd4+jrUNsOuL3sDxdQCCEs/WcCLC2yWGJib1uAkVn5MqDTQJdB4aSuN6ByPh
f86mc4CFupjF+BPwrEFPPlbNKYQP4adOjnXBvH/ckIdakHdQxHapO4fVrTItnMl9
Gw4pPCckPdVxZfhgPDuwCyAA/iTcFZV4eyTOXs1rUYxSQ6qQJXp/4g7W27NUm4o6
y96hg4fm5Z08HoX8JSBZc0qZUI7uNw8A0dyciatpOEWIJJPMlwSh4/MLyF0A45sz
QyU98fLWeq7m6Pvtig1Pl5bahXCKRURs/Y8MyHs7eXq1uvgo2NXkQkOI93mPj98T
Ns3edqD5ywa2DbNDpmNYPKC58xwvmTGIzg9w1qqoUT4mhU2BJrD6zshgirToNZQP
+02fpzBwagZZtrV34TihflMomQ0k21sieLqs2SInVCM1rNHTE6ZNzuxqReOb9/un
LIWpe2cg5RTePjt0FREICWM156o4KPDjatuHAEV/IVSJEdaBystwkcQF8uaV7L/v
TU31iPsSsMBj3n4dohVnWbaqh1e01xEKDHNr1Kt7hBucm1BFWvyWJVhFOfHB/IbK
7udyUerGEKGOyXjx7boaRlRGF6vFTvvKje6jsvUvYd2WhRIX4zKYQmDr4hK4paRp
j2xEI0C6KNqroCAcBNoHURixnGWLRPlpuNyynerQrUWZ2KCq62Wnb8p5ZsEcoHUv
Y/6V3p6h3pdSPVoqQpvc9XsQNN4lenKSp2L4/HCpUysHCRIQpYErczMDOpXZtJpJ
xRGPEqgfzQh5piZZcTNJFNzuip1dIx+qbl1naOEnWJc/hdR7vbO8JBkLa1i6zddz
5pfKKqm2f1LibpAFSIIr8bb5qyctngpbN9yaBnKtgB7rXlL63X2X/VMuLKHoq1sk
SYy+3VWgf5FjEZdlCpEhMKyfO80jCcEcO2UaBQi2MTJyETEHR8QOhxTc+rIaT12f
aD5cxbnSBlWElyFwtqCloh7M9FLYIfOMcFWAkoJLm9zQdaX/hoVo3ss5yKKzlgk+
oHRLf+W6HCA9vAX75ECStUz7I6H6nYBfmGj6YfGTpzotltAOhLqkkkerUVZXtELR
dLacSuw3jiJqIAZcM6ocPHfOhtnRwC6h73v7kyOi/7gIiheTPH7ehvj7qCQz/b79
maiQGzpB5Bt3P2YQA1hz2E4iU1VS0+/TOIh7W8pS7hO3jyUhPkgRqI/bytf9RuCC
x0mya7WGtofIadkWz73Wo0MUS3bTlJNRlUYBwlWBDKGABByWDkc5GrTdh0Z9l+PB
9zZRYbqzy9rrAo6aaqIGdbYKzxqS3OpLNstGbndqcwilGEjWR7Vsgqj2v/Y2VqrX
6JKYpjpetu1UCzSfUKwhhDjpQDni6jVQYUuAkIg2oTRD01iBXn7NOnq8cEqsbJtC
Vf7DUorsUvrNLJ+5oopPrp7ykRcPUSiJi6bV3H3oLK141ncF2r36txo+S5E2U/ZY
R8S0Yc56KKeWTdoP3qbOPDxs5p0xsBFf0gpPJBy++LGPQYDbsqX7H6jFCYqYLKIa
YpT1EbMwBPWVP8cAlMB/DObvMD42HGnJFz5FkAEpOyTkgcS+OkqxryrEEXLj7AzX
yA6QtEDLUOkj8mIbhrr2un2YcU6od1ywlMAS8SknBZhKNa1wKIVclgdcr/1ukvP1
Kx/YND34OgIT3npcy8QcZrCZu2oseVB4iHWNvTz5NrPRD3fY9HM2XQGDe14d4L53
vR0PEdO/e9hLGvAC5O4mUGnJDwuOPP9+73v3L7XWl1LqgEfYa7ijxEzGufI4pJSH
7+AS8qwJzBNb3cwVzALAIqGnnNpgWLnnDfutQfxLB4b3NnJzgM53pIJN/z5s8+ud
/tpAHhFqh5jdG1r2B9ZgMR5lT0RLS6xeLNm4oxDojOxIeGS6/twxpNzImYvjz3mM
mm6j1d3UyGoARcxREDwrZebAYNdh/47vt8Pv5vG2MGa5hXIY/akdsVXOvRclYH54
dlqRMzpIesBZgFoIXQJjhPWsBH4pp5XJXMp5IP0RQD+eMm3gj4I5+MU+W3lnpD2K
W8kcp6Ax2t2atAfD7Q01wVRKn+E/LxS3eiy5FX7Xo+Tb7QQTxoFuE5MgXm7RnnKH
DDJj/dzqEsuLSpTJoz4TDqz7Z5n7CX2bnnbqe3y1csC7wyza9Upk/zxTAoeyoqiA
xyDfQI+a9Lzd2ISRgfGy0p57zOIcnkFlZUYC1av8gHptRR0YB9gG23XSMH9txF9f
TrbpT1kJzIH4HOP0qWxZg8RsBDmts/fkRbla0zTNeDxkpAokyGGpIQbn+l7a0NbD
qCcPBnsEpynfdK285bCXrhM2HwM/dPvzkOhZxhFwmB8v6+gLkv/W0iWryWZ1t88J
mdn2Q452ah697Hv4JOjhnpCU8cmfrGktZN9VP6A7aZi3uL8nuZPEF9ZcIQSTlDRG
0lRGoelNuyUbzE3jVKdmuUzX6Bo8LZzPfRbJtnrf09Lko7ZR9IjFwXknKePr763P
8oPoaRgeifhn/s3H3Pk9pzprppfeUgZjX5WF1f797TtcFWw56uMeeROB8vzUvvCC
SfaEeyAfFTCMGmLkKOvAE+NVoWP9XjRj/QcKDUwyOYs/XfOkj9CewKIAvYXMr+pK
62yzFi0qBuySxdk0cdR4l/bROqzLgRPSY3bHs4ULpAkzmWMI5LB2FoZZf1oo4qf8
8wPIR4xCO9TeXdfH5GVvohUxv3A1S1umWuZ3um+6xdIqOnT1rc7QITkbN23NuRx8
DpmoHMqUDPUb0KKjjNqwhy2VxfrFR9T4A8XtBeNGggHUjqkD9fJC4pjYHZDueKYy
7N19bh841sJQPD0h9YEgzaZ7dKEUA2tEZ5j8seG2rMJUAzBJa+hON3zPs28po26U
CVXOuAtICjECTQP+hJqvUb7mQ/jiAhbiukj64ZOyeYspfTYXdfhiPMv2dOy0VAzU
gNhHUEr6SoKMhs+snyArytufO1h18KMuGJmV5rA/57m2kGBSaaLC+hXQxUSM0biG
sjD17JCwuI5mo5QmTqg+N/cVqj3x3DToQHHOIHkLUqOx0CX+cerf00JDEAbXqNFh
TnSv4nHDyRnDK0m4U+mrkjftCePeUxO7uwf8Ex7QlHZzJB+/EwBZfCZ2GDO5r+bH
q+6ggzyfrdIq4huDKFucAvmzn7wqVitcEDBbKnPEYlEpFOMUzYdOamwXhhcivBwo
idzxu47/J7q02HNIg9XkUWc5H7yDPNjxbSbUNqcf1ZTf4AJ0F09/kZXdd6Q9Vum2
/UHN8PKNhpLSM+SKljpHz0CJgxBwQQVdi6WDQQ4clz8mJ6qjzViSmj6a7hSFtA63
ZrmqV9cI1AVx4QJ3jaX+Wrgy5+acOQP/kxZjsg4T2qxZqQO9t1LmGvHqbQeQZmKw
oFM//ByECav3XaBP4SNk67aI7s3ex4jWPnD6LILUN34pjCB9zsnEYoE3LGowhpIo
pXEPwI30ppD4C4z3aR89bPUXlr7offMQg2CbvKl7V1JKBHXTxdKHZ0utop8sIEJY
5cRqQ9teuq+nbFDGesroF5F4fgC0ExOCAh2GoQGQ3SWjwmsFg19Gh7GjpY+DXK8p
ShYvJoBi1m+3X1iL14zuIHrCEnoWZxdqUjjfmTaLRnb72XX1iKJwlC63XTSpAEeL
4bK8kUSri/H/VjOu0da0VtNJMnBDMVoq+UhmPk/F24VTM6Fd11KQL2ObW2U5T50M
AS3jR8fOstEtmPvEYGKHNIoKEmzPmkOa0hMKPR2MHmvJyaravmBe2myDEAFMTC9o
rza//PJmx3p1p8jLHZpXd8qLznI5ex2unwcMYdmjD/JQU747x0Z7Uh9D2qYbXjpM
yUa14Q1P29rBUVAih5NkGyXVn0pEnUjDBxkhQXkzHrwRagXBKK6V8qswFOJp2XkR
4L5FIvot3oKWP+gnKgdYY0LZSlV1hzrmeXMqGwxSf56JvIBqRdl2wtXojxJP31Da
tFH5KZ2W1/rbUHEe7ORZvuqvD7ScUrwpbFfm50paTF80aSv+8m7hIafseh+TnvT9
IqCJet561PgUQ22klqsbhdq+y8ymrn29raS7iCUgQ4KpD56IPlpl2HU9hXeX2TSB
cUkOgnkpSPhsPqtg0/peDFWe+3Hq2NUn96+3mjhLNbvNrX7nmUT3ZN1xKI/OxR+E
jsZitgR5CtZ99Ccnb9YZ3xAh2QmF+sQXN6t/bAxNRFMRVBSnalZDaZa198iSviLB
dTSqkKoRslJRm+vzfkju9UMSn/wn2oLiOGPUOENJe+owwEWo0kdl5inhZYthj7OM
I5+v13EXMFBbvTgh9eDNvdQ8TgOki66LU5YJG1kvKibiJSC0vveJUpLDi7127aIW
WOJN/YAT97fFaWHrb/U+WGC0552gD5hBvmI8jNk7NhQuJp/oj1OWWHgjRhK5h1RY
+rtdeiU/fmBKEevdhspnijatGehbS33qIR+pLg0DuNam7T97YFUuM6sZNv0udBgQ
/qTiInkRlDl8qkAu+W4Fm+OcrHUS8JDUFHDfz++MZXWVjlaGP6DSF/zQe5L1XaJY
GFNMW2q11fD7Pl2GxejW18vHt5xFIPhEj1LkM94gduYC8U5BSinB3k8X84uahXPt
KizMYcvsLAVL4ozJqehmQc9kIjaOyuSzjRLT5ptloj5PIPxHUY34ffo9rqjJwAcb
jbuYEG1lmwgGxHATyj8cO/KWCqYwAvvzIEw+XfUHopNZpsjxIpT3Mct/tduRFXfp
unNwZ1SL8wQH4MZusSoXrlwgyCUIldLyY+y/ZsmwzOoAFFQ1O7UQROpV5lo+T0fh
MdrFfdDlS77Ddv7l6WeEpdsht6V0nAx8sOzOQYSquc0vPaEVtAFWAkkbjdbi+6nP
odlyswyWlB0sNrd/ftfic4Hd+Z1Vq8B46VyNdp/j4T8VYBrHYHfecYY4ADaawXlq
/RWVz4ikDV83Ad75Xn3RBmVwzurtGIdv2a7Bkax26VRQttOdshsY2sJaikwbep55
j4swZXHG67+iCrbTiRFdda/Oy5DjbHdxGTQyV48wNPEfTlA2bXKdvU/CeB/M0zuj
KbytT3HmPPdMmItZwuiXKds7V/uEuz/T2/RTZZf+sZ4/XOay0carcEE9u+k1E8yf
owVOGCPa40ho8/PIAKIFgsHmr8ayF4awB9igpMDo4I5Rmr2KCKqqH9lqn9+J7vdO
tB5l1/trc0gLvih9xobQxAeA1uCMzM1ZxJiRD70smfJa5Q9JrY+ylhLZd5S4rfYn
k3efj3TV+DKc1oEkvWseA4Zr+BasqrocZpZmgoXxnF/PJWvORT9sYjPvTX3J5Dq1
9LhlMCc7Zqp1RlOJ05idhzMaHYTNBVGVKoCBFygpoZzaDzeILV60yfxh9i870wxv
uVUfAXqm4/nHRuJVr3JG45R+8Z4x1ZUOa72IMmp9CqtyMMiXowpqyv/aIZlswQaQ
UnNDRPYzb23REhSTaNvZu0tKF8ij25MgtsrKEwen6O1436EJDvc2WLbz6VhEt8ze
3YyMghioNk1p3EKL2oVB0wFgzMaRNSGio6ycC6Yyf8fP+Hmrpgf4p6AE6D8qk2Zi
9pcxBD29SKo8dqsJuW19wZRwo9hRvR+En5NnIyAdJNN0r7q/ALKzO5VmeG0m8doV
4NdE/UgNcYy0W4VJjdxJ/mtIMvNpm/Lwdsumi1D49OB4LJZfdjEmuuQCK4uQtUvX
apv4NEZ47tA0R0yDcBJB1iTcmqvZCBh4jQ4wp3jo5qAtibW0qtFtTL367+N6j30m
CR5gUjOfdSLpBQErIcR5Ry3lH0zKkaJ/ZyHmrJLXGyjCzSITIHrdnEQXnkKCX0db
0WXfcn02efPpCeeHIXpiADUQuU00a91i9Q5FLdEUm7rTQfeFVIuYY8cEFQvwKLX2
EvuSzCMBTBvPoewSuYkqLx0tObxdTN4JkNmbqpM8XshQgASCKJ6Bgj9ygvLv2A04
RzcMEZJ+SlHuZHzV6sKvOEbwZbfcu+52E+HQSy+HnMZ5cvZSupnIjVACbhHt3e9F
P8VqXhzL9fcjcyOdIn/rYXTi5LItkyMZ0iD7PWXDcA0z+5Sr0dJSQv+k80DuWc/f
rex0V31XW66uaST0jt8HanKAjTtHjbsD3mUqh7Rq2X4Yjz3TLxJZi/iErsjSWrFk
2qQZ6mRlUaQEksU+/ChBnzKdoW9xsaOQOuygEA7gqsALgwHf7cmBHakABRMLY8S6
kzGNfVASMVoRGJAYBmKiGYVCCDM6xUbEZnzM3R2mTasp3nEz1qY4i9C6Yxy1ei62
e4FbNLioB6ozTNxopi7bb0+w430AAcjvDdfXbciwkDFo9IuL0OXxv6KNmIRomdXb
bhbn7D/jlX8xLUOO0KEbePcZwAQZY/znXPZZJZpLmA7tp9i/VT5iANTdOs//bwfc
fZEa9v/pEkfWwfBO/LETgn1GXBdkNrMglP3OeJAitdkM0GIrb/8lViQlGbT/iM5G
UzO8M1aBp0pYgK2VTz8kidY0aiA0TUGA9oz9uiaUvb/0gJdl+rgJOIJG5PIicmwV
NDTnHQBjc6guP8UqDk4o/8F2iaTXoryyQrnDh/Drf9u8SM1P6JJ8uyerh4Oth+Bv
64HReHjejZ4rfmKYfqh9sEMFgSEsmzHQzNdV0RMf/S2wz+oLlatanX1++apaer/M
tAG554NEGtJOJpd9ERsQMJqiwCvMJOhLfn7DSmgK1id4pHM5nL1UW772kBOUzFJF
6gRDZbauQ/J3o24liOW4iUqfI1K2TEWIqpIUYWX6JgRSvXg3ZK+m2pu0aJVgjB2Z
aRCKv6Yv9KsYM0PeUXlbmSKuE4l4ZtVzFL+KKoy09C0SMAZ/NAc0PY3aGiLQXeb2
MHhekYywKT05aFJJLXYOdD6EgkojaLgIkI0Dai8e3JK+DY03dJCJ4WH8tiJp/FIG
pmVcqWg1DSD66p7xzGfTvqXMqxrdspaoLxllqKpzUZKL0DknC1v/p7Dz67gJzR+j
jCpahH81bhAGEh+e9F1Y4eWqCya6gmWRIgxNYspCGD78Yr+SpvrKboarMq6psvaa
MV51iNA75Slxqzr5vqyIhA2QyjaavvUqV3wal2GjEYeLdU14va+wLI/8aWnigJpH
s+rZIKg5A6O3Z75zU+Bv/PQS5o+qQdGBcP01MSkrkt1fYHaXtGuk1QBTmyzpS0Nz
rZIXuBCuekuYLFTG9EJ07xIEnwKAl8G2vi1v1DLbPaNSeeC9MLaXOMF4fr8dngC4
6Wz1/ADK9zvAP7aPO9fURhcGLfXhKHSoWgsrNbZNQXrJvhRt8ye0DpkvmPOV33RJ
WyFu6CY6s/qqUR8ZTKOZJKxoGUfDTGcuCaUpDHD1ZtIP/T5Bk3wBC8CE+sLTIWRt
SXezezjinCgqEbKpmUvcS5E03ichzxaO3yc7VED4deMgiqrij+MnXhdCK8N0rNve
FooyfMjL0K8dTxmB1+N5yf/O5l2m6WmGkXJWnw92QA94oKT6BuVfPaDgCnzDFkJ8
Cg14h0LHzfNaBJndCNyslUkV6SD6R+/E05ciovyNDoMCYQcesd+SXdS+6toSu2j4
ilCWXI79D7jAB6cmN1zpj1i2mnRqdslEmXxYjl57Z7Rjf2ZT2zP69E863bvFitKh
r3XAse5fJGSSc1m9xlzZSwcHVRdSGZuM9tB7b72sNxepV4c8Rff9ZTaNVnxicCad
v6gI7ZmV+lBaa38z9xd7PDNafEAzMxSEyQ1eEiquq0lhTVucCQk/xIwo5KHc2IkQ
CohEkiIp2jdgjuXujXCMy4gt9ihXJATmot1iKcOzkS1IbiCJdoB13G4rnxs2uukZ
vSPoUAMhVNaT0eo7XHNCFobze9u3pIpMjrKp687tHB/cU8d6RjfHMWZZK5Sf1sXI
UCk+UMSkiHbm6257du5nI7Jd80c6fhW8BAbu/B+m8XDvoAdYPIHAOpQZ4khLy/LL
KdgtAmvWapQ1n/YtPCyugohS7NNuxG61VIqgfoDffTnRYiIoBXwkdZa9dylwJRUh
u6Dj/ot6gXtZdCmMojtQ4pUZFd9OX0zAxILMvKL8IB0xbCHXtrYBdbBE00Q4PBHr
2pCfMcH4hVPognZGM5oLxfIIvEob2Z7dwYywWFJGjpqn8lvosuePJXTu8b4zyS7g
WzLf9KqC1at0/RVlcDK+CFOUcCvi5ArHLt56z/5NJ6lpNuxe5aWeLJ/rxFJSYhd0
1OPch5hqvJ7tJeJiH9yvkhLbAzgMDVngaAEO6VHdeodK8jlTnADcNDjJlfTScOkj
+u3qS5sCEX2U/Ja1cT1QLvae8CN4NXCOvlpXlVqY5sk22vj/Wfw6uCv/bzHh4YKA
3Z9CMPILpSswuo3tBC6U6jnNjy5HzfJkNfvLYiUNSfONO1wBot/7SOOVZtsoGcZq
SdDz1qd93qzJtKAeOylckGVw1iiYaFD8KwUW1MWO7LNA9Lo7W1MVeVJgNfr8MP+l
LP+gHaRXD8KcOtbyGR/oLa/05Xf1lTY42MRQ7Y25gBjmoG2oX4wvLDWMD+ZTgB3B
Gyz8EFwKPN5ZyMEu9KWNqUEK7JtVpsq82sCswyp5aQFJK8mMK9EwNaOTb0k1aQ5/
01i5CXyf8sjBt9z5kGUVij96XuiVNxnzlBzvjOGKdyktyemQUCNGzrWmTEvBdpmC
gRhtFS71ABw8H7n7ut/L3qboLKQDUZNs+uNmyFSOLbfVIJhE+Ajx1foqK+oj0+aX
LIq+Qc9LjOXS0X5Qa8Uykk444GI2TJLtv6h78LKnCZNmxCHvI1Vzuh1XSmY/Ys2G
IcPNguHLIiXPFV3hjySi+v6Eo4FELojbMV3LhvYNrue4AMwOKWr9M4FpCVlngEeW
bxS4wctkPxieFkO1rM9siT1BxSOe2hLVQnjaR3dLIEfluwNJAs1WpOJV5LrmfQnS
2Yf+tOWobQ9t6M6N/U1+y9G+xZ595zrxB2q6gKIE2Lmhzh+Rkfy9Hwtppbo+peHk
lL43xeN2+6vci49vX4zJ+DvVkAp+1ez/BeKBsYJUs7o/vt5CjXlffBIkplAqSjVr
XH6catlt6whDZUAsG0ZIKE+wZ7OAyBax5tW9CFYmhSEmqDl14+n3dUjf9sZkkSWw
KwVi5UCb7N+on7oSdB70aaWkeFmqY6h/nBBETo4l00LWPc5f8LDNasT//hjmEJLM
yzrf2hEk4HjeDE5ITkjOUsWOFuXZM3sWLZPLj47OUYzbKsFWwpSevb9lVsQYb6JI
ikWISKjuGCHk/cFx4RjqXqDdQG8k+wMB/XwpijFUUqLMH1j5Uqb6NcnqXGWOSZER
fWSoQ9I8An6WdxFxAo2o+Ng9Vx1Ey/b7Q6av0UN0EuWw0cQsnFLeyL5rwAQWYJfs
kDpROr/J2TN/cEfOBff0pzRWyiEKhLaDb5YEtTOrFs22e8dSWuIAiqqCRqZPRnwY
ux7WZH1bprpvqutOh9P/rLZZ9DtMd+T/Jb29Xhus5ppHEaLK49vN/jEgZvp87jXQ
LEYVUaUGN5wj7SfiBulOGFa+snrJjC2a5rkqBqn+YZYlhaddeTtdaJjzCRk+zjmC
GaKhMQ82NQVgnaBhMvr4HAJJeGj2H5Ea75guK55U2Ex5y46/wkMMSBwWgevGZiAa
9QPO/QmzuSC27402VlMsxuwp6PkUuRP2Hhq4YvN4wSt4b8NwgkbpaiIO+gRUaX2B
szhDenYQ2dE+SYd04gKqtJRfzDJKTKJQY8HT0QN4xex3/umMpsylhcadZv/Zoco2
Ey7RtHSb+U6cXCYpZI2B+bXHwObV7Y5cDVOCydELN2wk2U8u5XCi9UMz3fXxX7zg
eGoE11BVUvd2DrUuun7GMkbvdJOz4YKBwo97xF7wkE8iX0pGpaBZDJNr+hHl4XxK
dMFqbdQOnUoQEzwhDeWcj95RSi0Hgg9UtImL6nJuNIKMxA2D5Ph5sFCHDfUNhqiL
H8ya+Er4o+p/KPd5t8DanyvWyWkwX/8Zpmk5G6U62iCDMGnoycQDtR2TWgeGBz4m
06nlWg1kct03zXazb4gTPW8+K7hZTj04ylhElOzxz+9KxMAGNJPQc6fzVivoLQsM
jci6i+WXrsVow7ijtG8za7+ZvMwwzRTwGgY/fJBPFx9wLicujAMtBZ+rfF20Dtpt
YoFw0avOGWDPqiFoFhvs1CrU+YLgMDXfYXDMWz7qg/WydK9DO3vu+DBF9WUcUS6m
2kdWGoJdaeZ9y7XrC97VZ5/KPscrYcZ9Zs7p4NDJ00djE543DfJUVBqpe7Uuj9zI
NOnL8UTO2yIlnK0HlxGrZvDk0soAwVNKMFKA/oVUOi1aHjnfPRG+geS/JB7AE2q0
YGAhUX4AkNke8DRZssnY9VmdQSwF88ZpofC+SMoCV8XqyxDZYj29tWYmOqFq+5/O
xzkMaRccCeybUdmi5TTkVr10AbMPU70jMmUtn+QLYtxjIfeMr3W6VZDW51bV7x0t
d7w/iuPbuOwWhi1SJJ7gG8opmgdAvQNcrXvL0E2Ava66U2HuVq1fcdQuB7Ey3GTK
s2IyS0VMYG3ZfyWTFTDBDvsmgP68mSSeLm5zHtLhA1x8wUhdsZ7crnyMP6jmpV67
qwKtoMM00pF9IpZqD7C8sHkQSK4nddeALUYn7CwZRm4oSKVcEXozneWxzxkSqh5T
ImnsLQGI0hHUdWYub3vja+ynqziWKamhVkwmNKBoolNWvgwX0KZ4Q6D+MIGfi2oA
wQjrpHJwfeceKoltFfOZn3680Bgrhj7C2noZPEJx6K5oYc8SZ5rZzwS8jgGKi+sw
OINbhdB7YayWPLys1PjhYsFibCOurS2cClupwZyuVCER3yoRrHmjcEStXT0b61OE
lyc1R/SZ244VBb6pkaLF7Uxe/Y3tJk4yDNPp6+lgUQfXTBovxLolKkptPebaOfn7
F0tT9VmfMEM+P1gco7LJJopDrQh5DJuKc/f57BuB0JmJhUD0EL02elhAEDcL0y55
244LgJY2IJAVZRzdBZ1SEKjk1a4UAvlYRYYckL/jbESf7P/s/Md1URd2sVWXHE7c
lY3+L0ijREtQ4FoMnPWmDrjMeQsZwYdE9nX2iF32SlRLnAtoVLeO1pPw2O3S+i9d
CJemHiga+bg0rhokecj8v3lcu5Yf1JK4egfztZidDR+3DBJ4Cg/wtI4XgilRC7xO
oXD8IFP/Pk4aaNuqL9ZvJBswIaqxHtt7ZgfGVnKRnbckz9ltGLtp5x+nKLmIZiRY
i0poJM+Lh8zxgz1tQwO3Q+Q6HL5Ux578GtwCNpfFZ7hwmNQTXKZF6XTTZXdqKKJq
UShbJ4Mg/xnoT5HlwuOWK8lwYhQIm6HlUHFjkErih5ZMGuizydyylF+1cb1lEO5o
05hWoYlWSLKowNrXZ3SoJSaugaWNf5arHVntOLX0BJKCSLHjEZ0a5Th12tJi4g0X
L5jVwC4kPbsEfDKTy8z8G6Wr9uGxKCAxteKRySVPlFcSl7YH50roT7DJu0tVwG+D
gLMueCSV8RKIegUk20zJD7clj+vTnEb92Ni3GlGe2CIzxkHKSReaiiUew+4J55wt
iWaV0EWw0lIWQrl4ji+x80IS5M42sQteiGbT9sI6R6YHtRcjdx3TTwCWlHdIxRoH
ugzNeB6+zvExC5MzO8Tbd9z6svEJ6YqdeFopB1lSEZsmLc6UXzerKbY7gChsBG50
5kVswfGY/V3GFw8EvGmKCR5bByJ/T5y0siwNwLaYySpi9oU0lzzjhWKF9u9cny7r
alY6GLsse2iHONH4pUqkEcpV8A2XWAcFac2ARTgmz3svf2HIYYOQZDRUOpUwxlli
91PxtQzr1m7TFDcmHpR942HENJ2CKP5XC/2v851DpE+HA4NDjnjjx+mCdcptrKnJ
EC1BHlUvT22EFWB3zDopQj4UiWDINGsD+VCn1R73I+YQM3tplSjtTPj+SP8+9QIo
AFbCNRCEQpkkYe93o9r/D6P0yzAqvM9/bXUtLDKAvygxjQjiVRZOsdSUmYkB6pux
bUzZ8i1O7vSVvVv0sN5QQB9Fq34c7lWlTi6b753oGbbfPUbxl5w9WKY3krDx6H8H
1o3cghAJ0IWD5BGt/U59uKN3L27jdBSZJFKQ9yMqqTy0lsWEoMiE337mGZITlXPg
DAG/5+i8+zCWkhue7qWQ8dJn+5kDY16tr7Ow+zOk8x0EzWPzDuJ8jUp0XCEcH75d
dduOROzL4wdRFNCzTGpI8CnOxH4igssXiwgtLQxKGQkoRFpT+xoBsVEBbwdEpx31
7RK8xHECC3PrLdxUz67O7b46GDBU7LtNx4WiBHTpZYod2Lr6pwiThQFpwWWjRoVU
u8DWk9YMHwtl7LG3MdluQQJfmGMeDXQ2PrFwgZVcMak638h0tdwz3XYzRVnSHd6F
oiiRcmds/ve8Idh/1HOFpzez1NXKSCOsz3s5f/2JCEFOHygJpM1zStnK2NF0tIFA
BdW1a5+sMpdX+Cw1qa619SS6YD3c/8XMDWqmZOb+ywtuo+pG/VabZOQEfcBOUHGu
b17khz/kvlvCAJAt9rL2Cq6E7sqVHTjPVwXbmCPR8MEPepS1NVxkDhYX+wTIp3AR
BCtu5WH800+xM2uApUH3sSrjMwVFtk0FJ+TRaLw6kWeNjmDMlDxZcY4daHcDlDI0
AbO79QxpEqGXiDb3ZhWQj5BUB3BH1u44wKhcpnJqANC9dkUK63xR8l3f6gyjLHB4
8N2qH71gTbC+6yHgU2y2+xZa6lsuILL66fNJzgrapq12iyr40t7fqjxCoNqaTqze
Et4SJSdcY4UIbX1dRdmB4+3rSLyYLctp1H95MfwvK5wlstA9QRa1cAt3kuEf780I
obmsVoRtEuJNXUbPwHpFPPDE4x8aJwyKAyDnuBncgj7pXTm+O7nVmJsceW+QCGsb
ETcAXO3tdWud/s4eAw/vSkrfjwz6srZyxK1WkspH3mQ4XyOfsEYmZK7pG8WKXflH
2AMnegFCa+oI95fAHkQuhGgzf1zNp4N7NHZSMAgKJc3Gq1nBk2q43uhu0ofAwk76
CjIqIn3Mb5cnj7BTQz64Tbuiq1Bt3g6G9jVDYaLKdsu5ArvI/52f5QeCA6TKWz/u
jzKY52GjA8YKehvbpTATKYaejV51E26B5D1onXEu/8rYXEA7gXRunsBSJoKUV+m4
Xv3vp0scfKZ5rNezi3qQrJy3uKyh6xq19nNcRo/ugHoq9i6tqGhn9rmaswC2wwmR
Ip8V82we+t/K7g0cqlx3YLfkmapqi9xTVNbDAc7m7QPhQc5Iuf3bFm61CP/0QGKm
SzUO4oopejvkKWAMN4rGTh4qopReriCLlKwdmTBfOCCA5rP6BcQJhQh/XMigBmFV
McwiIFksk61s9MN6gOO2sNYTZOamnzHBW3ew79YoSuHok1amJNL3d5DEtlqdj7Wf
XXP8LoHiBKQjdGQ5+fjY8/+Z9DPW5jl9IqaDsYM5UE+aM+d4Wx8BPw2zQ27K5y6A
vqUeJjs5Fkaql01BRJc+ZQjVk4yJ27bR5IGaonIE9iV1B7ZSNWOXWOocYv/+8ahG
Z2tHmLJH3zw4VnoPxxZSmCkMPxtjUEX+oENSq0HpmcQStwVFBoOAqe0y9uFKwjAD
cDetRkv02sOGRZfUQ6KrQy3VSCSy7ejocCesEMAk8Vv51mvkSh49PijnaMZkieDF
ODR4lEOl86VG/PTLB7zRkyJF7UvusbFE8sWxS6+jV0eem//rvM7mrJKz4cdC86T2
qewWrTun2r8BKlwLS1VgTTPRt2E86//whSlYgMqUiEDTA5Of3vOslx6aZtx2oTgq
M4c/2f+edoxeDJc0W2ZAfCJF+iLX2cyh545BjCCc0Q4QDXuwDMDmzb14O8yfVVE5
e2CTL6uXVonCFz8BhblzJjxosWLyCHe+oCzhm19U1aeNXVjvxKpqCOlCt626b65P
D/skFYMspzkWJKOZpkkj/bYoXcslTKiUDTkFvtxk+tqXzLPk0xn95BOQzExrKzVh
cjGomX3jzcT/NrGiyIFrmkNkFcJGaKyt/aofTOI5P22T07jyUAy/M/jJhacON6HO
KJO1rxtdpYO/ZfhSW0vhIrbkXH12Ar5oO5UBFFH3K+pY5go5BhqNe8mrh/udG52v
CJI8zp9XLgFINEmj2/k/Ln4yp/e+ScVdvYmWPiiolObLT3ZTmOgVCSIMkfCKX5Yn
EYee+A/KDkyQZGk5f4sByfFkz3wDYPUqqNachyJMFO5IN7D8Ri4m3df95Wz9W5Dv
OYIyAMO7CXJsMNle3lzwFvdHoDkdEjLfvHMaHJXQ7I8enjWu0fwoy7aiRRWk1Qwn
K8S991l5UOs4Szg95StGd2yrdXqc2Hx4uAJnMp1/U3teW8eps0mTA+b6W0az3/vD
RyAZkPkZkbdF3iDYbaDQmIJzfIac0tfheHueGv+THxvb/XtQziQuCnvELiSoW4Pw
rUbnKBtWogkx0aSdSvUspy7EjZbqCqPemdVkavv99WXbG6MsgpqrIljHrKF7KKAF
RN5/ALlEl4JvdsxRjtoiV0MOrdOGklt2mIO2gLzMPRK1OR1N0DRtXDTh5vplt9qc
92ArPaTLTTsSLy7D7O4pC3UjZCbgJmaABW6KK6Z38ht83juTuceD/PUxrh3ZuvdV
vWzPAfH+3c3iEwSltY7oOi2eocuP3UdqXXagUxS8jt3NoKXeDpgSiKxElv/aDklB
tQPzR8Xnxoskrelh8NAWTh0c3469fFcDWfhsg4FRtSjKobGbH5JuXdSnJiO5uzRJ
/Z5ZAGS7ho4/QC8y55gC7AR2XATgHNeOqQ7z5qwoeULggTLK3LHSOIFgptg76OrN
kMoooj3xO/4PncOZLfBjr8ZF+1de21LQxjI3HquzMt5Zp7N+l2EXSSYcFrAT6oZp
UoGY/XJGQZ97A0IwGqKKIpdsFQ08xyAimaCZFbtGxxroW87qPA+GTXkFutvjvPaM
BGn8/vXQkN6SXLJTfG2am4mt77t2wtenk/OyV8OBFTsnj/eYTy3BYgSf665dBdSN
iqcgTDZlA02ZTxE73YQyLEVA2DeyqrsRhmyNidRvw4vHLs3rR++v6mUX7SO8ZIfL
4Its+TiE2pqDm+1YYvgvPgj62WDfykOjuEcJ+52I2PhO6ULuxYNUPdbb7Ww0xKwl
IceC/PK7648DzfbtZelivG0Ciwb10UURY5bIeLPFOataJcTsj+r1MmXZFAHA5F4R
QE6O8RcwFwI6Bjlap0B3yb2JSeqJXnkAHBOmPR2H8PTC5Ry+LB2IUWA2Wg4OH162
ZxZVvO1XeeIqZJhlS0C7D7ZxDwWvo9lx/is23PXWc3mceLF2cKTeO1X75xJsLVUQ
GTHo/SyZMOTXusfGImrAoHJ//RHNwaKHP81A2ic8RI1QfecWuztiPhk11XVxlDEa
XtREfZvXlTuOJWQ5w8rDH8ip6lWgOM/nsJa5kJoShsAX+U1wKD68PnoQsGe/Ov3w
3rZ6EpZqmbuldTkkz2gcpp4RYAyPFPV8Aa71FESwUwW7uB7xT+Hfpw9iQIS4XIyK
l5QutaTrh1rngLFx/sjNu08Bkdpcm0nil4/xcrMFM7pzZVNsqh17QWXseN+kgiXq
bvkUh//ml4T4MShJZM4L1IgbUfAstyrLsRpj3Nrvmc1RLFb7iY50x5fnnGxovUgJ
3r41My5w7OxVHtZjjGMJI8axpwn0gcLwR79oPMTiX+owwtT/mEomiiRNQOjJEAdT
7jgg41qfoz8ulDx/dQ5KOIaxvzWiDHdYsV6PlmkGl9JOz/m1CNuF0OaTIv/mmWh7
nP7Kw7AnqobpXuqSP8ViOORmsyZwd7g6l0vZKeCJVXYLCFGkROos45goZMA/b9Nx
9YWf+LUoxl4J0j/ob1pnW33LOQfHKPyWBZtpyygq73CwR9jgyDjP/ID75KhlfhaR
BfD8nkd2Um3jBfGLDQ8meUlWXFGQ/yeOSluhnkOuxCUFr8IS8vzYQ1a5Kb+IIpHh
HHlc7YbEp3/GwlAkZJmrcA6KV5LvGcI2PxDxXgpC5JUfTJp7xHR+4hHLFRzd/490
lsffHDfz4FND5bxEaoNtsn+I3mF7I75JuNDnlzWB/hsP8PWxLlCQ5lHbE4Mj/lsK
dPgYyIhP9KdJ2G7KAz0bbZNMQ64t0VMOZmBNCGybW4juoNBYb4GkNqLx91MKQ7sE
qlF9xZclI1yNLtDoe2Z6T36U9x3s/GGBztzdaNGRxGSUKfoqB3km935zVW93gCmf
qMQCbVo0ul2K3t/Z/dCts+c4OCH8q3w0UJt/AkSjIqKciUQmmHiK2Wp2y7caf4oM
UFImXYeC5zx3mvgMAzve3cSD8A2HW6s9Y+7aZ3GHHGoY8mNFGjEBX9mnJLSN8y6T
nZKxrTA2O2Xg7LYq12C13/WTPqEdxDfA1RIxWkOv6pZ1rQ9sjF6JbbeI461PxOMw
+y5vXnVPk5e4U+hAAXlGLafusC1q1wAL4aJCZ/pgYPG9Ubp33j983gVIqm+rcBk7
aFgScxpEJB1x0Rq0j6Jukyih2S7pRPhzsk+bkDdCGRXdnnfxWo7Ub5MFgAVzo6YX
+K9dfpqnyDtUercVmp+xDtJmWXrADKJisQBWUnHeSZKBSuRXL91474Wpu6kscI0T
s5nxLxyzVCSjrndda602+/Os0xSra8d37Ld76uKAjBgdl8x5V3S4dWdsR2ZrsXvU
rOAv07HzY51q9FXraCJXXBtneeb98/YZznostgc6z47ldKGZZR9GOVpcX/QZGfuT
zr72TeY+OhEpAipoC6QV0vSZQTYLfL50mmDrY0ACU5DnJN+/ExurpGgWu2XmRJcU
xy1MLoN0AixtLJ3dSjF0GHF1oxFBy+Vzq5IG2J+LKlQVrj0UoFSEnO1dZ5swMl+v
rYlUvZwQ7pE2gIoJ8d61KijI9DUxuGC3yMxo/lT9oMQDbnqYOZyuQoOp/iZdzNRz
rhl/JIJUZLUmvXJv1XQ6FMckDv49DLBqYcEwt5u7nNbRB8tCCqAFdG03MEv90qBQ
gg8nNSfSyJ6opPccEMmkMSpSA03p1GG4woyMxSO6CRBQUTLgNVrwVaVPuKnkemt9
Fd2GGxL/udPQnxXi29gP8Vpln1cVtq1ZAWCG8Db0SGnmQQMWcHPJjvCkUs4sOzgL
XrrCSx60hW3I6qLR62o7rREKtfv5isw0fqBPVRs/Aq2QjT4CnQitkSwJGsQdoA3S
IRi+JbWaYRHJZ7BWIyD92KLUhSnVTqMD0Og+QT/fn5fpCfOPVVcVzyS/zROCjID8
LpwFoseZvPLExtz+lLcZw6KWae7ZMBMuKD8vhnQl3nRUiDanzhxoSEghK2TmPnny
ZtduimJ75aNOjqTqJGL5wPmW0c3jMgPfUG6E+2dzcyx18wN4JsPw/jof1+SZwEQq
yddft2EWH6DES8LYclVwFElPqETKeGJKQH2ay7xIAHqpIR8BNc/uGPvfDJF7PON6
5uJyWbDVt9XXCMm3L/RXiizcXt/u1wAJnd3X6pT74/ngiQkb7ZSe3uDk1X/DbLVn
snfPTrHcOIs6gIRhQapbdF1jI9SYXptden+eDKYazrZeBVOFg4GgahkHuqqtAKlk
RjLnPiiXWJgvs+j2vvcS6uqqWlarsWcuJU5WWOUQtusyxKRSHaZWa6//tSYOzlvH
P4J2GCOWOAhBYFVZp6IBz8EaT0vamXC0QNOrJYyODOFsHsdJ2KciJ1mR43rpnmfk
cP9DhomP4WY5y2CeNFnrZLbcfHQ6K1eqEEALj617GGbvrv0YHPKA/Nz5jbCQbdl8
ojydJCkdvBub2iG3d093ZVgVQciJdbhLKTJvrSZfD8i75WuASGWv6MJkoSF94DME
GUPqgl8uXm8xdbshcWPEFMl+j4VoF5w5Y2K1r0rx4GvVv4OQCVBnVuNdZzz+MXO3
uCbsTN3HyGAPivzCsdJGo/E2Pozkysy1uW+zw+YHCwSaLTAUMQTE+Iugk7fsYOW/
pAtdgmRfAPsfD+m5EwzZ5NBgz+XM5NC8BdhHPHjO06DlpmBDWZs2YUyS5ipHNYJE
wISdVVzffL0AfgpochJt/ZiorGTALyjz7SmdDx7DpGK1z7gRuAY2CmyfTXVx7Pq9
XSO+RWS6KUTj1wMYNMR+L6JlmQXCh1auew6E3fJo/ShF/LaFSzX4TNDs3SoHUqy2
TEvHYDCG91CzCCGvEA68kWLTNCULJfP1Dsu4cmEXJqUnzIT1ASYc7/3BhY+twJVC
Y3ZDuyM7CXObceelMZ3lZrm+vBsjqs3pIdP+XiVI+mA2UQLViAyr2Fwvkyts1e2N
Tq4/owG23uhOck4NwqCobGasvwvutYuPzGt2bbMHxIAOtkwElwgyn2Rd0LhCW1EE
0zfqyVUCKexWQ6VcW5GA2F7sitv/JdGmpnvrycEPNo1ioLteuGMFjyV544B9cDCO
SeC/zxvZ9foBb3SEdxyNb90F5E4En5bwnu8Ur3gZGLUSgTt91lqm3YvCme1Jp5fN
oEWawML92pTN/l1ezHJ7Gs2mVtvrEKdw0SBSRc82NIt/38jibkDg/lZkiTxI6+li
dOoge8Rd7j6JmMm8De8C3FMMvNXewCqFXcso7DTxbl24WralzrrLXKFJACmVRx/4
9f1f/qo4R7wjQXIftcYJpbx/kHKhWsLvw4n0YLeElh+nJoxx2JLixRS9Z7VWDCQl
ws7c/tIDulyFUX9r/mlKeAfckIb8C0TugHDZ0KiCKhPZh5AV3xWV0S6asIQkpILW
Ba3W4BAODl3aa67Y2H14QSc47nnK4LxCKv3ceYRg/AAlyIdpzvViUgKw05BuT0Kc
QT1AeEtRoz6SZA2KMjZRDnVc7FMBDnVe8a+m79K0wIFydSynFp+axJ6WvZ/wNzjG
kq66fnpCAPXWznZDyoQAFDwPkhei0ZFFQE3Q/9Jh8KFUtWESYKJGEMEHSFwOQMtU
Hd6pWdQ10hblScEi10SmPXxX3JUPu47pV5/MzqidTjj480EXppf0hfiRJvfaYY7Q
wBL5nWokN+RtnkDeo67VBFH2h9vMBGjo8mAQCRasw3Sg9Es5iSNnyVQf9+yD8il8
+wUbr8MmfY2qpzSp/M+EsDEc2EPyF9zPScBxe9ac8LdbhF8ePp9yQ9dGHPiR6PJv
FjPI8+hCxDRMZ9HdKUlTDR0bg2ELZxJjn6HPAsRfobio/p4CXTo2PZSC2U1Yvih1
ndj5xf3I8RVwAhYQjJbFL6VzJ+AF8pm8rjxwR/oUOOCdAaj7imxTPqhQnaKojHgD
o16lJYTTlwO6PmPrQcgBqZYfM2CjTe8Xa2tgVEnMB6axae1EZfg4kVSbvRMj7uec
I3ru86AmQb5HwwoYqZXT5wPeaQ3hFAJhMhreU3WeBIyTcNyIEP3Y2GBuBWVNOL1H
uAjg3ZPVcIAG850vGkzdnT0W9wdE7qr2RtJDU6pxb1XjjmcP6uYlg+UyoyvNOdSn
u/VJnWSFT7O1CjeQbGT3z4fdH8CsMiv0tSYMMljzd+syfr/KEPqwKw9jPd+tfKnt
UFI7//gHR7rdyPN/vgoG1OuhxFQFqa6tmBEOFds2pg+6dobnfMbvpflnlwv+kOY9
PvasAzImc/M2KdUhyKh7a7poOi7KDOwwnGR5NjpZVZHyDaYZpKRVEA/3YiJgXeKH
VHlkJdxqvEV4JZj82PO1Un4olt0nVPhxPUVTJsIUC9DpyZpMAPRXjGFhLXe4+SFB
35w2c8xVa4kcpl81NP1mCltNTwivUJ7aLBjvR7fI67T56+XS7z/4FeHP0Ls30sfA
LmUXuYMcYvd+UfHamfku/E79o1QJ/tYjjuDPTe1cNoQBKGIzkgqF81d2XF3AmQIF
EAfFEsMGFnzg+gGfLJ91uwiqvr0kTCWVkQWcYdnScNi+zFezrZLgiN/w2JuQV7s4
8DiU+XijwZvpCDTXL6fJpbpkr7PkQSAZ3I5i/1o7SLbumji2WYeZO9vFXXstLDG4
Ur0JfTpXos5JFT91vqYyzcGzH1rgoHXGpPz1WvObagHsQb7V9pj8EbpynczUmkBb
OP+yKGhbz6D9SQdAyfxr9tbSkwUI+EXYSOm5rsVVdOuI8KFuXd9ZeVxKIbIAbTV4
3SG+j4k/DYGdpDqpH+LZNZm97s2nhtJppHTRHQ+9SXM4QQSPmIPLIrdGXQDhRsoH
93oQoPvq4LUfwKcSZsGGmOqG3HNAquy3OSpqCjy3GpNgcb4sU4AzGcxnFQIRKQSF
71nxaO1AuCR0q4VN5UggU485N9Eb66CQfxvAgjv8Rzq7yceqRLO/2dnsZQ74CrX+
abiwtsFHGZQN9N6fCzCKqWnnzQe+cg+DRCnFELa3BoPxTg99LEhP+I0Xgw00PxAs
astUFSZQKc7bNLWwkuAnFYT7wPvWZZ3ceGxsBXF9+P2R9wFKrayOMIi8u49ktcWF
UAjqIJqBo/ssmn+epozIS+LUOhhJbqmqnVpJfPGRAp4Zl+/XHQtQWgCtpMPqPZkI
KxvxqBgG0UdTOSDV5Vn1b8GRkEsyw/GXDhR9YSZKiv3A4uGitbEnMehF2S7IohI/
BA5xomB5L/678oFVzJJ2GL/EcuoGs0JUmRTd6nvj9iXxDRcwbpyjm9CwBgNO7cU3
dshDCw6BI77Jg2v18gj114bduvdQvZ4VGC1kEqW9VNu2WgmQXkXANGHGmWJEE6tZ
4KA7bm/vrc8yCjUHfvBK5cH6JIo/pNd2FzxFYaMnRRFsjJvMJ6CgIie607IYPbU0
y0JnxXQp5HptU0uaPyUiPq/gU0o2qBnQf6yBVP5Cb/6plBFAY6eWXmRlsnTCTk5Z
SyRh1S0pm5LZMr3RYB4Xp/V41Kq6JvMRo7nnOvLCeEdeOkJrDR7DkhN11zRqPLCC
o47+rvhDnw64L1sotil6PpWOgRTsw2EAZ1DYuCHL8JC/eQ3GonaZWpNJl4bCbQta
hFgDuVGZzYSc13dW2/hE3hD10AQu0YULqpcuVc+GGfrYh17uyPM+W9hdAn35AAoD
uA8Do/e3hC31OAc54XLxp6f78WFWQnYiMyYeoacZYF+WBcm8HjSxXxmQaJ8TecTn
daf8VLYg9bbCDOtFTiOccVHJ8c+RdEorsnHMZ0g8OE4yBbLnN7Gx+4fTaY+3zC4I
wHYG5BiwdcK83/OACB4tBpB0/QiENLWKxesLUMVJtXw3qiWKoj3H7KssPfuCzhjx
NHzQ43JT1dTegn3Ozd1EWVRR9zEOeB81PzpkdPaxapCw3DDncFBmqAwjr81TD5dy
GV1mzCB3tL02sM62xtqaFLEcUfW1rDnZLwjTc+cZ8nrbrObOFfY8CGdAGAipo/Lg
O1ku7dzxmAj6u0pyxiGEE2YhId3Sc9ElZQVp+fwh1s5/sMgq2mcMl/Ax3QeZtpr3
cALjn6v2U+QTZN70nJBOQoXdU7cYZrqPhNbC+YkE3g4H7S26N663y9Nh7hZf6eGS
XFJL4Q3ufL41ZNpbShqpBEsbp68/ZOK8IjFsnVGn39m+aQNL9bJ8+eO29alfv967
PW/SXC/PkAQMHH+aN/DOpsy5pj8VD1bXN1qe1KrtSrqX97eUqJydG6xSpJ4h1uTm
VqcsAcaPW94Vhhv0UegSdrhQ757mfKx6UsO4mVlGJAtQdgtEKRDCgJbgy1NZFYw4
kLVA9rp1sVwMME/QECc2/YMwuIKemS+I6RKksXcIcB8sGvLOenvpPXD7776j4N53
RW5tMUFjo7aqjodCQWK2lLujo5FgqnCQDg/zwFtb9jFkTrsEMuORLNm7U9ukABe6
lcEeMgpBYztUnBVaGbEdsi2cCuhgpJ9WJhCU3Nk4Kb/d1ujIlCo56NUcuamYsnhs
IUVSzz9IjEz/e73/GkJEVYi7Yza/eBaOF8lwx2qAJRlCABS2KBf0ksL3Bq9atii3
GSjykCAnzQ3A+LnKtWRrwp8O/EcD/H8IAFT7eEU2H+lCa/58VnOp5nl9K42D4Sbh
7XE931lqgAR8PNnNLmgawfWoUaLgOA1PgU+sOHtiUb9T5Wb/zGxrMm9P5bc9apb8
RVr0St68Jqf8dKVqeCABWIbzzdHuBgtIB0Ui6b9fBxczbCTT5n7RWD9SZXkhjLlW
HG5xynUIAfXcctOjQMROlCBuqQS96n2MiOygYvBK/dHBps1lydRD8yQhlZZnOt33
KfnhrjXQav0uxBcRIqdeFwebnh9WBfR9L32TspqEu4R8qUpwKoRVwne8Y0HyegWo
3bxz2lkhyVM3W8KKlM5VZzdY5sQRPQaHEZL7oksdUflzHYYaIRnAQcL6Hdj7s9ga
ZJpTheKP1Z6D+zpUlSI/yo6V4bBrdzMol+sivqUVQr+iEhmDN5XnMnEoChdoOMuM
srTovuS3v4IYvCB4zLik8bE3WxOVvJJyvcBQly51EHOqVPxzf3c2tNiDoan3ztzM
K7UipdmzVCiM2cYN8ic4oTf3jIly4Mkm2CY0jhhSuwyxh4Fbk0+gXC4WpPVhLm9V
ll4kBggDdonp4YDt+0G+ANoGE8y4W5WESfzWgJQIwPfQyjuwYy18CY8TedPZD8W6
hADQ+ewo1bkW6EtPjXjUu/AoQRb2D1oEmcosFMkUx+TgsgSEuTDVtz4dUokECloF
m2NhWy01rgOguMFWhrd3ld6/Y++NbxynWclcSVRLQFIPSHiykpCGYy7a7EhYQGGO
zwVNJLso2nd1WLdDmJ146y/5DJFbSJW4BnlHTvvZoB1nbBBrqdLaOUTSVOwQbNw0
hUh2FgNkhsakxuVL6kQ0HrWiN/Yj9iXKkiaqovixJsxpztNKtCVOYdzPCwZa/T2D
wsNeWQb0kn/OXK4+mcYRDnM/bZD22J41AmbjSwpWpJJe+BTlVP3WhQyXKqNaKRQA
5CM/X6vc5B1Qk34hnhVwJyTUmc1nSwe5LXfK7G493m1VrNppSkKV5zFl8Yv2oDAD
CT2WZZNVHqXuAMHg4UeyBEfQoXh33A8S/M1TLsiV+g1+ocz5uftfwpoKE4yfZEcy
RZY//NSStSMxT5VMK4wZfju+BYAXTHRG4McUU93hG7jzLhOnbsNKR1g9OZKZFk/D
o65Y3MUzEZ6hvcbX60JnVOiyUhHZrYVwOUdTZfneupi1ntSE5NU2su2kitVCNovx
/kYvg6jNmABA5bNkmKUFK55khQoJGABw+im7oyHmDa7lsB97KCzmDGLh9b2oMsqt
ItIzu8LwfKoTQD5dyczUDT5QiFIhxKM8mVUS2RIelNnUpzvl3QCmZQbn2hnwaEP3
7pBoGVUdI2eXTvT0vtHbPf9DRGF8h8NVUfAgzIyviFw4OHi8d5t/NI9MB/GJPTuT
CMX7x/lDCrxJPVlvhmLsR/7R7hQCf3uSydFefPGGjl9pXKpRurwUZ73MKHt/6A7C
JqfcMuVFJJscwBMS2ZDmNMynmL+8d+lvv5DKJqIGpEFxXF+OV7+mJ1VmxMEmTFiz
296DqzdXJDzc6yYZDPzqca4C31tjIcWMpRn6p3Ozoz0gDRYD/CBCLVbFP4THvzFa
MJmUUznVTR6JTzb7Y5aQN+vm6xrRR0pLqoj+EQKfXHXphSbP9z4yJYl/CV25Jq3I
clSFmUpZIrtag88lWGLnwmbtui9vEzWzQIhifDRHXM0CZ/q1TU6KzoBGIEitGm2i
HPoCbYxlIzAThxasdRJPQgKVFukxsfyxBiFzj9tKEv9qWCsUybQuz+wBh7EULz5S
748YLlerGBef5n9AhFjbwIR7cfllUxN6jsoSmgPI+ozrPJ0GwnckAekdyuem9Z96
oJ4PlGdyVqLub2PC+qm0wnwtuXCn9/GivAGefL4RWm61JYLP2/teLmithXU4D1QN
CKnN/zAGSDQDUrXC33HZ5iDke4KNgJr6Ofy0GOiDRy2VmcV4qboVCTuAiD0ocSVh
wUc+/crbY/0Mq6duJwkXam17eNg5dFhwc9gZwRDCb3RSrNZRdqL6l/zvB8WnRlRK
XrSpK6L92MAO80mqidYaTpu3SJp9Oa/OmmTKXCaaRgi1B8i7ZflzHIkplZ/mS4Bq
BXANCOD3zQGP3BFt0v0goYTAreitN6FylWNiPXcFUYiuRGac67qyw/wxNXT0bxan
pupC0mkIQE71TktzInR2K9mEplvy4pxkvqlkKG6gMFD5cLYQyvdAsEUZrLebZqun
Yfv9I5TMC2yNS7AqaN86RLAjFjPXjHGgTr6GZR9h8L00W4/BR+XEj8eEs7NqhBKF
HuL0rs+YPx0g9SElk/Cag+QwQ6nzuX8SYZWE7kmBfwTveVd1e52Cv25i63wmUIkq
+xRbdNMI7FKqaaVUfMy05A/eqSpyJZlbYb9BVSA38WIcw0fJwLIdRHddPLwu63io
SbsZJOKIYRiUKmRjYE+vc6ZEXZI7cKs9SZB+U9AQvJQ5E7D0kgSAYqGQuOGwcTsZ
mtdY7cedx7PpLEXV0xIqZHeURa4d3HUeS4LR+nGKIlgLSiFrVfP5svBhX1XM/9/6
h5oMS422M1M5wK5mXP8XROKwFOtkAOiSf8B9lujOTUZnw7psTI84wXrAYtSzokSq
SYbQQLSAVkikA45MXaRT2VJMwXGe3fna8tkmHHxdZ83DeXZilqVW9cC4u+KEKJHR
6cLdBRwAYTvW/jggrGzezOnnuV5Hpg2Vo/kcagpiGda3kS1YjrgCNZCDkn/kGzG1
bqz2QOESiVr1eOUN85VrOWfzi/dJXNmWfbR02gw17fDyjf06yPxrvvb6LiB6LooE
IrXuYBL67vzEUWQLYA78iCX9S/SJMcUHioa7LEyc++ReCHzmA6/NAW4AwDMuAXOS
rvrRqturqv44rsv5FX1PKr17iYN8yF9pekeVT5YonAsKKdlK08TAOcIM2IOwzLox
0ocp8TPdCr5PtFt/1PXSz1ZDKc24rUqJSxQ6Ou4nA1GtEs/5BnlhpqgJjT+EKuDI
xf+U3+hRNtY3s3mfr0DKCuU7Ue+lAvf9MNWhFjDp4OByy9ueJK6wiqbkIZ2uX1dV
PdFheRjaP3MPmAhKtPztgVelZ4FmBKr5jmaTcIBWAXFpTMm5fjzMnBa9hBkj9rAC
CTzhdtEOnEIROKo4dPJHYIcXmhWcU9va4JXVj3wlK83m8yKNIeTqObAjnypj6DA0
g6pbErK+PKsgCBp4+IF/mAemoFOiExnJmRcB4Nr7KcZ75khrUSoJDxfpZaQAo3D/
t4ErIesByCvpIHJAbQyMGXDAGrMPAa5B5Zxon4iL6qmDEPRtDyNrfVPdmii7TU2H
j/lQ7ji4Qcbx7pqnpGHTPnum2Boj+b7eMevvI25SUnCk+lTh6OhtMe/XJbyn0d2V
mOAGx5lSZV6YPeP0s9K39mDnKRUjntAIb+i2EqHhqHzuapEenLliGNfD59ZvKEK9
G8uU3HZDv5VD2lP57Txe98kpjuDOcQYRcoyUFuy5ejBa0Bom7Vy2I3mmmJ57uaF3
eUapWCx9Yh9u+97yZaufhAfyA0evlFdWrkY8WjnnmZl85MGree/0TRylBMJX2M3y
Y+XwVTMfeu0i/sXbdikH7hu9SWGkwFNeZbOz05ZECgTvovqxDjz8zWe3d26IxJai
bQ7HKmsfP3S5dYvXfe4/oXrBu/y52YZTEmAFkHT4iUXKskebyPbYnb6onOpLT0cX
honmiYGbaS8asolqbeYJWvvo/MbQBvRQB/R40k0sj1e3s0ENGlbI8Z1nhzrAdpHj
AkCIXUzNakFK55ozJ1SjSg1XredAQ/UA/PtdK4RpseXgXkmqDp1hslYDW0Sw6UVK
7JA2K5SotbAGVpzxzmijfyuz3IjpPDcsVkB5UUHdPfi1BJTxwUGVfn67hcxdMcjx
ZyyG2soXkiAVQVoeCs+wqFdOIh9RoxDkDb3gPvSQpmortoa0SZAGZoS15BPU4BI4
B3nLyvKf4VVRS2YrHRerK7/CALQX6tDqZYj63Zsw06L4IP8vjefjCPJ26/Cels//
6u21/kJPzNZx5PPLTmKN5YnWQtyh3mBE2dA/BOS8fDzzPHL7T7OIlhmqWMMU0/xc
HjlbiCXvFEvotw4jMsLi5A8qOukDu5AXxh6nGSwfQsa2i/E5m7AccDWZBv+2KdvM
EXCGlFovGDH60pwvZKX00iq1izSKTnwmmzKo27PZlSq4hRvEiMsxwauWhjAObpBW
mkR8KaMRef7amzH3IwYRKAnVxiJI6Qm2PijN7YfjDhlNUoCAhQrLSjsb5wqTsazI
tG39m8uR3fIOEMlJET8ziFWqYtrVz6G0SH/jxLyukO2/AoU1kITH9MqQntRBcBQV
sK33A97jm3bfStAhD7d4GKOMoOY12MnZsTy60RUo9hhFgdf9Z+8X0VDa8fGUVrMA
ISiqNeLhcWXtsF0FBzSwp7BcMxtv6yMUUFc+poXj4fyIGu4WIHNHXEPXPlNWfuW4
nenTpJYqNuqFkuHn+7uTvU+CFFPuWtkq+KXecyudcih21zTgxMQ4FcR2xBVJ7OAl
qep9TlQB+6r+2ecXybPPEVGOaT1RD+3m6iIwjtzZhc4DIhzhNI/4QUiMp42DxTHu
IMnqYfL1QIPY4/IANiu9IxrfnQRpk96Xb18t8jB/uvGl7NrvwMoWy6hmli7xz0dV
+ZAzOlKLnINcUyXaM2fY6wxE3TNUcc2UcJyWltsYnKaMhwrSInmfVHFDUYc/K0xk
zwpHe6EtMZlAlZH1TaPslWUMqV1aNSEXq7gSopOxipc2maABs7OJ8IKFkH5XzXQY
1WzvAeGe/HTI/y2LPrA9z6xjuYUO1eLkf4UL7smepi1glVYH6Q/Ta2R1Rc4HlH4p
IVYnxMCRFNvo7XsR4TA4oUA6Oo8DFkYgslHjrrML04x7wMyEkgeDXfy/T8t2LsQZ
U86fsq/ylrDKtBq5aPSfz+SgKI+Blkk9aYMKGXQIehmiYAh411Y+yrgRgmvNhntZ
1Yla1wOU26rLXyvwiqiZ85W6vCUZLktaRLtSTy1wlT6EpTBXk/Q01c2CQ8lEDvB1
C4hAr8A/YKLCMl6I5L9YoJOCMdPHNQ6+xkWzgqeLSTwYcudXA6HHTyHMK/z10GF3
dztunTBtyhmwZz7d4AS5/7iHKEXhSdIw7i/PeWUy94FIQFbuXkK8nD+slgQHi/co
lWmLMBOlxUZxBL1bompjIf3KA2HQq0X2sAw7NjNFPXH0sGeEqmZ2RWlFYQZzLptp
BMIILv9E0EgoxrVgB/g6A+P8jBLQgQxAvtN0JV8vxzj/B7WGaOqdXeTlzJEWEfxA
+KclqLXe75ySHDEkMHbJsWCwlSj/h9o9yusVkdmdIfXgd9bDazupLdxQ9ycYqlKg
SynSzdheBqQqJiUkpsnEdNDmRB+wGqXzHyl3ckfIuWb9n42oYV/6YdVwX/9GD7YN
84fnjqWZ5dUci5N361BdDk8rn4xkK1QBBNN7sedIKArGyzhzasiAl301T2HEUZfb
AHFo8E3zVfD9b3I0lO8zKk+FYyJ0iA2Kz7/VFa0X3vKxz9RxEXuQbkApDokLC5pi
hcKVbiZHICpgIvLTA/z0+yIoEd0xAYa+W3wMppu4GjGbxjeRbOjs0L834QpKrU8a
i5QYZ2LSKUO1OxdbH1wOb5i5EYDpEr/89fVkCuvvwmPu8zV5Cb1Zcw73JtBqnVoh
+IX7zqiKHsc9u+j2t9doNEYOEQLWDMceFo5EbBD1VCNdsdeXQgh3GvMhF3IlJGcq
4XQEjWvRTqfbFPFjk7cruBTzhaPC0NkHwWIBkZSusoLsbxROh0ukIXvJ9Cn9HeFz
5PKKnp6M/JaP4/R72aYiPbOmpiJYUOIL6EP0dG9RZhbI79UjwbBgC5TqUH0xRK3O
8fT4ZdjMf+RloGxZcFf7H7v/IGW03V684DDKlYTK0JVK0NgFrXYcv8Yrq2kzosPx
j+JCv+9cCdlFwmgEfREtenUgKicmyvK8vnDINYnojNtLkAyLsERJ2nrONGYT2ZL7
7P6Rp2VhifZvta+bnK4B83gwa3ciJfI3zXFa6f8wg8wChNelDepfMRSr4NzpH+XT
XOUJsQr9i2ZG6PxIIZkstG98+kZ6FggDnhwyVdeLj6nXf3y5mIKsCBgB9QIOOqfa
Gd29ASeraKqjFtIpoCoOkD9I5AOD99eUwNmFKjug0QdB9JqTmbt7ER44c9a7ouqs
1jj1JHf4VuwOvYJw+qSEnx1h3DButa/Zs4ZpLNcS8ilq9QREEP10OEFuqibek4ys
xWIH8lz4K4zljJp3LVcGe+KYrfga7Sahg1DXP1mxtl51UApOFkMnUahsP/6xPK8Z
hmkvd+8drD65XrbCGQarupeY7ELQicimxCCi4rJ85du1ionYEyXxC3f8zwVjyHsJ
uZXzRB8zb8j0TWq8tKILxzc7Ov94pTWtFnoTLkvg+5AD6QDgsJQfZvAMS3wtpZBp
1uQwilcuaRc2VzX8wMMEow+Yx4aVDrj+o2tStR74DOsY/j3zturTQlg71MOOiKt1
4JGkUnbJsb9V1TbrnPxV5ampIy422rl4TZk7kPXKAZ2XHp9onXT8vRa7mAGv3U3p
sl8gCd7age+5DB/MfRLTGSJV7NljP45MqPQ7FqMkchMG9yyiGjzkBiErmVuHopgk
AkpjSQIJJjgqtKKxYn1I7GcDX6RnIFEl25Dsll+6T46oDAN/oaqZ2RQKxIyCfopf
IsGNRV+asFhOzyBDFZ/9mzMb1JyJHFZDxRFa7rut6GdUJywaTrGNIz9ZkLbEK7Xb
US4N8zi54Dh6GZ9E/wULlvj7VswTtNHg+voXnEFyHxo1Bf2fgkD46uXHjSwre5xv
G794LHiJ1Q5MrRb6KHx5u/cys92bv8OA8ewZW2ohp/xRnhPAjkpEghUHqYF+AXKL
5jh3vWENXIpavuWzCkywGM8tKT0k5Lecd9nOoQA7kWQnfZAy7AR3pCbVDvS82agU
qjd9bFs+eKjT3KWiSXSt3WMn5Wy+NRBJU8uqpjbsI+KJg/HXiykZF1PEGw4ScrhY
lu+CGSMHV6vf2/eS+iGQwkLNR1iTLKePaMpkworeRZq73fotPFcuAYugEbQfFSYI
V/jb4qWUZiAi/BW2rwWDYsAy+ndorR022xTUYNVVxZFi7PasHW6rAvg8LB2bD0Vv
QPgAZ9WO5mdtyl/D08a/P62OhjuiBR+WrosQV7kgNlx9f4MxW1ExdZ4j2Yx8i/4y
l1VTgoGWPg+9ALYVtfH/K6U3685/cZFrM+7nrrhgVpcNEzBtS8z7HVEneg5xVRok
Bzz+be9yYfskvrhGDGBTCoB3UFb8YeAfkwCxwqjOhs+cEiPu3sNPQFj0A6w4alcE
7VLLhXJXvR2sMKMIrJHsZVKjzAbk2tHeu6MQ5StoL18PlFWz0TvZLSxq0LCQvk06
HZvEaxXgzCsewSmUtltXNjzAzCiUyG8RxkUAVbDl6lhvJNYEob2IROikoDnO7mm6
c88hjvXBD2LMKh2lPzY93AioJLPDW+6kgkao44rPFTwvYw7AimMTH0cRJbOMOdNc
hEQKPg8OURWy48Ym7nPlw7+XPy4AkamuJnCVo0JXtLdwG8liYXr0XO6pGnyNJWLn
3hBYvp+2zuOb0pGQV+EdTZBZEnSZ9OmvPWfp8RjWd6BoxDAA6Tmc0AgQ5ra+qrHF
KA5Z0wfogFYTw7IYNEogQvIujJrLNwsrLmMVOSMr7fFJ5ppTZbKhFyWASDiKu6t4
/nEGOxX52oHnz9rs8BU3p4zYrRCerLADEEIByq/F03qKHPKq15kqnCsK05+BhjiZ
J6PtDkwuVg0N7F+ncTO/NzwUbIGI4r8NL+Sh7R1PAkJMCEdRZmIul4EQhl3BHA7Z
rnEtMemnTWD6YtB7fWFZ7msyJmrs2eEW45xMzguUSLU+7wzwGXkycW3d9b7h3v/U
VqT3iQE28t+Sh2CHg1vOxBBt1C48GjGbj961LBO6iA+mu/xJtqB3rmvRdUAFL7qB
fo8Z0TRG+krQoJNNqT0qseAD53XOEzpt6lGmdQuD2Nhf6yNRzfDb20/Vsji1+t3u
oV1IXqyKay3hOeUxWzDxr7NAVDK1NZKSrNNpEG/sZPTNdXU7n86+x38r/lac8x5O
XwEmJw3mK8nhNLwDq+YarFHDvIRgMGMxQ/cOUPN0pHdOVS69KK0oI9o5s0P/5wCJ
ogjHe1YvLnqBsuodrOGx3+gIWqXP61qXy5UtloJMmVjm4GyMzoM1KjX16AFKUVuV
s/2wMHYu4YSgug+c1SFuU7W/nwdlstYHwYRTrYpkVeYE7cfLjTtnUkjNUVDbsZTQ
rTz2VUYMfSbP2pGSBmNWGziWRDCjQPzCUECDoL4BgNk3SpGxwiXpiSIYZtXyLnAI
h5sWwdwERPM++wdarXB0D8ryhZU3B98lWR33VSUgboZTYvb++OuVHkNxiBf8SR/I
jbB0d7yBwmpRZGQqLobxqHSGNqovNRW4BgzsTrtyL393cne+THRDtGCcp7vVT2rL
bs6QgGyS8psTq2iMDnndII00aB67Ebyb3d6P3g/gUyPzzbRgrGQcfF57fbRK6rsA
P3C6jDPMupi24+2SdLlSNiNXoB3sw4/nePJ4szh5K/ubikLKd9Kni2ERYT9PgPPf
6P2hRTZQx/AiYsIolNP7HsllsuumcI/Tv9dLD69MvmQllbvNBiCLVUrNdM7ugKhC
SCoKcHMIluLP+826JSWj18+5RecR+K5Xwmt84N/3dgP7Qre0UmX486zeCZ1P+CJv
Spj/RYLFF8floVXups5C3RXrc5Z02NVqqMfOGnnAg1M/2Occ3r8xaYOw8DFYtKqL
h3sj5mxlAOvfy/kJJ6CxJOgUXc9tXibxtX6TOhg60Hj8s5BF5aJEQuoT4c6W8iui
EI+X1LQfSEwQkMCDa/JiSMRmnZ5USNWBnWFVDQLAjJ6yOj+V/jVo3yXy287c0Hcj
IU+13nW468eCi4usueyiudgADFZTASLkWmL57OMUJZh3XaGFdTo/3vArSuddGEEt
zVdL25Xw+sT5OZwy80Qf8TSIju1BI20IhZ6zyxn7Ag2xRbASlyyY/4AdpKb2rHR6
D8cWKkVj+4VQLiBNASqE9HH9PdXd6XuVwfUoBqacVfmkW27d5TwwWzvYBhreBHWO
MGOTnL2lw95osWHRREP/yZwsaCE4ityrdFjDrMqz8+lJI3ZGUtbYEKYytHy4JoML
I3lm0H2G9PnbZPvUKUgmlxWtXLdrL2Oiw8/ktVx+sPpLpC9QpaxjTdzkY4MqztUe
JUi3aJHN4DiXphMUIyo8dSzTQoCu0EAo0okrMH+K2oitxuIcFimYAEAiGA9MN8OI
kPTNDKZufnd1BMlPaXAYFUK28BBJ4Z0X202Od7CQoc8B92awN30Uhb49r4tnodbB
Jorgy6vZoC7dMMcxhUDPR2EMIvyJzo8Qwh9EJHQ9XO3fEYRmceAGmBhPIZc5hf8d
y2q67ivzE5HdBZo8yACuQmDQs02Ogb2LwXp9+83S7+4xAQPFwwvkFO053Jv3bP9e
8RDedhQfjPcyhz57GMpc2f/zBGf2KEQbVbQ51QfVtxBySR92Q6uga/zp9XpeERDd
ORjl4H1Wrkc0a1Rbh+EOtpJEqecGdxtWm4pISrvWdq2786f51jLMNZzHRidRWQ2/
BzuDiswmXmToZzBlZ1qcctN2udJNRzXjWN/T2T+L1J+F5E2xt0XEXXvL26gbT1Qu
tmvl1Iv40k7tLgMLpk0tB7pL5ZXMcaVzFrjKcEpIC/h6RdeI7Iy9Za/5CXgoaH8G
B7VIlIcE4eVR1P9Bg0v+Vo820Ma9dVy2YX/+ME0rSg/dUME45cjRVYUdHsLDsfDn
5RthNq41d2GHcbczvYwWcnmAs8s47bE/xDLLCh5LABPrkwjsvdI8tE19nTBpeosc
bKTfIlHhEj8Oors30/Eb+KN7rFIv7YcZ2mBxuW72lpicjHUIzBIZ7AX7wZgDYvET
eipDcrdBespfieC5r1XmPHmIsa0i3rVCiyzqsSFEwQoeQ5oVA0lm60We5ny4axvJ
WH4gDHWC/dthtMlqGJtwG2O/15atyVuv0jTOxMMB0zhNoDUTfkbWGzqfSm2IyPmT
eVaGChdjQE919zWGAE3G2l6J8WWzwY3TI+nNulD5ZqaLpw/p4GK2H4fIpxg8H3Or
tgd26wI6tmao9U/2rEho7cDCLCPCPbMKnl86wifm39+Xqw8LzG+lKAqPpZLfS+7u
y+ZZCkwXX9SRmpfv5UAJEkZ1wAO8b5IPDiaECmbriGwaaRqpqzLZYxSx3dk/eNQA
5ni2hVFVnM1Nc4gUp8C2YqFHwF0i3lSfpKmT5xceyUJIRuLo1yPGBop9DO7tHp/B
gZMUOiCnm2TXYhyxev0WRcNUholLZTd9AzwqPwwjqMRueLp3bSqsQnOh/W23Ong1
GrFyMncljnfoMXxX5hYjiSIjvjgIECFRkBsKpX9lRIgf35OU7YYOTxEiszzltU5r
AicxD8+t1fhPNPxTMXQHPPmNRJPD5yQCsJyDXsiAYBnPOY4G/lvmGZAGpI7DzivH
Y1kukAOjeNmdjSjQiyE0l5jhBo3BIkGDfZik0rGfsZh3KTk6YPkH91khBJWEfcTV
crNPCJ7O3ppno4YFjXDsd74o/l3eav9ygB0T8m3qzKE/1aUvOEOnbcPDN9UYUL8s
IufDtorFbKR5FN/vqmd8vf5tC8Oi129LQvcw4x3kwWFh8Y5DzGw4T5YrUlPM+2Qd
OBWbMX7Ry+zoxY+y47pYqLsaUV88gLcjp/jPn7zk/lfWHKI2RdAfVUWceOscSkIq
F7n3WGgjcH96xj5Dn2qlvNevKlQRaUFRMPGYiUxYVz+nUoXx64ZSPgxZjZJxLa/S
XtqI7B8rjQYXiaOAnqr53JM9acctO60wcz8hKNn4VueHLU9czE03xJUR+GNajqj7
Q5tkRI91i6perPWQy3VkItsis9auLah+Dxrd9X5Nd+dsW5HXjOZ9snBgSguZK06t
1G410INYxX7HlWF62wy4cTlKwH5jV8WJEhz9VrHQdLU5Il+v1kBlEppPDfy1PBUb
MnMj1qunigtNDfuDnOh4lbVN3b+X7zX239gk/UPBjtjdjt3nueh8IwjxIk2zW13S
pS7df1exr6DeeT3R86PBpUEyOreTuLgIKWXMFzNOxSWOIuBx0O4AnvgHzfiqwupF
ZMuk6nGoKVkOX1B+1o60tLmazI9o1sedq//MbLVTBMcv99xsxexl+7xEJZLgDR4H
TXNedleZK2iYpRl9RYfwQS1qa3ZwrGVTsPfVwiRwgTi2RnBDnmnFtYwwxi+BPZer
IGAnK+GQEZceR5sXbF32cY2dggfbKIBPekpHOZIT8BXiLUpYYFpKHFnk+l1611rL
U5oKVgpEbyZKmfb2EEFfVLmFpV2xjYP+rFwW0V595ahqGoWvf6Di0YqWA8GEH4hi
YZpT7kRx2g3TdgZ0uDGHlGQxIAzctYmoeT6VVIunrANGqJdU5Eh3S+bxJ1MthAti
zs6ZPcx6Q7b+pra1zXCopRzEkqWaUBqj0VornKKISlZdWPZOAIszA8NL7kc3MTD/
Yow0BPryIHRSeEk3tp8xhoyiT8PdODFTB8yCR9WBUGaV2LtXRP8htpmOBS4xMzPH
pqplyJeWnYG9/OznclUd7QjREp6rLpffKP3yIKXCtc33rQkb6B2oLXt41uWSLfcj
WgkqdzwAb7mkx9dYkhA/NOWjPuO0v3zuvRTTi7yqAUA7Ch40tzXJRk9j1IoX1CW0
1kLglkFVMQKhW5zdKxBp6X0IkXwH5b1S7fu90aR1FpWwu3aYh+eOHL/x4A7TN4ee
naK/JJYmm4AX9xUqB4bmGeFQVV8mNZOxVYJAiE8lx0l7uY7L/9GWvBNLilPKm8dX
ee+hhjvmSFPdGjjoT+WAeO/Vg5KSm25rZkZsH3v6AEBoCzRJoDuhnLagesiH3ysP
hXOdO2B1/581o0UoTepYcyvur4u0wJ3ohPsLgJ1wMt9qNSHRI4CyXf8MQwde1vMC
3KbHksoPoXQg14fV1cya9G+WyrWLAXXK9JH63xFjKKvp2SOsVysYC5G0c04oL3xR
AsbPfsMsHQVYxgPfIGIlRsOHJPb9b2mzqWPv8qaa18znfDPrFwHxrL8h+Kq66Nom
ZgR7wW2J3kmuWqsb71FkU6MO63pOqtW9Yi9XT9BrcLuJ+4+NhobD/E7r0KWYpsrr
w0kSOvqMF5fTwiwtvA+Yvpgq0aKw897xnuz/oNDIZdXSxk4p5vfhZjfgXk0FqjUT
H+EhEP+DH3VWyS4D6/O0uo7sgLs1moLojTdlQwF5S6ZHcMYWbxY1/3cvzIMwxtLI
g8rooCewsL7nU6tpZsGx0JORNb/kn0PRIAXCecq6WTwoudYZ5/pIV1XACeGgbPmr
CvjwI3TT8VPVLQI1BX2yGWI1zTDxnrpIAgkSG3Iz/pMfMx2RtEOwfoaGtr7olhJ7
Sqi0khwTODNF1r+YT6+JEcPgyQRlGbzrsheQJW4XhejqkPgV+momkyTDOCILczth
Vcb3pHHb3rVF12emtP6lSlSz0b2HTTauwFQ10+pFeGmIPrSa+Ryl0BPsNIynmgFF
zienWdH/2jIUz9EDepl7cA968n8QAMwo5Kq2q+kBxGb3lEGpuy4nhUMJD5Eq0IfY
uMlB6WYCNn9moQpwYXZ0YFgOI2hxYtSM70jkD4ZK37mtnig6bc/4QJZIIkTAjiJt
4+I4b0a4oLrPc5WTt4hSbtMjZBIlqnKgC2FGZB1TUeYzVb063byUJ7Ep1lwvcJJU
SOuCX1F6FjHctTOV7wr4HLVaBdngHr0iIrlsu7serJAswgZaCGar2H2NAL+WPGZh
P96Gw6Wr6/LmMzABWRTmcwkUcfsrNjihzpc/GCIi03HYci+L9OO1aRwEy8XtqBzZ
HT83lqdUm+zw26Y+HqOrJwDdz4LLKDa9d9H7xMLnzbzPzKup/nZab3bfZf1/r4cq
TS7v2RoGDbEbUsoCe7YzfxrT5Fdw8cHwgBqYrLjEHzUKYoijFBcIGLOLAsaLVvhY
bLiUCd+yWac+erMe50JQiasvsdWtyieDxU5KVN+o6pHpP2NIX8oOWMl8GnR8pW7H
JMUV2EYjRpSb+p5MDzgd+0lOrZR+oUVn8uzSHWy6YTXUqDLr0RAAQKmSWiMjDXBJ
IdQMUACuUPprkqP4GnARKGyHupsl/Xe2hqbczK7tmZ+Hggf56ycIejT8IPx25YwO
8NS78fiGZMIuqyvrzcLSdAPCDBaw1B36c6Bjpl5D3+OwbH21FyM0/tygioE/HBhV
jFUGuNaz2kNz9OVbsnmOTtz+RplqUflQ+XGtcVhKOLP1AexWYPVU8bJPPxpE7gm9
rqiq7IcB5Pd5tGBxS/fw1JXlGPU3/4thPy0N3S1+2x6cPLqL19xth3FswYCLwMV2
M7DE9BPFIDPV9g7vx03Jgg/2yNh3txiQk6ySGWgVNj48AdlHRK0IhPSW2orRr0dC
HPNuvuAxB3sDNgw9J18c8iiog2iMFs/Qr7ybda8awxX92405bhVSKMk8XMBkd3lq
SxgthQOVANsHqzqozdHdoQZIZqEAVgQeUbzb4Y1gJ56yuALKewiIQrkj1oRz6nDT
fSiz0g+YPEFBl0LKoTUf0ln+TV31HGoAYs3FG+5d1msmgkw60kgy7Ev+rPdXCe16
krzX6CjYZ2EE0fAj5v3TyNkTVuIM6gR16amdYb6EShXeGDA8uBj58tPL+afp6tsF
z/up52K9TzDNjboUQvYbNXVyFAipcv/aSgewjj1ZgV5iv9kKDNykICVuSB3nylUh
RJ7u84ePz7DW4f+qRGaFMvMj/fyNzay+odT7UK5m30SVizrZn2KS45J1j3M7Pvmn
QiETJrEQD/TDFomw/KXgvYBJOsPZk/kKhAoZwD9JHI7xUvpQJAPZbIhh6BJOWxOP
sAkmAWNA1/93aqS/2y2hQ1X6y7nLbWzkuFptEW5aNWXi1S80xKiA6aEYZE0Sw0oA
7OI8DZdHXhgqm2hg/VinSY3j/+u6mFjPcFiczdDMHL/MX77haSu3RpiedvAc/FTf
3xv64a8TloVKFMfna3FWHnuDCCq7w/wA31lNhJiFT0xsXSHZsyVfhvi4HVpOOKJY
DMxzUyOF+cb8YHs1vg5FiAqMVlvALJpTot40rGiAaADeMrZE3QsV0aoTeSngMy+8
qMVxGmz3oND6wJhIVz7UnB//FEWlxLa+9ITccRJIjeWlUCg85WzJonJXEx9DG4A2
X/PnHOh7/tJlVCpOMA8Ok2blVKEsXug8eRu3pmCXNpN/iuBS848x8UdPG6eQCQtc
v6rA90u7FIaJpyC7XeGPWcLXR9RiXplA/qDQQmnhlYQ3CH5G0iIji4gengJYdSGl
WOrYGg/PUzDrkqqmn/KCkuCQUZvDHAv21sXLob2uFT/2zFdVFYJl7dVAAEsaUJ8e
HNGG4WYQv3MxvT+WNTQAAnbaMnHuPc42Y1MGsK+6x/TCvjhPLobTjhp0F+BQKR6t
8q+Nnyrcz9d8a9fC5bW94q0+aVeAbhj5/0laljcD9+hcO/ceWHUcMSOHYc/ZZnvd
ldnf230u1uvDR3Pi0XkVwmJU4SDwgQWZ+WfUmuip35EBImeKKJc8xMDLiIGYwx5A
AHngsM02PmdWpfnmcwK3Bq9Tu5BXnwCsmktmI+9iZjD5uQDlrbmA1S7PMqm+ACF1
hhih2gDaauXG1F1Kxi5ckAiqln3XRg4omkhF+oBnhjxu09No5aW5R5aqIEid7Cd1
hI5ZvVFJNPkmbdSZpmz4D2jlW8ZN3XaGuRuttjBjZ8ajhcECHUaPZlfklpRgazwD
SOfpHTiFVsSOUBBQk6EkLsuRuDyIDhSYmsBc0EP69WY0IpvkyHykkQKR3tuTbjGb
PLzw/ycaw/At03YKX8/3s/1PRo42Dp/BZyKjoyGqVzE8ogZOh1hg4HXEj6q1uINf
xxawcXmzWrTVBLzOso8ou7Vq/8bcPUOjy2Yrkogssm/7fRAk49twLvhdj1KFgoDH
AbWD1XcEz1RkKF1D0nPvNDVMj8bHz6qJIpRwsM55lu0AKVNJ7LptRWu9vGFEgvW6
pnUw2ellAfv4fTYgUlSTwriVhOe8NH0XWdGzKPccfzM48+hl7rVmFZU4yBaKbuzi
N1ZKZVxM5g6gcu/XyB0J5+qjlosYRnQ+LOOMN8b4mSBa2IVcOrhAvceT0YQUNJHG
Ky0LgP7wz8NIF8aGgPOGgdggmJ8LqEHFNL3LrztN/IbO9yZfwd3RgUpxogdrkzkb
zWMfPt6U57S3RC+hJjsLXwQ+1E7SdNsO+C+S2q8ZYk4ZZ7lINIROvgbYXaXTSPc5
nMoCdTCX2AMQoyQeVq9H3YtUqJO7/STfBVKqcNUnSxUZJrQdB0frZDChwhjHnZCF
opYXA/7do0VChNvkXkGGholerWW+wqwiqfi56T2lyLeEQvyK3gCA2xUrXkzpRjnG
DiV2YZ+C3qEWvZfRmGry/yMHory6VMAhMmZTbgU8RnMEkUBkSEJ4XpRV2pKxdgPg
JxgC5SVddoUvwQbS0MmhyHJLUV4kWu8Z5dGwNzPz2PZMV8CkKYgjg8ctV6DWxIAR
FApxKq6kG6TC6j+rv6wpeA2qxTTSJR2Dnwxdka//2WXXdzSMO7vkm1RCTQn9Ey3f
PdosPzcBDm1CDDEq0GlLnpNL59nsylU0i5urooGEqJtNH7aqVT1m6AiPsqbuCYpL
dByql0m15jxXJLUuEclIWl3HnnxjtXsmGLh6E/7+Fn3IPXUavp+XzVE48oFIC69v
wCbckM0t026qygSSPPSWg804OjSvluDtXdcdaK4sidrW3bybAQHbVBkZ4bF5yY63
8KUCTTm6fvNyoI6ZMubXkZwPOwz+s7tE1QJPQz9qfQZm3tfRq0GK87kTN48K75km
bwpxPnNr2fI+49O1gvLKHVNcnAq76i6NHERzVk3D9jRgV3+LYJ3foWGPaRIirn5+
+/U5Wwj/NqSrCFkQ8TaONB8nNutu5NYEEUYCYQD/++TeesXNSlozLNGtnDA+3IVa
L1eU5tYSKt1Ln2doxrCUpPtD/US/vDej9byRE5MH9Ns8hCAg02ZLIEIb8yGnpuQ0
9FzBr+8u5O/BkhWlEi3r18StJEVB1LfMxi6rpHr/82F8u69pRwDEg7gjVGmnutYi
cNSBoOgpD68itL4eMoD5l5Y0mcbcaXyo6s+6sIEV7omT/VVI0AtJRRPCdWi0YZ06
Af6/S5dGQT0s5iy91nTKJ9ozHCR4PrS+EXOepannKJ1bU7uBPhsYCfDKiviDlzqj
YkW9iqklcGP605Jd48rAIPmE6dhxKlGNCTWMmt0yyDM1/k/Z3cnABeZ0SipF3J96
FSKmzWNB2Rh4y2sDLMu8LzCFF/JnnXiGhvqhIXPNCx6gkw5+IwWk3bh28KFONGId
l9s0JaAUo/x2si7xyAsk+aCLykpMqlJhqtbbAaYdJpLMygr0iC1FX8tc58+C/rjs
2iqlOrDNUq2Soq2Z9facmbXAqq0tt2o+YEvmtJur7e0IIRyOVy3kKx9LUMy8gFuJ
rBu96Dkk9mdt17LQnTwUKK7WKya6C7DE8boCmzX7q4C67rQiY2S0ipuMb/E6SfqP
2jQ3xBr/VIBle8NfP1rmU26FrSP+cxekfCdPOZ4+U9x5jcBnQVYWVZozJX++cSBs
f1sHkPuopBHIVvd+d/7++uYAF7hRJeWw9StW9y51JhcBnfrWxzOaeTJNlrgOI2X0
H8Y695dnjMm/2GrCL7m5rJsrX6snHffIafeB23gmgB1pLoV0ifuy8IglrGmqvyJm
+ZO5brlOlA0opeuVVRE6JiMFILeCszfrW8ASP8+bV9H4PCzED0ph6yrQs3EXb2gP
Hph/xbqLBVVmkqQPT9HHxxU1uPffghNi/ZUnjhTXenH9xM1mMuErsk+r5eZqqFif
JT9kfkG06rTQCtWDoxf41jitDX78CqOKhLoCjJYxLxlEOUZN8EUjMgUM6LveW62n
eALbmryx23xGPgKXFIiVbf2XOnRmAPx789gmlVyf8rfUql1KWf7wS+CzZx0DiJs/
ZjXJglsKzahhZWLLXvKlI7vYRVEOdhxuaRDy/SJUARbYXDjaMYMQtOl4esfJwU/k
hIq1xLtjfk382gWIuTVNmnViMEGLiroBJStwZTB069TJD+9Be52Ra0Fvbq/d30pe
RSUUdKYiULrrgGryVaAqRDXyLJlKqoGFc3LS7NC8vR8zTYKfRtEwAaMIx5XGdRDG
B2vGd2XQMAHt9IoTqbEsDk+xRavisIbaBLw+wjKRSfVlfwz623mJUZEve9E2a3kb
nC1L19JkAjh4pJhXbDgQ3Za0+ArrPA/zA0TuPAdYou7uT8U16HI8Ebauu3GOMAKa
1a9d24fjvwbucUiQYf18Y06hjpeBCVf4YpQwi2luo5EoLH2g6GBUWAKs+FFw5P+L
UBb6HhmjECmeKnao1qN0pmD/ILDAaJtlgoW71v8Z5sDal5DhZ1dLrRIdfFi4Rtz0
Kdpinud0ZN3i3YwqSIi7kdMHJBnOicCseE//8ZITg0Fj6aVVaCL5vmh75shnPenD
nVXuQBejV3MnC+evbMIGow9Ofirnl+tu7ME0o/0XyXUnR6lJU8+XuVYN8rn6w/pK
NR09J4uO2KL8lOs51Js946uUmzg2lIuqDUDTT8i/QgoPHQJ+1w4LbVlr4pqrCVat
bHsjayMaegoHFVzwksV5CRvEgzzd4taRU8c6CuYYV9i/RTKZvXUYf2f1skbDcpjD
wJFY0F3uAhPmI5DRzQrsI0WqkrbTdwETkE/A7k0+DndyVoVYJ+3xOXX+ntUp+Dmy
eT7x7UWlGqsu8CEkVp66buL9MGf8wAXMd8DSg/xu7zBc2L50NVXfuGS5KQYDIxeK
RKrqMUsb8x6PIcsSBq7Os0V2JUbuIOhNTLbVMll2dayuluBuxYxX4LyLFa8qp0l2
Y7dUFqM84ttsasTC6BteLjbjM91hl11x/PXtibmkmVPKDfAP1lfBVPJdHjYFDt7j
OQlwYNJxZM4+MSsiRrVwbWvkFtLtFr6vQw9V7+/+hfno1s9bY1H0LaQT/1GOrzwN
xPPdvYM5TBU2bIdC+rWBtyoys94BkSWZV7V9F6TknUvYUI/4Hyd6aH7JIKGVN7dG
fOK5UTHbnm7VM4Wr7SWZgN8xsiSjwLU1kAa6d8KTzWI6avKPHolnx/e96aPSvvCT
LT6RowCSoSIXLvFefmQD2ABJeyk4ae1XA7Q2oQpG8xe2xGl+yn7LboEcczPrhMSj
a9TtLlQFAQYsis+s+ed/A1CTf1iJ66auZct0LSfxcBGwc6aiQFGqXQcT53tTkyQa
AK9xn6ZztT9Z4KbjU2ZKWVs2uBottLny4DNiVNzKduwZ0HetXqj7bEBwjXaKkbv3
RR5oY0xKj41vs9e9sc0nmXc1k2oVIi2DVIbncUoUb9gXzx6EFfOUIsQFzog62nC3
klkLQ3WGe8o1otDBaGbmpKpAKreEv5JmOPSnltffOmvA2bxjS8SxPAv/KE9h4nNp
cR+xo32aHX8zL53wEe/8OqwoaIPrG7xkVUkCOI7azvdR772+dbAPI3+kFluOY7Qp
LX4efBFXTvlDuBo9gUsG3tFllUrwk5WCFlfOWlPS7dtF8qhiUMXQpgpV/0E+Mjet
Jlhler3kbnTQ/47M2u0skYBHDkTwqaBjH4hfTI488Sw5/oDAMT6ILmWK5iTdFJXm
q4vOWdTX/lhBcIL5hvEm/2+MfWgFprOdZzPp0M6dhtxQEJOeczpSB/UayJytGUGh
bZVyfpHYlSfZI8bM3qn5S39bjC6XPIrGlzuIqYiAWsjoq4Ugop41EouEw0lBAS3C
3oDfjrWA4XLnY4PynaTkztZ5djZ477+LbTuWu2XKUYDD4Idh5k92pGwaaCdqENu4
U/0nhzaHB22UsCNmusfl1tjneHjb9BSjPUVXDAAH0HMLkrg1Jmd7gqJoU3MzH7iW
CEQK1jbcdd8hj4RqwUG+DmvTjDKDpmAtGMCp5y4taeW5vewtcryWkWVksagv/jHV
yDQjOdsGPzeziYPZyuSNL+iW77lwX7W2q45RtiR1EfTrqFBiEKhxAubkctYQGwdv
80R7nGd6Jm7HI4W4pRXEUJHUlwP8x0oQ/mtMARE+INUjBYm37fb/lLKcdkZXXHzo
RVrVUc14R5ZbABcImgRz9cuaEAXr8Ccf36oAejytRHQ/ySP0poHJ2eV3fvcl69fz
QSIbncBXjV3oIKXqxUeVE2pjoaXONRysfnHDIbA+IuCF6n8V2PPUY0AiW6gMiMO7
IS1njkfXC8e/IZ5ptosUWPdIeItMdKm6ff4xw0QXGPytNI/u28a9ISykGWtgWekm
kco21lJpalqmqZsKw+9fvTFhh8EO0m6N/91OaRv+VjWM1xvpf+RKTa1C1BS26Q8E
dgvd5MxdeevrY6w/XX/yu9imzFjvIecicjnWZMAAIZOtYvDwnzQCponKetpP9xIK
UMkuPtrbBdGxHwspKtfTD8DFPb5ELy6H2V9hrJhJATwGJN1S9qvDxqG38LJikE5j
pMY2c7/j9qgbt8cdbny/vrpK10FklGq3m3iHDHkDrfw5JBXcQ6YiFqWYCvRktYKY
LVrPlsLrfGnpyPtkcgKqUF5l5nUR4s1qgUJ3ORJN6GtlPBEM90GiIfd76bTm5XjP
nxAl//jbDo6z9mRm+Itc/WOyV7ZrEUor5y7bJkpaPryTRjaUtsrU4GLWfLQJmcRa
qdY+L9fpu9LBBXrTw3YFyOgX13q+q3sTEKIYUNYQfDzurkIwtg4aODMvaYL7h7g/
+/cUxGcilSCq2BFXos29EFCrErsYo5fL43c06P/j1A/TbUNMHbSwtYHG586uuLMR
FI85GNg3fnw+cwQvoqd6k41gDWzEGM/MHyWPCE20DlHIUY8Xy1Tf6Jrkf0gAq3Ri
9HQU1zgFQCOaiE0R65vi4q4T78i+ITl6O7wS9dTDyu7i1MFAwAEi7P5EBUKRM87j
jMMPaC0MYuBJyhpc52IQxT63Qad79Ttxmccz4/QaZyP8LS1cFVcH8PNrhRtuq1IV
FUuIoGDGD4BJX9/hz5vSY/0VP+cDH8nne/mnAuYuVnqTtS2X3DTBnFrzuAv/OsVC
qMoNGEM7c7Vo8ozWHzd54dRtmAbkMnhaZgQsZLzbnsIxZzLru+bVH5X+xc2JSK5X
KQoP5tc60VFT+orJk4ilTDH+1y9U6PEeod723M4w5wVx/mtLLFRzevCHNVzOH/hV
AO62vX+NbPLC8qofgNFbCDnB/51B3TV9KwHtF9fwVse4rehEi3tpJNXJ0vDoWRCx
lx5akiV4U58ZF2oJFOixHC3ER0l5v7HZXf/Z3vGhB+44+I8sVJ0GRa4tuPtgp6SF
c3tJp4HmsVs0dZx3ae3fERmVXyA8ALmhj7BdRJJovx+DlsRwGx0shrYkISAurhRO
/EcGsB41/zOJYbBpnib6DBWn4spCUQoDjQTdGVqIC/TzyeE5HB68Gr8ZqTaDWteM
33d2Qk7pc+xxACBpiwK2DWFsy37KUdqgL+Vgvr5on0pop1z7vrNGqezXdjVZeyCN
GpKJ9IkHrFdGc9BBvY3iVbuSgrbXJ521G/0kxIx1LETOjAS5JHZUh1VEwn6MAflQ
3ZAXtNev4UBx/REE3AbvwVOvN5+dq4TE4kQ+qoCjDXN4ad/O22Y1h5btIcMGFgd2
3DGWPLXPYbg7fPbFeBBf7oZwAG4Li75h/5mtYrR855PnZ9uRLiQ4es/MrEjTqiBg
ob3CDkRa2qQ/v4wtWmMeE2zfpyKQnHUu9jhSR2oowTVxzRaxBGbzJ36XzGxSFpsD
2ts4BKNR647aiii/TPLbv8F+91osbdw4TIMa5jvC/1jRmoScBM6jtA+pJXN9IipI
yHxaccm5J0iirlkiiEzZuwpBPdxDenm2Vxl1T/oexBwoPRzHXEHuziuAVaF3QKAz
FzdFHloMWfrYWPqx8KUOClJQOglc/DLOysx0Rtvzy2BXahd7urRf8WUfEmL1AEYG
WehtN7fajjzbZWYqRioB7p/Xa24siVwnr5rGI/L1oaNDQHULXQ4JMXBKeAOqNYEZ
3pvt1x70n9vH47idSjRs4VR8VrKhoO1ufb1zOAnYY8fQ5DyvAp+8TUEGisSxoTim
0JbcOMPZZFs2tfvh8nGZq3J8svMALu7qPRVkH6rQcUfRmqDmTxmbvUXWJH07gevh
HagWHUso1Dhp2mGr4+4+69kHtUU26LHpX+Vhsycf8cjhx0HZbbsrbdnGIBkRkOSW
sIQ8LzpOT6J1Efmz1r5AMQjxjj2Pfdps4eKbdleEUsl/uRfiqr51oDE/l47minyG
tBtGwzixugankVd3oRTb18IGC6myXYtrwTncXpi883comeuHFwZRItOTBAaOoFNw
9IrG+p08B0/zcEigRuXXHJkMTAU0Z8qMNTTDYdLdDJQk0MX8o6nTDfKZj6k2ZV6y
MGsmoM+t5XymcQOZ9SoP1+cOvQ8hPSzKdwuWR16/qJndN7PZMpxdfwGymaLNlFZx
VxzZKoI3+LH+EsVOVA4XFRoRjnmEFkQu9qQyAAg322FevnlA7d/LHLxwqH1mmnU0
8SgmdcUsNrKJEHupEIV5KkaPzQ5ay/eOqg0hCphzR5h22EEDYYfKvlaK4J16HL8B
/djIbpyojWYD1HVbuGWzODv5q1bwXfGaWLR1L3v5SsltHrZUzUSU9lC+MQ3By+e2
1t7F7keT3F6CJNFERKgO8z2z36F4/hX7jmOjoWHKWCSl5iT3Ccvuz9Mm2MfqSmXB
UPI/Bw+uyzvLDix5bgXQ6rXllwMBQTDxoymMJ5sAH6iymy/f3cpJPyp08h2ovLfY
yfbbvyXeXHzQERKPGPfDutNHureJAEmOlYS8abIoMO0GruOPqVDfjNuV82TjcaRU
8/mdaJSkaaIZ3sHO0QBFjU9I6u0eHRCLxiMHSLmVcaYbTuKw9PSn6DSl65+pYXyw
j7gYDmq4gdiU/YyZGSYAIF16WWav7IB0cMtlNvo5fiFc3o4Pb06lJeBtAc6myD09
sAyfHm8EacPiEfdFemhPCztZFuWcCeOibjKl8NzurP338wca8syJXX5kDSvPA/G+
CdU1k3i+7UWc/EndUHHjAykxvA73hVfQzjnbkj/E5zpdKQa+l9CvY7mk3RfK6izS
lWclpQzw5+deEq6rv3Eo6GU4Yqs25QhHuuZetISkUYw3QNhqLeIp9BMDG+ZH85Dw
Tumuyj2T2vs7gUXljbi+fn7E8R6bM57yOg+RmigGUuOlOHPUmqMi4VCTHRRH/EJC
DmmgzIaqOmY7EVWOxn1oW5hhx5ctg31yPW9OvS4JmbBJtqP6zFrSZICJkx2fBhn+
ofgnjTUd39ZcR9zKOHrrHyjLU5I0FnDG+XBgcUS9y4z34LSl8rlDzvxWfsRIDMLQ
JjTlxhiSHWT6qhzN8XMuKi7TGlBItidj/mFOSWMRgM2rUPbwVHGFtnLlWp1lPbqc
UNBeLZPUEvmqgZiQaVcRnjr97EGNd/a6sAV4jeA/kupvfv623BKwAN47d6dWJiR/
PXx1l+siI5C280l1cYtn8mW0jzVI0V9vKJq5x2dSth3X5EdHC1j0+Jg3HM6TqUO9
q81bId9oF4CFGFAd5j3Ilc1H6kT64HYFc+gymS2zVpIzB2DaDFnSDFBD18Yf2oVn
qc7t4e8v/jDlDlKGYNc/B48MkcAc3ULZO7vFTx7Ggdd1eVeklQYYCrQ+YI9KWzlg
Kx9P2xzMPMg3wr+vFvRoA8T0bKmC0Dft5MxbyCqD0EuGjRzOcjt+hPpoHBkgvi1z
1SwnFkYZhxJqXpX4FzAX4Xs17cT5uQRdTmZAhUNsCmwouF8NiSgyduT6N4MsJ3ZG
jLn1uaRwtuBmWk54XarJrn5xdUt9TyDV3CR25/AcFNwp/aCH8PBrF2EwucXyC4o1
lS300BFVZT0gTOZXXfR8u7tFV7Ofv3L9r1kjW64+4oi3st1+IPHSrZHH/BxxD1S9
MBkjSg/hqRDg3JdLNyfNIYbjmpCpj++SJZ/uGelWj1Zz0mnnpTzCKNWtxDtBVTeb
Xx5IumbQEpTBGPB79b2piMB6jqiNicQKx1Jo7kV5X3A/M7VQXfUDmKBfBijD7nTz
EAzWDRxGOfbRWe/r9HeuCrHXrW5LlRypZIhMQ3+GSErbNL8MocepXAMxcdXuzAR/
6bAi6KysaYL8qatbJ963WPDaWsoVnNcCQci4LP3jCzO+z5oaRv2ttmb7Ld25CMjC
v8XI4L0B3iKUHGBTSONJuo98yJjb+xvBetHdV7JLudpAVdCWUfkWe7XHNhMIQvfy
D4+eEYMPw3vcquXA6mTwuGMTXDf2pF6IWqBMAw6fChIQZwCKhYPu6uaqKWeeH0mr
sx3gvQNymJxEkJmbdDqWWpGAg7v3iawihByXuDAZADF1rRk6LiKFhYYhVQ+CJOnL
ad5TlxU8zNRUFd190r5EfUHK12dq+3peJAwIT7k5IazCvHxLpUF3QwYklU3gjpQO
oNKuPoRiO1BT5TxqwMoV/u5Da2SkcKe42IUKSfgmkns2XzinS4LWji5M2UyUZrCi
AQ5NJLDbMjg3oKAbNyWQ10eQS4xXrWfVaYWGqVxIJ/4O2YEKiBOtJDOX72foNuhu
F0539DYy8CV79pWFAdVAAriVyvCCJRWVcIP4tXsh5LKM/sIPhhaRYCowgqwG6Y6G
ypdaYW2BXCsWaJsR3hsQfMK+Tjghx9+j/akBproZNCz32xoXP4sFWGzEqqXLGN2U
0gR86/7hPMU7aoFZ8RpZJbSYPsZ/btIKwjtOR+90VETvxaVhVQMv9OEfSrsL2QmB
rPnCBQ2W6B4NRjIBCM07DRR4mneCO4LWwdd3LcqzdW3sz6PzYTJ31gb73pbf8Knu
FI/8P48AA7AP88YHZfb2nLsvi3fR/zzFeJLjrLosTKWk1mEubxlFOeqEzi1x+ABw
Nq2INFdmraLXaDd21adJ5zxgSbH3dWEpkv1Daa9523BjQ6ShgAdjhIs/M8l7Lw5T
klirgqirzWgrU7NAXL+f4wjg8h/lEIX2CPmU+2o6hhXQpJx+2Tssi0dG20TQ7VT9
NMKZM6TyKXCQAN//6HYwj/De+jFst91/P3G4F1g7b6wPd09H1xEhPOW1Vh+TLzJh
iONEl5JVReI3ucv3/4LL94GsksrTcNEna6+zB6gQDPra81murDvAmOh94hvOg0GI
ECH82s84+hrBdhH9I2SH8irVmZhH3WYI9yFzSVuBD6rwHoKxjtRV4ZhRapUjJY1T
/5lEXTaopJr6XmE3wugbO9lEAZRa3l5ThrHxBliruL57nktIa8JShvefN0pXSyff
dsfEUKFJGOZWwhm/89aTyaNHjnI7WRArMhlLmLGF4O0T648ZbhbwfKr0xYp+MV3E
6BhUqBg/9LtC+7MFkKP2cXv7MZbnX36HJOmneMzvgv1x6jBTWKT3tabrBgPUUpLJ
sSlW4OSIMQpeRIc8qT6YxCKdHv+S9zo8QHgpTaaURPgORG7CrVxBX3i5SBfTlSGY
kywUVRKCdE8xNHt3UziZeZW+t0fITHmnv+dYkZCY4ixqsUsY6G+Exj5EecXqQ/e+
MSCtwLHfZpXc0N5mpNdZ8LjaBtPAHiWvSyKchgOklpUOoSNYRLHFleMSbjQNrwd4
mDMcx1b1/Fr2rtUDL+jb80MDFYZj8CiFcrVPPdqig2NG5kJtwvwSzpwx54LEiDKl
G2lRPXVJb+8P3ntdjFxppZQtZx2jTLDeP/gPumKggW+4snIv0gjoFW5VTLNP2ooI
XpoUQ29siOylNFnXBQVxf6OqKYA/l/0bRBgKreigVVW4h7kEMqWdcHJ8ae1/vZup
jAjeV62UN9VIuEdKbAD7tiVAGFUB6YtWAfmapSpUJlzX4ebMsqSLApKWjrfI0adc
x/9TZhnVkGQbYFLdZmvnYwz67hs8p7PYrT0EJBO8Lg29lQ/U+631F1jYWe6iklty
HlpEY3OCy6V7P/GWddXD/ewl68YTmlMgEVBF6WMYZrM1hGmlr7M9NePSaPljrIY3
Nm7/iRjqs+ljAcGZ3nVhy2x2G4WECKa4BxNtPP6GshbvKEpPJjOvwE1NU+19/wvJ
1zUkHHoZubS5uF8qw8z+xVIeaLhzt/7EMhtnF+h8c5+ALRf74QqM1Oh71mtqMkrz
sRHKRlYjSvBc+t359286/6eoQVRkcvy62BJBNru+nF6t8tFWQwcjm2zoUaIbTQ4g
K+1SCMe5D5iFzFZGryyZq8kIviaI6ZqnIyqd+cH1PKTKqxFpwm2ETuqcoQUMvA9j
GFDC1mKXfgBo5PiRb2XBLSL3gQtYs4ZaYG3kmU0UZc800wkpTr2hMu8vIrcSo8O0
7vT+6Nao289DhkCHbQFSwoHZoVvPkRWbuyRmxjBolmkLKHebJ0OfSEDknrByZlZq
AuEioNROQrGmtDUOn8Ign2uo4XR4Cn5BBZLHRQML5H6ighsiIUsxqMmnyHh9v7v2
k6S68Q3jWGj45SvuwsNWREo8DX1TT/yZ3LkpPVVEb7kCn8JHoFQi9yvLcGkLmPVe
LT1PvaHL6bS/RLtBgQut0ZTxY9wNFP3y7YGs5G+pxxaKuTLjD5e1J8UvkIMeoZFP
YxaaWudPG68HCDZ3o77YnF49vptKZVWb2Cg4Y4JMuitZBsqm8bfGrSiCwihKkzd9
QtI6XD6W/aM8bdKwbaqp45xvab5QpBdoWNQ1LNOCHV0UBMMgMgrH768zBBkf/ho2
NM+9YVTpwuHlTO1QLqzR5PLXobzb8cAAPqvMJnSa1bnNx0CvXrIkiQHMlgpeDwq5
qVo3wiFz9QDBhAVNVy6Qm36lO1O0WtMS6hOC0kk3RVx889xlEfTOEqYzA4A1v8dy
5oSlDziokxq/jHrjv75KHirYiEXVGI2T3Ju0oLtFra40t92KQsCXv/s7ccp0oMd6
PeEdxQ9IkyV4AXhNoIhFN2LcSN7qifXPcIrtC0PAVy06uEE05uwr2IPjlyIR7nCT
Hf1NyYigXQIxjI9iq/Vv1kt8LaJGJ+916GU2/A56pMMAzSiDmNMGH5RwoINUzRo2
JNxM5HoEv1WQVRf060atM8SYl0l1E6/2tVPFAK8sxn5FQJsHvr/4MaymanFgHoju
0mCv+KAWL846TEKxgS65RurSUY6sP9TwyToT2pYsivceLNWWzI3PoRdx+/6v2BL6
+1oQo4SuWRpKF9kHNvTF9FLN8YLqzhwRrUqUEzLBxOYD6YtPebWQflql0NB+aRVc
GPL9TzT6EXAavJCPKj0pbX+hwG6j0UgA2+U9cDwlqO4snOBtavlnROMAPTXvIkwK
5M8OVyxKtJTuFIXIi5aPg/oZHYacImOytQsIEmreVdl8Em607zjP0atppxtnZPPY
w479EHkNi/zwpS9qFnVkE7vZNO0xIMIE7Pzmi/YZm64pUFqNvU/jYwr73NjyiAyR
ie3tcpuvxpOm3LMjf056hs/ALktSkJHMu0DsjAAqyHG+onCPW9oRLsPqMfaQEH8r
tSgPg4Qp/LmOE9vO3I1z3Bwyb2Jnb4U6TuqCVQNYIK6qvLcRiDtNS0sEpiGOOQ/U
CevcW9pVQFr0GCAydQJY6D5ngNvYCGzlw+9Qm419kMXTWdYvJnKRz+HlnZm1F4rI
E4bmWHw6arbfcfHcZ9qf4eMPu/WiM5MO2f30IxKIs0B+YK8N1LvYa9bGGRQPoRgX
y7gvsmI9c6KQUG1W1Sop1cPoOm+wES5ShEu/PB6bMuQYYcS+aDm1B30Vv+hMd7GP
amrnHJTeuX1ohQYTR8P+O5RtVKipgXTUYOrmZqC/UXcbANP8lX+/dyHULfOmSsAn
UpOgVbOoDiu1jBbw1MsGq7IaVrRu0yjePgz6gpxKHWMHy90xbZr3eZsafDQAwCVl
IIivVestxW8W2rDkZzJd6AJKe1xL8wrv+05qK6NJ6rqvvdgHTHa1MBexY62ksI/O
inwBdwy6hmy8bHVgicR99X08Dhhk7WXwurrLYPJsLFPe9HTab07fZTFiYe+rT6zR
BMAI/Tr/xD0Vkmkfxt4/wqz9EsR/dfGXqGz9/52TG20xcbr7LxfKUi76t14sNpmR
E9sXsZ4hpWxKVgZKkR12Ut+cV9dru1gLhg7A6kASVgv/gSXDu6w1hOWo+TzuYAp1
dtTi7Fn5BPINW1+WpR7Dq0TkrCm6D58FYmMGcPUVYQ7VXw0DCQxq1wtu0C43HAMp
hAvb+qKwWz7EV48gtwk7FunAsYpD8O5Lsy6AbRrw379ACeKSEjKS7baS0pt7FG94
9/vLe+/8U7qn3paGUbfIO3m6rmD3F9QXWwWNTboBl5o6/rSRpjcujEpHgOmbXZwg
/MeIhFa2U6hB361YYQBy22ZZxdEdiVdmha03tCtprRaEHoBwbq/Jso7jxMFEPshn
9PCqFQ3sH1wfUSdOglc/DpQkXx/+531kvbWC7qO57CQa9o50gBW9VZYYvjxU2/pr
Ralw2SL+d1HIv+gS9XMF+gnGUKugFnL/qv5TfSyaRFhiqy7nl5dT7Rcnsv+31nJb
WGkSIV/suBtQVsjDK8+PpKU+4QQSv5y9RpkNgbrDjSA+02G3XyoQwPeNe2M4tPb+
SMZHFMKvpoEO1LV6gbONRmIDvM1rJJ7paIY4o1DNf7hBJxeGjPOBllCgxaW5iE8S
r5carYO41vFLeMfAiWfnMhXeCP1jt8w2Og3Fls+mmg8zTLHS0y6EYqVKg/wiprQZ
oxO2QKIFlJcPp7JtJkpo3tOqNagDvHsLVR1sTpLhY2Zg7qnT8aFkqlIy8eM1OsJV
MXrAI+FXYLIVsqSlNRZGW73g2dX4zmSlMC2G00+oc5uK0dpOV2zQwTAKPGs4YjDC
4ARutkDnvsOGljD/UsOoAi4w/eSLpZ2VZjieUGnLAYlcXyl4DC7B4wUdZDIAwS8R
nbZx76l/LCr304WmJeMKXXbHjvsz8LHCLM1/56s80PpPBQTfgFIG8oRIyN3881kl
oDSHxl9b/AhX3Ji/a9KaW7MiWq/H/GTLuzbIOWZemFO70xBtbrPwFhqxNGO3Tr1/
3kd53PlAqxkHHjJZwdHICjGL9oEVR22Nd95V68gkbWOvC2/X2HXqVUY/Yu5pRPQ6
KiGiQjwxOuF+aNZHug4jMj4bh2sroeLl6/7OgLOdWC6boXG8y50h9mlzZAyszOTP
UwCbrTDG9Tt5DBZPvd+gNmCh3/cvEOiUTY5Qhlv1CXWiBcezY6OylMTf0m8RGPrp
uot/nfb7pok3oWJDlSWahLjVtbe49sCvJQ6XdrZixis6A+nXtFveJmmmspYFaErv
ly3chv0eWMXqyWrRmJatTH6Ome9lVKHVSgRXVQvHE+pf2ZS/edeTnLQ8FUduVcIm
1oPNuAdL3N4KnQiQjYbKqYWvhbWRqScj9AKvQM3G1GCvLjWux7MXh1TqodBqZjJ8
MiiLNvowGpq77JN1aLb3isnmBEvyGDOeA+wSwsffcro0nT9yiz4gr0GOfxB/YiDU
QN2L92K2KJrRz41AFjcD3/jLvG81nHM+vRm5i4tkhh4FSg4PA9iueLcPhUJfnNzs
dyRqwdC3M3LdtmlatWMOx2MzfKBSgMgexiVxblaMLhZRZ/c9m+S97IEGZU2Zv5Dx
hJvOTfJgaQgHe9sMDyFWgiJCUtx1wnJbdFtsU+0luc+lR9c1qRybbKgv4dBT/i4r
tn8tiRwAT5KZAM7aX4qDBD9gWbQEwuiCZTNcJ0DIs0wYa+TDJ/GZlI1MEwTQhRAF
IEn9Uzq8DRGmK2pCpe6y99DWuXpfTI9+FF943Bjww3Dq+aJI+OFWgXBJOt7ZxO+A
v0oFnZj0xVXeydt12tpgOW3TU5veDBuuRL6m5pJEx+j0PkMPrV+VE9MRQSnIiilO
ngu55xSj/DgoT2gWfogR1yhHWFotQx2ag4rEHSgD4dSZ8uLXOHXKkTqdtpK4/MvL
QW6FioEymTRptRNRJAISJCekXjtIvMb9YNP4JT0FHne2XBtKMO+a3r3uG8vU0ebl
d8JLxtGnsCMfghzPKdEiSK83TylTo/lz40oO3TiDbk9qrFFECrDfweDGHzFSptWv
D6cgi3te+fm4GfTV6S9vIrv2vsPPdSskfGT27HZLaj58Ou0PCuProX6lE8tulwe6
2wbDNYK6LpfrbCmUpE20kdlQwJE87mWwPLX52NxnJMwXM5sgWdRfksBvFhpnUPlM
PyA1mvuLRPuoW74EuMZRzBtWewDi5ttREZdeT39ddVtZtoodJXYHBA24V5Pf+1B1
4ztOMmzayqXPcddRRSre3MCwnXAhf09NV71lWMPfik4K0ndxp0TfnbggaBAY+Ges
CfqYAPaLNnvWtt2Bylo2aQcyi6KXItRwbooBeF0DLOeWwAdqEj5wisiRMjtvMLJf
33sw/ZomZnwESLz5yHALf7ZeMl8p3k4P2JAKCDpFPsvvkCCSY3XReabQvogY8NwU
VhgsS9HFD/tSCmBF4YZoIDi0yMw0PQ+W6XiOxXuj/HzWM4mv46E9VhxJFkHNA1CU
x1hhrglbpBQeIo5AA8D9YwIwih1dwTlcYA0CE/rAHBEDXrsJ4cJwevkbKzq+G8za
N5Cf33eulnmMRNjciY36BGZkjImCJzkjmSCE3dl4He4RKAgt46vVW7smFhu/x/5U
Sjd7DrIOcUS22EHRnufVJbNxDm/ZXpRHHPNE0DftX4z3xcHtzegzW6RWsn2U4kk0
3ztn8tM98Ajoj9mDlbsgVv+Z2H5baHr5kz35ptaM+7++jXxfhNy35svN+IYfiN0Y
Df5nZe9yiNQQOlOU/YEKPRXeORX6uCKsK/7bENMgSAnfiJuLHSOSE1AHImf2Banm
RJzAtwcqhq2shk6Az5fvzc27smesT5Mfs12cO9q6yFZZ0AultCOmQfSx4KM7gsrk
s5rHDB3eN35ngHvSps54H5LjndPAT5p+nmdedUOkdc9OwqlH1gO/97uELbNtRWdc
dR4+hdfN0jKLXNdrokIvcPL4AHbDF3qzOYQ+D69BLlaemdKwFkH8aHwJas06/oM8
8iAbZpJeXBzewQ8TzfsCzmiKmN0fmIiJNZJRAn2PwH+f6ffDMZcqAyRYnU1pvbKa
KoG708jGCEGKG6sv1d7zrRG/XKZwZ0v+AXxUwCgPE1fjgB7+O8+lxvfX3PPNuRRs
wpnzFaar7ud2YftYrgLKvb9HZ465XhCcgNOJ3CFzL7X3qKTU/HMP1ghbEleNSvue
q0Z1NdLrg8t0n0ojtww/0Yeti3WpkJt+Ig7WVF5gk8+shFM5CioP6wi7Yo4mtGD4
X3DQ55kcx/EzrT8RlwTFDDVSZjbV9JAGfXBEhUxaX3X8+FlNSEhQ4bRy98RK/aj9
HkfuEUI4r4E7vQE4qSdq8SDRNIixBbsbOVtyUhx3g9foP8slPWWv7k2+cwgL6PKo
nSCW8Kgz3RVPWEpniaIhHjCXAwwoyiNZ/uWqe5jWAyHQPRy5ooPfsRodvOZi8/bo
1lQE9cazllWZhjQcJru5vTFHTcxT8IO5twffJOG+u5cODkvENCb5aGlyVsAbB8Rr
i2qj1LSSMnGqFYZQ72hH7nwGFb/7prR9rnec531QVYRRPtrMvqFd0k74bPUYFVmz
NOsIHbskU71dsK2H/ZzOvtdwHAPRQHLM/aCvh8UwKaZu/QZ7c0dznzA3C3uw5UHw
UiIxbyx0cbcoOWg1pIiQayXXKv8T//N2P0SOzwv84646ZHlUDKs2L6lDOQj6m1EZ
Z4ySY9SMqwnQe4WiST7pHh4ZT+GZU9fHl1X7Ob4HgaJ5Q4z5YTkyV6zzGNksUfDA
qZe+AC16QtzQiG39fSHBR/iYMvSC6zDV1VSQzDU2J10fZKNWhEAgnObzwOw+XO5A
SClKZ2l8XNTyA15Y62rmhzWHklsAcFF+tUhcVGko3gTJln9DPK1oRDO+yFnXJf1Z
yiixODPu3zenMeaK3TM+WuyE8plYgQ3N32RtbLKKB+Vp2jua45x7GvpfaVthm+EX
2zhXQo1aOynEkBW7lgQkdH3KrysFCk7D2OiocmZBjMTf48BG32+cvwX0qY4bWQWM
SC8LRENuob8Y+IYTrf8I5eEyfBxChtRSqcBVh8AJqg6sdA3KQNILgNhiiWvrdmH9
mmLiiZxTfs3/nujTs/nUsnf+OC700xPtXQEytxRWHxXvSZfHYULmeIZrJTjvcZeT
Di5yePQgza7vk0V7G/BjfS1m86zl4e4ZA73x9fuLNWkD2IWTiPssnrexRZrFApk2
RVhMwo90fKJf44CNpDoUtj4fGGe247PY/RfU93fVj2BxtAPSX9eeLUiwBaoMJI6N
F2igMhhFU97/x7ZgM+YfVBUph7Ahn/SPj3clKVIsIKvYPGZzTpbqoYStS206993X
TUBam4Hr2V7eknSWlTtdtPOrxWPZD8tzAUp3/hhgBjCfQCi1mBavw37ayVgAZ+zn
/quASu0ejO0LKXI21nMmbbFReI0KREDOdfX62N6Sjl2z6hVsTl6qVP9PyMoU0E14
x/hFJe5VqFGNr6YpYzM/Dd/j1TlL8lIsbVIlDgcjETVERXxQZgjVtTiZIWrdGf0v
Cnujgkfv30SKyuxnr00Ui4GmyBBA/l41j9kPoqhWNgeOS9PaiaaRfGUoyCmgUFTW
Q8Uca3NOB4b1rrKeCvphfVbaqBvde868qNBbVELEVaHlVvZuBJjexGBYmdcgARuA
tnKKnK9WBgucJ9U676LfexhYgI+GvdzuAWD3qLq4PgLBG+nuiir5WEuLy2T2FNuj
2A9dZfzCeJz07WzynXkpSZMPBZSUA/k2CifWbmAWevSL3iq7QKl/9kegfQ+jTooK
4ToH12KkTjM7FHFpyT6vpIzLCL0WqU3GCZie/0Q6uaXCxdF5M5AarOJHLvgTqIY3
GIp+bn262DlUdxcx17w+3VwjrBw3WXsO+1bMxrOLZQOL7K4dwRhbL0a/DWd9oXq1
wVHS/jX35Mos3JkMSndZX3/wegZpCSSMuhPwM4LOen24J2ROOXnRSYBvajhHsGkj
ZS700Shy9974uiReqlvPHN/EUebepkvT/7PYBhzrRbWDuqY5u0+VatdNyQz1volp
30eASEvEceRa2yrD/WjRQe8eTupW/st6C5ISIaSRmx9HUk6BuxvXwkgChx8Btw6u
TqEREZPapPPfytQDbTVrfXVeySI54q1mwUy4L6mDbFAOq0DWwY33HiwSb+HQb/gt
JGPW3NXFv0DEBugaXTZQ6RQIWBCZVwnEJcQ3XclxEupksL7X+d6667FStfVj+5Qo
mYIEHpbiKdRJepLW/jPV9WSkFdYHJk/QVEwnnLAL7SHqF7ovqTE9eLhprHy3TGDT
E92mbMWLTNBKRE7rzUG4DC4pqqfJ/42NE9y3FwKgwNYOdwuIWHX67Huj17UOTW57
9O25EH3+kOXdVJexT08MSchITT9LwQDehCJyLKc7bI2fTDVOCNOabgWYLOb+Zz/o
ysjkuwhkdi3DQr55cfIvh0RlglZxe5wkxuxBs0mVs+fnt/uTcq2LyJxvxarXPWyD
ST12WyXlCSNtCk6YyZBMOZt362BEpE9hAcHy5ZaGr7yiRSDEmP9RjYw7JGbOxlZ1
bY5eoudUl3LMzedHzjHvQNUzUAecCkoyN287fGdkGl8E6DMWlHlaMyzoClW6H/p9
crixI4cjeo9Afsde8GUF7Rr47v0J+OpB5kWD1mG28JDDdDqaptO8z2ASNhzdsVKa
1CcwiFmi97dzHHsRbnYRJ4stmr3OLOa8zBJu9A/jVsHuiScixUKpHALBD/a3YrAw
Wxp30GP6Up63UZoidoOrx7+PMfvN/91hauUZG4te8eztSM/ViJIpsQWyY/W7WSAJ
l4AI1hA9pUZLxgYJia1Re48FlVEjFBUPOYtrpVf6I3JR3M7NI48ZtWbvPaAdWOG+
oH/RK1F8D/SkW/MEcFFh+Px9o6daOmrWx4lZm3kD6549IaKTO5O2LARtJnqqpSq2
BnyvAZ9IQ1kCiUd98mkhsg+YG9/Q59fmEm4+UuNz6dVFf+avADST5vtq2O1BnvEm
aCSL9lYoOElZQW5uhjA6uFYGkLaK8ndZJZjkRprkC5Fcoq1m3SA4kryvBW5rUR1X
ZIyc1KBD4SK59hRasNiQ6gXj8a88g/KGYSlQPMAUeSL3gndGwXG5M5V9juolhKhM
0BfShO2gK1TbUhyZa73QFXuHBZFUtofs5KvqUiYG94W4BYTCZyRWE2b2wOS6zoOF
cx59xDL46Xvflc/3lL/8xHCq2fRfD/ubjJOTq3maFtqYThrrasBVrj9TTYUpgWzN
ews3WiCWLkDkBEemkL1fqr5OmTDY3Q3Kjqcfq2i4q7DMHVvPkyyy93CWxfSlmt9S
S2aXzaHF5iLt32dshZDg4wXB5nM4BXivJFz613cQiuqNehsmYsWApAwAhm98dIhj
PLQ5vKeR7lVCYLM3cOU9gUk1yfKBuY00GtaCSyg6LhCfUpFH2s8KGJsiQSOmaOeK
S4fKhp2fT4nIctZBELrOe51pLPifUeimsydzByVu11YFgIkSBozVEWdA0wHY+pvR
TD2iCwPIgSNIDA3OVs11ZgC2Ipvph8oCYjhD/ff8SzzvdZTe2EOW1ghLvIFWWiLN
iL7N1j+SwAzfn4OHIfbgNwpE5+6TSyzImcbhWoHz+Vc3xSvIuTF1WUDbcFTAdyON
BPdiJCDHeUQ/G1nCK+wURwyRiKsjz+zU/TwLtFLDLYN2FBd/lZyPEJH1bGJd4Hkf
ddArMpI9Zy8kipto7We8yhY+1nk8R8o6vWw2lK6ki9pSj9pts0wGjvfTSrJb298k
lu6g5A62jh7cK6WhSBQF69frG4/rslEepv1GxBtTenFmLXmmMlh5u2pAiu7iglMU
p005Xl7MWF0+ltW9N/Oc+puJN1DD3lF28KNfGVaaiHOUkmXVm8Vd3P9rhrg5s6G2
6o/PTXqu/vpU9vUswgtXKwnM2SISXdYX/tfFc7vhFZBVCq0i81oFmf2fZegCzpw5
oPtICnviudBfwxBVqbmyH1rt6o787WO+0CfPT/ser93pMsTYEkupAO2XysEuJJcH
Q3caUQLGBevwgOVKTWSFHiLPfvz+h8KsTI0mk7PflC+47W/vFB01pMzhRdSQ1n0J
iJirbefu3qPt9k1ifaSzRnRKH2QZ9SA6oeyuTcjw5csN0HZGJG0mSd5SYMXEJZNW
wCa2ViIjSmvrYgnjxagYmsjGZYotmr5m44P9uiJ9pxOvvBBISyBAohc4ZvsFwwJq
QCO8k5nb6L8bkrAdgx0IN4KMnksDivWs0inzpgfU61mzgtdkc7TvqZ7ZyQiRFCpa
h5tqDVXSZ0dErDgi3jTbdFYlKbZ+LeLzWrj9XV7YyNJYDcTqh9S1RywCML5DSOSX
yZSTzi6WxpDS/QZPFo/KhYwlEHtgPD+3yXtVAtI9iRU1YytsYAkYn72ipHpXXnAW
R1Z7bc4D+LFvpI5oYZwRzgpdMrhegMhPgMc8kt1jLs+OR+qyv2C09oS2pgTW4vrg
sE/S0PNCX3r4e8y4oOSX6tjtJxtR0fZ7rFSxsmD/61iKyBkMYsjNWugG1I2GzHgf
cbxy4/La0ZPdb7Md7zG7EdkIwF2RZxBCgRyBVdu+0MRLwjNB61FgfCtINY3+H5aL
nTcM9wzUJpino4nth3Q/PB8IpComDwLKodNg0lqQtIl+n1D1Rrf3znJlbtvPpyLn
V3XDce8PqXXNrIT9RxiL9eGWsgt4NPvyIOkIKP2mEWzvR7xrc4xxkR96t3/JJAXM
W5ZYlHb3KQhbBdL3L8n+6D02do0FmBIT9764zxthbI+jRHkrUFXQWYFO29Pz+hoL
C/Z/bzWWh75koDkcR/slJN4D+gC3Oh5pB4jzxL/uWI0/mcqvwJ72kRjY4Cc+561N
A4dl3tKjUxraQuxRj3VuRWfsKckTSaPEN17Oqkhk+jtwS5+D6+VX2PZk7f8Jh/pf
rPlYoKorZaNrO6sT9eLvJSROLccM3JsPEU5Y9e6SjcCMqHmwMLfx0JpCyp8+zoUK
fAfrHh9KKhQztXH7bIcWTOgXNcP6NbgJ3q1Le0ES202dA6fHNbxmUF47CtFvi73k
W/hekZ3DzTcRYxf1F/lUsv9y/J8RLdPJL515wBtyRGmjmZzirCYjYu98XXndgrm8
JKnC8btG9OrICkLMhxLXTcLEDOxt2df1E1P3ivif917pT9HDwoqWARoSlLIfFjgw
ydKgiSTgeapbvtnZpfJrXbe5fT+iyGfy+y2eiEGp7MFaOSkyMknmFqLl1jueyk4Z
PXgtYQMUM0279y1WCSMcsqkPvzlr6AZXdeiUfIVCxTOOZu8RjjcCFIMKGrLRg0Pi
vDTK+95xSFL2dbyk9kc/O6q/WFeS1LoeIp6jMuyz1HLOV6DW5zTB/QygA5PkMP26
0ahJqJtZkNxVnTiP7YE/6swqYPcEINza2gT58QYEUy3xC2EpAVSoCEboqCZ1cplu
pU6Cwx9P4jQDQBaa1bwhVnO9jOuVL9uYThdXljgqpleos3dVO8w5PZp7/AQ2oRiA
y2oqJnoWzI0eO6ujPWBUFXqgzEHq1lZIV9ZMpd+QDxYxqQKI27PGOdQty8a4Ijs0
hJ6VI1IbUZZXZtfp58ziqJ/wRD0wy1Sqb2VRIZYiHUu1dwvubvmEcoPasE//79Jj
0NBIlS3LaB7XD08c7WceXtUAU6EVuERv749dTEVVYdBH1ud2P1OkquVVl3lVSKDe
lS+WRgi/PctfD29EZKQsbvTF35zBZkZEVnR9jVwu+N7Rj5nEfOS2MmB28x9YSUaC
EI8vukPEx2COmJqHVhwIU/n7yDp4hb4XLbG4icsGbLNJZjgXNMV0is3O+uyjyEto
/7qbjRAkEVxuR9j6Af91DuMUwErwiUFgvU3CoZkaw9ewhWHp/UnPXjrkhh9kGlfa
bXF3fZB4PSCQCSOqsN4ogc8Wrc6IAXq8zC5yIUz37+AXfCpYTEViXxiWZiJ4ijsY
8kkzdzGm4l2yvCxXArc2pVMRCPB1GW6x0lRfsL2vWY2cirHd7115f8/JpAuALSSv
1lGCOv0KCs0G5MSwZB8G5N+M+XH0pKzOwk7dEWrbp5H9XCHZp2syaqtFvztWVs1U
CXZqYwVAtaw/dsbBnT2dFwbDKyrR3agZi4C9R68t4b5ttY0BvkmElHbyVJZJ10MG
8GJux8cx1A6YpZD145oL8EmPweaX9rUH7UFSHGY5ftFx04Gv4jtiD6GK1ychHWNc
SqDSljyXUBANY1mz6OHKvrFPgoWKpNl2bA0kbRrFltpU64jI7qO2du59AtExEleQ
cu2Us9vC6k15kh/XOGCiwN1+agod5WgufG+9/OLyO0BDIMGvZqXCUnjrWc+WZLUy
ZtbA3J6v3KN4IknLWySvVr/zhKG6fLY0Gy3/EqTqhRXQp6a8kdvF+bIXUVFkR+K4
0ODbyW+zC5Vd6UD1mZKxvKKfed2rKbbF3UcxY59QUYAOjHDmzX8Brb9d6svkPrBL
PGoWL7BzsmcYGEKCQRNtbima4oxeFarZTZuDYXmD+b63Q5ZifenUKwv2rHNhKfMW
pInYY4IweGq1oIelqe2azM1M756utaTnDm9iPPzB46g3rdfZvDyAhe8SOjj8+949
un3ut5cuMacMNb7FsbDLnrcTI4fWT8tiiH6kB1nHpou0j28po2u7UbP68vYa21OD
g3HJzjVKsleaespnMyC7jqO1knvRZ5tFuNcAN35ruXT73zeI/BWfG1fabPJz/r7K
XIMAS9VaeatepDNRXa/FK9ud0VnsHJzNmGVV1NiIif21KKVlvjmvAT7h2DqWKDY6
xkVEi235vz6vT2ZyC7U4MrSvHu+QN+3u3lNnzawwTCRztyGddUc2giuyy/jM0Cfz
+I+2mUa3h7vEbyKC/I16ILrnhpKl3SWIxj6yTcS2IzdJPmlBvzy3gi3auaIA069X
k5v+8FMbfFst/q65Ty//ouwjlL68EWQXzLQ8SN7N8mQ1rhgQo3BflGwjH9CpSA1U
9ZDXj0crl0UhZCO2SpRD9O5HQj7kbq2kJ2zUIcAzLzdbR8p4nDUhAYM6FAAR7vGj
N+zhN0bnkklxvgvp48BTsL2Ll+dScBs32OVsNfqzzAV+Vs3I+mfqF2uA6H4fehuO
SzylFZtOwDU4wQdXpR34bgu8eXLRR8e77PkFZN2w8PvCI0J7fhLdkWpZHrmLF8En
LDDx+UBuCL0YH53mK08RNrOnCeiPN7pTiZN9dA4UYL2Y5ZARjYoJRXf5KKHEQP3Y
ITDilMn43BEkpEMB8e2I86r4uV0i2WD+1+vXhAFK8u3bCfpcd+NRuL7K8m4WKBTI
Myf5jn356eYWj5ZMFp+4EtA9HmsUhfB9u9q3mqSad4/9gfsCjM+BlRjVYKKHULbr
GTsWzhH8uJ9w9UmR//HWHv5i7ERj4OFy8BExS3CIika7A9zJj29H9RA1yLarw2bI
4sKB/pBfPGMEYll8C/64jfEj6ALUw7Qc/D9borrd1BdhC9DhX4q8yNQhJmTu0uDL
YwtmNsRyerRwzi/vJ+SwtTOlBgypieZGsk2oTKMExTW2VBtcvJngstEFi4VNN7s0
zfPFdBtKGvgk4LQ+7AkwoBHSRM39NUAV+rl7NcMnhcBxzbNqicImpxq7HEGiFN5j
rC8Z6O/+vMXPYNwy6pbcYk2R6M5wvt/Hixu3S+jSfFUbiBA5X0kIgW53dqYCjKwn
sFMfJrLP2bazNSfmW8eiFUIAmomhTHcywn0c8Sm4fhgta8D9uFhvnvep6Z97UlWo
b4x/WHp5qsF8CI9Qc7B1iCl+SmrNeVgfMbp7rgBi0hzeBlmzRea2znOmYfVqquBM
AovnobzzmzEgpjHpoWmbECx6/aJGUSq8A03VToXIMOn62IUCIDEBB6mVwWe+3jFP
vBzP0vUYFGBKP569Q5pdi6cknpZ6AR96/G5ghfNJOoG95shqwXiNDQuCm0R/MZjp
IXLD9qvxEVXvLwmTc6rAOQlTalT63q6mZeNKDyRIKHXQHqvTqIi+oXTQz2kMpDsD
tU2/Gx5ZPcbkk26t2B+EjupyG2sPhJ4Vz4YGjNoX0sVtb1ChxHoq61fD57bjYJ9U
edcj/5vA51gJStpjahmx8UGU6TIPDO88nP2PZ878r5qh6ZpZodzLZoElJCbsXS1c
5IJUdAuk1E7Sdk848kmKBW7TVEOi+FWBTO6IzZOTQdwZ0hZ7qBH3UEfVzXBeZ3ut
OBrT6TAxhyi2OEYrD0xndtkVvuo7pZ1SdYBfNLX62AJp5YHuyVUkOEQ5kakTL1z3
qAaMF16zoZGng7PwGP0KZN0VcUHBMCmGosHV6j8aXwKws24YspoXSzrVayARD+E+
Wyj7avt/f5/JmaNKndrZmhZy7AI84BK3dbtdrSqCBdoUiHSxEbabOzq7D1H5z+7X
03b6+nlUVikBHyzVU2amGkgEGUsYgf3xqIqZNqfcvTamgTUz/iNSjByw+toqorvD
b+gjaJBzXCibZDyNH3uFlyYAHtNYeAOyvr5xWX503sWRP7BV+/PiQxXWmN5RTqrD
lqdCk64W3q2Rr9XcTVopk/ON1ah195R5onfMw5uZNrZkfRK1jxfxxmPuFxOLE/YK
nPwMPRbjbWetn/J3UUtyfu/KASSpGHh2byE1V/Okq/gBOt1aZs37YHWN5Fna6lvl
RgxC6SPp7u3usP6RWIJGupX3iYGJKBEYtpgppOld45ProB1a2Mzxv3+eGs0WIQ1Z
/f51yHacbhx/zKBdM6QQ7dIDLLiyYZWZ8EsSGaw6frdSy53bWJNzdCd2dZEJzg4r
wJE27ty7XQmtpSgXj6XewfQMy9LFuhN6GupZHxxprXVgi+Y2VRsP/TL4ioD2AmNV
UGc/ZayTQHpVLd94r96ATwkmBc6u77bH3Cyib4EucH2/Z/quPUpN2FKRBAcjlCBM
iOUu977HZLqOE9hvFTcixjowSyQaqdBNJeDoaRwSMpXSby648UiOOlW1lMtn0fjX
wpXTnYr9hXmELt6sUX2zTIIsrNukPTd8lezEzMN2ncHWaeUAnrVhCOZNqnr1F7X9
1t/gxcwFx4dDFKIKn/s3RcTgyEG+wd4QqxOshNwsh+R1kSnOrx7JCVZ9BHRQtx6m
ynaMlfu5yIJsDl/fC8il3NI4XfjKw/8WgKRTFjoelxvs+aj+qb6MYKEWbDqpP6ZZ
0RoRHL2rTDuN4vV/HydUpKlE93qy3hJ/mJ+lDamKH1wYCbPlZfWQUhpRw4Ug/Z6t
RzS5Q0zQvRPOcbwOwzQ7l+QDhuZBdl+Bm0XngvekELiFM6q70PeTOjyu4/HI9Giq
Od8d8jaJYoAPPlOrN3mkTNc7Z/58xZ26p6vR48aNphaOwg2Idb4krcpEU0vC11VR
TJToGeYiLJwGfcSGBRspc+NSLOgK+l5IyZpGJK83nDSBOPi7jANmh4m9ejDCdbjY
V3JOC+HWhZZ/8WJjDSpLi3Gp84ZbYwFVVWrPzkHNsAcl1YYORh/1FeNvEpAEgY0n
VR66V/D6sPzAe8g58MoJHuDWaQKiIp2j3tsQAzKavrvOcx+Yt0L+9eK4cmB9iW5X
j9K8ipBG4eOoY7JZgXZhVrT9Wbhhvzm5YUNYDmE3GBf85BLndgnJXQ195wkNuFVq
7xMcFFtbNJYnzi2OLK9d8edIqo4aLI37QuDYHavLR2Jbc3PaCR0QzDQBT5JYXN38
NIz2YT3p6m/PWJDfTqlTmL24T0gdzZqmv9D8h/0zqGDeU1iFizybDzH23gSzZSG7
W7W3rZOlvapsTx3vT+Kbt7Z53d3RV4/OBu1A1SGpzLNWHm3nqFmigAWH3v4JOUK0
Vvs9vVs6dS4csJfdRVp3lyHoStgdBH6Y3FA8BljAYmJuL7Lzk1+iElltwFQbp+3Q
Uo6MzfmTWFxqS9iZ/vb/KqVymmsKSkG4BZnmr4UR0vbTl0iBCKCyZBWDKLzo0eWe
Z7hUqfAcl3MJZ1gQ3VIrXqHjdvW8V3McrVlDmaArKzLpYNYU1RAc3a6Pstr2Y6ld
wi3JmpPaLbLoEdecgxnAL+lDC/mZOq5avylO9KWJzbvK4Ci+J69xtUZiehY5xDzI
dg8SkGN7l0uFuUaN9DzFbYmpT95Wkv2+ZaJ2VSDbC2wKmYQvM2YjF2BBF4uDSIM3
Oh5uuqo4MJ3HTZKnZzft/Q5TtMsf31BtKuXjZNf2VjTR68JtHX/q4hsIZnOq69y/
HL5WWg79jwrzGFEI+S7xJaa6hKVTLegl8uwepcWckiAiL4Hxf1sCans/d8quW5QL
wD31P+t0Bgh7a+omYHOI8vkjB3rlyqEVB9+MesUy0CGiQfONOjF1s2a4O/QNKyyR
Oz4Xq7edsK0VR+sC0SHw4pyecdS8X1dN/3r7wcHimBqPbRTm5nQgFhDeXH61kvP9
bUVaCOXVwBp9fexggWDb1qP3kJLg9uOYPkF/ojEZcH/f0wMvt9sSIW+3KQvUupDV
LctzsnKiNz5tOdpZ3AebzubhjK/NYmMYhVk4No7P+egdn0WQzrGc5fadiP5w5OS3
drHq1e1UJsI6gjEufm4WdGF7iil7e6UBZRdoPgCpyWV3XW5ahURaIZbRj6jnSzqk
ajXfKpDGYtok9IyoBa7XvXA7X5u+bykV/x0R3rwt9cg2F69ssJTYJ2hhBBBwyj0p
pH5VP6Tt55FP4Y9kP2xHFFeUT7j8f6h0l8f7Anrtn5Hwv/li5f+XC7mhsmldiy77
F3Kso36kK5KEajr8WdxoM06RRrlvn3MiIKYj2L4XeEJQUZwpUI1vPQOdnJNvu5Zj
N4hahvt5n5TAjGdTZUzN/w4TjtT+9p3wVIoRWjIT2VpLILBUjKc2zWjlmdHgmJ8O
uWVN95gXMEPyHgkGkyNu5kbG72iRQL2/kdXdm1D8d1Yb24QDZ9F7pA0z91jdl8J6
J6hrSmtZUYWg76PvOSqe7ra89PVWigIfN3BaD5N56ewsa2ObXzcnH+nkc7oAZ0Yq
Hyz5xSWYTcIbZtWkq3H+y7yqQ7Vvyk/uUT2iKNS5rKJ297a0THIveRZo/lj42Ts6
jkLc+CYA1MtgoBd1875UIbuyudw6vihlV6Al9swEQBbDN9DAOHVjak92fCt8CEtN
EX0ZBKHHcQiIzDwPGNs+VfLZg0nKxe91h6UhyYcJ5StNOFDdz8ryu5jg2vrSwF4y
Bd0uLqTThlZTEUjxKPpID2vHwEmEeoB0U43MGNS3fsq4w64dus5GtR8P56nEX1QY
QHh5bygs8xBBWUxv6KdtWOUXR4LyXdbgg+2i/OCA5mOWTu/fnoN54ARw2MCjmbnr
eNYCO2h/xTDXWsfKSvE2fG7VTAyXO5Q8S5S3bNZ8qJguA10gG3SXEvzh3m5Ych+Q
vEl7N5KGfMtCooTbtPzJ2UtTwH/vt4u6uxipMfuL5X0PSBKPraUqb+ryjS5M14jl
G2mDvok6q7NoBeN2zgN3xwI9EzMUO0hvjphJZAE6as6LsRGMqW0r7cCbG5A4kAls
0g/DXb9ZjJSBsUuOtIWrmzII0XbM0U3/5z8+2R5s20GRCWUtmBJXq8yQmaAxcd/0
SH9vRU3lRfGZyr89ctosKwg/+C6H7/xU0gXhmLgMcMx71oojXTsOpCW/ihoJvHs/
IA8m3YAbL8TifcGtD0mxPzpyBnGodoSTM+8PftV/AOEUR34F+tvSAcfT/8ECdIvc
MsmJ6+XDhSrsh/fzc0lcflafYUpQLqql6hNyU5ztXQG9eu9FSw16pn6D5CCF/GIW
vB7rGEehsD93BpecuqBcaBxz1pk6L2sFiqwfr0vC7tikDsAaltwvFl8lbhOaizbW
4B2DEhhPtgDWhhfNxoRSOXePc+ADY+MbwUmNRvSRD3mm+jcFz0dbi3Bm6rRXwx87
gEOJbwTe59sEY+otb/Qq+4CbJGFE28rUtVUf7DdPnuVTRUnZ9JTjtPhhsBvyhZbn
28ctPoyx1ZzS3DlzY8TbQI3hf5SuOLsEGj0KpGkeIFRfPlqg9GQSuc5e3nosXx+X
bWEO7rtg3GJAU+sEVxoo9ZU1t0EoymFXRcn2jzm3s7n3LS2nWS2FY8N3rAkWlQJj
bKUrOjq3c/xwezgM6SjzSB7beKQZFd304L8mmzS5/hqjB4UnB9eWIPgJoDo+Eafx
rDdgRwAGMBTIlQjH/I+IS9iceqzy5VP8WHpABIn4rENddnre9YXRto6wt0VAsZWV
3FqlXLbwJMfcyIEyfomgqwvLuDsqwqXhX8f3XHXRnKWeShKMq6UPbGU28T+poRRF
7wXXJ+zgJO4y2i1VCvsI35zUgPBDSqJyUFGgqFrYntKlzHAD27Ubw5CG5IwkZGKb
L3lgcUQL7QcyriD7ImGILsdINS20W/hRffGLJoWskDpaQ1/SSAw4sO7IGOjsE5OE
4wY8xQntaPDoYTl8Sco86UI7cu0DNOuGGUprjiksjDoPEZQ6hf5+4kwvOm/wX/lv
Qo+a5CuGBAsTWVpzHL8hSDowGzmrMfAbHtS9+S1003j386ktyXrTWKdn6N719TlU
1lj2m4p9kOzs5mA6x5rpW1Ok0M5rBTEdNrKJZWj5aycVnI0lht2GqIJi8A6z/+r2
QGoKkN/DLugxX/rqTywlHIK4OSRcjQ/cNCB+owbm2Ij98b4LFKUb21B4z8YfdfSc
U+VKMPSYM4D5jAe7MLxyMsrytoduTLftKMg2vgBGR/SKIDLeJSCKov3nYFju7pAq
+ikZD/p+nm5/Ebnf/fKYImAaYB2JlWf2Uk1hx4q175aOwkpgakvU4Onl4TE65d8O
2ZYqNQNwgOyOZR/X/eRjNPgo/CMH3bJE9UM/HcaFiC/c8418zOkTBHm6ksX+/bNT
qSLtUVQ0dH3Q5FvwPcewkgUh6UTQD6GfiT6PcoUAEB3dpPBo59WgNbo5S/A3avag
qj8I2Q8nhgTIRYAR3q1kZxNUfuTFGX/gWGTXaDQGmvGc7lGBJG0kOxMPaamg8l0L
z5EiJ4PUD9rNnHozTuv2aUT2cQPqjgV+ZTlRV9yFcnEFLSksL0aOPKJOJvUjKXKK
uLX+bkYObyQIpEJ6oSboPLJ7SB18Ba5RjrYG9eaGUrT6R196sYt/19crg7qUqtbK
y4oZEAclXzpbQBwIyAUVEcqolInHCJjK90vas3asEW8bTUh9dniFtKPe8WYf/4E7
HnSPLPhn+pwlAPQRqiiyr7KWOQ4YjH+hB5d7ck3+S4+n+D1IwdmdrKmvh0NvtoEO
8gboV37P+/vwbCc6/cgTiYWKBZ/lj1Krj+26rCD5SAJGokOIB7bxEMRQbfNuPZ7U
Urpppc5n4j2STiZshtBxAjEgtuJg+2qJZX3YR783axNppZmUJenntRUQq6JqkgGP
bDtzJbbzWhoFPuAqBFnyCgMEP4BGzYtYKgprzmAr3Mv8gJ0I35fx+UxorJ/cacP2
fdze0FYcQr4zOmVF76WdIjf0zPn8Ps6h4yCtq+hunhClu824N2U0IcMAB44130s6
Z2ltRBFG0JjSyQLKnpitUViKghieLAlCPjazLBuiPR8N0nq2+jiqszRBJZouaX8v
02Z9F+xGPI5n+j0DWplIdW6Sg/0fbD/Xg9xgFUq4PfwJMsDSSK/VUs2FHfwq0AcZ
nc6wiHik0/dBxDfmryBPkrK0V4lUN0GNuVROYJxjh/UQL5xuSoiXCB/kaVGfxNT5
QrhBJVliYqyW9q1x+yFWgKSu7vjaIEXZDQwyl4+6GnadsAJNVVfFrJ8ICahCLqgL
bIErAXj0pC/wICafVJR7z298JVDXJ3cThr1mG8BE0QfRHF5RYnheof38Nw0Vanuo
VeOOXKD3nkfkE4hakDnYJ2eHzWE8+3PcYWvLzxrBWx9a8ki/MI0jHDJb7hBL451L
PfSqd7Ulf0K/nWbFduUJzldhn94vfpp7Yu0Wo1zqF+5u2o6fKw0mZK2BKLJNjHns
yyM+4gH0ystbd/n6ufqIxsLNoOwM1lhn0U0KY6EweqgBnfOnxWjjL20I81k8sqVW
WzW+A3PB/mkzihLzaUYFSuGhx346N5ua8VXo3MdxMBAAnQ5MeVlFrPZxI5Kz63Cp
JX6SFlAoVkpCn+OfI/vXQr6xyQZcEZlo4K44GM9VknF43zt5ZjMKK26hL4X3cPVQ
WC5+CS48qGl9KriHCcb8qfWys+SqYkg1Y4e6W41BUXCPT5UNUl+G8TqSN8iqSuBH
Hb435wUm0lO1yyg5p0WB/NYp/T9ZBgq3Xs2NzW0O2RZDPQZJatC9OCO99Q0xIjau
Crcek9ucYUf+iO7yCXcpYGI2Ij9JzI2fcXDkxh/pcrx5EcXQuKjrWx9z3YEeznN4
T/ZF59zORMbGn57569nUV64ixOm1GHj9SewloGZ/Wm88a6T8LmxWBxubrcmbotbV
JAygWHdcbwYeqbH/fYR6pGhj0uGFb5K/db7J0l+aAJdfyr89m0BVfnwg1DeGUXDK
huzf4ooU+Y6nYtTaobBdwB5kSWj/gAQFckEgGa/VuVBDZOH8tsaE95IKryDKSa6h
9JrJC3aDKzkLGFpIN8lUyW4YbUPfB2hTJhUa7c1QIU9TiggSNsx2QJrJF3VUQ3pr
7I7YPrzDV04A5Y8CxIGsL6lIYYZRtJlp0NOZ2Ga2hdghDL0DJUJz6GQxER6atwb6
VXSN9cZVVvnT/KIroxwOKE5/QD0Pv9DTLRLJUQegOQw4I+nTcOc/fmHaC6cfITNj
mqHLFT5CUaMjasJjDWVrMUyJ2tPg8dxlWdiKuustzCklkywSEFlkPEy5XgtjjGoF
mpvuI15xS6qSlluEtat+Y+LqsmnzuRJtj3Ii/Fjgffu4cMERALH985DshCr0xpFz
bztnsoZ0G1anZr2yKDXCuAlscIROph6FAyw9CQwjzUpyQYO6sIEvUAxGUNilsqIq
igDqshd6SMZ+4Hrkgx2aCofhJAVKFZsP3JBdxg+Djixg1Q+J8fQ7emqJljfTc8u9
afuNxPzkBfvxsm5ujw1QKDKbQdRiPWigB5nMUdauzd3ooVyvmZIEhJ8GbdqGkBz3
RBKFyXodJlGJjL/QabQhl/iWDpjGY1n74s50ikB/61vRRJnhlcDCaRlyuPSkkln8
p8iTW6lppq2q/735vHxF8AmzYBGF91Ek3bloJcCF8HYxF5T84pV6KPcn5ZrXijc8
bhm15AbE7L64t2jCjk3QesYnJK15+CnqvCKuJNb3SPdHqogSbROrA/jQ+FLJ/tro
HwClXiGRlIYK/JVuC9IDy29ZnHmTcHxaBxvhjzXkjJVothQbmCBNikZCcpszIuvu
Ka1sOwaYnrUjeYt9d9koU2Z9e6eiJxn+izvO1ALZ59qCNDUOl6RpehrwKdVdliWz
poAdCZzRGsNFVvWU64jFq/J5xD58vKkH/+HyWF1MUbYuJPU9y6RGwTSHVS0IAtqX
Hap2KZM36GvcVZ5qkbaIPRwYG7bKTwtnEay2FqaVqJ4zjFL1PgmkVD3zBKWuuppq
mWXAO4KUwvCAQTp+ISTBeFXcVYzbxV7svfM/TyTNcMaAb9YJj0c3kjl6Hxu3NLra
hOZXbdf+XopbTusEvVckfpK2B8Al6e7Jl8aWpIc3O//K4veRkVBuKbdaEeD6qyDr
HtjpCmF3O5Sl1B5nHyZDp8AvIp+G20C3fr4DvDx95ic8PQSJTnzhKbEGfe19q7E1
L3onuuiZHH6jTe44GKrvpmb8epb27JTn+QmU+bc0/JSic9k3VYUwRRIwoJn9L57V
cREkzA2bLKCDAH2KNDf1acxIvCX7FDUWbxsppfUcyTBE957cOXmUwjj2pLuPeqWL
kEFK4LEb84FHwQl9f4w6kPzLyqrfuLpn2tcylqMIEJxhS+IHza96nD2FWQxS3df7
hzYPSZCHWI+KSlhXxCOH/t8g77jRKIHogSEsPbv78Oq28p1Fgv+/iCRdI83JuZ+p
9W9ZIbB/N8PHXNAf5K5dyCIJ44RfeN6l8/hAUejeypH1ZY0pXrCV7yRWrOamWVai
wsFje8/LCe7kUHev5faQm2tP5EdqKs3tHQqGNP8wKkc1LDlnwOosI57v9/ozs+5S
y1gMJdpVLqtFRHDOUK+UoFc/LphntHczcIdyOTDTA76bM2vUgBgkT5QXY3EMH9YN
eScKFC3KoiaZlSFWEeAcBDvw1kTWOuP3qqidDRZ7uMf4oLQEB0vrEVtzp3vxaIiD
Dcy6vVX+EZchwYgFgUiJIBbGMPY6nhVX98I1ijfBUj8idbJA40/xuhHMqa1IfiOn
faqWrEDh9GA4DtNJ8nPvL5djhiG+OjIFPnxI0aUSsXuZs/RQq/GHWIDlab5/azTB
5xj1LY5AfRyrr5cadEv6SyQgDS5Pr1E/sdK4Tb7B2Qo1xOsV4MV9K99GbA0MDx6J
BEnTWOiOTXGwyve+1U64H7KeJGskj054bu3eog3pZRRnpoam0IJfFTwEEB5eY7hW
CAh7D+onyWM4O2z1u2EQ3FVP45u3eH/FyPgEUjIYanPCwx8GlyLLeL6tqAzY5lKF
X6/S5n9tt5MLSOb/ldtVNBN3/r3gffsXdHBGPcZnEA32FtCCXDo6GtlqiMQT+of2
iSwJk1N9bodiQ0GQQAzHuyN6F8R4bSG5mLJP+9gKThaMNQAxnWpUf7Is63+hksnc
w38dAtJUpCGNQwuGvUt9UDcS5rftUl/osMP1wMBS/PoOH11S94rWiCjTrt4vqf69
51OOibkxO3Qs+OUI6vHhZ1/iso72Hjt7C/S5UQrMg7pitaa0KaKbTLSsQlLifp2Q
iPMtI416jMBzZjbW6cyQjNDvx1v1iSv6s8UhzVrtA4JNDG5drxtCULtpdMW2Q1S9
4AOH0l/BC/U2qZqnZ/f5OVNvdKqLbV9JPzLvgFTveXj3ZV5M3fFdVSD3OGpuCm2d
MPgsPedpHozmetsAwg67Yckr+tZjNaKANRWdWxG0e+phJdupWxxRKR1Fc6CAxsiB
AbHdTsa22ZD6FvAqHldkU18ijzQcYQtvGzaTdfP2kmawVIcnIczSJ3F0iAl28vYL
THNDGYRAvaj4aVbMNZ+gnaei7KgNS0avbreBoe2MtemJ393JXHo7fg2gjwCVMXsY
1NgYDY8wKygzgtj9bufCtMozkyc3DxedynrjE1lSQtn6G1eensBM28usVVW3XAUL
XFq+cIEl4Jiq1w3eo0dnat2eHHPPqeKuVDQHk06kY4D/21CSHJ5nplPC3alF3xLf
Cuv8MrgXpbPGFoeRWFXuO7NfbRQVlUHg5hCIwZHStY/OpxM7G3w9oznbmgMSmJ/0
m0vB+7ep5IrV9WJwDjHzlBJzgLubWe0xAf51A3N3nQeLGHy5bqwhUTFvT+bHoTII
oU2mtvwoYtFTR9UndPqU3nGqcGWylLLur9Yama30pOMyHKpiovrqv/Co6+o6xuky
p/+OZT5/uSAMPzyIwy1WNMT4kQykw8rf9mC9bJMdoyrKqFpFEBf7Az8qo438FQyx
ijqmRAUYe9IWK9XvdYqQnCz6zkMNQ4kBNUfqzOR2EytX1f8bbdCPYvAhdGqLiF70
N/5VZB1q9d4viLOSZDAC6DaHY+rzEQEfl2VC82+fLq9PVB9JOyHlJhPQCLvH3K8P
JMd1V29VHkb/1S1wNc3B3M2Yy4rFkH7jte+KWRA5EfXn/xwFl58+SPf/dMA0lDi1
C/rrQnSRlawFGyeLl8ezPi0QdFgHmMjUvFJRygVgfwK1nnyuNBP9fzyDK4uyKTYK
d2lgZIVSX0YFYzJnbqUK1Y4kebwYF4QlDZLqrwHRsmd1X5cAu6pjJGF6UCbAk4tm
8Vs+TFMM7797vEezC3sRecEMk6RTofs+a+CRw3C+bYHRv+OQwYrAGFazx0mCRPla
X+EeaxN0hTlKPEcQYCnt0md3rHd5QRCZQfGmRbBRO9assgSm5AhUqVVCOZob7nys
lpvr/mujB0io9i1QWw5L/SJG3W3At6gNtXe5IAyZGPz0mTFptmOtMLBiDEMIdQwr
raORgK23UUEfzvN6py2U+rZz8ZY9dUKTE9eJ/YxYDvb4EpwsPwsgd359J8WELTDp
GTOq/fvsBcJ/DPN3WwMOMO74e0urPLQnEUKUmjJ1VKikH6DMmCBiXZRrcAHYkv8D
Q96gcBCCAdrw3XbTcGSxxIjvWH9XzPbOjAj3c6duPyD+Jljj/4jnQrG/SVpYWglI
Pidpx2behosCv5s0FFawNsqtNaVDLiz9BNGzHqGIIGvA3T1IEbilkjYr9MS56BoL
Sv9eDNa72GO7cg3N4CwtS5htgtozh4+ULt3m5/wGJ+vzNANd1XNBgL4Tn/rbJoSA
36GKVRadPifJP4bwLaV6rAJlAdh8q3SNDWdQCD6MMun80AsXpu7a1l91891+1ShR
H1sUE9p9mWs650pgsmEogKLpx4CPtbGm7VL2BkDkKQCAAnFQTsrmAXM6W6eF9Ptk
ChhtVMNHo3qbruKOsFP7fGo/81ZiOpYK7HaU8u3TGqWwu6fr/zPtfoXbp7ISsomx
kODaAwLYAwW72tW1FlxAWzRqKooBmmZiakPfONuVWcD4XABhLkHU9pShKa4Wq5Ge
xjGWiVVZKwbCZ5dzZExSibhD2zcpujbh5c+ri23sjePvysH9kYwqPqF07B3ITNLh
60ydiCn5xZyr3eItHq+ZylCYpTRyteJuY1OmqX18jWQK2IQu95KB0hJQ91Z/oMpV
hPYN9AFzjn424eYjIgqXYVLs9qxm6lGHKzl7KVuRvxRWzgY8r7QvRWGP/DEd9RlV
XiiwXrp7LTP8XiIcZ6J8zsezvzw9+VsoB2eGghRqNPWIsRkcrSvULlbO9d1sU6vh
QrCrAtWEOzvH/bwaFFFfUM26g2imcr4V6vgbepPn5CkplESDVd46tfbgdRs4FMY4
DRrybc7CxRMQFVcCexhGa0BUCrPpDktt83vP6KHpH5B5pwxkskXKfspQg/96bVLR
NoUJT8FKgxncNtz+1wiwBrEEWNG3CxiWzliM3Fsts5pBlLuKWPtxgENuDOYs44MQ
EIyJjV84rhZrBwmfnDIYxcpfNF3FgJb+uECsF4ESwVFUZ09Jq2aFgWguJnMe87NT
cx5r4lwkBROixg9hKIep2hbAeAWkR/6jGWgKmncGDt/2eU4MBTFz+5NeW/Zdvtkm
CfuJ+9+/rGKkoi1nPIQpyoZ3qTbe/gbnczTpXjUPSx8C12ZLNbO6oAt/gcx7/6VN
GV5/aYDGrEVitNhsZAOcVCBttBBaAnOgcf7vpwm1Mq4JDDkVjdqDsHQxkww4X9ei
gGarTOurpFWhPB9uZ7SrRu3+XHq+x3Vn0mzsAUQopRjygm5OR62nPVvXA1DfKehL
Ra0+DOvf5buL2APQCf7cYKHSjGGH9HLB2/1un8lShzJ8/+KIAaDSZpvMgFhoqNAy
6CVANYChPgOQfYiZcxOQb2uhl+jNJYVYOxSyGpzPhNaAbLJIgVTxUobn1Uxiif51
ppCFEP8ySxOiJ27jY9yNJpSnsK0OYl1Ot1QCeMsGfeKXaWnz1SpR9HzKMO1HlPHf
EiZNg6azAkeIP5zOSjG2d0KEt+9zzEPRxkNEsh//HFcYT73W531xlu28oKXFMgbL
/WkhRyu3o9TH0jXuVxrxJ7RJUitlac0RKBXO6Rkm3sOvRrwvYiOiQ0o93WlHyjkJ
bW5PnA4XYkiC3rYvCyerRB4hhhGKXHOxoK3NW/+y1tFtKpTipYiJJFh1BZitbF3r
lWqCtTAKqcSf9bmX7FmcwgZCF4bUkLgTD9ARUKRroazSd0OCoiSfypFboA+QQJY6
hONSU73eh/IN0RvR9fujfs89DrDuMtGcYTrkeOhjHqPRZrhJIzlljg3CorFuStlI
3cd0iFQiLdojzbFFdizU9yVs3JhtuW+OkRKnqsHxRrhHQM+5+QAfo5CenvF04FDn
+9dQ0ElexzFs7utKoxQdVlMlj340MytfyNQyZxFfpJ5N1gnKdaGRaz1KBzMIlLvk
MAYOxjNcKDWkFFtRJAn38AbvDz2LmNJ2JZHHOXWhUBjcaIukDPtn1BLTeSmWR3Bt
3DQJItgkypMY27+hwOCG9g3knDxxb9ma/9D2EPGmjzC1D3+TOsVGAX6okUTWDPCQ
meLkt98CHPl8PRL9HYnVIAMO+ko5Yv2n2YYk2HIZobtaAV/x4mn+x96qE6XXX9t4
EeSCuNU8d+Cf1WnWN9d1fx0qzkkQ1XUnR0FfbTmxlG1oZQ3KNJQ/hkbOhQ17lnc8
YeTj2ddTIaESl0aeKGKyGuvheOMQlKyDi14dIvpeUH4cNTy6mTzX+8dEz4bz71bH
c3Go2npq455N/SE4hHlaYWDMPPwNh4IAkEjZVwzAqgVZ1NslGY6xc0MPlW/fE+9A
9QQRAo9gMky9D655c9aGhoSOHnFXfgi6FwBBez2xu3UPW5KyrCBDLPEt1jb+/+kd
YJJRDyVnFeS4dMFqesYHz1Xd/bdQ8K8Cj1QU3gQnoNC+Mkatk5J/SJPUEZS6ECAq
nYo7FGRg9OZQ/49YM85b1bIprhk5L46kK5EYIIw48XThdlbnPpSi04TmYB736v+6
vkHwpgO2ZfH60hjWDC8Gb26abvQhSloUNtVTCE6cSOrXtcqM13VcnLHm8xs7kYuM
aIPS0W0+mu0pCcn12n6iGCDzeHnTTlTsS407jlyFBAVfbXwU9J9a0JS+KbEw7zNd
tRqPU4a+rt9Q4D0ZARJQInGP9XXGyK9758ZdNdsVIYjgL1wRBeS89NcMpAyyVNwR
jb3r22Moo9YkcvsVk2ABMbCPAk9oHFcDva774CBqvTw/v+aslWqJ6ztOhdbN/CbV
c5Ck/ONeWhed9jUEJLpDJCyANxkF7Bg8Y6N59FHfxiWzrwdU40gL1bbTeiAnWYVE
I2hQGcNaaXrCb0MUahmeGe4WfYssxq3QvEieQRQ0ULbrgoQlRrL4M63ijSy5es94
MhmfSybBmd+I0iTmr1SxFmS349bB++z9NPOdEPOkqNs+qPrF99VUNhGgmZfMMhai
p2jSo7NrOp1dk/U2cfYDxkUSJKhRl1qxHv3NkAkUJUQjsDiJny513Y7q415RJAbQ
HSscXGBLomyvc5xTH+dNcqeVN67Y+nWYouE/YvznCywi+IDc79gofVeWpb8hlRxn
mkFtKyLIqBK9VdM3o+n5Ka4PoAHOlj6Adk3oWznsFy6/WPXv+Oa2pwPBM2pJG6JX
LUyufCAqRBCCSQMQdxlqH6oamREwyDqJn/d8fDvVwCuj/YDPuh50NNklj2rq/8ob
NQ98yh2RDfnd+DXMoC+EsjfJ0aA+QTszww33IYTRDGoIbJ5c5406l5/5hHhAXXSp
ET7Iccev2mM1CFyW/lAEjYacMIPO2Yh2ToszUc02x4Yh6YZ/S0qDFurHiFe8S+1U
N6biNXDmiava0xIfwmzo5dzmhZVv9hcGEQPEq22V31G+MoeKS5pRlj0+LKULvXhr
4L/jEtF3Zk10F/XvTvcnG1LXXfXdtjG6FqP4W3ODo7eNrtsUrscd3qx53hDg/2zy
4HMjGsT5ImDKYhtO0x8MLUa2Ap36zZzlQ2nBZSNnlYXKbl7GEvOyrrkhRZgngGsB
vFHpVUoDXco8wbx4ydwMhzKc3XDQ1xOEp9NiCW5acSP+Q7xotyWxPJM8QUgYjy0v
AUUlDwj5N+Sp3tAtB8ObLfK0cmJlIz+j0nXg0ZHHTRlQOB8DeCDffSt1Dvrkz5Ml
M+cvBF/U01gpDg/ZydBZ1BYXcB4OncR2j3K3o67sbJCLRZSwbEgT8/EqXGrN4rBS
jvE8B3kgeqThBHHZz6HNHsYUNqlxI5HHikrmRtYVB/xyeJBwcuU6lPNOLQgiMXm7
67TrL0de5su7XAheXaD6ivIdXXUA0pd5jnOI8aIYpm1M6xjmqHCxxc5ZZJRjdZ8A
GBH0cUOqSvEaU0iA3zD6+5igec88IAhNHhA61NTHJGOZK9pwlATie/nuIezPviFQ
bVHYMeO7umMfs/6cdfaK3IUmgWcU+1K2Ih3XRy0gjvDyNLo5zYdQV6/CdeOoCzNc
/tnouczlV9S7SkJqXjggtf/sT+//0CvR+1oyykPC7aT5Cf41kkALrJL+8Itgf7Ji
fTIq0NLQt9P2lRq/Qy00b+erGmupDTTJhYfp4MQufzOu/DiFF7/D9qny+DMuKhxY
tWrxwXmaqB0mq3C8EMINao92Xlyvtxvq7ijjHcas1qrRUoABaUw2BkULyQNH5g0P
de5or+GpT13LoKwzbSw7mHhOFrqWMu7yAVh0+CSQVY1eFSnK41k1fGQBUkzI7vgM
ha2wt0h0i5UeQXirH32bMDCGnP2B11jOcqqEuE41EbnXXD96/Lx4cJeXqZEWzRWl
L3EhrqOJ3Hj4AU+cgCrt1EbAIw6zu2jHJ25keIsDFCxSGkPMtUL2h2Wl0R6eE1fl
f8aE+OBulRlKeCXHSen9tc3lcK+Yvsunaz/Ssh6hKgM3KSFLt2BKCIJ2nCm+4ytN
BKalz8EuChsE4sX3xXDR0hPvdq6+llYsEvmEolx43Cy/mMl8HZ+re/PxZSgPhwN0
y+u3w3tiR8+/bLgPRaUUWJl0MHs8h1BkY3lb+tIk6/CT9SbQ1gkryoINoj1oN28F
es3HniOvxSU7ztn1oY4dGP/Tlkrkbe5MhuSr9iA2RLFH6hN+wL3aA79BkTGsAQkW
0hEzF0/Y8R2yRrf/Bo4rXVCHwNvdu8S3SP+HxmdBX1DgoM+uc7V3vsEUIBQfIwIY
6zoa13MjBXJ5NlEogQ1mS+bZj1iFF+P/Md9VTHcdoh/6XU/oPg3dvuFroVW12fUR
bez2/ikbCZOOSYBxC1uuQjCqgG2lOTERddOkBPNw4ZqI4BW1LZXAvSxQ0Z/8SxTZ
AF0qJZVPDjWHpyLztPMwEIA+6ZpOknSxf8tmoqTIGMLhlOO6B/P93p9SDEg9IVI0
WDBgVFA7CR87xPsW1psH5XZo5KK1K+iiNOPVHqednASmSS+8xbimheBPwqL4GdCy
69DTmZbL2RZzvnNdkZl4GxVG6j91gBoAvaRTomXOST7uy4hv+bRD4dghZu1yaJpE
FUzVej5BRJgtIs2oq56FK78oy5I9aRzOKtnTq3YoxkfuJe6H3d3lrTNXmTj4fH9d
MzfOs/o7EPc9w9BeLFCcPvVooCmb/SxcRdBuT+vxugO17cYORAgGMVlwOOZ6XBPr
he6BPgcW2R2yH5sMb9vWWAbxEnTw1ZPJZQC5ysj4ICy8Ct22gr+Miqjb40m7F75v
HFPlpK+wnZW437UiPcSf0xc0x5wwchVrmXM5mC2Tk+gxNZLghW8YHXiOVe8CuIbf
ZYZLC0zirILV5QWZRj/wV6d0ydrz8KyknaNKae0Ao0ycogYgrWX5VN6JqL0+w1+Y
4EVpWIVni+lQTXleQUs7rZHf3khmhQLDceYe4GHdF+9gjNnCnK/9jBDHn91alMjV
NKS8XFUBiBOt7WAylyziP0XIU6T7sJl61zgEU0sruoC9+ZrZztMyusOQ8nhDWTzJ
DQqjCoyb4l1R9R/1/3nFxlc9o4OA7TCvLgfDXvPX7QUNi55zapcKS3KCGKl/2QHb
Qxi+IoHk2rh0ED7t49IuLzFdSXIY8vRGsO8Vut1E3gJKYPJfeoQYVBYvoD41CT8O
xkOb8Ug23/0dELA0gdEcr7efvbIS2tNFUf+x69SQIfdOL8t+6fAmtikLNaOVzhaS
c+NjptLuEMJmA11KwrhYORqzf7cbP7CXx9zBjvKcOEkTBzk3ey/U4yjdybksl1J3
JwdvJ2xvUhniuLgcUzBAe59z0ehKL+gOgHpxr6RE28Wx3G3XdqMRiOpLqoSKgKEd
eOUiaa0nH1SDeY8rw01CeICb/3vAr2CMxTEYvctO7QAyRETo5P1UjgLpPDB21zcB
6bJQbuUQ5z+wX0NtsLG/sDTuBN6m6TccqbH2G36jFNWH1WdMbuKgp7MIoEDV5wM4
x724n82i7PI29OESReHWMrWzNWj4Z7duUuVyRjfqbwppTgg9GaxtyehVAY6OCyFS
jJWGu440wL2eJ46LHgqIJP7P9zCwd8SciOiM53Ib+tKNHhq/MXdeiwIlCRdAoKAw
YuO+kyulCHd1i70pS3M9Z73bVfLK1cxutd0oVUOOH+n+in/mySmqCmqwfsKAanaG
5BUvE9CPuHC6nCbjeNYwRqg7hjYMwHMUfU0LFuncP+ttjbT+gfbIgZAkYj/khv3z
fnY5FUfPKb/iDEJdOj0hw2MLbgd4+MqWFfSQTJrMX5UPPHjPXkA43jv/wKPrM5qo
5m3VPn1kattR+MykI/MY5hAErRX9zA5Hp6EzHrZcvd0K0MZjfNEIwnubr2A6IL/a
wzFMco2vBN53MQbd6sG3jFQvsVl663L8cdbJrPwZ8zZ7THX6apf+S51vCAPQtYhm
6a8bEDzjchePoS4wZUMHuigBuo+fKPe1xJiI/CXNjglEDuF9s+5v2D4tPlxGJUNP
a2+Z+9dB7oCGltrhz09CJsb3RqcjPwcOKN+3ptwAqdTlxCDaJdWIUmv9ChnWzDW2
KrrNpwZ6GFMZs1nbzpT3lbMnGmL3qzjVe3OAUHYKT0Gy+hNEhf4d7GWFmRDE8SAd
NcfUSLXFOGXDJMuJqOUQDe81LPM8fRL6+U9hA/LyABUG/2L2oXOv4GDl0hbOP0Sd
wGutB2ychkybrmXJ3XsVVFIeabtSUxfHkgnIaXENZZJiiyOrdveHKYCTeaRFU4LD
3bjVMo2rAxnpd5JfzCsgdCP4sb/hL322mC3VP9S7KWy+2ujPXHvbvpCwv/PGq7vf
1znL7pooDzUkg89Nh+BOMpB9r9OCAGNzEwMiNwiBxFpo3Hp6U9M6pnyZnPVUycd6
Jg+vR+RedPEdNAzTA81+O3SJf2AUz02KAk1f0RY+KXftMUGDkJRnDQbbE0Jaax28
IpLJpbW46jVj5kxSujNAwPPAsx7ubJDsGlZT59PnDhtIl+rHxo6ZrEYQQyBWUtwu
auPc90XKvYqfAhtO5WWYaDyFi4pT9kaQDSoUcm/mkQ8moiza7uvL3Ego4rFha5l/
bcUg3/yGSLMA3XWejXm1REPXlRpMBuhDYEjdsokOSbUGbyeXXUwpXTPMR96U82+U
2J5aFElP1bqiGajfyh4G/eu4ioiwWJ+QHdysOQZjIcm629ae5dQJ4SYjk+PTH5mw
A5U9F5ZlAaaJqE/yvMJ17vGPRNpYG804vVpLSncDImXO5+Dz9NEvye2aYMPRf12j
RSuxBQ0d4v+L6Emi7Scm9A9Gfc7M1GFuT6WYYLKCuWzSnGjAZxf+DzXf9MhMzodw
xFzPTjnvXZaGiPhUOkmR/STBXtP1IU97k+TXo+Tq1y3iJWol3fJbuFc1EWqpq0KG
49yc99tjC32+lRuIDCtV4VtHs9omhxfTdqRrnGMiiUAmqxYqgjHuQqe+R/G6ZJoH
N8DXP42irG07Ig3KJc9kW3F2IXFZABmm6lhflbgIoQq0505878Dz3eB7pz0sAOZD
bzs/7g+myQI+eG6WIP+FOhSOS/ZombGOWeVG90AxOd6AG1rOETE8IofuEkl5qfG/
L50y9VI2vO2KQXUmNnBIIIzc7L28JRpIq0ZCXz8tmRY/VfS104r0iPo7728b7L/L
gB+bV3BvHRlnekOORJ9gCeQGRvlvsDj0PyMflrFTIFyNKBl3eDXwUnTDlCxFowZR
c6Kg39U9e5UDs6JIsL5+lV1nHo/sagDF1V8+Qi0rL7JvNOC813CGzgIFcTRwOkcF
8fGrnzzwW4ttJ1h+D9ZrLJsZoUQnqAsdJlqpgft0fA3SQlsDza0P1hk60DH+lzDq
dbFCne0/1XqI+8THHxpJGDGAUDaEckV0mVgalf7QrrTTLL87BcXGK1kYBUbvFa+O
Q1UqjvQcpjF/Jkd3blDxW0ojRqEljmiv9V5wDj/qO8ytSpGVSt0CT4jcYvbS9u1D
fY3QJfqrBK/XSFhIad6n5006osOZuUrZdsGnE/sgXK/DeJNAgfh5HUJfRWFm+cUa
sQ2Xv9F2VLdac7C7xrqqf86dpLeiApG9Oxi8atW7pl7V+G0tEJLWTktSRVzMdGm5
csZAgD1NMM71wyaqmq+rG0McY2s0vHhDj1P1B8zVTJ8ujATFPMTv4wZowIODAL68
0jAjHXFr2fo7C5GA6kZjl2BTAj74qvwyr7AftEfuwYS813xOfl5+9nWdyCzHl+H2
o1+8GNPpG+L2mKdtXgyCZt8V962ABAt4fD1QuslJm1Cd0N/VS5pbrBnaKKg5JCDj
/wxsKZkZHVYga1gQak0BzyEhH6pzRqsMkW8mR4MOrMbGBXOuLAeSjvfvuYFgEALg
UEoybSLjmsIdjp3LQHd3Na1sR5Lz3Du3jy6Iwr4cWYq9jThEGC2ThljayFy7v6YX
V5ZVB/2JY8UHr1ykZ7tLMu2JyywiLKsIuIYG1AE2XKwZEuyPPDT4CS0ucL8ePYeP
n44QUYrdGXF6BcWVnbQtHkZJfTNdoJfokE7gKrWhndtQNbgGcKQlloKpkjBoJZQn
mSxka0+llzYhah/+hR6N4ZNviqTZTub+ff/juUAL40dKtktBxlu6uZXgwsQkdOrl
ZBtyOY10T2IvHbgbNV8ztkSy4hfb2PUUvFSHZtj8M3BWw93FqzuTg+Hy1+xp1cgz
N/FGNZfdOxpwJBjv/GPx7cwHjAsu2/tbFbsvzvTm+LY4ppP3i5m9pMta2/WUoPZL
wF5U6HMXd7ei8uTmnFV7sKO3PMprkXIPtymlphG5kyes9wAaxsD8exE3cf23Vs1b
QamhAetPiMDprUxCoj1qx6/qyQaxTNwX9HYRE/wpsZx7Po0AvXbfgGLdMS4zHPRU
mtV2n3zL6dTElU7unr/3XP4n5XFCfBNs1BgJ4BJDzfr7oDeS1S3gpxiKDL811+OY
bidpoo0DS7ZzGoX3JuOz9sUGxpt0CnJQdzV4VoCpO/g7ZRAxOIigjZjwRW7Q/KAD
g4ce823xvsFn5FzTPIaIsyB8c4kZS2NVsxNz06urs2mBlfs+612HybIHc8llWNPe
XeDBjd5JngZpWf2BCo1Ul5bcuOGaTfcrmcAHkcITjFpfT1UtKMjnKzc9L2oYHc7V
DZSUf4RQ5Z8iJuI/NTWQmg9KNyF48zd+dhJIiQrLFyca+4H3f8i07aub8Y1RjbnE
IYQLkZt+E58jkD0zAH0y7Ae77FifPpef7nCqrvmtpS281Y9SQNB57Sx3JBKH7H1P
CCogqdyEsffb6QEL3WKRhUeOEFWAhiwFCoPi90Sow2II+l9LF4We4yFDXZUMDpUd
pcvjbUCCT3X/T4CS6gEhTxDCDvZjH+hXxs/If7scgIILauCxEngHrbl5vtu2um6U
I8V4+O7DHjyYULfUY8TQfwpyBLHydzAgwdqkXZiVVAfYekfBw8Zsd+Fj5DmmuwIN
lkxaQUNAY44t2OnhmbZGGtcRc+JLU7IXTylYYLm7kwCAwME6kJdKvzmOkclnidml
BAm3aZJA4F7zDpazetzWobAdhITZM45jNuIJAR3IEbgQiMjDqChZfWaUq2rZykBo
TiaIgFm65a9xWsM+mDTo+xgHDdQUoJxLNXn2FAI3aSY4UpKDgj7bSE0PNDQPWsnH
bFuAnzsFUsAdtpZd0leai7zjzDlf1+fFADVzIFvgdU1I58OW0cAtYX3/+dKE0m5A
/jFqal53Kk/YfOGES3KWu0n1hjuRrUFSNBfWmlulMqVgh+3FyUqBbvPmFCsty7Ze
Ux88p/ySAgg0Gx/6tUlzFoZKx65nVCNbMFXxIT0OIEzxsXaoQkfh0tUt0WUQujTV
BfMpSthV4MqndAKBoZphK4O8WfCZGvUKEsVCXuqyIbJvxCRxBX/dmqO9++yurOcs
fUoOAwkDyB80UYTmaW5gNWAA2IBsXgkoushUD729mhmWw805ANI7su0Pf6vn0Wxq
1Jr8AHR03mje6hFNC59pSF1QHbD1tNOSVfS5awpJI/SEjdr+UYPFLlO2g2VVrFAZ
Le8KsLCm0BJ4w9UxPGsrBSEeH7DcqtDvrCBDi6epvymPc0BxnOW25L/D1bvVgLUC
hLuGoJl2eAvzQ8REA9rJ8eSWBDQEIzmAJG1sT/gZHsbg3g9GmC1Xf1foX5U7jCbs
W5Fr7Pm7dUbuF9lzqy/LhoUVvRY8lv6fC8lHiex1XX/3MUutyY09EpO1v2BwtmO6
DtA1jiGAaEYSh+OOAmeYEUTEkG/tTAJIwHw/atbd5SCf+RYq9NBvEy42tQehDRql
wrngHAeMWvdZsTKP9O6CLtGmk0Fzzf6FEenOdGh2CI8kuwdOd54Ma9xcZl/6xiTN
vIr4Q/CGm2n7x+xX5KtxGLnh3OMBcP7SHmJNTtxx+8xk/48NKB213fmcGF6BU1f+
WAtis4AnwUayJxaMC1gqfo6xmrnXU0ovuDyJReSRENpc67xXCBOhEHUVyOUWATTr
AsNEwRnZaihdg4SIeAMuw6b3d1xXpldMqaP5aRw3zGu8//67/KfoAbktnqpG9IVY
uSGrMqJ3elcIAC7ucWblCYyShtt+Q/d1E4cdBP0AErqlgwZq4BGNcVZ8Fyp6YP8z
/P+EwfVPuZqdRXYj9F1VQ0xbh8dOdXRjtOriqGewZ6O8r80cmU2RSQtthTEwVtYU
x083BabFICbkjo4VwlsMwotEtovmgTQCrfGrcMSWJCeeAqbRGOAT4A6NSourR6T4
mHqsFbHN+q844MLtR95MfRSPWASx+BaCe2QV971NR8RosAoa5YlxbjFTuHkSQ3WX
dNtcLH2J4zhGz9ayYSd4ub8wgV23np/PklxLLDi1mWy3oO2czHjLaoMB2rPICtS0
5OJjJPixgONArsURyoGS6vqa3ahv0KJvMs5gKjc9pmC5OOoLzyPH106JoR0BYkif
XnTTAqWpL4zGPRrsQXaT078GCT4rTjyCosMkNS/viCakidO3azXG+Yr70VEaTcXA
hC0BoXCD0jdZV8wRTxGXdDIJUsuk/EacLWA9+q0tSwtIaaz6788MEbV4viWUi1bT
XL5apjZDD7XuPADa/fvgYzYyswBafRIsNxiL+EfHC+onOCh0bu3PtTA+6wfONWZ4
RKV+ku8jAsvPUCBRNmkXbU/4HEl5TN/wmZucEdMwINN37eSxnwIULGxbmy7uhtpR
0IXdN2ZKs2H2j1qG1O62Whfgj37iIZ9gYchuyqsjM/1sAHsam3O6+9KGPhi2o42V
y2MkEC2uY9P3XupObWmSAKJQOIvDHamhPah3WEVnb0SgYDhix4yOyPVIiPjkW/Uy
mJRQ/F8y/X/DO7yRnbmNrvqeUhCW8x78PKa3rRqxFOxmJVy7Hqbgz3dV2j1q/xdk
b20fMUiqAmfaFx8mhSBd/qEJGUnyFSiWF3D13i0292HAnopMceHDVDpxfs8qjKxf
/NbR19eEOPfILjAFY0qbB3RYUCM4+aIBjZTGEK4xkxnIHi9Y3q7hOZNwTeEW+Z7D
9GtpjUkGKlBLWmiW9RvXIrjNHpog6QXq6sRCqLE8bss7kbXjZIv0GL0mWH1EiZWX
HihGeCSg1G/PM5AT+k5chaRzuajxL3ydLtvdu9RRkVlK5pSmO68Q1Vai64/XNOPK
QoliKuUxhAPG/U30K7PZqTKQVWg53oUQXwOnnkvCAyLGfc89+54oW1XiEwtI498I
9WFUL5xOEO0OljpD5rvikblgEk+z09xZ7IE8+dLTTp6gpGqjKry786uXgeuS7eoi
BkVz9F3a9MX3sZc6hQJJIay4Eo8V+i7GpOUD6i4gwlK8XJP2YDsEykl57D7hhc7L
xnxlgmWB3QrrRPDlyG8oXv3aFH4yNmMYMSqieGgtOBVaUYO6GBUneDouIQn9hVuG
4Mj7OBZLxRnjSQrVLD1rwBXkx5N4yjwSTPWkkPxK2ZhKjUOrt/z27/k0qQZckXlb
70RGMhLuP7k/Zakbl5hnQLOyPLXweaO1LSYAnZ6YOGA5G34rCV/T4Js1UYiPlx/U
lrOmm5mIuIvQ7eycXqPGpa7RYdk8dOHD8OuarOCgOUoS/o/RHYFOKumo3X3U7ky8
2otwQ3JuB9OTwFVoDFcMsMuwuu+eypb2iGOqGziD62Dwmjw7V/tlJG2mFO3vfAjy
GdMOVFhwP+U4UN42WOSZ9U9Wtll5k/zQjdhzURNvX/loAP62iQ8DHhtAyz8ktWD7
SRiSjwpDDanlcF8/ceOnbdlOHGnUaQE+zdFtWW5+aj2Dkxu4p++rUbCOs5yaTvfB
2VfIM2etXY0XhDHU0aCdICkkCo8VrnynMl/CaCMGDzZXja8jeVn5+I7yFJMiKwrY
gSqRTzsAv1Tg1pK4iTgG3bo6j6OykumzSOU1F8toZURTIOx/swKHrnR0vSSM5BtO
/Mz1n9pMH+7qBCGjsyJKvcr3dYw6jwrTtnzQ+DV5VzoB3itEeeeA5mMMk6o3ices
fgirFn9F3/yaYDqH5ami92bYmFsiFl/aRjM7d66FLvSv27EWV2kduD4COno+mQeh
1g/zYaPE7Wx4kUXET6bowvOBv4MbKGwkvQVLH4k9XdrG430w0I+v5ugy+LGgn42O
47eeISo6byjbVT9F3TapKv+dR4PlFNUyfSQ8EQc1GUf3eqfm51ZSIxkR6w5/fE5S
Ly7whEG1f+E4yArfrDD6J7YuzNpn54YLUXy8dGnNdmYyDaGVwAkhoQQ+M303ucUX
aHgS1BdbuFZQBvPlLzMi/LBcTfFMmhciwBmItlqSjN8dCRDYUDROh6zvcHPOhJ5l
zmIafJe9/QSEgsL3A1nwDbiTdwZi7jk2LK9fzI3QVvq806TycfEbVHcwDarAIuOC
URgKp+6BHlL6V1qqY5sB7LuhVCSIx7+Vt2WJgehaB/xHbMxSsbTO8FgHCBqo7XlL
K/KxpL1Ko6RhNBfZklqnrIkgJOH26Pcgg7/6aZR8cxaBY6+3s3yRvkaC5GoZ+H2e
ANskTO24Ej9FjrHtptCjjGTypaD6KbQahzqUrc5YsWcgnSYeDf5G2N90suiYuWZQ
+2XNE0lwXsY+ui25QrXnO/gT3Wx3AoA8V/Kpl8kPIDEjlOAzY9MhWiHljcx7V3w9
Ltt9+BTq3RISHSvHqkTu3U6UcFpGfLj+8pEdJ6tDxRjoV/yXTYKQrD9uDZJ7FmNv
JEAENdAHo00ysmkM0er75DUD1Z79MCq41mseG8OpwbsOSHcG1UDCWYAwOB+/wqNK
UpNyPhomlgt0VIVslMf3ugE8idNQCuGa5ZfQuY+c143xdUYDL9HaSdE254KxZh57
aLzmeykOqp+2Fef3Z9RS8tZQghk6ej42t7dzsH9uhN8ftVO3EZYSoH5etI3X03e0
8p8Q5q81q3gOkS5LbfWyTHSWOw+6vqEKVSLuG+Uyd5RgabkoPlU6LvBzE1LBcOpz
qOFtKis9nFOzb6Cu7WIkSJ4VMJiN3S+y3Vte4Hie3+G24tN6APPcymX+/lyAE1rZ
HxRpUjlidodxabz4Wr4pBXkZ3TkBNkSBH14YzLywVwvcw4TLqluGhjb3sXtTU5eg
xyhRRwFOegieK1zZvY+/fS3KyTgySSLMS+peXmoD5nA2qU72XGLi1XKN/N4bRfky
pUshg6F8TA6GYygtz0ECjktsukfhD1YSf83ZBqfsJgy6nmRxKZpxB/bAJO+AvOCZ
Oh5sFzXbtpjynzbtWmMbCJ7dShMPf3YavHlUmoxgsI2V/OCgNdvU4xpQFwj7ZJF6
SeFY4hRwkAiEkD3auVF/sJjnTZKUvQoI8GtmaxVepqB2vLfgO35IhbRb4bQUnj8x
wWUASnpir9+r9Fxuk+hOVpt5cQnXpuzfLEV849yEj3jjf4SSktAKmN2iZdbfBnVB
f8qevWWuz+tLZzFO+sKUh9Yzdh2cgh/+6fNx01pW5T4AluF8n/1j7uX5h1rfIxtT
lBVw1SNt3q91rEQKvFYHOqaTxYRxfvXgm3xXcCmDjtbRVHUhmOr1DyihzHzMhXNI
KZZSMaOEs3mL4+Gy7ZdGft4WMd6AmpMjuY/E8d0fYILyM+8ZghDsc/x61dJONejr
c1C/d0W5pWxyJvAdqRdFbV8tID5q3DvPZWB+kTcwSLRJLs2AMhhyWUUmSK8vRTkE
y0REBgKVbV6QrA4o+JK3uzgjWPdsVUVOYmpbKKj+E2Ldjb+lByjIulsxosqUc81x
KtYzSQjCdE31+erx/v2Ko86+Ssv+1Fr2FYa5lVBKHIEVGWq1w0hRXgwFKshRb2F3
h6lMCiy5PeMb9WWkaceMBsIcwKG1loyHVJOz0ISlsyMPLDc7P8PyYUEwZmDbEwrd
SvER57dtsiwUv6xvlqlPqYQDlFsxT/80eGRrjC6lLPEK8XZgauMmVDvC4z7kUVel
RUjTO42KU28jVS8cvfXbmOUd6WC/2e6A0iaDyCPJo0MnJOw3eqA7Fph8nkGVsX3Y
SudpHDVxxwplhGYcaXZmOqDvFvFwN9SQ3HaRjDSuae18sHsjc4EEZCn1eBRVtrVc
1iWm0IPoV0dZObNrSg+aqNwNUrzrs0gsLsQ6ZyFKDu15KP2Jex68mfnmW2zcdD4w
hg4JeioJAAEWHiu8B/XfYncGcVzYrkMk2SUyNWwSjynuTNqNxZViDYaiGr8xRG33
0SkhO77f8qvOsJ+oehqKS97M+oTUHO7XMVZ7TiDaUOBCdij7YtTfoVS5CV2+ail0
uh6ssPXiv05tgdVs6dVasuMrO1NlE+kIN+VAj/ZpgMl6SdczmPJL3/p41K6bBxoI
xfexwyhaYvIwstUVtPjq9bqHy59ZMV3A2bUZ/t/9Va8HmAtfZs47ZXKxKk2DzYXF
qYGmBfSuvODfRaxAh1sVEuczlWAAOd9ZVqz/dMj510w+G+JGAi+fhNhBfB7qIRWI
WHBlQ7DdsVLMqTA7bC91jH0FhJ1y8awtf14xE/9dghbSvo6AUHhkrCpcJDyw4g0f
BapGehnWrrKd07cz+cY2wjwHp3V8LyMD9J/rs4E+xu42VBsr75ZV9XyJD18wgkhu
XKITaJYA36Lg8EcV5H8wRf4mrq+jUXXTBHZR9RcDJK8oUktGo2fvBXpHrd2wK8Zz
3osCG3enZRYRN78cNlSyHS/yzXTbtQAxM1SH+HDuu7Jy8MUk/uLWs7+sEtkbS+KE
UgF+vAbZVVlfVnJzD2uer6/v1HDivJUqBLyiFpv3zIZQr50YC3UCDvqXgtGw9AvS
vFORCt67t/ApbQa8Nwl0ndwdRTBe8kNOqN6FRPDXhT9bl45ZF0+G+BptdcZBf672
TJIB+JePTyB8DC5erhV7JSWHFDSowR5M9sDSftiKEcr5k0nZ/W2i6KmjK6fvOHlh
9wxPNC/8z21pchbrOTEK3wesEExWm7l9vZbOHr4WLttvuiQBTXu2F3icRwZlMQWe
w+dif9rccR8ix6kQC1LZ7AMxIokhQ19Fd+L0hxt1pDsM6y1yePXa8DPZUB1crYQ2
hLJSQP62bCDErxbenorIKv6RhkbWBK3AcLLItVztTec8JpzJkJSSQ+WI2NX3VTNE
mxmN14It2ABvRbox06PBmyMdCDNN95RMEurn5Swk1qNggL7kXmV+N7dD/p7QlA/2
a29TR5XiFuGzjdBOscokZx6wQSJM22rKnVBc+gGW6C/FpisNjUzzzv8UssLZUTT9
iMP/CpUbzk+d7079RZ1eqVjau2ep0yRfwoepO6A7v07I8tCs0wbTr1ITHlBI8ws7
+huMuGKQxjDFHb3/w9fwi8OQIfmUXfTBBLLkpy1r1dHHR+MXhb288kKSFfTRCvLr
12sbAmUOGXh7BFBlP9pJwxX7RAtBH9jl3aeagOLv7Dr4LTDBYrlcmZO/nbgWu7C+
7XxYuF5clrtBXaPEJ3pIofLgxWR9/7wHDzFfjY8Rmfz0iwHCnvyxU8mBcvRSjWcx
rympvLT1pFUU4QTB0HMbgqyiMBfqC1s52EYbBUmzZ74TV5atVWNGMmDMQmj4J/b4
w3q0awFN4C5ezPK3noZGhhLM/19AOGD5zGsiH1JM27yXRTRbGd6TVUhTW+P9fCzs
gxSq+Si5nuaviHI/kID+O3K2K0cPdtdXE9vK63wgrYSEPNuG+SyUejEDuVhxfW6W
GnffaOU12JDsSX7UHxXOranooQmcxu27qJxrxGvoFgoQcXnihGMEptN6MiBBg91+
uEt+ev/fv6PFgv4EaHL6inE9Q3YrGJtGYgP4g1no3Iz/QVBXcp+yQO47AXqd4z6f
RqO03qgZC+RUIaUf3YpU9g35yAuzCeN9OG+aZzMbDN9zuyUfQSKmabtG8El8EAta
7dmHMs+7oecaTuoh1mHrCk2C5jwVEEHwR5PUhlBU6+tPjfZ8Q4L+4li3ZcTKRpD8
dRwYvJsB1GIKmQes9XPVYMuHIGvhxLWA7dDHvKDBklqYbAAPO3KMCs02oKiT0Wy0
zzuYVZEMsk8k4+bkdSWUAoAa1QDTheIzES4hRUShVq8eBKp4amThBHeUpeNKq6l7
pmuGB7tWkSYB6PZnIbyGr5/bfjtUTGmbN1BGHkklLR7yyMSWbpyCSfgYjPSf91bZ
BfTw9GLkOQE+IBlUktltXAU9y8EEA78GDm3VxqiFDOFc3XJRaDKSq++q1+eb1+El
/39+F+3V03Nv/sDi/Gvq5mij6t/HGkUFezuMFolGmoJk3unhBka7Bcc9isoo2Elh
64+zdxSWgmomY+iyJ8ZTuSsW52wlFCjzkEPfeVCjg9Pz0n9giW+t0XCduHuYS9Kk
DqPE0eqID9UERq+opaX5Dzde4yjWUBVcJj1EPZCQJgxt7ZnHQ0sDGGY3mH1Kdrmv
59BlECyUH1WsE7IVwE0Nd7VlSWPTXQ83Q69qzrMEZRVrBz4rc4nIPguyjBA/T6dH
Fn2LsSEj2DZAugSQ9VJzXEl+LxGElE7Ev/N7MMs5kSQy4f5JGi6FjmwfvtFIRx1J
8xYiTzdD5OJolBf3rGEEyi0JsIPKfOuVqz2bo8Fl0kmeS4Kt8Q3qNPmD9BgKGoGo
l/34riJYZJC9NpqCmqWgI8MvJp3r+KkNLZWU6AgkYzJyTjQES/D2qhNQTTLjzMVS
A0zmt+8ZYq5eZ4ElDY3nrNXi2YaJTdiVD5jIUeq5D3hLEKB/Xi0JLssqwwbG4I4O
19pAApbf2u3aP3RFnS9Di25npcclQ21/D4LJK0A5Ehzm5I8CJGZEz4ieiL1Y9WED
cAbtUY24hteh2htief5OOEREqD6v/3yS3l93rj9h2ACEqpIrgZ9HsdnWTDrRKH/y
H0gZA586/1ftmBer5hpSKiTNr/6NMFbGFwtgQ1YpElRWxxgGGhsTuAYMHS9l7hcd
rdBGudsrLQjGRRlHm6lddMjafxixzKuVxOb6ZVDxk+Xs4r5j1hHUgbp6a9nZrSLk
S0r5X+8ZBYNOMBKkQ8ORrpjlFSzPF1MuIhjJlOB497lGVMwNpkaxsRw2RVh7O2ZX
BaC+WbXPDDbgimxApBXsgdDd35MtfO/ul7xzynUcpRsa4aRex31hu6Sxc0X+9RrZ
1F4sVO9R2oNfnyK0Jokn0ljDxW/1jgO24YERRX7+T9dsFmJ2kYzl4K0+XKlUV4Xg
9Wa2gb6BCkgFvNUGbfsaZHhjAC+03k6bcurOsCKoco2MX1gX3YLUaogBD/ojApUk
JTSYjVBetWuWG/YSJR3Ux5fYZNPMaSEV9HFSVce2yp8uDwRzgxZ9lSxnixNhNH5h
9I4cOSwn+Zr63h/odg5ajh1LNYyvjbMf+s6hCnxLd3vihTbuXltmqNaVpHSWbwcp
VF/9WqNrWvhCPRnrVygYPYwXMWZmZopCDv5h7zybA0PS9vYPRu1GlUQUaBG10C2r
eei7WOpLyapO0fEuPkeo3t6wY5yh4RZG0hv3USYv3puam6iqVpGeOvAiggWC6vvK
mZ8HEFvHCiVMBHSxvp5m2i/nCR8/GQj8/uugb5wXxydKUPM2SG0V8t0cfVNQZmmN
KlftjUrH5bWBYFF/+D7Jomjxs2y6pPY6huG5XOgizFz3WVCkUR01EEEoZWOvDF82
ih/pU8b7c/Bo97gBlcl1mQJdE9acN+XZyaxB+7Nxu0KjFprRx7+RKayXarW634QY
lq0Yjb/mEx8T9g+WqQfwvCrrpMmmWBCsotLHGOweT9nHAijZFn83KkAPXkVzd8Wx
wH8FpjqWczXWGG3XKnGo4mqQQVxrDNTqxXG1w828b5VLijGDmX+/X10Rg+V53IGG
4q2gmHo3KOVLWefaa9rArnAEsibe09JFq04ByIc9uZmJ/r4WtYOg2GIxuV9LvKqK
QGjEPrEQILkvF9GSSz7e5rEt8qpGddbr+yDToACn93DWJwqc4nbvD/xc9gWUhYQ1
s38Ua/JS+e6iK9s0nIG0a2cI4m6Ixfy3xZVqu3yZ5MP2j9+70uqJk+VWmfKdcSah
9OzQ6HeKdOzs7MsHb8ITxBkUxZ7VzdWSaexRd1YtdZnsMlFlJSVUCPJjgWoSAojQ
YjsyohLq2jRUorOofe9b2QdnJJ7cr56t4W6VAdsEZmVv1Lp2fT/zqgG1VSeH/Nwu
uL9VRjIji3BJ/dnG+8NYFH13mxFTS+PGvqwx6DS6LwnJRmvK1TrdiaoYXp3vPKFy
OmC9SlwufzsWvq+CofntkeZWKOa0CboZV6mkOCysCVhUeWBqZdYvWzIEE0wNWYu0
wek8V1t5CtLp56uOLTKKeSCHKi8A/nqaAQOqvR9QxQyXV1FqzSPDkVeQCwsnprj5
enOHXQbZSiWw79Y3IohClrCH6cfqIV1YfGRrMMSspWLA04X0xGZos/KdWEfl5FHp
1QNJ95BLGA9GuYD9ieNKZmTBqgNXkzENRyYp1lK9VsjzJZ5Z2axTbRvwjz4hq8en
Quiv252eROPhW1Oj+ssu3SZWlzrCExXCP26eUbyE9uCiXzpmxr5FWHJoIkEbELOX
Y5zTAkWzxH5QiOnA9xxMCr1ynQZtEsOojFeCERrSMvokekK+fG9lSCZU3n5pnk6r
UJAOzRSiFxXznQl7U3GhbsuP4euVDv2H0RNLUYipiLbA7NH9CSYSFC5dOM5iYVM7
flyXjX0DX26XCAECjWMIspXQBtYbK6DABC+OnDmbN0oSewguxbFVbfSGIEIEVIui
BULDQzQclQAqQf5TGSZgsxw5quajHxjpUE3IGVBIQR7nt1V0LVVFOFgSGcWBNZ1v
g03Xzoz6NyEc8xqG/DAXNaaV5QTm5mutQ6TJZXBhyDiJnjhvbgRRMeZxGjD39+La
3r/qygaHtCh0Vi/EVxNsZXFLeUoYKRiEsfe4blLv1AyAeGQkrokJ/0Gvwoo9AmVV
jzopa545a/sw2aTVrjXDLtoJgPnRNNeFFDaBd6umRIU65nl0f8A9PFEItj1xS92u
0VaQEBGVCu86ZEcXHKIzaHSlX12TbAHKkfiBMsPspja93n4lkXrkoMQnf+w/touJ
jyq6mcsB/UuxrjzMF/q8e0k6IcXEcbnLR0FlA7P7NXr+pqG2NjS2xFD5/cQGYu6z
29Pi3CrBDZJsuJqYcnMOqUGS+BnrJIp7gL6Y2aZBuigwpwAy7IwurWFAoD0J3d39
wDdwHl2xhgfhPIj+H1iRSRHQwuO1HkIKTBgcxccgJcUPLgXxUjcZmBNhXp86JcLT
21lRz6OE653sTO3kVMt50em0tDMqdR8OiJc0x+RFuqt6zPjTIajCn048j5CLZtLD
BlRcer/ocDOyeO1kVgcBagkNydUuJnvkcFux9H6vW5ON4gxbtBgK1Y63TQVJsn6s
KKS7F3M/KoehakTHawi2gOkQlaj9T7byDCuk7Xc8VLYQ0PywMT8x4b0IYNG80bfi
I/qQ2sbRUSJ2cpusGcCyc1ThFyyVb9d0wUGtruT/DIX9/lrQ9zYBOdSfhdQ2QW9g
iascIfzogDdbPhUm9Ku3rRITCqox8TUojkYK5A+dXcZ3WDbXBtN0t+bOEuu6FLbB
WHo3Q3cBXcp+DMp95dKUK/CbHNWmIOMHF9I8togaU62AZ4akBHwOeBFqpzwtAPTu
tWFqBnzk13gcz2vb3pEznlZgGHY/Y3wN9cut/rd6JbJJihTbaWw2TcuDvhh8c3vu
bRppe4nPRpBUmZMgi751bYXxwN0jeGaPXQmILKkLJIYjs2mtug3wn8znZxskP9lj
GbPNU1IdC9CcokccgRp3KIqlCCSc2fhTXjuL5ArqR7Q4zXZt5ROLVKueeUWMLsct
Nf4aelJaKz2etqj2PIITbxhwmUflcuHvIXKZPY2wynTueOCPNz7e8RtCgq9la8Ud
i6mtdQgD72ICwU9tKGKbu0fRbs43ps7XG6HqbTxQoL3nibxOZVCO3IJd+c6P7/0n
69wDHJSMsgcUymm4t/gdak+iGs0opn7vCKwraTe0xgoIZsb0jnSc31kKGfe4knRF
IoGYG0xd+jsIQio9MQ6Q3axC8IU2kiyy8wtBpVZhJykf5k2N2pGx8IRGio2WhYvB
9JznjPamgkBPviOco/sGMef4h+MGibj3yL3v0iGw5v+wh6W5ukvpD1beY+w2XQJG
D1IkLVVKI5PaVcFLu57Fkf0hNeSRCuZmnn2eqw7sZ1JQHCW9IJ9xhfmOzzc3HESv
3y4KkM9HIpcpckxboZ6YDb1oW39STPvwx1Uk6xFCoIpTuEusYmeP9PqRNnWeeg9l
B2CXbCkmNPqwoWRSLehN4T6rd10II+RO6zg4psyjkTy6p4e7j3GIkniw/dE81kjG
sMtFQsbvOfEz9kzON/2Exhc6jLtNczxN3328MCOzQt61wFVBOmrT8Se9B+PnO1Sn
G+SRb+lvgDoMNSPPrzp7PiPV22HKUnwGKKMeQ/gBr0qFWnnpPurDzqqcnZ+QlYzX
1vLZqLKc1RRS1X4TrBEaGoC12xcKvZLGEKaZe+puLG3yo8v8FLtHQqGIuM28sl6l
AMoA+v1N9rXLX5m/m+pZYQhrUEBG78dgqc/N0kpIaS8GyUcWPcSsf80Yhro+oB1q
0Rw9dcy3oyEHSMcaY3gcL5rWc0WA/TRg3RY1IJunMCnz+cIgsapQwYia94WQqtOp
rlW3uUnDIe2D8GuPComjTV+tXPmbQqAuj72EeCbe95Oq6sPGZpSBnKz4ksIw/jyM
SPEs83q77JLFFaPttDAjsVa9BJQTIch+g7kg1TpaAVuS9bjfySqyDyzAnCFVPl8W
VoRuDOB5LioGPeQ/xlBu26R0NA+Zi/rmP48cBe+Auh3z7x3sxy9TpaHQ6D59MYQW
+jSEZs70oYJAu1lAzwtu6sldEm9ngpHPQeHJSBh4bOPsmUEszjApKWVjNNUPXCAu
j/U7aT7IpA4eqxPwONJXtFPUKpwa/xX3bD6B7vlznVUkOvc8KyVZeMywiWjPTG7f
zN13n7GHRT9zry2QpmITMJM5ll5AWT4ZK1hGSTfngLn97LAOCFGxzRoPCnaZJ6qn
4mWN6PGFCvJRjMdGqqNWg8SIaXs8xJ8tqMubH/3Xob7w4eyD/0axe+iiCczrT/L4
Mx9ZEZKT64Jx4E7VMHnO/+qP1tkKro5bQblpcOzt2zwXrdlN//1HJj4O500uIP+k
BZMjYPDtT6LFAL0UHMTWkJdDd70E+1xDbB5yb1a3tvlTQR5OhzcgFGj9EpRzxMWi
8torluKH9Ay6x7EIKoq3EN+y8CNF4J6MW2AVTJyVHQxsb6N8j0A7zctoQNfn1ObU
Io70D3eiMhONe7OzQ02qLpt2sS5p2U5zB5wOQTpaDxFW+4A3dMvypxyXzVNqiGxy
BfmYQESxOTX9c9wfqd6n4LGLogRbtxLJGcLYW0qk0MqriGTKPOH31A51O3gR1xNE
y1SBtoYlZMXDAgi9cOL5hPYwhzqrdfbYf4BnqQUqR6HqL1JDrNA8LTgUFfHLuTNi
UH2T1cvpQwkWj1H3Bj5jGseXFNv7cNJ6GGgW2HOc692f2LaecDh0v1d4vQQQ9L3G
cHqMS1Uau5AvmC2KSuhkfD5U42mkfGmhqkif0gVe8fQ6MKkihdwi65oUAOXlLqzu
klcP/d5vQ0cjUG+ZzMqLdF/qkBUpCMbO+iKTwPefcKPvuS7B7eju83PZxEVBVNpw
f+Bs1IR/I5R+bKNTs68AMh8KUTapmEzcZQP5e634n7Zn28IcMjXYgQjziu6AmVxJ
6QgsZTmErE2gItEKwneST3qK83qg0xJBm6GB9XbOKdSh1U/JlSi6Vep85sh9XK6s
HUHX/16C4PH1KTzNWRR0y+jLVFX9VtkD18VGE+O2zLlMdNvrroTqcssvj6N/dZOy
ON9S8PLfgJPXJy6JKDijLW83O1Za5zYfjdINy61Z5+34HCS0LSNDe5VKH91yVuj2
cRc65qWRoPyjDJZeYkktSUYfy3YxmCsjPpGo0PeFZzurefH3HdquRM2XeQMvBvDO
OKYeG7C6acwkfMOXkOR1YGRQSJHjNRoJIfulC0+1GD2rK1UNld2m6AxDww8YOAzR
Qi3TqPB2ZAD+n7bNvApcguet+9bRWDFl8jQAnXHa04LLG1V+kr+d7VUY3gjUN7rU
DwXfZJMj8PSY6tUyryhMhUU0nD6SF+a2iYParhFn8VwPFzLBUYK27558xP46zlO9
i8ojMwgPCw/Wk2t+uLyDOfzVbCg3o+tnCoQrVi3Py1JG5OPHbsTCUJTPpcYCwdgm
n/u9+SEOxn0ww02x01JBTyjbzfZXvZB1oOiB5MYo8Vrv7W1M6itPZ+yoaQ0wWkkW
8hYWd2SVPxGKjMPW0p33Vc6AOB4+zbFTu9RJFdF8OiBt4QLw/B4uGBggGrnwQT0/
0/j/nmKoiy1byxjlNFH+D6dINFYxkxWagdqg3WMsJ+AIdrRXnvv2tBr9VSFYXTr2
pyRa/18Kx7huJmWv6CxrR7RPS1EIji0IdWN+2W1Y+ti2Hbl34xUzHuMxVhpb9gfl
lJHiupi76h9HCL8EF9N/BP7IyR5ek0BaxQcbCU/tvCn3cLWzlPegw1SD0qLJlkdo
I3DG2zniH9hijgh4boKISNRSW5ro8oq+jeV2F8mZRu8h1tam64vd0lomG7Zvu0ZN
iQ+UoVw+ywnTCotKIxYHbJyFRj8oNVCZvT5INXjtDSPAxCnauEULj0pN3is7N14m
N2MTrhe/L9rcovzBxf2ytO6C4sNc/MRuBS6ITxbu+Q8C4yK8qcplkdSG0hyKvrCA
KflJ5GRvJk1TcKSO34YeCTv+qVCBTCAe/XHvS6ifL4qOywN/j+M3tOJOVCax45j4
x3qGCySDzI7BrWV8q93uSehaqdHljCs+EQT5fvyELYnKjQWU2NQBuzN5DFBScdSQ
OG13R/yFx35R8mghZjWQ4Bnj5wdp3BH5MHChUmHAsz2qNS10mB3YDQSdv2rJcqmE
v4Z3T/fzK2N1XFYx7wlHMSsE+WFAZ9tOQRkVLeuGsIhdQorgFK8xOm1eqdQm4tdA
3f10WcyY0kz3W06f69bi6e/P5vBywXu1qW1uRTaEuDM/G6C3aV/onl/g1gHVTvP5
I7zv6noOEhXjsRDH7mf49NjlTnyuD4IKMrKNQokLGikpr7dN1EEepc1XMcBDJuXA
/YWRP+VXOR4a89LmWKRWdmfErgQqzdgOsfHXxVUotguXFTb8azVupI9eDM4eKOL7
E58RE7e5BdPiS9dCT3aGDpxJIMdDHxyzA0m6VJB2GchqupFPR3S3PQGBPQZdG35R
jXuktk7VpzkV5TP9TBZZxobJfU7WTciKdrZOxUGHcLednwTupIJfO5PUTmg//S+S
/DUgkyQof0F+yHbQWH4hWyeSigQ/wEOtSl7sv0LJ0lpSyrM/LlIPdYlyFBmqRxe1
9hcUQlbp5K5fPpoW/N9ZSiqp4FBi0zWffDEnUkysHWXEYSkWtQxsnDQ4xSUl2/j4
FeFa3Iu5nOAiH1/gxsm6DoN9xQxT/TlnuxGbvhRhQGn/F/E0xjfpNxoh4gr2RRT6
4sS5oDSUP3RY6Rw9DldFey1G5f/ayApiXJwKM8+J6ME6WhpgGMMD8nxaggvnXvqY
s3nFHWAdD4/PiOw8coX3CFDEdyjCPeXyTAM+AjAWTI4VX89nI01KV/0UDg4w34/s
XqM65aQIsjK73R4djg/DAx4vqt9C+mRhRvGBA2SI5dTNIuNgS7FKjFj+Oa0zFYqb
4vAsHtsVmHzo3bjIp4HaAi+8WtM2iLlvXYl7EV00NcKUL5ylvks7ic2hbwPtt2bM
enFMLLOR8OXooYrtDZ4Zmii5IiCoaN6U6d9y9xMFz1y8/VSWNUA6z0Akgqt48JR/
h6D+LGUcQMwrf8GMxq2c4KWGf/d5synALgMwHP4ZZxfpYN7XP2tFkuUu2wiBeJPw
g6z8h6Egz05q9pgHH3SN9wlnKv41IUEoUyDpSs79Fq/+Knd+MugRfxWeP22nV7Y5
rYYl5hWSwrGeiDPboHgPnokh9r1ZWd6FmLs3qF30Vr4x9J4WK9J9UwNBfTvjPWsd
nmCoToZauOG4FtUcRyxdBy57nDZZB33J3rymq6yoUhOGkc3RiwqimD3WiAHrdZxz
qE0hKUIepvwZMH4QQcun9dAjzLcUjL720P2YM6RYXmuia8RfUbnPheleUlF+Aji2
zt6ryvBJn7QOVVBTcn0t45GCwbAHmuStyNnrJFVMXsNHC7F0v3AQcvp5fhDMcAW7
4VrFZevyMx66wUPJ84VXJcNV/ySL8iGoKYdlz/GLi95Pf9DwgsDPeBqD9AbdDYvC
cU738CDnk9pgTgj8zoY3BEF9UXqXgl/PiTm1pGKgLZZKzI8pI54y+fwZdD/m5r4Z
Fzqy/D+mJ76XYxRjOyjIXYhHUJGhpZVhzQmRZa9AXxhMW/l1h018MlKbXIaXFISr
JkH+i/IunNxYnmSdQGRG/8kLZf3JZnPYi57/2MFSzc79fV4IgjcWqo2+TDmfshZr
MWAr80lnEH7UAoaFeYThKuGyl5yG3sCc0QqALa5TO+a0sT/+yA7zPmjSuZYUg0VL
KEdNfrEM+GAcd2ACK7EkFcQCdP35Pnzu5PLd7NGF0u6PuVnk5k8HMmmMW1pmsboj
0yj01MDVWbrYcA6kjmQgxXJijpc/73C8fDJz1V/jKklEowCrn8RcDPjloYhCVk5O
Jeyd5C7jx6ZUOoSHi1MEoXbRvjQfoujM7aXZtAu9ee8glhpOhu02MPur6+ZpDOwo
rhfYePpeaPpci9eglxAr6aBNw1YKFQNf96BQiLzRxgfr/lZI/P5mQhdrWZ7e+tNA
tTtZR2L3hn3w5qZEqB7G4ziVjCd2VGD1DVLKfRrSG1FdWdVJ+Z3a5oGc0UdYfJdg
5ctEb8rhdkHfqFLn46eSPNb8FSVLJ5TFsTa4GttIVZLS0oIGSAWfoCGeMYaBDwmU
PpT4vaVnZO80pZyplR9+ARq9pQR689YeqlUoq9HMTFjwEqCeg+s0PYtu9X68rSJJ
o0TTe9n45x5uFlmbnVLWhpqEuQo6KeFlqP7+FjvNv9/F2xvj1cPgGArh2FG/zpQa
vmoVY8zSoe1OuoBS+VljOcmmeGAkOmezKsQG/XaKHyg2XDuVVWDumbKKYwQtLJp9
mq1wmqF538j8jodWhDeiJ9B7wCioE++5S/MJ/Rz5D9sxFajab+rJmN7/9uWWB52m
C7Hh+OKQPyE7aD35M1a/rq0ZIvUle8xlDiSMGHIaRIYldEDCsDbLS4fTDq2n0TFi
12NIB9TZ16iKlEBDYSGJfWIL+9SniEn2fxrSyJVLUJrGOeB0X0uDzKbkip8Uhowv
hPKPfMyv2u3BHuum9lyPip3tP6CF7eCslvSFHhR499a9BuPqCsUSQ6bK02nlHPCb
hdqyESVVpLGVCKNCsv+dgO6+JPEG+/TGu/lUp0DXkNXadwU9cqA5myngjvN+5Q1J
bHoR/Uvlyu45SRzAKxONxzlp9EdzPvDelyoVca13o7TjpiQV4H+fNV+scmUpn3cg
LCLR2o2Og/iM7oJ7fMfP8iWyVLOsU3A0a0I7FhfZ8ehrWsUTGtJexzpFkC/XGONo
1Ry8y+dInuWO9Z0iskEreNIj0UjE9x0sIPITNYbiYa1ZezMAM1qkh5dYFgcnQawI
E3YLBRm3EvralkS553tuf50W3wG2bkUgWXHO46Q41K9Qn9ZRa832jbpzE6yvktY8
Fc5MLjXv6px/G//QrlCpsXdTguItI0R+KMyspUedBE+Z07UIZ84+sUJ9csSNByi2
0DSMfsJ4TBVK5F/af89XeVJ1z9yobINVxA841FaBkdZ7YDCOu3Zcy/U/P2U2GeQb
I7bCYvdzlVCVyxtvIwmPdRVsGZMhMYmjwiTtX6RUR96QtqrVrLXHYG3WeGugXsP1
ofigp9HenuHiU6/NvBuP6Fc6dn+65/te+F/wixi2m6yTYP6ZottwStR+fkTH3EHS
RAsIv50agGKKBN1a06sKD1NdWiQm8PKkHieEf+qHOWQbRZzHLhFKbVmWH3cLz0jO
885bfIkClnImn2n7lo/2FCgucV7CcbavWSmpdeKXHCeuPR0BKtw8M9ma40bxO+Jw
uDhqjNtEXX18N2zGRwlTv4zgiSVGMnMUaYBrosCbrQ1wRq5S3sqxRTPX+iY0ht4u
erH32KOfMNkTLthj5KzBF2D+qy4H+1fAAM1KveRl8qWiUTOVsohwJyplJpyX6R8o
zCdukAkaRXuY/ZWK83uV43Y0muLSlTLUr/VwpwzNPkBinUajYYM1SMxrCn++Osp1
hcvKvwWjXnXdAVp1f+fXOcMUVk58p09td6/mF3/DB5OVik4uLQuK2ut8vBdkG0O6
slIZm3bTuxFfJNmfhMHhNjXNbhFBcsDfVzMbqaDntvURdX6WYfyDKvPKqFbtHj1O
cl5nUbC136quhYC566I+P5WP84Si8RO8/bylCzCtlXLUN7RZ8SOKt7a0cqyY2wnO
bUhI4S2AjPxOj0WyqdqBeg0h0iy2jRJ+IAvr4HTAqHJlCgrDG5hIZLOq9o7aqXIB
eF7zoJW9G0bdmh3Cdiq2tBoLDCcqv6ugWyxjhAVPyqHpXf9/XinhuyjNVNzl890G
GVHqnoHFl+bfnLqNAHr+sQM1kJ5/NgkXArRn4WJlIgyU42+vw94xvGUgPs20qK7r
+ICfpfbOc709V8oZIUC9hxWRClpW17amGMB+c3Z5Vcv90RVSK/Os+tPz7N5tbtXV
cDGtJT2TBykbDYpkaUZqhPyuMMuZdEbNs3a6bo2u5nUQN5Pk+GKzBdvcklrubIhP
HMMiD9ce277LKu3mhEDmVzzGS5HBin9qXJbnjSmbormjV56WgJvWyH09sSY0UPVK
BTYWFGLC3mzxT9Lt+aV1mDqtE16qsVuixuJWs4I4dtqRoPRlDmInpvd6EomqLZaY
XlOdapoKkLjX/oXJM4xu9mQuu2L5JCNqw0pplGcJjTqIEB04vS0JHaDcGk3ye1+T
qUiIhWxP/E1fc/YPE82ZPAd8FW45ZMT32R38ajtbuHg587/XMtk5FZbiuy8vy7SP
D6BKX3eC1+v1I2eirb3O50sJ3lSKIGYCsQDpJZYsfNSzmgnwShILQ78NYZIbdmRx
VEyMzhxfCr2SmNd2Ao8bnsGusF0sJReot8tcFOqwg29GMCZNJpS+CKtF8rIuGmCc
4DS3AQclU9ib6cOrDEbly76tTuJ4f33pMguaeNgwgHxbem8RVD0jEjwloJYROaFM
iZd5MoullsecDYR8TYrfdAW7Jmv2kUMxUdeT8xt9yC0FpH0g667UjXr0jwINS34J
XndZ5+Aeg/OXZvdTJTs9/afMFnDn/TvSbc5FrgIuCOJx8xKGo8lqFbiV6gocj/Ou
oBChWZHFoO+27qCtsX5TAPo6dzUsW1KptwZGoNeviXk/xIFK7gfE67c0GmVGpoSL
LDYpFY6Hhne05X+U+Y2qmIwEuNpfx59oUydSxFhm1AGg7W819Rt3wsC9OnTqVPrN
x7jbrWj9Id7YPryToscxoJFtee/P8DWcKhFxrI+I9u3OIbZ/Q6fR1fd8/LvDu0I4
XQYMUhmJEiemBORsjpJb72Fl4HkR6l9rJBCe7CgI4TJjAVaY1b+2bLCVucF6n5fT
DCFvRo/WYWjmOCHzWUsqN3M4oCCOtEZWsKUCTKW5Kp4P2v2g1Zd9wy0V7+pzotwL
K5FmA6fNpQKwLeWSz9+XpcEd1pl6EXRifyxxdueoE6yDxqxZwtEFVxc+kPuwkO9v
1rXR1rZgUBX8dQG89X1JglC1il8cYT5i5nXgex6X8NZXYLMON2senhfiuHSoa/xv
J2SqTFQmBRpYa9p1wY34Sf5tZ7OP9EYjl9PvXrca9LE6kIkJ7ioiUX9gpSkinon8
pQV53BPk2Y78sCiMyOD6ZzTQo88vGbRP+CR8VfgtDuaEk/qUgBoumUdOBx46T+Ch
D6l70OiJR1WX/PVSaN+e3rGXb2bLKNlcvAWlankHEVcw7GzCU+jmsQIDA/T3g/Nt
pPboyk43b/Z8MQniAe2CKK2KXxAIyv7LeqgUR1Wxxt9Hhwq84GwzMfQKEUYYPXMq
ZygzakEI5riaCY3ipAEJxLL0929CIucq6S+bKaXWtCbaD38Y6apXFNdOMQJPw9As
PjVaV23kSk64MueR/PYKYcsggdj2VGzgNAintVUQd8bnZX+8hQJWLuTUFraP+STH
KZ0I9bCxQIH52EVhnmS5e+D4w9/1YeK1TyjR8NsTa1WXrC1qU6uBnRpVjcfxSPwm
iNrRB/kuOEx57Nz7V0IjgXAe3Tk6+i7+OKLF+dWYcc46w+UG7MN6StcAjhpJWfAY
ysSw+deBi36O/SpigUYEmNrJr+CqJBhOSn6e8Ig6SWan3bo6Bq14oOJsk0lB6D1E
3FAvF7FKLGPq21XbzYs080ps0YJMVcZh2jmjOVQEwr3ngFxoKmdx8Ht+jmsOB5Sd
6mzXfpyF6R+yHA7crmgGX3e9v8REohIn0a6klwDiyxcPxdB6Okr5ZMdjYR4asbvs
EpqyPyrIdKZKaPpHaNsgvJUTaIOYNMslEZBiNOiSg+SwUudilsfVcjb04MzQhQOF
d4cal1NglNIiKEDZan6sllm4zO3SoFtmW3gY2n+7KrRKrgdsYsDdHlXtCcTlTwLi
D80ByBbwUDrOBOgHButVczD92+PdmZSZBMENv84Yi4ekMICNoLtMGn6XxaFzjSfS
+y4OneF9USH1qEAM1eJaApPnf0sXBq9YNrsK4lVjNyE4BSh5S/ENXdrSf6c5/9e2
8DFG5z4BWzgNRvnGFVj4yqNpr2b/O46nPdTiaBJ6JoEEIqNgh6lTxm0FpEcakl4l
e2zUhP2Xnh7G9uMVTD3GKZ7zUsz9X/y6SvsaaQbwdeV0TTemqznzz2YZcBbcC+wR
z1kt3dJxi7gs3mUfSU6PWpnM7ZGe1fhmkDBp8SXUb8vO/aD8aT1Dp0bpH3hCqXg5
3Gg+etsRVZW5KDhBciWPWZp3kNvxSvHqk0Aunmn5xrtokE5tWNm+917UyOOg7QCm
ZYU4miE/aNTqiq4rZHpt5eVIuLr7nNze5H6IAckC2hmnKCo956Sr0S9YoPelKM7u
nw4zEzfKkrWhuJo4llCK1nu5BmYKzb0/ekN8+yZIc1T31TqPWrbJaW2N5KTbfhmo
N6XFGGtUqQ8mH2DcRzH8K8XcEpsUjBKNHafPlRtUxneEhL1PZbPzUTAyfKD7Rh32
WgZckmkbLQwZhrXxQ8IM/RT8hxPa6DNkKQgXpgfTGdw0IyvqjR98eozkmcexLHMD
mPuOj85i/IR6KaEBi6xXryDiVcxOYgaYo0db5yl+KuAqSv9r3bQcebgJkPbKW8pr
fBzvMTueiU759TQ1rOgjTnCsYrZFbSo1wG2JAMODpbcfsnAiDr8qdC7oTE8rWDND
muCPK9WwfJ9A7NEp5cVgBRXgPt1My+kcBpkXY698/FkXrlcJ1VRNFtEvrjAjiS4a
cfjFISEFOvPVf9AWiLYWn2Qt+OzbO6fLNB3ufgiQwwLm87n18NAwhqFGLAEe4yxu
nAC18STMGv0P1kAUc51D1dS+q09zd5lUV58xX1Z/XVLVGHVcgJSUmYSq0lnA1l3t
Si2Cizgv+SI+chEkYYtg1INzJHNq9hojVw46coJhghPE8OXAOMpnDQ4CxLTkywAB
QjXUBbkptOT6TSZPFFpS4ASoGlCut7Vz3WneNEznd3eSPIIn8H41mXMmKGv/W0r5
Xo0DY7QDn0zb9ilg72vEVvtqS3lJF+Odnhp0noibTZAwcLIgD07up1y6MGRQfcgh
T6zZvTJP6NHQsD0zjWg1zlW5P8NEN4xZlFc0g4uMeGOoN7C7qHvuJoW71s57smmW
xCMi9e9lijO16ght5TbEjo5iL73n1eAy7a9QkhDBcdH28utmuCnSB6EPpotVSbw4
FFD2p0RJQLnNPZCYc+4V5B859P5D6K1h5/I6An/CDyqsFr7Z8ZyjxJ1eNfCyY+eg
NPqV+8LiVlBHkuHIBpEgwqhJ0109SJx2RMz7OocQ3ZqPeQMM+J2O2h70E6TVn/fA
dAuRBZ6f6LVKU4jzE4g9sdWCZ3UxqTxKXN5DC0ILCBquZYbcqzKiOBrK5/x4FsTV
VMOcOyXup0dgEX8dHbPw0XQUf2kY6hP8Dt/k35mJPOGA9QCK6WtbtMn33B4/fwwS
+D9uw/j3T2EotPhfuJ2VHcKoRM1ondiwB5+9f3KMP05CZWYAVXzvBDflaHZKlPna
gh2zsvKvMvndS0RzO0vJRdu+YJGvjvV/7R3hEtmw7zvNNrwxIPSgMOMWrfpqEDuc
jnqDA7MCcqXQ7ANg4BEbWJkpyE8eZAWxuH+niWYjmOrfD+9iAQbsnJBDEbcpEct6
phX+mZIxjmeMBGmT2mxvN7MNtR4tORdhCW9Eu4deNsp6/NkK0qRTOUSyMYT0fJ8W
+esB1jgk1QIsVcWqh+q7KYK2IEXsxbpEdRbsKwYCNBoP3vG6ssuoaBWZLs0PE8gb
2tz0w0gXvle30Qgm3ie1b8x8IkZBkJSBqZ/SiIujHTLh/koZQLsH6jrMHzQ1byrB
KiKN/qlNXswBgKEsKO1ku6JllJKKCxx7yIVZ4uen2umDyubcCi749vmRl3ZXN+X7
15U7ZVkMMHKHoLILrtxeQuzVGzsDs4MSK3EpBIlPhxEekvXIzuW0Ev6nQD/yCD/c
yHyde2b+aEfkkla9ilDMiFq3pI+2u427+km11RnV70jsESed2mwDJb1NQgjOUZak
hpQpaS7h65NJhewWPPIsFhPLLRs9h7gLtXPAvxh1E1iJFgHbxuKw0pS1FftieTfx
hmOFd68M15XxLl4Um4z9nSjB4PFh2kX1KWUviEEsh2/hKeSTvh8T7xc7VW6ot5CO
G8/xbGovW//c/JCYibsmudVG9nU1ejzY7YFfJ55Nq/UGPVyav2EBw14ykVid2w6x
jveeNh7osYhDviD4aNm/r7TwhbtGWLADF6szwQID1x8t58nbthKR0IicuRSSQ8DC
4VsgqGKHxXlEAKmZv6V5hMvzdTC9j7jkMng6gK3dR7C0cjtoVzyaZ3MECgtQu2k9
msJoPs8/T1WQVxcCr7s3ldoIwwbYhpk7S4uB0OMi+9OjZP2TGYGFzvDASDcRaNJI
3RckYDOxpcyMkVV9wKjFlIVz0b+wXKOvep3IpD2WDghdrLE66GqYQCF4pfkA4EFj
6uyM584ejH6GGPc0BD1aOwe09aMlA+XdoyrY5Mr0q9sBoPMzYNvtDh7CcJDxAy7v
vprzbYJYdIHmzhx9W0X5Ot3Bk+x8dympPc5SCX92IW9fPoZVrzsu3oGpUA1aB+XO
HJf5+uBZUqkth+GibbnERF/nho35bwlzlIp2tCrS2fbRubo7gI+A8byyeirDlDE4
7z9I6mawtt5qRtBR+GAvcNXKcgTVplRuZtTlJfdVrSA54wN7fTXFwHbrB3TW+9iY
mm4w1T6rfhwRHBhKRYy0Gjxi6ZtjcxVwxlzhmgGv2MmEz7tUxzVmIlYp85l85Snb
mfJkbxdpPFyclloQLxb5sybP23MYXzf/DtchMKJohAl4mX7Vf7HzDU9oksKoDYoO
/wOxXg75GNv0mT0SXqWqb1hnUV4uinjcBYd1zEDfeCV6SF65/bCfDeyn/epPWUTP
tMduSEra5M/pAsUOqcyFkhCUBvRwRmGyEfr/Ux2WsHoX3dPftHA9ToYvvvm7PIlG
0qiktJSKuEEcOa7NmSW6x/8Xm1i2ezQICCXXm6nwLJQeWYqRMDWEMzZhlesQfMrf
rRE5HO+x63Cov0APGjbrw9VQDbRO8rcNUHC4ldQJMxiiLdOUApiKUg6qnaF8Z19W
7VEpmMmeTxxAeK53NWmWaaTBtiiHBCuCBQl9SiOktBKgdgh21CuYcz6DS6oCXN91
NP4dti3TUukcZaGZRuCFd5Uev0fGNWQGbZeB9QeV7OULZnGtbixzvWpW8NVwC8I3
xcMkSkjTCT8URBQfK+oPjyYOelzLU8kiIPIPGgZc/WYLPWH2wQcVThdJ+jvtKUlm
55bKsXROSEF0CbmJCJJy2WJH18kfpH5N3oSP7Vr61fBE1Q7wxzDw6qWEGnS1BMEY
FWcKdtJJJJiMx67Qzoz91yLUFepNEt0ABGRN8zB8+JaM8APKwGoIz/fHtfeAwiVm
jKvadoqCC5bCTBCBYH+iRSup3ZK8iy9X4Wea41xS5VymaIfudKF2EPrR8o4+un9g
L+Ne7P1hzMl3BmONuF1vh3uvxQWWEw+YIoqEGCPxcO8xc/xno/9V0/NftOIdjeBz
mXcyGCGiT1ZUUCir8Y3b88jAMPxqMgw0iD0/696KXrQw5XqMhhkfcYeuxY3pRWMO
TdBYchGaOImlfyTI+Q9MH7AYCMo1oJKeuVW0eI1+5+AelesflUpPbnKz02Ns0qTp
0nR3d502iK4/LreYQdzluqt4H7ng1SWz0VpRlyTVugadAACRUgYh/hiMmRfGrjHT
nBIHJh55FUzwX2qR8Fm4CPXZD4tvxJzZg7NWDPjCn0Rc2e4k5Irgs8aFHy88iXBm
CLqMquP9Dz0ldOkOl10oKlK2nyAXa8AHuxQ5kcfzzRFnGB07DGjKu6PgG1otPvZI
Ddb3NlpdWs+HCvBJaMxgleKJf8uwupPr2tjSG1rEK1RW1FrUJ/V5TT9IlIMy+gb1
g9TG49AULTJfwZjuWYC9c/u4zL9GQX6P3ZFo7vqfeMFPHmUZli0LXkBGzAgf8zGW
9s7CdVHc2sWVGG+rTUJB3Z3IUZG9ajCG8G9jVKojnW/DFPYxO93YHukR+w2leEV0
nYDOa6oZHvxuq6o4+v3A/wNvsatrczMzT/YGp8MtDQspsxfeH4q10uzOoPZGN719
SBxNS3YXOVB6nMwcRz6HGa70SzM1VpthSZizwA5UovKB8K8YORa3WhME37QlMMWo
1ZkrdO/kU1Su2JXrFNjbaxDd9e5SiCft9pFhpsZP8gfs3y7Yd/MGxD6CSLYpA39b
xgWIQb8fgMRoCfUYu+CVeggLtLGYUjShKyUQJ2CZ6gagzPd6B/TmXJ9LQXIXvbi8
+fQ5kF934DTyqs0e+ryctq23hVEPr/98ZIVtW1mqY6orOV2A3m8LWbqC41UARkUt
cLE1Czin51d65Qbd4oUR0hOTXb29b5gIeoEOuKL0P+0YQOQdIWOtVLhZ7SPU/U0v
wCJFO8zZoD6V4SphlNK4Nl5KHPRXbaB2wZ9hMnpJ+z9X8o2/sv6Sikh8kRA3fhom
UN5Hp4Cno+91ozAT7z0r50msq+HjnTtU+xVh61jn4MdnEaSixmdQHp2p4oiiTu1x
KE8f2fC4Ygr47G0hpjTw7fEz0zydSFvRSB5G4ATz3UP8w/ghY0YVXjps9frdKcVh
2RfRoKe/4JXHF+XQZ23ioRN6rbToxDUsdRFhBoMyrLOnslxezr4tpxO450eaTh1d
G1MXpZO85LwMkiyIlYxf81Aq4Z3a0/y/Y5wFlHKtXkF4UlyPQ9ZC78P0LBjhplbH
z1nZEskMop39Me16G8rr24YjvzuHtdY4X2gYQwmhFaDtXTysfzbYf14wS8tjVclt
a7nRcl0fmKl2CySYpdBuhM4dRVLhDtKK3cVXj90hbLJDIkEJPSZ64+viWRVK1k9x
BkcAqYQrJxhZHjZLV/K14K6b/DahT9zly7jdm7t4JO8f3ypgm2h6Lb6Qekxmvh1S
SmoJedjm3a2VRDGYMaV/+o7MvN6arm6oRaBkEzO0GU9BT2nSweNtiKPa/eHWGAt/
SCKVaBNxzX6PwQE3t8P356rl/o1oCpvdOfR+1pcLI7QDc1gj7cveEPWiIP1BGjOe
Unce9TYi8drHg8cAAJBmVU6qryNoF2P8cWgHBSt0L6zNRhuPSvfC2/Am2YgksgCj
no16B0vodyChTAva0O9yIDKpeJA1rLNDqvm6PVkMUC3zM+yR0u4nOeuNuRKTvH1G
vNrR/qRCLWaSfdOIUFqKiTumS+Mo/VLmVlffIRUtQW/hBNIjFEeC+cAk9IYVaRRP
yHwCZ6iGGtPv1lQWH0N3a5dKp5RTBvWPB7j66wCYLjsyk5f1z8WnThZU+zo8JaXa
BDR0y5n8Gn42xOK7whIfH85c1GRegqLdbmJSvZ+pMc/01zqtQsjWs6srh6HzlG3R
a1WnPRtIBRE9EPRLXd6i6JbzxG0JO5YGmFlgk6+5cTfyKt8v3RYDVsWVyZFXmRZZ
pf3uNMuzS+r5SFx1Cw7d5sIzc70hoRbVmxcVvA0EKTz/3VmpzIw+OW6fWlfdJVoD
wKh4acccGgJSYLNiGSgsZS9JSXEkaE/scCahbTyveY6wct7rEdDCKpHgeYos7dHB
GX6CY/+JMGUOW1MoC7oAtsISOa061DZQjVkXl420E6UifT6/8OIC7p5TFGMUiyEg
fWJp5lcp+iR4LjtPa2EzY3yeB0L+DspQLleVAV/fQXZLW8Kkk5QzIGCxtd++hl1j
oSwfeqeHt7w0UGWpTU8QL+zGppMg/LWwYSwxyjlqJvJlXac5ktc78UPpmXZ7jKRX
lBecwWvgFcceNXzDbXU5ptwk99Lo42EYgcbkM0/FQ9eFyrRm+Ap8j33uZ7ZTKDhD
9sHh2U0MtwEz0J/VdWntcWVYj5EVA7OnELNH2guO6fGJtZXoRBqiRariaDUFPLdl
HbbQ03M9lW4jQ0sfMcNFHOZprtlB9BO8RQp/Exx6DmpKRyP6RV87yiEkp2KymCHy
V7gL+a0Hp542NqvGaKebeu4fueH2se5JfJWgqKqNtnXxVIn6XDmbOOh8ZaJIWjBr
m422j0jJKmQ0NLOFib1r/E99ucKQpkOe6k8XiMYAj03y8+3L+Z1l7N3AOhk8QyM0
/yqGYiNViKN9ZY0V4Ps4OzRURUZq5tVvJK3ibcYzxUuRZLLTSOHrumlhAIP72StT
3XRoSDAmf7z9nVkZF2KXD9Y7+E3geTl9WqoSiSSzouiufP4uAyDsij49n1XYQuu5
9ss8O7QXeba/IGTg2vELoqIaSqb2coFHyKvRD145oHsZAeOvbIVZFayII6MxPK+2
WF4l3c9/iWPcClEFy+fregMSRe5LJ9IWfJ09ITSagVsvgtbjAOl1Zy03+mbrDuE2
eiWdcmqX0NOHMDTxEV6ZnIV5TR33qh3JUGh179YZW0WbXKO0bGv6t0gkogLEyWYW
/EnWPG8GjaW/uti8i/CIGQ1ISe3IurMadmHjG8ADAFKAiMCbpNJCMUjqm+sf4jc3
TCdvd0TiHMSwFr8QGHIjZxLV7MsUe27rt0/HYOtkhifAwoDbi9wy9glnzsUOPg70
NSbbBBn3Kbk54iCd/7FGi7uFaCNYt9JbSP4zGOQaXzy0aZVDY5yIOvIk1AId0cNX
tpHGHkrTv7b9M4IxSjR6CsvYSbX539E0RGmRG2Hyn/X6E+BYSMRnBAwyJudm4WX/
IxCDEKvKEG+vppKdRWnbe8dHb2f9KKE2T/rIVHq/ePA/8jyAYgi0GFWtyFPDbaBw
GKBc7Z8K+kl6U026+6+HAwlhYIc2hBLF1y4tZcLw1yJPLVqqO41SQT7tnwsS6QfI
9EXPwgCY7yfGPCIPrk0ZrFLgG1QHl+tT/zmw+bJ0MqiXX39OG8iNQP3lLjGQfkl+
km9Hu981m8Rte7o5ohVqATivmRIVMOgSmd3b187Nm39JvReoEjbYGe+C9juDcosj
crJPV+wNIhACtb5vNCE+t4C8Kf8UV6zQEF369oUjtIMU/ufV+5LAOpQMjYk/I9rR
5IGtj1F3poGD23VViPVRqWHZmPVgqqcEt8Zd3eD1on9Xx6KjwKFtN3vm1deGitU1
q8JDK/1xVi8S5pIsrfmoywVIWE8bh1a0LVELJ607mIOX+UciQ/99UV+f7oZVftpa
mvz0FOPFI9FDJ53vVIbIlluNV6GdIZLVkUcMRuYLncRujpRA69kv2yjQNhsrDxL9
WvDnCVEivBz274KHaxzFM017YE0p1P3yVGJ+YAsnkSL85TknLgN99s7ChZF5JVb6
uZ9ZyeKpvZcWxBYsEmna0dDG0L7rrgjv4ejnvVaet7WNvh8o8965sTbXMlHTx5ln
1orjaz/Cdn6tzQm//8K9DLLwX1iuR083PPn1Qng568MUTJONtpDeVnZRC4r1udeK
irlfqG82bMvwxXkfwnPBa6Vv3iTCW35YzEe3A6Ke2hCQFTiK3IWVENP7K6bpdN72
Qs7ucVUVHHPtBOwD4npBPRg2Tk2Hy1cz2QECfGZPZHdCIkd9fwlkebTSqaSRHr71
kanqHJd+dHLiD2AtUap+jMReQstWEavuAXSvIXePuoY5XpYOxbJiSIQDS6fFMQXY
urgNx9YerlVOhd68zELNNAwmiklAsU/K2Mu6u3Y6nJR5SPXTxDqWxNtKEU6UuaZe
EuVgw4o/i50xAjSCnJvbBM31zxxSBl/cfn81whxjbx9afAyjIXHBu9liwBZpFjCU
f3AEsCcoBp7/AqhWuYzFTqt3KVQZn5fP12qWg2CBS0hbY5HXrGnpCz+G3/HuaBir
frHeNK/x+OlGOgI9EsMPIyyrwkgJLs4QjZJvbCkDRkqRki2UKCyJbOD6wDPX03Ma
QOJjqTmtV/+8+zMQ7aVRf6dxuqjlq7+ZqpjC7CIUSh45bolPsHf71/jif0fJSZ2K
xIUH0q/pbHqm+sfifZBexSuHMZFPZ4J0ECIpNXm9Jr7bR0KN0bHCSZNU3Co2c4oS
EkO5j5X4flPKCPU4PlOSXhVt0KCLPBwL7h4CzqqP+/47A2TLZ/65FCElRF1Xc1c/
XN5KTNsR7zQK27HPDz+dHccT0g7sbJvs/pqgH649plUmWlvNNhavZW4H1fX2OjsZ
2lxETGKDYvB//QLMcRkce/x70ghxWpYcr01XwRz3kRhxJhpx5rhM97cZ/5xrIc/j
tPBYj60+KTAXsvHYyg2f22vFPNlUv5oY2Uz3uzmGJ6tj1+aBw01nlyaqQMjFUz8A
4+GrlpIkFUeE8NELXaF+Ojgh/zV/3zBvDnPAhjfBgkJ1mbsh+6XCMBQxJsD9M6kA
MKzUgrH/Q/RhyVnmf5UQPaWyKJtIoXpFaUwirPd5wrKmAdAOJfp/LxS/hw8yeK+j
nkcnmXZ9lO/veBO/dahNzFt0g24fLS8plQ/+xZ8uWSEJu1gYeDJOyNXjbWMnPc0Y
BRrxfbfdDQ/cULX2Hl485KwkDhRRK5OZFK+WCtp/1GS9+3P8bg40OP3wFZf6peu4
IslqdFYz2gyyb9XSgton/FeDl0Z9FZlCAY+eRhP2mkJA/3NdVfJFZXIFjBZ1dJ6l
BxILXJd46SShGoyE3kn0TLMXrf7YkwrwdsWijxImr59QqZSXMFz8cOIKy4lOanbR
8SQzs4KTAD0QT62ffS8QoN7Bgqk4R5hxfxwJKvbnTLR8gOUhFkxZSeb6utZgpr7g
IRy5gLJ8mgbORzhfL+JXPwjavkK9DrrN0bikKobDm5QcJ6bQKSZ8yF1TbH24sCrX
jn7LrcgXnlQc3MhFlUmk3EK1B//PzOnsZe3uDvo31X5bNYD3Mqxs80pulwObqD4u
AU95duAT6BZMmn7XfpYPA0olcpMpGSau9C0YNTQynW0CA+ddPiDObdn9LYUMewMp
5IouVS+YkzR18FNpA/JopEgwVDJx2v+71HvCwBiogudDHKeqUgAsT44U+lGMDNgr
61mDBxerBsRLqtRZzhtvyqh5LpyfyrfBw0f/U4A5f8m6AVw6o2wjxaWi7QybGv6v
GmXMB0g1NquF8dbjMbVHAEIHgzOv5NRIjQVD17KqJWbxP1xvcByD9IeXwO7K8v49
zxb2Ci20XNawz6Scwlksi1audA//cFusiyXpaSbBU1yvReeEl04T1w4qZYAycmR5
z61Rh+swxdhEIrLl5aRFJgY4Ef77xO3RdpZv7ygAtUiR6HbyL9KnCdfQCNsq7Afm
bRa6/x0/pilLiYada2l4i0YfutgfzMc9c73VN3lXIlLxATS2zxSeHfYRaslg6yHF
I9Fn/DHRDeV7n6resHqSzYjTKI9zqc12qb6WrTSCNDX05n77IvnexXu8L8LrVnHT
dYWz0eWLpxxd9P1orz7whPdbg1QbGcPf0NIgJkXYUKSfvsthmxr4qmCE49KHdM8G
LUGfOALEvRE+pPqkNcvem94EA72G1JDgxIg61k3kyt5hna4qCfiJ2YKrOcXokot7
x+2DkUr4Y0d63ghygfLT40qChJsdLc4/Ixpj6Xq4ZQl3tFKwsd+RqViX+mTH403Q
y+9dUmxI9Z0j63FneeBEOgmwQhWqQT988iFiAbdeLXKtK2JnclHdTjYCEzlcluIu
67/OnIsmS1QJdkGz1+9sFLxtnkMFXDC2JrXgibjhiCzAy1Mai9+dCeFefJIhjU/g
hKkh8CHodf0D5p7jfoGJeasXKMGlAkwqfzvAnsiOFKAiJeGxt6hPzLZNWlf2SPIT
KSDpW2McIDHNFLk2R5O9+jCWjHGpen8sizMAazM5Xxja+LO1WcrxxjHDUIR6dwfN
iNdpjhdZmbOYsjCR0DW8RA+iWnn4X4GxIIW76adORrxO6gKAj3uCpMWGh9KmwjRx
H5Imh+BOs/B49TCsdM5X1X/3HM1g/fhAnOzylWVXF05tabz8icZc32ZBJ6vwCvK6
csze1Yn5ZeffI3KH2B6xbNTq0nMXgObCrwYMSWfekIzyaqb1RqAQOYIfrFFjXUkI
tcG3pohqMOzk1QRWwgv7qJG1vYbVD1DJSg0ELFStUfojnebrqGNSTUdb+/pp6BLZ
dDxkLQ1K9fQtlY/vs96vLVHh+ZAbtG02gC3kSMEIblT2ZXTZeztOTUEFovYIEERt
ZeYoaDveXfw1Em5J/xb3ZSjqI8DsA1hdyHZ4CnuqFs6UqhqIf1cCpooFIReciIgq
uMVeyaSOK2eSwKSncevjS4d1A5cOSR3S8BqPNSuPgHzcdsOoueASpxj0yEhQVlNs
wqXDjVaAw1vM6lnI8XBHaQAVz3i8u4JAnaGNlZLSBFMCfYN5rHSEcEdLbvP79lxT
dGtHn6yJazH225OiAnBLvmrqLcTSyhlZxas/dqJWDT0eBT0F5jSbcEv/uRQzCwcC
UwXACktr05pZv61/8t3yg9oi8rE5sIoIxi8yJ910Z3yEP2rUMBKnPDgH3hUU374B
Uqwf078EuEjSDk+pXtlR4xlXq86nqN36iSOy6W1Ma0YIGtLB0AuXOWY3Q20Ay7z6
+uph98TjTPw9L0Ks+UoSEJumbTf0d6+NoemqG827lo4bzeOaleO+FACY5fQTQeIM
kKhn0tiPqtiOm8UcyzI2mJRtewG/iDB5BU+v3DqCC5jKkwbTTtVGxMzuPIc5nig3
R/B7AXNAIjvvDWsb0fyLMLTRtxsVg8Fwa4nxrUhWSN/ympu51CIYWuPrC9Tdkaam
4wK89gzHUXYN5NAEfDYtZpouE/LmpXxz+i9mDSeJ29gHGBl9ErX/0DFVazyWLclU
fbnNEpw3G3D7s06CKOzyEjuS/fIFqpJjF0eDhMyNptV2FgYL4Puwf5vIAjDgeBXd
P871aWOSzexYECUg01xI7Kgmw4WdqhQ3KvQ4u/WQpNeUyoPXvpOF+onYOpZieVs0
SmHaSfEAx3k7sq+PODqLKtlFd6h+tqsuMTQiRhuc2ctGNGzQprC3vtOTqo8OaeXg
okvlzhLo3t1mFOoOkt3GP77A475nY2Eij7lZTKhdRIpUXZeShspHJqMxZ4Vw9KoW
wxa7Myjr+S8mO3HvPmnGKdRbguKi0/6n/DRijPu7F0/Psc/QBumGSt4grL3B/ToV
KVaBfFHwFxSC8U2Eqm3MHryP51wz1JB1pII3QEdtQY3aDOrtYVzEbTCfcowqda/e
6NGGmqtYdYqSyIdtso+UroAXz1MkzrcVsl/B9IjtGiABl5TXr5XVYH65KEz5xcbj
6qTs0qu+Eivv9BcisyyHWZHn/iF7ighMoBZtTFVWtrU/3ZAux8dLVukavt57g2d9
H6Gxm5AuJm3dxGh6Ma95t41TLAShdGq4Qccbwv72uuBHBeHeF7xzol1U0VnHGsqe
eSckqrg2HV+x4cfOL43huF2vPXGHdMK4cTi9GBvmOvvE4/wl46WSbWF5Ptf72dYt
AMR8hi+zIlMmD1YroEz+HA1hueqmSnoxS/YjarNzvdUWrNPVvTUbmzMMz66poUSX
rgl9DvQispvHlmatnDlwRiFki30rsTx6pz1Exk6Jo5F1Jr2YaAok3ke+9FtHl3SM
1If5drHTlX8C37dDY0xNBigz3PBSmDJRkZhYWSTMoAAKFFLoXQnPls6x79glp6KH
qKRSxGP/S+AnN3bON0Cu8p29jCn5HX++GqIEsKINgMU2hImK8mBtMGEH69dlhD5D
nVebd5WjpPMXZe1A5jLctJhYZf3Dz78P1o7QNaJBMcKjK4nmJw39ADkS4kk9iDtO
CMUqq0heU6u/VfzNVodoKMQp+96ipKH3A2//I12sFL6rMXO+cXlnKhE1zPKPnjeD
W6Qmr3VX3nLbf+xEt8ObuI2rnzw9s68zWDAzLqNFppwLVMXgGR3CRB1siAYEAOYi
zDxM5yBWwQVvT5OR7XYp9EMP2yl4GY2CL2/I0cM39kl+BXiDWOkPc0YHFHV6m28w
DfpXYXMz2li2kzUH9BbrLsxBuH5RR7D4Mb2HAJn/KokeVmO0yWkZ9sxiXRL5Gzc1
+QTsTbhNAHlc+XwArt9GQDjbISlmJhsnqHMIgh3JjtiVRKBGe15K66yk98ZnHakW
Hlrxc6Hq8d6+BWBOifCw06wmHXDxWdmNobVTY736nwJ4rcgTSWEGJAGRPtbwwAfW
gX050EfWYG6nSxcTRbkls2lmJzO1zXni5AloO/sk/SIjW5jCCId1zfT5d9w8DifP
a4KO7ml6ylorPvS4eTKzc/3w60ye6c/sb2g0SJGwd/rnZNPrx1n1BlAMKlEniLn3
Bxfx/vTUbivxwD958yVlxmBoFAF/gH/TRuzeclxarYyOuUjae07wRU/R2au49Ssa
GKZr46TTclYPto870KwF41fYtbB9743FXtELSyrb2oeH+1VIueRzdVhyg6nn24Kl
DjJNZIp4NwjcjrIpbm7p0vqGGmAMZm0sdPioKhwXt3kitq1FmjdyvQl3KpQplJcE
lP7wLfMB+DPcAXpDWqZjMkJ938OdUwY4OXbRU6FBTISgtga5BNdwteDpdTs6y1Ki
4BLGoLEhD5Dgqvr7cAlq+wc04YiI+v35Bpo9zInuX1DsGPQWboEvfnxuE36TFWck
9KWm5Q8Pp5YHH3GgTuw43rYmb6GLtm3mXJuFTbkl+JvW/tLCv8CoR7PPst2NFQlw
+QAmoDh+jNS60XRvRyp549eQcq7V/Mkp7ZBhSpreqE1LIgkPtvWDW/75w6kHKXHI
L6adBP9vxtXcDQudcQ4tAXXizfLzNXmmQ0oju0465njtKYre1aVucsEtc4SmcD2F
S73qn5wyRS16GTM+j816gn/a77NbhJ9KIurKZ/lJV6QKoVfv/VPLN360FQVCmMOY
v7U0OSXFU1ne2ePTzcZS+a8b6Mj4nDfF9YZd7inXPGj2dudwFJedUb/M2+DkODBs
oiuFR0bj/QK+XNUG5CI1SAVnBKdunmY54Si7ed6kkxncRwKxMS8gwEIqZlKqYl6G
n4E5Hnc3OnXbl3OiunVXvyRuFZeenkqFnbkfu9XLCmgC2zmwmu8/Nv+WPA0FsWIT
uvP8hOmkNhpclOQ2Ff1adXVxP7n+T7nI9AaoOEre96MWeVvpoli3ikBmzPocPt/D
iphOdRSmMit1R910HXHGAWauJCQP47KjE2HyiW1kxymaaKikb20vzBc+VbdCUdjw
+VyAb6K3h1sYtzwNqMuh8l2TpR5TBB5GFMbGUQ/HK/lcU7CJiru6yW71Saey2wYL
iS1+at591CTuoIehRgsyKBL3suoH6X46k6ENirAalYSO/TLURQT2z8GTCsZciRPW
u8Xu9mcJbJaMcsm7k1uhKh5c4TORJuY0CfWOX0xr2zsaG5m3V0n9fycHiNssUtgU
Ffi8DfkAonUegejqxnN4GBNvLI11S/UMwTfDztTBba25/crXk0MceV6tvZTJz7Ud
cZX4Fax8ChN7pz2acd2mIJL32yW187TXZVcBDXw9wTRrGmbmaigDqgXOKLKct8In
7Cx8DC8nwcb65+vyuxd+2Rj1COfrfWe2Y11nOwDG6e3lDxDlWPVwrtxbC7YdiL4Q
rWp9ZIf+xif7tAEnjN9sCRW22BfCFQfP0OGOiGMYdyNzheLp427enVaBPeq47qha
EcARjrbd/63RCrU46P+rUJcQBT8g+TaO+tBiostvFseJWh+2diqZS1FLf6AGrtpJ
TPOGsONb+LeRntpj5YsrxHowOkwzmhDKIrwBr8XfEX8f1XQW0m1NRULeYnZUMhS7
mfp+QbXebmIRjGal6FFPBmFW32w9Gb3jzrUS9wIZO3mW3DlBdVqKbLVWLPJ1fGtm
YTDXXWKTunqqKz1/2OpWetUxmNqHx5xX99eMFv8Fn1nf51EMQPY8JQuxyqts8D8t
ztBzeV5mCwUiyoUXt5LpUzFq/ulC8skDk80PgbMw2Nr+jfGFLPg1xeLRXaQBi/Lj
sIplT0Rv3MQ0fWojCrPZUWE5R+3J1CKmqyZLxEZ6VNtyz0EBXfok/d15ihjlRKR/
xpDX4S2CW0duF0fzpZM5Wmk4D1oRt/u7Sve+Q8ryFnWP2CufMwyoQ+z8iGyPaX8q
6aCzg0/BOt+Hmsc4gkRR/Ug/xSr/loiQWGVJoF8KhcFBSNoyyv/EWx2+ZouhtIxi
s1RL743O84JhWnEh0JI38b0GBQZTJsnwjjX3+bSNQ46GgVChMGj5HF3dK6ArWpAr
QLy0s+dNcuH5SER2nIzwoR9cvaPZVjn6I4QgnklalAPPLTnV8aPM+F6uIi0u5FKh
Nx1XdyqlNm8ueNT6aYicv6sf/Mwwf6HxV0UwdFT29qWi+B3gkg2JPg+/7/GD3s4s
/YMxe/3LZGbCVjijOq4hCSL2ZEroHAClhxwxzC7dFnxcDo8HBI9mUuaAxKgynJxr
E7fQKPD4+sne/6OL0peu0/+3HvmUF00KVcYzU7VW2aQ9geZ4NiftBv5z/zlgM+AZ
BCs0xvK/AapKDnsYBFalwVopQOn9tXr5iQhnmoJSug/+p7ZGLkFGVJSN+zcY56U/
I12GPiLc6uAxUktwR6KlpMqBJCh0OcZ19Bmbt1CWtVNaqMPSmKhSCIh8rhwQWHOw
/wSNeHoV+k1mp7rIPG71ELjGE3mPf+nYsh3xOjubiXbweueuRawthNuphY05Ztql
sNPCkRwEu52xed3KbGIMyhjpdQBe1KXRC/KyiQS4WkrJzkr/GW5lQ46p2Mi5054o
3Ei5ZrKqzJFpucl7wo+V4YxByL+nz8bZhzXOicjpf19X+CAveSfQLqXVVteeAvVZ
IUy19kQ3KXcU3JmB4uRUzIi//C6cXWlmpJv0C8lRV6j42y9YL2WD/3718UP9lUCD
7ME6x6Tyynte2jKirwTtQE8NYEOPvkOATTh41FSywcZvv+wJITqlCjUKL5JI5aLb
BIwOVYfq0++1cVFhT1nE5Wid8VoVOr0OZFA5BGeC6QPsYfw+ept9EMWzi+OT5mBp
kajOx5dbIMh1AcmogUN//78Tm0dHs8dP0ABr77QkWRh+oJ9/ACb3JG0jX4GUySCd
bfeplOLMxq1a/eGXe7YUcxM6XxC4k3vI/A4fnizplpVuP02XiuO8m/w/UIJIFiAB
Ys5+o6MtwtpTYGzl6lMfV7lY/jA0FxuORRttEeil0g/dvWOcCibdpcvLEcz7TaAa
ZTfoZd+IMMDlURCxB8NQ3bCD5VFDQBjYM6rdHBP/Gkz0I9uHXpkh4AfhTX8MORBs
ZUys+NQJvGmv7RXuKQfgK36D3a+2V1MXYfezSL38vhe4D1UJxnLt++b3HSAIZl4n
RVhYBNqkq9prfeapd/4HFOLb1HJRumtHgpdD+yN1ToWgTDDN7Pzrjpnfhjmu1t5s
KfbmSKRmTnlmlo404M/Mc3+6DN4OHVFCh9BrXEE1viRDY5KmvFtrBex94IAF+68g
FnOcLts8pqj3wktKHlUDvkY41LMbutaAaSfSHlItxm5yRsfLXDscdkuoT/uahHAn
O9vdH+IQnFoSAzBtI3Q50KgKPj577Y2KqtmSVK/HgWVxMHM58yAoBF5nyejofFwl
Uj3j4s5lCrC5ollDxUBOLdG4k0rv7VuZvsOnpRBPKa1qMmrExZcZEXrlGoZaoBsm
2owUZEn75VVgkST2+vegHeaYZBVJuFgpNDEFVydccwiCVX1xvDLbCtnCsLfWTxHH
ASXbDtcbohp5yL1uf6XotKV3eKGe7cTBnrLbRu/QpbUW6GBYNp6a5uL/dmeCAMub
+KL91fF5hfhtY792s2Xf+npFcAeQ9fYnfM4nYi7R2kb90rB299XFy14ATer1AlgW
HIapQcsKvSK7lZBjyrVPnSptf6guKEWEWmSucQUqJ8izejdXXT3T9XJdoSjjYYye
huDNVu7w0R18pcPhTmCNqCvpB8V4nD6DejULEREtOGSTe/3FQAVPm4Ri82ZOgmLq
/hD5ttz62xoKuasvgGZvd5LdkXOzv3+aTEmnS68q4b4SbX2RY5/PczIozaw3u/vK
GpSo+O8WHvFqF/HzPnby13+pw1IUbUqqSm8+ZVn7uE22lIVCyTa8umwFojdq6KW3
gpzPizAPW4iNNmmntErONUAUstCWc7OY2FbPyocam09ysGFgXC5J0GS+jkg+oxB7
tq+9MGu/rbDbPwLgbZSpdPg9XPnqCKeKyqRFb5qBdY0uiIejVaKcC2UyMCq/cAne
nKF2AdT3c1g0Jum/UNxYO+jt08YlNe77LdD351cY4kPsQn7DJSyf+UEuLqS8BRH3
NejZwqWHp+ko9HCsOYbGMQ/6MYBI4X03e3V8pTndNH//PSfCEAKDEY/7srcEyL4i
WvDnpkF4hdec/fKFAjOu4Uol8T9QROsvkHvLDsLq4PJzQaYQR441Iq6sWEU/8APp
z4GcStP95HVZIXu7rKrkaLUg5iJYjA1kdVVBhjEPzVpQi/HZUQ5ywIEG4xtO96QL
8TDb9VT1hVw5DD/8uvTp/5VFnQf1fiJQrNVXPL7iL28x3PP0Dn30iQ+wkH/DkPG6
2E55FJ1tx6/gS8GMcLfUELspoNl6+arjm+sYCE5XQPvbqxeDRxrrlGTn+W9e4N4G
r8WDwguHWLqrGnZ3cygIzh60agGORQZQdFQOEjvIPg789+q2HoyrXmJ+g5wW50HR
vdhJwBSh3hYz+HtnyCS4WL3p0sozEGwTL52jbf1ABb2L7gLl2IHan/8lWjVHadaA
Al91LoiIiB6P3yKcKjR9cym2YrkJjB1L1M6NkOktrCONASDIOXW1WvAuoy2SjSqg
tD/hoAX+TMX2umeFw8Nb5mMBhUQENiA28nB7W2JzkhcivlcDsMTrk/iWy5Qyf5NK
d3OxGNWk/QBS3EPNcXbchhIqde+gQWO6MgCRtJw5YMRNaQuPg50myHkzL7K4pUvx
xcwx8ILT6pjRKq4KsG0JTC/a6MedANekW8C7SoiRS0DvjxoS72oFdM88Myj8MidT
Xht09yGOhHHmo+53LSd7W8RxtyO4uX3TAv+5UoynpSvU4hGW2X3LQEGRmi+S+Zrt
omGzoA4LC9eTI+IyqX6SvsVtTXdkLKNFnYF5Smq5XinvA5JP+eU2QxbV7Jw+34bW
1f4nPMba2i5NsggjLJeJHc++VO43OzSndxjUUQGtLHi9V5mTOpYvaQ63Qe4iWBY/
2BnRfuLwK0IXCXYQtFARZOR0/IgOnBhbhZlC7um7WMiOT7CPK4rjOL8O4cGZExwZ
19bbmfewhZ+5BTirguYk0mgdQtlxac9lnqVMl0hlh+cCT4Vtz1djC65dnItcFM8j
xOTIgnd+Nqo5ryjZJLm9t9+G4hY0XbaEbWPrsx5/unsckLbPMUnKIObOguUEW+m4
/6Tlge5+9C+TAZtiEmqycOUB3M+gD+u/uzP8WG3nf/3q1Noevw3Y2xyM95lX0QfT
qPtSTnD7cw09sZ+MTYFyS5pWEWRHZr0JMA0NVNLOazVf3lin6gxkbS4gyUGHUGxQ
Cxjz4hvG5OPabogEiziP0I4ow8vZyY0ffT45XuMnLeGfq5o41MNIB/DRsSdkNcFa
2ieyjT7C3Mrq7EBPQOUsNgp/tA3UzWUVyLDGwzSfb1ZmhmJUAORU3oScxe9hz3d4
ileDUl11hjHyiYhdgfoPiDtwuQ6UukDt2OtX3SfgnNfpF8ufM69qlrBg/xugEv0i
hT4ULLzjfPtF5H5kqlaD9lpO6FwhD+DcRf/gtE64W/NfOVnz/H/GI5Qqz7KhlrYp
eOCFQXNBApZiAxMok/9djjBUVM+CLSU4WtQZtP2cAY8Stcklkp/+QlgMm9lShGJV
lXjuyvFFI9ALZK4tNvFwspeWb0oYqJgSChXgwKRNYnOwWn4JTd3SAFgf6RaOHNOS
0udJfLa3PSg6cc3C2Gos4wEAzLX8nvL8T3CmvlLfOHoOLl9BRL06jS7tsiC90Qtk
5t4bYuWUlvnOW8m/S6J6UfeFpKe8scQhwawHnV+CmivpQQPJypFrZCJULvPY8ClT
Hf7/hy44mL5WiSBMVRMkmFM1PVd+WtzoN4oTAXuWuewVI0US8NSJBsljOjSXAU5d
leEXwZMTnxkc1/mlKwyG6IdYW78l80KENBx1fM91f2l8WObKFRecOJiCuI861PJa
UFLEdGtPbH8TUWXCkjZTVkL/IH9vC6NVRrsKgqWYWsItD5PCgfkbrI9slD6mNFaA
Q33j5PKERPzjEB5w7+juSRP4tnfvxKCgaPMMCeS158ard6E+P27aAsK2lRw5cxjl
Kzeyb9+bFONRW8yvxliywznAd+CAmMTvgEeV4+OvW1/5spJpJGWdvhDxoO8y44AK
P9CF8UgGugmIU88kenGWI5gb3OSdzpqBeH2rCboio7IYskGM0bNxoiG6xVTlCQhc
MjktAgNQdiEvsPFx7qhQ9C/2lsMd/Ebom/s6Be89Vtc5S5WBbwmxo4AYhrWw0wjw
8KgLKvktZdTsHUffOT+8OhdyMQEdJN6NafReghCR7fB0vLoJAdLnjp/C89NNTVvl
ziABawI3Mr0bn7pnk75QUj70+F8k1LeYHLEi7uujhhtQHfE5b9QV1IDWiOl+Euum
5UF/vkIF0QyVXGDr0dBwIsbA137Lj2nQMSnSoy9mj4i0NWwWSg+XwfMKQ4zKGuab
8wE/UIPbbUjldXtnrZHtwQhuxAKd7OyF4REL+auS6kQ45jhRVMeoKFv7vVXQPw6y
KTjnr0FSlM1+akDyPVG31KwX+bsGYmQO7FU7rmXshsF6Rk/5vosO/WNFrEqmYb67
CmipwS2hl8HxBqtoLs70DonX+avkHUYV/RpIwp4Gq1w3uObs135vX1Vjh+WYTKzH
sUEubhO6TboaduxF+dn4yW/OtwqEvTqopRrHPb8+R8TGM+IPXZGJNLVoUUeO9uUq
s8y2DsI8TIUqI40xMoG64PZTVyA4QqbYT/BOGtIFbeR9wQgmkS/e18ovP75srOfO
jf2a470LDruG/WaRo7eqMeWCJ4CDYsSq1e6yLJsNw4TOXKZavLR07CYVZ08aCJvG
pBqWxZb5XvvpLDICI7rb0LvnOfOesbUHwMFek2CnbN8angAYHKNgm5Dnw6vsNsF+
9hgOINTI4q6+US66rW6LVuoeXaeRryoVxLNtaPdUF0FBNRy1nQi5nD2VXQh7dT3G
b06j4Wj5/Y0Ghkc/va5MLN1agExGQ36YybajTioDVu82r6ta7FalJMc9k3JVIicZ
W9YFLx5+/7aDM18O5msxxRTKca1QKkGnbu+LT+zVJZiZhdQK7+IsjweHBW7Rc3KO
Go6y3IqzNPSmRYCWczcc8V38YWB9JUR1bRUhrHUGe75YaM7qUkG3h44lIEVihpce
Hti1/6BYi56or8Hs+NwkSEz8V+nSuA7sVKrHMLeGkb2G751+l8UJpahCYo16h08C
ceHlVkaAjrOPzR/n///rLP8k2VcRZRyJ9g3+Ed0CP1ZUiH5wj7D6pUK1PBEdWrTQ
LNJR6+EjrezqX4DqujDVOPDR/eCoH51UZ9Xqms7thqNIpQwTAWKeMi1E03ebghA8
RCG1uE1UUJyBuoR/Vo/QqiHOvNDEHRclpAAsRDGotLCb9zY7HHDX2vN5ySLOY+lX
NGyag18PABXshZImMHOHKFTCvN5rOJ2qH+Zbrtku2QxIU1K3Vy/VkUC1jARtael8
JKylUtgfp3ArF+qN366c6u/X1NDKKFRuKGF4RZp+2oUGzOD84DF9k3NM/S+CKAjU
tVQCe3Q9qTqcBnfFsm3g3W3GDKAq1JFlePhbPaVjhquqNXmntgiLcz3RAUeIMvpU
gu7Iphs9x5lJ5gqkpJnR3H68DPa1pD+H1ZUe5WTk8xmwMVcNWIyqMsAiDao/5Adz
KZgffp4Dg/WDOeEnV+aDEAoK0QpGFuE759vPHMavk/Qe/Fimh5OWr2oq6lU+r4AM
X96cmiQ0oM+1XzsSyWmiP+XrbMxA5wEE5jndfLt09rshSblKrmerf9eYc9Bzr/VH
eSov2bM1zzkPw6VcZA46Tw2fJ9eJ+b11Zwdel/zGTLQ/qqbPCHfAtAaUTudwyuUV
DPKZ8TDiqaMBvMnWLX/atTi2JynaTz3cV7aSTd3ht0yPlAMATUiSnoMunOft6nja
JHhiwdgFdW53T2wxKKZxd0Y+4ceD78GM2Q4h9TqxklijAUq61rLmfnvUOmWO4qER
xSz0FUb1sVolvQIj0hsTB7oZD6RJQxgekUSRe5qG/soOvoc3xEcYLMtUE7nWBgKK
9f3oEl4zxDY3l/4UVQPCGEGg3AlmL7m6a6YyE8hp3CvrFtCvKnFP6gmS5gwWqLsK
q4OSssJUBqL/dr/uy5A1Dorn02ISb5O2WTH8bqUrl4t9d+ooU1GIJcbsNx4QnxXj
XPltXTY9BrECsPf7PeLuAnlkMVnnm9mFc9UO2awQ2CguAxVeSPxNXAJ8mk7P8wmh
Y17POBfjyOZOl4eIx4ucFp+CQCPYHQssxkPnTdo9KSDaMYD4PPKkrMdUS1JDK9t1
DSXtnq9yFYJCB1f2HDpDeu4XY13P8H57wORauniPNd9WNtk50twwgmyEpEnm+RQI
vZW2rKar9cbYdHsyuPUZ3ays2zJu8Ubg5KHjVHUFrZO1DXROcjufFAwNbwC3+Zlv
AeHVhfSxnCI3YE50yjrVl/W5pnnJKXPlaycVbCLuntrKc3L+7sVzyuqaVjp1HCcy
Ru60SYaHlrQsvXfM5Z2gulsBHYDyQWyrsoGTqJ3oyPbXN5Dqgz1JHRFKwedRG4FN
98omQ+yVi8y6zddS7FqruVvnx6KoN6Vp0iSyiK27QQxOwHzPsXqBNSpgONX0uO24
hMkHzeZE4LQcr+vy+0BMQzY1na6ObgmWEzU1DgrJ771clFtw1zRBmyGvT6NZWn8z
TUXv+VYPKrjZVi5wPM7LUt0PckXslxwMPKzC/oWAo+xv/D0WqY5+Wll3i8AJsij2
tDkg7NAHQ0gquQ+S1ktqB7avzD7JIABanuBjZNWnCvqWIOpKZAZzjPHrPLsPoTK9
G1XGzFtAwAMMNqj2qO2bHffYLeOVMx6MgkfgfY3Nt7G3P9CyllGvlartrVeDlALx
XdyGTZ3Xc/0wSX2eXX00rzR2pLCfRcuDw5mrXPK0uK3pKhcyBj0FncJ/Flm4aUdD
N+V4m+dwMKi9zrzuzPH3pfXxfTnPUS/19Ot2twxPKkVaRy/bcPy9Ts8XPpwshdkq
WzTnLjXXt9/CIHoD0IpJJGFepIYSN1aKr03DPOnBxN+urzoM3hZ5CQljp9isvGf6
k7ez1JRmgxHoFLZ/+1YsAhm2XOPCEiinKRNtJA3h6ov+c4I0LZqyz9eU/uVQ5QTl
c2KFmS076xki5t9j68CT2NvS0AUZVnrpGMwBMIUan52yy1wekwf0vSLKxvv/qNq9
3+aBnQpU6TmIfvxreUpN0OHA2WjtmEgIQ2OSXjyhSIEMVnlET8S36zkpwElDjCyK
OKJzEGW6auslnxTPQBZzfxEI5fhLiI04Fl6+5XWA9ZX3egZUZxlpT/LC/XawhoMQ
VtF19MrY2X2DnGajblzBZpF6uuRqGYrsJVrA1jkpJQflqr1JZh/afJJy53+5mXta
euJJQkUUAMvwiQE5iQKWrli14W37DJjDFZLMdet85sU/LxnJV7V+0WUvOj20HuoA
mehwEfvhiIZgg9zGOTNQnK+G9HPJ/ggKnESeK+tnYyElq7k7MLRyUZSP4tk9W/BW
cIKoKiBM5uvnwaK5BxARkJ6Guv0h3RcWmzYMfU6Ni0ef4zNrrlpWiYeZw9c2a6KP
I1fqWmW4zyYcYICIeBVjDK/cDiAeggjRbUANR7/3NM64uBHluy7HjALjyFXzYqzQ
hs43CP2/QqoECO7OxauZRN2E63Eywns13lWU86c533a3pIy9f9dEjEMkqiEumUsZ
Xc8RIVs6J4eHSSsVaS7snht5jwXVhlafVxThlmVnMjU3zFvQ6x+4sJpi6VTwX35f
Hlhm/LU5An6SrCo1ssebHqbqB1HOXH+vTCm3GF1Cl9b/tu2afFV3KH41KwSQoaRV
T2US9aGvfv1rSP3HKmbGMnFT3PW63T9YrMHlijzEzQBV4HZ7afIac1XxLy8eKtsC
wBJw9lu1Dfq23J0SGUvaQ3xpKfvuGnx+kiHwqDLKS56kXob/FqoQEuwDkNl7bbW8
Mi09RYScoRpLdYKvjXkZoP123pv3lnhqaWrJ/UfUkYnsKQmG1NLhswnkw6t85sYj
eXYKvoN/9w/m/JYnG4B+PMgeCgokDJSpqjHW+BVw3scrGa1k33enGcYaEcuCUfw1
lx89fxjqvM3zqB/1Ne1wokdy/4wOz9EgkTsHMe3mvYQ9U0W8+qiPpR6X4IT4pnx/
qw6ur5xXOvs4y1IlOZaoUrJ0/CBZdKMsbizzup9LmwRjbrgNlklwts7aQ1Du1p+v
GBVzgVqYC82lkQdTgelfym5OXrf0bLRAHzLvP0izP0PHY42Q4uzdVWOVXGW3TfAy
IUB34b6Xwows7C7SYEz5r3dIU5G610Zt2Hg0QGrit6VP63BOvKDte4Z7IBEjrPNw
xNmjljs4wFvZCcA8QEnpsSacp2BWYHY9V6Q6ZCUGkcZ8ZGMi6DztnUlomKErwl/x
ETfrhxcUv9P5Km2ABTrAiaV/12EyKueLzFpA6B3z0+e3U5YUeWYANmqmDKijjEUP
rm1o/SMJdyvVAYHrn06u4q7Ai91tt4pgH59EXrik6QGOeanwrbfP3OIend/INhN+
w/FFXUHeqAw2bwuUoidJyz+m3OpuQlySNbLdap1oofuIiNVWXQZmuPP/KNTbY2AC
NzoSxLvr90YbMPzoXmNZwdP2XIhexyemRORU3iYo/pC9qm7EQxQDEUz4tmJlVlcP
rra7rXzQ4odaLZrKyS1pRV5FafQZm1KlWHs5FID2S4CzZHtCALi5yqPw1q6V0ta+
Gcdtc8j8KWB//aUuYJkty4GLg9O6gH2nLftWpf6U8BvE1Lg3Y2H+6ye6Yj7XMP6q
fjrEmeSV39AAgqY5czelgyPu+2/CqMX9d/E0ZSlVDefHT4TxWBDEwHXIPdX/WFDU
U/Pt6ovtrN4PTjnP6O/jmUoifcuu2I2aK5vX7hIbndpMDIO2ain81vgI3jZca7O2
B6YyqbeXfczrOZ8nKEzSoI9wfJYcIJSH7C2WhoB8WR5r2T9B3oE9AfP7XXjl/6DA
JQxu6iA4bboIYgh67yhOy0JtKzwSBTobLQf6nIAx2tVxQznflmChZeCEbLP6lAMi
7u6yvg86VOjnMzuOyonfyIHJxQI6XWfawI6L8CqgUuvJymOTQQF7BqYnRAtemoOU
ZgbnyJFSAdoIjfhLXiXzkr7j46sVp+1kLGIzwy0WSuhnAsNMO8k3sJcr8HV0PyQj
iTtRpocv9T4ZjI8I/ISzrsCd4wovEzpb5K/BmUkekJ+DNWLzlWjyOCuDUaDJ2iHC
AUOQRQwWplmhDfQGmra1pAw2H4t0oz/TYnjledlk6yG6uP+fFr2Oue7wlXGNDmlN
PeMhlroWXx9ZlVcgZAveaD0lGjCFNZSBuHtOxfizsKyc05nVMfzvwtObHeeanotI
8vu7leOiGHoEZ6knsDtpAhSyDeS+t653G2qNaf9BV3cjVHfJn5eS1T/+OzPsMomI
Nugacps9QQ7bRfO+cwaJxKpnVRW6CRcPRjyXAGFU1W9C0AlGeI200Q1VA9AU1xnh
8HMqPz2tqLh04Orz0lvjZ5uy5S0PPx6e8axL/4AQS1HV3eCsCJaZWatAn+AEe4Je
bXW81Ow0jARpEeLm8Qc/lI3A1GtG7q0mrWZECEYOs7TQMXRsvF2h8yf43cEr4yo5
4pEO9a5dzOc3ezG0sajTfdhGzS9/fBsWTkPe16xagcM5LiftfiQiVumD2isAYOwt
e1nDwa55OWTezyfOD4s4r3iFOkCHcjFSI+LQWHBOQVx7hnrbn+SbCIXhJuoYfyY5
B3sr/a1LHIxpMwNBOkeIlR9pIFOu8FaQRHg+aQhennWDFbvLHWU7gPY/TKy0d4ZZ
H2Y4bq6Tl4tuc9eCm0ei5cQ3jtKM2+0HeKGC9AfezDf6rlXRxoHF7O6LqNJ36KSh
Xq7/mXbbTMEVotP1EVImLA4PLh4frJiDdwwFr1WBavGretkUwCXaL7jTfdKbfZ37
smRGda091YCNO1VPwgubHTsoOCjMhvQMyWtDOmdF2LrqfVoqbu7dLryfcdoFz0/J
VuB7wuxb1zINBWO6vY41hLGNhoTCkjZafC4N7L/YIaYPhssJxhGDXuBHTfWufs65
U1wy5wS05n0794UmoR82qgD3S2riu9FEUCKepbbOybTTVBcHSj6VrE9/1RMdItiP
lLxNxwOUFyO3yKjYAdriAqYUttEj/NVvrB9VUqQNq3P1vu+Sy2PvbNVYgeLdGEyf
LeIUrQwTwJTcMAUl1dEPQTsHChqXeCu6L69gZNEBDefDaPLkvmTbPF9iu35L0Qj8
MqgHu/b6MBSnYmvNSpJxprIDx9K3Sao649rI+R6sG3/1EXJgZhu5fXuVbRacaEAr
eyA0OYeMV5n4K9Nn9TU9K1wNoLWIkSPGhZLhoE9F1vcKRD7UrxawudJM08yIURHS
jBN9B3YAslzxqCCiWtlOLNysRslJH1DJ9qQHSpVHS6ckgtCJ4YuMboGY9/m5s6bE
Dmu/uscvf5ETqU8YMExJ4vj9s674TaP7LWbLn0Mlyc7fSEDTPHG4M7l9ymI44q+7
q+7RZ2tr7nt26ivmjZYMiwOmo2bf32ezKDaWNo8YETBQwSpODO3IwmQgxefnn1hU
4/xlosJlhGt3CkvE4R64lOXh5ks0ayUJ8LwtoyYv8BVGGN2cPKYKxwpJ+SEDQeoz
h4GciuWiFhmksmAtMEA3sUf4l9FyobZW8CKHSIlDDL/S/A1NTzQ+sZMovoF2ZWH0
IftegNJkR0DvIBLIS8IyGU42yAoH5En8tjkdLMzZVNt5KcLccYG1X9ch1ck7y8ue
/JpLsLA9hmR9csUOB2klgfrcc+/NXyi8vQ/PjI6aInWapis6lvUgXMRzmIjgGoxl
x9Ol1QbOxcMRFJ6PxiGcLrAOL9msHIsVzIH+Og/oge2hrUoF58Ce3rkdBRFupW3B
7ATBMYxf5IE1wqRAG+sLchGbRrLqcnjiEpfp088b4VxZTsQd+R00CooJZOhvcVsh
xVwte+BhPELSVudDy6Ry1TwztchDkzgldX2p/XEyIcRc7DtoFnNbaQoyETWJswPp
URCt0E7KmZk7AAyLCkFIMJJVUECs3WFPsJ0DI0X/zru0+Dq6Sq3jU7blNr2xrLqR
q16yXjtbsFZFyRY9NlrDxW5E3SpPCA8DyS7y1oHUwgWVGZOQRgNSilVCgkCokg9H
0KcG0PTUq5J0qpVJQDNQCW2uPTf2Ts15WTSFvVIjM/5IpbP2gUkhO9AagswzUHsc
LQWRKm3NgyFkq/wb8ZcHV4d8ykR0asqlS1/i+eZXg+H9+IlSFnfZxiHicSNzWWsG
CfUx2LK1EZnicMbI5B0wkHrsvpjOMIoCYN6XdkcagtpoF57JMyRdOKADqoRzk3zR
T3TrsvwljoMwUmhKnjudc468emFZAi4m4woONzgVV5/nbqiVbTeXOCoQ8HHXoTP/
CPf2aHtKdgs8eorxo+v5o5untjgYrsZmiGZSLpfZIcRtwGVuri2GU9x8HmZanrZW
HKc1wC6BHkShIstm1wk+bvlVXdbNTCUacN0gU9kjPZ4PxzeTxIj82dC4djbnpwv8
0pAaV/0JHVV2YsXgR59tyJvCojBMH8bhwxPKh4IhOUmY3gi5ZyfHgP/QLWGbAObr
5V/Tnl5Ra61JGSwgoyCP+iwCV/khrNCnUMAZl3RYT3hHxrbd3Be5VvvXQPBdGLL4
rj6em3kX2vFR5oj1w+C1sftTUnIhSw1c+VZzsid7E046OYCBgN+oWZ4GhpPQrbJF
j7tcIyvL8dhAn1s5nQwwsn3rFVKbell2V+4t5qKk5T6EiE36m0J4xhgav8auP8b5
7ilGSww2XpW9d3Lg/viWnqra6NQDNV6ANpy7ktCfp3rIr07Ni19ZMWe0wZGxYKeR
vRB+LEFPKTaKyS1zNj2z+lP+Jm2hxGczNHnBeysWrusz6DSSL74qlG0y8O1vzD2S
R7Wl5ey2xueFG4AAt1P6BEF2zSkF6uMa+19fNjVB/F//JDs1x2WQb6217oox9OWb
K3Q5oTAX38KmbQyyXoXX5VbpR8Ry6J+BtWNlhrJ+EZCzrjmN7/1woKI4vkwvYZ1c
lEZHsTF6bA5e1Q+Fjx9UCWtdpFrylpWDFdZAX9kAX3G4/18SQX6u6vAuwywEKOm2
fnwnZwGthVZdaUOm6qBJOKvcKJUWiN3nKxGegFjK0UD2Bqfa7qRkbEAkLlRsupFr
bKHoreHT2tVuAevnBwgxUOhEmW82bQ9eGGf3RX5Migx9CaUJ4NDjRy8kN/v7Mi0H
6HiWF9+s/WCESvwO0/Xn/aBnFFRAlx+POPTRif9ddMjrmiUOdL2Hit06WR+uMDrn
CGx8SlYHV3BcnVzARZNsRa+0EPccIVuvxypb5j6T1QjlxiuyoTcW4tycrNk+6ZKu
qYQ+9dfiqvIpD24tfvjRNq8dWObUSv4klsmSZEDZRuBraujJoTjxoOwuERWvMopC
FncBtZa/ScEdHHp78Te5VnjW7eKK10uote1YlKJKXa2k/uJbbw/2qyt/QG3fzR/M
dL7YM7RLMkpdXbNqjLa/wQtabPwiDT+IgUxd6x5AaR6dym319PJD2tUUjVOO/j4k
UUNP895AuUQPEn1phtcAjR/LKDndpevFQlIm95MogqMU+QLh5xULFfd2sQi6yDeJ
YaILeX71JFTcakx1c4L233p8lFqHGI4n9km1CWvi0E8i00wr5BDTB/9JZrRcjwaZ
R95hrdO125NGaSdnEDT9lTLAA9nyscf92mVoKCoK/PNu2AAv21tcGyNp2hQSIG+K
SANWo6yNrPctTmcfYmjafVgbdWN4ZLreYfcBDqXF+jSN/sRDyx8HdQ8cAo69NTll
8gs72lqR08ndJjJfe5ZrwZlpN41+FcTP+8H40WwSaunSviEZOreL3oqXByXOPHQ8
v5kGNSYGvWM8LSruJxpu44l1wwwYVuOV7CbCnq/jv4aLH4N2AKzMIQZjfOLvPuGF
wdfeg5C4ffGY9db9N06KkQBYS7iQ/loaZj93SB6u/cZxY88U7kV5Je7UioLX62+f
+mupwAErQ5UFDuhHixJvhGhXtVHsTYkrq305Z9r4+ohkVIhqxQEGN0CJ5gVx7N0Y
Q53bXSu1bHHviFniA4pQoBjTjYfSLRf2jQl2xOlB8HXw1Zg8xXaJzMx/IX86z4fv
0EydSpm3uiTpiZU/iGyKnU3y5NRgfOGGJjZNnqp5pJ4cd5wFzyMANCYDf4aB0ar9
X3g3jw8pFQBCrajxNBnf2nwqgsigClwUBjmQ5wCBpNITkGphvY70ejoZu55sqBcG
Nkk+pV6gpG5JUppBnovPLOHBSHyUOdRKC931axcN/KnhkdQ+YPenFhvRJqKEz09t
RwSKRAiM7YOMqLPsWUfck+lUFfisZ4yXk3Api4NThqpbS/oLtC1Ln3ARon3LdDQz
Bomfkf2xXh8Gt3CGJLTLgAtmW1+rq99V+E2SWJzrbcd1Li8XVSaCxR5ReVghRgzQ
li1zckrhmuyXmbHydmzoCl94dGTgha1R3QqBPQJKcKlNlgfxdPMQwa6l0GYRoneY
C1SlDfh3dKHGNCaJ3T1iTg4ixVrULKUSVVpCav0XYU1k5F6j2gWesljplJvfDqST
f6kK6clvN2xTQQt7AlL/urbg2kqKmydgfc0m77Vy8z4rKpW240QdFP0tGekNlgDg
ITNjmQA+9C5LpPqZg+hdRkeBRZTkmXc3vc0Ah2Whmn/A85aDIxHOBo03FDN/8obr
gzowCt4lksvis7hqe1jVz1I+uHtHDoyTk4054uefwKIfT3f0cj5dV05EHE0FS52w
F/afkvv6O8aMh2jK+6R9IOR6WzESB//cC0M17OCC1gZihG+Hc8J5nviNFmjxB5sC
NircycMxTiOORUm6h0aFjxHdUqRIF0LFuqYsEkvQ5iqDFPk8Gv/yDvpGzlAU3+RA
ngyj+yHv9hrKLcIqYB/5PC9ciDj/xqm+6vQrxeSjt5reYBtu+5OGDpl5oqJEVz42
VZDUuCbhfk/b2jnXTEaa4z2OR9kJ+lHG7BjW44p+Q5dU9eyqgtJP4GBLkulXDRUH
fNkIwHDrf9uVV3EM8BRGMSoJ1sGHY6T+Zignd/cqv6pL/Ji7H+P4nXjranEKy8jZ
gF8U5rFSggc4oVfIbMyKUllBYpAZaXVacJfXGtM3fFOmsiX+ogZkByUlGtS3f9j8
zc8p0zCMoW0eo2RoamiHW7ygo+bR6kkCbmCMtzv54NWaHr+ltLTyxobouUfrs/F9
3P/95QV24hbg7zj4eoRaKp32EpDGxMaB9CWqvHIerCsGun8GI97wyc+9jiDW2awV
LN+fFFvF8CbGK8y897kpr8swrrHvNTr1Vywd/lYSjhlCl2J7wl5l1kvR1hnKUE6v
eKcXbVJ1ytnY1JaaomBEmwcFOjz34lJ1OLSK32pP0n5APqKvdCXtogJwPWXgfTJo
y+UA9Ei48lFql9eFadwp7jVj5oCutgctCuLxuuz2Q7ZBRH/VGZDC+ZfANfBRgU+Z
F7lp7FZO5bI2VxS7sNbGld3K9aWPIKRm/knVT3ouyjVlYQq7/GnpM262/RkhYfB0
t+snROo5hwbReZu4bZx/Z8KcVmG9L6djMxB+ZmVOIJix8wZLxWwxYXgtupYMsDeN
Zw5K7wks0PAYNS4hJ2k2NBtiBjbizPbKBKhCDfzbnXtBxCPqFK5idSIE8hZK7AkJ
gJcWtjdRDEYYtix+elw5ghbjLv3zTcFtyZ3ehZ3gF8Ec3q6uEcMDLhj1LsXIUoSg
kCpO1re+IgvodOpfi3+UY7JwiZLAjYXyviHiLjn7Tj8FgzCgRDV44hN2hdxO+LZ9
BikLsmK6sxDadSRSTJecLZjwHYE0gId6UlOapgI7daHCy6U2PSmJx9B26+fqV8Y3
4SMHVpUO9dHYGtpPPkfvdLSSyW/UWn8cHuXhKYRUrTFIwyq8/DqZ8lr8Ep35y7jP
sIK5n9Yoi1VnaYjJ5BXZ1DnyKNVBazf6SoFcUJBH8PoqU1ut+AAowFLvjvl6tBgo
TqdHCJ+NNrYXkPrcUFN//I0AhGdsZhyYqgp42pb+ep9LtGvLjIuYdo7rwrD+YLb8
zBjQON4/DRFevMXwqK34LTMSQ702vQy2Kg++ORhwoDVw3e894/aMehdcA/ZOSBro
nu1ZJZiMLlv2uVD2eSojzR7Us7E8r8ae6di8Nb6NNP1npWA+5o4PHW4wlOpx9dbY
+DTxgMjl+cLI4Yjmq/Nl7636E5v3u2l+tJQ5xRLPOimsFiHQcaBViu8pCyn17N1V
J4ZjTpLjJuNLWcGx+jNuJd1SwFvaGed84aay4j8XRxX4ZOLDUIsQsi6tYnuWKj9F
XQqq9/v7g18yPJXjxpYACIoUlzOR27xGmSKVsiOxwSY/vm7ScARgLgW6R3+9U95q
NMOW74Et6BBP6JlI3k9xivAQ9fQYy6bGTY1YLiWVCfJecRQGfYpK+9IONfqEVSjt
KX2seL9hD/dSursGm0JDDYsAoqTOf2zg05gPnXF94OHFWax0T4OahpxzjbOzvTj6
Ic5N8RR9jen3rR7q8Uix7rIPXJAEWR3n+NgG/M4Qmo8qdsfvBMchVCJCUUlcDb9A
PDAdmz40ahVvgfJPnvph0+f0DpCx0ofP3SsUxtUY7CIVSVNNBlzZ/fi6oRAvVt1L
+S7BZXp7JsPWMK3XZk9c1I23xgLlqfwPTz38/zAa2mp8GzorT1IZisIwzRQBsk7W
W4AbIqxSSDbIZUyYeSwnGFqCtjwVReAXiiRzmwpbIqccwahSEaJqw4ObBgtya44r
q3cLexSIfV0amZCNxpdsa23UT4/3XajtKS6hqRpD83UKkTQA84Z3picQ8G42p9wY
jn96PCUznaIwRl3W2v7SbfYJaqGhsLNdlMPGOKMN4HVNFlZcbCPLA/+hdJBuAeD0
rhbYqc5SZ9fJ1TsJqBhy7CQNwpH53aqsg7MJwB5K879c9dmPwY9Nz+BAChmiE7kN
gDxq4jY0ncDMAS9q90kJYaYpdos+3H9m11H934W+IAeoRycZOChXQaOJHPPqX6Oh
i3KxeKZY+vsQwumwIF9X+DBLt0ags6ggAl2PRKev1ke2IlDNtDEjMcNR9RTha5pH
Al/6waKIsbM7SEc8b6GBzCrTaEtE5DX4NNNCb6/MCKz64mG5vYri5NcWd/QupLzj
N+0eeYrEDmACvSNSQtdnQyd6cgwc4TmmDTxYe/A28MMlopmkSTID25jKiZBUSZcC
dqM3yHDEVhi/324AjA9div0BpGIYh/QAEe5tkr5KU1W8g32Y4FReBrZJVhFqDeQf
7tOPc7u/ML2mwE51/FXENVo0Z6+e8cI1I+jYcjAoUpM4NpIYwZ5HrGhX8hIBSvV4
c7WHS22HBtrD9RGswkCnwFJag8hqQGq2FBhzVS7UUnLcVY1mk7+zpnEKfbqZ/Q2o
QJuZKWCohRSfs3RsSoTHraO6YfS18qJzoaAeNIeT3M85LC0oKm/hKosoZ/ETI1fL
Ow8wwu6FNml/38Xt8H2lQjVsryXv2ttzNVelvqvIbQko7Gf0jO/Ozs0c++e1ceM9
TNggNqnd46vOV06in6ghJQMoYDRrh6klWAAioYUniWSff8EEdpnZV7us0ISbcog4
s2YrDWcvlO0+eWkpl80weYwcXPV9M7Xb9uezYEhLa01/ArOGM4gdSmW4MUc7Xz3W
IL2jOOgsJd3qYsVQFm4aS0FGjPkPdDKs21/fLuWlT4GU6u5dvyn5AtNoRYTXJmKV
eEF/ppXji6Oq5BdO8bykfk5FpVyqPgDptqVqFoBubbwfOmhm6O6DjH9XP+GK6Mo5
0mxNHhO1EujOOiQAhnA/ffYtTRGmkQadEuUcNOLM42vVZP62C/34+tKr2n7eyBrn
8ovn0WpcCoY/exRw1snlH4GEDPGlEzLBTxGLZIwjXqnxWexEqNedCL6TE1BMjFfO
I3B59GSV6qpUSF558YBCMNsxIx85jCWIdqBORC4FJhRXbwKuWofrR9RmwzXFydYv
BhBM1qyo7N8y3fj7+iOEAu5B4TtObBoixzmpHBfzZsJqbg+6eAVFUyiGSICoXQlw
NNLHZsq5Mla7DfxTU8/lb4dGaBtgWJsqEE21olS9sbV9Qkos2RiZnnf2LV+T4pmS
TvE+HzYWRnBtVyiXIO/iZxKdJDYx13hucF8tRvNJRdUTnbKn7n3sHBmt1s64oPee
LSQcSnVhJA459ZeQNpFU7qsuveEk42HIqHA5gNuTGQrfIEfr8lY0Rr8AuYxJ0tCS
fSTYt+dLga0ZpkGauMP1birRXLaAQt460mEcOuXwypbS3Fkm328+HAuXwIzXXmo3
D67SzzBn4JnKeXCaxxtvrCUpdwop48o7Hwo+snzurbdwvgQO1DhPXh263AT9zpIL
Ly0BIzTnpzisRL3PFErZZMYOcqAWQheo0AouboWj3HQOX/QzgO2s/YcxKrT5uQ2D
udm7Cl3IbUsZa3j/xNfmv+9JQI3r25plS+H951E7r6aoHH3DY9DTeCdpC09RJv+j
VNygzFyIu2BQaE44pvi8Q2oYuIoeePdkfIYT6xJiyFtQt1GvvUmvM6vAz55nCF8g
hR5ZHmQXp0vMyaKjHoVWDgAl12m8t74onNCPnOubvbVVT0hb+WeXSUldLa1vQyNL
qrspii8qBON1GnbTJZmYm3LqXytRH+bJK5dTOWMqh54rBKEM2jCZ76BAyhWfxUi9
6ETWWqdXhetoVr0k5txJkNy0Ke1tLKo3/S7omwTvfdybcoxeom9QdLYajcdiYwvJ
HjjKXKqlNR4bGV0nQbMDlKBi0MFI2PRe/sMidZxey/s/5K6GvmpHUkomHgUJaO2F
aCVfykqWEkJnn4buiq8Xm4Ai/H+b22AnqW5pMArSqpeuLsh3TogaxMQNNL9kcTsP
K8LmlyCOuOdAMPsBuEAxHCE6qKMhBcIUcE82KVhh/rRcM3YkY0LQFxT7Xz4te6wx
d4rFRwckMwuIbowCN+cyM4HKHTeZFS59F0+gM5XnSxsdYo0uKpzrffDJmzlG8NPT
HIwjZ9V8RVrvlIo523JXuvwrXD+lMmt0fXlKkPAHhCy5g4vSFLPt6fnZxNWTzNFL
cD/uijMzGMuqTwO/Y9azNHYd462IWXpcNHNfPgMOVSL4svG84tr77U/VtVZbmufv
qZBNGRiBKZNkRtBwg9CDJPuF7AhFZtfgP+6kF14Dd0fkO0LHDQtxec1pL1VPvFrA
ZuWfheJS244yB+iIcrnL0yyNSl8VidGUFBCo42DXlYdRE2OrXLAW0orIt5CVR1Uq
7DZRdwysU+/ews93vNLV7ygtPiQCXWy0XF0g2+u6XxtAiB8yNYL7Q4tqnHmLTF7T
OwO/NE0O3Wn97vy6LbKRNG6QoCWdEecNzittnuyM49VmZ/AsRl70ja/ISedy0ePG
9t6TlOtc9UrBzvZ93sYDwQIsL5FW4F0B/ma0j/JbhFk1wAw+Ajqu/+8rluXz16Py
GRV1/Jt0xjtJm/8p3FJNXfacGqPhPP7InDtAqo/wMy6fvJEXr5e09zGvdKGK3Fcc
/TzbZMkdfyLx1KD8MyKdOz9vCMx1sV8JddNQMhKQCTsd9c5WbuGidgymsR/HAi0h
JWEfp8nXFOSZawVppTEudfeKEB1YPLdm34yKArYJURhsqnUFBX+i4NGuS4DHTt+1
d4IFYSKF89LrUWTTVfXM0R4mLGjlkRfWnScgkXfSElQNEoG9lq0/LsGPnjH4qDjB
asnjrRaU57XnQnzPULfDLImhl5xUyE5wBuqFuWBNmpoQOc6f2NagJns7t8XCpAQ4
ZD0KEhJ/5irWp+dcHS4ZFEZfj0MVxmdYbsCBAkfUPaJp56RnGQL6I8ppNJ+Ohbj1
jKKvqSOszu55YhOwIOInQ+Pc2qmZorkPxJ90OMQsxTqNfujFLySCbLyVIWuMhVhu
PrhgZZcu22BDBAubr/BDLFG6hnp+sO5Qz/DCFxWgTdlo32RzJT88Ecqegj8jGmui
oM+lY33JTA5plA1gFsqYqfIBn8xFODTHehlcqSLIXadytDgaTuqQl1IZVMES3PgJ
MuUHIdPRyuCx+NuNlzvssBNCDN90ne+QJelxI6OOyjhrj+rVN7HWRZ9BNo4XP65h
G+aBoNxLaBTJXAHef+QRfey2mF4g9zcxG0HEeK6jxwPkRFKUiHGRvzaiu71YzGKJ
Cox6+oE3QQNIe7pnqLGHVguHDrG+1kBaKDMKKAeVeycvivlipSCdV6kJJeKmIqfC
kmzuBqckprSjzddLaB4QNERK6nw1H+kFJG35IN8se4THK7/IPcJhyT682Eaa+INe
pE1FXl50Fcz+rHO6Qolw39F9/6etwf2a0R/NqKKJE+sYfl/ZJMFIm9+L+bOfRo4U
V3vqqamqsbzEfRaSWAUg/VIqYR/qXMLwFpcHUiG4bir47awpEzQJngvIToD1eoFg
Zgf2W7AlHrx21n1vAbNpL9G/bdlNmd8e4beqvTIDb/aN4nPcN1Ij0ckYWNAmXC+e
Z8gQXOICJqKz5o+gjSOmRHYsmUD1vrVfDdRV8SRFeTkBAtcdDtEQtcnHvv9EowGu
QkC5iTypM3Y9nc8Nad34nSUn/Veiowvyj7IZqeJTR/QpYJHFTj9QkPrAEABp+qdP
2IfVsKZaLtzbv6us8FWTxYc5aM9+HUMAUgz5uH5nQXFGCNH00CcGNCVFxZ4HYg4t
VWu1t7sLlVXw6+rKPCxLMgTpU+e+LbkCVIRDhB4ZpcoihBp5GHO3o2KYKs8xVRBe
TGJ1BrHJVT9FW/AyrGcTwJm3Cx7ewPlLtroTw+fMf2JQptSk0ewRUWQtgh59d9sx
o1tHeZv2TH37w/gbiHKrFVeYf3AhWh3uBCyP7TI33EOB8bmrKnN352NW4SZ03zOc
wq/EwZAxjh25iy/Wnr4WyhE62MkyNRIf+aXnB+DcRn6yoHlxMlsC1RsHz/r0dm0I
Nk7zBJFBqPGjEvQzmbCBe3zun9vyj4XWVJucGBID0aI9occT0kZPqHEXkhbuUnzS
lNqvZyD2aWkTRJmd7pDaEfYRXvzRHC6GnrsatbUlaNqIOy0w64ZXIZzyWnuolcIr
uY8Cs6k5lvHEdOOL9bZVxjfM2K5UbzT/+A4zkjWcFIGx0QPCvceqf5lPurzY33pW
z+gfww97IAv+iAVwItNf5DicUPSTon9m/wSzZb5oEWq43AfmEx9ZrZg62BLIEqLu
6uumvrlA9aRy3biIA5BNlCfUvQIjw33+3zwyIW8ZY8fQlvs4Wu2W0L99qBLrIfMA
fgglN9GstiJ+FuzILquwaBpLHuTltB7IDlfudOIGRmMUvZ0ooO6JbiXD2GQ/e4Uj
Jr0REKP5hh7VJi0EBNODyVHUi01RTmdEoyHl07XgUDuBSjSG5eHWGeMokXhU8Ts5
SDNwzKZHLTUd1N5WfNtTu+W4WvdyqNFeXCwDAcsrllhb0GJAh0QqswohMeRxFzv1
xjBHURLpJ9EOhQsx7U1tdG0JV1FUParyC0xoFFvAt2XLn5Jy0iVUVmY0bE7G3muZ
Zx6JYhPpeUqcg+2nk55hln0O2ICbm11+P8uL9uAbgOYPv0F12AN1HUsTm3hzOUXf
/EIlLerKpfm16Y2FvHkx1oQHIxkpXfL/FHR7wJtxmqzMvTCea4NWiom48rrnUkmm
8myYfPznfuoDGZ2sAiJe3EwqFtyalZ000tFHT4s7P4w4ew9hWOpRKFHV1b2VphRg
SEVtAihe6prxQgukQqh5ny+r8XugNZjgBpyUulIkoTL584r2w0PRO+RthhE7raKN
cDf2+ouoKRrIjHPM4b/WUjF4SyeTfSphx1CGXwo8D1gbzd+7M048R8x6aYfMn6U9
FESQMtG0bYFuBTrmt57bIvHbFCSFtMOAiXCFiZSfp1QH5ZrrZpBl9+yyrZ2ukdAt
JoZAd/LJWFI1qPWf4xVZsoW9LSFhiohhbn6/OcZFJ2YymOTc1rPHYMaG+ls0GOHC
DSPIItuJvlVH6iIm6Hr5gxBTygqgZLx6gl0tZrJ2MuYIoKBeuwFyPaewMCmSir9j
/JKOn+ljXkZzcRYVs3Vh9QKSn79UpGsH9UOS6dnK37E4EZN+gWNyYsvA6JPejbvA
GjcFjkQIUvV7TY6vFvZc9b0bKIwMwP84i9tCz9h6thpgyAxYg/WWbZpYm0PCpUmn
QYS8lA1OPDXIUbVPkacllvm2rSf9Jn+NpMBz5LtXs7AsEM5q6IaKfbwQTr1r0a1V
wz+UPUnEj7Xt6/efOce8qYGpKu7+LCclsc8aMhisFrxOCzktORcqKlitBtYERp9D
OSOcmso9FDhSI9xAz0UVMFWnsEgdbifn3wxIz3Y9qebmo3FuKYwLhtNiufKRGAVe
a2t7kVZJ49GdNyeQgF3E1SWH2UGlHWJ+uuq/1bDksQ/gFMw1vmUNt2Ng82F5QpyI
7Ghydx9/SiFB68VrHHiEqSP96XxhHKLnQUgd4VG+B82jFbVHs41LhVQtZhisGiGa
sju9r/FDvwkGghigdYv7I9aTslLhQ+GBEYf9v/5NH8nZVMyKYctwzfEQ+9dIW1d7
JEii4pNEpt8UPpQsSZwpPtnZmsGMMccktJCSR42MJ7yFvNl8dqojRajY4sTQXlHm
AJA0xuRgwAWqVLhiiR7KPkW9ydH7SARlC94Oxn776T9/XDJhj6CEy64QYhDiRqcX
Qyjh0glF9/YfTlPfmTzpiDVCuOe4qzIWeDdumiHMPiLXJAMFNHbx8D3rHwDE+hdI
jNDZWSt9FFKE9VN04KRqAWz3X4YUmn5+0WsLZzWXldTzCJ9Hqq+fTaHtKIVVgS0o
2azNxT/DPpPS1G1XZz7gClt0YKyD3tM1CM97eH+YKIJ6tL6YOpG5Oly9qb2IOgt2
W2G0tlL10euct9n+p7ByhXvBwMg4CweQXHhf8nWTHSQ+mqtT+y2WiKZfY51007fU
0omBZ6SYQwN9pogDVJ5KrcNUQXfwikqft3z2LCNIysrDfbSZjMF2oyI5NAQShWoD
X+AwbwdlP7305Jxdy0zncTY35trypSu7Mb2rFjKz5wG77oEdyfzKE6c4ZRmPcxjI
uVQ8qVvJpnH6qEKY2f0nHogxPBkxGe/G+L+XlZbslQyfnVSRooyryEyaJSzrVSli
cMt7oZFg5DL0vtYABBtZj+FdiRDiuruj0xgHuqwfaAijyChejTqRDzRZfwEHdkMQ
ICzWhYyZQf2gJO3YcNKPNJ6NzMMGzpJRfQArTRzQRlSym8SNMyJvLAM5C2uBLChu
dSTZwVzS+ItNolR9/ee9MdaZjalxF2jMP7j+d4KyzcBrxqNmF1TaHbrOBItvqmfF
JGZj+jFb/vnjqxkgp2RinX19AePswfjHIIJjeIHjPiIED4aAiQE7XQL5aWFsOBNA
qrVZjZb64c74Ir9seLI3uftL+7naUFaHzTFbeE3qlkC9HdvQ0Ju0+vaxAdnoscUQ
21meKkpjznkVeru6JniK1M26FvPoI9XYGb8Qo63zYYDTglXOx5PUCi0x+zm8Hx6E
iPLY8HnuBoFVzI8eQcV7N7DRVKWUNTTnRpMCODqgSvgDle5pgSuSJJXTaEtbnZz3
905WvnXLB6RYpsgU9KgoPG9vrpqezA/W0J3e3vEPG7jP0moGYyXehVha7AiS9wi8
foIRQVCWudqOeOq8lDhHIfzqW7EQ4/vS3EbFQdac8OObtQHNYb4dCPvHbDa3B8+J
GQv0I4itdY3ezUqRPptrmQjW3T8um49RbNczXxJCxDIgOTbp/ucV5zKVq8lkzR6X
mpEmwnNEEk9DNrjktm50Ij5QVgRgFxmeemjO40AIt2SPiVQ69DSM9quAH1CeuhmD
KQmit/y9aVfDkznqyq3uIuLvFclH6X0ene+YLba6Cdj/il3KBqgmDE4eXFziyhJO
k9fPX3VmnDun2Zoe3ni4cBuqxYrv7QRV04F+o9y5lprjVVqtiJq2x7jNe9x4BMtd
m2/bLsOZhmqq8aRfLZS3oOrYUklap+a7ghH+jRxksJ2gmuzMxoDsEBGVvleln9/Q
1ouikPJLBWvuLhMo3oEdI+HH23NdPlKWpZB8NouUrE3HppCzhOSma40txP4uBhSp
kJY4sLBpewk4fpS1iWovVFzUqYU3SaJ8r+06KNn0nRD4ALGoc5zMo/djMe8e41Mw
oSRBLVSFEGnfEhy8P97+aiG5lWf+H/9w6gDHAOqs59vusX/JIk7VGHmw5cDAKeSJ
ZCF0gOfkjpILVmlqkRKCxij+pmKNLLVpwilcFO9w+//vEdhEbjBFHDLByyMzZOiV
hBGerClwr+3BexrKpXVheSRURge3ZA1hBd/yr4SUv3KmLX9/4eryHYktK3PFY5fp
NILnSKwHyHI+F8i77DKjDj1gkt8ZdrSvzX+vZFmYBkwjMdkoZfF4zZceoj8nEeu3
jLn7Rciq0fwlfF5sxE299br28oJ8NTmHv2HTZ0LlwcEoRMf2tulZuaO/JVG2P82i
oXo/X7I2wm7+uum0xOUgKpsQY9MEPHtEAtPBuoT4I8J8HDtTvXDewTnyF6KZ5mXk
h73qPlqtYPz70RwXWKhuKv5opThmsX0HRo6cs625LaGhFy21lKPzDLTFQyJxDDCw
X4xfo4JwGWHHJ0HyysNKad11JADk41YQhAUdl3VKwea17GXnWaLFqe27n800oDF+
Wn+QZIOgt+1FGj519AO7Zl9UePaFF/BMLsCEVerI8wvcrxXs4uejcaZIyOcA2v/+
1qR0wodlWACa2YpHeeO5TxdHNVYGdE9rMTBajE1fPO62pHuTMyTblWclJ9S3dSOz
Kn72u1xX55BKqYWNjafXCu7L6lMPtlOKRySoplNNJizwc98P++Z6Q3Goc56JWQGl
/laoTyuIJDnl9n35Tu/RSehodc8y5akCHS6J81suJINSnaTOmtOHP7HYik5flt9v
t/654oLSukTi9klON7tpHIvRnKsw546HMtmOtA2EyI/0YFfrp7MOzvOyAmScGfGV
Pv+TjtnVjR0R2AYzrDwP58X8TrKEJfLnCykLvKXcEy/xeqH5dyiq8yAveEI/44CS
Ukvz9BfE9KJO4LlxNL0kqZK3YN1Cq3RuGOCLguhU4pwM+4ARvefpFdz+yWFQqhOS
PWVwvJw4jT/QSKSkCRoLyFRN4XNf53zfMobcWPieUSEEbWNLdGPdUxjEB/+NaJNL
JUbK421JywcPkbLJ/CLtb9GUpZHUimrx6I2vtPjWRF1T1kXG6CWGg22/ZHnbi99P
9PYyPwFcpWyCR8/aHgVQIWp1bh29M8AtY5M7x+k5yZPKPMeGpWj6luJE5ANWRH4i
xhHUMaDUr6stJVh/1rqYoZvpAVA/tvxRpmIWZJjCa/lRXMRLfmq4tOznJEXO6zzx
hbPY/eNnDlBI/j/P/+RATeQ4Ls/jSVjRky47YT7IBzZ/oZeCOpSeeihdNQrFZUFh
s7qMsNW7mdGBMfo4vTAJ3oQoQ4H740vtDzY4OhQ28Jt2qlAcC42TpVBnooVLflG/
KQxJUD8T7jJicgyC+gPEJmnut2VzhLslrTbkSLt8xlROPqmXs0e1zR48ZDKf3EHl
baWLMVje8gjC8XsxThrB5fVbzwBI26mUruqAQ/siNpBFTZSTZfIyZzGvpF8mnOlN
G/gpsNaIeV/omo2tyPrxhYa+6gxd96rXo+xgTPKJDP2vkMeM8fUob+WnNrPiekYv
9/PSycDesG+tAA9f+lqyhRrq+UBmtYjtRVl9wuHNLGkFxpejtkE2yvdpVtWxx3Sj
RxI7j7G0AAFSM8L/VoPgvZ458WyMLHgP69xSQscLNxB1LxfBCNnPSGwZKVjLxpwj
hPSWK5NPKaeHikSA69mmuF9nQI32qiSq4EQznJbJmg3lrDg8u20AYy44j1O16Yi6
Aq+A4pHOnX1l/66kzGEyhPrM+8Wb55YvEDoWpSBB7CkBJLVmKmnPye2L64BsyVA/
PvnxBCHVTnwSdmvGrzLv0o0F0flZKrrowbEWZ8Jd5OK9VBDL/vF8mMsMv0zvo6qp
uHXpUcTPcr8v/lbl13mEoPV1Umer3hwx/lkXh3hctKF68RN/XXG5DudvbMvGMjlV
k96eFOM7fe/ZdvELXggkYBBscdO9VaEKwmg3T4MEmO+OJmy8CxMNeP0NaBhi2EiD
ECNf1siAA0ZphfoK0zVmoL120RqAN+PCt9PFsWnlLbQu+UB7lQvxjbbZR+zPMspy
UFK81KKrEZqFTcjSWt4Px4Ox4iGlbzT3pCTm/TccZKjIY8Jl5oMRdIrdpmsKMrLW
F4zobwJEYzPv/KowV14/eZmXseXDccZklgOiHpfKAcdXd0hZoKjCQ8QGWrr1NTVv
Gdop0usPHzVKliXfgODmEj1nCP1kRIxmdYiFGF/7FRs5UYhaWdnlfdj6E45AFadc
4TyFc6i/XZM7h32NmpqjU2wcAn8qKUNFSV9CzNGO3OxQvCjagrShRdHME6Pja+op
9jH5w6suPy1qMSGsIVCwWHufs7ECILd1b0dCmZlrWCYlKGVSdeIOJWMmue0PAp0B
iZoPqdA1S67U4KJ6Alolu+30qgswpwRqtAH837zzgfjeOjG62eADMTUl1vSKaiBC
1BlCmL73uHrWHv9VMdQu0Y5sFOEwcDqrHeGqB5CgLlQu/FnacoNeOJg2aV+qjkEB
8ezVpPvYybztDMqYS7EKYT9Usm1K6CfjF4gcRnxqF0JBZecqkfJ+W05HIY7MXYpo
wln5xnCFrcfT0/vnqdM4IVtIXNZ/mFzm1QbKb2G4aDbwj5qCFt1FEI9n1gFFLjs8
/nZihJslaUeQxz3kpOJn5p73SfeLdXlqHkwB2hfcP6qtmTtUKFPvolOTsgPr/inA
CiIfYNavD8mRvwtZmJmhx8xUvAUsMTrSZZQKUqMm9E4rkHaoSpUSYB4AdzW81uR4
fq7I3O7jhBGVvx6gN2W2480yh9vjRK3Xfgb6I5ntE3HF3gAvpSj429HrJHoJ1Vkc
FpFTgco0xl0LsHaaSBbqELFK1CwkOGBUYbm/8t1bMV//G/EyvlMeNiAiI5pi/P2K
GGCC58zSekneaQEWPUl751cQY/RqbJdeg/xpVtFcrnxR8cwgt2EPGPA8iodfq35X
zcWfzwD21RYytBEf8qerFaAgbS7IzXpQ2SJYdF2nL21MUbaDmhDzL1V16PKmOL1z
dY6oe7AWogni7QZlM+kXCmPqa+Rpf7Y1HsxB5XUwHOF+JWinj4bK+NW0XMyaI/F7
8KiqT+y8nqNT0wKvZDkS4zQVb8WXpq4bjBfzyuOpnD/nT1JGhaRWZMriMmmBCtQZ
MAl/Eth5AIip2F+AjKCcH6WhBLK/E6w1dzgX5UVAujDhS7mRQAVD4PECp7JfzZBs
7soB45jdfBYyB9vIvAmXOOrxa3HIA+BxnzV/E6uTMhLNE7SlqjCprEtdoat8zsBy
3W//MYh+AJkGMbQJil8XQsZkZcYIjZs/4F/Qa8WOdD4ffBmdE2AxqBfyNtANT/g3
5SlSwm7eAxBkkUcJBGRfKThPEbGKMMzML8nvLEMKg0QryFUoyZWVdrFW3pqhE6rN
b1qgL41X+Pl7lSw+NfVkrH0NkJQDg4X6hdYgKIpxKS09JbKo8hFJZva8c3xfO05n
lgIC4ZYHRYfEAtvJSTOn02By6pEWSB96waCoEPemDt9hxzddZMdFcKUGujH/Y/iC
3aAq2/L8v8YJUcM3NqvyNpMzLRewT9ZHSOcOI0kNnddem3hMz8yqF+8bufNe0yCo
LNy6OWbadvWtx3/ttFVZeWn/J/n+oF3DVS0DXYO2je5bVYACr2QAKbuo6nRjTT2V
xRfK1oc7VzCdkn4rlKNS2XxFcyn0GpOMksiiIufRWnCewGgPdSK1gIu65bI5htlp
/0E1wJkc1OSS6+AirslvAheW0WPbivT/Zf3ueqV0pg9WFXFa0Adrw/hlrituKM21
QXDCuL1D+4YPcXz3hhzU0XWyql2YklyhEOvp0SfxvAyZcYr3UEYWcCj8O498rSrV
KXowDoiXyIoZqeuZQ5r9DDo62qe3zv5vAmkHss2FkjqoiUHjy4frgY59ConjAc1I
EEQmei4vDa/5CjwzFJXd4fhQG+Bm4XrlzdhmI05jVuVKeWxD1BEwGTLsd0lSgQbj
QwhzEEb9AA+OFZjqg3JA5gdMb2XsU8TS58ttIU/Q/zJg0PnB0asWfsYmQKqRa5iz
RE0HVrxRJxXgMMKRfk+1UISapxiMo94Wewi5Cqd1tTbZF+P6gbagU8edFBRA37cd
DtPufoumMhX2mStIXB5E/hDD2FGamw2MB9wL1x0AqSAqoFtMwhdzogXa/N+amjbw
X3NR5/Orfd2IX1CRG02ysFN2H3digRqnbIn0w18KFyZJ/bRjHeEDl4O1QcZ1vxDq
bYyVBtLthhaZnAUn352JBynvBXxhDeLKugxyXpAR/yFk8jmNuzD04VdSAdGt7F/H
SFWoJHV9IzHb1C1+z8gMzvsQyi7A84CYEZ3aDVISIuthNt+L8omWAtZ+CSJhRQtT
FtpfcNc4smrOjTeTsmvbSZqaZBgxA81dtmzvAvTBUy79+kZIjPBef01NfHoAUEZC
dBHbFmJH7J75iuXQ8wZaaky5W9+wNnVI4bF+T1WWl6spF62j3dQIwQwa4ssU9FxT
FB/oPGyhefU27FLRmw2nDo5xiM1VEESvrJysCZ00Ac5HS26HW4XP0osgQElG/nxR
G/etZ6R8CVqiXoRp3v/w02Ug1ns/E/hxIQ4b2PDCAd7r1t6zaPG4T2uYH9e+Ibvz
HRGmkeT81lavtJHZXrEjpuRj48wPy33IaAhU8IozhJTX87KM9hbOpOw8Z/l8zzjv
1mA7rJnLkUL8q+LiutoEg8Tt3oLt7hpWMxV2pZHCcCvmHWKhtwe5+mT2BWNdCXVf
fDGn4LkNYlt703xG+QxpBi1bLHGzE/qg3molPrX5lssOOm3YMJ/HBgM/h7wZazle
LFzqjgdYTpLC8dSHHB0BfyRu7xgAw1j7LzziX5qpMkT9khThHe0ibB3Kd6Vc4Rll
dpp4QICURdsnb4mcdN3knRTK7b2DsW4y+BZAUHumD9MhKEY8Fnqo9vJFfsNjadpk
b9wnuDNmDJ7ZSKiEZeG2JlUKDHNoKeyLQqYxwLDrGG7hoC2YPSOf0Sqy7xL3iUrp
1zB8JI4Zw3Z6MAG9ItJKuIaXdqE3ESRGG1T45b9MGw6uNFJ2rTZwzgxpagNZZwah
9KQ48FRPUiaAzn5zQKKIkUwNiu9XWG2bLoGT/0fFECgcVQ7B1Oy+YEFyGP5biTQf
kvThCwk9SZxLpUjYWcGO/n1zVqvRbgPQlTCzVS1mOYTSTibWr36MBdIphuOYuzXL
U7TlWEXWvf6WhQr9cZlyT98OjJMGiE43eJxTdKZfHnw1fqB7IDj77pML2PSzAs4m
xwSss71bUFSZ6AEhiRXhGZeyFp89sq3hmaWu91QHebQ6XAvyG7YRulnCbA2EbitZ
D4o03utIw5NQ+xeDQM3xCZKsRsmCRjmF4RaWImOP6e9dp5fBmg4U0sqrLxlTex2w
ShbUP7vrcN9A6Dau5kU3X81yjo7aa6pjK23pu/5+lqvnwUfdLOf5HfHh/hYHl01B
z+HGc8UEhDp6qZvWoIr2oe26AaBCQzUC1jHjE0Vio3IJASmqqQVZfhg/0PMI0YAr
hRaNdh3t+O9gS9xXgRw/54x1N5Fjxh8N9zJIG/cuuhk5HHZ9K0XcEsGLro+TsqVm
c0RXj22ykBf6Hs4D1jzboHrmkKpNstmkfG9aN0f0XrDNE9+lr4cjgNv2FM1vId86
qDwdbgwpX/FDlYSHJCEUybZGCwuJtqGVftOVbT0ZnXJ/G6p1OUrt3Wu3+Hp8zQB/
Xl+N8MfiM6qynAZxLW/vOwslb320cShlZNQF/ofJIwkwsWUZxJamzaFBRws7ZS39
nr94qHsnUX+wWM+BfT2XBn1sAdONzDaZJKiKqLAjxSYGpPZGMx22KffKKGdR1vWS
opw57FasYI3bXlny986ua60krk/SrJuYJq1eUHOqS2gCCels+Spo+ClgHJxA7VGW
Hi/dgC+DidlVHo3D+fKUQJ+/3ojoBuOaOF77fjL0rvB278/qyiQ5e8B+kRfsqGHZ
1kM2eVnznZhQ5EgS6sw6h4Tviih0BDAXVezeBHa808iYEZRRRlHPZpbnIzeOoO4w
FLTBbOh4mtvr7ZDYatCYUDnkmd08Uhd9+U8ruREmyyu7fYkbB3pupth3EVOJjoXC
wRdMXpa+0vFPGzjqUWvK8KbuqDoy9FGSNSQRCBM8jzWBixii+AM/vBMrVeXZ/DZr
wMTyXe68PV89fWSqtM1JKHM8oMwly9nhLXmHBHMR7Dqsx3hCrv5WGsUPe21pfXrp
Wti/x826Wt9YLHHMyunTCSNkjTCdvdULy1D9tH2YtU07dPUhSCWgxfA1nLAEs0sh
wycdsNbwCbRMFco4NDzNUwKnt+HnCIJoV7Koi+L0gQwcmSdT3lBtZZo6x6WRdq9j
vxgWCAKE6kAXSQSUCEt4L8FP1xsjkmUWpWQhtxV++l6YgzKzk+QJc3daRgs19qUT
rx1p7cFplKYV9mCn0vdbc8o4nRZU7VkEEuu1wl64vt3xIYcv5qG9uvbQtYtg/lfe
o84G0yVvdmkAbmm9JODxzFW9iwPqQuS2viDII5A1FcK5jAItEnkZrMDfw6m4Fm/+
HaIzw0m9HwGlsDCbLrkZKSMHlxMmdcDWBduKzgcMWgkZaMGnVB50A3rcOkDCRoIS
y/JzzwGjBTWgl6tXgW1HMhu1AWYdflLkjC9lk2JBLgnMZY3iap/iTYozkmaIV78N
79FSLd1laiJ6FK21P4ZffmCZcjYzgkSbVm780/+I275FCFeLiO77scuug6YhYvUg
FZ+kEc/7PtIMfI/5TtimOncVxP6a5FjJXB6bbO8yMCCbi851ueOykHxmeaC+RO7N
S27R/ZB+fgXHo6HvYHnMtKRfNUvabXT9IHeAggU2VavmY1/pkV6iphPqsBHkKDqk
JwC5onpuQpHPyAM1tu8EaJGNy6VN9CkfJ/nIDgI46iQwiMdURnKM3Vjc7WGAIEYo
Oz5xrXQCKsvVKWEl2Qnq9b+c5b1lRZTUGXhWiFn5tFVDJqF+38iIm9YKQKtsZZgo
iFCDK+KjWTqTI0fFJqEcGMywaC0Roim7GjNsRbdHQDSLOvDSk1fUkHaAyWK5Del8
ImhGCAXX6G3JHBfy2kSu3pvmEnrHDMlUmZW7VK1o/wntgSBvilO0Wasv9DwVSWLB
7Ag9yFD2LTUk8PlZbl8kRTWaQRa0PN57a4oCGGS27n0ZH/X/rE0u5VFDRkm02EJX
8LANcB4AYu1gRv0FX7vK1qYcwhfXU/NYHeQhIoD4w51O1mS7BRAxMPniavehDUAS
Xu3B3M9F82KbMGDL6Pkl79rwp2jJ6OwCNfKT0EVdAK2ip/R5rOnp53mVTpcEJoJ1
jFVKFTeGsjctPA+X7WkxLwv5R9Mf/ugF99mA5SvRBdvE9ikXgSypH6TW4vUx1/GW
o9HX+LHAIVdt5RJeDkIbfwxM44k/kYkprnc1FNFkm0298cNMDHorLWjuhQRXRn3i
Ku3URbJ7a8rd1VHmKI75VdSmmAFSRT9EuPPRBSwrgfo9otmi133dy9ZkHsq24gxz
1ninFVi7uL6UdHoRbarovAzdXUXN8AcpM7HtXTPQlJAIGlTqCFYi/ogBi/XScQ4J
hUZie33j6oYUQ6bGcxXTFyAlQIgJ+qja3TYNc5K8pA92wxNnBIRQ6Cq5UtoEZuYb
kSKHHrA7TnNqWgQCid22hAHg8sdFJVYJv3QPnJAoPso3P0X989Bhs5qnCjy4CzzH
uXJ3vTYcMYZ7F0uzwMUHwuSU/OS3/PxUIoEWPYWbjWz2wkbIYJj7k6QY3e3LDPh/
A/jbiI3PF0V42EOXlM6+iLieKxngrVPdUud+dbPJ0Sl2YF1mSdmT18iEPQ02dlaw
rN2x3ueCxtwBrJOZpexMR4rQhKSy1Qh68LBHGtlXXD+ot3ZaJPj/1BpsuvhSok61
Vk1kx3gzSI7EQKshvQJjbmdBcj/sz6WzP/xBrZwlNqOk1brTTjP5/BEithQ6IC0x
XoKwf7K6KGHHE311K9CEW6CS5gHbwkohs+8nzpR+JGFN0O5xc3t3EAGtjosjPgJ8
CUtA/2XaebN6xdge0AeWx5LeORP5GgZvsn2tWIfR3dVHRZT04KgryEadORh/tJPv
LxD5RCf4ar0qNSrvwb45+uBq/AX0H3Us0C9nN6YqgMVhPqA2u8gEe6iZ4V5R64/Y
QUi8DEWm8TIz1VpJCWXBFuDtmR6pLELwSAfdk69KG5DFKcAUABy1S/5PSGnkg+TY
6O1oIPhTzUvb9lOTfhsA17BOozseNAQuZKxz7TNtkM+GrnC0waOr3S3V4ye3Yd4V
s5gjd9MSpSbvFIdcVyuDCueAZicsf7maHgCy2Swz+XVP4N7Rfss11Gan9eCPADP8
WQkRr6J7FSEmFQ8w4qviVb5v1c9qG/5/p8SLsW0kast47TGjE312Wnnmgnu0sUSk
A06Rb7wFDGW+soNbC5YB8qOrIXO1S1GElxcl2IKK+MeMUU/O5a3RIBpfXgzia8/B
oXPLvrz7xEq7rEfR4aq+AwuXjEv5y22b7Hvm5jHyED6Mj7496kEJhHhXR17OeM3N
Ga0OXdz9fGjBqWRuN12wAc2flJwUzLAbrNVmDnMkB7VXoP04iEN6MjEREtSr8nd6
Kf+hk0n1mAJI/MeFpv4hIdKGgY7sYM+xe+s5j8+amHPVymgKOdoDJ2Ef5PB+fOxy
DfOBcuoStHEw/eds8OXEnL9z+n8cJyHSy9PXfO5obRhdnogvuyJFGe1yo6qmdT33
VGgGZrN7MLt1KIs1Vi53LGoa03UZpqHLSujcLgNHUFbNJqz34i/im0Tl/W6i11ri
qPDv5gtbhNJ2AI9pf/0hKsTFA7z61kCk+pKmdUdrsMlZAp3JY+AIzZ+vaAqCyFoV
QLEMX1X/yulJfks7sGOND40CQJVxvHk2s19qqDL4Sp7jl2AZtlS++x7G7yudIRJu
g+G3n6LVYMKX7XO0xkmtnwdDAIhp1f+IzttUdcfqygemJgw7513TSdex2A+XvQKu
T21VB/O7/evBkss0hYlFP91pP5u9ngozRsVt3/N6kiOz0HSkVICdv7YwxmuKVrcK
ElrT8dK7xv5mF6kD1FjHwj/E/57aJZ2EGxmzndhvrfIh6s6t0dHIz1Fyjg2BrZhu
VsBM+LgEd9Oj4gG5c1syg3imBbjFwXysAH6mkQAonW3vGQeJe17xskIQ5svMVR9+
4VjntzY4ywlfknHEzLj6zxHINhLCRwkK5zaposfL7sGmKc8FUi6tQZbfQfLy3d/W
Y3hWiAf9ls2rHSjFxc0yN7vKEwa1FPE04vABX6KjGGlC9Gwe48YK2AhxgdyEusFo
anIJT5UqBVEcZygmVhc4e88luecIAP3YXfWMOTjWUjH0qnmOvtJFm8ITwuiTF/xt
4lQEdonTuHM2u70uZ7zcNh7XAni1bmgNzG9abUXqTc4DXb7rNY+TZZF0SCOL65Vq
mP5t6oPfPU6oVVuIJRCBb9xt66AfzznbxE/sXR3bFsfOWD1QbX4l3GRS3SdBY9Q0
nZBOeVgVxSOJuGi0v2GI+V3wGhWlALoVZudnyNt4gK8i+AqvYYhmLJc7PJTHOE56
nSXBCah4LtOXt3rPyvf9CcCeiQ0U/SzecWO1Q8f36zpZEN8J+pFUqt0VyzGrNnlC
pI+v+fpB4Ky/lM76QmZWwaGJ6tPY8q7gZl+AMKILC6daYyv9G5aPzM8Nv2zJdMZ5
h/Hf4C+UgBM2bsj5+MN2hZWuXNhZpJUKacecaSO76ooVcVkixwqCtxpoY4U2qoP6
m0U5VWuWQJ8NPxyOS32cgqV6J0vyZC46Vh/QWkafaK1yhUJfZqWJc0qPg7U3Au6x
isoYjcmxiIwRt3TvWmbvkHT0MgcqEcvrRYqtz+Up/1y1Lan943cc60Sslqb4kmXw
Qy+M5OrncFJhwHZ+sIPXmlJXj5cD3F4LrljzrbdAwIL65KtwfJB4CLic3x5JqreD
hPjtWclayhIL6bsa3hJDMCx97vvGZRpwHW5TxrDIY6noMr0+ALCVHwCuaqBHcItC
ciZf891nbpvB4ACMMWDswF3l3F7eksBqsZ5zKEruy/E32Jfi1w6pmBbDusn3faWd
k/FdnBV+Im1f4hVQoyMvLtU5FnPUn087/wFG4TR+9Gb3CXpSPGQMddgudqnpthjo
6T+f0rkrAZCslYZm6ZESbj1LAfh7hRuDx+iE27TUHmWmvEpb8HKQ2/9zfw919Be5
mZcsDbvGB8bl3pFAK6G0jfumaxt3Op9BOODtjjBdrpqKjw2ka4vafkFzdazu9ru8
Q1QJnc3j5UWSR8cpndp/AqIfcEPgHcxQwLCod8ImlVwWVY11LcU20m+op7onJpG3
6ofi3p5UDHnJ3A72pRmpFf6XSjl5CyTiz/jAdlDIMwG3fukZvtAXYnQY/wywMA22
ai2aL9LowsIO/hj8Tu0frzcqYABapJA+cKsGwiJQ/iFGa0SoTtReUrkz+tqs4hfO
hs6qikAss5dLBpv3hRVzVXW3uyT9sL+q9i9xHmNPl2oT6Op7fjtduecy8t7hcDiz
MpQ3lUWmpmKLdC9tyghzRUEmHaOxxqu0JTzMkWi3KrprNFr2059iipeBeA0cAUhZ
0mZwwzVnRgINnK9Gk6LrbFkh3FW6u/ZT+mV67wlvqhwo/JH16Wxnm6nmaSCE3lvC
AHovCbJXCAL4Ioxk108DbMnsWefGjN73jpxKVm0vYhpmSCiJmVCibSAsP5SS4buk
rV4aQS7UspwQzSWzGrVq8JlZvNxWDofN022vZaPgFARa9dX0FwIQig/Hp1agRIiu
Y8ZhkhMCUW1uuu2CcHqeN7Jlt+9mW4midu8r3cVo8t09XsdNqvE4KNjMd0RP6DrQ
OMIrFH60iDJGlGioknDmy0uwYjpiveUl/pWF/NYOyWJkIvh5Ev362HVBRpuRsRgw
aM5yBIRetHUFU4+zILnmlNVRxrjuknta2LBcQB4OIYKmjyPG/SpBa4QcAwCWFHMs
2q7JIPQm3vno2m7yiB9IsXS9hzakbQ8NvFpwsSTf+maZWGDIEYxkemTPW2L3GHLT
pn64tSj+gIeAtc2DCujL29XNMmW36kFdJDqrFn6nKPUKn+nsu71n8AmxGTXaGTLF
Zbg9O/NZuSSDvlshYOlmlyITCoo/4NVvxVe8LcULxoFO2P2n4x7IaJzfKYY5T/Lk
J5/iwFR1njmbYTY5B5F+LaqzEzC0zLQSWWdFp685OxU3Jl7X9k+NDS0LzSuCjNSV
k8dHOZAVjKe7nD8niGUEx1V0y4PIPBAAcfcDe+t401DOIqRIi+UdLMZfpSVVjiwY
Binas/CStScQHRIXOe78Htsh8OC9x6+rnb+ZFaBmIlE9998yizut59vC4F0zCBLy
gkVfzHOyF6aPOO3jSEHRDtNkkwZM+GDitBQJD1rJk55ARZq/uSot372l2kBz+3Ba
/MbKuj3A9lFvWoXFCPa1dQEDaRDqI5oOEldfU26qmEVs7ZVjH/hnXo5UNan5/cbk
kLg5gRhl8LhDWemTNk2Vc6FGCHjGOZpzGWY4QRfZME1KoJTlTBa0EcUt49MgbUwX
p8h/G25fWuzOrU4zKnnvFHOLYdTA6lWR+wdxqXES1LsH0afReE7ImkPsdj4FJ55p
lDNldoCHZw9QHQIWChb7XFytsgHDANqb3MChbfLC6qu3azKOV1lgjrdX2rzUuPl6
mE33N2h/dYMvKOzXxMvjDc5LZtaTjXA1zGSVeZLmlQm8AMCrCvJClITNBPcowJvK
aq23UtT3d7wz/10x7VYxgUFcHZznlZbR/Om3L+EGI1HgSmew/UTUPGoXCqiUwh4D
kt6HmcafoK0E832s7HAKGc5NJB0puPPAK3V7fdIK3J0xUcI4uVf/8oOJ1LwcOdoo
2cO2ChBiM8CcKuqUulRbIf7GNsU4wEbKmfiol2xLzwz72e03bBgfrEr88roDQq5O
K5QFb2eYuqTKDKtFWKhTFDE8rF9mQ6Pug0M7P/cnMIbHYmAbxhLcINUmNF8F9oZR
o5PFcnq3Yp9nkDesGkhkr5KjR/cD9WTurcDPRiy4szYoscxiP/KD3VY6FnvFQLNi
hs/eMrLPtJYu1SYUHOfeeqJeWz5y+I2jiQFjQT2IUXn+jQE8XLFCKiz8vZN64hnu
1fIQfShgpdvBHCzIeVimv8MVu62qk6//UdxGf3LFdjGaZc1zQDFMgKet4F2KUQ3f
hdsvXOoW67LmI5nGlYKPZIl5Rjv/ZERciAP57t+Fl7rVb+IzRAt1Qp10EMdMfoc3
f+7RpGPp6zS3NByCa6ApySs+nmmelry50UMuoJl6s/3VgT/bs0wPbXHTId2Nc7h4
V4/aH86ufCwoBUEvSgYoMYuu6g8BG2nFpEMp3UudfeCXZXJGGfKdvrLfjsbul25i
3y56ODxTm/GT8XPd5hGbDIWuNLcBuSnNlgFysEqCiZoe0fYoO9qlgTg4mNBY/blP
kLiN1tVtKTDvBF74KB/CdHr9zGgISozr0DweIUq9kxGiDl3szc+frwInk3D3iYtq
Fw76pnq1qZBUnVqb2xyOChjS7SyQixrGghulxXzZhNXJoA7vRYhjIbw/daJ0xGVc
PhGyX819hx2mIhSufT+B4hcstfU5rk/5oaRlU+Cd6DQeGX6uWTU49ISGdnmvRkDC
zYwQJe1g9B4R+oOi9N7Q2sqfRJX/sM6RkJH3VLdG0EZbCuz9am8JiuN1YvNvR+ur
mbWJzQuUBBrCfsXibsOj36qd33sowsxR/i6KGo+9ZfoHZCb85eIJVK9cDkgq5j+1
C1LIXPUVzNUWSkfQBgVEI6F9ij13J9Y4K3O9SHDPRjOAyof4+f2D1lHDlf9oXZpr
LYzrqIinl1qjGT9gdyPDM0QE5GRTcRnP+0+4tPR49hmv0j1BxtFabl7OYiXdaufD
bQ+PXs26w4itq9e9yToESwJAX/6Hd8UkcVnjVPqDien3b37EucDtQ3QJh2exczZ4
uLPWeTaxqwqbvo+m2Aalc5p38MO2OV/G7gZiNYp1CnyQV67fdeiilOjQffKgFHqu
luM/Dy1358rbUByXzkbjJruBp/aRC6CXp+Scm3fOxtufLHRRXArFhPKz3hp1DyXf
NFffkPBa91b36wtsD31IxoZaMKa4tW+EyF0TQ/EIO+raraIRUYjeDFOMA6D9PezQ
cRHrQT46YDywLwGkYI5H+epPqQPtg2X7MzRRMZaCWTkYtv9y19o2keuLJrphA4Yx
I6yaBYNsD58+f6f3O8MFogRKNYTwRTcDLYMN7toOadqxVuJbBS6FjZcPXy/0XL6H
AmcXTQLtUHedwjs+aSgHmF3h8X1dHX/unnZ0TEZOCnTJBIIFdZMZE0SvD6Y0zIIQ
d+KU2lKcQPPMASZv2ENqwDzpyK2NPp14YJZCfHgvonrv7A18SQm+DA1dGsdBiJYF
pBpm+72jRB8/oJTMPCjl+CXG7PzxyKd2SdomdVM9LnJ/uilBei5rtG9khyHNrStW
a7tsDVP9aUxMQStHt4gnelw+Cof2zefO9dWlpyxly4pZFSjZc7RyYvY7VpwG43t1
EOMnaJvFTkwwgdAA3pANJB7FH7lJV7UDbp+fO3k1y00N1wdXxmSWRDV39HR7GIjm
xVrw2LoD+WXOmuWJq1ycjx1/4QFFIyu8+PB4zMuzH6caY/V4QtAxt/IQ6H4t82KS
1sHGnSJf4TOO4TaMbqR+/OnXpUtBPtbwfHb6wPo99b0TxHE+xqKMdQPuncTR7aLy
x2VgvjSGRdtH+2a53gzAZMZw1zCUMZbFNy4HXltPTLYqQYuiNeVpVWgaGdyLoEs7
roaGsbQ6itob/d6BjDTolek7742dKsRBAOwtFcgRBqcp39pQ1O+BTRt80ldFH37K
BfN4nsCglQ6J9sK89VODOOy3sTmDte4cKS0op3dCUwLaFcFDKqgNUy5hcpAS1aGj
kCxZcnZZEJg1nkudjtVBHRTMSetXWHYNw/8XV1Tve0oHHZpon20T7yKVRuNT/MH2
lAdzn0GCOAbL17Sq3p4YELoNmjTc335qLxnGyUCU+oID+Id4TAGr14WN3Scr2t2D
WdNXG4tL3LRfatOfJom9OCYk2ERjbreqOdgcIlCdwK4iExEqrji1HLnWsBP6DW5K
PU2rxakWMlLN63D4tOlHEJe+zn2f1RdwFRkQgzF8s+8c1FrwfGo3gV8FMFoULWyj
dyrj0PyUswa2Hqqso7c2u7K9+JAqAZJVu8gvnW53dT9PuTOQEZpfU9fEpX5ucGA5
5hSSAVk7Sf4UPbuGgs7/KgaCOsJTXjb3sJK1pWAZW2jnU/rFMYA2xSTzyvXqSzbD
wC4dFq9pnlDcccRN38XVw2YW6c7Spp02rOogUDJNB0yKQ0MYYgsmEuGMm7vxQ+31
/dOjlPd0vKUiiB10b2PNpIlIDUbFxA2KoHEmr3Lfe295gA/NRHvM8kpc9Rtg4OgF
Az7VVwFpKtwCFG/ynxT6QVm3vdv+ckHndeyikaNfglGsq+081gdcJwjwuJwyLmyV
umYfrdrUawyIdrsr6V/AjLDIaDJRRM0XVOaig93K7pm+ln5/4AXikUuscD4MYy0x
7ZIcSiuISQmqDNjRpSqZgpHEC/8EYs9Gi1iV4Ln4QxeRMjerMmPIzE2XB2ObHvWw
JVVtO8tewg3WKWNe969hcUGULg4dCZfrF/Hy5YyZ//9T2gDVCJ22RXncylXC5iqx
1ovKeD3LlHGHdIwyIaQu1Spr4rm0x89IxZkU+kvfT0AB8ijnV3ZXRrEwwDIQ8Cpw
Wxuthpj8w4dKgSW/PnZQMYPqcazIriX3xHDaHqLseFLkV+j+lx7WPhIO3tYEboz/
zCK9UrtR0FKmn0QnF8d2qARrBJmhznh9qpPg4RZoi77S3HIeCAasdwF0Z0T2jspe
sIS33ifayfdZFNrw2CIc+JAzh2Qj5TeTIRtTuDXc0oL4C08osp5D0Hml8maUPvRt
39bmSfov7SQGOcoSzICJZ8ZZWypM42DQjBO/bLzX2BSCxovevjH8qzyHQLwV2s+L
ymaSl0t1uoVK4+4ltfurkJ56Cm4Rt69VSVFcMiuFJJ/mkS/Akxe4/z5kgVglecEP
V0gvby0XvKynKkx2eGsg1n0JpEQHWaL29P7vp4hCdO6uKjT8XJMSYsI/PmzetSwv
Iagzvs6W8Yjv5gLaIAD/a5TpNHOadwKWTLVJqXgWbcTDVKRfirVzjDawL3W9NR4X
O1Ri8LuplrwixNwrDMs2iLRmISnHRa1rWpGHhiT4EI1DGjIJbceem1bGpOpG1T6q
Sx9i7Yg6rj1TGnn0piKfNeP9DzwhSvEiy5UpQtVhPMjAdGN+Xq6X6ZMfRERXsGzj
dk9DkQIvWqiqGR0pIttR5LnOTL5JFOEqIqNUsPYdmk3KocLcAaWF0ejI6FDv/pLe
bWvBy50dxzpw+B7g28FiaCni1QqvAnoUYC9jE1p/4jDJyaYzsNCy1yAFcLq3wGd6
bdviXpL9ugWCbD87szbkFD+yMpowVBRgGA4GElTJ5sUQyajFIYYpFoUZSkAkkkUw
E298DIxZTGH/clpKX4atMZeXdv1Fk4uTKZjzkr/FMwje/MQYUNz9Qqjt5NO6bbf0
gLJ8xGEu9kO0Dl4DeXFtwCi5WzUifTGpxL7JgW8/q5EAyFw7egkrD1pOLVcZRUCu
Xro4PsrBN6K4v0yjX5Mlkj3hwNwYPoh3WLdyi2d6Z513rNF/WUBptkb8I1jiOmZU
3e76JEM4VW4qndcArMrsBRp9uebAV18Q44UogP/3YVzX0MA2gUvK1pj8KIXl/GdJ
pMrQpWssbZQLPNqtkoWt36EG5WK8v8rVzhrnKYOdqA0YTvbt5kP2F1tfdY/iK6xP
lOuJc79VcpgHEq17c6xC6S39nO/JuZ9f4pF+dQLAI86UjIftXIuGbYt6/MKD2+E/
toZbCdBCwbYUgOJO1NTZPQywmUoIk3GsFP87x13eZKbhcl0Sr7MVrhhyzfzALbVj
tWCTUhXgONSkX0SXwtVvoAURoRN9DLM05zN27Ub4KOFFLj25HeuU0YgRkuEJHHj7
Hg3EYR/lpeD0XmXf6yBEjyLinjneR66ohmxVEmSGftH0DWZkc+azvrfC6UyzwFqY
myzCtllfUf4fVpfkvFZxMc/vEOlvCNRoBW9HbdLtnmkY2EZV3jYo1n+LwHdgYKVN
/I8A8euVBor9iD/7GG12P7kXbRka0uJhuazfiFEdFVfYHIOsdQIgUxdsAC+dDHih
EuckakKe4LKPTZIReLlHTkyI6EBdZTQzDUL5QjZptobxsBJc212fe4lwHDaJPa9P
ESJyPDMjAYK6gW35TTaVF04mPYc9LqOp79Inium4zidSsfhSw1+dW6mHZBkgirbV
8aBcf3bXWO5vAVaIvtIvmjy3X42iZy9vRsYqfs6/Gs82X9e8muDchMDpY8ZeQmy2
gxSf3RXoZ/7IyykRLTaq8A4SKGYO9Ds82vXj57jilklLzJyk+tLorfCrptPqoWBY
QK/TWnPj2SOBxwZrkHbG57tIFNUyvxn/vlKAOnvctOf/o+3fuopzZs1tsSoSwLS7
jm1qmk+ptZj/glTrHAsQYkIHArFgIeB/TUeKbh/MvZvtwIEv39CN5kpOAsmtBd3D
r+6+nrhGzIJt3zwkZ+GZRG9mDba53+PBfYtd4IiWNoLqW6nuD305VvS9CR+o861u
4TArgdqxoVH95FbO73BdQw1xlfaXLp10AjzI4TedUNli4TyVPlfRTm0iFmvkunyG
GchHubzHgrcLxpEgOFSykmwnR+SntVdr3g/p0CeVAiOPgTtooebNTpNvjtviKhmo
zyH6p+LLwgPnwHzn+rgt7fYWt+KKFxEhxJDD0u1k9/NudAFQA/OPPjg4QLc06IFj
98z8AlTWiyBdi/n4iJBTajD4Q3W4r9C9s3l+8+MXlqw7uY+YG4zWO0q8sX6qPAKf
kuROFv+G3lUgusrs9M9FwwRXNeu23QMYM69tiOO49GDyEcI1q39arCBSBJJreoM7
yUpWGYn+V/Tr5YM5WtE9g+S369J/LeOZ0J/gFmG274vx5YcLJfxQ7aXeFQFrYmjW
l5Pie0Qfm8FoWXImqmQSb7Ka0ezsELZ+1LftGfsOKjkQCwGkV53xK4azZ5lfeLy9
wEvCblcbDEYGBXneg5XkuWMzJnWivu68PxIhZi8EfyhoGoCydLZi8Zwt/8TAJdU4
ReAgr1dN5lbCt2N/qmXg6l+16Vx6GcsVdg7iv6vXF3k395Jt17D//wlWgZsrLsnf
/lGip6RzJG2bf+JKXMwBc8mBZolvFClynXv1skif6G4BV5HxRzQ7HIKAxy2NNoi4
QKbZwE4rJ17lO3CjYgVJkJg0nY5nY62uqOSEw/3lGP/h18JtrXflnprm7RtcpSyz
w6Oic2Ge/XIIpDmmwe53xq/QQwNhvbU3jUVc3/wC4+gloHZjjZE1PMbKja+EO+u5
YLhgddxwrXh0be8qbszRzsn1RrnghJ5sR9ZGCO0GdwWH2dtQyRr5PBzZjv0mTUWf
7CFY8oMBcnKMqkKqQlVZ0uApxE/+9DI+DSJinM3Xxh4mLQRS/vv0YjgFBUGtHLtf
TtAgT1ynls+hbR0J4C7BrD4xV9PNYZNGasZLc4dTPOQ+sBQYQ2+WBY00jBXzVMUI
fwHd8ILGTtwSLNXoSJu1hq79Pm8OSePc8GGQU5cyNCC1X5nUHynDMo249FeeMw/T
qFu8GpzwdcQNYu6cmchjavxs7owzf27cGul9RkusekhATweF45+3g/nlaZZ3CVFA
v+ozTUENc185Zi2mCPpg8Ne+rnThRcvRS06cdD4FPil6ebwSl7KykYv3KnigZpiq
IusomRLym8R1yWQZiPaB9KMZLfovBxgLcOdiR7+m62zolh0xw4HUWVGAoXMEP6n7
YcnrCrQRWefWuy/ia/f5w4om4fNRElUXsHEssT8mD9rg+0eRqlQyFtTJm+okoOvj
YMtvsF79jLnHNf0qErV0XgSgce2HHSceYpWPDYhR+WlcwZwS0BqqImECbTJO7w87
OVYoYxM1xi22jWKG3StXkduOuWcv9WbvC7gPbw/LKRJs5OsjGNmkqENd2QT5QaUP
/4WFzq1I9UdXT+N5OGlrTyWC6hf0iP1GpWw73bbvPV0fM62P841SPmaqPgq/Rgpk
XZiFdNwYWQcPhbg2/BdXfNfCSl05k8K2DZon2v6IJ7kRuDXzprCtOA1lwZMEfzvb
Dg7tcAR1VI8e9tE7FZ6rXpCEJ3I7gCpJM5DN61iCinZZvdK4KW2NIKOh/QfTLJHQ
39koGZ87tYe8TizYtZzXWz+rfLtHVUI7cJLGifnhywTyP6K7/E0vK3Ks33CfnDNz
ASYM+wIPNSUFPnT48UkWXlWpfmnFvooMPY92qzH8GE/g+ubaDjtWV+N99x9vB0Bt
sDAIGednqDXPBTWyWkgrLySqfSgW7jmhQaEDpXINvFfxtPWoZiSQdfsWuPn6lyFx
a7d2TQj49nukexORvpUXbS9yPZQW8NeZ3ceqbLTK2QciNI6lMT33OhZB5E705j86
/p932XyzBAENrqqQUOp87K6kWlN/3ynmkxMY6DyWja40WL5tmTpvQYFnionSL/MW
c8hIAnpPPB0UhZLtb0VFfL7q0UhCsi2Gv8NfsbgFTl1DVOSBPtuBWgK5OOXkL8vm
4PDtJy/dDOmY07i/enyx3Yk6QqhVklz5JhTbAsEfnhKuWKVUVr+6B/lC7+fetuve
kIAHmAvGSL4XGuekrXXUJU0/W2aJhTg/BKl4zXbRlC6nBT9VVkGqPZZGgjpYiGNs
OTwCi8nbAb+rl43P3ABYmVfeTQ3KVlvtF9ZE5mawmDQsf+jnzxgFlB6GUibf7xKf
fuMz2Y7hjDmf5JLuz8Ryy7AwSH/rZmyPLsSu/WATDAlUu468imxrR8t1NVuY5l8U
Re+53HPeGn92hZG7k4yHh44Kp4M3uYTsMJmJcojDHHHUnd/zsRvopwnvcN7zuC/T
ZPRuwr99eS3ZlpxAEUglkWVR7QtFIBudh9urmhvf/r+6NJz01BPrl+iJXGmNS3c/
hBvKiQ4oN4VQdI5daHHML0fB0pjfunZ3cvBsmE5cO9b024lNPe3Vw703fpBW9odo
ibpHKHjL45JEcjXIQFdjetq6O0NustovG0vi3ehD3XOuIU0cmIKbIcmrZ3q5P4Oe
jaYvZMJR3H+oGwoa2uXTSB+ictz5UOA584i4/sfK67SdjVhKPDW2ZThZ+pkrT4zo
ip/lXqaemOOxuQY0ydZ9pRzenU0JOdapzejtyITw3l0xQRI3jr3NRQvw5kGUUhGp
VhFSp4h7vgtmpmxh2cQzygw97r0r5taTLgugCATX4MI+YPl4V27aY5Q7g0X+ZEIS
x5VPNqjtvmS0Gv5xaCMTWdbaCXK7iD38Jhwc2Kpq5ChV03efjPYqFsK31pgvIvHe
zFdQHP9eCDhfDCsdjjhR43PvKiN/AXVxS6ApPE0clxEMTQ6ySr48Tn9Glp/KEJK0
2NUGQhN9j6s8Sc96WnLIx5FB1H0tCEC9YDuEbutQdITRDBAUn6rMANH5WQuRTynU
GTBl/rnt4jthHsOfjHWmCG7ZVW6R6aQZzDffwSnFA6uwaTHnADgRC9jPRVBjDTjh
ynEWP4zYdT+PHWgO9MNVsO5NXMmlGA/wLuekXqDvEitNiXGcuONqg48qB4+gOALw
adFcOvyYnqNVNAn7IadWReTpWsavOhDs42AK8WaDiaDHqkNbLw4l10Tm4VyDlTs8
fiFVifk+wdyxGmvPHAT+u7KG4jauZh6C8JVcGxTYGcZx0SdKVYULMi+412Y5Jy+/
oQzdLmAnLj18C2QqTfPkISA5dmDcKwF/+HkTDv3E3UD6xMOKVoO4Ycm1WGIAzZr8
6DQqGKNAIs4OI7rq3Myc+ue37S9vJap/52sXYRC76Kbaauv2/P7rwmXOVUY3YnK+
AhBPqdyFIaNWTSi4sTMX020KQ0taMJB2P/ekcL7FtIXQTaA0c14jfLuEldQ5Kk6V
nPE68SCjeNUw0xV6bAZw6pQ8DZFTPWohqzGzfFPVbKvKwEBp1D7m32JE3n5EMQk/
fANNLUM4ehaSBg2X+KQoQUc1f2LPwxvcMg0DRVDSa1vJfLpUPF5oPcLuFj+hDU0r
TgnqEbh86L6d6A73xHozAoXAFbZpltAOjcNq9WlSqSxvssruzIHJH4u1ab+oJzGk
CWZg9pvwHQj1K/y5Qxcl7eYEy8/1bAvdwVKP2J7y1tD1DVXPIG8EuQfwrryfzXth
sMs4d/OaWpB6412S3jhfKciDy+y4xuMI/rCNxPc2wl55QtP7/JFvgEOZsMJUr0dU
h0OdozVgIMfdrnHc4SHmLdOrCOHZJjAuRkS7HnlgNyQlw83HlNzGBDj1FL7r1SRH
fjfK2UcxdFxaSHEWvNhrJyIR9cQ1QaJfZmNyu3GCDVw2ywYzB3Kx3Ya4Ab17xfHg
fXTRWZG1dy0Z1zxncPLv3r2+wwTxIn+Xj6fNYvgc3JoSBbaT6JvXlAgubcEjT+Pe
cxtZpo6vkQ6uxoLZkf6l1S8TgBrEULX47niA5Hl1KLozLFZ2zXeXrynpGKa+9/qv
n5wPVgcpVLnv4/ZZDblAM2HIla9AWdj94ELwUXZkGbL4xVlFQTtpKfg9UkoUVxzP
EO3ZjNlCxSn+l96ffwurJI2U5TuVA6mD3tF3S8SY0vLfUqcZ63u/kDpGPUN9sYkF
dLyPbtcWlHi+yCB4swhky+44+yRZe1LIMthXqiB8P+Wu9uPHlw6MoFrSTkKEjz3e
GzfdyssoVgH48oJJmKUlrme7dmHQvLLSAVM5/Oj6yjJY7KKtXa6D1MSNa3wTRdYt
63C6N+1nC9erwN7nUiN+WY1rOTm0Sz2agsEE7OgycXHDOeJciU+hsyF2UR0y4WmV
brYnGU5YofYWwJRLb4ohYfokQJaeF/1r28M4YtLYid9uZzvmdfm3FtjGtqwhp6Ux
RQwHIpoYlitw1Wumyj/bXChlxR/afIDuFpfR47PDd950+aieEfX7JEi54K7DyMZq
lKfA28fXtZtl1syCAWGSuANlv954fUFR+6OyVc61E/iYBI60rw2MDIBepumWM+RB
OCsATb73Qavt4COHq6AJzMF0OAJVZGpB8Ytv0gSqXL2koeO6MvQ6LI1LzKaR8k18
4lJiaS7W5RD0gG37nxcR5p+a/UJf6fzKJk5P3w9+GhfTN2TKTZzin8OyeGxmdr4a
0LyDCq+JFOKqd/VWukfIZr3aPdNnqzA4mBwUO7F1dt4FcaZmnvcpE5si07oWu51y
jDdzn20Yb7iGQAN8KQxXF9yiMuNdl28ACaYm9wO6xfGN7c7YQKinTggacYjk/gW4
n6aDqENBvVNrHVVu1gWWzb1cfHnYho1HzsnceSi+EGJBnr/2PudJR/IdsLt2dwqB
mgCPAebLMk3QDaoL2GblLxHCE+IBTAkktsb838B2QkrfJUwsESMunOF7RcWIUOgY
wBiT8NkZGXdKh76A7/Olc7rqtgN6C36WNg/Qo2C1LNsB98/MUUV/1o6PI1+BUh9P
BMAt+NoC+5y7VHRmvLXtd+9NvXEl4RdR04Zw3tKoUpckLLg+0RCTRaC5YCUGk6IT
3diVCkM++QbUW2fNJePnjp7cxzR+9X/cxcsomJeYfGj9bZsTA0AtmxZkOkib5mKP
9WFk/IBZMSTqsNovk5HssIH6TukDaXzh0oxjdWNytqP+oHgtpfsc4kHhDbJZ0uRe
BQGb3CfgwayVa+pkguO8QRh+jxYC9//QzqFoBO5orAePfCgxICRmNA4Q8mcpJLvW
29E9PJlLKXzjz3gxDyZhC/jyUEwdtXzACvXKiJDPihl8SjBRqIe5F7pSRMAsrQIc
QVaETqzmhHpAMmh+bsgak2n4tZVTbOL+GIZQCVIYswCmr5xABDPaSP8yIgG8MKFs
Q9qGSMjIucD57pAmYxcPWtDba7NDA2qHtA3MrXgN3nMviF0zAxdKteh9SsC/1XnJ
Mpobm3qXdQLhGSmeK6O2/KWM4icoxYFzXgt1BgzrXcXdNvEZnvBNIzFSNcobT76h
iV5lyn8Zyx4Bm3N67NoZuPmqALS9PpKILktv0fzjDPng/D6Rqy+dXK324jH2zVGD
WlkpnC9O0UE3DJlPZ3pZbmwtOOF6CyBOaKgJKqGxkgEOfGjHxuoy4bMInsPtCbVj
vzmM7fwpxLGKDppKWXtT6oT1Hp4AdHHltrP+nmif/OSADS1KYIyAgrLh2IdrI+BO
lpZebUnblQZrsm1BI86ZcUDE90pfHOrjW4W1ahFpWSEKoGUjft1y78KF5EgJ5K8M
ieBZElkRIUndoM6YePLrX3oTyF2XWBxgMo/cIltLodHehPu0P8Oqm8IZGa7SQ9gk
jmIGZPY21zeVmfUHxehjAI8m92nUyntcooAzlRAv1R53zNySPpBp6R4PFMAJlKMS
GE++bs3CfJ5kyBAB6inG4ixp9YUkksG4ZAaUFV0r8/QzSqyessZs7oXUvK/cFYFd
GKTKveEuS05G6ZNPLowFCKn3y9+N6ugmHDCLSrJ+u/KJuiz0Mmb/l6xariP0FFZx
yKdixhLFNAwkc1F9RII7FoCPXIqowLPYhHkbNquAVhb1z1RaAWRnGk1BvlcCgd6m
2SzKMPohEp6wvhFticgcDgl3xWeDiYqX0yoll3VfHoRoPmyb/2Hg91qhq71xyDWE
q5Sg6vPItJac4mHCMATEii+0wc2Z72zvpyruAwJfIgIZWcohz+Qxq8h0rSQrBnvr
NsOu3j5Xlrbn10KabnPIZCFN/i/g3Lz+Jpo8KsytnXpxi00J3P+THCMUtXPe/v7a
0dPkqmYU3ou4fvur37cLf8jZCbpGpvsKSAH6OSTA5QDpY7jPV9jcNA/9UzsF6n5O
EhouaLdL3HIw+iCiAnzq6ctZXl/ICglILEDsMNFPCVsROVCzMDmwKYfe6pB7Mevl
X2v99rMg2h6IIIwdNXnoJzPdCLY8YAre2QFmf30eNBn1KnCPP478FiOoC9AR8+JB
8Pr5ofc1omBXdKXEQL3Glwqit46EJVPIT0UoVz5lB0kZ8WXhF/Qc3fHRerU/mTQu
rX+j6jPjpxQclZ8xNNm0zdjnwUMaxbku4ALJF0q01xQSYSp65pBXLPijM27JrDWS
ZDVSOjnJg7nH4Yw/CryaovDMtdC/lGhSgGm2qTQKR4IsdPrNoiMBSlWkLg/CM4fe
7W3G4qHZOVxvhSUfXFuobazamF2rjR7zpNHgO1PXamUC4YjAqx2ugvnh44AualXF
NTb8KSaXZxOqxvbeSLLJAvSERJn7IJ905PoHBPmatdQV9FCyQCHHHWW6JcOT1+Wv
o2hTWi/693pEYj7/6VotkYjIgqKgc0KUjOfO92YMEKHJZF/YhWjRINB1BqiGbPDQ
Kj1F5Wo+3cKjfiEdOYsFjKbZ7eUpV4GLyQ0IToqQdYk7uzKx3FhP+YlKu+8wcvF8
qd00rUcePLgqfckI7cqzoepc7lcWOUYyOC6U5aNEmSJHDERrMmp7rf6p94o+rCHs
uCbPztAvNsvVIRZPC45WoRi6nA7PbZAI/klYzYfeHPbUV73BiNkfAooY+mcuGK7a
iKjsHgtRmRF23BRcH4raUIyWY4YJ8CgI9/cg6JisM5PxFe6Q5YMvZiKaed/5NAE+
3LfIZ2FrfmRsK1O3JlBrCPAPR807eIGuekww6z+vXjHOAeV8M7iuEIVf7sAUlnRD
moxeRhkUYsuieA2usy3zUGLR9xnep6aQFo9J10BlCcrGSAhoRuXMUznnjMCIFOZ2
ijnSBjk/fRT2nHr2TJnlqZaGcKzuYuOmh5KjBlq8EbYpsSuH9xAsU/IgJlrHH32v
I8EnOoKGybzWvA//eIiwkktVZr2IdyCVkRtYzJT82CF7Sb0qJGb18oCNoyp6euxE
Cz+l3db+nSZqQgS9B4DQQkXag4uUK/aLDK9MNkUCfQjARRLZFV5U6dFcakIA/HJ/
Yw09ynBBUZud7eBK0RMVNeuDVwnaOby3pkX1io2hXnI16KIsag+v6QPO+xm9ZbsU
JmPP5RTmCfG8NdR0Da3EXG4bmpAvbmUm95Z8/81kglt2bAk3RuQcC0SSzzehuOJz
Mkr5JnKdNgJdEuoEpoDMiJ+ABYInBd0lR9xqM2zc6r/gutslkKRxRog4ufmDRvZP
VUwtcyXqWoJQ4ar5cGiE3ZDveip5+ydM0qpGrRh+yCaN6rOiJKIwfjFyG5hNKXzL
GGZZUJdB0VglxoDPqmixYmnVpGWvIr/2fTX68Xd3C72TTUflKPMd+D0EQrZXr1j1
Rg3oF7PSuwUQKx+vtdSnaFi1cfC/nxrBP5sG7m2leTZgQO5zI23sLDf52doAPPnI
r+yHJME0quM4DQOALTOURP7OcmIItAfhQKt2D8fu0Dsg/6G7lK827oz8eGASwluL
IiINfqJNB3qk3F7xDP60Js2HfRaaI9o09PwBfggytuyUrYSPIMi00oRYKGGa/RI+
x6EnCBKbAsjMxYC5K1lmLyKWzuLPIs9pzLqNYh6Qzs6vIbyqegPvhOHjIFyEngh8
GBZYePLxwxfMBlC6dmalvx9SQN3acJJYMvF10cQlzuRqNZfZwiTq41toPGCOxx/P
XxT45F251PQYpMBuQvcoAByF672B6JTeXUaYUtREVRSf/lrWOKSzxvh582rQO8bN
ZgxcgCBeV9a9M+UOoFLjAylQIGHH2TJMvE+vnhrwUtVy1cGzmpWuQlhEnRjn1+83
i/KViyM7aXhxleTC3b1LinN7ppC6QsPUQhkLDj6+F3lSvWL5bFi483op/6cscw9i
H1kJzj5BhhPY2MscsJ9nnoUnQZA/F7XVpUGznfC1n5hdi6TPPkseC8ZCUCF2P/M6
UvNVvx0GlL3h48j1wbHUYc0TOhMojLUuhY5zhJQAtIOwlmGKW10qkMbrA4SsFMNA
Rl41QHSM7k6Sxv8QEym0hmDU60k4qzjwldM85vUdDJ7D+6c9xLgcEh68CyQKWHlG
iLSv82ywhJ9whupxSR5PUb4nNV4W8D3NT5WFk4H8zP/1TcvX0kCmGMlgjAZvYCk0
U29esxU6X0slc1ypw3FA9p30DlUlC2BpBqHjx4SSGr2i7rjtmD+NxTLkpVBcYs5a
UAHTDQvtEkanauf+bQUbzCKVWyETUGqauhqLEP9RM123ZpBnbf8IyqqA1Pet3zhH
eGz5YPHCVAbPCx/CoEws84xq8PwkBjabeEgHsyxB4LX8HIoMEGKitCgYwg8Fp+BP
H0sLAeMnfrXK9+EZdkYc7rNVuwJSSoo7ROerc2LxreEbAfG9dfJ45IBi602exwek
sNaQs9e/FpYmmCI7K0z0+eI+Vk3/N4pH+XBjN8PWuzK3heHDdZMlVsNb9Tr1T/7C
0BxJsfON+hGisRH79CxXRkA1rj90Epl8leLK4JFtQVPnnlCKWoRJitS/cV4oYuQz
PvtcUuEUAIrNF8Jrg96FPhOMp9JGRSnenHkhHl5L4JzWXkFc4xxTQ5au5pMPtg3x
Eu6wLNVzC3Vdyi2g57Z7Pv9yiBw0VeJ0fS4OwpsdbUS9WG/qzfoLe7rbpeIl//Dv
fTR615XtVoq37e2SqsuNZA3qWLMqjQJYRKRngDwHagi45YwS/NlprVuJVwMolWRp
mu8xg/E59oNaDytJjaClwK++CsMhG8cETeP+6MND5cRMQphQC9c+kaUVcpmkt3TO
AfslE3So5in58TATfrtGC4iVIAKSpSyGZ7/sIZXPOnL62SFaoXsbZp4fE57jbFiZ
mMMCEjGIFo4igoHtLpAuPpM7ccAfV70WOmlClyNs7TJ/93qCTr+N2yjnjPrGmb0q
M0ZFOA3PzenVdQYQXDhgWzAKvT0giKjoH0N4zJxIcYYtCCcYGZXo6/alcH0dhTLv
3/if6WsXBA2ttpJO2gobvEboXA8+nK/hEGgBFajybwgcVbsIxNal1SX6YSdSLs9/
9LxDXXcpzHzdobU85SGn1+SAHH14d/QHEEsW1jUacLILG9TyQrugxoAByA5XIg37
30lkK9wuMbKNoFUNQmFGWdsLktAy9NV54GTdsiQyJifylGnyKsySl/yc5uTkgKX8
EELT0SSmV9H5JhdEwdLVWtUMZmCGja0Jez1N0CMGCbWczqNPjOn9aGZezurDR3Cx
f5cL7B/zqHxHKUnshP2JibjuHj7NZ0vGIo0roAc50ngdvSzmjJ9AfLXhdyCuGnkn
bllZft8rRiyudBGMy2rSV+aruayPx9Sx70bNf1L+Gx+n2fEv6e+vg8/23BScwncy
4cEBqGOvPAlRsCftXpf38UjeCrPatviC0HJCpl2nx5yggBDMtuF6sSmg9JIMwHBz
gl4vtbfyLPwg4S+H7XnLf7GwE3zKI1mMmc+U4cxJfNNX8DSK0Bt9N6/Yp1aklLbS
Lj4+XRaAFb8Tj+r4+oYoh99695kk/kO6SjTS1bqSF09xc+Ys4CwsY1buYhfu+sYP
Bx5/WBHvOPBS/xl0896o4eGqypiKT49a/NsYz35UkuiGiicBYvo5IClhYW3OZsvq
SyhG8cqXWTqpcB7Bk4AGFNc82TNMO3rOP5GI5Rn6PvMrRXshJPSCTSdy7Cf6bVz2
j/D4bZxeBhGo4jx18B9q3BTWPpOgfEIQ7iFdgjzcZ+LUN1W0aAbQHj4z4piBa20o
281Ah/z14yWYWWsPD4WEGV0x9GBn0BHiPQS7cNd9S951oemRf9PsuLzXqENp2kQR
1XxxpcvEcx12+ormxWLaGXjHuWJCxFTUlw7gKmhTWYrLProWoyo+5FjfmLLRxVdp
2vUkwNXEc7ttfjw7Gx9BkZLGOO+/Tc2ms48lORQ131cIyir1ZJNbVdtPuuHR0bH0
uaLpNFwcGEOZdr8hqpEz6M0a+AvLGBGbm6rsc65N5SKhOIllVU20zBrCV6W7g1fx
n4+WAhV4Kl/g/Btdaw3vQRlOYsoxe8yEaBpk4U7HkEIPnlZxve4OS6m1d/lOPoaG
huNL0JnxiIn2JUgYKj8SiLxUKBHiKt29uEj0+JijVi7wrSajRFFCNU/sBn/d3gTR
OiTZwMtjSMsCkSQ6mayjCdIIMhNIhUM3RrD+nisXzFlrMJhAEqmOLsnx8Lanhp1U
0tDcrkjuVi0MQMZ5gbPHeA4T+KaYyD99Y+3OyROS4IoqMddPmy8RUChkLlbYXdJt
B4LJoiGn87H4AA4l+Qc2nlfyM/+FGy41cKdkM1Kg2Eh6eoMYpakAqGuBYT6IPiZ2
wXi6wXnah/6yXFogpOdsYP1TJzPPaoUWpA82Vv8yj9Njs0jq3k1Mfof7kGhRJuTk
UHc6g/iJdavh2QGXBiNeJGSTZCJSBVRJcNEtJ/P9P3LdHjN1qAs/4F605udG7Whh
K21r8QdxdX+pWhDLc1slxjDkJrD+sx5Jo65v3u+12BPIycKov54hQ7Tb0+HmEo/w
GHDuJk3dep7QelhjAqeQpLuWnLX3FvJ0rmOFUnQ3wldaBdfyCw6k1OmO/9UOlW44
YPKZA9cVTf2t6MZNHmCRE5acws6yWwkksBDI9R4btWX0kbKY054U1TuY7yvYn6hm
gnzJ4K+mt5wUKqXBBKo1Aukeo7pkR8hdP608GeAyBhVDclWxvR9PRoRhBP5DDk4v
lnTqlqV9dzihNGU/+aIueXdryX6WZJDE/h37JmjLtZP6Om5oP3uuXAcngMYkdfZN
zzwoKHUk29sD2+p4c69qwsyZAkfhAcnxouvhgMZ6kc1Oyv3pGuyx3XuxQVNKbwUh
nO2GY6TyodiFfHhvO7EonH5GYACTkaUCyPXryBPnVS5OZtf/6QUiqxq7PKyAhlzI
XO+mSEtE3MnOD+Wj4TCwf/gI8WQF1GGCVk9FSd7TLYEyLT9/jQ9FxSys/Ptdew4p
kIqmAYAUs4vrSZxFzkgssxBJ5qUXRl8aDpPMilmLEAYbF5fld0HWn2QaLFgdf+VV
/tBPiCXQCc8Ymko/HjeQd1Ac8cmkF6OeMrFWXvaIuNh4ojYGdjV1INNw2hhovoRU
1bJnJUHzurS6bGEXLJMlSGTRNcwmyN45vSe1We7faaYM3HfpOHaJjrB1PHVtdfH/
M48Or6mlwKNEgzZTzyPvjLIjrEB135PMSwzAFb9rSig+kkaWCXQZbHemgvFatFW+
uYSrPBRcMAS/Xkz9ZaUYvru+bmHJhilz7WB7D5hutt67cs+qz4HEoh8JCBQBTFTl
gg/U+kUpROENV0p1E6PLTOf41HbuZWzyKxM3wnna2dK9FzOZGZ60SO+xPSZBAl+C
MNQtzX5Ss1TxKm3t8b6XL/9CtcMNW2n4m28IEZ9R7+8egLFRNkQEhWvM5MB7qpz/
x0A2O7TAeO6Y9i8avvCfDFRP1lr4/DW8b02mz/2G+03Rel2XgZdYaMEDgFTr5er2
SAl3swxabFhm7OkXj4v5gNLmu7djwC492tfqdI2N9hB6v3S5uzZV9vgaSJFuRgzi
4tzWdP1R2169MhYj23gF8ld17bSqdhiNsl8yqaM/eZQECBlyux/yI3lBcGtWez/8
aWX52dKyuFZg1pp0GdZGf86EVe5mftZlotgF7uLkuVkk/j3fzFfHlREsjsebNShj
wPuOANYltuqi6CP0RuAV2V5q8Bb9r6U4vqywd9rbyUPWG0/Dy97oagEmRoIqxSN4
3bVlO1mSP462p+tXrYWWobh+IWPjoczU2T1TVu97uxARbv6Bz9Wsa920Ny+dzIN/
CM36SFMtvxaORgqh5MYt3av/IdS9xkMqmkJHVoCQ2KHGgY2gt8oL5r3TNuu8b4E8
zO7pC7OXASQp8zTINX2FvQ3lPdXvJYvG6Bzyqyj+SiBpzcEXfTPAgGGKOkzmQ2CB
NogKw1/tQKqmmCbqDM0LKgLXhMSOVyDGitayCF1NKYLsg24UhBH1K89TOSLZXvqn
dBt6H3UL0yF/HVqR3ldZSCBOCFCPEXB1VxBeBUV24IgIM+XApL9H4OLMYJBxb1BF
4wz2YfbQqLFAZGiflV6+bi9Gh03OA0DunZGS0vEtAp2pn0z1HA58AWTXWqhraiT2
F9MADXPOxvuEnkoX6NnFkRwSmrVCveuFCQ5dsWj0ouUcyR3Cf0oWIj//NcBGMldd
FSdPOkZu82d7qfwBw4pLV3P9Z3wJSUDx5vXPYTy9cMTNu0XQuu+XZ09r8xysPBQj
YnT4o9zN/ltGtG/a6Ny20ofDTUuEglsKrIQucvrQfZhYoNsfKdA4zjn8hiJJUqhi
JdcXe/kVyr76URliPJAImsWJscfRrEIzknTKXPkVb5lWMaXMt1+WV9/s4gAjnKh9
z/qiUuo58drro+5nv5o43al2Zur7ptd4/ZpLhQHh9i6EWp8Ek8h8XIG+70g4avLv
M0K4zq0qSvuRX9LbOgy9QLzewhfYJWp+uehvEZ9effi5q2QLfCX9GdFwGtSWXBrY
I0Xh2nrycloOpXDXCLSU9jPjuxrV5jenSoHRVS7xN9sqAiIvxGLxZ70dWP4fJcTc
InwMZAd8jVKgEYprQubGVie7PuPSGRbHPKVw4dqEZWY4Fi3uCq2mKAa68Tf5b8el
k8F7val7mUBtJS+Mu6TXfqrlb2+Kn09rk9ME/uwcsRm3yAlrvlOz0uxe0Q726/RR
ZHF8ZH8/wguh+mfRQ2Ygovk5VovOQOvN03+YaX+dUW1ilbZSr0ZPJ/BaEdxFzype
40ZOudAONnG1J6bMCpVCR+6JD8ze8FPfTqTOoFbKfTT6mZMC43UJaAq48QbHZ/YZ
RaSrkQMC8fWUF/qP3eZ/UR/niqCpguQW3AJbicK3p7QuKw4tgIai+OGoaXLlkuC2
r/SoYwiAhbe2J9zoNstUogHflA7WjTdOmA9buxA4ZXigBg329hTwMMUE99zCTJ52
9fSWAKj24gMd/PqRb7Bb7ENXZU/pE0x1nuPSMnfr4EP+oOnpET4YOTgVoOQmmj1n
TRmNaMhUJaicMy2gCD8F89oeMG6TlEajyznvGfp53WjEqWmQyezyTQJLQ3NdXQjv
OyQrs0/fX+3q/XtXfkuaEbLn4ZH+S0nVEbA5wQ8OjguFDB04rD7WkT2illgHV3Ji
VTjPwKpqvjQdmHRiEFKEEcg0R/vpnZPKUw2pc3H2mkcJ/xEZbAzcCc0w981WW6p7
UcWpyXu89pCQRSmQhw0+vNVDSSihhyUWF+nXTRVaZyVFiLds7F3wWtp5xOhdTNcJ
ki7EfhO9Yj4IRoglp8LacHJjQcLGCKQUdMu+qMH29uy+5tVOkqpryQPZjlDnUoyJ
tG4QafSouWFSpK1BcTi7X7ETzFQxa7fPVglj+FBhysNp7kUS8XNEmmS7/oBqviho
FuqFMVSKsYXOob4msf2plSVyVW/PADSj6N3FANPnN23Yo9pi/TuW/Pyml+5rBtG2
fypmPz1JjiBzx5NwL4q5rGFyqnMrVPjBlqPUON7r554VG7LMHLfd3RcDqzQ7uMPj
oBZQuf4OXSV6VJ7UIv7OnH+VciiQ0Zw91n8xKZLA5frhf0Tz+0lPmzYaqHscdZvD
PxhpqCXcoziYCba/anAuxt+Am/vosJeDFgupvrUROjIWTnbvpOrfqcq8I7iwzUEM
43YG20EfNkuTm30/CchhKSYUI+9d7oSX7NaPpt52uIy8agSOG8bninj7LSbNOAi6
XKbJE3lve/HZB5jtOaj9Am303t+tifqheZdkTeXpNGIUu0dfPCJgPQIS6p1raMDO
di6aRbtBIpJqv94pERbLzEWBOWOX4cSwK19DM1aSWyuwbwgRgjBSWEg1vlPxZqPU
AzXiNrmNP2MeDHtzNZtHxfcaX1kHDmrDpT5rLz+LylQZ7IO/RnF4l7aD3LOkw0Um
//KY0ebWUIu2SffoVHM3KDYzJh2G2uBJz9aTZDkAXuRZbCWnGokUd4AnU5wLn7rH
coMW9m3+004plbRUPfs32nRyy9zzYd7NCqtp9c646aWw9ZY+uU1ZuI4wQCl9afde
/w1MKU1Psy+1M96fGKS67W9jVbEblPc0TEcWAdTPz/5Jd+btePtUcnD2Uh1bZzUc
8okCSGvBQEgDfmBQcj7u+Azd1y09RMeTOzDkwcqhraq8SwNR8ReuTUZBrjeerv2T
eGT+LYjPZ0eK2B+BNnoWaEnqRGo4WDLlnznDl60AgVRodbW3CPYqROHE1TZWQLRe
kuz39FvMzaGIOPD6iiBIdBsOD78Oj9LrfpYIgvFkReJKvNFg+ORje7yAFh6Zzgv0
leh/5gsWrfPQbSX59hxnTKMUHKQSCeR5xGrHwt0sfqnm6UI6h3TgmV0EijTCHkCj
YHMzxbwude6ZlPeEBmAZu0WJ+zZROR2a+eUVr2F7gdNDd3Mv8j2udmrHCbU7vVDq
JMBA+TxxoE+hgOuxqR6Hi+L+rOLjD2ptzbRhxfn9cd3XjjgwGXUzUoZPN3QhwYfG
yF0DIICXzkzQ861HOvHVaeDY7dfpp09j02p3uH2h0VluJ+6DdOAiD3PUV+Eudsp+
dIspTeQjh1RSvafqkR+iERpxesJcDFfVoOsnvr4fh8GJfJLIqJPak1iOL5jhQI17
5CiEzHzlV9DdCX8OEdmIFc8cJbyB/HC6/IcC0/thjZx4uQmo0Pb1OSNcRgcifddX
TtkR+cM0UpnqYydwXaw72DpgGV3O4dXHgkAqVMA6S6EgMZHiiJ4uSohGSb0vhhoW
bm9SWX/j/zmkUS1KRQikBJv+I/7ZCfXKEcQMtDnAPVLHim3EEX65bsgnT4sSNrVC
Q8LAVNfKc5dolXoaHRedyUmiv7U9OrSbyjNFg1rmL7Ucg0BQMUXV7owBC7/bkdS+
yQfWWTDXDIl7AU+0KUndTVX2+56AQiGwQsz6VqNeCP8pUnbRe4vABz0CRBm0E459
gc/TM2IQeftmlvh4niA282aubNbsaYPwVurQcyqiZ3yNI9kKmF7kHh1o3bLyn7It
izLgl306QvA0zH0f1svyb8YYdG0MXjSPzGgz5gkE2V/B2f+2fCPKJIFbA3m/vqwG
ksYqWr7DVibEsFausUtp0A9v6V3XMa6Co/Z3AgNAyvhOXWW9cf4KnbQeMtLdV/BB
HI7Y8dMFS6NAaILyiOrhkp5s+lp4qI1+Cd9IH+EpHPcL4kN/J7ixgsjGnS2J56XI
MrczZ1a7e5LyGSVZdava18nDsB+XCIXZRmQk8eO28INLxZuj9RNo0WMK+eUSyYiT
NSt5G4jd6D3MZjvCj2Q45bRSWUxfkmS3TKjBQtMp5dZXvIVYyLno1bBagK+RyGFC
WQ/U2HmmpX4UMSu5Q99Z2f7XmfSknhKFTLCOsNk6QDYOSt1hGhQaXEG5lJk2sgX+
PtA6dwYn7TmQeUVe7JRnCOVKRi5h/argNJ/1jjJeuaf5Feglt+fy1yyl4upHLJSn
mCEvntrobxM9e1NIccifcuP2wsxLRnl6mtTrbUbUmiXp9tDW8RHN/8CPd6c6sjLn
k2MC97E7BAQKuRBaB+8R9WWkzgWBQtWKimrA+txeWqY+Oaxazlz+2Oup3HlwzxQk
SoEiFJB7Ecb5lr6AN+pGpzFNNBFGd+YBO/en8weNBCREV9/2sh2KePQ8wswcSihe
E0fcIYekFs6aH1KDMUagO0pBnkpvMPak2EJqrK+fl33FCH7Do4XdxjUm1fYlA+LF
11PHMWFeglINhYpaL9FNOtNiNGjGHQgz1ne/qhqzNopC1v1T+5pzQiymZYrGzOgQ
+gSzOla7KO0gtoZn54VpbjUAmF+E5Y8pNd5ULLuuo7GI1rNqgWpu4YzCcjrnlibj
I9cVmnPkZ+H+QgZJnYzujr7NWBUn72RPOpZQR4VrhfbKAHMeV0ysxjUu+PJIdsDu
TQ+ezseIDTdHkjAdNNsYtGNU0EwVdiOcLzqp7Ib+2bLs2hZeVW2zunN/aRO7fntp
5GpHNgBOdsbfvokKj3vGTcnPwYPjC6paefih5+hW3vYbmijC9UES5cbGGQzNP23y
TppaSum903QDWfeZXl2I+ATvVnJntsB+lit92b/08Cz+Qr6wzJ6DpaiGBv+mJAke
DYcyM1JEnSFDBU5cVCJU2FqPtdBOoEgSXeYRfUU4Txazj+tSPB2c/8i2sQv7PvUr
vLKdDbtL83SJgnnp37Ia+87FtoOigDWnTXyidna9Ql6m6NfARYaV8gp/QSR1W87Y
xYvDi/IWx2jMD0uhwXfGZIf0rZA2GQrs3DQO+cd60tN1HV/ktfScXrhmTr/vIuM0
mFzsHbx1AQDhVb8WtVorlCNSMAb7136pEhPVUHhCBGEWkVEjlKBvxitDWaycyNKe
7sYf6VcKNP2feTadDVeoxLX+AHTVmom7YoutJf5IisdwL19Xz9uXD2bxgArWnlUC
Mbhj3B9ilyVEmUrwdrw9OqwAnWLAUYJy9GE2xix1UvMLFBoGJMV1DMFwbkD9kxN5
0fC3vNT2Pn97u2cPTXXw88x+0XK7QfTQwfIwALClCqafz0J3F8/WuxLGWaHBlxII
MzOYLyZ36ux0jlSB6U3VR0o6vkx04FceoAVjoksL1x5x7tk2FB3Rm6MOtrb3BkQj
4cuu5xrd2VDyyLM7F+D8l/Hr+gDcoY7K4k6FYISbwVzHk8JfkU39i8MH3kfVJNal
FvHAe1rXxqRJ+nfzyvByQdjBLmmx7u7c9iufqWtrE/TjykBTg4MN3NlrgU0jwW4T
8lPKqbgUbgccFCOCizhFo92+RpAGykzrKN332RiQcogXD79Jo/UNghh4ymVDomq+
LeQnJBrK25O/umqtrK+pz19nOnUXXC0ZlULOeSinn+w2xwGQapQ6YgESNzQQ3CDF
6CXhfR8pYxfsMauHjyXPtRt3bUJt1iHLfi9t9mBSy8vmiDZy0fJcqJ2G6mLjhDCT
cNluB0qydx2OKMu2fwXmNDroQgttM1wOxMYTJZg3JgWaghQtrsuRyVlJr6djDVOv
RUGuer2ExhLcxODmBV7GoQRYM6+Qrq63KcOgZK81yz7+kts5xySChafhHP3ns5a1
qp7ICFSxVBcPxsintB+iFE6hFdQemA69hQPER+NRE0jF4N4rML7TydWTCLU9qmNP
FQufSH3p0yIG0upKz3x4F6yep+v2xmeBNvfEQWwcbNjIDZSNd31W8kx4KT10O09N
YT4mh+XUsQBMRxPASq4eZMyT7FT0xiweKLqK+SHz4YvCt/F6in84j2kBDuQr60aa
3h0c8LjBIKDctWvlIMwytWec1lUaIZ8KxIFbG6jajTbWyyA19h30kx0ls1W/cc+I
vMIInqH7mx+Nn4gIIUSMDjk9OnPimap3olUk2Do5iEbkZ7hSBb1DIfs1s+W0LHUU
0bkHENwV8OCGzIBRLQyqX4hINLUUxVaSE7skHD6v/izTQklk5hqfHGUWZVURLmnZ
M0ai3ENxBPJNWIPEieiYOABV0dgugC2f0DTIYR3pK72wZH4ASYXOUuTdSy1wHzg0
hmniS8th0050RiXekX1QRllL5oq/ydsO233XoYxlDBzDnuVQc3RWbw5crSHkvVMQ
NasiKXYtmF2Uslqry0cp1K83ivgQS4PIofMe/WrQW30w+7DhH4K1IJzK76vrTVT7
iOxxoRX8E3Uff5ngoJNpJBWV2KR1A1Q+alZ2mAaE/L3aqgUoMVT/dukVI3NMEnQ/
AVkFzuHywLfDUnFao4W5Y7OykDHbgrXz3iehuG6WxSVx/d00yWp9VjrNMRi5Muxc
dU/iLf7hph4HijZB/hVevp0Ezg7IM6K9Ok8cs7ner+yzxW46RNXS+b6b0xtVqxvp
P36cCVNg4Unm92cODECseI17sZ8jwo7FVbuT49OHeaaiWdQbgrsXCr93L7yN0IX4
acd11quzbsaM7IXIvHDO2uOlCS1qIHK3AEjCFlqrPmZTfT7hkJEn1YKZm24coVZw
Y+rhwIewTVueMgjj68shzzoZS5qiy7XZwE5/hZxiE7fn+FmcE4TN4MjCAGxKeL92
wlcOuSUJHPrqjb5SOPxEIS+U1NJHlXf3UYwlRISvDR0zCxYEmNds7XEYFJ1EWKQh
EWqOGMjHQDY1YmSnaUGj/bp10UAV7pSVck8f5Lmn7bmsRQhztXdjlIQPh5XaMoJB
bYTnOaKnIw700dOeFNtSrSn/oY1kbPCyAZLFeBh041gF9jJshfJeKVReSub1+97S
TwhiJ1lnT8yw00k+Gyet5CfxNA9zyK9JU7ndyjabg2DqJ1+9UqyAbsuN25zkC8U1
0eEqGcF3wPTM7Si2YiKICgQ1GLHdullZ9j9HuxT1Gk+hBDG+h5neLbKxSV1FTBRo
kdmookzUzr1S8Nk1kHoTYRFCvGQHt6hNa7SJepjE3Y9lWMelcphO9Km7jBn8OFvY
qmaNl9Wr6fohXxRMP4n+nGNs3ax2RYC8SseFHEESXc0Bh6lsxb5glRDDhCzZTHE3
0GiBf6oe1pYbA8oJilHWFkwy8vk8Ln1F14s7yoalLEsOK9tNTzxvMjr/6zCXwz7z
4APngfPqLXGjX0KoJElTwbmnCTpThSFgcrvNvuQrus1nvKVRFsIb/KYU8BNKaBds
sglOnysyMRsea57fnSFB7TK536IhlglkhQR1sRGEHTEKmOQuU4KaOKyENbdJkYHx
JQtwNBHqD8MgihgPyNBW7xwjWPdixoYINs7qhQn4W8JmzfSa+dY6acINgFSE3e1J
79+dFL0w0Jrzf5RUgek1ZNYlcWz/MaLiShmBxqQyXMdomlKEyNcf4ncoKQTeihP9
8ODOmuA6CbrcxPJwSPEHJNgM7ltm0Wm0kS0v/E7b7S6mBeVO+1EuhuwlU3OlJd3k
Ka99TSNJYqTkz1QV8vPxNXZoB2TMDVnPCKLtWmfym9HeCzQFDE2rIsHiErkkVj8N
Ilcw5QYwP0tncdoB+D73tdTFPBj3kV1xcRBMMaPgGxJ+Sn71i3SEFRXRTsMkS9OE
4fpq50yhkUYmvFwqhY7CcUTR0nYHpvfvauBifxrrJ/iXlz/PwbpN6ecgBHmv/kxI
HrsGMy22okp322p5IAS5YjZP1kLF9VVCULbhsMGpKOMk6DnHXI3JnDFnq5EaDpi4
sCtBKzhT/+RulAHdjP1QbQYi/4UWzeUwQRDcTgNGePqB1mMmsvDUlq1YQIhayP6u
aM2OG9+OBZfHw/VnvHb2aBqdanbou7Gu9e713lyGHMw1PsZNKqta3NO7CLYY9zf+
63dMg7N0cdMX0DMAQ6EUZxnaxIGYvq2f3/tbH/Xxi2Ib3XBz694FYCykmy25Wjwz
pRtFHthswGwXAqOMA0LUObVy91m8AUQdJuOVMVJFFOJ9XwJC7FM/R21okG9hXV1o
jjU8vGwBHrFnETL9yDfxmSfggF13FwUfjWC1ioMfvikWKn7bNyayGdLla9RYfm0P
Qoyev0KH0H6VTmPqvyM25j7okVu7TU9b92Zs87so3F2zlqXNqOXkA2BrviSWmjjH
j6HmuiJSrz8i40qkP2oaUDKpXM0E6xUOyis/pe244V6FJi4LCp9lYU8WXLxJ5o/i
dcNOuBVYIVwArv021zOsrASMgW4+PNptLTeogjsomdRNaCFLhlgu+pHGxDTtWsk8
IGZSN3cgOUnzhxwGSDYodka8nC/9ys5xpmD5o3C43dEDtoHp3JJ/i7EnoT76ukHm
qlbodCyT7uKp86r9lshElhCqARBd1tvG41+12a01TEyWh7xHtGCWU2uSod83dAot
O9pIuUwGqd2slA52xyXqHVudRc46ibKiw4WXi5lpQGDW/wDsN4KESRHyqxeF8kJ+
cka8rgMap7GwvCOS/A7kjjCJuf5cesy4DdSz1eeQ2hN32qfpydA0UL/Fk4sz37NA
SY5N49Ek1frsDdwCuE+RE4r37GKlCTPmsntYxWFVxEQvPaDpc69mZLbjHC8PO0cv
+DJ4UuVni7NDEL76Wldllecd4p3lT1YUZcTX2gFzVXgwpRZ06tM25zeVF0PlnA8X
TJyrAHfiD3oCE0mDq/rJm5CvE2R6wqur6L6JrlmXErNOFx8xRr0Jn6tJfTbR4+2+
z8yUoGuyl8ArsT4nD++0sYdw+TCL/lxlcRll5RSjt8e4TH3o1CY2+sslx/DeVTAe
tG4C3SLp2QlsuYbLWF0Fej0nO3ZT9qJedkh8TGO5CobOsiN0muiYYtUv/PnAhnmc
ZASCsyd3ONjrFpwnv9HU/XbJHDV/Fd/89guilYfuODeKGcsM79VgXFmVNEYMr3wg
gh4g0U89pensn+BsjZEahXFTOInAuYg+FVvIm7TngcvAA28qRcoZx8fZdB9+dMFy
SXMpzs0PI6mBEajeF9P5asAl3a6mRKW3VPEq7UzpJ+14OGN/Pl+slvFBxOpGzDYe
N0vfEr/jxCGdZHKPAK0rgl+Zbrf71gxImpTNnHk8FRezuqTg32lg3vRsdp+7S3dM
j80sE7onQ+yWry+/jIEtz1cKJBpJuTB6O6O9ENFaj9xqZljpBpjEXSKwyMFOzl7r
vmPClpbHmao1kulJZL0pZmS47gOzNRRKxGHU2gu/AY7g9mz8zV7r/MiI1kVsaI2q
ScFo9qyJH9Rl5qyp5B/sO6ngPQ8ltjwhJ0ptV6eUJginCTHkhhvkXdMhoujaU05A
OPpZWK5geeLGMlKHn15AyYRxNnpYREjJrUoVrfLTHWIhHXGuiyQP6aJuxS7hnJPP
+yFqwX4yQhgfXnfhTA6DMURdWcNu9tSvXkP/8cn1Z8BZwPSqad3wF/x3V96SzNo7
lZ9dFCBOIOjUggejRoa/4RTx/JAwVGpByZGmGdx8DPUo8WPWvGYK2nLGc7egjIsS
nsjawXvfTZSPeQ4aAtqbc75PRr1XuoI9yfMFKju3mEsW01fldTl/frN0YfJd7uCP
hDZZld93ITcdoI+q994IwDhBud4kG9NXTeShTDNb6DeS3xkq3nKjC+UG5m++7zuh
gvReErR/dECVEXbJzPO2N4p7/AFaEux0Pl1xoGF42Nm/XqbhuR96FgTw5qJhvVnT
35q6gR+MGMNQS0L5aLMMJ6Kwn9eqlRNYvKjdzqmVLpbatplEvtUIMkbzmrLvhrVu
LgUAY61fJmcCcksQUUzA3RY0lC58OjnwIuE8M6fZDt9FAkCDtzfpS05swyfuTDGq
PJBCo/0/qgEn5NB80mCEcSYKn6wSr+CdkX8DavRL8MVY3VVOlgWJulE156k7dM4P
HI7vvxXCcySeIVisi1IO7tYkIPTaUD0irjYRtTL9xhN3XTXAQkGXb2l6fo6k+bd2
u1ryo8bR+GIBmkOFpDcP7hPMWS0j9//r+ytDtOf48kuAUDQM/rxCmreSTsA4Bfdx
E6y0qj1m/T9xrl7Sl/Jw+2+hf21CEl0ywTwE/GZuT4TLWNpFySI4KKZumQ9NblCc
afAEtWsiIz9H+/A7ZZwKf6zWXQsf0K6zpoCS9CLh2Kh4apezwn3a3h4aDLi3ox98
uokmSVqAkeR5V92vxtTlkYPodhBAWE1eT/q9DDkIEYBJpVtYIe54C6w8iVPXjOWX
JymXJIw8ozs7p/YJiWhjVTQKffaRfJixbI0oE8aLBJgJZYPP2IzSraPyQGGyzw/T
U7m/uz+LNfQWL3q13AN2aYRIxLOohS2iAPdCm/13avcFgthzobn1ELians8XlOuB
Xqt9SwUgKt61L94DtE6X+Dss6HkdUQxBpMLuOy4H9Y1xMJHSNtBVIM0VUWgd18Ha
/laRAIkLLTjThvJ2C8Ai9H4+ADO3/0jWOV6des+oKWy2r+WlnptMmfPjAMWYmdSo
Q52dUia5SLtYQLa4vNBxlvTfPiJPwI7E9K5MApBOFFTqSHkeEePhVbyDvunbYqeO
ZdURQ8TUcbrKbuc/7+JMs9bDnTGNX/vzdJXp53QLTgQuwOcnj2iWr3COrEUWfAEv
B75OUsXw9IVgdoS160nh1Ff41Mnqtnn6JmW7l5OiM2XQ/v9WEoF2/AZceaW5U290
q6bV1M+aglQUgeiPrUMuHi1T8+C3xhcpucgY/Cm4943BFC3h7+sNOOvvGGnp2LxN
ZXr8COrGhR4S1jdh3DQO8k1KgnFl/Xk5ctPattQiTEbOXzApKpU/rrutyKwp6cig
zZjAKx+Cz1l+EdkDdrhGk7MyysNy2woakPM47HeajAlKPpgX05h/ep/2RVX0P9S0
ZFyk0PKMfet4h7uL1kfNVQBuukST0wAtvXKFpcsrccjU72lAWRE46LigxTJwKgT5
7fOLFbEP6jRZa1/+Z9zFsqiGlcX+fBHGaaVF9AKUeCxqVEhCCTlyiPVNtrmtkHHJ
7vgmiZ8fJ3lZMSCgns42zfZ9BzdmUGwstimpV3+ef/OWuc/NwPuXXXj2rQ85GSJP
jElxx2v74wLhKTkLJ5ljUotZ6Y3gpwQIRgzokD+Uj0YnnFUpe+xKvJmNVrph+RUG
hP+Zh3YQ+mjh4A1+Cwnf7DID+UHAiZrSqiwyRZvXUu8WU661vPQ8GFlXzxNYeodx
CN0TX4pYhqNbpVyPgx+fsDAX3AehCly+tWofmjjqHkF4mjiL2h98l8B+QqGbdu8Y
RRGA5jXIjB+DGk2cl37bA+vAAycO0Idavlfxrmah87MsRmts/MdjS+RSCqhU1NYm
LrY2GjNJaxHUAAkV0xJbK7rXjuiBwIbrlfY/AvUAHXDriGMj9kJK+bR3VkW8K2xT
PARt6m4mKfDfUErstfS1rEQxdF9E23oAWdBavea6vDpN9yfB4QrztDK3AIQgMvET
tzQuP6HQ+PD9Qmro9kKQv7iX4AKfV70f8KisJMBK3PjfvhMGxLHQqEkFIzB9C1hS
73fzDQ0W+ifIBGZ2WcTbIpFQoY9yTXPtO5AcSTeQd1TjJvT82RT1ASzA3FUsQ5qM
FgHc8lDnn0S8owLUCzMWf1kiJuyN6yKqfoxs2y9kLNQsXxuwyIHRf4i9WL8TiHM+
Zb2h7RA1uaGc/mMoFlabc2rvFMeoQBLPQ0u76HVlqPaHAipVc4LI0eR3+QcGVmjT
AvOYDD0j8Q89wLnv31xCHBoTnf+tmOQFLUqEVO/ziO6VK+ZBVRdqv1vuq/0KD2iy
6C9l9QdKe7M2JmhCZ41MgGeecHkpZfsgwK/eRInvcLc7aNS+yIndHJbDpjYS8AwI
MRH3geal8GoXDIpqaBIszNgcwRLFPyg8u+ME5kIPLS4dShFMASO5UDkZkj5q29lJ
is4wfA6LnRcjzbl9OnVSrbDe5CsyuzeN+Lvboq2s7AOkmYDY/NrMiVEQQtkNVF7Z
kz/AOF3rzYl6A7/epPwpir7yysuklgXC31+ewI80fMI1yzlnHG2ht59CeAYhrkqb
vWsmNiGAmlpW6MXLEzkQARVlNCC/yCwZ2NIJ1uIhU+MGvm37KjZ9Vj4dvWGbl6vU
PGC9nHI49yyhZWFGj2b+XTXN4lqrWRJUwabtEQh0ao0c/I2S3xmO3BDvyqhNi8Y+
zh6Z1c7McB3TE8adU48vjPkv2piCKq6xf1xWDXNGL3oJSti3jlH0/NJi70Au0B+x
Rjc//TokpKWXgpLHuHlkir5TnBgetGqtekGUTHHSuxfVCknlWQC1/7Ie+MaSeEQL
Poy4ErWZz7OJuE/1Cm1Xz38RTRot+byf7knpnH63cdqnCyHxFv+dxmuTsJbrImbB
2ViKFURQgXuKtam4DDppPLaXez7vcvMYMHaXCHfju68RM58TEk5Hnxo58Hh9jTHL
EPgS2o77kE+YxeYdir4EbeOkCNEGNHwblQjhHfQP8/BsWgTQYnpuM7HYbLFxPJ9s
A/foCWghj+Taba7zWeEr1mhGWAAI/1wM3wyXHSswV8m6C1q98CvWLlXW+Ls+WrN0
XQ3he1fdhHVFtl84c23KpywFlXzDeMR4h6VuEaLNlTO5gq+uLrZah7TFWX54Ol0l
kSSNloPfgarOGCGuVPA/uKrvYBjN1F+u8plB9mRrcLnbphe2HtZkHKkrzVrNO7I4
Lqqg8esGoQ68MJ38GkPX/jrL3FzS7Yi7HdACCz1SN0SU2mnNSgEqa31WXSZxan+B
6uRmTwVYSVtwe0Xh44GzXvi1n/aoJ4zMXEAeQvsvfPxlTCsXaZ3P8hYtVOo/uVod
lGisazd+NabJWZw4pRVi9mJwiubyoODZ8rPEPTf1sD+w2lIMOLKT7nJVh9RAqCIr
6qAuUFhUdmAT9hzBRdCB1REFw7+pLiTi5VALNdnpIs/lVTI/YjmoE2XcPJCUi4rd
ZHCT2wDLwQMo80aWuvhMU75+tn9vgEUCTgQDt+T2FdlhA4gJ8UW5W+2azbo0flSz
8LMvhvZHvdTGrSeoILZgSVts+yrJjY9kmqtWvfRA+lCneU/+54O8Zxjjdqm4ARK7
sG+AcNGi+MGf5QxEUgc0mOXwSI5ZFoavJa2/SLTdG/7Z2poNufisT1EVrJhKJk5o
/qQqNZe55vkIkfrR+sw7fniMweND4ozenlqMCqgRUqi7EbF89yAYcwURoKoiEB54
I7dniS+4zAZT8tRDZAiJJ6pwIeubDDuwDYgh8R89mSVmYow1MXl7KHsj7ewq41+X
FB+dLS8y9uWZ0I4zyA/mHa37/Q/BMP+7WKPMKfAtm1dYh9p5DkKjT3lfoVePKU5x
zyfqhUF7yQlWI6mR7JKLCyiu9AjgUlQbxcxaFNLzrc0VUOomQcqHYdAPBq+uWUIq
xj6e36C6Qm+/BC7fvDwByY4Ax06FjiudH2TOlHOEd+2wJOMxgstJiMWH1/GqqPV1
XjcKSilFGW3L5+EAMNzHkeCeCWQW4agwTLrEKVbumxq8X3qaetOpBaLXdzN4Y5Tu
/gIsnNHsa08ehElNVbSib47Fd/sTArndkobeKfV/JcQio0vnrDIAkxksUGwbqxoA
HvOdMH4gx8hUcV/V35ebSNPcsC6NeihWS3Pgr9bDX10xxsiqai/YGFY2OEu8wBf1
atgkbtGTCrXHdScKr/GEhGR/DygoNG242ICLoouLHzeVwZTkxMypF+zMfWkDTCet
k7j1b8m6+qCEoHdt+9MVsjbbXBZb/lYhHD1idMP2ZiN6mbfcGpHQadIyl14f8UyF
XKGSBAlqj75I9RPVRWgSGv0B/PFqlmNRokMKgMFJpnCVV66avstUctBfSDZg05R2
GNUvPM/8rLPME+8zhlmZQZEAtN+/KmwKQrWKMG8d2K+bF3gd6egIcNgWyZnsslF2
u3yhkn5ASguaxWWE6eGBezx3j8UhCAbYQEHoXGTlCJXiQCk1k2uM1L3ZfrOINHCA
AgaWDhzXxoptubgXsRSPYQ0b+rRQxZL8KJzzdDq5RkNiRClNDtQ0sXzNNvvc7PGO
KHR31AfBcV4LiWcEpPwVN6juJecsqp1AOsu9rEuB8FGcp3YYIMnM7uWT5kHXAYQb
TGDwMB6eQGwClsgNIzM7cdep5PKFhhDwPVmfoa/7aM9z4cR8LzLvZMf9EX8RKWIx
NC9gzjFNUu2GI2RLEHSM9zP4xSkvkgChDJzq5R0A/aXst6mwC90SFgTTxF5JK/Bg
7C2mP5hR7J79+40TT83Od2ZO8khXpnINZ9CwyRc/fyTxqJoYA1RCZ2xJDw6jIvQO
YvEptUQ0Vkh4iC/ICBpaqWxjpHK/gwzhmXy22/V5bt6o0A7J3x77Zxf8enI9ahU3
+d9iPly5KMke0RwvDA/LlqyDtM0XSQ2MRcTHSsQJh2XwXq/Ne0QjB1/Gxti/nNOv
zN58oBhxEFt24e2Eld6HTmyXaMrDKOMVKXuZMa4y3xG4yRi6n2YSV66AxHTsayI/
ldYiUS4tVzfZVVh9CILhJ+yn6E/DA5Q5syXiq71wZmrZXm5eeVENAPaox88YVj1+
pmXG/YE6eJ37JSXK1cBy32K8pUvbjlYHHCAS1y18olA6BEAg6IhSQSW5Csxgfcxm
4CZMn3Ci5gNX1tQ6GFiRLeRxYzQCgN+I414R2TnOK6KvHjrYj8ke5nZz9nLfB3lG
jEhDw88lTNM3RHVlPVZX6lGlsh04hZTmxn+SiesWMskXKHSRdmqeG1ztcTl12hO/
XdlgUqLVpyv9i2AgiJSmiz9UUJrOVGcJkQcFhmlniRwXgC0pvC0zP/7w+aEdVh99
pV7rDKsY7wRI9R7PF/dpbP3KrNui9QHpkEV1A2JZZZn8bBI9DiJ0jVQXZuJF23iD
v8dWbdu+6LtojbA3uTsKjLQhJfASFWHvByo35DwuJtw46b+LKv9omeAugVd0BoqR
ZOtnpTaxYNl8MBxVwSJRAS5lPGaILwsF+wjHf0gdwdcMn/i72oO1wF/ZUkMf7eHD
5zp2p1TvpckWSBT6Dnv/iTA9stn6/rdnTh6KLx2oF+mS+OU7UO/13AuK7+2erIsS
paCdOxm8VPo29EYSwsTZIGDzB/DdO38AG8+LuopL2VdLwxPM1hc780Cva0IlBWbc
VZv5lzFcFKjZXMm/fWk38Hp56eqWRwhaulyu5WK1avOvq6x56d8xVurcvOE3uKWU
cM+VFlPcP3qey0p0xHyMXRcf+Eiy3lQkh2i0FuF2smG+WRMUlvESD8swUiXzrHIF
HHMyP//5/gxz2am2nwJUj2cKktJbJQPgOU02bq7hu9YE7AOez14XXGMvXpwN3li6
XnxGZtaCApMTeO7h3y9YGLlShr9ZB26LfJRkHRmBowwdn6bnImUgLKZYJG++m10p
yaH/JqpqfOizCf0HXo1znr6XR2exl3Q4bDcExY+UOX1OPmNDvRDDuKdUEorWlASD
JjdOf78EaRtSQI/ppwtDqJ6oIQbffuds5gK2Mzf8hArPi1bs3brksIZx6AMjlWjr
T/Y16clAZ4sIl+kFloKdI0oGU2CrsP+PlBRTqzjY33dlE0B0JsrUbJWAvMr0BIwj
u0HM/r830ZY83UBqIzawHzPm9/1A6guyfCVAOZ+zjxWe4/hq5LnO8yB5fT9MfN0u
nE5/eFwT50xVnunIjYTGkoOvJ/KT2TQ7Jm9Ti60FJAF68a+FAjB1uVGLghQwGqfe
MdpAcr1gWXsAVXey/PKsVSsLMQeoKhLDfv46VRTsUJkwY0Gk5GQdAtTnIfRh34L2
Xko7VtI48OOb5xTp4UD5+5k8/f7t6lsnqypvcU6wocY6hhUhP0DV7bFzPsW11HN1
eX5ctqkExbdkaqQ9qjgDXyLpfp5Jb4NyDeHaOM/h1gIlTmkBdAs0vsbaoTRdOSc6
u/pi9gjgPfmKzN+1fHu53yjhhdhqqKEeVVdIGbjXZEiO2Piq6VLGQkEd+Y/OQ8G+
jqjhdEeq7ZZkHPvkv1DtOQkhmbLbiz6b49dKBoyCXwPcn4TNcEzXQynwkXGOj9Jk
2u87cwWY9lR/08SnXPT9R0Hp6VzJf6vUDEvP49PK9t/Wn7n8MGlTtOUPqP7VSZ7c
Vg5ewDNnlPhyRr8wWsRmazAuG2JdE8+AF0AQF23ssnaqv/mNaIDjAawh3mHxDVow
9tMjLIa/zoWujDy+zGj9EUx8yKu4NCSbMpCxXqcOs1w8UmTC8Ui38H3TcsrnF5fS
o+J1pSpfUTnI0zCrbiL2hcpX/Mg8Uuk2lVfAHHx/fTlmyqZMR5Kq/FRoSgVsIsKa
dTXzr+7Sgqne/fo8rs3HyLAqKdoiPsuqNrjTGTpVtqsirJUwM9yMqJ+KjAm5fSba
/G3Az5FKWAbbSrsyEiO7YoUrcN6+G8jF1ofReniT/5RT+FsfqFjt1yy9KXByDosT
rb2fNzeiIc+pBqQ4iB9VU+CXYiQIs2N36ybBXRdeySV0vWOjUDlLIHJALPMQIO6Y
z9LspFYj6S/5LN4nfZPnsdaE1XH7UO5piKfUakDoqlGOMiTiLUsmhGNvp46UYwdY
eqnlUxYfMyKneyFgrd5V9/Qm73Nvrb4ZLmWOBnXbuUJK0NB+F0Rdi5iVWQAHOb7i
d+VFHhsVdyE1x3vMwvQqnzoqkXCphM3TkCcbMI46L7olyYP5elpiS3dnPu8X5wPv
3+ooYDLk7hwEzhqPwzecRoLmn5N9hgOAOli1QvUmqSEMuCPrEhLTDPSaRmuxOy39
vEZYY0eJe8rWNPk4dVnZraTB1k/yX4WGGXq2Mmj0OisLQINZDNn2Zhs103sEC9tW
7C7H1n/SdR1VRm+SFZ7KS1ixtnTtkCeufrLd6QSpEP7MctaJQkhEQsYJ0c4acpt9
r0MfQgO2T3nPpa3IseWt08XgUSdIYSzlfop7o9JaCTffVXvFVkWh4rHfdGlzue05
Nw8B37KJAOOflk/p5Z90Ly4jaNrFCtTPyHW326nFzSBmhb+jYsc9r4BSesvcWdYk
QzSmx0/n7Kg+AnOv8D27fdP31E/XW3vfuQItr9xV3Owu17BDwXqxBhc1li5cbp/y
tYJTIgj8tCUbiCzG8XH6q74Wp0Qt5Zmd1F52a18oa2Jg03lRhx1oYJpHR1HGDWmd
zMcYoX5Zvrssf2o5+PnbUrndTZKts1wjU0VnPRgp87NtDngkek2PSRRWmKcjn6mZ
jkX4Tow1YAx0tIXm4C+flPo+Dx+B4W1LShrbkJ0buoMnH9dqwxk9TWJY3ogN0pe6
3b/PcIjbPslWxW69bWPfM8Rf8TWTyuRhqfm1KIPVAZKY5rQvtRYy/mLSRPI5hHJG
l6Azykh9o9/8j7p4iSYP3pzt2tJNctUQZ8cSUFp6ql/yQUiU5clArb+MmZQ+2SP4
PdpAlEImEfWQNgT4BdcKCXrWSXSVSQF6AP0lW4nZRmW8GLoWN9qni9l/yi/j4N8h
roc03wFrn4TIAtXlRdbvR8UgQp9QacuEvGIlNenLwHqmabxn+dv4xeRQetJDg2uf
BYRQzZU+lv3KEB/l/Krr4HvmmGrvUKxBAnBksCy01pQvkRKupTuM4Wl9J+YkFh/f
JYa1e8OsT/fazj4RlrRzpuRBKLXrI0qHSFbG0lZm8HjbsBwi8QfmoIhLbNhJbb1T
rFksY+Enr6ylEht6yVP6/QpwAc7mqpNJiLRT0Ws6sxJGk1MvX40S9jDxZw/PJGka
kAsdNMSkHHRcC6DqdmLTJRy16SyaPUgCdGkL/hpQ+CXf2UfQYh1izDEvSIcEzTru
mnrykZA1cJFOObCpLaE5l3bPWX9XOtRHbMDpYA5U581vcs0Y26MUOKcSQHmPEs+B
wXF2mFF7GpX4Stqh6muLVMpVtjcVU+DUG2onzW20XbyXlus5ma46G45CGa3J0AQl
YzOEDmu4DBmiWvtqYE72YRRTcsg8CoxanxcSB35qlb2yL1BVqbJ0w/gW+sN0UsLc
pnp6YkzO9yHZ6mupAAZQCBh3Ovw5Mswvejofh3hbZaAstJ/0/3zj9fc9gG7WcTkz
ojmaKjD3fxH/XwSyanmpJ8Bh+MsGnnxzZU2Wd24lxWykvNNPUnhKX3aLegor/ER8
UqbEgrW3sfH7c92EY7nvBT7PDBOHND1EsenR7oulmBCB+33cbxgDYMhhljqZ4KLx
631F7QK+mUmfA9AcQzXQ5KFdQcZjsDmf/UCAOjgN5dfIHUzQ+CtdaoDUnwTLmYZv
Pc/CAqUa1m7QvUaRg8Qe2HNgHVU094Y4BUP2TymQeoEgLBjjswbVR0ClhLoU+4qp
olgOn0yaIDciQE7dEjBUxXUHV1RuUrgkFyfShUmWzQPpB2RGxcws0WlCWzMM9/h7
LEyZMPF3raMQTSKvYd1vkTleM1RpZL4tZGOCVveKOEfTJOGTxTSedfEFLV2YbsHJ
TvJkrbj+V0m659DLq3QGPq0etzF34locaQUBqqMyEnLlmS79A6+BFfmdnG8bwJ8p
pH4+J6nElHLm/UZG17UFY+2Vx+MOsE2pkbE02V5kVUdAWx4Ylq1PbqdmYuLhONE3
0iKA9OBTZ1Ue8Ezno9PO0S7SQ9djg7wxXkg96VpZlC9j+OD/UEFPSjlreMj0+Hao
ZS+0QHkSCh0D5jgy9jn4orqaOBY0TIblOhWk3t7HvhYmmAgTzLzLj5bAjG4qLh8k
2fYsVrSZEguh7HiLm4I5mhITLsNendWU+rApQh2ZggwOUkr7TBnjhViUChXUeMPY
NNX42h+m+jeDoCvDIKUnOZBbHhC0l2ZvK+z6CAbkqLB0lO39pnkpUjl+tVkpyi25
5HrNrLZS48DhQ1I3B/OtbejMUIhitp/XkZzgD6wuwLlHnXGxQbJMpY7Mg6mC0Kdl
n81+KYi5g1AFb7g7dAjpp3WOPJ/0kU4VoAcyixAwLfFyHSKNv7o86SLQjIEN+tkj
mHbioRVT7LN4yiqF6L/2pXY6+q0P/LPXkkIKw954PnbW4PDQd2Umrplgl+vtQkOw
ANy97SqjbCFouB+upGvbHdllFeS+fUJmtY04oH2of1omd/BIyDKkHDbktRq3QSn3
PugyhB8dohAg8mZRpfa6zBWhRPWwlsUW9JdoihWvTnvGRHJIqbq39+4f1JWSYvmJ
BjwjQeoU5F/+l0CBkMJkTqcT9zNV5ax/OeERjnAAJ/h8nGsTrvv8WZXp8eKHiFb7
A+zZT6P6s4+v/KDlX0mEx0+dR30yvjoSBg0uEx8pDz88d/+G5i/ErWeK/U+n14kJ
LBes5XPeO9JJv1uMsNhBTdFFt5Jrw1bqjD7mrOu8Bn7/kdHxx7a/WKTLBbl1GyZS
vuA8XsIAZYnmwBUGIXP0mMvtpkj/IwIuSkwrbC96N5KCnrUVWVGverovSJS6l04h
JL2vhkUDIQhkcsYbMG0zKYi10/45Tw42atyNVA6uQHIKF3p23U8i6tI04pNldkkY
DRMCLSsA+ChazvYR8au+u5AJ7fmfmqvtU3hsEhGermD5JceOJG9bDA1WccXw5FkY
G4IXetMpFKxjQtqBCUlIqRq/yxwMnINBfXYMOzl0i5vRxCB/OtuYcxz9oksMfRmf
71l2XUs0b0zV58owyMP22RsjJO6u46v5ih1cUYydidz0/ZI5wzx2RBx0J3Ir70te
GNhcc6BkmFVuk+AXxdQ8wTSXKsrYNZ1cPsey7ym6gSuVDTwliqsRtH4EMP1LDYvY
Y5AhvrpZdIF3TSpQ2DveGw82mcplCJI6yDzo/TQYgjJjCDItmaG+V8GLTBsV0nwQ
kUkGZmBEwtp6dwCwA9sTRf/JAkBrazP3LAR501iklHRorxfkrwT6vTaM0CcBMvsy
1ZhihHu8u6l7tlOixieLOmgBaHqhMn85ZNUcOd9Ob0Da5fH5dUbDq3q5lHrKD+CA
Pf0CL8TIxCR2kKy4ajKFgIKEJ8iDCDxWTN2+8x0T5m2SQGC5BogYi6hIlH53k2so
9+LC4sh9fXl9m8UMylYSPIzJ/hT9z19hydibFCC6OUzr0RDOb7ddfGTY4k3teHq2
GqZr3K6np/wo+qu92Gqylwp43tF4VG0LAXqwhr9X9J3ougRncFbxmh7OiErdcdWd
6oHOWeeItfPlN04pX/p4pEcv3INE1Iz9Q+JhMcFGGt6EqYBaAkvUxgwEbKOC9iQc
HgG3/KQqGVR1iY2cqwUwjkqV18xJZkAqEYXBnDR4TcdNndgRsUL1mk80NTR/XZnq
4127Y4nnDaRR8py1JIyuwciay3tC6AbbtOFxqjUcq7laWnjUxg+mBjxybfg+sIrS
LA3F247D1ZBtWtatutIIhLxgYn7FngRX3ZQ3MqmGZdi/jeh/Cyrh4gnxie/TlJhy
waFR0Rx556IILsjltNvN1kEuozEQnUP1nodlvfZJzZa+QL/wHQ6WpOXeOyr0p2yT
2axfkXsotIF7TjSwqiV9RXrDpU3r1hLTuV8OwqaupgV4ZWFx7uZmSGMw3GvOjMbk
PSolThP/agCXa4JZlTQ1uPIWNMNXlSSv7irCX/EaP4hwKSfOM8dOYPGG/2KIlSy7
mCG//slXPqtyCE+VStdZG3aNnVmtPKRn+7vPXG6CX4iUl4BWJh8j1bGekI3B85Jf
SSoS0213XGs9NlZXxdNNov5S5wQe83ivP8wDAQJQ+DIEsoiIQJ+N9ToGDDUbWk0c
qiefQG8gdRnZhIa5qAJSuc9YHi6IHYs/tvjGIhRWplJQlwpvNKgl5RyuKQQBVcP0
hxL+DT1hMckxKH/aANs7GNF0KaeN/ZA5z/0abp8H/KnAn3uuVJ9Pl4bc0XiKJme2
5LKpGIB0luxW+6RRUbBBNCLFavO/Rpetwy/aDY785oTL1clJdM9xGUpY7Nc+ql5n
dQ3JPdQx32JCJGKFwmleLYpLKu//ksRk4AaJj1mn3HIXqEyLclVWZnZ6zSvL6Ui9
jIFzGqu6qbU+otYGsT1vEm8XGUqx9B3vCVSLpxWn3+TRP5sbLrj1C6pwCunR4MOq
ekY0DogJMrL+X6uIq2HZQBzsmkGJFn3vUUKfp4ShvV98EdYCSbyKNKhPY5jLpIki
MKTxc93oe3c3tJHtD0UFW2W4FWumGRw3o/AsebQ9w6ZeXXCKRTKfW7KcxT4Tei5H
9lX4CxV6zhI1BjUhMnlVdMhFBHazXLF8WwFwH23KWkjhHarLK+2WI4b6j4rPyZd/
4Lc7od4cAiiL1N31wh54RXyXG90WP8G6z4lXLrSeA5XdMnjSfyD8dhmf3rfT/aDu
dLJbMMZTUakELbUFcIZyAMVibONBnJNGo7NrqdTYUXJ0NXuDhtWSU4lsLEw8QplT
F3P9JGd5i2oMt5LLpxnqiIfmDXnJxxA2iqso1UTFyAXAeCdswV8COOXyLXLJvtOd
lHFWLCkjAlLI815Pwjz6xym+t1hUQboNOEEbWUk6NzKt4472rv9/Kt5S6GMTJpb9
Jkp0k5SDYwFyrNNb91OHAsAoGmFkVLealmswZ3gK6fLc0brAEUkIVn7wvIW1kJMu
oea51MzmvrKGEECn06S0QtP2ROREwU75NOGUFP4cXsEAWHm6pwqeA4j7p5tuqEDw
okPp/PPWnKUTwXq/LyzPL+tGnTvxSH8NVUuNDnOFf3rN6wbG+tQh/4FdaZf+PrRp
R9aIL2NHr/VwpO2WAbLwS5NoCrt+yAA1HHdlnbmPAxXT+rXhSJuEXFm2nu8LeiMU
nI7dJKcifuGom5gdkjcGpdE9RRYidlRXWvC8Vu6g/D9FS/hhPMK7Jj99S+qfEFD/
k6k9fCGYffNm27sbktNesmHb2pPYBj+xEPaiZlvqDmhH241+nCXfR1mU9uLGq1nQ
Q8CherYJkaM9O/2fY5nb5uXG1O30hLKmlikhoZAsC/7V366Jrb5z3Knwmg6OhsQs
B+0lkYtlBXmy8FrcITFcnAEVwuKqui16H3RO2WPGcfaHYCbTjHwsWFQSMC0Pmvrs
Xhbf+RwJbIUiRVqhLs/kP0TNWubqfK0DH+tEceifHkO/YTnIFcRAm24++kOxVqBB
0UGSwgi4y6OZOl5J19JMIdTXBR1dGeF9gY6hKKZ73RhZFKbvs3IudoNhFd/OapZA
oZcty3Znofv7a64nj8pXyUHj4rUgKqGwAzqTyHYKhYTMA46v4MJWzd6jwVqqCgTO
g3QWt8hSUM0Aqqa0Kyqu42CDS5lfuCEqOUdrw703sRh3stf05mNBcNxq1FgSmuPY
Xmdd9XWxBrB4DX8GLfJ1kHJpGcJl3pU49/G74netAyKlDAbPzf2k61lFcJzPvW27
EVroGRMIiox9u2avcLRhVyv8EWNEouUdwoLCiWK01W7ag8oMMkB3FDjjvqe5HlEX
m7N3E8TNBjIgme292eT71p39CLzWYPMCMv1Xt256I2uyJtkqm6sIV//nsBu0RttH
I61PIB55i4sc9j526QMhDRH2l8HxBBOvfbCKiKyutW6+ZS8DTiHtX4c9IXfjDA62
/IhULgukZ9QhNFKd3XaZvkt7cCQkunXTje91KIFt3vQ77Sx/pq7OxjJp3e6DRAzl
0j5zVC+DeRFeU++9wv2fxmJc3447vG+3mmE87NxNBfvHwBOU9EHucdAVywrZ7KZf
1/EwaQRbefbv4frenvgdIOfDLfEiNNwXdf7Wk99JG9ScBCTrkuLS4+pWLli1s/gf
ls9yW84B92c6+yqTCKkv9x5v+EUSTeFa1vnRsNj7i612c0D5uEX9eJViAas369ME
rzehhKDtwQlUfFvoZS0sMTGg3FW1nEigL5ocIB4Bk0iBPCqtcDIIoII48owsjxDW
yYyBxqwRL78Upx9JpCm6Cv4x7n2Zw0aJHefuBaBll5EGcRkZie/ARzdW0/wYWViU
UslUebXu+yedIhNrlPe4dl0+0neF4O/UgoEPJjLFSV3qf+HyCuilnCEKFBHr0rmH
4VW9Zto379MtjixGeUChW9VVwobIvpCrbE5J4vW2zFKWnF0AwHWpk0Qp2ngBzi/t
ImNJow2hT9/WcqdX7YZtbQKiljXD6wfPgKPu/6SjxU7LLRsLNMcYeIFcqnJON7lN
mGaxphAKNM/BufuFRsrMiF17Cmj9rjLsYCP3pRbFFdXUgfvrwiCMmmyxpQqsK9ed
Q7w5zasTgBcs4nWxfffAZ4QFAuzF8Lx3PaH4xJhnJwhslfB8aB7aul1HJPXU9vWH
B/HQDg9c/i6l5L5Vbs5uwokJFvhSqoLiQ8oCBuX/KlRxdghYdB2R8YZDKz0pWLk5
0rZllqFHMguUuD12XvET8+TncnYnfhGR395pVs9IuLmAi7T3RtU7CqBjQDsXixvW
rYIX2gj8FKw/J0mPdPVDvnO0YSezVoupEHko7P3/teryVWvr3UU8R1qqQ5cAmd09
W+RkXO8lLS26qp6Uw2y5yjyFuSJr+JkB8il4F6tvzQttB4MVmWx232JrNwF4TZ6/
udU6PfkyC3U++YFGudlQ3d8kOAY3WGsoId2OYE/eqMZ12lDLWRcgIZndvJECBtTU
ndb/3QQtmU/kXynSWj0Yb2kwrrPIaK48Xv8BzCtXhXdeyQ4E4Nlnngw0F3KXckL4
p878fLVNzRfsVsh4YYfBwGzQiykPvmEmBqtHywaI4R7eV7730kTrLGJvmtLVgpcV
OvGh4h2SVKoy9f3RbWaM5jtYFTkFkGlX53KdvGYGrzYbLFosNzskdUhhD++yPQ3M
LneUyyUpOTnyhZt9NYYtD+Bza/D52ZyE2hYUpiv/FXsm3Ild5FgQxVLsmnLQb3NY
6P0prTwXmjOnNd3/xbGe0NleWb4V5/BLWC7UXH6mRItDun6AL9wXyDtO/juDO1Et
iAQ8rIiMjRtlcmUjr9ky15oNubHh8+LD4h97q6JUecdh1R+LZ/iDyVYcTC4sUtJv
Rx2G5N9vq/6zdLEblqeoXflM/ZWP7USlQa/3oJCWcV8Nx+8Cg5ceX5ql2QdRUYfJ
SN+9M1G309q6bE0tKrHBVQ+3J4eP1iaP7UIY64VfjRYrB9MNWG72U0V516H6jpR1
GZgOLvBcOvv5Kx38/KCgFwkvR9HsBXP/TIqkoP0FcXQd/YPMq8ms7AP2wcmWCqjH
CaiUOqbe0LcC4zt7HzmLNeWM8nX4fUs5zNdtMYroAJe7RttFl8jbLG6IrN/gNFb3
Ur3QK9fymg4dAZNTL46vqEeMH0llly3nH6NHAjyeqfAsDQLODYZr529cSg4s3y8r
tw/5DFfDzJpdMU3rMIrg57yrF8gDAC8+fAo1AAfDeXIu2cIulqGUPhSgmejEi31e
RPuCVQUCK1U4alZmK9nhZZXtzoNyjJUT6cEA5LxsutJrFxHzIjTzF+5AFuKMTiUn
VBnVbFIkzK6YKF9fd0pFOt0yleV5xLSEbFO8t47YGZZ09CPbLcTQ8KyugyGmRNJ9
PerdqEWuuQF3NM5/8tmgSKJNFil0t1FR+B8AHemkBoAE8tapyjBRsn+wSqgQCxN7
IODO5S3hc8jF1cdipDzxvFk/7rYZM7wewkhLRcaburVuBCfcdNklpXA+c2zHD8dQ
bUs/G/AXlrzc2qBmmpG8mo/fqy0nfc4jlAeFIl1Go1G1YJkXRGP1G1XTab6hEJo3
PVWSNcmWaVBwnMzdocrO4gcaDEHIrvoKhaGc6DM0B7BwZakYc70e2VPutNvTyi1U
eYGcfCMGEPNaJPfPn7oyygQef5YPnP62ha65xF4zRB/htexDwEp+J1iWIZh7Kd2C
Kk+tBH3jlwfL155oBFURe2N395/Z3BX/DmXLeVxlU3JW9MfwgzlIn0Xw/if0boEg
nmN7BDxF3RQvEMOqmRGfBCsH6pSvwAMElWO/syrVX+3h2GNMYgvySpfoPII05JUc
5P45mk9JkPqxif3Nlekf76anl3jJVz075O2I8c+1FUJ7fgVc3sqbX6AbKSYZnwmS
ApFIHqv/C8rfRcn853o3v9Wb8O1n3+V4VcpO5fuvg6F6up1yqSYxzqujyrCMgx/W
tXxOtnrF2zFmBdgI5rStJp44WSa1g/ZcvdBbk46MKoo2Hnd3Cg2UXyHCshZ66UKd
j6kIfD3OA88Lhe5AL6toKzXQWJo7BgodBsLR54L/2u0DvU1QMHGsS/hkOLSwd1Bt
YGkwULPszVJFSNYjKiIJGdIGaBfi7WPOIU7KLDhEHbsg+1seUOhCTEPeCWMblhZu
LYE8iQ+TW7OQIOueLMicPyK2k2ISiFt+n2Hd5mgY5BGh28fUwQ6txwPBTExY9ZW8
aIV+HgtTDRcSNrnvZegO8k6WH4bKPBxQhQw6Igc5hkpBavJ2yuQdu8ZpVNdgb82n
zMV4oVDDGPFA22vFUe6GTVNsHOiALv9yhFa1dvjanVoaQMBdmzgsMNu2ka3NOO+G
OfPCQkpGwIl1lxW5LxcSiewBWsNt2N14/A7s4lSCyYJ/w3M9BPfMJ8Uur6lTXf7A
au/7D6MX8aFtTaj/1jwF7lQtCWRUIN6lWgtSpe5ZKeEi5PniFHyGQK8QgMlh7T7u
WlMnWCdME8LKPJJPq0KR7AXZOu2RC+4CBsLYbaqlucqX0xs7lddKIqINrRh7aoUv
okVWp4bDu86is+Px78J0YMVNqLSM20mOFxH0lSrR1l6wWiWUlphB67rIbsvlojS4
sGg2v7lRjYTqgnNvLDRS0uxtQLZrX1fd/rkYPw8P+ezw0e7qKOri7AvbFFzVbWXI
fUD5xgftNR7mNC2k5FV6vuHgkXnlANvH9P0O73UWg1zc9E5eHSLWgQoMPmrm5Xgc
8X6gsKO1oZHXS+WP6xPnIFVE9YJGAvVWiHWTeuo7x2ZrFRlc8wpcnUcO4b312DdX
u5cAuVQ1ajpaaBN1rHlHVwzfHKhsmDbnLlD4BGK1xHSYaw8Mu/y+zuK/chjAiiqj
OIILj3s0H5z3DfOrwbpZX8YHAUWCbkMZQGQIUritFVoTmWh6ErVoqC3jVCe5y8My
sSef8Z2vLWYbAcjfx3DL7geD8Q4U2dU3Ect4S444kxs7sKn19Nu/lwlADX513f/y
C0LNnnp2JOV0202fFVUkJ0O7nvvehamJevDxTU+CBnn51f3f5Nbbsip7Nw9R3Sdy
mqmoplN+CaxVD2jHUowCjF6rlaOrdAWIaS/WnzGIQLH2bByTPuGaVKuaaYhRsQAs
SQfHAlB4jTAz59LDk1p3CUR4AeoG90/EMiJxOj8tu4GjsYWzDGcDuEa4r0AMm2vb
8J62EWy3J52HRzKMbaQWqgqE+3xxVF5fdUHYCzkAn5n7fh/N0vC7LErhOPd/NczP
/L/GFIX5lCGB80LP5CGCploKiMrD8jwv23BFkaO3MC/bjIYzKjHiXhUW+y2M9Ien
FX+1OFh2MaidJQI+k0S24mY6tnoz8pBM6zNlicQ8Ka7yqJyw10/E6h3G9sSCAz2X
E+he8sS2DQd561L13F5fCS/lPVKZ/W6AbEsQFgBoLgBnIzYuibnVqQ2fnNJZFvE7
dHKKM6q2nULNnsPQ7fWEb6VSF6CCcQ5YQaRoxpl4uPdl+hM0tr6tsdsgYqh+go/F
/gaKUPzCG7DxfO3Ad75m7Knr2b0GOjRuJtbXYjDs4PyBbDdDs/L4sikyPfEdzget
ak1JiUfx/XtcOl+qg9O5zjfrNGV52w/wXPHDQb+7c1TNcPoaOYWY1uDNhkmSwP/A
j85tVp9wX1jmz9rTnTnvWS4OutzYn75lf4PoXQbt8QAU54sRhwaeKeXuY4r1DJkG
k4jk7uXn1cX77DqcDOPyab73j74pYKtZCAtMYXAxRyCHtHBvgJn15Huruy4Xo2+C
h9jAy1q+JEV3QhLYWRoewtj6r2toKmkip8YTcvkpfhtDrc9pKl6216yg8uInXBqP
treFukWHmuVsA04GZ3g5KZYGtt3vKQztk7uivJchd4I9eqiEabSH+qxFraHXvXiy
Fs2TQiXSMjTczgS2Q0v1GN4P6E4aKVCLbgywW/OwIesP0Ges8Fe6KwccNlUrJG8N
l63oObi5qIrs0m9V6577MwYsXvV081wE3Cz5bx5yfi1T0+5tT2lvC5Skcu7NPkdN
e1awtM61jMNvhirTDuujF/aCxWGDKVHjVv6NmKrB5mBYqI4YnY3/nrdb+wdhDdb/
V58s+gX3TxgTeRuZ18MB+XT3v1KEj4XuHHpEMtStY/P9LLDx+8Hfx91KNVWy2NPT
UWcw3wtnxRcyCbnvZG2MF7VSk5ZuEonow3w9m88+2bK/1JZ7zaofv69notUycF5e
T0WQKC3dVYt6J+sWPbhJpEC95JyAIWGx0A/8lrwzVP5SH9uyx8ssZFrk0pV6RLvP
Z+jC4zQDK+UcAGzfP7SMrzAQNFXHpBrldypXqBSOeyr1pi4ihVdhW0HSrY4mmGZt
Bnu33GXrXJEhHH2TuJczRzpyb7wKx6qGWgodFgHl0qc3qvz4fMIsbf3Tcix8nh6h
PhC71bnUHs9ntjzCcCZBdHXNPy4edlYc7ZIJgywTFtzY8oIaedhO6Hf2qgVZWdSv
FhkMkHU/qzY5I5FMAXNNl6rl3aZ2fSNjWxUvTkYsm4f8SGqURJGbjJ7PoB3Gne3i
GI4o3oVVeAm7BnCxgfPoh/VjBcrHc2GVcxOseTgffUXZKW4uUCPfyxOkKEaNBCHn
HJmoI9fwClLbYG6IIb2+cDg1WEB37mYbILSMVoFGUosGzdM7poXR2jssVnsJcTh1
ClkFHDKnKcDd8EuZMjjFvCRiud54Zo36sCsapXSmo8zqNjoWkuTXtQacu4VDoKs8
O+f5pGqN4Nb6+4IawL+/MZ2/WolfSvphRTHdp8tCrZDHo3SmxMcKFWLV+oaFZkpV
dRn44ItZShELXy4JZU/tbxzstrB5Do8NOuaJ4/tF27m/H/Oiu1hvXBY5BkR1GeVv
eJOMOEnKMs8I36IxYkuV42HOK+8T0oSBjBu6bPerfzj6Jkaak09J30ET4U2cpDUR
ELgRSaQyoVK1uiMfhudGNsv8A/1HqykZ+URNXUZnwzbboFQsIJUTmTcBl78mOTyY
5Pjr1Xm6x58aDdAbTf6hqqc3aXQQfLG3gvIFkOkyhClE1KdONqu8PKKg1TzhYkmA
Mvf++8I3tfsEmq0sTCrWUBl2rXrYJTT6AgT3L8uTth6ENGfkPI4nHCTUaZIxOR8J
FDcBYUH41iJLUGEiJrTGIsVBI7mzrSIkxgTfY8tsAPkC2y20Zmh+NomWkPCRP5Q4
v1zOmBbwMPXEI3Qk2ZF7VoLNcwCQmdEHsBmjo+C+Q7JkOxArtiXJoyFPigRK9H5X
gAXAdvneERd/NGXQOsgAyNV2cXdO3fermjWMTQi6tsH/H8Ad8qkpMbAC0mX5uZ/h
6nfR388M6Vy4OV/aLKz0pEdBYx3/4G6AzMUxZvZO1N9XG4PIVp60HBuyC0MVmzNb
RU0oaJFF4cSmtAp+WU/VHICCqGuieBT3govwIH+8cff0jXnMCtPyvs6qgGuh6Uh/
UOiyZJ4fzvst4eRL+H+DtYfJhLQ2hemN3A+zBlFa8igHOG9iEboZCZ/M/l6Z0f9T
PIfWnrvFG3Bheb1Yo9/XICz3PdkiOnLQ6S16JMSmBwECLjnEs4KGJqJaaLMdoEzl
kjkTYZlOEFCDaGPZRm6d9R60UQTSKArnJUiNzSX9JNQfwo6cuwcQLjAumJ3mBgrf
HPwTNcuwj7OFPYIuEb/Q6aG0raa7dvDXwHIPGqJz8VonqJx7RM85/+ntYfWKJPHO
ATIHzYn/JSE03Pw8EUt6kNzJFov4l2nJegNZTJp1LhPBCQvn06I7GxletEIvvbA0
R//8Zs3TOyuKfZ9AidTlT/TVDqKQosxrgijAKovvKXM41nWCB76vy6arLdGQj/CN
RPt7DPpnVfV9O3bi4lk8L+MCbG57p27JHcF62pKwtToH6KbZ1cwKRT80xjNliisj
3673TQmk5q56Z5mDHquDOP1aAgmOv3/GBLB8E5V3PZ0ex3synchCOkiu+lx2Di/N
jdOHYB0j2bKKh7ddxTFXip4/pfFARo/JNT5+TJIw1lO/yAElJQI5559uCz76b75U
yxr4FoeR2j8tQzL6WtjiXgPhVvSCYmq8TYX5hodqsQu6FD57aQvwmbF/GjvzLP82
Sp60pRfziXudMWlwOtSc4F1Ff560WdGTB6al1Tuz26YvR0noPE0iDHKqKSt56Siy
C6m7ORRcAkVpbbUUp7oupTOG6UNuOlykJkhQdr17FIIxtvxF9ICWUJ4LO34+j85T
VK+tEZEtbU+F1xlFmIFKS705g1xBCCTjy6ETBbv7KhPqHSE8dKUXoW0rKDPKP0Mo
Ru8WTF4ypI1CG56RJj7arrSApNwNB7GcoygfCYzdgRr4tOHUbJKTYW8BCGYAmJID
dhpu/zK/4KUW8w2VUI6FpiDp+XKMeMJcUp+3k6c+kZ4zvpXq7+XQOU0phhAfnV8C
uJ3U8uXlTXVrv11UaBEeEeoenAD7VsFOi5DAdfq93hepqGvWWoC3FCn9FFQUJfVh
0LzOtPQukYoHDaQVZPfteZhbxVvgb6RopQdQJCDI7+3Yivy3loym8dSerNSSEKbr
udRGYjFTUrlOAmTpdOylD4b7URF42QIygTR3tjl/EfZjUwl+yNbiSVVS0iVDRORX
gZ5Yb39mvEEv4ic9+i0aHC4FDXm5diR3uGuvUrGOh9U64vXc7cmajSMtsJMgiA/z
qcCamGrkICXa5DenOgj6GwcKhMoA7FraP9NzSG97pbcsLlJ9ytlHYq69xnKw+Pp9
vbk8zVqFmoLt/3mW59TvXduzI8mTSnkLsaq3ds4Jdw0oB7i+glpeMCPAdZrUZmav
iA/0B3pTKtIGTMreZR4g2OyEQsQXsDsa9v+eq8TcFOVudkTiidsjaP7NtnlyMBGb
dyCSzEMBoJBFdJPI4NhHM0a4qZTlOHEbxyX/9bAO/1HnP5QvXTwnx6A6BfQh7s4N
07003uG0QDlFSEuNAsbhv3I5fJ3zCeta3HQ6iJo0ApsDh9hog+sW92a1GkW3+YUA
KFvS2IhwzYhAcYKPND48iE79BQ9UbzFI7ko8s29H2EtG+3OyJ3g08/jrfToW4A//
cSvKnUDufCPL2gmSl/f3pSMxPnnG2qqW243xu7tdnCSYrQ+PRh6MN0/bEByI4AAb
0bnWz0oGzjHASHCuUZCyUDPRUM77AQZPSviJOYsHPBQkCBRI9jvhfopOj+8LEYxp
K2EnjP6VSZfaqQ8Ejd3AsGlgLivcJerKJkHDS3HIvFsJoznXReheRlW2t6BUyVVo
bWLsweRfFeB4yI2sSZozGIIrs2o7xxxL81aWA3RihHEwFBCMTChAg5JrcM0gqUjG
oMIalmFDiJpXgCHRbNIeq37dnWhccW22vSxib9TLtXhqgEVGo+4XhfOrQrogqYBF
IEollNqd1rUCASJ3XqsGPdp7WOa95wCYhdY9sa6oPGiuDEcF6Cll1cgIfe8lfEXd
k1IGmF9BkKfU8SF3gm9WuIHfRdxQYhz53Z/uqn6ydNhDUrlK6v6rWCDheLux4Ky0
IS0CU6v5wNdY+v4JsoN7RIGPKvN4618sNVwVW/iG+P/7KY+dAyJAbEqGh4X3XaBZ
p6XE0j2bcZVG9N0Sf5jX6pd6cYya7lf7kKscuTFyeeUsgt5V+PjwR3X8RzX5FLS7
szuK2uRcrFylQRdYKuok1miNtpkcEXn+ZD/89nO+XoZKLlrQeT7+dkem14Qf4eJk
Niy4kES/pEG6rt6oHCWVfv4CcLzQKlwigu4JFHrzh7GyIPoElNLxHDGePol4xw3g
+GmGdMG8bQ7hdSwnwaE/fHpXwyS3XXBl0En6jKsGsOztI1L/DFTBSId/dHHJ88wE
AkLz5Spay9fuCZ6CSshlgBTk21SqqIM2LildmjngGhLbXJoUKOGkcNlV9ry9W+SH
bZr4rN8EUbcdCHyO+4ZFytmP68nkrZX31wZ4IeJGSUza7/WZdnwoE5qg7yQbKeaL
aRToJ6iq2DLNuLiCVbHEHDB6WLd+VZOWooQiwPQm9iljka4Pe3xA+UeDHYVlpuqh
8STCZxqC3fiVNcCPH8krKJ7UGEf2BCu3IubGiLwUWIh2yK90mlPSd41bYRDV2dRx
U+dkg2pXtBPQ9z1Mrd8ZXMTdOVL44nwrCdr9xA8rY7u3f0DonTkDNmAJn1Oi9vOE
gdU32YvvkBSy1vg+4zZBCPCgqxIexesvEaztbCTIdx8imuey+xr9cIEnpjlPfAuL
H3q4nHZQ6RHQ6+6qzc4ROsPpTu3iVvXvuCNYni/u2yNEjH9njzRyQE6uB9Z2tXLj
DBdnvj/ARH59ZoWKaW9+lOhOBbJKF0u/XJyDbVJOj6OEZLjjB23ybjEMi5leVHAv
gVXpJJeDk8KrlNBNuNmjVI68wihpzeY6/cKDiX1VGIfjW/LJQ2vgv+tbyZR1d4fu
EJkNn5GWQ3WMulj1CKKbZ4Prh6ia+fsLdRUy+QT3A3dS9RmjTUBORoVKuEnbdS0f
tWVumjJwH7ku72taMeDa5Wln/9A8PwIvUjqNIzTLx9yqs5jKprNrhkE3Q4Jp4YUK
22ANHRzkMYlbMCIuynDwKx68bFewtn2t18VrjZV/VruzjVZpbkx2j28dxjQC8pb0
WlXdn5CqBX1SzQ7pwxaLyWPKP6zhqxTjKrBdrlBc0Ubg1qy45uyDmsL8ruE2Ibjz
UopAVkgwxp29ILTmVQGGgGXH/L8+p39bmF7LzGRphG8o9wvQQ3+y6wwA2C++Vl7H
7H34pk/ng8NLmqnxs3iseeDBAGtwGM2Dja9RQZCIBERJYU9rpCn4AyL130hjybFL
CX+IE7eQvLRlgbBCeFQism8TEMn8wPce5Joq/hXUWMK36VYVkyJmZKWTTuwXIJMD
tbUXJJzXHBRIJmPYMX+hJZu5BWb3o1xVcudkWIwSl9jwbrs/V3SyYpVQ+MI4XGXX
9VfQfnqhBQCZGQJpMyL4yzv2c8dtnAP4PIQ6iWFINUYP6zLLh8CAIZ4MxpKmFbky
Wf/JcEgpP9+uh1W6mACp6Lmhv28KxKWv8MBXU3TIdmwk1pG/QqumzUdafVMQxggW
nUSxTQAPMOpJA1aBfnEr31bYDh0vTxOjrZntFMYczAH6HSTAel2j1o7r8tBWJ9i/
vamRSI0vEkrynJl/fd2PT7DZCCdHdgXe4up3VOE3Qag86q8+d6djjUmN6q7nQUct
VI7KkAn9a4QQMcecG4/jqhfvVh0q/A2U52CO6Rlo1TWmDvU3FObQb/D3yhwYxyx/
S6NUNwG8inqes4BlXSEtNthMZ8VYxgE0o60dfQwr5jPoP8ZVQ8p3ftu/8NSC7zpy
LxTWwkGKP4Omz4H3IODo832OBaznbOdAqfQvG7JIWDoV4+ShiWwB53FJfhbRZRzP
pflnD8WMIMi5/Q7kEFMKXGoIG8kDDHbO3WM6y2L7CSRrKhVmtzzwiNgzLa1UCD6h
xAAwBDmTxWxPLXx3kHK8ouUw3WkXlUh/VhFUiRkjN6rQW0Tjo6rao4dmCpVuDMSC
RDHNIZ66+HxyElDAZzJyFi1CMe3/7e2ZP/jhl6RDTMMqqRi95uA4XVXhp9KBfLVg
+XKyiFiRolDarTyx80Xb+gS6Yl+XCluQn1lHvRyDIn4GlKSJf9Odgx2vsKjIIFFP
Crl/QdyeZTpt2Gx7rrHUuMJcrcoAux2TFPza/g9Zyn6EwKqraHNY2QbpY8kGARHq
ijLkiaKPfY2zi7f6Ey4iKZFgCzsSqvY6vkeurZ8lo7Di8x/pDFPw6G+XrCWWzToG
/mNVZknIizmatQAt308g+G69a4O6fRJa3FrdmPHvg9Vg0PED5G1G0mY6QTXMfyxn
7e5R0a78lagR6TZ9JTFFyu4HC7b3EJ3NUw/ioNbzRvYzCnwt6b4l+0yWGdmFVkPK
+rdMY5hdfx7MnjCC3jC9xOIS0hl+YjJmWU6mDkI2vofeXU/81G02vB8klVbiL/Xi
bqQzzrAvunSYY34oDARKJXjaEASqJmixKv7y6sr5fqV7gj6cegJY18gre/2KMa8k
6RpjgQIVHB60Xn6wVsuG2gpFGhNW2lyM3feFNGtKhmRqdGioEm+BAqkgxvyCPmh9
Y3u+AU2/a+VaSS9dWionWCSzRlts9dfW3CrCPVvNxJ1EoD9Bngkyj5dY/UlbccQ6
patpqcot5jaBiyk7hb/nSClfIu05NguL3ApK7yJMm8SX3xcvqnVb388aMrfFwecE
+p1Tm9moHpJoGKIm9LklNE9zrjI/+NkIofrBjaCSkxj4hdqs8XFQ/LCud65oWz0K
HpGQp2Ii2Og420KpeYKjNvBJbdqLm8X/iNdX6UPyGBU/1G69HHeKAsoKIdZKsDMo
/qj6/TbePcUSEvG72asaKOohOYr5hxBSs9XcUfWhYf1jKUnqu1Awmhn2H4pX3jef
3bFErhcNYlbWTYoWo5WMnOnYam5rCCdubjg0i4FjKUgF80Ulqq8HnZPn4Bczaw3G
otm0dWs19BhIHEGsuDD3iyENfJdlIfeLxhDfMWXWJ2aAS/Pj2QKr7dDvr0skaiNV
MIQiiuKFyFuAgUOdpxl+hHs5aWSVwjUWKHexe4rNz+Q6qL/m+8we+JFbJaQ9yBJ/
NUZ6EmwHQCMD5J8NekLCUKjqa5FIN6Xs2yx30wjmhLrHBx5aMsrRaiguaNfeQ73h
+q6Lt4gxLl+JTXAAVyHnzfbjoUebAr6w/ih7s56Z4T9fVeQvMCKmm2vdn1FOzHY/
EMgxdEHTL2ya/USiDmkzDRov7qgeptat54YLdSlJ065s1rposOxGJhUUAnyNfiG2
s8RDKhQFxf0S1GoyW7fwm2hUZhI3G2ZGpFkR7FpArzBqU4q1lp2ITulU+z6OExfv
cDMK/9vruRvCBrYMlbZx4A8yxGBc696QeRVHnJpbL31mgKJuoCFFWrNwsPH8ahyX
QZXhexbe9KkuA91RueJGVHJnec6VS0YIBhQaLvxUhbhpDrPqevjF7NRbhi4fdptK
KxhwQzh+BkiQgI/7w9zbBD1lzx2tBbPJ0MaUDO6jMkm3jet9yflAQyPLmeYPFEGp
JP96ELrXqaqBCAD2e9s9gPtE/VinHddaLLGA4zyAQlIgn6FxiUaMIZq3xtDm2bA6
NA67kRW1PanFxCwanYMwzfrqTzpLKjm2VsHQTvDNWn99SlogLrkPhKuUNBVcvG1v
73pd/UF8oCoU9yxDRcgJXAzWY/nbi08EZGtpKHSwAzmhpOwrMFvQ6GcO9eYt1fuy
j2wo3Gtx9c4bjctPeJt02Kp402FNO7uJwy6PPYClxbjwH0OzcV161NOpJCd7qckz
Sj4zcqj83xTjt0NkLyV5pG3Bkv1nHH4t0IeWwRaa7lGkDYje9Tqcbe+t+DHrkuCD
KibA7es9Eq0kf8kq0pk1j4xDtySUh1LL4qlYrwZyfgwUYFVShlaWoE5xVbX5uN1T
RexdINt5D/MzKiiBswHwQmt8eI+cCkGk0Bf+KLPS0b+KZeKrCof88Ag10SFkOi9b
f7TvdXsk/Ljyj5t+n9ED3CPhyWfv6DDGj+ObGU6A+I340G3MyWIl6twBL6cuIEeR
WEF8vG8uHPu6ONAyroXCX8StviNrb95MX6VBHjH80CQy8V9tlgpThhkou8aziP46
rAwIXepSL3Ni/I0i2VdoHEsbNlK2qwFxup05Q5CFuTj4V8K9NgmOYsDXTilMhDSs
gzejh8aIHjs6JNkNDwD5aWYwgfBzZh/yt6Q67wWxqC92gfV+4uFJiPfF6kV1/P4d
LafCDuudW8UpSgs9MGXa3QeOQuQ+hqexPzNsosu7ZThEMaYDfTl7iw5RtAmu3qXl
6thUFe4/AJg8zqornGQR/Q9COFqgeVDVRQZ8ZEB3YJTZhd9R/e8KGiMQPKF+6sHf
YGeYtp3b/0Us59fWNiyd4ZiCRSMsi0UnITNObXVY3nl0EM5DAKJmBL7DA2n4kzYh
2nADA0BQTHVi/O3oRxW40w01rXZ8MK2G4e6W06pah/Ta9piPH6Nfm661pPHLDDcw
xaTli53S1EloPDxkBmqg9CuOSBwjpPng5901UaqtOlwiO3ucPUNHJVX2aBStmKNC
St6UdjdGHEOTfzTxBdS2ZZO8M5AB2OIaR73rm7ekEyhuYbqsyxc3gDxfmOgsqWYW
IE9uWJ35eFNEKNjFjMEpm2VyzjjgoBx62aY1GJacBGYdx8oMbxYG5LRQdX5QmUnz
747TuQYqPMElYBXONNSzIC0WLf2sxoJYjRUrCgMqRxBzfWjDdT5yOqH97ku7L1iG
2fHQTjyxWTYVKn8GUjmhTQv7gGNNwi3JZ3wgveu8oijLbTL/TH+nIn16BrDVB2i4
dMKsZeEXm/KacYS8MLeyzYwINu/+gdd+LjjCp7T6kecp/6cOjvkMA6nTj+AXDclW
ohIhnOIomMZPvSvR1bKFasAHgJHjQBT7js+JnmLxIgq+PMNZiv6uF5UHs2rnErvD
5B1qJqUtqPNS7C/jb7EOtN/1MD+0SbMz0plyCCBDqs2ej9ETA3H010NfkLWV8+Nw
WIKMPnExxsbZizWH1iRLGpnqBlixRzCbTo/VLOwrlvmy98TTNbxavT2e9XwZtbV1
YsMv7ZbrV+8Bc7s4gQ0IYHhj1ggym/BC/5Jg5eHkNNSCWqC0FbD+pODejE3fGBPj
Kaflf3EInfm1VSZOlrhZBxNAR/ap9rmNw7PmfSZ7zBk7UMFJxaJzyblPXILkQGzy
s4xhSK2aqeH/tpoZb/WE896CYkiHJnH6qc/HC0asSyyPALx4Km1ooynHzmwWa5m0
5fc5zgEzUn1JOBbpgfgcse3lAb0qQ2EDZ/88wStSyWYZpNDAP2xKO5SPwT5KongX
kQOykA7qBcZ52i/NHj8gLg8nN/rktr+x29uH1Pt9DDccUSjSEqiaB+hHwoLrugGu
YBsD4y7wLAkjzc8jwOTOtYLTVbbudUJWC1Hqm3ReBlt4UlK2L6+/RFLPamphARvx
5rTcY4lqkJb3rs2LC2lOZwi+I+P5bGfEY+OTM0VqctZvZ8aRI77hlxSElGt4YAHh
lIJTuH5g2PgHv8ZFOVnhttooYBJ8zFpE2Y52aCKD1iyj9JHbJ7iM907JFm52STLI
t5TLRDK59OJLfRlnTEugDYTrbjKLppdtgKWXK4O05F+0whHWX2hMqHRu2AUqWDBX
wax3bQLisGySyjvABdh3uc2AOItL24X2UBDvecTvXtjXaSeBSOfxZdZVBzyUHpgQ
5UMR6gOfpvE4cmuo8wxuKkPwnnpaHeoF/w0d4bU5YYB7/9kox14HxeKH5FzPWxxc
hfwz4XC0ErlV4o0xXdauPqPTGgvkG/Bgp7FWM2d1T1YM7v1InL3y4gmG8FyKQ6We
9cB61hWshKhWu3qffJWCH0UeZePBW9by/gWeykh4GkHbhW50QsL0VG843FBpU9A+
q05cf4Fl31pGhUh0BhA3x6kLqq88aQlV+PaHGxW5G6dVqzMcGufRmXW6VgH2tUFj
s778HhfEWS+qUHmwITX+oVPf0wHszccMcp3SP+ovHq2wjsZ8GXF9Qx9r02iD9eL1
DJWJJRNjAqps7iKwmuDBWKLLYZT6UiQQ91b5LSys1wS6Gu9ONks0e7MztM/4IOdl
5LJanWuSJ0o1kCKLlHCMVjt6+ZLiMHHwQKmREIEjIqCDKArBGQTGvbBTI5CvtADY
RGqPalO0nHcq884lY8OPtW4E6kmPcYioNZ+ncgP9S2ZojNQkUMHGPJwec/brem0i
X58JNU6bnmEQOPoZRWxYRpaH7AK0n8yA14KfIVovWf2QnFmkFzDRSD6hHsLEGzxG
DvUpt3qZYjQgRLCIpDra8RiS+vEkeK84TlAxca3LF3AWN/OCnuI0k48IJutejBay
gBDIwOpn7meydCjclay7M6/E8RpkTae/SwDPoIabmbP6B2hh7Y6yQnvRvZEQxciW
2T1UgqALFk0YLMzWtgNqkXWCMTg0kAFlguMWREBUhmqMEfrSRhMz3w35BvvmK9Kj
a0cIgN+MFUHyuBrQDR3K/ZYuY1hY6YnBlD3Ir4QjaZwP+0MpPdh0S70IIkbCXnVH
jHn7jB5j0Ez8DlAgssD4ZaxlUvhsLmqFJ3k17qt9EKlgNjOejvoKEDHb8s+lzb9n
V7SEzIqGqXYOGFg8fPpGlEg/OuchA1T7w8kHbvlPgXgeC2pArXkhVeK4Adjv3sYk
N+rbaxpiilXxbdZk9c3AHXteb5usj/mU1fVd/4nYPLz+ti60VELUw01adZj96tGh
Ar7LOgN+gtprNIe4ZYUOWnNJJPWfd9+TUIjG3lv7HBQkUcxW2vRuMNje2x6mo3EU
8+P/wah4BoqSYnWU7lE+PA6IH0OX5zciFUDydMVaVcs9yTqmUKiPSAZfBLWdfZNJ
s4YO88iGAGzUmjdHytPSMGw6CV/NktDkzF+LyxRSl3LerRfrvQKZyFkN22naMflg
ME/PuHwQ8w3P0m3tnX8Tt+2o5jaYEblHIBSknjbf+0fJJRUT9pGLN4pzKb6b5e2b
nzn94kACXXCCjQVJVzhZQnpbBQYvbOjjnhrFovCsnrvMgpTxs1Vt2mzMPOwoaARH
S7apTC/ofOQJ6n42QHfVlVKb4VhnuNOVVldNFQLdoyttKknvZ85omizZRYxxVhWZ
DwiW+UT1cv0jisYOo5/P4MpsFlHHzv5133b3tf/kzQHApV+bsK7xZ8OoYHGOoXyT
+CSM1iEgXydHORj4swPUqAVqcMhMzTcKW5yCP4HCOFz10/j8Pojp4Q3a+iC5yhLi
rgM8twK2WQyn8dsXFw2NAWN5sop+awVWMCebRN6D64Vql5PP9Qzgv1gwfu70vRh9
NcLQQkCn6m5tZ9iQopCko+N1e+taJNtwf0eHlwb7q06HWobdcRsq+H+JjZcoXCvf
Hr7GFxnpLy4y82Tg+Crm6UK6rKoPU/73CIjlYU0pc6jqWFWn05LdSqqqmsR/79sX
dneDpZYbCko4udrrl9p3Ttfoa2S0Ghf1fEGObcET2S6YGdlP06YILn+TginGbksW
CX1ntBiwNrnbjSLGDjv9HHowJ1Ec92Q4f6Ph++pFDfU9oxNvrypyCyH+zKuo0FdP
m2LAqg9GhjYDLMyX/9gelSyykY/7WLAn9tReCBN5jxHeIlznw6+0id5YN5Qe894i
a440ETZxUWiWLL2VbU5mZNnqgC3eCX6QVwdyZNtlQsouXUZKaUuKC4gZ15vyktTU
Gkpjp09jI61FmL4x2m75leYap8XOzywfcvTpJdkTCdDUanRK3QLZLMovdqusU/7D
qy4YjlVkSh1YpqtpRH2MRK1uzxFpSUJKFJk+w84hV7AgDGeGjzv1x1Lyn8cRApyM
I7g1pP8ZVLoqkEGVYVA350iBo8F5tCjm91kjD5uUI+AcgVBVMYCEtqZuLhDI+0hW
2vU4ame6VIvmiaj33m+Xe+KrVXbRNH+i0Ef8WviaCgF/QG7JExmqX9ynd/3+U6s4
czX0Gg19bbUFIwTAb8AnwcML9IQMoSHE6qswcAtq6RXkiRnlIdTkXhlVEBCfV7va
ssx00ADztbJvuXSc9afoUx6qXZdBukN3lYAWEyzIMaWU1Pq4yuX+03xSOM8p4m/p
ZKFCNicXOWOpT9s8LvA4VVOoHSDhclMj5W57ND3YDsJujrL18SYnGopT/Duj7P5Q
4xhxWPg4hoQC1fn5dNUogKLFh/SM4sqlpHlDvrIt/zYGVjGewfRNWQTbl9ka6ePk
Qsb/rVQCYZ851SNu7dSh+IUUkvSSNfoXuD4IV9MxDjdhegacSytQRgIshfaI8jFe
4tmvGj1DbNNx7IZY1iL/UtHSdo0cPrwk6M84jKWpAC9ltjh8ncZTCfuF76u717Cp
i6M4YkUswKyjpeHihxbo0/I/vfL08xtrhOLGqOkN0TvvzM7QDt/d+fdUkZyL/JXa
3qaWMainwnnOBuE8K0FeoF+YqmrKPDd0YBZpjs0rEQV87hRUV+z46pprQ4jL/1jQ
T5ZcAYpP1clFKBVoY7NMHynuwY0tUQIMIxENrLqQ6cx8cLURB1g6AfoXIhkj1MGy
VK18lQLscyMYvO2ZOcYen608MSW8Sz/lQT84VLh+bJnR6dlkSJeOCFsgyn/++8ds
TTZWj4EKPezQSZCMtkA+wVlNW4hcZsrj5hpkgg+c1yCEcJW9mpClF1QVIiqkbpK8
7Od+5iCBFamXpr6KRKr16i3VvlM+YQTtQs6uGgXAMZgXkm5Ii6N6Rn8SA6bnedt+
kobIRd8barxJ2G7T1Ara25LGypl+Hd626z+i6keIrwsD/d5AtQonp4cQUBevBQms
IcoS+uBVohpFTgLFNprzSWyeJZW8k9FhEj/N9AnDiAgQfLWZMN04qm+jVQJnN5fm
38lWJl5nIPMg80h34AK98gkJ7kvpnLDQqiD/d3+xGjNDbDJCPqIuLDBB7Y+2wPZn
08CIo4bV+4ZWS9JPiXWikyjvqCIs3sHIFZAKjQ60lS6mYeoIqI65hUUOQQirEF4h
rDSbLiBfXo2ogcpi8XYbIaY9YIMIhBq2mQkEZnweI/qJQYybb5drOm+DdxHv7XNb
vGj3qNKIfOocch1zrskf2Dgji8qeb5HJx3ptO0HtO2qDlM7tr95Jpbny5Nq8sUbK
zO9VkUMb9jxVH+5Vnn2N4awQan1wSO7jWCBnoMUbek17jrjNVocxh+bSYFmqcB3e
gBMm1ipjPhWO2C4S0ztol7+h+hdgZd9w4nVMYp7z8vtNxgZytWbH5KJpJibahSLc
n2H7ZLpqZxHy+vooMcoAeOpE8rOnhXHNzYKj6wG/a+YSTg2ZwEiQRr+cK+XSQ6Pb
wg1eJ4EjoUrUkDeb4s12v4vloX/AOuBGQJmzETGZg+rsxlZIMhXu0S9AOPZUGrLj
B9Q1hDF1UsZ2WWqorP3DnehjE99SfZ4+7BDtKd01ybW7CDnN0NpO7nEu7NbcY5va
hYLfH0K8GEkoW97UQhfVPodC2n37YVYi9Ankz6nX+41k58ky+JrwLmK9rIIfEQBA
3WDAnaAbLOr6nwGIpRVObRJeFPHc1cSInZ1df5aozQsqGQUU2qObz+72YpDOjAOh
JwGN6ZuFts4+9OtYp1Uj+8QEIxXev+Ty/Ba++g6JtOiyiVi0tOYUPzQL9JOjW8Xt
yiOrouUAIL0AgUdDzNKHiaapqhfaaHvnBElYRPDRXkZvjYw+lY5F1Z5oFmstvank
dSZPU4n8JkHyyUMZIS3uTL/efqun/U0aFQiuTwIOcQwj7wLHV2cy4DqPCbLSxXHY
YsVxKHCPOuuPApaWJeLhC/rFam7yYu2DLE/rqivBT6w6zK8u1KFMfG7bCv8Cndom
7lJdFTL/TvWsEfisXnimp0KlbNxtF6+PM0DZPZ9veuJpDfp6nyoKCQu4WVffIOCk
eDOYslaB74Qf7vg8YYt5ro2qoftFBvEpSJJ0ZsvmDUNCQ98LrjBm4yoyRZmV+7WP
A2rQpx3LasN8rhRwQVU8TG+iqIu5MhYOYDN2D+JScZvrDwdv7NqvvIlVari4H2sh
yPkg9cDrpnS0DB9bE1aGkxneL1Ptfuuh0eth/rhQ5y7Lwh/O1lR9yKjZGuOFKhb5
PMbQEobmKXv0QdcGf0teye9by83QKhb5rwO7kda/P19EtiQMG5EUSU10XggxIiDG
9nUHR2FpDGdQamhJSHCEREkZ9HjGGcb+yoUKdeh7e7fuCRT643hDd6jTMXiG356g
Q1K7YqQlRqV5u5+nB7BUqFX0Ftq4f9ONJ+/NmI+IZvVwLgQprJsH6e33Jf4ZR+9f
H4uTSk9bMQzg/uqdMlf63u0o5bF4A7Nr8sgwMVTb7KJ2Oe80oaWVhh6TD2F5KBWf
4ZMK5jQsOIVbejN4TSHo+bE37FeJQSoj6HEVL0ewt+t+w9oeVjhXpdHxj+IaQ20H
sbb89Kc9DfAYca/h7//JpKi9JOfBgHI07X8iasp5V4aJT2DPDRivzWOtbtNZojeB
NzLZSU+yhn690Bmanb80YtjM/axdn1Tck9ICUxNtMC0wXNCXk2HN+iu5R8RCJyyG
oJVFvFlPgF6cpYxGLZWA8xl1bkaVLOqVKNdk4uz9LQJJKjTkM4eum6jdjDlo7LCn
iGsdLNCh9TqaCx7szW1v67mYlx3UetWvl5tLc6WnNzYiuG6BmZ0Wqq1DtBUR1e3G
O/WoWBrUN4ulWPbBx2uYr4/6sVEfvPbBfXePXu15W1c76FmdjC7NQfQtgLZRt+na
mcSneTQqLNMmsTZTcTLtu+iUfR6QEDEbIUWhLuIcaFuHztZZFHk5DS9Fx1xaPQGq
S4g6ZR2WDGShRInCDjnZgxTTqH1EIGnTFoKMpN1jFFmo9UsSBBfNQ65Tlw8rc0jI
OeWi3BF8jtghLnQWuh2irx57F3W2piumoIq/XibAH5wD/nvCrtrYEESrz1s5CU38
CzjSrIkmdGw6Y0UDz8/2bQwcSlah+4yI86CzrnRg/Tmb1EpHHPagReX/JsYb/izy
W97+JU5bw9GkPERj7ZLDIXTwCaCxBSxcqOYv+hUBTR9QCUN/pS3u8Ee5V8H8dq6E
+3Mmlf2sZYB0yPJ3IzaVdmE7OCuRrdBqO+FsWK/O1niatkEvZq7CvNvIgZCzFkqP
T6L4n6AgfVudiFF0NPgskMGElH1vx5udoWgGZgpga4nSh13P9BCq7OPGRwTJbXKu
f/ivLP5rQHZWy3TaTGdkmrClzj3O4vgp8b8+8LsSOcPKqbOJ/HCrmqq9loPpzmxr
qUBp7IOEAk4kM1uEJiWpeqRAtTXUO46g7GsmnqdqOQKwiwfRSFTFiEKSvT4csWJF
zDaWWKeEYvO1oPm9M4XQUSx1UUky9JX2/3m0cEHQISudXl7jzjZn4C136z4S2MYZ
bM0578iOyorjpSsgyvP/JQxyQDpKTj8c+cQNQv2XFTpT4SmL7yaqPcFo1SUpXNIP
5yQp5p738ttB/BkTQc2Ge19w/EGEGXL9GC2pmdCGgOwx/iIlJuTzi3hQ8u53Azlq
D5Wnj6ViCm3Gi7d5LSQHM0R8fMOL8c2+J0EtNU2hFhmvFfn2COjnKHn5Tf1XRL5w
IDaq5dp5SKNEeDh260EbB3Bf/TC+ejpZw37awwRLRPrTekvqsiMwsNE/TwHVV5v+
c4+E8ANHt3LFimuOh+KjCXLufBoJSE8cJLG+mpXsUYTLYVzHrKykhJ1Qmn8FBWhT
3loOe5k5DM0G1R0/iJF66IIyIuZ23Z0L0SDvedPrvZ2PJjWbb+dQ+vfWeP5ZK0GO
h1B/qVkMVTsS+EFSodJhxRZkhp9qBXCn9WtvzGeqZlVVMEVJLmsdY1YzQFjJbu+V
ljHAsC38EIgdMhEaMfhQljrp2X/61+4no6SIpRgjn3MS1ZtePPBnCV8ejJlf7R0v
F0TTwir4Sm6B3pV3RhwLN8vT+/38R/GUHS5T8AP4PKAWhn6BzNkb9DeeRb1+abE5
oIhas4+HJl5p7lHk8Om61yW4u0rXaPV9Y87ZkjWPqw3NJELJDLKZsR6geaKlyb8y
wvT/ujRhMH6rVL6IU9Hgc2nkhZKo/bazhry4c9jCpdoeWh7fliboLv9WobWQ2fCF
8KGvDuiMLFdZ3YWOPEckZVLO14uq5ROU8uVNPIsb3QcEKgIwWcdBm6wuSPF9+87O
RyakAD5cZN1zJwAWfjrKchwqz51Md6i4oStf65wawUNYZaq2WrgQsY4EFmHJDSvT
dBaXN7vA0qDMy8260K+Uhr2G6IOP6eRHXMFSZTCQtdj8NBh+pjA72tBbOB8mNn2w
z/RFB6KpBzyixE5Xdwzjl8hFMw6vYDOTk+LfL16eFg3aIABQJIpLhQnn2h1kg2H/
N0QzXjvhCLRAKwDFzlonzam3zh/9FIBAQc7lZ9aLVVgVGlvjSq+dSxjc94R3PV3O
2rUVdeiaI4j5x4DX0Ydqfr9rl0eSfBePEBj0JEDf7cseABslq6nI82WK76tTF8q4
EqlSVrrlAusHH8TEYYutNGSUCoAOlHZI34VTMxymCIobGyaB3VjNwP6PfaqwkdiX
0JiWIN4gTweG8HMgk/XXSx6xeTVbw5dNmVBLjwGEsnqocHEqd676ORexJFcjVJtx
buq6szYUXCSG9NDTj4FSXt5ORXCjjdYLg3tG43RtiLsvteJsds7LA4XPOHIb+SxD
aJalzlyb/WGHb2ylVocKToLKg1McjXjNCUxGmEtiMoEKfy+WjEcJMizUE/m1PpR6
7rgGlbX7lpZLcgnVJCRDp7MJf/pcPacjWUKYNtovySGY7VDJjKefSIyzKD1lp5WK
klO9hc28CYNOThcFQZpQwvrbJsRQRQKr2dugl8I4vqcyao/AC/cBVS7PhVOzxutd
HQBF2j+xLNmlpqKEUi0iQfCoPk4PS78qdVmwCnKkMi2I3rpgTrzUG5y2aSswGpgh
CDdM9jz+Y17kNqWJkmev83Yn1tcF7EDxSOFHU3uGopIQj+A4woZm+hALz0RGUmxO
p8GZI9x19FW8O468QpXD1TcEU49eHLBj1zAWMW2J/qLMC5j4pBWRjVDnj65Tt2vC
zqieP4/c2c9ffUj8AAU23VQ7n318B8p5H31XTLQ+f7PtZtCXh93o5GibcY5kGv4/
BMa10b26ohtA5mAM1ctOz2c8MX/yjLiRrlRi9HnPXZvIBG1sy8WVxIsgyQclWG2h
lFM9UzCRYHY0VEU/AhSeqSH888r9EGH46+QzlyRqH8Md3r2i39WE0Cq41d96r7yq
3XAC6NAzAgR1SnDpzVt36fkHPbhQw8N/GD/qBNpT0kdI2+l0rWHcYZZGyuDD5vKL
SmmXZodAHmr2g3g7bU7e77s3CXTcTB7ZCrx4gQgeqDejDyAQQutTVApaKxnHg7in
42AHR+LzFsd8x+8tYYGExciHIrM3Fj16h3kUGv2MdFmeYzFB64PGFHvMHCerRlvl
I+hXSN/D8lR3wZI8U/ygapGNAx0QGXy+JsFW/Qt5qR96uuHvhTo8TDMTzNlvCBbK
oXnC82xMrri/kcAkm0MO+7zPqG8lRTnb1xCGBSa76kWFNCJ8g90UEVJNY3YC18Kn
2VIcSH5UNqWjs7ThsveFwnXhhhNE9QdJWxsYsLa4TI0b4xr8Oi/G1c3D/lphG8O3
PqAleziXJjDOmfldeZxiSljw0azuxh1V1i6HdJZwb7by5ciivSKX28Yq/V3nVGPT
jPf2eRC4IUvINK2OFjadzYzGLhTB8OX7fXx9rwFa4YUchnpa9znlgFydSgxDsX+9
+G6ou3DP7aCygjeWK9YTnpFsvIcZigwc3CYJLq9wBVT6/GmhfSNu/cc+BZ6Txuxi
GFS1VBhhHemCHHRtMo4BfBC5rPYjnFcVYvn35kvwgrgJJehVVE15rA5dix5ObgB8
GaygCuXGfJu/UYxAUd7xUzqdn29OA7BSTznzYDNdQqec+AZ8sJgaxx156DJArB1a
Nq+SUlrNEodljoJk0dEoYGVaNhu7riiS75ElYJcuTxSmQfOmSkxlkRCCzqB8QmS3
VdzfN7KuQaqLcj+gWxkvidXv+Y9kxGrNVfGScFozZgXvLtQ2nZIZ6HUt3Ja29Chg
kIt0dEYVieiiSIuM5e7p16Z2flTwdvuk5cduc6T00bXQKtrEc5Il7ICj766KPwRz
Gv4CSJocdbwFRFEhBfNEu10oiClcg29Ib2YpJlOU30bq4L4hRNOrpwiXvkXXOwg8
L+5E2bo8aLeqQDAo362RFT8c/sRSl6b4lH2FT9KRSQfZL1bEAbp9yXlpWzE9CVLv
n5blWg7+7pYbDD9OujxsqaAF6VutHloIX1BBXm/8YD7jfuPSaRoraTRur/uWhXEx
jRrZWXpoZEPMuxvAYXVpsoYq+H53UB7CAF/mWENywvExIrlFzIrU0EImKPkjMNow
x9C8I7qr2CyGYHVTJxWB2/OLw9tNQBpemFtMA/ciH4+oETCz6WK7X8Ev+005Pm8/
73LghqaePwpetTTIluKcZwoQ4NUNZNiIWGhq+j7nK9cFaK5J4ORjGvnCXE96AD8z
iPLbyJ2T5blvy3Xt6gwPpjO7cKFizFMZMattMBycDFLcEewB7JwLY/NaeerjAdYl
QKcmBAYmT+FLLyqQ6a2ps9tVg/LBZzq0XWki2Nf5o13v68bulTy/AqMVoPmtg509
MuYiWZFuoe3p6lhZdD8gdeHCCRsstRp8+tUVUjmanFTRaEpE1nzD8XSnlyd4GG6+
TU4yJA6R+Po8cLwB2+SK7pQwEm6NQrIDQTSXIYeJWI0IL2TSIIMSZj9MhtO4Ont8
Rpu1Vy+IoSb2AJnk1uidK8+BZ5w6tEaiXVTETIexg3VlAIlr8uGZh210nWCJL8d4
ux/jKDettxDjks4lZ6OHsx4m5sDUODXl5X9+mcqwuiOQgWukmOrhYhBt3NCFqoxg
odkEsdQLh1DCDpIonvcZeNjURRz3RdR+IvQNEocbjLRfSeq2o7dhT7EwurWeigAO
N50prdyiuzIoaF+k5/vo47PeE++IUHsHRF0RBN1fs9AqLU8kYfipQ75CbANL/gfV
T9GM4Ky+oCsodUfxYfcBRi/RT+INxWKd0PXdpJsGjf6IQqvBF0/RG4cmsiUyuLAN
kxCq+qGUJxbZc0WEBd129PFG1z3sDLee7YSUa5PiFBQztttaZcmn1rg6QbC/I0Xk
bptKgNAGG5zH8K2YWkxdUivaAbpKRBzJJ6ejhc/cjjpqRP9ptcrt2A5tXOeeRfps
x6wcNIO0UkWvZPBKwQwxCsmazoTAGmhI5evqiMWx3QE1hLXvRWECqIYhTpoSNs45
nnKjZoPkkTTFVNlTomtTW83w74PdvWDvsSWRv1lqZMx1Deh3Scm04Jqnm3oSn26b
M2ZVmrl2eBBMfXcyAyJfHnFBj9dwIKP3EAKyqXYQ69B4QdHSXUEeuV+4jlL9PopU
E9ob2Mde6qIa5PXR5/mRu8WCpFrTE1wmZ2VZaDYXUQ21OVGNI51I9jDK5NWg2Hj3
TVki3SmjGxeLUYlaQoL0vg8Jv1GiRHRBzEjCQzFFx06rsD+RCLXLUOuQ+OCHI15x
L8mwyKX9vlYOIGmplKH8FBzoCt37wP2OFHdg+te1HWb9WUx9s8wLM9sysU/FhAxK
eleWYBkGJiiff3w9lREPUy+5vkr4DYRNsrCvUuLQ/nSLupkywRWklKfVaf+0YLv9
59zHIG/2ss0SV/hfjPTYy2LevjOdciD1LpfrsdBSma1vDsJWfM+HpJi0yPq5mMfh
/uZOHkosWuxcLlsbVMQxrMaPm83cH39+ASzzLO+imSk4hCSi0qmq4KwuTQ7pjE7n
ypmSwvLNQ4u/eFjnp/gRfs6GQ9umssttZS92UUpU7AqdIHZclY4lNy+BypSvEbNS
OAf/3YxzLm7JUBsa5TlzQwSY8n5UnEz1HZnfWWc6MizryLcppSEpP5eNHKlV3A/E
MN2VTc1CCKUTeWac33X0kuYXk762ZmSQ0Up6bJQNR5xJXhEJbh+cDhk6LhV9vntP
T0k2unGFneEcDQA4Qspq++73JH9ggnuS+ZvXgWGYIgEjobQtGzgr5SCqznWeHXr6
5qA4h/lYXQ3Rj3S5MV2/eK7NIWloTuFOWws6FBokG9NXi9WRa+twsXS9UwdePjj6
OY0AwYG4IR115Gt8lxRuzvxUScpHCmXj9H3SssdC789MNMXdM8IWqXaHjbTKwhy6
EAeD+W+mGaRZaj4RvnU+KZR385xHDaaidcrMV4yl03zU+wZElQUTdwoagPNgX+4r
YZiMBNm1njfvD7fw0P713Rn7AXYU6g4aPmLC3TAa3refnqsH9CAJyI8OJQ7MYajr
KMS9UAPddzL0AMaJGgorZU6nYHePOPge2sGJ6bbPT0HdGEkzoaGWJveWMnTIe2ru
v8jQ/5ZHFIkYDdsUovIeD6sk4GL5yMXmIPuhh1J7cVECom+8paBI6NLHFivr4lEK
OYi6xY53BQRlNc0trLBAtV4jdIYhSlGbYaQEToshteDL+tGiO/anSmpxk33umb9K
4SvpmL/DgrYKyyIKIiKy7YTNAS/lN+m1po/sW672cObbTIDlLSrwmQBQ1WV4Tifd
2+x9f2lgoOWKzZu0iGEgZGFwZ/0eK43fji+D17+KBXq3eZ6rafaLUYjo2SNZnHWu
jLjZ7+nLdq43BKCnwhqgUfzVfn1P8eTyyPqL2hikw+Wjyx39TltkxBQ4sGG87rr2
WuB8GjRB+jEz+gRyMKyieX5/CXsqn/Wv5SAnnGBnLuEpRe3AeihHBoZD4zyfUtSB
x/ojjB6icEYSwGJhFQzwPfVyAMTVD/r2GYN7vpj6pmNWTh2S5cKFHmuZtJJGUF4p
DRfIRXlz8zJ/+sBqemTkuywJAHDB2MC7negKWiMXkiCWHOgHgD5RLXt0PFnLQYR7
Qe/2oZ6jX5lEVV5PJ9Ms1ILXgzArgGA5hWC5sxcnpIg5UeyzNwrQk8Kv/eJE5+Rg
krymVTJzVek/rBZOgPsFqthyZ+lJxDijcvK1kB0uXGZdaYnzZS36rsab7L/dzzCS
n5XGAoU6n1cM0RZvtaAB6tcM+8LH1sVHVrMQcgsLmubHYn55E8yWPWEjgRTUplno
mnrpGBE1PeZNOY5LPZrUhtDX7GRgqxpG0oW2e/DnxBii7wn482B7IqKWfMs8dcIn
FXg+24+LFrTsTRuierPKC9FG3x5dYGLfBLQ3Fyzu5WeCt91Any7i6LosTm8h6Mrj
2krxpsFBs2Q2Q05WHqsI3dqgoRcQ/1VA/+1w8IfvMudO7riDsCnKDFiZ9mT2xBuy
ouJLUewhsS244DR++rb9vIhBXkQu/vSyAJB6Z70J3rMLtR6D8yAcUhUSir8cNLq5
HCfLGXAHkGZfRI78tZjTNHKEbdL/UH3TOqv312HMkpK7V8Zz/vIWnkbNEP8t9Eiz
vB+BgtqWGDGoMEfv2V0SUf7O6Y1IjRWbxOCiTw2Jq3we3+QAYgfSmOegRaatZdIG
oa1ux6W3xy9HQ2iqlgksX2VJYHbBDBpU/Z3mzXFfJ++psao1nylt36e8H4Kx828x
t+K9UeEqL3vsSfihmTVj59h1c/KidhsCz3UZ9D8Vttxx2heJoGhUioc8LDxIt9tE
OSaqOy6U+f/+0fm7fI9uQJYTHAdiIY6TMJFt8MIxemooS82hXeqPGlUPe4Yldu1/
gLYLzDbeCswHq94vtjcQZP42bv8hpNFmguNzEmrQ4fuNOG9cAPwF5KVYtXwxfyqf
dBRu40/rj6xef0m35tZqylW+cmYZd5N1smp9QdZ1xLL6jQSMKoiU4POrT+HXBGqu
S3hA86VPBDL4bxbar9GTImssSykslUuZ/p2jkk5Qd+w5b0kZE23IjyWDAKlhbXBi
oDFxz18xMB+e69IhrcbalH5jyCut99lwh1A8/thKZrBOULOPE+NlQAje3cl+JY9h
IVYwQPi3Am8fkjgkds2tYd9cHkcePd7qlwh0oezC8tN808jc5ugKNb/GlBS3H6De
yvUQLxMzLQZUawfSayd4RrBOJXpuUI6yNotO+Uzl8mcVzGYw1yY4Q/lRxI7gEQQ8
jgly5tPrhiFukcwfaV3pdV37gM2jo7/7nwF1mDgD+fIjhl9XJNn34T+kMvw9+exM
nsd2NWgg+zFRY71H3J1/Sn9440ejtl4IbEOzWBmvR1H2YNwANWpKYYeI8YCZ79FS
RNq2XlINPXM4MZwCDf9CBCJGmAtf/h/I1KRAak2QmRxryQkXpWwjvALRpFbemgVt
WqgQNB1MMHQ+Q9PEHUbPteChwHAV6kD5zamqXcTtfpQ3DzzJsnC+NWEYwJraRjdT
7Fi+tWZIyhyphPcrNiPVNsoggqmHMGs8R4uTcTRKSBQKA+YB7EPBlKGUGw+auMKg
ltf/tyjQn4T+Nq4RBvCWQvgymaLBweiloHwYzvaxiQBnnb/khH7kIGrjICzv7DRO
0Cw9FU6nFDcfUHIzF5gAfDSbOf7YT3e9o2WNE4IcX7dqxccDbA0FQ411uzE6bOW2
hxuh1zMtXqbEI1ys+eYIe+FQCW4F8s1wHd2zIlEafiFf0vrfwFjxaheP+ygnnlc4
OQUk/ZO+c2GCzFxecbbsTRbQt7mNxkc3KORvbrUCU7YyONIYGWguehsUl35b7hhN
3r2QYJg5jaG2q86pXK0hKTvIj8tVidna7FTkpmCuDTdlgmREDveiuGyHfwYn5GIj
ohc7Bap3eAluau6nWmIPv5Cl0bj4b2cRplV+5yiHInxnxmujrIhybf+QfuB6zV1x
lM1wSxZmxroWsAw/Fc6Pc+Dw64k9OGpeRSRPIdj0FbZcdexI70/DaZF+m1xaYVlB
dpS5hfUBVLwZ6R3gq/Q7rwTolC46kV3uavTuDysFrUZBh1IKto5dtRhY0+5S93RH
D/5izl5DB6UcjwTB/Htn2h2NSLmHKT/1TC+3hEFPaiTgHroimn2kOeid3irKb3G8
VthUmIc55VrAxnEY2wMYicri89PnP85t6rPxyv+KSMOrRK/Ogjke6Y5Yd2gB9CBk
l1CTUubMCmav+rHMs/ez4Oh3jvVxoNc7ZVq79eW3D8GRIBuTm+XlgVVTJHYvkQc9
gh+l+YmhwTLtg8e0BEOUsJjGJp8goLvkMhphGEZj7bWSpNRyTnstjHFy29aNYsN2
opDqr83u/sb+dNCGKT/A5Iam9YOXwaqCx0sRlnvjImSQtWE05UqqRDJ5q1x4Z6It
idCU8kXpyvuGUAP4yD7SNdjVh5vCIxRiAYMsYWP7Oeo1pHHWpaU9LiBsI8nvD8+7
aF1qQbXIG+LnVJcRcB73Q0EcUkraHvu1vYE3ePalOT6JhdFsHhFo8xkZ/cTrc0Er
mFOq4W4cqN8MdfX4OkE+rRLhBMewckA9cV21f5rEtdnUL6PX5KRWd0u6qT+biT/B
OQVAGdTtJq1+z5OnhJLDQuCwouwUZClidkC8LZjPNm34PZS98bf1K4t4CnVfw5Dw
ItXUKvxVBb11o9gUuuc4WteVCA9j96GgwzEwDNXT6VA9nNHnoiremSF6wIOhIh0q
cMMO1Ocgz5XKc5v+3vY+G8UmAT+9wZG0446cd5qadDeXiaXvnY4+nC/r/R+YwuVz
Cb/VDKcJWlXHGT0hCGOu1qOEE85Tk+BQNQFIaiPQWa8P7wOAIrxz1cR8zF/Fncl2
fv1YFdFSoWNL2/P+U1tPtootzLDkbKn/ICFH/u86BdA/MOmFH1hp9TEvSnicnmkP
8y1sBQkjw6fvtd9Ic6HqoFB2kB32Ae+SCMmn+wKX++qoZmkQoAXB6YEBJLGD6jOI
/xELlfrQGaQCJLiGlTWQrCsb4T1OiwRAyDNlrJg1quCZH1+n3G4dR0YO84c6ihnI
zJlnYJj47gmTaVl16qTfZ9K3D9ffmOWiYgD3yB1qkzrIou08sBy85ErpX+65SxPt
IzuumN+PrrvikXZqtJAcn5imF7COTJxstt9wrLeqqQUnRo4KgBmZg83B8foFWhn/
PPy2QJ6j++hAXVjvdWzfbXwPIW5tI+N6OGWcK0lJDfZuhVT0kyTSP4US8tnaZ7d0
QFN7wgrdbg82xbBmEHtc0nnfqO2Q8G3a6sKs2P8BDbfi2yywSlJUv/yBij6NK9Xj
WGeNKzFadiW59uuoaTsGotNDdaJG04Ou/JPP5WSwVf+CpVnzLaUGfc+86DXbQN8a
aoLu6U0ApAvJ9MofnHh8a7m4ngkOn798RrSaYkeu1LpUaHYOc7n62IDzLSNfTHvn
YFIafeQAhLFO5jVHCh23vdG2wSnq9eL5PBwL9eODN8p3TvUbFLgYgVpVSCxdoCb9
gsvx0S1hWk645xefTbGuz3ltQIa0DpSrGQAlyVrpo3sfJWSNtHZj1lEVnn3sSH+V
f0VCB/4JAOu9sopTB136J9YSkIbz6CS4m544GlDJ3LfXP7sd+bXafg6NcMU4KQjd
8jNiRaj1vN/QbKBlAdHzkC0rXRsOWv7UYcMtY0JMNqCZBQQ5nWL2ZMUwU2sU3BR/
QST/wQW76iyi0SVI/IHx9J+uwM216FDocczWI56d0FtaI2A2sFHK2qiQxifnlvVs
7CFXGzvJl22kE7NIQSK1qeq0b8iazHgPAGDimfD9oZ+cToIL7KOgipl1iAQD37fP
zuR9BMSRAtGsbZGVLItXogE/Bwq4+VjcJZCK4zNBm4oCQJ5iKkrOe9Jn60BthAjJ
uJKttap/BffXyiVyLcbF0WZl2GlgeKUVoNPXDMpYEmOi8mBwC1t7zrmY3tIDxGVc
d1REOS/wC/FH9U9BrhQ4ytpFbAa/8q3Rn9BftkYhrN7GCY0aHYiYFJQ/BrxCy4Ae
b+RrTHdilqKt5Y8rAmwJfI/pvZ6YHWST2B/+quQ9lhh6QyT8axnm0W48urgWBJQG
XL6kv+rQAJ6l7xVnm8bDKLBjYOpBMGNuvITqR6nj+e3EEiRLqWqhSYfmMTPQL2ZO
EV+/6TYtVLlEhXq0HkVxs79aiqBk3/JlFK1uVPjRaabaYQE1scDCrYoCKIR8pQuh
J1Fi+1RQhxsdDcvWd+F2yd+O7uUFUllfZ1WahWtTdZftTxEcn4/vF4IpoPVo9wQa
SGkM/OAYi5op3BlxtdbYIZY+iW+1PrKm9fVyCCOf7tFqIvrwDaojIdUWRxphcwWP
S364UBerDr8j1tnzlrdnyy0jpQUPOB4q0FlQGAAX0bZKvxwSITri00dTOrkN6O9z
9AkYtLRfz5osd3w4+HB43Pao//8yRCoVdJ2HvfRF26Ew9qIK3dI8HpoF1lEKh2m2
RHWICLGb7yXpyQx61RrUepiwIVF4hFAN0SWe7bEDGdVQFB1bba1DtG1812zjHn6n
FXNvd8Vs+WN733xfQHHozhlfUqgxky8jv7eG/gbtQjo+h804HgIrnHKjAIGa+NA1
j8L2sw9WDHiuw1iAJZlaDKbQjfwopV2Xkes9Ym2TuoC49oCQC8Nku+Jh0qqazjds
TIINz0YstbHaU2ErFsfeAow47b+gCy5K8mhqOldSOKaIYuRM7PGYVoUGPOwfGX/8
/w1jYUdukjBLUHgUo87P5V2sysJqXuGT4q7ixRLqPJEd8Sm6IgT0zFNlW65EKl8Q
Ff7HW4irWQDwyIrsHU0s25JpecZOhY1TNN9Ki0veUwTKjMysOOqYAQyMAYDajfkn
C3SrKcI8ozDTCXpbQCPKuCsTXIKmB5Ga5rcW4DWmj/bN0N4EblebOEHke5bwfecO
HaygfT/ucXxLI5UPT71AvKF+T/3gH7te5wRpExCjequ+Y7hilvV6k3HFN9Yem+3x
R8VEjo0TQhWX8v9h1yAFR/vgV1TlFMmsGvGE8VxJH8usAeA+Co1zQMrrrPBfusiw
70QdS3Y8rt400P7JrbIz4uHAz2sh98uBAHr2AXVY7UavE87Y5SlbtZr6dWo5Kl1w
kM9cYWTPC6BHnsFdTJaaxjmeH6Cmp6yj37eV6aZnRKyU5bV28on1Lw5YlHf3rSLU
Ti32hJUTMNPqd9RjGMXz96PQMgJQecQsTG3X4jR9tkMASiK/zy7d/AAwjPAR/0+D
Z3bp8vZQ9ME3w3PE1EMsH6Ic26hLSmNVju+c/sFIvsiiVWUGE47JUFtOhazkNZOw
MPe/ALAAk5D/iv3LLmKkpxc58H+6orEX1b1F6AAddc3K/p9pH0kvxI/A4pFVDzea
nrk+b75IYJ3tzg5a//PwIZCtTMRt4u1KPqo04BA1FAfD2Fy749CyDab1gIneehPn
l75A+KjX5Bve1yuX4nAXsyQPy9lWtZWH3XClXieTQH2IgFoLXRn7sIZcaLA8gKOc
BzvbXgk58C8gp5akpDMyRi0/O+q6BeDA7b9IXU1OmM7JpMvNG6EKJByrgL2m9xNq
irSc2iX+DUjYP3aegDkmjwTAfDY1j9frwiRmFmpiAaFMXlivBJgCO1jzdHc0bPmc
203wD37poGaokfKKPiNXFIJqdBnYk91h3im55hk3DgWmzBoAykDXcTmXabw18Qob
vC55sIY8nM1fTePgPglRYxcU91Dutjd7x81o8gBu0kxxmkS0CBf/Ss3NSvc5alXc
axIf2BHD5Xy/9dN9JGgUYAUlqjBOYGGZ8qLU5213AQmC4Gh8UYMpK0mr0Kq1mDzW
dw/9V/ju//9QFZdJPT8nO24pbH7L0UsS5cAH2d5vLAM74D/kyXeWF/4ws0X4Ouly
oe9nGVCbYyHDfbu3XowtgzWFa4SBfnpFH70iRvBb2xv02/wLAc/Np459ErC2DC8u
9vjpGHI5R7GsDNprRuaHabRaXUt2/PSI1h97fMa4yTIGR6nGmrvuAmkmGkKFfKBD
E08o+BU5FKeNP/01KONw2KmgLv4N2HCe7X3Jn59zOi8iSjyzlUS//eklMRvywn/a
95ifwAgqUihmo3n7cGd5RygNTZ1zC36H+bupJObvL6ndcLDXeNwFQKNJl3gjkJrs
bo3bCOcR2ugaSa1gtZppqQJaF+fD6/qM1AYNM6BrnjET506kPTQsaON4OCunARWv
4iNC+3zpzBANw9G8rg2Vx7TfdBaMB+t1sKwAorutZJ7Hi4tZpJRLVQLrtAWvFFXS
5m6WpylDfLPo7Rnmani7EaDXd/4+8BVL8xe1R6Drs0RMJr7kmdjH+JheRwwtk2v1
6NgFLOwjcb5zXRbcmKN6EmXEhVwrXHF+yHYD3T1bsTSd9Pq5d4cVksWi6/Z8WICZ
ofx3wpgU8t/TymuOaLwwW7leGrokLcQFlpECEUqxGn6wZCqaAhmIXmKJvxzYYK46
ASrHbcKPSy4R5b2HdDHIZNfk8vCzedZtgYXTr+EJxvZ+pPGOKXoZZOkvjJPKCl4k
1D9uCS95eruSAx+B0kOPws2gW1Oh2r7ImHwGqkbv3nG7G8mJz7ohMneNwc2yyiID
mfdGFFJZzyAPUjN6AwHEDy3INs+ZOguZaQ2RJmfUq0/6MhV4Zy9Fm3uvWMDONzJ8
6p0sq6/Lhv51Nt9BOBcyyKdgrcELrp4Dfe1HCop7CHXYklrhBq0c75CA6/uKeb3H
q6P7YGdAHcaPg/cs1OBbVy66eViwsKKcniA5PG8hYWVyBN8+FF95BXc73dyGnCEq
BdQJeyrfihiDaeN/bI1+E5FZjGFuO6ZiL02tUZL30FhKBorPvrGawoJCKjjfnQzX
RgrAaBfLKXT/IhdcfyCN2xgAT3bJ5FkHcYSHP7Ryw0VQi/JyVq1rqt0G6TudSKN+
+BF4sAVu2/7+TkYIpSmPzxKZPYs/FxFnJkPreFzh3p4/hUNy3+3rb7dH/Tdl2MOf
PkTXH0x/NDSWMrbxiJ2kJQUpEVJsKk0IOKoPzzObOYxkwcPPTWw+C2LnBuTSIzPA
QMUC3I45ARrRbRpHc2YeFMPnsqINg0V/br1ko5HvGaPuUFrVD0od1/nQxyKBf1cQ
6mnOh6hGEsysi1X90DSyzUOhwoh7B6bbZVfLUmS4MiB3BwEOuxqaOBEH0aa4JN+m
231QbqpQPtUK3dKtE4fg+g1Yol7EHU+K93O3qUhiKh9LNamzPMkkKbSty00qXyGW
fyaaw5xvIZIhh5O1G6XN6PgHKIJiaVmLRVVvRHzv9onkG5TCKokr/e8NlG5pm8VT
9vpBaT/CQccYDxmPBe9us2sE286NOJBUFil6DdQUJodAbSao/fZP3MWhAIDrNLS0
q863Vl4THhJG6wNa4XcsMV+BXTvde5JbmNt1VLZUHGSkFZoYqNFPZjurRg0UF1uk
qHXQFglxAsHoWFcSbc9Ee4VHKv+JxRpOQAjhN4gsPrp24vBCZ6izAUGBRa8/3z6w
grQdKh56pSFbOOD+dhbNfQoP9SogP3k/YoGmC+Wack2ilCM7HPfCYvtT3jiupwm1
hhwkH8JGqDVobf6brsxmbJ0CG6ha1geamgQUucZsyapNHh/3XZXttco+z9qCI0Yv
BhMfOcEbWT5zvyg3Ctd5KK7uCBCRWCd8WAhhjAv1PT2UsBOi3xKbWwMsNBVN2flT
Fbn2gzt+Hd/mreftk2E5fnrSr8gJ6vg5+yqaLh2PaSkukG5A0tknI33i4/Q+l3kk
KOWrJL5Fy3vUcaEHSpvIk9keZ1aa9phKiyg4IWjTYf52ZHHIdL4vbJcvb2fyP/ao
8n4KubEES0LESyBR8XThIVGRxTxwofSQjxe7m5rMnjfY5QeF09kguyNCTbNo5wGw
6wgufP9XNTuk4vL7VDzcnMvIYoC3Ka4CQW5NUUGGTTawxGvdLfvS786GjTFp/4If
kk7umNub51qdw9zDhN+8xAWbPHgIPENuwnqRbSF2jZ2NLLy47v1W3GRZqw3Lfvda
TqGLHKJ9jism6Yrv+8PIKs9v8WqJMvaw57ynn+Br6Qdn6qzhC7ecgP05PBXRpjXK
8vhDJXF9dMPBsCV1/PDYOb4/anao7VDFHOUalmKa4dhjFAwFFedDdbaQE4hvIKe+
XoHfM6doHD7p0kpfau1CuWAnEVrGslUnnvOXjKFZzLy2eMY9nNlwn38TQxYayP8e
4ypkvQ4DUTz32ZaGuFXq7cb3jTSPry7ja6732r1bmIcwzSiApKJ7qr8c0YHr1JdA
OSjmfIA35PaB4AG9+6kypfCYJNdz4BBUmKrlVOhrXZz7PB/bdvqXCYSw1BUWandk
LncEF7fu7j1+4hDAuqaiBnex+tJUzx/yrW1utvNBrzZ/dZSct6Rr+FNausbqvU0S
NYFgHFxUuSbSmrnVSkSN/s1rnXT7KkVx2Sl9OIZJ3sNceoqlSm5ZbZbwMhlMGF+m
9PX59SZ6BOl2cYMd6e8YRQpiYypN9xiMArUdPkX0AKpoWEUGR+0Sh/09O2b4e5zK
ABoBSRu5kKYxUiruYRVJrFtMN86R3oo8wy24xipPYxwt8leWcudoRndlf9lMpVOd
0dsJkWnSFK7z4sxd5ZNCoHH6W6apeVfrDBgve5q9mztzTTqrk3BvDCG0fn0dWw7j
nyq3P0hNVw3Dr7PTUAgFdFkzgzAuUvEFJNHEO3hsYBJynJRrtolHO2lsjki4UMtU
T0PhftAZ4oaV2yxupmT2DwCBBhYBVsWadTsg0wZWJ2N+InA2yXfr+HTjkNayh30q
vHDVd9Fz6SUn7F4QoE/7aeB13YYFcYhc71VRfsRCdUjhFLx1gqJrdGCCKP0xazOG
FeN0e3WPiyphERtcPtqfkLvfJrDDgQDsgklqHnFNnK+eluTmgLLhpoL0zunz4r0t
/5wK6bsaOvTKR3ZHLVvXcKFCKfGmGjvaZJhY+f5uENnG/xAkgxc/7B0wSzrbmLGK
USr9QCPrE6v++0ErN1LVN54AIGnroX4MLn7lf8jK6C3U6GRmObAZiCp7CO+OhsGS
hXAL8z67tzHe+O5H6ahSJZXwwdjZQ4UYRHZDuMXrpaQ/3Y997ak778kqcwEmQsSr
ByyqYJQV5ZX9jXzJT0frFjudm0BcmXaQoHciuUFpgMmTr0TAHF7LyvxLpmh6ikyK
96z66Rv6JNCFDLVqW9WYvU/gWPgPTZKaWT3DOTEOOPXBRE4Oc5EEtiGeDe+z/Xcx
/waB7j3aqCoiwAwQlCH/RPpyYOqiAbyBWGE88EJlPb0jWa7dI/QZxnVTd9tExlNP
UmDffIEtwXCxySg+imnKZAnO/rs9Vqf4drE3OehB7DZMluNqOsLr7awcVBEvYBZV
/74loRxN8l+0qQTk2QoQy287xQis/3a/CX9arGvrgxV9/n8CWGBtqmvXfRz1Lmxw
CejcsmBp6DPjz5aKNGbyrJmCX5AOpTXx+WAfkjGKdOtF0NGkw79O8mtY/U3TybAU
LjmPWfU7y98nJfQQku1WDHqy6Ku5+ee7i9W7c19kxEIbvyo9Ke7nXKhobqtaOxP2
HkzpwRQsicqCkFBbV+zLY67rYqeVe+lPxZwdUtqhcUcqHjAVfj/5Bn9h8Ny66X16
ZIcI3nqRUWjP7V1Lkmw1J6c+InZ5+sYTFyEYV0VmBOIQP6/g5eemiiG7TMtKiDU5
BUQjJncGMIDhyUvDcMgXgcYlgwlSerYG3p8F/8dB/VWBEqtNcjaDAf8nxZh2F+SF
DQotxJvZB3loz8bQq1e7XuiMFwIB0onTGad4e0vWd3rqCeTPRaBX8EFgag/H39D5
GYrBhzEDB17uaxl+Aj42VuE/PPCNiFgcc1Dg0Z07OOp4VdhAAal8NRoQBzjc30F9
NJ9S9GrOGmtyFBVG8sx4uUbqqpLVMic5R0/liho92YNtGzbeN8U2hwJAGjgwr1yB
Y1IF8ndqp7/PzqIbcheX147wnUO69cbLWYoXVkIHr1TTHRKBDoBxu3gx/fmdt+VG
v6Bm45J535LYVQMS7W60oovPJ6AF59arow8boTl/oqGgV1bbMEDNclTt1CbZJ6uQ
L5d+d2DHcdrlHSCbHSRAVsqrHg5lfkrbEnsbkrvNRsJs5bDm68At7FbFbNhjrucb
vGPh4yG9Q/EtKZlG+Lq8hhknMyyOfdJoaQNoRA965N2qpw69Zp6O+nmeGNnV0FMa
PGb++M0c9GYgAJrV+LMJqPaLDkJdxNX4PO71C9Bwp2gWvGw7bQpoofkFY/v6/OkS
bBguiE1sX/pfnlcZZw+y+nqT/QOW/lzeDxL8JRi93zqTYBAakxat9RYG8iWNFi44
5Se78X/if973r/YZxRm3jeMUT5Z3QFxLXAawOWWJOv1XoY3i/avy+pWjcmksUI96
qatBBXrvIS67EDqLUM8x1VlGWH+lHhQlmfM81frKAmUNLZAaJ77FaDDNGMnwywHR
Zm4B4T7kGV6PGp5L+CzPrKDvJkvQ25cS9oexdQGKtD8QV9JB0CiZIuVYHM2JnllM
PvJyOKuBp2U7ouiVBv4V08/y9EB5vYkiO6+8+q3qttzQzt7rRmBBkQzceWt2kF/L
PEQCUTwikS/+8itbt19uT/1JqnNK6JpzxpYBA2/2a9VBBUNcNdcUUasz/DfUpdEd
UPI+kof+/w8e8NKfswd0jwDJgD8DRAgqVBtwF4OuDN/EZ/elobN5JT0/Z6TQJDCE
AXei4ubYKzQHM7fURQt3RfgZwrWXdcjx2c0mhRHxAyJSF4T/MVFL737Nh47dQgQ8
3GKzJhnHLthSgZDZvTseiZN1u9+XMEbgrLUMuCKTkTLLnDGE14NiQCtL/R1jEqhJ
jmVKgq/ugl0Hy0/HdE+BL3brSD5gNk6JITj9W6r70rmWVFG8wtXrm73whLg/gMkB
uXdDBJinQdUozyrtaj3ekZ5FwR0Yist7foE49L1jvbG7MMNTYUBLbhxsU+gEv5Zt
MNoONUhpc2Uy3dR2iDRE8OYfOWI3ORL56k3IJH/ehz2AkLSF1cTNFb/9pH0Qc9My
Sj1ZMfjnGYKyheez7PyX/ChnA1KZSKcArsjnU/cxDv5VvjFq7S/gNrcylLVcrUFQ
PRkyY+bXjm5XFLHL1u7ndlqiPvvZyy8aIiyMiB4iJhc8ysSAUqrANPcvOfYJDN1Z
+LFGbLA8PEo+TiVJQNnhTg6GWVEn/2Ez7bI0JUaTfVacRvWkcqG3VPB0+8z5h7xR
sKX60tz0n2ZgaFhAfRnj5IcN+H1wiU0VWMvNsuaGPufzJHmBiBq8PGTu7rvqR13M
Z0g8lahYJUJnuh4rSMpTMSsBdon5O2mtb42jYAWIQuXFKv3iMSfqPwCJ4MJRHTH+
PB5GGH1iCCLOus3cLLnYuSROPoOoBoV1Gz5GVGzWz/p+vTXChYiUa3K6tCRw9SH2
oKsYDvoHxlVxXy6Alw9jnqbRTGmi38S/WZ6Xr05/oj8yE9A6qiGsXIz4Bezd3PYE
e6QBuP2wFzZTA4TiK5xhgkcTgrUhTHnEozt554Oht9lxdCj7bKKL3xo9YI2GBwpy
2dbsz2h4Y1kuH4KE7YBSQz+Mx+MvcL97Vg5T5TD6QTfP7LTXLUHocZFLxHFjpUTa
yh3SlhTYe9ytlDxmUd4pSIjHrRR6qgO2/c6ZMzMvEoymu/AEAroQevp+OXmhOoP1
kd3DuI5ENi8tdAvG3TftxfXKrqI/TRQfNefWqrwVrWtnMRGLDlEYtQTBVF+YCUrU
yyPTKljFH37YbtHKBF3aWVzSHWyj71dFbK3hcKmW4mWd5azEyLXfLhF3YAtyzYiC
HCJhiNU4zzTPSqit/92DojA7MJwwut/xuZrt0rx8t7tS7njfYVBo9W2gUV0n1Qnh
o2dLtrbmDA1rHKPjoQFG1Cd26IBwttRpDthK3swxRHEVYGLkzFFF5gVEW72MDQNK
fL9lIvI880zt/30E3S0R2U9iiNq0R8bl0j1ofMZ+MWvcfSTMisxEvdV96d7nNpT3
aoLYQ0s/f+mahRkPer5ryaQnaBWKaVd3v5Fvcw9VXBJJ+f3c+Bt0AhuCn+DJcOlw
OzXmhq/ycESwXvo4EbMMp6J91q0q7ifhkbXRx1XIWRIbqozWHDxIBFopsGDRPD0k
QEAiWLgNPbiqSE1kj7YAZ8vP2YRE8KdiEyMqMUbrHl6YgEjAYWH5I7/ZeV4uuIcq
QhwLM0I711FFE3+TFk41l5s59Tx0ue2rj11bBT3MRYZYj/E5nBEXBdZGNGbmP4hd
yHAu1AyAWZgvmJSjXEAd1Tb8dVZhw33FGWkR3sK9BzkD4wMQu8OjY1fK/nV99wJW
cfVRpUoIvPTXzW8X7im8+RGfnm6eFuXoXI3tuZnCA874vCnE/yfiOfADWuR7pRd7
9pJDhuo32Cciyma6m9O+xzDGpNhyyQMQPoItBpiXkYETEwThw1PZpnP5TKe0evLW
QBusXL2hgQwdgkbKfZI8dRe34h1DwShqXCgst0WIUUHJzselGn3PYOL04Kf9RkSV
4G39IxLzf7uhhSyMTOhKKhGPYioOrPHpQhZQxjlXFHKqDabkoosBPiCFNaXGsnDK
vkTpC4Mcb9Ldn9RVslRbEEC+Ws3FFvW9bxdEEcBiNX+NoWtqZmyzug2arLEOngo3
4M7C3zW3ptgZA5LUoFbihqspTB6hYTJ+cuuiEpuYOsgiUdwUcbv1rXyeIZooidrH
orJxxD5ly814CmHzqc679y3oIDILj5N1stolChZ05/zO0wsbP8QtgHdXByk0cRUZ
1sVITHVbW3xJgG8lxTVXFiTHoBG7KlIy++zDtKUxAvlRTLnMNL2/PrFVV1+zZ4Ww
ZZNCVSVB+Bz40zbsKXpkD5csXxmALeQlMo1+Xr29PWUH2SQT93S5eLe8u8eGFJ2a
YFEhlV162/KO1FsMfAq662n5FFf8a9naox5oW5B35wazXFOEv/rROit1uNji7/MD
EdNutMw0nRKc/qdpBNWeNfrzvsUATjtX5ed3+Jqv9gzsEGCqOXLVhkH0U8kG+HYH
xWD8ctM1QS26fnm4cALjC3PMVChrAMSitboHmiyrGIcGZI9/E6DmmZyyRCYhi+8e
Strnma6OH8LHyrbl154EpbQrlWOwjW0mekqO8JfMku4NAHLMxjjwY/weUnX1V79J
55p4Y727lrmW38kwK2V84gelwjIKbucSjbr33fVouePrRC4pGH5XIQ+KlfsaK86u
QnoJ++VBj7ddZHkn+ntwD+8FIQ/DrMPGayaOhrWMszKifCUWpjF00Dpkb4rSQyTJ
eDnbZqqqBbMMuvsevfOSSKx/xDHtq4yeE0YBGr6TMW6M5nljwIyjlr96tqAjSV/r
SuiQUedKgpm+4de82im1gts/tU4beJof6zNXLgfpAhqr+VaXOC2d1rPLlG+rHVQs
/oB4UxBRI0iKTatBpOEOjDH3z8gyVQCWsUzJuBelyFUKw3/EJOqgrQ9CpFimvLuZ
nB+ef+fvoIKG+TExusbrDVCgGkHZLyhxQ3UIl1kNlY/rbjI05C5Ar79tFDyTzlXf
mvEOj1NHBDi9F7/GS2BxBncSnnEUtqiF386f7Db+7G4lgoUdB9Q+pVrnwmT4Zcy/
RXOgE82ldy/p1qmkcaXIFnINGHVs4+nlAuWSMDkUvM5BulZnzU0yGY211FcAQDaH
9k4c8IB3nsZYdLfISsLm3/wrTQhBL1+rtA2rSJxQBINQVc3bKxRU2fUvGXltMUuC
OFddjLkTTAi89XNbSWm0gZaWJeuZy0XzxTa5LpmlAGfxkCYJ8J3s6G12rxz/XWRH
DBX7+LJlFvuaBG507IijSlzKOSa8+Nkk+rE9Xyc2g1t4BVPA/qv2cVjYJK0/XAGi
xOjqpSgWMmYQoXEOnd13g4bufciu/MgEVqZuXmuwquzdaVOlFzD3/R4TTSsQO9pm
I0LQwzi6JyEikiRLXgkWMZ/0me9DLRC4yoihhgtxxLpFnl2kmDebq8b2Kd8bDvDN
XAuz5F+u8NIP0QoPKMAvSLb8lwEjue+xXyUqrI/3dmBQt/aLNlmDSmVaAnTNgCxj
E7cKStHN6KeYCxIylxszBGYFQTy3cp+amk/BRFbV6KhT7hC8UPnmRg7nA+bSs+Z9
YFEJwm9ETKpLjLYsiNniZ/rtyYEOyssPdh0WnTHYB18t3hygMPi2zZRerXfTMF3R
VOA2Yckogtln2Cho56F5XBHwtSBj+IMQj+7QrJB5vcFe1MFZ+Ejh59VKBfEUVVeI
wf0fYSL3fE4CldCrIUXTPSKWR1H146hBWnMoeMI0MV9ejV0R6FyXXW+0BmxP6jvA
ZJ6WqAj2jjgFon7N6u0okU2kgG3qqvF+64F6ZVrUZ7lrdjwhuV4FgDpbycybtF6T
JDy6a3ufGtrxhE6yqB++KtmXLF/0zOxK/FBUX1jpjtKKtDFqcYhJiTvKtzpJqmrq
tEpj7gWBUdaNsI1qiSwDsaR1WrAluOZOeVPZSuMpL8RCrOC8ExuzsYW/zbA0DcNy
9wQ9UrcNKkDyN6eOimiXzDeuWs87r7BoX811U+WaPD0gmfOdMu1dghVioCWlr7WM
61hMpBVEC/wAvPy01B0qh7u6XeklkDuu2HAjQUiP9TagHLbJLxA9GUugY2t4qUbO
56mK+dinVDxcCDwu5E5dYwEVcdBRfIYilZxiv/pUpCEg4a+Sq+QuBHaWVNT42wTg
dNMuKZDWxjDfcHK13W1NB20BSZt3EQIKdr6oS2iB6D0YfoY0D+GMJGa01NklgXFa
5e/wGbQmP76iCX4e7smilAFJmjWSEiWksdOzVEQbwF5nLl/voPNJ/Y7jD+D/3c49
sEqNnrBe+gYNDfUL1aukSjZdoquuLWAD9SASWRM1D6OGJIqqh8JbjIaxw63NPMqC
SBQ9nBb+DDsOVFkMPY7Z1QLLwV+3ovsEY8Enf0O/zhwcAdFsmvhcAkZCTLu5OI8M
+QT45J/t3CaEfq2KSwZsEFc0/Eq0fl/YYkCv1KqtTb/wTKcWfNcjMI3ycXiqJQT5
OQSm25pl8Qye4+ZkVfMofUxGTiziy5D5WusEOR+636eYxTMsEqKoIEKoG5TcC0Ay
8CIJqGPS+0GIBEI7BOHAHTOEEGbagDhZNdQpq2aaCSTQ7bgZ8c2KIhK26WNjAZ+c
wrX9Wm8Cl4lzfnh1iSp0xL3sQRpU4oAA+XQqYc1yLuIr3Pp93Gu8S2xRBiJxUPs0
s1rvb9NgAAd/bTVD1gYuyLPM4SDDZSlL1mp2nMzAeHtBqpiitmugRWoH+prNA6ea
1GP2crbaRiqj1BWnqoJO46+fOJVRBXtwYN2F1CemtwZK9CqKIYvLbUiaxpn59TcE
DVDpqMnlj8JDk1NZtdc+ToX0sOXV8ugigC7HOpaxdI7nWHPyjX+NvJKnYorMSE4l
39E5C9ScYg084js44l+iYkTtdRW9HeTEyD3aIOVI3FAGtLsE8OXjel9IHYdQYzLu
QjTIm82uHXWFdqq1Ue7PF/iPdwW1udNPgEsw4CE6TfocDlMz5U8kzmkM+CGKHJH5
xIw1z41UxMRjAirgnrGDI4bwKgBADLWtQWly7AvNPaAoOIRBp45gIv/sA9HevYXE
Ys5JAVB7k3pnQHEbfLmh/vU/At+vv3K1E7rWAuPO6Wq621YGOs+CV8lrs1pF31/V
weTvsHfLxhkNxYihHM64cMIu15fmMS2b4JnVG5/hhJbArviw0SRSHiOCTcC6iM7v
3WyMGTeZ29DJrnsnt2JH/gkzF+Nf4+Bv3Z8Dsjf7H2M1UERPzpJrk+lU5mLzxa09
wWgzNLfM4riG06hQR5JCIhSBkCq8CLEAJEYtq5Y9sVEwnCRi9NWICVV/kUPBEBus
4P9c/vEjPfD6PtGjzSp89StvFAoEdOYW1bJgqmFlzrR5bGZ8+RNdnCmZEw6S5fmf
RGw/U/J7Qz1McgzAaJC0BjsCpbWdn4m53Qr1EzZL+EABCi9sDz39Afu8V4f/wVkh
FxhFcMpq3v4kCezI+5cKgpEuVxpLwKJ9wk/CgPOZDsX59aH57/NA1irlTF6LFqD/
aqcJWwr7Kq662HOVyKt2bMS2SBSZCVnJ2zqyWeCIEwiY7wrI6zsaOE0J1gpJzpmO
zEUtVn0DCiowlPjsjcrzncRjFwV3MYlUIV7s1iEM+M1sk9Fp/SNWVXV//2NRF3iy
mJ3Uq5I7Ee9i8iV+gZocNlS9dMMsknCVR08pntqmUlU+ECGTq4Jh+zbilo7kTxvq
hv5YfnpiAQndcrmM4OeRBtIlQkj0iKQDIikGrBjcxASI6HeZdagir5EyOVNPev6y
VCpq+i6qKYoIDRePubwy9+G9Z8TqTdp/7f4vhZ+RMse+jq/spHFM6vsc+FZZrs1M
9loJ+fzU2cd3WB0E6Pp9qjZR7UenK3spXGX4uYGCbxTQ5MbWwOjDnky41LB9F8Lz
/SrhwHJXbV8l5PzNFxP5hv1iOYMpBGuOL29MXlgKhIZ6ASF5luGXZDBmfGq3N+2u
mTAOrmNatHXQ9TNBWR7X3SGAfrT2CCm4nwx4WAC8Iiu1oCe3FBrhK4hblzUy65Kg
lO36lxIF3t1Ox+hQ9vD6naGrHmUzcgSgunOae2ZkK30kp4ChSSi+2nmD50G8ZKhR
YmTnWdVEVpmpKopR9cQWkin7buadg8S8FB0Y/9/T04RNegXnrsBr0glXCwQ+5HZU
FWMnGqQQASVJmWhWuTLReucdgrky8gOV601IPVn74U8CNnM9JWwelDBwdnIm58nA
SQlSJ18BEs0nFPV5fdpVxep0TIXz8nRkxpyP5kl2uxIANQnnC5HCsBLJv1DeD5Qa
iAQEGON+otNRJQ3j1Y12ivVgQRk2/14o6ToeS1t7x8RKvMCWvbMbgID8DvHzE6zU
PX/1VFuM3hi0quTgSoxNevPtMHkO4c+2mLoJhj7bS1hUJG7S8NIJC9trD8jpgDKO
kFn+AR/F1wu5SlTJGEKLHKDHaKUEi8+UMFN3EbGDuThj5RKJpzJAV4vrT3ZIo5Nv
VUo8QcW4u+fpFLVtnvuLIRFUs8OZe+lipNxIKnl/oKs/dJZ0wf1vSfWWumItxSwZ
CQ7UFNQnuLKgrZf6yaoD7Qs3kIID+BseQECTwlwhzrGUyOHQBZD6qBt8n64UPhRO
AGKBvOyhyXFJUWmGxxbR9O9t/58z6eMOfkQCoqdS+9ztTGIGxQ20paeJjIEkD9BW
m9RitPFAsUQsxUD8d64sAUMYDm2GIhpoydcPeNXz+QiN8ElqXIFXSgTf501cPaOd
476s3EW7p/zIFGlXi6gTyS4j+f/TYcXmTm+ye+0RyeKNvzYTNdbgMMc20WSint23
wttB7FdFmbHqo1pgdS63athfQfjRovb2AHkafJ5w88mJwm7RcfvSVSI13yrLHS6z
hdS/dvcCRmdEzMi8W8hBZmo8PVtyUw0h2U+2BNcHvHDPU8tug5TAIj+H+zXkFLPY
g9ocza/J8DLhKkSpnWlOLFcv0gbxEM+8Nm+9YIeNwVmFu9VjrtcqxChyi8gHP60p
3GHe+BpICdLbg/UnPEI/TGcTftwWPrQ8KdaHYsANIjxqmAPJNpAnnqoTTswG53GJ
a0JWPkAxtftxSKqgWuhzgbh9dT4j1WNK+VPkMWg2lDiyT0B1uqul0mDSOrq7oGiu
onNnOiGXGNMI/ZsFhNLj2xZX2GmpuEKqhbKoobQ3xr7thNtIeqNivvb7XeQeBSIY
0c5u47ZAddsaJJz41L8aPlTX4TdVwcZD1zkeQaFUDirIPSBQWKXUKyiG0ZEwjTxx
BbS5fA/MP2A5MmQB+9VgmosgfSX4wchF4MKQ3kKRmRgtYHWWMI4i9vlzr6a6S/Ae
rch6HgW1gFo6o+rEleywWYmn/SRjNR5WUIAtt4b8xYOg0DipF4iNQkNENIuVJCYF
VlTc6rjSVGgjnietnK+GQ8ZwzfxkTW0ilNragJIiuQBp/iihcSxyZ9uRCd/tObiZ
MaJAK/KSeRJAy3lrhwWJY040CQ9qFVhPQLheq3dktILn5aazpsnBqJgKSm/lRqo5
qBRGKekVQX7NSrXlBxStMEJN8NGDGCakWXT4ba5tv/UKrcc1xttWNQ337UflXpfO
+GcPMzL6tkxP2ROjZViUv/hiCjXhJruLFr5OuPuY+/yWRODUuj+m2Z0RZ+ZZ8YEZ
Piu1pvYanjuPX6q07cg6rHl3EMAQhsFhVKsCMBu0OrKJ2o24FRDHoCubr1UcagcD
TkFc3JAXdocyaJ3QklTK+DEit3HAyPaBl4bPzXgYCgKAP5zVOSffe3lHiBO5Qy13
SIwoO6uf5A0Fq1MymFq+5H6mmuym9mYqzCIaWmuQGRpL8gverTG2eXSVeK8ePUw1
ggFaIDh/H0H2r0Y3ANw2fDj3846FD31woYyl550olXVOreKNQQpNGY3qPfnafBwr
M+FMCTokyZozbmF+p65n/zZ+HkAQaa8MZrGOS63ifGh+viDyRBuFk+W0DPcOUlu8
NLbAF2AOvcSUxTxa3loRFYTO0DqZBXFjISRbSSoPHlmkdKZ/PbAiPSLR1T8gmvJj
LnFme/xiIaI/q4/CYVjWv+PfjmVmXmW+yBQXvFoNdKgjGjlGnMbyqOSNHUA8jmCj
9LwqBN/yHlL/aMlO7nQngGfrzaAKlNtiCXAj/6dINDXnBjJtA2LiaDkiMiTLbFqo
RKmr5Y89tyZIO0lXejgtP1xHEMaH6Hyx98ZLUjYFOuvF4511ZiKaEJCekKU6iPyT
b+V3udNQEbTf0f7rE2I7o6H7tKJd07k1VH1YC7wvlefP2tYT88C4aoQNMBzXaNtE
G6ySOkq8p98/Pp74/0AZj/fHvZuhkj1XeloT9x0yJih4aHMF9QhAkZhPXvzS9byn
YpHHrmKF5wj60IVVWqynsJD9wMmaBHlRybCwX4DGNjJRh9dz4P71t2/xymvr5030
YLBp6q2ymn9YkKQj+wKY3fVXvfJ16ILvk321nahMxpZGBlef765R1syIo/YbzzJA
J66tLDvp9wqnr+ABXhz9Zlky3qVMIpbQnWJ3MWOXU0ej6UBhfoi8JD6TWCLwXFaC
zQcO93EJMLskRJ6+8XvKYqQ0JCbXpjpfwvY9mqb+Kw82Sd844OX0EPeTfv1mA8gp
7mXPHRc/cbxdg+Q23xvO8McubyA3Xfm5gJDhM7pX4wgga/h//zz6ca8y7nuNLldN
TLrTzBW/7BAj2CE54M8PYEcodCxFXYPb4NMYtQgC11UxmlU6FadNXNhkV0rQyD++
VQx/k+kQmuS4fkdqqb/i9UI/3gz7dEr5xF4Vxhfo9wuSv3SVNMLaEp/aFQKlyaud
qmzCNsPUNLkHkHIWm7s9OhlwF4c4N0MyAAN9CxOcxyQbqFQ0O/5AS0OgJaIELYJh
53ei1Im6rLCzPPKbMR/SLXoReHweFC8u53JXylhFx477dzmc5RWRousPwDZZHqga
cI6wg2/Nf+rElUSQYRoD3zXPqy1VZkjgoGrF85m3kCcp8cyu7sM4r9/fg7TQLvz0
dqqhZlMq+j4tM40hHMUxvImHpDHKH3SPX0d5FJWehYYGeWEBEfw5nH9tPPRYMWdd
ZMdeAzwdmqx6TUHsQnJXKO/3DddL9ZYuVcds7qrDJ4qzSUK9oFNQYwUoXgQK8NXV
lPMVhAW2Re5XkUH3xLTWg9dexE0OCvjQMhH+p23t2BGW3ITc0S3vd4iZ6GsHP9wL
MteXkIVANLU3V8XkQDkF3NHIjNrZuwJdZtrqhHIiRxBGUj9S/vcuBzZbgFLH9zXs
UYtvaqDsELnubR1KoG/JqFrhB3P0xeKKSbT6EAGx09EbOU82Zh9RuSt29fV0yf9I
6CXyydBzYcpjxzBMivHZgB3e3eRYmJxBPCQ7BOig9HzHkP6t6WSP1EDuixx69AE7
I53gBMh01sjJGqWg//FDQiouGk1AxSYfahvkZcjKPDUF6uNx/jvvbMkG2a8yKoJI
/9fdjo+5d9ytmEu/ccao6ZT2Fx9vEos75oLGGJArV7PbkcPsjl882TGpk/yZIwFT
GYR/MD/GpReaVsf1s+bQ8DCWrnBPYUxe2VhLr1bvBreWqwhDpDG1B5tOCO3fd+RI
n3Js1jGRsNjmd2/w79WS7gDA+01blTtSAHE59QQWrvemEhmincL0kToVSRNK1Evl
oPeeXr2ixQGbDF8m0UdnOGciS8l9G3UjG7LcUtwj8O+mRDXnkyA4gdvvb2bnOLws
Tzfw/paOgkov7GCido7xARFA+gnKikU6p2cDTaDO42JzElPS5bZStq7DaBU27/AN
sX003b4N4WD2WhPLoMq+CPzsMt9nBzK0PdcyHLSBGgmt5pI1KjvJ2sUIwGyBRxFx
Rjb99eyUGZoUROVGmTJOdaiwkzCnTOdmYUgZGwwAilT7MNY+p5OLUDdT/wOaGete
K+4EmpLNvoggWWKr+EC5MCRxATmGCMRND4aY2KVDpCyels86E0+YNgNzHfUGYJVY
nkKizulBnXHbMLXOwtxE/U78EVtMiRArYEaxYgv7sINv4PtvkQkRpykmxmYf4NmT
XdwOwfroGyX9PPuGMWK+1W5E+L6Pl89Q3kK8SHslsKAzqphLeH5dwAKZK2qcthNx
poS4UkA3lSSg6knmvKrzc2gaLSea2CWwHq6Hf87DpqgbSvP1GK0Dik6/8cpl0oaP
uiNOmwaTTeLO+5e2DGeQxIex6FS1OYVxNs0Mjbq2E3MXa7EWTjOZUnHMCafPFfrx
NXvC3jUx1rEXKXU6cR7C24RwZcn9J4TGLuQrlP9Y958bFEndzPXnpTIA0bwyPYLn
aEbVQiOMJ59YDEspZ29cJPLIyKvnHxUafrjfuH7mUGXm9lOsmu+lxj/1uxqXldrB
WVIMRGvA1OD+pdcfjeXL0fxZrTz1Agg2kJt81TLWY06hbdlHrf2/BNaLrlpE5fON
AqCDksR4C3cOHZmZHe9MHu53COVKg5mA+nABLX2W/7/Ruw8t2NnHEarlhpAoszLl
dhlHio72h1dE7MixPPG+EZrcz34NPNgqZA87bL+hOMjTBP/zEli7GT/cLaNq4vrE
q7ti+vl4qecfdpxwSfKdFV0RWlRQ6wIVW89ELmDAkKT2ltqs2H8AHZXwSQOknGtx
QURSa5tU+w1Mn/lasQoN73rV6Y1/LQVVafv/4XKSrr5DhJYv0L7vd1oS/iq/M7hV
nqj0rftVzCFI4ppa3nsdnIrP8WlBU8ozhxJDC4HG6uJzgJly7tUATQdEPU3dJYKH
yl3ygFylCniM/4vLCXaHZ/tWPE1eBiJR3pgF6oHe9cM4dOY2QnhaQ2TzQZZG60uF
Mh72MJq7EXHGykC+ZY+uMOCzj7kE4yCddOqFsPiOvh1A6dvd5twBAOGnqdY7i1FM
QkPP23mIcfZJak+/b0wEa7GJ0Pz+h8Pri7/lPymqw/5kP0zA4yfM5ek/YNGZKV6t
ek7XlZgeLWSiKwTZLeuuoLxHgG050N07w0HHu83t7/CU9YNFGlHNivrWRmKg5lM3
R8hfUHlTONKdINDYhBgS8bbHu/gSlwrQe5gZEsYy9ccY/dEnLEXoNrGTDtwBSS0U
bxnuEFrXHRzZX9mpv7rBVegYDSMEkxz4bDT9Q7Lw29qO7b+unKinY/CK5Ik24FSf
KqmWRgbHMOARyRJNJpub3v8OdGEJ8dGPZpeTkRktAj6m8UORBkhw+la9d4sdkcWV
xLzulSf7WtyUSNCFsvXuBtTIVzlZXyPo/m/l26xm1Bqhy5R2HS+yrXZa6lpVknu9
+y2Ap+aOnAnR2t7D75BlaqSa1l8zrRt8JA2BuLZtZGRdQwkI0vmFa5xMs6hmPfcz
ByxXgfd04MOUc8dxfbkxunRpRSDqqCmAP0KPBtnft0VVkhv1jX+Y0hb1jDn3/3lJ
NR3Rebft/hs58Ddr/R2XKgoaUwhaD1ffNE2+RABbiKjVQuxU2BZexMILY1x18NEt
+3h4zYIrck6SfLFoVPw/GF2OC2rw3OPVaMo+Nx35OJZ6k6xxl7fUwfINBlz15eI3
McVJyvRh3ks0RtStINl+PAXTBujWnSnvtbcLTmi2JVHrmPBx/tUNOaIyeaNlnCe8
JPZEA/ncNkYJiaREiBrmD37NdrbQK31aMH0Oa7k3Ve5qK9Iv064e4iFr+AdvXcFy
9GlxmP+NRqzRdPSTKlduFap2dnfWdF/t/rR/aZ0aGPNWreBq7cfQeZwFMi5mJE49
+TAQ9iECHngiPbpYyPIVKSD5ijkl6x4xoX1LhjtnwAqHdXppfMJpmeCXJmKQah2C
kR/HaNF70iRRmn4KFTlKI9OToflxagsWvb4lzaXG9Js7WoaZB2h/2GUw1uWnJKj3
LL7bhokCgoz1m19yGJ5JHkBik7lLvGgrN6avXAugNIfD65SRFWy3WF+xOz/EhlWA
FlVb8/f1rT3ZOCzsWzc9loK85+ym+Jqzd0wqy2k0f7wcQ+6qj5dIqwJx7pxtJgRA
EHW03Hf5gX5wlh+sLsnw7nNqEzMxpHUQffW9hwIDKvg5mRDOofsnrclQ8T/WePlt
d2XKnn1Vm859aMb1kPRhwVbR56sjkF57gNjEEvkDtkRHzkzD2nOmW4iy/Msr/EBJ
dL4Kg6Z6A3IMsJlGnUF32ZRH6JjBgnsYaUdSWbn75/kJiSeTyt65aa7B+bQYxmAf
QjFYJr/YNHrpFHe24qSrePBhGbhxdPd0P3tgZMLCU+H2X/SgydBD702SmaH1g7Xz
HTCmayXk6vPzzQbRoePTzER8Is3pqYUN99NPLIdnDCSUz8WEGqtzraU+WbHiIWrt
ogcGG01MpoFxXrCkjatcSCoN9gnyCmuMtf4NfoMeNoebws7cAc1XhnyxM1H6UIgE
LQBGt1E0pB2x0v00/ueSGxdU58hajkMAnCQs7GaqVb8fZ5P/GfSZ0rAF3JCtbBUZ
2a3SeteUeXYHjaDt4zb2t8Dt11eooeknEFD4TrbCJD6h2fBsAUWJxUMlR+JIHcjD
ka75a9k1JrHguB56hmUuFBmRWdo6lDOREssbgwT+7GDnUtqdA8dd7L9jvsPhjY6R
2KDm17DeGNbxk9LFueWkuEQQKxxyd8tw/8/leQlP36vvKtjiua9riJsKA8Q+MpXB
2jY0cP7UU3WTJ/0WddQ27czXGilqFDWOyUh9h6kdamhJdQcyhVtxC8OBBR1jb4DV
EA1nnErclbPP4xn9pxxnCP+IL6jeCxiTJUEouxSIrNg14deWexD/CtMU37FESKp8
GCoWWd+He+fB2S0LLXTDd6wgQa9XcFVl16zZ8AZNfIeZ+nbB2pyqDr81B1AyHfLn
FD6KyD8YDS1yUE6hDlH5OWiZW0qexInRQG0ePoEnKjU2GfE0LKdN/xrk82Ldmcuy
M78GDDJrU+xtHX1GSLEZvqH0DO3l6N/m47wao7DevhbNrpxNaMyUIklKcmLSIR9O
Z7fVc40J50a5Z/ieqcUOhFUR4x33O+4eUFmonPQg4NqWpF6TtGiJwGGjlLkrZ+3o
0EhPbyFrW66gCpc2hsmkWGwmnedIItkVBcBoyxkOqScSYIFlb0Rd3/azYKYSoMsa
vh6hXsYrneU/Aov8gkl4iKWRmgSNpfEv6CgpsmEVV83tPqoPFztNPilT44oKXKbk
22WJ97hrNV6ixPPcyMKm8OZ+i/BhXeTZfECD9G6hH9jAjL0b9RAwGg4qIuOZFV+g
Dut/css+1nJlRnwZgxhEwOBMJgg+2gLTJA2mjzRS7XEeVR2KRnmegcgLUzT/LznU
AxiuozdiGINA4sn8IdDykZZdwN4b3ePj9ugJeE3ZdloB5XT5jqtzuY5XmsXl02nD
pBLWqA6PV2TmXtSaWzC+u8fBfEI7oeCuUu32IpGXeHf9HZSwSufReXPiIcv8fDDz
9UjQ8VSjxWxa1A7jdBe54BL0BankPPj0FaK+A5z44PKpWt8gyES3GtWZYyVVhcGh
Z7gjXPHvuv7/K+RVmgCNWuTCAnL6FKTowlOnC7gtGj2mZ5v9tYBc2yc6KgpRslNc
Ofwh+q22vcqp4U1e1xr25TMnPM/mSl5UKcVg4tyY3jVREFblfF+ypehgQuulofIJ
610SPESH58y+dBx1sjwZOGyFXMr3aHl4+9t4qbv+gTKCXWq36B27eUAWzsRODd2o
NX0mdVNjwvbIXqFwLJwCvmT7t7TvP0ZzZHA1f+/09Aeha18GGTOXShuaI9GUv2A7
tHdsrYwRdv+sXQIRio1u2KjVFvq5Y/FdBHoziH4+tipJPlsHc9MUtBBQNa54+5K0
gVh2g8FsyGb82PFNvDzkjp+kEMSr+GQhNOnzpI7FpeDCg2WHUMOSV/ROBApBNAvX
Vi52TUnWHt8pNt+IMMVPTglVtzgySPDNs/RYuzu+wG0bC9JtD7dzCzSXTGhxUjNg
IFko57KJGbbb231Cob+rHy3x9vC5CDXDChgiR8Sr3XFEeSVxNavtuhTED7GIiBxL
8tfMjBHHP1SHEZFUpBrL2wJFth3yEwl8SuJbGLz0ea1Eg0ymjj+9UE6ezI08tabp
vcDY5Bw/HgLrmdju7vXGMNvVUsNaP8kDbKuJvy6f8sep7K13xdm4vI+Gq62DUb0D
xn7RARvdmMFHQzTdmQP++gwWnPVEsDbBbkxvESPKdeYFeqUow++IRLPa//iZArmG
NIEQX2en0QKcjBqHYNLdSQ5fOQBKuKj64SViy6+CXN2L737V/32X8oiU2kgGL/4b
cKWz9au4O7LAxl8ZatfuLqDQyF9D9Lbjj4yIthE4DuxjO2axHmS9lCnTbrE9bPQs
JcS1/eBX76SkSsQxfG6E+Kn0lE/6xQs36NVli4uVGhCzcFcMES28+r0wHiUDtDCo
dmwd3XVrI5QT70qF778vFoFziszcc9MwAXYPsYtRQhi+Gcfm50n2mpvL7qBYJthu
SJVa1eByQfNO2ymb75kn6n8ShbM7BZpaa/ffz8NJODelDKlWAl6Ut0cpnLtJazcI
XpAKwG0xhGrfNLDXoYWeUVP36KyUx6hz+UXWIXIlZgNRikeLhugmgzHlhv6Otsyv
OFaRZVfulBvcc5Q6vEnCtTwThpqB3mlYJmZxPBk7wkAwDENsx2zPzBjPi2qEIdv+
dmcoNYSPw4ddErAKIFHy6gf0O+GMDD4r+Wkl20N2+SXptWmDSomr6k2gsde+iu8s
LVkoInipLTRN+UB099k8VpUrK/vhrO4CWClirnngIXyoCe2CGu5S7oFCNGNwcKZm
iJNq2vY/YvmnMZioauagDrILsCONIujmBkpNbecPbfRYnX4lvQI1coG7Wc9jrHFW
yhJ78RiFSPU3ke1olACDDhrnAGRiMLEV0mjvJeOvZk30oJ/OjPCVv97fJSBsiQmL
G+KORVjJ5sEE1yHtq3A4d6oRLv7HAe0x6sP9n74sNTTSdRrSpacghf3ti1vUPWes
cy4xVTRlMV5ROYWtF+fVsxwDIxKPez+eh09m8bmmatfnRrlsH2uy+6QXcQjc9ylb
VkrD4AOgGcfZwDN2iDwVhJjPlggL/kcUa/lowEMzzubBAhdjpS7lNeyllZ44N5a7
tzkOmsI+ZMOas51boVYWI3fb3stIHHkNZmzinDum4blltU/FtvnufZnVutJOMauk
lubJPp3C6rYogNSIx0yVys0mlzh6Xbdunz7pDJ9+lFujUiE7MHk415SrYmuK2ALg
5/gTkaG4u5aEXF5wVqvU+o9e2tiGrtt1SUVcV9gEcQyozfx552VdLlSe0jypbrrS
ugtRrQHKiBiz+6ZbWLhfydDwaCOb93QZxTZYMOPx6cbpofQG6ZwBmibCRrsJMgC0
fpiQcPBxNd03f3Wrf1rrxu9Jh2yCStiDf/iXgkDEc2cXY7gDkYbwANvWh+urlRwp
+7UE4In+CfEaNF9i3HE8YqPR6WybOjuHHVxyKwAAI7isFV9zvOyFqTbQjwhNe61N
shPZLLa0joli1SBjx9P2S3PvS4bj3TQf5UFRgKS7iORkj3zu+HLHVwK10/Zup7MF
oLHvVI02c/v6AdI8abHfNoYJpglBDks+gLMkgTnJwGjm0iT+VS8dzVohwaAzbgrb
UYjPYSrRQdIXK3NbWSvSh5pBGx5UrEGoCItkiQFPji1qmeKA0ZcOGWVw1InP2frh
KyNJ7n3A8EdWCIxOmya8LsAZdE3yCCLiMPY9EurKVVRiOFacU/Sa21IPE5flyfoh
z1qpRnrl4QRfi9XuVjbW2+xsqEG3Jf9hIM4+6Wn35+Rf3PjKIcHQLceYIFjsTViB
zaYuAD17upI8wPgiU6l5cnRZawNw/gUEV34YqSdG+QB5h7aB2hsyYpbnxzj1YfLB
Y6AP6hhwLYTVMGawnj/OxqnNr1gun0qynuDygTqhnXUIGZI3x3uAwXKFqBCqI1Xl
cIyHoBGO+kT2ha8ipOeujTvzhaow4Bpon+RtvtM7fY/MkOCbN9oqj/S9hTVIplXI
0f0uxGsQdVj4ZFxJUnHSZSfBlMEPjhl5E0Dq6Aq31cy5yat7HG8hqvALtRYEhxZk
YGHRGOFTAOVojTjgrQnYoa6fm0gJ0kYB5qTOnAPujksQtTT4tlN9M2c9YaxqeNL0
RHwopbeWZ57u6bJ6BjZ8uY8w0BnXzLfu+pTymU1yK1qBAPiMew94eIb73W5md9sM
8GGrQpdvfjgArFM5PEAgR3M3+7geHNsHVxsQdwSQt8Lxt530jfWHUDsRNSZ3QJON
3wwOAVNeCKvTuJu7rD82kNbFEVnw+NKSqD0Rd8RC4DdRRNTzZrc+0lfBNZqM782d
RNvIwUH/JLEu8R+T+Vo+geb1hJSqrg2Jr5d0g1AMMZnT4DWeSwOXPDTNWQzoV0ga
MSqQI8XIxdfioDzD78UTSeqBdego4WrUDNIUGYQTFwVKJxGSt8dU7nPmIFXwDVO8
CTnq+n2ie3hcmvkOa995/7NyQ1KFGryAt4vZhPYAVYthayOSwJ0nN1xAX0yl8wr0
Y5e1FjU9M9ktAbUtZb1fvDWm3zoWhDYD9bgs6WOWimQlXsA72enR+K6TgZNRnS9l
rYuHkEBk8+ZQQ3G79VetGEVA38+LfoM7Bs/kkkU6XukgUhvFjQqMf5XYF8VacLxD
mLUnOunxfUl1RZksMQj7iue57Fr2t+1jZ5yG1qYF0bGu6XorF2QtrumFGVUfd6Tu
knbZUHeVLheqf+y0OMgaVZzssU3BQG9KdqX1/hQC36Xkpby43aur2LRQ01es+8ot
ckepvxN3AEVwaueOm+Zydr86cRO62BE6uZzC5LfZGBgIWu+KpzIuKjYVvkTLNXI2
/3GbxJGJoB4FxSZdtL5wpF5Fw/eiSQD6XzSGpII3gJEKiPc03yTXemFTevjrrTKi
y8bhNIvV1uNtG1LLfyo6TvELI8aiUeUjrNfUhb0RJjV3hFy9ZfQ8SnzAnV6mZrsW
5Io8tMWKhhpTh3JbJQkkJPp70LFz5j3Se0KECUKG/SSVNTPjNduKFaI6KJgRp+US
icO+s786bo3xjS2ej553Se2I0toEMfAFf/Mv+qXiHkoN+4TVYKsWznmRVNM/oyej
n4EgV54GgaC+R9z/5FkghSFMxNl5V9G65FXsfSZL5qdrjsXisWqn99Rf8PDvNsjD
ZbyBiXJmiwFcJGBjU/fbTq0lBe1uO67OjweYqkcO61II16/8CHr9lQxERezcW8TD
aWOu+cqLmMO8kctG+rDklOY1AFrA92jAuSxqx377VSMCXs5PQ8FVzp99swLvA2So
ZrEZPUIibtvkzoDwzW8510Y07fb4Re6DL+nQf9KxHnFrKbw8F8NN5MNLrEcjQXYa
HZe8bE0QX7aeSM2wSy2Wjsfp4Q2+W9RBajR49CkpcWq8OH4qwRsImxvlFm3Z27C2
hsKgTFbJAmJQVdYJLfq6K1xE57SoZERnwS7rU1mD1+3uxol+Wy3UOF0S9N/dm3i9
U7duplYnluRffoLERaHUA1ZkuBYnK+haKj/iVrgLgPHzjDYEaWZMS8t6tQQdknDo
/8WIdtH1zjzUXNiVd+XYT+j01pfzsoIXDK/W4kCvlP7+faQpvA7/PaqZA8uG3UlZ
C+4LWa+PiX002tsyek9d+Jpx0QLHDhaMGL3AXxz3rIp4W0lngdtG7IyLS44CI/LK
EmappBXw3bKwkgpFsg4zDxHk3cuFo+LlKGZgNBsE6arEMgJuSKBi71e3vHjxs+oM
N/ZX16IcALckIPnpEDtGwD4vfjVDzKcoGSX98uIHNMlnEP9UqJIQcexCBWKOV6/n
G+CBmujzVav3XbQFaYicmT8pS2srq8zt24yIVpRP7nGj/tNMaex6Nv+F3rrB5FfJ
YLnQorxqbHyxuVPU87TpPF1vFbbMPqvJNwmYL05PD1B+jpT9ZThHyQk52tRNZpTO
S+qYxmYigstWYGjZAE5191HwU6BS1oUthjRXQguP7FiYhFh7HDNZ4pOCB7UqvnBT
w14fBEUPh6visAcFyf7yp7RvDDL6APjmaYXRU01onKnW49cVrIhrFgEvQw3cGQTN
51I21UBfPh2bWjdhJyEmwPcqRfTctL1w3kkQbDkSruY/zTLcvZFVYaPeyj7Yuzma
E8QWyqVf0KmfgFYiG0dcWv5xaKa2uArbzqF3YbgSd0yreAHEq4WU17gFDJAZxeRx
leilu33FjLImtfCEjLNMkMKH88/It3TtLPIdwDJKXq1P+mEeH/x+jvkq83yrIPy6
ofDh8XjPoUCYJ+Ka9Re2qNzr7nYvqfIgoG7JOfw1C8lxRxDMpP+N3bVZki4HVlgv
UynAmGOpcjoxkORNWjUgXQj2dUYBVDiOSUNkY/G61YUSTEqPVD7punv8vw1uQsel
PungaU7i9SiXx6EGsN2myVhxxwiGKSAKoQMZGsqHlLuyNFxeHbikuXsEAU0nAKcB
wfmTqqSHQtfUWALz4vebSgXL5RUDE7hrkEpBQKv+FFJvmJ+igZFe1i2tDGOISMEr
i1kyeDo251mq2vuhQZRiIk7x2n2Uj6Q4EBrU7dmBEoWbZLKpXYLgNR7tDWTZCuFq
2wr8vTAs2qO3O2mSpVHw+YkMNNCqxQUkzws+FRtX8MYn91uL171IBQnAi10LKniC
rDGBxWDJNVaq5zl0avUJ2/gJ+12+lJk6xHBVbnZABuXJCwqAfSFSYqCWC9RnjWI6
KpMyKYopJrIKupBOsyV0FTj2qs7e8Dx2rawBdoSsqZjhCX3Au52alOV2IcH6UZHt
HpTXH8vbsv+LhgFQcIkXRfpVrvvbnhN/FEOYuzNumI7BXjgvbbIfBStjWV5dwdU/
Y7KBw3/SgVQ6kI2RmzpKDlmX6mKM7zPXfmME/1OTzmNRWHuay3c8DXlIFuL4aufD
caMFszqb2ZVfrzrTdwGtSZ2+Q4drH6pPRvBpaZpOKA4ApbpigO8JLfNg1mMwBUoh
D1ZqvtWHYTdCWe5dbt+2ZsKevSxj1qd19NTBJpF5MYISmrko/0MkfUMblZSBlzyK
RJ+EN2VmvKj0b9bpcQu3DGMGhAkT4R+JUDJcjq9PlEgsWzgXvbCgB5WnQRYZMIRq
wyDbl4QzHQ54pqvoYlLMJf00mPW5QbQmDzuoPoOZVVl/WzN9b4qzi7pn9aEayART
pPG8xGOp2DFgDPEmK5YILgENMP1hoxwOuwcpdpKY+J/Lo6WuT88DjYkqCAgENhzH
mwTt5llPXdokhl2F9TiPvfrPYJjuGhu1qFm88+HiYAKMiBgFUHzqGNDKUzyIQK/3
i6c6HSxB+XN9ynGa4q5lfUpKm4RG7Y0Xjd7CwQZ8dwG6ytZaQ7Y9RWA6bwTyx22m
VGgQ63NG4t+ODQ14jxQGFUXef1cblts1ZcCEtEU2RATuO8OMmjinR3Kzpu7ViF4Q
cit9fwG/b/TAyFmjDn5fLmstl3sGxgkf0qgkYVXWL2TayeCGCyCiYXBrleyEchvM
RXoH0kXI9DM3xqvKXvpJbEeB4hBEGc8PhZJWawm2EKGZi9nB7RT58fqVUuyHQtj7
jk+8rKjMn7BtAvI9OJEnyOdPSuohj/vZ+wraey6ySxqONmDvPc7HSd0gF+xsDJiu
J7QaJTmBkVYzdJ1Hl3012tDSC6Kv3Toax26ME8f3xcfpBgix2ZcbcbA1gD6ufJia
+Is5Q4OaSOuiZeUWIbm6IYsqE2cRxTBhZmDH8f7QCsZNsbdVrI+O09mz0stGq2dM
0F+RIMP2D682kCK5fZtJzy0gPeS1A3BtjLCA4qMvhe7F738cxP1DcRLZczOA+M7B
CCPXhGO49b9KjI83kbCix6BgfCkNYKXF0w/+Rjdq/DtIGZJKqyExzvHGuqSAcolJ
5s7DvDPVOrh9iK+g1aekQ1juvQsVg0t1AgF+HWuwhSNFUhaTAaIckDpYMtaqkjiH
pFOXQuGY9yvZlVw+DIqWYt9TU4urYYN1DFSODfGZ6rMYF/YuTntoMEbF9Mh4CqqR
kz/tT5E1jc+t0/2NcOKrdSftkd3Pv5K/dGCf8wveBgF8B82s9cfMGwybKPY4gGsR
09ps3VFKSpP1xCU+4w0KMWYifaeqNARnLgYPxlOdvry+65Msa3Rpg6jiNBQO/sY4
DxBRPvY6j8axPN7PNZX8LyQPF4tNzISB139QlLXY7iCGTZ4HPYl+OFVa7DKyHRza
xurrukMwgBlhdIf0ristSBn8Pr2pdwNPby5dKv758y18Ogys+qLuQwx763Usjl6h
gfCsivjViNX0XNF7RqLpbfXa25iwv7BXaYDAl/GTFCDp/+6KSQEmhUW4xvIqZXxb
DmaDAFCqtuIdwi3aVqy0U28L4Tk13ccMuK5OE1lvKDGnrRINzZ7itrlIrVD5kGcJ
NwPqGGvjGvstF4WtvoJohpy+8wXXazwUviUHPy/8SV5PbbWyClLHAhyevduFVTRM
ppsCcXpr+j1dooHz3kmKXuypJGS0msCETBKl0Bqgb1k2LqpUyO6opKsyD3yhy0kI
2O5nUQF4lbsTL5htkHdK0BjAp8JskMCn/EonZnwHNALaIqDp30wdvBDUvptmz6dF
g1dY2EzGYhv7ozM8eJkuKBcSocK3Rl4QDqmf8rH1s5fjpVHF0FRYaOQ2MUzDvQxj
PDijP9z8ixruZ6Ej04v6LqyyUg25grbFcdSBnbO1cEwVdAXzhliK/pYsHeJt7Ra5
hDtJr95VQN+9ZpgWoZ4jpg5HaJ/mpLKad6PTMs6w0yDLQe37qLqZM0RMuYowT0Vw
Bik1yyl0z5hD9tNpZH5gtvtZxnTEb0CtzCYZIHRbqQlZUQFHGxLdkxskxrSPdZhy
C5+orog/gP6+l7sfbc1R4pWrSqgXP0Hcs6b4olq7zN3pjwhVQ75iOWaISXyz1sfC
L0XC1egnI/hSH6Z3VZElo4AG/YVUKd3rg4FODz9AuwZ3ilHPSmmAbSPyHhvdoCoZ
p4HdU/PItCMbQsyvJHddn2/Kz5Tj1KP4+C+ysXoOASD+Suz4J1bXAf7eBa7Rg8JM
Zz/OePyj8G6tIYyRoBTVOdHXDRXYI4O2GzevwYTBverm8T2wHqsTBz3FCG41cHpP
kGtLc4dOyzU0M5QuRReyGlbt7jRs6mFA0Tyqj7H+HdxFO7xph51fE7paA4DYSnpV
yFKr/8sY16Utlu6Nj+NZApJ0zNQeVYx86u2pFAnNOssHzaFJp1ibwRGcdqsHQ5fu
b05n+oX6b+U6Vw5xOflmag8zaUxcJNoLZ8zSIy3ylH0XvR6Ht2Q2Sg24W3BteeRz
3MhlORxk3X12RJeDQYHhxQloZYWMKSGPQeF5qc2PhwyBl8QAJwITHWRhSde4fXUj
z9yUitPzqloHEIiyEqgQYdBtLQiF+kuVgOf8JY/D8SEPiiYl3dg1QGj9qz9s8fTx
b1Gh0uM+pJrLK2P4LAz99VlCHrjzKSVSHPRU0RtLHdOBT530HJ47vqU67OL7zwHg
e0jJs618HyRvYT2y0M1cLjKC0lcSiIhc9+TUGr+/DGosqUijff9Fz/O0o4iX2MKw
JWV6IRQgpxKumZDLVMEholF6jcosCEwqneP/fQyueaUQRakfc5NmEMaFbMl00UZP
u6eoPIAea8Q8VjrPAgKjcWWdlEdtQLUH8VZKiR69t6ayWwm0r4VsaTn1Fo3FPz5E
6H3fmMpzfUAf9h41BixemUn41d5ap0WYVIwYqx+ZZ2b2yJPp5j7AO0oILBiCTpwW
Ll3oSP4RxDXCGjYfAttHv990Ng2OOVSQBqgszQwSMRKZjuddozceFICAYe70GO5b
ZTMIEhUjBYj3py7z0o6nT4AdLSVgPkMXpZtiR1De8+lxqieeuCE5u53+vZ80Cuna
/8vQObFMhxLbcEYyLuDb0SHP6BjjdwYNrFMp6+WyzGrNHt5kEypKDAT5vH5Hb8jz
OS/dffCqtC11pPApZoS5rVXhkx2P5u3R9fOFq/zZ1LT9IUOWZ4ucbMSAN9dT72eG
st1fJc65MA1Igcxbim9e5de2BHw4SXQ9p+sNpyKLZJlUXjKJWiymYgLeRS3QdVTN
fr3nkmLblfiAZhGtCay4DYke1AM2yV64lo4bt0N6NFuH1BrJJnPfBcn1zFLuhFXU
8RrFNC5tpv4g1tMuK0dfY/FDbM5I6lEsJdvyj/ncxpBFMt/hbW0gSux4W3W0gJeT
ms6otRVVWojowt0JUqchSLsgTwWMwm41was/eGHa1S5iBazaXLfy9Q37sudA7dgD
QGxraj43EG3RW8vTUYQFVyaH09S0bMaO9fRMiv0joqHii6qQHORgaoX6gaFrU/Aa
drKv3b3d70vIhlWhC6pXTVshIQvvjV7jQyf+SxovTzSWOrjy5PV5r4pH2H9764//
6JXY7M4DDU0WGtlZgjsbs1ZFdTmhEbNdNgHpgbkgN8Cf/R70WTkBicELmRZWgepQ
Or4rT2Wq16Whq8Z+U+HAfkPep+9n3Y1ju7Qil7At3n70ALFvAyFWXxC5sou3gH1r
nf9lJUwWB9LPzHv6VogFYIoGwDX1rOrwHkATjQCq4YzColnJP2xMyJDbFv/poo+z
i36NLjzLGIvWNOXTUSJqFG5nGvJK2/rO5UyogmzVX5UyWwWdWkzfgtKm8Wt8G7On
DG9wxXz7Xz6F2/60NDG3Y269DPm2pEGIU/ZHJD8tgddn+NgpkEpeF7B385c9BiGL
jw0hmbfckooif7+G3sTDkwhOZ5Vmy/RCnuNi6hmRab6pp9rmlHcYYEFZwEd9sYta
NW7XyQ+3YultsYqaR2w+OjV2iVc31jvl9H9wIPfw706Bdrov+wQMgE7oflfyqX2a
5eQXHGOAHDyRF+LMuX4iWNqsg9zBCFC297zLJrMjFjEH+Ezio+I6pcSX3s7kmZTW
4euHAQzad5N5j6zc+nxjtVQwEQiZ108quppNJeMYXiwa8rUkZf6FFxtVhP1lyLvH
JjNA9jGBUgFwEUxVdAzz/7oEUnXG61obn7XJKy46o1nk0Dw65+IbcGzBPXaIE1y3
oMm70ouyaSwmENKxv7+asA/xObIDeoQZSRVcroK9GMwKns3lfiFz2oKzrFwD/Olz
Z2UqDUe8cQSEXF3cY+237lbAlSv54o2ZdZssEoL54KMP2VxaTAw21Fs49i2R/Wo9
7OZuGlyc3JR4ZIr2z4doh2wKBUc5H74RXJ7lN4hcIy5YFhPIVQkz4Knk0R8WNiZt
GdOoA0c7SeZ8Ytzw2rfBJl24cYuP4m+ZCK9qt0xdIc0/ps3Ii/gMxj//uGoUX7Iu
J/sQ4ypQucJXlGA2eGb17gOgnkgUQLcCFszE3T9Qr9cjETb6n0OZODnASuAvw3GM
uq1fxqxLJyWImgoZBdGkfS5I8lGD6KN3bGx8ixGrXI/Dd+FuJpr61GflWwa80PGc
mf7FpBUoZYQeHKMP3QlMED0U5NgrO47RqUKG2QDDIchkNVkmS2lDkmElngyThbO+
tqU3bjaTAlX/3tJQXJQSdOLlXIQPT7Dcr9p/JIE7WTmtk3q/dGd4dQFbJDlli/iy
UuKckIYuHwtrk1iZx9gNPdblyIy6eNTo4cwnC41tg4t0s/ReFOmzIwxJWetZrU97
+NzvXdM4oQxZNO66Xc0Y0gMhngw1SQY36ETKd4cvWFoes2rouMEbXCObHvKtY1Td
BADAPnHOtW0vvxBv4o643aZXcTmRG/TSFNylL5F/Cp5oykfSz7WFjZuH7bFP/d1F
2U7soy24Gi6eV2+dtgEFr1pkh09ubKjpsBATGNs+4wDGuBZkAgEZR7i+FdP2wtQg
lq8m4RyFhizBjRMeRrOYZTBZR3h6ukn+NWrlkLLBizZy/VgZHg6sc0LRIzIw9lAf
O1tvF0Dv54F9y6gS7V/5xtwCTgrn9p0TeizWHCW5YK1VyfREfjtpYsRS+kugNdnG
kqF0e9LZxQz2JHWUcF2R3J47a4K52v8yR7V7eN1g+duQiVYat8He17LIE6WeGHVW
UE/8c7Itx0Dyj0Aq2RCoRLfaT1AOKZNy0GF71+xd8Z1jSYtWmR8acNobt561DKyI
WG9oaYA/Rjm5pSz1O2g5oIDhLDqNWN0S16a3jsQNXUSg1psNL8S4M5yRvsb0TBN9
Jmb7Oi4tO5AN+/weUQtcJe53s28FpTpId6HbiNeaZhAacYNLsAcPFzx3LlF7L7zr
/oDmQ4HUlsD0eaP7m2lcqVHhJRdHjWNjBQuGkw66fNXcuVvZrWwWvA984rcttdt3
M58Qb/1K9L7pHDxBwS+Q0kwp81ClNJgfiS7X/PsSZskEjLh2+tQLfKlTK74DcV5s
XlbDw28cn9YQZw6wP+AUlsvqJsVZ8AUVB0kYbldVVD7QRDt99IjRbr/BBptSm/Rs
5no2dojNVHARDnO80ygCXwVaklhoCyLaFyCXJYSbYiFkcXPWMNVIeRTFmpzFQlwo
TJbABbOQvUA5zqPlgZUaqACdG07b7//rwdaDk7sfmbLXRAdm2R57wGLUBuvQE4uf
JM3ieWn9ykGCVdXP0GHx0P6f1eawykeSxcsMapyVm6elsIDpNG5RRP2cvh/nRbKx
5cqm/RM7Tc6YwjMfOwkRmWiSgXpWQEhnfpKLWQ/4JWX7mgl4/nP3+LTJMZ850Bi7
mFGHvSnsKXeP3qql03h2wSAKHy0y142KFkUaCyTSZTEisImDAWjLdanhUSyHePbs
2CGFVutnYjc35nluMdo3q81iLxYa+Bx23/GJLTEswLc7/MQfuc8gJseRotedTFj9
0rQaKJIVgLfQFhnc3kiVPc63MLiYn+wkK3+OiLqntFCrCr6jDfxivh8B4fDuovyk
6I3wHAfaY1o9lIjJRXgQotyZPB9scBuo0yqp4klfULAO7TPOb0GwsRbXKpxtF40x
yI4AQSe9MRqJNLHY8SbITnMffojnL4VfQmprG2rpYyAf8STqKMbQISWpm6sqzs6q
LCl8ipk0Xnyg8ELjBZUACrUXDmiuMmlhe9DKM5OhXDJtCjUn29jAKXbJwnnXQGHN
qEW0MzYeRIS1t5jwc9XlwZ9rZyOiK4WTddu72AAAdqsIebUNcK6zS2lyAgnKiiKS
rvHeO5/qI8VLEwnUWSzTcQc2NU7kPbA7DOrBIYPF9JuOi9Xnn4oqd3mkkhiL/Tcg
CwtYiVRAXWEU8jvFcZsC26ut8NY3xBY90xHPcLKhqHtHWK7YxupwuGdzveVsBPQb
5N29xgLxykkapumDbG2GNWnujP1VhW5LCLVC1myi4a5itpvZNrFsEK1Ig4XiAYhO
5tckOL1ds64DAzNuEUyJhdBV+wOvaoE0iFN3z7HPdXX1SsDIqV4i9XBe3socIS4a
b9wCmHawTF1wkv5JbhApB6F8f8CAreJRGpH0Lv0Da8msXaz7fnt8o/vMZAFzx6r8
IlgdIAKwrOrl02TKGArXsrcVhVXN4xvtEgJ1ijQ4zzjTkB16kjWRRP+lk9VRrPk5
QZnK4eXeVM02htRLSkaqVOQECk397M2Ad30GH87b3Ou9lyYFo4ODqbsXdQT3qfBW
QMNyNLDQANChxPm434m+v//G83HIsCsHXRnTWkuL9EA9p2468SlL9o/95msuTjBm
+2piqPbklpjOIinxatVGqLf7tXg6cnJiiPyR2nZ+1KZOvsIj+ezanLZZEjPcZ7B7
aSkj+anUcgIEgMva0fK7CPZsODcT6yPx+EVuFCql0xHeOk9jTO6TddJhuWDJ8aCn
b9swg8su+Zj0B9zdQ0utDCCvoUdVEl9CvCN7PrNY0EPFNXmQ7YQdcLDxrmIyK+06
KzwcSODc1l2/ooP1b/7Xfv88/WbXV4srWj99wILlQpza8cu8WxwOzRUhBka4trnK
TurJ4JLEMBmKrT4xvrFUPwpNjMHweonxrkdmrOcWU7RO5A6J6vfENV9YMde4NWwS
dk8lxxJ2NRrWa66DNED8MHughDywU+oIRjp/SOhxBMLjLROL8ZdtfsBl9H/U24vm
WyRDJ5bihW1KxciMMwJD4cYQ2ubO4H0oV8mDMwsc1eFQjZET6XJH1V0HKsuTpEA7
Nn4O3y+MlOSqCj68ApZ5Aad6+VakgaFo2Qt04TSBSvPFFlpRpyl9GpNwh+CI/+eN
3SL812FHlHOYbGWG9G3Ck9214K6OSHzNj7lW0UgDCyHzGj/+UmMNLLUN2S+TPGJ8
EPbBdlIrYp5TflMM7bE4AMtoFCV34Jf4FDUDa+b8RHGs7eH8THozJSo+NIzpK5iy
PFud7qnFG+IH8VwSl5+YXrjRO5nNPcALclce44naODTuF1h4eW25ZUg/Rw8hhvbv
bxn3gQcDz1xQRbHe5n66wxZhIhSr+kH1//a/LI1ey04pIAWrdyg8xSW5dWx6Yqhr
PlcS3nSXeWydmd3U92KavTU1a/1E4LSQZN9jqoW1Z0MiCQ0dUkjL80hXTgESqmn1
KK0GZa7ZtTsb6rR4F1NiUN4LAB81QbcMlbsq004YL6bxF5bv8Xa45mi7cYnrDSXe
+P+x2GSwa3z4y/9RC3Si+SeNwfcjeAR+9XbtU+O25VnnuI2ogAS80ffkjfHlVPtK
EduDqrOA4HMckmmINpcVQweTUKj3ZYqOMyJr1fQ6hPsfXaNneWeChUBtxOUgaAku
/j1mTEBpuiTd9KBSKm7uK5cF1dJVB4krta2tTfKzk1JZoJmRQuZQiqodS8IlyWLs
osgsTyf5PFZ3kbESDVmXmIVgJtrvUCDTYxE7p+mn5vrqmddFdDhgFpHi+SHGAlKb
9PYeYSEW/eeOKgnHHSn/iTUtXNybIgOCKa15oMyfqSoGfnwk6h/qKcksWFjO6U40
wUePkPHwoiXr36wvAzIYIKmM8kYSPmZYyAnRA4SKTffirgwEZqIYrEA4jTsa+Phb
EZTQdZy+xBr/T3U7Z1o2M4qHa3FIjXJ7XaSJ0VTjxjVbUqo/os6b1mNCu3wtey2p
yt96jP043POUoUe79Z9glnjqJifukYPzObg0L3ndxEkn/MRdm7aepEbXsmDA0ter
YmT/nUSx2QSWGto7fpO/xUBMA/8lsWMBRkFRsQgDm8SJQTKgEm1cWn3Pc1176Kwc
T+grnf9GZN6GOwdCCjBU4phDy/zoanvWOCMYdprp4vcWs57fgP9Z4LeRCdQ2UGA9
5iUr4QUNveEKesnZQPqWN4FhZzDXbZxgBhdSiupWsN0KSaYFQ11er6M5Ip9oV9B9
ag5Kj7gK+CXgFFBwT2Aoj518hJ7xfqRSIwip96SmSNnD8hAV+CcMxIvtKPqJKAxH
oCemY/Tmu8d8GphlPlLfiP4+FkSL2u+coFEAV6FkkE34p2tkx8MOlM7A5ppUx3qN
WPm5py/17tu2svG1FVwHxsp9ulkYS0lEUiXrIEnfkjmP2GtQdW9hhB0FCMCwzv+7
GxvL3zAwS5KdIGTY/pC5BRxOMg0YQ2BUxnh1fFiD94X9lkrzDjsPGJm8eKLezsY+
IB8zTVotOEyC57jyDolf+TKa/W2j1ipVNhR5LzOwaH/0I5XlMj3X+vXdTA1rSY5R
SSptJNQJLenvjp76tLF0n9lR2l0qOfnp6CKuJhxvEy+hMhlZvCliKBcDt2Aqbr3R
hTwBylWM+Xx5vYEF5GgqHHUpBgUctR+wypKGwIp9FueZQF+w5DG4aJx5wA9FTUFu
/CG9tYNf58K1DFdRElIxz9v5CG38Rix23s6vNOiCV8izsKDFLAhd+ej0FvtS4jp5
voH1AVrr4Vj5YiO7cds6WhPIl20Inw96H+TUAc2CsO0jkn2O35CCLBO+00OUBPt8
U/b4T2TTNN9+Io/uWOyyejZ1pV7bRLPTSPUBYR+N3VBVnwMfCyh59ZZwn+WW4qp+
lUAUGkAO6jeq9IQpoH85aHc3CEV6HetRjVguyDPRSiLeDYk5dlNv7CH+oH6z6BGq
ggP6kbHulf24BdDxD65h9ry5qYuA7Yd4UeElyUqBl6riKds1dVc34Vq3jvar9A9z
4K+2AEotT576wxVcYl+KU3PTjazjqERte6P+vQQiaiDKZLwy2irz6ZaxZa2NYEE3
FBcMS8q9bN0uuZUjMYd7/jjPhWyqCVPbPQvEfmTUvv+qtxBSKljJ4b80B2jsABYq
WqbMWqYR7oTC+fJQpmMeFBpbgpMNRoxyA+cjo5Gki1S6LJVL5pa15UGGbQBwsI9r
/rx8khLH4L0o0XwhjplcdvzqWp4CqTCUGEximcPwG5HTRATewFqWJ9dJLl/evZOd
OlgtZxo/xbtig32cDr8bOSgrQaU4rYXNTxPqphhFhilG3RVcIu/C1UZPJ2N31gOD
yADae8LLu7o7DQKUJYr7rSpoIy1kYqcoMH4AwBTBR3KoRPda32rpUA3nFpZv9bJ8
Ia8siTeXVigjVbjPAT1nrbqK9sCWAbo+DfWektXk0R/64FfGc0K2mJZb7WA9G/+V
+nG0at1NAVMK22noCLmbFw3+P54VQZKnWRzWKht0TaQTvdWbF4v6kZI5+C4k+07G
FtTQeVCaA+bgWh38jhQZi5xYJ2LYTiRSx56tngolGfTNvdvV55t5WZJMU5B8VIxg
Yg3cDjkvjDbImefvAAL7XPzXfzMMzYvbHOxBfJJiqnw4VX2wGWigz8Ltr2fERwUm
SBn7oNUUQLwh9A3Y/xIfNwqIQkbSu36t3Pf1sBUgkEfUHvryGVuqVRGZPvWKbIqX
d4/j6MRuhd5WOcEz6kZJ9wwcx3Mft+Fd2hh2UhEmapDsRLXjapwENdeO+1gBV85D
CENZZ/mqpg6hIpLJ0eyjxK7UPF1AJF2AtCj0Oyc7vSkn8GK0zOcXJOihPuH+3MQu
YAcqqJ9hZu7bxn5p0KVlCV85RZ3KGz2nnawhIQZsYgQO6Iy2GZ3j9bcxScM68keG
oC25NaAxl0xmpWD+8nf++Tldll6BNEvtca2hrWdXYPE14dQjtVfxVNcjOqN+badP
XMKmJ1pLW3IiB6B4D2UgreyAx+4FEakPyPWVTgvCimVCzEvpQ3eovtkYeqaUF3A3
GolEADrKxc1rdNWonjBaJLjaA40PUOeVft29IcE+x9qYBZGtw/GJ/uKxkGAgFkfn
GsA54QYmlnMsckNYj0nHutlVZlF7Qg1vFAxSVTbyLSr49hSKPFFGg+1OCDAKMNvD
YE3VG2xi0LyXMi61qmvMC5J/EPtjOrgeahu899qwerVJdIlT+r81P+EKBjS8smI9
fPUuo68DnIKIHXpQgGBkuSHzi8ZVOTOMhXY/5sfQ5l0Gp6Jz0gPWOmlW44WkBhrD
TfzPHD/2PLRD2olXNiIoOo24dzjkBlhEAP4F6boxOuXATOFnHUNiqjDr+W7PyrA+
BdP4Z2yYqSz1pVkROPoM8IZFah460cN9ws0t8u7gaai0SkGnSYNIbRigWcxctDFa
ZyvV0WCYbMNheYsatOwqDOV5mMGuK6Bu9Rlh3TPvHe/xaYS1TPMyLAOVqYPHQuBR
h7f5WkCX4RbUezygLzClbuiM6YpJbV62xF2C5UshkOUP5BiGyQkRX3if947DMuw3
rjyEm4WvxUVKZm9VRLp9WkskaN6o3FnX0JChCRiEhOnSeTBSwDqPDx8Yh1q6xl1D
IG0Fd6z7XjkGElWfwxrMNebh7cKj0J0mVm6bBRDGYb+jV4BGzMvsWeB1Q1DDnKjO
nV7xEou+mxU2fWAf8i8SQAf5AvuNJTAdja345DTwsKgNQ2RY82FaSxz5FdEdjwML
HMXFQRFOEVib2iDTr6gVxj2j2xOE/MmRHUxoYrkvrQm2KVNKXNQz9GHYTbyOJP8t
+Nz9eYFkLGp44HNdMcBPH1d5052tWyV3CemvVuiDvgyzpX3Uy+LCxZjoMhLwKAVe
vH7OfF8HtR0gVbZWJydQ6rTQBEHglHbUtIscEi5ZXT2Am6IWjoANm612YhLWYkGt
PL/dIYjVlGCD9e3OSfvXApRhEqAJaZB+yzyTUAi1zvLZLQV7gmvtQIvX1wpIIR3q
ShOW8PhOFyd84CT0ZozW0/SPm52wEGMCFA4ksHDL7ZUq3jIUKwJbwaDoGOsHHfhT
x49Zv1cFuC/zkTMsiOogOk+WhTfqup3Ek3zv+W986mLjYCCmUXzwdJBHX4FUwmpG
+tWih0blUiM7HutFABCYBsGYKE8oZx5c5CgmPhfUq/IKUDQiA9gs/mxPxfLfhrGK
jbm2plcIEXO0aNlUnJmjnbPQYfS9AF0L5QLKg/ssSysyQkS0AygatdcVnKgZUV0B
Y176v1BVQP7eadfH8k+CjS/2fT9KYMATf5vC9Xdev+SIyxGaTc7BKY+OnAprD+bi
pMtnraJKxA3nvqSea8rwo2x94IUuCa30nrpmIZ6p2imVLfv7NpcTVeJrayYCnOJC
3maw/R8n5Kxn4JDMgQo/w3tDRCSRqaVAHl5hsWJ+XAqaRoXcQFWipsTmrYyhKU89
mYhj4NabHyauk4x351VtUPog5bP2U+K39f559y3Aj/L/4Hh1BcQ4rsnm3rl5wH32
+Btc9Z2+Q4kIP6Ouotxln9hgaD6OLnyzx8TH7KuD9kt1O9Ipm9jRs/7WSoiDvJlR
uciGIolEXulQ9fOVSsMlFyubDgfR22hqxmuHEJjU8Dnr5ciMdBgVGURBrborbk0U
8XuBU6TfvaYDRuk/YsJVCRYDPEmaP4kRcDhuIOKUCNAm791M1//zd0+d9pqsF4NN
Nqiq0XFhvleaupQ4Dh9jMdZRdgGT/HIac2hh9KwqaoSoapFJrv4ry9cvFx6TifGf
OcKIMLYydtes632UoDNgIf17eJAUD45x2w1G3xk8Y0utfgwGXWQL95YB9I1vxfLL
8+5IVAR3ASNFXwPMiB8EL8JRKAkWcTRlQMqumcXM8oG4aDhtjheFs6mA1miwVf5/
+Ds7CAaT5OdGbQQc1SWZE64S7N1crHIcY70nNZLwwLmZQ9GxuQ3WyMe5oM1sNIqX
Ydu3IZU5/+EJXuHG0PjvdFoQVNu4Hn7Wmq96Gy3fz74Hvjb2U5fPz87HcoR5UyPq
h2B0PPe3nDzBWC1/0j/Dj7/+VUobho0qsgJvfSAQC9eEHpthmzA+UznEtZmeI/on
ED18inswTODFURQoLq8wd7uU2Ychnet9sB4uuKlzHx3D2uy0t+Ce6DKQ3kjVWMG1
D9qZKLwpEJgqwGvkPmimJ9MBkQZqou+isHxmLdgbvCa16C9HvOkXrNioGFEP2Fal
J62/ba8iLVZTdXbP0XK79zWr317mfVJ7zFqE4LXYTfIXp9kzcNW7rs9wyJPeuHGo
I188AHw5hNKS1kvJctvxoG8isRJx3e/a0DsfJ/KFytccweXETUT5L7FmC4LsUapm
aG2sXVfTomKvyVP95P2e6Zw+YuIwWKsaMtVxxfWFHu9vTdZFXGvie95epd8PP9Vr
tSWMId2EaJmIXauh8aynoC+WGAUWQ7V/hxrProf8MewVj6jFqZd1jjGaW6n9EhL2
M7y1h13fDvvHsowgr81yx079NMSrl3GpqRdtkOOKnm/nSJA7VYfqq5CUk8NWqg1x
PviQpZrM4RV5EANabmmg0p7uk2V3MD2/8Z8CfmLSqxCvVgFw2DoyWtZvjtzojdoE
WD4WhfqBlbmp3xC8kuckLuqbJJcaDwvudb19wh45u9hPuxXW69usQNy4S4DNSDfC
YnrB5GP3xg//NjUwPnp3MHEtsCdAw7IxvQKID33m9gg5wXJPUqf660aG+s6+4q5X
pWwk9IDiyCXdabdXv8X6X2x3wKvXPDjAWdsndLqakGqkVSN8X/NGv/H4Z9b/VXEX
XkecexsEvGV8tG2vA4qP3LFhPptyDZmFBAv9WcYC8WGRe7hqQ7mlLwCs3yEOO+02
2D3cBcHEnKBdPtPrwpYx0B1oZMLMBoTKMGavwM/bRRAPAVACGKowB2z44CmZ7XZV
C1F2+p+fnP7IR/iAMNsnynYBGX731JPMxs25u/v4JVJhJaGy0pX6KJmf1G6532Z4
AUzi1ksc6JeTXRrS/XAVptm7Y0sPhABgZfWd82pWE08qrvAgnYLtUZqyuPch6N1K
Pb5GnmQi8+04e4qbywa4pAauctiRMaKZ0XjbgOt6IlZmvJ303OzxU2NteEHYvp2O
cQCA+U656GNN9AJmzp+lfxA1g2ZCm0O+pvhrYQGQ79npzA4Ao8WvOrPQQiLHlDvY
XqD10YxAtB9hrXCaUQH0SUagJ4NxbaUIe8igqwWq70Cgs6RI2DRA2Bm27QpvPa3I
RcPVaWc/tGPS7UnFJw5B+9hd57L107nLUK8Ot2RDGF9R7RdGy7P2vJaVzqYIMQ5y
X2k0webyJ0tNhghPJkmjwV096KbyAGaNqib3R2sLfc7NrL33sM+k24PnGcN+aR6l
c2QteXWXaVHL9oTh8EXnQQBYIEsqputDAXfH9gjXuz+ZhIChSyLqpRkk520UmGWj
/21hKaQqHn5jkH+ZBiakqYFVpB1BCLxIId9qZJVkOxaOjo/k2MOAwvUr6dzhvfE+
ngBflpm1sEO3+J2BY93/NowXhB2XD03AJ0pq5uFt3GdnAPEvMSEJYi1+Sy3fR+lt
/tmhybfBhevIxnk9wFo4zwtT3/3fo9hLq6pVwkMS9SrnMj0Jv2WcJrWZ+rqf6YpE
GDBicZ173x0eTd3gOPzf5RSkoxBqoVi08U9P9pLIXIWQNnBbrn3mRNbihXts4ABk
bmfGNDLmwtDIXnwXD4JuzSz3+zJl1f9/HQtiFTB2QK7uKbhNTn4QVPC6iVx2AbLX
9FInMRZJs3vMlitI8GXwnFXvymPRZcji/UhbTbqsNbSTvrnF6c5EcvbZ2E1IMfo7
RgwrnuXi6eIVRxIDggqSvhS5uL39e+WVKrlxwSGyR2dLzPPz1N0swNOYTWSDcB3Q
wQ5pMF27PP8dVKvA5UUCGSsjPXXabu0N/qRdUmXIeR/Z2jIZ9k8My0OAWZLnb9RR
3Hz/19bH1IVHCnKbzgGhepXdxjkv5N7PjPJMwaY9hfSjjEDuQ+IF4F5s2XK6XNuE
8wBgsTQyNuQxzxmmrzlEVD9Kb4+ID9xjh1t6/WfYXjeFXmZMsiyShMfU6FVVJfk6
7NnqbSPnJBirmVpItP21BQCQ1b9Ql/99+/WGeK099auDljks7/d9zugS7/7xj0qH
q/oLglD4yia0AzlVLgISiugB2mtRpNd1GN0M19X91dGllQeR8xuAFdkdbnQaBN4Y
1JEs2F1ZSAcWNRXlRtDbLOFL3p2rn9h3dfNtcehOquplVSSrS13AAdlqFo78/7wi
P1e05c68IkXuEEgQ2bvYHyvR2xNVvtBOBte8tB/s6Z+eQI/6V8JxEAXhXj9zEdL4
fr9BUSakPDstmlS4od54Kgi24eQeM7Ka+tsQiIkvDgYz/f2hLWqSwTRge8r6AJGU
YpFp9LqvSnDglKWsFTl8LHPfMy84zjgLlBO4hzzu+mfbvu6hysCsLIzVJfxULROu
TbzmZtm6mhX7yl4xQxlfKf7Q7lCMHes05ryDtl/TTnz4OVB7CZbGTJPc9ITnQkN/
Ds9kF1G5gzGUg7oRcfTavoAPKkz9VZvXZfY+LYR+iGpMwqYA2UinOMDJywQ5d0QA
5wIWSFgqP8HKMtMZZdNWjiyVQ2mJ9l75NPsoS21phXCr922jhG2lds0AqOsQmtMn
NdU6hGd7IBZQpp7xH+0AmWzohw0vRMdwgwozIPtQHf7e/DMDzd/b4KVZMZ95JJaP
IBEGmulc65kz5hEQmVj+lTy8W5gFrZbYbxeHdeG7AdBclyvS4ah4A9OPBQmXfGje
0XXJyzGd6HCyaNuRcptz3HZnYjhmaA/yegenHkYiwug0VfmOzW+ibvKsxgp1uIyv
VU4ABhWj/ceqtz1dk6cb2eZWfcV54K1Dmw634zLx2gaFnWI/Lr1GWsm6CZ6+025V
ynwwjGxD84DPTBMp2mGX2PVOuSCc4GHAOE9PnZv5s3UwPOZILSBM+SxoBu8TJ54m
WsF60Dq/pqwjcgo/ZhXrUoLD5xbrT2otsWV58ckY7BZkPO89TW4mNIdusQYHh64V
szlaUckH5V9pvrTAUmLTEF7p5r08yuqLHrEt3ZFg+Q0djbr7AnTVbtQs6F/k58tB
xTfA8Ed+eromzj1bhLsXzzGL+ih1GIXkElD9BeA9WfSTkyGFp8eJrCy0qI9QCVgc
dmVsNvWxcZ04JD8wny3X/bFQj0H5yTIJGThkEqlsyYuWqn/xCoysBhj5VNDtAPyk
neTxr6Krljaiv1Gem5pOpLV7iOYl39/RZV5bxHSYqxX/pkFnMbWZsz06GowZu0nM
fYzYECIjMOt/yL+TmauqYO0IQsacPT2mwMDLKpVfulymBVz7yxsGtbCmxnN3H7oZ
aKkNchjvDPHF0SlprkruKyBOGlEPIoKX6Ml1YLhiT+Ah9ezTOzxzNufuTDpr7o4h
ETTGue7wULWA7FbBvMKlnlbW2b2XyT/UI3qT+gXkkSS8rMHJi0cIS2N6VlIjjHUk
YBUVp6gIgKUEWGOxBNgRWt7UXVvSk19baqPN9oqCM9eOxeq+f2cRbWvxttDw5WKK
U09mpLam4rqNPc8n+QDK13sSUEhVo99fet8f9PVvFd3dWWzU2T2eDpwFcLuRhLY4
WIOMyXWTLwd+7Yy75NEb0X8diRLUy6417MtB3ZKO8jE9z0/J17SH1cog3QvE1BWp
sqnTdUOU2Xi6wVt4kdbeLadfQuIsZclK4+803bVCVzyTP0qllwSGAriiZfYNPqYv
M3K/xlUvSr0MSKaltTIMXUux5LioWrh/cri6hvyM1RXvCisGDOtXyWnfqJMmCklL
mAJKV1/KjF0uE7poDl/G4DMcGiF6EZAQiJIw+MBemc0BzQwGG8et3G7kzFN65PEj
LuAeEtsjyyBBjUXVaW1NEm7k24w2LJyZLVjrXrF2Zsm0WxxMpapqtYLoEoeFmJZs
gjBROyHZboHWJKtg4mNjabVqVUT9WsHGxJZJbBcGgCqPJPpuepAruacv28uCFJUa
MTvgY0Np+PqiAO2OALpT18Wivy2N5bOfpN+4f/ON0XVN0otEpYvLRV/CWx7UlgLz
KtIizcfk0az7Um3N+DpyupLWujmowqPs8ZBnE0CrEMfzf0OM+6lQBk4bsuhsscY3
d0HUv5Ie43/aSIcchvvI9i4ec8oGx7BhTmRHEXWFmupuCfOBIKrgV09wmAe9qKTw
kPV4U4zwYvdJMGr89N5kn10Bl1rr7hc4uTLMJK+cyc9lbtOOVtWZSg3SXgAakzNc
QZ6orAIGPfxGcASvCA/j/tiGfne4Yg5ya/TrnBMbc0r59yAykcPqhYXYEON7r9ru
kmi4+WJkY0YPlW3DzYjBXMyTDfhvok4YKC7RTi8sOtC9nMhiLdUr/0RUKqtsclZ6
mvAHDllWpHdxTwbajPS2G8cOYWsOG7SV769Xi3kh6nyjTfprVgff/pRJDXO2mGZL
Hfr0WffyavyPkpkYF8KJu4a1to7tW54K+n30h6vAH1SVe8GIpwEm0ao1A/76kRs7
7sPQWaHNCO9QOBC1z5JFxwlSk8d3xTZFTtDkj0ewKReMNLwmOWCCD7OPOGHgfx11
asMiXptJkFBDFNsmpij2W7nB1hvVFjcU3l/WCQp2bXJQo2lghy5jzd/3ThLS00CO
yLJOidmGjG6XRW87/Txk24mj+3oWfgzHaRSvujG0JL2uZScCBQbzR8HmHJz8+sSF
hipUllAmofuBdF8nWLrmjpmmPwHjTe9Ym2MHpq2EMRTI8/JsEhxqzJ/JMfwKKxvZ
TH8lM4pjKawvYL8U/lTwLe9+ntCGRiNctb9VWJ0rn201fp1XLL3D/vpd7Q3/cTj3
m6JkhrOK0dVm9Cok/eQ+nRsqgJebTB7F6pmFDfFsDH5bfywmtaWyx6LNv0RSeun8
g50DWi4yoH6aJ2iDjz4XsSGqBTIBa+c50oeKvRaeRUWD4CpjVcU5hZGhQdqWEG+7
h1GvHGR1JcFV5kek1ksQ/cAWnKN5zGXSC82R+5032ceiUdW0Bn6aR/MCeAWCanuE
mmAZe3DfOow2fIbJBOPDz24YbahYQnP7+oRVSlbsOklAPYSTR8NMJAmNTSzQPFEP
r5EZ/WxOhWb3cQYoG6j61/2+W3UveqNL7P232kacjbn1FH6K9WQrs610uHvBXHOJ
TK2P/lTIez+6KJgpU257EaxEHl3yQ466EoxxLSCFO89R0bmhS7AVqipdl0xaHtlJ
uJSQtxu76DztgJX5efXmLZTf3IvXx0SFTDc62tkP8EesYq4b+e+I3XI8n/0cXmYG
Yt3uKyE0N0135W1mgiCG3NtDNrebwJ2QI+KZEp7rV+qbbHiQ1ro11foM/eF7Bqor
OnNub1u5Ly1GtOMfLqwE63N5grStYZKRgUzFLgzCNqkCKhNpehXqI21u/2UkSs/a
uXGnd3BC/vZLcImGuNPnBCxaoPSzSV08OgAXuv47sue7eoyYG+yF/ThpkcVFZ+jM
LrASD+4vMT2ld1Nilknvw8y0qrq4wByJKsdF78t73CbR4BYihXnG+Sat7dkVkadl
hmvaiOqPQBQ+rkdq+7jF4/EA4cVg+r9NVSCSXLWhMQDpjbhSalaURflJIFMpZxNO
xuY3rxtc6g2+hX6uClEOw7Q499oYpXSZP0WKdP+Y39v4RJrUJX/XUwp3p3Am52qs
54lncmxn9jQt5AuJMfigPkSfcW2hL7pmRJYYfKS67GntL50cR5lZNF/XGJVHFZ6p
9EVlmkM+MWadNYq4xLKltC3yDe604rcLB1kfGfDF+B7bHRBp3mjMIT1OMKZC2Tru
STxqLjsTmPWFcbxGuQpVZr8YaGL+SoUZbq4FmpkOjaw1zWpSP2OOO4S2793WyFqf
HFiJsEZq5g6PuLO1RfAyAOZyeUsXwKLMtnUXst9DX1zUkDCWYGhZ3a3SOf9TMyFp
Jf4hQwOhWxkTO3Ndb4lR2QEdaG/5RZs4xrwctoi+WwDssbCUfaRT4Z/D7KfM6ng+
a9oJjQCB+1CyNPkoRALDRR3/vXOWsy1lKSyCoz2AH5L7RphZXRhwv5FS4MJfdcyD
FyELI5W8xk3NkCGWDBQL7jaeOHz6bLlNBTTNR3u2Hw9Wxaaw2VhEowJOzxN2Brby
MPutlJQwRNbiFn3FRYHEGf8C592QzxD+VqIXWfryAIpO104l2Ih4EMFmgROpazaK
VJs7OVT3ub6KPW7dWkfX+NGt8SdvaXtuNaelVc9VWdcilFeb0nwfMZV0pKTKt0fa
ekgEGLG2Oaq6QFRllErgcIqJ/Xd6z9sz5mXno9Uh7DH+ui7l57LcIYIP05mOYrCP
l5BUhqnpCBSK6wnce6IHFNavPqubwdyKj9JYJ88B2xy+O5ANRqU2gwjeLXJ2Oek0
BmqtCAifPvVb3Q3qV628qwVuiBoHprn6D5PXN+nwoMeruD6Q71dz3P0c+PhZLBp6
d3L6guOKJYPCBfPU2d3Zbu2oORaKmsOt2XtV7JqkKLGqCRcCWlf9jpnC1tKyeGZW
Sd7iQfFhhBLj8UGV1XkaTrspVJozyQlxf1NygSh6/gO/u50l5onLLfDs1wNjJs2e
qxjuCoX1uV+f+mvZeiQLpKYYpCmP4u2bDcCmrSZf2lSNtcdmh+Yd5q5j2FhfbcDa
wWsbkKB1YZIKd0jLGg9+uuTaFrmvaDuoU7Cu1j8G9bMlqWXVSXPu0+kbuTRev2fQ
exGLmU9f9vTGu142c0mbZeFJVsH3QjqK3COvu38GuTQz5fwnT3aT/p5lHAjpU0RD
n5JMvhv6C/XELi4kfrfQPtDXOU8Pl5GzeZjivo/GB1Lyqf/vN33PsD+hqQDSU+Gy
I6WZNG45BWiKJLX+IB2KsUWOOucy2JujRrbGxlpfFv/CIt06k8tK39hHWZ25LnSE
iyDw3bDbqbOfOHsOwUS0GWa52RevWYDL+/ZmhlKwvPj75ecXEEyE6RTu7tmOuYs2
vYxsluHGN6pZ27wxMe91Xrgm7WlxaHr09mSQIJ7GKcDPLaBaSjVFfutaGbcMbmJ9
+W7w9zl5bDbwEhi9iob+NY+rqX8gikQjPyAHi2Ta7ZLW+BsfDtSTdeFOzsBMoMJP
8cI1JkzueViITWx9m402uzeSQA8+OSEcmShIcp2pKqf6YsU5WKQ79CfLco8mQJCm
9WNnucuvW1FYlzufj3Kg0nY3JoOoisjksAP+iNYynxKC1jRngtszQAtpKHWAdg1V
kNKBhjR5eaIF0wvLcK0XsaTAE5Prm7rwga8suUrbV3GoYlBAViDV7PpjTs1uuGX9
Eft7xh+TCkO8UXRgHc9RcZdHQQa2zqYQXQzkX4FF7YXzmfCtiX3Hm8yL8JZGK0ct
FAo4rspg6yuv+Y5mjwIsjtRdqK0XEFR4KC/dXu/sW8GGF3cTpqsQS9LRyIOfeU5Z
VTcdI1vbDIogsDrnCIieEgrAl5PEZWs7YBvsj+9z1FFnex4jWYEArRV9SyNLgqlK
KcghmehyNRjwGPq4kfOYgaBMeeJ7vC4IROSfWH39g1rThv84gVDKg+vMuizJ6fwn
K6UXrbg9EZEVLnO8iZ4aoF2P2ztRCUyDlgEqa1bA8k2Yl07gboYi61FFUziUQI34
38bMWDkHDGiAfGFlUuE0e38MXntKH50do36zdtaYD8zgYRahf/kJMNLCwV18j4H8
0I52pp41C5vypCRogZZBam8loMOoFr0Y56aDY5Ykq8Ry622GO+xp3+826EX+vbdd
jcH/6idBTtLgEaWenHYjIkGe+3dl1MuO8Z4tWqKO12F41AlUZBwpQNtvYUbfi0xr
/nP1p+Ph09HoelEzGqnEsGG2li2S1oDSq36w6V0iJPgyRqxt09TWM785nDMPj1eH
SKsDROsPRlTo74xUI7sLCl0kLKn2klk3lv2XfTHKA2rPnqE2rfoGryn96XZa0661
vXVezRVpKAtrk9cz9F2jMnKxhHIHsNTkxV3ZH3sRw1Z9qW8N+bC1n4O+24mX1cke
9GPa1Pp+GYV46wXuljrIaftdjOhhq9fi8U+Z9DfLC8dusY2gvlf03D/5UdxIw4Qt
QFAnNKY0N3d0lawedqLdOTKdjIUFw8DC02P8Y195ywSDlBkvSBvoUXidUpD8+1SD
aW8uEjhb7Ygvtej+3VItM/kHKHTXYstNWL+DCAOY5TYzIngf7I/Isc+lnE66BUjG
sJGHVhj/Pd5s+afpiSKabiyY9DSPPh/Yua/JViSihwBZY7D+v2N7jgrrrzTyxBRO
zMo7ZSL/c9syPMmqiJGBWkT13+2lNQU0KjqbcNUpp6PjwB66sngXakQtjkl9gWJq
ga/IBKQOgnL7VQIKyn8cgVL/4CzEAZ1fFZy+dE8oWBoC300pBZP5EbssuDSDZgU1
vpBzrEAAhn5YXj6JzRBOJml0P6ngZ+bohpIOpy7IB8KZ7JSJTg0cKkgKz3Ieg+pS
aUbSi9V3EpSjHT0GKWhqPBLX7yjsvQiOhSXwFX/YiPn/IJ3B2uf2X9ENGyZYo4FD
wDpBDSh8GWzd4vzj6v6jJs6MrD7N7oIFS6v7wO5UE+SLiXq4vpOrWE0q3BJhA8Gj
SIBtYCS6P+z9EQFBcHclWZUsApmaoCq2Z+93bbegb7tTRobPJQ4xTEhS3ocJUoTD
BUaxZ1ChnKHtLfWVSoNRxjNGaNqBUboRz7gzwhOD3wn35E1A+53qe1UmMuNe6H/k
MdlYy761rs0eUrDVak5so8eOsaz7OVHyjt6cC6ItRhUZX/+Lh4dVcTn8/CHRBhEl
5SjvVrNOvxfFif4GuoS1lR8OTh6AXU57WSUf7lhb8VhTs0Lj9KX0TXi1B/Umpj98
ZoruQAiqofoYKmj7c6PRozJcbLJurYBMKbtgaoOeGC32axAGFsMoKksRDsmiCUXs
L+UOob9IJBisnAY7QNFBrupfetzgbEH6VpF4GJ2VJEI81maHWS3kpm3SZ1kS0qpg
qK/R86CBqxrLBRlTH/iIHdefPrtWSEUBFgfGz0jMPikA7rnhlmGES6HZ8FReQTcQ
zmmK+WMXdbBZgUNoau79iWmAIuWqSRaCVXsGn27AHEyfA30csBxiLiY85uYA5vyS
Ku98zWkXnWz8wZ7IMU6hz6jjvpZ8KReWGr2IGFoUaSNHaoz4uF2isOL+qXx1Dutx
NYTCQtcNUiDK7tvdr/6NHCyCPkqPcNQmsGd8t1zKx7cshdgjqXK1X/lKB7K9yi8q
DwSJs3uAJvpI7SFK6ql9ccyF0qKhSBoVwdg9+ETrzUQKHv9SG/F2a5/uehCAkQtC
tyRIE0nlCQCrHUVRk76tUl6VItfr9eAqhfOCnT686FOsxHK8ISocksEc4ZZi4KKw
vH1j2NUY5vcivMoPmQXqrKVSLFMNFNQ6ZqlKMcGDijNF9+BJh/H0qFOHt/YdwGRg
FBJtKOehM1/SU28MEoQV+f68iWRdV4+WLtKLldxEik3cxIgZHlpFFGZFHK579Yw1
uA2ynwUFUVXZARuXv7n+6HAAN0LU9tnAE/epmY6t0RRa9IjjqD7nvZn/7oo5MkJ9
+pJmfMoPhlOMTW8XBZosbFabHonxskS4vdLXU1OlndqlOEyzMEtE7JuLoJk11V0d
6NSP/7bUdaeHXe6EEqSk7FbJvbMhp0VPEwGMPqyLKZf88QdTdFA7w9kG5MPaYtxb
7yNN24Pb85EojBezCgQSywl3PH5c9hM6Mj9P/3RUnPcBes0/m1alRF6baruwF2ZQ
P6131F+ONgLjydSfMcipK+JWSD7fnkJfGJJ388XtTT+REYFwds3KzygDIIKIzMPC
722hRfAeZyfMLHtalnGrU6ZzvroIBqKGKfcfzHLNtjw5mtdtFpXMBbg6/xmb5g7k
9DwgIl8CLtg2e0vKa8fhKpD34qg2HdEzAsxnzwQFs3Rj3WSy03NZ7GNIm2ykg0BZ
LcQyq5aAKRX+udN16M2WWyEq97D7ilGBnqN3/6Agqk73oK8ciEn95DUkRWWfmOPv
qf19d0Umwvjc8grxRUDHgEx3nEvXgI2ZyaBKNPJjgGHxmFRxWwV4kDlswNsKf/dD
7PV3Bhg+t7bDhcUMoNj0nU+v2r1ILHcvZnSg/TwclG68jalcLbcBtOFfMHu+bdDf
2Ymgz+tDqcTPFovsepX2+qa4Z6GsncF+CoqpuXosHRNUY/JYNQJMVQpHi6U7pnOe
6GbkLy7sNGf0UvEDfvO0M6GhLPBikYbo8Y+7rgkvIdFpjoPK7SNNgJ/fVDmOtxXZ
Z53sKmXfwPjjvWjihepIM/gYl4b6eHa4t02hY4Ouf1TlfZPozHKBKjDbaG9v8s/W
ANpp5Y8xvhaW4rwNzx44/imtBTaUKq5R5S89G/gL9Nn6jiOuukhC13HZ7ZkM02b1
1/xlHoCnajAKjBfIytmQEd61xJ9RxvBD/uwqs57hRkjqr9eYWN2vbnnodvp3H3+6
+WL7PszWohowmNqHp9f0TLHIkm+GvWq85LWkOT37DLzkHtYpKb9ympmhnn6Cd4II
YLZPwkt0ffFkkNb9NNfVdpX1qYOmWtNcX5jTLM5ubGZYfynkR4XP+XdoF6BzgWRw
ijh46oCnpKyKV6FZhgc0W00itR+npMhCCzmCwgSvRyvEr4dvILpuVU2GIKxlMKJX
dI71Z05QRFW6etRbNDwytHEkx/RvgZ5XLfsAKW8Dp86bz2eegZrac6WeEsgwYHbb
6bAcGvj2bioh71obmJT7iFcUzkb+++POfNRg+6bjjxbdDPg2uaw/g2kaMiOSC2Mu
j4xq01yebTqVWmyhKX65TWfYT4UHw9yPgnGnwt4LAmmWCO0ccgfEvKWnY38FhePO
LhOgRZVTmDrLELiP5IaL1LUpAVsm2dyQvjbnmR+N9JQXAn9QArmuwLm3v8LCmRgc
RsEhH/tKFVJE9H6ygPMuqBeu3d/w61zH5KZrV8ul95kod480HAdTuNO/MCJVWs/N
qyzoBQ2dwZFNE150VWIp2vHWZjc6VJH2zKTzlILHy2dKKeGEw9V/Pi2K4+jGz9H/
Zavf3lLhY28yCt9f4mJTavyPHUt5dg8XBc9EHfY2gJWoaX0R7/E6+i60kYXKbHdw
PVZ7qLU+WHX+4mznZqXjMPacXyfSFxU4LfpaWR3HkerkMnxXnyexf39VF/yZO0Z5
5QbQfe7GbZC5qwQvDQnCxQ9Wj/9jy544C0QPfg+4N18yrS5xz8nQXSaGRiGd6feH
C2JEs0uweio5AePRz0AMM3g9mPsjLSN4vtRAhecMZ/BFjHQC4mjo/Aq4C9Mv0Rtg
omZ2taf0nbdG9UqpBVm5fVIhHL78KgWghwKECWw4GG3ksDDudxX8GI3k7pR0h7Ss
+URTni7dK6sQSGgPlvllgnY8u8gUV+k5CCdbJ5ci87wJpH2cIueTzQQck6glIaJx
iPF5j+/UsNH/rQYaNwxS6QwNnRZubI7mMj2adJHDfRsVg94r4BnnGr1VmGcdpXxs
PUi8UByd5cugXuOJLvi/L0ONi5Qt8QLq1jQSI4s/A5XHk+BDElr0nfnQezjMAoiC
d2HbNDAnOapxYbxq9wpUBFsNavbsAYKO9ollUUUz1kV6i0WTWBMMuxAbwHPKldqT
lTO//WEiZ5MEUVX/EXzg7vjlhQNRUvAga6PlqNkr2FAyYjb0+rd5lIRxCirax2jR
5AzGD7yvda4T9/koB/B+U387hd0Bb04Mh7H1hHGoOLkTXb91V2O4eRMwxrZIQusQ
lenqxsizVsFZtM0BcryLGVkOB82kl2xJimZ59lIkuarKKC4lQxcrqTuXSYoNEwQn
uznsYF+Gq4qQPM4RTwKAWTZqawEFEh9oX/YJW+K6RgBZxZ1RuTJGq21eZH0H5szO
xk1QaNeTld4A2CNzoCzH4Qh8Fw41OUMXs6mczB8mUj4NGNMZbRiyp/LLWbkGxMdG
zVaowPhpB4IiEKa4rpYgsohfNHhyHqfkv/MqWPO+ybA65vJuGXeeeltT89l50WK1
ujOI/X33H/m6//lLSDJHWW9zYlYop3ClSSxxx61oGcpyGAcA/ljrTmDBcjfNgVip
XnQ9b8gybW7UGkcVg5eoiMdMnck5LgtOz7E+Bd9zF2h+CBmpjWZKWAo0Ma5qjr1x
zNcmG3hCT2TGbrb7Pw3GdwDbOJjlL7/vfMUfqeAHs3taq+WiBs2izOgtaT87Kezo
fZExLWGQf12ISWXAJoFv2eHWiSx6LJ0UvNOwNdI2rb9uYG90zCgiqqXlO5Zoqzf7
w1ZbdGcO91VFm+JqoEWwvO6EQetNKwkU7QnksMMPmYHqyVOsZ5nXDb+orQpgCB5T
8cUT1Q4NzJ0i33wRpGfvvAwrA9GxMx8+oQoAD0qyHLxG9iETvt6hUIgty9rZKpPZ
P//IcDkrrPHx7yzHwE8BggeE1ZN8dM7Urb9T+jaytyQlecbS5AfC2Vw1mWrkECQU
trb0jvi4hmfqiQ14G8JX8mPaR4avNNue3NtqM+U1uLo+WJQhK872PIGhaTpz4DuM
L1XN4OMXOmRVz1r0OUVRRY3J1waNELEgWFlpFkbi9T6yXE+4SZn2yWOIUmmbd4d4
6a0ihQ5bKEZyHU3Ab7Kpyb5h/oDKTGgimvSjCPjy69TLlHOV68jtAUi1yZskDCAA
POnGWrC+1eJ/LukmSxkZ4lRktT1vauX6jDwd/lviXBGMx6tXUf93euLuoBo8kzvL
gPzt9F/TnYHL1KXyloPOQmMDu26VYwHWTDcjCDQEOtF54ZxKQpUUze1ohfc89qDd
M4Huj0yp54oZOoCVEnBZPlyIhKGSQ7J8yXqyPeuiBq60TyFbx639udGCJntPoTQs
JPKqiDXRGLa9AdqFlXcWIJ3uPw6lEz8eRRvDCeTSxmbRtu+8OxJtA/NbgGdi+5KE
oBH3nJWA0r/cJoFm2+FVZ9OVdAgGQkEIDbhYrumfIuu2btUlYSs5YdnOMtOpUdy7
g+pLEONHSY8rHzJV45awjOjmCT4hR38CAT0UK+KNz8npJfxv88FTcKHIitfxnIFr
my5EaAW3Ysvs/Ya+bZ00y1BqCc6gwi/XgsxqQfMHAtft/rbvrqbltByls7xBT75M
zWovJJe+8j4c67jUEj/4wzeS0tUzAdR8Y0Ipo68xAY6GdL6WcW16I56yVS8fYG4h
YEHKp0/DrUyR/dGn93z6/hWeShi7CeC3huIfAf4KXy2wLJ+peJWdnvb8SsNst+mm
SNIs+7JvljVW7D0XXMH4bi8ohz27PJvN+goUXSY/qLpjmHcu163Qpexp3g/TAYet
P7pLn/RXLHtIdJKov38odQ8gV4x6SCXws+zJtgZtAXq0tdmECcmQ0wPXFE+Jl37K
ejsYgmT2Mtbw6Hs4mPkESlZ3U+SAuY5lPO84XTq8AUweJxxPIptgY4NCPTCs8Ql8
CSzNbuVwsG+BB7SoIA37nezbbIKlFCqwhb0qbZ7BwD18Ypp3gri7INbXFEhp9/Mg
Pv7XE+xSoG9f31iPbrJFKlqkBey7JRZqad/tBjqZweb/m/V1mBciD6J8ziGw0gXG
e+bzmb9cNI5ClGXqLUZL3kNORfnBHoWYxv070z9v2Ij4e7kCVwUs2U0UhbYLvB70
M86Zz9anEofx/px+PLdhuPiS/CCtzpgJh69wYvXmb5DPX0DRdZhcTYXpQWPZMEUQ
p1/QZVlkxThwi7s1xGutn+QODFidjy57qv+w9ej+wB1AuIte0JDU+bDOyHwTl7wv
0MRVpBoOfxJkgVWDE0uhT97Fj8jQr+4cB4XC68pcM4Ng0gGkKBWfJivYhQbMZuP3
kTwticxWgFgoJLvv7wq5EmulEfa1Cg2SwkAio8St/Ir6M+NGaXkqLM5g9C1cYkR9
aPgyUq7VMBFmVcYt9Cowq8qcCmWhxn32nH2acosNBoImrSWqRhTl8Y5LWrY57OgJ
xrbLHxufS3vKyyAdeFPIyAHjuj/d1QMFxKSCTDWtApcIVckqfjoSKIrInQNogADV
el20Bb1APrlLbmKQhw2kwzT1PV56/7rXTyaOG27Zn/EdUVjZPtfLdzYqidYaelg6
AkQvOck4aUKn79xE0WGSbENH/wdX9INRGXSh+MEP+Juz+TJqfkw3MRG3yf9+U3EE
w8nePUZmznGn6VL+Map2DBscXx+Racy1LY9qaZ7h/G06NssEjXLAJRFWQZ6rjEJS
1ePnHQj0lhk34edYFqTg6TTTITAqpqOIXCIaS22hE4sZ9OyNWNKLB2yeLKr1Evp0
ksq3/0PWW9M2SagqJb5Lu/nTAOZ4j1qaOAr2oHLevwY0EaCDiiT9wWaRU9Ezx53R
pCc4rsiEWugCwcT4xZ9PeoHjCm/uHJvHoxYTZg849MsKBECKAM0jD4Lp8b/SDCsc
weL1EbhX6JLuYPfIf9Q0JLAf8HgFBB+B93kXRqWyw57Y1ZtTexVL+mA9Ov6ZbcgP
Zl8fQ52cE4zH6QSXvyUPmAwh4iCrDeJSYnkWnswxtijtwyxGkbGcpS8ZaYwrlik1
qQ+zBH3qc7to4mM9IEUT21UDYt7zDzgI15Sre3+pz34zGqloaLLVCXVdn2UpXIfy
MANrWqTAfx4WIzKYgf1vTcZxLmNNlfxhCPhxDL7IBRe8GP3r7Z3mPRU8BbZb1qoX
Zk3lygll9n91/S9p6IAXA6QTCD45U9kRlhseb+TQwab54B6kmTRufk7ZTXv4R79s
pp/kKwql5bu/o2tVFAQrxa6zHrTZgP2GTLhQYK4nIrkmpD9VHP9gBBQhHUt7tcbh
EJE4P0ensn1f9pmAL6dFTohjGrDmLnyZusnOBOfxhV6Clc+lY+F1DLGA9g+l+SdE
c79QnHE8UwVq699j6tgLxGGGEvaVEwdCnrN6aobs5ftv815txUURXRYlDUvJjvxm
hD8CcBjk8n2D6CC74gMFNAiQGBGGc2myPt7HcD6oBSGha+IgASuxF7rFlurgAegM
qyGNYtcb/RbBKZ5DiZUOi+EkJGWJwrEehc6zc+AjhEVWicSyRYGjjrAwuHwh5S18
L6RG2gIiH+UvoRqbnV2NOAi/yNzXIbfWe/k0hngp061ArlcWy1Od0LEJ8xK/Lqwl
O22d2esY81026HCoTozzYclPsOYl1edhqdoN7BBO064eL4UgNV8lk+pRTjnmMWaD
FSr6+hpGy8K5sgm8sjAAjcxjG94IRAcbZC2eFK/8G1NPGZaUoj2O3OYDgE1FA5ES
/jY//827MFRWnEcQ9lae8wJHxAh/k+MJrUey/uw6iUX8+9MQdYZYlpqn+RQ1xGBn
O6KAIJmBfyfbEdi0ZLttpE6gTvFexlkMx2WkVngBU8WtohK3Xi/Gv1T+WFIivqDm
84kM+CrwuJRpdji7aOk3/s33YGds1UBL+bxUMGJnfpAhshplefY4nVO91v2wAFxm
hBKRM2P9pUgV1HPVwXz5y4WW1AB/PIFH9s2c9uvkdX78Vqd5Ji3GZOefbxPCDsFE
CyEGYDZfd9GsivxIv7SnqXZaKCOFEaD006QhlKBGVSxuqBCRhv2Y5XxsN62sDK9/
ii6iMLYvvQI4csEVjndfr6IcPw+TRq0ob854V2nFtGUq9YeBQ6grGkesy1vnhprd
OtAFg0yKI2/PAjw+cqSLqQsy2jtqQoIJtboh8CimqwEneSgY3rUJvVlN63rEOqZh
w30k3ZnP2Du/W3XXQ2S9ParEXFvn6yWO4nUybw//zELBb+1ZL+ek5FALGVOiBwxe
CgZga8QWF2O2cnJgVAuxMNWqwJRQv33m1pD9vOwXgvWxIVd3rHLyPHsE5G/4JOFb
xlZ32GScmzq8kPUVxsQFcVTNRoHZkq0yKCKq4oEzkXxI8ZBEsj2NKWzfG0lZmNSB
I+APrhBvPhKUn/2IFYnd5tAG4BphYKJnGANOAxR6QkGCeSJG4aParTFv9fa3HW5i
7FCPc0BbVazPrlrv1biez9NtoI6DIMiUzI6S+c0dKeEnX4DgDf1JqSh0e5FlujTt
rQLoeUsS/oOak0TgJURDw8heKjXsp3HWxSiw1ZVMRE7mbWv+w89FjZdTIRG1uNhb
uqwF41GZr3LJ3nIBfMHyaW32xCMQJE4keSXbo8ax7bLLIUx4DkRo09XY3+TJFs0C
Z55eIhAKsVUbcAQwgzq9MejMKimAaPzOgppcUTEvfR+LT4wulb4p06ILby0xjSrj
+DcNhNhVE4ZAwfO2nxCZV4XLRCGi5Bavte8Cy2mF0O0XmpBka01iOggpr4CZQLMn
uSe/SQs063jo6s+EqFk+8OktI+8hnoQq+7DsEbOIHST4Eh82I0x2TyKXThiFfGSO
UL+Mczzh93I6ttpAepa8BClai0R1BqMxYR84BpE6Vs1kl/FOMq08QS6/ATJuHnur
4rrtf3H+XWcxTLFCdJ2Pmo40cdIF7rQ54WkQAIcwl6Ouw9FUUFvYAZ6U1pa/+MzJ
Yg2Rc7+WckW3hU9CG6TNLg8LG1Aa9zuOhIaR1qZaTM3COxhCUFMgvcCU1zdeklUg
mv+4iCw8BX/0d4QPba1Rs0bbJJMMWpWUMu5iw8/J8gsRjYtfxoOaoK/LviP6+ekQ
+NAles2HmI9bIhQAY6WhrcBiL5Wjq8i0Xd9feNpU/pECiijDyU2WNQSYsQO9/szN
J4wizfB3xuh+ilO/6V56O+jqdLeQ3yDiJj/B5GGUCivelr9J3TiHUADPESIvYohH
Rc/RvcpzkqPGHGDel+WrDoi3KcmuHrHavlrWsYpzhUjq90rEB2N6kboIZ2DdL76x
ZThe9xRPa1us5RUKrGvtitKd9os3esPluL2PxdfeN3G9iiLAPPLXKbHwPzVwx8gW
cKGk+ZCkC7qeT55XIdE3FbSjJnfw+Xb8WxQ7RjYZEAhXaFUN9wIq9SD1Zh5vA6ym
i2ou1glRx6RwEMD/ni/b+QU2em1ZZhe4FjMjQ34JYK/RLupijQSPXTekHycehVdB
61XlMf9O6iX6/3YbiRtfr/knkMLu0fqajB9GuOxo/Yu2tWwcBbBh0p/i2ljbOWsm
C7l5HmiuYGVCoRCxh7+ntxVHu3plRmZLPipDrVMnQs472X9apKpv+0pU0c77MXxf
I/JWIi+etr0pKTf2tFAMUXLGEfBVkkpem7lW6uZvCdS1dC0AdxvIXL+ilQBZfTw5
UHtwW5AIu7AfI2mM30UaPdGAtleMykeX5J7C+Bkq+8jLnc0Taz0txvhZXZcxBBWH
LelTB1IWqij21YOs3liYL9S2y/ikW52TYFXncyoBShbNs4pXuFOmtqvd4aikWTDh
BQI9he/okpg80s8qkARqIpG/So2VzOgXIRGXz8F9e0gixMU/mK4sq9uJYPtUogiq
lSRT12ZqqWEBtETcYhCZ+DsnxaUClVMW+D+SXuHlUFjCvMKfx45+z8cMiNlx5uEd
vT2T5lNnLKppJ35PRbpF9naTh6LSa5RLM6em25zIcTOPnlrHHkZZyXNBiPmxZev+
U054j86MpHSpZJwxM7Y+uanig66+9QM5jNhavdErS5xDkg8mB7vTNcEEhQeW24CJ
ADWmny5hxDqYxtg4FlBXSgvtEYeGbQ+o1rKu1VCz8qafiWRWGf9vxPUy/K78v5+8
dE1YD4nGGhZYSdxS7oRtgdzY8G6G9g1MF/X+NL7Ns5/4YSMzcKwKMlrFyal36oTa
+5R9tIYKI8K5i0HGUDoX1fCFV4YCJORcQoOK2EVvgdfymls37WpITCQWr8dLS7ez
zOSY6fWjAA/MQV2S/qbma2nk5vZpviMHlEax1Ww1E/0rC+dCCQok6pmb+S2szVKI
59UiKLWJREh6uIzbbS8H590nFsdX/zhYEx8ADGXClut85o+SK2OiUumf+F++pM3t
GUFfVqjUA+EkO6K3rlaDQ9o3KBrahfhEEM5I53W5FT/bGdguE1C5mpWqQIICtxS/
oDOhg16XW2cnK9chBbMY+yW1O+zxljdCEnadLt52AmtNBel5R+isNBUiZ1wep4ku
Gwd7S/scaa7nUfPq93ShBlZyrjIkc5nHsllKhxn2RAirG4G+aRVzdmqyScuKHBSA
QuJxWCvfLbZJCkhNJ4OktEBAxb16/Zg2KA5n6QS3OEjCBB/gs+XOMS054PjvIN8+
A1bggBWuZMw2a5w+UMuaN00+EczDFqlR+2WK6pYPu++nzIzXS4a5+gQpUEpJeguk
KtnhShgx06rX7JoXKIyjjAXHutXYZTPETmUOGr7aWPRhZqsC096dp7bRiKXGQ2WR
rRbaQoCxxVdFMeaZTc3LyOWWnW+jptrIg1QBsk6Fmy1HClDeMBAOwnLZOIApOZmZ
Uh8aS2dijsnK95bYe44OdtEZ2AAe4EPX5RICtdmF4TfmTPULmpgFUkCp6ufPyOk8
BjQFcXbI0EeD41cu+owHIqmWeqAobENX2ZbBuJ5kQx9bJpr52+Bp7DrRU2KSVqz2
ZOVIDR4CIuEyMSTbBOdL1GxcPXrcXjQJWOqrd44IqxJltluVeUOeuHWPSXGgFrxA
EEKOecEuN0NvwmadZjjJUcvRRKZzcM97DgXqNiZf8HMv1Szc30AlyUkmlCv+T+8I
G7mBGgdfuH757G7HlIhoKmXtwWP78e50CBsIFZgurMFI37/OT5lb6dAxQyAXrSXP
4Tsy/KuTfGgySeslhnoI3GIzOYUVYma6r587aqqMCbYCaRyn1dpqcKIL1afplCNg
TQvlWh41CV3EH2YIxuoPhYSsbVau4KpVbbw+F2kQWvFM+YoL2D01ASaal2HRLQfu
7gACKMWzLLfA7vr+aQg2PAGSyWONDHh/JX2/Rkw2PP/512rAx9U63QNepNg+LBgb
aZWTgOSZjqBnT+0vkHkUycM0QeEe/UvKhg5wpQvIGvXDk+v1fFsgHk7WLzXXsmJ8
avkU30QNso0sSPSYW8kcfEo635dnOju9zAzfPEa0URqhgSPXLI/HXrxFoExy8jSx
ezqA/fGpSiEhjXe0AqQxY/l8fovtScEUZskBtPc1gj5W3+DpaJqj63ntwQAh74b4
hXdI04Lm0HddQ+p42awB3x7B8s+j7fyMJB3feISExAzvsZQ9AmeCKcM3V4SdNQdG
r/vY24Y/q430xXKnIG7dSXIExeRV0fzHQeZUFFvHax5tuD+P5jWTA783aCnjDpmE
gPPzZQyQu2GzC1xDAk6SwPOCHC3dv5zidsFPO+YeEE8Nc6MjZX74XktpltG8v9oi
9c/wjeu+0e86OqlQoxb4yU/JZd2jBiBXHHu0A96dC08fgVDO3vfJX9RNYfB4GIsC
mPtnF5C40t7uNzV+St0z2d6eT7/iAAVuNq2S3bMecIOGNd6GdzEPtMBvQiBVXcz2
EtlqzkiPUU9gZB3JZU2vR2LOO/1CxDS4ceWt/mRWqXo8+OpHe03/2O2fQakPbU/w
zYBLZhwGHfm9sz2v/ARL4NudK7iR36PL+U6FHW70QF6I9pkZAzogH5tMfb3Nr7xM
d4c1S4ZlWxeolz3uuP8laDdjg0RcjueWz5LgOzON6c5X8M59MeB29JuOyFtGgF3G
NcLLa0vi7Zug/gsny7WhuA3KwYyPJJW0IZEC5qKc2I6emc6HKcSxMdpdr9b8UVOm
T11rvbxyVnj0E8jUmR7SpT4tqvqjPWYOCSfHwx8QV2y1Cl+76PVXLo/qBHQuKlY1
jApT1njC41j3cjwDuVqLIR+O+XHv3BpYA5Nb/ttU0A+pvzfl1CCHyY+JfSQTR8HC
/OPeNI1T4E3FJG3Liz8aCZZPZqMQgOjdSgOxgplO9BYe2EdWP1jyoT8X9bjunqAU
chuTmN2kLU+sqhMkzJvVH84Q1ZxEpRfAMugHdG/mF+4SMGo7LUX92t1NLdAyThuL
pBD5utVs7oY9NksrfHhNZseinqCxD4m2QV53ayOMffzXdvRQxZERJmGvwQrRMToY
VF2swV2Gt5T4FzzNS0PdxDJAM6F6ECFzn77+wpy9TW87PbbeCmZqMExDRWYLKvjs
yTvH91AhVzdCVBHVz43D8rZTStkJsRBr0uRpymAG0fUlhvEnHWJRtKasunwFxCvv
wNDRs3OkW1d4GNKBXLTddu6BG7YHfgsYznT172t8l/740wyZx4p19lUxJef1mT7g
chjfW7tuV6XMatJemcoqFSC5Bl1/wEXBAgUlLfI7pszX3Dzwixzu1RHj01h12nPy
G0zjXkfExLPtr9CnBQmm8wcArxJxJycd2Ettg3IrmOsuvURkWGAE+KQJJnK/A9qX
/5Us4gWh2MYgONxwnXPIhHbLez2fl3hYJ4Hj3fp3mS0VouSywOO68cjUCXUjR+Kt
tc09RXm58OxXZPTarA4nRh4g9XUiijcgjlQzR5itiIak1Y9UBylS0Qk6gKHQ1amt
0NSdFD5MgaROIZvPPZZpsqIP15bieOtkZL1u5yo/+5WcF8bCKziEyF7ezsCa2y92
OPlpoHQ8RFXmTCvOImlY93OsIpKg3qYDsGPwiBr04KnZ1oE+iqToZL8DS8JmWM3Y
9nfj50KrcTe4XlFYVU87p63DyiWlrRAwfXISgp7XvaOdcfvFcRvNKXkH0bh4vfk8
zxKhdmPNJ0RwEMV/LqHqzzksDmnUh1rJE4zl6zM0Y49PYz7XQFdQCIKait7iK4AL
3REXJsk/4nkHBz0urjQS0A8aAfeYeF7+fKbw8PTeBQ+0CDIx1dROGnhOpCe5mRGI
8AJ7uTQtNyQfxCc6c6k0HjZ8SI0NikOyRG0W6drnlkkzd/yKjgCiUntux3mEyhd6
CEOnhK/rqPFKn2CTwyHJCVhiUNu2SaKDLGBKlP7MUo/FubHl70+R6DhQcakK060u
+eU1vLKZHQwHdxLeUOX73clQ8vsE5YwdtlLpulh3OkuJEMV3cOJ6LJk793S8jFWS
b/ujrNIqVwb45A1SGfM+RlJrGSSyoL24+qetq+v4TSvpPMCVMccBuwVhoBstaaME
l1oBgdmHZe5gY0tb8jHHS68Ws3biKUQOMpvMbzGa+bwgWzcvdSX38U3TUbBK7w0O
MWnKNT4pJe3+bxdLVesjzSlr78aNp8acbaspgy470W5m65vzu/pJO/rJCS3/1Zmb
592N6OPYJlJimO5KsIuOwk9b5143D/NIH7XJQO6DXT21V+e5jQlsEQwZDpOrANAj
XIwy15rEBlIcvtGOfSw6nc5lAC8Tl81qfs8/AWXSM3mEoPz+AtkyiekZ9S26Zbjk
xIxW6DROEk+9JUHxdCJjd03KEo0pJ6gA/ij5rO6b0hOCrMJRaNVy99nIo3wtPFfy
I/daYIIGJgvFue7CnR3DVZi2L2POEx/vSxhAtcGUr+18M3QXpSK4C1ps0xBtO52Q
2c8YbueUHNDaX0z/oRFGFECoVyV0kKZY5J65AeLioquJPe+G4G6W38eQY8UXC6TT
wFkLRY7HyqNCznte+is7u+stk/fsRZZq8v8Angkjcp/ssgRaJi82L/z00Al6fsxP
zdTX7w//uHTaUsseGn1S5XA5A1SwsZEXwF7bNeCCwxpqMufmjm5HHGD5YF3uVF7M
DfW9DhpoYCbe09uQHWOR9+Zo/vMUrA78qGoMnj8XL5QX9UR5bSn0vpZh7nKDPZok
LKoldhRwvq6oPlmfWqBiOp9PpA11MSF2goW08HMd7NNF+rSCyM+NzTf8sJV7lGw8
5LIYWvTDZHvRyHTXSm2zCoymoFvIis322Fse1uR8pDyohF9dy6ade/bV2/nzjI3t
5nuFE7sDkkG7Bw3DWJcgDBVJDT8atG4oWkXWnq+Q8OD82p5kgIZ+UVbLoKry0T1d
8GqWqD0K17BvCEYuxiiDYHE9PUQEaDZw9Dw4bu+/qFTHqR55TK/IA3CEeyNo55PN
IZ0rZw2ruEW/A9o8lZVg6LpPgnDQowKtTDUxOZqSZcF3OqL64MLOtzeVbDhtAZy7
Ig43TjFhOrsze3j17uya4xNZaBtSodM+CImaRtEfxzLyTVm3VOWp0gtSrzDSJhoU
NDyC4W0+aYFrKaeHbpDKJtoFqjnVllCAKgNErUCaRCvM+/+/HJxmdNyFwQ5T2aRG
D+NSfm0zI5fJb+zusAJiu6OZ0GkmltHlyfeJCfGoKSMvurnBvCPpxzItHgIvuQDP
meofXMQ7HO+nTKN5/VCFI4A+O/r5SFwygQpruRU/ADMWgFkS+5qUajSRC3hgnnUk
RsOG69xsdhGyJdm2LYtm1L3VJTxnA7s6oJE4L0Us9V3eD1JVs9psiGTZhn/GMh/3
W1fFnNpxQn81fKnphzLVx2rvOpHrtFWv/6uVWyUT4ZESKZxIAM/5vjrcFPmR0UCF
b7qKKchM1fomhiQq/NQSru0UErBbk6Q/Hc6UZK2uARkbcODzbonoESbazjJi7QAC
bB610bam9gZiVcmQ+b63FS5ULkonrXE2vAT4y0/JsuXWpk02yEpR4//D5RZfQ49s
bwN0/qCwRD2Sg/DPRSLbqv+4kFZCeCE+RNSTzkSmajWPQDQLNKZxQnrArqlcmZ+Z
mMNtbi+G+eTheBmUH4x77k93koFss4MNk9Uq4sqLHfO6s4L87etAd4Kbb9eTxtRx
Hlq6RT+oOvjycsF0N18hqYqGXIIjhxycbWQiLLKKNswwZMk1LdvovN7VdQv+wBTF
Jdrddsj567ypIkJ6a71ueWo1XZgW5u9DQTgqqqgVMN2UxlcDn0hBvyVmxewy7Rnh
8McxIJKtu81fSnW8Bk4gCRp9Fw7CAKW2md0M7/HZYXYi7Xi53Jo/SX9fA9TZvZ+F
dugROdVTZYAgXzFS0/mJHWwtSPAqx3P7dxYJI8n22G+BmKjluFHe8MRt1u1huzX6
y4ja4gnzvHSsayzIcScnohoAFOwz7Tw3fBjVmPJDTD7TH/ck+3DVqkU287e5qiTV
v8y0iwoSxxKurRG/hrrLDxsV1np6eTySfXp0VKRR9D3qzByNiiO0nIx1sTKBIjht
nRgC9nI9PZPh56eQ2idHR67TFjCypZwOSogkOrMfd4TQjv/5E9AGxEm6e0ea63ET
MJirCw9tswjfFhs3ISfSt62g+Qpeb2k4wi0m56CHQXHcO346phxobml1NKJCZ6x2
67wJuKLStLiaMyV1o7j6EZVycyAQRmxXegF86jlEvNMWZuaB+19/h7sWJ1gk9ZgX
0rzpIusm5UzZLIT/NcP7DaHvcyLXS1B3eDl9C3EwmaaM6fCAKHnX2fx38pwWdTcw
W30lDsIsg8MS31apaRGgfw68SV4VZED+UezxslV+cOzseAKBm4E3RYQYyQJktVie
GAq+8iC1371vMwP1w+DKFX3cQBQghtpJ7EIy6j37oFHK6izA8+xxDAC+8Xb6MVg+
Dx4+nA4cHwquhB8jSBQezkhSCiM06i8WIEgaJCZbEW5zlgs8T8isdxZm1f6ofg71
ked8aM5cr7G7F64ScrrnlYPQhorhfU6DI8nqXkse19oJ+yPeKI4hbVcayZweMrps
3Ovnloeh9M8YzqRpNovMMyOtpJKZ9D8MEBhNcZsFH1cUGjdjvfCjz/TdhZW1OcBb
e4MBslNRgK2jwfIRvUroy1z6wfheAiU7kBvRYu/gWLsLptJm0JDlmApD7A9dGLEh
YimGp+VZtxYSyl+c/ctqax3fUBXfGYiMga2VaVPR6E+f2+ymttKwse5jZPcY/EEF
uT/8w2SdJjnlK84OZQ+HdpM0fZ/vyaFr+V46LlqEU16orskQ8gI3rbDuoDo7Bwa/
MMYrBhRw0HQ1LwGmz3uwQOh2gLZexxC9h+hzfPetKHiWrMd4Km96AiZoTK5b8CJU
Aes2n79vdFx0n00RLdh1X7Gl/llxAwSAsIpt7BNkBbHdZhWc+HcdZdnwxK2TkEDi
RRu3IYBoErfAgM/EnZ0pNjMYQNQCHqP/ofkAWPE0Njmch/KshJRrLnweWAxvr4HQ
in/23sEu5EPXpQ7vWSGFzDpAJCwlgOki9m40zsKtIoEfjBj2s9pX49aNYbuLP1zN
RNIkx8fuXQfC7kNChOhiqT4fW9ufb+SPqf21OAxWtLNyIpD8N/IyGsdAgGpN05Xl
jgDzs2ruoHLuPv/m09xZ/wa1MemCgjXAUuRHMSdXoEweIOsCyfJ1BGqhW5F3fl8z
roUJ+8/CsOJgBBdjiM+dgwk4oqp6Y0/Q474466cv4OGPiASIAGM7bBupLZ6DdzJx
QlPggoppINOLwSNZUkIkGYRbJKUCpbbXHmVipmyObq2K/v94b0a5LYBUC44tBCO8
gyvxreAS5OqutgXAMT5+JsJGRXskRV6Fa6GOrRDioSe5yEiaYLaAW4UkYVHiBYqD
Ab4NULvGsZljL0HTlGNx59zsQAlg9qRr0GY53F2XngposLA/NXfQG3xl03phh9nW
5S/EFunWQtCWmV7hQtqHKiG7ld1PI2gEQPcHUUeOEgMzUOKOMvI1dZfEcWRLkK7E
4QwttRdOxVzyt7+G/cZ0fThujBlHkxZZ6qqzWCAafWhxGCIF8XNRbu1tTnlr38lO
2cxToBcFR7zmeD9Cj1ZrprQgrHiH/+LBhFbCDYlDwZpVK11fsu/PVwtzwR/n85U0
qjmAGxgo3qCrFNZr+VO+uGDx2+aOCvIpwsDDb+rrLt50BdxAGmrC9AGbgWbmkF19
dPLCIC9FCydnuEJpXsXRdr714wnl8CdVZ1rOo3I6ly+GIgEuiFDTvhE8B4FJkvnu
cmTQzMT6Wci+jv2aSSZxa0O3pfn074xlEgXL2hduKyjlGzsmXOqPdEHCIfyj47+b
xdZBRRMN7LlHMiPjf5ZxNjKK7MivR5iFBJZx9+o58Hu1w1fZJWSlWiTbNLADAI5j
BHzMsLRjj46817Rz9u/MlAjhCdFetrbs7GLzmJLQxPStyqRj6Y31vl+z4yz7vNt0
lTHTLByQn3f1ksiTjqVnEH9Ye9Atj45bqxgteEHNvYfgZIBp4x4X2/eKn69hWIfE
OTfZg2do2YGBBUcLF/P10GeUxGYFavVKN1O0jUltTWnQ/eebAIUoggCQvPsezMxW
yDt2MBh3Ya1Gl4ckeDqav2mpRtWVbu5cpJbiKd/1xuA3UndfOvU3ZgfpepoNz7/E
AV5dH6UkdqwMAn6IdsQmgzDL8fKEdoZSOH8pkfae9Xv4wN7YKMOHq/5LmwD9Qzm7
JnaIuOuKtLyg18hnCrs9bZW7lwlPW+L1+F8NKmMSsilqO6By3vwllvq9fijAWxxR
MhP/Z0+jbl/FMC+xMqtclantCCTyqZKjCQaTkG46EHpP8mSOZYbdlT9lSHbfndlb
iEVNWXovxkQV4h+vo+h41bDhWIGUuc28kyOW7s6bgLbnfZXXRS+ILwtaRw5ilg5z
NOAxtFoSm3WNB5m8LZhQwjBqn1Lkok7d/s/MVSCxbyKBYk99FN8leDk4/XviS8vg
lOP2VCZjoaWzbteMHXd37XLBEjO2H5b5CZ8OQ5XCZeGlifxLumbfDwVEp6TJCz8d
vvKnXi5MPsR0t6/ZTGvUnqxd0CAX7PuwdcVHN/VjYaCRCJwFyjB1JmjWgXufnK/w
QT4BwvfNpTzKAT4GQcQwv1TRo6AbqeTCaxiOXYXnhfG/Mxfpauv9MEVO6avfur4c
TYowB6ZN197ZJPT5vyRrenrXRzZfZiAjWkUkb0HreRiHgiy7t1GUyE/D9DKlwHm6
VlGNHukWCq2NKYEb4pJBL1yrei9qjcrBIbZxI0qMgyp92wdFGSN6b/lvqrxaZ0mO
k59LppeJywnjZZxFqH0VWnCdb0XvsEfec9XnIOj7gpES0JLIJxbQFM1VM5whY75l
HnFHwO0fdg8FVBbK76Dcyp5eAZXZ/zd5BuC51xmyuRuUFiQXddxrOz1PypPvhL94
QEpGC76xy4rn3lZbkfy30rz9R6aTzPMZALl9SJHTDAL2S6BjeIM+XO87CDrsllx0
A7auod/5L4oIIY2Q6w9rox9Bf+kVhAXPxaSxyY7Dc+fLn4pnqZ1t/KB8H1ZyYFBC
0BARf7Lcpxca2i5gQWUhl/U1dO1FoBlzfKU5PI7KJ/Nm3QhNHYXJRBoEt8ri6cnZ
PPOBsMyfwBHb1nKrLyzVPPahq11A2ZMN3ON+g+zRGehxqcB6pcSKCUQ9AP5CVKIc
OiIRlqL6OyL3PJ+/ZF+XrK8MTuLZuEDIGhX876yEmbXIRt3OvaX/3iOqadXaA7TR
0sdTHmDbIwSp34x545afdK2fPqR5g9/FNhdxKswVVmfLKYFewibmLn6jOW52xYH4
TBqSpkBezYwQX4uhb/9FGtrpsEcyWcm2FohiWtBldUel1hOQiaHEwVOcMLRYGVac
srkMhMScBrwXgY4kOFVMGCWvp+hTT4feSPBhJr2vqQz8/GE/2x+ZczevBurJawEa
VthyOhSOuqsbDSCoe6mpNVQbYdUqefg3Xx8s137oY3k2LO8b94xVln2j74wG9fFN
2k9WQ7jKu+5NoKtj5pKbHlZDFErr3alnt2nhBwrmGrpTbNyHuw6zEYuHNtIKLG1B
R0yUo1AXKJi44OjRV78FTDrRvSg94iOBxhRv0UIEENHm4HyRfq4Ps9urE9yJgtL8
HOsy0wmfxh8Bocho+f15yENd9odczWUt3C4ZS/O4RFs6h+adLo+T7X1X8AiLM376
czPFL9JbakxIyXDHc6/a5S4BKzoZmwKVl4stlW7EDpRJXmJiZOaM9P42YEsrxViL
vqZAiLl8tn3MS90AiXeacMKBukUkA+bJN2uNi/LxWu+U8fdHGSIo7H42irRAcgyG
Kt3CyBGwW2DWTUJClsUxuNNhkpurpU0lhVHtqoGcxgF544IRDYVSfOXwKMSnQ4gY
kYeedFJBxK/c6Hr8OINIoIffBr+hMEV6yEK07iAeNUG1Q6T9mmAPTvj8/wr0CLf+
Y54WlIC9pYbaYYgqXwtBUnIzLX7w/eg3DqLKogAk56c3h9Cov3j2zkew2DnKosaL
Z20Uh5RxEWBXfNUDhL7xEE6AZgmFV08zFEEJ8EXcUy7UK/ohBAVFI6Nl4YF//h2/
gMffOBnXQOOegJe4cSBNSM4fn8tWdbASvpCspFxLwa4he89FiTff+vpCJzb0UvkO
gBfzagoQOvxKXmT9hV9Wcce1FPKrtgSLhQ9lvBf56aTd2Y19PnKiBFMWSAsqP5+F
g9OwRj9taeThxhWfGZmwMkwNirgedNWlPJuVW1/lHomoGSUPJW0TZCUlVzFviL6o
xbOUzbWk2JzLfOsU3O/DV/Ip80lBTWJlaH1Jtlv51fe8XQrtcF+o81QvbRIWzm3c
WH5unibGWgdgdy1o/Bwdh7nXwqfCMzz9JTAcBcCFxSODtzMqmYoqcUDIG7MF06C0
t2YHJY4Q7GNTP7ni62XE0wEvQbSc0FZb7oPJ+lAaRAsay64mw5XV1rZpHe67OyDZ
Vco6LKfZYyaPS7nts7JzzcRt0buVnEPVcJHG1EMT8wNyLGHustls3n2m/9igE0xF
zQNbuaKGikgysKtqDp/49LZefgvbZOrPI8LyhjmsRLUFpadSQtMC8szAMQwJmwOi
5nCTIuQcBAsf2u4bvCqR/Si4LFxgflXbZWAXdZ/Tm50ildYDPoaxeox/Pq+XzSck
Nvm9PxCVR+Pu0O1rxTdfhbBKKohgS5gIUZPo8qxfB3n+jJ6HadvaMvtmYV/uVdUg
IVPbn4XulUn0A/WTIuJ4PEIcQpkGAjyXhgzDVC3R3okt7TIQws7X95Yw6wLuOdrl
NyCGGPiwDt4PtijVMf8zuVmaubaa0U4MKihLtBZxXSaQorYt7Zg6gPfhSaBHoGbq
2+wxkEiSAexxMwO6Ideq5OODI0yRxRDsfIDzDAJu0NG0md2SH1amVqgZ08qEp3Z2
vKYmmogBSY/ZwJE/PymD7O1SNMMmM75qNQ8k/JqZ1gRhd0FNshZrPXHCaLK7IHOP
oNC//nmDvQV18SwfWdvLzD35wBuDsUcw7ST05E+RUsu6Z5UUQ+3xTRAnqNtGjdGM
NgfC0RGOgXP5eBpDVgXjfViC5LJ3XFesCFMXPehGEg840DAMp9tWEyDAmQztm+De
HPmHk/76oGvcL8o0rsFagWyvRCVYhpQUHA6xoeIlah4mo4Xy/A9YhYzMlKJayDst
oQTpfg7lfpeRXuAweOx9DL0kpCxKU8+LjZy0Z/Qwa2mb9zYwDUcgpF3xAXRA2t8k
upXC4vjkou/iqX4/WxAbj2/sRXUVg8AJkhbFz5aalhRveilNOASwiqzsZX+dcJf4
OQ66QohlPfiDECBIZyNrrAr6R495279trjNOkWSASDmFOX+DeZVtyVul2O7iOT5o
HkDjT6Fg/o1dZVqc6WTnwbHrgH/kdQ8yiXdkhga1+uRBSHsq5WoQIgquXw/kjBbi
nQwi3MXtymo+I3DW5GxPD1WbC7efA1HpuwrLGFtF5rk2wFj6AoLLZpyE8bMWzyLD
N5bwSJv2OYqunqIsywz5HTr5o5t+R9u0paA4C5EXpiv9fqy+Nem1ZNx3RRNfGt8J
8aH0evCfel2J2MeG9OOLuSbcMtdEnDG9KQfgrxVwBQoshIKCSi2T1i715gj1r1YT
HVxLJWvwFOdHPZmDdkf2NtjQ/NRAkG+hdEI6mS/4houqNmSdwIUqQ6DXep7Fx9BG
/SYIMIVwmV+XrdzzLLcOrh0XDgTK7WGfnRKAMv1mbDoBypW2ZY2wcnjG6N0cck7t
Lw5TJfaofnyRQFwcF1h6iACLKaaMRe0GAD3XJ3H0lO0WMMEhqG72xyOvVUAp6hC/
SvduT43bA72Gt3oYBrUI+Lru3FRgjZ1HI4Mw0rpUdTXtlx9G1MYNGVKB0VDzxOrx
MCPBNuFm0hyZvbi9cFtjEeToL7yGvw707DBPPSutWqFGwcIc/1pJH5GQqK1ZvHPO
hM7KtVcecdGlghCgxQZhNhpDygu3Xoq6xul6V30cK+JI0r0vGzglx0ijPJW/Hs0J
bPx92wmUbx5CB+mdKJzHmIOc3FekskHDI2qN0eCtiUwB7zEMVysHuBBJ/2xEo17f
GlMMe02dfLpmj7lGrMVra0UryX0yiQdo05XnwHIgoE7UqFDPzRVhi1YDgAIgzi9d
08BrIiPUXzk/Nxk7Jl/a2yQCCbqr3TGF5TYqHfvQyGaKl60EmyeBm50hZaNQU/gk
Z0HxRUS2MnCFYe/cpJegsSn/nQxnL4l80DG5GYz8byn3jqgnlst/3SqN8uHz//B6
Ni0B1R2NuCYTntaRU+poJkY+mZjLDc6rkQZ/lXTovkfCg7mrM/jI199bX0IWRetb
xHjFB5Md3tYu033PiTEVSwxD6U7vOFundu/dB97a9itP+g81y3Mud3pY37lZNBwv
ZrMc3K6NzfwFFfye5yzuTqc1lPaNgG1Xpt6Fg7wnrc+KsSv7cbUzFl/XGNIXJzUv
uspc0+8ZUPntyzOTEIL/EM+/N4byh4+KOPwnr8o5iR5dZSncAGpdAYSe6ByFkEuy
AYhTm5H9sG7yLcZZVaJRLVH4zUfgYgSv7eCf5SHF/M1SnAOrzIuppE38kG9Pudwy
MGeRiRIgA+yVMdCqEvacAFxcqdUABzUaRkIVjXEjGR8LM7idt+57BQ7yXl7BFd1A
aFmooQRj927tIdg4qal1yIq8GEBU6LksY1sLYZdoe/GQrcksDxyDGnBkjThe4une
u2Qz7chJ9DCMiZoUdrWmmjO9lS67ib4wkmhO44yHJ16EZdU06sTp8uLihqbrEfW+
UH4jknV7KPCzN2J7be0LC6tI62p68sE3ZYJsy32pYQG9UhOayrdwVMns2K3Q64nA
FzQBLTSnNRnH1KsZvipf87rmgXcPukDDbJt3c1AOTQXD77Thv8RfjK/yEiLH2S4i
RJ3c74Q1yjqRGqERS6PvJHZN0573qzz9uU8JjE4kFoxCvNF/+83ioSRoyBrDkJMG
vCpSxjKi70go+xSEBvIzEuKpAzEFKqEIU+jfl2wMWTr6Mr1+jCxJqfW//LyNvenA
1oP3zMIYdu1Sxn/yzrHOw20w7kRoVB7wDI7xw9NhGdLgAe7c4GMz5VWKIaUDwGYM
JYGkse3aGUuwQ5Ej54dGF4UkhkRpRKBG6I1BicyRa6abkP5FZg2Is4s6zoRUDA15
mIY4cwISC3yDnOMUg/RW+7i9xvz2ahbjHC+ThvVYvbq2B9Tn6cR/1O+q7EVJecmK
zvw7/f8YcLGh3A+/PyU0uciXszUyD587yyS1gzRXdl32WnKmLjkfk13S6VM4X5kM
6C3pzWYUCqCPHB4lb4h+/FcQKCuKu5Bg8O++nVDZpyNe5UPXSOTTM7rj17iTcP97
xZgvmGjvUUoO02N8fOfgOO+hmLUX7y36t2PSP17offihyFJ2x1GdUamI9R9u6yN7
p5NCbgcLvSn9Tx+ZtNSsbOeBxDR0gwguKm+LzrbZHr86FiFN7CutvPzLqC8+IZJQ
jiVQZeHmTBscOk0p2h0U0Bhp9ANbz07ZIGy7DSzioQ2VyR2Lw5+mZRwtADrQ+YR3
h6wuQ8twj0jNKaN0QRgoySvQfE7JrjStj5tap0xt6WIcWyqmiBZDYLXSh3NHkkuB
hAzsyIYsz6BbVUNke6GUuO449FmkgHBW25J6RbBdgzjqZnUWJxs0f3kPW17nleRD
AHJd3SHsF4MD5amk3OCfLHpmtwj0hbQXhwtkkPSwRGRYYVJAu3yqzsJTHhWOc7wf
ceTmVkCIF8dgan/p/NtaJbeVVR6fqK5pg2HQhlzrS/fxd9zHTljp0VpAAMUj2KAp
Ly6HRnbQiPCCjvJkYOHJOkvLBvV+VPYC/k4MLgcf/757bwUyPl4fSxvmSTzCZZc8
JOrudj9qE/SRoOJ3LP0tK/pDAaJpqONxv3pYvzKlBqvG0RsC1adJw/Nkmy5xvaTx
4QstI3+iCR9Ce14PBfRxL8XQn4TQoC7HxBUZjnNZaV4oYQ8POseqemND6KDDyW8I
GYqleWaHgM8v5TbenlN9RAmnAP+d4pchAZrB8FEXEZl6L6dkGao/05NZ3/RfTT7+
QR/gbhd01ncppqM4nrjk3X46KwDd8gugJBKmWWMJmosfzE6hrCSDsnViCRiQnjUV
9rLRkAjPStxjQS9d+B07cSfkGGsV3WQNM9YVMQ4yGREVycxLSzf9hqHwvsrUmZ1q
Eq3fh3U0DbcIDCnT3YVM6/DGxW0wVAyOhhpzbTKe0hwjoJnlIs9k2x0Z5mJ/xqX6
xbfw/pv25w9Roqn4pxua7kMjr+7DB5Np93grc0ni41YHLuPwhXixU1BrIr54EWDE
qfPXHiQVpIoSpg19NrzPno06TzTN+V2kxLSxrrI4VzjrAIALHvGMWnBJRegN7+fq
vXOSyA9UcqJDsMT1hwWbiqqvdkuDA8/372WgelU2vZU1UjWhETWOqUIG4sj3KYXy
v2lr9MZZE+JS7xCVlekUmV40fR2VXwvIYtHvg7ffF1/rnfzXT0gFDzIO43wyn9bn
1uHTekOcgQaNNp8W4kJAQB9NT/qr2wdGMZf+bAPcddhJCXZuyXZV6sALUZOoXt/R
20eyJJ1zNreE52QPDHz0adwsGgfz+8dlFuVFXj9nC4XslrvYrDDBaIjQd7XeY0mE
JT2SWgm/gFS/5fWd0ae6SMZzqVjr/pzK3NSucf5pH/gmajP5UO8EUrGhVEar+lsk
Yc69aOiO5LWmzn3WlXR+bKIRu32PJMV9UYp/eVwH61b5UJayfuz0qikTPpyvutVB
0NuT3WjYa91nnIPU+JeBWl9l3/DE+KzYxQyqzCsM0dCqPQrr4OQiygAMyoblMaCD
dZH6z0uEDzohSDmdBq6rbCBTCq1iZR+4XosS3lvlLxruWFLRoc3T5vdfI+2JN5CP
sauBCWRUuYUV+Xa4kneDmrYmOWQvoX81CEcYaoIY6LxTmvwcIZ8GODCIfMJF19Ns
Od7jFtYmuPvU9+8O36t4JLq4vnAD6EKCeqixCFL0MjHevbE+EJ0Nqp8/fceShMZi
Y7oKAho9L8hRpZTPRkO9EkhYSTylxYhM/gig4hQ6uc5aFV3w4iVtiyA7B8UvAQHH
D8q0PgXSLsEi01q3S6S87Ib6bSMYpc3ReiqXPt1AkoIAc3XKDRGV0Pm3CsHXKRt4
vsi3Xh17qMCSOhkz6XZ1j/uPAQVn5vzdOBRTo6PxNaBHoHAIkll0Qy6hRW03HMJA
ov/65Lc+nYL53AVKv1R23NJb9L25kDejMJuYAYQcyuA2BWEurAr9yQ7X+TC0kjWj
2p/suk+teK2qCxHYNv6qULWoEfGa7gk+0vmTuFi7wzzhLVNmIS03T3ox75Ih6ISI
xG3UsUc0WoDrCxJbtQRpwDj4Cx6sc6oMMFM6D78U06G0aqoGupjtCahWJ1QBmf9n
BKMVga32XHbO0/V9089vAkE3ha2c8xcrZsoCHy8yNEhhH52aWJt6ddOwgQdwwXVQ
QPYoTuZCLEK7tmRTLpuzf+0SZdn/dw/S/xuiOOiIFM2jNBBgJAxIdjpp3G9UycDn
ahRLuu3Kwp89oLlpqq2LnTmon3OwYKL2JJZWbkic5r/sPrL6cXa94GlhUpKCh/MH
YYF2VGa0fWrjQDNXemssu7aCc42Z/LOMgYIPcEkPlZggm4dA3TbZX0jloEZFIbUF
N2xrmYcESVzX61dM/Rkwa3DLA8IFM/w3W2YPHGBnZ/e2FRN+mFuD0oCLKY1WfiHP
++NDeoxOm5ju0yuHwXSQ+Q7u/BgkLOXEBLpWAevUX+ZfHvhKoqs/kXvOiy/PCp4e
+kBceF9eAliusUYROicAiOca8hzXH4rxImJlmghueumv4k5RtGleVU5xyBGvDRrd
z+R+AgQFtUmlUlL1Gj3nGy5OOO27uU7N4lPIbYXhA/Ori3CBloIYEX1ngzivmPZq
gAoao3ALjrCsu2qRufMFFokid4os9XQYpdwoKjWNJLLLTEfdvOQM5xsf6cyx9UHu
MFvFW9TbXlbdTwdEE0HuyR6IOlALFqObF/F+uatXDGepivDmkCI6Ed+fmULzhUUQ
UP+/J56uxdvWWQx9cznNOG7yLGfhZV0MiDICKRqHwMjqWY6fzAQ7dnVxNQVTT9Yt
SRJJV2AMb2z8L5wi2Bs9HTAz8e0adABTR8MAYHkLpSXcOmU3LHm6RylxN0ikMpD0
IihdoWRnt8az70D9EMSNGEeycKK5f1+aFk1u+1uHs/XT9hmYDloRhBQu5LRcJbKY
BbB50cqQFTLW4dtjHW4ccz1XL9LO5XLuoetS+3bPL5E/s2NlzUpFnPrMtZXydiYv
NTod2UWreh5bZGmfrzgP9lBNHLZy8JetQklADTvH24j96Pzxz8lJvBupEn2V//vo
B15dkJbYYSbpZa54LWglF31iJdaeO380rbG0MToPK2a9xMGRwtucaFkggpgotLRj
0MCMGF7zG3uWBLAjWYlGcJVzVYSIvPL0nNL/8EIQD3Yc6Qi9cD6he232TC1p4XeL
/9netys56as0B5wA28GJzqJekkFeEbKj/68xs4Ur7DLJHIAEhSPFH4PR6YtFin0A
KO86RAd5x9Tov8UyHOmdOJj87v5EfbsZCSEvH8gOuVrgXEdWYoiuTaU3fofkzVCJ
BPaasY78auBYaEpSGOXJg1V8PFQwd5e8cCsXkfRgMl4gAgNVDM1m6sBYBQcVNnPY
0m+uEpb1/krHwW9KMlmUdFFGrk26eC2sCnOJZPdCGdHeLCA7f0Q/7Gwot1xYHoaj
u/zkS6XIPgvicEMeq/MbsLIxwrtc3jKFf0LeHpj4wuL60kf9wXX8ka7PsHc4wzv2
1SOl69Eb3raHD3uYhOsQ3/miIngnCjvpURJpFh4g4Tf294SC6V1SkB0baUF+TVcm
Niitvg2EjobOFAgP6ghggyH7+ZNKI2ZGeLqe1G6eotIGMj3q2KMk/v7vkUroO/hk
jxP4d2lL1jpG1jXpEueWThOfweX22cQcU4S0oPewKaY9fiaJuvhbKOjxf/qk3SIA
FF4WKgalXo5O8hRDVNZSMLjRtrtVKJCen5Ac1Yt3dnRi9VLiP7/6bPED21lwQC00
ebOmlBpVyBYIJOYyWuDA5SOqGjynczHiH9wGMioDFkG72M6V6wu0hRUCT5XjDREX
nf9Dq7dC/rrFIRR9rygjhma7czSPgb72f8zTPDGBCFXflAP1K/Y8SHfLHKiRp8sP
lD29tDbzTBzrtl11ddAsVxTPqc9e8vTdKuDWiKTCc/ky61zcjLLL0f3TBPn9Q+zA
JSAmwkIwNA3N7y+7jqjS/P8Iy4TH57/H3nKwfNv88b7SOkw1BnS0ACt7knjHxdei
NvlLXV2gmplFqjL0DLfKLLCqqyPiY6XdH4Fo+3mHPP0b5DCd17KUDNVsCzHU/mre
ojE84DLdlvHWMY75CQTVGBtRV1c2zrl11gz0J3GGnn1MZGLbN7hSPwhpm9uTiPjy
C4CtMYvU/lmnCb5V2Jn4Qk/V0+pTujMd7qKbGFmwTkuEaoUlzLXl8uQWb4S2z/xc
vAmoTwCxG/ZLU/5OoB8a0FmRI7u1nLA60LDyqE3CwaHsvLlYKWecCGNwJZgLrtDH
atM5ccWEFZcRXHFs1GuQb0+fVRC6BLaIr9V443+ble/GGuaGMOcv8ImUoGxPmpVV
oHUa+ulMExAFC7/dWmLik3bVXADhQCZii0kJR7s0HLtH6pAf37EeRw7mJHhhF0EY
Eaq/aF7xzN9ymA2UEOudKRwJMg1KL4QXMJfkL/iP8ii/5YB8xhbYOXMjMjKmrXqa
Kdja/91/OkYqx5lfv4uDiSqkZF4HnKlaW4TX5YLnUDwNk53PzS2Umst0sPwOLqa8
bp209y7QFT1moYISeRUSR8IFv+mGEC7MhVGSeC97VKfXu75wa+ugD9B6/LtEQKls
lTDjuyNZOvvNZlD+TVzwdQ8cSm+5lv0Rvw3u2qGCaTZSzTTogTb/t5RiaGGLsRn0
+3WC/H27GZaF2uTxtOWuoWZVToL6APYs3NokDzUwFyRew0XDTWmlGTPyifr7BvVT
1BzpHer85fTAo0ccv/9K/J5sDjAR+JgQcG8fxw3/LuIlH7JtYBPmULZivLfVn2Gb
JPL0YP92nFjCNRMX8X6HOinzraMNzqDKRViIuD/IS1qMLJvBGwPN04ktWpDfVcM0
kwvZTJ4c4shN5Rb3S7AuA7gEMfxAHbFNrYdyLhhS9b1UW58RT5Tslm1WfjxG2MwF
pe3/VkfSkGrCuJkkBbxe5JsM/y9IRN72DvQWWdQYPX4NPliBqAzG7fhKTsYXNSR6
uBWdKNRmNjSYZQSEw1DjYcfT56koRUIGpVpFe6HjRgbCKZ4TxEHLzXH7NzFVq5EM
iBCUsiXFK5vMOreXWV739Oj++KczPSgPGpO6RxMJK5s/XGBExv0ovvbSjv8SQMrK
3Ok5AzM7ywKWY8FPlVzfbYuIaX7PY6jSlqP/mS/tQzkguCxY13hoxACdK7a4CcAK
oBvt/YKpQrtGz/f35+nHH95ZpISHDe+2cz+QbEcFVj6Tq6dqsnazk6gcLUE7FDTJ
EeWaC3DvQGh5Cfe+Kef+GlqaySeFLECA7z0iplkeQMeF8jOGZtDGHOh6TuX0tBtt
0YQPL/tOfFuJONFqeCi71TJL455F1rQe7bxI9ZKX1ES2EIyxsmN6nBtkbcx61UNq
L9H9jNy100UrI3PETcFtuoN5WZE15cNZGxPuW3Is4uRQQqkXXvWMpJ+GXI2ifTY6
VW0bnuO49ajD9PM/fxZk3cWIddRsOC9nHJblu7D7SAlnwkv6oJu30CBzgVpUpRm8
H6U6ev5tdmruJ+jrE/kecyGJ/qSK+ZIhy35A1RQAhfkMgi8g23bXso0q3uM+ej11
hM1DAZSv0VsZvahAjXpYK8y29py9oCQ/oAuvzseYCWVo7QQLBNXuLx1gcWXZLGIy
y3I8xSE0qXJz2lK/lOwvShyDlAdAvZr3rZRSVRT+cAkPPf13m5SHgNBxFXCZ6Mal
XKH/gL5GRcSm3GH+R1yf9I1Ub7Vy8V3Y12iXAlok+sJ2suPycab6E/RZHrZeFhC4
NXYrOA2apxGyaaSax9rlDm/5LpNoiFuJReRpGRPhRrTKz/WgiWUEhW3xu1fbLcS/
1ggsR5ny5NBWYT7O/3Sz5QbQUqp2/4VIaiBT83M0b3fKFoliyUaRzdqWeUdSrgf3
NNe1juhhx24BYidFdo5fJBUkLDhFJnnmlYFftT4tJVC+JW84RPFxWS7WTfRu/KTP
cIUZpTY+f5s3y7kHsFfRDRh8elMyQrgxwP/Zma5QtALeG2zx49TrQEPcVsBWx75F
purrMSfrtgPIwV5pR6i758ByTd/l74BYWdZ9oHYdp0dF+IerD2HNHkktOVHg4wcO
SFtSmLWsOk3HgeYBibCxXpYRhu+P7LxFlbZ1ycCJQbzlaqEZ3CbdCG9Ppsn1dzt5
X4ByuwOIpr0mG/O+USmirLZ3LqwhUlIbpjhigHe5A7vOOeEJW26098zHC3AhVN4y
uEBRirkkXuMt9OseIwdXT17Mp36j3lIkF7/JpoqN/EI+JmIyUbUNEnssoKmq9oeG
f2RnfPYO3t5vpF0LPY7ujw4TSDMuEZI0WBxxJZsV+aZ4zSXadSE4+BzTssi+SwqM
iKIQW+txLP7ccFSebxrBni02UZ+nLGRl9lBL/em8xurTBYB3zzXwoFpFIbLbhR8u
U4lAP1jlL3v/AFl2cIViNDWiXzZm70LHHYn68AQTJMXYQ8I0zU+eU2URikZJdMbl
Y0bj1ODsJYdvJHh0494jJ9rGpN0F3ZNse1nj2L0JFMlCYohrYuEbIUPMkqSD1m5L
X14U9G/4h5EiFw7Wlcx6o5oPEb/bMp/a7gB9BqEsF2L7f2O/3C+S3F1QjZU4on5s
wfhG9wWmoX2YG89SCq7N71MRho4rV+MG7HVeRYBm5WnKSA8SKf+MeYoBQu8d9WGv
ueH8sVnwavRdsontvxr0+tl4VEf92ehW87m5wyXyc4HwzKblXVuIcG4fcqOVDTlA
lN7ACSmAabTZZEwSk9bGpijoDhLc3+N6foaLqriouyxa8u2RDKp+gohjuDA0aQOY
VbGPtBLmOfp7HKZ3XYD0krKybdm4SrdP6sqRdEfhfR+K4ioUym2Q5xOtMJKN00b6
yIeksevP9Kxk0lb2M9CG1BFuMpPWvayYGwLMsG7Ojx+nxtWDFOglrKDkREeKRKdG
H9q09+i98b7T7oNRh1xVXkuBbl+fWkuZq9mGyB4jp1ATUxL+x6RlsdWj+nr8qeKy
V1GrqauE+sFjD9gocfRAc23XlEw7tvLMXMar7Db/st+AO6S37oGhwuH4Om78WikQ
fFQwblXgb1xS2WLbdj8j+PbzmoKaVU/IwtlGftzNZVBLK/kJOme/amrdzSxyDj+B
OJH1UUIPg36KQORYBrIqPlJu40wRNiWhd1kR5mx67c+GOWTNi0ozvBYm+6HCHmGc
1PZY4tf9qIj03zy2U5+wKbMDZnpeg31iDZF87B4DGnBW7rON2wsZC83y2POwwHXO
e/wDeymkTBAGICa5R+b4EWFx8C0VM+696B0cq4l1QN1I8m4OkrMod6UBpbhEJlEA
f39aOFjMqOtzRBKcpi7HyrGb+R5DZnLRjptWCxmyeag923VbYmOlQUSTEhHOnacA
Q+TBRlWURtc7LY0nakQDHtgzZMdhPKjF2j7imeyOcJINWXFCSF5o3cUaCEn2WUMM
GQSAYuOb/+VvZmnjm5uD5f1K+Sv8G3m8ZXemZE2GHujiXloS29PSR3OV5rc45861
GA+wDj2hMHmWLaOdWGvF6LBYbanqq+lEyJfoVMRGcB2RRw8gGmB2C85YPuQ30FiJ
bgzEZ136wLGx8Bo3ERvmoLnu9h5u6Ma8lnUq/DYSmfiP8ulDsBLrAMJDDiZmS3CA
lz5/vcisAWFnLhf9nshcB7vnDjZ+C19vuTUfek/5teqUAMJRZwho8NAvPM0a6RA2
AK9EnYt4Vtz28EZoj49XWcs9moVnPoBnkC1ns7kIH/GlaA+VmjbNBzTMDyMnyc+S
vqn3uVptl60cmwQ+AO+WriJsRYT4+3xps+m0t+AeK3o6LYUtzPAIoKxHCQqruamh
ylcCR4wQjLA1ljCM6d7dlBFky3U7ODobZBkJAzUKpXS8UiGC0wY8RUh7c0uqFakl
hYORGn9Cg1dUzAlFTOTryRGJ68qVu75xgVcOV35Sme2h2uWi9RGm5P8AcAXBeZ8L
+HHZRxgEj6/7ZXZfe6QhlU7ridYTU5h/YjvpNChFXdC4gKa3FKiLVFE11kSRfrY+
Jmk+ZJXdK5ViVpCVXODRV0k10iZxrFSYn3OjVp3Z5heI8UxXvwZS2VxstpPhDyhC
JMoXUZomxhbQBabDTreMj+GOqtbz1g+Uc3XZ89Ee1/CPAicSOYrnzeaVIKkBGkH3
otPCXX2Yd/pVlVDNp42qd1nUQYEDqdFg78RO2ZJJW2bZGs4X+tYcPFyHyk4HTLEP
m/zhq252/nVf/v9EoGt77L4alKz55pSMGB8hF1Qqji44xV/mpSjvlJG318P/sDer
LYS8WBCPcICUssF63Y10uboY3596bj2/XUrfOAwZmZPyMJT/a6p9xaYyZiJkFBZw
UQ/tv38lEy45z/DffxsQvRx6cVyCMu7JIUpLvldZPCyyYN4WKnZrMWfImYd+o4EW
fYAEEaOzvaIvDt46Oblos+8uiSBqFmdqr9YhNLP1rZ5jXG0jL2/mlr4O7GBMKGu0
iHN7JlEBOoMX7Xf88zwMZLUJC18hNCim/OOIRkR7VQ2JJBlDTqmdowZKEU3OYHVH
DgvLPxOpClrfI1gxbasg+dPwWTKSD4GofXi4kQZWQbie0xjywu5FBDpeW4yF1MkK
MqUtDhmeA6O9/FRWwgEvd+kjVVabvau1XgT7hlLOigxTyWXmeYch2CIBJQXBYH1x
cssqCpfwdMiIh56pJoEntAi9/T9uIsyXsxYMdM23nnnvKQjfNAr/FbQDQ8DRgtn/
WBd0d9bJPLkzi2xbxG3mBi+NUBWXVFyVfqaPL1Q3fG5Eachk6QTgZe5JbPrpE8Z2
IgwTk0dCDKYTBwsMhHWwErrIr2gpuLbSS7K/xqJuZfxsO/9Gkwy8p/2EJYwRuif1
j+Tm/6355aTAFIZ3Mo8DfNqwhzSVus1iZGQt4R4TyR3kSgDrsABLw0oPNEBzh7/u
3VM1WzyaDfzg6DWsGeqFC9MNqFUf70NA+5lwta55ITMzSriNFjhIEfsge1Gs7SAd
Y8hxxw71+28JWznqB02l/EcHhVe47RJHb0NRoVWVGTYYga1sp4UcbTNusDcCSE7U
q+a/c4OpV/GmWjZBp6we5zMrEYR1NH0ryhQ11MzV4QqLPGZ3iJgQihwYgPNcgmDk
B+shN4KmtQXBQpT5/O2XgGW2Y3AnZjQJqGHpP5KqZJPQG2t4vZAWcTZtVoMuu8eK
T9Pnc5sqIZMpzHgaFQkkjCkcU76Q+EScZfuR0oAnzkc3ifsbkxfPuDteHy71jBuC
r25+PDe6DAUmIOwUc9oAvfuPiO4EhmJdKGGUzNUnwNGwCXKV5zyIffUOxpW5E4Dm
y3v997104nT/pRPKLK7RUZ+Im/fLKIYg8nGrmkDYrojM6Noj32P58YBOYTcqZX2j
J1LiEuJTnXB6XEoPh1MAYTOvXEnpUn5gQD3ghKY4ZH11493SuuZdK5AVYGhac/P4
ereyRpFZ71CmadeFxBFHISf7BAVR87G7Fcxss+Dm/bF9DQp6G1v1+fM06+Cz0VYH
aRCF0hHZOyH85XZFfuec1VKHZB32EW3PgElnvAG7Ba8WJyYacXRFO9JDEyHwSiCo
5jDW4NbMmTY6C5JFYAx7n4cXDUIDGI1Uu2Kmi7HdAuohSDzWu3etI9AsDqazAH7Q
/m+SCdk94c9VIjn6XYCeXWRZWtxROfVmNvXHhrkUgDd/rpTHHYBoJHE5oUDGCozd
gTUCXK6LglRAAh3rmh9Ici3XOSblg8EF4XB+Tdf+M9wvAjU8pi/viuOce/jvKKIb
Xli1r20iSVU9wMHyMVZqKb0I+gnGq+W43Jb0XA5ZqgtrkngHSFfJU3wROS8feilY
61aI19Xfq4vQ+OYkZ1KA/zWtY91o9w6Jjp+hTRU3EU76K7ZNcmARTRhKTkGRlZ1z
Ge38gKGETRwh/XnurOh8mPhBDCGIQGvOWJ5SNDAbGukDOr87irYOqXspKTn6j5n/
C8ZMLDSIRl6Fy3INsvD1LjJaapVNP8oYYb2dunH6bcFvMTA/PPjZy6Zm2JVCm19D
FRfbyMFqJm2OjuPVk2lWNTGXZDdOknDlkPISN3jXjFj2AtAYJYhxQFEtnc67He5Y
gIS+KRs+Dy2HdUX6USPd81Y91dZy4H/StuQl/Eny8q+HbSwvjY4AcAFktLMnZGxf
J/tHS5COuEe4zsSCn4e7bBdDe3WyKZ0zFCKX/5XU0N+6EkNSMfLdhIErz13L+BdL
9jUQ6W1lhC0IJrE65HzeabNtg5r+bBLYNKcTrhHHTyUlWySjmE8IYhbSPvQzgX8L
ZObqmdWUY7wVzQfpI5H1wTmU29Uyx6QZkFIdaDrxzhbDqOxQYSHKsUgk1c9v6Bgh
wuqKzcPrzuuKCbPsXjBcvfoe7rCxY3f6dCfut8jTCVB1sUhFfsUrj7Xs1N7of39G
0aBNN6GyDBjm71e18kr+LOJ48LXLvILJu/Pz6wE92NEaqbFUngSim3V0ZwGv/Gsb
Z0QgoNfCeTGKR93CPgsrGyYdx4xuSdI/JqQwxIn7gWeJuwFfoP//dgfFwZFFnbPK
1UbZz77ns34yBqNltN5LT75SBkTjZJXS2u8MllWhEc5p6lMLkwKsg+j9Rz/Ld0sd
wgYLrmKOan+vC9/69NIvOIeAp+N37HSU4XLgyToQu9P+J8m3uDAMRTK29xielEHR
zI2ig7+SY/nWaF3rVtlXeoPWC5nVkO3H+stD0aUwzC6kZ6dBsw4FOZx+3TO2+ST8
gIPe5w26UTeqS76Egq9FiE/2z2sTq8NfQjHVJo+MbYsBALgOHQFZNf6IEbS1n2hd
kgIxa2esqgRx2K7R7ApC/VmaVA6Fe2IelTt+2mvWJ+M9lTiDBpm0WiUAzxCeQjjH
L4D1xC0AgZM9FH/2oVKh5dg9CRAC4cWCZv3u9NJc/rQ9B7hjSvhpYdaNkGkB3pS/
U9kiHonNpaTdzC83vKp2O8Yj/zgtt3c6Mnu9dg7aljhkXIxtK2ZcQwCXEwY+YY+A
szm76SnsZCuFZQALJ/TCDfDowcPOadpV2zKV1cE5E6XdySa7k3QI7iaHnuPDBgF5
oK6tdf9Op4VLB77xZZ8z9agsv9a5g7siaP/kqNQuC+sYSKz8YPe+E+YgNB1fFDRV
R41LTooGCTETi1TJ1PUKHL9nAeLC31a6J1qK9j2KJC1IXIyslD0LJQfhDkh5rvIC
NeTuDTqj2YNANaBz9bN6Xj0dVFhMR1yED1IEuzXmSlJ5EzPffhoSODSxIXOJdVOF
uKWDfbadSG3gbf4M8wA3v73/50LaWdxpNi1N9kYcEi+gW/v8e7C5R/EQNktnOqUe
kB6lvyDmEw3pTmRnU2tjlIvLWFELbP0qdR/ywZIBkBgz0SfOApEhKcBe0cRxWt9/
NwkqsRiGZXqB1lpRUtji6OL06OmsgK2htgyNwr3N4LSVgoglJuErTZ9CnpMuBVUI
1XTGj8sMUevaXMHPQS8jLs6Wge/sxp5LzEzFd1/gkhMrznZA5pxNX2OlYxvUQeSp
iOcBJbxglvnc7QnQLzzFkKsMt6pCgDuG7hve4ex2GEK94abPCpwVAHbkxepcjsbt
MfHrbAZ0WPGOrkEidmHoAxzN+vCbcIzoRgVtCxJYT+bewoS+zZxnJqi5uMRdypBi
URI0zwf0S0VaFJ5jTjyKknztZxbp/Bs9GBW9EqvjeQbn/rEmTg5Riu7SVH1/61LR
zjjrtIElDxnvw/Iv3GReJV2buzcEpM4D5PBrdKWk51/psLYcwf/oqSM3BnoIpqLh
bMribBikUYNwwIFxnyF54WTLtXId2MWBMZ7Dd7HVnF4Z3Tj0Pcr9d0woxAu7nPkG
qS9OKi7xhJyh0Mk3Ckkjro+i8oIyb6c5m2P+JBiOuEL8V0vRx9hlnsjyuUBJ7dEL
GDizsheT+4B9Qp7HgypBY077Rhb1JM29tiRbUuQkz6H9bIBz1uto9BDypbu3vXdl
GOLbFYu8RReEgjYsP0IB4eDuxEJmivSDW/GMeSivRjlLW4r34g3gg8VnyURJzoQa
Jf9PN3QOe8q29qvyiEx2nEsGgBnvLMLy72gewLO2HnJv+vd8jeZNbKSX0efQxwD6
8TRRgkbxtWsYGeh2CQ64tMFnghDgv4fflhiMDe0u1rXeo2iJj62ZlXOeqKyifBkU
v29tWMTapvEwhsOzl1x+9kddms5yGRXfLRHxxB1iCEUFtbtWA0ekxOZW6GM7DehR
IMKFtudCohRsziDaYBZBMSab53kM4oAQUsFZpMgg3s8d6PP2RAtbTjBzWnsUm4+R
RkKaBxsTQ0ZFU97vr+cr3E9dOuyJxY8Qng2b61Y7UfcOrd6CIXwX/YIYqmm3UzNp
Bul1nNDLbJKUG2GxFZp1ynBslIGx0ixCFxCqlnHY6G4RbGn1SpNF3Q6XWgDjMElP
iv4TXqjWuH+Mi7GXkFYp202yR48PhqYsUbxEdOkkC9f0pfUsntT8oGqp1216H3UH
w5B6sC2dQprgjbQsjs1WsBLUhVPmMmLd0WULWkaIVZgy8JWfE4mKgderdMQsM4xn
zn4MM3SmgjBAcZHJoqBqE4wNOWBZyJVfnuK0RldEYitQTWLuvwNaaWdiusr84h1B
CaNpD+O9OLFRPdpc1Xir7FRYsS7//V3wBhCdV8v93Zk555kSMXdP7ghLgykqW3go
blQV2JxG4q2fyjs/qsbBeT0lF4rAtbA6EWIXvSgjfRJxC1zM9y8RrOb+GwVTR/Gq
7PuFnESjKH+mOP2hFKrvAWO8+Lx/dDn9G/Nk2ucx1K1y19rpUoHC+p6w9by2ClL5
uC+HhtDKdcPKtirFycRRNA2QyF6Qg7ATvdXzbskt6EfP1iKMBdaKgD5A1oBr16bM
wfjJDuvsUR6QyKns19VCjjT2abDZhLcTkF7VQO7GWvpFKwRsra2BjVmK1+n7Okh7
Ghy5rm9QEwpVKPptSfWaGPfGffGRqe7IsUEv/T+xxJ7YK5rRRp0n6UewCvIYCOAX
vCZIJnzk8VvgnYcoNMMzkzC/NFfs9HYSUsHzTiBBoADXT738HmL8lQOZkoZrL0iS
Wkw3wkY/UokQm8VIWBMdWcPGwTtvjWONmLoetRybeGJ7vMgimrOO5351eTJjgkI/
huX+hRXsK/bHwszkLM9BuUvgHh3C8A9r1tEc/65dXfr0KXvbO9xFJ63YtX4nsn65
KBpQG9rA7OWzUS6AKhxSG8Qd7yJXQqnXO6z3/ydL/4J6/K5Mbm4JywyHeaUKSv8K
+LJY14VUtAfn8uDpsJo2MhnD5uMWJ7rO5cwLDwboGYr69/iTcV74b1nbRP3J3R4e
E3qLH0zMaBpZbKuCqHtLdngPqsDDWLg3XlaZbuWnQ/QLZkXDwpNmaiI+s10nAnNu
yPnhcR1iiXk5OYxjDVQ9+tvcrt/ihH4KT5okZVIhWxHYhHSCoF244VASBlBLVZjl
axrXMzMSDIxczdxEDUtADL55eEK24HcHtZpW+bdaU3WjbwuJdYw5EC8U5BzF5YyH
SLnsInLVATEF2xCb6No7AnwQBEZ01zrb79FjBsJZlRbbPg6cmjzYDbb7drMjjfVU
lM4yrXUXCxyAv3u1bK09BUT5JMpHtYVyB8+OBb7i/8BCCEYrs5czYgu+huVmdA+q
ecDPiMJ9KvoZpwKnXv5Vd+y6/lLovxQYqA3ZmHhw4RKBfam7qEdTfn18oPW4hdtL
pEDAsa48qWla3NoYIWKVMnOKosWBZCisfoT+5K6UThT50lW0SnN/hWNTRivyEor9
+6qsvLpV0ld/OGcgaaFsWGwsOu/Dpi2wu2pvli4uuH0LmiCMYZ1YMtrvu4J78RZD
ucuqSt8UkxviRI0M08v6dKuWHZmFKNFACd687F33LmdT3XNWHhCgf7lauDliFKDB
K989pia64Lq89UW1CY/cWWhxflOQvw7bYvBYcqmbm4Qrr92Pzi+Md8WG+cPAUYHW
P3sf51fCEVMke1xjnKRy78XuTkHRyn9w1mQkQ+X0A2RNqVNX+VEEPw+NdGfSH6xY
kgA0zbgmLN1SuTAw343+MoZZnR44MoE+VIx5jn/3WqVx/dljhBWc2HM54skD9T0v
xDsdjwB3vl/IwUQabBq2O1tNDNWoW3UP5HTbYZk2f6HP0HNQdiR7g34tVq4onMi+
IKtqTbTRiVpSWVowIE6FZMGl3M/prbmDtcWmDTr/bH7oOEKNDel2kC6H/0iW4OEp
UWMJngWGAcS5hyv5pE7yngrtvWjGh5DzMj9AT4M4vlF7IrWrpzIzfCaFkLPlk0cH
hfpGDxopL3qN86jnVku6TnbWETeciE6hkn4sTS6APHpkFn8Fh5pq3gXff2W8PWKQ
QZ53JjAzLhdSa9tp80GPkcFSHk7POCtaJzNYmdGJmOCzmW6FinbS7TqKMScyssFZ
6WSVag+mTR67t/dqnwg4A377kbZTkJk3KCpxuuT3NirGBwqLro/V1t20AgaFLB0p
20CzoLM9opglITl9PZnxy75DjTDoazNkmbd7v4OtZ9gt4Y/s2SdjkSRqHpQRIIHO
C67AisEjFl5HNOHApedxJLnHFKkxiv9BuqjQmmG67AO9IBfLIUFTedeHAbrtvaKT
uRns8Zteah0kwASPYnrq2WI9/tPMq+rLjGD2cDYl1ExdArnQocnQ6HylArbnRXT0
q1N4pCuycNqgBnBkBDRf+rVq4IP3tYUVwLgAUK/yLM2FUpXcnzVYdbC3u5D1dZZw
TRKZD0nl3iE0QHGRrdMTzyUwuVCDEv3tM/FGRKPlikUsYtafYjwdurQSlIiKcqw1
qGx6K1Tjln/JA7fTlod0lAMPc4xK0KmwXofzXb1nInWoDKSYJ/z0Z50peJf6T2Lj
aH5C82mtwLdMDsHC7l5jU5e5Swr+lfWuAeF2mxNRVyUa64gHeJ/PJgPJ9GDZkFwX
SOwYA4Z6Uom1kGVeBGMZTCPkHLxJkFdA45iYy6agiMnoWveMasSkHcZ85bOFJeJj
2e9ZlIASG+RZH2kol+864d2GdNMeHMH8Fg08LPLZdhrEbVj9mYRf9GN2Q0ZR+2pS
6eEITPT4978hDVaZ/6mEwDcr9Ql/TMkBeSvIqEM4QZpBCWeVqanHXG/J4iWYeNSp
2w3WtzSHbi9ItdK+cW2DxTJkQJcnmVev6B1GhfVjkzBCql3bN5rQA23ABIL+6TvP
nqG9ILw+NMtR8c2hI8zg4DGHfkPl1bQHyfrjzfZMiFmh32vaoWdF+9qc8LFYHKjX
aX8Kx8OjJ+LO+I0Gwokbl+14mzP0Jer4rmDAAD00O4rDyCtvDr0dRApmwLwoLfT6
uEIlIrB0vitiX9SbEXzTrXGqEnEyByHSzuTSUS9Lwi77paHOUvPVX+D/0fG91lh0
+5WIdulTdqyU8szxlOV2B8crxKTJBGIPg7LEt5fIkq5ox3Sdaapv08FzlLh0qIrW
0WRsWchWslnZODn9jKSeCfpu00MCizQpIVc5UfIQgfqAv9dQqGBdW+e4bDd/qfIw
RYYn49fx2yAMBbrKuuQcIMiayRRd+wl2viYyDPmt7YjgcqzmXODXpnGch9VY3xQL
tSpVSXNaAW+GFnqCGA4RfM1sikEMEDv9SIbLlYO3TMly2aY2yQR+ZnEc59l+Zgl7
8TGAXwxSezGCFsBPe6zyc8VmWZzaSW/95ew0MtsTHWgyJv54hROshKFwKiGOPOj8
SR00FU37IySIxVrixSt3IEqNoCcIIblACx2YcYnWsuu39uz1cfwkJ1ev/fvBzDbj
0DvyjtYJiMLMVq1H4LKKS4UGXP7U4rPKwGTmKte1pOsAgIjRoFyh/7xmF+yl031N
wk5ZGQRa6Q99lzkZooPH+90MzdyZN3BpqYvunKb8S5uwjHkA9940YRGgwIXlJC+f
vV5yLwXyKZWTe0h0A29Fa9xb7QQ3Dpj6Fun3qWCT0J7+6yo6/mNoBCKegKdPZNVD
dmoLwi15hWxd7gKuSK0gB5rSQjbjowSO84Lza5UVijYAq5VeGTuvHNYkHWJadKW6
5Ib8Y9layLxqL9jyeSxWKP1ggJTDylqfyY0beDgKySbxjqALXiOS8Dr7+lePlt2n
A91U01BVvO+fXAMQZOj4PBJ3IoX4I/GYuZkn8Ftz9myDMB8IDepSvIwYWfMT0WuK
/HzUuPazMLKvKY97DLQ/VDqwS3NsWb+XMp6/Ge564/Jo7KE6er7lC7DMS3VX440e
VDyIrkJzxp8MWzgUUujZR63RaeVNyhTMK8As9g26AoNgJAH7btvtHJRFbTcRlWWW
4eO4z9u/PY9A3+7tmbeBaaOdBUMdR8eTEeME7+nzW3Pp2Y3f/XAWbbcOyafgk+x5
ee9Exz0nyjtiN0FR3T30msNFzogNIDHLOTAVR6QNMNZPd9K7HFPMxrXOBmrhByH+
REvKsoA8WcfrT+a9Z9xcZLKkF4J06huBAB1VyT4OdeGd8d2MYDcw1s1YzLGcTvKv
21XvRPJrNZIyKulc3FFFt5Mou/d2JduTcTq4l1zP1f9P51hCeT8B+ksf5QiMRJyY
/nzA5qjaICeFf1AUmTQzuoGwTmkpHScSxS1ZvBZ/qe9DrfhekxUMh6wtC/6bLxCy
ZWc3DF9srx1/zu+uIsAACU668qvzVthz1D0mW7QO+XJEwlkbghbrMubiRr3OiLA2
0lQcYcZfE4N7tjxBho63pE4yA0ZxXcReKbmeZLS15pomkdhjlHMvF3qGVo5694xE
FC/jT4X2X75pH3eBduC6/B30bDIeE+dBoErsq+vIXxVwUSDjDksHvb3Ba5iZj1P8
n6Pu5NmrSpPyJPGfXkWOzMvfUzTbtOCRbi0fZmBHJzPgI5m/+SNyfrnzcXueUGQl
aC+CxUUsXbQ7iBqa5IIU/BlZIkDOOsOiFbLZKnssaaCuLuyzGHIg2+NViivYqGTZ
vQ+biKerl+XZTjNTK7UNHyH/kCC9ZSZj/9/vzolVC82vuuEPVRqw5zVT4jhcWvYV
kS9PrysBh4DRpG4L8prtKIY7wpgANfe5QWQPFwQuZS9b8UXtht/jfajIXqxwPCJm
oQf9l/Lxz78BVMzxfuCrYlnRQm7lV4DFyBLQtEpSMIUtiYJMis7JXq4JlkK30WJk
B7GH6Hgy69vBGqt536GOJkwQKU4xJ4yzBl0cg+NM+mMU7y5vBcjCNCDmexUfoL/9
hsMugC+yT6FBtJMMX/GBOmnbZx0nt/yIxot1fqZroGr8TP20pyZ7XE8BzN3Fck6s
ua4N35zu250jq55A2M/+Noz90xwOT/SUWKZMK15bGlyx04BeAngs1zAJwASyT9YD
ZvpnzGEiNWnf8DRQkRJyjvRHMwORq4y8cHh7NP9w252p80yVlTGCpZzNulYJSx5j
69/gCvh6btitD+cPHb4rktp0JVuwX/NJvY788TjrTNXTEkxOUUiqnJInCqQkRoTV
mbgsxFp0SvSUkJ1qMEYbl4S0Q8Etm7aQZ5yXk0f37HpWSYevct5NXDCss005yrO1
TuRgbfrDEO4zyrPKDw7RVtIrTx+oSwvEhL5v70B7Aq7jypoD41Z6kJyrfSHB00bn
X8Dg/nR3V96xVCjR7Tyu3fu4U6f5BNYaq6/rAM4VnATGWcxCwbqLFjXNLJaoRZlw
oFwq+PeGE22J5a6hB6IGwS51lnQn0QZ9bZWDcNCaItyhl4u/wbF2Q1rJIc9ctO3J
Tsi38VJbluDNkVeaZixhubuzhPBtC9+8d+QB1rCjgrslzdJGYgu3AaMMw6Ho6vQ6
uB2ZEinsEMjq6uDrK3zDEn9fDFxjK/tG0+QePzqIbG5mK4szhvLNx2JQNpDD1/Hx
lv+KNQN6jQX9jCa6I5ZVAy3T3gOKUWFlTTfFXvMIifvAoqCcB5LO8rM60WXgfTp5
h+IYiPTxstrkFfFDiHz4gmR1kCaxLpuvRmrYIjbBhkQWHmXJVhMVagrJYiwVUOf1
Y1W7O/O0LwglIabqjVuDbEJIHrYjxb1eCw7kJ4ZTidXjkVeUB92H14VFjd44L+Du
K6REjPFwOO9A2uEJF6If9Z9OIqddoTHHjpbkSHG2N1ov4z/irNBW2YfMhf5Fz47e
+PmM0Kft/pwjXfVWMnjF2E64Eq5BnUE7RbMkq8eZrfguNPwy/PKwHDSjKDY4G2UV
4GXpSt6Bu9s7c083HSWg9dk/RV1Ki0NmabIPAnuxO2Z7zgjWZDS2TsIXlDk1tqPa
TFp66oJo2LLFc0eDeqPuA/D9idzxmZoNDXUzaO2ekbXJXIBE6Xizgue1qc+QHOOT
OmGa2TSU7riFCTMPQ028I1xknIJyFMJaMnEPfZwgH5oXLle/rd6pQIQEoAuiM+oh
yDwaeQb2lfPNbaT6I6pi7rnLofHT8DpeqhoT5Q+kwEU/Iku9LccgR/Kom1usPHW2
lxhgRwOhS9L8KStw1/CuQl6sFwxjfS1PTaRJQSdy1gtEg2VG7lbSO7YnDDrOM7Tb
YbwFOTZqq3j/Y47dBGP4aXk+KJhni+dJsMgfkFjw1jRUHHYR/z/qBGdjrlV9flqN
UHtpGnj5bX4t0qdICJk8Z8gtLJO0rPtIok/wiutKDVysk8bUz3PC/nTZCByi8t52
usqnJmPblhDFSw+wyfUVCq35cXTt1Zbo418taIZWxf2+UXyeBmXkbzzwgthcQUej
NrTbgLJWiue8/vl8MWsS3dkfV3u/NuK+mGZlYLKsGBoMb3m6POX9sVpGT7b9k6jD
vrtgaUFHL4DLtVxZFhZo83/4wsSoiOfmvw/JSMIXm7FIarkCE4P2z+JuS2r2q8oZ
0TTkQ/8fUnkfGjzSJ+UGVzq4V590DlGnODv170bXDHR4Fc2vMkAIBmTsVXKD4Xsw
p1E+D5UYHkFcVCYdflE+goxc7Wws0GHNpCXz+X75LO949cls/+1tQmHsXGvHILal
eJyzFOnCzikszSHiRKwVk4A53EJN7Y+qyK4oC0bFQca0sJK1aMUG2gNY4/uSF/kt
txJQ8tfqLG4Q5ZE5azRRX/CkZ/RWR6PaD13Ku3IgTKn0ymKd2oWIdkSJzSQacszg
tWOYHqPzCMuWCHOyUsOlpJrPyDXLLq9x+uUGxqyFF+CR5YgYEeUnZCEmuENcy7i8
ZWnm775jCnr5krSbcxyAcq3YFg7FIx2kR4cjqs3JtnSLUsDYyS0KFlKLyWNF3uKV
nwbyI99iwbpW3c6ZsCHNeGo0Rdq30tQ8KQfGPOqrlg2343WqZvJqF6RYz+A6QMyY
6JrgQ197qLT0im2wNr7PAvznF+2cxxa3jwX2OJo2HCSZ79Ykdkwk5eg1V+Obg6tE
RFulYagG2nzxq6UTKBBy5SxLz3FZe+iVPftG0+Vc4L2y53rUMHxBr8XlU3Gh+pOe
a/1r6dLQj3w2vyk/KKjAE8I65WT52evdDCu5ATF1tEAPWZo/lOqe6uyAhfrXwygk
wRRNNYLcHyqhJywZmnLX83tAd7Ef4YBOx24lR8h2kV8HmbHLjBPBOs2zif+7VzLe
ckzvsF5BeJUEv4pjDv6XMO6Ly859BoNkY397vnxxN9fjnSyfRtrtNLJKBF1THbTE
8cIhjC/9O0j3CwB4DCMcw88GoSzVxb5D40r0w46Wd7utTZasbkU73bArzQUfi9OL
Gjx6NRvH/BKexOtBEqNpq0zV9wdAwMAE/EJ2xJajHcJuBSv1mEebHumCMQFIuHTO
kOR4QMWcMMQ44+01QK6BhM6tiphJ8tBJ3Kw2Xt9aHIMuVDyRlI5aLE6JHg9yul9Z
KKF05Briwvy06FSqL57Vm+/arCbymbQG6EGaNw6di/XManGbMn/KskngYhKWiCNa
yq6C7afoXRO+WK3rJHipIN9Ex6ZRe7Iut8kvwTEsp3IV08JFsPJVGtIbDhBAFBBM
dVN2z3HAkxq8CBvHg52f2EQ8Hl7vzJxV97hxOB3n872XEfX5+d+3USvtKkCaMRtm
pV/mCwMUr0EiW5NWZ6Ceks4O5AHmdosAxleKB3JRKGPmKfkGmbY8gFxVMEFyUiXI
aaGykGoClhxQUh+nNgMCJbzPAodUIr+L/4QsC73HkVK2hj3si7XP30zfq8bDcj3e
Uv7Z4DRb3v86JP8e9uZaPqJV8QacPdXW6lRRqMlD+gjwPcgTd9p3uLS/df8JziKa
fYVVVa10nuZODAUGDk15xAJpdyKjZKuAvU1/Ib+ZCdDpENZaS43ik1j/cJQw2rVY
H8wFm2poQCpCFSvMEy6baVgIHHUoetM9Kghf91oqjnPpyuR1jtu1lhsYcO+qyOCk
lBwRlR2/8mq6DsFsDCqwX+jBJQX0EMaLC48mogsSfGXQPSM2BBJz6sr4kcYpGqe5
3I2A6FrdOk+V9KIImyksJoR2cxASI28LY+CbHcjwKYYjaFV6quDWUtYyMvQSQbST
D8nt0iPMEx+Zn4NBqiXFV4prOu+FY4h6l6u82aax2J2gq8ESeV22x+grvySpVojP
OgBlNI687Y83nnQeyauk/XnKC2nqnQYcZ/S+ta/krNDSdaYhAhE0CabT943R5D7m
MIdjDhOraqrjmexjScqE6ldyC/OmyE7Y03q4ygTzBjzECh7e0RevzHr1+YsJvZ/Q
5xWiCwsMpPHVImGSkqYM+Y3yUooTFsFZPumj8HDlmILzcSlbqgi0++5b5EIv/4n4
9htzp2bAZVDmhsV0TNpYwPxqwZ00v7HjHJbhwYZkEukL2r+DB7jRfSTc9uBGlhPC
tupSHzvJBwxw8u/662v8WK32HhVNe2c2XLWYFSrpB/lxUk1BSrHRGgoc/vbh65DO
/DbZaznyrFmZwyKwRmiXI8EeE8eb+l1yoFP5jsPJ1avR9vruy50BRAuTJvgJCy23
16Pd4IFF68ZDiOx+glIR/+21R8ffG3NT14WtoqhFgXzI1WCXkHu1hpwxDDpdzdk7
j9JHKwoHBBkposdLygQzFdMu/TJk0Pn/H6PU4yP2YueGA8tGUiwk9pRMt64EV7Yc
i+HNYtEnQGquD4ynyuBmwAqGAlXP+BCux1saPpy0oaGtwQW5pTWCT/yWcmcyqcFA
kUBjCDzskS+FxNA6c51VkvNMQh5wLcYoA64c78ocz/ns4JVYXB5CtVJNHH5l11R2
hZYURC+GydfL+hZVcSLNjZSY4ZCod+V7tTkHuM7jX2r0HC+viwTbQZ9mT77wHV+9
B1/uCLP8xnxI24n9nOra7k4T7OcTxzFS13Ntw/83eu8s8qOUyk6mmLDpOp5i0gpE
+Ymz3M1rqNzq2+5/x3bxadg/abvFVJSgwXLs4BuwghG71rvZGVRr1ytlQg6jTKXy
2yP2O5060SZNnEcrmROAz1EyjNMvA0si+SFndV+jXWf3y+mtL761tnDFWXvG0L8C
idsAlOTHJGwaDDvYh98MoOMGUK1mKiQLqAUSNyWPFmKY4BjOdcxdfRvNFxB3io2b
rhRpTTAsY59rB33NtlEkl4+utvWAkIMS2gTQdErf7xNbCCiDqsl9vVkcBBTMRCCm
vrP5CdjpBglpUoNJuYGoNzZB6x+PzCixJNf8GN99NsYjOU4L0yfHpHdcsotz3a4J
bi2CP61/WBnW/HGHglW+OfZ2JicaxCc5OVPnTh9Sd5UJ8o0h5jvgmIkCwFjPtXQJ
6pVqNaLG8w6gF0BG5mezpmp0+Lzv6QSQgJJuPTtRnlJ7JzDXcZKkSqf7Qq4cbEiT
GeivuNTq+T6V3Mc6B70M9eQNjEf/OtwoDgzpQKQZ1e12/qd0YV9p4dgvuDenq2Tu
Dh4lkmJCxmjHvqjB7ObuwpoE0BWIkej7CkT7iqQHvNEbP94xdWe+VKRZBy7oAtAk
xvteYJDUeJnrUX0UsmQ+RuyPhBMC/LBa6zwVDVY4/zGVr2FkhhgeIO36/XL9EUcb
DNR2e5SEex+o6pzWPtM7yDSifzeonn+/y6PjbmPSzu1SVuzWEI47MX9RDVe9GicG
M9JsHEbcLRRCTe12jsc2ioQS86ZOzeZPd9pAKGrvezcOVpKHzyVuVGMTLtG3h8Is
1MTCToudYyqmHY5k0fSkcRKLkFYGGodqG6/FSRCJ2A/tjpTkSsKh543LfdWi6AU6
V2DuRJtvpt4Lad/kQ8EnW7HKefIjD1lPMvchJVeE5fxVkTySSbVERZXsL2q5Qp/v
oErDiTG+IIMt6gIOt3v/O3kgg3c4ziyciirEoS/TIcY24I5aDxR95nRhZDQ1MUud
VKz75S6osfbxzG8x7EvKfHTmpdGaoqmjPK88RSN1u+ZL1XT7ASyFMXnfotC2S88R
C6MilSFa244tXWYXi4/YObSe3STb5pDJ5VGp83jl/WOIM0vxXL+VLRlSyJzRaCax
nK4DiWywVbypmznMVwEDxDa/7hCtLuvg/TNoalcbF74fkwOHUpNkUeliE/ln+bYH
OSPDt9as214gKEKVO5M4ZIV6ky7pIEe6kRBedWKD9WWFkHaBDWbHtF0+TAchKGVP
B5KE59PgAY+2XW9cIZZ3QXg41rcfPDGGDzQnqyVxfC1YrYkyYUTtuHjyX+14Isec
l1eTr+/j3wHL8D6MyTpWcnfbs4kzrsbSt/yMUdlLA5aiiGOK0FTMRoRAAYSxOKpQ
RveKyib0r9UHYC01PT5KaTrwBFjDXxqXNrEBcIvBmj1AaDPAtdKpmE/+VD3w8d1r
w3QBHhkHxsoGXoXE3Vs5KKcvMqThObJhODxicToYcaz3Tax+dwZq1dLHfB49KhQi
WJRWmUfN5PlzI340XX/iZonmJUe0qFWQqBXVniEZAEgeOdWt6SbylvwGb75bTDA6
nVtygzY3TtShpR7ifvDkg2gk3F4ky6LYv1YezD2t0LARppYGMS2XoYgT7rlUgUk7
ANyFvkf6U9D6EoDjNn5M/gP3M6wNafgianu65NkVL2FwA0yJTQFrFJ3j0okYhfv5
UdIwpZgU62mtKof7lHCRFOyctz4tGfXBrVM05+/pjGNW2KYRKiqx+ZJEWd/pC57s
5RzQCI2JGueVxFMYbMzo3vBj4s///w/cQkVoHN+zRLuaVe3+zkpIdgb3V39wLJ29
k2RQlxQNv88UiEGPugMK3aFWIAibQuBSEulaULfrNy1tY1Zs2oNvWhPkNLKjuQOw
jN0UlWnpEN/w3P/3I+5V9nLyWmwdo+uI/E5+x+HQnqsR0CmwCSZ8wmAlV30vfhjL
S3v/Qg97Dl0lnHLyB5TeEObRnrkOf9uMw5rwxE6OfmHacuRnjGBxJpStLMLruHep
G7rp36Mn3yipRXlldLDXtH0q4s6QDcxy43ahnlbfaf0zaeK4K/4Licq6F87ixzly
Ur57zIBuBgjSCaWtJc1VDsYTDRfjLBlhjSSeI79mMeKshFGW8kYk4h54u/l3IclP
5tl1BKDbSLctDJ591tWtkTbmkCRyvFxGmwFjDaqN1Qw53UYiF8SV+OCJ32QKywJ2
M3mvZ8XQmd5wtIy/ebHtmMhu8VatgtO4dnfhbuwEDJ9Ym2PAsztFr/AerPmC9j7x
o5WtfHbBPA5Zt8o39/JH+qjPALXO4rHtRMu5RYlasIHNYL0sEA25IcYesiFQ91YP
3JheCdKJ6tTEtAvWjUQIeQoYABKKHKfqEOXHpbzH7gOPEpg5AFUZ0/AC0BOe7vzz
Y05MtEVnj6ndqcrAIMOjA7QYWTo/DQnRRpYLQRadtbeqAiPI1DNHltjWFt0yjDJj
pgcJ9lxyRjueyFfeJsIJZAEqHwXK++cj28QvPS1cWsZUuIlFQMdakIkzP4qNF2hn
ZDG2t5c8G1rBcqTmNJLnmY95XBNIGwpvyfSzr7BNNtybJNk3omJREX8+GfZk2aFB
cso7l5Qq+8vVbzNvSMAzuLutZEIcPgPe2Y+Roj2f1DYDZP7dE/QNCawCcZLkbBL7
U3PPZ+zuoGIehlicHk8wtzw6Ed/Iumw7Wc0nl+nNvzWbQCg6YiSeJCW9iOzlqoj7
U+yN9zlBz0Bedsb58VBRiQiGyevVA6/06mWM1baM9nf1YVFKwSw+jipvODWwdCTn
Knq1eV4mhTyC3zf3J7vFrLUCl+3ATIXZPha5GjIwG93bYqdJrZCwk2/v8GDnDBLi
F9po0+Qxv+kyNgsZSvnnPqsLenpBZYuI2nkNnsgMVmNRla8IA7tVH52cm3XF3psd
XIQ0xXJOh7AvIhVt1SpW/VdNiOOicMcDmV58Ty747wf/x9V19+4tYuswKJoaMvXE
F1ltIaUaOmFVl/l8KxB1axoW+UyX4qPno4bY58xkfsTEPXGeDGnuzh1L5vIaTfjK
yzQrJ2U9w9B/5N7+6QihHked+qZB44Gskg3vl6jNz3WZg2cBE/0Lz5R0V+SU6GnO
2u/Kn4Ns6Gel5uajnCkQOVkq8yqvVEx/28O6MeHtTVgFBTzpyC80yTJSaoIWJxLb
BMcOLk/DAD0D0FHlFlzeT2ZgNSoKKn3Dgyw8jwTYx8/TAtsvxycWixr9RPDEf+VG
jZY6H5a6GH3QykTWo8t62WcBIB9femloxZy7urRweiinUdcDTb/R2enhKfSUPhx8
poPnxQCzqHxouSJCSNRiitxt6h+89fr2IxNtkFpevIf3i++rkUEydF1xJG7yEDWp
VLfoYvQi5ZEjzhGHfhMXDVWoOcI0hcEAJwy0D6hL6KwY6q7Z0pegummOo2jsHq19
uMQx/COZnNR6RUDB8jPaNuqesxZKSdbAN9ffMLVfL26B+EH+9penLL0SfBmK7Aio
OwxFvUr95SD4xpMfenrn8xnH94c5yj3+YRJQw6xvOdIoy8miTDUsQaargPS6bHky
fTvjaEwG/dlK2uvOu+d5l+6hK39DTAsiTLLWsZe3ScpChilDrZglQGqN5BrPJUV7
4jqA1nC5X+O1tND3YmvKaz7jCc8n3fSvHUTrWAanuDSroET/UTP59pISLDv4GtXs
+3VYhpq2Jl/gu8pugXpXcgpjRFFNIlM/B+VMl7WgLxqTpwyyLY5F74nm4VhUPbok
gW2NhcdTef7/lGyFTA1joO/ZezoJlh4lgQCiUt04xL3FbWB4Vnml7yTxcWjD6h3e
f5fPISNQfU4/vNmCVZqTJ+gfmG4+gH7QojCWl8G+rLdf67KJlsPToSkg36Ofi3h1
skG2LSYbh2V5VTQ7xLvneKqK+rX4d5WuIgLjA4f0KQ+oxqI2y0sw8ULwvctHBWsC
lcgXYxVA9YlYFt/Ja2DEyo0NqQGR7EiLsWjMX9CZNUK3L6wZnFONhPU9GCUZgY5o
QcOmLTSJfeAIaRy5kOw6rchUACEbl7JbeCRDUainFAo7unniDVuyW9s9TlY8JyMx
JfUUYQYvIP9boQDzXfSwD/0UTDjO+1WcinWKcRrAkIGJs37kc9Uxemjeh+4aiETO
n+HTGAZK1pRj5a2KfQG4nJSJF5T1X77bsJi6ipEYv8B2aJqUt7W5Pdi75/tvfd9b
T8jpbgvonOjlcFGAFYkCXMKUQknbtCR+fMhU5AvqXJ0M03h/qAsPScoB+fKvofjW
j2ZkVr266E4UHskFT8BuiSUAOlOOJ5yuCMGse4Tf4xb0ArWVRk5oecIg0IyEDKym
ZqJqCCdIl0qfd1PWsJ5Q5Pblw5DuNMa2haPWtWL6BlevGCBxQa99RfR5V8z5Fczb
U8v9ki3gpx8JebPiL+jqFThqsYazlZ+bGsXlRWnV7Jt4EWKhF1m3HqYPD7b1Heo0
bywvrBr6h/h+guImiJE0ifoRhf3yHbM62naEKbWD7MqxCdioG9zCouOc1SRwBLnD
Cim03wsbOs3yUpcY4HkoQ03irVXMS+vjZkkXt+t37S+KUK/8j0NS7Vsdk2zeXnxp
hfA+MpCHAYuzKp8lgDrNDbUFT9863Gxz0UEaSvFvd3tzjp07SxWgOKZsXV+omJRm
QthwKkNEynOuqE+6Gd/eIB7jOHDoOvRNjB98WezRvtOOtjiFGjgEj6gc3oEjuH38
ktoNCCxnuR8bwP4jNwJILTrJ85/cBfXl7I+t8VNg/JG0jAjEjk1dHoDt0JxOOXzK
56SpD0xyFu1Vln57IlfAQMRxEThUxXoQK+ojdhqLBcQia0zDOpFKXDcPoETH0IfC
3URupGtHmvYWhLV6UMTXmjqczLFdHwKpKCPGxfAEOhUwbcsCBnvXrB0VGS0GL/ax
llFrNJzxHdRs8A6u4nG6AqEnutCrmfW9k9E3RwCXvF8jFpYyqy9MpqOIr5DITgBd
h2Ya0H5BhHSG5dlrgo4tfWd9Ja6cgpoxT9rWSswq0yT+6UoGcXbH0Ybv4h3cRMDA
e76clb98lUaZUN0a+I54aL3k7PV12KAb+rBG3EQTt1HhIHrf2z9Ie25sQM8RrS2i
fAumeGvAbvulylELlJ3d5aSynxnh8xfApcKO4mG87xUU8ouKNTgQ7jQy8VVq9jDU
dsEdLuJLHtFNxaG1kui94AeT8F+19eat7jefF08gohldqkIrWUhiyJy4tsc1kOoh
4S/zjL8Px9Kn4fAaP1asNN2j6lFRM30RLOu5XtZuEXCBP+zSQUTD6g/t4SgootNd
Yc15A2E7BPZV3wGgpJBEIp3TSdYjAKq3jWu1HebSjq+kEsO2lsLoR4wS+82QqCek
qmC1pOBWUFjkl9aZ+rd+2jeSRPPSqgBTVuwk9uBryQ6O4hjbvixbFiBimwbmEsXf
ro5Dmc9wldeXNESm8r6c3YP29BG8bl9LPFLQLl93vnK6zqEnuSONjDBmglRUh33+
trG1U76ZC1ocHtKOg7jnRplV88jBHX7SQ8iPZZYPIvz+zymnhiyFM+AWtCx/im9Y
20hFET98VyVt/olaNxQiZdBAYgPg43Nux1NS4Aw5V/lLrh3BPjMMYUzJgphaQJNz
C31DDSbC2jN8T+1DLlMVz4UOnYUZbnMqyIbq+Rg8t0Jjg0yeyX/TtQZ5o6vDnORs
AY6x3u00AazAKZjCZBLHwLyPtWdSDfGfZDBkhraNpAj5JYncJJ8YnUASfytnzzLV
MQDJ/EVGoemtFcBOacYjTjgQhSAdY+oskukCu/w+MxgBRCi1JnlYKGpVCLqYP+Fn
ywVybrk/OmsX/igmQZK5TlQqYf9Fmlh68e/btAS3NSJ3oPCzfX4mTw0DQ4oT+mDV
BLBuZ8Iu+D1fOK9U9RLzLgfU1qBxncF1/NwEMoH9wYErsTDW31x79beJUlA6sKfM
R/15WvpjLZmWaiP8jbVWzrM7NFJJMxSTkEaqV5gruYn+Oq8slzxi+1Q9MKQrZxEd
K2kg36bb/zeSD7ZxXwKSGsT0Lck5OlzK0YatMbijjS/sewVfLCs1O69ukMejdKxK
hy6CfUFIwbcaDCiUcg+LDwH3ouwE617YvOvn1cmNokThWgYR6vdROW44EdmziL0B
ZyH+skT8PlZ380juyRPRz+WeztvUaioUcnddZUdzbnYYX7lv0xz8n8LzdFNKWvVO
YohV7O1h0Qoi66aJprwldkkfSAMRToiFLmD3Id7UNqRVDYkyVEbhdBYgqvvs9VAa
EJbfTjicwuEZ+Jz5yjkb0xxHT14CCJ9PzjeATpR4EXNpr4fsn/O8B0WQ7FEcodHW
B+ka6UN6ZInjI9xekSylN5MzDdgCdfDhHHV7jTfuTCl1BLdLrie1dJwQ3TxdVBVs
OLsMMC1rercMKDMTA0h0JwW34qGSa9bj0ZNZ6UKSV1Sksa3emD50LcDUjmc4iXfW
k6OTaKfpjPbwOg+j5s5fDRGnnQSxn7IPtLWhVKLCLC64uHDhh+4fJ2Fwu9bPeR9F
doxvkxEG2jcgMULtlYfwB4BbklsXbhR3t8zxDeahC5iqm3By2eCs8FCu24UJ7BJi
F5SHYePfeP4LX9Jt7Bl3tRrkZz5GzD1xUHIPzNeAgNfp03E0VOlFCPc9GOHWjg6R
VHp3CPr1P1d0Jh9b7KlSdeg5x3CIHuETmQIJgIg2BSttrovGenq9icV13UbVUH2x
Yk7kusXV1jT2R+z2lz6cWW7vHtSPZ+hWW1czFc10nzRHqkx0Uf62CSZ+J3jmK0hO
vk+zxUoHJi34ywHLnpeplY6GmNrRRAFQHmIfSH3lNxyAU1Srrn0iic6SwIS9zHbA
j8ZevYXaCwQmQtypooHt0+S7V1G3rInNgFZ5Gx4tkPFFocb2xRQP6k66jXCuAJO/
gYIOQM11bx3W0eOewOFD5N8Va8x5fQcobfeDegLODcBUCTO687LOo1rdYlb+URQW
zZHcf8TjljBq37ptvBgEmWMkCSKP6xcFIIFPc7k2nGyMAXUqDtZyf/lw5GrtAfW9
EqxsVnDcL8oohhRzrY6RwkOWSAf5c7nOfEYGVKMf1NRCMoXlvE4/4YZ1+XvN9Pzr
O4zyq4sEI/8G/XvUioYwwPlm3rkhCVWnwRgLEozTP5Byl/Vz8z1/fihX0626P0mJ
Z3Hq8rBfINi4gi/exYtuTrviScaV5x5H9RTvBP4qw4LRTZQVa6gvtGI8MWq7wpy/
MA0pnDMJF28sz+kV7XuVPjZ3c9vNHtXzlXTDyIgrvEfzuabD09ILKw7UlVmo+tOK
AwFekSvtie07qw8CIn7dMfpuS2cuLgLB/FFJDLkVHh6hx3hvdxmnUdTJOAHwNTz8
EOsdNvcfmWYccKF/vlUoMT63xqpDEMzW82jgNw96uV00voZpXnmUGs8J9e5kP9nO
2ezYhWEcZ0b1Wtft3LARetx2cs/N3ZT3huQJmlZCxFv6FX5pZGZEJkJNFOl22VXC
Gb5vWBwLkfVMO5lEi0VryZoWASR+LgF8vv0wB4prgfVX50DHU1IO48eXwOEiASC8
2hvp0hOYkT+LjlbxZvDogTubZvCSgu2du2J9RyNqoS7IBHtFsr37ESYLDpHaSY8e
suevPFGeNuTR0mGdugbjolNFzsrHKDAdpRZ8HfhOCwoVhO15DoBnHFxo2Ey7zuSd
YFZAnnmr4k73RO5VsnvHgDqjWzRrujXXDyQ4OB3in5UoGWPRllRGpeTol4vJ7DIL
ZNwlbi5KKR2A6TaAbDFmiIxKgJNjdla/9QqnnMc61qZfNjcbq3EZmmqW5qIdENmW
874I9R0oK5M5PIz2v0q39oqLlb7jjG4Ti0Q74VjKKSE/PnVgAeEi2qSjyxYGYPMK
32KIoRB+xWcFhEffR6tCJYNiGyfIr85MDyMkiMD97yN24QYQf8ETnnr83R56FBkn
fGY3aDRqR/jQ6hDbwygpKcv3VVJXfdXI1ZEm0pp8OlsSdxoeNxcZuUgDhqn0w8o1
DLdIpx9mtqgOIGeSHtmFnLrOUO0ur6NDZYGl4Aj5NvYayztfvJ1IFeJr5wNpSJVV
GJaOt11t9+j0aKNQO3TmOH1ve4lDzlNv6w1EVkI2ShO8Jmkc/jVZYJFA+AcE4VdR
dn8VegDU3A3a5InK5q0KDyKKlis05W6ynE9LFGyh4Rg7aYjLAugengFoi1y3P7L5
6rs2fIKjRbUGFw5rm90Vt3HtH1/n+XCPLsXe4NYByhIXpJz7sXDzHCHT7qFa9Ino
BoGIfdGJKzr9kExwMRqR96mWImtaU76M04OSjERrM2xK9CsXAxYSAuewslKS8HEE
Og/0FFFjkZXXMF/Ob/7NIvSIwb6S8yjf/ZZso+5diZpuOZjw+qhzklmTyVX6gqMg
aTATU2Qmgg1ykIYEMTDDppyBild0TcBCnLqjTDzdSWsyAlbjtbF5J/B/yrtbpR50
408VI/NStZpLh+2krCaTEPCdd206cdS3YNq8UiBQ3kP3Bky68Z+d1cCEaLF9ADiX
aB8WRVR06t/wanBDMM3Jc7sI1N6Y1NnnUCakhwWjtllKxVemr/0zU2fotjCrPYev
VDOJevRetY5ddLEt15fPdPEcK863pzI5rTjb5RhQUkIKRpYKT8iEf6KqXcqsHYws
WLTKu2WI0r0YbA4Sc6TomsU0XkSyO/9pTDzYNGS6gf3IBIhsTAp8CN+RoMMM/kN9
c+Gz5/RoATsUD4wL8YrM+4hdAmXrPz/z/qPMLCh8/gW5QOLWAyra8lF1ktVoLZLH
2+3+aoJ/EIG7bvedKSKFdIPSQ3UTklrXENuLauFbHtNxAPNsPVYDcyLRP1iruyLw
9T8asHpOB57WEiD22xLYpTncEx7mWz+xRraFG3e6ipMEwfuU0nNgq+NcGneOlfjc
P0MimO3H7uqud/jAucxyIRyHraeSClqtNy3g5hHK+NTvXR6guJMBJKGihs5Ytb03
c5MaB7TZlMGPZs0p9CAaGSKAlg/wlmKNvARTNhqBOhfWl8Fa2mk/FfbJQ9cTrvL9
W57rLmi9CLXQByyG7eX6e7NC9QGC7HSPH3Bz2fO7cQ8ubZWowUI43yLnDUwTpf6Q
ImCluTK28CXFphPlMAJkm9ykQlAxN9PTlcP5sAV/HnR26m6xsOsZnPA+B+yvBUZ0
DTvDZMiml9oA1+TlJCfp0UE4QxNbMSjI95NifSwvo/BYWkgXHpjCIwUDHQvMeUAY
7f/Mc+v8KbQbpTcNZUF26k84Lvjl1k3JgvTtWAZxN99/pJ4/pGraSpiqPIBf7QwF
3QHhIl5CIV7L0EO4bZGFrnAj1qq/bAlNr6JJe4fI8BjB1+P1hMTJDx7LF714ALRM
ySW0pv0QL5VXL2DXxH/9xhDuoVAeuHFhgdIh/kmIBTHj6ImT0damrtwGxq5LDqh5
7JW9wn/NDALu2nZXf7oQeQbGop6YUXE3NPFa2qtLoQXQ3a9l5uvDy0M7HsKv370m
ef9GeembLfV/qCoOq4l2yX59iVMKGdGhz+hLwgOwAgaRiZ4/m9ZTbYzX8Phh5Hy2
wwbA6ipaqYR2oJzztcCQRuVAlqs3sCmf0f2i+hMiE8JfrPc25j2NXrpdLazQ945h
ip4bPg8uurKNsI+ml9Z7jDpCtYM/xtqXWZ/vOtOl28q10PpOewql71S3skuNHNBp
SZjYP7U4VsFSJCqAbT1DtkMZy9BpkXOTGjyQFoSsoEFtrhO9LGPe/50NP4ET4ZPE
6KBHHYr0RUwrpzGLlJuhURw0ukFNQ2Zq4Hi9dC5L0KDwWwJ3YY4D5NFmKhcihbFu
Mc372snOPNCv/Rs+Rl3Lml+dfUvMfSlMcgq0Q5O8bfjrx+rxTumjmMNGasr1sehr
si2lmpHkf6EnZCjNOdZMDKtMDHBO3TXHZACUoAZrWJoMANMufwh9Wh/wbBcvE5KW
dEfKWyhNBuyGVRxa757MzZW9nnjUVmvV+kqSy97VEJNPzIeqZct0B1wqWw5K4ye9
pHXruDKd32+ekiBR1IxLbjIeY9BFHDb8V0zBkxluCttzaeNapBXMbb3NTkWxv8E7
l6kH+ip8AMsAbJZnxA6CG8W7V2c/XYI7PEVaqzTfPkT1dxxtXilrpNq+Oees4OOI
/ZODhRQOEVHZ2/KYWNjnmbtfC3A8wzGjDWQCrGXSo76RT8gJRYtEbKNd3qiMPS2D
MXaHSpINFXkOW+V2VmoWlVQhrwf0WGDvd/nfE0FPSNAJKDBfehl925f0CgwVJB41
F9K8o14TB+aO3zBw5hE+sB0BH96aKQtYifh4pg2o8txY2xzyOH3YJFFeKSrI4rLx
RBQMwtDArAQNsnpeE8YoTwB8IGEP+jNvEB1AbTmc54AajmAob+mQJKJMf5mWLpau
9ixzOdE7VJ4/20KIo7N5uLogkjfi9a3eemoWszrXAmQi3yCPyaWXessUQneX5wiE
RvFfBSip0PChx+m9o58UbbldeQggzAHp/4uTMSC6TD357jx3UZEZHTv88Y8ogoqE
LqCtCYdPGOZ//FwcRHBNorX5MkDFFK6LeReDBlNBp6FJZv2+V/lwi7xK3gwJb+SD
cr2fSyupNqZcBQfO22cEMLf5Kgm/xVOgYcROP17m2GkAXPC8SlVc1GelO56IcIGB
u3YDggSZD8ryhqxXxCuecYbfGAfPDdCtM0U7AduzwJoIgd/cv2juZIHP7FPRjIb/
sd2ZfhoV84Vx0lmcfyGT8qHGQVWFgaYwmJgmClC3zp/3H8lpUPi6xsKfSmgFNxSh
EdNbRadoftweqjYcpEFmYNiZxwPZf+IBVkVKsFGX+nVkVuuaLHIrHoCKOzB9RN/q
g0yRSnjZYoJ6tLat88C23oF+IGGWOEqZrc+2CC+s8NR2vkYxc7NVCRdYRnkCKs/y
mZvZK+/S+JF3CZPIXzE/TlGqjMFx/gw/AuVziaiFSJIvQiNrhMsukVX8BuH0nLUX
Z4GZO9cmzcRyCQWvPsjxzIotdSZMTRLWjzofFcNQ2HsEx/0iyhc4x+yqL0VIE3un
HY1GJP8n/+YC+JRu8wscYFEqlwvJxYdkmfFmMzd8LlRPpL0qMLXyFyw2mb7wKOsk
0fno3lIO2v/TY5TsZ35DnA3FceZg6ZOSNEoMmTSq4ORpNaIYBoyvgHq3vHnQ2UAh
dRzBC2RvrKsV36PRAL9gX93GKqaRBlCuMSRxowuvkTlc+kzUuLIxK1Ix/j3Hf72n
uNK6eissyKfIkFkL0oSHlYFuiWpGsO19bdJIqyS8Y3IIZaYCHiOnnmy9ZxsNG6lU
zPDf2P/Fu7si7PkgnGLJ4P8C9v+XWyBPGwmdfntX+5DYZNXgrZ7wxKDTx3Y18Hge
QpPRXgwocFhoaj/ABFQuPQl730eKhzeMH/BcGGkwuZqGhbBx81fsbP/9LWuU+8Nm
iB26b8C+E9+UbyI58CmX4QvdGbVPhgV6c+5ViGrqMEiLHd+2HAZko5ZcunDB5LJN
B294ojarLO43TiJS4w5onYN2RgkRxS+ZBN4h708nDnWHG1y3u27Za8DeBJnGvsG3
1xaBl8oedFoposngXwWV6tKKPJ9Y13lkZDyyCgfjFBbyFUdjxalu+pXj54udz85K
58u1S+3QYIeo25gBTJp3hpIU+b4wtKDHzNRDl2wP747/wHBapLBwFS7I//XSJ6IK
+++2r9uAwCQqd4YG4UwsG3xXkcFTVZxdhqYeX2YOruN9KnmcXF0HMxESxbBuHOsG
zFMvH8aN2HwxbJPPA6ejI1vBPrkkeCHr6MX/C4a8DoeBOACjPL4j/eWaZCcdT9hQ
v7DFbDQvbPs4guBaJpf9MtK1YRyPlJmFTiJegt2KQcWk54D9trjlzNEZEcjMRSfT
MbkvsySy3lzpNvb37K8/vRGAXprhVjCWx63LxvagnAs8ODYhR86m4bzqD6nM/TxM
vMMZPeHvGbQONGAsjMET5tvTM3PT5hZthmhcXG6AJ5A3c2JikOQXN7K7YYKIF4Ra
n2kJTCF2r7CzXQ5A4eONUoQRyrnjLTXK0yVLhRGaVH3cHPPlLN1M35RuNnsXizN2
SvtFcZgl+XgTd7/EsGvVjd2lPXVNPLyQaM+Lk05yI4wREHgACodIatwFF5b4y+tR
tjnjSZ/HQiDh+/ET3PNHCSJ+7FRilpe0h812jkrWOKPzqWnpYtIyDvm+6cGn1s4s
GaFvhgzfBZblmMEH4MCLpGZV6n+nprc+lLYNtmXSbLpUXqWWpat1FqY+Kaz62u0G
iihwcJy3jDd6GhyGDWK5J49TOZC/vaFSEIlcbBfekP2zrWRtkm9vUXUX6fetRTRW
5QKJ9WvFM7db25uF9Q5fo0nU/WznKOxUw6ShJazPZDVKkyqV7yMcBHnmjd3m0BHC
aORhL5lAXoGZZH2OLjyMc6Ly92K41G+UXM4zuaQtP8/PE4/oV+tATnQMIkl6fWPH
O6p0ZrlnMtPSJnttmeMP8o32jmxxkcWsYqrYeJKEcoSukGjGEvnyleMazHISiV21
fc4B9MLV/P3QYPeJ8Pif8henYy0PChed44GBSpyiiZrkJMQ577TEewKytFyxGZ1P
rAzH5eV2O04Fdj5MVDHKXqTnNaQQ2nWdjo75kXnPidymmVs+lhk6GlBP8+1zZPem
e0egpNpLiPKfzyi4yNl5R9BhmopJGV4AW9OhKSgjVzWRC4HLnn2+vZKRwCuKTPCY
lNJG5obn24pOLZzpRssrCBZEqCr4P7u3BE+ZDKbGCN16pu7sEBQv/v8uqex6G4bR
3wuQRsYLZP/1KdO8lEMdt1KUksvlw9+xd+cA6QiTjBXRbRfnNJURCWerbDwsj77d
f8xPvT+rvG5lcTIKNV2wVK4GoW4PD4OZaupOMnXi73HpTYw7jWrQ4aFwtp40uVkE
wbCf3oqbljZ4kCY5JWb7fK9MxvKJ7C3cX+amLicU9lpXhSpn6cbfHo/c9G7TJf2F
Gkw9NpYNzxNE3MGJ9flyRPfTl4tKJV5JMb7xLI2weNdET+AhCs+hd/TPOV4vsB5/
SN+rEnOBhYVFOycpwwatA5KjMRZ2GCQjBZjVzi6HynZj7VnjSsAmBbxL+MnvxBkj
o4MKHzJY3mKSY0602VwsTYyBykJRU48U+1EnCIlWhiJDq9gFd8isZ4Am1NZwzHn/
uDuFK558qhQFusTEg104N8iVK4Rm+kcgOGi8F6CwB3pKlgsOygPfpWm1KaTg/ASQ
M72QJBEZEmlXUfbEIQV68IiawEgvqMIWsnVRfyLs8Ywie+vVH4du2JCI7LlaAIGo
ccIFdfEzTTfkhukhDtQyoBkPOaa0k1x7GHrU8fd4Vt9rGYu9D680OAVp7wAcbuAl
+mciqGaXSirGkZoAV6WBz4lnjs9py/+9gCXUidFNTG6O+Af11/5z27k1o1NHcioc
DHgjoyNMapQTR03O7EO8nlhtM5YYiUUsFeG8HuJhaUxw+7PqckyBViphE5TObau1
TQElLXlwG9lwxQt2DAmgy2nn2oXq3PSNNR1F+/xsCDhcetRGwpMq4d3odVErTChc
KKYChaCultkhKct4hcHWqGBZJTo4lnkkYXKBzRbf/gevxP2AOzSAcd1Q6JbdRDU6
KYM69/c/JmijXGoK2CMFnoGb3w7JZuWbQGIfnNsasBm6mo/Uwv1zs9+cPBj7hxCu
eC6XFlKhkZN4e6PnxiF4+vWrxXzw2uqmK9uel7XIMmy1XRVIjNY6CROX38WmJO9l
KdOVUqGfrLjYHobCyp50XKZh3d0v7MQ1ZhUSWsyNaY+EfYJJwr5aweeIb/ph9L8K
stj6CAWMIRlNdEBpJDNg7kSUxw/XorxWPZXZ/2xmt3d3KxSBZIiP9VF4PU85UybD
Zfc1oOd9rNPydzgYpHv9j6Gdz2ii+n/vMilMOHQNbjk/flwEoMzp8JvcbqI/g2cm
jOz/vRY3rDHy3wT3LCEekyfV9Cse+KSx2CgEsCFdSpSF4FMZ0TBsdHNHGEeFFzyq
iDdNZKh4I4+rK26SRrPLaoOs5Rn7oD4wpi+9/It+0ggZs2fO+xIrwpT4+wALGgLY
lGM+ZD9yY/qYRSiutbV2eQ78pz7pQ0Cq6o9G/pOOWYHTRmYz5KehkEzTTgtNGa85
olALIM60BqNLljY5Gar9nsWH90/dPEHVXCDveFrul8qnNAXibj85FgUWZZKw0O9u
vNvzDr1Xn1gaErR+aARjz5ejUreYxLrKPn+0QAuCFliJOR8FHYij09+KLaJiJsCG
s9EmRHKc891q8E8YmixSAMTfKFqsScRMfBgp03bmM5s6A44OsymyrjRhj5LmVU7k
QlHl3esOEGSQm7MXFVHLxXTeBDeFkB1QDSGxeErYSvf2DQniLAcor5vmKhgEqpk0
GUJEf263Xbtt+qfUavivW3ft4YIGzcsTeLmIFPvBfwKtTyGDe24Y14NnopBEtSYJ
XyBKSYlRK4gRA1fYJd4Anfz0VQ5ZwWPVSbyNBdgbrQbn8gvVIBdi9EjX+vHZ1Uau
e4QyC3DGX38abu1EiBbxaXuMmy/E6N8QC3IkHiDb2WOWPxJRQrpSNQcMXvrGNMgX
LLZyTFDBsJ5n1xG3flUR9MzceQZslFDW0IN7hRYzBJp6PBtzM24YtAeyPe9WF0Xo
vCsydIv+ilGYVANyoI2A9fyMzXkluDRY+cXsdsVcbzlHsajV6A+ATVWDOC7C+xdc
g3GHeZI+mJ6uHu07snHKcDwsE0kLRlTPzcPRrRejIhoCEjRbW92sHQJJ2SU594rJ
xHpABV+vfFmkAKtd57Boql9niGKgBHDYI6p5SsyuzEwdTRpZIW+isXWOEGJKSsLM
sK32gETlO0TxsTiegEnlJvc6GnrDVD4Nw0SlBXm81Zz0eyVioEVuFaASj19Imz1n
9+Q83MwSFdK3SiZzgpiQ0dk1JDbGHLf0P07NyRNDGrgrfqynxs320HsN4ke5bOLh
mAsQXYRnS5cEzlB+bjtisjSuz5F9PB/GRa80eMQFN0L3hY/9Dqk30Hn36lPSf7a1
81OiA6LjHDsNoFwmLlo3GmybruHIGYo49gzHA6KPUZjSawkJ+B03qaE5lzfVQr2U
f5KIRjzEelZbyFtGL0NtgDhRQRNwwfx06kFlmwBFyxHpeGF/IUC2/IroBupWnTNh
7BJohdO5qYsfZBAMS8aqxbzU5au3wYDBhqDjBPx8DfpqcJAM7gN6JbigZR2uAl52
NJrNyEUuFhtDt5tevjDpL9H9xLff994+W4mJ6/PRuDe2xKmWyRTm8I8N4yP4k9rX
OZ5eiZ2If3xbxQ2Qt9LIJZZjuXuAXPOvd0F/y+BZsdptrpzsfNzAFeBwmMSy1ejp
yZ0cR8+lWrWLhxD4FDcS811CCOb9bXTnQaJmvhh4IWOblieTn3lV9sW/g8EbOJaT
zJ0I+13Md16rwWWwg4d3MJaB2WiQ4QnboRxe5sbHcFq1id2Uq+rILM5VGC9ebPH/
rM1xfvO67S8bmPhLlrRTlmNRBtBO0L3NbE/MwnHouW42tIOiO4V9LNty/sZV3c/G
du5qKIhFEfd/hvDiLjw1gb+tecPkz/QufugpcQ1FT1IugIzOWqm2u5U02Qr7TZyU
rxwFJXwsI/TYXvB8J6f9K4t71/DSBgDWo7gvjR34ADXXd3SaclM43iDd5lVKKHmG
1Mqka7QnAepZaBKsPMwf7AmEXKGHM5AwvPij5LgHEj7HYFcw1sZDFd3rXylJyQ5M
PbGKW16hfAlB2GdGJYXZzvtFxq8aCv+EdQEU7C0VOAMhsAzqABTlKEAexghA+Iqs
0JvVzxXiiN9Ni7z6gaI0vbxdjEEhrktVDtPfKAM/pbrdVxMnrc6aB9oqBZjyC/Bq
8eSkh62vr9LcqJ/R9LCs9G/2fm3ApBpTM3m9b3l94R9S2Loh1H2MqJE9kiIi96Aq
xFDD7qXaEvMf9ra2IUYkbTpFKQOoOS6IOyL7NPGq5IHu7P1mdL0/81sqB+RgGx2B
E7DEucwwFk9tGWjT2QbkPsV10NcZiGrhahFGO3MF/NHvXHjs6pJ1IQLasQ8gHeiz
sXFrB9SXE0w0PC0ZKfpvmJwQO7RbiCXKnxdqjBn5YNIMUxByWTuu9zwpmI1FjDPs
F33mErRZQbg23WpI6DyoQ+uiq/Lj8OE8yZX4w9aFyx+iKe2V6XkUSXVT9bLpn1z1
hR5svTeZcQ1mMCZwt7PYA9RtAPtHpCrvnOoGlJ4S7RnBs7GGDPluEJS0biuPimfx
KdiB5P4c16ygUR9cD2QOKvjuhmS5oDC1fzG4vvYCcLh9ay3T9oA16RxsnDoMTQmg
zbeavBIjUwfdQl3qYbNeNKSZgkCOPzVz9c3TMurryLYa3BjsTzEZhXv3w6l+Beb5
KoEY3gphqLnXbs3mfW/HkheWaWy5OFwD/228nKCCQQqmArkLDBGoyhItdJE3dMVE
RPSCqUhkLvXcakaGxj8sd8DOS8QV+fr3TBxpKcUiCHhdQYDZiKEGM8oAEbt+uXDZ
aKN6FbtoWuRtUVsGnFdS1nkXXtZksqesKtcOyhc8+96wTCvF8Pd5Llg4/ZmP6UYQ
/WnCGaLvnA0DNE9RHFs94c/G+67bjhwx7mo9A3RSDpoh+D4u2JlBWZdUflXOnXYI
2DmxjJDXsJR7VMyv2LLF2MmFOrG+c5keuDrdwlDHhUgfAUg5CaY1UAYVf3r1bxby
GzztvDZuiaQ4UyJopfnvfvyao++d1DxW8AabAltn7LOCwfTsKjh/Iz6iykEzQBvk
ei21almdERHNSPMPVxwJr7wanyJB3YSTjtQHM1RREWvbwqB6R3t+3SiWL2qv+MG3
n3iMuqFXip1dBVSqz/ZmRoI6LY5gYSG75etWI/Hn2A11RYgOSqW2ToiNqD/0bWZ0
/RlJe31uX9tTboMvbQjTqnq8D85ZMssWhHqRr+c6mxkA1a3BBT89oBwDkvk1xLrY
E8jyq58NPogFuuYKM99Bp2J9L6ankzatL5fxsSh1hlux6kXa6+xCRTy92U4NDDvP
uxyxZB6dHyCrTPnYB/To84G7UpJRgqXHFQtmbByip9ClT7kwSTwKQ4MJuu9Ui3vb
qfB7O8MEKqDem++8t69VumhEptiHdF5zb6MjoZvOltHRml9jufTYT0gZrPfC1M/z
3i1EypQ5LB7krbiq8Wi0wkovUgjkxm5kvLGQWAloTpiX43l6QzgaWShMsnBtmiJ+
8GzQ4NhPN+6fhXeDzvWA6zz/x3K7ipyR560n8oEc7CadtvN1iNRaNLArEH0ydQZX
1Uo1iTBU28ryWgw+E8lCrHFG7AisCK8XZSu2PMwX1EHle808f03QwCbw4xQf3wXm
uSSxgdaa8JKprK1Vz1UHoMwc1RFSo7n+C0P8l/PIllmF/+OAv6bP35PLAzSe5RIW
rVkeAlNjrA55SZMbPUwaBR4QGUTnUehf1+vbUV123bRyh/Jf4gCStx/ZWC9CWfmt
Kyt3QplEBiydm8HtLXGFTNUZ86svB59d30JoNnjAX2GoqYy8E8qBd8MuKfVGhY0P
6Ltlc1HhsfNdPYtRI6CqmIHEu53VgpvF6Nk6Hx9ITCq71uygOLrzViYe/+QVW4RZ
7qP+n6iiZZQTU3wMQcGi42jYjFMyPEY1pAqvousSTtWUSuC/MUeE3LnG6scVdr5T
DDJZZGGJEQSddRV0odZuVEKFAZfnWDA/afh808NEJSCZebkfVWHpmavdKbYT/BDw
NaNPd3mNv8wiaBFQ6gb83+ck6QQvlTIeoWmKzIX9BnYp8nVHvYndyZ82EVZQlpQv
XWiAj4qyJxsgPJ9oGhGvXDWAF2KZZ4bVUu7phRK2ZLotlSafuRBT4oRSF3yokQF0
nXor19Y8Au1RBv3V52yQzJVwkdtVmO/c+x8PXavo8o0Q5dWauKYPTd3zpWE7gHov
Z5nfQKlweuDWaBSCNm6oHu4HzN2L5KGdFGL9nYGj64Z39hu7OJVlfh0mb42t04v3
YZwiEM9rzRbPu+dRZxealAmgiIqB5iWiAiH/+aUPhgLwHp5GhciRLPwe5n8bJReK
3+1+reGERFPrwLWtdBtoVWDAzFk1glpsWECG3DMpe9rf7vwKj8/MkQKu0d7AQLm9
rk33Oe/mXyItLdguT2fLoprCP+8402swJNXM+j03CfOXyg4o9Ii/3fFTs3JjAgOG
Lh25hT78sFiJO1dIrid3XepgIMYOfTbAZmvbwEcD6/SR1BbBKeiaOMUgiikz9oZ6
xAdSuQONYi9/5nHdff/65+A7VteUF3NBCrSXQH1yNt0Li4mgCZUC7qapw3JKJtyZ
plibUHpaz+fbCyRpy+p/DQZyxfV0KvTBYAYfzvxuc6EISTbqnotUhYxyA5vCQEgl
kwjDr3OQXMx3Vmo7WHERA8FiF2+euA94H50GUJp2aAHf5DDL+SFwC2xslh3ZzjdH
U5mKyBLlY2G621PdyZlPmlFTcsIuhwvRHfs0EQbimPvgdzseh2lN/P6vmAVOLynT
wLFvvxP3B49ilPPHlmv7AmHbsFLXMg7upFj8y2uOzsuQgG1zmKoatqFtJ13NTUpv
ejXpuBn/WMu6TEZGenzqGIxdvVncbw1AO5INyZwShIKA2fUlbZOqFh337S0msdGc
3k8UcF6j013ls4Ilj2BJ5YQCJUw90H8TM/oUoTksPlwcPPk8YnwfHwFxfrIv8JIn
5t+YCA1KsY2H7cDBZLBg6HPrewCBu2EiusW+OZLk504Q4NYZnuJ5TUtj3XJaxJQp
NgncOkZu9gwHXpJknMewMAcX+8q9WZAc7CeLqTPf7CvJPJOXvNbW1dqoUnhFNCqn
p7dJ2RCZJIPrJfbrfPaKXYWKIcWYJlF6gHpW0RZf/esf4yEm9Vmop+lyJbRLhJcA
aT89jdM7jievH320FrCr5uFysOs/6ytpHpHvnO3fLGSxpYLTGiHUgR76iCmmKN67
jamxICy91kH36Jy9lDmyx6Ruy8pul9IcOagWSfBC1SD6hxF6u/z2ZZGiE4TRCsnY
m8UrZJBWQKR4+fGVH4VBu0/KNXnwggtbZyoIEeXVCVdrG3jtzwctKORTQIE0Kva+
DjpyG11iMsJaaNWTqwqwGEZGEUr1DK7L2OH2sUeNKy/lbIZ8Pg0fSDFxh1+f/08c
oYZPoXbxDjpDUhToiWMfEGEg5kB8wIapkJytK193xt1lY8krym8JTNFm1FUBvNni
u/mQlYCZZYu4Ds9kEBMlc26sj9tX/Rk8n5yG0KojbIZ26KiaCREz1MlxnpyT38g6
9vBKl205dHb8D9Ue/bLbBAtiW9qbQL1/ypU+oqJscBm/AYoa9PeGDSZyNaJxlJPO
bLIRKP6bD/cFjdk2KsJn7RbwWPDaDZdxG+K9nH7xuy2vV+u5Yiql8wTqT3OB7qGx
PNySKVaJydtHR0jhQyN06cNgUQhavVqZ7AXf3O2jOH8kihePu4U+16oxjY3UmTpa
gUb4UD4+aUsNVJC8MzEeFCgrGR7PiIIRUAKfj9hzh93vO52crLrGi+WwlhAcY5K3
RiZjES4rtaMOxtZbul1BPdDMwqbhBQG50cEZFHhDnuiMHHiibniqLUS1RAmB3iUx
Qy+OVHcK1lmKZstTC1342Z0FEP6ogpEOiV5tobsWjQLBnV214dYZ2GbkZbe4Eppw
1ikCb80LJ9P3dMWYj2/ySOivwoDXCTdZw+v3fwXLY/fu+xz9ZYjvuqtVZjY16Grf
OjHYfNogUsQrjV5ku7Wk9+3PuFQBsRlVF8UaFpUwJakACZAMldRZYvDWocXvbRjJ
O8kk9p1n/XPe6KnV3uzUGH1OxpQrAnY4CpnFDKXiBKA/L3OCMInOejGVYK5jj1FS
oFkJD4IME72Kd+8q8y0FQoj3KnW2HUj0iefJhh0HyeegWVsVIHWMS5U2mwjXHl2p
monr6U+xADQlfMTnkilGn95xE25/4F9//7HVG8d6cn1fN8PIlNdHYmwVw7lWnHW8
Rpif5Zdoz5nOLd/RJpLo/3y1El6oYAKdhmzuxXmkyXKJHmQdKwJdtwmiMZkM8+Lu
1t6KViGYeUSonFOCceCC2/AZyfMScm5jy4PZ3e/SH6C0o11dA9/9YbyL1Exeo4vF
lmlSodE/2ImhTyNomTtS0kiTT2MBsAv/9OXzUUmXkY2upUJcwxQNHJXlMjCC681I
2bnJ6ZUl476aOsuSXvxvJOGnLXQEKwIhIBLBKbvPqDpoB6mly4rJiys7KZI1SYi+
3Hxmle2ncV9Mwv9uea9Vd01neWvTTc4cj7/h2WCDl6p30+VjhGejCFP5oR5LtF1Q
fJ0fVrRY32WOh7y1eNhPYSIdjsIZK4h7izm/xD/NLpjsmIs1w1WIie/24F3CEYDm
GIVVvmY9wJzVMZ2IZKV3+nACB8J5s+PVT01HcHtJ/ypCXAIwiIzCrl8j5J0J+L8A
c00pKAqB/d6d5me6gWhYgke/wn5tBKn3Kd6iBl6TX1oV/Pz7L58z0X6Pg41SC90C
dv0+zpJMi7MqCrMfmRIU7VMhkzXZe8BwStafYKnypTbBu0iUTSNusfht4PS0RdCQ
avL83eN2hc1Lm6yJZkYCZUk4TMz3OYhMd8KoiNH7cCx2zzlG+tzRFTSKf3folG3u
8Mk9JqlA1zFZZalpcBUz5XLIJmZRSuOgouoPyK38PXzJnJb0QX08yUdheCLsbHkI
ehi8dvr2x+wjqEaXv8wsIizJO/QinM65ZLeZuXNQobytDswz/kGNA+vwSThqfqpD
MQ7zUphacPzWMcWVKPI+C1QIy4gY8LXsERgnfbdkhjpAa6okABdIyfD9LlT1MZ0q
4aNDXnIn2RTRzsiXPNnCuAg4lFuaTeGqdJoYzEXYfIPxnrt2ENVD3fPnPc7Y9STJ
aA565R9yr5XWZhKt1Tlr9gZEzbBfEbvTIqm8TmtecJCel0lPTlpRZ8+Gh5xMvAEG
B0pkog8CRNiWTL1/2WEYVY+DNpiFKRPDMrdxo+ZplteODymGoNky2yTnD5+oWKt9
OLzVc8xHftV1BgGcNQC8BPu4s/xOU3DqqkzwO7yBe4jKntkBPfrkVd36IXw9UfAo
P8CplasQ1pqxfK8jcCg80q9oloJMwHfWFTFVH0bhBalbJc+EA+A6xJBEXL6/aJoi
RwpYxZ5CSZJ0TyhPyDjuRzbE1v1fGNxhGGhhRIT+rDt8GoDuTksLTyrTNX+6htR+
Ee+SBoHRX1X7szpS+J+60Po9cbQE0g9AHTepVWIfI8mkwJzon1CV5IAF9y7pxI+w
MhNZc0qjArjXZ+9LeGaOCZ1reKddB8PzPLfLh8tdR7N6j/Nnc1qy3Q4adG14sgPv
8Iv9pNEq/FTKfi+1Y+LF09AxutRpnasDDWQ/MDlgTZNlTL32Hdr3VTuUfurds05w
vLfUkhm80lKmak6EEzGTiIoYJuS/w9YGl5VE3ZfaybqkktAN3n+phONbZYV81xcL
H9l3s05zLPOa/wy8WAEVRx1eItGwwvCaJONgw0v3zYxEWz3rrceh0QawnYWaU9ck
7bHnAPNpAaoxrbnrbNmtZnCHP9jbWHnWJ4OC8whXvybg67QNGq3F+LczLsppbtIy
qpcibBevtlSRAPyaBXwOvVEDpbGH62fSbRSvCeaWSqIDj/dtoHpLU77NGcO+6ZB+
9MR+crk8euI02+ro4kduaZ5EOcSWyRQdLdyRtokkWzVv2dBDeYYNGPNBCt7SJbX+
lblfvN0dJpReO32vGidNCJlbs0hyJ7VrDIryV4c4ThQisg3n9Y4QT3hXt5BvUA8a
KLK1NMsY0kS4DuDpqIIiiPM3/GiHHVBc3rl9J+7BrA5T4vaT8R9hziIEDfNcmCmj
YoaTgtMk9fU+fUCRbpRiF2DFbOrV76JXZAtoeEADzKzXKa9kbT310rtihBQmMeyN
Zqkudnuft5hyI+oqevKv5M+B8mPxaCSYD1DyoLfVL/9Ge9zsGD6067eL8PBzxS7A
xDBPiUfyCj6ijo1bbClfpexnZM25ssR42JEyib2gUUzoec1obD418/ndjwb3RWU6
e+1XW+jNyTKYd34Q+U0S8myrbntdi1lvB3uHhU0wpTf3gWisW5gguJq/kUlf/IDe
91a09Are7HvOiBqFFNROHkZInIEgrjLQ6PsteJEOe9LmEdHOTul0gVNYytPL+M8J
j9MQ/QYtA+BTysp4RLmsQRzHRsGqMU+mBPpvTXy5Ug45p152fU8EWJ11SnPpwCSz
Vm/lVKMpTn5UtKkcx+r0H+1BHrJL58QeVP1XMoq4SePnlRSiONR1DVIWCksd5tnt
rY5WPAdG7cLamFVLyT7gx+PBnSzxmQvdtEvPfC29O8VTNK/G5PwpfvuOcxw/Q0f9
gQ4ggiWtrURQqSSrFP5ysi6+zEepdFem0Aeq6lFd4pXSvaJe2S3UvczSooY8r6m+
kbb7Ym2J89K1kb/Fmh+ka91Bj2XVDz6riQFCG6q5tCLMUTqD4YV5N9YdC8jd0ODL
/FXxjzykya0xruzsaOFRQkd4GLtApzgUB8hRnus/Q9M882zdKPXY8DU1mA5JZn87
MUCL6GN3sQo2UNzu2zzZzllaE6W21P5FhIYjlP3W4baX3CT4pWwL2gyb3NSabdHj
KrW6sA7AqFDM07otuv9JQf9YA0mmCrbsk+0XxiE+d5Rp11YrHfLADm13CCST8Xbq
/YV2uKY3xvoLmFM2Fwff6XlsMihOMpZFd+bjjjn8uLppF/UkXU1LKC83i62U5WWb
/pY5eVjM/Gus2hJIgITUr2e6PdVm43iTveoXIrSsodKPuhRZj35rsQcRuxS7gVIc
bkACviXLVZ/wzEZ2Yn4o5dK0DixrUbrNRvoUSuGKwoe/UXgWqsG2UXNXHWUeFBuS
coCe2drgkASfXA1N7wLb+JWnrigko23J/T6ZY0N2ed5Rf8hi92hcATgCkQO8n0I3
78mOx4DSQRNOjHuLcek3CEpVvkix4lIVhUSY8FiHiMn3qtto0AK62a2GZkEDC5L6
y8fnWAGuxnhwvZRzYuvZSEs9Zg4ipm6aweUTc17K0jLtcpKS30uN7IA3XlSDGkqO
Hgy9OLj83DdLzCvBqROLPS8wWUs4J7PYn/ws3jgp2iCiw4XvxNFHE7galqEvAMZN
53jedAbkyZmEtkbGmRzOYhUT6lLk48KqOa0gsxwFPsH7AAczxhjBIs4P1Kj6iIRN
5e5FtNIRMYZs4XiB+COe9Ic3p/RNl4tAjWuA/rMfu/OBARpeDOGiQz8pptho9pRm
HCzfsHpeESGOW23iWVndto8f5yH1q3prIVbPMhlA8bJnSazMJS2WAiPWeKVxPYAb
eOrDc7uYvntD6nxClla68E7al4cRJn6o2s+A9m0DwGEPebEkwqHCc6czV63eU8iB
vspDXyuTxZfUnR3+VTV9TpcP+o2sCM7ZMdVKsKePpypuT3VZgHcZYBXXRUCGrGbf
ciMphPOZCObZHLIdR8qRPRFLkVHhBZXPtvHn/MOUjVY2m/CRWdKe5aMEwqa11OVK
SXjrWcTMYrgB8QqM2dezt5tMSl1gsOnc8I54wKqx7RG+MD8DNtmn9VoU8mgu5Knw
awMXXFkQQfkiJ1/JXiexDpdaCsNKII2AF07K5WW5YUr65SsmkU48i8S5h0iOupIh
Qa+bAcUr9eWhueFoPPwk+ATXncGiAALqGUOjXE+w2DK25aNqev7l81ZvEvLGrh1a
iKLG+jZdUrtHYCR35tvaE8lHy9Q739SannURl1gDqH6lB1VY75bDkU2U34k+MvXq
UqracMf5T6vMQG1j+tuYaTjxRglObsHpclxOtaiO48hdD8/5gZDmE7VmH/ZLatS1
wN1En/Hy5QHZaoY/KZPa3u+mVHyzWSwNXzSUXhT/SfkZjk7JQ4S8lEaKiFi6JbJH
C3qUOmqTuD8H/v1upwoTUuUOA3GfnaO9n5oNtR/omnZHU7aOo25/hv3ZdKdjvMm1
+Rq60qhxGM6drXbc4s5rNNM8mcSuzt8kMxKWIfGTmBY8Qroiaom2DYhqgtZkoOkW
EWYqqx0EUB033etdOy/2vbif8JH9o7SIG0Ub9pMPeph15rM6zE7SrjtRikH9/FmA
G+/D4d2eo8pM2mPmpPU8yBXxm+fO1WxSthRS+MozTasANtEO37sRC7jh7t74sK2S
1SKToy3GONHSUT0YkkgKP4KnQA8i5KWyqUtSOypO0KileR3IcYao/2ZMyay+HNUp
oSXfRgKb7aZg/A5JfCwImq1Gu/E/j0LqxihZXkNsYL94pLigZnZmJl7DZ1eGBPoN
HyuQowpgAiNbwBVo5rjVM/nIXTlHLf5aOiriGTssYBN0xAK5neG3KO3rN+XA4wpc
gi5pBBQRGIk8QBgAxhKBCjxFkmlH5ciHq8y0g2DZLauComLd+rHcBvEe5dmCd1iX
FmdoHb1KM1ZgaNtGWi+WnMy4rY2VDJgiJXLnTma2Pmsee4rBRf6dyD//b0plgREg
3YByHiXhKGSne+LMFLmND4qpK+eO14dNhDicM3dLBdYbOP4yVG2RrgBK/JA2ukvR
U/H7s2yNpquBlG8BESALOHsi3SfXQTaX8BbMjXYOfYVNrdo3oaddYwCYW3Nw5xcq
82c5GHaTD9FD45uUTvK/y4ytzERdT2eMTPOlArJrbPdV4FTaq+lOSOnn2uTJamB4
XM1qTt4/aOLJ+rF/+xhIcMCk0j3oDdA6CAs2YbjoGOgNWiHieusrNJujl47jWmlx
gi3CDRWUmRF2k8xnc8MnVN6F0sU4WP6qClUs7s2k246be/47e/3kr2oG6ypPPyTT
VtrFNRn/c7LwkYdlOfjkKJLk/AaW1pFlVI4bttboln+zaJE0KKPj301XRseOdesA
Mb2dQAv3eRtkmuigbCNQpRkIlS692XuK3cd9VIAw8WZWfQOe+X5R6fkA+yOvoA0P
zbdF5wvqb4LIwensqDTCAuDx+5AzwgYC9vmMHjM35AuiblxTfgnsdb5sTCBIHA2i
PY1gJ1YS3MNW46X1CmLQQ2X3NY+ycxv1xctmeA5AdzXUuHfZ69TEXbPnaeRtk46a
qyadhtduhiWc+YN+R20z64dcPdOm3eBw60fQHvjyxToazi/l6FOHADcZWORTYXcN
jtbfiX/r1bt/Sz7U3aGsB6gHIbOyJ1YuFlxygHzSlOXoGiGjNzqQigFo7h/COE7q
58c8GpANZcaKdc0Hw/D+umtNQTAsvdyblVDYXTtimo4LhsjWwr6qZ9wP3JpSx8z4
VgWV4U6A4qkefziQVAcO9bM5iNkgGBkx5qkdLhZkSIQ6LcxMRPJMD2RHVWQFrvAX
HVEiVKsHKxuzTP6hKn5ueBE3oPN7VTRkxWwgt77+jBf5YKa78hpvnXCaDIkmxWii
YIvc79sswLK4gFQkUM/Uq8MMqyFv9Swxxf72pw+aetDoWR5xNTItzVQD0AspZ/Zp
N1SrD5dfr1bIyW8RZpCRVp6cxldGiv8r/UQEWc5PYgJikeINaKncoBo9VAiLmIEC
UipLShzOFzml7JQPnwd7YEKivStVGfuLaqdxEyqhWe0ffqTg8UwlAOc0NS6fCPMn
J7w1sFXtPQish5g//jwjhiliB3iFhpNAlgxG9b13BmJ6nW/4j5ALn7A1NFxy1cUJ
5J5DlFyIzQxugf28IHWOCVkI+qBp2w3A53tcWni00LmXxvOyhN9GyqTWsL6gGb3B
ZjZh+IepE19OSHoFTSLeY+4ZMt0Xa5MIW2+AxefQvCI5S8tQI7yUQ2q1j2VJOseZ
pTecs/lEWGXBhS/trqzfBE6aUhblzDzeKYMrUTWErAtWdo0M0K/wGMGjYNlfpZmC
cuMcAZAEue/jn8CiWUbCu+akVo6BL1B7veMSQaRG9rZ+Gjrzc5YHNLwXvy8QnopQ
0+GveZaWq3+RALoA+sjKqnHCXbRDHPFev3Md3T/oiitrl+jnWOWqV4Vwtq2/WsIx
euiYzCaY9eNQ4zGE9HTo0Pu9855v9F3oBKiKmVreDCfJg2YnEdKSXK6ipm4huY59
TJHRJHiPerFdAGTuJFTkgo64tAtIVzH1i8KIFgQ7lpGW3d+8MUrbRCUcAo0ohOPL
R1g1MRsvNvDBarK1jkaIYFh4DphoDT9q6VrIbEwi/uJL/kFSVFDTWfOXYox9nzYx
IMnJ2fck8+pi1FBxM25GPmnZl95Zw8dhtOs1R4ykz04iYKG6yX/P5M5WHr5Dt2Q5
wNrGmF7N1A3xOk5YC9psrSYEl1RO//F7R8shxOz4V717x4VghzkBjTn7EIV71eXt
hbNEn5mg8nV5EvRwUVcgVVzysGZsx643ZWTnHq/78QzxoYc4NKHKhmxAxv4NR2TP
IXujcrmPhiuTudE0py1qbI0TP+meKz2SyRosN5coqtmdOXcdh6COEUPyvTMDCylK
gQG5iwnBjta2Mz+FAYI9Qr/+hYMw7CTYndmkN/fBu+r9PfSlD5/l5nnB5KEefXUp
M7KXQC0LXKjDizTCCg4VLdlUfAhOkRloZFnlXMi+aO84DDH/PUJVMs43wCMktsfp
wfLdK1aqGvXmXnc/PS6BPq/3J2vdRJ1/wJGD7lVWg8kLFG4K+lSFToGhCmm/BwWt
uI4nOMBZ9kBS7dHNPIjkL80rUo8B717ZXVzz7EhwjDYsaAQytSnm5dIMibIzQ2GS
Llrpl7x6N/K9Ei/lGmZZalUczf2Sd0xCqZ959MKGgyCSxmdF8VerJjhSnkNfQPLr
MsTiU9OwxuhZd46tejJrOedgmWJ8pjV2PMAn1PvOK4g+eAUDyWSz5oGOtabpCyEE
19Xy7XUOFjREdYm5wf4UmRTkChe6n/RbLtuAAlM/i2L4zw5Pz/2uagvKt9qyqPqn
KCmWIW277SMIQX4pZ6t8w8aKnHYgE7+r5RtINXE7ldpuN/oUYYbiNuvAgKcQBsvX
Dh70pkaSIlzx9kcOIr2X6MOGx4ibg0y1T55zBpxQfyknrbwh+5VMDdkbXrdel2cq
yZhvfD812frbp3wIRxYAGlaJM6AzEmGUNJflYIZCxSCXRLoDQNGxtz2gXxY6Wszt
jNq3/O89rptU8CISMWSQxOVgtYxsTbZbAA+VxyJSSulbCr6Vd6edYBF56+re3OKX
2pd5Mj5ZXoVj8xqVlqFnulFFn5MjAiJBwdokucHnOlo91eTdJCo0BIjGgEINpcXl
cIbg9Guh1ZtMXIt36RMoMY9YCHyC6HoqFGlWYjGTp6WFIZdyTyRYtV/Yr0DoYHfO
O5kJNZo4i5JLgSjE9Oaao2cTXrlAZEaGjA2fZTbLCDHFwXyfHbEJsBfabFf//bDm
OcmV5qlpfyficM5HYcah1/co5kjh9HX1V3S2RA/Qu4l1F8TPc3CXhbRZIMqtatwN
UNUAha/pJkgozYhiGrZb20v12XFCuGykBWJCnrQnGNDijoTRJ2Gx7kgetw+S+I47
5EQupIZTtwED5bxCiKOLzQVwXatZTgrGlvWsosEewtU9Ea9cbt/f7+MRDFKsvdkb
YgTgCf0/YRYZtvv85/T356FoVlDk0pVz1Xz8dwr+3sY7CBf0yfWqLMlZzjobDyMh
OjPmnLa7e6Q4zyPJqeIBzUkzt5SrBfvSDFtgjYQzenEKPlCjiiJrQcsooPLpkXBy
oHfEwWH7qx/xVDGo+kUj7fMIPZmXmScpbyada362ooDHjbu9Smuy8F3DgJzF5run
XWsa58Ly59LXqOyVlwVnoLYonvVVu+1FS6v5at3CyrwCmQoLJkqLN4vFRWtxp0gS
7mYFRMOw1gPa3U2xDoJIzm2x7P1KulmAW2RKvW6VwvEfALVA8tvJN33xcyX+CtnA
/C4rBlilGtC2Boq/2jcHJa4eK6QuExCHedg1D4A2p3kY7iSqneW9I1yS4xirvYWY
cPC9N4U8FtxVz88oz+zcafj6efxgitAZ72Lf3Cm4ASoQI72RgMc13EK3AbnkpXhd
BiA/QEnepu1npXz2eOtRVprS66FLMUiKM+mW3zUzxRW7xLBi0c0QpFdBTqStT2+5
DMW7hGqGWwTpwlQOmWB4TX2Fa3F8USm1eDWZJtEWhOu8foYeMaBwu9TbWVN7f1uD
CgDOZREZKUtvcr1tMC07bFJ213mjhFMCcjkfupxx+1P0xo7C8KLh7GAu/xNcvpME
eHOzACGiG/S5G10qTLwEcqXs4eFBFEnz5nGDbxA58+17w2v9pUF6Tmd9R4v7wm0D
XmyVncqYylQ136fYDRbjogs0TbNPOdWT88m1wJ57dqUYomT2m1c4weTn7YCGslHc
8mcf5jOf2O/k9Y9756RX/qh4mmgFzkje998SLy1naE7pxiC/N4GeB14/tQMwPe+x
EG9js2eR9CyFkB+6V3n7stt552hPnJWhF6+Ryh4X/5TYZVHiTWJn0Kk8Fiqm9ZW1
Pz5DBhsYo8vHv5+ioJSHOolRL8Z0pQgdttI3ik0WAA2Bk/e84kDA30zsme+GJfAn
5yrkbbEYo8YaC85lCJD8QyZVG126pWUnMg16XbGpvGbqzaXq2OXfD/TipAIrLNic
7D5TLXKKfLlstYLHuGH1uInLEUZ2Ir41zZv6nbDASZJP0KaTlT/YMttTYGs4m1oj
X2h3FVlaSLfLeAo6pVkMWMBaC6r8NZqHH3dGWuYJx58pxYJZJ2Pzwb8USTy8jv0V
dKUn8P8WbpctZvoTc/AkNQlxOkoym8wacL2olMHE4oK8h0NCdDmB9k3tRWlK70rP
qVqn/4O1K9GuieeUOZOyh2uQMwBePUvGxRwM2UUkYDoN25mwT8t6yUIE9pCYfaWt
WoqDlIv11+2dvFUiGTbOPYrMdFCE1yWIWq7olHmfJKioenaOL9YJMQ7p0KMxLJ2G
HkwC+Yrso4MMgBPhC0LCMvl9zUGdlZRvMd1WDZEfx3wnmjfNfTRhSAC7A9xlMM+W
HjEKtz0ZACuSWBqBFkCn0ELhDeyKudmnFAk/z5SZRkywbU+1GNDGYyVKGiKYfrqC
T85Uj6eoDKemN7FP/Aw375C0e/SyGZeOVgSthFesZ26fcPMAlzHT6Pf//vBdbVDj
9ildRxL7AVbz8Pv7kKf7xIaFNM4uSC+EVZ4tDneD99BnrkDr4VZb9mrMQEXdtjG/
yDheynR7qbKkd5Vy1GM7859Tu6cH8+N/vSSMR3d58ejrMgq+8OshSNK77m+V6zXU
DR2P2TghoVsZH5XfOlyEPUeH5Vs6fioYeIrh7yfIhvL7V2vM8V6OR+9++SJ25WF1
XJml88EsmkWVS1IVdvx0jasIR9zrmyjP7ZIFaWJuhEleBfu3yKnzcmiU+4gYLlTb
wxOJ/clguzeQ04RHG3CraSUEnRGqutY4rQarzmvsr4nQhWGTEXjogIw+TG1DjEMT
Sz3NJgGdir2RQO8RJSBFYkfeZH/+h3MUv6nzQ9shj49eqs2pqOJQuDDc7oekNr5A
kxFDpRBAQOfI6ZcBNEO0UosLDq1cQmcMn/6SrVPT4BgrRXiMgNcgE4c4cPub6tUg
xv+qGcI7TiymZrt1FjqATFA7J9xGLOoynzC72yKEPkRpMteS8KNKiznNSNyxhkep
6HGuCF2/sO9ZS8lv18XmmrnJZy1IyZipw7vV1d6+weTQL+C7xBV4wltSUke2qJDb
Nw6l5SMYzE8MyegCKxAoxiv7GOcQTunjFGWP4QreCEHjVvvidnA54AqFTXN6PD32
G2bC7LA6tPz5GoEbVDeaD4FcZ8wTape7hMyiJqDcuh4zfoRjMsTBBcV6WEd6vtfy
dsRSqX0dEr7TQQ6DcdaxKdkj6WJLq8ZKdakTNhC34XkF8G0lqWXTm0DEgrNL16sS
d8N5oeDUQGu74/DeE7l+ZNoYohZ42Uh/SL+YIIDIDpPVRqhgnN/AKqKzrEct5z8o
t43yAaBL0/R7SUM6mnSeD1sK1wTf0yyC2+M7g30sd69e1ySFypIfCfPwzr1O96Zh
Czks6bEKCW1TZUKRjVqsp3EnxfW5sp70JNKj1IQr+Noql2CKOeuGr/oww0hACmha
tQD7ltIt+qy/i8c6m0LwFSwXKvHwNkk01W3kNkUVVKKE2xUtHA15pqPfzL7PVG30
krzrrcpXDhJ2LOdDLn4rY5nQxRhliuzYDDZ831xxDrj7RH0ocRrw9dksRyuIENif
VaCX8SQ2HrSv9+KCJRxsDw41l472zgNhEM8eKlNeHv7nJ75eHzhydnl/LDS62Dpt
dJCgEVAD+VNWItFxJBK2grR3pSGW22NU1zyozFVQZInRMIgixDRTkPbUo9aDGYbx
fBKAn9nugAs0kadItqHgpyRdqnzTZBkXnDdPWfYNxsO0KpOoHTqZusabQQMBajzd
OH+/JMtsDsVxRF/YkUKf0J5ZsNe+pwr3Y6TcOFT8ZDctJ6hokjBi9CIu8vMGvrTm
gglvRoc922Gewa1+WtUdMFj8YiKtG0sqnTBCJ7D5G6YBQAwxtR4KG6iF7AoSbweJ
fvkxp5C5C4h6kENvMuQvZvEcY/ZDO+w8oe5WaaeJ/CylOmccqv3/T9ceJqAbI8OU
4cw6aHYhviCoV230f9itSD+mh3WUePh/SJjPUy+aHQ3j0o+DQyERnWDBXX0FWQEk
XeUVlBhrum48Nf0Tai3oRqpLws2k1GT6M7rQDzxhoNWB9n5hWb2y70afZBoYhQZJ
eoHBs9YCzt0tTbhP7ZYJudv2pdzpIKfUBJs44Anm3vLC40Px11uZ6GlL4LUpRmMI
LTwR/zdsIx4CU7b5Ka99iwLdeEUdfGXFDIZ6J2A6Nzvmtmgg7ebIeV8EHPvJ6Ums
UZGtNQHKRPgwMhUOLzuIJw/UgrbyDREbi2jF9OF0Y9c7xw1K35A9YxFrNXd04mYI
cFM5xTAV7e0stBd7S0LWv5LcDsQTOT92D5ULpHoT8IQCLC+gzQzpSyRmXfX5ZCfO
u7ekttTFGYfsGZ+Q+kAD6zzdmDJJ8125CVjrN0jgWfdU3ka/rVYr2E+E3UFmOXI9
cBPVkhwilkbaTG+d7HDHrLizyXvmKk5W8/lyIgctywDerNbJjhnQnAnkEC54cmE7
HlQk1ReDRnU97426oaLPq6ezlLddTNKzPSNjHE3Mk8593Wwl/tZ/b00ewTIkz7ma
wx32U4EI7YIFSz8gZcuTCEZyEOnntzrfqctYN5vVRzCozxjEFA3jt9NJZGEfNBiz
hhWC8S0EEy1c2ed2odb6mMDuJoNQJ2tD4z73ds7Q7bJdLdbNAJsDtzieGhrM/8SG
eVsXtUjjzwCV2spa9G7W+BVrE1dNhg1ZrIqepW9ErJC++D7fJAzi8gDsal6Zb4Z+
vIioG5ar4lKsyyMZt9wdXsh9S0Zlk1eU23yhCFdvo/fbfz8HI9cXeaoHed9cHmRl
1O/Ak5AjkvuUE908/deLYNvhxwZn5kquX+Qn9/v7mRzEMuC8tKXzzv84ZSL4jAMl
ma6bYWC84TCSu7mxfg7NWt3u1sOOkIKXlstrqHvZgSUz5QUhI9yLPOXQCuOXrOq8
tP4wRq7gEBZVUXC3UclHuLo0mv6XKErOsy1HVlSDblUXOuDNVSHx43AsoYeX5Vyk
S6OVMFr2kmyUHscwGnkI+o2+390CJ7UfrSziFKw0zPypUT/nfI0bjddqzhxcOQ7o
1aeujgnfyfPdA/QHQavMro3cB3U+MG0GAVX3rbHGBhSldJQ7lh49nduef8pw08FT
SN54qp7ND9KzLIvi+vGQ309wgmIFPYbhnpzf/FkN06ejWwo3qmY9IV+PJqfuvhde
Qa+O5/UWaU5mvmI/+1ey2rMiDUO0ptafoilj6K5Dja3du2FKyqm/YCPSySXiGKyI
OePDqf3YYQ6g767zuY/NZlNnXWLuxHpWwKZQ66bejxN+9tQIBumJL1/jlbBV4Suc
NT0vO7UZ6w2aKtR3MmHMqgU7/uxqepjegmiT8ne5RPIZGSTkm9KydYg244aYkijz
nhS7llKQnfB/t3bASjFURhZ8RRcmBiQkXuj+HSZH3lsEhnhsYiZ+epjhvKRzOg1f
hYQX6kwVLCpqFTyPxI7u9Sq7OkwdFf/FnkVxmmMprozOFWv6phgS+pdHhKcz3sMq
l3lBm9qWnrVOtVzeIAphW6boOSejlIy2wRrpDKHrx+hteN1zkMzcvtc6XOYZLKDA
bPwn8lVCO9/bEpcgnvuaw8vwq0fWqJ9utEY2xCXK1w2PIKUCL00ydION14ftsyrI
FHbPuszMRwz9ThXKLHMYRkyRFkBCK2O/2cQVEnV8jf6j9XAegpXLtLzaI07pGpVB
fvE7cn2fT5/raDzBeRjPV4yhUmR2+2RujNwHPVJmVlYQHu1EKhgp0HoWN3xMTdQK
mccgiycMn8GwtO1q9Q+kQZMv9UQ8yberGptT+fs1iKFcF2jsoSNj4RgROo9e31dS
OvlxCnBWNkA0e0hTsyclpp2tDsLDJHSph/GwuJ4YSEq8S+qKyddXf8hVTytSHQEL
GBxMYYHcss/mjKB1EF4jbmFgpSlS/ygeQ3ykzd3z8YiKZViw/C1uCtX4IgPe1pg4
yPXH57PryZ37QAMyI9baGKnyDdSE6QxHqtQCCpmYFretRJTqv5SJmGbAXzo8759Y
BGvPIHKLqW+myIgpNDQz5hm1T1CUuz0XtvaqtLtHGIkAQUYKAUrnrop5NxwPW2eL
dksyi/AE3T1Qz3ZD6hYXGpc88kSsz43dImF6pcVeGFjKpisAxyA/WMzChLOf4S8Q
9kzykNL5lr87oEfOdvEgjuieOU/oJJn2MMc7KrUv5DqMSXUIp20zmsBl9t9u254q
xKULnQYIN66Z9q2AZnY7lqNy93WbPoqTwWmom39jcAW84XQzoCRhrPWZMZEBJ+6o
DVGkiOju5eXN9aIj6qzL3bVXHSaLnN/X1Gx+q7PIeGRax8sRQQHlD9AvekJ30zAH
GDenkDW6q0kgScW93jlAGvPufDhxUAW2SbdnyEwFjD4wume5V2RieFQG4DgoD0h5
emrFkG2rfjn0mGpNjZGAkYoJqwGYyBA0bDMZOBWKN8tbMvppEY34Hfx5We4imIBP
ssJQsOVJY30HGbYOO/Ykk7J4VYs8mQo/ikumM1+hPWBni3ULHrhnssZfSqTkbq9u
rExUVwkxIQgeKSsvvX8NaOSsV6tUhyTaGEEw+TQ9QBK2dUO9pPcs7zT6cVWEqSsP
C7rWC7Yc+3JVobJXjpPETkKmQrWUdqtKCg2MgBkEDZH0LRGGsFXlSqZsOqOMdO9T
TJpgm2rPa9pSSVDjDc7kxkex+kK21NuDu/ndVEv9aENWbBPhaAbNVsAUk1aci0up
WkFH0cMagxDIzaO0EGoNMIEeAYYMj1525ws+z4KHbmWjw4RtQ8uAwpV+DFNXko7V
ESElHzIRpGS+4YOT7Ot48KjrXbxusA3xKoHZwj+5CBTvW4hUr2Hr76DjVFf1YgNE
9nn8ZClTVAB/OKsgLIwyYAETvVb0EbF/qqP2j4+Mvu6NvxaodyFt8tubNliQ1dho
FCA3p6cYUoSfhqDUSqwpU/YnWVlGOYwsSsLONyVgQrGK+oQz0NkVSVQWYUgbYNjJ
Rm3CJ1hJNLFoeXOUOVvd04D1DHRVtX3GUFh48dSisGYpWUXIzUa2HuSW/ohSX3ms
HsbWqVatKsScSwdKtNHCKScQ40XPG/svvwYgseJu2P1MIVm3u2n6bKVPTSwHT30z
Z7At7qC0jMoH/kwXVy6EuB7snsb3bqGOfHkdWGh9ZufBixDgykpwZ0WQiooiixhj
vLcu778+Ckna++GJBgqVgfyrcV72fr1tbsC/J3M4YZcNytfhZvOjXWcL+H4/nNaN
NEDipVfoQk3UrlxAQkQ0d1D/YRStsb4Qf6spLx9sdXAwirOr5AkOvp5XUzIEwa+c
VzyIBFsJbypKSYTyJacX2gpqrG55NWla2Vtp/twW4abRem1hZbe9e+Pfph2isrO5
sXRCkqSNiwFN7WAtYC8YYVIlPPI/r88YVa6xyn/Z5ow/Mrw0iAE/TGFSjFI13uvA
+QPdlkbCNt2ZAptjRbybqNStcrV7TD8NkHYodWCao4rY59MTdAGla9Cdppe57df9
Aoyc1mk3cHjHi8FPPfor0d9NvhA4oosvf6GvzdSVxruZ2SvnQPeyrNxEZMytLPCI
1s2sdIcOzzB14SLeqNIK62j3jsKFxByFTB9bWhdU73v54H2Zpn6vv4nZ+t/u9JH7
3V78iH25dc0nwldlkrpCUAF2aObO/LfXkCii7He2XClNb6IIuDj4tIji3nWaPEP6
LR/hmF1/ry/mjRGSpN7Gdh40R75/LavjQPRkSXDUik1vxSnLDpgvco/3ssHJvRI+
KRgFsN85cq1ADTp7FBxOT0r96wyRsODfqbOYPxgijCVRJnWYnMWDSQhfvTcudgzh
zCStmwC8UoaSNjWxKlXOQZVPbMyIJ1626tAbUBN09RQZ+4j1zPj17xKbUMV9No8a
HxWEkd84Cq5drFRx5Nma/GDNJ7CeMIjVO2W6I6SGZyoZR95v17LYQhfvm8FD3d/w
azzNxNPkz86LcS7u7gN/t3zaoU0naBgawUev/wOF2pC8XxQf4RgQ0tzghStLEDUP
evSvJ7RE5QTfvnfYmtKRH39rRf9UfmAjfvR76gyUVfWAjn9q8rGM3NKCRjG47sCI
+LJL3euubhoE65hB6R9EbqikH2qwiA8hoRBDlo5IBCiPaAdGL/4zPGLQkPbcCVB8
FpUKtl9kMlR1asWMfi1HTg3E1R4DxkX/BcO3nNZ1734+mgkIzkk9zGRGU0TB7Lmm
PVLEuCVqboz+3sFHlvrimy0FxZRPdtxe897L5VjsqBMcmpk+a4AHwxg+uoiSBgwn
cM70IraE+igicPj4MOqFRuYC9BTbF7tBIF2Ue+aATXpXm2B5uHiLj+pNYafxmLQH
DpZwtj+aRUZvCUwKZ/qy8UnYyRqDIAGEx4J3Tta/oaQPl56TTZ7qGZwWIXbf8qLS
dp4bGMY4tTiIuJnu7iJksM7Fe12ydEPuhSGSrGSh/GOveLY256ftGclq3yO8NXWa
GWQ68pyvKcjI8bSLzUDn+lon9shuEgA+drDxbZElP5NqaNzgo5vPPkSe6Zxums9L
YaDt3hYdPER7QJMqCwnWBxaAw+ESSXLd78QF5MgS8QueQ41ah+ij+ZpD/8clbW5c
dUoPwdmmgtn91RnbAKuDoiX7nkDa//meuosgaQshEZOv3LOpRNzNoLKEqTozauF9
DtAb4I5AWfo+F/Bf2XiO5WfsLNSVdyizeuGZ2V2ivjLTcJlo2X/Ga8mNA0S5p4Vc
je0XOwCzMSRuzamgumxjlsoGBeRWmyCjAI0T53OwOf090HAtaB0Zrz1WRmld/3ej
lsjVDT0Noh6gY9rwhTpi1gUPXw067FL76QKFzpY3efLd1annllUHJO4CNxSMhUFt
5B+n/5baA7ds0ndfg6Q8X8AtTBrTapjVZys3z0WlyE2HOQ17/qoaorsvx0aUn/T7
RYciLWdGlTCst0+gnh6+FfKAY1eqAjTTVZHQCdNQVTwF1ytfLRgHo+sfVKd9D5hm
m1yvhzKdk+HppeU4MX2NpAo35GdXaUHgoVoQ3feGvVw/KnVw4Ak7EO1lNDCrUy9f
8pp1PqH4m9n+Z0Q0l4qy1AxBqVn73QeRugUUCGDFO4pPH+dgySL3MgaOkCrZHLu/
skkHR4juUki7JaZJZycwnS0qfR3Hr41z6HLaqzH+Sxmy15TTzHfutR9K6Qliv4c4
6S3S2POCvvDIguP0lw2X3u+vEWoEQvYgn3MyJL23mGHNxjOsArnsvgaf95g399iH
5qz42p51UC1e8WVyLElPh7LpqyqvmdCBXFoiDuGQ+NsjmHdylJ/GBhTvnoyVbwfb
bXbTshp/Y8nxmy6cCjrEjbet8BOa1VdQ4iir9TlNFIzMEsvLNT6PD1EtmVB4BYO/
Dj/t74uO3LT4A2AMl7/FPQw2tYtYchwqrSPgbZ0yv9+9sFM3jem/4IyVstyk3y5A
H1xdJKQMI+ZLr/BdDE4jYJnlr3TIJX9XpNij6igNRIJ0yL+CBTP1d9vuqUpOX2/q
LFqXxaZ6f1ilYuCXz8rudBy8BMQncqbWjQ5zFWiGRJ/mHJ05MpcQlrd4EEpd4EOw
A5BL4A+ZKWN6423AqfTtIYdibMxMBL3nk0Q3hB3E76pY6Z/DaZo8GR+ufnHILM7g
i2RB2d0LVCy+d5OJmaJCQQyCJb9wQyEi4bxVvqQd59ot8m3YZCYid1fcxdYmId7o
3CNfL/vb2dRCVuyqH3oFT6ikOZ1LxEJOgjBcGO86AXLtB1cTcQk6oO028FJIEUO5
+kmA40A+qGD1iqqBnxIigSdSbMdCzeI35Jwsx3mWB1Ba5jivHIapZYmXsiH9vv4E
Mxjc8lw13tAcKvR9i8ZR02U7G8UDdedZQLwzBi5hfRo7qKhcv4J8OYdKaZQsiD2Z
Gr/mQLLmcEUI11RILsmc9Pjm5TTyB/FDdq4ZAab+r1lq5RrkYqhzZ/j00u5vXSkU
/Nko0njpVAbJnyRdsaScITD5LKbf7BEZd0JpZBDC4wQxCupky4Elx03Jz/p96rGb
5YQJYseIZTW/JnDp/Kj10EyA3/5i46gPmOSfvGiBhpM8KYysjedRBw/cQKMwHgmN
s0saoy/jQ2EVQj/VCpguJb9jZ880rhO788V0Sc1kuSjjNMiYV6A8yk1K1/lSM5M9
hjcyTGS6Hc4KIi49p9q0r6JUeq/OZ/ApGHnKP/lWLUpNsu6VsKey2fmFKw0lalrh
eTQHv54BUqIxfwc2bXnsG8onzUmmvShI5WQBe2+8leJNhbkNhwYUXO+7bXautEfr
wNvOo+hEG7QMwy5Dtg58JAAyt46cchd916i6d590tdoSzlDOejbEU7aqquaPO6WB
Rt41R+kMHy1cjlUvp2gu0ugck9TZwhR3DfKpJpQMqMxYF4ub+XDGlkGvbBTVj5tc
qj2mQxFkRFlh+Pg9sl5Q7eHAvuLFVCJfRcbElby6jWWHP6WR6iTZQ6bKOH4UMIgp
Je9UvZyicB4loHpkYfRYVw7W/v1Ev0kLQhm0s+9uJwz2UjfF37shZKduWLirKuBl
ULMTR+CtiwYgFfGRnH4UzFP1CeNrVr+rbcZhm+Ns97Ndx9zgsiMEBuca+gF80sow
a/ueoJPAElnQA/1dlVieSNME43bz8tRFK6PlawlQaTkpu1ViHzWbEWeZrqd4ifI8
9NbqY34gFG1J5xhyjCUEwZLAKwlvo4NEddKqrckFJdMLCc46anGDyI7xCArLWqRo
WXcpqr6LD3k0haGliePFVpz532o10PL947TGb/DrnfpioaHk2AiucUK+TTWtuX8V
A5MJWHaJsw2YTVX9FscgRA6RIP2JaitFKQwhQCb/D3s0ofzDuXsqT1GjE3ig280G
Xdo/mmodMBrn/zX7IIq6adg9r/qypobLQUlxq/v3ImHW2tl6Lfe88iRVQer4I5SK
QFtgalhDI18tisO92uumeLKzUHWxdVJAKooUEJZdE3/KrcvlZR86RyU5xBZfZW1N
qHTkY5jiMRl+z/8GOAoY/V8HxZDey4sAJiDd6R0cxVggjDVze7YZ+rh4OiYwer/P
eL07i7RDy8SToAufne/tSU21cWWnWVBvDGUIW4zkNXFvEi5Znd2e0KovDG/oCq3H
XxKfQFiAPDYMX6tPqL1UwjgUlLeRwpQVRpa/O8VEEVKvq4HWIlYUrxKR9lEadGbz
AjrlittETIvQacn7Tg/m+mcXEdjvne3iABNqNXpjWizBR8ysS9yR8i38OOdeEqz+
itbbj1SAouCdLY4Ws35q2orsfWU80a1/oZQ2mf66r2O6bI5sbScAkaNil2s3wSgq
HcJHbvxTvKNBJB67BPNrCRxv/RnD/69VZ6cQj6GwBJB81yv8ROz3/S69UQlI3X19
iTaaflsOrarMbj/tmQYN8vLfik+3fBxZU9sax1ecopp+o8eLQIKBcDsYV8cYA+xN
kcmfHACvphznsLZtkMt/G5XjQPYOaQkAWF3MXBJ3wVGxE5Xl+b70LRFGS2Ixh7ZP
rY7ewpaYU/HU95wEWB7hRSAK4PQb4HCjT8Mxb/RBpiPFuErq7nnDd45kdzfgK2dD
YET5n1Vko+fdGnYHmHaddtObwIdrCFQNT8TV4bC91SBgW0yWErkIbyF8G11IPBua
xFo0/PpQy+aBsdLBbqIUPlRrQKPkIk4bqqA10KdNkGb+CF/DBPyYb7AuebhT143Q
Ipi1EQWAaZkqOYxzm9D57581oG7jtGOfqnor77PECvC82wtTRTXfVg4X8p+4lde8
fBUBm3nU1iKGkWqkqmHSLqnKA+2lO2wxeobjlLUk+gqmaEP2Oq3NKRhNxzLibiC/
8kUslZfJ/l2Dl6pS6xHzssqm107YAZOXtnQOsArHrIjqG5T9pVjiZqATwNOTEbQI
vTJaTNlyKsB5S/oOHONuc/KKUuEE0w6M+A0fnTuNCyQ0b10xVY/gRNLvgDfRKeaX
49KLkczfPoNBqgtZNyJ9yGM9KdUczznZDJYXHxu52XOoT7qgSepM7BzhPbxJEOan
5guT6pVhdfQ2e0b+R78/uz7Tu1cyfAm59CKHY2Iwh7xe9MxhXfViu6VBIeZeGmtq
x/+JO2PvnSwxK5wla8J72zFeWe0v+mbX/riX3lgw9Pr8S7v4Vwp7PKqp2tijnz8b
HijUlX8NKOeWHSSP7bC3JwoGFraGpHVkf56wKGIrnO6jmCGHAnp3pIksdmlVs79k
kSEEusci5OKFz0nKcVa25hbwZHU51kq9446n6+lf/EC2SQYoxLotD1nK2AXDnCqt
J6lkY9ifjQmBGerql10UV7WUI9+mHPkeSrZu27e6mag2VOScmbVYl23SGOUMe5QV
kmQ/hT5s/ET/rJ4Y4OCrDIfEovby7bIsTxHCogAvUbi1XV+sTkpPQoRBqr1O2nEK
tEAzdHaImC0X/2+tmUG70qk9kPQXzDDxTYJ5OiiDHFrBCvBGHIE2twKk0Wzu8PEY
AsGcSS3JUgHRAlB4QyRjIKiEoXCtaIul8iY1vxQVwz3lMKqLTa2C2SvDfWwYGuBW
aDpaXlb0ioDXCEfoFggJ9nOh0L74SiAX/PWwTObXo1Rde2Z1Ff2m/AjIoGFsmg+I
uAuqebybF48504rl6+qY6Ub8x2FvKr7Nk0PW1aRgMQmffDSm71VKTs/vArZFm1hb
38PK7uRYKpmO4cEL36VPkLMzWB0i/eibObTdz/mKK9S9+Z9YzL8S9QkeKU3ax7BC
9qyCU/rS1Z1bFtU0B9PzQ1MBmZRmD0lhE/eDXtG8qkeqqfOUpkRkV3fczjJ7QyEQ
9zFhjjTJ6Ux5KUGDTmY7gJfWRhCIMOzrgJq2GMJYTdcFFIH9OQM4LQ0w5t5KrX/H
mpAFc7J5e58u8vSv6kQC39FREyumXxys+oOGSe4tG9pOPwMQrtV3kATUA3PtTwUP
KXwDzfukOBW7EAOX+EeUrQDHnJJVpfGG1/3pnE2e+MFG74xbRByzZWiRKMTMLayE
P0iHqRGdcIxASNt8rCu1Gh/zvwO2d9Dm3Hi9SATCV4daTUZfmIeyEG271eDztplN
VuOGpA/KO2HsUQefP0Nz9qmSl+x4zRZE+S3xjcaYHlsLkgumi+VistzXWHEXnytF
Hv1P1K5uC1ZRbbHpCG84MPhS0HIp3w3NBwW6RVoT1p9B7zM+SbuBbROha7TDwwAi
cAQwx83ws4XBvHjyU32vfBBRrOM3vmMSpcJGlwXaRsNt2+v7Q8Z0pke2amB5SAHX
I+sArhjstYocD0X+P2yQVrdLXUYgRcoOAuw+hExF0ruP7lH10TEURhJRV6mINP7q
P8j9ZSbgd2Gph0T0hDvRrrveOx8RSDyNqWbKp8z20Uwmzi1eq0TbNQONK4kCx6K0
6j0WM41CwdhOQdIO565DZjLnbbGDHYHxRLC54WcW6a5FeRVDZFRoAyMK3GrkzKwy
66Dlcjvwz4FLiizWOE4m2uSwWmKTBy4dmHjkYsUly7CBdcGfbRg82M47/aG4TjH1
IfKonczHCiTBzuCwHqP1ST1XFv+hAfa159r8A7G5TCZxHehh122JniVTxEaBMtVz
FT749KeWxx+YuDdmFXtYVCGuUiIYLR2Ol9MNgjVmyFgkoqflqRQuuH+aEK0mRgDh
HCCIFUVnm3ffaZbh4eydEYqACI5oI0ChV7KUtjc5/O7ISl12i7R/5y2RrctebiJG
rBUcYC+t4XWU2Aug1WZu7j0LkNyNDVjIWfulF8nGjxiNQxBbsuubc5VcmtKT6Ysk
TeWdBswbOAI0h6526iLWYdroB1PCOd9sWp0AolNpTap3QMBdbemSZr9vzJPtuYsa
OL5YJd0tGoO2FeJkljPIBC0pFjtJYfIBg5L5L9uq+uY5rNrogRAuLKBuFc7iXHaG
0sMGDfVTiHY6Mk2mjgsPVHiity9IeXV0U7nBhNhNd+GTAsHfGZ+Vq/lr8pYR+vnK
Oj1Zyx+ELyaXe8F2dS/Dy5dofJZ129uzBv+1LEQ37gqnjxj9OSJuKIjqW1LAaJlN
XkMbhSD+3lRVQfIfmoAKKV6sgje5FdtzRrxAVkLWTYGh3SFs4qFNUQgNuZ7Xn8YB
qQRZGcUtlt8YrB7FGKSWHao3SoTS09sQLNmZ4EJbSP7qBnnlldCjJBmKGz3XBnAl
ZrNoI605mIfZZhEGsdsoFCXGCaR6IQE7n7mdtYe2pZqFj1mVNBbp2P+Yph67nx+1
odCBZfRyz4V2wEfo9JiSvuadnDnP55ET7XQvR/drC9kD7MxB1ncofMDRhJuO/00x
8ocsbIJ/qYhfzcoBFlqz0m6eRIYXsrChIf/AWT+Zcjo+o2nQ+iOOsdO5DYfpf09I
0GB/et3+2R3PMf7Zlygu5r+lpxZX0jGyuOK+WHr0ZtqJJEIAdOTh0MUutTNg5pQE
j8YQU8W+yHo1PnyquMxwEo/Sq17SrJopIaWykl7Nz6gAylprgFR+ieWs94n+cpkk
Ja3GwAPdKx17CNthamPLvegpGIvAsy/iBSTV3Vn9mNHRgBPmb7hgHbhHaVZFLl1N
IbQfnPW9IuOEW/a8vzlAh2OPJGamusQ6qDSlXn1yoQkvfAiJTJPkdbkVsx1MCkv7
ksP38jZr7EKepWq5gs54is+ICTeu5DMh1UqVkS2gnAoNXT+sWtmOEa5uJT92Gk6r
zD54gcZIdieVMkvEndsPLumfk3hn+RbY6cvOH12e7c2aLTVxRq9/X1eyoDXoUXyO
McFG4yxidXqS8fpwrEF/1fT13+yy+1WeQNP035TOcZipoZ/EYFsoSfbeqxXWhZon
JQJcEPMRhmTrKbk7KTPLnWBZlTaJ6fGej2ntVr44U/UoKh5ZIIhe0DWMCf3/bQZT
wUcV3+YfCWHQ2HmVcj9IFauIxdTRi0J/smSnxABdoTuxlipR3Jl1fj9jnC3BE8Ro
USKZLEhOIo+uBAlz8uqVyocIeMyhMVRj1cbQTyD9MEwioDV0EOKH0vi07Tn1tiJ5
qbU4B8n8iRPXysHUSeksM6cdzLf2+9zA+PONa2SAGQH+eLUI2KbQXXBf6tqqyLPF
oT+dWtWPtb6/ryXzLeH0o7uYOvcpglR6ogv3a1T+s7J23h5cDr644Hd2iWGkZ0iG
2gKyMtLR8MThBDH8b7cMjtMMQMaWS0fPH18IQ1qvghkN0lMt2UzaeZB+lowzeRKM
kCvqKV5SjUSWfsq94K/q8g3d3OdysoaDk5mfwWNTBMWBKxhXSDQwmh4HO32nGRB4
CLeCXwtsHS5Z1P4ug8Q1IBsZOcZUYgoG9hbz3Rjxt7NrUxAFaq6m8DuRAU1nQ/RI
ndTp4GnV3e2kdZHOhnXdKWGmEMn45znby+hWpcuoaDc7XIqzx36v1JLMfWBnxl35
/xuJctIndYx5+i5qK4gwMtWX87Erri0+72iHHnQhw3hKCp8Z3+2PxhUXnqwt2XeS
3WKb0Ve+Bo8wUzuzl/HkZNheT+Zeil7ISAVOn3LK5Y7iPCFzgVn3ykd5gr2xFMuE
cMIMzNyfhB9gcQyh8zw/DzL2s4mJavXOxjFqdMvOApJe/ZmHVuBejru2ZaN2cOPq
QuHBzEkfT9Z/xuu47nQgA7ze2cmSXMn61uNN7dGX8p9wXeYCNYOYnRbbeeiSWiIc
GtgGXQ+lwDHH6zHkdJMll8/QmtDOcejfhuVnY3iRAvl6fxo090Sm8YA1aSlY3HR1
KTm0R+ERDkf+PLuGT/7HyYHEnGKmwW1ft8G09o/ceOO+yLX4HfFT5NxFUDp1ISgJ
2SgpmD3I3z0Sm7n18Lfsm7P3IcGaecyA/6j1qqQZJS/wieGh3VwuFbh2EOs+9g2m
4Bjfe8OiEmbCxiSNvye1QxG3ocz4nA7BtBi37SmuIyCuB4qiRCufBNO7N4AydKeB
3+o+jl4XECC/pnV2G4HllVL1o9mxn11vNEeBfGi9O7a00kFMJiVlZ2AZrf/jhi72
G85ucIb0o9DvefSArcLf1wk8mImZyNlElH1RoShdFqgdm7enxxDflIQWd+FChHYc
kHRjXWCDZS5JrBmHmv/AdQzW47d5RKiNS1eLOVYxaEiYTkUSBM506zIROjS7cBuE
FG7DBLC961hPZmI40cCEQ68WOoquyeOJpTzxyGUmnpTIpYHmdAkXz2V+GjiQT13E
pl88pCQSBVXc5hJkNzXNOXqzmIWbtiVQkPXoZS8k+5/Ghqb4PbkLVFamfjS66cul
PRprIGgbqdI+0+D5Ug0MqZEHOj+TGyXHBejvq3pd5ReHHHpUO8Y80jBAFWgTyS3Y
BqGZIczamPBqWmAE/12JSFyapfeju2pqlEZTwdKwjaFIBmEYSOyBfCHcSOys44sB
CUUZSDJXIsbn52zfSC79aeNcazzh1aqbLkco2VLXPw4ppjadKvgOBCWEXbvyw4yi
VLUFHb3+losh0hAQMiyXwm2qiV7edYio47Gx+GLxglbgvRE9mI8nOPGMikM4Jkiv
8nXcUhnGfeIXMIBYW4NJA/MhAv5LPL4QQ8+XiFQWP0Omzqx/gx0DTvwai5w6i9Vx
a+AkUwxvjg+kl/jbhU6RMMWNrpHHU69tb4LThm1Jx8obVGsJO6skYsDKdaQbXuAJ
0lNcrWNJLj/Nik/t2YOV2tM7PN7V9RnBOz4a/BxF0Cue5ClQvyS7bQOVCjSGFuE2
z/CtRy0Rqeg+OXOXJmjMF/ovTZshEsJ5rxs2AwXjewSUbS4wp78js65suPpFkYQH
RVc5FqM5r9k7S2CzIwyX88WXOqVrFRgh/XUfsYQYmW9YBzaPDMOPETXZA6ojxgpG
0sarHVZEB2zpmZvLUJewnYgqJ4/nrzoTDddWobmQRaTLa0PLMRFtfrJbiVfOarzx
Ze0VSclBcYKPuHNHq+5rV5k6xrP4nfpCLPq3Mrvfoi90Dogl9Z8NFKVU4UXBg/ry
yFipfQriov+tscByO2QwfvAyiI+YZfvLifsh5PZ71vgI8h2eedMAgEcV8nTrdM6I
HtH4M+GikE2SKOmXY0bFpmDWIZNbgFpS9lrUbTIMwRyJbMEazc6zy2rAZLhU19Zs
oMigFowqHcoFjiCEC5o20yGicJjDiIlkQ0FNTJt6K4lxHQmCE4vHMVFr/v4xris2
MUXWaCHibQYbKI2oTuqBRE1lI1bWjqZUKBH4ioBSZYF6Mm1DXMw6dyEC//hqnrri
lHUsUpmDlI8yFwAHl92+K+auc8KQS0sWtYNng/oHKDWFrA3sOSqdOCOTLGcFM885
DadWJRdbvxJUF/esXPAAZUecbdF0q8/lvfo0pEWLiyWPrv5spEJgcrcmsblpdeMQ
jmcv+hXsi3Niv7XPUsw/VsxGcxXaHQsGYBmQ8yVMrZ527Zc0bf/VIMR2rmeMvGp0
p8r3XyYm4TsYZzT4ZVc5Rf1t24kFWQOG1+fnqhNQqoZr7dAA7GupsqhyF12lBOVQ
an3LuNdFPu6igVvq6ig5RdDIA4/vDdBcHnk51aWAimxbp6CE0MQEkH9vqfUtzAmZ
wXaVUSqXvVFX6BZIKqmHlhnrZGZmeKNFz1Y/6CWcf75ioT4Rs4DiLT1tbhqv8SKp
bYhseZNuTfWXFL2dY5twr76j+81hK00U9ivrt2r8j82kzkRksb766kJ3fMIhwHlO
i0R8jO8qMBSYcAWcLsjrh3ZAzytcZbI2x3mOtGUSTmxlpB4iw1Bbk0QOF2lYPIER
k9K4Wlyq8C+MgOBqXJdawdIJri1Z6bgbaicfd/Szs2FEWYizU90JIr3xvAb2WO4+
/F7s2Jz2DB6wLRA+/PpgEL/b41kT0jbPp0+rUYQV8SKCCha4kfIopOZDOh1EULxi
RTJrnI8wZJraiHt1osfZNZYIi7WIdQR535moc24845lpdHWoP9LEwEaKnEF/mRci
z6KdqLirlAEVgn8JfisXwlseD06bH8uzMltoaMXGl3u59AZD/uOVOpw4lYJuHNqG
LPsbG+M84fVoYoUE19NgK+Zp1J9F+PrMnP71qeJvDvTKL2jE2sXry69lhT8h3RDK
5W+P+o2me2CMT44nuvQvFoOuGJjNYGBgZtOLPyw+lv3ZMl+bRLlkthSOPNg59NoK
y+rzA31fHECFNphPeI3eLYisQ1Ed4JkjFUBKJND2Lc69uTo0R7+Ojj7+uDuO8y/F
O3tYN/JoRgNNOOi3GpiXMD8cmRLRnK/DNMUgXTP5qfSBJidrfY3hmHqm9e0Lh3xn
WmRq2Rgw/Cn9kqp0+kK8+ONY0XTcr6efod0u7Mt8GoJpR0HUQ6elRV7Fs4e7uVmt
tlavCtRXY35edDcxDCwHfNMjpKyCmSEcFk4K8ZhMjsy+kqrq6T2O9leQYMz1e5XK
jKPK6rUfUMrzs5Wjn8GWWESCAB/z+NfuwbkAlGLUc3UKc2oXBBtwCcQogzroNDJF
h8Ho9TWzlQocxAF8dbGG3yicSDSjocnqS1WULlWAJrnBFNVhwoyyehbQYzB9vFf6
lCItOuRu64Pw3vlLju1bTSPrZhm7M3QcxsK1l5Pg0GcwzxBmRAM+jZfYUXYWoUUv
UBw4YbQadUSByBJdl3s91hOO2Xnc8Rkp+V9pdWtYoJP5gZ3zHCNAkL+M+57qT60A
E1nnwo+gXfYHlQPemGUoyGFuhrXgwpbTruFu+3B48c0mZy78vtm3b7je3a3gOYW2
Z+CiBhbIbl7jJdp1hkdTUk3aJBaPedutVopbakKDnDWPVBCJA7ZC4rSTYrFMRgmR
6KK0PfJEofb8jflkYuGYM5V2eGU2mP7FFsJqZ83e1dlxMrIN2BJsPoNzUpRrqrIx
y2dISh8VYif8fdTDV4Q13thpqYx7gq0vFxx9VX4VlUPVGhBFH20r5pA3AJn8QHu8
ynzO6b681Ulxo79mPeaysnNjr0H7Mc4sB5NvNV3UAA9GAfQzBDt4jGvZ7L0//54Q
Vl++3riep3dU0vXtixcAIgVGcDAlsyt96hRRj9uPbq4dGcFz3QPYzI88CkpGgqhT
FJ7ciNuIid+/Wed2w21BzCzztVOp2mVo7981WwcGV8TMWz/EI7mXsSr+r+ldFxzE
+7UfGBmqTeFYa6XmPFB/f9RQNzRPi3ZT3KzT+4BraDGyaCCQcigRuAF+fJ3rJwtB
SATEybY/DLhFVNZk21qSy76bJ9U7S2/LuTIdwjnJo5nhbdH45APng0GeHWYDGoD0
wD7lfRcFdUOerjB4wQXtxf2XSTd+7QWZFKnVaF2LzQQxwzihKMdFI+qhd1pWO59e
ij05ysH2o1gic+e7sqs1s1edSlaMczZyuI2H56bkADdOx+zFko94yEvs8EofeGak
BmUWVYiFQqgW65CBkeSrvTB89mVoQ/Wqr0J4zqFBMnwg2WYByFMXe0mv8qnf0Bkz
k1YpjVbeP0hZkCevGY67khidru+PJrAdGydwZKxtE+23R8lZet5cZmTcntIJFESA
KXzWhoLCWt0oE1iTL9LVlGale2/N/JbHcdJVQMy5e1XAIdjPrOGR6Q65M5jKxH8W
9W0Ap9v4TIUtbZ8f/doBSX9SAD7Y4bEoPsN3s/Ialepa6sF7+kIsqizn//MWubBL
nXoQsGV9xi16ji7aj29/SCTySvpFlf4DLAEgnrIUbB0AktYI237ZdUS2jVhn3KQC
AvXb5bdFFrqwrTHKqbo35M6Zn9z/4XO/Dj+Ro7PbxTkA9Igoge+mBpJX5te4ZUWT
/It67wH4vdBTshMNyyXuYtOsN3mRG6QIe3XSe23FUbJni2MrSCX8q6B0W+HTr1VS
wWoSBgZ2upWnwMD0B/clj2lxCA+ziH+s42OJ+KJYXoEF8ZlCZ3zODkMY7JSJFmGI
o/MxoHSoLQpNCGcgrP4LpLjdK0yItyrv4Jqzx6a1PwxDCrNZTHtzHTVXRaz4aZWC
kI6Zac8aCNS4gqd4SRoTdCvptHw/bkqyqKpNxw2X7c4bblsIj9/JpOWhDwGM+thD
FFti+RvOD0Ufg1W9gA9S5Qbakqs9nqIkQU4hos1MjoXpHgyC9tX/DyO2/bH1KuPK
uU7l3vhKJcAfVdUljJmZKh9I9ElyxEQe5y0+yX6Z8r9o2LcgrwxjHW94IroaG7yA
gI5tisYjchbI0odx/Vmp5MRESe7jdDegeUobU2C/inGDzjmf+waHkQl+pHkJhcx6
uH6FJsnxlRzqiqWkBaKHas7t5FeQMpIVhyUpxs9SRLXcrg71XltuGC54r8nAbdpu
+aUa4B6LRF2cwHGeUG6qyYDjJLk3i1BwWHWH0jkvonw0Q2Hev6Blo+bAseU6TLfx
vm+Y/OLLam2xx8J8UnpB2SqqXjIqiWK9X7mUDOqqRR9Lw1+L1rPHeNDxH1OmgSFv
kN9CB1O+BKtQnoQSNNOROYsqoOEnU3WOw1R1qd9KEFxtjook+LPrKfZ2nYFZggXD
Olfj3blBHNL0P3wpj/6uocC5B+Y19s0qGpJ+T3ztkF3hyKg3SjdxVAoixOJo20FW
0sBD9Dve7R5CMCZWS1gHe60DXEdelkYod20s6QyXAxjEVACzTDV3gG0drwlI7Bhs
Lv6krZP+uJowOKPOkv0E5i9PqV8Y+IyBF9A0JLIV9NB5HwDCg4jhmVIh7/txRk+2
denSHs3Z1cKEQUgs0K94kd7OvAsdwWCl9LBnRBDOLAbOsA1uegcqDqVmRGPWpLeM
0r77IyIoRBXGyWfh3j4IQrBIRbwiiIjG+6tYp0Hu0pPOacbLIwiZyJaem0Pu90qZ
uouLBrZNIzMWoGhjI2PsjdnbObuW4Fq3bTY2yHnqbMbgap+mnwu3hWXHAEJiUAp2
PjnSXXfJ+jqnlQXsBpF3qDo4XaKNFrZPmRkSuncS5rb8bGSK5m07AN49kRcOE9lw
VqKWU5zhIb2W2CY6YVulcD7vlwsuMF3xl24btHALN9/wIyjKjEhTXaAJ0XrbKDL0
cWYkY+Bj/2QxLNx82hxyxNMm7RdyRaZcMnzwIIUfuXtMb9Vvsa0GNSsiZv9Z8RpJ
3tjaf6c/FuiU+SxH6TPHSflXmN+oZLn8bf3B9RxFJG+2muu4Bf1c4c79yT4Fho9k
GGx9FZUk1QMMMdWHb0Qm5uZEGLvoHOfEJ65EvzPpN7Zjkn3F1r9p3KV9YZdMJI5U
fKT6WMaebwr2qvMLu8XS+MXTMessGFQs4FJDOK/WR46ytsq9hglUACxa0fI9PG+9
+1sDTj43aznpt7Qoov0OfJukdviQjafxL0Y1t1C2DaFCvv3IAgz26L6B5K1/6a9Q
qP6eilkpNQ5ZMVTgCPDFoFFdpTa+0+YZnaLZpOSV5GSIsb03pYktyqS517fZ7wpj
itrW3XNSshoK1VGZgTQsHPLx1Vmnp9EG9zoYyvp2Hvvv8bymc7orUVtOiXRCGUwS
961LAuVsRGcLBbz7eUnu/6NVOXdqlcNcBCoFv0lSO9VgwzptNcg7vkJEtrLznkEV
dvzuYjxZHA8BLUJ379g/a9QlnE77o6hIOr/xIqFRa0BCFI7pbUXVf5dDME1PL2rJ
QHAqgHL1/8K2LBdOFXJ0ece7vIn83US6v4cz7SEk04f6H9tW2ZKXfoZkdxQ4cy11
IYePQmJO+PPOkovnWMbAnYmgOUV3Hoff7QRFXTNfjyFkxLYvRqIEHBb/b4U3UFiI
rVkVR/XlXbnivagEMMixk4RtRHmz24w6xypn2tZzma49S+sOFH9Krg6A9IGp87/q
Lntj2nepIuEFzDfCLBqwBs09lKVH5cGOhvOvXHzWU9jWK0+rgfz1s2yAtdSjKf/a
sOV1o0GEiwPyALtbQyPjxgkXeh7T+yMTPYxOZrtcmX/GdWZnTWTTLCeazFaS/cIG
0LVoocy65Q+ftnRfjsY++hdejIpvgAUM6SRIG4GqFeK1lCFB9y6N1BdCkxgW8Q4o
rMT5z4zpO9VONzd4osj6sZag+o0GZBY7+C9uX9ZUbpoemqwUVUv5JnoEDivgJ56T
Topmwovj5grP/fb2SXG/5uxHMdMyexsx9Nxh2eOc2Lm0J8hVtSXg90Jkg7wRQoD6
C6w7nWQV1+9unudee84o1jHQMwDiPgW7NH5wev0g1EByg10lEIgVXmp0jwQD2QXF
GZDDQYlatDsPC1p6t0CrHi2xAdHcJsE/BxkA+AaZr3TKWJfrCogxeLHVNooYFVpp
nzMM/8jhnSaz+rJJUU9a3sHE8vySBWtOEO4fjcMOcIyHzUg3mKFdtQnpitgallUv
tKDx6/zH/wNghAEQroWbM1TOjrL2UTVMbo4wAYJMARniin3/A9oEtHlEiVJXzttI
81038bpzzmjzL2juvE0Qofp4NMQeFNSCNOUl+yQLj2VudMWEPFnSEt2ht+3K+hCQ
n02F9mcfgb6G3N1dfAuwWJClfzfxU4v7Ri3ANoP3hdTUCF+OfZ5nMCQ7RLL5vbEp
mTJM8dPZM99nfLBTNcztBKRJMQSOPaYAmU+V1mYz+gosyTNyzqkRLMg64YsWnsAz
4TIR+dDDua5QgkBeU9qp+/j14Qf53jyxXHDqEMiaXOs285AbIIokyIQUyNBVlPMK
T1czBZh3EltURqktZZAQ0nnfzxO//DEaZDBYB7FCuoPPasc2jD1NtjZmtTpnOZeA
AO+Sa6Y/Ovt0aCzETZk8uNV3ul0dXM0bVhXq9NBmjFWvEnkj4WdPV2KfU9IWlrTW
w4gKk+vAD+m3Cqzm3ynUfylXU8AMjziDylmoUE8qtBeTZebVz5NhTJa3In8W3qju
MQhgAiaY2kPc+2p5TexUU/x/G/eiE+AlHp9y+Ywz5cTxRDWtbSwg0owBSC6nyBxu
U1X55oCQrHABbNROmvqNflBjyvRCXVxeXutEH0wD50rUdTDMhWuMi4JonTgDoueW
huQTv92Ahyf71p2aMs55dGFp11Bba/DD8KG70O7Avo5VXSDrdakMY4xJuAf4hHy+
FVBu3pO3f3yxeVzeezGtkOdatVhJrN1qF1SNlgS1yRSCIom67HOlEfH6zueCRvN2
fOG7DbYEiPjvdu/YTl/jk6u56QFnv+7v1GyWfmBIjMCQVQs5nkvVzwY47m5z0NBg
LV/QmDSEAyiInZpilz3ztM269fulsD0i9hvwxkXtF6Aqpi3iGwWwRbA0uVdmTQM3
rgJQ3Oe1DUwmLQK55N/uMHbvZkMi2LkD6Db+O/xau5qcPfZ5uWKpY7saCmkQDN1S
XtYt3KfxHGeccDbwopHb2KNjnYGcsQSBfyIZwdjvM7QGe0KSTlslTd3iyy3NjYLM
gruM0evpB4GdTPHcS1cxyl1EA2CUoetr53XWqjemnA2Ujt36cjtY4ktbslx2T/w7
CxvpL9jkTaTipeqslWo5MGuDa5YWvleB4JHcYOsaphR4aiqw4cIIu3CA/++1UmCA
3Rq8VepQXdnEgbAWFBGbV/UXEkO3DhSpGHb8yn2BIrxw+Ldjb6amNLW+3RP/H81e
TwuYQXIlHo2ju5HgTrhYTnB8WdJ/hFbbCzRD44JTTwnBxgV0kjv/Qr0PnVBJq0Zm
6RjYvXSNUwMBppmBW+k4QEYKwm3Itl6mXhY7RYGZPZOzobM3OQl/uuQCheK9eCV6
mXzFMROENZFes1PucTCnaiF9fi2FGslS6xvPIXj37pxIXcog7wvNTzpFVK1TAgyf
o7R8yGVUH7PixKWoOOSp7wpnS2RD4JClfC9zulXidUEz2Jh+jP9XMWWvfUqX+1KU
5u334XX5GRlEelTc3Kxg07TwO3zm4APvBMH9l0nP65RfgLt2couW8E7Pz40WCXhp
E7tkjV2HWGk0FPqaGxB80XFt1vmtSjuSdHHR1QmNSMSj4iLVjuMJ6LoxdQ0Hx1XR
1im1rEbycvE2mZeM/fIwQfLli9OSekIF9AwdlaxlooiGZz9QzvfpwLy4tMNQWbxu
fRqUqclBnnKjtg3lZbO9TDcA/kq8iYCTtVRlXnvkpZlvQwBiiDD82TkIhPKmFeq7
NaUhypKHIq7RJWYd/GuZeswPFM81cSXPfduEI/Pp3T/w2wpXXrFyiKReOWcLDRrD
1YhHxsQ0843Bmfy36ViacQy899BKMFtbrG26jgME7w2/PfhvZs3ENXSQu+80k7ny
j+3MJybMOJEPLaJrWvX4gXhKGR79bYRrpBYjmQC9G8jgKsYyEFGN2rxxJnjJw85B
Sew2sjWnaf/BJ76wiu0Mm03GgoM5IJXnUpvxkYP6ZhTjSK1INXE/asLwe/vKA0tC
Dc5GDbtT/+KP9VwVGIMHNDj0ezJd8wFN0bFNMl4ii0lJqISB8MQt1l8UB0LJq0hD
odSN3ZuaSRgRuK0aMgQKbEPydjWFNxzJ1fH5gjD7ChWkAD0TKnSeIcVaEQp2blvp
oxnEYns3Zmy5Jx+VofvW/oWE4HoWmF2zE9/TXiZa+2QeEqi/6zFnFp7behqI+SOH
Qi6ag+m3KGmYq5pJ2FsCtQX3ijzVKBCTbBkXoP8/hjfNjH/adV3heI+JyEGYhOKJ
b6XyYgMWJqHHb8t5wigFBGdfmWSarjjKRSZzVn8KAfhAYjEf2ua7nwV70VVxqn87
oppkggJXhVPOo952Ob0qwW94E7PSvn6mCDCggc2nOIcorjNmGiL+KqfaHW2JGJXV
k4ZGiCRr62GJgHMP1mS/xBVDkEWLEysdpUlty3/tpeaexUzJs5bVBHC/q/ArTzw2
pCIgrHegC6J4MgKoDVJgvy/1jmP+jtop4zF2TkhOlZyWyRer2UulJeJxMk+wxBNf
nFjYRBmaphlNPOdjMVG9cIUp7KXxBU8cUyOBZFdb0/1xY6j0+yfaO/HIfN/uqeLA
jadb9ynO0IgEU7N6VXC6VgKELs/k81yISbjpqXFJsh19+bi4G+Uy9xv7uVD9tZiZ
fbydtXV+4QJj9F9O5UmVJLTOQi/wS4XSwQ4zkvrKLQLC8mmdIUE5UCY2DxHMHP1S
mOu+JXRyceXdxFmx7/L2lLbQpzjsTg113GQqpHLsV0UQ2YyPRnnC+mChAWOd2Dsf
x3LubFnaIOAOla6FH9UtTaKlL75EjNFRpB8CHaiVMTTUC1OabcBpPcpAoNlmYkJz
aQ95bPBpY9W3ZsxOWGIQqQBqDydAipDlWT5YVehPMIZ0EZ0phKxlnCHUCkotIfI6
BahyKdezvctElTRkw11HLoXOg5BXZDysy7tjlzNIBSAXh4u45/vtSHAxvnutyzRq
qxzmqoG4aMj/kKpY8oaNTmtcVjo5wwe+SHg0CKSGB85jHa1u8QLJ4YD6MsupBTQW
RrCSX9QqtArovA4kcB7UrzF94IHEw8MhSNv0Tiy4dJo6aKK2udYGy45/GUQJrXtP
vTBsnAG78ey47UIhEBQDRQU2fu726tYCrmYQOsR8dAvsi64zLqgxtOKNfmPwVx23
IjN3r2RAf/ChVXFfZvTqldVdGtBWDO4K26uIKh5XGNZNn/CdVaX5V2KaK8xWOCrI
WPFkuuD0T7ainmOwWFFSb8/kHCs8dRF44aXpTjYpVNJxTDwy+0Z+bzZdJp+Z2jpD
HT3v3LtYzSmGll2mzjlu84E/EOeHNdTMptNg/2hEGhDfswIX45ElGbo+p/gW6CLs
LgQuafd/v/hM+GbEIJJXC+Xaps/RUKgfpIsaS8So1jjReR20+hKZr1zIYexeVRLe
sF8Fbl6dkjl2GjXCOwoDyMu6c/OAFjXB41LoKHg8yIqD4n26mZ48fohqU1w1mCuZ
R8BsR3nmxpnjKoEz/QboHq0zZJQBLeOCqTXTc6eAbd5nIdBtRhu0uoHtGjbcbgrQ
K5am3R58SJ0u7z97msCr+e5J/2cXb7CqNyAqNbeQJfLl4mZodnyBsc8ndokCUgG0
/k6rgV+0XogwHB+yMcf1bqvsC3vIqc+EprPgmmJJ+upQ0ovqeyEcq4hnEAV9MQCI
ZrP0+ipmVdPTtHAIKieNw/Mfr/RyGFD9t4smE+4KONhnyPOlpOpYElMFwHWLYPFi
f1NzhmcV+wDwh8Z6zB55W9SK/B2aH6Q7I1osINbDAto3hPGYR+h3aYRfBC9KaDra
JigQQzeFKfWjZI5fx2GeXM1TKqTm8H7z9kVJldRlwHOrTFDX4EpOv/na4LOZwNrD
7u2NmWWa3Q4qZY3z6edzWWN+8jRr/6QhRj+1e2TXUbpEOr5eaHMpmy9Q/+2R6kot
H5TjM2ufprNCyaEYHG4CMukMQ51inEdOrB4AQEjqHPCvPUqL08EQmfGV1czdmjuW
fCWyKvyLGcbA6VpxjohU03TER+UYEM1xtWbC1ZxPIPZmoLr8Ps8V0om4harV1/Q/
5CiivcCY0zBF4cHqLQM77weIM6DPyr/k9h9WW3iLLvYcx9YKW3cl3JR0XQCnsjDU
YIX4y0uQHadBybR+6a2czKVTOywqIMTlk9NfVE+LW/+y6tml6+aOng4KgqXTI5OS
Oq2F6HU5WDGlRqJRK4pdMbgjftJOwv3MkNkRcG56vEgxONNGup4fa7PyLkHJo+LX
XaF3Rsfcg3nUmZKw+8oV9kkSbjjR9xRgG/j5rmPWHYdhfll6aFZx2EVhULcD+JUf
QmIkTAmiDJMRHMR0LeImvKHrMKWefIL2JmRwIL1aM9FdGztLoD3u7fM0MwuH9PFa
0QQTbNj9tWDk/GXJ+m9eR/sSeUYBbI+o5kyY3F+tDjm7VLHw17ObeEdVehgCqkF8
ZoOqFs0EMuWiZhGEvmFvoktffE1FgopMZcdUE2jExKvxc+vm+XOA2GgjonK/YDh/
a8B3sfc9OO0oBVjrg08a/rbtGkwAC6WdeikpDup+yww4Jy/2BhBbMxs47KAc4e58
4KHu0H55eAD4IR894bKTNpafq0fPKC1zWaYjxH1VScs7c/+AWr4qW2fi38BHvT/k
Rmt41P3Hd3SH0crh5yvLOzUYR3tgTv3DsLO1/BBGtGpTMCz8til3NlFR4I0tMinW
JGJzWlN1KXQntCpTliUjdcwfi+1PbsiMqtKO1heOEGZWSbeHJa5dGIBXOA1zKT2A
WFgzomV6AUEYXO3V8a30G1S33q0y9fFvH48iPJSan3BXZkLUvCXip2d7QjS2jSH+
eDGe7EdO7vCXu88lazyH0I45bq12i7h1f3fIspACZIfr8FIeZHlifCHb5tfgq+/n
ffDrcwFugAb2J6yJo9xumqg5f5ciq5vSjqLIKkInkPTatXlGJZlYdpcpMVSeIZYu
fluA/SR/rlqZMdcTGnOodc/qymtohRpRGTgFON9F4DWm9xV9PmWKM+cLk2UMgbVM
XlLyoSYxUYLXbQSiHL0J71JpXsBvJR2xkThoyDLrKDNQSNYaZ5I2cYIIl02KIhSw
Mg/Pdw8Uj3ybhDxkVUnnk8rihQOgmIcbFREWZlvEh8PSDctnT5it/6IVt5KIWAFZ
DnDs1bOnOOBpprqV5bd+Uh2CPHYxIjRmvaTSNPpzxb8cflZjc1kuJTXAR65BlHYU
BQFiyAwO3b+BrYUS0KTGXAm2BFcB4CAG2yVc5oLCBQUeyJVhm+APTvF59Y4FdBu6
XRI//tJrMvbi6cKpVYgogNZPOL1iTSC4o+0b1AyhjkosMO/bWumJAQbmSfSIuH0q
WZw9F0KBS01DGPB3lX6lUB1JcxX2wdkxsCi/tRE5cMytr6gZV7CYqMzUjgZMvCxu
ayKij308vE7v/Y3PfBFN4OBmnljPTng5DRDFkMLycJD6kPPpuTezG7qPtHQCYRP/
1kHlj4sxMnkczPFQQphyNXaI/BJvMRWdgslLeHHekmJAicW38t2IO7RF472tSfAZ
XcaS9JPrmdQ/DLWt5uNuc0OrIIulbKZ4lv9XQERtYizzjq5AzXxDtIIUgEd/KGup
Asn+/PXPoGy8iSMN/d0HMSyOviEXl2WiYAfrAwgo2kPl1eZVqJrasIh4tkvE+zgk
kifHHMzHTA8KU2WO7MCZkLZO3dc/sbxSiGXafjvvPpoAuL6AvMX6MLlal+xEJ7z5
iyt2oG2Fxe9sr+j/zmVPgT1QBNmHL0vfAZaa9xUMQiw24JAtKzYwUrsum/gWB+iX
ndegwo2vXOBAnLvvgeKbFhxBC0Tpgec7u6/+h+TUq6HhCzhHf9BJJ7JvGDOJb0Yj
NE7fgQskmSqwoXtpd5i+0DymqqKSiEBd8tlIujKBOO227tm4zcJdra5hurjxLXcy
MelUGoNyJUQ0N/f3chNajUK/h73xPH/Xr6FKBQy9/bVp0Q3/8/rCeeDwloX+BDQt
Z6BWJCJXqqmjxLILi6Bpq9g4sHZFVvGz1s5lxRpshJmRoKO9CidS2mxZ4EkVKFvd
F6TPlQ8WG0eB/hTYqTPFtwKqLUUeqwASCCj7pmvVINMZQzbwhDlOsVnb1H2cqkw9
/SEwHrcggiub+DtrE0AdqmSYKB5h9DYiKRfE/a8Hm6Vbh+WRbSMcHN4PMmrL2waK
2TkAN3zSmfAg9D7QbChdzmyyGD8/3w91QCp4KJZ+3CWmSE9Pe3UGK4cLcHPasQdI
K7FlwBobxaGR99QzMD9vggCb3eVUoe2Owl2tXvzUX5uWg/fCwCY27yhotOH52qvi
NaATzWQWjFPqfhb3pRTj7fpuCfnl1+0fyZ674OugmCgzUe4a515Z+naFDFEeygl+
4Sio6vWS/Y6y9S75plbYGazDqyLmoSaEEn4BY1EMgoNeF/X04+vlsfeEwZCoXHdd
5dhv7faSN7dyN/8duptxCsHOjaISA1hMV9Sth2I6r0/zITtp+qbtmePyPuJdSx/P
oUpes2+zu8cvvOuB4P/nURqUOmb3uEOQFXugIinUv+UHt0aWZPCMTYcuDvxA0DTD
2qQ1np2hVCpqYYsHfQHW3J809tzB0Y7kTuheHP1EqQA/eK0Y+21MKSWXgM1V56iZ
wWVcQwmJlMvCdUARNiVS5+rH4EYuvMgZ1ZUK9tZlZsn2Ru7qzYp8zybLfoqxIE8Y
EZ3actbkOHY6B8bijXkxjSUU7r+mYVg7gwdjDVAYy/9pG05FBKjOI1AX0hdgE7DW
ocLfPWlHpzpBug9TwIMHJSgA88Rd6jOwVMPlYR4/2tmHDxZFDIYY0UN9KY/go9+D
xhCqd7WXMocxehpKBXKLScTswmx7iEoAeCwSl0RLjCf/IH99bODVm5gVg0IKOWHI
i4tDNMQHVooKrREBjpwTFiodYacydOtYNeN0vONoErTau3ChBaOQbJc3fORmPeKZ
lia+Bt3o6zzCEMflOx2RZIevuAOm2EnxiUE/WfLVhaJ2ATv0Ssedgit7CSg908lo
6H4+9iKKj7pQ0sfxkgKn5CwBvPR6vvhRVeeCto3hHuxtsG88mLH6m+KbYvk3vg2g
6PIQDhtdDqIHe3mBLUtAPK1Jhu6RI0Nfkc3VGmvu9oIeNrhAP5n0QtIxTle8c3kk
55vNjSDm/esfeofUD1B2yamoWVMZnwirzbnzB00AlFr3qWh9yc6XSezcdxgmIOv0
r5P1qEkVJQd5sTpGckylaDZ8S26+3T/usBlXuv0eaY4aL4AX3Mdc8UR/FM+OKVOO
CUT7STw8JgWutMqpBpbCicq+jO+4Iql+nLL6VvVgt2s0oCb3nvy8hgScrp4a2CUI
vOJKL0nFANFkOeKIG257qqZhfF6iaFecG3dGnWO+JvnABXkGyovRbY+N7VjU1W1e
GFIq3EmcFfj8ZptjEz5thGyRMs7iRFkZRc03psDarTtLg2m6JLBndRFWnH/RnfWy
K7wW3YFcFy8QzGFTr1ZZcayw9vxPkD34DA3KxtOQ0hhZpw2T1JHFJZOjApE3vxBI
qOqF5ZJ0BG6koxpHgTuw2Up+BIbNsogDXhV71Di97xICQokBFB1MNt/+GGIYa8GS
ET4F329W0/118zLlRXmERBfMZ2I4eLQWdAIUkOsC1pfK6xeK3zH5X98du6SEisq9
Ywf6yzL5KHSlLidMOIg32iroaIJRoAulNuLPm3n6H//ej4wIXRUIDl8LfnrfAMN1
IgyTrHkoy1UbuhQ78kp5QNyxuglEt69mCVI8SycyzGZc3uSpwl8n5J8g/ZdH/VAP
j3imiJsjHWHkzd5i827X5HNiyj/BIp6YfhwQKWvVYhx6p7jGaIR4bvNePXCtG95x
KtUQ2HaI2dJSTFaLbC7EG1l5M878VG2GnYhNpghUBO9cWPs94chHwlTruKSuNS81
4+OYffhALlwHdqdWsK/41exvgeGlIdq7QuKeykYEeumQs4hsEBQvFQG9fMMVBmlw
ZCtwXsrAkIOiK8xmqFwi2LUEwsvepBUepe+4uKbsoIajdBQfPjHoJ9nL68GkJcQ3
FuVNlUI4gETwU/mQ2zEVS6ucRIfqGraRxeHqAY2OLuYN2SCBo2N/FZhEz8+zaA6E
35hum4bmTACfI6xnPjSk96goX5iTUSm6uUUNXS/gyMWDV9vA81ZtCEcROj1jnf5Y
7laC5QJ6gPtRBIh37WoWEPwvG0HoliaHuz9Ww/JvPUeudW8bTOptQSf2lnp/Th8Y
GAQYhvN7OyrrLcOZhXisvcoHXQDyaeqKzyPbjNDYcRTYQHKsnR1nfq6qS5Sh/hpK
epVS2+zEc9SQoABPJpWDFYu91sOj2RewJl1v2OTNg8T8FfqenQLGDbOXaK3fzhWv
Frube5ecdml6NOZdhNYJiTfCYtx/heFrgHzAlbL6poQ7QRkCN26KHFd9JfzomV5R
vx3LeCxFNfXfF4iba2IFsQNYtUjyWO7IAOsZTIBbEp9se9iOiemHmGxpVzENP3x6
EkWdnLP41UQgrip6E/ywDFoMUFxTKeO8/48Z79wEuUcRiEWz1GtqljmYj0vMcZ2n
N5qNCgQvofeS0T0gHhNaoQVBWOLj+fT5OAfqzDOgNSha6QOmWmrmu6t1SXDNBZJk
cXMrNBcDJYe7ysXlUXrzW+5+NpGrmMt5guHkO00WiyoZiosCohuoxX6dGxlRMcZs
FWnCXAbofp6o5T2QDWeQZ/q5i8pGIdZp3j7cUNJ+ZK+reYoGPsdHL9Ond196MnUg
9GBAhr3ZojMcM5wCIXUvjQ9YOnl4N5lxSB2m2DI0YiYi9oNrRkY5UjjOGX8U4EWq
SHANutygjO9pNTd7pfxoLA7p3tevyCUMqtJtHkLDhV5eKBRe2AjtMcjPB86Ejrn3
kTt/vtiRwO68iXIA8fEfhDm3Jrm6Fpe0qdVkMKOjsa/iMoytU4iiXbQJgQsN+HXu
6uqIDVHh8ZEC9R6N7TsEEqRg+9/mAOJUHTIl9aGKONPIYoS9v077qLcGMnxgl4GX
Qk/D/Hk4eyvu4rXzprP4dySZnzlF+XX2agM6CkBWTwa9EMdTexXeQC2UVdQYMMsc
T+ACt9gD1i/2hZCu9uowfx0wUygOHLindZn3ltJ5VKfy/SqcLvJl1dfdUEovOAQv
kiPDtTjvNWdxIOxCmK4QmCnxiEX6LIa/2IwYHGUBA3uHdpIvVdcuM7z8UHc5ZDPL
NFWPIxj2wW9CkIx4X64xxRozelpInT8LWQyRH0reaOwF5X6y1TRuxcdhUkGNAHMl
F3c/3rnoj0yBaQnD0zyXboWnKSLM5jebj6EiqH4iWhC9WNDRlP1hG57TLEpJz17A
mEakdC5ufuF1N2fPfGSYqEFB8SModCHMkUhCvu072TbsRXYFRJRD/fxwNxOzk1eM
N4czB0jVAncoIHAPgNNz86oMU++kXKuwAe7UV82ISMfPeBrUFV7kzwXMfK//AB8S
t3A6U8jSkLx7iuPpUh7vikeubUtP8VFSZBAa7pjQEdLxZPZwr8uRqjFG11K44Z1p
hUy8vMM4dSzNYhECkexXXPA52h8qzuqIx3IWCll09TgRsHHWMNT5he8vPdgGMCyH
zGREfbRMDsIJsSuZeWS8y61saPwiNIvXxkJU8fhTbox5JU3wV4VN6trWKQ3mfagE
SbDchZbkoiUHA744OoJyNHoA8wKiCl5qyNPurmboF3HdHv4c9v54m+/G0xDLqLmm
KLS2vkf6m6zBYdSYGxGifyJAwXtHsyeaaDXIn1tVfq59V05gWLghJWliBPHorwgU
mfSnr491pUPObzw1JP7EjmYu8ArFVWhb1rKPOXlwO+L+Hc/NDb/k1NvzHPvBNW1m
5N+RfhLvGxZqszD8msOdMCyHVy21A82NNNdSQt9N+Mhlr7bfK6zcromc6+eCucS4
N41Z8WOZGmZlKYWuPvNrPQ3HSPd9YMPwtr6SKQxGZdP50vvppYFWlNSJJPNm+U+p
RlT7cGmSyohRfv+IlocNOV94ZY2ViJTSbIUczSAyp8Ry9B3MjNsd4jSpyAu8u9i8
JU1JSSvZQV9kI5JHRZp98f+okhrE7FIvHe6oCopJVIPTFY1zVjqMsXvc6zVcYbzQ
vBF++tz/7zV7BcQaiDxxkI5LrhIRXNu8Q4BSMRehcMnAYNsUe00hrXSHPr6rEDr0
k+ECn/OJlM+ALb6yvxpe2/EuPahEdTOFytiI6ItrMWS0g8YGG+iFTez2aw4ai1Q3
h3rGVjRbrdkzC7Z+D5zPm1G6hNWs1X0BQTex3wI7fZ1VIYw6t0YK/SqHV5FMhypH
mFaCJ1CRE3hthc7rpSvpJLRX696XLSLfSPdzAQ979EWpnNt2RADUAB1lXCkyL+CC
xVMEgFpr5o5umX7LuzhKqtKTrHEmePsuVSsRI5feleKJ6cndyYuGe5LLYOPIYK71
AsQ50ruljSGW7ax99vkOREf7WF85XSRoHmObFsFZbSxYonyxjlGzoVijUAFfS557
i6omrOpJhUABSe1oZ0++4JG8ad9I/NVK8C+g9rU40+nYxrwDVU8mIxV87FK2vsDK
GV4jfI3dLKA75KZdrmPL8bAC5DaTBqvzNg3NXSZ1isKlfInNaO06GwIVcdpgrrxV
6NacjJp5eKVh/ZJR85d7eIe6C9w1Hq4m8B/fAVwLQrk2b8Ten8WF5pXRP4sgh2nu
9IP/NgBam1MVyCWFKYdmD/ppF9eUWceyHnKIPHDATYPDi92b/7043W7sFbu6LT+N
5X+5rtPXNnqUAci10rFU/fMNFfRcHe57s7elYeYPsoXle/2dBP8sBzFVx9+VA/4p
twFlqxHwS6Yd1ySz/phKrOmW6LAoYGaBfOVSqz7j7gZOB4Dl8ZpZ50LvXOyLtYwH
d0QoHj4CkC9tUNd/LOPwdFTMn76VfrpTcnbp0rrtmTBuPPgzGhbJ6a5/CEScA9OR
4q8O34oLQqlYRe//5Le2v2fxU72WVrVxvUyLP7k8b88mRZtVeYJ6HeRbsOHWVxLl
su8HAf8lJURCYiueoOSe34c57uzzQNOM0xelN8WC4gO8yq8OMscEiNiYOVwvCD/V
nUt5Na0BD8rdkbAeH1HSN7Jj6+bV2NySSzAyAQVVhd2A58MyS8HyrkcsSztOm87X
MtQVRs+qLr7a97b1gEz7AloVF7gABWAWqEwyOYxDtS+HyUq7fZxrFP8kJETs2NNa
c6wSE9SOqce+pJyU2JPgRZ+WPZNx6xUYyfD9A2j9/U5Z0gypcoDLTZX9+y6NkbFw
kQLzBqkGrgU3ba3m/QPElGUbwbvO6xdQPUGRY+bYTFNXNfNK1dZoxsU0ZXqr+0Pr
ZvbNdww+TyszhnxzhebRqfUFVHxhwF5an0kywJyjRaWXpn11GeJuFdJjeiVQchjV
Qp/Gj6ZtZFQyCQTYc5eR2Rv561O5hHZpfzrml3+Ep4BWnytzyJt/mzPUprHYaXTS
1AhFBxqEp/wNOwZJN6unfNUQNRXxCuKenCjDQgBvxiyGKVBa34LEMXxvyCdUIU6y
v3c/1M9QQs4+qoGHpCNs2LKxEpqZpVoYXbCM+pOKJwJqjrZrkEdjYk1JQgcUl+5e
r8uZOWsc8Ouq82cXVyn9UabPJMpetl0iPfI1sYlAvxCTHQVp7WcKeoWRmSJi7/SB
H73XXuWJgW5eDYQLbCEUxj5+8kyXfNNViGEMRkFKC68ZmcvXQoNFVxEDir3qUt6p
69gZr1qxQ5vTMETR+TGxilQw8ADm0fV4X53iJJMeYTmA/+CebnMq0e2VGP71QNAG
tAUhyRSe9s3MCAllzF9FSDk7u122KMq1tKmWi5X+X4bFolHS7lgI0pkXBvP4dad5
44N83UGia330tBegl7e5duWxqeeiWufe/WQTh7XErKTIoNx+g7Szp1EsXFBssSlY
L87B+q8siUplQ7bQGb8UkhScSmvsY6Nf+2D3k+WXZL6JHvHy4s+87ttOadIJnN9M
oHYqfn+HlrFAwmtjzm7Gg/ZMqcRdu/BWvkHaUvuKk+NmcJ6L3aX3YB+1aRIKZjGW
2PMcIFUkhJVY8FJ0Zg9JFonwOG29tiY+QmTEWtohwzCq0cOK+mkEylyZMPAXjnuV
GSEUMuyViXYKJN61560Q2i/ydl0LJ0WpNXn57T29H/5f5v/KSJPYWmoR+EMzYTrt
O6WXzs+/FwBzdeiboNuLSg3hGb/01y6ql/mhM7j9SYEG1dH0Y3SnK6YgwQoexNqE
sv5Ob8ySFvJdwjoJdaLcV+5Ln8TeDMmBA/+qs54BX1AATIs9qJ+/gsz1kEeyQH9E
Ur3Q0oOMitxK8+uYykz9rDYoRHkXG1lGy1EFaG42AdtcIIOwOCL6+Su4zW0ad7m0
UhocGOlhAjZ89KWjkc+4sk8EQ5s7Pz2IrsM/O1TeoLO48Vu3cS2wDzn3cy9vgRJ8
9NE6iIlHzw4xsSvITntoE8l9u9aHyx3h18MEdZ95bT/2/J9yluyaHnT8BCJdPP1O
nizEf5bS4Vdy32IMadnQk7kWWBOXyiZYR+qsAUtHXyDpZs5rdFbfr5txP34qvneo
zNOOrmsCXLLdz85bdwiKHsEy6gXboDx0lc2IZyHnIZBuMe81ZP5sJEbM0eepBk9h
NCqEOEOsev4IctdTVte7MlKz2HgDgn9fJoKbaK21/fedM+AIybaRHHcTRG6BKJNV
UWb5IoQDfihfvbVtqDjcHPpsP+rbx6K60ia1lQPkUKSNyFpS5uB/OiFMP1fMZ1BY
0g9z6Lg52gK4jfH+rluMdXeo57xSsPU1B2+L+BAQVy4aBeBWOYJDkRM/Ke4SGf5x
Qdb91ZK9HUVFj2qDkE+pjXEODFxmuNO/w4kBo9itpGHKsp5XIqG7xmvsN4jDCisj
sPIk05es3E3hZ4VqNsxlhsRXhtYGsCSTUGmh94Sw1hhxRdHKdHfAWepPBr2H3cN8
Rw9iefDrUNKeiDs91AnI3y0uetXdFuSRk5E0AA3alyiothmr2u1qHbstdm4b7vNv
8W9AiV8tacYar+FKkEsFXvkc99o6qo2RFCwCe2iIJYRTb8F7Z3EHz9pPXiDZc3Hc
mkRk7hLDdtU6h9nO/4V6S7a5ypuR6pxUA7FFF3VLkQJC1WrE9OFJDUn1eyef92U2
RcK+JwkJn7SsIb8QlshXeXF3e+4EnFXyH+Y94MAhsAW1Ynt+f9HXsEK89zPWDMXI
m7Ev9HC9kX2qs1EaNZJ/fNiaugloX+f4OlHwGCiCF/dKHmorFh/aTLuqAM4xzcU2
QhU3G6cZYvlZmgtW+Fougq6oItuGpgxAXNCmpEPWL+vMlRvjJyPFV6JnVK0Jbs6T
x1eRUjPE9N3DTrfbKxU3Eg+blNayl6PgK0LdgmXgm7SnRinzQVkXOxSaaYA2r5xw
AwIBfCazZLGb5LlrOfnImcj+CpE1iOAO3+kLj4Y8ZVcxN+LG7CFFCnckIrpeVXZ/
kBZK6iUAaMxLTD67aFPsl/Do3/HJvAWgPhnN/9KQg7l7kG6e8iNJhDUjaBPzYBRl
seDqXo8l8U9Hf9JwZY8kGssf2xSMoOMPWt3JPf+aRRMKJclEVFeE3zYM+HaFPr9Z
TiLMqFoY3hzcUm4ng5v4VuX8jO82FjkfCEVMxC6PAnUUMZMKbX3vS88fMeJtRwk+
++28DgU7SIsobSRRyIGkj5mRN2NILHbPGmZ2VaGb3+mwqwJJ9qrlgxzNPcRK8XHE
ksYbC8z1IPvDxxbzPLit/6MmvV85/xxLzga5fIIcNYxm15HBXQ+aRU4kpJ170Ot6
I5NFphtYs9xiAOjBAvUDS2b6To5aMe+uFb6mKoQjQ0bdEH7eK8GRmuMZ9LqulH44
TxRJI7f5QukvcZbimIe0LGtn3Jx8/LxXC3kUgYPeyJ44LiFa2kx+SrRnzakgx/c8
ATQnbMDQp77XBPkpWU4Iu/BRwqExznNURUtlLn4sILtF3YMhNpkR6Qmo2qWPpkIk
P51n2eOs6ZwlbigpOMmLD783K1WMM2mS5y0y+fU+r1mqpaQLPeWERsZwzp1iJVIg
0alt01CDegY8Au0+QditHEF2+XKAk02CVLLbTiqtBr3LXgkmFibglVaCAqVnvxb6
LfI11nOJP14Oh4wuH+w6VtQVyhmJSYLeZQUHa9cQD6LeS2zAzn9qsOTea6rR3i31
Wz1mJpUADKBidQR8+lHvFqwBt/C1M19To7FVygSQdbVL+SmNVBBmqFZPxZjHwaJE
2+lIM23i3Wz1JEyZrpXIuEaSB1ApYorl/ucW9SI/h0cdND/gfpyErtUWrYa2oB4G
eYiqXWnz4biG5z4C0gDQ4NeaJixe9/wnEDlwCG8orY+ThZfGwPWy176YkJh4EwRZ
7Ti2KsZu46ARAfqWMoM8v4x5gxyhzg0EbD+8Mcxh6bXyR8e07cXWm/FVVcOjJgke
FJQtqmw3JJek8/MPrgEfJDSVB06nScY1e03RewEd+faIoZ8dxZkeZXiS0utstFso
sUXGXyM2/oIr5cbNeYlFi34QXEJrzHWpXfPKpBUVw3Nid/oSwr00Mcl5SZcvgR+I
Tfvt6xNb6WYb42+vICj3+sXw7EeJMuD/a81ZkKBsLZsX04761RHozuys/ysJo0Z1
W4rYsJE8w5q1yAmTGjBHnpwzms/JpIU6PBlGa2Ui3/72Te4tGO9PPW5pShxX3HhP
HvmPIg7XE7X1qQdAy92kNlSzVzr24gGUf0iHfTgQsZp9QQxfgkdoNJ2GYUJ8LbK5
SoZL78hTlWsM/bFyOdZD+0KqPPFPDbDuGg/0Bsqg5hH8TxsYHhuAcegCu8yKtAFz
3VRpCPw3odEvyAg/DaMRAoq0QSjyYUig5YhjjldtmXyB4i7VbMiKv8qEZqBYSvRp
ArEAk+I8e1RBcVPNYGt4PrNdv9gMkfnPsJ8SkLznPxzJgM3r69iaCK1X6XQKgsce
11Kdl9QdJuVlF1Kel88xy4cuOi/PdVNgyx+R5GOE51QvKJO28S+zOCiTjrOyoNff
2NJdVISOKs0qV1rDW2kq3epleBrWF5wVV9a2kh19xkWJeO3Qtx+AWVfTFImV8xjm
nvgQ1lsl6bpIP45RF/ickO9J9un6U059HPOP1EgsN0XeJhQD1XWpTFGyRIZY75el
oq7tbeH61H2rcLy33RttN0XqCkPLA5W7cZyjFG8hskFz52xrdIexiOJhOHpRl1gm
i8j6jY1JRh4sVFjbUAhCaY36+QuHl026AJ3EVhHV7+G0SbkLP0S95hHZxaLze9de
nXj0b6D6r4Ukx3WO2Wl+lIguNMYjQKi9PuYT0bAtqQmm0dyPldZiD+1U3m/bILb3
QJ+CBRySpuChrUEtUikgKVuclZbffPBH3ydGxmA3fPHaWRpSTO5fs6yC4cB3Xd5c
lvoRCSYsIDNVweXiiaj3EI5KtIDb918uvRHruu3zEzLjN+B7uA45h52WOiXHXgXK
SmcCvSKo7n7BDwQuCTNsBKX3s0bMK8u/Sk4Il+gGzgcVqsSzjJ7iZkjg7qnaBxsw
yiBDhYSD4vMXWn0loW0MzHD31cHUlzqJ6XJOXeIsc/29cl5zveLaHqr8v+1lk+Vz
RdZaKD40MuMOK//N9NLtMHLMSjfZQ2IRax+aF6tHV4NSOwa6OKlwJQGb9DlkNONL
D1Be+UUBsseXZ55jo8TFqEoUBNEm6jFp9SfL3YHlH/hmpEDYMgQv/r0yDC+y8xMg
fN3cBmDptD8H0P/sL12kNg7h2qz8oF6PkKnC2r3YqSyyoosWgyTznFOfOUpMDq73
6BhycvO3XO4mDZhKkId+LuHr+ImWvgGB1TuYDDkoxbDiEh6T/XCCjar2GHNTpmgb
z0DzdiYVhCPnCzxClDvrxI2Qfri2Da+rxlH48EZBnQPeE9lpiNwnYTdOvRIF1ILH
eRbIGhVzQV37SIQZLapbRxT5C9p54c8FLFrKRmb/gaLfpPf+6yAsndy1K6UAR1AF
Rsyoa9Riss0YfnVRdadXCZnWrOKVhGm487PKnyvkHz6QMkugl8O32LcMQUGlhjsV
MBP/FrgdOk5poAuLrlRpKRnoM0u8RO9t7jrJL/tbTaSo0pnH7nP0sQSdZWqWRRuD
cfwbFlCqXk2crG3vumkirJKaT+q59gUJilJZ8nuq6N59Afy9Ruj3IlhG8XSxZ7Nl
7S0VsZOCxs1zfq48jCeHcoXrAPqK4s/9w7BgBNPeHwsiZdIAS4DY7aoIrQYu6Xwz
LWwdZNGkrI6SDAL+cxd9xMsUKua5/Uw/FBNS2PectDuYPOSGl2hFgygOf9JSKDxy
LqucJeIsmQGy/7clCfr+AW6AAtlf52X5+yn9EQceJPs6B3tbIP2/oIwJigfAGygY
BG6xhdUpKPVOEZ9y0PpQPnSwTyLU2iorUwXGboJ6e4DFt8XihhvvJxw0TEh0b/+9
XM3GVtzzNuseNzkbZLRxLqCN8VWW/+G88gTJAh4uZWBPwexg8PEKMoIEFscvgq60
6e+O5hQDTNkEnCrj36xqoIGANFRUht4NdJ5QCrqtl4Sp6keCiBy7c0dTybAYzSmo
HcT+m0LAXtN9SVXfEOUYk6AO/99gevdYKWwGKscUAURl6Xh3cgmsVqag3yZfLTkR
IwZnX6xiqLGkaSrg9f4sgt8GYOfmGYrkX1+i+rZxe9fiNQQs8h6SUbiZ6AhMyCnN
gXMESPCFg/IjuvnE2htYg/lSOHu8G0rVjmbYfQVybVbCELvsg0n/K4qOt+kFp9IV
3lB053u7sjPB57SG4aUSSI1bMjB9OJMcr39oWwU6NedXs5GJsO14AV0JVQOXZ9Vr
9QXCty5CQbMLhhwCbLcDMu98JKWUNrf1UL68U+jGIlvFycbXA8eK0VR4IdO5E85d
Bxa6iRT0mpLcDaTQy+BgVmPYFEZgb0EEgsnuy7eGxCRW7e8rlb4Wvn/JFACZiORa
fYMgRNV/UQE8GLAVyCyd9l8WbzO7oRvmjSGPvvp6kko70xujLZuOoMcjySwQktIN
RZBaSGOWuDtT3CvLRtQkP81JbIRvTVkU7oK1mfC5sFFfdiMPKAKWpTmd0P1fDztg
Pj5/OV6CgrXsWFzRkagb5fpe9eEffgjSxpZQ/gtbpgUE79k+of9rKvEFq2/uQl4E
ohl7NaRZkPGxrk0nNabMsuzWVTOpO7g2Lig/nZB0dqfDW+Hph9+2/woe7tEqTE4t
KqcM4+E3wknmNJVOd2AU+ZaIiLf38Ge8KLULZYd6nWXddyuzypWYoPH8sZet1E3X
i/SwbvPwYS1WuQQ1WCjKUyoqczpZI/IU0Stn0dqibbh7UGnLUFGJcMeNuu/DcrGz
zwVyTwn5nDah18nLHwJqtaBOfMOUbFR9Bywo+MsCBolGx+G83d1qoUrdFk07yZi3
ouDIwyf+1W+TUIc/hTQTyZkb7BVUEsGHSj5wWdMJYtP+AsfMt8oiEOtLP89u8rkv
+/Qzfxw0bFbwWpAjqUOTNVSnuMDeQ4SFUwcCS3manIgUafT0rEjw2azn9WBBymZF
OuX8+hPuKDQduiUx30eNl3i+gei9MOQenH0fQpmZjQP8RR9Pvd4G/KmJ3pMwvmy5
y5gvC+VnisY+D+u1QSVeq8/ATUljoon+d1j+kMp1Y5iAhRhLTVtNMU6Uul0LHZLN
FzB0ZqHAGhQLB5+CmfMn0PpMOJxl0DLPEmrbu4Foea1yuM0YO3qTafoqoGnKlkAU
GvjOIujZM+zsV6OTU3CkuSeRikYjD4788+xqUjGq0e/pZM3PgYZ/Z1+Et9cK8Ep/
8L69aaDKe+D3dm99wdnXfFp6ylLeQR6bcM+iRhJpZsjZURJo44Wob9GFpy0Eok7b
zK0fpdzDebajsWYOtdrQwqKwdF58IyX89tx6PNyPm2NMWILwOTHjgZa7i8ZckzGY
Xmnpw4Lnwsnuiwp9/ywG70FKGC2c5v3mXoaETABW+mBHPQljy25wuXoMB5QRhFg/
+JiNywASeAx2n11+qRU2tXusRWhy0rx8F5MyNKf2jt+vGrEVYO7bNze0cCErWtSH
2Fpj9ZGhKuzbSgDVKW0FxOyZMAivo5onFMUpD15pjUIeoxrubmx5FpfA8Heh6UsJ
vvdVSuissSkxAyAZssTn0Pw9WwimfGFWW6t/bySdp1+w9ai3DrnGBOAjs5bqpc4z
k+SVPt2WkRYLGALZ8FLu+mbtBHxd+wW+BME1vqkzI3InNqFSwzSkCZ9bsPxRxGhE
O3OHXdv4/CS+ZEXhFYBKG2nVPcKbkxx63FTRRCcn9ZiD3un2SQRCDW8NzDKYhvI7
CvTml+Q8SXIai5ZiNOLPb0sxSKltSHzwoc+LC6UEAJw4IBkFkMHNaezbHfc8917F
scdT/Os2RtHlCEqmQbjI2BGBThmG7o1dRsjyJlHahnW1ZRfiB9VeaAt2BCTRcN/V
HCkOLsTbN3sp7kfOKXxM0QkdwtcRy6C7V/9iAJUfaH67keQvJcQM+eSD8kaKG9Tj
kSh/i83EkR+eWQsRyKdHjMD/02VJ5v7Ynw5HLOpszueAZCr8PanxYdRfiNLMYMPm
UZxYsZBh2UzM/T8s9eARqodEjdFgvH1GucGM81i2Cy5dnhFFtQR6VjMEVnuHN8ET
abaQZKE2uEUheRuqQKvCqfND1NPBOpL0If5AwLyvF/1hZqebeRI2hbjC5Fhb61z/
Q6r+ZNhMw0SwgThVFwzjpemkUJiY6UIhnOWjFnw5kvUp4bVqNcYUPf0M/lwyIx/X
Pi0qJ3IKmWM/8yyIdgd5Crwai+0JWRTIPfvxrt9L6M5hqmoxborlunpNLOHHAeGO
+UiHYYzTBuC9ecSiD0ZJ9IitU0kSJo0B9U6Owlvl9uygFXb8yHXhpeKwHpb/bcBe
m+gvPFNBWsE0dUXXlyb9EryYjxjGeePtmS6sM4HnesimM4qmZmcps4kW7g4w5rnu
jZDsFsOQWxhFoUi3w9DwOE5zrt+NUBZmwxR7ABcq7HuGZpdyFsSSZ0Zawm8oEJg1
gVBw7KOm8564wjT+q5CIXgmUObuQHhXCWNsWwP92KV4nTKY36U9O+5AC7us7A5n7
rwtnpEHhfUeGxWH6QBEymWSabXa0gc7IMvRC8ul7kuCguHFWVyDOxrSkPDiGKUCt
dYPwstLz8Y4tyYaFVvgwiVCm/pENBVD9itDdMlsFJ5PnVjxKBsbOMdU3TaGv+bln
aYawgg/6FyMNBISQB5z5l+oKIjLIeFrzPE0Be9oEBAEa90P/M84rETkt6BPEtqbk
Blh0/mOkqekehqLpMpixbNZa3JOvaum9Tsfow0EdoWvamGyA7NXx3dtcDN0Pkbht
DsFe8yVrh/PDu2vaQ/NfHBSJ6xhf8Uoh+JPQzVsSpGt1LI6f233Pmjd65mcptpDR
RIErgSKsMl4Ipbkcfsi6X/Nzt8z9IlHHRv8AoC6G29KKAx308MP+nLdyeSvUi5uC
3+9GdnQ6anV78pzq3TY/Qb/RXKCv8KU6Yqhixaq5SGK0qO4jowWSQWqRF7MqwdQ7
jgPRE1nWeYKoqZC3VeeLIeuso0i1zUBxG7P/UwBoSlUBT/vxhmbuDgjt1LU8MelT
86y2bp4JIbcve74le4AJ2ssBY+FhUYTlclGB5MoyRVNTD9wWPGh0MMdTdxjsGOad
MSjlP/0ZbVii/eP4jxKK7BBq3lovzfvmyJBgFao9rsXZIZVAoL+3DKyDfjVEfMyw
I/+rJ/Q7wTcqC8wn1I61lijNR43QHWPYBMRp7jFsTlyBJmRv+g4j0OYXXp9Fq8uQ
7819EwVkhFgYAz8jDvp52nSVzLeyZ3IYBgZMfWNntvhK4/SrceZY3OMflmhpOYXJ
tvptBYjLWqyhEbxg/wP1pQininmuLBCehXFL01kBgdAdTwPG1xv+NMRbXkiwc24N
rhszFtzMWrlEWs6xOWVN9DQk5iNR8FilMKPkdZ/BsOGQCBP+G91nOpeEuvbs9OsK
SByMIzshqHrLYuTmdsiJlRdDy6L16TqRMpk5qN+yVWbkS8q8kFpYEFx/YGmYKHyr
siJlWl0XB8lDj9VY4Y8pPxyTZTrVkxCVNx/RzrK5VYfvbqyF6SdLs6P1+fs9hzTc
ekrWjXyVNpnhmp/Qyn/YSce0IxoWFNV8TkJNYzrL64SM/93RViCAbpkqO4DU1kK/
pDVLDPr2dB1gbGPU/HHcl2zpHnho5kwJQy7rMoYVVIj3zthkdPppxneWPasthRDQ
LAAsL5EV4bYmvRCuTpUm11wu12ruivirfbs488iKfdNr5nsuT+KAYoGR70I/st2f
LkHLAfug/3Y/t2pj8VYXJhd5tAsTBNBqW1EhJhC1Ec5kC83IIvjUfd3krmYbZ8L2
MJgaB9pO9dBWfEynv/fJM5wOmr1oZbMzMlyjtvdaJ9837VqKcl8nCNzcNGvLNpv+
IvDbHWI637awAV8fnG0jucLw5p8T69AnmEc6npd2GvMVWu0h0EVPP90/o4dz+zwt
dCaIDul0vuIGqDhXeEN3ZwjbU8TVQ0iNGkkicHmWJOpwwlkm6hstAnPkGxmq67cY
O/v9a25xxkHWy/t0TXW15A40pGEQn7BObZKOxm2wJYrncuCdSYTNocmStLjOng0i
JBxmN70Pr9p+NMMSOV0BN5dVPVo1ecnfy0Ns1BU/pjmgvnD6Ci7aB+Evxt5W5W2W
5+t0J+nYNp1TvduHkVyYAxNA34pKMLf7Z9LnU6oo19XGC9vMiXU0nKfKyX2HHgSR
noYnNbauCCd/iQl57azCGDHPQuR0ucGTuv55AioFhu4p/2ajmatlkvJkASqreHZt
ydAmD9u4afQx9Ju8V1jEPEqhiCeznDXdcxOlBShC8M2VNdFz31LIksBfT3mvRJn2
CMwLrGJfuNapVZfmv+zxyUoPi5t7+nhPUw1yOWVDRsGH2IXZF7J2sEUE0ESZba4E
dC7xzNpcnXuRS7SCnoMeGlaKKNJWAeT2X/yZlRfShvLpRouANzeRZkPXjyo8NrcC
8d1Zvn2HRfvxQfVB/mI2+o7LFEkxWmwSmquzaBM+kzs0kK5Bgrd+anXMrJYAuYKG
Ik9a4qQG1l8R/SdiInwA6QU/efxFjnavQiYYhhDBstK5dJ0WdP5TwJ4raweEsexD
FFEOL+7XgtnQhx3n7c/FL7kJE7i/weuBfLf3TYk6frZHtKVzaNtDrA1JmPSed43e
wC5Pn4BzfPZw/9I2nqxYSrLpirs7swRTCiEkNHGa6To9a7dzlvSZikpvfRgFHD1z
vd6Rl3ZE7fNGa2q+CYguAT/aBrIHaScFB7QreteQPMERxkXxMRkkyVNRb5+4esYA
ZYzErdiO8z2xcc+aeHBC+xfICgTE2rT79GjLN71kOQz42pn1NLN9w/r4xYpy1i9l
BN/wc5EbMC0G2rzPMJPMJJRiWWn/9ZIm0VS1uPhaGvicwxf5RBd3X9RPDS/zbe0D
+BUUyobSiIaErIv/qRFg2cdJBn2ZlmgrdHnBqlc09lzDLAl8M9SB8LRcKfh/2J8/
1H3ECig8sPT/559m2JZ3cR0eEtblzlv1e+mframO9eruQHKmXXUI7iGUJFCcfYfW
NRXwzhdGsA6MNQ3gRX2Le0mRb8jZJTAzzF4HO3tyiMUxClX9iVJSU0XhiVkIrkV5
xVNvBLU0XbQQksW24jwMQTuQaxFHi6uTz6CIVu2B5FJfNn7uEDD9jVvuL5xxosJj
5XNBSp1KbJ1nIZ2IXFtNY7EK/UIysKfAEsDDhyC4KVLxTLWl6mbj4DWCAhHo9v+0
i2kJZ2WKR39evk81Q4CDxUajaROgDkc5+moBg7HcnH8jXqKKpXXCd1UrDHuperjd
T9mgOKYtTKzSEDVapzUiGjjVECuEvCg9g6K67RiqwCwNV7o+Ehls8Fl/DYUWORRA
60z+tp5MKPJ1dOOrJKg4c+Ur7WSq3CCVqKJY7ce3929HgUXiCn/UcUT1XzB8N+Iw
iOOfynbIZWqyiWu2MTog+hYgJg3fUxQ0AdxCVpl7ZBerhvh55VBj+cYXKDriwsm3
VnMWjIUghZ99bVxd8W4LzNykbfzbDcATZAt7v+llgg6tRKgJ0H1oeegPNUnA5RZb
M59+4jQlRRTBEOweKjhLKr0eTf1bV/h30QTCCADDhbHO2HyvVaInh1EalBq//jS1
gDmEYYreF+xpm6ggqfuukpN3yzJqCjaCRtFPRdj1j7V41ac4nJSZeLVLvTk9YEW+
jDAXlM+Z0EzkYii2BILiFuj858IuHbWYwpaX6hUZDajcOFp9hnV+BhDGS+3O8GwJ
6JnbTB0+4ok5jpfMHKgB2DXh9mqsgt9mnKrUKLvETd3tSv0nCy2/se+fh4pjCfi4
9fx0S4vTzYYKZSXAtDJ+NYr6JXRfvBejR62i2R9HSmI7zsbK/G6oQBnCZygNJWkE
sZYzAHMkYwkUBQfS4MfTShGTNJQfil2WFtbMTXcDUUQvfjwAKUUOGNCtLka/7vKp
MXukFXWb14chgUjOHF51wC/NbpbO3xJOHVWF4eXDSadhcuQsYjfxAUa5jgnPMZrS
IKJAx9PO/xrl05OyQQ1K0sfB6u/6qpalp4YL6D6CaVBGoPt3Ypf2iTBg5aYtVTkT
mWlpkWfF2hPKR2W3LdptRCcoNcgKKUofoLUQg+YIyN+0blsahpUXb3O20zFemE7m
DZng04tEda9V95Yk41iddFcErAaL8Hsim4scQA5OMEEA97luiIlcL34WzooPBM7S
4PrYqzFdmCqQ5eJdD0QfoWZR3Zwhg0MSQdjR8RHm4X7R8H0Ps9ycjmRLTjy3FSW0
5HY9TprDNyKKfiPDO0hzwApF8brOTbQ7k6RMofnqdizALER2ETKOWBiybS3dfiiQ
I6/E4CSQ8E/mXZCBLvR7ufflT2Br+mMJpiTcKmCv1JXIh8HuXlqnZL/d7W6YYlNS
9KmdnpouIytJ+lLou4adNDefXD9lyQPJShUZEyB/ps5td5SM3GoGUaJ4YVyCiNtf
vCFzPvPQR5Oa2rxg4isfPcdihND3YDCv8RNlEImkoTyQ1c/iqxT1R4dSN1VoSKGF
drmvO95zVjvAD3oJbqLgn2U1ADGmiadoDrL7RNgIF1vd51QKlifGQTgNzgxRUmHf
s8MIJDLHj8p8U1LL9i5FVGhCu7SmpSw+XShe+ZKJXPVJCxIF+rMhZThUfXMF3IjP
NBnjHDXKwky59anphNa9JLxTeyFbV3jmd1dCILMTQFLdnpnw/OU9sC9tKnzF9Lsp
dpq0H3Wc2904NenSFCVikCj0k459xc/HtFtfC/o3XiKVsm2v6RRiOhUDD/15AJSD
cFk5b+8y8tZENcgpqGnPlCgztuwQDNR+w9extsSqpjPSxbQDG63Mdk3hSLcE+6hX
cZzdT+SAPSZoFo1ZaMCLzbhYGGp8s2HXFbcTuNbn+kx6CFAHUxw26UZFPEfksJba
Tb5qyEY0dSeVCNLuAbvvxfVzB96fYFT1bVsvFsiLyRKLuuct7oCpdl96PJVHx91x
XZNmqBppWDMHUUGaE10bE7gCNGIzhQHI/okbhv7wSrHQ1ZjnrqwNw/MRd0o/dI0x
Zf0LSFQmkCx28PCsTp+KLhnLkMKtwa+KEpVDUw1Q0ognpOGYq/i9Ce5fiLqyjCc8
GVVUaO+c5DGMwAJbQXVf1b1GYo2jB8x25g8F6JnVT37bA/6FZJanPVD2ntgFDDgX
XnEIXOzQu2vG3PqaIIRWSvMXRww+EiqOC0HCKNywHd0/7NfblQXfAqo5g1fbQiix
Acc7N+YkwOsrYChLuSFiR6+xNamj8v1j9IF015FiHyqN9hgy8mE5MClhSQRCxak5
27JvK1Hrt9QUwshVOGTIrJjofejDKx0vi3uSWQkYotURtMVNEG9+7qGxki71mapy
FIcJLd3Ti8gEDQ8uPGwKIbXSa6cGk9NEzDZRzhEN6scxrHIlIksAhwzfCjbqZoSf
5UQCz07zKiJb7CuiSqkI4lKbGk6T2Fxdha9sgSCem+h1X/sxxOucp0eMuQwGWIjj
IQnXvl2a1qBDxWwvGVR6tClpalI4zSLkjwup77aFvEfhjtjBQiVqmvyO/uYNlrsd
+uWTPAqLUUX5DfTz7vPybHuftaj5ABhtqRjKP19TK+RVVOwQqqX6M7l1G+7w25zr
B19TQH/5McpEaoVhv1Q156qSfAuNeIKcGJotfYmqwibA824YreMUnvlfYF8VGSme
cCqe2rPdRCeG3NsB9pmoWQReL/Hog+ltoONZFJRD5yTgI4RsR6dYatkeu2/uCKl1
jaAx7cPichggWoGgibwQBUmsx790I/JfaCtwasJeaFoi4pLUmtUpYrDEtfK3bh5u
qZQt7HkqyGxokZaO3s08DpoOtPUJvDfqEGVhISGiwLMD4De1JnDmKiKRPMYRCKTf
MnHyUhdx4nyFObRIhy5LtcqqEZf7Bcm07qFkKUgKxB+DUrapq78ifu6XYsHV34w1
jkmMR/vkAZUBTBlxiwIUTW6XoN41/DrGJfJJcce18CzLkk7i6Q1Fr/50jOs8GviC
1AAx/fOtKeBV3H8nCd5k1hN59lw6GUkWVJkw2XxchL7GWecWCxit6dBUvdBdUZgI
7y6zWxY7wVFkvk9iIvky4CUMB9lfAjMGaZYWPbc2EAg1ZGoAveLb5kYwCYwft2WR
aPIjMu/MNL3T5/Sv8AnxeuGGMo29OwHpgba9jwT6FUzKeQRFHD26J0GzmaRYo4u4
8Jx9TduT6Fo2U1NgkdjDQVUg2kgW+eq0CRaas/D1g+mSY1j2i2qzihppBEw48Nta
OozYPaKYP8R7CPNaYjDIDWjD/QLkNWcMVII0PkkpjyBtNs6kMxL85evuKqXUvIjJ
bbAEdCW8f2Q8raGMxyzZkUxtX7kljwLtRaTgKfAGD5TTOs12riNqh1JA39S3aH4D
1/CaWOz1HDTIp1PNKWjsTmbF7uRbL5+gLBRrOUVjjw/HSk9DF7a1SQyoh7J8k5Aa
KVliZR+8EKCE7G/utkMwY4EuZIoCkQVZgsDA4h+D3XMwGHiVM43ebMeOpvMfqLLk
W9qbVwVoKiNtXEMBZPmhMZIO06KA5xlURWqcFHWebLBcFOfE74FoSQd9zLQDu/KX
2NM7bO9hhMFMWAgiRIzF61O1lPjYq2st34+Vybsk0fDc2A4xsnGrnGvH1uRQ6OkZ
A2Xfa/HeGvKIp181FvfGCFppUNNS+VuRjWo3cp7k6K6Jvp+kyU8QiMb1R/I1k6NV
TaVGcNzuqg5FXkVxWuW2SsYGuzHa5V7AePdz0X0eyN+zIxWFKhIZ8MAgMVldrfqI
0/t8aZzEOAUF/nTz597IJHR0kbzaZ2MYQ58IiSlWXvK8y23coYO7sNfAUy+GGE1d
ySPSaTU6bt65ng4D8zwTiPw+HG/F/fcZamTNpcnBD7X9aEApVj+RgIdz91Rr8kLh
UxghaP6R799R0FFH5cc/DdGAg3lGtu5luGt5qqgnZAxgrNJ1eFxG4A+f712pEopi
H7KcAKPhEVueTSoz0eLnGoRqFcoC8TvF1JZ/IGDV/kffmQHftZz8wmKjqHXfAj7z
ssAi3wQsLzavNyxc/p830dtLhRMUkS4CFI+J80qRr11kuLbTWxsNn7Z6sh1EAAHy
cvs25Omga2v7Pe55/oby4bBPXDD8+jD3yhSIvdDZLvsmD9d9Q4+Dq2exGJ7teHrV
6tMHuWJCyrv4kDCElsynXJQWWW5n42rPU5CHE23+Dl7NFheXxMTTEIR0Qk0CvPdF
hdME0GGL/b9aWiLkAX6uk0yAmNj0Qv/BwvSQ+jfVUamQ01+KFRchphaGLHZCzgjq
+QjtYOyhaSmixjT0DFhvMGPZkUrosfGO2xA41nDTmpD7Ay8UvJMa7q0nGYsSb9mK
RuisXU+VC18b8d3quWWrEu7RE+NoDjJnYIrSdLdDQ3FOa0eYe+ftk2d32MCjUoGb
MPmQyzFxnH7Dmkb6OLJ5jToKo8PxR98Ux4CaTdRk7Y7TqfD2BnQcu9O54X1zOmeR
lh6Oq6e1n9V4xh12C9x+ebxfIEqQWcsZs45GM1nopZ2SFMw3KKbslyI8GpK8yd/n
y0lDtTmtMisJVM+LAp4NPxMIiQt8+w3HVo4PvkHaCTXAhOGUYptSwwFxY/WI3HNz
Fznx1O63lgV0nwUKKgHih+w+0+DFtDouI/DVsyBKDqZvNr6bqpGKQnXGl5lnbJb0
QXzlECthFHDY0XRfCPcENgZarbrExd1TXxopjIAIKVKRfJSwu76CHv5MVD+QfizP
qerQncZTJ9o0KpG2PFk6FRDzb45ot9Akl0n4l4iNvibIH/8TjDBE9v7XN/1H4M4y
o2WgxNGObKgSPK8AKhIxkDTxMHKd6GSwUxW8qy/z3KJqdlFuBF8zFvCwWfxcTDZZ
BKjIGlbNK9INmQUnYJOwnAdFyIpV582utflJg6jv0OlSbOazmyE4k5JThNSjoWdy
a9thbmdNgSKvpEReQxciZHDaO4JjcsCkFHtp9EGsExY99HoS/jzkg2gUHbjbw+Mj
1FadWhTaVutnetvbRy9MvfSZ1uMHKzEn2nEJgQM+/tYF+tOZ2ca45vuNj/PqOIP5
FUtnLP8XeKVSPmypg722UUqVFpND5WiyyYYQzCObLu6XRFK9V5VqJkDYwpnKu06p
Fn/XQQXp1wCg4eFACT4kFoexXZnOmrr2uym0JcAUXFkUWaA6Rjf4N1c2IKcHxaMO
x64vK15N+EbxYjbNtNf2wjg7aXAyUv1/W2US+Wxvq1EbD0QnHd4SHwLnKaN5eZMo
/eGcNqviw9auTYq1nehmSvAWE1x+zMTBmcQ1Uw6uq0lo01fM4ZjpD6BNPfaDM4B0
MEZJbML+Qq8hb9zTH9pOV2Mp/ZYFq8R6SNEOQpw9qrhPvzG0Tfw5NNHnOMN0J9cI
IAn67mu5l6gLmid7xUE329MRpqJC1s3TZYwI1pZ+rXxnRnsKeOBlapM6VRXsT/Kh
id2UrRf4wJHxaL34yYkIJ0YASj7EJBTRiEB3p/mmROWSqNzAEVSGA4UjeCYDZytr
hcQL5kHD1tzQ2wNpwTPkKhqdmq/eZlvHCQjZ/0PSqUo+tRDGxIoefmDuhUOSForT
n4OvDD3Y0f78fLsiJOozUr3rcsWU416H6jb7XdUZP9mHwn3XE/Okq6U3BU5IbeaS
OpTrha0vJkjqIZYBikSMaAEoNk7uSQhlHa5Oj3iD4rvRnTsxi7x4/31e+nVpTuMG
h0jYW7MVcauD7Wkuk8NMh5zWInuDsl+5276Ga02PHAi2VFsYTgeY0kpC9IWsiuNY
A9wh09U3etUcNv6kcefOmjolM9/Q+/SpO88Ca15jfhjEyStVg3aa7mx9fyQWq+FD
KnvXrkEnfIBRUvkAQgSq670kjYOnKFYE3/NpQXiNJh0u35Gh1QofsM3l53W7sH6j
4U9DjivqSocLhOn+1jFaMiGIjQ39of92UL6QczmLwMKQ2S/YDVoHxWnhQ+m+Vyjb
ybMt9m4M2IrxQUil9jFl2kmcR+ptXN9MifDyWHJPYVVyq6evUKfTisugomg2uJth
I12IRl8JszgPUMY8czxAKvV+4iEWd9SR7CYmZrs2L3w4XlLQrF0RaDuhEDey8Es9
yCroI45T0gO0cG8DP4HtIADF6SsrHcgj6nEhbQTVYmWv7BdlhDDHnmd9RhA0wk2q
ACDMVU9T3m15g3LCLHGez2TjNDsuA2LmZROj+yXC8dx93CATATqFsxrXppG56OIG
uCv8hSDZ5PTP+fD6otqhXZ6WZaJn8SAUIfULHG3/LxcQ9vN9uKfrfpz48/21YVcU
ftQXsqlkkD36/mYi3rjagIwebUEEWlylTjRxVbxhSP3V6xtnaSIaoBpN1hHYbn+1
mm7PCFNwDIhMr+VekTbfK6oRz3vAkxa1JaBrBI3EpHUp4FFAys4XB4wZJczg1gpY
sbnMlU2iuB3jl25q2BNrROB35fSbrv8wiuTewQd1HY4jwx0ygWbOL/D0/oYoBKrE
9TPKw0BN08vLj8RRjMh8iSDNvQ+VYDMTQkuVUq9Sw2Na28ApMP59L0q8YJJdMHLz
VU7kMYXs+Rvr+SfuXxsiqaSnkpkq+gQcy3LwqtrGX0H73BnA0kTGwt6u1b9qBKH4
K1ftQFX5BwQT2tsNo1UNfIOWEfQR0RT9xLzE9V7ITl1hif76Rrr38gRyil98m/O1
wTfObbaQy/7AlmuHACS8CRrYGjNQvKhLi+/WN0lnpOYBmEMTYivBNcP6QQwfJA3b
cebV8OrPbJXkBnzapZDbJqvWjNgUupiNru2SY2ESIMyMBRsaykMrb/NFPMfI9wKm
qJpdIwpg3mTSC+N7FLHrDCjy1jr61cWCUvlzLy9MLVp2lYicYrNE5TcrOk+yu3WN
FTBP9rsZCO4f1yUl4XwJDoHVN14h+L8ukBLaGrYA/fxxuET6LI/q+Pd1QoYoSnY8
/JpNEU6KKmis6SAdFKH+LiLhZQiIitIedqj7nhf6Vw2nj0nZ7k2hESCoJmxvMTf0
QbmasAPED5NCjYwV6HRdvS3WsQQZFSssah86A1VJst7PzMtFDLQ+hkOg1/8CnHSB
IPC+oOoXLsAmgf0QnRsXNcbQ5Mv/+dnq4kuPq/KxU1QpN6BU9LFJ5ErVkB5kGBmz
Q3VotNzmDIX102fDms9byjVtdDepwVL98RbnbQP+wiXV1u88qwjw126D/AJRKUnl
VeMAPwwFViMUiF4fTZzBSJeGtuX1pRU4lPmS1Nm2opJcViYPEAZPPlc4V/F4LF54
N57ZqUsma5YsYW3R6OXRhAwTy0IXw4vTSHFryQZfylfGSUpuViBEELwyoFcPCeca
uSfmPP4uhLR8BMqi6oquUNkZC/qhhjdz3HY2JJxdhfitifUXFFF2WGqoonigauBG
lcL5AeY9P3tmRGeJ2+mF9+nfzyWzXMVu5PaZrwTMdv3MhukIAHKUsORFzch6CVac
YUh9nCUdL5B5JVLWcrNHu6KrWxZnYz2muF38C8Vedg1rbi9wmWzpFbzNQVSdxLvL
mLDohh2tC579v8rlo8Hu8+hNiZz9R3VUNaLoOXGESUEJbSCH5EX4fJ/f6vpKR4Xs
2DK0wmaYGtNqDT+QSb5CJyu2hovAvB0jlui/eYLqPxFVfq0Kig5RqTLfxFsFORps
YUz0B5jA6qgfSi2r4ekyRKeAMF9UO28ln2/R5qFAy9oZ3GW/Af1A/x6FZzTjgtCT
70p38QXno+hAgB/O4B9I4DejsRDSbA/CBmmAWS95qRPQSj0pvl2wK7fUzwxy+aBm
cTvReCsOEb4p2YfkoQlPxrODHgt3tds0mKL5WkHSfXaXMHbd4YKSWScuHgQ4UGVe
s6g0ryBUlm8+XwwakyCDwvvv8GHemBt0NdxMPk6UzcLm8Q34/uzlaST4YujeeyOf
zAJheSW+Qpb5hzF+XnPBOLDYbc5pVO6QJmo898b5OOjZdORgxX986P7kBQbDjN/k
o1DfeSGxWW1A6N2q+TrBrK8rjdxoduf3+WPrvq7vf3jIUUOcf3jluY/lO0jHyFGv
TENCY19y/LiPFqOV8vLfCgdch7iAMOe5n0V4otRsjI/x9OFh+6k+TFmJ1R8OAESN
1EMWmbmiw1MBUIxfat0ROXhWHq1SmQO8RhWYcYhoE0G0YSM805fTJ9ZXdihIBK5I
nByIRL44VeMSERJC0OKSS3cmr7qdqRq2ka+oZJ63CNnKkYd1lqUWE8g/H+QWecrj
6ZiCCgplDfW7Ql4RA8u1vjbvx6kSJMipTlG7ch2MqYkTUKSfgNql6GyhO4sq7FhM
vwh8C+SuA/MNCox7D7GIXw4LBetaykRAE2jXYiEY4cZ16OMnvn3UC2nQuSP68b3i
pt9oRkidpobOP0iMq/B2pWhEKU1B6+0IK0BesP4adIHzyLU1drMRig7wG61u6ITe
nI8vC0G2iSi9irhk0RCTpvqwsy4CmfzteJUV7xA9nNVQg4kAefWf26pKmIt+lSFa
C1XM6VZI+kTPDPpsW1nwJCrZFgPwnDRMPfJ36BV1jiZszjGHFgqHN2blt3++VsIb
Pml8AyGH66doJRIq055wX4XguBvx+gDX1g/B15DmYl4nL/6v1AmThJGNsbyttNTZ
oYlvTXJrpq34ylwOW1tWsq6g5ADOQCax/QWgf5rFoP5S/oDUnzN6GSrfSd2nNJJy
TD1YlB4wwJpH06aAVMmoVgpTSoKu08S7n9iPBbJV39URrFb/uV3Z0j+PDr1cU8y7
VXrowzjUPJEg4iPGcPK+oUN/kCPiYX1l0uK+pzVaKQyHShx9b3dyI9/5N2SiCaDQ
CqHUpcJjANESkTY/GGh6p4Pu7X5F3KrtCu5Szfxv2+uXZEIanV6ziTFzcYQT7Y3P
YqD2qkSiw1PgC1iLQrNh4Aq6LlXwGhCeWd2xp6S2/8WBO7cJvWoFpjKgeRRhf8QK
GuY8VwQYQ+jqPg6Mn3m4NL7nri5KlzNqNHAF2Kkmcnb6xZxqIuY+W9vMuoxUZnbo
vjiKjZ9oYx15p2vlJOLrVrFtKlJ+5vKXuQUhvaI/BN1n5i+XxuyLVndOE6uSuzMg
GmFv8TaZYhBjx6mmivwJyBpG98Y/Z7W1gyiYhRry5kuEYBopXDMGwFGKiQWchbEe
+YF2dMQZBXfyI3aXcNHu3TnuQIUU1w+A66opJWi+RPtQ7LNQDwfKyCJXF7kUBJ4n
b8G6CP9DKNRaZxxRPFU33e/Y5/y8tyU4xfSiVJ3i3qXGNqFV8T4c/HoznlAWwvPt
TH6bXDUnq/lsjIyzALDSZzjBWlPfnQsPckyt6UP5lxf4aoo9xFueAX+6AN9IjyZx
oRj6Nbb5p1tDW9fhApOVIX2IVE50PctMmwZkcwq3FH/kBok58i7W2Erq058zK95s
W3KWozJjk47ZYGBEhCbvT0WpFzYbbGhzRTClEZzkV8kJgAcHKuBep1cmawXWwsop
wTEfoljoXAvtHB4GaHY0aDMIC7Nj3BaG/VB/KY4CAmj7QGANr9dvjX5ViPb7EiOd
gj10OidUL0S1hTJUQOcc6b/f8w3Rc8Sxil2bSvDdERrQtks0RyClujqtQ9dCrHZ4
c2qOWqjjuqMbhxnhT1muJulRopFlv0X2ICyVMsdFXZ0pjJe9Va51VortmTMMwdvT
2HYwB4PtFs4cAgjy0caWNAqaCMGz9UJ0VCAHlSv0X2pmUdbCDCdD+xmo5Zcwe1WG
GD/kHwnwwf6QP8Brk6daRnWXj8byEX7MWnHAxeYvhtEKJGOehNDeu5nXEzb49RWq
AT+9/93MaLfDMd03vEB1//F7q1/aoxLp/e6tWlyp5h5o4QCK9oobzC57+LYI82JT
pmHe5OWQN7mhtxKsv6rll4c+ulcb5ksPkN/ArpEsM94S5JQ3MrEDxNY5r3qmBl/i
rei/7AhY2I6xwN0GT4l9yfyg2XypNZGDL028KJZFKrmDdH1BDNU68q1a9P+5IxsD
WJtg7+O5+4nykbE0nGq6Y/ZdO3B4+f6OtNO2eoe8NunaAV71QVmORjfHkXIqehhq
0TnoJsC8JP9svdSVmRT7Smk4hvhg0ZAjVbkB22UzYPJv71rxu+UsBTGEMTF777nC
zqWA98FbRgiTv+G0AiacHjHVvchiKoLEvlyPJCYmJ7jm7XDs0kiEoCA8lrAOMoq0
3n44zc6eic7I0NfI/UV7eMQjdoJiAUBmnYesdwo2PwVVgacwKAJnGILQi6JoT/+z
WB/24NUVhrDL3ktNdcCFBsMuiqbBnAmgOheA7RnbzBf4ZSyxv9gk3YPzh4krszrs
WGA+aXX/jHMG78Ei5mwLCF/pj7jO0YkOM2ETFI4ET20oHMfIR7qTL5kgMYStdKF0
jHF9bJyYZXettYWtpFzLbSrjnrrrc/d13frv4xYA4SX4KQ5lcRSUZwOyntb4kVHV
euceNHTyfofH0TPP6+utctPMlrl3nNJlYMlyYlIgnEpQHqzwITnap5KQFhKYPV6K
H3R9Dp+G/GSktw3v8FxSI9PPpcSrxgF6ZaJ6Brhh+WSOQBu3qjz4RIqx0wD+lblh
RAGiyDdAZbSilybsDWVs880n4VnKbTImpMRu6Wzm0TUqnuN4Xb5DEZ85rASF2Bdl
8jCiVrRf3alSBycbI4zsvXufA8Nb3xymqeXTZRpVKYSvCUHA7xTbX8euBJUpyIs9
D3kygT+Hy9yHTEUp2i3AbzGtMWwRS3F/IfAYucZq0CpKovPi18Mwxg4jnNczbqJY
Z8kMv1JjbXfeOVEPfcNnoOZCfD89HtaBxImZK9jTQW6FDLwYEobabf6SEqYJ80le
to8cmHU9D6OJh1Fco4v4fCEzyCACi3aX5Mc/WiSF3oVyRe+c6e178GAX9VxIHNPn
Ejn6HNVKN6f5SzSWVzXNv2GiY1Zs7I6OQJscKpmqmj/998afJHwqHcKosOpIRLMf
qbzK4QnsRhCv5luNPgXLVQD/LlCV8DUHZyUn14fsN5Usa31iTcTZhcqCuLoxo0Pg
6/BnjMX8vDXsRNOr7fBeLrpvF4Kv4ovvQxiXkc+KIDWr4JDKxNEpMYOt8Q+++B/W
wvldUroNtlNAfc9YReDeA+GDSLBG19X1B8rN4ulc5IIFItV6Mo/4qetGbqUjl0Ie
GGHVaTpFHeidnts4PWUt+nAJ+fzsNNtz9R8vVX8nQXfgBALVaqV8Ja/2vaxvqVIk
mUMScK0rdcecn/aMgGXGCtarxgckZgmHD3fc6CXurwi6YKQ0TGwv5k3h6QZcmi0v
Eutz8XZVXoozRnAQwFL8H0F8SyO8Bl2Quf2GKwOS6A1fnnLzt/StO7PpeLyXNrcW
3GlS+4No51koDhRlt93NjQWyMlLUtVRIzzBRgZI6bwi9XpeYWg3HjVRzcj6NV3B6
mTHFcX0QxG9oJluf2+sWsK9sL2+orP1lrWm83566a0b962qCnBkDz3qbYtLIDDgL
jvDlF/SLTGJKhEfZM/whF3eD1iz2WDdk5Jau8l2CwGFTvrLtqTRAka+KfjXcspha
tCXMRhmnPnkmeIEnn0H51xPisJqta5VdI9JS4bDNebNo2LmygQGUtBL78JbbY0eR
OeFJpTvPFCjzkq1tiA6OFcxGsyGEAU1L1aMvhw4CwBNgYMAwKUCwPZPQmEkfZK5V
kabXl4YEuNBNY4aSUi6hFFvf+kDgczpXPs9Rk39O+/0CTpdh/ivnMP+0fvkCB08G
KDap+5DUzQqjRGL+2awFAXv4G1WOyzOTXkn3zW9SpQQ6dSnzXzl5I/S+iuxCYImy
O03s09q+wUfwanPJKg39rczBIPXokcPrzpuh2TPdMARw6unk4IDb+KrY062x7m2D
7zxqoLWuKICAHaMsI/kS20vafpFauD13dIn/PCF3SP84OZgTGrn+vxLLv0Y9JZnr
m3o7yBQihmH7m5Nl377eq1X4B6gBln+OLKntHv33IBdkx3+b88DjB43thH+sxA5h
+ncvIlCiD/LCgC8Ev146OsZmWgAEacrX3NoEK49Uy2R+JCxv1bVA87hVUH+rUj3C
GDHtAgHHXwdzOHSOmYqmevLp3z3qjI8S68q75Alh3B87XtfZ17V/FnvyuYb4I7QS
Q4Awh+fPCo0oIvzcBVSoJVrkgaFZfj2GRm2W5uVsvFPxhaWPGysesF20srbHo/Rg
oPV4eMu4LciTQGlTgsgME2Y3QAvU9vV+RhFM+JOgkVXLnru7OY9NsS22cYanfUrr
8Y1cJdcrs6TLzn/MK4ItKZRiA0lqwDuaYA/u3GX3M8cUIS35RTcPiUShR26j6tzD
y/+4VMOyJR1QGpe/b5VaRuG0BeS3FkeI0VP0m6rDemx1SY/BdbDzBAQa86jOJ8Dz
EEyGUHQnuqKJwvXSORxIVkhXAUMjmhE5cKeuw9g8zngvNazXvyIl5aGOnMAAJeVc
RTpqhIUCU9MTMSRAR6PAvTKXo6ENMdi8vso/1MrT06g1QU+J1efHHiAjplljb3TX
6XVZ0IdUG9QOhtiEhJIPnR1EqKp6mZUVnea+qscx8grP9otfhHV9BA6zihlqQhYE
eyNAf5nbWDa9qF6GROrd3dCp5/MtkVW/M1v+cw+941Ri7fpAnpX9pb9hQDCOeXZf
AaMPvqH6H3CLqy4Fr3gCDBNRfQq/Zm/xxnRr4zU0m8w7wUxe4sM8S9jfmlSoM1ad
IHPnca3hqsLvzpjXUf0D73Z8Dg863BlC5eDdTbN9HfctztdfyD2AHuKuinShqejD
INZUm2OpdzSuSQktOCQnEv782wTydnHWAIel+MAWxBoh/E73sX+VrRQwanDL5vAa
u3G2n5XyHngPps0pF4gVxESCBZWhKAgDwej8omcmHyl5NZiihwR4g4IhA4FPPB7p
5PNYRM36iwul955tTSoduO5seOb6E4RSHu0K1OppGqXBuXY5Bw7fFqGXMQoZwXKe
XDBSci87jEFlIOF8y96VMyCLOaTKzSreJGgCTbYVMy/fdECV4u4JZ/ue5LhBTKJZ
u+yCcteFwSMYdagaiL1Pgn3bEavs591agB1mMP82q4LrF09/t8LlZDLvNMj7AcWj
TRH6sJ+ycCn8Npohsthl5m8whBhRpMbZKpaxTwuXzaDZg1z1fnqregAl7OFbvZrW
Uds+tWSoupIkTJ8BP2Lhoe5clUq6y+BKZMKaa4lWLArgxAoZbpUav4QBVW5HClur
6SEA2fulCVF82e1myEvdLL4uR8fmRBnejYZuWFCIP7uuBvSEWF3GBr2hvVFQVCtU
9WD+yTMxlubReixPmbUZx876ChJhFaVtbmzva3Dx8TQWtD8OQSli5llaP9y6Y4PB
HWMDWiwFlFydmA/xpZd2beIn0XZ1fow6UQMFdguREnopCy8QmJ7+h91foOA+jb0N
SqW3jxI9E7jo0tSahQts3B71YwK/PJwhg6FtqwDrb8TCJ5p6b3hqmz5M7HFdvTvl
e733NFBMsN4qyLxHObctrJm/2ZgLDZh63/kiKIYiQEKBouDcgG0emUluHkefafV5
TcrmfKhtVfZBxT8rLgjWyYRvrVpiDiVG5yqmH4WVRnuha41wm0unv/3za0geMdBp
d4INS6CaZUtbyjWVDH5hMnQXR2ysGbPEvVeJDM+3aMo90vLR930jP90xMJ7Ffr19
Qq1e8Nl0BxqVEntw18mMvnCExww/+SwHvF0FTshkX5goc56vZH62HV/zrOEF8+bN
xlpD+d0kz6Ih2GHQ2gMztorEesVEjRUDx7s314sKzXxo4/V9W6uybUUtTwM9+GiL
V3TLYwEFZPn/TE0r0ZWJ0p0UX+nuers4Ds48V1SNhkDKutFpjVp11ycdo2Da05Nt
GJp26FWu4FbCkimnJKl3RI8J33V4hIxtNYlYdcd6ggWRylohocTvJoB4CQqvWyww
QmueO1SwHVXGCNUMrbEtFDiGZOOShewLe0334PqcRrctfk8lSdqepZEbVrv03lza
DdvZ170vvI1RvMEGK/z+f0gBO5/nSeUV7bLGcAcZZnYsfvqTsOFLkRtA2/wtTxfy
0R558BmQtL5aukvEe21ZOCKXDhg3yjthFwA/sVU6/7frlKzOOnYUzZn0GObqJtK1
7PL/h5eCo53u0rfwp1eqoKmRyl6wWwynstRZ9wbhuxnvwrRRRbTmsXeQlyynELO/
h5VJ60MulVzT+ukYmH0tbJuqpwovNzDKHsWrb6QsznbgAR+GFPziGVJ0e4zZBUJe
hK1nPfk6HYGkV4mUibn+JhpgSI4797WmS/4o7NoxBZYsz+YYdWhlsMHuVxTId8Mj
aBXzPwgfK9/T8gIpl9O3ByQe3daBu9P72Qzyh/nixvf4lmfzUkEnjJ+t0cyTomUZ
wBaxr8onLhmZgaIZZoiDNChQ6hd/9eixQo324aCmabayp1EFqWwf0p1xY0DVnW3B
AdJmh4RF20JbIgfkvGk4bU+Y573hq9qudru5rvlYhlv9Hm6ajen46WM66b93u0DZ
buIvzflEWSmClKvtJUUGwjMw3+qpGycm8VHiLQGbigaHw6YF9G3DcnKah+vZJxlz
hibC1+1CV6a2MWcIr6a2ypPKHvCNdCV8ubCmiUVd1UbckwKfmTFANCTuegv1AK8F
PLXTIWxMyIhhPLFH9Si2vH6g9+iP6XalLe0p+czummirqW3ToWM8KpSdt7RFNBHy
Od6BvdMtIUz0dlmYPDA2nzv/xRJDZzuHWBSINTHGYxoWUWpvgbCSBdhEGpRHHhat
CWWJUkRU0nXoWNksCkSr5qOrLJGXsLbD2tIYBL1Dx0k2mPgQBray5j0sasqkxgjE
hMXh5K4cUXMOdl/OQ/7T813Gz4h3hpLpd40lZs46CMOFaeqE0sx0vL+XI8rFSxjM
yHpg1pT6jNyR6y9kFj/knE4MERXuV3ziQkYS27zBFOMb11fkoQfjvLdV3bin0sXS
PTCaHBbNe7sqi7uZwM0YbbM1O1hKJYxa2FEyEymiQum55dTh2JHZPnjimsIqLWcz
cwanb9OETjiMgiQw9w2lEaJbYRRO8nEHNiheGVR3B9Lzvfqn5Yra6y8Jke4ibtMy
c51n+op11wiCal1nZVLjTZ1IHqOciYskxYRP714qaSBPyBKk+v0SZgbCZS55mvVM
wC19tiuAU8jL1T3WfoI/0CAxV6xn+8K2OpjqTN1m8CMW9lmx3WWkEIDlBFdLVBLV
ssoYKJ/cn4A+m1yQSWmcCsylXwMSAMG197Zg/Tfq1MP/bV9rKIIdzgiBNWq+pUJl
j5h6hNkOyN6NTcgNqHbyp91MFjTo3Faq03VCVPs6voaSAqrhO/K5F6CmEeYQ4hpm
WG81ibCY1Euzgdtvwz1bChynJ5xLj6L4dFUr9BmhTOVmIT7Y2vWELfcJmGP4ITvw
tGEWMdplT1QlStrtWxScR4s8VkJQuEboWycdPHQKsxOOAk0n9GAE8cC98qs/CUHp
Pp3TAmovwHq3BRHV1lLDjDu/KIJ55ducwKQvoWzb5bpK8rr1GaB1RLuPMMY6UnA3
aRGQMY4T5OG28G0q+cyqi8f0Acoki6Ml/AAxLXy3oGH8SN/gKAKbnXX56EMkaoZo
JMKS8kdkZSOWE0AkQlPcWXMLc7LrT/BxK33Lu9C/EkV/E/PnijD9JxDnxUtdmmb2
tWuyM0tnf7h9deE1DfZm7B6Ob/5K5tpzRvQj/RQmFU5vIVZpOcIAmnHH9MOmrVnk
1GwhnqhyWXpVmq4LUOllW8EkuN7N2tD0Ng2UBxHbv0GouFB6vMaEf49K57EktRmk
lviH6Iafik+BzRG4O8tjJs6wO7DIkuFtPMJ6qwUDYPx1lGlQnKgVZYRQZgWoEvhk
rLHnvpOndoJHN8h/KzpCCUQWQuS19vKjFACZ12uGbr8zkOLJDY2GF9z+XpOHa6lW
RMVfqbSAGJSzEvjhfrhiXfdZcqgVT/ttZZFZeknX9mcENe5sC0oi6a5V8vLG0U22
gqLu5wUY2IXv15AKNV4PNHTogiuahx03ZacelRw1qGg+fgZhnNm9HgpZWqfQ1UU8
YOPfYcdfcJK+stVez2VTBmq7Z8aduNuzI+euD9rzi0FLjkEcy++MBuZReVJneoeG
Gzrogj6q+bOcq4J88MWmXU8b97CkFUrUJui8eEeT8og1N28jK09vneuc+mpyNjMS
dLyJ3LYbVaG8EDXsN4sN//eBSUQskWgtPUe05k786KT3dOV6pGIPqPHFnKEwPFEF
Q3BfONWgx0jbNugINCqD8W7Kd31rYrHqoV+NEzk8q7NhP7dnE5OGN1WEaLeENDF7
C1tPc2hB/PxE0B18uCPACPlV9FS3I2oXm9gCfnXp5hjIrtJNR9v7aGO4Sbm0YAzx
PVcoI148q8AuhhILf6PbUpY+rNYxB5N/N521WvpJx4WuztoSCaM95nBtt7jAQU4T
XqNdIjzuC4QzLdFRObXqvnyuQYlozYxgInsqSVmdQqvPYIKD7HHrpfyM75/gjqD+
KjEGcVKRYrf2KPDdkjYdSKqz1pqR0TqJu7KimoKpVHk/tEALxjUY7Zjg+Ln/0nJX
m5nl2JaMS0i/pV1OD5uBKfU45MkVFlSGFyxZh98sIyVtPW/rNaJR5IOup7zGJ81o
B4SDKjUT0aBtB6bkPP67R1o+0UImLzBmgHHxR6nZcUo+8GYlWqDLbAcmEH+LrzOM
FWVFy28NwVwZ0QcqjWmOy8ddWSx7cT7HMRxsOrEgq7qBgFgFnKxeh9GgMExNVtdf
i+bTx2kJowedIh8FnuSf3u1ID3pIPFEjUWah3Znocg0xfR1oCj6/OL+pDCf2OCt6
dPL23mb95xgb39mtHOPlSdGL+W1KjpQdeCLMa3Tsec++WA6BBWkxGnB8H6QegBsd
77Xj79LGj9UwcD1vuDXcdSLt+6UFQLBs2b9BgK+gSyDyTJvNKyUScoQrfP1R+j10
rUhZcHCCJ1Ni+Bae2dTHQG1VZBf7kaOnZ5bbsKkh5cId9JTnarNsR9/2irsBLphF
oLLWmix9Px94LrBWRQIqjwegcxgio5SbpfZbnxYEglbB7wtlZ38PgQ/ayA0mPsoS
EB/Wu6wD5iQGOlcvtn/hTxuajFCmL3rmIyOMFefFy43OR7GQ90T1E1b8hRdFfhkN
eupt+q5ehcWVqXwXm2fFJDAUOVBSzludMONrX1Fsplw9BhyuU70GLwDWP1O7DXmo
34oPofMpPu+BM0xnywiqSnAYC1GbM7eqIGGyMt2mdtLtuYMIUiCEkeFPyliO1XUt
TtxX9HVDNKKDhSX+boICUmo3FuIdxP/sKZFf7gZ0t4++oftAbA5E0yOxnE19mMMD
bjOeZn8r4kEVcWiJ9Rj3JPd2wg7UWB1zqbDLCxnWEwvcEhcoEDH3rq8HoZFDn1It
B9Ae6mzuJtOldW6hmtcVjt3jNoi2IsXV/GnH7hRZ6FZKrq2medIsUoXO4ceOImEl
fbQ2+Sqgf4+wIbQa+P9OQ1vLrIjCFwo/DbvIuVxpfAXK0pEMu569AlORjsRuoKTB
kYSt1bW5yAkIeOoOeKRszMm3vmV5Is2AZkij2t2irQWFlWr88D0SPwux/AWef07Q
B0rdQ1ceFUU4qzaKF+M8QxD6qyitd8muPQ25d5Px623QDQKo1OvY2J45zZ2vvglf
LM909qNSE6Xwblk4d6reN9F9lM4e/aUlFyS2eujDuDYrPjksjUqCpDf6B3y0om73
rAmUSq5Cq7S5qqRAgWAOxSygbHC7sLffUfDFIkmcfd4JtiqVm5Pp0gexTdTPY8vJ
vaisHTfL0cm7jJ27uIWTxWGmFIuXzpoVVl2zdsW6DMm3hCdfZybDFO3ilAz5DLGZ
CiO/zNF5C5nX6Md0L9ZOWxlv5Sp0KEdmRQMrk8U5Vl7Y1CWWKkEzwturA4zfdady
yMEtwTar/Tsi9BXjsuFYg2PTjPCAl7U12bT9glDcrD8Hx0QN+whRJOVPqhSrOmsi
9GL+GXCxTXoQ0enNlDnE4MadVbArX0kUXLLWJrhxrWWaMhyQK7vWJ6kAf6VZf1CJ
Ao8MXw0yR8Xldo1aqBcJ8Xk8MzK4ZasfroziyR9jRC5M3mHPDel34rQNM1AAysnQ
30fgkFaLNMYUEzpI2pSOK1bQcg/HJ6CN5SF6Dx4s25hvMkZASQV4JW4HbJVjOona
26BXYVb1A/Tzpa80WZVwOCT/qS3CQ5cWK8cRrX+UPkYEZ/IxuvBcePcq1i4u97Bx
nu3iIy/EE37mlJEEVPMsx3rj5RUdCW+vP6Mde6w5Nb0Bri4nTA770Rwf4zMF3dXd
pkLN1JNqG54gaFm9wAP7Yyt0MYcPaOz4SDHqzB6CcdxpFd8fMOqXI8ICDo8Bu2yu
F4K72nIMnayVDXpiOOzlyeO8hkKXmL1AiLLQfiGLk1eZCDbJTNg1UCr36TIaR2kj
csBzNVEn+feoQ2px3c0A6O6+YukkIchqyUFlEdJBDg8KgX9i2xPXYknXJCQhFtJR
JC01SjH9oJ9aUiTwUr5DpIsTw/kK+E+kfrpQZ1/WtGJWdNZsucWAvZWQCz9c8zA8
jxwmNhJk7Ub7NzorgTl7oVXb8mTqlg/G3a4m57HsITdftyshqAOWo8m89IBqa28v
Ui4VaEwShQc7U+94GoX94CnImzHyoUUhlxBQcAjj+1Msil3OvFvjirjTZiB24ZPz
Urvi+qp1g+QK2OZdPPFJbhtsgug3+41fHiqfPKNLaTK5a0H5VdD0o0ja8p+gnNC4
z+LbdcSQjtqLPJVCHeQ7kaKzbAQg4Vi51ISjkVFC92c7wpdeHWRBdeTK3dP8ZquU
SrrCBmDHUJCAqV39DKRrq33ubrqGgAg2xijyvkurIbZMtTP5FRD06QIoWsHWuNeG
7p1RTCDdv1mo7+dm+q8k/X85hhmXFD6bKhfZoN17gr7g+YC1Sf0zDMjVV+WgCKN1
yrm+wv7MfjKipj+odCwLh7YvKG1DwmmvZ2EpYBzzREJLxMd5S8Bh7zbaz4q9+9fw
uqq4orPeFC/CH90A1Yw9Bu2tjkuJ2QIaFED0/GVq6k/SFphD4K0XjcLLDo0OAXuT
JJhQTzA82OGp5c9BGcFbbI4JxBSW/fDLKPSmC2jbKGLItoz9X7QhpzjyAMMmaagW
6nea8XBEC7GflrRxHsWVvX2iA6wCt/V1qXDNh9Tp+IEcYdWAqDb0h2//jL8PTPab
avCLWZHRjQNNrTxvm/GPtj1gtkQfLm/9Mj7797m2W3OkkFUTZATBV4o5mdWFFxwh
NkD8F5VXtmTz0NUduR3TLC5mlDtSrV2SAlJGU1aVGNfvhPZsbpB4+GmBs4KM7fRV
9MMg6qkRGT2hXaMtWwW1ZZpvcW+3nfkeP1oRJVgDnBZdxSqzf7Eqgwj+XiBwXuxi
sHstuHuyEDZaU9Jf7uC2B/okJvRvf4P47N76IY5Y7RgMC6l250qo584qv4ZKKj6S
y0WoEk0TIE6hYrQkGulRaRqLObBf3vj+p2EiSol26Xtdhh3UDeWASEEFbIvmXhbt
XaX5wwqx6Mt5PoFuBP1g8XHp+nSPri+B2Po1ykeGssb24hgws6mz/6oEVQpqdtY3
V/BYdJyN32LR2wBcF10c/3DpMGxdvZ+GxGsMUpGriO7pDXvfoQdJfYMWpXz8Q5Ac
4p/vJi3fK3WHgwuwRFslT6sXkfdChIkXyUVCsAs4NmWB+LpEoF6K6fXMpQThk5PD
0c+IYYoQ9YZDQw3GwWdq9slRG7fuaV6EbL/ouzSUsPQbz6pNAc5zTB+jKMSwj/oD
Vghz3gOvZQpeyPpt9+/5Gxe6eQ0LA7WVHcUJl5yPeOaqNPbkVFlndzzt94/gtV72
QNwDGHnTi0EZ/djnpj+osLOYGYawzNIGfKJgz0SjyTXt2ai8W7nBiOETsOfVo7Mk
H6rXJolDIy/kY9pI59dDBRjwqSkkdly6kDytZwM9hgCiXZApDIshiDZ/9rhL9M9e
Tv417ePLhNFmF0sj6D74qPBSMIvMAngkQd8DZQqJE7xUZApZaNNaySuOTSQCO7HH
AojyY2rVym1zDH9kZu4wpvZPvJmR2zdlOGUnK5pv8E3HSTJj9dOCtSdrj0qZZ9U6
5sbxBVV9YgzBTWWJWOyb9kuyhN51QogPUTLPkN95ci+1Nuk0uE5bA8PqFFq0eBpf
BrW3/62IH/22SztBDaiSp0G57YprFbDS3XBHNSFXFWT0v6IMgdETdd0S84RkGDo8
VdKNrWLaUKL0YNoAPyfx/PWZfeR7TQ2Jud+A7ZwKn09efjJSUFaIXsVt+3vzs4Hw
5AnS3I1thW1HoL7uXxt+MNZMcuqUGT9THri3W4Mmm4DmXTlvmcy9Eo39p5QgzLQr
oNvOLpl/7mM4JRRdt5rHp6sVp1gSvj6xz8G2ZKMkpnbjlIxrR2AvkcOb6jbcEEfQ
LGjePS8TLaOwaBUoux1dmgYlkaaaHmhzEiagX7eNBwHyXMBXGyyxSG3J/9bDoFNG
EgAMVgghC7MBDohaXGMNMzU0Ut/YVlJjUMPlKOOj4qV0M6saEIj6kZKXfYNXBuj/
NF9ENFzVFRss1dezfNIIMhqRp961jxcpezdBG9KU9tbjgjBwLHWaBpYyREBrVhuT
F5p1gonoyYTqxNenm9sqiyiplK0PRkOI/+gxfn56aE2y6UhKTAxkqF3FGaPTbrMl
IyrNv8uM86mdY8QoGkLdsey04yFXeS06w+M8EbF17kXquA5OX+pXkXFNcZQ6ZFkc
Eu4/XHcgALjesjFZ4rTzOcTVXtM2f4WpvFbckiguDFQ9DKehDU6vDCdo+QOPWPdd
6rc5EBL/+9Y6UbZo9bu8KcXAtM7HIJRNkuVt85mAvuKVy4YWY4AJt4/e5u4ElxrJ
Vy5uKy0yM2RoMyVMNR+PQSj/A+vnGR20s+Zp5MojfdkS9UwB7UniReKCH4t9B9qb
040mrFEINl/JNWpPzQOlMFkgetPmznQKu7sc+lzirPkHviY3ORRDDqZvVinWxQlS
6luWaF3Q6azuMyr/M2U7H8jhZYk0Khi0WLY46ptXJ+NgHQ6biBux4H4eW/k73+47
pjJjp75qJOkDpL/LZYNcOd6bcmt1u1muQFG3HHHUutpB7/9CabBcdxdT+G3sloia
Pre/+67OqksN1DzdnnIB3VoFKj+JdIZN0pGGPy+eXgiG7GWgv6Lk6VT3SsmbQdas
FlLPDufXhukiawFb/wNEc4eD714JN9YaB1BqeH732u9PN4UkrLAi+/DavhVXBxAD
XvjNieLcAiuam7O2pxY7q1nxNV+vwvdc+MdEoeLO3WNtmlPISeOiaqRGhy69rO8u
yjwyDuC4G0U7UEq7phmEv8TTW73q8BBTsGem6n+HyU4FFd/0Ogiz/7yx5z/zStG9
KgP70Y+u0pYZr0Wl68+P98SN+WRKusfCe7D4hPtcga5D008QLpEa/iuoT09EQw+Q
J5Hdtrg8ZLU6CGlOiA0gQ4KT20GisOiRJRrZL+IjCbfqkjMBFSWRBUp5YosImsB5
lJ5sIQcRLp0F+XQbMG9yPQbPz7oG4tj9RawTk8DvIVHkuKT0S6KcGJiKtb/64SZs
cPwzEaBaQZxGM1isgxP9VmMkW2vA7eR8eGY1obou93O274NeYZ0322+N6OWuBZEl
9o8y4B8pdRRywhUFA2hWrl2hVWTRuI6+g7JGtF2qsukKFAD4Onxe6wlmqFfiHi0i
ijR8aIgyFDbzQswsc/d5ufCQVtGMFxvbEUv6y4qGaB2yWSngdsng611nPy6NEJBo
Rhn1AcguWdKyyjWM+0QBBkDonM40+GifZNMD9Tb75WLvEBfXZCBY5F2WAq2zcbI0
o3+Ni9RvHzYXNRU8WJcAEJ8AjszD+OyUgsYJU1axOktNRgmg9FUx0syLxQloXayi
AEhKsa4gQkw5CRuaCr5scQ6Rowgk2xiNG+dP1nQrRbI2MFXrFdNPIZONwfxg9KvD
zw6gQuJujGFNBFqj0RZn/z8eiyiVn61J2DHGcOISGKPGH/YNu+mIKFWmHJdH2i68
95h01jKLEx6k2KX+R4AgjFD8GTqdwok+OzaDS14LYFC6KrSqoWexmbH5JQPuRn3n
VeMY/+YcWUDoWx0RWE+UwXAf9k16SyTJxFwZSFIPfNgGTwMiVRFjspUdSFQPfUZw
fhGjKS8D15GdSsbFIUlJ0UO5/rs5eLUGdQFrtYtqzov2b8cc+Q/4DsY8dkfh+uu3
exrT2nzUOir21YIPGUynmxOCMi8Ou00rqCB57JTwmiZ9HHiA0iMFXDZQyGLMaeGl
p63C5SB5ZY2wYzlVi4/D7v0KB1sv/suiqYpOkADcSs3VALxlrH1r1iI4Y89q3MMg
WftWk5EF4S5XU4nXtZVGCrrR4FEV7GpgtzPMm1SOOSRXj6DWShP5Zg3HEpV00TZS
ATEzh962Zh/PlwiqrK+cL5RLy+GEnxzgaT30tFE5NqKiFcon9Gfjc6QRRz0ytqyq
pU0LWibOdBOcg6L1VFAnYixYLuMx0YfB6TwR/7t8Nq4fErYKW7qp+D3GcmEzNBx7
eUFPZ2ped74KYenrSqHY9aMFb0Hdq6JhyL/8AbEEYWdU3+hwSvrtzdW0QaeJ/CHW
nQA9ONu3Kwj0J9W8/I7f6LnMLjP77cNcsCh+tnXGahqU+kbchE0y2E5MaAJ2ba41
S+jOTcqxppo6+y3R9rGuiIXVBAHGOdOFnxHFfaiwnwv7rmcHe2bA+MPY2sJvEfQ7
eGaJYr1QnmtaLQJY1kHgYtiqrjXBfQlMTMhgPFG4SzhKxf42jHXvut8jrn5Iisve
NFdqkUeeXFpRGiaGSSzBO9dnGih8iBDl57qZJSnKjKyAoZnDW14osHp2Y48g0EZF
M2VucIoipHazFXbqwwu5SVOcs4qg3GnTHNhF+vtf45pqjJCvjZ+ItNNZ/ZyuKzK1
8QqihczGGshxYYzzU0sR1pmPFa+jZl5MhkFi/Bmjivm7WmM7jZSXjGcloApUX3oz
1qYDAXj8gvdOEFuKXbvXfogICOYT6dj8O7mLXK9VRYqyz21JeaAl6OrPZpLeT/Ab
tfhhBi5a9MqVzDDE1ssmi6PO87VUaqy2/l1eNiQFUFO4XPD7n2potEVqpAEznYeR
h4oxb9HtBdimEPLEzLfQjqAFkrL+Hj08BUK1WoWnlcRlV6eU5htOY0H4lghh2idg
u9nIaoyczIFUuFw05AIFlhjV8LfUGEyrNIBPfL1Heuz02S4b9cfgIKKZ9YvV/GLi
6sWZpiP7h0I41bY3WzFfD7VMc8Cm82LI/0mxuTbOiqQVN7yjnpxq2tHyvr6JDfPv
cw4avHEzUhhvb08h+Da3+7I3fcxCkJfuGiM9dvo+pkFC+5RwLfDB8LojU/W/0lwY
8FX4+apKqbH00IzcFpesV07/CmxuMERzH7WuvvWKdF9rBSMjF5hxHEbuSFgbNKl9
mbbyeumWZ+ujTqVKmW92Z74jSFxWAHZx3UJGcKfzCpiZV+QmJB0x2YX6qPIOLEPa
RjF1RlBBI4HQ51Uw3/KFX+EkUeDkDn4kJfIrR98SrFKnVaLJ5rWMBUklJDJqwXMQ
luXH3A/shWmYffuOoOyWR7lJ6+EoZ7+LTNntn85rbec6s0jCLC9EqMXLgXY744iJ
/SS9sssJjZmYaUXC9Wbp27bhuOcShg/F4+attoyPiml29hHhQ73WbeaRSMlcb+jq
j1zvApiIBRR/Fvv1pqoXmNZfMTdjpxaeDryDl8DZ34wv5dl6ipWzG2IG/fpxzS+Y
tMmCb28sl28KNJyioS4QCvL0DutzYsA7yw1uiyQ4bdFLOtJjxwNfzWrhV+avMjFw
rqwaSlJpCw3XGe7cqxAJogfRCgX2SVK9BoafiLdkNExyjJ4tLnBpamSVHRGK76lk
/yvNpx7LDFbr+BpMHkUU0LV/eYpyuNupCSxbxtI/vcY8wXJq6wxmDY4B3+u0FooE
khL+r4QL75pelGOSKw63I9EdqEQkNOe6vbp/aoIynxp2sZ9NZVxSnrW72jnh9Ncu
QM581QrJqdvCKUsH9nxtgDWrX8RppzY/Pf9lNsPm5AtaYTuZrK9XYohp9QDLJVLy
HlIgni8tgDdr/noEBNJGrkS3Z6CveVdxsa1mEaG8EireXN/ZK83h4/mqUaNiRqgr
MxBot/h5r5sLJMLQ+n62mA2arClp6KK6OkpDl+i8+2TI0X7ydLTbhm35GmfAZqUj
iBMqb9WdRZLoO/dT5MQv9rZHGFdGbSGngwzPjsmgTyyqhIKyEs2lNBhiU2TZy/BF
2tLzrbQficGbxK9PIrEjgNVTx9kDvbrgDLlyxeuowlMskj6CcGN5SHcOlOLuvZeS
XrkLPnIKf8Tbhb1IX+bsFf69dpBO3P4xxCGnu4cfl4gTMAPLq/Tlstdty7vQ6uFD
eebtXnbnaXi9k/Xyd50nuuV/g+oLTnForwsvPpL5+W7dGXjJEnsjYAw//vq6ZStN
XzSRuzMNw4tB8jMReUiiQKut1AXeO+bNNnhffqUuOd3Dpm1UYKyltjN1ktM1/T+7
WFEF1uj1pYGTz/UTa0Piw+lMOjqFlRgDd50fnr8giW39vsaULIAoZODgLa0bagYV
DkfIs0gTzSlbow9M56759pzLrRHOs+FRT6QfAM4ajKsqKWoy2crVR5CknKqFjshn
9/YEiMWXAWzWnIL0fxOGGskUfBEgadRt+PN08Z5k5hIgEWYm/MFiWxhfBTstYjN2
4i8akAjRciky97ZwgLxrZJnUBWDKiBOFZNnuwjN7M0gsWZLd7EPFWVl2izp7UaHk
Z7I++PTX+ha4tGnt/6GpJhA4vXRPpSb+CA2A8IjavXd9H+ISCPxELqVS/OQMNyIv
gI9lLBleFioocyZD2PGkWUZ7Hxtx8m5ZXSB8tgInkJQJjTpuVxN7gVmjjFV9o09n
g9x99izOA8YnV77kgevZ17HIxlokagTdwkDBaU+gZtz4b3AgUlfCGPQYFaHpn1M3
1fuft1hJbXh3lSTbu/bQaBjgcypBnKbjBb8I21C28j45w+OsvuXEENViblk9PnIn
gd3EvcfqQY1yvKsrzcrvjaVy2VsEeH9u8DQ7u4nfwzh5pIA5lCF3bGzh3z40Lhyg
RvEkTy7Q0uPhruj2QLj4aQLG5MM4tOVAG2TMy7Vyy90AIhXmD0Rc5SgztlHjKCNG
1k3B+Y00iBqdKtSLOVRr0uMV7NkbMs/5sxPe0Ywbupbu+HGKsMw2zoEvpwPf1tO0
vexr4mHZykBRw2FpvblpXRVteYcLpm35vG7Di0M+OjGf5Zk6a3g6rf2qKFyA1Tds
8C2FdMuB5TkehTbCFnmeKuSmQgbmMKphWsJ7XORWB2PoxuIyBtpVKwGe97sKKe/d
NBXet9rD5enof0gMkgLLYfQ8toXbiAW7NtSXBnAvSMTVpEnVrO4Gse4Dq06LwQ8a
5bIaZfJ1IINx1PRMNDyVQ57ZYLFbj0l7WudKG+M6Z/i6DF4KMZ+vc2V3zOIHiDaN
kM3KOQiUWBBmLiruyOfvLNnjvZRutLHWTcPgd5BIsH8+t2z087CEg9bKptcX2PqY
c3qVUSEh649oTYBIAWJtodwzyW/M2WLf6d62aEuvPI8ZtdrNKNeDZiN2VQZGGF0Y
BSssm3J8iqSulOgW1AKdXqnQmPvqfF1iymT73vjvewsp/ri//mfW4I4ltaC26FC9
l/g98jnf1fMzhwHhpBEVTbbpj+I7X65iPj+yR0FEuXW8mTIgUNZExISETA8eKViK
QvEAsedVKAjK+pFqakSy6LHS7jEZ6VMGHNnk5tnjeLIyNgvZbg8YvH0/Od7ixsG1
gbgw/h0PyUFeBG+uQrA3QQ+yxbnssmbkMV5PqxXsAh5hyjv8IfO+2oMJIsVOJy4v
l1BwHZBDZO5f3l78S6/yxOrbaHFRjaKQEI92Nf3UwI6OwpLhbFBsFce9AE1dAi12
unClY77MtW8oyqJvy/qrMBaPbsl+1rSKl5FwpQ3PpqEBInoBeHCgN7P4TGCpcBzh
2JgpptbZVE+QvmJLoffA3tMhFdlfo6I0rHdrNJA/eCMxtaeRn5S9NLkudBMNYk5K
1vBJQjk5Q7fDh8EpDIMOmSLrmPXLVhobVEqSsQeQzyGqlM9PgC+8R0zfKqm4GdJc
dD/pDykKqcdnznpFrju6nophTnZLU/parCs1oV4prx0KdiZ5VJxMGeEmW1PYEk1F
vv5MWHnq8wRpvaxJhkPV32r2bTouPXxDm1gBpiCuy8NIio8FKz72SBF37WQL4tGk
oDrZjFKeFyrevodQQjpxBOrTYbsVtGAl/t+XYmtosvkxlj+JxbG5EesgJd6pP/uI
vdmZkK1OInu7ORuxoH73WKnI4eDIZfXsca3ffScLfWdPtzp+56kpEMHB6BDZNYOo
RXY3N0C2K2lKwKOKMDSK5u2P+FCsKxP3yV8gMNN7uoORLtCKC1aSBzHRPob6geDL
cW9T5ZxGfS+DWMUCuE7zbPROY9X+QsHDtM87+CBdTWRgshHas+LaBVkPTu+UCWxk
M39fNAXz8EKEq7XewEj7XiTcunhkeZ8zi2S5hOuVR94HR0WZLuwKbF0RWIjMUq9e
foYZVtPiRYXI9FyrTixUMMYUX0Rem/gXU1xKRmlowuekgyIXaQ6TYBW7WLflkffN
4nRZgbBzMrKLNWH5ZSbNMPAq3k7YSJNVM/hLG8Io+OSzdd6upPzE7Y/WB2kArFyC
vdmNBdAj+JfNdTD8vWDrqDW1LG/nntBo3px1vNQqR4S7goBALnT7IcaxlJxcWrkQ
ZmJC4ekpQ9EU0MKnV+4M/lSGddHsRuVRjOdgGqTnX0qyi7Hc3oyFU0jS3QAkBS/m
noFFsLo73jIwNXIYNIX1fMqCBrB3c2uhRsTWQfEmA5A5m6Z0YBED7ZYfINg9WHLN
n5dRZJ/VzI+t5CXnV2yXAOF4KZGO0dycqdl1MylfgCL7n+kbkPDuEcBmZmPMxmZw
r+T4tvJ3x9HnqpjgNS8YNO2WdWzFuSF3M/LtCsfstxcvNrbVhaCOnlcjtsWjN+E1
uRhuTwWZGQHBoL5VSjFMvYQ5MayMnN70++1h6AVM+OHumTwslJgxbTdxIImVK9jA
4DvjS8F8bap3rB1DZQ44IoMX603Vo9qmFUfNzUafgUkCoLR8ll0/ULbqiq4ROjh0
pU6fY2yfrLLx2xTaFJUyQ2ibCM0UoYVh/rT3o19ntMPGVF+Mszde/VaZFeDmFARh
a/Z0LQf5GxHeZr2+578x/GyE6+AxizZotiv+P2ggaxgT6lW9kxH5HoheRaRfLW6L
IxhQnqAKfWc7rExh9NgK2k/eJugZSbnoa5bbHIS8ABHCD0eZbxBp8HaUvzGwEWf3
BEb5CoyL2HkyEKV2PfAWCoKD5jHzPrJl56NdGXPLgkuJZAGk8L/WMTD7L5QhcyLw
xdSJfJ6mMD/jusC7zn7DWe48g/SZejzJIxuEDWSPuSaLJdLlnzeAIR1lH+qreypf
zLLgGgQkOSaxnDvGTNS1EMRFk5CdvJAgAYppQfbu6X3pbVNxsFeENJ0xlEEIRuot
iknxwSm2tgFDkT2bC9r9lKR05TSzLPea/RMJfr17aBFV1mIqQEx0HiZVIYMLlq0T
NB0a6IOOggfhC1juT1I/sPpnIDAaKvdB11rzHsYCrwgq7VXsbviIpBZ13LtfRFXo
JMxhTG9zcxtVYpiyPImnCnAK7Xtv6tisNg6vacCu8a/wacZ2TgdDCTxwf4dyKxUN
3abxQ+KDWGQ5mGziMWJ7aiWM4icL0b1rtd/8U4+8P6JwkUBdztPsxoUHJIB79W95
1TYCEJxjbB5BxPC/TjmRo5Io3udTrbeC4/mpEsISPumhhPXDeTmpUIvX04WLsTZM
fcC9menYUOKgaCofDEHHT1UyksEUg9LEsGtcrIMTADg9mTER1mAA0GTm3+bpX7iL
kWI5Pg+PX6ydOchkLvpnmIiM2SE3LGZSfGRI1dlCKXVbislarX1VQ1JtGzR0MG8N
WFQYhh/6ZTg0OxSZj7JLCMclohkizAIdviR51OQtgZOzKbGASRyrXXA354y5FKII
VH4/p1sInFaaNOr4gJ0mrESuZwAzLeFmwo2258omGJ0zYi8S4OkZdyEicZKyMwuS
xaGzrH0yiP0YIOX3IflTgQsnCgNMNxcouxrh9eeHibfH7r10fDGPlOAO0QAwyUrM
xI1n2CAhdYGR+1Ta/sNrskFsN9CeuPKCbKQeMGcXWJ+PVR4sFNmPb/2aJJnIxM3R
ua2/wjkh0jHg6XrzODwxdNeBUPuhII5DdIT+wlTvE5+sO2eaMPf9n+p3luilxdZ6
7SMZZwo6HBaOcLm1AnXFY9b8UDjzNr999aFVh5gLU/cciUzNQCp/5//GXjFnevFh
82VbzTuQgVrtQrCKXZqm3SBATp8nJ1uxSasN1hTANZDpT4ZTqQXdyKKUXBXNXZgp
PHeRu3qPe84gDufLqYFESXJQxsmjPLBqAPGIfaKiNsiCFqo4dJFIHCX4qI2o8YQb
SGNrP05Z2J5ax/rMTchyBcHyGTKuFYaVXZRCqvoItZjaDFxJWm5YlTm2xRyaCsk3
bbebrcbNcVGMGS2hw/0QCNku//7sKYokk/9tDmvlv2U4+IB2Vte7i5+7Lo/ko60x
IfEzfJ05vaMABxB0G2MuscNj1Y7kpIld49YDO8Gmz1VflVQhBr2q3o3418NKPyyQ
oaez9ynoaO524JOLtVxOeODT3AJcQERF8IKq+eca9HUnGtw5Kmmz87j2ajFRhMst
aBjnpHz/ZkAv67ojzf3zHV4nc6Pj56yh2wWfTnR735AoS0M7FcgxGu7Sq691tcz9
OBvWMjgw9BWMFIQk/p6fwoCNodbYIv/tOOJG14q+KQLHMx8oYeasIU4Sf1U4NFxD
ixbYfHOmezQ7dd3wHYTac5d2LVLrJA19UVZsn4GOpvDJjA+TdtGEE1vknr2ELzwQ
4L86vII7FN6V57VLLIKuHBV2PxySQlhgGdP9ml3w3jQUIlPh5vtljZsOyQic1OG5
AlkKaRqTHgEAdnYuUGY47/ltUQwafMjHkxxVOE2bc4t7EGu9lWBm9aqNtJvCRtyM
hUvvkmyF1/1k2mZNBUj3TGB92GHg18ku36cCKIrWeF4poceWJU5ZagrwaVdr/YPd
ihPgoct629M0Ro/2UWdx1WYbRc1tYJ1T2bEtC2ep+MhZqrsX5BGJ69GJHuXlhdMt
UKDYSDkTIelJoAKOVQg29jUeUIRXfe3TSBkaq5KYVlg/FMhj1jtDxKE3ARkkcCh8
mhbyE1bqf6vMSkLwXhmMmka1gJouxtsHsDrTrSqyXQ9ScZ9IAEvZOolQ/rU7pkNU
GWmh3DPb7HzgTDofHLXqeZCVZZCV+ZA+W36NklbZgGVzffyDQGQd2MX52GyC3uLj
cR/hhrbYTEuzYeA4fCYXrPHLVv6ab1Ka4RdrIXeemjqplGjfjqudB3XvY4Hwr2vA
5Dx2og1Wz/+2q4YRkizs/4akqtl+i8sgFynKZ25zepEmHH93oVnySA53stclmbFI
dWTW9pZuK/10PfH53oXtwduIm71m52EU/jTcxjR7HtdSmQIfEOTb2JHjX+JRfynI
Cz0qMbU7QGC444s6HKZVXIhSqKiKrziVEm2bZgAn0yYi5eaygKAq+djFuP70g6Yk
lCRzBv0PDlVzbHrelA1NoheTeWT51jnR1icULMaBMG0mbJNChnssM4Hshy71LJgq
iYwX8fgCCMOF/pFHurJOSJnB870SR27SidwaGHAEsIkX5MuYBoUM8uyMt3xNNUbJ
W3nN/5nOvV51VS04O4jUV9ghp8f9CZeOhxOHbAaF9WJ6llXSWf47EPv1EAkEBbdJ
V/buk900F3/Rs/tox0T29gyXU3+pDfLYWgpiT8xAAYb4IBR0lzlzOASBP1z6vjBH
mtOUIDw/12iFhW20HbsapwQbnB51KAfadxbFXmQyf4BrziOny4Q7VsA8dZqfi7Vs
p36LkgM+IMHtqqp1KZHE31hnBTtJxVbAD8RcuXDt57l10ZxP/toFOf6RMYBemKwH
l2g+t/kSqz91jzAbLYIuiDANWp08WtmiE4bUuvoIkxrnGvYw50y3y/GdL3FbFS9l
1D2vF2gVUpKQW+4z/15IntgWXYGzwNjsvVhs4d8T0wJDK1a9FIJD/QVHgvHkHdCE
8W5Gc8gy1ufixyPzblk5RHSN7zov02unurJ+bGnFCksxCOG8hJ+yRybEvDvAfz0K
F5metxHNtGUN6qiUqQLVa2TVZjrgY5Wek2bfpWFwHGz6E487K7EabzgFtTVwMYrL
vAhw68V4Yr1aKi+xWDyqyrs+lQwPFQ/oHXR62xystWQuQ0uOwoCqEB5UrdqFh91P
QLqx0pNwVTzy568fqDdzkXcsojIiSDrggM2piYjDle+3tI3NS0pdlpV1LFRv11sx
c+mat3CLu0Tv57Uqk/2b/5GH+sbMbJ3mHmEyTA6GIvN8v1krleFLheOrMyV+fguZ
XhQy/2OO7HGxJl8i3gpWj0JTh/mPXMD5fxLcYTj9Q063mc2YPQ2xo5BhORl+/nvJ
T/3p2XKNw9a4ubRk88sWP/QQwAUXij5ncd5SxH3eN8xlz+I3OlpOkNUBgFrbE9bc
7LBOzUfMFNdVQTuh6CyNzpNJHKW7TJ4kdy6ZfDoP6lRpFqQWRjXsWgI8tv+PVQ8C
XSr8CsrZtfTYQ1QhEGza3JL29ZQxZ4SCNcmpoaaOAgFRo8G7XdJuRTgbHXhyhfok
8c/S55jJSQ731nryOqSSaEmLnjoS73g1czmIbGmfbw3A3PRDOuegvqXBTvh4tsD3
hNLA/Wjz0+VPQzgUF0ewZTZfpm004CTZsQj1db1qaFGCDYNam1zm7eYBNYUEzd+t
IRqrEqOYLR2e2pzVj9Lt7m6T9LzxTSIsa+0BIhpTNdKGUZSenkIeaFj5ZfnRmx1P
C+nLB2wXZ1rbSlGbsf517iRlacKENRQHu9jcEJ3f0Qf8TZBslLQwoOctqJ9YxDsQ
Y4BD3Uq8U9iM64lg0N4Va4FmNj1NdWaHqSzLNjpM4PHPt4/a1hYEKgcuuWesO5kK
oU07sG7HtC86dtEYhkVd5zNBrzYaNVjXvXYu1B7EXLiHYlWY1BnurmGQtY1Bq6K5
pKgRkIzOI6UKyQV4CJ+edt+O4H45FUwSN3lZRbX253WZ7INX9rv1V5ZjaHmiflwD
du+BSvtgNB1oDY4Pv1z0mJ7EWRntd0kdOlA2XsKxLY5RuVxxTJ05QOfVg8HAXMVu
nNCMJuSk6+GFQcSCVdDK4erEjK0KgndMzzv9meKAVF+92wfkHylRr0hv2+qGjm3f
Gk44UyBSLMs8qaDVk2x4zJzWpcUtcICUm2OA7gB5rkl5w5az1dUlwiucFc0eJhVF
q+GGZSOxRQaHhJLC6XcI6jmRU7W+ZzHSP/VYNLqfDlCO9GEYeosBLLWUhXevbZOP
Pm7F+SSeVcaiDTOsMM78Qpbk1ek45Abie91wESYi1IlOXM+SRMlpek/x3k67pDJR
wad7TeymttE0HgmnCS/lutJPDvtXyHQuY3MY6AJjuZf+/TWWQNKPpW8OWfOeWQMr
3zar5A1ipRnNj7h2TxJNpu2WgtDj1cwKvmdz9UIkUEiwckzYd3D+qftodLunsMrT
WAMr37VGnr/znKKeHUqMY1IWIZSpbfzEZO2fgIgErnwvxYmt08d53CsT5SUwCcFX
KSyzeUiaUcYBEE98Lh3HrGp0M5ajvoFrpmY8LPJYceJIIcT9Q30L8UvB/MCKNE/y
EA+CXZunAHOFalvyU51Mwx2uaVV8GVcCkSswmi9a3s1HBGphZRVFbd6HbdxgCf+z
rUm3XalZRe+QeYQXLDUgYxMOJ/eFDd1Fr55QicjmvnI85Re6BH0q+Xn/GKtouerF
z3MfJyrUhVKI3/hgHDGz7cZqb5xQRqhPCXEHz5f4ejcBbBBWmjgRbIQRp8WuUA/a
R1H4ESIXj9YOOeKQH0H4Dt4tv4wyrwmZeiSavxOK0bIPEoxl4nn5oo+mj4OfzH12
Gc6YGtDedvGfjoH0xGvSUMBbkgi7IQjDHWN2DN4TgTAyxMTarHyoZ0H7Md1vrbH7
cFM36hn/Kf5WsrQn9vGkZJQOgT80s3pi2d66uU/+Q/Jo26b7cQ5XpNBt4y1f/1BM
0aG68bIKbESpFStUegsIOCX3W9i5D3YnPW4W/nf+tnVS33ynKLIFKQzHs8WYPL+4
aFfP61S3LD3+qEOztHT3TuxYWHS3apVFXxHQlVJgDWBwFhDC3ESSxEG1cIte/Vnq
YjtgEdjcsPAMbN8a2GyP2CE5TNEdhNRQHX62pW8qIy1/G6vT4MAwq/cro4JQ3+7y
geSfzql5JCo/2ZnZY3cylcND+dMbEE0qzvFJx33bwpzgEdw+xqCRYA0KJ+rrS1WI
6K5R7kql90YWGoXNgB599zueT0RlQtqWXWF50TqiCWCwaYNTkCxQujl1xC39Q5A2
Z1cIBfa/fjK+WrfUhaZuoc6NNHkrKlnxZULt2fYuhrp2zFmVv1xlkUKKKCCOmx/S
Cgsl2LmbgN5PyTyikWqnqqDDfiqbtpyC7Omktt5GrnFrGiTxTayGTQuXy2xTyU6D
yBeUsMqmEfJDb/y0PJwgDhtIOqvitTG5GS9m3/hBAxb7TwKhjNcCHjz2bMZPqTtc
/DWPIn9JoRr25DoCkV77o3Sqf3hBLcYN0onSunyYoUYni7A7TEQi0s/QB9MQ56GY
WIcaw4DG3hw0vjKlZ5njFgqA4mjWpHvrpUS3A35Q/GHXXQqZ0P4IhOZPbAEJXLTv
naVUClRujEw9jwxow4dWa28ZyNo29feCRLAMSDnYZlyVhSNlaRRYdpdMyrvhXRXl
R6hpKQV24iQQORqTpzHJTtGL95PwSM8ardndl5dUaCN3/u1GMyy1eJBLHEIgI1oY
c7Vw8kzsSLLgwKdE2OLgUhavZ0E2SSlCD2QKb7Z4rSau5c/BVAcY41i4nkEqkEyy
v3bCIx1F8f/hNnBmbNR3fiPnch95M4VmtEVgs3kYtskPfgiPoIK9De94qNDgXVRv
ValCesbDpDkPdpEztC/8MIsx+GNT0RsZEbR4k/cFnfGwgtNOv9oTThQtVvWIKmFj
f236jsl4Q5obOm4V9/E5pmQDzMfcywXmmGh+UzLmIwhHabQhAJDQrIErd41J2LQj
6OqluITFl/yjaLITmNtJeHXQP71P6tCIrCuEMU6UWXvOfotUjUIOeJIhKRLprwY7
br5iovtXUcq2o+WqFvdjmCh7F0tZqHcKsDHe7wkPJwDDjnKZ5MCGAhV3g7zgVsUI
PktnBzfmyz8IE6Tq1KdVPG7nJKL3K6flMPHhHNSs2BWjVeamS3gUo3RSoCua1V3c
eJj1FvOO9GNYH/l7TVfYYjC04a+o1f6cWrlDsHPTvHtL+e/CbyhCB3ncUorxI8rt
F9ehhBuquMpfnGB2Nmha4+VFfiq5v8OM+PquBBGJHXIq+i7xMDsFI6L81Vk8NJcA
u+UvYAlenYTq1lMK3s5aAbEVfoc36Br+F01tdhdexqEGvMrmTZm+xLxbfrjXdbk6
TI8aWUe4XxjcP/lkeHGTV+KWJTUiNUm/SiLVpdmEzcL4obfAqtuypKX2/wXQXFjQ
YPOKeeipX9UzfW+XGPWROspHfUMekUAjD98eM+nvpIO77zJTzOyussT3CDLlBSvi
MnxO8ZKREqOD2dB+hvol0C04+kRgTpuPdioIkFmZ0nBkVU3T8J/o4X4QRl/BKuHZ
bAN9alhn9l0Ws5utm0g6x0Sc4BQcHrviim7hvjH9eq5k+CmouhUOAJ/Wxin9ystn
bYFKvZxbq2lD9nrRBYVbpp1bdyjW73GPQzJVcjP1nQb6OO6n5a74JMgK/Melkq+m
/VGbqMH74zs5cY6/vP/PoTez0u67mqZUHZI7EXK+6pt9J43zXz5Rt5TZBsfp0BYv
3swsiIEnPFE4YV4OkPN3wGYKl0811GdSkXrxBKeCOsBC/ztpOpRBFQvE9aJDJPXF
ZaS/T+AaMziwqIQY8I3+Fn2nBp54Rccyi0gsBeLBfhIWtHNF9Nh0qNWCCGP3WNuS
9fsR+U89di35Wrr7I605hNyRoQ6TnGhmIiTcuETQGFa5LYkNjCX4bEf/93BVDTlH
zswr101KqJpfB9XwpXYIWD2aKm8ujR9Qr+ufml78owm1ZfFyLbGWRQG0oxtASGON
FQwPRpqE9IZVYkins5vKBpN8RBzKQ+3tEo/601BiNZMHGWutTA+fI/mCfuTFq093
dhz1sNSRWrV0l2IxplSIFtMbshKRRK+qCz+OMnHz3tX7axEx5E/MWR9AQkJWHkBR
6wW/AQkFZbLms7efCXiNJrTOaTbJTTVfCGBy7r6aqWynlNbOqdpndy79FmmU1xBa
mqxnNjxm8IZdVveVrvFV78jWx9CTqfBwqZnOI+wmdgg1QEZjy+1RWaQq8FX113fT
0UQC27qQW3BEVEQItQerD/YqFLa6psmUkvStGK2shLTKCiPyzptGmViiB6DS2cB7
GWyiAawJ4Xhphxsc9839Lp9wJSfQi2WITBgKUluQBtaWvISS7vcgbMPduEwyQtcJ
SE2cu/W3ttJiwVxRa0tRZDQOkHPWwASmMr6nToeTPyGoBMm1r6UVUI9LH97xmUoW
+R3dGOOU5ntU8LMoxOaiksG+4RcBeXt9X7SQidFP4E3EhFWgxPlESzcBhf5OCh8w
YiougYvXE2tETkiz/C/X1RC/ejAOxn3W5Q+OuVT7uIUkglOjkPqzBU1winOWfzvl
IBED7gVEHcazNGcJUV06NWF91PuqMcVOBL0WYJz196mU2blTpf8F0a6pm7solOLD
z1G9+v/b1HQ0UlQ3ejv2NN92JQQmRkyuh64qgCh439talfGVp3bt0x/k32iB256M
Dkin77P1c8vo6Rnx46/pOSRFrS7Tuzi1UhEOAnvWUZLPoOBXuLbs+dX7oY+lTUAE
V9hZ3arSfX3M9b6sAF/xbq+ntXqLTFnjJn0SHqE1idWuJzCMUfNww/nXNfx33pBL
gdKJ7BfQYqOIYwMe5v72wYjYkkeYcW9eoE49+ey2BPKxU9YIF+jKjdp95wSEn3OM
yRinP4r0LdJvQy6dCbVqt/8Jf1SNLsQQ6kaIKJFvL8lLWGHWq5sUsQeYAEkyUc7k
kiSUo78ans5wgf/u0GfFS0MRJQml32K/uD/q1ZKMOpbe+rzj6YnJ5y8FruqtnYlq
DQCkchYK1TyMhoepU+JSOiTr29b/cT35FuDqzWEBAJ9dqmbW3iu7MuidH4FYYIqG
a4Ub3dgq9+6PPziecAbMK3QCb+CKzZMBx5avnGoSSshq1fv+HN8ZNgPfV8A5wUZ0
8V5Q7oInqXOaszue48c7t4TFQlseat3IuccGGtnwEXv/BN1CelDl9QbPzPCFwb/S
Ay3ezoiKF0cbbwkukQXtt8GkomDw3alAdAzkGVc3GwxE9hK4VULY1Edfi/J6Xw/Z
PLabb5mF4kdcJq9nWnPw5j9yvtYBivdrOTClxgKEC5VOVKxsfDllnruk/wgmSl15
P1bPRYi+P68clR/zrgctHA6S2kGayoVJvHXfmmu6X9rixo4rQF1TPZ9fBRtw0l8M
Q2c9GOykffML+LGv1LZZCT4ldfkm/3ZIIZfVDa6WC24pLGrFfLXJYJqV0181LT0F
bG/1l8/uIGFUfNiEvoC9KPUflrpIYR8eS5bBLcMDzJDBVqPtFoMw2y3hcaidwlNG
fuRTQYIXd42uTKlTMR6bbTlmlRqrbjOLkygOBvqxMZuU7UMLRerFinzhDvydY3uj
JkPMn/yO4mVytEDd95bQVBT7f8VhidXk0U+2nzxm4Fy/rGYrvlmId8kZ8fZIs9B8
CeGQRbJ8zzNX7HkFS0uXn07QdumYOJLm570g2MBQ266QUav1JO8GoNgoMLYtIFob
BtU+1IT5SyLmUYV5c6QmGbTvhunzQS1OZWrX04eokmOn9od8L+2mWeFjrgVolLtg
z6xJspICO3DlwR3pCXNeaz4rB13DHGL23FNFlqcUA3sxO6F7wkWaqWhb6XDoZC6b
IsAp83MQ4DMCjBT+m0lKY4Zkk+I4GtoHaWYatZFFaDAi4XxhQNURfnUFNk4taYR2
HdZ7aE1bty0ELDeBjsAq+hMgndJapu1MiagVLK3O9OOmqneMOGMmTLSmJBEPMweD
olmfJMlpnEDYwQDYbC4V9+rdslaptL5SKGUDsM1LJKRxYQu49PMoozaiRDA0faiW
ei4f7CUm3DVZAM6bVN3mY4ToMjyOhec5VRIHt23yYM2GmH12G323u4M3GE5uludX
XBcUd9TX/OfEGA64UWjd29Q39wYd06szMQnLJvbc6V53yui5ohMLsL5Ek13fOPAd
Q3sd5A8XWpYyKYydMZzXzmq4V8RfZJD3xuEBfWZbMyF35kOk3BF6x738NL8zFMql
ywpcsGb9PmupJemtLoD1OPZOGr44mz6hxYPH5J9gBPbbNnOYBkLl8sAC82l5cC4F
hUL3/l3F01lMonej8r++nqqskTmn4wqR4InYdUyyMSyoQ6R/wg87Vfxw0uVM9OUX
fFI/wzRlNlYrxiZ4Y6JFmxfZV5hSNm5J/2o0ou9ae5tjiBpAICTIOqWheq3TZexr
qiCV/EacnAbSDsZS9NF+npVAQgsg2lAZiSmYH19R/LJ0rkPb6KSUGg/t8q3NhqM0
5EKF4ewJ3QwwyG9M6DVi8Cpwthf+VbPrX4wDm/wOolm2QyR8jdmyaJpWFpElBZxS
x2o6VOg2c/dZD9K1t34R5/y992BIXAV5LTdDqPb8PimUGB+WBsmXPrFG9jfyStrf
kiSNKdzAe8E7wZbOHfP7xhZL1TIQypzWu7ItEC20tuE/em8g8IjVMP1QRO3XZ2kq
Ic6F0V+jzD+Gr2RnACIgy83691vtBL+/6Z10ls/eQQrNJl1yQ6Bh3tj3hdru1VYL
QXF/gKrJ+hWtX/cAK9gJLGDZABrRxIG1+sOuc9IAkiZq50BzH3mUG3VMnFoZxQrW
mDSbZzCewNJht7m3433UZjalaJSpaPPogALBzBAZiq7ItjjRiNtmSotJCamTByB4
QFVkVhOeebFeR3OKGra6C9V3YYdPIHCE4CZhGxgRItJGxV/hHOCJ4Eb1RNqHiPN3
7ypt1TDe+Ar+4glfRLMK5LA7K15K182/+Y6B294su06KdxOwBFXd/4xG6ERYwG8w
IeSoyVqxEpVvbFB2/5CQxmDSFjXPC/A12/5ZWBlxCJYTfOwsvD0WQmKN6OjYIb4G
MPldweZwXNokIgs+Gi8YFxsKpvcF08jZjDpgFnoc3gscWSM/Wm2UPLLPAsvHV/Ac
B73/oe1haw1sZeKxHG4wbmRP5n6MsHn7fk8gz6F/tdXMc1Bnqf8qFzpw+Z6O4Qlf
RD1BE54JP/Ezylz4LHwzFODEiDTwSZCL4FzE0zi8AQIAa5FQa5bsilNnpF031kWF
pEg/BdWv3fTJWwnHUh8McS1VdJUqjmP4a7ILDmGpTVlZJqS3l4uBkBpbjZxxkDQq
dHlxCGDAElZXnqCjfdlNeIKmYGsjuCRQYWx4BV96IQ7k8hzrl5c5eqCZ16q4Urr0
xjqK+wiRDSDAvTwtbRT0nyXlt1NjUPsDSFzuOFB651/v+RLi72MlJOsuyvKZxi9k
E59BPA9//2SQG2WDW1pLEcXPetXdz/KSveTNORI2bn8b+Nh0Wb4v4p5AH/+BQuxv
X7I8VRYUooFST3xSWU5+tc5p1Ev3hV4Pq8sB1Et5x1oNzD0PZlzJfHScjVJd04Vr
+uQ8l0hKkz+Ji9EYjldH7TOaHH8vW5lrK/LzkecuVeu6GW0KsQ9GLofMg9rHAUBO
ps9NftbEhV/KSFcrAF+GYSrMtXdF8NVCSloucskXhcSTLCHk9kOoj3cAZAbNcx6x
hOFq+CfdH0iqNZpyXfSaLblVCUGWapww0Lp33KbUfm/+PXFiNl0wspIatgLjNyPu
Vtrg4pfP4mhQM4W7SW7drFC4fz/taEOyyS9LyCTyr3hOXTiZP62fjnyhnQ5rQT/L
7fFgiPDwSp3ldcgqggikSlV9NbZaBcWRrMXinHwzks2+2Uu6UsonNLzLp0RLST+4
huoVlc5nEEMfUySE9J0YbhKXjPELv9iiq92vSDYFF5njOjJ3WNbDsDLR3TOrMBwi
M5mAYXCO2IdAyhFhWaSa59OOoUncUWR1vexOyRR07L0mNQDh1FgXay4X7rV8OisE
KVgR5XIGjcN13bkTTWS7fhQ5domFPWFZhH0Yy/umIhVsv7TF5KEeICaOtlBd/D7F
J+zUAUVz03oFKkH9wacnLr1Ns96ONcCg83mpp+W+KmaEaQky4v0pNMzaRsHTGITU
JVmBOzhh7D2AJ966c4c62Ro5Mcm+B7ub0eiDqxYERIPswvp6AqRVmQyAD/S5xSUG
zHYUOm6SoY2O2UJ613mlnWXPK8ff83oA6h1jWeNzul/aYlx9KUxJ7t1cMoBe15/z
wGeTPOWOUbE5xTV2mzzju6IVdyeIxIXcAX7Si4Gc7FZvQLMBlxYg6zuc6NvwdPNs
1JTAnTqsZw24psnGD9+GyB/s++UMNmREkTTN/1khKGDDEgaXKHShtxksfBaOlsse
3hNIABH4WMuKFh9aKFWwPWZIcBfroKJTzjeinzTczOPfX7ZWitKI4sDwePGE3NQ0
cJKF/Iblo5zPrr/zPtZWTWGZpuiIoCoenN6GbqpVbxSakJqHc2X52zlPkUJYDEGZ
UrvGwcOCtvIod/OTPe9gvnwMUjbzezZC2kxGTAdsgnpzEogpWBcRXElzu4FlM2RB
ey6UVg1NU1FQiyjdc1CfmPfQxGXyqnSr0+QWT2JBk15z5YeFAzvb+D2IrfUvERdy
qAQSVFxeuYrd+sasHA6PqfVtsISDApk1Lysp145+6sUh7ikmcVvbJaeEiLapVwKv
k1Oc6kgwNtR7gXHEgl+sJB/GjTtjSX6xXWtGxXrZUTKMNh4eluYojImiWN+omHoU
PZxhSCYklbbXKPou9EwwSgUG/yY6mbCFqA6VilI7viJDIBc5786xcekHHu6U0Rpy
6yT0b9fKWXjzeW/ErmTcEX6+8uo9ujKGnThMZ3xLJgrnXqSO/QNExLdDSDQcqFEP
WUjWVUInIrM+K0Xl1A32dai4odocyBgaAQqsaNQoAF2rWvGnVUxPfMWinfgziOyP
fs192/g0zUpBwtID0BY2cDkkvPNa+y7iV/Ft1UWV3x7EP0zSHMVfPgtnSnbvU+Uw
VDMgGxqwvRpVD/mef5GbrxuoLsGMU2s1MMup6KZPsBeMwk1n9L15Ayr/i+xOe1Uy
XPO7Y2sMRXkSBufWWSlwX4fM6KTzvM2auL0FuP4QA+YJiLyyhGfmvpQcIb7r22zl
iz+A/cyNENwOZgBUuSAjY3Awjrl9ovUF7hqepsFyHBwLJIAgXYXgqC5o08YUxx35
Jts5lozpwoPtYxZb5vsSzIFnkbChQNap7YbJG3brrr3vZ8lq5ULVCvC7QsAxjb5U
APW9px+2TPmS8OXxDmGPBsojiOOYypbLacy0VQIcPJru0q/smocdTeigzIyOvvIJ
cmaywS4GiHm3Fm6mfJEZfGuahaJ/Xl+EcTZggD0uTmjLJb7mcG+EvnE3qWwza96m
Rm/POeCblno5PaiVQEtZA9xr27v4GRjRJHNctQR1GB2xpQMJ9Q2urmgz3rIZsVgQ
L83tXy2tbT+KDdytsb5bflXha7cDyAE56pUmLDs5nO+MV59WV2YM7XThgTtjugnN
8stZGmO8mhc/gc7XwQoo7c3ytc15/m7wddJ1CBAJOajb0VqBP5QhJOvfcE22zkeV
1LJH1aK0mBYaPbJVdFCwHDb1aji+N8LOilhc/lkZ7NaIVkPU0Lb6iz+TlrKI3E7H
2didMh/YXHAXBMz4R1XAC/VG/V4TSC6zgyqZTE6XwkgUL/ovdCBICe4AwN3BTmjS
UloMZ6+OM8WHb4tGpgDvrvkInDYRtjwsgIrZ4EspT44ywmZVBOZD6FUZ1Y4tTsq+
PYiJG8Rjwvq4JljlVWSho6zkPQV2+85UesapM8WZWin6AP94C2DByuHzNxxX72do
npTU3UbwzlBEfeyUrBDubZmH+r0OdnLcEGtpU3soqRukOd9tmjvnRgfm4DbB9lxz
gfkD3WVpHNLpZH5Vg+k4AQcmwvsmWOZ7fZA8jBz2TD91c11q3ojcALQhCihUzzxL
eYUqE1iiwpnnbKKPmzG1NE0nAjJgqsxNE1NrlQQiiLY5vHMlM6VcKbYqzAWBV7W8
u35nt1gVP5i+a/NwBDHFD90RC24Na66Kizfl1o6q97C6vSD46POLBNUUUIIrYSw3
BZ/VmxZ+W7EXEdufvmW3CyacUfO8yuPceRC/K3oYE8O7Zze+FQSn1XrNhrT+VB9g
h3A+jyUNYHdUvVYNA+bsfKtvQ3QQcZlmPJ4J0VTg5jlqNh031A2mZchqvrCqvlvL
VOgmecG9cFl7M5ixQsJTWexyDiOVfGKeKT+3w8keHEvYyu0gPf65YjD6ewzdI7uc
3k6rj8Mu2UMFoyzgIz54iB3XvvWks7aI5x6uOXe85OwkQe9+rYafXZ20ptjCNqom
ZYIx0YZeuFwICNxZ2qqJdBf54MEMC5ZjY/JCI4TSH6VCIhOf9rf34gufXYuY0oaJ
gW65ecrjnKqnaYdMvO+KX7NWTBrEMvMmRlP6Y2GjfByYj6vBziEMLCuS9PrWF2jR
mX42p8HAToUMbeRR4cxAF+P7JE2J3IVl5S/6tEhKRvdkLUNEfIGJe3X/Q5UTz2PD
1VgwitoZSY6vSg2QUc/8d6Sn/QAp9jVhbjD+z0o5TnOz45NdD46yWCkQ6uBzmA9Z
jocm3POLVacddk44EDEgu1LJxjKZOMtPiHBfEzk1b5YMPErmV2DQ4OQhSvsFScVu
+v3owdUlXfcESnQTi1IivarxZkM59N23z5skGKcm7iCPz57fsrCIzXbPHXCiHNq8
OD/cAL4WqgghsbVx0rJbkdnMkYl9RHcGdczhnqK2EftLYUX9wcKPRIFTm3ejRsjM
iqN3OqxZ4zG+4eATLEGk8vhdS+0WvSexbprXRcrUfkXS8uMkoGWd7oeqIJRr9JBl
eFnBR8oIdCfwgv15Pk15jv4AExSJ4WoEPADc4XUbYcrxMNicgmMDyxkwMvor1eKv
nJ+urepoErAmmyOqsIU+xiOoWRH8SfgrN1XcAGRfpwLfnTInCladCzS0FFhYdLZl
DQQ4wZ/54Zs7wwBBFIPoUyPWZiigTJkmSdX9hMOtkzKozyfwPzk4dOur7IAgI4fA
Em+F86jtZiTNGLaVI49KGRCYtny6RqRY/Mi1XEUdF41tHeRuY+JvJB4qmtDtC5I4
hban/zF90JRORP6fAonrS9Hh2B8hzrhXBefu91z+A1UCLw5UZaFOcrgQKOGA+OgY
Kys0J6S2IXumH09LX0rV4Aoq5THEKZx7N3KG7jc7r9v9Z1XGV1fVbiBHIedv+pd9
47IHMVeClPjEgjIflFBRnA9wnwnziFCeWiUrBKLKUlUP2UUlwq3i5iqEvNszEHpk
PBW+hZHQYnIw303hVaUniHIzrbQbUcdD/bHH0LvlW6sKC4T4IBZcbKyNz0TPpXs2
6Ng1EQ7QL85dhGfKPLDYceFaS1XaeOtCyCbtmUP4YgBxWKJQkHeBvzBX+sDVR8bR
oRlirZIjwbOJ+UD3QZ1+MPVBih8+kbPGOLPBRGHWuekjl1xpTN3PvhAKxLm+N85i
EmDcKHXS3GTpAs3YMcoPzSl5saNCABJXoXOCJ0xOSZVp2ooDHLXG/6pT6XnGEhGh
jJbz2VzVQVQOlit5JWAE0lR6qYmImy2w7jAMwv2jJRl80RJYDrp+gsamLxRMnTLh
Hgt5mR2pMw3QHR6jSCdI5Av4ul9YBkb5+8BNZcn6vQiHIlCE17+wsgQp193mKexw
BQEDqa3/orGsUKfGErd83k/2VeImT7+FtxvMZoBUBSSf5RkQHhRAfdSr7/9w2Jrq
Uvh/BWb9O0TgreOpGSAcF1jxmqDNvewFsHeY/ygEJ82W1l6D+ClymLvfZ/RJjbjv
hqmRnIi501TxaaYy1LeTanAcWt+CPwf4SnNzpKpTKVbEB0L4duMBfPmfrwYyjvGX
e946bGTt7x0f4EnlQ0fnMt85oC3jfZ//oDJU+emJ0kl+v+BJSUR/GR1g6CcML3GJ
IwotRzFySL/IJGcg8oE+oii3WUDARVCpWmKhISrG1A2c1ehE2hyoQxUMQtIddhBX
P5KfdSK5bEFtHz8ftd8bgPxdS+GP2pNXPyyIIThipBPKEou9UlJTmw1guSC+YY6s
cdvtFsmykVOFm4mnlM+e98NW4e+xB+2pmmiyjcCKic9qWkXFaPTX6IjRGyznnCja
u+n+AH3ZRKOb6Vu/ZasLqiTL1fvDXz7lkSnGIotOaYWu7k9/agzQ64te2ob74t9v
trXmW0HOF5aBP//amJLsIXZcx2hwV8A6Dj55gfvRak1XKgmgvornVFlBjCT40RcY
lucw4TuLUwm/gvhTacFA0qFHxtAVfTBZuCTBFPzJz2uzocPlikRLSQESY27sLOdO
NffJI82tDmXCB6bsFozIYqpr4NdVITBAKQl7m+sg/LD7ktNdeM8cXBtKgGxlMZGL
D29ii07K2MRZLXWVDe/avqEMAmApHUzs1Q6aD0PLtyQ5bRbH3yqsXBlUgmu4QNVD
SEQU6UtZEKtRZiTWKUsUvIjHjyDgTMHHIn6RdV3zGHxpIWBkK3wsBNr+9VjLlBgT
FsmsBqm+WyW9bCSrCSd5Rr4wzc73zDeNkqNFGcH+juSX6ltA0dUVUR7GpXHrmT/1
M1VgAyiqYWSFWSaWaMNYhD1IM4r97GLXcPLAKqBYbpCzuc6Aqw1tKwYPCiBo8D8y
p74RxUsItzyXd0fgz00g/DbPJycfCvJlFO2GvN6TqyAU8zE9dYTcL0lh8Z1V22vZ
6Y9RIFkj+LeoGcA1PmvfBeEsUIgUVtcAhiXmKGzDvvulEUNsCQ8UR5UeRbaYV2Tm
6DW2UshZNZHfZA9uqwapcA2UfJU7H2mcEvxMploreiESUjaZ/D5VKqaXG+hSg0vE
iMoUxHN7UQhVgBJeiMQpq7u2GfRUGLuCtu0X8e7sNwH3gry7jN+nqDwkt0yZDBYz
W/eyT2+om4RggeIBmJm1uz4XhbP5SO1B29sJ19V5A1iJjpCzwrmkTl4Htm8nxtrk
I7+e7tFMbvmqSD32K9EKM75UYDjVRE7SzhJuhJ4VsX8yVddt3IIuihLKsiElXnwR
vDOlUL/T4Chcd+W7qGj6q0J3o43sJex/YgUSf1thX3e0RSYHCBPugMm/nI9WJmWX
g/46RgkLzYV3nd4knRhMCOXJ5Gn5BAIXeyaBYFw/orFpBKbht4ojIHmaueEIlTkW
aRuqTeLeVJieAghfL9T7+M9PujwiY3bMDxG5iV44G6Ybhuuf8M5vvhLrWjJthoZE
Ipj613dQan8njcTUJppr6yWx9yyJuXTWnyrb1P788QKdr/aIcxJi0Fd7pubu2buU
HIdNbtad9udwezf1Csf8ePeC6N7QcoGVm93rn+40NlN/g2HxCkX5O9FxD33qfNY+
nSyX8jFfst7ANbq79CIvNn30JjAKkamLOZJINxk9XZBlmr8WNIBDasiBaJCKk6xy
/drlrs5uylZgMJLik71q/stFvI9YiR4qI4OxcNdUAeqcf3/cWldEY53+6PvmOLWJ
vd3W8iPhbVOAR3/n1ZiSXf5sOA84FuNsnjkHceA9Q4Q9ZGoyfzeMjZS2eFqTTroy
3qRv8i9qbZxK3mzvRc6HEHC9siisORuPbiYXQ61jSBHxPfgsgozkTOTp2iNyt69c
blPQ9mEzo85PoyMeI+sPjxAHOnonSq1EjZIqfni01h+1L6luANX/tDjkPGfwxQVM
iHXeG/n3Vezk7jZoG9/9WnxORN+9SLDAW7zxK2GQZ5qv06H6v3mXWl2RLuVrNkpY
XqALhbERZWHt4EIjWXnJYQKsGBWWOFh1Pw5HS0zeoDLYXW7w9sao0yAqu+FoTAWA
VYqPmXRga4vfC9N7+b+++MPUZkUyI5bXIDF92jCadlrhrHfJ7ichymW0W29whmzy
Kn1VQ6nJaORoQtQsWbZtZyayz3cplml4K8EqCaZSRbk53z07Lr9VwqDCvdlTcvTF
MtiELRmucQDbsajpof6k0qeqdrVrEDCSQZBReXkrAY/lIIh7YXiei6Yhowf0hcI5
cR/OlrS5IGG2OpW5kzeEprqOfAnvct52BUGTeZFBweV1VUtyKxMbS7qyWrJLS4fW
xb+kyzwJLN7vEG0huYBni33ECtN3kXu1eXdX1oiC+pRNZu3Zvt6QNOiI/NiqEj5u
dr5Ec/1MeKgAtbONxPFrmm38ziv5ONezk9RhyLm5Bk+z2PwwBFhOpVj3uQFbqup7
nFPlbYu1IRoDNuMJbFWORmro1NqbN0xqQqGEvJju/cWOJ/2whlEbTWKwgPUas53c
4vc2C+JYR0euvYAjaddFcI62284p85mU66LubsPceDvgLHIAcPrc2uVOoq9/5RFT
EP91xyQ5zI80sSn004Oqg8penlzoNIpvJu/+KfDHRc5zO44F5DJg/T2cPec6mDAM
I/yw6ndoSUS0ZhyWkjZ4YQB/j6gv33+zu7E3XcRWXzg4abwHaKKvKsGzU9UBpYZw
+nHfsPSzQbXQlEqSYJ6Wq+1JEE9NcDbQXtFmBQjgwIKYaMS09dNCUb/8LkeNln0h
dqh2qz7nBJtTmokzVthSkmKFtdGR7K8hS08shWOYgbWNY4uEci2GWtkf5bOGLg7Y
cOAinePptVel7gscTw9UGqwrDJBeJh5IV96r5sJ7rsAi40r+vbE1KglD+n2KdQZh
fwoR8Bx7lGYm2Eg2qJBG95u4uWFmJx8poSHqzoAKA/6yKuCva5Tk7fodQMcrA1Tz
IwXOc9U5kNHBd6cWVqZx4TxkDhQTZn810I5CpZNOH4oM8zV+Yegwe9zMqjynB/hp
ApugeJPeDYgEBoGOoQJ9yaAzb28rkdnTrMfO+YYplD7lrx41FgxA1jIYR63F2/rN
8n8MTC1c9LQ0+iRICErKEa2I5/pvQtfjHZf5KdIoas5zhTD9GSX63eyMIldsB6lt
G81h+Ba9zH/kt7wG/xm1/qN7/TotnSQSwnv5aPKZ/mkw43xarOFXNDp5A4VDaOlH
5CnlEfAs5/3Fum14j0X34723ooqdNUHdnR2hX6PmtvCoLJkJLYT0pOeEyYTsgSGI
St2bD5UzWpXIHdssVAzwdxNQoJ1RHflndlndBL+N8tEF/Wqing79FaveswrKvXJR
k0shECYzT06/UpvvXLzBD8Q+ZVU35ZztCmvLTQXbLcYdBJncsf9FrosSlr5QGcrA
5haLeml+hoE6MsnBQ3ulOFfuxtHFqc4sLOrNX7ad3l90bDaHiqsOc1QWINC/7ijh
Q3BPlYVX+h+mPFZqspPNkXpmpdGxlkiyO32Wfc8UyNjzMiwe6WjzJSArBMGMiTln
rh2COnGcCQJT3IyMX5JEaRpsMPZH/HhXYTcmL8uQ5qFfmBc/oCLgftdQKU6pXy8x
I/fEdHor59o0w6cvAzssgRgks/KNDqBwQqGVK/MlmKNGqPuj3SuNglCNF7KwhmLn
nHxjqyKLkLR/rbaArMtwzSCgVGGHJl43BTMX+8B1b6H2LDEEh1gWVv+AkDBr6wjB
yUA2HdJNxgy59jmt+t6He2iK1QaqyhMH3vcrj2sVJyRbwmJKtwudOxpsGylLjDk4
MEVboYeBM0hlg+LsiNRn4aPwIydGY3waNDfc0DFQcVF/aMH3akPXCw1DtJzk0vzj
Q6qvHLuMcmOXyaPa4ICT3UQYEUYhSWpMQmtMsaLdRjdsm6PXMudE/jyrfT2osAcY
mbi4Fr+v7d81yp+qUyt9CjheS19cM5XiPYRsaEAUzWb1eS4kf7NjAUk0jCxLdrtu
uB2OoAAKMl5oQdphkolkNKuDQqXVoBBZ6C2NH2ZTZQNlN9XPUvApuuCpeBhgIMGE
ArP5RZBQolmZ6JEGW/UBMpRoFv1Hy1C6BSacmUsYPSAaMOgp+QBkA8GCMOMCGY4F
OgwlbBMJ6+qvcZN23I1Dhfn+M4hV2v5YKJRaxwl610c2e3fh87Wd0QEjmCsnnE2E
mPAWbRUYJ7sgwcf6hNJnJ9kFUi/d9yvY5iby5s2+HounHZQDQhHBbBCHLlVuYSHa
+QdnVCKzyKAkT+o6qFkyl7lOXMXzxRCP9f3ZBPXbwTIH5DWLHeaNNfcFE24lZ1pa
YbhKK0kEJ8n21gijkrYAvFz72LalBVmUM4FGhU5OS4Uiz0Gz+zzvDoygGK1OV3nN
ahkpUeG0ACVoUw5tCxbS8Im3XfpxwOU7cdD1K9DrBIJ3/9HZWz0k5Fstit947x9I
gWBIpbAHgWl0ClmZC5Tey6k7L4hH8ROYtRYRHiC4qTpneQeTanFpe+wuxU8iv9T9
wrRIXVz5Gd7wnrXrdh12S5HaOjrd+a8kTlHN13nVyN6ehtefQRfP11534SFavO7F
riPDJ4WUVp8yaMMaKuRw7tm0EGPQ4ditbropqLKM4gJ+TZVyXV2qlX314lgU4yk+
iTWgla1ichKWehsOL2ksh7onAIhx55LQ8x4wKKBH6FS/EvsxIeWLrh1lMaAKpxcy
RklYZZFKi/egGo1Nh3855oG57eo1+e8oq+owyo/c9mE1QjAwiLGXbii88hjSXF8y
INW8do54S0ukYWHBBjaBI+7VtP/H57+8Tx1UA9PrqhZpZqTn43/y22G1259Isimn
jUe4I3rrwhb2n79efNKnQ4t0kwzeFSEOVFYae/PJlaZWnQJtygBbGpQHBRdRgohC
f4AhAlLUVx/Necc6yXbKxqp4CLGQcxW7w7LO+FCLRdVBAKYzqRt8vYBwlp/VpGsP
uUuyOLtVhRawfRNq03QkmtPlyjNrv/fMN272+GlS8TaMD/4GhNga2Y57VFK09eb4
YfqPV0Q9xOUpbNG6uF1C/wm2ONwk46lJSZN0ZadXxR2Bm19oq890KA4NzFTUn4qV
NFgeVGtEGeUAA1UTEZutJqh76Kgsx0GSYO6VgC9Rmezf2Lrm/TqODxRS88HVooJQ
awQ4v6yMevV+jogV4lUv2hh8L2b1MZz21y/0tK9I0nC1icS7ZJabIr/mlPERQTsW
PNloXMoj8MG+YT3pOVFpatV3LPBnUD8qxpxvCZ/pHQWMA/5OAlJ8H+VS0TNywAbk
t8A/GGvt076F8r9UTs5lzV67P91LA7x9M1u09JA8VOYhD2wlNdEWwUn9BsMjSR+8
3K31xawTgu+HILdtxDawBfYLPEu+kGHNu5WuJUX+QVYEYX7fCx4v1v1FJcJbtsWk
3VewqJCOenVmun9P9NIGpga+RHRGNgIaRhO2MAaQ8moHF6vrI0CGh1HdSc7IkjMQ
yA1XtXa8lTYmrUIKe7RnFgVUgAJVkb+4COT+GNFLLxH6xRImB+lZ9Hh44Xdw13Ew
7dMV+fibyUhrxynKy69mDvnRF/LA6U8/yQ0iRf08u3n9Mall9+c7nNieXT6cvgdF
gS2F4NHBF54VKTI0LqRsyzGokKcMyYay6d2eSRa32QQ7pU1C7mDDQ6OxoXvG7ysB
DMgO3nJ21vCTTl44ISLYOFhX5T8vY7Ti4oQX16rj8D5aSxwnAkXIifBAfb69bZOD
tVgPKg010oJbNd9aXIzZkFQCEzKOKVhnge80x9mQb7TJYbXJzTe7/bueq9a7GYdZ
+37tKLoiltOWcdJUUZMChKRvRakdHzPEuIOY3b+WAGQupuD5ev2IuL3WjxAI/rz4
a0WrSLp8ygeoFgszHOAxTksYD/vWEc4MADjrp/hhLw7O9TATffhQDoVEgE9x050X
mt2PKUMGlB6Mw/lPQRl8tQKQq+rZIPJOjkvnad1wAJR1kWbiQ9bxrFjKuOckuoo5
2EbvndB+5QASIkxLXl+cZF0f/72e1ZPA0Gf8WGxNfEbMiT7f4kZUlxa3eyKQ+sHP
ES3j9wbWevIQbS6Ez6/PUgeH1De8aT/CdPVRPrWTGMAaOHCNRAv5SgMe7SfldERC
pUDjbRnY8bv3dnFIxSobqK9gEeThY9PE95SVhNPxovdDloq8OyKpQiwG7pTdxuS3
HUydfw5JY10Sen5Oo2iRYKul/7lBrjG8ez5Jv7pHoIld8vtNz4WaBfPesgdH/bJh
2B5VUgh5Uhecn8wEAX7JZb8h/mVwURu0LyeKkzP/8ibkOD/EfQGgXsbmq6LzTABS
0HmVBoDtgpiuOp2y4g2LK5hx8N3Zwmz6J4QEw4CTjLYbsW+oTJQnXzp2TUR6rt7G
AEBHNLJz+C6lBrnG36B+YkT9oy9RD5hv153tPwfj9dLH85iAmctIV1jpizhl4yRX
rRiXC697wh84zYU/4AGdsnsH8RT+8mRQ+z+QxaIjdqHr5eQVIh+aUkmLAwrDV8V0
mXu552rN79QdvluEE5QsHhtscP1lnAamMzGB1rj/zdchVyz9cYOaNaW6lp/Xp3hz
08OCkEotJBc7DKxDIn4y3v+i3H0J/fBEC1rlHSBaq6nfdWKkKwV7BrW7r66isnX/
OfB2H9cL8HczlIvPLquuQsB/gHDb/cGfkWRC0ifFRENEptrl34oxxRmkJ2HNAzNl
2Qgzc+z/WiEw9+zSNKRI064UsnPwX4Tiy+ODs7f0KowSVCWBl9EQ4FExSmjS1Sxo
v8mg/3yfQ59efzYpWgbz8YEFU4MoewQLr0BImyfAM78rJy7D1DqfZjh8W1vLSzFY
XYWyOyKqgBKuF6osy9de9pBplGmB9mmWkpmKx/LAtViQzWGeNHuMa/pYvcv4qRvy
Qxr8eoyqs2uZ28RNS25K8ezqZEj7rPwxZEiQXdgYyWKtPm/FE2wJimSUXnxXqN80
wi5ZI9a6Ik6y/0uD9X7S/wnIkFVgdxh4RTGtItoosUyUs24c1McpNiuqhc3qhQbZ
/VNKQhx+g9kqoOTXLRoeJo78viWFD6OaRx7JJ/UtU651y/pEHi3uIhMm4Kw9y3D3
4+orCtw4ClrUcrjTCQq0tcBxXbzewFrcIge5E0BML7/2GLXGVgtUNvYPsXZ0Dd52
XlINx63JsIO7UU2b3xiscRXmHpXNy9Bb0oZIwC1xNuesc4AuXh3wv/KG/20enrjx
LCFCfpy3UNLpUvmRPqID27kGUM5K3SgydIae4t7wKN0GQzfY1cWGuhKvP96hKSpI
mRXqN/+4pv193h1ZHnqmgh5eiyTDQrI1+BkHiQdrmL3aD4MXXezuuaTclpz10DX7
fHyiqrgGYiNOAUp5fI2Hz46n+6f0+6xFX5Z95wUaMA3lZadbVrKRlsSnwi+dFViS
5ZLUx16o9cTr44eqNGBMkl9tMDB9C/JaMg1rxp1eCC7xE7oGhVhDu18isJ65miyp
uMRWb6EyfEnQFpFXF2mEJQIogWFmILtHxyWpgTIxWtT5QIpyNbrCtQ1W9mAlDZIw
yl8sAP/ZrMCXu4SlJ9kdz/e2UOjrO1tKXkQ9DOi3dUYfVt8fsJgyXRm2Ogto00KW
AewtAy2vCxAPmd+bEAOplvpALIkoUTzYaWDsPZnJhEvONK7NurCQBtACetOLsmGv
nYateFxIVOVHhHBOk7JyyKsPiWmvdClQ9kTaYgjLeUIvvRHJwrZaIGNOaSnSjKmJ
C+tr0en/6mMsbZob2sX98HgFw3ZYdXGmcAk+N1FQP2KDaSulrT9T8LXNbcvWeYJP
XegUgNqydmBAvsgqBg7jESQ0XhLnMzxlGIgu4zasEmdxTuELa7UllSLVprLBsGea
V1rJt3DOnf8gHj+ghkAR8mUSGif7ymrFCkWx+CVyy0zqSycIdKFICa+89Xa8eL03
bS3FZyJ/+7MPUAbgGrheCHq8zXBDdl6GtP9ZyZN1VWx83Vpd9Gu0yyu7FEaKqN5I
o+0PmZkEpo4X4UoWC8rKER2hM30dN3JrcVgwXdKrIevaYYnW3DFsSdmo4sZFSTeq
fit1ICFts6XVjPqvV3/PrLvqMQy2zMHLUGPb4SmsNu4HFLmDBrjK881TbOQYsjA7
lgrBsRjn6CieB/vpvdICMti/QThiF3ybG3Mxt/54oare3qqoOD9RtYfVlGCRWKcF
EoZ+UqQUykq779CI1CnpJhCuCibpgIhg49yxfB6CQnzSHFFpdYS5lbYxjOx3uO5V
B3ESGXr6OIwRj4VVy7khBGoXhq+ARvyxXyjykBXmrZmhXM1ujaABu/28/uH9J7Re
VTddmZTE/+qtgEi5c1iWd2aPaBtprV8Q8leg5ydWpaGAoUUBaMUi/OzlDGvlAkjQ
wpEPkvK9vBsQobTNMipqP4gClgQw8v29QW/wCyZgbOVL0mLqMGpZTmpmNdzEcDUc
4q0oap+7vFfGeutkZ9GMHkKoAJ0/KhcGOh/AXWwf1wQqJaawpJL1bNruKAIGRC6G
J4GosiaC8k8AEfY3hVag9yoXmIw640eZFWQ50asvMZZlsBKynoVYTd6TnHWKIbex
5epll7La/5Y8CIEikf02rUS0rEYXR7GSD4xf5BJ1NzcZlsuiA6Z/EfX6tAYkewye
7h8HZjbPBzUlfRR94V/yyJQqGLrGWoVJ5We0hAWJpqiUQhAiQep2M6IdnEB2J/JT
EicMVMGLk3eM3CwedHyVCqRnNfUm+9N7utn1juzYT+bPTds7CMOZh7vXMlV4jtqK
aPEPzG3VRSY8JDmcY8cmNrbV2uUHaXcc9ewB0J63Xx6ghzfsxgU275HEGAYv3yh6
J87oXkPZ/0WoKoh3JY1QBD8vd1PgQ6wP7LaWDU17f3u5tcXk+gg1PhspliAdFfst
hkkx1IvU9l+KLwrbIf/razX/hVm/v5LC2p57o05BjISt8XoYx7KR7uJJbYoP4UJr
XnPMcyyqIZoZsH/XjrIjilG/FiI012kbX5d0ENJdmNmB6PaCO3oRkGIidMevq4O8
0AAYNbo8KetLh7M1W7CYKAwkoygw1r7CS/hj/R8hLYviip0lV0OJr3XX18XEDDkC
PX8VqVpmL114dmQ33D/K7y98tMhOpK8BiMUIsH2+bMrjdEJkBf66xQ7jprXzdSfl
/Atz53M7yNtf7q7+wLF6UL9VaWEE0jFBFgvIerds+DHHuSUyADD6D+tiZIepKTs6
/hi88dZMinSIEl80XqTN/aXrYvA9u38ssoZ6bYPA7qvV36snBfQJmAg8B5ZP6bxD
vddn52UxE9vnTHe5ppYqK8+lPtdR8uncbu8sxpyz74wUB30v/FDfLBMZ5f67JZA0
LCNJT9ByQe1cHZ3xky4GsxhAwnyhKBJesg+RHplDAR3mqVddaQjLd1SsJMTwxgXz
EBgCW0eZ5RkzXG8S7hIP78y/QhZy2aHvWef2VOHpm64Cd7xSUXR4aUKD3vR/ZyXz
x6bZi92AYMk+fdN8shxQBRTZwSzFh4o0Yl1VOaUAccQOeDPu7vOY07+J8dHk9RZn
fnz+qKORxxufVPh9q8rgHBZ4j9yuJQhJVWmnTrZHqq9J/zcRISPUdvXyVcDHORJT
qcT8BAbHCz4Bm/FCGOI9ZIf28JNvuCXEgGFt2LHVKYNKtEM8PtZ5RoJ7uH6QOErT
gYgQENjWwOHL7GlvVf4y5zijtReAZEZDkWqm8c1SeTlgMHqzWAdRyAhZ96mlTnom
EriSetFLo3R2lJr0pB7Wm+QKy0vA/icsnPebb/MQGooOgQ+MPqvHX1vFn/imlpeo
CtgGo8mrc2bt4WnxCV9NcnIW7fyWfagwvhMpjelIr7PrVRAukd3XuV+vHg2wZJMw
RK+PPASckGUcyqaB9pYKNb/TRxqB912QFXJA6P78EYNUxp0DfA7Q+zrWHf93H+s0
IpTzx+uVp8Wuw3fTPz2nZZwmnbERFUf++gWcrbXjrBUicDJiMyyUxROzDoskcU90
HB8mcF1iv9fRwLsXQ77j26jkB6oF2YkRTIE5Xs6xw3BQJOtHq8AloNxNAKca16Gc
IL9hsbwSJwA/PiXIRetu3pfpVoBiKH0N8TVcsseoT0cdirTuNgTCKfmXlbTybN6e
YMB6vi8IbCrfWhWNJu75W36H2e4R3G4rPeMEd3dl5RD2QurIepFRsxN6r923KDgf
Hdqvw074ijaPi+ueur1LWaWqCOoj6HSxcayvLuE6eqxN9GHtco0qhGToXLD4dtIn
NHlehZOD7EZfOVXdTFD7cYlu3RKXwnkVcUcLzrzgwJeNm0XZM7p/3+SHPyubWtRl
p9Ny/I1PxEW2F1ZnYbrlUCBOkG9UCl731fGtkWUhmrg0SLbd6e55VmyCInlJnOKG
s9xjHzF55g5gh6JipaEGKG88UNqXR+Tjg/eH21ZFCe7Y40p0VzEPhVQZIYYxHuWd
LUZrYS3/kh3TbTrsa0WyWzcoy8c0QLAkbIrfwYvkGrPXiGe/H9MsLMbDClc+UlwI
jHnAqQxzgu1j1tvl2xYmmJE28rBT2gzLzJ5y7lbKLFAvX4I5mSRk81cX5T5PBLmW
MHNcQs8Y+618UZ1yzBp8CwXpDnBkVl7nDI7uXbkKCxWRI462pReJMGNhpwt1y4W+
j7AmB2qvOTWyiMruQFIF9svYvyKaUlmVWAcVzx1vWWnmS4RUh9GHvD7E3CzC9nn9
v+TVPnobsKZ1p/Cchkvv1Lv9fA+urnV246KBydp0DF8iw8Cs3D39APdxM2h8yZoi
AELuKmYsBsUFhPZti7x6ak5wjOIZQHrUeM4iczlPa+EvY6KXNLzr1VUjYb95x8Df
z8CS+tMp4rz0I7g66DiaHJYNVujtPEvcItazpImY/VUmtxg7aYDeTChyykl11aoK
1NzzjgatZuBplUAj9TzOiegBbtiuxAYbQiKyPqG4aH2WQ3XTWkzljperhlRPIpWX
H4X+uxxUPsEIBjINXk5W7IYmASGF1C2A/rTlpFb5yR51rVpCOIfBBU/PrQC1ppzv
tg86/KNx0Qg/QRaFm48r8YDHeYyyjKRwliKu0PR5yTPkluw+UfI+piy1TuylRqLg
Cm3zjRh1ZzjOseVBbfahMVWYhlXcLMlTwxYikFtQZurweYyFS5VDumN3Sd/um7Bp
Z1S++FhsWX2HSHS35cxV/VuD7fBesi9WHB7OnsRhRe3pJ5LAJB9tvlvL2HM7pBcd
AufiIVGvgQRZSPHgMCLQvRJi0dRjVb7ZTWgNjy3ZbYIZoy0HgRa5W0cJqoPmxeCH
ur+jPWR/g/JP7z8ZStxX1Ci/ystSSb+Ek8yZzrlBKFDG/GYPiu9NM+cm9SioFeuO
LxwpAMRx0kPmSLBYLjXV305kfwLNjizXm4BLoederAlWuCq8zc4qMhh0op9E/bOT
LHgx6MnEGmm3I66JfeWu4kRqQEH9n4gERXOEZYQ7rbBxSz8TnNWwefkdVPh44esO
rICzImuWc9KF4QJapfiB5TboYKlkjxYqC8ICTw86ybBq1v40XprBQhfQzZBEwsCe
bqS6fWh2TEC1gNPnQFF6MM/KQ5uBX64CNe47zG6t8J5e/eT6S5W82t/ffhcXo2EX
ClXazr2qxCNfTvi7gC7Kg8Os+/DAVs/nuE8M25YOS61eNvt3F3h+5Pie5x5YA3c1
+s4DEaTuDFFcbUUfQhZ4OsGI8VDoVPZSpXfJhyMLL00izSNsrhMnGXBuuOs48KjW
1JWueYjlK8iF/1Mcf1llgSh5aMTZDduEfIDjy3uyPErFpVcdsX+0+gTqsQWgBqah
EDbAEEwtfS4AHUhSZEX65todOOt3wZd3t3DkYWJhUlDtzzetHKn3RRVRxXCfdYn9
UD6JNOq6YzrhFeiZzYUB67mC9+KzjH62xXIre2IdjOxIb2q8eMuJzkp+TRCOGVJq
LyMlwkl1nErVDEmqcLhIf2dKKuZg1xJbhPs8O0bqaGQQOd+rsbjdjlh5kQrmpISi
4AA5c5RHxCGlaipNtS0J9UgZb04uZH4iC2FaaaI7RmcTejo0oVkXLIARajOiNbLx
GUG5HxY9MnKjsSPoar3u0U/aeuC2BkyzlesyJtAI19ypGzOB6LVfOOp9rD/Vfdsg
0VlTI7NkFIFNGtiSKJL3Oiq2bEA3m/l7Aa0BcOFGuzcjKUIL0QyGJzoaP0EAenTu
0DenP5CZ7CMb008xgBfhlu0WiLoHRcVPoUP7DkodWUYWcO0LZMGqNlvolSsS0oiH
XqcXKuVsoQe0qRT0+pGjV2GvcgvFY7Jr9x2eYyMNVZam6WSG0x8pZHNu2Bnk7kzD
uVBDvYfLvIL4GhvASukI8c/CriqUzzI/ixfBRcx5Z9OD+lGjmvioeKrZZM47Rh3G
dY+w3wV6MX1qcmSLS3i5hq2R2w35pjXL0sygZivaHh/Ik9i7wu1G4P4pvc4x3IhT
QrjsUlDAwh+8id34ArtKnHKlLHmNGd7gvJQbxkSqSIk4c36UAK+9XcEW+IcoUtlt
vOG06zmlrdOSv38KKic68ewe5g/Y3qGe4Ba7PNqM9ZdwLE4M3dZS3jYFFljSDda2
NV2O8ZB4wlU0GqWtOWBJnAaHOztkgLP0MYFChUh594Nu4SYSM5O2RirzYZMCR7AB
w8xlKfJadlzFKsDMrCmP2eVQc5NDpzGuhnkDtcC53fTczadkJCpr6izqwEqyM2BE
jJKQkw7YqcSk8aYIQcvO2oDkmNwEASNtkBP08Zo0VfZWOx8ba9qHP4VK9M8JCsaS
gaxg03MBc/HcqjovhPUvkq5yjVkqyrDVE52V0lqYIRvELQXv1S0TSTgGMNaOZPUE
t+NUQAPoIYTen++Yy4v0bZE/0DgjfgTe6xerXaoPn90qniBI0uU+2cf3IUKL3d9x
z6MK1KkMYoEhzC1FDI0WertL7IABeqXMq9B34zhasPmwEkc05nV+7nxlBJjyYdVB
m2j+wrvGCsGrF9+kafGQA0gGtY9AyVO5Q4erVesgO9kr4SCTxS8yAtUepiLxJu9/
e95jV60uwvHtqv55UAeHJM3+wZPM+6yxY2H+cYIiEv3IWUxNuPWQRDBbDX6Uv7iu
W/Rkhl+l+RG3xC8YSLukORpgadWuHr/uVksW8eEgOuVd7wsH/+ry/An4AN91dX/3
wv5ke+gua5XXxBRq9r5Io6V38xYI0PMtIci8oRZtwYFU67IMCBxhn4XD/u9+LQ0b
hZbgk9lZ8ZYpRXhvO/huwW5y//2WwMj43X5vhs0QuCzmJMEi3chPLQkmAlMo0iz3
7Pvb9nTFDuCcTXA7GP33mKD5BlgVRn+TtSprTlqw3J3XQVYufoITifyk37zfRoJ7
sh0iFrs/EQOz7AWBbkEGR80CTntKUCchFO6mFa2OJw9O1NhMKQdGMpsJZLCZfLpZ
EsPzoFRZD0aCfAxgLDWzotP5/VpD3ENVsCulONhcA2rM9gJsxUpSYkt2/KeL0p+c
c878qKSTBkEcUJyr78xRqPaYE+8XAwxY4VEd71aZ7Tj3YqR0yLmWjqHwk1hqQ0zQ
u3Ywwv0lj0PpsvjnTFMLCUICMMFsxG0qbqQKtycfLKznEI9VaadmAqbIaXYXZC88
QdsyqPlhYzWUJWY1sPG/+ViIyi101GdRGJRbofL9b64OCkuptRXKsjkWjHCZWSpO
JUNntX97u8DobtlinKFpEzB4BFN/0w2/NyGB9NnU+VFn3qmsEqVFNJ4wfTaP2ae9
gK4y3wm0bn3ZftNHxYt5idK0MtepkBP8lLt3nRaIs2WF3btd/n7NROqeRc6wYU9s
1TKzOMcT4Bqv4cdse5ZTh0hBeLJrvSI9C0KK9ijIWJRANHJzE5A4xZVJ7tL5j4ND
7F9kmo804nIvU11EyFru1lKuYDg/VYy1mTthjr9dxgQhofTamGwuMoySaJHbvXsO
py2mWzoyFmh6bx57dOpzdPq51Om8HJ2gfsoF8bCH1RLKBwYBLZoBxJtYg+d6R0Gq
GkTKcYc2pfeWCjlm+N1dYBPjFBkBdMKVygCl37ptxuSC7dweDfFTwWOTlJbwHwRH
O6Ttfm2g8DJJhooyuGshTfNtlKtT/6iWpJmu+jhpSjfGBbY9PngUR76TbbmR2DgR
vOomWurG/rekkCT5GxdZF2IkxQONWR7Ohhd0vHe375owX4KkH83U7XiKWlkBCIS4
zrGK22hVydVrinibIS8UUdXk6GXhvjE5SUuerTwZZQm/VYIBcQwzVkFhadoCU0zs
tpk9AI9JkVUFATgAVcKE8fo9NLHrZnNEEZsuNwa3IH2ME43IGIr8PrZWUwT8fi6d
Ti/kz3Ytn01PWrg5eCXxCO0xqhzFI43DZA9CfUsBvN0Nuk5UAqXQxzUHHdhk6qrG
4PfgTs/UWvfKlFEo6iEmA8e0n1GCaVHiBizfmoR2Lly8vnvRXGvU90M1BpaBoNNd
1h8ZDyrzvM/64wVjeOjpyTK38rjTcRSjoC6oIaerCxgTdHghz+eiCiiARWmg39OD
dho/DR6By0zJ0Rqkem48OMQjIvdJZ2o9bukqxfLkzx9gpaKnznfl+A+45vYQyt1l
O1zxdwHIT1lGCW9s/JOsqqIatGnmMTR3+5cVhzk59G9GKBceb6V3sX7NyIy/OB/+
7vmRW1GDghlgRI408o5PgKmiLIXKeiBmcEeD1d43fajXRHyMHsk+fMVLP08VlNi6
yQeZVNxt+5N3ovRriP/cVfINKY8AVzHzevtltMqKNlRuLd04bnJoIG9tUOXJ5Pev
9QkqDtK+sHjOLI91/kuGo5tzVsHdjJVoDWpkvs4OGu8EoMMXOS/NH2kTttukheND
CQ9OJ+VL16jGdEjdZoRfeTHXdnEnSB2w+//kVI9QE0J8MW24gyOhT99R843bZz+t
Y10KUz+ItEZJf0CAfMD1eiHeT/TiRfUyBjXh0NkdEzhunmP8e/IbPABgUdP6+YZz
5K3xAlkOD+r7OU8USH594yzURl+M+w/MdAcWc3AZaC9DvVIM/1GXXQ1xe0umR6bW
vWviyBWV7qIDJKc/nBiwm9JQC8+EJI4chWLP3Df2h7jxedGMesBItdDKmkE5KdTJ
wajZmL0fS5XoaUpy4Kytgytjso0vHuTObzIAEGBuFUAazV/1hA0mriMzBneG0BuS
8gNjGjs0Gqq2cwsIYTbaioXtETZAwGFB7wS4OqZqAAZ3t2dAScffehk82x8AoVzz
HmWv8LtxSnHdd67lCzn2AaNO8lfgZciJ6bVpPhco6QfB4pSMARkLgVWh/fsAYl3i
kVWoM766tIPoQWco1yP2KYJKh5sGvwKdO0U57/G+ZGK31m33sI1jrsdZJRK1DQi6
yjiHHClLbhXAnAUngVf8Kr0BWAL1670PoDh4ob+NdTMhVy/ZBXR3wzAfWCMEF6G5
BxO4wVjQKobMxbi7tp6nGx385i34EKkO6BV2EjyAtwWi9Zi5JIywF8ajQTRZFQox
IrS77owkMUVlUybNM5erzLZYCGNaUZ6Qq9/w5LYXJmpoNuakkGlStYKsKtYTgZXO
Xo+1ahs3vNK+bKRENRRcPglbc1jH4SfInI8888HYaVLSs1VXsBVEfrVkCI8PCFjk
4px/gXbc2NK5k/V5f55jBpyJU8VFTJxq+mRDiroTTzjwD1LTf5Ex0azKPGXN/AGa
7n6Xgn3/UwO3WjOEohKblZLo5eTGMQ08Y1nChWQKcjASFmLXU8bhFUkXaQ7YBjLx
gZ47hCv/iUZdS0TyJZE8YBgr1v2rICcuTAMyOSSNbGx505fmUPX00gyCVvHtOjrw
h+w7Fk9icl5IPL6DcyKYTiAYdXZXWQ/pKE/2o16hWLm6OKJJAotacgetm6ZhgpCU
2YzRncrQnmfUi8vJUjtM3Sq8hLcYM5Lt7IZ+bF3PIMGgfvGllaxY/1lJPlaDcqxn
VOvB3pA07lddnoLYZ/v3jgsAITXRNtRzFO0Tsvyl41GOb90D6iig2Fkwk1NRwyFv
qBcjjYhJycsxHje8/MJ+JepQWzhYsdYROMMCS15oRPjRU8h232HU4ZGPe62pyZ2i
WIk/lOqh9f4g0cEGTKRoZ+tMaO7NrMPHf4KWAyB1vqBP0VJfbb0v4KKYNDOYShJT
PCRd0FsSvQGPnhohRYwIxq+XcIJUHZwRyVx9l4J/0WT2/JBq1MoFKNGOSSqu2Hw6
tioKndSrWzlaKH4JHXVBkXDi1dd141YbrCcveLGd+WRX3ntEyS+KvM8ZjQcIjPcx
HsRELEf0wNMcMZryxJgd2gkS1cRxqevsQ+7iQc24VWUrIwe3+cnueaO61QSTb8fK
yWltNP/c2uZ11OVID5ll0/NduMT2ni16To2RwYhiVhC8pdcYzfposF2GEEvq5J6W
aGg/lkZ9eZjwr3Hj9Rn+wc5TEvSsKqSw3a9u52K0irYu3oD2X/f7MLDJMRcDuEd7
zf+51aZ4IpELCFYRMjcOpiylRfYK6cL9jaPlbwQHV1GdOSQmE4fQoomgZgC92Cel
yePvOwDji33xUXQsLmOW1Xouh2jwTsgqmAxw/9ciSTQ+crez3ky4ZxhHdZlZvXcS
KK0t+SNcX0XCCdl+meVKWpwJdIG5gcROczJqM1bpDLrou/XvGpiXuiI2yyIKA33r
KMlp0rR/e3BmEIjkluG4k5yc/KtYiwl9atS3QB4gg8dtOjWZ7w9sT0T/7e7E3GHV
1y/N1K2CAuzKmpTjMCSBj+ItWaHA3nRLQ02bECGxWgz1EqmQOuVHr4MquqX9WmWB
fJhtoEAIRkmvosURWRzgzQP87IVis9TQyOzEpko/KN46rg0e4638aji8tgucEpm8
UdAd4QBKie8FG0PSeJDWDEKD05MjwXiBPZVVYg7wQDZeiBuUw8wEkGH0b7Y/nDcC
V/Da+2ji0iIY5rjV9ZKMjv9orvUIVMWe8Cq/NNQjAaRNvSe93BVl3cBGDqj2oWm/
rKOfGTABLvHNHhtn4JHHFC4rMrGKwF49sEZVoccxSgwv++Ww9VmnzJsPAQh149i2
eGFQQk5kHBHldMtsyW9PXsww8bJQwYORyIrJt41YteBMc4cydJFat4f/cJXcek5G
5A0B7geK2t3W+o7U51C+hUJUNZDtTYolsb0NEaey44zofkzGgxvR8vWjsXMlqJ3Q
ZFNsY53VHsTzMKHHPVed1rRuK19h81Vnu9fd5tdUKHD4PYiq6Y+Qa3I2a4CAMPs1
j7bZfID4fUQ7vI6W/fMsC99fSWMzyGVy1E6iH2NatqDz4cI7n4WmqXoKdmKib0Wd
MyM1iuFKRqT/q9BSc4a92oapjpBYn7IqThGyYEehk4Bum392hEgZs9u4qLBpx9ME
pSznFpsSfc1eiUg2Qd1I460o5dqo3xvx1jI3toyrfpggE+uO3ROSwDZi+K3+0kDe
rMCNR54XSpVmPhdSZLdCqVllcU5JgK203jo6eD8SoXDRdU9wX6z+WCXLl0a96C9q
nvV4FE2EnjRi1UTyw7hkbJaY0MBfyUZFcDoWLlGCv31bQxWpKEivH3JEKycLziNQ
PcNLumRT9TLVEGzGs2Exf5raM9VEGU0qRiZ3asOrKMwBZZcZ1N3FdAN1uoQIXu1P
Aect7TmF/VJlSsLP6pfOQym5sr+eo7XGdGWaDgBAvbTdaO1CDUqJJuEjxkaDVC+y
yisSS+JvhnJSgkpJ1r7EMwVVSdfY8j76xxpRSdo994xpdPIbuT7UHfJnUZdtLM1w
lsSZzSAxGk3t16vybLan/hcsJtx1H1tjlMQpbump6OCENC/Tgxlj9Symf48pgom2
nRBJaGYejSAYaGjmES9rWAGsFoo5SUXF67eUjohqzMQABsUGi+vrPuHgWwBwwxeO
3ole44yfecia4vEzrkuAr2bL5Q5lfZul06zf8lOznvGYRKyDmsFw3s8y4zkBlcbk
B6HR2vNFQ8QJA0IU29I+OtUMwS9PE5BSpAiDX99Ja4K7N7EVUxxthjqoESsLFhln
rqvFvWZXyJ7w4zwE5g9Tk6K+O0XR0Gdu3ucCL5hJ9UnJpZCpk97U5uPWDRsNDf4K
n7fAnCFR9LLcmflEjPovPjH7jub+F1/ihfdboQ6j4fj8D86UwOJTKmPpZATqp7TH
MXhIHBan5k8perIDx7KkIc93DIndR2OfRzL1eWH9WpkihTqk2dpohwMQSbEcQflf
2lqBS8jbGo9PGdqRmbJ8E4a1KCVsaABWTmwg0a21YGfhc8AEQAbs9tfkbn/ynYsW
DvSfeA3xg5bS6CNhKU5TqBQDgmPACi931sAHUpXNKQwqaITrMGGmiKnMYWWNGiwW
7nTGS3YkxrrSMr261zDzy0ci6kgU9sUC0qeIaph1mry6ub5m6pM/i3M7h2w9tFfW
uEKiA71rDG393RpNC0Qm+mdkS2LSOo1Y1+/DNrCusQiYCo49QFzetjRayRIdhp7k
qSNOTYKw7JLQHEUvLv82Om7wTc6mNWoSXA3bkm5LPYCCv8IAWOPKcz4/htCH2nPU
5vThdcYciA+9n2ouLq8oxzVcBdlDwMQb1guSXBd9lrbwovzvLqd5Yr4QNUE2A5Ba
4YfqxdjGkY41E3pA4k+JSX77ynuNMp0X3zup0u0LD7M3Ii6pIsvyWVgYni2HgiGM
pyHQRGKlBRu9oT+eppcQoJoHb80Q7En6eOEHoe7gNLrkTS3/d2G48S3ha00a3jg3
r9G31PEm97Q4sRefeTMDTyhttd3/fUZL7hcJgCPNbHKLugWgKvy9HKOBD+LDMIJt
zfPBG1V4fHK9knc4jJ/H0Km/YAuhwzMgxwV0Ij45MdWVYraDc5ShbxnrfuDsZeKZ
nQuJ1lR1GdyhtBBdFgx7WBEwihBCdjRaavne8vzZh5wxpHfnTq2Skz60YeGkesKi
F1z6B92H5eSpx7YiwD7GLs+9QOZyDbUo5Amx8VsotpoBlp0J+loDjcOWbq96P6RB
8VUkg4U6KctN6vlG3zzmCghkR1ZOysQI5EnpTQZ2/oaIicdu7xmjWWrOnTMY4dxD
6AQq82gTp/JfNiMTv0YB/WdCVwimCkuZyK3gSLYpZ4YwqfxTgdHoNGpuURhWW0Da
P1+9Sncgnr+J4SaLO2YeKcGNcp1H+/0EwpP3ffioDMfwMJPNwjQFNRSIpc3al1ct
7HMekfDdIkab9lPCAyb3osymt8ZlY7KZlKO3+Hy9QMB/KV0SqQPd4ovJHYFGAoSH
+RB1QGqiq87+HSoIRElu9lTYXZbOQRw9IlOhPeRJUyCyrkG3mvwGHApkf+HjPTYd
zAS+RwIiTaeN4F+jWWWVPtCCH7Igku5/I1+SHSbIV8lxbt1CnhzY7aAb+jguuo1N
Oiy193sOtVOgULdH7Y7ztPW8R/aKXTBAbPBTpspHQ5Z3iftr8Om+KxE1WJYZ61wU
BoXTMr+tJLq+5qOdShs6B35da0FerDahe/73WFHSTxVDp/DOeK4p46vYlIqNajKS
WkJIiwq1yuijtT7r5bgwf/qzGWWcrNKlQdIzftTiiQYM4LKSaXsH4ldZGKcXeDw0
3SpuDWxqOeIYBHFTfSw+9OgDcUY4Q+jCdxlrDtdDcKZecFMqZphvX0nsQ0lMZXY5
j5ohpz4PfJsCpjohqmZoya70zrbx9S8HIuX/fbVVIaYrXf1NRyTSgm5i8V3Jxlgg
OABtgpELsW/MVltX2bu2++rlpjgo0iUEhBYbNQV2vwDdLOabQzsX4SyA/jTiqB4r
l5Qj0n128A5oXhGST7x56iCcKQLAuqvJYcLAqD6pzouAgotNXEFI01RVzGlRl6i0
xzT/4V5FBbK113KuzV3RmIXbbV+2bew5e9RDlLAGhQpLWgNNzPHXKxY8D5jr4WoL
hWGf4icYkbIvvtI6Y+iweCz++heLxEymWDrLkJizkmFBrZ97sa1t+iW+37HJH/ob
6l9Wo4AT+oiV17WploTDnUWQNwjmVk46PXCjyitxVnss5qoXNuJs8KkR9UKfGauS
U/kuqdxQMhBEz4hCe6ssH087SK6YRz3U9y1BEjtKYNR+XBBB7XNcSlVHC6evKqRc
c34Z7mWDHqKNWmoC7bnx8IypN4mK9rZC21Q431pkafswWNT03JLVtWUn9jy52M9B
DjNqTlLwfFtcuCWkfU+JTuBl5HEpOqmXA1q5CndZduNeNGAIigH4UAsMZp7G3Esr
ir8SYjXHE+NK+5y/skQumWs49Y3tMBwUKYLIfrzkbDaCpA0Pff3qzNUOdnX2vMnm
Xnv9hwqhoQgfy8sLAP0/h/gl28Z1LvmVtw2xIGDNchGXCaPWrRxGbFA4268YBmBC
+goE23c8DrPgBEIfi1w6b4C3X1j/pQY3KfcPExx5hXN5xsZYRTxijTfWN7pAx0ZW
HjyhO1rhgUSRUUoio4VRv0LKKCE6zRIo3mkT8GHvSMN1UzmYVoZRrQvy2M8BUXz6
guX1CN3HlgTSlMyeCnsNqI188Gzu41XsS0Gb0TfnUr6rgqSEwhh/KxgVTGd49ghi
96Z/SdIhImNJOYJdmi+J0oPIFhprMhOdnL7USvgaTpk6gmN6VHREk59QyQUACUqw
7KUmNPq8/QLNGfq4r9ZUk/lqhcSVPsIa2Clsu6Mi397e7VQuBHLWmdqAz8aZVyPv
QERZP+O04OJ9fl7ji/k7Vlrd6pYbM/lYZRsAO5zE/E6mn2oSAUDTzsmIZxQXvgJG
KNjFJVJjE+dfJx4hp2fCXMGqfaCx/rgYP6WAnuhtK7Guck9R/+C+4IDYxcWRu8Qh
GAP1zEJEt2ilPcxLpGYoVRDmCW6SgbX4zOltImEy1mX2QmmLZmssg/AId9pldePI
VpYU/etoJs95DHCdt+kWAHHAy3tgeq8t6iwuOgPaB3D3xeiDkguN0/8HmcJ1ENGy
KYJDMgkSkYg/je4kn1QkFtayJ2TSrbvImCNfTASLgnefZ1ECWFhapSFxMDV2aYG2
UzT+HLYz/jsUncObWuo4FtPpAOtGYHcEa+4DZYwcoZv+MRNHhdedsWX3aW/mWW+l
cUpzc+vhHemxOfje3BbR3Vu4fRgPWuCTAYfplOJpo9EwdXItqtw6X1p9MimhhcpV
vvxfC5YBs9Hx8lOmjjRFDNnCXAVl01l9lgFoGh4PjZTFTQqLQADGwTTK2tjL39o1
LIGRRSrcxEotKUunUNx4JpEYVdmgoaYJ4sDUdL2gl1KMo3868nPGpOMLMKI2Vzwr
JWoR1sEfgq3wDrD0u+FVqC7WD5kGcG2/AezOHc1VUyjgUPu7ijmFrwCYYEAErd8I
vzw6hSvaezExL5bSIv6vwje6BKpuz+2BIAgChkAmgb5KyDA0uWNm7bjeWXRMuthe
TM+sNRozfrcZZn+YAcK+N2a23QB6s3T0NO8dLdgaKm7DwQ2iJ3weWVBUph9r2QZb
Ihnu6OFLTJ/ymntVex2ms3tII5uEnvRf51oJ3IKhhUVgMCT5vUuHP09ykIVxtpNr
4sl5QcRJTrzmMiZG7TRkApB0uwF+/l5sssePQlgasei3WyItmbV1SNJ4uE9B07MO
Ts5O20TQS7M8Iq5Llxfd03FtgsaG5Nckr7u9JHXwAR/i2l2C5q4jvqnDq7QwCbNr
hVvRrM2FB62120EiSIqfB8LWwQ5wdVALiAQI8XXyUSK4C800aCawXW9b+8QJAOsU
kg973t9mpgWR9ILLmJoittFwfnZGpvx74kamHRNOnXqiet+5T4NngO5qh+0ZyR/2
HqvaIlcgGbdLewNmf9ZytF34D/LfeBKchHm4J7Gwq4E+IshdUlgzgWCyKVWAq1mu
BXBeW1LYPKSmlzHArEXeeTsbagt1NX5pihPG2e8IeFYwTnjfBRLuBAbqJoip5l2N
0fWmCrWCBZuM06e+FJV0nSjMEFUi6CtiO5XIIH4L1apJwllMCqC/mteqcHcIiQYL
COJfb2Jf20UL/bX8UHci/QeBlQyBDcrLVsWNQhQc6nvO9CsUozYVYvnYdQ+0yevh
Mc/DVGQ6bYlrIgANyJ5wMCLr/vmzH3DZ055qlAFYe07jqfPVAAScph3szLCQZA74
e6P3i9Eh06D0RLYsRhoqo9n9fzNVycl4tu1BuwflWdrA6ziCszEpSLKzETF99qOQ
QJujOm9Q9N6aTqT9ADOmTXDSsyLfJ2fJXcQGTj5S8+mMvB1cOiEh/YtpQWjiafTK
NMA0RbJq5D1jf2O8tXBV2qo/pPJAZfoGKoZ3QqkQr5OI4CXRcA+SbA8onz+95ROR
TZxOddAZiRYseCDLRuCB/6DdBjTE2uDFbKvU0/nwp18RmwXPalCOeK7L00oXb9Da
ZKMGNIya0Gabd6rGX8FUbBcwwy1rZOO7fsrM99v7fJQMGAOtxYK7/q0XdnbfCjUy
vsr+MotoQ05wNjDr4FvBA6R3uCEnNX5h9dTQwFvgaJQF1pXfNcEEJlsgndi2XOCb
8i75Zcp2RWANOr6ecCKSB64WtPfIvBSLeJuGA8vWLmEtIK04tkoDtHUVuk+54XqB
a9b9a/CfgTuqyGKLAyAXO7VEXjWJP/1fyLAFIJi6B4kAtnWJtKY0E9P0qiwWdLSj
uL4AsLiTEuBZVmcpFhAjiuj7e7hpQwJ9upjgKgMLLpVWSSNiNQZ3+aHQTsxPPOn3
C6cAFJGqk3XSvVLjT1mKYY5aV3ka6icbk0A+bQTSSOvJefyggp3rJs5g9YtYgFsb
+PVvsezCbZDZAj3xdfbbe3tvGjACimyBX6Pv+rTxldziVHKZl8lpocNZa2BrdmVk
27T/oiMlm+fv/WujXLZgUn4V6KTDluo+KvMsrc3fWvfvcF4xCbk7a8BAV8JMtoZ4
99F/INzMymU6RZczd28VYil2Id8pHB5z6VV5et9iTmfFSThDbK0lp0JdCeMAVahB
jzpHXb+SulRllt/4QyDn32jABVg7mfkFse3udZgeBo7upsEu9c7HiMusPq3cQxxf
8OKR9InTLBbNqfpu99ZlcAq05UbT4HQ4S29A0aFH5N596JcCyT7DFzexCJMZj/R9
U6iFaMZDR0ImnW+GW3gZZsukUd+e9uBt7BRJ8kK2kOuZwVRNre+vfeTgdoOHJrz/
jS/1+SevOQXF1isjKloxexh0wocU408HXWo/0ZaExV9RdMKjkiH38FtQP/GYnstX
SWEa8Y9Seq2H5oAcEBfXEaQqp7Z6Rt7gvl2ZYlSzcISs0O4uTJ6r2To9X9Jjk34t
6phU7wGCq/+GppUZ+RgpVoGCZbxU6lkEwKYE9EzVSBYar9rsYX/FickdusLi1Vb3
N1Xq8Z1VPlMv6ixOGQ5wzKk+QPSvk7sLzJPw6DYtXpjwvl4gu1Qm5I0ChKjVw7Cb
bpzLEzQz1fDsOG4tos2DnqcVYpDnnaBojnDVVKLX5L3C1EyMAK8La05M6+y+eHd1
bkw3Eeq28+Hk99dCYX0SAEKRPRqKNffryMlYf51N6h6vyTr8G5HZgdeOtNDPIVSy
CdNy1C8nhsPcJiX6nCUJDScgEmLb8tuHqNH9r4G+7530128m4K2yMAwNmSlbnHlr
s1Vzb2M1SdcnxLPfHyl+fw7Vf5/qtQWulLiq3qoJomudECd5gMiif7Qr7ILTH/wm
zT/pwSef2kvUzEHZEFZE5co9JWPMsUzaSF23X4F9Bwjgh8YN1Q3niGx8kGN9X/Db
MKIrvWP/x6hrpu5W4tsli2jhjnD5C9oZZxUWgr35xpULlv8zqgnBA3CQ0BtVVvAz
SOyYhL9DaRbwo3uZa9b3MMskFe8VDUmSey29j021zIo1hVeUPY/f/yuWWOyJyw8U
+pR5qXm0VWiSXjf3gqzq0W2jayyMMbiPgv6fSmabLb7ECxhF+G8WmUAqipM71jY8
bI5gh5X2HUEFdkn8n3l3SZiGjhxzhSj05Fiv7j2hM49lVVmbIGAJo4ThbEBb2lVD
zS1SrIS/Bmyr/UzAcKE0QRlWpjP8LBu6JCGycvWMQYaVFdpdcWc2hrAIFnAnJF35
SLLjqn9SIs7OtRLbT85C0sYgj/A1Q2YHb+2CC3Tt5T3ce4j1Jv2WbwXlMl4KWIke
XdQSfkb+Nzjp2/kLdLMpkxGfMBsAy9CFeNz1s6ANCAOJhNYFZehZFnv0pJYLSOUH
F81Te76ajQ8w6kf/0Lmuz7zXwUdiKlGkIzCMMHq3pr4JQ9j4F6d4d58fGjhty2lK
CXqVGEjvcb+XzoUHXwTMN/blRhN2uqgQaM9LNbiFrTor34ghY8sZv88VajmqyXOb
6YinUfb7sw+JAe612xcZPlde7Uon72tLwvviU4STGXBUWfBg/NozEUewNAYiWVF9
7W3lc+TywQInK0da4jv40/W5wfhTeLe0e3XcvUKLQvyg7ly/DHDlw/05t1xcXZ1t
VVRNWBNkzb8zTIV3ZFlcnRxk+u+pLdyay2tzrDX5V9fuFQfFtbKBe1DTvCGPryum
+PwZdC1XtmwaVANZd/qRs/XyjynfknKDbpaH/Fvl8E2lIurgN0uaStc1aRC/2qOT
sk8yAW+O1lbPUP+xfgTqWar60btgMNZKvMxFokBhZNfHwa+NWFmqDDwvH/rJG/JV
QYFsNPSUCuo/inmZNAyq0H6+2kOyNcyU8jn57FtRq2yXM0/NDeJ6e+14krXvGsT4
CpYWBUgPDzrJGObXmj1uB6iu+fXrrtdi+WHrmj0KNV+Vs8cGSUB99GoPGqlNi87h
5+YEcUA3ctzPGtKfLHLoLPUskufAhI2Z+ceyY/IUKDJ5Td4uzW6cXaOWr5QNhn9q
RlWJiIObfkX8Euzs3wvIqxPEfQ/lLagJqq0PoAdQNx+fk/Qqwgcrf3pIc6O7gEIL
wVagIMssLPYjz7A8+sU3TzbbollS8ALsgEBrISD3qwVh2mM9CqtbjykjSXpzVHQ2
GoPpoKSEn2OZO3Pzb09rUHDTU0zOfhR7EMTdksUC3YHdSqLkkTiN5fJGukPbthf0
IyOHx21fvpjTlyXXmz6cLHgLWwZnX8yv/H1GsSzmCtKOcLO/o0YdYpsLJp8hHWL/
fGGywVz3OvufFfbG1BjP9g2hu93JtnVtSWgRhAEWIdf2Sxy10j8nKG+xweYCBgQ2
YZbuI6ugjRZuzaqv11Jg+KCF6QJGqZMBAXqxhxxLz9ynG/y+UqWOahzE2oq/5Htl
weoOr7j6ngtZkzwvxhYFoWjo2pxkXEwOs8OHw4Lw1reDqB0RgYoUvGUIYIUAudBL
NMy8k4RoIUiTWw+jBSZZWHVs1qj0ghvNh4jdrAB4j+MvK3/2/3tizwfGO40zj14i
Z4ybT/w8jiGVM+61vaJmtMI8v+PQ4uTaSXDhKN347OdqS4rmm+9tAyvdz2CJEPr5
ROOJ7Mr458v6zF0LW3HUgcyb0EAL6nh3oxAiknT4JWSzXSTTvXuOOYcsmUVu4+9C
BbDyUVi5VYCMo5Aj7N0D/zmpIjgStVnhuMMcr/Gk2GE1VcDQkb8NU9UjLFksLRRq
n3xhtnrSFch2R4FzzYSAmc3ZVM4hsngSTooLuhZ84Wmy7cnFBaq+AJsg/mHMXkV6
/Wkv8ZqP1z3Fb0a+Pzh4pz0BTNarPAfW+igmWZF5wyy90TzIWcxHPXVpzHGwhBCS
NQyQwz3tJm75TpfoPJBzH1fopiH7OIn4kGUKbNVX98tj52UhGjpnck64qjEVW/86
Ob82wgH6K0Be9VlyQPjretc12x2iScBgw4Nt9ktLYLue2yeU/Y1Fg1dKhME56JNT
2PzrpcmXt1Bf4SZsGplqtu2veo76wVLXv+zvfMX/ZubsPfH6pdBn3Dv/3tCBnj0i
XStHE0CaOHz3rdebLjlPgCRFOQKoeQgPooSJzzZB8OB56WVSXAvV3sWBn3hmBahi
e88v0Z0mdZs+JxvsMZG2d/kSlgkOvNlymIu5nP0wQvd+ZYfQt4Ho2L/uisqFiQ8g
p8DYBVnmGmGe4elrSGS1EtPhLrx3AM9/GjbXtpjdxz+5t26JrteeSB7d18p0l148
QkDWwFDXo5mLiBLrICJ3KjNIhkiAYJfGoNEWS3g2HbbJgzcs9kVNUUAFrEQYi8JR
t1jyeMKTWHw9CMQNF71lScWuaWASaFmABimvy/yVwckl6SHrtpk6rc14PfGWdho2
NRls5tfB+uwTqLkeihhp3Sx1XJvzTDx/azuc032JxIVkYusOith8d7W8Zn7UK7V7
JcaJe/4jBqAAoDuz5N37yITvtOCHdrCMVzRXpYOeZl2rxCDGnzKMv3TvdDfI9Rcj
kfItV3VAjSKaneEjMQnXW9Mof0j+Dyb2InWI75mTHJ2ZjqHSVri0kZgpmCOERvVX
YTD3WrnOa7C/CEr5/gA3ZEqiwR7ega/MRQoLOgl4A04wSA8CKNEknIR0erIWjgMt
Sr0NRm3OqPyDnkqpa8lFAhnexc6xj9zYk2apo9kHDdtZtKNR6Rsf5gxM3IaVYz6n
bLf5DZ1uUdvLJv22K/i7QnKnxzrSyzSmTLzg8o7+UiFL6tt7jZEl00GjVyvjdoNi
tzwK45SLhqggHu+9LXYL+K/ywBMiTKpt7TNphdB/jyxWxTymdGBotUQugesuza/B
Q5aiIb6cXILXqa9D+gBrJKI1aOW62shCyDW6o6TndZpeh05NQkFVAOxQO7sKG7ei
spcbMbdR6KbQY2vmnBnS9DyRla+jMxQiV51E1T2bCDvZaO+uP0QDFGVpSgqLXsEN
FWM9LORypsS1sSqof/EtKEgwCv8eE0GE9ApKUHv+O+rAmBV9U9WHcXixF5IwM30a
ecnPCzp97oHPes7S5HBOuiE2NbjIU8aYFa5SzR+Qf7ECAjnjDOzIslvHXI5N9geI
IxdFOiQOXVmbu1mTSTWTODXUeJEmMGh1SQAQDIZ73pz/UP4x8g38GSE5nrjfW2Hs
DfY2nTEbVu9RqJgJjmgW+Am6q/1npFYtFCWIzIu/y524J+1Jz5VbtyCurBxnGrqo
WkYo7hBDCK6WNdm8gnfdM802Xyk3Oq1qGAj92hKY/uIF9aO5rbys9/vU0DyG65c2
ns4hmUMlS8rFm8gzde7NyLEciNFjStOQtwgxbOtL25Dj9fGbYlt8uVABRc6xb18k
4lGy5IViw81cDjf+GjJYp7dDUbSAPxcbvSAHZ/PvachiJQAA0lenb3NhWXqW7noP
EaydRhHyr+LdC4D3GUfb1gA35vs3VgbQ+Kg3I9AB6yT87A5Rt0DhFYPyFR+7xAH7
PmOeq34XqXqfD+wUZv/BZmFQAeWhHVFffJ+oB5AkMS9eIWlYL48mT00SuqkIzQEm
1eKcBYoj0nZlf/zAKeYUZ06XN5+sTzmJJz9ZqvhRYBnf9j1Rch5zduNsgMVD6l22
wZGYg8YBI3FsxVHYWdRbywIT1Qacxp8kKuTiztz/9wsF/xBrUxh2hpga0u25ijDo
cQRs0xxBWwkv9askJrsThIm8XwlQ+GF+mPW3Pla7AoJsFuIITJKvDY5MRZ9ZE6jZ
n2U+oRJldb9aufKeELLrnyXAZ+m3mAhyAf0N6E7lKpBcyM7h5WzzmtA8PmSYMvBF
oXcUNEOcDfbC6WcFlA2R98bMLQTDGXp9dRSSGHt7gomlhp4e8JZ0kAEIN6HrTilz
aXcVOxNqe9f/8fqGmWzBBVh87wDFcajO48id3MOb4TKa3ScyZdpVUf0n2Cj5JktO
JeiVu1AwDVxuylBtH/YdooWHWu4SpmgSeeJ0OkKv7+SLdK6cJ2HUxtPevQklS7r6
IAGtuDCkN3FUpxgbk6KgGDH//xsy215BgcTK9eoLahWhjnWMpueVr6QAPM9SAeEO
VFS7OHwSa3o36e9Vv2W9WNJNBMtqPtJy9R4PAAbHoKw/cTOBghOUj59tlzHy9Ruk
/WFTlJJhejjmufOl6jQUCvi5pu8V/gqSmg5Ri55pBzM4zYdxHCm5pAJJ19PHGME3
sAaU7RrHqKgSYevjaV8rSMaTgB3cdYW9oOKz4NMD4pQtd6TqnXX6aEQ3Xov6lQcD
n95YXT7tJxYN3zOyYUm4u9wa9HbhswNFPMr5DzMsMj5Uiow3PS2PULEvqIVhFwDB
6uOA8JO1y6Fqb1acTj2oDPEbqFQVskRftRdxkhyuuo32USlE0cViUFF+uuhQyFCI
FaGXVOuKkgz1vm5JLCY2Iii/oFtou6lRC7yGpLqtev4VMS12kNf1HJsq5K2ijE5v
7p/uKjZ5sMyxp13Z7NP82cWVpF1VFL1I/LrhZWO6zI2HZURcwj6iRspbBLgv10lX
1gpFexej712SkhNvkd5IL+T6ghk7caJBuYeeAPjK/SbGyIFfNpWjg7hdurjfTiJB
ghuL6ahbT6OBdczyfaqUb/R8F6gRqY44sPH2/bFFCTq6A1hWeq2zPe+BrdmbVhp5
5BZAIn/rLSrUb9nvVCQ8O7a1AEhny9vV9KZGQe41QQ/mhQ0leNgVqhYf0aAiVZ2D
ebDQfYE8+hND9OdyllKwZuiNGiWWgQlctQrReidcv77qi0OgL1OyyFYkeZJI2CJz
57FQyDShgp/Happzi+weaMPBnsTKINl6RPifiisGyJUZfyL6LxqCxIdV/1fBciLL
MNc2eCWKWmMAHmFjp8Jc706duzYrZ+7bqTuiwvYkMiorlnLphQ8mQ/WKq40gSsjd
N7UcPK+TMRJNodt3NX9oOn5iLOjXVTvqb3m0aYFMefJ6RFDJ808ObBgFID/mp5I6
0A+yTZbZTxROzisj8WBGGwREuacUR1o4XvwNmyHChV+zC/qyEJ0MeOCtRmJjOrnz
y6kp1guW4g4PmTXU/VE4y7du83XyYwRLR0QCFGoMbSNmBaDO2EnKIfv0r8LMG4Pc
RMXCYhNiqKkkpXbpJ5k+aWkfnD4kSKNyv9BRWxuk4SgB2WHmT6Zzc/S+8mcCnFNz
hlasoCAdT8AqnQ+GAJLHG9K6PqqQXQPNzFSTK2PYQ1IQYflGWj9ofdFqO8gfezZ6
AZoE4WA3G2b7KKR2N0Kledo6riaQgkDt768mko1VemtytsO/6lcKhuPpvYqEQMX8
VkAGrzasGMKS0TdjzQcecxI8EKVEi1FAyGVSpJLkxf/Jxnwxd/mF9M0ly9qAOITP
6TyZhSgr3+1wqPkAdeFBSE3+qHVQOUYY/iK31Jc3ZXJOHK2ECwGNgQrlcLHGoyXg
XYumIMBr8tbABRa9XDz/tk1nfsT3hPGHqZU9JQfrOe7o6AO4HN+0LV5sn3ccaAu6
uwFS2EKu9AnkamNPBPyPHGQY9fUHmUEcDg9nsNYevMdGjA61KyyDGrmehGpSpqDv
KjsixV+1H2VPTDX/ukA2gJ1P/CzCJpZ9IUVs8fv4M5jxCpAxVJDkDVVx+konA7mm
er9Afqi2+CRZDQN8TrzSCPvz1A46VruMbhpfykHS4hPFpbVtUYpPCllKk/KyEDIj
JhAWRJWxLgLCKlV2tBrQE7+9Rxjqo+J6W8MA8oI4evRQVie8SN8tZzwRVUuUECa4
oSv7/dFStCTg0Bwim3MeTT5t4JoBkB2oPrLyLfdlhQWswZEE9OxIobtDSRsP3X+k
yTUVCiajX8+4AtHXJAGcd+2Yt/hfY94RAuLM7lyZHptXHTo8x/hH3upZC9MuleQ2
KKbVHMukuBDa3yjt9JwK5pwzs2KXXUWSmPdb/CQ+RBL5qRRViNYVLnjh2bBxkWtF
k0wgo5e0Z3GaeaOCYYg4jPJII2tq6wWeNM04Z5qxwpt8Smvb/jGyciDgAI+2hRC/
UMiQ6+8EV7MFVrzkDK/2LHYW50Lv1b+B78PvSwLVdGwfBR74wGCfmbi3xL6ts+ka
jtIg6RRyW1F3eLPuNeTCttut1TYi3Tyf0wp5rWxcoA2ZrFKKBXZoLYEBaZ+K2Ute
O/FDG8GNq6pfAF2UUSFSyHRNeqXaoMrPKmfHNn5vSAnMuZ0ah2oTEeqVyu0Xj+xU
cdahUGdYaZKkkEtPaBDZauiPtP18zIOoPbRyHjAMGhwcOyxwe482h7sPehzeq0MS
fL+TidGrrFxG3IPoIUQhvBmetn3HiUDuByunOHjUnbIQhrnH89LMPzhN93eGsgQs
3UPO3Vr07mDu6h4hsoa4EbXKi4xIKelZQfnAG37K+3g2a9vB9kJd0nTzT9IKMJ8L
zaYeiIUzsUM5pB6dfJ5De234xTzM7wSZVaF2+vPFNvxrhsgx+Sdq7u5vmyvFZpEK
sm7q/84eaLldEo4Iuxu7O+NuBwJg+DZ11lNwJtACd/zRD+LS5KSKDO70YnLH1+za
z1ZIZDJe4p9nxc+xBoYV4nNxbb9knuBSBiNAZeIqh3eJZujq7zIpCoFP9thjmOuV
XH6VDS6+onT6uQ+yfgP/MQV3XYhx3Gw7mUVHLZBR6yCgDJySwXMZsRSw0qN6w1Kd
JGRB1KGvrxtmoaOCDVpjDMjVod0RuKs6EK3iQnSk+AvkYWuMF4bh5Lu3bJUz6W9I
4S0ekN2XsiPxYSQwBIAuUcIXpESshdRXJOtoeaIpHnT74mS3Ji86/GhCtmIsPn/D
ci6pI6lP/DoJ3JFgc/KeBbJV0u2b4Budgbq2Z9AbdKMwU2ciIe5b7boyeo1tjWbU
7ILnbg2cRILGB0tsHwl3boiJi91BkBB67SyafIlZg9zF/tL9GyVjiNU6cldP9Adb
pJQZjwDXyMSGI7JIpC//50aqQW4cJxnckjPrIcDsB83bbc9bFr91xmUY0i8ZlMfC
Zd7DOWcZnAzk0Zo6gIsH9EzioEqivYqFxriEf2V7n/GkSg8012vt7xpI/14YT10d
oNA2VY1CxofLkQR6YmsbwjkEzCUHx3H9C2LjBeWYMWd2XLCpBYM1i6uiCVEFE9Bu
LlP4KdG53yLrK+Tt2iWg2Tm+8NXOz1ReFVAoq270pYhlh8IOoJbcDWrddxisvTuw
gOyLsUY8A7Jy+5wX8XD4XbarNgyu7meTkEbDNWdHczeyfsBP0H9qLymjfQ1EuAKZ
7Ws71ZYWStZViaTmx4H5Blaz6uVX03EhgOG3nkw59Ew6fDxBin7u3qW++CEmcgWI
AKneIGwS2Pa6MTS5pOrV3SGfcid8hcxPLYGUyKY2KChOTihgpN6QmdOD6+q74Kvb
jkT8Zi1ZBuZM3ysyVCT8cE1lFZegHz8rXKO//NCumxuzThI3IW/xWpAIZGPtHeix
pSpKhbOxZF+COQ7labrRMVuins26bhWhJNYMHU5JP63NjcsSCae78rVf2mJLsVA2
TGEHQYsgmMeeZ3cAh+2zonzzTtxVdm06A01z/lXpS7zIzG8AT6pR1xD8AU9XSKSr
ZdHkVl55kdA3l2gl8GnjFla6M+FCAdxWmTCt5X9tOvpeK0iGjvtBl0C2ECZ5V32K
VdtjXX9gXJmJfXGV9pe5kEYQTfw3YQVzgxDMLK0i81vh+oE0uBpesrzW93Y43MtI
t8XWLd9wj9DqgfwoGz3xV8yM69q2mFuTUYzmb+UtPCTLK5JDFE3rWZjjxinAerlL
EGlWy+QEPCZM5CE/6S9Dkn67hF/gMjk7nowjLQPDa53N9ig5Tl3PgiDFurzSQ28f
maLxFSNa67jDXi2wkusYspN/GnVcnn+T2dZRfgKAnaWUO0OW2E4tegWbdTtl6WGZ
WAO1z1bo1rQKW2REz/0xmHm7/CiaT1N36EHPtxH66JkJ70hPKi7omgpAHsK9dZj8
7wMXGlePgpfh04sb4OpC9HwNrFsEG9WlA8r7HvJISTAS8SyGeHl2dbXcsKp9gDAW
jhJkOEYpWAgYNxosO7Z9AEQ/osGCqM6sXke1bXfTktmrz/oQlVMPz3luy6Ee6cQu
cqgr5aJsHj+HYn/leBVMVZ0MOs7+WaVxDvDiRQpJet5TgoBrQ/UWx3IJFFeL3Uje
j7wQCH4hr5lJE+BjGvnnQo6Ij5HB9c6ocLZ0/MfdnO7LNTn3jenBypvEO2YiyEIN
8Zo/a28BUo+CPmIZxfndTdlaoOyG+sibe3ZIW1GXvd+OMP+g9ymcO0RVDDcKBPPP
bwIHcayZWU2m0IKdRew/EiCtngd3gdcK33oi4KKLuQsze/SEIqyt+MW8ivtrr4ii
xTd3tJzcVxd1f7SXFP1FPLin4jNI4GLgiaeaM4Zf+AeStcjrnAyQ7U4luMdflELw
Qy2xiuEakI+0B/5vNXIE2dxKcAfYmTJjXhmvnQe47ZyFKOaeMjN9YAs0eLjca9my
f+gDVhtINmFes0AICqtnJtDlWh3ilXUe3fD1NdJvPo8MgqGaeLI419lxf2djwF0e
0vCQdwJ+veaZoNsD8h1VZcUIJHy+nd/Qvib5cN17n57c+Dy6JZn1YIXZVNdCRLZI
UNc5kiUpAY9aIyBN654SDYU2nptaXxeCO9oc+xVQN/LaHwQu5V4voQa8whTX3XFa
OyZm1aHogCFlosaY9voiVKepexc4YQImVNVXaFZbJO2lFKYcu3cos6WB25tlutVl
SAQ1uvsl2RxPGPbSkPikkFXVYQRUcNwPOfKanbBvO26tAaRk85aaCIjOqHjV+et3
0SFPojtevEbG3+zyMGzSGZVnR8e1D2/3TVxBVlSCtq6zESQQoUA0p3uP/XQopDCm
u7imYrHapQt20fYZptvLkudN/FjNpSN6Bzu5hduMTQUP/x6Ca0jPmX17enbv9D1u
+YJdIaUevoIxpDhAxzn/1cvYfF6lrX/wuFxwdlSKneeN3M9Q4v0DhZcU2ls8YJs7
BwTfTZ5Qqiz8+r+1sjlRibE6ppdBK/FhGn+usvjPRQPLP2jjVSjDC8aZWFzSO8dQ
EGBfyl9RdNWWrLD6ATyVk1WzhJSyhmSRCEKkTUaMRG9eLY7IyJPn9xWeD4PVYli1
dWygCR/ltidLkYa7uyCR0O6bgdtIJAzPGLU90s+hDiRQ7AtqRN9hkUNpCIYPJTmw
S3JAx7B1LglQt2cW+UK/uyNBacafmNPHat1+a+c4vC+ubQUCyW1SNUVpbDiBYmRC
6uPYtW1W+DUu926/4fMPmD1IZOTsSifbbZSnrZc+2k5GKOsGgy3KwLl2QHXpMnny
vg/7gB8AavZd4Q1fW4rxjCPC0zlHwDCujahtCh9fHHVHeb1ufzlu6LE2sc8Ukpxj
eRluzR9Xr6W3zv4MIvsJeGgxvuTOifR3kLYlqxm3qcm85ogFXLPTrX9ofrHaL5uX
qkyONGUDntEh1sM1jRDqI2qFVm64z+YezQ2Ow2ZxL9UdwIbxfRSuIZAVWLf1sg/P
m8Vg6fqzhzdGgX9weCFLjeYkcrkGrpUy4W1Lp/Pw7zKQQefcQJzif5jQYCfwQJau
XIpHLk6CRsTny8z6tFcNNAUWpC+W3wy4S1aBKn+s0GHWsBXDnE7G62VbGLjalBsA
fbNEzD4QOAA8GdFfAeacq+APgqNm9mz1cuNtaWZnKPCeEsrRvLx3/qtaBrNk7zTZ
dTIeFd/TxAeo/qzfYmWf1FK0ec0RweaINuv2tgnLNoxyXP5VDw80mto5c/nPYAPn
F//FEcKbucANukbG6Qb/ShICd+9miCNmhKIse520RMFGaLn5786iT1yaODTAVb0r
we4JBIVSFlx2SWQDNC4snjXp5xakRouGx71QazPgOeq2AK0LebAkUA6uqSqGXAB8
zsXytivtABxrToWTVpAcY0vLvEQuh5y0uT1b+tu2eG+bXKCIwN3HvkxUjPpAi4d8
cMUcrUH8w3mmCIDRTCsyhCjFIcy4jNB8JKdloUDENJTbBJagkl75v38LiUV9D6f+
6QoMnUO1w6Pw86h/N+7MsVdwNuKDN5Q7SQ1vCLVxE+s6f17CMQIl7Y42Is67aO+m
iK1jFP5ei5FMi85XNSUILErxi0hAVN9BPi5UmO/pIT8sJ3yCvrtoAv+zQDhS/GLH
ZSDP3KDtfptNEeQHzkugCS0n1PH+vO2IOY2bN5zlR2b+pot4ozhh0ZqYZIfVqULe
ioP6hXQsdTN17+9F52E3nMK63AsVuYTw01eucT04lyXwDaN2nTpaasnk58pZSDso
Thf636OyVkYQZLBnAs2u36sQhFXZuRGYI5F2l1r9n/0eVOeQlEaSsnCY7fov3WHm
n5mwIeC3FQinZnsOf6DPFRBYtkoXZk/W9RcIMQS1UapW797RPEss8QYzXiGoWya3
P7tDXrmfeWZiWM17ynaKWZyF/GTsI1pU/5GQdX0t1AHKqASjoyQ7hKijRhyR6hNP
4Xu0V8fMjKqsSqtggaPoCg5jiOKJY8sxRt9S2+2sFEekUxdgXzEsE+fQSdhyJEse
gIPMrweG3EQtI3SEIt6555JwQbLzLL7ng718gNYUINGe7vthB8bl+RtToghtB9PM
E4dXOfKYxT6UrmslbTYIAGl0fi0ImxVMi85br/XB46Xkw0PtfAFFWHGCfhKGtvwc
fPFos+AFQ3i4FpVC129GFwhHY8mOYkLcQr2R8qHPwuzxUT9DAbWwcz/0r2rjZl41
68ez02ayQy6I0/j0IGzmNsKe8GZFE+zZ02jPLOCifKrBeEPRMXTeLkHIuA3Lyqq9
Uf7fAWbInu+UP5GrWC2doUpY4WPabEOywKIIlGpH5MknZPz6/veU7nMhhLCv19mj
cWHTt5FSgmjO4CcK+Is+axDeAXuQ/sOaOfLXzVU7I4/3ZOOmogbOJ1emnlZfg8RB
eX9bO0FUxKAKeKEekiyf2UKPXRGYY/hLW/f8gaX/a8SKtmtJWg2jorhuHsamDtsp
1VgAuz7Hc2311FN51dFKM9Sv0ms7CY2AwkWqx/Wje/WBBrhXaes+R+yrVzNkg8LF
3aqQZbB8buddAPV4Uor5+j088fdtV3Dz3XXcqOE4fpFBTPF0ZzjNh3NfwsiaX8/m
6AE1A7CfDT0NL3ee+PhHyxKqNu58QQBlpo0jNbO2Y0sbiECxjpdJVuJ0RNVdpRE0
97+pFh3JI2WJJWI+4mga/QRgeCp0iqUpX8kwnzEEVlWO9mqe0ZHHZDCpAPPQ3Q3e
m4JyZeoMp+0X9mgD78xsnMBv4s6TR97rXsVRuNmgIjnf6Mm8TUuviAgSXXeN/s/M
1Y9UGHmEMgOJ/tgdd7IeoP+zr0nDPZjOQ+LaSWnyjMbSiSZjLNkEIjoYPoayzf0r
ZxjtQM6jcxsj0lBDvmv2Zvmw7hBLUejn78VauDDvWX41mhsLcxJNdB2kISIkZkkP
Bj+zwYH2bMd4KcTuhe0eSYEgXpvHJnagy93eK4EU+XxW5OMr7qMomaxnVYru79YC
ZVSWprcdAfd9rMW2PjgUFVwqtuLZrf8Np/6wvzgQJQZ1O8YyKM5TZYqXdavsTibs
YCQFlEwJG/x6bBbgluGjmRC6DQ8TtN+az7oWcfdkiJw9VoyLOpORk4XAKEkkJ73y
aMKmm6BM6tyUq1c/Fl/YLOAydNsBbloBpRkoTrfU5JSgu3KoddwZUOys7ZZUECTB
/OalyqPF/VUEb7gfDa9fF+emDLN2ePol8SDgH9s4xnUUeKVwDcO21MMMh9CMS3Nr
mBrGwhZf7453WmuvlIkS0E7AD73TTntbV6H927e07F+RbdbV43QEKtiCKv/hZD4r
jBrSO5EnkIUTjs9Y/GuvRPJ3bLN8rjLm7JXgIcIYEWqOnFk5xqtjiA55fci4oztG
u4tSmLocM+mWsIYTHE8j/XHKvI7EJEUmRoNopL292BcPKeb0JQuWasuyJyc32bse
yrr477WeLsJVGn/uvNPF0nP3P0UQ6INeHHaWbtXsKP53TQ6VSg+76Sb5QySdrdon
2qS7t1ImyYRjMg10Izmn1uVpOPtKfd2frMcSxg48KKb8v2a4Jkso3sAIpjP1+4OC
ZBrlU8NTanvZ7Bi4oOb/IzwNxBFr9UIw53zMher9HPTiqEnBIfsqmEmWH6Y2K3Gh
5mEtWg2L/G40pYAOnBIdhGvpFIkOiMKSnmOm9lWe0zy9gq+lhvB9thJPaNhBETtp
YDi9wejzxdsz/UUaLFPiLonfii7GGxxaoXRtbYyLq31jp0gkHuPbHYtaYqnWCrEr
DBo5cFFljeivJGifC8K3c4zZ7I4aaOIu3ccO5/6Y6ICfS+Ovw19tVlEoZXnV2zd/
rGb2xXIMSqBMb3nbsCGt66wqEi7A4+f+IR2Icphjr2dZZE+Q0rD3rQa8VsJeDRFI
5xF/v092TIkGQsIuSk8KWVn3p0L7HX7tQ6gSdFPldpL6bxbUmy8q5TSgiShY6HfD
P1kaHf+pE/3iuWRqOrbV2a7uiQp9Yvti8t6YPaJPEXX6a122cgmXThtVWBpec64R
TFT6MFXtbL7Zry+aLkyzilb38kG+gnKNvIazNt+qnqSDDeddcGObHavy3G7qKVrZ
hQxl/f+L7hY3BwRjgbD0RHRPRVVkttA1Nt9+ZOAKQjIfbW+kXc7Vad53/ikPSJZz
m65DCbqTKJEHKpar2biaqHu0hf9S9yEPGAuzFS9EcxLe4qNEKcXHtBAMCZb2+KZd
ktc9ihtgBRORFQq2ZjYHlgtyCem8W51XssPBTLNVdCiXj22WcaD1Ewy2IlvxYDVp
z+9vMy2K2DI/sOr7oPPpQZMhE07D7cLSSH1YAXJUZkvgaKWWxQ7rGGczcqP2zmCQ
WSc2p6dOOUTFOG1UC2rEiU0rzk0GDsH9bfmFnokH3tiCx1EUoMquiF524P7kCycD
TWmCu7EobstrxxJuPw5TM+8faKbYmGlyi/pXogToysp3meX71JlS2bgibf1KFEDJ
QlLmK7sP1YA6snobs+StoWwaZ2fcyebrkJoMm5vrpTHYJMnZJv/JGXFJ646ujExk
Z5BkdDaLUlQDHtqrlKK+G8Z3CVEVbzZxpHIBDF0T7F9z0Y+ez0HW9815NIY1xyxx
Q7ClaxpsGqFxCJFZ7dUljq9QUwcTTFcM+5RVqMvHIdM1ysLY1BjoAk8Acc/fjw9n
0m1Rh4OXNDRanDAE0kMzewCscxJb86GKrLOsNb6a0KucJp4lBAcZzpjDD2USLnvb
a+YpPytRe0H6TKPdbbgj+WXkJCgI8gjZuzoKhoNkiOG4uQsfqnhAqFBM3CfqtWBt
rMTb1OCZgQMJZK9SntQDvGn5Mdzy8gyhfJ35Ch9SEDkOgvZnGjc45+cEfgnF6vqJ
oCt8F/w1AP36UMjkxg/kg9vAOtAhH9qMVAau38MDv64fSx+EY1nnLPz4W4w/7JK0
zWWokgFbExZKHVr1PrhAHbVaUZ37GZg4BRiyVUQ8qZ/3Gn+8+VLJ0+LtLgcbuVpz
7P76Gm9IynZ58jAf8u5mM0pwF/N+SFeNWIYeGU6p0tVsobd1Ga2+ypXRgJR/Mm0b
dU07OgkkKUqq+tkpsAG4NZ2eKsw3UfxwwLz+8jLjOOr3bQMzFwywODjkHq41BmNv
1QyyhbD3LfiqJMLhjikUTnn7AcvpbX7JV1wCqgevDunEOqkIb6ZabitymT5HnGFY
8vYimeT3LFn6FZORgXEsvjYiWsf4M4fmt+l5Kca/i4FtZqQQ0bpovHjXjKT3DDEQ
PrDMslSXTqgpvcjvxToMcIQywTp94oYxx4lalisX26oktnjTloLxpzSLvh7ywku4
CaIXx6eV1+HcDWjA9LoR0ckJuMdQq4AthRhZ98OV5LjzVOk1lsoUAq2nTq+oE7oC
JJfxNPtNqWCWYB0derxpq0vCurIhC5Y687+2Ii0HKYNYaStiS5D3ZNqj7cHCUrIN
6O40xrDRbSbJl93VX31KofBE1gLfwAl/zVMt0e+ZwKXug4QwJVyGBugo4iMB+j8G
KFr3IinuED+NmJTn/erJFkrVZ072OF2wLWdQoE6B6P1yeiEimhMLJE4g0Ta2FZEm
1nDSpBJx0fQFWg1mlHVNwcFLIcz8pHdMmFRLifQn+TZALpqDzxh/5cV3JXYZBUbk
1To0e+jS2jjBFNsIkI1JPwTKJ9QiPDuferVCa0oH0w2t332rTTt7Y3T8ezkTgGOB
jS4TnbM69lRcAS9fx4IehwfaOC3/3qIoldKYujPP5D6QGwNbm/JvNG9ShrRHctiz
zPY6lDUaIjTbw+SeT6jDTDvy6rg+L2TvDt3uglpkUh+HOmkyrdve5LDxe34rAd1B
P7mdllWh5ry1xV0tt88OwSKmt4dop3hTVHS6BrGnEG7lfODHilTHTVvu1bLdJ7GY
7rUwiPLj5gLW6PFgB7yxDh83N5TTDrqmHQtxwllMmkynMbA0bW3Vq8bVc3M3eYFC
OHGHqpt3aiR5D27rycoq4prDae2z1Tylw+5MYhn8puw7DXv2KUoWTLEuTxI/PIjQ
PmrbR0fsXoJxoeBuYlNkin4/g8IzMTp0hMHL3093vV5hZhYDxnVxeNqeXeWwZGeO
odcHf10tgc3EibxKV/LU4FzHpToyYsig38uBsNpDTmPzeufeK9S/bsnKESbg2Fef
i6Zmo1fJZkGltoWtTrg3uR6Wza7cz8wh1829nje/XwZZemek1Jl54RrEBDSDiL1I
x24Smur0QpIVC3eaahN4tj1PG8F7sV8XAyo8HAQae6EnLSvkQLV+AzxYG0sF68K5
Y1svhbJyr+OmYUvDsXXRDgdx1vsVT8pWFHfohJYtKI7JVZIMehqMX/F88IS2b2AT
xXo341n55EwTakSQgl5i+1ILf55OIMZDiZa0G7KCx/RTIJNWBcn0xjItYmx1UgLW
roOiGuuLr6Fp8tsyfDuwclBGeGi8aSjjO8bfeU5XfZjxgoQ/jdicmW8HPBu41RPk
EQJNx8/7HcUC78mZDX7JeZdR+K13c2wZsMor3AqGF6f6h4VR60pFvkUVgO2zRAf8
DDWEvGv6Y5KgsVddyqeLOn08OsMvDgXKEc2oifQLT1O3+nHdJMpgMXh0pPsASTdG
ei0o4HfrG6Ee/rhHYhUqL61B+lVjqteCDjYRs/eapBfBdA9ML1cJshAodJa+8Ipl
JiO9Pz4nnMCJ3S5E8jdQP4thPYmccZRqM8Z1KJ+Ylrpc1DA+w723IJTGEsG4drKC
UsPjCRiKK4Fn2L6VV5ee0F/YXATUvXmYbxUeGL6ZpyIK5E0GBV2MBdiuQfuOC62K
HFWmb5Py3g7cOJeF7rcpDcpznxN/zIy5Zj58Z/aci1jYRLQx8t6Wkq2z2WNI1vS4
x+H617AY1P1/hRX/eUHWLUAO5ZMhtdpkABTov+XLVRbK29ZYmaLlCVkkGx1pjTXC
JBp/QJUeBfrF3A9f4jhHjKaL7YozPs1koAbuQbfXEN9qa04hX2fTL9nzrZS2xHQ8
bXjedCuB2PHyUw1ubJIViluhX8jqh2xnrkZ/QeQFK1rZyCt92Bj7qI31dsnpo7Sy
jGjqGxLOUbxEYmnukf8Se+kOgK426BNHU+mAn50S25FMhScLIYccSOAOuGHNafkS
JMIKtLuSsRjKr4Wmyk79kYfflf6EiCmTvbiTpS2ZUuZcY0/XXat/xBh211H9/e27
8udxOZFntIilepKgInt4q6VXdcyVStyv7tKENDalnOhkyjfhi2ggc9/d55+OZGKL
0BwjzsssLXZ5JzZRu9IedfybB1+160EskEAYpnewMIr7DAhIp+j1CR2XqzuGAGYC
R+vftPhshTgZuVQsQYXwTz0GDhIMA9XhqiO0FSIZNqzdt4xzIeldJ9Gh+l7L/OqQ
azAh/xSzkw9iumvZWH8nnUhbI3nO2D9ouu9B9LJCTvbtButbIeO+BQKMPwXUVwQQ
IIlDoZvH0YuJiBfgrEx5Nv90n4Ure/SCYOb//8TyA1gcoS3elsOXc604D2z0MPj0
+Gjpk5mijxRZefPxMJz0GhR9dHzUOpc0JZsADDZpyFFbayJgOF7HAgQiuc599p4l
QVynOv3BrorvmZtftJcnzRdYeI2WBrflq+fttKUKWBfeV33hLPt3WRzpxqiz1ZMN
skiVLCNbTcxcf/D8sV2r2+I295ZUGgyBEiaXEcKp7YFkBbR6egvKxMNId04oEYyM
xAgQwBeWe27EuD2pVitErMUmhc5twa7YusEiFxX/0PHZ7LORe8+L99nJBoS/I9jC
9GfSpmPAzkXtM2QH1V1CV8hdzTFuJrU8EsHEP+pkjjXCxR1nX7GiYv+q0BE4rj3o
Kqq5WNS+Z4UahUV7Q94iP17vAaCUhyipylEDxuKhxNeONmLEae7hyYiiLY0nbg4N
+/psYBcKdCFDg+flvGsvlw6JQPRSAnOeh5zx038X4z3F2g9l/1w9THxFRlzouR/Y
usDug4fJsMqn1c+zE6xzu7dDhjhUjLrHdE5zFNMPxyxICu5mPgMpLwKs/BmbsWIU
z0z2KvVmajODrjtJjPtKEDjf7L4hOnCbZmuDVJyuFvEIPFKQO9Ksv903eg80tS8w
/JirbgnA4naBklI2bHnzzOj9LcRqqOo7thbnd8meSPDUuMAGGsylY5LpyEnORlmB
o1g8/Iuv8bmEJdbUwBYSyblntLjXVJ52T9nR/0X2yHzze0r0hnD0RmJJMNpHdY9J
cz+fU5zKzCabi2MjTcKS59ia5n7SkP6/TL1qBqHeMZbu8yyg8ZHllQDiCiCWn0wi
vIyY0ORccteh4xiVV+Q+3n4HxiZF1TpQfxcB+J/dtQjdHDbjb8/zT4SH9HYlfl0w
zGFjYPINi/2HS5zdDybMjnJj+Zd1dO/L4baXocTW9pwrqFzIMYp1+tz82C9LJgAt
fkx2nRfoFeHp+lkFGPP6IbCeV7oPP7UkID2PcEaMohYZcQw3N+CcyUWw0WKZA5T7
ZlamnEwZQnFOkcZqzeZYL1xTjjLhOfiwJ3La4hWxlpRT6dJeDqiiPIvtR7NtUL1l
lpeEoCeO0nZh7EYvb4lebYI1xcmcrmj1X8hljyvHf+ms7vzLRP0FQpaIxzW5R/ze
sVMxTskvfl2/2bQkpW0EOXOWwxH0/dxpHcKcdn6NEnUL4iibOJzUdkz+NdGd+vRj
+We9RBrD28qlTNCyz3AKeNnUC7ei+H58qgR8eAjKR2sWjtni3Us2smk/WStS+RU3
Vxfb7u+rfNsSZYOdReUnUQK8AYbaH9AJPfcwlssLVLj6gZ+ohvosORyYwdS/jAXA
27DcSrSKd/ZM7D8pp+WE26s5Iue1S1uqJk5GRV6bR8+Hp0sM6N1i0KH03qcEShUo
vMpRmvP1pbCTU1Jn3wZjo+w+mrmWx7e07UmizC133ONTAAaw46ZH12emQ7MZT/xb
nAxBMQm/zD4Cc2kDnwgV0pSZSuok0mVWih/zpmKAn2HWtX1qp+eoFkc+edIhmKl8
6SanFNaoRW+INsFKU7Lum1CgSwxnOXA0TDr1VrLhpJYrCxpXdJXDzBTi22KTCxws
bApYN4Gu4+8aAJK9EmpPguTuAS7Oy7aC9Y+HPa84Ue10Mo4QKMEbIeK0WyiIWU+/
6vDHbipYplRrRyYTOUpjVZEyWqe+g+wG0YdOnZheE7zNWRKhgAV3wH1xy+Sxw1ce
wb9RRtc/9phmXsuoqboiFi4EhZraZqDW83NNTBZTnjVKZ4x/yf/U8K/Pv9YZn+13
hUps/ReckDFCZW1GzT+y1bWnx4wwNN+wWsO1tazRyJGoJq7FvKTOyeIHcAlrxoFx
07F3MmYf66x9YOs/+9FG+xx2KO9wl8mbMXlM6xJd+KFccNhPS+6HIzgFcC9ZhgCx
s8E3cBUVwTnGfVVX2esqf7/GPoGjurAzXp7T+LA2fh9NAZ9fYLJLCxJHKoWuX1G5
PpK9B/78jkMKB89zkM6o8hDaPi10RWl4CrdVHEt2oVoDCqhwrMhxoOkYmEr5MJI+
Tid7R6KmN0zdW+3QAdmPDzeu/wb27zPN+JbK7u2HjFiKi7V7Ef84qTZp3IKBF5St
7RvY+Kq4SvvevNKqXRwnjDyfarU3NN4Hpc4jnqB+FW7UpAvJJILPdfuTioAsB1qy
goRVZb8ejhdiDooFJNDLxB0GOxoh7jjfZiWIoVC7VPXAQydwelyS+gdR1xKZuE9y
016h5EAnGvIV/Bauf7Wa7yJiqlqJZ6ViMTEHsvEOc77rA49XuvhSq9NbOz8jqxAB
Am1Q09LbuC/ps6ov/fzBSaKFjRrdjf4IytXZJHCzBiGvZiX1Y+OIka2OXMMD09gR
TWv9hWe2Jw2AEDMdc4ZtLkNYQ4XkwGTLID35klDfNpLMF6oRNZKyS4t0jcd+hK/i
rkVCAjzQtLTJjBY4YaGa1UE39CpghIkQiOS8nGL2+F04jw/FCixRgnsCJf3GX2H/
mD6oMdrNF8TLs5HbDz5Io6WEXraTD6pSd30B1q0QftOtmzO8NZAjylfX7YgcXbwn
LDvJUVBoL/AdcrKumxXk/zj7QQoxSjgejcVFez4QXUg5YUUF+ZkynIDPofChMiu0
QDAhOoNd1JivUApaC/7Wepq3eqIOjWWEVAyT3Nc+uoPMYhlzkBsRui2uXvEaGDgJ
ANjocgN/W1x115uKWXhFfeSehh/pWOko2w5N/hNRApaJbx9BFjSgwgebwJHZUdHz
HLJEkeoiHs+aKMK0zwRU3pTqZ9MPwjoZmt/5Om2Mz54YTXWtdhBVxDR7q9CFXQpG
PO3Ii7xybWqC6xIsUhEU4lazSucD5TCWqpzl9i2kUoffpehzGCMU8dGA3lphhGpf
fEKU3QHBmW3LKCt+nnGrvwoHgf9fY45u8I5vD2Y1B6+uK0HosCkbcYHYlDRu7fmc
MyuSNWB1o1md3MY9D5z3CSBwx7Ja5XO6PbP0WR5Rsg4PNV2ao9gS0GPsbi93/87M
qNhiwfN5mCeOABGuQ6IAzifdUPD2krvgYbfLDIA6EYzeCQmZBuHdnw7zejqL5n9w
cALxyNQCQaouIohAFbXgAKIj5Bw9M8eYwL58qlVBt6j/kezqL/SkjGtspg/hjmG5
/5GOBTmOT0LQKmICezrWsTbbxlJLH0wRF3TgNBtHL+4lpIl+5MoKTJQv+SGAruM2
hdVk5jjhznKlD6x3s3A/x9v8/pqy7ae2trCFT6K9+tIDVTRhTeuLkHWce62XtRa3
Cnzz1kvdt5FnIsLoOBmZ6rKHL0yC6fuLMhB6vP3vkFfdgNseuYMadkyM5f1P4F44
RhA3XQbsSJXa5r/5J1P5/+r3V1ddyz1S73n8WjpiCHr4mhlMcofX2QC8DkIV0VC/
vo24RFSPlzHs1fsmjJ3wFPJ9DkUCgpK4h7fuSsl013WRZwYzRLETSLtUxuiI/gS4
gTVxK6CV2Icgb2IpkufR2RYRxZZI6qiuqE92IVtzbBArK75UZ8NEnsmkXOirzc4Y
5WHXJNAjS47jYLGS++mGccHiGHK43LKQVnfaG+1hHWJ6XetkPtJvp7LKMBDigWo5
AIHWZPmFdBtJxFKwOuj6k6exToRWOvzDyO2XExffeErgamoZ43EV3kGsp+vLik2X
P24tMdMXWHdkfHwlv5Ydm8fXoZ7/VQkyBMUbH2kDDSTKU/apAKMc69zF7V9KRPll
QKcpj/BtCZ47LdL1o4EPWnMoEAjLfPp7f/YXJtYLHIvzuvPkFYqJrO0RStR4i+fo
JK2ppqcjKGzlJCWhIToSrcT1tHJykK1YNW6FCCE9KTtFtd7AlRZI8PF71CHyKCyl
jYNK9wCjM19wRaFRapD7BpRb/+T8OvwcXK3Cf/U438rliLqVjUAaqewOx5i3N9Sp
QOadFvKEcoh0YbZwyBZvD72o10OBlhK7/XqkKMcaiCf3mJN/h7ldCrIqIUJkiBN8
EdoVgcrYkO/ECCjJ1/7YikQ5rarfdFr7LIbrOwfdsQ23W3PNJgPBFAntp16wEZLN
JoWLuSleUB1IuHUmTJce6VLRcPb8JM/tH4gU23En0r1ytWK+d3mxqjf51yxrTJJX
+7GmCaitA3w5C131r8AaxUfL7vfUbYrDkVDUdVr21+JtUj9ihm4PkMftRM4UZkKo
rcmVN5ucYzwYGSYzrrb9o8cVJOxEdMLbtd15vf2iVh2+a+FG8xvHLX3G5KLpPX0f
9a79RV+j+ND3yeBX57eMJQEYFEkurHI4xUOfGzSZlph1IFso2MdE7ANotK2vOUr+
RQodRWsTkPbP13gHuiVDvp0RFzqw85tLEcqI+J7IWpEP8YGrYVE9UWc2mq+MCNH7
r5sr/nb+k9/d8RizfbPMGXYgHSMZ+50ERSgc02aN1l6FYuHYuzm6RHas3dlZovXA
qFH+IO0ZrWl867aUZMbkivEAeJv305oDXAoQ5qOo//kHaEMda82kp4VTh9iOH5Jm
2pP7k+ERusSpJbCYyCRGSTMi73yZvlaBdED9n4cmu8Z7xFGYNfNfy6oqvQUfkHlT
mZujO0QdQ48zrToBu6WRnhfwyl2UMf8QwUAr+fOdjE57/D64QuKLPGtYk7qX/7dt
4z7fST777Z8TnwH1OLhOjU24WCczgQh8tD57bR2YqRBgGzGEVA5040N4ZC+g/ruL
CI/6KvjVb5e/VW1YOfOJ3Kg4L1sA/pdufIG+INuLFXdJgGhZL7iNLNkuJmZZ9o92
qVBtUbX9vak70Qk19k7+msBOBGYv0zCh5UKq6ZUeKSgK3Jp/aMlhDoOHfo0NSPGi
OECFe1M6hDnoYB7W8yoqRWR6i2VL6nu3VofoYiRvBlGIqo8doCqkL/Il02HiEFUr
vM7GrsGmOtVngCx0PswpXMdcTDWcEIZtwW64ICGZ3H2nSTevIzSANjQt/cn0S+bd
uJ0VM4+NmCN/dYLC2+LPmyXO4U8AxSe2X58FNgcF/1VaYNpSmRsDlF6zNxn6VkQo
AD+s2ClahR7TZ8yzBsrGq1F9qQhlVH3Gas9WyJKuqafcV/b2qCWW5talcDoppryw
asQbFm9H4BRPuilVOgf8bEZIaJlXeopLugavsjfK2sFnzMBX3ZHF8k7E6cH/12yT
w5UWNWcQhLOU9n32IsA67zCi8z2hVQh4mOlDihOOfXxXiKdyf8k1Nqwe7caHvJ4G
nyBubInLlcKoFGCi7MmPXojC26iwxNohUqSfjO78vQOCEnSmIocCyFVrLMbwBh70
ixm+SsD7heYm8Ag8nXuC7mEc22jA6kbPyK7JvdNo1shAP6CrExdxI01Az5AeTjyb
MONYsNTRX58idjEVNdb2RYAJpxowmDR9rbWRUm2BLV26lNIXXRMZcjZkR57Fr1FM
ZM3G8l9J+rQUOhhmd22L0DDwbVCDg3Xq9HQPz2Oi7UVFU6vbW4ZY26D4aL998KW6
ltAtliJGcR+DI4WFHPgwn8BK+EGDApXT1gouxhQIDBQwi3EvrB4XPx58RxF98qpX
iLqmrTzu17xZejFsGyrLbg/uVGa55P7Y6bdGylUOkO0shgqd8HPfIoSPeQQtpFbg
Hq+dNeHzPHlDTiewX1L0Ya6KO+d71LhGh1Ra8cB294c11PLQD5K1DzcFDTFldp9l
/8D0rqcojhmPogrErk/xefejXMFeBSxlNAwP5+DJFfnK1jy3fUncQkRmWTzLC/eM
SezDTGBtljCka9KSQmgj+eCszgdpxuPW2/Fl0xaDL/YgPrxlCfMVI4lHP3kyg/dY
k905YsH82qf0HZ0MPaYVe6y5j9LRBwNcVMvSpHjJWA5k/8r8xuLrwsKPHq7eBG0K
dCSL8zB7FrzSRZZ4ZZbQ/0YWajqEXAryBs85YFTLgkkbYDMiDZ2/55S5q5sBqjtr
9jemkWnlUWi196H/WdKoWwPTr1sGXMEpUwOOhmFB2oPM8s/rqNbCXUb6u/a+b+QY
bCtr/R0RGAhsvE7mYrqH+A8UMnVZiZIijRFpB8aDXyT+Pdvie5ccsJxpV2jK1UV/
3HLsNTGf9N+Eo7gAwySqPx6JplQTIygsEylsnqBOi8yLmDWLMhso0tfLzBJ2tkyU
+bWeuF/gkARhY4aIYXujSAyQ46i0A5BjtzxxdEs7gqrGVpx7MmeZQuCVNW0O1U7k
PWtGbQeFIXICGvmnc+bTDVxdYKNTfd+GF79o+p0Dwd3ePB35qTnCxo3bldMCwBPG
0Kol1J3BIwB128AqL3I404fn9B9GKZxhAqj9HvzfhscjO2p4oYi5XwzY/r6rCSWX
K8m706JKPcEZryMd5imZBFTKdoTkxMiMKhD1ozSbpsGvLIOKH5iimI2FUc/kZTe4
yuJR/qWNe2HvzsrwpJyBgwMvoaZ8zmLiLiI1iiaQ/YK3wxsQtAzf6MxgbTvVE8FT
Ap/7FbC2MY3OhALwPhYjRObn2PEnZ+6YCiNBbWg9tU4i+cM11WIpVfol6a2Wze2G
4qH0fHvHlfp56QRywPXrd3Co4UyVWK7HjUus4/ZRIrxLWoB9jBzBV78rmM/1K5hY
0Ct3AReWQ7NHK3EnC+nxsMoo/0Tto/UpraXVT46vmEwZMgWjDeUo4e5FQzfFvlJV
b/iR5+MUBzitmm27vQMAXdGKi9IKR3GaBrkCUQtHFS9Rc+v7lNmnmeUYLpCqQJKp
mC3zsQ+r4kNNTaBBzrmF3rFBuFqXQ+tg2/uod1cuEai4pJWABSRnYy/VbfXc2uAU
+OKqrSo3wSosmo8UE7MOInNp4z3Y6P/NL8uYUFDgzTO62Nng2hipwYNBuN0eK/Fo
5dt1P/mgOFhfICM97cXEAyD+AwteYcXZVUc1DRuk9z3q2F5uRaF9ewNFBJcf1xPV
J1a7fUsztn8Lnq+Jnx4Kj3Z2gkDoEjnBahYyYRwvKyPNDQpkEHrLsQmf7ez3wiIi
vUlu4fGduyfDjqqCdtHRlwYfE710hhhBuv1NOCyFJYJzloXVEbWJ/r75CsOMYTfR
F/oOCuHhzpmxmvANrqmc7MnFAg9sO7h0qHl0tDPAAD1sm0uV0FxogLpUqfM381Nv
axPGyEfqAg3atzXIKxMaRH/5gi4wa97eFa/0HpKl606OlJhz+W+eanjwdWg4l0ME
c6+ey1iLz6YT5zoNspSmbm/hJ4GC4oP4aOc262uQMfmM9QWpWTxOCoQvGCPtAfhu
F48gOtgNB9F5cxyQyjSVHbVTODalIwDXVxaFWEjz10eHFnEXkNvMxQChrqXNw2iI
dkVDDelT4K+L2ASS70FWzlA5oDHy1/X6lvZ2QGo0AouS6uYRYeenvRITYM3mWeVp
tuuH5kjuXotnaWZMEYf2DVe/Pxfftx/i0s3Z2enIDvs2xDAherS6Re2YosUqOalp
jZFcbUcuZmxoA1MGk11r5nd1m88xWcC42Xreg3ph2hmn0t4s+yEJ3/79RHDVZMZi
6V+9IYVhEc0j6fSrDz77Mnv7BCW/uIMMa4hpl/4IrDja2AMfXjA2k0Bblpacwyt8
PcsSRvADgP3OXv7um3kGAoiyy4hFdo4D+v2Z8nI6EcmtmQLaPbSqWZ/ITEjHXP4D
VC4MDOdHqUcfUOuYbwTKotlD3VzrycV1oY9+aWsf2HwuM3O/L054gPz03w5RpycN
lOIv1DpbgykdzXLxBSPQaRFShrWWkn9g0gB4gMvd/msDeSXw39xuTFU6dAU1gPLS
rKF5M0rKjMGw0FfuE8CXEqFTC2xAs6/1rdEyi/ZepMCM/l5AGRqVlkuwLzcYi9p0
2xOKRzIFbuVxVyiKqcWHX5AW2SqdRyT6Wt8VwJMLeZDrEYrrJewHg7FO3eYAZyPB
pQwuGHNqWdst4813cI4o3St6+P7EyUsZb3uf8iYcksp2Zd9RY8VuyxEr2eoVfbya
cW78LrclH9RefaOA3wETNaCgjmY1pdV0/4i26U8C8UzaMkEJMlXUo+w83ptr9az/
rw/XSSjl+kXk4ohMybZBOUd0GdKW+cmt4kKJVxesn4YTCkXuuy5j/Gi8mRl+t9AY
Da9fm0oGZkjOgsjh/Bn6XYCAl6yNcAzDEXmFVKbMqSu2HiGoBMaiD/g97ODZBId2
MfT2elqqVkDlkPOuUdCHJGkA6Eeh2sw6y95bRVMsLo9O0m0+KOvFb9a2QP4QjuzW
yoer46vMW4a6gQ8ij/fCwT8bkWyU2VufzLQg7hAK8I2KQ+12E/nH4Qx09mUKaZZo
DQgjpVU/MP51Il506fW0jJY5ws91YOMOjvFG0F6v4kgZwnUNASIPu1jFmcscITFd
oGOINtLuL9oDN4HvIyLKiilU/9CBMWh1z9h9k71sl4UiL9CpDAXnSZYMbi2ItWUR
tEloDtsPdKmuvu11740tVN4qZR74h7+MwYZOcoI2pQbaWHGVMLzABbciwGZnEuNu
8NqyZQdQeLXcS54nDcbCFsP2d5+4/p4c7uE4e3M6fWYMkxoy/9XPSkQ+FpXrmRGy
Ei7Le7RDCOzHXaumARlRc/bQGmuWGDmnBliEkEeQiE1mvaZPuLLM58Hryyx1Gl3Z
+QWOhcAq7jZsRhbV9t2wjXxSDgrvB07lQ+big5i0ggZmB9a0RzhAqTW3vzQhhfpj
0FOkZb5r5xk0tGHIeg7kxgFo+P/rbG3ys54dXfoM2b2n22xED/QDqybLsVDnpps1
SCNSvFm+lO7GDTQ4fufrICMp1LE+iFzhh46vq3JcW2Ej5ya+Fwi4ol7qkJPJne1w
QyJZczVuUIgvGE+UTIRzpgG/o5HK2AHGuaTCDxQpZ0EwEeveVyaP3WzAX+NRH4Ed
Lw8YB66oRX/jWuvqgwN+QXPjIpKFS34QUOh+uyS9mgWtaUg2q3VUc1R+kLDZIaAJ
cWAEdL7WV+h6lL1p++m6CWxE9qPqdDjJzi+faq9ytgfav9TjtaYcWrYMDVhQSAR1
EQAGwC6v/iz4YzE03YzBucQFTE/8fzNuC5ufWqrrtpe4CY4ESZhlHIYB7pjZHGZq
U2bEz9lNrhq3IiV4LET5tExl7Jk8wbToBprYgDxexyevA092ofQKxy6URELLbzpS
iFjbuyJ19dxAVjd2shUX7cx948fl5buty+ZG8XF40pSSl51NHW0S6AArqlAXv9ES
e6PMONwzLUqWKOyKitaVk2dAOnX7WPBMmqS+hg6SdNb6l/ejwoN0Ljyp5TBueGE3
zMefRbuvtX1jKZLQUeD/6EXCqBbaEyMsS73Ou2gXudKB5dISXEJUBWWddKo8gP9s
Ugt2i0hp5ASarktStLugUCHWLuXLa6zYMnu883gNX146Vw65WICk4SYgjknxz/sr
KFuZbRGtAlar0gz2d0vBrD5IacJntNZiONbALyiZoZSzQgX1Qsk4MGZlyHbcK45f
vhEEaTPUs2hYH36FBcc1dT01/i3yTGErgQ45ORnkw4ftSts+fL4K2mzoheSp4uU+
2xZve3TaSVilHgh0OApkAv3l6kYydFazvljy/KPkWrtlyxdyoqcQsV1tZ2K7UNra
4CMH9A0Hslj7QJ9eP53UWIuNQOT3sBIto2kT4Xp2o1qYfpZVVb4AkDkBDlnC0Grr
ehoLLpwGPZ0E3lp3bxgRGi8Sxr0hBeX0czRA8TgU7kb+IsbZq+FS4h54kqtM7SpA
oY4MiisqnxticpveW6XS7kugG8KIwyS1NPLcQiRFZDaomkTNNS+Y4ztWZz/NGZSJ
ZxAhNlr3J46n5oITnSESlyMfm/N2UDl87zVKTLYQbq2VevVMDBI4ZlpwVYXQEkwX
lzRE3TFYmbp0kMgFf2DLB/42uCJtLu9h+jeJpiLbX5GXRNbJTvOkvbQWbWxl0ZpZ
AYxY3yw0EY1t+yQqDED0re/kj665VrT8LqZonm3X6kK9GEfV3tVMAM7sl9ORjhZj
lbxQtrqZx7hVpF3For6oH0kFTS5K55qOLMe2hj46/GHSBzFl3t8HxyzLhOy1Iaa7
MVbEQXut4lpZGyP2seSqclhq+9B3Kfap0uSzpjbkWisH2f58PlTtglfpo+kybLRN
REtQZwtvfWGb7YIsQgHxQp7Pg7f6wJ0mA2OU7rTAqA8q3cLEFL9fNhizamccELxO
Bk1K3USBINuUt2kiuXbnqJCbliXVn1CCMkbO4r9oRFtgg+eyReruZ8mGGASg8Z0v
SintZ/xRh63C9DVRncMCone8yvbEJUjXmZPeKPDqbF/3fUmQDXDK9zfN08o2Ivux
IsWFkrsYqiVC6bi1oCRmG2P7cLNY7aOE6NR75XBt/gXdw1Sv8kKgfx1FG+VRP3FQ
KmnLPWI3rLv8ummp2VMKnCiU6snelY4B8xQ4d11xE6OfYXeM8CQ9FcmWwCBUrPFn
vnutz0gSZEQ/UvMFd0S6oeXnmam79DqBFCuRQiK2fG+a/+4NkFv6KSQbxxSQesKy
5CUdQQU0R4cm3mHYfMA9H7AkW+ZKhKM93On7+KHimDuwUvNaZfUUgFP9iZO4E7g6
E1NZm1JpzWC6aZkktfxOyAZGnNxpmmdJ9mwz2lw+9tdYMBZ6aqVt7HcdJ7DLuM5h
rKpWxU/XblLBPiMhVCkcqxKyLsc6hZvm+BY+E1IpFStXccBktjSQKspljiraz3BZ
aZSv8UzCzWwr00hmjtouLpoHNGPGjWQ6Rrknne7G78pMiebkAC0wi2fbunqukMWY
qzR852zYN5AeHHkR5n+8apfuMB+KnHKFULuiCfx0ALtIte7g2GT18Inx+wC4NFwJ
GicUaKwUGzIp7Jj4fsszXkmMwyc3YC1kT5gma0sTR8avU8oDUivH5EQYh2VRUuxI
eHRdQBEarnS4gkkH7oQwXl50hUz5bhexi9RkGQu73anHS5S5bmiHqIWYwC5Wes1a
IyGWhycQE4JRIAuGqLJwklCLHQqqzWPCHvrTi1DqaocKvIINu2gU9w/qmV7i0Fhf
cDX5qLKVtQQMaJs8dTUnXE9F242vOSsTKCBNifIrQiRCm14QR/MJMqODCqi3/3/1
deA/lTyDcVds7kfvHcmh8g/nymtwvJ2+E2JToK5pbZF12S0g7W+0VFlTGsDjo9I0
CHDL9olJTpr7xL1SLXitZC6UrU7cEldMDs5+/7yRbKBtdq/4hfTrvm6lhddwUA6d
h9A62zAxvNaR5+6Gc9AF8ETOLy7hQ5cRsbYJPxux1fn92TJvAT/26Zrum/SicWEI
V90eJwIB4hdUfFfCs81I7Mm8XZlwCB1yPOn3jSLaahrGSZMya7tN7T+yvx7E/Z0e
wTkTXBb4x3KhDCSCuaAk5qDTj16o6q/VUZpyJqte453XdnHYXMdS9lXrdPSxs9wg
5iUPYyVw4tCJZfH3OPo49TEBD3uNjHjMhEIsE1c4U5D4q553nZsc+cPg6ULHHMuy
D3mrcphMhxu8c9PrCdUNQlBWjZ1znZ8eZqhin1hmfdhyVL+opkn7y+zNehvXmw1o
6KaUB0uJRX2cg3uIHM9ctIFPuRNXxY8v9nGtu5xgBR2EP7Rw5cYfghnANO8w9a9S
dq1P8AOr74qI8IgOQ0p4IKCpj+QAlMThIGnJ7PwkuilmBdwMxlPsHo/zIzkgPHNH
q7AE6nuxd0/J8fiwfUud+XY1Nk62pB7v7cB1QtEVz6nkRJWQEu6f+dN5q6OyRoPh
MyWPHtRAmmfWPZNK5Lcn15tmYrNa5pT1ZDRNQ4k/wqkDLcpxmSYrm/+XMaN2rvNN
GDsjp9wuW/vZac7PehhPsblKY3Qsw8uqF520+GizFMOUun5Xv4o5VTvGMPHVFLpz
s8h3BCGvVWyPfXnB+yJgWUFDSTHYc/92ma0dx1AWx+6udoufWOs2fnpB/a3DEHPI
13k15PzFZlPYtGCRMqoHg3ZQuVGVoAGpwBYNg/bu5+4A9BlPtBEIrWgbfVxck8nN
aOfy6+N7TegDTqdoMc1pJFISOrq6kVyUdUdeDWezSgjVqF+zYVwmMbH7Abvv7vIu
vAVsWUU0Wu+7Qz1yx3KPEmdGztVcWaE8fijicKJZF1axfLF52/uriUn/IfR3dBy5
9/9CCUsKa7v7eRdEGwPzE+GvENMvF4PICfAag4Hu6KmW7d+/JPCZWK5M4lXg1ryH
6j24V/T/D5uGYVcqNVBNxDn8V48mZG4rkVs+/cbiDdY2wUZod588k0hZwOmFn3yq
51Cq60dtwFhiIlYf0w3mrWghtKDXX2tRq55VZqyejqyJ/qJPpRVZd0H7IEIMtZsN
ArVWKX23+lxkmboS1f3fZea3uWC9dzYvrpEvyyo58CPAttm2Qf1N92vnF/lLXwTq
4gvQtvK5S6HLhhyKyXrrQYQQ6xU3qO42//HuvO1JyWDpp4MAfXV6hq7AmNyLbLgj
ksnJhBTS9zGQadZffub+j4OJ2ycxt3NQ0+CsosaElZWwx8IWE5Wp6EqABpqu7PQk
/gJcbTVb/m+J9XviOOpACzw8UO6tmU4BmIUXfeJU6ix2L6Yz+cQO56+n1IcTv7ff
ixQovdBqTLSy/Z0GaK7ZK/ZILgdqjFSRurfIYNS/6lgnF0mgLu2Ug92nIjC+kare
XFAMFIaxjQwFegkwWN0rPSeA0cnAcP2UI3exS1ixNmj+aiCYZFN3hPROV9KccZL6
oi3/KBIvI0P+UYv2GAvQaChBm7f0rERb9F6WzYVFNrfEkfGVfuIZvHAETYWaI+4I
dNNyZw0nH3tgqq1oH7Y3a9gezcjpskROfMFiyN4Jdpdw/+Dfqzl4Me5RCP/ntR3t
ZvOxD+EgvCtOViEG9ykMUJT+ZFMJDEMGbCJHWZj99npsYZTJK7oOOOWmGU7TG1K7
v2C2/uzTCM4PzxgDRX4TPK6LiEfuBD38LgTChQrUt4I4QmMRjhQ+zd3sw5eqB2pT
NiIEBD+vBkxs4ZnoXmV4H3lVUYX7ZMhqxMQwb/dKBgbr6FbScRRDGS2s3hNCUqkQ
YotaXApHeIc7G4fUS4KZGnW1JiOKp+Dqlr96Q2bb+BleOIe8nbgKtKB8zzl9O1sx
A++MO0sg8fCLcIB7gMbRSqCnwDaM9vyHEwKI805RZVxCNZ958t0aJ1SpaMXfNOmj
4cXAS45ZJNmneqvjX5xS0L+oRG57K5+joLzagkPdRnz9/YTQSXfwK1FV5ndhIuqX
MFmFa9sLiTOmVzUEAFM4muMJ7X90W05gVzVl1zLWiB9u2xAXJ1bQc5mUfl3iS8PD
2H/GzyMduohxv+1+p5ameknHxxoUAZ5WRXFkgoHA5Aa3WyRbUmBzzXL4jDKxFLFh
bfJvFkgHieSTKGlOysbLZ7gB6SVrSn+T6Q3iG4hg3FlkGsf6lWrKM7zZaERyAgLG
5SBp1H32Oqzj0mhPYSOEZAHFrpQpOJ7QKZnrN4wrTbWahLclVOpaHTOoXiuWbnAV
pxPvd4uCHh1jQvwEmNMSQ5496ecUqWnr33hGVFsgG8y2Glto1pTF6gqAy1FlqIWG
9irj2fImBlqdB+1JNOeuIQ4s0BSMbKtU/BvumpNwCaq7DUYGZn2K/tjXCcW/fCnm
pHZU0qFe5exYXpvNvugKs0MMNOH3aBOHdYavef3y1qmnCFiM4SnxzX74chlza19E
JYxHKvwWRPC6JNbb1I+QIav7xxlu/x18SuaL7FnPy688MvwQXY7TQP7TyEKWXla9
lRkAjHq8X2afVKkLDPohisqK/oam28g1veuMitdCxgFq5dwFs/He9qjTMKEsVM9U
lv89hYhTGsIgP42CM9BEk7dZF9gvWm17if5IARudwkNLmBQPEXlAxchB5PIFMnzC
XIJA3VeSp0wfTJuipGahMKU4M/RCatNGH+Lmhhtmib3KIwQ0LOybU6k3IPY7g6kU
lDZ1bL3ChjbAm6j4RP0fW20MBCstIHQvBmQyne6l1D0VFWoOlh5Zc+QuttMEjHBz
3rvLlnMr+/N0afK4TKwtdc3r32grFZuTPY32+bMRq3weL4XCQ33vRUJQND72zIyQ
9nGbFYK4oPulfPNdX6e55SZzp3xAdSqfIWbHzyiZO/bPa5Mul/QV+3PU1q4m7Mbl
veBvYeT5Wwb3PblFjB78F5C+HwY355Ndr6QawN0JTuK/NG+o3rR3AMLENXUwLoij
oxBoUOs39FpTjCwi5MzqLzblrBbqIA7pAamskBSyhydtEbmR43CK8wCXhdFAMJy/
1CypIe1IzQhzLqYu7Gdvgj9U0tzw+iJrOvrjZqFHtKUgQ99ZdzDaF9+tTYYHUAaQ
r8XtJ8ng8S1pQn8ZhTWM8kK4uzWSnd238djn7HVw3kNG1LP/fYIYQH/89P3+w1Kz
RDlZcbjrvy6KPjyCqD53vKmh0WrgQw56HMRRaB3vdHtrv4RAqhTnBiJZqH5ppD4B
qVt2yOFcAadz10RxkwgfhX5iLw5GvGdiN1HXj9F9pxuc5l3I0eErFYxkQMWPeTvG
5TrrGjK1/rlnVB5rd8b7HsSlajoS5w5c/wak4+c4Uw20ISM0BwzKOaSPyzBa8IUc
Rtv9TgzATSvyzrUWsYJda2d2nPKugPmfPthPBmQ9O3345xvBnIs1UZu9iIOBGyXu
LVPAQup1257zLBjqu8On1r//vK7VrqViGSZ4ZcM0QRhi5cVxfRu1XVIca5Cbaluc
WNWAHjY1BQZzh2MJdhGmr5b3Zjdp3m+HxNsqvxuBwxdqQqSpVC+7YcknaR3FDda0
NNsgEmurTXTxeLf/33a9pp1HOJGyRqiQV8P2ULJmCwroXhguaRtgJz/J4XvKXiU3
7c11FgKv3sLcdc3vGuYoxC+i3RtRMQkkZRr9phB5Gdm7J5tzeW/PPhkASmYB4+lQ
gnSjmWOQ1y5Rd/7lG3d4kO0KyQIAU2qDaTYuRQLR4fX0ZD14Pb7drEKtvwCjQO/W
dS4y6jKeaxAqv2KJ5sLg86qF5kZkEaEoRUsluyQDT2N7qaic3xDpGLk6zRCnf+nq
jfy/ZsvCnsfa3ocrXuesPQmf4GxMNkK5xt81MQGBzbkv6tdIdOE/if2qqaN7U4U9
R0lgzrf3k2Gu8d6p2jY4z+ZKX/xJrlV6NfF05hjRCk52vtGjww2tTVhkxyLwrQ0h
ArL6Bd2FH/f7ZWVaR4PIY2MW6XRKbFsyZi1ZgDP4rUOJTJBA+Qr08Nlou0PRmZDg
SXprT7KWJuzapICWCtvCY/59bB8LUQc6UualWSivozfv3lOn1EQVug1ntxHQQLLE
DyFh/5IBG7uzpl9mG9DnguYsAt0Rdbd/cjSNTZ7+80t99eQh7VO190GzmMp+R28v
FO6T1751pM6A9MhlfEc8FB2/X0116bk650XOLdLTJXcen5wpOTULN0NkJckPjkQS
pwpeCm8kXrkbTrnDxW3hQbqEByjUxaNoivXMlq5UMnQ2YgwXsaQ6xTlpRhbwLC+r
T66uRprHLjN3oDUa3e7mhinRAj0Ao0PWxdZD3l/P5+m5DGws0F+VPWGu4tC5nI+p
rVPAWerGQOAWoaIr7f5wVhhyO2jk6nj3Yr8Sr1Ci0O6eBybJidiFWovBu1MFjRnZ
Pgaj+tJkQoJbOUd/7AliJz6Y9olERs8v+6T8z6qxyUH+Ebvz8Cu6nYH156d+SJtR
FbXotRKiQyfemzCBF2tUd35F/VOFr3PTD3Bsw7Yk1dtkcuGhjVqHwJuc1z8dK1MX
VD+ozMjCaT7D6yhwPqwNgqpcNZEZgmXFn9nBOiPHklcrmVhVokjnPLRM9OnI8Fns
gfP7XOTbx/nNRJFgPRGARUhMC3mQqGaNG5EU+A+ypMK7tONfTqUCMgZMPr+WmGsV
UpYlzzE1874i3pr0/tsSU0AFYZz50DGsifFTNlx0hiMeUmRxj5tG4ClbTLX0jcPb
3RqFcJ3Aiwj/w0qq84kshN1DrCQivxp/WWlMtgRIISjZrYbp8USJavmk88fa6gea
UuYGplU1K0WvAHGpftaJpzSF0oZmCDap4MvIHV376pkUE7nbPCdh76RupvSh3i2c
s4YSUPo5+5O3rvBnPLW2JnKbT3hsVBzpFVQrVB6Pg/VSSkFqCG+L9+9S1/DgYRom
TqZfeHI94cuBL56DMH5lGcOCbSIyxXhq9YNuJQleJJGK/UUONN6/1W13TlwhmYCf
yyzuKMn9TnbVqsuBvHojcer1p0aUGJZOfDtzArwAZFRc58T5Wo+3+1ADT2RCY/EO
BIQ/SoHFH9LgbtfdKHIPrG45hBy2v7X5T5CGYoG19UKzTwCUzgcSB0q4CjLBBubE
bXSiw7c1TsyzkMyRyRDqXQvMNPSRxJjBIZTmU01eiXj5v/imfe9Kz7bEBhpW1Zyz
M8sGRmXNfDVi0ZSigIQP3tKSo5Q4U0Pd9YBvrMzrdrQZzhNac9F1mG2YGpisqIKK
aqnvcATAdVKVmI5m/F/RFulbLcrjWtU3/kr8fL/c43hrhcnWgGIkakP/imIRFNUf
WR2J8rwuX+rRKjieWOnIQP+VATNHFqQnoj8l3JjaVTZ82tWiw1DkytPQ+v+b3JF2
llNB3C4+nlesbPttfQZ+Va+PEAxsEds/32VzynGdcsQi07GdhlMJNBxzY+kfsIsT
GVwBFX3swb+ijvmzU/9al6OQELEKPshERmyn66136ITB0Dewt5flFuNZyGDSjNtN
zNmTKLArgE+j1UQhotKC83TGY2OoZ6eJYe2KZV6+jxGuC7kuP26/UJ5K90hk49c2
k696Uqr7ClVn3jqUbjDrO24NtdKen6aZdhz58ZWEZo01FhPQ5WbHlKmwlXJTXSLV
gdx/Ju/6fMGGUWC/STe6Wi93pLAuUG+affFK+/nj9FPvZnYRJJyUNL8Kxu7aSS54
3hrILlt7ucia2uNL1uFvBNLB++BdcgFYd6sRihmGuMn6fT65Ajfp4Vz6vCxiXt9V
lD41NeJLQSeIzm8OvHoJCs/QoEe3oLuR76YNT1G6ndzvEiE27kdhixjJhcJRNsC8
qCNrIjN50as+fvOGuFpdStgn3pO9wTmVJqoQBERjxd8sPCDMSAzZEu14otVzrf38
FsBWuiYhsrpDnt5dF6r2cGKMZ9t7FcKvu4+J8X19GzYMLZM1FX9ld7q1mLZZlErH
O+8dTP+cDVHlUDPaIH9UCgbOE7w5tj/2ViQ+fugWPqUvXwnECwxS08JlCnh17vgk
bulhE4rdDy8EfPjxTl+YgxZf8/bWtjPRJaC14jWUd7YwTFoOA6LqaM/buHAarWvi
TjtemUQ/7BDa36BDxmMYpn1FLrOv+GB8S6XBExkjo0K+0zorpYhATxHNMXb+k4Gj
dvr6fJKAx/DVz2wgN7L01L4jHqyCrxufC8YO0kWMmpnRvjgPvAjUf+05vWku0NLY
Njx9G7jL6zVgwM08+qAmJhAps1kBpkHasgd9ir8c17Gl7A0uhoGIUi48Yx/yorZ5
LheuvNSPhypsXYRSkQq2CBq1UjCZaXGf1kLtFrClv6ooLpVnS1IVFWT7cNsWtjuM
j1L9QtOCFOOaEUtlD5cd3sp6lEvGJVDejh1P+j1drRByseyjLQpc+B15C/nI7J5r
sjm/lD2BveGnoLbeWnmvcCf7tYuKpqx6PNPEOEs/kmMIHDxqDiYdww2pYgi0h9FB
1p+pqXdF409/F67zRavPlTGl2I8E/Yj5Fhy9YrRK1sOLMJMmy6snr50EyOxvxeXm
xtr7uJruEd1IWNR86PKgzkghnxs860FJJD06Gl5OhJaFMZ9V3RqR+er4CG3MwUxP
ag/qQxfcnQpb0YC4lzKtPHDZHvEkvBv/zZ1D3j+kWFhm6wrsO2aWHrIp6uP24TIl
j8CRVgIsF/WNqHGhps6wAiCLmpKpIE7Y++4sM5fJjyc7JY/XWiiojlxftogSnBhd
qXguxAxciODrxGaUJsZP/637+vR2hF/kjAE7cx96Hh80Gr9vnqDC20TZc6lSK+DG
T9O9tlt+KoTODQd3bEad9bYJxMp0RzMCKLsPgYI0T4XV6iwGDGPJYNi1WW2E5RCx
ZL3YIW37w5h0zgHn4kDhnrp0RIsazLm8HXskLzcBgFVwUEBcWiNmUv5xhqby5WRN
OEa36rZ3Y0YclWoJtTm7oQSMVYR99ODEumpCAhZ/pU9alLTMrHl9SQJ58rVbwSBk
70YdvG6XNlGsGC0Tl4Zlyoua1STo3F6xrZQl90ZmSeh9qAhy5d6RggLmtAnQTzmY
iQboMOaRuKNeM3hVZHpzwn+SNtHKaVwJ9Ljj590hiM1ydLGWAn6VfNBOZJkLmcSm
B3DAj789+6NAt/AueCNLV1uC9WlUhKYtEj7KC8EaeZFW0LmQr1coIDdTwWut2RRi
qWbv8i2FshfpBVF6T/LsN1adax1c8NlxJu2mM9x13+ejMfnzgvjX1rF5L4mw3vEw
wiBNjQ/KCkpcuk/F9IbWBYCaBg1T/Eooo16dYKEAkAbyf29YNw/9A6V1Ny9nxJlM
fmHZSS3OQ/ZXkoSKQAVMOhzYMToLhoKj3AABx5/Vxx2zb5WtcriZYwJCXJJ4D85M
bYsltRVsQgQTz1/QZ+DbHJhEa0Y1KZ//izf2nAti+XgI5eMXo+JVFom7gWHAvNfV
Xj/E2x2ICc+UXgnNdjAT7w5BciTIrwlyLesr3QBVtGxcA4gUQNv5CD8fT2g+bAb1
CDPCtGnDladXRFbZs1AqMc/RA+5EHFP8NnnjD8+btobOqqrE7oDbau0czX0QN3By
qggVG0YPwD/w7TAySS6/UdGBMeGpGHoS8kI+1HSsvRWEG2bGP32ZIm2lBEmoQhsQ
eQB8iL4v8Doe184TrPshtaJVHmRbhkTkregRDcfxoNw8t8z7zlKibDzhHb94LX2x
ip1clGCd9p+oklUe9YfMN5xo2EXUBH5KaQ+iowdPCv+F9lVoCVy/SDF0WyTQE3Y3
mrPyAEJBqUX2USDaIqtkEfYNCpUsGoxW5YiDPhOwEL1t/Z5EZAVyM18cSgcZJ588
INWo4LFxn7Y9tXGs6BBixnR3k95qX2mngc1d1L6FQIab/kitfb/kTpdOGBfxfShu
Bv1K29+LG1tIo3T7rKaZidFXfB6ZlhUP0vkP3XGthtSZCgL7gdOR4dup5qia3MAE
qNHEwUCiPXIWRZPHURzTcPGsdujLCi8RCp9lOkgssfqBq/ADLp4SU81t9cXXln1C
SBzaOfXOqEjziT919Qe6CWkekMuwRckjix/0O9fYahv5N6oxUQhqZZwbyCjfNH6J
2KZR1zSYgbErBgJUkklg5fHZ1izjZjlYMp1+Q16732wARXxbMagN/B2Pk18sphdt
2M2XCP1TkE4/oArI4TObs6+5rj2mfbRBwEBOdn0NCOu7QR1ixPkYKBVLsv1Cctha
scL0rCVxrq6deXl+lN3u5JwX5O0d2FmYhX4HWOCWU62EgwFRtGfuBmwZs0zqzDNH
BQCBxLKGIhE+jjf9UzSeYRAhTwZZua7PUdBZCyVJ3gYbPgjP+tXDa6xOeJeIwK5B
do7F3kjYgWEemXJn9rn75ENfJNlURMSJv+Ul88ffCSbMzinxM9t10oaQidXX8toE
8xZpND/9OQUMRiaOQvajdEk4dUdDwaagN7cBRp9GORBpJtyZDzUiqHTZb73SSjDg
qqzL+zTQNdTJl1UBh1DSnDi2KGW2HuoTiv+nHfCEjgF8rwsNYFZ/KI0EYkA1U1mV
wzo5o4nXvcKxWOJBm4teKsosLMY8revJFzCtV9+qQIPlGWckp2z5svrOjEFL/pJi
aAl262gTMyiLcXwmJ9lk4ltQLm9A6YM9Q9UF7DakSSR+oXSalOi65x32qQCA6Zvh
PwzRRM5veHFuSVxokQhZtwCnYOh0XDTKt16WzyTxuwSy+PdeNeYJJHb7uwX7EwwC
8w2oa+0+IL6uN+UwgH8C4/wICRssQpBfoeOsiVtdxAaQgkIHjrXpftwhaYdpNs/+
aTRgfc4ypexHCifZPPa0QDvEY/u6Nwa1ZwoCLhs+fmHjJ75o0E/+20so2AheaQet
GEizLa5T0J6L5Qive+05iC2T6boa7QDbrjIUmxsDM3DnC5oM4iSDc+0mLITsx3SA
aSTbyRGIyFnJYS98oqDyu+dstcUri2L4i2R1eCLc50sEwDjf8Y5PXLnF9mGMN32Z
lPz1ID0odJunEMbwQdap8nJ+bv9tZE44oYVCIPB2MRqLyjkeJLKVpdmyFtgyGyJD
iimsyLqPU84dYUtDdbrFRK2N5U6A8ObT4jH0Xf7K4DLd/BS5WAyJ+ZqN49ynWfLM
aJD1Wl5fUfCitFyTIMFQXiFxuDgiaLOyzYM6Dm4wpE7gyq5C40J/kxbbyrL18/9I
+KOYW1iccSSo8OTC/tEztinhtdqsmrp+icDbCRQpI0gy01obBM3PmBqNAi6VG2yn
9nX3S8Hxh7ZFAEE6uwwsFWh3A1zZcRqN6It19tFUv3XT66eszzPUqv/1NKcnaZOR
9SB5RCbwOMu/QI0KFAEVULDf+U6fu3gWLBT2B7HHbyAt65i3bdfODSfMdpIwsZPM
Oz0gO3TR9XgwEe4B9a4aO94h4V/FXfkc1/eKIi1/A9BMSDz7hpC39rJum+8D1I8Y
TCQ5aHWCyMEoGIH9cPJ754pTTcharIzIHIP4QaH2jBgWdM5sXuvCVB78VkEYXFOW
sfXaL2GWx0eDE6owKQJxYSkNBJcRXGWeZNkVNkVXgrgrx+cl5H9MnhABoHME/UMO
+Jz2eCSkjdlxwSL7l4mAks2FyY2pDFInNZcEtHEmeNw2LIBexb7yqaYk4WUYfaRI
c31UTXSOAkIBdA9eJS4eXshxSg8Mc0A3A6pW9Ru5k4O/iNMqjhKT/BO3I+TodXCj
Fg7embfLoTsKK6kJD0eTPs0rhJM18/3DIdPpNP0UEVhLakVrA+BHLPWe/+9BWHhC
ZVm+HqjV4riGlF0g9tQwQ57qlCQrQ3r+Ks7to3aYd8qTYiVQEu9d+LKFOQOpdC6A
SaabdQ3+p+G4hvKOz8rkNdEYlN3JKaQOw09dnu5IRZFlWM6AFQFQkFgLHMmL65c8
k6tmoSQ6lyIiIwATw5GRoHKXuphUTTskxTkveCUWoEvSnkG6mqI3r1OcgSL4pzME
1hNZa0K7xPD7JPg+9Y3haMmhkXx1b0gAUqYKGt2L1vM5jT7rzVZ5JWubmKBrU8AK
QLKVdSWw17m7S1pcyEI3IUvaiOY/ND9F5l69+/6fNAfKz9A7yV7/4x9ltHvicrgp
JeBBASXNqgM8qziCVwUladA8PZK77Gcin+t52l2wRY6V0JVcXM6VCGQ4uSZ6rHGf
b0i+mBBMzvjr/xbG/wsPbzTrjL0s2yWtkn5+68UQOFcBTK6w8Qx7yCPalbhOuNb2
yoic1abTbt3Lx8prFOXVSimE2jmmfr+qosb+ornKbxD8aS9p2NrbHd94BWsgvmdD
dluj/vt1gVJHkFGZ9fPCE4RYSESpQAFa4hudrx5SUcJR1oYZ89IuhW9zqFZ5rntC
V4o6DFnKAXlsAwiITyR/gx2msUBrM7WagHhIXz9HLxI+2D/hRNBHRIzoH7rMVg8Y
9GjLu3zlknK9tWQLF0YhIyvIG0eeJVRz+7aGslBU9yiPzuBkj28ZogkFPMcoox8b
Ji3Vn1dHbqexQgC2RSG2Z8hmZhCy+KlhfXXtvzo/rRVcLbRcr79RwQMqEYpp3LGG
ybBBUJDgbpQ4XhSH6mySdiPVE2t2aglpmKw97IJBJtHTzmxghgwWPkF4SHQVn2bZ
1UOVBaUcJ/OOVD+J88WhdfEDqaQvsBXAEEwcrIqfMavOuIsW8zhK0J8h4BKVWNqR
wQsh/3nUleP07I35fEvWFWb2kfT8fqjI0mPKduwlmYjTwil0Xzvhkyo3yvye4/uo
CRhan89Fwbe8yva1Itqw9xmUyQk6s/wxZ6983mMVoXLBiUl325Q2EzL5vnD+pzPO
COWNUisRtY0iP/FoBw0kgKNHpKz+h9Xk4q7zAIbtnruCsatzE7uvg/8aGV9AVQnl
oewOiRFEs/nTIPdY+SfEsucrCngBbNsORGQYA7KoNw0unrDKJ4e0pFH8USmEkNNs
7gIGbh9UlsDj4DsqX0XK24MKTsJYibkfuf/7noViZjppNTCnsQNewmGkNOcJ3r/+
SXsq+hTxkkLv9+FgqeFY+oeGFSwREdFfsG4bJ8pI8Cki8+wMAursV1pbK9I0S+87
dL6eej4uV7epAQGXWd7JI7IUZHYjqgzcjO/X3NHwZttAW6v5gp7h4qqUZ49g1kdI
pkl1Y+qMeC0YsL28WBDtTnAtS78nYCcL2lysWfG4mbPEO7e+kL3usbj42jVT98NX
SDAJ1X80qmjQlDv8ruH6jkLE4mDbRV+ysO76YjwrqugnEX1x/LFZTXvpq7Hd7FF5
Np7Pp4mHMHK3NxdN2qzWIq2kvQNI5xa2uE2pg2YC5xI24Q6CABmluyYdvNjji8nq
96puJ5eFe633xs0gx+cdrrTk3ESlUgY2xxmok1iroHBkfuQqpNqok6USayFyYrfY
KgbpFiYPe4ZVX8xEDPi6/xf/FJKYqYOcR6WmstD54gnPcHyMTKl1b6Q/IvWd5tKi
Bm2AnAZ9CQfLApQv623vD2xqvITu/tzC2+srwouoFMP86qli3jyrLs7cqcwyJdGO
dt0pfOaKzTMTCe23wbyejt1rxIp0Sia5JtJDvAZ14M4arz5iRUPCOGuDbQqCXmX5
fPn5/jgRusLtp0Q5/+7VlubX8rz1VnteWAigbZ/5lKpra3zlxh/onLJcJiharcSZ
TzMbCrCN0Jgb60DxbZ3yA/iKegxHNU+0+EfYzNL2AizLEqRQd1kEkoRksGxTgF0F
csL/z5FaVJg6YovaZWN+SJITQQ2gkj3HwmbK62YBMHWzIUv91wDBPatrK4TjXsci
uiqR6dwtj2UlIniUh6FqvIcrI5ehTbbwuvluEtNe4p3q1GFJiexU7Bs4/sZaNV8b
MaMXJjI5Xsq2s7T8+fMqwK+V3SEviyymVM6poTHEipe1CrG4KyS4beJSt3MMKm+6
2Pp3ov3cSURvI0vcxhZ828yZv6RZDI+3Yoo90K2D6zlpDkMWlo3zLzw+0nR+cClN
m1YYUFeu7GYvh30EVokBJAYLvn/KtP4K8vVidJZTGa5tXlWys4hkVLMTxer5iLxJ
JuB36QG0gm+xUW/yBg1la4wFFTi0oGUQ0DgsGSZOdL9YEeGIN4vuaq3lWHKJKYnV
YsRNKBtDSz+FEHaDq4EYK61zZ21J8qgk0M2mtQBvZhwNoyGvFVVpLolOOxQGps7S
8uGH8EClcCG7BVOo7YVzxzCkmD9HnMNkucnQyRThvMu56rTBBAf6PYJfunJzNXs3
ynFddCWEHYfTEABxW71xARepYI3m60JMexrGc0Uac4tqZp825uqFl2avBsb1woLr
bfr6ZgYlVobD1M0xg9uBTo+nfETlMW4r13LNAuYEQjtoVrIIM2Il52gdpRDj5+u2
YOKwQrm1/AyjXXzqOIsIwZsnFdGXrQIbtHITAF9A0t/zVQt5kZ9iwZmEljQf0mZw
0YY2i9EhKL1v1IFwKEPgEoW0L+JVeCbgUgHnJDxnwJk/iU+UupV1p04wUFqBXRMN
k8HggC6tstTsoK44eJB2hm+hZ2EoSOgAJHTUrMT8+U9kgCZmfyv6BkhMqBotA6m+
vDcdOzN5QD2q9wRU43ul01fCaPfnDdkj4Ik1nDeKECejAQF8yQFkpiNzrWSsoEUS
j/7uf5ozisItA6zSO2f310KWASVOpV6Q3FY5poS0exRqMg4Bl2lMuTwjrEfItlsy
nWz6RJR19n9H1ObJKRgn2flxwqZ+eOmEaeISzccxqoimeCJa5vgGm99p+v6p1W9V
TxuFFQjj32yqpUXVlilcbgAwFG5zFbyyveB6Oof4nHLSGp1Gu9vi8cXVX6h8XubM
nJQMWesW6pQ1kmaRP2ekRQqe1w9w+yuZh0TzKzsL3hLxt55EE62UkihLwRNSQPMj
VgMfSKCiqyPCRJPAEBZ5sXiqTv0GhfR7y1JHBH0mA++2wDJWC5rtbft8rHd8ej7x
sFpx9VDEnXpKTUsqN8Jr4PS9ZDYy+srB2rA+TaqoF/Lj3MwCnoPlS13595cZnoLK
aQNooQxtw7P8u8s7uMT1P75ZcxvQg3mSu4ty2cFfUZb2Tf913iVaqjc/dcd8LtjG
FSmRLHdE5kVXzC6aa9qgoTzraE/l6Oe/im5eRnIPl0D70gHUv05Mixv+e68Dn34u
l29JV/w2I6BWJAkHLjKTLuThlER2AG3iebal24Byt2sxClHav9FsHSVjCE+Q7frU
lIOKvOfP0SF0Z2YwiSiitBz3B85LQO5XB+3adUJUVCbjLNUFHIc8l3AuFbTD1jti
A0de8deqSTbCLRGj/kibA5wuFRU5fXE+2fLGzCDwrJ1hSbK0PUnnidHiGt+xghtA
o2ywr0NUz63gbQfcDY2QQEmMX7ZIk/yBA1VOSLEud0DQRX/+eykO1vmJpxh5B8B4
vyBh6WSSU8g/XO5JksapjbJKAP3ReRUtyXpABAEiQnk+UCJNJKBpyVnE+hLUjfcb
wyGgVcNfSr2wS1muT7jnxY5eeXhdQ25oTbvdQbhB5zxjy5W+cdJVLyxYFp8kU603
epkQEp2Vny+ywQDQtH8yRZSKBxLGOamgMUvQZ4myvT6DzQh98j8Rat5dh0AOAoXd
75f9Muym4etlVxrbYSDnC4STlfGMCaLJhHQyLQkNs5PxAdUuNIOw+cXF6Q3PguJV
ZOXSOFQJP5Xi37UuAc5X9b13aGoyLcb9BVxmvbxwlXf5ZLFc21eT7wkmJl+sqp/W
MCj0de9BpXIipSfMZiMY4Lc02Meers9G2ZbzgxK+k7aDTpxcxDrqEk/d30TOTvDA
MEihrXmWYVkrw736mui77OVpLU4O7rRPzJF0dXzK8eglb0H+RF2FI/mkG00mEPfQ
fw2gPE3EhbIM5NV4WZ1nW9OKQ0ImtgUtgeor2b0aK2DkHdULbObCzkHyp7Vfv5Sv
fuNaTE1/pBVmtXoktDlCDzq3pQGK3HRQIXRC9YFHr5g4C7C7cVvDg7Qjjkxtl46O
a3n6p+GGHoJkbdTgum4L5U+kn6opyfpeSxLgOR32B3Jqsy8z6FIXDM3+pCiSyBt1
o32XZYrazrXR+8tT9mDU3aYIM/cJ5XjFlxJLseoKSkByAVp3+4yb54xwmZIPGS3s
pHP1UPE0PvZF4ezm8HUyraDeGNl9bXlfzNx4oPb1cNieRaghMl5jHvJquC9BZLy0
okdvy2zEPnf8hN3xzYxArP4vQWlzkHXfTfeJckZ0U3kVfG13x0TeQs/iplrk10vB
BTznEVI+4RAiMC0nFhnDTJ3UIP80OcwjpdfnvksbxK7I3juIrokE7PE5BxafTM+c
mse1f++BngFD0ONWRaS0k0KvjhHT+C4k/nUIQndyuYLd33LlvUHgSjfv54LuT7j+
AaoZiLLj2kTuAry+E7gcgBmiT5yn1uPaOAn7Y5KmBn0N7kNhBn0GmvDARjUQgATH
7Z63Msw0n6EUolznsGwox5lmwLpm8Na5iI3IT5atSGf3queRu6YY8T57ZqHAalag
qnq57HhHgL6/q2FaG5SZ3Wk/nnxwFdo0gB2hzvi70KvukBcJefCqu0fe0gQI+Ad4
NXPG1OKPNg4Ej+iWJ+M3rT3H5kibn5VYoDjClK0b3ko930LjUhN3hu7JxSdK/1OS
Wj2xk4plyrJIz8hkHXxElVZ2hAUw4Wim90ku5eVn3IiB3Od92yASNHa8v6axJc4w
5jq/uMWkcCETNvBHw041b7bWo9ZvmU3kFzbNrTBYQEtTFm/KHJoOCuNTs9mokJFj
ABUzWoiZ4JNHQy2AtM9ps7zkOcMj8SbTNGppfFxWcmSpQGR8pWKwQduBOb3X/sw0
V1kSUYkH7hzVF8SlAHqD3pYtmkxYdkN8diX2CyKQwaLz6t5NIHDJ+778gLwxJ7g3
KQ13uzxPGG2dcE1twZ1QymLzH/9BDKPnkCFuSKCXcfY0eJ1X0rgFv1AgsmpScvgg
pG4NjlKAqndp7WvrQfE8N7xbhQC6OZnpVjrqGl+3ioGU8hGTIc41rd0IbykKUQRZ
gS/pBRH+sbUNI/9Kdb9zuVuBGnPqiu9YT131gxWV7sLq9WIkkGqqL//97fTaW91D
AXBcc9CvglIGNi9UlsBGELiDXXU6rsBKJDpU6DvkhSR71nqmeP3rnBd/xHrNebKx
5yY62qD7jjjKhTpkvi8J/ouWzGzYHHwtGDccQwlbqUmxhoSKlVIK/jnOuUQLkA1T
CNASZb1LazJcsgRg70x1MrehNi+GSBn6BDeIOOcKky+i3uWrj+2vQ7EbZJ75BDh7
dOtsgeaN1Kw1DsBG3wLDeSZrskxcqq3To4l03LRqmyJ4dOhIjIs7hGIr/3B+Ic4H
DYPk8L20q7fkHM4dylQFQUTiyvQ+p9evR6cI974dWqjVMuy9WZsN0K7fwmUCIaPu
RyYWr6vdgCmWFfJvn+vQIIQJNzAIj+sfTheVBf9GibnF6cXcaKPtniMTnhWy3/F2
T2slrBZvHbqp8jl3CEHa1q4UgtsJ0vQ9SX/3NQdO5uMGSf57L2Hn1lJwl1LnBTvc
BBlIpvvZIn0XXTH+oU27EAy2/efC2HAhsalxp9UCFNLc5G5Ehgd3HMXuVWUrjc+4
/mMWDt+gMS8GGA+GOIJf+801RshrblZ7eNepkzokGddIsQDZHGfUwuZLnNFy2lBe
nJ/2OgBTrAzl3K19FvGFAgGxIQOmmYPjxCA3f8Mibg3DSwqx5fSwg0pGQs3/RwiG
bznoGRgdvQ09P1d0StPq5AxXBGnRv/yabYt3+XV4Lh8Ij2AY9+72Q1AcvXdu+Rrm
z9bOWcLJke4f/u7Ph0mkNJupoBf11pG2PYQyof8e5MPTUPmqhxdIPjlHxr8p2lrN
Ac9pAH87AVmjyGKnQaBMc/fR+JD6A7qI1ceDcrMyPOTyEJxbuzwL5XAOxJz7YfuK
bMTyt1X/gPeGIOaKp7/DpBvkj3+oksWx7S5aQV/+Jmis0+4mcQp/s65605L50P9P
FYTGltm/dF1QIfzeRYRgpsAFUzJKf/7ahVOrMZULsz7MAzu54JdiAPqjVqJLyRiA
M5vG6FBaJ2TeA0V0m6Fo1D9dD1oOqiRxP+ejrIbUHen5KZCp+iWPU0E6yOzthoy0
eFZB5wj8YAvWoECnyOQzMVV9ubzk4E9YSqb8Ub/zxrIG/wqFWxPppl04wVorwtS0
juUQS/8X5JtJQa2An+IQQGAMLVxXXZdsRNGj+d1aOakX8HC+O8MKTntDOfKjbGjS
pSD5OelYGwrng3IhqyMUWdXcLWbOFnO7Ll8s6yUl4j3R+uVgKDMkiwuc/6J87uI8
TIAxJWMqO6lmX4BBpBQvRsSswef0vHy3lry753MHyhCF4/1xmHeUS3uF0uiz0soo
VLg2OYWBxDHddH5Y93uAR7CvHjPhTh9/kuUeopL7Bl2MU2EaDOb9vHCL36vRKkaE
aZcGjcfQEZUVG4c+/ahq8TmEPGl/JJnIyEHpLuiNZ2Vruh/boZjwiFi93YPDEwbE
Ddr9rVVPuFXDyQ9BJpI0tW7D0UiLwWLrqGVGWKcbseLVm3bxd36oasKojDuYNLqx
CuA+KnrTKzK8Xq0H/0wslFJXHcBxrNaDTaHqb2LGPROkZgrrjAXNZsUMVHsHj576
K3pcpuMWqffC8jshYiaQY6SAl7vIKZNEupN27p4D39J4Igvnw9eMMK5KMFxp31ak
FhZpUmUF2sVyd6onlrwitLf3H5bh95zDYduwzessMTar/NT1xodVh8r32TvIoYFD
KjJLIqUYEOxL11iQ8Ro8kHFa/9Xio2mhYndRgfpJEBisDRqw5l3Gqj12ub2kxUwB
PMTwUfNMhhf7tvOGPZojof4kwSvEh+GdyFBaCFLGeyLxpdfyEoxwdbVhUr88Avm7
e4V6siMKSHFiP3wePufSybvF39EVoIi8kniqs+1vMujt5Ery+OK5gKwO/iQKhIWg
EJM4EVi8FGj8llS45NiC+SzMtmw73LcwyCY0P8jFCr4UK5kO3pEtxsLozFIwEfFo
bNITAQDgGiFxs5BpddwAlMJnit/vfGp97DGPNlvLVH7zHFbkyaxOKgoqnnSdT+EH
0pKLD0AgUQHljEcn/cA2VWcgtb66MrT6gUK0tw0xlcdBBZmWD06EBThJzEKvQ/QG
lUPtTwymADaNFNYmh2ijt51iLC5L2L4zosfaIzHIo1Rp1/muornam9W1zsfkAld3
7JzJoSvxNqtfZiIZPFfAeHb8Y71SRfKxlyjgUj5cTD6pSby00EpqlLDOXCjQ41OX
ArArVdofBhz7jyrFjaQFDxoz/axcU4ONphVf/NArWPx89WH3aJPc/stoRfuaKPKb
B//e8wM8BryWp5kunHU4bXrETOmhzpnf/OKv1CVoDRJLsJ1G2eh179CivlTaDUaA
f1gpbM4s/ygL15AT/VRMv4EMPvyFBYXxwl2rnWBXvye8wC0m6Bwf8M2bW+oCKee+
+sGmyvIDTwIPC4JGskwKizLqXRkTYu+CBP6Y54CpOKXTTc4lfxQvc00rVfiWECT2
gI19RFwvQUWzwmlUh0Jcc4Ht9k4UsWOV+ROkrThhsKqs++8NB3XYR6sWClVYa/JD
jC8sY/bubsRcOsjlVK9MsXw4MoRAYlpYqK+LEUSemEoNZY3A6u45UUfhwz35AqLb
tpYNV8jZPX6dOzqx6QwdaSArMUcMmPDjXZ2DoyH1HU/Wb1hfHMZbi72jAGKyATX9
9J/MQwEf365KjOOi0MYFACJ3+kVmxWIgrRNTiYHnPrHymsqoINK2EygeRGpcNk6j
XI4AdlvqluCatEXyLMQZRU6X2awez/7hTykgfRz9sm4mbz1QutpbnXC4LMHSG3I6
Uvk3teT7o8XS5OjMZIiHeKq+yl+LXeCUqZVlr+c/vzS32uhy7IUbxvv9LvfYs17+
X6DaphB+Lbd6eHoZENDFX34KMCKpUQFW0hdWQNw3uk6pwgUTzpcALUyxOhcpZzP/
JFyBIwpFvFQ1eZ+HyDJ8EmmsvdwvzHfP3xlNvWjVf91vZ8lPnJwqamGBLA9qYT+b
1YEiDQ6+SHmrTAsM705H0kC6LoWUSR2LPIxh0JQgufW5Bwfs/c7A1MQTgPmQvfzW
norV440t1xzKST8o7YId5kB53gskkS4sj4tXBXXf3tJoQZPW+WxyuNwnGdoC79kL
P7ZskzTHZZivRfPskpZps3Pfb+pd+bb7bsrRftugh7St1QrsBNYO/NF67+hjNjlY
mO26gU/n2TTIRe4mD8BA73yYYaIuCi0LuAe8/pDXiu/TC/bHqBtDAVHv3svAWUg3
b7OmYzKJ+J+jbo8BuxcnlEc/fBV6P07NRgXK211M2zIUdMRa9pd09E4KZNzbW/da
nyiJBQTQ42+JgGN4Ey3v/Ja3YHIUUjuHyiz6BibNituku6wH0juWuuCivjAeDwvy
V/13qD2aH2be2tunceAMkMLdF0B/p8UQVCvS3gzbXWEIpS3HkEz11IFa5/jYJl7z
g+Rin26CNFNpZadLK2tXwfww9YVAVxYSNzz09Sb9nBFJCx745KFHp6b2NlpaVek9
5QR2DONRDU+hdaAeMkbH83nfs7CPRn9+EA20RCoqG7mynNHGxliHY8lAS7eUbwxf
VCPD/DkVgs5Q0OQHSVcfzGgssgCgwx7wP+TzOYJRUwXwrYYHVfGjOcxT+nNgMkRB
o4YQayy9sFnH7XkLbxpvI15MGZWfakjfazotdZNDVEyFOTLeLRtjeDSu+Ds5TZRA
8erlqD6fWyqjHbV8Q0JN2parRrzUGWmz9M7x3SCRKG7wPvZDJBvNOjD6n6rV/iyp
ApaLbGbJAGSoXT+0iezII0nyJl6Hu7PWSaVIOdwS5YnDikXwvhM4lzTCo0QTQAyb
FA9V4y0uWrYOgm0c+S77o/dovBHoHNMyhaNChkqoGWU0Ec1BbHowGZehv84UzFxn
6aVy7WoUhcBBimm1lpHFJ3Gf2HKMEoOarI10SDq5IH/yCS+sFW+5l9kpQPRNWWA0
TNQRWLj10t3zY4VEABehT9Ekwd7scS+vPD+Hpk87a7ANejRh7yDOHkj/aCIYty8h
b6rAlFo1q41r3NgwXXcsd6tjGWA6UGPVpURz+IUkimJLaMi2eyh6lxFT9ouhEp52
6dXqObRgHAv84K1fxkAlEq+dOF866tcWu9w4+/5P8QDpK9K3e2VOiAecZv1vwFn5
fG66cc0PZhliYTIJoQvuZoLz5HZBZHKFagDGbv1zN0389vSnYPThDJmz+WaE3Z7E
ymf4+/R5VKdyoU1gJtn0ZyIMuQyPC8G//9a4qIVrxHPDgOTaSnQ46BbqQge+NFh/
c67Cqj26Xno2jcI38Qk/kv8twNR6rqKxhokX3EAO78NsfTTUlHSXDjqUEO+vpihQ
G5uny55MA2DcB5DrQSjl5Vo/qmP6vw58x5szGD5Qkssx1ajLol3Zb3rxVwukwEQu
Mm7A9Nhfs1Cg8oCetUr6FJbog86r/vVxwS/+W1OQeBpudwJRLQr4XDU8x80mzspV
viQ0ImCUuZ1wnwzz3nGoIj4INIdJBgYj5/q7RYlrEiLXYsXNADjPQ6R7QyMuAQiU
lp3RCLNJAPGN4Kfr7WkywNs7vnjYT08s37//OzD+JK3twwGtG9aFVK4k1y9UEHh8
IzCrU0tmQ9C2qO0gBMtXwzhYPaCWm6YcKJ5nLYiS5Le/oHgKbTwDTWkhO7wf0g01
QybOTS1qH15DgrEtyNEMFVCBWljGncBbbV6fiGZ1yNvnCCzIjabJHw6RiPKABHqB
KgMYhaKu7junqMkC4spL699rdQZVi0/iuC20QUWSLLJ1mG0dQJBejDAk8PMMdBU0
fFCJfuMPtVCQntR404jnev/en5GoYwNQvB6w3JnjHxi/SOlIWOzBosxmrxn0S9o2
6zpAuw8kbDlHGJgG+zG+1SA5q77FXWY2S9Z6UrEhqqdYBSdV//IukZRYHGiQBFjc
t2kKoW6vznSByWncglx9cpHnGJzjjII8sg+YTZ6OGVozPEum815nKUAqUsHJ/bw4
f41BnGfLkT5TJRo2Ut+8Uv56HaCXTg6x2JSqANXCiZ5q2EVnfuFw2Qx8aP6j1dF4
R2zpGp+iOmxsKHshLncfIt6LH65bfwPS9ff3CjyQys10NKSdcq+aAdM0k2A0sLPl
kYoSwVacbmmooGtUgxqGMi3+4ghBdw/7IaSsq5hRo5aaNU+953+JlJbwCUEpR8H7
44DW1abaYfxdPPsFYqeHZXYQ3VwhrZtyynuQ0KTMloKNB3Hz1MuvplF22REzMpui
VEsisFQm+o4F3dBzvOO7heZ3+a5tNzb8RbHkgHq+4I0p4QL37jBlT6NWzwqZ85KA
bm7202Cptpd9QCXVRt40VT00HcZFQ38J8wnI6miCckoJbm08vHpX5RK8qK/NP2Vo
hr7RcFvFqTzegC3K15pUPe0Q9ofnRmOzYniF79MhXaHatRchp51IU06yWdbDKxsr
axM0AmBuuh8NJ/D7HAxPOR3nuFC7NYbZLQkrBrMSVtvz/94oYM9NBCjA4ugtLgjh
uGnMXlsKf35VsJZNZm/tPr9y8PYapG77hF6xme6ZrBkbyolunVB4fqOm8BCgUIgV
371bVAf/1mQfMkOveMcFQYzo3jRBd8J72pH3XeoJyA+v+EBcTjBRCNrldmeIKub4
PzEmXMnPapyZnaqK4PQ5YSiJqvHeYW3P6085imF27sdW9+tb4Sg/qQ4i9jQI3NRK
E+37GCJs0/sLeV33g5ivPK/8xiTXbq1aBdCUIyAvTRNJuzgTLesVRDhdggC4AsnL
1udrLeIYAj4g5hZYkf4kjtJrynlSfmhUrFn9WHfdvCNAhgnzirjCr8PubHuUnAlV
f+8VqqiZuQ+FcqBOlfBhgdJ0kSkyBABdvE2eUFg8UJ5E4/DMY346s/u1wy95oKbM
ulKpLdVm7/dyLEAn9OD7akdMzA1zzaOEBRaZLrJ93qQpO1DdUD6DAAddqD5nD+/N
cOV34Rq/0Jr02EhKtfoe7XEuyLORNztSokCGET5k/ZWiropiBmxYoY5dZxanGD4r
7COEdzTQ/F4LCIlaD1IJowZ4HJYEjPK7QDw805wR21g3PqL62Pe8LGjLjvHJ2mEJ
15rifVa6WsHv1W9ONkvQgVkvf/LcC1wFd5F0UUbve26b/PBImYsoByqNWJjJhSAI
uLXdITw1mLt3vInIUnGlC4dXy6rb3KJs28jQmoi4suEUudth7oLcngu4hf+MjJGc
MgydcSlr20QsG/UaFynUacdlfQtQVYHtFLGi7hzhRaHQSWS8Z/nma0qGD51t/ueg
1EdIjsgppgVSC6hWbQY8uCSb1+Bfm4rAQRdQw4NmTys3PltaDEAPc3mDzuZetBZS
2SPG9NljPtyU69sHiW/8lIWKzCwAMAsPaFBkz2O0vZmwje4VgAtOVlHegsjQXp4k
8Kw14y05o5GdxKz81yKSDSXZg78RZTFfdkEYEmTswNaYBxkeSYcZHvPyIdmW0T1C
JWbWgN8QOcUxgmVWjUkaUWk/4QjID31KXl/rykR/F3O4+8jmgoiq309mLXnJ3Shr
sdlIGCE3dyTWRKaBt+3JAX8JMyD4cyziQvWe1zJQG3om4yRQagFZTBq1KuNC3Srt
DIYcUDXey9px4VNDDVXwC/K8tICSCy835cPHpRmILZoBJ1FisVJQTsdhLTMHX7aC
SS86WCUsVTls7eYmnma3lzFJxUjAdPmJHHvezMuUzr42D9bWv6NlQ1gsyf0cK7hj
3gaBagE7K7eaQHNnFqr6+2RFkMcSd+BeaAknm75NWPMmgvovtc4/lWf5d+fPgEN7
s+phNzrBGwC8V2SJpzz2MbxJgx0q6T6zwN1/xtQZZrdPG64FZw6KFQ2DtryWNsf0
9v27dpsaHK+qcqzK86zb6ey62eVpUmNleFD07G+WbqN3USF4j7uqQuZrXuuYbvT3
Vp4n6Y/b/nKsgVJuZqfSpOXYv4+j+3TO5u1eegjNDRqcwK5WtMMR7USSMwnKZN3T
gj+IKxsHfcZ3tXF3619xlKKrUAr3KWmGZNMmGMcqyLOyTBgX/ScgLNRNLS1GL6aP
ezrCVKU2STBbYoSsrQ7W6gyVxaFXX37nNZbMSppjWuPw/Hi6oU1/u/QskbmtmbNh
TBvpqNuHsl4rWkji2jN/OcLoTwTPyyJFhM7P0IEqubQMS84Mgui++IZh6Ppa7YFc
NiAeh8qfPTIVL7LVctbDRDjNLLu89+1bTiw//RYFj7w1DXTHiKhOcz0Axf9uKBld
/fcFaMRJA43SsizF/+dWKKorfmnsw06tl+ETomLryN9IyxiSjK6LKWJMMCWzZoN8
ZWzArtVRK5aWzJsG+rh/uDzBBBCFwwbpJsiYzQ7lelXTseP+Swu9nObbxqQ6VdpA
vWbcR1ZEl/od8q3RGYPBjBFxOnKxDJlbOvvyG2Rm+WiOPmoxtEmY0/dfvztGMJCH
DYmJ33tY5cBlq9F3afu9p8gUyuIHQb/T/ZMCWqmsTQIk5TZzTGyjbU02quBuCHYp
VQpNwu/ttTRd1nF6+wLex0evB+g5HzHcX4YlqPnksZuPqfM0SrLyeStGF9j2vCbF
+9SyC1zaCwGefPGITl4DUBqrPuir2p2F9UP6r7z8CXsfk3D2VyY+8WpJny4Zumw9
AMHmWXNpimHOxVfK87wPLED4CIT9/OVOkHhiwppa7hW2nv3rug2z49WZYtK485ty
CPaEpRFWr/no5CBFWjCpu/CtlIhxple/tSGfOoEVGCUgyVbjI32Eq5xeeswVkdUl
DGkEhSoPEPVUTiLXnbpz/7AADyWqcdgCk+td0Yi7hn9KntXze/Gr2saY4fMaZ/kk
SK6Z+mxwfICtyo4x8iw9VzZ0MSeUFQXuOXqfeWzPorRlJsQSXD0urXXSXPRIcsb2
eyR3jmI7HivTKwW5O/F3p6pyjnNTd3sU6JPMrvL+iGW47wmga/VElwbVEPCljFoC
0fCMKg2XbZNEeom1F4oFVa7ln/p7wy7YSDcOaxtsY6bTPE+li5WbjWlmqR51mZ5/
sfXMdqI0hTwPC/IHDnyEsncmTOjePzps57DCbrtyPnAkgWw7XyJ+0FF+l7bmHSi6
vGFoHN7PO2p0yJL+hVoiGtoXfkUOVYntvISJsX1qSzomF3CYMjquTNtQRSV8DcWL
723pm4ViY748VisZDqQ88BdalxpnBVFIuszsSwbGbqVfYR9xd4ySCGZouCcXgNrl
Upn9s6qLTE7EH9T4XC8XwtWbuz3j2t+CEDoZVcYhsxHWQjC2+QQEGy8khuBuSjJp
jLgvRP4evps0gOn+qWy9zzPjpBIlFEEWE15ZKJzjpydp4Od923tzQ8AxT03SfNi/
4mnC7D8JEYt3BLCj/p/4WZ0RrdXzR8dVkiQdYmoXHmMHS9tu2o+lNIeQFVnXpDnt
R+foXOwV9gXvbcKm52IhuQ+UW9OQRcTxwsdL6zIyn6RRnXlT+lg/1dVn+FH/+VVM
9nK5/SACN+pukTO4bpNfM5zzG+Klmc/Riuz//9PsMOp24yJpLDwh/zcRkzW6wego
PwpiYA091KYAFxABdvks6aMXvFbJQzsrxojXae9QScqf2fK50DhphPzuBg9SqWrr
8LNKZL/nqKXWfosIpUE+0dnNZfBaTPz7vb5HAc4oBEe8+2qB0ko6+xvP+Nvwx3Iw
urxlxUFVVbbuMl+72wwZ5Ll+j6WaaO4IEZhklbVhn7NvI89GBWkk7q26Ud13wwlP
sr5KW9HeI9TVK8yh4v4SnD9TRJHhuTS9W8ol6MTx0Gt13p/bdSfrEp3FvgnDVNV/
lMA7hsv96jJzacM4bM4jpazZyaT+R0fdEDtvJP4c3aZQD4KdRIs2Xd8WCyxrv/uN
6npB+3f5q/wl08gzl8yA78HGPNt+ZVcRFJC2ANffLjq/00XrwxiY5h4FzcWJTbM/
bubOgTGskhGyR6N/9QQ80t9sfsi6PR0BFSt92CYQPxyqrZRV8w/VLZC1MQUEambH
ujVZE6L5fGNd7A2yCAbqhp55SToN2BtIfoo9BYVIqYqi+TGfqFuYIFL1dYRedSK4
xapZuO3BcwfGn2NSNPL8Q7hLtZlnNNfjUg9UpEan6RwJ6qezwN5O/q7T3G+XdNJF
1qCXIejmCnqz11Ez65GKbO5sFTayRxFY8YW/ruJpbxY0+KWn9WlH0qvm4aXyia6M
uQN5ZnFRIoOI8iSCmg/Lxc1FzEY0dm7e4ZXwtVM4xhrFBozT8iyxHZD6YoozsIUn
h564bgiAYQpXT9G1Ag3PIbelN1dYrnyeaTrpSCpnc2w3E9FScvvybnfvOmBDL/2t
il1vinMuSstTTNybqSKkCEe2Zh3gmddzA6UoYOpRQ5dXJnsY9TaIoavIhMIv+aME
Bkgh/kvaEqnFtHZMBDMsiDhbgq3199cxq7AO2sWb25ZvtMznnEBmHQyiUYH2Kluz
yA3YQW4gMUTbxFdjRdQtMLFnngL3JpYEEkqgzDX+xuzEiYgaAvF5oVQd8uuJdVco
ej2vtIe4SC2c+oBZZcYrDlTkzTtA6IoqrREWOFOLf4Do3EylNBWQFqDKYwZkmU54
NgcJUMw8nsuKsEani8/rZ8kaDquBFOd2ntiWJWBEAeUy6NOh64EKuiuR6bwArREb
irCIx//HXAgAJRbdNveak5NzmtW2O/ZKb7toUoJSsUHw7z8UBtT0y+9tzV41J8dc
3vTbQvMMHMCFi5yWKiJqnj11/foEzr9CXNK561cVbhtExso0c96fAp0m6dk/UVlT
K8ZlJweyxsT2TMp+5LzvqRxPKuUm4Jz2O1Ike7cdKzeadcyJ9tyzfaJRtVlRB391
UYIb+kHxR1u25ig5aTSiTtei+jTIVxrAS3LD5r77GYDId8+AKUQKpcVHyDYdX+UQ
Ebdr9fCoOfE/dxPS66SEhwW9ajfpIpinuFAwBqw3HM+DM6pkLD/M6qtzZp8DFd4D
2HzJXHa3zA5sxYGekXiqastXQ06TLRuP2Jlf194cqJo98mABkDbVRofymGzeRlZv
31WrD5ROfLkeu51i6RGt5S3ik0u/OXZ6EiCM/fHbdm6Yy1R8MiGzx3sD9qzMXIE+
XOV73WUvi0ELSgDmkuuVOUcmlClxZA8LhYim+dwUx7tilI69tJ6webj+mIUJrZ3N
vLVERHQcMUp1ah+i4mTGB91aHjrjN7aLrucw9jzStusYYVKgD+lsCCN2rRe2IRgz
oVpS+775f5ggKo5+Ul5L/r1sLggz6zTcpGc2TerQwBriQVMXs/1MuJ33l3cyV1v3
CIGhTZO3IZRrjKLx1Q2hGTr/wlMINOWwFtRPTGh21KkylQUpE2VRVdXPjn5mADyc
9Z0KXC5XJIzt6JEqrQaWlopSYac+pa3bGmOXv/KXycnSquCgBl+7G32imgJO2sH4
pu8adYiK8acpEr0EsbBrwuUpz7/CBRIepwbmhFqthujuVtBShSRnAvKFHofu0Wt1
EfPC2rlrT7EX8BXb/MekzWdFMrZUB/XBO22uF4/rDB2qFPl/lHLe2Ge2gleM05dc
Kkjz/RWF6rGKVPjWvRe/X5FmHCXXc9JZZtTZn6tuqeElcCgI2fj6qv4a0TdAfnTZ
VhO+xD8xcEReWs+Ic9I2eobus9s0kGvZaft3DZwsOoVmb7HrBHJIzqtzErNyt+R5
Iu/ab1GcBtXcDNhpqR7GJfOtInq9AIH/dk/POb3Pd/NSNj7wFUAjDH+Ov40+wGWi
ixT6GsT8HGGCUHDf8/MrOsSO2hhFMS1oXwGJf168vY0r0+ja6QISIiQGD9K8p88u
vlBnV029o0vE5pMe7up15xGtEHbKV/3/g14Opdfq+v8CCQTvl8x+jsrBAP3gv+5F
8xm5CEoAUNNZRMfjeuyoYx65+gCCh1cgEtuHsvcQI+Epy03NYPm/nEtgl2gPjeo0
KjkVEHpy+J/tFJEMQ1ymJFhFTEpACVJVpAnNHI58475OxLuOsr7HndLBOLB7hpU/
paXQmUqTU1o061aGX4t1iqa5puPqYeqAXXPNWWnkpKpwVdhGOKmdyT3F4QuHQneM
OaxU1jJ8rzYCnZwf+JF8imcaRKZ9rOKSoiWry2ksY5MaR3buiRwPezo1nfR3wi7q
bQwhACOhivrNTwvo+AW0Fy08sJZ6GpTc22kOwEzoUDPiorU+hos/T7r9Ar+EgUvR
2/ZOqJYrKfsOL4hdnzy3U6dNuv8ooca7Yp8pf837l8+9ZBnf2aTqzwKqY5dH/I5K
eWb9eW7uKEeE4uzo4gLViAEBAL4wuRNzWztZh7uDP973G+TUnowLEc3mYjhXJKQx
Aw5VIfdvfFVA225Fmjxlb9ILNYqwEFVmzKN6NU6MDncFA7E6832ZFA3QQ2638uoI
wHNquEh9v0p8YOxRBB2ArUeVnhTtnswDn+PZyqVQWZjs9lAKR2qFLS7bfP3zyOqa
HiGYqJKRDiJdGh+5YaMzKbxkG45YSndK5seWURqgj+VFriJEXyBm3t6he3xdRHqp
WMDS9KJfuwAgDcIoCPozkU1UFKl/WQb7OpCCEuPLZkqdcBYlk9XKbo/1DuWQc+dV
LG+Bw/Y+VTGcQgjqmZ30kheh7PZ5WPMevv1L7XCc4PqK9ouIGE9kiVnP1WvDXSfC
9nZnjNVaJFukKxdi9uVta83hw2rHXs0/GDCCxk7laKt9G9Wub7M9APSl3gXJvXuS
yc2FwIXyabVy1jDnqkfUNuEyrosJ/Q/EyeHLtituHpu+S7yhaeW5kVZSTaBZ8WAW
1T8UWn33Cob0Bn0eBVOXL2P/ARvyygslYqsY6BYf8WG58tL3uQ3cxj7L3C3goYac
TfQlQQz/SUdl9gDLdHP9AQILQryr5MzsqEC4eEJzFNUTdeLt2og3aAs2tn++3onN
N0LnUxLyuv42I4P4D7xxT3kNMXQKNz1WhwxmkFN2wTND2Dgf8m4J5sKz6UrMDx5z
9FLDhcpc2jkyAjOxFGtGWNaSFCciEjnNxqG40V/rUwIoOWUYV0MD94vj1wnP70W5
J1B3bdkEFNy76JNQ1WJS/cBiyCmM+JGU1StxCuvFeZFVdkUmNxMhuwLnLWT41uz0
uG7+nPfFcrksEchgTZblQTFbY78VPJnq8CZTqIp8DVwbV5syI5hgyUpT2mxcGNMK
SylBmwmL2u50XQRmKIymbCDiuQq4FhI8T+2BpbwyzNTCdM/2rPbw9zOeEr9wolFe
CxqzsVP4bRNg97CcPOw+tpGpHgw314hHcWKpf2BiooJCx5m9ND7z/+F8GqkSzsGh
eewZ9zLS5NGNe0JGk3pv4L8uBQDW8UzQNNu4CZA3b/WzcTDS1XMiD0zfNVOyF6Jk
Y7Bhbvz3YK4YFEykQCzSsg1Ulrlr4O/2WHOJfxcM9wNw8sEeKd20bdCvCQOJ1BHi
o76Qnf8K3avwFP1Qo+VdMFtzSd+mA7Bzh6hdQwP6kdFI1F105cCBZrThiR92PnM1
DNLBj/f90aGwbk1lvtaEdUx1Nn0XSxEJFpxuma37r0jncPT2rTe8V4JDeNCZ54ZE
zCRSvJTBweigo3XPsCSqHy7ZP/CTJdihRBWl9NxcuLBzTdfWoUgCXfxtVbc15P+G
Cp5irYABAeHSJSK4bkSYAp3dyEvnF2qyeUSFdXo5SYojub7LxKu5qvwJOW2eQNCF
aKIC6qX1ngoLympQlnboIGBSj9sXpK1Dhhw7Rwpi4l7zk5Li4DQvLErekMTnRmR4
9/jzr+EAXjQs7TYXfQybn8oLQKNNjeXkIMXt5rsGZ2p3cZu8I5sDYRnEEyHlZ80U
RuVk6rtpPBJtL7aS7vsb7xdhiMr75ALQPzD8ZD4NYBK/JgLfWqBpQToKYgTCZhsM
iFIEY+yORQylQmdawN1b3MMvwfhjH0ME2d/p1nX0YFFuVL080nt5YqzfwIt+k9VX
2pVPhB0dmNxBW+ITxYw63kE5OdOITRwfRGExxLp28fWTZErsu0B7Eb2+G1NY4HsY
ARnpod3SGZx/MSwnoYs4Ohhf/zwzFQvWm4uQXttqKXaJKWzhgelYo/SOqRxOE7fx
FD79qCbIw8YBFMknxLJacr4C+MKsKOhJaWGC+PF95Hv2TnTg/JIIVhtvcPvUKv0X
IDP6L5uYPWoWElsEu5+lchBOprcSU/8jkKKfp0ujdzIASayUCj/jI44f/RZC7rjx
OSXazoN/7jeeQspW+xAXtGuhFnzKKl5LRWjY00F5+ewG1ntEENL7iNCYNFoMqesN
9eRsLgnODNR4eXYH11243pF0IDQwvDTk5QpYukrHMrY6/GqW3Mku9EnkeKKr6zdA
VlICf1bL+Ja2A+GFZZwZsJcvFe1VJtpB1NtBEu9QrZqWGNfukL1AS0hmXi/K/j+H
bzd8mIq6FjqAOu6B8pvo9yUd9z4f5HFV80/U1amR8p6/eh6ZspFLkbVLp4s2XqPl
eRZ1hoD0diOQd33YJGBUcpgvACr5XwzKcNQHFgVMHSHGgda1MYhwO/c5gozplpRK
fgVeurxylK3Mk1R5Ubjp1KoLoQmhdNXShP/BM9Jc3Dnd9HNEgWdpGfY5RdY+bGfJ
X5phqpex8BkKuYcxSc1TqT2J0xSx1yJe4UYkQybUoZAKcYXWswXL8Rv+vxCLQ2Dj
JsssT9KsaWYRd3Jy+0dGuxke3LQlCOEPmCm/WO8KjLZQ+CoLSV3gtdIDgiOgB4jl
u6K491XCxONgfoNEaTZwRhpV0TAcw0P0ti4POVPszw5v3YjvAc1Te2+VqqEESS/b
KC7F0O+iqzh7A64IVranggLyd/640K3MxhD/tnMPngTDu1nJBRyJ+XgeUHI/mOd/
VG9ffKrbueT8msniTsi45OTBaIycPuAdQT2Rrwrj+A79IRa8ZSr1KM3zuCAZBCKc
++myLxSjEQFY266jZSqI3kkjz1/Rog3qiCVS1+MfFuziXpVblfnCe5+l4eog5ekV
n/G8775NLIoESWQkqQ9zHteJ83ErtkOvd/s4VIXgT9DwJAmn/5BY3G6fVLxtzj9P
jNaZVQ9Bh4wgReq6zN/yxBcUw9zXY59U7lGBhqEBFPw3xx7XmXIozCFApsodupv2
MDb/mCfZdhrj7E2+49rnRA70Kw7taRCRXESTykNXZL28/P1ykJ4f/x2X2PjbqdX5
FhCYhbd3GLyqdd/w7tJi2kanXjdrr4MZu2HQ/AMFMtTAoef2Vu/L5V/JjSKoqgDy
LnbYtUs6FBbmdASj8KbHtaMucE5eMAWs/yuabFlUhelvR0pq3GJoGgwzXZKHGOFj
oxwm32w2z5PA6ia6z4JowJUfTiqvF8YRnMV/Jgy5Lbj7TIZLpA15gmSQfov3sAV0
mwDZ/tI04DPH6IRHS0aON8SCtT6c2XjDjCxi1uSawS/BYYmY9cQ1v9nf+fpchnKp
NdzUgiye9xxornc4hujYqq+463K2fQ9+VkyoO8nK+htM7bwE8dU3zEVYaZ94GE3b
Ha7Ei0Fvl+6+BrJyQssFk51P8U4LHQtCuSbj31UuqtPQsKY35bqhyCBkbnxMWWyZ
q6MhhUSJrN4kaALMBr7S5nCIujMArUcIW/QzEgF3bOImzFZkNb4Gz1fQ4d+JeP5h
dk1763TFdjXQ7cJHdR0LoS6hXW70ZuHUKVRxw4E3+Qr9Oi7rrFBDCP1td6VEmwiC
BfJd22c+a5PnBpXCdvBAWnANWGiSSvMhkY/oJcenJrShf9mRQ/z8REAqoNp1kgso
WTYZL/9aHqST+HL8BQ3qKSdgniGsZCFle/JHww/F5eFAml/KWmak7FvQ01HEjqfV
ByKlIlm77FWWNsuz9xaXOwvsJ2ievNN7Kx0iLGO4MtYwkSCd9w75DacVNIWG45RV
gR25MmD1TNdlOBdeNWGbgzfAsVxjZhPWPc/UDmtuNgvn3LthPZrQmo/cM86pqSPV
zO3PWNX4wGTmtoVyiW0kpDsmfsBp3PoULavhJk9hT4RkKPtgjakgfjcd/XUY+U00
cGutkdrg+9R6gVVXqs4fNH/JKo5K68BOT3bQQasNNXf+fvndTKIZtw4KXXVX4h4C
8SIPu5M7dpNRs1wfWH0uS2DRVdWAiIAtS2BaiiCIWNAxX8M5/dve2soY0zhsWzxt
gs/3rcggK/nv9eXlTctg/xV7fxEThjC6nvECPASmtT9/gRv/3oiUYPwbzvQq8ixW
84kMiSIZK3CfEBKfMdMCJxUc5Q6+cViFG0YoM1FV+upOFAkhs+26wamH6INDfNVJ
Rp2L5Yt4vq40BejJMEeDh0JbZ95+DL3S/Ln9VAegWn3H3aHyyvNimw+VANT+9FzK
3TppYhjQES8XioCdNkx9w5zeN1EPeAi28M0+2JrEPJh5tMRbkMJUvOItAiJf/YjZ
VCgc8JrYPrVuSj2oPQABIYmU9ZXeuMGgz6jT2dpRDL1fHNFwi9wG/rj5o5O6zcnK
E8mFPLsDpmOgL0dN71A6K2N5QT+yWsNeDo2RsMRwK0JeSZlJ7WpSxXl7ld7EODiq
D3cfIu81fsBc5XT2ErEJ6ONrdhjLGXKUi0a4u40KtvjKIgmC/HRJwkYQnW4/4H2m
inA6wB6xzcLKX1Pg2VPQx9VpUoNe+qK55qwjFz3eBoHKt9/GhBlldK8o2Bk2W3v7
9W3hiRaW+Ehqp9BvhtBTvBwUSHUUNod9WFP/9oLjWE6p5CJInbctny2SzUzqr400
+YvEJe0ZKLmXLgx5jWX3BYrEPfLRt7zQuzDLjys03aUwud/luYZmdpqhvfnZOW63
gJHDu19/B4KQsWSsVchVF08SwsNfpyezqmwUwCO8RSiY6UhBXsN7n5IKwbcnD6On
5yFVeEXDjq0+acs3+IiHtquHlrcqnFsdF5cYCB6vvWPqt7oRUkJpjGxwNhYv3bsW
2LCaX7gi2L9Ri4cUu10RQ40TnNkWUYdbXMUvup3GzSiBc6+iKAGX/ovpB/02LB4P
0KZf7H56uOUbrhFzJFwiWhwS4DMVC6PArbhTjmIXui8icYyZV+RLut1YrDcZJ2sR
xLRtugGNYCQ5QC5sYBSJpPvxZ/VDfDvPdWxfK1nGkJsp/eFDthNUDEnjH5c/Fd49
CBMiFffA6vgeFJ4qcn495p51oRsTNJwhjrOhl1o9XhMkQGCR83pWJHMGUIDuOUI2
ovMq4K43KY4CnHzTwqGkZy2N0WgdJTPbgieVb+Vux0LzfdCB9OYXXLIg2945Vjo4
w8S7PD2x8MKp/6GUG/i6rng1ZR9XjkJUas7h4Ly/8CYmBvnOdGmtfe6E1TjX3cMZ
CqtLfHTGgjc5tzAvq56USP497H4du/IS9TAX88TCbZVEBTKVLpcaispOPOJPUs0K
IZ5/WfFh5cb5hk0PXs7xgGWh47u/zoTq3dfOf5nUIpYDiup17CCiu521vWBCfTFl
eSfA2GVbGRHSr7xzqMQthegxjdxj0CktNwO3r+9pvhJuRYK/h1F+NnVBPtcTEBpq
/0wI9yoXwYAHBoBlzuk/3qq+lSFizTivmTuUE3cq0y3CNoBGdUxvZg2U5htq2RVV
aADcp1y6RD4qUbdEnCQt6l36iaUFMwkGfvVUl7BKLYunyTrDNxsYZTyb7CieEvvm
Wv2Me0/yvj92nUmz5dyyT190tfeO2iTo/9SSN7SmeEOdCoKdGyBemA3OG+i2x9Hw
lj+IIOt+Lxcdh8p9iKudqR62r0wm6yCW2N0n3zCn+oXRQ8XcImZtjxFBe/kjg7A6
vO39qqjDMDAd2O+H13IAUe1w1DJlRtJ4z8yxrM1hmNcrM7WWGkFDJwbgWTjmCbHO
U5TCy6mkSrfiQ7lfMEI1WvUtv9lRr2sEurSXJ62pIoj2RCcjHndELTxvppMJ+Hmv
DNvX6TZbHgwx5REvR6FaM8cJEbNi5QY91pib1QU8kLmvNDssjZXSUXhjHizCa8uq
HKTAP4F1K1JPoxRzoJOpWAbK/nNl0hFmpki3MuwqBNBB9fhhzJ/Yfyd2qZFnxFCb
+rSjhTmu8iOFh96xNArXoYAwQfeX/xVOBeerjLjX9VjLVDXTJFep+U5XvqwwEzRA
4sHDj3XfcNDnulTGE2ohQMaGTGJOsimT8FeHtTEpG99jFQ2wHXcsH/JMvojTesVk
TEgB25Gt7h2WGZ3ZBsRZGFAze4ThtS8Za41oo+lqUlmflz2IP9YCXVu3Hp3bLSbQ
XAhm5H5dkF06ubM7ZhMtZlZW//RWq/MT9vOTU6xPKxZRwtK+NPH4Mqzfn1wPXb2R
II97hER74mTR5Tr68g/wjTVmglmF1kY1QnrDP4/495hGc667uoOV0b9zIy9EbaqQ
dtQfQXrVXG0SHJtedkMEzpSh3TmvkXCt3CLg2uSjLzVvpowRRJIoldxd89PHgYrO
1c36fWD0qZLeKH4qmeKZdBq5q1Au+2EgQH7vJkVWTa8dAdAHnoYWevjxe22RQymG
jkmeltdmSuKqw74D2E5+DuXHPz0WT2p74XeJGrfeCg91t2GUSOeLPD0yYHEjtnGs
7EzA/sJru8xRiRRZ2IwH3tY2yojWdsjAAYrdhi6Tact27JORSdMrhWoZh2dKGzBu
hoFv6K5gAHMWPXYAQ73bsQ0ONASdlf5ndW2bzSmoxl0UyKEGoZpWFDfTOR75q4Qw
kugNxjNaxidZgQy4joUtWxao9FuAV3hdlH8DaFVmjVZtfqmjdBstRbe49u1QXMLi
+Me5TI0yrUP0gzwIR8ffZ2EH+KO4NDbuJhudFeVvHBObY6nUtHBckJUzMC5M77IP
k4uHtl/zEh6iRlF12/01/jKLKk5NP8IaXBOYeN8yZ/AIJ1iy4DZnRsZzlV5MuchU
BitgB/5/MBrt8Q5A19o9zESoD5SxC6/nYsVcHs6dzCZOyRacI56bzXOsWQuzZ+qB
M2Qq2/c76v93tZF0KTIyDU60ivQoFl129TzykOQWW6Tt9pBtKmabL2MwA4KUxTk9
XoonhjYDqh+LpEX5fvWxq8493QrxS9C/eNRTfDGYAOIEN9we2EyEEAAnkBN6uteZ
1SY3pNe8roCbU0UoAvzsVTvsFmIRrYSdZg8YNmtg0wm3IcbacEACoE/0RjxNqZJW
mmklqQewwGpKonuUW84VbJNdsn8k4WCvDwXgGAiG3U7MUgFVL116FjYharPE2Npm
tb5p5Jgo9C14Fq2APu/rD3Xju/rA7ZJp56FWlVuAd2nAxnemFZfropw1UJjG8YuL
Gmr4xAp4Qqzlh+Y2ZKT9fevujTzKotqrGUIvAQpwsFhFsD6tOkwgY+Ur6APWQgjg
BkM8QJG8R8yHVUfg9LSk8Uc08RhNd0EXzcz6RodQ7Az5m95X+hEo0htkVYyD62dS
YUdmMI8GlDwbvmK4HArRaoSYZRxzi48nWBrfzDIELxYrl/Du4tsAyLCpEsv2RCR8
JuQaPV+uOEtHnxwUONdzcWE9v7rmxMQbcNcn65xDqwzWA+ATuyJ39f+KYC4m+TCF
r9OUfjrqNtym8sb9mCqc7NOSk7RyVsl4hoNYLraJxmubwqXGvFrGOeGxkfH3L4om
/C5mdydjtc5Lbiea6s1zu/K478pSIRKdFrciugIHTuLOcftpOTMGMRsWYVpv90R2
B1FwGPd7ITq2bJPzdPBLF64hkn24uG1gdDhcS9hjypYnwFSU2OfTNDUUlHwIG8PB
Iiy9WT1lFVT2icJNn7+KennjRifYcfjLi7siiMAq+aeTg3mieoPoA/oDQL2GYkD2
ebpKZ53r6Ag7qlrQSRX6aC0Zcqfy51azipqPwl+310NWrqYhyte5RaBvtTh7+O6r
e9aktqO0h6jBp1tQcmuwUgeOsclrATQP+QIT9iy50AiqMVDCA0jjOGKGmUz/Y78J
k/xc3SX2IPRRAou5pUTWkAwND/HzKkcoDub+elt9j3L5AuJAZqstukS7kvKro9jL
HxE/l5jEArzZHyey6HHPG96yjPUR7UFBDCyuf4ML8GQLmdsrAQAKb4LbJSh4qDLz
Eip8Auy1GqAlubTSJIeVsUS5S+CVKdxzfFTHadgeK2OUprNaX0BHLvsiLvnrHS2H
KGh0vAP3hqlC/KpIRP4GS9FwVkpLp/BiykLwVt5+SG/cCJTXEXIxpIAE/IUbww8M
R+qtPtwHX30BCdowPCzLUXLnmnmSNFSGqwzOQcna1XtlnLby+NGJual4LlKvI7v2
wygmGZLRg0x4MaPkN4bwGwZ3HrVt11cE7QewmKOmcIkL6kNYKB+sL0fadSzFZs1Q
LXXcjXIlCDXT+qH6W+kcnEdLNWxfxiMCsKfmN3Ofx6e5otgFI0dg4rEuI5Gf1EW/
r1XdCY6MBZ3rXuwX2/SHz0spjlSNJqmqHoMjnnCIL7AgyeyP0FbqXbS19LfkHv+m
eCEPdRL3vwo53qzX4eUSV86xnFv2ktWTXKLA+htlR6/uZaFZ69Sb9TelMz6WREMb
B9iLVgtH74HS8L/Tx5AT7qRg1PqRlrYtAKgyChgWYjY9rkPBI5v7mJeGVqgFbDYP
oLb3l1Ux1Mo+cy6G7z9K+gdVdq63OoiShvOHmqK9n1WP3zEy6oWI0xja/fhVfkj6
ateh9RfeMZYRh3ZY+Iyl2z9UAe8LKhzXyBpGqQ34TnrzPdS/5qOyKtFrDJ+b0ur9
euEj/7rpE46RuSdLd1UFLQhfBgqAdqdbuG80m6eZxjqNSfzpXOZWtLWetBl+WaFw
pcuhY1wMB/O/3kxgU1qzaB77e2A9ELug8PFjyaCSWijf533Cxn2sr1qfwXf2Zvx5
PeLWQ8VRnrUpQV0oZOVkx2+3L7GnfhLD43mz0yqjQ06jC57xJtNzAvS4bfY0Jp++
V1hsH9U/+FsWixqclHnmnie//GXkRL6z4XqMQzAXQRzbGqXnPvvToZu2GS8nnQm2
DBf7yYUVGNMFwPUE7JVMWSzKMJnJA2wt4D9sdVVBSV2/tgU+IIlS4QyJh8VwN1aW
3AkDAUl1LpMrXIloOfGzj2oV2c8T0IdlOyaxdSiAA7qlxV2NsZs2KCdnCR8b89un
qdrL5Rz/PBCqcaxc3rGq6J7iZ+flvat0bn1NoF8xqsc95gXhsGfveh77VyFNga7n
WEU1TCihJDlt3YNR3vacnfENbBkXMT9XNcp0kCoOKJNwhVyGaKpHo/1ie1B/S36O
d8Ab2rYU+zs2IwjqPOsXK38HBgQZSQzq4JoBexYeYGa+lnShJsigKxROjJv1mRFA
jhv5lPmJv6k+HeMr1wHar8N2zRCHmKQXm2wP+HfSj+NDbcGwdwyNL16xH4mr8+S4
wDjfyH95VKjaOKFpPn6SIlleQjylMHjsk3pR5Pck33nqVAJjxYGuVIEIxGcjifU/
kyg71IH3CaVoBJ5f2fhNh3WFZNEs6WZcUB6IU0yYJAQuZEYhIrQYh9I7u3J9Feev
BaY5Um8D9UKLPc4RbVeB51QKTAk4vS7VWOWfsX3eKTRkvXiAIRawMsRi1+9jNwS+
ij1I+jZLkvB55buF3DGph2SBLSyDMgn7d7M7QXv86uJvvXWIgf8fOuSKOBj23KKF
+fXmJ5ZqvJGpkBDuYohD/ln3a4Bxw4a4nfGEypqK1NWI8riNFNpUQvNqXhE7Qwo3
B5Tewbm4TZenyI8Dk6wbldVcprpxybF7kUqtHcHNieK9y6fbCSUSpg0JmqgmzohD
XRlVrh2uQ/Hl0znAsnOriApwHdeWlPevxtJ/PKS0h5AlKIW7baCqNwGQzdb/Kxmo
z89Je9Wrrh+VuRxn9QnY8JdqwNcFyjfkbIu69VinKq1FaRIx8JkUayuGFnTrwDM4
bgwn/wtMA3TrYjdfDZAxV8enxeRC1WJhn/fz7kWmtAebazFyGbGtlTTOi/6oTI9m
7KJqTJV0CZ0b3MT55DPWWb+yzX5T0qOAwTGZ9DnlV+a4bxxy0gKDbVCEtex8II+k
pEdydC73sBFmxUfdyGHcsguw+RPsQVqnf9V6D0pC3o6A5gpgIT2UG/IyPRYnZgIz
amry4iH2YgL5f7DBWH6nhLj/lE+7B2dPgsjsoGwwsVWU7KiwbNhRIxPt4U5K/7BM
2uRmQmm7hYix6OM+o5e3yHEdNDcZ7diIMF0rzHPxoYjWX9ZirF+EZDh7rRxYzxmd
fyWso7QYbji0r+V6YKiZ1q6U8BYorWJKAOLSmwvkKvUVP4O4lxDsIw7TfzZ//sq2
WTMBxC/Qo7ELX4kI4r5kZ2MtEak00MnimcIx0oMSqxEUMwUDNRzx3wZyPIKXvxyx
7PGEaBo1pMYoByTJ9UjNhG6glpSaJr+IoS46dN3y5d6+vfE//BETBlySSp/eN7rK
qnRCT7c97yx6I6ZrVgThVcRM5vKx/kgdOoibfAFtaxjMZ8p5ngGmvt1nu1oN0Moj
+tuRdmF1SxOG7XvgfhhUFf5Kh4X4LVAHz2hJLNYWgAMYcuECo3P9kvW/7t4b3gQR
Re83TbtHA6aY2DdbuM4GsHX6j0KCo5V3eRP4BGHrGmuv4p8fDJQE9yDl9psyBOTb
DjBTGCYad1TtuRh7tIYBoByL1TjcXggoPgZ5snWQul0I6qj0YZlyN3Nz/DABjfCy
cApPzdekLkxGuL6Wq/H3QwBME82YvtiZgb0c05N1P3f8FsaKf6rITGR6kC0k5KAB
vOFXiJn/9wDzIboP1gyp4Ke9khdpJ+NrHJqNuYid2tD0XXolsTTG91adQMWpWgzQ
rI56mzsOcUSn3yEX8GwRMCbTIPH8MkX+La2XltcQd1rT+K83xWyogDrdhao1umXF
8QvE7vmpuYWI+TF0gdf8nsH74tf8vBINhs2VqzKRzwL4V1bR0KrwBhPK/8zWMeuK
HB3C1JZZ2qUAYpN8cm4+eBcu6byXe0oUUFvUp4VhdOkiz0jgWJsbWCMYbcRFmgIV
EcISQO0nvsyDUzkyyebe1uPF6VegxHBLcmI9DXyUrPNGVAHYAWFjbWzWOw/tLI3G
4iJ/cePqSuIyGFEJZPkRXU5C+OVzFCxyLWn0AkTf7nVkUpPhyxNAPJU/Zzp/JmwB
IAZ3bDHFYSw8vtplcCerUNYwMPVapK4Rz6kauyRAJvvpt9fw+RlnvMoZ58wrPk7U
2r/WeyLxpoHjYbFeqKdaaPHf7Ro95pCAvxSHDK+efIQWoQZ6Jx335ewwCmjBM4TX
rMZzIVn6HaYdbf6iYyNb7Z6XbToPBVm4IKtZd8gB3ZrnBYNPbooNgXMN61JFdf7J
NN7WypQvT4ISlr5TZ/2o1EPhHIKlEN1sUFxxg0YC5WiostcNHZjDQmC8rgpW+Q5U
MKtZmnUOoIbSmkXW3gb2ITtDRiwFXy7bY8f2NJOQReBN9WNrMfxj14oACUp24b7F
Y7RXkszQJpRAZiO7eX+X4DlSY5YhB4B8LeoAT8AxZIHRHBG7HU3EBbSTjhq0UNT7
d/ll63LvylWwPlOxOsnO0h7v7A97KoYLpcFqpWmTKQM5myr1ieLoulFW7/0m8WIi
1bS8dpm5st4vbSLQjT8m4J22QiDkzgr3sgczSvc1u+ylnBH3iEzk+YC+ooyKqZtv
TM/AjdXZAhs7X1kmVcOsiG0uX4gKdReqp43fynOA3a2v0cWrvA+uRP520aljH+d8
zB/xlyVLoVCRXx5T6k/Qos/2iCICDzz8zf9oPNcD4A6140xLRAB097gd8+1HAWO5
wPlAGKD6lMZ9mvtzpWLS6LmpKoFMIHTDM0dQm7YGAn/4p3HGbttkiF8PBLr8kGDT
6VDJ1jLG9TwBy9tj5Wpj0zimrZt+gZk1xi0Q8CfY9238aa9iU0uaHIoMF2tAziMP
2J5DFzvMjkwFCpvRNO23KvtdbbX1ea/w5ww7lLqZ7vwzLhcXhSX90Hov1l26Spi8
0DXVcQkUTq85vpVIzthkauouetQciWM4g9aJHF3I/Q4oUlDJ7aglvSWqeBN7vNiR
wVMDcwPdgse193DDPg6e11NpIgo5LArhWIlV5OqfHCawX5tTJcGUJY1r0392Lxos
fCjq2ejIYpClHljr1illcU0cH5WmN3AkchfQzg0Exmwue1saaL+CFmDBaQNPpeuO
0QsBcZh8EQgQuEwLo0hfA7hatRo/hxBTX1flDw35Pa7I9/wrjQErCQvyCw/ary9C
c2diUOrtAtfvtuQD3VhYUyKchqkfYLLIcFFI5Vo1PbChlo1/Lomnl1VNERaCM5NA
iRnWlxr22e+yUR/e6TM/zJIOoSr1dyk0kNTqxvUn8ZgD+zmKAj03vWqghY4q2Z9C
oE/xAHLYJ1ZFo8+2RC1636JIpb0UAaJ6hnp447+Kp4LADEQpcGSx7TP09qaQazKt
YS+Vjjlad6wWoF0eg7jbBr6xq889SZLl+tXOpsc6RjT89JPzYIyCtkLo2QDLEv/M
BdkRHUtZs3TP8K5JEkGiI6d8Yn+OiImSnJlhfmU3nXS1t+wMu2C+vE/Jh4AZW0DX
gsKDMHLJExQZkchomlaMPZ3EBrEzB6U5qu+2IQB/sTtdsL0+aFMcXDYbmolBckNA
sQEYVQ4/VgV8Ml0uBl5HbW6116bYsSR6ReqomqvjIy6U3Z3I0gyJtBEI2UQQt8Y3
0AbMD5gTgsir9nhugrwhX+ALvxtVF5hln9wRZfDWuYGtk4oCAyPvGXDb2kqNkiLy
mWOwQa1V6ZQQAW5OmGfh+HB2lUMbcxK9YpeUl+IiY268yhgbIKDoZODgSXCITzZ6
TuMhTQRazTyKLZcODHw7PESdV3j1ZjSZLaEzmQ3pOob0xJ7M2b55QfZGPAaGg55E
RXvP7ROSDietSoB8kxb+shlEYwzRnI/HGVSu5FW8tWoCOKPJaIcCvktGGiL4nMsZ
msbOfgIw7SRlQynPBdeHtwJduQuwu/rTJfnzQdonXqElUm6KvN/dT17QZnd7SkVn
xHrZZ/qh9olAU0JZ7/kSU4EQqhYV5n9EnotMAduy9BaMP9Q1RzPnc3dISjXknb5R
e8oQfqxZeclWq+rGZhAPMJJ2ZoTGPcVK9xQ+R4pyxC+P7uvIgwlQetqzwEGMBmb3
eS02uGgDfIp035B7wCQPdmsvyrKsEnwZSO6iiOf67RY/yf5WPEywiQyfuiL49CrX
i4Phu/PL+GPlIKK+z1BdcuD9Tr/WKg9dc9WmeF6L4bgaIgee1oJtpIW68H0mHKxo
4QeXJScqBooX9Ph6bEpDFfT12uDYH9Fg65NaNMmzj5caNMFiO7++VzR8LZkBYKEu
R8bOKN1mXt+uTbqQKWjwV4aqtfiFYX+EBX0zamTLesxtZtR4CinpESYMxY53Ys5g
OmwihvfdJCJjE0R9EErsJl9brtyMYmG1obRGZUE7Zcw0eTXrlWe+QGWCno+o6tjA
L2C4zkGBSMS4IH7lD2m92KtzUCoYIysd1ajCAEv2fNIOg4cZX81AU2q/zHnLUNSd
EkiMKW4gXYtURVE8pNgV7m4ApBuuQWiqpIJngvuBENZIEqwWb96n7ndLS3sFp+Qe
Ox3jATWZ22GW5E1x3d9LqXj2alPo8GRceNiAtQqv9kPpI2JznQaS7wA61wBzq/AS
RHyvsp+svPmD5/Bq0GdB6aVY1Q1J2OaOWF5R9niIP90mrMU2qGuMZOtnFq4a9Mu9
70qnhWF3aKMTWMEc5C3EZfeBSHNdocuS1AUUr595TtbEGPr26eaDEgvE4CMW1Qzk
Zy3qEcB1p/aX2FoD8jG4mrAxQg+kwu7/W5mFiqztqJ4Vqh0WsolTvOoyXjOME1sU
py9OzbANpWV9U1EoCEJt2LPYm3Ie3ivYBZWvY2bLbq0mrEH/iUUIEad9GnVVYfhQ
xnDDtrxdBGMvurS8IjQyBuB8qfGoFwITAhGgINiZUzoQsjij2wI7Sj6+dYr7FwDl
N602Gu/yp0jWhwMce5ivq9kXcGqXankHWFfDQxltvCzxJjV7rGvF67XfPA8qik4s
IiKJ/F7YQDq6n/IVsdSAFox0zhmzzXajHzfH2UPL4gxbD9EiFrnw+29BLj0+L+Lj
3Yn1c0F81PzvKQESbIB/pZnb2S1a9JfiM/qy75NaRGQ/jaQeab0PIH7uG8FXqj7Q
kHpKffa3VKKCumfBG3JumgO2z1X2zSABlYfWO6zW9YtKzMJJWOjgHAfMH8HZMoMb
I1jjLEp0A8kf4PZlyPr+o4lAEKdcRjbgmT7RdecmsV5OW2mjhWVYjhNWavjiVSn2
KduJ4pKXeRKOyNUv9PyGuF8salau2o0/KWXSb6c43xaPWi1qnzjf8m8e8DxUp8Ww
/nH8skrySfiBFQ3qZx/rrKRS7R/sm9fhv+OXVuQoiGM+WeqfrVsLeoNN7RtfHkXT
kGnq3Weg7+GNaK++Hyb4qzA5T+ugnAGJVA+ezyxYrN1wOEzlT4rHv6bBWo7Oaxtv
TmWJlDhkTCmrQkcSugg11SNpa94thc3367YL33vr2IerRyKd7lmi1f+erfuTKJ/3
peBvNuv5/0H7a1zmggDfePj374dpGSXnyKXpTNzwPonPTVAMEJSWRWCbivndkJJx
Bkxdhg+k4cjTN8xTtZjXiPwhZYcVJYZyj0QjS24M935PPq8egQJmldYiO5veAp7Y
N/KWy8yWWOlSp0/e3Udjcq26/wW+8cx+sW5k9hVyV3dz034AT1ZLH/J1vRNkiV3o
pj0HpJfKYIrL6WdtXXNTKVgR+B5fv0WXBRE+WZsX2Grr/3Jn/3KL7ko2y2nWq5/n
B4KubWYK0iyNYODAOGjk+XOItTFtuO2IcF2NwcdblsWWgy0T025HK3L3PPnnVb/V
3JkxZJZbU7fHT0ifgi4rx6YXpUEcnH7HSwyVb98P0JAwr04HfD6Qth7EAUcNHGmu
QAnwkP1EuqLGkO1GtYcwRuVsd4P/GnM/hxguG/SQOWWfN+wtxjKGvqcTN4/fyBDh
HDvmLc9bA3uaDBYsiGEzGuZxGiLmrvMECjx3mLh6pHTsw8b5PZUKuO/ka+oHEpuJ
tx+RlU6X0DpQQWPq/3h4hcPFV8P1HZk7vQpTuaOyOYVhCVYTOxnBTQoYMZjm2n3u
wu7nE2Z5lMndmOVZSymebAuLsvHi7Jci6PyZJGLUYdLP6ZBZmsNKP9y+GKe6o1sp
izmyakGBEWWiIgfQ7vSB82dRxTkWcNqHgApsGu+vX0l4n6IuP1EhN7UcusC+pNY2
GIWbfL9HzBxo3OPHKZYK2c8oPvWwxufE2wrPAKNMZN66dPNLOy83yTq3dCw3nWLJ
x2wg+K49dGRTBRfxJcg2eMO150IG2Uhr7I2ZH25hkWKgHdQmNx1USk9ySsiJFYTy
Z8mMJ+vGlfa/8+6SBj0f/M//WRG9n6/uIIFwtKrbaXxwc3XE0IF90wXRqqzIOfbF
Dn1SXC2UhTL3RKFrBTOKLDT7sAkt32r8j9xjXykV0skuzoYJdDYigcgNp6UdL6Iy
sTW6N6C03i9FF/SyrWnxGdopEq8w/aDppTS/WKl8/BT2OJRmXPGon50Menh/SeCX
Ud6OKeJk7vfsfOTfR4QEnF0zWVEFgVgf8mQ6e6P8sGVyhqSQVple2IgFCrbcyzOV
BUzaazZQi9iVROnZu+E+pydlIfzZnfJmfLutQl2BeOrpBpQy6V67cjMs+qaTDXvr
TtnOtvx/onoc+d4cREIqfIddpaI2jN6a/tPrntrVURYUHrbqQ6+aQUjPo5YYhYQ/
R3sCht+62j03ExjfryWrBgojNL7hi6sE1lwJXjWj6K66pNiFrd73EoqnXgVWemwz
74FTZ75cJI5jnRDFxbiaS2EekzFxIdzMHxhS6mC8CkG+42teA1eGtWwq6lAjCur8
nK5SGKoCKEBSZ2Why3/RE3W0ta31+jYTSfsir3Qsd0lEQ9BImmOm0vc0E7sXNC9g
txhKTFPuUe9u4hC1VgZNEQjmc9urmMl9tCpfAjGjaZC20cjYWKP9ZtHJ9WuUDfY+
wCkrh3InA9cPbOXxvUDfkWb7nNAdSEHMMnFRP9kGAGrV146z3/e566M4MqI4UaRM
QE+d9DsnXXRT5x9EtPe5vHyEa0J1X7yBfbu3/AZsEpf0aOMXAv3vOeRHGH/4WFqK
INhZP5CxYkzilZ671k7nhMviI4sQRMWjnoVhP4ym3Qqkp3y764NuPuTahCj47nCM
Q16yFsITEQDzKnXSxFNpD632Ipy6IfYJq68YfBSjiGqKZfql5zTyOCzISm9P87AP
BRSvrspeX+0c29Kl9cKrXq7pulexF5zHkJuUz3rAArvmV7VJcSeML4UHNVMeT/uJ
T/E4+QTjLnfCzwPhGA5WP4dvavR92tcTaQH7EmZYvsl/yI/h1kJcqNIdCRqdHxPB
EByVYj2C93KA6nNK/wRzN6CixDgbFZajNWAVpc4RZ22jvyvvRBcyZ2bRsu1gCjAL
vVCWW7cd4GWwa1yOYyIULEXb6RVfVmsZghwXZ4MwhRYjrl4NLduJV3xYY2D1Bp37
TVcuhLeEmgK35dTT4smxfpZQaBEGzz0cwDXCoFSU5ghig1dHLvrueogKqbMmxONm
DisulOHhRHRdLiTE+TCChTzq9dnaQQA1RCQcmxA8IPjyKBbU7J1kcjNpJMzt2kAA
T76TGDvT+H7O9XwCEbxguHYcUUtHGpu8HXIofid9fjqcJCKd3It9/p+Hc/onP5YV
JBjlSpDUnATMhvUaXFkloJGsZwuWmZC820Ji40n0GpBecSeYN04k8zYq0ENWZcHk
DWYoWi1dv69FkAIzWaWnzsu/dr/vcZdE7br9k/UWUNo6F/mQqm7DIOk4u8kxF4uc
cR0smSOyysveTKtZU7ryoU3ak5MTl6AHm+bGQjkAVAKK2txiPhhh2U2HoTHn/GmU
Z7e4cszVwK1OIvnQ/XgLbsQJry9fWtUgJi1W35eWxb91+yuOVlpYL1zyxYratAqD
PyNz/f6CAcL02Zw4HI9WpalwndzBZoNDKC4pjNUXr9I2Kw17kI26Ddh5jdwshG+H
kMCunzB4sMZxVuMwiUqCRlFmG2i+gXwyhfTryv477XHWBE4DoyVIIusrzCp56nIS
YCZdvhhq82cfCtdDvuC2Yv+KU8mxirVPDA4bSOS+lzclFqYm65HR7j3iTSwB6Bje
J7Wg+QyzNyipqJPFOrCEfKKlz9nZs/xUTMxDKWs85gClyphynBv48/4nX3VXFUL9
rB0qsBJNses5bZ57ffe6qZSEwQ/WNXSBy+WKUaLa1xMUZmBgjKnwXPNT4+qv2Kdx
cnBykSLk4Ao/HMgRt0x37C1n2wQnNYUAAg7KrxeY7F7Lbt+tdUN/pPbs/LEdJUnY
JsZKAuUU0YSHTiI8VW0kJrTDOlO0KtjlRVKpv4KcLlRhBN1ouTEGs3HPBxuDp6Vb
cD84Y8zuGjq8iOtPTM9uNQ0OpoccHnCWnY1lznnE68zlq8JS4kaDkPrJwOD7tGnn
X9xO76zqV/u2MdnWfR1AcBQW7pymumd3uYCA2CpFT+pZlXryS71En0CZx/bCC+rb
awOK1SsYvbS5eTzsEoAkQVMiDf9JgJhneaoyCYWOQ9eVowMvWG10JFZD81aRl7Vq
IwPheLyxw5FyPGJNMpKOCf+05yUdDgw1COUcnfN+/wPv+JDNZxm/8ctGggoN511V
wZQeIOQOPiwuZUin5K2IrsSHFzl6g2ONELkUvwSH2rNN2LmPYLjbJPItVrDg34UM
zJhY26aH/AXzmiBUmaeEAUK2ewaTo0PD/bOEL6v+Th9Js7FVVFUpNjmKoBPfHpJd
RaqKBmVYu5JjSVii1Izf84YIub2qTeo6GbwIDxeLdLIohzbw12nKq2kZXlTsUleN
hfV1v7NefG9FF5LRt3brAySiZLIZNrDZs15Bz6DCGqW4hC2AVIjQ2h+9S5pA5wBz
+VVJ4O+ROzClPC9fXSNoNXaFl527PfbzBOuqvFYHFIcrU5Qz3jorZJRYKVZxbwOs
fRVDLeLe6Y0GefDNVuoazSMCEj026k09rxfkhn7eGDDSMeqCUICJj0Sz+3hFZ1YW
7E1drDVuJ9cyiKA7BQJumiByL+u63YxHXa8Dsb7FmOSWmrJZFXdhn4Ok04XwZLdm
CnFZdtdWzmq6WMTpuEI41gzUUAGsFwYh89FMgd9y5mQf/zeevG5ziAgkcGBhbn2Z
9reiVxT7cfrObgqqypMyUMCP41Hz/FJ04SymrKFGmuYj+72WqUmvmuCBkBKMMFCZ
sUBMcPGJsBhDNW5GouQe3+v0NlPWoPrO45MEHiXP7YTxqTm29B9QZigoRcoyhXCu
EmosnXLSilPmRn5+imNDKcGYe6JmH29wRtqWeLJKwaCknsr78gLwLflqu62DhSQk
yXWn7FZLCbpyasQ1SGdRZz9nkKx2EKi2qpyi3bPn/35BGNRREK9zAGwAhbBcHH/a
d5WhdkOn70eMQtYgryC6gFvmtPRLD8jQZFBjLS35AeCiBGB8ZMu+8kUJ7VIjHlBx
b+KJB4MKaGfZg2g7IIkKXJ6o7bxwp9XmD99ngpH8WcgcFG1LVCELBKr4z268pihK
W96AwjTKImmrBjzp9weB9EfocHH4u09zngVr6fMumbajma/fNgxMAJyEdAAPTeeR
RZmjA14bg9EG2JD3QFfatOESCs0ZUcwsQHY/YhGdRuot3SnpZpRdI10OmawVQEvf
m+zsrpTSMQjSaxFVEE8X2GwZh3DSb5UVeibcM+VTHAq+L2e0VqnexK6Ec4xuQETH
SgDuyN2YdJQRFKyRihTTdWDQJatdIfMzB1OwRnPoRKtrZi+3QyD8gLOkxs9CFW9T
Aj2EoP+KNCOFKkHB+R2q9pa9RHkyyUCUMNevgKIjSzPP4g1CXEothQE3TMpPvcFB
4dlbg/6lL19BksdNnvreCzO75GCW0Pt8SKNdyGdd5xB8WPjJl041DEETkkC4fc7O
GnP/Ig5+sQNpx3MsNjGReQr9MHKIc7xxn+peW48TbeFLUm7ChZKXVh1pfXjDXqaF
RUm/Z5uMZcFHu3q80B7PnajYWHYAFm09gvmry4cN7V3gEGnr1bUYBrczyDvEZYi8
jP7ubofwvTa8U5H8GQ79r14aeJbR//fk/Lel1MonZtsWIIAqndH9p8yndgdyV19F
AB8WtvtyoMyyP0LkFI+sKimZESvUl4D9IT8mVlcpKUhf3To/7teveWBbM2zmkfP4
89nA0mw/8aAABujdBK5xa2qED2Ndf+r5sW2dJqzS4Nwjgh22n2GipMEN88XmnKJe
z3Ut/3gOMvWiqTvSEMCbhsAmgZyLOxyLR4he8xS3rnLWcP51xMXM9xGFMLgqX8XQ
1EERFwyw0956zxWYFoBUtC2Z8USNbbWWZowTod9HLAdm/l7/u4CLnx0O7v5iSTLo
EpVXQuC87SbihczYEoZqYtSMGDYTfOSS049K5zO/ULKUrOQZAN2Xg6JZCEida6tM
GJ0gP7VAIHB3Dx/yuvwga9RZstsxGxOaFhidB0HgULGMyLY4C6uHocSiSFJGcsck
s4c9vlH8CSY+DF0Wb1+geysFKFNZ7QoDDHdhVJOt/brg0LP7mbIVAdrk16uC2Yuz
g7VhFafEIhrr81p6balQdh4zJ+EunUS0Zjq5Gi2XxA9LCn8wFrw8gAdlea4qXrxk
OsXrPgOUDTxt1hNfkRtkQr5U83CLERgQejhYOkFxd9F4N2IgpS6BwZOCCK6FTaq/
owXaM3wOAKiY82uQxYsfNx/6Ym0zm8Az0h7BbNs0YtLjh9XdqkYGoXSGszl2EE1W
hDIgkTVsWyvS9AOkxSzbovxc3G34NillZX8ns9jogrPRA1QsFl45DliYw77FqK+w
ozSL06EhXoxxPdPlhZYZQhZZeLOQZpwDHkw/fZcvrPK2lAiy2Vsfv2FBQXU7M+uh
MjqYSqxz70gh1BCjyXgEZmmmIKtId7yMuOi51qsm+2qyVHG3GmfgG3KT4Y0Cslmt
P30pDv5vyXjZLMeQj/KC7nBYn+oFc4n03FCcsEy8YzWYoHhda5VtV0fKuZ4wuluq
2Yg6mPRVCX98eCtv69ugJNgzeNub+D8+j6MZwdTt3VNPJZPPEhSGnFYRtoYAfjpu
6ZxRFa19gZOVRJilbWoCw0AG0LzD+HvUIns0c3xZPq9n0VyXGkIApmxaFxqg7wnr
/0RjqI7G3+dcJS+PLring63+YLe8cVtABwTPixXorwaiZDjCkfet51Y6b55B1nmt
KhWdSC8mI+nyeK6344damfY3g1mDe6NXVmQJfwZ+SfuNQ9MhJLJABFRSm3AVpcVo
XPQ7EkR9av9VTF5NY0eNBD5OtaIGrmN/kcBebAPaWX7BC05GEcnvKxNU0X8axVd8
Cw7gCy1tbGqCVPqgXvUvFWiV5AhWyu4HpRI+gI+T3Xfv81p3W7WJiIMpSIzHNR2z
CmHuV9q11nPq98qBuOJQbpytK94pFCEYSzafEusrzCImtcnaz95s/+1+HaXiyHq6
2wfckPoxgBkbeg/s2xyLFL+rV1QLeeP1u0TKj1K0wi0od9bB8MnHDJqnfLiOgV7t
nBcKcezCC2fg2m7gbwB9sfKR++SuyYADalLuJ0ILQJt2vuV3kfl+ogdQCJoJ67NU
hXt1V2i2xUGDL8vU7s6vgIoaAMDVal1gGrcDWZI8vpLq0v2yYyw3pfRJ676k0PQr
fHaYxxnf3RRdn1D+k5A77v5nPrDZxeVSThVhJ6grxBKhmiOUWxZXfde9dGOXGeDa
F3nrSYqfcP7IZY1M26MaC9dkJR+wbxaRClsdEo2eOIe8Zv5X6rwNLkKGWY9uLdrv
4KJbhvOzPgM0kAJqMu6E6R3HvDhJsPD9TzVBa/sG6nEut6hwYCyhQRmjEKjiplWw
RG4AD/+GZs6XdsN9+463Mg5nlYvRiIEjGIZyBIuRIn0RQQU1sxWo4HvyssfR7WmL
C0psiFinNTCZTuOuczAyCoFzgm8YAHUiyYrCoUzehOqrvdNREthfKf1fZXWOCSTw
zUsRCEJ60FagfhL29J7X6Fgg5SUhAM8E93FV1CvmNBfmGQTSf+Uwl4+9u/jOXvQu
RtblulyOm5zWAXnelZdzCs83LgLUE92T+j7piHFFhkWJQoEAduojW7OuknmZ8lDf
hnXR1ggcJuDLz4s6DBl3TQ9MzhbrmHC3fN0kVwSIACyPq261bdNG0Elcn7xRWEH7
mnxcQCsKoy8buygq2XklD2tIbUhgevdqW+6764JLAWsTp8dUetlWZMZn4CSqw8XX
4RSgo9dtWX1JNKTdhrp2pHHX7Z3W5IAbQqTH3+ypbMuimi+DlTuzXFYNFGRdoTBi
qI0Bi9s8l1loKP3Fat1VQNygoGn6Qtz5LRB2vjaRAPSQyxHAFOsajgZTx6jNAi+7
BX+k84c/jQI55ylK3CsueNC82FHmYfuEOLjoRMPLWVvJqz61ppQTlWtrv2ybJJLe
h3xaUNFd9TazZdUcpJQpp/hyj007avcCesxtIBv2cdKoFRDRpc7hzypoEmtQd67D
K6hRAYkeuwT4M6O5UFExyH6IlvTJu6J1Wu0IXQm56v1FO3kdp0eK4coYsdzkiNlI
uo3acuWLRg1vqm5WQHR6TK68JyvBkjK58LehjMhlVNLR57O3pfodrxoz9YcHG8z7
Q8oXqBzli5WkYaj2ap2Mhi5IY9l89ceFL7CirON6g2eEeqAf9JQ55wnm4j51Lv3X
XdeU1SnC8OX621GhCI4hUqHzzJezwhkLevWfEwpnFQrDu5OMlnJJi2TRukJ8R3NO
N+QZbg9zxaWAblbyFf9K5Dv+LG0KPYmff63E2YUjwnBKVEh0pxmWFayPQp/CuWn1
ggWqdJSosdjXHmV6b16ic8jfA7rhI8B0n//dMJIy8GMmCdQjKRH5qAt5U+m6b+fh
tmAsUVlRTbys3lTbX3MkY0i60a0CiMtfr+13yJqQNrh9ZKGUtsYT1CRG/GckaU5j
fCXREdeTyLhcnaZLnRGW5LBjHBWX43gV7HdC2BHeDtrg/4gf0f/KcCWhfz1DcVvm
33u+LIUXoJT0h/vLtsaypAvjbThfh4sL57HpdB+RuGG40FJyfrGDlgUJBUvFvw4i
BJ7gQe/I3KECL+4TmeYt5ad4+twiBwEcdgMelG7Paj4wSf1AXzTe6IPT9kPWtRfg
8H7/fUnhVkCJfWmibtg263YnpcrWNwhqM12N2ouMFpTOaUhhUjEJ+fVNRvXoSKkA
a83jQtnZWIrpCW93EF5rcSw/mGxWpIYmtCprOBcy1vb8t9Dpg1N6OkioclGWqgBD
VqHcoEaDz9q8T342ftCu0w1VKJaPdoOlfSOuXPXSLCrwunbvsGUviaratZyLTIYt
orB/9vtyRtLlgsuSjSoPyERl6Tu+EkuOwHfzRmsYG+LdiQdV9iZll/hrPDpVoAPd
iDlPwH4okTCr73DrHve4N32khCWBILiNn4cA8MBwTs25xmaBvbEQ0hNLQ+NSdQ0/
jRF88rp8lRR09E1LJsT0+nOQO9w/+ORKAdyXr610SkDWm6S4Iwii+Bo9buJNUr90
XRVuQKaKJPQ48U1wji0hUF7RM+FNwb0NOJD5F42HU4uAg1KP7rYZPL2UaEz24Be8
lFh2DdIQG4nvb1JO2iaF3LPSWXVEPdp8qUCesRorYDDSpowc6AkjzIccGFxR3/Ro
wAxBaznpm2Z9PfTmM/radajihoko+ZP4CJsCDp/7vkKn3oNZ6hzUToyV995wsrey
boGPpHTZgsrAfi5G3aTg5SQjDqqPMWwPq4r1c9MXLDngk1fl+shi05Qt0m8DfgJ0
7ARahRbF8wQwSVdyn7Tndvf9Yhggx/wF7oR+Mn7ttn9l3UhN8qrQb2cDnEEIT4Tj
iWr7QmLHuRRxJB24g4hzLt+wsKCdV5vZNiVjR8JfZaj8dISn3ebhWg/ivQxm0E8G
YZ6Ny6BfFN/eQKYqb17oF8RlDCHCoA5dQe1yn06UswWWvm2HEtVmVMz/BGjBPMlv
2oJmgqohKPZPkbtZMF8S4E/pYFGMI+YXCCqbfUjDyWKb5ybnbVOtrQa9nk46lRr4
O71ajgc5PqRwFb9U+BjUSb+e0jrRRXr3N7QbShusWUUvDFVFu29w2jzvX0Fk5OyT
idwzbkK3HsMTJTcE6TR/yGMh2LZzTaMbB+zlsEGiEQV65IKEn7HKvJUAvBDiKxk4
QOvMvfS/RKItJFIsuwq4QJoRII0G2j/yJixAwfXVpImI79iOduCa+9yaZ3mdQCSM
83uc+8pW3CDRBOajuYR8EAvNqvZaA/JTfvpDjBcKVk7vmgJuAKYhhKJ469WKa9pf
hFJlBqfI0OoOCTdTq8NtK7hFzyt59dXSl71UVP62ja7SlzE2UaNgE8FL4eCogxWb
KqehPsXiD7SccYq3WrT3LiEe8tzCkZRDthZOnWvyP7tmOhZWFcPmiWpljHlvyqm4
rmp8FpkJcV6xO8iago7LHrVG5oDto9k1tJSaQASphttYonulYItV8sNDMasq8Y3p
ATmRwo+lI06+HNtyiF9MljN1QAkkJ1sDnunAC8OwdtA0qPiZsqJ8lb6BqmKcYo5j
0WkuWMZjGEYf0tgablCk5pJ7fIHpaicy47k6/Je4j6CAIoKb6/vAswV5LF6r+PP/
MN6AxcsL706vyeEOZOd+gfSnddnET/wLb5fosxfUMMVjnzyf92pRyt2IglJV7UzK
rmTxUj8U27orBcz9it4PfTg+IcSw4264X1edV9+YKAqh9uuRkuc5Y+6zho0NT9vD
r6HW/jadG3EziDvqiI4NDSWzY0ihHY+xr078dXrol5y76Hy2Ca89L94OkXaxrpLH
qmxVqxV5j73cG9JKDnqkdgnktwedOZKM8js8eLHoFJq88nr5bAiVGyQtyLC8WMYJ
R8j/eVy6BTcpsRDcu87NpMT8z9U5E7LE/Sqdq48DtAgqhFIMTjBjPFwI6E5X8/ZL
uRGit/MowbByHcedLLFFaQe4uL3S+WOHC3uaOTVdVt+p90VOWJRwxPPfIt2fIHEr
lsVrsLUEvkgC7ecum03OHZDRPqs7BUqdARIFWlCBsfcqznKwJdV8LORanUKGSZqN
CWFEcIRIuiVOasrZlGOAW/dl3PALquguC16+blarOoxI0mLcOrhCoYSYyEVY4MZw
VvfDslijm4ymudBomH9/hi5dUWTfE2fx91rFbToCn0rCKXp4Y2QO+MXAAWvt8Ht+
KcVLa3uq49JZmxhLM51BeXeM459ylFTEX+TsHiE/zCkCm/A0uTSGriWUBRyLl93G
fbGBOBm7La7s7PUIIoy5OszKw5w6iHybLlf2Uo6dLXsVctoj0+LC+1kbRCUPD4gb
h1jxUuwNnRJE95dTUH0FEhPEgAXaJ0/Bw0vToI5ZDbr7m1hRveW5dG96Ms26vqHa
UwWZ5tN+GfM7/kgOrs2ZFZ3tcbuNnVD/kSw5YMsCgz1Fza+svkmSEqFHVY7HTGVI
Bngg1sA3/35sqJbz8smLbf2E1gm1RA/ZLz2e3vjZ6JOe4Gx7LFqJwJyuYBd2/CgG
H74/KVfbdfVaEnLkusCCots62Jl0wlQnJhBAy4PUnBg4wrm/yQ1fckPM2UMdJ8Cn
IjSHKR9UVGbLk2tw5bGJKSSEVoH5zpUUWZ8+nWEjE2Uel1+c0rcBD1pbDRnljcqe
apEnZu2O1DWr+bx8CR7vtdjeuVbKEAHcxaFhUCeEZqLzTu0KlXR1oHFb1pt7o9vO
CiE9YQnbCm/2poQ0sYuZGy1/Wwj1uq8l4YeEBN17NH471p1otGlmAyNZKzQGQK+f
2en38iO295Fi/VEi7iABmNYXKnorPhpPLMyGYWytfRP3j47nHnS8bEViHEuyJYXe
iGKSH2KF/z/JLK8dQXX0zyetmd7jNe373b8fjqwJdR7yy2MWMtusEyROvL0mcChu
6bpWsRVC0DlFWZrQakVJKL+cE8QRTnwB7acZ3ie8KC8V2rcB2LNqGSiGjOOGfSbO
iCezCW+gmn/IfoscvOwIzCd4F/S3/SSJQGLxvf40OFQSxfSZa1vtju225R75Kyl4
ycDLJLlsoX8tF8WmASFVIR4tpsMqwbLDaeztkfnPIwtQrDriJTP6Bk+mkD1aqZWD
ljYpo+vh4AtbIJ2KBttXZ8KL0grco7GdLL9ZwUDYe8/U/9taD5sk+2ocC2sdI2Um
JFzo6XqHJNqoRX7R+EX36h/05oJ1KIf8ClwxT609VtFUD1qxCWkQB2Dc7mb3eefc
lAv6d+HLibPqH2pOn8wqz8kOLIM+k85p5t+V8xS2tKCf+n9D4cdGdr0x1iX5L80k
I5g0fjNVGs1n1N+y46BHSTzPcQpU77AzlQA+Wu2gf+CRhxaYPDy6Hm4JVyhlp8dv
u3jR3I4pmVijLA/YdHxDr63z4DV04+HIQKhke30xU0BFp/PgGm6trB22LXaAPrGv
4xod6tO4n77Ckd69ceuNvMTM8KiTAwVjZ3oEMWIUwVRpAGgjHMOm2/larhL+V3JC
YZpejbmKaQpwpv90ILB3xzGyYJDU3avLmAA8JpbJZ43zcWi3lfLbWEWrtntY/qh8
F1Yx0tV38z6ITKc6kUlVMmUoeSofB8eliLaQAYOC0hpnsAS9RBDpD5Q4R0Bp3vFT
XA/CxN8uWr6OG8r7GaYp6H3iubIJPIM5Xoz1/dAUP2nizMqa6sKtLmwcv5BW1dIE
6juiMS82k/0uxI7pl/T1yljjxhgM7RGWwX4vZWGwJz9eQQRdqQjG729HaTxTS9t/
VbFq33ywQIo8mt9wqdjbhChwkgHyhBfFjpMnVdTYpK47CgzBhE2Uw/Ky8LH+jqle
2eBR422gobe/td1JaFgVaHgEg+qTJXCWfV3VzWLvRQUY6KlqaxIi3Ev+NU4SvvUk
LdQor48jB/ZreHjQdCRtfjDbZyIULDGrrLwlqEPw0uKt99ayijyzaWYViN/4yCmq
HhvbvHnSJ1EZWAVmEJ4bDDA0FHG5oOWbZAgFWuR9KIBwlkQk4A3b41iSq4v4RXQX
0jH9Q0EP5O8G3dkkI3vTXQZmARbzabvReO0Ai6tizq5UUniFa4b0pIp2iG0FJgrd
K3qvuVCHHPYIEXbiLJnkrLf/3YVvYRAAuT298/9grosxAmMrlNNRFwIYiPnIh76G
nS2Hn7ONLLFGWNawu2Ddu+f83mOiO9/nafkiiA2Pv/0+YtpeTDuOOs2DWC5toJFO
ff8eppg1lpuQLgdZ2qJzireRVilnpmUL5w2nGDyxTQb4+6MBfmsxCcDvHholhPTI
63/I52QTFrWYNIPhvEptIIGHc8+Pyu09ca4f3Lme0VqNWVgCOLEvBtxr9ArkvOJY
OnVmCLtkgc3GgfF4cP/T2Q0rU5sc/Ds1ZkRlIFiskrwntB1h8VpCzsF+zN9K78El
X53rusU59sZggiZlXX1emF5Gy5+XoTjUtLRRCZMjeVAN6oWCsAT51Duz6H9LdhBk
5USxuFHUfSaToflmrmamE+suVbr2M1g5IpQilSvmqdWe4lzbxhOq4c4yqOy1G6b1
hKpjv5wYHxb1v9u5n+anhz7RRJz1tYMpwyrrxz6H13h0ngLma3VnbSOFfqbGF4v0
e8RbynKGFmrbfKorDDrd8UlD5B8FZQtU40iaXZYGGefPxTTyEKGRGB27FqumUKdW
ntXxLpjmu9SM9FFJc38VGQqdkhfidz5soWADzgEWLhtUt5rXyeS41319pchsYG6o
WjEiuS+hrJx+ORIaxqasRiAzKQptBUB0qj5HhPeDcWyjb55UA/LeNG6XPJV0mayA
2fHplFavXEKY3lRZBoNubQNqyKduj+ASIm0q5zcYw2GtxESsFZPEpilMiy7gidvT
r8piFW3aOOvqbsw7AuinUhINIBT7M1wuB5ruhWAxJz9kTkOsYlkLP+xEhDiYmM5V
mUhbSVTH9fGDeC8Wb3lgbtQTnzJ2RHEbhvWinYUViZ0wuPkscmJIHXhVAe7RCfNw
FZa4tQHBGOjKKhMvbUdGpcFscKcdADMnJ7m0L+doRIKUbsLfr0evlCtOK4k54FcV
JORau3oRexNJWUvbpu43um5QFunJHv+ffSqOU+6QHGer2ELgls1NpdhnYnn5oY3l
fBYHGB0kNA7eWq2DdSVP77u4Ol6ScwLrt1syeqRiEr1MN/Iy4sBmRwkgPyhYlFLI
8UIOcDEyCOMBfgpGHJ3roXuDaRyqQa4goWSSUEYfg/nVydvoh3BDL4WrCPRwsScM
64UjTu4F3MDHDpfGzTaSzb62koHlBLojf/t5xE1pG1fbvp5jFCQ3/Q+34pLIDjXn
KinA5t5DDDpP0GeD5FHu09HcuXgql/fRFlbsrqpTqb1btwBB2MHh5BcLddS42ZPn
9DhFmF7eRLhMruQrfA4Htm4qam2XafNHPJhJWLygntwDwSKh5htZ66EgvJ+odIco
lFAcSlofJCjzus78JTAQ1OIrS8O20Rxb4xgdNw43IH9uUFHsyGmbiAR4Dl+anmAc
VbRhyCeRdoUzhC1/tHbKsPq4eJdIqvAZcXK1J0URFwyIkGQ4YrqyikH79NhYvgsS
I10oGEjojnWqbZtsz5wpXr5fQbanY0y2nzQnKeMm896DzX2UaCOFW0a/Y6b+TnpP
keyHoNHSIUTLH1u4YHo8JRtZsX85hB3SbZmzkYvxQ7EHgTBMv/RnPqDNfsK4fnPe
G5TcwynqoyF/N7ynz7A45PXHPeuVXK6BoX8AtIT0WSExo0MEVXiZVvL1Zg3mb00P
OJNmhN+Yw6SdZk1rklLXSojb2vzKlUMwdTsiV2eOkVJQFq+QVvYsyvet1WXp/r0s
NdkZq8IBOYgoibd0cY3bywM2WKT876fBdK2Vdk6cvsgbYtiRqn5+J1GHfU/2YuDm
ffKNxt7wTymWIa1cGkvY3IYlvkZ5QN6/avsDPhuPvY/+KSHlRYG1eC0Z+TtYJXv3
CV6iDHbYQ7S2wPBLEtJOlcGrEpOEgFN6V6moIuUGjPEz7JDbPxhFm0l21P9hAVIr
1c1r0xsZb0T3ndCgtLIe6W2XqVwNhJWYswwIgTj7K+g8t1oEmOUMWkZOuIpDz7A9
5G667Dn87HjdVKD9lZ+oGnGlzj9RQpTzWUhD42yL/lzyTnV9LnPP7oo2XCDpMTps
Tu56MkDCJRBxqXMc5sOBoOsXg5qy5B3NodoxP18xsPmv8dAw709YzbVRVe8z9/Wu
C5b+Wrvg+fXw8EECoI1rhBk8aGg19rNDdGd6/yzNObY6ImkYY8uEAsEBvwI3WolG
G7iFaOA8FktMyVT0O2SlZlarHfyFkoPBKtYEBsysVo/XACY8E6a/4qvtBTzzeUDl
ew0avOiuHHEzJy3KlggL3OzsgrTljjKRpj6pwfcDcKI8RzEtrek2tcDr8fc6EZ/8
L8MDHp1cb+0qVNt6UlfkH6+5He+eUwZSFLiTivmWPhOz/WW5McfQi6Szs64gHw0+
cFEh4SsGPfLUSTmkSH3L9mrBQmwdPwY588eyhnphyPwXY25G+yyVwMuLtUCE/bZP
soz+5hIk87vTJ3DePERNN2mksm28HQ5bbkCaNNcQm7u2CeD6f1DCuaPPiwDUpzbj
C1QpnMqGicY8865nnAAEHbp0jcOh5FN64pcR+xUkpCRMZxyAxJtmUwXkBTouohzP
rSN1BWSqRfv1zd+EJrY3OxHGZty3ebGmFnv3IQUxxErH1xGyzLplmidpvyr5iW4X
krgByobT71ehMxA6qQQDpAJBaO31yAzXLLkmTM7sfFWclZbb4zWxNk4FjiFu565r
W+H6WBIQxA0y1g9oOaoCfc6wG+JtbAudjRrZHuOi20LbDXtt2/4yaN27uTIy3zuh
/LKTWRKfuX/unOwfKoioGw4N5osZWZP5kQalD7cSeb4Kc1XH/AwEroLQ6v9nWNb0
dNEldw5ZE6CmeptR9RGXtWgpgJrY+9dwOscinIZeP1eJT/tg0S+0ATv+3vfI3x9h
/RYbZcz4K06VE/wc1W5DhFPzDf9JIC45rLerGJ9uzjRacCYJjRZa5ZI0+Rx9Ae6K
MUvSbQ3h9cAQsbFbxpiWYS2EK4UXAidgdqNOh0/OP2e2ZyMDhlY523fyHv53ZKt1
2dOYySNK40S0TE7ITJ3MSNwDGRcLl4agZIm4rjpQHlpdXz4if7bkmeTgKZ/gxsOf
eNjCK+KHYxBkF4x3/UTpShrUr00b7yp4paKku+Z2S/qx8JstgZ4MYiMEs6MR3M3L
MC0/LCHwhdImGrpfLdagFIAcfUJWcYkSkkZfCkeDVfHDIZB4LXyNpgBlKl+w4FI4
4e7+ztmcTohjBYZWPojgE05gcn7G01gNgFAhCj8Sx7G6OHxjVwrMpvvuhzWLs3L+
k0N4fNRBYpOJ+sEg53FySqzwAt2T+jcz96xKNtXBG99wqO5R1/ASoknDDz/BQSFs
1Id9DCfZrs9pDkM5C4Q+1++CX5ae2vG+rq9c00mrwFu7t8uHR83qIHN7cyrw5zBX
hcqSCeHVhGplYbeY+JMBY+pULEwTPLGuwLAzyJecaTGa8hf781WTIDP0QtP1fzis
aXz7RLaGWTicWIQOh6hWt+Bc1At93X7RqiD04kRg7zX2qtpSOL67GKH2PsT4Qt/K
ym5Ulsl2iR9/TCUyBjofRkfLwWtYfJyDLWiU6nVUPm15o/L2REeGYBOgIbwZrvNn
D5UE3adwzstbRBE58gohtwmE1RqKvRyHaqGU2bGGp5BeLnFQ4Gi1SrMZBmyXNPLa
bnrsjyOTFCWj/Wm8fAHDIR9wdx2E58B955XdpZMGq1LOXupRxqBpFmKv8Zbh1JAu
fCIP091uBTf+hCLN2nlrBs8hac7K154P4NRwuPTUNe/hBfd3mCCR2CdTOwAol2vi
rr2eEtkiNoPt/SNrTV6a/QHRWl77w3l+4es/kB1bK/pWv6Hd21BKk+MUQ+It9zCQ
xpaCr5SpeT1/eh2OYRFNq70BZv2oS5PZtMD9Wyd63DN4bY20POy5fUyPCZhyzNOM
wvvnDxAvtve3CvRPoxwDLKAS+a9yxpVUysXNMDQ8Oce4UJ/li4fy5OV/CMyMNKbR
eDNG2tgMl7Vkzh01DOtuFyuH0Ao0ZwxyLUSGK5duhYowCcRCGhotnuq7KcCcrwCb
e3TkGOXXXHh5cjDu1d+KTvKKP7C0H0YU6XjJGr6gaM/CyyiufWxDkXsa7g1NrMh/
khqkJb/XYhWaRYrkY5XLhNjiVlPG6wBrnpg1Z7P/5PMvlWYIjI9nxqc7xK8HfrhH
ickYVXogicFz3tJnynR9oEZ2Pozx5JbdEoq1BNgUuqPCpWYUTWccsLwvWRe6ChGU
vxtkK9UXU8+2pItUIRi1v59Et+r9y2JyLTbHKWvYpKzAQZRpca7+xQ6/iHdmvOp6
nZqUDHI+dzC6rpIomVJomW6Ug/fSp6yQ9RicWGNrepBf7c+uJrkW4nikDfFL208f
6Aa0eq0sNgnWdA+MulJc9IulZcrZ40eWb9GhHSzMeyxVFqp5rZbsk9x49GrIxNDc
jm8AIld90PK1EyCXMR2Ut4BTZYuIuKRo83+tBO7RS8iStBX3BsWj2PZZTfzNjzlg
U5Hk+WoK/dIA16Wjfohs2A2BKLORc1uFigh/kXaLPy+qD3M3i6nOLi1spXk7jSKY
TwOLWPIbxbfpRr+X0Cr5XIonGx5PSJhTH4TFREcfSbADGW4E38vSLYZGcqN/aOuh
d8S2Z1UBW0Rmq4/L+RrPMWte+1xuiNB5ambxeNR7hrp79sBvI+VLU6fPv74EOADd
iDyVKrixxztsbxekAbzmxVs9XIbPa1lHLooxdfC//o3VHnTRo4qDXrwtanWhWWMS
NrqaLRy8mmaeVCGyq0mJOOgH/THamyRv/oDAY2ZxuN8HfP/g8T2QCzZTCxrURUR5
FH2D9nUyfXzJEgbN4RKWNav7yxjIYTRm9911zocEhf8cc/gtuROyiJjH+S2UhbjY
C2wi8Ot2LZK9HL/NZKExmQW/F9Fbs77dyyTPqsh2uMiO/vIA206YhWLchfApoDL3
W/lHIH7FEQQAMOSAXAPe51NtD6duUbNv7GAjJBxyF27yc7Y7R4rPKUU6q/pG/swg
/2FWZa14EcJgwBZBhekOXhmxhkeKDPxmBzrQh0iNYQSWrjDyBtESzyFTn43U1ZEK
/CiXbjbsRRxMIEDz/DI0NiGNwirNf8rqt5iFNkY94ROuJPfKfru+j60g48ftTeCr
3lycdz1/xmkTcxjFVmEvEgUIx4Ucb6Z2RS3VhI+5kI6/tFJ7kqNsaccQ8oitJEl5
lRxUhmM7I+tvddh4KuCPBrIyqpCUogDA0QR5zxgaM2wqb5TnZ/INq8ejzy6zZ65e
b8JoInrqY2EqXvJjEG2jQnieBy09oiW42+1kltxcTopLuuf0tYEua1USD8sCZIJv
NJ4fOYq/deVBSI2JRqzoYMcTglZHVu6W/R6r2+Khu3M19QsWKO0MgBzlv0W9w+7f
EWmjmFh/a9Fu1VxJr5rBtwmu3XtGZhf/X17ocwVNVUfJJqWrL50RTA8974/XPYOD
87kOVATIn4dGpcWwIfAo1W0W/ZYZEp9KRfOneY4f03ycQOYYhIq19QWqIA0OuHpG
mjFT6PKi6KQVOUnWI3J1telW5I8+QFhxR85K3Cd9SlWbdo2oKymerqafvAR48q0j
txmfbyx3DBhpf2OnZmqK3GzpRBxLNFolDqAUL25EF2YlJr+ZcP6YThGM+U4W0OnP
LGZZ5MYYToKjE6AxRV6rGeuZXkTY+86le4GjdPYaqIBlX1GyyC5/jNikMbEqHpHE
jSFiL0Z/L2DetKTuIDpArmqBfYHTIw7CptG4rppSxwTShLS1j9eLgeCE3WQJXLrt
cMCwnoLMbKkdaChzyNp6lgRXAZTj6AseW7RL2QCcvpPy5c8rkaTeuMLoIWo2pxRJ
06PTD3kfiaSzx1CpGXdwu4TDzj+ve8OvCvBhHcwFXeLSlhH2W0XaMlIh+dCLGEMv
kjnn7hZ9682WNOhUbnNkp+JHjWge9RZGkcLWD4fr4bHijEyqfpbDqVWgPCHLUE/U
prY08GJpaDnRHPvwnUpsyevSGLTP2VQ6zo20MfZXR+M/NLHGnOM47Ms+IYPhFCCE
kAEaPXBzg8IpWTVEyAYf3nkqTMBhz5fJBl8PPL15Y1EBDH4UWKb985V8K6HBONqa
1/Om9udVQkRUTnKMbESBnWGjwQxGSzJezErp/WubkqSpkCWOL0n+bGm7v61MvD0D
khwRdqM5/PcCuiTv1NydHDB+fHX7/VO3Y02Bg+ClsrbQRM5QAsjDTWowzgn7h4ul
MfHXSNJtxjfwZ1/aI9sGyuojKCC4j9niLG5ea4elcGn6LSyRzXd4Eguy80uHb3mK
gG8BzS1Jgt7AYLORuR2SoTcN67mHgq92EmsN0WCayeepOZZB+bcWSxl+Vsdv2p6H
ZDRVsS8LZsVtciqXIqUcVP1WcNEpFjYc9Z1IaZn+EigqH2iy6p/n3Gj7wvEdhqte
JGCVGWgb+hjv4fuYhC3SHKJffSoZugKhYflH38dlrKgcNobcgzaDVrONsIlqxyrJ
riDPF3XZENOynDIhYxbnV1Sxj4SSc7NCk/h9rlQfCXkYXJCcMSNcjj8RW64Zz9uR
z3/4g+/W2czey+0qcjPO0KP7SInNdY5yfgjYv7/6LMrL+Y5dbjoFyK4mcd9NWRNI
R54pLH5LuMt69Z7MpyRY/rLjX0v4ariAkZhTEl6b8kL23tPlKYFiVDv0isHLMUXe
jSgxbT60juJCO5Hv+zjZNJUjB+imrRF7lFef391rDq1aG3UJ26Roqne3nKKUYXNg
3dzYD7RzdnZ39f2+MwMsHs0kXLw5DKGyUPoR2Zw+wp5O6IySru/HKQVkTPNtrtrq
2jx9VlI+n/M93Z+KpYcseZDFd+uZNqbI0jd76wpZUqXrrYfvDvklfrfz8+d5YdRj
lwK6loUKisqmwSdW3UF58kSTYd16Hl6rJXy/ow71VTO1a7cSoaRVmeKqgp+MNW8C
WgxAT/AB94fAz4Ti5vHi5SYGjpTxlt5XmHhrCIi29+pwH02Ax1Ar3W0JdUCekxNs
rfuiFYfwmGEQnwQl+7whqpPdICI2Weu0yAVTKYmXfmrQV5XjnaMGPTnPA1H1Z7mw
QdmN7b130hNmrMn8SwjeGARMQ4u8oUUXUwtncNFJm5wapbg0dM/czHAE0qmGlIfA
wYiAH28KxJiWV2TfXdrvYlJkgfWJIAQOuUoyP/SSi45lAIoH0rl0TtHIDcyirkSM
G2VoiK0J5Y76EvxONpB5R1PnLjG47k9bMMN4yJk0or12WBBQ5yVCYmRsVp8QMyZO
G9r3zLL/op9IjTgb9dcKw8Ml4vk/U8/aVopMZalLq09+BYqwrd5mmyLY+eiEj7wo
tGWLrYFKUrKUVxoxj7ojUSM3O3CESJ0jOGdZ1YTPBFLQN5wrzcjQ+KRYOZaP3aQT
eoxXHYweIiXuIzBvOLgrMg0jQQpBjPiGLJfQ8M0QlKYfNvjoNjBRrgViMQ8a/W60
un/919gMzqXrQaYULEsrNQKl5ZrtjZLMSN0fdh+jYet+07qp9RdO5yzx6UcmAODg
JeNCKZSi396PhxTiMyParQmBSR0anz1SmdrYz+Ygh6Sf3vy7PjARUl18M/fYnQRr
KLn5hHF2MbQoBYaauFny1/ihKwOmWQeWp8hd797YkB0QxGITOXzlZGagjXYVnkPu
Xaoy47+SRfzJoh4SFw+JiOKacPsX3OjNRNKh2/0wz0aych5wnk+vbJb3+AmV8PyO
KNFZESI3j8pX6Bup0XKwtEkduinQ0U48KD5klZ6ol0r31j8n9xPJjffRAjFPqEVU
f5cos5JRYIhT0tWrppZfnYoyMtopGf0m681bsunpBFYpYCkrHmNSKgqF7l4odLgD
UCtkQfvPAyEz/aphgKPZOxsqW/eLNcNzHB1M1htZGb7Sh2wyuAstj4yhN3tasVk/
vjcsIAFbGVRGYePuF8LfWAZcCuLBgc9Db+axdQlK1hiIQFPxMO5Zbtp7Mz842w0t
YlsuQn943GpgQEfn9tatHE8KLFuaFB5oKCV+/sVLnYSnt3FNCdiDIKkSs9tc6ZN3
FGlfyXg+hK4jfUUk+fKyaZt/gUNQMKR0g3ukPaLZjrH7q3nLdMyPq5rCIVyc79fn
8A9KWfQjX0i79ym+Lj7CKN3PXNeG4WZ5gqg3xqRLVh+Dv5HhJq3JbwfOXrQuuYoc
GfExzKpOl7iXeTKDo+lJ7+TA2pOOq4JJiIKUR486PEae8GTjESYbkoP9WoWVgIfk
XjEd2ClP9wuu3RjRDjCDT6bBjAqCyemFLKpFfA4GLBN7fWhvptMhVrfGjaOKEA2e
/xpdaZN8TWG9N4RkKRvRrKM52cpcgF2mBsb5Zr67Vv6E2/9BFIbCI8ZteXI2yvz3
u2Pt0qd9Wk/0wibfIn68jxAp68W2QP1FefWxHO7gTihV+PpdQuIBS9bLPR4EnmXG
kVEjWRPJmxmtfLdXtIt6wfEC0RbAbg338YMD75j7dWbTYWBgiTnO1MXWAbkgXw4k
0tCEl9gxcQi4Fl5+/kQY169LqOpN3+ohN7NCH6U6hhDJYi5cSG7SSewyh8VSs9Lp
YEI+ejC4N0SOmCuVYZf6W80r3iwJ9kF2rSnvfiOPABYuyRYlPz07AcMs+SKbrDEH
173x1SQCS7Xz5d9gF2asT/fYgOmJqnmq4LWWQSoqoUJwM1phJZg/OoV+EufNNIAS
LqxmKHGAuPk2J3lvih/myearp/APBeWJ8MwANuQhrKqmC/2A70SYeoa3O819yAW1
eZ0aMacmihSYMXZiHi/SClgaeozf/DxxyJv3hPJRYwBSxWU47G+QjzYXV1Sj/xDs
EAROCriJ6UUlVsA+JqAKfIuxPqBmUXaGJ3vwNTSAw5N0bGN8RCdUXsbifRrU2EVr
YEwP/74Fgj9wqQo7JX6dE8cEYhj0Dx86BwEdbANkxhJ0+/m6Sq+zAkdBSIzh4aMF
werFMaoMh/lrQBXH3HKYEW9Uv1jHQsxJqFMK55XOfK/B6iKniiCFPh+KXOEw8mhn
X2yJMQdWiOPdxgu13EN/P7Sh+vpkuefF3RppgzbIGS1gmG96TjXrcxRWy9uMVi2T
AACaQfYmdOC9//dHlEr+MhwtIBlsmezyu7nADZu22ZLZHyHyPCsEbYPOg3YmEUtn
q0OtOdzGzUAbIjHQFuHhNUH9OS60NsTEx4umPJLtzGIGHyGHNlgYkUuCllpS1lkT
VOUNjuNZhuOi+FLvuREL7g9wRdQayFlRZ+CbgdVfxU6kBFlWO8d5EtjS/TUTVygs
Lfmo6keVsF4VAxJUR7Jda2fdX5iqeFoX9wgxUAJTsVa0go9EcYc8MXOSriCMg+vV
DNunk8u/lt0JkhrxXnGlIl2DsU8GUfOJ2Y1ra2LM/mLtEXd7CVC2h47fheAudvnQ
jNjW//HddL3PFqj86rX7A4tGoFKo81of95pXtPixPuxmbWY9zHYMdTUb9LunBsSB
K16Kxif1acpOoSL6UIpDoB6uFs2u127BBfpwbBrdkhLMOnxcfveWDDULpfREOfpJ
7trpJrMek8DNsSyE3822/rwqOj7hNjDlL1ZaGFbwaLvNuqPbQpgOwzGkKG9i3eNH
mwD6OITdjgQupU+pv6RpERTJckyx7JXmNx26QiFNCIX70j83Zts/hOh/anR2Wgu8
qFyqfUE+jIuoyXv9z27gdaEo1aUjHoFQUa7hyCdCIrs0OfIe5lg1sZ8qte47QWFg
ZyYQ3PQ+JBHOVdYxXrrz7h423BkNPa67/tm9bYjMGkyZkTH9/KF/8eGqpqn5cpOl
1afv1Pf0gg14Sn1Ti1O7vhk77B46RS2+YWpWrBNbmW5zsFMhg+GdJ3Y7N787enZx
8KjyOyqyIOCVpcdPoRRrR1DA8MKv3Zg+LzIkNj6LE0Mc2rT9sQEVmxV6TAijhhWB
GKH02b2huzgsKkWPj/bxpFabt9m7MFnrTyAqwtB+7i9Qrhf4x57WJznJmzlosxea
lCOCMEJcC6doFDcGwgQLFLhUP1YPrp2XNHQzGv+8ymt81umc32o3kIQF8HJCkUYl
vzLLimK5JxKW5sfyv2LG07Owjwp+jmA9UTlyN9EHX/bCPw4TCWzYgFxdp18AjVja
L3gftnDe/6QplfubvtjY5PCiEet5tvP9BgUNeNBpsRS8w8464Rgry0JklGRMdaxc
rB513ijo4UA+trhD+fxFiKXqJnwR/nTrFybO5nAjQ8R4HjrEiREnFi5tdywzN9a0
G/XmFuRXCzRpXjepJ9vFJV2MGU9XAU8TeW3ymuuxpUi/PDITOyPGLzjRQjsXehTg
XNQi57quQNRja2exRpgAoJZpQk4QdS8JB19l1Qdk7Ctru4wbTJcIEPiXoQSMADMe
jitQ8Ks522ongdliBys4tfcSeAHUE6qhC4IBqvjZlTpoidDDusF9ZubXWk1iWBt6
uyt+HSrCL+2t5bYPJVFA5mKPiT0u/dyCvWEKS8wK0wAmM5XDOGdkiESedr42bZhN
R6PHVgEPXTcMk6Hc6PBg72kSqGqqlvbBhHfJGCSgmbIaTz3N0Gt+k2/n2AECIOnm
Lp7+WB9N2zCCAt8LXF1vY9clIw+EWYDv3DowjDqaUeW/eZG3xm3mGjwckvTX00dz
DQEZcpyrw0OOj7ltQBX9u5umaJKvA9OsivqlmcIqHOdXC+9K6RAxLxdENqg4EIFf
2futBdunzv5B5ynURAY7cuPL8ZhhulTaPPNouoEnb0oABuanj6h0NzRsY/r4yPML
hAD1DHQP23VqkUijQx7YqFhKoCw9x743+nsRBMtxMotxpzg3+/uQOzrYxU4ahG9Z
HBP3E6y3PCEVWEOv6VvBwpqUCzeNSnN6GKECDMGfk7STPywMW9M1MV5Uv+qTLTY1
6vtBFOm9KxO9vk+WLVW54GyuRR+0PqiJEL0kqn9ZYFagnKr7PMhsCD5oY5zEgxdp
lZ2S96m1TpgbzIliE+HLH7z+k+qjC3TrhVpepIu4VZnw5doIkacWLxAyU8FexPoH
jGE6mIgyFDkDs+BvY9HxwDzr63sbG1Ryh8P0PVBWROzbczvIu6ULz71NZBFC2eAo
OyGdOwG+DG9ZwAwI3TR2j2z1W/+vylWv/DHSxyENOBCFXvgDfDKq2iXByIzqpDGY
0yrRTEtVAn/u6JE/c6GVugLHeuiEkZ0gWP94gr/Mfe53w2JmEcRcrb67lF3jhQyN
36YBgoW71WKPp5Z1CJTq539kOmMmoqrH31GYYS7BrT/8CbFDI1s871z+n8NIFUEn
REpJyT0EPq+efd9ffNuI4ddE/+5zrTPnxH6IQP9eU64xGYzYkvJggh4XJTc+Hxr9
ZDprw7pdURAri3jL843QTxim46CD54j+ZE3sazIXHDqAPeLbtkdqo9T4x5Hzo3NT
oNr6o/f7M93Ius7Yw70exxQE3u154j7JXsGggNXZouyuO2mp6wH79C0Ae6zpJ6aR
/VNHh5VHicxSO9WICmEoZhhSi6qLUQDSBo1bybhcOIZlzQvL7NZlfzuJTMsr2n5a
pGcAqm+PixkvyhETeYQx5PXcFlxnVqyguXMam6sqMVqwthBA88E5MMgECkJ/XieT
XQbZOXibMGbXv7bNb08pawtL4W+1juXp67LBbJe3YPPMPaYrIHfPPiS274PFHjFV
geiKS9Y7o1xMJ+VGP6Z6a1Ubhv155B18MnyHHPEfR4X1FLCL4LgE08ZsNv8xA+jT
kDiqOK6lc6/9q/VPOfnFUdVSwjvGql4jzzkCfymSg604IEnaZ24vRuQAsnGUnuLg
bPrqUMCVa1rn8xwFAYSYl7qE1E6lPUY/A7F659g3nwiQnt/XqsFjKQ01hf7zLIXf
dxQBytPOes8LikIqjgQxriQI+5yCEwPT2IvBxeuwAFGlY9+q/WHA1ybfvhjLvgG3
4K2UiNlVRoye8yhz+gUQhKaVIITKA3LsgxoLIp1MHSjhnsmFHMM0vDbn0W04twKr
aJ6vUVLB+CGryr1K2z3s2po6aK53qiAw3QL9/bgKc51YLLxbstyrvYMI+av7jxMp
yfzET9VuSOljOrQHPBpyvBuX2jSVS7HYjsWP6qEnpXFzKdtjlgUXTbRS4M94ozB1
Z2VlRXoB9nm19D8oHgXTv3qyQIBSvo+q0v9FtfQlRbiy88csgj6s74Uh630cGME9
TbDA6VBaP2wbimooBNgy0o3nLrSzt2PSsuV/iYfXUuVgy8MMPHVqfMrmcMH00KWd
BavvKLZTW4nirdM9x+l6je0oKcGrB1tvqX1OKE7DgAS+8qDYelf6Q/uvRBrJFQYs
kcD/N5MDQPiCkGETHp6V7yhpGUdPJV5L+8OflsGC73Y3GmiYsU7Un898rC9Sp1aA
PXLRvoR+//TbxS3Pld082q6/iLDfTeKIRw/3O7FKonwqNpXxqSzF0xmw3GutAFjc
q2rdyQCrb783p0+n4ul6af4goack2BYbgAAXJts8EDUyF3Sb5ifqhZsDiLdNb0xg
znT2RZRxZvZg4z5tqLtv1fdP08bqLOzrtKpV3hx7KpyoYKYsDZSz8Ej+8ZkHuhCe
4D1ap8rS0U+jxFENB67pFOpSk+y9NXnZKY+857S4Uqo5knb/oUOU+9XRvYVHEPDI
gC6DnppfRAHRuCBf1aYZuLoIpxyLC9CXxqzKBmcNbHseXdai/BlmKGNboWaaMyC5
o7b332iB431hTQvVIYtgPp3wlQ/Ohlo5YCdfiAmEud9j7QLI5gcKAGECzdUjJrCP
kShjHoihXgxgcIxII0NK79l06VLdkMJ4mCcs53xOf6cmr0N+Wl3LrXuInURGh4QI
yczeTEasEin3vB92pPdje6XN4JCNcfMHZIndH78I+2udYpUtqU/iKbtFj9EoZlUR
IxfHXRY7AhmI03glJ8KWyqQU2yCJT51dsTDuK1cd4wHbHZjxcs1kLKtl/vLQ1vTU
OPJ0+xa5VR4gc9oualzWepJkNEdVRaa1bxHlMhCoWmCxQT2SYWKx+8GnpcGevOMo
isxLCzmNJDWp7wl7R9SMwM/lnMotZtKlai9F6UTmCn90jQiKDOUWhVbcI1bkCSAC
J1lh8+meYKuKuoI8Y4r9Dq4QOVrVBssM/C7T5MK+IppFUtCJ6uxjG+8gHyOyDrls
ZuXqbjfOjzw/PpqvjEc4lEwJgyZooHz81tA7nEOTZLrcB1kwVDEBGqiTqmAehLi/
oAhq0Rp23Zk3X9xtScWAKfv5ncURNxaO/zQeISnLpdVQN2cNkShLZ/mXuO1VasdZ
xhCSSzEjPiPEpowhCD3Ewy0L1C1/vYHa2a8PgCRd6Kg332oQZfuR1ff64t0fFbUK
NTFOFma3MNs30oi33UOEecwGJX8FiV3EExlbndHtIXEXLWx4b2C0SbVvu8Vv6p9X
fQ6dtwORLv6tBDRTxPZcJttRXZrdtn/LNzEaGi8ySmXA0fuk734A/FrdSJfo4Dlw
W6HBK2X6Fb4D1+A1L6lokiW2JkZIb7EJdyUkxkb0K4DjAvzG0VRd1k4whUskBna7
R+CCTLVIZ0QUlYaZuYgGkSdNndDGcRkA+AFCst35JfyHlbXT0CZ8HBoxHcQBWoYO
s/pz9zDs6arxAJ1WZVGKtP3lbY3J5CKlIuNm1cNsBDOmTxHT2OOjuy3O7i+ZjlHv
p+jP+fQ3msjgYaOCH+T5Ehrif9eoGyxd3hIzyA/XAecRz1qkPA1wSGDjcl3XBYnx
nnA75b09dNUuTV5iUgNX+gloIxpwkz/z6P6NAAgsory8GuR4csFMbCywHDiU7Osu
uXmxHiPISpuYrKJHAVgwcBseIXVR9pzV5n511vofGvgSeKJpthdg1ychbhOfsf5l
aoF0eX4YuywSdX2bBk8Ja0wwS7vYUKI6uk0403RrSd9N7vouwh4UXzS1+h+txeLD
Fcl8GvI4apgOyqEg6bHu59mGdmRiT/WwNDckBYFeErr9HOWVoMTEYPnB7Fl56t3G
BFM56zp02K2PPZpHRnvbkR1SdWhXlrAJjKzMByBZ3d4clFQyVPRLdGhpX0epiGWb
fqVfJv+xwHQOT+rTuuZ+nmVAXRKEzH7sOYMlHfNRlXf783fqlJha7V5g5kPCo1+W
NVvyv+vUy8YshS2Dn3xQrWDBAukT1m0T+s6iubsv5Vh9DwxNQBcsxEeHGbmwuGjC
scArLwHxNaIVuoy5WDCxzVHMpN+T7E8dSG8Bs8x4tmbgrRJWwB1AOYYzoRncefCE
LvO2l5mK68Ad2R2XI18fNEfMDBJae8Sp1JhzCjapjftcHkLGhUfCahNNtOmr4vEZ
q2zIcdN6EXx0gW6rsWZuDsBtDCeUTlflU1p7w8wRLuvagGl3646n2nYZgjf1CjEF
VxUr0N1h/a2toiapzlRmasOxDKCh5C5gsRCGIINzFVSvS4ownAmtkUqSK3lIPwJy
MXqb9ugQMcAiPJu/r0NXCudCEB05DjOy7DQjZoxald6OKrUaZnDXoop6I9Mr3RIT
yR/QqgCq5BUCqvl2dSp4DISnlmafZQd4FhroSYKPUK35+RC7gnWbEiMS9MEIBgt+
utRHwBJoSt2+RtKgOUCL/Hfbt3azg2w2eqQ0CngVdaqh5YW1//s0KUObfe2bLS74
DUeqtP/5b7a4Vb7+06X9jQxkM6W0tC1eHU+xcSB6tSzh3+U8b1bV/kO9fr1ToIyD
Qn896sqI1475IYJbP6PxAvZHkqhJd7hJ7YfpBNig+SbVc0jGPPnQ70kIV2p1IhO/
2bPtDktYjQQWMzl7397uU8xjJoUYVUXoLjOsGO0j+VL/9DSwYmoawkY6E0clpQLX
Vy50owGDgG+qgW5Q6ho2meP2iDZEg7djOMis5GCkWL8mpxIzxCas5vBRGw8Vvmhz
E3Bc8NJjlpE9Cr4ob0U/TFnGzx6yuRQ+SJrJ32zDlC8q0tHCXAHLeUCnk1RpNDuh
fmh0+DibfQuLXNeARCKYiiAXN3eMq0xwSnZbDcWRs4gAnwgSHJqACOcfrzwVKvzU
F36YJ23/7QXsZjmJzBP71pqpjCll5LHhzvVloWPla2AV8uciu/C8KLlre/hHOlj/
cAITIHyVVxqduuINNOvAcO7P8j2YaU5zpb3HnSQcnXJ1E5VaVOF6ah6NRH4XONJv
GKx6e9wpx/EvGXpp6Ks9JHCJcPikb68jY38lSG/EedEOHQGtTL0GDGvGf86ARDJa
liYXuOrth7qminAXy51ZI32vSOJuIzhHcWAy0l/pwjie0KXfCxTGnc3GuGdAgXYi
dfZZGEUkOAxPcquALDmQIWVAbrPL44NMAFtb4B3zo+seie2VUSgltSWC5OM5gXs6
jglaJMouUiIuomRcoBvut4Ili9I1ZtlfOtvJsTbcMPJK2ZbCzw5fUJnTkURA8H3k
IvDa0ZSDRiosGrPVcagzHH/zHA0YUBnYEPZ7Q6vs1A28QbSj3M4kJjdCVfW65NwZ
Et3gQdGEosEG6asIWyMxoSzp6uFTCr5MjIEJ4X53g/RXIRI6eWH21ATQfhSup9Yy
2K3RUKBKXe8/dh8zZQtJ0oI1Hs9PI33Wvpxa16uIynajhpxscll/U1p36UeinXyZ
30Xzj280aQEL7m+XgSNfN7+hCRhROxtSKjFCz3GVDxVo/T7cqA2DPGjQ5aSY6nbH
Hcc0EuD5WHl8c1tNlDbhrI5kn8sQ8YptrDlON1G3qN2552V5menp1lTKA51ke16j
dDOufWbGVFty0VZczRbp3+mdBko9QumaekqVtUgChsDbUntZBAQx9fGygmtcqp23
E7im5rWG3WF34xdyXJii9TJDRWmSQ6zuyBZhkGP5oyqqfCQwSJxbnlj4NAHgueKQ
WcgF5S8Iz0uFiwP2cC0QVAEv/NAFA3TmA5BRrMWP1Hl1cbYOKU+vzGIm1jNUwbKB
lAP8r3NecfuD6Zc1Nub5eRuaaRtPtVaHG6sFY8rgn2Y1VPjt8SZYnGTpK5cSMz7V
C6WRUgI52Sm+KItCQDs4HdIEQuNDDJk29NbYDEYYJLBZCGcvcmGnA/gPMZNOUBD/
M5qYr+iAPnWQCE1hHo12VZUnjln8AtAIvRsI13cdddo+y8yO2GSBbY4j4dWnYivT
eITBN6xztuHj/cJfwGm7wrxnRq485+zyUOeqDtphR4KadrxACqy0zDfrTNDhxYCK
DDcNqkr13MlPyKXtz69cpr4+dht5bvn4GuRLT6VOuDRelOeH/4nYS0snxgubkPLl
fTRp8jtVrlXvjU+6dvEFR2zLG3E4+8tlPRh12mlCT901fR+9oGfIG4gP9Wdzpzff
jfn5rpFCNWB7vS0JeGsmuRwIOsola41YGSyXoOM7RrtZ34aroBAeln2pOlobvhrx
3DEtuIBL9kCp6aWa7eM9CQ5MCwHPRdyHzacAc7PUOcIyElb5e0pQ+2A2EwbTwQUR
tcyeAjGWuts7p2w0YAbcvnQOcbiTyFCvJ133I5ah1hJkTBYG0lDUCsjs2qKW8twI
OR42yskrzOhq47yLzYK/vnzQeGRGgf4Ag8Qhwa/GRzxYXN6UZDbj1mA7rOJ3NlRP
Kz/gNzfJksR35/LShr/832nPnwBLlaiOo8or0w22E0F8uAn1jS2cOubUhlSlegVg
9wD0oW6tnBWZ9cy3ZM20exb5bWrsEqa94QX+v/wKLuCu6SdeFxBsFJmlSTeeXoq1
nreyMTWojt56HtIngCjoHnXeECbEfhrbb0djW6wi/vBiXYReWsIowpTEpli0lmPc
6MQGr0W7Qsg6+IW/r1LJkMUoGB+oUKTXaRxK+I0ZiievXXCiap8c3GzCH8XdCdaw
9MxGcLvTa9XAzDnobHmv9sMroeke1nPYazTBmvWhZ9n6NzyHH9RBhE9vIkwbfehe
5sASiTL4ns549lIk9JUytY08W0XgmnBAxgsQfq6pMdFoCQxBZNWFs8ezmUrfV/Fu
iD1UjCtSwZH4ExEXS/PQvver8PIQfkYhDeZX5SKP34H12thzwC8V0+oNL/h5OOWF
4+rnN9S+CBrEEPL9L91CDAA/DepSd7seZGgCq//nBLB3F/qolONDa00KYm7lShLy
G23fNQndrRwQxK0PSv6AZiMU1J4m0sf+Vo6ixfsmsraEHDnfu/Gos1kpF5Sbu1mc
vI/FXKpN14RnJAUMjfj7WRjVEP/5CLQz/m/Yjk32VnXsDfiU3+bQLF4y13TlXk8n
LDPfnD2kY/IQQsMPfeoHN9yW87NXoA8mmna8X0EVSN/qgDDe5FnjfIv93t9FEHyZ
2OBuqz5FHoSI6am3ZIzmK3fv04DzSoork2/vJ5uz96TME/SmqJYoA7TB7MNMqQCm
WPxgt11u4wF5ROZ6bBUbCInUR8qNSubPZpgYehfHKOIgoYfDQsySqNOOZH286Q/y
9aELITqmnGR9iss/3qBs4Ni2vjWHIZ+OOGY6Bht22D1+1QglC4I2mh/Z3E6M4RiO
tiBR48PQmGhCry07Rz3rXU5RdjqkXIxPFZjVInZaERCiEwTWJBPxe1mXDoxQ803b
G1YWBU0YL0xaf+gTLyjibG5BP1xcjVA3+g8lT6qoTeSe3/E3m+1euimkcr+1b4PX
WJItL4sssGbvt+WhC2igcFo77w0swLTIjxn1N6SoQbZVVFizyA4d+f8dLX6LH8YI
elXwTTDAPsuvfUvM0LHCtfUyeavbpC3ueTPe5JLohXt7i3wckg721ZljBJgHrFb3
esKDK+wHQIITzMbE4ilh90u9Nmqdxa71OIhzBmDxNZGQ+/vTKevGpkCHuoQ5dCQF
I7hlwmB1NdTijZyswp5Md+77wh/jGx5up/i/dS9/cNHM9GQ1/Z6uiZe+R46ZeQlR
8AFdcB7XCr+BVqp6zh9vpwbNLabefX+2hDpaQc4hXgJMNzZO6vvFptc57nLI2YoZ
Fp3iCWbcBu6YedQ0G/+/ej2CnyWHhOv/aHd/mjeqFKoR3b7HpHLFG/EqmDaWQoVJ
o1ewSvWphcICiZ0DDLbw397uCGhOfyEW5RFpBnGYyugwB9Ya8fPMJ0Rd5xAv9I+l
twHwYHmy0iyseUB+DgD8v3mYOPWhKbmzcuJpBRnVT8Q2iYb1FvvceYZxzSC5SSYb
GmMopQY5bpwG3RcElG2vf/63FXoXAFycm8p23udcLVghL9qZSiK6uZvtG4igm4lp
wgA3yPBlo8Q7NUvqjVXCzNIOCgh3Ow4i/vW4+6NualljUU9WyrdgUe153JYoRCyf
6HJyFUQGAtVm1U3vMvqVND0/lTU50ryMfOc7LS8fy/EeLncP6QwnOAiWrCXyQ7En
kzxdvm3a67nrGlGhkGMkM/Oitr46WipUbjIR9tcP+oivnlM3qK4C29LNOH9VxrbJ
oPCat4wQOe5OqeP1GJzpp6pOKnK6i40p+vHWsuJLDK2iJzps+ni27tntZQEQLRR0
tec5q0t2CP/deicnA4w+pgLEISHthbEOLSplUWQd7mWxsQ8/HTXduAEZEpk5Yz1i
/WTbohAwPlxUJe8VkS7qJ2UJpqCublBrB2nRoKmMG1fSW+MJLGckhrav9aV1gVER
Doa3lFMMifMSfhyDSIrPuj41YiLEoKqgcX56uHAgJv7mM/a0ZO8loXOyCl0d+flX
wBOSRi+RvE4kuuwL+U7bsy75llO8RQydbAsc9/iwOxnlh5srtZTpSRgHFK4UGAD5
bxZp+Ndxnz/3kxsHa5s+6bzar4UWHEZXgksyfUicyY0AOgmLEBUzRc3wsYR/LwdG
LFrnItUslqVMUu6uumIV6aLyx0MU/E3sOsf9I6Dk7AfD8iOxtmkSthp4h92nOaMm
uQ3OsZRRfu88aiPrTHYmGicJcbcsCIa0sFPYu/gEN7xqBe8HQLLSwYEmQOhIEldq
FE/PEKRqUXq9KsPIsGpVPWCxEZWSwWp4caqzg54PXHnHHRwnZMyXhj6CmOaPSz5b
tKUWtSG0EuALfcbC5NuX6YvMRboHU4I3rDQSIt7KiHINfrB44zu4uXMeHBrV+iwo
6tWTAUJTqOD4wLYBfwsKaPcOnGeMnDL3Uc2I4+fwI6Tn5Us+gdK94UYVFlKaKMcK
lYZe1b6xIGSds8ChpzhEHTCZybweSSUs3AN0iI/2MJM/V1YF7926ruGHFCdyK3Zo
GMB3FDDbPp9GU8l4TN+7L20wzLhl3VYpDBaus3oC24+R1o/xBqHcEqmpkO3zs+6a
6SvmkKgdv301xXdGCbe9CxWni37hDM+ilhbEWa7ZzP1wZYad8DB+MTxarIGoJlqz
7MRa8Py0rim4SPjpYGfFANkN1qDF/q9v5iUwFkOiVQfiJVGm2OfmO7+Qku8IKOcZ
k0Vqf9nJe4OtjlYM5x0geP0Efm3lRkQVtKoGLMtwbyjbPRsfeXVcYkkSYZ9Vax2d
gWui6rcn7z1+cSB1bzrJrN/4uph7WUn5zcLujQ3YcNQ2BCausS5dAm76cj/iWBBx
ne8qR2nzrYLvspN5WutSV/5pljtzozPy7srfRBuKicksNENzaPsJAMydinD/Wqeu
rVRZ8fc0oLENclK0F4nhDBT3lAewSq4nRwpIql7ijOzvdZ4BAWcFNFSzAW5Cj7tK
n/qwneaVieBV5sLCN+apco4BlrsGxU8O8IIBb7rHpHyPjULd5hdsVu5MGmdPXJyR
KVgngv4fb6UeSGhSfbxyU139yHGg00HOrIO5A7/qImJTq5gDNVRVUIN1YVMiAnQE
JHzRRUX5kbROY7aA/6nfid0/D23pH4J40XPyezc597Cp9KBDtGy4Wufxe22QHYf5
bHNwP0DxLg9X/7nsARlk2/GSz6wNO8lYWc7pPe4TlUfDyf9iSXVsEELD4S8DtYFJ
4nS1lbmV+okHFEfwfBhdPeyFDFQm4rrmteGFbIINVXd+WMucGBb0A07Wbbkimdn2
0pAWfv442k74TuWV241gBCrDqKIcFRaJoq6f0Q/dUvRyxX5XjAIEzl/BTZO1dDZX
cITkYPriSrfr1aImH7MR+dr5ywVylBTXIB4Nr8NWuBElNLWJIWuki7TgEa3UNBoI
doDFaHMNbC4Wi+u27x30pbQ0IaOHRyLJKccOwo/78fuEmI7yOeGqdUHAtpekhCiu
6fKQK7RonpupIbvftyfj7GyV9Iqj+qTc0WJx6k+Ug20H8zXxQ8jEazB4jlYRosjc
gGzbLrRkaOoo5XCfnmYcbVmeUl6g6KCld0lv5UDTqPzLBU4yJcFGQZ81sgeNXtTb
82kxFdGZRaz/ZHjJfoX3qdPN8K2SE+BU2vQT/SEABdpnwyk05WW0B9SgJ9lncl4w
brW2B+yWvKAkCNa4wDiedI/GyZ1i5AGywxFpkZZjSKdAIGR9u0YmygUstJZ7wzQY
9kf5zEFnkwYwaQ38cLDHYEWmX5nzY+53Lwb/x1F4/rZVKtlAqWomRx4DMbFxs/DC
ylK3nqPD/zF2tkTqI/tD5LLg/q8BQRHCaQlQRe64h6mWjmeuBdedim944EaTeaYg
WCC4+Dkv9XreAZWAPt/IkNCkLCrU9d8GpwGiyMKRXA0rfwlAOLIkOQ1KeHYhQeCH
ec1LyXkwyE9c0Y0Pmz9B3bvztCGHru/1e9caPYyy9JiuzIjm3zs2Kq8JiHaEOafb
ha03kWSVcn/NkehUmxoCyz6BzayM3qt9CG6g1ZCukjBP5pno1gDEUI6cvmNiEKn5
yxiXLEtY7YXIMWednJpgRzP2LYKS9d3JXmYWl0eJPsGBrP9NDlO6o+1Q5oOteSdW
22mRX8217LgvS7Ci0RXw79DB6uq5uPHLW3fnoDv8qrz3UmOrb4L4musayWEe/8pn
xJfuVz9IcnoxMqjlj5RCn+IC/5qATiAcJp49qDyMwDCUXTG4TqyrM68Uo+wEVPBO
vySNiajqtMFkUAaihAGwqjNMIHJ98AvnYsIGH0b4uhxDu+1gXWYzmXpQ1046Mbmh
+M8CKHR/VsruyHVhCV+vVh1cR8BNy8AUm0wpuMLcHf/WnTChehxLQ0EKw0gu2qIc
a7btN7GVoeIsvfONW/M6pE9T6c1tjBOYOzU9V6GhI4zkXNHztZFrVO3BhZ6Mb8uZ
6ynVKj8UtKg+Y8kKAwLR1rEgqWdHDm6eXV8bhv/POeS8om3hfJsrMoe4lUxdifd+
6DO2g3oP1O3ycdBq/qBsag2aur6GLlwS4Dr+l4KieI92TB0w+eXfPAmREW1ZOZhW
FUmPQMEiHJGAcg4/PLf2wUQdGGE01xrQvP0MO9Pm7Plwz0vhaNesvEA/TASHeBu/
+Ufornbn9mRd/WZ/6dREgIQ7EoZnFEMerF88BUa++vaRdJp6QIu8BB5o6IROmkIu
v+Ll6VO007Pe7upSaUWrf1GPX4AS6mO7PSsv3kqW3I4BBrknFnoyQ6hvo9EhF7Tp
k+R3Mb18Dp5+VU6nOEOpdEBlZ7JsBhp0ym+t8UiQNOVAApOhIgACU8hrd3w9gzFI
2JUqoOWblFyTrBLXWEVWRD2seE0UaWOIJ8jhLZ24ae6JQPs6/ZJvFH5inmCXO+qs
7KyclUVbPfGkpN0vMJXCmrOG3cMWsGCmB2SvLz4zZ4XA+w10nnPaRtDX+6zgwR1/
WYatIDxj4/WINUvb/HertjX8M3iFXEcfg2yIK62j370v9gwvx/7ICGty8KyEjuIQ
jyCPmJzFj289Bh7Vvrr/kWIH7JjovlEt4Mexy0200XYIFy2NvAuACYGFxz5QoW2Y
HPSPwCYrbi0vCKp75pwkFMVo8Q763Pmx7ql71w1mpdUzlCeFR0mw0dJsDP6ihU5y
yQiatm/HplITql7V5mhAeBcaXo3syntV+3Ok2sd8eUAISt2qrIe6COg/pXi8UgYh
ur5e4ZUz2dSAeJGvrJMK1Doa+FlVJ4a2MFd2N4wVhOxqcX6GXQEKXvla7lzKtX+w
XHgFaacXfew5W65+ux8V32Th/ofcrrfvKmGXiqcsdBr/e5QYQsL6JLE4wt6/UVn4
GJL4TL4s3hbYyrPt8/JzS2/8LgtW4M186wTo/JskCfxk7U4DFrBnXcOnCHJ5bhJr
XzmVnpPr06hYuxzBwhkEcYPMQAHRI9Xrv6vbX6oyh+Scwp/lMx9+FHm6tIwBxgLC
SjrBuPStSNOwBF0ZxuNY3nTYa0EYw9SlqP4JxS95kZJ8GmjEOQWMUCSOqtk3XK/+
xi8NCZwKAWHSFGHMLGIpbhms0cRG1qJ6QexwfBHMM02bCXEOy5WazDcUhie3voCd
mUnyLjGArYWUhor9K8yW/vS7cKTm2nAGVb2d33lg7U/l6ZcF+c6vNFBxtk/tZbJc
60Zqy9qU42R+QUM39Q0ChRahQ6BAixMguuvCaDBPALSD9VE5gIgRMzmRJ5Wvnve6
UOwcpT2zdZjb4cjVixfX4enTtgoOmUsIZPs6I5OGO8MX5nXjuMu4IjHPYudJQ7DP
nQxnuwsX8v4LAJ+JqYdXL38bhrs98W33J7kQigFfM5Y8Lzgn5C1Pia96vadtJlwE
pD7y6Bb/LPcBerRrp6u1KxdIJdg+VeODMOgFQVvn7v8ga6RBwo6Ly8tbOrilkJEV
CJN7GDuqI/YJOtaK+cJ37UFDZLuuVG4OFwovkkfb/q0elz2s6Xn4OBXmHTrzDsen
hOhLB7Q8KwArQvIIoA0H4BBRLGEEaBasQY8/Hjwg36l+K/oq48ZpDYuokCK82cy1
hqbZIhB3QiZWqhUIlXuHFI4DfoRmwSo9xQjP3uekuGmSqG7nosYmge/VXWMORDbp
1t4GxXBz7JmJq1sb353L7Cm6i5543Nhrlg8HLmymSlHwzKrpjQhfri0AgPmwSGGa
VhUxYa3ChC0vhI059Ta7m6rkJKHKbiifnonxS5sYAo0OEgMAUaq3LaP8EzTpoPto
BPuX8QcvwJU1huFQ1oxyvclUeUNIHyUuzMByDiXmUmSNpWp7jL+fMCLOwnGGlycO
Jxv3rRk6cz5jOPoz43A9hN4GO1zzGE2oTj3WL/o3ZdHnvuBpCwn/0ovAOLXAOxK7
mrSCPPT8YMuFcMCFWauYWC8GXvbxHT2/yzq3TwSlG29Rsd6C4MKUZlY5/6jrVNOz
dW6gV7z6XU9UVaGz4RIQBUHfwLd6rBW/iC6RUlBQn9zlOG9UHa7ALNm3YyPh+Ra2
AZ1DaYXEfuA/H6s/Al3VQjETaTV/xTeRWioMaHIirNXSPczm580FGkNzmidWUin7
lmLcM1Mu0wWacCU+x6fA+6jola0JlvO2z5eoAekgBAhPqgKBT6YPOMbJcIYfxpT1
JRl0XbQYYUuhEyO2OTFbniUO2D1BEwVAqOfZFRmF7Sx1vc0fr3xFSrwrAWWJyFfP
nRiQiCdWx7SiXwtsM9NrY21Zt8wojW50pN1pDSno7sdZ/HftDA8WULfChW4w/CIq
ieBwg1NCygc2txyYLNnfYv04tz5YmABecnplgZNT0d0imQYN0oAeEF0W6W1iafzZ
CncNNnz6brluccUgT88uBvObP+BKPhZnBl+EvUjifmGplKH/RbayFgZt9lM7rDo+
vX9E53PcTJ69fw6dRDlVLNd63Sd+urXRZaSHhTtnUvaH7q1GzU4J/jNe4KhR0TFI
L/atB/uauteraShps5Ru4VyUNhnIRAnbivnSe6ntl8ur65ouIM7XQzIgkuSWYrHr
IXLkVGq6R4f8fpP2fyjbfmcUIMS2LwJxUiXejoEj3T2p7bxPUnXXHlOUFMbumT4Z
D6p8qrvoEoJrtNRVIHXyY3JiF7dAhquc4jLJRTVW2AEYjg2DlQ9h80PX1AdIb1ZY
3drxGmegGleEGnJsYbpVKFtV6KO/WEax0RSC0ygnuxAJkELSMctSzv6m5ceG7FZA
O83Ktej1ykQEwolB8q30ZpZkBPmbxB8HPZrBcu5Ncys+8cc06hd4/7TG30r4SF6N
dT54nAoKwMBVca7xxwwgTknpeG+ZQsxobHQWfBiLje7qyOyLofJERSbzcD6byLKb
lgQmvohhT/hWOQ31AFG+nsPYf/YlX6rBKwtt63dWZC1N/Q6ILJ90dq6KUfrW+D1K
f9ZjG9mR0cw5HEppY0sp3Kf/tAinWsiaM4zFHOJ93fuMDLBK0+ZHh/tRe4K5goVI
ErdpNFRgQnw4zqwZ6C1vWDtNQgQLIwjX+cKLHDBddeMyoPqd4I5ow1QIg1xbEYhc
zZnyW9ohqWst4wfryVEWntfi2oLpCs1vyEQ5U6XkgIvFgdL/xXF49ZgGTC8TVK2E
4OSyuDs2ZIt1F9i9hWTUFcPGJyrfvb3MFBfYpLb9XXaWM9DBNCN6TNFO0Kq3Oeaf
Vwvnvr7N/7yWEkTDPbOMqta3s0WmBteLsxycqe+v9f2SpubXoMxGqU7aHZpGcjpP
cnWhea1TDR92Y8L0parDEIgjGW88ZrbFgcOibZUZoEgYatDHS/aXBt6It4ydSmAv
MehzhhBWZpeuw/EU+MEhUsAvWBpVfvpmIpgtj40NPSizGrOc+urVRpsKEPPJx+g/
pH4i7zv+9rxUCNpgLPcArHAvmibYEC9iyNE/MjM75fYe5Mzhl/TAxBZLg+YaPake
Nn1+9xSp1fhkeZ62Ni4KGdvdoqTvtoek3Pz0/bZ6vc7NCNcKioTKA0NZqLONC7XQ
LxtT/r9s5xodSJF8gXqynKOzXFUsVZH+wW/jeKuS9mqfnlEBWr9YaBLrx/mlb71R
6lLYS3NcFm/+xyjJDQ4UhGScKetBJSVyKm7/EAnrwlIEp6Zq75rczwbsMPM9+MP/
//t044vbiTTbEeHtbG4jALjopsHzhDjq63QOF5rT55cm/2c20VFPblMQeZJkYexm
Q6NHi40meyxg0KY9jbq3B3Vic6OmcdAifGsouHyLhjyNmwM5tDCU3BNxKLVVND36
EAiZHDhXHPsVha6MZhtljFuZAEvYichenCHiDfWzErR60BIUQVahIataV93o2mxp
3TjoxOLlKCMqM3mDA83KzGOwAIb+O0M1xHsmlyTyqQejmYCheJrmVT0KOK/R0xqz
64C4fMvK1yI+0uexenx6pYN+7kwQBisMU9CuvP/1nYbLvCdWeFvk4A0a5r5YkHLc
CcmA1A04OKPXRNu9QtR1GIILFRNdGk3fxx5qdCfsQZZGrKt9aXbAWfOKeIofzMVM
DOG8GSSeE9LrMqwnnGLEO/FCCOWeJUiICTgNTuqgJgbS4zcLL1jJ2ppHKofJVers
3C829iBVQjVx3eiRUsqbm+VhNHHYP2TR25CB0/8JEncQvGCmS2z9fiq61r/YFv04
oSivkW3TNrSl7hcSSt1z8POfkr7k6BmTRpfNox2V8ZQtfgomy8nvJH33u/aGR3h9
/nejsHkOMuxsrCPvrqhyoUPczJce7UO5/xq7yNDv9Po48krWDGDG0NK95sogNJNb
eD2J7qFvoNLsK9pCA4OP9mHlC3WEbYuwj3BF582Ymqeo94IksnpE09hBBbBCvJMB
pqMhOXzq9yGZrPFRDxGLgv8takhyW+YxMIqQdjMVYt0DD4WRp8DJj0E+2GiJkzUE
fnoX3WPRw9NL4NjXCGlet9SLgawCGsqkN/GzXKlSJPyiJJTL7EmOEBq2Zm/EnxxT
xQIU3VE8QZnyzaEAJSnibe1JFfdYJjrLXHvYCCLP85LR8oizRStbOYAbslESZ2au
SyXPt9MvnYNpz9VSP+aTk2nXG9cTs8Hw5oRcJF1A5Wsxjd7YgeluzCuXN/QRicGh
tEzibsQ+IB4cWJAI+7Vli9Fj6dtBUw2MyZsL61BG1nby6MtlggRax6cfgUXxTqMT
iWM53ElKVyQ1Yba5TRfe4d2OJi2zreZ4sl6S/6dMK20IuzE7JC7dlU77Yzb0em17
i7vB69qoGXrKu/G1pM0otK9ELggYoIQpoAXiMr1mjjySufEG+AN89r0nz5biD4zJ
lK+4F6B7jObuaJVxN2h9xX7tW0uRzxf7G+Q5XJOZVOQJr97v0w/YW1PR3VCpJeqa
VXCz0ukgN5nF2wgXjhBrVIIa0FWZshRwru6vURX2eLrOucYu5LtQYSulccKMHt91
/8lhr8/tRzgc7vPAAyMiqFam9rHmuD592ydrUxgvH7Y0i+XpQSd/ZpAa5T9BCyNd
LgriBr8S/0SDbD2OYJwZX0oqHaRP4o2mrJ1w24kGTuThcz0Wj2voX0U5nzv709YU
55RznKCF1nRlwWpOY7pXgseOEpo4G7hjvs+6fJO6+mlkzBLcQ1/nDEPNq1j+BO49
zNy007Zp6pD4tYlsDpk+RfACbc7qB64EX6AWq+XA7Rl1mMlCw6BzMJcrvjKWu9Vt
9Q6ZYn/iCQNt1lI9xuKCg4vtoq+yVdX/DHasmpLb42aev3ub3yG3osoR7g/wSUhr
VFrmu+MpcLTMZfVjifOZ1Ufg2UplGqqcwZeopxV5jcSAyq8MooDpLmzJ6vwK9W/w
CRgGDldHfT82IU/PRl5XWyo0LV+jUrFdCvwfwNH9SN1f48tnFmQsAhhuETLN4HsT
MJ8XDZezVlM5COkrLMxOJIH5UM2fUV6HIgI+7aTyv9qi7Moqn8y0m8A5Fxab+5uv
4mweXwZkgCJiN/5RDX3Y4DDuSeV6H4NWsnjDC/a1ULws1qwtttU/LjPB82yI9aGK
6ccYIVt/5JZGz1OP0MPsFArCCSJO3IXFq+AJzM5zXFvE+XD1fIx2l/XGGHtoI90h
sLr/sBggr1ms0WmzyLXiDlCa0OT9fsrSCsBN8oIR5omcAzFts9i9/strrHWCGTbP
OpQuS9crF00rs+NCZwy9TcA1eU/sP2t5qOh2TU1fu0fAlwsY+B3GoGCD/cdAmJn9
jLLxOFkU8RDXLbnPo6mrXeEmJkKePFFizYB1dUbfa+SWnIzCedbjJusxmEzr3Sui
cMYxlA92wIq4lLc6LzhGrIIHUxx9x7ADfQ4bMM/IwPWQFd1hybVatwd1124JuBMk
nDz46fOaY6cWqwjw/wUsbYWAF4lSDAYgmeAsCUTWzFo0XwtQ4bKWixmal3TOUXCl
Tl6syK+XO5msBv+34o+CUdMogRrAMXhkqjYxiR5fleFoGLhgMmwzNqrZQ1E0u76n
uJyi07j1rOfi0gE5gUvlQTV3AbTOs2uemesqTkJNM1sUA8CF1fFtRrVOaFhKlkUR
bheEX1nIO6c9ufhI926bM7G9oVMbEw2G9m2qYXrUVm4olgePMOCNCTMxfFLgDBUz
+QKJmNo1FqADJNSxhH2d6fLliWHyl+i+XxLLW9PpxO9CnCW5BjxuAzOim/WMzZ1q
elQVq7cqxffKCshO/Iy07Rq82kfZ3qkIsWfw2QKVTZ+G87GKxuCCGrbYqUAQQWcY
dZmJ1vN1FmF6Zmbq+BmMjK06Yg2dTowANIREPDLvYi8trcUV4DyVXJZOKvwidfn9
Le5jIQBjW/OwZXFe77Nmlv6Y9KByWj5Ifmx+EMf6L4VuAqJNmT0lzah5ER5SPg3p
EhKiqEAjJM0rDc2AmYcnQA04oWL8JP7wq2Mp5iWv2aBQzpTmseIrQMjvLzEr6/86
/k4wRczMgG9VjOvkZc0BJG2agG+H56tdWITLY6lAtIpeBinSDQBKgHutTOiww+Vp
AfCrIqF0Pl78MI5jxgnSEcGL9PR9NG1aXRSik7khUrXBfStVCytW6BvnKP/PEZRV
smBod40rHM6JdSoMeSEJ+vYvTT4R98hPNv943w6CbAZbVRPvEibevHTj3bEy94qZ
pCa2wU+p0UZTiHQak4WpfxYEKvNxh3TacNqZ/TO2gQvirBnesVnSRjj7zpD4jooU
Y1p/+yTTAdSB0O2PmhhuHdCQJBw5lZyN9yciYhMNA10dx76stVLsuYjzqhCwZmfN
/upaOyqDqgWoUuth3ZB0mRK9C4d16+ste0oX9v/02muekntRH183A2Ffcj3GktdZ
kwYOE5akXiW51id6O77yCbv8LVxvRMqrcc15uKAsyzxz+wH+tx0hMXeD48NJU1Lj
dm3Lg/O48M9o6nueolJqnyFzm5Le/gTbKW5XUlfrYZOgnLcpLJ140osSb1wsBGro
F3kAa2aq1G1b7z7kQVYpm1SVv/eBxeWtP9uV2BNWGCrNU7NtkTp6L0IYE8Sucw5N
+yKuhdwpkB/b1uLzhfcyGIJvCGupWU1C/UHEf9c9CBxi9V2p8WjHyJ5Gcl1QW7fN
HDg4k8mnYky7jYAECGTEvAYCTCigbezRyIWt4sMrhCVJ1+1Muvxcq92udfSw0bZM
7K0/kym7VF9e0AM9PJapAr8ksRpI+3vmMdmUpYytbLb2c05x86w2JygwMDORg8DU
xdEQyvXKCizyNjHrj0LeGw5EBXAx78T2rSXzKiP80ign2xPWQANAmOEl7YNYLKDh
weszyr1TMitG1epb94luYcPVbMZdnKwxGRj/7S5EGrVWvuhmkcJBT/fNRymC5CiP
SpI+O8xB7nDStfPQoA773mgfjcs9+KeHAR63Bu0F0C25UeiQK44VZeoKCDrUNq0Y
xNQ1V+jCPNrZGCkTzCgEyPSJ+ZKHXWyIcLP8VmekaanTdSDcCnsr/YROuWSVKxkj
310voeM1oHfEciGIYFjefb0i46MaVZtj06q7l0TEnZIafx04r5OcCc/pIfX3vQrW
Kn9uDbCJtrYX/Zws0Oqgnp6Q7Aqj5r09iz88EQhpP+dGF9DjxTU28uFLGW4vjoNl
bflJoGy1LqDeO08IOL73uRyOlc/9kcai7t6hc+PvmsqvhfBea4/ov4KwqpgrosCO
q4vlSzCxeBlLeyBsla+S5LvpoEcJ7TsRfyn/lATSntbincaPnHRTYMt0dKnFhK2J
UBzrrtSzqcHiL9f69ilhVmFldtwQMcF+uAR4Z2D0Mgm8KzhU2vyVIy3sx2+S00LQ
CvMUKB8PJZUw2pu1m0EvHs+9GM0LhZ99gm3x7rWHatwFIfKaOl3fXlUuYLa0HeSY
XhPzQV29QbPEIxc6O2xFfvzB+7ibesCYf8NpsCs6fDMKmZe2/nPeGmWDZCLwiDE3
VQiJ6pdhunUiUzp4S4+lD7zrxyOqHgaXZVOJMBqyH1+atlEUWgi9TsLAzjJrdEeN
a/f8OQ2o8jjh32bHmKoQiup78iXIubZv/YgbYEm2I2ziBtD8F4EDEtAztwS1cg2b
couGrogVC4kniIwm7lkTz21+hs22kmiIghGwRQOYARR6dRgrfVWJL2vWnxsWtLR0
vhxkuwE7H+0V7Nn25ru/9V9iKWuYmeC4kB4fNctrIDhW8OIC5YQ6zpBTgWoVCT0C
TVJvES2+E/ojOZ2ojoFCkHWDNeSI8NyUnOWVkkWodVgVtpa3k0qilm0RKMH3J0wt
KZ9gan3yuLSXD9Euvsp6GwZONZEaZk9Pb9aSxhiOOzxM7uguCyP8lAsC8SwUA5zs
J3/CHNiCfcMrXZ2O6jDhLXeIslBveRKdQZbNuV6bx+w2R2wDlZDw6JoCdBsU0soz
JzkUJ96PDca7hoVKOxpEgzH9+jNL0In7xhFavo+Q39rFvpWp2CnO7hmNlP252Pan
QRdWATECZs6Sn/3tyojE+Njqf6zo1TiKX2bI0B5ewiFvlqt4rVi/VoVJnGBOoFsM
s+VyxUQ7+4deOlXvA2PTVEcOQNxUWGDrXT08c35sS2Qm0hbYGLYbzOoOgdFpmAgh
XW6h2JFjIOrJpeZAj6zeyjqaVqlOLIWWtSCWPqDJ3+Lsv/OmBbmnICmudtXuzRy2
EB7O2ADJxTApPlvurnGxIIuhVhv3rYm2IhlbmRBfjXg0wvgz/OGqwNZVnwgo2jQ4
YnEBp9JbI5JUQFUD1HgLdSMBWvfiv6QyGY5VJt5lMxbfACK/4uWY1jq+IQAO2IeS
Yd+NLfOvxcuJJXuzBh8/tuf1ua75b3EoNk4uEV+KaG59NYB24x2yKAdywkZXwM3R
kj73UMzegPEoN3gkEbrbkas72PDi80Zi00RP5kMFCxVRw4N9qinUeP+3vjVU6QWM
0CNDKzJ7EkIM9G+90pMrt5n/9zrn9rZMGr4obrh2ljUod5F3rEf2sDR6LT7eUfyI
XndK8ugg4rmTvG0dwsMbYwnJI1PSurC/mYunGHFgdaJ07Z/gSM4uN+jE8/rDfRrS
fEKp9op/zk836EriAB4mAELjeB7+oWSzYogSn+Sc9OQFDQz99dTfbAh1a/6nOUqF
xNgI34JYHS+IWNrBlZDqM7VbTxlEXdnstiHl91ZrVQStJig/1i67Lw11+bcpCDyB
18qomXleDT00mMhEc+/qtAj07IA7xmj1oWHueBBafCSxcLYoBxTFmx9urdsB7LTa
x0EEn7JjgiY1TLIJHjguyzHiQIF7pbtJGfgocjia6hC6ZSlRLnd4ewASv+FlnUfv
VddF2EZUUG6Btp/tJ8BWDYt/OqkpHWKc6BNJiOR/2N8FbPFGhzeCfFjGobaJeX5E
radUTCOAGec7IN0VH3x4mSNVUnMwuywyqh9FZhKjAosGnxjgaDY4pAFHn4T+Kgy+
b5OeI/yu1PwL3Wo/drlox7LCz6tUXBYHrj/QjwvewxR+dc9PayBfW+W821YU0oel
YKmCGGc2qojSLlNcvSYpQkik6KTYpE2kkRJiut53tBMcQNjfN6A00E/bp3Syo4PF
NulWHGasjPRfaVg58bwGmD0SvsU4VVxsbefKcDtG4h2lrzf/iJSsGMIUhrchm0aD
0m/y/SxlQock3oHOumq6bJwCrA89J8eLDXR9tSwz38fRjNbC+SehJSWnYCH2sW4K
8BdSKcGCgRQg9nA5t/BXxyvC4my6yLmIqKR6R07/QhvZ3t8i267WGgeHp3mTORrc
q0Q5sPHZE0P+Y8OASlk7sF5zbjTm+Mz87NtCpNf3auPVx/golrYvCJOJWGc2CAFL
rii+y5e/BnhPOIRSRhPvY+yVCBaCRzAUoHQ1yBr3iNSy7EPiPdfVMVU+NivKw7C6
ZrXtB7lrRE6Gom5hea8D26AoSyKw+92nixq/VPIjOpurAsJst7yHNEgI9nPpO3Bv
flpm/H2PYik1XK2cpyAKZVU1TNz9ctAcMnDRLx+BBl+kzVlr9b2fEAYYWuPyX+/V
H/X++9rwFSWBm0s/sfeY6cIqbpqpA9i4f4BPYKyvCKhmKy27x1U4h9d3VnXRt/CM
YgdpN+WS2WzbP8krzlSIgPDbYrcEmhgbqlVpoia+zky/CG6F+yDVX+Vsa894fF7h
/Q4JM2bHeycp2c+22bWMJTeQFdiMeci/4SP7Ypc5vERP14mGgVgUPNsiu5oxDn0S
pWUx+UsnWaRj17ZSkh72B7om53p/jyrkFNNWaNpfZ9TZIFOMX8aw7Q8ywZoWwhIE
HQD/UyFqJmtNHW+l/Blu/XycJm43ZNbgqjC4PfSssUqTmFCNk3HDvBRz0pXQzAwh
HlGx5+wcKlh84DdPNfxbKa2DZX9bEL6oqlUha3ZBnrRTHgls+fv6dHJQ2QztrWjf
IzM7OLPorxtKJF4dzGC1OOUH7+SptxyUtKzI1+DG6R1sy2acUW5rwSes16zJ7J+9
4OAaL0F03rOzS3FG59pCorFTtg3sZUPnJxuTsR7s/k8ixFrCANmhHsNAmoqI9Bkw
LfIXZOriUQMjFqrkfUu/+eBXngFl1DSP8q4P9gttdiLMFsgcliiW/evDCzrOEKzJ
CVf8SJp7X2kQDclujUZomakHekQMQBUKW8F9mFJA40CCBEH3jt6R7m+0pGAi6WTV
Wg3sU/JueyoARKZtC8sYVdtnPhYkCMKywiAEw4a6cJUeGegImoRRM55dloGmEnZX
E094neTTQc6dqHn17eV+kSFgzzIzvWHf3QBGZCxJz1fux9v+bX5MwcMakeNJI/Iv
iCjIaP7HXnnG8EMj07JApnvYsX1B4rm4Rmk+yQf4IJbSSGZHGn1UJDHx7Q1M0Q/9
ORDkrQpEvUpeF4pd8C0pQOlJRmD2S3WH2HxPMsPW7Axtx42YrP4RvsfrhzRxGIX3
l4UE/5mKBcl/e2/6gqDDmi1+8Dz+T60gX7TOnGFRkBdmY+PqTXZ/AaP2ALMK/7KC
afDcHowjmdOmfxnWdjcvRs3BrE5rInjPDGMLreViTouaYqVXHZEWEcoNEtN21R/x
CxpYlqMHqKuI0s5RpjgECvN57+0++axG8LLaIghIymgK4wSGn1qUUjlJQtfK8T8K
Wy5TaY6JkPxDz7TBqLY9cf2eNJ1YHGgRVOuQ2pCVM59d7TQaonm31gHsoDEkVYYJ
z6MN62tUt9Pf98Mm2Hl3pYlRTg4naKUuWbNwvi9SEqhK8vx7MmrjGsi7AjOxNupC
FEuVdaw07lYrH2zHMNAiM0NGk4aysKjEOwJa9/cPFDQzkci8fpajlRIa01TMCw3d
blhDrqzKoKhEzB+p/pakkkZQ7adqvTl+8Dkis69aL2Tr4YbbZlj4m0Y0E7irCLjK
PqPwHB/j/Xe0RD45zmnoVBSienr4EbyQMc3JFHzB/k1MqpG0dEPDEWhOLwdI26wm
Nk/pKfASKOxLokkYas3zjcBrCcn3qnR8m5IFgJE3f5NYJYuKdSve7cXjjQoUzbRA
VYUmJGw/ktOZFEG8cJ+hHNSxbZUDRmLQ+BOu6l2xVW3TPvMI6ZuW97XPRQjKMwXY
lkwyZn9OieK5kt0Of0GPLsd6gV+LlstHyfLWN3nw8UvOgCAMGP9ZyNT5y00Vux7M
CuOt0WA920k3sRDcfXYcIVzgNW8h4swKg3E4IvjkQ60RWxLlJpGX21unvYVHBmjR
p2UP6KLf02KeZ9GTidg1MFUQVZJpWdFrjnDEP8D+M9qh0l34q/IIIYzK8KgmJFW9
faFUSgqtZFr/Z1kSVtqWfg7bsHCNz9RrZhK/1Soz/f1U59nD6ZeIE5mB7t8kJLZF
Tttuc8uf8ou6EQTbVxTRl3up+/CkG6rpVVhpSmNnSLuOngsApC+3uzKJkNVx79Rl
/KGM9Yn4fxNljNvNuldOTZ+IuiO/irMAEnlGXZdgvmrVrSvdxHXvk7AFR2iHB+sW
hHJXj7X+ls1PgthyZ+x63aDn8o6sgudD2OxGH4eVtICY+UmTByMn4B/URWE05Rhm
4KIYE9eVNWpbsLms0NoHyFAlLCbpvLhPCHm/iCJ4tiOF4TcrvSS66+dxfj8vc5zb
PVKGP7rOaM5h02i4+4rFen4x64njeo0XXfH3ZeyrA4i+82B3bduJIRJtBLQAZG2q
PP3IkGyoyYVI/JTbTIlpXdLKv0KMb7zq6JayIl63zzAgMInsYEgzG5CiRpiX70pA
579KBMiMyLOXvm0AZKZ9InIsAPFqm9EjdoHzrkTrWFuZ45CEpva/qo4cD/YKlhE1
41xn9SvXZepiHzxPnptMhRnez4yZOnKUXg5xFy2VunuZXEJ+2mRvs5JpEuUpN1JT
snemE+xDACQ2ljX7ZTYCoocLNVhqAjzworoZAyG2KbL6wR09d86HZ9TUBlKeqRA5
lVfN9anBnxJfJacbM661pjQjRTkEqTN/OIeKnQ9ABeKrI9l7Pv0z/qeyS9xNYUro
nfTYveBAXcSClzVI8n3GnPecqH4FgIeKcp1qRNeXz7N/AbQdEkAPGrg9si15rdwJ
DQ/z/SThfbax/mmAH434nxOpIiuLneSphXxB2rLTJlXSqGu7BXrAYADi5fLBnrjB
I/fSuXh5afVxWl20uczoDLFVG+zspkfrCOEYRK9Ijys0p+lUcXpkif+Bfu0Ni4ZV
DD3DnbBP6wTTyOzExneiV3ggBDiYT/mc1wKG840b5/f3h9Krvomyp7piKhd05yZD
o7aN/y8USLM9Y8IPTnCdG1615QnkvsVL3qMEQR9nqyYi9ord6tYQAvP83qAwxkVl
fsVWWOvG6nGf26vhXDAelLV3TX2eWO4/WicLkjHFgnlUhcv4ei9mt1XUHKVYg0ft
2NgdiVc2IU80GyM3OQnlEKzSXHFfysJP2FcIAtSTeCJKjbpcnMfVD0nsROHfDF0D
gpnJn191r7ACKG+oZhLZHH2tGcWVfvii4HoRn/8qKa+qLiU5d7XjFov4jxN4phtv
70RURn8whk/giv7SBd9TkQaxK+tGNKw4YbgffmcOwrLayT33anuCZi2oXpFJxCyX
j5B8b2yI0CR3RpC4vFmm0dQgS5qpB3RbPYz8t2bCjxgUpYeWyPLILa+Y69VZG7aI
xYAodgAIF9YBZm9o4CMWXZ19KdvNMrJ/d0usoxJM/QYKIaDR9rqrOUPWDQjX0YGc
QM+z66OO1rU+7ggvyc9+pkIZv4GKbgacHXnIvwC0KynRt7t+qq9y483eGnukSV5/
z6Prnj5Uk4dj9b+RZBU6+CTnqiZ0pG5LXGmjEHed47HkRpt43TFeR64MhoE45Gxp
DZI8+iS/ZnfAowjt/tM9NX3aocPCgo5Gg8ju94n1u0pHeBihsH/bjD+MxUOjPktc
0Bhu7dlVbmajPyQjaF7rDgJnFNWPHdPmxL3eJfZPrhmR+5eGmyCub0f5roSOhuG/
xQdA8Gq/J7RNqm6OQ3hxj/Rl8u3a2L2yJUrWXAFVDcW7XlKSfNW3mumFU7CY2PuM
dHLLbgxKljN1RZDqXtdqX+R7D1ZdXMZvWwIhcevXLo2NcWkykDfc2PFOEwgsy9vj
zuEMAfU8SZ3R+uAZ8B4b3CpQC1MPpdAWXmeQE+xGM2fPETlSu78rKkpyDQa/TnXC
T8LFW2tk6WA3A17n9ZuGZgJlR2Y9/I4MEsOAryT+wPs+S6AsoAnGEEm4GRkh3Uve
aX7R/fKUnqKg91+GYk9bkU7dv/SVNJYcQ56l7xES3Wd88muHxY+BXUimLGIUrVgV
XRfKQlZMADgO46dlBgx/Hl6lxtU2RuMmUf+lGJFPtxhuKIYpKRKzmd16SLCGLdnh
Fb4lwc0/XdguX40agHjDeinetLh51al/DU045HUfDYBlespwYrc61/Kj8lkh/PRU
jTxXeHn3FZplYemvJ3cqrxIcNIonO8WS560xqxhz0G5eWQB4WrjzcABkmRy2zkeq
a/yVslDKm9rRJ7n/1LU8gVMxw2OFPBLGRXHuDGW/ovjoON9kPf+f/liJBDrlzhJ5
40h0fGIzM/j10Ra5RKkwtSghUT3J/nqfTSbfQ2JVsDpOpeTBVKK07G3milAWE+2o
q+1aPU5lswxsimfCWeQDxjQGBBFWqdNxhDCMW3aVc/Qs1TtqQdzJDLUaN2sRCW1O
0lyD+vHNPvPXPuMJoghCC2JGbTL+6l306TN80YiOdTYfNtF9vAyB2n4MgVvNze/M
NO0YlbTByUqJB7gbWt5usXIs4Taep/QL2z9Zup/yiPxYg9hIbgQyn/Cb6+b2xOWV
3qp3pYs91b6AOHnCoC+Ul3xB9BRMje6TJ4/YCzYURY40YVqmU+yJ0SCisZqBV3Wt
nfcNaU2n0RFe0Eg2L5SY6h2cU7HIvMHzWRI7jLeQCltp4TYx5GEp+VRrnUMunsbd
nzIQ4JQhy6X/tGx1wEu7TyJEntpb+azd5zAmgWzONAvFc3sBsZij0Du8UBa3VTF8
218WMRT1XoYqt8EWLisiSTjNd82BmIt1Z+aVKAIhX88leh1eOGIRmL8gHh72xwIo
Gpu2oO6/hCQeWTaKDRkqM8mkIAPA0INLV7xg4ylJ7MHY0btnfELWfIOAC+do8Lt8
SZKb04iE8IrqYPHJIIxYz6F+ZopImX8WWE3/w4KqRLaB5E3/uuVXYm7zymYW6xpx
sL0K4mPFi6RpdeBYHOCn7nFx6yWGyjTw54BY/eYkr7pjwc/ORUdy3GGy6o9AzTXq
ta9M97MKsLjJn/dSaZoKKIFy8otn1gDK64r9lLckq8KWxRsqo5S8oaz2JbzF6kVo
7Cri2TzSDyKBH69P+j9LOfiDGFvX3X1xPtNfln28Cj6/uu9KOiqNw1V5CKPri+AW
KgQMNP8DGOnYNqIBgXAKUCUQTb2FwdKmGxW/296ZuPh2iKyxYA5Ob/QW2VW2ubLb
XBwH3gPV0NG7jvvKhixivktm6XrfH4kmIcv3HwjBbuwv//XfoqkqdPccZE8xiyRm
03xS83N1H/UKmCslHEfHmtFmPi9QEOLiHWV07gPWbTGi6xYilEyaEt8DFE9GZSO1
j85uHdXYZ6ECrJd7l8TF4ELv8/q1epNcKuvJUH05ayJLjLAAhWvaSrp1AigbY6Dq
STx5RhQU7iwovD7ND64LV0l5/p8FTzBpDEHgm+8YG2R/dVqVdMGHEbr6pdNm3jfd
/3E8Zp6D9+gKztSXhNHPHcfVA2wceGIvJ7IAMXwFGUwWg5hBP+J64nZcul9SXFDl
RlQxOzMinJ8b8kSlY8gNESgVxEXRQBvcMd1VyACAdoiYt57T8mf8RQihS6qwWuxF
zn54OGTjDEWtK+FHRPoZfMbM6N4y0orh/qohDKway7eIa+ejilFDEb3XSo9BCEum
5TCq1M36G+onZ9QEvMFfRUc611W6FtMpgJgas8Zn/FyzNGpxwMaQ1h6vKvNW2Mf8
5cWg5t9N4a7xaDPtg0b18gv3GA1ENwD3HiOpT/lmplJ4QiHZWVqI65qsmLdcDFeC
gIvYLsH490+3SN4GE2YbaRTtndikGs7nCGtkfpwE930J3E35PdBKsIRHpZvEAxAq
BiFBNcWVV98s3lPNLMFTYKdvg84BwPorlWw7GavrA95yW79/prIwxNqtCbsu4RyI
JOIiEZBlDO7dzPCeBL0l/0bf8l777fFUJEFpLBd4hu19o+Sn56ZKLnb2YK9+F6D0
IMm85aVwOICOW5Ja258/OWYWwCwMXIJaoy5mQ/ITUsz60p3n2tteTUi1dudg8kAd
UCBJPUnrWod9YQqAlj0ZxPF+ZKPzVs85IrjAA49NGKMQJ0cn93T5ehaHiCVHhb1n
4I84ou/P0HcreEhhHz1oOM+9QR7m/K8FZ54HiYzpjLg8zHCUT4qkgo1sSLtXbxMi
0lcM/Lp10SiD+9UJzKgaen8/y3SXoNmgocPciS5ljMdjq0x+oVwogO3vp1ELhzqx
ja3bmucY1Ow4OheGRj9+4ImcBUVse2tfG4dnjPqw+Sw+iOgCUF89LZRNCwfmXKNy
L2fkoDnwxKdAwNeGxQY4vHNuVBo7sPxignzucdlbjppR9mkNh7/vHKCoqR5LcB+0
AgxHqe5EdGZbavtZQJXRNzAZag0QC+whtfl5vfkdh23/9kJ7ASejCpEVcV4vxTBD
nn6CCKv9BybZavwIEZfEhlPmI+yKMcRhBysq+ebgb64a47tNEGJznbNpMsoY55eI
j0HLmdGthMd+7FkyERD12eoj008lUaNk84cGa/5FTFZOGCJYMFKrW87xTRbvbWeg
1GFapXGsktndFoBRNKubaotL91xrlgrgxiOvhbnxWzg346vm/n86/puibfYzPwGj
CgplaQ2o3vmubbnKv5qxfiUda2yNY0NGruSHAOUVP94XAUut3inHeDbQFENPFZYR
OrB9/LoIqWeLA22Uy9rGsHBC3rOY+eE7YSARfhOC+GAhLYGpLk82C8NdfrWnHAZd
MzPqNWK8/gm9ozdl8iNzk21y5/y9JpOLLqDyUP+FXmgTWT1rwN36VWZ7vKQTHnAk
/7zLzGY9IEI5hu7AHlwyBSxf3zQ2O7mSSo+UM7um1RzoicokWIBoX0tEoum8jAvQ
AB7w/W3BLHg7zStLeJ5Xn9ABuwkfKg0Uik4vFb+Fb+Xc4LGgbCMLJwplWopNzpDB
0PcrvqkrYdjFaDDjukmDIN7aXYBiCklhO6EYL+gxkQ5bqknUZPr3Yb+S7o7M1+Qf
9vSWJQ9Li85xp0O0TwgGD4V/JDBvU4ER/E+TaxjPL3Fu5hyGt6NoFH6atbCbTIEX
lHT43FMWxQCaDuq4UDzQ0z6OMU6ckw5kLbcZlX8MTkv2HJ5v2AV6UlXRY+r7VAhF
P7OEW43Y34TcdyOLJ1dR7YqqhbXnLBfAAb6/cGeVxBW5NWQQcmdKIeFntassa0xD
6vu9Rn8AO2jUBtu9HGkK/M5aQ4RkY1CGtLZiAcpo0BoLKFi6g1looucldCXlE8pO
Q4vjXfbQILULx8J3qWGXnDbI4tkMBQp1N4g/9PfNJj1rtkPXQFk0mfNsoUGQlmPz
JcEc/IOKg2udfaMdRPrkP/im2N0be5GsGv9uXl1PcnITFrfxAdFCUQ4+cHH8qbn0
flPaD/DjpPep+uv97oMUcpNf5g5A5MQU8YDoPyisrMgXVpNvdk0C9DY17MLD52Xr
XYZ0dcEdddebBTQ+XTTxsnsKHwEUhsM6Xcw25okKmPni6s6gsdkuavT/9AbEwVO/
sQfy9oJ9p8ZjmLDShMe1tKwNz1JbEcoo8exEXqwCfLnzK/1pFDA14fDbyfjkFM+b
6kiFBVKN0moW7AArjVRk9D8EP/Hg79cuRTWF5WB/85q27HG3VH8BbXNU2MX4+tUv
PPbMMf1Z2HBd6inj0gSMsRn5ts7ihFuS08LF5dZdFW6gtrDwXk6vW972tbadI/aQ
8zJ9FocDEf022ChE79u2OvV8Oz9WjGRiRRRB51b1PfHQgJf+LCvOWyGymuJ8qIio
Tk6zuL/kUh/thGo4YbCRaqOOFOVgFjzvQnt9WUdXvNydK67GGKHGcdfi4RUylkqm
L+yCeAY+Psl8l/zenbior7fXyoU8QKhC/CrUxR1XWPyC5P03AMfvqn+25+mnsJHW
E1N9xlEPFngEYDkoImyF2nR+rxs4QfQBueUvsx2yyrqeMf56REmz/gFqzPIgM4PY
BrQIXzxyYVxF9T47AxHj1f8Wshf7Z2LjZOauc3w9RMby85CyHv6WOQsMUHBFvvVx
WpIG2sqa54NIwo6rzyJ7Lgky+7YD3o+hydPi1MAIfKF2QIlrk4+UYkbSBX/Hb/KZ
vxyWJxYupoUD8jM7Vxi7OMFJbNizIIhRAaxlmQuB/gJXdAyC9CscC0GZx8xpdTwX
PW0BjcmUANlDgsq+kaLDK48uRRZQ93y0sJcUL+okqEtiysiFNbu2ESdHaBJSFltg
0OumyJeMJlChfJgIya7cE5uRP0MKNxWf060jUPIVpCj4eAZUklYTD0GjJ2oVuZJo
FAXrTOpeSKoF+Dz2ddYpi3U2rVN53cCDOqKLd+jdvVa2tkyY1VwwhjZCw1mMuvSY
p/p7vB7KnM09YsiRdukAsU0PrYlouvVtSACzRJgCgORNYShctW6zSGpNo6BMF4Lo
jplY3VqJEqfhNFkIuPkkEt69QCZkly/lktWxuQMVMjJHlmd487FTNrdszq40QSh6
DzpXwEuYLt7Y8rNaBZIB8ZVD0Lft+FkJnBetxotPb6+yNgqiW83BMLMn5b7Lb9UF
diIKh9owXaLfFhuQuMkUkpyXPKq2dy0YCFzLrRoNfMCZ81HfHnTm262YAdSPeO8V
OfNSSFP5il1MFJFOxfJhhgIaX1lo+ZpVQR9cPyZwXJwHDe5itet8Pndp++sChpwT
ZgnufjfHvojFoTzW74MIwDSlNSfYqvTSnzw6gQHxN1dPPzyXZSOx+MhdcNyFjLAd
0+Y3KJyM/zHY0mUAXWJvqyc+TkVya8FLUYIGSsQvSOIMC7XWXYYdTGuGopS9tzoT
XuAVcJfyTp/IFZHO3UXfUb8BUTdaUsv0ocif+K83LBz0Gm/5Qlz51NaEJG/w5kS7
ia3b6JvGEWm+OuisjfUacxUMPMg3PzlOkzzU6N43SxSXzhCQGGcuGPnUZ+e4PQUe
qfAfZWZps7yBbY2EwVqC1k7Icon8MNrVrF2RNLsX3hhhiHuXJxgvcKIX0IcnIJ6e
nd0dQQShSPK5DPAGoFOrTYl7NQFhRWoLcdcbaz4OXNi34xgMAu6D4dN6/sZ/w6TZ
gMtDHhG4UitS1bqEC5x1XPzYNrCoEYoM7TjFzvNgoTPjqmlKm+Uz8ba5q99M+u0d
SXCLNB3ojgqbs8lP2Y1iBuRzATvr5TOOmgDseP6Ls0wF8b/HWKifFO1a+BqABYJ9
ZJuiRnPtv4qNsM7n9NkIMjwUOdDVuLjx/4Ro4miyispjoOYB9KUk09mgUsyDOgaS
xrTyisKq3ya33WqIRdEj0WbaJyOIEd5n+ZOqH3OyJE8COcMeoP4wTzidQJVDrB+z
B+KdTfwqo76oQrWLOSS1vHybyD5NQL5FjhETSYttiDPbTOzEmUMYUtc9e7XLurmP
5dYt4+Mht4zBkJ42Ai23O+a0yifA8QAOhsEzcZs83tlgZ1xW1bM6KnA77dkudLCQ
6iTZRmUcytpeiOq/hulOi1rYN5HDAIj1RaL9ghOhUATg2qfFAkqF8xGqQmp5qNl1
y3NRrImgAS0joFHEnqPZR2XOqPmszU14KVlYbQ6oi12bD4TYfEsa8rJCpPTzcbiC
1nPiddx3oX0xZT0Ptdr+iYkL9kdmUCYMi6FDJvfNjkBO7pRXqPDYvkNB3b0Ah1nw
NRC/MVgoga8cRJh8vqX7YrWMDvcLSRi1p0ZBupEW7WmrIKm1MtyeUHTlmA3EReY5
vMMw3ez13BqJ7CNPqg8+Jyh0ezF2yYrI6Spgn4CMmbTjOab3AZj87qHSyKUVZGU6
EFwtKpU+7WIliT3Y12w+Zq2OEfjZjyuBNaXp5ykczZVXkWVmzx/2KMzor6Dpx9AN
8jqThexj/RoHhfytzNiCRFavQu+2Vdwm5cD33VVlybD1dKuKwjPif9JEnVzpK2PW
+fwhdC5Jinh4htY3rou2yd9D61r+emTsJZHh0J/j2JwE2zyfvN3qPL+g1cbDxKnP
NsEKvYvBP1P1mZixtBMztzOh7YtnEDwOdAQhMBHzzLwuoFp2yUaTHIs+2uGKdmC6
8qISkcmG+CIcX1yMAVvddWS8rvlkeHcOMSbr8YW3PFtFJfRIFkR1jXVYOHtdX0NB
xvQPEqn8qVc0ubb+99cAYfa8fAddAhVkierYfXOuBT1Jz8ZcW2kheXMPPxJK5jeZ
xYB9Vr0KJNGgluXY8DGMY+FF+U9i+Ps7CGEos7gXOimUu6sJ1iJFnCGYCa54kwHI
mhOT7J4+Nzi1jQbCyV2rkRhtncaPwXxNfMJydLqWQJXS+Sz+Xf5LN/Imc7wK3cb8
e8X014juaDpuOWVqJUtBUn5ooNjpWtZiOpl3eKpBfhkUrl0Zf2L62RI66EhxGFXo
gTY+jBidGQP27OWFvTlZP20wkfwQ0DsUk82kk3fgJVnedLxyNl+lLifnGWy5mrGw
frEFfQBvXHJpkOgrbslWl57t91JrmNhHQbkD83J892ER/FoX7zM6aJMGujb+1jRA
JasfqwuTBT18e4yaQO8OAn9Y3xz6+N9Nr2Ouo8Xn60t53yTCjRr2Iu0KkD6Dkp5S
LlrMhPJCo0pUHxLZi6pKfxNqKRopQh00EYV/oKA5lLLnAiqQH/7rBlPg/I2RJGZ7
DZX4VLGqCRg4t9gGKYkRxC15xaiSIrCGd0tnPw3dGFfghMEIGBnqdALxEJBsJPAd
09N60MLNPpo13LDnwNRzAbnoA+MBERBDpuSwa3kckS3w6njOl0FzphE786IkImbd
aRZAk8DTtqbLOQUaORFG+b+YvNAYGoNvVNJ2GHrNdq8U10WnJ6opSy46WWtNcVkU
ectNpWaUUxSp8bNtmrEIMZuSFAOnzoo0ARaWqtsRAmvb6fu0hkQSAu0Ftz4Mu8Fl
319J4d7EVQlpaB/1crkgEuU5OlfummAdWTCjRRG+4n3UfU6EarB2mGUKolmDqqef
Vch9Ypq/9NtVZ6du8o2K914OyJx+KggirXz39xo8CMyZnn/Q1H2rY3Bz6QBP9vQP
gbpHlWjeAJCtyIxOL0HCWjfqcWgyvBNzalfsQ2EoDwRTVxYByYleqsVuFVzA4RCq
7NdmHqPG5BBeXruSDJRp94BAP/VWgtBXyOteCMLTdbXnpmiyNhvMFmMAEoG8HuzO
InRp5Eix5rcu2E7ffZ5KnVatUJGXqrTQPUFCOW4v78uLToq8JTGl2G4+wWjSEEp4
5+ocPp0azZD+b+rmjVDiA7ujCCkRQeOkYsBI/MQ/FyF/GG0Qec1yQN5CFFLAJL3l
sBW31pOYXMsZvBEC6Lracgra6xhN2pKJI6BxDsxaXqTDv3QNpxHVw1/ERnWqD9Sg
IYpliOCUP4ygpYvRpo0S7Bhth3RumQosMDzBIK+46R+Ir/+jfjyK+k/Lm0SgyfHC
2a/mYiQMuXuodJqAgbAKrcclbXv8RHG7MTDKqUyF11netbLwGJKkm3SKB35Lb7rr
v19qjmXVEApLScULYxRSi1H9L6spCaYUSHB61/Tu89Uq9lhx1uO1ZRbiNbUwBX2p
vnwAihMYdxiLYpRhSLr/RunHR+kCw1jXVJsA8te6KcZH6EthJqPStTt3mdWOVX+5
8aBAOlI5SPKPlYwj/wEci5DPnRT1sioznJ5nCY7wwOtP/OP8xv3uDiO6srfWCT39
B+5mSAFN/9WvkC1H9MfkN6LoSu1EeAjCztqUbLRXjARgNUjilAoLvPszGt9Hkf4P
qCaQzQT73Yl9br24qsIhMby/6mDkRSJDHfeQ1qovd5GthM67h58N8YevG7EX4GMv
8WHul4ugO7gr6G6UhaK0ihdoEsBd6szJVEDD5uab060Xl3svNr060DFwfzGOghPF
K1om6JWF9WOMn4PaQwm7JgSCGnYDzZA6OcbPSNI7miJT3mFxPCt4FtXiSbbqmPZb
Ee/FEeXf21HgjY+ueTMDkJ/KuUZWy2sEhvu6uRbdZZWNx9EmcWxwFIUBQAkbC5Hq
ZusBJOWg92C9c+yH345jpe8gBkRxyJSNpWRa2ESKvLgDqk4La77cYpGew4qGKl+q
UVRknq8ji1ddhH94z4lztkKYgtcXd9j5y150uNAexmLqJsFcrpK7aPQlA04KbQUE
QnqUNxhPS1/5ij3uk2mYitQm2yQ6BufzXzO/fX8OyOM1UziS9q7zagJ5+AKSMnIN
IT+p6zJW0JV/J/ln6D3KIFtkjU+22fXbcMaqFJk36dAPsdVmpo0kXMjB7YVdzuyV
2us/wJSVVe2AI+SfUeYLg4DxPCzdqKNnyIlVp837gM5icLf3Jt95N2/o6hCsTUgE
exJBDSdbjBYVRWeJ9Oj+Jcb9RXBm258GsehEygzwMFTv40CtmCz2Tq6F83++87pD
yo/xISHuqb3Zd2jd0en0JgtS6gTUpvZKpyvf1dpz0RNFC291KtdLWVUVu95TEWc6
UAg0r+XikHWTVfoxPYyY26PheaGLchiDQpoEJG1r44z7JxpcowTcDQEodeBDQ43h
XJns4CD95tve9bu8Mw6P+WV2JNBbNGoPgTvxq+xqAj7mjVnPzPyKrAwOL+YX6qOe
viNv/0G422NdezwVnI+O7YXdp40ADWFZInEFAEaMMfPG215EyJzlFT7ue0ENbn/3
/eYB5f1bxrMyPtmEWbH8nS2EZUJI4pnsiEIrs10CqtvboVzlgvCfBcMeB7EnxLlP
oLQlbqEyy4uGnIXwn2gkUs7fNtTfMwICM31qnckExIzPLtMYcQrULu4evXyR0jlH
xnEBGwKpct0+ZyIwZ3G839xD7k6uOOgeajfajyDbKifAMhQuBgBjJizEcSBHn3Y2
+S75yCbIQ1PFBFdjmQp290fCSvuCPYD5UDaJc5UedPpIHyhFWYlMcmWg/PB2EHKu
7yiGmtTnno2ga2kX/Rj0jypkFaFwoLD6ak7Ga6npRNEydG8w5yhJmKs7vvo3c+fe
9cyHP7Rwk03iBAjiBpvOyyuM2mjCRfUlStXmYorvTdw3yKJejuMM2z8m1wqgDSHk
hZ2fAusKfgoap7S833azLhoUB0cY3QoegC3+ereTkcF2DdntRUcGcyo5vVchvb+I
WjGKYr5Fxlr6R96MxD5CGp5DF3Y03+dkARz2X0bsb34U2azmQyhdb4V+YiW7T6N4
rfwbqxMKkwQHTzWhq0N7tJdebho1rPPNa0ZYGEf4WRXggKJ59yPC3nPBdIhgZySU
PDkeAAHErTRCOr/AQ5svgcL6I42kNgSpSQxbVZsCJMKNs8NvaCNkqBdPmEHk6mZd
3xQLS5ok2aWnofmcx+X8BVzpVLTCwq4N/kXyaG6hN5ksbX2c/09tdv3+cVxcrBHP
4sN0mBWI/1LnJKY33xxqDCTLSQEMG18dAN5OY4XxLHBMLFUaE/mpYYzcNjmaC202
bFkH6bMXg0EUaLwa0o61IEuv+zLXIUj906V1S4QZNzyoYfnwOht2xopf9ni3a58u
orcXradZgtlVFhrhcxCzJxt/PGQ4TTQvAIYMALvRZ1Clqjogq3NRVOACHVdU2X+2
Ub1QDOM58KAjLCx+NtU1BOdlcthpyR5BDZCTagh3e9jAcp/bmkOtf6/tiJug7g1p
fAsy3WeV71Jfbn3yt+GMLyXZ8oUqHy6P/ciIh+AsgZBX2LwuSNFwQL7flEjRebzL
o9Zb5yw2EmiHJ5kWeWwj7MXhQZ8b9A190EU4A9r0K8VRf4Fgg8Nuv16TDV+9CAAV
xDrTNNKeq57mh6WKvJgzc3P9lfRMq5P9S6eQVEoVKIuDXqeKkYk8mcefA1IR7INC
xlcfLMot4AV4eME8K5CcZwaEGvOew1r2LLX9yRBtuokz+1AcaLaOuNWbseBi11PR
xYA/cwlsc5+IYPEuI2iuZ9Evm5bxBuBj9xQhb37xg+Czu8RbcUHvVrt+mNNRVjNH
YSOZiNN3y4iX2B/IQcZ3HL4O0IJTTHfCaLtfVXqm3lpkrCPW1p4J6v5wXlS2E6oR
Z63LVqD+YcJYOtqZShEdJAsW9B4t15/L1llpPrRnSb6TOcFqxQgQM3xuhbUUgc/t
t04O2PbwGbaNx8N6Z6UV6dbezK/GWra9rZ1yfNMIC+SabpR46uw+wq3y8QsDlyTX
LVdnAWg7wp38PYKjXxHoczwRa9z8XdD13R1bh00auEiiQiVBnqUBEjyT3uNxGgcE
uKw3M5u/dKfURV2nP0btRih2exkag6QLrs5heDfL2xaLYQD3wrhW6ZyiQXkX0x4y
TQ/9oIbL1WkzujkdWHAjKFLBOBisY8jLssHIMyom5RwDcqgU1kLLsIJ5EwPrA8lw
kSkt31JxQ6FHFpVJVOwVtGoU/I5lkSH7kVRNGde87gd+jubwkTTaX5g29PsUbId7
HEFnK/WXQiaHVYl3eAzT6vvkrTxY/zwQSCiEW8paTaVczkDio9Wz7K6e1dXXs0y7
YjW8u/dYG86jKCJOANsjdfWYUbTdncwhZyOTzy+omQ+9M7zhY+lfEg/T2SJlXWaT
a0lwOmxz6zuXW0uyTMMydC3VZn+d98FTq5f8S/P/gHUTGVbo6tqG5BG73z9MZA4E
SUfMP2sqERPCqBts9yMBgYpYbZE53keS6Hs1EoxXLJ+XMQU7xjfJqzORB/FVgOL+
gH28mg/VzaVAb8WJR72u3abzytWuzXik/arn4D4zHEoZTVgXzpGQqfwrSsdiMsqV
sCTs7LxRYxzI1Y4/zG/vMjqYNDw/p7aDsywqspZinMY9AsBYMvcEEV+KyztrdkBl
+JjlW/6FMKlc6ZTtkJlWPGf60/AfkT3DpvpNnm/doCsXcI3sbcLJ+2dR4CDWbney
061Nr/dV96QPXkxEjMvKvji4k77Zi/l8siHnEBsGT+Lv5GDvWp3HMc6UokuT7tCi
Hq15BEobWQuz6ZgUJ/3rnf95OEYGis0jVt5hDolWIIPMXZB7khIBRo96II2xV1cv
P76hneG/hEbmiuWEJa1XLE3yJFBikKY/UCnyl/c8MGhsNInKSMTrdlQFVC0/4QgS
01p14v0m8pbbsmc2I0ibe7XxPYEQw19hzpKcO53h6gQcDKxH6m60KbVWZW/URH+5
GumUuaZcggX1sDnvAy3rA2KIyMVZIvJ7dBncjM4sUtzEp+mJY0VerjL32H9yX4Py
SSWLD1LX7NIj5+BoOCpgOAFWZor7jBW1w2K+aQIB5mFb8LXYDlSwuBl4Vkd+8fIr
sy4DaY44xNq/NLUSZKyHsop8J9tJ9xn6uVjJ3MOm+ILL4036Uv75/3+CxQPnWTXA
Y5pFAoOqtDwFZnY0LZnVbEhdLTRJdOJ+IAeKix8fQpZ0ZGWWppEOhlDMFUKEGoQx
2vIUTggpA44rtlukfaSRq0ORGlbtwH0rAt7pvOykMoBy6lWkgv+sF/87pFuas/EF
l3EmAzKZ1iIQTiaZexlzFqUWsma7k6G8tC0L6v7Fyw1ypsz8tIIhkwI73SityaUh
KVN4o2bA4bxe+XlLyfRg6OZTyJVTLDYPVu8yHtCHwl9opIAIX7AwNDb1OehSgTlg
IFvfbuIOT+6AS7qh8OJeozxwGUt5zBO467eOIY6t/J/hvMCIW1GBDWLwEb7yd5p/
+Q9VAOGHEh9kexioExWirUGD22oqGZAZfdEaq+OWqHp8hi3OZ0Lgnbq70t/4FDPy
zDBDCp47ErY8wXyeypxCTqkhtBLH6+8mqOFB012ZAFx/je8lGf+Lmzp2kU+itsfr
tqj3vkbBJHycNjpANa99rZAt/EmQ+VPTOS26m4bHbssHhwvLC7CgLU4KP1aiWk3d
AnwHQqlGDzKu/6vENWmbqtIzZx9qkS2wfpImSAR2LvmrkVv2AlfiXd8AvEPqZWCB
KQO+wvWPdzLjNOcktWQO7GhEi5EHsD+nzyN6dSYT/q+ka5jpO0K+Twu/BolNmPwc
Xc9A0uAn5mw8sHpVMONtVmnufT9bI/9GIXmpiBbBmR4XzOLBqyjK0L5tcM8+lEWt
YW2EYUQvvy4LK8Ts9l9OhT2P6WyEWWP3ruhsfK/8J61a/vHVoiGxYEjo6sGPUt6X
OaXipxQgHNS53ABHl/xxHzoRpm9c/GPRpVfhISiygG6HEK2lo1B5rRRTJxGpXWeJ
IYxZDDlVKsrF9Z/QEo7DP0ku4W+aTX+BoXiO5G5IHJbLBfEImWLq/Kodnp2u8hhx
MpG88qYua5ZKDQzM+im7KLkQOVlgYTK6mO+btZpQD5pC+03uYMY+sUI0xzIdOggJ
bIdXoOQteUeGheY+yTLjrUWaAISP6PjEjkN0LwDYe66MkdkJNORXs3zWbd4AwLTf
4yLQdVS7/w4DpGacLESooJkweU+yGXFVf1EWOXgssEdWxyls2VW76Wgbm73HpvwW
Qk6LrRbWRCjWa2aDzAoANR/+YTYwuahreqVNB9LFW4rIBZ3nyGzaiuFEHi8/ldzw
GR7bZHFOfHi6JGFMoqtL8SsfjUkF7NTPP0Rfc1ysBNHlHRfDW+ilD31ZPWMNlQtg
reavB2th7+Tdr0PxLVUrIiMzo6TgaGfQ/z+UocJuCvOuXFoFGkukEQCyOUeGp2yQ
4u31zEJwpVoLw30Hg44DJaQvH8jdEv/uhNQHtPMW3JCwX/UMTqLBtosGQbNWkZu0
mLzg7PKVSqGvXXoR2wb9lImGJQLP/PcyMOU/tW1o93ajt+1c/EPPsqeOwYTQBVVL
7/cOCeCUrrftW71I3PkpSQScCHrSFsjeLnut6sehGTtTmoyB+myBnJF4EnKsq6yR
Yh/DUdlnffyIrG8tba0S7fxdu/lZMWFedp853XO/Lc6Ubfw3zEr19T7PwydZFo8o
muaserajGdDYgCJrLMlIl5vhicNCVLgZAMXqzhCEMXDcMIhZvS0brxMpnLkyk3pd
rO3ytt3ndSWXaP1L/O1LQFxSe4Opi01EDblpP0VkYBio3oufAfJ7NwdYnW6rxjJI
Y4bkMEp1Bm34QmYVAEBRSnSct+VeHJ7XC3FLqJQ9kM8NlJE8hZTsth8hHw4GE20e
133jEWk1xL8HHMsQB1Mj9tVR/DELyIz/McDahMcv5iF7XyT+U9Ph6FOfjgP7l+iU
Tuzy6JtyR4Eme5x1CWK0XvwTa54H2VJOqqq8jznO52Zpiv2zID9ooGGhOEkLUruG
WxzmKNRQXwkEuzDG5tdZfxKoMBAlgCF7xKjbhLRKqGd6PX4IzBMEhp8j9FUuoaEb
wOMMaSFg8RXltxOdUrqPnETNBXA116OCETZM0Gp+rkoumO7YBwYSCZFEzUeZtkTS
uHhPIDThEQ4g/dd9v0jQMu8jERHpekvQPsRP3nftKnu2ZltjO5zsPUI1BuaLvs3i
uTQ1ILY1QJI/PRINbGQxJCnL0lhP58zOQu7INuCRRo9t/fO3g3CwDwEKgst3QF+5
acD8v8qQ5XNZkBDY2vaPb0oD6L1XopwsAZmqPgAjfzXV1Shg+1PGl0tbQo+6ZcFH
sj/y00HLIiSUuDXBtBSSOBdIDxqKpVoxNNkqLujiQOow88bWNDy/OzrcO78/MeAV
qVee2Q/YbHz4p8oZyQoVZ4bvpax4hQtpbBG4XTEUpA+EOnHXOkv1zWPL8tNRrg+8
QwGlshLIqp3nYjZlhToaosclaH2h2nRBUqFspYdticehna7Xcvh1fjk82LnX9e4d
CwsZwr6FghAFlxXc2ErEMhxtHomSsiUraZya8nnnvwsilCs3FZJNFyQS/I0eXyuG
Gz3sikkN9rJTOlxveDasMxLy3bi+sIp3zK0mrie7KG7+tokUW27lBNxSBlBznFkD
z+sxOjjJ3ULByeVUqDKhwwQtfdLmZChKOQkTeJ5HnczU+44Qh1l/sMhkmL0uuIq+
GP5FtyCrzErs90QPCwQAqpvhdzFsS7EE/mW8UwKuSf7RJvvIs0Nlu/oNRcygzjdf
5EJ7LoSHWniuERscNx3BAuykcqA1Sln3uEKdwFy/tJt9Ic5o8abm7asLw9sA0N9s
rcJq67psp1eitEw5i1gXft4Ax18LkvejKABHCN+ovX/007m5s68nI7UzU66KOILK
Xywc1IVOc2xEDhfVNHmpmvF7PvaA5R3jL7XcJqn0k4Am8ITU0G/jYVfxpoQwcFuH
L56A8BSn4HtWucUjIbWFLQgvPzkBWsmEyPsObukHwbTRhG8tpuBfj9YET/QSao40
sCamPUeSZQ03wfUxbPeJvbrgSqtrz6jgg6Epj1EIQk7oJM9P6NSOfBiImPOA371f
ZYSnzkEIgMu5S5Ug6JaVJVVZIi8EHXrhjo5EJchemCYKtHJeY1UVUALysjkIaciD
Jv6uvSRUzKzvJqutZX34W9+D7HR3QmCCGaa/QaqdlFws5OVj61mTjJnMYO1fvpxr
jdl+6sfR8a6zBaHBBQwJRVBNxIppMzNkMiRZtZVmG6Dj4G1erfmaqTrttyEw+qJ3
zh52yMP76/pRlmjvYNZtL48kbzyRCeUBiVwgw8mphANGmHe/wnAywbwZkwqgAOKR
tBqhvozZQIkG5Gzfw2oOBu/XKl2K/5qCDO9hqTrXn5onNJXp4wbuZaSjkeBB4thW
7T9F5UnkBODb8TX29RcoSOBUQlClUsp375GqFZRQ6PsOwnEn4u4/e2ckr5O2tvXV
cIADn5fiiPJj757YHRCvgPiEvvxV9H0L3Uxu7CnWY74WQeuv/XCSdSHZa5PG0obc
YeW0PpN8SfSiclYOYk0NeGCXAXyhoHkjc6JRkMWE3IjLPQc6HDmr+AJGuu4ulrAu
amDQzNb9AYbOnEa3JFK+0xPDitbv7QGhtsgJZiqcbxu2xe/+x9PBssqS59Qpct7d
RBP+r1mxCPB1Ha/hiMWw5HSL6iEcaecmZokguNn0gUh7UMhSD0/XP8nLy/RT3/Zf
VccmqBhl/i26+T6NN/ba0W+qtugfg0xZjGh1o+4Y6yXak8H41VYlkJ5aBKE/pEgB
m0fAPRjTqqPazus59b9PZWyDkBU1VYN6d7Y6TobZaIupoIWWX8kx098bTFVqLthj
+ScY5uZYdRe7J71xWo3MJ1OBX0FDiiRDhuxVXXRnAfgpl3H/yR1u5I6fmwqFEmAK
kqUVSSC/ywb6tqteDzYE0SjH/8K2k79Mw90o+g1RkOio5Mxjv337CGDJNOIffUSa
InFx2WX6OeabfLp64/uLP3X4+3BccZugkWXZnemA1J+TkyHrt1TRNjepCFZ7nRwv
cWr/VrLOTAm4F9QICZswkSjxCzV94o/QWF0W8fgBjxcYVNZHC0KD+1tjpg1PJvSz
e8Dsq5iNNpELbxlQ2QjkRbLrpys6WQKf4mr3CARsuZZIKrwO1CyMEAs/hsAMzKcU
M+ZMdFlW++sFuAjV2nuLEkZL/JDKX+91fkQ82zMnaCdaEIeia7ccXBlJxdyXYugO
N7NcKnbMB/2vuaIEbOWC2SMnl8mWtNsN75klQalicqo8VAccWUr8CoqMyF9STeBz
vpNiLYinxPqfEcJvDq9ftorHLl63I59mheT4kC/0eL9XKAc9ue6CrBv6nOcZ9sym
ekjUGkRTPPFnS3MO2VmDR9PfWzqBxbMQ2S7Xpz8o1sEZdoRku5vUXFevNOeWS7Zj
neooew+sNJ9er8/qBS1Vg0xjxQa9iYdxKIi5PgtMR20fA/6AenJf1FMWKD6Mj4a8
Mb3LR2Tf2gqS5mODs1RC/JivqlxPnnGi8qx3MRZl59UZ543yuqoCFDxdM9/yfeA0
8QShJ4i0Sz1qzgVGIRzW2HZ/lKMT5sQYPjfwlMg5h21DFePec5zSJN9R7nOY/dL0
CwTqvF391fUhnsE+dpsB1LEwqW221JHA7bBeRw31J2OZmm4RaqXBS2FkHwPVE1t3
2IK8Rb/7rVOsaOghVsWUhMLYWa3Se/OE19ie5t0g422XeTtjX/NoEm6Iqu7aYBPM
85mzRrgzdLRnz2IUzGb8a3w0hmlnVf0DLHlZOMX4ZbOQpe3YKltp4JODtZOx5OtF
o0tBaLU+jOqIFpP9eb2+ZSsIyznOSucFTRO+umL/5nYokv1Aj7yuQ8bLbfJCVjZq
QO2ZE8jgPCNsv4gi3PUz+68Cjk/Ibs05VKXZNUSWZcYg8KtZZNrfTuVqyX9qRq4W
t0CllTyUSTnk83pr85xKinHE/JCM4UAiI8uUSq6XGWz///y2mBJQTWkW1lr9ZNpN
9KcE5Z2QFPWb7Zciv9REWgMQVKwoGX/O3ahsMsbUFr/v/m6BB/GTfNy44tv0IBgI
7hU14XROz6HrgjLXIV+YSCzwiCfFx4r4PJYjHcHm0buxB1tMCHiYZ8LLkdPn7CKG
LHkIhQq71b8K77AI8TAJjC+VSfBO1F+uuvKwq4K44MvuT2WMg9x5O46ykATw9DUi
aUqGqjHsngFJE1UfSCCSKJIdc+rHge/TqToAeR3pp4PgZNhTuTOA42jedBMJZsVr
FS6oJQ5K2TO4LG55/JAeY28QTciuNQkFPY2Jr9B675ROij06gnwOVL1DzqEQx/OE
zPJ6lhzcxDSk+3BNgT19xNGXkTL0Tu0ALYjTgxA62RIH876mHLMgi/M2gw99Ws1q
LQ/uA3VxU3CA/38FpkCISnoMMm4Z6QdCDntsqyqFGLa/qj/wEJtjTY26fBSleE4D
685qqmrBmN0fkoaqeWNxFKYBcKsQu784mM8iVD/f4ejkiZ+UJ/FvPRl1tHmLCicI
1pdF9zQ3mwUw4p9X3A5LSTKWG9RSvVyyddm+2a6kq8LCI7Az9kWB/oiiWoQfT5IV
/coB3SNcrAdVBFuM3ujifQJ9o2gTus2i6S9HamQmtFmnxJNRu/xRtWgCE4EL4PqG
F5YLTYN6nsmuFruk2vgpSpA4fPLktfISdS4W7svVAbQ8qiBH1qPP7DVhcoF/W65M
gh4ZTrXgg/SYONKj6vM+KC/2CQVtgveZievQiypqCoZ1mVYKNbnHPyDQM+Bz1PSo
4/xc0vEk8dJ1jm+ZFuuaOrQm1PgTVt+B16aCVuddUrNLicB/hKRrfGVrYqIE+UYM
KizHP/jZ5VxYi/Nx7BuehkknDxopwSuzvBJ+Tb5OBuPOBRpz/uSxqVt97/tnjaao
Gbv5j3md35hlPPPBu43T7UfztHGNZVhn0pBj8APcZhWFONLDdoZzi5UqYtd9LRSc
PT/QNXYuVZW7Rlxvge1XQcWytHXekcClRO+E1yTrFIgzPFJsGYfD9x/0dQcwix5F
JOPq2o+OAsPM54zwqxOOKFk2os/bIF56kXVxYO2OJUl8u+iEj5p5Wl31Au9tH4fH
Pg4T7ISAvljewqYnHuf42vSpo18aHBF4AUAqtrFlo0hNpZq0lwMsqhg81fXMPm/E
OtAavY9NLNXtIftRtVkDi9FF73y62TzFfitAVE5zI3lOpJbLh0ABPnjXTGgZmAsH
EH4GVWk68f3HWG6r+LlrIBIB3AeWZxgMjeH1yaNBVJ/RXsJZBPeTWubMZ6MaS+tm
p4vlzN/Pc9kt4AtD6ZKXiYjRT5b7ar4tlz3HfsfH4IrRJsOKK4Nhmsy0QcsqcM6H
EACHAOUftN6KTY2XylEgi4ITb52lTpnr4YpSz1ZDL9RYn0o1azSq1ckTa8QFmvKl
DWUT98zOjrlto/Uppg0M2PLaUevojVYPioHMnnHaXMALFjQNGwpITHj1yfsHOnt0
8fJYb4EErzd0mYgADatxF2flDupUoQYdpXBJGU2yJNVIb9ee1YVd0QiuDsPZu8wI
Sn3jHCy/lbWo5MYTbNnPCIUdUPSckC+vC3P1Yygr9z3Q6uTog7jTJN8xYyDvAOHJ
/FubNoLGHROHHJP5OIcW/VpD5aXmMqwgytEyG4YoiVI9/WIqliEhJqT4oFvZOD5s
0xzILRidv/q/TYlCwEuoBspEi1WSVqFRil8jV6Ugo46l4ZJF4DadehtX9zHP5pzo
r0y+dyMN34BG2yTviIr8o3DrbtBCjCS7utPqrps0o5XS4kb8ejd7Yn6EMtJqyEOo
7LjhCul3oFYWlV92/znLybth5660A5+s8zeZp7kjIzJ2xVj3CM0TKp4UvFO/m8g/
EQ/ugF8mxrbM0HTcj+EeM2rXZIv1h47yMcwprA9x61MeVLuQN5WOxAh9SNacRmoN
uZNxV0ubvgwjiMsYjovLquB8urZCumgG7PX/+rf+r8iApsJQBob4nksN1zlF3Cu+
hZgbnRrfhNkk1rwe2/P9CseMBVuCR91fOEV7LWtHUoMKX5bg0t6T/telFFopKn24
nWYR7g8as6sgVos60zw17aIiXA0dfVNnWeJ5VxxmD/KG5ySQOMDEAH8i5UTm4h+z
qyBQ+FoszEanRk+gLD3rPzdhWKI6a8IgigzcTYbGxmdLi4O3imK85wQjwr8THhPK
iHAvoiYWH2pNVZfdl7V7WWS2gqtVz1d9Nafj4FRkrt3v0vSu9HtVAehfIBrHi+cs
PXi5lPJ4H0pkuISaeDGMdcRW9D0v5P8NFA1CVwEXZ5/nOetXTDZJH5i+rjmxkMCA
WX7fjAq0U57NilWMT5lvcWODaK4du6ZxUSQbAECkyapsxS5uCViIKnsXSZtxHAQo
h1zdGyUZtG2+x+oeUG4Zf4a0zZWTL3u1JXIN2NB6KN+YB+MSKUGxyhy5lioeVvNi
1EPNJqODKKIx4M4/6z47zwDgFDUpjr2pEdpRMC9ZgcIU86l+Wt7OBlAxciBAHbYD
IRQ3MboWDG29+RCh1HBGjq7bQZHojUBWXPCfsdDyq6752RKe02czCezEqEn8N1rh
YYJO+RTV9qw8uwPxBMm9Y4b5D3aOj644dKroLiyIglmDov2bhCpHT7Xtw0ckQ1cW
YaGw7cYlRt+BNAW8MYX3VQ39k1fE59M4/cSXnQjTeciYaxkpkU4JADP4AFmTleio
7wPVsJg3BRK3Ncqir442t/J4VyK8v/wCe65F02oSs0A5zWZ3hJoI1omWJiUdra/9
ExXXcH6CdFqVeJrSO5JZTo0WFb0H1f+mWhsLuuKyVcnDX+qZ6XgekSaZ4S9bwyBa
I03BIKGjv5ehv/D0sDqXO/Y/QXmQMblqo+J3sZZbCRptj/IURYVOijHL/8ttrZqN
d8wv+4mkVidjTdSRV5lddBBN4fEmA1A23FtBadJhOUTBSqte4k6tV63zhqxKY6i6
5s0PR0r7mvRc0gcNJnTCgNScQh9GBnnthCuC7/NKAatAe5iX1al/aTbAMsEcrQRG
bYI697f+oPtFP1a9u/i3P9zXpQGhAhLZnuGmlYGZPMOKpuua++kk+JjUjorO1+qE
hpCp+rFApik/5uaBbOB5rtxYXbfLKtmkTIAtPsZS8VNlvQHsqQDsRppN27Df2U4l
QoU3Sn4X2rrs5IW2ripquZVQlOyxB7kKfYyllwN2EWEgDO0Raz+XPiWZ6FABdUOG
FwjeNRpWoKAslykLcPEzvz2vi4f3NgvDNeVVpzzxUV65aYsh9ARuQ8e40SXCIZA5
YVLr5GCecszKqq656i4xB1SeouiO77gUg8uYuyR9EPqzwpwxIpxUBT5gep57oQL9
qL70bTJ6Y7dq1Tplra0n6iDRt8O0TCdkhLNQE3kMucvOTeJazZR8sbQ50EBbb6dz
4w3U185jhvdsI9v2shiOGxWpTREInHvGl6batPoon5SXQxNHMWJhkpfl/r34V3xL
rRaVCWg6t9++N4NXzHgNP2gJxOzLtRU+NLTMtvBJlR60uzUXJTEozVpD/j2uP5fJ
/6OgCwpu9jRGxP5uGTsbDYENvc2mNF3WZR+FpD0evGmK2ItM9HSsSISZHaXOfVp4
yLaFa0dYY4NKt4m2qTeQ7/ScMGwxljFV+CX1cgYEaQdnkcqGub2yCC0+hPlOG9oA
Prlh7qebcFC2rk3l3JRxS1F+tMb3xR8gBqnbN03558NBBSL4Yp0b7jBykCPjOpkT
ww/iP106ZL+vvv5HIl+y/6I7mw6+UvbgRwlu2D7I3O1RNpetLsIg1YVgqHrb08Of
AlFFVOxZJXK9HjsIDfHvvFm4Oqz4J2NOJoF/JMuTFv1Wm1uBaMDunxbJOWmL3cK1
NOxQ9moHWGyhNQUcv3KXXKXoxp+7cZoXkyDpWBR0zDu5zEK77BmzdE/sJfLFghDX
pm9fesMeZkjFvVZe6XCxzBIjIxeg8m9jHwD7S65nfWp1sxM9d3Dm5bmxHsSReoCD
LgRS7Rx2K0pleYcKw3pm5I6gyzpfZEn0whZn9yloVn/JQ8UjJ9Jj45TzalssVJmK
s+4/7gtuBENlpn2NfTqWJmHY0rgECvFj/3RA6JMLwpJYG6Hf9KJTablBKi7NfDQu
1fUV+vUQ9UtW7trX8azzLZinvsAxfzcR8pw+yj5qVUTUDmRQFsQfac8asoOkxIYI
ApoQwx9iRPyXy2QkyN/bm+ENMcP5pHjdLD81b1pfYfyRzqJeTR2L3dy4uLz7V7WS
xlB9rTg5tmGuKdgRsW5O1oSP9Rccpjci+KKS+n12Wx0iMpj5t1BUFf6WzFwo8W8w
LD2fhRpQYpP/w0GhjDIwVEK/RLShFSfZX5vIV6DQjNa1gOppAvEwo0ZILBx5aCE/
vD1Ln3rnblbDDl8qwqxjQwn1U0GaInZhLAnEvt5h+rWCZ1H1N2MdT98z7VZnB60P
a+caL5ty1MvclhoQsEVz8khr/uHpdv2tURGlW9hAiAMJlrqDN4+wy2RACT/Hh9V6
Io8vFUjO27EFzzSLE25VVI4b4PF/6Yf5aaaO+gzHnPbDShubCxuhKoOPfrmc0NOm
OLNqcHvtKrZroWr7EzXuTouHqdrjxRzVxKL0DjHVL/0OEhcPgFuonab+bN4sUVHH
1tplsD9czZQdsHvBw/eR2WJkZ1dJskHBxIxlSDcPYTUhHeChre0ObwsjRwRlRhzn
hX7Sub6whA3o76+09p92Qu4t2SXSIp25aWstsvZcm7RN+7ixvzTCKtjt44xxCOm4
IyDEdYliXfYL5EPTdpfl1KBMJiOgAuLpwoLwXwc687ZIj07vg0hgdheEXYpeLj2h
9KCJZCxzquI9U2evxylBTmWf7erJi0XO3+x0wnzLvq5cCmJ5nvQWgGWDE/joo/X9
/DZGXM0HECb7ir+EQeTRbK6R+e95O55c/ULRnJZ+Tb3kk0KNm+kJROFz4cx7V77p
W8iYX7B8bVC/Wbsd+HCuf24H7PWKAcZpt1ZFAqWhPCMYcobTd82EuwiiWKg7sX0S
Txb7/hhyGo3otWVW3JHQMETIvNN+KnTjrpih8gakmrHfOEjiW1ugc8rqiOLHVOmT
7pww4KTmULKcrJnx5gcE/cmnBZQq+vjp8J2fBspW+DtzzZlWijMTG4o9R+D08nuT
DgSWPgyCzIJ9Fs4an3FAwpZXu/QLNVk+NQRBsucmQV6vV/wv4Dplm5O1O/NwsXNc
+yTQC9NrtdzxH8d0lyRizpjp1fFjzu/QiNY3gl8pC9/QntoBx13BPY/TUktpUXLZ
F7N2RtaK+61Khi0J4vZ2DSEQO6xDOwZ4gDlBUt9rQvrC1A9/XqjsaaoHpYpiAXS1
7SRCK3nbdhoIWkl2wNd9xx1dn5Y/zVtgG7sNisK8tEN/wFUNEvRHlyliJ+11FtBt
VZyQFMGG0jeLLrcVfnBdNDYu0spD5rMjSKefSA1g+RUJNufk9qImSFkH9kMQOd0n
2oYDVAGszA5lroXXzO8mBccBYODSwgWKwd2f+CI13eXu6m6VaChAkQO1Mfm1ysur
1Apft89/k9XWf7Pg8PzgOPiy88ue2DWc2pmbfeAFuGE+JzERzsK37FGt/Sb3qpD/
ETaqj3JLkg2ClJKPlCjZtLZkt+F292Ku1RhL5k7KfC8602AgMl8fWLEs0zUt8QFW
FYywE8hpVt857tjpHaQbZ4bKZpLByl+qbi4JH18eDmPPBLLH+X70L6QRBZvoTcmJ
3bqkToAJ8QRl1JjwZILC3KqabAbqvinEbK6yO7VZs4rE0kJP9DfaF5E0mxzjBfcR
9oazZy1mciWeZalyk5xMMbp77t+1APrfXMJrJsx8eHeuz050R8UeavW6+zUaF3DG
WbVuacR7Xx2ELIYx4IjkELNomqn8u6jXjFu+bg6IuCpYRuI47OJUsVwlkOM/mNU+
ZT9djGH+HD+cWNooJ64Hw1xt4XQ1/h+XAyRx2/0JODIZQFIgJBnF3DN3nJpyK0Lm
JBu9DfOnoVHaH0GvaBuD9AqnI7fASrQv9vTrddAEA9xaIhBy2PTITco73dCEYCK3
hlngyjXe25fMpzeiL7GzTDcDPLejghm7tj2Id5e1eNEKq2Z8vIA9lV3As64d7F9N
Ph0jKBZbjrAyCV4/CoUeeBrH6p6+xiTgkni/6RLyYYAU+Y5x30sdsfp3fRRp0CYI
H41OJGdbIk4+8hu4dw3iZ5wg9ClGLKgVUCpx4j7cTFKsuBBdcy/mZqHi36m3A2/s
9DVuhXNdxLyJJ8jyGoVEqzEfJ98Wp+SEVlzszV92kM4ZTEP3Gd12IP2tzo075/2a
amUzqzMwjyLVv8B1wglpfuvWHKlsntl7hUpVqftyZBEXTYgHVup3MqodYOHm8hfm
cD1YprCJyV6Qey5RlETFO0o5W1OaNXFyhEjzTHQUeG2WNaDcdpWNFX+Ta1jpBwaa
VrhEmhroxoEWimWXnF7BKO3lSjXtLNVV4pzrUouxpEZmYwjOzpvk0rnYct5SBx1v
c/GRqc983TIiVyLXUlbVX6rhR5M169jFZg2UfHTbeQM/LI/vQVckGDskPr+RDml+
APEvmp9kBM6tShCYWrIM6b5cLJCgyT5FtAxeSkHLeCjwMoAyVls+VvsaN26HWs0x
Tvx/84S8aaJyROOQ5zvnCtJcxHBq4OuEX6V5P8/TxmnzrPOPn/aUFF94EAWDPexq
G0tQXHZyUJIPhGzwAkSEQGlYdGHb5uw1JgEOhm/vqk3aGPUt9MX1Y9wBqB/rwauv
7HEsxsR8RTpywsY/jHSz0ny1eF9NDwlbNWu4I5kit45WrYVPfMTSc3bzwHFV6zVG
VnJj0Nxi62Ut8tH50LrkWjET7MylhK91gGn0QFVzavciJ4r6XrMAMz0pWxpQdfSU
epNIrAZ+U9E/mgDwC/LkgQGeHEao/Lf3GkwqJKtQXY7aGjlCUoeYhKeceU1a0OCF
mt9pDwhNyp16XQkf7GVdoBMHN2tsCtT9QFnpGVmSAg6mGUh+1mX/t9YS0prMMiqX
GcPJfSLoUZitPE4SsFnauSXajXZ58iZoMoLamiy45m4DDGreErMCi3Lh5FSvUU6V
wvLxD0OAEw3lwCIXDPrgdYPBcaI6FXSZ+9BEALFn3NkEWblmhkiyr8YxoFs/guFL
i/Gjn9PWURXiGvYG6s2hJaGQDR4agM9C/2byJsVrIgmprmiDCK2F9kp8oSJv3CsF
JXTHHvUXX0bddexemnnpW1GgEsdtJ0Y20jYwWtrCmEm5eaEygwac+dHOFFwZbOZH
7KTsoB3B+SdpwEdycCeXbh98GrMjhvQI2kSXtW8LKNIck2AJm0npRWBhf1y8LrOP
lsP139NsPiwehWVug6lP1aOw/FYBm9u1l+vAXVr5GddAmewKLmA1vfF7aP7PTItb
fToUAMM4p/Rg2/2BYfu+yblPugBTW25K0ujcW85nHHzF4syrbzNWPXc8oKWNEHt4
ZiVK22luspMlrjOdXHQIUu/mvnzEJnFfsoItMjeIrgbmbgZcQTD00E7j3nag9SpJ
hBVMZCJR6vSAP/eNrJwKfh6ke8zfzJw6CbIg+R6IOtTAide0j7MXK5Aw47AFo0o+
8n4eYh1wdIrYNJTYM5DrsRyI8FBMuYPf8BujwMPTTdYxPwsgFHLH7XB702mSpw+M
3D3s5s8h7juQob/xi2U3CcRMiJT7MnpuL8hgEHgIlWwWUdDyaKLJQOca8pXdhLQZ
KbN5ilEJ/nvx03X7AfVMMU1BD2iH+O1Fy4hMksxNZRG/h2b3HNJP2Vdev1PbTABp
C57UTuY5AFe72Uz6DIGF/BNI3/AIFWotTwaIHXFqcJdZ71xwxolUEhZNFP9Lh9UQ
kCNnthnpxmnhs8PXVuaMZseZaYrQrkgQqMibgyEV8zUSlp44vyv3QVnLVyogLuvY
XU+ll6W9fSkDcYDhrSLses5skq44el5YG2B54/VHLPLG8BerneSkkflNig22G/5I
a5XPVbt5CwZRg1Qy069WsVkAlmMkKL518adfSjCoI4VqAWs7NjpdmJJT/iMHUOe5
139SefM21yhE/lCMKCI08/zJugr4MhymwgFe0OakuHB6/3s3s7hlnxYNVIg2wa+/
HOay3uGtEKwVvUPFKlw/td9yD6lYkTuWZQQp3rzsWFAw39HIGZfWLosotKdh8yhM
iPqstcgzKkWuTarChd/N7BXSMVijVBYnu4cLll2xZT2/2n2ong67csHo9tFuTa85
0/xXP/Xn0ibeaCSCebINtgK3r6BOo0ucZc7PB7mmIMRCz8OAyyWDkO5j9UzwIZh3
92axC5YSYZs5zOBoAhXM1b6E0Hyy0TBLIpX0YgGCEvvjzu2HKvkBkdtu2JEF2PVx
QjkXU1Z6hBh463Jc2MEgvIlSUJ/2Wpvh8e6nY2q8yt1QoOYRTN9eTjigbRAkvgAx
QOV6k073ycae5RgMEU9Rjt5pN8Ygfdm+VdKEqX0vaRTBmPe41ZtX0nxm4ScHlFIm
G59g3oTOjaBs9b2if3VSy3LTrkjtmKURAEjIy9RjS/EqwKTvSUm0bGdwT2aNlF0j
WYBgD83kA4OHVP6DbMoKh3YMWujfrLUbSXe9fsuKlS2o2NH4Bxz4ipjWkZFjTV26
1RNroDwq4ez8anTbERHDemTLA/DUuKz5U31p+WvPay77+TWpGhefPLIgXDRMnJs4
+lmWp+KV5KT8QXqyDAHgLvJHdqokSPoV+EDa0Jb6+vlAJAuOOwdQ5alf9XIo1p5T
Gb7VRecevUJRAhqlHe+ty/J5rFni3FCDem/+dTRfBdqh7falaFtIpeVDBjyaCEIK
NLgkzqmkwjl68fsw2N9FWJmLqXU54AV6+V6bU+n92orZVucR8aIlQPCKreL9m75h
YlWQoc/z1pRwOvPZ1sEv9pfhpI9zcLAmOXKlSnGVlPbV1l6dIW6595QftDfFToyP
V5PVWBFIN7LVqaewFO/P2JLNS5o+3w9dZ3cPY3nSgS5DJu3KU5+qq2DmyvCNRnYO
U0ROxC8PbE8afB6PKa9hT6xuHh1V0j+WI4ao45iX1EZP0I9nWPgbVsnnuw9Pezcn
0GBJboaI2BWh5l36tBTVHA1Q2YVMILVQzaT30EOMuphuidN1vUbLoXj6LFoYhm2R
FmGqcLQGywxXXdKKD00ocOIxU5OOC3hCFUDZQTTnbMhu96ghuD02frVSEVWh8dwz
RW1Z7ZZ4fHIzKYvrVT6yfxEFI9p+BPomi8ki2gv99GeWpRipO1Hz+llQjw/glAIR
1jlompr8LpgPrB8aG8QMM5/EFMDZxXto1Stlo3Bnndug7x/M9ajNDg2j6gWTAjTT
RjcIR40y4URN/p9D3eUjOPPx9c4X948gDcu4GEBcMlRYReOtFlMpkn05XaOmM1kb
fwcdJmcbBNylQW/Gfx2aAgxUteJeHMhkPGxNToxeUMVjYzI9NY84u+UwBPsg++Qv
VJK7iLjI1bwjGoHQp1CK0bsjqLbKQzp1t4KjQoB28JA0o1ZSqxm6oAfR+A5fVZIz
TE5d5QGl3TRPo+moq3jMGc2pNh42pc3s3cLZiesbReDVOVqy+AXmN6eUCUQ9urVk
rzmufoeYwEknKPyFRRHbDbdvgHqqzou3FV3dJzSt3AemmTzZ/brl4d/Nf+tdOr66
n7IMHmP5gp/ZjJe+lVRdsvl6LHgAbyiUHDLqPuS8dFrlrPtu45U2X9WnLmcAphSx
fXDoe5m9WmXMYntPtY2DEEHzha1pnJPD/aHZ/MaLLfU+FBHD5C8HvrARUlItZOnP
BI0ThP7inpW24YMZwfCvqCf4Pod53MpXqO4bfubYYSUZ3QTbACirvTOBCzrLQ4JV
BgqPySyFxiplT7MDT78C3C7fey5LacIqDPrUB8hKgvtq10ld1vHKgy1k54X2yP/Q
3zvw9PXm4azUR4V2Sj2c6tMxeWSro15XxGdzNKc2cDgQwhrzSnXuAgvtXdIxG6BL
fu+wg3WdvueukUO7A9Wx145t8xBnYOVt0o43UV09L1x/iTOHnqsPA+PqAceRIBwg
tFFaa9AHi/oGOyaANhPmYuU9hh0ycXQqy+dMM/0HMBjg72nqkagxjRlIDNZWJoc6
6v/guGjUxBB/ufoleI7oi93lSJ5wNV6sxiCehwCaLCPt7jRCC1l/HtrbdIPHDzC2
6K+ZBjm/QYI3+7FZPOe4f2MrFZegEqOJOtce4w/6LjnTZWUhRqFgaPC+wWvDTGgK
CROCf2H93JCqBNpy/K33pqghpf2BhsYuFAUAdHzJmjvBBlIA339oUyQDooTvTvEJ
tFIxMO1GhdrocgdN49x1loG+Astt9unPIx7vSfiMUY7Z6ctCD87V/FUzFn3jaqYP
jPC7aSsLr1TdjiwTjRAgnQkSZ7CRg9YBw2lYT4Kt/0B2AdQaQ0XcnTFAIVzlAQ6W
RJ0rHpTj3RylCnRrxVjT6h+xPX6t8nPsaG/WLakYCg8s3MzWiFT9TjAqhQGORgsJ
nVQ2Vsz6xGJi1wEBW+mXvR5xxZoflOAIaqBL25EI8mEYftL5ZRnAL9Afc/7YzENj
1wO7w1XfcKXXl03u4D7PTYzp6P/uC61n7azBQoXx+Rm41eJl9v2iGkxAXFtBJBlU
1PldNhSGU1m0o09/hihCMe3ZWCMA8ZcDEa7qLWbT7Zqbb3e45iysMXh8hde3gMud
qM6Hp15KWuLH/wrlbqmd+0t7olKR13D6FOT9/A9umCn8DedNk8J4MmeKfVngAkZW
/0rnw7bAwaXoAf3d5QF/x51Qso9hC6NIcBKvF5ULIKhbmK4nbT5hjtbIJ7YB6bg0
zfWyfIlOg0gUUb8PVTlLkZ3hmTv9bxHlNGbgfwKMJUSp7ZGK4jjO1iiRKeaEwwIu
O3Fv4tH10StmFBVXDUakuLt8R/vClkrqRPopjZqvJ9IXbkUiCGSL17MPPr6dYBJo
U59+3rMnTKoVsG3gdHrLzCTX2uT2p4T0sJOVCiVlrUfsHqMxFWJKUUZkLAc7U1ak
UQAeHwQ53VR5RcN8kYjloJCqr7ODgpPmKfbeW9cY+IN8S5zyJ3t2h0mBfF49bpVI
cuWpqEL5ZkuAkUsGmNVlnuyoiL0txCQ9OQaCBIj/Xk23+1DTV7ol7F9YoRkrdHRx
xlRCPxs0hb3RBc8KR5ZIetVbgV3n8wABU+1pDz53Elx1o7voETi1iWgqIcsSYMnz
Ba3XxxbLbcU7fM1I7hIe55Z48/i5I8y8gnFZxmUaxqzhjNopilGjBIyv5zQq90qa
ozQkD8I6ZQn9N9jYScZYlRPoQq6xKN9AcFYiO2MwW4k+qSlh+ThmNtQZXz7W6ozb
v58L2wGKEp/ofeF9CMNKZJjevW5eujK1kU3eIgkp6ie7tMO7ItY7rM19G5Vg4O0H
a8h/TaGaEmTxZQmdNbxZszuywtTed0WUy4yhdWn+FWRJBdfcZSPuxBut5J9o/95V
NLThX4jh6/WI4PK71XKYPKhlASD8a3pCY03ULTq3hcxVY4XtYmEO8EJ3arrcMmHF
aZNV+QgcbGO5GhfmSRPaOkUTeu3IvF71xfn6DgrRcWebCZlJnBu2dVXcx68JeqkW
rj4gLOlomMVUEA2cBDiHsroz9WmczGztKDIeBuanZOWp0ulXaasMY/eDkZKSu5n+
V06KQh/F1h82w1j0qsXSrOus+/siuWQRdgAaTAFYOv6fayS0T4GuLrE5UBEVKx54
aVeOxOaouEk19Zpp90G7iV51KTZMWyOjPOkL1XiCrhdeECAJFFdVatfMb8LPXTUg
EBaJ3Q5637U3U7oNO90+8RE4GTYvDL2b9tD7UdKT8kDyr8jCLalLUrVRkbpuYq/6
lFKQIVK6UugdaltlBz1r6gKXZORhW0z6QAL7mkZNNri9QkCEp/7CY0QpZaYds9eK
kPaDGVZLo8M5anmQEpgoCGk4GuSrLxjwBIztWhhz6c9iH/uBeJEcZ2gFLG2cFIXu
VbijPvArvSSWidY15EyWtgElH2KsxSncxEp0prvE4922mEXnnnN4TU5mrCC/8MBC
loUV3WJm4s46PuNgnqlxNVQjVcuozzy8wpNQE46IiLs2cugbPrOhE+QCvhimuZkH
HA1luw2YQ18+2slZZiekSBHzTrRH7EcqlzMxIUsVuK3aGrdImM3w/F4y9AHus+Kp
FrdYreAwaJ3Q4J+L+QceUUFjZ6hCvb4MjtI7xaKfp6c1Mf+YTsDeejvXeOstPN2Q
ENSXvV6OOFvt1q9vUyJZ+QVNZbylwr5pHWNQK5MKcR/VO72DQGXkZORx/XNtC33C
ipet7kEjxBQAUdnii/3qPEqpALEmuNzDN7cX/DsZKlUtV9F2lHiNaR+/i1uouKvc
/WJZhDX+jnbS8QxL/JuYR4gSWz0vs6tTPPFy/PwfGiswEH6XYwBCV9K9nQBqY0kq
ItZFvQt8lTCrsdzsS2DP2TdHbtTe/zUaP+nI/OGXbQEZeMfasDye8Miy0UyqcUSs
pYoIFJYO2sOuxkKnVLSC6tBNzPoIM9mV9QEPJ+GJcHBP8mWgO0jNMTgUkJMBUVnA
ul7OZxrCYwackbMoYHWNEe3UcK39NblBD6BRP5s0jEfYdUNox3rBrzIB0eokbRaD
MyYSiyBOTZ/2dKX5M/HIdIRRTTzuifDjfHgpwyccSPZV5eyuAg03Zid24xjh/bip
qlqVTpCEm2N15WTFF8xl55u17VM7LdCFN9sZRX+Q3VQU6ka4+Nlqs1+2eEqSZixC
K1hbzDPilFyQbifJVT6WAjKGZOqYJjBBwATMJX8j5FB7BYQ6DB6rGogliKl/U8c4
nnXGAO77hyZXzS9Eu/poAIRkZzPVCMwUZrN/IbMqMmbZxQsc9rK/ACX9SDq4J7A4
uRzL6PBl7nV2TPK024YZodIRZ1fHWQveTrpdWQYYY+sW2jmNZlC5hPk7L+Hp9xVN
VgKHW9dJgwlxVqydA7SrJ/tqun4YeGy9eJq8LMsPF+WRwBQEEliwn0YztVmjCsPN
vfG41G/3cpncs2qNhUrMCuctwh2+/WcCpRydovhlTDfdRuOy4uUss0EQtnorZ4Bh
MhFeKzVCPNKAVSuDLBDjEp7nzBzqCtTFM5npv6S86p2jAsgwDpUbD4Gkkt1Z905+
wavVcfGkj3YVbxHCyWBlw5nw4WTju+9nDQvGHj8opGtYp9UIa9braCJVs7ULUNPf
/MiKIz2Hm1cPWoW0YCgK+mG2zI3aqeV6gTskYRlu4Yd/dxH3qGaziZXikN1pqehI
3NjNmwXqfW6hpvBaSdd4mcMod+f8vMfJznvr7SNCCWMPbwG2N89rVgx7+Oz4oXt6
64dpIrqnmUyBSN5pmtu+FB4yKcgBOYG5+NIhwuQdi5PMfzzZlRCzW3qBAKnazV9X
PZRBCo5+uO5mFSGtNiamK2ygEYvayVvTwTKE4X0o5n82Ajb9mj2YUHlwG/NYz5JB
ek9oxRD2CJgkr3DwUnAXlVoMvFyNgNPqaEn0r2fkoxYmH1+R8TMD4282qOdKiT4K
3SJ/EkPIOwI0Vl/YTiTZzyZ8by8MZ3T93x/20ixLhHyqy1p8pwXEYDp+9qKNT9/Y
FSCgmGXk/8fqkU+uEZt/VveBsGr4a+m2sL3aSkFIzzjkGbFqr//p6RDsQLnras2N
8cW7BnIKXIHIyqfbQ/jMPxxRuPWcKOhIQE9mFwYQJI1E6M10h46lSuUTn8xNXHEQ
2hwiXV3IykoncImITYr93uhOl4IvsLQVvBczdU9XNkFo2PJAZtJzSgB5UG3bZWrW
vVjtaZvwLV2A6ht/AWef6u2bdAsDg0iNMHXETffzYoVQiKHg/Pu9euK1banz+fZS
L+RtpaUMoDcQxpOYFkUI+gpOhr55EB3VhzhvzAu91XTqXuCM6CsR/Ve2c3ordKak
+O+GxsGKOUcO4ozkzvf0vbyk5HJWyFwTIFtr11SuUjojgGBs7VSik+Y8SrWhA+TQ
jISRUS76MnfK6jM3lq4OzLTg9duitFOI7UZF1l313VlCSRtv2xBub3mpFFTrBk7p
cEGEzGgWJRPsl0XHuX5bBuf79e9WHog+vDZyg8X4fMcyoRSfKLi4xfE27dArr+b7
iQoDJKvg4kRynqTWfVPC9QbhADbI6sEzBnW9ity8JIXzKdb9SmbI8S5WWHAqawbS
TrrviiJ6ngDkvrFfBnPHpBGQfuvzTNwLOfNpyZ2MGpqJfwgj73+w/Da35VFEqNv0
gjsP1HB8zXQpJDCCO21jgilWqBbiBKjt7+BCVxLUT5gxHQBoyXk1d5xmFyA4gZ/4
q4xmzTgUjgTQ3AKpy0YN/CnwgN3BQHSrxMvZRA8VyFYW4uBocC+/fQYz8WeD4iKm
SRcawQy72brTx3z5Ii8UP/P6yCw0RG8Nbr2wX4Dz3Wbmd12YZLgIGbAPHBEEZGhv
EQz1dw8b2Ux8U656+0FDxxx/Wc6/0WiQ8Uc4Y/2ML22HtzalGMQi1cQa3QmQZrou
yi0DzdmLa/w7gPKs10uqLPIGn8DSyoBwf1pwODj4PUi1NAebqIiJUJ5v8ZZED58h
eKTVHLJkKVgQea0hySoS6QLy7C91IUp43Byb2D4FjmKexL1+x8ltNnKXBrfms+HP
jF79jaMs9TxY3cuDFHRirJC4uNiP9zK6Q3/kZGVBkSLoNQVKWAbqr9mKrcdul15q
UqHrpP7i+HzLqGJGQqskBCH6QLaCWo/mzpPaTrL5k41CEavVu8blUKDpQCpYfvu7
H3hVa5e/I8DcTEaY80aynRLI6xm8llu6BDZvfJw82YwZiWLwn0h/w2wqXUav4UDy
diUX/MWQaY88h0GGY+LT/WDnyILC4lX/cVScVjC5I05Iz/pF3wN+Vh+RKSUO3JuO
KhJeMlk7MUhrbVoIyBVZ+Aq3KsSQRo5zkwUm7bxgiJkm+c2GnQNREBIfeXrLM9B3
noEob9pLi3O5094Ip+ofLJ/EsQp/MvYZctOqDRNYdg9EEk3y505Y2y+8gWJjChaL
D1vRF9hAA6p2GvgoKKK/ZVLtdKLw12wBHcI1l3fRbUks/2MAPMYL1FjzYok34Z1z
Pe1ckhUUV7qJA2k7KJymFS04s9Of4zaf7ImYTXGNcQGsMXZQOLBWdUJ4t64aPafc
SwGwXAnDRoH8iPtPVcxiQ/xywhu0X/rFaiga3UT1KZIR8qHtMh226QVLXxGckTr6
6LQg7Eu/aCG163qRi4v3UjanWSMNT+xhkN1nYhye0chNV5pZ0uiR1yLl3K8ePOvb
XCuxcomDR9fYeHhf/r2XClIe5TsrZOZVRWpjeH6hYG/TMUVq4WRJiKjHzE8dg2Wu
+p/2lsFD+nyvttD9P6JakXmVllqng4Q/YNaujWZBKz1/7YMLxYIofWqmCBrhsoy4
NpPbFy9rjY3LMU3T3+GN6MNs1UBRtCAgj143jWnWILsE438DObfYKCshfnLshXbG
bJf+tFNLGM5ZpiaMb/GyhqtT3B+zUUsyNqPgYY65KIJVz7BDU65YHg23RJIL5zIG
jycKfSVNCNqPL0otjnk1cBM+9DV3oVWDiaJlc7pORlBd9+bAzx2AyBAgIXriHedU
MJoRXkLdk7nFF9uRZlY8z3QVcMwRYNUcSUPA7KKbYgyMfkPgtbM/LvBl0Ml9wYu3
ISrDfeJiNs9xy86ovrCuiOGKKLnfDwHMJMeGKj3HWFTMHPBad3ADV0hIVnrCd8rS
eWUUj/46zy+Io6HruLxQCfwDy9tw6QnLLU+XwR2RpkXcB8MZ9cRZsGGAec2rnQtp
ADLcTFkBLgMmAQSzS1GfMosgOTzO2gz1Z7cMmO6CR5sZpjAxbEMma2rehOFjDkn4
9hlQOojS1ngoH7BREZ2qTkK4xEFkWmAcCnv3zvsSeIoVh2mSRAmxNu0KPG34D8mP
Qvc0o4sUXStu9AZSCVauNhdhp9+/WW4UXnO6/LOdT2r6Wy6P0Pk12nuo4JglZNZd
Ny/ocbRcQsYtwZF/0916wQcbdMg8oK/9GuJRZaqLlJkN2m7OZVTdgne7CYbf6eE/
PRvFehJq0NowqVt2sjoitHtYT1DL4aZxXheBUdWwL0lYiP2R9bI9u32udZplTOok
6zgtcXrH0RQaaOpMzDfVi8YWRF0XpqBFkEsQbEhq28X60SQ7ARBXjZB5GUkuPGyG
vGDw3L21D/EIXGJqIkVInwpsMPj9JD+s1uZDAg8B54QlEtLvZZwNdQ2WeoKb3/sD
MbR1kG7HsWkNvFp6cmA1vjFis+nm8x2clX1AI5wTts0LKv8BdHREvlQxXJhP65x9
gDScJNc8lVeWvq8DKNE1zQzv5Vq13M1GfSdbmzagZb9+S57+Hr3FoHQDl8wm8fhk
BLKYvtj97f32rt2JbsXie9zWsTamRnEXqjur8/EzV/+8/G3GSoYYNrj0V81zat4h
GzYDS3UaL9giKveCM7+k1T0zbAniP1O8QKOZIMeWmngMpFXXkEsODvgTLl061+Cs
4DHr+Ib9fF1076dxfxceMbrRj0fs6qkkvSwQNt2kMU3pK19mDMOXdnswm0yxjazX
exr7QbJPxpnU/ai7rJhcIRShhXG6E5T0nk82CT5oQAH6nNlre9GNWFxV8IjAsCTz
ajyjk88ovZmCwfRDJ+CcdLqcDHiASKKoMZGCHvnR6gJQpOa/lLbhiRnr15YBARXO
aGpl7NfaI+mU8jlmZ7Tz+BXI4F7Omq886/qSNI3MTf+UMNNbHNI0gAz4RQW3Wo7Y
Z0Tqxof6r+K6BgMLN0FZY9lL90aJKCoFSS6e0vxHkMFJOoT6Znhtndm5yUO8j0BY
Fu2Sh2W//8cnfDm5n+q+momrhSZnXLXiM+blCFN21h9sK6U2N+XNjO/QV9xBem5V
Lie2eXx7cJ7qTAj3CByHnIxuSDi6WSulCwmzgsNl524JrEZ/lS+8dSPsivVFo2CX
EGYxuDg5DDW/xwkdvogz2xiZrxfYtxgzA/InRe1s5XyTc/5VbXutKf863WDWsJs5
RsGSUSa+MyWYAYP2QAqBN5sUGDv5MJV3OrP1sKCod6Egp2+KZyORgoMXQJdj7mCB
bKQOJdRkVlrMcjH23VBCORyG8iXGl3Gzsrha73WtV/hDmenAzvvEQzrdghlDneQ+
Lri3O/gnPsFhoqd352Zj5glADoXMkWoV2tkEue46Sa2twMZh+x9lGNOXRSe6mzbb
BUGi5VKsCyCnLvqqItHwR/fE+EKBniQXPN5TTljQc6lT6ZTSpIVId0MIllZSbZrc
LlafpKmjHYV6rVDiAFXgrWtNgZFUkitk6legUE6BtIOtosYe5DZxxxT9VO/f1D+g
5xTmDR/ibPPo9z2o4vtGKZ6pZ+7KXUWN33w1WX6fo7obkFsIWSS1XbfAmg7vWTuo
/1lZOjrMTPjEzJ5ErOTUAxWOzj6SchZGGrYa4DGg+FWynY1/a6+RZswaJUqAW+jE
lAAahATswl6+Ijil8S+a2WVkqOCMt1N34VrsfHxUaAgqOD4kF1O2rl2s4KCezPPY
G3m7HTu0vkt3HC0aA14AFjpxyc4QTmcCcgxOfqSs7oyowWunqXSz1qSpu6707YV8
VAIBdaZAPvJm8T1rxja6FlvgRC2oVfFByMWNVjLE5Rhjw8CA051gh4+sikKjg8yQ
R7aTG73J5Y9XVnWWmd9H2oEja34RcSRMqXJePZmN7MYqsk/HJka8240de0nEz8u7
xwQF9w37d7lTelh5CarwajnbSxPhTBRFEP/En7piQT4VmOtxWMBk+Pn14StirLQx
X/KHzms/CShH4mp71/304In3egDJ0vyLSLq302O8cQGpFCIN6wnYQjcoGmKTjs0k
bHDqdEktUNFwBUcwpH3BrHUfmYYuN8wiZyjOWoYa5qq/gcQjKK0AQO1Z7fRtqhpe
vleUL/0a+964m8S4tEPEQKFGLFBa9XhiNk4R5x50wy0Msf+VivCdf4pFNH/5Xe4z
xihT/aOjhOeXm0lIk0BDGlSoE7msyc8okgdc4rEvkO2KT9OHtBcsBryfA+cQdlnl
fqqy1+9/ZhBrl1fpORL9rfI8C0aoNsoEB33hbERgxIXqaTu83vDNool21k+bhhwf
5/kG5t7rO4bSMcLgyejsfjySt9LuuYT8uCbZG+XctDcxg9dAthYRvW9FZsRkbc+z
Ujo8Z0WIyKrbY5Op5QGKZ/Sons6fNWycp2dWBAe0AnoABQQhaz0C1eh5e+RBIN7F
JRIFAvjgCswDYr1KC+aQQWeh7ONJwl0sKLoEqKVhROOpRv1qPXSOlHr0N0zPRPgG
tRZaj2UYxeNUDGZxWiu6cBYuNd9X2SlX9jewm5BV3XpJ9Pk3jMdqOBozNStDpbrl
/llFk+dLaQIMzr72xnCrXSOeok3KnpGgjsoJ7fwC6/eptxCMBbzgFkZF4xW1FTq8
E5PNN8TqLIqp2KtTUXoAYVlFjEDKYbeMWRF+1SQOB/MgN+ZP1cwD7eYvy/kUwqob
SuWLCsss0X2zv7bq1/eS2n0NcRabspFxp5tV0rFp3BSfzdSPB43+YMg7uUdTQKIN
UOP2EKFvCzD8VE7XCcOcAA3YCZfruo/izJ+INy2plW9YpteHv4KPnAROUFYGksWN
oiBoz8XSebFW7qz6AVj4LRexzBdPntmDt+B34d7mvUJ20nFi6nC2uDXnKelur5P/
voWlkQSxjoB4jnJXrKcPFjpj/Ip34ArL69fDxqbHkf1tpH0jJtOyVnjAy9NiMoBS
y3sYMGD3cjnGDsyoDF5J7GLdSne85kEH0M+lmOAVMiKx52FW5negAVvj8JRntLlu
v14SaeqblE9X6TTATgENcMJROiw7u+icJERPi7FTmYYGAUOrtaT+Ta/HV1Zq6W6Y
5/SW4f9Kg8D4MhPz/jh0ndrz6z5BVcrGm1HK5bVwXnX1WiehHMfh+vbTE1rixOlm
RSbWJJZnoLdyFtusYEFcSeYv6JL87OTRRDQAjfBYzvI77YrsMDxa6vgPgQlBtOZq
JYdtYAC5srmY4inVxwFebhamhsX3mEp2zPujba/fudbh5t5QAcfBbsVpwze9bN9E
J7izjyc+mO/JgSaI8DNDacRA3X5lMdWBocoSJZdElRzwoSdRdxx0z/IJZJGxnGVw
hzHc4nHIPUr0TPEqDrM1k5Ri6UHui7lWilh1Px0hRGFrayDHmjUyFlKehJcmDBm6
g2y3/iohPdOykK1JomLwJcVLb0PMIkuqwn+aRvcM6tRRYzAhF77gwAVSl759g3ys
n0XMMhzZhYJCoP49DA0TlZVLKwXlGWAw27CttSIutQiKlDDFaNUd1/31BkZ5qcY/
bJmAJhCQ9JqkCeaHAMzPFWy2wU9DnnVyyquTweDyNXlBDoraTBWj4K7ZdZUMn3ET
rEhUr0B76m5WM76KFuuvkI8jhRrYW+9vLIp0YbsvCqHKnoZIKuvmPwcKGIUrckt/
bUdnmsIbsuBNWF3fTpgf2caUJml/8mR1pJVnXDT1AVtaGAMmT8bNec4IwdfV8KzJ
cpM//ac2MuA6x+RRwAyESHnhyg7tQx7NI6Cd+bKzHqjJtQbdU1Zv/1mnOoJl3WuG
bU1OWQu0CAoRFheovhrGROFjMlzc8DKembcBUW4iHEZwYTQC16QbcYDQcrnsdGWW
AfP5plAtEKOtjamR4UTLtKTRGwylOMiyi/hV+K5s4jBMdW6zoEs3jEg0XAL/qXlC
HDN1FhWUJ4G2zMAh6WqEViwoiH+7tiGMkx8HdVM1p0jrNq+QJa2oU8870rU4w06B
LidqtApwfLN9l1cG0QzSbnWA9sRhcR0cct7N8llooE2/kpsp5DN5ZItSsuyO5+YT
pTIU0fGbiAuIm7VMgtfMj3wg3Ef4wDLB40HYbi+G71yZWOM78v/Es/+lF7QR5BpS
toDep2jNVcbTU2aii4WLapXsZVMFJhif04nDrrnTURWzVCNkKhQUDSOw9nSZcGjs
YFHSO5Nlt3BfZmfHIwTYkGgzb64fxrqdx4rErOvxesZxRmd1dNUu7FK0kFAgVVtb
IZfo6xxMj0NnyH9QqdGi9FCW77DZ+04/hrGySEJi4TBany8jYrKpACJESU8lM5+4
TBHvcOnIwxJDipUkvj6Q+jwHa8bqTR8hmpNCFLV2Xop1p7ZIjx3eFv0nDKzJXUcR
C0+4b3SsodmBi4ZQLu2IE5B3YPcB0XKfkTP2LwWxrZg4zeCf1BJTRQNtGEj/kO0F
rJDi0aQ5GEtUIHwFxr126p+fTxWToArzc+vPPSCWWo5PlOn7mLb07wXXLu9J9jNP
T/fJjx/dRGkuis3kluRHv/Av3NFP4VGCbvOGlUc3iGSNqlx8boclj2Br3AGsB7fY
u8gPhZV6U3XpNuebMBx10kWO6LUu7Yg0hSlSW5QaEp7bSBjk5EM4/lz4+w39Ossa
EoCh0BZHwaK/BC6CRO0UJS1tQCBEQ3zwqH0n9JodnQuuQElwKxcxSuxDvL5Wk+yc
Sn4tjWMSzKVvPXIsUAHlSvGBWbsN9yF66Hkbu/YpjFvnQINmw08RpUWvUN2GvyAK
a9+m4fR75wVNSlXVjVfPl1Ii4w594ynLEVw3MBsKN4NrBEhp8K96vkrz7kGBN+SB
BOL1Vif6R0cYwWzARu5JYzGywAfkttl1FFXjGZjsJjEP9vju/DNx+IaUS7po9oxX
870xyJG3KVbMEHliBR2OqCH8hIopDuSu7zeUhldnT1b/Flxj0d0tYPWcFifzzI19
GmKoVU9/VKyAPBRDLPadXkda5Zi/4XXHp3YdARxe9fdnnnkHdYENvV9StRv/bbPR
l/6iVePspmeLNuzyu8nJ9yHmCMz/BqtPy6+5Q0rXYNJ60MR73syo2dSfEkxYil+M
mz/hHOefzsG7J7a73VFP6ku4cruI3z8SKcleXxKva8eY//6/w/6m0QyQg810onfy
fQsEFySsPqlXMWO4oUALMnp9vQKwbrneRx0j62b49jfLdq/dJPENA6JlQ+iU37Dg
lRHCB7mnjKIb+VTjjv+x1UntV4tvUz82NBNpa8MwkzQ0hl1Q8xJ5buJAp2nv4opY
GPybBbLoYn88PrvjIEqIaY9F+AkHqZxHLCLz94CJadUxYm327NKdXwuUo9q7ixRs
w2+wetvxfgu9rLAv8m9PzTSxE2FxU1naY1J9dsEQlJrwTAawNa+/EyecZjsbS/+/
V00lhCWz1tM1kpGkw19zYqxQ5K6OiUhriA1UL0sea7EOHESFh3e5qGrjcRYvH5u3
AgYEF07LotinI46j0mgymTGTF6j7eBbmd9fnc+Akd4TZzwUeZTMn99FMp6wSkPLc
jUaVOQhsPHzCRxuzTXWb5TxuPfqv9LfKUwu5a3YwD/LrlpEZfmN6NDoZdkWlfwHn
F8XIlujNWLcO28IS6NwUbh7H0N/DQUyTyACBPcy7txoYGQgRxObpQsp0t4BnWrOE
EdPEgVZAj6zv/XCfpwhQo0zQZY1jmcMKSE7aY4lyEcoBqjw7zBQkgl5SoAhVcznU
VN0+JQahng/Nuyrp4heykw/bqk5WxYoHqlFbqz+oEtZMKchGHU3g8VRGNihsE4yS
ZNDZ3h189xz5B8O4IIyjFI55+pIzZqYaG6ayJ5gf9zxLYJUWZ8M1tG5Wq47rL/ec
KVwSP7coubGaBGzVGaBuKaeeg+tKYZrJZuDfTHvxhq45E1LTXMRalF0dlji+WWz8
JycCmZ4OfZgvRtq2ukiES/FilX+T37Fu1Yxb+iCcBa3A6Cwe54cHaAZpsrBCaeI8
uuMFZP5zWYXQUY0Q406jCUqG9U0UyI6rS8bUFbtdOhMdhDrwxCCibfIoSMKyqzMV
ur5zYCH+HpOlGIpviTgtb7dGWU+xFwRKeSVgCu4XbryD1rusCHNkyihW02b2Cdaj
3rfXD6M0Vmr+Z88jgn2Pi8tM9InZeqJXxIrMQyXghDimcFd+OGnws/YP606akMlf
iLx6J/ugVLMYCBZHevxahp77h2Ks9RTepCvEVFwW4FP7rclnegQ7FCyNVnJF91KZ
3OKjegMy8nRdwpVJTEpZL9JzMqK5CU619iepd0UO/6XGKfSe3+yMF4zXO0CIi2DI
aMJQGxF0f3tivRgZMKxY5uZsN+eSEtRvW9fcqFVu0a7lh26QtLpCUsOzSBfRzrsy
Oc+EOPHIooChpYER4kiZ/0vKva36QaRM2JqdM1rejFRqc2J8gx3X3pjSa5PADdrY
KPTVCIoNPh2QxeWDPZPfto+Ooo9dptfaH3Jp898qKnY8w9Qmy2pGMvZtLnd/EIJV
SLxC3rJh0qVmchYHAbL6rVuzi2pFxqbgI17KJdhSXYDwng+TMXylKDoM13lGjwI9
1NJQotqGiuzCHYaxD13hLl6LoLcpmBLchhMsj5W8LkYklnj1Y0u2qwydCbFw2B1q
JKQCuAjloc0EqcfrtVRr7sg5cS7U3uxFdy38O5L7J4PcUVecikFe4KFsieBRcHiW
FF/Y/yW0L8lpZrjYKI8bfX69rQ/JRrpFR0gN4zvFFAmTGVcH+10nr3KhH/0yyxsl
MBK/a7wrPUsCrzNPfPuqzS7eYJSfLSDVw6GHytDbaOGXtq51qhmm1tVNdDzNZqjQ
e4pSBmntqxKiuqoGkR+FAX+hlIMyPZlk+d8aa0v3W9OdwMg9WsPIFUIjL2pBso99
uBqfOpyXoWMHVGlcUcaSdC/1IPCi+SxosVooePJc5PKL+QjS6wT/RUWX323LSdtZ
OyGP3cU9JRds8J5wVN21FTGvkUgXTDGQqscV5VoRUfHosaUyh5VESROz5JFJAuI8
Tycz5GrQBCzzrz3NV0vIJ8tfYYHJUGxrbnzV7VL9KmqqlBRz3LI67vIFcDEdFs/j
jyDdDZ19b0L02L4CSt/6xrTMoyMXh2n141zS0oCvPwA6EiakrK/Zw0jvKXrjbzGv
2f7g0GX1ZvmuJsk0OPD+LtInd7h+lETLiV5FVwLsDi8y0LYZ/mzMADW52VO3z6xs
RvkmousOhXBeTBLHDENFwvP9p3mCL0ueipOUP3sE6gSPYwNO4DGxbKR2n6Rog7Om
lBGo3VfzdHTm1KKNh2hwbmdtRY2Md+p5qfJRb8SD+GBpIdqBRodFqS/DJx8Z/zZr
q3zl1EhHZ7ovmmfEavSgnQGz2l3El3P9nMX5x89YZ0DStzHajriqe5E1R1lsoP+S
iW25YhynyuWhZ1F5rLiowcE1rlsULJdDaojLtrjGNyU2Dd60nlA/xt5ucrk8TKU6
kmBHJHy6wdMOQ7bTlkwEgsZnTlkkgH5S1eFBaY9tw34HI8r/2ERm5seMr20wy/6D
zBrVVQm+t8TbCEOzFhYGDjwuze+kBDYpkZqKUv9yMLkP7S9IxjlnQfHTyJ1/GaFi
G15wRzIusf+lT9+NX/La3b09qJuWqs+qKA4p+y70U6HBH5ZvScDs3GnagyhiehRy
fmxiRzsokt7YUvrVNpxdGnRMS+aSDyCG5EMmOonsjuYj/HpKi9O99T2Ym/N+rLZA
p/rrNEJ/GjUHMhC/1jG3uhTUyk3i+s6WKLxluZ4A/kUpRPjykRjuoCY30VyfnH4x
yO9sqAWDM9cIkij0qvHGup6o+gaCjPCdX4iu/mNksLsx4zXh1AaVeFP5FspQkwF6
thHbOZbjOJuq5tYhdJeHpUAzfX3l3sQ/O7V/n5dJaIfeAhyVhPjKGRDqdydfM47T
0UXMhPNqICq776TD31slhbwypLjW1cHRPfhitAWPjwM2y//fZpFuf66TxxR4TgV9
B4E9IqxMlgk+AR/XEv6n8P8Mq33SFnJtzGJ+iYrVOZX6MPE0GIsj0OxZWMm1EXQ5
DXkML1n1BxgXXmkGu99wpQ0gW3P25k5d3I2efQPP4TQSu+J1X3Y5c7ym1lojmcTH
upk9ueWSqsEiYlz/Hol2fLwlmY2GgpFBWm/bAnaIyJXCs/s3KSIGB1piiSFJ9+P1
JMvlXkm4qa3q5JeQ8OQ81ojomMMR2uFX4jp7jsKD0SgJ+6SFNRXStff3KqGS7q1z
M3RH9IWD5VKHfLfeVnq9M186l2n9BPVx/YJ3Al4ueL+cschq1QHZniDZ9sQOaniz
ebWk4m3ug0J19x3FCcJNitfXbb+/9Oak6U7yBrJK9PxBDdFmEJw/tGyjDEJvFqt2
FFrKer7CF7CCuoNKvvJ4qmDijQscy1SfVfyERpke7zOPGbJ4x1nOzXJwY4ExX59d
SB3KfW6K1Q7eKqO/D6wAWCuExr7ykRIQH/l2D2sPhDius6ufvKqOj5PSk8bY1HnZ
I2tjywSIO94BQg/g5nn9NjZhcT533w3ucbE7268RyfUDdMtp8WKzmVCfriBETI2Z
WsDtebvRFyR95FhUIHsrnxLPjC6fXK9SWGaF/9beT7SM6SveVdov7G3zawka+KFY
qxxk0FhWqDfiRdzIUni/Rizdf63RhopszT0wdQM2IdcVSIlUXYUcrEheMYNx2m61
ayyXoQ/mbOw4ksfjlNRdTI+mz8M5jkkxn+LCdNPGqOAlrJ21cBmR9gdO/d+Lkn1+
w3aowRSCskb8jKHy7h0b/vwS1vyqgVrc8oypQfHXBiJ/sB3k8IuIi6Lc/TOvoVGa
oQJ+Dko6VVAgT8bV1edRa5XwCLvZ9ZlMl5AaIpfNMYwIJF0LgKVFCW+cRePjia6D
AWPfebhak7DFobm8EgIZ/jGY7FQferaCGy/UvW+ks0qrZkFyaO6kaVsDbVsTBvLo
Zz1uVItpvtvx4BWqiDrpwEBkEKMHyFR+zGyJbG11wPfUJ/iRjYqxOqrZNEXvBaQh
12+/1dW6JUX3N070x6KOYzKQJCi9KUSbHKEMBCX1Ks3mu2fDABlU/XwQpAO8e0B4
VzRQ8AFdWSbJfGA2kjC5A1P5rPGW8x/kXKh6l4pvrME9mrA1t86uM5+JrlEJ3ti5
B1cLuyA1OMFUYTrvoq62X2mNDlGhVpQb8w18qnQH6Df3Hrfze+B/bRBzYBDzkRhp
GOqbJrGLkNKo5nbVQBdkNIv2isZFFW1J6ZlbqDWow8bMl7LF/hNySxCt1lzQ2/6a
WY4tRuMhpj0AgqCNHxd5hGCA8yyC1Q/f05gGxQpPB9ARBtbfiUzuNp6eNVq04frz
xm69nc07FWrL3S6Cx24ucdzTtp6lYuAt1fawKVVRUW6v66xS9rhGsOGvzQfs6ooL
rzybIcgDLU6q+eUWMqMf74dO+JkJMoHD9BFjYwvcZ1MexBds1xYa7EtXl416/Rsc
ls1qmaTnZcUwqM4yEBSQoWooRN3Fl6xuL/C7QgmITL5T42mw+eRFctQHKmqCT882
pU7esIITzfAjJVpvNjlUfjZFBl8mPemX9YECAypV5buqY5fvWievbc+nSxy+at3N
Hq2tS0h3PAzR+SQI7wIy9lJsJsv6gRgVPZ1U8deBgQLWWxvVJ7b7xf5QuyvsF1pK
EUUJyb4WrcO6+4JCKJ1i/Z5l3jD5sVHrpMvG6iHOnqFu8XE2wYiapPbhx4Qv/Nz5
ZzZt+Lt+VBAMN7exQuAMGrkMf83i7wuMRqK97Y/jWjRJTap3xgm8yRxjFguC2stH
pc+H6AVGWN1U59ejKLwk0uAgw2k9nU8QFTT+6MPt+LSUt3Y9fqwxTjDoT3K8qegJ
G9ZurcyzTvM5H1Rt1PzQ3rSsnhU3Pwa3W6gz86UQrguHSjZQiaZHqMh8Udd8UVEN
Zn6fLhguBFjxVIfHdLIAJCqTp4Wqg21YgAWLoxu8G38xbq+MsazmJkrNHQLpGrrf
jqzSVwPhyXAUTvHYUeXxq0GQXUxRaND5JBQjBwnTfHqsW24yJE5KewUb7LtukBLH
i1ktIOae8AHYLJxZ461oilo9zMHtPZpvQc8A+jJfVvStRGLTGVsSLj+gk/Xc1bbe
S1/VZQCIha5SClyrQwlFvSwUWWYTqpVnJ/Mqw+x57pUNdpC/G2FYilDb4xngy9IA
a1hsY4rsb95zk/rIcQJjZO+31nT4vV7qrwwJnH+jaMDCw4qK/4cQI6sH9v1cpVpk
4AuXx8jVZymVs1XJXAKHWyi6m2Hs1Yaj7ivX3dkvP7Wjxl6NTPa8a5Dw6+SIsY7q
tuz1kZbCkHVsNY159nd5puAQlBTV/fBLaBVK2FWMgiUgHRrsV7P3zCYKH6gIK3C0
cdnxTwR74j66U+2E5RANhuGrMMbNYuEeSxAATxvQoV7biJEm3yFgxZZmpNjinKy/
w3dRUqULp45iJawD369QBOjQ/xC1i9eyVTb9JZi4pL0y+TelVSZWpuO16+Z8CCzr
ZyZ+mTiWlTZOaYgTwdVstiUZyIYpLpFTvs8MG2vRf8JLSLp+ifqbvumdA0JUo2Dj
JSCR4cvfm5bGEEWMClEoGH0wy2ae+7FoktTCM856XHzH6DLUq3p9Zdb7nKT/DAC9
+4qJ+mKy3ON2AiuUW15pdh/r6eTo636FoDOTxVj+TnfgZC/DxPaERadNNH+UmBiU
YMou73dTbDT4R1Lvh6DN1/vyAcDUDJMnXlE2aZQX8LoIuh2hGzkOnkG3TGlDU1HK
VJ7BYGrTdzHI9mQQMRA1RAOIDnZ1X4dt1eQOWtdqhhh1hlGzc1PCX5655qz1clcJ
qCFfkIMt5qXnH4bDsb1mbSGQPqMovmPWtRNKY7HCu3NWqI3o+XR+kRT9iHKU34AI
ewfsVmOkNBjVklDtfFzj2/XDhMODmDHanpjED2XsgGn2lBiyPpqcDvdVfVXs0gO3
kc8g29sMny+Jkd8SqX72vQhgM7i4VOKjzc7GfWaT8Y9edaSihJIwxzsbGlKic3ap
Phywgj7WnV2dmcUFfZaCJvXY8rRWtYKgiXpjgysLPJ1elPz5EhxymACw887RPZya
h40PCEyPUPIC/3qR3fDQPDcSFoGbg+TRwQIUmkTcivdZOxPVWR70xVLVPu6Rhezp
PBWG5Mv34bc6UulJ+RDc90m2bRaO5TTdf0Q33cwMuwv629pncQphXfAS7FEjScn0
tknKWodcp3/9qyKqkYcQrWBKAiKkc2NL3tgtzuU9BzV+hb2D60CBojW3boRq2HNi
C8aV7uCcQ+aRqclqdGf8+1xOenjx68I7fiwj5VYYPdEHMPu0HEox0rFzJIZ6LiPV
8omGLsUx20C0B5eiNPryISyP2nFdW6MmD6Ia+if6rmXOu3PAGjtTPSn04x5QyZdi
1NZAG4CjBrIBXPfsUdVoRleV0D4A0KpwsMcL9fmlHXwRbqHe45IoEyiZXn/3R7B9
nGtBN5grnJAKryd26atcQg/sjW0NEAE+Ue/tQ/gn49zJ2YV5yEPv3P4kBlnk5DzJ
dm7cGDVZsrWAWikssQdBgMpT2DtbcgavMhRn86cPmq9emQxNnFXiD3QKeA24U072
Yj9rwlkh7XDRxfTR4QxQgl5xLgldrB4rWAtvNndKBFFAWEdMwvFq+kgQ6umQNkEM
Ghm9WhL+/eZ2JnyJmELOLVC8nD4Jv074TixbwZdyO+diwszP7Iiefk3wMuLx4hBc
vhf4o2GHYCY7Hy2QzsWfFhnqTgDBp7TIwBKu85rOZDckcjkPj0wBN1UbvKYt/xou
OJq841HVXzy2DkG1ThqEOzy90Yg+bF/y8DNTy9F8o17yrl2XOJakWOqORZlRplgB
5EpedU1Xx84IzSvF66o/L4ll3z9Rqu8A5M6dHm98frR04MEFS4uwt7c4s4RG8bVC
lpHmgPg02J3fl4XU/kIks2xu12ZfL1S7ywJjZ99KHaHWLauXPl2z8EGhN4abPajL
uTtYSSUrUGqnGv4uQOqsRNWXJmNn9jLbIJs/3RbUxepl9yggrO1ZAHuhTzNJRxgX
JVlqbh70CcCO/SoK68gRkVbviQyRZKMccPi5lUHoi3B1j2MvsfGqDwXgHs9s3v0j
Jy+RJaeiLsl9aFYtBuTJoWl3zs0ETi+t8LAKPoTr73dUo3AoFDsgXX4FsorK5v/2
ltz3nm4x5ZtW2kuVXYIfQtrS2Fc4+BWcmRV2o3UlhUqi7mi+lQbR7oqabfnH5nCB
cTfZEPPnGZniHy67saDpzOme90ijkxICbcs7FR2df1s81keZjywW+587V0Wjt9Eu
JjeC4oHLlnigfCHeyBvBYVF7NqAm7vTlQCeE9FjUEjm6YToLo6VYPNkyBeUSnakM
G5XS28BhhcHadfe4JxaeVOg7wAt/tK3FxKgesRTK1Q6EVHexSUUGr9X40ETiKkIL
/P/k90dl4ZsOKLviKL+QfOCuFlWy+vaYLKmGciJaL0jT36WNaAcy3vspx4glcC4B
u7m4I+hVsU8IWb13hHFzU9Ya33t5ul3VERdZJn+OeFpeyW9QeVzG0o3N/6gMEQVa
UciohTPlbNL1K40NCjEow0Uz1PjrO6+sYcQ/p/oBebGTckuqT9zo3Ss2eNGvpGo1
nFf9ttLi1ANVEX/cTXjUu4wKwWtyEJ7N/jKvfGB1aKcp0LrEItj7rY1AkihWXsj6
YN06mWHa26G8HD9VKY4vL8qEZImlnM+kdDWlTNpzGyJJEdrxQTKU2u+i9Nx8cWzr
vvh4V8yfSG+mM60F+Lmt70bAt+HQWlLvD2oLeYZDPHmxfQOe/LddHjiwVw9BQr35
EPJvz9/VJyCM7b+34zusxM+MpNANF7d28ZB4wUK/tVlzupWUGHOphxqLh1/rkWY8
CQaMHMa9kSV4TAc6a2RvAW/r3ZjvnyzlbK+id/WBDvnzNE2WCRnWEor/1D9oa3ZC
LHQ568NsoILby8Pqzh90jw0iaHcR5r0FSNEXFJc0oFm6vux6rap9Rtvttuxta0Cg
7KhWKmm/PlgBEOHbQJp3JLjCPlcwGt+8ZQHAR6gT0TvM15bBFxkqVd1JtgFvS9zu
3F5yVvZ4Bftv0l7kFTTc41/Gd9+KEv+lHf7GgFc29mUQWh1nELY5ctqPY7ooBarq
dnB5A3qXttp/wqMzmU9chYD7Bsz6U8hKiREzSuZ+XS6z8697McMOQlBx2S85IbTu
qn+Y2O2Wh/8XPblKeHNZ54JIGwc0GTkotwObScgPcm1CxkfHSKO0l0eejXz4sHZd
pHYLcll6rIznnvhzBxOtWlsU0u54nDaPf0UbFS48fLJXlcbP4ehRf5o+ZIJT0McA
ypQVoj7PMoPHSE71kQfE5/B3AT40mAPg9Idd63nj4jKzvDjT8enriDhZNrISY6F5
esJgDNQfPwuwvQ880M84SZnkj8Rkgji4VzsgoKK3Z3tijOSlU3Qy8Vp+w3yL8+V6
CNdarzhsJgUof/jzFu9wLf4XLqguXvFCgDStkELFHh76LTec/MXYoRQX6IwKCCw1
uH2lgPtNPStITnxvTF/6hRA4sFnorlYxTF2Ur7zH5WQILLoey8pv+RGkqub+Bi4I
80LauMY3mwRq+wmomWWTTtQm7AzQ53ShqT1O6yRBQzo37esxr5PNizuVorRErq0y
tdHzpqTp1053VOMfGM0lb3noUEwplzBJkRKgjsQ1fAS8hXjn2lFBu9IJpWLn2Jc+
6Pl7IyGyMNnKGApUjBh9ijMTonctefKEjsZNQcshmWR/Ek+R/4+srDT1OXR82/8z
5Zq19tdbB15wkhyAy1TiUpdsDB36S3oOlM/mXZoeV01Sgr9gKbdwGrVgBVAdQNGs
ZUXWNyvHen7SmFKKkR4J0YATjPwIkfpaLyL5uz2wUco2tQfWWXs1pLRTshFPIn/D
BuTDn93o9BXAorutfou8BGXGhpqHyBhUAAlAR9nL4jmV42wSn6KzYrIWnBqJP+GM
WlPy7HEZ0bWlUMOIcufM07+0ubm9IHsAKz9tdkS7xtJGBj+dbyw0ciHNqNrAFUZ3
eRtPaQ2mnUmKzxVb3AEGKwRNP6MA2EUzZi6p8Vd8vxcj4K2K1YDU5uWgjlyoa2tj
sRjiG/sZu7akYzoqRDhezfBZuHSKLUeJshjJHYfSyGUljysDm/pzRG70lMqcs3wM
rryLUCaBFwgMCwVug54/Jn35gYsbZSbR8Q5IeUWBd8IK+6gxbLA8l+YvJ1KvgFri
gaHkxsF8iJ3bHcj5cN23VUpX7BmGkjTtbkjsNncYM9HgiwEyHHP2dk3D/k8AXGw+
XWDMVH5JgFvrwSNUJo5sD4tMJk4urlYpBfhgG3JuXI2ziuf40PNTBpsKBVKx1UPJ
V07OrdLmmHmSgUNyrP1ueXbFwt7TxSOtzURy+zvwQT0JBoAAj03TSaLnL6E8YdXa
z+RBmwZiT8QDEtBDu32b05HYHvoNfoWUJ55RMsIeWY1eyM7mEdZaYLrnw/KQHdhR
msFKZMle5t4TtHa1ZAClBLyW1RWampV8WMQBw6se6D+SJtXBRVe/l5XCSTId2g0B
TyFrE5d95Hpq/01jEP+iAcMUQbBAGUZwAylkwamJvjiPIzu5CFSnD/ctusLsm9ae
i3IZUJGturQ3lTqRrywfgs9R6xFXc6qN2srusN/ISerAra9omuHWuAKajXXLyz+6
Mf77u+NzLQKEZYxa3VXnAV8oFhAElbE6dqLtSPytfa19yfpDR3824jIfslCwvJyV
7h1oNillpfIpvn6HiFuVIJVPKVwxYZa9ZyxF3lF37SFC1rYN1xjRqMsAzZFN4TTH
9yJ9AzMD/43nctszz4VXAeMw2cHLdgL558oxQ/o3t2CufwXTpc6KVGTnBJSpYHmv
ws3WiJpFE7YcEI4v2X/i9uML7xrVuKN2PylVxbnzsWesenqT40HXZS0E6Tu/4aGT
glId+BXAd8Wv/PeF+V1wUf4exQlUu6toWfobsHPxUaQ0KK5Nudh5kkMTBoUh8ES4
oK2WRoQazH4tApk5c8CdgJlMcPIgN8lP53gZE7sU8GDrAFPSqrtR8tyGpsVZ28gj
KmiEzmtTD/zT9ItYTPFLDvWyttlp/zLycj3sst79AOuyu7zU5e12WkZiW3VN2ToB
rLpOJrqLykSYj9qE+RkUBVhu1YXKcsCjRrsakfuXZfNPAGZszJJL+lgFPUyBaQeT
tODPUiSaIoZZLMWaZcgE77CS73qH8Y7vhhLwES494xTtfAfj6G5kv8aq79jwjsYb
55bKjWrQpNwt5o+JNlsO5YVVyCiIwQn2IGRcy0UEpHrbL21RQb8NMSkYoW7He9Pv
/LyQ0P0D8x3DnxDZjylTjjQbbAaCmXu3hHXNYGWsLY9ob33ougI4UsrlnOnxJkhq
0plGHdAI2HPimMUIUFgBx7sueKTkdSy1gsDfuAoCQ60nTcVN6dGcujIyYq7jsete
1FP45isM/qzu7Jabbac5xJBVWWzC92M9cuawF1ogTH3hxE7YY3Vb30XvntHqD/E8
1UP8v7FN814VG2XAlE8jGlK/H+655I2C41nHuTSk6HC/BphHUaoXusnvme5g+hY/
g9hCUDSU/gyXqgzwaAmMb4ED4qMBwqYOGEBCJxEmpRiSWjqdsjXTQ1YixQ5xyi1l
Yj6h18J57+wBrJ5h73AU4XhXfYNL5NVegMqGz9/r4xW5kiwaBhGyp6xAgy0u1imS
3zKcemS9d8x/078+j5JFo8PDomWUdCrot2qv9tVAMu8hccwURYOzwId7wyk7nprE
vmibr86nUjaM/eTLJhCi2hhpwztoa9RfyK2EajnZt0/2pdAN5Z3AGG41Qnxo5yGA
hmXxsK/e3PhrEf+XUEInTjLxENCHnMDUgz4b1nreE5/pyXvsWNrxcGxeK+ceUrwM
CW8UbpZtuSxK2ROmnAAbKzEN7MdRJu64YucxtsCrqznBg2EGA7303TfR+Nr25SL/
FUD1hrtsE8lf9nZ5gq2h/e4OwvaNxhIcjI3quNrWtCotq5wOa0/RY/OGwdimaMLn
5GIBxYHedTOsQuBbmB7EfJrqbnwUuqd8h+8/p0T6MSBKWaTGkHTl34D8e9dY9JRd
n/Mw+F5QPpHcLHUwUrdVNPvkDJZB5XEM6/qoql1z0DjmracdXEpKBS6lu9PwQkqu
rHkmMT+ABMy5C3hHTpDK8LR1IaLw5d8SYUZPllHq7dVwEH9rGIYlaTzHj2YAPNiv
NFfwGtuhJJPsNIXMCkOP16bGNHmab3lASHjuVQ0vlTSDOvBrVMegrRLk+zcD1sdX
IOYMNVZt5jplc6mC42RvtZUE0RO1y30PkAHbhXi7R0+ZLQDq61s0N9i9dh6kmz0f
nDU38s+WA+R03UeZsPmE31OUIccnTrwt48ah6vJ4FOdCdH8CAvjsvAhCQlxugytP
sxgDdhLYpv0sRlAelKAkrETymtlwW7+acOYzfUJv/dbjA7AnY4meZ1izzUccoVab
HS6XFiDX5GlVlw8H1g0OU4le+Snt4+hBH9fmE1kTmTVGRS4Cmo4zUpG9GOXbFwa1
fq9BH3rFNgtRLQsccbDiGbiRrd5M3Wusl9saSvPhiIOjYQujmvlJxctn24oWFdRf
LCD+hgsTWQjv3Oa8fRTu/0mRKysJCQ7rmiYnXhlP1e6vBUQ/Ax7PG9MioZRH9VPl
t0GMpwljK9vEhGiutizxCG8HNX00ljpjLasmsNGzFrk5LVgSGYhaQXPSHjLcVYGO
DHzKU838p7LzJsoZ/TlgDBfFER0OrvvjQWxmDGHEEuGuwD0kxN4okoCmOf/mNUHg
TzVFfddrwzZD1C3yWzTUI0sm+J7RHKFrerpCMzC5u3auuN9n0XEkeOXcdj+AGqZ/
PG0ZprN9YGOXgg83P5VBzKEMwptB7IeKqs1mJCDu7uW+TfxS2ucJqWt0EoqITC10
FiPKpPK5k4iWF2iKb0cmbGGiWUI1ebdBNlYeixMxmWF2UB8rnIm3755J85vakkcj
e8sbcZhSGKX5SOijOUByHc8GGbkZAhNRbeI6ckQXeiSqYALCUAMTyELmqLVI2uXC
kV26KjaGVV98pQlSgXX6qyLStglMrCw5A8/klwMXFAO7P+vXrjC8t42YNm5oFkmk
mEwPssudh9/XEouL8PojMXo7d8NNnWt4dsMx4NIcMiU9v/UPulEb1ePHcR0uNRQj
t2YawFtu5DGRaOeoGpKHj/luKTiNO7j6tYv9gbKaHYtJQjYN0817vcdjCEvRAyg7
dIK7aDOFPfkaY6dCs0mhXtt0BnQLYb7D9E/QNSzvx5jK9eac2wfNZNW7MZ8L3qVz
McOPy5l6IDb3hG0kryC53kpc8aHCIPk37FEXF+N6eJBOdgJAtAadqt4/ECIv0TR8
h5pPN+G1u0pQmkgwaSL27VpW4LjK0WqfrDvGR7+iFfmhynrWDIvlY1IONGLNbsLp
wSkjTRw7zHuDZwLfIqNILE02+dkjXcbxfJlajdM+rUoEDGcVeYNFsgP/chAlmyZ4
eTqqZxOMHBMppcW4eBMpf6vzbcP8z9cUGk7R8wwbbiitKSUCVA3kajZOFQV8wj//
w9gP6hKzZtYgY0KMoBokleOQNGO9WscqprgIztUG4zBA5nb3EtypV5Uj5f7bfnXk
DlkTIt0WSL+VKaHnbMLG7nT9JvBGtj0gK28cbhsuUj/seuMKvIMH0Iz5L66f1mkz
iZ4HUoHJNTTPHlun42iG+oWXBCHJRLaCyY4bEZdyvsEAoUnhQxdSO+UpP9NY9pni
u9M0bKn0WS68peQ1nyFcu/XMUFlgnO7XIE0EnF4HaOhOYd5bL/NiuUizVHX7Cnqz
QCdgnezSvT4fDbsz9vNhplCnAeK4ceQ/McxIQTK1bTlbEePQ4xAylfvEjnN9kyIV
gkmEHmk0b5rhfeTQHkSme2rcEjyp9BUI7o6cUvrj4Av2vznakyj8rg01o0ebV4nm
R4LaTHqgoDwfOrCWB2OqGONtLGpL0eUM/MRnacYor1mtdxzFqnNyssqpLUSS2+Zt
Q1cChNWHZOoNeZ7Yc0cAuiLRd37X4P33abqwxbGDr5M2nowvUVuWF55cmv2fiGQ9
rBg9+NnARi2OAjs7qfTI31sXCR1oJrvVgVumiWs5Bi6OJkVyZk6xIDlygFfTGLT3
M8ewPnp1EFnEPQqnZMogs7xFTjOnEcVoaRwYBTunlhcVIpTAfDu7ilDys3UriyV+
rFk/jVBoSTxTzgKeocIvscPkl0iN3ByO/934du0b8HFP2IANL58k/ZglujBDMUQc
Fyq1rQDUVkXPp/83B2tOc6yKepHwC1PUqaWLfVTb4FZa3tVlJ/L4quEZ6fU9eoYh
Etkhrno03bN70FDTwWlLnnDgmZARxBLtcSVW1C637tCtmc4mXr54wSqT9gMSG0S1
kBRQCMqwoj0s3kRzQT6QA0x9pwYzD7u/B83fY3WxIyNkwW3O5gNYXXhgIvmwhNpl
F5ATEg9vUdqzGdsGPnCjgTVx3CgazPAx1qQnBa6KxSP2dNACRn1w0mSEDt8yb1gk
riIP5sYum+xHWMLiJrzustzqnJk6FKykagbdCGt5LumYcYC6Q6HPAxQWxgw7tRGI
Q618osMz/D/Jr2+nFSec1bxc90TvNRqSeeq7Hrj8xxbcf5kHWvcx4vrXLKAJh1p1
zXFstelv337IK9qW8M2pn1fT1kHqNOUSLu22hv2L3swTSh8giKZtvdkiFaZwdPzj
6Yj9MO91yMBjNPVigMv+J3mSrfpeHN06IEEfEqfVANLZq9Hsx6r+/Vss7XEuMHwZ
vOGA5pOFXk4ofj+p0Js3mF1I/DsSs9SNRDKVmGozXz0lZWp3p8Vn9PWfHXuH++89
CSi8KZfPKvLzcqW/R91V8kPZeCwDrMgy9KV8FikbqqIYhl8Ihcy+QnbJcOx23nMF
P8IcZXByvD5NR77QFDurdLzlcjjwDyRRnEdF/k9fHOqBViHopS7SrRomIgREDTJN
cFdIhAHLTBooF4ae2FRDZNx1DbVDVhAL5xuv3xfvbEa6CAlxdCU5BmbNSMzZrnLE
w8K1nevvkzI1IxXLIcmSW1mw2jeDI4FjnNbMMg3mGWNI+J4V0YRfI+yvNdRCnKIu
PTwsgs8zi//Rwd96kV95aqZrEBqSDGdduELkNyermYFYFx1jkUDG9ty5Xsoaut4L
0UQf8rUuy+hhBilED/uViHu88K9b/Tee0u5v+V55UQp9tgRXsSbbs5yJaJuaT7I2
3ZGhbmIaiwfvgsRKXdHAwNAgNvJeFIumfvCdsVn3+/ctuW+t8HOn4XhLWzjuQdeU
zu/VOyu9JwgvouP89mMQzKprFA3SVuUasqmlG1nJmzXsK+2KiRh0pp4FpEhDp5vo
V4V4RzGoZ1vto2L64mNgHteFagH19FPe2ZR98c0AYUHEQTSfSh0Kz08kH+sbDvUq
cGf/DJlX/IEtfF4dwllXJD2DQOc0pTvUfU2Ud0+ze54zJcsblWHmPVwU/fqi+kEE
n8H3hN0N8RWvYhMR40AiI5U6DKsOUYfMLwcGlWpdm28KvEyRyb+6N9QMWn/jSBTj
gsbc2zjivpVkNVxZXzbdeAt3Q1gqDWHezMse9w3uD7QAPh3Jiq5sTf+7J7Q969xT
Wczr8v4bWhdj6pMtXYFwb8Yca4XV5GfKibE2bKG8GXEcDpVlYRU8XWdcMfr8T2oz
RFTObKvg76ccjAJB3gbVOw0cg+98ryU/FDzYgLiFWpa0eaMfFw0ZSoDHuqP6LQeI
6zyX8FSv18dh2HICtmNJXj6nTi93qhl/yFzB1uu7Q+SnHsTgRb6IBXuzNYbsqT5H
TTrcqaAM3S2pHZEaCDpbxmsnOwYrMIrq6+zzsVXv4wakXHEAcHVIMdwt5foZi1FU
0y2BjywSE9dxjwPIUjZ44/HI801epKBa2zL3YOig3PQ8aUNk5nZYB+vtIAgcx1h1
Z7m5ghe0BQr7YxeqG/nTfziPWx01zZvajn63qYAqL5EfLuIZbQ8HHWCNkbUKjxUx
SKJf49UhlljjgH9Qk8WW66MeMLaVfIJ39HrUScJNdrmxr7sq+/tm8ioX25C/pQdd
jGuW3hR61oiaEqgB8JHGAWDZ+ID1YUcbEckB60rfL5Gjvf5EgiJItyicYyNL8ExS
O10GHr81T4FRxlnXQPT1vJ0waJ9HXP8xUoSR+gzq/bLLRux4VGVy2fOOig5/2Ern
NpUJEdI7dCBbLM7nfamy81mmvGuNBMqSTrfjpJJobWMsSzcoNXBIn+ych9v5Lj9c
O4FMv4WL9PORg/KNi8uHwLkiapB1Yx0+/Y/qPLGSUAWdzmMTG/y1EAHe3CmRDGd2
fzQEztj7tcC2MOILkSlQIijRjtaR4Wz9PU3PnRnK6rt6OrPrP6349kb2tl5eom1x
/VI6zCzIMvDSayntSZBo3frSKw+1PWlmZXS/TpgYKUaceIoY5YgefgTRCUErRLya
LoPbVHLOHvxbNI81eQM8IGX2FZrakuf0fYxlo+B/AjvK5U4wV2omBnFJp6BW7KO7
eBUcRqF0NTKNZ3852DgSlNYFxS3oiVJTVb/b41um/Omj+0dPg84bLzp3u9oXe7LN
Cuay2xONNYRFdzdGNsVjg1WXrmnFsK1T+6TnExN8jbsAAkFjxfxJUGi/oYs0E/QD
aUzVLhwDqpL39DnVT5hdQUumvuzG9ktOKnLrbPkvl47Rg7y3gOJI3RVtoWg9qD9u
aArxe1ANRDbmN2IP3tTipBn7wxbKx/96Z4nRgVwh3UMZ1lj6bAmKvyGGRZ2m/XKZ
/7l9JkRfoTMt0ah1xZ1vhAjJbU01nME8/j+jiV0lD3+w2Q4tTJj9nyCZQTJ6vrlr
2HKxzgbXLbVxpjhxK9oSV31T970j/AYlhHX7gi9ji8qzm3EVuRRz6Ytyddl52Q2b
y2SOXHKI7bzXAPPSPkoZv2RfLA6mJFr93g1vzw+yAPnlfC2PVSSSj/qny/D/rMIr
RwsujflhqC9oq90dxFVb7topj9YmfiYcQ6touEB+sNiWiX+vwtN/fpgWCAR2VrNZ
bHBgC8lvxDEOYtdhNNMXkWIga0KNZXMhIwvvxPNH/egod8mn2Ay/IZM25WnLLSVE
YUfP6rvcS6tu3Lh6A1ta2HHAiGwVLz1rt/SkNEb6j7QfMfidJnF4R60hCFATmMcJ
+pd/BqPpa5bfkV50TOjdG9pT4xguR6Bsi89I2NIYFD4VfZuKqj7h6mHX6VFKeQuk
+kwuRPtBiDs6Dvv8KOAPWoF5nP5whyJPupHCrkRRKBQhSZC3wdyEaoOV1lniFq1w
E/VgqaAbh221b5OQ97k4JGcSo7BZaQDz/EKoa2NL7zHc9OFPzgD0dtgF2yd19VRI
4PTEJJaTq3IWxlD32yX5sj8O0IR3tah73heuCr64sagUkltGz+TPq93rL/++Irkt
QgrzAp+xWtnLDOx6hlK/SrEhsgKD1mUZf8VaaQscZ+Rdmn1rPe/rbuwaiKb9mGz3
PEVh4a1lYEUkUwebR+NfwWn7czZWhzUf4CtNrwKJmnKt9B5kco4YhhrnFgJlrmEW
md2lHH3YH6m8qod0Is3hwnpypxAOXI4QZ9h2UhnhYOKUxlCsbCzqxvSSt8zeMDrb
+BVrNGYybFqP8oHOsEFkWRbbb0zt65+mFqcNsHmEGjAO6ScmtDiZkMlw38Z18Yfr
iUqQOtRvd/Rx0M8uVKjBCC3JwdylZ1ZQkiTzPubBAi6y6yH/OW1etfIWpcmz+PCs
tJzh35/8IHXW7X7oOznBKmeiRqOPsYMC+llNlEtt+NdO9RlZEZz2fBOo2k71UbL9
+82bjxogKJpo/kY9FZUNgDpmUdip6ftxkUB5fmOwjbm1fg9MAPoJE7fUPug/CsnK
1cwsCncBmeSQ7cBVoBRNabe7UiZPpIg/Qzv3svklXrRa8MaRYGJEeIM15IEptsGs
GbCj2WJUvRBy2iFYNW4aD69dOtChfoNZnoI55dVmkDkgUQDHizxbt3+wEux9BQ6a
zZKo9jHerdqC4K8b4AHtLc4KIolQx8wi9Z2rxKCuwGoEPuKx6Z5XL3C6FqJNiTSt
0YD41Tol6H6e2yh9iftqLSgtPZQsn14tPd7mj+rbXk5iZPlvT9La7FeE38VgKh6H
V+91r6oBovZKr6evAxqgA72285yTOHli+t5ZmLSHAbKVNGTy45ueiGljt9c+f1Ty
AWpWx0XXJN3XjwutSmMzXIFslkaiILnyprEhCHFEzmZfsPWHuXz0dmUXPly7adAo
WNy5NYYr+CELZPEKdyJFSld3FgRO1eOPxLOuk4MlfSi2fwR1bwZ7exBTs3esnRRp
Abu7WsgD9HShlthvbYPEihgr8lIeMGVZqvf5u0eZRPRlBbSbrTry0e7JvyIRzrHU
HXWnsneGBsNhVp1Gee9nH8Ky16OREVBfqh5T39BA00t+Rf0qjNawtGM87zw87vUi
yGxKMrXWYm5xydZBiwDEEZVD34E1temH3NAkDcFsi4kQadFZbPVW34HhidFWaCQG
6DqyHxvOmo+fOSvxD4NxQecT9RjfGlaXZ3RaS9N/Ro7XCIT2xBVqN7wh+p8aapbr
Fv7E56LmL+jaKgwvz7hiN4bZYThpm+P0KIFwp2q2jdBv4B97jpucB8yjaoqKWVgG
3KkNJX24cdiVhxFYCZtzqHYMRQVGup0a3c9bykX/1PkLIdDd+2ZJ012A2lxAjUzN
T/YtOFyv9wcHzg/iv/wlSJrSGwm/l09ad5xXMnDMwQtGfVAXLlkX0V6dCrr3aDmC
HsA/+PVbmQ1n0W5WK8H8q5UgYZgk99x23PxZPrbywaT0cOR3vF76UPtBBghPAc+b
4ERjPfvQ6T/cDNumxP1WmSml2jVSR6PWiQmfQ/5v57BejCeqyMJ8Jinj7Pj51NkU
ifGd70FxNCMmsgtAOF3gV98W+16ZlVRYBKTP+O7XpEY0FGXxrfutIZF1tUkn5pc0
2MZWy1gNMxJSNcdFEpx+Gt0zLfSe/LiTDsyvHTjGbLNv8Aso8bEChrDcYYrstrUx
mjiWEo5kF9QKgXp4p/+R2+e0N20W4Cml6+piiMcIpA88/yeVewGmcAw6cyQEYoKj
nkt1UGG4rBHCUzsAqbadUfhiLVMg0uoYYgvB1b+EwkznnnmRF6kCw1gbUAzmtGxO
/9xNfWd+A/ylemItJKLLYA81VE7F4fG7xUqMKwRJw+6UZsgAke+fl3KeVpFKvHN2
0UzrB7kPGRbF2BX5Ul38aewHEu135LBbxCvJKEEqbEXZspcqQHHLfSF0K4zhDDkz
AsXhyC0aizGn6YsJFB2EwCaqOBTog3xEeptsc/5SLQEWBqPdfuR614K0gfVgKN9t
y5Rd2wIXGSmWfuilp8xSTxNXcmXGA7EBddBjddADwh4Qi2iT0blAWfTs4TDY9FJB
DkmRFNXpmchj0yzR3Ur6Q3jO9bHOJ/AY06jtibzLNo/4TIsTNoAOAQfxYEWBYPzk
l38VEI45+Q5itXwA0MCRyIPgQO6GnNfH7iSwUACqvnH/9QRp96Toxsp6XJI5JI8g
+73R45Bel4Qk/R93VCPHhMTv8x1wZF4hvVaEd5zvTpWd15t0Z7kNmm3Q4MFe8RUB
KhJmMzneYjn+iF+jNdh1L1/x4TlFXg+aOMD3IFfi736bmgTTTU24L6RzLE283qPX
r3XqfRzdAFrOU7dpmxtAJmO2rkWg4X5bdQ+WyDdzHNSmy58GhFxCSA5hhlSDXAI0
ZPKyAWG6ymkxdH/S40ICR4Quk+FC2CbMdr2MDwxwaqfDtpfOKeIybcCHkVBxVH7B
kRBz8vxPw3BPLUFxHV+VYhrx/fxbFPfX/fBxShEQKMbDrsoiZH/+pO+Fx1cCT13w
otO1ptu8DsHu5M+HIqhLZ/U5/YSs93iM7a49bRH3H0QrxAflPo4oDTCNx+qpHCqv
rXiFY3i1amX+0IgPNxL8ltTl+zg/6W8GcYEBXJlDuyaqLqsP5DJw2t3O2oXi/Xvf
APyv4t7kqqF4HrGIs1pTAtdpMChfFpuBeZ3E0Ply9I0N8VmzZrXjbmmM6ZwSqAuP
6c/7MfvptU5GPS+TxrbsT3sJ2dGnELIgrzTnfBhvTHNVkjVXHEUYgp9Jf7xzx7d6
WbH8lmV6/APRNugxGVWvgnvJNtiDSIRhe4ATZkZms/+sshZaW1QxxR04x783WNz4
fGOgvFunWonCRqr0U4cCdqeTwZy5iYocTn0xeNfMIYgqxRV86J3kkGp4BXOZ4Qbh
AC4p4JHtEYrW/CG5Qo+v9GpLI2ceRSSWrqeYhqzU7Dw84y3hBupKezI9aREQJtDW
3oLXYlYU7U0ETbxcP5uCpt9LVCDkoaJogbA7KeYeI9iuEJ6VioeVruRMBS+z73wA
4IZvlaSP9GCjfMiZMgc/o9G6j/olqONDn9iOTXbthgozXpDwXFRR4YWPVHbS7Tv1
G+c677PWepWanx7VFqN+r51Sn6qwHCVV/2FcuR4JNevtuwkcVikZoWhYTCHcPGBb
gOucGBPDY3dLDvQ5XeOhlTQpgcd3aa+iUdH8OEtLarVDBHgFru+1kgI3hjq9txUK
bd8019vB/mbeenccl5dlvALGMuoSMIu7jNSR22V1oT0tS+vGwXBFiRVzK5zEXa5a
eeYjXYzeZgvJIcOOro7H8N/15d3gT0YSUr5t7bZWyxMFXtsd8d/9ddAcET4BBeGO
Pnq9dJOev66916SdGnnsysQxLzvO1T7ob150jnuRqL3Keg3fCslic5H21T+000LL
6W5Zo/fv+tXm/lZ32S6EqqVC5XYxC33kBrbzdESvm/d5l15WS33k8jPmh9Y90FzI
HLfhUxoylQSmueFrkpD9AF/R2MzdN6UBmEuTK6KQ6KtVDdsK93v22cp45gZcqHnS
r4LYJ9BgFqp9Lk9/8uGz1rNqQKHyKCmSBmvwlpER38u1sVrpqoDjCBxu54iItXBm
tOSnt78SNu5XXZgxbduF7uREG6J1PTJ2w/XBAojst1WSQiOZTxO/DyDWYxf8Dnna
jbXVs4Gupvg45+uMtDoBePlpArqrxLDnKebRvsPs6js4nmlhz+GX0vEQRjX9ITxB
Hwd7OjUhPnplxZT11BPBVjyaM3Xf0MANJl4+T5Wj6uCBICS79XN/hznAkKb+BR8M
t/un1qjqs3t6ghW5hwbZLiYS9FVUtpM0/AvR9Kf05OSNAXQuzSTyCRHo8cvwjjAk
+4aAjPvuWeVm1z9VmIS8yUA/Xk2mOKUlGG/vxhS9iEtzo6Jhx70idSqxrejupk/4
YKVmCUhvnTzwGBAIUcORdG8kS8fQkPeMdxtYZseQ2PZQGoY1P1MhNc+E2lmMYywx
naRsy4mLEgh1oYg2HIWDYZrzeDfHvZ9uxDi1sOPhq6lV1PDyU3y61nshsHnDehzc
Ls6TEBQt0auKCwcDSnvyL3700slaw8CyfxCjrWVYHLf8U9XGj6PICL3Sp+yasT9n
zv7s6fhdS93k7txw/HlpuEjLWdrCGgOpKs0biCZeI30QaM4EmQejEFnJurrCNaVd
3nzq5H4U3ELFuK1mJOuzu7n9sIkmDAavc9LL1n/GOf4/kAwhl2gLDMkK10zoMBwx
v0UueOxarxa25zaK4PVYCClhWkflyeNtAykaf2sksL70jE1beDnOeaFQotwQ/eK2
Bu7sZFwjVsMiAU4kEz6iJicGpuOzSa2jCjaq9rhrXT0ExOHD1Vj5WaZ3zavl2ZcH
vbD9aBmEPLf+4uBR2iMquiU8tCvHGV+/d4z7myW4nzfvbJzd9kQx2P8D6w0nU44t
KpVgMeC9uIhcu3HAE+Okan/V7Gnjo5UatHC+26GVIRjuELF+pM8gkwiUCy034SQI
E9vsM35QGnychoYAGLEq7M/y3QrfzeNV4oYi8FgTs9dMYx1anQuxfKite/6M/R4i
HudAyHRXU6VncP0KFoulRnX4WN6W+DsUKXsp8HiZBbQSZcOLmLFMiWb46DZ3v+PI
kW5yE1UF1IaRn7gxB07FiEY9o0Lq9eFacFDFFH6+rZGHHOmUsXx926lrkw0Cs7eB
yRoA13Gh0GWd57/vLsAvO34jxiUV5n2czLjZ1vZaAJxBdJ0QTu+5+ZKkvqmE06Fl
TzXeRZODJ3b/MCEBFIQOA8v0pQ9VS+arth/sxIUgCMO2hxD1wirP8LDN+8dUaQYd
mC9pw5Sx75xw0wkQF8WziEjh65hs7Jw7LilI8h0/07aMVnuGJu15Wvx0z7ONTlPB
QcbmIoMDr1RteOtOuCVzoEjZNxIkk+Y1z0vsLPCAXv+F3ARrDPW9+YVx519hYkwx
IF4Yd58VJFfRJo4v5y2aK3oawEWOli9tgQhriO3PNOrmv7iaSuLLDsKg3ZA1fBnK
Vdd0jI+oFsUMtQooc2plzZPXe1Va4OpaBe5vXcK3Q2W/5eIE3ZoJJgirVajJTqrQ
+yESk5Pwk5oMbDBNOx5UmAHgxiTVCz9DF712kadxfROMCgXw2OQZVgYCNX4H6Mjl
8YgyQKl8fU+ZoBRSSdLHEDBoY7rWjQtpZBClb4ILJbseon4gN+NyCE5CjxewNIXK
+6HpLDCy1BoAyDFFbEe8CtspvoXE+dtYArPIAzWxLO1P6kXIm1RY9vSUiwmLKSQq
UF30IGGBuxDxKsZpqR6LcpP5kQAyJ4qYNRcmVEQ4Lk0R7YLXrrGO2v8ViJY/da4N
XGm+4Xfgq6JV5Cm5bh6eEH8/ykqURl7RXtK63Ch7bx3sMPz6HLQsAgyszxL1hg/E
TKesA5YofHuhCWFdpVlSmOga5eJ1H1meliRvY3J5IWhtb8w7UYdluBcvN1ilwWkT
iUNhe0DE0Eoa+4gV+1yWNpvt8hQvEumqGztxeo+h3fDTGZq4l4dFPm7VS/vfAlgv
JiQ12QQs8lnZnA1x+gwtRngXEl9BF9eHbG9GDE5JDsTVJ4YAc5XFbZOiwPOILPFH
C/J0V5vjdqVOtI1Ch1prq4vylzjs16oSkhvF6SUcf8oeZpIP8UY6ASUu9nFtDNf2
IBw+WGydjWfvslnb5oLS/F01UW1WSLqSSXnQY3n/0amIJ3o/hmPcQLvEPCP+pC0c
ngGAIYa0jPhZLK/yFbqi4PUgnrF/tndABR/+uRrQYcUhGhf5YfB6eIFIGeU6lMqK
R82OQ0vSB4J62E9soWArHcPzTaKgkKswFYLISFInAiDYBsKCJHMFwGpeYcC7JqI/
QPIdHiZIcbqahewHIhugkUTzdDApiJbQXzeOl0Jx7quvqYD9mRPgs7C+Np4ovIrd
8dAulLXCvLQnh6AYdnXCpVMSD6wVZiqC7yk7s3UgtSsABhOSYwK1BexHshiDCDu7
TGbF+EnhL/yRJ1XHQrv0U/c4oYRT2x6Q0AEzoHxRihaLJk3p2rtwzeNrfVQC38rn
wN35teRNjH2Lzb8YQcMPCqt8E1aed6SXdLSI3L+BBIoH1P9AUYlvoYcoSNrGmcbt
ocAeATJ3TKZfU8f5E5XLh6pbWW8/jnNCRiTz7qoePs4T50vEQYzkugfHpKXlRraP
N2+BXcvpF4OMFpJ9zmy1riGxDcQlA6y958pqF0DMrpl6iWU52uwkRwxrV36o3i9s
F+ZWDnEWBl8Hi20ow1ekZbaXOh9nc3tbwbBtwcJm6KPvZ5rpJNVsJXfn6hkziOML
MMd6TLPjmBkVbcLXLkPrvgjxPZpKgq0SYck24fxB5qGPnAdcdO6wWujxHCMKGx4H
BTzsv8DGw4ORWk2hRNsFuozG77pUO8cvBTDRZvhrkdGwJxHn2TDENJv9qaRqx3jq
U6DGVONd1kVN9x1Y/MpQCf7fUMFhM+2+GYuMORZVBVz34J7tckkC+R7OvPeWbMbZ
TbCXCB2QkE59fETqIKX96MQSvotHpuLJO0dA0VkmFP0RV6GTPa52AWR151gSa29m
kEFPq0P3Yis6a6mkan+yxc5/3Mn5Qrl2IHUPkG4/ydU3Bj8Rww9ewDnNYI3sru1W
U/Wv9IiD5QaaHyQT2iLa4oyHoK3ol/6RyvFX2ySOKKSD9NOo0VGC8yhVGNz/ajC1
VdJQBImwjqk4zl9SkdIJaR8flEV6oTHeFpKJUjKWYl0JRhW+ims8CuagBTx24zW4
ZiLsXJ54LKOfhCmeZ9HE43EX8jTSNXzZBxfJEKCRvFD3iIepxJBt2IIQH6+dGdKg
AUzqCxd3ppdIkZvFs1cY/LNdRXLSF5ZHuBKvRj1JTPkjzRd1qV7rXSMIVAi7Zly8
PkeGXZrPssV2o9deLUh9DnIfUj/TvAzXmbvrI2h43L0GHMGsv+VkygD3S16FTawB
i5L3sKmM5Lx0bq/ELdeu7ca5HrcEqzuZlBSA/fYGsX19zZP/3+pLMQMD6vgvr2Hv
ppgiC5aAdKoaj1fDvxARXKxM/em7yRyyheN+5YR427vS+rI271i6Y5+tf2fIzMme
B3D94dtPw9FpsYA3Bsf1Vnt+GDqskPkUot2tfDS/X4B+m8Ra1cIqIxUrTJ0S+GHx
ia7VVX4Wq61Vp4rG9g9W2XO76kJzo5n+3+s1v49h4zYYWSq/GlVau+kPrbex6ZiJ
LD7kUo9DOifnlFzWgZiJlMwB473tqdk9Hwb/VAqxQImewemiCXJJro1udFpYd0Za
+6ml8cU5Aax+xtwRkxfAbILQ+6Zp1qYle6K772lIwQ+zDIDlaKSBf1gUWsiKljhP
8TLzeLsTuSG84UR+LHcnfrjkDslTx+jiD6Lw1jF00oE5b1YBV/JVTlbYBoQI5fra
1pAIVc1KunHXATyYFnVXtmOaJes0NdYP19TuB/2zCHiNrhBjL6IdkMog8Oul4E7+
ZSIo6y76GvwHdXzXW3Jzft32vTz2uZVpeHCFvWYKV/xvUDB41R0ZFBjVAxJHtqny
Wa9nR0VDp4SfjGYJAno73lVsH1lY1oasCJGj/Z+dpJzlgw53Zwk5yWKee0V5+DDA
VO4eR4w0QecWUDKTUxlPGCD3EfHoSHOmVgLBLdnZQEdF7yDfixdOy7ubYraxI9np
xgYjjeM0Sy02zBT/Uqu3qhEcP7ObcNLZuRjZNCU0HCjU9q5HTFzftCXk6An4wO9K
Pi37SIJsyRdB86PTrcmKW5ehtZsfPrywaMayS7Bzkq7304f5CV7wag3kslHYNq55
PZVuf6msnFW5ekWGDUhrQc86UuXl8PVh5WVR7XYqoj/xuCpjpTRBEEVrmMTagSbM
KylERtpDGP8QD07UvTu5yAqeS8SY3qw5+jbJD0it7Wg2Cg3HOUD1Jouy+Q6kR/h6
P9wm92/oPUDEYsjwl+X3fbMcdnjj2VE8yoIhLex0gWfrgokjP5ZmASlkKmIkTakq
itKjmK+tKi1SCaJO9zNsCEjFd5yhjMD8MtgnKP56rlnn1KpGjCcqae5n/fY/fVqk
UIUD+/ZAkbxq4wC2PPJAY5kMhQGzleK2+dHy1lMG6ccfhUESDvSyTsShnD9LJgX0
jaZ4BXOui/L+dDipJ+sCidmcsDEvOzvgKoPFEzxL9hJaCNy2x0VIf6Gx4zF6zob9
2sqJ2I0/QG676gtru3qK56VSixWJxRku2t7xeTQsulZm/Rq8+RelQabH/gpV/ZeY
bNR63zKHxcHPPikXaybdXNU1lSuoqbqdNiVG44YN1JL4B6ZpGYLSb5dIel+Jusbq
BHuDBeSf28JSZ5jnnujW7fAnYBlMSmxYfh3oP8k0vEIn6aHUiHsYDzGbS3Awe53j
Z2XwV2KWosxFVRX07CcwzFvkO2SAHwHjCYeoVyWyrU09k9Jn2Wol7ZDCFs0nc8/4
n2gvTU/Z/UBTMCNk6zfDbM4AeT1Eh5Qwcf7s5wuWsLo4/4CAbz/lfi8FASw1UqrU
jhAyvkd1RfpROiMYIRR6IATKSEApI8QdgQrsKxkbTtr02Q9ctiQzcVKsnEz+V2Kw
Wtwm5sTNAa2U1fMZZXmoj6V8WbnpQSsrWeoP+rjspPIUsGwu6rmm/l+BDRQBfgUY
/A+yHfo76suFUyCZpDyxQIswl+ATInl6c3NGG2pmxJvMg9+bMpFFa/WrV5yP1m+e
5lewg6g1v5NQWeolHlcOduPW+m9wX+Ncvf6OLt8dIsE/esHoxp2DvwVkRzcKzk0B
bhB7tfIVvkrfnx6h5qEC7GpceRNNL14IV9UhbU8fGnPuzJhow2BVjY/7EJTG4WDh
l3jLoiR+PNYWZSFsMrn2Tsp2DJurj485tRVweQs2aXVFs6GZKdBsSoukz6z+EK47
6R+SqG035FB/gdQcGrbXf7ooOQ0aIlskzfwz8X1ttwPKdN2l0JhquRNXfOhmSF0q
icM6/byeZBF0FQ3Oji/U290ruRqEcKHAM9Y9T7BgzSCVJ0qH0KP1/xWAO3lWOOy9
m7/6pbVhOmjrHIo/9n0i1Ic72Ew6xAjBlr2PnlcqAHVtgqyqn20DR3frdo20p1WO
IZZQ3OvdUnDrpsr7caPClswdjYG2vIYRcUEEXA6d/lT6TTEolfcw2DpYooemkRmj
ZfYPOl0n6p40XILL7Uwm3LKACRodjwVlNkHg5qN4ocSwF4ZfE4DK8i+Jw3pX6JNE
AOFAiMKtabaWfdzpvYMOaQeAorCTQYPepY1K20Y5YeAv90m39rqU9S7QJ/5HMjK7
fxem25YDEEZfUjqg+y8ga297i9Z19/UihCgPbaq4wzl52W8ZVM6y2a010K524Lnr
QNuuejekfH8cenVH19j0A3BPfMGzz13u40tc2QB5nGTivKK4go6eMTbWSBxHZd6U
pQEzQnC32+Wc3TNjEfIsxvj58OpBylmAeFwLwAvKMz189cgarWwt+hQbhq0wb1o7
LuERAeML5eXvZ/2IRz9JIYpvBNOZcQvsn6TEF1Y8jwzum/4xUwa87GpSyw3nNsg2
aCL/hIlAn/Y5Hk2JI/mj779Yi9BfxTscog3fi8MDD+MhZA0CC8PSoi89f5DZzesm
AN1ejm8602OaUggZ7diuNzTZ0N3KoACMDpZqhMP+WHWsKJmhb+HTFky7XhsVnSax
/jj3EMT6OILYWE5aH5f1mP5Pd8jM4JdSCIFoJQZDzhWDnnDKu3R6QPAj7ql0LFO5
3Z2q5ZlweTRS7NRjlHpHw5PNvv9UgC0xKEped7dLIjnWb1xG9UfoOx/7XJEsn9BA
VIjuzqdZm9qJYaIUTki/V9hfi80XEQWHdPaS5pXicDzHPhS0pOB8l2mUVPqKTkth
Q9OL0rEejtfVOxOAuau7NNBUFmilyGVSKBdK0dg8AvdDf//WP9tYOeyiLhQfm9uU
Zri7u26hBhA2BniLAz2/dhmQM8yVnQKrxhdAZJjI0m6WMFSQzu2R6nKECk3R5DVh
w1wwu2K/m3WTozekl9z87yWb+cgxkAx+bRGA3entIzySedo00u/6rqb49jHuWlKn
vQlOW6qbCvUiEaxukU6mguxwePxRtXR8x7o2d5yXPIUr77VX58yrnvleLe573FFj
L8G75h9yZElSGdFOhtHJbg23/5e+8iiy015h8oDJSmYrqN0bkzDq8dXv/Gg/3ERV
wB0mjCzLLwutpC1fCNAS87mlIJQDssXe/0t87ijBR6yV+pStUjptY4Lhf/GGNBW1
xRj15N9pOgPttPFsJaBvFJPp93LBd65HAIMB7bWGMtRRFv3nBT5bgJCUBz1xWHte
Pu5fyqJOvFXxShRF+Vhoy6Q4lvFC9WwSCE3GTl1HGGTKRXXa8yF++Dq2EL98oSWA
uiUnkQZ60Uuj0Or8DXUPyIoS/RqJ7e0IgjkHZpqipaNpX6rm2LEIha+bPGUhgRBs
hMTblTNtDzhTy9HuaRKvK/PJy0fL00x8cMQvmujrwTvPu3Ofm+cdNLGfAkNuyLk6
YwsybgfiGlUjFgG+2S1LuvqkGGZhoL1lj9Mafxx/s5Xt+qY7eABYfe789wOFc6qg
auKIXanI+H6yLluKw7TmIbqMxixRF8SWXm79/fNiuKd7RdCtQNDQzZDggk2hrnOP
l3lb5oW28u+/GffvUQJs2gAkLM88WJKX/jWDGWsCKUHemwLj6EyalXipEJFAhPAp
/15lKGMFwtpIPf1JSRl+GIWbcVasFExuUny5RKzs5AUw/UVmABgqGwewoZ4xNoz7
kM6MB973pBBIa7P+D5cWhsHHNmxfc4VT80/u69qftSJc13gieZEaLTMduQzp50Jh
PL+Ok5zfP1LTsbn40OpzCABFZSUA7otwJ0/28SsVg2WNJ1YkVMFYM3FWFq2megvJ
5V20ppt/uZyRQq6S470yMX8Ep93qbgoW/vA60LPs00wWdVZsApnhjYrUgNeewdlz
lN+W4pJHRGLFFR3QRarp+cm8ByPJLE5WuKoNBnUkwN3cbBq0pP7xXhNDe/2xAZvE
JOJM6k2ids0veqNlLruo/3ftNmqQNCI82e708094lc6m+CTCz59wGEHEJLAsDBWd
/sP3WX1FEuF9oezb4D3iyLJKYOyfEAeCwoBuSlQq1dhVcZLHN3JumK0IfbkD5zRY
R0ebBp/Xcp1lNpEEBk/nH2paG+S+TGwIj2NJFiUKLx0HAu0A2VIBALAJ60y53CDa
wVW9Cy2TtV4LGHM9H/xR9EtfCY2XPZYy/jbJz1LtZXdWErfQtqATKI1yXajXxjAc
8HGNO86ksosIb7wq4c+6h9V9KGwaEG9drGIF1EoXkAX9Kk6okg8hBvIHcIUT04sk
lDanltz7vBK/l+zs50dg87IfM4Ru+yrToT0XTXa8EisXuwuxQNbXhB9DSyNPstk9
DlE2CvJYajg1HLZxpC01+Qw73OjeMXPrNLu3/WPXcMuL02Qmx2ZPGtG1cuILF5o7
FPTCln4dqj37rSB90aYOUk5RWrdnXAH0ProU1L9OYJgo+ZksGhAUlt9aUjTkffXz
7w4yA+LGXb9px5a4JWX8C9pPWIKUc1qExHiO3DypGKx9MwgF6TAMpW64OlhF6VYK
Zs5Zf3hmJPIqWlKynvjsqazRyB/o6aPoQHeHpCQTgYydm3z+UMonshlHCig6f7yn
OtjTjdTHQsqsFjQfYIrsiVbaejAvavMqi8YhO8SwiKl2CIpzav/9YPKOzBOGLl5L
wSytVbe1B8GYS3DZk0miOYA/maIx8oI/1nX+6vSDDsmeoX1go0riIncfE+CYeCoX
7kNJ7PVEXAmAjUcIDYH7ROjf3o3xcc+ZpB6aI2DSN4rvggaGPVSB6xIuLXzVThUy
QXdAIEnJDzmCxkLU9HFn05m29dkWDsueRakN+BganYr0sNOTUthNL5Z4wExwZcdZ
s/xzl7azpZREioBWJeNQoqDUTizcBwmgYnUx8SwnvIApu2WB+9TB3YHWbDS22wIM
aNfkrOLz+LNqxnykQjWl75sT6XvnOFy9lotlxn8LsvfvxihiTBNT47KYNQabndNf
pRFhJc1OaHx2z3sDBOHpM7RBUAtTdBzO+4c/yYUGx8ZfOyuHVmtpc4ubfDwMqQrD
38SQl6lxDg45mLVFSqo5hdu4r3Ii0xqdf7LIXcfCdxR+1jKq42ipuJ8mi8OH6hkF
9D6fkmjOkFSrEZU71iqJyR40BGAPqiFw0rD+cgeiCWH+4xK+EYRkA2LxGu0rvGFV
YmdtF9VMmSAf+Vnz0Ml6XO668JGFNsM5oNevNBOMQ5mnd/W/5Fj6mwx8JeAkkGUH
wJtGnfFRZTOOQ/z3lE+oHgcWmDYlxetDFz2YafAYdDC3/tbqPIC3DUU+dbL38WEu
kJYMGQAI7JAzQwpOeyx1DnpCB0QXgwk95XnUhLf59MRLrxbLbbpam+EI+wKIL7eE
MQ8BQzPFWBnnLMCbxHB5QvhVv/06aUMcjZ+za/1Zulip6aVyPt/s+WcRAD80H9j9
X5vVGJPRV3ZgNQBSvq5GthtXmD+RB6Byo9Y2FVl6sFqXn2AZ/H4CKuz5Zr8B3XNp
GZqBZDfZQc3zMulT/fYwUWZqG/24a4CaJ/ll48Vf0070Nh+zHTg7YpTZDi6MPWDP
SBN4AszkSkaMBuEZI6NKkQ2yi7So2mpRKhzyK/zg7PpCwv/zoHlJZh/EXrOVB1zm
GOAXSexcrhScSzd5layptS0AsVdktwAMjJsezUbzmeYdGWGB6ukAFAPumc62sXfC
Cx3rSrdmSo7ZZiWyWYnga1aWMTPikkFu5iBnVUv2in8T6keLm1nr24tFWwK+7VbD
r3KxUOPW/VuQgTnl6E28AFbWWtk3dPQ1p/9vEGWZy9OLH/WQQqGTmjXyEaj0tB9T
x1paAYFsEpuOMSwZTOH26p3+OazhKr4igcFyO7MOBxX8ZvjZpemSnJnZtao7Yvau
rKJccosN4/RdfWkXoLkO9B3be1shct7MkRjbWErGvP3tahl2jrMJ2RhUOltx4XCM
Ree8y+JyE5rsBMhtlcG0IgtWXigA6y1MtbQgbiOSAhLXlwWmEDbjpV+y7oBYgdpb
NyPyxBHUBYRuOVqfjRrHKGFn1DunNT4NIvfHgWw1RdObAHysDQNore57w/0ycw8r
yo8Fy4KSWM+t/l8M1EhxotnS8oUgCau8yTSosJlTh22GcSRPUvlGIpdAi6f9ijIS
KFuW8STfzyaLf9LCagWD7nr4bqlkX95H5lyDuWdwrzVYoRutMXjITraWQOQO1mKV
VQfDImTnMQsGLhCGr4RKblxPWkWpwQ5RsHfQarj/CZaRCDLem5poMpqzzZIO+xky
m9ts0oluLAyACM9BdHtzMk6uYrHdWg3Xwh0CedjAtIFMBnwXmKMPgxvdI1HMTFPg
jtvegA4M6KfE04NE+OGE3jTkF8RWdepjiURAUFMDKn4OHvZBuBFcHPEQStl1BiTN
TrcQ6XjV9N7mRJ3gN5uNU2R3gGKSkTd5G9yqXbDg+ZN0Y6xy8OoyHbZO59ip3Tlm
iw1mF47WkijMu2FHBlqXi9VYzWr22gBAoWcEhi3Rd8P8m/2NbHUuyigufZdzM7QW
x4VLtd6WZz/S3mPfOpRstRSSkZ7upX6NB9tlmqdPnr84N77Eza0kWPaqT7BDoy2r
uQdSP+A0KaHlDXZ70iZskOrjWOjJeQKd7RznwwYjvsqefKBCAZuT0rCuI2ExXlih
efJamOG/76MlypII0/8psYsTC65xO3gRdpONXLMr7tJG2vs1RcDP26nrd4AskSjC
i27Hgv0fQtfGl52cWOYDV6I25aHB+vsmK1rMDdHTKCHfxoxeIQ0XLW5JdGbNZsfr
jV7i6k3Moyv316nDjsIErKfzDeaVCL7Ntqr8PnpJNCbeCpAUJWU7shgkPTS3UvQB
tRsVwOpKu6Sd6UrHNRM1957KbvtAofezIrFT2kfQ5+Qk4UdQaHbKfE/iK8Jiw5a7
CKGPueGnfFPwgYgOIsYsZpUM57t5B11qdaVwXu/4JaDXW8VaRXZtyy26lYTXIEsi
KlXmQO07CnbfcF0GOoGP3GCTv9JotF5qXLNkzJri3wfdRiuccHCt9thvcCHmR3V6
HL2TSds8qwSAraqv5SJiIx9OIvqx6ncGjKylwViQHuifaKyRH4PDfq2DlLSog7RA
EnRv9s2Thz2fQu4qkT7GCgDht70FOP688rVJYKsJ1qCy8okQhb65R8sQiECRzSYC
u35nGn4rGPw4ORsWhLBJw6uqyOTVwOXZxTfwqZl1w9qTxupFkrcuqNpGllZh/V67
Pmrl7eZQcHxm/eivkUo4MrVQOnuV2nYVK/9PBJg+xAHMzlKIYjBYD0RygPJDvhlU
lqBzKB1XeGYTFNXFTqxRC48dTXwm+tu1c4pO8nQK9NgIyQkbRUc5W5h+EnObjYY3
Ri19BNEloAI8NcT44XQuxoUwRpDn4gEoCwPDHRwIC1CRL89qSnQmDFBeRel1bZrv
0VRUXUH14pVHY3k6qF5q3PPeVqK70TeTG1UhBdD0xTFsTwdvQzxctu+Cmm2EONMe
PKruqZLDjH5cMKTtqWa0MpaDpSMS49pPLnUbOjKJyDSkmsX2QQneTej//2TDVA8i
q3QV1jWY/N+nubNUNIZucbHZ3pxWxmz2UDBkyuYC9viMuMN5LuYErk8+kCzepUxH
6u1peLxn4PKvoRiY3/Yc7iqkdnCTp+x542NQEfpqeTEKG/sc1t9YzkIh9051Xnhj
Fu94J3cE5Rwz8p5Vm2/HnGBlQoepF37taQOVYKIo0F1deuQ2dSIj2PTgfgrEfDjI
bRTrxXQl+YAxd8mPT+Q3IFEfCE+2UgB8hhop01NtEiSclJ3ofMPNFCt2LEg5BCfN
wa2CpwzKxxDW//OhFSygS7yVWKYnmuQ9aCvqXoJzhv1H1MWW2Dxw1iXOIk4Qgwes
R4n4VRs4fIjAn2WGwglitlUmVVrdKx2dG8IRXsoNpybjXM1xg0+aNGy6CQKYCsoc
cNO9vVTzOfFph6JLQNoCnFn+Ous/emws4Ot25bf/wdpGEwOYMrQdODrlnYxQRgL2
3U8qo1X3HR69I/EuYfJ9Bzg3fZ6y2GqmboPBzNv2xBj3UHFcBXqJfbg3PzsyxNIm
+uV0M7t6AGq0EfCZ7aJPXhn5lVYqtK7WRN0S4XbFS9ZZ42scfAMq3nxcaX7fdVxQ
o4cYamVYOtokQsiHAOAkCvWJedqgJYMPF6JqNZE0jkFn9ubggWOQDNk8silK4bPB
cajM4Jxgnj7sGmogP3KXGUSoJ3OAdLn8BMPBgCAx0/Wgl5/TUZYPjzNLsStYDGzH
JuYF+PMjiZS4qWgiQoERMwfETjH6EY0m5pnw+G94rZxgyvnMf+Jrl1R3zIJ8u1eo
bevWyhhC1JAdJKYElxvZ8Kkj+4XYu69YLYMcFDE2ro3TjJOxXJco6n0Z+yt/pk24
hMgPocPqvoZ5O3EpnFRJWGq26L7hI+NBZzDgvAd3DBXsd3OCP44Iy8KcYqRBUOmB
4kI7zdQzVwJi3x4haXYukU9WpQOfVJFVqPgTmw5OjEg9+RjPe3DA/3Hrb0Oq30fV
l0GrYygxU2MwosJ14+dakR7OKUXIk6Zpfjv0bq8d/vk+Et1Q0lo3wu/UegUmAj49
xNsIoXpHTT7v52o9pK/6bXtg0iaG4Ws924CBezA5RLKceXVHbxardWO5yTsEXb9m
q7Xa6o6vWMLsoyTNtBBC2nARW4kdhXEMrgAWSXamnw1+827PCgKHWYLIJxmwYceG
r6QgcttsWjbqH5j3Wl449BiEIc8mDsY0s6P73tQ98iYZgSDmdT+pmTXoZKbc6Wfe
BvVER+2jXCscn99F2E8+b6Ad/onEe0trvXmigOITkmU33CYtiyZfZ+s00QS/sRYJ
pH+mghU0zO63Y6j+7CehdvmJS0ju2kImYMLsTw303sQYLXqE6Bu3uiKWDfAqU6Q9
1O44KRfXqCBtNGfCAcIO5yMQ0jgcN6Xl3yp1KjadnvdWpBzrBw45jw+6kBZoGNbX
NP7hsIlkFWe44vh9on/E1TyjGqYUtjpZwkWJ1pwGgoplFJ1+0jpaJEOXb/++PlFz
4Qxl2iZrR9zIzeFhHZNlCV3H6UEJE/br+QlTPNEZHci/MGS9kfdwEpDXqe3kUTHp
GPO5QpTeCtHsFftUMVddqyHXNURpItyJUT8tk+j5rX3p2F0upsXPRs6R4rSi3v3z
UXie61AXjkfSi/qvlbxrKbvzXElZ/RgSASyagZMmhIXnw526WzOjZ5dMGaUakpAz
hnNYJCXvJ/xtXlqgR7viBZyBkwl3rABiLUxIMUsNshc7unGy7ROHd82XPR7E02qL
OcHs4e2LwpjUqX8fd6cFoNs6FTiwqBQbs0TwRv9ebS7c+RmMsr/G+eJoinFFIQ9/
7aqKATjQ5i1E1NmvnWmFzzlIYTRshBM2U9+k3j102Hmy0WNaUSs9eroZWHYztzMx
ohYu0b/t+8jn3pvTuTPbgbEwMW9C1DhWud6A6zA3XO8DAT/S9o0GL9NBInD/wnR4
xcVkhE1FVy/EUFu7dfvkpjo5MoMACGLh41hrfGZP9Ezrv6SiTtSBIGb4qfrROaBE
geVfFfqoCeRIeedwXk7Kw69A3BkgS+L5LpGIq1G7BcQCpnAXLEyssLqPH1qDW8Xo
10PAECI1PtT2TD9wxa2EVSfgGBodp4fBPp2ODhPpQ5wcMBCT3s4nIJHAt+UiNf7j
3915fc+kgCimSVUnc38WompyKlqjXUF0K+l87jOwucbUsIYHczVri9gdZ7QyIhOU
LA8BezdYTJXNlpQxJPWtmF2GBs2BJUUmihPxLg/HBwWkqIJowzNUy8QZI1fHCDc6
6WKkLBjuiOlR3Jq9teSfreyDnEwA9vcWR0fD85x3daQnCz/lM/62+nsty8RLPtdg
6WcLxwlWJ6H89bOrGHtQvTnTLU7DWY5JqseqGEEHph8ptH1a5Qyk43JtfHeVV+R1
XtdT1wFEEzpPurulrHIdURSBlFXBOcitJWC+SkHLfp1CFdamSeeCP44VH1KdYy48
arwgxcoEv1YL5LUX2c8GGnUq4FdQg7KAmfUvmLVH4OsIoWT266qtkqcKX8YeNLO6
tyApra3E2jaWqIGJXf4bn5KkQ6QfapnwKCNPiVboEDdP79S6U6fCjJ612o5ALBJ/
KDbcWi9JFSprg2SAzjrA8C6Sf1R3zTRtKSk567ts3VfGUhM9W6eQR1BJDhvDEag2
FFaGbn2s0i+P8DypZZDGObcJL02qHdIiyERmoSCaqSck5x4+8BUH+eaWlIKHtPkQ
4dpqPH08sFAKiH/2zr0iddz9k7mBsa1khvT24Pl4EbYrcTXSAlK9SZ8tz8ZBghGV
nKG8Ehz08fu9a4EcqwLM3MGzeHlvr9BFY+lVlNNUWtcwGvP5VETp8Zbs7s11rF0v
gPVo1o8pWFFGjfD77nLBxBPYsIqeomIsR7Dl3Rg22qUIQKFfG0SU9FwXiIFfHUjg
Pk/nOAVKUFVyIyqXs8VyfHzH1Ednr9qo8QaKS/KpJ4ayjnBCiisT/NVIa6aXqGSI
hNvwQgt6McUjI/XdpLeiV8F5mo/GFY8VHR1GAGXJ0BzP+BB+F9SVzftzbdgNqDZN
LpPI8eAyctd05VFMZVUahHj5zbO0+AeG7nBkKiNBz+wpTVX1zQmIxfQVSAlC1l9C
CI9PUiTtkNZcsrhGaFNDGkRuUk39wdHyg/FLCKJTjaxE5w/1qSwgVZCrpMFIDtp6
WWFT3tI6ekoju0xmeReQdE/bT83DCjeSXcDOkEGwImvsKM1r3EbfAzPPCmfcwUUT
TtQnkskJf2GYGsM28g6rEi3FOy40oMu2QVXUJqmJy5AfWOy0nhwATvgY4In9ERAr
MHTqEiCA0DA1i8F33mvM9+vctLzprjCGTy4cqeukAIwsKt+2RgbYo9SgGmDcwcxM
IdI1A/hhinoGVzo0z+2lZPrqTmLoo8dEyioWcdEdxdzaAlVqFCbgPlfBfpVVlXMD
OaPUcXj3Of/8BV4GJaOSATBVJa1TP3z6e1Krors8tU5EL7lLkFhD9ZX94ly3jLeA
vVw9DAzWo7JxLCGxDlXloDQ/URH99Yfdc6aaQyv4CK8ahy7U7F0S/XNPtQUET5Il
LvUj2gfnb722oW35qpNUlEj4zlIpHJ/rylC4E+Vs1SsXnoDt2hPV5QLq/3zyp6lZ
rI5dibcd6CobAx27ksWY0aUEV1F7A1yyTAPftTOmcTm+2xYcJoky48AxocEkepjB
0qT2jiipWXdnpJslDWB0OCszv/qdq0wj6kyXVjDSqh8G5uUArM/k+F49vfd/Ez47
GtZv6InJuU4stBCEhAE9c/XXGx2p5j0wCkSw6aFodWgQE17mL9Jk9iJ3LQAiYK+m
Sldv20AMOdK0q9xzdRj74HWOJ78S/sL6DlKK+mRuFbrnVtHe244B7GxkbaIre2LP
usK1GEK+itV09BR1jB2L6BCZXFbnZU7kfWx4AMoSj7jO5jKbvknBPRT523rfs4O/
MonQV8tc6BVfatE/m4zWm15+KszXHqo0iQxCfpqdjp6ezX5sMT4lvDbdfWS8IMBM
lD/vOZer9wSR85K4C0/7Dp+ZNf2zFukEmaJqm9DJTVbRb1wG9udGwPXJnsZPitEX
6tF1QDZyBnVTHEnDRCN2H7GeaND1b0ub4urkGO05nN40o+7UFVWWISVFRBYX9Kjf
6C8Y5t9EVRwZFhBhPMZ9vS8VF5FJG7Wq77ToD9ysxf/w9TeHq+lZ6j0MtngyrQee
05AiqHDnc8NymucOIUUC9MO18OlqXLNu2+EpnzSg7zJXLgd3JrPIN2pIVFTCFFFl
4tE2new8o74daG9m3OhfGdQpfhKY6st9NjkiTV5UV4nFXK4v5Cl+UslTfMA7EkJ5
Ap2aFUISzVKm1XwwN2snwPxKCEuv8jQga+TCgPPZzwv8M/APg6Oz/kT0Kwowj7OE
M7MenPElbSCWh3Heu9VjiE3pBr+V13rmYcWTtyKxSzvPQ34Vvy5f+gY7TrCjEFZ+
InA3A4x1HunbZXygW7YemPNZGh7VqLX0O6adfY7d4n+GXcIryg0koQ2uATDD1bpt
83Y9qzLjEAVjvWktr1ciWZSRFq41tIeaaY9O3dtHSLzjZ5wNW7JES0bPdb3qralv
N7rIgqg3QnQKqwuoHzUaCOlhwhBjIcp7GGNWBygeCt3emj46ZyevgXEQ0REczI92
z5YtMhpdz1OxxIWTXLZWIYn4cEKRFdJcEMLaY9agjjmaBU3L/atbIqkTDDKDimt4
yWfKuwNxhBh5iO5BQgfvpIyOEqIO6tJbH55vZCDnnQAZAbff6D2OLafaiOcQZ63+
VnwhKS41dTn1sswm/b78R5chA2qCyWabx919BonrhHmQX7rs2lIuktUC7rGX7a0w
iyfkEIesQ1/axQ0t0VV5XnUuNAxT92JNBNN4Pr6nFy0hCCcfpv+5XRQI0HyvedMX
NhNAvxhzlgo8yWSvjkZT8qQzHIaJYXKi1j/CDaiAayHM+MShjyGflts+AruB50oo
20mzys7fMVmg+xNf89bytR3+V7IHX57j0AIogMkAX2TQtwwvuL5ugMoy2Hc+J16k
R7Ihep5KGhXjwbhDGs5IQSwb+mZZzjMZ5tPB2UXi7yHHm96v49VsXQMr6G3xe5Yi
EcOlmOK7RHBKlUTo1xhl6nTCPBIWjb1QWqbFzQDWEDDY/1+/OX6UKcz8QzBzf+FA
0sXcIfRTcadS0LyYa08oTo8f8hZukVAdpCa2zPlDigkf5gKsac3bWgWTd3t5M98e
oFEDYBD3USBM1hHvRityw7EyvMkP3mr3EIN4wp5ggNj7RsiGoofhskkrIGvKFKKE
RfDw8b8pDT5EgjEEeuFfOjZTE3pUSfXRxjZaUwDGvQqGyxI+7Ke8LucLBU+FR1zg
Qir14BYgkO/Jx/0zy6DUy2EaoS8Z6hkB+1iAC2zPJBdXcA6S1r0H9J5p9zAFYAuk
T4f8e8ycN++lPVR9w43Ko0oUfc9RnebGfsNR8XRt8o/cDKdjVHobnpU/Xk+blfRl
VJjW/sn0gawMd7lhk/S04rfVuORefbaZB83pSr/tnlZviDgvg6/cF2IjKJAYfYnH
nyS9AWRnSG4wf/SP/tllQf+yXWwRGFthtnAtTIaXZRLMxFptsAdKRm8STPxnsGyq
DnGpV0dboU5xIEdC/pgTIANULh8j5/uN6hVmuOpkHNrXDpKraAoo6Mjq0yurb9Mf
o8GYMfue/2IJVdsGkYlrHNqq1Qm5T3F3ZgRXIV+qCEdxFATcFMlkOaSmLYj85+ya
9QJwQYH6Rd0EuiU7x4pfpW1EsPlrV//XbVmaH7vxmyJW3P2Z9MEJYOXfUSV3g8au
SM7PGg04iG39UQY4v+5vksiNHEGl5Q/NPjV+O1kysJomfP6GxmaaCN+2RZLZ/dNa
eSEB+Rkkrl0MUFU5ADYBn53fbQDs3WIwBRY9l66glHpvX5KiO3f88aoOD9n/eo4b
GlbUj2JE4365DbLhNdmG7gzgOsOIK42/CkE/vNjggHVQtq8kptS+WJfBsKWcQIw3
rKb46BD22BMQ9/XEFqfgBJ9tD+zenYQEwJVzhJ6v8BPbu/G0bRZSFhpbntRS/5qz
QtBoOUbF6f9PQjTC/vKWWYR8YWzy9eoxVnVSumdqtotSh+63wYb1ZHgNO2M0Zwel
NPnQirRSNXJ73U9rwT1AIe1I7bdJfZ9OGxK0Bf1BtLTtPqNN/kWjDtWnrhmtOSUS
27vFg6sKOVuSN5RYevIJDE+SkC9RVRe+qXcOfzpgvrW3Sg/vMVR9ZzlHP2lx0nGw
ygUn9erBGYgi9r6Kp4KRZdLtdQj1eEfEzdvuaxCWb3JslYq6tRJMHVM997cBHA81
utcBtyUdUbT3zncpmSn06D2nUlyersmflGYLt3wbc4lKlKP2nSmJuzk+JD6Ca3Gb
m4HOWOp7KvSzlH97jlxfq61DfFD3gR4HaEKUSU4oGM09NqFcpr+Nc/kMwxOHn1qL
1lEm1wmAvA/1AHoiRRyYL8qAScKo5XnqcOWvpg2yiNSSbyKVUV0iZQxKEQSRG3Qz
djAMmWTD1PF5TmtyR6+eGPyKAYk+QXDbBJcfZKYTi08oqI2SZXmzrDhZIRbwy5Sr
4zIvSDRt7Qb46gT4D0+gQMcx3YzuzTeZIuRMPYXYbiCMohPZD17/mphAGkGSaxLE
N/0TH6Iq+jood4kl3/oh1tDCFajvn89CQ+uY84J46Qisv643KyaaFRA2DRUtwxTz
+o0oLY/uiJRq7DSGGY850bEVYNsXnIex0jyuO3Y3qfiS4QROArlcDkz3vGiFfxU9
tbiMbiVgCDzfKFGStJf2QSVsPXU0buadWIF3NmgNS96w/tSaomhzJtzbFaO3VvCj
eY6W6JEHt8mwHNLNtOdLUobn123mldmHJsqAvA9NMNLtNWstDXiIca5xzFm1o25e
SJnsO5KGQowwGQo+N9tgiuEnFrF7kZwKsI1X18uWLvcbQ3cDxYDUdTYaz0gnOQpF
2yaG4VwiSz75XM5QzURs50RhR7v1UrfIZCJ+KSbgJh/IgF7o9+RK0ltRu4zlBv1r
J4/zQiCMhT8S42iVHKSXJlu4/Xy/fs+AF+HmQ3a0q1WpVJlWn3ZL4bHxLyw0C/aW
Cebd9RxX/w9GRrXOZsAygxbRS+iXHh95iSNZCdoiT0TzMCwX7RO4MsRE3ETjHqvW
kfWM1pkX0X4SpGK7i9DXjrcLCUWsFo4CEtE1R8oWVtsjOskJ5k+tVjEB0wgifA36
+eUpksTcVCsF71mCzSNS/J/7FWo0eiYRHtoaifzLmn1Zsh5AOon8/pLQUS4hEe60
ARkxDUk2WANYDu7lKmOW2XyLTa2uAcR0fZ6HIK6wJA4u8/lp6kwKb4BYAdeeoKiW
h1gOOOeQRlTC6ZqGLksaqXRlFh4x14YydY+R2b+v6MnQtKVSHkfA6D0zPD9VaVM4
TgKAL9Sunma3ha89mn93sEtzFOgXZbB2elahX6iW9Xsid51snknivbqA/wcQzp+e
88B+35fvq+3N83thuXe64tf3yHssBZ0mQumFCEXH9R1dlzxW6kFycR7Onh+TXGSn
P/mwFQzSVQiGsUBFCWh1MkAy3uBaxsM9IkZ69luCWA1nB6b/aODE98nR+2jkNpUN
7QSb9yf0v8Hx51M1TYEuNIHoQfDVNv0pfABjp/CY0g56epgB8SNT71nlpStLr9Jn
/ru5j0sU2pOzhIi+bWYvIhJDmy6kSZ9j9VFlnd9v/Rgu79weXuCeaqvfRB+GN1rG
kaOBaMo+cstNXWLke4y2agHpsSSwUO2tOPVJOyZjV6QVjVPVjwPpxVFltnDGlOPc
R8ovZ0tF6YxsGvsQn0rUoVNln985sGB1NjoU44rBRBh67/RLJNu0yXo1er+wIA3N
0EI8GOrL7zbjk+30JNLgX224o377/MQRUFYbgmevhi3QYVxJMZEBOcWO5LT4+HLK
F6abxmtrWyhOtzj85JxfBxYUrYeOoVYtQ4o+Ti9BOgs/MWNmNg9/ru/caItvVXSe
DkNABQMKfHscNNZxaj1Y3rxtGY6lfLPnnmYhb16yH9qcMIujliPV6RtdZkI0NmdL
ePYqOIw+iFeaw2EK0bVjUoTbkt+rEwjDRpyRgzCBvx0tJhki77dUUlSIbqI8kcSj
IvWwrJRVjTIEMsZyGMgh1k1JC+hKQiMli8aXlD1BDxTJOC3pKvIVcOOwSXieelXz
hZSqvw69BmBVpsdsjXyQl7TDFS9Gd1kO4twIwX/TsxJ2k8W5+of6Y0jR2TpDGlwl
2FnE7za7VC8lQdlkM3d1CuKIe9fQMErG/uJHDH7lUa8/c6FvXDdoKqm+ykbmkKyh
ILDVqbktaJX5UFgRpiJP3Tm3sk9wZJCjtbg5LYLqItK6racInfYFAYr+pREanCFg
5LxjdBQ0l3Io5VDdAaNZBlktsiUkdWvQ3Io7fqkI86/RY/iztl9zrQgQEpQ3ix5n
WBn0Wip2b6AkiM6elu5eCWiOGaAohy5l73ybuv0MC9+2oAYJKOgP6mpq41Ld2KsP
boJsmPGuDnEdiwwVt/sobUK5/Nl5Ai4HmP3UC4TUrdJNywWpo4DF0qgwbb7UF4wu
xVy/RNgse3QCzfF9XXkLEQGs+Q8vD0x3zajxdMHwOgWy93FEkraqPNZITSn+SnBC
pVxqz+n13I5wPB8eh0Ab+LYrZIL23OYrjEcjEryPqjd2JXMV/gion3r6LpVamt7N
p+WjGdy7Cr0NxzqXxhfrwUqX38iSM5pMlZhem8BwqxcOw/pIcNO6ygE1gWQjF9Gf
W4L5+55W2SfON/nhxS29yhQ2Sh8HcJ1v5HglDNH6PxASY/cGo43E6rfGWAFbcMRf
FqqBEx5ohXDzpcNhA2zMOh3VFnticDXq5iH74OxBxqhEYFXk4VtrX7W4LCod4fAb
GJgNO70XKadEJcAnbW6pgVN5UBiMYRF6u+2aj9SsPJLCFI3gsy4HV3BTqkYKEl5h
a3APdFobxgBKdemf9TQf7EB1c3EMNqlKuYFoQin+I0rYHMZLzVUGLsF7ddb3ghx2
UM4pUIME6uh1bemMdp+GlteLV9TOQFbMugBRGbc2KZka78LB/TTVjbVhWjlWA4rj
2YySHjs9PEWogg4zt6V4Jeew92LO5DefWuUXp5I67VqG4W8Pi0nYeSk/KCO8AVvd
WyORusDuySihc4EZIEadTvruSxhEhtZunhdDhjc0462aWzX3L4KYVHAoMwsNnPrG
h6n3F2XM7XBdq/ip2XDjIL9ACFrnUltRB8RMRIKeQEXc9CC5VFb7qUTSMewyu1QE
aacx5pijdGOAHIzr2KOaIpGP6xxRRqWcm32DKpeqsVevAJCG5eNaTtDDwPzyxYx/
JAJOfxZe4aWlCRpZ/hbadgDwP9Qwgo+9LymgWX01sObQ9828yLKTxo9WNCHL52el
dd7FqkWcteXSJIXDqZYo9DCV0CjOE5P/QDezihi/nVHXVXaGEbU3RRjfEz3YHE2X
LZNCXXab3CWMOCRTdQOByJNT+IKTGl+nrgMZcRcG+zuLz0ZTEnvyE3qQCyKnuvpg
dvtA4+0RVkr8UaIfGvOB5WuS+6vbYjk0Zw5r1sEpI8y6p4KB2EwMhe4+c580NgMD
o++HgHxZQNxmzXP2bfk9JkzTMVG999TpIELF7x3JM74nzc9zTQ1xo9hQBS3ptc41
ROJiOCxB8BulllBm+4sbMNvpXdaYfx30NN/gIIYDZn63OeISQUnOw51i1l58sy2p
wPw4J6lqndaSoZjV8H3Hg5vEikzR0H88/stE7N0+8veImL48T/9eOSa0AhPRyaoE
iRwm/6CO71Qt2mtfRitHCB3JGPOZlum8HgtgMqFcPaGPU0HtQA6wssoYnspHDvf4
+WJj7hB3oxYcjFXK3ONxVvgOe9zzbjFHfTSM8nERl3oXi6B+hTMg46AAjT5XEg8e
QSwj61kiPPq04fksjOkuPyR9JTGBhf8yZkibUbVX0Ii3SZQNUEyDJtTEfID/4y+f
x5XqW1hw8I1I9olxq80NFvwh7o2EofS2LeRJtRajZ/A+dDZ4MtQFjjifPEiTfoWU
F/36jLVLQsFsXvrcxrPn+kbCQdgm326UzgoJrkNJVV7To1MnvhnsFVD5lyfYNWWb
w1xqCWUgh1SqAhpO8MJ3qgfkH+2aTZeqdsFaLHyOETMdMLryItgMSfi0oyt4NLxa
6hag1qZnWXv9APG9rHQVoYm0gUG/y1TRmShS+oz78dWMyqyOb+uY3MKq9A22WcTS
9WRN5tcGf4Rm6XmCdfTl9FC9wDdaMtnx5ia726pONieLE8RvBFrxTdMRDDdNRLS0
GmvVr75Oe9O00LaRUJaLiro+r9Ys4w7/Cfq4mQgwgkKoYoGglgaNL5+NF/Fz5Mhg
7HlRRcIdhnyEwHvuoKz2eMdrDK+V+ulrXWOGGd0TW9ppmgyFPcAcq0r3n/C/SSRP
ZlSX+mGocJ5zAUFnMG276mk3YFGNabzwJ29LQj2Y7n4rZPB/8LPnEJB3ZK0e7S9X
VCXQcq7rqH8mLqAT4KOmJuVEw83xc4stOfbUrPi5ZdxZfbDDkELDQgg6LujJhyGO
3KCO/I1zHVo8bB+uAnM9lrS1SSEKQfAyBcdGbrvCtrurNICqQJbZC0hYXNBvCX/8
Ha8s2W67kPJTYdsPDWhtAjuMGZJUsCoPOf6fY3iBQ4iWoak/3q2zWGZV59zR6aPE
VMnlVL52WYlXnWPcT7LAXJMJVo6wTAf4xuxBSy9yvIPCfoRowh0m5nLp5kwDz+EA
nBm158NYruivlWbDv4yYNlM4k7ii/8elucUhKy14T2fNfVHBsPD2vbRrc6YIhfjV
skCcrSL3B9i8bK8yC/bl7hwEM7MEUFduOh30xyrLiJXTLqRoP5yXTUfnCyL4LYF+
k9Mrzhzkdfkbny6izGg2/+hGYmRqDY8ierMOLtrYwhoMmyIBfMUrPJHcaQ1fnMlG
pPCKtPMyOALYGN9dl9ldMPsrREwdUC45y37kSGICOxIzibd2oe19hqiIE+SfG/0b
GTJOTPeDchjS7oI11/bIZ/v68seGBPk8dnLIiShp+F2opbmjk6fjCIgo+JbRoUZz
tgJJr2jlqUu+ypBD9CCbZ87PkuJobVPMN4ZZVNFNAno+S8jvQX+QghBDY2rTuy8x
Rb87z8BGQCItkaCAbchU+UvnQwGbbFpk7gnVcirQvlRelraV8lB9F6OeNfFmaT3G
7s6SluKj1ohV2CGeidekOVAPqlgUOEeTP/zSR0F0QXuTRtoHU4uF4pkialWpxeVL
rgZryqNF3R+5RAZPHegqkORwJZk/5J/Odknrsnr531DVpx+QMO/GK//0cWxzej6p
HvUxghCZxc31iGzxCJFTRNzJn20emHNy9QeaVoBXoGdLYG4OHbDgbDe+OrpYw9p+
Af1+iIQNcpV1oiTEdnNPoQ2XfUa2hIFwd+nxKjimz9eDrojegQuNEtsvDNTj609P
OTX1x3ADFNJ+ys3fBFLS1+63JhvQzaN8Ih7D/PFvnDiy0Lr9IDsADxf2bxcZo+Ki
5xDlNcEXsZKF3CVbzWRyHga+Ir8g7ZyE0bNvTZNP7Rv8LzF/UdMN9TW4bajuB0lY
/0J/3lRoIbFBnwcgFQmxegJ/y2Xm0m/doUF3Bbn57c14lpfbdKkySKVAy7MVMIuI
d3hVOX0O82xqOw/t8LP7BYcxCZHJtLrzowPHvCv4odann7rBIdADzSVc0j1R+niy
cvt9W20O/H1oMxqPCq2Dh04q+0J0TCEeiPHCV84SbHeQbCpsLqP/A8ejE7cYrRjQ
zm30+hIn5pvwrQkWnx3DrEVUg7bgE0R5icJmxrA2+nBuJOUPgNyblRaFBBPBRugg
9KJLj98a2BEtT3QTZjzIe7KK02vhUXa3OwwT1OjE2DdEcaerywB5UgjR8j66HbV9
bNk/AVfMN+pGkQj7epuq17qfpUkeTn2eqh2zdmtbsZaP2IxsbvS9OV6kJbZ65TG1
xZ4HzPTKs9dX7htrvCgrPQchYftzKxH+rNi8uNo5phMzBm3d5M6zHbUdQ+M7bqmh
5gmPoXwXUyl5SGj1RnVaVvpO4bQ5u3lC+cMNnaR5GbsOHOR7LMLM0ThcQMJ65R1k
1aSGRBP6Dl2TkjD7E5ZkE/FAa/Yrcl/ovTBWxsG/UGrcLR5XYrM2CEgI+5UwGjzc
N/tlUjlrjUOIsw99/jAx0SS4HLAuOxuPZmHcYnoPXmFDIwaoEI6YnufiOgr/uCQu
7FXSoi14/8BP13SftACY2QheiVMC8sT1CovYAjxnBWnWUJqxQa34rBGimoGE3ejU
20niPsrKvQ2DYF4Vy+up+geJf+BmkgbWbDZWKJlMtMOgMIMpkwCwnjBFFYgkv11T
gyf3MStAZcc2u/15TwxMsAzrl3sNtC71T4f11phXgkWT7T0bllAhgYbrdmJtbMDo
D6Why7QlKL0jzDFwTkuJCIv3ctH5wo2mCfQU3ZKgXocAbzHge709z3FcUxaLn2fH
TcPw2bJLlexC2HTcQ+O3yScIXvbJicze6ypRxTKUibn64HxP/hVgj5SVY0TrlWB4
6QUUFVW2AxrWCrvlwStcOKuRq7E745ZNVcB6WVxx4XatP8CNSrNJMbn8hQLI5MjL
OyjYLmr7ZpdHwJLzI9pCDDqsTGIiJ1nOJ26VYS8aPSr4zjc8FNSiNykykNLsryeb
mvdwIVRfg1u0ULr/tH6yApBkMsPzcDYqqr5IHqhv1fJGM3CGA91uXyO5f+iFHobx
7A++VDQ2N6nLnvVBMe0g4HwEYDPYK+P9xF/+jXqNE9lbjThuebhwn2nMleLsieXF
EB9mklZcVfqYsYeqrg5c+KyVq5WZQG2N6DlSzvXdEaId/6755fEF9xAEp6+JebnO
5cwSnzJEqxGWeU3KLUsvRMr6/GfuFkqIQWSa2niRgCF73pVLbqP2CjaJ0j24k2sP
8S27oHtAb19LqG7MewOQQjWKbqildnBYUXQBix2Uod9oE/cV0n62BPrnJ+BcnAjQ
2sCj+vzugIhYFCPU5+WBSclWuX7nkhfA5i0hrzkhS60rngLBu5MH8YsGwEGJUsRg
4lJM2C2KylCQkoVHAFFSneU8B+y1Y0Cz6ZYMe0h09qcDzr/7jOrKmKA6a3KiJYKV
4mZrmhvQ5QE2iMQ+09LdfO1RiVe/yi5yTwJiUEPDeL8I7cElVWdrUcZ4hmQ6ORFq
HyMX3Wr5cdE/gag/nuYauCnHEzj0LyO1ZAoxwTdPHxTIe+IR1EOjfncowqWX1Rfj
4imiMvGh/pq24DSZlJuw0iOSHJRcSIApERT3R6s9OyZ3aD/XIJF8x47AzosWIzJE
aoqw68LMYJhvGqJxVThxtzgYn79EF+v8JegbDH3smG7VuNMj8UrBt2shidNttGFh
U0uyt7J+AdwbvRf0l0Mk0ckZ6RxZ3NEDO5gOfP+cdhA+qL7drXUBqtYZnnq5BcH6
myWNa3lfl+e3hUjv0H1zXw2VzDgESeP44bqGiYawd+y2P/tUugDR5waey5pfdhYS
LA9Ba23Lr1vWGPbIUFo+o+SFIvgFdExzlErdrH/X+iUtHHfmE7dkMoyej9E4q0xw
xl17Whsom/Hyr665a7oN2tPnQnUdclpgtV2KAlSROOpV/QwibKwB0J3Leu4ZyCXj
m1tk7JYurzpUNLy1ZqHjMaJUt1TIfzepSDiIxAp8+Q0yFoTB3e7GnoeEnN0beviK
ySH1hFnLwg9jh67lM7/1hlfPiOxUupp3CehjtUNsFL89FGLfUQhtlj+gMfgx5N7B
pCTMEUFH+D1XxPNsH3p4SYYo81t6+lrqa6Qste7Ok1Nc6G2ZEh42qTe9STVW0Uvp
T0niWcxGWEUIBjFxlEuMkGeybXvmk9bAJjv9MsVmiI7Wc4aQrTOEFG4eF1R8lbDF
wuwGMzm3RI7x4ZoqJUaeofHFDF5lSokLoZ0FbSdrHpRlNiDsq64c6+mHekWNx9Zz
dNHNMDTeWx/bKR+9C8BOVE/C6zOy7BjFjgLPmqRAH2Y/4fV/2EXGsQISfhA03gbg
amcm2EmeI7xgkZd4GRYtPSymMm4xUupdyWJRU+iAPst7vWuywEwvMl7DCFvqsANh
GfuSKkFn9/GDiz5x9p4unAhiK7PZBZXy1Q8WcqkV6a6luKiG0ytbuDmZahSEz5kp
1OtdJc1WUbYdhE3tU1qhirQ00lEGRIZHoOCJDmzMjUP7q6AaTEMTXt5VhcN9hnJw
TgbJx2VxkSmtam49ZeXbSuCbAUXlFa58gsZNxDjajfkOyv0dTozSvz0pjQ6vQl5T
7JuCz6DyuMv8D4g5IYvKrguUs6voEdW6U6FzE6YEeMFzvSaQOUK6xXHiAd/FzpKM
I8Zjmvc+MjlVDTeoqR7bM1kXtIw3LumLMWjz3GVWsDJhB2V/yKb6JVeSHe/K2q04
powbKDBOZ0M/T4WM29KSb9cHWYX4mx1ztN9zm3Xo2c/B6ckRh9CM7UfakwAcUoZF
YBDv2BhEuox9Zl9kwYhUJiY2+KSm+zlPKb6DbH0ABcNOJ4H584W8T+EI0F4mNu+c
UUKmtlsqg97RO6voHdCa3+LS/JIpPvy/wzqEdSDzQHr0pNQHiVaKduRWAlbbOxkc
1KI3wV2gWhWOhvpJi7gw05jGh/jFTMscAAxM2N55pVebFonGTbUKF1ssOIOTVcms
XgVYx10K/7eXBgYKv2KGMm0Tg0LlnmtY9MYiC2nTywfD/tQ50MdbTIFxnLXvBSDU
uM78KirNWsVpuuIIsOn97cqoZE8xTiSdPIZ31wlSkNjnjKS9AaE1uBUIxDca902r
llhlKMwsr5jJBFB/mpA71DnA7M1vdysqXG4h8j4mluUoR2uoeUm+EVsr8qbKLoay
E+xpW4eOHyOzFdge3Ae5N+qw9vQogPGfxyyxYsTejNxs8oro2Os6cPTp0NgwUB06
hXsWCt+AV0wqaAQrXgmEpaqnl3aWFrrR+ZCDp1AU1FiNF1x8hfFX8j9R2WLMBeUZ
Q46CtcdNi4oUtAu/IWKSqarGHzaMZCRoSvGWzmc+weB3uDPC+KJPqScs+pkhM3Cc
69D9xwH+AK1p4Dt7LScDuGF+BufyawmiYV86hqeL1TjaEn0XEWwo/9gla67OXxpM
stkcKK4cuczuYxZRkibkcBGIzDAvpPcz1nZJVWjN4HWpzLGyl8gTqfDpt+d30CSd
vmQcB7no/G6YvvSZ3F6wyKqhAR9Fge5uPQJmaHKW7kUOlUgNlL9LU4m8kDeuEVp4
hi0PSvYUwKm1b2tzwCDFMGK0CM9ln/JL+C1TfaoRzm6NyCmpPJQFDdhYtfoNlRb5
WrS1VstK3a3QXeU5BMOG0GxrUWOXJ3sS0voRE2FIlYR7WShOeqFCNExezqUoiegZ
OyxULflLjctTC+PctsKmcBaE3DHTMhnqZLKljXY1vT2HtGzBbHC3ghMb8fhk73jS
ukLSEEr60UcF/kxjNSjUU9FQqKWFJnyvhaMYRZi25jbyuaDhvF/qZRa+gzZujdMN
IRHeeWt7AP6FWVIL+nmcuw8AfGpUEySKAZC6lhahgERYhkyGpb1/PKi8qVYcATWp
C8iRum+oYIecwYObLjWtTMCNCqB++oTiuWW0/Oi8tXZ8Pc3gEysUww9Gl8Wf799B
nVJ/7Q2PjW6k31eJ5BypNl/v7WSwRui6pvW5wzCbf0Jj2XL/taxhxySQX2jJUVln
q0BY0hQ3T0fsWz9TvkhfUFh+lrlc8hLg5qSieBVdLt8oiyv4Z46N6ZWU4sAiy0Fr
abwTMZS5N9sBklOiyMx9F11gec33b/NjZWvsrj0ioWlUEBleFFO0xVctrDIdOzkx
+ZVhfeFQhZdz6QTBcEEt5t0SChrWirLqx5MjbvwuVJ03JB3QVyJHt/IZv81nX+y+
Uf8OgozMSRIzz5YWxlsPdMm/m2jdUF10eT/VorYob1Y2bXzwUJF/nUXqJg6wnGa0
H7t5CCVjSHs2Q1uixEABx71n5zaXXcSY/ZBbkzKD2njbSkX5xvydmDaYIPqnhDbR
25pQo31bULn1e3s2ea2TVtu9SR1hBBqKTdA2UbzfhRWOJ4amx124XUw73M1EVnR9
sJmsonf12I2SbW4KDy6/vARfNDyDDyWIYb8cJ3jxvITvX9hn4gZQi1jCtfkdAfXi
k8Lgq+K0yvrI7mtYKQn5c/Uqn7DsYxmADhqIyNMN5EDt/TxDg46LeRkJVn4tFb/u
7rJ60fnd5PXkAYW7QsxT9ekFQ2KSewnLmEYnBhi21yfxNrfU614AYj7okNwuE1tU
F7GWjkyf5OdmCXCLhu7s1FgSlpjyF4GGb3dEd7J0cCUXIGAVuQ3eE6YR1BDMYJ0r
MtFrUcwiUQegTSkUUbXwVjNPwUy0qVZz7gF28o9IZxouW00a/UyFJ/wulSThZx0F
s31C34GTqdDiZLaQQNdcifVukUjhh8Blb4BpgRVSulY0CLDtKjUn0LDQqqCoE8b0
VNjPc6o+xvLt4tknSbemcz22RmIQFCldcpMG5d6a/G5FclBR+7l2WD8shSk4sHe/
qf29eiG1+TfG3COceq0buROW/oz35iQ2ru9DfSheKx6BElnQfxIsF9r53JRYmjJZ
qRjJoSOAKXvYsTu9l7H/6hNqnlLzRBC4aY2Y0XWJX6iw9xkykfG4JxPMC8rBn6nG
t0HEH6uEqBxUj066emTSRFiQhHE2DW3YCPenieu63vdOIdvPUp6lUoPDzdR9/B/+
/snsZR3d1UNDdW1Vj9CehtgVheGl0tKDpJzVPnOUM5f/SAeZt/0RsiSyLRd8rBx6
KXowQJFnbVryNoI++FuIRGs7yRdCaez1b7ig2w3Aj51dMrw+Mpjw5u0HRFb3X68v
eJ6C9X9GDoFeDFVMD0K4b7m3gKlySGs0JWmcGIOrOMBJX39WKlfnr6q13esaPXOH
L+Nl0xiPgx+bjspn/DyhKbuqNRllkYH5wE+p48X7I091QxbqmE7OsaHdDigsXNSK
xkgiIDEabgGvBH5hCrSzOS6Qz58IS+TfZuAVrbsCDK3jomxwO1PwNDWajKOW2sCN
ahqqz9An5FZhTtTfgr3RuFcOOaWSZFgBZwrycOQLfw1IgLs90m5DJOzPaI/hZUdc
LmMzvC5pfi3aeG1BpN2Vc4BJh/vEqcKaXlIWz/o/HVyuNcplGHcLOSwZnvLeRt49
2wZJIHybkh2MvuyzWs4Z3O9rFa42dis9UeuxEFu34hlrKtsb7o/ndEQMz7Z324v4
FXxzCr7gKf+4nBCoFFf+b5DgE6iQpCWfSl8AXjzZlGCu6bfblX9iNG83EQGg2Q4A
MddPjKYie558uMsIwojqiPSHzSCKyHRdEODU5F1ZzMf6J526JFtnyeDxEEfnG8LU
KfhhRBzYcAa5zOLoF2zkUicqlJqnus4AvHDUyAW7LR28hMRF04oBrVeD04ICc/mL
YY3B0eRmr45g7/4VQVJ+KquYv3i1E3Zk2kIvN1KLupG7uPxrqHmeR9Hn2Y69s6XZ
GcrlK1tU+eshlC6KNCiY2Dc5CDxKPmHGAFQS9X98SY6AXbyvpaKi06u7Dujg0bZD
sU985ejxYxk7aBbUdyW4JOPHdiTdQAh2KqgPC7g/g6fFCUXAk00UqdGWwKg0R7oV
NbmXPOMmceaDusC/37zsZn846Epfv0ar030SWSTgoOq2AT6GbulEB+mkGJyqoVwE
QJgAfabjFqv/n6AAUsoMR93DqhAONVwbPOwh2sCEHA5WBjoRUl20YA0QOcLCO/ix
x3lGSJ5ZS+P7UP46afLJSRYQ86SbhQGHtHb5K6bsaAIsJiG1h2GLXw46JsLRhwBs
F2pM1TMX0kjcosBNpE8rFr77adixUTYXvT02oJPvaCbzeV5tk9qZcDj1W2/W+Gtx
W4gcvooCC0MHcWG3tsHzXiWWpAKmRCpQzsvWHQJt5jgZaDIyFBiDIKgxR3jJqzqu
JJd8GSRYDZL1TbzSWY8KAeo+LaId7IRhq95n6Pdz4ofPVT92nro4Tx4vnaQiZIgt
eQLR1MT5qTcr2I0hFfROit2a5JjT2D7q4TVT+Ds4InB5WjYLSYM9vR4ecuim4KAN
ywNRHz4jOAR5jwanHVmVFmFBVyCfzrLj6Ly1c2M0G/JG7E1WOS+yeYCr2LLZahw+
nHAoOJn/uznXD9a4ICuwM2+Z0J5m2crhROQks8wZbxk4peRLR/RpcvHGKiJQcD0u
upiaI0yX0vJ8m2M14h0xePAogXSgkNKrvH/8NLjHRPcFCqyFGlaJ5eWtNm+nf9rn
+4QIkxn9nEGumFG87wEnMHCxY951AGvmlonLaKIaF2MEP6yB3gAa/6SRz8xoR8FO
h3CGJRCpTsj+gN0CmGgwJDRgnhS/sLVl0D5DYUc/YHAwgGNTTQldm6f/+2nM4pg2
cn/Jud2QvlKwYkpNCRzS+xshn6c8ho4lF/3/SCkkntq76/Q/rRQM1rZNag+wjEiS
qowT1sukZJ1gy/O/5W9RSPDOSNFa+xqDEFswPBppa0Psm+dpWBlv1nQWsgJ54zYZ
QbjOeVU4ptwlj2QuI4eOFXs/KRysFBX9MzNYtXxqx/CqcORPTfLn0kOR47/lBDec
qeGE0SzDxr9PxWLeEt3DBaaMpJ1OtEmi1ml/Qvs2KliyRoVQmvPj1s4jf+4VDoch
RLeUKX8ctaqA3YQUo9UxeNC358ix/hkDg8HNhADdA7Z9neXHjjRXXJ9y3fJw8bHg
Du9Z5bozHpu3za221QtHhmmxpXUHch8+bzIHj59ep0K3pnffuhwtAxPcHtdFMTvj
2/aLDkRBqqClPgBCxYb6i0apAymvwsFJpdcbxYl3PLLQRKRsLf45EUnEPH3X6V3y
EIP1A17/vtIWm3GcuteUQDpBV39bPrJIF3nN3zmcP18ktARaHR+3imJDmzJcpenW
v+vcoK9w8s4jruzEBGZmMCDCFDF6HRi3Zn4r696TB9KS5vuJcomA7bI67jvYNY34
NhYuSm8HTQHcPMHMPg//ocpE5jip8cPJKt/5w7GdgulC3OrcY3eLlV5T/TyahBEs
4qobgBgL0Q6D+p2G8vZmTJlePmbVasLolIF+O7rSsB3xVIIvbX6SR+FoZ3jG+nli
bsCZMPVK/PFLf3hqOBLzLWUhFeQZillApbdRkYjXfnpbpCjR47NDbuIJ6lkfYM/K
D2aVB4OaD72yWYceZKxrvAwiKblcBaWmzLE507nxqgvgroB6yGTsGL9GXYDsVV2Z
FECSCMYYGeQitYAzwcN9+B6SfXj1RuhiwSPdTgptxeHEnuvZUIcac812Eivs5o9S
T9l6Y/ew5R0rGMS5aSXfEF7SYddPvYssCT4odYG1l6LuegiM7yqS42PVP/RO39uY
9NvlTCLGJN2mbVLWvwW3Hl+V6Zok/vNHF/k/FuteGqWkm6X1j/srjb/oti+bkhAc
q1bmP+1VMClFAiDYDe644Qx/29HOaP8kGmtr/Y5vHL5QMfGqFL1fhg92yEWpp2+l
F6cI21HZv+UtiVYOruU7HIWgkdHUr7A2vxLCIrv+x155d1tHB5GJ2WBTNMFeoEp+
PndBtyBsLzdwQszKzPSb4gW1rBq+7g7szyJI0Vboc8KSdLq74LOn8ZtzWnaPcA0l
yGzMO6kQ1atzFBCd4UXI6FtRL85FWZxf4vNSpit4b1g5yhY9+rtLwyq0YWBwQJkl
VD3PxURkiYsHi+FraefzZTt8onagMJhofUtouUdmROQ2mq7K8cbSJkqp/xyMaTVE
vsmlkHMwwgln8S68ngQK5z+6WHOKIFf2hxuKfs6w4Y98qb+52/NBKakJbE65WuOt
/wxBtLNKlfKXwtTlARUtEA7DF8rOAnSR1HFGu3hhvxq77CcKEnrN3PEEhiIvzE0J
DdgDX0MTqI6kYW2lFn5C/HGGEcDdT0X0ii8r7EgTVnp0vicpmJfkliUg2fbLX5uh
ctH3g4Lo//jv2jG0ZwfLk/gstUV0erL75eZnZelAwR03XKmNIVrSblNSpKXK6TMm
Y1suqB69ihakPTvA00L6LPI2ooJnPVSQyN6ggsoTQhxrB25dS/jIY28jvpNOUXtP
GpLb2XDZEMV+4J+P/TBA830Fm+Cc0R5Wq7BgAOIQf76vKQtRI5zr4yluKqhuuPXv
Lfq+0Ix4q/9g29WALSNikHMXUifGi38voOV/timvfLSimmjIb1VLu6e/43hl/g2F
8wEtk+Qwj7kX/89AWCOj2yu8VptrCPrKVQe4wFQMChxpYcNJJ5BFid9CEECNqjm1
3WRHfPQ3oS9k7KEf63/ykZEVAruiWvUTtfpKYMpC3A74wwkW3PeVLFWI8Bz6RaaB
AdTiz0Kemhai8uCBOJs5T6gOVYwLwUOW7/JYOY3uxEOSVgez9DWKROj5PfRMshx3
avYqv6sdrHr/3oIH9Mnm1AGVyjjVQRh1odhXeN1AsaEG2B94Q8zdbXJC831BeJ8e
K2LNvQ/H9vAo7rHMEfgUaAMOS9pSNzGfK8VwgG1LrXLURyCU9cuDGxypU/Kf/w11
UbyEqmAtTw4Feg1ZPqJ60glYS2RelvvoOmhc2nkuVs5hg2F7mOwJZ9KYfsLEtNjS
nnpPnfXCgcEzWtGNywedqxfPKUt8inqSE3aGtyoJaYL95L++HoSq2s8vFR+PHY7m
2eS1/ie5I95D6mDZTdJcVXmSCdMIpNddX8nKHXaf8HeYSNs3hfqKr1cAfGfHyMLL
8A4mDdudqlrNyPYUgPC8cSCltj48TooOnbYBpZH8jwqF3akMd5NXUQYGcpi1V4F1
G2MFSWVAF+3E6DFnePRU+50JoitAzoCZp6VZHmJpx1Q95391zeXSG0xR8VhOuWRk
Yzr2JhtveYCdpchpCI2WGku9GlOOLHUXwkelZ+UPnZF5s31VkDoYG3rXgMkkht8K
t3uLqy72LBQmjUbAImt62nftJIvJ5nPe0ZRbODG6CFAbbGXBJZguxXdJKZb3EYwy
G8p5oHcfcIm0jUn2SDXSV4K7ZeJtimVkY675b7DWmKEYcU38BU36OBvIwflevCmX
9yfH0gCrxe19xDRYwgQ9yjg1oJjYDERSUyiy8R9hobKYiq/MWBIuQUq5V5jkMvtt
+k5AfinkYjXj1SuHyLJBuueJWULz5JppRMCdD8hVM7kD/u5lPyPWP5q0T0hn3QR6
ZTe/aPrkl2hFW1Xs+46OaFad1UQPB1CHPE4mfwrdVC7YqenVcCyPa+LtpbaynI4E
YrvQALK0ws7BFzJ/ziYWx9Vt7z0IAeaOKi1gEvVJWDArXUx5/mOID2ovFFdz6dgb
c6KPcT56RRMhpuh9PP+LGAj/IAZLbc9TXSepnsMt3vH8xFE7G2pZxTpmlW9AmOz2
Q43zTZlY6zLnSaskHB3MsOMEyMT2PaFqtwL1qmPwppr+93mpSnuut7X49yXX35kH
UhYMeFASraHm1cYRTqAvzr8JXsy0PreVCkA3OeBbNPXI33TfWfKNOQL0kebAn/U8
D40LLFAvZTT+kcuqUAxf1ANmuoHQjMAuUzwWt90FkT558Cd5sc5k48bQ9WSuEd7d
ZyJ25oUg3RwnDSIxiEUk9m/HayDiE1+4MeXwD3U+YCLqtGFLggQ494vBHDtlGa0k
co65ciAKvIAl5qY10v0Rc/UVLGvD+Mte2iS7T/sWEIsIgSEoqCvqftuwSDx6tVko
45UaDDjkf0greMsFgtyy9L7u4Dm3LskmtkdAAsJy0iS2fFcsuV8UmfaLuFf5IIQ/
3Oy849BjWnUJwY+86Z+/tTiXhjABXtsXQgegPB/5STO66c+wzPfiut5nIhLA8cTx
qyP7UPChYzzxlDYbaBSkH9n10DEzUUTQfeBspGsKFdLPvS9fHumeT4F4ecWCevtf
CsUIIO7EJJQMoKwUlpVn85eBLor98i9HnZKRfPxS2E8S28pKTGPJFGnLbs2eYSlx
FT2McrzDp5QRhoyDG12Dqv7ExsvrLJKJ+Y7ImNaeKOz+0RGlW6ZhGA9KUCXyeAt8
QA0aqwNQERRxqbZSrdpFmEREyS03w0v/VFct+2yDn6gnFuU2IXfWZX+a4sB62s4I
hm75dIvaioQv/A8nRq7JgMuInk3k4tDv9TaHRgJZbzPGmZSrK9R0cFRXF3vYRWcF
cEuq5FlgvWvBBhaCwly+Lc7xlwsFYq7fHu+3oWiD5/w1M4NMFXhnXPW69DgLxYJY
PdLSdyv4GKLWZN2s1fcbDgXSUgXh/WMPG1Hz+8wKGFtoOokTems0WfpK7OVjPKlN
yyr11AAl7V//YgkvcRh2SUEn1XXGbAQ77w5nKe+u37bffmOoUNL87tP7dwIP6BiN
KFF8AsPPeBFQJNFW5mUfkn/BstR5IfYAkFWtUpnqhWhI8q6nLVBWsadmU6nszijJ
IYzROHothWJJjKxZV3mZCTqX/8XDrnJjhkp47w+qQGelYzPsdMi+5EZy19Rrlo4t
bHo9p2VSigSynUeQO5VNOr89Hedsl+zcY0FVu6BZxrWaGx5fPfLhVIxsZv31b5FZ
reLPbV5cm33rpnimVIi5elpR2j66oRfgtUyyjCAI83ySI3MSk7nzl6iop/1uLBQk
RFTCYwkJwIa5rkM/8eKcxAQFwA7wnMR+cdoDdcBAbYVeW5YIEe1Pii16kbxwEsA0
giXVLDYegnnod4Ksz32ZypCbsNbvw2YpvAEuKX6dipYXdu+06QhgsitF2z4ph8Yn
7PyjDlQEDPwuk+eoo8ueRbwdJumMExMhghXrz6SG8cxKz+lcC8gmQn8ue66Xf3W/
l9Y9J7M34A79dfuqN6NmZiJIBCxX2DTCGJwrnytMJPiEwu35BIi7L0VrS5GfhWLe
5zhVDJvUtGzzmawmlDsZkGWjAbmhgTF4egc2Ty3S2s1VtlebHrwcAZsnXEKAU5FJ
WLQYZUTYrqfR3t6YMnr4pcs/O26fwo8glsMzpC/ThZqTXQwbd2cOaq2FwLEo0RTK
jQlcXi2/tBerK3HuSoGPBNvR2mtJPXC/W7BFyAK/Kx1cJSt3htKoz9vzEE4kcV1B
9YPVDosvq9b1JHr0NCvd42WbbDwlwPYU9kA0OLl2+RyTQuBUkBgRWIS6lR/LNpmY
obzD/rt/KkTReTBZXDFf6zkNdj9J5niSKcE2ihnjNyHz7AahAO+gOaO2Ng0uNCzP
c2mo6fqyrcI7Ps8ZTP8hrcEHecsuXXXEn5HKXQV/vyTEc48t61GT3gGkYwyETctm
0byGKStHVwGBXMUnH7RAHF14D8upr2E6HXnu1bgYUMI/il5nDwzcmaqbMICWgmxj
l5Wk+hQFLSuM0/6i1dZ/YMjtGzaHarFUE42NvCiWhev5kDsd132Tu/HxmGmoXSUa
W0Yy1+GICIYlZ92Cdbzvh7V54zKfpctEWimGCO14SywqpipVp3bb8NLdbX9cgcQ/
9M5+eYvbMvcv7We/EgJj4DjfBsv984tyPWbsufJx3BKrC2jJph82L+Msns+Gy6dE
hn6Ve10rfJZkqXa9qky5IMOWy43pjIlaoE9CDa7CgviefmoLDrqYyjlWLlqzqTwr
RAmmOtM7DLZAVnAdZdSjgwvOR9PRwod3CiVer/ddtjTFveUxQqD/nnpiZ741CbcP
gjiv92M9FAmfojgHNQlm6+fSXpBG8gvRaIbuHBtYRHne87ijouBFEYSercRHnIkO
RV04JBrg++8GPvVtmO02HgEr8FQ9MvpWMpo6JrWq22mm2/kqdMHGXw3uO7f1kQiF
n14Qx0/0acSBaL8JT2WYxC8nVhkrA4kGQhZzXA1k+wdEC557TI/HdWtyLCg3umXn
CKhVngK2DYa7KkQvilHCRVRPTWAOPj5TRCblTClzegsSuMueH2pRidOykjk3XAqc
ZoG83qclXLBlIUgq3m4HZzajmMw5KtRCqOyZJ1eo/yfKRmGh/kwJtjg+5izNtOTD
TI+iPajN7vbfSge554GYLoxlDpw1d9zMQOm/lYZ+GWQWMuUnkGgzbHToj6C/dQ1G
SSvg00nsNTdldA+GdbIMxDPOfzGqv5rQqnIvogzzls2hAtUNz807Wg0Ma6LcrwZz
V+HZEwvu7EWUDilmyV7F2PMaaJB+CgWVnVFgS4LZ9taGDn5ZRXQ0Zjj/HjSR+tme
NRc4BJ/WDdhSsYI8ViSnNlyrFgxZZijEVt+f+x+pes4mY/hK68a3JgrrS1QNyKwG
YJsocgvz+aNMZok25IhZ47to0843MSIacs+0GsJThjvpqvVQZNoqHUbTUgYKkjeu
8LVuOvlAbZGc6eVsEVv9hTGIdWrurbZTtWHrvgQ7p874h7JTQUKp9wvimAB9XFIT
QvIk2Ct2b+mnDRl+62t6E4u3HIkvn7aedq28CRERJoihSQqh5IOZ+noqx3mooxq7
QKNjsQMgiZhkQVg3mKN3dX79NMv8hVmgOH6AdntGPMuwLw37Wk0TYfkB8jFzCDZh
jAGe7LdMA1FocqyNKwkjqXfMCszMRMqzkRUqjzSFkA8VS0X0e/NXJCAeSVjLNjkT
7K2JM37V4GTxqAGBYvWzvBEr3vdeUWvfjfSA5RIbo1Tpl10eG+qOLfm8pa9K/UDn
8j9WAjI5l4b+PRA65utd9yrymQgAJ65MU1p4AjgrqxIi0h6mcKK4U8tS6WbKFG4A
7VjWE1k8A83m3TpDMryTyZAzk2bU8+hzPC1U9FTPHdYbdQHDaGt7Bhi9aM5inV7x
WVe3rs/6NHkIKFPEG2tm8F0E2deBeFIg6GqyE9JC8WHE7WLMvcw5KLTQ6992qhqi
a2avgRVJUofgVwv6ie+HF79R1STufFLhcajVzgMM9P4jtg1rAjyOok2Z/wBO2Ui8
P+XKbGf447oBtHwJd0N1u2PqeLAP5SAYV8tHpzQqjgqhnfVGaP05r4k7GKEQMse/
gH8c3QC3jtTIfPrf67uSK8mR0KAZSUFQTW8GbnAHohXDgaX7U4inPOPlG+8NvVqC
2GRQ1SwZdPEBz2Z0NoNPvdHEZ30e8h6+QTEjsFurEZntC0DTmMkByhHOm0K3x4iZ
bG5zRuL6i8khh6oug9fPtbI43qDj6nIptrT8z1rGTyj1mQSickT8Z+Eq8FEh4L40
mg8L4IKW1n3WAPJ/2YcC/keQm6BeFhA/qbZ+SKhhaAX9thfy7qCbWWoz0HFMNgU+
EI4MCwORS7RMTTyT0qUN4ueovi+fxFjWqpgHLkPdVq6d5Gbw/eMTVXiCxBTwocrW
ebZweIhMg0NLpgmC150UzsXROVG4a8mMRUPL7YPSI84WwwWOna2ddjB3Wlpm4WY2
paMDSoxswogfKTtOU8jR0NpZ88u7AC4q+k/+rgtyjJQ37tQRJZPQNtb2QQbDOt9w
Md9OYAJ4bdO+Oy8IU2KO7Dt0sa/wtqe7FnbWpF57WmMujRWAJSEnKo+BuT7GN7Ck
XsuBH8hdXoyBxpBoPMD2ws/byA8rPwEzH3cdpxN3BU1GOBzT37eVaPEfGRP2kAuc
eu+xxnEGWGJ+11nybn+MUXp3VC2hOuG80dxY0iGsOCysBxIUXBMJYmTaIxRehpQ0
a6DbN4CEqPv2pHsCc6sohBSaKucHIARiNvz5is8rsTCYYc5rGzXwhNhbuDi1qBWU
hSbY8ssoPqLsY3xIlhV1IP2EiaVjJcJpJW4Mc3kh+vyh/G7o7fQRMYdxj0e0K29P
9LGLUXt7LccEiUUEbRD/tLVjDVLdQT3D0CpLV8CctSUT4E4BzGim5nET4Wno8x6y
xcW3B+M71+ILHNVpuAbPswwp4U4jYZJl+kstGF202yC2+Pv05q+VYqr6BQTukQxm
NKohLSfEwdZC9itr0SIkI1VMPz02MV6mDQ3MzE8lp+ajGndEMNeL9zNF4aRdf0dZ
Qog4IRBoH7fC+7qHEedGuqIiYo7GQWEgo8zejDR77hMO2WFnPfQifW1HlwaNB0lm
qJQ8XBX8WgY/I7GstxxDip4nGdCzwoSXua3Q8PKBn6TyHAJn0b4uss3aS73ZmeFX
AH6gtpwAlPbV4wXn2UHjp81VjHFCXtIF99q94gfdEOtsOlk8QzqsMKRN1iSrYxbz
IxTuWubNFJjR2Hnpv6tu7FaB1Npw9AWYQtWX+OkIkSgtif208+W5UbEKY3vPMySY
Eg+EzQDIICvHu9DDa1mUuCyHxHrpw/2TUeHIzgD4Ap5/c8VOy57PeB35+R9kUjbv
rF53T4xIDBuun857LefQY01ifPaMaPWDAtaKKhC1Ziaa9KJy+dVEfFTVP24aUM6S
JoRKVlkWsHQDwdR9imMnm5Q5bC00DEmhEFRhJma6onDx3Gs2Vsq46KJ4m6Qns6zy
q3+ZSaaj+ynxyA8Cnydn0nSdZgKZfJhHVtJyb+e8fQM078mW1xCVfxYP6R2lZB2Q
VN+lizzEcYRXK0ocrjOdi4HccQRGuM5oRw+xKcK329VJLxILgRjgkHsrGdS3gtTk
9e0Nuuc5LS/I9dF9c40Drm46J4pywXER49icvIQ/BirD8VPo6LfcurD6R85CvB8Z
6fTi8SccHTR0xsBnohIUJzpAgssAxBXbkSrAKwjV2fBCoNp6GdPrpH2qyhlFvGfQ
HIsuapSaxBCZ4k6vrh0nIsFsVQDF7b4qfOLCQM17rg7lN756eMYuGgwj12s9l9v7
PkGbQdePj/sevziTg51tpNTubOOdIeGtD8dRIe6sCQj8KI/4NdSk3SK04OV5zgfx
w8rTsJ+v6uqlJkXYctpWn90QddEEI0TPc0rQk6htHrU9BbHbKeCLztcyJiBddN/N
g0AyeVPzwCYTiTZgR92HWbvLZUuHtvV1LFXQ+PqWM8c1rwQfY6dDo84a/UAIKuZr
uH1JaJDbOf3YBzkKslwPmmaNwiVULKl+hFJMnFvvc1JCBBFlH56Mj5/RLm+TWWNG
8SnUdstYzQ2xL7ggz763gztcctWM9T061S0HFN1xc6whQqHADfJiM1xIdyuvkOT2
jopfu5Y8MqxLDCf3EbDviBVSRkb+5AbDUfvcolRwvEAv1EBceZHPHFy0JJMeV7kw
NZbo9h41PBGcHbUt8+wH0ueZUWbE864Cv4xAM9J61Lxm1pmHvFlcL/qAAcf8xEEj
+EryQa0KbYdr7fPPBfYZUY55dLhZhnBgcAxo3CJs1JzXX2ysLGnOTuR+9uktJknQ
ugxhTFYR2uX09Io3JwjQsSf7yBhoOROOxQTJDWv7pE1/8DJuZC1hR8uBX1xczw/F
+7ecfq198U1pb6cQfUGK71M22E0R1zWo2UBgaw9LXZ1XiFbrFaZ0GeQ26KaM6bEY
isqLQ93MwBYD0toqAwLaA9DO8ilQk7Pr26BunoBJn3TjyoxUuJi3yBifCSCl4kdO
BGhqdlN31ZhZuO4Mdxa2q5K2iRrdYd9o1Awo+TNrdlTV8y62R/FHgO2HX4DaSu8X
/x3O2sOE4Eao2MeLNCoPn4uA2r+f4Ovz1mE45BgL4bajCEd73yXHVDFe//P8+wLY
lrlkH9+fXEqIr6UR2Rs+0V3ZFENyL5VQeayor1sKPEesnhnWOgmCGupf8PsQVbyc
TgbErWKoNjXKeJkkyLWBMulfZpXoud1tF8GR1+Resf5zA5/OZhjBRoIY0AHbUoMS
FdL4y20t5ZATwFH18QkjdPyalNka+4a0rrnF2dt0BBc2M1W5EjcTLE4kXHIGhXJw
RDE+7DWQA+cD1hRZEfSK0iod9Z/ChhgDxsF8EiaOol/V19+RNJJasCH6fchbgpEx
jUcvknwlrKA2FRrAaicJq6PNG4eEXkN1yETl8c7JeDcnIcrd6ZhrZJoWjxtqAguw
3QRuGGGP9tR6c2k3K3l3vv53FJty7VkxoKi9FL5TZD8GpBQDtksTWurtiDVTcv08
VSZRoPy0AbScs55Da7GQh9ol9R+qh0WXncWxfqZXGPuW9AoGHnFS0wh9SlVTz4LK
+qStCc4WJVTzmYyltUaZCPL8gZf1E7ZP1cU+QZLousfbNWYfzgGUJdBLwdsQ0WP9
XNerfianaerKgBNRMbDSaSnHMER41kaorHzGwxt5AhmzMHKlpwOtCQLicNljxeUw
tpXEPqjOXz2L+zSZZyoMJdqKqM5MG1wUOZQrm0ADt91o2DtmGI/lnnO/H1XsB8fv
PmopyKjlXaKLycz/5yZ5kPkALwiRImVPFkdAn0wdx4llX+8XqLfi4O8MjdxKz1iv
CCVw2WAq9jaDarEUljjNNY2yksfq+2Jv3qljdh2/ZagzyXxt88vv7pJRPKXYIcvH
QhGVt6TX2XO0+jNjXW/vfvQHa6mUEXtWXHMtORPUA2fRcMQaAw+acr0smv8KpwhG
BJHiHCHjdzAJpolXs3WajeLb5V7s/jtcFBi7DFW+pWSig0PS0YzPoUnT5EcsC2E/
UQGi1uG+G48ghknCq6g8VyIdQJMXLql7KwnWWXGteIAP92VJOSU8mBLxtXe094WP
0YchErSmiGJL5/Q6cGKLb3XtGSmw4EBcbK1KKwdDC8kzvbk23zMwFWH0v7YwJJqM
ciGGb4F/7q1CvmYpKBtHGhjhyWtguNJeNCuF/6wvvN9Wt9OFydc8pTOd8VnalhLx
Qth+qhFCn8/EmP2UL9kecWq+RzWyKtOjRrfx4/U8M0MGzuEvSivtdCssd5MdaYOV
VhuEMd1Wku595GXh66miLOgv9Ovb61micER++a/7rfQva935ypXJ71lRPyTSDATq
ID+iC9wWY0V4ic9NCZiE/e/JdgmLrId1DE2tSbNKatI0UFP0X70WGOCaxsppxCoy
5YNf9Yf1bSACb9lxlhleMb8xaYI2pc2sQ1HELiDTL9m//MsN1IUi6gckdS7ZYsWb
z8aGN1LNvMcNPX08eU0zlMSGEvScaNNrDjDWBjAkhVdOcJMPaIE9gSE/RlN6JeoA
+iTy1AIgSxkEdIYokcFzkUDQ3Ob1Pk+7S47VF48hmPgFR/rgvu6kL8KZ5haxYt4z
l+CJ0EomQIRZsli4uCfJeLD5donhtxREik0Cn3WJoxX7Bjpd3N7wDHiLcG5uK8N+
zvhGy84zyaL6u7XLVfPKnoyUFsZ6NeROH8/Pn4odZmLR9LvMW3Xyd0HpsTWh2V/c
qksFiKB+/HjpQ5I488GjsEDhXEHBBnIwZKmIgpbXu+YFzMhvm3bp8YlfcrExJlGm
Ner75vxVmuQHXl/6DrMHHDxyNP4CbcbZ6qWwOQOPa5xM2YsMz9DUZMZe2SjGCHCb
+3kg3V5GUFWoNIaXHgvpBIYnkyeAP/zLHT/owisbRvdwMn7dTNzW63UiLOBZ1AdY
vIHR61E1BFmrXoUexw22+zPku0xU6zXwr2nZIf2zF+m0va3aj5Bs/2g0KOV9JysI
SQyEYNuUDJBdslG/vES85nPIyc8DoqNh0HVWKLtwLWx7ki2cDEJlb+kSEU6DHyEv
VlkmphHRDN3t4mm1r48nuFQsasyerZjUl30/7L680d+KkBSPtkPuUqKQGZsJ1Odu
o/A5sD51uHNqN86T0WuWCkS4urV2l6XGJHu6MxY5AZKh6YOe8yyIm31WBTeuJDlt
32YzJ+usamY2k0nx/278mZA37w6qxEpXSXwFfPVxXJ749ycCQjivPlDIM+PqBEn9
c99lt5N1Ao4spic8GjwyzFPK4a8Dm8m9OAs59RlxR98s4uLEhn8qbkNndYCdnxrk
eGNL+woFXP8DkAUQiXu4te9TASfr0fuoWyffv65YTie3MS8+64zoNsFova4NDens
eUrmUojzPxdU4sA2zhTrgVuKFbPiIBzV5LaDxU2le3SSdYJj/HF3pvlNNiNs+7YH
vjqlPidIeZPe/wkUThB/PhZqtK11E0rTB6x3cKnsLm22S/S6DUBHci2gNaQaWB1U
e6hheypluEhnNmywf/ozkCc25nUjQkfCWELjtETEGfz5X15GsBw1w509mod4/6MD
g+hnGRPf+K4m+KBvm/J6o/by1ls4UWnjPeLPiDteDDnIVNAkxY+I3iaMbmZW+gIU
AtNrc7IFRq3+8mf4vFciS5oMIi3+wRT5PjtU6Ai+WQWeC4dxQG3NIF1vZgseI+GW
5O9BDAuUwiAs7T6t0cRtibkOtN8JzQzvQ1EWU9tg5GitoA45swjqe/BEGvPcWeCC
KXr1jVFASqYfOSO7PaLeYqA2e0z4Z1spRleKUfPa5WdT/Rn9Mir4b6ug5uppl/u0
NGAgb4bqSiPLrju8f47EOeBj5jgWNCk1ZK5hg1qnRcLzspxCQ3e9ttsxEdXWAMNz
HFmQKoR9X7LzzyEbW+uURfMmZmm6Ox9+9YmCYUAAzs7FuMpu1oR4XtdmpGdyFZif
gnoKqvEpg9tnO8gfpq+d4P0WSrkr4QoDBb4jiaIiJH4rPWUXHJRg3bmfJ1/RsCt5
Rw7t7jxEhtaNL6e4Xr2VJqzJDsGVBrB6MEBA1MpTGzZeXXD0x+9VU7HMJLNR8115
YVP29P99RlxIX4kcLCbcTGgyrsUzQU9M79Hv60W7fSIXsznAyc726SKMj1NfC3P6
HVSGllX8CwNTYDrrBm5uJeOt7+MPa7q+nfdgOEUIBM6Y+GqHHxW0HfmJGkigMHAM
OmXc9htFvYMAIFkkawUEOMQphcuFhffCG0ZMF/QGjaC87J9MflzOHq3pJMNQW5sU
395JxJSUNFsfR49qyXkC4R6bRqJW55EOYxQ+qTrXm05bd6I3U1nwMyKGKyhqdLkL
i7t7ZZ0NgyDQnkZHXf6kucrjsx/0MG9VXdNuWk78/T5mzjHtWqu7j8bYw7wu662V
kYkyeGCaq892Eb3hlAKmur5D18DpcyRjEIbXebZ+EjTw1rU5/XGiJOKV/7ow4i3C
Y3wnomflcAo7a7GbI8vnzLU4vPCw8s3zwt7YhLk8w4tUCiTMEzZgFpFoMvNNQhMP
zq8KavVb+aSZs/nsA7S3PVOnTpVrC1A9jVJGspoyS5MYMxAFrZSxz/HqCmgXP4u1
9U2K4TE7bnYnhEWpx4ItK0YwzymiOtSG2ugxwlyz8dpnrZBszig6/cpawqmp3MYa
mTSFLb5sJpNgeu1ScGrV0PfjvxNM/0/MYG7nlXgWMfX1XpQQKjIr+umTg/9fh1WY
duW5dsYFXehnJg5+1xYvEyHqzm//Mh+eleEfNdWOClPh2FUKsoD5gA4fh5T2amQO
uK1b6l780Uj3y5OKSSy45/KbsvPcdvYxgQ7q3N18qRhplMx8Fo/Mt1VIfQPWagrk
5dJI1qdWj7XPhMt7X/90ikjQe1ExRwumO+A30nMmPwONaU5g0cujHXJ3UdJyLceF
pK448yjxAB/zhRXEhC/xrPxn8d6A8BEuDXXurfjCbqY4UBDlcvGDnzWMllTIG0c6
T+vROh0ZL9ebvfdBMndpLtxG53eayGDdl+j+O/1T6Khyy6pOVSdVRBT4J9gkFezl
OZ6Ij6mIBwpeY4l/eVz3QwO8zHAuTYwabEsLojdGwjErxYs2c9WiEq58Dvyq/H5S
tkdc5AH2B6tUiNf143/zZmkr+7fycI0RIvL/KPnyKUUD2OzV691LqUvZM389osad
qQGFY57WOarI6T5NVRYaKHMiuUDeZeb3BK6+3E9rHRL+j3RJ17O9O9a9QZthYaAV
32uKWXTZNBYkKTR++XXbKwlFVDQgKKs6HcUxk1ZmPpYD8DZfL77V1VCSbukR2DQ1
ROnbOts1KHLB9W/yN7VWRM2BUwGhhSQpWhkwySa1KGcqU/c9wdE02lujNfT8v01D
ZMVCgWewf7124JSPf0JpE42RJ6QOtyUrXXqgpfeYnBToa4Wz11ntJJTsNLrHxskg
CYoG9WEy1lVwUY65k2d+Y7mcZMZ94zLQXkijv7WmbQsBOy/346LFZM9bwrg7hMnQ
RrApynsVEbzDIWs3WTJRy+GvZz3J8Nn2s0IO6nA4LYFEnOfNcH2+72QaiypfqFzr
Ws6xL+Gk26b9eH6BkHMnKQHbXbPexuSU92NqSoSaJqrcM1I8KRZyjC2QO6asURKi
C4n1znc5D+myhhsanGiseDrPGDqPXQBvhkgT2FjKBXJi5GsE61deei0zjjqWXKOZ
MStJauc/gp/be29Fn2bNnhIVfQBm3LUOH/nbDfttFVuNKQI+PaWdhrQzM4xrcb4r
HMzl0qV65dWW7IXEcElAskzvf3U+h8Z0reP4F64A3tSeqZvlLKc4uHHFF0pRQXD6
rqM9XU4unxzabNkPFOkh2HJ19QTNsMpdFUzF0btAC47rC1r9CyhPM0daqNtDQ0Z6
Ln8XxhAPUsZuTyTmcNvhEdJA3zb9MNV/R998jz02cQdZ87KRbjBpuDfG/Co2i9e0
qxJMnKnh26M06JSHguwiU6eT5Qtr8iIVJbACgkPczYPRIEMyUfFnWSwiGQHc/Q4A
Fx3I14PeM1fBaSxLZEQ7185WDgd1+TFDhcNIyOgKQ2tOt9a62/b9n/yCq8wsU0TA
DCEL9tXbxQDKl4887vDLUvZ9O3qU2ROZoWYXs80MaiqtkbMqcy05nzX3URTL1isg
SLjCsK3HoLJ0zZeC0V+Y5aEhm8cRBeVGo4853XNKsFQ1Cwy89YMWJ14gsR6qZsS+
PWv5wOocQvr3LqgpnjCJRtiytAbuMlz1GbcXEX+ZKweuwxbQWfc0AICpea5bw9Cl
4Q75IcIGxSNKo5V428IkowfuTSEnkhLJEFTGzymjJUxRcvq0rxOFHIPBD7YB3zMg
OKKkcmeBymJIi/n486wVmzKIfKIqwzobvSWZ2Lv0qfq+w+vKYdypXZdUsMxG5wQ1
4SYpiN+ZpdHFF5zYOyLc6+OHsAfm4/4DzsFOL7cVdZiS1NisbDY9vk+ptmfy/0KK
6NnKUWx7MYjhKVRo0G4bgC2DLLdxLt43CkyhMw3V6que85vhAPbFa1mP/IpdMSxh
Vd2FvTBMLt/1KKIahhFgkDDPmwDZ4OHCjkhw5C26EGbvwjDiXjvNW+ZJG7SA7Byz
0QHv8rMACQ3U1hL4IJ1XN0T6Bwt3zGrRmsE/FK9IIKkjjQAWV5q+/dHVoiVdVLlc
Bqu3fhMdauLB8Ays6vDe1pzGRJRjt1c0iL/8Ua2jUTOEgUciUNSNJAXFQ5qJHi/Y
HgqgLLc34BFLu0SKJeDXx7cHz1PGjuAOwcrzCfOBkL85foLU3wuByeaxnX/mflWt
Qzfx+SA1jEp2oiEbu1gyjwRdyLvhvK/SOoF5F334TPGmLP5Xfa4Oynp3xcCNLJXr
aa6Q8bKtU9S1JABUuaH9VdUryqfVcHxiWQbPik2I5GQ3LQa3p/vPcPhGXOYvv3AY
gGrDn13bGASQOHJtyV/d5zWv+fmnliyAGqUo5BfEo/B6hTSBf/7SliWPY7VgZX/D
FfCK6UWU9MyzX+Ds2LSXzC/YBOvQTrcUtcOcCm3fiUInNnvuVhSWu2ZmzxhSve/6
KzA+GeDlKp0p76fibCdUwOE4Klg8MHQPl83zyJXve51PnryaNBouodhFlrdfLI4w
R0NPO5hh45AUmUOqohsh+b0M28J5li5a8CJCQwBUNrBioi1A+tSk/Nq50fvs7PP4
+tyMAUmcuX6xt2oFG1lBxv7Pryw1w5X+PubmE/PHUrWNqcVhcdx8TmiSULqsOIi4
6V7rFZNde4ANuCKn80e6ynXOWRRhuuj17nlXaAoyojNyxcXFAQ6cni4XyIL6KTn7
c3gdIrgTeD8xTT3nuyHr3jMzCT1w7CazANV8OqTmWVwcp6v01Gw6urgeKPMKsMq/
jLYovErNycorygoWNsYul+WwzDXfmo+lfi9Y8Jq2BxkZAtyuwsRWk/ni72fWRyOj
7sUmkPQxI7fcPf8sts9Yrc9aMM8fc+IZdgobnVun9R1xeYSD/enoPBUWLLddMgnH
tn77MeM1oCGO8OBNh2j329gmNDrcI/nhZZ1jUKHCKahOR7bikwfU3JoY0dp7/lWb
bH4LR77GYhUbKovN24UHhOUXt/Rz8lNFIe6kHaswzVOOc35GUgGhwgueNokzsPHH
RmQE3nOzHTHNJuxZpFdUF7sPdojT4YznxW+DAIYiFIfG1Xul56mLLHm1Npz3BNp9
rcEpt0QyJiIGu2BFpAOWqKUrHBlILMT+aRRYXUlyZeBJIXTgrMZVja0Vk+QTqAnb
8pxKVYEk8tnZ3NBm3QnILqen5DqL66nPKLQ9hGcrDVvH/jR34C9xluc3G59KhEWZ
iGrLE2wy2NACknnxc5H6BIQE5XaocQSzs5hRJdqObmBgNh+SoUErE5H/unI1wDqA
/T2E84HC/rGj8cs64uPm+JdOSQ66u5T93lh7dhGSYWOzJBSSEjlgMv1H5wocBspZ
KxTCsKK8JTMpC0L9wCF2xH71D0l02y5MKO/voL7DWePnjOyRV40LLsKs7LyqbSwO
g2pC5QpuYZeMW5pYJSD+B1/ClYoBlenMvA5cw3TgZztmji/nR2XMuNZ5U9eILM0l
h+accuMArcSNe4eOE1o4dwVp5+IjM4ozJ2RI/YjzL0nP5rp8Q9TcUWNxeKx3lLAP
4UC0Bc6e//bhO/cksEo1KCUF5/lThi2o+hsQvrfAb879yu2E20BHzCXvG/Yj2KDl
NHHlwsUwWtiiCEMPWR4NSKAcEIsXI5FkRKgIugsvKty9qZXUhjlNZp1vW5gqx2ka
6RaXPQhpvO7hMts9jiCJpQsE14w47j6+xIPofTunqCKY/wvCUkN4tatgXsOjVDR6
MZ0UDwB7sPIW7HcpBcmLVySanFTU31P+dYL59wxx8FvxpidPRA7vNth2wpHazHwq
m5zNE0VBYLG53pdFpEjoJxIIITLhMYy5DOYJi05W71DKKQuDGL5DOlLkQTG/wB7T
4wpcCmiTwM9VrEJRKG+4a88BLDxa4anM7ddCdJSSdI0HcrhTTvypPD3GcAR8xc/l
kgpFLLRvfDjc4t8/rXSptU6ZEQLVHdVMve2HFF3wLXxmPJYVfzoHVlrxW8xfcPDH
E4WNZF6EU8xe9DYEsq514JESaHKKxODFTCyS3YzFojTHWzC5VmRQ41pTx7EFCyAM
ud7O6hfvSfhcb+rVdbIIXJGQ1qO/7n+qK2IWR1lCIVxk8o6DWaX4wwHjtucSU2MF
p/pJz3UnDwcg5XDYL7b5mAfb/kYF5eK3yD6kSIpFkqMj1QK6fS3GIaNiiPTGi9vu
hsI431GchGRSOZimJGfR9NUNdy5Qbek9Y9qbUhzW506999jtv5EEj4jNoHuzazik
tPSee4uixFB72WTBilsVDKLtFManxqrM+PgIvvfIW8HLIggM2wkClcmRkW0PvEJE
WV8kEhBXIqVj6/BDX4niNrsUj2WCrAtxOUCEmJ3DKXz4xEu0D0bFT0B/BzV8pBtd
MBOViSO6hz6IqFDu76R6lU+33Fn4ZoL3kBVHb6GMK2MX534PvYBZMa4vJjLPZF+T
6rhHSbZtb4Y3gCVIwji1DFqs+EY0tKNVYlmt7FhbDr7em3p1SseTtaBaD1Gv22DG
1qOMT99gY2eWYZBx98Gb0xdi5e/llrz3S1gkMhFm9L8s1WbfzEiIdcU7vPa4waX5
pUDHncZx6MqgW7i8O6voGOX4aJcUj/dSbfvYslEI2L+aD82PK+ARj1nw5bWCjv9H
jmSn5IRRXOGZeURoUNEJNSg4+MmYyvalUrOPRAmzScJRYbgXnMZTGQKqogQ7B0Xx
r67GsxRZzbA2YnXnWpsAL1hXoXfNwaHqFPEQjlkxiLF6Xwx75JI2R29JgPewSYuU
Qa914jo+GBE7U3rXBr+xg/qcL476AYEROrJlFqm9+DLX7PD+lA18KlRrz4yRwksp
M7EXruFnwR6krextfgT7M0pRaXWL/9PfOOk/2Uf5kXHP0CDD9cU1RRC9NCmHY+7f
e11ych+gd4zaG7CIt36KGHtq91FiOgXGtKYhAvvwi5D7aVuc1fq4FH0jwNo3mF8e
JIOTxjRP7nmjCw6N1WbS/AvqJfUhNbBY8j00YA+ZhZwyyd5+R29E/RG7aYkVs0mZ
IMHjKf07dsx/Jr0AWwYRsFeT6yPcO8AX39z9HtRu2NXKfVCCOTECLK65QmePOsoP
fhzKFiWDzk7/U/LTjIRvjZZFx8ud8oaOShtI8ySN5qhJujQE5RyEQaoPtevSMq2K
D13K12HGdLXJPR58TzQKW1sQQO+pHsdorUCI23jM8L75sAWDU6cJrJwLqOoHYVUk
4ADQhAqglxiupbh5+RPvcenFcg0HPsYEv1JCwlYuYUa83UxXSNWyP68MYsdX90f5
hT67RwepKVmlaqRnZDyUDQoQVT1OgxjhjYYzTg8eQLdkIGjGkIGGZRG+LL/4+3tU
Ku0Z7xXzoCtpkHoDo9LkJxk43dZPL3EZ2ytKzubtdL4tOksflKsHTqY6MZJpOTfo
gV/E5Ri3Y4Ov4+e0ogB6d82CvshCm230GeJ+mn0djO6Vx0/l3Zkd5Wp1JZxku+ZB
Dhj0t5jkY+NBFfIegmfNAr1a8lB0SxA9MUPiz9Z/1BmQb/Axa01Yu/mFwzjDl47B
Zot/13GslReQG9+7IcoDmhrda3tr8a4twja/2BE/P57JF+y2oXvjWo9XOj9DIhYg
GLHz3tzdNarh0aM/m8zvAHvfDQRg0WtSFMp9SfdCZ+SMGYeO+plnxOe/VDuSHJqV
NSu+yh2LkYdz8YDi0spciXiUibarKP2ne5WGu9XmoDS0YsDdSmW1mpqoYgO8rIT/
suzK5aRlWNGGR2D5dzhwtgoKmfEOpL6kaePLRv8R8Q4ZD6LqntyE9hqKIdCiVuG9
V06ow3xqTfGRybTxnCgxQkq7qv2lArd2ZaAStByX7iC5vRYLyCdoB8159LRx816K
0bUq+BOJhMWo0LakFdeOS/VjNPLTykcCFxKk7qGESJGUBtKdz6XBs2YQK93Ki9T7
a5R1ghDxQh6CrT2RkS7B+tZcryArTzqhllydmFYc23Q3Y4W9NG+WnmfzrN2msrtn
1rGclfkrLU2aWsJfxWmAdS8umIlgh+R2mgCLQIIDho6UPTbxnJOA4pm204ameRzy
C3OTSkfpmjZAVBwwsK9nOQFS6hvYSYN9TnQKqBMokUNTCW5ueiohtRKfxZev+qSo
dvP1IxpA1N4uhdBCH910sg2RgN8g2v0tLbihpJjwp1Rb3jXzF9974fdfseXJHpmp
iGb89rHEphwfRJpUE5MN+xu8zKNxGynHSrX1+rST6dpnhUTgrxJPYZNljaJkhH1R
QhUIXFvd//i8hrZ4JUxjeyVfS7CEZ0YXAS4aZxj4+yL6l4+DiZEg9OWDdgwKjfsn
9lUkB8yt67lbrFoYbodgWbjXSSAR6xpfryd9icLOeaCPMkkdqNQXPOE5Rg+tKLTG
8boMqrmXB7YFXvYPxI+rQO2eNtLlpW/h+AgTzNhyW+au0huh1qW+JMuPXQ0NKatj
IiOAHdaxWwONZ2QLaDXJiEapOnoo7BizZ6b8U7p3u/SsGq8o2O7dAcd9tl2GLUEN
u7TegGfTMk9Gm+TrbXrqT/DgjkDKkQjGJ3T9HnUDkQL8mJZsbHWGwVeqyx3TI+x5
/unjv9XG9RjsI9UVLRIi2hcmVmEiVNeij1KlYHxMC9Dz3kzobDtiMp3I2ohiac7L
8rozYyH2jaMcvHEkMNxhf6DRw98aARRrHxB2BwbxlEopti2ajXbGnGEb8mCDFbiT
ynT+AdulvJriVZSMS4FNS9ozA1ftGVrbuS0zPEfe3U7vIcnSSLlqHgvuwxDCpZSv
7YKhq1gQKXxoW3QJXzuH+NXqtEz111fzsEcD/lLVvg0xs5sb8F1MoYj8kzNstYOc
1m6uZSWMSDwA5Vo63CxWZjeqaKHQjrWERFHxcmhHn7vpvusFQCTaSuZxxTkT5cEZ
bwAmPUCgj32ehe+jcC+Xybm06vIfmZfc3/5v1coPxaPXl98gdJRlyoA4MUbYyVY4
2RUiZhbb+M412zuDutoOtTo4J1nImmfb7xsTYBJrJPG9Q4kY2JfE1r0WkGBC/eX6
4jGfhcNUUxVy48vm6q51tVVNa5041La6ZZi+HfiGjilxuPGD7D+OQNazwETT1zTQ
KM1AAkz7ke8frVTaR9mxjs3pZWOX9DhsL0a7qL6TZ9WZQr70xbSpHc37k0m6VcuM
28Axg06zVIyADge5gEahetFeGgC3EgvMtXebUAKZjS6Fawnw8SSaf7Xi4z7fDnIO
nMIEOGVJq+sWJsA54CKa8oizCwho7t7n7h7V5h7gMREwRcMCqJ1olV9aUV6wvKDv
xgTyKz/y1235xPy1YSE5ApJDjKN3OvMvfmLU5uLebzTIx3Pdm6FaHoNcr86O5IWy
IxyOKLzwkuCRux6RzUvfI42rATv9yLtDWfl7da5VKvXAtFNRuW/kwjW6EnWCaEkC
jfInvElQMrtPBRjvMPgW3SUpIZV0Wr04HTEkcRMxTCLO9kR5tiTIapj2qbHfXeEM
uiZYfpo51efm1yKrkGfqt57wbWdsGzv5V4gbkoLXAYzhlkWOecazfBvAjFpToIj5
Q2soY54AfBlHNOzGTjQp24hSOTMQztYZicTPSXbKidozOV4PE0LtST3comJKYRXQ
tJAJlJOQHkX5yPdFLx/wJ8Mgba/fHruhii1Ww6r8uOmCw6Tpj8CzugDEYYO5+yk/
OWJFc7OCRpe4BMVa8b/K0A4ZQapC3kgyXykLOtlKf/dfrzKwAH2DADQIMSnFIm5n
VQu5KVTa+0sIDA2ch3o+VvgNHfRzgWwJ0//YPbGil7lR77qjTdC61oY6FZ2vInfg
ptmn7B6ybgaLPePSKeavsY+Yur//dlV0XlQw06LunY7AD1C1JnJlNt0NTUEN/Wg7
LvR028ZDuPAy0ACxQArEAIlMUXnB20zTrHwyvj6ouNbxuioiglr2IFlBPHLwZ5rc
mzp7JhFt8aaH1Is/5p2tZk2/4A9AGtYWUrx9r67bd488krYYna27BXK/raf6EeIr
I79mSlEKPpELyAF5A12F8vLNyz2/QAyB+O0/28RA6RZIZlRudacGXsIDZLPMjtMj
Xkw9jJngVv1nauT0lDhEOEcB/kbbUlWuC8ZIx/a5ASJX56iQkD0aKZZkCaxbAVMx
IXQs32hYhcI6GG4fQ4wn01UGVkVs+2rPEu3nLU0qUPIsosP2Tp/dvI0p+ekhAHrS
kgtppXJdjFBjYY9eKkeZ0qhbeFel9XWyqMX+c2KzokWGhPZeaF3R9Oo52jg220kO
W/nZqvtOV+VQ8SQQYtiX7DLt/QXAaVON2HPMPy6ulqgsl4w9M697zbQQS0y/8O3J
iUAI0nkx76t/CGMpf7EW/ECgPeAQFQQV30Yj2U8EcJt70BGr8gNkKvkOtyPXISVu
KnZO62ieK+fXRpnbq0kILKOHWKCYaqEOwcheBA5ccPzH0JxwDTJjXSP+2nnaXPQK
tEwLgRO1srTdG3GIemas17zQrjI/wcdsh28y3/+/nM47W1cmfHmmBF5OsvDligtx
hbTxQxzA7iZ+jV24FCw3jA0m2HZBs3esCV3L1SZqAJe9SAkcCjVwchUk1JKGG6Bq
cTSTIj8njtg2BWnFuO8Vq9VL1feJiWXNgxV6XEpARXehYIVZSUi++5HsHcU7J3G3
MyMN9s5bCntK230IyL/l3HxrUd7WGoKRHa/DUm1nQeX2NTTPbmhwj0IzZ8W/7mzN
/hfWUhVSybjNr7KJ1N5Gx5/bNuDleo2eBhICF9NMVQys0+AQUY9Cy9ZW4kf3k1h5
ua4FUd8l7KD1MfOLZEWeZYyKxFJipCezCK7vLW+EPO9hi2aSuPh63iwHV2D/vCeX
bHrd9Lt94c/+voa1MvcQo8HFILv1pUsm8xKRFH+Vl55l3tBIWOBR038wT0GorHiH
zzONcGmHtNk6SMRmz72YHr9aZNEusi3qLuY9v+snaL+6h3gwj4XGStAcf5AIhBB5
JY8iebLOfpQuc3DwJ8kfLKVNfR+khyuIVk3LC2Xqdue6YSgdTYkwdaB9lAMJRPVv
2+iWtMPzmn8oU8N8agalQPfL9Bo2ACdJkxWkK9GRrQWP6JWGsXsGH8aSvqKKpdxa
USjBTv9xaL9YSIhI/Jy2L0af5UlWHIFpeg5xbmyXS9IxmtZlsnACcPtnDRg73AzJ
TZKZV9Ln88nO7giQzSePbokNqMkneWsunwtNXNoaISKLOW23kRCNnk/xlH//tF0x
X6asDxTmOB2JKcrKw/OOi1u+BdIXyd4gIlU9LDtyxx5Wov2iOjjgiVdXjUVBKd6s
8iYbN0WA+a6WT7p0IDDU4MBqic/g8YjaD5MnzTcOcfHIiyNDEZERpjAVBRDpKwut
OYsl1I3dKW1TXeT8UEvfjqmPjjKHF94eWD3RbH9L1lxRi6lEQ8dlAkAGyLzZk0dD
owDv9fqUfqYeYU/iMoyEUGFVLlMZvSlPfzzEndVnL2nhKHyXDqlvaMpJlmRvDOYR
yswVS7zkuqQ8oOxzfzWjQbH+fzoUNvTXPM+zgQQHjkOS97pZsu1xoRmiaZXwFS3/
UyrAKErgw/rcMYHmVuEgkeycPgBWO76n+LMdYjKjW+LEhVYo8K6e5zpV/oiqHJ+z
61y/z9iFBOpYDvnjYWN5U3kNzYEuzpJgUElR/O9/bCXd2nRRKlLrsvNwjQaBXFue
JO6YMr6JJFL+04IDO/zxFLzzhxbNobTlM3tUq4c03znWQt2EUQxeVGzZeVcpnglZ
rWrRQAMgo/zlrhyeAl7ikQcwILeY/r2+QGw+ChqKcFWgj5iP0mkNHirCkJEzlZSq
S1OxEw+L/l97pIlpwHnHJdSQJv7CPuK5On7uTyOAN7lmb5zI5szxEst/6cDtSUg7
20QxopR7gr5VfYXqG7T54tNeZ9KashV+B766fTjBPb2ltHZBPxWbvf3vz0TOPUmc
F5VmRb/koE941zI1KQEiFCcXx0PyD9eGnEeEq+i1vKPGHI/X5hs0iBBOedVJnQjv
rUiaqLhZRUCPr/Fiq+EqX98TMbD4a1Mub2j/UH8AMfvNcuGKGMf75byyx7yRjjFE
hDWQBeSRXQcsVRxKQk/B4BT849HwGkenvrC6cMOiCb6bWE+iGsQ5CnUrkZQf4DGe
ZmfE4Rmw+llkC45frr2X/5Is5+yPVGw4E02nc3qeP8AhFwPEF7n3L/T5euxarv88
+Nz6z9KG5EMtz1eKjELau977aJFau4zJJLfIeR2nBMsWwu/ITVkbRO6vI04XhBqa
pH0ZHzjN1Ax9VX1Ufznx558WsOnFS2G3lq3+2WtoypJQqpMN2mbzm9pZYCBBxg9t
/7M1ro6r9fC3wa0EjQ4CufTE8WYs9oFc0V/x0V3Fqd8hZxxwYjM0orLmJQil+ZA8
1w7PmCtCM3dt2H4DFJwPT4J3X6v0/cQ+OsOtcmKZ/yO1moDvL6XSQlIOTsRBTnr9
bJFHuTSwdI2Du1AmZJs1FgiyuuGoOyxCNPBGyk+shnbE3HMxqBqxtSYZ1e0pKh9V
a4vrXuMaZ9MxJAnwdlvfhXYzQDMI0k9RYP7LricTM6+VcCnZk4Xv7NSY2hb+w7rL
mh3dXsouhIDEkSMwf1szDtldHlpxuAWa7u/y8r6+cG+hmP5mTFN+M+a2dVVPj/3b
FUhtffsB2e85DM1hYsoE4ANoj25arixLWMKcP5+vKfJjkLkA5R3uJeCHJ8miE1f+
YrsvwodiR7k6qlvHK6iKNODU2/HM6Tdr27hXXK5fL+r/3VKDHTGIuAJc6gR+30lK
xriAF/zdZlkGUIwkYvnAWR8htTEgPjnKJ9/jJhrNjOCr3PhTjZjtti39Qn776/7G
5Do8mHgF8XWhiIWCpcIFLrVF+mrKS4QIgFlsg2ZIDW+9XZ08oTU5qv90j2UBnBnP
iD4dXSglnFr45+McVSieKtQJigsABczx6psl+Fu0oYPGLpItx1sacSxLM3fDTTMk
Z0diGRXMNzL7u0leSF1sywGcgtNKQrNUi4yR8USRIFhlZ1T2QbVdtSTBXEAJRJMj
zBpmMajwQZB1rWPYnw1npGeDZ8LP40+6WaOUnodDi/9CKFn0DRh2NNTmyCXb/Trw
d1Yc8iZ7BSmt2Qk2RgjQA4KKRAbbdYNrELEwwZZ9/38zokGBvvtBq96zVb9PCZE1
kTmdMZjJFK8U0o4iLVJ/GbcWDP8QjGBO3XToX5KtG22E7SUxReKRXlp3xhkXxMW8
xC2FAl8Nu9tbsQ/4JMoKXw/rQ8I+7NbbY3pYLF1QEfKNze1fFnSe3ApVUNmbB/pc
KToLFGg1vhnJ/Onaxeb1dIDA5Ht153KsVOnXAWW6ruLCfsZOWcB+FTi0wpKY899c
uzBxM/TmRjJli+BVf2plxDGPBLChlbHqxj9h+smbW6RFGSs2fBk8CC8BvbDjp1GR
HPEJ6eFuzp87w9KH19d2uCUVrfvXbuat8wZ4n1tmzH0tRrkmOo1rDJpkpbDoyza0
xG5BPXCW8WqcwxxieCbn/FtRuckuL2DF043Mzsygp0o3m74N4TUnQdLSmIpxLn6p
1zLA83hcsfmBthXfOlYohY8G7XdIdPq1Gb4EjIK1o/QlZZ8LeDwkefOZO2sywdm/
6mYcKHfE/g7vWjr0zPjLXf/W/eW8RxX3m+r1ULhKyM4CVJnk4KPkNyF3jkb75v+g
yL7PutY9LPoa8K2bXY85uMicIpk21KGDOq/iiAMcn7N2UV+sRnieNzDVlOKF0gQN
4stDyMju8HcA18Gwio8pcCugJOxaZQmULz3G3u5VTt4Q8e8LcnF8CFS02QmvfVRc
QO7PW75e/zEHzchjGQJy4qTDGx4gQc4k4mfzJ5lDpsjgF4HjW19nhwMr5oz/qiEe
mpbF7389kD7VfvXTOMnHEeAgnpAbCZ96XQzysQ1FbEXdJSH6eZQ0VXyC13w+fmhd
2WE26/DDmTTCfgN8vwXk9KujyuAfw/qSps9cAFOHv9ce2w2LTKHXQ34J0ovDER/7
XwtsOlcfLQZe1wl16urI+wX5L6F6Ks9Kjz3dExIm1iByQsmCh8How5p8Zx+HbTrA
9eNY1cnzZdY8wCtXBF4DYKorzk1mFaJkqCrd6Umt/eWEtYjXywjzVzovjX86bU3a
bZDRiFTAqNQBqkP6sfG1Dd9Z7e52pZnyHks/PQgG+tH+YEbr6n/HHIjyNjf2Z4Fn
ogbTjQ5vDRFaBj/Ehd1TeR2FEOlOQfF1914aSyFYN0zheh5/MIDqsSEdYnSZ00Io
SlEh75pKwPQWU5Y/5l1V3Pj00mdxzE1raQqARwmJv+b6+un/wEz226sB+l7Gu56i
0RC1Bsy6XM3rxBJhvfTCAtGOyjslyRGn6CnlsbfZlDbN7VVr+nGBDHx3N5qbDXbw
8lOvyhlha7R6po8PZwMmcg5/Or/PXOUazg/FKfYcRznMVrorXneWnj7cWwgewnP5
poWWyrPLVNgwmn2LHiL5Ta4R6XeodNFSG+RgmiZ4av/7G/MVPFTMvYiE+UyB94yu
NQp4U4Rb1iFj3SzEbdv8Ys+xEEq+q0pYa/xGVr+I51RWSxZi0QiJBL3zbZsHXsYP
dsfCoRLqWMrFwixCzkZdikAruDExyfFEkJgx+ySJ1p8f0AjUkCFXNqosVwhjKp9B
d6PPadrMgJrdnPZ31ietq1fsGYrco1qeIfereyrLwp/d8VIDl7yx4rqeDDYp+PZD
2fSgVRi/BdwL1zTSZsvGfA5fbb4BHkGWbkjaO+GUeVqNLYx2Mt80HEzMaQanrfT4
K1rrbdJRKgZw+FmuG+dKTf7T9mMeh53Y/ZKbHetaHB4mXRuaoGIVXf8A7M3D98Pw
cAuxN2iNRqrwijhqMvnQXb1kJuz8EBoJNyrfdIAaETf1+tCTvhvo1a6qSl3xyHrj
IAcISmP3ilZN6xz/m8r6a6ok6C1o6yLETdynArnfpqpWKFOIIKlB3yJkRQq/XMSg
zxQozwp6KJCJIySpINrLY8iiYhSPuOYHnChSceOgPycbE31tvamUUSpYxEg61Nup
JJqmm17Sl4/uUehuPrx96c8sdKFHt31E29NCVWs6wh1Lf6jdgRrWh1kPINCHedC4
uCj/PmrstBOcSOEVO1p2jevHwmYcP6GkJ07QRLB+7v0U6RftbNvoccyAMcnmPo/t
rhBn7EOovYbXBUInmsHDzt/uwwLmDMDXFpnh4cjlz5qkUI9D3L+v+IcZNAr3ro21
E5c8pKxnQmJI+T2aFeoT68JLo9d2Sd6lYpg3Tuk+hul7CptNicfeGHN+bfQY+QEM
q46kR6GUCrd3RrRSyOM62abNKW3Kag27CqtvkKDntQH8T3h/52nQeoBJ41Tvy9Hw
Qmc9D0UnY2i8T4hnBOn60FXqTkzJR3JlNkADN0P/yDAyXYEJdBTn1YSSkC++u4K0
8+rIHfrEp9C2BZjYuv7Bd11x9VAquKE2dZCOElqty/V2xZK9FwTNiQT9KNYzt9OS
k9gJ0a2eGXkIsfnHlvAUR+D4iC+7BZFCr/j4cLzwmfFoj7NGImFax/y7Rqo8eWhY
IhmWv6SU5DznUb7n53tpvG1wMncL01dwdsOmk9qk1hcMZYjRTPXr45bXLwFhOaIt
uS75EMLIanCcoqTbVi0hFTZQJR9KdD5kS/jNkFY0NO/fWWpROk/UK6JfUXSxRnkA
6byEAfAqRZIlsSWtjBPHSomhblcQ6Q1wbI/VKkHKom2laPf1x+aPoXjPhRFgV/fV
6oWkkzzzImIIDslJ2wSNLZKDeqSwV3zKxq9EVO38HdmoKeEXjYBCMRO4V1oPLD2t
hVjRd68PitNc934YO7RY+jQs2kyOHeq6C9Qf1vEYCna7FE0Kw9KwguV5C3kLiXj7
FTSFj66gdKKRrhxF9uMGShNF6el+DVjo4fiE+lXMMWsj0PK0ewhgJsp8eDnj4cGp
viuX5/RTVt0og9ANUNE0C4TrGeuqukpJCG0o1AIeg0sEzZbFqh9/D5lw3OxprRwr
NedJr7quU6VYWN5RXQRbAwv5e+oihptQw1CZGEhGl9tVPDKW466TN3GNp3+s91lo
3sjkN7D7+Wb68TMnY/C2Ra5Qi8KXziaHlcCjzd8K0ytXzL0GcHeipnxpl2Q0Wh+F
vdMlpN8V6tOmDr7SVNkR/N2IyWT30byaD2OFkCLCHONnQGPALtmlPdDj0dsj2Bli
FD3PbuGhbDZVDdTu9S0SS65ZsCO+7JRWdpo0PVfHj06m53qCXMgpL6olRA0Bk5nR
YXrNSWsCwKXM+VC27b7nLVfd/QlCfqcq/j3YusSAvTCNLL9dSPEatAsxe3cvi0Dh
xBxMrbqQFBrkxzQHOJeO1wyH8pn0d12xBWruDFCb7FcZhbzyB/TAx+mWGxYE5c74
oAybUoPJYhlkN8xlMyFbARAt99M88WMqW6QN2fe3AxTn0seNPwDbbFqV0EmYbUiF
lAR4fzzztaCpFPNBQiLw+i+FYAXiVxdwWneaxRKiiM+f4B9jCetYeSC2XinApJab
7nm2YSwmSq/pvhsO/5vgwkyZEAYyWRgfBrtg2OhKtGjyi1jQmcBblHHzUzi2hXNy
tJYrD1IhCqQVRB+rYojGOrCd33GZd3Y95ulvlyg/KGSHl0hYbCqJGubDeQmbg//o
qY0di7myUfPjA49RUDmBcWT21RE++yLPgrWBcWZXvsoYNE0woNW/BAnV2mIFTy1B
al/x6sg65mwAKSVu6PjNWAOdsghorYG66nLffajUqfXVBwYylnWCblzxNwDv/TmR
EmnsRfP4GkfLuqa8FCPC4QTfiPiMEdmgJx3F6qEvZeNhcFdSu6eVU4mgKuCoa61p
wdtNQOx2ELiLPEtUYyyjU1kgBE5RKf54crrg+N2QzGNmCWB+97QOZQ/fClhpFxzU
hsz1WcVggKVy212zBp/8Rwu44p4S9ORDzIePSPgin0Z8k6eN/tSPovlglGMAF3p/
PCBfVe/O9xCCWAF2aCdQowShMRUJKQHuTQ4cy/yca0B+ebAjHyJT/ALuBlQbpVaY
YWS8B16aMZjDfPtCMaqH6S5oM8U363z/aTLaL/QAVw10WkbFWQYdwi0qT9yQgDaK
j0QMx0dJuPiUoM4blsAaiheqz2KA+kdrpa2+ERYpOCIdlT81P7QoHujQTv08S3X7
Kgw0NNWvKCF3yj85bIlH9tDNxJFBJX6ryJhJQEIETAzJprB4e8/9q+NlykR4lwwU
KhlVKCFJULM/ChQPiGuz9muDCzCaNabS9odGJKAid063TSdx5P6S9EJJI5Ka53Wt
jVAituIRWc/brC8aoB3kb8JEx43+i7QXcBu317CPyfsuRnqcE5YNA9b9E6yufzXh
e38NcY2seFgws1NkWWs3oIWhb++gMENNOaA447EVQOW4HBowcYPb5Pjf9r32+xEJ
ZjPtHff5oKENNBbdB2nNzKqHcSrltJ+Pji/pYSQjx9sY/hilKFmSkk2AOi+lr4AU
JFaZQYTmVFVZskf83KnwJ9VaAu8grboeIr5wrzNTrzQzYsCLbleLafwl3dFflzR0
YmgPM3oBX+7TjpzMseYiZmDrlm5ezohgQcyfaLldgruWKwC4qOCMirBoWDBC8dti
2Td0DKwknLWtxPkENgP0snqn01VxRk4gbyR0Nz5OerB/Dsb9iIZXq5iAvrQcIPMI
IY/MGN1RlSwa0a2fJdvfBTcOgILTmLgFqilYiVShL6M64SciLovS0ylam6DH0Xjs
BfNAIle9sOClGTi/Tp8LEyRzpXyHOPiXPUQA+gMVZFg4OeryDz1klAU6ZeWsfX+e
c6RIcLateTxmCfmA7Ducx8NuEtzODDQdEOUWn0g+CR2LDTfJwg/5WiNY4SveLZJN
Efx5HLj0DwX8coJzVSfFWGSHSXSnokhDfIztGrQYPvKW1v0XlaekSLmhq45WQBhZ
2qfa2rlxO3DRmgzkk9Ak/rpX9Q+vSWXVyJI2HGJYRJI8w18/eEdd/MCREaAZXkgF
jlebT0jUcOJCXGcz6EmMG+EHPnDOQKauMXBmALph7anUpoP8I8VwzfT5KeDErkkV
plN3zmTgRX51Guxs+NxX+RVEPhM+kpKsMGo2IRj8+wn3jpOCkEgaEDJWFyoiKbkY
8HpYtlNa2s173u7aIouyAeubDoBApc2kPY6TK042Km8gol3+C6I88vI+cGrDzBHj
Fg2WkPiyLdbuapcmeUUhBGL/bBJG5bzgXqFMcNXfEYS1hy8sa4NW1RtTLOW+zier
G3whWpH0kDAr9qKHKWHVqBqA8GdgF7byjjDSzuS0RDB8hNv3b/zppG3LY7mJcjzt
v2peonZGD9cfJesgrzD7dsWIA1R0mEfhFRnCrO/p3XPixocyTZc38hfXAHvITj2G
t92srzbzx7k2LhRcepSpBrkQGAGu8DD5ffjI2HQgovZj3Q5v7OyMq9i5xzaZzo4J
phME/5E7a+ifPydROyDpxf88Kl4zwn+iZYo12s/Ti6VH7shw86W8VfKjlVsxBcv4
Qil/7icZVgxJzhzSQjj1bEU96lb/hKMQ1QFMviKQfVYqAikE4eX0K/fXEkfJrymD
jUgH+RwEcyW0jzSU66sgSxEOH/BzNBK2cN6+qf+T6dCzLg2jw+eJD7Rmsw6Z66xE
8E95J40WQvH6Bpfnhx1BRCm9em9rr/PB3RYsB44RIUwKsF0P4QlLtPY+CpdTAP7u
6IeKXE9EJzOfHb7A77yDkZDL/5vvWZi+c+ueB8BDagb9xLbgl7Fh0/bhiG7fWEO0
tfhWmoaySdxCYIDyBKxJHEVWE2M3WbKDfLcvawgNa6saG6c9Ew2ZrvaS+uB37xi6
zO14q1mvp26YQDsJTaWf61KIf/5Yf+UvcjPmHKBJBHrciY4NhTmTjT7Rah0uaKJC
rRgXju+Qtkplk+XjZDXvTc4orO0Oe/TuQu4acFK9G1L2qeAjZRbBrHBBJrwsDcgB
zx79Zr8WmD6x2NL2PkcqEAECaqCYP9lG3zGLiQ+0JsO076qzKAFjAz7/pffr07FY
NCQQQxO1HQm+Vlf0i7z/1LSOY2xNU7TiElu8ImOupCVIdC9pRSzFe+CmkKobr3gm
fTm1Jc7p4GIYeVoxXCCaCQdes+lDOGIALOOxQPPPf5MKiZiUPf/Vwm97Rvalm8Ju
BQUvwR7GJF2RqmzF80jNL5+UGx04+v8Elc5qzTFJE7DilH33pjKJ8Chb29PknlNU
NqqN/rpXijPw9P8fkl+Ohehn1yyrlORwHIeIsd0GP3yG9dv4GX+vWNqahtHJQzeY
3jCvu4JD2gTC2GgOmXP/Fc0etnaWYqlPkyHPV6kw6FyjwCI3sVblX5A14kMr6l6n
0NVxj8sNx5uJflOu5SUzfgBUDCjMqcvHOv3he4A82EShcS/3z3V4LLN3aOYg8t1c
3EsB629WKQZlVKrKRugYkEZmh8WrPIAfzP5Bc2neBcq4CbuabFC00Rb8nLhK5/R4
McRLujlLK4MIne4M7iwuxkL8R8Bui04OLgUIOYV117hfnjCe+upSQ8kNE4ZMDR1t
yXcBmpZpHhJdDhb5jvAhAZp5XQIddChU5YifJRq/H12kFwbYm3ovml3UtHP0o2hU
hMgxu9HixedAah2dwFKJR0MJYSCLtEYpv8RY3g1YBypGHXygVYCBhQ8Ft3VocZa0
W7UG5S/Oy45wsMG6Twp2F3rzcu1k/1TJuk4ZV9GkwQFoAqa2O9pqI/XRvxIaxZ1Q
prX30Zx0z7BO289ZKole/K0tyEtuK5Yyf7ThHqKgWD5adrdc0ICn3+9xPkkw9FnZ
5IF1oWcZsL+Mu8V6ejZ/Bhw4pF/MAgm0aLK1cSg7mqw6ibNiXbsimtXd5KDpQbn/
9/r9/lU1AfSg6M+eo4Y+5LTOs0aC5mUpEqzYb+j76dpPNXFTr/v7qDz8XtdEtH+U
G1SONKLdPc3tP6sXH/7pr9BPSDAfpX95pQLw0og1V29HDjYGH3sxzGylSqwM5kQF
MFMoHSlunIQgbIrJeQX4QeM9XUuODq4Qn7O5UcnS9HtbzeHBlB1mbMLK0bLQvKkY
ex1WE6+4aEgXvz2pQFqBmGIHfHHBWuCU0274sGB9YHspYXcNsX7SLoreCfXHiAiG
RTI/hxB2z8KROAizn4SgubTyGL/yUUtmmXE2zgo+bisowaDkgEzJfgQsqXwr8hU/
chnLQMIJqpVEcuDw7//g16BmulzLTWtX3mkpxPJkV7S+kVjtoH4bff74OsQyrhEU
Ug2q2sxLQOht9cTy3ZtuTEndPUdD78dz5XDIQWMuNTu1qS0+/va2WJ9kTu+3D+5J
7EVF0o4VtdCw1oK3/HS+IgIcmzfv3E+tNeDwP+jO6Ywl/CHgHC3Of1u+ByZCIGzJ
COOEICDC/DltqkX2fRvSm/wHdn6L8lwL0rHjtR0OyzfVtrwdMV050bkd2tSxlhLZ
49yZZtYnX3mhxpXQjM4bVVq7d/ErEYGntmVecd8IJpMXWDcTnF+Pxze6aSV+Bmy7
yHqqS6S+P65Rt6M/h/H3d8J/1nbBKSp0I0mWm1eVfGqSrkyCh6Lb+rEOFDphxbfX
l/fUY1Ie7PjHAZPmjNBU+DtzkjOKDLVf00kvQCLndKnyrPSKFFY09mdSOJCFq5Im
f2C5lInK8tiRp/Ta4kYTEAPV4a+EXplbOlkEyQWpe7p2LNipW/u7Zht878P+Zpps
xPAp+p+4GPIET0zg+0pX33x2bFt6tUSWVHR2mFn6IkTf/tRnEKOfQTz0M0gSvOHi
Ufbic85BqYC7Ne99RxD8usF3gccb6L73RbdSayHck0K/D4cDAKEPfLWI98afzeKV
ejwya6r8LycCbNq6WjU9Q65VkAwQymE3xznGeiFTQ7dOBI89FtTyO/lKc93aJ9Q3
33nNDU4wwNN1EVBG5axaahuOw4D2OaUCT0l9q4C31bYN6uMYEkDFqpAMI2fvwuYQ
oRZG8DUcrHhQrFTBlHTKfGpj/MorakoLhC3Z7nBUsAzY30hXahSHKFaA4ReJdpRB
xItuOvLsmJDYOkLm3OhnRq3sEIPNrmufBFW8baYnYmTCdcqByZ+Bj0KvIUszpSAP
DVN5zh5feXewuTvLH4PFcEIF0otQLGQMcXXyKxBatb1oEvRqhV7c7pnmH/r/fqDJ
mewHDGafAlGf8Wsz8UaPuGrpqYqyozkyNlwyuGuQVBoPfQvEk9YJBajAFtSn++Mv
/G2kDJR/nclDtmAr0rQtifENWv0H3M+y8mvdKMi3wkDlRMC+YHY0fmyUZyipOvsM
u0ACKV9WYYd6ViTa7sNb7IcK2kUjRFQkQT1NZ3SBt0nDsFahya8RjQwnWlA50OUE
CCdf/ccwuwZCVX1SZrt+MKZ7n+RktLGrwnK9CFNMJpaV883iU3/1cNFVGCwkCz99
5UH9sj6ExrdSS7BXLmHcdc4wOCl9++xfGcaaXkkvctODSnQQgwuFlIQn84MWPTOK
uHd513t4hUqbmY12WXTrDCTdu/fS0U6qZ+rERNHc+SnaimkOef69T63PCR8waCum
wDSUQUL9blTE4vylFZZJ10ICIdsJi9LaGqyPWPdYRE/GgXQJBMbBRrdWEeOH6HGp
/kr9UXPXNyEhj+Rjy8Cha0heaVETRigvn/HR0HmLpJS5lzVsU5RI4SGavazRXduP
LXUNdczipnKCz7kM9ycDMW5WRfgTNc0+OwlHXrrS+2QH8chd4ALyf+Ols5WXKU1O
lv71dq3IwO7+A6iGke7/PrsapDQW2qTL+PhoB7BUZgiXJNigOK4bfsANR5WRnYk/
qBqSWR2U6KYnWMaOEAIVe2w1rND+wPYma+GKUgwJYoFyju79tjQYSra5OpCE7R4H
Np23b1oP6zFiwZz98BoV5iFygr2Pfk4ZQqYeVl+ztQyIyJfv/HA2oxOfzQqjx40s
8+Cg6NRXfBSdzGbzyAmf7HwdDNiXVRmBRhLBwsfGa1+Ef9BSDKy0j5ybYoBHUcWi
/b2I+jK0QUQ9J47yrfId1Ol4w5+QSLT+Kaq2Pe9lBrTCVorTvCP45uIppiX3qw+J
RhOiZHn9ceq6ZyaEb6OkazvVmHvUVVgQ62R32maa4XzKQFL5xxaDHuJ4QqOdxyGj
H/Dd7w/Okw2TwAUmaNzmKVtNTbjTKj1V9vs29EVZw3Jvn53u8vQkdWGlM2HE6Xk0
qDb+RADdlPR7MMA3TikmQuOfPRTj3ivav2qhn6rgjoNZpB0M1AR2PLb3d9u2giEq
EL6HPSSPF91e/uIZMVlQborYviwKvM+ei4JWZsxFAVprD2odesiV7cskf49x+8sL
feDhLNaXqQPFTTpXrwEQNXyeESbcM306YH7NPt/gYhyOlKBO28gfBYFgaYjs7D1Q
Cyhko+lecwxu1mRkidU3pKfvpHrgoyYExFgYKAQlAP0XZXFXOvtFSk8RYb+nTOe7
dcwasV2mUHHcPNJ+NFG2yEId+pXrenPF5RcXfKM9LEtmk6IvwiGXlxjD3yhMngWd
DZZP0OyK1cWRmGYl0jpgz0/K+SuvQzhAmu0q9YHXarooEk8AMi7azZgLDTUSEQa3
6J4RKgtom28JA68Gl7DgzhNy18yA004c90Nd5mdIhtNIl4kz4hk6WiVQRrT6YtPB
yYX2zE0ekzOETuqOMv93Xu9mnoh9wYg0wEtUyAeCI4J1JmKqqI/Co+Qu3MNYR/gd
0rCRqmgF4TOJF3/CdxUw5BbJoN28V9sj7oGu0UOeTC0XjGRdeTQRf1j5lYAM/BHY
Qi3BZy0FwIaOp2qBar5PZwLvlVIwZ7MnhFSK4ViL/SbDmwkRFCbkPN7JPEdbvxYQ
M+DfXOPEeDWS+/KCsVatcHrAU+vwigEMyDeamn+fFGxAg0eCHMWzoGwKS1jqF9Qy
eq3UjmLVAtBFyDGT0qCUVzMSvlPs82k89V71hN/l0owQXZ6QMg2aVgt2QsMbZWVA
z/+n3/j+nqLlt6b5RxJkHysvV+94hPdG8IN0NBFxDC/zCiLj+VvIPVBucf1pw3yi
oyodz4O+fJDuVZIygYQb4egl+reVwlJFXjnQUdRhUP+kFELTwJx6Q/8OmiGdBFrQ
4NfX5uht4cxwX4JvzOtDOKPHwEpcggq0GUgHJ1EyR5qVKgqXpXf7xJLlYs7QlJKI
P69WJJsT0872d5nKehBc6AyEvZyRp+tiZMh1mYqV+Uu+ts8JMFFnSlaUPL6E1NPq
cO3OYDPRjqOewT5pug8uFHNLlmvLqw2FlW1vt4r/mF4oRsf62iKn2SuhYX2Qv5wy
pz7XZhatAILKeEv3cLvCUAz+y82tqR0sfWxpZT0zNXPq4rQ17stsAk1b6BmbR71+
Fu5xnDcvx2kglCqIqyuLdbmnpao91IH2vVZkkvjJsjRL47654rQL5ttKQWZhj3As
gb5Dyq1u5TT07onkfEPrCg7sV4qgmy9AV86US3YtE6z6BO9+MB2+CSvqNgZqnie2
5e+quF7o33XdDdmJsUXFQjGzuZxEOg6GWSCMQtfRZbmsdwT2tqZSd5+2cJHNG6kl
kCeDXBTbeWip1epF8FF+/6vNWeRtY7DHqnnJoF7LSVCTzlLeXvW1pP4oSfGhWecn
hyfHW0uiC38uS6IBqCu4O/V9CWla4rVEJY4I2Ki9DBujh0ASONpEZfCfyCt27fVr
lwu7mh7jQmk6W5FgCy0i2BloaJI5gWPbC5qUmccpe82zC/Gfh7ZFxXvnARq7NW2V
QtdJ4xC4i7EckPExY7xsibf6wPOtkLrxmQew/XZNjUEWcKmNQfJ+NTfL25tnDthR
JBbEKXxoF4WzjX+TYfIh0E583KMGwCq0v64koZJ4tE6SzRWbH26e1TgIuB/355Vu
LRMP7MrMmd6BakzQAS5tQ0gW/BQVdmfCqT4Y9PwTFE2OOhehMJpw57iiSxJKXY8J
0ezPUPRnQSyhJY8pBq/kvQnO9lxREJ6H4rj15oszMZmlVqdD8+VKg7a4Obiw/b6B
vtvUHrMXhi/2/TSbSRhTVM5vHPfAG+U4KwzX6/0vx35r/tCkLrvJSzrd6WULbQBu
QPHQXd7eV9uk5MSA73NdbR6FINbgbpJtZp/vyDAG4tzUUYjGZxEL+8iJ+9bD/I+2
h6Yd3W/+lD/icv39yEIF7chhjwGmbZCwn3PLlP6txRzdRL41EDTyh66UUQM/+FOP
As9gqP7NitwCRPd3ub+aSklOtUjNJWjMd1iRxQrJ7mGUoN5nTW1++PK1FqiidwUn
Z1nc8pnAcoUHpy9m7FcDICu9TRjauRPEGqb9XrWNPWyyf17KUg0qhN0E/L8JyZKY
r7z4GVdEJaQfxRXs6mkfxKUAfL3dpS3PE0Mg+5JO9opwImgud4C4ERDGebrHo3VF
PvShzmx6aP1njJtwcOwwJpooY7DSfC/TBviazMqYiboMdehiEnsgx/3lgyl7fifk
AMPhYWhkZlfULhVSOEymmStkx90OX9PK55t0V75pDBJ5EIqHuUvmpVdV5m+weJ7R
uBbTFDw3/e9ll/b4E0bXpeIiMXgh8Pym69lTDrjfSPGT1BGhpxeHUmJkLQzjnvhZ
2g8SmKVSSWbZkmuKLEJYgrTaEoaZ89ydGC89LF3UH1D2/0apiQ9lO/JFpQmAm+AJ
jkjf+WAsoO5tVjFrQBFRJZJiHxk8rJjvfkh20wMyQd+1E+gXg51YIAXLv2y+sqYV
Amd9JI+prxcHhfhtczsViJc8cH6xWyQTddv9HdGtJxUrEFhaTkevaDBpkhzMFp8M
V9tsFowi4dWL+66bZf6HO/C7h604Bht67t+3gnWLo6bl6+NjnIdXAWIhq6x0oTT5
iAYCI49JyK2Y6h9wRL8RHQMvVOYMEbO8an9oT5wDrTphnMSFp20jCQCaSwR8Ngmf
cwPaB6CPOtlnBhGWH/ax5bCtOmuvalO3p1TXfng4ntTCTD8LaPdNFdDEieNSlrO8
IvEH+L3qM5RqtheznODO3TJFcYbr/syRyGEf4YZyC2OWZc732pVbc+g6qEvDxYf+
5w/9vtLmNC5R+nKoT0ipFopKHFAZ69UPrHhbmh5dhoUNsiRGzajHkbot0xjL++VA
aW43dQ+xKUKSKg7ZEhz5d8H2mATmvKHkDroofTrCc7/jmpMJsJ0LPMXX3UWcUgiN
hLO9cNxKws0bFD5tO+K/jerW6ucmKnveiFtUsF66/Pq9fRlGnbGu3MY3KbdQaqHE
Z/+dbVW+m9Nkh+uq86k4fLFOCBGTmtTSh7e56BuUUP/JwSZz4E6brXCIVzPKUpMG
+2BwNP79/xonTVnRYNZ0KEn6q5IkeZHJP2xQDMgwSF/9XCrglU7puScqEm5Xw5HZ
geIoRm9w2UYBac8d5D3DXQCMjPhcttex/Z4ofM90CNrrtWbQjW19M10p0fFC7VKr
FR6qxkXngOnzwk2xxW5vCQpxDBDZvCp65NxZkS4FowGag8XJ7YB2a1iuoAABDBhp
BoqRo17yfj6Ri3nAyKDy0W3mKkeTZey3YwREVdundRarHyj+0WvK+ZdF0TBP1B3Y
y0SKup6YXiabYu2gWf04dOy6jhQZhEsOwUb9Ei9PNOyHHkFxuHTiC71OAzDw/bXp
yI1OAbnpknomfWK7iYmnCNniaW+InlEh0SvERv9VZ2l7CMkjciJNgwnTubNTL4/h
qWGiENGhCnK+8+QU7GpLeT8EWWr5iSqNDhZn9xj0eeTMJZVnVZEtgsfuuHwQFr0B
so889JK4XDiEpUI7vSz+BZEwV0LEEhqFP52NEwzNvHYpVLei6f8qFUzRgs23u5RV
evJX8jJLLS4JdaLna/sK+RMtqe7B0p6lrZpc3DrYIn4WiF7gywvYPj8YWjFFqQdp
5XS7ioIb9qAldOV0rT7jReqNooubYletpNTxXzaUKqsMb2jAvzFqyB2uNMW2nCSt
UfSB8XEm3JkEFMgz7YD/EOgPhB9zWLlghz34/tmGFYSfj5HpE2WJgTdx1xpRAjDa
dNvfT672SixCYdqLFI09G+fPJV3vV3lW7ic0hB0+ucSzmmKYaGppxXzc6ndPXKd9
hW75elED20K1vzparQCV6A551syoF05YSK1sOUr1T8BvN5EZG61efKR56r00mdtP
cUiNNR/jAq9/KqsmKPWDIHMHTdtnpWj8rBz4jjB+/ikGv6cBYPudnjIa7EEdaV7t
jM7oBex4HRRjTlVanCMwnukfi4CJrvrn9XmZ8wVOps8gI9m0t0a+v0dEhU1kyKPb
YXcWx5ov73k0QhhHdWAQJMpNJ8bdAmnkOpjCOzw3bNlQ+gcgs7NBa7hv/nUR+CAe
WtesN43PICfzzDO9OyQ4x8e0zeR2zE+dcVWUeaP4dF+mpEwP+IsNWSLWPycuOiws
X/TtI6/mroKmTWM1SHiWh5QkH2QRWMFDOXpqLWOdW1oH7lQ4Odvi9nTUblx7Hn0I
zeJ821Mr8dyvhpBCMno4/v+jebgNdVEjnRB03xjinIcMPrOGbUK71WFrlPESEMk8
lSrkiQNstcb5B++0wxaIzGY7MAjy69Mre/Z6ciAWwRlc/K2c7yK3sb9IbfLlTGL4
oj3bX3JjlD+g9OOHSo2k8R7dvzlTnOuMvMf6dyDUdg/V7H4EXqcjDREhWcz7qMJz
1ellk7tIaoaIIRkuoepHpE/4P7oxYGAdVUOVFeRJmj6vVRZwSNcXhrlTeAeawfWP
DJRAwF0yGOiXeEhSwoXCpuOIp6xB7JT+3W8FnBWImDaZAzn2YzuF8+pT8anclPpv
hmLImwcPq7sRjfsmk5+rgQg8QpXX7VoEGQy70Y1NvqpwgVytfvM9LhCLAl1MFmOg
KmvdT/O6qiOE0J/L1bM+TCiX1YZJ1AZ6jB0J2NEmLpNVrg/StNz/fmVpY3Vx69RK
r9ExQ4QiV+BADBAJOEyfQ2FmfCl4JsOba+3Zq/MNhMOHRvv2s7T0+EV3fhrim8c2
3p3KZXIfTh5G8ER8aQlPB0H8K8fkWvd3oiJRQG9w0xLWDPyG2sZOpSMCN6ExYpZe
qv667/ZH3IYrmP9P+w89WOQ35bdwXAfGfXKZiCNrjphBW3EUKTs0QkWq3y8Pvx96
RUxH/aejM1l+8CgQEyXjw6wNtGpflCODds7OpLROxTKwT8QFRLlbd0tNnwcYUUhy
Jb31PUUh0f7kPRj8nVewNIMrZGOsm0nNKOfe3Uj9MH1nQFq9046mdG2R3c/3GkRO
BQdeXHtfofgazmxMpdLJsJxtIE/34Rtc2xIrNK7ttdlLjn812R+yFOG4nREVV51O
KRvko5t2THug5CXw4J8Wv5f/q/qyiLCXygNgS4+Y6YGhDfvfVMDvE94JoGas9AL6
kiBULm02Z7H5/oL192sIqZTwn3RuQDm0RlZyZRLCB+muFtFj9PTWtS4JlzI4DEFg
6IG1n/5KHVCF0HiisMa5EA8L7rvCGipny83jR4sfYubRv2jxyurxCX5+4I9e+XIE
gg9AWyyzCXtXlSNNJiSpyKYjMNLAP33O3oAwuZkI8e0p/UYZf2fYn3RhRhwhsI0W
1IquiuPX8KtchBr+3ReAlraVAkuJ81MHdsWfFJfqo01cQPghV7ifBxOlxV0iMs2g
f21H+Bo53cCQ6dpCiNviFgmS8nHgu2y858F2fxOdjAbYOozBzCekHS3m/2uqIzA8
UqSdGG/JXcDvZOdH2BdgNm1tt4h/Una/xXTFQqvyH5qYvFM8/6cKnjcf4I+C62I4
/AUD9O+tsBeZVvy1lnuShHj93qsGk5Xzh2+9ejdkjM07lPAIvLylk6lxmE9a0J+E
uMvXeJ/rzZDnb6BJajAiUXYsQo0uAtnaK7Lv6xZEXLErM0JkTtx4YbdPZJ5FVrxk
h8+266QXRimP3VbR6VsBInbzNIvYBlYYH9L7WV3l66uXjY3Y5VobolY0XWfA5WV1
ExSQKD1kfLbIILlJ49VIE5cPyPru7hPoSv3+EMBviCQvBl7C7+1+ckhJ6joVI7T2
NYGk9WYmKEV7P+nqootgvx9AsK+EiWhqes+K7ZPuf34il7YWNtujaGcUz3RwGc8d
TNxb3w4vsXmkDvwc4wjovFVSi19fT6PoAFKZs6zdU9k2n3ucu5VotgTPJi1GyPdr
vNsf4tyduA/MBgSBZVi98uyBusXjZnuzdUvYhBZPspXQI+nCoVEG9/bfJvIswTwj
rVsH+D2+KL0z/hQmKj/HidHYTa8sZ2stkZiofJvDffxxVZ7P9JYt7HtYRTG+jOk6
xdpCWdZ0PA6PGvo7CGpGv55j2yEqwe8yepW5AJFnvKHDrd+n23xPBQnbJibBmM5n
5PJOsoCzsDUYCKTtc/5+fyw0pXhmV+toQiUX+DNEZOsIJZYKD4DXVWQa5a//V4+Q
j80uluFcnm64pDMc64wU+hHk5XRjcEP3PBeS5PRPpADamjmLYl8+y+CI/BUfYdWA
UF5fZ2xWdaaxQqRAUaf77EdNE+rvTMcH9m3UJ2LGOgHDlLaY9hFJxMH8ansZmLRX
blRzVlONh+1SmnaTfQHJFj/2gSTxEusRpWcxv/gF5xzzgJtMFkAeLhaY/FGkcupc
lgb1y3CZ9DamiAygsRfNXYo+abyMPXLLyAO5+wEpl/9ePwaMyHbrWPOjRX5gD3Pq
JvRb89AegVqM7JwSgnWjUgqQ4uoGrv7MrP95N9Qwo2GULgv88WT82rYf5HBCbMNZ
1Ndnwbh7HneCBU8h3V+qwQgevc0rD39lvNF5kiizPZJ6HRo+5IdHWFtjQHKglSMQ
YJZd/vfFDlaOFoUG1RvucMRSFW0t6VnoEe7Bvdub4mvJBXEApgNE+u/BfMxaAJCf
mgeIw92ayJO86KGfCiFhjIfBeJFsO2M9NRtgQJDui2OYCB/t8Eee7HPCxh/l3Cqv
Dsr963Nxo/eCuDSUxe838BB1gi4Pq35AezpuHpRZ1Q43ItxBcM3ruynoN/DyvV3N
AbIzXvAzECYj/ZMd+pJyV3aCfazFID5m3wn/fVMxf9Nq5xPtaG/n4k7nBdGVVz17
XCkLtuXcXYWkY5gNDlgCxAdrTawSIZeOjwEOI5PPGVzSkgcsAMroEUfxK26T+RKc
dItl6X9cUuK+12/aO91OBBtoDddN72d6foqlqwfoOtGHHovPuUmpvnASrdCyymCe
tOyLv4QDJ7X2LYg+aRGiXsr7cRT6hv0xm3Zz9tDdiddGoNgwnvp1EHTpySvkkyzD
irnMLkQ3lPGnISKl/9ziAiwU6b7HSAmLibA2AKTH3gUvT56EHvq+SQxsbKhpZjKk
2p8T42ibYjGj10be6vPvt6ETZWKTgLgOgeNpEx6+SY7Pwn31Lw1L9gnC96dtu/0c
IWIV13jy+oE6j2jHvwzHCoaLnqFeML7RLldGJS/zd4huDNr4JtwGXQkHDUPZEMKt
kgN69CToyb8tczx+u1y5SmkB9cJyTe5WftHD1zB9dM9M254T4rYEOa3G48Gzxf/x
pNiw8NLQvXS/0+LzCt5BkWVMopy/F7EMHENVqFOckKb0jl7PsSdtOiFDLN6fZEon
6ZXhLn/nRqMvK6G5ouK2a3bEaQAWUVzc4LCrb1I004CVeqMHbfHtFjyzDt/SJqDr
033vtQXzxJ/vqKLe4QEIJyRNcipf8iPvevPx+enjUf8PFFIPx7mm8l98pejn6d7W
K6MA8F8w+JliqANHK0ki0bTcy1Kt1VQf2cw8JouJ9LT/lMoE9ceMkACrUGKjzOJl
gE2Q8GrbmDQdS/8VLsQUd+5asX9e/MZZXqh9tuLlvJfBivsXD8dbAc23lxMxd0ys
icgRghyCn6UuCOTjoXN7WXQ80rQwODlceBxlqrj8QiSDWOYl/kJeXdJziFi2M6LH
A2kjhh3pPfXNIUIvud/4ue9BXsuM0J5kGIz5MMCp+DZsXAbfFQMiuyMIMy/bEHe7
3OcSXR64Rh1WaMZDy9uB9fAY8rHg+dGjTsJuVqRbGQVOlbsaROt82eoSRlVUvpMk
qr2V6cP1W4h0Ap0VeDzmppPdPNtIRqJQm0EO9hkx12COCKGuyO124NEj9bOePsdT
1gW5MV6NRarEjLEwVariKYKHcPyyAzTi5TzeYAtywPt5f6f5mvXlKyufWNa4aFv2
xSIilw5sYFQPSWLjxsiiD5Kmy/eN57lFmf8NUAiydqX1L4KxH6OhZb/L2Khq+F5R
7TqTFgj/vuRyCskZKsc74kkyqCTM80xXgAQBfzm37ng3BlAk6YaOkFZCsSkQi1np
O2hdR3/q3qqGNR1R+yTYNiMY5EGm5zFd282i+TZuhXSHEbtZRzkLZ332Vwss/Dbo
SDzrV7w/xGoishN10bk2/vHPLR765Bw/UA0iZfPgy8Tm9xCs7Wr04rWI3RsHnnsA
LyuEc5FBN1FB/S7uDRfcNCwlnwAOgF/bI2KuZ7cwhdFLpbiIdfcqV14oyhsKlAmz
xFY6B8Ov+FHatMcRbRR6aSX2nURpEvPRy9PYx8ZETl5kMm8eHcjezdilepeK5Jva
DYliwq0CCTW53sjRczyrWLOQVm+OA+LNljQu0hSaGSyeVmNKem9dzl3MgiBb3wju
KWy/IUC/FZUHrRo4DPpDI+9UT6v2Hg4OiB5S543dKtChn6EdfUi71BDTwQHtjDUL
XyW4C/JPypoGYHuiAmRt3UCpYHDCtNP0/igd+YYJwPENp5ljs70zX1iGIYovFYse
yys/l+pKLurs4fy7R5xDU6H2TpYBiEB5qwQqG+AZtuFn0IlpuMdu+GcDsKMfQx4K
hju+cbU5MuXgLNNMJkbijtOU95JGOXmVb38Ne9Dv4ClsIpYGd6XN5wmk+0ls0Lve
vSnnKok5Wc1d+OjWqNfYRulpSX7sAYILz2xdKS9+EFXi0CCYTmBoIBP29/xlPPKb
AsMdWWJ4bIv2o6DHU3MJ485z3smaeXeJ0Zt2S2vsU1NuaiVSwphhuPvjvGREyiZn
pZvTGV2bAPKniUkrzXiDQYLvcI0N9tY1svJb3cfi8xL94fIdmZftcRvHC3hhO5fy
UJv74oaTy+K00GrOyy3jYhjgGeFpLaiHSJjDJ13AYoJzx7Ixmwv7tkQtGX0Q54oX
zl/YFiQGfSdFSv3JfGHwnWpOnf/VsAuPbFD3Wq4qQIpAqb5OyHYmz7aHWmcBw8IJ
euEMQP980gtNTyht8mzcKftqdeamxU0bkJZjMabt6YsaDftAdZzU98aTXqcrHytp
EO/NP9csqOhXd7HsLPVTCYGerCDgg/2/Cgnv2RucGcUE+cgAm5fx9idG9kC/EUFe
FAnQCssOMrOMAfuuhKXbHhxGuymOrtSD8lsu76J/XyQ+fBTyvIqjmKwWcK4SVXne
ZwyoKuwJtt4Me3S2hPFm3T6dJA71jHizfo6q+fLwF4RCcUSIn9kxjk07N3Tpe5w5
nSV2z232gmC4mcX9+pyOgGk6TSOeFhkx2jBgot6RNLSCEx+IaoGIizvmqqtLtX5O
4pPOQmysS2zRqXc7bOn9Icswc+fBugs1L5OWMAp2C4dL836i8RSWZyAM5yVN3A6P
yu1nOCjd8UJpvT3SQSY8aTlWUA1lVEaZUIew3io+8r3gvMjG3ZLXY9LM9o2dPnQU
Et/arHlTIFv2fxrfWq9Yi6rLCmW7ZJ71IVKaoj4rXbDVzQUQ62kteC4ewrb7Jruk
rr/cc1en8+4CowDOe6tEXKxx91Jugmcj2GYMufvW78/TkRZ1Ssc+//XAEJwvou/Q
mYJKqZzOqETLfUKLV2YS4Pduz36Db3BxMLijQZ2CIfSBp52C0la1nv4+WD0Lxrfh
Y6MxiGjZEfEkqiTwKiNGz8jGmrxwgYfXE22p1T1+f5CsCSHIZhWgUu4om+eBdAOw
sWoys3ZVuUlbqSmbyIJBFPdfwyMNdoR1uFzIKp7V/e4WucICqQZMegm6eXMRe9Oe
2Dpl6JHbHUQTpQBI1H9ChIvJ3L0t96Rtz9ay8VlFr93hJOJLxL1NloP8NX9Y6UZ8
oDpEzmnvZm+GHjHkfHsfyE9EfVY4g2KieuLZW8CAihS3hM8hkRBdO5226ww9Bnqb
NUkk4RVjfUdljfI/V4mUqx1gbety5VXLmHqc2UBEQSC76BM+4r+751xhIGfz6C2K
9TguAzcB7u1J5orr/G98+hiN1SpO+lyxFANrb1y1TmI9NfB+F+rPSzmSRG19qfXF
HB8ngMdUKh1FrqGCS21OCCa6LP0rtXA+857GgWmFXk4LVd/5CPirw3ZsPgYcmLle
eThSEwp8htdo1mP7HC5wT4y5wfzJP85G8BgnAf/mvAzrv4yV10r/ikSwmA2We1DP
HLm7VmoBa2MQjYpWnnEBTajEjUu0iu/jXpaJhr38thfs7x2mANqL9sSrT+cjqTd/
wU6izMM75hGiCqOTpoJVdZnTg4uHL98YAM96LWXe5KvbbOfNC2OWUV0V/e9cCjBV
XyGnbVIeJeO7UFOTZDQE+G/JKIROS5C2dRODX3XYls2PtSk8YWLEAoh/EQLxpitx
rxnpt1z0+IN3wgCj+dUsVNTT3/L/0NfkW1BwtzIMqg+KFTN252+D/A+D73ytnT/2
2mR+A5yikS3G1OlyExzJu0PxSBC5PUwBYwuQioGLLHwNDM18AlyR8aHQmMUdEU9Q
XIYGTeGQNwu+ySa729bmv9sHDzLQArqM97SJ01iwPSof3+6Ia89fxVnjchvRfxPh
MsXhx2xmiQK2zlxJPtJuNIDhhJSea+ULkzeXkhPhB6ypfMhvZ9i6TznaS/+VDwaJ
JKJEjVhDa/dWek6T01TU5rsMASJRTWisp/uT8q5ZjR5gdIlPmMv1bofZVJNTq7hS
4KKFjyJlEzIn110uqnQv1/jm5zbBt9Fb2B9wtOls5MQ2Zu1gYt6TfBcogMI53r9U
i/nvB75qpqJpSprcIL8iT8iYBcQ4RrVaIDy2nGvHN4b8rpWWvuGlGftS5PCnapun
hVNytd8TtJ6HJs/k4E0xyVfSf9nehtY7Kc8PNA5vymYf+cBdvIHuAeJhNBNw08PX
pHmiU5WodzUvowUy1FJQuIW5I1NvTDwS80eG0UZewKxVFaT1D2c0jdfoZl3YWooT
Wbs5yZRM+llkbyApkFGMhgglkdrpJcsi8cJC5H0db7DR+ApPEm8sv4kWCaXm5amD
GG+jmazpYk13ogT3WnCAV3TdHvuBHL1tNahJ6boDASGm0CW/V/0j0L1JaQlIOlGD
GJZ7BzCi4bfFOvLki4pkvUDzh1d8248daap5VXSxL52/hDsg+3TiGLwXfDfdy/BF
rmHIji7qORDjtUemb+a7VztCpRFf22Rhu8Ffo3Fkz9FRhY4msXv5OG6Gd5hJaefd
VRoVI4ZJTkFO5q9WZket77jxX0WIV4SK9QmdYWcDEwewtl8E6lwQ4jSdjR2AbKSo
9SrvP4zPoerfqpymSVXMab1jkEbjqvunojAK0algQQm6HMnR0IuyOGJiXjCuc21D
hZkvegfJK/UbAjDOnlrIvVNdt5Upm8ZVaKMH5ljBkVaiiMdGARq5sEVnS7NJZqtO
vxXkO3XYhyETyKDJpio1kkSztQa0iM6gBLcbGIK0YkAopIrvM59zPTKUwJi2fmI5
2blM5GPPXA9t0qX2uZ9FhKqpKECIMTmpmf1fiNiX17ccd7ahnGydaNGhFEVNIvYn
84syrcI0DJyf03Swz7QlgjueF30DLSSDBcP96srgiL1BfxkadLUiojycUaj2EpF/
Yq+mzo+kD74b81lrLhy1FxxYuxBKGr62oLHj81pBVe7fhjJQ5h640hQLIA0MD5XV
yjzUeKEpdAG0M/bF1UqwqQTclvCFVuQIvUWf0n+jtPctTPJGrZy+0eP8MmpYNymQ
UB9/qAgwLNe8f0ww/M9ZuHKOB0jVx4z+f4GsnpQyXkLcnNnkri2jpkidCvCa8f1l
yflx3sqwdjjC68dymoAyK4oJXbDaD3LG1mG3AL2jmssbH/VJatxSKB9UYTsecqmr
8OBzQMGR6+1/9xAbRcD3ZrjfjwJYbq84TO5/SZ/xOf1UVN98CZgnzhVG1vGa9lDr
kmsJoWuYyn/+iiVGZErS2VhZiHEfCMdTFYt27O+1L2xKQyDMnbJ6E6YwXWH3eF8c
wHJKGx6BgNEkfCgHGKmt8Ouh0MO3FtyLJbHSZRJStmj5JDPih7aNzaLGcWcpf6NX
3ye7/FJkhTT+DLqvKaYHd74mO3WCFEfKrPabMKxOoosZDbgablZe+kjzuiwHG3gq
bv5ak1xND50H//taBdFwxFTwZjAaS1SG5JCtt+M9LLTnGJfwL6FrT3ITo84NZCkN
zZwZyItf5IyV3kf3DQBu5JpcxanBSK6oWTQOXUguVThkfGkDYirGj9Oi9rlxMMto
ODTTStGCKHgj+5FT5fO5LZaZ8t9MjZTAxWFv3lJHo2rt5S2S5aiRQs3fnl+oc91d
p2ID/oZx8z3hwGDjNRVY/pEP84BJHDHs32tvtZQTfjgAS5LnPScZDnNV3KmicbFa
8Z5SW7FW3upHYTyuD/q846vcFHbNxOFPwj6ni0d4wFD44Pjk27YvzsYmdSe0NgKC
8XGn23aSdvv8Wva09ApodGW/ZeG5t5CVfHPvBCUP22mt2JnzPK0pIbfRBUPZRoxe
EHkTOLRQUyrVkNfGnNJT4gHT1o26MLm9UJ5RiQR4wY8eP1H9AA2fALU2aF5BuOex
Z7wepf+AlKvZcSphIIsc7oQ2lJl1iq23RJywA2UFw0ZXIgxzF+v3zHDJYRyiZOHX
9Rk4gDh55m5jiEbuQxyNeZrwnrKzPJHozMEa88BRzPTHFD1Ys2/7HxpTGwLcW+GO
Am8dpu+uhXBUZyUkaI/F85RVFGxYZycwrJonBuA45i4YttkpJUIkTaFUYyRfjUS+
2kPf3l+91D6NawbV5uTOyJ7OREhbUAEbYj9d0NbuYFqfaUC+nUTG/sti+urJROMy
mSDDXZnqOJVcYIjEOArUNTXecIUCBzrj7GZVua8oDpZNjzzhoHzcJ1iZtkzxW43s
FskjPNP+dh6y0MtB1mDm/OrbAcxAtTRD3UkOeCoeHnd+czQ/lPFam0soF2Z9Ocuw
BdEuvil+WW9C4pEjLpozMD1SkuqQE2GBYq8rnd9j6mX/X5p/aqdBrmikQrsjlsur
MuWJ9P+ssQXbyoOviIj8ZDg18U8Mmemjc7mt13RXyzRfhlWV8hlDaWM2sSXSBNlr
16pI5Vmw9x8Ka4UxjPyCY2t+vB9CfEEnkFAUnvSPMp9eA+XDXsTSmhIg5vs8D5PT
lRO6dM6pOxavXyjzfE+QMuW7kNbbQewTQG4n94alsaer/5qMB1gX6MpfpBwLe4lo
n3W9G0KVbfNwVNWMqT/dkaxL3WPYnSfkMur5nAWbb6rO3bfegXr7a2mSpcjyngVF
uXBtMznahVMpWOkHDPU8n//8ejxBiIJHlrnvavzxNvfs/iophYqAclOu/05JUW7p
VqfO6pOw0TZ9w/5gq+xDUnZbdlXQgGVMZW7OGpPwpmwT3xD8sss8qMaGXAHzC62w
8L2rQte75wkcOGTWtcIXbcPLHGqo1RgHpvFw0C/NTh7fxH792l4TT7I6hIVK+ccU
KEXQfkrF4f3K0OeWN2WEvjop+EW6bdvD4GSfY76xngtJP1jTTkGMrEbTPWfw464N
y/gnEEh48c72jDs/K8TJjBQ3+H8mpsuxsgcCAxlKAMqbIiPM1S0835/5ctAEWnL2
57mSKPMZ/jEsfUrvf4dF2S0gSrFbI1zVhlbDBJQWkm3TNOmkrKZ2MHHELbeGFPar
HsCUCrDoq8eD7n1dDf1MULxH5yVT806oWnqf/t5b9c6Ik5cAnXSTo+lBAw6mGtkm
ILISC3QEDpygtehqtb8W5ghzZhF4rwAAwTyQGyJ3UApQSvuqUMOtlpg+Pi3ov4pR
Km9A0BOq8iD79n5/etnczxOLwVnYRH7QpU+UkxX3/TuH8kaTBk7G6EGuyF5YUjU7
8qowpFofYmKu7UMef/ZOS40MEwodzOGFUCZmptwnq57wmi1lQ7MLo+L4/Ht4nP13
DB6OSHqbwqXrIzJ9XRP10seMBqnY/HzZzUlZEZhlMIppFLc+cLfsz5PO8etgbHZZ
3k2CBqho7IfecID+8vB+QBfuox8iCVaVpVKLvqiu/p2CP4szMTBx58ta8H01ql++
2YvaC/3+hs7Mu9Od1XDhkv67xkMsObAbegS3c6bTHFZtDSUbF6gwknlR5iXY3Z1Q
CQa7ABlRfEaZ4an3s6rNU7qZ551vlqDueCAtgLTJMAuZJQkcCRtxYTVQIt1g9NZR
/zvLJ4pyJ7VodMLvuf0YmCROHUe0kat0589fCxhdmqctrmUW8bsmp6w1kXwMHPae
JEGQqm1W/RLOw5jFT2kPDAWgIa5fVY2FC3loc1tB1FclPKA9Fjc99j+3Mah8Jvyd
/e3PAOi9Yu4QnW+Sku3qv2qISig/elfP2W0YgXqa2g69uU71xsK4rNqt5yZiSPaI
Cm4ZpkuafewFqW1qt5QuA5PF9XJXEL9aj+7Vz4FmA2zGLaeS5wsYZuiZHdwVN/Z7
8jUd4tJWcB2Oh87Ob3wGZonDktZ4AO8Gry5bTS12ecu5M6jOA1w2F4Vcfexe+tJr
WLFK2wY0jyTWrAmawbU3xJUXt6ZGlgNgYzHLogMEmkp907/lT3FITut69P3OG3IA
0d48Bc2WGuKz0hD7MQIcSurwMhb0Kp7XI3oQhAPmYndy/S5xn/8/fkZnTtSnzyeD
QqRlYppjENWmA82NC4bY9EQYczdeBiI0Y1kzKLQH0euwBJEp0ebomGUj7JvXpUuh
8xKaKBDSdg2+7rvJ4+6YHVDfIqXQRiGHs96NqpFjIggOEaDXcnLbS69QEs2enWw3
xydAwHui72eVUNaYjLQmOTNsRndkeq8BHDPn2dVjVJcnEtMxRWgFjsdgDTno/6Ma
sSrKPvLuxRSBnT/uhpJHdWd5XKaBlxSodZXtYrmTYv24eXMJhDGuE2Ejh9OTcjNB
xR9+ond+vFOv8KKF29nH7EChyK7ZoPZvVpuLhpLD6EwVRqGzSGW9zGRZjDxlxOit
0ou/7d6Zyn0aTHrTZrcIKbd786gQtkZS3snj7lPyKhMFkp3RW5qzRuJZpb012SWz
9zXB938cBBjNjNIgY7CpYABxO4iNEwBGY+ilct03hKSEmXf2xBh6JrNAmbMAMR7R
eKRPRCNTBrwMIDKW95LhObby+14f8SsTHar+EYj7ejSy7nw51rJsepR3j63n7nKX
pIfpGGMseowPSBfOUy47ty3Ttzj7y183SbQU8qFDRtdDPrMIeeKhcDHmaySj7s4t
LJ8fzmvCcpX9dA2bANf8LovA1FbWczEpNWPpjp1bbRa4G4sDnNmI0QaSRNUwePPR
wZz9wtnLrhjH9elGNzkkLUH4PQxDl/4Krhy+aYizlraHc+04Khrxwj13HasuGw2q
dRfG3CJom6W/EOvbPTznC1E4gJ6mXCSHb6ebuo7/tRd15ecw+iq58dgupv8Bp04p
TLKPgR5Fw+nEFalmATUIN/5GB2DiJt5LE5GXe0Znkid69DW65RC60AnPXyjP0FNd
imeugIK9d8ZxVfKW3RqG7PCnwathnQwk7jyNlDRQSH9C3YDY5CwKHK3OF6/Y6bPm
Z2ngWZG/lFiXkuLipCjEx/nZVUSFy/xXo3kADsSKqLddFR8d8hYnkuwd34XqpQCv
jrwAHSMmzfcpjoIExYRVy8CIRl2n+uamSTkAhTOg67pAuqf9JQhDr+lH5E98pcLp
pjZsuQlLu+qWdTb4aSUeu+eLIOBR2wGcMKbHBneBt1XQqIWwMO1fDL87ckpQEZUP
69ePaf5glZP0VQCVGyCNeX8kDOKjGx0lC6DjTQbdAfvHXbr1jR6eqLCUCe7ulgEb
jazK6yt7tqiaC6MgxMWaHcaK+caGdpynLP39lCipaekIe02lWDa8D63LqTE3X450
ozRsOU+emdMCi6BL6r6pIvNjd8cmMTxitqflSGZyxv5UFExACDtjAXHbNLWvJPLP
Tgped+S5QNo1wXytgnoRDbpKqWyWSSpeZJ2iHUD4qvVGY8bHIX7hNFhzbsp5om/2
b4VyXw5E4OJo7Q6p6nj4PQugkXPWO5DNBfiiQQZXmWKIGZ7vdisJ43+pc3KIAMIU
HOnz0ABjO14JBz6ojF/+9pxtBFNXaKlePQlXXOZhdkz6rxFPlHKqDcpfJNORhpXp
y0a0HKIPaz1RS++7sKuRFg/nZPtCMl1z2/WIwA/TekH9oeO7GxXFSFA4KFDgZoWK
kEOaHKa+HwbpfS7Ux2YjCTsmWQEGUrNhHGO6945VS03K6II3FjAeNvNLWwaof8wJ
Bwq5fbWBruZhkVexpUckMLjbtZtG1eKtyipmfomq3rwg0hCAbgqnsVRRMuxB+nsv
BVWongdCmPjDB2xEhz3+U2Vf5dhMJz97lV6st3rR/cfn/ve7Qd5b+u/Mech4Rk+u
0uym2P9I+yj+8XCE+a/EbsBKqGB20B8zWWGq0Epbg4K3AJMWk9bZMJh0pZIoTqNW
792X3VRqqyCBKA7OZ7RZ8+B4I5a7liJqNYOubwC8I9jRtBKC2k/vfATDv9Bf9Yu5
EF6k5tNJJXFG5qlJAn0RmLUMplS2kOQ8zsEQYcLhaS1MIFl/QQC3BDq7zD5hrDqT
Pvb8QwzZa6nAe38QaHPC3VfI4hnTxzsIcBLCgU44E+HneNIS+bp6FAlFWvj/jdPt
Ns0Prf7dGCZZPuyVrWP5gsHzQrMt6SOtBgiWyrMBknAaeRHL7xkpkO4D4dK7j6T4
tQzl/uPi30CKv3aeT+S5bNwqMIh3bA5LITlGj3p/sZ66dQFQuJ6hgQJcjknXA8/s
QCI7yMaxp3YG3HUEcEnvuaq60WcZl7UquyQPfcq4ukwWIlaNlERMF9ZEfwULXY7U
p4UaGHUzVP5MwoPnnmTTXzg+NidMzCHotQldzNTq4u4QHm7hl8DBjVpdUmCSrZeY
SK7Yixn0Dym7AQ3+rKCAIhzAhsu0NlSxdLVyUNI6OD302QaZv06RXjwHf17F4Q4k
S4ly/yMjY7x6GInHLrYR9uvoe8YIr5YKpq9KY4s+vvWkO4wOF+JvbhWnJPFgEBNf
ajsGKiesFkyGJVBbh9EvugTqhRymjua+0JWyfHexGd+NGNUE586km0Bh162JZSz6
8FhHeH9G+tRetVnN5bASzZcOdUR4TGqlhb1qsmwpZ+8/SPGefHYmEx/rpFxu3z+I
dPR576ilEV4x4+B24z9WpEldSrSg3FK8VSM7UIa/LE4l18DEthBGsIBRFLRlRO9E
czXXx08+qDdKu7Wh6nPAOS7SVt3uvsmiPlhCrAzli7KPDwOOxD1RVoGrgrnMF6d9
E59x9/aZo4+yy1zWkQNgmVgbymO3YTAQNo1Ra0p8VxSJtiF2YWIldkEQ47jCaLOU
RypqNRgQkZ+FxeH7Ckg5AS+WwRWIJOlqrBPlo3I6VJqqf6aFEFc8L6j1Trvcfsbo
WDYO4NOr55r4Dlu2grihInYX3/Dzwo6h8sNKUo8e6OJX2c4svT4v3SVQgOHiJA5B
H/YZwQTlGz5vTN/ijMKd+bcgF5SSrMJhh9jRgR7qaSJ/X7wG5s10vW/JMYxG6e2X
quP5kWNi03n3nlQCfvX1+xkpVZodUCHtOx7Qdmz9jiziVYKTxs/gIbRAJeD3guk0
Mhe48DIT0BjHdD45QdB8xIAc38/DGp+7d8vfrjFcLnJOwehX5JQj11G305OqbKhN
cSaOYkuYT9d78+zTjGCp6CRRmBNZEM3By+zwV7tcxCrlJduqsDCASbUzFIlOFhLR
Oo34ek+9ipy2jeRcey/G6C/5LXvOQj3Y0k1yZu6BeQce4iuBYmjBTUxb4GjZdnHp
ZPjjecs3hj73/7OTKQFK9SK/qxkOmrnlzSQxfaOVcOF91XwUPkSXrMPU4K4CHKVd
ccRyfh4MkhPYvp18ADgtum9/Sm3vF3nb/5CSImeqtQ5yXLx7kdKwAZZJ2vFMzgFP
kTMx4HIoXhls2R/0b4DborkIWZY0xkru6TrSBAGUHU/VoltoQ9wSa9BUIfiu7YdT
+PzHlN1sKKYCzojhhuTe2g4NyFgiTFS7BbBBDMZK3U4y+6TR86xQhXdt6GIxuIXL
P5fkE7tK0O3qSJHE+JiMWU8+vjJJQ6RnKV4WUojojpEbM7Vfn91vtvwwlxGIX6fA
ozQIMrILYQC8xFZdax+u3t5l/uqg/b7oZmXSj2dXA63yLFPqJnr4Dnk/IWBEvIna
OR4QPJ87H2HCW18q38sxAAqIHpOIjcuDZnQEoqKaB8a6DSaeNJcwPn69jRZ+u+wt
lsuk7H0p5uuXhWRkOhyow+Auj6/2yfJoMmSJ/fW5fLsNmW9ny9SY0EJAM9FFbWE2
3uqavGi1AvF18VQcrLJ4XH3yC6GYGVjxljoBi35i9tUkj1dEzY6rER1p8q9Hebg+
X/0r2HzN6O4hskgIpIGKlNHyS0dSDr7IbeQ5pi5Zyf/1B3qsovjohrjS77KACdWS
Zg1pptqxJjFZCQ6gkxfmuiydDEUEHDx50oDAakmiOLi1Tp3UOObC8RRSK28Jx8IO
A+G0gLY7emHWzKahLifiTRen6ImQpwK59ZhKvcvm58n08TRDrWDUcUWay7SrIyFm
A/coUYgW0hDQmmrfTzcMCQlx/oXkn1Nh9YjjDqyUtYp2FTyGCh9G77uSib5i0cVb
PJLjkazG8znCCKBmzTzde9DFZzp64woJHXVHnJHHA7UjBP/kRRLdpKDPkAsT0wF6
eVSxz3OAo3JgjHakydFYpTiYp2IhRJenHscmpPdrFjz+ftZE9AOtdeIqhwoGzTmS
HUNAJ+QRchrFYps7iF/W8/NC+F8Q+lCn3zTsnAqjxndbaOw6OlDel29E3RR3HsBE
QlGDWC/z66A4FIiJEVkHCHl80ojkvq2U50xDBE7BcqmHMs9PbrKv7/GFeaDZi+WW
O96if3gCShR/j4JJIZuSqmTmcj+Sy26kfhXTAKsVaXmtqfB2/zv06Entv7hMS88+
kanI85b3AqetQZKKQ9xjqlFo7s21zhUpBh1tyE5x8pWEhX+XQC+wtOAIwcoC7zFE
rmfgG+HuCgdextFYqMGZXVy9OJq3Gp7OadkiagDyydqNXXLYfdFJOrJLHUK6wA07
X9M0JXJ/ySYMv7ImKVAc6eWB++SaZS1zS/abt+kyxZtAbIXzSkRXSshdY6TKSJB0
yNp/s54nlwodqp8QIfdvPSn1eTTkXPwpctTg9KGRyfd1ggy5eWkDYP3MxKbFwlj0
3ZcV9eGh6g1YNhwaSKhN56odXcuonN8hi6U31UznmIBI4BVMXbZOjLngNpIb84Ts
cS3OXTWVpE92irSG+LyHwH/K8OK6efABGRIzOr4X2p9f93fOgA/O4hshrVtkTXQ5
S/DxF3cqfx8j3ZcTeTdf2345TabMgGl7K52Y7HH1pJ3zGTHOs7OImVAWrQsO3qIl
jxNENpUAYHPbY99+7oroZHNS9ycIYljsYObdcosb8bxxpQ2HyutC/pLZByUVTOM0
jYevHcHKbzjOHm4OnImOY9Sh1gR9mKXFn+ovrgItVdWsMJd/onTT3Fzlh3WXnLY+
xhF0m6t2fgzlyJ3coeBOgSrz5LKhKryBvuaV5BDIs+raDIw8jkEGklvt8NcrioJV
DEyg6TotOKHLF2mkZTROPcq+zXRlkaYa99unee1vuxTRB/xzmEMwl0KjeIGkbvIl
heb6MTFzO72VZxJPKjFz0ZubQQn4qDVe1oFgcM//Dsg/d3AfeQ2a7eOuv+XP+aul
CcTzQH4tRKdJV1wHBYoIdQHFIgP2S4ka9CrkKOTqFO9ErZYfAGEy5U6g5jdQmY6d
wnK+ti2mVJ22LeBWVpQlGmCEOoAbYkT6lrKVRbZwIuGSXnkL9oYeIH7RoXJg3ADI
PvZiIR6PW1in0hct5fgWNYuYFOyaB1pBFIvNgfWvek0qvQFJd2ehuzU4EFZlWNMe
wPVVuvqzloInn01XBTrYyKFlS98K1UaFUYNmXbOV9FmTfpRg89Y5jFC00IP1jIsS
HOj1euDma4lhHvfsWWdFQQks14V2s43qfNJE78z4NbcHTQQSc5UER8dW5N0JKMlM
fPDUgGeBEpQzFh1wT3MPrxrBBXbUrRyoOSf4gET9BTvB8nRewwRJYwabWhC53CdL
zSOoktZZ6oumaQrRD6XJ2mrTLU48KGY56n+BOl3EXfyAAlAe/KntUEkOK7q1I90J
9FKY4/JLmaui7jEcGQtQpe6W8Oq3azihb4itBsukNGSZdKiXsaEmHVI+EPovuI9h
vVVAdQXFLnjLhE7ToVqjOxIi1LFJwxs6VbNT62jgh5xakA0ZWTn7bL59Q2tM7zES
QxkAMLatfZSlIA76p+LeELgTG9PPf7XRGX+LAyFeBL7wSuaR5kqhmHemAPqnfN2n
f4XWGAC/uoYq8FMXWmzANmWr0FLa6+Vf6aF0pb3gGUU11P0A57OG0lWbWbHOohqv
g3wG9J4UajIGugBcD/E86mTjSFy2AeSCE53OgTuJ+S5OpUloFLzv5HV7NV/SuQsp
WygGTvkY6wUjCG3JPanQed5BKu26S5rxJfOJ9CVDBUgvv69tTMfwoK9NLAudHLri
OOoo1HuA24NgKlvd1PT7dTs5PxVErIhU2SrGO0Y4HEBiBtEuPUPJbZxTIL6Wn61U
3epio35SWi2/8I2m8XOvV50YsE6ZBtYln0irxkIaJ4BM3131o4urOpG5e8hW7Dcz
8hrTLJIRDmS/DI2OtexorvhXKYvnx6lA8v7CLak59S5U1rKKN5huB3D4+p2bRG0+
6eSRPpWU0BvhHLQJbi32aDezqIDPmigOzN+LuTMj6vDcKvAb3IBnxPIDYqFinOiN
cemZhFHfaUE4/2K7pQDW5CHNU0EbLLHaQxC6Y4YYJ2RnlT2zP1rf/DX/wjz6v86H
cgF1jBImT8UcND5Q9xjnd3GJPg8Bmz4cNglxmiedlXxyJzo2EHOOgz2YvIhYlCvG
Ll8lJJEJc1I4jtKOxzeRWUeVfpTMgOHdR3vs+53Cyyr3uGZbUabzwvX8cFEF1/yM
uqQYlr4vGcAcfZjxGA6kvlhhHYSTEvaB53Lnz+Mfexd4fgm7+S8Q1/TX8yfH0paP
rsEUnheJZ2AERON/a85pr7+4PieqFnmXT2Zo2pLi/s5D5bITA91/dg/ypwokQ59H
miGAlHHbV1JZzC7IM+vRmMMxFeGmSZuDk3jN0uwp93p+I5v/AZE/fY5jVFVNaSja
I+BvB9AEGe8ygU82+lfaqBmsHGrX7iOdW/D3g1YUkbRfFG3aQYc9eGnbXQprWNxE
YGoAjjz00r4pSh5CKpzPpyEE0e9kt6CjLXx23mUgav7RIvxgleVmi4HwWKTTj2gh
55mJcJPRYaF0mDFBq7/e1wiN3WhieSWpwtWWO8BtYpo9Vqb2s3zo0M5VW/SlPj2t
YxheZR8nfNdcZ45KSWOFxqz8DSeoZqmAfonJ77Z2z7P/UkvAiD4fMeNzaUkwV1pS
c2yxUXrbIAX2neBYMD7rIpzasxoE2qZA582a4oWqC13OhRf62nSU96rkElODHpWL
SrfsJssonwtKVAY5spxc2+OjzQMobRgKunY/FzjPZ1w7utHfNFSPw13DoNGziLJX
sY0JtAT/c7KHoIJs0ba8kW3XZxVPBSuTEngCHOOLDHfpvuJcdafcWEilWlmxsxMg
cX9I3/quJ8KFrc/ichHBNH2sXbuBTnmwPZBqQj82L0tGJeRRHrlZNbZe4l5gUt98
jiNHkkb4Z2pashjNr+OX841qYokNhHh5vnKJ7nBmnD3OtCBUtTzU9LLABU5E1uSy
9PDPOPWAK+utlNuDRwCxd2OpkvXFXyBMRUhGGftZXvDJ4MWHLHdWZgG1mYAyScjO
GSfqdsCVRJ6+2akcCs2p53A8kn5waGXrz2xW7ctQZ0oj3GCX2/AkPpF8h2V0Klz2
+T1O9YdVW4kqLN9s4a3cH+WQOkyjBetkdPHnh8mXB+ItN5sy+A+mXes0Yyz8nezu
lYRwVYw2cRa/8P32UrlX/BD7WfWdZCPb5Ctn5W3kpanDpXLt7spGPXjNrVfr8BkQ
JFv9+2c7C3kmUDgmr5zVZTKCmefLWP0WubW01XKXJ/tARB39TXBhfQ3dyl4f6og8
zLCtfAPCmeNVlvWdY69uhyMadNtzYJD44ldnfPgTS2yi3I6OcpvKHY8hQZZVlbor
9gzo/4vuAaLNNAHtpKvF5QNcXGsmNV3Vv7do4x54e/LpLcaeO9aE/55CnwE2A1Ni
1hiRpzZQx+P03kibCtNlfEKkj4quPxDqX1FLPYeoopfc5XKytyB+TNhk1I0t5fQD
cmLtkRjiXbVOjp30O5kgr38IUYQW1aKCC9cGfX3G0f8ZIqzEfiQPfwU93sL+HKOI
T5ERKNo5z1vOIea23ZE0BkkKI3nJ3QhC201l38azbdqipsbDoVKBYVYdbMyxpTr6
sjbtjPyHhxjvB+zeY3+6Tg+puw7FytodQP3vHZRErbrNNeXNSnZggUzctqhy3veJ
Egzkerw4NitehCnx8/r6J0jE3rQjULXarAS6CZnPopgfpHSj9r+yu94Fv1RRq1ib
BY5jkjMwJE265kLkuasahCL/vdE4tjIXjPIfBAgu4C6EnLhRvSUDPBjc8rEXa0Az
E65pBGpZIC7RTVux7iCCP/sWniM9fHFnbXTsXsxF/+3VveBNCOFkWIvc4wg14SNG
u6Mwg0Ol+HNKJ9YFAfiUn4XbO6geRZBFMdUoPrLnyyZCR6airr1TBZmq+Lc1LzVS
/bDEZb1pn1IO7QSJAhCvqSNYxAp/QRMQAbZC/LyOE9SPsUcecjXwzoKTaxTE1uiF
ZhcP+c6vOsI4MxwBz5iUQi7QLH/fcey3BVUOp5+TUjXNainsu+gLa342ey4BA9it
uqpA8kJACEqsG/Jy1Cl3JMBcZO3/YU8JkY5420vJ0cJmk1e1s3GvnBfRGc6pVUfP
hGO/8T5X4MqxZatNDBEooZXY239xzAiaa59yOHZC1HvkO7S5f/HJKs14tzzRbffI
EXCiodM3FduYjyvsN9goPqlVC2drilylL0C+q2u1sG0YaRFSljKWyr6njto9Bun+
R/mFqDedBhqKbxderEGkrjaKh/I/LQtYH/edIiUKZbx52WXOI0jbmYGDG8cpMwDb
CUlgGoqIRHSHP2JoiqjmenIj2aes3P7bChwARlxgmIJv1ISge7HShnOoX26toqHv
+R7drDPkWXAzGfXNxAmRZn4aVsG4xVMTtymuwD3V1jqZpaFSZOUltW12lr5XyB8v
FG+JP3LHaRv2ylWVbrpcZiTszQw7758WV85v6ZvbIi354FywBvCYLrcVVH47kAY4
A7vXTTctaTTNztshamxMNwqri+zEurHdQaEiIt8vI4k1a1xujDxVI3DyZyk5/t45
46JTpzc7fSlgxOjs7ej91NSnKiOOAoKfyG7g3CIR6hyDZn5qjRq3+WORIG/yctwG
VFgr6GOwWejFS6NJbaG0avZnAhqVdHpI9sqBfS4Hh2ebJd+okFtqQNXVI8fgfaxt
2in48eV4jVVChAVzhLaaXMgbR7Pa0JtMUi5Ob3WpjQUCWqF2t7Mbw7nspDuvHIMM
vTvGyht8Arc6J6bQ1ukEsCPq+kAK8j/xqfiYpB+wgzk3x7AZ5ehqadzSrORquJPY
g1QTNxYpM0TeXbStahYLIhzqCPVEPgjlkTc42m3k4z0ZkvbFIkcL8tx2jYTO+u3D
Ms7Yf1+O/Wxu1h84C/EK6rT8otl8cmDOUmjsF4paUzkuabAGUm9EeEgrL1OUQ5pJ
ib2yegwKhETZly5Xu3Nuq+cIaj8RecMZ3dTdY2uW3KPhMWRmObyLdrrCdOKHqvPP
0oN4O/A0dAvQvU4Jb/Wj0gj7IMEM9y/h+bmj0oSMOzKq4eNmQuHFqmdPJiPqEa9F
qrCIhHKZMso0xjyfN+JGQMtd8eNAId4Q+MIeOtg533JoSGqqiAeg+uOyfqRPuND9
rQSrV4cnJdaFt6tYA9OFJ6KCkR/j5+CvxF8FWUlPeypZazsv1cPeFt3N/ncB1G/W
0d+miXjkXTGH9Ofxxo4e0X8EapfpTbfRpDHirpvVI1DCqob01soHr7M4KMW87zi5
Vkl4Aw3eWpipA2Ee3Rt70JR5b1JZiJWxiIazNdXbrU8ueGw2+eS7sEJXkX71bP5S
fRTJznwmMUdppfm/u1Q5fHFrB7Nxnvap/pfUUDlIGhmqDh1eDs/O+bZoUafX0h4q
VbxJ+Q6gzdcP4lPUbnt8hmSzrrA1Lz97G8Jpsn+IYZhbSag9VarwhNZOVSrBoy+z
Ly2uWeMqaiF9QHv77gpGiWHVy7yeKZ15W1aaGzsq3FvQBMUjtj2HQ56WEPcBC4jC
w7b4eeF5gKZd7XSzfNd3xfXmWC2Ik1kkO5d03WEjs08XORoLjLWUud9NyWVG1ioW
+kAUrqmmKB+HkJS1ZU7uDvlKA3W3FfMkIjOXaZ/qk6TGrCyxcefGUg0xfKRabbCj
Byd+ENkTAMsLDRzuFFwiExtPbEv/PQUGzWLTGUDd90gQbWyZ7kPbXbhR42206JPi
18xzNGODKDGou3QkdWmylY3I/Kvw4/J6q1t1Bt+tzX8jZcPg7+Mk2i0RThEHnbOz
Tkbyz5+ItUcVDvezB8GEnZUV25o3OaldRsIy4G9039KDuEvXyyA2EtvWkPLuEtvl
lG4zPvhl4gkXHBqsDqhycpmAK4ZV725A6eQ/6GcyjFsM1wYmLmgIjnENl8mIm5lX
B+MzENVFQGAZp655/mkW1EBshck4FixuErduSzdKeCbduEt2dDqH7nYT/vH8/zXV
I51NELP7Y94IhYdH0Kf80EMYnuOxOYVRJ3H25C6A6FhO343g4bnouqzvCqL+qq/z
O1ePdxaabfXAiiSjoRaNtJ0onPwEgan6kVtGW6J1UFA+eT7ZskdGy8TVYlPWXln0
iuh4kHjRO7PDZvJhA6YbCaBf/j3gYVL0Qv7Or9HbXII6KoDFnOpvMiiqSe9ezat8
37g5UC/dmdigL9FrXf10FaTk1lrW7BtjMEfuE+6Lw7OUoUlcLZNi7nWkGdRfjbCG
loqzSdGb6CbwVebfuT1v3KUybqeL0X7NlhOLgviPLxDPmPVy4isI2BQHHNvsvLkp
B0pTbVGdWVmQJkpnnmITzhU3bedvMxXBmyzdQUlkvFkONCH23SsnB48LTmegOw3l
HTqK4ufo4PFaMFaL/0yy9ods3Kgv+3LdTJLE6bJZzaJhI9f9pqWhLQmcP3ejwNqS
m3mrgoBrnt42NbbVqYXNk2rDv+9+PSKdmH+xgZCwVXc9iQ90ipwwcgzQstipM/96
T5R0tehG5SIccqanOWKvlfZJW2a81/nclUhktrpfiXP9Q9Yq0E0JRbqObx/oHVf2
GDY+AWyS7iQhv0Qw9t/k1YDV5ioeEE4dKQ3pYuyOG9XbRi+dAhWeIDpmm9UuO/FK
+I/GUeeuPkTkNtEiyBkeNgQsiLHKlj4sepH3Ze4Pydavx3Zv2cmZXbLiIeKWtofp
HwTIxwv3yECa8arFcv4+vsEjyF88v8OK1Vi/zOllzrUIlTOIyyg2mKjBvWGVuixe
WT9dsBaxKv+iaM/MUmRRwKyQvLu9S0OrQT8IZJ3l1rOgLKG9IX7/R7BmjiVVFIT1
IAhQXowibbPhl62IM3XxPnY95tFCUbVe+k17AtxT96TvID3wBuQXD5TIRUcafPZQ
DCY7IwDOv9IImomfEdXjosQzn24vJ9QAJE2yE7Fw9U0ygb+0628IbLWQduYgxDXU
SJjgaDi83sPh2BS1O5o+b7O19uR92ngRmoz9iMq8TsX8VBHuAXRZaunhjFg08qSB
GeWI7DXFhWReRm2Wcpx+1kPSsKFQXGQspI1FLt1fBsHmqro4BX/chSUrt2d+hXwN
xODqLhVRN/kR/yU6VWgnfXOzRlTpPkqMSoV69KcPhwuH62XB10k7hFdBiRslrT5A
9GbrBpv/0XIq/uv6zsPYZ9CtjEw+tzjZcMdrclMQWCTLbgR8ecSnI3duPrjKUGno
RoY3lU/V9JMPvlrkatZNgj+RPE2GOf4cvYTc9VXDh9gQixNf9jYcdNTBH2x0sB/Q
t8yQn4PiSlwiJ6Ly5lmNqBZmwVT+qwenDm34qhyC+oL0hkzDRLJMpGxaHzzPbU9x
QJF44k1ftyzTa7+hILgbSxD7qggOucwAbN2GprekOblGcEbVqKhm3PLjtJriKtXE
qbfA5CFJqHS3/3eR5CZdtCkwyPrrQzZN1RlN+G/1WELZArbpbmcdwDyTweXxm1d5
CZDZkvVuGWhcSkVHjd7+5wwFFBJDSzPQLy0/LfYlgJmVrW4ETg88dW4PfpA9x5ue
/dzfK+oDem0WLN/bIjjbgP0YxG2P15Iknz9pKgrGOfHdv6HUcyYzmTjG3OcAawCc
JTp4DcikQ7x9mfiqBfkkLRTOJKy6V6KTmr3FtyV6Dl9/TP6HEPIVsVLq9jwp+L7O
kH4OWuhGfuqEZorL4aF7MLY/dGe23vt9IG77lcai2EOEyw01XUYNRBCYzuKO1xA4
ixTnbDqo4PxNCwdETi/ZDlLXGmt8qFZACVFWf23X+xGsTE/iUcYIuMHNJdcr5M7p
YRrnstlQnhNBuq2W50X7NAWah4oqFrGXVzdh7IHQ8cPU6KYR6UlMsuaLM3/eCGum
TuUu+Dfxo2kEDfWcRJDNdlpGAfbDMIivu5T6whWoFWn72+PnAudVevqhEIppjEAR
RBEccIHplF3gHyIbjmGK6L9uG/Yb2ccLtNqDRTb3MvYAPUKlOlkjR/9Izy2f5/jJ
DmOojU8tvqEMFsItRoJW2Y501d/EhGeIO13xP9VVDClc8CB6ZuKxpgS3AmJnFqQQ
DWZJ7RMkbELtyjR5lcGbAYK1LJaX+SyNIDDKvJGeGj8XUJsWpvenhXbmbZVO9gwi
18l9/+dF0Qq35W/IlxMfkXRboSAkrl6zRm/NKuupJodkGWw7eB9FERdy2HB8kvFC
G5DUSxWTNONAFjVJeACvxa77dP8ZFIJ/BzjDSfmT18aNFLyJUuLN1RKMq7al7Eg3
kzF8SHNCoYkrC0Xu1v8KtnkX0E+oq1vN2fT2RCIPHsvqrevbdY6zMwV/NS3CCbl2
WTPj1+emlhOMby3L2kzQPxDePtEzY8OFRyxG2AexnARbgApeKV8Z7FkHDcfUHhhv
WBo7DwZ8LiLsuZayuMyo9LMjfIFAGM4JTF6QP5+Yp6kTeRHKFpMo9SWAk24krfvw
k+HN1lm5pIh4bA8NYKzjafIFbfar5pGkp2pDLIoe9lDOXq2JDXBSNXqBp1ePjoDD
kKUaHtHHrpI1YBja2t6POcba07fEW5sugonj8Gu2VcZb4LXtlIdOeamBXHnxUu9X
nVCC8DDLejePtfp+ROPQh/fzEs2YKJ2KvfCQMrd6O8KJWaXfIxk1pN6TONehKDgB
olCnzcQti2VLO/jsheRKRXWvG1cLh5UP2vuqbO7gedwwfeq7H1EOD2pEj58x4aB5
DCKYqvapfV6FsjV1G3SOjf68DL6jdGWXGgtD9yKsgYlJ2C84RWXwPv6tqTcaEeUf
oFU/czBl+zs/jhxqUU3JNSMN9yvzP6+Kk22kBTQGD9/bBoDp+IjnlA5mSF5x3ILX
tDMtefgdVtSwQuuTYvHlmmllpopksp+Ufs3LTdIr9lf8L46XrNTMF+DT0rJZmzkT
P4pCZ/HZOeXw+Fm8idHVFOxfVwsAr1bGaN7TtPtvtnT8kYsSrzKr5g7i1z3TGMbD
iZ3h1nuGwiBlNSVgVBn/sgN3WYnCbYjbKfeR3HDelYSvotiz2KbozX11HCAMNEqs
wHNS3tgTx45XZtEGipHFY+8Kfmoz2aaKDP6a5QFNhWgZCXdvfw4MUbOkXIeANTzR
wyB4O1fCWRv+AoRYx2+QUMJDffSwTnejQ1gYkZotcm4SKZ8+K8z+TaQ5WFLSUIUH
S/7mRAhsN3XL2sZ2iemY455hd1fS0yk183c1ZDWi9ad9q1lwr+Z0wtrMjcGqElcD
uNBYj0K6NGfPG24UyTaGzvKlxcDOWCPqqaZQltiOMTQ+/MiFKKjfeVvDSVnQr+iv
0QkscuMQ/4sKn0NOGhPXeu/MUv7WKXLWnX2fofcdLrZUZcu171eIYiWqd+CtoJJi
bbFA5BXDB0Isp+uD31GjrbYu+4FN4qdWzy3iBiVt5J5mm9pwgdn6pr9lLuiN/BiB
/hKxMAB+9Z3+IpGUYT8q4zx2W52fw0f2cJxupPKwLXl12+sokS6KuIPip5o7pNHB
lCAwuP2sgK0ZK5AjtrHysYFEYpAEuvdazrU7Osn6Obmcgzkh8twinnhl7DqYzvDp
Ps9EW/5cQ2fMrC6cTYNi9TxFiDgky9if1ajC9l72kL6ukvxngkNvVpKhwvJXULqB
5F9hFsDnF0GcALKfnjy53t80AUmEKERIFfY8NiM8LpcqaRJ8JSYiM/8dgSW058xo
ct34VKe8YJXIZd1X50vcFuTCoD7AGWVk51XzTBQCBvutSKCi3sfbRVBtSot2DOMD
sa+qIuVPieEbEbS2m6b8jQUVaJGB5zzojc5eoGl0GE8CoXHbLl4kbag3RqrEvjWc
6FUhnKU8Z7V6MB1b/JPg7/KQSqhYKbo1iCd0dnh1aJk3z9ERop77fLrRNEGLEsYT
TZ/t9jQ6qPoTrSFsVLg3hP1i6GOWza+A15X4M9R4CIroSWx3CBdZAe6bNBFnqCbu
IZZOeOxF8qO6vbZBW00CmRmfFPDmJA2vlk1VCckGIn3lnI0zMFZg+nIbnucGpnQ8
JGdNTfPgcsnK43pO583xJP1RmcTxaqIsWMffowQG517XSimfqNwpFf2ttyrDciQT
4JVtnOEWhklmXzztDduufGNWNRO1qFHWJOgGKRm10zHTtfZvDv+PY8+ejKwHPCls
kNAyvS8xo24vuIXo5FMf9i7jeKu9gSNCahbYCT14+Vuy5fh4PLpX9405Gi3fyOLw
1tvP6bJHzH+zznBA1rCk7Pci50aNGNdwWjyQ2tvbbvYhIUNHspR4oh9OpqjKVX5O
vwhRm8gKQO0uA22zfRRL7h9aXSbc/OCmB6rumRJ9TQXm9tufRwgQH3XwqzfimlM4
2v5TvJRnxk/fNfmC8sURLUfvdAag7+kLQpHYTsCuqDviahHtHkxbAxGrv+FQvsuf
h5vavCCTy3IqrvnwFHJbRC4a6YTsikYamSjkoIVlQaCXQd/weFii81UGEFfJBp0f
CX4pwgNFR+zc052/Xu2kcBBUjE+IS3TH2mOpnAwTVk+GrfQUih5on6aZEfmbrTV4
Gd2kfQOmis+BjIEE/PgQSYXog2Cgd558WOnbpK3ngEEnvfMu7VhKk6nj+ai8ywlE
M/68HZSC66rAf81P0zbzTlG2zrOxXiU7mv4QknbuuKCyMdvxF8I4gAwunsdQj5qJ
ZU+mFvBWX/qvsvVouI/WrqE06mYIgsGzAtY1FWTpUXQ0kDIw1J84+23tfjEh//Id
6epAnVgEcWf2gH19WgZKddySQQO0vJfVKV3kd9DiW5hY2gvVT645ntNIIB7oj+Lo
biBDM0hWbHBi+gjK4cHKlOZ/5W4tfqi4/mECBrFcZq2VPkoZYvGyo0L00EqZJLZq
bjc5Zs5QNFPxWXL5ykk4s1i9B/v5SEJ7u314ojzJrk87SQzDLKH39cKZoO+I6uQG
IsFiMX088dJp6llapHIP0JfrYGTBN7rEwkYkU9gAkOSDDnW9rpkrtFEclSBAg9m7
K0jZvsbHdqM+sj4ARqLjueD1+03jzKVHGMgEkWcpPYCslhGw/LJAuNi7yeGcDqoI
RvRY/6fM9s0zCjkl7QT1FVS7L9ivRVXgsv9hKV0/zFUE9j8le7zt2M8zSOjmwyDq
rQhWGUOR3QPWKzM9fM7ll50IDB+sfD/pWiIRwOywoUT/l3xusLGzQHiRwpATowk4
3w2i15rPv0yzoFwe5LaXuehxHjs7R3dKQZlJBMEgAEOwQE5P5gvQ3AfPZIN8a77v
1TdMVLtt1H9SipIP/Vqe11RoK8aXEoFuZLyYK83E2OpOQsZmOYJVOhDzoZYOKsQi
t95BqYbhRRH+QKnpUrwd3NSO84YR5UysyM0zTm8sLQTV8VpwI4WH9QWwuXjIvgKU
Z9CapeI18efikoxlosqDgjFASPwzDlwtguq9Zp2gMxjEZokVj3CAEUfah37FcyI4
SxCr78R1Wdl0unIPzC9NbkL5C6DSyYA1WsDHHcQ7U82ZX5FOMfvRLYR7Cj/eW8XL
WSpcnGHLsbmAovGDgM4dhThF4U6yaLIioyMyEmbQ+FQECm+N1+rR3Xi1jhLAuw+U
NgAuU8ZbdBE2+kXh6+Oe6EvfPLk1+fKjo61BK1D03wh2EYy6dns91jFYCc/hZD24
QisekFVuacD8ZKNH8Szd87TO49ZL1DNeWwSNkQkC4kDz7oCsYMFIFI+k/P4LAmXW
+qHwYNbZjOpLcMQKHqWmucvBSXTl7H1nciuwBZo497EWqu+lO8ZmJIcjp+vgXC/L
6m35AA0TJy5a7nXEh/TvalYdeOK+mk5psDIuNtA7O7gkn+B6y8aHKYBcrFVKB+oj
0GKNrKqWB/N5ISdj7vTLZFWATqXabwJHBXX4zX8x4bFBjhks4UXHhdavbIvkLjDQ
YaHXgOa8c6+Qb1gSESjUa2aBaqUMjgLc4zqtOzZV1MytTJYGYr4p9BgsDdKmyi8S
oa+H2HrnqsIbiauyIyjuRkSEVaQHZugU6/o3MjeQl6oXffTBa6teo2z90qd6Il+J
/1x79Pr+WHLXdx5meSyl6RCc4NHD9Jv24xYfvvfvv3Bl3li0GNFl2D81AqbxuxmX
ZV05hP4+RX+uucbTkPI0z/ma20ae5DsggmPJPjWhy/qreDORqGlwDDW2qk4cWFTT
rIOaQucHyR9TG4zS6uFBczrHL4aG7K/yoOtGnm33MtMVoegbktomHDUnfDZKbBdn
0F6xiGFO/fL42XV9nbFR4KgMHRCzFpGsGWEdQ1Y54N2YPOel/DGNPfVktwPA6xcB
5en3H2h0cqhmv7cLKJvHyaTIKy0WX4NI7bWuEx2c0mHVC41bBKO7M1+s7pPCOfMh
pY71cByC40Idde87ZZ40xaBSocqDbaYFTezV1683gqMu/7Ph1I0fWSTeobj12Csm
N5r1GifqnuS1/IVBZJYSre3gSz09jl9Nl8N8WrXaO9LbXP9Y5drLUgx0JaQG+px3
vODwXh5mCiMWtg0VCB9oIh0JUOOxDN5fmYAw/MZPcoLuOZVdBB8G6rRXWaqojoT1
oT3Q93QSUF+13xoCx8vn0bp0RpcW9zcbdkfdI4HftPB502wkyIF+Fj51acHSekW7
kHnGzOJLwrzcmRV6cON6sEwwBMDoUa5ifb78GrNiZWGjIklZGTxWtPsSqJHlZyUB
gj+3llTc0lT72OSE2dwM+5qOuAjV0I+FBiN+xBZQGk18AA0xJXkuMM4HKKKCwzAn
6MeqPKntZI1oOptauS4CdGn5Ud1M/vbnjChFnIXpMXYIJ5ft2QouEFV9f1MImaJe
c4+D28oY26SrRbPShr6IKCZ1D2kqTvRt9r1FBxBw7yghkl83AZyVA+pKX1R6lIdn
aHYvFd/uqes1KWbxEartR8Y37IK+zH7U61eaIv/a93w+gDrcL/z+6vEwUZRgWBw+
39qc5ubrpCRr4ay/BxCDpUlboe+QbMEShtuCVpkrZDAp1UCckdSNzZ7Jqc/uczAU
Wwqa/HevNILptdAmCPyqLd6NyktJiuth8Wj2ZF013fjtBBgXy43brXkGIwhuBi3s
x9loEHbDltF+t39aZl+g0N1Qbku5+Ajwsjj5nRM40b5Rhl5i9pNvCfCfDYgUW7zz
TXutRXqsCH2YW/xWmKs2eGWAmFSl4BdzwOpEZC++0nAVyD7d5w2kvxsosF/zUqxs
6ljhF/8dOxCoFJzKBQCigrMs+58IoWMoxjlNaLRSSvtIZ8yI4DtoO6Qi9/nYo99o
7G4iN3PA2HwIS/wlL5x0S9++71b1a9fDaJDlMa8W+D5axk2XCbGQZfFLz0HGtLBe
37dPCNN6Jc0mUwC1btyo68mCCLcD1kp00sYicOpr/JcFxrBZWpCRoGDlDe33gfmX
aift1ggmfMYuj98SKIQH6nqBNJQtn+iox2u5muFeyoOvvPqnjJ/9ODwpzAzBoKaE
afScwg9PXvk519GaGrn0fQ3NiA/WbnIydeuHgggZ/OZ2VTHyWejaU6jEFiikjyEe
xSXpIkZ/h09zzxROvqpov64dYZj570vbyNCshFk4DzGWnYPsWz/gzo/m1iyUDzSL
E7+S0GSLDh8qEK9xq/CSyw2KFlYhJCbOJKN2ODhjlJ5pkgXeaXYWSCMq0ow7a2vs
46F261MSui3BC2pgsfD6h44cQHaw5+tgY4qqUzOoYC4lejg8TAxnQGqkz+sJfG4v
paJ934LeJ0pKULKp1YX3PgQq0nc3A7/BhB/xv9NgTmL/NrRRU3/uDPceTfqJqRA6
CcyVrR7PeX+5i03OUqNnIuzbT2Xxc9/YU69H+vNs8aUlegp1ROw07WlSiNYe9YQB
bRjAtw8APR0lGJSKUQwT+eCmQt1b9OvXKF38yj3J+2YQaYG6peYBVu3G0iSHUKyt
kPeFn1/CboOnzB4DZUo6a/EPqduhx/UMC1onGJ/FGA+i9Uug/evS1hCo94lS0zv3
Ew/cSV0/2N645utyha/09XENHId5rOLO+McflED0h9pj/SaH0rhrESzvd6jPvnSS
mDAUixvnM++4iwBphAsda0AQTvuDJLYRYchm604nHerqqgnGxE+GCjjle0QfW7c2
2FUYTxeT1n8STBsNUX/nfft9Stlj7bzGflQgaVQNymQCN8P+ZihorDXFZLDGi6BL
EgWIgIDWChYLjEYBQz+UxXqZ6O8lNwSu0dcmK8ViihcgHceLJnEa+Gmfwlf7z4el
MV4Uv+ubNcE2/WFbp9XTPwOUPKQUPfZgJmvPVrsIycbmJvV9w1CfVFMVlo2s26+p
8xjOJlVLx8mj3aQXb1OFiNDq5cPGiqvPdBaes2VtMbAUQJD70dTWwnlx6ePQTrdA
nSPdlZRLrNuyIY6WmJkivinrpjv4oNUHPxEPffaAXvPcg9bJRjxbvtK1cIGH52tJ
dh+/llDmHkSe2z/IBsy2xsdQqiUMETj9SCUyrtznrcsyUOakmShoRUqJL5bBb02D
Uqo5PqSEuACMvvIow93xVAKGlsff9DlnbH4SYJ5K9usSyJR+1/HyO0EW9n6qOuTV
mvdjqgSD0BRNvqDEbaf9AOmi2CrpKACQr9PWHKklm7b9X2OPGAOePUg0bY53jwe7
wxYHWyl+nJqRK4OF4tiswynejob/sUzl70fAqQz1OTKJu0oPTGq/mkZQMkDuKoyE
dFbAHTqc1xi1bHnbZzHcn9aZGs1H2vbBxYrpg04dPZ2jtmcQrWO4aRtNsEY2wuKI
7JZrt0Z4minTlsmYJyVPu5ejiRkZwVyYl7NqomDFmaLqfFGoiizrkJDHxB6BPKf5
bpe3RtNbZkgvSmGyYw4NCEiE4cZmvZzyB4K88cguJwDMPYrdRwUEbM2rOQgk4IXn
ubLHA/9Civ/G9OJbZJyOwi0hrL16IZDMj0fQhSIsPG4NMLaZjtF1HX6W+K7gXIs8
MtNm1dwTj+IYsxMG4RfA0wwC0pFFnIHhBj149b4Y2XgEROHJEUxQIoHUAhKlaaJ/
DZUFzmyum2liapyn2W/39zYn0IS3+LnsRe2OuJGtFGzkKciOKL7Igh4CHo5sDEX+
aqUbY1K5TCURrxOBEDqAm9ArWXbDnSQQxlhdWt7HcrJPF0TNl6YRXEeW1H/tU0Ef
pYj/BNY2yZjFjcPyZpmwz0cbNO6SyvJdA25kV6t/0j/pUKvWpXrAp7z4aRHCWsMW
3HE+ZM0r7zlm1IsIe/TvjJ6NA+pa+2C3SJcIFp0/FgUqqiIgbQVTKOxPhsJKpuzE
OW8hdPJLhWgH5vhLbraPzMbGOgK6CYIcRtzc0F1NqfVfZ0dPQ7kmxF3sfRZuvjHv
VkYp/LqVFLBBac9dICbzrrmylytjH1lbKoFt02/Nahgq4HWwt2/tYC7UuGZwyQoa
nG3Nl3FEFaA2r5HpQxpJiWQ0kBmKVTNeXl3yhPNYMAlYXRw+ZsjrMX0NKQ6iPcxO
d7z7BNsRB3gblQkmPxhxJ/LXILR56GCfpF5wyYleHAFfoQV7kLo4mbsevAGEJGSM
4tB6k0Eh31QX2f1JISx9KVHdha/YOPy/XvhUCzGB9YTTsLppIoLq7y9I8zaGmuAs
3ojPgZ3FdcD2UBkeC1xdrRJgXPn/jRrk81EAFhpAPgbfHlEPgHgUdGwiLDme4RjH
nj6nyy2a+QHtOWpqAsTpnd2tAe6auzc7G/dwLmrHUpEa1MKVraQzs+SQt3Tk/nS2
B4MyEqotAWk0/goFr1515BOObnD0rCGQV7I6IQzx+5VCuFR9bu4rytWXrRhlyOrx
aTdMAPRsthEoU+imMsYNxVbuHFpremOjJkHb8exSweZ/kf9Mzicsjxab5h0JcSl8
/9FgIc/W8Fg1iZBKdxEltp9D6rlLVBz8eOrYfS69ShXw+Ph9NCVTzxFEnnc9hQmA
eZtYjHvg5C+ZMePd1rqNbxZ+0LGQkwOV3AYHf4pXaxsZJOOmoyxVgtBoFFh4piwW
+kcXY82JyXzn/+CGIU1mnCVFm1zMKEc+DKMDDI37b1unNmD23CW/n5rIEMraHnxx
LhOdIJzmZQp0pUcvUPpMiDoyr/GiY92LM3ModMYfET9NLjObBn0fVx6Z/IpVFAKq
MQweSMHIWpvkLQxsk32JGmL4ek/0FT6zf3aYlNnZpn0/g/xN0O8L1v3V9ACad/Y8
2a4tpM1T4QPCu8pTHtmvNGtybFN28TnaFjagUuM9yVGTKuDaakjNNEZNFnY339l0
wlR+F+Pd02BSPfjBBUHZkFidRtlSi/KXIzmllOpbdZVssYb2WzAdZEThpOoiauyi
nMkphux3DVwAtDnfOt+wSfi3MuMY15gCgLKcnvANDu2FJ64gQiv0kNVvmlrm7XyL
ugPqc1q75HlbI+8CyWt46wVMImhEw1nzOvolkPoWcBDSOK3O61jDB/eyqs5tpwnN
TDJPU4BL9AuwNghP3ZhtiVjFZ/mOiVA2lPb1wopiXx0JFAMBjp3TLuTWsuRh5HcM
+CvdTN+52/MEe819pFlJaVgPBXBrt4w5AQReBuve099JYTm3TXKBjkofqWLwhu/f
23etRrZvrkBP36qHbOGwAXwOJaKh4QzZbZ20G67q7/kFALCj6JFAhCOTYS4WoGr/
JAjhYxth9Xx0xZO98YqWBwbRHDGANI632nESyH3aVtrX+aU2FfCBwIZsgs8ZoaRo
RWKkziWIhFDbQnV/JSLeYBKTPW7Iz/JjQZkvGUBDxBkhwIy2sxq9jqjq0CciPXoL
FTs0fl7qwiyL/tmNe9nd2nfpt53FHvj2NhZhLUM29y2WrkdsLiDIEY3GplNjwRBD
vvmPnv8eA0SdKS2Uv2B3C+nbIqfVFtlLJkWVmvXoJ7126SPHyGR5WzMedpqy0sW7
ZcbG8VrlXi+gGE0Ao09zhR0za9wRlZ8PgCGSNZXpe7PythcQLPX0ROO7Drpo61Hj
7d0NgrU/ARS1cG3kKG0fcomhYeKe/Q9QL5tL2lsfniXrholKMLe8fwM2BNdKAQlh
2DOKeJoOe9hj/UEAbaahTYeAXaRplKxwDTZ947Y3/4DdC7moohgES8hm3NLnOLqj
bRADzzvPyYMbvbPW1N890TadrxmC5+z+qQtngj3pakpfhI6KMGgY+hR6iVyGnV2x
pkwThvYh9xm3eycwXD1bqdwY5+hig7pLpJObO+JxtM4dWbg8rZuVKJsFFfCdeYH9
1oxTZ849WUKY+ejT/odUm5E0PxHezAWiLe64+88SgXiIeE+lwMxMlVEyzmWJyjlT
G7Op4DnRGpyExygL7GC0eqfWUdEl+rq5TlvEvwWDDmtFwsWWGSqpNstZxbWEJurF
5HSTgxpHUmxjRm1rjDRxO5za2z6EYTZknq+wuMxal7nIoUSX0Nozus1ppJSVcBwr
z9+RGq1BON0ZE3sECq4gILCTsxJwt+C3MGvm7MvDbIJv9YqDgLFSdoiymklXS6xB
glZYuP56MmlwrYyHWPUcGOUmddov4Vz/R34vIKWnWMkfFk/BsgDsgISdlBi0dgAc
PrNVb8Iy3PyftFiugnSKLB68E+99ZguabBj2MnsOvZsveO2es1qkPAea18U2xnVf
+62HvQFabww/ub8ZqFdrchTQF+aaz6S6Y5InuIzmViZrAyLg6rNLYfDnvTqcCEop
JnuyHzOmZCQdsRkysadroTVUnwJA1BwIOoz5OwUcoE1IWwTGVsGTd9W4A1J9IjTX
kIvnIeeIFgf3ebBt5Y9kL3PrpN0pO9PGw05gnni16ybRdl0hZ91IXq+k26vHmnQ6
IaHCgtOSXz23Sdz4JpgEUsnIv0GxgSi0JWPBSvkj0E5ez1B1+U2EKvMKlKG/1qRP
9ZSBMJEkqSn/WL054e7e0y9d3YmeKf+cod9PGrAYDzV5lU44l6i9WrvJqhKcRIKA
sbbuY6RfldU4Vd0GaH+ZS4VtPgoqeQsKZ5nOHjagtKfNwgV9L+ESjOu8qvXYQhfP
ajx8MacZmg3v+fEU8T3eQyecdMdvOJ9alGfGS+aNF0aptU0daYxwDEx990vqwAPR
lZ4/U3VQ2I4jKZ853mw18z3XrGHqph+1ktna64UCUHrOe/QF1/MmHeWtapEh10aQ
s0ZT0TeldgWKTaJjhBEJn1jghnlH0hYTZz+uPuBnZNLT8eRp3IiBC/bXOeKKedVt
3j6hCEWXz1dMs2I6esLjcaHRudP/BpgrR7sdTAAZ3hGuePpjUiOcIcH7xDqnpvCt
NJeRLRZZCS3uh2XZyEmBej96hGC2PbVlZdpEHbBrWl4rgI/jyD9Uuz/42eB6twfO
oq4c/xi4F0RlIZRVd9tVjNR+S8hcuxgI+QZOaRsdZVEf7iuB/zqaa3LQAV2DmIiZ
5ycclggViOrI6grDpfEenPNnFnLfRszUDJmon0j/8gPm5L6875tDwH62ZQEmGniW
4W8+PomLp6sja+Kgnr3Me+VBH75VnQuJA0U2lBvg1R8e+1nq3u1M4oioFuEc0ugn
pqQK+4b5rWlFcO1mYeGpyXe+T3FPSbbfAtVyM5RL0l0/K1e10iLdOcSQLX4xCYv0
jJpSaVZmqCovs8+axbfVnrmO5r4KxLMJBRTWnnBUYxcNhqwVh4Lp8q37DCCR/Oj5
3+iFbMxaFnECooQ/CXdhMpsHSpYoNm+pv43ikIiRSfDzR2kSVrD7JttkJwNbYrdg
9nwtdjwLHcNc1RDSZB/EVYjbm7dYJn78w577YIDOsB7pbL83oPWcqYQue52DXRiy
9hex77+1xoIkKN62sCX8QCn7yY26e0KLEtNH/JVdgNM2d+VXDl+9qAnoetSQXKRf
e1vryIwdixZ6ig3FPBYIvJtsjC2IRGKworTlG2B+cMfFym6pGJuZbBJ8zebn71l2
piWsiFYpzDGBRbwC1PHtOhCvlOJTe/cwNWXyxbZ2j50pyF7WHTqvAJ8YOuFjmY3N
lHjyscKx9H6Che39X0LVdANraVb+Q9Gl1IqsxltKSkuvTBTv8W5GKWcY0WuMdUbh
Fwg+MpeBamA/L7RGZvxR4Tuv5cz+viclGy01dbDzSKxI2nQlywINGvhowIS2g0/e
jeEaXl/+lgBzVI5lGtM9F28srCkioVpvQntik5B7BzqaXPK3Toqpjxdl17KZf7gF
NLJJ0i6Aaw436AZbyCL33TrsAN9xiEHZYLvkkeZtxS3pGre0Ty/Lo1OBG4kA4IDi
lTX3k1gREfhDtsUX4bMJdqFK+MepGrKaxTE1m0rCn182aIvw3hgZK5mOZCceei6E
jSth7FujFibibvPTiU+0AVgOFCBpk7JQApj2DZT96ZdFiG0xGUEJcdNRJyUxrq6l
UmYMhC1f584rz90nHllHX3/zH0+vHMZ1t5YpXejx8twYSxAGK3rNJ9tMrLEiMFpE
nxaOB8LHEJ5fEaRujhvXBQa+w8w1pvRAKEq9cRNs+ZsTohvQkBzDOr7EEG+ZXbyD
Ti9tzYVSNVFr4ZPUx+e550kGJd2piEop7WyRb2AxNvSyNcCys5aj1Z+rqKtBizlp
0WlfjJywXgzYT7CRNoiRObTbAieQIOMhpxYyYeTeBiGMGWwguGBbbU8S/vligI6z
bdFGY9dFPRTRldUMVi2myXIVZ+rLjS69nuAq6RxGDGnwiBgteEztW3XZh8jir5uq
Dvhr9GmeM9INjuqZ1aOXPFpQrAxMBhhddbA78Ka6sGPOW/yHr1o165NyeHpLSVxn
qlN8YE3XQRCkw2Ok0UPlNCXI8EWmcVfEfCMx1DPL1e+9tsnh7XWpud115TITicdB
CDPJOeEjTsav3aj37vtPRlIPlKjWajb3l6wlAo/2Xs9MpTXZsA2MsPUgsdw3oOE7
kDx52ZkypubCT+3RK+c/4vAFriMLrzCaEg1tbwSp3no6dFivhIBJ9nzv1jEWUD5T
1XNsYlXCDn3p8lhlWVFOn4kM9VlXSBhnKNCPoKp5NKMWE6stFMEdYN970C8uwVKP
s3yqibfN7pBAot/Y6u9i+4WmaDDDAUGpLRzD2TbefAW3QazrNHr/rLrmVbizledC
oL6xDQBZlfIjY4GcrJbWnyHLbtA8THFxE1hh89/AszhRLP4iug6Yr51RWEubZ5xa
vh1oLfY+eImqklaq4VNe+7Yi09sOi56U+V2AeFG0b4WUDEhly3ymoIsUfd2yfXPx
KXLmwnA4BLfoJT+dKfoPMtTE0ka5DqRtd9coy9Y/eYO0Vj+V559ReFYUYSmB6xaM
rkq5UPeL08gREgzKokC46EuruTxHo6FNKb9zg/pqAtvWd5/GA2puat0kddArRl6Z
6kKqZI+AD3BAGU09INYPHKWwGK6BElKtaf2Lpbiq1OmbrlVRuj5k6ODxegiTOBv3
DJLzrr0bSV2GA773L6sW1pI0FZiww/L0kWKmbRY919OVB/F9t4lc0gH3gpYAFA8V
nMKEvr41kI20KaSeTvWWVbD6pS8E43LXMMnpSi2Y/wsK6ozacpSTYTkRdcp30Aet
9FDwiRQG0qgeHnaXDP90PXERzSA7pXELdtCGf3Doy7ZPCwBhYq/jp1H1F9B7/F0v
J6k1bPiKOX5mYUSiHMi4K6ngb0wpe57xoZoWe0V77DSico9Qu4cAd17kJ5JIuKv7
NXTbXjnARWnuzfJcILHDjr17GfjAybSx4vlR2a0QCAMLXrDPmtRMWW4R4fVH4uQk
fxE/AZQpDTTBSTmRmxjV5Ut4CZ9+oFcJZFzdeGlY4hJ2juEb1qg0tknHpv8857h2
XWKuDeW3JT5RK1Wnk41RYVv33qmuFxWZePeTTu7Bv47juzxg7Wfhmoi7JDbp21i2
jHtONAVCsKUTFanWH/3qZCr1+jA1/wetjCBHm6I/SF7fR3Jwhmep0hG9RDpNmi5c
I/o/c4a1IKSjEsa3pQ1x0pebvXtYXywOa2vPtj2z4J6+cHAhXAuiOUPZd9W+awMm
ZF8WHwmVWsDcv+wxCNMGd+zYBdVDR7NeQ+w1OH3cmDlY2aIPa4vsAJadc4oB7Ibo
BK/0OFjSnhkIc4LC3khr7/QNCjgGNhiYEpGlFUlBdBhkMCHYZg1So6iULT/RoNH8
Kf54DpCq4zaLgwJ/t1yrD4X1w3zK/sQLmLgwV4wrx/v2NZhDK4E8pgl4z+GrpOBt
cjWNXyaKCrm731Omr09ygsQDdcdtjuzzOaYGCDrIDbSWsU0FX0ecBpjcJFl/zsDE
aANBaQyUjhWugmg9ISMBunlYxRiW8xzwFtf+FC59iwkCB3TNLn42CmB6A19+gG2y
ucWlli8UJG3ROCdzfpeY0dTZ/Hrf1wfCU851OiJ4jhc1+a4iWfYoxsJbUH5+8G5l
mMi0ZoS9YCinfSzBJignE5vkxFJcH/z1KkLZzHftGuj3aEuiUZJpoY4ja4g80NGf
q3W18cETfukvEWwS9UTGf+wVesilDcaRRm6wsweLj3hs+T7vw1NywK2Fz3rccxq0
LFff2fwXuhCiSDR99F7LKRlNcYc5IL3nG5Zu23yVC4oKvrgdG7YdgyPdDajPzczk
Z7UOaYFmgbEeiE82vCRYPRWzNpj9uTrMWE3juE8TluHed8RB2Y/c7NOpxBUKvmwQ
MdbOi6VpL+SEZbxMItpcSvB+beA8NAZBjqH+QOG7Ovseq9Ig95lL1DfkebjLQF91
uFC8xo1Sv9gQsXFnE/CkEYViN3EeIv2QyaNEMPhV3/7wUyZ8XhIL+R0VKTS+t/Hv
LS4ZD7YdfLnYiG8f4RYa06W085gYBIz9U02oNzqDzLvItldE6YUhGVZboJd/cXGD
6EdaiV5CUiQtK5etnW9yHHq4t1CyWofxKTeGaqdCh41eWHJv9Ray/cJEo6dq0L2t
eb8BXyhdS+z8ubDC4RsiFRgtEOu+oyW8GUWLbATvXuEJ8enNU7NZ6ouhW6xUa7j7
N3VqfPu2jTng8GWWUm4agfLuZsEwFfI1y74AXw+WTyKFf6LVK2kBjra7WpZlSip+
9vWVLJyaMY91C4GvjZx8Jbfbc6u/M1Aoy9t37ofYq+WiU2fLWzgIdWCTQ2MLACV2
U0bA5Cx2rvNLZUtxYTL8sOpnaSLLzMDDHG2IL1IEegX/h2y4Vwc2wmR/465wAz5s
MApvDd0LTAwAH2Lr5HMVDCfZkBSpS/iHJJpkO4Q5Mp7fS5VwpZNCDIhb9d+XUI6K
hX1BJKIcwxNa3js4M/p0erUg0FwVKK2Sr0/TWArFYYQZekF4Z6fQBEj1Jl1A/ke6
x+FpsuOrIqM42oLk9atXRJFLkv8/ocB5KHzoDrLThzkLLr/MXQ2sXgGwIwslPQUv
mJK+lep/YE1T8g3CaKUJ0ICggKBLcCB0RC4cEI20dB5q58bDojy0VOsVk0QG+iOp
7JSOpanWvCQlByx0OlHH27TMW75IXbMN71neBD5qEcAarqpUkxlalR32z09RgtWE
Pt93V5LR62txaEATrECL42BdO1cEH8pNlNmlUqqH4MHxNekg1GcRJhiafVFymn5H
A+Gesh62kEOfwKwFPk1+LjTtgymUzS0q8YRRq1bnVl9UBKbc3VEsIl29xRrFEv6u
ZoKQJFdh+SmyZCfDSNKiuCFRnmzlUDAWQT8PMHQWph6AVBlu0vefZ3J3MuhCNMOg
Ul4ouwcNrE5WKHJj8YStXN/TAA61fyqIryChRWc8+8DoPF48KrSCpKl5xIXgfSok
FXVweg/IayHn+GtAVDM5fUzluTrDrnwucQkZoUGbfqMJHo9a0jcRfKXQPjB27e3F
5WPl2wOPCpvdu5qTBNZzYXMJ0lEYyS9ykkeGRjbfgAt7Xy6cI1jRmLjUsvRvt2GY
PwQ7hhDrkaPvuWIEEy5lDf9AQRWCin2adXQx17MkO9Mk6+iUwbUc60gmrKFdbJEw
stf+dr5BxjBGhDsONlNZtxVDsA5lVnnYchLBUt0oezD8cHlVdpofb0DIunTAD1GO
Un2a0Tdyg5WJ0tq5q8VLhtVmCZx2/eeoi2d6T96RxHKXM/vPPX6ol/au/qgvdl0G
EOk50NMOBo3kveEzO3NSwgN6leJhjOmnb1r1pLF4zWQbzoiEe/serhwV8o6/jVbB
CyuSpRSBWxbJbowCuwOc/uUaN1QCrEznrbSoaXUTOhmeEkBpotT5hWTLvkNAi7CK
UBphZYnEoZvz6lae6R1dMmzwQLfKgrViDbcS9XBxjkntVZxGTfKVfVav6dPJHW8v
wIZF03ljFQP9Eu4TofO2SEOG/S5ipNW8/z5ppGfEP/9Otq332RPZBHKRshuqtfYT
bkK6jbdD2f/Cd4ipN7RHMVQq8GXWYZDu+gOx5PZAtJbbw7ETa6f5XvB3L8inpFnM
YCcceCCqw4TTnELPeiXs0jbXvDl7BwEI7LRfxiWOis8t8ruwtNLd3QRBfvubqdH6
PB2akjXi0tS6ADa5jWs3O5BnXMNQa6CjYCD8QMCorB+hBZ6kzl73Hulf/7987I+R
YbTfG9OehYC/GOL4vkZ2UrItroEP4k44MmvfJK57ZY+8mDsOvuBFEB1qihXXwVpR
7eGdB4eItRBve599u3NF5M7Ms5n9kO6DOHL1XHvBimTnjogUf8QwYVg/6RNMq09A
0HMyaVtZTL31xRSkBFSOPHYyXULC3jZe+vS+ggj+oCT3PrBfzsBjgyh0wNQfuKoq
KnLJz0akFbJ+LtnkwOGoVqRp2v4wQFuahMe38lj0gi8hgR4THUCNl3+5Wd56gS8+
bYpajZJag/NcNpShaRk/nqPEQYMmz5tQ4Wd9C8+zaDoXnCekBP6vL3l4YTbHyDRu
7K+4ZAmmvbWQUXXgIyVgjBrm87a+Boq1DITXxmbKw0f4h5rUkQJbH/J+CrMNA+dg
4bpU5Qvt2lTIBLbX0umpNlxuDgS3qe63paScn4LOgP2h7XFfFgpA4AndD3G8f6kn
9VTQ0dGPRJGV6xVdWjxsapiVJTLqfZvJ6xrm+2BsGoUd3++QwkH5HQbq9gSUs2cC
S2Ih77NhevGxPWPWaX0/gOHeWKpRTRpLU4FLeqEeTDw/e7j1SBl5SsIgBCQYla/k
6+V8uiQvUD4roPAqD2KiTHRZpBE1D//xo+qUYM2BlTXyBSfcbYElbBeTdkk8E7zB
1KGZ3EXyymGk2IAIyfa84naKayZy/gIwa3gApJqYSyOgYkoR4Tw4eCALMaZ661rt
w50nWVmM22f/VLGuYbKpEm2e38KEc6fnr9hy7x/a+GtE3eF8AGdTyGCwS6Zi3ybK
SAd6JQ24sqHovRw8sGkyjSiEVpf0wNxD4yRukXC08i+pZHNN+pbbpsgMwAyEk8q7
a2ihhay308KlhmNYmj5MZ4fWCxqRnFGqg175QH1FQd+haEhVn6GD/RDaUdL82fuh
2GhbS9jRwHulFr3zFriZN7DFChzo5yCh5YmGipKUofdyGSqJL1ON9K6Ke0t8MXXF
WcyDdQ2w4DZor9XFzYIlrLjP1Ji/bg7+IPmHQrgijvVI+N2UZDPpC88ccbb3LD4r
9R8Nd+TRc19L3uBlFDt+dj5kDXGr9x7megqtAkx+8XM+MU38o+5VxJRVg0DgNArS
EPbxrIDiJzHnZrasDQ5f+CW1bUlmWVJBaUcznTs6+4k630Wom13SXtIMq1g7Z9CC
X+1u/3RAxWd13wzaVFbs1gej4Ioz9Ub9DHb5RW6jOnL0hnJmqi4Ihu1bj0BAFyF3
J/ULHQ0eavNWa/k+3gNSrUmFfzTwJQp7Hb4YYuR/zSHMz1o5o6/KMoNLOhWyPnn3
OWqRmfLFErscVA/hkHc7/L7SdSi4ZDiEcpMiGp3wCQc4p2PNImALuoDh6TcvJQVR
7roVZx0r/UgrclUeS3CporYrVVSxdxSx5vugClUkXTe6HHGsK+bBCpihYYbATYFf
+YOuJ3FjLLTMJbrbwlXafBZlPW7WgBcOO8LhFRMp0d/mMHowXA/MyibCU9Yfxl6B
AGAuNprH3MHjj1lOP8/jOyEPJeNZ7YOHf/D8TSswcpC/6N0xJhOw9hZjn1U1N5PL
2CPc7vgswLC15eNIQZVFOs4HAE6VOu7GohIEFoT/HkfG9MH9k0P3vBmJXcboh2pX
k/lMJILIiG2TV8kFYejeH0j5AGQ+v13x0xI97iPJpMSIPewmrjQBMz8DooLSluZP
nRCq15W88vUQKaL+q+e25eVEvpoHELnM46w8qoQXnOPBE7oOuCx6U95O5pusOunm
b7rDvFbjD8dxinNFf6/BWHbRPgCb5gmr5i8ZH0COYmmcCW9Q9w61EfHLLEkqotpt
idYPmURBqv8WJrMwL9Ib+ILOo9jI3366hAqZQjPghCi4zkFTqfT7DzsqHK6CI8aV
jJb3BMhMIEwgS4qpK+Em0TciNVPv6LheHgOLhJVLK48LlDMPzVJ4zcrgls3tmfGh
VO+CigOTUp0N+jVZlzJyerqbFGEQpOsHTTGeC117N9nmC7LPp7gQBQAGMMM5O+dI
3Eqc4K0/DduaQlWFYLCjz8qSHGXje4Sc/bvIdB7/4SbgWiwcMWTF9SwBtUYKSpiL
9Jl7MVCIo5mDJbk0o1cpY1jh7MpZ3jwvRqJUUYsVEMLy5CpN2mGggv49dZ5yRHNy
2NV6Kav0lU4YTfOHTBJ06kRDwIkml7TsOpq1qD3jFQ+zXtJtNYy0hnXj+0k9WR/r
P4BLGxUvgZ25QGvslUOFdquu5bgXb5zZR4CyCwz7ODuXNU/4GXrZ08ihiYMTYcu/
kzgAY9KmvH6WYQTSNFhb6af0b7+FmgmTIp9iaeA/sj+xTr0yJOoE/MpYwQn+jgg3
kU3P/idmfBD+8hHTKDBBcoBonKt6VfbpmPCILwa57qaJCnErwEFVw7tNWZnRV+Ug
zw/tO7Hz3wPeT5MGnDRcmYdjhlvFw7vjEqgN44yaqZNlPS1+rm3TRp2STHCJKaSS
jw2vzwTYd1OR+N5t3+jFBG04/w9jj9PvdihHwWMHKHwXrm68f9QcNlal9oWx5aPi
8N7MPaHM+43b/K3kd0TsnTYZHJNjSq9Y2T7VkQ3FoalJcVgFBzy6ygD0Pr06Xj3S
L5RPby3CIvcbgV6dm3kgmutqUBb08ekv+rX4RMstksOGWJSRyHePrr0TsAWrTgOj
q24eIBMgXGrqzJUC6B9zhFfQyY0PZEJcWElFXeDOwxTqSyLadsvYKN0OyHk+qP0L
EYXs4IjqOEaMTbhBrrD2V1IqUwb+Wv5atMc9VgUfrTE9buRZDszi9bciYGQ5l06k
F7alObYLGblgCj37LW3DGmsKeKNDPp2mw+G3k+5C63newy4kGwyr5N65r/Cl2e2t
+glDZnTWm8qMdPTOQa09LFmqn5rTDZF4LHRGJ88RukIJWlPpZ0+Qh+SAyhBb9CY/
JFwwsw068La5bWDQJU1M96jvKMudcXUQUvaPeO03afr1LIfVm4CRv96fJfb6eKPg
l0s3zx4iP+Gb6nK2tPcWdHENmpqLhlifTxxh/x/gGN6w89gE2HEeVWmXGulXH0lS
nUvz+Xqj7NyOPeRnm7RcBeKYkR/7npMSwup75GUH7aCkNlKc4sB5h9J+cqyPBuH4
nW6HqRlb69tZMjAou8kkFb4CwJq+ShsDSlY3kbzhLm3P9yopXRpEtP04TbfUUITi
y6kFjc21nxFg1BLtH5DGwFC8ShGp/YvD2IhuCLAKvveEkCpE0kOtFQ+MW0ZZvKxQ
iRpfxiZvWAdEFvTcZGl5jj2cfGrvTpB5JSh/NXyxbLdd5rv2otM8z/tv2Hv7C9rg
wMhU1Zzzy/HKGlx49daC8twN4vf+OpLLV/fOKAuOaGnIOj+i0gfT7OYmxfFP8jeA
MWzhopA97vv4ZvnoEqOuIdPjUTOXDPNs3cw6MLBn1GnqaZ3AEI2AUJTOAZ+UmVgZ
Y5LN9PbrQiv3xVzAZBvhvBE2YrlHecQQDq6T9chlqhqs75ngRYmK7JBj05ysLLeB
zDrwPM+FaJc2GMCqWP2U3NYnKGk5lScFb0rN4yVYwIZxQ7MM+eFpTZd5FDJqaiIT
5noBTWLxyq+mfN/Guo1LrZICUenkKKkdzH29rXAmuf/g+Zm1gBnSEr4QzDLGJnLT
0bF8Bu8ChG4Aakprqxp88LddYlihgpKsBCqi3jxJwkfzufxmUaTBJYPklAgswayY
Uk9Ql0Id4e8GaDBm0kZ5/RkaXNTRTpNVXFh4hE7+V7qMSoySd3xXwg8f5gOerkvM
U32tDFyb4V/r8oJtEKnWt0XV1zDj1SqFwSl28uvypgbC/SIiJ7llB5M8ZIngLKlA
PAg/FdWU9KD5EWZfAQgxKfGcEj5wdRGBW5+2N5tue6qosxLTqPS9Q+COedZvWx9R
hAxoxDnB1W3eAxx2ttT19yNF+SMGJh0LQiQOgbeoEvvUTlQoOqwBlTjEa9tLilfs
EHrHwnX5/O1DYq+PyaHoOTD33JWA+KUUR2BlW5be23pEMeE+kBSfhMjQcom3miPV
hIWAPq4ADdOXOhuJkRSKzIdC8xtnjtNDgvgdUAzLjBPE7Bd0w2qB9amUM0zD3Uuq
NN+HNgZYnA1EdQK5yC0ZnsFrCBk26mqdREE/q9DCDV9QCRa16+7mP8mFPL5kwzW0
VWbKeYq9ePm1600TeOotlPhg18wl8xE23DQE/546CI+fUGyOIF7ALX0b+MD39598
FTmJiU53T9g02nZ+/Xnz4cWvaCCrZC/E9Jgx/f9T3wDJCfYVPjlJ3TZE8ziyrK+P
+YcXSKJb2MqhiZVJ77okl7MxkEiP6HPA7SitjdPPZ7B8KSdWcAbT57xSWwL87+mP
U1k8SnKuvaJsMWmN5+1W6sCbRjkzjkTE5vBxDEgPygqILvINTzQVDroaYz1XbOh1
3ihp4iRSpVVvRJ1JaHSN7arJQNkrZ8I2thebuPrzpFN3vZ9NYE0ZtPAj3/Ib6cAK
dpkLnCsMrgiZYFc9hKaqkflQAV3lV80zNQVMlDjWoKeTB2jDt++i9TmICnYi2lSg
r9x7dLhpxYAykSEET5WvRPzZTXAX5v7LaNC07qyJOF/QaimaYq1K5+kixXj8RvmS
TgNj0OfIGAYqs98JHHjpTTZCKvHJm+aO5weLUyeoul1+KFkRkT3AHlFo6tTI8dmy
Ky25nYSphl5j6R12UmqX53pW6bP+Ky1HziL2Hv1naqJU+1nVxF+z2iG45NBdXf5A
kqitFcgZWMIahiNChSREdVJsVhHdMEhT8P79nxdfXvaoO3CqVjOCB4/CPbn727eq
oYbKZTkix/7uBMGmQo/9/xXdN38KmV7l8AgfCXpSvVN2bTYVA40IPUb+Edx+aPKT
4SrHVptzSWk4txwEW2KbQ+WaLcXs0aC6TM8bnIgY+Ce4CmGdbpn8ilFiSJFv9GdL
6UcJolopYWy33mtBO43CoLiV6lhg8c7ntJ5XTeqLT935pPR183YAD5u8VFOgVFKY
lEVS7rwmiVUiD4RpxY6gH7k/sspNNcwqAJ1F2QiTe6EKr+ma4oFP4YmOytR+cFcA
uFOUlWzD4HSqnX4b0xvjm+mh/qlRMutKe0UQ8LxYzp1uYIOJalz4mGXKe8SvIkM1
Q3aFor+NWamm6mojBY6qrx6UBy0fgyCP5kccc3mSDaqmvxHRi61Qs0bZwbObjyuP
TyAMAVmJtXVwZAs/PJsRbWGrsollomhxPtPAfH6hjEwy+sLCZVmxl7dn9rMk5SY3
Y/Mpfaf74bj6VnutjXAHWUb8hOA2f1EajTYtA6wGEz34m0XHA0TkLz+L/9jg9CO+
i1XwoSuCWLBX8avPBL/SrkfVDlDz+QovrEgsDTW7Q4144gyNzPsdtTf+bYXvFlvv
NUidoqNLUx8w84hbN/KpGPpGull+QUPQ3UB43XY4l9Pae0OSYiPqOnwstGnVxU4K
E6K9ubRCMrVigcR2AhO75EiyL28WvmWnoMMsi1rliKOsj1Wf59EiFUVD4NI+p5Of
/BI7nILIX2g5b7MJ6Aq73hp+tFaahy8KqZCSj4SKuQgrntnQDwZB0i/WRzQ8DJnx
yzPAV8jS7sRJgmnsJErOfyonop201Xqt1opyLTz66m/AJZbUvMwG7I8CCiypwOL4
2zl7uyXg+Bl5kTupAHEUd5f5kY+8R475LoQGeDeuw9KLBknj+T5H19qWwzCspwYJ
0ypSCOsAk5ff0Cn/KsKc8qK57vhi7f7n7WcB2aC9nPHjqPxGmm4oozMiN2chDS3y
Z3J2uha0lXz9IZMYdy/XGtDzy5U6Db07azk/7QY24ZIgB0jsjLyHPemBvZfhSpD2
1xKfCOYzMOGG8bvKLIpaaZigWevGKEJQIqIGK+98pApz7UUY/mo93txJl4q3scV/
PQfQusGU6R6H2ZPo1YjYsWRDW97X/LBK8IkbI0d/wYtKKAhKsxD3yJtA2DhwNG15
gjdbvQXT18bajTmeZ+u3BsZoaN+BnP41abBOfUrhzLcZha9tHMJy61cogGnFDPop
OtUAf/nWlf/NO81os1hbAmHp+QgMMRuSeHUaH8g/Nt2rNfMuR5WNhp/2axOvqxcV
nqvQoeeM0tgrvCO4Szt1FCrO2/5OjCEGhtv+om9k3pOg9SgM0Fa1toaCaQyFT8Vo
XkiQLXYxkYzYAVyRlGWu63mZ3KuYzkoRnrY8fj1LBDy2M2Lg/QJ1tJvsqn8nxqc4
Wu6a2PAQg4ixo0Ql5Wvin2ta3wUdjH/hKf4RUZNnrX4f/EsID87kH+V7K/Kt95/P
zVrNbV6WMB/YpILLmVrENMCMpS318YEdGWS6U+IdGdRQ3SDKn9aQ/7YnfWae4dVG
AqTnCWRaF57Xm5I62OuVV1SNg8xMzwErAPsNzI3Q+5Cts+hO6htmVhw6uOx11Bkf
tuqxBJPNQaDTULyBgTcdUqGZ2t80HjBW9P1ZncAp9ReHoGDiwrl2lpB3CaYpCggW
nXNBcN9LMDDDqBI5uazHj/unCi3CKw5H/A1lj1DAbN4bM7m3/5s/kIoEx4S++AjQ
dAc3hGX1wWu7YZYem7lkWFRL2GwLYk6RGGVjSuxXqEamrspVYq03/fPG0BFNeaLC
b+mKPKGThAtVJCRSSRjOr8B4/fICA0HO0YAu49v9PxbCMwI2W5G+78ENb0nckrdZ
y/ch6M0ufj7IA6gFGtLUBRTgLHpTIK6o2S1XWHUDFfx6OXMfUIWmm5l3n9mLC8cv
RsZ0ILn3dQ4BwZvhoBtUla8HDpYhqF8nPhlQPcjJL89lM010Jfb9GM8TQNr+KgRQ
DgzP2bBCzA1gM61d33jrqWPzYqGe+ngdjYDAaRV7QYjW8Vao2FRFYxQBS1SCQXDG
pHXlF6w8IoyuAFj4YGn4caMs81Ht8M2UA42VHfV2dvh+jdkh7DDCMtfnB1QOx+tb
6L/8K36a02vgs+bIFH1j3/hEPa+eZM/e3cPlKBwMQMUDwfRdqftDzsXZ1xsHMz42
51ZJ1+D+TDaW3yagN3bg1NTFKyM4w+FGwsX7IyMp41tP8ESzQLlccqCUpjZLVvEQ
FJmlTozk+u2dLsg8TQaMM7t1MJlIkeOvOw9Db8bQ6plcoZ9OntLNCTv6vWn+87aY
n3NROEo7JZQ9MekqSYJo6bLRjAYGnmSg9UzdFHUnHc06E5E5G5pk8szajIlUM3gK
P7zGnGqYUnkHd0CFqotl2nBNdfmoQWMYTmkHjp4dz3jvl8AAQmbla5IltnnzCDke
7QoLMH8CxjGwVYDQxzJag4jGc0IczcrIUsmx71eY9yRv+hCot9J/dkYJTvs5yUPB
NYCyJ+Gx5NIMUhxqSQoUi4Nsv+y0Zj+4aRNJqLhweVP5wYb/ZqKnfL2Rk5SSMOXY
zWDcRsZ0N4VoCMe5cwql11rPuzWAhHSWqfTDlux8EBJEPWeOuXBvs3smV06Cg0zd
a8+Z5S++eaF2IUtCPWCT3H6eDm//LQrWxEjsBQIz0Iz7ptn2vFdRr/YsxB8D5srf
I9Cdaoo+Gip/TxB/cVK+Lwts8ENYJ2n5V5abSz2Pc2eeUbQPSlmFqEbaUDFxTdVK
GgER7++Q00lHS0CB+VxbnaK3EXD9z0cjJwGy5HaK8SE2dwQrpHTGHqrWAexFCXr4
MTWEVzgSTsLHOv+PdqSrMouvIYh28sUYmkh4ALlxQXmAoWnBWbouv3miz3KI5OIQ
Bh4ol1CyW6G/NiLWVmhOAKYfjMOqj4NajNBSS024UXsI13Im3tMzjSZtFdQPR72n
M+KxFVwiPNOLm847fnej36SVUsHkiaXftTZg4Zn1TJXlSptqBxFbDLamam31hcG/
H+2pKxFqMMbCzeOMpdyJPo6jVn9HFiXt/k7EuCmw5L2AVR5M5VuEo4tZT85pGVzW
iV8vqsAIEQaH0pRQP+4TMidoDPijC17+kh0aWNaYemFFfFlbbZif/9eiQCrXfnoM
cWpm4OTXsFYgTuGTkf+PVIQaQEI8Kz5cdn4qE4gWeG+oNJi+VRYQK3R/Qz3+WoMB
l3hvHqUbCBImOYWiYQt/pwj+HqSFStxa8ou5YssvAieLhHBxcqSY0XrKY+kWHrKH
rD0tepwp8yauHHoYZ+qixWQ/tDoTmTt3GBkEn/AOB+/bGaluZekiYapEKK12e45u
3kzIboEiNfFa7qNAtcMnr1zdsE6Ev61wJGvoUykSR6CqUUetwbfozLenLBJ6R74B
OXdS8+IgDSHQsWZaDYIm9rtI9Zvdqbl+/qYG19jn7HOzT8c54MBkv+UWzO9E+Jy5
luUCqYct7P6RcT0P/yI+BmVPE01l/Spbn1LhF+lzYJTLarrNDvEnTBzUPDIOBmS6
DmT7kn0tyDP1v6bqKppRru1ZduntBOSaLhAGY8gSthlHO3Xk27cmiVUYIchqg8Ao
+oufhZBV1VDZPZawOaKMsEoVs9Zws2eWJKPDT//Q9zgfQrLltpDIr1oXaZQkXTPw
FTmlE87JOn2OMXOX2nP2jkzGt0wV88GKyuuMUw2Hl0deSSG1LMZKKJNtlu3LSISz
1nehAlr0pJSdgsJVIuQa3aY6cbX2aNjjLeWJH3dJ4elEM7OOZEYwUZk6+smhJQIJ
Q7EO1X4ovEXL98a8FA3q11XPya0THDjo1TJHCTQjZcvZ3EUo8BFYmpkRHqp7DPYO
4ol3ApQYjSTNaeymBsqER8c0xulaNlmfIQMd9VOFfpjnY4c9UUDIscjCXwAvo6Cv
vIF0BfSKkqRVlkbsBq6USBuK2TYQ8muj+Yy+75zb2nvmYwoht8tUT92ATa3UCUFi
9kVmU75qTFEz8PpBXYNqjOlND/FPFDZB8PTMmZmBqPiifjxoBhvseXcx8TuF+X7Z
QaIvkxmavty5+xpnJSyLXCjt8yYiqVnlAYqZaR0PzQloZQRtQOjW0q2UBmIXnkZY
CNoeBJV3QI1bTNKrZt2HK9uQHFo30bES7NPOMZFeicCY5IEGQ1SvWd08BIj6qpjQ
idsmwF5RBfGjIdOkh4AuAIcEYEA23Uk9gSM0olwMOno/2dSpPQzVprWAPVCnzoWF
VZ3YHYy5hhkkvrvOUUBF85OneG5XQjcYtVAC0uyxB2JDqQ3PbliFec2ajp7kOspS
R8FPau5bvmRBZxBRx7ewJx331d4P5XCwdRoT8NRQx+CqrW3uodeodTU/BmpjVQU9
pn5IBgHB7WMTi1r3XNSHiZiSlW0G3z8IB9Fbtx7vsWtarUaaeCG1caDSDVujRE70
SV9FRHVMn3XGoLcIWwkHQrnhGQMrJ3MRi3rDOuwlrg/Zs6H61SwNzfOEVQCFWJd2
Z42PvwJsxniskfk5XDHAhq/BUY9tSxBD1bnwYOfRIWxy2XeECUuqSuaMrM6BFvdN
kPYWsUTrZ0iEzCEApBcu/6hyk4OgrPQaqdjCVjUcIBIP68M/GFrC+GY10/PxJOiV
hPBat+eqMkxuhc0YTTJDEyXgdGA2kgtk3pNQm8lYi6v4xjwZKXy+hv9kYEJwcDob
Aon+4zm6wKmbgkcNlUUXx7Gnfqod1DVcg2Zh7X05AX9mlmaXaYTqg/wGSZqMKFQv
DRNENvpbA9nL0KizUzxqhKiU8ZAyrjMkvtAeqJnu/wV/wSZPuFsrSGv1nyIDV9WT
Co8yTtb32wg/VzCTIEIqmSZG+sCLIycF/vBbT7yY/3dFxvuC0ufuVwCCPO1Bi6Pu
+QESvxwK/ZdIrkWFnjua8FRrmm2863Cvnsj4ajIcXf30Wi8yvpgkRxE1KAW15brO
ovn9zLY4cJ8lPGdnY1C18mXZkGBcrFy5VwSpF+aNZfJpT8WZZ8muHlLA0Ri4s5+q
WiC6976o/9W2jb5c227UaFdDFwlZ3ejXxQNR4/0XYnjzkiGU5PQRRdWQaxR9VbG4
9fqteOKhbNrY5T9OB+RrxPxmpy8e+SiiW3gYMfR9+HUXLuKvYmsKre/UvoQNFM66
ZZVfX00NNDk9jBrfcOCAoBJz5wfgh+8UA/nzxP0pvcOOM/MGdKu/idWCAHBaQPDh
rrm/hn3D9ZJINDynj+uzh7FKR7d76rw3W3cx/61Qj95XBCt+rYcHCu3kR6bKP/Hf
8s+FbEk0O4kufv//dyNVvnpYPCBuqI5+iN7iu9fHCJJTMKmxKu2GnoxwL0prMS1G
eWbVzO2cippsEKqdfVa6Br8kKP1M5zfDy2snGXCQVpnl2FnyDQdBVskecIJAsZpz
oyuFC/xFQ/+IGaT4TmU4Igrobi87ljUWd8bLgoS2IGzS9HOtgIrX255z4Ebc5qtI
/HOCZYJaM+YpZtaAiYMWB/tIbBYlzwukfFjBNPc3yGIRRY09HjJHablrl8IPI9fq
igwnpryvlp3d2EstU9Azq3PmZgHlqzV4Up9lVH76/ohBp3X52k11aWV8O2aS0q7K
LsGMLFID+vQ3M5xrMfko5TZfW2FU8DVaM2lgyj3/VPqFwJ26eJJKQn1/i0fvWtwb
SoCphxZAh5KGnS1Rp+TQCEATGUnARBQQXlai/woiUlW78rKOsjlddflV2iMlf+dm
jEtY2Js24N5ROG2zcPo7v3/StxzXFFy1C+tHwOuzxaagBZeoamWS/Wnw3ejSEqc3
vN5yRw4oPimEEVC/QHYWVDfGRiGVzK684W10cHW4PpHrDisBIest5vuk0ptUhQ6Z
enoGCZE6bKNm04FTcb7p4Ht/9RgIsDuaeSlJy/lJVn8DAG5yQGcB8HjRCUWctaXB
v5NauC1emD+aIJ1gGFU9uMdyPIQoedKxWI0jBs1fijp+d/G6xvY8wEMMmIDzTzoY
ILUi4a6+nqS7SM7I1Ot3kmTsiM9XgoeZHddHCyJAc6DO+ui5OGm+GNeQy3TIn/ZY
VShdHFjnNg1bbNsDOUk4kQFPOISech+OmIkGcgNsTo/xDUYBlYs31FsymyOvJ+aI
0QQfDkzsdqZXTak+45JatADrdrus1vml7fKdpBqudhgWaXyVBAtwkdXGTTz/atqk
ht8Fkt0yreyB8NPYEi9WyolFlBggOxx2QFJ8riz7QoMK8QgLTite8y6xZDHEQUxG
NLEPvNu/u/WRi9yPv4l4O1LYl+jPa9RkgxzPToGm0JW4bDmcMogpyGGt5kQBjZzE
WOUNdAdwAvmh/h6zMdMfs9CtQCE5SUz90lN1E5HpCi6kxSCHLenZszwlDYP4/X8o
LwWU5gyffaiwbU1ds4qfG7gt/snqv64aIRQ2zFArnIHvATPPdbL3pOAAtGrFRLV8
mbamlzOR5KJN3gLQFSV6L4+RegzZxiG6QdFUv+YGKh49TPa9oeup2GwRqTzgj6RC
ffzvOgQxhQF6PNIlDWCTWQLaiXX5LE/myczQfWuVlbAqANT4kcq9aUuxF6Qb7aqm
ssoAFLmRl6tIIsOoPXSS9BLnEAV3uqVGFzPtW7QOWWfF1fhiTB9XLECGASAIuZ8v
FyaN/3NFCMxVIimlK9KcpEeSk/QDYOee1+fG0/18KV5kAOuh/AhP9HIa06kl4xA4
O9ZnwHwHKCnopWeNSckbIj+qrgHg2HikrLpXeodqm+/qDfRVoUv9xIeVYu2gu8Gm
yJpneZSMWFGff5kyD8Cqup/MYo2RwoULYgIRG4z3qIFS7tUigtHBh0RH13GdPkAL
DlMTYnTJby0/PrdeDEeD6q9C5y2m+atJurJ/6xAIcz5M2KvlmOfvjKFPbnnRVgRU
forewRbkkuYU53Io7Q/N15yZcBPA4eXASpCilPlK4ioGZW+3F110iaGzlgMahTkw
65KbwZdGrIOynJchqlSQS+0mDr7FQ/4K4HTKJkDDyyNlMto7Gxz7oI5OCjO2rxcg
MDFMvP0mUg2CsSOc5jFubIbpstJrCjt9JPDiQ2af2JUjC6aNnhIAVBqtmg4nthcR
KnjyNR294dFmSK329Ub8oYGpuVAfOEuYT+57VisVco/DrXX6O8f5mu8Hhz2dj+Ld
ivP2X6HbYX/h46r5b8isSryGfiQRTsMH8SnpU92BdQWN+uWlHiP3u5kBEoBqG1YA
P4y2cm0GR6PblQf05Vb4sLfF/grSZSf3RXgu+Z895zlyM9SD4YPIGe2Z/o3E0DFp
M12C/99cKZeQQjtZ/ECpjjMK1cudtxoxph+wKI6qCdupm4Cs34rTOF0xQliumi9J
xY8vaQRk2KprnJ4TiD0ZKJRoKxLYypB28VPxw3qrEMNE2nj7Zftn8uDxsb03oM7k
CSjyfInTvdJ972KNcO7zW3GK8l9URFXNah15CSsA6zipBEHG9YOEpulbAVnvIgAe
uifHBdBZDstCKTaSxks7dRNV/GF13AaaeCF/F5C2hiMlANM13mr1urdxB86zvLx6
ej85CzUCYXOfgYzVxWQlre5gRno46CtGnNe7maL9OzumIxriKp3Dvm9znso7qdBU
5d0DpF08QHOeprG0K6iMzw6BfwbQ3H5ncs30s/xVoWzVs/CyNESE0h+HbTVQwwTn
iDttn7lVeN0fmuLs/x5oYnMii40FFlFFcyINKZwmf3v6vJqxKmcvw5LaxYy0s/lV
DhewgKDzEn1Rmtvu5WW85yakZ4i8E6qRAxTHnF2udExOVPVkJqQYXb81aCEcwGFp
diMvYGN6vR2kRJzmLr3DYIC4y4tMQLjN1h+A/yd99TVixHYvOhOXEaWCJZKowFYJ
jCUO59XttEE+eebgVGalYsKXrZe8esjFlSH+jc1Ofg+wPy9gLe6PrnyUGiBLozRY
sOpzqtEDa1TKCRmp3Byw1K/fsuj9Ua/TmHsHTpT84qGJgLr7H+7Zqq50edskgzmj
Ajx3JHI5jv1w/dlAbfgqtNeHAyS50ENLTziF5XItySNp5BP7GUYb+lRJje+A7kip
IsF8i4mwzx0f68lofsTBcB/GQIX1jVMlOYjHKonrt2Nng/J4aw+JOGopBVZvoX/r
Le1zuKeUxfl2pDEc4gDAPh/VKTgTFEFwDh75PLFx9XOeYupn8did1g2OUBpBSFlw
upkg2TYa/ot7ShBb4Ir9LAu6f+AFa3O9YpYDWxuciUT6+id3acjMCDRcLPOsGuN4
XMTP7hkHHtTVgV9E/wRSSrPx7BlV8XrbclDifCM/cU/Kgm0R8YcYoIjEE5nRCtEG
dna0TxSCOA2wE//mx8mxn297cD9zRzaJKF+0ks5TL0bQw0XCYRIMXrtBadTRoOOk
Pl2SNFfF96mqDDUKJCm7L/YVGqvdmNO6bH9fdmnpwym4uWXHRDzk0SQByf9o+Oio
LM8cAB8I2w8a+FK806FYTShg9htSwtAWIfTftlDsjLoBM1TM/gC9x1n0rSFbNFpD
jawvPwzVDiiYSHncIF+/QqwsH4CDbgOPFyEQk0Ax8SiDttG28xUtq8Jqubzp1Wgx
0hIKj+XI6VkEdcWsmP/bVHoOWgt93oVUwa5AN9VfXCcrhdcI8JdVLmOZVcSuRsG1
ZJUVDeMd0ift+LRAKAhjFOeGYJe7G32GFVyIMKvxg5+SD/SVtcGqkyLcFbboHann
qJ/e1JXfCpZNoMKzbtYJ650irgoXfhQQkF4Mc87fsdxevu1cYJmZoZg1vDos0jfl
G/KiFyU0fHSj8g4sV070EP08TK+h2JtenfBDAX/A1ik4JEzxUO8hmfNJzeXv6K/v
Cf55u0SI3ArzotoSoxQydOQQjrs5EiKVG3iImjXpXtHKMFqwW5bxPri89I23i4WY
PrtE5G6lna58Lbi4oJCkNVUrnM5Gh61KrxkuCaTz8nFZmILvu7yTne5hgkJfTJGE
55+b+zSqI9/f0LOK1rOXUjgX6MYaoNIeO8vzzCh4C9OQZm2ZHAa+qaqzyf+LD35T
N4k/StcYGn27hKaiETnvGUjIdQd4DrAD9oiCXQFn0pwTmt6LbEWgPB/ZU913puxn
LS1rQtXog3qP7uecVuyoa9HSATESwUlvwt7jW0rfkCRH5cru12mDf/z55nzBO4xs
R09PT/mCOsUmeSOXMnDzk8FiWDBRXZUg7Fr2Ammss2jsZbl3Iifr/yxiROKtQnVM
6UtnbrY4gUl69mBTsVg/SphW40nHQldWaztmh5nNfebpQUCsBn7mucUN0uNs/fk+
kNAqaz0XruuDV2MiXvaBnr8eSye2WENIp8TbU6XKAu/o4BrmKD4+HiNlzwS9xir0
OhuQHVqb4aYWdOqSFPkOtzYPv/0+W4tOR4eGKxSfImaTzC9Ot0g8R4UqPbi7xGs4
mBdmQv2JbIu44L3IOs3XnTTApNswW0iD4lI63hQ6RryWvkJQTokpfJtU4NsUWhcb
6Awoc+eIOS40w/zrdl9eL8ucCv3tz6Jfc+5NSdgA4jd14Fkl4Ebn9hM2tb2ob2oO
k3NjEwrpick6ZsqgEQ631PcBYL0eu8ylBVX86YOBTxr22BCCit9Vfiro4tQwTSNn
puvf338++ejFUWPRLwuFFhdvSGgRQd+eLEXlWMJEf4CDofyaBBojt1AqK1W5tJd2
LO36oE+FyugxnFSUG6Vhw3+Z87fVVXwubPuf/ye9nuJSGlmcKMfD9g4T2xQU3d8h
GM5qC4QiMWpL7J0hiRs2rNEZi+rjaztKjnfM6ex0YiPWw4Hw1w6oaEPZS79x01qt
abRuuZ+zZIFb9aeAmeruwBBevQoBbr3BHWpAbM5YgZ4edGp12FXxa0Qh6kCYG1jb
Y0LVQvkvn3Incwq7eIgbdL7b29a1KAXjq02Rq3CM2fyKv7MGIroLTHSY5nHR+Vvn
ZLRU9Nuj94lAFZaFeKYahJlnmqDh2XXWnvENxlSZsKUP9T137XNDDBJrSrsNp6LZ
mx2vKrWZBJn6xqzILZ1eu5SMSftcKaH0yfEjmWjOJ8jzlpMqYN1Q+KqmKSIWkyPL
9b4JTQGTtIQ2P0w7xLFPnvKZn+t3/rlDjaGtbXhzGQnRSIpNYijKP3liXdng7GVh
NqPB8b0lYyyPVRZ0U4flSYd8nqZGuTM1OXgaw9P3HhSxBPf6yrlX9V7SiuZUGkgn
jUsjYZ7ISD0bYr8vWWa0PTuNaDnU2DnONrcbXqJRme24WUQeRcDrtkXYUmfMsNUq
4RimKm+bSsYV0nptWkPhhV4QUAVxwDuTdWsz5e2+Hs203FJ0PZuCSJGnUDD/ClGM
LhRRCO10QVrVXqMV0ORR39VOt1+q4pyxsj9AEcV3FK7iM46Num5FFOIyHyl4RjXS
XWuj9ZF7ny4P79vfnuHuzwghsbKL3H8nlapLSURj6mmzXlitkW8APyyZtz839pFS
/s4fnVM5r0GKaOY5BBahbyZdYEudvhQi+OZEoVvRsiOLvFciNQKO9J2DnLvbt+Xw
7YHgwS2/t+TGBs3fWwVMi4oekYAIflF/jM9SQHyqNcDYcIMAG99i2sH/l527Qniz
yal9Hh+lRCcj/lpjhdLKlE3Rl5XQjlzar1gvU1vlyE89FZUQRgjEAUe1qIVT5FS+
1b1t/roEKI6aKBKaAqcBrg3LyEtsgyYAkgmRl0j7ySXsKuuqJlk81TqPRKGfybB2
F932pfsj5cdsUusWjwFO5B1OGI6k8fTFDK8gSBKX+hze6yUZU9YwPqVLSGLAuykW
W+LWkg7SZ2WHQoiiHMyfxvdWLvSOHC48fsc+jjmgrpdRJEOdjZiqc2hTM9c+38aT
dgNuEmtaTkJScTPbfjpqToEaaRenXQutItAKyj901D6l60hHCGrRtU77nDa6HaFJ
FLSBnkZdUlMdKIoh/zemCD+6HimLEzOs+R3I0Fg7/nr5rXwhrVIpZVSd69NJBr5G
Qi1PNt6uXfxD8td+drOObv0RNIdxcCxGdMLKX6RAu9jUWtKYWoxqphd+aYTH31i/
HARDaabJq/aczylF0rbD8AQvGu4aEK/VoK5Xqj1aWZsQAwMI3tYEKMynkP2PJFz0
bv+QBGksqTNUAf4WUVKKEgIWyXVEB+7YD6FYiiNB7Ipr9vn8lBr1561hz3zJtNok
6FXEEP/w8WYdw7KBQZPjmpY+NSCQQ0gJ04lH5LCgK6yR+mE6jvlPF/PEElJ+wvqY
FkRKCkc+eOLy7EAFc0sFdznoIHyEVMzu5F59M140zhlGmVJqoKfdnucOK2fEkx7d
bLFofvSy5PjXLGQvF6uISyYyL6UR3EBKDboAHsu2Djjd8OenzBKFuOIKArQDItt2
9dDw2W25RnLLPVTPSb+iZyriL9+4nsrGluLFKmGf47Q2x0CW4PHgoOdX7q+c8t+4
bvTSYMFiQmVJvkYF4+3p59pfMA/bsOuDhg1xX0uJugMvh4Q7OsMl4U/9fcj+O0DR
bxD1g4Qhrjt5032LnyU4C7cz7VNiI7vOHZqFOpadzGIYZmCFJU2KxJFQ6AMwbUxp
2LpaH55UNn9HTg2hW/55Pluaa/5mgV4LpfMbuVN6oqL8eb4Awcsv+YvXgYjIUHXl
1Ua+/q/XOKD3YoVAq4HacS1UpbD+VaS79J+8S5tZ5tbO63Kza2YlkvKi3u/10VOD
pRl//hqsqCwzjezx3aHzGvIsZ7c1PMUYIKNbxIE8LepW6i20rFZXAY0FLx5PWjaK
v2lOwO+4LDrT2faa4hKUktLzLf0cAA75AQuRrSZ5N+vqMGC9lkUnt5Q+0tnR+0fK
iydk6USk8r16MU/KPJUduktvGr1yYa+h9+0yekPKi2YsSnQoYcAnHvJJd9nU8Hg8
dQ7kQXAz6q2xxYw9h4e8p7A02YjxOzfluW9YtT+RJM4YkVUj5Pf3dY1u+DoOHL/n
yZs6Px4TYmTC2lbjA1IdYfdeK/F0SKwRgsbmr0EySUFj5EV96V4Y4qckAqD33n7Z
Pz+Lya0krhsTWl/GLWvtM2x1BzGg7rA0LB8sVFTD5aEg0tzNW2wlHnNl6zIUG/nB
fNHNWD4GE+30TfncMEVB+pnjuf8liEscZsXFxtl+0gJ1uEqvXGYom+WF3Vm6Ge6w
vtapEbYoP1pMKPG8K8PJp1aijrkN9NCG52ltnmqVD9ToLzz/uAywHaOKO/zIyPC1
um9IdqClUIEl0vyLcFJgZs74rBHQNpbUGu8Ymu/2xCCwzCd3bCUr+09wPmu16993
2Hk0/4oQV5bH9eu1ERSGzfxB7fB9oNvnblYx1f1NGkbaVN4eo3kU2SdgctJsLuAl
w2SwkWFRa6tGzlt0+bDwSyTuO4y/H4rlJ5foeWMUylpCbLq4caqJIEVLQl4H9xZN
ZZdA6xyFfQcVrtUyMyEcCkQIsu8zCdn64oZCA2+/BuxFvdeqEsc5Sv4+Mn6MbBXd
kkW7W2gWkNMXRPBgbfBhcfL3YlXJ0aHqLrKa0zrJa6Y8cacte7qia7LOtOguNLHR
XHDe/8YHH4EWJsZ5s7vPkD1rDA8hflPi1HMJnrrEByD0rRXCf1rESxA52TkQ6O5R
n5na8STABNwAkJgs1W0d9e1YohquPadmN/h1ygZHvLHbECIWywZEVXo5/cjl5rUR
n9ALmQ+YGEN/VeQ+Jhpwj6+XBl2eOOy7hkDhfLZz+atlwrOMNIVvVkWxfqSXGqcl
zuVpB3DMVaeEhcVrVYREruwuzFu4+i8AKa+3fDarUCuxrGRqzSG/VpCt5CK22QvM
pkILVySUxQQBicfe/iO3c1a/BkmsdWrBz+ScqZxD4x6wa+HJ3hiZiWXXTofEr8v2
H109YkJMlOMMHowhWEZJjhuOAp5Od8Ff7jwzrw5bM5fvt7fpG8T4MxWdMI1Q9GAJ
cA4yq4jKx/ZUyEEG1v8UZKVPt5CsCz0AfoSV3lkgraglqTe8K+pTYX+aM/IrJ81P
9VEPrqTtrbAyZNuesrlu62o6L2QBxyrM1MOoQFzVbZ95oWH6/nLDKsFIn5SDp7EK
bwGirCuAmcaEryjsBNNoSdr/7RaM0OURV/Git3cT90LXDBK59wWaJ5L4ZhJ3J6FK
OvVljfIjSkKT/wT4+4Qju/DZY7oRlj0gYqTzNcrrTu1u6JNbHaR3o/6Bfqx6alHS
RM6qg2axBz4iP6I9xXXpvqb9lQesfUJ2aAtdCWAwaDx0abUODJAYAEaRmBdvu4w9
mCwTWW88cDnEK60z2is7v53lBIHq0OJc7Owhi2vXnQAcEYocgkHaUTiWIoZFp67c
D35CDWjFTXRSrsPNt8s7Wu9U24Dir5pNtp2Ld2VSGFoGh63BAyw6OQvhFz4QzCQS
hmp9h7YVB6gln3J5WkeVi1Y4a5hpOcHJ/7krp3XJ+VHcsM8h6pgZF6RGN/XZlSe+
6QbdzjfDBuJGhg5WbX5iAv7Q5qjRrPZFyhKG+pEzLMpW7+vvYog9DbfJshyqAETF
NWJ2AMU+TVWIwsCU47LjcWJBsQLwjviiXohnMu3ssGm+dS1Kk7tUGMjsBm/qrY2j
nj7BiaX1zcZMeGQIDvwjJPwhgFO5OV0SuqDTcC2erSKzYFiAW7m7lFp0XfQQ7r+X
XbNXO0Ld+pW4SPaw3HGehLYwB+v22o4HE0GuIZLfUxCU24rSy+tOPDMI8MpeV+PI
clvaWwrnFFgdA5x5x/iQ/mpbZ4N12rKWjKKtjiJZiKra4kPrBF69+I/CD8jqnfuY
J9i5rZ1rPVg0lpN+5OEhBlY4vq+htGxkgtN2q0NM73dWPFzC72K5MCySxnEkJH1S
aWp+mFhi6jRTK3kECtEetrRB4aRcNyfDHEtLsnMMU9hy89NH/lBz+6A6SURtNLMY
CuumKDSLuqug8SzA6GnuQlA2RwxpZuBZR2fpBtEjU5JHhzC1U/Mo/x0Bv3NBSAIO
slzg23jXipp+wec9egdWk385xj5GO634EXdBYHCeVj/o9NrBbG3aTS+3qZZKK2W/
K+210mTGvPCVGeEFtvTK8yGdy9GESAcnE/HFACQQkdA8MTOrH+l58A2Gybufm9bv
kohwHYLnzBA3iJ7pVT3PR4JRvIN1t0lzC/GYCZl9v2aF2oqY80dctXL/jnOBV18G
qFRQfNaxO+1+V69LI31kVhBdilLjuzIZJZS3Mdj6j8+9cGwXn1mlJuUDnRXCpolM
pp/b9cH/ca3EpEkK6u8IL57zdlPMqyDj2KA80/+mrR3K0jL1/ERUiTjXV9Rw7lOA
DzHWiie7lE6+48hecLiLTiNyljyaHGQkc+ZUpYpUjNFEaDvtCrniV8ieFSR5cvKL
KC5ISH3T/8qgkuUTZfjQYGRHiizmUWy7/2ttvF/7e6WE/VY/GzMmlwmnb+u40hT/
gEh0MR0ZAB3hroQ3/RosGP80XyQAF05EELA4P99jq3cBRlHE5Vcp/xWDYXE7bJCD
uvqxDWX4GEKuTZVyDAiRuKzWLHGOlDY47lcQ+gq3Km9qi/RfyrgAjA31hAMqCOqr
tDxxfqzRJwAXHTxQRqPhEEZGL8eKvgKPrL+g4w0l5gLrct/I/d2jx8QeU4O4vWbs
T6j2mTj1s5ixN3wVKwzRN3yj5Ti2XG2Aw9TqwSws/gPF4rDth9ngGaw8lVRg28jd
ckApG+KzEL1sTcZzy5EfUzBovbBqFhMymQy/mNKNsZeN6gl+iyBKJ0EfdnWiIwNB
2njBfA9zfLg6APl5rIguOFwnCbUb9WWTNgIAtGHqsHLQSoATpIwCD5INxia6piUw
iFTf1h2ecxGnsSFXVEnOTZayC38QC6dhfSHAvCHGgzWapUsRqzkEHjw87T6iMOBW
zZp3Yq9zHZWMxULU4yPxtE+yo0dw4mKfB+PTUy8kbCjVhaak77FdlKEeLDx1jsje
c4OO37xWXctPx52szgkEjUNUS6og2WNfszjPehMgwDyHQTawZs57zuSyp7OXYS3N
w/V3OME93kdE12PAiQ2kPf+yogAqqqtM+rQmSzc4N/1U3EKRnNtX2aA6Vib64gdj
QMsrAxyOMM/+Hcwfd9kKepOrV7SvebbU4/AvoMnoiyJB6BeEtk2i7mRAkzgd4NOO
rnB/uVcmaydQmmj39bALTrk2xozgAmE37cwdbaeNZoZLOt7pxulPjytdv2Mdgavi
a+ltOyVK8VMXHhERHyAV5nHGnvSU7cVAx3xXHLi5FIOpq0WjERyXnweqXblCvlHi
s5CksCM/52az33ERZoH+rUQrQt6wwJUBwzqaMpHFcu+ekWbXU1QZbD7g6UMjyb81
dBjuRX8ZM+3hVJjVfvlqYDb0eNZdxBa61Ho/L+qwVNellm+388rOrY3FRCP7kPFQ
yzRsmX8yomSzwM8ZSMdqqh6Nd6NqbQhDYhgRKGdA/CbRt7Rlfwu63mO4d+RKu4uF
Ie/Fro1uys2eveaK9JObcP5F3CkOOiiObZh0++6aQ9HqkgNYRZP3tX5RjIRPJWLh
hxe7ajj8cJsWEFx16ucPBvPs9Mz8UepHrt0FytrZYmPCDeHTnMwg80/tl8tJnKUy
VqZtaNVRamjVjI2QgpAfzmJUAH/fF7AQGOxd0T0MO/te5tu69S6FH1dusswUpeUN
LYLy6B7vgHDC0SIMyNNiysWQP4pbDyBTu71XTC4hTlUWBRIR7NoUbKEdlIK6vv2I
YnGd7LgfVasVDHo9n3g8gbR7B2/A6iuiwBZTX3i/RcX1CprPiSCAHyTQFm1rXEKq
WgWG8zw9Y1m4KrMaV5aYPQ+SClIXzh66wsCqMOuTS0TqzUSCqHLRm3hmPhfK72mM
Mb1MD39ak6oUQPhqAmCuyp7Emsv0Gn5LPnQ24UHBU86Ljc0k3ph86drx708KxQU6
3ZTJ8L8E58fQDVti1E+Nj0DiV+kwtYbpGoJxpXPX22ELGdNHvnRqzR/DkbBWIlKB
AMIpp5AC49oxjp/xsJ9D9OY1TNy9AZoIn/cjYccKeJM5dUxZJZnL7efzG3jXlLLB
idaUUoaHGuqm6t+lt7GoSzSOIzCAz8rD+M/1r8x1bj+FSynfwhXdKDX/20HOAolC
sICmKlLWAEHZcDAcZWLmqqyAJ2yyrDs5bfi/gSxK2NWmQi1vXQINgsJ1t0TTd7YF
XXBw0WGMeHxifsV82Egaf9vOuV4z5PMHrUM37uW2xvFRbj9shtV3miFtfzAKnRmC
eC70ziLYY/9zj1dFmLxuHvG3I3jV5NHf7bkMfVUSblnZ8+RABmp8gb0E/bkumrnG
SM6Xnwo60PAPzLtySxFJvRDF4897M5IJmlCG3EHrDpiGPi1+Z1jpzCI66OTE7P1l
MFvazkpFHl8X2lglK3UZUrAIYk3AwAVq5a41fc4vxg3t5njApGCHUxZ4oopILtRy
nvv5I7NN8P9GzCObG3nVyrNdQUbDuKoMoZQ/6vfPswVMB/lXj2M6P+8k9Hgea3uc
p/4wY2q31Os/H93r5LVVtUoYP7FrR9BuGFyiZr4f+2rCt1EadfwWpmiwiiFAOuj3
ShsOg0jOdjd31KjWhpCHXsn+IBetDDRltmpURqaPMDbEhkjjYc40m50N0OfpI3Gg
XKcMrgWIppOHSd3jwqq/TC2mbXRFunCvvfAWZ4yoaMbcjjn/YMq2cPDCoGfXLKar
VZVJTKuy7VKySUn1nQD+tTXgSUSGDziZm1+DaW+0NvahR4M9fnqi1K2ZgxILA5sX
R/5xbxydTFoHsDf2elPJNsRFyVLmCipfJxmxXcx2VWJTwVg3diWWB1aFh5LspRj7
71FaeEt5YJoqbQRQaLkJzXlnxmw21Ybfxj7rvKPdgrCVH141CKWPW3EKDVpm07+4
EbWJCcZUltMYTJohHmcSiX1Tf7m/ceFWTUbwe0Vj11p/0JE5TODqUuAJSH6G1HXG
ZRqTq6ySLbsYjBPy0HEzV0uJ/i0G/W8KV9LOrLWlrTzGDVYL7gPvOgaj6AxtYaoU
7k2PQmcRwnoim4MyigMCSVQiunoDAdwj5oP/snQcmPdVPxNHtFC/DJGyt/OJ/e+S
iC1u2qH3PmMM1QYrxsXfMjjx+QPWVB17iF+uuQIOXWsI0rBl59N/XFhIQFgFhdzZ
DmZmlym1XyjXVHKtdXP5+rxcZPnSiAPRkStM9+ZKTusPEVTYoBAe1EBt0WZc5e1E
he5F7oLOqPB000BIDFzHpdMTxkE6+jESXP0YY4OBIm6eo8mkz37FdWUcAwR6lASF
jeWBgWknOrFjCwtnjOm918GrOhgPHHzHUabKO8uvnT4Jz7pB0vtIZo+Kxo7demAd
ReCdk2YBoN2RIg1Te2X6dX7eu01wSVN3xA6AYp+6imX7ERsT5+6R5hphE2lnnhyi
NGk2t2p9XbYmOtjwUwNCU46DbF973jUlwcOaB4cUW2CW2U28VUqTC9cPpyI9qz/3
4vJ7H7x6/vLlXB8rO5fHRdECIF1Dj9wR/ZtSKhERCFGKPduGgie+6LiveoBPDFWx
lM3aSIw1L4xgaQIRWfdDfDLLuBnvEHNtAt1/uvD44S5ibqAlPZGccOHQGO8nRHY3
WcZtFfpLhXrZFI3BV3PsshjB1ztTUpBNhvyqfTJFuNU4HoJl89nRMDMDeUjRVfu2
8QS03LHIg9aATAYMqSbVy+H7/HW4qZI0RzKfTFkBJBTamTcpWx6EXFdNpQ3qyTp3
TtnphS8ZU3BizN4RcQ54PCPbSo/e4R2LpZTofdu9/9epU0SJKGbTkgrP3cxi9AeY
qPfch/kngcwDrn3mPh7We/nITsKsVROJ9KDhCAHSJ8jPPCif9TCXK8ByOd9zGrnm
i8rzlN47KUea+XlIkscq0K22bu5bp+uFNeX53jtl3YHO4RKfjZPZzgpU6g9oubdB
fdVafqbJxO6g5n07JhxwDuFWEM1XaajmalORbDIplWsTHLnG7yY5lzrYbrIQaarD
jpsT7Fsf+D1tj2QOupD4IwMc1ke7R1WxbxD++4Re+bzWsoxKnyGsUdmVyqLbNJJq
vyHKUswiV4DVci1TZOdgblUvbnlJm3GqhAyVh7FnY7Pw9nVnibugg0d9OZ702XK+
k4FyOk/pD3Qe4Eas+NAtuugIq9rPvMKXjARjLORkfP1z39QqyU2DdzM5ciPwkkrR
Xo6xAey8ZiFO7CWszFweiccX9ARDsR/evdhkyZhdheoVPCMtfdCp6pg+V3+cIpLL
3YaWkAJl3JXri2IREH8P+dne4OcRTN2mX89+9SGqjrOpZEL101IdDXWHT0u2Y42T
gZH+mpbKM+Sm9aWPfBSgqR9yy213mU4SERWf2J9/qftoG5ImPskm6b9LROuw99WB
1jWsSwPx85raukfISEmCImfF4l2Sb2yL24tQCuL4o0oXYmj47veeZQIFf3QznKux
ATkWjjAjjPDgSuhIH9eC0ETCpOF/ju90QnO3Kx2igmSiFzcCRWh3cO0ylA4i8+6g
GAIn5ABfY1+Emvp3P7F0ggrdTz/khnhtsrsRWbV1SDGyEL0SZqDD6P/KQx9lHIG1
cYORSnu1qYKp36hn08xk9tmDetrUA7xiQRrn0j8QzH3Rwy+J/QNELdGbvtu8YlMR
d/MyvT1eShiiZDlJxZbTQebiioJEmDAVrj5IjN6wcdsgWXds4L1xfg2/CkH4Figy
T0o8p+s0Pr9H0hF9o/Oz0e1sC+dBH9z61VepqGo0PusibA7+szh2wOhkEeFJolg2
aEC4z/q0b/46L02TlGy5XwVElxnlWCxuw6wT3e4ce6VTD846cqKqDqdNDBmidsUe
kWevYjzXmLxxz9I1sWzD6MjWhr29A9GITDlZZsPFMZDG8v8tQkl+drmxzt/0HJQ7
5n3XO0g63pqTbNQqyUPuhOsyjMet9xeRDPNVusKkKNkQEzHCmQ5pEmpNG/rEc1Bh
3vfKL8avmY87z6wj60gKWnRr6gGJBOizrddxL3raYtrtA7lb5c11KpfVgUUAzGfS
tnNVzf6dU20Shplythn45P+oL37mhLiz2KRgJ8sU2SddYq6KznOZ18BNJfddmGhu
EZrFjY5hDoU0h/WboIcHH1uxl2grl0AwCDeCUhJtLfc6fJ2hWV2Z4pQCzIMNvtMV
QcAMsEGbdH+Hw96Ud4hpQUQ9EIm5yRDmm1/um8hJH7rkFuz8cM3ujDWbKk04666O
5EehS9zM1nqMkkEoGX9twtpgcxcpG8jMmWf8F2Ith448bMKPpzxIYpLvXw8i0J7o
mvAjquXfhlilqf5+KAESUzkucM6L6M+l0qXItS1ncd1B6mM+m0SKoDEukCsd+/1n
N2vyP1Jx0AZK2qSeZlTdsVD8+Iq98FMIb2EQlDEc6ciN0m1DjuaI8/pSLS00IDgG
H+sRT+FHlLLwpbeN3dxN9u+LdXji8xwaSsgQ3znbYiH4kEXAUNXwLsOvqPU0/WDL
NfMR3zLlwsW2Jm9ZEDRZIWIAPuiKkeSwz7E+4yh9exvGqcZQs7GcKrvwebqn9QYL
Rp7cYPYA4KasH7D+ca1I3+keg/BRiEUb5WhIZa92UuR+Vy0nMYQ+BMDV+r3mW509
ihnH90ZMHjqdXb3gtGw3XrkHkfsudKmy8ifG5QOdoI5UUi5Bh3B/6CmrYAvkMQw5
d09UAFqs/XSmaaElo4qe4s+byl8YPzUFwmW1Gd78nRGX1TMf5h1zLkXx3LnTKDJ0
W6Na5jElSfRUI8IfQKbmSbeZ4dR/IxitktFERGan4L7V/yG0fjgQsJBODmVmNW+1
eUZqsrxceiB1v5fdHKWJ6rT3ODpEDv7c4+o1uZ+03J3lHeWVgSWZh6AVaC3K/Dw/
b4nOHyCdmHe59Q2XUfywibyuR2+ihKVHUWpZ1bemFzupHJEsG3/8SkVuxt2o8Mgd
6B6F7e3FidnofW9L3QJSoekB2Nfm/LGu0ZUVKHinuNsOpSABsbthbL3d2vv5mqes
60lnQRt+0UkTrIi5kgsbpbD70xYSRAsc9JVYZhfQnAA06296JmJzfwkR1Zec+otg
IYCDszgexuHgc+w1OeKGqtNLfZQwVBpQF1rSpaMB6x5E/D0EG2EqNa4j4L3F9BK5
QE2oieYMaeRBfCyzNOlHG4qNGe83oWQLDaYXxYgCJJfSbAqoI6zBmlnNzdXOCJM8
vicbX4+Hfbi0xdDSzKa0EZJnvC8I2v7ddG8GzYGFcwJCJURCMSNDjOGuCeYxs7Ag
6WMCGM/nEAGh6RRmCcpDn6Votw7bFkhs/BXV2BSOVZceJDutvIK1FxqgdV4Fd8FE
RPrkqTyMii7u0PcZa6g1TSFL2L8xwQMd+dcQou8AcnvFV6mq8Zgm03RLjlxZtkXi
1cJ/aXIMnRipL6IAo5oisZN0qAB1RMO0kniSFzcHd2/ZdvC+pOzw917UN9BGJ4Ii
JMjefzo0LvqcCLYdQPsVlYXCYyotbiqnl2/MNU0GldHRH1AfJRl8gSnYrPjOD5fS
el24ySvUoLQhZAAKXdyzqgZ7COgaIwEfpFyNahBXIsCvdERyus5AzRYNiobBikGV
a4Fid3gsARSOX8ohjUXbE+BWrZ/l5yTn5YkDzWXjGM1ARtUDlvYkGH7B+zdxrFNs
AeHnXmUYHkjSVrExAdYHouigwoJZte3P5ikaBNQS9Dal/tUUyLY/M8bxHuD1FS7Q
II93q5lHHsmhAw5nRo016WRrFrc89A4Jx+sds8g0IXEUgZrg1LwfHkvamvYQImMr
qamVTI3Tz5cTH9uHgNVwb3gMBfZ7V35GoYmz0/pWpf5b79rHIHBJQAFV0Z+2nfPM
kvHEqNDr/lmyN7R9FKX4vR3nJpe6x30YrLm/QqI0MOqVrnyZaaw7lTRxIeb/lDZr
ShKqqU84Jvnw3OS6wus4pZC9bKZp82hadSlF/aicDjxOeIJIlqQseXSNl7s1EduT
ZqJt8H3RPh7o2nm8rZqMfzFEu9LITchYE1cTJYeoXusCF2lRoNE84ydioEsEpNHZ
M/CQcfc/g8vs1xXW0sjJJ6xVM8TjUP0I1X1LKl5wy7JhXk0IsySvxC68ohslkjcq
3+7QNFaMok8ffdpqFQZ3H4ki8GMxRWEgC5iV/EcxM+7abiXcga+NSXAmfAIRWQyy
XpkgiIg70/v45RQ4uLY2qG46WRQfIG3riB3y6p5jqP0xziWCfwW4fsNlE+8or+Td
gJMnSZ4ipY3u2+RYZcbQUnweZcYUMVtPlniirl2shQnXINhRfL4M1DKTN7pamZy8
ZM45XO5yN4nY/OgH45lKip0G0YqrtCU9yYickrmAtzaALV+/wdOkzPX10JOAGswS
TVTcbvAt+GmmXiRijxztb+cNSJmY74xp8zBqmarhHzO1zsMuwrhzjTiVFrUiTht6
pZN6k09yRN7wtsIqINqcvyvljRoXCrG/7c+D9nw6xdxyCEr998h8iAiEb2c5AxJ8
VSzDNlopHaoi4/phQFfZPx7y5GbdOYuQrKhFAkSlUhatjWM+YP3XvkZOgLU45Uan
yGfH8YA2Y+qSMMtWd8KA6K91Oh7qTZFB7sVQUdh+MFyB+X5DdO20eWNUUgZFndmc
2bVp4JHr2fhymXv4dOClWB1/Wx4kcXDabUrvcSiUd1XqKJzC0IFomnG1Ya1kSy4E
zGWKgQ0je2sYX+uScrOTKMEWIfOvJWwNFFfbeX0uIbciDJyo28Y6cF+v/0WM4Fep
LP/tuCqR88GoLgKjqRLqFkUzhJ+wiuu93TpK3pyMyBnaWKoQPUO7CRt+VUC7HOui
sOCQ8sp1kSauHchuNYhvOncQo3ZEgbpzSTcm5hSw4HC68kxoxWYB5ieF0KQwt4fx
NsQ/CFXJM7Wi4AwMVpGpQHhbb2+ie605XHgHabyVCBI84bp4bWKdb9p11Ly9aa5B
Mz4MRNTjZRLrwSTuZCMTORSzv66WcPoVzEB3sfHlWuSVRgu0uW9AQLheagSPceD8
hks+KjFzCkP8KQDnJj1SfUkfNJQZaVVqjEy2KPQBZm/sDq/JAnI4hHJAI5FDl5qC
hchfvpGobAiykJ2KZBvfkHSjeC/gnb/SIJ9PFvG6TkjnwmYLtsFqoxswomZiL4rX
PnuHXcsBl5JtFTrVClLYlXV+T1e1YDMWWqm1q4PpJtg6QTmA5jp2YBgg7f+MMyhv
Ej/yNvgbfSa1yqqUj04TBgFrIqdW2H2p6//0V/CB9M2kBTp9x8H5o9JVXE4uwoIo
WbXlC6IcDowzqvOwsqaVG7LLa1wgURi/lh264DBeB7a2JemT5N5+fAUvH1Det9F3
nuMhE0Faw5tb4M+PVzMwQLXBoWNBfZMXDIJH7oJ6bgAUqKQFlHbjbIPQlFyDhiA1
VzUoSenH/Whs2zs8kPMspsAeRjCz6dhWF7lFYMLNGc1U8zAK1yQc9dGVHn8M2nAr
FurgBNN0d0v9K5cJm28+k1HHSjViRVCJyjMuihhtgkfl3XSt6u0mR3EmyWiqsxfE
HZV0nL95Sd9lFslXXI81uEHy/I+MFdmEAZjxolMYb5uSRRiO53Or148V2GEuWGdG
e3Wxt99trYHEOgrgLiun1wkWZ6FTBmDFJUX6fnxFuunlWOKmUvQoDAA1lLjLyYnj
Wa9V3L9fnSzt3qrhayDMOLYkgBGVrkTFDtm7nOBc0cApCmLwKMmAQ3n7UWRQGU5O
+yTNbZZT4pUAC2naDsamDGD3B13ryOpScSFIfZqkUQBOtaE2BvFlFUg69yQ+jJy3
8WSOncSspHbi0BEeGg8jmU+nfwTdGosBZfVZXebk/AZPRYR6m0rVP+l7nS1iJtdK
JgKnUSjmS4UFUBHDYD79fICYwM91SLac+ZtJDsvkQyhny1vmdHS44PfixW3qNFgi
YSbaj4rklhnNtiqAl8DCQ7XUIEms6gC7038RMRdQ0u5qRTkOa5OE/y2RECJW2wyp
A0OvW8e1CnrJ84U2jL0BQw7SSy1n3Nn5jzKGrUWgAEh0xhrc2/mXXm8Ehf6I6pFH
i+bocfY2eD30AQ+mOqxSncmpuUyXVjBIy98dZCPVXxuaB9jHrDeuDbpBiI8a2bcs
59Ne3jN9nM5nfRUvSFh5i7RcEBiLob17zz0JFMdJ4N33UL3IR4SUBWxMToXIM9mS
hjC9NIJoSQ/i2AKVX6qrCB6wqmGCYGMeVNvxfuP42UzerUUCaXAiqBbWZvhO+Pu3
+mYf6A8kuM8VXeOGGtPH0b8OWPOY19fiIlvnOcFP4rqW95MSymuSxQBtxDL29Lph
847Qx+yS4Fj4MOxnnVO69V7pctJXNhkg7J/MbxmmabqxTzA1uzGRsXRrQY8qLfLF
80aSl3t8sbDAkQbje1oaI0jSxh4xuM3gfYJWaBXAx83PjEbLwocM8L+IRir/wCkU
8aguTppqntflnpFCWqe8DMBMHby1ftWVI8/ZpTN6U3H2YEyQHFTSMPnQRytI3aLM
EYvTpYzVu+/EXcL5eGVTuXj0VtolGZUEjv7T52YajpAGf7u1Uregqg8KCs8MqXzz
Mg0329vTDqdfSLx2d7izn0Q9unA4mDaFPuK+JzNmTAzOlGH/2h9Q4fIQj/yVpogh
Q5f5xjnzFbCwEw/2UOOjNAXf8zsTWiY4Nq8vnCnBaWV7v6j8AOz6yks6LoAHiKlc
yd/0IwA+zTkqDKnnbJZWcQlA727NFJCV1jNPKQyO/s65Yhk7DLshPDuKw3UTak/k
vANEs2rJ9DCh6y/1V81jOPxJoBRSDiG4LAd9m8Dq4r+pbdZ6A6BbohuWERFbgtxx
rx2AjVLK2r5ygHvtJdoO2EELkwqlDMXt4vI0BU98hiIqU0if65/RZA+xo7em05GJ
ucTX0dTlboKdyNRgn5oL7dQhA7Wjlx+rnGTSgtr9nx6TIrmBFTWjVNl1C+GXdSG+
nLuNPjaizboF/EP5AHyu7EBuCmSo7d2xUorVj8WLkcehRM3HLIRKEaD1dLQiOlz8
k8TntfubCTnMy6sbYERLGfzjz9OCmMCyLQNrl0FhEBuW5xHdd16JKAC+vs1HVt4P
+sli3Bsy3o9JY8agSx+gCob+Jf/cQM+8VR/u4N8tmxF3LxIQUJUy0ZALbH0crOhH
SHfvTk1fHPzlxLdWeTZVIioHcFYO/R5y9uXofF0HA8V5vxEjmhuMyDQmb+kTTSJz
JkQNY2t3tqdszE0CrONW+7ToaREqMJwYFN+1g0ZkkV+ZU42xRAinW/EaayDok8th
lECbg1wDXO+JkwWs9jBgEp97ryDJA2d//+NeTvPOzI6omJry4VcsyK46oOZCCUO+
RqYKThVGT1lk3bq8e8yRL5yhCdqEyjJBC/Ipe5CG1eHqDSQzgjSzBk9FUN9SWW1J
Gj3LY/HP/WqKLShfGIfLLMYwUiiEEOpUNUk4vQkdF/5mG81DP/0dOJ38CMVRvOaP
JhEkGZNJr5ENOej09eFnd57MlEQ4/z0qxiWQRuObp2lZ3PaxJ8vsdSZc8OfXSw08
+da3+AHgC67a2f0Rp96fdhib+3qgbWTupVK3LiD+Te6WWG+DOlJDAMzNSOjMWD9b
3gS6sXcnZCYk7oV2qfDmyRFoA1iRSiop2U5yYpthyxvpkTRO/To8lZsrNfFHGly0
yKOthgvufvjnFo8i5Gh7w9f5oofonJ6WhmA9Bh0M4ZYGot1tRXGlTcY7ffUwz23t
TtG3MeLA4XR3CUJrOo757gULfHDlhbL/LUAcoTOlhPIWIidgbCt/NljY89xTlI1R
sVtYDgRuLr7qk54Sx9M4xRv+JCLXBrZrMo1wFGOhJEoH4MbEwZaJjUsag+bKmc9y
zmwpz9oWMKAgitTa4hCC3lxgpLgoLikgdFcscZ0WT0HafmxkZhgJaSPaiLn8Hkz1
RSCt0b2wxjdVojubXEsWupxZ41dh+kO1Gy7aXL+7nWT2DPrrQc7IsyvLkuAY65ZV
f46H4PM3ro/8Yyssv62KbXHVUuSBgc4N9mZqkhA9mvVrdHJK4XovPDk+I8UntriC
8lZWd3bPvJujh5jQdfDdzJ+HyYKlTxywiq1ap4C7oGZINDw29+1DMqkeixAUaiDL
O6JaRQfxMEaH3x3oduARQV0+Yy0cEPzUB40o2U++WVXRBzL1Su6YbdK4AIqUjnas
qUtNrZRZOKpwRJTasIDagJliHXUTFAwRk5djKWyBvLTa4EiqGFCwQP6/OKsASD0U
SgFxnDwvV9VialMVOyiumv6HaM3altg6hJIFCn6wZQi+AEV4J5FOc44Mnlzv+i79
GLqhoZjh87hdkEWyc1U6tcPBWgTMAm1ve+jlXluoDXo95N59+qUPWWwxQ1HdbGT8
T2utqDoMTqhywxXHH5+gQd4F5AoECFQGIcsFezlTr4jdmcFa8S8ZkkJD5FegJQpw
P4Rw26tDY6xMuSF0Ic03Xd7jAxaXNJMd4K674MseAhsmnr+3VRQZWHIojGSssIfo
sWcxRkcJVj3zWq2rNXxYGmPHae3YmRKdyVgYUV9u5i2WSFpV/vQzTGnW0265LIRr
IquLEwiLYZNFkWxHLwSunWGstqbp1rNoFTgHwjIZv68ntPNTSPma6V/DR6nRuCvJ
90bdg8bWuc8Ws5AugzQjZ7rVVw1hMPac64vPq7FdR/yc/gwqbVQcNrgUy88MegGc
39C5PUo2MiiUs+CnBgOVPSe90Vbfzd4XmUHuR8gPwThiHYDDyr2JvLI1BWtfzbw4
NROLW6h6A0igz8Fy2GivLx4i4TfjFxaG2yDtC535oz0iZdKZJUCf0fhKxplUGgmM
fq+pU5E36R+hsK8OnWmBTHLfSm79mp99lyfC+6CMyhopFn22PF8ycdyKJBFgW6PC
L6VZhbVhy/91qayEV1sYiBrY7enYbP5ZhLvB+XHKWG58AOBrnoB1HUCEJi04d/Uc
QxhXBgA2i5biJavkkdVqkh/ozJfcVIy6ySxh/gspaDmKQiyKBkt+Tz61Y2LSfnhe
Uxam7p4vHvhVWQsCeF2m0fbBxAZghkEvdlxRBsrXDaaYZt6va1GCs0sX9fzCNIVC
Mp0KFQDe4d4p1Gy3GmrnDd4XBXAFWzuCPpjSV4IdvjouuHvqTsdlZ+vNgqk133tK
opeMmSdKoa/E07tUoGtk7Umb0RWixoBWUJbQ1aBm58Wkz2oR7WPdYhz54IyaESKe
OIV3h4VKdfrOMyf43kcpxfN7ChXeWcTAKCIwgPdsKigcVmU78mJcK2dm+stLtDSh
v8m6nZ/iRAiEl05fvfjp87ZSy/c6WoP4lZXSh0nkANG3cTIkm1DSXbNjTMQnF24L
53k16AonwHIqqNPoA5nqzGmifVRhS1iBvLbB5TEISYzkh8oqYJ7nYAvaKtLEQt1W
urnyXGnYPBFNF7fnElleCWGvIufdoL6tz0El42vudVw3AeRgKSRQYl0PcUFZZKwH
kzMcjJ5t+VDnhkoI8RNpTH7Xc/vuEXWKPbMRMYO5D4+ApOBnOB/xmQgh8kIQFJZB
2eYoGqSx1IHqW/giQK0b2J98xzYZp88UruhTkdCCQXJ1IL7TCOo/qmCKFe/4PDjm
AEDsc0kVY5BtMbqEcMcEF+3qr0sAK7o2C2MovKlfxcTm7laMmhl5XzAl5PFGKHlJ
11kKig40VRnt3caeaszSVq62H0kZzEeSTh2BaxiuAaFBwQq9cUMbi7RwGes6VCbp
2MSUD1kREa47G1u/rwajYCHiEPrRDMDyyc4b8y/b4ceF5Dgyc5Zve/74QpzaruUY
9sjRQbvshANb7zezbGhuMspFpUsPqsmziZovIEFz4odyyfKyaJClrXzp/qF5NGc9
RKN6SUMLWN5wwZtuKAvZkH3Ds4yGVJ6gdM9rdKH1hADU6Vv4CrUnNnfJ9gqMxnI1
+KLFHtNXEMPxtrCYoelkkxt5zUkDrCCQ7WkZMukY6U2kE0MNqBKuyF5ozUJsiuxg
TrHj/pg7p5OuSpTXc+nKdv6TwO5x5AJyojaq1oVCRPfredAw7PG1pXmZh4OHQ2pD
UJXtYcooCqyQOqPdQX18rmFqYLDdSjoz6Ci6jLtUkSTE7TwdpHa4tPnDRJCvGZz6
R/SUJGCyDqZr3qFqwGaXD2j3Bha5wAcKF+UFhcSqkTpQio/yzJoWPKgZ+8ptp3U1
TgDRWlkER3wL0a3rf5FKsYGqPgakCEN1OPtaj+ug45K7RJFFWA1tVuvUFDVrki2n
EMT3PYXyyGVVjrmehUqkOjDoJ83Rd0s1w484bRLJSgvHn5Gv/GR38ShDIag5OWdl
elJbj63NvxFwa4ZH4zHEjCQH63kr9H/BeiEwP3V+D126u9IjGlmtNkgmcBkbYTgq
yq/VpCuc9QXCVnE0UWooOwn0bCFJyyj8Ha1umPNIluu4OMpmkT1Lt8/w4YJEfb9P
2+SPWifGhqBAV+2+ASDDFmG+aNkVmV7j2zZQ8EupoWRt0YF6Ze94uPib32/A8V3G
tpYu6Oa7kq2FHDaynG9wgqcWFmFWMzMWkXP3LxhX22ZHPCdsZWRvKsj+9HRp1ly2
v9+ab7aax0HQPmBn7/CKzac6Gh2jBbQPmxPzqcU6tC9iow9cFdbEYwVTXY/+sgWa
yz9GVZZmPqPsJpOD4T8MM0kBicLHz3XaymVs/mlB8kbC8lnhzYZsZUovZimiY4b1
LqVWDMVlJpuhhCQUxtPy1KRm74ATbbO2q2PvTnJLktc1lqgOpih9P+mPPqFNtlTS
uORxJuK1/dojnOr/qAWaVTjjHimHvk6+hqPsaE52oTqKssIOp3Qyk1PZYBqJSgp7
ea3fTu73u0uHQzvp9Xt04MXRUXm/fx3k8+sWg3WaxTw73jeNAG/6QthMSB4G6jv0
q/+gn4mNNGfTyYfimkAKcyv/q8xj8n/cbm9ytEEhCDLSFz369jQFg2cSMOwjkpi9
cAbSQbai1lisfHwRHTag2Azo6KS5kCkbX9IaLF0HuFBZT05uDiEsjt2eGekxNbD8
jzKby0IQVMy4dNGzzaQFpQh4Z9XnrCvAiT1aHP23yFAvUJ2NaMmUCjhuBwL05oNr
+vYKliLwc5UnUxEyffeDDLV+vONuQneUHYNQZc3Ru9Ht7bRLRoKUmsrG0n5F8Fy+
ec4DB7oyFSLeJIBTiD/DjiLjdJHVHnMYShDGn26lKAHqRSeMzL6cF42B4fwTWAU2
jKWJJVORdnm0PEc3CsVJgh6OlyJ97ehkfRKRSQBpnsRUJKAQ7AaiS59K23r9N7RR
vGfSWdSAtsImgfK8+kxFHRsddyV/U6zi3ENYwhPTIWlC2Mjy4skW3l1R997Mioaq
hLXZYHk6vtDf7vRmaP/RHooiSsyOR0ydeT9eVj/Q3C03MMMEoO/YNEqpYLtqcHie
5K4VubSxtLPiUNnJ0yUogLhxuLspklupesEuJl3s7XFR8mopmCZNHMmV/EgDcUIz
tZJiIjCKS4m2+zxTBAwNT6PXdUkKCJuWfa2MV090GIu0SQxPnpb7I7uKt/ImRRni
E/USjulPoHAJc2ADhEuP/vorbO1gyS5amj4wii7wtcwF6TMuQ9dcbqShli3RjvGd
Z6tpL7RpNYi/+ZQg3eW/FrZPVnICO6le7j5QdcqE8ypndE/2nQ+s0sLK3LeMNpmP
PNeZ144raHti4VOw+P5bXJoZFTZvnyMF0RfYx8mU3I9Xshho+5BnH62kEsL2aEPU
iVxjXAdFpYQ5tEZCVCjMbClSWLARqPIPK45kwnB5E4Ql9k7alKIOMA20CWA1a/5q
oS6UMudtqBzKkQxvMaMaY097bnxAvCaP+OIc6K/RLYVk8Svlr5mhEjjZN+jY6mjy
PnzEtRXF3WFeWnnigs0MuAeEAJFza2ol36x+GZ9a16K6d+MuvJPvm+tO03FVKkAv
atk4GrVZvomlVjmmx0FFoYRz7VzRtl2A2mvB6LYOFKebpjAYm42clTAIoATIf0jU
syk3x2j6s9Y7mvGudINe/HO//ceKJYIuoMUgWlMHwP0/zXYixLMlOO0bk53GQ9TQ
rxEPAoAfXHQgksTVnxBBQ7/N96VvV+slzmrXukmmM25TbJFVnP2o84N4TZJ85HHL
meEcbXoIe3ju83YdeAF6adJqti6b12sOi0lNJJa9104J3dC5mxkc4ri9q4tFRnpy
LOSEnAXVJHmNKbGAQsH8SivW60xKFJnLZpTko4BQ7X/cY6nvqfQKg2gboiVV/m8g
k21XorY8HgMnecI+wNqyxFhcOV10VHO01uU5UKZD84lASWnkAjiHRx351agtvJL7
Mc62NaNCUQTNJxZTQYPC5OVGFijys4hwtV+4X2I4tgUgY4msfiecESq5A7nhSGPV
jbdict+UgDnI9LWoWysVlgufgl3mKhET4EJdKRcA6OIEvQp9Dulf3kLKYvvjziGF
teJG5lX092BEm0fqZSQE4Bpue3zQL0L0Ur2ZITnYCPnyscUUeLM1GKjwR0ZH7fdm
+nGy3hE68gorObmUXxmkxFShM46IgBrNxBbcyy2qWeQiRHHh5QckZN2NrVsLdVJz
LHjQYJs1PnYsPhaApwOyQxrwiRbHl9DvujfG04capdi1tPMtiJ+lfaXijQrBuZeY
LNzDITeSntpMrcPaDqCOC33lHO5w6WptxMlZK5eOMc+3xXmhf2A6s1hn3DnSxXrQ
Op2p9U5FukWU62acpyWprzGy18dL+CT1wA7DnuCgBm1Ph8QwvsazsSQ/AdoAuuSR
hacdbDyMvTwOYdPeqCwse5CSyPFzNG6SBAri06WjSUh1H7zkjyGyZC6rsYyAYFy0
3/N6CQuRGCQGzC4HNsepL4+cDwrWx9sEIo+zbxlMmNfP/6FJyCLdkTIKPHuH+kIY
tQuW5JDgtF5QBKqqTLsThIU+GmB8bC2mU98nWAO67GcMM7vdqPV3tBdrr00fPt8S
qFe7f8QI3tMI9qx/yuU9F3OZ1nj/5B3jK5cmrj2jO4jklA565lXugkTwzoMWvkJ5
Y6ca2VQhTLcFw4wSURLdMBVR1kO7vpzWfBEuVuy9vS4A7msvOMwajJqEBP7cVWUc
0d2SXPcaDhQ86n1cRsswfxvcQ4zezWqvimVTcEgn8AWfyam3tysnImy68/d1+Ydh
eY3whmvCAFzumJvysC9Xzs67RlIRxfSDmRtKWaj7KUCtU6IRYnDLZz2fvgS7hFkb
CTbKryGN2DLTqdVta/MSw1Y2rAQsFiS/53Oq1DR62xw6U1WLl18eu1ae5MGV31p1
7zflahZEJc9HWs1K0xLRGyZSC0UKJ4SQUAJ+V/8FJACWztSqv48Osa8/QDqBxA5h
yvcOWKg2EDIeMwZDuQ9uLhjFUvSY0w3discTAIibseNCxpuS82Fj+gIxOn1GH3vy
GeuGz8IfPuOIfhj8AwSRs/nIRxfSRkKf3xt4wqhqgXJDUmIxZfK2he7M+1zBIE6y
g0tZlnjeBPPdNngLRuX6Xogj6wgbdB4Lu03h0b96AN9p+iYxpWbqO5tP+uNHtoxx
l1fRJERbowqWPTDotaJDvQbl7HJFfBPTBjXlxQxjLYA9FdON/GX5D+SpZqTHChAj
Rd0JUYycWw7xqcYaJFBr20CblPihLmaAeVVsIwCjjYrbDHtVqfJOSBgRgZMeZGXj
qgL3xYasmc/jejB4xPy8CdZeP2aNuhguPQrH43i0CxRJf6OMH+Iz13t/jfU5zhd8
YEP0B992OtJ8Ozz8KTZnXLj5DMSW9niMKwy7U/Fi1ne/fE43IWznWu4zabXNaQbR
3L34kOrinDZ6qc92jP96mg7p6R0gaWe7rJKCum7imLPzZy+L9ac2ujlWQ0UPoC3Y
RhL1tk15O4t+LlLIcqfOGNQpSNQkj++1pDV4AHnJ4n+FF2SX6dy5/YqSeBH0Im/l
GoOor8jf8iTUjv1IvTiL1zaMwkQgqEOGe7vmCqFtlAHGM80glR9WbCxNsh/xxJER
ztXVToamnwX/dGuV1t1lCFMNiWyJB5CDmd53si+rK3D9xiNtNRxqC0o2mzapUvps
8KN6XKX8j0z1VnAWqcb81eDyP+PuFh3xursvsSoRrwEqLm0S5sqT++dPbM8kNIA+
31WFnSCCytjMrg2+tCFZmgWMkJ23N/zjXGscXDvDqg7axya+EQ9ByF+z6gpFjIYn
KVltFhaz9VFJ2FnmsF6/KRfRCb2/zUPhwmSSzTppl8gij6vyeAVbUz2fegto86OR
wXZcnlI19Z+G1KgYiI+vC49Ipl9XHPV7mGFLx9F0nAOG7gkZOp0lDCNqbwlB575x
lE7R4V2uE0cdC/92Ufbf9aIexAUuKJw7Jdy7v2VgC3+p792BFbETOmBLCZWCNTGU
8Y9Wxp4+pKC8P1fZEDfTDvVbwoWWhwCj+ZRW2FUUKqCbPoUWansnME0X51yeANWU
EPUlHnF31QyUKUwiN1oBoxhtqMHW2J3sjkfathtBy0pP948Y5WBC4+xKILQDswIk
Ev4F0h3+OmLPSqojTFo30jjwpMuIp4S3CqTH18O4Lq7WN5TJ9cZgL5uRG6V0Code
Va/KFTnXd4MYpgvrvVSSzYwoZq19EDpXEUdY4u8tNSmu3ThTqCWbePgZFIHbgsvu
Qd7cUEAT4oTgVvxWG3rpFUBPSHaJqWf5vcJzeFCc1YSxU69zvCoadbwl0iWGZOXc
ggLQbZkriWD/JYNE2cmF2tXFQo3HH2IUBQJqWiCwjuIYdRTwRtiZVeUgq6luFh8n
9GL8SnesTyVqeh4g1Eypz6PfO3zqYgj6UfexRe2Ix5YpCx4IGxVObQGxHHwul1/M
1lbxBKJemvBpLnsqTFuLyQhuvnWgjvu8521NH5G26F5lXjy093JD5BvbnMJ//8Nm
aogevN9i+xboPMoKH04DvjELDfeN90OMQydAZcuBNHXH44Af/nTGcfLqrQlhGjlR
pPhKO23KPbcKlvP7We5ms3zUWjCl+alSwhXJIKgfJ8IB8R89jhS+dYnzBHsATw4B
7O5Je2OMdeJkx1k7WE/3i67TyH10CM4/AEV2XwfY7mVKe49Gq1JNGZ4ag8K0no3N
6U5cX0zAd9AUirPj/ii/vu04m2BSlz0mobccVCdp1oKkTvgwzeWlLDsQWSj6BriW
INULbX2QDtl/9Z7Suk+JSu5axYMMjTWfublaIEqjQZANlUqbqxAGkHqUo/PDC+l9
N5UK8eh+QeicamPq/6+hWXuwzpedtoMnGnHH6DxNYawVS4hB44Uai2kTyBWQPyle
Wt7Sanm0D2U1A6nZS2Ts4WncCrhE3jDS9hwbceHabSidoHEG3AyDBzzgJzn0r1uq
7oP+UReHWNtqnnLcyr4MEz2lDsLau+UcsEZheXBvGrA/q3ATstSRgh7kQHhBuNT4
Nw+fm4wnk7oGYQvhTtssEOWUEOiYJk0O4qx9E2XQ3vIok5uDQ09H0fKUgbu2GGBE
NKvAt0AsgNLLBSYYpZp9VH82pt+4nrptURFj7FeXjR2zVYKLx//cyo0vuv3V+6V9
alkZcmcD2X+C5pcbvvaNvWFYRNebaVB/pbh8reL3hYFKvZ9i0yb0vElJN8kHi8QA
LCrdcGtafdpsHlC/Ra/vGXRtUY06oqjgwCnt7FKK6kt147l/GPAipvsysp84QT86
yVq9GAz7/++AxftYTjlTSkg8OR6gY0V8WIrykZveUQLX7sbmxwVcFMo5W5+9I9GE
GPInKMAslPYyqOxNtzxXtzVo9jUTZPLE2SqDFcE1NChuMfh4VOqyI5+l4GAZDiVY
joBk3h0xcNIt3225gqrAl9LdvKJTDEGNZnJTFyDQgXGeNRStzAGO1xWF4mF0mAC+
oenOPITTWcXDmFQXIRf/OPH+3rWBhsicSUtkKMFyH8aCNP4egxNXelZrrP8pwoXE
KXwAzswECN0ym+TThMWSgha96+Db/C5GU/mo92e7oBMJtvagtviEojX7Ukv/23RU
DcvTfcMwta6X4HSmYQPCYEP8dWX3+UhODDp1nBvZIKeOUxPvRk6SES5ejib+0Ile
hCGyExJhsS6rGVwDZafwXx7JI0Hc2QUNNS5bX6Wfnp71cZzLw6ouj7oKO2uv48W0
ZyoV7RZCrqVJvs8AU7mGeMka7uMq55YJ3DtP7d0hxDYN0jo1uX+8z1gIzQFyhGR9
VUR2r6HoEwvUEODyB/KKz0RgOKoqRNXkqeCzW60seYAeG9FL1LMDDY7p53sBtiR/
Z8Oenb8IuHpfYct2N/9r8xu8OYLJA04C9lFlHfIo/Oiju14h4RW8kWCaLnByvZcK
T6GKs3cfFW+yLMxPgI4AnWSF78Hkqu9s/01BrGSwPASQgwWpRfvhX5yp4hR87PBF
GgOb9TSxWANA/isa/u/ONpTS4L1aTbaSFBf9uEAgdAutJFz4PxOchUnPX9DI6wmJ
OIEwYSMzZHES9BOFYZhxgBWxJQ3cSua3ElT8hUgBRyaKMk1L16CiIQgaiHXNF/+g
ZGBiWRFhML4BHAW3aZs2rogrOZKg5wOWhGqAlRZFRgAiTprBU7L9ly2sakvYZ2Au
KhTpJafViHYJ17eePvXIWY+37QKHvrnNt+Uz9Rj/Basi0Nlz8Cy1hLHm4n4zXUx0
QcF10xRuOtR8B9hzAsC7ztBTbt1IUTFM0A4CNG7EqQKQjYKGi5RKJWgSrEAz2GEl
Rw06s/+2WsOgMeUbf/OE5y6A97gu0PN3tVQrGhTNqTzAqr+rzctegwpW8wJCP34v
Si6AaX7ZScEMqaAQ/5ancAa5981V+asVYb97Yi6hJb4WX6lWTYoAy44hWpVSEgQ/
P9z2d4uPAv7bMx4CADV2fZtNwa2M7WFLW92s5gimFy+XadKr/3W7QebCmO1k9YKP
BWQyzXMiyj1lM6xUbJmK60Ar7S+rIRwYbNNADyB3/Xh8negX5AoWCY3WnJAYBRLM
JNOP4rMOGZgxjDHPJtjg78EoV4C/w7hlNbC/kqh1Q84uvpNEQSe5PBlDTAVNX6Wb
HMd9zIVMBU3AsB280l7uHrQUZ3K01sFAvXZp5eL7Tfzc2FI1R1FAp8CdFaw72H6U
4Bvof7tW29Jb2BrEGu74YfEO3NhSElAeUbbDKWi4aTIYsmHiJLwYZbWNWqsv7zgB
PKMFpLzN3We7TqhTqYf+OnWzD4q4QogbeBYwWmny7m5f60v7u/Wkdci0oORHPyqL
DhxifkpfAekqkOlSeGjSjX/ItyMu7l5FwtFdPzO3Sh1lHG/dbBcZ5oWEbrsedJcB
RMLiQBAPGQAla3UyYvUaD3lIum+ZMx4TCFye6nGZNeOOgtTqvQXHA7CVzPMohCFC
tC2sKP3kUNPepO3n2ssxYrb9X/X1EVxWUi3gtaeTRKXpYwWJXjiK4sf1V0AnYRji
fS8I0HgxzmQpGK94Se87+IzBzJKKdzbtzghEkqjl1YbIHKlXFIE4J4agnvAIHH3B
sbjr3/G4LUu8jCAal346943wu/GbmNXlzd7pVMpFKMwkB+uIqVEh9LJg2NMvvuUV
T39vtQbuDXvaZ8yr1LPIl+d8NwFvwq8QUXmmXZYh1/ksDt5qM1zXhgfq66kWUQFG
QDekpF2VpmyQpIbx/nKZuV5gXpLVRhEuiyHK+mg/+vbFakKLL5UFGCduU/vh1Jnq
+Wxwtn+9kzZlcnJGUw4mZtQ02KsoaupU9bSZgXOsmcdKr+F5nphheaI9amUPbz0e
HyE9WGNGX2v0/7No/4ECXgX+QupyoRiAuT+dgP5ulfsh/ZXiU3dPwCwWZVtSMsqi
5D2K2UL6uLB2uGXal0cXbvYI8nlKkZ9DjTZUz6eyXdt7eEY29P83gR2YayqQ1h/b
ypi/NeIEjUYF/hvcS97pDI4dRzLKlD1YPAbq/SEuMlxjDu1QIsifYtryFADv843+
/DAbpT8O6Vdb0FevJwBTXQpnu7l4hy4mdpY9sD4+a2lTRYEtdts0RsJ0x2hrMH0v
lWDPiXCBs9zIso2eHix/gVQEOD7lPGKepyHdu5DPUqKjs4zi8r250S1/MxIllQWN
uxiRpmkKB1q8WBXlzlLnvk9yHR/VdUye7li+hrcq8DOL7i+qBPPaTeMvJD/ZbmNO
y1C2AFhENuRI+YumspjmLxKqB13v9hdWgfcVWr1qXLpnNu4PGEr3fTNOuk3eNhXv
Yl1USLctXhsDTMwpUTngTbJWC8pVYcd5KgsWMk46ldSZB1hjLlwpPnmiBvP6xeY8
lFF4sd0x4inh6t6vTVSSEproLU72iDN3QxOrhgu+5bfwUaAO2JcQGiATHS/trgna
w+oeEFgbSwAvA6hIoPnsfCpwRFfWUZCYGbhqO7FSG5J4LzZfIph6+/vslZS1sWeZ
4Yhw6hGRPLdHppVlK7kJvfuuAFDQli2a5MIvn8xsKlfrKc8VGweivGdqy83jBOmm
qkXH05hfROWYc0iMFoN9CRPYb66gXWXDn2G6HiL8Q+rkUe7CPpnCwgbeWPSEOqJn
+1vUR13btEG7+NvD1kvf1Ry8gUvE2p5UKkJkW/OD7Ri78ygsLAMGCWe0lmWteKqa
fGiBwM5YT5ZeaeFK9hFmOA++LiyMkto4cIty/qICHnLC3IN6Pgve0+ND8LGSIWQ0
bPJvbxZn0QWDYkoFp3FVKnhPbcQTpsYNWln5Y8JzkFRtISmZrtYAlcjczGBlmLag
RS7IBeZlwLpB3GM0IUIG5ptYB3PvjugveFi+nmjIzEJ+ZGFM9got3sfsRWuO7QSn
04JIknHC99p44V0NLX6rkrUx4Ll39jjwrc7WjQVoq4LjfszKXEeRbFYDSZK6w8+B
8LvDnsjDH2evkawPhPRU7Zz3hmzm/vBhRzNbnHOt0Zpk8GWUrYr/9AF8+3NwaB5A
TnFSYclxEdtxtBJGCjYgkvCKehSYBm70k3bnl34+okTOnpwuD8nRix/P83eO08Jf
KSvZoxTExnxoO0aJES801BE7rGG8bBXKsHanzPbCQTOE+WOWmkYVJSfY5GLcQBzv
7qBKARqONdiyDkVr3Wg4A7CMIwnRfHT25seRwPjg9zWwAf5gyDbporh0FPhdFuyc
1+lcrmUbMYmgVlFtHOUK0zVy8wD54zXjlowWKisNvnMb7C52JClckI1nDJ3oqLq3
jDWxgN7MOMvYYBfQwbe4VNduGCotOIANmC1T8tMhP9Si70PpnLiY0J8nShPIc0JA
YvsxmYg9BTY+fugFtDF1P4lXfdVqOL36x9q0/WYvnyGGMMsFIOsRyHfl8qYjhznW
g1bq3CPY9Tz3gdp/MUj/VbyNISKhJn8TfLRvpHlQkRuSo+ZCnG1WwEx2URnEzeb9
k8Jui3qqAzlCWOu8O8YfXko0tE5/X+6CwK2blCBthqI8SSbxXz4LiyV78rzhflKZ
FYLfAs1ICX8qfpyY5XPXWLpmIwYOgJfxKDPueMht89M41jS/6e7NIy05p2Y/iRCd
ExQC7lXZfbca1r7N5sE2/RLXcE/VlP4wItk8jHTx1bEK9cwRCjS0pvfN/I4QaISA
tsyskj561j8+olP9JWEo5VS0eTuUdtiJklwb1KOSXPVmwbqavFwDQW6hpOfNjLhu
h8U/paO9bguCflcjicVHZZ9aJreV08VYHXHvF4waVkX3NH2yI2EVcoZEAhAADGMz
eTXGOhj6bV+ABh1rouTYVZCducZw2hLmICdhGqNupy5ax3Bg4VJfqGw3ZfIAfsP9
7qmErDpJF3gmF9EP+ByKQff86SQ1I3cbg91nnrF/w+I9r5Th7pRX93ariLYnqs8D
Hw9sWCYkmDT5Ci5A8RJCtEzp4jsbuA2zoHicDZ9UAz5qfIDvqpjzFZRnQTtCC/JH
LkQKjUXFDOHczJjs4yNhKq5M/ThPdqRmhGeiqDRlt8E2mgQYOpzNRWfuAbCZ3Wl+
FS0wgqrobnQWzE+tAtjd/ghObF1VBQUBQ8/NQf9erd6yTaygY1c4Bp4nUHmuz6lG
5liAP7GtWo08bScLDHNZPem83J4zKGyiOm+ZPqZER2jnGXg8Uwsq1m54NgJ4b2kH
kvoeY3W0q3vrpAcweDYxAPcfzRpi90T5mY52BladUJXqiSdUPmEflIWC9DNeCi7G
bylqhmiaBZ7lrK6ouGbyoG4qJDSBPcawazZa0vAt+7hgyz3xGwp5hieqgqUJiJ/P
33kGi5uvQI698KBpmhWWY2bYs8s4FuPtapROHS8SeInuNBSsuZTKt9UdtmahOdCa
+8GQW6CLs6I/QA6pg2pehaCV4N+2Rm5lY4YJMe4QtHp0h28neikNo+aLB/miK+xk
0omhn3NI9SL/OSNVegWMGiheTWVcWyP1SMFNxHwCgNZ+bkHx1eOOSHPIBI4u/jeh
dKiGeNIG4jVQgx2v+bL6bYbBdQQv0+5+RrFc/FY5c6dfWdVtmGsEms0iX67g5yIb
OZh/pbn5RboRoCftlyUG1hJlq+8Xe503uPbsLhNLlDX4Te7+2Vh4qPhoVkoCK4wq
cFw13XGou7gxOTpi/576k18X65zdLXX9BSx+tJ85UwtB9nY6jSEwNic6JRJ+pKex
N4LzsXvgkJt8cBdetuKxzSHsL8vqPcl411t+Ef90eypbY+eY7BEcyn/3WU0RazqL
l9nDNFFjkoc/+M5E1C4B+O/9v+BhdJiuHQa+30ZoUhLq+K6NEeO/JcJZURG+tnTV
VveT+68bLMv1kbOiEZUu75Y9F8/hQgihWsYch8GoVmTgyACiE2soUqRTsdENXGTd
rUSP8onFjv7Joyj7ryGIYqxpl5UZBcXiYfH1QiatgBWXgOuPpx5aERaoIZqVuB7C
iNvHV9Awx0n7bW9+faWI5aBsumoKw+dK0K0zkBRSHU7KZqwcmvLZtKFUanbIEQUF
WyDb+4JmhimYL5Oery2nlnzwA6kM2lyfEjvBVib0hrlWvTe8Kqxq+63XxkZ96ozc
MqJ7sQXyGJZPsYzTmh7Tg1fgUbHp5LtcNcXcJYHhx3VifBVy+TUKWqaC/NPnBoSg
Er6HyskPRGW9yqYwCkjViWJK4+bwu6TlV71ERn8uNMACAawFOCpM0Ph/Mz+sC//d
vX3anGkiFEWJ1W2YP1ndO07Gc1weLxVI1+Dcm7fovGB/q5V8fxIUQb/58BA2JYov
mq/8d3chUzpJCnpJL7CumR28A2wX4nEm3AZ1yILZYg//fYuyiL2Q9SzXh1EncHsH
xmlqQpNJzGKPm4I8aMKsCbLvLVTjljSbvibx0+rTbg+HsPD8Uv57EGeHA8XO0tzP
CdYHjUkrGP8JNMFPTzOnXrmLEJsdFjud+ExGaS1DwRLVg8vqCiSn/3HfAC2kJdyV
Ow3Ie85DKfTtbfYtGpXU9HeUL3tJuz4uX4/VIYJO7/xOZLhE7svBU2m/oT+PApdz
3WhU17q8lkDv7FaTBxbOqjia4WbmlS6DLNT4AgzNavbTWJfsyez+V2aZE7LU8QIB
tHr8YOTYohh656NFwisPZbfhIPjndgfaQNyU8VksBcjY53VTAQlEomnfCAl6s4o1
rLlFgPJd4eB8TkLYGovhqewbeTd1A2Nk6BxSqOCcANpgB5QUjqvWmltXnAsoA+db
xK262mmeM2LLRdkzA4i6eGxTR4YH9zXHNvf5Vgjlnm2NATOrV3a56MS0meZ9uUCB
ErD12evMskONZcCgQcaPbcba9vO2PYXAnN/veAzypsGO0VSte6r7BxYe7ZZznSUh
XClHIz/rQYxZpRDS1fROgz2kiRhKxi0liNZLQ2lZem/bHGn0ZlS0NNOkih2ME+yo
2KFZP6jqD59+btdUvRtCrh8qaSEo+ER7BnNO5qmISV1tCqS9/Q5xccVOEXZ4msEW
nQsZlnLHtnfFG5hWK0JVA+opu+EV3VvBceu1/y45AhfFPRhGqpBiw0MFHXM3YORd
M+XTgdoSYUU6FpT7FJpsIt57lVfKaqFqLCRmQi5yvJgouIKtRgDUpTtEGC1dWAQN
72sxQyyEbGh59XG0l+mrMFnMfrTkSzchDaxZ8WgRsoBKXLZJ8zJzmuuvcgsxxgBA
UWfcATqQ1hXXUFBzu94RIDj1zdnl9ABPQjNpWquuhFSGawNic3ntpcCejPSSJ9Pf
ngLOO8uIxO73nCh3Le961aj79VQqLe0IQYeJ/0ToLODIOpAT+E7IpdDyNb8Y8ZIY
TrxX7jxcGkFWth2MC/yVJxkdayqi5CZ4QuzDMpWIQgy1zJOBF4/+YxKvq96C7LP1
AVmlsESWAjLtyhiTpFhUXfwKFwmzSWT26rPymiecpOYZ7RTmzCDeoafgjCoYG/7Y
hTLv3Tk/ApC12ILvwPRLz44NOOMAbD0IL4GZ2XYjpP9Z96JpNktbOsO9IqTYEuWS
Bf5TTWpQidKkht+cxBhKNe8Tsfy0B7rCZDs8/6hpzdwsi3A69AcajSz4Ox/M7wdQ
wlRPPeo1uyPLaPfalkT7dbXZZtNscJi4wcRLzIkv5dwSe71iDSZnUIgeF8K4LfN1
X5oEn47J6lesTIGnUHEHDh9FtDOIY+/sVOr/BYo3WnT763Ss87i9aD9Qlt6HeasC
0Nd9Kv6sqPoMfLx8GV/sz/ic2pvjCt6wQUG9w4YryWISHVXbn0DENK9pYx0csvGw
J73CTu1ZgHToRwl7XeAKgELTTGPJERWJIduDfmDWAIzpbK0IOH3rViPDhA2zNSlm
rMuqjq0RJcGVbTUBXCeFQgArJMBt0tyUmVrLBgZSBK2fGXlSwPkubaeGQPJa6hHX
Xd9joDA0gVa2Hz6eWOP76UybkOQXI67JhYiOo0tYwg1wz9B8MBTAF7icHvKI7f2d
8+ydSvaGIethmDIxSQbMvWqWLvqZRs4FUdhgXhUKH22DfM9D+R/ov00wpiMjTiD7
bE2PjftlaVL7ZYV5q5cAqgmdfpLFZ4MZDZuA2rw2w2XRoMCQig8xZjBzYcNxQH8C
4ZcMgON7HHMLeASzIXNr7pfviB8Z2+pkBvrNHWzGWZ1W/v50BmU1TDUB/Nu+YZ8s
yVtsj6WjVV4InZUYsMRzEJMPn3o4nwt7WXrbzq3g96Fh+rbB818R0JnICbAtEdFK
8zR/uek8EjSdthBKm9DGYjY58J+52CrrUcYjlmYYhr7xWvIFolfIo9m4TjwkNRLx
kyMfGUdue383YbkKIFWUYPkE4GH120+O9aQvUJe3tKmLAZGAJir8wwFi4FnoJjGB
K+sUO5BNNgrvnKyqEFyxm7wp4F/RCYGcdqLyKvdNBNpXwcMHDfPCJfLTTPxeINcx
pU0VMHGW7C27gXXbMhcunqIr3QnDbXn8y8hiCoJOLKqp3EiSmh6P6v1lcQl3/ZJ+
KB/j7GaiKJjnxfRry6npOBTWgILYdyrwVFihUUWL/sutsVE3Ac7sSRLahE8N31A/
US8Gkj2/r3I+zQ/QMV5kkt70OMdXZPSkEAP5q8YqcAwwAwuumyS0TWG9+jmvAM+F
EM9zVNfH/OEGt71u7LYvnKNdHxAiHz0JcXvax5uDQiCqrHPWmRHwRk6w91en3lGy
9ZE8MwF0vbQrLSk3i7qnoeIMS83bO9OUA7yRXqUw0jUG5HFQjQSGrOA347ybbaz7
coAy1Y+mi1HxlbvJhX5BWSXVWZZQiI+t4bHgRT6xRm1T7/HZh9QtNEcQ8OxUk7Cr
FYdi988IJbI7V/CAwebnsvlKyWn5kwvAdersF3+ioMkVHydGr/yfG5bDHPAgTCHE
U9r/MDBvcmv6Z7ccXb1oZCahhFELffb6O9E51LLcUR7/T1UZ0Gt0Nyx6eOpOV1M/
z09tq172RM+D3aa8bQEAnVPvc0BJ5aMRuSX1xrXBfVnIIFxat49U73B9fg65VJdF
rA2b2hyqvSq1WIxSRdlSCPdqem2HzQdHxxCoUp2J4CTc8cDHD+LXQI6EKxbQyZ9N
7sG1pE1fgXPqPlJ+uJMMCm4YrN9EbIjREcSfJORxf/pbInKJ0oMVUdQ1IHMrm1Ub
MqGajvGHKeGqxR0MFwL6VzAiVtbiqDirRiLb+/Q1a+hKLKB1QT7rM7dn7QT5qP2X
HXrEF7p4cPDdrduuSUjk+u3hQuGJ62S5Z3vtVCxYVKL3NDCWbJ2+8DBD25tKqnDG
bM7SukhLFrO4kkBrJXPRj8Hp3vxeuKNW8FQO11DPxV6sDOsMAE2DLMbq3rQYs9sw
/l52I7x6kZAIiHEIfZSLDVRrjynap1tP/+MBUuhNvpA7sB+4YvPoFW+96dHgF8ES
mYR4TIcA9kkWjJq6PPmZrPILW8xukiSypYaTdljnFqd2DhIBeffmOo7OI4mw1OO7
yvZXYEz9EthaE734XGth2ilMLjTMm2sU7/3qEI+s3ZB8oLc44TJXBpmlxcCXA8+k
DzvjzWlhT0IvaWqLoRVUdGQT9KMKC07z0DpQgK65NscZ2yhJEQ9RxbXRR8XKjDmg
8o5kDwja1HLtaNpUhm98NbsUrNb3glS1ZM/HXGsD6mlsqAZs9eETYZIa8eMBufCG
cJzW4OZqhF/cfp5pT5y1riTra7A0SFLeqmO7+hXb5yJOr/sNo+A35OpeieHgXpOD
GZwPY9F0yLCm8YfJAVA7uDTPVtfbsBU1l6KJZiiu6y98glI6qSB49e07HM/tlHzi
+GCqZkQeKEUVtfOMHmE57p6SNoVjNuNApmDy89aDsWsYMkZdVHfrXtEYLdxakouA
sWlVk2ceK5J/N7jl8DdOa+refg8KNYkS7Bp2maFltgEZ/hbTnPfZWlrYGfp+1d19
HlYDta7KKI7AfJPP3DtQY5n0TgAcMUUQovvACAvXD/j9BiHh/aoDQ8zhBe5vofzn
5XtUTWFtVLbMwjTtre0kIroDp+gplkkOhQ1Mzoh44ncPg7YdSwqlTMPt8kNC62Z2
lt+sfy4Ru5tQHtSNnrxhwriYA4rLsho4/uad/eUJlSMLJvpiNROGlmtGwHz8RLG3
wQyMOKW13ELMUA9wH/qCLtzTFwEz4f4cWWiA/y9uAzI/vLfIJHdVXTqfuamhXxJh
Bil6P+BPeCidgITxByOQ5EVQv0he+yUG49oC/Za86N9NWMWkLh3Tfi+4c3lYoJCF
rNl6f0vd1Up0BKfdbI46xZRo3Y2OPqKXCSgIrdMDCkYTrjSl+gpobBh5rOqyoNaS
NKBIFvsZ6h320fBjtm+OupfMF8G0axrUT/TrBeNb58tbmnqM74oASQNCqWd00xbR
jzd5B+IzXi1OsANrrBSYJ33R84hOiIVyLsv8O27/Zz4pgV5XXyO7BCSxrPF8w5BR
XuzlIsXHp8ofpGy9F+9BnQeZer31v431ejYyvqZ58zrP5M4wswzpdNONCppdb20w
fC3V7P5FQArCFNuacTucDt2FD0MGHN/4H0VENAjxpCeBB03BwnV5d5NcUUK9simR
ljXfze2kZGg/PPPaJerd7+AmukLwSUkF/C5eSDnxfrXT8gQ1ji1eaGMwRYh5IQAB
MIFzhXrQtYlEm3tIFIxBkvbk6EC1zn8BWS2qUDW2IoIu1Tmt1NcKEjAgYzKUBrmP
AEJohdbuyDAGFega3OfKC5SmZeXGF0k1umF+FjPRcp+Ci0NSeH0txZh+mN76pXmJ
VQR1Inq/aGBgSYGwbY6yUGv7hxq5ExsPODsXn64W7SjhdZCT+JXGxBzu7xZ0SSKF
rz+hsWr/HNT7h7K94SD4eyfEyKGI5wPiPC4nxxhp//zzL+CJ2mcRtbwc4oIB1Ay7
TWWS+9OwRzM3jFXJjMbZrNybMKnwjFvDUxwICT7dhoHcsXxa1bY4DhhfBG4Su6qK
qXDTuI0itoZ5rNRpt3dU5NwPjzIt2Jc8ybA0Zm1BW9o+AvvuZJtBaoxDlBJ9GAuV
6LDoQJGdkoOBuEkfr/LqqCa4kFc8WreUwBP9YKaKtHEa7UZB7goFVbICdYWHcaqN
4mat/0IL7FFpD5eI8B1gwEu2nUHesSMqAl+HybYEhuZcpH6pdc+au04TX69ohTpD
Ui7EMw+C6uCxgE4RXbonu+ju6PPci1b1uNezaQszs0apikK8wGvxrLItpifRocvT
96soeUfW+NQDQASYjtTxQqfTcooROF/Pr9g4ex9VLEdVuAZW3tNbxdHuYwBja4di
m67M9x6edgqtVpWalELKW5OiXOwloaZC2bywfryYc8+t7yGUvTTteD4xxDPqHQiA
vLSn7v84HxfZrfMQbPFVmuDnh3et/Dp6jIvnErhlFQ6/PDVhYLzf9eXrYVu/4BLu
oXjlHKPydU9J0lLlonPlUQ3th0rktdGFd6PlGVM23PKg0c+kFAA7Rjz4MhFRgn9O
n9Vr2BkymZq2xRb/xEv/1F+eWSPqkM98nVVQ9QSQ01zkrAb9JdLOw+a4ZdVrIqUp
R4wZ8Pre3FuFjM4qd+yYLVG6S2x0V7z3F6LzLL3zauIRXwgrjBpiZvBGtvUKyhn8
nBaJnZMaC4Ke16FEL/QrtNLvExZHA5SiigWfy48Q1gNfhSM+c/Ejei6BKQ5k2eHs
eHT2p6i5PEaeMPCYEKx9FpmqFynsDMf0T+dCAyIFqy7K8Z+4m/6gNFTkV5M7A4el
dejyC9OeL/lbTkgIkVFEWGeDX+4wKEYLDbTo16eCFurG7WpDoOfyidoHoZZl1OCY
xUKlJf1IZNQnBH7aBR/nSWSjo3/r6E6xYe+OZMNIiBntYnyM0lHzBZ1GsHbHRJ4n
IshusqV35zy1Wt/hQ1nfV/zVMaA9MsQ+j7t0bf8flsLmM8a38M8i795kxk5h5ksy
ghPXb9Qb6EahwLwxoV3kz7wRB1CW9hRdccUNYVW7hM0bOg8WHWaRZ/UsAAUkfzZX
CTzJo+Xy8BWPUgumG8dQbvvIxjIllvF3sIH76j61BvYvB+UI/g0CU/rssl13sZ+l
CUyy21N9yyjEfRmIL5pUuMdJif5MQ6PbdscJGu1rWivWVOgKZLrtj8qLm0YYkZMT
DImhPWuyWWxuoYO/Fd+Kpzcp+cDY1btSq8CVQ1ZvzXnqQNPue5hekAm+jomJ32FL
11Iyg2WUoPOFCSEIM7fmS5weaGysBnXCBgAdSGOCbPknWB4Qj4gaiCBszUMksRAL
zfvY9js8+UUFAA14hL01WsCmdlB5x1LCXZ6jFk3uD4RWQR2h86nQNI4rTjovilPr
sTU8QEmmsMiskxYEH7DV67TyzBC+JYSIXfPvst6HVPPEJsoO68iiQJl58laKq1ad
NF+nSqGppbS7rHj8msiQyIdmH1H05Iitd0RUdKEc3JBUKxbN2LWSMDQMyuV1mrsc
sXH0Tjiw3BgOUgE3v+91TABS0XlMS2JJPvBnEZO3Fb3Qb7QKOf703N5e+x5guIDL
82Nk6a6vFvFSrSR8glj1n8zu/6c6C0HwCXWh3IrRcOMqF+DBtEr5zr/b/sJnGSdh
aOGnXbwn6GTdwY0LlAo/5MNEA6lQR4ITPoh8xXaO8Jm7Gh04qbb0cw2ZnWsQTuKK
CCIvWid3ddArsYR/wrduu8wqvHVtQz3Q7j+7QMjsIwF2mSIx+yF6Esy8mWnLCExz
ZIHSvRYGaajNxmxFtdY5DGsJxOhjErsStsaMj/So47YWDVcpwNhsqGsRLArvej5H
898S6RaGq7DqWI/vUb+WOSERkDaNnrpwn1fwCheRcxVHbme4LFS0nJ6KPu5x10Hg
uvD6X7NDGFlS5hF0PPV6j4iZ7YNftdlX8yN7q9O1BVgKxY8Hm8PrdPTwKY3STD25
guth036x5OheUxgTuZcFRXXwbS5IVK/CC8fbMR98lQQbZ7rKuUN2eL6Y/zhK83Wl
s9cI6Zo0idbOqlMajHNQ1AAupFbkSXJz1vhTaU3dAQIDKFUBhK/MnN1+FHUv8pyo
od9MIQTQzcamHbo90+daRlYxemu1ZPpgz8uO+HjtMP+6dUyA5UoGYMZfT+RTIRaa
aDawzsjdchNIP7RIxcvkRUJd9fod1lkooClD7Do9Kdky5kuq1vLL2x77qbyaYRm7
D0chpIn6xcTp0NNorcLC+u4vcAgGExHbakUcHXLzsMWnji09IoSdYi0JMN2tQ8hw
DrGghBxbU9bHfoNLyKA7eX4oiygrLe70kN7i4V/Ft2cVB2TweCuyJgOZM7BAwbYI
4dGMlNu83pJcQRH7Bf20tV05c0cZKym95pcVNjEg8/ETjuUk09mQ0rex8d+jeFUW
xTCJfTcqWWyjGIhjnvw13G7zpJh9ffmUj//n/We/4VcesKdva4WKp5nd2NJyGe6c
3Fq8/VpvWckT9L/JZztuA5SuEatAFsqOUh1k6FuAd7iJsQdbVlBAGoqEWzdvQmqD
Fj0WyUWNdcGoQVvulYbhVhrimEN7dKTDSXLxUAKN8h9zGYgKNor3HGDsYfHnTPlS
JpPvZFGPV3N5ArFrgrlfibyNDeHJsnCNioWs1XiCEZ9AwduOCxMA31OHMpbhfsH/
j9LDHPWjRsvKPvQ/go4DzG1otqNkrxGO8dZXgIiW1XOcRAb8p10BxZyTzrxq0VlO
veK1HZ9XzjoJXIlwlx7LXDGU3BrJcYvKjivny0b7aWaR7AbZuW1wdU74tm/OMWcU
xDrons4SBUnUZiQC9pVFW8HFC3O1vYhUx/HV7Sw1fLaW9yZpw1XCGgH4Z8o/JF/N
6po/1VdM9ozHeCdV4WXEv9A2am4Ae8TeVyBXIv+pjpM8bhrPaqozcPjDwNWowp+x
YbLM6ddxX+M2djzlepqxNz9klFlywgrBDPM7UGp8uyH6S62rvMf4ydJ3SJTozEZt
DE1wCp705aoLDJqiVjFzySH7MuIA8XG3+s5czRZqIKy5SxbXJsRfw7RMoMGsm0sk
ZRGdQKQyVoWHcfmNcGYUDE1O88C6BIFSojUJG9alj3jPLgJZyY0aGPwYeQh8CiAG
pzJN4zPwb7xv07s3Ynk28G7/3GXcizPCYQ5pykRKOIkEiI/h+XxCgY8fGOH9OK6F
bRddVJlCGUI3kK2yI9oGJuOpVKfA9nQxYf1XPDPc6+Bpu1SQfUw4b+OcqQDjh0pk
1alN4KwzgRYnVjQFzymuyjwQdzL46OLlwSLRhxibXRDQZP0kiAmf3dadStADIutR
EiuV4EhXzoeHz0SocekbjbCYyH820eUJFaaQlB2dUF6/kE9pNGQ6hxJZAjlUnBXt
1OZVwXWX5wWskh4WHFzdCX1eMXEGRYreohWVX85NPiI9/T1yOnscUad00yteR5Mo
Kp0Nn7iRtOXKCEpAFcnL7/M8OEuwocHdaESwTVKJv0xzCfdZsp4IOu5R33AZs2Is
uiXgTp5Oo0RFv4JCtwXrm/oo2cECG5vjy3tuBJ1JjfZtktCYe6Tz9n+fxLJeGWOu
DJA1ces9E8wAEjcEai3HUdJvvdPl7fkdKxj2b0XGVhnqRBooeEsVRQ2MJHJsBh8O
C5Z2bJIXi1u+o/zKfoGbZtRRyKkT3P2mq36lFftzcNC+JwAyzO2WbCf3j1V5Ex5g
MNxhT6dGhaFbkaOSgktkzF47LJJqFoi8BK5wIPnAjOZ4c6qDgf901z8LTFIvvbCO
2fgrODVYgyfDvx2wGMNbDC7/Pr+bhObtCxIydonhDUEbRkVvxBZLR8LAU8i5xMFg
US30RFlUK/O5S0ADgM3we+wM2zHL0yNVi8taNvDn+nSOE5+DB4EjaEOkWdjkc1Vv
po+dUBVHXPEsYytd/22hEe/lUMGg3bwM8yXUyo6Jm2KTtjPYUYWzxrNNu2v2vJrp
yQVQLpVn4GUIXJ7SQX14ix91Tl+1/RoH2eA6Iil5e6Wk1KXgqOykQyKZOIBp8yHr
rXyoQOMmJKAjOCUj1e+nbKDlUkRyGz6mB8MN2zAbAKgCkRPMTpNxJ3aLsm5kaB6E
GH3jwtKH0jQzeITDmJ8SM8oNEGw+VIFlmr6ZdJKklKwUEASByGvPIhTHya0oDi/h
pAWEyMtggjfnPZ7Dss5dc023XTvf73a9cHBA8SWZJAoD0yTTzv7CDTHVTMt6Qt0+
YyLtSw/ZDaaNHyMV5DgIgMmyv0HG0Mp2Dnl7rkEagT+iitcz19LpUoYzFDusSpsZ
dbhtud/mXURBG75FKI0MMWQmpIwpE5j//K7c1icXRLOI9hzwRp0mYsm8eprwh3nJ
vFznziTFdITD2Lzhu1MkDqCjrvaVLpkdpSwzNmzbdvMX2ywT15habXQXOBxz3P8L
ApOFTFqW81Qmb/sstdpbTZ3rQfAQKElQHsJer8FffErsFhW0OvWPmfsaUXS+OJX+
ObQ6qU5mgK9QUdneJFcsqXs8zNKWLCnx7G8ER3tvWtLW8i8PAhINdhVtYK8+3iu/
DtWhjjdDtlzvA8ms+/H2sKPTWWEB2O3o7YripUOUIIK12CbFbHNjpPX34D5gIesH
Q3Tm9FDpgI9Aw/+IUpKDKDro78dAv1Tp+eezyYY3N96EsMSbk5ON5LxvJhMwA5jg
YTMqvjLLD335TuVpwhgiR9GYKVIa14BOEwsYoBupizVhcVtgcInmTox30qzVcIdR
k+hE899pE9wndvSaaYvO1o8EamNTFgso46k7rvMbeEXETffi5Ka13hIxyauIBjF1
xeaBNQrY6xdb4Zp2pwDQ16PSo62mVkT3XDDXfvFPJb4KCnRTYJmNp+364gllhTLZ
i6HMqbYTYk0qMWFGYBOQEBkVrJBUcCAGIAfEyFZvL3//EF8kPD+EoARMVJmJYo8Z
rksv9n+elTj6TY2uZW5Yf+VkpbeaybvWSy8O7FJ9vRZj1T6BG+lnD+XHWT36jOxf
vma/BRCW63PILkcfAZbxjtD00mMnhVRH52yJx2mZMpEI3mWWfAle52jQvxAykAr7
g8Q2nDclcDR5DgFiPTTyyJGic2qtdlIsvKMwu0y6rLX1ngVeh5Bs4aH7XUHxSyH+
yxiEP39NyoSTIC/uMcdtFPrkaBe6dqPyrw/+ZAb+330FczwUfTEwkjrN0JO5hHQH
CvjhTj0dCltfEM0e8f99xVf+b56BLkpQ8kbHCExW0WLGbRgdyKz8m8koB76grcLV
IDzRLUXA17QQAe59AhrwWD66H2rCtLvWS9HTgJFWsC56hon06DjPBxMxN4vOGo5F
aL5E0WTa3UIzUtRh0OEJ19bVuH0aaUyqmeYvMCpxVwFCVpIuDTe6fJ9ydsSxanUx
rgzArAs8ARyWYRKxEVWiUK2h+s65QHdSgslq5Zk+A1fKBJoJ5C+Ev5S6BQe+XzBA
wbRtgfbEnBH5sifVFE4tY1pEA7YRGMtKZMnixw/32blbeJOtLPDHWRRGsvr8jIe2
yGKA+zoM2HYEBnqtdXbKxaGzFtPwCIvc6LdJxBvW3f9BnKFnyJRpulZRWkFvzoGJ
Mfn3t1BskhKQZdzYvakixTa+rqqFF2odbi7f/YZe4sTOJ6/F7iS+7NUkLmBnhWAs
8UAUqPON7rY+VvCTP2n083xOtLCfZQbAvXY7fnzsmpAcbBK2K3HKeV/cBIBwU+Py
YZsnRmjjvEoNVaz+2402oOSP4DR6PwcRz4rTPvycRRYu26Zu3zu8LZbtTeC5IE6j
ftaHJ4ODTvJMvq9X7xaBFWVSLCQrPhyGx/b36LRSP6AS5msqFczxnsGO1nX12kSI
OuE4NBuEU8TT0e1u7GjyKgELZK7Lq/CHTFo4tMdFrFRDDbT8YwmZuA+OFJwVUgX/
ZdY9S+Fh26ftz8milfhH+nTT/pEvGKGDGmtbqfusDrILa1BuTegAvtKiVu56a5gH
IDjLa4xe3O/dreOXdUew2QGTYtGwzjcbldbrt2BgBKxKsglRgeeuzs4a/rxK/aOU
Amr0qkioTzSfjOnQMUG7FUT+hzYTAsKigwlx4CiVdfzhuH6wUYy/LdpVE8OCr81o
gWzdgSCCrWIsHX4tf4N7VDiobvdqAmUuNFg4DDk+vfIE4ny2ulQrxKvJHCg8Qv7O
c3ewNd4JmKn0D+pbhO/cXMrB8vxmRBnWJvqVJrZ5i5aa32Y/IMaW9LKzzBcqdtcl
SQzo+XMPzMu8XbI/xI5/YdXRb94gTi6w5q8vBDkiM1ZacQKEen88b9SiLI7mLIwc
MX017GimxS9ZVLvRJP0PUuSn2JaSh8HxGsJbIoHraL94UDiiXAQUUCYFL0hdjy2f
zfW5TdtI44aE+wNJaCarrXsM5RmULX6miVLbEm18WczluqUdyrQ7msurliHsGVJV
C085z4lA298pkGNl1SKTOwxGpJmGRPNBMPQErxHcdYvGPN80s6y9cKEOjtf/zwWq
skC+H8jKrdFDsEE/xLx9DClhQVR9LFsBfyOJbe7XmGnDOJcCv3DhlAI9NybZMvik
NIztthkms5EPHytoa7Y4Kfgd8qMqbc4aDxisie2ZDE+iImnTzj7b0iFMkMujVauw
V/mqVChh7b3hX+7KT9wXTAuJMgvJSHsRte+QfknXHr5IK3a0rT3/xMz1FMDlOGcx
hvdqJXidiNnMX8z0QzoC9PXnyK3uIk/7HrvG8y97UfsUJWjjtmmNsiVHvHFs3ao8
ixpkPwfJLJkrQ1YAAIRPP/Nfa8PvFc1+ej+8tf9n6QF0wAn0wuCbdst3VUDKrMF6
vh97oudzIn/0TP38UTOj98eZtaw+J+C6Eo0XPyQrjplHlZLov1gdvHpUbDt/69VE
KSZNOmjwXT/B/wZh3eGPo65pSzadt7NDrFD1mM5kGw6htXKE407CZ3Ro2ruzRvQH
BdrAF427ghZk16aLB+nigy08/WmT71ALEKjqJy0PgH4J5md/WutdtYWlMZdOgi0p
o5005UFkGvssZCWKg13GDYSObtbISOIFJa2fHySkGzIzr+Sof9OIXgiMVt2x+LsV
GnFnwPB+HvLr3SRo4UboeNRYNIrYkwBrEzIPgSxwyCiEhRJHosxEBtBezBELg+3Z
SoR4FpEoABpdRHVf+sXMyF3CmPwRqD0UaNePuteVjbIhlu6/uQDbZyXiNbDSxYnO
sol/rPBITwTXRAdUVP+SFqW9XwjIjFYwz8RN7T3LeIhuCjbNzRfOHbzw7zg75wNh
8wonFzUq+T9sIB0WgxCYgW2uHpr2pZFHENCn3UYTa3KmhlyIR0E2kiiLk1TdkNrD
21Q+k4qNPJ0uW34f4qdp+L3fyemxUek0KidsRJDYbv3AykbUSzgTWnkVrnuT4BSr
EWSn4YnrCGdiW3r+BkIkvcKXR5a1X9Q+5BD2r6m3uG5dkf2gHZ19y6L1YiG5RXs4
ArhuS1qJpRx5gK5FjtumRw7q8dJaSr6cKlLtWsA9EWQCS5wlggprbwwaN8dkp3N8
8C86TW3RJm9XIFx2i/uOCze7vMjX+JFbx4Gzjz8Nh9LsViR4K94sF/Rntcy8wlaQ
WMOYsJYPWrx7QMygSHqiBTeGPCUOcAnmf+hvAi6NR/CG5FOtu1ZkdgY5WQseeUmR
vDDtd80qa7nVD4MtnoUOaCnl/XQNqUo7+02RIsVnAXHGe2OzafYsGMVDDQhaaZLO
geBxot1mOShGxuHwnATdi/oJqvVQ4DMKVmYZGjg5EdIKzTDLag5EWft6Tf6IA1i2
wH6NDyJkwteQobgyn7KozdQ8V365kPmmbY3nMBY+u3t6SL5/SuVjZZVOD2ednd4G
BSX8QTXEgLzMEcUcRFmwsk8n8fOGcWZq459IE0OZ236J5rAydVH1D1728VjvX4xs
XLop+eXkWkNTPV+wgX+QrAUVWlcXFX8ClHCSKdQKxD6aF09cQIlHi0+xUfu0j7Pp
BJfbzKe7NuTnF/ZLNG34Om7zW6ngiuo6MTzSJE2vhhsCUNrxfYdSTrNVsC726XZV
rArdjg1QEczoddk4vTT7tH7k7XPw5ey3LMPUiaWIZn0L6C0t+KFKaNnyXK1XRrVM
xct5+IkBkK3EVeyyIrqp29DJ1d1OIvCT/hZKGO/9Qf1NqIHEESR7YrpIl71GFihR
NQ6jaBG7fzFVjZXRiULUDrlXUeyy+cw5OWg1jLIsE6y1CzDYEbh4DYpO6JQDeU/5
71zqDjF9ZhGZ5v7VYapV3Um79pP9i303jjbQOXo6wMr/0mr8T1f4kUzXO7Y3TdTo
q9/LLzWgx37xG+fsr5e/RaEmxz7vOAzT3lypC0NPpopz8/T9bctlvMBKt03bunB0
M7KtvgHGIBRY0SWRFjSG09vh2CiFyv8WPHnAS6HImrDrSg2y3sN4yjFkYRCXrhlb
XB2th2WjfVRTkbMAOHESnbC594dHa5+jaAERw2sElV0DVoxypmbEsVRotKpgbAoQ
ht/Ywsb5hra6ZiqL+Y+QOdu+01muhzcmpfrSqebqON2FClXqbjKNOJ2pMR/BpHCo
RCTn/ovgkZLdxGq0eD69NEtFUqPleW2WweriI2zWp3xxInFhxRb74wurDo8w8hqI
6z9l0aTCdbY9pp9xG7TcASAgKK7V42qKSxXSb28Z8hQflpy1uBYAluxkOphCNH1R
PyQECYtWzKyzHc8LFpnXZwNndoceqXqlgMi3435MWuiSKAenFjWhLzDHUJ/u3hHR
KNZHO3Rd8SZfZ7bquBwnjuZASHrZFMNq/rwa0EOG5MJcwX4gadvoe0r84qMlY/ho
wQhwKDGlwvozI8v49X8DaILgDJVZ7gFh9js3k7DpPXXaYQteMKpDCagEHsieNfEr
QLmb0NdSwv5eK/JANV2GJeS9NKbZp6P27veIdTNbM64pdYDiA2xtmyEZOl5K7+9E
WlcRYK2ZPm9wz5t5Ql6r0jD6I5HD6uPM6UuPjf9fh5dBcjWAOG4yVmaHPwXArW0e
E7r/S3ry56x90Tk+yHkPAvYElBLHknOoBos7G/E87nZDtd10TqdTt2lsOPA9Ppjn
QoGo79UPOXBL+At8HCzSxwht2lzZJykeGvqbuS4Uk42AbuTSdF7Kvi7d9bV4adt4
vLipeqKt9l5ttHIs40iYOmDD0e2YYFPBScnw64I3JeTRl/kTmIsoLirY4KWe0dxt
Gnj5087Pf+DJlaGUn92xvUMUagL2FP6pzHbXe58wu2Fx5lJYcPZU9ei0qgwQ+GWR
tABRwS90PgxyXfDXyRDKQtn4hq9bH++/GSC7zWv5KbqLzpcWvdgrwSfM8mztouKV
AG+1QwXgyDBQVyjQzPtPtGTENReVTXQInyF4VLEBFCOwzl5iS+r97+8mP78GjdFm
Va9ufBRJPjOP7PLpwo+B0f0bls8nI1nCRkx+0/o3A6WhqrgeBPkMYz+tab9GTvMJ
izkgdD49DJ8NOxwsbXDuHUYCeB6ylJ6bREjIbd8z3+redQrZ/ETOmwd0qik10y6y
rmYT3OQbap3gun1ASvwQ1FuPiI6bd3zm3GC3yvWkwJC7EylhDrED1LGWDIMkv+1V
smPsb7KShUDofq2LqYNpe+0sZkZjB3Wp6/oe4lgmZpDzPy1OnRy+rYv3bF0JNRyx
Kb61D2WbEm7f+A0EFoBFJnlmb6VTtyXYverv1/7Jmt2mp1Ic3jZam/LKHixGi02q
aFpLMMv8eLP7eU5uyXda7om3C9pmjmNl1NL1OOt3cUkthzCbioErS19ouy3y1Gyl
maMCanNsd3QPLsSUhZGxDkk8bZv3ZfMPv6tDjF52mRs41SDpCkD/i2iw1sKiklvL
81D19p3SPaAhFJLSJyXWqR5h8W2evX3r+BmTh66hho0sBmQsW1ei2LtAzsbDcuEV
H3LoGZhg7+BhXl8GQlvAlVUlMRT5Ir8ibEngAe3dfzerCURwrJMbPTB3Zru0BtMa
dzFe7tCPtnTIJ0KxLqB+dZBY5+cPIyLO90EbGz4kNwJTKd7xSl2sKM+Pa6FNHoLO
l2BThHq7onfin9jBrhjoUWsGJXcZqHtBpdSwRhXkQXAvlZ+bxeGyAKzpoDX7HS9D
/Iv6As4E+VS5yYhrRDbjV+778fDUuFKofQIDtv5an/clRujtiY+ZLyuul9gWAzER
dTiaRJVnSuZkpyTiBM7z6E6gD+bsZJgNKYwqjvlcXINz7PqzZFdhWEOIgXZuLUUr
laS2uNaG/IgdryHKYcQWxOcSGufgw6gsIgyxcG5jh0mUGwJjLMM5SA8m6QIa0Wxc
l4MKeOwRQ+AAxb6q7YTXZxUh+R21ISiDQ1z3fW9zzJE8bgTWrI3+jbYgPtU55ljL
CfEx/vrcNeibbbieqzCJ9nXovf1P3le09B4JxzgTwhBvdWr0DRlga7DXrraSZrRk
XfN3cSMRHmX97drYltkUhlA2jo5rrVEuyBM9Sbjm6jQS63ECpNO6DPk6MydkP/JS
6eT1Qd5lj2OyYzEa2u+gkDOowpE7vv0XpeVbXmAHu27kNLz2hd06XHFz8Vc9wg8f
3nS9WDl5V7yFSXGkGnmXA2M52iv5F2MCeP3oRgqDPsxQtvMeDnLdKP4rdcgIchER
SlkZ3nmqAYyuytK2PgMt3x6yUZhFLqCj/7FiXFgY8oDE2hG0mbAwLsLPSqYbvFdb
7+YUmyQCyxeHfr/MEv9pURKa2pcu21naP3Ro1yyTYitvpCE377Z6C7muZm5MY3Ce
MqHtGSXD/a/FqKsr8sF6NZymEnKhrcFrqgWX4EYYg4I8czhTOaW0ELxOTRyYz1nY
d92Il7rSXu7Rup5nPi4lqnXpUCERpbAUpFFDrQtpEwme3VHlQe98cZlXlSq9TrFE
y7Sx1MvbtZOVZwKHQ0T5r4E8+2TLG7RvNZEhb+h9w1xWIslCL0wWBRFxTeTi0w2R
BoNmvLt+E5UQmmt4/NpfsHUaDLOjFWTKDMj5zHcnC8CsHawU2EEoCSVELnaafJuA
mL30cVk3obAvIg7Tm+KeutdvASFKacrq7rypbZFQXeoIhZ9zZdi63x5pTifSwCc4
yLg8Q84bGufYGzfOAyrRwJKa5rlEP92kHNuHaFbNAOrcs1Uc8VKg+S3VnVMDVI9s
eFAd5H9DGzEJICWqyEl5fdCY6QBu1dBBDs1uZYDGHj5KSW9+tFQhP1BAn8z0E6CY
zph6MPsVYTmk3Xne65JXlMufb30a7VuPfacI17hIqH9N8X4iDIW68V+wvMfS/QqA
Latsi2hTqFkfERHqS9fNhpYkRNLAC1hjKv0Hd0x8XieK9BmSXYXNLhlmTsvNY7TW
Gq5b0/MPmTenbKaHDx67yrYqTfQg7zJCs182jGHLH427tB7gxN7OhC2/gj5YvQYJ
QUC60o/rfOoObGEJPp08XIrA6LQZ6LgSbuuWkoyNTY4DG7qqbF2UGZ6sg8d74NlA
hIgGsaIbOA2WTRkSGLI376Nam2bYGNHFFdZB+7CmH5xjyeme2Thz+3ZbdYhHEfsD
4DiBApsWOgp0Mo2AUWyV16GP7y16LG2MDSfUpMGaCqdrI6tIJE6je3LGiRIXdtWY
+DaZdD5+gK7JTSzZaeGUN1ok39qefGZjW6TLunS4MRPKKcUr2esKeyvvlrJJxlWg
4TGL9MDTY8fz3VbcHthlYMaPylUjGF4lIxIotw38C/v/Fi+Q0qps5xFYiSgUkVnk
EA3ty7FXxxJzVCHOzfOHMvH7jyeBXCvAZX6j3uugxiASk0HEjIhXSbVPZV5mVUM9
Obts9hKe52qotRHplb0Lh/Ejw2byHXwR8ZYu2pPYDijcEIB11sbfyyDb+kbBsgdq
v/D7GSt6D0cYG//ulbOTrp3ZohyWpVNb5Y7YZi2EhrlgCFAtcCWUfPC5v9WT43qA
Ov+r66F7PtayTz/v+GsGttwwLGt8mT/U3L7jpM4pH3AIaaB4Lyq0PmQm2QOBJhis
etmO8zlwZrtwrTHSEymjJTBJV2P98ZCndchpkbY4+lkJNIY3RyC8CbdSfJafS3ie
csK2vvxWoEJ++VE4IRSFma04q+OiqdsBXFtf/GBcuKJI5NJV4Hl8DAMsZMMINF3h
lYiP8zV5kTbcQsOeMvQHvUqhl+yG/VWe+TKUb4C+OoGvNi1Y7t1sb+ep5dQJa8jm
RMyxQFcSq5konoVTP7J80luvHMFwO6Dkx7kyNRQgwT3MSILvNW7hFffw4jAGxg1U
tmQf8kmA6QKJQ47lbcqGk6uTNIFHvluC7Bdb+/WXa5yODizW34cHDPr0hx7ekuwp
8QY+h8kWjfeSG048vEf6+F8kqQQDZ2CAjKjxVH+bAd/YaAuZ720gNPOGbRoYECOJ
2K4xx2EXBBSmbp2J/aka3Rs4F+4wVWs3TlBO2NXkOBAjazEfRcSV0DXsG39t86ik
DfXrsMuk3PMOh0ft8hyue2qrsju+zS8NH/ZZJmAMvt8QClwvd2vOfjfKfQTILDg4
5f1OhUcHolfYJKTpz2X9jhh0kk/bT/KVMeOCyn2awyIUv8ykpMTXeyWbsdPw42Eq
5plmqMm9aCCl0DPrHdLCw+ej7llvkWQcOEhm18CN7uGUGJFKD6QWt3vgHPi1l7hp
YN9RUDzODbZEpjL9dcvT41Ds/h4URVI99rETqVt7pqxQOTO+2rok6ujI5kBuYUes
siQQBEbhgEI4rQUsCDWnyeQwqOEGw8n3FwWIZ04pRVX/q+GIOiOSzPUasUpomrYh
bVDzQ2sbLD6MLwU07v2wm6/WJxFQLTi4ZjR+LE2Y5GA/0nHH5qzD+HE87VdMr72h
hvng7+8T2gnhI/LiHoFYOD3+O5hgrbDd6lLbbeMva4kUrQgnIZJHqMa48PLETXRM
ahkIj6OsatUU3qvDIuHYncUKLsZJMGI+ayPIBpdpep1wYs7/Q4+ZxHcks13RhfaN
fsIrgLYYgHjdbcA82iA3u57E/GsAv59DamD81p7//tFcuOcin5YzU4ttUq9r6q3/
O2H1POQjGgDS436dzMtIcJ+MHcdpK2qLPULelKTW0/si+FqkszSmb1OIZpeL/lXt
If54MPtJLZPoyFwPLkuX5cuJBp4xkw2m7+KOhnwyXORFdktN+uaxBjMUROGfSnHJ
5IkAvR3WyiYeOlNpHkAog+i5xTcjcb988+KeHduku1vow+kRzuXua3o/g24J6Ddk
SnAoxIY6LVu+nlmnGoN4c8zyTfbHIhjoQwumx3nG81bUw8NBaSKrEVMc9q5f+b1w
tdmE72XHxiU7x85lvzWjm1VJvW93yKQUvqB5W8vJczzlQiPpZMdmRJ2U7tkOlBa7
GYyfWSUgAmz7GHPhOCgmVx7zOIOl8KjT+Bnc8hc18TUX01qu1Mjd2UNCQ7XmfYn0
mbRieMToem4G9RH8bL+vEMcDnM+pf0NrGE6eXcr7dV8vJf1ZEGNohbbFh+brRjqp
LEDWsXO33CQ0cl5p8VMWhN7bcKz09u6hS2PP377yHu4iv2oBIr0atxQh35BFnf6/
ZqhPkLVWM1h3if0OtKmPYo+1viUEP7fj0ROKpd+CUjFI/eoxJTJlAvfM7cDtu48z
cD9NMmjbHhuDkdM3qF13CqPGzCX7seCSFaH/AK1Jdpjwckkh2M7p+lY1XUxWcgKu
qFDwhcPQ39Q2cUyR9e0JGMj3A2rOx6pFMxGE7EWMq/FbbsTpwXhkwcIyaVewTaEd
Qe0Cqbqbia+Vj5thMTmuXhMdZqVskY2rpofmlHEfF8iGBcsrlGfIHQf1T7LhPGwG
ZNKKdVgfpgBBlA95gKhsgDDJRgwhhLhfxcywtHzCr8tChYOqp+96hLBQwfDoIWAj
BQwV1T5nxpQh/EbPFHxlNkYYGl1hjLTa1J6pBuv80mTAV61oNaepOtADbeDi+WuI
vO4tWceofc0zuLi3kp5WpgjkLvJoR7fwHwzTTzAqGZgkQctWNV2ZSgMTAWCMKKbb
2blPq1QemSNV7M31QKLnQeDeQCrQT1gvt4RpBXlxga2sVQo+AlGPf8kHPBOEG+wQ
MWW0BrKvhU5+QU5MLdL5Ley38eUGODMpsdl2o6Qt62F9miUxqN8nMnPop+QduFdp
QZ2RBkdOYb4sopG6rABx8sufXtMZta2o8yVXdvbdyc/XkwLCRza96ABurpu+EZZF
MoaV5Bp0I8f6SBQEulMsRlt/AZ4pmiLr3RhiI8G8wAXF+KjlNwjdSL2Jd6BMPwV6
vlAwfX9fiByB7wPYS8bdUVPxZ6mu2lKGpo7nimvvT39QUPUvwkO4HA6E0SgRxerd
IF6WqvAX8O5jL4Rp8AXsrzUGhSb+dfnkCZ8SPoO+7EzCpcaRNLM0TQNtMnzpfP2y
bzwnrs7MCjs2wZamve2iM03MojIJ+VGtIZv6vtNZ+rO2FsEJ9LQxW03P0k/CSOUi
9g88RbHK6BeetCzzsrrYvtrL1qHKHgAhIkMUISuXa87L+wckOuaQHlu1Xbn3zpd+
94lsP39ORfwbP/cbZJbikCs8yJV+4C43o9hC2eir1DOwqez1etF//d81cs1VeVS1
pcur1QKa3EzPK9YT6LwGlgyvIP2dq1NFtISIQI+eIXCIxJGxroB1EtX3dH6ZrhVY
XeOTDpY3JVACHTFRdvZXTR/HzDrXqg1dUirr2xXOR043g2N2RinYBS/kvOkt6HLI
NbvYLFbAFA/rqLImSHQ2ZZ0SAjrv4X+pENvHrKheID7AnZFpPXZ+xjzOPxRtqgss
WR2SccL7n7J+cezuowoGFbdQIj0nX5PCI5NEizC/A2s+GkFD/BaxQKZNCE/VrIt+
xzGv405Rzyym42b1y6bZbrHgdFOPCPMG80bjpauihshomqawWu/Nv6HwqXp286QC
LGG/8VILq3ahefHYDlApNI1XWteIb478VrHx+QmVjCn2g6ClVb7+d2uN4i7SMybP
p3BITDupY0aOf5FZfnMXmlnvL8d4rtYsh1+4mm2+QtIWZBn5Z6xIDP4hYmWZhPNd
PvFPGQRS6ENYk+Lxk/yyb3yVuk9Yq2X9Pf+IP8EAP4pzEKWrRLtsqbssxWiGRiY/
emWfHrnJtC5vgWSLzc06GozH1ur7Vtztz1Xa9HiMbS6/87gKcy3cEAWAKIVjuGP6
DQNl6XrmvxFb3SMBqe3BAhp5ZVkxOD+E0nFX39d+q/SXqBEBtzZnGv0633fIv9dU
JtIi2wZMhs9HegDhOB7PuBOe1I4qHracamn1ZCFCPHxKBrtP03fGrysm650NG6n5
StrlhUCESJULNiZ3daXzFSGRcTO2aVNWWBoLsiznOyTU0SlzPRdHR0o5oN58sN3w
by1eMF1/PdPIcVvz/4ZXEDF/I7aI8vGqKD7vmbKwjx6WK6wua0YMgiaGJg/QijhB
q2ks1+Wc6Lgnb+ssgGufdfBDCJyb3SplZsLCy++LYy/lo2Kf39RPoXZZpQdWy5PQ
wR55SEuXduCtoMu5Lwp6O7nN97kc33fnYSrDBljmn/3+gFeeUIJ5Zy07DHDfBr63
f0qyhOu5oGjns6ctmps9i22ENJx9SGeY8++Ya916MO6Ie2kbAcm6+80OVNFZXXEP
Bl2ksd1xwfZwkS6s4pptsB2EHvAx9lh2x9tHsS6ytE4B4tFUu+CBbZLRn1Yrc3H0
QsbIX9N3HZQ8HZrEzL2MVur07pPJu6fiOgiVfDzfNENL4P0z9wNWJnO62OqTw0Eh
TQI5/zYcIUEG/QlO03VmQOyCQjYCQ3pxbOLcAMTmybyPLockKEKWNzZ/EypL0wXB
idutQAzwe9bpVqCpQAym7fKBIP/xeg7APbD9UYKBJ5PgxsKH9anhOgbmwMlGslQv
hRXMjhMnh2ejiVU0xeGyxZTIy8DWEH0gQOKyPhW0HaIvgwkADZM9e+QNC2QkheBS
i3Gjf9wFhK+rUsw3b2+326UAH3uuFtgUx3TDvGb4/Ts9bPzWCYkN7tYADoMuvj6S
01xQ0qQVAhH73rsFetZR6cTcoih27i3gncG9ZEWJQkdLVBjrHUT4NAvA53BHGYKH
7WBv1abWXBjQ5zoDXc6XO+47U8Y6gMQ1Q0MEFyfUFK/bXOUXbhD2lpa0vGUM4PwC
teRVB+A8ydWuZLcYT3yL8nozN0gdk3oIH2xxXRKdd9FBbE7Ni3G/9S9yOls8tdDh
0nQa9VDulxG6uj0s81h0aafCIu0htkcreH/dF/tp6COZn2d1/NyhLueEPQBGAdwa
iJuhakO5RnoJoHiTamnvxBsfDG4vyqXV+6evhHa52aWTnupKFfG8JO41rBGDFEOK
s69SfSyWbLgZwT0JiTlNW/N6xhKCe02Z1NUAglT+UitsF4d/5/maLMyHz2nuRemg
CC8wir5IKC0D+D7SLkj9ZjgDAHpk5Jk1eshHitE3GSiVrztvnmom/ih7MQyTqJ4O
QBr/ZWSEzawZu2Q910A6a+XlVmNVuHHjJYIaYnkGoo1yQ5kg90+0QJz8DEHR75PD
odSzmcaEWsvucq+HjWe0MxqVHzbUFMYC5m3xPNmXEfJA7fyY00uw6eWBMXkdgXVc
y+ZFitdM77JZ99WtrKJ5wAanYTJR9SjL3+uwAYLEAmoYePZHssmQ0DMjbgbFAZKy
cFJiWCNF4hVmMna2HeGiUuA2rct5FBjk/I3GXzVuyeKKsRTDPpZn3lJWJ7onrP0s
YmgIQAVJPkCulCTCleYaAoF+uVdPOsCe6PaxFcPlYv6CP2b61l0XAcysOM1apCL0
kKeFIaotfBF7UQszxNvPDnB4B1v0I5KD4i0mFoJhehspkEOlEXqTIe0npsexVtPC
pbxHcn9PAUZBcWepgbv6PHxIwcNeVpSkdSTi4tt9oBaUcWU0nn2ARhedHxiIcqeM
3Qlh/udgZRfznwgjifnToG9Wjyy1SzCd36W088JryZFvduxt/mXR6724UtHZTWDx
B8lUhLmmTQ0GDi+ZPBuIW74Kg3jCPtTs3KDrE20kla/qT8dphaEjkYONT/OGV0F0
ZalNlqjZWjzmlXqmqVx+LluQy9E0CON5VVEU9WlzPbgJ/KQ/zMTncpnur3+y9F/Z
pd06fDQIwBVHF1wShMWcD/ZQ+9B8alVcwVF7LWUWHZ4+aPdVaGga2ibNsF5KjN8J
psrQ+ATJboGMD27yV4SPIF2iW5oFy3PP+Yk0rZmSCpQ1AY9bbklU5x+kN37jCkVU
C7V13NMBD9KOkJJBz7hEro/zrb49kN3+5rQB+OiflInZC2Ir9Csq1cElYaMCT+hn
ws5q2icuv9cfPt8hlawv6NvnekhRwO/5t7z0sUe8XMApVI+gNsvsDFYQV5R3jjKb
UYxd5tH00jTOrFzvAZ/v2DwPV02fMORcM/MqfUcCU0EDCYxlPZ5mqFIpUg8Za6MO
s2hCFQd6C/9NRnmbzNUnhL86RI9EPQIsq92Ni3hw9cNq+49gyX598qgJ+Lp1mKfZ
qjMG31NePLaZ9KUdbNHhitsYwUttEZjQ3iYxrskSwneD0EhSMrGwFgFfrAYL6hxa
9/O580rCrpQgJJUqLGxKaMfyxkQRRcyFTXxLZQlIqZYGa4UIu0swXP7aTWRklAKq
QSDwTObM6c7Sd7AB4vQrzFJWU5PdWBUBqyXECr7UdL250vCOOmjs/7Wo79aiUqfD
uY1qwwlavZvdUS1PWijPneG3+9+moK7HNqwdu2At4TXd8WulI/QuADpze/1ByrJH
1f3dMPYIu3BIxW1wWOKRQmvaKZUZH0/oL3h2w743WoTwUjs23+IYAYW5TtOG7zbY
PdbzUuIdzS05qlHj2MJFovqFppxprfAIpoC3rrL47uvwPYmvvRuuu25smmh4CZ4u
dSgtOV3SS1Qg+hoYyJ8+fEwDomldsNXARbvxSA7umNQMsYvUKU13P6aUhNUd+FQJ
E6qbjTeE+SBXl26cQvjiCrhEPwztl+uoJg9/QaB6ufzV+2ynKAnW6Sxp7y15iNOZ
LyJI48W9qXOf2w65FVRDMKiqGXx2fVzKzxFh5nIJJ0RKIiWrohdIFQB+CS4macyA
v/WP7EVYtRHiZA+sAVhkcEowM5obJufrW1W8YLvucr9QSFIzZu2YR8Yxypxy6jyP
c83ChoMS6EQzUVfEMf4lD7TknIpQ3c/y3wOgy4FPZA47db/6iQDT/kaINmPahU5C
CtJ5C449owRCdQAZ4asWaL+VHjK3s5bUkE/oWQusm8mSFke3e5ExU1cmGyrouwCR
itB2uKekiAnmAgWdz+HLSfQ5WhE578mfH4/56Qt5qDgkAdaP3+VNuJDCMi8w6ZC4
oc4N9End88ud0NE2MyxEXLt0cYN1wMpoelg432bp64uThBYMICcKsv2n4oProH/m
bw/EL7xJlQwaVwj+SBK82HVyBshnyI+wfBXFBDZhM/6vYLDKxYvkuM/0q+ZRTIXF
U2Z3iafrEUoJrQnX09bCkfZ+8OKMIydNpDQPrecLbTGrpLtarXtSjgen7wru5f0+
HAzEA0qShAvaYyoYNSavL9Ox/pgWVC1U3FkfIjhsGLEuQmGU5tDEuLI8uT8b2wKn
BHDaOcHOaDLXoNKzWKG50zU/bSbVtLdlg/BYasIbYIzGs+oxF3eYU109TEljJUwr
X0dlbuS9ovme3dYx3uJdnDOZQ3sXlYA1w0x/H1YqfO+Rxn7Xw1WKVuJrhkFqioYR
N6ZDZMkM7g8NLg/fC98qHQLhdYzF3gMlK4AJr9NPTA4y8j0D9ASU+3b2uiy3s8vW
DasMysEKkVQh56TRuHVyvOIYOmZOLwlJ1SklhANRpCGE67AInBTCMzEh0E+czgzw
4kdhpM2Rzyda82mrNoVvDFmpSyBsm6oPxROFWRKPb8yysj1a4tQG9+qJ1E4reh/+
2YOibbi0pwf7iuUy+0LW+pMPVUJsRA8S2pweI+uDeGLRuYkxZEoWh02plAJ6dHac
b3SOon8GsiXDcWtnnCfZxiE9aZ0+rL+MuFkA5USNn2Rbhpa9Z04l6SH+d0cinqnG
t1xpcdE1VmyTYPftNDE3NCgohEJEptJdkOAXol+7mBHADNEQpe+ethxBjjeOHyXX
dV7WMIf9NYnSz2ILnWlIXS/4nae5ABbwH8PHnNglCNpE3DNsvn9y92vYMhSef1s6
O5dzF0/vJ7Lhy5AxT4YhdlJOvOHo5spBYbPeBdl/RYSkfmijsJwMdSibL3SUS3Li
o7DIMEELwplTw7qGAhlOzfozClbwZVWhfdXctZttCgreY4qj5WtcSQYC3tPsuW0X
o5lc31hheH3bU+NIeO0gt4grVXp88KvMnH0nQp656D+x473WHSajQr7V88aUKWpg
OitupSJpmG57QYxZSAUvzxmWc1g271DeppT/bb6vmIjP/v3CoFGw1Im2DtS0ZzJf
42GbAeEbCTfJTgXqvAlwj8hD/XOEfegfmPW1NA+bCzw0SdaAG5LiNM5dgtPEHvZz
xqRFG+Je+z3Pr7Ozfu2wvkiIjGBMf599OgPGSea5qcY59C2bJMcMifi4J2uKkFl/
ZOvawAqSacGH02ny75tmnnb3plawA1n6hvFujKuJa0vd2wYnmYA+CLQrnYm5wEyB
joXtSjikjKo8OLP22uneq1PenAx+p5fiKlgv90LXOwv4/ttv5K7lQzpF0L7tp3Rx
a7kVfZfvTOVmxOAFGVSFZIN7y0iGuWwHBcRNvSxpU5bQJYBieEPenKnkrSDMZZuF
vopxLsRNqWWZpOn8PvHtJUCvsnYuwqFr4FhMdlc56iMkMZxagtNFFJ7iCupfWhTB
XuKwRFpBifNT5t0SBOJCtGZKtD1AJ6Rm/8LfzB+13KgrzgsOAL9VrCOdttrc4l4A
ERkRKYhvjpPDC5aCmWAtbDrK/6TwwuOElTBj58Um6G1urMBIPRM6eS8y5ZI1XKjs
vJpm/qUIQJUXoj6StbeGU6RGnWzwOGIT2/NChkKa8EIG3lGzXE8MNUly3CQSAysE
tM/TZOaNqJ4lf9VcGfkA1hkgotDhXHHgHj1mPKyWslOlBOIHCvrMv/uYKgWUdeX8
DuM0TZ1aNzuRY5IjSEV+m3KswgtjeuTZbWE0Y4pg/VggLYIhwrfcSztwTjYFtwyb
rrraF/uZq7PYdNBVgoeeLFH6Ct4P2dqOH02s+emPWW7lQJM2OqDUbh/e0F594+Cr
hPb8PtyPcBuCE9V5RhKkDMp7r2H3Yoz6ILLVuGkgIvCn+ypXH8Nu+Qv7WsOF97Em
GF22BE+gSx2b2IqQCdhIwhD5bqe10iOvButxxsAwNdnf7nh9Wc6bhBIG+qwQOwyX
w2L2W8JKz7RqQCUHstUTYoEyHfz3QMCIepmOEhN4Di7vzF/Y70d2YboaXXNYdd84
V6NqkotY2jhYTflFr7MpN+5nRtlusxzzWsu5N7hGiSJBk32N0OTDBpxxHiGy2n0j
evMfpoy/c7EaZtg3KlEHiFzcmDin1O6nwdGko4xHQkyTpIAlkRQASIjzQiWXmT/i
EyR2/Zgc7JJP1HB8wFXgq2uQTlrBZz2NU2IT73Ki4MtjvoCCZ2OuF7yddYx9zVFT
K6WSF986+hvKZned3O8jibtUQZcQXbQtYtufnuVNqa77E25RiSACJ5fpq5lPRs41
NMKHTkt1OxD+Up7b6Va9AfCqjzvz6XnZyOwoDWAhNkfSAHr3cdqK3yj+i3eUQFEy
+cKl+oYKog8ljiqsl+4iaJH+bT1KOe+fzDKB1iT4XT31rk0kDQcm9yNBWpg4kEid
lfv08HmHo3I9gi0kgj8QfpnY3opATGxdYZO6effQ2yH7cS/MWCvCUFD0RV3Q+LkN
R1x74Gd50MD+YzIlwDdCXb4msA6mgX0R/tIIA71bAY7F9xFXc8XQ+oE+eEg6tQa3
FYxlsbjmiPovMORsEPoiHFHvtyMIvL2lW9esgrFWNeyZAJJXqcThh/xl2+HaMDF4
H1aNLOYsSddK0nEDdYaD1Re8Ntb9UP00A1XiBJOgMgyzh8ukCUqyRc20AHQEZY6H
Ih9tox3iz7aS3WBugk5XvHDCX0Cz5+DwBtSiSFbl5pm3fVf5HCrxl3Z5CNci4PAd
Ym3ePsHlSNBL6sa5gsTMIFcpZOr2qV+bl5BJ4btfg3nCQKa9ejxCgmNGi/LtUMpI
jjY46tNpUNFn26+/tAzDPvjFC2GI03M6EMCaZpwZHFfAg6HoM6XnbYnU0g4nM6kN
21FFSAQC9l157VmnoyzgG2rarcDRQChVEgrWrl4sTuh04j9GAfbaXM0cug2R+ecj
1BOFmAbHHhXuEOMIvihpdSY9Z7tsd4SCMNHJbjCvlhOfY77digoTjBZKnFBQPshr
WeSeY4UeKIF1lhXGPyBebd3v3bzh8qayKDLfn3BjGeowqKyiDtcIYg5MdgUTCOof
U8epeSsXV9gxBXVFNTRxOjwy6gdLmq2a71c8U1UCoAuXEgEMeZ0PnSd4PqptaVGK
PWr2egfPilX/WBch9q6Dr8uH3YaEPoOIKZg+XP8TtYxFl4SW1YQGIDdzVj3SEpp/
vkXGsf2ZnVLEwtVyGqfOYK6xKItruZ2fRcF6CBvLlIHm5WejMtcCc+p/MxzVOaBG
yPislnjhyvMC7CGqNkKI6BHmQ8pTvJJGsraA30znLY98juwB4z3Vjs4eVCr5yudW
AjofycXQm3BqO0R4UefdADmVDSs9z7ic7STp/JstjEQG3kpG8IBB1TUBuY88L/W1
6NG7067NOZoXEHNnBRk3VRBRovZ67rL41aChxxqPickVwWEe/onTOSbWDK7SLNcZ
TepOZrC1skubhWhktwWy5KkAYV3k+FX1xbW6ZosfeyPYIAccW3LliArK06nMSiFx
jyJg5FGcGgvVbzG+/zr2SsqvID/0VzgWDSo4CD9JoYnP8Fv1q6BZi2dDfl5qjQDX
Aj/w0mI7cit9fS/sGQQxKMKPEh2IheZWywlCVVKto5aD+9e0oov0O+RWn8Z7k2h9
8zd8Z8TYlcRQ0w/np0qYX6RdMej6Tfshp5Mso1bJ0DQe79UUg7tdX5QdMogf9eGW
gp7NRRjN7i9lj9F5TEVfEAMyB95FkhoU622bNVOZKc2nMI6PqU0vpB2bnimyXaLT
6hNeKf2bxhUi27vEyKm0s4N4W3rzjtE+FlSHa6mVLYCOKUw0HdyeOxiGFQ6MpvNn
SELirKkE++6bVe1gn1oHJcnIZG9S97MILjd+1ga7DkTfQ7UTmGG1S8LVKHiJ66NC
Z2B6SQ167OjtT+rUN8dpAuzAPTtrWP9UwKo9EfvHH9Aq1g6uyA2QV38QlBJTZGOH
8KOsTobHrZU5ZZcN/x/yygZtWToSFdA1oB0vMf85AXX/6n88l+/+w4TvAPbwWP86
Z8FjG6f+tG12HDReqDKnKj8OSOI+zb4zINxf6vfIQWPAJw2rN7r0gys88VFFQfeV
EsGJEItJ+MBYbWF+xmD7SdfvvTi6BQOEyzp+QuumFrEMO01JkHPKZmz6fh4Gpe0s
MnSu1SL0DvfUGDvjyAH98wzIK8RkAxpcJgcZQ0ikrjwsrlOZrYDiCnIyWhpf9ZY4
gfbbZABDxl9fV0gslZIXkRCDwnwqNByADfY38ghv1Dp7rIfFmNUCwZAYKunraUtx
wxVDK0HdBH4zvMJdCm6hZlysfYHsITr+nErVARNv0dtZQiO4AukV80n3BDDHpdWp
403j33e1280771JfsgnyTmfub1xLx6FpKiys0gClJlFGp1T/NwHhfNPtGWW5RWPy
4Qhq/lz/Wnp7ZQ6vJ0oaFTD58HiNza4PJstFzWrJ4n8ArCLYqz5Xix4BIE5RUIvx
AHgfj0LLmFnjCYCcF2185etR78k4Ht3bbfnimG0dIj5CUoYPZjRdqdeqLeOijVj0
hhn3jqK7ttsq9swnyf5TfyTfNX5bV6j7QJ/BVe7CNmP8HH2f0qR2MaLgb9AjAmz4
+P+Kjbp8u2YfIwbGnE2gBbfRYO5i2gvqv37sate2bRb3fjaRDEsGeEHe6h4Ej/LB
vUwJxgwvINrNfEVPBMK4tGLeNJYKUCSjs/dei1yI+aXzQEnWzSWL4yXMU52sL3VE
rlOxYEx0MF730i/6lMoCzbChjWhEuGRMQoNzXgV4EzrX7JmFZycg2ObQRb8l58vX
88ABQq7dSEP7EtBf1En+AOHVyUZwlmv8NOSyXMmmUh1+CRj3fl9ShNdNaOGo7NoG
24lEDXh67zLL/3OGng1BBofSvK8/SnTHa9vFi843V6/X7cun9tmTt6J2LN8Uhn7e
XlVPNzU/mI4SELctapS3mwpn1LaIGSyD15SDYs5NiFLDmVfofMjjmvidAmxzhoPj
1KXOVtsyZHBX+Xex/xVDmd0j+6g5WY80HprEs/CgPF38dHXad1u7Ah9vyb+UAcpp
ZUmB8tZmZ5LfVFioPqhcsTgKQ4mxyDQy5irQiWzAWKVQzW6xKpDMkcD8vEKdRxsw
oxOmGA3oMQxzfPVp2Ea/QBvuM5cCF85gMdVank6mZvBO3Ngkp3TJ5HhgYoHFLD0+
DG5jTlyalkIf74TN4Xl3sPZ4PLmR2eDalfIjGw3lceSME4awaxmuR3ugDeUwdiTM
0RcLQBgM8lgduRpS6W3xvVqVI7bMiugtVNTzCNXIRc7JSGqNqs+550yC0wpWeZZ6
rbwtExN4MzFaOa7oIhb3m5gFWgGmJeZGKRIi0JhTWqsS4PoQ+Uj2sA4jaZKb2i3x
2AIf9KbzUWa0INDn1TpNVJvrOsjPcuGyjaTdqbNCDCGDIQY386ZfS+8j8B+ljQLS
bB3CViLqKjIkJ4lAK9O48trH9Ik9ralF+MnE09m4C5jny93585G0gC36l/whzzeJ
xREiLFVjzae6PHt8TPIPskc3pjf0Ae1E0OuefZHbif3fLLb/vOJ5Oyk7GeGXVszb
um2k4Vycq3Gtqf/q6v0E5TRBYqyed4aZKhGVV5+yYIDFtxzA3/R8pv0MGkYZM9Ft
iS4hWz+OzGGzID8dUpC+vmCuVp+t9ZDPyZ1cT5QTPUsi2qtaoOPvyVUoJHxMtvtS
l8whqZi+ab2FJ11yg/ZfGsjUynyiiYdRNbCurBoKv1a6WC2HmzMHNKV9cSvHZibp
MVgc6Rc7C4/qZS+oCZiirQfrLw7hmqDSu57lflWr7iFt0Zo1e+qlXOopAu0rqS3p
D00oFyGvpJRKvXy+ls1rsTl8CZ8P+ZpsUWa1pYFx5YPSH0DO2G/ZYrrHZFmhTMHL
Hqv4HOX7yOTglDLM2CSlNmmKKFmajSsL45hY2ulj2D4yComLgr27bRCncG/KfB1u
HqYF7G61K9MG1fUqjuDKpR+Ps91YbHqScRNYneCdQZjaxJo9LaM/ajcf79nLIALi
4IclBLHJte3qnDk+TXRZiOE3BW/phFrXDBQDdY518I1s+JgaVcjpxwNEM9XzYaZU
MqS53W3vomLcvcPFV2qvhvmWaWcoLhfZIQflwtXH3gJtIBd01Hux+/8TUFGTqeop
sbd5L3xKWjKaHa5uJKI8S3awx0+9UxIMr9tSVPidEj7PVZxZKx3wvYuws00roxRs
BKedLRQHHA5cVYA2xFU9+vb0e/SjpRo3s9G9Wj8w7Z0IXQQSSRIJLLfZhnZp3o5/
D2KmSMKyYJpFxt5i6hjf9JMrIifhR4nWj8IS8Q75VRkvR6ma5ac1hypmu4t/X5t9
HW0PBsfy5gd0IlhHDreq8kcB6UqBSKZtwTIrPu2CJyT2NiFvqqWm6G01ehy49X47
nu92w46BDTsF/7p5icb+JbabLv388i78ZB4tPFERNqu94sQ7HxjZ5EyuJGzh97nF
ZbKNgXvdZvAigqg/VoPPsSDzZpr71fGwjhAhmKHTrCJSiTZ911/MBHfboCyRD0DG
kzE3sjQMOFr9o85suPIJ+SyANldvEaVevskkUC4YW9GfTg/rJeYMhXxfaYwtodvW
rzJtY11ktunSJBI1qHozXwUeThF/phwoGTd/6zH/e2sHTVGksq2UZiWGfMupr5IJ
qPVh/CfZXQIdufzDCxl3RKb7L6/2JfGc4U/TgVEsl/PYAl/VPwmTMRaVj1M0klaF
Awr3tixLCut4IQxFrsyJSyYvo9ADi3ig4bolO9n8UFUPJSgadGF0obi5qu1iPXIT
81Pnr0iDndygaJbEuy9Q+6WACfX4mG+oMaAFowcSng/H7U3J+2DSELJIpDa2MAZ1
NHo6L7SJhcdieDlGuXNPq3V1beTtagCUDVBcJm5P3v9I3WvMoAz5t3pu4iJpXt9K
bGDOIbowv7za5gkaSNfKxcl9mOAx6zccEdULfjrn/rMo7Wzv5fZ+g13qdN7h8BBG
S+jiKAv7E2qEuZ12HXpzc5+DaNBUyjcWS0gI4u9M2WHHnZ3U/r+7LoxrKB4Vfv/H
pA+uKBeGFbmNU+0BGB796jvzUiznfkoS8fGRghgzywGoG6c0mqBVrZXeP2As8Hei
ic8QoGwf5qLUgV4ePSRkgMlO06UWXIaN5sTTTOL/7kqXPW0HlDmvc14fX9DJJkyw
NN0Gpyzatt42OIS/stQV8Xs3BzxrEiVIecyokOWipdqiu6tWJcJGicDqddSfgR53
eIwweipJxL4sDngzcHGBL+XXcS9+XxaeRnHMxOYHvOzOJK3nrE0soLBwr1MKPIkE
cvFTSEz2PrvgPQjYnus/OgYwT3iWDZROZarXZH+tNBhJrRzyGR3qqPeIhsqmRf3t
UXxJnv/8rAS27+g88AWlePSP1tIFlA906l+rQHF3YJOvC3lL8Urq//TkYTOH7sy2
eY7J6045jTVvAC1lT1ytwJJMOpMj5dJCbz9jZymIfO8WMedciEwg6eVe7TBFCEwQ
TyeYHYMsFWMZfKI0d7ghYU+w0vmquPGwQMm99SfsSzM+8TiUReasttNUeZI7FOWm
la/MF+0tKRA0q5DoyB25ra1pLgTV1OJr2qJH9qGcKj3seXJUkvkvCQ2Au8909V4G
ronEfaxa1v2ltAnVeRqclLrk2UcEx9T05VnyCowCWk3bM3c4TzOUyUrMrf10Yf7X
lRugN7M8YxrM/1JRktPyk23Z3V6/74mwlrRgWf0Vyng/p/lDGiZuRpzaVZsNKWuz
sfCmB+yNQsE4yUb5d9RpmJlNG21HBM09anDQKXoSQjXM9o1bj3aazVNLqf7lMtlw
kqyhNg0cWqwwQ/8Dv+Clh0t7sEXKlNW0mTP9CFWkgyrNbPamtaAQmLOddY5glqal
7PGRs4yfgmgVWFUYWLkEUwDktDTdCjZDSq8Fc0xj+gH630LeNaR9W/881hVLGdWE
qVDc81rdKm0hqHUKWnxnG20tn8g0/J6+QfNRAxXMuJLiRT+TBX1y8ti5sqXQgJg3
/eUG2Seu0xYC2y+mJqhjSD4tcyJnodgPkuDN4pSXoO0V9ogFmbwiV/4lybELXp5X
aW3yj3rcdUh0uxsL+20u03oY06gQCYaEme1iobqiKq98ycSoYV5S/yp0zr4GDTWQ
/HZ1XUDKTNXmUh4obcSIs/jv4cXGkWMES7MTqfSxi6hG4VzC/zF+gni0NxMLh5Sd
Y3HpXwSbtBIe6eyh6/1gXnAYz2annxa1/DOMQxgXa9nRsaLpxUk66ntaXrkAhIuw
RyLEtKDMgrY1dzPuVQDYUBmDC8Z8M2Z/NLjeCC6APjxBVQT9Un9Ih6X34+YAybXz
jW52PH2gTp5Jfmfo6jfsyJp94QryWFL89V78sv/RAGuMAXS7+LUzAXX3IBbmH0aC
z7TZG2+KJxuRlFovwCUSvVaNSuc/eAIbZ0iZz3LB586f8GXlKA9Sd165Uae1/LI3
8Y02SzsVAdVqob4l9LZ53YfuICnZlAy8AOtcHAZAyk8uovo87IYykjB40l6Rttjm
boy9TpIL/7yGdnkk4vx8IS9TTYokaX6zo0LWcCXpx8aKl4iPRLtTgZWQ1q5354FN
wuAThzCrFLxaSoGebNoOQii+w/bUByE0g6+XUhIkW+9Hz4hJ/ZWCGLWIrsc+qIxi
pJT6z7COI44nl8ByL/peKanX42T1lqjNgzQMvYdaoLF8ExNmqSk/YlarubDDCPGU
Us5nodPGJiWgdRMDcnE1zaZkOkjUTLdHMCJHwrf4QleyU7UbEqRL2BOzg36Eu6WB
o6SJvG83f8ILEkLpvfCSd/KzuyWPiLz9PHolzVtczI7qkHG8gM9yddoC/onKDlkP
IxGaXvwaVORzTPBxADy2skRhZJSioSuP7rhhai8J8YwnvHPfYF5HkXO4CeYi6QVT
NGRSpaqWHA/+ehsz6WqUFAXFKmsybcmAhBacnKHmajg0F+WoYpT4CG9BUT+Bzl4e
3K72uvzsUusA+/8I2isIdgPAVFIkxnamTWqTCo7gUvLAugyPfCLl97Nf0G7jzu0U
GTETkuTC3c7WtJuOpxC42KdkTL29/hj3+T4x3aoVZ3rzbETyXmAkzN8fd6LACBnR
hV79tHPKDx8zrZsNsB8Kb8DNVv/ZMOPg75ObRNKF5nX6sJ1ml8VOncFy0C1/JTik
0yp1OMl9GMNZAyZp+w9sDRzv1KM3NF06rca/H/gVO0MEZ1I7F51v4lZt1dn0Rqm8
bBHK5uL/05fYJkNZu2oGPJ6JY6OEZZXSioC1BjDl9/+t/h9n/cwZWvTyBGL9h4DY
t1FZcgPGRxBVTeIWv2h81ZwRjtAYQSRwgSdwi7OCbL8ePi9U5ALKYuimS0vNo3pa
aBsrH0xvYpMBpIODYh5eG28bOCPeDm2Pa59WA4RJwnn37K0WAwwcdRPLcmPNR1KW
8pjhDYS4GX1e48LJBeQl1a2EMBAb5tMh31ZwT2dPsXO8qZrgymfscuOS0fnjSZSV
jyGgdoRPKHnfCJgVi3yFOYmLEqahTAldiRmEQ2tqWPCIfNQyEQNuKUiSkD4hpR/r
Rk+uouvnPBlY10w2eCN2RuusKGKANE3EUSKEjZUNYKyW2SZs4oEEFpLrIbF1BO6n
dDa9ge/CjY/TYKVrMfzpzd+5QvvsKm0EmfvUx1jpHdnC1YgnRmgbaM/43+QQswEz
ysNVA+hwvmy4SNsuLY/1gWjKgLJQ8jFkM1vkUXdEBciWUcyX4XnewJJalpyXslf+
P6TkXwGH0td9l107cDTqX8qaHX3hLWMSizBLqCEpRUCv1YdPqpjJZJs/d2d3w6F2
NY3cOjYgO0TM/jRpeNW1J6xlsViDCjC8uI+E2VmCpluOENBr+BDTvfBNQkoh6H0h
WYg7/44Qy/xbAI6mAjMxZIRKftSPDiToaiBlw6V83kbruEqR/lEM3ypASv4bBBVa
mG8dZ+kr1kWMpy6dat/e1V8++tT8o0BildsCTvlxi3Dmjfm2ZY84iYyYFVnXGz7P
/eXHlrObSUc8d/ddbZ8vQGacrs3euvlD8D1RlKmLQ/H6WR/Br6VDnDxxom/KrUz0
xLxxu3XtQ3OsnOgKSYBgg4Sian8lWhcVNG2K7sW45Dg9M4xUOF2fJaR8XkU3AwG4
0Dxwji9GZFC0F3WbyolFIKml7uUblVfcBXZbW4ItuaSYeeu2lWXgD0aC14n9aRFA
4UqkPugg/KHQLRSKg9k5g9fchJwHq/k8BQkICqx5h7dB9fcI72whmhJi6MPliGGy
O52PqWqryDnoox4rCE/838vRbXnR47szsdMGp38RYeVga2mFeFBVv/0QYs66Ad1v
aQocCypp4cjGJT4bYl+GQ6Y2/wV1yj9QryemypbfKMCwbLlczMB1/1sVJuZWEV/8
RA7cqNkhYyYmxN5QW9fx5yQ/u89hKfnW7KHiyy3JJ6dEHNAvRaQd13O25TWVaRyV
LKVhbp27OCF/pZrxZibfVOQNGghBJne2evTq/DRmq8EbBXzmhAo32MtE4qsMs/di
U+42ObR9upID1K075f2G1EHApynP3gzSa8gcv78Lv+1OQ04m5dO9qJ3Upd2LVEWU
AKol8LepukVaKfVY6PQrUDnnfnH6BhJuxWmSISQSizmgZQRbzhkDrP8cTu3DnLS2
9bu7lAQiL97SNVF8fS27oCz6Lhag9JfVFMDInFx8nTVFQCfQrtMa6wY/aeZsMHs3
QqBH9IrEX1O145+k46IMpEWGgWvS7BSqTk23HeKab9yERDRMJTT0DbkBY8hD5Err
OBauMuA8fM+ClUXuA55Co4sjwiz/EeC+gmmtUHML0tgrK+8hoVBH9u2+RXFC/qno
uUujd+mdxw50u38oOJK9qoskBoXBTAo3Wa8Z89wpJPx/OzeRneUsKCBzXOvzfIsR
wNSjxmLrHwPLYByNWgiK1KbidTb30Q5ZakJVL0ZRE7XHzekADu9kabGVaRfSJ56d
ZbIMfLHiplZZJIwio3sIN50v+24kRR2/cehVqGqUu0+fBTchZvAlkfxWxeQRiFIj
p8ZqoOXUBiWWDDtvE9HdBc6guc0P/E5ng8LedNmsEIxBlW+pm+bLQzMCG40idhh3
snVe+uNHmN3y5916oIrr73caZmiuY03RYdQA0hs4zLBD9AITd2YY2o3V6Z10u/Ci
HlsI6vtqhbwKTGPvA58wZG0XmCY5ZUdF8Q5ub3Zv5a/kNqPVfzCqbzT/czquraen
igdpMN12jTzdy+ntgNc5QN9in2/gilkPLO2ghn+L0Hwluu5nAa8Bj27erRQ03emj
oemEvn/Rzr0OGxJP9G39KEwHukkMHmOpmUi3c0oEwFrhcUfzyQ6BHpR5QiL26nT4
/m+XuLqUXfQBxdO/bUv5lATohbpM6F8KBIPDdIENqBnOEZ8xzLteukgpozoIPQiH
K/09TF99BXw6mmHpX/Tv7hZUPOFEEV0aDWcABsNgArMWWhxjMuFSUUycBvMT+278
7Kbmj4HhjCG9buqc2qEFLxllf1UtR8wnXNqC26qavjDQYUkYKipWTCs7PIOsRCem
S5cCjbZTyZomnR3kduKel+yWCWTyOnWlfPGRIaXozzWwAEAM4n+l4fkhhs+fsmAy
TFgPr2UlC3bcoDsxyDo5hZkK68oh1Dj0sLSxq+8DLFgpfmA5jWg7FXZmaHPD0U4l
ShJhFgLSlkhZSuhMicFFKXdlf6XYSxbZ+RGb8pV/hqAcvGiBob/TM2HB16CZqiY0
wji1dlzBCj5JOBcjHLsWni71qFjH/s2BOf3onDxzZiFHbWjCU+Z5WHmYDsFzYU4c
ZoiYBy4gRjqqdePquXM0/iD6fhJnv1Bfpb/O9kS6DsU0Q9XnuWdcU04n3HmO6f6R
5ha2/sq4kSDLcqrabrpNSRDt1qhE0Dx2Uc3JOYRIHnEFSALYUG3HNV5n2IfDi5mW
iXyvuoPtXPxLKEaB+g4+kJi5PRnWuQcDICZSoqpocl/nEmU6ziYJx506nIQtJje8
Rk1TsAn6OXiVN4X0iK8AJRIkMxWqVHNPHllArtvnXm8xpBD9O7TBBo4W5iYfgCpw
BnZb2vfMXWz94f3ZI27DZFgBh/Po/jj9dK8EEXoglDd8cEf4p6rjWMrwXJgmqIWG
lvxx2ow7AhVLc3JTPjiqePtE2xUheKDdp3RPyAwFeVNnu0fwP+zUq2E6z7zWGak/
B4Ns6GZiRLOqTNnUmXibUQQL2edcJ/6jdrsFtmgKmXU7KBlF6vI2R+4sOR5VYmjz
zqmG88/s3C5DQ+OJev8Si7uTS9Pq9SflUMnpGNCs4rsN1nlSSCKdRusFljKSvxFw
qlR5pOf8Y/Cjqyqr9QwXalQM5mCUOCoNFAcM71pouuwbxYsrQRjt+Ul6CRf6oQPw
0TbvVHdAdYDbuJ88Zy6yv3NPjswistR6MXh1R2DcdxCoddsKaGWSYwkMbs+krixF
jdCsnkb613KRl5GxX7AeI1fExdn4+05vhEImoluL+DcXk2RMFkh/afgK3uhu0cFs
bdmi6uykFCB+F+WscsTD/Kl62lYKMh8YE06PlYAPGHOc5UpuVu05AFRkFYEBEW3t
8mL//dX2tm/mJeKlvFi3iK4ofkk3KWPV4X8shvCO07g/wo/7t6K3zy3EAntYxzCz
mZW6d8nGaeF0z8/7gkVpFWkj0fyctAvVabVBx1MyJHx/nCAH/Zx0ONseMx+XN3k3
523ZnGLKNc2DnXtj1BGy0TKRhFHH3AX4kIPpYRhBNjLbFo34MtoGcWoVlqJAnkOA
Um30qCyx9ytKzklzmJCpm/ccgV2GjhMDQ+oHJArnwl2mC3FzJNs1a0M96kQj0kiK
kNlFGc2OpXfmHEYW70W3+YKign8HVP9Lp2LxuuCaCA5C/qYH9oFLXs6zYhidZk9v
V3xrmlIEUikCwCPYrE9/JWvEMDg4s4ItcIx7+YOR2FWiv9CGM3jNg1Naw0+l1H3U
miDDDVxxmocirzLe+jedy64EmhPU+2vcoIVNQZ3Ehks8F0fShaOiySQ3TpD8MSqM
HoVO25FHHqzrBBfsQXT6FeJkgQccbRL/XbLQRMOiZbzIE9NCxa87kmEHQzd6pVYE
ZMtW243aDqIf1qPdSAg2HAJFhfF4QsJpnKX7G47fEjD5ojq00Xt3+HuSU/h1nlgb
WGMM3C9deAmcaCAJKjW6E1KZYHuXXuXmIx2YUHxzFXD3qmrT9RaU/LiY181zi9D+
cwTfmszF2MpIJVpjlZ2hSWNkJCqCY14mO/FGl9dcki7w24JJ+0O9S8MNQaBTT0fA
JoGGGxRrczgfvd3U5ZDxX0/sLqkuyJKMQhPsrMHRspfJFOVge5NExVJZdGg59vvA
GQuOQSMLdPynuWFZArHrW3IWZ8Br8+XyCDYsgz1c9YEdGwhEc0Y08opJ5XZqMZxc
/Q4oKMPcCH+s2+qinxckif6jCF0V1odDZNff4NDUg/yP0OcRHsuWhyGJfERY4ctS
AWkWvecQr4eQ+LpAEoyyF68SiXH6IwMZLS1gHmp7HFcaeFPSdKlBXPjZ66DHEtk8
l4thxXiVq9rRylr9cIOV8XPV8+EYriJVl/57IWNYYFUTNuKdOaC4chCT9/JRUO3W
fV3UDt/e4JUqlWb97tXpOccB5xwcBcCacd+gp43MJCn3/JjMhZs1FhSC3DsBlw+S
O+VNjvM86I8d3IGX6cqFJ5JCM54AnVCdbBkjvbLidD/TQIDYE14ToqRsUuSRLz2B
REhxJa0Vgh32wt4waZdESgkt0qCAjeVCT4ZNlLICCP1xp6HT9NxV8CYtNuyfY+vn
gZsBYYnz0aiAntKFR6gof55oebQkvYY7wAwkZVcNhiMJvrYfUXBJnUaNajOc5riX
nqXRlXmCV4hAy5VyMvAGrw1elG/toNhUYBty5sbtNpoEH4Eb6rKVjVRMQeZOCruP
t13qdQwG64S+V1uyoq3gflmI6WUEB+AOyXfyYU2NwVVaLbBLEYXB41lflnumYrYb
LGlg6gYlUEHXejzDEWnCi6xhN5Tu0KDsT2ztIw7U+tnyOS/1nPdS3yJOSgx96LRP
CAntv0M8211gm1RLmlbsjA1UYtBMGFdqthPr6wjIhcPYZFNb51W2Pqy2CbgbpIO8
eXyhpLtj2gjHgHS/BUlukTXvOl9lij1Eqbl606krqhv9rGRGGHMCE5OyPBSXHEwY
sxAefXXvU4UltUXrdIQdPupm8DyfQT+rLQQD7kxvfBUXNGbznM+OXM55w2XC2lhE
6R0AN/m+UEVHLyKRf0n0W7LcM7+gRm/eUnv6ZbtesgXV70EqAYRp5VyJffqfFNsw
y/wIKAib3wzGLtD/75Ld++DGRLqyhh/IACD7hYo5NSWQzRaz2+G6afvs8b/mRLs7
c5BRJhjK84el44hqLoN+KwT0LIcwzrVJTmWPTCQ/DGsv7i7B3ZZYBj9ffLjy+OgS
15SoSSNgxxeD0/4qLbdp7gf7gO6KN4SAdq7MN9XigJVe3sswd/acWvppzZaH57qR
2lMK/wzincqp5hOK0kvYuc7o+aPnUeWTyv0flX5eWNnQLqdpYoWBVUsdnguSvBuj
t8Xpj9/CC+2/EPjfJxdMkTkOXzRYXa91R6V3LceYBeYAF/sl7NwUcfxQ3hCakEwP
BEjjV6Mro4/CbPglOtvSmaIXFVzr7xqzbYKPHUciQlHnd40mC9PoTWVtOr2i8L2+
rNn7qc8e5KTh+p3reTuP0gY2/R4VHlTzItiX7E5LxNiQwkZbFyFnQ3uxTLlWsaAl
szkQPf+zD+t2bxVCoXYVDJJgC5o1v1/UJV2jZBzu2U8IzUTzyq2Pxfkg7U/9kOLD
40xOX2SkI3OGqw+v78eE7g8aEyjl43l5a7Gj5upGxvDw4He6yeMPGwSduvtopYJu
wC20NxbyZ8wNWNWh1h9Cw2uB0ahteLrUXEezke0HJpVusOO7dAQbaE4ps3aCWsfn
leUsL0HmHbWSvLDYOqM+rcFCSUrqc5/eIPpOA8D1kAEjUXcJKJdoUWceoM2Mj84s
bjYS2Nhe9aM/+dotdhh2yLtA3BZYfcJtEgeqm9aI8HhjBNCpO4NAPucIw2f0NcQP
pZ2J02mYj/IwidzYdDnJPoqZIgndXGoEfsI56h7tpw7GUaiTGtks+LoP9eVAG5CA
3b1E0I0SwWpTBNlNwvsE9Q+ljOIxyFyUMDNLE1+CRhWL65QZQfuPET46F2bQIL3/
6u1Sjr5LcZR49IJxRTmnp6hw+g0WEmSjRTTQOG/pl8H+RoeoRY0D7X4wUSm6JRhb
ecKzQ7FOKL6YjMiVKVG8QNgjqzgljR6d3ace6AaweZ8masiLIjPz1yqEybm+ixsp
gC1pY4cj6irbYikpX8stIt11Lmsvm8j2Z5KSDNGj9zaM/9hjrJZTCzbVWIHWjB7L
ttvO/P224YpPkUCS6layOdZRU0auJGIcWecVZlUCggw8uK4ndGZ03+yq7YHfVA/V
uEablSLUveeXwLc25EqUlK8NMZIaPpjLumGhU36HAtgcVB0WqZd7cT/Vcf/dSCAR
ZMNqcY6dn0lPU+X2LRyh30+Ez2FX7NYeZnmMPxzHDzzxlGboQ/jHuVT6qFWW9Hqr
tWIq2ozWOCU5+ZTvmwoKsGs3Gc8cQ+WVVE1aCB2gAjnsGZKCIm5dvJWfXbqNa+Nh
j+z87RYzv2tn/MDRDFLDzxdvUGgQBbYT45fgzQp0ICByLundLnPA/mp120JRK/nI
+J34pSou6x2eT0Y4iA1iKKHKpifBHO1ZlrjcPnjNX4/GOhIKxS/7oTQFj1Y3mUKy
niDDPKhDZeEpxNCCa8EMwkb8ufG7JA/p0kutNP+pCOFDDPDCSiHYkXR09Ttllyf8
keceM1MMNfRgIeNL+tgWivysQn2yNqP4xzCAJz8VsUFnc8uc+dVzv07Iso5ieCer
3jXhFTFqs+xMu5nIat9UtNzqFD0PYWIMKfWPOqSgROnv0XCv+UZGNBNIE2nz65eK
dx65c53YlGElWIPxoSycz0xREiuxsziyiTUB3MdsiS4g7kSZmpZNmp1sIECl5Dgj
wn1FFOEWA+ni9Ts+uvzz+eUHQv1G/Uu3JZLEdReSuOYWPmQlyk+uwqTzkFa7Ym4p
UQlFVLz4WJBln20YY5WXelPjvpslj7T9efRxKeg8I62ntqjHLURuGCq46IeFvE6l
Ei6ErmJztcMePwJkUdbnr55p+ZqEhBZ7aLWnO5ReZ3QjfcZM2fsAdk5FgAvMP97Q
XKZqr7uQ4AU8gkUXdfHShPbSD5W20ivSZvoHQ0V88q4KtlKu2D982xq7PNtzWPf7
nNqzZDFtlhttbyUmGrog6a3YBBSjp+rphcjuzrLvmKU2MEVr7Wg4i0hoLZHwlDtj
rpGdPCZDpFgZsKzBwlQUpDBkw7qDlwoJMVq3Af5XcNjJ/zpSP0gHgjTlmWVBLxiR
o/kOoBC9Nv7zn6XVvKbdQj5woiinOllmIcS8C3xVH0b2ifMfEuuPByN/T6xDj6Nx
WD9BQROTNiapp2EQ9lnazvPshYy0dXcntXv076+UNzOzY0F+isSi+zPKaTIWPaIP
mIZYokhKR9ixAlGWFdKKJHBfeOA3z804sHrViS62b/StE87Ap7yBACoRcaUxFT3g
y7AVatzWSwzAz+I7YlJx93qMEe6gX+bM98gBVKDoDmtBnMOyqyrjfwuYOupQGzqz
8QrrAcIgkU+mx4eQFLwRz/tjrCAwUSz3S/N2BUa13WLZQN6ZkRMNVkkq0OSf0Fxm
d8hbPZ9+avYCiS5LySFhDOIrHxiILMeL3cTRiGS6vVbftaV3MI8/N5RvjUH5vN4c
7xlMN7CuqbDpLpyr9Bj/zR5RvnCo8zwmavaZx0v4OrHAyp787zUQwx5BtG8awvxr
iVqG1W5j4MlRctkVis2MdpS8LXXHUD8xxq5u5c4JKxVF5bYrHyPt55NN6YCvrf8F
UeMuuCIDBeUoUEx6ZnCvqK8jGhgoxgE9NBLp6LdtF59UCTwft8NG1+a45Myc2GVz
x0cJxQ29Gh8zY5b50DQWvzJNi/RPYuX688L5+U0dAdUSnSOqbZw+I64yvuQX/tU7
JPFmluWrYVrUgssZWc6nVGoqL20D6fhegMORNBZmW8p1yajYehfWGoepOn1PqwDO
XmioBDQVHmkS2d39oKoFNkPY93VyUoIbyjRjn56ryU7pf3taZQb0YUf3IcnjqEHs
Q+BNUi7eTGf1FktEcKvUj7wM3/tuNgdgpZMz20rDIrQESaWdHwFLPn1Lf90dMUT3
WVxSXqXQNUlKSL/kGwKZeKQRrOuADoWewunj/7Y+nzlTic3mc1+07h5VDX8iGtld
w4t6tey9ehrOvuv37DAxiFcnBeWTn4Kl6rmvzuA0gMFo6rXCwF6C+/lAvMjovOuv
P5Qbh2cg17n93kcmEqIZwXQb/4Weggn4JYj8WSX1Aako+c51UeNP6i/wA4QxhWDw
Uty6C/U92A7qlPNm5/H/De3Qh8IZRjz256nLTK3zEUIm8hXvu4X22Uvo1LJVMhPO
VjhrPqZz5jWJskdXq3ItxEwHrevfjhgiJvyRA30aAkPCv/gsbd5SBtw0Lwj92Swg
KK1IDN35Jve9oZg8kX7Ctx+Ub5JUkqNgky+vR4D2NMLsIOE3QWYdKdgZIz5xFGhT
Am+tRccHafFWP2vgYKjN6o7psfqWR1Df/xck0PsQjf98TyRJoI5NgjDpdLeLGhEt
iGbYOiYR8gUe5NJAqPeShvGJFOkvD4c/3MPuGRDiwB1RqdlHwhqCVucdsLcDJyK4
k4OgWN1Zk/kuRJLUaJSYETDB2Buf7Hh+OfUlAYbt8WGqEYatipzTTwu15+2XQD4g
Rbl50VPdm/+OHYPTQ1m0wu8qzgAN8OjIWo0Q2eW0gtxqEWRmHbT6YY3U+E1q5U+E
SQ2GURZRvJYfG0Y9Qw1KS5kQ63BDUEJe4SsRwqir6tHugSIgHlYhMIpbjqRQGCuy
ZMr5fDwtGYVj/ElIsgfNf340H5ndBFzVvpkBboL5UK/pGiRBM1AiuP5gE2G6HZgg
hi4zvT+XmRSfMfAPxKtYb6JoWjrXdp5nyzTKAmoJb2PXYhTl7n1Ta8yr45xYKQfm
63fFyyhZBkk8gSosyCh1kxnauedtUzERbAQtP9NKqrCg+SlGFAIF2h1xW9GxFWel
rb94HCoeYKESEvyb3aCwoW7qdRkAVCAKQYWeTc2wpnChXzZbZeMi9NyRURaAiyKo
VxQQtmDM7kP5WydCMn5Xo9JUBQPnk3lUNk8MvnnAtIIQqVVZt3FvjCRiE8ab63/C
jrK//RewtIipY5RpyEEoIJOwZppKhfPBOt1OysOvLyKttFTc5F9D/C/sqtND9PIo
Ronl2QT2G7HnFGD+JBx/jhpGx3kwQvukIyKKKZ+pAHDTcDAuv03LNK56eM/WEFiz
NQKDLhJLrDug3SvR7lgorIbjYfg6DRq0zi3vYhoqGMwJqf/otv/DGIeh0hoRKuKU
shWV0dTv0Dm88gjezwMpNwVZpSqgpcu7Pnc1RUf7M4+A86QhEac4wj4Sdp2GBR6p
9TKyQZeCkuq2dXLragokr7Fdyc9qBDRqyx3Gay/ZhN9wgRaRfrzqQ29FQfqwlUy7
XfFNhktJAMGSQXPfGqtuvmt4ZeeN4naPZY72a5rW04UwfosyzaFAP0G0VKKfRvjp
KjNIg4mCgyegIyRZdXeYErZOQj1K2m+ZugxFhnE+K+39mjiKKViHl6MOEtfAqjPt
ND8zvuaLaPG2EMDhOKkerMw+GUbvfZ+Z613Nmx/SCrwMIUyG5s+W/oI987mmMpN5
eoqBEVZN+vg85UBh/ehOIKB266FKjQe4hRYTqT4vVjknJ5YUDWzOejQGKgRST3av
mVsrAjqt4+nq8aJGKDf3V1c8oIyQR+pOafCVRuHDVRQRcHXK/2ZOJRpOwaKpvTym
ogS5/x43tJWRUmph7s6yij1cS+wOXNVJVIOJOvTaaZYZcS8ueOCK1GvSV0QqDqu7
axc1ajePa3//rkCbGPBzKpiHpuUMZSvLIlBnt/5pn6HeMJrqjkM0iaHDAyOaXMkL
upEP7MDlf8sebMWKCDR+Iha7R9k296ChGIZEP5X1cL+j+7YkGqGEbLs+B7gqO7+G
rPeAqG8dwokGGj437XRvvZDpoQDYOjaApkAO/wRfMIxPqZloqVVJpXvl1y3WziVV
Bsi9c24tFzbY0lvEqz/rxHxWERtRWFZqK1OAgrdtnQbsgjbdurT08FZD4vyLfAF9
i5k5zmmnmO2eXG452uX0mjEfg7scIKUkCdw/cNPFQymEUEmh4wSF5ww/5qxuOcJx
DUWmC8noJZT967ykA18D8Xpb9pdX/DCdBW7MgmeZIwJY0dDWKfNLHWZY+CmEmekD
5FKc/+wGqRAMcoVXWlChg2BtSk9rWvdrkK+Qi+pJcpQMKM9siCFkk1Xi9NwXbMKM
YNgU43BM3QWedHTrb0hcb6pgL/d6mEpYhNDarK/8Csxxz1S+LDwiJJAcWf26iwuG
zJESrsXy5tRJxwsz6YsH/ly8UIEcYrbUgVktPUGCGbGtut40Ny+ocGYZqickHA/k
9j4wzvGGaYHCLPrwxNqveoVjXH2+PaP5dRrqb5SKF7Ie0vlxKy8SJtAh4JagEUE4
3DRebiaHpu1hZbs30drKWCC1GV5IoFpfsJpKIRTFU4xgmZbIcMsKPMXgaWEXFVcU
tH8gV62uMLXyhWT5bdH8b65OKgpXlGY6lMKnOntnGeJ4xizj9KunHyG0twYUFfWX
RsJJgafsOxMZohTzYqF9KS6GO1A+dP+wmiQqY7r2B0XeghCapmaVp/n+4B6iiXIa
gv0HgZnMdIU72Oe8LryoU8MjVc/C+f+cd/1avCXfXLqlAf75tjZhVRal0NJ7pz8y
OUNgHXDJpmSXUI/flAedtKUsn1VWQIbVnJLmBlKkXw1SrZNa7YhweILSrFNkYHOP
i8KgRXn85Qf30meyBv0K6Ip1f5HvyKRGp2PjwVM6+SR0ZpzKeZATeTrbdMsUOst4
m+MXWyYRQ75vVwyhhwVeJIcaxqxeRylHM02GL14xjU5Ka1tgBTW7AbTvDCtrkKg/
X/GJSvXFlvUy+iAJdzpdcnjRSJmTxKW3hYT1y70/SW1nJH75BQV4atE0cunosWb8
F1C8/sK+Iy/jTBZB6XHPfeDieO2nsInuxny6TYk60L+POfDgX9qjaHJi6mGoi9Kg
wQJtjm61TD/qwJ/ZIEMFZZYY1MIMZmAT5EEOUZwnfyCSdt7os+GTVQwE9xhCUtnt
81GjAXPvdE11KyWc9qLFcpSyYebnN33p3867WbytM+ggx6EiTnbOfrpQTZinTdFs
hNOeK8wCCQqE4Nlo3wM+jKqkV78KKFBGtpQmbIWS815qFykE93wbDQ2pvbz7Ukbh
YePUWDfr0cm5m2m/kuiAqpWW9F2br+S9IqdepJSScctxPmKffpEQSm0t/UajUP0W
WPoyHu+t0umKGS2H+btp+IsC8E9Zp3JvaICK8A8vUVYbjJc5En0k0Teo/lCEQ8At
VgY7pb7MCyMDodE6K4if67OB1E2HBhdHy5oPZNi5IVTAlT/xV7q0ZnSBgaaSzb9d
unxAIlSjOeidWyqcBS/ZP/TUPI3M1xs3zsnY4iS3r80iIjoA7vaB+BcUf9nbFwVC
vZbXEodQoSHMcCYzupKClD+f7mOwKyoaOqNVXbPPyoBOl0OniWw/Q36Zey77gxhQ
FejsRveMjWOk8aAdo0D1FOJEUfs6JXj2sReV6kLiOAXKzxJH6D6yb9xnZnq1HodV
3soxaKio7IRVtytbet+CCLK5pDyAnDLsPdPVclvYxkyJBBr+J2TjJXZdS6ljrfse
6nZEsDIZcnuRZfPHf9bZ0KIrVJtbT++F/co3lGuOnIz57hctLf0a4ofEqCUvI+PP
b7IdhA5ylNgnCNsQOmdfmRi1hu9/tXQpfgN9j5xgjP3emsch8suz1DFkP5C0W7Hm
v/MbbPz6+9S02kyRZg+Zia6jk83BebVvVuER1/9TONeWfQ1OIfF90PVzjDXd2/2F
0r/xOh3mNsgEX6/WLTr1X2EojFCU4psjY8pEQwXf/BraJUAucGnNjC0lSD7F7pIk
i1UIOObI9sLS2z/JPlE+V+N76lGHZ1qhBrgzWu9TM3hge64krsD/2VsHnkBeijz5
NVRMuACjoqif+12Fl7vc7j8vipjIXmrpAB18gQ7ybrMeVeyZewmdB8GxeMRt0fTU
kJMUBdCkOtmOlvRcpGOkjxFkB+Y6IqnFZD8+cSjT2QAFBJvMXce2J1/wxFdSVM/p
oIlzfi0gA5u16bG7TbJwe8xMbqWiFuf3/q6lT9xJI9JoobK+xqOj4tN3cpX9qrIC
5T6TsssK3W9FU7ndRhHHRrcSnvAY68F9RPSrDdIl1+0KOTALhF0qtzaIPNvGDWvw
IvGjWaw/aQ+KHQ9MZdA2g/ZffGmtk3I3qyub0SCXJlrYvoF7CU2se8Tu2ROqHe6/
I22iVOW5Pp5WL+OqVZfi76yd6prYaxsn48ll7AU4wI3yvi48Csti4ZtG+znj8OL7
W+uPEBcElKzFARkKYmoL2MWJ2MdiV8pVVN9vqDtDglpHPdb+DHcBQh5g7hjZWfca
LEh40FC/KYkLnjLApPp2Zv2sPqKGd5nrJdHRDOULMZsUNnQf+J+gpa34O7bKcThJ
6m08ngenTrqBcnrFRWMcXxhW5+/ofL4E0FuuWL186zcT5tuHzdKvhmoZ1OABJQ6d
sAlQkHAcn1uICBgRd7qDfDDPV/uoWFK5HJdMV4w1tCHYA3dj6Rrmgpxrn7aHMstt
R3m0GRbpblLHgUabv+k/dQROqml5VxGZZzrQDMT2gHLlx95rRlCh/Z/GNc1/zP4R
MetOpO+94G1PqyM/REbBFqvJsALku7Ks8m1N++TZQv5otw/OIe97wK6dG4hwo/Xr
6j8BgtULwtkjVyFxJFyGJ51xsbLRC5zEgGihBLLMmoj3UP2+KUIHSvLF0VwpscGk
RUuXZMTE/vWI7/TyCQdFXqdbN7cdRLsZJo2lAaiO61E3U/fnpVc70yUnTGGHsmab
NPT2yMhCGnNmUIzXzlKXwlnOsVJduvgFQZNXwVbiII2ZbGsJT6qESbKEkdzDYSOH
Fo2uZMj/a5WE1GdGPnGNeHikzDJ+c3PTz20o2VR6vQQiGBElzAjYFl0tMG3dHA20
6U1zEzT8zyo9xyGhmL/PMx8bqwUhor/AZ9QkNPvXDsCJgcHUWXzw3I7UsChtsn1g
rQyms3b22O9DjAAcRQJe91RH9ISBOu7IWB8ORDsNltM9YQLXiTi25QB+ax75TOP9
+8PH9j8/T4WFzG/YIhA6QN6YS5hKNjdmZd0E999iZ/O2wDbPDaSpSO0MzwqI0iU6
SwHOtbVSet5h9tP5Qq64QKfqrLc5LlJujygyoBRS2QZVLq5EAHYIJ+OBE79n55YQ
a7NIS9a1xmtcqvnScdT29Qu0WxiR90wwGLl0p4g8jgBae7SCdshqOWEFUb11mL8K
Mi2siw7fIoA7hCqwhz0SYOimAGaVC9dtale1ZSPFgbh703sVItP7GcusVcY8spB0
Z7k/SC7pX9rOTvWg2BWJJbsng200J4IhVARkTFuKs6TBXwUf61bkcNUBP1JAWdAw
UQpmZXD/tAtWGVfNCtqaneopG//PAaW5W38DrZ/UkXtQcdV7oYIE8Y5yhXNuHsds
sCQFSPKdrfi/IMqssAsrECYJb5fnyUlQipnhhFiyulPwbv18RzVm2eE4+uom8WZG
ZOc+RkuicRnELjZ0E5IHAaK0TayDpq+zkPD/4s1LkzrbvSiQCK/lefOeIHVPrWOd
Yjd0zCUtwRIZz1T85mvUsFe3HuquyWq5IPI2JkQ1f8rqFfuJlYXs+jrQDtYkAiMB
bsxUCSCxkfYfoH8xn7ykTI7ly6lWH8CHQMfhF/eFd/19F+3pW8jH2A5Im0/LdW0n
st35GJiNjAknjhob2p2epycJaGYhSOzMmQTWuKzpNd8GZyOvZlLWoJymMAIijf9a
FrUI0Z/gM+gE9aTBh5jxAVITyLoknkq9FxQndJtg0STjg6FUBZ5dQVwXDScQ+Zl9
KpCR/uT5Pnpe+5W0JFJfBsLoiLl3XjBwCQkB8A8+wNi8GOmmHBOgtsIhHsBMMj4R
aVBj1MLp19v7cR6AjHXcvqIxK+ZhQCX9vwLfc0VAnVNKlSSol8tduwkRv+gmnLoG
w9sKDQLMdB8mFXcLW0Zgnx2WmrhX7GkilPYjWOSERt3gP8vAKcMzhm6KmmbAQPbQ
TTVZ7Zc4rnXTW0thcvevM1jdmnOy8KN2u9lv9PpmmfX/Vs7QNRRjv3gDEVJUtEru
LotqPYZKdoXhNpYasdIU2DeWJYMdWdM9fgNZynvKdcKfFN17elTkOavdyM1vI9K3
IpXnnb4moEYODUO6yko6fjGBFKJU99dKQPysfASLLlee+LeyBxe/0Z+WlmpaQykM
PLYvpBQfxkeqrO+AweIIqKHHI3VBB8vp+fCr5wClIU4xcnRU5zZcKDvv5yLO2np/
6CGYFxm89b1h7Y0mtwpMgChPNCs70bNw6YffHMiGr3k+5WkagYPom7E4S2d/yRFz
DIikrN2P85UAXiczwWIyBCpziL6le8cJ2dT6KCzikLlfnWA2Hvnh/mm5n5xdGXh5
SPV93rFODuq3Do7ES52mvNKG4Xj/lwhvU+DwIUPC1YDO7Wz4caTgmnuNRCpLsfib
tMhd5ESz6/VRqMaDHSEXk5oIsx1LymsRMoEOIJCpr4hAivZ3uJdRf1y/HVtZPj9+
nZGUXDhsDHP1lZUiIj8o+TIBTAF7ixjUt+8/mOkqFGMyM+T3555KLaq6FEr4al7k
kBvKZD62izvHmWDl+7fwyxFGPAxH2RhsWXmb/tvybNUqLLzrNY1pflbE2cYBqrk8
kfLqY8YpmslxogWfNAQrhdNMQtlAt2K9kTVYR0hmn42djsNQMFRCl8SKyhA30hEb
imI7uFS6eXztmVyAtVP0ravc4irFnziojbhwOE0LGn9ZQYfKqAHVDoKQSKYETETE
6suJdp0WCdZzgPLn8OhB0RZqVppCWdMDdrT2yrfGEsDoosrarKyAQjsLwEHwJqTv
jJPV++MSAGzeZTKwuNNnatjcMDkhImEiyT1hH7f071rGmIoQ6p8n69vT3U19bBbf
b6SD+CbQR1L8lzfVkONWUHYJksYKfKy3xSuSzJsEqsr1T4AGws/6IqZTcf8jzg0f
ZbAdYYDfqJll0A6z8bQix/c/+TiNeCg4ZffXhXmtOe/Wp+0lycdeDwJ7/7dPo800
7JlSvnpqB36KWztB+oJOVxHOBypgeaw7d4gvExohw4A86uZz0gUQl7iLuYAX0yHM
CiHhaqiAwahPjOIE/il4BZoABmUMc1gLaaeGIsbX3nVT6N9gAIwD50IfRkG4cYsY
dFzAI0doqLakhjISmDCGE7wlY+0jens8Gf1YPcc1LCta4c8pc2Kan1IT8OuMgVSF
jNfvkNvKNqopMkq4RKWcDKk9wVcK2LebzZfUtkz+GVodA3sVHgVTyaOZBpaflD81
hz6coqBrj/ejRg+/jHgjxWapOXHtXqYyAcxK1aTVGYbDWee9TLaMPS9ZbUbOf/Ug
0JsIU9d/XpvncY5QyMNtvqaFYxuFtNjZQc4d1woxLm1BBmUQkJvyArwjgj4h1JQn
yXPkS3Od3KcyhqbDLxPCSkcMkFElwF/IZOTqXndPiw0cjToTcqvqoqTZvccyUblP
8JqWo8ttH8fmyYf6kPgrO8O2Prhhkkt3NxBJ9Q7684KJX422r2+4fjLFVRrcHsqw
Emkn3U0l7yXkHEqz+sdXX6Ik+WJP+OVDzZ36zP/sOGGVi3/CX+nfyTmFKQsMwOQ0
XHDbmyz/1XugW66dIbrwzrG712GmcgY3gOogvZ9w9nw/aPbxEZZa/yQoU9wm9xb7
p8gkEnMDre0Zs5ZQKNw3Za1x3I0Sp/pOWD9esgGzsvTrQ96iJQmOkGJUuR70mFGD
idbHfN9abo/K8DRYNcwSuFWJ1hZM0Nl8O9+L4ijsBRrQsOBrAA9qgNvT47gCo6rD
WxajVJJwxlj7KSy/3LjegnFGcLcyMeBipmoCybgIwT94eVRrlIDBkCAHFTQquZ8S
yXRY3NzaOK17P7XQbEFJ/AvVp50AzMkZsvGd3fuY6xF+fBJOn9xtDJd5Y+u9okvl
X0UOiUyUcIMxwgxD5JJ98KBtGni0kHn7MfxCZMeP3wpvXul6/9EUdBsR6kD/dCUP
FRGexWzA1xzJcLz9J2x0pWFGNrkd56JD5KZUON34vr/gRJWD1lHVWYIyeyzRJb3e
E4kVODWgtlEyrBMt3j1xn5tHJXIrAwfTQqn8LYjpboHuucRt2AIl87YqMpFhrg3u
V/Ev/toCaFlZj+NUxLJtGr1p3FXHPXBhkBi3tUbom+Jt1VNrb5AxGJPWMDhVrKDT
d0iGWNs7yseyV5szvIHDHCNoIJ+r13wYZ6qRhJLBff48iQFryJf0A7lRHCl5a2a7
Ab8AD1V7sNN8ufW08DEytzeROpdBJN14VBD8iw7WFFzv7VGyM1etcdOt3LPNoBxS
6Cg993JSrDsv22DqSZOKM2wskfksqI22tJ7TKo5gsoDietqRdpiyeOTAweLN5sJ+
2UdSYIggCEB3ugfcHm2p9tN0KJZyCzTZ2bQJminThpeZwy2DBSnhPXeI2urQrg/p
r74e9mDXxqJb/IuSYm2awAkdK3rg/1Y9XyhreX6eMJ7wTKW0dVDjBsoHCkdz7X2s
QhiuOuI9s0NVTPdZMqI40KfvKrLfLa1Mwx7/Ak3t8Dsfy0dy4keHPiSowKjqR8Ie
IkGJFn6PefxjQ1Sw4MjC3jAg1QOdyHfYbEgZmWxgoSgf1qNYE7/ojtEHmsyzSvsa
MUrbKaCMXXssxfSdaiFydAMKK1OAgQR3mBu7PvCjUDqauoq64fKYO8CxYi9gthL3
ux+fUxGpo8Ay4zL5o3IMKt8t3RATNdtzvKkAuaGa+kzFiaYpswdmYp8Y2fqVsFt4
WTlXxuatfmqc8fjh7TWVDVs2O/O6i5eZSwRdTPZvATPNSan3dx65K6Bd3l/Lvy6+
OHpMcKc6zgYKhBSVA2e5hl7wa/tvm2marEzK8M3TYBv6KvVqLdNlkH69JUq1x+e9
NWa8owYUtLZtWM6I78G9KmbNwBLz92zD75Gp+Nf2Za0WVIYOKEKuJd8f0EdnBxiR
fNbnHvO2w8BpMNfp4pOnKBqtyO8Y7oprXCG5CHVU/HsWYA3UU67+r6FAWdAijHb1
7D9qNiy5kFE7U7XkSz9yR9XxWgw0w7E+a4W7GzbtoWUyYVoAA6CtgUEbqbyv0uvB
+s0KBazQqyi5SyXSfARsqYkU6WaCJ5BdGRdT2PjhZyPoUKTPiTO8nbpL5y2SmOAx
iKz9DxMGEytyPqLMQiXZuX2ujJFWy4DhZodi+kaog58ryVF5UXWI15gN7dbHALQ3
eHbQrBSeXTHMdMPk5nt0iciknZyzbO2LJylnAw7R3IRvvUGCzWbR8jbAh+5DUXfR
qqJu89wfAHXIdY1+uWsazv2WtBOkSCUBSp7AVwA16BJLGaRmSzK5mf0rLqClt2KV
KjluKlCuTmHzCBCukuvoTtrdGum6re1dw1II+IFTkzLAmqw25dWpLUeNi5JBvxIk
26rcYdkrsWyCM4PGxoofX0GUCPvNYfihQF6LVbwH+l29SHVtRh6VuDRC1OOZZEGC
FSROhLdQyNerFecj84afGo2Zs/Vejl52z284++Bye8f0PcaQ5nCGvFpFQaZB5CvU
4iGqSdhJvz3zif+ZJEz2VL2VIUjI2OOy8KIO9IYlWyFDIGEYcsfdhqpzsKwx7dko
5lyUD18UdZE7DsnabRp1rnDf7y3ufo+Pv38xQYlpCdujO7npuoq2EKKRpYXm3jWp
y67kEFGnU6oG5WW4rb2BhrVDoCbCl/zIxZ77k18U3gPrkLg9TVAxxWkKX+jykiC1
o5ybjKaYKzAfxZno3Hmax62XiTKdnBPG63XwlTAczldDrfBOLc6phVf2usiPloIG
ZOLGE1SDLtFFpvzmc06SCWh/rXNZ5JPiWSOnHIl46ZX44MHadgT6o56w6MgN6C7t
UEhyxvuwyZtEZH9R6mg7xO8VMn9eNY2dk1J9JfmJYtedn3SW9sSYkOIidqC4Vj7+
kGuuXi7ix5Y7uHvisrWM88NtPT+pIefpIbeWP7uy2C5nykRyK/SnjBrjXgdYY1qS
3S36r32B2nBLZfSy+QZAPDqNRcAuy6KkfSRsMte25gNrYUfRL4RiPvhiyNMOfzS8
nFEGzL6sklPwQXnqMxHMDIXazYg+1zRClAXt0KgvBLOawbyhLODqgqZ3+LVVClQH
selXk2+lKvt3s35ZiODlPY9jy9dEDr8DikoNRcT30YBdH98zDeKrIq65RfQVmxnT
7uePJLTUO8VK0VC4aT+hAoknDHxBawGEZOuEzYuLn54nIP2604np0ZdgDu2KDrms
KMpciz07Mszw2/r0Cq63csGWBli4Su3COM54u1LORaPKHBcH2IdqJrQcL5RtFb3N
g0HAKVXznVOo6ALfB9rw6zZJkSWbtQaq/tNFkukKg9DSuQO2EXNFRWECOHTwujXV
83uXvyB5nTUZUA8RpWw77nR2+YljfDjt9yPvQL0DLNnigAXbkjfW77Kf5B+hCAQT
PstRZqUdJLqG9TvjjS9bJteG60xKRIpz8YQt/bbJvgJBK0LRG4Uy3uUglje/B2i0
P6Kerfi4QjcHNi+1OvBNNMisO1g1KlQsN+uI1/iWhBbrdWq4oIq/z6hIkHim7yg4
QyAfOg0PjTrmBRTHIweHseNh3Gx62cM5mZ8NH33kYbZBSX8nDhUlmEO8RMRE1y/8
cQwujuZg1czDI+CzoeRFrn/Qsp+IKssnkZnBWAOtAtkL/OCHF+ULRPLCSdNahRV9
v7rcsvfrV+xDlfSRPEQXwGXnPbXasIg6Q/RB2UfoAB4MK1R5YwuLvJQBdAJpGpge
nIeuTg+sOwgmCbNNHe4vvchlKMyzdVWj0bHMGW/n+6xl2QE599SkPzbhmNokrr+0
iFZlbDv4YbO3WNFOjGDPfTJ//yNntIbg2zvJEv5AZ1JcEKFMDDrZlIXvS/7IcVQR
/F8rIvDbTspYJ8CR+UP/QkVlKapqwdXiCn0NJHIi+SdUzCTpx40wHXIWWdSgdQfp
kFKlxmUDBheJ/RyjW+LY+lpKOqv5C4M9Rdn40342nwJo9aBvGENAWBeSw8Ex1DAH
2BTa5pnm26RRNNq+fFwnD7TBNOq9OwVeIv8y7QhmyaECgrz7rGUs9J8bsu1Hvc5+
I1UpVwAt2CkUxMMQxzPCpfsGqJ2u3iEYDvxpCyH4TtVOs7hUvyYoECKvTvOkRiT2
ECjkkqHaZRtYqFv+f70Kzs3XucIqFpcYErValydSdF6w0V9b7+41EwWR3grzuDm8
uWm81IWYKmqqijZDHsgx0+otfeDSW0QlsFQqyTOLb1v05IxBc0g5qV3AWPD2b0Vu
XTKL7qdGmCAtGC9Pbfmp+fl7tRKPfX+fF6cXnXKmnk7U4N7FB1vxjvFOI7r79vvj
/r0eL1HkFHtNYUKU4kE1gTV4rVVPgtnd1vE+nPS5LV8N1ZSM49PmwnKPi+U3zUYZ
z4i99DDDciCQsVaEJkhUQoOnj2rzol1/QTwyWnIS074/qQptFFSOcJ03O/YjPsRS
DsxDh8jY5Su64jUERWZPHuGj0xG83yNzIZwEi7tj+Dg9l0dMQ8DLsCOh3jwCe4di
/uMuIw2OOrds7u18bOwkG+buXwq5MMnzM+iKYi2B8mMm3YaBwwwltE+ERTJrZiAu
hV7befalRYEiFhKxBgba3/GS1I4XcFnMn6xgvDJGvyIyzoK6kEY385ME7R2H98Ru
OGPOgUUiW7WmLX+KXTsUogaznHZ46omqeBwRyXlHMMVUu6J2tNz3WwY/jfdunL/A
HGKKBhKs5BeevWYDKbrS9sUm9QNGpLFfWU9eCY50dJuIN3mWLqywLA4Rty0UGwVv
XlqxoJ8nqs9DUo2SwZP2V71C9O3PzUQTzBe5EvS0D0u/lo6aTzS3TV0Tj5+xYAVj
dnAE5x4ITZidvnrrOa66LWN6/NvS8WXndEn1JblumWDqmwz9qcxr7Wrl8FfQoUGt
N+fpqNOX6KJu2I4QllYlUjJ3YMyCl2VnxPX//9JFPMKcBi4OMBsrsjiBnfZ2xybH
a01vIGb7vPGVkHcZV59tFSTlbNAz5hcBEoMyso1Xb4U2Zb7k46I1oBNT7UMMihUH
c/WxYQlq7H80OdtHJeiTrsrQbhLyLpFskmKfOpDy52u1mP6YWPnjFajtXybft4A2
zw89ifv03yc5mCdokfPtm0BIDnqqZ7bRELezGQw3hJj57/u0cC2db52ycmO/Ji27
IenAGJv3JTzgCLgTJI/WLhJaxIJZvwJimMvf5OluJJ8NlVWV4FLQlERrdwM9B0Qt
5n0nfAAdZNI44WenZapEsjmssnI9vKCN4o6jS4esqYFwQLNDUm4/u/x4jz+MFIDW
iiDdY2N+kkJTFdOz0JNzs8EvGhwsvIrXT9Apd1mTk+Uw08x8lmja9O4XQalN7hcL
X+4wwBsR10bKsx1Ddwhj2R4Dz7aX315PzDN8oglH+KKgGgLyiqzOq/yl+U9hjeCO
ONycptqsnEvIWKHsYOTVcs5UyTNMNUvAbh6gLx0xaefoDeNdACrG9/t3eYBZDK5K
yDI5PC6jMM+3tzMSvjCRNT0e0dkKuYqTvyk232VSgHd3UTsR9rnAhBXgQ3VbVib/
KV30EFL6ylMXAu0KbMABzhMvOWdL/Uz/jp+D0fmXU7JtpkmciTbpxWdjtfs6wFN+
uKarhVhysDh1mLeCCSN1m4rbhDlo0NG370YOP/O9BGfQWhnS2OUMSdll1imHSMHT
PYxV5PZ7yMdFwRJVzPi/7vvpuOYp+2DJHDdXYXd6IEPADrR+rzlTLA4Vo81t6gPE
PCw3vRpApeU3zIaFyUPF7y6Tq0qecqpUZl6FRBfjsENGsZIsZwM+T2yKL6KaTkzo
84GcnuuieJW3kUelPzkVCovNGMpGpb0M9LFsbQ6wAfNv+FTh4iS/oBqTZbbEKIPB
tmZKpc0NlzY2to/lPfC1lTZSweJkIOn14sM/YwlJeBtQkYQcALgq498gCwgUpByC
JXXF0xkGmb19K8+JjWifBGbvUGeedDHOmm4bcaPoTyLKBpsAnRcygWQrw26jYN9M
vQcFhxvCFqDY0fvNI5/5fQiOA3BVK2EuiBYnBy7M+yfdfKQ1UR/XmxBE1WcRmP6h
f+YwqE2fJI/vtoY8fH4b2OiiI8xg7jzDeU3z6AxewkaJ+JqSqZ1pBEZHaNtfvhJo
Q7w5SUGsqyRooaC0EWsXOuxybJoagouWgS4SJuVk+JtQAClewowY9UlYKu0wKVle
9yAdlhNClnmSTZGOAyVVmX50NTH5imnGj9wn2AGNMU8vGZve5AehGOgZ7adOwSsc
9U9NPpHWAJ8OnTbiZKXp8YiWdOAQPqxpbx/5SBFklCg7zuDs6mEOrijxSSWJN6gz
YFpwsj0sM76B/pNAeFARkbZAmU2SznPN0pjxDDxie3W7ISi8IkZIzbCAJUBQ2cLH
QGB9BM9aoPtEBblEYDE9EWrCS2musBdPENwOSm7G0qw8pmAzYFoCvIZM0HxcdjoP
eeE8rmmVgcdllBXsrk5gi7gykoTCJRvJtxNak1/7mRwNZYiGCdzt28eaO5T7eUYk
MnZF3sMydv26Ftr33UJXTDeG2XTRf0IStNKFcwL2//Nn7+FFk48Cd4GQ87jRazID
1hD7b321/SPuRiFjmMLHKVBHJWdLrDs718rQgkXBYMJ4Pt2jSJB4c3SmZycU+yeE
Ad1OyH1Q1CKtkuVwQbu4nDxbs9kJeY2GkQ6W5WIkOEMumhSi/2p4MxZkO8Ah7avt
OloqM2eI7UQGE8t+y5qrpTpkctRX1Q5mdfDvMQaaWDIqPoWssPMjMMcuK7tjCm/u
6P8FrkAPzadV0e/+vmjeeVPbFD5AuXtb9HeA/Mysj+5Jhp0btTQ++XEMV5Vnpmha
w4HqY2gRPlH5AVSaokV8eUzUonsn9cM6jH8UdxlrUIseeDmN2XLiy5g04XJBDU7d
cS0lVDdotpIvQJDZaBV8upVjru7ifZghlixhQIAv5VBI5L116cDc5Oj9Nv1UvpYK
sqnOsJFXrU1Nt+Dtp1xdJk96AQtj8ZkRAgiNOM0CMvjWa5JGhiRyzpIsEHG/Ki1u
wAz8OeZtY3j3LtsFwz6Bo9JzUUoG2IxfG/YbPMyqgZ/NuXu2/mJjjE1OPaN85oyt
XMernCR4QAYsba/I4oi/Kn8kwRRhOnwv/52+gjuG89s0BEqjmizdiMkZ9Wb8Ji8K
V0KlvWFnyfqZe2Imryn9AKKbL5qr3bFVKMi9gcOuXkBCVqS9LTT3dJ2QySoWi7+t
biLjHXMPEOryfaRfF7UEEtXhpeD5AcP2zsMWypKIH41gY3m4T/6QzfMden+Bs2vZ
en79hlghUDKoPijBFt/kUF6n6qi3M+ryz7SqoVpNip193BuR5CuJ5qbRdotaLRHX
3KHSgmCb1UPL7VnIL78wDXihs/owCeqM+fA7O4NgB+WlUybia40d0o5octviUGyc
5OHIij94A73BvBg4rkZdjRESUuD1GNvQvoi7bAGDZ3wXFdIoAnaIME9+bWfG7/gS
C108eqI7/i8dRAsETUiDC0OnPci6yomJvcVKqXpJ1oKVom/SgSIVUfRDPlfjMaVn
oS3XKyLw7eIUPzvmM0+xQOthK9/2GAsv9ATDfp2PJVTlQWjNfHDmakwH+H8bAZoT
kH5n4d+IQ2C5efk20qukHgh/1bblDCD4hzVy2Ynk4G/k+lZJEIPxDOj7WHSSIeBk
AR/s7kpH4N8Kc2HspKVT9D6J6qk5/l6UF/WKPXQwewq9YIR1i4di7OTtiMbyXBex
0v9eYBqNNheJa5MJtiHKr3ZNCYt73epcwV1CN+2Wv/d5qJZFEHF8N8Ui+ScuJMtC
pdlrq+pOAOqiOEYmF1TvSefz65PCxjMLw6Q9kSYXuN3JSLcEwUVg+8MW6FrVYOom
vd3LNvQ/jhA8LYACWj1u/t3ByLyX4I4RxHUOOvW9MbdT9TC4tWbrqb6KQLQMUbCR
aLd9mxCgx9oZKMplGOJnmTtay4rfy05sSfM3B30eicyVvlcLXp9Y+FGwLk2992mT
WVrsfCUm4Z9FNP8ny3veg97PZBhZj7OZSse+i06i4Aj4Hr393rNmJjCEvRiweyfE
UgcTBZNGy+9eP7ejsszYkhF2/+DZ3GytykeAI+DRJCr1mFF2xrZ6kZbZBFUHPk26
ZVJHQTb/GhpdP8NH4MK9igNNIP3LXUxayWIUn5vgRKPjNzNs6TCIawNL5kPNXdkj
0Tv0b/kqTLHefEcfCNko1lN7ebzzxYaeIj+GimT46/pmp9Ukkq9UnJQNOg8jErdw
6JqBJX/FmFgjaigrg+CMamyXbcJUH5uqIy1eRSfEObgN2uV9KNZO1vrggJ/IE/CG
s+XKDIlHf/Yu8dDWeTn1Mvr2h7cHQK5Hjd4bdytdelbg7px9G9PyKRD/zG+Kls1k
wXEv8MG3I/vzNYOSiy/RusUOd2CL+YJiHMJHsYgekkHeIqQdQhvpHWH0IbS3n5OE
pwZcaHWDrY/qO6vjVklHejpMpFxBRwHgFwQe1+exUcfts6b/oDbBeKzd96HaQjpe
pkJ4or71OSZkIfxGnm3drXv+K7fKYlHkcSICQDx23J/Ac1Rb9QFUY+Q2DvbisPeO
qlJN1Cot6lPvx3sdy6Q/WTejbqrh7/MOM9UX+2wtSCB6rro4NC1YwInVplye3NNJ
qBNkqkuPrVDbivdGJ2+LPHxEhJAyeAve/eN7mEw++gnAr1WUPEduoRA8wDy4K30D
70JlgRhALppG9TPHoizezhZtRgHw4/Z5iiby8EInh3zXkYPSzrOSttD6/OKs53mZ
AGZntj3sFyCjwuFNW7VX/VVRhOm6vQeAs5KBorgI7L2bq9vJQSNKAurOYoyQ28rQ
+c5nRpK/f9KfYqHTfrJdVX3zL03XhovcAQN2ApPRY2fHsypQHgRS/5YWVIMnu8tu
tLHhNY6593OfezhWtfsB+sPzVbcJFb5xxRBPCz2Tbc4JW1xzFCfL8IV1FB8Z/OBl
cWyDYqBw7LCIK7S6/XX0yGqKO6UqVNvz8TEFTmXqG4h6feYrl+v3Aiat5rTY3MmK
ZxvjZbKG2M9LR7eucTzjXYqgFygVFv9NAnYJoXiuMH8oOp7WtytrIRNg0ZPQCvDM
r6Fsas8udevWFmBtreAKtirjs+VaHQzPhM5DOLJvowGbnEG1jANRl6f04J4Qbbhc
B6DJFy3ksm+KZ6XMhE/UO4vmkO8aiMcMaEgkCi3EWYIR7pdyNuMef5gd0bS6Rm9F
1tM27tKicBFbBHhoOTH+tRUcejbtJs86Cj6sAa6wfM/lpDgIQ4+qoKV31nSVQMkc
2ocbJlo/rFyHOWYL3dIcNmjhNmnAeb90Hf7hrN0lkX70Fb36HoOP9zjgdxK14I2s
HCHNABziWgMc/B1VzpC1U3nVfnxU9qX9nmRnHoXIpqjg6JbBwvtB8FsR0ESwm0Be
4tVUgUtyPLjo8+fzOTPrVLNoQznOtQ58t02cYBMCRX5b8+uIhcW+VQEvyWqHwz9p
AgdyfatUT15R7CiHC+WTHvBH+dpwwNsfawJW8XTgrrMRDiMwW7W2+aro6pkBQpFZ
h1J4zWA8a+5e/fCIJvJnwikLhjGEwP8XuY7v4klyFCh53aDu5p3Qx/WpMbDsvWHu
92dLZcYQtCrZsmLf/KgALnD2dfLyQlZSWIkX0JzBopHJVqr+ZPSDRhRsJxsq5/Io
x4uT8B8K0ryo2PcAtmQc9MTBanYqtqc45KAe/mR/GgWNsMHg+1jb/11gfNqafMbz
YQPvLgAhUsmPf0Rn+wbCKmetR0mCItRrzFXIZdOtn6rm+02liFESSq3fnNvL2i8w
0dQRiw65sUqcyPhnTOsGuIhAaO0VNnIBYgh0yMGpN7TlxNiorWQqtgwiqrn6oDTq
CaPpsx+7HpBonHsoGOa6rrTEbfF7/O0Br4HmRGDRIiY4KDcB/vBpLYE2O/WA+h/A
jTJ0jlM5sNWIk7kv4Y19zjvb2jVdSYYHx1qhCIz2vFLMZVfYIT58Ou/1bCBWNOuU
EXFcCSSrohFnB64lvURtkRAjYzWHMsv8Sk8580M+uKjemISBYBdbuquYRVvcFp2p
MzSdc98Mh6JywpyfTE9TfUViq4IkoLssL+k/8UQIe3KF+QL0SQmOKVI/zFDlW47e
qbimVtodN7rv4m0zEKQbp+lI/isOhQCdFLCsApj9+I54ApblizaU/5y1aEOI6UNq
C9sxpofM0eW6ojHG+u8ecQllDYxk+SWKiK+eaeda8R0UQiI7RvQ7GfeEAXaIJrMy
W/pVHMG4Cpc5WVByhwbLd7N0Nd04+DvqF+lNYbUnckfeJwllQSPM7y5ZSzNZmYOT
A1+ZxpR/QP+c4B3RoTo1NauLj22L2/8iAkj7czx/Ix43dPWRMglS94piBI+1OXuV
w1pxXNQDwbV5xOx6UKClyVXgGpsnkSD9k+jL9ZlvBWd5JLroiChqY8PpqBtC/Lfe
esjep1BFohI9/EnG3h0oDyF7Z4dbmWKqxZTpR14JoM+82m8YB8gxd2FXw5aLFb1j
JBWRiXalKR3kNSU5E4fRKRRithObTF10T1PpFnPlrLKtFnXLG+dHFOqVEg8XNjHF
9RM+CdMxbkO+SpIyUcNLu/pPzk3Sv5DPJDTHjjdGTB3QYOdMQakjZxUz+puO12VW
GnwHjpnq4Jo56vGpzAGYMgkTFUYjqKP8rLOz/V3xvw6l8Yf4vqfee1BWoi6iJVz1
dNeeRjRTgANmNxjAoqZdg7/LWK3SFVQpCBS2mTfPdIBwoG+qdDFFkAccpiJh1gaB
RF/Lw4GKgIRhvD0R0dBHjIVXLwQyCyNGyClsqIx02w0chE//dgb1q11tMljhsQs8
63O0mlDsFGXe5sNzINxxLj2SK7wUevIlFqJgf6pr841sKWqnwg1RRkQX+0Kbl8mc
aMPKpc8poEIiNTsS8mXolu5xVE9obKxonPUoMM9zlGQMSlkmPArysTyiwt9m7zyM
HzIdFvIGm8OnKObL9m79i85wVMcIA8fueDGnH+MlSmjiYFSCpNMIkcQIVO6asaV3
SSzk8888OBF6t+z+qm7GN2kHrC7XkPsy7CP6u0AJSFTlIJRld6bIBySL5gaN8LTg
hMTgMoNynI3e1lR8J/QPy6WEBgoP54D4xWxTvRu6Rz8zeNpqbStS550r+KJ1fTBf
F+YmeV1TWsEvh+ZM5SE7JUsiYmXQCTjNNwHJHMHhP1n1CUEkw9WowXn4yppC6r86
+0Vzk9H6xvPgV9KZWdS/d5bY8lGfHEvLgbCQHU1swLpDHXiXnOAe7v5C8trEXFsr
PYbu/C0TzWLoETL/27eqwCpCBMMDM4CvPy4lSuPkz9KyraqK9fmCwn0OujIKaLHj
PakCiWOtvLUVi/tMNDJqdAlmOebfNbxjCjXZX50TZolCjbY+C6TQ2xg6mgF1JQz3
fr2Cp94IIvWP4hmSNjHZ516rLakJtL/YAPVThlSUHTRlxu3ZE9O2UKzsPbtiRN/7
Scsck0znv8wo/xH8cpytStRxb0GmDWbn3gfSwso96JIyrBz41w8vewogXMp055+t
mCLY0nTsmddsRL62tKX3OXWJNvXx7Afv8nkgDym40D4Jz/i8IbjcsjzmKyEzpAaU
3trPqSwf1IlVqYW919c+r+ylWceyd7G6OjlH7s75vferF9EPCBHosQmX+vL84h/T
saG3nMoUBtd42ubMGC+8MLGG9e2KGtZct48TC1GWr4uvqxoIBUWtWGE486vcxMVq
hGlBY6+E9bq6XZDET4zdvDq8e90eJ4ymXXoyLF63iBWL5YO9cJEXQNcCsAJlfBn0
ljF8G3jLJ8rvTTW9zqsiJcrxLUSQ1lVGliVYStl0+81UYuQD7kRepuW0s/yEyZ1R
C1H08TtnXQy5yW/ZkPiEdJOP4p8O/5PZ5Jw/dV4DbH2XjckIz1QD/bHKK0RiHOBL
IMeEXFzZDdKIfewvuCrFbZDUHENrVKO9QN1MJzEPefRTCscSjPdeCwTBIDwiq3xj
sDNvEE9a5X603ORdffYx9h4SkOjcbJ3F3XJFhK7xV6WRM7nf/FbO7x0BO5AxMgZe
PqUbKauIX4/qUIKicIQgieYBi5+c+F4s0VUtw6YHn650BgsQMrq0GLFOedVpghBi
UoN96YI2UaD7r2YHLv7pfb3rs1gKXO+jB32qeTfGwtjtne/YD/qBmI0lNzboSILr
Hi29bxzdxAIjEk/YtXXayXUg9fgi6kPIhuRwk4UAhv7nldv7KJrQ6og/9/sSfUd4
tqOH4Nqyb/NtFMS1sHXh3ZLVkpUlM3OiDu3NiN/XlaDkqhtBzyVhuyq81TW0IiGZ
7xZ5gxJ4K9wd0UyL6zkls18sRAxHJjyFupDcG2Xfdd7yiX5oCThKOtyaNq8mDb1W
bJ+itG75XWcH4CQjAaBjr9MGttFJr/qwNjBezuL/demzKUkPIVpKZeqXCoYAObzx
hUJ0yUb3sH1mU1JCQTEjgej7DXHsDP7Tu+jHTFw7n67LUMES2/VbVfjVBpv8sgVK
3HVaokwYb21r9649AzrPoogYT9BSwQdV5OptYFzP17LfiCNalVBArIk6uMZ2iQxG
46JmriuDNxyemmzlL6yA3tbbv2S/0WRyJqnRwmh1r97f6pEyRbrjwyoTv1QnBQJs
jJj0GRejNuhW8uKIk9wW5hUsxvxWWUjMEVbKnIjjdAJ4U0KZMvk3cEubZACjsVKL
xE/Yad8Qptr9qwzwj4G1cdXJIOtNkNud7P+ZxD6ovrzW7R1/oemOH6gckWkviogH
grp2kj3wBT6/iv6m2D93mk9JdzaViaCJQgocWIkdpFC5sp81dp8xFcOlbS5kAIyi
16/Fj12GKmP0uoZbrCgp7izJmEtCeWS0WtoYS142+eFDqlg0ZNK1XJvMgvbUC4Wl
/rECTvaoFjE1rqtHBY4repVZVxL2rAT66KpTbXlvUOZdkmlwnfzUUFbJM0cuncBl
umOWNiAVBTK9eKvfgi7dvRQ9AdtpDw2oKxKz/u+V4httQTCwJoUaH8+wzzVN0WMx
SMgBY4zWfx25+imiFOu/OUsUYgr7o7HPvz9qJVBNAe+pzbF69qOkm5N5npfK3XAB
QpgkHcyHZHFdK/vxEzNxJ0VyULuX1oYjv03zPFG/lpTsm8HTbmQUudB8vRUEsD10
1/Fpmu7BbBGtg2m71mxad/aUnUeZNLO7RA9JM36wfwva8VXH4gvPNq09C7oLWYLy
NPeA0wljciur/OLFBOoRzgT36esrXX97SqYbXIVnxmyTT/ogftMY+xoSW9AJNOBe
G88IH6lpscdk+kaaFWayLf8yOGKMayrTF+47VyAMRVpBxo8yA4v5Zh+tvaVdMbLR
NSuC7yjCtpvn4bSYsNlbpGBZT+gprNmz6ykYeq6KhTB7qdDygRo6MBdo+xWLM1hb
SQZATh/HfJjXqJaD2VYjilHygFBGKaGPAUfmI3SlU2zwFrzJqUBSlJ+WGyhCM+HD
O5yhzCEFC143i2X4s5l1c91c2z9d5oGrykA+lylAsAF2Wh7T0OrGFR/7QYmL74SW
ckg/XCHWhdenSPaiW+jF5b+DidDikZI3Dhh8W4Vo9RCFPlsVXv1txFsSRAHRx/0I
Ui9cmlf+4dauhDriGleryMOdu7LbKpk7o15+5Rg4ysPaea7LPYtKlMjFeuBDr4gS
RZYid+mjWOfwLjp6qCbb2/ViJKu4anjvKZGYM2KshQiBiu6RfwMM4hfFTqyYgLqf
ylpwjP8t8ZsxJVjXnSqjd161ljVVUkxJA6S0nJk7Zhd/qShdcb1ALnOe5iXb0OSR
//LyQz2es87cp0MnsPRQavQAAwErCEj+f9k4my/0uJBBacbLvLWORHHTapohwqr/
FN0RsJkISkIIiWfjk5wbkRIiPXTdWgAdt1jPBrs8bOOI7kRcNUzcNJ5pscMaZsfD
D4WrBH9Y0OPF/OzdolmTaPyRiuhB8GB9F1XppcMzm9H7o47G3rSNOYMALQ8dBG/P
p3sp3clai6ZMqtsdE41t4ZyUFV8NmnDvSnPP9VWg+YkRaursTzG0hRwkSJ6DiiTn
6pm+cqtN3LpBkR4xJ7KAQKwEvup69uaU8BWOnLUx4FTE9+JmuVH5l1swGXzIU9pn
+DXeZ2oS9eR6wtMQlW2dVwJ133uCuPMvnxZFb31CLXIfYZq40IXA/VJBIiUC8xf9
H+BPvdCrTlfjJiJBC1pKr8baDIaA5cwi9n7OfaUN9P3SkcfwHfGFW7waZH0FfYF7
9EsF2JRZgA3FxzsMkFhyZI+ZNe/obZ8TF9O6aCkH6gWMjoydwGbzKiFRdbzONqyT
K9XtvIT8TDgPb8a6KBc2ctb6SGJo11p0c/aUT5lpFz9tq5s9YOTC3UMfbbObzmZj
jKKvtgtqD4jsDO1hS53bYqy9kRPD6NGfDVy2z087SK04r3ra0of36jz91pBb1Gb2
dHzlefID91bimfugDweJK5I6OjRSu87z3sTK93g7R9OCyTmOxS6rtp9j9MRj/uzH
ILQa2oRnmrq++Zuk2mHbvpa7QAy6CT9vK/ruAoCBqrIXN3Q0xMpvXFJ77z9KzlwM
gx8mQ6LI4QxsnunQrKWNGmWA2uBh6xXzg2yOroM8p1tb7qjJOjBjsVOD2HrGzKYA
5QwHRO3XCFni0+32akz6pL19k1KefKPqkDEap5wzl2gGtuvy9RnpQzz3RIJs8Say
wfxBvrlQDkrt+YHlzTBTxyLYQOEoto9ntRcC9jjcf9IkZwi3xbhvSN/Bds9yxvt6
3GvY+JsA5UfKGII984x5yNUtXlyEKuhIAZ2RNxCcOn4WRMGTIsl7gNqFOv2zzXce
uk0PHlOGPh9PX7vMyWjRF5ppcclQddDrdijFQqEzdgwWhJPjAy6G+Jhgq2uGxB/x
5VPxFoHRzl9D7IzFqoUgm6WB2pr1qjGx4zanIeChwok45EUKpg3biY4Gd3DoflCO
bJ8E6mPaEWKMYShfjP//hrwhNmHIPTbfuMbxeJHe55e/yHMQFFW6RRMTyVz0Cjkx
jMCsuxbfTJrift/eCaFXwm5OdlfB2jNI91D0IQibuU4ihs/KyUgDyZYrlJUkLepv
Oh0uTCknZHz0iOYEmXj6Tg+JIbo52DQdNrlrLPHP+zku77ApuayljPzaGbv/D3mH
9PwFg4TIlKHbhuIN4/FqB4XXVlu4lFxm7vUsYMegriVtUuABspciwtd3XWSaLuoa
fT8MkkYXuyNGKj8V9bijGqiFK8fqqdl32K/NAYUHTjM++qHLl283CSLB4jEuXjRb
eCIn6TMG3w8fht0nwpmx2AI+5zkwxa9QKoa8xp6y9Gf+vGjT4B3KvC1EFIHSW0wY
RWWCF08Vbx2BGuzGVdQWhmSTNgrC5QXqHy668TEfGihiBdnCOjbQ1tgT3L5Ql1Eu
r4VtHhYqTVQOQfbYhDFrwXAEMr2iM/qfI8hLNdvwdOQpRf1hxoJRAfELZ1moJjNQ
5XdbqeW+wer3xpeahqSU+z3tyt9YUg0Yo287AZWee3epHj49VX6ZmFcEfEUOUSmI
xNyJSnvkzloaa0ZuePOAACwpB5bjBS5fGz2T04TRk92xrWlNW+WA7sUPYE5UmCT4
pEzWc/jLxtn31LJe3rDnkFNxi3Zg2AtJIp5xlH6WwycqbPR8xmI8N0NktVFAQ7/p
bl0OHaU1et7vFp9Bym+YKVy8B/89FZ/x8J+XEWP9oSOsi/eYY1Fa/ebQraGG6kph
P16AnJG+1y/HWVbzEbjMAcz/PS+LcVnlgbhQ09r0wl75MvHcrgh54r4DML7XwvIV
gXX1YprJM1n4dYQ81KJMacRIE8qtKRNFJsUlPVtnX/MQ41UByBu5P17NUfTuudwN
/2S1501xpKaCaYwfj5/Imp8+yNLe5PeMr7SfsWXFkm3ph07xo4iCYsCOZVjP9q/B
BHXalh31b2HyyIdlhn24nOAvu5HJLTpj8oMuL/zMdeLwTXqlqTAzgsPt4DQ36zPZ
tmMo9x4oyoQlvg7Xdz3ZbXEmGdSezMHZgyQzEQscfG4M4ikFhed3/9nvajuAm7fr
GBTIbdttzJwVofoF/8DIl/IzfdIY1WIgInjQOj9HuTwYKx88dycJmvZjDl23+dfm
vw5VeXQmCJSsZI7OFNqnCFqOCbFF187KrxQLBblAfGH8VMHAtxYH1BaW20qYTH/V
BbzJTwAkVFOpRioL6qMlgMbOCMsvJhqCuT5gY3fx3r49iSW1nGRWR0w6OMV9bBl+
kPyYJbik9pRnuaqn9CeSE2w+eu1rlnWzLrYfmK8/Eb89PVeZ0aHbJ9uoH6uChnDi
eJ6lnwHlxdxRu4VvaYih43MRrISYiXb94nzw9wrWTrnq8UZf0xU+ZIqizQsQgu/W
RD5bUD1WumjsWymWqR3AUPSu0gJzXchhQ4ZFKXOEkfi1uXfR/TwtjqyKyc/ZM5wC
0zL15GAlNiaO2UjAxL+If7DrkM1ghzhiUSYe6Bk8I3RyOR+9TO71JmWb5NShUYYg
PXPQJQ9HN4UGy7Jx2/pCd9mksabnG2xMv8ARmU0v8iJTMaj6o0VAxUPDLC52hDvd
Kjsmsy9twtfLdYgmYdhYluECxgBDCspe+Frm/PfHd/TB/yyZPnlxXx7zKik/zSLv
Dg5oyeMTS/Vuodf/pVkOhLG2EeclbVf88twB1wYlW8/Yd41YzkotPlFk7BgN9/w9
h04XFsDMSNDR4zNdlDxlwa36IW+SKwd9KQI19ATexAItDA9vmgd9zTumabIlavfP
3hvdH49iFOpGW2rSg2Jm24sZrvHieBJNEZ1FDBAPNwQ9tI7/0pbKLFAXYixm/vTl
gjiViulzWduyZEGj/FMhGOroaE3bkLqgcZ3oTma4CZh+VwYr+t9lsDpHrrJb3mwe
bUptrnmI5mTjU0nXgcf238KGCh4kURTTD4tw66JdGAZW7OFL8ogbGzsdu0FAQdgO
7FncMBEUYU76JQpRm4PlKOgAZQ3rVbuWYeNMFQ29MsVIAVVQiHN50BByO5NsUjIk
IBpq1HOtrkTYX6AvTuJkqmy6ChK+2l9IPedh0gO15HPFDeM0r/E+sLhtY72vlum8
+jPOXbgmParorTlAuqcPCTZIaGsR8gMlz2zq+azLS+QZHebgqr8VkoCMUkrNG9oe
BtDhkm/sdAeDxItfpb7dSCc20ew6tY7eBrtYJN+grS4BMvCFhlQdQV+twJBxnvNy
9MgjuYevHFcjS3M+CDyrNAECtx+/ZtmqIHYTrwFtV4Gw1XoTjxOWlKTRDFhoqMwm
I5st2/9RVyFOEas36qeUNACou6INv6UPy3q/zt93EjW05nfLZE4XnFK/3GZKDVVq
6Lz7vvgrCbTkjn2Nn3RWR50zO1KyxUHIk+h2ELlTo70RsD6kzZCvqs8k9nL9vsoz
6mNZgbt9A6/2JeV0AnN8rdq5JxLiiRIzclLOfuMGW1uukCh8rHCSQzI4CpZm3B/x
MD3R6fMlew0320mTikEx1BUFKd7PLqtCdoWoivBDyn16B8HB6QjcctsOg2f1ZcAO
/U964EDRShuYjvfeLBxEGrBVX2tPoSQ/ikZQMFONmWe4bP8RMOsnsSj+JULOpnPq
RKbV5FdZlbAYNuOQsrpyrLH3nOz139LAwkA5zkqWLoU7It7xs32Uai2qiqt5z3fH
bDdRU/KBUUZf4fajucMHAYxPxE53puiH3YGhqfHv41PJr25jDGGYJ6E9NNrpPt3h
DGVfCw7BC3Yh5nA4OFlycUdmHjQQDORTYMfYv220XIlcI9wU8drnftLSeqHV5/dQ
+VnETE7h0hrdumn1SNmReqbgOqXNasCik+ySK8rfZArFkDln//vybI6mQ6AXN2ZK
no19MQB0uAGIhwuIjLbH89iRHiRHZBxiZNFFZDqhQeBl+zNwaC6N01rXvjJ2QoQU
F8bMNt1o9yD1Uq0U5q4epOZpRIRivlG984XtA4CnS1TOGD/s68P66vWhUg+z4mab
wtforAzavLYrAAhQ3sn37zwQNDcBKkHiMDEO1UlpJs5UZ0uLlS7gHmO/0VqfDYPZ
+x3lEeFxX1kp5gevsgAocZPv7omAay2UWLAW4jkKftn7tTgQep0evmN0eZWZEDNm
lmo5faJEetR+xq+fsUNnECFyB8n6SyXmUR/actegmY8wGvkIUMkrYZ0btHebpboh
jQmN4fa1uRKFejNQyAjoaVPiBXILkioTAiSuMf68eR6oZRt8HGQM3WWp7M1QG2sv
Bw0zc/dAVaRfRpvxB03DrMHJeEyhZsZwFXTcU8TYBkG+ZehLMLXEH62DYP0oicik
Y37cLvCI5V47HEiYyoB3Mfm1xjv1szFwdGGB19zZnsLOFh0hcz2v0WNbBYoyEGmu
SO7eZnh2eZwyhoXKKk5PxzlXOFxpBfATomAngXP8hqLbViH0iyPxYscePT9R7piV
DzYKpsBE33/iSDclbmZOrZj0raVkaB8GrNF3wH6deVUZwJMlsss3xIiwebhZuxpN
1wnPXq489WuIuSnSTxv24NeuY5LkDNtANn5PKjP2OCDFXfjyL8HYhAea2CfSEOVp
xIZ3rnaO8RGobBeFCSTxUEF0HoLd/QwT4zA9/Rjg8xp4opRV/uiGXYWJYa8XRsl3
2jGiZAyPOYIYMgiOxfNMi5azv3P9/PRG445Hh5dm3LpYKe4uaz9kJtlxaN12/Aco
pYe0OVzWT7nNsEi8SbXmSPnF9LOlNLteNHNWFXlW2/1sR+kZ0yNnM9/EEf/oCD9a
BhMhwpVxCGhVgwpA18Oq3ldLxvgubasyFVaypmRi6gK1iqbtG+RlLk4YMerZobc/
cYEcwc4F73cL7VlRsW32dyOgT2JA/azShs2EvW4FedFsyJfahrDzypL7NzGBWXkE
NvtV0Kxje8DcUggpfJasmK017y+srt0XkK6SiybmxRIaNyILUKlbKMK6jjGpr4BV
gn0rquJhf4TLwsw2KKY1PC4EQbwDDvGLX826dc9waoi7YOL4HpOXhHvkydx4hYIa
CeTF1hlnu+oa4M80z0kfjUjMsHMy2fSKIpq/u6lgFWklOjtm7xb2TomQ+eYbTmnv
sB5pTSVnyx7n2RESEImVRfsp7bMoibsXa8NhZMknnzh85Epk2jUfyTbSBUlWDrF8
0ay879ydOnvHOsC317QXmRA6r0IKfW/AxEo1SNdKillh/UQEAvELqGz2qycTPUDJ
TAlQ5xnz+MoDRmQ2XlbLOJLz4Hs9O4gnbpbIjBo4wwdeAlJp4rGzBs4ct8If8YyW
BudSTHd78qgtlnVG9Co3pDiygIg1Em1qa9aBtVbVYXog0sre4i50VlhDX52u4jmx
YrH5VMlnyNFybUCXnqDGLoNW/6XmTxXIGgBylsEeRzs33bW8O7NaMuac4z7XFrL5
VEdSgkxU2V85oYzvBkxZj0ogLj+aFPkG1iq5ADm4twHmF7vYLXHW6ABFTyxsI3vU
ozWLuXXB/dvOlpMdSDbnJQdNN27v0VhUHzEMToeQ99dVlPgH8QIHp8rb5CGnHDkW
2mGFl/ST1uKFn4aIiv+ziQNxLl+dfXX9Hm7WrCamE/XEYdO52+f/B2NrPmVG78w1
D0Y3Ed8OxwirWOLFl/uNjPygD8ySCD3TsJSmmHyZkJw0OmPxVgKN3cNdwao1rV6Y
518j9NbeMxZ0Pw3XIW1g7GPLGiWFGvGK37db5zgMuft1PIg+1Xca+t5rDELZNrt/
0gXf6gulMTsgrTxDGmPemlk8+LoOI0hSiUypMJh7iVoEojiapuUb9m+nLZlH5Ubb
O4QOiH65fkz+UxPyHT/lj9tIx2OMPJ7H0C23GHijoGft9nUe0zYjn+Qbcg1b+4Rq
mziZB3JVHPjERj4UfcYc4uhbT2gsb0eaozC4hicpb4gvYT2csZvSWxaOFafUo04N
qzhdJx9U+lWOimbRQnTbq1WqgOsgShoYaOXsymWYw1JQ6BsfU9aJGbaMWgld1xz1
NKNXx+atJ9D+ZeXeI9l1u8JKtu3sLLk3usas23eXcT06BnAw/0LspdcrCOE+Cp6X
ga8YE6yGg+2SYgKWFz8NZ/LLL/o1Gt8pVTKIPr0f1vaZCVUMUpctv9dVsr33vCBU
N59pmRjf4pnwlBEa4oT0z5Mmtrxgt62kwNb1it32Zp8+8FfoIwDRvpEzZce17u4I
FFlU2fxOYJRjrrOK32NIKiacRZ2cCAUQ8nCEFbfZklkugMOj0jCCmf9hkPR3bfLw
0nUGOMvGrdzSUWxND35RF+XjjpMCy8sJwhdxhgf3V0OrKzGvRJw8RHzYmEOvJBDF
o4UVkkchhlAeoYnyRtGGCReMKqafkI4HeDNC0GI5laolOHe/oOhF/ddkcEr8Mg42
xefXroF4+DCDjMGTLS03AB+uhEPC/LgTVih91uEx6plV1wfGnWKNPgd5DjBglJ4T
LPaKWrszJVeHtpYurRT2SEOrEH+PvyuPbohnsIl5cH1scZQ/R8rBzdax3FpGs+TD
5NgS1SMXUTrlM3M7GI32gQRHz+aecdVfjfIdyoi2dZpf1gJsYOW942ecMKuxc403
x24Onqq8N7WHf7j92kjqxgJrtwtHXigEvgIlNbrcAGmqG/g0L4n+O6kXqbdAGpN2
oMTI4jpELiL2IVJMClbzHp8O8A927MinP7KPOb224HisLKGMKkx3aHCd/iNyqhT4
py4QPbDOFMxUkIo1fHvUvvuxs40IYQ+U1/5Nf/nOt71CLV3RnVUR0jRlyLvbDcK0
iGJiolB0Ld9n1POxyZQRXzc4xT9Hl3MSedFF808ny0HIPxs0yANUcUR4Uv+IZTsg
rG84s/vLRZ6kLpD3V8L9R1sgOstN/qgQADC7xSkibUKx/Cmuj3tfPqIrkONb50Y+
/42n15Y2WNyUDqNmi6GfwK4FCWBgUCJrkQBFxT7p3GGwvveCdf6uZ09qnDoxThHW
c4RzkU2d4QIeAELVmRYVYErB2aVuu08B+O/xMoK73s4+Gwqv33s0DSmQNLKV7p0Z
cRBtRiUZUrry+E1+3v+Ld1izO9q/I0veb85r53p4ubpgyk0lkB0LNpOZcWWrZGny
qn1cYFN9+LegB7UWruoxzgS7lZRZQ2GvMh3s0VFpu4JF1UAO03uRI1bKiGGINbOv
w9lAyB+jZcrfOKmFSAp/HBPOGIip4LksZElLWyrjdSq/iV0EMH2m++O6fYzJUxXv
8P8zFgtWPICE8qVYU862Lw3Z6tCkiwJPTiDwSh8VWy6YFfRQ/4aX775brFx2jtQM
p1tBqiuR+lyOstFWSw9YFVvixaWNMyQVFClcBPjtGjqyetHKMQqiI9Fsb6qH8MUM
Q8LHyJfCp3DcLpgP6BCV7piIjE2Q1LuXOxIAA36ZKWO98AIHD7bY7mS9eMNh78mq
iTyurQDI25aB/JnReAU4h6PgxdbejumP4yUw57FMsCLjmtzpgptR2yS0WZVxk9YS
9kehPwmLZdSzM0z+0bYd5eFEaPo5MUVAxUTBAZqeywYx8fPen1d2mmeSx3pHCU9J
XSkJFPjIUXx+j+UfsJXUmVCQ1n0zv1k+pd5h07GkVZhO40XkwRKjnWGOCdZ2r109
eHcWGjjLvG/nhF5B2SZRIKg/DPx09PwNEYXwoJPIfc48kV5G9BpXvAjN/TgFaT/W
hyhiITZSHo4ZcpiXMnYTeTme19II2saDQgDvsQJeZPBI/sr4CyPO5I7SlDDxG7Tb
o5siNBq56bExounmDfoID8Mukrkq7RygR1DGlmZCWiwCDbxOqB+2OEN2V3CVdyIu
Rdkx2mnB2xlNtMxspUKvvIFKbedWeinRu/EhuB7ygCU1nT+L3EblHxyu90tJlMmd
6wFqQfmvcGXymxLa4/pCaZi838nF3zdSOt/yCqMrqxJhZIScogf1Kflexe4rhka8
PVHnz1OLDM8PcBt0V3KYehmS4HD+HNe22O+C1FIZgDoB7lEPvpQj3UyyLuzr/xSt
ttgZ4+pbvdyn4FRH37yYntnaayYKlZ5N/eOZFLZJ5xQ/TjDIpuPKn6Lix47fM1Hb
b24MCRw1r6xUCYg6O6WXdzewt3yC6AY/iS+hsGpfMOGFh9yEN/JZC782DIol+L5f
GQhQQOf5cGdT+1KHMBGMptK2BEn/UEx08RWhq6/IejlGC3vT5xwAQ+gpDg9na90O
oIs1/oYCyrA1EmWniAFu2p1wBZ9l4UJ+wFuWof4hA5mz4W9FEZmxeOuYRFH+ulDk
e4TA+SsYld7Nd16R7rBpMjmrEG/gIefcvjSOhFH6XfjD5wR5GiwRXWNcTtXSczH7
mgnZcWvBb+Xx9nCQAYv8jIRWnXVZv4AkWpOZ1m4KhV0oDcJ66IP9nM3UtqBVxCy5
mSg5To5u1Jd0orE16rNXx7fR8vV6btEC8cGwAes8f5FqiB+0ynW2g+cTgs0Kfo8u
zH9kiATxi8z4Vh0UBAv7pl+0ZxV1mfSo/2RagVwzDHhzEnxgtco98kO9nFrGhlWR
txJmVc+rxbF3k/qTRuib8SHs/3jlXhlE1COziaaXEhh3RVnTg1S7L1x1amNteNo0
amwA3UUEN/ddEOUwYvtgvUkLTz55TFuF91nNc5dob94q5GKdRT+AX5hoxlvIcohn
DkKCNOS7VaQ+FmhQdvTi3TOPbHBdLdmhA1S3HOZCFIUn58ec1/nV3No8rrJWwRCq
ti9bxsO4ANDnKPwfl7oHVvcdrAhV9Cg+KOkiyPOAVHy3ugkywaFwHlUi/YG6fTWo
oGOudYhZHzGDQftUQZ4xg19DMFYXQqjfm86CUHRCjyuKPhWMyZZaXF8dPPkK+Obu
hOCFlW/M6yPk2BwdsH+Ox0DTrfwPJW4u906DLh0GdbRVSEhQ8JmvKml7Dqwtyi2l
9vYw7x+JpWKDM/BqKOsze3I4i5XI/8cBE6GbkOCogZAIhnDZDbOt67Y1Bad02ZDe
or/qBsp4ocS3k9unUeXsdkyF6RRggfYUxRMjIiuVj9LOP6V1mou0lADwJ6ALuehi
HieM2ggiLUUcf0ii1AT4ziczSaUcqmIOPgvnhdVA/CiK1v3BzF9PetPjg9d5I33+
RyQF3ypidY90X+4DMA9DfzToIDs5jq18Tkhpj/2DtsTNB3wq7ScAgxPB5BY8p51o
QVTgy2+2+RR/aGlrfhIELGjBdjgwmMYvIqR9jjeJPPc7PfgcIJGbfi6TK5HvLD+9
Bf/j06qBpJklb5z07tX4pym6APY2A8TzbI+ET5+kWprv1Ss1hk4FJ4qVy96v1QM0
hVcHF6HK3GnQUEtlmsGqY7B1z+mgDKgNmw+gqhhq0pUe3qVWlbbTQOfxBOVOVnm9
McHQIaxGabF+i/MJE9CwGqPgSnY7W24RoZi3r3dthu/Hx2mvpTAfZqIQt70ww16F
Me29mEwwL1WQDh7OR4LCqAwnfHvoMfhDjQyBkqFsSvYpkgIdIAOkLiNyReZkB+ev
ytz5RWVSMyqq04gx+wjlOvrNppZtNzANhOjm+ATXyH6MZABmoXHhJiWw1/xvOyoC
P0mXzWM8qzJOZ5ju/5s0ZmQr8X50+p1eSmzKrvWwA0557U9PBS1Az/TdTETPyECw
77BaUbwxfmOYVtBTz0UpEzmemNoBziHXaivEzKgQW9OFCDFMcnT1rwbGSGznQN5K
QPK4v+tVlQjmNtP9KPecrV6ub4ziSpHHYQpJC+9glYhs7afj6CyDO0IORxYV3Kdj
tD16ixbyMzbahrYtXADtLWP2vEVBMk1TD14lMVTE9vl56vU8igEjBguu4G3/o1ZQ
NSDgSoMWrnoupA4fMdCN6AnsFKvAR/x34L5RRc10Mm5+azdNJHXIrmtkvKcaWjwg
W6MmkJ2E2kkqYH6i1xy34v3cS+JKdT96xvCiAje3U8biy34T6ogncjxW8BUAbYvk
SCsOaC2/uVwDuUiC67455FYERZakYauVII+8GljYyXh1V7wn2Ftk4quefkBdBw2k
+dqAfRGGkqw0Ox55TOU9ssCcXU9mcFRtVbvPv7FFUIo/e1Kx6SRjuIFy9Z2Tvubf
53DB0pTB63lDvIKbYRIlBCZdaiGUprEBe1NR2Lug1I/6yd9xtCZTaWFqp47+znGR
8wBtzm9aySuxmGDUcg8X22+VnlVK9HBXCvvrr3vis0u7ho6QAh2gjRtCaPQoi1zQ
GXCNEkkM6HpvJMMcnzhb/9XSWMYHQZ9f721/G1y7KczbNwCwOTwCb2iddhPscwO/
qEBxvBf2I2Slb6wdzaOVibufWb99BjiETo4B9KlNjS77bJwCh370VScUssKbFP8S
fYkSdKedE8UiyKXFbnWl8l9z3xo+UnRY9bomIMuMSSgnlXfmMU1Pc/a+UnG++XRi
wRhOkZlYI+N8lfFy/0oNiOu8rIW+U9LhqiVMhNI39GyISsROEC0uN2Xc+B74vDeB
Vkzook560aXsMzVrAzkCee/W0FClhKJnWrDF7EtV6sCRxBJU3bPeJIoUt+65iCbk
5GDL62lWbk1nmAzuzU1BZO2Vk6GutqDLlo/fGhlGHSqJpHKSFqrFpNf6RK0H4zS1
QGXx/qIBlLqXfySGs/wj6PtdwNGSWLZ4kGTa3+BoEmjDnzXIrj/jBYNe73iiVs0l
ojG5H2EuCqdtE+8GpqkoRcZwY5p3hIWlHNdaG1qg5rZi4RQDQNCs35bi0QNz5mB5
8u6OqA22Ej1smI47UpATCexdk3ooNUxBedJPTmCoIPgTY4d7viNJ7EEItu/VPcQR
QGDnI4onKcKVpeBEi9V/+zMA4S4+q2VA28XK5yuV/e5TplseFuGTiyjCFThFU/lp
CoslJQFxDb9iIfInGDQBUEOod/dcMpEfvJMzZz3I4gGdLGlSP8qATL505F7OCMwr
3BjHyKHv+D7HZWRJwK9wYAawTLVqpzFsvG/LAzS2l1UUdu2IZm2/O7+zFTU7knLs
9v7uk/FWroWJmpyoJLpxswAfkOlRgZBQuk2dGKz75POadVzd7VJx287aUlfGP7JY
Y41y6wPbJKMZzuoi3AmgdJZyxRm98q9ai/ltiyYNQnmnjOjyYQ5k5awpJxuEVwso
+iOi/EFnXnT5SI/JMiR8WU6z24EXTw05PQq7BcZ0Z6hbBK5DmhFWJfnJMPBjLDUk
M9BQZgTOr379wlZ/dmDthP/O0mCFhfZxjGZaZn6Yu6GC5x+HD0ZJQRjenVYccH7E
kAZaa84XVyya1Dtv7q6Cmd69BxrOHgkaBZC7nR14WYij7Y6azqBQ2EIcXzrAfslp
DKezETVEaDtcV9JT6LaXyy7S4YFKZSpe6Es1YUaA1ImphXtADplUTZXqokrZ0Ue1
STC3WvOe7jTTHWRn5SKWAKZcatus5Qde6mG6RuQ7zeZB5UBf1/PFy3gQNpP3TE15
75M8PS4j4RtRZWKbgLSm+4vKKbIes/cMmpB4PtMk2YNPziqenZH6/5b/QSSjZHKR
Ggo4HnPRU1v/NS9DhKh8RNfLWxSQdlq6Kbb4WwJoLir3cCKEUrBrFaWrDX+QnBBa
BKP3K0TbBnYU9RVJqaG0y+bEqBp9h4Div1ft0tpji1mMbHNXVb9C3t6TWoZ4xc50
z+vygWonr+gGR/7r0Mmc1icazzhOKDJvAyRHfOM3R3pgtyg4NUndPg/xPlJoC/FM
lUauXFbLDeQaLBojRBQIZ9bG7okA2UfEBMYhChuKXiJN3/5AwI4A2wQmL/SR/PQG
fssmznAKYc7iWqweiYTNgpxflm0pLEsNUTfasZxvsupfYBYPDRGah7xSDPUpeOkh
NVlp3d+hz6jrSCxAz9sijP4aUCzvw9+doTtiOT4BkPsoYYnEF4I/ONKiFO10coeI
A0EnBd8gVhOcr+4/DaHQhgvbBUAZh02PaBucbGaGDmCLpdU8Xx6gYk4veW3xXAJA
IP1NnszKo+qWFLTLxxVAPGqd3yuPBGCupQG19QrJ2UY/Uo2T9bVpgFWwQjkWZlfq
E426KuPKKhh+2saGF++PAo1s0zvlYEKSnPk16fXfPd0L5pYRpJyzv/ZXWuicpTl+
L/LhOt4UVxShS5NhuGbAP4KZ9d6it0sZkXddRquHEj9EB70jnVVNPAb5VEYVzvh8
UAH16HeDAL8mKLwEhWOQ6A0FezmUSGwft/DpQMFZ0cjRnwQteFwGmb4NSzGNW74c
M2vKU12/aKbWGFgVFj7CBZJXqNJzcmCpOBZBF8fu6LDunsT9JYC8hKBbPu18VylE
rh7ATNTKMzm7wSvpvngTsMXEaFO5M+fHgUf1c1QrbsKPqQFfERCpoQi+b9FoYX0+
yFqKv33yhiKvO7+KV3gyPELCBbfTOsqzj5We/g5h66cmXGg3JshYSQbJKkX86szI
tTyjr/1KJSJMXiwG7lBolD1T1OaSWW0G+Q9XDTR8TnYVDBRPc6ufke+5/rVZIXeU
o5/XLV9miKUhmhnhwt8wZy3KPotjewZeFOvlMEHB3EvgjuxwAVCq7pY0WMFsQomd
Qqv6NoZEzozdzETrONbSHwqpmJ3KhVMEfN3L72IO2XyNYnnBAG9mgdEYSHxEXQx4
HLqhi3m1UZi5G1GpOnYrNwZHIpvTqf8ULUjHrDviCkG67KmL2S5kBe81AqNIOvYb
TE4SeN1PO7TPbhf8HpGOn8V1d3ZSV25EFseq0jSMbmVXpVDUJBQfDtmBNn495FMd
IsRasmjMQdmkYy4KP95O6k+rSTn9HzoLba2ANgY9Zas4xEZOZ3P9IYvBghGVn/JU
1icydJ99i/1pGsJiC1RQmOkX0D/IrVGAB2oTfn4bPXvt+6oSDLbjbnKGPNnmk86z
VWJNj1x+j7V6Vh9pbUujdd+2miOjz7RDgyxfIBZpnBLioUfYJ6K9SDnKFAHdBBw7
TU5esiiIPdjsRmeifXAM8HUEA3ofsf9NZ4ULdKP6LU12LkRmp+MrQUtRJPoBi+5V
2meAYmWtleC/T+Bkmi8Q4qnN0caxdBHrgfxwvMaAtOzaSqu1sHlHu6D2ISLLNw/p
MRVErVAT0LpCD+b+2kGrD+9O/wtorKkpbkAAHhcQLH/d0V+pkkYhszogycfbmvmk
on4zP9QR0SPSZqS4J7DjMF4yN33dmj+OPzBfLF72JaCbTdFKsQaIYrAwTjg4fviu
GWZ+CJ6V9n9JeKAk/Gv+2lz2md96+99xSrxY/iwOk5xLaAYavyhFXG18xHaNbuoj
QGVvmbi3YODS/V4hpcOTZffnA1Fisop32G4EmNnzVTPc/vm2XSNdh+eXZrE2kwsq
vxjn0c8BbDppd9f+zWa+I0qTNjp0k7DzkoMZj9PM6yxbzlp7nWjC1JuaYI7rbATX
W5NZH/ehu9kB5ESkTAxiR7G8VbYM+FuCLEVR2gsZ/nYYbyQc7Edn6uhrYu5sPH6u
7PSJ5W+NYDyqoiMQZ6CA7gCnWVJFLBMyLpH3LLtcWR0lNMSbGObevR1Lo9amW1eY
fvuH23IUmp3LJiQfjiaWMHn97o0NkuP9kK2RT9wsXriYbRBd4ES8A2yYeup1gbtQ
jHN+PknAYQMnHFVqgvhVWZkWAke7D9k5jB6BZsGXXIDLSf5g/2MBMvsctq5pCXKD
YS84ymPR1SZYyBfVClKpKTWNs1hmDityRUVsFtVyCaq5FYoXl2SAClwlZ1qwLx9T
RHQ/cduB1bmBujAnIJQnt7xOs0fBWdE1sX+sna4R/idxTsHzAKbNhuxDd7MZphcY
amiPfTs5/icf0jlM0MlGJUyLbyEBBusCXYxmqXOrE+XFx7yctMM1tt1s6PiTcotN
aygY3Xyd4BNxuJYkazOU+CTpkvLWtrySVPGaltoJvVGxzu03MgSmX5/yO0NnSV3o
ulXnXX5OEbTvHSQwO0vaKHayltRRYS96tT8NkLMN2V69iDh8ixoG/+yyqaK+ZPka
kj7LoCVDu6i0mB7XyAKjwXdNjByKkYjmn1REMggzpLEQ48BONEVrwJ9G3ljxgb6y
KQdVmf5oDs+rIxSiM30ZTXUEgPSa/GwGoreQBulv82hxoPMwkfwTnTnQDpMkKMbs
ozbaFiKmFh+892mHYtaM9RFSrPcbA4aAA4jDQwwVF4lHtNXZAWfmWKphNYsr2pJh
x0UfhF3VYL9aWYZsYRrKaHztSLHO/pwBjAyxR71WMYo13y/LLDi31IzMBKAI5/Sp
I9jh4IDUNIdvErdzJ9WQDKuFSm3qKg490Uwr7g6oNrzuktur4L1SVP94qTDrlc+6
4MYDQjRq3K8L2rCA3fkbJ1FpNHMKD5N8FWOziL9ftaqx/H7wxwQ5QdctOhOY6HDU
fTD79JdKa9SUSDUKdvfh5UnID4nVtGOF6/rqj7jDY1rsVufZisrKZaIF/LoTbHW7
Vg8ghjzwivZ05+yB84040Oldst3K9p0eM0EL++u8kVe9C5x4imDrBZUY+EIrfkh5
9eXBBxw+Xrnt4eW3MNWqoXR0/ljRRxZNpSiBYQ2Gu28D2dbgKDRE9j8XSv7aQufz
JfwnkOt0gI29Oj5KiQPL6uCweqbjVUaid4nrSieQWzA8KQwwwknLYVDUADob8MM0
1E24Zxs2r0y4bbfXRIDLRazPCNlMUsfp5JlguxRkZ7D8j/adaw3UHfqDFF0mqfv5
LOlaxImftNp2TbBAJpq3VaMyP4F7AGnee7Hx4DbpFtthHZrx//ScVgoiC14WdLqX
eoBSQ0wq2ApQ8n0gzZ4viJN9FYr/IKM8xp7dEAJK+YVub56cimQtMLSDJE7CNNNV
UqkfgWQsyPodqcWGOqp3NNK+kEyVEF2uV53xdqaJ4Vd0vYLNbPYblzm2Q6ODRO6S
qK3d+G30wudnvRh/CewgAVoOugDqPKpt8fmS1tAF4FjtNjPsAas5uAJ+8pxIQjsF
WKAKldMnuARXY99ZKX3NbZUi9eZAOgRBZ9Qt1ZgpgK5koeyTPuvLfrKMY4gURyyF
tp+JqQvvcU8TPV0B4o9KjmL9ZO29qubgbbmov+KCa9dR8RLsNbxyLl3mkzXXgPu4
JVPMLFICeDHk0RTMlMl/4jwJ9Uc8GtRIJFig9XgELOaKMS3wIHSf18qaA8e3bJOR
29AYkxNxU4s1rpGL/JscmyFETyksmA1HMaNHlyF0lj5k/+G9l1iHHeqB4ep8A2b/
duMit+1lWkUf7u48RDGSYbAA40PdHY0tLWCrRppidKhi2Kf38sVBQDChmhw4jHPU
JTRBvdgOVZTcF07khR6/fKQlM0xeSbvz5MPvp7O9LPgNjhg1BWssaSrnRz0Fn0gy
QyMOx9M9MogwHukxgl1D3iqHR514m8D0oRfYR/5JXWKf201dvC9q+4wiQ/UuCEMq
JIJgM+/B2YNwThE3+txPSw8irmattepKIHs39eJqUgsk96tgSnEdaeYA1T/uOHpL
ui/fbVrR/qH3ddJAY0p6EY/606bo8eHnEQkVOdblsecJ7L6Mj2Oiiqp2RW1wmlVu
+xugoGPf+b3kRbs5eCrUdWX2vCoiIon6mWu72FHvoWf2gYdeC1t4zilkmPwQoXFq
g77BBJto5I7n2n0a7z52ZuEj6fE+aRwUpMCWoc3ee++vQve+SSGHO4KtKRvLcqwR
VWqXlHrZQbu6fjz8lCTbTbRAQg+ykUBYdDPcVa7mEvOlGurF/Ctb6Vwc2KXJsN3F
HBPUNdp3dP2iCN9TDfg9h5qidOdtKDJm5VoEb7gnyCo1Ok5VAI9IV7PHijkH3WsA
zEObVAeSEOSaUGBLMZCpZ/Dy4yteRVAPU6b5Ds0jJ89WRJLcD8NHCl0Y7zSOHUG5
JtZqrgVGWPHTBD7xNIyHxolwLJBcVjSDEyzTpWYxj+Z9diuKTQlx0yxq1OcPLFpW
LBSSI2eAJd44eLMDRZOLFWSi0zJZkGndrc8R75QULAPlBkK9b9r+urEtXFy8IWvd
zPOLJapfWIH9fTkvac52FdYjOQfc67d7QjcniiPhfXkgbTGBD/dMSnGXcnQQE0tF
CDN59QkIRTM7rnKFGAI2XFjWooZZZR6LQ8DfaH8qze8bHtMevSduVnCb4vzi8i02
gt5ODEpCzfAgCN15ndh2//su7g3siF0iZCVbaXZILQZcDjVa9ZtXmTSqPAcFAJeP
JecDiKt3fkVZoytKxrtSOmiIh31U9NGXd90/oHYvMSmU/2kgkGGG/CS56jwBjAfH
pL/yOMJRahBzDHyZipndEu4fxNbj97bX9kQkliUpHnz7+wEGJg2AI9Ws3UDf5NSH
6vtYLkUXBO5okN88r8YTYrQtS51ha4r3rFb9lWPs+3vWpJTU35FpraoALyFLCTFO
iEXU91ay04nlFTu/zVT5lYeXwbQaRw3Bj3p6x0LtSEwRy9+SxnsDWDFg+2UbAKUL
CDuOVgOm+Jh7sQ/s20lLJYuq0gVcOsi6wCeI073F5Kz4Fka0a7uc0KOR37zctCLQ
mYIi8OlvuDif8G/BfcQFw8PZulgXWyGiokj5e+gP7zJrYIRRXGRRLzrUSykLXLCT
ernZuXW7anC58U9RQ2dQQkklBO6x1n6HX41qDGkHoXOK0BuswB30StA/sZ5jrKXo
TyMPrfxEFnkHvHNs7EbBNgPiGs6P8VmvVwGa/FrRv2ybcxnVExreAu//x8LfBx8Y
iyL9BoW7RQ8Qa23cMZIzuAlNnZPg/WDtcR2622Y4pT+8PBtVp8VFN46RBOWijJ1C
ELkJVsO9MHGBMq979LBDIQIOY+K1HHIVQn2dlzD0e4QObxy76j+FhiBF7YzeOUpb
pPLAkbrWApu1bu0IxALO8wPaYb7FvMn3+i3kWXyT84cVN+3y+aspNyctJdcxZR+u
uErFywK8Rhgi6bVAIdBGbk2LW/uD0jkfKoVLf8wbqtqjhMWR3mJDaVRDhyQmm2ka
ycxFu9hrjq6NJKAIQoSgVRHhKFXQ03eZmWb0EDrGX6Wrb8C7Pf1Eq1SbtopJwu4v
7sxFsXM6nfd+vqnrnYoP9mGYGM6IfYCrl5DjnPU+TJzMH8Aj/XnVICdpGGmeWjeX
zACCefVk5eg97Np4JRkso8PzeXxIpxq8+OjuSIKJuozgsEIG4hIqmRF8Arw6FTjw
kZEM0iJefjvueG2KDp7ZEYoChCg4Osrv4vgycjodaRo7MXguSbXuihkKZ8pzncCG
urIFzVvTxhR+fOPqici4QI+ESO79dAgi3elLAUsGJzEoEdbumJJGfyuD1bORL7IT
TL88+UNN/9vSBx4KOv0uY44DivJjH1S+j8nZGvWon1LsPWirj6kanpQfZRFAFiNR
9cc4+fL5oRgimIvvPzcMCUx7tM0T920hsZW1telEB3arbpIejz4ylRlNiAAb1I4S
DfSmdGNIno9Zi+76jEmulk/ei9C3xMsRgemc31p2YhlV7F6ZmyxUjmNLT1eKIfov
kpYyjKdDHqLQYW+wDdxJa6X25bHRi5yCv8y/FgppW4/wXpI34XzS26QPSBfkD7fp
1rNAWiWSe0ENp2rPGJ3Fn0ijEMdryQaQvhyxlRkbSTuE4RUw3qcUoby8yJO7IMNl
XlV1MDd4KTt3ccPY4FvN+8sLV07bMVJ2YQJjLtHIxfSVFHAczXsTDq7QsfJCLYZW
oIR7sOxcW3o1ti0bF/DfLIaD1p2xi2W6jU1RTm+nI+jf9Rd3b5epgu4i6r37nupA
gQpulGbb0PeuF5PDSc0WkbiN8ZnkZnl9cig8o8+dMpueMDhDbkh8mz5VmLb7xxHf
8FYgUfeLDHsY1TA4YyR4w8GGlbFcd4Oc0j/0KMPN+STGyqKbX3+I1Q0QBkaEtzFI
VLnMIYmrsCppwhO8MQejOMJ481HxkdJEdvYd4nUayK9OII1YxNIIug4xJ6czmEDz
aHlku4afPTbzLHFYu5twhnClCOmBGm1i+KktXPQH8NESKMFqEc6ptcSOPPqbfxZq
DXFYpa3zsANAYLaRkTTnISLsBis0TW7yOmsfVFemDltfQosNuF81gIsZQ7D8u34a
MWx62qDSqgwGtLj+q16AMf5qJPXjYsoObfR5mLnXXfCi1jRJcbedTWFTMgbw21Vh
mpb40I0tci3Ld/iGs5EHq1pDY8cpa+L3wisx0oKQP0gFXZ1d9WD68HZbvT0u2zU2
KB7SZMR6hSkE3NN6jULlLb+ZIk8PcCDGWKLjXxM4KJ5LefaUg+fBAQl2rQC6WWYt
FKw8d4quq7c5+rA6hxZKmt1VNdGjY8GHPEzv7wS+oGVwU7GSs8hxN0lFO5A5P83R
JERbjLeBrEC8XTbU8YrmQFQxtR5I2/+SgSlFCP/hfJJfLUB8pAX4ktljKopQtBDt
0bAQ1sHUXP+m1bR/IJPUxtQqoYMbzaUcbioP50EvpANCkicmhNmjQWZrh1BkYLia
YkrzoOWYqzp0AKqYvLNp8Nomjqb8ENZb5QHqmjwswWF0qnN8qtbSzIK2lANUOWiP
YSIf90KuoynEioiOenLUKZg+FWJvPKYWfCfcMHiWxRW/LFBbim5iqAC7VFLm5Ul3
g1j8F7L9qAUOzaSoM3ovVke2GAV+6XxvqyI7y+FJMNdBjfFb/YxDR8EJVB364Lxd
XrvMlxKu+X0oo9qTrKBCmjcX8MTuw1j9RefDwAbgH831jg+drlGFg2eKOyRRv5PK
7GLUhIa4V/QFxDdTvmwNIuVMzdsfpQHvMRzlhPBjiMa+pGyVogBjNBJLwzlluk6j
829057z13jm0jsmJW1YeCtrgPy29rHGZ/vndI6dtxCVwzY0KgOOlEw/a9enc6a7O
0LjhzdZhz9AG9AsMYa1+Yu8NHK/E6zDpjuRaERIdn8JxJBkPB0pHG2ZxGlLXWfmx
x7LQ2hqFJKkrqAlIKwcqqx2BygKBUK6wHdsXF6ILJMRCu2q1IW7BL7XuE9KcTsOm
sx0P0/bh0HBiQ81CBu7jIZT2i7Ke9ZULkrwX5qBUCfhNEm5ReWvHXDOg4duGbj4S
6FCfyZKRBmbRankEvZI3fRSEmUIK1ba3E6auNEApBfZYfGNkASXOi+wK6fFwT0NS
+GFcPGDqLyY8J5FT0p0l+bmRTwl0Z+lWktVKuY/Qzyeh6iAxJXn0296HM9QdDB1L
Iwairm3EVxfyDum6rnd7GQYYGXsac9I/4BuV4/2wRtwrQna/Xadyjiukh7F0Txc4
/cHJEAbpZ2w519dIYCA580bDW6YaTONXeTYDSzElRzK0+cWVtlJy/3Rdk959qe7l
K4O/kqdVqflPmDXydE3xi8Y+qmeuvZ8wXKodFzL0KSYjAvhbxI9ymSncxZ9yicgn
pB6TGkt5k2oBRsXeWUxehVrhYi8ryFzcE4/hcMv7AcnczIQEModEvRxqEvrjAHHn
5HE/vNuNkTKgJipC10zWxBruKSKZ+2cBbeu0Rwb1fe61Nc0i+h+2Qup4xVi7hz8f
siYEqsBMfAqZe1mT8l02v7MSeQubiA4Wk6KTtplBDqCxHB2m1PY22lsXcyySs+tb
3JMiNof9Z1cuP7JAcaG8/GI+GRh8ap99eA8O4yb5BVJjnb/A2OuDqm6303m1xaj8
/XuaA9mSnPftvPdvwEB40XFQ8pCA7P7Rz0PW+q6pQBEQeeDU5HE0egoc5TFUVWqB
H9hfDg873Y/Qslde48FvSXU3OV9zdgBPE7KCC36/Z2LMPZR3ztQERcQcfeEUcDzX
n6517+S+fRfjJnPmm/nl4GnI1fY4KHn4Ns0LwagwndfsDTaUFNU6D3gVQVMBhfYr
+l2TJ5/iLEPYr/5+byUHlN5jUhpa47IfB+UfwpuWwPg5MGSS0mhnzKyEJ5nkkndu
ZJEsuZmRxp5n++IzVDMrEIfp7L5mOLk6bXIYHthE7ms4eonQmp+GhIYC3vHJSutK
nDDFQeXwpMwTu7P6aZ5NARWvrn5D7QCfz5ysvByjMXfuxy6i+IVvkgFHn3qiCcbR
qmMOEmor+16UAXVpQqSLkFumv6rL+Ck4ylOQGRpGxlmV5PcGpMUnbQiBoKzCh2eF
n75/GogY7t3I/d79fvzW28HTC1Jbjcrnj2VddOGBf4PaeS93J7h8ol4eFWt+cGRm
u8tVUx53qVJKpndMsSEqiNGNEhad1RqXkwmj7Eu3EUVtyfRA9k7YOs47B4Wk6L7/
PldcDzNA3IuIeaL69olYC6OVSm79Xgc2DoEaDnD0UcUpaRkRBwRwR4EFcDjrSf09
XMKl5f/1N1PGvuXJxnXU9KsTPYNfhASiHnMdwWZoSKoNaqTmOCYBba9b8ndpYFcZ
C2imbDa3hRTwcJ1esziRXDy2y5sdWyE5LcoQ+5CFxMh/PPU4hx3jxM7uqccCurE2
1B4d8Qnh5AjdbvMie0FdDoPiMoUN8/fVx92hZNDU2E7zRh6a6F57kPV/nNlqMfXH
mE6j0qj0E/C+gePQX8R28bqoFZJzdKZ8xnb+BXIMpLtqyqk8nmVFxOpKwwn1swJD
6IWkZBDadanyaUye0n2MzkcAXAHAnC1Qc6M5NwnOb/hSNnL2mKcgB4BkM7Si6RP/
dzivXyrRY8eQAxRAMUJ0Oojflbtu+MZnZ5qH5Z2cyrWFY9rXXH21Rk5QkKc+fPiX
a6IBVNbujVPeeYyzK9uWg/ibYQUQZfKVn55Q/BHlNTX+LyjZJSbPLLQB0/DAboQv
nABhxjzZ4vDsk/VQ4qFXOdZJI/ClDfk+1rgQFouEchG1CToLo9+eZZGBvlbdVvQA
7sokdY5TCuUzc7iLETExkD6MJF5otTh0mqSAy70uCKtf8jKaZe2pmjCBIWyBYxQP
4OWEgPKBbeFz6QYoVhfImaz/uObn+vt0Uhbf0V9wEsr+DycKQjaO/UaxgwfPhHBw
0TXAe/T/QvpX8NsplBkqAtWsCPkiqFdjuIxZ9ID9OEKc9/U3QzHU5eQ1uGtPjInP
+rebM+aX5+eghgmTstQfr9GBfQGMlMY7WrmRP+6rgG04I6PG67+0XF9UCbrUQVDc
hDFNzHsFDwZWyOkCJ3QyrzZURZ93u6rw+XsXOQXWpfDmjkz0b41XASQStNdfhjq4
67Q+mFuld5zQY2voDe0dh9+tk9mDF8fP57/Wl3OYIN5T/Hz8tMAxd6wGXGqOx69z
E3aQy1kJiWCijzYZlY/f/Q/aNIAornIHGzaANWVHmgMHDYXYmscv9/60OK4humEq
LW7iM2YB5TpVnEanghrZ7Z3U+jr5JeL3DUdYuymki0kktbUDpUlLtQZ7KBZABFtX
XfMj5X+67NtkOCZtnGmm0+Uwa+YdGLJ1cdhbaVY3SFgeI9cmlr/V6oti1ez26T2k
FiUWEg6C5WoA4kyJJ1eRupUR32ZKZHQZxHkEC0qGbFxz+wmy+2dk3IAV79WQMcwf
EaFtijlcZ6R9zou43HcbbR7RBZfzEH8SApKoywWcydoQyjCaBa+Bm56TqCKJMdDy
EvvUn7lxtBjM8dxdylX53xTMxVdZOd66TYkbFWrYpNzHQY+mhoganJf7z7VsdOy5
uwW3uxJ/g8FSQRJX0r5MUmGwlQql8Ki2e0W8xUGHCbTrk+1ZunvFZuSVYzBi9WOz
L5DaMju0uLRKSeBWZ8anDlSxdoPrLgQvoch/gqjM/plPAP2P5h50vjXwo0D/qcXI
A+DvWEqyhWjUNDDRdiuoMOdy22WEZRSFUXYpSm+bfl/+5OV4q+g1FiSQdAevw+R/
uVqLu4LOabovBngxzfg026FTBJuzCoztsm92+3zHWKxvYh1ummrR1nFBeyE2CJgZ
BPsewXoI8sFe+HqrZ/xGjss8AYMoZC+6bDAyOmjdJEpS5f9/m5Dz9Kt+oLr8Ka1C
g7cPt0uZECL3hj8vDg0Yet1NdadIvMYclVdbbls8Rxp81u7UoxCg8f0qKMilY1t3
d4Fha6ORXn+g3UH21aNzT5/L9mdoMBMqpKgxOZ4pPmPNxd0fJw4lvtmbEbSSCC4p
18OsZkEHoCSV0xJ+pSLjYc/1yY1de70JcIA1KhzaIavZb+ZvoVz0VeujLMJHFjAj
WiX+nDJOJ5/EWmUbJmubL6KF9EGKNwYMb8XF9h8OEorUuv+8XeKdraBNqbxz19m0
kw1RoUskU4y3/eHIYy3ngs7ocSzPej0mzKEWMNEJP4l70B3TJb9YoYMbtvEkHm+k
XeZDbY7uw4St1aWT0mnbb9nikWrz9FcwbHUSBJIkT+16B8Xa1EVOiz1sPHjO2Hb/
dGoMO+RmUx+Uh8aaIspGN0/R2qhhvKoHgLJhklM97gknwyq5iNsszxrPnci4/wkT
X8igzZk2K4SyJ9i1NPqNIZSrDtVE0fff+hzHIwqkvwvQW6TDiDvqa4VxyZ1UD2iy
GoKQOqKP2QdWtU+hzLkKHsIpUOeUkiVD4DlJb/JXH+Z3OQReld6e4NwUSgPO6LbO
foxCdrGj49k7+0sI9kXyassjgg1a7AVALij42dLivRhrX6rFMjJq5Sn2G7mmQYt3
sdGCtP7jjKll5NkupzK021ucu3KtopU6lJ9ES315HH5ujHaPi9pkukEdVAwHTGZq
1+TdqYp2WovPyNOrUHx20W1BFCBU1sEY79rnBlsQ1b7djrHQZxlfW1zPqIjNlJkD
s1/C1pp8Q3oJ/D6/PVipouS0cPlt/BfxAkFA9uYXuFKnP98994K3mDs4660xstCn
nGTw86MgGCWRD6b0veJs8thAamyJcnLoSez2CZpxB9rF5oIH6wqJXr91vXto1nfx
jC0rO/R1qotBbTSP2VJi8c4UgS01DNhT45kMReBRs///qz3/m+rFR1SLl2wrVT08
lM2krVi+i8VsNrQnlLXirOQflHP6Y09LirEJDw5ps91NzkUe9AMaFcHpXquAIVjm
RP2auDGRMOR7ac3MFxmm7KxuneFJEVidjDHV1kq2UpysofIU1JkACWgGSGdE8rAT
U/egkLt0ZqfMJPq0tBxwqJSedSrC8hsyh0RT6e8DfQsFJx8lb/mQ0hpUqwr+2M5e
uaacc/OHQis1QlxyDDrd42THfGWPGfa5/deeHxbnoYCt4E2bjsfnMOpI0o1E/Llk
bOgHP+MyyyiXOfuU4Y7yTF9T7DDF1zPEcNRX6Ac7Q/4DbdmHtTyj526kPg55646a
FR3rlzmI1i2XoXeHZtWFGNaK4X3oGYZy9pTpgb4F4Gchzv1IN0LGlaz6j+jkjvnu
mSNhdLMw5RuaRy/MkTITStwqBxkcwJlfsG9/MMBiELYdeDTMHer2O+O4o+3jCVm5
Dtzdwv8dmReU2jI023m4CuUiUibptFz3wqY/eOrtn+JjVrTqhASov/32WIE4bAs8
l2IKCq80Rr4YV1Z3iwWokLSqrugylX5XzxGjmalEGGoUhqyyyK3TeLb2gQCbYxNM
7DN2CuUmMEosVXRg1riFL/2Pa3qmipwkWg8urYZLp3obrP9vNY6gbEmkKpd4AHLp
PMmiqOGKajm/pzNjSkh4+ZDZUCRHqsRaLt/KhhBng0LUje164YVXyzuSSZ7coHS2
rXnzzP+Ukw52kr1zVdmKcSm4/KG6DpK2+bikXkStcdypzLGL+vhtDi9vySb2ePMb
2c8DG22Tff055eVK02oDFANqroqM7PDjG3HZuiU/m1NwJkmnhjDR/bWlH6gCwKDF
6mFst32e7cNmW9xJzczizcwHXNEGk/Si8mAFpcU/Zm6WiSRB2qNt/32/fkvgMQtb
v7vXs+dvCRJrguxcKxntP2k8Bz7B9IrI4BfEt+u9BJJvXZjCQXoGaLbCbDxw1Wyl
/zgGgt2fQnckcTp+9GFX7HlDhpwSjXXbLWe9vyOcgQaJbk6xodfJTILUkDSQbtNS
z+Fq75mq+PmM/qUlL1mu6Qov/b5OOyTkJisoz68Fk2eAXbpiLN2JG4qxwfoWOAXI
YXMW199AgtWkjGAjlcznQir0M1eLOQc8R6qvoySitSVJqHobmabTZdFI6DsLC4Rd
JdzLe66qAJQB2CiK4El1Qg1D6IFK+kNtuRAbTfhPHJ2aWFe9KLpVW00qJVh8ZTHF
e4NDNajd14QUmA5ozuvHmUdmNZhb6DvG33k00aI1Vhcl+HIgPDuhXhtfbEcEW0ut
B89exxFKaW4+jMV4KMI0JD9QMvSqmYykAK8s/3p9fW7Dil7ZVhi3W/F2buLddJi1
O/AffuxWepHYnGWCR4tyVm4ku/GpE3b88fla4+NlzSpabUVKtkgEtFdZvD2HqH5I
G/SiTTe1kVngXIL04Fxflef3MM5TSCZlKSXGzUOGrCz+kt2CdHuP0KtBGQbPVqvm
I2dHJwb85RxWnNWHTsn/QeiE4hDRFQa1/6p0OvU5LnOQWHme2z9QBm9m62oZevow
fUPX9ZIVMYkl09cAhhu+iQVOkpX2Kd6M79YvGjSCH9VcM5MdxWo39paooFMfZwhv
mxaOyRvxhb6kSVsLhWty0kD3tK3cC9d3JKMWMUslv98SmqrKlGkG7lF6sFr7MIGv
6cWQ+2pUGyHaCfv60BCzQUBYoqled01q5jkcRjpnFEsV56wpM1tZkwjnW1L0aBJB
gRf+ENMWlETvLJS8B4nHuf4j1TSgDZ66YvOO0dHAmo3ASdmNQDmMlI6N/5rDoeNd
wLx4Z7kxj8CJ/jW/KVHcwkI9MChxGgSoFwvE+H6dlYhSI+rdoFZKrndNCR3EsjRq
KIAoloydAVFkLDfDOrM8bc6neRYMtV1ER/aETPJuZK4DItwFpBGd9Hady+SJY+oh
JF8bLZ9UkCXDMRxs9d0Ins8/57fwy0YjVFYXGtVDsF7voHZD7RktB0nN2B2aC0ek
uq7SUIKJYVuScIwfGm8LtapkgAHh+02JZjkXxVjOncHek+MDkH6DD/yZwzmF9jkY
TjFEu50dlNKF1rRO+yU0UCtZ2rEeBpjK5a0lzLXl//cPfpyOduHYeTaygW3wY9pa
0C3orjOYWDpTkAGswwCQOTu5hl8vcY9AV/zBcKYRiak1Zz9mb2PPMWnWQNBi/3v6
FG1zuYq03UE5DeWbDDA9doHPMhx9s0DGUxyeH0qLLW/KQ0c7PQGrnZoii82diVh6
TpYTD7IBWNXmmA67jvvDAAzHYDN1tmjOSo1lFl2196trrJrIJ8zuoZr3YUztzrSy
MEc5xbIXdT7jCrguNASxJoJv40YfVd3MSbgVLWczbQS8CjxSOX7+D57ZZxL4dVlq
qiU7X4OIrnKIV2i9cSxjTyWkqwDtvvwJ6IukGAwRd9WdY237xMY1HFy1mhhSDHJb
cxOiEiWOE/GsbuX2NJas7XBZqc4pMO+iUNW6rrkasfNIXN2uahB1eWlURWbvK2A+
Xutp36nK7OPuUOp5ywRCxmFDNhAKDlNtvQbqMkZUTnQHqjH4idc2yhRGA50OyLMf
lN8f5iS8rjmX9fFxMaUaYAxTryZlYcOmgbDb/loHEM1Ky4j2MgB5cKtJ2l1Ek6wh
872GupoJvKA2NeTkQbbXxZBUaJQ7/tBuIRWc+mwbgZ16CPbjZqVddHfp31+SpWwL
ClEJk2vD/yYft0fd5lLIibMGZDRktWaXupnaGx/pKKub3NO7o2dqb+Lux3pEYSj7
9AW/xH09N1NlIg3XlK4OrUe4Axpo3Wc2SKAzmoX1JjZJjurc9VZPcoAKIHUH+2F0
sC3cnEYFJtLkXhBAy9b5ykKQ7nGjOc9+RPud5QQ2TSr17cxUiKf2ZblFvaYrXQaH
X5uLU1DJpkdz9+6YWAcFe+hdYzKE/KZYp0k046tuLdoMAldwr5DsNvRbKVS1TgBX
Wep8El0YaweumBvyiE825wRObGX/h/GX067bkst5Y4C978Ssb1+N0Vc8jKZPoEXb
vVCuE535Jhii78GpojdkLWPq0gkhicWR9uSAez0nPQzwABUmqvWCZ0dsoR3anLoa
M2cYdZe+YR3aIctd19oijKXMZ5fPhUr4KpL8MBuI//o9bCxF4KpeYI/MQP0G2jyc
ehIoxQNZ82SLX1c5eIBl85g2gMe/hn2KVhX8/w1uMmKWIj9safwRAs04c9CRfqX5
5uPufp24VcDM6IcmpxK/iBnXuLwQf/Ox4TGjUWeB5rrmUY7OprgKyl0yWccSjIip
7ByX00V/xrpIk+oglrOx3hWm1LPAqZJ3nn3gl71MkwmZKq+LTvhCypBBVDN0HudE
nufriYD6NeLwP3Uh1OLtRFIu/XzUvfGccflQoTCmTk0QohAFQ+jZP2pORhzwq9fD
eDnuv3iUc0HRNT0qJRVYXVP21JVC8EUv8YOT8qXe7oW9z+xTdv54su9Uxv6tG88g
9HILTRioocuHn++rta6Aq6fS/+69R51VHnwIk7O+Oez2sZ5evrIAqatYQDdWCwSy
Lcz45H9QHxQnoeiAp3LZr2RCS6kXAMCRkWKm4M4XlcLAJSWSNfWNzYYT9cZHCDXe
KWMQyKDbJZsONJ34FvzSXe9mbELcHb91nT6C7Pmy0T01RZOoKizaS1ilUBYBMEWN
kyOeoA9zaP+DauiDwsMATNY0NTVWJjSSr7+atUYlmPZga7GitfSmS5F5/cYYkHdV
2KLAaJFb7wdO6CXVj3YWiX6wl+79zx+USej8qypOhf/yaOo0/Aj9eYOLi2v+zPvy
chs1jn6iGzca60y9okIaDmiYYuoaRsDg+uMJWS8Sx1HKJ5wbCwZsdKGDUk8w4Zze
NhtGnremDuzdSZHBX8F4dp0XIPFjzt6DEeXskE3yfAt8kS//knIJxiMrvq9h8bqI
3uL2ZUbkOYN9YWKzNX10Z720rHM7chusl5oJe6RxZESEHXR/qmMX0J/QCJbHsBKl
Q2mXr9muQ2tkUe10oygMXwOXqyUnFpbMdFrow4DCaK3soGiekdnqU+lxak//6ybW
mKBsTFRvcJa+0gZPxZIp0Av3oJdR6X6k4bl0P4rQPozy7U3lMJQkmBwg5LwMI9dD
/vSho52PawWX/qqduHLb3LLj3qX6u4xPVZBb2pAk8TH/ga+EN/kvujnXpgwdekd0
aufUd2cLsUjoKAt2ZfFG7+qpJQ7+mQvKiHnzhnilTjRH7BVEW6z3OdauNDPqrRl0
1DGLWFgSt04wh5nROPNnqzLNS9no3uchR9a2fBFjiPIc2pF6OLZhbc1m9mh7dSnX
93yYifR81HcHapAQo2eHQZ5+bju0vfbqOYPQnsVBOm6kJLVBKXt/f+rFWDQJvMob
JqZCiybLXB4eI7qtvYhC5YvoZkzdX2wVx/+CGgmDG6/myn6mgRiLeq60V7TCIDKn
erjkAK1+HMnFUkewhlOXxguegzQKF5tRGxPp6Y93CydgtGVx5k+89FDoc5/Zxyt+
+R1hts+jT48Pf9GrWCGmDZU7J8A6WTriq5SodNMFTH/PxwHXvEFax32ZSRQvnrjd
heQmqWLMqumGagVXftmZI2U/f52dfcUCVcG6I+tOMPjBWRwdXq6cEzv9TMeGbFUB
qxQwbrY4lAvDOhrHpfiKDZK7pZMFBsJI1gam/0Pi9tq64xcgn6/YJ1DnIDpN+2bA
VlcC+hRv25e8wRs4gBnZ0AK38FtkCP/l+srrA5Fe11rJaG8SDhml1xw3U+OTBI82
sYVQ/dOnntjvU+EMCY17jEPY6tniscv2iqHehwYyG/azYiXDbaGDAZMXa0hFZuhS
WXRicVR7i37Zy5ZK9CcOeMWwwxbh0S0gCq2T+XdoUlTij04AJSlQVj3uGiKREmiG
BFcZTRh8S/iiVpH1forP0a4KWl3Mt7Y5qKSW/88igTZPk9J/635wRy5MPHpLs7eW
xNLMW9wIet4azI+d1xQdSKOA2zezvGEtPTbPU0DAWXj+Onv2EsOBxO02NAFS0WoD
vOYbjjD1KopMTMY48uJi4eMxM94q3FNbdWqkr9s1KnpdVn2QYumsLelvlYY3ExNT
Lxx3Z63/6kUPNqRuKKjOJNggvgXHofbNdmM5bbqarBB3WeyX7KcLyTH47r4An46c
+i6/K5CHgvFmtaLxNNONB3Qr2Kj2gmlAp67XTv9k726FaDxKcWKULhj9keK4YeQO
n6ubq0Cth2tWJPU9VZRqeilYCNSW2evG6bYrwJTsmErtlj55u8SfRpgVUpA4qX2j
JCxBIow7GB13Zh/Z7TpjW5tBSEvJP4kQgcfYyqRuqMrbG7gaXwLsK3wpmhEpn0FL
Oy6UebLdSZwnhKmjCLLc2BoJGIx8U/75Q4H4AsYdkWciG2A8QtepT04bvZrTMND7
BbGiZJnx2H84SyVaT+uVRMPfFKvJqJOx6Fv5Psy6kKgSF1P00SliFYmbSbjbfGsw
G7brXJcqa9AIyJofsvD5wo64Qa8yna0FMJYAf6/W1YZjv3WbiXTMb0UZt0uxeml+
WB+P+cAcp6NGUSncNtNXXtsEGUHXnb3wvKWj4g3CL4PTFLkN3a8Q+i/TnSiGqSyj
t3CQccrQrHVoMmPSeRnswh41rxgs0aZC4m1gUVS+4URKV3DToG+TRvVgFDy35oH3
kzlDZBBrNEBXu2XewSxE3TagEW6kZzfAE6+LKW+Hq2ywHbpLr/x61SDeFeihtwdl
oN/8pFooN7iehoAAmhUVLZdDGcfz3dCFreeK0C1/p3eVxUmmjIqVEVYc7OHajmIe
8hyyLxACEFsRmvAHDF670DZM2q7LTmnWSkxr//KZokFo1jQXoeG+t7whvC3U6EBU
FdlRKHvTikYDNB6o2TPC/wpw5hh+RlVSXUXWKu79PY4nrW+vIN+3WjAVNJx9eEin
Qm3WRZu/5ALtmwrq3e8FInS9JJ0BuQ4WUn2CjH2FxXErbJKsNUVU1Sz5/zn9tegR
vxv6QqoU2WP8Jk4SrxjzaODkSv+qIP2y5P7SGHRqf10ODeKp7QhxaeHp4cQij+9r
+/EixDSyzxln7slZyaCUqxGajRtNMZke7cD2rDVbYcSxHoc5n3cPDI2V4MxEASI1
zqdBSeUmHIwtB4uq6kHRC3mlbLSQa5KOz0bjSNi35vYK6XnvWWtTGDn0WQ66Sthj
nUYHsjPgnlCmKnrle4dJAFmybhyNWwucZZtT1zpCW5g44/5nQklaH+MkQCHp6cfv
0Vm3gkqu0+rCHuiVjljaNdJzgsaxXuKUOm04PlXWekvKgPpwlCpO+P/4UdEUQX+m
Yhlc0qNwUGbRCu/JE2nf2jDHtZjNpLzNEeW0oXgDtvcwMwMOZbALv9vv/aVR8UVQ
uLi8oVU5yj436Rjz5yWgtSpgX9Nbtbb5ACI3WdyhpQJnmz+6WF7b+sFPQJqjJiNc
snaQdqTnbYtxChOykJheFklG8tjDhWhLR1ETqaaaHre+odtQZYadsKDYOdyLcoq0
y395HYbKFgpHI5NDPnfSXyr5yfmDJvcDSV3yrJjILfq2ADyw1eOtAenyhyCngvO1
rO9A8JsrnLY1aVrwXeaTCTUKQPrRyg1WJWs3j6MuYvQR/hcx0AIawPzq/CF3VwHj
8oETem73UqZ9lrPGSxe3SDpWa+Q/wggvQrIkwtZ7qK4roaxZQPSoaCehIjji/HCP
t//MpuygjQDtObB59wlhCVT2scySVkFfEkkpm2zQJg4hCC6OnE2iumWn/gtdldOt
r3wc5/haPPSyUC0CozMTmdI7V7490eUccM4oGWxfAnqGI3qeLWta1P0gdqfBPuNf
UllchePxGqGq/CqIng0QYKWDgGEicYxFQi1HFNxWcx1RB7iPpB/THSvUvBp1pPbA
jZVddIgI2QC4OSDBJbZF70Ja+JgPUGd5ItzDzLXe6U7SnE4hsesWRnPKcpKBjFu+
u66cO6elT409FXszz+k6w40WEz5dhfnLz055sGhm6tw/BfgZY8QKHGO9BkEsOavZ
M+gpHfYJbSzwNabOSxjN/HDCjJnJ6UjE0WIzwy0VFrGDL2+meRW8C51RzEfjLizr
H/0cAJrlSwWcjDRfC3Dw7KmviuSzAsWHLb4vW+9N6Ic8pvThyFExBlhAvu9WtdvC
6A1ALvl24fjhw7frqeungbh4EkBBQRPSX+45MTAg+dhp2CSKHHvbUvvNse3K9NdG
hbl0uXzQWUrqNymXTkVCahsqYsk2D17S0Oz4Mk8FJPnroWYxhHHI8fyyWn8yg2p7
O9tC2QVN+VjFUfA5xL88C8bDduB8ipYTmcJwjq8ZlAf6LuMONQhqcyitjh0uClVr
ATaBUt696cMBg3dGc0TbVQirAHCvSodDeynLF+tcZ19yNoSdI0W4NwHNrrquBNhS
i2WMvUREW5XZIJYNIVsqrErPfHAud8G6kAeR+lSNLHskxQCZwcrSomiw3QZbkloD
bqbfjIndsccuO/+yUHGhON+Gd5a+q9kPMJF9FlgvcBUjWVCNSnWRNnx1cqcU+4E+
VnMH6DYzCke+celoj1PDlfJLJYyQsTI17Nh+am689Cm9K8MTLhfyuQ7VsLt6mFSG
k0jxdQsyd/e5k3v/qsuPPd5+YUC15YmP3LHshXgmJhoIUUPd3K5+3aBw9Z3Ivvon
FbOS5aru4D1kcjNCSgfPuWAZoGItN78TZya0+7+73HJ+aAtBejtveIrGM3QRecJJ
PzaATiASS2gkHTUfWhyWW1HQ7gbAs0Z+CkwWJkNawUD1dIi5LddQcDG4nfZ9kv4M
iRVoMAYzFVhTM0wiQFVv5LdPixCLe2PwDLTs8xSmSSOqxoIZF0ChLquiSL7d/81i
Ufgi73ooJJFJqbY3QIs9ww8cLFWRjoDowco+kEENhR/pynPTYk8XUPGBAEsL9SMW
49cMOezq4p/3Ua7PBNLXbV+j8zy3k/b8fuWtw4em/MrM8FGyi2KYmued9i8moHA4
JzXWDzckvLHxPt56D1g0JCmEZp/6y3zx9YRZeQrVMfpAz68m5OAwnJ37/hvSb0LT
QiKzrzU1jvvl55b3MlSDIvDL7lvGHXD5A66frvkK0F2gTi7+LSg+k2/689joTH22
K5spbLTkepI9sWKd0hFURrS+H01+MebvwgTWDt+mtwtG7qOjxlvo05pY2NDTJjpk
oLfi52vFWgxLp74wqeakbZDYXj/muzT+UEAiN/clFxqLrbt8zYswQaGNoXq9tBZ0
PODGWKSz2o+MrpWSHqo6JSdxGL86HkLFUMJlI4pc4FLxBrYhnAyOPzcI1ecFHMlA
rFOT26lXSypPQ2WRd/bfso9p1boPXI/eGd6GetWEQ8x0KA0dBXRSk9OtZZmAkF8L
qVlwA8S09s4HLsL5eLc1KDu7jumOEQrif7eopdTL4IBwzHWUqQMfneEU31KiRw+P
qe8/HOpXSJZ2yqx9bsRH0jj6EW4iHQkdgpZBwCrSRIzk8tcFGG2SM70XQJNwDN9+
FVNVtX9O7TWyWXs4bxWw9R2zSGlU7VsolkSXuV4fcAkxmDapvhFZBEd6A6pJGDjz
nXW94kMTIscFOSdj72VQvYqPUh5OFwxLveOhv2rkfl2d5C3m0APtIkqOVmNkUyWp
S7zEyJ/UB3o3SjzsFIkiqc7332EMdwG35GQofkLdr0jeGMftQM93QfeLeh/GBWtA
oJ960/8Bs+ei5vRp6B+gMzaPZAW30gXCbAIRYprVviOV7VacZN6kk9vLzVLOQffc
zAKEId+sLpDE0/zQVUvpPqsG7RvIXDaVbqdpR82+Hb7n1loSlU/1CfUUnBG2DMk3
8L7f5nnRsGf8sci3+aFNbSxTPHKH4f8VXlPA277p/3IJPuyRZPntHtNkItRwQ8nw
ufxeHzmPIlbxGLkPYFskpDuRYA4vugfw1jTUt5DaaXb3XSqQUZwzcujHh71PJbG/
kROrMPMYz2gIIPtFCHRinXCg/tEmvcys+bmDS99ARZ7PF14vF2j5umGoNSWjAd1k
m9BFBsj5yq0zTb35/DeCFeuvXYh2luH1pPss/HLsQRGk23dnxkC6EoXvFiOxjHyS
W3rN5iqHwXnNLT1Kl+Pr1x7q1RRVBWDkXm6ymCQOAnmFgWXXQVCIpPg7igxog+hx
gGc3lh5DIUnjEBS3YAjvZ6EOl9aAZyELMvUxwKR7NEx6FDZZXXRp9KbJ0VUCac+S
5E+Ms2W54WEiIxxFt5uym27+q0JdSWjCIOVnPgFSZiSaRrSgXW1rvIVrKt3hX6Cy
si4CJnov+Jej1iAMqRK4CTeEBcMeCKvReh4qWc0a9WTJMYtFSNmttNQQd5neJ/eT
Jve/5jItMjNu6yKyhLqsV0bewafCw1dcmysJ4cdqkS8b5A6NtPtbP3/OMUftju3a
PLKSn1cIRJ4TfYlTgIDmbSDbc0m6Pk4ZqB1NqnqYX/pFyCSTLiMDyLG//pqYfkOB
Q3rpJgWGzymfM10LIuUl9ZTAnQpEvPYvADe6NSufRL7v71HAYZgMZq1M4BpRx+/O
0V8FCxtHsQE5Itt/PdDrG6R+gPmWLnOqVbHftLjXXoaorvcc2DnKqJ3zy5XRgHc7
DTzODV8yliau4/EiBu6EDc9kSMaaOSSWFBO8DFlrB2KrSq4YG0usZuaZ531G2pER
O2sQmF64r+Nv069MoRBuTPatqj9J+Rsv24aOv/CEm8tGjl6DmHr7JM0oCJXEBr4R
tzdMA+r8Zw5rMNk23LSD4KN0h8cmTUPkDm9WFwKCqy608iKrhg8bNKaTD0LG/W9Y
xvVwAoh8LU5NnMJdgRS6OhT8rw7wZwgMZgVkfBIn09VT9+aHfAjkJvGp3EEu7ZFO
hr7Etaz9LUT9k8JcK2KPUUYuGmmMJkaxJhVR7pqHRTaxRUH2RAa+Jy6Gn9TnIsyo
ZvjiIFRep2G2rdNTWDJ7fEZqPx8F3CXGISkxjghSAjfpclfjNGyMyC2SBa3fba7V
8Ff0CzBBgWb7z6rz4biBFIVKDwOVWzNNMM8pCQmvQVB14d1+sEB2uhamY6jyqcjL
NpkmqId33jfjFm71p2/Yh88XSiscxQlvYV4lvs4hmKg9Pn4cYxY8R/79dDyFzvLk
JMKSriqRt+2F5RB6hg0D59wWjHkJBTy0H0eLrs84uQNKwVUk6UJ0sXAvLCz+kh4i
dDcbwm+Wxn2rRdTEhe0SgpILfAViwC16uHDE6trdjQx7Fk2wOZLwIJMa35IqRyTX
TOKdtrvuXovQFr+4x11aa9gdHDkM9kenD0QuvwN6xexzRDg+apd9d+xnu/2TauSL
Ap344VpbbRC9d0zaa9wOG0sFgwRUp096JmiP/CaV7Rl6HFUEDr2eD4grGzCeHjiD
hr6NYnUXqbXLNtCpQG7rJXBv+B1Y660saln2txr+oLXROqFBKsPS1U+uSsziYAHU
gxR4l3tIpwRM49MoBQhd71Z2d0slUFo77jXtHk37Ces/3yw5BYRlHt0P9s+F1oPo
0WV+ai0Z0tq4uATqywC7hk3sz2XVcT4a9kmtZ/DAqQsWurtCQaH8aSoRwQ0NM627
UVL90BErI5qAkuA2BzVKHANybxM0T6jzmc+WUINLyFY7VNwjCp7mNxMtP44OcMY9
Qg0GJ3jLA5AJgVJdLq3nVIZQkCqF47pDjoeC9mDPusUTbWOwiX2fJD6cygjAaKyX
UGqo6t41Or8BGleqF7ics9L1gpI+U/3b8Wqls72+LGWWj/Oyz2q9ixbcPBQfN2Qy
pcA3jo3NBwKjjXKjzOHSGWYnHiVQ6Tp8pxV4PDRdTt9s6C9hk9r8eYqXA1G/r4Mo
xosrS1xuhpwEHaTnApL3tKxHnkbmKqnaUimhH5AQ//5asZAvU+knVEH+ZuK8Cvb0
s1R2f/H53YmgwzGB96aj3ICMVc4pwqaVP1SqvwZYE/UXUlrmkMXVKLOXBzZAKDBL
5WWBce2t/oSDQ/Thxzj1nUVUhJeLT05Jb+F0wZVk+cR5ZFwKSf/tl1Xo1WpCngNe
1w3qvqmJaJAbKp2BRj+FZPyMya9iSjfeKEiaz6JgA8eTryo4by4E8fjirAzFyzkh
ZmBkl2HjpDXCoTyIQWMa1Q7mI/2z/KbOi+ngnNEtzdX4Z9mmxrfPuDMg1R29qT41
1Zn8qVne25XmrYY8qGAFFjjHY/hUlgWmhpY17f0aabNs8FGoFfv/KedBGMAu4ZU4
e26nN7xLZ6LnbKUqDQM0iKc6UzwG+jJbGsu1tWgA5DPp0rL4fRi3Nnc9Dg9KQZw5
COha3DCi/jBF9Ds6Rb0BmpZn5g9OmSA1YufFP9CAdhqT6+pbdys4W5TKxLR+OEUT
QkhXAL5WNeSKqeflrbIuIZdAlkUaFVbdVmCGZ8CxGp1moWtx54Gew6W78fftifpN
CCYWl7jbWMY05nr3X3DykMQP++bfLTyAxzznP12GLewgJApJRlfaI9swyUeuo8Fp
qeJ6iJGY7GnNZ7NuaBFgr57LF0zHP+Omb5/zvVZzqJOlMLBM2atDSTH5jDcKEJzV
qaEMTj6c6+04QMQzizlzFD+A3bBm41oXCD11sTP3yKGP87qRTL28dP9a7svePU3x
/LYNqlUaUsweVNbD1H+Yv3W8OwUfobGieOmziTCTTyt9DUqoNK8MdM/WXZZEObBb
V1kd8XY/gRjnwJf7Gwv2KpLRzCSJ7uw2fbG54mthoo5Ne9wMX/vw4ThGeZicSlzG
ibqKV10uFGMChafuwYYU0zF0aKMgZ830QuOZVdNve40uggibZKjf3bd9E2hajbEU
NzaVdW5YRKvav/yc7rmO9p6YJ36c9cJp79J4ybW9gQCJq1M0mlN6Bffmpa5s9IYI
BnjbM8sOYLOdHymhb+WCaXr7dS4kCvwIPfvcVlK01ZccZasw73brZVU9aLWbcPsq
tqeI75Hq4li0DtP+FX8yYvlat+3TJl80TO4qh9xnnmmmEPXW8aCVpZB3soy5Z0xv
SeOgMFlt/mhUN6BXG/0lLF/yIl+XFp0rrGemStb1cnFyfBqAjudFVUkgvSB04kGJ
5V0DmGx0KC6Jyw3Pe4h9MFDKj3Q6plwW2WM+PMFzeMoWzLKl2qnEhqfkV40sKBFl
lO3rF6XL6zVOcpJyfJrdqdrE8dMekjEJiP/jwOM6pt6ZB/0AdrSMRDOr/FtVyuJ4
gujFE0Or4RlCqb3GdyoiGiqnsbv5fEJ2l5U04xjohReJHHm/vPkGs67ei6uh9No5
OzFWQriAtJCbQvlU/wH56Q8HZLwCDP4xAyIZEIGNFu5P8SRtqzB68k1rqLGXwIZh
PdoCiQGrChd1iCgAkuwbgRFfbZ5wjTFWYnoVFOYj3ufnH93VzmjT4pZwXYGj2RDn
uplf51ZCFoaPSFpw7m0T5RKTN86tkFQpyd7yCRCyC94tMPKQbeoGpUhyvrpmwCe0
bA/NjLNoZN58X0je2c3lhpXt7PgxkU8/FJ6DvIAqkh1R2pzCZ64R+5u7nADX3GeK
YXz2fbV7sbQ/n6LI4FK/wVbji6nnm545PzK2RQOSLIQcs9Fr6UEnPM1aFZJMO/Me
N0ZXrPSF6Te8j9MEVAmAbGJi2pS0pmE3Fqi3SnekGC+vREmMVNu6T5/vR21z31Pl
5y9W6uo72zl56q6okabwurKS12fU9igcbNN6RXTsnOuYdmnAH2MKP8HHUTXzzVmr
sonuXVeLb2vYw612K3ZI5zcMA4WoSAfEZPoIYqNtniLZ/Xd7UmRwPesjqjxs3vBw
QS3FFtabfWJnxH1rqSPTE+cv9o/lU9SoDZzA+QyTmd4z/hYl1s7DiJ4B+0UpTxID
G5M5Wuk18ChUZijiSf5HGlTOQMEaKtrvRd+ZHFsCtIQEDlh0bpvh5CL18hJqBd6s
M8rx0ceTFmBsh1UqGrE3YjMcfuodGr9q7eK4RNsYDkXa2kEndtce0GVycM1yH6oI
6spTKVp91008xbZzxElEhLoMkUkd6U4wcOw6kBzlsFgaNaLUgFdIVPrpXJvVrBSu
7vI+BfbAA9v3PEx04P0JfZPB7VeYWaynVRM6pMMTj4EAn5zJx7Ir1gD1d7XNuKH1
fEc8873V69B3jVqElfaCd3bfSwPeAF6RzkMsb+WDVooAiJI/w6pbFHV0WhvwDjR5
OtBYgB7FwlbkhpjLtBTbli017cQyYPFcnqjj+9ZPCD076FFIPkegsIsJIrPLYm/v
CK7KPoINwfGRVmEiLfTNt9Fe+d/ArqdMeEknNo4iZVPyFxDTJHk3s+Pnt3mdOACN
1tFGSkRi6E0KBcPLItwXm1Sz8zc+jjj7Vool6h/5IKoIArfG3vdaEd0rbv0BDxkq
Mpmw95MKDr/tODvwn/jplDfsRkyKFZsppw3487cLymLdUjcicJg9icFT9KvRhb8k
Vrlxl846bO4b8URmWyI8KrYlHrT4wfMatMC2aXWrvBkDu/LdFjmAtsmneTC3cCAP
TDp96YcdLbLbaKFAZOilXevXASzLjQqCuDc2fnTav7v3UAgqxyxsorwMhtMp+oDj
T9JkFsNqkHPMN6zE4N7mJstSWBpHznGIw4Sn25dbCbP1KdgTYVsxO8JQqdqY7rFY
bgvltD0T4eNAZKmHFAJpAiKGhUUyhJv2ooquUgOFsFk7tuaUxyjKIQBM5YOMaj3N
/zGPIyw6PW3WrSYqJSIul+kWZIy5dg7Hg4akt7kdGUSOjVbNyDyZgJJwUt+L3af8
HVhyD8YXI9b3saP0RmbS3W6m3CcMtmk9kVSZgS0JzLometgVFupyC240IbWrcVCO
oR6nLxgnRXFydc/Xwrt/3YYLqlTKMnaSBrKWZz+5xacLZkcE0d36TiY0rlidRYhR
bxgpMXQrbVPz+sVlJhhzTR+2orpycMYinnndNyhFxx8nchj0sdTGWTyGlPkOXqAK
6MZPsD1Q4n0uiTPzFxaFLahFrF/bJYiHwU8ed8ScEOm4uowof/4ByFR3uRHTQce3
ju7KZ1Y2Kw6Qjo8D4grGlTESb4qXPcMLt4zRWXJRZ7Sn9drLM3Nkx2IECSjTEQSh
6zQspn6if5dzpZTc0L23cDtclsNj10FpCxfflnylxXqq6K/d6fWGLdkHmbXLr3Iu
jOVyTor4EFBChzfcN6aDpHPm1NMg2S7yiJIrIud9zgm4UIAsQoTRh+XbPGOw9qSt
yFc4pzb3FBsw3YwF12CkCt0ZuLnqX4NC+ImuNeNGHYBFy69QPLDY1cdX6gi/uOcS
OT7W7buhjNv99X4xfTE56gq/fNhou3CUUEkk9LmceW1/4XRbfjgonxmavaHKGFJx
z2c5uIqsoGuFq6EsRBPKImATQdc5NZj9YtVBNzX2IZn83ZRfumLS/rP2NeseMMgL
69mLf10tG+sBx6WFkF8CWdUJpsmnEeJikHArZNm1sFoOiJoO5ZSG15JiumbCRGfv
rmn9WvEcBkD93FfFeCqjL6nl+TrprLqA52DR40pkQgsAmEPLOoK6fS3/zkU+blcB
yVBKsDk5Y31FBmfvDiX2a68q8VifCle31pegqIOUBiGlZf+Ai7oPoK8s35PgED96
2RSCUNBrBRY50DnXSnLnZ9iVnvcjGcB0nN4sk7MA2OwWFrHNoUjga4xRV+gfNGDx
XzcguQ9+UTLN5V0nwqtdaFxF0U/Gtl44sOGClLJpxC584yvIsT8W3guWTrkEgnEO
qFlDU548zv8GBXbvED9KlPUaiSl3k7keN1hWw7ft84qCioSo2i8CNtCEdiurxynJ
nju5Mh4yk7Kksux/P1shdFLrcmC2OWtO1eYfXZL2FBwwl9ee2K5YJm2a83fK1uNy
lILRdJyq7eXmx07TdkM34BKvHYinQ6XYN8mjESO+m1QLbOwBRdGDlU7JH4MugH8p
7OkDpugwEcsN3IsPZjg1PRXU8q25mJi/kFNDCmDTI5jNkhWNZUqCvyrXih3P6wuK
GGYndhGyfoitiocewTutmyFqv0wkfzLJvQRMf6CHWBNjeuEjX7HL++0vnjOrUpmg
fBXNpW339kVHv75L8WtvCmDqKCIag15hAcsvsWSYcMCOyw+R9kSB+bkv23fxvx9B
PM30UC4r8PNFG4zl5I2inUKSJXKz38m1vfF6mj6YbHQ/8myiFuh1ffI5qy8R5jsX
wxsGdY32dWC3LkiykXYEbbWb+ZJJ9MLGe9LS1TqMf9Dz+O6cNg9fMbRaO6IbcIFf
DQhiROToeOaVOgBqkjhd8RiJ/l/QzhyuFLw23+GuW57yPWX3AaRaH8zYk1+yoVQ+
hnzwZicMAfb9VJuL1+E78TFqbq+Bw2RTYH4FYougXk9pLYZ2VAvEZ4PALN3isZw9
+DU+DsTF/at6BiEEA9vFBGmGv+S/c6/g7K85/2xxISK03MJZqkbd3V/w4Y9ZCXxY
lXa7rWo9RfUxrdRWG+RKTH3aeT9hz9OHUuyjm2ntm9dYqLD9mkYESCchY175hbQ+
nE1/E+Ay+BJE9epfmB/uxRYb1b9uwnWQ0L0kBkSmxi5+yE3HfDZBt69GwZ5sU4uq
omC67vtHGdPafeYM7pO7agnWS1fN+p4Btpo/83e0j5C2kj3k6fvo6qTqK8m8adPO
EeFdC8knRLCAqzih3GacLTRn8gCCJOv4B70WX5dVeYR5X18dSe2nDR5lBsD5vhol
fh+tcgIZjsqhjNqEvSbxSaau4h3ss01BSpQ03x553atjZ8N5K/gXlGnbrFVItS7X
+EuXTl6sl4XjYHfwF2QBnUePwHEtSg1wZfdTnFZ02MnmJSSktjWqEBXNRVn6KLrY
ogxEIJmqitr94C2fLoyQJiz5vMIh+gwxIxAcUeTwjMy6Gk7u8n1sJRfDeuIxk0sq
ckC7ecJRihq4CzMYzL7Vst8q7SupCwdXjs01LUF0ryHHagq5v/gaYawXwkdeLvdw
RBuoseGxtiu7z6XrEGDBCTxYdJpU/7SanzH/BLcEhQOM1JEJr69He8oVIcfAhsfk
Sxm6DmIGfjfgbwR7Zkr6y9jrGQw0H5LNoCZaw8qISRZ3EsTQ+iCokvV2hcUiW+Kk
PkYgwQ3N8HpfGKOamY8QiggTEoOQnmDyNPOCIINFfDnpxJtMnEvUrLO1Dq4JrrGK
tJl2UPm9WCvqe/oHVdpk/Wf/bXFWe412jGIzjBDBoTBB10WBjQ3hcTOllPNHRKL7
31wZZblIzLsfsPv11PQz7Fn+vNokko+TN7OX26/+BzIVdiPcgGBXp9r6ElLf+Q6j
U6XmV3TIZi3nnzpl1pH7xKSVUJBBs5UW/7IRfift/CcYtV17ybmOyNeTU067B7wT
yzeqPtuCHwUryjhkWkGPQgpJb5X2sneV8BFZEJaVf5fZm6DATcTa7siCRTf7KJhZ
j3G0hrlFT9bO0xPTASaNgsXqX+WNQb1qtlUD4rFaUlBHmLttv9MAZxYlhntf7SX4
5c4Y0luZTclN/xoYM7CXOUQgQXJN5HG+M++ag3mb/FDfIgzSYTR5kb4XdbNsXCRN
mZORw4+M2SR8w19gxCMyzZLomVh2dbLBsuJ3ICcEUJGDhwjP882MipnFNgzqkJkJ
p6Hh/t34zeON7N8ewJ4TCMY/0zgFNXRIyec3lc8SNS/Rqm7UK1oHyJPZ5s592LBV
RMTYhAm8Gz08rOaJ4o/cspgnAh2LzLKTcX/MA079r/PdA6zf31kf/fcJbJihCo9B
bQn0gK65oVE5Mqzi0A3LZXzrBu2xTa/aQpgaJe2rxFFqw+RdH/tJQm0tikerQ2AP
jDIS34IYgIIOhEd0+a1Nn5yMNzVvXMyceAynTUEwKdWhT7Ms6KZ26R1UEC90Avps
0YhLcXsA4+ns7J4zTAtTOc2Qc/zVKOYdhtPWv4yyfakYWID4adCuXCEyldWHF11f
xcSlm2wuAirBwPQf3YymcOFt66e9MejWwL+Se3RwzNWCo2GolDpfeOfRjjJ/vIFQ
op4pFkgYf4PpBlSoKtQZkPMLqJKmdy9ru2EBgLhEZ4nTZdg52/dWt2iBUGG+sY1+
pSPv6gk/3mspgKDnsUjlVy4GneHb9VVGrjI8D/kswGYnbu88U9b1qPjY92mEPAgO
5+dEltB0SP1JNo2Cxpw4Y4fdxt017dQ47AXL1aSKezUIIS+Qrk2/oqUjd/lZCnGN
SPNivFdy5axtyVzYIWpaj3B9FMC/tAtUdvFu6WlfuRV3zN45NeJB2CsMb8rL+GS5
VwxI8uO5bEj49GlGCulCcvaQXbGRJCjC/gAuxLQFx+hkUFMUsxvEKJNwFxgRQ1hE
7TmXm7t0eklT3GPczff9H1dEYPsQHv9nSYJccB1DImenI9zBfQMzQoJlrTQZiANG
OWJsB6mX6UxoaWs9R32kRm2scjgGLL3L9HMk3TY6tlf6x80f4MWAobN4aTvpG0ox
J52YBqm1OnT/VOvX8ku69HMqPJSdKtSWsAZhWd1ueIEe7koHp81UWzOCXiFgd2HD
H5RA4vnzQ8b0gDjHaQLp/jY0oDjYVtiEOKOeOkU+0rWoewN/E8JW2JCmmOX88wg+
1GCLv/qlis2JCe4t6uPDRfB8NIqDt012JlrjI70cdj7U92hdPlAEFSCE0/tgj8dK
ZGuv18IMBJG8i1HK2DzXxfpfablJ4/301RQft9jPgvXGlIKp+xtk/Izitspq1bg1
HqI7Z8CuOgtuWfCOkoz5apwmEANTyNQYPO9ktgkffFVqHzD4UkKF/pfv4dWI+juB
I30sByAzN4FMeP3jPiQFIW22KJFXIIeqHRjUAPJd9Q1ig4z6cE/eIIexj2AvNCOn
WuUvilNe07euDuSid/vvrP1Jnc/RdkZwiFiBgEQpRE0SREQL0aN5pT4+USP/ek/H
7tk62JSLFz1NCb2sMGWW5QBYHjjjBbkJwWMpSeBoCSftpfmYp+oDOhcIoNcFfOit
AXKwAgTQVNxwm40FPCVfojaan3YQp08qJQYSQrE7zVhqxMwimkGzLEYQSh9xoKSi
XGX0Ha60xs2SMod7TSyq4PIXsGn2x7qo9Tq32q/3Nff5RS3ZYU/wAMfAFRgH8nxn
Ezs3aV7/jNrP5cCVC3gqpQHTZCB0cjDhEFsfxGfEsxVinddUO5MIyKe9BLJs5/us
OGGv/QDHLEU4Nc/BAfACDBflbT/kC/jKy0+4pOOLP1S1PC/2AhHW8YiEGx6JqqM9
w/HtfkzS6YdHfpzR5i1d310PXZ6EBf/OXlmh6N3EuYIFyf+WJWNIsivDvyvTxdhi
szM0gZhzS5xNr6austFK4NCByHjwoh9whsyY8guytxxSlXHdmcQ0KYDJK8VCDifi
0CTCON1TlSfR2nRyqloE79YSFbn4jI161ul7FM4NAeT/WwGeF95ljMFHH6wqTCpP
EBJAttGdfQO1BRuD8coWZbjC4GWZIS3/RwqQaNbLUXMIrmFGOBd0wiyGB1t0kPem
JeH8VTCOpHM/p7gtC+iiYDrj6FIluHrCtBexFMHA17dNXQolAO6s28n8FIaEenHq
G9E9d3da2nwrgz3Rg/u2dLqh314I+JR21bjJetuGMOYw7+gwX55hTDQBNaFVOwzR
+mvqNoEdwbn320VTftlfaPr9xtBcgKSHBVykXArigUZmobYDv6qp7mcSyMKlJpYg
fQ6+A2GzPzhe8RsmYEksJ2FuVznJA5aBh08eMf8vpw395Oc6Os6NX0eUo5sPQV8M
cblEkagdnXAWF0y/NHf8y1aLCDun1XUrd7JN3ehz0Gvr+dr9ddQsI+E9sY4KmPWJ
A4Iwg29aYnlpdKWrhZu1nquUMO+hs4hRimmow2ezdRHVvvQUoEzA/nZYqkcz9S8v
NNB3ypH39OfkwqDt+5AzAFn78GLVmKmnvkO2Fx30Dk8Vbh5CKZ+V9RvfEEJjZxf7
drHVL08ayK9ywRhwxf31bz49WFWaxrDeMWUGvWNU0wfxiDT4++P2xq/NFQW+P54b
VawZdtnB2g75IVBQ/XJKj0Y6/cJpJ51Qhacm9zW3hJVrNuwB4PjXXZNos1x3NUAj
yh+TxuXurp5j70h9FocgbmGo1Z6Ig7ob1ki00gOyVHLZzN310cP/UeSwfDW3j8es
U5fGCaPMq+8BlnwDK5/b/kk5O+3LDIXNFCWYYr0bIx+s2e93sxRWJ7POOBmGVuN7
/Fi+Yslg7Q9WM6/T8JDeA990ai5KG5/J1WgyFGISohZYUWnZorDV6MJXS7e6uoG3
f4kzzGGg43QI6rCkJ6DVceY5aDm9v7IOIQo7xQ3CVtpQAzAJ91zdU8KbDXt4qACf
PN2JDMJPcG+u0B/xbd+MRMnwOsNCzmYm3YPYuIqOXYLb6ysHsFBak2WBShN6VzDr
c8Lt57+Ydd8V8XHHVceJM2yEUno6ObbUc8rwex1/EDQ8lbSm4dVZrO5f/vnQN9kI
UF7Zl3bTk+eW9tO8tPLmUj9Jv2nf0G5iuPW2WmsXb6CIcuGFKiM1yz6WJY4M0OOR
zWUPkFaRkvDvn9lpk9tuZct3iMr6XmRz95fAB/GObvtkxKRLjOyTOIY2qETXv3t/
P/vTr8blMR4p/bv3ML8jmXY7SdXwkZvwU7BIbikElOJjBcj2PSi4kNPOV71oMIMA
YAiLCPLX4+Hvy2njXhVsZpfKZS9thrO9j/Nzz1kSC8sxNuwducZaTe9XnyVDJiKu
CPYZdXEbEtqyg4zLQUGtLWQJRzSVuweOWHIIWgI+NGen4kiwSGpWqYr0zQhpzj5S
ZHdHOi/OrZtVIKjZ/ZH+X4vzVgtgyNnbzUMK2VTko5qlg3JquA+pnDEMlhWq33Wc
IOfuDFRUhrjb6oPPE1LVLNN6keBWCfRvcsjfdmEuyaftsn3b0jHZ7cs1Y4AQwN7T
Umr8qfHiLf+Ri/UmK+qBzlHjh+D5yKXVPXCvLp14B42EfBPirgAPQlksLnD3XbwG
9XBjGqwzlIHf8tDAD/V1rdvo3YHLUiSvILa7RgtfFpYAW9wnV2jRF1/PxMGYA4Rt
Ogp/oHO001cTkkUvQ4JmfWdMtKz/Ks5Z9X5zkchb6s6Kst78POCGX+5z5k146BWP
A7dm3PpowFaMC2nzX3DRSrVQJCg2gY6/vvMNF2YIN6YHe+Df5HiTXWWRSHr54X8P
jDrc5ErinP3DrGI6nRbwiHUT9txm48KXLfLGrc/z12Rp6Wf2LSfh7m7IHujrVq5y
d5qdghQANL3l7JJImamtL9qkEBWO9TqQfnP44eXtyjjutyUGRunhD6vh/obUrc7u
F/fmluF74cPFItrIiglFmRMWcqt7ZNR59u52CIORZ7b4LCRElpT6jtyk2Inv2Ygm
/N6FHOMpheKIF3xiJyqS+yZTVF1veOaNCQi6QZysGKd2lrVmt+oMItW2PvLlC9Ag
IlHoegD3cAgEu2uP93kIY4dewZ5iHudxFderDsttgxdAIhrzDTpJrF1hQbsl2FKM
k7rpberGjugo98wfMQC8II4Gji/7HyM3h3DlIxAUWKBZYEYEXfOdvo7d8lHUDcwM
OMrLR/VAZa+6fSc/yCLNPLc5Q23FHsYiKa5xe+DNGvPXzsuAH81Lmqvi/6E1+gAN
WQx9TxfbJxPH+jfRDG5PNjW3WAxcUWlhl0dhVktqQVoik/aZodrQwkHFiecbVYzc
C0oXzTCNzWgy/MqC+2Lb5ACIJ9fBY+fBYDUflFRDduTC6nAv1UkuCFxMJq8ssqop
hItpGX3ovHjbenf7Nv3u5ER4O6Kh3iuTk76Ew3QKDoa5mylfQsO3CA8PP/XCmvsJ
Uti+Rc5zAYyRJrZdn0ykAlAWK2botiSKyLxPekXPRt5gbEnNVC0CSAHZmSzM4keF
7MNEzUG/lty+uT20U9BGEzsnqMX6Dx+L5PeeqfwJ5eTTCFQY7hiX6vIOBOODJBoT
lKqGs0ZMk20MmvLWsHX6Uqua2WQnwypkgY8hiJ605uKrABvcEQ0t7kPhRV5bL/4p
4DbKAVCrs7ICzLuk6ECncXdBI5XPZBoziKN9gBynaro120e0hzHZ59CL7WwYtVX/
2drpSY0sdCRUB59RUNFtD0y8zbBdkVS2qThLRmH0DGk7dm+CzRIy/klXlMKOp09d
bFyljKDNdkgbblLrEmCkbXGyq3cEH/uk4DkpR1tb+iUF6Z978t3fCDr4BsBGihGW
txcDkg+WN0xpmWEwqrV5JZNCq5kkPFidcqb0AvrsQFm9C5asCGBHhCgBw62fIa6y
GOd5PHQ2WHbQItQ3Fo8nyI96wGxBCbBFG3h3HbZkeAiDUT5Ce5NTuZS9/RTLxt2p
LDS+YdA7txWbJC7Qt/duWdj4Um/CR/XaAh+Psx3ba8QJNp6NR7MqVtNxLj3dN5J1
7yVRQFemP6wLPa3tgLTRmKaQkLHElI5LJWO4/CiDHf9YG3t9JiFuTMIwDnKYvKIV
dWPJAKxH2CriyIbmWyOSM6mrJq5xRerPS1RoYB/bHXLjwv5tHgoknuna6lax3cAw
gy1r+FasMInfqkFSmO4EbS+LRO6Og9vQkChO0ZJuCP4sa7kTsW1E1VGj2rbSTcJD
z16GtG7LOyLRVyDlp+R3M+SLUekF+UyxxlIASSpb9bpuvQ3Gj1x/hvREbKSvWPYa
zKlxlVLCrqryAJnl18K3lBmJOmE0zSO7Comjdp/uxkVMq2vIHSI1AAAFYYJJM2JK
OY/V3AQLpvMPCjfS2fY7nH/6Ii4EhblhPleuvofb6W6w212olOfjyweLZeDRIs2D
lKpMY312qo/UHDB2RzzcaMuIkbg7ZsEAdau4YvCc3de5/cipb6XgtIsLU1vBV297
OTyoZ0+GhWMDwo0iDCP2fBa2AW+iiIlfMXZ88NyDc6p9cMSk0hnPHjpN+AojzhzX
k5YhQhREq68Vpnq0qggfKMaGd1AOYZg9D8RVRVPYfMnOduqX2FjTpiQyBTEvO85R
DFjKvX5UX/PJM/Qsb6pdwgRVgNP/e1crNUs3vKmo/qI3t73qCeSrUM+rYQJomW/9
uOs+ifbKL6UHGICutTEGGzXp7EPosKjVpXW1o7q1mHN4QELx/3+vaM27Uv4yY0PV
hIEl+DeZt5ilLsub1swf0l52VJBgODJjyhabDoa7hWvpewmdll4YQXUgHRrhlcvH
Tqw+LWk6q0ClLnufX01ALDLDW99DNkuefLG1kvQ/hdA4fADP7jd7RHbRznFLAjHz
3HyKN1M7VoWGP0f7TZ9pPvG16chFySbGPwcZUs3Kj+eowr84Mk5n1bw8+X6LP0E6
xXCoikSOjgnVZscspw6K8StGwlL0uG3kgr9xzRgT+KJEnGDLVjcmb1kSWwbl+iSY
NzAv/nceKKTWQnaXSrUm6O5gBvLz6/Gb2ie1Qwn/HEYMO7RLcTd193gczOVye26K
zlVqxrSRdPBakkZvCNl5ClqRTT77PZ77wGdGk/8g4arlCSyxBJ53XDdZXiLzrSQ+
WLE9b5xdlFQcAiK0uNy0D91/KRokHeLXVyevJhvo4VJiJV2vjW5YGP/w9L3tofag
wdAUnYSTp1d1Ku6HN2l4gyYg4m9uM5MmzLdfGLqsX/AYv7vXpk5aur55OiqRxdtz
I5WpDl+5N+b+Nlore7mNijA2OI3+DtaRxHIOWw0n/+ecolO0a4zSljGlCPmwJ/vb
I4KvUYx+J4iqzAOXtzn/PA4dcXtFEpTtUFVDB7IeAADZ9X+e0riPYbogijZhb6Nv
ULLw62UZgQWFrU8r1rkulumpKP1yVBLng8AE650QjQJF8SmQo/mhmtl9ifWGWViL
aISYBuD4GbW7DBSMV72zAwUSZOxPrUgre+ME596zE00A1RvfESVePPF+bxfG5ULe
nqeF3qM+mg6TDMW6i0jZznrv5Fak3O4ZUnMUG+zvSHgYGCJQyXMaCpnnof8bKYGL
6buRKEX+wTfdgYLM7JKZp0o9mQcL6cwwzdEC2ONxquQHqCVrxPog8U493vaGqH1c
TTv+Zqi7nw5Zyg5ZOOqhzFHo3cwKFfyWhSfrDhh32ID+7zOLv7y6HW5v0ll27zby
lO0t9iSJ+9gIexXIPP+thYjFvci1supSD/cckPWaBFKB0AAQM8UUlmhfvocC9DvJ
xWVXs7stXi0XSKNuVMB3moVu60fhGpfQZGeDnsSqkVQtYfMA0golPFP6cwxTd5b5
XMeylOalPQ4yiomS4gcYugRD1ibZ+jjYtSqaAPp/2Mv07bPRWUg2uQv0/glAzBEc
Ts2u+ZSTxvSvq383h155KweucbJzM1jii5TbNUouf+91AREh3Szd1bWvBrrW1yne
CqUXms4rxh/tQeFGu/7bzwcSbJH2px4STSjd+YALiq85j6wMQVxdlnmpeZeb+DgD
XlLrCyKpxeVU2yPbBPmvSOzSG+NjDXBJ5YMwYenCKjXgdXtzmkCx35Qab0e4mIE9
KF69XAqKrDavKBcTIpL/OZxswpVVVlUaKFNMfeEeDCVv/bBMvlA2wUaQoBiOf0Zx
vorZAOvi3iw9nmnel7dhniTqH3B67gc3JzE+mfth/FlTsA6qIshP5dCf6Hk3PAZA
GohxA4m61Risfe+cxLks1w7pCLUilgf+44nptPHxpUI9B18+G+4vgCoaiHCuNHtF
UYflf6z08X/oDVtbl94PjPjsBgKzeIj5pJdhzFDfyaUYU/yeVCe63B3Ntw+Opd6E
ddiSHMTt6ceGEpy+VyAsPdt+bvPbaFzQyyQMQQFWbfq2cuz2FhRzb8eOCNOqOYTh
Gb9QOpUiMUIMq3o+2NbdeSjwc0iZquI9YdorP4F5WH9r1aXXKmfUmQzIPYG+D35+
zbahccnviojCGNyE9Wj80uZWOrAEX9pVdi2BDhhmHmStU2vZkVmh3UGncgRY3gAr
ReXqmI4vvl92aavoCOPWWhdcSdDjbj+pHA+VoJmH1lw7KUlpWJ405n69EUQFz2ps
eYfSZzyPNxpw/8RHe0GxBjnJ1s7hgKP4reQiFpErO7RYFQH3yvEf0U10c2qAD7UN
hRcM5KqmJzv1H5QmVDm3YUxzQ1PkevRmch0vS8AEops5ZA4jtROkOAZIgAeuVCj9
vRrkIvZAUezvM2kyaA81N6cZysSssPum9rQIujvJlE20AxxFsv5WJPeQVSyGg0Ha
HuSPovRRs7rFwQHjlUq3R9nmobU8AFHDmm2czvyJ5CHXekTE9mqCr9WP3xjcc3kA
9BHu5sbt1Meh+dmqbPiaVsinL2Glm1DHy2FFH+PasSu4L88Ng+Yr1bhuOfz2T7ts
k9+zjKPoNmMvHECcAYIw87tvz1VpF088YaPR9HspH6er0oPpR0NBxhLP2C33wQTO
4MybjoZ8VSDzF9I09wywBeRgnGJcgUB10tiQ6fNHZYWLZKpn8OyVzuNcago++J5x
ebuwMe+m7s9jR3haCFnAKzH1gK1E4tZ2kJo3luwnWBvNGx3awIKTEwMjVz83pqyR
ayKCnx0UhKwnIrwutB4lzwx2+a9yymHX0tIX9SxJVXMTXhmQBFTNabs7de0MVZPD
NZtpHJgRKOaUPYbVid9mMmtVdRsK0Ac5fRlxTAPbfkfnqgrW/eV+XNeW/wESRdZ8
xDMI0HC36Lgd5MqfAZv/CniJDykpCpE+eo4yye/XAxT2A9+FkJofYFLdICkVbJkF
DTMZNI/IYslO6BcuOd6/KI3ZshsyySdcsOPmwAcZDiWHL4uThQrmTBbDW2apdmXV
ErocIWZQ2f41PtyJioRAUj4fxvDMfMv04UnVhyaRig6iwANXPK7z6/rpAex12w4b
qM53sBUxQd037nlYysW1ACDNdHLovXP9s5YvjdVri4xHWhebQm0nzzeLXGtyRgym
D1dx7/2jVSBOK5uJJfeWbGb6FDdKyNyteQV4Y97H3WtV8k5MkQbYTplYu4l3Zvli
7GxXXD3+8iNOcV010ZqeVzlbL7CEpM0OsTDqCALYvOutTcnuxIevs1QwVpukO85M
jr91ibyhHlWg4ffNalCtbFGJAq6Lgix7SppPTeSzMiGOicdwOKee4JGJQNsBDTtt
0TW/R4Ut3Pc39CC11l9iuQinKLIEQFcxtHfn+dBtJdrzyPxN2OA6xrW3ygNtAxfy
Oz6H/0JfvNNpls78DyydQ7qnlwX/6JJDlYENGZWOp9WbVuK5Xyx727jMOgoVkkTr
g4tBTAt6Z0mA2g5VWcDYZRcQPHOswubbwVfnhdXPaMi5W8SZZ23gbFbxuOCBsSe9
DTQKSBs/3wXHk2aYUx5qmvof/WtLRbK0CBptj6bvFslsaUyS+9W8CT9bFFt3cJVf
5u18MvFDZ7tBCFCNe+pu7jZzALJE3tswNKNJcBqfngPddvjOUTgBpVQlQ7oq3aVG
pHZXAu0iPP4F1tIR0rozkJZf2KJeMyVQB+Uf9ZT2DxHWfoc4jShraZmuIh8UJ1Ad
Y8/LfMaRd/C6DhV3oQS0RQjoTQ9KAe2qT7VKKDs7xIjhHhAeoii3vYuKeNNZv5Cf
ZHtH6hVdneoVk5J8niaUoFX5Fd9zHlmhVXn4xFjn/CBCLtlOcEMRBDlbGDBoLxCt
s9SjTybv6gfhKjyi4VaRxHTbYOANxjXDL9WgSEe3GDB/A4ma9WOH6gudFlv5iJ+k
ePZ6bOQfwk9VDUx5C8quRIBpnQxgbQw3VUn21Cfq0hB6QJVNUzw/MrmSaH3WvDV9
mXNjTjy2crODWjlX2sI0SvvdCukBytZdOLchkm5s4MNaINdJuSnWJEnxAg1CQUhU
+UI+htAJYSHjTXqjY+LpRqliUYyftK6LBxq28hT7ZaQ/SfGhuR7kYOobBm0ZMK1G
hvgKwc8VGHe3wp+NJqO0Zt9UUR2FXM87o1OPnUh5glXvy1pTucRZjEat02ZUa/hi
UjUMVcxZphcArHR5EsA3BzJroL29FOb430CMs++LgawxSwnSoPjwyoi2SoeLwiI7
GYr8IGmyPqLQs28vzGIDxHXg3ftgWQ1H2DC2xFRKmS4PpGlY2axKSnN9g40zOAe8
vE7IFmoKjVHcAW4ujO251vqCrkqfUr+r9mBKxy2z7NyXo0wCBh2kRSHg94TvUlzb
iHXbTf8Z4zv/C6rNBsNbSGIelKN7oseTKFXbICsXnVMmu5IH+eZY8pR/+BoGALO6
jWibPZakaJhM/84O2v7XFAL7NoLdMQxItEsimPTzvCcBo226fiOG54YlehtgFRos
lQB8DJvsD85mTZ5tmwpUUfx5Xy+3HICUq2qugUifLIjL03wKmxlEW9gnmG9B9+v7
Tf5yHNILIepgzvzrjjjdjzWvTLFvxOJ7y+Lf7zOqh60Jc32zNYDLE0S8yajhLaK5
hbs+sfJs2NvqRyLKMfgiXIS8GSR/xUuht/wuhzEgNzJro8UdhrBLhoTi6muAcDDO
xCRuS3GUx5UQGY39A2P6o+zokV+pimZyiMhURaSKbvbVX+rUcSYKDqYLhICOw6AC
lCwFhzrDoJmeyW5bHGAo4F54/KhknD3z22YfQdyIRJNjoYyF5gCGgfM6PDL+4unH
w6Qka9vpreL8vOB6SmJCjcAbKitHZz3CymP3IDGa1e4laqzEH+r/SsXVqnxXerbA
DLVqwHm//FBDxLjKoykUePgzFSbciXQYJrWS+mmFVR9xqEPyA2wYR8P5sHrsOe7w
jEOZX5ZQyn0b0nXFwphUMfndVFMzH1tyTQjak1bbo8nwN+xvnGDoTMbCHZpoWYXb
HEK+DD8Es9YQWxfTgFpDRzygfymqtLiXTWUt2jVfmlFxa0HhMTaMoTFBknD1eM1j
5LVfnYZukIuxq/ksrDOlXau4UfUOp4BPIy2ILbFPGcJkqcefYuU3A9F6RQ9YDlCs
tMR3DC4MS0OkHfyD+9jlqh0tKWsm8X+bH5JE/dkFzXwoWPPacgUzbUuo1DgbeqfU
1JA39mk9iEdCCBQiFlYok1m1rMtNwhyTjTlw8K3om+RYmnbxH9o/smmUW4HWfMW8
QwPiodPQ4dNp+Oq9LNAttG/Pf/5z0OeajvMobxdiENnvT+502UZDhI3AYzHfJHjx
VaRy9/C9JqjgUSbOhb6jk7Pingje7aZfn3yjhRF7j11UNiI2rky35BRYtjajw407
J2roSjPYIDwS/WDHheONyWeU2raeyEi9uUQ7M14BhVPvfVw3gQ3bcteuGfym2xYt
luqxsxhg/x+kpQm5XTmwPobnZwcOEQoW2BMiPGjh7jz15njI6sJ1GEb1szFgGw9S
VN0D9W1ExpecHMQzryDIUuaCOznYudBLUNknWCrevRKX9ua/K66ozQikp+Si3/AT
6pCeQOTzrRSjUcr+TrFmWQtn5kn4ZKwEIT5eL4XEahL/xxnuSj8u5sBXNIfW6lh8
q9lD8SQ2dqJoUS3otqw2oNUs8cU5Eol2xIT1a806ZPU4EBPR2PZuHwEIf4IyjJ1N
ZntVyXVmqY7Ac0eOuz+txoKpHnPOcn8vGQal/ecPVOhoqcj/ZUVSN6SFxuxSVjr5
bBuBHJZ93gdfGw/UIl72MB566v1vP9jlVl7KGXP9OX+dTHzNzjPilG6p0Eyjh3QU
9rfcpPxINOv07Bl4ldPuXPd+5FCo4YSavlaTFhzfriuq+7F6cFVvQERl4lHYV42C
iIte30fbhwzpG+4iTRlQr9iwYbKz7inUenJMbBhHa6HkRaSHMys0kHogbQtMIszV
r9usVFXy8rJEztd8u2L24u+jy5isEm5s6jHo5ErB/eMKz1CgtNyaYcRnUIrNOoUD
Y/45v8wgWXQoa9MR469YsIxBSLkIwegpXr8XxpWG8rLaG4NOyo/o61xFWTsNW5kl
P6chpxN2f+b/kQ13rocdUnQgyxUuf6/50dhvOHC8uvx3JEkBOLOXeHE/u7+bREFN
g93TAvhVF5OSEdf4pdLqnPHb5JbpwIHnItK10Fv6ohLMaPwFmEKeT5vwG25NN3li
HBeANrp7eKXLUQVl7gd6HoGnFPUHIPB19kdkyKT/BJ4gSMZEI6/zU97w5EaAXTEd
gIJr6aQ5EHu8TXUnxevKMg9oHZlJjXIG/X1F6fcyaAmGMhZGwYVnOrPFfT+UPTKQ
17XeY52uTG+5ggC0RVYjcvrEfgaE75tYTwDyRAfnJX1xUGOWEoaypDmcfFhUVeIC
JMYrNWyG1aoBiaIJJez/fTg8HhVs3DMjGeSoC3//NVP9/4L0OyiuCWDhWawpTnZo
Tf8h5cU10C2vYOIyWjpUHT8uPhexV8fr1FYZnam51skiLAnVrQCXNnaPYP9Qgshy
YWzA7ehDBL/A0KXcgINmdP5Ff6Q6fkY9d70g01MYSS61ajBp6cgaZaafPSHPwbEL
F1OhUli3RTGFoIej53VAcu+qIOv/MBrrUKpViKmpSJvywPC0twN+UElFMqfAvF6D
/MgROUPUWxGK0szpm0BhnR95TIDJ1Up3BXagPo6nq1S3LKTWkqC4rkk2F++AQ7mZ
IiJqxdAumxstz5biCTcqg3tZhjLut60so0tSmiB5t1bBUBjcN8noY/gYEFqDjyi2
2E/te8Y7ITQWHiTDnwnaYqVhqQX1lFg3UTTJiKJxloxFBRw7ckzJ8nY4eA0M65B7
MEzDaiVzAB2lvMSKij7WJW7xqmpCqFNQVNgbbKFjZEn+XmAs55xREutTLuetxQJh
nH/9Mt6LiEzG+7WHd+FCGhHYaEDzF4jMZv3PELGPcgtZxzw6z3xy9Rm77bmN/pEE
NnKqPqTJSAyLkVRfrmdStihgJ+zNTIXr3uN72u0hoV0SzEtnlD9mpsFQcVIBRnGC
U2zo3lSCY/RhivJeMt/t7H4yGusMW/vdffgQcBBYKhbjbJ84JXX6UOzWwkTWY6up
7OWiNB2PVRizOTB1tA9QYUri8GW85bJkZ1flpVC33xuoi0z2yUMAaEpYM9kl+ZrH
cFr1m0HvHbrEDUH+1OZzDxJSO0KnA7bCrxJpDFqCUQSbo0U4ZfEDP6ehrqQBDuoa
HfqTNcZxYZ8ir6gkDIMCkf80YVyJGVKTL9RLS1beFKPB9C+CmGQ6AjVtwKt+XbbR
Cy1ejB1CyONbt/k+uLw96r2bsB5augGTISJEFimFl2otaGop2dCFOz+1FwUvgwuj
OdICHy5i2z2jPPpX/VLOq0j4bG0i5ovuXtZ32Pr1AegjhsQLC8QanG/m2n7uwsPn
GvgEJsQvuKQmYTH12B358CY9b+DroEJnZzOhBl2rW0ga75Lg4uAP9XKWtCGCYROK
dPhQ3B3G3qNL4uFVgZxNJTZKyyqYMH4v6qWYYMpeWdj/g01kBZ+AmYE+0dRO0+5m
KEmd7QQz81k0v1DkUBQwfTuzsktlm8eoHrKeURr5dRdjlGL4BlA0G7MgUQm2dQVL
nIFxRXI+RiTzcLYr6Pg887BYc/hCQRK5yKo9CqThLitHKgekKH6XZwUv9+WzOxC5
dyU2wRFql3vG+1NlDI2ND92vrAnOh3PrxXUM34t9rahkRgcw5irL3PBjgYDa6KRu
zw7z7uHhES15TEk1syiji77qmmwAvCg1OqMad8SajKrur4Ha3q2aspyGe6I9Fb1M
8NclrF8S9D6AzvMULExTDwnccG5ET36KZJ/YPOGGPjRxu5J1BI7TPvlwX+TfC5+O
4+jy7IL7HMcSrkhCArwwD4oUpa0Y1doogablb9rst2wB/foUv8NiXwa4C+X4nRNO
UNyrJ897FTkmTI6Rz8QsOUILoV4qHOqQiV5amEKczWdp4ow/M2IvxabgzboE5oeZ
IzXDxuGiV2/aa6qM/XLLw+oAgHdRSkCweU4gLrNQR4GxasddpjSxwt1jiquKuxed
e8dc8Xr7svXbpmSMivUFetx7xsMKKQKZ0ufLCP+0beMW23yhxLGNnm2IWsqOEVUC
tkM6eOM0qILsQfaPnT0RT7JndkhaShpGa2SrGu91GrYDPLakvbnciQweBjX+B/su
qbQM0GNE2LADdCHNq7Y2NtHRfoj3dHlLsT4wdddvw58vZT5XK+6HjH9T/ULRKRyM
0rnp0W9FauuqFcSh+cOF4auxlcavjNK8jRDqIWIHeDgaepxSJDgz9CuKQFvLZ3DR
DW/uqjTOE6CjVvPNX7+T3iC0VXJy/dHB7Qx4r6KPA2Hy0HmeKgJSlOvx4BEYYrcO
S6XM1jSoR7DYy5ATtvmMbrj7BpbyUtLq1jrv5UwhICfxoljnOJGHx2kcAt8hZPtM
pDCVy0wz8h03kGXj8ZfOrrKYBDPoijilDcC57XQ85YOxJWfNybX38sjGfwkDm4iN
zEtSwvwvEnVF/MERaX+T36x0LlsRc0smDa3ZLfzDq00A0WsjxroyjWk+jw8wyfWu
iuo8Z8iN5njtt2nnU43WA7sKYjaXy5tPU/vDcsZNElKxbdOPk+tMFY41NihNrWuy
3iksGN8x8h99dIa9Ou7SQ59+6oJYTwwFH8QzQf2xy3JVi50k66v3wOwyesNnkoTz
eVs3g9Eg3bEuFJEfag/Ln/YZuZqLRxNiG1yz/vJpAC/sqcgYKgwvhnLe2wm9sGjh
z9vfXmUMALbe99UqglHhBz9y1UywB7ILhYzQdwL70yjAYPF72L4TM+AOzj3M2TIj
4Z7g9yZFzg0UbgCizwiTrqzO6zucn2ntPa8lUXH4+7FHBWggEozBrfkdVjh0qKyh
2VWd26MlVX8LMunhpp4apGSFcOF6zj5WP1AFOZhRnYwi/4767FG5t2LV0fIazKfN
l5lZFkm233t5qWoPSfxhV0fgps3xQeSMSLQK+pdANne8nZH9sNH7aJPuL5tEWDas
xYTZAr0BhXTh1ppemPjhnCfRjXwR0gulSNrGbI8v5gacB2P56Cis/Z/WdPqZyDhI
xgxROOJ9o6J6NJlaPrW5cNeXmI0GBRjDRI4aJxmvLG16KRLljMVCpiYef1XeUwRY
2VWmabZABuihqI27USowpmJO24SGxb3uS0C6F1XZLepRlQm9pwcjY4O3yPatK2OZ
5qgajHqosg+2xm8yFSq19qu66w4BjyBAy330QjgU0+UrpoTU9Ioqp5pg96pYDifR
MGz2Tw5uhfd4zYJsvFatxFOWgazLW7+m4qLAhsIQbmGhjmcjZBjPgqDRwCBVTxJc
kEnIdVUP4UIaX1Byp47719maI4GR1FuA/uptR2YOQM9xAww4oM86K8A2b0XmqpHO
VIy6wicfR6tG9q0dFD017Oo4gxf3IuzQN2vc9H2B16BU/frK2rT4/GW3B0ZGQGKA
ZM6l9DR2ACDMpnm5/VOfmblDDYEC52VBUS4jESfgSHWvag/Zjk8UwHY2/gLt++xG
ekV5Wqt9kOK+qXxvHobVdEzC3HIfXG33lIXsOA6/fg05rnX0XExMX4qvX4xIudYY
yOHsLHxBnWyTMgXZ77zsaspKZOXcOsoY+yY0diCsP6TnvGXn1mNxMKp6RhlPwgXL
IZMw4xAGdGrbNkHrl25+cppi20e9oV7o1sxrunxM7OfTl6uHi8TdUZIQuprwtMbO
xhLiHWuGYBvtn8EVBEJz68JIGm4Dgczsf1aNkhMgrMEhRCfws7P5He1DFS/g/D8e
0NJ6jQIgXF6HtSTyjJtUSSwnrlaIdK7Qs0+R8tG3iMnIkpuSUT7I/O5YT4u0R5LJ
r6uMfS7heUS/AkNAVebQToBLllZV0JqZ5cilQyWynwj/AyzfLCGKezXt1Nx1h+u5
o2BZru5GEI4SlGUJWGpCaEhsIxNRXQTrQVksS5y59lA2tS6QpzulYY4hrdv+NMsq
bnCKAplFB6J/5+mIK9SnI+sDGnqN+b/EmcctD+FDkVebk2oOh/lJEZgz9p1ZUJzM
Q2xcaCKcNYIX0nBxxgc9rFbqfJPaBc8gwz6ivMGLBBkF29Ik8lJUc+ogDZG+XkGC
frI9aMGEBAvQK7rr6nztNoLgdlRYX7RNzPtssXTsE6AtlobTEvznzuPP7/0h6qXu
PMPGAT2j2+j95AvXdzY34sDpZc6+s5HBbklrn+G5Tzdm4jPBB72I3qe2bFvjkQLu
A+k19vVsM23l0kQh2tIFwHYO3CzwVHDQA7ymh5eIknAxHWJaa3tOiQhY+oxh3v/c
2cZRf2i2HOslAdP37iFeg+IcDyXzfkoQrJMm4IEPJ+huHUVeElLi20diifloARbC
y16AVka9ahvJEgMfTPO59mc+74GcxDx1tfd2COLIE1k4CrTpUCCp9mEEFx40cHJp
Yx2U+v+kWPSv13QjGD2QXzLn1Nc77xWWcZS0LgXsqEDpZq5nSFNqMpsXX+xK2puV
Mg4S9whbY5WH+b1zUJnxtAq6NcZe2pt81lKOMyDT8wVcvOw3wga0z27f5ULxRD9l
w4XRQOn038M8Zv59AmY7MIANCrfIrHPrFoZzgEX9f/8awg8lJll3AXSEcKcaVPql
XceXfSt9qYA2g7KaXtTN6mle65eN4t+nFk3uwYBj3a/jVfWH3S4qPmzKrxInU1Ik
62eOdsJiIUMLyMK2nsdZLAteS77AMzS0JBcwY5MLM3W27UCxio9pM8sviaa2b/Dh
/JRaOuEJ0CgCowr4PK6BsnzJLAgT3vXtp4w9ZPSO+qR1MgQfgciYZm1OMHGUgFG1
pWCh6Y7J6MD31S1ZMp4Nf9KNJRLa9vrTtxppsTykqgQcqFK7AU2HuovH2FMsLLpY
nU3C6CxOvcbepHDj7f+Ezgf2q2/e4LefMH+Zd5fk+n7yYYjRdyH6oMe0w1okcQoj
1wFUSW3BvL57bDSnhmOMaUOAjiUWnY9KvhVEuGIVUSJtgN5W8W7y8ou89kUyQK1+
xEc92gH/HTXuz+hbcnD+J5+FgvFLddZ1s16hnmghXXWo7jXkspKWoZg4Zoswowt0
Pn9dj7wK9oz8UXiC8dbT9wsjs0wZGlRbBz7yRzzr5xs3HVYkKq6wO1N/8j9T7yRb
Ve6jR9GdDT+uehIAXiojLYKWH/pxLplV+5sKPmtBaqrbbPEJdU05wKsVydRwBLbo
5wmkn9AoCnk5EDzzUvpidKu+NTP6yeOoBFbTlKdWqeX4iUpku3TNEbvWVWx25Gpv
I7XuPpqrTGHC47Y9Y2Ol620XI13SSJN8lbxlFtwxKtPPjEwhEfLP8qqhOHnLmEqd
dZWTgfFiJIG/8lFRuTqQOKwTEpDzl0IOIwk1yEMAqiu45U5bW3Vv6iuWvhqraun0
Pdaa1XLEBBA4SVT3pxzrXMxCfdRSQjN1u4pZkFzscojSSQSeDP1mSiyooz7XtzDS
gBZI0heo6kFbluj4eF2kd1vBXxIjuMTRCO3JxeiFZuIxUMhnMn7b4nTgMYtovYQP
q3JEys8UNWLlbxyo/v0k7mWYEPjg0MSxhnlAckYCSRUYyCVVCFpMkZGSV+77CTeR
CtfMsihLbqUjYor7lJ8gWw4BsKproI1a1Xptyc6Jp8ZUp8QdDVqecfY7aU08s61g
vhzCcwcFMIFW+LXtCTxozxgQAg64wbWza+jWcMyEFYyT9qyI7zyTkfDSgAO6IWrv
SEy6xQ1MV4hcRChwxhzmRjibjXDr6fdScVprRZW5fBZyyXUW7SNos6EwKE22qjMD
ljcBBLbodnK17sSGgP/THfJ7KinUUWRziPPmc3ox9sBuWr00FD4LNSa/QosjYawD
6L19i4Xl5h5X+mXLvuR0AwNYwRD44vNIJ73W4boA4JpWn6DKeZ5kCtatB0TrUQGE
jl1dwAapywL0WF6JWiOc/8l0dTi1tM9jYcwSgpxVqJDj27g4KLevBdevXBTveYG0
pFi763zQbnnRmR+wc/DmRjOk02v0npiSBLpM4z5LdSECIywzdsLyIWiy6HIeXZIG
bLF8egi6ZvgVBVW/T/K3D3UAM9oxQGbBdK8vXYNJNKDFVhexfdjmh9CFJPmfuEO3
i6NrVdcmhSxdz5wRGHo2og5sEniCgl/DSXLCNWXnldTdk9apdAiVYM78X69mJ49i
ABNpeiZ41aFw6vcLHE0oGMLzh8Hr/NmtFg0p7fTowRE9B5uvok4Q+UgcI8uagufR
GzJ1Z0QbMrBBblAsO9gqF/serEW6C++xXuZRGzJaHdE2K/AByGKfo7I8X2Clkk5I
Ph4cOPGeaeiCurC8ujIPeIgKa3cOk1yJlIoaZ/clvSNAeGLiMvnHrkEXZaoEl/2w
oLlVSblb7vrCw1FxTkp2g4F9omCZX2ky9A32c53O0ZmYJ3tsZEZAnmTuywPyhGdM
LFwmiMyYODeALnAslOYaeZQnKYk4igKjAb4keKoO2buiguN4AFJFhOIiTCL6eIdM
9CWlbUFI0bzSpbrKXxa0jxY2gCi2gWxxlCHN2h16F+XaLzvwQrdzhKgB1QQK5SN4
JAqk62m1A4WtY+jtFVIzudFnbO5v8GCHpgA1/FGMccAsiX+9Imch6gWHtDQMyqSQ
/hy0Bo/KmVuitMzC78pibT+WZL/RnnO/55+0X9hvcUQbaTOCu/S9jlS1mB5a1PPN
lK/KGXGcO66qOzDOLznOFMVkD4aZvf94IKrDHtUAJLtuUJHo3PDPXqIImRs5pNis
5VCSgXj9gbJtlQxSi/VuvZOH9IZ8UtUEtPFXoAFNanjI3pUzih587vnWW/mqdlDD
eHDXmGjGVcLXxf9UZEe8a0WQ0uxiD3htLys/80ZKeno4hP4taSNhepBO4HzgwZ8v
EECTabG+F8PKg8BWLicBogohO+0c1+bOSleSj/1TogfVQEn6N6a18RmW5M504A2f
suNU3mLavuCwZ5rgYuwK5Hl4qpwHZ9oTNlZyIfFL29hLvIYzIai7GyxPM4T1q4k0
iIj0ZUlUataaoe/wUst2WKl/L9VYx/bRwHrrb185CLHIijVC2dHzTiXoftttNm/K
sIvgi9qxWOj15SnUjHOHQ7YuM8KZn7a9ZTb98BkUQ6H7s3i84dJWy6VpJxS5l38j
YslD1P0iW7VnORRe0dTWYxPtpMtsxhp4dIxXruNsJgmZ6FQNgVhZ0XL0WioYAFXt
JrcMvRHfMOA7uP0tPTojHLxmxgRoQkHy/49aik5wd80dtcfmsjUNptF8CNXdgIqx
k5mhWd+2lqZh233Ep08wtvlcCCUqbpZySTwZM/4JdW4FoSYPAwPG6oXhNpUs4TFa
QddEF7s1/TWO/L8XByleDnpcVWymrfgrIKSt9rwr8haY2RCGvytP+3HwNCLuGsP+
PPBP82XKUwQbSyVSysf7DmmA77WQwi7N0eWcxMS75+LbrT1xuJpmZom+cF4O6sJU
8ZNJ7fjyPDbq/PwTO1EknFhU744/3Wq1zqeyDX07TfYnzL+QYxzA+WensRIfFE6f
DQZuXUluVs6kMYWJtcypjoMf4tMpoQBTWoyU86uPpEuyXVBzVINX7iavMCXt3Lgc
TvqnqEStM2W6V3wC2pWkQUf29qel4/51LbPaXx5RnZPp1R2v7pGOLy0chA2hG9Dm
U3DKMzzsy04zOlwOrFKiLFo93ZD582LxyEH4RaDn2B9ko3LLvFA7UurkuJoucmj4
At43fpNYEsH5ZWAViPKcXbUVFfpi84B9WTsSiX4313AC1PnLwg4jAKW05wU12qoz
kpiFgG3SZq65Q3VcobGepFHTE7UjOAm8aqsmiMVuY46ME40JUBVbAftCCD1v2u4E
n1hs+WeA8b6qM2BQDanfjv/giF40kTmQPqimrOQ/rFByzIJZtkuQ1E7dXsttChXF
3KI+M6fgZSNODVFFwAclex9PA/aX4P8WXZXjWhh7wxxyM6yh7bo5fOE6jxdln+bL
9TTAqYdBOWBqB6WL29l1aBAYDik7rgYJIRhmAvYLTS/UfdaopQyq5UzoLeLh7bI9
FQ1xEHtWNOj0maWr/jjJnT591pwHUFs1kYl95iRwQ9btdcIF6JHs6izOCbrqp43M
lMKZBPh9UF58PejkeqgfL3BDJ0ynd2i9VJtyAg+mS05H2tfhnRBrfQIaP9zvdGpo
Dw3RRfg1+2D1Gdcg7QtTcC8/jGHAW/S2MN7xRXIi/5pdd1onVSnzsQ5+x5WRFFRC
VRR0vL7WdqHNg8NbT7GHT2r9sBfQzjmlhjLTHUcrydMoJrx0bJayNW62XVtSpSm9
Ib5xw7I+DwrE+vufbo9GIzU1Okneenx6DCr2bV8/hlLYMYB0uJw1aEnxxY/BnKoe
6pUCG2UjsG+/3dXT5GBNzgMfuYq2gPfRCYQQV+z7i7KQOYTRUAcIFE/O74X0mjKv
agLDWcXYzFCHg4lT1QgtcTvxC/f7Zs40RaPhijjzbCCoFtUGyZZRNdkDNgNVeQyA
nPBpaKPooQU9XXBf8Hn9z23Up71PlXnGPrj6JtGxpv+P+mqsFO4P6Yoy68TQ4oeP
bD701oC+1kgGH8TKOhtiYw0iuPvM1HxeVFDVJFnybpGsapdQILVSWGNLNg+wN1Z/
XWAizcacAmYWuxtjVMsZZ7fu6EWWQbFiGqxaPabH26RmkAGarDUkj0OFSd61YzFs
Bxxz1lfceRzcXwFxtAMWv+GfnwFQo/eMW+rnHivDW2ONDHEKcv9VGl/lT9aiMvys
UQSXCdfjjYM5k0ZjZOT/SkIfhafshtc5d7ODUXwuxkSlDhWyNuk9FsZUa84TaVT1
Ygcyo2oY0BU8OjPXObBEFVZt0yQFl9qjq2eO4EC668sO/woX/JZdr5XumCEsOGD+
WQ0i8p/5hNVVkxLXTWEsVv63seyEPTlxEuTHztYtLy2wAj0E1p4A1lU2akKLDlSl
KnXHCbxZlXoKfBsqbOl8RI7mIKNLrWrumZLTZER1/1z9rP1lX1sb37F7lPGrpxnf
utHOXjFPNk0lDLbBlyNqimiL5rxg3c4+Fdh10e8raZqW1fcYA7aLAAmPkmsRqgdU
nXiwEoAk1fR7YzQIIsjlds1TsMHiYNaw1w0aeMIyDYOwYky19/c/62NFadhMh3C7
bP/i1kZHHqWY8AMk188gAiaAG5F0jCfKD2Tah/8oPJgvjTnGrkoofsdMCDvOLfOL
/EGK12b3WjkHYljrcamnkAjxwME+JkPMTp0DDFaJGFufA1mhzeUGvwB1rT+pbpqo
iAJssEDPet5w8v9j549VseRLXy5TKaGPE+5fLT9Bmn7CmxtOM5ZOLxDLiust1AMF
Y5KUBk7UK1TiPzkPDd442PN2uguULGUnLivXKDslYcv2uKStgMR8FyEmp/Tmr1+J
MUdgrTlXjruc9vhlPi4FnVus/wJT8O+eyw7rr/EWqYmA/0/m2mG61SrrpVPkOJxM
zNaBsyLtPF2z1lcpXScms58/Vx3OsOkebHwQ4m92KxI8y+DXrDFg1JvmsBk/7ROx
L4O0HQsuJq6sb5wUKrPMeHWG88afKxfl8+yWM9ozt6DSxp4+5KXwh9TudmakLkwM
J9M3tJy6yE0DxZfQSXe6RC1Zjek3Qnt5xNtfKi8nQCGVh0TiA1KsgDLrq75HOgr2
xvgUTVJZG0ExRPdAIh90r/OpVn6KCy25oq5AO2SR3izQSWUKr5iVibxPeBTpXE5o
Sl+35aDy+L3HS3/sLKIgRzIOQn/1nDs55IpjmdixoC8l0btmOXQSLf2QayNV6yGx
yEiNNHA/nuhGOTrJTviClZHcrLwmOQxNKUwQrLiFpYXtcG4Mh+crVQNPnwBJkaKg
UYMsH7JZ6KubtwLOX/r03lPyVAbGtjBZ5z4CH6F2DTP/KXsb2qvX9cBeQLMma38P
MCfwAFHhR69HeNB9Fg+O8bPdPk29IATtzwIDytxGX4ivZ70XeT2wCIMIdOvajsGD
p3uR2/pzDJNKqBjE4NQw6g60naLFaw0qvhB6o6z/M1VP51tmpb3atzcyawC3Ykn1
ZHCB+vnFeCZqKiUn2/FQy9K+cxMKDyUhwo2K67R0SP3zZwco2o0q0zrauEHLgzX5
YohGyYj62WnJTXdy5iwn2MtMMfs13+cz2IXnt1/QXeVUgAov2XHA/D8x0lnic8Ci
0xn0HF9CHw1+Ng13Eu6HRT6L/XZqYSjgmEyPyPfaCQIC0YJSJuZa61HKtamKdb5E
qJMwmoDVjjvYPciJVeZDJEdwFCDo+AwqB+i5SMzRZw4BbNvoMdtpakKi17C1rCV2
xcNKkNt2KN5BwzohZybx1PesI+Jf9VVvEqFbpIi1eYCNPJk8Fap6kRMadP0kc5sr
0bjRSZ9S3/KjHdGAGVst4+ykifOGQA8BiQisk5yvI/pa65eyu61OF5RfhthAvjCH
Y7wgrFTgXp3BC0X7I56rTil3Yrw8/lmfYAMXRhPqvtDEaIBvmACQNK844EXy3kjt
XgBQIXgxYHptiHg14ihWDKeItAU2Qhv9kTt9Z74k160XiMzPv7xzeumFEmSBzFk/
C11Tj4Utme6yku5CZjnJuNaqgEktEyMQSxH7Dbj2uFmelVx5uiaZX1phmJGKUrQY
Zno671byf9MaHuhFyjo5j5IrD0RJDphGEjNQX5/z0KNQVL0arpYxYBXPdfwppTVy
s7mMxhGq5mwGX8rf626QTx++17LRubr5y257H+jOlcxDfOtyYKtgjdWVnh+bvRfm
L0Eunb9tXV6mtloEMjTWKrOOAay7SksHkVbkCDsF74l/5ape/lEnBBh8oLGuavJJ
Xzap+06VWD5a9WjQsiieffTINhPT1R5by1tWXpCJMvZvJWMmN8VrdRgffE2Bq55Z
dXkn3lrz4LagtZzqYRrwMyIv6hNZhmcOUirBC5G0dD7V6Ny4xfK9gOT6QG+dpeCM
RE8+HzPrMTCRbaWruAu8z5ovkl6aXmTuZMEI9zEw5M5evltEe+dBN69GS36HKnDe
C7Th3h5NB07ADw6PiXVVHkYi/W48EuBEOKruE8UvAKFZcChSh98VIManM9IO/LJl
605h+GotSgKnfFK2AbDC3kEtdumVYjvZ1caCWD4XuGwjMi7NGNStnPTkM9yFtkf5
gkqoMBl9Yva9yceAgRf/i+ABtMy2xegICE3O8R9Y8M7RYdDh8ydqLJJ/ViQ03CDP
JMz3SC0Lo7cva52VHEV4/tfb18f6I+inBSPlCQYA3xPRJqDokE14f1pOk//CxmRM
StIvBBHckVGilu7QTR46sQArf1ns7N045m8eQm+xt3TA75af7iL4OjiHhJbHEfDD
KDear0w8mJhgtdQfV7+BDCqYOj61AtL1sjtgyRtz99ZOjl1n86Ol6Fleb706KHxr
7L1CEtUG54ogK5I0nYaXpc+yH+cKGNAZF1sNAzvnN6wiTkqAiIQ3aHIYsiHlUgj7
ZpYbMYnRqMI4qjmePoKd/N2H9j5UcE8Nwuw0KTsTprB2eBDKN4Pcy/esV0LCv5PE
XncV2Hua3vjY/44h+dNbdAor1ozX7Pv8cVg/MKpq95GNo2DNTh+lKUiUYxQ1SAox
JPRZzzZSP9IL76DAK/8HjzFtJyHAFwVTNDDEYY1SLxeYckTlR1hNKDR5ItRmeVe5
iH08Tk8Ioe0prKdTRHth7B3RJJNgX/rKSalShqqWYGk/HJnFMIsd/UY1uMK3ivi0
++6Ce7rvX2C9EZS7cxMX0y9mvJ06stbb72dQ4mArGXN9361fyYRJZRNVlDNEt9s+
vDnTwBZY6d7lArVLAqy/DTCruTrUR+sS10uZw1jIQ61rl2onMoAQEt1Sfse8Qsck
H7EiFT3JgBEtw3Fu69zRVbyAPu4MLnBvEp5KSN/QgsnV/wWzhfp1iOV0bHsjIUVm
twxOImVVL7iDmnN9P5QQMaoML16hHL734TGqKJSi5ueXHm4tWsxeE3QDpiPJjNaw
ItTSqk03RCc9TTLgkgTxesEGIsJYjaSPagHIdNxFpoe4aqsgTn1smpQ1xkd/EBoA
LR3jTgv/zvUHpg8Do5SF+9wlG05WuS93ZGNPdI7Uyk9nA+mwgy5sa86tbtXje9ue
7e62F3h98XhX4UBMsgl7lJE/Afva/kfsgHKzQvxjPjTA9vt28IH1kjH+X/ZgDIZN
ZE6V+25XHOgBvmf8WeLO5QCe2RR2q0EyO2u4X+q+QYSpJVkXYWSNV+NSj/qEaU+Z
g9RqBRSBa5NCuMSmmj857SW7dU41qjMwmezNN3ZsiPyxyEwFPo2I6MEXCt4paKDQ
UKtHCb+rAJ20tofHrSQNM6/B1ca/j+rkdUBLyVFpdM43cRXXqbnDb05Xd3qsvD0T
3D25wvmpLqmWn7tGmrVQQrpO8nfNPAG6RzQCgBwMmKfRd9jbpTQjrjWB6wa9l41/
XYdh2t6bfyEW7XFlTW67fRnvBU/b4Wv9bhOmuyA8/y0lb8hLwBAw1YH2ahBG9o39
SuSYj1R2pzIDoxp7zdb2VGtxjDBlj5paLkimEnwuGiVLMRkE1FZ2w7+xpZVg28bq
pWztdbTAlJdMm+mb6kvGcUOvEr2QnD8UjXt8LH731ChLayryp7MFBl4MZGq5Khb7
v3h77PP63ViRXUEagDiExceb9vY2zzahalwDzjNBkSd0WDrMIijjMkexDg9tsN2+
rbMgGac7DfVZTF0AL8aq9g8gZOf/YvCWycBAZk6ZvUweMg23W4GU5UlAGrWe+d0U
Xq8WmYwl33h/oMM8eD9HW2txDJz2VopkNcT7S7rHYr6STi3qL0QbhSSDJ8D1tCdY
kCdOizj+DuJc8QAahgEt3Rf2duqC/vsDyXKxuhdHGAqi9YR6S65/94FEKiMEW3Fv
CbT2/98RDfYRkhQEYl5GQo5Hrs1HKdCuPX9rQSrv3OeHwX3zCx4OTw9/fXZOjsE7
TVbZ8Z7K9TqTPx5vz+5AtQ+2d3xC05Uo36/GBFk+2d+5y+0kI19dCTQLBvv6KF16
zvEkyS7IK+2fbpGDIuTi3ttYbY+GzaUB1G5FIxFAR2axvaUWfgCpgU7ip033LPqe
OeKoxAq2iET3ykw7yFM/aRVP2CpUJMFC23k4kVUMipohR09hguHLyt6ziuOly2Hm
PBtg11Dz6GYRyc1/rwtJNdyhdOT1C4PwbSj73IsvcCeq0U4x96nmbbcOtUJ5pNbV
paP9Q+SFiwpkbSYo/bq2RBPAhHoD7ej4T/CLJgoB2mE7mqBmSn3jPMnonuei03PL
ECzuL4jU7sHS1zIbzDEzYXpakup6La7FzGa9bOfjRnpCl2aoDRiyt6SfDq3nZ/2V
C8lkZd4RdEb+8oBvIm2okDUEbqk1r1LhRCvpSBk/PHB77RB/tM2W6mSek03/ZjXg
cmK5BMifQj12enSra/znvMtn2VVghbXpkkrA8Z5FVyV2KwyPFMG5QHzAh//XJf/A
JAZWw41RaYyXCOqUswmEyTPJOnWrVh/Q0t/SggaxbI6beNsOJD+9YdJAj58zlMAY
7lGsiJkmDG9PoZewv8G7eHChW8g9gydbO1Ax8bNVZtemBk1Mwes2Iry1xRBjPBbA
/FR6ai6tjuJRXLQW+zVONCsnWCAWwSYIusDFyjdEwQ3JZhymcqsllu5mlBc/X+x5
a9sCFa5KBVmB6Xq+6zt6s37ysNo7n3u3lO6oQq6Ugt5uP8DvPjp0EBtQLZraHStj
tMfXRVHDaPUCOSrrhFdBaN6dko0s6/FLp7Z9DIFIKFfKX23LNa5XWqpA7Kcd+TSc
v0CC3h1d9RV7CpeH2U23sw5n+IEGHmKpXrScFrqNSI1jY7A/kPVY8Vzu2p7nTZN0
ryj/JKMEnpV1rwAq0GQ24F/ZzobqgtCGTss4SNBooWWD9DkizUGma17Rdqn2ev2O
uCkc2P+Z9TCmeXHVninRzm1BotMLew54dmA7H7FUp+XPwNljNotymjspysuUnKPh
wYuNhAy5uZkOM1CeEmyrs11+pPAykfUE4qabpaSxoD1JGWN7mMU00/XGGm2wHVMN
Qvs5D7xZe3IHKaEr5r14acQmeCI/eBT6/JQtoF6yq1X1334t5bp2DfHYkH3jfT//
1pb+ZKeR0b8t7de7XMN0Q6pW1Gaa0HeUJV+8PsogZTDj5woiqwhqKSDg5bsLqEyy
lvM0y5WvGde21SpszaiVCAugY+DApSWDxvTw6vrTxfpgKd8M4i+/LiNFVkESA2e4
sorvtYdQeZ7cFgsMBYljcG1XLoLzDQmDqiML5kGLeSt6ptEV0GyTPYqbnKkKkoYr
DvMQZ605JLh5n0rVIQ935L6/+Li9TR8kr4BS6tCB8g2dchgO2xSYcG/ou8oA357Y
r9peR4SwuIdR1GgLvjSllU9+H62vQxbY3qupErZyXHWs5PA9xflv36Kbh1x3xUNM
iZRW8bGVvlBt+5rM0yqiymWc1k6UAlDxw+R5zRrQSPPkAwBq59A/+LC5pm020Q6Q
54dX/RyOmCmUKr/Iyi6pWRqS18CH3q2oududKdB/jIFylUFC8fhB5QdNhaDDuytK
ouhOgTTh1wBsCD4MMoMgUWOJz7SpO0Lz2Dcp4/pzWu1p04B6o9UzJdciBfz1Abwk
7OlqTtQHWShLvZFFrYgTbp31CipoqVfJmCdAjhz3hI6rMFkAxNIRsVFs8M3CkwGH
jOBDtHtoS6qYonJPbXKeORXwVT/NKaCXfSHB2nDQGTXJ44QUlvpL/IU7sJ54zjdt
oofxHFHXbAmkai0yOWaWTdNgFZq1256NvPJ6ZnxlQzuoeez5Ao5dSvRf7vXbfnGz
Lxx4FpZTS6/BcP3fhW0b2gY1NeT994BvO/hodtKLeDQeUB7aYz+qf0QyqdAUbSSV
iK09P3oePN5xSLGkT0PqdrZkFhY652usehZZoxWeLCIZv2c179rCOgwRslQeYVP9
Uk2VxTDngYrk+Ck3NjoReKdLBYQIzRdLLusbNaR6Fv+cTcK8lMN5WKv1lKSYvIiZ
LbmJUgYX5+KccZLWHg8a7VbDPZEjqNaOrIC3mHOUI/NLK9rkyVH/g8GjC49lFrCs
Cyj2yLfeF4E9t8bg7Rd6ssu424H4Ai629BYIt6aRa1WIO14r8fV1ASvadhyTe7wo
KwtYBTnRhZRJqSPiumFsUH6f2FL2e8s4vzioAUlN3HQi3udlE9cdvcYBv3rp9foJ
qRPdh7HnYB8N1a/t2JndXybm1529BtGdfnf3AVC7qNhx+6k9bZg3MNgAsd4dtMzr
WWJZEgGSFZVIa+dZaTMgnfoLGADX7BarcwcxNZONsDRPYMjUxle50umfQJZly7YD
vcJcBhAtY7U91dS5lYUCcm5cn14KHGqGSKze4LJM4yPxcTkidlAmr/Vke3cBIYAb
5tU2qobYYOBhM+orN/fHz2oByDxqmO2gS+xpC9WXNcxJ+mCLtB8f1eNiY8HxU4U2
UQS5AMzx3VqIB0NwH5mJWNYc89XfqO5icD4lXSDHZMm7yLOkAWmkhZq5S9inyJDP
OEwU+T1wRgMHkBouuSRSL07yXuEI7/rteGRP+z9cNt/lwAOfMeNoMG9aUPImIQjc
YQ0sBO6Q4G84Fn0FVPWdXI3RIkXVMW8892MUZMAXSP3ZyWAfvSPrDjOySdDcB4ch
tDYxMFrvaYj1l11zTVICgSwyBkfxwJS8guRUB1FBqpa1e6l5DCnSFsLOipoIe6yI
8pKtn6wMiuku+wxHJqI0ODQn8lmeqSwRsY8IVplX1Q5Ulex4E1NJFPEdFEbjVDvw
kWmWCyDoRCiWxkBQwBqiCK+jFRySAdgGN3wEvvM09SfF7kWQBqgjDHKXr9MmGR7o
HlBZMEO+nT5Hydrzg+PQw1zZqv0p31/rGUjOmkDQuK0UwfmMrQleccQ7v5yvKjQL
YGcaqg14WPn0lZ4hRAX8XdDtKUgKbwux+PPC5hgIaJeWG8CD50hoV4Gx6hw02BPk
FfNgQbfJ4DDEKX7ZGaVAqbndbLLqgUU8ebMht4HXyJBm8IOXFAR84WeaIH5ved1k
q76/Zjruz/zJCKe3nPAWTqlN9bOap3rkQVhV4drqChK8liIyCdtRK5WfbdiKlrhA
A+vIbdIYlDXBYCVeEuMWIr5sCF0y0SnJEuSCeKYOVxX9nAKawqSaBeJ8qXkDHxIL
J7obysQUG8GmDs+j8T9RKi1Oql6ZjcQnb8pp0lY0MZoBm4hbAbcexRRsaAfS8byB
4NSnrhi+ot0k3mFfef4Bm4H9+8oLupmWPj4KEYqenDHL2YzpRkbp+wmQq2bpUmQu
KM97d5n4p1FIdsfNMxh6BsqNfrmu6F+0MmBdje39SNfuwJgHf2DyDkeeTkSli2hf
kc7T1rbJd/tun1BPq7EDSVTZ6Y9sswR6wv4VqAmnYtmPb1zxiMhKOUs/frV6+bsv
U1+GLOomZs+4GvjoVrgKTjafAfen5oTus3FDpkU8Wa1xS6+IGGIeLg51nC1afjfQ
88LzbTC/yL9N7VADOugBkv8TpdLf7Cowc32JQumaZ5axt37mwHfUdGxdJQ97f8XF
urfGWOKL2Lt3/0IL/2LcgLZhfibUI5pTlSVBuOH008viD6dOIw+iIg8xGRkqdeMW
vT8MlfVxI/p0oFwgURO69SnAOLBwxB8vDGdBakNGwMTvwjXgwuCVa+5slnxcFjtW
D298P8lt1358inLUJU07zXocDTQE3w9BrR2tBkXqp90hwx9MtySXActNX68YhPjm
qUtn3jN5wwTfA6KnrcjIAE6alYmlUGg+hMuSz6zLYjq4kCSu+CH8fPLxcyryItXj
C78Yk6AlLnk/c2if227yCFrZ80k1bkzVNtD3UON4g70kmMSnATuftn6Uhh20fmIE
gPW0SGJFytes8+BHgp5vpnwBjudnGGva5oD4N3/wkIlKqpU8X2IQuMH25dlJx5dm
VWtQArFnUN9Zc3od3JccIC6R9/c2fgbu/uDIqA52fueGjNmhCFiMymS+5gGQ6Yv2
/aU4OXX0KrYrzoANrCZE1b/JQpKlPdpUKE1fMyRrpj9/MwCJJkD6Rmprbl2QbVkr
+oqWXZxj9UY5MZwlf7Fk+sjQWSXlzffY1Ouvec0IHxAf9r3z7dFo/pyea5g//EM1
11poIY8CzUpnOdu0VBS902qYvkq6aC4P5JPORha4ykt3kTzlIbhSoNWZBmsONRS6
0deDQ2fOaWZcctQ4zxupzzQN0UcuC6N6U/eEcnLdShhLk1v7W5XfkQw+FlnHEMaZ
0enJVq78yrR8H+v9FzE53BQjf3eKWqhxB/K6zPB/C/ewdtaUxVeagPLYmH9I7SNy
cz0+aaDprbPhvHsW/3MJuNd/+it7fLmOOiQQ7bp9nJCAU2tlOEWcnikCg85ZG+mt
zhBNpETYoEHqIgsBYYOMja3c+Bfcx6X2kqN7sVoCp6BKOaga7EVS14x6sa/0Ik9Q
URlcIRQOcGs+bDddB9Doem/g4yOB8D6Uxo45YjZkI9vmirYPH+v0r7OfYy3ekx2P
YBQYuEPNKR/L4mIORyKejjZEdsj3bFO/RE1FjNTBKvoeYYVUeNMXlHDJML1/wo1R
l4eO4cOBpgg6mbkSryoXIc+czlF2MGTAYcDNMJ19lVDftmkZZn9/gQGdLSxglQg1
owk1YvGm/Nn2PQ0ArCz6fuSU4GzMwg+K5a8+Yy8mseWKGdEr1nJeBXfEgOiDC8rD
CoDVbdiOf7ZFXzcF2JOvBAGzsZCgifAu5rCm5qsTeRnc6cBnaE4CTGqq+s+cfZfg
02pqi68eZJobj96mJf+uHm3e/WQoPEV3FCYEmEDpnYwpH6wTmELfTbE5G6IXrtjL
BmluvPxjOzkmcgny672hmWo//2zB6qfQCXQ17sQHYTzOONko+cHod6WLlkSzGEGd
fsLi5pbPLDVOV+yuydv6FWWDTlLJ2hWVpwHyZhyZu/nSASFD0CwglAIto4vU2DMw
GIgt7HaNw9mZt48H50DB+MIRLZSkDyRrgkA0Yxe6zD2BzAD9vUkUq8w1YCOgD5Ob
FpLhfcSOTnkFilv2wGtLQrxfeLaGT6+TzaC/0gPnPDqu/bAdHfyeD7xCGtn2k7rx
5tpWOAt+n8BvcjY9Hx20j11zSw1Oo/b3wY/rvCIN9emdlWm8iIcdRCL7brXvMZtO
vsfWDnxwscmCy57Bxd8IMS5el8OjlQY1Whgsr63Ph2t9E4PZx/cMF9hx4tU+qYIy
p2w9myI4tPS2GeNb8JP0I8T/bx3o4KmUTOt7nFa19HmW6Uo7VSsR7hWfagcDpDpL
0t7oDKTU+LgY5a+hsF9eEEPNAoZJupz1sTrm2xGCo9vB3iSrOmvDHWFTZwCeAzyj
KsvwLGwQuTgdr9IY8ASR76vQ+uz0QTK79V/NA1kJjIHnNp5UG7FPZtMOPy8+oBvg
SM5urYY/q/k6iiZCW5a4HDFyWwK7pQtcJdKzDgvjpAM3oQrZDXoSR2OijVnQHHG7
Z/YOJvw0P/VDh/peEhzGTNDvgoCzcyA+4Vzi/WKs9jENGSVyQeWqoxKDblQ+kO8B
JGwpJt7BZ6KLGUkRYMxZjlXGRVk0Zw82yHmffAgq+CWVdXVD2M40/kjn/Cv/uoDj
TqftpiLqaGzR2pC1hjs/9udv5bGq9LbCByozHO07m7Ageh6tm2NABgbItL6vkrI5
C4YZd80I02sDsI0oVqkFi+9MWiWHrXjDDw9YmCSWQ1KmGMGFHW2qYFH3RLSpw29S
ayef24IC0661Octz4IS75drr4jFqyLR3/56fSHbecH1wmk3C9icOdeby7rD+jrwN
9E+r1g8ujMgfInKkPGPvG6l1RB599YdkCiTOABQW3IjFbuDcKydqd9r6BVxOwSbS
v1Wfu0yemXvwfw9bwVZTK4n3/HFug9d6mEcSMo4laG+JDZpljuXk5Vn9N5kd6OnO
NQklOt3z3FvOTComISV9FhqBaXTBpxDMrlZDwFmqtGKIVWCuv9EiHA7vK1wPqn+g
KXaSlatR8USDosT6pGbopBPpC5Tqx8nDFN7Zp7ZpR7LaouocJ0FLDpPy0Y4Fp/VH
cSFNx/B9VsTstCqYKln9jkoAuS6aDtTOO9FSOFA3rV3Iuhr3dj69djmjHKixM9Ka
8boBIGlVLrFfieV5/G2Cv/uGQAyQUKVq63eny+55Bw3GaCx86zevSu8YDVXALtEY
4aSa5Rew68gmJLS40PigtPseH4pmgusN6xMsCGotzmzzjzVxPhufjfkmTAKs5FzR
URmpCfdHlzSunu15phLdklCfrWGVNBhmdjhXBmz5Ny/o0YJZU70sSHrzNShwAcdy
XMGcbWne6oSmxX1wzOY/KoP58oagfqdDhnKflIB5i4k9w2/mhG+FS3de2fv729Ay
TroDgtKkIiUrLKhi5DMPVWuLSHDewNz5Ood1F+AVM+HWpfVNdZ6e7Y0Te853il2V
CWdQVfOotBSpAE0VcezHzPRHFbo6o5rXzvOQotg8xdXDfu1ckyEg3dhUry8eEPc2
ETPO517iaJapako/W88rpPMmGwJKYHv/3AZAZ2REFoXZm1kvzycuQX5j6TuF9ncW
FOK4DSBt8GF9EXVlhZGcG2uFo5TQdD3DV/6ggu7nU4ZtKXycj6SrKYVj9oiDobsG
liKQzhAc/uzC6htbZokU5DpP1ePR/8jqZ3XGUja2rV78aQH1rt1kx7wj3WeM79jr
q188/cUI/fpFCWOjTJk2eUI/GdhRqcv8eGySaOTuhRGOa0q7WNnqJZo4kt5lbc8o
CaXuhugEn0TXKHU/gBZF4VUk9n514pbAWUHQHDzs5m1B6yYoLFOgWE5RTZOBruKr
82xv4EQtsODcJUtP+gTdvkX5DHzkyqUpecUPXg/9GllquvLk744jG0KjaABieNq1
YLbdxbj+NHJZ+F49OBLmeRF2qvnlH8UQVR/WDCmheQ+jYfsa7u6EQqKrrx559UDM
26ucGdk1rrUuwda2c2OqBT7euFi4+5Stgk9t8YWQUfObC5c7mrHTnYFSN1DV3N39
cDhN1tlBHg7fA/tX9/vEKaZecRJAbBeiG9zKjJDRLq6aRmLoyHZ1eg/plZ+FkMJz
arHwKGnbSqLIaRH8Bs6c5l1AX/PMobJc6if4/agL6FQxlWOpc9/QQBU4gDbh2KCq
tBOTAo0zaBUnX7eWqvyQc/vdrrT8ofyRgAGTWp3NHkHZkIqny3Bkjg6R3B5kj6hF
7MRIrA9zRBPG2zuMG9igkeRLyF3eb9fwrr9hC72fxmpwzeT7EE7F4UzTO7DnQ65I
QIDATyGcWbTOjcDBq8nM6d6VUW1tEn0uQ4LedeUsdodR7zI3rAkjxWOyqF7H5sih
CqkoovWUau68RMpUwMf9i96kw7/e6f4GVt0fOJ8OKztzhJw78pPc1lfjRQH4Jjfx
Y8kWyIGLnjMtttOIwEaOdExUNCx/yB9b8pBn5jI1ZccOx7qkr3wYGpepoJNV/7G8
W+gGNB3LJl0lVGoQfxbbdm+KsYVB6Onk0AwpmhtL1KViTPbmDy6l7sqPdb1Oz/gf
S2l9j8GaYXdzsOGdHuxa4lUstWfvXtI4/Q0IVoZ94zmf2FeOmzH/ye1S1tyt7h6i
q+s8k8icNPgVBQGA+YpMXTFksG9QclusIIy3QuRqlKpFPY1PVb+2X6IAFZ1N8V1f
qUGk4NQ5Up+nKKgI6FdN1cf374p4tx8TvXMaBomz1uBryMvg7x7LFJh3zXNeUEaD
fN9ffRd814r9LY2gJeCXknRrJT6PTxht0LY2+YgzCI6W1woIVoKPP1dEc5OVIgtH
hpxA/FUD6waWZRcpqu3kGCd9s6/qSnD5lVDgu4zk0Sh38XotleAuWlE/+isnWOCe
zlR8Tk1XMRuhk+GvLL981gD7LmtDV3hlyR9Ts6NBRTyT8QJ5ZIv0tqtydQsplYr5
sVhm3yKvp0j2gLZ/qfnzB6+scGKcrjENQaPnPMjovW69JOgVlT1hdnu0Z2OH4B1h
AQQrf/D/0oF5SzS7KxoOX6kwsyJpHES9lZn8Uq/ZiokBL4+CyLqWCXnwtNCLi/g5
+kUjm3IdQ/r1qDc35a+D0wvP2H+iZ04jvF5qbu1lPlFAxh+In65lYn3JTSdz7oXO
M23UQjgFshQ1d5RTQOkLYKkfGY8C64/azWXbO+TFqMnWYZxOGQHCz9J1OeaerJE4
gWJyHPr7KBubf3g8JJzvl2VnN3iEqYeA5qY7ki91euDJcUe8xbY9L2bVuLTwO6Pe
jlKh4Fg4eWRwHBFsyfMVJZ66ZtChINBSCDfUtvK+QGSJfbMXFhdANdKTGPZa1/UG
jPW7AWYCc7aGKU+CS1Ofvd9GQRbroL65vkmDxleSDEkONOXnGldwqjOXSk8xkPqv
bTeZXtx9j5PsqJVIGql6xUU+daSMUg+zd/TVq5NHu5FhHijAo2lFAL+c4xtrqESW
8MLErh7gu2UEXTlwCwiXH1c0vSoMGFWZ9jGLpEkI9obTkZ2/1XAieFdk8Pt64SPD
kC4/bCb2fFGBRWKI6ktz3MoZyI6h+Fx0vNY78o2p/cvTv+53TkxH/ZZ3RWOamtsy
dZhmqGUuZmaSPvX38e0xT9FqzvvP1QB985pKhr7aie8RC+5jLINp0ElmNCes7H6v
IMH8lDEQiVbFPJUuU9CgKS3Bd/POfclvbju0HnT1eT8pNGucMGYNzI4RQ0OfEaIe
AITxqHAbpPrXlClfAW5E+sth0NuF0fnBKbKNtZh0zGJUpAuz0gGlIKCb/jHA2WUM
Eot7gngILRlIhAsAq7pu0Uw5GKOi5bjPgrO40AjQU6gJnXc0DLtg4EbVHXn0bznd
rxLx2wSWQVMuHcu57TgKYE6bhkiYBf2Y8vDbi6Eea0JeNjb5lF5mknRQQTA4dvkF
npk5u2mOdSdhhgYOcvHrF3tYg+rBxd3LxU5tSyfv+/D/0TEL8avjonlC4h5+mp6F
YKBh/tJnEnnNo0koa1bb78mZzMTrSk7u/NZmfsJIApeJoOPWzmCR3rECgAO6aaF9
8Hc7vjnkQhzecjYUG58ynaeOIYsUBzt1+X/7uQzzwDHwbPymV8Ra9LL0EYgMdHjq
ay1B9w0LZT5qS/3ah84GkQx4BCDk+jLLiO6dwAX5hvsh7TGj4lLJaxM1ls4f8kpe
NyOCUm8I2AOiEjZbqJndFB8s0WpLFHvOO9FEvazKFfWAnMK5T/QXnF/2mFekOkoE
34fbA0FpBMYJb8+o4CAH15S/QHKEwxnTmLc3MD53CiZEbMZmo28pRXGWuxwMmH0J
Njg+iuhdV8c33e0uW4l2RCUe7byBmLfW44Cd090Ojc+eUNPaLu4QgPnR8Txi1xLB
bbksgEXiAdRGET1mYCLoqM8KoNyQbfQ8vz1cgNPVG+jwFJq69IEUksvK7bId+Y/u
K4JWtAMiCzjIK5q9NYi/L/2Qey1Be4TpFo7lZs4g9ICDr8O6MHozKeUdhwaFU7CZ
unBuOiEDpZUrO6tNmsNqEcxRZHUgfHVfgrlntuomYrnFvu+UUDqKCJ1fn0jNPDve
Im2TPGdGjEZ6P33sGsUv5Jw2at05TVXD5L10HhRFMyWFjpRcfndS78TKNO7nTo1L
GfLwoymp0/JNFpiADXI7qYmKKZd2wvTyeGkMx6UxYWlpjtXCRTI4pZMp4HpJoRO1
grnR31XNV4pix8M8NfRjWK1P4gA0rRH8TH8Bjs+5qjumHWFvBKuzwayCn4US3Cq5
yJcbLm9MkTCpzrtUhfABT/DZEdk8kZRIv5HqR8MclN7eEOJuXK475ZjYuntc1l2j
pol9OwKXOoVXv+cMRgaYCtG+PZKrL4rJVdaCNaqLrpc2RbS0UXujfK3RE6kksPNR
XERwt316Eq8RWsEHN9USZnvhfNQzu7MEX94rZLQIAfS09zZK6XMqoFN7JXr3tN5G
iFBFcShGWSPuRmCMzLlyWF531VIdzT/R4JVNjWVSw1Ce97TPgWCfEqvUmzqbXyQ4
WWADzvoDEt8jvtRlAPFCUAoCY214E+M5Q0uixfUpBJ+/R1ibdNXJmhAOn+HTKBzV
B4fWW/Jm/t/U8+0e2IzbG8H8c30WEpLDWBuivJMAEfnaffTpav0vYnP1ZcAvYya4
uYIgsH5frBrTD1Mg1vPuNuD4pUuUO6tOPIBoDaTtxnoyK4JqytiQFPSf13alxKgq
NreGJeDXcH3hN/W4BUJCU0zb24LNyrBrDao8nGkUUcKIfbHlSPXuB63LS6Qgi2NC
V85bTpjQ7eNPNvLYcCOf90LWdnl/Emp+n+lsI4Md96kBXWdmOqhXJDpYEhwiSa6O
lAea5or+4xHSfpoQ1/zdTow+mQElTygKYLB/GCoORjSeSDxmUWEDgqqUgU2cOMDF
9qvxqEZQVEVzLWvAnLTwj2/y2bHDjuEVyGBz7f21niqJPbk+eQrceaSo2vcNGPVN
O8ZUzr1c/25u5RCoH7ZqCZmdoPgPLMOD0pvXWrl2yj8E53EnBcZrVmYRqglLlL+M
Q4kec/fSf7TPIQc62DFMj5zyZ3Ts8o4bVv0k9Bjhi9obT6EOss+lOrlgf1ZYeZKW
Tf6uLbI5YcHaFz0FkvpDQ0DpX8vSV/6N3jFCikuCYm/xC2kuo3yHGmy6QX3mMOiy
CzGltq5JHRuDwgbeSxEOR6XGjuW049Wu8AcF7gJYpW5y9W3NbpYv0ru4OJudMksc
7u+aX7NUm5uTOKlkbhKXG1st9sSugi4GmIb/RoyNYC/aMA5QCz5Mu4xlz3/MSWAW
sgfeWV33Ou3rNCZKB3CS70aPh+1GLhTd+uyoL8ua59lUwKOyeMGpxhWW5RH2BXeJ
u9RKRC9dlWR0erakz7Mz4sj8qZct22Q0oHrg0ehpvdftyLpDgpXpRPx/i8GUSkjG
AZCDC6KeH+y+FY9qVdfkgEEN7LuRBlAUwLVOiWNwjdtxRE3LtF3/yDD9qyEdY70/
E+tI4ce//Dc0bIxfXKiGxFb0gi/r37lvaR9MKO81gBnflGjLneizrNwqa9s2szvA
KgtgXmO0De1l45pBYowjZBEXCTl17dV1PB6D+8d7wmu85gQexnMuvtnjllz7LJNH
xuCsm1Q7UbIw9xD2URuSZMsfuCu8MCm2rSXjWNu+MmwpnpfYiddwgoQN05iR3uqz
FBVYstM8s0eKZ2niLYD69yU9Hh8Ut92z0Wt6IU4CVLOkiGIVT2Jrhigtx7Vt3dtZ
S7wyRGeyEKkKoUvGzhf2auI3Zj0GQwdE3IG5ArDFCnE2UnhCgO8AyrUBg6BAxXll
qgo1WY/cWLbayLDLh64uSu3Av+ZjxtLHieVlOPCd7G7oOOQ6n0XdbQFEBQGYLXrB
9Uea5ItnaBd0dcO9+EutFCHg1SPvEQfIP9Z5bXX/Q7FJCm792+JL5QSTYLB1WYND
2Pajlsz5T+LWg6khe//MImGDkyib0eQva/puRHmtg8jP4DKeT/uFFCQ5aB5xnC4s
7Vk7Gjw1NyyOmaiupeeEPy/wUF62KeLghb0meeMUdCIW3sYikrQJ4/gF0J4gt0a4
KG9SItMmRuuZ4Kk3EevlurQwqJRo8bLACGfrrU8jnr4/xmqrCBDlNQeSsNs8OMO/
vSpfa2qAR9EoyddwrTRbC5Np4qAFPQXNmcTxlq04RlQIsdQdiZVfXf5uhHmO5GWt
cMP++1DEUmxsLAGUTqsJtZN+wmO7IKXvsC+HpntUj4LiE+MYhHLEyw5aPMQWYQKt
w32++gQNZDmwW4vTcASubArFLiJoqTJqIfrTa+4cmWvhbHCH3TmJG9rkT7YWHnOc
e8aroRfoXP5chDYQ2e/kym6Gdyo+qosUqtbiH1we8iH4YYiOKNT9YcY7a+bvb8x5
UDhCPRW/4wB8B2NqFoPLGEPGq9ZqLjmpZrvFS0Vixzd6id37RzeI30iq2VFuIf+4
rYP/m/AFCN57I0LDM1hBJ5KAvShFm5hdUCoVQCAy5FdLxSAnTWt1obRQLVopas1e
vEXDwL7AJqN/upSh+1Yvh/AqMUYhM95mpyetodoHDNNoTS01K7bsnbJT8+G03Y3c
t6EY91TMVITa9dOz/HSLpuae/kqbBH6hWR8UpPoQu1Pd1U++rPFdH1RUiqft7R97
aDdNGjsRniykfIooGnLi6IdVyFlB+545vRPyQP7/y8yAXDgmsFJ+n9EswI4JLnhO
a9HI/r5Az3NCv1c8/TrFxlHmOC3Gco9EUUVKsMJiC5mI7r8MFS7D5B3DnkDWUdE2
Y1EZTqRvzvcnKloAweaxHkqnjk7fNYz0xuONROsxJxs/+n/TtL3daQ7ptcUTHYOQ
Xzwkb3e6QnqQ0/ICuYIk5nF6Rh0Pz7su2mbNTXlMq+6e77982x+3BOfLEj760Srn
rSDWyykrMQBjQfox/8GpcBfBEAKVIwoKvqeyOV5Jd16llfSlZeKvB9dpAR4M/Lt0
pbL7bkrgjyg6r15OQL4y0AdGUCjnK8uPkty4qVPZ/2BHA2dj041+4nakpRyb6L1j
Ue6vMSzlfg0Ve4G/xNTzPclurh9qJNAKuW3uw9G8GgaY0ClOSzN/yfhw3CSOUkdT
BRfioWy9BBH5UVS93Bz1TJl3UfVli/USZf909tu3y1PdKZoU0TP2H0jABKylgQWq
r7rEyaA41Ogb5g8RqvYMhczlhay8NWebRLqceh9rliuQ3Snc1CGLj2vcMRO+ds2e
NyWtTHuvdDl6f0jO1FOGWxqUmcPhQogztGtKweEmHQ5bfW6X0RxMpb3YJwgC3thc
5xvw9m9OdD6UJgGBIJS6SO12RvJv85hjGCUpQliI9DUmAM88y/hBTTl3zRvZLsDZ
4P0mIoXbEniRskmxB7DEn6lomuPu+EX7a9EgTt9PW+CNkiBQaWUFtsSmk8Z4lTzx
buD4oh3C4RF9N7pu9sjkpgREF2K7ApPNWiktvbIXQ/jcBpL7IKmnLKsYXHtC5eGD
V8jgWRSRf3zYJLRBUE6fdzo46k7M7Qkz3ykbD7fX5n+Cd4LmfSCn1vwI9P/t7d/i
iSir2cZL4kK57Zet7Cy+ZDOZrqse0dsTKnZ4hBgzmiUVV+CJgIL6WhYCoYHi0Nq7
/jkgVfI5ZqT5WuVWOHvN4MdytDe/v5bFSS0+3ja+mfxvMA2ecBChtlUjP706AJPl
RRbDEBHwyF9DZMybMGySOqYGOjfaLDZsbYRdpklhX+fju8P1u4b//8WWHQWQdQ4m
HQcDfsxNK/QMJqAehPVaEaPDGxHW/WkhUv+GQVNGiRObBqWWn/+6eOzyBVkNNlax
1XCKIN4arFL9AySvYmu09iyqezbrXwc8bZHuTdW2cUz3WOEAaC83A+CGHiD/Yevq
uxmxJCIJP+HZ2BiqK+CQUP9HtgwcK0lcmMvlHqDwQUK89mmZLvGskfsmKjjNYiPX
X54QKBq7ufivaSXAe/1JBu6lCIOSVuRfz5Txuw3ZVhQFSaI3Hha7F8LBCUVYUVnQ
ZswXH2mXUaxCwplyuAu54n/NwcS9dHLlFA27CYFPP6fhHry5d+y8BdjAm7/69LOM
rMIvm+Ee4UUzYMbkhw2Aqe6NhLD4CX+ZVFEmlXjBGRCjvp7w/n4yP39+EPfb9mEl
d/9LunsrO5eHIqXDz7koCXgw2VS7IbRQRTJRCxZO8ykp+eP1+FfRlzga7iK0pFm5
+ZNTLZI/jjRrITx4Xz91SsWPSmML2S6nX/YIg5qlpqggwjFj8k6pP3tzWNuUuWVT
szr1Vlx10lNPDgKhoPtjuFs3noVduffooYkd5JdJWNy3A+E2NS/oh4tpKaQ0ImHz
TPZkMmwt1UJU27tfl05rAkL3z/bzGQFIG2a0QNteERCkg6LNNccN3LstwNo9QYpJ
WY2ImQVZjpmZy6UHzQjTTHrD2Eh5tErPoDOFTRGK5EIHsqe4brKr8Na7P8wg6YBk
2m+0KhbCn9BIQi5QLPetMxRMCNc1IsuOYp4eOBCSXDlAcGcvcFfXnBN2ix/BH5aG
4U4SvUGnU0OrDHRn6/48MTdz1aDqVTOK+LU22x1u/pdFG4kaMOWlaSzIqzXa5lYY
3qYvAW8EsDB3oX2e1J0ZwNgP77+6FmHOWOH0GQcMk9tCmarNwf6/W320O9KhYuuu
WDU4Iqs+UfGeyPjR8QLbmpgXqCJzkunUfdmEKfcqdYwFCvglGvCLrLwx6/hBO0PI
uJyXBNpQaaDGcwkz+dOjkdDjnfyh9hCjWzTcIV5aqPyuSFkxgwuySz26sWgDNQIN
RfybBusnMqH3o7guPjyhuKmwayH88PNEhdK25HGYgWpIfH1pCA82RbxoWDhizZJa
EOHXcrbgg5oqXN2AY4OBCSTxsTg5gXZwGG+UOGsSfyG68e2rMBh5IRI5mbIyIv6K
p2KXJ6SyOZskAo/FOeaTBedTgFeFjwAgv/ROfA88oxPoQmkjc8oX78eul9AoY4Qk
yGBP3JdB/fWOPnbKtOMhgF94hV1lIuGjR/r9GKsymirWhbILmvQJ4EL4CXB/hFJ8
dFxhg5hIY7fkR2HpUkP1UXmHUiysDTxttvfcJsTURSaKxWud8I2RMPEYJ+IFZ4ZH
PyAteSmtYxgNetyZmfSrZlMDUK4C+TjhmDGivrXgdvWCNoExXhOgEsbXkK9G6KuD
5Gdy8Zx2hkv2ktwJbX3KVXepvdz6vHY0trhljfcPKHbz/tj/ss/bp9TAXquchwix
HvuJbnubSmwxbBDNU71HfdIPMzyyAD09wljFlNuIfHkMu1nLugM0FjoKCRox+UTM
uLt7WmLC27zFBN8IbLN7m+7TGnlKdPfytFgZqM8a591+Oigxk1zt5n8U04WCMlv/
REMuPcoctxEoaFkl/sBeAiztePDoGsbaXSKrqPOjYcl67q1evtxWwBVxjpBnjToJ
7R/ciOI47JOjdFPq37woIE4SA83g4A1IROMPp0GMaNtkMCpycq7ScodX7efT9yia
RiiFxcb5gwtT0qD1vnGHxXYZLq5CwlZddss3LeCss2rnoFO7pxNzWWJcvbXnEccx
Xti3HEV4ejShLQhmwemw+TCBVO7Tm/dvqRZvkmjgwIiScifGrJ3qZ3PnDzQG1nx8
d0Ecjdbvrmc2V7VxuxEgDyzRQ6KZtI3hHPFdAZLdkugefg8IHdN5LKQ+6y9X0qS+
9+MiaZjza0mrn8hSYeLvPF4KBvj45ga/l8uhMD6vQTR5g+0B01q136+k/PV23Q5v
cLGsjsdJb5yYHzREMPDTYaRU+fGKA0wPb+2ggI8BV9SBsNvFwZL5tDVNLx8AMXeQ
JY+2A68umpCAXgieZVX70vn6RsBuGe/vd5LcxpZts42Muj/vmTJzqAOI0NN11EFH
YCcoXtxf2fzOgn+43EmzcNiwCrRoYcqRfPRol6pyHmqAdXXaXF1dXpAUH6e56RqT
8ia2vD+4gTWSdwIU5u7A6XXDMxqW6pu0YxMErl2qASCxr+XbL0P5RBSR2q2/9TJL
ztcmychumklh1IS0Mi1XTpiKb3huTfum8cP5bFVAk8iJGRbZS9fCnicAsXt2XasB
9lrQsDIoxZrZMxdR8Bwo0Wx9zOMTgfD7MjRsto8Ky+wJatUk8cEJQl3xBNzygC2y
Hb73508R39PlwIXsUHXDE8jljPrb4iZCNbOmuSIK0YDufYb0ffkibKCzDZeL3O3Z
BcIYTgZx5NXaA2caUcV3D09gLYuhbPUhbV8oSfgkDMds3tYm8z1QUjFNXfgO40lL
7Bb3BK/wecJuKJYqvEouyClabFoHkZLTlQ/hvSVh0VzZNO1agyZSuZeVwXnVRI94
lWi7cMTgKsz4Syynkdcu2hkxr/vQWX/lYZzEkhM+OLFAhSKyG9g4x2fgA+WPEuFa
/xE3akoEH+AtaGyqonvB16u6tMhPktkZAx1s4XPneaiSVJGXdnsjxH6VMvft7Wzn
lp8Y6+/gUWr1v5vmvPQ7PsMJ78Papdc6fLXv7pXQGUpkJ1e5TnPk+vlwnRAqeopi
IqsBpTNg4NQMbr/CP/DW9cs6pCTZORujFyilSsHNxrPInk5pY18a6POw5iLUVb38
LY3v3dn8pj3qZ1wpiyBZq5pSe+Tpx4nii9hIP0WHj0Sg8FFfXvkzP9uSM0RvBg6D
7YDueLWuVQJr4o0W03FFFqL4GYR9Cl6lPGiwfNtLSLY/lDL2Bs8n66loSSDOT2Bo
fuAXtdOPTilh1mHOAZp71XJLhMVtycQ/757EzcZZ82rwOvcWtaTBA7dxQvS5AJ2+
wIYfhSRv+JKIX9h9S99xFDVmaIqGovvaRAVZ5tzHlE8bLz61a99s9rHT7sSxvpjh
dHvZozhjsRNQplpXyOfwV9wWWpTiv++tfR+5fS8vBcFNrUOUggPu6Zw+XMVPbPRb
r0s9oUG+WHw+LwzwsxNcZmveuT1yyQKBcjTZeqNGyrBZ1NCnJCzPvMs9NzENsZ8U
7wRqFmp1L1+wYVWr30OmkTOQE6WprvD/tGYUo/KGG143CgJqfMn3Ezf6rG4pKnGa
njyJbHZ6jR4RHOYlv/G/qXhMYHxiPPxETle39dgLG8YicwuVqzsffqkou7AaUJS/
nE/jGcD7OW1f1qKf9VBu+fRh51msR8Ufh1vf0gGestGanbhKQ1lMG0X2OXkCkWbB
yppzqNShgIsZ7U9k6EPiNzC8Ry35PUvMd9uEu1XF+GNE5i1YYvEQPhEUj0k7Ba0G
H6bOq9SJ2mvBQEjlblFrMR1sQeC+yK4rWHJ3CYBSJW03i9VfrmBK3IOOivJHtovO
SRjGlQHW9CUQS8rplAQn7myLjzIfxcdZlAet3TWf+6w8Fluazx1y1Yj+wmUJLp7T
Hw2k+Wm6yAmOnzFgMKfgrm/ZMxHlI1VY3amCh14C1aQoaSmb7kz4gR5ADZ0P9eOE
PHrGr/ZMbRmW7A1/oWyXSYuI39DHS6e82lUWAZE2gXjnctk3pqogPL4IgTcFEYmg
EhCvsZjnQNsSD/WKckDg+XayqFyZLGgNGi6pcOrGNAQfVT1y8DRVwVkXG7mZVO0j
GD8XgdxKl+3u66VEDYMUODnCaNZCk2E38U9ep51rXgeIzjN1unFyfg+m+IGf0pvG
zDbekwdxlXoch8cmrmvCQwf7A771Ofle8TvFzrgqyMx+w7LF5kLxcHpZ2D0R0oSh
NXu6CArr6Avk4wDYqWcb2KqD7KwWwJZ2npGZQgZHvfC+rFtI1s4VIxuhmsFml3q6
gzFpPqcYqA3KQti+kH5t9bHDb5iauH+iRP3hObVv1oeqWbq2rvSttBUk0BaAbx4o
oAPbe3KOOjObK3UVTlGeX0Rhg94dyUrEpjtIHXHGVG8IVoE+3mHWnisWkIiN9Aec
yX+FXoTiPVXvQfrZ2E5kHWsbKKT1eCAN8hq++E4LpKJwUW3g4NE/hVmIeQwefgoO
gc/XcJvezT4D+MtFXIQbXMSHjFL+eYbWy1tK2E5d4naWJnNdSRndWax2yo+Uwyu2
99dLcVw+fdIQc8WHvapQoDKsxv88rmHMiDY+p2Sfy0B3dHmAs8BZsZWCRbyD6zeq
jaM9lWmxBhYYepsJ57vIjpWP88x5wagpMuTOv5XFAX4aBpGoFptJcDOrnBsYJgeG
I5vyZqqI8A43YSqDN2ALMTu7lcnAPQ2oU1pxIgSOmtTL8deca40sZcxiQSAIvX0V
1p8+rPr4qC9EHF7QVjDG8hFqxCkTNk5Cs3Upfqf4lOc/HHTqj1rzYKHNFUvktX9M
N5hW9ZGpSNqnkRRrhkXP7TDxRf2kM47FeYHVWZGZrcRjrtrrPvo+touD2osd5al5
xDpY3iAdwuUF/wnXojWg0z5M3bpjrlFRx384Dr7Qqt6bM5CEbx+mQOBP/nq/y1Mc
kqLCT5M/cPy4s0zGB6JSxcZpDK+bkbMLD7GopYvPy0rli3EIVp6d7K/HWgaVFFTe
YTnT416ebcJNSMzqM1GpQPE+ZURkAUrd02CylC3a1OFkM98u3rstE8cKSz1squFW
0i15tqq0Nzz0NMHOW0SpnVtTHZjSM2tSwYZoOeTSYRPPh1KfrClBAHyvJMmSQkTB
ntnQGpiLvDpgQHJlVfNLapHxd1DQLrfgnh+tQ6OeAqIqcnlDKlASGUVEQ2YjoJaa
PsF6zTz3sqdnbRTthUEhiRBagDDAUGkcdhEqy0NSUmlM2xynX9n0qiV2AU/xoDwY
c+laDLno1FoqHTpEFZaoobvBK958J/UFfX/Sa72IP2n6XAFjvI4Q+/DBfr68xFrs
zzT9p/AtxUDIm6dWCE+9Bk9axluYcaJrLHMhS0h7v3rlf1Hq6kxit0lez+dc6Z9B
sTGfiCoiDC2yTJYWt5LgznwzFgtI89zILAcEU3XQKc8DKmvS7DZYTuz29Zq4CvHu
/2IAumnnwtJoDhGYF6HeczJREJlDlXpgLom28po6q/+Uufb2gHcu7OIz12+Pg5SS
kGddAwOIqE22zAojSLWCvb+ssMxTjV0sMQc5uc35epgjWWQlAesPHpnFWNw4+y9Y
up1AL44F7dLECOK4S8gVCpANWoO5fvm1+8rjieK+/9+QHv/IQy81b5bHmhvC+oF1
JKRYwYYoiL235ZOllY/BycROaefTHj4iarUnr1Hrx32uRhEWc9zBHWG8dvzTueEN
NnnvDZn65OWQorg2lg7HbMft2i29fBzouXwRJ8QGNK5IbghrNcyRL0wc2IGw1XXp
K2wYBABxeFFeepxEltMENDSBa58ebiqo47MVvu7p3FvdaZS/tIvIK++16e+wu8KM
rW37C8DiWOwxVwXOUY/fExmoqblV4oaoUO3zwa0qzA2j4I+/PiW3xBozGY6UKlqA
+nZTZtBKM1eTLO498tVdgB5mpd8oezyECTsK9yDmXOSkZK8So9XMWN3L15ozxaxH
AsBuWISbr5D6mKQqg2tgLDytxV4QYX7gqjiRlseQVmaPsTnwWzdveQbMDxttMHki
rUKsJbq/sDp3gwe5TyZba/Gr0QbqjUaINCIxEojT7dDh7VOCdM+4kqhBvXLrWmcD
1g+T0YtosoOhPUimORnY8vH9w1CG6m+MqlbwDhL0lj46pjNgoASa0kIwUvnf21ZA
eX97zGCl79GL/OXWX3YGZnPJK/JK4sMmSpKh4JgSTxqTOelNyuCvn072Wv+rhOqI
SwfHBqhmHHpCiG9SzUbJOe7oL3iA1lRMtSXI+FrduZWEpkfmPxTMj8JUEkLpLUZ2
3M9BHyeahy4Map7mNMrnlJbtaz6eTQDbvvtU9XC3frGsnj894DFwYZojme6uzSZB
Cxo66RYO1Wg6DSV13JPJAiIJTis0gcsSaNxWpoIJ086wBNt6qoW2U4AfxMF25PJz
N41FZq9ygAgLEZpmQcMX0gaZbPjh8i/jaqImK0TATrs1fOsXySK7VgjTznjuYo8/
qVGz2DY2t2FpJZenh3oti4xnR8CWIF+0GlTV+LVQ3VdYqtUo3eDEKl5ZBwn4SEln
ygRXVJrg0W5ue/vLlXOibs1A7oNNl/HHHIuHZjyquCp4FoCRdQDQACBhHFQbrHkC
/puq7eF43cT5DAjjpkXtDZQtJI10u15I2zWAp4CprM2Xpi2nX8t+F4lrq08ZuSkF
jvQcD9wVrUR4lEKgRzKiexyPAuYu0zSqE+n9cfTlKBS+99aGWnCG4LkBpLBf+170
lKyHVHCTZZ8DWvxTYfbu0vrTk/XtFSTva+PC/IyqKw9gMtku6xn1+2OoAOOA0Kvc
lVwZ0okRP+UqJkkVeaWRsuwkY16Nwa+H4Gv/h/gXrvFky5RC53PiDD0N3vxUWz56
fdBTNSodrDJxRbipClLrwqRWiGbfzMFyeuyfzYFkbjONAJ87SUJpJv5fuvkGy4BM
4ep/PTbcmEak3HLBfMGVJgtzvrIC4dGUZHVW2nbbu9zyb+Hu9aUXYaTWizAjKn1O
RsK7jnURW8IP1ABL1Oc1mMUCLFuZgzMAZ9A0uFSKlem5DfTE03mxNW2GleuXXtXt
mquzvvqb4yWaGR3ZY3SuZysSIaSHHHf0SchLQlhwUQfcqpxRrwgGteiqv4oYh3KM
iRCTpL/xK8iZ1cGQtuoCMM9d3UAXNTd39gbjQhTYRmAHwoI5zlg72Zu3R4sutayR
idF/qs9xr3W43+TZAK2IncZYGUVJsuCFQ+jCdjqVfxDlwka7ll1eWoK6ga+/rriS
dQpNdYi9VvH/O7fsQ3EN9IenKMgvyu+DyksyF6Fmsg7jnz1tbY4pqspqFSEbUVRk
VNsYqYbvRZvFv5TtwbUXd1pyCHWgvcjrrKmt1xdiuUDkCSGxpkxY9oC8LGSyHTWQ
LEl7Xx+GKCRd0rRcYtdcWhODl6n3qH2jzO4M/zmZpLNM/aZcTkl/vce1GXZOsJ+j
8KCQmptH3bPKInv8HZYM7QXt3S+3jrPoGaQUba9P7tSQO+ThkXg0RbmKr7QDgl85
4b9ctSTmwkCCe+1A2VY9UbaGwqAzY+3HJTjkeVcRd8tNCFZt4h7KV+senPvN36kq
EXyCTNW+MZUuJOlkPlUdRHpoF7vUeTal2JYsv90yt0hyt12gV8N5C7YI8nEJI9QX
n06+u25f86+iEbiOTb8AgpTUWh+3YHlzwC4Mo0sSr6nW4WBeKFiRIf1kKwW0w2+R
31+w5iUE7YlEVH2QqpQ0LLRCtCK5KO+Nlh5oBWx/37uZddFDZ2O70Eoh7IRJLZJ+
0uAOyHuTXueKqF9CD6dYSOCbYcNhrfzq0Aalmbe+K5lbxEk8tkHVcTDHexlS5K/Q
TWG1I8HcbkzAPEIoWS9S907rOkvqhfqYu1tUHiTN14uOH1CYi6gkES+tUIJEe5Wh
cfi/Uj8GzQtG7XgP/95Ew4AoHaSM8WoLYxPSFl4gGMArzslwDjYTPEDIz3VR0but
PNImnwuFtyskmbl4Aq3S608FbePMO3eJWXQ9oabhXCyR+4wL6Ig1T94l3WC9zm7y
0BHf91wJy8w7TValHx9CZmH9fIgDqhCtgSZ1GlZPsgpgcP1Ksi7/P5jWVsn4nL0/
ABPuCK90GoAlQH5/Z2YO3cQG+MDiGPk6YSGreozh3D8lSvyVFCWjhWnD1NiRdHBU
SvWWHYdS1IBnWApBe1uOaspuM38uKdlKalDFTEcFypu3+KKPt9+gzYP4N/UVNaap
ahbAGMqppQAHkcalhDX3SENeZsY2l+AhKZafERzciVAEZhXKSCA/tqQBjALdQ/pN
Cub2KM3A9lH1vcg35NFIuBRIvIV7O30rQRKpXFJhRxsB8bJaRGyLNBMESvpWFHmF
gVDBQ8nFJvm+xiOunUsDMXS8GQ8kGAylbTxMCn6plXcEsMEPeH0JklmnsK5r+czp
ghoGfFt4CsORTqBXVWuWth5PCQ+ZPXXkQRcSO1zRLGodsOd/yY3BAWwm7TKCB8yw
C4a9A4uQIsBJliCvyO8NzDA6DC4E1OgM7cB48UKgpJiJ+MD/M9VR3P5pqBA/L3Zd
8Y49ZjOq13qv8XxXb0zJrLLFTmqBUwJHkI1RJUhH5VTfeSqnWk/DHk7JtQ8enCi7
ckm+vf4WMEYlsxCdGnYndX7W0RCieCe+WnLHN1bhbaiUNBUPGFklKBCaAX5ncESd
ydMTdhwfapdlsesLISgBwAaVYTpcNYTWmenZ5en4mWMzTh9FIugF+3ME11k4ohWN
KngmJTkYMB1YC4515ipebeuxIP3BoXFzPs+KVUvs9MHhl1YqdcGiOOhnlaRl2LZJ
yKiLa4TYB8CGB5TffmCloJZ0yujLW+6yJVjSyXqPVdxXkHXM4wAMXKZMTZQhS+Pn
y87HtEpvV7wlk/1MqjglqjPdIhnlE23HfaXhJ8BBjQK+YPP8HQQJBMhiWlFJucH0
F81TM0TKg3TTzzig55DPQZGBYounVfqkTfhznLoKbJ0zYE9LqJyCSmfpz9Bu9gUB
Kp/FivYCifpL2/rvco/HusG8KModn5AKKLMrxFgaKyIIVeJnZq8mqx/PgM+kZUzk
Wx6KnxcMlAjIZlY2MI59RLo6d22OtBRCRqpu7L5MQGMQVnLRX3PVs4KUZchMhXfq
7lwlK96Zrf9QbNBRhFv8DK/5J+oaoTQweWyp0GRnbVny5dYy45NvCdOma7/DGNZR
zpYXrNq3mH8qVORfJa3RE+wDkLcH4xFJt0TOSzoefVh75kJpxDWv5hF0i/zrWxht
ZsM4mBUjpfzDgc20zN4h1T6PKlSWm4sJCcANQjgQXvqXn9HiHtZ5ZTbcu/JaW7b7
ECcY8xJ3986iU6XAYh1++p15FJ7AmV7ATgJXv7nY6RP3bUzS2wGAXJdchEJVc4uA
TlbKiEobhuKEU9n+ZzNPrHA+dIadZuj3p10gDwmWN9Cuv8/fvmlWy4JLRBhUreBK
iZG2NHIpWomYXqsG6eAN67FKPm5xRgT63lU5uoLzTue3lX4Sv7bXkQMJZ34QaggY
rWwhg0hnbYP0r8LSa5W6vpIIPqNxHI6Q5g7900MEc1h6UbGi3Tp9ax6Fr0Ngztyp
rAOCnj6ty2vOyJVGGRdrHtPAYwytHdaaiG3qDBk2SjCMmPpAWKUfRiG8GH4Ps4w/
AmZwATIq5j3Ep6r5lR48B1SQd0EoklcuG7hHgxp3AuFh9G0d+ODt4KvsKO00Qj2M
1PSHG87NUJk4Fp6G2nbL0wU3iSIrW7cDEeuxW+2CgxaoOvWcpc5KGt9yX6r1GpmZ
sKhPFkT/nWddislQEbYU2kH9A9yULsyfdIsluELjWw5APH0ZK2lPJbuiE5zpMriT
Mx3o0kS0DozScoukVrnr/RRiuUynriNw86bLR+o7Kjm/ytCHwKhtKXZjSuFU9kF/
jM/ZaSZwJkUo6FGeV3EIxXj7oOtUmvTihORV1mpzUZRAIK29Jz4haZyRbtotP1xE
3BzI4xaNWKqvDnbYZxm9E1yh3SXhLIsSyEQ+4ZhEvAFv+du0Xpoux1wzOEovWlTS
AHLHL+ur2IpfMTOy9Aa0eLS3SJW1xEej87LfIXCspsF6RjOTzHlT7tAyiPo+SwBs
dvN9Zf7QMQWIsr4rhwL14co1V/L8Ar0RDBnvL0lAJmMXAfamknBmaSKOttlxsA57
YeGxxkz+NBbhIWotoUWAWZeB7koklci5P9omPFvDSEnqHK/4WIbps67/F29zfkE6
6ZDgfpuWQZE8m7wPh2i6TcLiJ3tn1P086TWa3iv8jpNrpwry8gEz1QB2C+7RvThE
ABToE4k5bwouRlnfCqFA99kjcyElvaeMMyLKLYrCpEtltwKkbn5Nv1LeeD7z5RNG
1HcAx8sNchQ/MOFePtHNVl4J/bBTLWaeJmJCpuQhA1d/8BxVt5ro2WwIYI+uC4mo
dQZemKw5QXSZj2USYBkjhaoVdiSdx/YI1XZ9zYMC4SIJ7O1olulTuondIw3T6QF9
4OekiAdeYgcJi69DEvAQP/XaQVNOCRxtitut90yoepYDvqHbEWwuDZ6Cbcdsytxh
FJsMYZClETud9hj2RY3gkIMRyGoVnFrHtRjnJiKdSMDd1PzBH6wQ9KfndlLZhLpx
gaaaBBvYYVfUI03VsiXP3xLfevojfjsTCCSdj0p4B8LSMKkVnSypnSnSYBWZtj1X
CjuJVeRtDhKXYe5Qpm+UANGKzY8vkK1btXA8Mk4+bAMS/oEw21MqloYRy9jKB+Bh
A9r8fiaFaRBrlld39GZtJmBIHwrhNQKQWwgpwXhkmpBzGLjfZTWgktF23dwcVVyt
YZzgB3SJGRIdml4ymvyXTLO8fYVHcrrGLy33D/rJ+M2+55hbdHgAo6cHxCu521l4
7NUpfKKVe0M+NxNG5TQWt/LF1yeGFIi9MvOG6oeB3Wdczru7uTosoWSKYIMqIC8i
OodA2ASsqHswUIi3H7ZwOZTVKrkh7IxGXfqxDQzBo1jCpaB0i4ZUOt0Fuo84Y7Xt
JRAw6pUU7ecitgSdaWL482tKWkXmxQgTd3qUEyxBn2JhNjKqjj9NLJajPr0nTHyE
drxw6MOc95X2qVWtffXzYSMcRYAD0e7swIBQZwZ2hdWgKeTX/hs8Y+ovbJv+KRQ+
B24QF1axBXf90KmGAOecWwSO96KURGEVKcfRpzucdrYsUeCnSRFeaojCAnVoUv/g
zWhkGgUpDOFX2FOlGLeZlDnFd6rhXhydD/h6WHG2CKcdeUBTydBR71FV6+gMEVSA
sjHK42V89UZFfu4S5uf6zYq86+sbNeYkVoyBAzCgOba+SOQLQSvKdBlgb70I8TEw
wi9A5M4rJtrxks+UZ1dWtsvfEjQVrKnttOrHfjHg6N6Kmv6qmOEIPycmhD1PdodK
k/xG2iK11qQHs9kNmEPPBW9LoyFyE7ko/VM33Xf95JPmVnuf+NeKhgzsvCwb2cef
a7p31Y2VRScClFwONUQ3cpwacgxOjUsm8STapIJY/lEbi/pb3LPAAcSso+5Pu1kX
5QuXdUS8UDIVQr29Tjfuew5eCPpjEGMKgMQylI3U8AaeuECv3VTBWzhIchuj6SEy
Lmp/OYSFhls4sboY8XA/s/uowPAmmB4gaBcglVj5jmHmj8dGksXdNSEXPbTPsB6h
B2rrg8e+SnTNJJ9BkCbIfGRbTks3kZ0FrhC4Ci5OMFiFszUAvxPFYmO9IFTh708X
EcDM7F7h0O4AnxBi4NtIMRITasxIVHW5Wow+cfy3a67wIyYktQ8shATYL0mu8UGl
VnzEbc8Dtd4fLO5AstV+Sa20o8AnTvysEwZZnisB97n9pO+fSxAveCbWh6vOjzDK
JEORMCGPzOUWS4XmFalpAgiJSTBrRHURB/lNzadvaoZBWI52VAnRcFVz9+PRoF3g
0A9dmtW/nEBddSinbuwOzJhblmyO3QU6rPMPvffbDR2EtUFHCDMRKnWQr2lUdOKg
0QlZSDWcpyJeiD9picRCLJGnjAlgJ7SkQt07FJQAEr9IwKw2OO2ySS3Jmp0fmKw1
bNQCzvK1WlW1GXsO0Faa9KOTqtS7XbT3aU4CEEtTD0nQoIRYG0poQsgNmuwSz2r9
FyZtHRpBZwhOKjOIF1Di25Qt1EFo3dom+0ycY90e2LGZtMRxqRd76JF08XZFRt4Y
rFPHzegYwthD0rEWAwG4nPMhcYM+XrguuLZEAm+01NdYsbmbtdREPLiwbqDH4g4l
w44miBkAZ1q8x2By1KE4JolDZAQHx3KS+zPhnYDr3X8e/2hpBIB6JEqOtZfqbIY6
TVvnRwIi0B5KzKoqVQbbVcsqUhEuf3rhnhHn/nkq4Cq01KYFq5LbfezqiuEpvlQp
H54kNv61HG8p9jLikxg3Z7O71fpZMcUzOv34Q5zZq25lBBtgu/cqSqW/P98hvHGU
qCQWXMQmJqmeKMwhUw5ZCe6mjvwRRsbbnNa7CbFf2JXoo5g0HItMS/NUoRre7WfT
LvgLiFUBYUE8lhJDdSvNaZUjBRJUuaYKaeO6aAtG6TJL5FzAA107a6TGSSzXTpYA
vXEm7mMiuNLQI2H25vIFH6Lqxrt1HRM9oRuri8KNKZ8sGqnibnnsVTLJSxr0+FZH
CWQ+b47RSJskJ2jpMpuPGdeFMtfcCRUticjWRMgWXclGk0+OnhFmai9c9C9Cc/2P
Er2AzouxdBgbm6n+nL3vKCvIjv8npsx+egq+gGDHCsG2zYkNrgFRooEWBdLt1T0p
thh7LoNCOV1HtpsCN8DHlh1OZDuQaRgVKrgpLlsrP/2fQhXeZRjn9zahoIgjisoA
xbGQ1YtpGctXpVxF/yytMXqcqBbMrkvxKEMEOGh6aUsAL2uYpOh/POmB53LzCllw
6WeACaptQ9fxfkxUlzPr6geSzhSMl3x8cW8KB+9JU6VHR92yBxryZDNIaEX/N7Hh
Usc5jLhBpa696KI7ySpBZRCmGNzq4vZjBvlIVxYyS6ziZFCHUtV35EnbBMbhbbFT
0J1VD7d3HIZoK9TH+N6HzGQaUCtc7HLMokSg/Moa5b5XlIiBS06LePsA81B2zrYg
OQaNpRa52QmYt0HQ5Ip1LfjfRPAmFDF5UkoFqzbwl7AqyBO871DY6aShzTNUK2gt
Nv+MtSSJXCMaSVCtfcAzXYdkArFAS42s0V1GqVqKL0pVOv1EU5i1FuIyJeuChgaB
nPnqssuAFOOh8FwtJLLO3Dqqd65gBdry02oRPnGlGbdnsePTyQhLR6fhzJKjpPa3
ZsnPze6J/w7XyfEkeVdLlHWLEtwZEYwixp5MRB3g8voI73K8ZTG3O6Z7w27Vyymn
ngQlS+iZuKFzVfLDEbQYgTmfiajugrqnRm+tSyqe5soIiPKztBvnyccL0WdWu4VS
vjblaKL9Hlm1Da5G9ZxlEQZ0ZM4nXKa0cc43I8ajlZI4O4gq6Oic/Kci76Ffr5Zu
1ek2mqTPsR3En7wCSB3x6hxsM09j0ghqyT2VhM/0jnv7QBc6/QTy1zRqniAsyCZt
LjGpOKGJOMaJdIeOWf5E1E0F295WdzkqyLzmKFv6sky/wPY9pGUDng375fbsYJSH
4DzS1oAepFR4mTNiNzxK5uYaX+pjWIqZT6NUfIccltsMNCkoh9NaLMcMsvdYxFh7
3baFNcy4JUiJzzVvAWK+HQaHU20Vo79S6SCSBps64csg+nVgdDvnKcKtKNrpsP2b
q38UQ3EGsII4qxdEMDL5q9bi7GK7FrHEu2Cui339leFSBBfG5sndCRijFukSZ9Rn
rPF6xUAGKHQf0Kxhwvm4WlhrG48rD0wsH24jMNVm4rdLM6keOhzf6/1/RESAaqMY
rMSlFohZNRdV8e5KxQuQQJAlTgWN9+47PPzupQdJOpMwkBnQlQZe+sQWWoJEusmF
HelTwv41AZAqArM4YAy8JTp+QH/GzTnnsnvVYvXUYsy7WPFC2vtoyEYGL/hOa5bl
sxDUSu3EbppkB9IDbqAORFQFAMC6nHky7OaOytLGx0wSGdeZQ6yoPypqwBdRm82/
5G3JGiQZ+6tw0t8bTZpca2Nlbm09155elGLx+Sv793KTO3L8MLXHlptr5RA+uJlF
3C06JVEmNHsK/gV3A/v/bbckAe5khkzEdOkyStgf4SvzNuGwO5J+kLb9J102ACAo
aF7G9pZQLWkEpKou52uMF+lodvujmFqdCrWYEu51k5Kae9rKbJhjFxU8Fio1Uwzl
kfguLGHIaiPZ7vcvYDtU3jNAv0XzmYy4gOkZEBygdwn076utcRqpbCnsh4YpJOA2
PPopx2TKcKjjIaQpFu3lJe1AxP4sGxDcF65jMHjDatJlknkFN72/ToJjoaCH6Lpx
FAw4CcamXQfRJy4Om+EkhEtNV/JAFGnNladpdDRyW/FY3w08jegIT50t+kNh2GiQ
o9BZSXr+sKfEH7t+Paq7maEBHTe7h6VBbYsJ62GUNUl5rr1AcmnLyG0qt5lp+lnX
sIebekwL/i6urSxWva3c5fgTBie4AVtXhLPHi+Fchd5tTTrPIsV25KjNFN0CsAxl
NEPGix/+1Xfpk/YyfSorMMXfoeBBMckulLNelC2LfFM4HQviPLaVqzLzDckZzY9m
XsvvrrZBRPKovZG/2Mce5+HfMzrG/SCvM/7SAaZuDKwo45jScuMQlKTuRiT2GSFk
p+GvYui+99e2aDF7IhzjCKGsPzfRsKmwfL7VaP/4VgawsPZXU0wmOq4KfbpdCyld
hjmqaqc1Ci1b6chMs+HjMB+0osfwoyw7i9q4nl4Q/qUZVEbnHKTtJkMPcYZZAcxt
sIBorsMrqyS8xdVUtKZz/m4t+/LWzzpi6HnSHs+VMW1gzb1ocvKhXmFFnkL1W670
NGgdqPn6bpTXdhW1hdI9K7YnLcMPFPUVMZJ8pCafqYaULIW4LToSSFSLcJOjkZDQ
YQfq6Mg0XmkNigGZDb3ma9ET8U/t4M9Vz+4gOa/DeWgyKXUZshwcQWwFU5XxfrBS
sYv+qsyIGaBKbI4Opi5tlJ4dSViJAGnA9vmq4Ns7OJPo9LISuUhx/AVTEFu6TUJh
j+P0ia5tZeK5HK9zhIHSsjdsHiPCptxP9YV30TzBKJfraCVB0YjgnbGPWSGjlfQs
cKfBpTQxmkjr9JIVJ/sJO/Tob0VvT4cF7da8MkGbG8cJEwUcZjjGcqmILVDsbYAj
oG6iCKlkZ6ug82+oj1bAoTbmq1i1HnfOH7GJs1eBRBG44XtocgaD4tiljHyheVaH
yfqHMtLHcIGzn5CatMitbtbD9sesZNfIJlYEa/9C1sCxgBHpk4+xFwqgAjuo93kp
C4WDRWpGOBz1CImWvCcZFPt6uwDD2sW83ZAXHd39CnAKY5Azvu/NuzFkwm1oYe5x
qvw9Ha02PUKPzE8dx2/86cKJavMwImfkDpsUs/xfjP0Beeej4DdeGuU33Fvdebex
i3Rm3CtVvbyeiqiDpucoF0F21yO0NVKoaWsgd436ZkhSMfF/klbdUOnv6PZqPR+U
0jZpl+chcA3oIFcKwfawIqBiBc0Zqty6x78pD9r/TFcmML2jBEKOlpcJQKbLYwSW
hTHHFcS6VoYH1UdN8VrlC2GVI4f/EH9ImPgbnesllHQsgMEEdfGJn9s7eNed6NwJ
B9kSMqhtEgsRYCnxFFJytEpw27YR5SGkzgScj9IhruON9Jg2Mk8AWuy6WtL3hhmw
hLAzc70sVm01hnSxCbfKjNw/mfqJnEoZKD8uxmIc3M69r88WeLejApVp3oL6zudU
tRivmBIiC+Kuw/7yEGL9iqiDnAlhU85azZduIAraSqHL1rrsHqDl0sC8ECr3AO/x
LLh5sXPkO252yD6lBf8Je4tirkAbqPK+PbHYK2eZVTwt8dsX8UAo1X2u8UTZ5CVE
7f49Tx70+87D7S7IhLqLEoUuSBkwKaw7EtXMuE/gNtmZC3mQt2XbxNRedQzXNvbF
gXv7XB1bgeholqXgZpd3CCMJ5jjFpvch4J5mKv8VNeO7rLghDZyky+4jjZlHYOAZ
JvC+VFYeXtAKogZl9Ul/fTYsLrAefsgLHCrCJ/mygLkyAk3V6r+gj/sNtxbDf7wQ
mUJ5YrezB5TyRjdeNap2FRNFW/HEw+rqmyU5T3Zxh/u4fee1QAhAeoGgg7wTI6Vr
W3ldhWbTbluXotfkgZqhH2cU1zqKfDd9PcBUl6w+p+eg9hS28t0v0wcb0fY6nWP0
ZlCHs8k4M+V1UtxCDsFUEYjzGsFMtq0d83JEk0xXT0vhS3w6zZeTU12Ikts4ftw8
oGTIkib81kiZu9nUqQi7OKoiSrxLSxU1gpksafXavwkHjukAkVdDgbY1eBbQjFvQ
33UVJvHOJoAers/9H9Qn/Fx93YLRA/bTQGdNU1ww10jByg6AnJfKM61xsW7WN/kB
MIkNn9s3t0MQKtcEpc1NoqgN9pf9rOiRL7FKW4/2dLBe77dgQKf4u9DwapnXvv3y
YcGAGeOCYy1ys8/imD3RlOFjbHMMtupVzPSnw/ri96iJFFTmnLdwHlBZ+OLeslyP
Bck/NuvYDNdRBnZrKNTq6fgWkJ5rvPVjhxGcyUlbuqpmSsAkJWpoZlCp5qlYxO24
kpZKLpgS3kyel+haBBT3NrhJbf1COAOuxpv7OUm9jp+Ziqix6JosROiHeLXhZOgO
A4+JAOrk7Eh9+Vybng1G1cU4bqMXgS56CApfHewYbF7pMRGc38PwznSWE1YdEsi4
ASoY6e96nheQi8KK57x/oR1rSyS2tDolxTRcpsIZOSPt7VstnF7EAY/2mjt8irO6
F2J6S1A8QYa/34cEIhDxxPMPTlN7a8qz8LjkI78xz+TH2/Zo11wfsCdzCPEpvLOg
gRIV2qQAfXWMzQZVoLfiGvr8hUxSx3EBZtHkHrAQ+Ddw/Xu/ASsNYDxWYDyS+jT5
nK+Qds8jBlrOvBvc8NeZp2DWQ17K7IQwyxTP0tobKHaUCNA07y7kb83QRePb0204
kHJ9fqqjayLj+L0/gEM2FX6Hkjlnm02WZbhCxKeEVbKpV8b1VJjVuIRRw7eUD2Zb
vFzKII4k7wjWZhHPD1bifVKMGaHsGbUXJ29LX5lz+kZXjNvQFMyGGA6WAhv5v7Vu
4GEPbYMqD9dNHQQIGpsojYGOSoeUSgFKNIvLEfMG4mBzqO0NzWOUHE1L4IBJZxOv
GFvdY1rrh/O+czuiK9UZKPawuI9/jjlauffhWum8ItD+qbBk6yPvdSdjxBsgcM4i
A+XjshZUySZVid8lnE2CZGhYR0YhMSBll0CccqnL181TqTw1MPmxwAHklL4Csrhk
m4ypgkYwnNSFPHrXmBb1okdQLmBGTrbIP2Sfn0MjhXiDzYkGMDmfj4daitP4XooA
64e6dUYLhhWEQaUlrfbusV1NDhLhewFPrxtjdT8OjPB+kZlZex5SLtL7hKmCF+bN
pvMQkpA9tDRw3gXW3ajB+gSysZRj/VTtLkrLb2bxDVeVcAjp2VDwa93s/nxJrjS1
jkIefrySJw+7wzveMk4E0QcJ+k/olxq0jb7zSuCS+9nWI44BLpjAu6XzIefy61Ev
XgFr46vmTYvAyaLtvx75SF8huRRNNHMvktpyRwwYO21dtG/LPW2gmCf3aVypwuoQ
bcUzkCTsmHkMa2nd+QTvQNt01f7iH7XVjkUhmtyFrUJGiMIb0adjSvXY02MLie4R
nQmly93qQDfHvzAAHBT01BpOorpAOJ16zYziTr4+Em4cCsJFXN1Tt0BQTmQgRlMl
XzpPZOsJ+B6sV8/vKqnnaMUof8TZRxtbAQwnjRBR6c2eAQUKQy/C+OCpDoURndL3
gy3aMX0iFo9hx+NVsKX3xtfeBe8S5n2ld07HVeMTH6sOYxk0p8L+nwLOZY/GEvh4
vZ3KPL1plveGQNhqyT5Mp5ImZATUKCqGfxDjIhPPw9H/0t52MTJLnUIr+YIempiP
FjnLmOw51dQe9skuT/s6Z2e6S7Kv+yfwGQF0eax5wUmgXT8hh/zvjmRcPmdXb2Bg
kK4nw4R3FFMYKoj5Dz0kGQbltLr6+Y25lK8oKlJjcAx5O+FHjL/0WIrA+2ZxFSzJ
8bJGC780SfbbTGbXcm0auSxSNhX9Z5Bm++xG3ovclUw1f7SJvBQUCj5Eh6bIMVaa
cWt3+LB8yYnwI1IWxBX/GAbsLtXZ/JGkooevggfDXrTMvlbCaoNSGN5/Vmomuy6D
2zcfhOeQ4pTDBr6fNJRkbkVtjzO3N+b1q8GhAN39SUVIdmsh8+LDH3PsHk6iuKQT
k0VO8IhYoTVI/CC4/0nhcBijDNNAdgrpnm3EYXfu0CcZqGhqTK84mQhD0/MZIlFz
HFgJeO/a9+r1DnlLT/sxN4D3bfbm2geXqoET+gJJ6UhwNqyw5j9Y4UdI2XwodCf8
Gk2ScU6z5DcEOQVPcxzBapTNcLH4DFmPec4m0sV1kGQ9/KEk0VHlh6rEZFegfakJ
IVufPOc3qQH4O9GhlH8YQItTfVml9cpaVWDU1lyaXACCK97epkpemKFdFc62hBhD
tmnRv2PS6Wj4Yq9JG/f8o+P07LpXkuxA2mD8FyP7PAiGtnUCV3bhPJIp5OvU9cRK
q+voQq+mkREkFDbUWZWJ1gWtCb9mXyC0NwLAIj6m0L4NPDHSDCgMBuXL2gMoITaZ
RMTrot/CGDHuE+061ffNvc5dIfetmEmNmACckcKgeDizAag0jrJ5Drhbo86/i1vG
L8jLcNt2k/P2F9vY89SeShT/Rsu6M1ezEOYoKbrqsxpivRplHU2WWWZ2JhLAdo76
+Bpo8uRQ/7OcCdUWycuu0ZnirPEohfBuw6RHQa2YzrGc4+3CtfmV7MtvGIjB59tV
1HctOw7+wck1vt5LnzkLlls/A1i5VUSpRc+9z14X3nFmTWmP2KUO602xMavlDLqx
qH8j5vdUqiFM2Z2tB/SF7bFkQ97AcmLCdOHpuv3HNXeWZz0p8Lpu2QDerDiuxcOb
YoLKXGqWPBxCRVqd+rFuqyMkI7fQxDbNVh4RsMR31Enj0MXabmxb/Y7826rnvg00
rZ1HPwaiu/+DRO7Vy1l9Vp/yOqbWrcJYRqvbjyt3NsQk7JWm/K4EEOfo1V20b7Gl
fqcWfvRUv6khF+pbLTRbS5o6r/MBJTM8gi90nzI82Rn0Cbm02wCmfwPFzKH9DAAY
rx72dSIF+Hgbdvbt2iXu3p6zHT226+VMbqqakkpnc1r5Sp9UBf6+fGPuzLI5PezA
4BECMgPFNcjSgb3YHVswy1XLEsZJcLJEwrl8Fx4rvqR5fwVkJ1AG/u/5TNdPEXz+
hVncBf0myHWgCAcAA9InwxbjeVCHXkbc5zr/TlMR4ZEOOzqA4e+R8G+QoPf3yQVt
6bWR+Rr80Ec3nrofJW8eVBSGgtnkDtTar/2Iks0PyKrZi1U4+xfVuySg5kny11eT
ulpbm052V2BamZaC3v+Vdm5wO3o96oStIBgOtMZ98fpAj2y7ndwKMRbkbjFdrPvh
DBNM9vjN9vvdGwEc1iS55Z8w3k6gUgOgYuAS9CvZbqJcnlOI+0UjWt85JIQVGVTF
/Yi4DJcJx9cLCTCMNs8ATQBBEHE/ErL9oGV0PZCaej8arTpjnDV5dcHWWFtJktwv
znYkv8hJ5PfkuWO5wKF3hum2nPtjXqfi/8qrkl69VM9IZqH59O8lriZki2Hq2ado
Fs0QI7Ykck2hGQTGfFRKc8zLerLgpRPbWUgvPvpRdEYlHJBk9G2NZWw/NGUlxHB6
TT9MAZxDIrotwmADkUYDRE5wUTBncTfkS8mo8BpJSzB076lhCk5Qi2Ew8C/jd0mL
6Hp4R00VC9gmvQU1ySPM4BgvkiclUYmYZYcDw+VnaTv09o5zcEeD84OjrziO0wC6
hZlFEqAf2sFP2rxt4wF1kuLwLOzPU17PjVggMu38qipAeI0dYFhGhdElZV146mrC
cSO6/85jLgJF4WzfYrAN8Km22aaFMCGMJedvV8buaHN8qc21oqjh+zTUbijOnG2F
rlJKlUf7a7azik89NrW8kCX/eCU3cvGq9Lq43o/oWVol2ySpKwxr64CJcqamsCFY
IKQ9QkBUOUseUA4c69S9VySroeniR44rM4PchDAjbTi5A7sRzpTekH5adGXyyQeJ
sdUWzcfYu44nflVTYO8ixgedmZ6EyB4Ae3x+dFd97bthg1p3B+3x2yKOOh2SGOoO
rt3AYf7m3h2J6RtesCIaQo4OWkZmbVy7UIfUfiwePsWLao0JUnf4tx6wPxK0vyS1
2LBsNa4D4cGKYsqUn11+AU+OJjAuGXSjMVqZO8mMyAEJLp2wD8AuzK5ncQMM+TpH
hS5o0vAYPMbTxUm0v815dnAKqANRZ2xUgSq8KdlZFVBOdf8XsVcI4ZOd0P3aClmP
47+iKBbklTBMeBYx8e0k7g/F6qNXgjLvcgWkHku3SOvP528yXPfS7j4esAd1FeIw
9hbVes7uG5TNJza+RSSc1RJ1kLHr8U8v0JP4o1iZYXwUPfuU+mQeX+WnlhAel+Hj
vl6REh/f71JwZjS/e4gPkOvzXQATfAwjNMcUpcb4B4Z8iJtZP7pWCQpDzzqnxAK6
fP1R370ganS+MlSvi+kelA/xTNGPpHvUZIBcnrVORd0iuSxuwSEarrHpY+z96scU
nfesMuNkQweWG8D6RoQwhllNUPZEHuBDCSLMFKi72OiDB9EmTPVNUBVRtZwNvryN
X5Ai5s4/sLk1iB/+vVCkLgghKqmrnQy6/lElhTFpc1VqDj9ZpLmyWRs2Q2LXYcp8
p9Eg7611Wxg6fp8mwPxrr8UDaVII3i7eDN/OoYfuu6zflPHdnudAcB7ehYr6QvdC
o1dDHIw00mCURUQZ5c4bnpxZa0U/sa06YsxjMBee3fq2hERECQPhcRkcLNKwwisS
Ht/zj1rHvUoX5MJluZBUPRpo0jNzvZmPTYNRzcK4QU7atjfEyIK8AfFKPj+/zwwH
lp0B8bZDeTzyXgy+fs/JhbLoRzk+ZfX41QFxQo40wv2AJBxQVuIpqSqqJECVbLCq
xq9KVBhtda9WE/c2OpcKBTkVuZEEKH5lLZ21uWcAZSAm8n8j9s3yoT1m5anapgcQ
a17JhL2s1LhnLOPhpa0jM0azAG3fsgHTAafMJfxZY/cY7U285+E3Vcdn4hfJP2EK
YNhIYEr7NhbxHz2c0nWWJrUgrkB/r3D1rzb/4JRUwhSnZfncoBKnEOIO8Z75to/4
7/lYnPZC4BZtdAD+cIl2VpTM0TgV6EOrhuwXPJMnlunU737d/Zzlmv44eu58Mdo8
XZw4o73ncbyqa0ZrK94dzYT2vC2W4s+ZS4vlp7lEdG2GF/NnuJqxEKfzODNbWymI
UgT3Y3OTwrkxgD0a44bqtuXda+sH2cm4SiNX6+5ZslCTO5okXISOlucJvZqeuvSk
SOa1UJRJxkf9bCJmYPXaLvwjXLlQU8fH0qo3XowM+LjydCr9YG1n6papP/Qv9Sbt
KqbiaNYSPW/uhb1t7kC99GgUcrE8CpJWMRf2t7zsoxVZB9l3cq6jT5HWzMoG5pBd
cf3JcM2eePWE6x6tm/15w39z80A15IBTvcJXRxkvwKvQ3g6oFw8o2LXKfQmmrGKS
cu8eXnUaBe2jlGFjannDFPhos8qkyh0NO5D0M2xasWyToejHtiF8lsCrXuECeXK8
FvaIzbk/UU7g/QDvXxjRCxMEhwpWfy69ujMrZNno89N4OFbLav29lUeTU57hBhsE
Tu4ql0LtFCBZm06A0kDvMu8nB9e+ykZJqHWzXJKF+TEijMZWrAT//8ZtVXSrM4dO
2z2gpeyKhUCcHBZTI8EuB/BO/cJxeeg2ltEBkDmNHCT++jjdg1CcjlXqqitCta0v
0EcTgoWkvFHPJ2BuASwQt+ZBB91n0NSBJdqujKKJq3ulxMaqhJ3yL4VlKFEY5lSk
Bd2wcdWQqFegscLST5sVZKi5+yKbLjt+3IGhSO6O/KP6GsVIvyW5w1fwQ2j1YrTs
R9b1SJ69SGdOE75e6RfwNevAa9M/AZ2B/ABbdWm/mCgLEJXJaGNVm4SEXlLV5v8I
coX6hIPlS0odM1gomUdj2jnv/L7vMsHMwrlClFE0hIjZqoKNXESudBOk78uOCC0N
kSPeJM2zZdV4UXnNG8sNMigP+nbpUgsnriLl2B0SyRKF6NkTA4LZTNJBNjqUDA/r
v04N9sYvPOC0TKfzq9KDBt1GHRUHv4hYCqWaoHavibG0YweeN0z8+LuEWtxzyAny
BOopQ9+8ivWbL9kU+nWkbssXHBlvq3TD1Fcr5oOezhejY3sWo/bnn04NhV9bOxRV
UNTgWIsWM5LPk4HmvuG/ozrX1jGB/pTZZS1uSX+Vo0ueEgD4ZW3d7J9Gf9am7bN+
1G3Y1rZuDLo/+PUZekd3VK0t+4ehpOPcfFOL9lgEl+QhPS+Ana9VyqcJpw+mMuHK
D2tZhfnGMeSq9nUmkUN6e34jdHnswhdku59U5HfoNGS+mY9PH3LxwGdsifFgxgGM
k7MJpKS1X1XvngjIw6elOjRLYdDnCVw/pph7ib2m2J1g+zzfwU8n/KxGhrTi3kU+
yYFcqiKAB5qxjV1pIj2JntBSVfEsYeuYxV77R5n3Z51ppXPgFOPjy19wtvr3+YEp
acN9+Yq66GydEgjnySBN4vei2TtJAgTRqQdldoUXRIx7fm6UgxM3tWqtHSAVQO2o
cdiL1XG6s62/wspKCyrKKBPxeT59nyDA6NeO7GJ6Jfp2qZNDMWv0aWO+Z/NzlBB/
XGOrp7Z1ssDYPGikHz09RvlYCbh7mTP3RfnQVZmm+syX1sWIzPlf/y4ItT2YXCPI
QSETcWv+L8Rw0+TXcV6PGsvB2n1CmO1Se/jxCWtk0r5KtIsPYvyTIMjhjIC3yob+
zMS4ZNmZQIKnorSF9OrSYRRqv983urh13PNW0Fprp/98E08nHC4T5Cm9ntafJku5
BY4VicnuA/plye0ybz92qTQ6nXwNArQjFOXSWSaqkNYVCpgCRj1z7gwZsICvhN8P
HpkNZ4uxaS/ya9HlW0N+kKHIRWIIWhr5/GAPYCs4oYcZaYoHZC5uyq88POTcXUGP
O6dQk4XGw35jkL0IYXxHQG7x2Er12DxWrwh7T6PTRFYDp5bT7E/VLQnwT1PnZbFu
jbAHEWhMd5QU9qvrAraH4SJ3aK0gH/tv7xiCzTDHQvuX/TXTAgH8JsCzlXDxc240
+4i1q/ZrbFCMBbw4e/t8Tm53H5NhbwFtDAMY5Er07h3H6iVxklIA2zFE9Kvic8g3
gWc83uGQLtR3KlSkwuebcNmjYyAsOIkREM9TRPQlhyTKFdxYYLO6uOQJgQ2/4mcl
+Cq1+CgeIcu2FLlk9SXcUI3A3JPEU4cilTO16/3So++pP7Ba9DgDuaRzrr7kDRGW
vf3TyEx/+2M5NhVydb+UGFy07rzlFPOXbA4ae2GuVnp6aY/vapBmQUkmYQwnxWNn
PWJ+6quaZ3kK5+JofbVLCPpiKRoeNCDD8LAV+hTWAjB8QQ3CvbWP3zyeUs3flu1D
FeUH3I5nPmRCjRYUcBJk+mwl07/NxRvkFYa5c/ddLSO4GcBvOMNvzYP6rK75OjAn
TfD9k2fh/6R1UiR0Bs9yfB92138g+YK24ApJo5DqaY9+Oh705ttfwURGDF+Xn1a4
y7EQ2EyGLgabYqbYF5JMjzAOsJfmoNh/raJlnsqNK+iFuY0y4723hIA4Om2V8JAB
Wm7iW4zSTJ1X5BvysFlFtdBYKRKaZm2tweZjWC817iHp9bBf9t9UqUexq/Zb0iiu
rrZtLvufhh3eyq8mTgCobpwpanS4manC0d7l19dXi7hMc1L0skI4HC4VtwPTbWJf
vdOPzcwrRLkfa6+ugMz3p8yicczR0/qFWjh+XVgM2lrDplZfjjUKGBgMy/uFyvB9
ZWVDbd2RfHenJCxIv33wmS0s4jy4SZtmzN0PKtipE6dWWl5zkgGlqzdw4f+nZINP
MHZl2ICLMx2YGFZblHrjDrFZTTndNDtP+e148GdMVMNoo70BEtfS5H0tEaHDBJ2E
fxWRetr6y9lPNm19swsWnZNXf7fX1MpYQT5M5okiQ3hC8F/rn6knlNCuI9mLSCtj
TEqNgyo+aQVL3MnGdoXTrLTMK6Xv2xSEemlBdhGoyzIlt0uxadxw+/31oluiz1UC
HHs8oAL+ajk+NAwwD6jRKVrvXMCtTDhAkyrfrtHo+kqMJf9IN5zKdrYIWq0NrXrs
sCmviDn+b7RbQg5/x0d1RSffB6YlNe5aswJrJbainsO5sN7RS0kg4jVjlgdQOkPq
RjjuatKtLusPpks2APlES3/4bKTwoiiGLFCwbx63HTm0XxIOofcUNNZpCa7RSjmE
TVGfyCY57aEf1L7xxl4Lqs5nxKsDs3VuVgCm6h6841J0VWwRdHkOhae8S1LjqP49
XfW5Epi498vdupEoLeIbiHF0xRe7CF0xco/esqfrn73SwpAkv/uwwtCe5vz5qYgM
LTC9Sqn+HQ3KKCNJDYr5tAjFMH30p7qnH8oxaB4O4LKgq4y9W+sMsYY53Aa489rI
osaxHoBRRiHqFqoaLKz723Um+fK12RrVPGslclYYWhWZ3IFkP44vzfr60Zi+Wa/n
YwOQiSMMr4lmOujn6I/w1DY3zUcuqDQnafsjVTUno2gkjWYGl4+o5vJURvv4ExO/
h8EcTFg/fB90gDJtQ87VzlliPSyp7np/4BOmEol5lnrfNqltJDwPbF30Yo+pVK4z
pm6BqH7RibYBBnrL+XD8BCF8/CjWQGaumtaGY1j0V5SDYWHNQaJ8joQHoyko1a9I
Eq4Xi3XCxs0n/XsFCxZIoYpyJyu/Jbx2fa5T2AGMdX7XKWPufpvYJ3k/3CC2fSsw
T/a2AHT8c7gWU064x3IVBqf8zzFsxadXe5ksq5l61TbW3OuwlvC/e+j3t5eEeUl9
RtZILagskhiqmAt5TTun6b18k4uha2tNETDrL936wYCAK5xFQhiOcb5vlP+xQbt6
+dNdDm7P37lEdMI44x7a6ntp20EfqgE9GxkafrxOw06YAl8XQok/DoQY1v3WnvlR
BX2K8yD/8FM/ci4zFeSm9+2yrvFVJ6VqOteGHdd65osh3cmD+7QxbZg1vY0S0gcZ
KUKjywJeEgSreH7BZg7lQdAo+xaExCdPoqTIAL007WT+WyGVoKhKn1jMFLLpQ8pz
KwjPKlmVWszAYYKRbgriV0UrcwV3q2pDIlR8w/f9XYCgXFQWQQFhBmkcOyM54Xvl
ZocOs5/IzrHlhMxzWbf4pVeka5z+lHfvH0m2ocCtfueOAdHO2LqLEZ1CSFsJzOmX
Q0O6M+Vvx31sKpy7ghRFP9AGLeEodKcnowoO6+O6a6fkTEFFc3VLcR+/L4uSjGIP
FPX0LhNRERHbwC4mk8bjvgHLV5eozzpTa1cXETGMK56eMnqCPPNpRgTHIDiQ2CSy
gcuEt3y31SPIscK649Sy6TzNJMlVtRufRmOMl5xmoW260jIGTIr8Yk2qgzoZcphb
wT+sG2CxBObJZpuoNGHHQVFPisdhqbErX6q1v0FtlCKGsN9bDDu2c4wOBnJFTJEG
TTyPav7Hu3iuq2ckqzZfmMPB6wfXpUCeP2Gk4eepFQDHEKtRtWLJHGP5seoCPPoR
TfL3tdVe/R9KfeHbvOEaJE5nF1mIDkZv3uzbhJHhK4oV2c1O18UZoEtDZn3hsmwR
eTSvvI9ERtid7Mbo+aci67LNzZ1ce6DKHPjOQskrY6bz9bFjgkHK34T7ox4tWujy
iWSYZ6qgkfx/yckceSpXLXXLZ1UytAxiUa2RhkeydAibO5IObTrzRYV1oZIE66hx
Dpysb0RxrZwNNWTxzebv8QafOaphuY8gW0WNCm/nRAhexzenQGbBiWsLQ5Fmnom4
8RvD3/VFykv4/MYbrrJrTfULdzTmkWH8zekqTAdECaOpduibGBruVMW8uCg0XT5l
F4oWeYVEbzZah+WvOQIHCEXYt8pbzNxzw+XgS71s2iSXbxXxCpOjwYMhFGBFF4fH
zrd4Phaz6yTab2dFBRgKYY+c8C5Ufo1Vf05BUxM5FNVSiWIEoCtuG22wwmqoGk28
VbVXI4JjWHEPaPQ7PMeCsBISydPXlkDJN5C96fkzJH1NYwvBG+xoubhwvRpHSY1U
tklNKLc8As49w+9MYF+kUR7wkNWeZxizcbDCTHEndEvV6AgWIgNff5aVzb6Bty0k
19uM6+Ujrp8AP2Z31bH8TRHBR7JhG+6bW6W2da+fTrRF6CcrBD2nOH6t62gtzYPi
njL9mq8/s4jc36aFSNdrUFIT7wFxtc2kc8lP9DdtSD2+U+mO1Os6tW6Ucb9FLekv
jm8mP+370e26K6HhQS07Zkpg9MIILreqwUlXybG67qyWqQqWbrJDWxAFMwz/SjLg
PPJ0OrWnQaBK4HYw+4ACPPPudDc+gbt/d5pMvCWf2QPbPZKZxabGubeVRJkVKadl
MZhZzfCQtoi4UFOnAgHvEIMPbWHE3U9xCQHrkg7TLy3jE/WrtC2Kl0t4BACCIe01
VWvoxJvod4MDV5/7U9HmAVkW4BBN+Tovo9/VP3jNFH3rRPeGpC1cbXq3aZrwEttj
qi6iEQKdm2kDJkpC+j1tswMLZO/WiH4BZJd9nrZUNwzS1VrAPGY+DqIHWgfLR0xj
JAUq/qjtiwHFtXFe+sC67ZrUQ8HeRR4y2Edf5p9D3IgKBwIvdRuQ5bcuRH9nR+i2
8jS/ajOGI84ZDkqqhYoBaNOpFGvurKj0Gt98xmMNYmG8byyIjp1KUYofV3Rw87qW
78bo2Cf/buKFiAtAK4SQOPf8HZdhkYgk74UKyHNgymB/T+ORefDe3uW1xgr2TYkv
pTiwyt8zzlNR4+QnDY0FZ+fkwmpMdZSwD4l7F3/QAUg46BhnM+h3LBVFhNXnQAp/
LVHIBQhgEADqrg1GiwFVY7rSK8CfTjlfnrfoz+8JzJWnb7AF0QLxZxmN0Ewfc9+K
FJDcbibRCLmP9MMzVGTxEfxve28AiVCsz74NjB31HmzE4ueRH36R3hsCvtt/Swa4
0vuA7UvGexhl+m4BQR+I7/HPHQJmV/ia5jfsAiemYvhN5jRJubt53gKygXM29luR
KQolf4yO+aAEKBTUGqJalGkneVNRHq5yACPkACazBbSwyubA1haBjbhn/hc/6wm/
xT122qzyA96t1htbo19Cymb1geQD747imnaRTgFtlsHHHGmxRJoITEOD+8IRkn2F
FpdOvHmv00dwi2j4LqbMHrvDkRj9ErBDcEdBfQocMGXgsm+xMBCrPjnShbmsGOJG
VaRiP8BXyubID0oOnM9t1ZxIi8ZLpU6W1LrdbxZe8OmjosyVn05pC7eDTkZf0Ch4
VwBvzMv4FResDIEdSZVpstAT/zkeLe/8SdD85Kqxbq3sa+QAdnjFeUhDIqtL1A6R
mvxu2qWJyY5n218QXhOu7cSeUttSA3AGK59C8zZHApCzr3fNzkl32PchmuYpb4zr
GbFzFphC3m0NI7n/FTyPI6Jrg30Mpb2dhJARSU6USWIAbgoBrEtL7dYcf7BDQT1R
8JGvR3jBSzDDKPW9F/l9UBvn4P8ly+5yWoRFyOqZPfUYoMkvxyYQ2gHKimme7DY1
nMqJ+yHM4leNlJjsoKpARgTIBbhESgSSdqxHh3pHSBJjNZi3S6+Y6tb4EYTC3V0s
AhkKZdFn3qkPA6z+DDSdZGCi1rdAib+z+zt0cdezlVHy2UP6hzcTxhXRGMKlFzen
wGH7oMVKNi9d1f2/Exll4SK2xhQXrLeMj/nKt/cFlcw99i1Ry4EUmKjIB8WzJh/X
EY6+QNPD9AVOoEgc9gKSyl3wvftHwLIpTIUPRJ1iClUm4P/W5d4b40ve68CbzUO/
PzqqdXJFxGqxQdHuorTVI4lOTqZPK5uvjUA6rQTz/SsK6nj/AImlRYdHfA9QWso2
HWkDoWn8wdA9+2aboohYLkayvRUZBSmy3faGABDbHgL1K+2BKz9w7sK/LEvUzxlk
34KUcLrovUOH4mHqxIYCqyFJiMYIQYt/QctlHaZxgPObgXKZifIMtqkIsDMlPPHp
BP4zSJpK7fffyLclLTnseXo7iJGiEoZ3tEL9e3wJOLGvmcYiNEgu/X5LOBzUrLBy
X7IgixtNpsayt4iXdG1fpMfhKmnRP/qE1eRnDYMy6s6v8dpbClTb1W0wtwsCPFlW
DBIrlaJpkAw0bCbtXuGfpTKzkCUHmcvMGebH1jyKp2/FeOM2VIjlH90bgd0JPj4q
MlJdSj0lgSvep9xLSGelpASTog3aN4o+8DSQ6T7jwKKnWkxVDSDNoRrUcq1DVQG1
hty4zYTFWe2+RKDLsCjJfp3D2+evCKRust3e2v79Q6FGo8fWbeumVBN+xaOM3VIt
owxrWTXkSOAGtcQFueEAqkbG4UFfm7mKiXABCszhzdTf/e/vPsIms8sYbGoqUhuK
voN2jHmbcv7b3BSB7DNQlm+d+pKg3YpABD1kIZ/uaLTO/e5JmXC9eI13tQAzOhKN
8MdtmpT+gc3//q1wXbMfVdGo1PAo9LRySnH7YjpY+98Ifq3kyWrDyLkyNx/3g8PZ
PPuaJ4DIoSgzRnKW6T1maOhVTa52HmXADQN7DATWOebrIxraNLeSom4rIm35oDLd
xvNovXH44W0TKzoqNrri5acrg0SwZSyEoEWCd9MvU63pAlCk3NY6HgNcOgjsBxjH
l2RsMJNu43X61kSo0q6R3kvFIFSBd/vNk2YYzyQgXgn4yv123QOYJd/+OUBN6BFx
OxE8BKKGNZ8R3CwETtd6m64RAEtlITS+1xM8hsylcOD2ELuE2ltT45UiRDG44hPM
KVMcr50+iTnV7yf8EUr6Q9GoC2D9eRA72Gv7bFaNmtwe0ki9LwOYpFnONjSFZrZ8
lZepks8J0w6nk1LFX8UGS9LFmQZ/wKCUAoUs7OyLXKmPdePLnQ5eq1dKo8P7ZDVd
8fDZ68uA+K8juDZdxkY/CwvwZ78Cp2FqMM/FlGPK7KdunXwWUrhp/mSB6xsyEInd
gijT2oc6q3YD3mEGd4mNPAFpCglrG8IQmqSgtqsfmscswI7DiUGe31GyDPjJdgS/
2sMpam8KRnAk8sKul38OFQpqmP9rB0jXEwkuod5hxP0/PWLwl54alwK0FvK69jSQ
wKQH3ZEnB/rmc2YqqWmuAdfgJ8EXRYlmQu2HUbfxepRqgzaDATbJszKkeJmoczY9
qAnmaJTQYbyq3QwIYRcXiDk0kjXZDgFMRa5V2FbVN/9VTuTdigBl5w+U+zoyzfao
3q5g5HNhhQwXGU/Qr4ZxZxSsWYbL/Q7qgd0zR3/Qgov93c04DgXLhrl1sc0nCu5s
OWg6xsa7ak7sjtOhOnnFwPx92LgRMYrIf2Xopnl8dJBCA+/Trq9Yb7wb/MzpqSyA
braKOHaHN+IYZYdxhgpKKShFs3L9yULzKMaouz2S3WuCTAhMf0Wks8wiBX37YDPe
KjfqgElQ2T51mbFtjB0Wxbp7xpCq74w4HY9k20fcBsBYIMZaUmmQNfaVtV/EY75G
+FyhpYl+6TvKpQLecEOjGoWqM2HlsL6mszYbC86N5OkIepTdGus5Q0pQxQWf83Lh
5h6B5QUvZFfEFfIiI2i23PE0WJECkiXq73ci/bkUMHL4xd2O69hdkgt+H/drsX6C
ZwzuTWnfKw9hYd4dv1XYreHmvxcTYE9Pxny6AynovXCgnwuTCJiCUuOptm9UgXEw
NpazQMkK8gUd+6pQT3jxX+EVCAl+s2fZlAvqCJuCYNYb4YORrfdMY/CObXkP/fnZ
Wrtt2Hu1rj/s+SkXqMCYWaNsX8Zie/6DRzs6Fr9VetUr7j3Z/bwdAvckX8961AJ1
v2qVlsD8/J9DYp3tsouxZ+v/KBZaCyrlS/QhD6XVB3l5Wh3SDWMFvCxcx4y4oNLf
5ySzsHnVfA6D0idUbbnr/NU8DYUmFfntteeu6YTEc49Gad+XmvT+aYOd4tA9xwFT
m29ixsCuY0weSG0eUmqiHBM2pdSCO7ZwBGLF2IUD7rBqDvZ9MoelMyjwTbkQ44VI
j4cNSp4Hl7w/bp0qDDWdON1ZFTDRZs8wMpcy8fpvHwkqoR6InYkzHbsEsZ4OuqE1
Zo9gXYhPRzmMMrfSWzs/SDnhV+IdLVZDtHJFzeaAStQrPGTKVYD0eNcJ5jg/0bmK
Ot/WpHlN8YmSDHehXZJ0qGD4fA86LRk4tku8ybNd1NRmSIdFWajFQK2JFg4fByp1
KV58HYebmHkTytxyOEppCXc1ay+Ckxx1FfC3k4UgeFFoAMzpQhjvvkZaFqE9T8nB
rFJcZzkIN2qhMs1PPQEaCyk9TAgKrAF1Xm6rdSR/GrCs9yji5016S1eW7VLGecFW
/+EpglPWEFZEfiSCPMlyUSAaUrNPrKlaRXRIu+C5jeeV4d11XjZD+PT5gmxrTJ/R
+LFmVMoUP4yYuGznMQtfStLbZydrlfn2f6dLfIiL26bCCrZvCyMMLUf6Ud9Qy2lf
ULIzsgrdjRV/cilADukoa0NaR3dnLCwUn77iJ33GjrCzMsT1RwO9FOIDyAKYq4l8
sWxg15QFQS8Pm/4LA1yTlW/r2CaixRCZhGm5PJQ6yyUAwK/tp3pher6bi18JMFSQ
ZuZavr3Vd+InIixXy2GZI6S7WKRysMSbcWZdvTQO0nPyUgTec5Q+8CIhjG594a5h
ptjJo/NZ44rKpnXtdVww995C/Q7qnCUKECp4R1P/+FNw+9rPU3ZOtPo649rzI6u2
MYFtP3sApMmqp+SMbuHscF24gKy6I09QLoOsxqB8vczRwogPk2Kci0X6vdV4A+s6
zoYiXGuQonMZVsoLj1U3OT/XF0f6zCvfa5iz+5eBouzNPlHlnanz+IPFz7FUlf7J
OUTr4uKA0u897USQkAsXK83oIkdNRvAM2yewL8zYRQDTRqfsbZRhJqZ/vRBO6N6W
nhxyT716Hao/fkpmnzRkbRPWyEGZrFYdeVnsanowD7LczAoiOXulzmwqTKX5BK4W
rVh7fUS9JEjh9B8yjbEyonFjrdfubGuQt5GfRSfLhK7OInpJ8EJeAh0d5T18YIJg
9HZ0piob+5bScAThEADuPWnFwm0Pq9u0TxUn4MeKRyUTVFUSNZMxcSSEECVc66yQ
u/jcdESNMX5b+zFm73yA38DbC8AFHGC8WNdNNZkCE8UBMAvAWwsJZ93dVt/gNrB1
wKGrZ2/B5+t+st3kPsu7l0J1jSW1KDMZ4rlYJzY7kRXS0n83g2/xLR+v6KMB7PWl
AgwIe5AlcKY+Rv0L8nvSYn7xKsxCsGFOCTu5CAnlByN342Hy99X4scoQ21X3LIoD
YJN8Ts01wDo1aYG8iXsiSS9unw2WBaUfEjg4VWjwwn0pbUwdqoNRf4pH85AH1hD3
evkm+GV0XiRDCJxfPY3svcbd2PCiqK9cDdy5Wl/cFA9x72uORlTiCxIQnmEO5zv2
S08UQCcNjkgTijT59sBZtgYBvjqKKdLyvxIqL/LhIB/ZhRzTtK6ieLRNdQWy9EFk
cqPLvQJM8rJgWJj5W2MBBroNlqNplaBL98NfGvEpVORf3UbLCalSHr7jqCtYJiDj
jglmTyIMIJ7PcX4D39fQ4XKiPQTABEYyA7fCh7S/Qbm1RqR6niY0fTIZovGrpO1b
dmC3saQFzen8UiNIhwQRpnnKf6GIqOxzhMdpJ8TS6erGWm4tcWNcMzC3AEUysFH1
klmETVKV6mIX7Q/x/nsLT/D8lvZobvgAwCVucflUcm/fXqjeHCxVgF2RkGm8RJmf
abM2jpQfjUnBTsQpbrEF5bvcEwSSv0BuSzl48FkXXxShEm3o++9vnLuaTyJ+IXEN
wIYACxUqKUxZoYvHXftxUK2sA5M65ZrqTvkn0nIsbBLu8cx89Qdkm100Mzdn+ITM
ecRq6jv9IHLK+zAmuR9cCc+4NlqckDC9U36GH7L8hTOJup0JGx4wlpWxR4n3/bh3
1Nc1/ed4l8ngiPI5dklE7/jhw+b5gf9wZBOj2MNLRD05rR47l8GAI3VWCOxoBq9t
6J8jcT9TcbMrLBMYC2DHMHyIvdWzfZ70TU0nCnpnHTRcJgpDWxjSJfA5w9AGETlh
pibjKf/6RR7GCziXnuQcoZuHu27HEif/1cP65HcLxb6RYI0c4DzaTtIK+4R1SwXi
NnR+TtaImJkyrbbXevAAcP4Y9qhktEKjJoDyJGaVm+bimGnDle3PqqAxw6BIGLOX
6Tb/CELzcZtIYMBMvl8pnm+CzxnIx1vuDK/wrqO8hR30Wz/sxiXxa6OKvrqMbcmr
6LobDpdhazbVnGDpuvVWY392WVIsqiMCW9mk2qEFhSWSd328fvsDasWwqY8DkEib
7E/RAriV5QotVcBxosSBIZpqNFDppWJpVjmikwrNbIhEUseFvOfW9i6NyUALhT8G
FX/rG0TkIypmoHoN/Oa/3v/LH+UvA2auX63/XyLCLcP66ofQqbGnkk8j0V3D4KXs
DoAzBtj5UKxGp2ds9iP9akwxSh2znrNxU6j6dg25zbjkOEt7HDP7lwVUXKg/TEJG
pSqAKpuZYVztv3R7p1NbI1vQCCFEYajU011snM0aQnW9SVP3glsw82Ru6R4P543E
2oL7oBxCMesbXmUgI5je8DAdRzs8a6leGEI3t2Pc1UaUXtGhJg8CzN5TSr/+Nkzl
mIpWtS3R1lbiZsvvjoCFS08631TYsH/OCxF47fXsKNVQW7nNiu46N4kx5CGPCulv
l8ry0w4qkSy1X9RqnuKgpkt+txC4inP0CR85hTWDvAqhsVkB7uxFTWU/wVAnTP1q
xK44pxAkC+bVq0QiO3j78D9+mAZl70igQCrCEJSzFtCO5I2Dxaisxy2pYTgzbhqk
MVTAW9NuM7a+6axb50zyKlDtSAx3E9NvrbrGulkxvnmIVSaTNh7RBKbdmDEKhOY5
lY44AdPKWaHNlA0wzFnw/EDhv/UBH8lek+0zEz95mdMizZwHAlJWH0jDlnqacAWK
LCzFLZZ3cXdOVCnafAUW+DkWvDiUmhI7ECGKfr68lEqeGgtFJEif4zkhwKhHUfv1
DlcKswlCODVHSgavoSv1GLfX7vnWt4g+wBD1xMjig8wExwvqjQjwrfTM7B+8Xhuw
YEK/wzhJV0blFJnOorOioYBPIkvuAYxCps5+R9HRXTQwxQcezRoMM15kbajhqcu5
Ejd9ghbDp+iK7glSCzY06aZ+em5E+NMwhfJgbJ5YuUm2bpFQctOfnDcpyiP2vL2f
97hrW/UI6rEF3+Mo1SbrfmfpBatI1efPsMHOy8Lb0UZD0dHdZDNvdb6peFQLXhPK
FCR5QXgVI4mWBAXMTWs2xmzx2eM3vmCBUWGKcmsyrzZ4kQq6EEdVfX0synvqBLvs
HnzXKMj/FZOt4ef/KOJJJWL8C2Vty4Iq9a3J4SmnKJ6GngGWd9p15Lj88G2Ak3PJ
Z8NCvzUxOtLUajd+4n3EAraQJirkhrsft7Q63TpDOS++y36KjGgtc2HuYvGxPsZo
190yzH7FxpLUT8HBFWlQ+m5gQ2nwQv0yci/D7BetZA8QypKlS4FBT+hjCZFpdKD/
e+sCQcGRkhYAA5F6aLoEyB9UawVB8fYxdKbXdXZ9RbqJ0YTTFn9NG5U0VO+Gxflb
brHr3GrJQt1WbyXtLoP1Y5GKzu4Mc7U1inxhkAQGbpyttZKIHjDeKyWNRyH3dGEM
c0t77aqvZWDA+9TW8Rc4Dnq6JDpDWOeuA44rQw6hFqyNtAJNG/pLWCYm+bEzOd2g
UtBsJSmEY/ENJDVmGNB8gx70dhYhH1QCQVdkofAFuhBPjQgWp930aKOYzghXvufQ
i+uqnjM3xOaoSdfiyr5kemuuGL3TKIUBQyFGTdW4PgVzPTPv+NOANbzzZBhKx5+j
Q8DV9Mk9ceIxYRM2/mZGIMKdsNJpTcADo9Q9/AUDuRfrm7k4CZmGjWjdV0+presY
vFjbLTp4nNy5QsfhxcLhJpcdVEEI3QUhoIKFOp2/wRAczxdNoJzgyOk3Mmey1PdR
0hkpiB4qQGQjTUQvKy4hbSDLm/1BiofSz4OcXTHw+dScOJIgR8FvzNta5apbjXbT
m4O2hops2/aGQcm+xffGAGthsqpPQg51w4XXzPRjm+XAfzp9FrJlceYa10T51cs4
gfd1NQqk8IAlwOyyLm7Wz6nc68pSzV5aHsYXFKP4lzXimFVQcvKEknO9U52RltMy
b7/vmIdSqNaPhAW5Do91NrhXYuzBDBYcSAU9RfXGPNzjSZ/peqlpHpHvdQ+pbJ59
d8cKtfJiStYxyLIuIxwRpF0URO9kCL9zpHvbzoIADagNTVLKEXeNmCFgQsG6Lrp9
ceoEh+XAaY8ZdjI3N+HeHgFcONM1lIXyCEFP8oCHihnrTMgeWwCaizATAxJLhs0c
p/OVoinn60H3FQG9TDJbumOFCh5+9TqVZaGjDA0AZlY3ARgZEciyFe3PsHqyW0ky
ULEWGE6YIt8GvnAqFef4jyVPKF5Wbbkon+9ZonI3YGQxPrtqLGuDW/rW5X55lBAQ
3HoQDDfTjMWy5wT9Ct1q+e8q9IEWD2OIxD/2KJYq0vLP7Jvw3ehtjJuD+v/q112z
4pYdUk2vHoY1pBCOkkmDPyxo+MDH5BF9nsqfOIXiLomsKWmvMgUztXUgIUEfHdZ3
tlhV8egopiyQ/SFzUD/6Q4SAv+i7UEUI3uADEaSTbDdZ+jqWdlDmGd4L6RtPeish
AcHsYhLbD5JVrsjjomAI6xz8DTwyf5gv0Wwt/AYSAVBulgQRyRHyqAHHrX0j6pgy
i0MO/J9605/zsrVGjRB7MZQ6fTazpWKcYETzPL5ZGZWJpvARaBakM5w6hl2EpCFl
Z4hNKwHVGzzqZxqplHbZYMym4NXHLQdliSvaFvzUV9NKndIHYD0IXKFExDqauf+/
htAjoxEnSaQB5EiWr/CVm3YH0ICQ+iXKSenbtO0Dcr6XTyXGn/s4+dhc/qmT4j23
QtSiKufo5c4Bq1N9Y8q5uFnA1275vrl/lONRvokQ/jfkOgxZVxgDtwtqUZmwtby3
/R6QDJOxhMqWbMnvUtGtSAhV/HJ/qwbROUZqc7RafgNpUT3+o+eosLmNvZBxeFIN
+lU1D4+vjh/SBqbqyjf4uNQYBy8OiCyIDyYgHhKNiIzAKTQCwk49sbHy5bfx2jwr
4xZPHCCGOaEJq6a0JZWTvPqu5WROJyltDF3RQe4aJWfwNK7M8ibjzfvTlE71koLF
FB9rjTAgmHpaZfzUo6wGO2PTRVTBK8/rLbRcsNMGefDjWxDII9yaKaqulCX6gf9b
G+7WEtPZukJPF7IX8pTJfabnYo2FVcFEGJ+sI+a3otLeVSjtJDELw7ItIKciwPRJ
A8xtYIpg2xcDIH5J7/2+R3oyyANij+sFo7UHDx/J9LbEpFxqVoJu0HAabqeQZiz1
Vxtf+Gp6lvEuU+g6W8wFWcMpbIya1NG7wpGWbwg+9adqSI1st28JyLVqXk2DLgqL
+CPIUH0ogYgP2c5tIrjOmZ/iYgnGxczy74Oi3SWoGih1NN3UqZBRh/m9//zpgR8J
SVJJ/EdcdZOKPKn9nFhSjJgOODI4xWt9OUjRxoxH3xc5eU7Fe3Ck4eXxfV6+FKS7
RYq7kJpxrOgyJn2+oA4JcSvmJQU4/1p4X3vRDfbJ4Oo2AAi2cRr5VllLn9rpRHEy
QqpEF4v0bXS2XhRpK6OM0ZtL8cbHP9y4+Xk6tCFKy/CvhJxQb/0An3evGMIA7Gie
OIRXXhhi3Lac8hb3Nt3m1DwXMET77vJQIk5qXS0RrIdvAtPwK9k2YAtItHwI+B4V
IyQ4CyNiEtr53iSWPKw0H5EpSo5O4fdABIte4Nt1MohC8iOIWBl6zJ2UuUa9vald
Qd8AHFys7GQqilvics53VYIMJs4HixEuXQg9X20n9VGkncE+8S8z1IQlFCWkSlsg
Z0NoWDDdfyDauMAHXAntb5cIrajKbRAFQV1Lv12TmwVxPwLWECyml00Y3FZAt5yS
dcSTo7YaHv2HgWgufzxocYGnt7wxvHyYyZ4lTNF7shbgVccK4OC5jmDNZLCiRy9K
je4ja97qHQNWybKS3A8WQK0E6CJFIdsmarhLQ/QWRX7zP6SVaKrExJDWMBWOGmhx
8N6w+iKnpByc/UMcqGSrvhkoybjtZ1ZCUK2Tikz9+7SOxrXA6nZOkhEjLD/ramMz
XpXCrznFUvm5hxKFYsBbcIsHvsAoYUL7DRUJqYyVrC/gDVyT0+nYiEO/TX1EvEFI
2/hYYCL0Eq1QpMfxgqqdcOcXlNbQ/fOZw9iIn4QYeXHKxxl2hZDLvU1H8OKfgZ3m
FsxYt6WHo0N9Bz/Uv2Xr00nHJ5nkl43t/karRDgv8bGl9feQuxnIkY5nEuS5eZ6o
Apkl7QwQ7lfyuyakU1WNbzl9HqrAVWgZ3pKguC3SlNL7hZ0o3/K032qUkc8DlD+r
/Z1DIRkbYmHB6GfyW16Afwq1VHeBuKF3iol9+DEROt1oTq4ntWzFv5dpew64cjMz
6Di/o5PWRwcb0qsU9tQibYXe9MP28kmwFvD9bQWTI03Hop6Io3rquq9E4zF9qmml
YM5Jm54Gve9f6FiwDO14XXXI8t+282imgLg+mLf6LS00bbqDwD959JUAkwBdWcG1
uQ6tXjM8QdKD9aHAA5Ftma+0dLYxDNPHHCbDwNSvgjS0XfTlSxmVCoKgTv5HRTv3
AEXcrAznqEFRk8NFtsmtticpLVhJRZ7lB2zEHV1cD9CJzG+oPoC13Kb+ibbxVrwC
IaNmD9HixYZwpy9oOPLxClbdSraM9Ru60ek594K5oJs3RZrytHjKxcNbsIyWKVSm
X/y1l7HiUTexN/9GyXA/XorEmlo2XpxNhlgldEt0/Z2p16kyPzcQGK0QdrBLnpY1
LC1/vNS1gGMY3KNlzjmnyF+JppPDO0pBFUiWmR4ClTA+fD4UqFhc2b46zX2bqJCq
u1z2KNU++sKAHFuvJTjfGNaPuW/PNN/Di+NNswyKH1fOtdAbqtiSUzgt1iQwRffH
ywH80lMRLwRnyX5zo0eIIEf5clGgYC9PkxUo+FubnJM8sASn3FsPIWXAwEeOlspR
lw8/Cxbs1PNLbbdJxOt/7ceSZQS69kQ6ZYQGQnZi1uC+YThUy1R0Fh8VnMTcorAY
7bU5iNrYAUuSyc0VB4Kzmlyr5qsI9CxQGGLRuz/Ya+Y4rRFswAHINVwNMyypyCYY
bMKYyKs+Ovyl9yA25M98QztfBK0ChrHzPfK0gG9dJoeGfG1Fo3vZ9OamC16qdn8P
6rfl+fFmpRTac8DBAmsWvlvmTsjHoeJ1ENUmdwitqnnDdbKDvUyHL83u3lkUNcCV
nYRFzcRqRNsQPFd+s2dRJaDCJhuOjZq2UC0rW91RVZW86xHNn5fK8gAcSpFf22MF
oI95SPFo/lthm3h690++I3TH0F6Q6/2OEjihu/Ch3AlNNge2RGmrIa+H9Mr3zxH7
j+gB/rfQHQOy1gmElw7Ba6be8/wB15JQdsdS9NpZoGlVSnao527bKitpF2zXNaPG
AC6nBjV0hzSlyk+wMHZxqQBYoPHTN7HVUMZra2jQoNet+87kaIywMufl2uTS26+I
Hgu+0CKk/MdT0r6qed1Hqxr+bRViEtmPKw/GG22rbE/0DgJ9EjEI7gdDseFXvQg7
7sXHYs7m2vUeiFH1PTiqj8A1wB6nSr1HP4tFeSCvFivslPzUWAyGll2CavpT+rUe
JhrRg4+QquczLHQL7xIXaTUtkgDTV+oFNDz8pZOaaTz56CCF+sGyhBNoExPlfT6L
YDXtcmvKNHzRcPZmVr7YmghbMbPgKbz15XlKli9CDPOAveuW/s0RbOFnsAjMCQK+
WKvtNF3BEVY9gOzZ5TolDztY8A7Xq3iFIjXOi9pEDuKyYBGczVih+7K+o7nWQg0/
zpYYh9nFnFPZSa4DFbK4qrmTquFJUq0G9nQ5vzlKkMNY8230AMTL6aPGSsCaDcoi
Q21Bi6nyjQy3v8X03XH1qNQSWHXHMPDIA/8cYR2AyB4pQmRTSn5qrSSOl+ZE32wK
WnM6EkAyEg4DSR+xlkghUal0oCtzsUHLV6LfEHi6bg1tZ4SxgIXyWdXE95J8ZBhQ
RJwQK4NMrq7SOEZfcGVe4VubDHph97DGB9SJL1/y6XPmZZtSIUvMxzZp5aN4dK20
oRJPUdc2ASxOReWHvsYfrsGRRwgMNwBykkM+cpX17GDGr8xfOcJ4ku5fUJmWWsCN
bnIaicN4rKSr4nrWkl1cMl5I9ut7cB8qgBoN1AF2CH3CBvwZ0TinJXSJcoFE2jU2
6AN2vd6yhmB3vpDsFz2PaLW/NL07kjfz8B3Gxb62JGL2v+pBc7V3IDgWQoO1iu2I
2oPHGcGGFCP/TEZpQjYtD7LNox4wGvetIOKw8cMT8c1nKzasArRaB+wByXfUnWZB
KCUWrDUbSh92XTSEkd/osMbvKuLBS0jmBhBwSCbRBqbZ94BcjGsV0GC8BxdJ4RtX
lLgrYOuHKNVx1dKoKK1j/12UY6mrkRQe06VoHf8kSOakCUDYlM2gFaD1FtmAVxKa
G46YIQ0DmU/0qIKWiRpjDp7bzUoOyA0+9462S70sadJbDlSJaSYxFPyLaSqbi3EW
L4GlH9nj1oBtm7BRJ4+24cY8A4wXKoFgGTBAl4jWx66OXD9gLNnq6yGvHKGS7m89
0Wfo/W0jXJmC1xgi7OX4eJWSfVdU0waZyBjuMBzSZmgEj4qnbTFGIwrm4QAAeViZ
5QJ+azdJLQONYNLS4BUrvWYe7eD7KsVoaPCpj0H6f0eAFTPRvRGyLAu470k4BIGc
80hO40Q1zA9KfKj96/MF1wQvd9K1XFASy9XqCPbta9Os2dLG+DkK5sxr9EaL3WrF
t85yebJUTpwuqHP/Xou3zkh9wSjY4itm34aJFVcTa/eIsTG99c3/DFz1UP6aoMgp
rgGl4M090DC9MpFCMEV7Mw7Qt/67V+Zt57aoLiYPlxMxn8YSCNXWBhEUxviv3R7W
r8tWIKgWum0HSByellNpbNHGjpfuYKNfgHF7I9o/Hz3Lq3He6aHse/a3rgYrUren
2WW6+ZE88szpjA8phfRRosQ6vgF69ZYPEv/NolbYPokQ9LhGo6m1DwbFCWPGJJOT
BzgVI0DsPSWMT8xcpNEjm7itmgNa3CwNj0L4+AEV9Y9pemOkSuOSonYLgExH2rji
e4qaz+03pbNMffS1J2cDPYAsnjpZQHRIXwQZRtYgK/8JIdlJ0E9MqF6LuK7wqscY
VR6SNvLnaHvtvzlGjVRgdABgfSWujkFlPErJgB/sTOpsCLUtJvVgGfeIFPC/ZSXV
MPYHs6Pc46UEdoByoQuD0+iPWwhO69r14aSgTb/B+l1fH4v0ugtnJ8gm0oBRioDu
S7p78dkmW2guRCtB84yeU4dnDTCQfcS5fs2elhcuVHT7EZVjljotmBdIKXXvweAG
kynIPFq1/9v0EGCKoW/rS9GUVQ6SKWuKxrBjyipAyviY/NdMuXpTBh9Im/e3iTie
lCzjqmCn+iIgzqVGwA7XO+Mp875CEbfYzHdWPUAKT6dl874ZOvoA8TnnyQAt7/Gl
/9G1PlQnX6k5UKMpmouzMl1rVd5FXUzCcQM+8Kfhu3RMZmI+IcSK4l6FhwCKh/Ey
+7qAozt4/mtKJNFr5HBljuO5Io/r9msuETZnhsn9SFabz3LnNSb3Ds5iOSDX2+NP
Zh5BbdQw582pkni7tkHcti8EItnTpv+Pwvr73KQXy1vsgQueZN5xWh4GM6m/uz7u
eWWrrqKBu60/QwKFIFrRjRGjkCHRbAzUZIrIUzlhzYKfpQSSiC0Q2hHBOKe8DMgj
Jw1h6v1Vpsh37phhCNizJUb/x8+IjdssqSmXLjBELR9LROCh9FdCcXuJ4SAzR/0m
1weHiTrACwgByXvIeGqoKcwnzsp7JrsNAKOf28tHkbHE5EhSQjeEEGx/UAvg/60q
AZW0WMI6xo78T11++LT5idLbdugNDvU8FasNddNHMr6TO+wnAnlBeTkb4VWJ/40w
/trQ6Zk4pBrUFr8rxgCU0h6gk/BhF2V0LhbL718jUzhPHxg/rxmQXh9nHyu+RTdv
CT7Q/YPU86acyIlUngq4Cs1OiMxCuaBoQDTTL+ztv0ZBNsCqCjy6fAUeatop0VPx
SecONRhTa/zpyoSgIz4KJ4hZpWXum87TEQgTvAfT+VGu9jJeSe34LaQnRJFN+Vww
gjGTnEYPlRjy4jMLgVf8fH/LJsuWvQT9V0vOsqIoQfo+KwgC04HXEAk/n4hA/XBl
oeo+QXvFfD94LHi7WDBfwdsi7acwu14lxKxkCWi5uwy04pJf0gUb44FhD8lfNXv7
zcXRCy+GudE7rtubFiP815RyylY/+nMuaRoAYbLhKzS1n4v0fsqlakXLUcqps2sI
HTuk1dWnQsKvmRz4uYnH21zSzSFflhQeSR9XX8gWH5/WMDbydmVX6RAszpbzrG6c
mg0GwdAt7iUf4IMmlivsQtUhroZhkVBKJk82YUu/2qHeIs7G0qqXCI1WItPoStqM
hI0ex+n+T9YqyKOqIZTww4buMLiPRjB4ICTE2QsXnch064OKJ5ViTFyLlmCvZs/y
vRMMPFvWoBcEO8s1UbDR11yNtVhfvFDjrvSLuvggIE/l9PUfaoZAHo+GydA6CuuL
sSraCzo6K7/BEP23rWsb2N28LJGpkNgQp91qOwiX48Wwx1yHjbKi0VPjDohRUBwV
Cu/4baY8NJE29F67KnvVWSIqW9O0XpTcTJGoqPARm2xhoLobSfHEbI4osQE5E6Za
7W9Tz0sY1Mm5uDqpFIZ9nM7N7b5jaWbEttOIdg1aLdoBP2Bb3ooPFkHVLjlRI0b+
o5YdmSgQzdkoAAY9Uz67qivrFUKMZvae97WE2TA8pNPsaxFBuwTVahwImLcKRnkn
Vrw0Mmt0i6pBGUrrFYNvAmJmwcs1YtgaG/1qVnXDYR0sHjX4yCYkbcqy3+LC/ufc
DiE8pcDbV3xAwxYbD4JkFE+4k4U/hpc1RepfiOg0NtgrIrnRfcgzEBaVyWFZY2T8
P0noE8ZKPbdgCOZzJbv5zsyx1myKrvDMDeVmak1ySZ9tnei2cMcHce5GJt6Neest
Tq1n7qoYT7tpNztfCapxr8STYWhHR1o7h2qLJRNxyQbMOfb0fp4iB9sK+Y9zp/ua
VvP2ur1oqbRijUnJdpoSQAkfq9Fqt0prtbvMWswhs723dcNjAgzR2g5AEBDKIrNj
InFKXrnvD7ijRSk6RNUm6I6MUR2vNSSG2Gybk/o4P7MAZn//KPrADGYCtodNnS8V
+BCsmwistPIy28DfGckXANIMAu8phdq1ZL5DtJjz/9coKEOix1zGDpUYqRfShzn4
G3Ixl8QQFA23l8pTjXQEe0cEsTcFiMRVTbKWmzwKknIold+L2i8TxLnPYePFkmpb
E7VKnvr9mMAj/KQtpWrXeLgTs57E2apFGo0pFQaBod69R0Kq/1xgoKoaYJ/Xp7HX
aVZaBJHFq8fZeMm5LXK30daLS/hVnAdhp8LvY4FbsYY6IUdl08uQ0VSKN7nW5cbz
5PSFi/zhUbQGzBihVTdN+imKHXIKcH8NSvCRt9xsoTOctk1InwCpz94XrpjFJwlW
Hzxz3ufZDOmw0NrZyGlqnsgmIXaTEgp7e4AAoQQx1wW+yWjo6yLFq1HvFqgGVc8A
VTW62wbycKxY9lYRj71bzMKrsmE05dbbnIB4jAVVzsbIptlGK0Q+PLGTHLBep1ys
wR0vJIg0lKKZIJttQlKEJiAvxs3dWXenHUs55JYEahbO2T6KuMacIgA/v3My/NV9
ZqBvocZAI+ic2ZV0XGXb7W8+42eDMrUq2SMBvpBvqDsLeSNQYIUiE0R6EycQQrVM
+wNRrymPI3k9le8AXxK4bInclSff+3eCYhPcJHv6ZkdYnqyErPFXbEs3dtIiLoGY
GlNzmSHdK+wE/jefOJETR6X6geML8dIaDsDkPB0uHT+6mHOH3el4FYgBgsA2kE4i
FHHpJCBHMXpuUEseHnm2CGDZKAJhpIrm932c4eZ1oBrmNCjRQKYh9R+t7Py82HRz
XAasbCEk4zwZjdqGhd4uB8lBWnFyCPTDGYoxX3ZrBLlBUE952Ye6SbLli1wxw9fH
JerkEHX8rwr3u/stZwx3yn/ieJi1wJHmRngQMJ0s5UKOpUxCO3k+mscM+2W7P3Th
7+3bgsjijzyGMn386d8skUwBZNgoIhpxuEZFWa/gFndb3Va/zAZOjkNHQ661+/H3
5eBZXbzYgMRPhmahQK9I12NBTRGCSaruJeNjEtAaW8OLtZIMqcmDz9hczV8vwtXj
L3NtafljF6MaXsxSentBhXZRxO92SITo8H/TEp13w0qdXnxRnaHbWg6Z3eDkmgbX
pFyBW5+8ofpO6jlyKzCA2VLfww5EOpQmXGOCYIjNUHEkR9y0whdQUAdEzGtPo2fz
8tKGTbtM5Gv5c9W2UwGLXeF/rZqRGLYSRZMml/Aol0tRB9vPXeQ/o79qKB/0nyM5
AAFKfuxNn+77S7z9+ri9TARN85wR9k7OBocsAuuhnjdXtVSfC2oUqvSgsjIf2o4z
FrExjNXt5k5v27ra7GP1Tf/xC10GMbNCh4Kum+HbNDROi3hLr0Fcmpxs3KWhbGMT
8K0uvOYH4ojYoc3JYcO1WZOCvBubFhLhmbitjvfzggJvG30JEtH0E6Q6TGCG+0z6
A6kmRcB3ARh2XRcnhOkw5S7UhFjM7b6k+2cl+bHb5JK52B1Tj37T933q7UEWGYS1
upNYKj19QiO4se3M5ZDiRZ981EmApFLXzsrM9cAa3wtXFj11C8d9gGs/B8rlWoCS
Hzef4EBkuR/4tUyOcrBocSd0O6GSU4EozzmZPwbV5jgorfwrb2DFpJJP3pPkDjPB
q354FZAMBdsHdmvWYHsg8Tce97ljVLNnAyW77bsE8TfVLEAA6FDyGf14SQDAfhj3
ZzNbMImeHVJRuqa5Cj5GzGO89spI3cgAxhbtWlJr8A1tGVtQC3sDV7zmexgEUaXc
UU1O/RNjYCmPMsl8bMeaIYb+HenWFiPF/x65Xj84KGe/nH6SMlE4LZNMh2Z9i6I9
B98irkq8pbK7A8Pxg8oEtUf1Thjh6t+Ik0/enbv7GnBoOqnsKGN3l1z/p77xlH51
1jhCWBIjRnKbXsFd9nWys3ctBciK5n5SR4BLHzfLZG+5fOX9N6pAeGmxMrkG68yX
UzFYHyaRtrcDprVeugVHSuvxsBLOnS4w4io3E1zzf85nE3ZV5ZGWEH0l2nCflT37
TDmGj7pQy2Kn/Xi9yIBi9OIQnqBMBQoItS6RVZgiSX4M9QOxG7QmL8+IzCPhfKjp
cVQ3oKONCEnOsPJOLw4RDq4pk2iH+wvqufsID7WmpulGMQT25QS+CCLvzqqSuSUn
vChw3FizZxnR5lW5j0wuGkkKeC+Anzb6Nmc8hS5YVPVONoV0iHYXmXnWvQmdR56+
GUAS/9myYpI6/UR/dKdPthJdxD0Hz3q1FM2DoXBqnnMupy3qlzBbE2VTNKwmvWxZ
4pbaC40DgMLJg2oVZl5vI9S+ou55SPI2S4Jq4UeU9Zf70CQrD1HyXI90R3hPY4Wc
7lpRHQsux9Jt82m+w/L17KgFZZ4/0ErfUfi10rFWxgFXZq/C5dvDA9TdmEHaRayH
5i9lQzj4OVoJQ6UtpmgAnSfZqOq9/IpJFKIs8x7bpzrBvaANmKsAwHzDTq4OvhtX
qorWkiTPUSvzm4x6qttkYfGYzy+tJwwlOicUFg2Thp2Kpscx/ekvDnibe70uSVuk
VRmUuHOl0itxmOm02dSesRhiOMj4FcrREHqJP82N09wOZW1DX+NCvdMcQ2Ay7o/a
UiBgXIdO12kxtGZtedvM+XCVPbjd288QKbcyVy5R8sfnmxZ90L5hiY6HkVJrWY8p
J4hMaoHE+W2GYDhpRprbcW3cjVr53jgkscWsF28hWAoIydWYFL8iKyVwpYB5Ayph
JCaf2Wegvme0H0cpmFrmXVN5hBhAkNAb84amE72HQxSTL9dPAFaEiRqFXaawgTCg
zmSwOF4t/7cNYiIFnxeTZOX4zEhYyNwIcLClNRRXHMoyi9gmHWAlq6B7AjCh6a9N
BYz1XLINMtbs2/n+mTbkVV4sVIAiot3Wrj3V1xu+TqTuIGQo3pknAHyDVv3caWKr
/DeRyOkEVwCccMETHJ468f8P3Sakem55yNAP+scmx1uRvM8ETEL/tY0G0vdmqTuq
zRojvK+MEop1C3d5vUsvqGGYClJWxNxXePXWIbt0Y3S8myD4IXPpBKtUSr4yRPE4
RlwUGo1UPC9TSunsv0/oYkVa/2UT2cByfWr5Qm8ZGJU1imKcuLLlIR98P2Vl9nky
X1yzZGSPU5R7TZHOkWYBx6kkwad1E5zVHwIfV6dd+vydnpm7N7U76/ZWVwfFwtNJ
/jURNLuV3No7BZscnf43eLA+S+CPm6EfOSbBTQucOOq3kR+E0BZHrEE2LmQkAYi5
PRD+hgQnpijqQ4AZBTeGtwuSz2IC17pxmr0hH1p833ky7NH42AU3BG3vQeMRe+fq
Jb94/QcUfnQoa+uQbb7/88xS7aJo4pCox+OUGNYusgOKOa3JqTez0bB3pgR78dkQ
klTwQwIari2eeNXczI6nS553km7UYtIXNXmxsJ1wwwRCtfQID6Bqvao3Pap/Jyk7
3sffea6/iemAw+jVX1fp5OlhxM8Y2IAt7R8ilB6nY5IdDPrboBm/clUw0vkNI7Lk
ZQePT6mGZDTl8P9nuTdcmmNYE8swMBUBvAhVhnw7cXbSYVGZeAVGNiOblF7o8Gj3
+GuCPxw06I4GhwiGkqlAezkAL5t8Ro8AG3RSjjDey/HdJD5pIF0IOplG0XwapC2E
m59ESL5HBx13Y4kpyeGLkGkv/F28T2UnPAV+oZJy7O5wxqlbs6OazrjlOsh1AIqI
50jKATEah/IJVu23CHdNk7p4basQBweDu4Bz+XOcECGDqmAsup6T1xjkHmuRjbEW
/mGtjXR4eGblClb6AkxlVP7/8sRaBb2AA0pPtNxdNZw0glI33vnJ7q9g5pjUlunt
pL9jQ3N2ZyXsNbbCDZoFgP0RIGySWaapLh8rERh5d79GhpJ0cu9ifbgWoXMG3Z1S
JxzRKpsCdQUaH4Xi3bk1q7MY0ZMCkJIIdxJpl+j3kWOxuNOVjKrFRfkMSLLzL8J0
sa0aigIo6ZMplhIaPzpza2mwbSqOhqddju2h2Lb5xeFsTaQinLK8KxgpKGrehNjX
z4wB7m+MvJcX+tStE8Io8eIqnXmeps0STF/IftfBfoxlpPwLojjavjDxk7++zIG/
bWbHX+5yRwWDyrpGXOW5l499Ynnxh73x4fwaGDbafUkL3JS4x0TL0edpe7c5ccaI
pOd0LaYhTNHKfN7GYZgzXfAXvNDrq/V//b1Mv3J3qdZOBjfpokteC3LWFbIlLDAC
UdHNN+tOXgbuLWCgnryJfOCk5WpQDJ4M8jqD4z2xVi6bEhnO7SlkD9NeujPF1Yx2
ADCVGEEI+34aqsyWa190n3Quwan7urjUNL1r6cKQHeCOOa5oOKzV31ssbVgRODRB
GiUFKY4hmK6VTR5f03jtD/707V8TAG5CtZlhgK8A/2twPcCVqIvDt229Uof7A19m
KpubpI4OjzzMts9nDtDl0nmvKl5GeeWs6jfJB6D8QlY3uI3Nz0fPr6g3i04Ofnjp
xtpE9u3ca9QlRoOaeyHhTMKnlbctsvrOL24prOJ4BCanMG5WjCCQAGUvVDZg1zw3
tu+NOZxPDtrVc61AHNQwE7vxoLx3YziT1r5I3VEB40m7xrW1edz4uGBlLu4G9IJ4
CyiODFC07yD7UVYXD+k32YoWen131GOwhbZgxSNpJL49NxAZsy9ERfaCoIgzDRu8
WBpIqe22CeHQPnHDTtywbxAtaJe4AhbNWJLVu8ltCZFI9A1iCadZyOHk0T3sje74
nExUe4fMc8+/d7UsNSSyMOLQuUSj0PSnDk5UjCuFLXzBKaGxrj+rRUlDoU+1/Dls
g4AiOs/glcRBFJqVv9Sno4LHi2mJChfE7Qq8aJgnrlxW3wlFCeX1jBfgASk/+BXS
Af7U/TTwZRtmb88hD7En5EeV9pkWFBXKiduLOszLTv8d5SEZgA4ZdfD7cXUVzuFI
ggf59h32HLR3xk8lW+YH5LIoLDiMtjYCo/VcLpNnhi/dOaWEMP7waDXoCPqDxQsn
61V7sWKgwiB2zGH6C0oVHYg4qp/T4zci5h/Fn/Pz4EVNBRqVaPxLnvlDPjfRpv6i
RRaLvM3RBZ+nn79HGIw0ZXCjv/9cvU/jcETd+TTyFhMxi3OGx4tqCNUJUoXawOVb
Fl17T2K21LG6dexTeGvroaoE0kx9YPICMjKzCm2uHSKZtGoSVZM6UNmlGrvMbXZH
qbnYgZJGPFcBkaUuxFxM/6A4L1bwZXeckWH7a6Qic57mCrnUi/F+dIZZCCfD0Ax4
TuH/skwwzno4OBCprQrLrTdx7VFy/oQF6fc9fEhqxU7PfFZjS3xajhxtnGlqI135
IH8i59fo30X2qTCzOefmEJt4kVsplKoU2SwDodVDB0QR7WK+76nt1s7Xty9pm9hX
F/LFsVDxbGY6Ih3CzQcPnQb6uwLoq9OEb7IsASSPlhJgM8aNIBLzxB77SdluSRcf
iKbH2jBFKo3nIImtr3oEcGlMQ83osO9Ifm4HTVuGgC5r0mXqZM7aIcbeN6vZymNQ
vjt4BdyrIGKFzSqgvbPTWABbXdhP73GtuRpARETHsetsFLEthxpN4tuJYZsPvh6L
5xTti13UaUaLFPRcT5og2UtpuwjOn+08b1w2BZWOqf5IsvMHJh6KPQtBjHT9awFN
tTiUlnD6PSAXJ9Qh0F3O+YhCnulI9e51aib8QNzn4awudXFOYd1g5FLhY5hyiCYi
cvQEoarAu1iEHJfG8L0K2EBVpNSEA8EFiIXnhNw5tbS2xUs9T3KbooGxkj/pnxP7
6WF+4yFdK/paNIAqBUnMbCpDLcLgtQo3cz1g2nLzp/U5pERveUGYMHcyh/s7yTOa
D83NJp9+NOGuG13H126uqgBtIT5c383Kbs3b+HsAFah2W+nhtW6H6EbIv6x80ZBZ
OlbHn474sd1YuxM4ofpu9O0ny7eoY9c+pxr5HTwFZ8R4l0Nhu6upjI6UIFRZp52R
Xz6fXU3AgVhypjXoQAV//Wwwb2KiPUZnm+R5HwzRU3XrgXmZ2GdSrv+635EPLbhw
UPiciiC2RXf+x7pS+ISIadVxnAZLwC/LRrIQ1NdYdxa6qHXbGJegDBmufYbcKzK9
NVdwzLIovsa1GX3GDcNvBC9fmFdSGoMsDWjFpOI1s/OCe8pBVHuazLsVKjwghePP
mvhH1pNQTyFqEd5yQew5O4nWP6+Lm2lRtPUCWge3VxSOavF1glHzY0i8GXS5+/V3
kKMr/mzKi5apUiJTht1N8ZjENFZ00ca3U1J+iDSJqm5WQKYVnPMZ5/gvm4QHr08q
gJhDm9cbb9PllrM4QO7tLSKr4PrtgLa4zfC6zkegnfuyLz867hv6qT4Rui0uv7EO
x0NPgPFyn02oIGueQbK82/TJNalkmGy6SYyjSrY0wbRoM27DgYwe2BctN/X4nA3W
ZkzzYd9YOzoOdQHAvDoVMmYahVEHXquivA5B7Q49toVZPM0z3337nzIOGstzasvb
DuVlUo0eMlbyEptsJuwc7XvsTU2+3IQPsdebJOADguGAtrizz1gTwaZDjCSv+i6M
R8/++Di3VZ8tnpJHr1JIgFwXyf4vnitAmhTD/iH1+HqYOec6cz6WAgPwdh/D/n7p
+804GiAlYJ9aY/CkW1k/DW76Wpb575ZMgvUlhzCh0YK5vvrRUmVFxPiwB41N7+3c
OhMNO9b3JaGbo/U0SSZN9xTyDI6fJYPPjYWWMWPkq5y7RH2+dZP2R/aocOWDmsEy
wT6kQBvszEI9g1ZEEDuglnATQPthvjomcVivjBN6/ffACTg+1iTVo6Gp3I1V3Pd1
kAWHLzs6Bo2FskseOPoIkz2wApDLS+nQolh8lvQ8SaHQj53UXVt94umHXpzVGz5e
whSmeo/FkRPK8NAoXtlGj7sBwklXzR3UsDUK6/JXW4KoEiVmc2opyH4IlPVrZPCg
duLrBXS/BUOIJ1hoh7+wwSZS4mN9XiucOq9W6qdgq0aZCyxmxaiox/S0UYprss4B
dPSI3A4r0n0p/39AJbLs0zH00qTGsxQzaSy/L6U1OHu2hZQnAxYlhyyfiQ8GGwG5
D5HYQ0BxG5VOxCGH8Pcw84xBKaE4ptdUnlfEDuPCXyzfn+di5h0X26EU6PZH9fpE
MzinUUIZsMHINGlqALP+ijWMEkPWY9AV4bEHT8sYjkN+nNho2B7x6M2F3BgWlBph
tE/hpH+kuYmH+nwX4t/Q1SXgHB+s/I5ikTKu9ciGdq0AtKVLcVdBuajIXA/it9cO
sgUq9bhTXAvmNoeEZufBqNG9SWZqbQCreQ/DYiwwYaeEZkQQP3w2N/JlksGs7Rlj
kH8yaYZLsVZ1VDYoyQMx69loDBqInqqY+1mMNPg3wnUIQ+RRJbGlB9ZqKgiyOhWk
TmpQQUZKpgk/gQMkxtcYwLC/sGAZSbnceW7Lhvom3APlmJg0SgAa95RxyGge0B2d
AW5bupP1/DZCMQ2zRGaJFjaU4j67+2itz11mqQC3wWnLugUW5/b8Y+MUdl+QY6Np
n8kHQm7uWKDHwxS1gi5e0FL6btoRZeC+8mo1TpneLt4F1LKHmBSbFDEG5ITongFM
gCIfrc8vfxub1kEwQoDnJB41hnV7uIxosrflArJFpT6jt9Au26UFQ/5I8acD3FIb
glyoIAzAp1H+p5RjrccVjjuydhxvInJK31Q3QTqoQZxZrSi0qMtGvgbj7ffXha5w
lK2Rx8nkQVXM6joIvyAujh3Vb1SmGyKjtM+S6kM3YDHQ5nZTu/CYe5LRUiwkaHkW
AmSzykuWTwJWJ3NlkplSPpjrMZIJSx4e+DlxqTzAEDLCWHPK7zRRp//coB8HhnNg
j6u/cULRsks1E7+rz/XGYOrYft6FCd9/klvrXPC/apOvm5EADUeUOu+TljiwwCWE
qtImTvnzu5l8cRBVAHO7Kn5yFGIPxAV2T702YIIxuKwo2I+tyKtY29OT3LqQSz/6
V44VNLvNdH4U5QT6CcYiNO1Jeh3ML2ytoqXbJwrAw+sjWZ6jv2fr3QyN4bIIBE0I
X+tOgMyDIQbARiw66C1666wGObXKt7pWArpQuH9dYvLKkMj+GKojFD+Dt6R2kn2w
QU7KakFo7nKPFtJv0d0kClRyFAzOr6oUYlwM40hoZ1L7TnqL6+90rtLioJA3aYnK
hKAocQgdoK5Rg2f5CSZABuQNaOdZklU+rrh7lIDRaswkIAj1apjHrgBrUbNlTXow
NtU/RlIDK7NQ0RrtRNAHhMMqULy2j5cmfRRxHx1duL3uJkYkgyWVGcTpElbkYcCy
eonWPIkk48dkME2m+hDh0dQisuLBKqZXr0y0SxiEbnKjmwZa3/U5C9a1rLVNzwOL
S93s41jtfAs3kjs3VegoaW1BJGzpneQZFwlAEvVf3K6e49tU/nzaGN/R+xDwARee
HSr1uIZmY84u3YjxZaqFOgG8hut6XJjXUmaGkubCpjHA4wF+lxmRyuGJNc+NUcS/
pK/ZYw4vMBxoHei5gma06GqvQfTjbWdOQ6MPMCD5ZOgOwLR9v1bdG1sy+aELjUvX
YQmPNWNgfatz98RrAjlF5od4Vvp0F+InKPsfvAIFynoL+It10mJTLOh5vDq8M2rj
dP8xKfSihimiUt76MAzMsq5AIIz5QB+1+xrqIdqZwJGGX6nX+mi5TMKPEPzoB2ps
4q3lrfAUU5iWWiubSWQplrt5o0ecfdGGEF0d2IcRi86w7/oZAP69uTaBOyD3YoGa
BONW7QxBglCp7P5EXQRzUW5H+jCJs4fFJ+3CpgdYa767DKNgrFOJ/BSg6z519dJN
/HNbtKSze6ThDX78SsgpYQJ4MIfqVkG59lEowl8YdDEQaHSL7cD0vM8ONOevoZKX
UH41EAGum/APjnZfH/5Drb31R8vPB4V0wPl96cXzZkvez9MXdMYWO+cYlLjedYRV
/O0Lxc0qnyjbHwHptuX0okWOJ8200oE6COG7v9FIgn7Jf1TQOOiHfhDYiW4NTOMv
+tqUNBuHkSqgmsDFyq00y8L+sKGpW9WNeoLQ3k/DXKvdQNEsca+hXpG9zXPpOjf9
aV4KG5P3C1leu0l8xmVQ1BXQHflscDVB5tb8qOtbkdHbgY7Ct6VZuils0Yec9ck2
NPImaYrDWxNp7cmYIyb69lFaAMiCE5LgWhTbT9yVgzy3X/pbf4oBfHkBi7AvvEvX
kTg79BnjxXat8lUJmJH11wsbkDg4G8J9kyfRxEXUILfAApP409NmSTVh7Y9hYH5A
t5fxCIwRY72dFa18ZjEnODbn4lEKkbj9hJOWk7QQPmMbaFOqvVD5orDcpAEV3182
QimjoBzFDQja0tHAj03VM+VsG3399FjX7R3Oq+OjxFKvXy4uetzOT7YADCKYiLpE
MG1NujaAAC28z+wm45w1WVH7RpaMCsICL+s38WNA5aWvjlcKj6TUeiXMJFbpunm+
mZZVxUCaxnFW66WzL3u9Nc8cu6+8zlaHIBfcR5fvP6fqdLa8GjIGlo6j7FbjmEff
9ORzX1hqAmhyW2kxrB3SZVo04KsGEdJ71XIPWNP5JLRyOa91GOgczPc6ylR6V0Bq
FxX1CeFte/8gpaFBodV7XWfyrLe+y5N35zOfJtYYWBgQpLlSHCFlMsxIGUjd1Wsd
5N1v0Ez/3iKmLBGB/ZSEsjZ8TlYrNMsnTdCxmVAuGR6+sNrFMnSNmTbelCgpGvhU
qX0epVoCaOuE2QRKitI4PqAL0w4dx70tvOt9T9e8VUyjp/cwL5XIeyefl/eqw23t
07++nVhcJZNWFyQEkwIIWDy2mRR9B22E6n1LCYqfHwOpWP1fycqitKveXitxPDH1
YXHcFhQOp1NoG2KNVEmK5R9lZovVFWwYhm5ENAbk8FS9oUkDwta5gpsHeNErIEEt
FxSCF9f60GuKz1z/yzwdAgx4qPxd3hDjiThEFtpVEKkFRiLwgX+WIL1pJdPvUO2c
J7+I2zHp59Xr4TzV2pycCKg5RHfc13Xz0miNQ7DqJ11paeFSOE2VisEw+WT7ittt
gvaJMN+IEEof4ws7bATQc6FRgH2W/8vmGmghMn77DYGsVD6UgDOi/HvyNg5G2oxd
l9wlu2uvEWnMTMY5CkJEjdDN38Ef0pau0bTtArUCIZgx4I9T2FmcGbLgT+FFo3WA
fRNf4dt8kYMiuuazushBgcyildHMdejlAJQmGHr2uyUTn5daowSmUYEpQEsxcsQt
AHUIcvUzRrW8YkLJsaar4LC5jLzGQJmB4gwe0nDzHoaaoK0DX7sRHKQ/6dMXW2C6
uOdINMHjtjvrf5/O7UuvqqeO4irC5ACG+UPeB4cLhoxw7oWZA26pDBco6PG6NoeX
5ygJyE/65/loV8UNYZX/Ang7V+YKFqMN/1ez+lx12E6+KuTnePrvXyLbk1icetGa
SS7sEIUN3CWlQe/d3Ugwvtq9nUWZEwlHoNOO5pfwdByK5a1bInItgv2drZjG01Ti
UZdGynmp/XAAGgg28ndAswkxGfVW1gOVqyDF16Aa4AfpoPMHM+6JVpy7XvwVUH08
fdCAcVnql3b2VUPf9Hxu17yJoHcKZkal7NNB2MeFGSg25bzvi1x3GYE0u4ULrUsY
wGy5HXSLkZzk382Sme2PyukccqUr0DsMxhE2qKZsiLM1D1pa0y5klGChIsMIRiyy
83/0UnMW0Vu5KTluaIrsadRbq5pC6AZbLyN0zHwupQmQT1ydGpiFpFO1Y7JhS8nT
8oU8nQlohh2Z1+qp8LGEd3iTMBZMERL5nrzSELrjaw4Fowny00CBvp4viCVN/IN2
/A+StQ4ADzNlR6h13CGGKBDTC9hm/h4ioJ5og6qZfA8Ji+chHzHjUR9ADWSVbUPP
G9mPi4zw8pmnE72ebDJLYFdWHb4hQJrT6/mS+QbYvOThIoYlMZHgs3OUZFCkCjcV
OSmKbHF5cs58I+7V5uhdXjeB3QyBoM/iaFOscbIauhqEuKTJP9T7bYoyXnBvoAKW
AGobLnBo5efZ32GnCumcR6Lmc6FT8vKeqEZTuw3osNsqnpgjbY/KMnsFbSxUsX0a
FmsHBm5eBY8825SmfVoB9IVjp+SWlcapiSJkBSFbbUboQ5WP1DUBRHun9kWDe+y/
dzGrnnsF9Gr/lK9/kSNjYFgqt4Qo1/i6dz6AJNCgr/WCi2FntSojBBM0IqJYMTjR
wdTLs6/4bjmXnNQOJ4nitJKC1gZ/L0442UxPgQ/RV9SRvRsy61+rdoWT7wgIVF5K
AdbrrICgrQK1wktOYjpKwGAT9TjNvceZKc0GcAF6+wV2f4s117+vKO75DyawtO5H
Je/JeJzAI1RazrniJPdsMl/MZIBGV3xXZMiHTQqb5oqb9caL/IS1rtCLYj3SgkmF
UwFmN2Q/hQACGmQQ15qFTMZamCUf0oj0QF3IME5U2R2SPbOq91C1BIhg7nhRulWZ
NO/qJhlk9ae/E3h/8VcfQAHeZW5gY/bLVBiDkmUW0Swbfmpe9KAKoLZtP5fbnZvF
58uqXl+3nSrSrOSzyyUt+7D1Knpj2j+46m3X15tqxxNihqccbMSMeS44FWrqfdJ4
4vZqkppfVAubzng7JhTt1dUJE69DFugd3mp/r1NAjVB5fOtFaU3PyZoutwrp/5ln
jz7O50v8yi5cvAfLWTLGnRKdFW6v9uEiOYrIELuysSnq5PY2BQ5JPx6cJrvRkIgO
i0sE/jN7GFazlgiGyn6kwLAOyEKObN4lGUboBhWzmE3w3qmPFakzRTucUFb0r6V9
Llk1LLiJlsdiMjEMQur90Yazm0bmdnOrFoBaW5ZjaMfu/TcdEQz7Kz+VNexhomdD
Q8DBAaQYWOTo0/t0L7tDD4ED5BexvpKs252TDu7uMqX5FEzGyEgZRhDyR1HJ78TX
Gl6cqGqIiqjvH0wiGrZkCGmY3ZG3/qV2X6PRyaAJyYgR4/Q6uLWTzG/awHAWixYT
qxNIZCZZo10AJ3WjLnOTbM0vUSDFcGybwxbTFvR+QJQxl4yDmV0saey03KvAfRbO
/Tq1JNLUc/2h8G+xvMFkE8UR91++OU6EVqk2Z/XKWe/zfAQ3LPCjHfpch5r3MvSu
z0yVaH0tLq0wJY8LZYMmOq7Wp62vhkdLT9gKHTWjsc2qt08HMP0xfEgj4mkvPNfQ
f/aXEt4KdIxxRTKZUHhxvURE+H3x9XLfAHkYyv0l3ESt47eAbUtNdCuII+5CbZCQ
rbTrka/4bTHHzGlf3WOPDgVbb5iLk/eimS82VZGBIEFhF5Cgso6vTcNB+w6GhUEi
m6O32MjuSwExUNCaXy04/pIQP5YI8ekjJ7341UpoKTrQnVuhJM8o+WknOhi6H/4Z
iUmsLZ9YkHH/8HhceYL4B9yPmQ3v8EiiQWoAAp8JpLpz6p/RisMCSIasnKe5V+FI
y7F3Zzao4DFVkgwjFoimEZU5Pjnpm0E63Zyii2DBcjfzRQmlWYRXNLoZFanfuMJb
NvCH6Qtzut3GMQfRTpP4ifLH9kurzwaR7u2IZTAD+HkVw3UcIjo1utEDcqArIBTo
9lo4SfBX04pnoRGpu+9HeQKb/RNWO5gcgccv51cuIG8Wi2Oj6/DnywYP3RAwMhZH
xzM35lm03wySLwUmqMAKmIFmmb4sDe7JDvBD08hSyjjydWzLN3ID2rT0rDqukTJ0
sZTufb6KGPHnO3pTv/Fem3PbdnqGZ5XSlyykq3bYZPG2t3ClskMEg6Do7xQJCBzq
EpmAymcwJgLmMz32wqHmmyItG2X512ugQIzX4vKn/bc+bCN5zOW6RFMHBgQMdpi5
auCO5uV3SFDUAYO8mLac+YssgGVUcS7hwdtMtHA8Je3tyxR8i02gBymq5CU9dS6E
7eMkxARPkRQtUPNQg7P9yLZSKAqz4zYMupdIb/qHnWb9ffSAwYIJzipE06781n5S
sKgHjRLLHj/PoZ8qntPqP4VpOg2YqZ6vf3y9D5aA0gYbYZlhPiOXJl0ty8ixwlh8
er8ZG85UXW7bBvNba8Q3L347M+0/I9fAi6x7N39dDlXQUJqD8O1nu9gegTPws7dw
0ptNFcS7fGeCA93W2EQKnBxC3KjgsRNRXjcC9BxUw1RK61V/aJqB2JZyIEIFUi/V
LiRf+9SYeYlBs8LIURKwgL7cVuOf1miFaO18Nct81ZAHwFGxZ6JSRo7kXWAAYu/P
4UQErFTHD09enSu5gcsqLFz4VL8kKVs+MRObaoc5NTIFkUjAhkcn/ydESxUPhUUB
3Ce0LnGfA4olny4qawqnnLlipFO4zT3cM5UkIc5ZmLKWaxqw9XcPKAi73JbUIiyg
Nk8OaF5QWHhLKS0dWSD+sHjGeXRieXw2c0c8DggFbLldLdFFADq38LZF/u9ASPfm
Gxa3RQq2KjNWa95WbPLzD7fSdt8CjcuB2cBRdoXyIgOx+YZ1zOpuEzdyH+Ge/3oJ
xmxp1eg32QorQ3Bw/iWVZWjtr6ogVhU/uV9FK8Wnd86EijA/R/uBMO8uDSLQsM2d
dnjV52EgOlFWwTcoYlR8GdRgYyw5hyqeie3+s4Tk3q46dL5kRFsdfPFidnBrtZK5
4TvcDCu2wqO7Xa2hncvqM8efKhMGNlmw+7cN28Qc6xNAaAlf7zxlL/XwQxAIbOw5
IjC2/CST+/UW0LrLmCHEX7B4ElfV+J3+GYnKMdSfYHfNlFoKXrILHQxB7o/3UNHa
NzdBC17l26ShQJz/hLiEwAgpZ+4H/DR21uoXFZLsSWUaiH+yEgwswjU5cDNmQVqp
lFqhC1ujSHH/dO1Ncu1b1c0wZZb7J2BCGaf3uWi+X459gSmncCrSp+5HlJuuGVQE
EPs0joprslK0cPaECRnxeHsMeH+8OvzjNYBEhgAJxJnaH3TdMnKJWAMvKTDxpJAS
x/1FKJMq0diFaTZpx/wbuv7Y9sn7YLrkHLCt9/f9yvk2oUqZmuQ4wu66PE8Bj+ay
TrwC7PG1uddFdMD1XpcdSdGHEQrw9NwrLlScNwXnlxOjZJnByd+tUVQrc2SfPHId
I19m/isyr65YMHUfWFxzMh08dGl17I2DD3DTBEOs97u6Has++v1Jaeq8vGhWIGqd
OgVYGNub6dcqUZVohfsqLyArslizefWrfIBk2649FlzSoUYytoUjP2EFExEcnF/4
6E8HA9ZE5oj7gzCfg0veMihm3k/FVahg1PwvfzF+SICeSUNN948NQC2M0gCII3F6
VZNb8msLL0IdxUUQQVONoQpTJLdq1o61vzSXGl0Q3I8dolw4QDJ/fmT7TKvKb9qQ
ZLxM8IqcV5GkMYO8M+wu0zdLMmQtPYx7X6L/hP/FFCXL/GR1N0KNw+hHAJNCh4cN
P5q4NMSbylLlIfPkvIPevtRTEGwE+qJymv/BXH5bj5Z8RmSZyIkg3mG6MpWHLdxh
1hrf7ilx1+47qjICyqWEIIR+XHJfycwSUn0RrLnORAvSde5Tr8J5O+P4nFieO7Dx
mMaJzsRKFjhWcVKLmgadtPek8bAZuOCBwNK36DkN56FCkTn7+Q47EcCPwbSKhXPw
z8+xc1fRbZE/2LiYK9v8SmWQmJtXF56fxI4K6Z9KDBAOIymY+hHBp0WUb37xUTKE
/vWIdoXz8VvpZoi6h73tjY+MxD+MzVWrw90l/Z1OfLsRH3lDQwa7il4UplSQlraD
+HtYLEXClE9eSgeJK3LBLBHhQAay+4GfMBZ9wQ1b2Tu63oqy8k9l3jnBvPZPUA/r
+ZDayqn8lQNf9GQEOtbFt7quLikDdFiEvNt0cj6GnMico04phVpihdRf4OGuF9V6
aXOw1NqT5PtJyMAtvZqMCIbKuj74J/LT97AtpEh/DSMC1QnE42GG4tRK46vQ0Q+9
/+VN3dAn9+hCZE1T3nbEfivweqx2lo13bSsGLFZwa9skGuZgg7cn4L7x8k33oQKV
zDAlPfiTyNvfskdzoyfa7yf/cZTURquaaNBg9byj/3A3lMAVGlTOi23UAgBnbYuC
j1RsMPnLaXx9fO2lzrHs1cUvC0jUq57K87t+3LJaH2h5S1zkmze1eWTSv3Hm8Uoq
RvC1jJW/ecmlcQjgcpp+qidIZhliq9E2/ei3tXjYfT+fM34Ps8I7/1SBp/w+TQfC
IdFUGHUsnBahwhiOGUfBL36rLCU9xSZ7nzO5sL+EkprbiQWr38TOQ6GU8AahbbJW
lwnCIBS2ItulMcRg4TmLgPG4tu6Rc668lwAIWsqPXFR7P5N+kKnFAs+2rkua09HO
239XGnA7m1CwX7MqloQm7aVHTFUU2AdvsvoAAlGHdIGmW5U3g3/3No8hvdl81GGn
ITAM5WeUKUX7T/UPyZigp8fu/aBu6TZLoYkSUk7MHa4EgpA5eabRMDea92BjLEjf
1QQsIjLJGzOPO/1MRp5rAHrD8QoePc0kkD/KWYMDI5qNjQRVhw/PHFTOFg8QYIjp
IJNCPbuF0ZxC55lr5VW7LaXY/RX8U+jcaZp8cJLQx16ptNPd0m74ksjYJIYfiR+s
X74SblDC7vrRLexEPAnkmWDYl2PDD6W9pklbW1bbHXsm2dC9nhrmTPFOe9oGSMhp
CnePlZxbDdw7+1Y5jEWttgMBPxUX9SOj27xmIF6qcwdeTlFO81+LotIXkBnm4b+l
rEytTiKJFw/Zv5ODvVwMx6OGMUcL3jSVkchOS7/i0oeBMAxA3Fqh8dWsOQxBRMzY
GUJ9jIDXfZh67lURWQSTAb963pJT8o7KBGK+eV2YTWM8+avyfG+u/VkVZ4HQNaR/
pGlZ9tfjDzYnAEKyRkD3D4P+dozPlJFG505SbzKjNwPObQxAquN89q4WwY8otDVx
sWL2hAzl4peyZbcTztjx2l0duRuTHVf0BGHdjfFO3lbNM9mJMAIaWi7u/IOiW18u
VYO2VKSijABxFW4R61SYbprAM6ZkW0LcJPRMrZ/wydTyftlzG2s7Lljxi74SI7c7
dW4Zpg2RH/Wp+NvNEL+tZdZnZ1DbPQJPqWHnSDpcR48MUKbNpRWzCxH+VCffFnFv
spbo83p7mSs+nVeqDlPpMVu1rPE5TtQSiFeVp4GP+NS+ItuO1kI/6m4jp0lpOnV8
IBTr22R1q3LETxfZf7kzfWFDwD4frIVPs4J5ywu8tAAwl3G78XjxdXXuS8NYzWBX
anBrDjybv6nzmj9A8D+8I4Bs1m+qRLgfMUmutcwuoQ6NUXrhWSrgakGHA4no/N5N
kcoTFhrrZqryo5+Mj7XXFLxT0HFV5byhwX2TZ12zkuIBKIOmdHqW2E1lI07Vhma2
qduAm8jZB0UYJ2IkOGqfCZLPLtGcsa7XB3owKS8kXlzhygh1tf7AK9oxvjpuzlOh
ChjJ/8WlCCbeaIY+0Fu2Hd+Y5D5xCd/TA+gbwX9cBRBarZKSFQ7tqsAhnRBfak1g
uKTMIUC6c7skG7IIz803nDRXO9gOgq7Q8AdAR6vMd8Y9WhEHa6Y7ux5M8ZNF/UC3
B5mo8xz5ftF8Yga06rdPp5OBV2lp5v/h+51wFZetQX1+bI5sjLhYZESthR3EqxFJ
2TN0yX2Pyy8xTYcw7ajXlY6b+xeXcq9TAmg+H3Lc+8KHfwKBT4GOZEr9bfIaiyz8
vsise7QYuba9mGtpbnSfZDjjTWcFafZBCdXIV09MMD/WqjThBcA5H+0Fg9qmsDzN
PQor5S41uxowXAswjUVhmM/1RCJrZb8QCFhC/aZPoL/W0Y2TzPvlIdXiWOVqoSAd
+zhghCwk/3OzfY9dDfxf/oVkMeXjo8YbKJUXOCQJQ4/Ei2j/nfjTw2TzMx2Uz2bY
JQFbofh9ZX5cCQYahGA7HW0yEOs4b4IJVTpbqzHpGlq/u/r+A6TeItffChIq+JEE
fXEuWF+jbvfzUOmbYTxhx7BkMrcOZGtPa5+BP3Ya477T9ZFA2koghABAKn/EuITX
VO2C2pNtmnZHl2q4Qtc/fvqgmoNHJl9vEbsmIc6NhtqcZp+XSKywLjcF1J0YUssd
Dm3teclvtCm8LSH13q/OIBqqZgsGDG9w9VmEEo7MhXjwCQmzVR7K5AMVEsa5oTX6
9NyJIahBJJQtbnaz3qmiG7Lq34bUgPdH9os73GY74ZpWGGwrgnHt+5VattNxGWSz
V0EE32cmVBRFMTREVoBMwotCgat0nKC6cIpohYxvdK9FoMsUcqw/uxq/0tjIg3C1
GKN+JZfqcdddS06Av/ApRS+wYtQLUQiOrNDq0m9DqtU0HybXacocKlhyosSaAEFd
05Kd7n2zw2I4o86HMvQwYEh3Mq/Zw6odD/cJ/AdEh+tNXkoR2oH7L/NWx5cZE8ck
r3jf6Htcef5oqiegQjlxpxrrLzqFA/+7I7ZOf1qa+WzSJ7DLyZrqfOygpP13ABI/
GPEZ2deb11v9r5kkE2Wov85+ILN+SBaE2jKQN70aJyT2TKJTlkR9w72P+aZUqJNe
d+iIWXKWU02kFkLvvQNVx3/uDlpGJfOFmSpOviXUdz81aYSD4PquNBq2fnEftywY
P4GKqRQh0SBzgRb5dIU2/QIIvNKtyzdgVoMQhjCCAZjZxknNeFZI6T61Et18BX8k
6kGPwqYKBtzuyP7pQDk7QuFbXI+LMT8swLr2S++XKNLvdayn7KXVFSCZFvfMpT7Z
MErYX/MN+g52sU4X+2ixztH/eyS5PhoOmFl/WMOlngJP5QikUdA/4kKIKv14no8A
Kj8LvdK7ZuetZ1ujk9Y+hUD+3khyZ5UKWHW2GIn2A2+uRwjoYdEZwEmxqF617KpE
KY785JCxsjJrKmCPA9DMvfk2kZMGDcaHFi6Zsg3fKYCwT7dh5ttPxlywgu2h/B2s
tvqo8Nuu31/8vcHa2JowyKg4OSsMMohxEm7SNZffSmnRSMqx5O9oocHwiLYkkSeS
l27LpWyWDF4EiseLoxDb7UWdjJmfVXpE3BW0NCTrHvIeCpAHgYutDbPiBtJJnw3c
sRb1VLECs0B/4b+gBK06LERZiJJsUKW+sahSkDx1tjWa7DrLPDMBG/Bv8GodCQYu
GDyDJfpk18Gc7td+cgGUZvzQwcNHFcrWT3uv0k+sGMM1ikZhtS/2a6Dr5Ly5FF3p
VG5DJESmJoW5yVdXOBlePi1no5IHjqtUAl4H0Uua8QKLDK3QZEluRRboJ5Qwyraf
PgXND+hMxCkVNvMwrx8uUz4ynf3wt3X2R1FTtsw2YVEbS3MsB7cWDq6BGvadp0Lk
QNX7hDkaIpBWohUF8IebeKch9lzE1fw9y7kisVotXQV3cTW+gkOCSav3GFA6mqoO
OUrfI0sYK4sbQYyepFS+oHCcMCvdYnWEdnB2CdG3De3lCpVmwN3RG86NChyNajxs
5Q9PZCHFL1CVq9ICU2FLGrc/EiiqaNIlzdTlE4aQHGAfNqaJbd5hfd96p9DmuEG0
+wnymSUeLzTwMbkd+hRmxiKI9IbqLkwIhzxsNMl8Rke6zr/G2/MNGnf1k6flytLf
Ez/puEThqKCWljZszVr6lygBuHT1VVyuOVwLBKw24BAMB/GMkq7/aeAwM6xRneB2
xVOgjtzBNBbKdF8TxRQsw/4YXEWIEoUAaZBpXXy2j1XU3qhIcpltrLQJqKzMfufk
kALxyiSbMmzn55y+HPnK/I86NdfAOzwxHTtCK8CPnqiBK1zsVcAgcIkjc++10nds
ioi+g8hVKq+2vOXIRTjI15iXDxXYSy2zcEkc7tbmdwYkkuqqP/DcMURKMfvFTk8a
X6HYHmuGhOHr7IAsBf5w500TCDmbGKOKDE5fpcBOHJASRylSL7Hxzl95N1Ocjd2e
dAHlmZQivaQ0CANVydGQstU4AdQp8wX5wmjfLXZn0Oni4TFpe2mG8UTsi4C9z20U
tJHDq9c4HsFz2TvVVo6GVPKb3nNFxjgBE9fsDWHAAGRkHMfKf035+DWTFRG51Ek0
ZSNHnEvCXsYV7oAi+n3UoPIY2Qp6ejKDNsqsvqDrRmmzwuso2ahsPSeReTFfrZeN
x95grQ5Ncifwtcoz1JGaOedXid9QuOn14T+Oz1UVxOB3CORNSag1/+gnBiFLkXU/
TNuEEuAHyakCiUd6ree0yIOwjX22qG/2LIBvsBwNFXqQYXv3Gttpnkp7cSZcySMk
gi1zxCMy6tVyWr6u+T5TZ6Zg4EGKF3Rk+YVZz9UGolbFfEkYfI8oSl/YedvL0llQ
hoOU+wSL27wlmL5lLgLa/KPScy28HRL+pZ9UNaBHDoU/5MM6EqfYgwsxr6XmufdV
f/c4d/dO99ondVWnTXnIsxLJubSJjjDes4+C4tlfwgwD/R80p992hrJ/je3Pk9Y4
stx0i3uWeZ0iYy4beFmLh82CS8GeB+qFcA6A+nei7bofaN68XlDr7iWzL1h6QY8U
cZ8B5AUjQr4j0uJ52/D1kj++v8AtHr4Jrqp20hjeAhyCs6uEHImr5UPZPUlHHhWX
eEUCkTmW2zWQfdak0kcmOnDQIVy3pF12AcqTVAnk6GevybRPUtnZrb/VWdTnsBmA
t7qMzxbZbmq2GD3cosflmQtkST8YMWi/jh3frZrBvhLdriSXdJ4XHHybpeFR+VWi
BZk5KOPFmdbnHT7hamz/Qgu9kwAnmKuR+1Q25oO1Y5sAYg6ZhlRHzLz7KE0t/i+7
1dBX7pH8rlFeoXsCsLxAz7RYMRfxgDUasZSokHDGs6+GRVjh04Ie1XazSlAgxmNx
XtjRJJ4eaEXiap9RyFeZftgrI6DdSmz8PqMOS/1m1HH3O66Sn1R2tPPbJg0fB9eY
t6w1Zf/dYL5i6THvumGrNv9q+u7eo05Jb+lMjggpBzlMr2+x4833jAvyJgl2qfR/
87yb62uJoygeALTv3tnJmAqLkO3jOwRKVRKI8TCkJS41iGJWWAVHsZWdJArpaKwz
i6ghbmDtIZoQRfEAGMlLoFO3GWhz+r8tZBsy7x+fU06EZt5dLDIqOoeaqNSP5vqs
Cij/iCXlMpmCdalfk4LPNpIsCZALylj9pvFxyqoTwTrOZgq2FG9did2HDcpHDM6N
IXmYVfSRnMAbz35BQlqAKUCJvRnvYT4P1NC1oNr2ol0wCwUIdSdYavHc617bssni
qaYwor2CBhXqgnbF9rQsuC7UuYqWtGM/9YBRk3h8m8dQhJDRuuHCPuA3/dqdYpTI
LjairiMTjTU0R4toFPcBulBnnbuiKtcHn7HUc/QRhZ3Gpt3i9nu2pbw2z+tarnpF
8sIUjh2PnPcrZZPdMhd917E9dmog3CGV/edvTgbPltP7l1SsEM5uyKSRMXhWEnan
GgmvM6luwQpmr0Ji6LwD6746Hp7KUZr0UxgOoQ6lR4hgwMNYuPU6rKyFttEi+DzK
tSd4lGLjX9nM1drN/u9NF45IXRpS/buyzILtfWlIVFbnZnRfwWcwYTJ21QPT3FS8
yJyEnejgjGKBDfUUHIRcHUC1jYaSJrCpJcNfxsqzEwIws6b2C5gpM6viQqjL8uAG
dVKviI1aQHdycymqgz7WtZKa7mH3/r4lMAveZ2I3gYgsaLJ/el41v3EB+AHTLf0V
vd5u/npaHuujy3QufjL1J/bVzcyIccgz0Mwku8/xHWNMk+KHJEmqlE5CCBKPNkod
S+cEYtsr+Y3YgbQZymelg+xoEViBniWsNSDnydGZf1HJSLTFI/qOMVR8/5OZO6tr
h5tVNBSfF1LkUy7xAobn6wzAnYKPfx7ND66jmCSHg7wJp1oQUn2BmBQC08Re2bSW
DGi3YnfC0NTf96E14BZQsADlD7xcBMF+pzaOlsObQ5s+eG3Y8wyXlzV13EfjrThR
94Q3H+trPAvokBKzLQO2wULTEyoQMgIcZBPfb7fQ3GZFwSPfG1FpzTFzot1+p76u
YXYvwuZE+WmWPZTVxRND781BlEAZH8wWt88bNTZs+uBTTX7ZRl6oqi2zBDWqaVCn
7+o52ECWMfQfS+LM8caX7Mlj/gmGAdPFXLBhNJqwPz+bfWstsZgDyR3S+OBLpc13
augA6pRDrBXJReVIPzQI35OA7N3GeEslSngBeiA32oVn4YBPJBIK1uDIv8MgfRjb
LdpDFxo2oQ07/cyhVzzkX1EHzHwHDn3ITnQ2/BsOugZ7thvFtEeUBvwNf/Pn6O3i
+4UMdtGS+AQ1xjgkPM+8HHwIV3xQtj1N2CXBQ9F/CKJdBLMhtcY0I0XOR48pdj4g
nk3bKBBl+XRJP+CmJPGo+zASSPYsAXbgRSqK/MdnNiyOiAvqeAZb6SegCoHZn+m6
unL3Na8dPuwb6AIIATsW4BM721seB0SWiSej1dqe6ovkHvquIIKnOXsfTwSjfszZ
GH8XXumDfxsf43JULvTE+PfhP/WgMI4WXWDBZ/0tJwFbKH8+1FK12YdVIJ3nO9ae
yjHRlbQ9antMG+rcydasPEWVOiCx0N/ItXDIQgnPnf6lGVEaoiSLt0e/zRjvL5gI
oFpFpOUD/BpBlOgm2juWqI14c+TpyIO69FUe0R+JLWQBnrBiD/By1tMk3vIzyout
c/xj/vOCwW+O+mnAi8hhR3EPeuXlckkGQI5a1252ofTkh/WQqK2EDuSVdXdsMLBN
C/7R75egwnNUAHc9fFc+ggMZCynm1NYqanfTojjJi+zBqucGoZz/XeyLlca0x6ya
br4wjY9PQyFuOKbQ+cqQjPNtfP7zXeIFz3cFdxRvQUAZ2LjWE1HdydqXkvnW33Ww
UoHkYXiirD25gHkufdA5uW5Yx1LxVy9Vmx3hcclGiLVyRmDlyHUbtroIptrESSUD
rJdUkmwRtmDLImmt8gblFj9JxHfAjIn5A+Y7/uuMzomse0KGkZ9PLUGQ32R9pANb
OZMpARWaG5KCfqKT1d19kC725wpG+iZnrmDfkPTqC2VOmooiE2WMzblOBBSjVuYT
fzeY9TcUSqhRoNBQFq4CDulEPxdOLXUNwJvjkT7F4msQ8RcVqBNsWzZHKnhXPbVn
MJYRNXywhsqDaF+wZkwWFd5CO9rT6RKvBUwZqLP+aYCmba0tBvfyDTF2ceQ+/6K9
NYHVDIiI/bt56hufoi4F9BTtzGcv8bWv2BI4XWE2T63YRsJTYvF+Uu+8oOlRucEO
ym6wvpuA/BbHi6OJSIjffi7XFHKYp/uJrK62LADTKVUZzzXCLvWbotV2NAWiFqWY
BUej0o68MAsj/LP3rm3nDI+uT9rUL63P/HPVvEmWVmumUZYtF/0lXxp8HXrGZJWe
ARDTqlowli8EayaK2HvQ2auS8MWnShqOpFglZkhE4m03SBmX/qgAyEeK9tDxhWq1
3l1SaNVgi4Sno7Sk7rLRYe7OEDP9+aAmevPK6FWbEV3HsQEXh01YBm9TAJJl+fbP
5zKjwZb5oO/yRAyO7DQjxIXllBgpzR8VrficYvfSnCq495CasRKeOyDAdYsNXiIs
TYd0Go7ltNDWcYJsTWLo4nDfsKzvh4stZYSzE2TTFPi+SHgkic13JFLKs67zqWzO
mWDuRVQlcGNQ/0Ni3SV8cT1zVKnV3aHnN0cT32qnWQT7F/qMoFPPTzeiYEkRyCdy
bIIHz+xu4VP+i02OSAcVU2mSj/1IxeaIf2JJShvrobObuDrH9IHv/GJoC15X7TdZ
1CYQbpwbFbmP9wtLYYXg/C4A7PvbeOZd26ArBl2Vrjuo8S0ZE6zj+mbvX7aJtxDW
+M8pJxeULZaJWw2FT/kQYJEXAReW2SpfwMYYi92L0qQSsFaTalR8hbe5Hi6IcaDC
0ZiL7Hb5s4kT+K47U/N25eigohpCDhyZfvQ74a2aupTa2mkNghF+9OQ4YPWh0qFN
QO+XTJkGKOLnHMFjjkbY0/A0y2SUJh3540G7qonisc5e9PFJn/tTC7dSEzLHZuGm
cTMZix8vbUqXMNvej27EX9A85w+W7yRkqlyIlE/vafe+p9CHM0DTSAVZxKNf39Q7
TAmjSKKcaUCjU4kGVxuJ4CZdPIlKWCJvVhYIwdgw4kW9fvrqrEsfGIy2U42qrbUn
91dSNHpSG7Ppn+pGje9HBUaVh1snLLqzKJsZ1dpbuWWEsV4IOT70QF9cJUy5mSmQ
ldqQW1x1Y4TCK2b0WmEbEGEibIJT7IDg2rvuLBVqMH3VEEBAJF3mHsP8yQDsTfPm
12Lb7baaI8zZ/GpNcyi+cnZX0R7A4tZSloANzSK4L8lQnKFJNfZ7Pre6EaE3cCyd
zKXt4TSmkBpKdzuP+/jxK4hmnlxw+QXNBpvxcLNsAW5Qw4IDBgJ352lM57OXPz6x
ASCEaCZUj9uipuNlfHx88YGkgs9OyKbwJ1FnsP16ccoaCpLGQZSgXXMsO+9BGi7L
HmBKms6Kza3hqkpUD523UKbcysZEdGt5p2jGtgzAtHlCuu0uR1gjct77fD2QuDpA
pDdaCF+6iSPty2cCAr76bsp5E/ylvezjgc58AKYoCP5GDNhapH+JYJxpQhmQR1W0
ExVICMGo1j6WBbGzVtOs4ipVfXTVxBSZs1KI6F6VuC4mp6hJFdNyFK9uGckT7sMY
l57jJLRop/j4XXey9+PA0GeGZH9zOxCWT+boXng2+SaKS/df8ip9LIspb9wV7SH4
62iK10uhlJ665Kyxp0BUQ1izNH/HWbFTJWjB+pHGQx/iPKo4VMTT035IHG2v9J3K
Ze25KBE9aRIq/TWnZM4ieRmvQ0PNGE63ZhzPWxtIuHf2rRC4UumED8sPrlqI3qQK
Lh0LNwMdbJriihWqQDT25xp07NlGxf9pdr45dS+vFvKo+/JA7e+nC6C3PfjxrjVT
ETO9LCrxjZ8YUwtojnRT0HqQSfFePwk1HYXx8BwH5e1xDHInUwtE/Kn0Ih7x5N0W
+bFAekN+6tHOa2e3nEqrHf13w36Zvv/6bAScslu2+Fystlj/EMEwy2dfROJ5bHjz
Bm2J5FDas8HHAltP/yUAtO1jTY6loUA8OqezCS7h3JlvaHWRarOT/9oTdTDDhTjU
OmuwcwUUZ5uq/7cJWXR3lBL8dsspH0o5zlho4ke52OP7Z2xzjLz44vAKMKlalhMN
70nFEiTDuAI18SRZoc6UNWVBCprx9waC//IrRBynb+qVWupZUVHipd8pqgNvslfL
kQbxrRqfdEN164ACHF1T//iS16dkzzgvqCI24IYKNkS23iKDDNOyMRDkbB13KGgo
q7m6LDr3s0Um8qY1lCtmkVfvf1smC+vGOa9Vow6eOXuTqv5NSF5u4Y+4wUtbEAH9
d8suzkyTDhYIrFTYbK3inFj2+FaSUq5YWT6SZtps4Oe1DW/wM+9zp1RiDsKyE3wp
MYdugRSVIu4J00+bOAw5kSHcTCODS5s8DtVLnjYSpjfpxn6JNF7wbj3A6IFRff/s
LUuV2qFUdOaEzOHyIZ3WLASYy9JOAZNpP2r+Hu/K1UNv/dM7HUI8DQZoQLmgJkVm
vLlVjZMH6TFI1dA94PsnyPlBNQgRsQ1a44O/RyMcVTfHdyyfobkThO1LvMY3LJe9
r5FJpzP63t7uiOAKytycbkp1h8io5U+ODD13tnkzzcftFYT1YQpOIXDLStziRxYT
Pvvqgs5U7nKwd3+YPqPjQg6IQjNA30JY0nqIuGYdfYNmP4k/D/lz0LgQQ5Bsktc3
iGGsGCYCXfHqBkKvOK7M5y4MKKmoLrkBMZsc6aOpvdaXkumXmGEhhnpNZROwt8RR
YHiiHQgHZKBV1fEHDIyanrDZNSSCT+YPh0nYFKFcRSd9USRIFLMpMoBHYnlt78ys
gIEYOmW//5cL/YZxdPhls2tZed41pdy7lmBJUJ/52RkomXKjxdUB5XpWCZVZF1l0
NQUMi36FmNfnWn9qBeZh2a++xOXqyT6hF9yoABXjQgQgL675byngPkHXrEaBzMSA
IUOpiV4d01pg36OqXOmsyCkR3M3OvmLLCwo1k+QIF6j/YN+6uHMIuYPG6wfFaNx7
9IKsz7kVuKc064vVt1fK4buO5btdfPRwRHO8NQ1zJkVhl1kQjAHGsEBKH1UI/1ii
r7zFT83z1kt9rWXAKohSc6f8VKvobY3zMLdMScx342LrPB9zeDghpLJUc3Igl0Mb
Qah6rQvFlUwlHUkdpgCFSWvkewT6G+XAoH3cjDMaq6PjZDUZ/Gaa/CAap7ZQZX+o
7NyMFz7sBnAlsTLF0GzmxT0/YRo+RA9Cs/crZ3+q5Cn2SVdEvO4bwDPPGrR1WkGN
SYnQzGPjwkT2n5ZzwkD+dyzlUjbzZrqmOSpRa2tFM8xcLsPkWIKfPdhetmm2XRXU
vxxEx1pn4igtiuDtFTFXFSNcYtHMqoWjvWAtOwcbE+SO2w24RtcOxkKLnI6hKKgG
ZVPPXQg48uWsl6kSyqw/fkMbmWMEadH1ueOSrJcPj+i6HGMKzclNQUXu5ecWgGTt
kvKjlrNKyAhQ3aT7mLl04ht/qpYcMgz3DuVbclVyrcQrLbJCPIG2lbkuL2bXntRr
UmQlqQi/61JgMBPQBZCVYAF3332xAI9j+cHdligDkh4frDVY8/3Pr0Revsbhp1wo
AJ2IsltyWH936eOzDEnuKEkvlYtlQ85RNz+7Z6QQUIC5tjKQ/19Red8o6XYdU3XZ
nlxs5an24uPJbYqyAXPFiI15o4GnasWleV4pjhFyldjgxCkwI1Oku+Lpog3kfq49
sie3Sq4vTuV9ZVNFnO0G3N1FrKxTQu1OlABKwGnj581Z2Xx7wwyK89h4omQ/gkVD
4PXIAacPdZneep2KIA3i4Zk2NgVc1OjX7p5Kt/wAAsNDjB8axEzCDDHJ/mHPl1sn
3E5eayIf3NXzC4QOh6hsYUl5Db7J14T+h6HtyyTNCBX9O2xdQjTEPFw6On6uZFN3
F4hnQ+KsADkxsjlkFnU7pczAjXgvMDgAqSiQvipdEvLEfPrtwzJUbfyBWes/rYcd
YsovwZf3KrsehZbXWqIMIXjiyTYbJkmwC50cmtg+7EumN/lt4FG8BDdFdy7Vvg+C
OM/Q/Z0Dpm110Ij6vDbiK7brQRqcjL+f9kx+Xu3mZhO582vlsC5tuu8p95a9Y1Mj
ceQyx+Sg4j0oEhm/A0i5WJOEipghZtI90v6LTUI1Wiq8KWa7jNEbcIILtk8gO8UF
+NYEmpFV0O8mDu5IWdQeZ2sJBfPZ+WePyAQzFKVNMVCZu11DvaILI8LNbDTn/PYF
O9yA1PiRgYSmq/GHakhtaDpG2tH5BuQoyuQw+yHifVuu5BxlRuPV98T6TwwghU9g
8XVS27jXfulohU0J4sviLTEM68IAsItxQbFDS+b1aokgIM4+vhV5Bs1SZGz2zaeE
bJWfAO6XZnd8t7J17bG+NekevaL+ZwWATgXmdNpfhK878goufNZFNClw/yoGFrO+
1x8uczrLeTQDTow3UYzC2AFmtgVZifxp/ueQyAhQEMfjJBotl18emcobCB0SRsvg
+1f759m11tkFUXJvFbc4K5aOqkUsQUnkEaJCX/TJpW80nVo06w442TVI8+6L0S0J
Etl8p300aQBRHqgfmPufm4QAUN2O2U01KokbcaheW4ooTJ7GJDZg0NCnVeuFBA19
3z9+caRlft4dej8QCHiLcYi+7OG7WGm3p6++DUhe5mpVchoSsZp+FtiAf9GiXFBn
xijhIMi/YHOS9egy7Z6WAwhqhWWqVj9ELwRdazN3XKBFE/f1g0rTcvn1mSI6zlwc
W9kMSIFJ1IIhct4dPn2m/v/5tbxp41Pbq48R0SHA07PpSfX2YTB530wD218jL0TC
F7GMxaVAUeaLQLcd1B4CGdLb21wM5EvXzsYyvOD3EGAnjsb4ceDYA0yZtDOeWNRq
4Xn7aa5xWfDDHZSrcBik8rBH7dCGT3rKv69Ao5aF6VKhZD8H06S7p+Kzk+21S/Ju
pYKLEfiCeqzMKhTyBCv0cRKX0myPUUvQQ798zhkMee7L2PNaDTmIRtYgYUCoMLy1
E2WCU9MlJiASHdi/1AsXfoyno6usCPTPD/hDXZ7sXPe1D+aH+XlI2sebS7K4t1DG
69NRxQOhbcjCUSryASCuDCPIoYVJ9TD81m32y1AvGCpsOqB0XCs7BjZCcilyDTXE
AZ9tayn+fLiW6HuTogCB/nnHX4uSz5ixHDsGkkxsJ13/jFuZUZ7kKl2bBEmRdx4d
pNOYrh/jwWYKEwmoDhG6iwea3BAX0e+jwr0i3UBTI06gu5NSSU0qcwDyJlsuilLh
80HwrRR4GFiW/DaPxNhSvztW2EIadbHaaQN8qCIU2whkKV+fSuUqj2amMK06Ub9b
6bQUbbgxoJ2u8PMGjLmO7Bpuyue44rUIpPKgqKMHGX0a/OM3qS7aH5g/LrQTfPbw
gbUGDdfkg5TomB6HZBXS8o9SJiuozGXf58UMScnAJHYsju3A0GCvgjmSqS+byOht
bb0drEQV+0XhzbcTi72GSkzMyR7nNmg0cR8Bn/ji9Dwx1x320SzlqgWczO482rWI
zryNcjRy4mwdXb3cFL8oi/2C330Xxog1wis/u/mONZ5mHpwEHKIxDpmKAK7odMsm
ZAMbVRUh5m/PH2m80WIVFU5hh4S9QNEvcwFELBsw52Ogj8jb4yLWIJtxHJpRZBHA
gquswyQynN+Xz06sEJw6KZiDm01TxW7IYCx/SrDnmkeMD3dFvb93QtE52ybKVE7Z
bwCMNLMWU3I9bclzKwZAEehY4n7wSkMCxVSTWDCRQ5qMkZNnT7PtxXJEsIimrq+M
IfCaSCRr3XM2Nh+4owYjS/caLefdCJ3zona1G9lD+JVKWFs3lxbjESvS05ny7Ons
ClkvpShLonGs8XyYMkIpxOzG47I+OAWFHIspCKT8Mh7wCppzj0YkwbEjCds6agSr
K/W+7ifWh0Jc02MhmO+ZHZ/ZxRr+fQaz2oqqOYaq1DAzNjx471a7A5RRRXOHhtpb
+KHltV00Xf41e/m+GEMVlscG15DI+cZ2v0vjBBqtN9WUD0hqq36XAcdZYFU90/Zl
lZXOqdBq69Qxit/Rkm0KK+G+GW+n7HlFvytvpHBTCSSaPZCYq6uOzqEvuM98Dfm3
zZYV0NUZ+A4MjEWetpmr0kp5+V+VoIpFLQe1kyQZ0MxUyg6lf3OpHXzVqF5RTyyW
jQCTiUtSfm/CsJdcin5S+55I+w5Uws61/J9wi7EuYyzyGyPuz44xgXp6hnoPu+Jq
3y9rPIjCwy6qvZVcllMyW+f5IX3awp2Zfl666yAkC5pejeIElwgAnU89wT42Dmvr
Ch0/o9KsthF0c99Q9FjX5a2TreIlpnkqyNaYxmA0zZY0mDUCC2uG6o1FdSOZDddq
e+jRohXiwvSyKp0HN+kI8GLPMgsbk7R2wzo2dVy23ZGN1FBb0kiHfnLLAUoXkL7b
/fKj+Z+qadrZ/AzOPp8zpsyWhc5399+E7dUwNjlbnTQkrvbgdx+ThfsViVD8G9s8
WwQBwQXh9cojhncW7QVnj4nUr0FulcwaTtwONfRsYnXryQinbvCKTsvbMHf27OEZ
twG4Fg1thC71ScO+dv8U/LaYoY2Fc2+xXb9kZw5VUQPF27ZIyTHP5cuDl5qpQuFR
9oNQndfsqB+umTI8bI0LuHT0vfVpwlITPCMIEs5n9W9u0Mfn+zmJ0boXJyVKle+5
EWy+ToANjaNEloGcCUfHT3KxdEw8ZxOpCKEWuxnZEW2QkOjYVtBJ3MUoW++JXEoK
MjaSQ2F7JYuL5k+24QNxHMmj8WbKKrOfHW1wL112QcY8ZCRJ2M2uIcig8yJPvQOx
/VGsca7bZ9tU8avASDXgCjlBT2vu1n3l66KTpWqSqYSUBhwyKpWC6e7ps/EHePXw
1Y5Aa9a2fGCx5l5WqBqWmRz4LS2iGawDCzxjmV8eqnUtJGXh8t6/vq4RkvSAUwe+
N014XqB5jqKdZUy7MoDqGawXw0V+YvPpt0CEAt8it/CM5RK3SMHS+vscNCLsCi9H
FeER0BIHbRx75/XIcRopObugxu7y9mMF0hmoOruJ75M91oAIDZRW1jMDWyei+vu6
sYRHDr1ZsRAML/YVgLQC6dcWU57OILwMBXHCtQYXR6F0XwtqgSKbuVS780dZvba6
QrHAyeMmor0/EcnQe6B7yAPd/fhbbS6ImaXwzohWZJ+iHcD7hpmJyLFAaZ7+cTmT
s8LxYwu3kRC7k4EKZGcNivqcVv0XUZPoXAUIlI4iOYf5BjGaKuC1CDU1VLzD+lU2
PhaHiFIcKvj10PaBEBUo7xSx9ak/h1qxeGcGL7dTYaV+t6DokkPwLKSpVKCqEVDW
nvtQxRnxp//jry5qC6aPR8GSSAD3Gdg4ECohupOfAXI+xDQtATNugDKx2Y1Y1MiU
GtuvS1/jwdnrY9lq8heI63ik6nSDU1gjAHoUEC5/pk0K1aVEYVyWUD0MmUhlY6dg
6N0lszGbN/Al/Icj6jV9zxfQxoIVSFSVyOBNMH4YyQhA0ncRQMuT+Gzy0E3SV2Ea
UBCbvj8ooi3Z4FFaHSEvauZvCVfKofLO+SEd99XlMpoSbNNhuUWKvGqhm7YcWhK7
3XoUFUQ7FxUgh2FXKGOM7O5ssP8uVYtLTnHOkV9vDqNJlffaTUpz9jyPws9BHq4V
QcToYuK1G2e/P5sOTt3lU4imvO0n9stJT6GuoDrj6MW+8GZiVdr00AwKxo2xylnW
OrsvUL2RkPqzMCVaipmVtQfMplYBzmRgkiX9MlpJ1tmqA2CDsG/hwiVPsV2yDF+B
9gf3KyK0oYSvPEjTQEP0xTSjn5GpA9ju+pux/CrYVSd76zfzB/XWcfbLnwsIos62
SlviqUofegydFdQ7o4W7soKO5GfLBjCHd5frZiLI4YuCNh9ft/nq/jrZaqUmXyb+
wGG/Jltl/ciwZ4YXzaxBFKlOgAiQkb7NrP4FO1Q8ZAKCWSxHVVB7Q8ntC6Q07Tml
MERhhaDkpMBdrezTz3TuwG9piPF77O8UdLuNrl6AWKAUEbccySnToa8EtzHcGjZo
0B3bglIRmc1uvtrZRa3Ki2SAXjYfajubqjJdBQHA9tMiuumKQ4s5L7Fz/tbUjiVO
0+giN0jRCf3dqlmWuEG8gNinSCI7uL5md1/eZ53jQ//kJtRak5gnXtUvSO3zTGWj
tgBKlAMA8s9sTJBVpD8EfUf7Jus+P0iyeDIcAeRPawD4Gi884Og1IRF9B6IxN8h+
4td9rhRz8CB3ouBGIFECybo1PtL/5EqaqhvS6y+njRUh3i8QZczKKoBKVATcYA5D
tPX33Ow1iQFYdinyb2VZTGQXp2qvHA1AMF2UaK93RoE20ETEeN/B+/i4SsUvyNtF
639X1RuPPiEdQYm+nttKHhmyKyZO7Ftq0FP+8GtjJ+aQ75tejd6+N96pDbn7xEqV
VcHat1hxlebqPuGjLv72Yh4vCjRtu6iNgewBwPhdn2f9j8bIOZmdqhiH8n4TJUpZ
Wc5UprHoe3GSFx3nC8V8wI0ptHmVMGagyLML2cfnImSkSIUgwYKnJs5ZnRTiyy06
LBVwo4P7sCgrP0XIUlsU/4wSePu3GVJc/T0J2dkYo3rlCSIJb/5Joxu4bm9NFCI4
jQ2m0kXJzAmCtTwh6RQVGOxZ/UCqMUl/R+d2oc3DSqqg1WOAWh792jgJVa1MjmmT
qZ6NS/U+bFmBZGIvUS0PGzBLzxmpMF5TKSsEh5G4NBSqhplndrVGq1DaGlnSyCAP
POr4ltDmD0EOiJZC8GgR1e6bLMEoCWgF8ZbVf4dDaH2SbsGG0LMeaWgxz5aM3ZsU
qtu88ZL8E5+RNd3nb+fAMENj8Fy0UoOuc6KcBHmDXl4SD3tltYkDBSr7wiME/51G
QVZ+5h6YiwAoKhAkMrkc3vGvvt6bMYDZVr0c/pmCK4tq0ncopDhxl0dduR0S/jfQ
XJ/EHHpu0CiTmTjbyF02NKLjgO/ZhsP9wCq55h5+CZepepWAueT7XeBdqzG/vPh3
1aVih2ru8q/1tYWuh+w6NHRymp3QovhZhoQdo2e5ojHJEdptX+ONtEQoNjpTmDwB
Mjp699RMYDqZ9e5ilacu4537S+B7VzgmNmtngYRm+MEtuuoOJ0oK46XHxQkOW+jT
9vB7ZHDvMrbT4s4rlJTdwiLWEozcsKdqKysfxnSF4ekMCbwmuSbjiJTU+46Q4rKK
ji9YeOY8EmJjAus8SdsCxwfhEv1XfEYC8cBglalDMgjl3oCBTuU+3cSC+3X11faF
J0FplEWNaHqgcegqQnwgPq71AjwWkQgNNftOXIeT3+DXs6nJ30alZRCFBW51HNtq
67fIbyXUKQ0gL2LO4SDHgbxkNzuiM8t+yLkT2o5oGUByCNHjBmVDCMjwlSJwpoaW
ynog9lvPiEwYClOYfQHR0ElwOuStqGRXY52T7F8ZL5iXuwV7yTboodlGQEMNhZeN
osEi9sD7h2tArG9MWucRdQLMIji4aAKEI3/ZO1E3KhBOlTXiJNlut9+ERqMOkqir
UPRFAdi52urc+6kGe+lCiKi1UOKcgpJBeqOIuuAwWso9FW/hLipFebqvbvwleys1
+J2lmfhEesk63cWifWsXSDO0t9sVGlPYBsJsTZmO7mzOeGDTIwBnAgf0fwGE9Vpn
MSfoyDB7Omx4EOPNNftAaOkkEjxvRYA4Jz6WHXE1gWG0gV/FNWRUQk+SoktXII1E
JQJDJA8wpH1XVaGUT2gJIxQ35Jn3hwXB5YI043wQQHEIPChpF2bBEV9FTuxzvyim
Y/QyVDCJPbtCzX0wZNLOghvaIW2Olp/snD5m1eZEd9wItC42LaOqvfTob+JFDbIS
JIgIVcqF+uASUdZ5qcAiHQ3NXaweMfUvPQvVp60gUUM/3GQfWsWuUhiY6brlYkLI
55nWF5Thsf/1OZDiKOypy2UouGubP9CvgrqkNquQQuJBaoPn+lNbjdEAYlIp6Y4l
ftT4RjmPR8HkJkHwhh6CpYPotnU/nPtUwF+VgPXxb14a5mmrOvgI6WwTmEJDHqHR
6wO1jtesWq5vVc4qcs1pqQJanJ9Vq1yxoOBt9eYN8GGT8EW8o7GQSwi1AM0VWTHO
ss3WbQCZU80V3X8e5rcd7ceJcuAZy2PV/zkEICmE7HAJMxIbBod2WAOttSu3d2xQ
MRcUXI/hcQ6tI7puYlZwb7r8bw0VgdKUI3M4W89a4z6OsHcJy3XOk7DlorrpNcJQ
NUn9bG2vJHtOvudsUWhN5z8+zlrfdsDxuyZWtWZ4Lk6MU7tt6ii5HqTU44amgawu
ycq0BNvDv6wx44wjJd6nB8etDd2ys98HQaxCVVZpH5cU4lqBTol8WBJBvsgHpTK4
r3RUL8QOwsL58kJ7W9zJfL3CzPkp6FNs4WiaIBxVfJAoXZNrwOV96PZAyoBA3v/f
tiEhrzga4B814C9a19gpwuyBqM5cZZ8Kdi0Uxa0+TYugJaajlrq80i8mGfI1P24D
fq2WqiCCYd/NfENxsYWnZzN02kV9uz8W2KkFwCWyCiMrAHb+O/b+jRLbfXaKzpLd
0DTS3CXu2cSBr44DjAUjeohvnyI/Gr4gj7ameCwTbZuKEN2rGqrJaTmVucLrDzjL
JAl40/bmIyskJz83UTvnS/AzgzB/d7j8R8G7qKfq67g30Y7HmbDETd3E+//+08W6
StLmJDwKCcotZerSj3GwoZ9EcNwlLcNP/a86yFhtz3CyKe1zhbqJHywNiFe/alLL
hnBPwQM/mj7t6EZcCWthyqVzERju8LAo8CcXHBKYY34RwnaU3BlOO5d+FfJ7FVl7
zAJ/CSbOPM7rO2jWEquf+gU2ltQSwyEbGZMx8towG4REVHSA7FIv1pIQ/q1QsxTp
L+7c+raTg6o3983E4IT8GwlQl//x+soRaMMPfyJ71qEmpwDDvJMQOTp8Fhci+aAy
QNhSEOyqV/HiRGWOIb+yToOEdO4sgoTVzFykIP/u3uwV89e5xBYDLpo2/e+MjcEd
/H2yOMvR1ncx8MdD6M+P5KcUZVqh/VR5E7/jjDhMILUWvloJCcTRgZKXaMIu2qwt
stg54G7tBqQbw8unM0Bll8sF/dWyp+s8htOuzXRIbNniTIV/EsNmyhsXe6/uJVoH
zFCCrn9/59qs/Ml71A88jUb1ziuLZfOr8z+A9m6o2ef8S93kwQdWeTjC0OytPzgW
YulGWVHQMf/Do5l70l72vWvVtRDclHkWQlAjDnW8OOLtvdFtY/RRCtjKzrJ9Hi2o
06MtkLvbnc2EHGksoFy38h+G27jnTEoS2ChEHBjnatzBTPigVWGoJ9U1F7hwCU7v
JqIC04cyQGpCuFnP+jFD2CznFNP8Nc31VavRCeIYVJ7k7fEqJaISJ55DJxHHn//c
BG6qPMBrC9JllpKS2MjrqQatrGh1JCs7gHSUWOF7Mb7/mTyFO495gJbE8ehXEDsZ
3yKIRSDVdk/NiGNVD6ilHCl3ZmY7PlHSrvSyIBDNnJppTY1cEHH6pMdqqswFXy1f
3opMYuEfhuO7yNWyGKYdts4t/8opWKDDj1L3aMDqbFUDIqLoMCvIE1l2WNgUykew
Ilqf7folCvuHoQ1dQamVH4Vlt+feLSAg9SoI+PYOGxdHsJgssVimt+6FIUa+43/j
hlYHrn9kOxECR5tafCcXHHm/iu0tX4xE7mdzMIadfbYH02e3TSiKLOxNP0pgnCFl
gt9E+xR2jI2QO6qv3ssoTDp6UxyOqaDTNCu59U5k7HRKgQcTxowN/0l3Phw8pjpw
R5gPobgiv8OYe7OlPmI2SPvLaO3sEMPbdYzzbuIP/hr+TKE9jqMHTevu1QbJnnpm
Vm+BKCTFPCFNIIza6bzaC27jFmrvfDJXKFd5fmTT3uU1+CPD9TZW6c3rQrZQu7pg
4zSd60liP4HENNUwBlXvXX5SVkmB4uHglxCrBFQNVOqHjbEKUXVOhe8aw0axQ3Ct
gfs0mw36AE1MzjNrrNgyR9Bzf8JKWEeNHqPMNfLP2zGNg1uUEM6E4d+hj3pDQdRc
0F3rgN2LgzgV5FaeZgZ7/5wBBo+kYgM49YinMepXw+FnKYPlgtSGYARu5SqvukhM
xmukIAiMB29OxXO9BU363Dozo3F+sP9KOnS7ORL41yjSwfed948jThAEyXCM0jhu
xbuIww77khfQ0HbrYY8hyEVKfiMolC2Snt2EewDYe65BSJuTjxhERj8WxIZBfxr5
/NWfhzeGgiO5Xc0ZOomkjfVQU+bOHZIU1ttUhAB5H5ZO5FgTuz+XLTukGW5e6krS
IBRbTVV/DS4XqbhNR2VUqWEQJBMXofm8R2G1a/KTALTO0InS0G628Qc9ZRWani6P
1cJpZO8WXOi0+o39wSxi3cKCb5ZlsBw1kzIm25M4+wYrdRzu2dDIcxqyIakyLbqx
wG/pjs7b5Fjahkz7VNBkyicTH99fJVwjGHCp82lCnCXGSkDc6Q5FfX2O4HAMlyIZ
ulIyuvEFEjHAYuqNTXraQP6dzYrhl99GzoTOoahnpJRyIaUV0rHd4NydbGDy0x0u
u7TR2XKSchmp0XshYsT1VbNZ3yw6VpIAKd+d2/xr8BaIa8oe3CnBHG4j0YSgoMXz
nnY/LEjTC+vocZfVoMfSglFZhgYkR7rbXvHnuDW5uMlYTF5xbR2mGr7tgjbkUkeY
wIsNeGLp71iGRk8O5Xa5h3A7M89xgqexPsZVve4dlWH1/C4LXId69BJ36xIYQigx
at61Otnc2+zNBbO1MQJrujulamNIfnDYgLlnKAifn2k+zZe1yZfCxJoa1rSs64qN
JbXMa2uPGdMx5F/rqJq+dWZappHfJTUWuNIMi2AbqYmI3zQbz2xG00gHRbg3R5iw
mLs/0Iw6ZDYqBlOKhOsdJ0z35QoYMoy1yOhUPNb50UMfBD35zhq+Phn/OFb1Qnkf
cCUneBU9n6OuMiLqBi7Oro2JXGbnguNsPLy+opCvz7PHcv5GphGBSWtjdNntmeI0
A4mevb/HeL5LpE7jop7MBEk1foqrNDBYfyzqwirJmiS4pBMng6E6OSwdClPYm9TR
0YtWPHWddII/VqBdA9v7hQg5GPsKtXulMQpeIgBzkv6BRFeMmtdO+1WA3mpC8Eg9
czj4L9m1yJ6TqfLvxwsFGRCHTtHCfvIgIDemsIBQF7fCfO3qP4FCqHgN3Lt4J7Ve
KGkINSqcSpTY/6rxBddK/ExQr/tpXsNZKHUm1Dt2fSw7fwoUpUWvYoncj5aENh+6
PT2yQ2Vj2dGw+BVOtiQ1Q/XDdDyaQLODm/e4kAjBh+3m9uxNm3QEFDWjFCyrzt1a
VOeBy0gda6kXp/7llpBKLtnaaFp3hK9sJWRduQGf11Vgj7RdjceBAMW2YFaeaxS8
QCDgk5aHhZIPBh4Sg5hYMQjiGLRe41Qpc9rBdAJ4RxuwBgKBuHNrBXv8U+Wce2WH
P/l2cl3HFUIYa2qJd48CVuZlUJUR4FkvDaQPtCxRqqf6e0WVdiZH31xujf2NtQGy
ryWoQXZdDz0xAoWl1vzwuYnL1TSXkpjwNR7LyoUqqt8TuCYTj7W3OL1dl7FeeV5W
n7PqYU5cTACRMESOiaYquWKw66NSSSesgPaHWcvcHl6K8+G011AMWujVifB8HhsK
ck4fWwi2SXWYGnoBx//7xdRliovO25eP05bjHaNvOvM504/I7wr+ApFFaaZK8rXs
dqiD+gfZg6vJ+dpzuw7gSuwqLTAEg6K+3RSL7p8Fslz+9CmBaep+EHT7W1yZ3Fvz
4zDZftRcmJTlO3sqqmEWna0/PDJCzAkik5iDrvkV2GHl/Xwl3TSVxFZxoK2GW9FO
HZ/qx0XM9vjHVwQPE86YgIFbq1GRmQ3f1+oqbJYLQPzcpGwZ6WEE609n5iwp5p0n
zZ3oDupxkKrRQQp9gEHZDkPkIbadm3NY7MU7ZJ4hTn6sUbbj3Ikkj+zej+zcBDY2
KE262BGsG5Jb9xlFtbrRIGkbhAoucxvjkp4uhjvtZyr0HPbStwuclOiP4osKJUH0
UuEKfjh/ZV4agPaJKnm7ZEUVVM+OBnQTNpgPYQh7v34UiwpA9LXSzZH1TJKrPVo8
NPhFI+nsNKAMit1yr4gkoDfZK/y7tPbreTxVS3cZXs/zpRnihrswVre8ES9RkXdy
5UKP0d9NyQow7JoqIt99v2Y2SE/F+lGq5uRkfBP6z+UX7pjkn1GcaWT3AXUM7sGn
YnHyThKdZBS4gU0Kzvk1dBI4ZU0C9Vin18lmXItuHvmT6slI40WGu1E3GxgsR/86
+xM5eW+qIQzXUAXsSTTrLBs7EH2N3eat9LtrhcFW3lkVjKiwy0ZxOhpD9LDS3IzR
+fcOzvmbGVQ5oIrvbgs3A8wEHvgP+p151eiGTx3K2mZj+w6oEKFNQCdp5sONDp3T
sEBKhwFZZlzzFBbGr9QxQIucvsJzpzBktc3f0P8sp8cTB23ygBhHGVVJfl186zBE
GqMUlcfedDPmdSJt3muAND2YYZ0XI7ZEd+HzmRPUj51V23yxlTP+f/YwTx97ovXU
nh6EahRwUCVEF3v4pxlYtSv5T/lZYs1a6c+uySMZlF0LkBpoaULh1niRhZgy7kQU
Ind2KbYYPaiBkY9p+GVYNdmikb5jsoy252fI53mcJSI36lpvaVGYU9iRYV9AhM76
MXAynwtK3Rzp0pXCePFD/Zdf1iMM5Oik4n8eEWk0c33xZiyU1d3ZfERJeMVbjw/I
7ek7AI3ImGzVLSMrDzBtMBnsTUWtrX1X5j9u/0vsmsXSMRxT1WxP5jhME5YSyu8e
QRBeQmyjIvDsCnL/JmRxpw8qiDnEVM4+dk0o4Ejx4B8l4TzOGQ01PVckrGGgBWAC
WLNpywyhDGUURMxvZRPoKKTDkzuFwhRoGhlEPxq8q3izYxrikRUTwmq5ggKyH+Hi
75rdPoUBE4VJRUUCnmIAX6c6P14AvWPivSYhFZaNystnXF/xNUO/STjwhoUgBtuj
WEOJIx00Xda9EFYXOrSVzATBHeCJ/ho+R61mEZRfIeP/DlLnJG8CbsCEQlojNEED
alqaL8Pm81GhLyqTyGB9oc0Y+lYVwgmZ+Ai7oIpUglhTvLLqNPCUggcak62uzmxX
Q/1r1Ca7Qx31nxva9mTmPOMb6sTT1TqxU7P/TJDvQVvMo0TGa0yPFVbxIhV/cKJE
KOPp9ijIF3cmBvI+gAsMb0E/cr8pi+GqnY41ecYguX/ImLPRUj+w76kRtAgLjuXM
H0dFOX2hytdQMXmN0tfa5Ujcsv/rUVYABWQa7MO/oLmWOmBDA/xikRl06ut6T0GT
uuBLLoG05PIbvEbLqaSXMy6TO7L/EPL4tz0Od6lwJ5+ufPKkxryyLxgnY3qDzYsJ
ET7Y6Qodxruw8qMfPXwCpZrnnofg1C9lv0eqMH3P7rKPGSImPmek0xNft52/zccq
2Roz4oy/h5LXgduxGFATUQseNNHi6gYwUce0uASFpGbJ6OA8KnSkY0bZjr0urT04
V6Y4ugGKpA9wC1CFUgX3+BlxVLsi/tE3DMUDPlh6FLvnjWe43YY+NMAGUObUBOTr
1WneZaAXYaLtT6WHP18AFWvYNzCXsVIUIj0swFyCo9eC4kLJ5JSk5txCnJcjtoiL
jUKbyaMIcIvnkxybDRaN9y3kMndQaq9NzPhIm6zXOTy1w5xvIaHnBr5760bgYz5S
GwCLi3uNuOXLgfiSVoUIpLS0xd1FT+IGDVDbAcWfEvIipskuMFpE+O0wMQkzY8+/
EqK8TXqZqYPnWQuKVpHz6SOOX2lT+SI1qF2LVL9lwa4KagUG3WnyhDfBX0t/E0Qm
MPnwNx7W299kMPXBkuxegA+Xvw2M9ED9Rc+ZgOQxR2RiDoVOJ66RN6nHaLyAQE0e
0AGwkR8MRXyXtmhfZxqb4ylPfBd+gIVb/fLDrLp1OAfVob2VHnEKB69RZ/ph4ys3
38xISRZJSRBe1VDOM/IUJveoKlCUsU4mk0xAZ0fClFPJJOAvvem9PsMhZ5yBFEZr
vJHb+wOSrfk/EtNVhsoOkGSNdzAsmiu7JfWwhpMdF7vDjXAzhKl6bwMjcYnGmRni
v3yaMMR1qkq4am8lrUWEjF76bcuGMTZfQWD0w9NfZZXkxcrXJtIcOkkJKwtWEOta
c13PScc/EsPB4Eo/QeTEukl75OKmJQsjucbpzDWrt3CEbTgEQB6lSNLBKenxAoXX
jrsu2NgMjctsFsVYz83eYaX1j99ajx2sL3fphbdSULQWBzIZS6dLrzRrlejDLiB8
joD0G4BoFgpP7n8oNPev3mBT4GZ30bPtunyp8sXAKV1FWrrNEGATZxxouVh6jqxO
cx8zcLXbI3bJ/XLzcbwnpS+M59q72z/bTmmQgQg8Gg1rXJu6ECuIR6DRTG4RMidg
c9GHKFef3Kd/I2p0C1cGwaSrWcsiSD9Hd7JRq2Q2HaIpW6BBy8eS0EDsIZwJQCtX
x9Gy+pY8asw5WvgwY6+oZE+0wA77XrAZXIzQOyV9bUKaSEZSd3LlyiumM7BawXre
rHxgXpyemcYWZB80vR7QsGSVbkJJkZmRu/2BK54dxvPTiNta/KiOvW+NrlTn+gP1
+gCszaQLQjRnm15B1GLN5oVilbh2YgSQ762+JfC1LHHhJ7E0VWrFSAg6vGiEF4Nu
vIZVfeEjdl2bNExElEJoL7ulj2TZzOvBdOxciuudsJSxOtgGn2xeKXEQKfKHtUyu
bngydErpoPIXEQnpPn0VVlmpXW62EUmObm6+AFfkEsjIDj5+7p2c7gi6rrdWYian
T8nggeB8SUlRqsgDAwg02HZgPKKteuuIRnLM8CpdAAj82yxJEdCT6jtsmqKl0XXY
6UnvdBLSZoLlXEevM/1wnREFU58nUl9c1iM9aqAip/7DFePNRbrc+iXkZWId2Xvj
3FDYiQOjdYh60G4o3raUVY9ElGKDpXyBFxPgekTYC82cuWxM3sDGNrZHckeYN26L
yCF7hKc50Zlmo+VTf1kxP8we4OiIb1XzwdDPm6j97MXvjZ90AHrNuWcsECFWo2K/
YKYxeeeWkCzsmlNaRngfCR52lcOFri2EYQhGsiZkOVD/r9kiIcdyhOsIeswprZGe
qKH0jpm5qM3+46VFAUfg4HICqRaRPdbrKkzyPv3X3AA6VDCz68SFc3MVlhBxOGbT
mXWEWUvsIJu0OXyF2X2RQrY4VjS3vker4LbE8zQiV25VM/dKINVarO3C1+17CanQ
kKE0mCKFRDLV5MwqjIMfLkJpvbjTUPeBZy9JVfPWW9zvdbAJ/kmIXM2LuTlSBe0B
q2dIOasxpt6QiRtwnGr40HkZKL/0nukpa1oeIj4Tn0rMpAvhZq5IH4AJ5soywDJA
CYEr22ZR3Kx1s/6HUNuQ7p5QtkmKJMpUZev9iVjo8yTSMn1zJbcHKbzJOeY02y1x
MsHMCRaAtMwq4kxtXCeCnc7d/vT2oob8fIXp8xgLdq07nf9v+/wd0LICKfHJL0W3
e9I1FJ2kXsAROWWU4C8XwtT7Yg35lJvZjnqs3LcMCtoPQ8Gz5r3sRT8j+sNKkOnp
4LZ143G9Cnm9U2KVkfdPju3jRiX1dyhBdArywAMgzIrhW68geuvFUhVmEkXV3lEy
f4knnGlcOsyXe4XjeGGPScDN9D9ReIZPRhx365f1DjPksKf61FJUI6SDRO+ptES8
+K3bDk0u40I8A2FHU1uahe6BSnzDznAd9Vsw4Bp1f6rh4CcwZ+JlsmSz8NjK+ceC
6EKF7e3xvV1+L0ZXl3AHmA+Z4KoSna48eK41xhZg49tSn+cdNlkgTDQxh/xmjU6z
RcXacKgM7ybei7wqTYxpapiruuVTX1yQuz1z3tOf/CuBAUTg7Nob6XcdNzbjEGuQ
gfjA5efLww3cgX6j9rrtSqLJSpbFpwcJpaGFXFg4gHk0+sMLTK3CMmn4JX40txHX
DFFW6ZbJmWlVvKsx5TwXjdWNBjU7EMnLEGkvfYpxAEJcIhnShChVeHY/N9yA+mF4
Jm7ZsJsRufIV7JANmNbCYYOERrK4fAMh7DRessRvlChVmOItw7tYZFkbwdcKR265
miL8WGTLSblmZWqoR4xcd9cQ3jP4HCLpoEU4sfQ186odqCRg1lZEh5ozXwXe7qqy
klg058btXiNEaE4b/9vdbCfPOicJhB/ov8FqIn8PhATABFxBtfVOloQXRBFepFHm
JHayDSBmjDI1gJwSLkHYjNkdEoJux7XAYO2Y4ETmRzT5A5GtctzlWOSPUUxqb0qA
lfiZjYwvRGzVkPFyXq2fcGaSC0GcjKuHlnIDzXpXZYmtfWF9i+RjTdyJMLihaAhQ
CE7R4+UIctCyfKnAXDQMhviUnl6wISDeHoumUirSCL+gbcGJFF1mn85ZsSKuWDv/
AgN+KT4WPNwDYuD+BHZU2Inl5VRKZ/I/hOsnTyDI6J/ORY/+WAtB89Ve2+VKDsaH
ypmU4ZWSpz51eGQnUd6HnZEuYO/Yo0DEGnT/FG/fgVKPdvYvCNSOO3wPVzSzqyNH
SUhQJTLidd/410IVCCtXIplE1TrCPqFZjzHFChEAeBfJRNmC3JtMj3hAcd/rzHGz
vwvkhTOX/MIMbrKkCLEqOWVdoURuI1a/sS0GDBGsE3Den9mKYK51HWRrmtextohU
Mx7uDhMTn/eL3M8y9jaERRkMmdO42/SMjD6Rvp26B5hFgjJyaKVLVKLNFVT9BHSU
9qVAEoq2w79UQoFGCac6fKV2ndLdJ4R3ETURbQOmmNPeCyEAkj2AM+m+wWh/OwfL
4Yb0Np89F2OSe8aob4JLPYRywQ8zV9JGtTlkmTK+255kykm6Hm+ukXWFxMgoaEJJ
zK2ODgsCtdJYdxKVdsi73PmQuCrmw38RR+7hSbj6knQXLAJR3sVPklCKov2PbodV
BD8szPYQsFTmZ8C5kcTy0lLz2ousIEesrjdEYrcdBEVQjmgmtLTNxNnhxNjYxHbm
7SCLIQ2N34hF5WFEKO0X1dQwQS6bMjSPoWQc5jPJeMcBigJmMqNZWqWS6T/7joRl
r3RucCa3sO7RyudF1KbM4OqWa5QdGPZGEnwg4EYpRrQO1Q+orSBaQFCZ6/KLz8Yl
w+4n5+Gvxb+kn36RwhpRymsoAzYwHa5N/8IcAqJsusIxC29Tf2YcPZhNCaTHZh6j
xWT51M20gn2uFOGSWXCqc6odcVLZ3Tbmrg7pZDIYqUrNiAbY4pLBculQeSN67r0q
Kib+PgecxbUmrj+jnTAJObeOPot1K7lKMEYuxZ+sNxx5ve6G0ombEawuMilTKo/8
FgziPllrrk52KnokPB81fxcuUOmbQZo0rZdUS7hBbuYOD/KTYk0gOeo23DAGMmzH
WQ3npVyCuEz20stoIr1b/6HEwuX/9SDBzrHFc2mTCAwHc8s8Qz5CTxdud7UC8c0Z
Hqk99Vn1p1Nf3yUPyMc8vJkiwSG5UOOx7JksuQYa19x9XKG53b4MJuCQtNGfcwcX
tjQLwBKT9zNk7XKbvX++O98qk6/BB9OsyZ/KJWGqQFRrEj7MjxIlV3SdGIlpjZ6J
czWt93YWCbVZ+VZ0rPsWI+aokdGaizz/x2p1d3I5FFVLd+YyNdVPMj5qdWtOTyHB
equBTsuGbkHpWSGyYNUoMROhOpNHIm9af2akWHnMamz9UN5VJ9LWvSjTDqk20+cy
pHfxydEqjG2K3QIVVogMk4VSliWlCfdMmuC56TghgsjogO8kQrdJe9zsZptllPrd
Fv7r46wEIpkUoIawqnXsURa+6B8w3F4gf7nB4UPkbTbeppypll4/TpspHXosq/xE
7yzaswyIjIb0o6s+iQxPSEqxJEJbQbBmESKr12HXR5E4oTNT1dorl3P1XttLTTTV
wmW+b0F7MJO6dVTgSTFpVKZtculV9fSglRLaHbHv+FSixXreX2O2YZW00qdzLLh2
v2jS7SEAjwgVSQtfVpMbtCXTWygSH/EBi4ywu0frSaoMuWQkopPKq4OArRY3HUeP
Gjo+8cc6Is6QfBp00ess1tRbfbVXv6KZixhbDuahXu8MWYNqHuDd7sG1dnREe1GS
kZN+ElmlBkOB7KXU6T1Sv9xM/dFfBQqpcf+8EqFmzYEgGVyErmbs0vLGqouZWt9w
/mKj8MGBl2Y6WVZgep6bYwtCAbOkqxt1NRrLQZhh9Hhv0GHvuLn6QTDBjsvn6UL+
dD/rSWzvRcHvVYqH9ntK5nQwE8M6ltIQSVnOG6Z37L1noaxoGUcUWc88UZXR+mQE
hKhL9j9iMEb5zKfTVSa0QSWiI9FW+bySd2hvIEoRvtZDYHdBzmlnVjMbzUGIDN3m
Y1BrztVug5PJ38Qa5aQP/3YzAaSjDp0Ka/DDXh3eInAiwmqT3VIW89pVIZithCtI
Ge2b+uwHqHlTUFDBKARd7jQLjaAJwQ5BvCBQALmeWb6Dm7KLQolU6DEnFv/9sKny
d/7Rna9xl2dhIbtzF4m4wEJ7AgEUlWBrzkLIriKCf0IAs/aYtettoXNiRDv+cUPL
sb6BqjisViEGzomMdLZSHxhgYY0C/VkhrikSDYMt9DVcbdUjVZKhS2qxa0Vln/bS
7tA9aqCX6e9n5TKbf/Cmzkgd9rWhVK679g2EQMh4VAuMpPyXb1J2MEtD0Fkl4qV8
f5WybJYRW1Sosfb2m7N8tqF0Yod4Eo4llMHxaQJtP5cMSyYrTbbkV2GUjI9h9B0u
bIygiYqytlL09YghJFSXDH60Zrvcx5CWOw6cqaN0HXsiHdQtvmT/U3SCUVKtzUEW
gCDxtL1FqglPzj7G/BJvpFn8l1LYN3MLmkdj3B4LXCdlHesXm5XrJwCO9skqGL8/
1sP40ik50HIKbwRrmtg2GsAFsoe8zT18GR7/+VmN1YXpVttOq7D4uoV1jKFoICiF
2M5d4LAzD8LIJM6qHugJDk0pXc6XM1ojBAsoLHlFe/5jVkxVOkbWcbonn+7X/p4A
9gT6tvIWHbIEZFBnaYnaO4RTAAR1GJGpxM4cV3YzhWVD2KZeIeLooVB38pAzEN8k
GPkNEftWoYvDTqDeC+TR/rRmZDwRqgnlXX08sZyCHuMTf/ljRHuK0rwAiFZ0Tq3m
ZM0a5xwtQblJZ3+obbH8nFs6G45bgnZgB3l0o0mn6MyECLFV/w+W6bcb+Q9j+T3D
FeqZOfihv+d5II5JvnHG8YNyhQAgIy7M6rvZ8d6MuYnxd/tWVEPOU1GAywgJ55ev
Jf79ysssKQskXE6Gj3XzDpozv6ja0oAx2F1yeD3yq/wk6OrIr0R+G1GzOTte5GZI
0rrz7DaZ/AlA1JOp84RK3+sup6eKj1nuw+2lNLnVknX/hAZhe4bqsZAYyDEpIyQY
YgOnqJPaaBBJLEzTKHcHJkoreMgI1UtY2hvuuxVCrLwIyI5igpImtq1peHyaX7ly
RT3bahO3e2Oqchi0qB5Kdy4e4Oxw98I4RKjvH1Xa84zBaBSRVCmz8omUdlP/+Nez
C5VsUSuBSOr5o27BGBv4FlrMV2SVBgiRVAhQHgZCBScGojoMAEZ7KeXAKqSeIpkL
PDzeJEMv/dg8cthweYCSYigLVxZGhtMm6xQvoatLfB+gSVdDiW9XVtDtAav/9Ep+
j/g9HKJCCX1h8AXb2b6WHt0+R5K749ukIQwhhUAHCsZmMPNEctGvMQ4Pg9gzfmNw
t++0L6BhMluVkWPOSLYVqUSev34Q6J2geAhGf37TBeCi2BX0zYfNc2AqQHudVJN3
4M2cY+jP0G9gZz60LWsqm7XPGXJQPxBgFnJnWMqEjjZGJaHPs7HFoT/nLfQem+ST
ve6UkE4dqJNHRlJmMwv6al6B21U5fvoO9uwg73IEPh8Z1iF41eAV+JhIirks2INe
idRZSmwduRJBJ6JrhlFaGjeVcXEC0ZqyWrz4paPna6MGrDLWx5R/yrYmw+U5VmWQ
VAlsgP0XN58fDsqWBe//be7kAw2Z1b9GFoL6Pr8RgIe5+1i+/44wC/2Ba8KBDKeC
Q9f75Xv1bisUGQqwvft8To2w/ZTvq2sXro3bnk3DpQLlUSG+6RXlWK86n6NEexAX
FYYLBeQTMFXBQgqi7Gx0lEyPFKb6w8uz/Kvn3pf93vvgKw13E+135sgFPjXFFfHK
0fx3vNH0YpLpMIcT5KCRFKZmK0oq65ec8S3ucaLI8cN4rhwQ8+4/RIHAnVymhwIP
X7ixpj+vqCyJELN+tuWzCU/EHtUGmW/GF/BmVaLstBim2sgvV2YiieLEfPQf1+60
figIiT5k0NdnRHOK4TKdC9JeP2qPvFsycwOJ3bzrNH/1JXeCV4AG7gRa7U0wMLgJ
jCNaOHdfldscJvXeObmDUZyN0O5vehh+I08dwngFLLmBKkNYzQakc6Htlu300u+L
7txIh9yWbMIZx3pxHc0PZLbqZGU1Pmd6D3oeG4Hkdxy+c6Duk94TbRui38uTl/Ha
uDXbSWc+58cndewSQtC5d2XigaYV5Y1E2CUP//Nac8YmK4nJPnCGl5nYIVEZf4mM
+rKFJXzEl7koZAtBAT8zKEYhlS7tK7c1GIu/b/U1a9iwP3Q8K55uwsPZ5UZrEr6s
6ahMhvwC/BGvdMYvVaeZLic6szF0FhcqU9kzt7/cEA8XqUsCF3tBrGx4K1NjXoI+
HKic5uneZRtaLpdA/eQfMD0a37IHNiaU1AhO52N3Fslhfd7zjjWsk0kFG7WQjYes
GMkKaHmnyALLdNWDZ/TTJNH9n/wsLxJDSKsBawvtiw+qmrYdwxVa7H12+qJbnhel
8ktv2m1kAEtPNp8qIQfxDKoeMoHGnKwNUsRkmLEE+AVIpy4uSXi3E8JDlODmg8Cr
nn7wHB5fDvoB8e6/GP4Hm4rsE5yVJ0FZDvtYr2lIdsqZ/3zOzXz6V4Vx/ES9WiO6
oXwSv3Ilt9QhyJIFADL1lunlaOmV6hMME1h5wJOCIab3PCyCH2e6cIKC0xmZkvEC
q0gBzTIZYGrLbYREQ+OLeIwwE98fI7xWotmIrNEaZ96niQlZlGbqWYcM240fMX57
CudMvcXNxxZVvOkJyZ6GSxvR0c4IfX87SYMPyydw8hOikf0/i9XadrZhwDKRuOHQ
Ma8EVKqZFqIdXwck0G8O7GW0Azne0l2Jhvcr6XJ1oNd04IJ6s9jfsMJXEFBWIbb7
51qb3PQ1b6hNMsyMsVS27xv+xmP20HWdl+PQdJYcAjNkkgeV1q/iw2QNzs5a16Vl
iBUJWJtlcmlyIqjP9yYpdgafEb2JWC2LS5eZ4ItOhjnzCf/erBNPSG3/kMZdCR21
plxKWAkUf8uLf2TaMrtnMJpcpGo8SADs3hJnLblzGx7UH+4/SJGdc/atrtinzjom
ITh4feVSj01cmiwTUlDnnjlt48wYmUbKwC0R7DEmShNnqkJ/xlpM91bya/9WQdhg
5NrbVPu1Lz+0xb+aY7UC5iVzZwTMIE3wncvNxh6egWKTgWXxlRlOFek+LxZIM0oI
m/vSanIxyY5qsNwUVo3kG55ej+L5xBbxHIo6LVfcV4aGSsIXbjGv6AHRlb3wgAhG
zMmbLkc5CTm5dDdqJyn9x4a7WhuAU7vw4agJpLb81Qv41hRhscUuruzC2HG72qyS
oFobkvOr4NlWu2Tkvldj2lbIwINSWLewGWWTIgtZr8EE0HuJrsemuIq15q03kNvJ
hCQrzVatO7HCDs0S/y2u0+nloMLpdry10T8Ah7lHqTapORCGllfM/IvRBaV0aoq0
mYKsip4wft0nKAtHIotgsgzp6lpWv4WUT4VOa2tdMWsd8J587ZdVq8JgOrgF925X
5+lAP3duCyaWS+vToAz25VRf8argNSyorEkeEKVR3ncX07/oTab3Hbx2RFwRUGSZ
zb2mW1zaapEiccr+9NeaZi1wh7hPQ0rKXolOEIegNeRtmVX1sJZsRHUNr5ncYwBz
UYiKyLKLgQRK7ofhHJlpy5/P+Ujc9Epq8SFbE+GFXoN87PSzPEKplrlNyFqYNzho
KlUURRLQZxUANpoFdpstjvoId4ox2zYuZyVq4+7nZkxTJ9lbmSulwB6TNsRqdPDq
SckjUQ8AgNScEn2saeevpmWHiuH7tdUP24zV2RWsiTRMeODtfwzLbxx/VVWZRR+L
mCNtx32fvWaqtXOmAymaQKnwEoKRtSZ8slxwyh7+E/pdxi+wPx6j8IdZrLOJ7afB
BVa3022zW7R5sihnK2ocCh/8vcyXL6I9/7OnLwh5DtQtBvUE2YbAMJ2CRYN3Kg76
dZF62Txn51djlBpMRawMbQRZ9aeL2hKKdQ33hpivwJlDuHE7ApTAFmUuB7E6yXxH
E/WWID4ZYXy+mdsPqVlNfkmBabqvKi37MX1JAmmIR5YDui17Vkzsbk6Ga5Gh/s7C
i1XFTdQpNMXoLmmeytFZLXKj3aGZ9rcjFmSiYf8frr2Qwh3IEdIKMYilEsOLJmWr
j533zYBbuoX6t32+wgXZcpDZtIk23ORLVMQHSFU/rYMyp0HxBqahoSAMdnCxcwxt
g28RQIhOiR8A0s9oeMgDNkPttPf77a1AijBanYi8zD1VUk4jz5LTqe1FfhMrxcD0
dpYqShxQAqWiafCDVGE8xhnJxDvkDkyKtJiGY2icumbNma7fg4RqstajE2Ug4ggL
JIrx0K+IV03TN9FjI9DBvvcGA3mdXvND++8LcZC+POf6Iw6DmnF1c+sw5KwW1cVA
IN9cngU1BNvjaeJgozpSbaacSXA4ncKp6ET5XRkkhRu+vfDw4/8bh67be8DfcZOs
UAYzh73mW43Z/vgxUmYTeg34VIgypBOj0EH79mRfedy3WeorHSt9FMyfFDEG2be6
hrAEOa2umrK9kum6dHhwpZbtsh88VNEA7kTGesmihZTDandaxeEw2AoUA7AJ8w2g
0iBCGHeH1lBRJTswCXnCYhKygL+vBN2gWXjcMZJY5JTqMrgHUooek6TVQT0Y2DuY
zdgK78yEROVzEsIsb0R3S/3n+WRW38L2HBc0pTooLKWj+Ne3dYCzQiixldencxp3
ieCagZedD7JUG7VC2VsGBmbq6DV/6y5jMiOxiPNvGBEOTxfGGkj+FfjyXb9JR3GA
qFrObDVAkN97V/yXTYMUgH4BJBancnnReHMQfDfgUM8LifyshM/fdGdYPf7BSxWU
+r4Klgtlx23Wlqo7t0RQ3YOfA69aociLgHEHg1AVdZIYPl7nyedX7oUOXFCrrIrm
O0jQG7oMIU+KYh8kX4H0L75lH5+SwVGQeIUdvJbMp9UhlldlQtwsToY/bGBpOOoG
IFEOxvfcIIUNTLR8qIWfFThI7ZpfyXBrKPRcD3uijnY37nlSvIqewZnVL3jb8oDz
1NNoAq3MMNZh6DKLgmWSa6c8HvagdnyQELe+0WVDX5Zh/UKeEHcsXvPS06iFaWe8
2cCS5Dz7LiFQxTta6A++DSSoR+jcYldRcWyqjuScdXh+VDvibacKsKHBItqy65GM
+9+tU0xlqApBxxkI9QmayYEig7KvIkXaV42IOJql9wqP99EXIJiGYc2YIRHklOW3
womZRixoCzd4tfm7FEhgTeQ57qmZWx8IZ3axfk0uGaenKJlmy89kN/CXHBGUobvO
IB+QElttpRk0a8z1cM2PpCxeU3FS9hwRiBnqtIF3dm3pBjLWu7p/HnHfWabBcg1F
wPvuiMOxLMSdlOTJvrqqgchKdtsSHNhrtRZnjggtsxGyFJt9mKAE4bfP+FDTZsFc
jdCv0ni6OGELY442m91EAmLysKGoFqNhaPAsaJkJT+ew346XeT86M21iTFm7VnQj
GDklxl+xYpvSLfSZDWoobmk5tnPx3sWyP8prfRYjdBYB85XpFpGrJfdoXEqS+hJ1
ICU4y8fbKCqWghM86Pc3O15bmd9dTKaDh2JUCV4UWX/1P1pWpzvwCj8yIKau9fLo
/3XEGUgpqjFZXsXnMWGpqZohsCo8VpIn4fV1AIn+JPNkn9aa34MNRcu6TDHp7E0n
D+zSj783Vyz8O98QXvtYIUT6i0qih4VRlDQDbANakI/hPfGensOCTqB5vlhKQntV
mU5vZN9r6B7U7H7KgVdndf90JKgy5TE37vnbXd7xnMTlWZFI/Uz6QFFNQgipXWxQ
N9iZyZnjTE2K1xvSat2Vq5iWflgffd9yRc/ZDOkTe30DmXpX605VA9clGrtq9JnF
3QFmzbHwToZodBQl/lGMl1aMfKTWPF94NdfT+7vJDUeMWuOQ3VPHDgzzJO/QMhp7
9f3nnbzS8H5XVG2r79mZuKuloLmIZSX1j3xJwVCy9YNCai1u16kV9HlWHoPEN3Wu
9EjD5OASMGWcVZA3fQ1hv8aWItMLKDxPmjB1AyZXjTy97gbYMMF/Bj9avndVvLeD
jpYtJMzu/acBXzyD3XZ+FGCz5l94c9SIsUNyrOF6cXix7+QqIFuVbRFH1UNAmeko
RRniR7FQbL1uSTJJ26TeO2R87AX1bHfhe0L8Jsp02iwBCLM5herFPloozHVrS7ol
gvSL6EtC2gAX5xN3XCddd1ygr7K0wtQvOggdap2c3GEkngyYEUvVyBWimytYAqVJ
J01Z/vYjrQN4BXvGqFcVY3s50ZfIW49bpQ68+INQKXFWsdgPYDgjk98gtyWVQsjM
uTYyt4Z9BjvRFUogPMTJSm6Ava5ifcO5zJanakPiUA0FGUkgiTHM2dTapRnl61dW
ZV6ZTqHcr8z4M56KG4UPpheSg9aXbFJ2taSnvUVfP2tmq4v42mkm5sev02plYpDF
B+ZNePz99mUEM3Rz+h+tbebOjEmaZLQJg3LRt/ZZotwntNteGae8Qti6VPSEGJOT
EA5gg0XOuQqxhksZDL5+tat6SAF6c7iNng0yKF7+DxjMXbPpY0Maf7l0Tcqq46MH
CZCGAHwzrZVkhgvGJRuNEg9YgJsc6MMsoymHqpCFkecESW9ayVVsKTAZeMm01QDm
T4segZE4VTauELznSGnMe+KjveCn1M1FgVS24VbB+cc8/DADMh4B6d5X4GnQn8Fo
rykDha8DpAiyffmqNm6u9bUZjsDp7Iep0cdrPYZWJrzQRsH2jnCa6seoku85hri5
JPT4E9deReS76PZtkso2JKQI+Z1wQmI2QrYH0Is4omTsjeE9V84ziGJRPXnyGGk5
uPbobbYy5t3CPISo6pH2790dkWm/et66Jl2hilLJ7G33DzqSalW3tVZW6kw2oSX1
8NKwNVea6EGIfc84TdnXqd9kTUB+splE2o4Y5BlZ2aZ1Z43t0WViRFbu7iA0rbKf
IR8ws3qI1DRnhCEKU+ZMVzJj7fqMeU0mYcj32N2b5b9RuZjyX2HTnHuMTY6NCzj9
TH4MjWj7H/wbOBw2qdfgyxH8z0ioh258NDxAKyhO9C2I5WSTbUasXI/+kyunlwee
T6p+nlZ7pC3QCPjcWCnO5EtaNDCkMCGAJZT3xrSQXZMSDeHhaifQdsuOa/goORMC
ai8UAovnJuwtZTIcl24k2NF3cSyJhjmsNclvF6clSc6mXPm660o2NV9VpRtCZfBe
YBlDXg+GIHD+w/mHnOtJFzEG5Qa0d5XrXNNwTZsh/ftHjA7lUBZp6hDHw3lq1zHM
Nv7uTUI79bCvWzyPoub5UtSeBsf3IxFwoIO2ZLy+Mtnwm7o77NprjmMZJy//qm7O
VR3BiG1KIMynopWyy7haTMZZvH3zFwM+7TEF5EqL01VFUdoq6O/KLvCU95p3h7hF
UvpcZLJfziIAVdgfA6FmH5PdG8hbdUy4yZXd6viz1E0UrzF22ua+nH4TSJkieMqH
DacIWyc57SeO2n7tXmr7oFNM9HkDAMU1YMnXxthnE5aLG2nW05EDNrlAacTbDnYF
J2CeM88Mk2F8WzGrfjNPstgwUUfanP3TSQ/FqXaVz+DeEPQbNquayriWPOS6IcGX
BISvxFNHl4AQovjgBPyo8CsvhchmSDeOoH8wjMlvfqzLj8xh2y+WJdAqFjIJZCjA
DHuocPnhG9umPlH7bP/2nbqB124neiamSqYKe23jrB8bjTJaVNll+fyLGRE5FO6Y
QW0J07nQ1zRhMGmH/8CPeoOIhtfL2d1q5Veb4N3RLq+xIPlNEi1IWDDi9BVnhADp
x2c5cjqomXtCAs+2HjD1jmWSOhoaT+YlhOLZw+z5lNZ17DWzMEYY/60nQiPNamff
oDRo+q2OFXknlZGGKhChf4s0aWDRzdG5QFa6wPdli0l1VXfVZDIYFrQpdH6P+RX9
vYg00VjA7Q8ytEvxOdgGvvVIAbsLSKfTa7v2bH3uM6CfQFjfeG5TiWiF3S3TI/jI
sp8EDpjng1rZUsETLFXtXOcJtrwB6ow2jAcmLIC6x5ZvFJC/jSnp73h9NlPiJ/zf
Uf8Ht0fll0xy4hyMFrWbXERkQl++pU6siHZvTIzSSdAp001XoBCYmEJQVFbPwYli
9RtASrRrwmiH4oP+p8G1PEGb1cX8sX74cIel1K2anFI2oeCkL1ZQgHMfAJguosIv
3QNhSQAEgwVwyZJXCp0P1LA0f93Ljl2ogOsg3he2WU+JGEosdK8X8gOmx9OkuvI1
aBBjrfTsJiEPF47jxw8w/oxC+iTiMp+IyNFk/JK9uoELT7b2HJATM4KzRb6zlrQw
bGWCwMDi/j0/xIgyMYoA0ZGe2caZyKAEVozbfJnb2kXOZpb4EgK/Fktl49Xz9vBS
UtNl+5SPXFj5NTtoQQ4DvwZIXk7WNfwDKT+iiVrA1FF/TFXcEM1EaG4eb08u8fpj
VN8g/XczPdceGHDvV2pp0dR61AEkIQrfszPWqB/OA+BlpQMC6KnLbxReIOdRdRpL
ejTxpqas4sWAH4u6FSLu18BOERqeJSyf4ufLwU2/tm+eidR7KcyJZLmqWMnaqPAE
518K1mI2GzIJso9LaiSrAhC/CXLWmouxQGSDlnHQ6w/vHaMOo6U356Bdts+wJf5D
docjvNs3UrclbkqRLpCSdAyU1wRfrkulu4qp2HQCrA3UisbO/x5g86qgYPQx2V3d
czunQssu8PRiA67z3gUcLJWwkKCuftX8DKOxtEUqpDtFBrmOQLcbisbX4hVVPMMB
iXgWLT7Gt8Szs2+LlmFQ05bxgjDrJmadDPdjKa/UxNuh6lxS9LNA3xJKlK9QG4aU
+X7FMu57Qvh86bo9dPHpnF+MlrA5PZctb6Bl7MIyyEGFvdZ3InDCOX8oaMxhKxnG
2PBVFE4Qu5jjmGcNcNrS0nFvpuTN4j+p9J7FmGJWwi8O8Wx8fqFVShgCyB4P8bxe
R6Bi9KwcxruzrpY/bUwOpPbMlDnvyWtbV84DQNceLHpI4TtWzLKlF66POt42fN48
r2fPHTq7oQYonjzpVLiFNmtJzfTvc24VsjqCZ1DCPryNrPwpEQnaq3k1cyQcsc5/
aiuAqCyy4ekrVmIHjI8xcgtQt7lwi3d+mc57lxzbINdY9YkbPTPcNZRMHJ0t+G4Q
FiLEr5tu5BsNi3/WKi4ikae0aCkoOmZgTxeErhLmqUAWcMS4ErJLwthFp3MpPUyo
5jMtPNHBGAULley3JSonGi6RPs42Ido7nrwkFkZ1JP1lNrX+D2KEj9p6HnVdEWhK
DnmddpSDjO2ysio4Li4VmDlkFuqZ1jSTkfuNJyqmCe8WUkJKSBbGoeooHego7jL9
+CYLccFLa6rridJ2m9WKH2cMsvafP5+HqEy8fkSv+Cacpe0yY2cEJGpACtCTxPX9
cEvoHUNF0+HkDqb5odnnayAGwqf9+7krfZyScFRnKlZ+AtVoQlQCNA7tXQIKRJvB
rTMFYPwatdcQMgZCWmOfqwSH+73Rnp52QwbrEnocy0ORg7BHYEGYhbNW67QCqJB8
V0glwhNgmheeZSBz/H2ELZCne0JIYWcXG4sRycq2d5IugkWlc6bsz7jzAkkhDzVX
JfggB1jBhnlSiXj29Ek41PzIQjCbL8MHbuigLwr1FukyomIzVC0LGU8/4JPWSWNQ
yOvkwxmCh7vTMB8MkzHTEechjXojX/1HcifcD0x4PYsdhjYLn193IzrlADi5h41I
qmF5GsLsnHJeqwfr1kXeLXKohxtkejDjbcLkkZpEvYwKulWa+UH8a6oGghXeGY4y
z7sge+ZRPtZOHmprFeC6bv+Nt/apMmXccc5zqOoKr2O1LySYhHF1NQyC6U8ezK79
wrRl90NwKi4Z05bXEy07IPwgvnEM86Xjms78BN+GrkkXdCYzgsn2LsQFtiBq/aof
X2Bp0u5YxD3ywFIc1m3ifAGnMIm4WEVDGbO+eISdU7VceD9yaV1NCP4xEXDmUrQQ
u5bZukCWaldYf/AJfBO1tIlanbfj9gqRD24zoHdFyN0R/4ZdKUMJClcwddihuEVO
YNrRK2Z3w562TZsNywD9smT6rNRg340hWCMkWoZoJVyqPML5U5S/oWVBKlLD9Ygl
L4kZgon0hjjVMww/ztOeBwf+Zv6MD02/xSZVMi5RJgrQIa6vSB6jKoEdXAU7d8sz
Xwkg6RBGJNscFNLpyYAlFkeswr+Z2eskWl82BFAcQKD6ioJ5lNV7ZNJPMCZgxRLI
MrDxqlE7cipyVmCEFLZGOCDGtrk/CKusN6Zm0IJ2yMPJgTuOyf2ykWJBcpF96LJ/
qcItFtiHaXv8YrIw/nHlOXfMnM6p7Vij4aTcICt0Q5u00EMW4piR3JEQ95c2OZwp
On7C0i54a406IxNUXh22fxdmigacDGaaA4y7UTSCRcQ6HgfUcxqZkk3M48MylhOG
zxHto8JZeI9axiAMAkav+80yrKH66zI5vehgT6LFw72RdDGNuHlCA3b1bw2AfPzE
2v9SlSv5j/g56c3AkHJ/8+/TRsJoC4Z80vrUIcoOMUr5VyoDG1zw4U6Wy3Vw6dZK
eWXIh76Piba2A52zVSNgNyBgQdhqmVX3kKyJNTwEwISAJKoOZLWC2ad9/klwC168
kEQLXlaAVKKdBDYr0Kw6aOV7/8ytwGGhSkogNEncriN2VQwXHrtWofRCjm9k6dzJ
SXMohHcFU7YdgXrbbeT5tdAxKix2gpc3yLLPgwpw5KDBv69botDi4385rtck04IN
IN8+M2bdYmYK9st78LFoJPXZdYaGzVnXRpL20m/eHReNlZQIbEiaJs3TNjRwmMk5
RNu31+GyWrG5pwECdSaT1rk8FEpcXexJUscqPivbaP0h/fmAhrSoxHCS74Li2cTW
DvNZYg1Nk9Bbnt4Hh/P/9c9sHwt0DEVxOhQadXvXW+GOy3w//G+WJ0J9EKJ2DV99
O02fhaeu8i9tsmpGYm1dN4sN42WgLdI4joLejh7t8h+b3k3y6wJ7AW3A226vS8M3
74q+w3F8WV2lhcAmPEyYQz2Vp8Wu7IvW0RMV47VViXJlbqmCoZLps6MeUG3L3Qax
Xmf01Q09L6x94N72oHdqTV6gKkRGTXfFEIYVIFItkmUUWKnwMqMO0xgAi79+JRzU
aPo+N4TwmF+YvXzQb6Xc+meGnaiU4kUdFRuv2BkPwpRQKpPEfCMK6b08iJTgqH84
paSDYh8kqHPUvkPNvKQ/7QorO+xrIE1xfief/pn8fus08SlSkDvcfxLnMusPTNJ9
+U3OJATcGhfSo7C/b57B1Wfp78hEmF7Xcb3eTQKbYgUdRDdBFWW8ya/CwOomkwyG
mPzxMTRYySj1YPORkwsMwY7HG9R/46WM8kRt77g369rW8TLYS1duT8skciLiRdAh
aHPmGjjqKSZltVsZsIa5HAgWaZTdAJuKIP5gYI7EoUAcwlTqmIDeCqTj9LUlsTqw
GLEhx7QbRKv4GaEPUfoQYvotH7wVH3tOO4lLrVnEDiWolx6B+vbQWRtbxYwiv+US
1qMVY9wblrBRXOZ6usgxwLXRNkc4C27UhdbtI6P4YdwkQkd8uNzeF8uRrQEPWiol
KySVS3kBWgCJCT7s1Z4dBgou/jXQj0Shtcd+OnTXpESOMCU4Eo6kK8yEmMwy1CE1
VcnPUmwoR2hYNnlcXMN9j7LVkgHCjNQwlOtEuMOAXekNsQ/nwmEcZeZj/tPqnxlp
BE1p0/rIYSbX5fZAnKMO7Xr+uVh6XtelnuwPOSB6LHUflCmIPoTlNjbCL0fdRplS
90KkbhChiFLLCWClaKAzTBuyFclngfimaX+pdzDLSC5oBxsR0U8tVuAbk6FpGTPG
CdAIaMwwgyT+5HapuQItC2goD1dsXwumly3XEC093fMWdIJxw/5G6eOd/Hh01OTu
i6pcXgr2kjhGP1L76UhLotVkn7qrT6zhdW5FEvoViAtZEScKomwauQAXv/RfwGEG
m9QDIelfioTqGFfo531mmlgZdI5DKhd+wtKLBoJQZlimDYvfVCJ1+7A6aTPabnmJ
GIw53mjJMGhqTiB8rmcw7hLSIbty0n+KSIe5Zk1tWfacSAn2SBg2li9tDaqtiiqr
AZhgaweOdaqP5xWRZB4awqaeIm6QTV49inxLz7vG6ZDCoAgsN8eYMddlbbR0RFpx
ryB005//V6ayxhs0Jqdtz9Td/i+kXuJy71s4K7JW8uM2FUYlBpX/YWBgS8EG/nny
Mq6UIG9MCKuUygh2XVee+ll1z6/Qta1R+1F9EhDcuCxOmiIm86FaLbx4dGHnv28l
CFKgBgfqh7JDo96tfpKo4GAh6jPGXu1Ebw6NvRN3xUQAa1b+iIGhtz9iPOUIVUaV
q8OA5M5cd/jvqc52v7U91Ywpi2mT6fHLIudB9YN7dou/CVp5kEVRBmEDDwtgMaM+
e+XxMTdBx76ehrC7rLAVBZq83W0E4T9nv8bIFCohh8WA2lNwaSddTBVW4WL5sSkk
1DPXrcJRy7DqE3YbSNrFFsott6MEhGlluNsqnmhLu3tV69a/Ve7LYwFS5Gf7xmMn
RDYwKrwYBvu46XFHN8i60oxd2RI4tYCjGXhalPS+1sAzF8C65CCajRNEpolDYamW
bRTAjiB8QsnUCbPnGHACacf+HUswby/V52rvbweCpKcvCbSqmS4Wa+m9o5JHijZR
ekdsrKYZHq1y9IpfTuDXPB7DQwQFLhJyO+FrBWxqnn00Ie+2DhojxNF7378JbSGD
lfYttzU19qvJ/XVlJfbE6mHivlzJeFGbfjpEb0ahYwI5v+tCzE6FGvnhWZ8L9nBB
kgacVemhJNhh9oWrf/+Vy48aaI253znR0HJxzi8HhKN3rX4n1qPpsXxdfLRrGFQk
MmF4Of/7lA7VOr2aO3TO771GgIWKFWvtQiC1H5zT059M7sEIgWNRvu8JuaeEV4oo
bEw/QtmMnqo1z4/6tqofr+oE6nmye7i0euYQK+AYcs2fyM+n58RYfJ/V3BKCllTO
HbTgsL08iyma/xnKn6Gkc+nGt7TSbiDRh+2pIoOL50uB/ycwcBFPtmfzhvGLVLsF
lhkNsv1R9ti8iqojTOGgc7ppucFLNz8mbqdg2vec2joEN88m50qgWqA2zxyJW08a
nlJ9PeksSbbvJ8+mgY7HT+ex+qFPY1hB9L5WqJgWdxL6ryEyO+ojhlGo8DcQtLG2
EXR5miyoQOnnY5WhLokbK9yWbspSbt6E8ngwCsm+iqcxUiM9J0p+EwaJRLNjeAZR
LgdKBbzbXkByx8FkxP1tujnlaPrOh2fsOgtoZUyuZdLDm5MTpHM5OnlgQ1htyRuK
V6srpbvDgqmkT9AJifbkmx7BlnUjbfBykG7MBgk+igwaW+7JvyyNvArq6BoZ3wN1
jvclwNf+G+xbIEhYzcwBYVamwgLBmP9yULD574eu3sJaAWXP2DBkZWyK9KxvoMXL
dOSmvtMpz1hRmvdR76HHOy+NLlMV+op9vViZCOuqL7x88SYTX1gGPTNKslJv22Uv
2eIFKmCWZ3N4v1EJaSePUo/yno+GaxqE9srH8JWxHXTBvRNX2PeLex7pO1vHggGk
yW3UKstmP5a0ShA8gjom+FOluZsmkEP8ghHR46QSD9zEPN3syC7sRTF/rNUcxog1
s7A35wTAensGTfkaBYDP66l6Xt60PDMwqxcXgc8Wvmi3Em1IjadQk1cHdqZWvt93
8+DhpDUN+iHaIpYCOYncMrgoYW0j8eUDp+1mGQN1RduReMj+Ki+JejjRKIYrFEzD
Wh9jinnlTh9OaVWWiUHYCT/vOWFl/PNFru+IXJel8mKV8PNvAVAeZsHoewkm8jXa
37ZQ79Cey6IfOyQiudO8DwmueJPjgxA/dWTJhYosATOsTGoDLiQprwuOnupk0MGB
vb2tw2+Mh7LANexgSkhbczx6AKvWYPVJbCitWfQtO0a9C6cHBWpNvTVvTYHk6D/i
ZEBJFYneLOndTtE/9XlWkb8j0RH+C/SlAm3Oe0CnYOZqkcIV476tzub8eVwuU75/
5dmCyFC5avZxehipAIiO6qC/wFXD3VwWm3s1TtWPxAtLHDbaJl3LgFsCPgXpc6LF
RCnVfB5hen+TYtIxLN7GBp8cOFX+b+C6GCUHkeEp2mUDDxN36gbgdyj0oquQW6tY
VRhiiJwWXLQgFUXVd4Y0vQsH6udKo/ReSe4sLda1ZDCZ+CMDQQjmtk6oHWOASu3/
3nTiDNgRoAriRVOvIDRvTGPmR8QLKEQbkVqLIIo2KEuCmxJWW5aIPUUIqtP+LWdZ
f3Znoe0ijmb38bx3r5Fk9YePcsg1ggK75HMD153stFhCyNsIgdgXwPBfGYbs8y6D
jw/50YBFk/moqfwGlTYQpH4QyCfG5V+XY96VFKlbjBcMg2aVPfXvqRDOwISGF5rg
gUn18oXI49JX4gwvyT7OJ3Qf+Gfw7GGMmVUUWdJ9bDDoSIMnEjAsqAHQrPFhYBR0
SHWOdYOinc5VtoxMlmmM3blyLd5adq6T4u5WSp73Da8twjVbqH3QXtfNGfOuKUIv
Ov4bvmsWUzKTqyl+Jx4p0wd8bQVZrQxqyCQL2Mhn1XzfuoYKzJ7m+M02UPV4YTMB
TE1NVNcWgBiEuyL4LzIwlHGc0Go7C663e1BlwgMjudO0x78/ZHJpx8lj390xMBpw
H5E19eAwB90O2v+yPiNd7B4q95hOb7kyJyKMRq6UkVUrvEEJ9fxKu9kfbevWO4Td
c5csmIn6wWNEcRTlRhbX/AlMhjrcPX0jd7UnLMmTQgZQySG4ajxi0Akd3fPGYKOd
JVfJeCSCMChyakqXB7H3P0CfxEC3SNXbgnJGliiub0i0DsB8JmUHUGBmUcGKCL56
fl3FOARxw5AME8RWbZxIyezSAolUjtfE57DQF8iLs5HWX2i6wFi9qnvD2i9Z/06k
EcD5V8Y6IqRg62aH8On0dFAcVKeGt3T0ymHw2DwkWH+DiUaW5hsyN03t3NZuX/vc
x2Apb1Qpm9pVzF8GVNHVdwdDiRSFXElq5WhLzKVDpmG2fNs/Xlb1eYRzgbCP7NYV
kXnkU4lmre8AHcUlgFG+tnYxbwX/fXGHy3zU2SNB5DZC+wE4EwKfOPSeoBoh3vf9
mrwwJ4wkehQZFS/ADhJ3hKggSWcFaCEuyX52UHRJAASIpGme+jAhgHKvnUJdKRL5
XOUhwY/m+g1kTIMIMUh/ykbKea2KcKx/MzG87VppDiZASf+aSJkZHctKQaBr/gAJ
RFrmRTmyYp7M7L8CLIToigBKez0Pub6cWAc9nTfZaVbs4MVvFBrjR1RY8WMUzFNC
BxRY2eHDRwpjm5DBt1b76eAhxe04O4BzjWLobmAMRYGT5oy22G/muT0WpBcuURp3
uyqF2ai17wAgA12xbgRcviTw/pS6IgAEk6AWUJQUZgpJFeFEOV6XWAROhh1IDjcg
DGoO1zLVybtyfLmtcgwyxHHVJ4u4lgXyiMK++vSv2HF4noZK4R20/XEI1B64cFTh
s/VK3qsBuXLWMagcfYFmf55cjhKgU34Cd1TrnGJx+U+rviO5UhLGF/bcmI8K4H45
dM6aLb+wQO1596GHjJnUbgp/gTdEglsZXiUJQktAFKJOhI7qU0rMNaV26tra9vyj
j9rfYRyq2aNNJG0KVeKXuo8iZOEtk1UBuXes+FAvNVy5yw+UxrV61FCUJuGdHNg6
kiwcoSezGHKYtyai9MzpnKTUEf/3UI21ImYiou2tbbQJHDTa1G8ITF7DEWGbAKVZ
s6aR/RVSkRkCd9cxTGhyR88yV9FCTxMcnRnPWFLcqv/xb49z2OZZE8zXAc5FbIvh
4Ty9VavrpbTyxlJkDKuF21EtzgoZDLeuloBlaaQgO/RhscgMEiRwhY6l/MuY69qJ
v07o3aCe+NSI3XcTCxBXaWkXRMRQb+EpuoATvSlXBs2jhkYDeodV/C2r+YhxLYem
wBADLE2k3b04jFOe6sWjKIuic8dguhqKvqWMKGyHfftbWCTJAzuf21fP4+6PvmMv
+c1ejVwKdHL1jQz2j+vNLbF7be8hZgHah8wIsNz6qP/iYAmcTB/4jZa3KL4KRV14
/fHVdloeLaXIcWwhDIAls8IADjx6qApz++CtYVynHzBFHYfNCK2fzmcargb2lQ3n
YK7Fusf1Py9eGUwxRsAsh0dVc7Bcvllr56C9lezMFk/u77X8h6D8sNuBaMyaS45B
+StMU3ea5fLz3wJ4u/V8tcoJJS9O8p4+0hkoi73XjaVPSZfPHq5ybtnINaRoXg7w
2MXgermBUUqwTNMmR41VuF9xrbTiUlRPlLspLPzhwFq3T+NEeIgKh9BuGWDB2dF1
a06Iu0jKxo7D/cLzE83zZI2+zoG+noUeH9bTyswSMiNyqZSv3lcIWOJOurIMg4KT
H2aGwW3zRXdcDwdcRa5x9R021VUiaTgYeb2Nekt2tC1fQzEF9vFs9ptVILVFssDN
UNX+9aDtbd6Yxed86iEJk1+QVVdMODShEiFqnBocJpokzvAdUZTa+IKIpfV4iAlw
McX61AVTSvXwDj8FgtljBWlACigOzpDSFvakXyM60DhVTjDFtRcDjFBCXYdgr2Sk
Ia39E8x71IhiZ7z7NTEvaKxusFvqiLdYLE8edCdBTJKniRDcq6vYEVG+zZfyoOsY
j+29wYk7gQFfIAkagKiZJ5BwHyZQmBysDC0ZIubEbcTHYQeq6XdLR+WYQwOhK1Bb
mJt/6XUzSeQLuc7xqqffF8vfFbGNJ95UisRtAhCbfad61O7VvuOx6HZAm/tc7peI
SELaU+ziwHN8yJ7+ykYm4Rf0OPbfnd/9916Jsi/47/R1Xdgo3koAGSrbThyDMrNb
3uZYkZM3A8tBW1OKlsjx9UEEgC1lV+UQsu82vdKf6I84JPDShSmnmvRbZmAAqQ3q
BwQsqkk6+htyDINOGfukqVepUNNQRX/xF6Ju1+fsdj/g/IcW1VacFZEqsFwzzPiU
J9onLr16m7zudnzAU7U4+7TRZQ/eKPXo10fjJilhfuzFctq4L/Q7m8Lxs77F0GcA
d4NtPa1atODInuF9Wyl1O7XDz83AiYHaWw8jpD3Wgf78011Yggtd4O8pRqNXC5kH
KzfRaIIvwdGMh+Ftb0LvWZrOWfjhjU6GW9GLpm4yyvlY6+o7Qw78Av4hQHNJVEMh
kAacrXpazkSXzOFUYG3bEF6IQT0vQ46WYN+RrNH1VhfofSwaBFRf0ixRs5aBtL22
jQezRFqxnefrYjC1K+UUKexQMbyZ0HIUXxL8CVies9JJDxnG0X2AYmRIjibZ/GrJ
o1KQ8IQvPSLb4xlGaFkDdj1l5UWV+yN1bqFvO6Bv8gzlUA/6XZ/uG3YG05I25Q+r
TiMn25T8/1MGl+nJ+hlMMU00ws/IvOheUH9aYjhvbNKjciLSoXakzTmsNaib2yP6
ONUxcaF4R8Tl4wXDtH/DDylL1Des64n6YPVTfDZur6JSIPPbdbYXxDrAVU6dZoZB
l18knAzYTkDwYniT7S4AIRmKHTyyw2lpqItLspP299ZfdKbdDV/GlvZ7XRmWDSdX
o/XOeUralWrT2MTAhzhgZJSQ8/Sl8UtX/8AnNs2Jg+quN64JtBzQOr4vfGlMPETh
WsiCc+GMCa5CVfd8NlgatVnGqBTSdBkEKYvAow12mtp07xLl8zTvEAVsgJ1WDiqi
11B+Iy9ZScy2jPqXJ97pu1nTy3teZ2WCKhIus8irCfCHoDvv3AhfWyI8CuDBk7dD
o99IJ1dVVHrsfNML60BrBntqz5hz4ROjNLtWVw3119dOwkVtEsLx2I7v6VDT8/LD
6cPNdK3uMd46pcrw6PGqh8rPLiy89xNXcGIuZIi7a4bOx5KpiZN9EZqzq22V+XkO
8PQkcE13M/zOOjWrtGwiMEv/hZAbQZBbo6KZTdSzXTLo+pPTl1tkhAyYg/ltPq9K
XNjWMdVAVGoti35bqjUMb8lXGw8hS+DHV0+rvIlpgWDco/YnWkTOIW5DiUFNKa8e
hdTQmgH+tT6/Orm+M0tiv5p3x7/bJBrjC5XcMXaSE6mDlPM43OPkxWo/aYpy9zPr
9Ha2Y+5rTq13vZOKgQxxxbVT5bAdEBqtPk9X1EpcLzpDSH9DIwM3SKM4oXizoI+n
ikQQpmM9fPbM95N/o1jAi48BfkVC7wE2zjNqKFZNHpXlAs1lJruAzsSJqyliWUvf
coR+0iVqDr8UZOBgLU2FCs7iV3a9sI+BvbcnEwu8iG/C1Bn/lBi4fv/diIo1XjkT
+/qRGnmGzluvhvbjVxWbshn9BbscQYDV3rTAD5+/bW0XVrArsv1JM6tCC65DsyUJ
BMwLSRol9K0p36c9Yio349w+qf4gCRz4YSFnr2rSViaqiRkZP9PhonZXWWFoUqDC
0I8aT/yTLZzniP27Zg9+TtAx8Nly1ziGrMyYvTpG+IHZD8+8tbnaNtHyw1TeCBIF
2OQRX37Ob8TTVzyWNCttWgyqTIk2dBsF8CEFKFhfUWJ+EUvBr8QydDgKvP4lKi/c
jpPNjyOylD7uiH2PT+5QYBz3sUHazIEdVIH2mxTcT3XdTXMLhhAICSP+JTv7GhRy
4bF7N8+tvJ5iTZUfTxeQSoJAUJLxIVW4hL43cxpylAsfJbCi+H2BI0FmIjFvGLwm
HMDKD9DBt41nq2pBojyZNhDu4hKsG4uG1yBgqsG18ujEvGtpLHsk2qUrc09Aw6fv
/umGeVV1dEn/IgvqCcbH4TG3eq8PxbyNIArTizIXZecQfnrs5pMGKGYzTZSwnH3Y
RPU21QDodfWxP90K0TnA9/8xmw56sqz1k5fy5bDBcHudb+MfPpjpQuvg46kvzYs1
i6q3YffqoDIV+m5EW2vxllQdIgzxoU9To2+jPfYe3OqvEhap7VOn2OXVRtkG35nw
7jqXTI+QLyF2sMpJMdC6CwVrtirDRtef2wFiZaFuvf4NjpHmLXlGj/BSa8tCOGzB
4XKbbfRiBjlxBVAoF5iT02Cfym5xCyZBHA6EhAM2/9UBN0HbMLtT0bjhnC0eBvwE
CRJzqZcj3aPwBfVCcjKfKlu44EHDID1D0Y2mvxjoyMgSRF5it63kUSpjJLQMKtoY
pHmiOuZ+zTgzYfah+bnP9Plnme8BdaA8HnrIwCDP42kRQaePR8aEBxjmXN+9YgVB
JG0hMMJXhB0G8FcbMoH979D9fU3dohc2OsUim45Yq0PDGf95sWXshdlJoIb8Vo/p
Df0E2zm2ZQLFjpVnKlu8qJICYzh0prQ6KclFPFtnpDYhi1dWjg54oK7+DO+nLWA8
K+tavuKgjAdNC4MXEdR0S9kYiKdQOQdLMI8mQ6T3yMyS1VGKME+IROVtVT/Sd5Ml
zVLOb/oGqNMUcgEa+P5IGjWiR79vf7NUknOdvJqu/JnR6NX/O8kZIii3lg3aOQe1
n+4e5ChmLFA4PO6Iyyi+8iNduT78ZlbfFcepp0Cg8Etaw9T2ESWgf38vN9dVfB8n
gmPYLD69bmadIF5BJSCs7NTDyKJ78/bErpcxMKWAsbJJ1nSR4Ba4T046AnWF6sqv
//MJxFbEgB4qbk6jDpe8ho1V4oGEmZTh0/27J6RHJ7AcbFODxcFDm5Zr/heXlVQi
ePsL72unOyN8RNP1wt5V7UzYlaZsNwUk9XJR1SK96icNIkamFjT+Vj7SiuoEpp6K
NgRzo8EdGimZPemE+I5RVg9ONtqgNEF791NsYa6YTY1mw4LCdfe7+oF73kvnHXIc
enl/NnMpjslAwrNeR2mj3wwzb3bLBkNSetJvKf+TaspSxi961N4VHGc0iLCLxnSu
8jsVF8T3c9J6PcfRbA0iG0PR+8PCH8swpZzRufvrufm0KbxAhnvAArgJDj0hhVs3
T+HMjpUWrjChqwh36NFslBUR6za7VsHgNwTGVDH3l1CKr0ID4sx+gG1oJV54stL3
kc7sg4ZqhiIOPD69SyeHiHFNV3fSjuQyOV0/q6Prv2xR8TPxeWqT01qxOdfRZNZu
Wa90lrmcVClIBc5j9lOj+8qSKpYFFIKlUtOLjmElNxi5ZkpqGzeFAOSmVRinyYha
/k5Zz/O2W9dRE4olGlxlUdR1kTGp+9CHRWhUMfZIMNhVsreDaA77va+Kb7xfRiDH
ov3+3FaMODYlv1SviuQoc7/zTuRc8GnaAHHNnJYcA6lWqOBw16RE52DkL0Ftt74m
0ygphY2+i6NM3TbrSsyGPewADp/HiFqdYrWCd4Ixre56lJ8FFrJ/68ieUArXgd2O
UKcZPVQSe9EsgNxqZ0QFSE/fLGgYXRwyuTnmDPIoSKTM0vqno+jEB4XAEgHrtm6o
5IsK007PyJEJeJeE6SZWFno4SBZ6FyTfleBfermh9G8n9hItR2Qla4CmirUwIz8S
Re8zyBAPG5GAiQfFwNlMIVYk1rvYVsANhxWYRqEM10CQXiQ2LYEWv6NnWU/q5XUN
y5UOCuIbgMVY+wvJ3NUL/BvE8UH55jjxJqXcx78zxlnAOfuLSFay4akqudzPZJre
cF8B+iqdNqA7npS4Qb8KA4NBcu3GqBk7lrFV9uz+SEQ3DhFVbj8xvHwggaTqOhDO
sCS5jFbopDaQRp2sBLrGBCsKJvQy/wVutaDOw/v+xzuQR2rBpEq0BWlq6yuVbwKx
Jvr/ORxuT7JIZITlVQHMB9kzUYv31QPwaUAkVwHKhk/yuxWHmc6C3QDN/VShQC0L
Aa/gUdN56R3vmJvIb2XIy1EUPIHuDM8Hw5sdpCOq+DcjXib+H+zVDBxD0Gl5y7u5
XDSnlTAtwdCrfRBJYTnQjJxty+L7bqQ3NkBx0u1eepxRYgKRurtGi3T7UFmkPu7L
sTxgt0PxnSNLQrv7AmAgq00/3Do/401tdYZWudAiUVFquYRSdzPrlh3X9GUaKkfr
l/uBJVYr9TpICP8+PHL2Djg2DKl/sWupWSMvGAF/1BxqGnHfI1kOKXQi8S4KAF5l
PzEiiVZW7erfs66jC1UzSqZkiG7Bt34gLBUGg3SkE3e7hI7yjcjqBENfJV56ZLi6
iyxTqIgxnzaQjek0JY5LB4ZbYIu4mKufpCuCnDy3tHaa/XzPPUwsa0CRAiyIVg+G
1lTN9e8A3hslSDEYTUVa+5szHsO9jFERu5ttzmF1CTXWN30sev7obffvLUuJNBkJ
Ji2/5o73MXLor6W4wADFnOpIfUIPQYl1aXISU7aIvGGFST9O3OCLKh1NWtnOd2Ze
tkZC58bZsLcAz9Q76EdeeRkTHNiatdyAuxC66z+WLYnrTPLTx1rz+wSgpzrw5B10
48D2pDC2L8X81hEn0F0u+mdHaDkICMB0WtjG+TBly1ZbXch8HEnM+2zpdkfUsDMw
Sw6/fKdh+qh+2I088spw0oKlesPm+1ws2orSR34e1zEWnho1Sxjd8GN+58vWrzJr
yIPGtpDvfO6SXFB3mWraxPRrimug79eZpErdO3zSLNAg5pop5Kff7IrQ06ImCE9q
RLCypZSTqpHBCL8uJULVIQr6psrAdbRP2gHaL+cS4fd2VuKNzmpc7UxpFBvbLN60
UFGpUBwD+K0mvONCwZ6bff1yC1XL63rWHTQtr0ntz2/FsyyumY/0o+99sOe+0AZS
+63oSks9cqoLh3sJW2SsUV6MFCHTkhmTBxKOiJGd6byE00G9Fn90ZlcXb7ZYbOFI
7LC21wW+BkBNzrsW33PMkas71bhs2bBZE+SI4/PezHQ6BSZARiTXfYKsJBXzsIDm
y9hzzlm5LdJCyjNOFNT2oncL+nDe3Dn/WQqCNEzL+QjE0IE0rZwh1YjWYPAtPgQo
eYbnJe6O5Pd7SnpZsR8tRixBQPmE+M4NppRnQThGf3E0Gw8Wfdzq+Rlb6F/dWsHl
PRe8e7Q+fAbw6GA7VRNMdSmyg1eTMmWs325THyClgo7RIAF/n/2LHcYsLWkCVe6e
kV9nJQhHar+H0+7iL0+jokljiybEdqqaKz/sixS3r5ZigevVpivPk9U79jJB1Wzi
nrepeMppkLHsolrOHmlukr4v8i7PBEhuH04kPOmdrE3AcQGKOIE7SUu4DMrSxEEk
MOJ2pXywah8tboPzGngi5rcgIL5QAtxQtyQCh2HeXV6vqJfQ7KEXl1tlDbNo57NL
4Yr9NTUl+Qy4JklK/l8Tku3hJWgxRLZZSbybIdN1EDMpHuUyK5zyOY9vjPjye9Ih
9oisFe+eLj4AWFwhutT3acRz4R9Xx9sA15PSmiTQYJAR0/BZDnXwKGTsRMRjlkL3
uFFCPioQ5Xy9iVmA9Dd+Rz3B9+e/5OotV73Rmp2ibrROqzaUa/b9dgQBrrINcff2
dcoojtgvUxdOXczZ1WvOLTvSlSUvS+5T6eSC6f9Al7fN8XW+08Nd82lpKH0BnmoL
Wynwk8/ohQX+1pbkAjnwpNnAJF7PiWiOy62r5uAD6WF4sg22uZkc7l+Eq0E9pSxl
RTqPXUUcrvlboFX+67Y4Ug8F3sdDzKzcbRK318q+SLNw8lQ5NX8d+d/7vo6d0yJF
8R6RFRDdCfVLqscsHmBaUUGLPvUe5/ihyJeWSen64iup8kUCmmWQ3Zqg0nchApVp
rbLuRk9ysr9Av7zZxkCvSzWJvzIaLzlwuh1nKEZ5ojLvKHjI4FjmKarEvDk/gwIr
SqknvJt2m/yI7pjuEI8GfvIKsgkGq1ZEjVEh6ZALffhaWbQgPlE30xOSiRhUwpaG
TB8B+ywrk+CLxqzUFYhg9Io1dTLE71gv3DeIlPShCJxrWSKFVh8lUoz6A3irVXFJ
sAlRtUSxVLdHKHDhSE/98Xk0YMOuHdMebHXpL9ifMZvDZ31Ted1hg1TMrUPheNXn
Pjyyg7AaG38miEfh/CoRQM8YdJPjrFRLMa6Wiae9GOHofg1F5Y4y5egglp+wf4ue
hSH5YccgDi20dvCs/nAHjJZLBHpOp7IFcIJohPFlxw1U7wD4gLChScnxeWhrQND2
KjKJzdD+GSvW+bSJPSXekZ8zlqb47pujKtBt283s8YKP9c9o3vZPYVnYZ73zjQVv
/ESyUL8D7bdSv6SJkNAVwcwfWGvVhpcVYZIqw8a9I06gHHP5bfAlvXFjua97l2iC
yxoeBWuoWnWKPnfpJW/RG43EZP5ATs44zMivLW0uLJ42Xmi9QMNr3u097psoIhBu
IsfFJI1+KaNrDT+KFB6DwVPh9VmwcZ9nB214MpLmuaOfVgL44p8ALNnDhm7rew39
GlLMDfndT0Y/YfOyMqnPTI0bS1UHi0ZZSVWF4NvqVMhZ1xThrHm07/5xBWsJo0Nx
jdl2MWyxMTfHEhZq536HWfDb3B2uLiRNOuYXwTDBUO90XhzXqsmbi25+ZecGLbW1
EzxNz/5lbH0vCtVAWpmVBaNQIn/zImRKtes4oLW2LkfsW+QuLTNrBY40MaWqN6PZ
sYvh+eiaGtICsvtMnt9GD+n9h1isPO2parxysMDe3+RplYnrsBVly4/mheauebHU
7VG1urFflj1na1N9dbdTOnYmM5fN2mgFACeCtRE0Ad1cyp5SAdowROefTsHCmCki
fRcXv8WewK55lk+RnAkB9jKxyTHKW7+/YIRe3nkd1kChRtwhdnKOqeoyFrn4q/Xh
eQ0voqKfE4wAAHamJbrf/A8veAV178qIC9iftIaGdMDpnbkQS9XnGzH9xJ2MLZxM
PVkR/D6iyY9x7ZwHtgxoNEJgcA+Zn9HwEjVQOtCj4YLLPH1klpR5Thswo5qpl51u
Dduu8J327xOoG0/NLoinH87chjlady9DJ1G/qInqBoM0j6IDoK0xVCSEz9GnGz8J
N4EaU37srn6FH8gsaCjPKpaMW2yLvTBSUmI8FKjJW12Iv9uAbB7kicRWSbUUf8jB
7DtRbqOswVHtFIId4mk6tPEXAua87hL+e0a91ni6s2npT5ONaQgkM86T0C1/sDYg
ox+1uiH/VDjF+/BZSCE3kQa7aB5Yg+orRHH7g1lm9HW/aTVfbmJwf0b94xf3GxU1
+1fFkCDxrp87nseivUhgvHI5U0ocs0BZJJ/aj51ggLtRkq8YD01xoEYXQJFDjmNt
nvUgxZap9qyq6WqR4V73845oD3PtUHnMgqge4Zn4baI8sTd8bW7MR53HKQZQg96b
YUVNrReiB6aBI2mup5khJRDOrAkce6Kh0ZKH4x7vp3am8Uz3JX8eqqgtpT/D8o8I
6XX3dsjTJ0qBl05UkwEBNYYqnQR3VZqjvjWc4BXSvAZArThV4oVllcI9kxhzI3mm
M+u/c6HgqkmfcZJ7IYUzkh1xS+poYxXonMs2qv/+OV7F7UOkARbuVu8dO4TSVKXm
qtSbRN40Inbrbz6pBHmX2mruMc4/17BYi2/084O5CSebOiIOhpYR6D9YjCOqaHGw
xbQP49M5iYGWTobcRBgdFqZrL6S7UrEbxwWyav98c9nbkivazP+PU6mCBH949R71
/txVDZWk7jx3JDZgi/CiTnmbjAWNtK4g/xwnOKHGWWX2nJgGJG75wWNqWzIKBYo/
EuT+VZY5XOFYbpZLdpi/bzT/l3un31UsSyRKdrhggahZLKjD7vfXinhvW88z4pAC
QAD2/APLZ8FKjoUV/d6K05sC4w3DYxQg1PdJVFHSDNZmF0+kHFagZ1U0XTKSEmwq
OkBe3PKKDOYWVKAGe/AyC3vS03WIxs7yOqToc0431Rlf8gg6d1tHIsvlVuJSuolP
GR3FJd8uusJDJTpS5QA6ITnXHWHWqavsT6bXqT+52IWNReXhL/Lhgr1ESE5O9Dsd
O0Pt/GNWYDndcUPJTS8pLTfF71SssrGkMKSQX2cPxc+BsXC28lGZ1zpudtw8lXFU
3iIzOdr3P/7/EMEStBjhix9sY80+RVLTtpAtbeKxW49jytXkEEsehkmYKA9BoYm2
W+cCbLz7cJHcHvYc0IL9unLX/JP3pEcWNhHUCzM/WdtkcTjaAzuYfSaEJJbrXTkM
Y9YVJc0b1mzAdLDWTSIZh3XFdxCkRi6BosEGhjuHNWoLVf9z+8oCBI6qYANGFpi+
b7ffAhUD+ZXX5FrVeVCYFh3JBdocwsmM93LAjqTP7Nbnt6OsOv9JpTIPh45Y7cq0
aDLLCBEc/qVji7d++9xA7ACE/xtcAdSQmy+JlIieHgEcM3ec/fFe16BNRYJCnBKR
8xkqeAQHeI9qZB0H27gUMazOoCcscE5C8gxwfaJ9zCScw1QMI3Z8XBzb/bGvw31h
YnXRp5PK96iENFKMBOWV6dazcO2O5XXcRmwV8zobU6agC4ChHVKbh35PGeMXWN58
SP7UyMzBO6CJ/S6f3i4/ZiYpms6qSoNI2t0Yebq3Nvu1wzBcKAwF3x2JRKYQumhr
uuUgp2Yh4yHdaHmUvr0k5EHqKccDEcNHMc4At++FdVzw7spqfNNbuuCO8e1iYwI6
LBtqJ0wI/g0ruPWyU+9MG1/C2mcLBO2eks5Lt3Gizd+E7/AQ842zumKrEFQ6ORsJ
nyQv2ezm1yj9o55GgBuFC9FDqCeqj1REmhLH1e9EAShjrbBdGr3FzkSyu5B/siK+
18yTJ797QO06dAxlvH5ximMIjN/rh1IXJfKN6q+9nwCaJwv+tEZonMbM6VVZcMct
x5a7SwZ59LB9+UHj/13a2TkNp/cQPKpO2HETc0hMQ76kHuPAiTIxMSG8TAgGzcTE
XD074xYNY+Zigfm66rVxhZao3jHB5WP5zUDGZ2XqJHoCEW2aXyML0N2DcQsWKj0+
QXpANfKozDAXSCg8888Le11fm41M1cemcm8EwQY3Xa9Kc1YAcCTW3zqjj2oLAt5n
tjSMjjjSLlleF3PyGyQ5arxuBTaJG6gX/WbnbDbSxqMrVO5erJE2zYMaGmLIQkMp
bYcVU1D0ieOkSwo0YW+6HZJNk++ep+NK/lOFii/PmcZ1G3ud76HxajrnhdIu/rgu
EsAdMcKwhLIpC97XTxQ6FYF+pmEK3Wyv7SGbZ6hYg2i5q7/OEWTNULIIkecCfiw3
34enxgO21ceddbpuj/psQdsfQWUU6CHzAjfPh400er5vl2rLRKaz95bmMXk1vj8w
/HxxNJqvKy4GAACEuhrZZ9XtXIvpnAFtFqPdClKmIudcuPbknZOzbjTyHnCHofa8
1ozE1a4HLhTA9Ls2IvIzC9Lp7adhs97tQqoqL5t8cIyPbLv34YcI7JWXzHopvhhC
5OG4FOhMV4ph60lhDDtx5amRT46W42llc4ertEgpct7toDkbmPDzQ8TYxR7Gy2vD
MIQs+3vtcMBafkmC1cpO1Usjfms+kxp7l3QLW3ZWRp4vffrBDC27Uk6h+SYNgLV5
u4M33giqfExFoLNFMXgMAHfxTwkXN+ylfxIACXHwjMp91EE354IPltdWs8zqkyK+
Y2bbCtG6dhylN6p+fO4TdF4IN2pRDm9rpLmG/A1csfgixPzGprvmEg+NHlDn+Dw8
UC0SGZcWVpu0Lz8VYp/cQ0dYxQS2bJM4g6XTSEY1lBkEJu+3QfHw2TPuViTGxVZw
sD1Ep/3Q7Ys5L+jNcyHYMQgXS0VfDOKq1uF8WDi2CL8vOiGVqG5eY+6xZD+4Uh/F
gimhjgKamidJe9AWXlfhGNFrl5tmFf11dechqBh6OG+UhwCBc/KNKvKrj8hMlMdj
SJxYLyeVIXLPf225NUVFXt+owuD36ubUnTl+yx8wrqPNNb5DKC6H+vsi5C8P0RJP
/qLG3Pi9F4zdTnBw0l7kqpT/eGhKRkciZMHkm+VoI6gsQg2tEy99dLnz3cAcoOlu
/8dWvz7jpxjbDQALCnOjFk93cIc1/YqvcLxlaFaUjFdX2RCa0CjtkJEXrH+3ieOg
itHUTcEVL0Ff/AfT3qZB44lVhQQPwYUYyY+iQnP+/8Dhy6vzMHipjAWaZ8mv/TPi
c7cbWTwybIRTxCVXteeY8Jv6sOCgwNGMiddJpymfx73sXgoXczEdhcx8ZhFEZVYF
ybMUnDYMtkJrOpWsDlHmH5Ugj/tWoBG89rAo5B/RmCVbU8nQliedBCvx4eZ5EV9e
LtkqvLDbLXIukHkVQkX2LbH61a7hZl1PKLBto3ggHyQsWvgbt9qQx89hvnP9iJEY
vkmjEl0lnNmxAC8qhHKKw997moS4AAfHNVf69SpuYXhj5uft2ukyOf09/TFAim+h
+zdCUUdOduAGUnK1ztYz0mGLZYDsIkQM0tmlGQxhIcwsc8TEZYcoDRMC+echk1OZ
bHqvpT41ogsNze3FQZIsBXwjDIj3RX+JtB64Cr0SGtB4ZNYxVsAh1qPx4RjsMalp
j3nXpv1sdo+Afjsfc1dA5AuJuGhv8mXT87q6Yq2+NxUhtj3oaLHX1OtUJeSFAUvK
6iIOSxywbROaQkJ60adwulpSyUc6dg0HHectplmzHGMDeMQZVpwoG+oqjdD0OJCK
+EVSGCX0io7cqoexmVKlwYwHdCQcC3RZ+ted8DsZrf1MUAPt95aDyMKgwsAlV+Ni
CwFDjEQASAOOA0abrZeIeeGn3nEAgHH+t0VUCXuBdVYoXvUI+vwQdm16irLfYTlA
g9YBRomEIoVe5YeHJZ2JRBtJtJ0AXMDnzukos8ktaJ/J2wamBWevTUXBsIKtlfV7
0TpZOoBadCzzzAWPy8bKhKANDaevaI7ZC6L0g8y4hd6mxKdmPc3Z1PCm+8iAZh9B
Dd1fbImvzruYCibn2AZNE7KYI7IJdu7EB9DyX8fKj+4Ph6xv/XI9QbX+oynkTHdv
e3BO2X15CbBpa2KlSdRjnSIjPqrFvqVc4e/7umsaUwVC4LcUp3GQWgcQ0kKIdBCb
fahtC46EiRJHMNWVuC9rYsHv3ptk24Q9xodjeFpmdvbGwjTuXWnjkI9ESzpyZnuG
EmYy0+I7DpB/bYm2A3LbtrTvb/LGg/I7g4tTjG84Pv8Wb1hLoiRbC7JEKIQ2qink
7Z/l3JlXbiV0PQ3GI2gLf7G8iJug9ZSs+ClErxiczTJpiM32sMXd3MwR4aKs9cL7
BxHN0DfccWzbw8Svo9OmXN80R2qO2N5Nv5k57nDKktngildtw9EBFZ43DgbPwHSJ
3ng8C56g5osJaWKJtnv4a0HEaanEpm/R0Mu1LnFsnmHBhVx4999G6nQBnwOd5hYi
Za6EguAkoCT+F3va1lEDuwzyIzYGlmEQTpRzsCJ8yJRJ5taBQZZe2s9E2ta9Mnxo
U1w+07gqMFrm8g/u6syiX/joPKCxsp+02tTzDV2uoaENY7MRDcHFZFUulhTKfpNP
EhYrUoe1Z2e+A8xHEKYA7kZcQzzPUbtjrGlgmk5tTiOJk61mZCmX/Ufjxgn8dB5x
b5xsRJSFdjYJ8z9ihUNBL1hRvrpY5SN4/48qcDYIy1zDvx0cDdX0QeMflCWydDbo
R6pJreLtBXgpREh1b23dO8gzBZXVpQVbDxNL9RfMg9eU7xSCn/512SY7ordJcnJx
tdRybSubLrhAh+SIdMu5chMj6fZMT+twj/9XjDCL9+JIL/SCHwYLBVvMio3A85AE
xNl9UERuNJ+NxN8lEGAUEngIqFWaN92UmhwtTriHlsON6tjM9pF7MVTBB8Agd3Dr
sut+BBrsj2AQbVdd8xRt5zQBA/Hlo4m5KH6gwjgV3RD6/u416uRZJG7nx+/CKo3S
JK4dCPfa+eQQcZE1aIY5o6ALUhdNCdMTDEaw34aVWq/WEtq+5hxwhFUnWSLb002/
R9XgPlOqnEb6O4u+KYxJgzx8CRDb5zTOs0pyyzNjxToJ58gPh2oByKz5ot+TqgSj
l90RebV/0taaVFqLhCYRSY7+W+QRsrELjnF+C7UZyxndZB88QZAzL49/7FIpWH8u
6h8DnsNTJLpJIyvIWOWg23SQCJIcokCACb/Qulr7C03JzEaeW6A6mtkFuVIUacrr
yzPb1TC/KXgrdIG+8qCwF99OZIYS9/2Bn2pzPaoQ3DxU1fcStkecR0BrQ/BVfQS1
Axl4b9Ryl/OuiVztkLVyjQgFxzpzbvN5jPYUEDwryq3aZRSKwWPTAXIUr4Y5gtsf
I0ZDaLHZH7GoK0R3x2014EaUyesn2JXL7k+IJGCRE/6Mq++9JETRcrmOMxN7G6CH
okNgubESFz8gHz2uKZ0IvKn5jjiQimaI7ArMhIcRb2sOvrTTnBwbvBUY03DjBGG+
XjzjhBYfYd26LoJhoJvKhDH9mh5XMab0+hHCx8nIRXLe+bh2BzbE9RT+q5ZhOoiJ
zhUZRv38HwTKNiZVQdHpADxULS1I9D+jEWvqKeABs7dgI0kUVC8avSlkENT+UpBV
IGfvBRSuAXjE8M89R31l/zwkqiFZCESI8Tt2y3gEpYNZ0YkqCC1ijfnsU8OjeEIz
4iAtD/S7oWQsSboZKYyAU8WELkkFLEUa6OPeZp4+LsRxshQaIpsFaVY4iYORC61L
E/MrUnwtgNSMO1VOPI9on4qwUxJ/NOA+MrrcpNaBtxbI5mj7rc057GP/a9qdZYQQ
bi2Ohthgzl8wn/MQS2GnbGWDSvC+iagJJLQw8zJRrSSyGgwR20GqS/TYrwEJeVoW
tZ+FW/4lzhgeZH0WeJwrtA+NPL+SGc6TSsCIdf/k84gsXWjQowgI2XMSzkEVYS8F
c/RyeJ7bHhPdhde3FzvZRivM9HDQZRdZ32X9waimyXK+euja2GibwRJ+XVguCA6r
i1+qr+A/P/P9VBGqNI5Wt5ghBudtX87+Re1/gyIcE5nY16/d70k8KLxrrf748jDq
w8zhj2ly2A2QimHdpS/LCiWbFDVvDMz7j+eqLhynKSLKP1N2Q6Qg0aUT+G5kLEA5
rMVyF8GCZkwS4tbczRsM6bwJmU0GUU17qOp2OtWLBsIS+HEsYM5+WiDGaqtSZF0Z
mlquNEzp0eWhZ1zTD/EV6rxtFYj3EGnfH5CsTsHlCltL+OzclLJPEgBb+0Z5ZhQd
XIuCjoul57odJRRlr67/fdIMSQqypxJXfS/mXn7KAFGbECSvOpy9nX1n2UrhL62O
AxxoOu35xdPOpij1B4AsWfXk5BK/SBD2UMTq2aIrL7xlAgmlrDWx/LhSIixtIFqZ
m/JaHj9zNSS2wjbCbjTDGljzfkrIPcBNS3H4/vXIC4JhLgGjX0KRECatbn8AvK4e
f4QwU7Z68HQnXHPwAlq0xwZJbQ2jljxdYeZQOFqdisqJDxxTIkuRdagr73QYnr6c
13U9JqW4YAWc+NslfMnz0hD4crnSotTvTs1tn6gQwwuQ8NORcyAXeT5sAM80DM5y
vnFCh4AaXwG3CAElsNMIkwFrmx5ryPLt3J75rCLMP9EmB0nEPSVIt1OAnoCuarY3
SWAKcb9W4whSznWIUzOExdxM37jQ/ZO7QPUXXnMtlRj1Y8fmEN+D8DaGEoOtnfMB
rogDDatNvA5qb4PGvQNlfDrwb0E4ivZgSm/945VoeijalwvGgXlJT9QXNCaV0+w3
+c/vZoes4sh2cwAFRQ899atCZyjzCqG/NrCnmJPm6ewgm8OSrESatGgtJFTBDec0
K7r05PKaXMZ4C4xbFf25zu/AdhBY9LqE1RLDfCC+fu/ov6JWgtXHU264JRcZI3tA
EcTNCl4sfx/P2l/TkxbRWxBg7q5sKPuj2jsxXnGH7iXdlxrB5NLKontHsRa8GJ4m
ArO3l2rp3qjBgPklvFgKUNSlr0T+IhjNvMokPGLnkf30bLMi68jZJwgzKVThpGAF
Ib1fto6QvGQSWAsF5y22G8bE7/PsEkcnDhNI0gP/ei8CYvkrLjY6kCpM1uEpRnom
Vkpk/Sx8MRNqB7RSSO1tXC3Ip7lqkgoj3CGN0MKvEkCR9zVBQEOB7+ERuaOAaLIr
XVYGA+achC3bhepw4b5vxU2VeQNqe9IedxqtWMaz5i7uRFFCkq+EU6C4byN+xxOo
oUhrk161XljWDrgFPbAMTUv9m1Vms3gw1FYNxx52hTv+V27GbNNWm85rgjz1B/rW
xVQUNuxtpwCWg2QK71nUTnsL1bCKdfg6+oXQEVXhLEXKVOMmujgr19h5JhKoYj0w
AcDjBnribXf1m1ILSzNO5POZTZi6Asu7lpVhLPPYJv38elSAgFKAEx7tV6X0l8vC
X5DqRmwD/8IL/iwWQ2y8yak1Wn9Sj5cFWdVsJqdqc3ODrTyqlIYEhEmR9Kq149cO
uNSHiIo4ezeGvDe4A9Gg9/YppGOiqGtM+4jjQgTdEw1dfYP3YvKdsxgBXEygha2p
1POmuUP86JWQw1KrcHQSYOKp6WztRqrXuVZIeh3gCkNEscmfbITIy7BY8LuOytwQ
l5vpcbTEbK8kl1WoPPQVrP4WpsjuPkV6040VL032oiRDiupk+SJaJGeh6FU38du3
TctvHBewGQczOgB13S6XSRQbfwckNnw/zT10wXkLKDTo4BcWLsgalqeRlnhA6uKc
M5H6IyncKvJiq8dbuSgQzZqwJhot48NusLcCuPuwiMYVqDYlLy1anMBCwJoCZ7UU
ylwnceLFEhmELpGQLILS8FvQz2uhA6oblvrhIQL5tDXGqALyywV6T070GwVSSjzi
lLdVHfGWLxLNeGCzuxjVtabUElbyZcXSlxWcN4LSt/jr4VvL+bb3ECiR3dv+Yq//
oFhZ8NvTZQDAX9yKi3W9b6zjQaCi7IlkkvywkIj7hbHD4WoZ++rzpSznbSx6YY2h
sqIMyjsBLnW8dpJFw8hzlOwYOSTtNLCHwM56FpBd+MhIdWIndImkxL55BLCjRRCK
GBSYQejdUf0FkPgMuaqVWgno8lXGDshQ6P+rHVP9e5a1m4M5SR7lCSF1qeb6DZm0
ERpOLgx3zCPBxF/qwSr2IUcBOFdTPU6ApOblGjSunHnTlTdy+e8DFMoNHyTTOwJ5
ILTzc/aw9uKMXwcBZf8xsDW/FaJMYYBVJKct0S+IpB7q/RKwRCr/zJaYw69q7sy7
bq94V4eCntIsqnUuy/LvmhJbEW/TtacyLyIQLHTBw6UJmHdeq63dTzapmEF9/e+c
2yMZp5+mQetXC76Rjy72Kh3Ay6/mPjhpN5lN/w2aPuwO3+CAtj+Wm7F/zerg2UgI
tJTLbdlEEXCLLpwbfRJP7NdmzRsqJR4PusowAWm1AuejSawFjt+7zK7SgF2ODrgJ
buoCafUtkJoM8h22X+P2+lC8QHSlgpYT6lTRCQpnlArdXpzhDxZf3c6mOTRcmCv1
eQQL9EP1FxYsqOPKm5shZGLwcfcafqU99qbkOv9X10RedIu4x2Ze2RTUtXQmX6jl
7el1c87v7kneh/KtlzkioEfW5iV6gqVOc9/3HcdeOGmqLUXXk+ecbL4wN96xX+gj
pGcCEmvVS05927wzPCgG4Zkdm191V2ASiJUAOB7zal29bG3OEwum7w6Ht2TIn3+C
SrKvxOfM1XCpVw+Uqnw3P7irdym7EroizdTgPOKyr5cbwWVkEQUIqFBf6kazwUQV
eZFKtchMniUoD6WhpbAnpbmUz5N1gXv1KW0Shq2epTg93dKivVk47lnA0eTPurk4
N5xS4GM/t8kK1h7v/GMaqhSePqw+LIe9/ojRLs4sYw91kJceJ9CadgLHgiNUqjmX
NTX2MTyTwb4sIccnla3E3VZPIN0/1OidIZJQCyL84Obg+u9zOfpMm8wkshfYVoaB
6xUwdMGm/hZlI5MF7euwr43snXWbmjGDaBWStlebjOO/tijk5Sq2R/xg7s3KLb+2
AVuI/ez4qdxLBt3O+7U9+CjjaOnaTH2EpRw/T5lX8qi7dWJFK0JyY0lZkIAapnFT
orfxTqGyjzPMhesheLP+ivrI8rsGXSTHqh+kVK8WXdc/SzBnFq6gd4pBU8+uMqvY
oQZlnpyxACRsOLPHvR7NGv63EN/YPOz++HUaLQAALP6UdEPlrMrrhJgsgNFyFA0z
Nk6yIzKb7NZ+j1yGMCU1HSqNWx+Tz+frpSeP3yxtpSiFn+Ir/P76zkJ4icX/Ku9Y
y9W+1MwhXaG3Kj+jdXKv5htaAhRw76jI79PglxAk13o3uvKIQV8Ejbn+2MjGZPh6
bb4j73VpmX14Uvx5Pv7wYh5wt3ogCcE3aDt81zST3JQsRXF+5buZxo19iLPTQ8da
mz8UUcDRshUG+287C35pXk+ui11hJbvouQBQujR2Ue1Bgh2FN4a+3gNwUUW6o6Au
GFGAcEJbfQ3mjwu1WLzgfXvuo95RKdpn5TgGMFZBFG8kVIogy3NNLOOXZ9FXN3u4
TYNnXYBFMgSx6k507fj8X3nlh4MoyDVLG3/W3YQI9/CcraoM9FYh7l3gI6uCc0uy
pb037JOI2zlAyD9IRNGBNWGGuI3JUkExBjysg+5wWUXcmK+9IrgkPyFl+X/UojXr
UnLtXQ3fD410Y8OWFHg9ObwaGVm61Uq0STnlfEJ6MVq/lirvF2qLLa9IUuHFi6EK
NOJY7bRVWo64WD5k+RccFXv2a94/jSry2FtX8OrkNvta9JGb757xu1zw4ZNX7XeX
UH7loauF9w5nrhWwBV655t89kKCcbIN1CXGrtrlJE1WaNF7kIN46TpTtGWEBZYcO
fTardXxRN484D/1kXdd+gV+C0akP7iIFihTjiphpJk3U3sbMwwi+w+aML9jeZ/XI
VDTFlx+4+2we8w/WaJE/xs21XlqDvrSlI8ARYPmRhJrL8DWyPBx4f9suBKNfKhlK
u6bihBVLr3jl3Cpx+FWyWAaUqOuXTiPPS4IIOnhPeX/oaD7yaZGpWcmnyV68YeUi
+YmsqoyHiYPFVFOVavxEA8Xxm/ZU/VpGs7We3R66duCtNwTm+zmUPpME3EGKR483
tW6oHCWDArvnes4BAJEC4/9xxU/ECmakm3oW0EWnugdlaIrys2rBgAOvCNQVGm8M
zRpJ9UXNzooaXBwPuMSqdZ0X0p0oNhujXs25BUuHfyDcfjG8waVAIr0ErrZh5uk0
ugh/oGkvxJEYACiJ6EINhi+AwP3b+um4HvVSvBJ5MSij6duEJDSMpW+Bn6QpSA1B
gN4lYsgIqLSPOn1FhquFF07I1pza7yBsnKIkqPkgXybdcqSBGfJj93ASyU/v75X8
VfulJi6RYnj7cwEfeL265oF29A8SZdLiQF3w11KDK0hB2u4fwyT53WMHWT2pzcNg
xMdwxq4xT9fAwuAY5NaqZwfK1KRDYigzw5gEaHE0swTb+0x+LLPVx/jDhwMDJ7Tc
UtQbxe7G84hc8TgSbVgbMX3RaPIgtTrwoZMWXuDEpEE+eFB1dL/Vx+qJ6yiNT2i5
aoBZ+tmC090FPC+MbC/6uhXjzu5UunkTohettEY2Ti1u0O5atJXzrbGIomL4MtEw
Rfw6ooz8/4q1q+shVIuOaJ1Rk6OfdXmypWFO2B+RIMcOUpt9EcgGom8LGqu6DABB
YUx2x0vK04U5IGjzL5Cf4gSauteT9/10jjXGSOIOytNBHoJsNoT3d4rl4XVslOIq
uN+CtwTImH3KPlGM5227DlKuqtSaokNdaXuVtXY1WcvJcCMGLbZ5zO/wO7H58he2
ShCBn2KZV+k6BLRdiZK2xEH/qPswHRO3qy78vZUENMaKREfwVVg6NjH1Z/0L0NzK
2DbEEJFL9bqsFo/i1u15PBkEIpOeVMB4eDYyxVZE0DxPksnpTqkodhTgmBSQoKUn
QchoHtR03RmXqw7mWWnL66XNb/9PwvUeZipXKvbCocDt88dO1nuZ2nZqYG5Lh6sj
JC1UHxPR8JSc9ly711w/gvC6UjknxVTZ1wGmz8KDGKUZjt29KfwqS2ND90sOF/lq
smAYknMlVMJOhs7G4NmSqPIUM0t24UvxsFPd5WvDa0K219tdV5FSdbMlyCPC0tF1
oW47j37nbEBiZ126nfLmgV1Z0WroVgY+3k5Z0V6vUCVcJ3s2TEumVQWanF8jxQh/
+cYpJ3LOTsPB2UhEjrQcPQLuvLXLxQNhmWWt6aYtdIy0ql+nAgQ4pQbDbVxfJJ+s
Z/0cfzOTj0NENA0j00S2/fgFBZlaX0DzcRxgFmWuytKOlDRjnXASYfZoyTXBLiqR
mLE4197opU8u0CMQXbM1/bv/rvltJ1R99/Q9HEDLMCV8IvujAdDl/0sooi+qJKDA
SOQn+Z9iyl3LBHPcZ8bhsOnlwm2E/DsmADxFvMU++lEdExccbeYOcJuggt1ae7pk
n9xcCizEgA+mo3bD5jqcYGxQ+570vQvlPaCSI7mi7Z525BY0iJF4Sn+SGsNgGm7O
mUs6lZ0E1Gg677q2SkbvCHNEf1N6nVgoWwhvtcbg5Iba++pUsQPjoM7chUfqtY/t
Nbgm3C3EGbJ6fQiQmp6t9YcxY3ikgPLV0LrcSJuObyVnDbsGgkP0eOuThLXORJyL
Ai2e4GEXCR2UndH6Q56Us+3SduMttlnRbiPFer8yEjePQiz4e1IQ5XKIX5WZfllL
8zn+8mGmzBgkNUwkakgwMtWJkCPP2oauzl2HZEHi5iBXUJwpjo4mCNu1jnih/B+v
iEYlzWuxXCZ7RkZ/bliU11ok0syYEBt3aBNAg+IrvojWkZgF+WD/46cDriV6L3BB
2or//IuzWFosHH3A+aLxNhkzru76uvUcW9k2yeBk1f050XEpWB/mpu8aXsFp3iua
myDAFqPWoy/E/NPEZqqiOYQHfgowEJQjMRv9G2IE0n/XeWM4+LdTbrlQOSwLQhs2
CZs8Bfcmzs+s6fkoUYtR4m8nlRla1N1WPAldOfOQ7WJIgiFTgg8K//jz6XVKykGh
m69yflIY32e110IBc2GcKeHDo8/rFSsIDTV5SejaC7BbyEPzCXrCzZ1Lri7rs0kZ
Z1J9crdTl3qDNpVqF/k2lcWHi0GQxKqXJsvZkqZsP+LvKaMhjfvoOWI8S4g1Sje6
PkZRQNOtu2hnMzDQtGCJm8aTxmRmoxzsIMmSKbjh91B/de3GKaq9VSuaEGM3WkN1
K1OMZ1qYLeAaCV7QSEZ+R1VzyeHY5ijZNcbWU1cVxFJLafwBxNfnyFTVoWxnIhxb
P7QijukgCkndPCDwmHEJbf1ooGwPt8w3fituY0Mz79QCSj9au86PFBy/smByzgwt
aPfPO4uW5fansGLI9f7666ynkcYet1T7vg+t31PTjlLH9A2IyBP4Lf0Fe4qyKF2R
dnVIXUziLj2pqwFtPfh53aM+oEUXWdsdzC0MOzt2o/XBSnXfnifjbOoaEB7pO+wZ
cObgKYY2Zd731ec2S+uGeviaYxQS4AyAl05P000yWqRewjNRDCwrAyp5kMEWl7Z7
JN3duB885WTzMs7PhBxjTT6BnXKNhqSLp8vZIW/V4ttJFIiNbLIYApvKthI3cpf7
re7PTQse0J+CCblY6uxY+XJwDElZPO4a/evsX0DX89oCa1mYZCX6svCVFA5cHwIO
G+WOeAfcT/VQXFz/lC2ghpvCTgO2EEwqVbReCk7tJorTDya+YS9eJEzCSVrHKFe2
W5mOWn7rb5nEp+L9baLlvdyvE/rnJil7vlgx71LizEGbBHfh9KMt2KzzQlxuDYPp
IylvGFofftRgD2QAP36yhX48QclmooAa7Dk3evRw1b42Dz2HIO4rCxPaZNDuB3bz
Gq52nn6A6WoTe4qIwuI8XeSfd9g4U7BG030fg2/5mUJwQToxgMuJtlegldqS/O2C
IkPnaf4ggBV0FhRxOw5q46kjJ49RvzBJxtEkQFS3DTE8et4616o6gQF8yWFYB+DF
5NOAtArD3XcjCmIQw67KYOPgZbiH+WZ9KG3U7ikP6hI4gwgiFnS6IqreVs+vdE8e
fk47Oej4Cnvj8me4iktwXeIYfh4uN5J4fysjc+ZLq2NguEi/Ivzoq46NsCbLqRmy
IMSIS9lgh67Lc8ozhZyi66TBup+pU1kVDWX1+G2QWSlyY5Al3Vpe8AEyxJMaDfBr
EOpkwGOABAOnQr0lyIr5SU1Hlaads3L5182Rh97we17w/DBDmNWMBG1xWTxmlrVr
1WbBzykZ3J4yu8I5R4qeYx02w/eUPv5TrrE2OEpDM1tb/CSJTwWDiUduUg0qSQkk
f9AY5YeWxCqBTkbqlKpuAdAJvql6wE6L+EhhhuofUTdCtiZMWwTWNs+xbv35qUUy
VyHRjYGkJsAorB77h8MdTkH+/AQYqV0TRcRmGJEEwxDze/816bOYLsThj3HOC/ck
1VLXOXRnbMF8reqCPkPvJkPle/E8PICSgGpwCe9mTVFrG7Sg4BZ/a+65zb9Q2gG3
QK8f0mCoAKbZng++r64jq5T9oVnb9kt5rikXOvBS8uq584wYA/r1mpuiKkgwsheS
RYKmKDDrlv1a6qk3t7YwsQJIjtcunWuPSxlMjBEwrW4DpWVrh7qCI57JMi2snXg2
civGa7S/IhTNUPiL3u5uYZE+1AT1mRLjZbU6AUVnDnvIRzcjXToiAWXzQlal4UPT
txJrdgRbIzP3vRoGTwH7zXnNI4oIYGsZAjsR92koB95DInuSiINaXzJesU2oho9A
p+W/epCGlLapKK2DXutleye14B3rdg3PYdPjS+ynlus0X5bH/B6g8rg+dA7d8qEJ
nvAPeQoGzj9hWKUqM7iNk+F8D0KS6VJKplqRf8m4h4v9DEDgyhoPwNM2NuPwCIOO
ZFUvktwoCnpDvZLLIynmCezMHalq8ON4j+yRiVNuLrg0LGP6DpgkYxN5igyaTwuI
cJ1QhHJgqln3kYvvOFCYkfHlSSw50pKTH/LRPDHJ2YwmowoCHHvKDssE61sYzMDo
NR1gN/jKcdha4W+IarH1/z3AeYqEDN+Tf2xxbRH3d0NAbc1aV5sXhlCwlPZuI9tu
wI5S0m65sGCYWJZ7BO/1XisxI5f69z7iPWI6nF61fV38PFl2sc4nIkaNIafh7IjJ
OnT4Xpfluwii1IqBWrLxx45Eytk1nXWOvGWKC+bM7x4UeVXB70uchzzux01SOCWa
dWiLdo2ZM/0H7+94bwuQVhSd4bt3A6VY60eGG5pxFaXZIbFqlGEFjFzFBPvguli2
YIXeC8LtKWc9ebcCYOGnC2AY8FkhnYBESkKRBWyYrVD1UCn7CjZoPml01tAc3ujQ
hkl7xiTFHwN0aFdWunTHSG201rAC2CE+TiX/STnGRpALSj7SAu+dQttgw7Qpy97y
TltC26NYUSQd0fk8Yx8Y5ANgj2Q0VS1/S3ayZVBKOG9ZLkzKhrdykqVhpSypodig
XbsY20W9mta8n1K3QF8l/Y35bgnmUOd28+JmsX645i78fg7Ue7EsDplrWcITFYSY
+vJBxt5c4o1yqvA/pcCpXRHQZ5TI378JdSQsoe6B7jKN4n0uGT8Nwx/aj39XjGv8
I1/305LpfDtDRn+z7Nx4De+3SHnKUAuCnz96hOhhg8EdwYCY+Mrc6YMMlCULKR4E
MnNhRuoovEyQe279clwFDy2Ncv2LefEaZ5IxGXr0fFlCr0odyJvWUFLefmxUnm9U
Ut4E0PuVl3937CCp2ssyUUn4PAczFjziiL7H0Qe/+5MkzfKpq/Kgjq/874nNOBxm
DtdxCF2pvzAnDI/50Y9QOlTe6v19OFUi3Qx7foqyLxYiTDhjbTwyDN3kXI/7cK4J
uiMESgzKv8HAo+gNkN+YfKrKU1UjATdXWEUqw7ZxADdU0T6r9S4tgTBGmXifW5Xi
hj1AfABFPB0D7Re8pRs18Va3VHjGN0vsRUuk173inyfY8QRuU8deCWMh4q6N04+9
QVvyNoaDmH8Aks80pt01QNlDdjbqXoZ7loSsqT+jlXwkNIvv9ugJDjOEiI1hrvTV
OGz2/1iElfSe/HeEnrZiGYVKPrtS3HXBdGNhff78mkpdDDRnYKMoN4XWFGl7nbzO
5c4KqKE31U+W0cbCvs5EKQxok7pYQoqVYS9Hd01qiDcRzCUAahm2bJohO66XvYcc
x6yKH73pCUgJ5xPu4b4K11w642ZUu38VaQboIJskOIULCx3kmmsNyT5W0gve0tEM
J6CA7Khv0mBm83UTuWdZIvdTkToy5aiOrt20pugK4oqurZgHxXF2A4u+Q0Yh2d7A
7zBUgW5BJSi4rxK93YCwbGeYOeBPgX32UeQqdFonx1gZeuS3RquWt95kwU9aoxhl
Dq4J+bIz/NNiAqBuUFvnldLhK4J/ZhJnzGiOmU0+lbe3OegdJNXkCbG1HnhpQwJU
+92DFj20kUpKLHcmc6qF5aigbJr6og95A1R/7W6qHvts8OBXmKiJuI21IXx0+Rzh
HlSnqZK8VhtIUhYa1qtyTvs9ie3kgzFazLunKpCJgesY8ambQDpCd5T9pb94YA+6
Gc1FFgqgtywESZYI9Jo3XeSW5uxCss4KAH6Rhw5zcJnnXwj6MwcFoVEhxsb8b1fH
rSlsfgo4VQ51LcCmS/Xm7lL9MIU+5IKcwB4O4GoW5rw3DjtUu9uW8c4ml3aHQ4Sd
ykvIbw8GlwTE2ByCjX2Rte1XP5u5HPFXL1p9YNcwqoaVgHQUHKS80XvrN6K3sVba
N/mpc30Jz3NFJHFFXwI3dK8TRno8RO9pPYM7WCJhsMi7ykoDYt2A3qtFLRfmNBDJ
CPuKUeRXmYp0lyNZRWBbZC/t7tMBVNq1Frt0Y7teA1TJS3JlIIPMZdJoKC+gYVNB
XP2HhxjoKg/aC3T+dRW2okS30u4QaSy3sR1h7XXkX3zvjDwFLxDBe/A32QwKP0Cs
NdAPWNau+CVmjyn2AAEYf+LGIMe5BUAPwcWA6TVmBKZM9r30e3S8bwEXl/SCuoaQ
1mJ7gw/cf8+zkHKnczv42mjx/MbYV5L6OG1y0ZegVMI0rtr6MsT86A3ywNQPjmk7
DA4zk2eDE9YY62GxXCeW/Le0Pd4LVlcbLAF8PWZOhowo8ccgUSmImSxYe2XXQy9B
/GO6tUA5umRngfQItC/OMs7Np97qMzZxtt9h7xdoT6MrWoDWZrjVOkhltxW0pA1i
EXQtlqK/o53cdNqW3Xwpl1cBOLUMZ2ld5YG4GxAEnssq2wNmHdhJBW75tevCXgf/
Ztd7B/syKG5Joa/HllDv5RDRFps/wMbFe8ey4VJ1u9d/KaAEGwIsJcZtZYmWTjYZ
GyKcc00zUtF+prC8oYZcxSHuMDLrorGsqw8M1TfzaCOjAeXySGZIS0jOQkE0i3gA
XItrqirevJmOF02Vh+ruSeDyZuj5i5tqzmJpC9n3ABdel2ySDZimZedtdntvdpFb
mpLOFAY1HnaWprStJdoRYvCXrcDRM62klzaJj0bf98KJKAl8QCR+hWcCpMEs8FQB
9ckHebDNMXHBBQ+qaTpAw5ylQsBrx2godeEdsmONg7topD9qGKr2EReA4RLtM1wK
GBb7JuhV8+BJZ+jdVaKD29W5CFQ326j49yBldfUCknAylFw4DnIhtPGduz3iCyN3
snouvPGTPKxw6KXtBDb3rO1Va9lbQ2BWXReLkWXlRbBeFGfpHXw39co7JRJWrdtq
QOtBdqaSaBEoAEpsFSsFURDdV85M/FodAj5jbfuq5h+1A1STmRERn8JOCSMTgvAP
+UV+ZV+8e7x24CwQHwIbtgljyu9l42+PScg+x9I6/g+4xYsLdsgKTolPxmNv8LW4
QLr4+nbSwVQmPwNsDgVKHHx3PeJhugSXoAHzjPcg8QF28esdbZChw/U704eshnOi
61tivHgXoAlon0L2pH5TQYhdKrE4kP7D0d5pb+m4FJ4Oo7T+siOXbp6ycqvefXgj
+i75/PFOjp9OgHC0ZqFLuL/hBq6Cg6b+AKf0aRU4ke7onIJSJ778yzKCDMZ2+4y/
NfwRUj6H1RvBNV5+OyqOisRJML8sq09fmjWG/wSYATMjaMAiGGP7eLBa/XJOLvdw
KkOhtPLlzYW1tYsDQnAk1xt9efPmFHiz6O/QRpHlc+2Fw72kOm4pIy6dA+lLK5gj
d4NhXg2i7E6QnpPQGkXtoPfwX1aFXVh+vJKu8QujfbrdifZZ+8Bh1QKZE9fbbRy+
wIBVKQdZqLH2vJlPyjbH7yIJe3O1YtXZH8M7pUPwZ542OSmIPKxAb61Vvzp84+yi
k5o3KRC7WClaLbJoVBO8C18NrJotQZnwR9v6tAx3NGz2dPJO+PGhKT3FkQDmh3V8
ul7PmkWKOX7zjAUUWtFLCSWaYMDP1j6FdPDhctA/Tajv9CIpDHQnqSiF/SnYV+vU
5nHoDLo3XIpWxMQ5GMCn+vCc1LKZL7qJhNyrlww9KBl7A6NF0uVAoTKt048zhtNb
IzS4+3jCz4S7W/t5vkBdKG6q5mrOajSam0ibfuAsXbad30/BD1AN+XbGg68VHc9U
2wu4I4W7TeDjk1gDz0z+Dpvov8RUpHSsV8ReXYYTlyixv+yUbhS5vsgPXROqk4NS
42P18yRPvMW6UB3lJ/mQigp5gyFK0CFSWB4TJ9mSJa4ZOMvl+zVLQ8NxGX1CUeIq
foAgzCH9ZP8eeaOZJgqZhPNl7O7+y9RcfTXtUnFIfXrK9MJPOHJG8E867iiRbg6J
jswqxU5V2RL3H+YWZQ7glSfi57PyVn5RZf9CdnZZ+GLFoXMUxxUoSLh1XGm9leDU
K35NTXqUQsR8OrZ2H4Ysq3VBj68insXo+UfCoPabLyWtxVROZCWC0BrsgOdUiI72
rzT4sIsrhD+g3PfCqj76iI3kR2txbmqeVZvTAn3fwpGZcxXaFi/ydkiKKcpYNqfQ
Y0cBckKKyoX+vdsZ00EAFgtdBf5wfO9VcYrrVztTPXAf10GJZN8bQjO8BluZdiV6
jUc6ELQaJYgUyKbPDmJF9uv4izHP+q6lV16DnWZg3kf2rwR/dfGEzsoJTkLYdKSa
sHANRzBT4VTgVtORUzMbBS0GruQKeOCWFJla9h687oAveXs+aOOWStQBvsgWcMn5
9hXQdcMbK+wSePXe0RaQIJCECSo87gaud/mubHcN7IHp4Y/KwV+ejrMUAUH4/ZCL
hnNGG3m6E99ZKMeVlfOREZeZ6K0MzQpUcj0nG0QBdIQy4a590WgjHw9SqoO3yhjY
YqM/wshSk3tTHN0MvgeFRoXkPPta2nib0nFAeh1lHb4nl3oQCApNFriYv9AYGsX/
A2Y6ZYq9GkLpog5/LtTcK7wLaTOJwCU7vng5h96VK1mSkNgGpQ9bFfIxicqWDbiT
uMnIMuMX57otonEKVQndWycjQc9B9UxGcGmwMUMn472dVcpYUnsA0RDa+LfOfi73
LAAeP7+M3jMNZTuC/8YYdD2zSyfOonKheWLqo40TsMJxI+hwGN4ckRZArt6zAZ8N
tr1vkTDpu4MHO8JN8FEAONFfUXq3x6ADjH9fIW/o5kOzzuS+PFhcyxAf6ALbTrGN
4PwNO3WZyhA8FcBomr0EU7jrUozDnKa/6DR2Yu8+RxO3ltmZn+KEhTYSlTyDOoH8
TDP5xdwDuwc45Gb2gwZOwv9lLUDV8xk8GCiDtN6ObOQ9OMvRfFIbtQgCBSRI08AC
rHqQHzfmcjYUFe7h5NjPcXp3y01pftcGsQEpQ7MERI1twBNzbRPr+Nl9zLRpyjmB
dT330BbX898EhCbrzKYYLKazb5ZMCDCA6EqCYNh7XwoTFnTEkTIXTnu2UFIN1/z8
Dgpf0aenU/fFf/RffS9v5InObr92gds8U6VPh663EfBkQXlWE3QtSHoQ+7bfHqKx
IYifttK8NnuBOZ4SaHQSzTzniHuqKSIaYKGz8pbErET50ewhKTsepCKXHnWSkdtZ
EANCvfMYi0ODfs9ktK8YFoNB7liU0Y1Y7FRDec6a4smYgbs2JPlrC2YsZ9JV2onj
zlpL5m4YTOP6sAydvoNcMbd+qUVNLMB2+6r+GY6vnq0Usd1Q9M9cAn8GJf6Ua0vL
2tWogxbUuTSVrXq1w30VJu1gawM3/xYozZ8F9Ihfd+W5hWkr1htgUwzH43A7lY7X
oOWsxqumSAjoQDolh48FdmrwWFQGjIxwfkPoVni61cMeHhyhbfPv0kNTpTHWdEkQ
z5aEoMj60r2c12qOiVgsFNUM5+SHR5l/cjki5+krZ9NcmeBxngmk6RwAKewyF8n2
UmUaguktf+Bp+liGpviHlFWA3/30Sp4oUq7f0KdMm1YKM2CIcGoEiNzt8nphnBRR
QDezzgy4yllUtMTfw2cumgS98XvF37IgTWmVGzndLEoi1favYVowI58R9+KviLvj
+0GJg/IY7wi6cr19LJblN/qE8dB9lnL1StTMeneSo6nPXGgukCulKwmd6XyPlGFC
QPM9/zvoSZ/ES43WVaqhJfspAnaglDLBdHQslL0PDn70XSDdC/naJd8FL32452jh
rPZQqDoZwc9epcPApef2Jdg58wN/jWhhbzgdDSTElEfaPPywdmwrZgLP7qgzxWO5
ut2swDt/RzCQfJ8Heu9to6qJOzWb3vipephIsoc2Rp56Ux3rXv5sqlfgtORaWS/Y
GmVAIJ0yYcj0lw0Z+7vjGUpH1SyJJKiEASvKpUtSHFviATmMDQ9J0HjKJdP6y3JA
hyPHwszeAJRO3JdenZKPvvEAdojjGp6NpIPQEI1mCbbOokY5YpUBqi/shUTFMC4D
wxSR1uzDmY5iYbN0O1rVhwl6m3CJgwygoWyEv+v4xZIlGwDHmmpzU7Ba0A2CE3Z9
3ghpnK9hAYiFLs/C6wDX0UT97YtkIJ+9rj7Y/FoOM4h7TLGq1YygzK5xMLcd+n02
s86N+7N8rWIGdvOi3kxFJdn3OyrosMgT9TTsU43HAC72xqbi+t1fGz2eVUaNm9mA
FXFdInQ+YLpZCcN86LBzKrL7WKV+vaRSWGRuuiVPF4ZN8rM3w+pOhT7/xPTlxjVR
jxcI9Au4c5oLeXxfE2GI1i6csTnAz7GM2Uv2N3e2Ivbq9W06FgtCTBCsSYbbohFy
AuUcrHM3JLwSYl/8Sc6WJI91+4ZHwk/nHTt7a9jX/dJbFZL3vyKCBmANNecKdtHN
rQm8logXG7QzFoKs0eUa8qRQV93i75tIlOJkphIajQOl+06RfKTJTyRvQ5a1HYvp
g/bHxNkfc3U7ee2ITZSMZZpuJnAeJqkA/Jw2Q85qHycuFygTF+vZop7n1rg5aODA
Po382jXM+VLOACzCRGVYdpdPM2KOvu2f85M1DvRCK0raOxWiMY2kZnOcCjuM8KvA
NGrlK+jUmS8y3P8hF0Y3PccLwcv5CS3ws1N2nIEBUaaLC6283738QYqjZB0cT8aK
pGXTUUBI0jlhGLPoTn60e1cjd2Rb3ZZ+XY1cZxPZVzQDTTgxCMmD7wtPpjro4P0r
5SCk55sYFFG2DJL0IEZdMzILV/5i96wY291QepxRnj95F5ZAEcmpkDTVQZ/tTbAt
JMo6BEaCYF+m6S4GJIgBoQt330ZqcAcj/eT63yvGr33SxpsB2gWm61P/z2NAdzFM
qOEkbgdaXYNHWA855y2sKrKu+v6oxStTOVhPYnHmiHUnIgbvMI4fIkyw4sVEQyRC
Eui+BEC3v2g8cAi1R5HZ5fAckY/PZMIBWkSWwXWCiKvtbiiL/B8LTPx406gjakEq
GrgJ9yvN5VwuyQLK6KEXng1ylUG9vJZQxljwB7UDdMe9fuTTYEsY/q8HXWXJK7kj
4uGmdfzj8MfaoG6xRETBATnKfF+d56do+/SsEEnT2MQAC5bvQDPRTPS3DF3LnNDc
dq1J6Nq565lzLphY0RaqrgrAw/9fmpRek47Nmky/9v6k8pEECw7s1mT5F20F/pHG
DRj4pEU2iWqwaEo8WqGo1akREOMo3NsJU6QPKdlYN5QbwcnoHbSM/CXjEWMe6whq
Mj6j6tHL/JzpKzctWOJL+iuS6i8J0SspUX6y3CkkNPJ0setyZrO6UdNMP1YGTaVb
HKL2znbYiS7TSS4zNWymSFK7PXtjlJzoynn83rB/IqS9f0e4TlDKVvXPZF19vZeL
bnR1oUtKDRz/B5rqo65Zg5khCnnyJgC/1DD/vXLZe5gx+BahrHqz+QJdRYnP/Wj4
RLCKmZRehjiiA115w6jpyjlgXdtZeyGt5pBTkG8yb76/vTYADilR0lNur5StCWLx
I9kT5RoZZlj9iuC7vJZStz39P3mqmLG+W+BKGjvcXb8d130vZKG7D54ps1Gp2FJ+
vyTTyTBjaISJC5AEkJg+Id0ewyb5eXwHEZTiyLKVF+Ys6nzTtSvJUUJFXWupV9qu
0T+AZPQKsHwdw2v3n3HGRrDfL6rVoKfKdy7H3OJo+14Thm4d4GiZRA8wUAn9v/zZ
Gu/Xbp9dtVRfZNRkIeoLh/Z2OShWrAUWJFsyoLUmNw55By5SdqHh8++9E/nAvC6s
cYgEFijYqOiI9bje1dVnl8SIAAA9GwrPIeSL/xW1HmBHe+8MhJmU/fSvAZCX/w9v
taRTjiDyRHiScxQgWRjx8fAxNNbGtr2aD5WXUa1AGGzKEZo/X9WoyhVN0b/MWMw5
PIvcnwS/+6PHPIiM59Xff+a0qWi2Ffx6a1o5vx6eyyl7AAHBpwCJreoRzS5jmanc
jK9oPYCY0X3hCr6Om9vWIvze5IBsnWJ/NvOSv2Bq07vAx+ccjSCfW2S00IRNkOkp
DduNc+62L6NxKJmRj/w+zC3enPVLyeNNPu/KjIcGTwG002tzwWrHaR/VoBmqm9/O
WXS5SxvwevjtmU+GK2AQrQ869phR9aP+onjFD1gYOQtljRZK6HDqIBxARz3d//9z
pM4PbKjf/hYTum5UQrMFyOw+yhwNoqLiKa220AyC/y7WM1ZcyQxpIo7V5gJ1WREM
u31Z2BsJrIu955mqij+ZTnHf6RK3WGVB8wLaXABUkrfRaCMNn37QThz3Vo7vwydq
KdSdJnwUwvjH+G5hbtkda0/EjFEnkSSadNxvu6vqSkYIef0Mh+4trc6Q9b912ruu
6stbOZmq3cmCkkKehskbKJVwu3Vp/Ny/cl7N4mzFntGlM9iOJxvjGD7TwTaGuG85
syHYVq0sJBcD7hCYgm1PdDUVBMNVtbqIRitxlXt+dCdjYg+PWnJO8zgOQaOuNruZ
lzdj2MlUdC1Sa7MLCK2/Ro88KUdshmkjECHjJPgPxktsCEa2HwQa1nEpDATNk9B8
Fhjw0OnhHfCluW2mVLz16jzGOUXpa/YMIot+eW1dux4rr2KGtdxVl8Scd7lJdKIY
y6EcuyYn9IAoVPgAWYqMcdiaayp9SaTDzg8kKnMvTyz7pUKfBmmzgaOc9xYL4GqK
i8SDyeKxqeUZ4lZQJVaq0BLOxURGrtDsaDujAquTpAOvenj9sKnApyNniERb0QoN
2OorgzMNrm8YZCmIm/GQoDWlRXsqH0VVi7Hl859/DEnSx2ZWOO0Dt8Lz6y/lkUup
xMq2HxzGIIQvWg9pFLpD+tEvMpubrFhsDf/4CMiR5McDKB14XNWWb5JBMYihD7lz
vSvthVE1khLgcrJuSABOSlcIU27AulAhefnuYCKaibuoXSaC9Thl9sI6SLOfMCye
EsJTiVGBBkwIuyGYtYQiy8FnkG+O7+Hjw/nSHs2FUIxW+OmMjWhF+pUH+owa3koA
j+w9O2fkRsQto0A3sg+h9MThCgvc+Gm+LQL+JXWtIx04Zx3TK5zhPfc+ZlH1r78N
VtBiNUC25jK1UKQdI+/c6/6faNQylDmbySQ3FT+KGNkpcPoUnC47czKAkyUK5wVx
iFZSol3PUNSYJzEc3EBYZkgfS5Ae3jjGPXSqgM+K5iQVr3r77c79QjIKbpjV31MC
KT2o2QFZ3LnS+8GMEEZTu7aSBo3UJ/GVMye6yruf4G3X+2m6ZvEKsZT3So1HGQ+1
z6na0zlt1L7oKwVGTK0u2Wyc85ErttmsDTOFCsNKtXiSar07C2Xd3DHakJjhLvwH
xJqayWqZ0kxk2x+ti8Pn7FvywvFm/XssVDsSl6P8Nl+kE9TuMeq3xVzCgSlafQAp
MBZODT2Y+UQ79sAuzEvz6RHl9fPYZ0Ep7Dp3jJYIb0cbTl6IFOSfmwIDUncOTun+
Nwucuq3mtW6LP01Gljl5oQKzxpE+hhtxrLR9MHeLamg0Qa/78UVo6hi8fbO9iCze
GW2ZBUJHCK3Xw7BfuaVz5RqbXgvhnHLLZT+TP/h4tLwH8UgSru9WDkfY+imKf/5P
/5hQ0YKt+WyyIzuJ7BDIfAqHGYqdYtDM+9nJI9pk5IxeahojEGl9I999O3qprqnv
Jcxqdpc6MJzeNGuZi9KGPWRUX3Gw2odQaqerr7gtyt0nf6TwE5m+w7rYKs5u6dDo
4MMh/udjt9KscmOcRm/ZKcyfTUz5+iVv6O/Pv4wRdy/C8UGJXKTSD3NMkmK3Tw9j
NJC8ikafvKMNC/Jv6UG/QIIllc/oSC06410VXXt5Ot7v3iJAqFGfagBNu5vFTrGw
r2TuCm3nYIByiuL7csipJZ5gI2knj7sJmaU2H9UCoh8X/RHyDqgBXR/q9EFXgkqP
NaXx69j8m28eAUpq9QLVuvWCFnQQiW+Yxz0Fb6ymfG4ssFeCV29nbuZzUPvrGDHw
mC4d/onxlJKAP3lG3E/ZmqQFm3SuOCNO56RWefFUsYianpkNPQcjTc5kcletc6+e
9DMGke0pfeU9ZijUPDW6YdKOxX4jFivbPLBfcqFOf1bI38DepCZsUxk9uKxsnwz8
tJfHl1+oIistN5xtU1DuJYvwGq7kTeo2kofIdzk8XJJTCOzZFPJlTjzHfDtQgui2
e3H8SoyMGdypIuvWNKwmrtj0SdaAHsob2X5u0Y95DjytNA6KlpI+YXUPX/0LgCLn
uYkbNLPFvfLtj7xj65Cc65lfJ6M75Qi4Dcds65cshnbkuN19VDMBBIasQlMbWI2C
fV01FhugmpzMzvggsJJD3bacGU3lUvtuphBHZ+oUjeLzjBcxPmsXBQaObh59Uce0
V/5CMse8ClzMJBKcD2rrQF73mLqoY/annEHs3/v8z380u6fCQennHNfw3ZexOVN5
68bo3MYBz7aqPJ1+NFsJTNZipU6Snz/S2GPQr3TiohaGEYEdYzSV3DfV8zpzGVzt
Hy1Hj4cwI4iTHriqU/+f24RymltT+GRlZ9x50ATNrickD/M7MLiHwCFhKdzVYdWS
PEFnDYgODUE/Raqy3+mCW+9rC7x/TxsibXgG4ejZ8T0bHlqzDZ2NeBGse/gKpQJI
fSomI0y8Ef4HKbJP8MKpuGLfBkE9ZYjevq3rpo/pqKBPn1dOc3c0cmkpk2qoSFzv
Ycq7orAcLhmI5vdPNdmKwzIuqVXLdR16VqaLHyvpVmBu5RvJjBcUv7hrGx40cikZ
V4sj4kQYCy6ZY5arpYvMsbqSeLEdhLH7rGw/0vbkG0KFwXf94ttG9h6nOb8JsFGL
3zgQ8QP920s2Br0arf39rfeLCYn011GOjx6HbG/aOHmZWh5neR63B8DCwU5aoyuq
yZ/aQkUXS1YzEG6PlfeCJeX96IYtDaB5zjxoZuT3cdKrDtDUtnS9g7ovFX21ibhm
DZxBz9xYVXmQHMs87UuYTbLsp/XzZxJHDR2665ERU2CtNt6wBrBCm2E8YKyWSHB3
qvIKWDcphafkXi2z+HBxoXzrUQqNrMXrmE4tj70Ew2iY1nfpvwJLV65zw8hFZWao
ji6P/EvnTFNUewDfNTnsg1KGHIqFbg159jOVucNFNU2RRQ0nQR+nWVVT1YYdc7Bl
uVaqqgSycAq//erB7DZcfvYGiL1ebd7VeG347uhHHBLoyo74d79PkBFWO2EoTzRI
DUvvoYqMwq4oiKiy7ZE6B7iq7/nmoWW4NJeKFeHzzB64SL12opXdG6VLX5fCtZJ/
TSPW8Y/tXsWTJiJ0UJAo8G0a+4VxvCAjE4wrdctO9YCy2YVWRb1FqvG7kHfMKWTE
qS6Sxlo3JgIzLy//tK6liKxNdIxZ5lmnJyvsJFHOY4Pj5AR8SD+ToO0fv5mz8kpY
2wp0WIIb89xnsh52dUpwETLbS+ztkvGmRUEomjgifLdYvyZHo+5PBML33CAvK1bT
qUjNcNvvL7MJAR2bXDmCO/dX6KjW04VGpNGnmNQZJW/5xgn+RqmoDOWCye/X7nIq
zXdpKwm7X05PR8oFgKjG4/b/hjVWC0V0cZLCr5qwCcwo8+/Uzi+AXSgKEbIE7VLA
mvxRJlvrMhEFlPcqBO/hdqMpX+dNsWckmLONlcyrmODJ13FX816MOfXJkbSS1O8P
KU30alyc+9YGUWFdjnmytZ81fLgszhV94TuE35nXYAvFw7f6m6Dr/uo3yOfoFXHd
VY2+pg6uimQ0FKb8tDB3sngmekS4ejRYXoKpF9dYTApWtHgGiE8oG3Cr9P8fIlUl
Y+AY2iHMq9p0ZK3O0BJdEWfcueiJmLrXsSmEbBis7Mf/xW74TdEATfo5Oqd8Fknv
4DYjLXjCs7KXLwfl6saa7i55ktxQ+vZg6IWo0pXeEZFn1bQyNjv4I9DHVCLKZAQH
Ap6/r3VtLTN8ZwUSmQtUjstl1XwQ7oyp9DWwbenaq79/PB+TONG/C4Tsn95ilJZz
gaQMlm+nbfZzFfov+mK4cKpnnx/b/UfvxnUHxAmfm6VXzao5AFk67SKQAEY4gZnK
1BAVbXbuAdd/f/bVxn+ZKmCG8i5O5XB16Vfq3MWHMIWAEcjNvAAMqglz+o2JWxMj
BNPVFsJ2OzkwaViZNkCTnC1EqU+qNsXiXQuMXOlr5MAZCMRFh5RZSa1b0AEvigge
hbQ1zJp/jgOFcK4aH+P748zr0VLaeqovi9FtDuqxG4xbzIfZ8gUA25U1NtCaNljl
UFjIFpFCv8AwlQUlFvwC3VEERYYJ8exkz4fFrSsGrnsyZXmB0E7Ai5uXq1xxrdC/
0yKQ0AHbk8hg44pIeZGfSHrikNP994NzfdyhDjzN4lRTbTPE0tSeJe7tXpI/1m3g
A9IAfSEm/lCh/1c0ugiGyWMDonrwgQ+CF8LRZ45f8sG++y312pvZJcOEK29yE4rx
Pk+LXMJWjz4l8OG1nxW0TJe7CfZl+ddqmAXh4LpI/a2C1wYKeo+ClnDqfUjuie2b
IaKKRxmiFIziwHjjW2uSpOdlIbwWOfcoaH/20hy6j+Rkfgy0fN1yWI/7GIa0FRW5
IAwLr2OJ7ZBceNfuKZkUsCR/ggKmOrE8/kKXWzTXz7s0cMbopAfFC4gr2VOW+xPC
EfTBmzdlSx7rP1tYUnAwV8motQABtnRIR5yanDi5+5WLLcu/74YI5RE7/jzPucOv
1pMbcT9R7JIcTdcvi+3qzHDHeWUnlJOxeZD/RuM2SkgyrQA4wOp2l4BaAxVFU0l2
VmkYe3T7/dD/+/aDMhVDNRDi0H0uGNgwq45BpF5Z6QB4UmzVRhdciAs0YNb+Ou37
/xzFGzgQDHvrmxeQpFrjBzNOpPkEA8doRoIAiqhssuOKL4DigTS7O0GbYua4gGBu
k772nU0war86O1NYgUyIAUGXocoqJUuzHPUZrWunn8NzD+QxYsomEV/xZvaEtrXa
3BiqcvL0QN7O9N6kS74ZPPNlMeuGXpA086uyQAx9ukaRLymN/Feu2/sj6v5f6HKq
cJvZ99aXFTjHgX2zxbRlsylsZTtuaNi9r1jLEB6p7gkxKU/ix+TLpv0AK9ElMN+j
hr7F9Pey92iZuVImYAIhqiIJNUSpb0ZsRi5v9jVrJrPWu4/g2agP0pLMPkXshdHW
zuMkif0p68r9uBnW635vMFqzNeThjCnV7XqA+a16cb/B4Yn3iaowIAXZNjYwoqRT
JR/9bYzoSK1vt24A33QTDYUJbnXdR7i4bed0t2ewlQUHJ1+E8qcHRaVuxSVgSEhB
Lh0Zy4sU3oZ69+bPGSg9p6Wikf7o+jWWk/Nx0aaa543Ldzvq7nJkdPupyK6+yudf
PnQ/aRiAaArFj3Poz87hILF+ZI8s5gjwk/lsapKCwLqE2V5Sc7Aq9v/d+ri/lxJB
Af66uYYWYBpsMdMYE6r7KkVADWAjkvZQWMemLgD+frUUvaRQ/g8tp2/CiF/MPf2E
dOcFiwzB1JMnZSTDGNedIQltpeUThub5G3xFslHHia9MzP0lLcwOzSjdP7oC7zq4
afhBcjbyo24U+AOqU4IEwtIOATjkAjlsQzrtCWIoJ39/G5n5/+4/SP95Rl/9ESch
23dnqgIhwW6zpjXYtIa+xYJMrWCN2lowCeNfidRoRPMy0fFJhto15GbO2qMKYfQO
RXakvSM9xaeYC+4oDOdwLWGaKw5tbn8ANrn+zQPh38vudA0TEgO8f/9Af9jy61Sa
Ucip1ALOjkZ+HIFmF2iO5XPQJZ15u49T4FkoIDdTJKds9/K4WIvR2sWRzUsr/rOZ
JxiPJV548ZKXB6W8hVLJB1zIEyJVn1T2rcUL72kGbFGpno3ggrpCsxze6CQn+YJG
bojB7U/CyZ2z7+zDbQj+O5MqSxrOCsyjq7iHexdSZ2EVbrsPNpfoAdTDJx8tXsmG
EnFropwp5U8mS6m9JWE4uAGm0Z3pw2iv30GDnPKBsp6WSlsmPB+fAcHfCiSQw+6n
91IitYZ8tImUCI3PcF44THjgiLqVMM+79Y2OGlnKx4HgZ2xKml2/hnfLshchDXad
O41A8gJO7Xp32IPDqAjr21cvRdym5unJYghG1DZ+KJ3QNLX3PiVRs+VcsArXx60D
fhAI++dR7E/Snl/xpk0OCq1hasRvDb6lXcxaFGQL0QO64KrospgnSiKUbnj5sHOe
JTByILqws8zJChImPgWCv6oay3fxRur2DrfSsGcTV0pIyEvd37uIghnSFl+fBaCk
MjSprCMyaURhjPP0YciVu3Jx8WYzL3WGmspmFxoYBgkiy6eHl3HePRkKMHPxXidG
+dJplmTXZRbAt82oT2J2JWrnh5psTykP6odB/w5gzvmCheVB1tG5w5Lm9xK+lzxK
1cmJBad/dKjTo6F0DIejzgqr+XbNQIlU5PNFkHevnp6HM6QhFzT4TE/DFRDM0K9T
0Uxar3Ftc3MqITWCD/yhrdh873iSbUl15TLN/TxsBm3aRn4d7dolKYj+EnqXQc69
s1glNb96B2yb4iG2oDSEaK1V7kPr8MMiP+AntnHmY1uf6DpPWEB/28eG3GFhmWhr
uCax2nH1tegQVX6gVhdB4nCcF9qFJkMKT7T1ORaB29AnYgGWA8Qsda9792oXy1hB
7qBVNON173Lwmbjq1QdrT1gjO6nHY2ZP1jPc5oD3KKe37q2rpL1Rdd+CDenwPyYV
uNwMoaouh5zZKB+Nqr1K2mp2PVT5nPXO/j636nQuDoPsxLbNUixViUwjnISWu3ip
23Jlnv+zdSX+wPwHlzRSVOH7JbbKNxT94+2Xc3jINqUuf/h1UkQ8mKKMnhdon9Kf
lOARP4Ji4RLRC8Fa73YvXLVBEu5fGZIk3Y4Sr2uf61QfvhKBz90VjDCsA+QWCUbf
Y2TbjoospBb9pWaJnedOtfZodz9S91lqyS087xiLbMpNvvR8ivHef2ZUOHcCCAcL
g1chDNEH2DYdHPFKRpFwvtqDMSgX82y7MxMIhS7GECVt984KJo26arwl0VOHuhIN
WketTrAx1OFbC+Z75zWh/XrHTd3ov3ehXE4xEf/dIF4CZmBVuFtUGXcNRCZxDhU0
YAzpaIHF5RiQAqS5U4gcW1jPDpRypvveXe2kZnapij+qvYBI9JwCEK2hQQ63ybsH
LXTotyKIMYFasPGKvIBtuB4D+0GdkXGIcYjg/SK/2/Y72qybpYzSvwXzP30wYojb
dFBl4jrxPlnWuFeqHLH/07PDUu8U++Dn0meiIn9ySDkohYNdDI4OWSVUgQJZjUTZ
tDj5t9+XyWLHTTqRzfN36nOsvG45irQL9VwRhW76lyHikIFB0Nj+twxkyrdguhDg
3r98nrYuBP58byozcp1rt/jTbVTW3CCHY3bfwCuezmMmZFb0J8pY6Y+4sIzQj8qz
qJRhGna854L+6fpsAdREp6zTSLitqo6ua18SE3FqFsd3nC+jPcVdP+e2p7+7bj6u
JaSqAwZJudmnV8Znltwd4QO+T59cDzGAWPfnI7hydJk7z93GUot4g3I46mHYgTLH
xu/s73i273FwSXeEvIPqlZJFx2UhqsQQKmi0hZ8U42nGBPVl1tTgmqLjEsKa+q+J
JomqldmVplTKQPkPi5oQQhoMcztuCdEcPz1dhwm2/JmIgmkWGMJoh8kR4LxeR4C8
DkjYdTDEnfd7FKtXqd0xwd01znyxhu6wYIKvuECkwk0HUokEkLHBBt/kqXckuH4s
MOCwBWB8c/0fXa1WyzWEh9V+vWN9AQ188mrhy9Pp09Z5OE2nDRYnL7kXi2r34jPt
DLa8xtqNIXjwL2U3ul657Y5sW8bjaQtah8UZngqN4+zLK/gU7AtjIKqYzeL3jtYP
RMrDtDmPMrh76UNZ0YskDHJ/l1NTg3LJajVcxB8xfrWdOaSsZgMbddowwzvn98DF
I69AwpVg2nQP5BDd+oDgadyI43Gd9mDUR9FH9hQbfJlTVwHjr7k2f6jzbJtPABRj
eWXPe6rFjmny7NRDsrJ1xTFMiLejbyM7uss40dY9g64si9hRqjS3PBQOFtCk/ckM
yIc/iGPuOO4TSl1RBs0UIxH5jN4wALzrGfMiy8M9/rOdl+RWPXecPhj6RqZGyHcY
apz+oq8brylzZeFMlkZ1gY+rHV2HSitxBeiuDpR3spS8KcJmknA9/p4jB5j0+MCK
FrOan2RWAMn+slo8vGMF1461vTbjP9En3VrlJXcdgkeAuh9iCZzu5bzVtcsh3ZGY
+dat3+u+3fzBl89FwOaLLYjqflYNvfCwZuIw90fO64iP2on8unyKdu1XipcScaZV
TJRj58SlmpvevyLcuwa2l8Xqj7leqCtgKCUArz3fpRDhke6PGl2LZKox9utzvQZ0
TBucyfIaG8EgqNj7xjejFJJ3N9KP4DzYU7GtMHrMt6BTvB6oenuzKfO/fEvVgXu7
Y9Vgr6RNUj71CjgFggSe0T5yLprxF7D7KJpNnJ4PdjaMJFJ+n9uxdW/vGaYZhhQc
kB2KZsgOHBJ7dhMNh9D1JG24npwUVUokSLNIKFSh0I869uxO2Ui3eDZTI3A5v1wZ
UNtMEcqWB9UQl1LMGAkGZuehipAjL8kFlfmpn31DvsGSL721ieaeDziO/dIrGjtY
+ISfjuaRARiAr9hj3eB/X7MfDWTkaay4iMb2QBw7kKuPvG3T62DYl6L/RQGvFNBU
3l+P0i1OtdvAjScSv+FUHsPdeU38lRQA9KkNVOMw0VD505fDYCXvWbgAaRF3bgKk
owWRMfAYfQe3sHpONWt0tg+stecbza13THkQSq9oEVMN0M1eo4WlRTfin6ANVKan
vZc8jIWgMkI2NXRuQQnCRazb8kCnC+izSLARFcgif1gyewe+cfg8p3Sg1gU9QsiT
2Lgv9LZ0v9yHVgHKcTycOn5in+vYm4jKYciVQ1FG/5SNDZl4Bd60YoYDvjBVzXmB
5PXupL4+FARM2Yab7s0R494/C+U/IayBfssTeAvJ4PzT3i3OI2xKaDjjAS+vIe+x
vtnh0Dxf6KlHmJNkQKMUhJtaq3CTWriJ5n7cN0YpaH9P+R9X54AsVAaJZEUOBGDh
AAqnOUeAS7gESCbV4wg40gPvazwAQpJElnpq+E4iCx6ApYm9rZRcwuogUKzzdEZ8
0qnlOf0mZHlj6EuYo/y9MH9AlAEG076Wp4bG2F/+L2ddxjDe28+rXTRMUy4nhVOn
bIEQDHf+2HrskKlwUGeez/Owx2uFm0MH1I3iwfUqPekLdcqV2TDbeQqYAl7yDbIa
aPatD+0+d/2Qu2uq/wxD8yXH4uFT1uDk7YgQXaAw5TUuwfUnVIM5Eh0NEgUHZxZj
SaHhhLAfmraqUdYgIiTZZZes7nCpdhWRtQxkf5D44EtiItROTCXqybECrWVII/QX
xROQw4fhkLJrN078zLjrTgZLPvwfGs03lXip+9YtAg68hk6nNGaisYTNf9m8v/nm
CgoYwAvKfwlfCb1ujY8hxPrXW1m/Rq1uFiBJYDEmUwohpw0ZjFWOTJ/Kb+wS+qSG
lIoe1L7P9Vq1XBo7rvp+xwhXHkXtCGBgMpMyjAeM104AU3n1Nv0xhZYeINJMG9B5
iaju4g5rZeC/1fO2P5mz2zvD3JBBei/Is4zdd/QqwicLrOWvYXTEzIOnWE0bG83t
F6ZzHJoH/c7do4fmGu8S+y9Nsu7DGdl44OvyKODQhb80JDTV5avG/WP4DLOuF5D7
/Q0S9mh00bXc6QXk50tsNUUlZ0Zt6FjMpfJ45iQEU0aCYqJTBF7s6qXIra73HL3m
nRw6n4QJko1E0g+/zApg49D6hlF52p+kltDnu2FqaYmLaVQAgkK9BShDIg1Av45F
JRaVjXMUaYc7JYg2YZncnxBxsdcy7+QlG4x69ZvY8UW/apFPyxAyVw27LF6ugmOA
iKzRSe48SM3MuCAGWmy/ST2PoQMYOWpKdbLHD4V1AD36ffyCwkCVvH8WrWeSw40n
eIMdXKEbKBSNv5wfxYpHeYt6Uzhgd3tKDbRCnLxq5By2LgxEUFKFd1ZJp+SZVRRf
CLYHC0ZgO8sQ8UmU35xkP/QECHhVP6doKIVRGLyuuP4T31hooiKcnVjqyzfs01MM
wbKOJCfGqV4hdfKWh4Uy/DgRSpFhtOwVp6Sp6cEjM/zI8ph8b5KKX/7U4juwQul1
COeEdD+MkoL7m5PKn9u8BJVhb0DvmM3zV645w4bEakJOZq5UZtSs7xjZyha9wh6V
Ol523f1eLRJsqlrH1/8WvHPHmyKKBNuW955zgujA+7jyH3e8qL4PGbC/RAZuzzt1
4o+B26FHm08q5K1J1ImbJqvFyN04Eyv/yXuBlwfV/krHxHLb3Wo0fIqrVablM5Oz
JdlDmw6ZBA4uIU+JmQek+gWBHWmMa753qiOXNmnqpbqBw6dKjw77hoMvVnVCgN6L
Pmt/PdGOW7f4cMIcIebQAinKqk9iWxXUjOUjSZiu9y6YAnAcUbJJ/AEeBLg71ghK
EvN1zEGMmnLW0VwEtVwu/MIpDxQIDneIR58H4vh+QZVJEo3qLhaWjcJJ2Ce+NYW6
osszD1uWMTTtgUWVwUokOc027g8EWF0tFo+Dft4WC7TKfqcBSFrSZ1q6qcMofkT3
qcJIuL5Gf1q2K1JkxvyQ2DIBSMGcTMKhdFepwVfq0oG1DvoYJNmk7GLtjz8yTypJ
QkXpdvP4rJUPOW3QZF5ISGI/Du3dR0rX3MojGosfi5C0sFZbESzHmUodBqHWpAbT
fznWaVTjaXqK6TqeFFSrQh7C/I36rr+G1T0xPOKLUfYP4McKBDMMfUnT5dVZfdwW
N7aLM1DCE7tbfndsi2mGYwv2UdnjhGVeLP22On4jnajMVYaF3pCPv7GIRtl+wThR
ZbrAa3TYC/27/QQdyPyX81pJ2dylSwUGD1PdDq2bRfXtbcCypXZZXsxurLHYwPSW
ox9ZVfmvPNZ2NE6QvjKjwhStVDp98C6rDQo0OIUW6nvF69sTCm7othTg+C7v9Qv/
UWrf22O1pksYVRfzTgAr+rQhoHTp0RBwr6KUc8M+JZeEWn34NfGVuUAn4hRysRJg
eysIHfGE4Q2eSZvVpUCsYqBKmV3YdmWPIt1P/2GVFgBau3bQRNd+LPGklskmUxlT
dp8gu/NQ1bo2+XANmZAND6fF23RWlqc1+Xak2r6tLfeQsT2tUNd5Xx9NFmGnVY/2
NEjE5amphRdP52662on7j43k7miRsOa2iodMMvwM3yaZHSc9VkxSDbk+QYzSxfCG
xnXq2K1Fdejz8bl48LSLH8nWmpJ1ScOmSuKVusVBtnN26srHPikNIUyMsPBqYnJs
UkJNyBbhidnPeSl29gufImbA3wqDsdnrmLJNQyVfXV7zjJRfdxmoYcdM8oNNKp2O
Mt6Nb02u3waHfSB8rzQJQvh52Qj2W5dMWh6y+Zl79JZLxvlt2SJx/qAnDXKF6hbt
OJMxfny96dcYXDMywLdOh9f4FKAW8tjr/QygS0S89t20PjXLUsRNEiyHOoav723O
F1m+N2+q/v0OpBls9IqpScVVbfi0chlDNaMuz3+YIOVeCD4Mjr4hk2jpSsN5iASI
QquzN4wbpgzg9/Dem6VPnD7br7Ml6j3iWuq0gFpTdfIGCW34AvKZyp7fQwy7omIo
X9PNJsZITTViB0kbOc2jIj4544Kd2rexvkjuIMy5Y0umBoTtUEo4ZD9rGY4f2rcJ
Zrq+hwtXSnRhyLLaaDpIA8XTvmBLDG3fYYhzFSRskNvd5MmgtyEPa3n/BeqiT5UK
X8XhDI+IHEGMpcb/aXYnDimKWepSF7jojoSXl7S9j1Rj20TvNqcrP5S7k90fPnLd
9w4vBGjBY1Ln8+XIWD8utCvCP4Oubcut7k/1WOSpUNZKsy09Qc5jdUBlYH0x2H8h
+Ur4tQIffrAe/VaG9VvvO0SS9LNqTNN9rFBymRJfOZ23LES7K5kUThGlrTliEtSE
1Ju2QD3BoZFc1Fc84sXUArSBmAxEYPidXMRZBFf/psNeZzL7Ju9PwG38I7vW3KxF
L7tfzCZkHUmmGmem+zS47Zrd/nlPMli+qmU82A60OORODiEOemXlJXFUocHSCYLu
ZrnZILZ5mx1yCCUaGHB1vDAS+R6Qfro8G9y/RFYo6O0zgSN9TaiM7zSyLwlkMFMU
AGiTwHbb4vQmSgq6u1H1svSVqMVaKIhtZaSho52YQLZDicv3kgyerUe24BqUiYz5
30iVQ7DgSsP0E/m0fXP7DnJSnVDnr4Gu31Ka2BYBtCpa/pSxF9SJsdVLoPW1kwcE
6x+HDDB6zNaebUrh7HwOCYD30sQDtkw2fnlgCAR73yEw5FVutm2/2nUaDYMRYwFa
PbXAFG1FYdZ/9DqGvz6dfGw5e1avZAaX19uJ1MMVsqJKcVsHo7F0P4FT00u6/0AT
uE9oAM7Q5AvJQbzNYO7c+t7ju7QSfaNYhC2SVxJYt+b3DePf9QMubOaWHfgB0F8Q
jXAz4Fs2Wc0MKI4o3zwdKr9+G8Y5j8B6tS70njLk04NTqkNAet/40p4NkQDfkb4H
SzoocB36fPkLR3YUscbrfe571eM2dTGC2PSXfDbdw2MHcqjR12HtQjDllH5alDI6
wTRllCpsr/uwdzkvlpg5lGgXKsJ4WzHvNaHxqwVN+pB0CXUdFKKkECwfaF9kyVnT
Z8t0Si/6PwQ7+WuWnTAgEZp68bbEDiv+g3+3Ionygdw2rJndLyfOXthHAzpuMxA4
LhKoCENVDEupUEvB5qPiI9L+nb18W+f5UF0+MQEc1dbYlbbDg/yhxB4a/yS8PEWo
ksDonrHb3haGVBIGjnNw4t+WnnakaOU3PpSS4gD6VQk8rEVa0aaCRno1YZp66zju
zq8BdFoMBkPNMOIUU8T5tKYK8xIpr2kWZzZ1QqlOxLDPkyNxwn2u9B9yBAhiMoII
/hHS5Ij/yMSnDihKYDlCFlRLtJSgLy0bvRtnXiSrOUE4kpZJuiz25nm/QM+tFACg
tbhdcXju2QGbqufx7FWHQ86+Sm/9AYCBNZzaL2/g9Wx51ifZO2nwB/dRb3ZaZrr1
GopXQdaCecn0mNyae08muiU+R4/ytHvoyOP8NFmKdVMjlj0+h4WB+aLLFJFCpeV/
GtjQPet1Kp5R+fUyDTvGfJhCcYVtv+Ild0GHOjm6oXZETTvTfEHKG7H48YJoIxSr
/LpEbXIOJZpK9kDc2QGhcp1o/djhCXwaxUzpGDoW+nYIsCivYm5FjMsETlrWmZ8g
lbR6hEoujNVK1UpsR3KVIZH6o4cG2IGUSILt8eQTPukL0p0/SN078FfWgMwk8GBd
BnL8egfV67IdJ3bTQ3tqlLA8CveoAz0NleGtGhGJNN5wAK1ndgVYP8jHbm5m+z5f
0OSm+50uidtLg4N9BfPSVQZNFxLJKhVRRuSPkih4iuQT96T5YSQJ99Z1zQkq80dp
/2lDpd0ZW8YCt4hu+1/Zm/kzSUbA49l8Soh/nCKIjKZaVpj/t9SzSHtIZIT3oVeb
6N20o6OeZ4D6/ceymHIFqIXDjP+fi8xIP0L8teN0IJrkpzufAHLMoKkbfVNy0aTH
xnIdx+SAQz074Zrt1HSxPhHY6HX3uXwt6J79g273VytiLCGHdXClg7hycBTUDv34
f3Zs7M10LwacraucH0XVMeYZznRlBahfkPCyhQEA7bDSqw4K60yqNwq17+3IamTs
gYF4hb+L53rxbAyoywP6bDI/b+/CXWhfK/5MrR4hAxBrBt1RVV56BUlAK/y7wt2p
gU+jUC5lS6ksJY0ssmIyW5NNTt7lSRj3H26srfczYkEh6QPP0j/qdmnQyMnh8JcP
HWENbodBvai5CbGTY2LGCIEHyyKttcU5/WBpzk9KAPHO/ZO27IVDfyigUQSl5s4w
x6IaJKzyACU0BL5mt/z5mMKsyByTBJDPW0Weoy2AsfpBszn75T3daMVBx97LCfJ4
3jDacGU6AhRyWDf4tmSiGrFn9zZPLNHnaoaBMNtxG09yY96mO2vf/b31eiMERSQ0
yj4sCCljVvSTMIkf1gA2JPGgZnTuJUH5M+thfLsXp6PCS6GXJC/iAkyyRw8Y1qQZ
Ev1Dl3k/EVDMAPEuu0zHbLCNzUEb5dGgKUpZ4mCwXqViqf6WKkTgshEEFbmmbUse
Am1B0vt8PH0VuS4b8NJciLwVWPnPBu/RR2hjhCL5S1FduCrR/OXAJXlLHzl2vFiN
P90tebrAEEDHUJQLQSOHN21hLzNWGlazwkm/GcCe/asih17jRZwBuE5jG1MvvrbX
Amro9V9DBYIgziX+1GGZsBIdziSzEbdVSOepdxCxZhhxFE70aNpAS+Ea7LuPLhCk
twEud4CB91bf3iYhCxZ9dTuVw1SyqzqiraHRYoTlNihIpb5gdD4kf1s5Y/YnPA3X
uoSGGiCG8lD0/jmSIoKAC5TeVn6dN5QEKov1aRJi2KpKWfyS60MnlADotGI/CDLn
A/7ZqguBSb4MsoW5N4h4nHWtMVHgbFyNXgqh4PIEzMTOyPVmSnAdlB+i98ujduAx
OzsdrWIyL7lMT4ECxxROi8V0z2OwtzsWh78tQ1ZXZ0tEMHg6QT/zB+HK94zN9EJT
+leus/fhon03rZxFKTLVpS4bw4eiWDTFdtq0/aDaawPtk//q0Udi7x078Ew62BpL
1CNpzVECZ7EqOKDB4Q0nHIzB4yw6jqqs/HTZrUMGkIFZbAoVsQcANxMvErhChnRc
6THKh82rvXgP6hSC/u62YaLcl9W4jjhGJiyYiSPa+M/j5ZHdWw79osBa9WyxPp5G
oT9FkOrPRUxPrjbhQmeH0qXxPIVEqffh7r5AfvYUoZY1RhOTlPzKpVs80NWm4ynu
XfwRLvVPun1wFuucy2G0a35nDRqiKvzz2g7smgjqxf6IukAiglr3SRAr6nGTyHAI
HYPLnJ9DU7NvdaUh3Eb4j1QBZgwx7xzLOJCxZlRiWdlW+dOu1d3549DdCglSK09P
7jBZKiGJOqmp2jyJvCvj9keHmtoi0HUQXsBIkCAF1v1KeW4rZMLyyYWAjjaW1sym
K8mhrGSOrsNoJfiu4RpIOldase9GpHRlKujTyUt4TFb73Equ9rWJkoIYZgww+7Ni
PCrlDJ/pk/0nIooibVIENME3ROsozlZONZFPs0cf6M36IDU6WT1Psom035tHMEoJ
b4iV2ze7lUENLlddAyzcRGSvRiYiXlHG+dv9ztr+lS8pjscLMT+V7v7C2q/mRcQi
EUT2Wc6WL2u4y00MRpWEcaWA4bp20M9/WkNieIMZhFQ5zV7YwhJmsDD2nFDf2qNr
Yy52QmcPk5zt5Uuz1q8HdPk8TSge3/s+/AQiqgVWkI+mO5NH03y9Z9W2gg9Lu0zs
oolkKsvOvzVSFhmSjef2Lf6URBnsIyA7qghF93OnFIZMhshT+k+hr5ORtiuVCoqz
TS4+zCn2ueOcVJM3yrbwl3bcX/TlB4dY+lJUCIz3i9eQN7gc+FohU4H6ZFNzKsun
YWYRhLqDw3nOAiOod+sk+hRXrzYOmpP4qYFewEn442HuuVcIzPhV+nEHTLJeLQQG
7bi7dHeqp4IDzweX/62r6QF4WrYZq5grA0m6Wd1PpuBBMGQAgnXpfFnCWbMM9q9A
BXzansd69JdcYae9n7QzNlF2ykBAtOKXRVEYRZDsd6933GcuUXFtSXgbJXCLAB1O
vDYmlR548IxWPtBWqxJW/xYT1NihFK7Y3ggdDy7gf+VsW+eUvbmlWBu7J0NsZYKH
ghx49PG3gPsU53d4p5sfDKtBPe+ejgu21p/GAN+LsDSDRnS5DlVzhgnjClDgmC10
ov+Oc0byEHmlQel37tET9A1uYDNpC5rvqOb/S6INTtset1cV0C7Iq1rHpELa3Ui4
neFl/CkFuIiD0s3FWnFHiNR/xzxqbLrI45viEMTdEFu4xBfsORY59+sL9hDy5m02
h6hmPWVFxJ8fDKjog1WBmcbPHDwrr1N7B1IXn2HAaSZZqmtk/OZuhyWQghZm1wPQ
Ma/+kPvgt0F7pYhztu/96h7WF1S6yZtYeA7BjHrbc76du+UHzg8JDSsXMR+amkYc
llx82vAdMezzyuk4EaNbWceVsYPcvb8yztOeqfiXKzznW0Ic7Y11WOblZ9lX4HOX
CA5gabhbRApiqdqWJ3kjOJJFzJvCr6v4+2ApZMh2JtgYIDdpbZJft+NWZ4oS9L6g
z6PgcEs5BRVrngInJeE4Ej+1n706ZSTUV/Q6n3vl92qvKezJqli9iuJL39TSE87w
A8PSJAiJRnib5zmGJVYXYbWDHHErPWTsfdd4KxjV1BJcfnPE6DJQg2gmrrlFrfGD
dBYeFXVTl5NBPXZUtkJdNH+rj/kI1A3vPGXKEj6mFJTsLP1KQ0cZnobqaAAkjcC8
7P83WtxRv8RvB3PZWFC/gEIZDV8ks3ZH0IScKm8/chnf0nZoJ5v5+pxlVwgj+uqh
rA5iCIdT67LyY8gLr5TC2ZEN7lb5UO/PY/ePi1ukpRh5nko017uldoV0qopnDsOL
3bX5CiIiLYtTV6UJbz+nV6/VI8KilqR12/XHHqDgU8E2f0LzbIVbjY3oLjjjab2S
eqacO6YC+NtOjmpItNLVHQWiiEqNR4d3/gXAg19qKf+Zl+vo+Gcvv2X4jGidjCIp
fmCuGpdGNDfEKTPW59b1QsTRRyVgKhlPs7b3D20PNCya6ufwT3Eb88lbgN/+d78u
p/Ph78Q5MOCuvLhcTBAGN6osy7ZfVl6EOw4bduJftWcVOAhFSUtqO/NwgaU8LhQ4
FY3cNZFE66FAkPbZBTlXb5yMH7V1jjDL5gPcVQizhoPOrHuzsAMj6V2DuJfT6crW
JkVcoRnf5LRfbzLPAiJBBLkzuSoMXReycnaasrRM5/pr5Bk+lhnU1ujzuApUnRof
pJ8NLrguYapJArxMFbju51tODdIMHg7ABOYhK0jmJuoHKmOccY4Gc9jTfMhHZvvP
fUkB32yB2C7/NPZJ6CrbxoOGJ6sIjUVeH8pV34h+0fqsLF9fgHk8i9sycMETsB2N
zPKV0BSHUlwBdqi+8TuIjv3+pupINWYudYbvXzXWK8oVfcTAIDg9LYskJ1nVjVYX
xYhxQq3p3jlFr7rtiefdPshRriayAVHLeBacAkgMmrYu94Sg8dHo/R0HlkbXG2W6
RQu/P7wfi+8frKY+JxbCXFYPNW7ahw8eBEFevdc1tWOglG3c2vuofDhPNs+PuEyF
cMBa9tP4eCgf0QaIFnRYrpW7q2umQMckOu6+TBNcxgD44xvcOty27mFgtdetucL6
Yq/tY2eU9kSXedybMrPqttr/iMpezbWz/23fr1sRb/V4RRJ9Hokvu0h6/OCvTShC
cs2GfJJ+4I9ECZsnTVSys4gp11xIsIo/mFmwaQe9jo4l8YlVkjqNcKlIWwfvFF52
rXnvBMkuz5xwEciOMtioz2mWJeo0Vz4N1bsIhj/5D/+cvtW7CodhC0srMoW8mPsy
t+tA8L0a4cJfXmjHOAd4yxFcGet2kmLefe1dVragd/LyhkDawDwcTEYv8wz2eovQ
brLQlA4eBChCqCg6qQaiUlbY/q3zCJ2T3kxPi2yu/M1fctKstG0qzNp94kon9BkI
AlaDXqZARnlTcov3SbeVZwtVFCXD3cq+kyG3JowbMGbGKozfZ8b7BXgbsr+EVgQK
243CnConZc7z6JeXeHTrRPvXunDT5gbYu2C/s/xYfm/okRdDobR0Voo898Dlluu4
9seCnHGU0FbvlPNvesupZmk3ZQ5nf59pyEPN7nJrJrA17UKJ2YPOyOQT8HiQCP07
B9OL/joRI3eesKNTxum2/ZcX6MDYxjsfa/634pRlynla05iiJ7zuh1bXD1670T5i
fHEpMIPO60fi8Sy8FGTE2NX5aztFWs5l+EXLCBEaWyUoCJ2BmQ10dxY3TJop8n79
K+ct/WtbeXUQokTGCqF7GRnhh7FTZKC8ELBNowwkGHuvv1zo+CSB4mzPQw8JDhMz
aA0N33+1rM6auR2GCCXJ9gEJ9WB/MnC5y0yBpZZyE2sl7p0o2Bbjx4hJVVB06PJ/
WuOoIbEJuD6kcGpRXxWpXUu6JE/jmXLQ1Y9ZNyVq69dX6xwhHrZHbe680+4cx/3v
fmNdr8dCHOKZI2vdyvi4pI6Ip3AhO99138IBg6vF44Xeb0yhqCWljCrBb8KMFCgV
GYVzOMGzl4gOBdZca82370frob9lmJsGNn6XyyFRMLR86wMxpnKshp1oBJFPargP
l06Dx7V2dfdeVM0BYofGZ57/iM2Rsqo73IYMsbmhcswdJVMs5yyQrq0CPHOnHo+G
B1t97Jps5ql7191SPGlw9T5l2iKIauofTR0212vpFpDZe4BbJ0Zsks5HDWDe1iPU
L1akmMijUCB7iT+QloNzgfMkXVkWx+Y1Xp+bN0fzxffCH3nrDEX9ov+TVeTikL78
+F9RRcKY/R7yyZ1cTSU2p5/ueRi4nASuOLgj9ihpzYLxAZnz+xph/7Mhj/+KQ7nu
6iMg3AOfFHpOpOkFTxnOUhA/Q17KiT2MG8Yzv4qQzgAO7VHO4HJiahIDZrjRYZLF
XoAqRjPBXfSLgwzlUEKfe5iRNxCy2tCDmzL6zKGgyi6hYroSIROFEMqpRuDR2HEU
Hw8575dCToymmOMyLC6lkbtzfybzUCA9IP5nFtCbPoOaLN6heYYm2qyOYANr3Xw5
cFcEqfWOzW2zlsGnBt1npAzojFqInKAMgeWyDeDYryKg6UNlfPE8kO+J11ftNWUF
4JvVpNAOT5JHHh/lp8JA0cHU32TMT1p+v0128CeZKoAUlIJMgBXN5fiiWPN3mfuj
zA3ua5/FpCucsGSYjeYOSQWPNsPX4TXV1/bCuM3uFhXQTRcJzZ54jG8NU8dsPY66
qj8G0M5qbRq3ZUXPCSih4yr2AzWMWndpfr+N1aVenBjH0dlaC59si2a5SS5aiKhD
surXDxKfOkPc3P0Jd9OhuJ5H+YKjN6RqIMvRjP/i7x9Kz9hswc7JNluabdlnEAKI
VE+7b721IL4X2X4TMCr+damSF/s61JxczmjwqcrQV+lSZHRyP1pOK3AzlZTfi2L+
44KAIYOhkXoLUnIApc6eOBmyC4QCTqziYiPuh/ZnI65w/bb4GmVqMAWfsWaaUmwe
6qIuWd0BekkH6riNbPBkQtJTIj1lm97d2ZyKYO06m5Er6GHtTzcyxyocgJMMfE1E
1sg5vTJHIZdPuyfwEj2jqeh4ruM19Cf5oUNv1JqLN2lvXs/selBXn4oA4ad1FsTd
P0CJ8kTpPl61GFTQwCZo2zV/RXCJisq0y5jUT+0pijhScKKmJ7gpxmMfeiODbYxj
y4wGd2+0WDQqpO++EADQwLdvNQkucJXIWdWOz0s46szU8ynONdyCmQNAUXTVwuIb
I01XQkWrPYKqEjlP106FfKRZJ5FPEx4jEyeQOesDdlYQTs+4V+14hL42CsCK8FTj
bnv5GDQ3ByEjD9UGohG5mwqhR5/JK42Ba1NBsp/JF+6fcM3wMuCAGa911abgErGW
sLJ6AKiCcOIW9US1IQd6w4E4uopNImrCIwxA3UsAYP3dzVt/IrtT7B3Jy2XpgvrB
bQVElvA2JynkDtOtSnDmf0JGJJJoNQosyAVGjeq19UjFkLPtzDnJiRlR3HcmKyHj
vxjxFoaUJJWq8QEgTPXQuihMcbXDnnbA6eZnhN0zuedz37wWbdtkMYoYacUpUGCw
qlJrhgT2HXCb/mePHfD2JWhYosAkLmuxaJ+7RXuRwZTpsQCObJJFmPC2RNIGCprh
2FhY+c7Y2o2915fQf2ExGYPdvVW41B0iwH4HM5NcwSdmzu4NMePa3I+vEDopZQZC
TcT1nISeFQlcD3tBChkYbsVM2588HLioyiZNvK4Jhub+LOb8ETENWg3cafHBJbn7
ryH4SkHpnu1/mBKHIMklsFouYfLSmx7WNDbsotIuenUq6E2rrz3TAxcYF6I6MDfO
8Cr56kuZd9Jc6JeGSJXOuvyoFJqviQnOwM70X7ZTGInZ868ruKZBAEOitxs+c4u5
fEHIlHqcjCZ/7nzBlZ9HlNHSZgogWbMKLWUuhhWQNdX/GLqub7aoCl+waW41KpB3
8xKdYpyWtsJVl0ZaRMTeSrsNW5cURxURIW11lKB7m8+Rx3tkiZOwg3OSPpmSbaqa
JjGdwvBqNQUpA1IHGfjyBgSp7ts4o9dWBE8Mb8P0e5ehCJ6LwXVfySiVG8CLMiSu
JwwsYYswtG0k9Zl/44nRXqg2uqIe52i/q4s8MXd8/n7ENK35EEFmubfaladgMQAj
jXbosiHccXzgpkw5D92aeK635wmlGcQbEOFV7liZMjuljzDpSnzoeMuiGNNeqFlk
uyARpP/YAf6h5rSLja9mbSHSo0fqHXH/Gt5GKbR//wn52oK52hCorrvrpwLgnEjs
YefrFpECGL6h+H9eLkK19ZK5yjwznnhcwS2o6PQO4rUzqIHsQvR7OaNM0tR0liPG
LcSIVannQMPlADG0UUAvybcWlsDUUuD5LrCgk7tspIuBZV5TBmwQCdujlP2TDJEr
gDFRhM7oZhkfg5CksgTfxuNn3KI6Gablkns6zHAUvXT0pQMomIVnDa0DdpGGSH0h
cSikgOUWcqN0cJ1c1pHci2D+plkj7kLQgx8tBwWMq/F6YbNkXk/ZVTX+OzAlc9Aa
GvMpGQtwPf9st20QumikoMsB4riziHwYGZB4gDKID/xsbqjn/qdaUv0L/wY3CqCG
EIwcNuWO/h6KO5GpEBwJXklWqvSXQ6ZTyvk6eFjSCd4yce1t1880lH8mm6/jztNQ
dwpao9yxDHmlMol4IUOJTDcMMvINPyZctOD5t95vQwQkmvL8JJRrqQy9hpPlpZ0L
5LQZh8Xa6NYkA6hnuSOErOXz6vz4BUnvpRHMzkiEYUyYdMyUO17TeG2In4Cs6+vA
R86JeowfHXVtWrib1y07nuh3h86oBaoekSBsDqhOJZJEHp66a33+gcQJxl1aKmJ6
netr5PjnPYs6dbYXPFwPZlyA2FX9Kmt3vfSFCzMq+tdcsVh/fFazWxmYIRqy2LYD
cWvhKeH/B4Rx7QELO05kKG3pZcPV+vhTxhO1DA8Bk2+vq26pmjbAd2U2DcEnIDYO
6gf05NoeDEJmj8b0hHemDKox0hQds6bJMFpnOBPAJyhhYDr3/83D7KZ1N9vJsP0J
FJOlf2Q2QzpuFnRmQWhcGya9hjEY0wSBFpRaQDquMk0DMOqutPxYcpxjw4o7uGI0
X13is9JTT5GkxSEMh7BR84vl9uwlmXGMvBaZi9CqadLELIpiyJ/EySX55zf0n9YC
tRDzMS2B/YOBJeib68Uhpw2NvhXcSh9KQ4+LZM74PEDaai6spAhy5Z63Yrx2am0i
5NBZ4QaFmqlMZ1tK+/LGMEa5kH0QPOnl0g+GADV+iivKlQ4rjGYlRzc6IG3oR2ZV
AET7iM5Ife4w/zcwuQBsBiNEsz61GqzTste520mREeISF+3+mz5hvxUhbmiihjVn
uj1mruAlGFsx8ml+5oUWuZHudrtqt3nqXqM+gjYFdTe/HJsejZO4+F0Z5qjLtWO5
L3Ntlapi3SuxlSpRIyaTIwyda2Vc66HxVXsiHmaHnynnbbjSZCX7hjgX4iz/klIP
UMFIYQUMUu/FaLvv9MypQQ1rlj/3bI/biD0zYfOTgAnXqIIug3LcWHsRcmNEdu77
3RLmhykS1TJjnFZhP4RMNVsVUb0OfFc6Z5aDf4v2JUqFWbXHWBRZFsms/wn8w9yF
TlxSUYLpdfWv/jjsIJ2gXzUl9xndyV3KtDaKiKR9kRS4q+FDEVlbEchoWycpRSBr
XCYtFcboNKrkn6TQM0ySDBJPO22Lb4x+ykr1LLRNF/OkkByLq7xDJgmRnWtMIRaB
mxMH0UtjCQpPOgqDfnIGcytnBrCaET398rQwWijeaw4U2ymt1od9lOzL0GoMRKiz
PUA7OHt3T2SpLecRsdCBvDnq4/AhEzgtsRbz52A5PYTY6Wu61raaPCf31EsG6UbI
507JYPEftFXYCtCX1tWZjG1MaMobMvzVn9m/RdBT7FHZ2H3uAJxfvu9FtgTMsC+d
hjpjkmCPSML65VsBb0BrsMss5Xcg4ShLPFVFEGUfo/JLOEBPVcn6BWIKOyQEYCGJ
rxASkQ4Etk6uv4N5RMzoBFPeztvbNWR6qDZOjbXc/7UQNNj+2Xo3TbuXCJ8fgh4b
l2vU+8MnDmUQB4EjTHRMe52H5mTV7JzpoAaQsRmjHS9Yse8k00fHZDtKTUiweous
lKQmJiJXzv5imcOrXmt5GjmZiTt4GkdsmF3cQhMd1wmlQIMC5QR5qc7IdleetOiZ
MHx3RnLAsaFzOZvOLptAPbClOwUU4CVEC2uD+8ZcW6MbRhY0mBqxEGGuw8TR8FKo
JjAzAQIplXM45Efsv7tr+lLf5CQuMm2CD7Nq5e3y7bJl3feizTzAJ+t5MKSrGJkV
kbBiLKCkJT5lCtAI+XlJSVeMsQxenippiwjU3pwJqcEl3P3yN2p6k4vQFhmIFnVE
0mGcf42xbz8n4AK0rRCsBzS+8Y9uN/IEdXunT6q3DCOr5jOTbToDi2+XMn/K+/b2
PoJu3vxdK1gr9BruLNljJZ667kvkLX03GbtXUkMAZXmBH+3kLy6UL4r4JyeEQVny
K1vvKmdrjem8tRbEQVv71jyIvNQ0ofBG2X1tooGEsvRTU7TujX1/iYW5tM5tB9k0
2nx5zirbTbx7TxH4BzPlKRmZ+qNa3FV0FRccnYBacUpEloADLrypYElIhroHzbrS
yW1rKXqbwj/d/p3/NLEGYT0fQkteyaOZse3QqRvyzssPOyZSLmjcPH1fKCpKGYBt
LFcW5RSJt0VEmQRM6EQOkcgn+9iLl1eU9iQswSI9SJeYpC5Y27+8OUQAIR6dt+A4
tOHNZJfKW57vTXkqScI+JKDoPkOx7q9tDtulb7gWAoBmm2pLRFg5udPEOwb5jyvO
oUtqP7TcZYN72jaVbDusaz87OB3m5PRcVfw6ZC5cuXR2AOd5YlsvxWc/iFzDRP2W
rze58MP0dOCMzv46wW+Qq+KEwI+ghfwRrBu1ZFVGA8pgmusiDDLOD+YiBbXOaiT4
fq4I2tqykhkVk79pBWE0eI2lx/x5kZtvKmBbybnt17PMhdcvrpOprzHUlVA6uFnE
qom2UeZvXvHQcs7vkjKeqhaVcld4bWW9umoBmWzsNuOXwV/RYIopiPx/qK4VSZ4i
LRKU5Cw7NYSmzJAGYJ7TwhVRsRi1dgE5Ibpv8DEiDfLEMAacyuySpgeajj+Z7KeV
58AmJ2Q1ODM4LMc9yagOJo0hSX64S3zNsvTiheTG0D55jmXe92mMUcug8Hahv2UD
p+DuH5z75gFfNmeusVXydThwbAuwt4bSJ8s7w571iBDGofCRlqbbI2/FKXavMCEe
NnDFYpr9xLR4vqmGzKcI67EB4Gyu7s+dpvFD1lEz3DmN4xmoWtD9kkDWJs+ClBTD
tdC3ihYX3jedgiqprHsUBt2VN+eC38h11IAMm1KTcd/dCItFj96E0nFR2x7xlWnH
Nt2qRwHfkVg/Nl3Xdiru3nYmfXY2L8DzgDaHwf1eDH2OaIY/zkk7nCJaAjtGHw9a
kM7/O7QTDNvK1m3I744yb3wKvAAjdlcUlhWKq5p4sH1ctAKhPw9C78s1z5Z0CZ+V
N2sbXDFgNtuTBMvMQwbV0/LiQ0ccKLxRHT79tHzZgtsIkkGXFY73+OgT6tlQLPYb
Vzaop9Lc3H7eN9DN1VpAGdlbxc8wDWdT6b5T8xi1hemk3HX07dTjvdbc7zlZPWEd
KFFIcRugHjCKX5kL/Xvydc/rI1UL35KVaYza0jQ1MZdF6kPkvgZ+t+rtJsFnIkLY
8PMtevKemHz4NUs+5lnMxLg6tUWK4Lvt+TGUH7uoscNCRkcgyR8XPTKccCaXY8hF
C4SAla6djMyRcr0bUfDSA8bWyrd0TqMfJj9iWY+oAd5GbQ/1Kr1GL55hXlrfENC/
wRYL+0XgrJUuC822D8okSDl7fjjNGPoS8Vea6w8LNFBK82Q28hAdauIZbfwbeuRP
JqVOyrfwXciGQaERFCsNfwaUG0NIueuiDD01XuOv0h3uaghHBXXR3m7lXHB7WS0k
ljHYA3cQPVk3wK6Puipzt2PI47406hFNOAA+IGCC7HCx2UQXZPRJzpI7QTu6RQSF
6BVyy4Y6OZqTm+upEhzlQJh5OEqo4frW+XszY45jlB7MU8w1+y4lTp5Ng4pGoBxF
F8dQSyR12Wl5XNuaSqlIa0ywf8TUbr741/RFbF47rpGK7hi2+UCuUypO8MnHGFVi
HVzNfkTVDpCIqM/fXoL4iNghpn0ACJrpawHGqT75QWJcLzqGVQWIZU+YRYKm/rlE
bhNUpe+SUttgLJjn7zH4M8IolxdUN0gAd8d6CGDHwH2JXRIOuqMCKuhTSOT07jxf
48JhMSQveNAvedDz4JN9Rs5ywDL0ejoKFutrJWjhaT65RU8H6ZsidydyQRFkw/Pz
65P6BQ2pSkBJPM4H/2b7sBQm/oZUqjsrOxEeslh2SSn4NB9fEoMC+qWimZlxsQwJ
9R0r6xsNp0N+JxcmyKX3x7sxwFo48c9RY3WvFq7chPevhfp7ks8DJ2gKoauRit8k
WT/eyKLUCWWDJUsISBXmX5kcwrIuBjEG2/wpOh1HFAOYOmFRdRp5oe9TQ5RbmBhh
Alwury+TZxp5fQJ7zGlFzIulN5CGPv1FBmOuPKRRrpbSXD072kJAgrWPQ79f+uCw
6Hv5HdI0pB+QBzTElBc1pP9K5yY3Vf8GFbkjqzpH1XEl9uW40mP/1v4iFj1eD9l1
qAEe5dMit+Na1K4arcl5B1VeP+5S8b6bzYMk0dXWBkzv3bG+9MRz7zCwHSi4xjuT
BiG2/5jXxO3KLlTmSbmp2X8wSkIN7bD10IiocSgzmSPbmNsoTB/5bRS23EQVUezL
t5+Ph8yRcHQR8xIrB7eqYtjlotIvrxfAo86c6IK3RP2gA80PulN30Qg8iLIU2xpY
/FJ8L7NaJA2AG2I7rcEFhITGi3dXkVlndmNzvw6ZQrOgIpkb5BWoR0WUAX24v2hH
vSABd2Kpl1ZOjoW9i5rZ0yZanGstGVIU0CWaJHtlhzQeXZU2jzft52dsOJQ2ULqT
PBaCLQ1LK6Lj0zY2AkmwBjBpM47Ugi+mwCEaKNZQoni7J+5sNStOF8xnF7lb/1jT
HQPjpm6vVX+XhjEV+awW9wBNsNM3PCW0nuAosTQU2WNn5AYDR/PK0nHzDPKvX6Zs
RwtRfqqHNFkzA6cwLFej6OhGolPNSQWaut4ThcPJWadbRSLnr87OBSK85x2tcaw1
a30UZO+QTiFUUAAMaiEnSoPC2eoH7DjxvuqKmjQ95Wvb0SFuzntpDNCfoUDIDr3d
iGAfkrR35pFs7KkxnoG4auPn4Ur51XSGLVUJDTyEC+ers/9GzzvFeGNjpnmDGIkC
mqlsNpsKQzJLKzmFzTl9Imh91hlEFHCK2r1aWcMOnDUQDMwphKsRzbh8FZ21esyZ
ggh0HxVuNvcn+QuC721k83LGmZXJ977FGla4Oi79R/tiy2sP7PDIwXsBkwRj4Kkg
57qX67KK2oLXnZcJmpL+JWBN92SS7XI+WZfundefjE8GaomxxDgmr7l/YOLXasm9
0Jwv2XeYLuu+WW9LCnsXz6T0bjdAa/kITsBeZxbYD8pXFy/cVEsYWaRn3AuPuk10
sX3qa34itqOB6/Gb3BJODZHXGNWxoqUFXD1p6he7La9oiW89xYo6uwJb/ywhCT/O
0BDNcxOP8J3/VD1hWyn8HErIvbb6p+CT6aCijtBlObXTorDveHGypHsZenDrFQqm
DnDG6dqogW8tBEp/ISeHCi6D2PBH6XcKK2aeSSZlgFo+xugngVMd8HD/eyFRKyXD
OrayM6VvIM06fSxVcS8nmigWYymbB8Gz/nKqYxdR9UvwpGJ3GBn/63FQDNtANCCK
Zs/ap/796lBaacA+DINZ+2vTBvkDXdHvIbkY2da9/it55ilR/pJTwrAZ2feTLgzZ
rNaMv0k34Htu6ptn5aIYy8Ve/ZFcdYKvvpEghoc/tkDJxEUmtefoPaD/FfWfZjNi
8epZP/jVHW0WToTze4Wyjchd3CnmtWp6sL/oI/KDGO9u9xtH4VKDmkksMWcH8H5f
UhjxzEsGr1Xs1Vs7PX8oh9uLzIHkg9HYocdfvqa1DPB8FWr1lWTOFK9PBFgxsAia
sKuPjweMSbwsPgPgjULrm96TUOdsX2ZyD26EXUJsF7K2s5KCogL50h1X1zHpferL
SsvVmrvuvbXEoM9dfqVhdPVtn0FUvOUIai0tO5B5DsKCWxdThe+ElyOl0CwQ4ILx
DCpohh7CNKlrwYm1UiAk+OLJI0CjidPLanToVDNpsfmhcd3CE7G3tSJF90H2uUGG
lw0jBL/htZILjgs79Ivf7qQcSCaLs76AnEgX79O0aaoG3rlAWUnI8uKhrtTNW4qe
FOfRrPJkuQVkIQTuOfB618aVD7l5uwytTqT9D4GBBE41A3/yoBBQyn0pePWbOsa/
hR7KBL1+RE6Oxzqn2zkC2vTMEJGs2ghC7a5gQxfGDxCZ4LnNKDAuwGjPiLu7vfJ4
1J8ZpC0jjX7jE5mAAKdwd/J0e8ExbG6/v5Uk6yREzMYinpyyFXXrjWJ0FhA54mfq
j9zIBcSRvoCWsdKEYxT80/XE7zO5uveeWG8vMSbFiW60sz4bfD0DEDvOmmC0xgBn
XRCJvIz14QPipPNdwuCdugV04iHqZoM8DcmPOWC0c5K7O3T8Qv8rM47DClIcIc8B
UBOfhNc6QN6Ec1BEiqWHyQVrPfxCJ62+9TdcokaJpH4m5YTuLeLRzEErS89n4Uw7
JuupafsvbezGrJDmZh6+hSfUqJpKvAUzLbLqcZUHxLuRHTR/ZnnAvjjBdODfDvj9
ARAmJaOJPlD1RqTS8uVF2IB9azzJdkDMbOAT9HtBu6LFeGsIzP3jsCGF5pLRslJq
9BRhdzVHhuF7H1mcp276N/STFtztkLsaFMuYT6ZGPK1ETDB+TZOBRUlYYUl44HBv
FEfjdsAqAcW1RQrS9JAcbs01HAvzM+jilfS0ePr7Nq/QuHXfS5Dc0PR4X1rhVr+O
s/cjS9uWM3O6YSzS/EwK+w0g4U/q53B+8/4U0F5xYv0HAfkXnMT0wH1cIJvhT117
f6ex/MP3MvK8EkbFMcWVlec9ub9laCCY+4wrY2h2UPXdSM/vCY48MTStpvJYfMs5
U3IQl+qC0DXLG4W4StEV1i01BnafkzX/GzzL6JApoF962+5SCccQtWbelCpqs2ed
o7rAc+HNUwIIF2fagee4jpsCCBSwQnHBw/TWxhgAxkdPNqV1coN892n7B6CtqGYP
8+VTfnXMnxR44n7YdcPjDvGL0BL4wYQehhU06VRjRA2T01Rq+Q5Q8RUdRTuZ5Xiw
VGy00EN6fw3rZVVexiC+dA18xJJQnMkKjpKkMI3wD4QVM8N50UnXGeQBAmL8gTwZ
0BlDseEUSE/kfiz7FnpiWWLwWgYKeopCgpbstPC5pIAKjqtkxRQNUd/iShQrUhFc
VQOAJI15udSocoCSXVHS8lDSkKSq63pudkMfwK5ocS6XwnPkItVA1utO2NbGSHSN
+LbfX3J9jcBr9PUc0DUs66lOv3lj0MtTxq6z8uwX2xttMJAlomnN5bXPpDfVPlsk
xhXuaI31CtgefRfWIBkYajGVYBkiOu9dbbwCtFTLgncA55CjkaEN0w1zK/dAKY8h
15/1i1VWPhXkrRRdbkpaBZiUafgv+1TndhD4VTcuH6929Gw1jKsoYbTpc/+ZGITT
mHXknMDFAlmatqCmUvydpD7mogTggfoMy31z9CuRqe8WN3AL3kml+2Co5er84Hp7
/Q8aQcYwcZc7B+pUPADrprcOtsZe95EMhrJV6mVYqJZkwmPBtfq+lVN0YTGLRXxs
YDb8JMfjVYG0rVJBVU4abR5u2GEYAuAHj02TwDv3DkRTmLWwZG5560qUQ3LhqtAs
Sw0kLgXSCJsY9hu247oYVLWVH9D0SMkvR7Q0VP0x3NtMBtjY46IDa4shRDcDDpR3
d6XiNhIPVi6sU7hQIdTLVYjqKavuNMSlif7H/86eiuSHCr/vyBv7U9Cp98LvVEuA
VlM1MY1xaJRfA+LEjf+ixfsZjFVolPamno91ZQ8aCFChpU0H/VTCvAmXIGxrawFj
Kga6675PFBgTFi4h3F3W56/kXjOCtaPHTOTa9Q7yQyVZ0SBw2IfU+clMZkSgmmnl
A0dJX9B1F9RWtQycDNP1aenQy992/yOGIi2cdRLpdp2FFAZ4PyC41FQ9t222UVD8
XvK6wgIQ2+WCO3ZU+W8MfGnnuYvE6sS7bPiOWZcrITUZuOi+r5nOjJpOsfRHigq0
mwC5LIIDDwle9okLm9wICxUJOebxUNfktipge1So5eQNSJzRBM0uGKZpRBJKs2eI
9X5urVFT8sMh+fC6V+NnKV6hGt+BWNnw8ukHw+XL0ZYniY251n2UFYGYygBlzW5E
LAtdT/mpJJ7pCzk+OikzAm4w0P0I5L4i2fQQCo4psbMDTaQlkV79r4BLBuejIGxE
GPTEt7/hlxxxDwG2Hq8GF0J8iBHtR3pBLrx7gGPtAbmSP/mvGOqXnXWZbtQgsIfi
GGDvqoqEe2C7LLfUjELuNCq+/slE4ruB4bJuHJEdEbP64dqTML2iW/faBm+8nrOG
nCWeljHCcv+FE1DwwRpp61ojDq6qnTvzm0nnVVaboctNi0K9P6HqJ5eEAAw92GvU
PvPlVAbQz9rk7J6GvsukXUznaScHQwuiakwagFg2Aif83TG74wW0qmfJN690L7DN
JtRGTmHD5hPB6096q9b4S/S3ibHrNk5GN/5OQdvz9SqrVhOGcdiNqp+tKInmBsAx
j1dl67JI4Yh5/DBrxbjOrgVwrgvv/MVTX5QG6j5ihFcr9HmnCZjDEVPyvCH4DFAv
cY6jhjNdNhy5Wc3Rjz1LAWPclPUQmP6tpn8/arjt7w/menrVzZNIdmA2wzngNtRw
Df/43XexO4AB8aQKE7v0ehlW4IUG3OyP4VuSezI6MKjdq02IrFHhuJWUdhaIu+ww
HceOsDOJynKyuKOuyfmQfO7GPUB9tDTqTREqCma/H3AJYY1SVJEvCzkWiNVMYpCE
rNa0DojVHenFeShI+YIFZYPpRiqzA+eHiN+c+dGYvoUq6cPQphfuwPWXd9R+Yknj
KDLsUr2v95IGu85SlgbfoN+aYiRn/sFCmRmssOcV9OqVbo0FZ/X+mNKrQJZNB9uR
E5Ey7OCqT51wYzazdFqd0W5mRL1koI4RjupEMfcxnw7AboJNDLm6ek2LFwupUmVh
KHdOSDk0xAlkYsSFnnREIuadFG0L4JDzLFhJQM9K3a6Lm0GzPvxvbn5wm/2BpNZE
xoCiXaGle8mQ10ZT3nqr3FfUNDdwaXpRJuyIBwzSVJirXlL7nJrtfF7UxyplQgYe
BreQnjmFBFnnBAKIJ2KuT9UmlqRlM1EhEfTuR6qmESo1SDBsLN+IdmZ4r2TLq2lI
CUU/0w81wq6FssOvQbpicfiU/JPnOnicppR0itBbwP1P6nlIxO1QcR4tI+rgMoGa
DLYaMTmUsYUCOCcL4LHqv/DFYZsuXm6UvEqvk8XVbkkrKJYBl+OG+kJM/ArAdMtU
TXoELVH4H+ZsEjQLO3ttQfKxGd/v2RgwEXzJnO8xBnI2R79c5HyhQ6VYZr2GLMNU
aVijarHMWE5vRtiPgIOhV0Jhk2KjsDY8hVgicOZzvIH5a9A24/6mcjRoPNZ4QdQj
xQWjsFy3KUXcKvv71UqYreTPpWUcKlf+sKnZWl5oioBf9q3Hh+wYzhBUb5qRIKjO
R6MDQQSK22w8e+GMdiD90HrZWaAHAf7Qii2IBF7hGPKenXMBuYJplQZisYJBkwyX
UJZyBHsl2D80FRfDA+NMmr3sbHReVCcTPLgrfcoP2EXQQ+F2JteRvwp2KbpgPfbH
1NlAuZ/C2Voz4OTwUv5oJfwxCaTr7Ag7J36MWLxDiVLa15QlWLB+YSXpZPsgcdCr
ci8d1KU4LN7KvuSGlUTytqKgmErirkTtmlqJeVpJ9Scr9gPXWvo6XjtBTeZxMrt3
K/2o9peD3DmXhRmro6PDd/xq+TgZlsSKr4PiMCWCNpQp3GkAhJ9q8jhjQUA9Ha/s
JjsLhcQVwkZZDN46N+kVbBAcPZN8XxPK57U9jwBzEC52u23zkcCfSonznp/stHaG
5xLK/D26adsxik468/hylMUYcrkkoCP+b7q3KL5Yzy767yZnWTnxekP0V24Ydgm7
Ikc9h9x4HHaZGJV5WOAvm5CRjunVN52PmYf0Iv/2WA8TLj1Edy5JxQlIPOvtZh+6
BmVlyu3N1Qwu/vzV1GfQf8QrwJJwn/6zxzgkId1AJoCE7ddq9DaBE4+qsn49oYp9
jPoUJcuMtym6S6Bh2iS8F8OvFWdGOjI7HFFMUpYTTcAURqeEco2irhhf4y1fKnj4
vfFwOpTAr+QO/ommbQv0c2k7RW+GQyzhDbXzvledN1BfVKZMOJJzJdYVVVzSrFzG
uD98WU6noAJedPUhnhGey1nusr/8zGC3pTAcxFjSYfRZWuTn4vao6UHEDzP3K4li
MVRxsVm8wQcH8//XKo3OqrJs+LHAN68JPqLIL0sKTMQcbDT1f922OKZqeogJ/ML7
i/OKhnklWPh7lN3Jl/U0Y0K6QNy9xlMbDIyC0bQA6mXY1+9x/AjOjQMcPg6HCEfl
57qyOp93nDPOOn9Xq6Y1meCWRRIOEgUKMMP54CRj6czVzDDEzl89BAC1Ny4J3HFg
saft2HceDbaPyJSzJ6b07cvKFzB9NSr4em+8XKfwrFpoSjA7IEANhHnpYfxs4Vhs
Ec7sqoowGQTEXob38qDJZRhuAjnEYAFlptSy2oHMenrrncuZQXHWBwVw5VTHaWeO
XntpIQEbxVyTxpEYld4vJsrkQ7xeF8ma0CeCVC8GHzrDT2xqg3lSwSiWoj3XdAzd
1X4l2hDTYT4iLqaRnuHyfMIOG4JNUreAOEFR0jAnsGpBcFxu3oWbPpJ0I3KH95dr
rBlL7NVnj44hIZxS4Dog43KV93eBlcikEF91S82aRh2NFHalEKxdbZk2p8khrKy9
RuT60H8hCrhvsFImpHYUL5IuCM/1qxUZ6Zk+c4Fj+nZdwaIVmEJemEkwH9+qiTqa
FyHduU60G9z76T63eKO49/MYzUzOXxu89xQgIhDsDcpK3Dn/A2T8H65Hrp1ADuKd
qkG4JHrRpzEvfJygpRpB43fIPzyg9VusFvdq2q+jvrMuyBTB6siQGO7LVfyW9URF
E48pKnV/jrb2M0IBMpwC/o3gsGjf2fLcpv4MxNh9Y9VJ4w04VyeSIQzOf6auVcMw
cadQDR8IAw9ExQFEyDu7VdwMv7T9pAAD1Y88X1c52ngZlJJe6B6QDUlH2pS6YwAP
JBQRj/Nqr6YojXCp563q7sjc5I2Qp5OSdhtomAAe2LnIi/YHK23I4Gloky8TaA2J
uL7V+8WO1L9TmsovC6qsq7RiReIhn3GzYgDrAtvI7eySmbthIathhjJS2JpXKR3+
Odr50RWy4rxl0+p0p0R1MO2zMJMr6P90Fvlt7KBhOD3QGV88ELxGrRKNMt0jnu4I
M3bVSdM7MzMRm/Y2hdb9kd4Dsx1d0uMlIMefyAZq1TSBRRKaNvw8AT18uEFna6e/
PinvqgVeRs7frhBQ/cUcPaf6XA0g4hooCYWzCvRnDNnsF1t9Ldd9m3dbqG4I1F7R
cqWBuDBrzn0nqW9frF6T4I4mqC+oKKpavcEyyQ69QUujLIFvVViWmRSkFRRs/ll+
XEy8OJEqfunw8UXEh1kC/KqoMAfEP0oFGrMFslbTOtDBwAjCMDcbXj9EmAWtUq1j
p8LDzPa/BiHg7S1L6malFTiVPzOvRjWtGLSIhhfP6kzqYMdNtsu/LKyEwt1SxVlQ
QkXJTEQ6wJEGKr8NfpCxbyie1BAwXWxAldEL+qh5MEEKBVPJYZRzxEN1Crk5IB/P
37K/s3Y1z0tC33mbxU2wLlr5x3/ZB4KLpluxtm+JgfBlNhSSb1490XlOxB7oCTf5
issH55lyqyXn8Zf6qtLyQueiwtbxJ19fV0/jGG0geb0y/VAUlzLzL54EJEHKaeCf
SehacOBqH774fc5GHWQVN3DdrsVkJuqL4suCc93Ws3rQH/65t16DND3gznFn/TSD
mhd3WiGhWpSWsKoinLiKJScnNxGvNDZc40Gfqmp1VZwQsxpw2jRYRE+sZrApqqrY
Ei2yVjR+IAoGzjCpvR7v9MPbQGUTuJyrcObMrvn2hHMAazwm8w6D6TiqkgiemM8g
brPvfqwO1PUyZKxH9E7yyn5vfQFhYCk/xTaPo3yz0YKYbtLSKSWyDEBB29+ssvCP
hyhhLARoW4XV5OHKT04YtMamPq9EoxpFFSKIaJzDsp2CtjMXITjRyJdiSIoxA7FN
kmLKV58dK/wUJgN4+ARTrTNrXr+MNHWq1cBWmpbQRALkO/h/Yb52qjySGGEEQDum
AUag4mDpsvxquGvTYfLwV9S5PAaY1w/SRh78vmOeBd+/CO5Kpx+ARiWHOKmQUShS
sLILsfp0Lygl1Zg5yUdulk1jZQwTRbla6c7EaWPsM7dVe4ycR1+539+C5QEdEUB9
/FKeTuj/JVYB+0jjntgpWpQxLPIkQ/ECRKGXf8C3NCg75mchyKnzCeuJ/ufG02w0
wzXTQXRkRAWihrBP4bfb+D4QCPvGWlYEfoPKeSfjeZKKLz8VqCDCRSWpghWmB+ID
2c8UGmnBUIpgQwWxWZnURqUMeVsprd7Vo0hlax4HxZrEN5pMunR5+0Gso040aFVU
apalXM0Mv5+gwrwwRX489miEHI6Nec7HsrZ3O+z1L97UI51gKyaleAWWk7llqiWp
drqjoFH7Fvnts7VGe86biPv8wONkKkL1fY1Tw3ngCnK3RYxuqOtqhSpQEUdgHj60
jB19zqAkXs6OpcO1Pd8ncM4wg/kpXYUHgSgRPr6rhUm0EH5fPPO+fHi0INGZh8BD
52gGouXSUIuwcYtN40vrPrpHSiBgn4oEsiJ5kTJ2aGwLJ9XoJoH1ByMIcPqxiic5
pqIQ4A6OmQcv/VVet0waO//hE5le4aJOXRBmVn++1fTy4YjjbGSiYeUjoXo2Wg1y
TOFotCql64RS8r99OOCEr9ysu+OaLnFhsyZe0BUMIKCWIvyc0n0Qn3bqbzJuYwdh
lqNPMqbNQpQ6mzrKvyP9mzWFEu8TTKaSHqbfK9roN5QIiY7cAD07z+13diFSCgm5
wnblmwCKAL2mIaoS1p1dQxoimY8VPV65U3nSSId+B/xz6VxRkvtArR8l3sweHIp7
KGnp8Ze9pWJROaSTcLVTPI7gUssXcsm1CbHtHAUPj59L9j9ZjhEiiD64ApGWqCq2
GM///BnUueinRqQXru8+rcO0VmDoStlfYwBmbvC6q5WJDtDu5Aub2fQDR1kiUhTY
BmlNvJvamzhhECJV3CbugpdEQE0+fDPFAxMxK96mV5G3Qr6a1zKNprcuTc7d6eKx
V4Kek28pzTOHw37qgyV95KR6YCE/3P4kscly6YNaROdbtovG7QhBkCqWhcwMLOUJ
K/b17wdJcJ8tqKswxmHC35mCKMJr4GF2F9E2OtPWwqci7eedo6cRCoCcHGb5FVOy
1QnpK+Ypc55bAamdI+I/WML0ebWU+wquFK1EpzZOaC3Fz9J/wsCRCMRcJVf8BpNO
chI7IA7HcQmTKjz0h2qv4KgZ/SZGL/uIaoZJ5Q56a+Yj5slDfqvlyPZSLTmczBEB
EQ6kekV0q2LSJ4rWEtqrpGRw0GfAmhrBUlAJMphUASvlCz7OMysFM3L/gMl4CaHC
8wWGXAs/IBv/Pxj1FyBoqJmTxxI7MTT2FZQ0BolQrmukcTWC/JVv72PQY7f00Hpx
uc3uug1FYcj+QpyhvbpUxqQB5EvSAr2CdhWNxES5sTdkhxDlNZd9a0geZpk4G2gi
khFhqLq7AVE0yzczK85HA0gV9Y0TkG8zWb4a0LCPpG1mvfGAQTyKmm4Ud+5yckAi
m1nt2kK7emkz71MsfnXFk0DqFBRj2dg/0PRG7J+Jm9howsHtxDvdB48l+LEyD7lt
mKrdwbHHBVsjLodiqgg0kfOV3Co+6Tmu4Sjq4MMO4WZAGWwQBsoba7wajX+F1Ws8
ga8vsRy9NGP/RnNjytiHio3Kjs5NjwId9wbSNYsn8hqakWJYx0VxAi5+lb5ic3vm
EteFIzZgfa/pC6BWtuTivruUs+AU5pgHL3LIw3WK5e6I867uePvdsCZKf50egnDt
PJGnFCtFvM4cdKvdnwtR3bSZcIPmgJGfU5xahUEbm4HRCmUi5VmVBrbIZRMsWmSf
BE8l/wwJ+MjMpiheownEnTyWc/xsbaZ7caYXQSgogPWoKHjkATdBP2kx+H7Eqwci
7sRFstBt7x84XPmXIvjWw3J08aHvE7qvO8FX3rSPpieW4UDLEmIewQP8Qrs5/+mU
cMczRVBL/ejBwdhoibmDpRQmJOlZOwSZ3/S9wuYURzvYxUjxToLjaBWJmbSU3wUo
/Fo+LH70l1lahoXrgd0yZiHeL5Kh2znzun2EvlyJkipfOkz8wcEXg76KAdEey8mq
tBn5gB8ZvV3FS1NikW0WnzLL89zOJAH+lAB/6HYvVnz51RAqfFi06+GqZ2cDxG/l
oN+XeQLSb1ID/Hg3l8unB2gedh6QBIcb/XihqasO5SU3IptRZjMDhsIv5BmJTK4D
unFQmHMM6uQ9UA6uWRLXVnVArlV3b0WLDflmU0jJWy4TajYt3WPjeBr2EuQVJEY5
IOzRUsIolIX7OtxlBLyUIgic6ACZj0j/JfZwhNFDVZdKgjJSWA9XtbKADGtFckSZ
fsN2S43SumYUjtG5p0LVW/alN7jdUujcTdI168v4bq5yu5+3sdjcoyeb2fkIstCA
suxhPVfFgTfQ17prgas+CK3YhczujEJ4hpFEtdns9zuBvErhIqqAKBtYU2koVstz
eJepr5LszejlpqBknbvuxTurkm/FDbGDkeN/elknRLz9EnNEObYZba8Eycp66jbG
vXtwBjeobyOFBUqnOmRgu3UmvK2bvsVRfugcKJi29VvP9QEiK1rP3nBqPfOTjWSE
KK1BvTM4UZARa40kRrgxczT2UPjSHHmCUguVFqrO5SXhFIZT1+4dEQqtdfakpqwh
huRZ+XmEi5TM9AsKaI5P6lqa1+OqVRxifscGZU5722cyhWY0JHGr/e6aK8NGh5q4
5JDRxoXTE5zDQajUZ/SwI9zpnbEp4RMXuNQM6Fo/8LVwK0mQBaPTv/zsZ9jXR98p
H93sSkMzp/sH7ItDrFdHyYzZOEzYydYjwIj+EDrMBybHWIgHObZ7r2CZpFHGjvJE
bPHVckd/Lq0aaZi9Apvr7nWBi7am2zqL8BD2L9/xbnA2/6tNapaOmxjY50WnGOpd
hu8TiCpVm5gqpP7jrnwe/SkVcrSYUj6mRS7JVUace76oVLbGG7iC9BednwPIR15D
309DFyfMjvobgRL4sKRhKbM50rT4VYz3mJtTKlMU6L/WGzyrK0vAkAIbU1jfzN46
pynZhX3VkNpqrQWSzT3Bfk8ljqxLg4h8NZuGE/2EQshj3sUAwn4jOYiE1INNhk2x
QbryqU2lDJPPVqGpDtxYgZVGog+1LljeOcVR2E35MZ1eb5Ivms0Am1lbYZLOSzni
4KkGl89U1EFWxHA6VMryEjfaVC0uGP3LzyJNFQsqPExrPC8idXJeQv7rMxlbDobo
UOKqZH7D5CkY1lDTUDI/Oku7313KiOHys02Ha4df6wPDW7klG2RV74Iumh4cp1mx
gQsG4gxYOedC8UPmGvNHIanjol8UV2w5ZtCzCiIVt3rlEY+QA90l2/f62id2zLzF
0gpC/nueknM61HcMlNr9SMaKEaDv0Gr6fyRTu0cDhbIFT3Fv/ZefDekNmJMS5w51
rigtzyEeowkpWmbh3oLyKUr+f3nW+x9NUlKcFns78ypjsDMwEUo/aKfnA1dwbdZ5
gFG8pLIezPPzuPmkJ1OQSJZsQi5Wh1caY6krXlibvt2e5I24ekPhOHc94pN5XKN9
Lkozx7Rp6EdCpXBuPz1XtIjcoP337WyAINImnsJNE/fVkFBioOTSVYhkioxU44OW
0/7ZnYkfwcGjO3h76n0pFUEqUK18a1zIsg9hhZH/TnPar+9R5U+0ZvjNfqc0N7xa
Ppit6FlrNUakleCNYZ7QB2BvrxW/l6LMzIk90abA2mezIv0Sw/Hbe5PQVqlerdFb
eNAkNHVlNC8RlpGveU8opv/cER342eID9HX0rXQ47GuY/CvZG6vnBDZfF0rhwOIO
9bVFJXsTCET9RrzXxtCHJYFMjhcCj/GGumejULYbGnj/UZ7Y2mSY+kfdburgtLuN
yTWcIgQ4iBeyq6OWru/sB5Q5Rqw5wNYTbRl9IWKYW/1sijRJ1tA4n0pJxJIEITNb
5q6fA/U+7sG8iJ1lilnSJUpkg0aU6RC5UZAe0Svk2WzWTPq0QWFe7iYBZHSQ/8Wb
t6lQLicG4NJlWQWIyxgqHtvhuUvByYMq4ZhuyrXYPZe5nUfo1ZuTG/uP3HBlUFKI
2ALQJuMomxDUuSN891Rvb6KcZUYE6zfyt/jUV/qzxLTTDt6QTjnu2YKNdvIe4S5N
m4eaHYPATAc5h/gyGqidqOt0xPD9t9kabtov8+HWPavpbjzWyZAMPh9LfAQfh0YB
qQGTx6muZWaD8TKpsF2sbcApRlXLxVOGg86bX/wmyxJOM6KhhrMthFdpVTo8q/Rv
rWfHe4kEWeHl+rWqVINNuvrgMTpry9TU6Mju0+LaNqHKQ7gilzsI61eIPTWvHctq
/oPDuaQtsD+LlaJmL6gioFC+9CvrNXUkpyOAODOk5PWnrvG4Oi+ojqwZCfpKKpVa
BBJYZZTrdVYWF0+xI9EpyBnog+9oE0Sj5PRCSvi+3FgooyTqXlLNM3p8hZjyScbU
sh5XeX8RxV5L+UOzn/cjjDZJuK1Fcqj1NUqF5q+qjwnTLAwbCTm6LJjYOaqynC5w
yklPBD3SvLM0fUL9kZbf+077Ni77Tt88ugH/XETMA4ygsuiod9+IlhWC0jgg1UDX
bJtbT6eCuBIs7/GmSiU3+3SpTT9fl1rA1J/K4q1HJCl5JPH6iEs6tmL7X9oT9Ks2
v8v00t6+z/5ZLtHrcH3KcYhh/XU1K6n8aPQXWJymKt35wGMiwcLQJiT/dofCF6b1
QVTCPz3s3aiyr9PJb6YfccOhwB8FVvJDgU+TriCdniW/FyjT3wv8+96bmX7Cz620
+dacTZaDopYSfY0aDh3OW9G+LKgLUjT1cbmYMAJQq3G7wSszBKxWlA3/E5LAGEaS
f2IhjDunoJTkO5YOYudmj85ZaNJRK2NIQMlCHQpCcG0S/LbCDBfwAvJ9S0fCZ4Sf
YGfb5nJmr/Rg+EgcwfIXQQglr2aL9UMw+rXkEdQsGTAI5bp5hwIsNRoWJ94YKSg7
67Hc6Ugq+bKXlkuOm0y7FuibtZ1UsbtYeTL6BFdI8sLB26G0NqGw/qqZO2hoFp8H
5TgeGdcLcdySA+Sh7XZFIV22iZcnQ7m8tedt9L2DPyT0Id0kH+BNU/8HV1BKDXLJ
LIJU6Hv9/Mis/UwkDYx8ER5/QsdKL8Pbfnf7nupkai30cxHXjUDj1xoHVz4n86Og
/LyxWNkXmyJsVrrWo+fwMMxqAs+VMF41vZoNkm2SRVGxBjCi1tYgpU6p4gEprPU2
TZwAPwl6gN+/Cx+gJ1wBHHukXlZ8g1kecl17Zo/x8KJ1ZrZeWPnctJAbNKEKGi1N
6xpQIUu9CAEgsFn4SW7hsPI3ezQmnX1JAAF1y0CJYLJ2Jtlv3tYuYaXW/toKNWWb
e47QvN/vMRvy30N6EBmrT0HTaWv6lxoa4pJozTvGF/KowNj01WGD0k9SXgUqayoK
hi4gx4BMyVxkrgXYVP9iBVt4xppPCVr6yn+hLj/PXq9bzvOz2TU6FBiIPwzsFaMN
68aBfzlAMTXbMUjqmyWhtOL0KQQZB+MV6HS2GhDyh8kl6aEjQaDHZx2o3FZ53LuL
OTKpXMMwLURTQweU1loIe0z6SnUiRfux5HajwqqWlg8K78T2oMnZVV4nB8ZU6t9y
D9zVyVxhnRoMTRG6Z7WHZ6CpcmjRfonjuyArh8Q9EiyWfCAag1m4a9WQRxI42gGP
CrnUMtz78/yqx2vxw/3s/xTnqvUGGlgJ6yyUuM5nwKfs09hRaM0rD1qtxYaeGJ8M
lQKVvw34HdIGEPzifF7wFYuPeflBBeTftZLljrraIbxva/AQY849smoaEw3JgGXn
uPQsAbOtmrymh5Iko8XiThD3SgAz1U9M0RNbAcZjNN2SavSIltAS27zzfWSKiuk9
rVfQ862HFMnWzflAseOZFEjs87RChVqhuLnJUasqQkXW/VOPJHbHRrPwxsx3WNta
rJQH5g3vir7tSaB1nU7rttXGBHIW8yeFg3o4NVR8rIEWVFOSkBORIrfzIrICmp94
wPKAY8LFCXofVVaOiGtpJ54hgJzabI0vQXWA6TWbpm9fAYxZoy9gpv9xQb6tQ9F2
koO0NaAIJNAv2xQKcoZCnd15Ds7/y4XMlEqVk6+O39gKJDRD8wicpzW+1NDPtFBy
TyxWIdkMgJVOT4O3WVF5CkdtcYPcLFisE7Dk3/+YHasr0RCajO+V4pqueistZx0E
yystYchCDmjhfLvpB2xVRv3Zc8ykjsbvko3S/q8wJeYwiMIiZi80PqONISJySwAr
q59YqJil9uYGiFs2temAkj12V0XSH6ZKkYVP88dHtCkWGQOvGesNwXAj9qTwilCn
zHA09nlBee9bUH6zU1ePbYCmbYEDv66FdFHmx5JPHJwDXI9eTdreUDb+v2AjimXU
5u0njPf+1XSROZsvaN6nUbxfHfhSWlGrd4zFVdPvLfjOYuycSqoob4fcwFgWaUfA
p+67syH55Li4TNhxWQvRlfT6T/pGYTV3WnQeL+jr8H6ldAnYhWxVNImBEVKaVa5d
9MCgFS+a57ZxMkXIBVnesxfEG5FTWrccTqMZPqmvdbzdtKbsWUl4Ure8nbWWUWFD
pOX8ucfQYxX+ebPWF89vHU43P2eOFtz+TcAT6S98YGbOEjujvKwZPhlYrmvI5FJ2
QcGsQVhE2Xj6CxqzLK+jWwy+sbF/eTmfvnAYwILpiZ9stHlshir4lEw5+kHkHDsK
I/JnXjeWk9FDX+jmqBHFt50Rj8jD3A4SCm4Snlt1YW4JPKp/F1KiWwiIjlmh+CxY
QZqxz7e8uORZIWMCtB5egOKGzqjZA795HvloDL2AijCLSAGXwPL+c6lcmo503SwB
AyWnzdoJsi8nuJVDFDVjj2NuIwZELJGoEJ6vu2JyTpU7t4B6RGyyl1rVDZ9CV6wn
g94NyNszaNQN61NCDEEZRRgT5arsQRVNnT7RPCn+iCWMdGAVE99w6IkZgApIY4DH
Kvh+xwTMCpcnFTSjQOgOgHSjPtEr+zPV7P5KnBKSsTtMOXqlyeNmT2ykIuVO1jph
LFGiuclBWttcOMPxeeCyDSqV9B3RydimMBMkGLfGYWBHI3Vztk++tTjfn1rYPFHq
fz5qVAqdjQL1SiNDW+xftdnrC2BbWzJEMnRbr4+DbAPYrz2IaFbc7L1hAPUpj6dA
WkncaPVNmXUp610zQ19QPjuVOToecp+UxJyPB6+lMhCof0yId85kHLjT1FZqE7wK
XnB6L1w0SWiGLzKBeqBTVFf4y//SdVf/nFOiyBZ08hm2bjhQWmD4VmXhvst0X+vl
J+6kMmGpc/hKA91Tv7C7fdBz0eR4ewD/S9CNonAH9jHdSdxNYTHxRnWJmAvVfhmV
K8XLT6LiSqeEre7NMpe3mEhZlv0+i6ZGO8nQbwmm7qheaJx4W7dn75owd/DoRK61
J8Nu59LiU8X91nEBaipz/laKXmH7RMdIoffV1ZATZ8JGIGCAZABzhxaefqeuX9Aq
niGC6rjun2dGguuRtVbiLNLUVU1veOLk9GBW/L4rS7QzT5BIlzBVXCkwTzW8tTsS
XToR2gTxME0Y7ZOYKPd59KNJuNCNuL1SZx5GrCgQLXF5MxOZ7u9GkpsLYYTOOjDv
vMQx+aGBA0tyqcPE+p1tawBw87MdCN9mVbmGXAg0pByirgNsrJ1vELe5PJenu2/c
nBF2w5y6CwPsaKEDJsk2o4JWx5LLigel3HAe/ljXZWOCODiJECxcf6Zmncyq4DVL
sttS1YPOO0+ctG9mx/AZes01MFKDsh6bOuJ5Iv/TvF9n6f3LMq1/3b+dZCLdYa8m
8VdVriAamiSUYElhQZ2JDzqoqBmfc42Ko0OL16bZUk64YEl7AbhgHwteu8ol60RN
VbfmQ+yEaX2+0ahbwbujmYH09847AGlucPohbEir7cimfVuuEVdYPNMpJXAZF9oc
cEt5MmrULpdRYYBZWfYrk1GAb9wK+4wu29uEw8+4CgVEA3DuPlUkP175Uh5FXRUO
o8vzAJhyjTMuvokvOYogWNhcm71Fi2ddzMu7YnZQySAVCrPW4xpNkwrPjfwtABMy
GU1xLI9LX3io5ur5NvW7KJMbFinCMl/LrFTIvmpI/SFgion+xBPVAhS/vUd81Bua
BtHp69O2f/ew2kMycBHRr0WzQcaTKjsoXVHboIo263bG367NgpN9x68b5XtYsjwQ
7ycj9EO4VJhMZO1AJf/UZgDmKgk8eONOgJ6hek+JV9v+L2uvc2c46YbFQxa/OiQ2
fYaaES4NggBGoX6ORbRoXe5FFgm+49z2/VW7shRrxLUqZKrTjNfI8Xfzn3r23Xxj
swDo6yLpnNnbDj1EGXuhMYOWzrwDsYOnZuKAHcQuHvEtg7ULA9+3Cw5KyuAOdt4w
qjG3CzVI0MuY/xqqaHL+MKQLvYWz0e2yS0LpYNKVqhNiraUOMK59Nt/Xhwl63W8S
dS15CqMpmgd0c31LJ/KToCFMdGuSyG5I42Rl4ppDfM/Ca7DxYS6otffyagXjVXuE
25RL6whXl3F+1DUxJVVeDZ/l6lmpTv4/Iytpc9t8BItMnJ0htaHM7LZZAQk6o34Q
BuvkZgJ+HMlwRZN7MoMwrqgQ6XqbIQ5HbhSv0vNY2sFmfkbAYahaKB+/I9RucIAp
hgFYs2cVlmvWo6Bf0f5oEg8tMLq/UVTu9imEA+l8cmbDXRGpKxsICrj9qMuuRFgs
m5B43eXN7L0wH+8kbVlUDPrC5vzx6AaaZ2FpKScrgkF//HHDZdCvBeipQd22WuAT
aR1xGU0vujGPCuu3GJ0qrT5tnZQnSO9GxeH2sbi9Ju61Rc7lCpKFEWRoLrL5ijF4
u9oT4p5ep7kuyPhHXSp2VbdgLutqhzmFF32U8AJyGkzCGi6fq9uL5UzjxpC9VvcL
9BC3Ir80Az5p4xgXngopuSVFeiA+a0+rlXzlTXQk3r1HmLoefR35IR8fTO1NC1RY
2vZX45ZlX/5bNrPMM7ZE2m+p911vGFnMdr5VCXm1z1tJLHdmQxPSrU7PMoug/9Eh
/vJHgTR5fV9fUyeiulWOSZ6LUxYcaxJYqBgNgYfMfiLnXXcEtwFMxGc5ZVx/nZJZ
/iAQiSu+ZDC80MbLgZPCTmy0oVzi4oaqZNdded3sTtVG0Ne2aVxvmWJ21xm4IMW1
Q7Q7qQFQokGfcZ8Ym/oQES5ASB4F/YkhExCq/cKyYTQ/QPK2IYi00/+LTm8ozUiM
2u1ZcB7El07B4P2FfcFg5fY7XahljIL8RkoCmR458bqxarO0S0tPwHqvBQtehizp
7096VnLc3pv1y+4O7a/R8mo2q2pHve1wT4yiDma1xsdcMJ/nRGU7QbfyI48449dw
T/8gh/E94cJJAa1vmMTpMXbTfssddHBLMA7yi81dfmko15Gu19fG0ioQ8AXPtoN7
3z5L6fcwEYKrRX7x+xi/LESxV1aK3Aii1p4o9q2/92kIyPCRjmr4ZWHAicGeKxOE
Ee3+9IfI7PpaUEpbmANkkY4Z/5AS1zkqDVzUSrPJp7JgBaDz5KHep4aonkohje0N
Yfu3AYH+fjlW6Y9eXKeCdhcnkoaD6+Z04X/6uMBdMrHYL3MUvodFert+GIaJGB9z
XYDPOb66b2qcJeQOSHhkKyGVQ5jyZbnRtRHvK1FUpTsXEMjcgkFOYOw7zre44saF
APSKfr8AvoK6YnGyIGmgn4El0+43ktV93DMTLxTNctfO1ZNwNwWxRWicogXbuhke
lKEsOqgNJJTnaqp2dFcetaiEF7StygToCGcYyt5s5oYRA4WT5YhmqryuypJ2P9no
+GzI3f3U8dIQmAJo+fc/lItpIyxfE7ZS6uMpN2p+s7jvcIH7+e8ZaQPYNFXFPBXY
4hdbOXVy2Cu7YiRsOQKAsc73GThP2f4ISjhnBfrO39iSvIaRKhlYB4uCiANoL0Kk
JJHxtmfFMKGjKkRiTFSPcGrBCOlZISFySdNexDGYRLQo3eqDn+BGzfwFImMEqVva
TLmzGDOv9NPTeM7trYc1ub5KKgFXIDMo3LYmWuKmF+Fypd3guo9nbz7vyXH4ksmw
UUqPM9Ba+966zuf/IHTL3cZNzTZagJPvXMdMK80q+B09YaY6ncE0ViTqMggg6yqL
nOku9cmSOXjUJUmlkO8dNz3koZF7zcuVr/6Ir4qugIWJILrbm+i/xrLnK3YxlRGc
KMNTQqi/EW2oXcdZMbB8wk1u8DrWPzN9Wxx5T9ttf2KMsiLmxBYsXjAEkfrBeQkk
Ia03XELnuc8eRiINs11JgMHNhePGULWQv8eS3CyjzNa2cvycbmHknYemN4RZY668
YT8IG/g8Mpn8PR8rpNtLqVF2ANtOcJw8dCANYa6Cr+idV+yqZFYtQ2j6td7gJrPc
Duyqex6/VshARM/B7m/+1ZhX8KonCC095krSpFadUEjPFqCie2DgvBdclP9zP65t
ZEg8vayjebbNYpT4toYf5e817sC2tEhSJAET/5jxOioJGO2WfA2aufPG7I/FQMF9
C/Mjzgf6Vp/3VXOPn+uG5L/1GU1QVDUSFGn7GGgsj3YFTF7aFtNkbZJn7hwuJK1i
Zz6Xrgtr2JTI6jJ4fFGpijgsa4Ng7n2UWAVZJXE3i2kh1we8DrvqNNhEWcYByTLu
pHm/4p+Qnb0cy5X2FObT7IkgdDF7zvhTUjxcY5NHsCdV0v/wEMbMEXKoUHdzZdpr
5pGrAnVCbaLl832D6qYoCBLOCFvvZ7qmHECne1KaYW3ih0iCWy6JgvfxRTVxDDvu
+E8pes3vWkAPXWhbDBO+vnaYAYmKQSkH245XScuIaZ+JMH+SuwtNqh7xS+IKBLA1
DYCSOSxUANy0vuViYHZsdHwKhJaak7CccGAXCCcngwobzTF7sxd9SZmH3I+5VZqT
SOIFVJgGrR8W5mLr3wIludAKwyM56bqSmk/0nMhiOEJupaAEIdvVef9henti2/9K
IaJ9g7YD/K9KuZVS3R04++F+vhg/kP94uV07jaOzLkD9NUv7w0MziuEwzLarEpd+
lkBnBNNPpBIw5WvtDwxnzAuHMimZm9tAssRzZTRWfj5Qqd5Ont8vcW7GuFul+HEY
+dXWuGCKGS1zWeNpOsHe6sJJdroqaFC4JbyrRYZTy36mS+Pj0Xs2FVX+mjK5Xv01
BvD2WMh3bvNo/HIKj57eJAgRVk/Jj0dQo04z2c44LXDKIlGs/g5UnYN8iKKDWlDn
Zi6XvlMrKf1niCFWh3Tc1Dkgg7vd202bkWqdus5z1wwIzjoVtLZTPK2G8dM3RyJf
KdwBtWMOikxMWZsST0OIeRn3D5aSZcu++IWoPYWMZO5MdKU8xJGUSv8CbHmdpQOT
oBtSWppWya9e2P9OsD54Kn5RI0s4OTGyIJeSKgg4wKwZn+0ycNs9YtE+8oMjS6IK
e7aUsE8AFKBlGXp+4JoEtaa5KcqHQ2zRBiaihPgzqRadgCaQVpapMRBKI1S1eN7F
Wm+kVVlgwxgVTQy67sjRZiqZHqIQLlOgOs9ppq6FLsTeLyBRtXWfbi1BtY+AnbyG
DE6NxDY/APYblA5c4oxq4592SR95nXkRS7Ct3hbPZjZn563vgNtnv1KEQDZMK5QX
sSoNBrawVYDBRcezyXUAAIpD/gAek5WAO288dElMutZqQlUsY/eJDZplmhKU9Ibt
GHx4neR1CzAU2rxvuJGQFQFuNyZPVlkk4tmq4oMP2Pbxu4vYyqFEPJyVfSmsRxsb
rE52pQMLaEZkMx5Of+c2kjhPj5Lb93PNijatMyk7nGyrg2Zyi7bzhR4t53/5b6V4
xBz5gDpkh8sXqeZZ1/f0VMngje9NBpmLPdhFVN503tSnyh5MnlsIeUfip9K02q1j
EzssqqcGE+wvpGPw55+1+fXJ3LryAbRpqCSOS75E0ok5pFBr8ajW1iXrVqpfAWLN
NHNiFBlZEXCH7XffEF/qbi2hiHJvzUUEYk1gma52R8DO9OyjKkelBHuVa/5dGiBF
deqav8hXPrJqTt01BPdLPunvu3NEa0FoPZKWqDaytROS20KhrcLfmixw+JOcsIRF
qfFfPayHb1ZtbZMnkYa3lvdDPBJkemqZmVazdNzwxlCpXH3ig2fbL9B7mLu14hn8
drTAtz2OGsz9MXMC3LDEQcwC6XmM8zGDvArRdEFYKVYtkoKz4ZVkRr+vzLlKklx0
4MADfIcMlczItn+RxkiUDDFUCZ8Q5S735vNHZAGDhRe8BIGHXVahqqdzExMIFU0W
03vOlNUdMnpwrXTFsij8EMsYqnbpB9Q25+fhWECNXhLfHcEKNuKbDKtJ8KiVKOqs
srmr09ABpDeW/YVsVnPGeaY/NH9XtVCQrGPTszsHl7Bf+YRMSW+XScZn75VxdINc
R1hB6rnzswYtbSK0NkRYIa37tzJK8+4/ZKDnFmHUYAC01uvcwXvvWNGqOfQ0b/By
+TDbQxncSbmD3OB9Nzi8uFNZIQwJnv9aOcP/MJdB1EVBzectaqGNmRbsgONXldFd
4S/k6UCGw5GZ9EoTsXnY0jVcjzs4lzTKNJHmSL21vgp5y1LydwXVeYzc0IDcOVxU
2NePRmODga0qF0HmSHtJssQk+77BCBOTfvNVdsw0xMa65MxINEfDB4B14cCmAh9v
RtbLk5aDybEvHBBQJXcZ/11Q1k8LLcyDoOlBMGi/Td8piGSoo6KxwFmxWHAYccGj
r6UDYnr9jTx1U7ESPVnGDB3UhcDCCuJWts7P/oZSdKx4wkWerFRG06glXfNu2zVm
pquRJQn9rHT4MgvQOLQKlLL7z5k06Zf6FNymWsND8VmbH11PMvdicvskSZP/OwiD
sizWgYC79zM3aX8tiFU47/kRKFsUOFz6/2PHOLgS7K4p5ETfS4hnryTVFqXulfdS
PQ5N1TfttIZfKp9lm6YnylXz265d4c7J54c0c/eyFx0kKU+dB04/xffICI1zpRaM
LIItw6bbkHkXRHJYtD/ID09Vmq6fnS15K6MgGAnIi1sAl9JinHHU+R26ceFN+R8L
J+px/+LcPWH7qP4TEMFX93at2kQo70ds/Lo74PaIboJkQ7cbvIRLNy8zWbnK6/sX
egMA+h+drMoBL7+2f7xUfitOvGJsFW2ZxAzvWS4qDjp1OJg7VwKxhOXYUQ6RuzWL
wREbWmfMtMq+O35hfosmYqebwVTK5aud0tUg7hjLU5JV5FMrsyORqdz3+k+y3Iwj
yS7HB68VdPmyo/Gm0/77trSy8TNQE05QIJYnuI49fcyixHWIC63x3jHB6S0mRUer
OidWGMXNTpL/2glSkGECWw+1jnBkOwssxezw2ujRK6uT+RqMcCV5QJ/hCN4lNR2r
eOm7gQrBAIQ7tS5RWIMumIfTM9B23xlunH+Vc7pybWEJ+Fpc30u6ykGkdYXvFL8p
HEplylCUrRwTX0606sgmx+RQQuVp/csHdBYQcM3OBZ+pXI6C67vScfNYjaNDorsB
RvAMecueEF00ra4TIoYUM2G/ffOuUoXqA1wta6QABxtHZ/jjoMZzeNNCVA2KDtl7
9UuYqyKt2EJS07sd3ig/zjBNvFFtTxb3ry1ROolE1eEcMtdxbZid/4oJOHqRFU5O
wefiM9UzGqEk5wZlisOpjozkfAeU1khwWwC3G2xh9BsFpvau4Mps7Ct4bCnnEcwJ
qiy/RdNHsJjvWNncl3WG8R2lUMXl3CCttCOKWILiAwa5zKOAzf7bZ7HilqV4bozT
jYuJxDpt4XlfA4xIab64P+mz7GlWkeXN2kGHpOF0I/3DlXixyFXRKOxdwGjN7Vhn
EHjYZ8T1XqKmBjjVUFLl8Qp6jBukzzSY2uh4zDJPyvYFU/EdmhzZDpre+Ds/ZOyP
PtIqst1ke80TColvthGx6dKOh7k2huZ8pylsVbmaCpDp5vNrJVryR31/LUcbH9q3
fPZYVj32/XmX+UQNNvCZ3E29O2SWeywk1XhCTmbRIZ/q6LB/jYVs63Ww4MxGm0tv
s8G/eEA81t6yXL05b+rReQQYqqePaSrnIsKnoLRbarHGed+S2etZPo5ruNT9Gfs3
hLudS/FCGYJyDzLf8YQq9QatcJM0SPjd5ruVJ5gPHyFXQKjkY0hSRG0sATaYyltB
VngDGi4ryVU92VKGDE7jBDyHgj1Jt+RZiE5H6GyWCPU9A8YSRdoyXsgvFIc3Qiw4
knCCXWKLnVYhv3VgEh0TIsMxjxObUpHx1vr7xhg3hZA9MHL7HDYH3ir8ZdPTNex0
QYnZ5rj1X5zi7rECkzqjOJiVZK2JyWHP+wB+cgGvgxHcMhOSXMId9K8FCBum3+2l
2JV+obbnFjy7KGA5NKegvmmOdKWuHROKFgTwWNxws1M3Oo31xjecorBJQSy1Nlb8
0z4pFfL6x/J9XZ6jdKwE5v/TWHnq2CKF9/pNzZQxzE9+LAiqUodttbBw32JMwIOv
2wwfxXwFHmtfWSUQCJ5ltgLKvizpG/8ZxLRwJVSqWoOes1K01umOsrdX6P/56J1/
XI8QgU25H0UhMO9v3AUozUSj6cAyZFzJzfYYWFtBDLwuU8NBgArHz7Qy+5t1Adun
R0UHuJoS9+PLQ9e44QkU88uJKXvkrXlRlinYEotvS1twa3X8JgZ7XkXSuFHTbwJ3
9a+Okxr7roc4jyWQdvaW1LgAkPukoGrRtqbqCWqoJ7xRQRp5IxD986GERcpCsb0e
VzqcqwjeVmWuYxtT2EkSWCwvH3QgJRu9t89BXNAdquFIxih3db5qUluArR0vm75e
2y7tTqnD8VVYzFGWjOP/Mb9EdVq5K0yc4Ju/G1NG4dNTFVjNhq9dDObaJDPSXVsu
UB1GrDaQ4J/nmlFijVoQyXGgDyiEp1/U9coFtBWoA7Te4CxqBHVns6dilZayZZ3P
dx8sXRplaPNxthw3OfM3iJ+Cp/U9xoTYGLRs+1RtRZJJn38O0GlvDmO802EezcHx
i/CaAEAwZVEj6Cfir7UXgXuj8sYxXwIoovGiCoBmJQqZB1rR3dqHldnsLXoLaJAe
5wPSN3yR4aDlMF8Ri/ZEyTaYR/4O02fFgxM5txVrqqcFDuGLybCtCh6LhQGhrQm5
/1L95Mpuk8Ql6sw8dXCBbQCbv57/bG6oPRgWyQTjqXqLZxvVe5CH2jq3QUev9sI8
Lo0EnD7F5gqrBWHyZJyrOniUds06B8rhP6dXYUTY++BDLWUDLxkgGd1UtykV25no
gZlboF1vwssf2pFYPR2ucEHILIaNWjQ75yigEsFu/QxqM0QK4xm2katQN7M3X7vI
ZP78Kf84tmM4IkhhakW45youL7goapvG6sm5QUJ6St+/+1SI+S31QkRfUaEvho/v
aWpX+ca9berns5JZ/UyyqO/YQ037lrM/S5q5Us5Yv/qWylTrgmtu0a/IO6S894N+
ykuh/oHOm8j9Y+miYTS6kxXgBArjLUL+xh4SoCxwRSX4CbOJiEMBifFVzUkKiLsl
BX84AHnb2Mq9vY6w9NkDXgmkjuKTDxL98K1WMeaUhog8spymGhqysIOgXUEbrFLe
sl6mgp7ggbzYt72WMwXrGsRY1E5Zyxw5/gft3gKTKMlAz1jqWGEgP5PCinVs1u5E
qxWqKLo3qAWFwk464Ffgo/THWVnwZVjG/5HKHNug9g5cAewS2+17ToowIqH+XlC6
r9vVLjwdISXla9BP2jxsyS0Vxfjl3K5hdaY1PywlQvH+cp2mhTzYiZdN+TXQKDWd
s1lf0+oT1ZBkpAqYWQiBEXJBg6Oqa79Z492ssJvv1o+2+9f89fasesmbfoo8Ool0
9C3uRzje8bSUDKJa4AVAwQuxkkukwSRHI4CtoIW8O0eJK2LFFwUCNrQP1ymDM1fm
ftYJAyOs77+PbaGwPAc4ZvFudoF1qeywVhGBdWWjwuhKDcJQKZWAt5ADgiKn4uc8
WRj4Qs5Htps8/60exrRpweDGpiJ5Kjjmd7HboHcAo4OA6dP+Jh1zoYpq8rVQG8yn
cFFoJ8KUNsPbh+bk2TbqqDk8OL9RXdlrTAq5hBMtl8patEUT+5I8/EtS8e4ZjcfQ
aos7BJZzanFadYFCnPXYiJR1KX29lPJNSTVDyEeuLXjpRKR46eLKe4DFCeTXGxPs
0bEskP78Rq1wfa3SrwsJKlM1gHMdpdqH//fwxxRHd88rKNzABQLohEsPX9CYNjxL
dpkDdQ7sirCfZzQQWMCOIO6JqorA90YL1kwh4la2gszD11+ubOgj8PloKIgslNVn
OKpKZwcCyQMYA3u8rXns7c0wIuvw1i/zHL13LN2tf3JaFDKLrxIYtaN63ufqbrtq
iubun5D546K1RycVCZNsEWM9hRWb/kEVOkdhRPCw370DT8vAzS3mrNKdrJ+WIgSP
zhbUArLqkZCdEbZ9a06SSFi+Y/YuOvWBz6uGOyNQe1T4Ty/anPEhA7PbhgQ6mRLz
MBuFe8MccM7IJ6IKRtOy25WvQCp0vZXTr3itWR2hIpqZZwx4JdsOvaoJlgmA1sPA
S33zMwzvgjtLISRLencSpBFpL+vopnOGAr0coreCWpqepcc3CqAZ5gJyPXYwMgDF
p2B1ss+0p/kTY2aWs0RMhamRwbXVqhyBqQqbSbTcNtCxQKTjrPi7P85NMOMEWNJ8
GUA1Dm8WOSg8TTMs/Ts0KZQFdyUL7w3k/U+E9gKdaHUzHsxKrcJeLAc47S48xQip
W3oSy9JIzZEtsbPmtW/PmtO8VnLrP3voh/RKBaTGWjCC/y1P8auKR3hR23hl/woz
AWcH+eee+F36kXJmeNhewecAWFJdyqzbnYBW/j0y/ZOoKY/wz8uQwLsUkRdTLp/1
SRziwytDWemYQPdZbIhDJvFsZJBJBblHGSxQvnzSgP/MMmFFR+a+bK4SOR6biHTh
b0v64upl4hE0aLUUOiL8zCbxOTtETRzarF44dp9ho8gvamzopgPG6x+tb3hU6lR7
mDicw417+V2BLsp8+p0HOTS8qyjcyT5M9/pXe+qYwsrcJpaE2odkGitaZ8FtN8AV
CtMNEtk9uOZ1i3ceBNlZwuSRhPOq5Pv0rrUO4Lrv93xEuUhUfSoPNf74pFY/qrL+
7CZgo5q+U/2IIN0oSaaCbkAywK5PAgfEFA1pc3H0PyeBwlwrZ+9JIjyNEgFr3OwV
ty0mIcvK0wY79ZMyCPYx3uwqsAbGGFBekRdvo9vlyfCQCLnhm/vH7WGmfLtrX89w
1qS9O4I/ngdbHiD5SO9AeicwAOjRxcbPD49aqyVY3vAXK4S/ic0fIgDC64vS76SF
4NbxyItdOkv0Fx7mDCc+8TOwCUke+QKkA6oQGMIGX+v9opFzLyvPYGj8etQqA57y
8LlEIG6L1yFX/npvBfuntIt7xdc+UuvrGNBJfcJ6m7QRm0MQ1O21DqwTAUfzsyiA
rPbsJwUHChOR8NtYUOy7iCu4Umy+VPl9meCtXzrXnTLQ/SB8FHEkot0EaSRjAlaw
ZozdpHUQamj5BVB9G+7qUiSZz832DaAANTS1BJ3P8D/3C87lpMEKiEIUeTqDmnO6
EgZmC1GygZf+9LqoaUA7jCQ3e+njJ6WMrkOXCWnm+Zk2bdrsBnOXnVUF6EPZ/H7i
vWfLXou0E/jmfk8CBx/fmrYPB6Dy6Y2QNWHKgpmbNk4mBuwMDxaEGxA6+56kuzfJ
DHH1sUzDHYl4kbWX0+Z6dc5gcZkltK7CJEE1G+TF2+JQP8gX4M6rKbTy/wHPT/nO
/p60KinPaTH8NKkX9OIY6Z+xyBgkQGs2jzzauOb6lnDb2G8U3YVC5HjCbeCa0fTU
XdKg5f2T4igqijcHKxaGAsxRKdSXqagV+XYAuxyakwq7aVsy3WSq7OS2Onnf1lI6
p532cG2dqjSkk6Q3w+cr53HB7W7QcYLZBVTE75zthNnqGq7y1UqDEP9pmAtBaYMY
M8ObSSQDsV7mZUdpeTe2iiH/2xQfNpQyFO0Zah6l6cPxVqZFfNXKxEyyrTSlCaYY
4e20yw0K2fbr/rjZ04AWB61PX5JTXjiLVR27BjG73hXDoE/oFKgMSMiAIhiiH0s5
lYg34NXItrNvZLjdW1Dt79ppq3gYVkeJ0IMYvLl/CcN3bxae8KquSJR4BrwKjMyI
2ZyeN52Da5Rmv+2GAR+xOLNhmkMyjQXtQuDJXW1izDU944zsaQqr9SMuhv6zDkCl
yXYBrYpNb60x3ZyKNwy/qAieEmUV4wCcjGAybblDvToItbYwraP2sDKy5Ldbxeb4
bCc0fN2P/khmTu+XwCuZ3henUyXbC2/PUqBAbnu2PgIkT3Yh07hcUJt4PsPUji2v
9S3jKD0WSAYem672xgomPqfnjAtyh5cQxPX4fC8WT/kuJ3JU8WPQhvyRCqOjP0Gk
QKzdGdbYlGOgB2RmM1R/2+qlqc3w8ka8DvtzHItaCqH5CfdS0rg5Ya3gFpqdbcmO
HopdnarGkDuR32wCilnRx3PTVgZmIP0la5rU0QGgc8t4soIqlOUsfkkA/q/0Cihv
OvLhIRu7gb26tvVSgY42uss/ggM+B6rOWnRbzfH1JBwekx5tQbV8YcN3XbYNoOOD
2lawi2Q9d0BUIoUqXba7xefDS3DJrlRp4qjYomb9JAZQj7JW8UZ+HyK0sREnFtiP
3G5jo9w1Djz3a4RBrSBCua8WSD1iwwiTSkp/uRN536mX+AH50N3TV0w4nu1PQD5g
O8/AjY2905Tk2Fguib3d/5n47eDQdq8hLTcuf+XQHNp1GpBD2Xhx3j2NvezJ4OO/
Aci627X/da9HI02dtjveOzlPXwLXJ8HdwcItYP6136EqOjh/7yoTFd18jzIEWOeg
AAybEawLE9Q3ez2Qzau+tw13JM7hMkaDS0vPhe0gJ6xTCFAy+VuW7t+SVzcAbfyK
K1dxwhSmZySYLZ3dwgSFVX8xRlwNk8CJBgDPuMl934tnyPry11Cuvatp2DRIWGvp
rPdc50O8JTTGYBnIJBnhZTsfemyVV2kCdDeiHV3HxyLgbM1KosnVeUf83NNWSPtZ
xr482ENgr9p5etwr69D7l7iQ+QzxnR4J5lL8HPpxrbOGYj0KpMS0H3CWbJi8gX16
OMQS10w48XAn0umb/Xuarxmu7aHF3FX4kmB96Rt52Bx5CjxVyEd8dg95ghkkPrZj
44TqGzpWHjy0/sPRI4H1blyas1t3f8InxAnrwhqDDd1LFf2Ljsb/5VDc77RuE618
hzKWVXSAkhVP+5/IQSSJ2d9h3R/x1QqRMxy6ZsLIGzn6kT/zdX2XiRaVvSMZzuRr
DGsfWaGwHPLzspll9hol3U5YdD+bfz4AVMqOLhvskOXc4ecqirQWYy6tBNvtTLQb
S4tCN2EH68qnviYE2VIjHl9qd6Yq+zOvlSsunHFUPVjSuLXsDE5LrfmMg2sLKUIE
Jt7Vd+ZsNXatb3ZAF/lwIb6Tb6SWrO+D9nQleh4l9PncNR9wNTRDO0Mh7o2REM5Z
nAtsoMJUqP2n/dF6JQmnUeSTvGFOAjXOe6fsuuRJPDGcxxZg9eWc7FxhqL0OxnoX
Oal3Rmqrxp2pUG6tMyVdFndmKBxqcIwJfZEweNN/IVGiC2rnQCEmsjUo1U0HKVnQ
giupsDPioib6c9or0c++CjK72/nYfgShNSj+pwc+8KWs+8iPl120is+P7oD3lA8O
24X4B7Ieoun8uj8cFQyO4l/5No5FQ/19IahTIiw2bFde5y0eH9ZV7t0b90w26woT
BpxhhdHyJ1CGntbuu4ieqLYHpaFduj0cLsl/n4lfxtapL1UwFZoq10BiIlmvYpTe
n4hbqMB3OeP6annvyr+Qn7OOREY/+ZydmxbTfzXnOsl4vglxNz0wWvRRBx2tjZO5
6weYDP0SzfKYpZvDA+YgG0u6pLrlbDxfQJlvYFEpbJS+bRj/yBgEBfmhhuklZwC+
ZJ0vYkxwAvzFr9R0lhNyUHrCKO0x7Os1rUn66XOlgrG1vzN5OxAA2C4xLxJOzFJz
CyClSAm3EUHHKBkAROaWgKaLTTgSS8Teq9sQc/Crjbra/nMjPECbh2w06M29oyLT
vN4Zd7ap2HX5nmPD/vocVAyTzvl4xJ4iIIiH/xwtE/ePvVi2jiGWHKWm+J1tWjUP
XvOQUzd07Wj0h5Uo5wNF0emnlwlsGBEDz32be87rTsRcJGATwB8Q8ijzZmHTPEVW
NF1NUobW7vs6nvccZgTgjJYAs8hnzh9djQ26VK0fN6TU2YBg8u6Wweyg0tw/1hSq
uNSOs+q2eFtOTNBWnmzpChx7BVzRIF1d2mAWm6b9BIgpTa/C0rhLOKOhqaCbPKcf
0tHYB3PmKyyx9UoQJI6eJjYW9N54zYgtB+C9XXelR9T9okRmL5goHx+HZoBwGyeC
GJ1n0oD8db0lYodV/UQk5R6ajcaRgH95GLY6q8Fi2N9IdV/mQAsR+EX8AQDvXr/N
UHtmTRxdFRyyTeDGKFAfbQxxc/jIHFU4gAGpi08U4m4bdd11HSYepfjMv6nQ0Yhw
OdU1GurNUjGz31Asid/juGp8yWLgwip51ASkG4LVZ4pkrsBBK1TbFIR4tEOwXFWi
s48bnnecYw/Lxvu2mC/KLhB6/OyWrjEaUi0/kFBScAsk7r3GOa5/AZ8UkfbFlvqZ
uXVGOrV0VMuaq/Qxe1qmC4LuGsUfGT2dEeE1uTvhsP2kIQXJbPj9WqBFiYn5f7Ya
kdH4Bf/mzO9X9Jw/pL6/uQpfL3XZyKKah1zn6M9cgrKNzTqoj/2SIUtreEiFObou
Dq0tbkBh1fo15nWlTwjm2xqNWPLwso3HEVisNKcDGPN+GqJsOpk1S6+ZVqn0RQ3u
UJYHYl1bLQEyosKRgXGTEzOjyWtg6peC6V0s/9kS+C/RhOa7XeFqX+KUi+e1dB0X
j4HW4DjwV47CfJlIECBG7NxllHqilOXlD7fSKwT6+zaRmzI52jmk9ktJQxJ0NlCk
FmRdxSBVHcoYlt+IcZkD0Ge0wxKXG0Vo4iyG+1PryRvonoiBcbdxKQqlhyEZEcO7
sorRBWsB0jAG0MymEn8J0njX8UgnhSL0P1H2NqruSY+AT2hwDAST3HJgXjhtrn+l
Pqbm6utTwmZPNHnSuq2vamE5k/KwWvpEfaf1UGhrjDxIEy4I+kxQm6ICcvyfjai+
stXOGnYePS8OEfGovgi3wiH+7d7dWH2mx414A10waKBzUG4X/Jwfg4DdwaQmepvU
o7gZV3jFHJh+ccjVCIbXjG2G5JcLheSz2Ba/AYEaf/RyBWa8c1eo37LFak12/Hw/
3OQ7Pl3RWynR5rwJUpGEr9c/YEh2gN3DRe5GqodFTwM15JYB4P2w/QuOvn2onlto
ZmAiiPrdB4XIlLh9egQx3swjA6ExTjr2jgFAO0jwqekGbvKyDhV/jI9t2WZZxIFB
HVYVp0KdHtMpbrNNMs++T/CvXFwTbhponZlrpJX94ZcZJOJ1LiC46KwBKFyBlP1h
xrf6B1UZcrlEcNj84CQ4G/oAEKMZ/rEoGsbkZ/inS4AV5K2zfn72xC1XCJlWK0xL
iYEmfc3Rfieps+EgFgF5UwVF+G8SzCnAmjHz3KF7RkXH6tAua5zvE7cYbijmgDsG
7IIRZfe6WLNpTN6GPSqrAy5DJWsq4fYp2t4Y4hIhrjRvfsYvLf5XX8JpMFh5jyXZ
g21iMa0zHBHGGWa8xfViBPpYsraZJoC9qnKPjh22wzfWfk+QtZR9LVECuXCTjOp1
QW+qJv2KGTauD+SyAVjSSqKykRVz6rO4aCjf/7vrxLYePkSfwQ554nvnmrLZP2FI
y7zeYcMfKQoe07z2aamRfchyEJOBHn+uHk2CSiPRvybRQVPAgrzte7D8Xe6yO3by
x/JMcVqftOBSEXlT7GELSz4SRKHuq3KruHbARpe1llyFBV7o5uFTrGHXGO05KS+/
5NhCeyo4pbxFJolL9kdGH3LAsNfnFagd6IHEXs/PbSOvCZYcBn4usE7omgmTI2Fk
uHgEc6wKSHf4na752n45XBP2dnQ8zbS7VTOxATKGcW7mDG67dfZj04soBVRpDAGS
qyeMRZ76u83B/kunyrQz17FUIWpFBBOIbP25aY+M0FjQu/bArC5bPDaW894A9iXj
sSErHtKesQFIXsUf0Mg+ZRs9GEqJvXe6rFv9IzwF/Z+nXMMPiiJ9FtqXyTQGpcCT
u93Z8I2rMKGpLQukYLQh5RYa3VLk04Oq10IFKw168Qi205gUbGsF5X0hFOa3w87b
gShZIr3QD3beFhcbGvMwmu2wh8JOHkxxUXCGEPKoSkGEcDsPLJLYZJLlC4dIY4l1
ZUvEDxdEkR6bLzw1UFEbVgOssQbFDbNuR5QDPc68TGusqPAvrH9zDSP4v8zJi5JS
BeB+oIHXu2e97bEjbr2rCATWn7nYQ0N8iwWHn2+WJVuO1aKtf4wA4Yp2K/NizHGF
KBaaHxI7Bu3yxBafN/4fyNYVJ8GHMtpiugko7I/ijeP6ZGX59wEK4uxk5JfSRMRw
uSRYx6pG46tZpcjYt1PxYKOTiIMYxXYeXPMYkjwAQd/ELsJ73XDO2LlmiUY5N6fj
Vs0YvmPP1JvQeLAiGCQ83F1OPCZmMiIJA75ZL3Wsm8RK41QOq6+DXy+ztoi5ZBko
d4AL29VKAnHutU3tdeRoYA5eLSr54cD8tderWsR+Gn4/xmON4Rercu8l0wZsIhmF
lP/SlpRcQp/6wT+EHgeRpFno6umekHzZgzKgf5y4mDAnkjXwvHzWkXvQqE+b+N/P
5gLN+Lxm5jvUsLs2QVyJqJKnzIioRTJd680496Z91//4Lh6Ll79SzNnLF0lvtJwx
zA/2MUMwK44wBTiEDHd83Q8oiB+STWVvp+R8KJVh0hk5ln71F3pbdVel08GIv8LD
lSqmBwzm8EuGQyff/Dg5LmjZWBSmm1vcJ9D1I8bBApqTed1P6aRT5o6JtEUgASfp
Bp6IcvVyiyxbe6RxUHr2khkjW85H+bErE46hpDXrOdQZXB0S+FPGIRQscJDha5/6
zheiZ+jMFb4K7qp6jJ5vxJY3bBlq8/hts57Nf6pX8o+cbBc41+yBl215p9SKIn6s
BwLGOQ6CbfPEF5lQlrS3O+M53qjk5mZTH3XSrti1zIIuIFCFi4RW1czZJOxs2Yk3
rK+bAzIRbj+t8by+DLkrVs1WkIRL7FneLlrHFnWu3Qb+DU9Lwbvc+gUvbrNR5j5i
2A+lvkY5AhTLFLcs2hx9qUiUSJXAKsADuUrO/CVp54J8cgZzYHRL3W0D2XJn759G
QZjn877FNqwDNUIbhLp6dboJchWSDljWi6szeey02mcu8vQcHU3elVN5wwscLlMK
O9GIhUDmu7BCQPev+IpSXNQKqpQwbimsLu3n1kIQamOWuBDGWt6sfFcCvYWnuzpT
tlrlh+fLTmM50v5YlPCFhfb0xSMk2ccY5RtMHO/0VvytnVtvDZBqSoWMR1G7Daao
ybOnWmTdphVmkIiVE9nTnKZ5+AbqB5EMrGwpLQKXGjzAD8MpTZXTUGyC+E9G53if
W8YDEBNiqaRePfPzE82KoSrnN12l8cquv4uq/obxyWGNmFsd4W/xolu/igZND0HB
NajEEmnR8Ir9GeRDp2zD2NsTkR0CQ8TzejWHC5bSb2XlniCNMwfSSMkanmoFaJmU
n8kT3vZ6POc8wVYKGkCl8bral0nOBg3CuLCI9PR9sPOgPbk/zs/+73/8m4B8Qkcc
o6d8K+Mwinb9FdK9UnBv9NzZ/a/Mm2wcB0kL5nYLSwmYkKRQ0UbePCseiHTqdnYG
sA7/ly8Z1Gl9bdjiV27Nf+UY4jrU+IMlS3iuZtDGeS/QjQ7nndQtBCPaojntIqYe
upM2d4MknTiZnQnRbFJ2bofIrZc6WSi0s8Uf19etaSq63WNkw3SxhUVc1bbcZFVX
fB8hry/qH5yBG0rg5IpeS/IPv2ehY1EdIT+pXpkB4G5sH0t94XMAbu8OtkRi7Nw+
qvrN+6LCmk1Ru5Ci44aGouUSVapjjvhk8IP29jb5NwNTbnWezJDai7skaVPe4kg0
0rQhfTNe6KwZH7UspMJuql5FcNJjM/EQgJBtAzco9K6o5ukPlpN/1pZwQ710lNvi
ocamdppqhKKOKhgFj5jrUuo5EaUCSNXaqB3PZCQJSCqHlPCWbAGRV5Ij1s+ipB7T
nC3F/isrdn3/17G5Cgu1aNbbMCXfolyZCZ7C8vkNBnjRNW4Q+AqNBEzZyrolEE4M
xbt+ljrQlahLBCYoB5XqQJ1KQlxECpkK9vHSoBqQemSRw2NJvmVXahoPqWn6VQzc
TFcK1BzPa3IXfO4QshiPPXZK3qB6KDLviyfHh/ym57AQ2TKy01ZmyaV/odsOnLQs
dzbBjSnJIb75G5d+WFsCi/03p5g2AA+iI6SFCk1TCPRyiPG4f2LShOW8LVW4dOln
QTkTbT4ylmFCKwqkKiT2rx9Oy3O8OwPElkIpw5uRqO15NwESjqJ658qxyyYOBQ7Z
X+qIWTzDlTOtjLKM8QSdNsKcIDwSycxO7JbEn5JOsy2b5zRpNB/AKTViYLJPOhGF
WZ3h2Gjg9mt4ckLWnz1qfw75V6nkMMs3VMm7P18JmusHVb5vA1BrN+DzsONbZY7W
fJ5VjYIBmnnOBqhe68NDb/LX9gzibRjbAMVcJueimUhr1vczN91vU6ILxsgKwy8n
RGHKcJV8/z3FxtGnTK9Q7BnXXx6YVTv/McEHaxuKOSM7/QxPDUNZEANisKTOWUWL
65OjFhh2c9oYUVmwDL58mclQiexj4ggQOA9RrSTfJHy2+mb2XhYYFVDgqopC1r9p
ENMEwF2C0OBdGIgzaQ0BNQL+lM5/Jzs2/9+UxAQRjuU551J5fzuX8aIxTg06VIfG
wsO8ndxrmj++JJFGpJ0/GuTIscenc7NaH3u/vr7ILhAI1ynfazTJACz3zcnvolQm
B2gve1O4vn4MD/TDYMZ6d5CodiLZPTI5s3VIZ+cqR2MMVntqccuHmWO5YrhP+2P4
6QS6zW/dnr7siUlvA+JM8aqwSjMMC8eIDERQJI12J7RMKD/go/ZHWHhhUv9VzEjH
L6/zM4Dzo5tb7tMbRXtDYVjzu375rj56ZTDeXpB/0yA7x7q7u91fZagVJzavQCuB
XKFQIFi0PWDC4F4Ix51i16RvgJzuGTqYOdbCcNq1ZFaHYGxgG2MjJc2BtywF90Zj
ImHuAuHCaAEnC5N9te/7JxSuRwZ+EAhcaG1bFVYOF5uKcMhJrCFB5M4nl00XKe3J
NUY5iNCHkeSygRoRLkSeKcXYBLKrddrkC46f57ojly530n+voliVvgp/t0tdFBId
h4/N9pl5ywipciskhHIv93CMrfxxX13qrPn/QA4xugOGmuQQrQkzDosq0OHk1eo7
O8EdA2mNzeizacv2sw96QcPvLs00xTO7YB0JK4Hwrm2XTO9OlG7I0FUlDeyDvPw5
u3ni7ddGkgDfIHGpNB5TWiz9vh9k7ShUEixWkyC/C5+J5yYWEXXStFiH827xoozx
4aAdxWE8YzbnfrKXLhXGFtN8Ldka0pgG1OViUWjeewvAmwAMIidxS6DFoz/OZuim
0D8jYUfGrAGjw4D6CQ5aj6gtJCrTujzN2ZqbhKDC8obbw5+JwPcaGD6rv0x3Cnmp
SA4Fucz6+m7Fb5XM9/HCztctwgvfrSHohCSzSSo0L6ufDTXrPcom/PJJgCLHI5Uf
wE5eXJxuSRbRhuY0vzOpQ9kHNosO0WzsPm9TiClijFS48JftADZ75c0UYRCuiQ0W
Y+5A7WI9M5H04vwenwudES2sN31hVojcHHiLfv+mFHqw80orFdTaXLhM6mJxdlHr
9OpemoYXy6jYcjqUfDUi8bVYvWqCCvqB6y/IHFEs7MlUFOOsU46MaV4dAUfsU4KV
XLK0cIyj7eY05JWUmJ6Zl+BmV1JV6nc2Rf8BPM+jBfNbq7Ymbs/gkBDbMWPslaAO
ee4umKcChsgQuKQcjmKDlrYne9aVWmWLG5D4XZG5Q2PeoDnk3xGp2VWH/D2m9zMZ
EaSwLAFSx6TOFr5XzVLoT5OnAVAQ4b3uXcLnP4ekChFrFJehN2F1FJ4NTu+9oJxA
No3fH7X303kT4d9n495j59l8l1lwzs8uBAMz1YPk9fByflnZS7wFz2gYBoWshxvI
7hlbnBfNRBeLhx5bNmCPpLtOVVUrFD7Jl28V0RBcT8mn9hWaBSaasmZD0Wt5Y4U4
5Elyf9GB5FTQmWgDVrIl/F46lVpSULFt+l6HDBV5cPlJ6pu30HM4T0ejr9UKSq1G
QHIApkR6jr2IMwXsmYixVafKVpXOMFQ0jzQ6ttAdJXB/fh7Stx5tXwjvfNUEgHU2
OiBCqW40vuOMwW/UP9Sq1gTKUGqME8hW1j/69yNyUbVEZIMdJJQg5NDd0Hnnix1G
xgfc8stFdAbmZ29kWXOwpL8ik93CH2WmRV/qMOrzJf4hyv1CQ64RV/8dVDERbfOR
YmknXHP5zrzXscmJAzZxRJK1uwSmfrsFjH8VkQrn/xCwzyzeYfObPudP5qe/bzGw
H+nq8NuEI1g2lbO26JNFHVL42D1i43NZVBMWBkDYyKPw6WnKCSQkTx7/4n3iezZ4
f72pj5XDIggn8ceogXlagNem4ktrHiecv7//K2qkYQh+1qI/intaj30BTEFTbtbY
pN4tNA15ErNWur3roueYMfSlrJvnwSdCwrV+vIHDBBoUxEAZItZtIGM9QGgXG/9d
EpMwXJnJQ2PEe3yUWx2acxna/UH+jkS3Lpmn2FGaEtkmXOpqoRyI7j6iMhKcMcX+
XObKkGXCKYQbDfDJCdOuC/Yk0Y12PDrziQBsiHQzYwjkLW1EixJ1Cw2JH8wHGv4R
wzSlTjhHQmgPnx2BFJqB1zkZUf6PkRrZiU0N9SoKN1Zszm4YwKpQVS8l6hldT+H3
WvPbWqojV7dJyEXO8f+D6H6/OFFA5bEjEH//XiyJiPTH/rAzH+tCCWws+u2AE/xU
RmcTnSLO4vjX4dM2yitaTsIX6g6vaAjrZz8gzLdAGXvQmIuNBk22ONh3hnYsRSzr
FLVBv911d0PScAW/p0Qz8NwLwdAN6cijyFOAF8zj45h82PzZiP/SC1yenXK6yXY8
1XMLmCe216pBT7M6e0MuvOKjpfz4Ym5QyZC46o9lfJmn854hHRu0EQpzf97CLZQ8
fjDUyCaYJTgaw24IUyxAP4XA7qgsYLtrMc9CuM1OhNdDDrFND3OmM6AN440Od3F4
abMMHxw4oQ8NDhEWfF7+8NxW3rilqIxjMEEh08XiV0NgJt8cQkdK/vOrmoAo7mJx
gDbvY+Ghxzy9mOw5pOJiRYb1OFUxL35/PsfSmFReeYuwl6imu78sMITFUxLE/pn1
u8IQgkgtcsjFfgSeztdN0amXvPdx08Ov9DmEYT3jKMrqJ+drnp+KybzQau0wYG5i
8NxZ47Bf0rr06YZhs2mbqaPHxQ/RfZIEVWyfRGcmToF9KOc8g3tAO1kWGzohA8IE
AXYtVmHPFcG/3+pXLeJ3ig/CAI8/xZ3cqUc/2AwU8xnC/GPT8Q+wo3ABKNuYxHLf
RniT2BdYtcvcbHWj1mz58eg0p0zptukYzmFL+JKGY3P336BYFQR4OQq29LoTcy9D
IMwr5lZPyPIwLvM08Rg1cQqy/rCiZ4iOfTE2mYU69yZbRoiD9VBg3zKqWpIjS+fO
Vq0FT1+lTdhYkwb46tkthr8YLpaifnn/JxN5IYf2pAMNSb4qDWbe2siJ+eV76Jae
A2pqNDabD68TU4J2D0oWDp3KwNSD6sTFe6B/v7+lTQKUfapuMSVh+8ES4JggASP3
3bjnK63dRLXldkxWo++SOJ+a+HfW+ms0POGZd6ghubLPVXLbvwERIn0DCSt0/plh
+GbLRwzN+vh9Kfw0m1g7hhQvO8TmO9vYD0YdZnB+fXMk8nS38QTa13zRYlTLpgWL
HChXximyGobm7rK8MGrjrsvyAC6/m8H2x24Pw0ZvyyAcuEaxnQDD+Dcd0jdXJ127
uai+/jWAXovjUHd1xf+yCHe6lQASCr0/8eK95ulQCxidT6by1xUaT+4H1HB2WP+l
GJ/41xyZEeUITuPglY9v8Ycy6udzjZB5qYaaHsQSIYEiJNEe6vw7LLlHRv0UOKR/
Qr+oa29G2TjLauMCkxfjVE9xP6l+75a2iaPFhSTby4ZVAyx5S7XIEQ3vD+MmyfxP
GRm4qW5Z0XT2fjrKK+jvADIV+GOpAqsd0xnnLt9RG2ekBMqCyjT2lDU5pOvpTZTK
xQOyDg+D1DwAoV6FaNeYALShXEvTMYuE5rue9L9yhdP/+ZLEXA+isE8kvodEsz/L
QtX+4R90mDH9jb9e4OFm7sNKIx0c4rJ0FDJVr2cRfM2Usabn9V0J1PE9vuXVpo4Q
cjruecPC1IKX3UY1wSEdqKNeOOkuYRixPhJaQscIbGXNE4pYoygMOK+khp0Vvko2
ywJXpBkGJgMxjouhIvi74YzNsrzxXLQDYzET3u0BLcfCW8wMaLgLhntjNPHqwpwn
xTcdfQIcTIA6CtFUDb5E+/nh5ojp5DH8vU8NRryhOwdAdSZyL1nux86LSu1TTzo0
QKh1QfDxDujAgE6/TRq5cUI1Y+X1O2QXP8BKfk3sV2NovNRIUKo4cNdnoNyhAffA
Cf3wyJgPqL18o1Vg4iI+U4Elzed3tbyxxWCgdEQc/JiCTIxdtEfjRsGmmN3TU2F6
+gQ5+YdLLdcgtVBxn818852JO7pn9dUPRf6NOAImE2wZRaRmeJfzrmEXNtUu+Ivu
m/NWYM6EX6D4WH5aj0kkk/y9igpVEg2b9tFTWma+dlUb1rvmCq2Brgx5bVQHf3iW
ou2APcs6gENoAHBOiY+XZynGjcw14BMvQktqmDvoakxzb03Qvjm/ZIGDlbflqj+7
4TJAfd5bWkc29ZVkNAJYGIGc6HeGHYe6FhJFT7d/6/Uhf9qcaGFUI9IuUoI+uSr9
YNT51eocQawCcyU0tNPfpxdekYb4/XfkltCkhhWYz7od2HxfJk8JPfVKTT0Mat/u
ECgm/YNYnr1aovcGH0WcPrOJ9E7F/Yq0NEYmu9iKc56MMKlCOjR6vjChsw1zwrLE
mkz/cGuILAhW5AdSRYTfqlxm9/ZoNx5ntKi0jKDWTdACmW5WPG7iavhAZhTzvMoe
tGswq5ihfgYwVykbV800eg5ayrSQXuHQ1qbzDyTz0tPzgeiUvchWKLn0X+w1aMul
PChdh/RUNYl7SS59MnRHbP9uCpGuq49p12ian6xlgTomF7isA1fKoIqoBEVCIGdA
Q+/d2aIst0mwF8DY5NDmVmBDxwJDnEXW/GX9c25i56rfZtNpTPsqU5xa+RGM7tO8
rVb405+GpYQmlnyFKnoq1EDM1tZQfyAsFO5g+gwTCMMhTLWZ/bwmacEiuWGMHLMH
B3gtnL3wvugelLA42A1qoNi+5JteH9V6IOFM8aZnZLsqwcBcuhFCG2o8qv6RNN/N
vPXgr6NPCAbFcEa8KdzDE5udoC6NVjycnxuv95goatZmJEb26vznQ5Kz9x+Rbu8a
RIwBkj3PXBlVrVnPoK+sCXdVJh/yu/y+O3mZ/NeHzFh/TkhHam0XyL4h7/pAVNsi
82YykWTY+kekQg7yR0BOd7R88iefa8dtV/NtPBNzXEvSvjY//U4eYC3r1x3P1RRh
5pXT6LFJKLCqWsuKDbLWAkRsWH/LpYjZ3rKIuCu8OzcKJHOWOCRTWEmTT32nxhNQ
tOO1UvSVEk+WAjTj7LYCnrN/of0AAiXacZuZiJyHsucPkquPCixW4ZGyrMehljVJ
cqycJDA8QFWfGoLsgoJaqwpeFGAIBZGtF8/UP5YQxiB2DE90cfvdiiE4uKGNnu8n
TFccqvxTpGYvm62fht9VRm0xzEToB8V289/RWjGJE2JXX8qUPNEFRV0xngEWbt0N
B0uXOej9NbbANbykxGojkhehzVU6Hp9f9srB17m605n0VsRblzgMHWcZRGZoo3Ex
n/YvNoVa2or1Dt5gEzpAPNRuVKm7tkupkis5zRUMh6dPe+62lH6cNCOQ31KXZSLT
qag7T+8e4BakobTkXojsfI7K56mtoRYVDhE0fjPDdrKMAhy7kgnOodCkEoHh8fRP
gZAAWgQb1cxm4Iq+FV059iGE95oEiQg7QMYJ1d7iQqhknsKTwpKZ1uE6y2DhLD1Y
DH26ZEnKK5qCow+878bfmm7boaDtYL9kob2ILo6QGpsaD17RgG+mt2gWYtT5xbBJ
bAMNnJp8VfNzUg0XTPvLazlr+V9WUL+MFrY+tZt9feAdYGTIqTOroA8vYmoGSXqV
2XIt4nLDbaBjReos0XBdRpkYC9CaKw2CbQeXRd5wcJCJCyfaVGti1FrJZgytS5BT
NB39fIcqf9k3xHoX0cM9rqGoW1BTnhB/PfFHkK+BY3Y/EFgymndIB0rEPmQGtnD/
EXpN1JZ1iu3wuj6svNg8JhoTYxTJqJVqatSTI/Rt8PHNfVt96pK5BInk/u3aFwuo
0klC/vxnUX9eTRQVUDRRqx7fSW+aIfKGSmqgrPhRQKymtkVStfvFPH7/et6c7J5m
D0dvbJe7HQohOUSerdX9rHpVOkwAyRQ0ofJdmlwjgH2FtDImTa85qXs1qUW6+ggK
RXxVxosSAAazwZTosFLuaPr7FVk0EXsYvr4i+uo49Wmg2Y40b4+8dbOAhoB9D4Fi
940HCoAdQ+tv79uVQ/pVgVI9kwoCyXpSUkmDi5me6Ew9QhESYnyuJ1slCnVvAluc
zt5PWdJ78VnXNkne+G/UWIKnqHims58TVERR/XybxLrSSajtU95qLEcgPhZggE6+
q9IQOfpiPQFdtCb/A4YpadOu8eUyiEfttYVfo6Ra3tXadKzJ+xM2BaNSsDa6pyYN
mm1ytsn8CqMusjS7Xz/Drqgiq89Y/q80ILourHZ1o1zwLVJXZtIWvdr4PeaLAjc+
zScX0nX4tdKaTvz7p+jZ4/Ifz0+ZgpT0Gr3bBTIjtz67y4sPq21RQs5t6Ax9VBvY
vmf/XlopNXb9aDYwS9zvVq+4JYwm2Y6VuDKBLuixVC2uczkEwNVRof+vT/V26iQz
L26z9nNXp9R5NSigGIgjOQGuzR4XJmbeVbzlGkcSvXLPLf+58K0zPYwsUS9kTVo9
ULbUD4D1HMxlFVe5AA3y+bp8H2JQc7WQXIutGx6eEiKPTPsNFBaWG3GrPMU7VXgc
og6zxskUOAfKxVxVLlX6o/RllfwsHQVl14z79v4cp1LoF/69GYly6MeL+K74I+BX
Fd7QMfm0+o3ZEOW66nxBEB1QAvdMvDIglhoFrn9jBippStIVApoanA8B1wNT2UIR
XJ/1BhtnglOInZ+hBm9S3MCM/Nik1nEUyvVNE67/3/EjW9MhXXWGaWequma8OEsV
rmSzibCWwLHKJW5F0glYD7HIVrHD5HL6o6zQWRY9HtoJR4FyQ13lfSVKkToC3YJr
c7DGmxSY9QJtTVf0G5cDw299xpspdqSg64cKSfokGgTA2WfGwhLGkUGdiYUB5r6u
0VDBaCL7jpZj46iHkUUEwMpWVI1eTNkF9Y4ev7VjS1PCR24VpmyP/AtSj/tb0gr7
KV02nM1p9OOdwyU+UP19P2fPVhIlIXxweQMqNp0n6LLh2tiowh8+yTLUesPF8Tus
ZT+zJcgjWWeqZ/cxJvnFUEDWf8YSYMTl8Z+UA7TeWeetrO3zIoCggJrqlfW6qEtO
11ZKjDHApkuXDafKZ3nAGOsj1ZjfBlGozvRuiiDbQLrYzLRS7YBuiZDfYQqNeU0g
xGiMMBQPdyjdqbBe/38riiqhrRz6le0eIZiKPm/7RSM+vF6hMRrjTfgUy3nVjWZ3
88AgoyeRquqLKlnvRsNy2olIO8Wg7z0DswWO8W8LTsYTdvdAEspd74LtHicGdbRj
J/i2k8SQoIMKkjxXy80aNJn3J3qtZSbxSYcFTSwL2v5cwFfnR2RRKMOoLMMhhraQ
o/xqhbwj98utMZGT0ZRgVZyETp9aI8fasMhanda8ZEJNInkZdTjmQkHgaFHKXZQn
3CfhRnv8XA9KJISUcAfJ9B7JYncUUEaNE6cOhkGC+GdwIncoIXC+XfFrV2fWiwq6
2t6Bm0PnpQ6Eud4ZsNCLbYYMduCS5dgxccWPnld19MuzDzr2ADMJUGOEgXv078YN
uw4UkHjziUWEPcbeIUwGVtMfLTR/F1NEBNP3dC9DB+n7TR/l8GJdOF/AUx474Cop
9M5b3ZdP7Tq0UQGDpTp/m33luufKGcg4kZgx/grfyXE+oIKzB/qE2kcWvH5txwBM
gF2/0ZTTA80wHMiHgW9gXA+sibn2TNES65C7LL9iFfxtzPAXTiYQrRMODY5knuCD
hQ+/WLqRnImuEo2goyhNA0wsnKSV9eXEHbr/Bdeph35cxVh4txnvdY7Z83U8aQgh
t/rMHTAeT220c5WjaU51uySE5xSeZuXlsGR2bdFAQHI7nQV7HtbFeJNMvWuIwM19
MgeRohbx6oh8rJV5RR6z+H3YEORkCzZAhxwdQVoXDs0qLj9rKoDW3iG8ilbTQuwe
INjgEyF20tkK44HTR9+G7Moji/eT3iZiJyRmaJwfyt7KjfHODJydhwUb+9wWEAf8
nASaMwhmWpEk3UZAu9pHE79ygQFhGITcB1ErlYStCIZzMlkNJHAvRkl4L/5TQP3J
K33DhSw5UzO20boQ0g3s1zuFmFOhTkkN8yvdgfhPOrr43L2Yk6rkSHgmqUCaGIk5
cT4CkK3k/M7gW/UkecS4lo2nb2E7CwYyCo12Q67+TAoxn+86rDTs2LqUodG9A22K
P4i41VOGTv6dOZ85mnGY7EAz5IyaT1XD+8pQDofdDrmC+RrZiZit3C2lheZRtX/W
uKrHvXT1oANnzboXN/o7AlsGTb3PKgE5wz3Djy9gwsQ652vpRee528+eLHl8/y+d
salcVmkMNNQrRGrinSpmAUoSDNWPedcuPeWrmonOWtMUjXkGu6ZrbrhTuvApigyP
nQRc43WTLbBbawGPe1fgucR8/TMCJ47GMI4GAI8sq+c/+v3ev7/OcXYZjI8VkQOl
UO7IloHqS/0t8rXTOlrGniTP+Yl/a3DuML0Y6QVPaImtBXleudsZ64qckkAYhbh4
2M93mbWXxBu2rDlMbRa/bdG0RhphfijEZCjIZqxtCwyoMjHAjYSSLHFhB7ibcEGQ
yzXEV5kIhjAySgkbMTzC1F80iA8/6D1jhZMEzrRq/ZlBwkKLfjGObS5aAprEXWlM
XUspNhArKi5FBDNIjCPyCOvuYt7jK8k7aAwVWTCQa+ZYyMrZy3ocBSdYsYlAiYXC
nDpLA6TrRNSPiBc8rueSYWyuPi5BNdETjOxnktJFP5yCkOegkO8ziKuQe1qk6EBr
QGb+xagzG4t2l9C609LVzjNGiLYssjbZ0B9gbo5yhoGOFHg0wrdEgsePNqakmlnr
4I2fpDTTAtFSyQ7CZXmH4pevIFtjXJmdi+use7d2tjytICm/aVoLjre4tpJ5n/XA
P2CgBqbTmZflGeH7ky6tVTCeH30+c8zrfG5fCXqdP39hYVj7E4PIWk/uy7F9p/JY
S6hM9u4m6OZu+H3qc026Q/WJlIni8iW74eceXfy+YPwcwpwZnVX1g22H1OSyAqcC
BNjfznntgy0s/9ejsBp1qDuyhEe3bPJOojTz4IaFGuhY7Xt+dAps8XnsGG+yajX1
eShqbdKG2MNn0rzOWT+wxPMRu0wRz9AssPTK459/4/0cHz4UHEej4rLlBEKQYXKj
zBUfQr38ZlB3huWgHkZU2GofNjZuXa71WBTa1D+/J2nMCakeXemWYnA8qpPDL5En
VPvLCn5hFDoYD5rMiviJ541gPAlrMLNiY0Isuipqxbs5HbnOd5/X3v8Yj+z3cWKY
T4KE07HesaMFfjUUxO5Zc71VDxf04lgB+m5juIaMDNkCM3Y8FZ5Lyu8WUfzJUM9T
7Y+tcWZnYSd3lrLSc75hEYqUsixnvSAG0mMIuUWd0Q7w4HHqtIGjDn/Kg8KHO3Vo
UD6jGVb5wEjoZ3spJP2ihFUy+d4zcAE7LzbmHNj/2VR6DCKlZUN9HxaJf0PyaDcH
3VZ6N2b3rcIzCmXhRKWCmo26gTyed5KhJPdiSuwsrEgod8HIdR2rn3lJz/8q6RPc
V5gCmQ+wZN4UlR/e7wiH5Lc9BduZCj/igikOTnBy/ZZJd+LgQCR9GJbRdffId0Q8
BOfQaAUsd12g37b3axrFN5FGMjX1qkYXSHMZK/S4djYpsXG7VvHt3mD6Owt3deKg
83vxc8jN/Y+fuO8SOAtqSYYFkb+qXmkI31qns6SDoF/4iuoSQhFgauWn2uCqQYcs
RwV1LXspiCn3M7XbAp+sTk9QnUMx4myJOJ4IqB5NR2a48RCGuXJO6EXyw8feW/8s
f0pWQFck6lfN320bCrhS6NbSsz8ehfvqiPbPdxhJBn67nestXdttx/QiApirdv6D
URyCHCxDEibs751XdPFgD+MwU/rjBirhVGSuc2RsfskDlnlnt1yQmJoHpS3IwryX
ag8XMHwS7qcdOTe5Cn77kdoCRcexgmEDqf/4oHniz8st05dyKGdD3PWeOa4SSUMa
SUJWcVKwsIUGbgLyaYz7/vIX0yJ16RxqIgAlMyvXLV9SlbfooiLCE360wUJSIrAI
mWrFbTCEmaYndtCDP8g4nAM/rnH7ttGsjNlySbSe80WR9fCA9frBofdIt159UQZg
+9PKPCi10hBGOQ2Z5sQFPXhAPhHtX11JgKeLjMB35yvmwZ6IadxBJ7i5V2xMlk3n
YZa95z505oB7FLCm/r9pxoSsYpz8TZbsx3FTB+TEicjBQcgnkYGvFc64Wgsj6Ani
6+uwVrEqoX97X5TvfgDACFQQwvj03TjytnBk873ySq6Xwa1hjNMRmm/NfvYAGWR8
IPDWus6cRUY2vYNOsclV+USwlsoVNMab5P1OL/JnJa3lpzecEKimX2hDzjb6VtTu
J+plBy6mjm8wqea8c8IW6ABYpbTN9kvtq8NKQDcOh4evDPp0b67Ma1mBNCELdyUG
cOVaN46kGZBF6f1aUH+bWF9U7TKkzhTQAbQoX//56NusGfeB56+AhS5dnMLwPVF6
4aPS5n+5B7a9Hp91ygLgtuIVsib+e0V/VMjQKFdwwJhszaTOcBUOcFPYZGvJ9na9
A0NViQ/VzIcaNBOJlJjFPg9i2Zbu0BsAn4sFKFHVYH3ymS+0xua5MSqWkngprt2l
Z0D5L5P0ipfmcfL1DrYt6Q837tMYBlL03cG99duoVknwJGU3rA5LNL4A4O9Q81Df
6hA2Z38jf7KiaVF+lI6KcZ2bWMeieSKZ5hvJ1EZvh3zJAt1CjUndyPN2GN71LP+9
MF392Oixgnu8p1rKnPkayEXqe2B12s2LIbicRsm2udU2cIow8ncgk6oo+2K/2DlV
oJwaNNSJlul/fNP2QTc/PdiDg/NHxpAVXUU25wfzvpgdUV+jR7bqdV6N0GLIUmWp
T0VRr+iFQSWuof3XFthq5mK39qqadjypspWPgAj5OwkQrM55KY6/8tAGNfFiJG47
PSSaq08K5iIRfwhynsi7dwu36TFxu8ywNPJSNSMlNFjgoO1x6sifB07MHr+UQaiR
KWIwcZUqMITVwDs8QXf7UnFX22Z8HvH4Q5QeogocBJ3zcXxSC9+0VF0GKRNERYQE
UHuVfZUZChhWS/C0/wUcbtgflJHE715oxLw0BfoWvKARHAdG4MFz9BNMJBVXcyyC
eHYKh5iznSRgrMtDLBiNOvVr7MyQjFyPoe24GKYOXCimiLsJlLc12GmaAY/JFvss
L1yOKyjwEfi57ONwlBHFraryP304tvWmAKTYoOuKzF3+qwiXQO5F6NwhBgzetkuV
gDZ4NGCI6u3YJPIxdkPJh2RwYRR2rE0TfH/X9aCTehiGt4OhyeEawZ+krMF6Nhay
fAUXPtVCNTcV4t9MqZ+D1XZC3OMs6LnH2cuI284lr8mmuWzIsZ5ug07Q/USjjISS
XeBhmXnHUMnF09vpKF+87v10Mzd8AFSzJkwcFplHhm3enzdISAYRb4V8hCKCD0mj
MpXw/+te1ETNeaPTi0I4iSGmWApr2SVE/Wy3PldQ3UVElG0j5SLaGnmedMM11QX4
zik6xRGxJrZ2Ewf7ElJC69kcoa3f5BRmWDKYMudKyghsZwOwC90DHoyjLdWuFO7H
DU3j3y+rQudQsRcT+lHGH9PGIPr4YCs6FKUnoD9ba2mx/avlOdfB2BhXsenzhYyk
Wzlt//lT0qxTru//6paFtHx79RcOp9Spv8nyaJVrCJVUByFXL/1sfr/7rZ9p3ebU
/TsaScrFwb9EJKsLopX1151rilhsPQ+upDyysqJhVTkChHoYBUcfR3lPxl4B39x8
1lNdzQhaPP0YbBZcf0a/F4+M//smQZQ89W/0F1xQ911SDxCDHGQKwPnRzHY7cvqu
D1+1hh0i7NLkOS/DQAlnEkafxw0TOLOP0kUsmEmcbVsiJjCGsqrrFaZfMuyl7TMZ
ESh8jubHj6hiLKv+CJZ2z3J2BlZmNSRLiJAdBJ9NoVxrpGgAQR6Gwqv5yRBLSOB4
TxVJCqKe8UkMlM+vFAL1SfJQsFtO8BySR5GFKzl4c+8mEWTBBB/od0s3cwe4LHE6
QxvhXdxL6gYKN04JvHl+ePv0bMdWiFopWrXJCvIgXgI++9uo7FdWWEDtVuLNmwCI
Dz9irygfN+K8+Bw+vaRcRYp9acScfPnVcB+E0kqWlbc3YKm/aNwXHHwxg/Q+05pA
LI5WGdI6Hgzi7iJ0/UX+lQX6S0L47bvja03jZ7nMSk/8ECQMTjHIqn8Dj8p9xTJk
YCCXKY5eMPQhNTtQS045JFLljC73IIppe2PrnpHNcIdtxMUjb0Y1cyCs0276d9Kn
ZacGn/CaCh2NqXZeGcuI+g/xy64AXknL1GSE0b2evZw4BNBauHoS506zrKH8od3L
YttMQg+ciQnFT6c43R4O42eM5E1mHmYL9r9RyXurXZUrYXpZ1ecK4ynj5U1u5Thc
rxJdEZfiLm3QVP1xm+vf67VUkdeiC0m8Ta6yqZMM/hzdyVrRIO0EoSRa0KlLN3QD
sq/eL7c6sauMqPXnbw88d0EOZbgbeXsoHrzFzlbNyHr51HNQKrrnX6uKC72hQ/t0
7CzdnU7B3y5TakXTwiBxdo+qcWcmPNwkJWWO9SUPKwXDolEZXQQXnJo2ajqGszJi
xLnFCBu6NooT05Jx903cnJhSjMiNQCe5PQmqQcUo2FfAXfiTvN4vQLBHkWbp9duv
zc+e97m6VymKKtchAY+06dYQW58dfDp8ajPvT7ZD6XJWOV8PBiBaZ6saqGV1b2x/
Ar7xr3VzUYlX0SwcycCYAcL7Sg+SyRZViyE/sPoBrh5P4bKtq038VNkd2fNLiMsT
URBPpQTwtxzo/BZ737NQOnBlCjJMaUy8YeqO1AKdg1oth3CZN4ePls7JY610j4A0
eyfGMAsrPd1OZM9XdCuR+fIa1ScwZGAL7bbnDQK9orDW8E23/Joo9KWyJHNWAVWM
w4ZSeHzo3QNvzM9i6NLumXijf9RKquwz90WpaoVel+fibBKpA2uUlo1KsL6O6eae
JSuJ495OItFRkUM7qceInwi9gmEfcmcXYFJ3GxklO7UUAYLk0DV0aMoPykGLAAxv
uQRxDr2gikoiiweFYqtkmCqSQa1KkTfodW45zwYmWzeR5yg7aBBjfSRqb1VH4ddk
pnBMuwnEK/TgebLjAWOETStoq5dBK9zA2kcZfEccO4i7aPmnp++7MM4fQi4hrukv
pM3oujDUtRTS5klTZOjuM+XjRxOFEqjyS6n+i3zfFvVpLFlZ16uDllbCYuUgHKfl
kMrDvCzKr5KtzoWrIi5/pi8vwz3UcxhBx4exQdbJrLy1UeIzHaU4tmvR4TdtnjEQ
9gS7RktqXOZkkRITiCvK+BEl0cEG8DLcfa021gUvrb9msCXF9wi+5gside2nX/zC
tvyQS14LerfQb8QCRyfH2uQCi0AnmHGOy6mIVtY9MY3MJRDOnXU3OEC/7YnZf8v9
Z0h7qiNRN8/SCJ6oelZxjLBAtyVu3dYDgyU4c4O8W0L2CGeUDqw0/CXhzHMuFNUo
4gRx3xFRkzLRgOwGifNTd2UEob7jJA8/sT1y1CZyCuvq7uek3Ug78S3S/IAsCfp0
oI5gw1MGJmWBQpMjjJmwMXg390bW9u0ZczoJD9AXsDqm57eCzntqaEjw02lDqx5q
584HMKfndEJUszogZaoJ47cGhDkts/CEgcg2K6UOh6FrsIwQ69aVytkGDwwyZ0R/
s9fdn1O6PH8OAML4A6pLZfSgt26H6O3hEnogYnKYB0qZ33PPo1PdKDvCqtISRCUQ
qO/OuX9r+cx75/TR/IfzDNQt6qzA/MJ9P15ZDP3LarO+Ca79DcHfIYp+qBau5pxA
9y8IvyNTOKAtKohvcqXxwVackDFkb1oa+yfdWvGtF3zv4gjLIkbUSYV7TO0QlhCS
MsAO8Qw6Gz3NvaKECX3aEmsw7nemmd39lMK3/6nn8Qw57/pDz2rX0wA/JMNpXPHi
BhASOOVJrZn0ul+XUpi6W+v1XACcRGQmxvOhocmno6UYEO0DO6+nm9Ksgv3bQXe4
rSdoXNjoZq4yow381MpTfNeXlrHvarMsJtKsqNaJmicI8Yd/sqqxCkLlCRBrJFBS
5uSDuBO2niHFDQD0a3BOOrLEX3t/R0ORu99HfuyyzWck7THb8QWXB2/h8EKzwcvf
5+nUL/dSNGC4kGGgxpwBAas1PHnH9+RD3me59W78054EdMRwpO4O5zSHNc2gtY30
z8vrKGAS4VCz6MTl8tX6yR1ktW1PZC4xaEToXY5zYGVFsCkOfYKuV5uJs7VQGoXL
i/0kKxJA1omwGu8qzWVqdWCfKKYGX+iU0yD4uMH8BWKQ6w077547zxX4Wr7+xJ8b
hr/kANK/mKh+eqpHYRZaY2bccwngxAwZ/Msf6zJaxARqjcfVCtYEUxgj0wlklbqL
Yg5tdjKSRc14OjvWwDwDVB0dPLCd0qFU66B1kY0cqTcdhbKSSqTajeoQkIp+QUHt
NA3RbutFsf5i0N3omPZzwbEWok5w9RTGxs+W9JYURtdZ6Wm88p575yI1anS7/hZH
Q18xRB0PkupCwAbpPjl2GgCCWqaLgj6I5lZ5Ai4C4bEDfvvnP943m4IIj968ir+t
XxCWASWMHeF6wQePV0Pyrc0d66viNP72YYaFffHGXJUigIHhKd3HGuYFiyi17tgw
tzPzkB6XcItmZzpWTkLnXOWucNx7Xr0o4b1KTTBzjE1HMIYz2XR1xZIsfBcoMtaV
f+sm8OfBakhzG64/o8gcnGS5dAIzqsu6Y+1arnb5n+BabsaL0VOWZT+kC/Heqe10
Lx9+b/KUsfYi9ZCxH86tIxbcEBFdBqS8ZIBZiuM05JiGGOVZuenCbpwqZ1PiTTc9
nnV0mKR4UWZABbACFTY3CZdexwkG7lwfRcrGBHPmQvnzzv7CKZW0C7P+xvgBFIFl
sCf1CmR0SMGpwqwatpfNyAwTpQ0anNqJLUf2W4a2s4zaZOzqKpfTgTo6Vvs5Ch5x
TeX/tKcAZL/9sVYnzkxY7fZG0djqwKSSw1IKnjWehv77SGmlzxBcAzQHsEBVUlco
AK9bsh5Mmd/UvRblmBca/Sr/NVHWdDK/C6/qRfwi8VQZrWN0vwVnj0GIQ1Wc2/Ri
kzErbu2uFKWFPlJrI9EmE+du1UQu+ba5OYJMa6OH1lmYCvk2Lg7SvzofTmPMQ63/
o5gnq2PkuFdM/DJrA0CKTGmjtB7mD24Cbd6y7SElMaR0akTsfW9fHNB/sBeht+4n
VVrWe1A/y11ZOgkK4/yUUbIqWEIULnUt4sMD0hZOI9Mghe1+g9Ier1mMrFJaUg8l
1NMeFK6JTtCDA0iJ+QP/+2N56jpW2J797CTnazNHwcumeR+Ta2K0gtPTOx+JEAGa
cOWnxSsk/gavILow2+O8jscAFdNX7D2eR+t0O8ftBJSpftmeHpyEFWDz2nFBcFSg
rxQae/yCIE3Ae3lEi95pZyyLf7fQf2vmGjI1TucF51BKwwHOo/4lG7OFBglBIiKH
xUsgHBIMQ1nDxs/xNAfZ/QzloMC5Np71eWlHXOt+fSz0pLpfkiOahoEyJQlh1ITc
QHhIEH7mawPm20dHlHYfrYYAcgc4CF/3qBLB9y5YTduHFumBHoRhmxEDQuIy2YHX
HmI3KLDCtZOVZiBbs5PZwJ6ZbFZz2RzZE3YbQXZGaTOtGit2NLgL93wr7Bee4xR7
O+0O9dH4H77FtDPb6UkXK6+WBJJqoTU4TQ7tPPThZgBC/uThIXsFu73VWvcpiS6v
nV3Ojutixk4rr4GvzrkB1onJCwd0KfkuOXkR8clJLx0ymaOyuVgNippgT82Unh4B
4zGTf41BJPxMUVVJZRgWCgAcsqAupSGn04aUrkePPcQgPLadp3kSYdqGtBADV+q1
nfH3vYQD/oC2kUBSVL9d/Meoj4VvIQpDof9aRHnJxOX/hvdzyHTF5bsLNqhPfNtv
uGoqMS3diq25gQDD0aQI77J6eLFTuwUbDcvnh7mGmbIy6bX9MV3yeNQIikh0ibfP
NUyBS6fr39bnEzgx0HdyUkqizTfSsRWiGm7Ok8MNPtYccX/nby3ykQqndJSRIPQh
2Bp87qNqx8PVJRa12bIQXcVUyiiqQxGUmkYJz8D4v+mjMNMJC1QyQuC8FavNvFAn
07vYlneGd0yFzjg/wklEimIexhc9PtB7yNWaIMA/QWxSn99pIiGCpXn6oCswHxZQ
iAJIpvQhCI0P3+CO2D9PvfWXhFU9ai8SwOWqouOeVM9hksj//QqBJNtiOrHpfI6G
JAvacuYCjd4zlQIqBAKDFTcwkqQZtNnJ8JBNDTRGTssEIKhIINYoRFZd0T6GYjTA
OiYctNSsf5gHzDTfmrTQ/3A3djnvL1qyLUSq6LGk3JlnmJMR6orWqj+NKygIBiBl
2Va+qfDETgPYApPQ0Edjm+fHbJwRMuHFS5DRweaL9uh7AwwIWR142GKyHZq4m5/O
V6fcAf2ELAMaeq6wcn0K2/kUxbvv8nGpxk5dkcBkuqAKsKV3TbTLej/l64bmHPjT
CmGspSH6ze6G4FpjExNJTBjNoe9QgKxYJPJIU0Y83Aid6ygeGDGk2oKLNJixwbKq
NOrDw7IymouGE8vLtcX9/si6KhMAYmlAj7qMRBvx3JqM5gl3czrG5rAQspFmsCJf
2Er5artvOatoHFRWEm4DkJB2fUFtWEznkD+PEyo99JR6rUeyjSpq7m5WPSZh73M0
Yd8AYBnsEyb7EYmBBr32Ge4hmcXWy84u+XhZImClbGDuaXG97pggIUzYDQmf3t+s
oF52PFlDNkIHHBnBINL7DdWgGUSzIdC13xKyq10HLLkDbqq3RTS2X61UaREgIPsw
lpoCRxu4brMj3A1lKtb6IL9bBri5mUXu4LH9AXdbZ8Qn/kae6+5qvbdUvtV97GCN
maB8yjW1TFJ1yfMY8YYxON5WfmzxDnUl5teLr2xRMSCkedoQ5RpSG4J3e8ZNETIg
jbpf5Ts3Gj4kl6hXCdHc63rFwUfBxWfnRppqcn3CGvXpG4UXlWCKW6ILaW7ru09V
imbrPI/ibDXq2Hcc8FuBwFmqmR9Zq26s3jSiiMdLJMzMXOjnZBrC+Wvvev8E1Zyd
ll4fI1MwspUZGy9aGOriUeX8ec6ST8FtgvJc3wLESwMcdv1ZLOLEC1WzwYvDZmES
2UGUuru2+rkVjjVEg46MWH4Nzjh0S1ifsXU7K1jEEETU4FSLrJiV/DRIACSYEIIn
rI+0U6WeSnFlCfaWxC4q2aqPIGV4o5lfcsKBWFyHrsVfFgSt7Qg0nJekEUKMNF9+
I/57E0XWe99pMcYPwURzQaKqAOhzQvMLoQRlHxmIib9GIJ6tHnGnCGnuae+cVShN
l3rVxYvgTEjgOmw/WCdWU/pZws4PfPUQ6BrdZmNWiLaOD6VxwzEc7uIyg7F1P0M0
xyd13XC/k55wRp/OjQi/epvfn9LgKg1PqrRn+BskjCPgZHDcAi4XNUYXtPk8pof2
gKuZjdEhG8Bq1lJRI2V1YwRHMuWyhnIE5wL0usQHQ9ZIMda24bkAgou/6brplMSv
CjiAk2whlPSF7IoD2Ibl6BAnUKQEPMbeEFGX9LFXewJYWhm65ifqHSrhUaZaILia
5nQRiV+H8J02iAlbzMriLnqp2YcngHNlOtroTuPyQWkXDP98hZB3xBLJP0m+c8S2
RxmLspByGzZIKGb99afj5hpmv+sMHszO1guMzgA9bgOiNJVSBDdeYFmc3F1TLV1c
Rl6LlEojlD77u8wEVN6qy0YMAGQg1cFNaQevfxhiChcIlLZ29Bf6bKfVtaktFvTe
8BuX0Ln6XRNlwCatY88/MOTMv0GsAkB/3h9JkLR6L47d+SUjWTeFvFZuMHKQO5dL
+s9IHnJ7Ncqo40xlM8LFdBy7iLfs9GHnMFkKD19Bo4tIrX+Two9JxdfhAn4/cp3V
vAYrAFTUh8vDeFngMzS8cLpUSVs1xdbVhHBSS02VPrhRmPtaQBsPqe748kNgXFNN
GirPwunQ9BZnCBd1zIL5kYwoFvcYE1dxvN3w4opIDdkIlU3iI6l+775FeuBY1NyC
dA3KBmwv+9HsWXfdd70RGsXmTk1B2dfW+dF8m08DNmzDlRm/W95dLAj4xSd4IOII
79Vl6/SGIxsp++8ikERzzofQ7r9V8zEJOTuQb03EjnLzu/Yv5ZEW5RVdS7VQAEkJ
pgucAgPosKL1iiKvb5wvhJE/JzxIm+tkSi/O/K7cAFmMC8ibsWPRl2WeXupOjbM6
PSm7wL/SOGuq9bjDSJS1mWO/DImmj638ILRbUBC4HOS+GjTnTd67Afory/jT3ZS8
Rx0lNVdyVf7MXLaOj1YgfLouFegTC3qyetGuNlEnmw7REdoLaQP/vKJ+4N+u9OeO
mgKUn+5GtSAq92STt+UH5cAQxDHkak1YEFJVfWxBcgf335/xGqrMDyJ31pJ/KrW2
ROeQdjNIB4cm5KUBcmfPdis7eYtOHP7DwKHIH05Hh8YrcenZdyg3RtgOTw79o5fw
v1CGPN5qcyqWegv1pfBlzGGVWBBOOagThGshIC4GqEY5GEgYLYPCa+HSd8DDFTX1
4uRZybwxDBz6nbKq5bkAHs/tqXI1Rzwc4j4qTlvLKvjXS76eJqYZP3vZnym+tWBZ
nRCCnklRz67D+NyHsilg73yi5vAccE2yxIEIk7ydb02GdvVwr3DXqfNymUXq/1pv
z0qybSD8Km4LJZZwSF/letHnMAczpbHO/91c+RheZHGr4essunrTZqEB9a1QYXay
FE+KsDkTl9Dj1zRLpxpRL8bQIxisv5LRhseTo3EyywKHKIGwPQQWLgQ5yInAWgVb
x0lVUjQBo9YP1HhNR/T7zPJZuNeMzrizZJiGXXGqbL+GHxrUGdHqOy80QP/XN+AK
8nOfvklKkWNv2V2oCcYZJTRIbkQyKwDDnZhk9Wv4/a0aK6BynOwj7lM7cUGUmdzO
gLV3OO17iXvWncymUzHDRpI7fmml1RwYc2AQgjdO44ZkxZybZGTZZ5oSxRfH9vN2
9VDhievj48FZdFVE2QkdMilQxsEd5yGbw+H6lPn5OYV57G+vrBTBFvE1hJn57Kaq
ipLPNXwjLAUIkKgWnEPHUM+/YMFrxPf7YiR5FEtc6EGEWutxjySVZOdU0eW3xBei
kipaY6zEBngbbTD7Si4Cb3gk+XeNh86WqKxd7jjw2U4x/7xkk/2N6HqucUMJZC6c
QOTXRlIhCDkfBxKWFh0XLZMV7Niqzk1wN0qf5ZkOx40zbxKNY+jj6N+25Jz3EDnm
T4Y0G0JDJZhj2hboFwHf8BI7vpl7sd+CHafBxW4y9SshByetUuQRzFrs6VakmPYU
WnA4M41AuWpd8TZXJhoof5qc+rycpY+q94ikzeJRNn7dlMWWY1AWHy8U00snEXwX
qvzWdvS3izXU3/hTGjlzGH51ovYZue0/YG/bpYJMHYnColcOyoeGY2/eQiQalA2r
yMaYqEJVq6KN4yN9a1hFI+DlHUH5oCvKe4pJpYp/1VemA9RYSwDBDp0kKw/Q3A2f
EZR/OrOJPUfd3ZqqN7v25K8fe2OUKdwMyD3e3E5tpX/YwA6WLlXfvGURI8SrOaik
KaQuXqgsd7dAJhHdAkn+3/rVPY+yfOHXsYgNR0pis0EGAFU78v4RfFwPWb0yfHVS
vlJuDmCProqdF/7+vYzIfIn6eKeJvRte7t8sxnBsbt3dzoe8LKpfjsoUTAqb9Pxf
yMor6BjjhvNI36FRCdiYDki/1y3zcs1RkA79KwnziPPvzI2Jkx+Z8yObuWeQVYIV
wJD2+d0KR6mThM3rEGBUwa/JUq1L6eV86j21ImV+2bj8mCmX67xJJsjeFPKvqXir
Veks8O0WXsh+J7rJsXYEHbu+kdMyUkmA/vVjKAqy8leQYZSjoeyrCt/bU9WM7bC8
T6V/mYcMzYgqBzT+UjeI5acE4HNTFgavdworezWhHSnKwqaQnaxQcwevqILnihEp
miFmACRpsjdtKMbPXtIIRM2h7oMxNl7nQrEcaReYnGPXjS8lvLxH059whNcX0RlV
OqWziZ60Ew8lUAfB1MdV++BfadXbX1FFIYlvChYh++QqlsnogC4SklwV+VcUmT76
l4FJO9zyMNLa+zzsBVyYeMybX6RwKVfXTnLosgDMLuENjblN+6TigBohDLGXclVw
J2sEdtz1ASXbtjrb0RJkxkyKjUpotaB4QaEM0gTIpoXYsHUts+bJb9xkp0n07vAn
En6t2UwXZ8vKxzupkau5slHhE4FdRLzVvCdx9+nXmmuQ+N0qSKa0wKt6ekOhPLZ4
CWHw1FrGRcXIqf0dHGLfLaL2GUeBRyt0fNcwPauiQKTvGbQ9aOP8UjZajTpFGA7P
0ykEjbSvNO9bwTKu+YLhIyjes+v2xLGbhNcB/Fr4dE9g//NdZvl2J5aGWEEUkT1f
qstgaK243KhGt3LDA2qkp3U+rP/BsfohUxQUh4S1CGzvSNc/NCvT8cdOfOnJ27qn
QRqQJW5FtxAq3pJX4arSufjE06mXmXQ97gl/cfNhQu8QhyXdBPNwus/MOI+nnwDR
6sqMX6FQGwFZuBDajH64Rc+B7AQZqqB/S8f6/NdyH/fJb2w+HVlB02nkAujwK4ni
2QcZ5YDARAiNtsBpOADjrbsS7XWpcI0z50uPODNkiWzhYoRuh1CkMtXAi2rNaC6N
WCrohrtGzBk+Sj24QgUo9QnMirOwLjAGqgHJl5RnyNp99yXLBMecc6Bx0Q1eRd5y
LviaVnRK5L759k+7LRmozYWXdOOcxq6gZFuN10b/aESqczmWE/q7Ej6eaJ7waJBp
O0Mly2KJe082nMUnIogbTtze/DTBDfkBaFrXJ9f7fLgTzYW+dBA+n9PId/IgLFnC
p1fRmgT0HhQywkUoq2cDaJfPG6BoCElKZX/0+MIlt8RKrLNJFl0AS6joI8CZ/dqw
4noCkZLE1AAB+AKm0OHI4odvzIf2YqY8LJTJrZ0/ujquznbBI/z+Cg52bDamA/tY
4x0UDe6vFeio4vY/TZ1hkrm848jjdWVyhDTPjbn6eTILMirPugchslOQDWpRkgaj
KVD+wxjSUTh870OgxvbnLiRaWrlelrDGwbf7myzVZTisAKVo1bNOPntXDKuDiF1a
YsAzgGEjtSGWVfvqe2v5TSyiIbxu9+O5LJkcUkMxgk/tEdIcE4fg0TklMPIAGp/H
yLCT5EeU056abM++eFC9nsPGXat746cvOvRQBsmyJJyLPNtHxovAH9YwifvvPWfs
PxuV+49/r4Z3gtVoZjKZdsCGczB+sxcfdn9d1iAFfaQ46EcCadcw5wdR+z0sIjHW
xDxr8iQtrwkZPncdSi2t06/o6buIGgzCsHai9hJzsdWRdqaQUUkjbT+GLQMIWZ/m
hFqXJSzD/GW2so1TpvxQdu8yBCKOvR7LkxhpUX00+y4XGybgpHd6mmHz6iYPkEYo
KgaY52HHO8Rx1DQom8I50xwwT74xO92e7CQCCClvkFk5OAKY0XJPY7j1C4Ngi8J+
KwQOqEDkupGKCJA5qTfy+MVVvgxS1vVyouY8GkD8VDzuN9zjjBf/gFra7FXAgzRt
N3oZ1I+Js72GF+lL/KYKfnAu3AYFaxaPG8EKJuERkA9Jm2m5p5Y7NyCfeAngMylA
FOM9Mn4Jja8lIlHYMUn1ML2d3ruon00XIYVBMY6tTJ7K5Nl8YfIj22UGJURjKba2
1Gm20MLZihQgmR6mSm7fvjStG9EyzqKmDT86HtiPxBexBZeWCS5tuaMfyCgeCbv0
FJ/3K+ChtUClQKqPG4KAjtzQVBXHd+5i8L+Ir/vK1NnBUKXeeqYRUOxYoImd60Bi
u5e992sP2YG0GzD6IpQSL7l6nmj2nlAM3AMVrVdNFoY0Eq4gzKYmq3raoZ6t/4av
plLG+1cnvkBUeRjZb1E4bI2I5mlThXxMVMEECPF/R0Wm9P9FvFT4Lod33G3MWn7D
gb32ii+HfiL2H5JPB7a9cgsIH/tDDeDIij69mFIxpNHayt+BdT58VeehGIp2KlIa
28+Hdpy30Cbf76hlJCFwV591L5GqBi2GHm19Yu4qN/eZFK4+DKwo6aX4LzqphaJs
AF2paU1WluIDxWX6NSLXeGuploCSD5eHBnTsb25NSpernbzHzpqt14DmgkdozFFy
9rEvhdQHCjatNPuBjkOP+pazxae+Gxoh9cwOse0836NdKoij4lqOXVl/RkVjpaGE
wHxIbYjUYzwVlmuR/oZbHC1pcXem/TUdKYRHv+jPojUsyj7R2zpcIoyQ07WMnIEt
8m7/cqof1JTosFpiJ/eRLjNabgiesw2w3hWgY45zZSffcxfxU7ps8HfdEteV+8XF
Dj0hYBW2LJ8uEHHG9iXedmDtGP9vr8vj+u+RBNkhgVjiBLHrafsGn20CBKv3LHDi
4+PvFpmoZibQxxXTbmiTvhl7RlNT5stZuuLYl/Q8KvLRKslz/nJcp0/hmDoAnu2c
ShhVRqB4FPgOrlUoKumeFDmtvAcs23YAaMKoYwr0xTiNq9Z6YDQWOF2o3l1zKg+u
b9vXr3cn02NSKWLugeLDnSOKhQL9tMiJMcus70Pb9UOJKWfhRdvq/BTZXuII8td6
2hC7HRXl6YVsBh2RA3qhojl2uO48F7Y2z//9hArZZ9BvucPdwRaT1ruVmcDkFr2R
UqtH3iyCqHBcgcnmgfTfF6tq9GU7TuAnBE9i06u3m3hwWEYP0aW+ZmyxAInF70yC
h7SzQNx68pQYxvp9ulYB18O5rETjVp/QdPgZn31leEVnOBIjKxtPt9WwrNDCsnxS
cUrPVW3+QdRcfugKUGZN6YfXHvivSBRDweJWeLNOFx3czSrYd4lWv+WNPjMMzD/t
O8CEq4j4WlncG/TtzLFXRsSwGA+s5Lx+LMppU9rjkAtQ4mgKKH/Elo3W10Acofr1
EbPKwKKW9PPzpYHmz4dVlZLzxtnzTd9htohMUnkoTTBSt/PVvglaJd6pcYAXm1rY
Cj0siki2d5pUqsF0qqxYCUafOXhF45X1jHCm9SY55kHGqfEKpKdOGxdVpCbeADI7
bW3NebOflQlDqs5QDd/FRDV20GSpzPLC7wJVNU0Uoz1KBgPjGNsKKE2+lrxWnMYT
jfKY5uHZmM7idx/BIE7glxoeJAsKATd5ghMxJ/EV5ZxMRFW4Zid52g6y5y2jTeAR
lb32OVaPCT3CZmvsxxV3k6fkdz4h86Jkg3F+1Nuj3RlefQ2SUIx86kch6tqUnMHR
VUYyI1jkaT7FFEVnqPfYb3FtUdMjhhwdvlma55QrWz3ZQ6QBELtvT35oHmhoVIkS
WPVhLdpJgVnnEugFhnknezBQJwJ+6oQKEuyY/xchQZAlRrgFVIgAforFmt01W+H2
yRCCVDHefmDJKWGpKhLsUYla0dH0KRtZh9IbP9nSWuo7VNPrOMSo2hKq7NNx/o1d
12JIWYxPmHob0pyhgHY+N72bSg69mFrxWw9mFeXf/ME3+EIXUcJG31h6erY4NBAq
58V3Yg93ObmN+K50B2GsItfEjJUJa+XrSNkhqjHMwxLGO5RIX27VfxlZ/Rmo9/hG
VOmpk4OjiPebacJ67oduUwd3kYN5R7voGOaNO53YtsiFMRhNDhJgIGC4Eic8/lez
a6BmHtxJp1j2wuKEUMODAhxoLDNFwi6xj7UBRJyxlSOh94+I6y3I50x9ASL5cgxo
ERc9uUmV2tbrkY7JGQpk9De2pa6S6xHjfwuWKLKmvVoEJ5bAd4vGgCs29hc5JaPN
TkBwIa+4mOEGCvduWOt9D2/CSOxnA140cz5+VlT6FlUQfzBdjteV+lU19EJHR2JL
8EQeQh7LM1SBY55TJnwuYEmigf5eEzkAAyofh8020JG0FBVGCv0G5hG0NOuAj4Fh
m1XECiNbfj+xzpAvb0ce8QFgHODOnxGNT/pDdrF7+w1C3IvVAwg/FOIp5p/qmbd4
P4LW8Jvr5L+ocPRs0JswC7rDa2RjSTEJlBIAMiUEqNNAHM0xObe/qyDwvQ88RTrW
jHUMYBO17sOLGhlT3ZG92VMds4TbflA2gxdwMNwsgmoSmsD9hqQ8vg+59ObgBdR4
mlk3MBb170OaeGEpqPymiSMogstI+hGJe8KP6fpAUwZ6ebf5UPmwzDFb6EeUVY9D
yo8aCicfiazvymzIVkVmeN9jUIIa370aah94MipCc2QDEc43WD+n+eBltIvvkt1G
DN4GkDzrKxiaM0Gi8h0lP+AKZ8d35WFapPp6joohqsRnbORqOykThy9U+5bHumzw
fGwuPONnxAnKbQIF/FCF0GYRPVlJh2QsAbNHU1va0RvcQxujNI0a6iCVKO0NIlEN
DVlgCQku35KIykdc2IZ0w1gzaF8DcX7sd65RSpAG2Grpij1bknCLmjVs2aRGkPaT
0jPd0u8yENs1wmidhUmSUkj0eQHq42W1aSOa05EqJKalRIAmkkjWzpTOeXZOMvac
IaU39KS1tfXgjqLxD6GLOIDrYb9kVZnemtXtKR9DgJIR1e6s5x6M3aCe3YDRJh6C
NMFPBD90GJstY0aZKVlf3uDmZmE+mJaNjtrkxvdIpHWiJzmazlXYavGlffr8IFwi
Raz0U6T9/Q+ffVGA/TqAUgpsuderaamPkaWlaoIup6TFAzSXy5AA5PbgZfD8+rgy
1BjIqc182agNgxH9ekn/Ah2dM9VnRKmN5Dns5Y7hpf4s8d96oX51kaM+IcvGw/WV
DWgkwDJId1cT3UmM8OkVKUppcs/PYAI9GNGDn5J/Ps9U2EA/KouDVviTB0EYO9ff
1jijStxmnWQu7zvmcOKiLMJFcLr05eL/6VV8aaEZgjUw2qO2KWm6lLx8TwgsgmBp
g7G7tPMfk+c9661HyDSB6yXEbthegvGG6dDXYBoiiO+6f6Wvz66q2xC/cXcDcwRB
GJJezg7Gx84VIUpJyiQGkAuUIZWPuElcdGu2G2tyWl001DQ/A6P6X15jOt69ydEu
qj9hI0P9l2wWAvOs2GfNvJc1Md+1hCLgfHlbo9HAbOst1kZ/vhu5Ak6VZCaXLv+C
VKjo1EDYK/o+hyuYd9KLv5dlUg09IqeHKLhltS+DE6+wZ89Pi0PRG97C5H+TSOn1
+d4nhfu/05DrakBcJ3ttLo3/4VfL72qG1ckZ05tFQT9TwJlsYQE/YdXsK+VFAQb0
spWkAVC51Nt4DO+YynrO8g9lEaRqqBmWRqyyHQCGOr4+YCWAzNgJ8194xiYqiVWi
g4ms6Oe2ZEAvGjeXd9sJGEwUwUs6tKQv62Cu5hw7zy/dxAPfTj6Rk3HFjy48SPgR
JcAbJlQzGoUG12Iora/hGAR/9YQWDKkkbTgEZH46ChgcTivmlxL1tX9KmPXrjed2
TDeDC/EvIVJSrh6E2Fz+kcIfj00mXWbUiIdTsNiggH+0zYsFJzpx8Nmlqq0L/LM6
61HgAnnhMN//DD4P2SYfqI/WTLh6QFfxqkkrkwqWzjkAfrUFhmB1LB5fngjO220E
nj2tlWqMR86VXQS0QWeYnrNs0dU8fVz6XgYJCbGcT/4y+xTlvXe33nSdDDKtBgSQ
GH4RId+COFWg01y4uBBVWrafPX7GxnQ6YGvb6ekhmwQ+fq5nZkyHewsTxhyl3hzE
9/AjzY3dWa9hEzqxVF2fDsTs6lfay2ca9aKZpr9oumgGBNnv+/CPk/eLx5Jt9SaD
NdVY+LTe0dwr5uE1kYrBKL6JfgIUlPCSH4mJZoTadrvwr1TmqHJgcBlYnLU15ES5
bjxTrei1UZ7A1Kcx4UhOa9YSwOG8W4IZOfsg7LBF61Mb7DXujlleOS3hUbNrSN9j
Bo1YlYDbbBIXHaCXUlAxXGg1+kNXYj0UHesaUfQJDYFPvfWlpHTUMO0Fgft6Q+jX
D0c2+uhx7F3QUd/g8QXdX+jhYJqQM4lGO/0Nl2BOZO4lmXHzRxPIW4X1+QZsedTc
CVSapQT5g7GZYuQYs3sKh57SgCRq3GZqr+upxNprny3VrFJVPmGMwtT8sKJ1VmZb
n8xODZyJFYhd6tTEZ4mE9KkOBGPlbKMzWMYUB7hHYcGmRIuI8QAN7nKaYf/ATs32
Pj7w6/jE7MfunNo8Xh5YoTwVp1wW6bjUZCq/SRu08MXbX7zgx/vDW4tcRrPKjd0k
y8k35nSASsQFOEVavR0rSRm/sXUu+5aFEl4nlvdR8wckIlXChFqYUIEMcjZETY2Y
wvkbjfRcz1BG8hIOGqEFix0tnlmV90ptH4wsOxXCwtPqgbfBoixurmp9tEsvKn+w
RT4hIfxibB9i5Rk7PA1OCvqxCR1QPUcwjPkbCwh8+5u5nFdNQJIYVTfWdEHJHdtJ
r2sAFWeCmzOOVNOwF9BTGzayW25iCAfK+2J1OGtrclYvVgNbZie0q4Vi88dNur4y
oP/pXNk8YnKSx026Shs+++wxlFhxmu67+jk1B8vj7p/OHEneG095lA/7PzJZHYMl
PtFzsVkCpWgsyPwCNEAoAEQf9Y21R2SfKD1AjDKvUGYLZgFRZ+Y/a52xVLY0bWHw
UcFHpH5KEzb8CXKvKEqT8eY7WMf0X4SAhrcDV1JFn35vNJum6wo+VfXir38JLsat
mdxi2ETnn56x1g0PRNNqytuUVH8/Rm0MYCRxLLkS3x8BPs75ah1hkOKDaG6whmtA
NIkLoKk0s67SBd/2Be4ScJdIjMs/nHpQ3jl4sAl6+0cQD0P9WvQCNkjyRo8Fsngl
S8DNzsP724dp3Evlq71dVRsoxOmV2kVm9a8vNjr02vvUwrHudifvBUkbP7f/2GZR
dyBRHx9I6etIDxVuMtngmZsKRYyOodEooJAw3mFy2b8NijykyIkS1YTxfrE46O8E
qjcDK8JOAghIVqWMCQXq/8llr1nj9sW+z0hcaNHTKUTD8iYKeP3/uknD6M+DZQJf
efUxz0XClq8nA1OeeJ/phRs/633zDQpn/mtpDqarCxjjf1dPf/d/qBLgTt0nUBuF
xNX7zL4vSNliw73QgDBbbbi/d1k87TLB1OXojJH/QbmyCfW68HyPUtAWR23u76/x
GShNgg7c5Kw9SwfFsX9FIyB1tAhQrZtTau1aJPu7d7aW8qDgZUVXkvJkNpUoNUUs
pXxrOWzo09TxjeNTXro64Epwqfn4Pe2vOpM4C2XPNYmJ2gd7q+EujZr7vXgy3Md0
eft2QSjwoLaZoXjPbYgcLibgMaN5ZJce9idbKGVXv3/jkSXLitxPDaRl9RwB1lvo
0B8trCczcg3DqiHhQ2nmZV1GFjwdhjRqzfCw3kVJutC+gerVXc38wNsxNz7Y2lOq
jP8lbfKy5h4OpWmnQiGITodcPPmFGIaFqUVf0b/4OMY2Gfioxdy/zTfIK8/S1PyD
A/8RskROQiprekXc2OZq1Rx4H6A0bHehC9aqN5XbEoDMm/Pf97BIkb0OFbRaye4y
f2A34w0eSno0+NYDPFYu3AxcE65B6zMBjOThxzKUxL6qVwd1gGnpjux5gKJ69HTV
EyV7nIauNr9V+QcvuQ3RvvpQjE50t53XGMFwIG+cqY03cgHa6gOV96oXMPZtYd1H
ohDw9cchgMEwZm3+225EN8RcOCHUbYJoIeNTyS10eHrD7wMZWlC6w72QquYEYatl
Jly2+YbYHEtmBtMw3cz+kJsAO9+BvR/nuX8ifkXTJ1FW7h76vs7EaLDxnEpJk7T2
mhP4/u707hBzj0pLVfWxnatlCm910nX7tYmpN4SyU8cKBfg0BPyY/sreT4zvq0MV
aseLxoU1AyT6MZWXgXuXZy05gWDtBpvZfkFUESm5Vqyt2o5gohKMVuVnQJqpZk1T
+dSAbL1D/wmTPHkwvMOq7J5aWkvgr3eatL6Y62/7QAHluMxB6KxSrcJloiofor4L
aV3dMWn26Pvwz+GIuF3SM/0/IbU8ee6myDskoVbZTiYNkVKNvJ4SL11MJHf/qBjx
jjLhZQ6KgcH7U3UaN/R4AzDKi2cSLmBqoQdBctdoR+i2zHPuswL16K3NIKYyC4m0
4t2dTK/Wvu4SC8mf8rFxOzsajqiBWrz9r5Bp3tjQ3OqVc1p2fB3w4/lLoTKIZcZT
x7K6vTAT/KcX+1QqQHlJDrCAHHKkqL/1AZlYLKJ3eAmVqjNO6zSf5HLIr3FzmAO3
nPEYmAUxm9TPPuYkdw2a/ULPYj7VEZ1j+01deuTgHqHqP680y/RqD5R2L9CzTdLm
JnmlxZUeyI0//FwU6FVIfnympvYqZEGeUpAfFc4Uh42uaudeh2o2q9ejxvvITlNA
fFIQaTFC0vEjt4CDwANSNqGf0NUjNb2gHCg3NlDX/RUbg0CL2qoXSa0FD7wzg6zs
2qN8nMX41wMfO3aKZZu0D0R0rPPTPoFauDBJWXiLihD/BtEy4zy93hQKH7u1Gsyu
teH3Srs/3Fm07/rcd7qC+AwhOsERazGCyao9F25mjwDEsmyjXyBVwJ+vEqlSJ8mS
00i5KSIBKBUW7rc6DPFqEEQTLNnufvGZk5c9X+m8NkWhU7HWV/er9yOX4yJ8CYGx
Bfkj0WSgLIaAzFXOiSr9icxx1IcSxJfoHbl+CpnzRngIOhr+qAFcRkuO/KjlWemh
QahEJTWxZELeEMPIUos6Z5pdGatU0qk1PnrPejyOfvbLGqZmEZb2UBfvZd/yVlsC
uo8wkuq+976F/ZJc5WoCKycaSvyT0FNmtftxnxqYh5/AYX7scUXl7UoIgoz2ivy4
+3XYPY/JGJCAsByapXzbAgNbAK8Z5S3jbemMhNZeVeBW8XbgwuRiY91fWhbf1Dma
I87SYIwk2Ovp260w+j9OOB/zJyG8hbbDEHAzipcLuBtY26taBRgEZ8WQk4Kgd7ha
tiy/lmmV2EyezRXxrZDE4xN7HtZeZRUkAnDKIYVqJQ11wT/fglCtg/laltg6zM2P
2Z1crLdGlThez5cX/kB5xrNna/aHA0QgPEVUI69HRn8PYTcpIsYPQlChg5Fvr+HU
UvbOdxlotBLzMgv45O2gm9sfO7+O6hDk23kRVYOSgCvQJddjUN4GPreApVcPoGDL
BRGYrHkq4WjgBM1EI0N6Vbhmksi4ZbXzTBhyUztRNSSt1pdQxS8o4IzBiORkAPmt
sjNEhBvPCb1aJ+CM2cqyCi0V7p7PuxCNvyvExXvfW6t2dBgA8oo+/iCSHE/2lly1
uyqy9HJyQkW1JGG5rxf58aB/GfKcMrc9a4a/Z8hk6KcICzvxwSpG/I7RumNnY94z
UnsWxrh/XPDqKduxM3GW0nT96DfPt4s9jOaPiVr42FglQ+XLAWKn2M2LpmS1wfQA
tNoSjXkO+u7h5DQJkA7m6qve9a3D8F+7GM4WNfKLVskWe5kieAXTnsp/HlHO6MbZ
g+rIZ4SVoNFmII4kE9qwvwk8knLSN8znC6fvFLUGVVk83XhMquQAtICo3neayVQH
JeQA7h5oJ+Vr9KoUyaFNV7sTGueqO2Jd24iC2UwyiozQ5qSNQYmArcu+j1KoBjE0
C5768Q7CmSO8DTewizYOsCdd0R9o7gO7DfOXwlsr9v1unTCsObxavL+mYVRsbxk0
0g6I4L95FhV3cc1ZtakIWEB0eEC65XTmw+Ln6/7iWISiIzaQ4fVopaTb4P4A3FEo
temQAGuCR0m6bdcBL3Cb0g6Fi8zfL6GbOKbb4S/agPdfrZTpYw9o8XHCdaHo3qdB
AeqKelttuQSqLtdC095x7bKHLMZQhc4SQBX9OyQV6oF9QLJweRMUXjswTGaCEMMs
tdTXeSli6LIdYdlmPdI9LIz+cxGoDc0aLeUVcJhUVrEs0qK8s438GfiNzw4UbxOW
fTV18NzQIATebQlgFh9/UyRVFl+w9j38kjTnSsNPgE9Hv9GQjFZL8ilh/B7D6KB7
ehM5sKTiGc3rggWmNb9jUBKgsX/RB0/tpaM7KG9EuHN6iTsvkY04nheNoTdSch7D
d9JP4Bfm3kVBUSDuKioT/BP7N6JLebQSUAz4IE8ORk5uHvqSe/lbrQL5xfRhtkJq
zjqQeD4YIe7WY4XbO6fp3oXIjg8hFvlZzgtvuzJUMlBi35VHrf0lxqSb6PSaC28U
B3RBnXsf/32B+/op2odS25TlCb4xvhwx3qUnNqtph3iQ+I3hImRctEEP3zdQCIIL
1TELfp9hZZFKfzk0cmRjMv2Mmvj7h0OuqtiFVGA7OjxrhdpeqK+nxScdTiWBLu+n
9gvGIbj0XtWnsYN/8AeMtyPX0n5n1biMSYSBoGOc0Fh+NwFy0blXksvvn5yMiZ6h
lqR/WM9Yn9vNVQa0IaAZ2/T5fQUQCFoJbfHnXH5V+a/x9/7bTLboGPmikgaddfvf
eiP/cvTTtGFenPFjJ/Fy/7DSPG3PcyKvLXQRKl3bf1/m2F+obl9KSRwi6+eCXbAq
2/S453m6HFvIeKrfHYL24lt7lYq2McBpVuGRKJS/h9LK4vawG59ted9rJtbc+U7N
4tD+kCEEHp55G3xTcsJ+dp5h7YvTOA0mh+jtA9/To5tazaOGUL/Aq7EnooPkrGQR
oekrfz+q1/68hwa54T3eSNypYRhZ2K2w7XbQbyPsyO2gqKqvwqw24EouEnEEMunh
Zf8t5Y8qi6XDt3F+sLCipIoFqLgYLBtwPt9SJUPD6u6l9iU6PQfk/kcSdEm/3/8O
TbdpngQpqwV0m9DBlXa0JMeoLgvUlVJf9UW9Dq+mhW0c12Pmeig6KTf321nIb/uX
UkmsBeGHIKnyr8PygkX+9UPAKrjLYg/s6+TKgHnJr8s2+qXo42iyMue67HnFNMNj
5ScOZAjcW0eSK14TeSNmeyzuXOtvh9w9XEM7V2csHXA7wDJ9FEisQA5Luzw+0hEI
WGt2gN3TvCOQcfjE0qzt/j2J9PDN/lhFn1urnQW5SxrgZUv7grexPY9MorGb6/H+
0TLUZAwSp3SXsS3tQTfTzQ+BNiZnFcgPWydxAZaNWOWu90dvwNBDGAXkJIVBw6Nq
OMswEBh9QWvktyJOeb1ysAkbJnzH8H4un5QwzXWRpbQbNR0ZVYoYhSPF1Ay6hJBI
UcbWss5C3FSqD0kzV85ZBQ9l0Yj/AIMJR34I4byjhtQnWjY5QkkuJY4UtdzhIxmC
+UQUTInW7bhp4HNSgdq4kuW2/awgriu7dOnyOpbuDY1/24bvSHslm0AYdMOhSqKK
rV/gMvJmDynMb8f9tGtIXFlRRz9oxin89e30NswLJNxpxl2u6jySPjewj2MjuQ/E
CbqEdO7TUaBHlOvtHuEsyLzHcPy7+eG+4FhzpeORB1r33rSIk01N9LzRsQYCVB9P
W/EeHURIqdlEWgCfQs/LDzME0b/w68kFcjCwT+UwKK+qDGQQ+Jj9qFE2nv2JdAkB
s7kiTHJMPmzXYJe5XfQd+ub4OO0Olv/OZc24VITcDsb2smxtmInUDinqPgT8FZ/L
3kO74FTjOXVsQjtMxg4W4QfS2LcrHw0uZ84NE5lEHjwCK6zMk51Cas5jsIPwf0TJ
eAN0I6ZVQoYBFYsat/jaDnlEd+1V8SSAvVrxB0tAcMwxI4Q8CEu+MalQKv2P/rnQ
kQvQZq9F0NMmR9oq8P+iQbeCQEBfefN5rU45r3HglfQnr6shn3yOts06J/hI6cro
TiRqX/rO1HsYSIHA1Ja17PumDysEpelkeWrAox72rIYtlGt+TFneJWZxdtq9TXh2
LWjTDWlZZIgF0Fi7VnyV7uawBaDeqN8OtmPnVNTn39drX8glOuIqFiioud7TT94W
vY4n6a/C2Dy5hxf526A7Vb0zgem8NvlGmQjmOraSxm5Ka7A0Tmq4N9+3/EDB/jXw
VS6VJizdSARiheimXtxWtnqgwhu83O7Oc6oL5TTqA0sQ8R4S7OD8IELQW8kG+KFa
gqQyjE7Fp4P4V2D9AWMS5vzfk/YsN7k6rfxQRDIANKtuO6NAtufaWnCvTokAOCwt
AveMb0lh1GFcm+pemAahyg1j/GuxU5kwYJYwhxF+SGIyJhy45Td6fTh7hKg4rinj
3mGwtENTUUHicwlYTVz4nlv+zm8P3zRbnk2zoNNc/Iy/u+bGK4O6LtSWr9m2ojWL
/xWS9s05KDazU0Apfe+4MzlTtOddanBBHLLb+lZNa4eqbOKGQ150nOXdCI8rLx5K
WtC26rcHsYBvDqoFc7ZYXM/f9B8w4HPEb4B3tUVQ6rBxPiRTzBSMe+mI8Dr63GdE
FpbpCuM1Wz3cluGQxciFDOQXbwGK4R1nJM67Q0CC4vkiJSCub2aM+HDA4h/9V7Og
BJND7SaSCcPhxHVgXJfYBVZGWzia/2ROD1+VaClWyowWl697KefgGAxSxWoBv3Ow
8SHM75yZptb/IpUYSm5fKw6Dq4Ur+drXtIgOUK20NAPK/uF2REjaxNoSgl2hJKMI
AFDVN29DlkJNXBUWGCzCXOsPOmRszhX3DkfDNP90zWndWUuJJbPDDWn1pM1mHJCl
YjjZED4YKdfLUssXzZIPJ1K55zJmXCjtjoU88f0+2dThGxdOHG6Ow7VfrThEtGO0
EM7NLp5c/ON+oUMiZgEmCGxFkUnJZosFnlj/ylfSJi8Bbhe4GTs5v2rxgtT4P13i
RCo7Q7sDkiztkwvagV3EZ+p+Uc9Q/OjNxHIHXpgY750msOpqPpkVExL+ozbRumWO
w8GtWr7e0/DUACnIcHVX+Os0UJKxCciYbl5c73mox6Pvu6W+J+JAp8b4OLjWf3Bg
TavX8yprh28uEAs8t9p3tryi0azYv8YEtbclnHroGAJDxgTNZ/0lN23xvHbYDUQ1
YpO2YjVVGST2TSGuH30+4Wq1OWCey5klq+IyeVfygV2UAFW+inMjPCwwLF5KyxIR
4aNWtPCaMbN9i80bxUp2Fh1tQj+sfG924WOzoprLGCyrq56Wp9zI+mlbszAl9kwx
EQ/CdSdNip5v2vJwcXJUkf8S/umGWwzOjjNeidISlwVntpP2VaRxsIf29QK27rEw
gp2MPhEDJY/rV3UUL7ZHk0gshNBRvg9I6CylyHPou6SWRBXW6q0ojHu10XB3NYxR
c+udadtmqFy8KuQiUrcD+e2AGyV20jOmi5kG8guKc16uL3LOvIRZbuXc1FRJafvu
NHDwXYGIUGpRo/LCE0MItkiv1JwWXKhqoayfla4TdYfb6jMatKnWm7dAyawckNsj
Vky1lkgCyjBQOGBoqbiwg5RWAxtPy4NGXgGjuWSkZMWuyK9WBDLOn3fNO4KFDNtb
MDP29KmV3PhhnHH/CIBTdClZPqV50J19quGDVeFI5t/oD+lz7nIkJTYC/x9IOcDP
IxgtqVbCDs5cQ6tpu5ZuVRT4M3EGcVWXnN4gFd/S4OACpl0qmfGrE+5rRfczel2V
QeLReEzSnrtfOaZ1i37lkjORnSYsfhelNj2lMpSK5aTWtUauBiYQQnADqNeU7lRg
HHdkzCemkjsZFZDpqSH4bUMCWyxTOx3rmGsP3D4PQ+/QfJqQ6i3iNl/jOhqhidwv
PiAe28KwiPzvQF8IQ6oWUeYbaewDMeMSFslcNCMpH7j62eal8G8UVt9jZAWh7vyq
j3QE/rn7YYeydOQE6kT0381dEwjOcOh8e9orasEC5jFeGtJG2ZGhjaUUXhZUTDA0
1sQm7ZUZK2Alhu6kTaQ4TKnFerin3AmDC8CxGMqCiBpXRu5dxnJlKy/saVWdP+sQ
JBI7nt6f8EIU/uFFX/JX4GF2w24OIYYZ6NhFXKlu/pcewl4RhrmMWDXDxNpQz2g2
pHPcShhy/8BJ5XuXmo62Nisv9edr9w/xH8GOSDJUwmjRTWQ6Om39AoWaxQOr/j1F
wO7bPJCLRs7QXnU1iKWGmrB422gBDoGkQGVYtazUZYObyOQVkvegJszipOmKFrQp
PkbADRLuMHBJz8tUS4D9xTUPXf7IeCTQn4HJ4KNaiqVUIvK+LMpdVbR0+cTx7rgA
PMBQjGJw7xN7d67g1zdxnbm781DslkZQWxuUO8qWBaj48AUuokpT1P+A5AZwlmdG
6sfsKp+/hLJbGIREQgmsP2Dl2lH5bsNcxewJVkeh8gTw1W6j/YpHAD706kbV0KWU
jgE4Ki+fP0ZljZ3aFSF6gvTd4ZehQw0OivhifdAZ60ayHHBhnQkS9aTpzVR1DbMH
SIyZI3xz5Fzfn4jSYwRlkHe8USUmm/ToBSuRaY/ebPyZiYGtIggQKEGFlDe7Mzjy
okrfSfU9FK3G99flQj9AqoNs7s3R4nFS4Zi/BJFulMm2xpK3cJUR5oi7jM6XmcHu
Nj/uiVA8wOpcn5g/5J1qLJ4VDdRRc2fkdpeZtouVYVcnsGd0rJcF91033nev6B1m
oq+JHl8sW4lkvxbmHkvrIwDptET+0xcsHjX9WNxn1JATq6SzvQy8nfuYsgTb31nK
wBmUqGw+Kpvv/vjn7pFxq3ojkCmvUYz8obQxUp76EoBgFn0FY5x1wjA7tfFqFZgn
woQzrqy9N6y5sVAC2pHogVeQCjITAxh2QXaYPcjYrd9MmD/eX7DJmRmp6KaT71l6
eERTmY3aShQUsFrBCuBxLFrdM7fWXgXUTtX8OkrdTBmmT8qBWt6qTj6xuuWuwPcE
vfN3eyW5xeAgsjYI2oZfnypR7GzTzanrBxfbRHIvlVheBTS6rnWDRScnVhq7U+6K
Ue50Fbu81WOtgI9wJ07V69gb0DFyOAsh5cpoXxXg1YcxTdzv2lNy31EalOCyw1bD
71DTRtiJWiArDIgGuDFLkH2AZbXFIdjOCmUVu9F78bYApZtZm4fY0y6KEY7C59u/
+zHuKXZzaCl4eV4H7FO3YKneMjV371DxZYcB2sUB6aHa5ijjDzklmk/6mOU8W3ad
Z62TQKe4MtTvLwjiq6CtPVAFg9w76RC/2E/Q1NED+UzsfHAlTkgsg68Uxq9u9YsH
zviAv4k6J9gxtJhycKWY4Qn9JuTlyUKGjNDIG/bWsseApQR7fGo6bqlubfCBfCxz
0S5UR7yJj6grzsYbc3rAL+v54ORQBI7BS4UlNq3zWo46Yaad7e7zLxHYNY931bCr
a8pibzDr08St59tOA5lkZjZaZt2vHKV5oV+Hu2rOpubNU4C/oGXp9/gWneeY/6Vs
LHGaAzlFMosfxxKsjqy4enTQr4gxC6PDAL3AbwooJF9uWFiHxHuIi6zf8iL5O9R6
QSpiXMkQcXGlgRx9qaMT0Iny0dDkkL3iqI6OB5gCRUnz/SrALuvhfW5H3I9El5Tf
nSCvssJW4KCVRKpOujRUGY1ifADXw0bFgsWmlhuz4CCj8DsPe4jrt/40I7fZujJ8
mY3aWzSCsX9swxst+gdimgi3DO02nkbsNQ0qYM5S1/i92qaATPOhlzn0aQE9utCy
zaMns++UuJPlQzDq4ItR5eEMSK9L3PWDSt8idVtFglEAV3/s1+ADQn/LvCJHAXjN
dGvUS/kR4tpxax9d9jC4Mgi8D7T2pHTOjJGZ7V4+nicUBe5uS/B2W4MxAFsEQyOI
GSB1OJmpfCmEuH8jOZad5Ysc9c14VHmpK4K1mNPE+iwxedEqDC7m4f63tizxjYfO
vgI4PRTEheCv3vqYZvzbM6HmCEoDlScYndMX7wnpVVuE1xj8ZlDuRbwiEUf2yKgX
BRZJLZgp+22cjCM/qTq9strYRDfAbuOFF3ezhIHQAL5MHbJwYpVxBIpM4y9w5SOJ
wiAtYu8KojhXs0WIA/nHGBGDASNUVfPhKisBYBuug7TaYMBopBTVnhflRnJWpJc2
KgEG9TeYlbozt/tcw5QKVubeiI8GrdON7fGlIFCBVQI8F0pDokPyTNVXHRgQpKva
6+sld9xDYXWkyO0PdeCZkAoxvHK6Vpa61y4wHaNFZkXvkoxfGvqHcV+poWeQRE6w
t1E0exTyq8c1JLPDH+rj3f7ucNjRkn1PrRubckOuOCv15WWRS4tv6vCBZHHYms16
7M5CIwqFJAnHxrDCfU0yy8G/CHB6EVH8yZKO+tsNiJbj102hFV/8nes4Vam2PoGB
OnUzPoc6Zw645kPfSlZBc8SOpI9xJeV3gZXInB4XJmemi3yajNFlzgpRPJYTD6NT
QsuPllScV3eXE7aLOE/x/krQiqB8C6ECQ6ppOnAkpjEyiHUUWiDIkiowhhgoDsRU
LrYj9eCG3SvS0Xz9LrX9/yhM+IEf5boK1hgIUAoQYJgEPnQqljQqyN2/7RMug0S8
SZjhN23asUHYUgYFTA3VNzr5rrpOwGFE1tg4pGup55eLGc4yKIrmimaqG6VBk0TG
fZW9GhU7+vAc2ezM0oPOHsUNqY/IDHmJeuLsdTd0ie5Gi0Eu0CXk9+0XnQ2YJru9
5zOpzQ9Ns8AJH7E8sImAuuCQhjKMO444zneAPyNZEJuk6Z5Jge8PiQzCBhfp4Cw6
Lq9kOBEmH3uUsOAau4q1R3k98LDyOKM/1PX7ToNKsLC0oyjEa6v0kpz1nlD40/bp
b+YP0UtxG5C3SwPsN1RHdZS6opNCeqyGT1DN6t6h3eEVAhs6DpmTf9Mk3oSIqEtC
fa56RO/E5M8RWVqN9MwsvpXVdKxk0Ig3KOKjGakJUBwqFSfUNXkm+2gIeYZbYPdX
3XkK2JxIt8O46xfscpfREanctVx+7h1wYb/ibzvJxrbR5eRIptY0Lmbhdyuzoktt
4teEULKcPpfoxMAergzsqJQl9DFJwKX+BELYEPhGa1iXuMJPE5tjPIGfMFkRaW0n
2LAhPssVtZ40BGg5oxqrqS6qAyOYGes84So4MivVUzFrXDIVo5um65wGOBKRfwNs
DGgb7OwiHLoGZPG3vFtE68NXUGyXSNaA1BCBZ+mKyuEITRLof7Bfkbf1PtBrvr1h
6mzazXr2mUxGVCxfapQOUWpdeaUdWvw+72V3lTktv8fQ9KNOuPthhi8J/+JWsYSw
ibvNg1vgiUHdVESxc1YTai1AX5i+MIPBg2FMhqOTXV7f5mysRGUX/3oHFlcKZS+Q
R0Fbhh/uct8G4uO4wlU5K7RN4be/13fnQvLdyPCtIe1SLh8BGTAwEw8EFxg+qhCr
Tzfeh85mtn6XMKKKc77pyK+X98fXBfrAa8XtkYsQEE2/dxE67N92CSde68fyA1mh
CfOJM72RH1TzKquRwVunwlWLPZTJt7ew7EBqNkxYG8L6oHILlKLhsrmBi3TVlIwI
lYamAaF3x0MF2E8RYTaQI1RqjeaysfGpUD26rOXhl68VJJlUS250XSktVPn/A17x
kGllIvxMsmSrWNqAhfej/ZtkLQw3ZLPyG5cSC4jSNaZdDFIZ/vzKcV1YSnMYG+k8
6KEMiEuwUUWZltep/C1AY2XIgxmYcMznVom2ClXYeyEcblhqirBC9A7ytfjnOU0u
C5vG/gO+I/6zAh+FgXWcJu92mWm2V5HQm2qnrhMmjh/xrm20buc3HAfJPBAO3lm1
cr2IB43Y7SryPCzS+sUdQFfKQkzNm8yazrEo4wvop7cvTN+eMQT2p0lfZ2RZGiKN
YE0tqa74hCCwpX31WArk/rYxypHcYxjvsmCO/tT/A/rf0/fdErL9j5IxfJitLwmz
2pByD/4Qlm/8L5kYr9OtfdnnFUyS2D22PAXuCwSviJuglWaXY4sCN2P2aIOdY7T8
hYiRbNrUFCsW+H6y7+4ejO/zc1TpQMH5iq45SRJO0wrhRLswSVTvDd4RPb1sulUQ
bhWCKTl2ftimyy3xNc28XiULyA/Q1tN0F4U4W7khPc5bUYuFVd7nNtol8CbsdBPC
xxi9tFuvFXKlG7pXuC8a1kIInCP4u7aQMf8Ab4ZsfC2EQoRF4LbrP4JbK5syAYui
XBkaNMu8W5Ltc88AgYBS5Sl+xsTTIVzv1OHYT1tx4jEvjgz5Sh/gfeC/XfEE9bAg
ccHpJHYQc9brJsp6TyL6Bcmuuu4PrSW6Cn2Hlw3XvXFSawQ8GTL11kKh2IADjsWq
ec74nIl09yF/alZcT0Nvq5iRFRvbmHU+p5uRqQPBfXdogj1u2iDDf4qMi5XDyekw
uPTNueDkg+6tXIDPCrr3mOjtBY2PGO9bexAzWspOvFykfXzPsOi8G+JjphfLnxW/
vUcEswB86fmNDtEZA9DrDGnH8KgAxta3ntF4bMyoRBE7Ue5jhaBQ/rzHa1Ynm69r
UbVl2aeOWX/TYvY7R3iKRT2W/eRFF6Tppit4NHnH9TNzWJ2bK2392naFeXwUUINK
RgvWlqshtqsdOgV5xlr6+X7GfFrGWNXNepJwYiX6p2Mwuz7bN/pnvwrI/d0/5eV7
ZffOg2gSF9dAIqKYOQBXL9HUd9h20ZVik+onHTMzat9ceV7YknGqrri/QyPt6JJI
/AqM2t4uzi2ysykn6N2UZ+bXnVBWBXVP8jaTZg7V7P36DubNfuYgkJmJpu4zMWCI
GV2QYSNRBlegW2NpgE8AF1+1dMCgmNnvhB2ZY9Mxmgsb7+P+AJBgKsIXD7sB3UKG
arsDulRz0D8UVhnQNArTJgfZvUOlYv5dPseE7LM8E+65wzYnlgPcoCgG32Z/U1Al
ZDIDyhGLscD24vr97+9xsx4gKVmURB7AVCeHMwrwDEGoWoFR1LHrI//KRVTl7veN
0/xrbpXvNHOJWMXNi4/M+cWvWehuxlhzjlDlFsDTT8EyylO5w5YTi0loroOciJcO
7D+1eZgFEL5l6KBQQ4KOmBgp7uPndD8xZ886m7WtbKvHt72TilIugYr3BXuBcMD/
TGw5tVm62fXMF5KR0OD8YxCre96dpyOZss1VlCSR7IYPMM5AFlMLrleqMtqr4kiV
rEVlGyF2h2ybp/s30p45kY92K8My/pUjtIBRN1Uj1VPP0WMue4nQluYvoA2hL7uc
rvYvBripQ8so+T06dIzvKutFiHMHQSdlZY3ppumV4ZGC6dveT6wfCfk5QYYbm2HS
JRovOGXy+cl4UaEz5W1/SbZh+AV3y/BM3zY/Drn2QuZv0UbUw1PWPddw0Yg2i69B
V8B2qWqDrukFcQE2SX+8KA9UqxSH7J9PkpdvyILX5noykwK5LaIeI98C03I303im
a4yESyoJ9FIFQ10U+HDm1ECxrneDTvUd4VJyYAu+aW8zFkutMTO6kd1iqWMH4WuT
RFDWWL86CYhcxBXF+CCSy66QD3YcIMPdBZEhgplBBihhzZ7YptFLoapZHcARZngo
q3PzN3pKNpBdOFQanHTR5+vDfjVHGYRBn2RanpnCjUxhe8MSWpBP9/aXhdVacX/5
uTqJkMoQ3k0Hw4yNH/z9iXT5OfPRFozTU2UYsYFPDy/DJhTke5X1qFP8Bahf67pG
7zqLPwUMe1JWUcQxf5Kn8ka5WgVR+/JXr81Sf6TeQLWPqlGpYClaUiBPt3epSzTQ
CVuda/DidfwbZg/Y5NYE/sci5rXoiFA/20cbdJJdT6duIqOZHFJDj0IXZxZ7x7Mj
vOg9lsJ150gvoUFJkB+BXZGk74bK9ydvbimlk+qxeSDLDlwTIzVDQLQzIzQ9b611
2PPSFhbsQ96zALv1cht897KTAglNBxE9wP8qxYsBFH61ByRwrkxdWIlSY0dFgOO3
qkFzfXz3A+jyhovIbqRli2nbYOJbkw0U6asB/tnh9yy6ru74FH78ogGWOZubCZe7
6FYw6kMhblq0BAEyyzqKhl7u65m306nz7pcZzM4J7a8nE+7xnLmi6Jfh3/GOJ4IL
E7cgthaxDAJx1aYxAx/1gvYzWeowaAPMOjtljYeSmc8nh6p6lclwwPOjnWQRaZta
7/MJt3Y8VaeSfD8O4eO3oaK2r5sparFJOMTlhFZYxGVjX9ShT5c4E1NWlitT97aM
cx46O7xhGNNB9AQy9pMJsp/Znj/gKdvKM/0JrQIgJa/r5YhpvED1Lt3rBHTnuFVU
P/QehWqPGsny8KoqaIP/zpreetf6H7GXjH90l3zjsKVBxkySsgsz0C0eugpgsEG9
wAgkLPpI8nKCBYIR8Qs57SOl2fveYWdR3BmAwwqxK+0BKLxN+KuHH9rwMEcA+/PP
pDEmn1lV7ucqMLyZqTzqaFgvLvtpLbesXOALrKyWc9f/jlSGXV6g/DwmKVlE+vYS
qSDW/Tk8I026gIVyx3rxXMZA7kqRClhNHN6qZzokVkWTkKlQoNyJ14hDclkgNEj3
EitutuRpvlEC1Rz6pELzBK7NAq9Bj0PW5vz2q2y3NcGdQhb7fW5aCEfgqzJm1+aY
LdphvpVFkuqV9ujvV1ArzQeMaAe9sa7XzsHuqwslCq1yFPawbruN1XgIBUle9BKk
U83Ngx+IDVUxUS0+e5Y5qUNclKTyBCKXu02bCg30x6ABk8ss0/pxOYdjP36UGkId
IW+NdTSEZnaUeMyWDTC3yr55j93Pg5bVC4/CS6dcdaDComu8kwk7XkF80lGcEu6y
1lMdJnKLQ/IUVy3vklwRukagaf5vV0BnYEIgRisKlgG0Bo7Hoo2Qqss/LjWXja2k
v/YjHNlB81bzRf+FM2K+M37KEwIxrk+H768gInQxeUKWW4c23O9W2cm8mpDtBQwC
429QOqTP2V1YTSJEmhgY+alUV8gtYEwWw5+8UyxO49IOC6UwxI8JdG127V1cpQM/
3ThWPqB+qU1CZyMJIZtotOojSwN9/BGcIH2LG+j+EbGok8h/q3EFKw9gRITJzPBT
cH3/VzQq+b0RjUrXmXk4Blz+YJOJoTT0kMai1kc8hHK2mDskriL7nF9dyhY9NnQg
OkZc5LIbGfu1ITc91Oh8RumM1VaajFnTMYtRL9Qoza5ztr1dymBk/oR/xQJP7kd1
ThiBQq7MFRVoTbpZuvmSuNkWZrBNPFnq9sEaNvPcsgCpCVl/MD3BOpwFyCOWN/iX
UoFeh0l1ZSmtJotvLVf/3lvah6U8mjJtQI3+xL7nIXRVbSBxtFckiQhOwKo4kJHg
28kxD4YPZjD03wiZpkAiBja66PH/U1B+COq89tKlRvteUxgy9HYZyPiyr3DS2x4n
xF0uJT32PU7rs9PTIOYVzMebn6STjYnE4bSvZnxmQQYhSBLybNowUpoFnMYuLkaI
0Hox5eg7AqSGR71y3XcbU4cItweoOFtofrdeoVUtjt9m+GxX39SDyLvxtK+QPt+J
3sXM1snIzDBe2kw2Pk7NwN6yGF2Hu+mO5c5gwgtFRyitKFVHs4Qg7Gb+8UrLPXSU
FUbTZZ+WKCYlgX9h2sHlV6Zg8oolK0BOIMHqT+xGKIYTxWNI3FxnwsNa+Vn1+HYr
Vp3TO1CuVQTU8iZlTjOc32mhAFL/3k6Eo3gFmNpVa/sfdtY6+tAwuYMkbqnRn0qz
iFfvId82AslUmy7aRAsZX8m+BN7Zl6NJEyZw+nphw1jz7NH5K9qPQi4JUkT1tM17
THsADHlG9sgQiDZJxOhKtJXAPsiOIgPrBISMXg5zgajMh7Uv0uLenDBzVn5cOraj
LnUTQYJcZfjnOnIfSwVnus5AmCYfBn+HnDk7adKyk6PXNmG5pLDV6PuRECzi5E44
7YreDi2Ohnq1DXkLmRkhXhizxBsjD9N9fpwG5SAhcePNH+Ua6AfePa5B7ix8dcg+
jV/mkNhqVn7x1EKdfgGx6roWI9J7SSpyde90OAOkbdTtUnh5f59TL+ceMjXZd6YZ
4+ECI8LaF/NWGIFzpiEA/TSn/LOR991chm7kDUu9n+vzKb9dd6VwhEdM1cFwAlJX
ICds3peegH6vK6JXX37sgnPViC3VrB9SbuBpD8hGKd7GaAgpbNhTPlD0vX678hwN
oYe5DpNoqaM23qD7+7xxkCBSSK7mfyHsKMxe3QpLF9ogIeeblBX3Sm1vajJgdOXf
WJxs8sSk8721l5lGRJQQnbvgyJ7u5XZ5N/M2flazZKCwNC+tMt0sKyXwk6YQOUFx
rBWgf5eX/FMpSQ3CT8pLI8hWIW0uBlyQ5CV2hxzQlEHLhbLoac9YchcXLW/scBdc
8hrigvsDaHeQQVMyhDXPInm5L9ij1UYSdydZALEKfoSmcNVGYHRcmGzCCbBDx8PW
r/Fkr4MzZ+Xf1ZFOSMLcHofp45n4fi01WaV3iAl2stpQnAk1vuNAz8r50qYdX3W3
w8Qk7+kMWTJzrF4td4ENG6ZEpJtOhgHXgwKtoL0HKUmuCIksoOp/h8AIhTop26VN
oZy6+bZNouEbRiVfDGY0f1mjNbltu3RAcVhMmQ0nL5gFHzy8jXsaEjshwD8EhjjC
gbcInxhRT6xrW1Jpoddgd4vRgXlhw8L9iDusix/pYqG2qtvllZazU9uk5rBmLiQF
WtQdUu3KKDc/sP9W5Ka5rgbzMyDWyIZNyZm2u2eFnRWPdHfqyvxTFFWcLo/3CvyS
U1MU2mlpFe2lUZTZ6vHlsE2/kt6xBVK3O3A549wMP6cZNfBbVDkCRIUtYoPm6H7S
aqH60jH9JSb2lK0syHyrU6iQISLl2Dx+xOBIJ6sya1aK52fvxbCIzrEm5Hq9L/lG
WThoC0GJp9iRGw+gHBVfy5sDojPflyMO14D08hgCetQFDiUw+UPeskrh/fWCje9/
AD4wDsCPFIPqsZhtS27CB8wdxO7YYjWnZ4GPapfBGKd/pkmMdwq636Ct8O8nHGXk
gUci84JEu9fm9HNC5BaT4jY4+HnHJBSDrQsz0gl9mKdcqUq2M/QFsEBbDtaRv3oC
gNx3dtL8vsQ7cOfNeWmKGbOMt6y/K97TaEqi0s0Nfuo/XoROwMG8VEbhijuL6fDG
IL+Fk08wFqf+K0xYx2xGNU/01PrzwJpEw8B8Q0RcBQ5KXWyag3dNrMQFTzfBioDd
Q887wiaTIyyfS3wps4/4BwLHOhGtdego9g1LtHWf45rq+gBzFFhrLztwPZijLG7b
p23KJ1d9D8uC708Ed1rIpxDlHAhd3OVZn6GTZR9PSbsoE+ncnKbG6XYtuRsdJ+iN
bDb8pfGqd5B6Ys21ZRKRYPFhLKfRfKRp717F7aJLVNttzTPiTtCatbYAh/CHhsqu
aubaTz/YlNms457AnJCix4n7o9vIF3W8z4gylEebUbkWPFyPeYWs9/l/CCFhwiKm
1BlALViMjhB4xJ+9i/gfvMXLyeDeZ6dJXbYGJBKk64WPKGmu1qEGbOQgaE1waalm
RWfPzDQkuZcBGuSXKf4kxTjXGHIO91MzGXPQ8FzVeUD1Xk1JFVNOI1dqjlx8/9Ij
i69LgFTidQiXgstN8ZGEuvhwcCe3M22Ejw0WGJHFsG8bT+yb/yohNbiap8UwUfrj
ZxjSbdIaKUL0/80ik9f2fiDtewo11HmghEQG2F/s/pBxXmJEhHIVldEzH8TATSdB
4ciottUAEPfMPPZZUuRa9K/wt/4BJhS+UjijodAqIgVXPoisGSc/4Kw4745BNr7d
O+JLNL3ZfYwyeMz7lpf+xPOO9VkAHlGqfj8nzZJj9dup+LNlsT5KmT+BRj1SFwkj
olCpb2YkYZbMWVVWqI0+srM/sux0hqTi6TmKlzP5Q9kQ51In/Wz0u7Po1RLfgK6k
x7UBUhj6dJcb9/xHKpAdS0aQzwZL8cDoQIvu88d1ERXiQnHxuBSffrUcaTGa/JjN
r8TRJ7A0Pzveqpu+N1uNzK6Yf77qHUbugA8urP/q15cu+2ktKVLxihiMP+28IapH
aNPWpwCnYNQ/EYHfHwnz8aXfFnXiY4xcPghlIyhpx9g1KA+Z0m7zXtTG9rT0SNlN
v3LD6NOBa4KOZpUhpxytTfeWFeagJPwg41CsU3BDoGjisiUfMbXdTyga7CQ2/sSq
2p7KX9hzAuhagW9rGyKpqTW1myPqNio6xGWsYC3SkKno/JKZ6Y44AhZMdL2UEPN/
e8U6wlbwKQl00fiTzZZqq1MaXnnrgX1ixEc+jZwrA16n1xKeHWijAR0a/CiYCQwE
Vy2BPKPJUWJlcQlrn9A7vzgsakRNP5giY4aQyXKz7c6z6m3nIJ4Evzxr8pujR6zV
7g8GbPL1DzNutWu9IY0U4UOF5emLjdCnF8PsfyLqU2KmI6czbCzjiJz3Q5nZUjPm
M+sAkVntKS9ZdNVeZQjgAMkxXv9a/2cDrcV47JpJOeAHOOM6sfT+Fku4BxmgvOSY
fBFReLr4m3wQMvNj3X8H6bf6xJeN7ievJDfwqzFrsAkfR9WCiitEJ88h8iScu5zJ
lGb/X2ZcHJ5IaTh18jrt1ZMAU0IKOtoLGX9GqevQKePPJrHqmwa7U3A37+o7d519
Qbx+UwDl2ajVB1e0UzXV0a/aNQ3rKZeLaFJ3oIBTztvQkauPeSdZ79r7+/8Ztjl0
yNpWVy0ZAWxDi8ThY7rPrcKMY+NxUC5e5jZXaUNPzes18gh62AUeYRDZH/qFGHNG
mgC+7ARkHHWcsBtoPPJ4zRAiVNl4ajQuLFPag19bWWvlqTJ/ylfgRj/biy+aYdvK
zrGFAp+Ev0EsPSYYFLCgH5poski6e7gk6XkvsiKDXZff7zBjJYgIB6dRyGMVEUlh
Iiy/QZXShNyGHxagRH+NvoqAVW9fjUUFbgso3tdwTtbK8i4uay12if7U00qFR7c7
9z4+cjdKQJJOl4S2OazouIfqedxAX40HsjkI5oBUt6BBnh3wUIf34sEhwy1IV83c
HNciQqpCUvWQysv927XcQLayMVSX49fT020u9BDZmBMGNbyChfsq0yvX+FSoBLBi
QtbnGP3y0yfK4v3aLAWwnyDvL7YUqV5/4ePr/64D7rIJDxzwW3Qz09sMMafHFt3m
HuXR/grJubas1qa4ddipVUKIezXnq5pB0Jn0rFBqKgyLVModzRc6hLZl0SYsgoBm
CU54l5BTragYjaAA/xk+sLbufZT7FKOJ5Xha8T9RwrvR4fMOqR7FSzS8C5ulWF1z
DQnM5N1SKes4Say1N9HhAhlDTBGW4PuQdTE/1tjz3+KbUt97V4luMhmQpPFlsMVK
1GUaE8zlC3HT9MVo0QdpN7gfTso6klb4FzcOXA35rPrWOlypVzLxD5iICK78cNSP
rTAThhDHNPYogRfWkD2UquIIC96Ee+CiNbhjvo6Dbo4YQwWuhasFSvO27lNqZcly
CJBUGllOuVE6/oMle+gHEYU10Fyxoi4ceMjCoXLCvcghlY5AdyozyE1UMq8cJhPJ
Yue/fCY6t2dSzUpo1et2SX8tQIqmiLKqGvG5OHtxURPxyhBJ+s314laLKWdPBbka
AQQYVNOqIbHxcyMy+wnmmJ4ej2ShtDqRN7vOxP1VR0o4IIvkoMGscRxyk2uI4vjF
Lj1EleccB+uLqZCAK/7tO+es/TgQt6qXUx8/TZoNnVpvdRrzb7CryfqCLGQUtR6g
1SCpKZ+UpBTcpSOuJCv27izxkKmXr19xVoy419Otuj4kioDqxVx4VfxpfQ4J3EAd
bvb/gH5cPxXGu+bF0N2crCeBiwTsA//QxEAuqo3pf4A2hVaI3ed/tiMP8KZdXYlW
iHbbyE14vQUU2e5HaatKFmTVM5P/4KJBF2DEbQFC9TjvB6n/x70VIZ1GlBmehAM0
uPdCfUe5bn5/C/mgBWsAcFm/grpEul//cSha4fTdJcneyEXp0JvNXKa31iEdYtZ1
VO8+cDsgGX1mPqNF0kRHyRXMElwfipvRiL2HCLAFUNLNYkbcwk0iOO4hwuWmqDQW
ImEAcWsnOd+iWDXuPpNn99Q33Gd9H1hm2d6E5JO/WGOJqWnxo+CfdAbqOJ56aUtx
3Ie64Nus+wm1S6W7lumIRKrX1ZFroNWaU5XNJEyYIoH4PufGwm0aAbKJo++Mcyxw
jV2p/ZpZd4IFma51cOXgxNYoMJ9p6PEWArIwDYItBe7M/Tc7ZnL4/9pOqlsgLXs7
wgKn23+zyMWILmMDI48y62pyRda9BYt4iZMkz2ptCVzFXqUx+Pb4xH6AJKt1G4sO
7PLJlp5MB8pSyDiCCO4ViTSCDWAQzzKAFZxagbV0yJQFV70o5gvYfV4+w23a0Dzp
KNzvp5N4hF2pWUN+BoVY7yqr/aNcS3hOn09R6ghbMTaVDgTIPCdC9AnXV4gZkfbZ
iCYUd0feEwoiofX7450+MjeGptzFodSN4ib4a3Hn6mkHjY1CsQdtikuzjp0JaEO9
ZVElZBwOY/7tvncAJtc+8PvP+ZMnjd3seUkP25Pj0EuJ7KieByNnEUrI+i4p7vEn
OlsxWwKgyaw7Wz4vFMHTsJM2x1i+9wX34Wa392xoQBj6LHzYx0c9wvKG6eRsXUwQ
0kUL2JbeoTB1XdKgogLgBPkhWwHRIIYEsEIvk7xJ2MUaPApwzbm0mzzNFPlyfewc
yIY9/jMHMPF17Lb6bd+rnHoxv51idZurD/V0Xh3Ddq8K45spDjmkVYvkU9WSdXx/
6cTAwcs/zkIHfF1s+CoE/tmkfEOhaVGZkyZLmvTOt2ltwpjsAHTgoKLLCa/XJloH
uuuB06h1sdA0AlOYjrVw6FWCU1djhsjmnC3LbCB+1830YksAq2eU3jEaTSrNgZEe
XSaPfzp89i5wzYZkwROZ+rlyt7onYJN4o9jmoaRhJH0R5PUDwqc7WcdwvZJSxMJ0
tRi3EEVThfg8uPSl4wL0ibmnNZGWoqZKT7liVjAtmHZc8M3ivoviJmAIwBokOzss
yDpPRM85gswTyJctvLMoS5K6l+cD95eA5esgk599zxSgrnNPTZGVPy7e8sXlTrzM
6pyhZCWiyuA0Mnr3yzRys1z0ET1Tm15QGqobYFc8MSuMRxPC0mCV45LLEiBK8oG5
mxll99Rx6liZugSRd1Trx9ZcrN9LtMfsYBmfQu3boTlF803F5ZIq6N1ekz2of7fS
/9KmtGFe0oI5ecKa8m1g4yI50zT05p3PnQbCKizMT8S2yJGPTXfN6dWrAt57H1lD
6QnSxEX5KExvJ/5m32h024aEmdt+UjuSok4j2lu97UFA0Z2XUhupI4ItMwloLVeV
tZ+5iy/79LzONNDAyRImliuSYqxTZwBvbtncZS3rp/C4CPfT3Gi251wbnTemNdU/
GOlePLLTWLqUP0nrWdZhslgo0sxpefrgPIR6HwH1UDeQBd8QSQFeu5Bt6TCfQ/yw
ITaTq9iUlw5Jp0KCJkJp0Rh4Cfxi1RTmojhW5fyJPHdZPbdLkeIZZrcCXHV0aId+
Lqt3857FXsgl1oh1doh+saNF5byJdZbLJghaAX/kgLlTKRhtXTTMzQzNJhGk5HdO
AeCL2p3tGPnTbp6D3Yqd4HLVAwKJ7XXarKXbrAi1bOgMJ16p10tViIoM6E22XkzF
fe8tmnU6ncqJVPnj6XlND3BhGszMQxF+uSA72gFkBgs+5HNp6FJr77fP4z5mg1uS
20ojAk/jmPjg7om3C2rJ4FpDwZTVdbdujolxJvtY1Ei0PaLSG0gUZizWszr023E0
MU2qVRuVXskMTzPl1uDxrMJvZPLxZ+O1ymLB7InWyEBU/SfeIW8FiDUsUagwnSgE
t0UNZct/wpEnExEnpCz+vYcWVxnp7OhXfRiULj8p3zxRc22C4X+OQdMsrPhFZuYt
6KUx+uB6nNritJSihqHIyn8dEBbKqUHLrJtoN0jRXkl4GU09YhSDpJSB4uryQJ7U
MVc0yI+occkxNroLnX0bxJ6anHndtKlm2K4+mn9dgioJAU/UHzjBV9mlDW1klIve
C0t2G3la5Kh9wFPqbN8VS1SI3NA5dLdtx/mS+Y09AUexBrcZn2zuey2zgSsZH/En
OThyxEfb4KPhTLPgSYbUyQbl7MsYSrRgyg8nMsSEBPfUwD2JV0zMTNdeWFcbRH+E
Ns63Wg8kF8JYLnQkh4cqWAMSSTe5djioezSTIhpLLFerChDwsJMO/bvHuWeom3hp
y1N/lRny5dpAN63Oi4z0jABkWjINzWPYxNx8lqmmObNK/5XyamCxC2tA4yXAj1q/
3zEQGa9hIvV9GvbYafE+Hlnh/rhlsYqixyUsWVCxleh60FyOsBXunui5iiuSUbrA
lrUBbOEb4pc13VQgw3LTopmcYJyUaPpfhZO9QYW1rUWUmEoyLzOBcosX/tpIbqiL
2v6Um/bgHUDU/iOfldOP+Jh9fGEd20umHJ1FaqnB9Ijko5c7B+vAIAIatcvR+LLZ
yn3aOJQxIbdmiq+99Hb1o09py6CGYUPyMwKEwGW27NdTpSqXwFXxKB7dJGBRUrMC
BK1aXFLdV7nGsTYdOcOADSYhbx5B/MyCAjcB3pV7JlMPp7zffquyNEDEZtwnb7vf
utIhl9iC/byEJV5YQK03N6/C9vmpnvXV0A5ugwyUn6rZI865l/sU4EQOahItV1wi
7KSA7y/siaMOiuaKy5t7vxYKbSR041ckWsuLsuj1rb6FfPGoL0UpW+ShSNNIpgCI
d3OLsBA3qsHTwU418Xakj/mCRs2JhlPgIR9KZox8MeZkUMMHqQv3FAHjmBQKnAsb
iGwhgUMpuHwgt1IdFLHAyEvKR16wZo+0vc+B5aKlIT3GGe7qHVqWhTJkFeEeNvhB
6jyJmzdJVoVuF6zCOD+swDuE4NZgivZecVdUaQVMWV3jZbj/681lkQNIjM5mwhxg
de8z/vch12shbGvwNqp05noiiXbVQEPXML52b+5RB5P4q+Hl2uluFXLTdfitaq1O
JT58/SB+oE5tNVlFXIHua1Xsgyn4loQz+7Z5htp0JLqPYVcRPwCpUjX2r6C9j3A4
PA4KwqDeOkud1msXn8vD40x/BrvWs80OxURmEZOzzfgVDYwcOfktBcMCug6nY3uA
RJF4/oroQN2X959PjjEguimfBYjabV6xhX3RwiU9trwBpFLgda3iQrq7+apKE53k
qSCvzj605n7n38tpmlrVGy1HkNmqwpteprg1++cc1YxPkTda38GBgN61lBIPQs0i
f4xlB4eDTSSLNITWsAI0MdL03JLa2Gk5i0zb7UqMDhP7NSmrvHjkUXRG4r4rr8Vp
XOU4+9Y5RvDSE17IxP6pWwulmKN8g5LOseBKNNaeJc51XFV2O+jww+/5m/pMs50m
1CEQT307EmdgHgCoEV6zPZMst6u4Qvp+NhNDuXlyydGn1WEnCySmOfNegnArUa2N
yVTKraCwP1wuLvV9mzlksehugwm2bRE785EdN9JRmDZlfptyG7TtoFJC6QphPF34
Wwn/UZnDFqREmDuMEzSnSEw0flo6ldDIVtj1Dwf6wRPt3v0O7Zy8uZo0KkZZXb5q
Uo6Xk/PnuwdD1a1iv6XVI/t2A9+dfbeDLy7Wps3ruuFvmjjsOjHPtgnpKtI4FL5e
ZXu9OLaD8/3rx9ohvRkYNWWWGIig4GGQqcvg06yWmgSgNS+YYojULAQ28D8cd4Zh
OC2LQ9AP1xcx58gN5sHr2F6ktwtpKw9yWzuqK29Qwqv3md+T0VR382gqelvI/5Id
bfhEQmxWDGm/OalLlLCXyqWRDojXvMzTtP/jqm5BJHDerWiVlNRuV1nNceSuVJb1
APdmeolcJKsj2HS6HoBRkF+/49Dbplbpcei3loC2+5GUU5ZhDwN22cr34Tpf2B43
aKT6am2i9lrNo5gTGpdzm6Z4IvvwgaU4w41xUBwkRfF0TXl1Vqmr1YJk8YcxknMV
TY3+OTSOxTd+TGorw1gBrhrZx0KOnEQeCxtYUSST68DnqURx6X7U8ocJ9OoUN2Rv
Ml7jnL97o3KFlJ1oEPaW1rL4N1vf8Km1fWHMwG2PBQ4YLaMZXWKX6zG0tX5qW068
cuGQPfrBxte7iYz3ipwsIxWJWGqxLiuSUTyeYpdUrKD+lU9TDJJvTLbMp+f5O+U3
xXK4qWCd82abXJQsHazGwTJhoeKuaNB9HnVjS0bWdJTBHEsgkLj1LIc8AnD2QS4d
uCigmzAPnvk/HPPO0EWQZuBIs2QR4Gq6+pAMLOILHpl4hi9l/H1wqOT8SElW6j9m
NVxg1htIc4Q9AXFpljCuZs1H9aqEnfMpnTSqzMPSkw7y0R8825oGcO8BUgp85ktw
m+6h3PNGqfJHvV4+v6jHXCqHzRYaIyjv7ZdEQUvIb/K4LeF4FRx0KHAwFS89yiEM
HsOAibAiy/w46pS2hK766++Y1lj36j5OVIu74HyjqA7H/KMZ0ajYDdH94bk3L2Am
bOYv69Yw7VaZ1cgBSTted597XJ0D1Re9SwiYIkU6HfcF5kwJPPG44ILbE/IWBC4l
7ey5nG5eJ2k4V4vOlI4eN/2IYtHg0cgQvb3LidreB8UnC5hIkyGMDkWoGkdhoiER
jujgOs7Hf35e8w5rNWPsH0FLpcFEFnW5hYorDv2lWsvtIJObfOOR5VzQdz7VhvWI
l2oUbJTmcXwHyUiksvshyGdnseKbY5HHFALzOgIff3vUCqB5aDrsE0XM6V6QKYv5
XOwofzGLuS3VYdZa9OWBzgHH1zlChmp86IYxxDgN6jeyp8kStbrvWPyBcjZ4Ssy8
LybS8xn9RSkw+E2hEEQ8mssJg0QahU47GBKK9YqUQgejBxlAuTDF8i+NCFDagrW2
JoCiAiInNHjMVt69jU6FDlHtiUJA1lY45rJiPVR0ARbwpMR+//7aaKjUnNTbJ9w6
7EmE4AyKQbNn+5Nxf3ZlxR4KIbxWYJNQId5oXK4aQm9dZJ0KlYXd+WoghhynM0GB
55YkQ5beYmSWOsuvtgN5/U3YQaj7KVKLAPrX6aor4DdKoW4t/TcT5tLDLiliXgfQ
OnQD1Og8gnTOwwuUWl3F1m4bZSlX5AF6JSS7N8HdowGg+Z8tVX6u1CwChSkQSPLW
YnPV0kaaCm5+T7Q9HsjXl08LMqwlUox/7DWKVK7+w0aS/bQOa8TpBM6UXd8HUGKz
SNgpmM55XvhxAgE3naU8dzwGVuvgptPSfXc3/+3MB9ZyyoASv4UkGVzqOTNJQpMb
xaNoVHJ22AuFT+DLo2XUExo6uUQIU8A92FJ4TwRUJ1AGuv79i0801ng2X5yEM92O
vk7xGusjhP4RfJUIWIRt31vWofEH/wtpqBAbthVPdq7SlaS4O+Pgx4IJJaZ8Noq9
kG99n3l1a4cCYVtjdhjxLY2EsmUt00LEOYZnV7V1qTP6+S2Az3upIGnbvHjDLKKY
GqUqyI0K3qJ3hmAdzHimDM42pXyDxbCpeKDqvV26I8rdfwRGLQsWi74XtsWbSAit
3p0x7iHSY602g1gpwq7iGttLQf4ZwFPDP9eYo57e3t2Ix9FZ+xCWwf5hmerjnxS/
cktz0LNsH60HXdkn9Cw94sjC4g2lOS/Pyf71NL3NU/q9gWcIOTgFbLfuff3cOJcM
i2vO4mtC7Ie+Htllz8gsLY+cHG76a248sd6MyZqZqpxb1zvl5ZdR18982dTWQDoz
JhqefuxB5RlgUPMqQpIK5EZPXdoF9/aCJDtTSLMNw8Zt55CxSQcn5WdG3S6/8clY
KgCg0fR2pV8kHaFpEKx/xLM9fvsEYI3vvtTQqJ58DdIWFvkYGSi4vgaXbPR/9/El
y7FAl2sM7QMmKPcH691LisIBFH1aqZ3JC9dEVBQuAo2ayHioi+AqF7RO7FLcYO1P
WYUeSBWTPN767a/h805zYGRkuoNhRpUDQxBk3adrvMpK2dGVjFdhuyqwOF3eddfl
9aDpKb/YCHaeQhFACJZhbMXq5lzJXhuF5YtLx/c3szHzbzeL27FfJNfvDBZSIR2b
h1iQOroH4Vt70L8PO+x0iEye5zTe/h7Pvy/BMg+YBc6JbfKVKKg6iowFq291FXoM
I2g7uc6lEWySIbNzRaJqHJxkZWQjAxI1wcCpPY+kgcox9oZgwOaNGbTpav2a+tH4
nkWRRamX7gTgDUeHI0emBf8jFGI9rg5+9E1vgV3eJbb9V+mzKcEDlvf2IlTKonY7
YkqP/02tXMP9qMDdJ0+ssksl14aLyQ0zmb7Qkw0Q2v4bE/X805zM+7cRf9MD5jn5
1JbPfm+PG7+1lNBM2WuWeTkBpRAcwNQOyV/VPmF721mlAWjkep/fxTVUDnFJgqTh
1/tYKYXMuos384v05qe7upMMVOU/bCU+ySAONyxx0tlD/wOKmwzWePQbw1pobi0g
lR9XdhrDxX0tjnstT0XxOrqBoku7GBXP6OZGqjiwiubzweBJfa8cTJvMp4xHMhaw
TzBaVJXquoSnaUYxO5yrixeDBjGygyFToqHOi4JRb1Ddt+KmKCHEdVrGv62bZLnb
Lim3AIqMan5CE3LUAMotiosLNiCk3EzXbrkgDizQxJhm5bcHhC2ZIORlF/V2bzeY
Ox/3yzEKAjA2lDrPiO8hH4u5ZOh6oIvZDsDgYtmB6iibpp15NlToOTCYMkKNU73x
rQ/xa1qt/0epY3MN6uHaRbXGPeqNPT/isSVFSnRPo13XsZXri3irp+HLclEXagPS
H9G5wS5W1V7TeNi7R/re4GCkHOxhz4KSxPOBcX1eJy2q2g8eBs6uH0OgYJrDvIv8
DMj3OPjDB66YVRpxHmhyQYAb+KDN4SvJZjIBf0j7mZIIot6dL2i0ms7IpzTDmlEG
xJALw5k/1Ac8OI1QQTson11cOnMxISM2R+Ra4yGClMZ+jp3G+SLQ0w8e1DvlchMV
RB4XVerh8cwjoQXymnDTnU5ZDUq1dLmgwFEP063lu5liavmYuTbXCm0ultgLguRD
DeKeSF5fc0sf48U7MZYekaci118gPaPG2XtwxfQMLmEc7RXP5TqZlCSrOZGPqjz1
TZyfkngb1FE9sEy4aqyWfCNLI8OSN8dk4WdjoT5mlgCb4ANKmbT0VZRsoEPTshWI
NK0BSOOYTX7PTX5/g7Zqu/hdGvFJN8oYuLvqjEut1rdq2Zrjl3E85h8XSJqYjMPt
fmDwuQ50wWjGLCybFEtStJRxYXuD71RrcoWsvXjmAEZdkxljpwV0+WLsu1dS1mJa
KWC7dkRVaaIVDjRE/C8ZPJ80Mnx9Z0yFNiRJius1paaThSJCMbQWH8Mp8wV4qmk/
rzZch9o2Sv0+7nOJW0dFo/vbRFFqcDl7JsnDkhqgP+IC0mwEd9e0G22zWhAzUecr
ALd5PAEsPPD9kASr3J7KrmhFKrRWtIYGAHFmJTaWD25LjulkI8VKfvy1fB2q/sxQ
jOrsgJMSRvauW5QAsUrcAiC1rL073TS4eT4YFHriFc8b3bVl14so9dlK2iZqJOfm
YvInYAZP1dseLxxtZGR+2+hcD2NsMshrrqeF6RkrnK+WsHwe1w+fXIixjuecvnJy
4z9GLpyqvtzGox+Fw8pN79WPyK7M58iM6ja0+1ROhYlNP8bNap0KEAaVYubzvawG
+t3wtu6Q2L6UytTlrCEx+/PeE/E6JTJyoNYjSAomExDHWGEw4v8NN6v+SAxIHPgP
Gq6Rku2dttGIGsJXOUvqUB4C9+K18Z8GwajvOZVxc8F0tsu/uWAq/Wntrt8WxMfr
8EnC0VU2GiO2vrOMuqUq/M3Bkc4xnQbZ/KDO6bD3wdnJk0aFP2t3fBXiXuJEztJ2
38hEKC2cZVoEy/RMae88USNOQN1amUoxVz2TAXRe+Bb+y3bz5bvwLeXn/aIk6oCy
Sw7IghFgHtLL2URv4dGzFPQJ7kgvH8tjOaE3kn1/+Rxbp/soMwDOtYW6TTiicALR
GeGhy2T+sbS71Q5qM6R3iLbZioLgTgJJUr63tub0sqp7RJ27+UW0dM8AJ4JJ4LoW
bz2iKa6xOuKiKzGXnoNguf0LzUPjS8SgBusMVF2tMcgr4kaXrI8j3lj40mLDgQQQ
TdjJdu41QQ4YuaT57Po89bVJbE7xiYPYS9kjt9xVQyYHy+VrdSRy+pHQ/kqMNUec
0VAbf+9Gn0KFHHYlJE0fyQljgeONf/vLFFxgL7+3oKFBeAMOyKhtZIbYZoFy0hoe
iDx8eIFK8HtrqdDCpyJ48T+NCG7It9kt6VJHFlPk59O/Z4g4Qhv4be0H3oF6xmCr
Yhc0nPTpDvhtJSaX6nQrYOnf0aAsg4jMPTOSS+RnKbVn4TdPb0VERkdYRKx1S79n
B2xTFslytEj3WiVUut/2qERjesMSSYrWVZmZXZHkDkyUBammNqIz7BqKQwo2Fd2b
ppQUqO7Aty5OoumtrgjFjc/kk7mlz53Y8dg0EGnkS4NwewVbnXwp3Rd5oVc2L9oE
iP9qnlGh2P1u8SOV5AJVhpko73CmzanRMmfY8tBJrnwOLK7fWEGoKJwtdENaGwDr
ThkWBWS/BnISiLlkp8GxRi/du4ZGnUIqiaQI4SCsRKzVgCRAyWeh6EVheQOOWHTB
GoXuRk22I2KXb2tC0mUX5TOBXi8Es7rfT0KL1lnjmNx3Q9W8JiqeJ+qURUea0NoN
vfiO9cPbSpgOYyK2feR3LQgaS2AAorNCVxy4ggl9EnJxsYMVfrIvb1FnfEyLcu8o
CnurBXBtOXTpm0GrLwsGZxVC+RjGLUZwV+62aw0BrdkA7skoNODRklN3XLhqshiz
u7S0XYv8GVZcrN73Jv5z+Nqm+GWICwA8X1BzSCNEpJ9tog6jJw4i71pTG0SpnmA0
0AjQb01RdwYxij9Yb5gKoFUIvlGFqLejvoibLdSqoaz9LblbciE7fo7EhFhnjgz2
Mh9gb25a0VliMfzthzlxpU/QwQZgLU1ALH4zR2cXoVImFZuiJy3rNcMoleA2Rgoq
zPeoZHR5jOTm8G4d0ez3hgjdWEcGH+sOZyQLtlAmJy3g42C0uJuLYphbIAtfBJVO
+EUck+kkl3jzbanh+q6ZcflAb3TPUXZHYLA1OglQsbauRWYNNfE0ha+yZXLOtIMh
bdNXlucUzHHPNzml47Cvf65xamCt1uoYVno+J284JTEUDwdX919zKeuHOIYKRms7
OFj2Ux7N5wm34McnPUFd6bM00NDrLLYzzpuZtTJ3iy5Xeu3QhA+DnhjINHM0XVAu
T0mdm8PdqYj4dMaNjhD9g9XSZ2QngZOjyw3a+Qho6HmKy6wBl2Nd0LQbKC7S4UsY
ks4mzusS7VD3oNyM0PkMIVO1j4XKbGv1H8+ge0BKkrWQ2azKNVNmMRaDoSQbAmzs
t6drEOch/qvuYHljy6GD2QVPmXrof5kPlHmbvXE7QOFFtrd3woo+Rf3qq3qjN45O
8sh5F7CSZaK9B9cdTX7k3zR7tUIfQMxcCnuDC47gOeIbSWhS7V8SZguDPNcyJZWu
nYW1YCe5Z/qv6Rofye24smRXD8IMGivEPNempOa2WjCxk8Rmo6SVE5TjiZWt0Y1V
3m+ORb8xxXGO8UcRfcmqVXENLGsPV7SYE4crv6voxbmSec2JxSdpJj5Ck8fvqFOS
cWpbLqfwJSRBbj98KQQCSPwAWYf9Rr6V6dyvFx9RobDySWYHyyvKUN48uivgSYdh
B1Wz5hrnq/kklOanARZWyhKsG3fmuoV/xMHtmR32mFT5F/EksLKSzi6cw9lRTs2f
6advnLZLksbqXyB0FzhrtzDvh5gMtPMo1fVEoRUY0u6yPyGxTW5QIDWnPyezimTy
ijmXrJF7A3gi/kCrPVanqmTP1PmLqJYtgl9GdbBzhgXRl/zEj18fwTTcmeY9MfgR
TigBdoGLYPQhk1oOpemofsYmFHz5aB2R5ay1omVhGlHIdiKDHS+C6tlhf+bsMqFf
cQ6+DV2X5h2/iYV5a7Xkdne65C+S/80OouHSJBKtJ0Tt3wMDQZen/aWSGtGUewaz
K3Vv2UtAWVhScZVzg+/csA2vipZTNghoBeLXwCnmeMY8kCPXacmzIVh9MZcFp/4y
fyhGV5pj4oezwbGHv52M30G4hrs+B3dxghEWGruQlW44eqXozWchfrPUMnj2bP/b
f+ie8bwSZriSxJsEt0wEXWxaaThx9BbooiizXNxFaQxevj3Zd1Z/Da1o3IIWRbvK
lSTldrySdMQnI2dj/Aoc27NFphNAR2Utm6nNqLvnkIhztbPZRozAXRJcqaJxHINC
HH494di2o2TVO+7YQBPJ61yfD6Azpp0hZhN/5uqp3UqyLB82tiZ8c6vZ9pwNq+vu
pbGIJ4aQ7eT1bBsPRQohkGHDPpEEK8pPnFxxXd8/3BlPTpYJATbmiKonq+Ya1y7B
GwarH0vqykvCrjSE0/6zgjVyj+R2Zl43cBvpTGtZgsGAEl4oUeCdtAixbOUQkmXY
LMBHyiKG/GtEaGE0/Qju97IZzr64NXvEJ7Nz2rudGj158hHbkApPkVAIAvpoL8vF
iLOkFc2noZAFrkDvkVOGM3Ha2vczChInzm1/kjXXaeObWms7tTfYalfntYTbKYcw
dVrLTeYVZhULNu2l86TZLfTAJzO4kW7JzRtVXQcFyMdut3VuFdHAPdYcMBnxsx9q
SvT1zpA+hLw9j7g6uOAg7HFyag08HLJ/jU2rZzfpCaPEzI1bjo4VLAfyloP4Fhpk
FYvL6O//LucdhOCyGicBJ723wzTqyhfZD8f3ws+1ohwFqlcd0S8y8wnDj1/gnCoy
VhVWnZcN8/GwQ736TwuoQvAW0uUP1KQ2+d4QwtT2a7g/PuvZS57EWKEEZ7On7uKv
62cbkTuRr62wnp9V90e6+CP/TxrIVNo+NYSxpQLcw1xGtIvwnqOFGjMwDvSCFEiL
4+YjOcNEhb6U7Nf0b38w/EmRR/fRZCsA8hMjKQ99B9S1cdWfw24OjuRs1llPrLjv
Mclnly/GD4APmliV04h9R/6d+qXUiqAIniLFPiF20Xf9dtfAXNxC6JS2LyvDGJuS
tNUVCtKpsfmtyU0fN6+fip/7ayoSNfOSgum5d1yDjB1RXtMnNdAEjmsi7p7sbFDU
zVWYcTes4biJmq3Lpg5vnrE3nRlpC6iOBaYWpS3HbNc1RVAgIwNQ8oNAKzCF0JYs
6ByiVA4MRaMzRpUqRQZ6SYccWsC8JGweS8+BVniVRY452titnWVjJFB51mis0Uty
VcXXAC4o3YWhWYDwq7HWbis+3vGfRXBxFFRYOz+yozbgWF/8iSU8iGD0arQHPved
72K7k/NSNDolXluyHdCJ8N08CWrXLKgBV2CupF44wTRz4e+DMzaWz4i5djURo9OS
Mrd9L71E6+6fb4OrF2XK+B5d+iqii45+LENiOz8WfebZDpQLfRtMOLfRYsbfUDzs
14N3eo36gczoHAmAPHQTNT4DmdpsPm/3+UqTnaJ+cacOw2hDOUZKfC60ABo4Sau1
WxmQ3FdouvQUDChbtoKBFISpjxZdrz3Y5+43Y2hmTN/ZNaYbJcgH42z8zIytOoqO
XE5UbZRuDGoUeOjqHVeD5yIbCekq/ra76FfZssSfkRrEaGXDTi9ARtBVYJU2ygTy
iI9DtRydXZhdE21iOBTquyfL1Yv4GJXRljJZi8Hg1dy1/HZJoQE0Ie+Pqm6bFtoO
beGgN1fdh3eIbXtPbHccg2J4/L+85+jJzOQv32dOe9B0SdhDwTC0xKwH16z7qUrB
DCpBZbZ5IXHodvhTXokxmQSUSqEWAr+y/nDlSJfBHGWEYkXCp0XCm21ky/8S13u9
9o2DU2Vkp7RjrHyl2ckY5FTZeeowAocTpJlp0t4WuFfYSxqB/3LCbTJMWbFfPDto
TE3yyELYHZXBAnqJTEAmP/9qB3ZO1uMOYzBKXYRZ2hK3u80G8qRXWO6TkRPTipzz
QzaW65QP63V3PrwjLZV1Fh+Bh4BK3oggRd1uOoPuXMqyPhN8BRF8q6zikA87Z5sj
+eC72wJ+XYmgj1gAYA2Zg3b/l0Gib/rsHZI+KAbeC3+Z4IsiA5EsrgXqc8hO40gh
xwpa8j9nmekc5/klj3mv2NeQfpXutAuaPEVH9kBFQ1ep1HNn90x/dxn6Bg40Tjvu
DnOvMgA8xvZWpnftHs8ofiq2Ide3ve/WRVMEdqp0Fr/M18xmBWzcsyvPRNTcQp2n
U7+thls1aqZaoiScS0CUuDCAlg6GTaN1dkOZMkxXXRyNC/LY4lG4Q39OV3IMDjm+
aLZvxGL9QWZUK5cFqfq/5INLlhNwKTVNmx4bOzTs+IsPzGwN0AvcEfpU0ggAuG3y
EakUd31BTmskSN6sXv4WORuF4RmUzfsnMe/mis6T6z0CDSsAuRjufXRhxaqETJZM
neKqTRggflwXq7ls2XYZlmqmzRof4dlfE6Tw8DcjSyOwz6uXkW5XFqapBVMKkiI4
8SuH3qdTa4EwNaEPdcg7/J+R/W7mEv2aRwesNQ+AjNJj6ZykW0Wi0M0KARqTFiTA
uVrphrvLcnyv38IRhjQq7WjwyrYQZ/9cLdNhMOeNnKqcLa0gJTfPO4DMLRGdF1Xu
JHUdq/a9Sm/zp/EQvy8H0ORXzHjvVXPmB+gRBLkfh3sPCztYHDcheNgLl75MnPeq
y1rVQa1x6QwJcKkRgmQnnSAJaUkVRYvJlPKxXQzJ6aSGjcbP1+v2GfcNIk0sHJ06
UQljHgKTFqRbs/GaVFoJbD9lv7auRL1dinHabzaiyLWdkzffdJHSipBkVjA2GJHb
oqJ0ZSPPRq17a1YEAtc4jjhRWKsX26IqTuVd6Vdgk9V6JMUO3mLUGTI81ahisIV2
25MGTbfvpiV+cdRqyuPfTE2xZNK87r3g1Hwn4zBEu3OckW+Jgv7rmY+rhh+AvYNe
2C2+EHX5oko4OPAiX0d8Ijx3Qm/fzyRxWsmQeyyBXQ1w3hplx1oj2+y0SPBFZY/7
ApMYSvyV9ljoWG9949Hy/AcBl4d6vEY8o++AUZptm5eC8Oflck2FD9hcdrNA6Ctq
pXD8BvU1j2+a2Y+xwQ5vocyUeR8n58c8HMC3a56txpe/HyBQlcgE2CSNxN4zTcoW
Xj0xdMCA/+7ySzecSusUdOYikHQ6UIZqF+TvKlWk5ycGoazOL/0vYZra/tnMif1R
Kkx0cKylhMEhUktmvINtTcOBTDygylIWmm2anjDNTJtHHXP53JLc/0tSCpTVN/NM
U81nSFWQMROVXjSAWGEAi6hzK5GBM6w1o0jsG0ERNOZkv29u1+8/o0AqhvNnwj6t
VWEfn+e3niW/uaVqA2GkmG+45oh/2HBHIJhZO8FMRtIjVUtO1+prJmHW2c5NkBd2
skF1oWwMOsPYwctX9zbufezDSbPx1TNEGZJ1FkF/W59z/vwOiqINJsbTxxG1WMrN
dhzYoZPXJceR5JbDCQjuO/srgGuqvrZwMnlCKWd72AX7n1aCiwXLEkb7du/RIH0x
C4iIPRGRcyF+7BpgTv3j6+fGgd0PjWANwlbQ4OzdzqnQKCtDskvV1SWMM4rwygvH
KseBTtRauNaXL8PhqFE/oMdZbrRWffVQ5RKy+AF+yNF2D7zF8XgY3TY4sDgomr/p
HzZLgHC+JNAqvX70QkBtfpAmHUYS146vLwQQ0WoFMFxrshaXLZi9bV4h0Uv1oB++
H9c+zoHvGDyMPpT+DcjfYyl3thJ5wy2h3N1dRF2fGmfUVDQEwp9V0df7yR2o/ZcK
Wt257qlfT37mIRA1m3WqSKM6Q4xZjE+q5EXWJ5EAxT402NrF1fqnPSoShEx+SVvp
tiOzPyA0Xl5+aUrAwb1dKlHO9Bs1NLFZn5QU2X+9sBZPUqPx3l1uB9YljgzRTrJ5
0EwB6HwK0Ei3Ik9vA3PVu97URZ2LpKBme5gZuxmWx+laDo9/OXK9OSnfs/xNaKLu
u4L64dwINdtE8obNj4B8AizDaZhOmdPOunJ1XuzH6KRpiLhzgAKuOFyoxxgTHwWH
nX+JeqHi9XNkPh6eXqcBPp1lnzN5d6qbsTdiHU+ko61FYsBSBoW4UwQvIVi2Lvya
V8udFpwvkH8vUY0COKNsWfb3l5pPSNrQfkAxDik3WKriOYGZhk8wtXgFxAd1+kJU
VhKFS9O+1qs7vauAYU1Zb0STD9R+XpjNam73ZmO0zH9QOpZ3W/s5TIc8dxTlv/7b
J7CNVgVDLvxGCzgvJwUtvxfizzWbbXZcHdYTqV+zz3MrEljv6GdH8XvtD5NHDzlp
7xyj7CP74DC1sG0j5Op8IhnOx8mmTW7imPRyuJVcz/2PWkMTG5caADveHcvkax5q
v56vbSgEQAr1nRH2E8zyDs5VurJRr2O4J1VEdKfjH1XeJbWwHz9MqGLLen9BHXL2
ObStf7wtnJPnrTf2mzV0m/scYpbhNQUcJalvYmLEq++O/SOrKJ2vwXrRZhIgNrxA
hBIbIkpjzEJ9NhNQrJ/q/sgRkSR6bYtVTvr2VVBH2Nf+jjmsHtVywsFrGQlHtPYw
1tJelGIgigWObFxa4/cMUaSdDgm/+PhAd0bbfgqha9IFA4SL4WYj298i36t3mwxk
ih+Gxpc+2BhpEKAa5l4Xdy9h9ozXaWm1DfJ6Kgau57xh28cmN3yOWkr+NA5BqFkx
FFDBSSPSnMNVXF1R6SG3pXDOGHvvifjgXwnAaxBl+wc4DGM0yoYoFLE0Iwclud9p
jK9fVVhKWJJwHo3fqj3yYy61RTomHpAcAaWrLrbLvC/REeYgNJmnptX8guuV2AWH
RoyHdBCW6sUtnS7xmA2cMLDEpmD/vEwYJ76AsL4RIZfqf0dE0lPb92G5KuIQQ2iC
4avR47NqKSezRq9nm/+aFJT6G+jKyl4BLB64IaSs5t2X4fCe2476DMusL0f0yiqz
/bNJbc4bsWjEYbLeGJgNwtYbtwSCItswNt1EauGZ6tOWrbSlI5yYHT4shdjgVLgr
3bVzVqhwJ/KRquLy7V0C5PywhkAm8N180OYK8slVrFNnqMGLeAQsDL7Nry0mSvDx
SXhyb2rQNGrhfilmRsmv3nTBWYtW+j62ak6dGXP7yUYylzN8guYNBp1BpylHTDZM
gdhSGwpTkmfLBpO6jcy1MS7mktFve6Y4x3Us0AcHGoO3ein0vTDvxiyn3JQBsVIR
KEUdle+1722MHfkhdRIq9QZKljFweq6sWpJPMlyG1DkEfZpvIJbeeFpO3S5OIqo2
bSMtWhAHqWwpwyrbuzeBHb5ucqCdC4G/zdvlD57oWSILWAsQa8ki6XCnVq6nmxAF
9kAir1df567YbY0SofotE/oU4Fv1dj/AVSq49MLSlq6HutBt4O9HMO02t0ldNPnl
QltBirq8e+FzNbsD42ua3fzp05HURTdbcs2WEMttPBG3h0ETArujq4B3HCA/71oZ
yTJo81Z0h3ujFYr3fcx/cNtq7XWBVj9VXCObsa0wZhZtNZcze9A9ZTMPq/84Zr7w
4Y3NsrK4vSSCRXF7nk9Ar2+r/eIK3A7stKx9ft8/TI0li3wqi2VMMfxEBBbw7lxN
PWOBniut8RO0uvqSarDbMMekk9Ahdg1DkF5qHoMdM6uoi4AO5pYY8buTPG5hu3Uu
8TODnlRPswXK2+dTdVtZn74GmqhDOEKawGTkPTD53Y8VapnpMQa4BbddLqNP+HEc
4MX2tbRWFccpzDEiuLvkybzAhtwWx6Y7bM0/bVPWWCRr8zV71Y58jw7JzzaUFOmu
/tKM0oBMxvE792dOjveY7yl/F+gRmHs4em0wJ1rimOCjYgrFD0pXS8sXVy8UGnEI
7RghpogAD6q8rT5tTuqG4BdTVuKnfjrGxcb/I+vHKipzskcCCDCwsfBDyeBy083z
ODfNf3wrAy5GxVYNVz2k4OG3/8Pb8qzI4U7QvgI5AnnnH+NuVQQoF4vPyIv3xGK+
IWg7lWTgYhZH0WBvF7C8hTWTauXY+BXcGOnEWfbNMSJdkNLK5bikMrum7UoqFJuK
1zEbnp/BDc9LuXVDTvk6hjx8kbzJMvxd5BA/BKKzqjIx/+H2KegHZ/QDMZMPkefw
ulGEezxOn8kM6gT/oiQ2Ty5UzT+tR+PokzRqtg7vQW2aDN3gpwqe2v0V4Sf5km34
qNxiUec7QPM7iZh8NKSriAWeNu2+JGhtWyDPmMEcBnDF/ek02uiwocgi1LO9PFS7
36tzfzm9O+GVIkCxjA59f8Cnf41689WWdMrnu7r/TTgRI1XRPmLkrPoSZOKpUgjg
S1PdbOYmyYVqyoeFMnsvq964M7u1dnihfVuQrhTbhRoTbS4VsRcN+oF2PN94Y4Fm
0KFjtFSWq44BpcVBJIhVbQksAi81qBtJ77tqzDvDtjJebxY9jBn9dX3DP5ZrII5E
wyv3hSD7HnjjySrDDU9Ht5zG5UxDArTc+4/Um74PmdDXUUQX7mmayQAfUko2M4re
edevR90RjDf9UdSxZROJg1iwDyH4c5MuVnfGqNosrBRUmnVTsqzkK+twP/RV94NH
67Vgci8zRYAvCHpX4oSkUDyZmoNUiJmlzzoIgEDqW6zDJ8efOpzYyvjevEmrvqCE
nOwYx95kUxoG9dpnBZ45SQEiT979WIk5GORZzOK59Ws8/dJF8hmVeIz0Zz5aUpld
/MDy9MzBwzZdBwJRZAgi0zv3SF1vXYW2HZy5EInznGUQjN4GtMKsnXh2uiJABLIS
HmfDUCG0T4rgxojvBb6ABz9RRNNKhTFYYrNAdioKOTjFbnpa8JEpyBtqHpqc9uii
wXn1IlEr9FuqvMfpo8LS1opYZ7Hi7UnXkH2jrtJp6bj0JQYntUF8mGaHpsW9l31i
3OtrQeS2pozWHzUJ0CJKDJX64InkHGWrWARdp0p/O148U99Gy3JG4ktIkPs+sI+6
H/dIQ1Enht6OcxrAMlmvM8j2kQOiFphuxS+/gX+upwyw3a+id+yuIPOiCqEPoddU
IpZ2HFdz0NMCEPWFIgVfWhsQjI4MOeiPSlZaiI/tEAgvqhAhqLmljxz9uSWonxfe
QAqynPatmn2NlJlyK8VbBwtniyQDfP9kCBguHpLqd3oJszeFAeVJ+IF+8KOYeixb
NihfgY3ddvvHf+s5u85fedPsztfKifHCR8cC5f7PiUi0gVkQNbNh1DoXaeQNQoau
KAYO1FN81nfY9eFF54x95KD1P8y6GSdQ+vv5WKvOkGJ2h0cO0YSI5D0h4tYuU/nJ
VN1VtQApJOmpuZ3qJfqoqF2l2ii3mJD+7uIXhclsvlAh5FLiy6FLC37f4BhXqbNU
/Agc6opHXYzVLSvaGKfQvTvQdNjdxA9oUDGzp7AM28YETv/+Ber0K6++5Tk5WaZK
SpLS9BrRPMJ8qXT2yLjIQ8Ci+fcvyDg0XzapCdaidyVzoNcFh0L30ZedXhUbaNeB
avYcJj/s817nvpTstxilhYGPpzKuA8QFzXOpPk8tJJRMCRF5mBmXPgwS4AAnpSIx
FCUgGGl3TpG557tPXtL68crsvedkbe47oSMMcg2KDPN/bG3cSrpMzu1mprJQD19P
hZgvd0zmS97sD+YGmYF26mYagbk/frnoYIvn/qiuVonXISDtde1zc2wJflXQ0qFF
9LMNnGSx4HYfW+CmHffnl1b82Nu8lto9SbAQ/O5QsLp/XJ3lChfXPuVCa3Crt4Ts
nt7Zcts6LL+/iHeNi6A+sWUO671lfSHU5QbKLRdg5Pgdeg48LIqC91Z1XghPU0qN
QWq/0ADj84YNp7TLax9zvhTvu1Oc+/l3QDXZVu29pFGoi3wTkhk8TlB241vF5ToJ
IA4tVueWuoRRn4gGGxij0BqE0g36NIYaay7QZRtq1azu6h389+eLwOhaT33LnJPw
SQfRR1+Tne8zSfHkpzZ0L3vDaoXC1ZD/NI4PLv5ExFaRdfaayp3evT0mHgqDT2nu
bnT+ivIpjPs/o8o8XI9xfx2ve9HPAbMaFjoWEMJFEWR90zKeK3yGoiPZDe3lFIeU
uT5K+m7WnHCXXP2+drrDYBbd5wsOu5sgMTgBu/1Bh7TspjrHwq2sevJnKGL+cukb
8+UvJCgMUvmYEEbYdGiZ6+HaJbMIOA9vV4geFPGDAuiZOgIp0atalJPFKg5WbUj8
IgRy6jWBk7OlrkTXDe+VcU0cKIgF3A5F+jNJjDCXScmP9V46MHpr+sTW7msMT/bU
g6TRYqnMeDPYHKUivTe9tFGGujzmY90P7jAfqYZNSaul1U0XmFaPzOt8dlbQAf6n
jeDVJ2ErFGcCr34dArpwTMfaTtcBshYnb5XHB06We6UMUKgRB8BDqi1hp1XBm5Vx
gSgZgC29CW9Ti5o04mAGVq0Mvawta1uAIfzy3paiv5l5f85/glZNZtXJF5PeQDSR
psZjfWU7hdKztXaFF+HwQqdS8FV7LqnF56rrpNZG07n+erlQUU6AyRYwxY3YNOo0
WRE06YDwDiaz0keXb3mvOFUtvniCPfWX+LykVtVjP96D/d1RG6lFYWyTn6nVHI5b
vyHw8cTUTkANtVi6OAxwlGscJXOvLVcwVpb07W21vhA1pgXQc56otp9rbTVwQ24Q
10tiBjNEskj+QxsH7olXC5R0ch6+RTG2RhKjfoxcjTMsfM8gKNV7vZN3xEXozjjD
xPygiFmmrxQSZD2wPrlaOSx1sneexkPQtUAU7vP5bzc/UBL3sXBzXzXvj3Z1Zn0i
O8SMMFnNHzPAqzYfRnSu0KBfe2VyBBFWjP660O7YmdSuOMrzatwd+pvUS2m4CFMC
y+U+XbKwFfT3i7XRGBcvbj2SCG3m5kwVpZeUSpTGaEkFaXvuW0jbe5fU/IGil2B/
ViPARbJATaR1NMGPb6H45CZnz19lFZ1N1ZVLM+8uj8TRJwNQuPe3ny8xQvGXdNIH
ghseMAQ+SFHEaKz/kuJTlmlQ+We8tck6CSUxlULJ+f8D/XLiZMS8PUASe5L2+O4r
faq/15m9pOGQVILjRHuqr5cmZSq3yzFOPh7exkCG38WUh1JoT/0i328UUSBhvwcS
d+9t0jg7tEnZ1M+iEpPCf7UL3r23nwYVPdZVMVzh3/SJ0ygiXKUMzeIicbrKMveX
2rGPV8btuodggjtWZQZro8CXa29XsOS15zYvcVKleToh+3hpXTCMzJfSYHWYzdaP
Fq94xhWL6hONPMmmrnf4RGTtluq9233bi1f+/HEtF/xGAcDT1w3TPj7iXAO4KtVB
ISjASzauUooSpGmT3jgZhH9ySAHSFlRf2Ar9BWYHJyS3FNIwGAI+YLYU+otlGonn
3GrlJu9EaK6qtYKwIi9LcQ2cmbEYrxTuYnoZc7wnUiavdlS0Z1qJCLKmvt3nXAMI
/RQ7jQLLuE1SYlWLrny4XId7BtRhVBQiAbFsTDgCuqwTVciHhfnhldx/LkobZmPp
zc5bNN4SjBudjBzIA7XieX/mJ03GIvkxO3wz1MHChTxnSvjB7j97AkmZy/Wj6zPK
cSwuPC/vxbziZFaHMKwgCPTc5j+/Wm9Er0c8WIkYAUudvkXFR3JkPhRhu/c0KGuK
Akf3qT3GwiIGjhRg8w+GIQatpuhXJgni3+K3z0Q9G1pr9tSwEoT09TfqfQ0SHgz9
Dhe/Eyv3XmNou3rqDzZCdgxUR/+ebr5DwF8vj7TrUZZCFP0F3OUBOHBMI1Mbq83q
PAd03Hk7UW7vUpNFNr3ikrErHKnklEdSyzGcRT6j/mNnjty35Q87RGZOK0ckp3zH
ml2QtMQvU1o4E6ZdUq9raokN+rNUPLJi5vIBVYfe+H/Y7Hm/vyPRsL3SjrTSo4Le
fGN7FdLeUSgp5o7B5WjSpsI+/iHC57bZayWiuAry3S3EogD8d+Gm15CA/2hfNuKT
cbMq4wzyshjwTQ/dltqaLxixUw4/zV4eMjnult8wLY0n1mMg0EChegnJ5DpQEi3x
0DZRdmCopj0c3h4DorEdNCDYBfIlRFvFDr/WKOpeXUopJKE22SVfLUseRZD5Ynxr
9nEq32Pss4e1EJ6gbK0pPo6hLu8qtr7SFcFYiKn7XfG2v3NvsxB1rcqtgRACw6mF
vReu7jjCaFJ9f4HnJB2CBgjcDv6JbWOHTI/xVNXd0Nhx6OqaHqkfvBil27sLhw1q
5MKLqDnZc3U2ENrzfysfghYAtB92kUcSyJqTB+nA9kEpdZ4JNEl9Co2r1glbMvKP
2k316thKtCmWs+zsM68VV4YycPK827J1C3ppWpa3GP/J6gSHiqlAT6/nD+DxG7Kf
EM76x/KVlV16cgIyr8iu2kSTl8aMcqfYRabtUXkKj5Abk27N763FDHg0IooQeQRV
CK8b4O+BlP+J2IbydsSL3zkJvud58MTywzaSOPzjkk/kDPvj4HXKs1xEDLnr9p1V
dzqir2B4LmFhkytjg06Hq4wPSRXH9tlKSNnJ9alBcL6EjA6TR+8SKae3negfXNPM
/BJdkYI7SBHlh+Kz9Lqvc83FPpPKhiFL6BZmA8ksA1xMq6Sy9hNctBmdbMutUTVn
t+8XGrdySqXewHbnHPbiBzamMkpEV4jvA0T1U/PNBAQpmGzEpqU7lB03FoHuoHJz
kXT7u4Oo9B1/7BejCMg2aQAcs9NeBGRvY34AUBv7Pp3U1pi/38psJUn74KUGkNNe
PMKX4cIA7KKr/2oy2rXvJC98U4Wz6/3iRNm00HO97dQmNgRVwFDYpD0iWCWRgRju
NMWDtVoiL9Fm8LIUuJB2ZJ2i0k0PkXZ0PFE/ewrIUMoSjUVDxl7Rsuw7r3XmR/7C
FwUBlSRDYPC6MwD8CZZlFkKLDZl3Vq8ah6KE9baTP5QeCVzg1pkgx5ZjMOjQ/CLk
50/XY7YMI5nf1MYTUs+Q0QF2HziLOB1hBQYeywqyYGJmXYR3N0jQGWSHn1NmLk22
nH8SBVjeWV0BI+WOhNOUa8LlxRkN9iWsJ0B30YbbqZvaIR5reFXaVfl2/3vg5mKK
0R4/2sKZ+sjI8ddPK6ANXPj/X1Q8GdsP2ShJWTKirIplrVuFhpgPrWuwOh640lMw
cv1m17NNXIKCZiviQYAGEd6X08EsywN/h9SlP3LrMy8yzWMoFOqjrsMglFZOkx12
YLs6D9PCZLn8YtBOoq2miM2+9euHzVLa1EWV0YL5KD5oTAApH/L7GTaznLg3zL2a
GqODPSfkEP6+zLNZdutf2cbO1ewe5Slf+Eb2jhWtB+S0mxwZEls5O7blaymSG9TM
CQHBvYkIXb6BIKNYs5fNErLa16jRVg8Q46eCMVv+O92OgKTB8wC+2iuJHny2Np/9
HMUBzdiFtNPbglmgtqXcolVw4ipW2kzSNxV1zBhpNeY4M/zjEfXG5u180417QOdj
8T1qpb+g037Sj/HMq6bus0i0fwZvTMYT0LvmdrLVBXMDKo4+x1AePJvF+OlTXiY9
W68tUlyskhVCnVTxc5nfMXVGmYPtmDFe/6jWBZU4nzyGxiAK8bVVJZvCbb0zu7yk
/qtAefxMvoidq8mhHsGw2NufmD6GUVMwBfoOszK4oN6CZJxSAafzr7yVLy25NBdj
xumRsbCF5X4zOYf4tKIW/dlyk4NaPJI0SOeshtM3Q6wBESfe5gjPsK5jaXT9OqsC
pyjL8IHKlL6zDaKYZlPe56xr1YLzzdHJyTOsACkDS5SIvUPR+DdLNtUHDcE5jPYb
WG1+PdN0xwh+0RrDBWYj9/Gzwmdj/7Iz67fe1EAAD7oki6M33VY8UyQ0bQqlFS46
ghpbdRLEkaxWm1fY3mQZ1TASukNH1T5qIiG+VFBHkeu4WiYgjlfqTJj1Sobyo7Ki
JQnghU7/6Hj6T3X/ajR+1L+QniOF5p2h7GIehkHqjRl1HwKA72bP7hJwT34p9mga
fleuWKLo03COYJiPg+0j7i6r7IApNYlzmjqe0x39ilJGZl5+ySGquCjtlfvWQng9
KIN/J1cVBlZ0dwr4lJ1mBxBdavpopJVkt5AfrPOeQATs7NnuWv+08nOVF2H/KBk2
CDNZE9J7LO9aDPYzbLG/92idZ3BQj8ApcfcoHLSTc+M7wqIFz41Uq9ixb3RsN/y9
EuNgRMH9DVCQ/9m21gsQD6orQxcagibSudRnxJ/Ucrd92ZLw48kLoeDUmdHGax54
aD4tHNL+WE/oR67yznDDI4+HBGeB9dgecRq3LOnHwZK0Of+reU+/dVz7vF993PDX
zW24chytbOMP5xgB093mRBnyAel9JYgQ8L8Bt+D+ofSClazjpepSc0YBYF+HtNe0
DaKwExIINY00Dw2FxSMDIOc5D2tV9QKBVQYXFW0Mr/oYLvNssrK6bR7edY+wvIhT
cif2Z79OEidaM7OxeUIwMVCPcXLNuiFLTTK+NRUlNoUCaiQAkB8cnwAm5NQ73G6X
a3mCvaF+crH5fC4opn+W6MaWjt7uR0sEPl1Wa4PaX7SCbud7c4wGu0RgeSi2SBqu
Hy3xRxukBF6QNIbp91F+tc3XOQN4QpPAIQRBX68YOKGSOn+kfo4f4uGNQvOo9wYt
z5dDyGVrWVfj5WkvMFtLBiJXQmPE0pvPwhLGJmh7N/2VKsMAKyQbPp7pNsLQvwlC
IN1KRmQUCVYy9SV/NHAptIYnHER+7HefWzhuWZOVKHGp2j/UKmJ3vSIdMC9sJvb3
bc6t6+9HMgdRk0igt0h8AvgFmVf1qXHn3cj9udLM9gaxzF77hQ50Oscdjbixj7qt
ISIUdIFuzc/PBQwiRwBjZbKGCQ+XTALDOvQjfAif6lcZnQ1d3jIKmoDL4fmJT0d5
ACzLiU+7wJ6Qwg51Srx3H8Jy3nS5rWPodgi2EdWMXc3Ab2krO7G3LUv6jKeUa4GL
z0IRsfWF1yNvEbE82zOeDnrVKpldUnd/SFDoejT02UBoqrtsT3ROl9rMPIBU/yWq
OKgfSYXb8UeoGvknn71p0YWx7bqMubnnkJbbTyxbkDns2ER8PpKDBnQ315ogr7dz
lfqz7vfV3eGOngLVbyrIfHzyV6Sm9Es4OmzMaaMCXAyosdHUKEJ32pfTHsu4bsIU
iayYDpBY/H6AiHPm1W4b7PZFzzk5yX/auVcgIX/l75/kwU8Xd/tFR4+UABVDsBQI
DWbAuSKkac0n0Jsn6SwquHh3QbeYfXNYJiYLFbA/6c2b/mq8povTuzCc4ITYuGx9
oYn1Q4qMNZBUOK4heBPm//nfywFqcQ5BsjVNkUGFi5ntC5fYbKn/+d5CMNAV/gb1
Rq/Dn/+Hsjlg5Fv/doqNls/gPXW13sefHWvXtg3QimmKg3lCmKPvfRgZnIS2UUgb
GPGuwJs4AHhecKFY5st0zvHhuwPh0d1DieTfS4go52PVEA/tUF1tTbQCDn0SLP5z
ZPWipS0s72c0mKZuhlDc/eBLvVee07GsJf6GS5oI5asgEf975q7Cb9HBvT4OxlNi
3Mvdx4P9EFpnlOlgNcGWui+/ufeDbHojIWJVLV1H1ljQ9YKvr43q468KTvKnsJ01
9EA57QwTwTUk+SPzx9B5y/j/+0uJrSARcIcOmI82BlqwFRnV/eLvk0uToG3Cv4If
/vO+LmBgrzpci/1bLGehZEYy7VJxCw83oMwQMr9CnFm8+dlM2cCx+G8GU+bE02zt
tpJ4tZYl4H5evMvZE2qXvkozGkxZ07QgEUz1sfDXVlsuC+6EKD2oq5kGeodNjTD/
sK1Qxbz2WF5GfMTKIxigaUrGg0oVa30fuvtxaAOOM2RMclYwgdVC+utM+yaJAXyO
DZRp8VHSoV4Sj0ek+crqBTOgnJ8405kFJW3i+ldsPIFKPYyNpnY/odRY8rzc11Y8
CFXOkWkZp8PX9qHeuH3iUnoOiAvJPKVGXXqECyp3C2N0PGAJoMIOp9FgnE/X2/5E
UFQUFpmI4cxEMTrulQ7w18NpQI6mq+4lqX4eNfHsDfbiXmCdbows3rs/Yxeb18Zt
mW49ryn2qD0Fq0ZDMoW7cmpWbpoScTp5YClL8gQHFVU3F64/XDB+cBUfchr5HImV
hlL7T5/DtDWprsE0Cj6izHPmSwPM/ueiWOH2f10UQVI9cR4Rk7kUBO78LtoHetNg
xAokrax8u+d+n0ShHzdI8SpwPdhQw8prEswPO9R+enLNl0EiAJPXN+e4kG3q0D8X
pTmQd8DCtTX0a0vyCqwpwdpCBVfwzF/K4Pn2sj1RDOqB9rr1xpSbhTn4IX0jx67h
Iw1mmQM1w6TMki/pA1lTplp0gSVlKCWLjOd6hlWCqX1WapFWCpsCx0/cZJyJb8D8
yaauNCcpJKwSNMrgbKH62HGNMjqzdM9MQ52f2zSG4196h1pFqGZGddhNH7U6izL0
/zYGap/hfO3Z57dVBzOdnOklsjOs0okJMg5CptqyTL00YFRuliJBlTgsOXIAywSs
Ek6zcCz7NaVorRRaZDysfcEAed6n5T+zKX2ESlOc7YaG8OxiwbeOeX5WiOM53Na7
JI6nWAW1JjqonEkYzM9Hp3E8wp5SqZDl09Sv7MOFmsUWfhM2iBJbvhGS2Xo/rEZP
mSxyRCbap6oSrJfTNMmyOiXvmlCpC3p2GtimtATOTbQ5cJTgoxYoR9wqD4u6iHvU
VXFw4aNCLUhhJdbA/RmMlCqGYJvFdECTnfmb8hXCCwhJJRmLvgBRp4FODyp2x0ca
qLDsTcQaNJOpGOdJCyGu2sxmPMWygNsAMyokgqPZ1i9amS0c06/BNkDajDC3JdK7
Uh2Kzmd8krkiDG8Q4Mt7CNSB2hgD+PfKBBvMYvvsvDIoZIbLcjLzCSnNTkmZEldU
UHbt7g0o3Ohjhbd3no5hO3Q+RmrUTID8p+YhePiVMpZC0Elb/9mIcSP/n/QTJcy1
nwwg02/4IKMeE/j/TqfxNf6DYGMm8LeKG139FIYz7dBwco9G94ZeBjMei3NQj6Y2
cn804viyBGgKmQckpGwHl5gUE3u5/hGaMdiCl5fg5z+6R3WkuZf2YxtWtlAWBnIT
Gl9juzMVZD2sGtin13r3Jg4j9rq6UrcbEsbMBD/OKpabCMWqry+/05U4L028al24
OOVGZNBtNhN9JnlWIsLjuyN0mmU57QHgyIguHsoirW/9ZS+mnGVQ9rSb/vT0mjdC
oO+4OPrXGiubQau7kkjM2LI8ZZToWk8mlzt3BnNhSE019CJgesLMhD1O98A0xtlm
OnoipPfrnFpA2rdJCH6duRl1mLMfQomsewALiyIMtcn1f2CdpSOxHEaYE4ZKD71O
BZ4XuN4ErJpfsA2QM9qrJ6v7X0iup174UFwbbQMoPhlEnZV6Mf3UBD/szNswwl06
qOchoSmVVFNOsxQK/LsRdDEmgnytXMmTp0yH3PDY/jxxIbNgrMuH7rM7YzWhZiSx
1lsnnCzUWna5ZQpndMIg8Kp4rqLa7qvMlgfP0d8UDoA0uAWZ1jo0hqsZnXEyZYq6
GOc79UzVArZCI/Gy3+jqAJQk7E+9VQJ5WhJr5DHqpbPkzuW6AOdG7A6L+olaK2Xj
dsG1H+TFofYHUaLoVvfsoswORfxiNNK1Fvnhh0bMm5RENNNJMm+kKc1tQOF/7edK
Cf47cr14EZMAswkxARHIXHi4dG9vHPgDcVdDadg1R4Wb8nXcTUoQ5UwBovOnxSl4
8+gE24n8Uw+O6AWVg2gcR0XB92ubgfd47q3lOA5ku/4qw42pfNqqE7VI2pYTLbLG
6f1ArUQJwug5AGneaJfHYHbeLkv8TAOsQbwRYqTmq8GqzfxAdBM8AXaXVpdBe7Xf
nFvPrcby/t1PhG83Xrw3h3byFsdmcNJtEI+2oGNJIpkKsVG0YXVnkgs27eosFFby
Whktnhb3HTWm+X1ZrZk6t4Q3Uv7W53YoV9m8w3PvjDXcVq66h7BvWRlhq/jIXhzL
gc2NT8Z+PezY6HhfH72WCywqmj152y0GPoV+qbjwz4ABA2jNkCnvC6quL1YMy2VC
+C4cm1fy1o90iSIoDqXzwn+uWxBIBZWVDbgLgW/TTPL3fA0EybQwdP5ZIRILvHHD
OBzqNFBvt+0t9gxRfO6MMkDlLYzCEok/+GaamHR0/QQIL5wUwytIz80kvqoxZZxP
QAzWZ90+NNbE48q4rYW1Fenszb6XfIUVRhlcCxR1katrALHsUyySjgM/oGRTTASA
PpcgovU5WHhu4MHG6pJOjmkwh/b14trjhbAgVWtJLzo5ZZe9W0FUH/Wq+qjoe3VS
ltbDOxBEQSyG/WdMNJPMYSyMrgT2JOvbqLDddfIOr5LsDxwLfcWx4I481CjVCijd
UKX5OJ0w5ocFl8eMINkesQ38iUnO0+SSXXxQamFwposBL00h3PoAiqZ5zzHM1whG
iStM4jZkVTRRgXaI+u1m6XOViffVjHSBEdcCJcBE4AjrGIw5rSaWiwa/VnrpTNv2
mEWKWkLYHVc0sUZESPbenJb5jk5WpJP0CDLrKMwuOESTAkggxxBFO78N6/eax58v
sp4JCOKxNC13sUsM7mo/FhwBZLDf0FyQVd0UoXeZ1D/vk4qf7Chpvr3DgwPgLzyH
EFDEe8mlHQo1vAuBPkqNm4ulDF7dWzBWumFYfkXVZSbv2aZbmFkQDH8xRZ3/hSH8
25vxTuHykwthkrX49LWjbbN0BmCS2zBFsYiFzZkj5NCV6oFZBlvLavTn91/4VWF8
PWXwt18jHQS0FRZpgF6cqvfp9IR5QxCJTbwhNF/I94T1sLQKkxPew9rbR4DXJxYB
JH7k4t+tG/wFDAim4gzBOiKavSsRw7qI6e/EgBgmpa1yxl0jqVMBvHigh000bto4
wWwesk4Zr+gUuNTx/27/6mb4zqvNaFC9A1ZITP9dFlsB9vJ7sLbsKmDPEIq72GCm
qoJ47EqYU2qQ9o9u9Nob2zyoglJQ04ZZVGIN28R7VVA0ZhQOpJz3XtEMb4Gc+AyM
rg5SgJxRETPbjFtk6+mMVRs0bpt59w1J1O9EIWXNpsgIB0hGbp69l6SIChGbFlWa
VdmKDLc+ieGQma7qhGnsOIg0kKyCpjjSE7pOXeqdHC/sqqg0ydQRpW0zuKhcjPmU
2T/d9l9ZqrBcXKi2vuwziokC4tYx7lGREGCVYNPWu7wVOFZbGgXlppGgAWcT3Ycu
XMaTo42V1L9LRotxKHHdZLpyT0h3hHB/uKLFDIf9+5RwWxOLtBpGjpylMdzZTTK1
HYcyVHcwa8e0x7s3zfKfWZeERnR87oLHaIVroM73MLUmiDJF8IwiL/87nY/JUGjd
PrrUe3Pi2JZNThRLJzHXq1ybAoFd1Ht+rBOXneG98wDiB0y0XWrt4iP+oYfez+8N
KiSm5S9A+6q1PdDfmx+dE4pzQ5JC2BwNQBrycQtK6B1vgByV39dkeS5oXJgXbBXb
94ZAEAfxzKUVjcjGIdLUu1v+PER4T3Td1JqqB+juplzGQ91hpsUs6rwfTUSOM10U
zg2Nlk6k81RnYp/7mlxKswi7yWzzO7hpCFEodLRd6ME1KuYMS0R1SCzJcd4x0kEg
onCoYzZ6p/aU+3xPDPo5zPzvyi7ksU9uKaNGVHCTW/81fAVOQeMu8q2htMW0OGoO
qVY+HkQrJJrpFGobq3G0WvH6BkWhDT8CYkIcuSBF65oHRnh3Yvf9w1R+eHfFOZ/s
ulzgbDOslhAwzT7Rfk77JxYBxOY5ki65MeomBasf0A3jU9v5SPOxOm4YpuwpISDE
JofridbTY9/ibFit4ieYnYuPQe4vy8wOYD1CV+ql0R1GSVdKg95xmVu7lqjMTm+P
Xo+dzKjbvSiMJagGHQhiYA6dawIAEvQ2S9C1M6da+X47R4eZZR0jWCevE0BgKrJN
IfALp+TGxR0n9EKypAJlcJ9vtAYTfa+ro1U7SXkdoV7AAmAddBSwvB/WjofjLdGk
sx4sT7IZtVXzxlHJO/wHEz5cun37+NBCfU/pbS6PqZ/WYrRyB01/CUlYLhxpEjFy
BnY6AifdeamIY34Q74ulJYc0ayOgC864Bnq7oowIKYSjo6Q6V2Ha1oCr0RuwLvzo
SCXeASHPRgSFyRGuEMtv/LnjgkPlxSkaVPQuHhltKh/nUJmKNaIVxrZk8+VNcvBX
FIikX3sK+ICyeFnBo+osZRjeiS7lqL90T3Qd3bBYLJEo/iqVe8ViL2IFd8IZyTfR
UJhLIBGqAnGb1rdfHJH0DrhJb9fIJNGp8XD1s9yqqcjW8OWYqUakV7dm8BhIXVlI
yNFigZaZm+vL4ntoJ5IC/6Ik1Gg2cgpW44dcv91E5YWSwbpgk1fB7bmuUsczDmhK
2mI1Ivzwvfdf0L6z4Zhkc1u0lQoG+NomYoGMBr/11ap4N7dcfn5okknkzO47M0FK
eunvBjZz46g52SjtQgy7miu9nqcw3CjuU2I35FFC1GmA4RNROJHCW0sH81yZTJjc
IURyzCaaQ6NbUeHgkM0rbXQ//G18ntPbwohJPvnIipmUovop84fzK3SAzvGtm7mB
/4oQEOqIC2oWduS91q0d/KLxQwVYThWkKYrMTTxz62CaOZXmUJWTrPAMUYVUlV6o
BtQkfjVOH/gg60YhlL2fUCe1flm6FSgelz5rmMagDpahIhsAASz3UBI/p7bVIDwn
FDimQfVnpH4MhVPKFT3WGmqpOAjafKDdrYBLmzvNg/FppgorQpQqUEDWl5M7zCU+
SgIBoNj+rlpOQ5F526tbUuQMXzHwvfrnntsa+YvQpIM8j2MtQRVZxa0L54ZUnXlZ
lw0EcjZzmUSh/hq3JDjTBMwa+oYLEO4O/5XTlcZFWp89/YbgMvZI1deXsKyksQg3
NZAXyrEoq9Ep+QYF2xkeh9xnwbuSzkzGl2FzOlKAdkvRIqWhKJtHQ08oADgSEcnF
HHxBITnniIHcMR1lLcWuhGn+vmf9KyS9Em9sFqgTMOcoJR+c3daPUbXHmn0sT+gm
zfXk5sMDUjDslta/2VVgPaRxipxsiHVpUQLztInmSnGs/l4VQ+FO9kPRTPobvX/r
eUZID70fLeZi/tIjIaekCDV7RKrubf+ANo7rUs4FozVFJHGffvWYn3MvtCVaB3Vz
2dyyT9evDaiilVynTcYsbcQ47k7eoCXXxxHz6VS95noNg4MlWssWNeWcNLxGsdiK
qrMRZsWxeJSmNdsqJmeuNIoElvYILL+CylA+6rtB6Unjp6OJH/fTf/8OaSe4ueMz
EWb8CWiGIS0tjajbjv6W/KnuessqKWg8ee6PdU43FFU0wX1qkLqQQ5RMILtro18r
yNp0SOsUUSWad6YsQMMdGb1BFf6J/OQmJ+QlQtzEVNglupHueNfN3qOyCt3lCkLR
Mc7FswhzTl7PGpBpUp+JqYPGsHfhzRaKLIVq94iTMm+6U7e/aXDF/4E9BqzMriJm
ql0Rci6dkwAWPIJAZBsN90xU3Hmrb3vrsMbeTFjpTMGib6HZa2Y/aLt6TQAcYmMg
MniGconVG2Zk0Au++GE6ClWWGjD7Z5K/dvDh0LrpMoNczT2HVh0SsijtRQTBpwCs
9wQuCL9jW2ceLhHxSapyVyZQa91EHjAgek38SjhWBSTOZKLCWq2SULVtOi4gzEzz
xh4hth4TYOhEuCxnXk/HX6Uk/pWEhzWXZ+/11vhUelbiiQfViyETKhVmeQcwI2zE
zjFG5CEPYOkYscytYwpDPPCockOB14Xu+iBOtpYnFdNZv7abOdpV3heVUmS8DXry
OTjhqg5TtuJNML+Zl9Z8ijfruO33znIbRLAUv8l5PHDIfrAkbhGhHJAgLb/YdOiU
GVafuOCg6kDgxY2gF52D60BvLvVPeRJPDimhYH/TPyNnqfQcKs7T/cuA5ru1sJY9
7dqlP2u3raqCNPJJVf5dhHj+osgHhnPvWN7tbElL83i6C3pardjky7srcVmjIbct
AoJY7GdNivm6CSSmbhhgnnfzBxwm1pcUtFCVhFv8HJ8abHwsxsvfpFkmCCacYY7e
fPBSfX0RieZ6zu5f89IgJUsFVgHUpdMIV+PJhLKLoTuw0s22vzhirMEVuCPB4D9l
umcIhIMHEyVEa8N29zDapBI6fMLyc/dp+WdHN6jLTxvcxiUpg8IVWIXo1Ofsu5YM
Qx5DpNxIfK+Z14PGwnIkjmt5b08UTle1+djqAiL043sL6VYPKWUBEGbWUj9vBrSB
i/6wfgqtvcKCaRe5yvxuue6D9EfwHl7PgreESoHVV3EnJiKCWoALTNalN/CShA8n
b8PKMTCGG4R44ipxVqKNv2bE7rdJdnRl81pfwZZRvkCaZOOYw0QQVXMzfo0VHGFQ
htjJZFdkNEBDkTPWeH/x+VPpLw9RIugZmEQO+O6fGbljbVd2nBOW/wqlYeCwQmA+
91LMPLXDvY4OUq5hW5UVZtnm8dIGkWS/MvDRWQ3U+IhiY6h304/oA4fbUY4aNBQA
Ir/FxQo5DP3nlc0vXF2aMX+TjrA4fO/wsj833KFsfbCzPNRkgjWHknXx7ocCQIr+
NJMy25Mu/L1whwZ9XQfxQYFS92k2zfBTRZn0MwH5s4mX7NBeh/IWEJ9W7+B+dtUc
P/+YAD/npjIIYNykGLijSJ3pdMxrHE/M9lI8s/yvBaok3fT05MJGrtKezMrF+THs
3lRNYOlnmJsEzl5js50Ao9wgmddJa9J8mPZRskx6lp91eBYg9674aE5qV+e21sv6
U8Ir/BvpgXPDj0LaZDF9MRVyzLY+LPXEc0BK8pET7R8+yi6+uo/kfl/Bic2FwSTu
rfw+JVfXAKfM5J5PMPYrsxVIMaufgEmmEt1xS2nqQypgg6JutTWKJRBuSCM9GiND
3r1lI9h3RBJt1epdFxanqvTiMEkviuiIGpm40SLbbi8h6zmdCIQjruzdjA2ZbqoU
jNhtyHzeN/HGGCgm3y6WfW6GoVbM7h1/Dc9OCHKHP0v9m6NHZzwYK+J5LIDd3ZyJ
TeucOlLaH06EttnlEsBJnSCiRgHLCD0JkiZCQag/5Xci284h0GgYYh6yKQBKAMrq
JdRV+BrL1nPCGdjGmkYilJhsgVmE/rhu89UO94QNFWe4WNRsE7u8Y16Pd9AFM/dG
RDvaY5pQET6BXTI1fBMnB5AdBEiJLVyN/hLl+VRmmIJnHYUZnB9Iz25twgbw5EZG
bJsrjRcVmx7abDTN3bawP9ICqKb46NTxWT4pRGJIxpXOhBae+kdSLfE7qXGSgDdQ
Q7DluFs3dK+XETqZhDP0TJSkmbQ8GF0ov68pERSwaHrQahtD/MAvTU2puQNhSVAZ
QBIMWIuTI6KTcMSudD/bXzxnbyxZFlFmKkoGXZShyMluQuLww4XCTsX0VYoxsTre
GKdtYUvGjpYDAGWucaBXOhDvMYf5ReolFMpcFf47HWNDQTX1ceF7uaVr01WOmC/4
3UX3iIO0E+M2dVJ+1mJXOfUhRFLFwpETggeXLAdHxSPYor82NOX2JYzQstaNAz/G
kW/Y82ToMDfRmwQY+g8MopDjTMRIqSWI2mqTo99JRqLn7UQgfoPvOrBkG4v3Hfv4
CTtGCyrnF99e+Jq6FCl9xCygRSIxIc6FomBoUL6wFTgnGF9OsTahCi0zoMPYVgUs
xLqufHGBB98zuy0Um5iC8oxEPlyyAAelNBwilEx6bcpA0Mfp7+5X3Vb7sl6bvEvf
hzxLT0dx6F1S+joQJK0B9geINgiz0T/Li1+ZRTRSXYRr2VfcC6QY08p7ZeoHESPr
aLlBeiggdIhOmSBQ8xPb8LVkPalM2T9a2LPrUZkC9NReJ2kirDm/8Vw0RugeWUMQ
Tg/SMt4eS8ycuGArigCj/hLIaJuvpu5kDUJJbo3+SE4ob77dvNsi15uos+nLHJLD
6bz+TTRlO7w6AGJSqMn+KXMy4RJNTrP93Vr3/9jzAYeFQIHgXzyNeK13f3leweDP
ITDol4vtwjPhZ5ysWON4QApYYJplqQOKry50DTvGaX7iwbeIo/lUNWhdPIE5gbOx
4ILynnkPvc+4wUIjDJRMmSpmL5c6jSE/H1F0APMHB+RB3Rkb4zoeOK4ch8P8lV87
OMBLxWf/WcbuJ2egNBBNjtMYSpaQzY0awq8/jQUwXbz2R2eCaPbs/JTjBwu24Xgs
66CXPWil3C78wzVkeCAs/0W8zignT7D6Fr0ntKwXy1SyZ4A6dHhoFdOQaGXFTF2s
TDQctC0swc91TKqKlhAruidFNOm1h/XUnbOHvIGDnJjKkGTqgsuyIhY+jRSAN3Cz
HD5L40A1uWtEzixvwJQoaZa3yG37yjFCg9kso6CZKixfP8FNar2usn0Y+2izUQP2
trN2h5rAy4kHRKCZ3HTBNuq62HMFYDOkiXkncoh4vWJYfvqp2JfzcAT4sW+pBSY3
xkuG6Z2hlzT7PggDQZgUG0Ua0dApo9ZFSNdo9c0l7wDfr0B5TGhtFC7Co1ZpaDU/
9EAsupOP0S9mHXC+ikrJwy7T0k/4W7Ln0qZ5bfc1Qy7U7Zq73XRD/p8GrOpWTuSf
tlkBY2dpoOzEAeHj7zcgY4wNn7HnQc/wHiLhLP/uSMecdtjj2PYNFtpmrBbi7exH
9jxyQtvBZgV9viLjutVAYJcP66b34CPgEqfRSXbKkYS1hiNNOCO4Knz1qcnWxuVa
9Rm7aL3rxBPAXI7hJPZOINmruHERYT5c6GNE8n/Qj1Zsqq2Qj0qNebTXpi0mvddq
vhi/K6jr174VJjOzS8ZK+QIJsKggQXmupVjlOtXlMB/EO440YBpGzbkFf2p2VeQH
uaEGF0VcpkKiPpbMxnv8MR/dmgtiUgiRyCftKYEbtfppN3WwRmoww+nKU531NpRR
c4uOxACYjc2c1GxY7G7vAYFZc07KxGVzx6c+UIKe4Dr1VYGm0qTDjT5HGJH92UEH
YTOqKMGV9i7WbP8EQaH1aJUS94RmCcqjd4yKGJdTH9NOmV2vpbQ3IEpnNszAkFle
0L2ioI0OhEjJ1ZRF5kM3GMtpKp/MG1Q08z8QEAH4kWpkGvAsGVcYN/0RFDs38/76
+TBF68MuWJvSMoId5mBec2rd3wlEwGTBT2ZnkStoY/oHhilrWpC9Cm9or2lSUnCi
IUAOWxMxraJYrblIg4bEwUj8zZ+nUqRoC15Cg+kv+FSVTPSoWzFonKYwIog90Uog
4yEVy7gh8EgESdkzyxvRDwUWFzcMvy377DAZumACWxl1FZaIiqk4J3MLbr1hmQbp
OOFn4CSqU5lq71JeTmjfRkbtTUDD1eGjU9EOiATgTqgsRLnVZWUNiRsr6QeRoaTC
nA1CvMiEhnRTVwwXzp14MN6LsSbjLZo6+s1JXqO4leHWa1sxmASoMIRn3pv54vHp
lpIQ4ZcTNQmDgcX9bshEWXW9QJgi9gneN41jLE+a0UR8YS1sl91sPLvlf4KMD7+7
u8qWaFaaZsp89iYb+Lq+6TfuxUweu8kPLrwNdRYJLYns5zS4/EfXIlRvkJ5fcP/4
e8k4yn457XkvT3+rikWLfqxhI/lhR+GD3tX6JW+VUfkNO2jqmjdor8T5toWzCvPw
D2YlloLhhyik4fyoM49yTPg0lWWzjXNswmxlAIvW4t/02BSKo9nns5GX8sztPoL4
7N4TJl1pvYL75SqlijKTwoa+8iSoKZBo/WfFxk/YX76L2gpvh2YVeYAgC56iw0jO
TV1gHEK4EdByDQYX7ViJtiK2SqXVrb5nyyGuF1sMnBG/Z4TB/lBWoZ+2KVkMHTuJ
nkZNIAsFF6/nVYSdU5HxDOPUFxQawlgrTTmO82sz64Xgu8YcutCyucNJveO/OnCf
FDkE30Z7jm34AwDVhXt1hU2D6dRup66cSk1cpQX5QLl6DOiNi1/WxOUzEemKTBXv
c/E0U+cD2rR3+sodhClV9GvXKIQltWwU6RY0uYf9pAjfPh5JtQgGg3DrtTLMkYP9
pf9ozb92Aq6IP4EPSYX6P7dPwXx6pB9fRzP/IOkLZfcEvTK6xh0193hV/R1yEjeg
2dIh+mVh4JxTeGuSFKcK7PwvGlKLJqCKQU5ELCS7SD7wP4d7lpKFnXtPh1WW9ust
xSzxsDu0HZ+HLoZFBWzEMlWAgIZaQThaUclJWwUpbWhXXpMY4dbJc7xNHrhpvWPq
AKwCVzG97pMeoE+Z5od31YXTuavaU2Jpaywyl8RQiN3r8HWW+0kj58b0PHFELqm9
JbaWT3MQnEExSC5FVwilZBqXPUG0EWQOHhObAhtECujlC8jkqKGTRY9kFJsGDwKL
U43Qv2K3+upNntrAvco2WXS9oMNYTdCFAiBaYy+1FlRe0zwUAWGL8UjrEX+q4oAd
WBAtPJlfm7PpCHcwbisYgeP3e5lz7mFCoO3+C8bdfTdfg9V966mX6x9SaAdblba0
rWNe4xatFOf0DadeoVieZ5FYN4oYhv/UhFF68sxCt0n1X/uk9mS1FyEWJ07v90Kp
Pc1JN1SzV6S0ai3E7g6eCZeZoKNa/J+FY9HxW1vKirMNAazxRLd2rQSAXtdUSeUi
SpWB9jffPJN4wQjAGMRoxpZt+19x/0JPRfWII91f7TnloIE6pefgUGQOjQhmGnhs
1TSYgaspg2qz35wdEpdVYdkSKFnsCoShCAymBT5KBqOqQRXuX7kLiBNB/W48ZHyU
gb4r0/t+dw/cVv+Od0DpD1ee2P6+Tcz2ldLL1qGoMxNqhDT3hB//SxTMNiGIzDsp
eqWSkxEJmuS/hoC09MXfkwwh9yUIAOm6yoSboYkgnOkIFQFKAGntJIhnmmDT7CPh
Epftl1QIMtJWHpPnTMzEkxovg5b8hxC2FTFpmqU2Mzyj/AjmPg+zNImb0/GeB6ZM
dNcRn95zEOIf6l8My7tJ8doRV5cXD49A/qBx1Q7MWBq07AqrZkRcSl+dSP1GrCJU
Zw4Ih7AhZeLC4Y2kKUwyONYdFKx1JHCKAney1gn0p4qRry/XwzJKADgyB1H+qh5V
lDF1yoRkQz9CnPfuJ98VrVT+TRfSQBu2n3/7Ii6rzwcxZpPMJS74vOXk2xS/FHDp
UmkgM0AIWaXypXWYDDkDX3yvc3aADDBDw2LgYvYwUMUxpzV5LEQaqBmnk2YNnWfl
OT+h3WjlPixsTgh1oxf3P5T36MROtfwXBciukm3e1xkr7z0uRqm73NMgiXC+LZeO
tkJgdmqEAOw4cTzMwuoy1zG8g1wyq6VBlgtnkZ5mq0gczWu8M9S13Ah7BMHmZpOL
Ijy9hxJMoiRVCennfJ2vV0YXYzKXzqnmhZbJmeVrpkV7YHpLV1mn3YGTX87ctXIT
KZrOHJUTa1c81BnLFcFojLQnWWsERHvGiDUBDM+6FK7+wOqmhNEjReQ24UQdOXag
4RqlvHKzxLwxU2oHQPasS8bG543kGx/SpxNbjtwE5Ov4O1af6OGasZvRMqhF/wPo
hmatVBjU4pvIx3BWvSh3ibcXxVy1Paed4EQnD7JhvT//QMIOm0P02BcMJ8bjoJES
vtm0H71pTiSua2I8CDOzOVNXqVZaqEfuPJXZccABo/Z6cLkSOoRomEEqzaHoKmPQ
6xSs6cxK5BqOQYOjDjitLAOR5oHRTValW2vd1zRg4Vnrh79HUX18Cp9h8EA82DEl
XzzaAp4cbscILM9zC95zRo60kBmBxtcmrVioQkYY5MUDECcayR/sg7wVhtaiFLxZ
3rBzorW4pvKODerwtLTiiWt2m7l5fiVP18ZtWlXn28dQM1Y8sWh0F186A8+gnXvj
s8zNn/xaARweyumq9omerTIOEdYgQnQz+Y4BKFegWxD2PMk2a2sgYDfjK2nKDk8d
mh0H0jxjsxBIU+lkUMrTajHNPgBBgYSURuw9++3z0VAJWnviPt3GgjlXQjvb/V96
1RLAGXC4QXcsd86Sb7hpk5+SB+0IQL/q3q4WhZdufjaQb8Zjo9wd8YyDfIjOeiMJ
9/DGY582k3EP3T7YQ9R7a6B8r+Uo6UKRrJtkVF/IKZ1iKY67sRF4szoYIDS24o8Q
HvcG3g9hJagPuDq/t0cqY2te0rRdcToScQ3s6tjMGr0PomUf1Sz0i4fe00XusP4n
JCI/b8inaPylCbflb4IGwFbgJdmMIF617nXHy7oRvPvTJhxEGbsA9TuESnD9D1ow
aK5bRhZpCT6wBIh+slKafQimFkelRf/otKyCrVMMuc1N7Nbq0SIMZqa0WfN7HSyH
YhwWKgW6g2Fd7NbcKVjAan008nBH0Hu0qWu3bRtwXvqqRavB3PbzzFfiAw7spKiL
2wbbo2j6NxWWpjd2HkxxXadXckl2my8tkqI2lftTTTFYif8ejK1WxThDobCnTD8l
zBRMp6kKYNW4gIV9ZBmzyBc2MtsiMYr0hiz1w1qD9HCwuWV5yvv0OZdjGrmo24fa
OFVhRKM9GBKAF4B37M1BH6nLTnH1qMxAHn0mfIEwfxJU/vcfOGIWVNm0RqqMf9NR
J7GD6eLk7a1d8SsfYpZ6lHTFuF6x0+e+a1M82ysFTE6NYSSjV5euo4jpvRTLgy/W
PxfaEvHzWHsiqBtG3czT3KvUocJHEMmI028i3F7ln7q/FERM9H7dnnia5C7vZilA
sBwJ1u9rM5Wp20pEkBCj6w1Js4LiHHq55yBcFdesSDm4weVOuZRKwNe+Yjz68VfH
Ijs9NTkW4WRqA7zGmNJGdzoBpvAyh61XBkttjzvgym4QfpynStExtxfwQilMc3Xg
+EduwAimgzUz+rxBoGFcJlizn8VG2Mt+iwbrQGg52atidcDIDBy/sr3ped04awBt
/ZXwYkOsKBbdzKIrMR0g/UAGUcHpGQqbCQsdQbwaI9uXenciTv/TQGQGMTfD6HSg
AvE3loqsXo5NcnRZdAq95MFFIuN6p4zKHSkP3AdUy36+xFB8z58y51QhBARLoXMd
IO7ylgjtBJs9J5737ajoMEWvgllXW6DYeM9e7lugqM8jwCN03/K6TiJG0eM0yeW0
+ucMMT04DtHruLE5lEvqBVnkFAFc1UGXCNPkwUOSgEVzJqsmQbuOyu3E9SeJbADN
wRFh27E7E7STvDTYBHheyWm0nwENlUcrKB1gdpp1wM+4qDg+ubmbWi477Mpe2eon
t3AhswolwS8xM/BrFUYLyUfbcJOD4fn9R+KJc1edk0FsnY5vD4T/YX1JjVnpjzBk
w6CvPrwhtew9ZIHS6A915Tpz973zOegFjnHhEPq6YOYae5ens3KHH/WbEsLbh68P
NFN2k6b/ZKoYfFT11DNTHQOyWaz2EzgDZ9KM42g9BKqtLigr5WFg6qk4nA1diOO0
6Ti3g9F3AaRGuWA2zatJoJ8FWeFYKLshZpBlY7V7Px1yJGMMArDm3wHt/0MKapcP
zEYH7D/F1WKX48gxb6aXyrjUqWY5CixanqPH4wd2GE1otLWbupkIwgedSNhUkhDu
im25TQkivdic6mtUBK0DMUGh5lSm3wjnM64b6Ib+7s8s8FOS3OksQzItOO/Bq4a7
idiqkl+Zn7wMt9Op4YHKeW0HOj15yWBe8B7u6lLtub+4M9Q5+KND9pYu+kPxIXML
O7mdcoF2mW7z5N7+2WMC2L6eHxpo3snuVQriy2ckm6d5SgS6YSL5sC27dVkHSloG
G7cDN50yVEY3NZw9P0nytxB5taFS90cUb3p5WaYYfRNuwAYtfBPDiwX4u0kDiUat
9CUBp7fimhqNJvUBcuGETCWR6Y4hLLS0S19972vmtoPWS7FRnYpv93nMq1EgsRgc
63aAUxfGWewFtyj0s7laexjrtsbC1z/xDxNuPhHLIAhZCVujcc/KI7BynvM3w/+G
5sDowN3dv3UnmbQ7QtpDh3S0/Mj87CBVDT9wfMDwtc3xNsExpoS2qCATUvq8lp8E
b1lHhnKtprCKs4uK7Zxu/wMus4CSKBynEFmrInpXVI0F+FH7CPUi6c4DZ8gJ0PQ5
FNwo20UWNZJ6XjFkhaOYdzG0XNt4U7hm78NnyoeAFABPmmMyVQZreGqXSpl+odB1
0ZXDQWzrk6enu/iwVHeNCIk0bse+qo3DBTt/VusKYXmpvChCv2pQyZBFGTSKpwL0
R/gIUEiIKozLSW/baPfj7uQHuWEaMOEh3LVPeu8a69q+8plG60y8TUv+FiVjRcXw
sZtPu2VsBBInz0rXQmUYMG8pmUO2c0MHKAolTtlUCqFaVzWOHlh/9l2gODiCeuze
8CYGfWBNEKJiPBtCBgJxEiqU4p+kc6RBRPFOwViLDtJobMcpH7/9m+vwmRsydPXx
Exc6MSZvEvAh3QaHEc2YVqvxlaOd4mCs7X6PJdnUMvKRnXidB1j1yMUWWjyrE7s5
Vj5cvnc8usuW6V0fU+BRBSsvoFuSXC7OyKTzFDOJi5x3ndSX3j2pDPcSzGLqyIJk
t1yvnsREsjc1yhjScfmoVIRtAMOcqVY8LFt594VWTzvjLT0Rn83tW2NHY3X+EZS1
a3YXkea4sPnmgqo9oWv+FB3e8XONKutmWs+I3fQjukxMcaHs60bsVUyE0tUm2M44
MQR2qCqx3bEn2JAOr2Az8VTuzjyMEvS+G3uFAt5JbyvUkVsb9NBiW0g+Ofr/2Ydj
75+K0GvXCuoigeR2nVWGETx11GXvS9p1HvIUKT7oSWeYaKZvhTg5Y/hgQuC+fCvk
U0bxoQfhLZ/WaNlP1uMUkujs9dSfQuKZLw1Qz7cUT3Oj/aAewK278G8VS5dB3dgU
8KB6kU7fpFVblq0OFp4a8nebkE5oaDIJn5leMWyOVrccT/Pa5TommA6ywQIczGdT
ua5zqZ6FXkgKH3KvcDJOsfV14GNiGzVIqAmL1yfqB4luRFAQk3XKrU4GLciJo18e
OiOvNI+d2wyw1H7jfSy3myAWHShEvOCDNEn+YE/NnHON5tx/pMKCuJkrKQjGfsvv
+Ewco4zb4kDy8f/bEQjcRN0AL/FX5BtZX3Crbpkrn5HgoOhPNjzEYbf05Z2/nSgg
KuujSW7ldILmmVE69Rw838q7i9LUGm88ptvEj4jsWDvSVgy7Gr3AWqWVBYY2A/pd
dl6DlLcA/Amg+c72wgbPvrn22DmscTBojkf4w4h2iMfvzKWevytG2PZoBXHR/zq8
amXL55XDnd1RVXeEYoVerTGQQKuOrR3bvdE6kIfrd/8UXwPNsNV2nR0bITfFFJNm
OzxqgqJeKi9eANOI/0jTqJiaaU4rte0YvOwpotUiTwCbNIf0VVazjklZ5Z+v2Xav
mlAeDRZb0AAwSA6dPk/oXVYhBC1Z+pbBIYoozUgI/WR33iupdnEz6+yl6+geoy3n
krfyRQ005GqeCZKkp6pFiQNyZdw7x0reKHZzwarGOWXTLfQenc5DafBr/cnBlON8
vzh7FByk+ujv3P630DUVUJVTrrosdK4fIx2x8bz5a6r7DMVH9xhmEYr4LmXT2EIU
favG74T+1jpZXhkHe6Nty5fX0nf+jPh1mFWyPmXXxVE19zipc7IN7s5okZpvL1ap
kZ46AFnQHG7GD+mhoGLYccI3Xqt0xDqBlGsn74SjIw/IQhSe7/Khv0JBo5vvfPmo
aesPpBC89wN2zQe8ZFdMIzcO6IC3+z/Aj0mudCHdAMwp1NLMpNzgJyy5K+f0/Mru
PG9ZJ/DElhZXph7sm0nzfIrOGjSYY/hOW2DXq73Dcl6eqJN5wk6YYqNEeExmCEdg
rAemiWE6RS/jtSB88ZgwpkQ0IN1gZXJS/OVriGr0vmDxiO74cqVesYJTyyG0pP7w
P3qnIJyIIbwcz7Dtg2Cencm5i9XmJPv+x9ixxu3VxhJhcrwzFKNwnzDZbWkJVzoj
NSBfpg9MCS4+viTkOUAoXdoKjjRPTG+O3N6heu+1/PFN+P526jNNfl4eofFjqo+v
wnnKyzdJ+W9RpXn0gQfSuKaVs5b+4LezVLNpRDK67FmQicBANtEcQHRIbZUd8aEF
8lt9f4B6VP22xJDPsSorO5si2GfFpWRGoSYgptj94Bi8iLdVr59v6flStWR5CDbG
vSv+QeCCtVn9VU8NHic2T4C0CaFMq4LzQ4ejD5n4YkDvW1v+5EJwBABIATgHZzku
rQpmX/k/WZwA8qI1NK9QeuZiPela2TNwHPvL577Q9+hmzhclK1kQDZEXnkyeu8aX
CpaR6T1ke17MaLwsev3gkOmokUsJCiRAvCRNjx3v9KUHMJIDMR/oR6JEn2xiiaiP
IFmocc5aP0EB9SEAfthUhqctYcZNX5W/KPSgqV4U0hs0uCMcDqyzPdqq/4rvmvwY
+Nl+rewgffMXfkl3PwZcFig6oAQtr/PuHPIdDe+b+V3J8wY+ohpBvhGgw4orphn/
bHaQ19/l/mYMPO9+3QMnXLcUCL1kRM+nXb5i5CLQEt3PdlToHTCaOshCq/bdTEuU
5zsMdFki+EJXRo1jVNue0HSnx9uyEeM3LkpOi/hNpViCqJka+1eoNqJzxNCZsLt8
7oHF0wSgqQWwCUbRN+BNv2qOgbwH6ir2b3+NNVdtmA2WuJyMjmzJCWTGy8WY5W2A
qt2pAbIpBaKWVYkyL8BE/Y+64IXzkzbEOc0Wb7P2Ttjlt5iW9eQmNIzNftE3ZR1n
LcIvQ3hcFfraAVLK9cNgQCprGimPPhhsoWN52xThqwcOCRIM9FbKUXx2fmvRoqC3
CNxqwFzJK/nLzTRd297MgNvPm4SR3mGZ82rqxbNadeDC2VJ+Ieoh1qpIIPKAsuI1
2X0PuMfGPIFhgtySDDxQkSEVyXlog7Z4MDxG/0CLFliq3ONTbJ3jtuFg/v/f5b+3
RjDKjjG32V019TSElANWDv5YPjnGy676UfeeyKOP3hPhTj8PBcVY3SU7iqtrVkXv
oxesp8rQ/PuzM3sumuCnPzWwTuNap3e/JwfE8HhzzJp0jiOONz2Hdt3NKvCjV4im
R9rn0z+Gy1RLY6dsj+V+FmWHufhGIzM7tmC3QMyh9VqO2j0sJl+nsmQwYjG/RePa
xPmRSqI/n6SssNcWtn+Puo7eI/s7g+065njE8CcJuZHb/yFct4esG9r7KLY09WN2
6a3unA+5/rn7XFPSXh2dfJYU9TtffIoiVH4S3UN1qcj0sJiWaahVoHE1vXgnCXcE
Ml2x0VaOzPf9OQWu7Sxc4GhAvacaxLlWpeMOsxn0Dt1ryulk+xyGu3rSbX1KkPtb
ZeNu6laP3wzzs9ChPsX+yv7rsPrHeIOzKGsFg+fQcOPkxCRUgD6/9MHsH/k7D1hg
RfhMv29HYGzu8+a25kNpcdkPodIrC3G9dk6cDjDcx+57wYgdknMCi39hhcAx/XDC
bFL/uHbOY1Z6D1A38cEsaMTguhdxM8/dps/D1Ijn1C4f9PzxM8H4Yjlr99d8/R/g
2M7qOrlXWwgZO/kOezVyuwJZV66QSKQVUM43LXDC8FPj8f3kv1zv7qWJCw1bJ4Ew
+lUOMMq6sHSS4g1IGYUN/CHCoAUM7gtoPotz3TE7+LuPqowSQFeUZIe9kXqSut3V
CAbYPIPyJWtmgGoEYQQT1mjt/ZihFq17SNCAb9hz/XpE8mD+/t1JvBM3IBQsr/aB
f+sPzLfG9mvkC5nj7lT108FdYv6CZVg5ZP+HM8yifoO0/Qxs5qaxUaQycttXbYR6
uolVkybfh293m6N+oPzil0rtjnX6VZDFolytW6MToqMIIz+kU+GMTkrxXuEiztzD
lCghHvbgUkZkwk3w449s/Lw9CYkdsA41V3y37uYfQhP4AKnuPwAWAtGobnofLDUI
nki0/5ldrQHPDvPfMacpQd13bDJlwcaKhLlJ/4Byq2bnwywuMy5e0NhAIPpoombx
/YJF/YZo4N4pMHxJzwNMrEByyDxULxLfYqu+dH8JK48BvocQF2bnPCfN/wXzugax
Hu+xIL8rj8AKfc6p3bymgL40WEIch/2DG4y4u7tki01ukXR8RDrXennxwE/goRO7
ubu0wmvFzrZMROWz6INnsPNcmnVYIR4IEd1s/wyVxQfteXfXJjX88Uf1HSvNQsgk
wSGXkGFLNefubq7wF/JQDbBISZO9m/DdGEyRt0z32B7gA4VXpvAE1SQ1dV4fCMgw
FgsIh9Aj1/yayxVIULGVCbc3ijdGuseNVDlfZ2qr2xMD6qzGSaaMXcuHRAbpFwKp
VQS0mYY+dQo3PhD4ZuQjkF6Y1WTG44yfe3UXAEFz0IljV13vFnKUV1X6q53a1+rr
yGDpTpFbldoFKmOUE5R60APheUMjaAl7n7wjcDwcoVrWE2OSkfPzr+nWv5z88EPZ
8IdSRLOuNVKO1QHVOf7B23FVrSLkqD7tfyg7opQabHZOZBW9eiRCaH8hEcDCCX4z
xDVBJ923VzObhYF9Nxm2pwVQ8jjYtjBLqeYCHaRVErt3BV6zxXkhjdE1IuxMvXqy
0rLL+mqdwMtrmIcOf8aFDqOUo9ybVJTLPSRoQJ+V3j0aYZbEPUCKFBZF3tSm+5Y6
hFDr5nB8Q2dsvSoyKDrV/VRF01RT35amLekKHvdOU/CHx7QJntw26gyzlXhDhSY/
oVL/lG9aANH9MwV4egYben15LVT85cI07Kk2o+Ky1CXmp3xOv6klOgANluNaI7QF
GVqq/YQODoWdsUjco9s50BOPq6ZAFnCnSGXYpTI9T16keDPh48IwlCRuz/OtD6Nl
y9gWFY8RH5bP8ObguZI27Dn6upkjBF3nqEIpHi73nB3zGm8WewI2wloXlTPtt1Nw
39jU6mOXrVwYujAYSG7qvZl6y/IviwopKImW3MzhbXorEbUQ9cIdjgb6QtBXn1m1
q5CGjbAir2uQr2xQl9pLxpPqoNbwKUgY87g+woEsgouXobZI29GXU6YYViGnGRBJ
Av5s2gyiS2XT01AmOkVjkyZe2LByPyrjnvh4ut/vyT91pieYCAxvtrjm9FQE67wF
WlZhlVG3reDeR9KNUDU6099eNIMLmOvg8ILYBFd4QDktatth0gONZ5nkoIcmn86h
tvhhpXtoR93s8nTFy/OEl2SFPvDvI1hPXQ+887ZUBVGFczldB7Qsy1U+xQ4YWmZS
CpRw4DSfiFQAyTUlwAstWG79cvLoL8vMbYQ8Ut3PybbnAaeLMi5uI0LHSoq6+VTH
WVG6KFEv3FwymJxQwnEcqnCpNEn0KtDu/xKQPL/h+lVthtCjyDu3FEyoNS0fCRaj
rSaeehfKP31y87WcjbZJOKIHpA5XFIwtaX1037EpmJ92eOkNf+gEkWABg5Ebxq+b
p6K+m7pjX12Z9vXu1/fsPfF25LpCWEmQnfpikiT+eCGZcg4MVvRI/cxFmRynhXMN
FyVzYJGIz32G9PYfMD36PlI/MoH2nma3AsxUrnNPkG6kCHBv26TA6H0KfGlTONBk
yjcoI0cC/mBkccRSUwfP7ynjZ+RCYP3WWGbeawnZaFm581oHYpY6LdDlcM4aIRSy
nRYL3CYeTwntCDe76z0Ufm5HvbcAceMQkwO/zRMCQ8q+F3o5ciThsYSpjunuKnkr
eFiYxmExSoT0kRgyGL4OPTHi7g9gobLSEnbsWdlTPgTwq9/UjYuGg0Dww0CRbLg4
ngE3tDcwNFpO5d12iOHRT/TBsn5voUf1+Z/ZfA4Fi72oFIzJf9ad0tDYk10rmTdL
CPC+K0ALaBV3sPzirB6ZufBN0cqeHWMvvNGk4VahrQBHIl6Fb1lVcc80HJ/2QvkM
0zYw5w5uqRO2glKU+NLST7068EfUYgtYUFzM+jCoLm95koWRn/hU5pHZC8fnhqaA
2evs7kMKgKfhCmtoCHmVHKUM7j5EEdOyUNd1ew0dtHSyXCiW+XFQb4bSl8yj/wHv
tiF/VFe3pfoP8K/XzyJE+eKbxyILsoXhnjLOOThrOOtzNxoA1bXilWs2DO9Gg20/
y8Cz8Z7kCDFGTJEGgc12L3RO5hJWIh65OB3GADeUWwO30V9uKr4suvc5cFMhy7vC
2ySOXUMM//RVTGXoJcMbaxRA68TAXCQxMsIO1I9wrsB79U3MIW37Tuu4NSwFDo7l
FoTGFG+iqWPDmVy3aI6Xa8n9XQuQ8J8UHogXEEf5U19agDnVVgkWFYMUIapCwxe5
HncqWMjRoJuPc7cTVAQ/jIYNMkOHEUKLtMf/RzZ9aLbKeZ1Uc3m2/RLQUSQAmT9b
9TwIIBYgwshJemHE/e8u/Lh052hRBYqq/SQvHS3uTElPGSIeoDCjUv9EOfwVCPlx
A2oFTqjo+7mBWc/H86XG4KEhTkjNbrtN1pOJbSWngr8vEiZqZeFfXdSJOjjfCHYw
9jt0ZwcWC6kVFlDRuPVcX7y/3CKW/8AuFE8gMETsAv15T0AM5XppyF2wXOdT4yqw
bVCE8N34gzWS8XknaDU4Tdg9EKX2/cCY7oCmgCgUiJFoB9Kuk7HDwfjxgHrlwamD
TcSH64j5gID82xxTyU8fNU0DLv5Sa3cI9/jZmL+JJcokmGRjf/MbLpZXsbdfwDmr
OdGtFPPgdl/JVnNNrYdRbJcLQ+BYNEnX+HoBSMVOG42RwNVUFKCyy58Joh4G9g4e
KSDwVzlhujV7Z2vAGi8xraag1EbM/SLenS1EIv0QR7M+/eOsQXU2NYbuGfLbqirO
7LrtiBvDXjWSnYETIgwG0fGNNpVRU3JCaPYcphALV19YWS6mO+20duCarv8iSjnb
eEy9dZRhp6AKczw6/FjU12XoS7GDMGSH+buez1bdhYkYuwabZ5ux9dv3mAaK2l1K
j5iMv4v3JyUmhijkm0jTZgSwhsEzQnLUeVeHvbziz7wfl+MeosD0YqMACDCkO1Ln
1t8dEh8w4ZRE+g8uDpjSxglfq6mFE8h8OCLD5ffYvshZ+BE+HIFYs4qNfRslBXDF
lk/zAaq4Snhrpz4CFQl5hW0QQzE+83DUtzyCn59Vun6AgiD2x9SSxFbwdLYhUnJ5
tyOF4MPzLlc2wAJoCXT/GRtIo/24592bsuz2st8J4xANUJ1GCviOFNbwcvIoUe9x
rPHho4uxXC+VS5p/t68ebPrfmisAKqTVnitn+Rw82Rt0q6xdatlApWhXgkuCDHDI
6u/HNajg/9whn3dlI4+UXr1I6GuRntA7xKnan9RPa2vD0ZAv4hXWz+4Aga3TKFYc
Hpwd68ZuxBBbn5BHOMtn+cj9YN843XHg0AnlEIO0WrslDUCAB88nyZrjyaWE7t5m
hoVm6j36J7bMhc8Y5CQbGePg0HzoC0ul3Vceg5+Em5eSTMOWCUM6i8tJjQqRzudx
UvAx9cXQ15TQnWVh2dVGQ5olgcUp7AFgsJlktao5xRCAQmebhRnxa7miv41bL8QP
hkBx+ZfkEJ5DYGZaX2lIeGlkx/FO69NXf5BGdaf7MHn+bhcm5I7sEAYB8zSseTQl
LBaHFMM79CwZTqwToHxRqh9qbs+Qku49l88ffIRC8op3i3SHFCnOqF9GEGHGX5IF
/uaCMFzuhIpvtOuZjNbNMZE4w18MUMfI/zLChB4ymtsCbIZ1Kr1YGMEZcnDfnnXC
8qjbdZR6NN97JPgm7EsA/TSmzdHW5i9hLQyOmN5imGk+PGKaqwE4N+KO5OyctVif
579wpyCsjqoIfPAWFRgAYJqACCgXAYAKHVdXjxOKuwod6B3q/CD/lQNit7pI640k
RuUp/B12Coff0tCJX2msCjZX6mC2TTLXcrgMentGgm+/YnkoyNhggV5KpN8mEAN1
Rq7u5+uqMfSA62lWcCo4g+FpxArXD18RJk6By9Ubj4rFjAFivqQkz3VUI55litwh
uq4fEK8KJoopSTjUabYX2MBbgSSLUB2tf9EXcEDxlAm0gna8jMCUHQ7zClTG381L
T5E6W0aZHyZWcTSgTR6KPvxTkVq4C51/nQorM+/RqCfdlau1QqKjAhWb+tBAzDlh
hpcWvShkEXXrp2xSCWFY9hO6ntirRpl1ogMvpJOoTVssCXrt5ZsfTQLArb7IlOOw
SI7RflZQQM33yAt1BjXnUUqTjIvFYjcW18C3PwzC0g9gziXLQD9f+7zQ4GA6zWBa
ZPxfUbvx8zag9lF2NCQ+SMsxBprdG8gUrwMbtYtRQj2QJuYaC8OYY5owZ63jfgm8
T+Ptn8JPRQ7q+qkf0kjry0sru5Mh9cB6WYdGeQOSAabY8ODacL8TykMAbdpSL5fp
iLIsNP38tSANc8vfUu6qrvjgURvtTMV4YrHJi+caHKctoJFceDcXCl6TR0Nve+Um
0qsFpVVNSGbPeh+2hjyY9uU7CyTvtVFOd2uz3w47yU/UdHHLE95MvCFD2LM+9ouT
aXQfLonuAAbRm3hQJ5OiFwzsyTns2V59Ls/Y61MVhWO5NP9Y/p+aJM03E5AqtC+0
e1qRemiIVDZOrQzS467Vodjps2fxMeVA0fvZCxR9CXauxXOCwJNL0PMLXJDVGSZR
kgj5NHGWpmmi234n05Qxlx367vg3WzoBE61qBy82lk+E1afuQ54OhvuqLWFg/rNW
QzK4+ypKVzvnHgoQwRkMoIrrrIx1mHMLPiJVi2An8UEvUqaM1tev5+GwF/1Po0Ix
AzmIFiYKVrMVDL08K52fek/fSPMbmrxQ+dqxZu4O+0UbkAb9Rg6jwcaRK2Qjl5a0
wLX15OW6d7El75RW17gah6KTBgcHPQnpHPigRbSR2k6OG1l5Dvzi2yTlABELHKH8
+jQIfpUuDVjEc8x6zQKoga8w3CnTynX1DGTTDSGd2UfB0U8n8ZtpDWhB7wBrjD1b
z/TvlemqPtBOf2NNETkevkB3f2rQOpWN77c5Yyj+Qo9rhdbCie7pZtS40Iq2CyHr
0PLmlGMnItPsK/XROyprk8IHc+12culFyquQHwfQM/gUeLIRCktR6zqTPYwsf9t/
Tl6OkU22QODXalvHzUszoQ5gHof5Eoepbx1w5joIPr2LpmicXonjr6skGM9aZssh
l670FV//5InNDnwzVhZvYLacyKMoqdd7t4b9mEyt+ofxE71Ov2pBO9zSvp8+5ay4
ICJWzwp3pPs4MeqrvPtpOY3sRKqSCJ2ua5WpkBSj5zRp7XUCnB2ttqUpav//0WWT
Gn5OxuniJL4VriUyNAJoXehmSzzC7EtnSNIH8T0Wtjp2SJzR/pi1KVvxxT/aIjpA
jdwEAM2OBns0RrlqFibNA22hENU80NpfclJz89OU9L4POgtZLxB7Ly+JGy3WAZcx
xFnSyLoLmhSXTfQ+1YUWII4NSkNuXetlUnQRyifFjRIyIfs/4s/yWV2mQFmNoDIJ
AeGlsKr2PcFUBhfTHeHOpZkmU2F+vZOCBgMn3hXKxozdD+TJKd3VlJg4iNKTXlbl
3IngRQw7PteqTfWR+rIvxDWTqalil8d/uvJPpgN9+Eh8/7Gs6o23skxrqgAP+6Ho
weLs4EJZ52ks8RH2jhVwaE9tqOKREqF9PGhEwuDAVFC9f9BNr1vZxRXFOSe9L5Jt
bpD3hMFO/A1MS0AHpxGcqBIKH6aAu4XQMz/nNA/9mSbcTZMf9MShFvKeoj12REZs
bnzeW/icfDjYGzb1vS0n162SVkFjY6leotwP6a6FpC5OS0iktHdwVtEOaeV4zyHf
FyTG+cSaMFR9ylMnawXyOM6DOBnvSNIcKQpWE/5ozFNjEz5a8WYcmkl30aVrkTI3
fk6I+lwltwKN/cxi/NVkLk5XSuwlHhvsdovm474I5vDMk9mJAvjDOfOZsGjBpQjH
WiitzUXNyUnzFZRfWIYfQK2ogbOf4oHK9XFgSxc4Rc6wIEfIlm61LtpZzAtMCrEB
wxy4Arqb3AwJU8A/GMGwgFQuv9+a8G2Ko31TaKpfc3ofyfl5G1fUGvIi1i1PxUHS
CIMhshpAmWSNJ/sxqZY/JbhScCuNC0LzG0xOkElVSubtbixt2pQuH5KjOJDXrY33
xfX3E/Lv7RztfyXy7/GYUMBQE/q/38rUdjFC+svp6fCQqo1N/6UzEdLm9K/j/Y83
bA3Ep+tLF8DqORffQpRoeoquCtqiwSvJfPAgqdis9zi0mFsDxDKL23XTH9wT3u2Q
wg2i7jJetNimNzoTNjCLhzifAAWIbCkz2mZnh45IEkP7TmuFh8fhHO8bGIe9CIkz
CavXxxbHAyY+GLtVjrM7aCiVPR2erg+ZjAqA4UMP/YHM8PuxDh2DTQe2kTarytB8
4gYmd1K/gwP+vrSSNq4Qu+XX2KvyqfqURzd0AUwKHq1qARLv3Uj8QRSAcfqLrIwa
7B+04y8k8y3/S7eP+KbzohoOBztjAIoHFXkcZnKhNT437smmznPb1SjLGbUd1uGb
JSX6rA0AUl10liTM3yWrjQaflcgnbhCQl2d/fvdNZEqwICLPa33XG76veT6Kpv0B
nwLqG3DSmfugEl6tsuu5esm52N16M9z7qNlk+IRYmAU1LF5I6A0cMIHx/M6QHut4
n39BAzRJKqX353CF5Yi/m5G4woigNlW+AcxuquYdkZZEHkmtZjdeEPrFXiMKONB+
qCy9q+2BjWdP3YBQ+5RM0Ika/Ie93HUCzIAPBClbCdzNx7JGn/1oxv8MjbgvOFQ4
6YJ3cS05coF3tB4pbFTOi4pZdP83woyw4rQvNrgGsQ/uP9Otg9S1mI7NONtsF/2N
oY9abX95Eor4+oZOuq/Jq5jGeKeEDxFUnNHRZBH3facKuEMXBakpGW3NUnvbx4l/
IggAGBKUS7kt+ieZF0gpL9RxSw/auyZkgl+PqnX84itd2oud4usUyvEvcfQaryMx
uVMe9wfwZLXaEo/JidCCEkpYp5QOqEXdp5MLyXhuCoBfSbuy00Du028j/lob0uu0
BX0sm+NirdFyrPCrnMaa3800CDGanHnSBVThd/5uupGl2UUSXmuOas3abwz2gscC
+L/DJReAjKvk6aCxY13TONbmGxHXvxkE0JXN7F95Mm2xoAz1L/IeBr7JxiOQekE2
4kE+nesXTlm11LOGwW6d6Z6LImyNWxosclievwrkAPr6/aRv4VAAdDU/KIqtZro7
h6B2R7csuXouU+PM24KYyN1M+d4y8HwM4eqeA4eDNR0DxJL3e/S2cBoYxK82jIwv
TVOa7vpWBccgluX2+915qhbehuGwWxqoiPB/ev4snOZBAIKs6bIXaQl5ll9fxTco
cxc4esV3Wc3ZFiGaLs0iqMEhMKoPKjlZmUiXYSP9g/xUuTKt5vCtFyr5BYElWv7k
yDaNXsQrwym8HBfhnJBUpe41cpmaDftVeVrQKAQ+lDw27OSf3WpckBV76Gy5r9Yi
5YhRLb5KkyOtJy6xjF8gsWWUA4OU6BJlvTCBJrshMjipVTeUNhNV56zMI9ewPrfi
vmgi+KXAgsxvUWpJ9BFWIY+wkl2HRBpqTUP/Da80Il+dWRUl12nwu5ufsUn6HzOy
W/gwHLezxTMbsngg7/ibVtlT6N/crICwri41/BdLsyfj0wkyESp9QVZHUFdt51NO
1bCowuMkVPMFZcon1J2NLwhv3xlIIzOyaAC5U5XwRyQp3SVZY2YAhITO7ZVRZZid
q4a6rGP2p78yq4iLo0uASUpycta/GofEQ2McwQR0KzZrGa0kmRRbQebDd8Jz3CGl
YtDGFp/xdWxHf7h8U91RhZHJTD9xMkQf6ZdL8akevRUMCkqYixUsei8tR4il9OE7
PXDWlwaOtFWiu70rZTy1Sk+3+0a7cD6YH+0Bl8ePM20Eyfx60AYjz28QwB4eWOoj
rXdcnVXGAy54nkqFLHrJME3enke3wDBI3r2Q2U+7nToPjMdxIccQkMVXQtWm7d0W
S57xhO5JSn1EH+EvxN1D8ekLamb9cz4mvtX68IEi0MhpcFLFZRiRB+ruYP2Oq/k6
Qi2RZdMhcmTdtP93nOKNZRXGuSNRGLq8Hpu8cmFrj90brRJipIcusgr5ZZhSJvoK
MXNTFW+0AtSeMxIxG5sHXvv9O4+JQGCZ9huaQH8fQgNWT9VTSxkY5dnjtU9H4q3z
EgeXmKshAOZ0ERy8+l8p9tZTvEuCLG1k+b81ZJKaqBL2ktD4NC54/IlrV2Syu4dT
kRJ4t+R7GqijrgPjSO/C5lWohVtjB+VEpAG/tzmI5e16SFW5LquDaYS8x3V00S6p
SGxwXt0079IxfHxztf6Qf7RA7QJ9i/Q6e5bS/Qpodmz6Lq+ifih8lWvTo5g9UOkp
u2ELLiymx+omyVMgmcPeXRTzbXWO/TpyDiJcGfGIP4/6YII8G+TotldYh7r3YjQt
r5+g5N39gLwkeA982uJPj8OU/3liBR+DjkBs2ocsXojH8QaFihEiPKfQ9m+bPXWy
ZGQTUMuQo7/SC88EuusMrpLH9rmi+6lyngSLg+utBC5sbvOoFIOeW0c7XPyYIDVW
h9OHvOF6uj99zu9fNETHcz8unAjXiCK8tX5XKWV4hupRp9FseQLltsDMhmEPwHin
BwBwBj13v9Ld2U8tQYt8Qh+l18MUZ7t9NIIV30XoRH/CRE8Dxl+hPbpYtlsAnQUf
wMzAN3lMZrElQRv5Hi+q/Yid03sxpVT4D3i+56WyIB7C7eqD29QAPc3q/qRRiOxc
9x0vJznfB8jocdUM0CTyXI769d22EEq7KYqDtqXQUhIR0YM8T+nLtZA3ezXcfIMy
mAQGsqaFIAnxaFQ9KVRquBua2vtelU6SxJo1uI5Rb06NihP5TM+BMvqYQu74tSv+
WjPNLLtvSybGb8dplCaQcCpsFUnH9KZssOxYUSLx6w7urDgVmh07VfenSlp9W//H
IQZBhBd0NbH/Cd78rrImiDwRqfmwIK2S4u+t6C5J5tyY/FX7L5P6d58KRcZahBfy
dm1B6OV0IGLEw5aRiaqUAbO5gjT/2bN+zL21YExn1rFqN4QeNuKhp4cnSCW6bpYq
Kj3jp8v94rSTdxvbnXIZfYiKtS0Gjy4FmuMfrtjGLxiSaGrENj65JO43eR2NULnM
qHd+jIK7BCaUhOhfmxGujRAzqbbD/JCu/RGb4ky03Hm1a1uoEbedeoaT7yu1j8Tp
rbq0/D7Fv5H7xsOTvXim4SFq7aI+hWHZ5hzQTRcgP3U6Pg3r6SW2YYWiix2UqRfD
n2sz/0hzqyDpwPolET64BwiBFXyaaD+e9T/ZuNnnNjq/nXq0ZvOHmePY2uilNgTb
b/wq0rZFi5s13tUoeomYM72DjzU5sTKmgusNoTu5CxcvdH50J/5hpznpQWoiwFdV
1CmU8iIYQjbNl9z1TrUXN2EQQn8Z3FyliJ/+UsJ9folIp4RhkY/73hM4vTgrqaUC
sRXpW2Gn43tNfpK27maysPyjee3zzaR5u5qIYHHJGdfZezYeOyKgAohIh3InhNI3
/K87/Cr6GcMbnA6oJlK5EpSSxDBrMMV76lvjpDL6oDbx7w2gDv/4Nbypwl7nQ854
JlBjxdPikAaWNPNMVknCYEd8KOM34JkuUQEbV6+ZULrmxkvX0LnhSGdxbTtN1/wN
Ax02iNS/7tLgsoLEzRd2c0vDsekorOAMvrzX433BSjYjsEjjXUgG4bDGMe/Yer6b
vhHllobPvRs5BLVKxKiBbMN+FY0d/QhZf3H1RzgcRiFeYgFHo/mOKzkeFmesYhCQ
WMrrk1ZJsgniI+7swIR/4kF8LpkbGdSQ/go+g+tPVyL4Fa9PlBHEg/wrMg1kB4B5
s5Fv7swgSA+XZvRVAhe4nduqiD9DzRXG+yYPyGzCRZLI3IsM99rHkNqe4nsDqsC3
DsiWtj3xdCvEsAihu8YG14ScAGn7/JAXuANTwZdls6/zCeDrPAniiNtYj4o9o/gJ
9JUVTk4aWaXSR6W9v86+/Hnj+u3qWsNTwisY3zxuvr8FIT2rdNs3iUQ3Y3wcssAU
DMSmZfRFovvs1A4IWrQGMs0WcEZGqFUeAFDsjfGx+4T9d0fpT+Nrcu6N13iMJLom
+NKUth6bjW+hCT1vaYqLRudG9YALhQMa7i/jvsQoUmwKLwsGDAfLQ4TTMc63pxPp
taivxuiyIXpYuTH0yDYI1VKcdotdGyzZer0XL0GPcE4AQMynDxnJ67TPO/A8UcU+
PFyzUpDuWhPTSkasFWFf1EqkIOlyRzc++vbvL+0oQVSyiD7ztSScpkckHmAaFjTk
YkJJ8iNcsT8+GV8XxXGYltkc3W8LvcMG5Cg//HU1QRKaJRVfW2IuXdUnYMXmisQH
NwJg7YzdzSl0e+4UrzIgR93kRkMkDHXqeb7PjR3Vn9mVhsOkHOq0wL6XXMe0VGAK
hcyn0x15vsxW/LX96okpg9c6+ETr8ZHuTeMahFyEHOCZ4x+vwP9GvgBLJTV2GjzD
HFIZV0HgUz9ONPJzea3XauzPj1PwNK4Tm42AAr3cnA7whn6Y7UCCl1HMZ+KqTsKg
ZwTF3h9wNs+OAVFT5dFWuxUJsYPbpB1ed4EIJTEJJA1L/JkDENVmYMRDdM4eCb3c
d6PhX+6QJI4NAXTJiS27Q+LwPEI6Y1tFm6OXqVYY7F0MpzUUwDCQpM4ed9Zhie85
H7NrRnixP7bV2DAI1J1AUTLy0zkcLQ8C9W0TUmUdghhNShlVpyh4FLaMrRkmokZo
9OFYRyTxnmIDWzD6rZdvUExKyTcGvnPKNFUPCVeyRNR7d4+HyUcASRrwaIjwKbDZ
YNOVeQaO+qTMS3+A/QWXrScjhuJW0AFahxZAWHlNFPOdy2y5f/B3g//P4n1EGXfT
gfyILHWMBZEo5lq66MjfrQygcCJZkGpFJESsFSlFLD7D2YrpT1k7OCUKeWKMsmb0
pO9yVgch928OF5Hz4/vI+gowD6KBS8dvT5yCv2IC+8QCYkFg+eVOgjhRk11N0YX5
z9nNfy98IacWOIZXgfaQh8G5PQfdSVFRLcZOg4nhzTzJtOsAG/LzCZ7Ik7b7ScEc
N+o24opBfaAj0vTSFnQN0dhnWCcPZX6MROm+k1/NFmndjXG4tzlCFOiZWHXEOi1w
cq4ENCqJHX2gL1RYMfSaG+Z9tdQnEElBji0jKFPmlD3v3DPkmoHiA2jsij5zVaoD
IBY9wLXzFtpnm/EaHjb2zFiLoMnccH13MNEfbTyKAf8+hvx5EMn/faKLlNk5kp3j
nlCTdx96TPmeiD0qC4LBCKYvDnqcUTgA5cb/1cHmtWnVjDybO5UWiPBQKKVaQovU
1VYZzP3cyx57ABBmhWkJDHrQMEiZ4E8uqO1zJ/5kNTAtRtBqlRqJ9d3UAWEa00XE
hEQBD6z252wmxXudCQ49/KPO+sR2IamFma0KPifG8BWJc4le941FwO77RGP5Fg7X
SssO5TjdyLXbFdeuQYCxWMzx71lLPhPSoS2WJiu29i4s2geuc/6/wA76FaaX7f/C
LkaSxbusjQVHdz3VxTpRWBRN0eNcTdnK2Cx0ybB/Las3kTXgELVny1Le5Xc/aJ0m
2t7ju4nBved0PwNCR0cDE4zXr41dL4HJiHRaZBSoFpGZtSHXKWrZ84W4CcwsNV6s
1ynxQ8GhY5hnD329ByaMVdol1G7ppffadSfUgxGIn+oW0ob3XtUNPKQd4IYczlU3
C2+n/pfsUr0BlRRZdyLdioDNR8loQ00PeLN9Qm0RNmgaPAcqPlxAQTf+VCvJCAVN
145I4iijQINpF4TZ/xD2PEls3rTQAP9M5U8pZKgW+hMhz+LAwrrQmz2dEBcqqHKk
x/4CNuKaJQnhuZaST2zRw21p7S3HG/wm71nmGoecwDqIyo1lD+6cwxoAsS60oz7F
XTkSnnuz1tlGo/8IfojouDjwUsL1lTS8A9va0V1yhfd8V4MUbeuIxvW/Mkcl8E9Z
9cv/6C6US1e+GkplZtFp2/8hn7+/uon7nbeCrC9WJANqdTuJxLFnurrFOdTRg95w
BSkjRgrRr2I6N0FHc0UOte0Q5lW63++dJVd4dTEX7JRY2O6L3uV/JpioZxqT3BAf
/Qd7QgJH/IamYkkaLZ5K5CUwA8KiNw5hwPpZslprCex3fhsS+ibdYnL/DqNmZZyS
NoGZXWXYucrsqydleL3i12wyKBwP8c3Ls2P8Qut/LeAKmnqGwnroybeAfCA1vMi3
oWDK+ixwfiqH6xYgojwD8laZcYj2k+OpPsfU770xDWdhdVgGSLmSUSDT3vmsb8Cn
l+R2sr7qtSNYG48arApmis12185Ta2Uk0f2OvzbBmosH0ZbPaLng4jh0vOqng8qz
ygHepTVoJO3uzuV+AsSl9oS8zhhe4bRFKd51cL6YDjl1ptZANKjL1LhdPJ5k96Ez
6pBnEuuCRpdAM5OJXJ4uxdEo5Su9Qto2sJRmxqFAmrVcwbOE/pzID6H3DbeyOD4G
eieLRqub2UFDS8A0Vv+ERhBXharR//9CqcEa/cBCWuisVZ8lyP3QY2G7iN/wl11E
dXOhe0fgWzsOwel3ZNC+G5ZE1p3CEOXSqhHSJxvE7P2mjBtY76VJV251vUvQdsIT
eJflIpyKmXa4lXIGNw8c2o/ZJ1ZeRBjoC6og4n6s+/qtlDxpGynUdmckAxFnCHOM
KaNOc8AUDqrmsjR/4gv7Cdm4JO8FFgDhrLALmJq4vKTsUsKUZBiz7UAKTPMwzGI7
LxOR1VVfnhjAxozHqasYARyUDZXIuyqhbJCrkXdb8jNOshqV7Vf7h11/Owy7kY8q
nqwu+Wa0ZwjoyaYdFSuiA4iPwPhFJMzrdXI6nDdczhpwKJLHPNdJH+laJFCISSHb
/Ir5ypKdgePIu6EZxPgHBoJZ7J6MHWHvvVHOgKP90AO/4iGUxVO/WkbK7N2HsjUs
Hk+xupLY8B4jwOZOIVBRZHBzZGX5G0DjQcZ4Awjjs8gxJwGcoiDkWiuQzfMWvA3R
CW17D4FEzKWkyMofq2OTPeWAHNlAIBTI7kZkRrOyTjpsB7HCjuHwnNnTxdv1TsX2
1Q9HeGp+w2ywlaI780XRC+wRFecjswHtnZRyRAoezOLxddhsxDoypeK4FEVV0WH4
BXGZnNYKENm9y6pB93ppuOkclltrHI4ZSn7rq0VwvvmO0H14TxyOAmqhSTiXw4A3
j/U4ghyxdBPwO0s6FSNHLbn+VpJ3dyfMYbHaXsorHf6PFQJh/Ox1Cql4WnHO/LSI
clEmgS+YT422/7HiAzCmXBDZLfOwBe+1Yr6tuwDURvhlsWkDXa4IoJXekQq6L6GZ
JQPiz8IMqt6sDdI/aZMtOIYJNQ/tOF6l3sFF+2ughrShIWGPhIf8tNZXKq6ACpBq
vxZ9zcDk3fbKPFNx9nccncVsSGPOh4dp2HehBAHy0VhHgDjQhaemZ5UMUdn3PsdO
1YeJORmdyKDr6kAAz+DnjuQkzLHa+e/rUU0cKHQ4sAASRAV4XuOO9Y+o+aMoeh2f
8denVQnUHeGqf+35B/hY0oiWiViHru7p24q4XpRgDQaid9NAUrBXtS0l7+45kkcV
xjFGjNbUVTrurSSi/mTCzDfObwADIZFpGE9OtHIvOrXtAv2lK+FyMhdGfM4xiI6J
JFfHjyvjBnGpNpI8PcMlNsRN0pBcpVc2rDaNzXtqNvP/JymOnZZR3f3V0yXNHYsu
20YFJzCxcYpSNsf5xg00CCddj2hXlXSpN8yAcxtj4DY1GTQIKPzikx2OXhFYsuZQ
lS8+cfgyy/+VBp1wcE8k9w4z/ledD6TK+Rxm32JLdSo5ojrdxKUJxU50mHEcO7pj
S3cu8fhnn2PmC5X24ZsrqqDF4WdwNxWRsju1iDGmcQeVeDuYLxpw7sCUzCtx0zDv
uDH/4F6HMB/c+RAnhXgU52r1T7cDwi7gzWf75Y3htdFmt2SyQb5EEf8Z3JTm1tqV
b+zs5zx8toeYXZifrefHth6yqcohWkVRU6mNw0e8HT1i3nW89VLpdT+sWzAFdRj3
FtAC8haMqPvVMkgdyz7Y/4NAWquQJhfJwrF6m6fMZY6J8RLKTvZZNoFoB4+y+0KT
CVzsUQFsX27y4jhwElPQnA4KM1D2R/BZz1KbMQa2FXqz9KV/CwVgSCOpKkiI4HE+
CQKrZZQpaOicIPvKI6zKtWuL2USfvfEHecfk1SjVq8UrzVTUfXKLjvOgmFe8atBz
XJvHurTPydpBxfrPVGlxZT5hdNRHAAHsD9uFd+/x5TvWcrPiijAvpSe3PdkT6tV5
13ZNScKDDE3z+jESLSI+pVvr+JhTV7yS7S/xIMd7KoVbdTJoUbeNtKV09S5bMJt0
bhclD+YQnouLYbvA5WGg9kZOoUEkq8dyVk7HZISb7jg1pOq+dJQSoaYkwKgQxPQK
ZncqY/ONHQWi03c0RTdLMIck1K2MWjsJgvMEnTNx4U1cKQmXiCqZ6l5OkWchGQ65
AyQLSz9vkn6UKmh8v6FwHM0Dao+pJnaD7hutuloh8mTxENKd/6oOWgusO3xonxzV
haoMLTudHMgPrxqklfdOPPGbrnaQsKEZMaelhuTiyQMbKi+YtCS09zK519FvpxRR
LPjzfeY/I7k4tFCr0FOMoq9PC8rylNWzvaqanbS0lISKqVWRweoN5onYDB7eGyym
rJ+1s9dZTSJZKyCC8T0D+DZW3epL9ih2iC5pkB0/y+3V5dT01pv2eHkrbdNOv8LZ
wOKLrVY+zs1xiLhRyXvJQ8GjdjB7KSQ727nF3cHJ0Mtqd1hLMEfdSiulV8wNuHcb
LkCygoCmq0kflNOglF5OIBoHSatQ2yNcAA6NiZAg100yetSyHDGg8SsbSfoK4/Ml
ErMOiqBu1g+NGYzKDOVDj27lpM6rhiO9pBvdahGS6XyEpkcXsmyiDQhfPVJiCG7s
A3Xr8K7a7rCDYDplOigeH/eEWxbiwUm1tES+iIY+TYSPOPh6P3KhjVMd6PKPxDxE
vLMxAx4nz8D3uryy9pjBQdi8cGQhZ+cTlCOnrIeGHbs9ifsUMdHzNM8alGweux/v
428BeHrtcGDh/AktvvvFORGhxhwkTQw2njJKDTqNoZ6KDXCYKoBY+RSCKeYmnQEo
Z4+JBscTOQ+N9RvCk9zmGF2yFi1JLMPEI2THEBLa8t0Dbq5Mmy0ulHpAHEmABI7T
1wgnq6tHxzVlT+uVpwnYcMMKDwoEeTewhOPNZWfNq3uciD9Hvq0qhC6Iq8hlLges
dpkiUUPzkfrZcmYZJxjopuGof+z6VuDf4kePBMY/MT6S5LCCCkfqMxaEJK8SsdgQ
wwZR9nbA3LhCEUMNdhaUnAsgiOFkyZ37W5MJQHcqzXepW3AQ4J4vSzboTxvt2dsr
2tES1Kd+4D7fjjGTS2CgKmJIVNJqHIUgbT45NKlzIVgSf4auq7RQSwROkiCZUUkW
HQkwg5JmJQ32UAHafh+wItNaGa3gYXanff7KSRPUgpPQDaXu2XesQooqPXze32s/
RDX835icBXc5S+HU/ujlv4h8q8Q9TKd+o0WH44ggEHnM1CpBPRMBOxmQfYgzVqkQ
YuNLirnYodbBDr2ARh/zKx/WbQRW8rdysg4qzy9UNJLKP6akzupByxteJdgSUEvf
BQ3EbUttGkscYCLdpC9X3o2rNiTjvg+ZuX/bI7kZuMZ8Ptbl968t6NjyaeZRg+SQ
ktqoZYiqiT530I5BmAM+sj+nXV1tNx9gbiDa7RJewZ2VCT6nESdEBa+DEPrnfQ5p
GMQalTJ+F/OxCA9NikIxsQlyIjJ+n3u/nX2eatmulwOAAaK1F5rMFjyznYr+iOc+
eHtI9v6ygOgpsqRbE7lrolzp5aguMPel1DVqF3RXEUKZ61GdDh212L08ASWzo1O+
MZ4+q9ZkgheKn0Wilau6YJpq1fPN90hs3Ij9WJOgUCrsDkbEZ5zNcoCoQ1h1N26R
6P8wgZdz3mSjgsS29JmG8ti7JRPvEMrIub1achD4BGb+yW9Klv8Q7ezoKltqloV1
TghusyknfwifLmDRyivTW0HEBfjHjCrLOUeIE6r1NjP5XIZDMBStDEzCB+aS2xhm
DnkSxoWMm5YLwQ3flKD1k3ao3cETyTrhEHICAyG1mUpG+Vt1QWHtXjX8SYCz0GLa
7bpUCMIHFe/V/pWTOP4sN1zyfJpLCz9UzCCVmSd75mITe8ac/oz+UWVsuhBT0Nmg
/Vd7cp4YJH94E8N4YdQ0G7wacmrTpTMQ101hdFqJhtcAbQaNiddjE8+JUDWFZplG
N25O5WB/VVyIfIywZUGC067/+GBBegpxdwP1yJz1SFcGnUD9rzyE3PcgOJU8qCTY
En6yH3F7svHNLmPFemQSckOkSh6ktnSCtHBI7dyniejZbunOoEhF5RQjCnaVkpk7
EW8dzjyenwzzPa4+8VbReQUPiBcIUAJkyjDA/RJquOn7gLBYWPcVSS8vAp2/4MFZ
BSvtijHqfkN7OxffUtZnaVtk5Qe0yF+9ZtOca7km8HNo8tT+OEr4SoGkkiXGiBPv
SdFC+GL9/Skcqx+Dalc6yfcbjZ/H5VuQJZzHYWtHXEgMcc1hEWetZrpE87pKLb7v
X+7XUZbsLeK7Ad/H7J33yuHyK6L6d2Z8Y+L3P5b2m1t46SwqMg4s+vtFmKev83IX
kudWKqwc7FxPEcSozXBY8xXhL9lteVHylogwD/9Ema6uHIGxqgKjNsG2DmdGYnpM
zKYUEs/fSH5rKPHuCCeP+v9NmrLfYeyVVhAQrmnFyl9IHRzWHzHi/oo+tIQU2g+M
QJ88AtTPYHpGTaBaagI6V5hDoePBJYr5WFY5e5J0mTD3DndjSOb2TIhKF9kse5dj
lI/6PwkoZeHVz/qYL7SQ140azG9ZR5sWQBE+PK7b27GzQP5y1eSoI0IdjJ2yxZ9W
VrvmWNKJ+NRHH1jH2m5bEQuPhgMnOmDd9tkhJU6O4vNfT69onaWNFrXO2eMbFpS2
JcCas5vyMJN5tTfzSSKiMEU66zk+D2Kt7FZLb6uC3H+qg2PH+mzuOa3zIReO8dOb
iyNmDcJIJQCeGI59/Fki633DXyYMB+59Rgmg3X/99NVM17VJjvuY3TSlg9aUkXV/
AApSmvF+APaDGGMvxnKFl1Ta+kIrOM/49+yd4JT4t03jmkVmFVGs8gL/Wb28Vrao
J/bL+CxTHZdbz92AvTWrX60ldBiPEpjkpTmiwHU2z3FnFeue0oO3bHg0uHPNdSi9
33aYaBv+L08U6kPoRDDfD9X4Ds1+J7Z7FafCGavID49CdVPWvpeZyKc/ZflGs0Lj
wbkLGvVrOct8BsjxqadxJwpltkmiz5Foyy8j+OktCM9oU8XXPRpCW4mmZv/+r/hY
58gzcqIae/ZlfSQ/T2rKlzyf2lMYZH0/xPINdL9gmMRyKEoHP3J2jbI8ZxUJZ5KZ
6bKfFuGgf35RnPXnHidyiqfkCiCfDN0wlWFp3UvwuOSZI1OotrIQCOrYMvxLo1KP
44xi7PeLARQLyttMQxS1rQ3JmJdPGmysV7V6T53M1/jn9agYfJrGMh/75pzPSem7
3WCPOZeXkZb2XwLvrq5I1NUYj+hqFwlONQLEEWtEGVHG/ckwIehD6EU7P6eaBWJk
g4QeKg0ePPfzO0d312+6G7Gn+PK79vtiHOMfxN+XurTs9RzbpX9hfrTBGtnxPV1r
ICMrvyWY+OtLZIyCpuIsywKwCUjMFtdwE2emUf/jo8Uq6Nt5QL5NshOID+Ggd0Dn
uZcYQLM1/m5qaVJ0Xh1mQwtpsY8nmyJ5AsejXDtOQIur+1GmG25cdyAKfOLCxf+y
gZKAOkBGndRybpOFIDIsBMoxp3GMA5JUeatWr9yNqpaPoNFg1nG3yOF3SjAuK65c
Xvv3KUmaNw93cP88JPuGmV7RMbdVgM+FlxzeGcAZk4kfnvKXYRg36cAtRQQ2ul8d
VPxekCK1cnqzWg/YwwZPlDGwybJAeG62GuySozYeAEc9rY3BFZzaBSFc9vNXVC3I
G/SNJck0MuaF9vZGP2gQbnPv8/+wRrLI9KXgn6+CuuZF+yXY+ljmPCK07e6WZ2cs
0dwiZ6Fmr6eaYuh/w8BvT8X1wrbpRXsfc1YjKbxHr5Zko4qAQS7Ijf/aEpGOOlrM
BsZadvDHrcu0Nzl3fMw0LKyPceS2AV13uLSPybUmXn4es0ATOPIGhoZVM0cjwBKH
LH75x8howHJqNyDgpVCanZ45bXe4lSyX3SaYFtOPjPHripQ2CFHoEIYtUNjph9XI
5riB79yyI/C79jwJR9dJcw+0bBKRA0QfQqP5F/p4FZyjuDj1pUeyO8O4+68LhRZx
Rr+0kNMQtiHVae6qSoQxk2LAcGcstbNTkAdyaNkrXo+aQrDh3eNbmRqjBKRfA8qp
xjo/6CnLgau/4mgwKsUr8OTvqX2YBl7BCBSD5B/rrvvWHmoPfQ6V7be9VW4OGTvR
G/FvFAfTYANBEKHFkt7ggED+fakhTTliwP2jtsPnbzPM8ex9ENIVyZJNvGOtuUVG
v31Y3xdIvnS4AIdd6xNmCo3KLh/U3p2OiZKSZ+mAa6m3Q+nyANKYLBxqad8Q1oaV
outM7ogoFsH9BzR6aXVqbImksDsvLqS1mH0YX+0rF4XCLWNTpkPqExyM63aj/p0v
Mb9cvu96XN86mV6LWYybJx6K32wqvnjf/PAw1FBV3Gow9OatKS0fSwWLhPjCz8bw
j/chVsIGl4mejMG7uhPUSs6r+Io5GoPue8cIlyfwuaYVI7VkSyPW9IQ4YQzJPqJn
NWsU6bmrBK1Zr2hse1KIOj7Hkr7RFUyQXXvUSB7LI1RClnOBFdfkNuUWYY85gFej
Xf8romNoDsTN4KiG6qE3m2AxOFbxI8X77U5hJlZMYIU1VVaGI+KPN4Fx19Vi+zsq
U81fWU9pz7xB/iyTYPWZRNmX1mMO9LxSqUgWTxY+KyRYSNHOT/psenfN7e1Hj+YA
nEY7GHfcB9DS8Qwz8AyhiyjOHMwh3V5JbglzvN0xWrgirdy8fzHUdDn0PSeFswIb
tUzeh9xR2nqtPQf5xJ7EIYw+UfFkRpwnXJ1ErSxMSEfWVe18DnRgL69xOMJlevLu
Tkr12Gneh+j6S6NweKG8iCrqZ1MKyp/oNN/Zty3ovAuDYzmbU12SPqn40kdfYaGk
PMh2/r+B04VQxd040ZizvVoWpSX928WSvGsvq33lUQJYMrBaYZn+sM/x5i1qd9Nz
f0lbkkQ5DhRUju2fmNkB8Ktq5W1Dn5evGcyx6uiamVOU6zNo8K/vv4k3OfkWD8SX
e4KLKUecleS4rs9KIid7I6YaitZB7KgElXbmH18jLU64lOb2cb8Oer5bxbO6hxI5
Jy3xi0kx/TjYtRMcmSf/NF1BbocfJJdk1QCTIiM90Y+UGRUKLyXB1PZdEB0lQ7EE
NBpzjCLQzXtrdN4221t4nZoW+fKBR5I93iBwhfg24zooKOXFUAbCDChSdemcgRds
zBFNZNhVICYY23egOgGUmjBK6STVgGPCwJobYOG6R842LTi8OSfzXRaHUGffvPNS
6d6kWOwUk0QeDe5XPn0sp/QErfqwMI7sLIHK9KUEi5P4HJyoZ5khOwDFthuu4e67
Fx9K+ndUUTa/E3wSD9r1hZzTx04KxvWDqeITJUlBWGBUmPdPJA/iKUmARalDPrtQ
uIw3RpXryKcfaoBo3ZIlZUYsKk3DC97tE2IrdaEf2oFTa6Gzqdih5kxLGeawX3YZ
QzQb9HzZqfuW2mZl54a2Ata+c654bo9iEdDisD0c08wwHPw6og0mXQxmVwmsy2jQ
8bIoLoRgNqJmX3Y1NUs6hsN5KuLEkMVoBe4Az+l//DjeszfyofShKMBeGXGqfJv2
eel26f4KVIoVFC5dKGUsmnlbtAXSb8set0AXFBO89qIlPNn97tKQQ6rjNcKuFOnv
ocuSI4XOvX5pQSgqkvmfSDIvbZwgO5gUNhCvtqWh3lJCNpFAfkc5foss869c2q7C
tHC3yGSnkXNL9ZCRxZCAPn78b/eGacyUiu8AJQeam/xK7cJZtNDmvm24k3FAC9Mp
uCrSrN3wEMIruYiWtD6Icx8Z/PfX1sYNvKGvMEkr0DlsbO/yhBlVLzCn4TKBbiZT
8LoJWyCnN6hn/SW34WMoB7wrxLPB3MzW7zfvZ7WIC6Swni6nFNo3fki8dfVk21yw
PDn7FqCzmYqyVSXcr8GL8csCspTtVZy+0bk8cCPvv+9Hr0GWUWKbO9iXO9VKjzyw
8SNsRT5/rlYYbDdPjCnhXEm6BcGTjzIyeq15sxSr5MFAvIGZ8HHt1M+OmMKcVhXC
ENjHD02qFjThKBlgevRuva/7/pVXL4qjsR6KAf3OFZVX1lGA91OUwkaw8V3keUNe
VeDnJPi+n47TGDbg4JwTErb/rKErO/+QxJhd7XdN1XB6RyYJnXAlGWErQggpxhXA
4L7KRVzzfrjMSidx0AZUT6ylXAD55LEOPLesi+atUUK2Aao8+pCgy8PXE23/dYsk
eNOS7jWxLzY8VZkXS2l8wm44TFxtW4TdyH/ZZAxZSSmc01Bf/pq6s993BUA+RlD+
fbRWRUBZVzSqhSivS89s2l/Uquub0NEWR+hWTPYm/+cTDJWpifuYu+PCqOie3vwJ
O64h8qtmY+cr8PNTxqBQr+VTGaGBucjInXUAn4xBpG6277tpdc1mF3O8xWhm2F6S
9vHV4mmWWvDV+KTBC0zEM2PZyLuaSREddWn8q/lLYZJMFfVv/nVrKQipC24+V7eo
fsug4d086bb+Ea8gRXDiTdJFy7dhQwmhX6joe8jsaavDaEzWL2UC1GBEmIM6iiJG
jRg6UDVOD+N+u7GSVS04sZLWXZ0bPYFm1fA3/MOGbVDbQcGrU+sO3LuoLp72NKAt
u8042hu5ESyfh6XkymYA0elXoD88HNj5X0lN57X81FnFUeLNrHiSOzoDT/Ze5lUc
95KGYFweAq6JX30nkcZ1BehdoKZcZrVvjOpTpCqEcx2R1pHvEu5v839cmssbAsdx
sSYxMGAkaauKxRJJi0UuIkxe6CzMSbU4a8lSjHhWHFB8AWjuqts+31paHDNAiRt/
AE/Z8RJPuKqlt9H9EYGvIApBge5eC/8WQoXuNDVbD7r5RcvMzHIEMCvKS5Gb15g/
QIHnLTqeP2EbokobtHCp06IeFrQswWZjFOHj3ih2ByROEWc7Izvqa21QQYWGPFU2
zzUOwb3YTpopEmfRauYEKquiB2a0ar9sA2G+VZbLW79/2xs5vV8R7dMwl6uCYyiK
llN6hpC31svlIRTUZizWffu4WKRp+zszG38bMv53WNSw0RyGOMdwH06g90cq+05M
R3sB21veTsqyLDRSboJj0vsSBsj9Q8F/zCN+gduTOeYoA6P2R2nDQEuCFsO0CT9b
tZD8ZyxDsBIztqPjXcQVLw24gjFlh+x0KgLhJPs9NfoVeWpe4N9jnlifpqJTLZOM
54tl+C8hUYwR7RC3NYtWdXYfymTaEzSLcvfFXmnRePnke9xLyrn32RQjhLeuZzko
dhqOVpHtCYWy6XtNNuqhWWT1TIHT+no3qMt8Wugp75fLcHmd0Lx9/xzzSPSuD5gK
5PfO58/nPmGjDtOa1srqWMLwe9/mBIeOr/7KdPjeOQR3wuxTlgHxRPj8jbWDvgNf
Z42wVU07nd3/nbHd9AZHZHwGrrjXWGuCcOgZkPkmWKP42F35acpwKAAt9lXVHg7l
LXwZgrUZxFC5K3FMYsn61vQCDbCqZ+IejqkB8tBs/WhTSRrJNkPTrZQlIqNOeUsk
anTNbsCutHCXoKKHyqWZOC0XcX2EGZxl7VxtAwsgV90VrlYtYbK3blWNYShgsA3C
YFv7fQFzneea02LOPIuCRsbklpq50woiKROV4NFJUS2UOMMWNqiMFJy9l2Qc024i
q6FuJxgv3DRgDSFHBmfYBACEgxZotsHeCR4yvIjI4YstrMWnuFN1zch6oUdy54hC
a3kTOjIt3K17glvXeBaselEPQfveE5YG9iN9ojMBj8GYph2lsOqPwfeEM5BCOEbT
QG2jLBv2GdcpPIYGcThWW/uvbySe3m5FG6zQtmdimD4b5b3TWtufyaMPq+JRBGY0
MlwrHvuVSQCltmxdPCb9GYYnVHvjMTJ5Lov1CKOmqi5l0w+uMf0ZdBDNnpZFuakG
QbA3UOgOiZrlzjdfhqBqM6s9DMBVeZ/np+eBmWBnKIS3DQAu8aWisuJ+ek0HL/Mf
SpQJlwQee0cNg3j96bZrYoiZFWzkAGF1tagIDeUXmRo836aJfqbpCs9dkFPxCkVL
XrkQwFW6+j6ij4Z2TUbpbOhihLE2YCC52Kk5g9aHIfcYza1mGv/RamD7Uj7+8g9y
YaEAP61r7Jze7QQFNBajONkjOEu5bEdkMGwt/GHwrqonEZUe/X099bpHXrOqQ8HK
yI6wvue8tYWYdo9kKbwWsny1J5GhGyy4aJKU+bolDMaQ/eUOKPA0oDtdmnO9ILgP
ISNtqIWEJ3DyCaXLENK55ZtKLzlaSh9J9n2gsyo4QaxC7EiFTABFno+q4/QL0aBE
h6Gvh/AoIu2XNeKxNfZnH/bN/oSHu297rCNUd5wkxWoJ/nImuCIwfdmgOAYuLpHr
+AEUL8jgobHjnrGVIjL++3Czwg/oKbDq0g2xl2RTWQoVI0M6ouvF262/1ekjJcS7
b0khd9xFkTKZGQYsIvVRTKu8XQrBqH0JeewNzqxvHUoW2OGc70rciRXE1bsDVnrb
wN0uFXln2KDkvFgBX263MyeNmZI1O2aYeXq6jPpu3DjP1nz3kdYCi0in8ZrQzmFk
tUyVfjmlMzcbKeoloQDaXJT1EI7u2PVWRs9ZV0Xm5NoHXZw5biOajw56Zqgvy7M9
TIAdCV9B82b7DYNsTOAepNDtebLQr8ZGigLXBTFNphn2SJFLNvaHrMsBhTeAsUgk
DrRPp+TRZUDw0f74SnideQrrnCiRYsEqZxEy2fyAakmWvXMe5YvX6krZl2skd2fl
zZCMjkhqaDPM2GUdSs8A4Z4q9rZK6ZvTyYN5v9XjxB7xps4NOMdxna8v3xhZdcj3
uZlFryZeJB/1Wsc/QouXxhlBlVUSSRzAJbED0V6860dLqGolcTj1R0sgduHIWm0E
3vAgmAbxp0WGfM+unI8k7FX1Bwc1Lm16O/org9izXVQx0FX3Ayt06wIQgHXPYRt7
zdXFnWsT7eAq5XjXxC7YpQMAHnj4yM9QdT+tHre2GDLGMA7Wk8kDTemU8Atof+1/
lGyXzbws+YLELRzmpcK43nIZ+92OOH2H574+JGqmWeOH8lFxx9Tiks91HYQUNw1X
eb7iULrZXaMYuFGXg0NtqGy8XfRr0wj5wDy/Pt+T25CTKAQOguQfp0QiXy3GPtIv
NrZ40RtnpcQe6+qYk2PTH6Arn5zeDT1vC0dMxJU+QQl8AkevQcEI+TpQbdz99Sbz
Ir+AzC9h959Ug9wyNg7ceKtOdUT2AgjaqyNEhWcH2dLpTmoz7dvRGDppzHzWzSyf
7oVi96DHPz376ElS/H1eSa/xfwnkkL8ITs9hLflHbP79ZwWkk5t7U1sWPPWrps0I
5vKcTiTVsUw5SR6BK77Wq6pANLICJ3DCJuUWkVZmv3setWIUnJtPgMT1CcmeT252
+AmMAxFLDYzR1IJC/01FlSICN38EZ7ofzdszorL9lGpyjiERNgEUQmpg6ZpJHQCb
bQSHIz3CVDE/FXL5QYYwR7JBnk13HLSupJLa4AVuyNyFcElEMNtmiAyIJc8sC897
F8WRaxeCtr8kkDNClbGdmEvj21U7IAwEzBztwkRdNsSVN1XEYG8fhnubpCE3V1zA
OuiP7YhqlVaJ6X61zdGxG/zPwqrYbbzRIZzTCezkRBfDJ6CizIjShB3kWRE8mxcv
/89v7c/rVEeWRxNOjlhsyTvstr97cCMOnRebifP9Ivvudy7jw9ekRVTe4sC7eRRO
pF9FiABCLvTauiE4g8cbraytNWTzbog3iy4FLlxs0PIiRdaahvQTd51rsPCu+iX1
gapKo8/VAyMP9qxjtjiUXfdB0PiC4iUKgUeLXcwg3bK5kQ6/kcUs6t7RG4RbIPYE
9PZIoXUIjQZbt+zDk467BEXhz4EJzWKvmnNEvx6mYewuogVuctbG5r0mq5SLC5gL
m96NVBIwe1E7wer6Ii24+q1lhLF8OIRnShA4YK6/RkeBsrCJd9vjWZhSRb3br+On
MXl4iAhMFwZOKfHTQDLbHsY8b5pwiR7l9T6Sh+ms/lArwnDwWqrm6gbimG6QR4xB
//5p5UfmeLFQX7H5DTOt3edLdNjxtQPJVO7eA98HKMymneKJJRMj9jcy6VNl+ruG
r1nVjFOmAo4l1gEZTTIbLNYqghNrmUf6KNSwjcFMG3/ve//w48JOv23Imcp9fFlV
B5s5okzL5CoRb5bSoV54KVrndpsh3kmFnEwp8ITl4H6b8trgmqDiPKz0VDgJk7xN
dr6cMx4S0a05jWnUTHn9gat2Wv995NEWGqDPeSrD8yNf5YZwq9gOOkpm0hyfk8yx
EyWxwLXWHdPyaTljn1iQ8mGJ51XhWGlU6HpnI30aKm+Z/qcY+79BMVNyHPPf7Iso
Fz4gMn0YTzweR0cXzO2gFR427XybLCT9oI5FHl3x0ofF7rX/QCTF4F+a286dS2z+
J8fDqmD1l/NGdIF+9fa3FVrtFy9kGl+bcnZjB/ja0kVZrDWBAuvsTZsC0f8MDXoX
TflRfhzVl0oaMZc00TqY/KKfjB9gaOrjCQRsJDN/zpwkj0pmmKaMLkgnM5oxQmaM
CqraTaGEqR77W+CyMEXDLm7FVVixexs1i+wtWjUeEDHNln0+aaQXTLsbEjE7WMJt
9V8sQUM2yITHDViyoOx/LSx5HgTXDJL8tUT3ATZVrZpg/VDrwIOKBRxW/UueEg49
OGbr3XS/fnDqLFikUdfOZVsYV5CoaJZR1tKjvf0vd3VNgkiqOUpLRmnNxsHRJhY6
KwwIj+Dcdz9c+lJCf5zaEoWU2zhYYeVIW7faG3xj02iN83G3IVw6+XWQCC0q1zp/
YCGbNZvt8Do8lSAgBVXYMsIpYrx2HC7EO2g9pkJxoTBbMBx/RUzj3oMuPoV62C1w
Jkr/FHqROWOHThL6vTY3EURNlvQUY50A/TQgt7chYO3EADW6dnNYqRX1CVEcxgok
mE38wFcfVCOjOg4cu3CIOw2a7DxcvpT7I/0lWwvkiPz02qkW04KD2PAD7Ax8sXv8
UofmntSfyE35kdvPL0B/S+LPI381xoDr4BnbEWIOseCgNBhhIKvr7LsbCggF0Zgc
4n95E1nXhgExQGlI6jnS6wm+9+HKrhuYTHsQlUHUtHbiDaOyk7016muXNQGzdnFC
5gH2yf+W7iWUd9KCu7rQCOIEWbgm/+fUtgF+mLfZMfd2hQpwXKrsfahqS9XXmsJv
B3FccI9MW4zbU/06h0QYLHYfMBUgT7eMUfy1zCCo7pVLuaL0cghP0P6xcuQ9w4jF
qbOT9f+m9OdPPLe5lI4qYwTlRLHMjF2l665+46W4r2LRMBBFIa+OCJLbuTXC4nzk
Br+VTueHkpNbgm7ZkdAulfjjdWs15tpXLDmQaGgssM5RstAWcFKL8bPZaqPX2fg3
fgxOlVqtjBFvGMXQEKXSoABHGIZWL8NTtEgff1c0vatkA+DpiabPmcfqMZOnC0eQ
eDKf3AS4VPUpA2l/a9TCKK3DKfJHHGkD1PF7j5kcH9ROm4C/yv0d2XWwMB57BxUX
rSeIsLiLFNhb56Ciocz8VU4FdaTVUbo1YWxpkINPE/4+DycgONzy9YAU5KL/Xghc
6ll69T2TDx1tZiQU2QJke51EiMlD4/yBfYcii0o/jum38b4kToiFCBnxvUVvZbgD
bSFHhZaRAnhZzg1u1P8IrnCKAOpTFt3W+IPzTn7DpH4XBjwHvo2C0JqbvXPFmuo2
3Aa2fy45rHuol5RMqd0qg+2Qx9MuQu/AAgd3tO8+8iRGhJC5XyDQZeY5vrwIWRhu
zStm4r/onF+1mztA8sybVL7VIIjz0c/jHul43tCEQnUNgrF4olP1lMGQZtxHX8Qm
5B0jdayiPdQjyUZ3OWoDxaXh8JL1sRxonuZDFpMUVPd50qnXkes0TKZfiLiw1Sn6
iKfi3sGxYIE2JzBG9or2SEndEDE0jhM+D2bO9iyKZarQXUoerbkAMXbJaSdmAEvF
rxq22URNjKGstdnrgFyR8/Z5G+7Tk8SZV+e6XUm1LSFqMXyNz4fMLZTqmfnwm236
NcWrbRVlh5wuzwHtZx6Bnyuhuz9WMh2w95DD72K01ciUqYQyQGIGJ5uczY1u/f+p
S1JwIhJVJmyON4epc8PibG2Dk7RfMpUGJE/aRr5oeq7Bz+kIs5P+GFOQrXRqC0SE
sBllkpu6Bsd+T74ffVBcNiItTPr9hAjSomFjTqPw78ng/JeDJxjlLEtEH+cAn48z
d6lpKDXpzkHuqLVDreMbJCOToaQD9HLMDBFDX2mVBf7mHe5ZSBI15u7GcZAOasSf
PPsVBgSsw27lCI3znwhBzdHmM4J4stSCANF3liuyfVqQkHw59nGsZmt5wkY/SUZa
0qaq9IR+ddGG1jMLBE8nSisZjdq7LF/B/bGfseAj6hjXHqwMyX45KYbUU76mqJAW
7PGR+rHSModWLYR7kqBjmXQAe1nz1fgLp+ug0kXK5QgMKyZLrddnqkqARixb0o/y
z/Rz/J/FaYDSd0uaK0NWkttiW6WKIFmnweWOcsfjzHL6WukjojiNV0VgNJIJ1gVD
UEqul1r76KwBHnzF+yw0DIGEnxeqn0yD2vEDuQ3mz1R//l7vtTzn/g7FKUc4kM6P
JPcmmfj3QWTo+6mBqqgrDBomfbIMkA+xQcWOcdj+JnkhMJRyi5qNCjaFQSihewWL
TP3ydI0v+2J32Fnd0ITqrB1dDlWVSZv2nSvd/LgCu+jX4WSguedNohf7BtVReycS
UtoJfvD/taeTDzsxdV204w/Ol6lDPO2ckpuu8oiB+hSDaYcASlcDtAlIJ8sh0o2E
EI2Fy4d/OYVtjcoilrhyyeuWeMkCYQshJlreUTBlpw2r7RpCowwabzfQhG90GHCr
uY35eLNvLU6tlfFbFhklxfSzRPbKYBug0RCP43qsAjS9O2w7GHYfIIqgfNg68fcT
HswoKyZNNNnh+Kt+qDn14pwn5m56lBRPrhcMcpaCojNeTALcKxuGG+ftBUPgy7Ou
sYj4UrP8OidLIAuALb4kyKJ4VjI5hmBQuLhqH3NMQc1Qd0QSUb6GoQ0mqaWepvpx
Up7sEy6dF93y7d0/Mfhw6IRgCvOyxeM0bDC87WoDWL987ZjX28cyNOymE3dW5sCu
9tOV6UzrxdIN2KynUpBZ4XK56swmMt0d2no3tsenv/GR9qBNT/Cx3ukEFCEzxCTi
nMIgShqUV3yZNduDfdlv0HFENOv9WAcsMz5LmLc7tUQOt9jtm/J/G/RvxRIqWmSo
AyGUR5u6aPqBeMnWs9Ky8ViOXhtnPbJ0jc1lljI8VA/xhRA0jBFMESzwMLHENOwF
fd4/ji+ljeS0LGtGwBpypRFgxIw1ni3wvwMwokIdGiTCb33RuJLKhDzzI5wXNI6C
66h3oqTWOLqDv6j9hidUHhn462mMmqjEU16Qb/9Pg0dYvuVc/QhmCyf1jruA86TH
y+kFEgHyOA3ND27mCXF4pwLW7pYbwf/PO70SyBchSjoXW70BXmyHAICO72qBpzSK
fmG8medKChwDz2rRAS81f7g7BaSxV2BrkAC2+nLiCY/POVcuKk8Xg5nnxWAk7ZuN
NM9lqqNdjS1Ien6Kj5GkEWWZxStX+Xb5Qgy4BzQNxJs2GxUjA2jF0tlyratmmdvy
IlTjP88VXc3jbokyeaWKERGr43IFChGa+wEIGI3Er1W+bn+buYnPojXb7biHqRGM
UZ2VqhFEHf2tujt8mCMVHWHnje8vEdmi42l9zQgP4QbW+1nYDfiFhmUzan1UNFS2
QxCHkcuGF3NO+4JoIu9L/u/r3qejWD8qRXed1l811p5z8uHclrRQzF8rDKHRkzIT
rXdhlTVv4w9Z6KGCjRqZgkXTwuAMnlMCbv7XbJePKln28nskQWBGMUTs8YlmG2hZ
pnyYzP4OEflCYeX93DPQkGT0YodLyaRXQ+U466EJO2UAOfW43BGIlUTX0Eeg8K96
pW6IYtbYAPwC7jLn2YlZ5LlKqvgNTodLbAgLyhkFNeRtpP3es/uCiGHGM3QvAdwj
nsaOv6NwXw1TuT2bE8aks3HITVg1yuNIHcqZBoc9tvxl6ZAn6KtaNoAbSDMkUiny
dJASOLXT3nE1CDoBDYqqvr2JleVi9RwETnTYb5faIA3rS8lwvqnFv8k8ilhrKnPd
xTj7yoUlPf2+AIhdK34oELC/nTqJLOKEzCxaPzhgtStnl1mrCPfDFrY11S6bCUzb
J1g3AtUTX51st8yMgSL+fVIDObf5sUB8VKZdXUK92RT+vLh1D83NWjyqMXc1fh7w
+/MTE41/h9bsVEPcD+6HcDC/trOdyQgwGLp1ufx8x6nMfvQSeABTqfdm0nH8blN3
QBU8ztwRLZAQv2mWtsL8c4YmG6UEKEneAe60E3+I6frZrIevzcPHQbVjXisy6D/r
EM0k8hGxcVO1ow1hOajRQJw2jGmY2Jl0QZeU09kJSsYk9N//JlUFYS37+kbImDX4
M+NWN91aXjkuFfVMdUX20y99seyjXwy14m27/X/vasGI0qb4Zg1ncavwfU7M+Wl/
HjseCQ4MUSCRsipoQRHZD9V44MnQO/p2fYXUrr1/ieB+y+lOcB1tZsia8cJLhK9r
WmiFZWdY2fPiOoIfRsGFPOR8eNICtVTaIcenufDRegcMD1TbF5vWe3jR9BYZMXeO
UwIV9cnceLm/n32emwT+cKxSnuxZeX6qggmnSXy7yvYrf5Ie36BhzE4NfC6GVGIp
sKO6JKfQD+BHG8wFocExgWTiRywuVSUCBrse1I9laFBnzQUaETaaz2QSJQLdzS5U
mUre7JOzSCamNphHavDkE7XnMA6MuTLmZYqLMCMUGxAsYX0SjVnhhcCafSKTB0eu
eIr0a2PUR/iq9tsyr1XKlgsumS5vJXT4q8kAbnNLTQM4PamL+cG/jxZQCo0uSyDA
6TLlYuabn/069AtVSFjlqr4yT0mCYfE2C6Q68t0LyR6IY/wAH+c8ilWLP+IeHMqu
ecZsbrT+Ipc3B/K60mGMZSbLNUqjLmdq/Xy1EcFHX6192yDwuCqMjJV2Lek2cRH+
4AUWqzr78aBOvvhVskWdh99PeD54cBUgLlJds18JM4RaS0YtfUOrhoIvji2o4H8n
VQnAuP3J/O7SAmp7VWI8trZXHJAre5fgNhjuufo3TG9H15Y7r4v3qqAkkFi4fLcK
BnhaUWqOEYdG+0B92TI1iXvzWtDIkCiJzhFgqvp3E3QTbcifitcC7rw0lhOtG5rz
bZnuxoSQp3kbG1U8MeJ6uPu9ijG8plEzUdqyAgBEGi3go+HblxOdQRYH32oF1RkB
ei1EntHCqFlkO6aFInqOZB7juX7s11dZ6ymxHqBeKyFk6wb7TDwJ0NATUu68yQLP
2Y/ifQSvppGWOl18A38dMC1BMXhtztpFzJP49zLvh0g9PX/AZFvM3Y9CcEROKKxl
cggjsOM0XqkOctwZGz6ZEhlxhNyvI88DxJ1bRgyRoNdohkHjOLmo4jsHh3IPmNzv
6dndP3pGz7i39Bna7Ug7a+kORu4ndcOBn1MKSbfJC9rIMln5g66qbV3OYgOU0NcC
68R/ZBgXd2zBzkJtkZbHM6kdocgFtV/1/36WcZjAsppns3MEoUGCJuiEhO5SKWHR
LNEDFf/9es6PBK1V2wCL39zbAh5l3UQWTpx4SpkTwJqgQRp/dVndo9notEMyj44M
0XA6b0fhVhppWFHBR0oJqIdJ6bbl50OGNy2aXEV00iI1zqim0nJZuz2fZJAxuEVD
Gcaa2jVK1jvWB5mj5Ztz1AZgAkoV5GvyGR3UDhherPksLJUROQAMHJ4gOyNTPZ6i
iq1ptXvqtEMUcL+JRy6S2SAVmb0+C5DM9OUbZpUhHPvPKl8pvBGsEpksyOyTBYnK
mbt41aWJipWARfrtxiBHFjq70s7GJlMz5HvWAJQIzEhkbbrT2RsgEa2w36BBT30/
lBvfcCak5W5ad4Nk1DKYaLR0AJQhmMJm69L+4obP41dpP3gEVaD7ixqfeP4sX/xG
FBb5k0ig8UHH5f9wo1SIv9r403KS06AWuw5w8BYUmnGL2SS1uzSJUqOKagMuB/Z0
GQJv+wKLJ4w8PPcZQi3+2zOcgXd1HN9+KV0qosfAKG49p6GG6gN/aOr5GssKesYp
iWzXGWcwchZhqdMg15oxxlcoOKRnl5/abu/NxCTIRqmZpnNRQWeEHl6zQlIyAMTt
RyF3R/OH1w659qZup0oRRnggiMqutN/ss/oT+1Qy7ePH/4ErUIIN/6y48dXOUCQ6
rvS5a9flpQkATRrjwVh06ATs/1mWaD1mPp6seyFQQ6FhjFsrtA0xpyqyi20+2Qpa
/vKW3JlDbxAeFNSiEkE6Uia+hYYz0/75IhLu/efuAKpW7G2uMkS5JjP0grc1XHrA
Dxl89PPiplAckBGdhLIjrHnns1eToDKz1wOpDNBE2SpQP6koZY9XVADsZ7kJeDe7
qRPTTvHhUuevz63CfhEIY2DjISVyGLu9KNDxhOFyyfGqkXkogT+Hq81w1C7gFKi6
pNRXf43pYMtkCVoGzFM3eZpCeGRhpr0ZPTYN5XHcOp22fLGD8yYepM5eHEmnhP4W
pPD3xaD7oY7N2g3GgLwYci5geKlldqvbDeHcdE6EF6PVQ9cuj+dHHqYIhNWrZ7W1
SEmFq9nZRGtluSIswnlwS8OpcQCDpCQEQhltqVDM8hVv/k05Mqk8I7Sk1rie3Z1S
CL41+ZUJIHqV2i/SBoSQvQmfbKrhxUfIo/kiL9qpcvEN0785uZCJFoExTVgOtyRK
h5whNpa8pskMoLko20ILM6Bj5FoOYEkCSTgfurGpqhJOMFF8ZqPgE3NIJvJffqmi
Qe/5ejzSdv1HMje5sUg/V421kEXxsqvG+UO3IsB5Itnx+DPruJ/iwbo9eWyolaNn
XRIY5svAGWhC3JRG5dtnXKaD+sqedm/RH0qTCPkaSaMavyJM997WXGlbOplPjiMt
fjcu+p2gr5swfQTTjRJ/1c65Wy3XvceYl6AKJDprdU2jex+UgT2YUS7UQ06PG3rr
Vjq40zqYWuViyn9r7ucQ3ZhlmawLQMJRqR9RU7S5i8oO7+RIaIzF0qsDXqADOZsm
91HQkhwuOws+buF7kVwA18shaQub/8tA20VkXmT6gXE9TM3x5KDCYTU2aZQGKSZg
ZiuhwROOIQvASD6TU6KsSPK4D2cAPHHc9jruXDjvHK28mOzf8kgGLXjmjanDNAOo
cDZgtQ0WRDFfH25WC5EDYI4ONn0IhDa4bQ+RCwXM1G1jaf4ecyjR01oxmYwKFJZu
l+YCwMVO6rFCJw0wbQDckRKipLPpvHFEKIN+zHguX4AbBHeAY6HlfLSFEhXW8lxK
BrvtBfosFz854n6WdYddVjfMgH0NbfSZ6F/Z2Q9nIB6qvDiR7m/mVzwSGpYJ4q7Y
Vah7MStLbGh+v7jB5FlB6dj1XIi1PmtNsmVjKr7GPZ9lbw7UcX5fj1kUmgY0fdpY
1pISL5BBBrjw8lHa090z3WXW8wfT2LXsQtoVNrDlOTE02qtysdHhACdsAvcBDEwh
XDhn8VOQhbdAUQo5NaOFOiGaIyc31l5uzblhGNpeKvk6Hony/RTsWzxN3diH6A+I
2d8tXNWJzkc7LvWgeP7HVxJ6MmUK2tryPmdAMQqsBE4zYchxh8r5fTMXs/Bv8CTm
ghDAprQVuq1yWq/34Tl/0YHHFxeyI1gLAe7fQgTCn2DgL3cFVEsx9UrhB+RySpZH
1EJC307A9ACO3fy+D+6bDFiCH0IbKhAh49jXRQSUWB/E8BR10EHIs45WxrSCmkmS
f88crQ7vFU8/R41a+lyQct0yxckQGTnPY7aSzX5lOJFTXIfyEn9ATfCae43J7oNA
osEjifRjHhVP5hcWLswvJBbCNcFDxaAqyfA17KVYc4v9S+rmTJR50qToekvt07xd
idN2ZSn3qVG2vSIN0637xyppNAMLvbcugY9pencUTamaUYCuMC1bKVL6QODvx4uZ
+GGk84YyFtVoQQ+jE7q5Y5ypEO/iWyFJ3gprwheTV/FMHkRBflrUdV0JG0Q/qEyg
b2pMlQXNMr/df+dt6eM1bn4qfctuHjz+DEs91kNz4sFXqxGfLzsJLBDSB01bRgxz
35L2YzapFkK6UBakOdWIyPLWuwm8+hrtiTnh7XX76p0IxfAs+5h9p/pdVjHx+zQD
1rA3yYfpFJX+NRumGfQwO5oLD6Ah8/CSpwhOjtKW5h29rDpHaKxliACHZ8DTaHme
SQypa0JI2zbeQI19lsWuMzhjGjKfiyZnizPC3aqkU9ASrCZ4lcMwgEA7Es9+9V1J
S77cyRYQN2xzq1c2qO5iLjuFjj2HRN6SXCp3DZApqY0lh+tqtTXGvtcapkGv3SnN
g5jbpR4H6taf+W/3Zh9TkjL/tFgSDqQS1G+Qn3tIL5Vs8u3+i7/GAjBGVDHVYC2+
kgjzsqMB6ieFZroAhXBQ1RokqE/6i+iAZfeD2I6lt4EZyqYM7h/SFbPPQkON3o7m
FS1JvdKgj+d3i4newRnNMy7nS3CUZ3rVkhEk/n7TdsE7Z+B3gZwAFUxAFqCALrF6
4nq+tuiCrM7xphgE1KvmpBBGYDlDe+6T9cYKFcFu8rtKVLIiY10bt2FpgkxtrR+W
trNPk7fT0Cq8MJzIcfKKeCT8p73oCSBplgqMh/xocxBFxVEkyDhLR2i/M2rv9QYY
Ctfm7hEGkIbnRCjKAHqagiOi/iF0+hfNZfjjcocyevGVcqwbd+NOFzf9H0FBwAwh
xH6YgEYImLVjIV5bRG54EZQhzb6L5EommJyHQQdserw67fgl1+oiyDRpVLc8U0E8
ZkmoIPnpx22VZc2+YHQX1m8gNRpKDaqq9GQpKRRpxKDYrFU7LeR1waA4zBmzqA+D
++98vyuxtkm+WiC76PiZuwMDG1llI97AdEojLewwUwkwWwnPIaxAM+1ChuejpFXm
+eZC7tmASxG/mLJIZ5u+Qc/KdF3xlxeP3zlSc+sDigH2eXURStzHZcdKdMZKYP5C
N6717BZqp7jhogi+vduh+RXrCqkCIGQ1ENbHettpg3TA2XCcmRQ5GK7EF+NDENZP
AthXc8jOsZOPsXsmHwuz14k9wYUAR7dFnszwy3teKlGSgpEc4YiJCXb+tsQTOeSY
qnCyHSF8ii2a7iJ+XmNKeCxQ9MGDv5Qn7BsxGR+QxyNQ+PYgspBgLkLjG9ceRu9H
8WWOK17CJYZegpFzEUT523lBZdE3y3WK+j1d43ME9Z8kg/uUgGXz0ejsvaF9R6Ch
0gtCQwvUCELW6yEflJyEaWHDT073yrWTJpWBokOW6vplblnuUkMf8RT7PRGMUS1w
xPO+WnIweLW0qQ7fKcMaKOH+KD7iKcIKzARjVbK18ZbrJgqJfpKiNr0KL0zXef4S
1ofx2QrVkYW3VkYU7YiZ3m7SevpcdLolOAB+sDhtfeM6ow7CZjuJRj4BC1CoHLn3
SN1M9Qgo+pl5uZMYPQ31PMPaHbE1SvBqt/niLHl5gT/cdLBR/bpG7yZticNZgo4f
ylALnUMznKhFZOlzHuyKLNFZP4tzZNR3/pXemFfm/fqIJ7gV254gQxdfuhmz2naI
TTZbDe2Lx81XHhFjmAMIwzDmZgT0tb6Z0HYKC7zDRnW8BcgXi5U7ghxrYKnSdbEG
jWT4siylr0t9C4NtmLHIsd8IyJRZe4wLvedmGjXoSnaQbSibKTBqeWJWcWylOmg6
RQvHK1L1w4NOMSe7szv6lFlDQ3j1QNkKGmMnhWdEDJzwwmROLt3PiPWRAUXaSQUy
qj2I0NOiHvq8eGgB5xar+pBBCT7ypU/0E641ghIFYpRZ7Ngtf7EI/y2u+R/wnxVD
tghe7Zned/tN/xiYv0SjrMPr2a2fjzEIk1SvzC7L8zftYZDTwLRDeDLQgsQN0DfN
S6KWU/Rq7MAQaQ67mKbe5VgUGnpcOYIWEOugRs7qp6qzLOfp/FWNuL0/6ijfMCdj
mcOFnX6bVvTOr3Oi+S/XSj9zSJ8yqK6Mw8k+pXfdAUP+7qJcsG0WbvYdsI9bD/Ql
7dVvrHAPWzn0D9+D9bREkY8ka64WqmQLvla4yrt7a1X3YGJIcFx/++u4ls/P8+ri
fNJZqyAgjJGjAZ8AcH1G6BDqO77ycuugOadf6VlA2dwK5JrfPSgUlAKkYsJppkAZ
AbvfpMjP0YG+D6GheY9QbI5beTDyEBKHAKrWT78GXkQ6Akmjitlt93mokQISFFsL
bEkVzAw/HS32YhPltFoOz8fvG4Bx0O8DslYCOAJQue1JZrk0dNePDYJzYAURQq30
K1a4GsEck2/eNOJco6ppXSsog1zb0gdSDauaf9vPZpAzcFeZlrM/PzFsTpkhtIa4
KdFPxLoFvGysMaqtvc4lToUnudgLkPRuy2bRX4q7sCnl9elxRLl6J7EL13o38Pn5
6Jeq+cnt+ajkxgnk5VHeTwwiSi3yb+mrvWLAJe/cLWjZFxfNBtFyJsRJRDLufS7T
AwdQualrs3twX9Lh4SO2yHBtW76/cQhk+XyVIwZ49LVQZt/edWrtwRZd2urNaRVN
NXEuf3dfS+CaF7ri3n7MUbcYKgmaX4EIYQvCXLpOmQx4xCKQ5/oyDFLJFn50ph33
E8xavDHEVsWWqcmfSQeSzzEcmWQk9SZDmrGnyD+g+kNbnVUpJf/4UOV3vkW5uVW7
zdYoBmsCzV2o+RWhl0fdhD45OVDbMRiWwOC1+dl+FZxpDshgLf2c7SBXckGRNUjL
V8AwQM9JKQxz98e0SSv8Vyd/anaB+47aSfJC9a1Sro3Y8JpGPlmCvr1yRQR1rq6F
buWWesmo1QkqFzOlyqg5IcxIl/MsofP1RjOcxHvDnaGYKMXaJ14Amn6vjz+mclt6
SO6mGJJAKCF66brGN+i342m0EF33lCWLPNoAWABp/MkM0gVX0BmCpXOHZEqZcklf
9H2fyaPrzz/kQwMsgBFtGF1u/yqB3gtNR/J1JqcarsnSd5XV2LH40tLAB92HdBDJ
x8vqN/I6uwoRp8UN6oMMbl9enEe/13w+cXm+Yx8j3n72xeTkjIfSTEVnA9yBoz05
2s+ekHAsHaEB1wb64S/kEDeWlNUl9B4EJ8sLCzHeG+J59sZU2oaUb2sB4I+55krJ
xwZHm57uO+kH9k8mgxZPYVhnTsui6rHyqCMXvZkEfH329ktDMK3r6B2uEXWmj2V9
I8K3P6e3nNSdxKq/e5KWI0vRIBrkjcGdY15C26OxXfhliaAKrxUf0snuNPRizCnU
cthpG0Nx1ckKIs6IYgdoPowNJYiFh50lnhbptSIKy0p6z9mxqdMeHl4LcIRCkE/+
u0bO5a3fxus318C6RrxHS8gjoJ0VLdq18YBihZ33J6d5JZOyUrBLs186GqEbiXNI
1gMUfWhlumUe9U20Xd5A57lGs8itZam3ifS5S0zrmi5yr+FrpOjFEwuG7aJc3DKA
0wfR6XZzMZEsCcAcTkoapbwb53smB9n8vx4WfXjS5dYZaeqrdg2XMj13wzRhwHZp
S22mnZODK+sgOJH7082gZM4N+eb+Xjy0gd60IgVJSGnqG2VCOzqW2Iz6mG3DEiA8
e1y8nlQdBRIH2sJWpLAvPT0zmNb4cv3YKPQc36yaUPXPMsEud/JVcFLay0M6f8G3
TUdoPQabIbGhruwbvNoJb43HGt6mpr1aqF3aC3DPdo4abrjl0qaX0pCnxrw5hJQ3
F0KH8m/Yz5lpDg7DRWfy87L4jPtXqsr+u17whnCy5N9nmRic+eZY5J+JObDXHccZ
FHrgduOyR9kh9a3fvpU38njsbvdne7F5bVdUfxqJpJiDsQJQOOEThiJe+fmpLENp
P/VYatJKQltDzl08Vm3FpzZzmzwm/78/9SK3QLpFoRqyJE+LBYGpfe4Ayv3Sjpj6
ctLgAe/Qpw55kYKGmcNb/+Q07ap1FpZizDsxQGFIIiGMOSUZGlKG0mJnyt2InyYN
YZ4RZYq6pyNGwKy3rXnUyBxiQGZSVxIZBkYu3B+si7NQHm9If3mZz4UE4bpDdOA4
VYdDm4HFkv9VgIteZTSffDSoHY+gb4JNEpF7qqac4lJ5K3uINlTD94wUurCwezmm
H4Cg+RJPkO43Mi631J/bxatSfegcEq0M9Y+72GcseJkLU6JmKtjYQB0tRq7zoo/0
4II8JDmRTn7DC7Y0YufikDvQ6xLsC9zkmKp3ybh1UaYudl1+NWGgrUiMgXPQMdQW
2ggnPo/iThDP7jxYEnsE0fFkFOPbAk2jVMrTAGu8MB7L4qGBwNynekU4XisId+kq
MhGv3MhbN1fsn0MRZLHG8QWYpUtCpZUvTt7kv/ssEsbs9SfVF/DKob2DLk3uZsNn
Rht4f078Aedv0fTm0u2Vwl3I6c2aDJdi3OY1wsj9iQq4wPl/r3ooU0HZkqaBG/FP
ONfc0HLgg7pMpu63KfrVSNRsVKfca+kK0ZtMz+DYlKs6d69xzGz4bLsXdSOSGu6t
da6EqOwIrwj/zeBuldzaItqD/ZBfWrZ5OkZeqwrEWwHzrnNNJWWntoxQ9NHonTKj
oePmdYWjXogAJKwKpTneItHmQ7x2wwhX9C4DigYRE566Wybu8M9A8eWsjUWRHsih
nCm26n31FpVqmQNqChRyXW5g/+sZabfruJ2M2/kydE+qkgi8Btn8Q6vKjQ2smhzh
Rmxn2dtATFg16fnGf0qImn+m1MHDAKfYtc+CMUbnkbcm2AIU4LN7b1CxPAaB/h0N
b49BgHQU0CfMkRPn635GzAAIWlRwacQ9SyiGt3UBWcSMcEArB6Vy6iDpMdlBizuf
9Qi9377F/rJ5kIYlKry5PAwGA7xkBW5bAUqJdJuDi/eV6t0GdtzOniTwRVIPpccr
JMtG/aTX+FnjeaCmPbmXqHeeeb1hFYOBS4Ot/XcLegG/qJ4OuM8+5acyn169q4vj
fXAgNGo2AVTU6wFhoCCxGMxKF/7P9xuWY/AA3R/3p7MuxL8i1WEOsjcT8AKwblwK
SvoXU9dt9ZaHNDsMEleql/KzUUpRvocUlWwRVrBouSDHMcPA4V5ODyrxbem6UcQ6
MY0eRD/f8L73VxMbU1mlh4i4s0Heni+r1HFsM1xUA6uocQi7DXMC0+FPaNpmDNzD
8PFntb1T4S95nVLkyyDr1h0WeAir9/P8BF8yurH0mjpB0wTHJeT/N6hPiC9730yJ
SK+4FaaSPk6kiM9z2vdEw+6/ECAM+PPfCaPZXuwmc7v2zKP7OHUwDsfOY5cytzh/
y0WsC090H8TLuDcJV0G+IWaZKEyZckdzP23+bhQH2v2Td3/HvTy6EbKBo5WXjAiA
TSE3wfqXlHUQcTpJuY8OsgAkms7/sF6HlqpftZUm4+QGntjOgX1qOzHekcJvMcVn
Iw7Y4mkkvTiT0yc5I6JSNWq0weFzCFBkN3/Ub1eQnNpVjnfRlDEN3G83S1s0rdbO
NyEWzdTbZ/hGIDcMITbxYE+9b7oEnFYJNePR0Rgcu/xbp+vdGUSUisQr2FqOQR6d
T8cFk4jA6VLix4gmq8AunBiys/fJ5UR+2UyhoKmGJCugvp1cps+MF6yyRfhS2eGx
pw4nHXXVhOPIVgLHhSSLuTVqkYg2xulfOFziBZWBySozfsNYkbbwwktVbGD/CyCW
x1/DXBw7UhcuBdYuPZOrpVnjQpraPpxaR/0OoFURr0GjIp4RWdUlluWK+l8JoXPt
J+jHEeh4M8CnBlVVJ4NtmsL57WHqUSWXMKwL7sicm2BF9Qj6+tj7O9Y7VgX8t418
0IzQf/Ld+Y08MbGVjWQ/D1wXUTt0nyXlnSx3MGYxPEhDtpBkY9MzUHX95XN0+q3Q
coxQzQKh32KZmtRDKQFE3LXqP+yI4Bvpl7iUdqHhxNMmZwzVCEpyjOX6maorgyXU
QFh2GDXflA6O0vv7Vo9yzkJUTZqrO/4WHqfVhmFDYEYuOvvWf9zvoNWgVML2O3yD
PIJyuCLL8qUpu6/jJEbJwjapyHLAfC6kGZW+1uG6cKFtCIetcbR4GdC73cVxCiFP
qa9X24vT4TVeI0Gd30S8Wr2Q7l1ysnBc0gJ7xvYaT6+sjsHM2TG/WEXFH4FRlKh2
TCA2qfzMKvXBZ7TLz3IT1tzoIuHG5RPE+1Gi1kF6cnPONMns7ra9cnHIGb+S/+U0
fTbgRZ9G18jlNDHWcNY0KIYglR3hnBMUIOn3RJy+XcNs4vlScjfBs+CKRQnVmEXx
l8pD5o6jpG2hr9uM0GWyRUH/emijwx40kbvaRNGcBhQCwtIezDkUJkNas9bejgei
2AAhjGJwwVdoRIDRJZ5Sp9aRvEySrrdp/dpW6PPJFPeiYEaZ6I3HAtb0DM7DCg7z
kbH9oW91bBmWjtGIHG+liy8nVS31tPkoHGIAPZQzayNggvic6+y7F3hTvldFBac5
jTpUOQfdIdLb8X1wlDpZcTgtpWJAKgQ1mJsQyP7asvoLxzv9AQGQFBNdMKTQnTwD
MKVn8XIFTkBdytncm882Eos9/hmjIV3szxVc8ih2HZRuNr4INLSiPF0yL1xkujk+
713LnBMTP5E53XkslE8C9noWC39zQ/BqRyXFRIrM3X1FDWYe1fNLyR3XtsVmBwqu
FAm4pvlXMiq5LfSlg5w/rGgeCW3iEgE98KRIgw/390bd2G2qYn3C0YHcvwIlVx9F
uyrKRG2SO82YHwBi34JeMgobidFbB9JhypZd8fQtJu53uKP/75DmmUzRBv49HOVs
jgjQdu89NnwQe79onDGs7/rSt+REX7E8Q8+6zzkZieYQIkf7Fbr0AeafI0gWPRsi
dnKodPQt5Al+tVBqFF+AmkLyJuhnm2fn/ZU18jzar7LHpq8IljiN3j1SogQlvW0y
o4QpA5fUw/Ooww4bit7c8wSZpnLfvqjOo1dMPWpLDRnBz1ceTAVvFgPMimv0NFC7
D70AqSULc7t5q//9Iv5kw/msfNQqjtrV0NxdRjtcZorx5D50gRv6N4uksclBXoYN
m8hwHFJKvw8VceEg/xEyMxP3at2g15gMg8OfJ6MjCU3ljde7Nry86SnLrnD6sWqy
GAvK3NxfhnBYpuFKqtnEt0FZdfXxBTvbTilxZLCwZsKrmvbawDotvpB0Iu28dgPp
qBdfnT3HTUDEN607NMsDa4lTDhSwtlYHTn2GcmIldTMKuSCsWW4xBqchiDdOfJvK
wFTNg3z7oINLNtbx5dv55pUPUgSzAHxH+7PUz8JY5rjjCChiA5qnlAHH+J4F08fZ
VWNKajmT4IQTkbS13AkMz+8qqyyvPTCJZ2ZFBsOpxCezQ55+FzoXHkObnii+Jfg8
ntIST5qlTiDIWCNnZuKPMioWwfGmF6nCqQYK43WO977zx+6kJ9B9RXPIvSUK7Dco
8qzlylCShXyFoCyGWWkpez48wDy8qOyBKABXb5WFgDZJRwxmbDpbN74dkV/UtKv6
7c57W3wUYfLDk+WuFVqFd3vLjoTR8vOzuGJ3z3EqMZCJTGcbfqlfkbb2JhfUarTQ
OzQj6OGJJgGpEA3wP5we2VHaQXCW+o/02Fi/QaFuOT9m2tsUiAp+SP0IgIZMnESl
4kQXLglRmnwIWqaaGRC6L9Y4NB3E6UMTYQsf0TbxBBj9stw2rn6WrzBSgmp9KMGv
VHJ/nYu/r7gmf1WD4Pz/jBAey2xCOCYjj916m6OtVItWv3ZszgYC+fNnK+6bM+0o
NquwSo8hfTF/bmaZaMQ2yTzHDtmLK40wQ4SvhDdjFWsgvqPSZVD48tTd9skSGUpD
sv2c5nUjbKbN1ENBYLa3zKq0JdPgOEM3/oGzArevpreX+c8nDkbwdihB3fnjwQIo
O1sAGtPUPDRnq3YNgdehGHb4RrLZqf1lPaY9nP/Z4LIXZWM+o7ZjF4ne9kMMndbx
OwPauSsVVuYEskTO8mxJtJDV5/nqIhp1Wxg7VkP2kPhIluZersENVuz84hY7jAeK
3gHFZFlxmjz8Hd00LUkoTBttVLU+lbOm/tO6CQvTTXO0MmiU6Vh1TwOvhg05A2/E
rPOKb48F7/F778dsce0acAo0M2vtFpy1BrNMMRH1C5Zq0lj7oKP1Ti1XqTuAXr6b
g/AiwfohF+P4/KCfhcQQSRicB9yJycoHC69q+FtwN2Ai5DGk2b0zEBIRjaAxcrXC
1GoVR9bSh2xOOqcM5jMpvQMPfSPONhC6M02Z0wsU9OuRvGk155gH1wnvm2f7Wjmb
foZVVoYLKf3WCf7dc6jRW/kBZJ1m74sCQYSBiksMLH+0ytvP4OoY+hEpD2dA2EJ3
J5bQieLLtXXEc8wHgm19GW11+/Eke+nzjA1OyL3wSe+P74BMqen8b9NUbZ2kMXiK
BFhapc3S/brrBJfJPJcEIr45EvyOl9meMMVa3Spy/wk9sBzdshhTJwWGU0xhznxO
IyfGDrWDI+ntsY7Eq61F0JoEgFKboAVA3jFqLysvzgtPclzyoZPveOusvU7DHQJF
5PI46RQhC7tq9NRck9aXh+yGJFspkIU1m/OYxE0SQMTPTg2zHRado5LwXJk3HXdq
wMqAaxJ9aMLz2ZjL1aXWyrL9wAB6VgpWLO+Syu3uyjQ4vUDsdpjYr1xtVKFEZcO0
NH5MyhA72EQk+vqB56U7ZcKGbnj5QPRlSUsx3hCVlH6lwDpDOX/qZCgASePrahwg
wYTaLx9Wl8gbk47tw7VquXehYFrNsK2SPJU69zZy/MpXcE8F4nzj5Ff+LLZfracC
q3EOJgEx7ATLNx49SihyG6OC1LUPW1C/44weIpuXsQil9aIj9DRgIoErNu7YerWs
xIDmW2dhyqpdSoPHRturb6CYxXZVwQO+qWixgTAg8AsODKInLfkw3Zs/yGJEWan8
kU+H5pL4xNOuYJDdjEWguUGetllm2PwmK6yw8EMcIxW74WEQAuTqUAcnVmDXm9Sa
i1xVQF0Dkxi9fDPjwvxIPa4t+gM/okWY9q2Gw4qRqPcjyAB2txWJc4T4yt03LCk+
xH3M3X+NEZVdCu+vUYBL8ON+nAnRG/TbJyH1GXWaJftY2DL85/Lo2m530HMnhlGX
OZePBPENwt8EdrVcdVEtzbAb6BCnjRk6vt//q+AMj1rH5Vormd3rRW5xs4pCSVH7
vOArfy3n8oH0bi7moMiAShTbD6PswpaWQbxjD3fFB+TR4DmCL2/xPaIdT02wMN+P
WUJae0yDp1SEuNTNBkXSm7K5+jpiHZSX3YpGl0W354h5+4mHDgKB3bkZ9s9BQwO2
jo3rHsSxS3465G+RSNX/xowS69HIb0TVPCrH0S/ewgiyLNwiB/coeb8M/2ZXPTXJ
aES9aCeob39bzxSeSVj8/ZYvE9V7CeN1VaXxOc2wznT/jXviDL3OQ3cDpwG55Vl7
Xu5oBDO49EACvKM0l617buWqB5VRQn/VjV3qRGsXveBClvrHKUkGdUZ8fIOQpkH0
6tfcH75EbC+fjZkUZvM57HAyPDcWuZkfQRQt9UdHLg0mln2C1cJYMlOLFIMXhYQn
wMCHgXxO6H4zpUi2KiYGziwkMeLOzOd7g5kG+H741vf+FNuLR1p2tt01mLKeUcIJ
5mJlEOp4IJpbYSH9vecCvGbyXTPkTRR5td1f+U+vcFpwnntt/RDKNfHxQtqxudZ9
bjr2ADSE0wStauKzX8+/brtPj1p6ZxO3vqq7jr+SHYO6lAh3MmU9hpDDPxivyl1r
UO3RWsZzBEaeIenCQe9FJAZUPSr7jj8DEXdh2ihTW3fcsKXd4k7iOrFISTqoR4T0
ncHM2B/CxxfGH3l5ZQAEcWp3CNt36eu/GE6Y2IOyQi1xZneSU78wl6kw+jAt0HB9
NQTeTiw54kXW1aI9lEmEKI+9delRdmZzobmIAbHD/0jvK/zTF/zvfkGEaeYeQS+F
r1vwYrETTMKttUV+7rtfa4gwj3zbwItRnp7zdWWWh3TgpsFxYJHn5NpGvbim/pkF
skhb20DfKIqbik3yGsyBx1HwZyGkCHqnST7o/v/HstroiCpjnkKn0fTNHHHjZ5SX
mVuTkyLTqKkyFveXB8Fxnsua1UkHzRVY7LXLddvoamwSPsMHhXa88qzkUFa7kSSr
LpIWa+QJyc6g72Ah0UndYXGBESkbbNRzeQKE5etOLFrUPYYwiKQ5ElDuC51mwW18
JPFEFc3PCUTCJE2VwGTsjDLwlZ3W/ydbl9VFQAzOR9lNbRWoWTt644TGimICBr2W
/eXxVrB5CuJY11dyq1qymXP54qmf4/vmGi0zTbfoFAoiXZAjrFIof+cB8y3oykZh
dTRt6YvFBmORjesCpR1kYjWrLLvHzyrd6qY5d++sc441mBTAE/pmH2YiofP9MKv3
09fKV6kXinUM/HcrikrdeakEKWOTBfx+OmUj5uTb3CeeO/vKKoqqjjRog53sSkfP
m/JQcbY8ShK9uUkzPgK+lzWjnBrj07+On7LTZj2s73HJb7QpJiBWl140ma2o1Nae
/T5txNGqGoO9yvcsp4KHzgwGxptGXzFM0z9pu5H5QDwLsD1HP0YXICBfBvC5ELzf
wX2GsFzsP8kxvGueXAsNJPfTFozdR4IKxstQNzh/7IkFPIvFzn2h35j0Cxj0eMAx
Z9BTxXvZH48qBLi2ROJ+TZ8UYc9olwGfBtR0nbWKZeKJCoHD0M7uHU6PFDIiQnkP
ptQ9ja6oewYxGKsoDyfhLokbqJD+s2nGZxGiVmbMEQ3jPu1X9Yi9oHJxsEe0PlX3
qDcfc6Fg22Py/mFr01K2gtcimtsAw42fuxKgbTCb36RTh7jRwG3qI7pb0Qy2gn0q
7q/AaTCl76bXpV5ZGTHw0DDreNHjfLQAkIa9AoWT5U2sHXF91RcxFXSmjLpji27h
Z/Xc4BTpmcw4XmDeN3d3wAsQpPT8grMx0Mg9ZdrzQj6f4FgYH8vceNu8OJ5Vb4qy
AW48WhGoSr7DoL50bzUwS0obSfg4VkLw3RMTauaNpo9qnmCGlVujk6Oo524ExExF
5B6fCyoGeNfJDpeIVKh9aBbonW+0G9XmFzIsLXkYjLCA2aLb7+qfMeziXEzeiGFe
g5Zf6IXcNA8ld6V/qRZoyUv7Yac5J1QH8BABUHQ3SHK9tdl+ZB62DALKMoOLtSuI
hAnx9S9xI7t30TvhfjWwEswFgwUmexQABdBtHKmWn2+fgW1dvMoD8/+PvyzQvXcP
E6dX1u++HOLoUrC5yTo9mnoYAgDdBu6iU6ArcDlGc5AFp7ooWDzeDL8OdHRCDTk8
9l+Y2dxfhPwF955kTBr5pPAzV/MEA1+YPZB4PbuxlOnUrXK2IKG9Ue1+Yu4icvOp
t73DRQtA3TV4ofk7SrfoBoCnA8ZJttJlNy8NgaBoETc+O4yBs6f0PIWShm1xw1dP
PO+Ek2du6OKk5xOH9VSf2BWFzcZcZ31nntD+a7SZvxnQyD1v5DD3JGhnwpBXr09i
rC2nG39qczYdsHWABT7/OCVu7nyOFOiEzxCs+RW2uypunriLBfX1qD7xrGS9fMmH
8Ov1hGD14fZSD21vqYVGZvOnf3uW+rIlkh7FHTMbeYPhvWa5EpNJJavQ8FoIRBOI
jNtr/QvSQEqCyHKd0YHYxZRjjBhadmLN9/ELOs+3zYb8YLYizjalHJOutCqVooJX
BFTHPXPkPRfJTJTlhT0Fbr1Im32sYPFRvfYSAqo4eITHMytPjAS0czQOGW+VNvpx
G1Mmq40NLQNvIZwmfd1SFWe423IKO4GuIPug/lqtB98qbUqjPTSFaCzgeVwwdgXS
rljQy6LvuiQ2eOTqCHTWziRtNw2vTrONLXxWxWbGSeCI8L5QR5iacOpzmx6kjthY
Ti4CcNsxduVyT7ZT68VTT2c3Ts/KeCd7IsL5kz7cAbfYYjw+MK27kSV2h7E6TwH9
77CPtM4InjhaEAMt6p2gjjpZWUuKGQS3u2OeAC+tawg3NWuDy3gj1n/q2c2FSl0U
P2yoTy6CQ1sMuqNnwxeAV2i6ZMz9MdLT8aV7FwhRPJ2mloMEgkhqwBTF4JMUoIgR
yINHF7WRYp48kBL5GgRvftINFP+4DjZNnJFcKqI4GeuIuy8hlb4UQdD21/fjH3gs
zNlr4s1Boz5x5OLaMnLpOYut26w3s1y4ElSISqSTP7DMDjcM0KvXlsPKYrFP+kyo
rk8dQ9KymBkg55l36x49aLpnZXfbZA4MCSUlwiZo+ccstqcquwx/bx43Ah3nqMdv
qiQ3F65/mKngvEcfy37n/hJ4M0fISoc3w51saryqkzw7nBTB7opR4ytwMX1mKrNp
3xEa/ZZ19g7K/zWmr9lITmHHsvAmVxgOu0YkV+0KI87DTGeZwGtuIvrSwQ++AsEp
mmAZSHTldAKouktkxldc9cK7z5DUunqKnxx5aYb7GfOQd9HCGAI6apTMwdaEITAZ
7OCJahvFMkp+z1KmGFh8crPvTLJ6xoKVb6IKSOjFD7265LULWxi6a6QnMfl1TXwx
4CUfG+ovkQBeatr4leUNkS6m5QzLIIgO/nRZnRcSVm0c4hvV2JoztAv4AFcuaZM8
KYH1+T8YFYk+5Ht40qycUyVi389Lv1sMyVEvcMnpn1FFzAFmM3c1QWUOkTDe7aXX
V0daxub9wnBp4XJYtDvVKPi5D7Qf2Iw6UiLsOCwVQNGQu4AyHU3KQ2BFPLGJeTTZ
8udeWOWiss/c8oiKFrgjTOyvwWrFtmUKbK0npt+IhcisxQZrMbO0civIKJ8J04sy
SFkOX5TvcrjkxsYpcdnWHuYYc2pKVXcrvv3Av+t9Ml5e1cvubvB5jqICfhP7g9XW
YGuVi5Wal1XKM5OykJxNzsfj4YOTPJ8wumvJ97qfAYyZbUEE1z1Tpfv4jvZuCwRD
D4FRVAyrNRHu/YhW+R0KYHowf8ykbR8Ar0ZlEbEjjq8dXs30FZcjdgXRZZPYr5ij
Zx8Hrz5lpFh1cK71tF1esBmy6M3zRPlwcGpwWBPxUgbfak04VB1n2t1YUMaW85yu
Yl3FUU0jELgNBjDyYkO4wJ4Ch3e4JKmgpSwGAaXMGBg/J8OsnSPm+RbTu3a8ZDui
lOKABbQfaEtFixK4fgGbh/7Yqyl/LrjUtJXJTcI5ROnNnT57V1fhKBSmFh916w6u
BtjOucu6JUtHBCVNH885coROwRC+s3ZULrlvWg57q+BgeMIPovWpOPII+35weUBm
UplUCxGME+0U1gT7mnGFABZl+yRxh1Mm+WXefEJI8cukUz+FdaNVi/ACMiEs8oPx
DWq4LqxQb/MJlJtHbDLoYCFUA/StE+/dYSpMAn/uKzysbvBQ0JUWYchepYLu3IdH
Kl633ol9XNk04/lX/+k7JdKfu0aS+Oelsou2DkTOAZuEIpcFf9wj+oE1Am3Gv6ue
Llxj8jWWK55ll/mM2UcYzxPIf6t/EeAysLiO44Jr+6z8xALwlcZPjfwrbP/FLomg
GnRf/tJ6r6OaC8ifK2hIycFSxNJnCRWJHBGAqIZlmJ412Yt8ELKTjDEldYlVzJ+U
0uCad6K8YX3xCncghkZiCpvG1NEHR/9WE0ucSt3h9QhsXkkUFz72cpDULEneRNpN
w4s0pCFb/cn3RjyqT6qiKf5/Or4VXBSUFIWGBfI5UCB4TQV/sDhMWYeGSbuazbTm
Xtdksiko+n94eJK2crW1DrJjTeSCR1G/av176t91xkI6wS2jXWEmMZPXQ4EqyiRa
DRKOcOnRu8bzh4qQ1eSLF3zfirArjyqWVkzf5Hm8QB/MIGo0re/yB0QbTnV8b3mF
abBbgIG4H/7OI6vJPdVoDs5sLPKMjZCzR6zLNFoE5QFO9W9Qj7dQe8IaGoQA+gSY
MC/M28Q3sBMswPmiQ0MniOsqZbTA8t7mqwebuUCZkJtuqcYxqx8D9dw5nGIlzOK5
QQJFdPMpVLQDvOFII3xFGeWcVRZf2VUv2wz1uYtTnY8IhNxuQ8ruxSHaYPJ57Wr3
pGShWtK6pNytWp6BlKSAdGXzj++wOaUvdDhZiluHHch2fHvDrm4m3yTxSvUs19s0
wco7CgEv39IbdsO0HaAWA0yKmGon9udt0OZ2/eKELhXDIMYqD9nYR1ZMKsv3aula
lQhNPKDlMufISDPbrY9xDmojSC9QgiqgA7iHMs5bhD1V0w4q+EF2C5ybBnI0X3PT
5Xsupoq/NNz3/bEdsBacdCJxVJVDVkglBwIb58oewMYP3Tp6ZmqXmP1voroKcRhv
WNlfswtmce6Ljm9Aq8cv5X90EuvuR93YOGRybJ7Y7LbgE+nlXaojP4pfinendhfx
UJD8r/dCxA4fo62L8i7kDazEoznzhAYFoSu+EAGgb/MKZcCFEYtgMCs3qjFWaMkr
21lWGgmJPIVH7wGn9JBkeA+sN+JK9YqzQQnEsy2HaaGBs53Wv01ncLioYfkRSbLU
Ya2juOQLcLuDKZ4X++AfrpeWQxqnavqZ+er5cFzyFo7zS3yZGa/8qdSeHOUH4Xnf
jqG5oOiw1fk2MxzVhL7u9VHhtmafOvxsBjZmZIXTL5pe/1x/Ea8Q7aJPp/Yrzovr
0Y1ei3/mWwcrk+/tBer0mSRxpAX+cKSuLYEl4rsCULPfvRwH97rnWjVLf6L+J6il
oYPGpg4N9Z+Mn3Pv3stwI9nF+3vodiKLZvi24vGZ96bSCj6a+b9mrY22pm9CaxoF
sklvRgzqV4thCJUfR/UpzO+HMFNW6wqtwU14S25bB5nws2bdymBmqLFAJBmEKLi/
jaY9eSEsQH9WDSE0IcTCW5WOz8qm5sINrQYdFrdQMAe4SJZUfm1V968KHt2zVMPg
iwgQy6zh1LTcZ+ChPb05kAJ612CBBlGLsWpetoTbXGeei10OCzOq2i4qpSVbWegS
vXu5SLkpXb6qSV3x2UGYVOG2tyhNpfMCM+ZoFYAln+Chy+vzDaSwUIjwGyTLLlBU
XpnfEWuOmpOk3ie4p/Nkb9WFfmP3iPPVwvakiZzHd/DM9NZjXGDxYn4wLXO5Uudl
4FdPctO6D2VVqzwN51ZsAlq+4Zwi1HUHO6vtvjSeyWdEm/AWXYpISmW++H1RfWM3
iWyaisvGtn0xZYXYtAoVS2ULaOSRaLU083CiQn4qAkdHXwT9TTSk/yKs02zrQZFa
2yitNaktFKRoFPZSee1BYtSaP3+qSeulS405Obfs1WWDGzzmRuobs8NvmnC/bseh
rZ/Khn+gm0kCGPg53ikuNiECnyTbu4MPNnvZ28tzfWOirDTm7w+eirip7r1+LrYz
41Hjc/kJwbdDM3TqQxh5QrHX3oT+Now4mo+yPBRglm8eA7iDLJ2e7LAuyR1OpTPX
/8vY13XGkYmHSwzacnpV7Y9ywVCAEDlCBkdo7WssCW6Rs6YFP5BcpB8cRTGQOoFI
/kOZB95nyg7+jRngTFvVo4HtHAMzHbIfgWtAr5PLjkLewS9FfHhbiwtTgNUOprcv
OY61TaMEV4DIPaY4DuH2ebJ5fq0P8tDG4B6mDN9rht6HF5rKQpNa0OZebGBOoMAj
mqiXPUgCIO/KQvQwBwHK/LUPlyKvRysUNc9MvnNirR73HvdAOg4/h95ORghRVRvI
T9yBcPO5iIN9qDrokgnGnk4GpNVqhlltrq54W+nlg9lpA7VF1HMuWGCVPGf4NM3V
h9/MLUn+h69mX81U1LHC1H+nM/n7+HCVflgOBZjMpXskAK9rqWk79R9JnrjGjmCd
xKCgXTMewpPojWigeL4zd/N/KAYymhphYccWlAxWrGgOQurHvMM92UFqpfPTd5nU
B474ADtEZaCQHXt8BxqFzn0+eedoCG18lbwW/FLBsYU1AUI84VIp/C4Jr8dO67QV
qL6PeexcrQarBDmqRLLszZHeRNwbTV+UC/Aif2uoqAxTK7HCBNjhBKNPMAqbIvMh
XVEp6IdelXEJlxBkBA8IQjxji9cMWrCZRpye1OJUjiDijqYhvZbFQKV5lQ9n5ZU2
MqHsjEvoC+RmzYT0noi2GAhjBb3axUs73Xbo8dOgt1v3hfnNZ/VLtAf8muZzqynI
oLfbL7Xr8cypnblKd+aOgf/xRpgmC1hdSUYShdPXvFzijijTi19RrdTUH/GxyhzA
NIxfgNAw0FU3yUIe17GpSQe9N6WG6t7CCnv3MyEyjILz3apXRXvmSqisDs8Qh8IG
qhXoVgSrhqv2B+7K4bChihlnyjrGKcu+X82N/Dg8+NSubgGLQgIAip/mAptT9iw2
za9ezfmis1j48bsK/iY8FpshwnJQHUBzB/d+BrDmwbykRCEnrR1G6qMtz92YE735
dY0/DrRYoak5lRUFO2ojhH5fTP+t5XpDuBK4Oq41mBJlr+Xzxk1FoyzXpToo9qB7
B858adqiAzpc425qOmsJ4aPjhQKhfSjBwIeMrNEkWBmuKWwOBtYXK0X2Z3dywKz/
AmUU3FSdvbmYW75r4ISRTniLRqatBp4O65yHQlfhiDsCoi3hgMsVdEoVpb4f9Z8Z
HJk6L6olDaziStH5hrmf5JP59iOf0R1rQxrN2SD5bAMiyFHSPlS7lpHAO0sZJiuE
WJQpBYYnR7FsGwy1xGAARiWX/v8LrzY4zP2AxG1xEhfC5cZ5ylk6uO0c6LAqsczD
iXGNAKTb0jiQoctrCdAPR7aMFZHspsNt6bQXrv5s0R9rQOm4WzwR3O9alosHbtM3
96jktx33iQmfFccLgIixfndzYV8sVJd51rjEyTRPqf/+MaAm/xEcfPxd1dSOqQVM
YjWhtiIkvkfXn67DRiFygumFin87LnPBdS9p1whuxjaSx/fVUF+zUTHWBZL7Qa+3
5blCDNDaUhKcahjqyj/ZCtuM5mBy/YXiUReokCcbKyJ3MvNgcTX+UiPehl/6j2FQ
qTfRmw2gaOLmZ125ZPb1uBjFGiwADHRi3PyFFO5QV6BCykkcbVNQHbvSp9uZMhAI
5d/rjTtdhlWqZUBCdoBsbvDn+1lA3In+A++MMvjf53Px4TTDgbMVHMxhOSN2s/Dc
N4ynomgq8//WTdFnhwcVc5xF323rXsWpkzxvb6u5M8USmGGsJboBt9MQs8mMv4ES
xAtwdcKnM+YsHTaCKOhd+HfrGzfoyKo7xwElSRHKnWyiREb4HHw+XtZnu/zkA4jX
mgRLsunJP5QAOUscLKC1ypNCOcYUoRGi5loo9iK50/bVftrk4GqX0C3ZSx0ft8k/
jud81imO1jTU42KnoUurYVdftx9grr9Zktwd7h9FvF4bkiWmJ6sLnT2tq2ClqQVK
LJVvtpf+JES3Cu1JBYsC14tIEuGkfyvmpPlPrjzT6UoP35DQdgigGx/UePm7m3jN
eOFjlqMwqPem56sD0HRhYOjZVPm6C7cO44f/OVo4l8r2pgHBd1c575k+0TCwT86i
yplMDq7R/+h3PgRK3rg4RNY+2Mi/6WJJYK6ShkWp6H1UK8ZiR0bQpx1rYDhDpgIK
WRrRxiwxZDOSMiVpSu5GKwGKNYzc6vHOnW9pGbDj1hGwUBYZNW9KMZMLic0sspl6
05yIy9xpheDvSRxdxGPjgLUzQS+cNSICrpnuUTl332yTLRaLGtUMWQHkLjiugQyM
/1mTHPHK9XfdOQWgWVOyixVWjUgGYbcp1VOsKF+QYFt++Tb6UF8i+wusWGsnMeaK
6PJT9vLJ4bjMsn4Drlyps9qrpzU3imoextDF0KaYlHoucwWBko9WULPDOxsSeTAA
XQtVqcOC9vN1HxnKcNIAO03w3YkOI6L79hFxB0WIf/B/zYHo3AcwMKe/cam+DHWD
FOLkXUERhC3jU59fjPdlyNdhRPSNnx9E4Sess4DQoJStcTCXXN+ClpC+4zAFMhZr
faEzTutVfAftE49MJ9gW7WkC7mVA8rPhlr4d323LhRg5/VqsKAcOAcQl060iLv/D
z7anwRtb70tA/iZIQDpFPA2FxaGCPc28uQSK9sZx5O3168OBPaEURUTdkwDbCGgA
IrTlwhrmoRSUqiGkhhJzDfi+cNt42820KMSl3TOSWmCxiKh1+DImdsxXpOENtsLn
ynKCP8eCWVS2mi7VTBHdyKi5wzNgF1POjaTK98CKjHzP5o8TYTXiX1sLmlZJn3i+
84n7uFTOJWq8Gn3H9Bpc2Sk8ewdVkhMXZtUqohGLMvLtxL+MWDg+tBMUW2fdMzTL
+64boF6B61aPP98m2urx0HlGWOc8Rl2wNEgxE4aADeuhyPEYUI+jxSRpAvktPN/Q
lIo1lYkkfbzZEpK8ZxzEGqLAXPQC/euBkDZPoDV/0CbTP1PBukJzJySJ8MCOPUY0
mve9rtqi15vVMKwh6RD8aJMxvVpJy+Xmz5yNu2GKA4Bj5B/Z4og4jUNtQMbt4967
dG9VPwaDfclK/J4Xgm3ApHvKyRYMLZBOGs80fszHPU6L9m9Tt8t/W92YLd5kQgrZ
ELEuQ4cQyJDJa82FxXG+WSqNt+lLcvVM9A/h43L8Pq3/MhcEOJj48/cPPgiP955k
EFPjOwHyy+kBslN4ydw4kmv3uk+09r+wqKNHblOfcfYSg/9sgFH0QtCCmpu4n2V3
YtC0uT5EDMcnLoKkFveQzuPDDAWzgOYNPR+1Je0CM6pMaTsU6dTMy3bX3YiLMK7W
K5GjKSdYIuL9FWWzRTQm+GrJz09Cp0Ne60b6Xnk9kfG5L376nAC9yoVh1EHa3iIK
gd0HmH7qNQXVfYsRhpClc4efPVJu1z+tnq49Y+tYJGb1JBlq3w/dvCk7JsIAVdIi
b6ZIk53StTjZnYPOmV8zsYl4nqO1mxPTKDiNm+gSxtjiQ4D7SAx2Fj8SA6Ikq/nm
D+1wxMcwJ83y1V/g1052yJTiC1H66Ml3a0x9Q4081pYspp4hXpy38K9V0/vDETNQ
cPseXWuzxL7JYbJG2oLo5IcW0fjCnFhQmZJHFxvWF57TzAkxUhGOBy55jIO3+t/h
FagxbWvmNjMLL/1VaPLjHP713Ty+gU4seXbyL/xyjzfu8HLAuZwEfs5MSWR83JAt
4GXW/II593KoWJMUqVacbJTFwA2/ke/lglhG2NYDgZDABREG6GqFckbUnaozoty5
6JuIBTFUNdL1O0+wobYzuf44MoPmps9ZM4tyykr2WBbAyfrsZBNaFQzTPDOQDW/m
x59xap7uh3/jXdXUHeGDo7bMzP0Cye0YSF08pCpLyi6pWEnZqw5/Zjke3D5vjhAj
oF4n1G3OIDykaFyRd5tE5N6NcvK8VtxDINB3TRDPSl+PWMXkShnN5FEQRa/sPx5k
w+a7c6dxK6lqyjggt2kil3Lcrdfj/he/VTAtYZBAO4raCSPt37CtVRGCqiwraH/W
/Q1V/T5B+ByzPuu/8EsFJs1fCabh4ZRXYqvvu0SpYu+o2u9s08+WKu9oWLHzttaA
5MwtX9xp2hy5VeSitaG0YBcWfm1v8CvZBuvkTWbIarcN+OY7/f1gJslcNkiml3cc
SHdxd2pX+2aoqwX4Gg3sChWEIpGK3fyzwN0AkXsSKNFpzm47fz+WIlb4+X0Thp6u
LM2z15KgXDk+0GYxKcJ+dTtxiQNeVoRH2PEejZ6RI08kv2grmuuMGyHNHEaatPzg
T4nTiiMGAmjsNKT7Or/hwWBdsog06t4PVG0OoATe+ENzQ0r4zq9J5cv0AeKvb1Uo
rqZ/dYO/d0rnCBy3Qcx67Hmu/DAqnTeHsyphD/izp8bY+xZFqkVWDPHPTcMpADmw
EqibkaFkFL8Cwzc8Th7gi8OpDoUfqs7nIiNDq/sAPrb6nMDf8ZR3rh0bFyxPhV4E
4jRhi/Mm9sb/ThgcMRPDPKdbLrnkbcXufJHeRoQAs3iPCJdbSgsYD4kf6mI7TR7R
QLzmCO1Lhbn6ae6Vz4oCesH+13UUWABqJQ4eUe6/Qn++wIA+Cxi4KiPbJFh2E7OJ
njV3K5Nx4xnacTvBRRVZxmQAkuQ211YlV09pUOSHRUJdegRtVh8ZE4buwg3S1Zn4
9JJ7JSxUPdx/ZlccPJgVlQSSibUvprK3LCI7eQgdku+oz6etvrhWgmyrKuwAdnsx
ZUxpxvyc/iB7ey7Iqxt0HIEz2929/8bRQpF3pLhXqAuv4d3aGlFh9mK4CCCEq00f
/bkjJG0F7oPLEuvN+IhHQ4O8yGuHSz+NSPjlldes6BLfqwxPTXlFvntyGZ3dXGSA
8xgjdsqJypJtwp0yKrRE2NXzkifw4aXgoPDCtAYyIJr97zUSVPS5FneluL38iv7R
5y+W0dYt2CW3thy2Zh8HHzpR8VsvXYYWSHwPLK2DXxx0AjeQhQAWKx4/PDk3iWOA
htnb8BzQKhYPFQ5ZLxV15NEtUxW1Xq6ADFS7L6S9CHq8F6SH6RZJ+dR6b9KS6ZU4
KjD9kp6AFwdfUU2W1eOBE0CkK6sZgCFum0DwSlKALmxmTaV2VnyIdTiEB85moMBI
9/L637EiC81n4mEtwztUSxdfbnomWi2H3uTSpVde/hycqzZ3H6Is1AzVtBfGM9/P
ouL03LBLpNdU/GIpjJgMRO0dGNS0m3VGikpQkyU/zxZRCq5O8NB8a1oBtfe1qY7R
9sdM5NnZGbr55lJyLIS/htSpQ2h3EpnHfcZBPDmisaQ7UeMJmnsD2+Mp9rCGh/hx
6lVlky1dKO8g/T4zQag0/tf3fgpvLtlW74jQJCUYhhUj3S4geZGBcVnByvNa5145
sJHEcVvCQ8ouPIVnV5btLSb32vWXaiswNLQ4oQXNQjCmol1sQ1FJuqrdivEMhojM
Mt01tBjMZ5tPM16lCBOfAgIkGdF2JFnccKQouyS2kXKfvFKvbaxI381dGc9oLU4b
zIx5JsHP8sunXmjVt5rT3xd7CvM4UxwNNxicuVUA/r81Xz0NZs5yg4rrMRrFQ4NF
HOLSqDZZANABkyGfpyQPgQPnNWuDZ2VR70dcyFvUKVIwtC6W08idgzgqa6A5I4ML
n4XLggoZ2RjptmK1ZSo8+Ia6K5WGjNOZnJagxUzWw8vMfPIKakaLe17fstwBUSZS
sUeCdJrxXGFgZmWfYic29dpc8OHvefD8tpuzf7tJIt90RYqbD3BLRqgDTfdIRAis
DKb6mpRI5cnftKKomaSRT65StBu4gOhTHI5ibB24cEusiK1twPpq2tCiB7zHOZ34
O9TPuajLWFKzCXQEFU1sRZinRYMUyD6fl+hVifcmgQ0PCGxPGPly+MtVaUtlm+CB
nJD1zY2eEQX8ocytciBthUmyIrlwxbzI1dfePCMqdWPpaf+EqFIr5HXL9+Maxt8R
K/2llkyKnHUp4iGNxV7bHdFxc3PjYX2ozVtS/v6Ew6EFRCxdAbx5QjyOBu6LhbzL
WhYaJTWICItoQdou3vBe7JaR98ur6x9ahnTjnMa2e4IF7tKC9b0/XpBvfFzUy3Tw
37C1O/D3oTlG4Ms/zrAyMiWlgQbxOnF2sRYpm6Fc9o+9gpTuqx8SAJFOq1ilQEcp
0/qVkSm7prndcxa93san3VmgXYA2JYQzvdf5o8jN435f+0/wkm1zg9V/0CINtnBH
nnR5my6lZ+E8jtV+NNt0wEQ80K0/RJ8701ikktOOwO79oqdWFaFLGUn1s1Hw4ruC
PK4PLgzz3kupvAS7xKsPLteoEm/hGV+9gXQdWRgmKVqURrMGe7clfEOHoDw0Zozv
FqCW2+kZJHc5u9Xr+KC+oKEjJQMRu846Hb8dNuN3UcBcYjCVULZB0KinmCMa61yX
zdbRZfAq1k23w8zWqxbcZB3kW87IQ/cnLm+h+DKtItw+L6/HOHJqvd2rqdraPrdC
TkR3nwkNF1oZbSTUhyBQeix8zstHDNgOmJeSN+LEHE9XbS92sN90EWg7a/1pxK+6
WiDyE/EMUbrsxrJuQQjButR2yexrg20i+Jx3ench/mav7N0+GztJ1Ij8zItmhaCq
WaHUp2IVu63k6jf1SbT0JrJeTsuGcNVq4AcyN6o4DMyheN4rTgHX9xTb7yEhnmJd
B3/jqP2OAmfTaA3QcxxbtIQi4Ly/IFV0105zEf5h0whhD2LP205oGHOz2EJKCoEm
u8Hi0sJv163o+JpWh9I3vBLJkOZbj8ZxGaeIC/0ebmHpeIcsuuOgkqEZR2+7/vlo
REOh7OWshIPmPQzXb4NWm50O+WYXOp5qCIAvfowt4XeyRrqIU9lu1qkDbLUhJIbK
i8Zpxi3zKmNXAGcY6h6IQm44150T36nApgD1dci5EH1gp3SE9vptPxwm+t1iFiyv
AlFMkFi0wulifugUW2vXpLsjvKuB6sC5QsaAPwuT2YzNLBvDsoMg2Twm8uPcrJcV
TqEX6vN46N4FEEX53urRmT/6XqH27bZZ/4JU8E3igUv3ScdrBqeGViI+UMxwjox3
qnVhkuKBCx1hGdmRMGIKfoVW+iFOkunp6ysTlZ1/kVUFqnzwwkjR4rPktteljdGb
4Kxlx416kojFL01Zdj7EKRPjFZvfSkueW9tc4UMhWD6dzVfEl94ochh9gvzaCLR5
9GhxmmuLlz7s9mkEvU9V2Rtka/c+rEIljLpHDpnV+WtyrYiqM+RYfvI80BCSTFEw
JKOim0G79o/o1oZhS3qx+iMCdyo2aHQimShInnK5cFLR8Ac22B3pPhCPK74HCmD0
wQ5JNLQt0bh9FMwog0bqXg6uG92fDZAev0cQOTuP1mpxQL9TXYI3/7/3Z84N7ny+
ikQUl7yDuF5wjNyxZfV9ScqyYQB/P9jm3gqacZlQzymJev/UMx5qsdA+OJiy/TxG
oCxv55Kap0x1/5hD/5R+npdOesFXTSBSUQYppnHgja6YyDCSNkmk4cELPNg3gqJx
MWCa2N4fY2vvI7SzSOTHWEoqY12MtKiCBK4zsMfm86s8b2o90aBkv4rKD94S6PIr
Vppj0toYT9KSdMVA0jSHDnX27OoQd3p5luvjFHi26RZ2G7+/vBD/Jvyknqtytcmg
2GrY+KN0TLlyp+Y5CGA0FS2leSipebCiSCX37G44KvPu9tOz62MkdEgSmDI03N9s
ucS6LCcqMjncxX+WTcKIz01LfDg1e8ANYPwHX5fGljZ+lTp242QKPZi01+uFYzcj
V/lrmELe6XYly2ybpIjyEIbTY5A4a31pqrGOmwevWEwIRtYoslDMgy53ZgGYRllK
/lf8l5WbopXfAalDJu3KJHiewPLg6CJiSTFYtQCRUBFTvBFm+Gwy76+jfskSZZ7R
YCvNs6lZik44rKZksNzBHGIar7tdG4vQWhdGpZYU1BEyNGh6O/fB/83/6g9+ylq2
Qy06JH+9uDKxkgGNQAkOv4uHTNy3haDCtkLsXxy1R9gbXuY5f3EZgxQLBOCv8KaD
fwKyOTCVxBQPvYV8NcDc4htL2DkBPQtzFkrLFEv71pqp/yLL8JLBsvEVJX/c0uMD
mDGB4dmiPmY0gTgyjOZr7a9MJhYAjlCT64z8rImj2olSvLb2p6pRxOKm36XGhpwr
ntvJOTLJeEfAtl0mYoHr1qTDj84EcJ36CWNu9K7eiB6TOrZgvz+Tnh0o7YlKEPKY
n1WoVJFTTVuFpagybFyiN+IDsrgr2deK56osVZSPUbBSHkFfVVOSNk7MyBIFe5Sx
MFFGfJLCePCMaWACflNLnqimMk+8UZ9EWRfxkS6qwTLdY38pazopNUEB4T85CdQ8
hhv9AB+Le1PQ7dDLR7nXGh6xaUgoNm6hipH0ZgVb/Gb2U4gIE0U6oZwdg2rttum+
g8GCkXem2Nmmukn27QGPuX/LDrHfohmaDX+Cmno+lgjiOSdWHqp7Xm/Emq+xaBAn
DA9qEvetKwGrN3ur9SMi9PAonIt5lV4kdjDzccXqhjRoACYKF8khVO77GQHkd24Q
Pp4ncs2vYvjedoCVHK+BWDo6UNLbKDRXWYIzF9B7W2OxDuXyafirswoY+fB4ZyeS
MZK6Ewz1fiY4upEwEKFG1DdGy0wRYTFfz8oEJh3CqMqLIynlGMegIAcsPIQ/Sl9Y
UNJDbRhry3w7IbwP4tKA7YyaxOzPidgFEgUeUDJPelzX0FR50GE+1z4tzKedEwcM
PnNaT2kT/CLwtUhHHj1IohPSxwClQkFG3umCuXts58Fj5oAP45A5Vg69eFyStdcF
1bZ50KkDriVo5hIcgrzDIRvEhPrfzc9nDF+PSBbANdqadnAgo1/0sJJTgNcrnA4w
8iGaxJc3AL2cljDYdYvIccEx8Zj3XevcDnDxd/IXJZ+ZRU9dp8qdTNhtIbvG/Y3Y
wvToZB8YOsWXa1OJCGTyndE5BQ9773MPtqIq89ixU1PIPhnRHpAIn6O2ztTrkdTE
n6GEvO2GE4g7C+r3pJVFUeILWySPVs9zoSTzoXiPlSVCUdRe7T2JcyqoO9CU1lYk
R0cuj7wCUz6SiQtV2hzzpMpYeQhbTmI7j6ifuE+pES7Mu6A+AlXxM/JKmghmJll3
6s5lvJFZS2S+hzCQ5G7/Ruq1dYxe3DF0NSgKkOhv8IedLUBsSMO1ZM7dWcsy9wPB
ykFMzhqZsGY60+8gWXS1qnUYwmFXrbQSU8xD7kxZG0zk8lCKZXYnwsd3lsSwg5cM
u7pYfSsHg3v584N9bfC1T6A1vT1k14P/Wm/aNVNmyQLrkZIoUfiCK7yIbVgXbnvu
bSg4AuuSKKuv7aVGagOs7vIUU14l6Ps9SQHWFuKQt8DpNNZ/SiRHw37m5c2GYDL4
sPbp62qNN3SDU43bRX3Mj1REzGkdaZGuX6PQAliQFF3Fu9oJ+oJTGt6Yc8j8WlgH
zY0DshmwEyE9WJ9q02Mkdi/JuPe+NBmKPppp9AOU7rIg4dCIMH4CgIV6LG+Mupre
j3uQg9EG6AsLbobhPSUvkpdG+RtvVcyLHUgw5ZLgegqRUygXSH4hNz6SHNx+je8+
ldhiVTHlwxYS6Orqf+79NzWHngvkiBJ5v/vUcWAvlYVGgJvFv51gUYd6P8OiSL1m
kgaqy4NADFHySDA70dT1bobDxceWSLxmPMxvxsTYUKUK2DVwSbkx2u09H7N3CKIB
jYH2l/f26DbeNOMAyThR3wPhYqk14wZSnlMOZvMTNB6l3kxFT6snlyBPzOXNpMA6
5ZhrqQ5M1Xx/+LAmbpuuRW4ZlbfZbLSD6VW99EkUjQCO41sU7kr8jVxVnZfsrCG6
2C1MiaUF/y7Jb0cnBb82rgcbE7XvaOZkeky05rftVk4MDb59lCyOfGbNlLJJ1C1x
Igxk8wqRTlr/rDcefhf9GYX/z2058MaYQemI7R8LszuztJd/JBM9eW2sK6qz1+qT
Bizupb+JQLGpngLeUbMZ+eHChVKtwFL75Xgf2PUVRon7DLEzyWsFI98gAMJeLb+m
INhlnBrQgGt5VyYEfbJq/aOq/AQIqyAZ+7Jda5KTR+VNPsqr0cHzugwuU9kHbZHJ
T1wfKFsPtNr0MnhyjwwNWgA+egUT9PZTcFKjWnK8e0IkYhWKOFJ8UiCmPBZsOU3+
kILw5L/BN12Waerh81WByntrzyYQ/DqlWldmtU2UL9inUdtn2UA7BjMNZfN9c4rI
FWad9qOqgp18rkbcw3OxsG3aF61KMpR4PQnphUaZpTAHBxgaMr/vFtbFgtzF7q64
vhoT9RZjZtoVMtv2/e0XoFvhb14i84YvoE6fS5aNT9jL2hETDH1QR5wRTHom5RmL
Bu/hTdSLxZnDYIDXpv4LqqNqXJ86X81fWhZ7waLitUkumISBTxHAiSMef/SD6nNb
csNt+uTqWOvHx6j8+ALEDg2HghnY4FDCDBKfOo4YN5xNRhWgNXL4vdGL+L300d7Z
C2ss2Cz7YLy7hTL7jmnouiTd6XPcIfb1TRwo+GGZldObHuxat6+wrYSNMyAdX8yL
pCjCmWDY1hMYeH5hpRYHLc3593Ul8OLif27jQJd+EkeMpwt9WLleb4ZdSxipQSmj
TYLGhF3+u68o74187rif7UxNkUGpf4f+DH6d+80axbIyqZm5tqHEk4BkcsXivL2G
Mq80yGTn3ENVFPdEEsXx3DfTJQOoCMjHewqwBihkz2K6tB9qugth+I+S/+x7koiJ
L9bP195AMnsU3Z60FPftbm8J837LQtT9UvnGzvc9kdxD9a4+pAKfNUFcY2cakK2j
qVNWTHBCbTdZp5anc3QbyVlR0ulZEOF/EAT3EKXoOkrdh4GL7Xfn0qPex+p2xhyH
fEvDi66iydALbXmLF7U51UmJjircDwsnT1jVNLxbIi92UewMH745WWnkviWk9W+a
UIupR1tsr7r7q0dTBu+mn8ti42Xf3tiQVEHtLdsFC9JJ5zmU9QS8FEj3y69J40hl
oAcYf6e3+BSiM3RM6T9wgQZj2xpTfMbrckL9j1Ap6gmWsgSvl6GdSz7NQUhJZ6U0
npTywqLrCx8rZ7eMRXZ11VNJN9r7IaTZRPNmgBN7uihmCB+wagtQXv79L7VrbZjD
7HBRN/u6VLUVqxlulxo4cOgDGWC1H2akdT4/LK/omvmuPmruDa1f6NV3y13z+PYU
at8cYf5qMsMtB130xsrnwo0z4JlljnVraJhxqEKkNRisHijUT3vd1c8YGlopWZoe
jCNqqDoDkjLrAWyWagIc5tDshzyviz+acckVbiBZIP66WOTm4Ne+1oFV/pZq0Unn
te7dqokynrraponhMuuIBcyvDOkMOHCUmjLkpq+O5cctOd5vi9cpzOAeGXDZhtVl
0VQ7KyOOZts1iuElj9ltGUPhrrpwu6432qOKVc+XMbsgXAWnmOeD7M96jC4pu9FI
3RegPaScQKXEZ8i4+XIYcEWp5G30bbDKmUWaoiSB0owJEa0u2JSPRIH+vLYrqAnm
lbUoyJYmPRPvZr417VX20FT3rETGjK3Thr7qEh4A5O0oP5ikFKkar1dMDriAtr7h
hoCMM6d1f3gPuszgSMG1n2SdnFuP93Kv5IBjSwVpzf0Td5sVM9fnH48W7w4fSu7u
U6GfODh6yogYbLBWQh/Y9o9W6LiJhr2VUy8WhSmYK9c/m5KKZy2ijAXrNS+ui/Sm
9Q5OWVOA9uW1KdOc8oS8Q21nR1LHQTOes9JCqFL7/oRMkVrhFiVtZrml8n9B7lK/
e0zyrHHieA4oRtJFo1B6nAS/P9DkDgykueLHNc7TBlsR5ur91ipIBNy/3c5SyRPx
dPw7ecTtOgrZJa+BdA5eG5wG3CpKd2phsgVaMfcTpjSdWOfAe2UGc+at6YW/PsoV
lU24FiK/9/GwsjY0mTuHUu/H6fEBD3NcxqrZTbBXO1/EfKCOm+naRXOI7zXotHO7
xjaFgU9Tn1Sf3fPnFJ/AXSqDuCwC7kh9DxQCOqErIoFOXbpJwkg8A+It45GafLD6
YBUQEyCsr2/EwHd9evcu/vC4DgaWtGaBq2OHBGZ3qlxCb2WoqPjD7Eq45j9Gg/f7
6FyxKNWDETb8yZGXwKNfto4d/f5SRzIWmEAGsWm1pLW9rzlEzBYOgH1aP9DXaF0c
jhLPpPu1WXsmSEWmz1bMgYJCRWp4+6s1RSeF5MhoJ7JX1v1L8ssH15TiyanISNeq
O8bbMlr5AA6ZvJtjag6bv4qa9zcY1oG7LoLIzq/xXSBoeBaFOld7almG3If2q7dQ
EHMcuJo9qz+qExR+d92IS3IS0fRPu1RHSSKYmesDxDdCJRobS+1bsfMh1YQG838E
/dOlTMvcF53EhheT8ssDPreHKa9DyMtSY08ls3a1TcVPBEQe9L+HNeYPX3wqFrNh
NISZP+mdr3jvaUk75B4ejxg1NLAxb9p7shUHTPacvKNM1/EqFzVLW1OZCI6ut/DU
BgsEpGGOWKiY6qTlH3PMz9ribpGbcdR/5pI+StiaqAEsNcSRiGFASrdNWGht+gl/
JBvCKEhn2AQjUIXwb/AyoQiIcOlfqtD29A6nJOHyfLyoVGi2AJvL+bpiq/4N6JAT
W2+/lEprv3KHwMuH3F7si8IbGJ8zsMUJNkdxW9v2EUjxNuZDY8Gl1ryU21nVNfL9
ySOKsdrOu+E8H5M9yLX66ZEchMsSg4zAXE5OSGr9ZqhVFlm90lNcLXo1mfypQhO2
sJ/FJ5s9ks0Kkm0UsZ8ROpsxn5Uy8TzrSMz0GqwnpSMH8Kb74Dkj70YB5vz9e9QQ
P0rt3VO2q8R5fQ4J6oS/6UNcARhYDIblFjiHOzaFf1mR29fzrlAUa6MRmhbJ61YG
QSsHPUgR3n1VSl2MQ8RtwKPVd0PNXr9LAJLOW6LuaCa4dNsG3BbYkj+qwgZoy1xh
8EWsBSQ7is7ALjPEQ0W4kWrTzMJv7gKSW/4FZphdOYOPVdryghgKptsxEK6eYA5q
FevCKf1z6uepJ/FHIF+gMIFkc80Xk9EDriwRuIjV0OcjCnXDGsqeq7xEAxLfe+di
w2v569rAJiofISFNDhnlKSKeGZK1RM9SiN81yZMpRsZrjjOpiWEHEzMGUsymNYED
UvKw+MWEljV7Qc4JleauwJN/WeiLd8sOMzFuwMR8zl8jDymWJS6AfmiG68mR0LJM
v2rEFhCdk/x6LWoB5NDT0QKdr6i4V+N0TmQyDpKBCrCy7INlvIr35QADZISd4+fC
MAjSNbCqBeNbjXE8o3t/sY9GQ1tn8nZiHJkw1eCmFka5XG+Pq5SNR0qtUGot3gL+
a+4dnOC5gKXCExmdPtvrzit1lhHUg58ER0URcJGRlw67GdtoKmnWNNf8yPa8I8d9
oTz9OlIUtVyqiy6EoMsaD7ohCTN6GYBxY2qA+k5QJ52LQPXRQvzO2562s0b0euhK
gVi6ok35Go5lCRYQ/OjiUvlfPsebUQyWtbw4cqiZ1dT2a2+kTXDxYNr5k+O9cYW8
DCDdr5c8ygrvfY5tAyZIiQjw/ggNHWrcWu8otpm1Vs8A3vsf3w7cWOuBYscO3T45
SbAmZp4XkSxsxP9426VEZaXRX8LJsjYfqc+orX6IckN9hrybzaEMAqp+BhVkhPQj
ktmmy7lfCUrAko3iudyOtuHAeUEUHE8VQ08Gj4zXyg4mXpYX6zn3Ml+gsgdm5cpJ
zSVnKa+aVZbnEUmXOsfMHYzxQ0rxY3WfGLwAQQHGgpwEXuAWiryueW+Yl42JAFjc
rCRgwK0iBuKJ7a5/5ozR7qBoa/GpScfYRRYyPlvvacNqktgobp5FSbEnmwAvzRU/
F2A1VV46bbQIVJWzdyOBKHz1VTwkihv4q0D+BnIxhasX9TbImMauciJ6TXFoui5i
y4mqf5eTGYDIPAeTYMTL91i/4dQUp+5+jLMNwMvvAnYWqFnNIqI3s7JzwcM1sv8Q
8t6qjegAoxyIZxEtC7ITqoFk9wD4YcKccSxEniDSif3tudWFkB/+zujg0Ex2xTet
cgfNlLZM0DyLa0zulITO3S6wWiQrmgL+Uy/iSm554C+fZ3vyCnxN0bnXu8+TlP9f
xUFetUlFPTjNCUbDrg3IHJyN6qYuidjFNRVWaWKZTUuAHUhyMctyz5VVei8bZR5v
8bh8Hn68qVbvLTIQvrhyNEZjDyg3vXYLy08eY4Imma9ezWiTG1xfFVQNDygTO+QW
1LzezSJvK+3oS5OGLIOlHkj3dM/JQ0FPmXTom4fcifCSdm8dLoJ2pIBnnG6R/rcu
+0PDJicttZ7OrmrgICuhlqhfctVeg7yuyx4PnAm2MkMQ9ShQXqKPR3xxa0Ena2sw
zZp8PcvcSRYZ9nHRESRHKh+C/1skSKp7Tl5nripH9AJDmuXEx+l8Dg0hmJ8Ddnyy
2Y0UORZZBwq1urxQEWK20mgUTU/ofXhgj3+jKFkpmAG/VCfd/01JH5AcVjcSB79e
6hd07f4bJ5Rpvu/DwPDAgBHnD4lETsZLg7u27M26Zc57peJjMgiC+EN+mu+RQG0F
l6F/aeiBpXBTDkYnRTT1kPjebSfIomAElKenSr8JxLC/j+wNROqoeZsWFCNzuG6P
dpHxvvzHzGS3/R2fFGgE6HMuVMK47GYqeG/pU6SKnbP7pZ+zkXezEVXgqIImZlOH
hkZ4zJlaL3lMIHNLXe2ZBMcxJj7kDzDPUmJGEeW0R8z0aKOzy/S3/dZ83vVreYPN
fQ/6SMK8Z12B4ynQgR1vbku1QCiZBg4tf8T3vw7fB8xgd3tYDze+T2bZUq9LaJIZ
xp9SiK0WhN9pKcpHEgEew5ZVsDkQ0r71bJz8c5mF+XBeBXniIbF3V2h5rccIF/Hv
rJ9lMYZ5x57WhNBFddA7BQMsWjxsidiNFbsNiH+8SNs07sJ2IbJccBuimc1j4CEU
dKzz7KpXF7gUqr9m9PDH9VBTNkjQEH85HGig6lEjdufj7EZOf4V9R/zkK+QP+fSH
h3cz86e6iowuKkOnMBylpfBk9BPeXYwgvHk9rRsJRBziRIJ443CXDwPsEK7VwNgW
aslalE/XrwAVFUQsuYISKOy3iF6Jwj0JhvWWpLrzD5BC3YnlApAmSwtov6Cl/ZDm
sgZJs1+0PWoH5TPytCZmI7BDfYSkQBJhPEboLZRn2JPei3mgw6E+Ob8tNrSpwRTV
FVpGPxLqoIjyj8GvgGBe+AYQtMfgWLfEbKEx540AKu0hgJZa4MHAKStYOr9a7T1H
MhAxzJpZXfAGNLl/5q5whBQyZ2chjLbXi6c36reDaSC2rtfqiL0xLqg1m4bpbG72
En/yqWTzqrncr0MEVy2EeAXRnKCME5VatWTWovQ6nbXbSXmtJG/vvtc2Grzd/+xN
QAAfY466ZUuWqw5CS0Q3Orq6QeOBkGJGDbi7SbN5ojjVd4bsaVCBMMzMQxin0bec
m5n0hTCg6adTToG28s9CLYWZWqlWpoPNWfFw0KMqqbtxx1pyK3j1hdnd/aDDupE0
PlhNiaeWO35luSZGfBClOQ80CBBxZAORS/AaFbMjKIoynlcJab7761hiQFmQtBkq
L9qffrhpZ2VLJ1GEDgipU1GaOtvtEdn+pISQwgUM045PiHZBekV5jru8ugEIoLst
Gz6HkbYZuhd8yXk4clnEePyTkv7tULGrJwoi3p5SDEz0wDf0/k9vZRJ70kEgY0CJ
3ukgorV0LX0/dbT/p9mqP+MLFez7bBrCXD1y++72yd2ixFXz2jHqBv3J+TACFvOm
sGuKFktCmKQD4U0QDBSP8pAqPqOmeYBvKkMLmOd49cCEQf4b+r1xZ2ll17hqcKJi
x6F6SKFRKP54UU7EyUg5UBc47uaLG/vnqlXiJJHsCrN5EaB2Gi98Nydtz/BdyeOJ
Toax2rSPcoHa1pulvjfFfK4bgs+fWjGTSVVTwhazm56jF696bpTp8rJnbnkGSfkc
zgdL4Gm6xkJJD10rbt501ZAlIAsJdgZDUVuGE9x3Ua4RPYkyBUSvZpCiHLe7xoSC
W/k0C86ie453XVcqnKORxzRuONjni3syOI0+laeyA7DBKnrPmpIVwrMFjENng3/0
FDIScUt7/yRSflHlXSLKmmG1bbXAcOJTuAiHhWSpHLBWytaluAb0iS4S3rNGpg+R
bEWJL2T+IdgssIc/aCzdLqYwpZRJN+N05Qwy3M0436srLZTU9NtWrGSFAzydQY7v
tHqQyCEk6NuS5Mg67QudbjW2JthA/25vIZlfy1YVk0SqaDKRBSAqUkV1ugruHxFq
2NdYGfII7kGIu1uDMe2IPIaCXzFRlkIr/weXzbdb1WAZxkiSQVkxJD5Z/h5C68LQ
iV6WoaDxJWf1tagKhyfFOR6M9tkH/Umdk9mBT8vzmtsQggvVyJy1+sQyvZAtKuVA
SdqwgQUqqUTU1jQnL1BbaYu8jE8rROjVhRamaRModyrVGHCpr2m4rgPhrlvQbpiR
kp4sj4irm/0Dz94Zk3P+CbKY7KD1K8GQ9e4rDwVM3TGqMzdLnlSFtudm91vkg8Tb
Jhp7EGvwEj5JCzAfMbMM8LzRr3pXYAzeYv2/+j9d57SjhI8DZmO48Lz3KRfeoRjP
lzzalRsyR4+bRQxoGdUwY83I3LmZ5OcZXDoYjSdKZD45Dfr3B9IaA+mV+EWcqM/c
Osmg+tevlEjcRZNQg/O72Eb7oswbJyvqNfgt26mej/CP8S0pQj01wa4YTl+SMw2I
h3p7ixTtqn0OPBWhRYdVaNt0tAcIGipJD5KC2z1T7y6QmJRqNDVy3CAMBo/zzBdn
OglXhAeCcrKjIrvnqYFWwcfXQHZrB7Bab98kYAfN4Sb0SKX/H3KNbqPWiR3ozt+9
BMDFBnn7wPLqKk+QDwRm8ZWegkuL5bm15BQowMYSTBgE7XgQzMOYU31TnbgEe5R7
7/1V/9EyWhdhrjhXa2DXjXK6oVnS4jgJvSCczzC6i5UYmRjN7leMXlMqpp5CnDtE
nd+MTMSUsd3Y+NbzDFVGS9SaccBU4ZneM9Csr01ai8GEKa86rzghJgBArpmNk4+Y
gjCcoE0+YW4LNUi5k8qDwrpt3VltaFwixxIUvQ2TlZCot8490GSArkt71Q1w4Ka+
DnEmChGin0Yu1A/sytx+8TTl9lZMtMOBpmHE9+mvDMoo9gnwBX3cJWOMTE2+mkNd
4oFgg3zHflJGloaDFxAAdNhYmoXIIzlkp/9j5CiDawssnxIQPxfHMlXjZfsySULT
malj/MNccxiholQqOJT1WlewwHpwvluGFLLpr2Jn5B56NQasUAoGq9wptOvsMom0
l0ds50yra5djEKUaME5MkpIkGs6YMXiBARWRpWs3YJ2U6cGFyxMsgdNE2Wjsqqcm
ZMyHT69sxnMkZDim37CdZ9+1PnHxs2XZaerI+4S9MFLrSXjEdnhz96z5AQ4dxvbJ
71JbcGa2GUTTLVZ00wlP1cGLTbLXZ3b0Ou1iKWPkAQVcZuCPC8232hjSNZ/TaVky
obFGLlZ/LS7hSSdpLkMvupZOTqlXF1MbgQdtStHdApewqUZx4YnW3oK54JfxoVrW
MBqfrR5kg7GccPPr1+4W8I4m6v4A2sKExUsG0GV4vcOb4pSOmmQUA5JT9LbtHguL
PDPMvuPG50yO6fH0HQMOngjUFbh5qlvHHos8664GimfFlE34laiyknAsr6ovEsMM
Ca+5qZJd/Sa/eU2gXf5BCH5VDziVLW3t6zTEV9dGgVPc/mYNEBtcThdyNhi/SKW5
xtfPpBva0FNcwwvFZph+AKpGowNrbSvuh4xNHsMSXC3u+e7jwUtX9bWLtGE2VHcP
iAyFs9KSOwPsrtP09qVX5Xr9EmPkyUxIogDI3AAxAeYSuyXWco8YIHaQXeF1vG72
/ZKETmFJESMXMMR6sy/Sbqnwmlx7doYz7MPDuDhspyqTnOsjlF65hNjb3ApimQDD
VljH0TnkGsKeWWjdmYZZVv8dfB3xJhHK+C/z8LIPnewUQtS/PaNE3QnH4w5VeeCo
ycwTc32mC4W+hcA6egAxQii8cIz/CK9cjUTyAK7j2uTM7HajNCzpQVW3PDLp20HJ
TdSVMrqUml2dLAXh6qGLORtiDIl0FYgXV4JMYuFAwIDYbXcSvbHKwqe/f8VVaqGt
TIKS5fbzui7lkXlkRP/PejoCf/e68AOxMsjrt3DhlKYKtu9gVuO+2+/Gwq20Nfo3
tCk+rnX6jyQE+UNwAsOllshn+hqiyqWjOPxil5bV3l6K1v/ICMhw5++1mKGovGNB
XKaUVhIijP5kwPDCEgn3BFKwTn3FyMxUpvRXmTDBzG3JVV5CpKOHiZHVIFgnMLVZ
PqPEpi20XCFAEI0jSU5UhZGumdKKV/r/bE1N7SbBe2Ih/hT4tTFnzTVs2VB90fRk
O7GXErbenNJWm4M71CCGC2zZeIrlw1UP2sdAzte4rrCGkR/Vm7tk7fdNXQJAL0NZ
to7KfoQ253q9OQS6kdkk5j19jqBk8hOI2iQQwEMLR2yQGotMT0HxFgFVYHbofg06
3D+h1DCvPhzgCRp563FdyvXe30Jjq6Ht/w/vSmP5tdAdUXEuZ7HRU6MTqhp36HsH
Bq3fKJbho4n799fLNU3gURNHi1mC5oNyhss5+EKP91YR67IqwLTZ+4Zw/AQQUeY2
ry4+X7mYPtKn7GyD4oIRgk4ZOIE5HlgrlIsBPOGymVTtzjfyzyJwBKvDAfo2iS7J
YyMKvcF00qQj/vgCPDJmYUJziSf55o69yWQoM/bGiz8bGALQMxaVamGWRl7Ny1Lr
djxYv7WXd2e0qM+s6MIZuFMIJ6+WScePC5LuxNlngOOHe6sjizmBe7lSLea4Zgr8
NvV73SPoPxg9I/7X6SNm7465RBT+etCGdiBHp3QzErN+i9dI7Ex3v1g3GKT2VuFk
CVYaIufkhJgaehJet+WyYyrOe0L5RKU5e9zQbzOqbqVzqcFk+r9wvGiXyExafBFF
r0IAcdvPr9IexRMz/HCREDfNPMIzce9puz9bcCJpdCnI0m+h0m48Q8vTejn8RTZ1
SKes7vwqIEbacYX7dJ1eFLkTgPQP8md1E10H3xAWvEKIsK2Fh+B4kbmPNmN0DFBV
ploL+vfvJQ1BiQQEGKQ5A05S/MnD/oRIFowkqPcCxMXj8RTJjT4xV6vOs/SOpcUF
G4nSOuqQooZDUU+iy7dYTIbJUJaTOBy72q25AhIuC6qmCgGVGAglWZB3yXZ8CGJt
a42S7NdMiZlulEQvjXM3kwulDxxwIwJaFxNbzuhn+wsI5GpnOHuuOZo8oQ8XKDCv
WdWVrqgFFRuDNCm3FyHvsj+jpULqtxMY8b7fK4ChmzYIBWfMfLFUuA+uZ4i1+JpZ
3K2w7D/GXV4T60mu9NsPyVNfhuWh9Z6VbyvL0stzSm2TozuKEQtNStIiLorssNJh
tGjozR5RkQqHOkHHFmW5LUyO0KNzSPZmJXlravMXtnEWfRaP04EmA9BOcJIbcQap
IePD2rQh0mmL2uC2mCd/L9RsQAUpyYmltr4x/JNpl16KmZdaO65XUiwpPH34JmJ4
CYQf5MiRR86cvqLGv0flFzP4P8gs9HqqTrXlwVdaV1Sij87wKCHHF7ZIajiGOtNE
sDIEaH2bKD+GuKyCad3wfqYgM9Lxo8uevENuh4IAHOiDZ+lAnfYH3bofaQLz1LUa
OVg8g4bxsnG7v+x22h2XKeiv8/GGWrgPLJ2xA2y8wek2zXN6Z9sWZcDKlmCusPrR
M8ieNeFdl5EaaHmNRjlYpjsZUzzCF7IigxmiandsJ9ewtgHSUhtvq7V/zUc8WHUz
vSfjv8YVRiVaCYLATnWX8PBGw+EafdOs4XPVmxuIeeJqTQZzWXHfo6p0OKi94oQ7
uanzaciVjNxvQorS7qLA3KDmlg0wPyqehbGGjBCBVVII1DHi+a80yEFizenWWPzm
F0PLftfnBmtKkv794dstj9yx8Ov9tp3vJgd3LRx5mQegQ1Bx0g2u4xzBjtKLg1ff
AydiCCj2YZlRzmEZqFOwqLQxvsVA5nbH039ErYb/yYr7+ZV5EziS674ViehYgbXE
Io2SIx86YIZuOKGaH5G6f1+XHjrb2N+TGTEaft+X3eSABr6H0y4Vz5PNURM5RTq/
w3iUIubeHQAsepiFjSpmbgAu3w3S11XPHjde39H19sYDyhVK83l9jZG7LYkibxMg
HwWPtBkpfB6FpkX7BpwajGG82ayGZRalUO4C1m3OVsejDBCqzhjkDPWAa/s+cpAX
9W8/PbojD0Kad4keOOpPBeAIpig29Saq4veeKaTGDs1kVCUUVRL6xQwyN7yj6O8S
tX2JoHcFBZkKlU594AcTtIFFV5ukvKtOlTYY7r0+iYzRmdtES75OIjmzwxqT4yTz
yworjGu+N3leoBqR5kOWnRNPcWniWjFatok/akwB5qXgznrTeyFRha2B4nqkhaEA
cONrkpkcxEbxuN5L++4ZR2+72imbvc37hZKtpLjqLT8nkPvC8mlDACAUrnhpHSvG
VfBvdcI/OK8KMvW+Kv9e3zXUdH4d77USUO2wpoiKt9bcDdtIDXqNqg90XV0KvHmn
1pLLBRj4FsBddU9RDSvZhgsQ1r50MwoQg04S3f01NwRCmyJhKAN3z8wQyUz0qlv+
NKUutWjdqw05hRNxbmI71oWL4X2veCNxuJGM4Rnx54037c/GJJst/QhXuY+dZvF/
cE95P1WLwPC4nte8+OxgzxMuwf/dPee+tzT/PHNvvCTrBw+BiRTEUt6SBsedU2lF
kdsXX/KNgSR60DIx5rVIHwSquWcVI9892Gav7a5RpbbrGxYaThtSSsMC2Q3HZgDo
BqWJgT9W5ILZ+H7wJwXfppQwoJ+4CxW31vY7MdepnapceasysV/xNPikAycZv6GA
UB6xcywMwCVxxBO+aa5U8gKa3WKxMSjcP6LeacgAD0d1bz2+1fsI4pjyT4f91G/f
IOdhR+FmC/1LFXs+4paEbZBDxXuiqX9Dan242IkOCxBAKnO6BUnAG7GD77WrJg6u
mlaAYFO5eRSs1MuDs65tIIzcxJWCxCd6lbzzGNXMFnp40xibPdBiInMVwNmrnAxo
Ol6y4klDVk1nOz4zbnKNwj9E6qw5Mt9IWY/U6/1rCqrR3aAkU+nf9Nlelzh/wOMP
BC/xyyfZo/TdrNmP6ENgimTG1BH10CElbBTl5Bv09yZIajc6LkahHJarVYu7QHu1
DDHBot9pgYbpAmoYmO3AQ8Qxegxq0tcooeAyFVe0DNgq8TKfnz7LGPniV2yVAJTr
16x9fPwH1qzEE1nbuA40pHkc1mo5B8A4EnqVRPOtptD0Xv1yoKmx/6qz75AoOh1s
ddaYzcUCwB4A/GtMqj5OXkptb/wXjlyjDqxh98AIn5g/Jfaup0MvR5yTvy40a4tn
8+ovwfi89+CY+zNcZC3oJF8vb72Gsg2M+jNYmzU7SXm1xes7XQB+01gzvL6vYK1F
9dQd5gZD0dEFJiZf7uwjLn4dek1O9YVn05QHkvA8KolW61qcSmTIDS+W6/ckg+8r
QQU03h4a/639xjP2gkTEKnd8o7+OWhCLGpvcjdfRpKJ/d6UewTlNfQ229QIHhJ8J
E7Np4cxpKHzBwXKCgLt/TKGTbNqg8jYW2fib/j7d5sgRxm/iwev9GHqC70rz7BQP
AvmSC/OoTgY96qanKfU1t0+H08yz/WS6bXhT35V9KpV9XlUCy2Wt0XgqWT3bo3CB
nqG1spw8Nju5+6W3g/hM2kqLQkNj+USkhiDtsaBue+7TCz5fSDCKai48WwzV3Cw0
LT+TlXi9AsqFuAkeKcpvi4iz8TKbN8NR07vn+qhVtYfnXqHJtGF/OKOuALT2UJkn
vhnvNr45tlwWrgZq4TdckdAiOxGFv7+Q5XDhjGtBioawvbGuttluk5OvWv8Fjitk
S/Jk3tXHdA6FxA/W41Ixi5TO4vCU2Rasqbvwy5thRz+69pj7Oh1+i3XK3XwAfUxD
W2eiM4fy139YsZLFW1/U1hz/izcPSwpxnWuyXvkYMDR8O9i7qZDQnQUU+vB0OjnN
vYzhRPsJwHqWUHZ18eVh4V8ptG3rfpeDb5U46jaC2p3nkSKf5+AK5I37b6Jygv7t
YjAvbvUMiz6n4EbsjnpmAnpBGpti9gNPm8nytvbwL8FcRdvXU1Mk/WYeQaD3xUi2
S0FgJVTvT/S52BcN70rjD20mYjlwiGHBaThZj8ET/ZY2hxzq7rkbXzlDqi6YWpmn
rWk6KSr0NstOSaiPG7Yqie9FW2wWMQdcEfoogG97Aa3oczWQRpPtgsr+zGAN0E4f
ZWmvCMh/0+B1+r0uwlafjIe8ZEgFT4PboDTR4OT9rKBFEZMj/X3DljdgBbUB+iFg
8YEMEhbTnjbmbtlVwJzLmw0NCqWW92rEiDCtWpulwxWwcJdCrnyR9V304gZorqo+
SecDRPyth7kARRfagQGrLqMlO1qgZ1aB2dDfr347fIyz0uAzJpipCPd7mmJWJp+N
CmKQ1UXYgdPYTajbaJWNADeMPRKON+UiZOeuKsXI6i3zmqb3S2vdu59X5JhEbrzV
2N1VHI7F/0qubxgVfnbMFkWs9/Uv3wxln4VVVKUpNAjmVQRrVfecNaNInMRbqJJp
sZrWufeCDB3/quzaH/x8qOKIeaODgfnGzli5PMkwKxpHRAExk7K7ru7Vj0jEDawe
O3ZrQXHJbqeIGWx/LUFFfzrEy/7PoRgpmsNDy3GNAk7gIbe5GQFoKRelWCFome7e
hWH28749mEJ/kIwHzrcbwmIKuMIsQGsdLe2jZzCNWctiSMmlxYz1FJ6E/uwEk2jQ
zYz+zmArwqXLcmPKarec9O2ZuNqyFJ2ifWhKOX5fG767LELtDDYlHrTT3zeO4ou6
kvuv7xEGQrskJr8Y53y+vR0L4dk2VISF1rhDxr1w0LF6T1nmrwT64ZsRQxrw0Ldv
9X58M+zwVSDuvb6d8SpYSGUDR4R60S/zfj8tOjF/dHA0+kpFJBnO+PA7cPzZdrFj
omcCrxP6psTcOD9i+mSB9ihjdneFYxrWZrTkkjK1i9QiIIzP26PPj9JypygaVz4j
YyDtD8TkU5zfR/nVmYmTd6P/MMtyuurPT+rXGy/QKpgIr/Y0pD+X8YMA5deUthwn
CwE6Ze9lbI4AqYLisC7c8sphykfqjcbR6VBraUNGBc5L43DY1tzed5z30cXIiwyv
z6DkxqMDos/NunoRuejll5GmW7pFPRIz8f8z5BTunyi45/4/dRzyo/fGI36d6TJx
CnS9FPjGGMVtc/XGlH+BLNUs9JmDT27xcF4VapWdMo/jlG6NoDDEvV78xwpsOUXd
A+6HRQ0F+MDUl2Dc7NWmaZryiDWN6cwwJXhJK2CA21eJjw9CIeXuyXdewXIwWbmG
Gz+pyoNoI0gQ2q3oLppEOg+AkkQlbd6gBlipy5VgMhCN/Cvs+LeNHgCBOIey7D2S
/cOA4fRKEhs1SW3igQBO5sIoyy6nbaotDvZj+3jAXcIBXu4E69nyFA7BVAVZ6SRc
gWPyZcdh88x6iwHnLqxnULx6AZMty0KIjkhtrBMWFcSEbSWrxzkei0dXsbgV6N0R
zyl2yLIsT29xwlnicgCEk+7W8dVKVnIvus+Y+Sw1I7o5RmH/UP6JeQZKcQ4BB/iJ
ZSeVnct6qX9Ji0QXSOlorG4W1JqoM3FaCXNnasYTkyjEdPtwwBrIWV/zjvZUr6Ou
TjwIPexh7jJp5Ynt2sjnhAQASeF+eGj0TGhxX8+ShQAOs2U+KvWz8LeQ69x2jU05
gZVQ3+Jr9dx7/ViDAPNHiBki20Fat7wbfm+sJPAXciT4F3EfM1eralRCmyFdGl+g
BO5l2/fSEgXv9qVxe/P82RWkQchyHe/xmZaTIHAXb26bKIFJgEuE2SPaEvf4EgO8
pb5V79WY26MX1uPbX5xyCRaKWBTmGGAWoc6BiY/ReLDjwweN8RSSwqpyZnjh0QGx
HaNtpVf3cOEWtOY3J/t0uORShyRPxoyGD5fVSDDeo28WQuaCLDe4ny80XWcB1umQ
hLn6g8p0Xvqqr/170a1sdWkKozcRhdK0L44+bSlSte/cUSfPhCRfp90TmIcqFl7n
UzW68M1DSPb+qGz+jM2VCR7zELuP6BNs5CbIToKOvAx3XbebqUks0BJ6mfk1HAnL
4kGYwuPRIZuZLAJ51zT/DEualsEn6PiyoJAONH5FvyzdpuKUS521CaPwjKRK7M/y
CUl3X5mwH72ia5QF7gbrg6e6Mkb9yTW6zj8UnY+QgKK1qJ8blYkxkeSU1UqcN3QD
7bOAJ3+7xfnVz59X4Q2q54ZgSQhIzq+sOq4Y5lEEYYMjr0k9dURv60NNXwjT3DZ1
Sjy23pshKFmlmhG39Cbuw4LqiEyL0C8/nLjhNZHL7EGF2jrqmYVavsfrxfERSSc2
tjUlluLcDayGOsQvGv/UEKWBSNtkfZ4Fh58bKois/auhFojLTP//g6ohEjT3lfl/
mU0ZMU5oWGtls3EGAGVUqspNVmp43Qv6Gpo6h3EA606ygzjZtXclE0z6Pv58mjS6
pqqTRSoiEJbCqdWPRoAi/0VfM6rQ1E7izXnnTb5ohgV2KVlCLpFnKJMveWrOiOAF
Sy6mYz/Qi+U16hnneZP9uFS64LbFwMmzTr1NhTMhPlSG3Eyuz7RkY0/+tgcTh+N0
kHfFD1Z+pi8MYAkxpztsAEfl262wSIp4w5oem7DhyBTJqwRAjzi7+1h/KSP7cJYZ
EMlcHbdxDyMqsG//o9iZ9+4UuQUOuJbDzpp7ZMfUcpNVpqakbAa8TSkEzD2st6Oc
ROXUTDyLOLvg0YtWzBBynT+LDWTDL2jSRsaB0Mm0qC/KoCsuY0d6jf3HaFMmvNWm
xyoRMCdrEnKBvR4bArgj/NtLlq44EK1E615L5XrVc+uzDq1ReNFb5vLVLjasMqCf
cnh6oj6Kp4MxlJM/F+OyqAbcK0Jd5HZLUMtvZNRIaheEC3WDpneKqsRrldCs3cMS
VBbe0ruku7LpTgrHksuCoesm0CjETkqwEyx22KzDo6X0wkPgL6unXh4fcYt35kqE
8WMy8hXBPIB5CjpgBMkqUs42PrY4/QsucPFCTRJMCrWpuBRACunULCmJ5/uQ7kC4
AZV8Jc2XBfSkrCZlYS06PCVthv8UjC7tasaogVfRU3m8ipYVGId+wM/wQbxwTD2g
llbYElMZklpeNmGXw8ywiZU9RobV0Hv4Js5XR9qm5Mtmu4upq9bqlsEfY6EWmaNZ
6aYMTQr9BCpS4uMj5UYR1BL56cgAciepxpDkKBQHApvWshIuqR/2+ZsGubyuxf9w
tVFp7bAq86FNYbrkTepSsCsyLVoUey2m7JyFp+L0sQ99juaKZ+41+pvtf7RdmBw8
RV07d4gBSZylqKZgpRqTd9itBU3TZ1uaIueRyLq9pG7QYdTC0BhUBOM2J79igvCY
2VSAPxFsB5JMnaJ296nvI0H0yX5gxhFFDsFYIbX2Rj0TS6tsRNTuLt4AXVuU0V9S
IJJnLj654EowoIUhYmtGfh5M+0lKCX+EfCQpjxhx2SSy3JPH/OBkKLojLdnC7XRE
JhEuCwEonzxeZ3fYd76r/7J/dpCA/vyiN0MUFcvEPkPBVKN9Pv6ve9mFmJNl8CFQ
WYq4gh+qiZPsEfAyrxHW50SqMWTq4pazSrnu2jy/SAJcqqB4PcOyB6aD90f4IIkS
xgrCxWOIE+Tjr3PpZ2axOmREeG5+3i2WyYYHy61BOxaDUPha2p/MB8K9QUXVsX1M
sDiJE+LI6lz7ce+KMfcZ6LLcPk1xNIPbwdkOKgebDpUf12DkwTNpWakk+HJsVaJ6
1PHDmAhAW6Kw825AYoFUvV2OTaUX65qPO69S+/TGPMT/YcWqsw/0KVyEbbAhwXi3
KWRhLFDPtvR2pZa3cLhD2zjHMFJTc4XF5cPety2QLKEvf3fZqgRd8nsj7q32erzs
818opnE4xFFXhM6VgX/E+WZlO0NSV/JYbNalIfe84+DXznR7bpInLKB/TG35f/ci
Oyl9GfVSzaOhJZxyXqJTgOxmgmcGR5/R33us6137D3Mi0jVc8yO1R+S00HSNQGgi
MjSOq6uWD0/C12v5Ikz2iIMnI2uUJzzTvBHbLN1dvVhLSwT5i5y77bOztFNko0w8
7TRdnNBWXPGrs07tx+jRxFCR3Vd174U+adg2N3eD5b3kPcVTVZeHWtK+obPSAF2i
LPyRPoS0jnNS8jQz6GAzSYxK12img4dEGPV5j46G8bIoN/GKc7H88qS7R792RBCB
tb/6lktQTIB0oeViVmGbRgKCwgt7NMrsMw6qQq8om9XAEuYOVzmp7DDEb/s94WwW
Pw0NMV+3oUI7Rv5AzXshO1BjDUdxkMQ1vqHDeLAyxKcZsV9tAVoFp1Bvx+Ut5lEt
nUAPUXE+uWUmVIUf1sL/GXLqBoMEPyElQL+lfTjMB4D3GEDoaXirKvTop5q1z/Se
03PEbpeU9xiGfK1/+5gUOBDlWvUe0cPTy2xrqjQrMSKZMO5XtC49bEWlbR/rm2RL
uHwbarvUP6KD+UkYdZ989bbHT1F85t/9o8YK/g9JAgQ+YCNmc9k++VJOvBccM22f
MKEiMj2UPZzp4Q2TY7o808roTu7C362PrQzOHRkL5xqFo9rmN9OirV0HGV8yz7cu
1iUBT2SEMXREAAX84WPRJ+SX1a8FUFUlqe2HBEEvfz/btCNdfCMtQpfCS6tRx1FZ
GWEpgmh+XuzGmxbnXz7VIpCHITxtGDudDrZNFRQjNnTwYxsFY4I7lm3HUE6aM1IU
F85ukMH2m7VPb76hnHSuOVaOiJg183iJmhuHk5n4zr2xWEnl6SQTe5WuEirEx9Yj
8mw3ilvVujg1uD3dnHKiw24jSIfXHm/dDe4yaV20lkYhJUgsL1nSUGIsrDvVNO7p
xsuAmEeUWvkmB8jHIwHanp/Vqk66bderxJPevGOLS6O0XFZdLu2r76rZG7XdV1eL
pbHtBXyu/ile3Qo61k4Z7YVHZvdEamU3Hh5Pk9WPxwSs+fom7HTvbPsOvIhJAKoY
BbDadHU1OO+D89k3VmyTSSTag1XgyC4bGn4EzwbhVyqCEOMsnts6npLySfJqhdH5
KgAnaVmYIAMtGHathl1ixPcUB6A7BpejPMZIxKYKEg1jNm56BCD/2gxWbqPpC+N8
d/5Lqu30bfR87eYKBsIX3gQ10+MgpX9foM2rrTKFyxI8Rhjwc2CXpqLS4C/o8RE3
g94kmFUZlhqZJUlsAMMi6PcAjcf/xjPn5ZI2ENrLKj87XSl3a4XNu3KpoOuiXsmT
c+/dP6sTjdXJfylimIx96C42sarz6GSalpGACiSUS9K4tdFiTIdJktujSVEI5a4e
1gmhht6FnE3xFfK/65J6DmEVXnBCidbZT2G1cXmu9ZG0vrx+SFJcek9+6+4kNESP
iBi0RQ4eU4pXfqCYt24fXHeBXSrAmZBuPYooUe+DRZFVxn5dv61fvF39FmvXdcnr
VlzGKEXUF0HkzH0C711CYCOOzhsoXadAyG70GYGsk+mPS3A//xPbeO0bW9o/zUn+
KyIBQq/XHebtcmq2G7KL8ZWgSjFGblcCuLk19zSud+k1W1KDM1TkMOXbqGIVGaCJ
0Oog8HdLTTkLm4dPEqurbgaQD+BEzjbvC5ye6DnTJ5qh93042o5yYyeKpamxvsPH
dVqCl/bLFg8iVv6TNAU4EV+lMWw6+U0YX6B3FdVOGByduMgmHdP5RCpCY4c9a4Ld
dAjMvU9rir6kC/Ggw6H9WPn/ncDUjbI7UP7wAv9kVDslBMM1QVkYaWBhBIOMjfzX
TVY1leIZkIKKN9PePi4R5p8HjQ29SmmcV2W5U9mzYkhssdSPA9eI4+7zK8BAwN47
OLF7znTwKk/0PvmR2E1Hauy7eq7RqEA8dmbZe9kMvROYsrrUrMLbdAp7PT9uQuWu
Acp25idj9D7iiXjAWuVgtohSAoI5CKbBBUN/ww+I7W/hucv+73gOzbjEoRY+Mepl
rFnmtMbfP6hEfcu216oSiXwEyTTezu+NuTPepZBXavZtb6WKTFijCHQXt0/cbuNt
RRi/IvZlKv1fmWcS61La4P1k08X6bSRHLSHdmf+uJTSfjRAqDLumaS93Tn5r8DZg
q5ztBOCxHF4s6x69+ZVhLykcwMEfZWzWm05eUQSlDMU1dVXOxaSTeYT9PCUL0Z2z
3ZI+othOVvbf00hxD9h+ip+/LmyRuMhwNN9XHe9mjI8c7/e+mo9O+Sq6nLR4c14E
YKt/T0bxPrjZIn1KF0DRGoNQ5TbE7AUGk6CNFVb+7I9a+MFMVnheIeOvL21TYgct
cg4cYQhkw58VjZifAZ4DhZfvYypFaFDjoB4Q06HuECXT7tnqRGzCAvzn1KV5Z0aU
1wyxclwddFBTrVwX9dcb+Nz1stDG2wW8rK5TLLoC+BLRkagw/dtmApaXTwK4QrUx
HOBsu8ZbLoFWhs5yxBfEfetQRwAIlpFsQdscyMPb7RXz3FWHZDj1/TTjJqCZTx59
aKrrbIoDtrGX0zil5rJ580lmrX/YYlfVGUUEPFXXhrSJxrtSbADQvcQVSt7JoUk1
wexV6Hm3cKW8CqesaqEIpcgHvGMMbEiCyHbq4nQdib5Bu2JFLhSvg/7MvgqyA4oX
p0jcNtcTjzxpm68Ofbon5MRY3CSD3uIgSA1Iu6A/jjmDlLvizP50rDBG3u4M2BBt
G1Y2kdI71Hn27S+ch/YAD9FlmoKJNlfyQxwPOeicBeAHqrrjr2gzY7SWXFJg/00a
HyujkNLB9nqXTDf62dCvgzObZQkBf+I5BDPazuiepDkKMsuJRs4y+dW32p6eEqfb
WYoX6fZtnV+rJaRSTn1ow0OwRp5kl0KJSDtrsWjMjvnWoBXvqc5qs4nlNDoicIoo
856NCDjgu1LTa0d7T37strAmJm22QQab7WNIRVtDUkZ90VM2IuK0xvbXLkWHvdWQ
oISiIMhKu/Lqlvf7wgwSrjtQ0YOajaVUpIcZ/dcgVU2tu7cuZXhq/PUvdXjtX6t1
Rvb3K5DNw7fw54SXEWcIc20IyZ3AhKHKTrcnMAJ3SZjeFDhyPsJ6rzOTEH373Qjp
jK7laW/hoA9Kai8b5XqZ0YHzg4ZXdceob0mIsNHtQdkwu5C+2qhsL76WlwacOzr5
GIL54QWq9KS94kmuDunVMcw9CIS6oDhBo93hwmWvfbi/fB3THTNI+SUVCMVJyk4n
rqZuZQjsk/PEjofZyNRP5Q4ZcXNBkTvYCqla9hwPho/tArg8x3A9DV90Qw0LZRpS
1ONerpp2JTvVqpShtRA6b21ZYb+jgIBhkq4MZvjRKRJxwMZw2BfP+xgWmWaQbqv/
67ao/aQjsUPFpT3YTRAz0XkLa6PAUdtbSAD6SNsgLRGeVfiglTEUO1BVwgE0MaU7
mLD34qAksSqvObGZDBdxARErc95a/mcYtM5TVyMIzMdZpPYxYWbrg9lr1S69oJNG
aL2Uonp6CvqH2xxYIWEPL8Lxvg220RIwvAG00RkZ626yo8v6M9k82X9EjnFoAPwN
GbAt4lPWfPSWKhB2nQkc8a0sNht2p6++QbPAyynRf8+VTFlY0A1LGG5OvS9tbaJA
hDK2ol/UiTwKHVmqbiQ2S8XmrItRgREDJVOEVdDXssxmghcPeYEMYmGiEPnYgpGk
A91k2f5ggjdtJvAIGGV8h09HYCjC6u9f6QNZmiAE5AK5jZudoHr/7wC4kuKzFaAz
WZqRWoWzr20UXtcv7PG6IvLjWlbs+uQ5yi2gQWq+mwIobCwyxOUVVuQcN6vDvmu4
wLFYfMMBKIcmfDa8sa2HsvMSmJbMnlb7eCMvhHrcsix+SSKgW31hrIXj0XLYfxhK
2XjVI4RjPkhn/oqDKAOx9SKMRNVZeB7+vq549z64o3ZdCoHOEBN2hI27yAInF2Hr
pnGcDAevfm57MN8jT/W/QnkZCw0n5kibARp+f/v+X1Z3Rs4dsGhFQ80aN1uOcP9Q
+WBMjk/mqCF7EKY+cdWvIWppYmLL7ZPerl8mqyjfwEq154q1v+nJl95Q6fSfTmov
J1I6coB7FOt09sQn89ZKJnmPmUtekwDX94hBDoS8NFQPL3MBy8Snw4+22uzu50VN
Nzqr/I6NNQbolKZPP6Fz2YNkkafD/fMxqt7aPgGtsXo3MJfMg8qCcvCheCTUVW6t
oUgX2jo7shRZ4bNh80y04pfycUAVb8HDpZiu8SG4ipDwQ2SZ/XciSU2EPXEaJmpR
1DN358gmuykreqkuFIPq4qIs7O92ruwcH7V2A7NR7Nl0sOAqL+J2lnv4oh47YbL8
7pdRwrAn0at4QFKyM3khl8VgaID0XWjGaE5jc7doiRaT9zj1sF+tBbcx64BJGjAt
iZ21rsCaOk7LNIB+k+WMET6mYtO+cIOKsq3GVmJxcsIqgVSI2dpJ1u/T2ZbqsyP3
Qnw0le5jInnhModLthRg8eJk7wnh5chRaDyLP90MOm7bFNES2dim+lPaMVznLxOB
1Frz6TRJyIWhU3PLvaxVxH8ehE+16YO65iMpv3vLN2Viqt+9K7se2K2E7s7tarFZ
ZpagyH86NZ2NNvDtxnc1nzbpV+7/Crg1ttafvgFA0rE2FZUfPzOyENekau5g9I1L
KWn7AoQf1/tkiEwV7dBpIq/NJh9nN2GpBHtxAUPnh+XCUhcdx4+dyeeAcVSnUArX
6/5Fc9pdXVwJfGp2Zc93XrHa3kn+7Z1jTNnt8SSH80ZpnqqU60f/zpNlrCMoUPyQ
FHC0Yrl0s6KGfAPR+CofGVI74d2BeekOJRhCJKoZlyVfTG9QGMyA63QItU9Auk7p
OUdPhWNfl1JZQfIrK19nGf0ZW8tob/bvKWB//mJUPScDalZaSE0FJUYWPDW52ffc
GzBSH1VfEI8fcqWlvvV2EaXAFMxirCZJQY5lWbanplBBqsfYjLv4DRrMMIQCPU/k
AQON2oG9AthjeC0QwzBudZxOm9WUuA6pnQ/DQI/791XszfoP7N9xadvQKCsgFNfx
lLVegVrziyFD9eOjva+ynzERbQBVRtROq5axoOlGNvj1gY3ceDuVkwjH6KALxDD1
rz8PIPegtHZ3JEGoxj8N0z4DPEo1jGWY1hmYSMb8kioLlhEiklhOpdm1R+3GOVxj
1tpYh0oDSAFGWMppU/7Lim30ulLA9Pj64r+5bcDbDSJybFmOWt9MpxwWo99y+fmN
sXUcE1S9MJWqw4JKFHMGlQNlsWPOYnvI4czj7MriATx5dOH9phtGjxmV+56JgwZo
BXL93F8B06BdGMB9twSCsRvrAOCy96A4/hiCylcpZ8rV03w3RozzD+veo6c0O44I
uTG37vC+R9hPsLMsAV7+8IRo+V46OJ+SCViFkkdwC22b6fXe91a8R2kqdU6U6tt9
7VOJ6NmLEDEPM/PM6CoEFhiBLLI+8c5HuRr+M/DDQt94akScL90C8Fr+JmpPjpSR
odWniN/z8aB7m8c8Dy8EflhYlvPogAHRQuLcUtLDxD/i/TKIfe8ScBPwgRuxZ002
ujunkjoAViUk/U33MLN1m0rHrcWeK3aQ3jZzOl/SZV7HgzQybV072lMFXif6x7g9
QvvOwheviKXKHS89/lJhzuXH11PhhqHUm3sfpT0Pl47XNwLY1EL7HDD+KhEFmdlb
Z5XIsr48v9NybQmoHM2nW1gh8pXWapF1fmgvwM6KTPQgUVBJmmuxpvYO21WeIAT4
2EnYSH0poSKDI/6gUSqxoBfKTzM2JnxXaJfWzwHw4BFkLMYV5pI1zkQwyJHIHsIK
F4WdxZvK2ExpEMkiCbfQzV9EoHJQXf5fMzADxkXs7jyZed1UipNx9bw6jksIIhAj
EFX6XO3+D80il//3gQNZov3fcHNmnbnuN0KdmMb2rRC5o6IMHxA74mOQOf8eskFo
qWT6VepSyLLXKfF60t7apD8yBs55vXzSZFq+Wx9aFeNypPy+nGbSCOEf5P3QMkGW
R7mE0G7/b0C8W3cwfJaeZR7057L2V9hAuPsOJMFroUd8Osmj3/MCZuY/XYdexakI
v63XpS9+4u7tTW/fiN8iI42BRVn19Hvr0wWoZvhCRS735f9vzVNMnQf/ApBy7m2D
UGDzxtWPbPIQ5ZWBW0B93ELtpap2zF2UhsDE7hb9VC9kwIO6Tkx1RwAi5MoL7WKg
dbh4oDi1HD0LxybBRY0nXO8+aApToAlPrWD0RefZVqxfwLzPpYzYChSbTLSxqH51
lYhd9eq7SZmQ2EaMkorwPE97Htaw+Uhvi54qlzPS8jD0hdhTmaCsbqBa345NnIQ6
Zod19xeUKrtgtPChpjAbqUq3qrbIoljs6L1r6WuDYBEGvGixS5lwKsiZlL0lX2Kn
hap1BT2pb+KNTnFEbVvXe4axNQoeRUSJL6jlSsWISbAkiDv/xRMfyCGTgAupFsbU
D/T3oFee5Zl7lc+qx9zIQdAOi/QisF+vWxquEptCVxWHw8aGiWaefoKseF+VWXNC
Hd3rJNldTKGSj7fuBUy6XM/jVG+sMaVBJbU/Svpf6PksIqXlauJDYaruT3Dg0U/H
8Zc6L5ejhVi1jKpDx0AN0OXBUu4ivxSN2pLG3sDPLs8Po5iOCfVQN0FgONQwu9UK
ZOEd0DF7LjrjNz/23VWul3t+DttlKl7/FzoUoEf9wpmdsDMaO88I7GJ+ojzFycFg
HM5nI5lXOzUWf9Vn8Bx1TENUw7TUjq9F8FNCRewhCy8xjWRj0PKFYRGN4aUqQNxV
HCAtx2p5B70+Q6qeitMKMfhMs8d6k1wcdY5zAL9btOmC4HKj2jhAsEXsKwH9sW/N
rPj9h/xgRaUWPdEACmtCDFv7QYPHsVXacNJPzQq8s/4dL4qHzQkzgiSV4xJ46lCZ
yqQY0la+l0hFOm3cJjZ7+J5dAea2EABI6ajmL/guYnUeSOYFIXqL0qxlLlMnEnNq
1lKv0P0cJdXRTAsFx5Uv+wEDToIwyKuS4xDfOKVW9O+gnOYpTue87+Y2R8NzaHk1
bRCj/L4Yk63DFK3fKL2QYaVv00nC7E0y6QYnl6tOzmEUfYye/Nbcyxxsv17s797K
Jlw+n3xRtQcCBJSR2Onu15WEnw5OWk40pK9XDOtIy29oqt10aCOF7dDD/BwqVDXE
2x+dl5XMCIuLCAlHHEE8owjJfYjYPJL8oeE+GE9g3qveqb+fw0UF8LwGmwo11JQU
ftGb+iv+MQNJqDPgvcHExRS1xDKxKHy22VCMlGmKsgMKydW/G3zBVnw/0OotTwhn
RdpAjRlnMVNSFOQlqYR/Nh6mo/aI0Tmx0zc23AJFb/VKZK9w/JG3LPZZyzTUqTaK
ZjyjFkSbLuOqJWnMpPiuIGHyu9ZEvzVSDgWuiWQYp43v3SWVOw9pLoON2m6jZTwJ
TAxplqHHzoVAcl/20s2fjzy6RHunocQxF8MoIU9UnmNm0cIo0yASluBALhSobfuM
UwKRc3VGnBbLd6Drq2L/luON1lOKRvaJ8xLE00NvhkPULzgWxGnRS4jkBbiXaAqj
NKS1ykcMDwqgOMmxa92vCUeZ45SFgoDlGVZDqkUhGZOnZiYpTPJaGXi+sM+nGqPW
FluIQycaIWYtN9nd6w6/4NgxYbEtzdNZOKJ1tniJwQPh7FhB2VJU4LLMYSDliY2R
R0Wc1oo0oUEW9S/2qQ3Jo8F7E0IYDg4dxPEPgxN1F679hwhJOPFz0Dr/T3NR2Pna
NmUjealQJDl3IE/zSnrqd6AjvWr473SEZS4DNZmYr59MLXlm44L0Nk0/wOKTLov1
GsHd65JNR79riLzcKaJSGzYvJCJWNucC5XbH29+hr/UgyQcuJi62GwK5zxBBbCWq
/Zhqhbo4az3Lb+3Ij0GcxHb3R4JKPTdjVYSyGEMw5ErzRNOqh2FcZzeBpFv3I9Ha
DfvHAgnizeg9H1BHSeDnA7ZNRv+O/g6hPQu5+SFjR/MixcmgcM+78O8MAk46okcd
Vvg1Ol7dQWe5ARtBXnFFxn+GfUKkpO6Gt3fJ0bBZdCHZb6KGsCp1zFw/3bavoy8g
vlng2g/6BCHKeIhdKU8LiY7wq8T4X6K9oQVX7OhYRe/RAx1SWFsWqKRlyZhmJ+7t
lTkxQO/2kPSsjI8DLtKdreCY8FdEgXT5Tj0n1Ph+jkrDfLSZbUnkBPrSw80RYpV0
9ffEISnNuIj3v9yaQOWy8OSCs9FdlTSMTdF3jOOme17WifHcEoC+vl7ZOEeZ0bas
q2qWTgdrj4xlD7r9eTt1lXt0Du7wZH6QAWngKHkJC+HFOXNDTLo/XIChwqNMhbCs
vDzHEfXwOa7Tjht0tgRArU+FJ17Ma+jIfG7k//ci6EsDSju9elXY/8jSJsZ3kBNj
Wpi+GuBN0h2vJaZ+1a0UrTzzjQPH84eATvAKTHoE0woO1vWeL0SIIkil4rrYUJ23
VteUXPFV0/rRsyCrmZcO3e7R6O4mmgjI1yPk9hzUdsIgMZ+0wwrQFCn/VoMyGOWQ
DjdqgkExsxYBB77Nvrp3FFuIuziZuvF/a6qJ8Xga/ncwC8Y1upKQ5Yl3fzRjM7fg
a6nBd962nB9qdKSiiLc8SaSCiM7zglJB1zhv0ld6P7mzH6XEbCxNcR6UXqQR3CDG
ANBJAdvVFmlkxi8E085rNBwE0CH7qsB0/XC4ZxaXM5J9hD/cxHWU3TTjjtJxFFXg
EQG7XKAAYNimkrh2+bgz0+oFpMt73S7EBbn9F9dI48KIl0mzvES+9XsVagwjv78Y
vCSWDQ9BxU+W+r/V4qYcPs4W1JFLmbdVun7yq2MquiWn4BhSJKUKbviKjabuG7wb
2ozFCVgaOa8aej0wuS8SSHfNw8rvIvUxsRxvfetObcWa1t2f2Nxz33sVsrjzOfVO
mwHr5/Ob3vR5f5bd20vNv8Lgigoi7QU070vfVirMCg43ek6SAY9faUuzyYNh2dKS
3ZMaV998UhgDZDw8eSYE9IUa7nIEqeQvsYtNtjan/aHelMUWhLoGbHH0DeU6rBdC
JB5RaX8gAejkJtZOlcqAYTazLsn2RApvMOCs/6gwDzJ+uYb/RE0XKT2oz448WtbW
fVjbq5eMzPR4stcWBjwsoRWVHCrvxeT3E/pEGjc5q09L37vSxucU3p46feeA2Zgu
rnjnthlQh/2TZLB3FyWpA32+YAf1LZvEl9WeM7UJ4M0rn+TebzcClfbVATAoBq4J
1eP1+KzhO2RjkbnFvgwYXQlnGVdJef63S5vI19N759naJreI9iAOloboe3rtT09y
PEGnf58eRuCWmcwNtJ18KiQZhGi8fjHgFKq4iya6EqBGnXe85a6h0WS2Q7VFuFqn
Istdj5i0sB5Nf1oAOkD4DAzbxT3dKg2Moj1i8ck009sOxxxsMwkzk3PVvoN989+k
MD8pZkWIUeWIhX8d00/gAFMMEV0nsvRm1s11FlBl9WDo/zboqtZJjpBZbXULRHQ6
RcbyfO1EmkfbeCsldrPCw1waEtl2UTMxnhd6a3ns+NKqRhbh8gTnVp1ArmN4b/fe
WI0uFvzE/YRE6yAhBdqxQQsu5jWM7OQAon4UWC9B360LC8mRU7GI0Bgzs+NUoYFM
0tWjCqeUOddTKVBKVc9IlGRtNQKnYRQtGi7zdoSeNnFWOxLPOSkkCHZVID4/0iH4
6RZlTzN9KX/N6SMeVHNp/0JqhIg/CItXrdvXsVA7KXbu0n1W1VWayNygQlmRU+2L
PPlY100ojoYXDsDuhnOryAYgd6FzkuoRbmocs7U9nkagusKT3pEwEg/M7MDsW5Z2
sjEzcCzy+VvZ/DaasHybpKMaBFlHr49x1VvD84bMKmiTZW91O4tA856VWTTwV5DA
2qBeaw0zvmRCMFblVp1KdWLN0k2lvVYqFviORhh20GVTSsFsf9BWIyPE37Ydg+Yn
7Dv1N9DQJfhir7iR49wExc1d9X6F1xhn96VNPiQ4wGwh4BeS/qEnAV/mlo4x7gA1
Em+FsUlebiE+B9Ew33UMF84BgqPwFzS5ml+ZBoGNh65ojoyyc99m2PVZfuzrH+co
hGDaJCvvxqn8598+vYsEnirVH2LFLNQEQykrQ4MDgOBD+BYNg8cM1r1vYd4efgzz
IDhq8R6pry5x8pZwygGLaG98SI9tJAYL2p98DZ+8eYJhldN0dPg4ocGgc/kczF0F
+IuBWnXTmatEH1wzSXKvJOTKlNgRuVDixzPinSyAuO7Yr/cYwmbkJrSBUeCaW2i+
exQWNhpDPFydmyImOXvFP2Ie61PD5oRMnLgJ5LPD5hCfyTGbmuXfbkaQ2bdrkfiL
xyZld/3RHLxIL35z43ZT2GINy4NaiSb2zOp9Dtt5bVttm2UmFCZ2GPkDfM6K1Jjg
1GZGJ9BxW92KixN7gSSoJ+dAOvKBuovDItXV1vhZRNA3g3reaFFEzcYrLouQLHf4
41bhD5knYrI9zQW0jU22f0erHcZg8HOnAxJ3tjiQwoZv0FIDqb4bfVdtrAwtOv5e
Q9L57ubbkwebLUIDOFuHPYD+KK/iQUZEss6DwYNlYWOFf8ISszANXyJQtUDsoiI0
TZYUXhM9xzmgdceYQHR+dqRhSCyIWqb/vBHfqQ2dKTKIa/PIObiGt5JbX2ke2yCS
tKZ6k42xnM5Otxx8/B/ykG6pMs87xEl5mUHh4FWpaqYGluB5MzykLRgbr8U2U8fA
Sv/liLxl+5SnNsIC+RQXPvISCZt33H7uBoNhdmmL5KAmX+q1l58vY9wSj0sQDjlM
fBmuZLX55DQMdixidOoN0Y5kHamOQMCEvN8o76+JGv26FTIkFH+Cd0hTenpD9trK
DBLBf2DOQo95W1Jfa5u/SWdAYhT5zfWF76dAkAWgyWr7Jo6A8j0Vp/Fr+wvEuq9W
ste6FU286upUVF7/JpoB5wCxskNeJAg2whycEWGia7IiwGSe1Lu629R2VejMRdHi
8whCEda7SDdmigLFeTqrsd9fo0AO1TBW7SgvCrsrP6HaZaKA4j7i408C43KsZyZY
lh6Tvuo4osRn0n47R0Vv4fW4FeHyewAh5prYhqpoOpE4lA7jvltgfikFacYK0PyX
npT9+bWJkZ1fsIAHT/X02F718rGRxwdXkQ6vdxD9fyl+0zlLtTZmZPpwHFPsr8UM
IqFMYDTcGsTBeudg54dniRvJZG2CNA81ZfBqju7sZ9ZywbgMeXD5m4La+755h9OB
cuwyQnUDUHo0UIxEZPoUT37It/FM3+d2LK46Iwe9cUjXprrosyZZTCmogcVFgAoN
7O89zDrNEW/UEdm/Nacg3QTUEyskF9odCCMSWGNzMsB43rk4DivY5bAMjsXpsAk3
NvaZjSRirmcPdGYXjX0g9dcbB/MstAWn8RMZcvdRf0eFR7pP9e1aF3yCW0hsbJRF
0Cu8Ckf7hIoaJGslzaOjgDurZUs9fz2I/LomWtujsf3BI9HBe6iiJs3b8XDUwnf9
dHHaLhad7ypMUIcqmeLPuM91RnTp5BAQV26yAwCHeqqIFf29nz87qPvj7QGeMAwB
cIdzqHTC8y0nGVYBwwbn2rEWrGn4N8HOSt1sx/znjHUmNwHwyApcurQlaOLx8bK+
7+QmOJkMS7KauqdmbgP/sDj12dGs6kMJqAnVIBGvYQo3kZypUraBAGZRfv9b1QWz
/GwvEfU2mYRpR8nYWVLNmHOc/JF48dXrxb92zZhP7sMtK0eDKCyDy2gJtdnqTA8z
UrNvZvckRQxqi4NvvgIRpcIObi7hWzBg/pM0IrwlbOo89i72fMmSVtMHTJHIYKnd
tw2lcjOS//u4KweNfFp4jaEWW+Vf5SlAC745FApQgcQKlQxBOtcM+EKsumSyg7Fn
1JenaNddZE8l4jlquwBxH+KTaJqjRtZtT4cjB0rLuHONOa8Dbzk/A4goo51snotr
TFnOfK2rL6wTVvKv0ChbWPRdspf5CDbuy3bQLfeIpMd8hA1D+JOcy0fuWNs+rbmc
8xlnQmPXKdyNCA6pYGTwjBEhlWdfVxR+XrxJmiS9y9U0f6AGqvihG+38nJrlPBl7
VprWBXU+SawT3J9govIYsjbhD8JDq2pIDwyYC/IOoDzrbfRV9GmxLcIpA8vmaCGl
dtE6lohVhYb9cw8BsqeGdi+4YBGkNVn0U4zpyA77ma2Sq2uxipDw477jH0eCwCsM
TcVQ6ayQ4YkmkKUYN/U8tPGXfFOA3zwJfjsH7/phoCXE64MX+wee36Orb7s6X8Nj
gm1aYzXxL2kfW6GcLXGX+RIXIW186204deeU3q7Xe+r4GBjReVXvUGOoS5Zu8uWR
AyjH6IOapo/Yuv4tze3/bjYMP9+9lT+h3w7GJjEmhvDD2GFy5gZfEIDb+TB4OKXL
2el3ZVr91jOE9LPTsxU3bJP8UOF+QbaMISri2a7ZFcAIjm2vEabv1Sab7HR/4uwD
OA63wn+VbT5JH4BiHF6sskT1tA2XFEsCDcOOF6jY1qCfDNf97CYgnRkdG3RDpPue
BjtbgnkxWWQsYpqMkjzDtWhMPlyF8mCs203x5Kr8qhse2Lkoc1gXs3y/T1WnzzSi
3GITQ05SPz1zVrFhj/5M07HCvokFMdTk6j1FKIxufY5WQsIEodCCCKnmJviAo2/y
dUkslPFoUuadV2yaWWC8aTwIFFlqXNhr72nxodJhdKvOZWvRXMx4OIX4UmybYf8M
cmveEFPefDiKy+D/V4wsHu/dkqHAacb1mKsEevSJM0MhATJBhwUWog7vKF6oINX0
bJLl+ZMANvSv4x5MNxTzf3GvGdOjNsUcRsx3wQAYmRw5MpJ+pXELVu/QsKLY0m8f
jnwXQroBcTmfD1t0NK19MES3L620dr0SDjOfRTvlqTDlXEAZjPrK2K9KqYtt1taN
LzVHJC9uLGecBBYsvVIt4goCozhy5rCfDPfNmS7IBFcYJVltcWVhXVuVdyeyx/mb
ql6vPYt8lF1eu92cvwKnJmIW2HKCwVyPIDUSyrNGVqG6hTTsYF8nQyCeGEBkLlPH
hWkm3MC/iUMjVsSZjRjHqxsau4qtSqVLZXso9d4V0cUVKVLxZDwNLBaWkvcXtapC
l5ePrOPOniNsgsKqBkiAZFZeV5t/+3pczr1SiqnKWOzgIKgpdj90V6T4erWCk50u
wQa+I7/l8tEf97K/O6937eFxOIagyPdS/7gwUZFeuelXgmX6I1anTi7nbIBmA8UU
aGncDfgZOLeLUIRBx9A71wLzttP9XTD8K5hPJS+5jzhti3oEYwgBin9ZvIVj6JPp
U/fzGIjBqR17NeuEdW+XoLg6+ZYEeM9GlF/EsUvoDQUhC0OSsQUhEkuDLU+GF/lk
2hHMoueFDj3h6HdTCVLsc7hdxwhpiB1Ji1v3/V01o3pyJZTptqb/4/30BLrO31iF
r9231YMCjr879ywUUQGsv/ejgUBuQF7jTtGZ4SyjgDBtn8b0+atHMTd3g2HuMDIb
jr3xALEGUBlfqTeOr3Bsq/L4JfyK49x/aoPtnPeEepCgsGWmO3I/9tLu2x8eNWYp
Sw5W8OKLyu+MPxQ3pMey6oqinVi9Oq/aBjHM1J9GqZc/jXt/SWIgVU4qKhdI+AGr
yxb3aLORQxNTN1ZVh1UlYknkQ9G3a7r0nz1iaiOwtV9GG1/lkgPHj5mRG3d1HgMg
IQN3n7IE5ANP6KQjQfGbzH5RXN473KB/b1oJDiXcAhOJxNZRdbIG7+8snndXwplF
oj1O0ElhsoDQ2q5VEHxTeGJXimRGzEQkoDuPAdTen+pi30MIx7rxbU2caxZpN3pv
PBZRAq440CP8ndQeJVwYAxPZFdsL7b6NtsHeCeJ5P6Rhv2/qS6MPxHO53QDAG7pY
6xZU5+XLi7jqb9hviCM+mfCjBZC5wHFFvXco+8FMEIAgPkeUd+TOHJ3Q9kVqfbrP
4Tc5bids/eD3gf7uD+EN0bWqrUwzLNuoEv2wRWD3vdSg39uXeJxHD23r4j3oxNil
eWarEHNIefVRe/WuawzuDkihUBh9+CFqOFEHlK/LqAHPozZ6UnYfBr8GMFT5bJyd
THlExrpaNjsBD2ltn2SKYrFi1Wy2aHmX/FRsqKGJJ2lxoGrTHIzjn1O16q4nlACY
Ieks01QvHRJooVec+76/75fvKGrBZdYpSVZyBo9tbORHX5+IO1edd1ZtB8r0+Erx
FAx8qUIQhhimKrBKYnuzVwLbrd8T7rfgCZUR+AkCL6JrU7dRHOXut4Ged4w8Hzwr
m2o7Z8mbMMjcBJC2sutpp9JMX3CTMpKhGWl39YlLRo91UomZYW2MxlcR57H/ei1A
1xyD65l1OQ2BYl6cePEhiXAU+gj+CFO5pjktK2hUrNKApTASSINDfHLYxV4k/ZyT
wsLPKoWHYR7fzGGJmfFYwJ62a+HPie3zlmO4o5EhkTROvVRhz5e+BOSmh1WsjQJi
eMN/dOdSKdjexuX7CzDVBdg4a+UNbrqkdGTAh026qbEf9F9vzJLYjzSBd+YTu5Pg
xXyZAURmMg2dbphniVDYV4W2l+MWo6Jb+Y+Zwm3WGlPWdL1UnAgbFFLKqa2u93+c
dpQ6KX/RurmjXva6x5HfGmKdk9NcI2wUw47rSxpJLVogQXKLmn4MWIKmm06yvV0q
W8lePReLhaRmChSV2iPn4qyTQ6Pj2djaFC7sQhKKPhOgNQd+dAnXOYlz1fv+mkdd
qlcA7CWskQ6oXhEJLvRcdLEf2vn7jHV6eR3ZekEsBa2HtRDNQ1yhmgtUImr124rM
zpnIPEl3dL8fFkD2+rC4ub+TIR2OwFfXpGHua/WsCAdvfLLShVa2vjFpjNEGh7hP
yQO+AywtopOChBSb57Nh+EUAstQ42NMr96ynpXHM/ftrG5/iIad0uroP597MbVLN
rfw1vC/wxe5azidhhOJJwlQL5QU2M0hdEIYfRsVUAWmaWyO9ABoyqUEs8/P3GrE7
Se7shdqwvPotZSeTztwV80oPzwUkKDjE2mTwdMcmtiVTOuWB85H7bZ71ALgV24KR
nq6ucSSmDC5ihJRPkkDr7cTryzQMf0VxoggnqJZZthryrGKFBXfamvRoYHyzO+EG
g/lvtwQwcSHc9MTxCaZn3P6Pgorrjhul5kD6rK1om0fUr1yG0noF4eMuhV2z9LSQ
JJpSUJhGdRDxPdMdnmTmfusv5L6j5pS2XDCmyKcgnoOi97l8CsDKDUgCE12ME3XG
VuClm0FH7UjZB2Q6OuNnVyQ1kKUny83DJswVviWP/RMvS3Hee+WJDTTSX8PKa04Y
yXP96W3/ZDmF/HbY247TAuIzlj+q7y/+8jFsiiqTkCOFS1VxHZCt/OjIkz/1zJZ2
8BS+sECzDPmu5TMhuAc2j0Qh5aklkeDjC0O+P/KpM50krF5P73dgnmFGin7dKmwV
9QCChgIY78c1PSdzGXQUYQ1fRJb/h/ytSIhvcuLByZwM0LZ/waS4DtgKqGdWxeog
G0eqHiXQKcwQLk8MHjZGXsfvOSJ/xTVd86ciUey8ugrMVZBWg+o+2CBY1/0YfCc/
TUUTFGDtaHxvmi6QRU6cavM/DzBVbtRBsXmu8UW2UC8q3VLMt1LmSQ1MXO6A3Otc
ovK5SKE4Och/bL+PmiyTEdUf4h3YSAPuicgwPCsr04Z5ZEIFy5MlmYZJRUI21qWH
yFLgzb6KVPMZjONAOgH5U/Nd5dl2BUSTRjSzlWv2bciQ+E6YxZV/G4k8Ezf3clzh
yJhsUc9Ygl5Z3v0e9j9va9FphZYeTNQyb3i4kYh/rAgU9OhRgsHQ7mOfZp6nRtgk
ABUYPz8w1VIXqzD87b4LomPHVgq22n/GXX7ofjo8E7MBB5SviZJ1UejWasxkKgcf
B895bwChB7/UgtwZq192aSIaZLx9evGAJK+sYJ9kpzx6NGqELHjZit1lIA5TFgQZ
/+CidSxqwpMWfxnaPqY/nddiZOFBb2Ob4YWVXsfuC0MQsngm81ii97990xXosraw
Eqh9q9tlkm9I/fDwJk7am2lE5lu31TqNBm6HWPCeJArj6NDXhMvtMDVwPDx2OB4/
z+URVTBb/KK1S8nBA0JbYomiAjEIj2iKK3z9QSpL9mcbU11Gw/vvg+9ZwMR0JvN7
9bluitK+FMjDlfMrNRi7c7Gu7UfGkK4pdugR+dny69jyEtx3cjIVFKxlQ85nIrCV
n9Dq0DB5XYlEMaVSiNBc5XmEKg+W0t8s6hKMPDf0zlDZynwU4UDXlER0AmmALa9F
zBBmhNyTYK211l6jewKsW5NFx2vJVXWl4iwCyMeVCEm5PEjyC7xrIinppoD6zWrq
KdCcPE1J/jf5Qql064oAZm07zOkz9DDysaV7uGAy6PfOuHJF+NhW0x2sod0yfUke
1R/lPhmmonzLFHuk4RZg2YfdsIkMW1JJMN+0wKB4kzdSpOZ+MAEY9YrVkOtMXZNK
UMqVP0RBYf8758OirRdVErw1zUz5vEJGOLJDGauYXBf3rs/ynmtLHFyXCRfWthoK
GaeZ4NoGvvipHw5V+iD5u6JaOSGObDnCAixoBKD7+QtH1HSsV1cA9l/zV9a3+xMP
hVMk5RtdlCoYe+hyaDp4lm9gbqGz4om4Mrsret4yjBQBPS2PcfMv15fdFM9Eoxb/
uSO0nLS0+csqfsygKKsRNHJxhGje72NlXjtlWWJ9AG9b+AqfYdcS2U55eBAjt2dZ
AQoExeQFQ+NiigxpZTkkJLAHqcNo8AjhrG+iOncEwBx4+bi0utpU54uXc+QI9NLo
T3nODW4SlV6WCjNyVAKrM1tKcXOrFxZutBGaK3TmyrmVl2w1nECwRcaeTrNz2Pmb
7b9FIoqdEpIm1jLR/YT4TaFudLrMThi6jxjffyiijji9DQG3FodCGOmlAUs9wQRO
ePpUJ2cb+lpLdF/I+L/TsGz/JuGBlzKhzLzoWa8apmNeYbPcxhwNn9K2ygYkwCNh
v12DYD8OJ1EqyKGzK/JiAevOiCeRbiHfQGlnjIEv2tTUmtqip2bpFXVwwroM0oNG
H5j8oFLCASV8bu5EpYMB4PiuxAj2YMHXchAQCi1WdqTdRx3Geni0GdEw99Riuxkh
VY3KF5fZmxFsGzcJe3FFL7NvId+z47myAvNLY1GLLJfLWriB7v/p7F/ICf3n2cKV
SRcTos1OmmegJciUZO0WQ74/AA8oq4IZDe2UlsXupALH+ooG7PolYAlayJdNJWk8
Ixttzrju/bf0S5SWzC2SZ0hKDK/X427iLZfi6YDRxlo8xJM/ltP2nErwcVMGNYiH
s58gweZYxZTvvOLCC1LWJZgKmECq1PLr9Gd9vMylVcsl6VWPueGg6HIPBOA/USee
q8Lb8+C81zmSig0TZrjI17fAPbCIir6E0FFs/uDaj/0vQYU7wAMjyYav4IBQHoo7
1UsWuL1EwOXtgaCmRzfUxam4VEwXe5wipO+1b7e6OwUGE63rdTwBMK41e479q4pV
5k8k+Yp1D0FZB1ZoK6B5B73gGNTRT7nVQ3zcVUxyjLRwfT5t9SGTeJRkeVplYFDQ
54En91secJtopZCVZ5F0r3rXy3hZzhHEFNnFlwa3AgkdTcT9skAPQ1xjdLW1dY4Q
N77NXgFsjy6NuvERjvpLHs1RU3wNS4VUrlyLgXGm6rq+4qvcuU2XHZ15MaBx0wXv
rojeokyyuSGymN/y7f0cdwYTxgAhyc1N3D4dNSbmTusAosa9UOEMVFnXD8R08llp
PawX82zgLO4qaGiJEGrHYcu7Ar3MRWTfPNXmEkxbIGDJnwB7hTxwmQVl9RR1HjHo
YEujnJFQQXRn1YALXBmEvJG0DBsklTOFlqbXQRmPxRkDTUzDsZD97L1V/kz4M34r
WvxRxhViiA4H51UCiydVfuL4TERjAOFN6ySSVstwwzBip6fj+Or8aIkRoZ7L9aD7
1wpzcvChESvvX6Z9lQ6T+4bGDh9MsleCO86uIJ5WrLkwCyvcRm+jjsIAqJgNi9HM
4LI5V1h5FkvmzSa4EOSIvw0EefhGWmqEIkbDxQi4A4eddgtAOuxs+4wTD8Jq5n7l
UP2m9eGWcePJvz1YaOXegxd5LNZLFU7niAtI5quXGp0l56UTVgTPYgx29ZKxBWjR
8wjLjk2BHMf3ArXA4Bz34zF3mdQur42/yF8Lxg1omNf0FQzxHfyevm+MBDG6ITXk
/CoUvfN05bJ474rL+pY2jCaDqjhudg4p0bQ/pGtWrdG+6+toV10KGxeTw0Q+OFAN
BQ3Hw6dSNc+zVfeh9HID/hQBjOMgVpdEmlhy1UFsi0/OIc1qCy6kYXlgnbXHeijp
maOVMbG0TNXUP9DZhWZznl55rHEEl9ZLSEnDMji4T1fFu2BkAJk9FRekSLRGPYPu
UuX9LFbBHTcCBlEU5Qw+fnGLzTE5xmLNBawZbdhbigX81IuCqrQxZvfGRnLJhCTC
j8xz6ylaoahXOiE0HrJBGwRvDI3k7U7XjbLSjj6a4DQTpY0BKuE2qDGAvtfHKECl
d7cTHQ6XxpkgUlB8uJGT+Mz30NQm2gGG/0e/vpwJIjDV1dtR0WjiEd0lsuuZFw+Y
5xn7ZmUv00gBEoysp0/24STCvbO8k3pwqnk6xVdE66XGRKIGdp9bShlLFEbu9j97
R/AlrTnYXmIg20KKaDGOAbE+MMmpfoYBK1er9NVsO6MGy+ZDfiCK7LzKIj/c0l0n
KyyswQhIN5ib0JvhzbfQA4iJtv/vg7VOKBVAORsY0V0d76LTCTE9QEGR68JSZP2p
151jYNomLQC5RPTUvxf+wfUyjGmg6w/eGHet4kQs22bbvFw6z2uOseTZ+F1HJ07n
XRUj3OLzs3iAXAgOZA7kjsh5McQ2sJP9SJ6GH8nga5b5ac6mgGBHQwmFWkRuwnN3
zzoYS2Vwigb4YQ91r7I8xipoJnUjpA08H3+thp21xz2gwDvVGAGF7/M92UdInVt0
zy+gDiEXHcgUBwRcI5TCt5tmKKeNzqZeMRLgtPfXRW4ktDOXZshan0WHKsRYvZIP
xdhr/BfBj0Y9AcR366W9q0MP8Eg0pQHi8KGWLPne61sjsjksmQkEhVk5qnDiiXZo
iX/6ACaLQFGnirk4HUazJbWt1+yrVpRRYaXqofy7gdALFhlm+352ftndiSDe89MA
Wbw3unG62RM9CNNBkiTIbCu1HsgRchHqHkXn9jzCzPyk7Yg2dg9/F582QQ4Br15j
XqapLnFDx3Nb9IJi8DlTawTQf19qEpBJ44SsJUCuOSVP9i7Ro5Zi9FdFkLq8a8DY
xKTKqxPhKS3Ls+XgNonCNZ/aWjXjpzR4X/OjfOXkTnumSxAXbRWqRdDDgslnQqMN
w/lbwWXlI5OPM8OD0ywZhDkjBdbVbgX+fiU1pxRwSvlWp+96yY+QfHin5w+9L0fS
Mp2aSp/2cMTTVUpMmVcXlJkZuN5JiuthIPPNO7WpC0N2StnuwoGFCeL5kofXzM3T
rzwW8fM4trslLEEXz9OOKM6up/hsGtO3QjnJUmXUR/k8ylWfuBFxdaIYsLJiFCgp
QkPfxrmCXDXvBRIONpnS8R4+LYxIeZSAYjyhCYBPtr2hikNREzvwKQoIy/Nrudeb
ob/H/miSBjHG0g6KYSRWfCXPft+xEYCXFCvdgfFgUvigR2HLZGglFQ3xfn/7Ev0F
yQBxGKWp3f/Gy5sA/po7DS9X7pIW6CL85sY28ungt8vRaXFCRlaGP8ABX3AMTIVy
iwC5Wlo5e0FE4FJ+0Q03z1T0IixRZYbkiTxjomSNqLGHlQwUIkL74paPs9lYVg4Q
RpA0BJDq8EokEtYCuXuqK1URUlsYjKGQD7v1p+UtbmYnvsjsIkqdkgOUL8PnVYx0
noHLkGf0dVCUexbFeGFlUuBL/OrBtznY4ARU0rGy59jfxrxrQePxXhIX3dlOnKuO
uvTR/jdeCtpwD1qejXeAGv1glEyGerO3EPTaELzm+6YPcdPUiwaQ2XnnhRGNn9kg
SZyGAZ1Wqy470WFJlkRrGZdrfKLYn6dLGf2kdVO5DXIwEgtPooZ10JknjGSBso3z
lLvm/siYNDtB2745rfqCvJUmNyGllf1WTFdhuEfIy7EeOntBshYjIEFtdIZkM4RL
JKxpZVLNtjyJ2Ra/3R1sqnXBvFeORAnz23gNhWUZ1tkwdiV63AFg9qqLhGqRP8kr
KNNZpiEaPnsBwBMwgvnoKCXtZJBtr2zhSsYSSnJ0A7UyPPT1n1bRLMMFJCUSwCPl
ipjr9XAp/iYdUbmL/ZkqGhMO+nQd7aHEc7smMRQl8E3mv4fnN9hzAh5ZYoEKAolJ
09LIKZmoIvnOt5lJoUlTOP3P7PD55DZc+CaiQ8PdQlOdA1JAKd1uCjqPRf60xY24
5Mn60DNdM8Fp6KFVOysR0uqju5QNYtTbKlYyHl9KnNgMixI/3pmZqdV886ee9TRN
XpO5ySIFT2C1CSnCJIN174rr2wY4o9N652iMnjwRW81i7yH9dS2Q5FrYZCPpxr88
yOq/s6XUMH+HtPFgsbOtgslfnAa+gXxlv+m/wf8vBzlkyWz66nvvBVFhWDG0Jj/6
oBcpUY+dIHYJSpYv18pdmWVHmAwRNHWua+tlajiwaiC2JQgVTeL/ZATkHpiXWwmN
gaIxEBjo3uKS8d8FWvWlpVdk+Vl+86w2gcF5kAcURBsuMpM1JTXSr7RBBS2NO9C2
UaBw4YiwOQArH+XZm5SV6oYYEG8IYaFr13BAElnxcitOIB/36IAi7YIPh13UV7Uc
e8XeuqT1OKujpbsNhepBDmnH+1jH+P3G6hy0Lzj2rCapUIKv9KmmOAvbF3ZEPW/z
SdLjVDo3T+1beObs/+7ZsHsCa2maSevewQSpBY/xzTJBE+cLpxZJmRU4iieH9Kt5
w8pgyY9yIahKimbDBizp/OlWS/6J/yUVryevST8LXkF6LdVNCULKbTy+CACJ7IwO
ycQeHVfsWAYFH4b2qszTGqR1XfkCEx0MicVQzPnINizQUrr45D0ga9bmehlBQADr
8hYWikHXZufQoq4BQKs6xSlKf7An0VSJMQG19fuiIZ6Ar/wVS8ISfVm8B3/Cruc7
xSxOa+T5g4BfG53XFMVReVC3vHu68P6AuTZbQ/iwS01rkwD6mO7IvCvQg7vxg1lV
GG/x24UtNjBq9jqU8vLtyg7smEXVem6Vbk6hT2DmFXs+ZA8evhrBNZ830Q/20WAv
TufXke6/NCofdlDlqBo9Gyy97YjQRJ83qpO6GxeQfTRv7FbcpZTCtKsMclwEQvrD
p5ewYx0MI0IfYYYGuH2YqUCTHdMrzSxOgbYgX8FtBpLg06LvxcJYxhVqvJHIfp6x
SffwZtS0lEHGp79a3pMwBc/wE9GCnZ9rpNh+DW/19ba5gOII/vcNekznuFenxllb
HV1V619NyQRCWZ0j1Y7JI+taPBXHsmF7sjvmuWjBwyzIiYkYLKEgMH0J8xRlzxQY
M3czvuvx/NUnpy0p8ocfqV/RnZlxmHHVK7aa/9Z6euA9fqDr3wyy7hn7SlyaujEO
wOu6P6ACwKta1CgD27912xmkR2HGJxhjJzOavUL0hQHzHpV7mzFQcT4lt1hR9Uhk
E+RHNNFum4xD2AmKsWUBa6UktLT3N2Ma7OMlhUsWaQXq/fVQBzioFoMGdODo1W5V
z70mBvvaFQvsAogKGPfFaQ/LqpPH0TyoKVWTWWhsNHSJA9bxiwQqoeJ0e5IWZV3u
4KaElyG9JMxd4AJLvbp2/RAiQOdxJPLnDo7rQ3+jMpXEg8bda6ovO3ziBhPoVXIL
3KNMClRZoga4JnmQsrcZRvI49es4hyhoqWnOpYfMS5rvgpEXuO2CMBCJHoNJGcaR
FBFb+h+V1lrU6aTiZRez2vizKLmVMsNJZGSsDwLjOIXVyGUbrRYjtU2dsoGmu4bn
tVLtBDBzFsI91W0DvSMTxvEEW29AtNj/zJIxbX0ZUJdiRXXQ3Ph6dH1/H5J7jbEU
zx1bTK+W8G+J3eDI0eyS0QwOQ6d4jrmuA8Xonmt0QeyAFSyP9r+Ln8Vo24PGmr5B
ZR4QRN9BWAQ/9icF0dhyGizSiEnk3pHw2dvM1Wc4ZnHiUGgvrsDUJQTzUNlPpncL
e794zAMPtIKT5N+5xz1QSgg5dvHaYx4XRlOMQik95enlpspX5iSlx2RkxL4bTyLP
DASMyGIsSL/hp47gCGlF+t5Qs2wv1rEOgf1fyL6RB3CFD4ZBK8x6/jHJibiQ9POD
1vcW7KPbrOzXb9BYJHyPtZ29yRHVv7Yr2edAvLc8XxjNOwOib7Odnyoq0JqJxXZY
LnpIygG8Xugq2nGmtKJ8YovNMLja2M+d9gla0Hwrli1GZYZ1DFOyRur8Cc/3Ixcr
PH6m4x5uwTPalsS2wml+RIRRJ5R2qV9SR+b13+RLZ6c0nnTXuTODDvAX4gkBM38x
9qCF3KBEeScLv2t5wLYESzQ6RGJyep3YeSabP97v+6B3R7O9zvqQhx+weiyiCH+L
wP2YpU0BxENKNedKipuOnabUb/DV70sJUXp7uBFEpvrdM+U5VvxUqoRj+7fviqa6
8Tb8ayWQvlvXF355A15KXusOgOuklX3eooouKcwpuPO2M3AyGViI31BGbYme2fWf
i3wPrdQsXxtq4ngDpsMfJ4wWUbIw/WWswfC3fD+ylkTrt8QK1gHEgm7xtXuvXZuI
XU0Ycg5lPmzHc9yZ54nm2fCvWPGZR6dT6mqvVwDBCeMXeT0lldpLSkF/8Ue5/Mfe
N6tcYq+Yq7tHw3A6eQ/WN1+QwR9umJUfxwEaNGUoptnfKxTv09pOIiDfFln2q3dd
MNnwPV3RHDjfein/VoqeaWJTTgkvMP9cJtdUrLrR5c/0h16y8R0XYPIuluYfgjzU
/Zt28DnXVNghlECIIdFmzpcBk4KJwLF1arVlFAdRNc/L8JH9736f0hSku8Ts00ir
BWAdH5D7PFcIxqzN7aGFLxTNanoUFVl00TiDq4w8Q6MHS0cG80Wu71Yy9o6yJlu6
oCZFje+xH7hMd07F1rQk/P57smdJF4q420bbrl+fNSX+ZlysDsaw0DP790l8Zs4P
fNFBMZ5/DTEGVuL8ZDKSY7o6ihbi9AuL0BwUxWR3reBRI8BiQrkW7mxE2/yjFNl8
lGVXG3H6EdSC6DKWxp19gY3mq9bey2gGjyhjxLIx8bvyZhvK+OjI4tgMdrps4rT2
K4BJkxqnr3NHnjYCCHSRz0wmEyGya8OiCnFarVlk5jAMEnikRCywlLsx1ffw/g6s
sKv8XLwvRJg+i+7luEPfpRPAOOgWtP3UCIFNOtkJ0TOSf6iJ2Al+X8XAia0uFftC
6uv4DzTlu1W0mjhoZRtnkvMY1QK+cgKoKhPIcAe7sN5AjzXj6gIERLcBaI/bG/YD
BZRtmPwSdjUoppcRxH1AyqUhdwoxgkhFms1i6Cp18odU8LAfrt6IigwoRosthZY9
dtml4PFUeEtJGwma0BeR8fsbFeYTBjWIQxb7oKcY2spzb9Z8qQ5rQbry1Rjz65Yd
lO5mwUvSGZucY9VVraNwc/FCdAbaWQxweXKuo4iCU2xreZMSEef8Xrd/C6I1sL4V
PjYt2E1yaNJM2S/Y/ViP/akx8fTKya6BV4e8iEtFGClU5Z5kIPGx9WK14fKvWU9Y
Xo1Tbd1l3GUtdcCn3/fkKbNJyinZGWvDMD6Tu8z1+ALe1tSb6XrTySrGcbwm6xZz
oS7BOZM4JV9EZBGbUns5CdullXv7GPS62Gb0Ga2an5PytWvd16MyM5qqnJe+8WPq
ZIt9UsWz02UcoygmTmz0T3QW4lzvIu3LQi5ECvIViSFiaH0nmh2Fa+TgOQ3QPTEU
xEc4uQdBVXNnVcn/NFi92wFXTCuS/5wU6sVqAKywmgJQo7MAVBHJ8LubZCvN9Yqg
piaj21I7u41anFtqCIJeeia/zZPU6vKcuun5qg4EU7v0DZvwfp3/oIDV3R6ZGqvz
KRtijQPedKC1q1gaLJW9Q07AXBrhEZzru28OAtOyS5ATieGeOpI/C7j8CSqlY+xb
DgynswDsgY2vIYzUi6fDsiNPPf9H5uQFG7eG+oYwoFJ+FgS49P41ZlHGZESuSg7X
AVyRWRIFOh18/2FFp8M4DLICTL9M/tpUh0LlnGE9lvCh4N9RtwEYlrdUAYiWIrNV
aI4rBzRQ4EXYwcSVSXn6kEdY6rOF74W20tzJh003WLxboRWGI6h0AaDjJQn9PCjm
CtZbCFvZAvIplAvD0nM/+oXZZGnvU4cVrTl92ZwC1lEIizBFwNcJET+9oG0+IGGv
1gUWv0Tw5MfG9NbbQLbY5eW6Eb3zJF2lQPb/9yUVHLeu0AsF+W1DnWw3NPC0f/UA
DhqB9ohk4G2e7169lF75KvF1Hrfde28s7cb32n5NadvfQo5Q0rb20h0O5gm2x8ie
5act0W2Z3apgeZX3Hzb/xjHmbNcxLApR8In+k97uC2StehPCVqjYOByWh+gXVV2+
ASK6iVmgqiS8iio7QrFeNsWBnVA7hnlwzwckMRAexOUiVmmsTQvoUFTh6zTn1Yq4
JZT7Rrd8LcG3oeXtbDDaIJIa19mYQcdGqvHa3GD8x6gUFEJXTHk9F9KNACKAdX1G
/JZllzHKEEsV2TGYXe1+LkrTQgnzHC/2nGOXBkeXqhTY52Us4XvZTCdxpREpUP5F
ICiG57vQrua2tutOke8H5peNPmwcwkSB45GnF8pVxIq6DKKw/RAfuZ3acWQ/3H1H
4se3w22Agoe+aU8WjQiwwLptn7FUsQhD3smlYJpOjGX44zavhaSiyLU/e8N7aUBj
lZTod6cPYDAztphH6WJ2xkVpUfJWYu84iaYn3mthEzW4azRt5lA3fE1G6LHwdSu/
c43SQoseZ4W3UfpUDyEF4NdrctVSznHUxfNCAjUXjfaMRW/7oueOgW9unHuCJPjE
mUeuFDVjuTtMpQh5xeDVEK1jKunHnrYnfdrbYEDhaR4h1voq/AqT1oKf83Yc6FGX
xhOzzn8YZI/y257Oejf/7cPMpVajf5ayx0hLzTCEewBdxSFktlVGlrqIeDjJQfVx
t/owfjC6bSmXubFZRqoKZJOixeoMJyqhad4pOeU+xhqgFswCEYLGjylUoka7Y4Gy
03LeZP/SNKOKXGJUAxRh8xZqo5RXM7mx/AMjki3LlXafqeIU3YFMGW60ypp44HeY
zWwbUP49UC/G2XH9B7RWQt3qtzdVJUr3ISjZKSvCn1wJuBgWHIovlaCE5HHEKD/o
73enYrXj+p5mIA8Oy7OcjKqqwusiE1RUA2KBz56w0ICKBysYYr8C5FUXnKMVh9er
OrRr+odn93OGxO1cKeqlkxXKEcrhzUK3g63oh7lt1Sg6pQTvwFN7o4wsbf5dOExP
doCB9rUjdaeNrZoV2JDmxjkvMIrfZUnSTp0qzLogfh+QSEOxVe62JfPDiGPuke3C
TYcyUUdcNraTU4dazv97PCMtee3z9JWuI6C2qvQLCEsx5lDYa5kmgwZ30vk8s+r4
rE9gM5rx/s/08ucDKpmjRTQhw4L3QWSk1oVD2ELHEPHACWVCbQynSu0CKLyZrDEP
5EIpZAfAPvIPmw6rI2BgjtQ2S+TbhJugqKxsNOzt9Jfl0OISVocg/OIXXydZbH4O
HWOZv96CN6H2CGTApG4uKpIPM1u0RvaM0YWjIUYftcuHnh5Puz01Pywy5P/cfUmr
D0Y5w6IEocNz7111/QhWVsqihVeJIFaRo/BoeJleaBb369lEhJZR404P9Cz6ZmWG
+ifFPdwGgvRI4D/xKX1too8fEZaZic1gewAmyRT7i3qT1puSHzBBC5GZXtWWuHA+
w/vnr1eRUq+D54XR4JyfOoTfPutKmagWgzoAH1WvUNzChdG9ksBo0OPOmdORLXVI
UdMYJY7v/V5fwYno2F5BZQ6XcohsLnB/Ii2J6Kls5k31aYfNn/vtiq8BZsaV5Mhx
HOLDppDcIl4076WOl+EnDeIlU6k+DOFrEpsD9uLtlnMnJ+yzaadxWjg6IlKDNLMf
qP+bKIww5LU2dV5vUlPRm7BqsFunw9EYM+2cpDAVXW3/XRVuBeZEAg1bnHgIMfkC
CGLELAoAAUOTPM0YxAyY1ZUYZs774dqbxEaDVJFSeQnReSSqILp31rTVa66akPqk
2jIm09cZqrfl/6k1BhS/3fl8hwBdD/xvvZ/YarhYqCo9OsGEHPEbjTKcc1+FCkvo
79BZmERUHlwIhtHUCHsr/nNj9o8YWy+qtPXWCrLxBdDvGFH1QA+zSBUeq8lgvu7z
h4Rj16IGOJFbNWZF7XCm4F3cFBhIGQFl1BNkDFpkl72gtzvKsmgoIjzBSluYfXbD
n53VUpQpcHfPThZ7yCjCWQ7DzcROxnieUIa15eXM7xZ5JHdIDL9XtBV5YT24mZ8J
xJsMlIno1qYkdPij0X7VLaGvlXv9RdJjGCGS8jq41NbsudgEJ3AwPzd5jujrAnor
Vwto2/sLjJOCVyAPLjffibsRmaIwfDM1meEx78n0knV84FZbAg+JLA4nj4PgBLbd
YR8TPy/EEHTXAMcCsmFuN2sXUc7HtxK4MCtbTSyEVZO+4BDVB8pMw4jgSCip0kZS
dRgqBx77+OFhiDdpHlbgnxviWo+h4vPcKE65EqaqhXadwErapndpCiqjEIwgy31O
ZEsn6jh29JRiiHFz8SA3ghL+/Vf8Gw6usrpS4XPqOfk6MnT5zf0BzK4Cny6Nmft+
jZuktsW1mU8ZyxTRc/8fDQBg788oVOb2r2/uNh1JimD6DGpu4HNwsKEzmyBlQXz3
i1q9MJ1bfoYfKocL/92Al7MfgCtL/1JgZ84EnOuaumf3w9TxLBhWHz9p9lxqFuIx
i+rGW8uIvPJgscnQYU7eWmID2WejGKlSy3k6133k8HjjBaXCayszl9emogATRp2T
+nYQmRH3c0WjJJJAhaZriRpvSxpup/6AHGjXrjzVtCJPc4uSz5dc+NKasEJl9GQ4
1HCcDA86JzxlAJP96+WO/vjorKLCw0/mz48NcheXjiuwWzvZA8DtjHSD4l+zOkcG
R+lWQrf6Cq9B26Rv0PBKCN5xUfKqtfiXP4FI9hnzI7OAhagAjBWr9MQ041s948qy
iw+v8QUrPwGI99gh+PFiUHh5Q/pKY6CJt/6g72TuVngVexMyei07BCiJCNowBiW6
0nD/QYbnwDEMQMowfhHQBE+dkH6fr7LgjnCbXb9x3lEK+JSVy2K4KZPjCjWuNOqi
435nqyciPPDzmsiz+87q6d1k/2LoopI5GWlzwhLY69mngVfdZNmU4OMd8Kj7FXqa
n3scSVCzjXPSnSSYevuzBx7Q7VTDyKMtmIZz/GRbLlHsEDTlBrIUnBL3TssSyJI5
hh9UzI8NBmhg/IsUPav6WOGQ5ZOGlVuJb1s38sF/L0SFfivWrgRWBVEt7riXJRX8
jRGu/5QS4V/h7VmiD5X0QgHavrM/h7kfWkBKp+hZiK4Qb0xvYckgY5HSAZvGXhfQ
tdxbwpVLJzxDZOSVR7bm1r//9YUWUZJMIRpHrrNfFOYyuwoJrR0frbOTcfHl/1s3
OyZ/YuMOMz5pdaGMDvI5kFYbRDt891ny7lRSRCBiWVMHE/YZ8Z67Gskv58TTpPIK
ASomxYF8hBsrmHTDcw/PYfagrDuF0LlHKja7qH89jIDCuMwW1Aic+WqMJaxAc3KB
zbt1mmSCfd7heULyc2JSHFfnoKeCf5yILIjC4w8xZ+hKTsEoj6lBdJ2yWCG2mTCI
H/rdt5GVnXZZEA6M/qjTb9dJOnWHUPdRFNjZ8dyp2Sfudj5wH1gHixFSggE/LOZa
Gz4cTbkyWu+zHr3peKpvTW8oToBIHHCoKdNk3LDO1UvCBhgPRttoSP17/0GfFHB2
mfCZbTme+WbK/6DSwA+mKSgid/12xX/3FDVuIRUd9FCCLLQy95kqYmXlXIEj2sm1
7/WPnTPy8oAdyunodh9mBr0O+vk11mT6FX3P7y+iq7aE+0ShYakVUEQEgm2phgqq
hVffU3LFBKd2IuJ4zf5BTK06NwaVLt7cHAVaHb5yzU0IkMlw9si3M837WF4hb9a/
zNu8bWcaPsNWnm8C/Wh6ld4fyXLgp6tsKVsG1t8f763ABc7uXttpyWCjJqDgaj2G
Eqpr3bQMrPLvitJAYsSpxwvMBfMpJRz6q4HmlAVZKjYPLa94PI49QrAmd94RLnhn
vzZgRldqUpTGxUM0JqOV5Q9ifVXSxCJClNNcR22fLxniGm3nileDphrqAz/piVcD
iCLs26AqdYPT/8SD11GfMgUfjgDCn9erY8LaDUU1RcdFum5E/geIFHYN0HL1hLKF
h0VuBzsWnQhmkoMruwwdpfoHUun6wy3uRHDoDhp6VG/sPKqRIxvmZMEEQYWof0li
COjjLJN+3exaY7VqlkedB6vynLw1lVEsHmY87SP0iS682mAnZeKxWgioRLMZcbkx
EyW85B04EuNI4NJIJFxTCF/x20O7TKUhFwqqxk3HPMO5j1MQfgo3PMJkBFlDZ3BS
53sDi13mM8jH3wYUBF5t/LgTyUhCSvQ2jFVdMMgik+/Z+A6+9s+lWSAu1IoZzQCn
5hcJZY5PA2n1bxFsx2gB7olCuipc9grXmuWm6AHBnapmrta//VDvPykY0Z5/M5qD
1nrQTd/F8ryK63JJr9/zgZMDSPqMB0xf3CCYmW4b3jgRBzZ0kuNU66e5LTp/v1l+
DZbTCxTQ4/OC4YzvkBI93fwphUzmzcdw5YN1XodGD4yF+OFerOW7h1g5zKYy1HBG
i+1jhmmpfncktnNKnaLotXezaXl0hsWz7VKaH6OIiY80bsHj6IghjWk1pS2rjaIY
DdAAR+gzRW/l45R4TH2lgIX1ebXXND1fhAFyj/Sona8BNoDN/lsVDXpkD82KS0Xu
deMggkJqeRgZONHPgGiPgnM4IEeVmZvfXgpN16qYoZTUnVYqVOBCwmkdGJCY2ONv
sNhl+UNbZ3rJ/4MEaqBUVEpt19uMCn8udD2uBCF6PtJ5JZDx1zIkwOa8mmJFYwpX
A+vHl0OdPGEZF2jKi3fgIVhFDCM7FGGOp/4r36Mp3maWWuUhS1sym2rFi41AGZVF
tqDa2g+njc2t/2ORHzc81niR9bqdVUoSbV5gaCP9wqHhA+WfLlcoiSulxsBIm51v
5jDzjk9dplyVoQ8qvr6sUI6nuQcWps7ufy+V2DeC9I5L0AhrID8jyyD6i2D6cFX/
DsEJq0GJolgsvrMwOs/3SZuhhSoE7H8SIYPlaQkJBhI+LjzQ3QWcr3+Yh+v1s+67
nqdzgIaildrDOp2d/YdtmG8FDe22rDHoadCWbvs1Hmv66O3uYyAeHwucl2VZybCU
ZjyZvLQhecXqUByQ1MFpC9m6cG98Zrao7D+IXRVLKL7ew7w1KrS6Vq27zMxoJRTN
Reo3DF+2zjOYLAlVtN1qncjFMALXGvaUy1cd7Pec33pLQMJFpJIWLVX+pkL3Xuga
FzPkKR3XqmjXTjpLcgQq4aOgp43lL3Aft/xHTI3SBKN3XjQOo6G+I+dZ6/0PGl7V
FFaEhzZW8kM/utdSqEKvx7pt1Qkgllz9UuuXbf9rCTG2fqEJOGsLyipAWecIdNm3
9ojp6tl1J1Q7v05IWrIkBMck39agvkJPQA8Tp9TwQZY5RVKbaY8Mj2gcBnGhyioH
D6E8t0wXoRU0eRryqY6/1v6SbbdWlrGFSRAnNrPGyeo6FUsyb/KTNERVBvz7/kEL
JkKow+Vk0wL8wS9LQJvpZ5TNWawvUpFcHuxRLqrbf5Em5wDB5TDikX2j6g0kIKIM
fwhfn4KOljA7np1fj+xx82hJeFP3E9B6Vq4LaguMi6UQDehEdurmaiNY0cgoUe1s
P05WGFkdvZmBbRx5VO9/XKqYKMSUMpkzuKOeTXriR87tnN3Y5Ks0cSvfs97vPZB9
VRxuMsQ17LVL1AF/0HgUv2FOAocWHVi6eX5TozCqRLCmJQWPdYOMLMxwl8lvzjK3
wbnytBRIjjCULHvUAKitPcAdbsk/shKcCaGl6oza/4xGVgmviWJ1rhlCYLqB/1FM
sBtW/6p/7YnbqCyMQ3pbsKdOVlssY09kYvbj6wyURwxyhiX8WdK7VHg1CyoWqiG0
mA7/wUpZq21UJSU7kVZ2/SohW2gzo8jhRP041QcCr7Zv4xi2Plg9qW9mMpUre/oZ
krg80SUBcqznZ4iHY+IZ1S8n9wMmWP3QemHAeBVM/phiFn7FSuxn2C/W+8WNKhOP
SpwPGMTfpDkhy42J7Fr8mZnKw7NkMj8/JWghLeeu8duL/nsqIu5cDzxOw7SXfxa4
A7lVVveCQ+1GDJvRp09SzojHqc3k2yQ6hcolzD4l5vFUEudkW3RUaNcRS2P3G7Cx
PSvI0B/Bj90vMQtFIeb/om8qpGb0Dcv19Srx36vR3dJQJfjAthDfFZ9n90c9rZxg
hZ8vmaayZT+7SQ10mRc+facVVGGMTSzEiYEnGIgKoK+eRlosuIPV+611CtXye2ub
rQZb7DblqrtqpLA1ljiQwvFiSqVh6h18Bew9uSwYJpjEAXkmEGtLtqzYbTd6OJ9j
D4UW77FWWyMl7A2RNDv91WuFw6YAnSo2CcsR10rcJgbAdK1t4I/pr6wf67OIkOTL
eXsW/ifKPiyeYeLcuhnCWixFHFDfbkQAK+pbm2V1Fo6aWCbWQA/Q/tBP+Cw4d5nL
ZKmt++FYJ5XHUe4C8XpQen8yduDDkAghSnUT5avBwZ1peoMcJjHg5cuw2MnPCMT/
SJOUPpVBnhTmCNdZmiU3qZjHW5iZ7Ns5hHl/shjUc/2sCw+SfTtqGoQ4TRyG6DHM
EBoNCMnZ0kgjGs1/3eFEZXuuPG5FZxU29XcXHmeImvuIzdWhMvnHmz14wZSj9Ay3
13yaBsk4cnNIl/aEGCAQmsBbNXBKLtNh6tC0cmfLpQXuONRe5Y0l0xJ3ZjQjV0Nj
MNj1vk7yulXZmsbh5nrpB4WeOoIXMTuoGwCfQWaZNJHHwF2+7yZQoLT0WQidW3Rl
Swt8TN1eYQT0rooP/W9iiR8iDA1BAa5d2NUC0jJr9YQtgii4i76pdHmQ/4BhixlD
EZ4/7FkzokrGfcR5uv/m9rMwUXeUAtcR/gJ1gSyJoFuSqP18gseE64uxBdxeOI3W
bq8VT4hcf+mjb82WRmzNEJTtlYSFNOXRATc0yrVhBdc6D28YVXybxfwq1gy72ARW
T4v544vc62JqnoWA/mrtLUp2fLphFFnKXpcuu8RYykOmr7o7Y3QprxnHAZYgAjz+
w2ngx7HjWkhW/P3s2lXHmDHQI8CUCCenTx88ZMyi1yROLVIRGG9omU4bsf2TC1ov
MrBtyUVqZkZCiFECRI3cV/GXjV5bGQm/SoZNQw93u2AMboSh7PvvzoB5DitpQCwY
HX8CVvqzvVtJrgjIh+a5XEep2yUwVoeS70YRes/qs88hDOH8jEeWLiQBYWhdE27Z
kmKP9T9AHXD4wqg7iYbvylt4o2Rwtf9W4cq6Kb/1i4GIT/2pf3jdNoYpINLhRtGm
a7mzufR0s1q5fpJsRJ/jKjL8TXMsrT0o7ortVxzbMHfREtrYaUGVjTbaf+aH7nEU
HjH/kPGKPfzbHxStwFhKOA0v40cTXt3IVberoyKdO5tCRtr0UloFYzagG85AiS2m
ibyxHsbRnkf+Zf9mOQ6/Sgx3oB7jhW1WlfUwlBrvA30wxqhfBTNU+0QCPaOVu/WS
Fo943+dTAdrfzZ06uWx+5gnW+ykDhB4JhOAIwKCQ5/MTVlP1q2uCQ7yFojSmqRvV
ev9XBprgBQhcZh3WGjR+ls8a8Xw/WcvmOPaBoZbwFVjHZh2OxPTmYsivxE8jrjo+
R1VcL39E1v1xubt0tyLeT4F4iWXURcVtulSe9qWS3vxC96xPJvjINPieLT0FoJg2
Br8GgIfPIwEYM9ZhFtNNeSOAy1Hp9UCWyjDf/CinMB4b5m/7X83QYFFipKTOwJVk
Lg3hhdgOauNxNWxR9bPdtENuZz2BNm9sx8L1c4K6wC0isOYDrAWA0tlAYpzOM0/m
+XWnaXxzi0BcGMMlWiVY0WEX8moGlzw80kjQmxTy9x9Nm2y77dqWjslAJTqr3P50
l5VK3t6luedQSRPn9uXg7sDuWwaUuhodRqp7VSiG0SksRNJrCSNoZEzjhqf/ZQFG
Ofms6F+CEU4jz7vMkFMKa/CDfZurqdbfmucfvIXKYvNoZz7ud32XYcb16gDx1k13
91nva1JifaeYihNCPobSJ7ODNB6Z/u1yA2eUIDe4zpVwOmpixgLahXX/f4gVc2aI
8A8g7+aZ6smfSV8BOZyFHGqp3F6TaCBiYVqVmwj35tssGZGGxHlQ2AEErPhVtqvR
9a0JaLEiNKODzTBnWiNyklHgrdzMLa8FiHnFpszqb9xNDMF1++WRgy0kRM1oaq55
XUfPQAfzd6N+HI/hosP7FAvBxhLDX2v2Dyueya1CKGZGxGPmTaD22kASDn4Deuq6
8DTv7GHABqsBg35a3kDpSGKtAXQz2gm1lyzgsXRh1TV+nUEmz+Mr7ROdI/ZLx8t5
zGtTa0foojQDL3Pamm8+EDHw1tLLwY9lMgY4rNQyYwaJk5ogauwpPit5eo+0yuIv
3tji9bz5u3LNm/JaFlTUUW2V6tkga/lUUXUpy9oOHGJ4weVAt11UJ9JNKnnMMBv3
NKSFNZv/oMmJ3dNXVz7PKv8TvtEpnlzEEZA5tzzYnmz09vrKBjOXiqumHmvh9tzp
eoHKoKVrW7PgptLnutzol8VEqfZxIo901feZg8QbL905FxVYOlGAJM12ATxaoIDM
1H7wobXQrVnUYG9rCTB8PDjCZhm1QmbrzugNlYyBzuk57Hr5N/DMjoT2RbtCTP9H
Wv0C3VjPsdg5m/H0wPbWUrCn/CQxeO3eAA7OepIudg2vGmQLfbJMANRWaZ+ASMPw
X/LdKZYYyECzvieDCO2qyYLVDk/XGXs7MuRacHBoOL9DaEH5zP8u+BQEL0dCnuue
fc/Raa1tebRCvY3R4AgcTrt9NPt+Yd3KHlluc89ovqkkgmFRQ12vymzp4AvV70Ci
6allvX6vNX4y9vAkWuelfDHTUm6Fapn/W4iUoVtGxYcSAuV350lFVF+zPXA/zER1
Nx1vp3NBAr78Oc3WKcumu3ieJjN8ixDPuFTSrKDBzgtBxSNTtSA4X/d/mK8BGFsk
pflOyJG0T/G6brhOSejwoojz/J2y9+a622Bqj5q/KiIy/V6iVrrbkoBeR1t2xXTo
OcU2hG9H4wUUp5mg4K1qMch9tKSfyEVxsVN8y6c4ltsTU4WEYVmBxLh5o0CVnusY
ZCv7xNH33nBSWTnlmUbkLcOLUkDuW3sh8EwkoRRwu4okCcPG5lx7p4KEvYV9Dbl6
cByB/ghDIUSE5fqx0A79t9xsVSoE6Ibh5QfIiEPIMgDkTHOR3F0F6L+ChxtkWnrx
QWWxSS7JI6JPOJ+6H//6EJs+9rQCw3Uk6L33/zWzngVwpI2UJitmw/rG2nWV0R4e
1D4Ulvb896VQnY6ggqs6psRJgAYWgqWmtER2OpS+/BQEqsZQ6P09qzpwZSj2EOvn
WYtWK9TcwzUuHZJTRoZAK9/Rz6k3sOSkLq4yz3gNiTyS6o+4sX4Mp2qas9xM/EPM
ynJ37xUqM/pJcNK+plyYTLiXDpIGPxrleewBEYabP1GCARV79rCHze3Pv89fbDAU
gPExJD37gvpAGYIgoQ1XfvrmN+lQpL1h/7aPhMSxZKhgzbNeoPG0OxfHGQwp3i+F
nIZw4T9UBS9Y2IxixjezNFpTXtIIikoY53KWdjtQ6lHVNdtRzC1Jbq8owqHuvhHz
x3Ic1GnPcVHNi/H7glDNYFaNhBx4ORBWdr2EvC2a5y1u5Uhget8J1EK8uuOe4kcj
Y2tNUagurH4Wi3ryTKsqmYdZzbkOXtTqyElg4WniiD/ZJ4EjqUgS+7FLOxUm8AYg
L98QWaFYuLuVGziOSMJha00OsThzfJ95ZbPfA6bHESP6oDuWtYkmR66WwhPCUIKw
gmprhhG7g5wpivGfiEOwl3sMZ+C3n8n6nQNgeV5uz6MKRNLuMG412g1ncZW1DijX
6jCDTEgc6CmyHAK95osSCVFL/X5pPwG9uMpt/qjByWfn1nmNmrSlIfvkn1adtBPA
e2Hau90uCvCjilqIyOxG0gkQNryC5wqXqwdbfjoHNzn0lhq9d5pmahX3q0yQSdo1
mUZMZxKnlYmQy/lzBVKKbgnLAPsKeqmvlqcWlYgRE13djgDwsPIIeeqGolQTN12R
NH3PkgzPgV5UqNgYMXDLlLOw9VQXHI9vfAA6H1dfwpR7/NblLcwfLhBYEDKrCBiI
NMqe1RzRYiMcqHW7ZaQ+2hBZ9z8DG2mqnhVt6rRJM1Q5SqaSo+qreU6TQmhL7atO
K2gZsFBP6sHN4XgaPLqEEy6DD+dGtG7S3+AIx05qfCS6W0QoqS78rKeecBdhrboe
IPkPzgx+/ncu3Ua6B4YSExX8Bd7f1oy1osWgTQhOHe0ToaZdjhMzxJv7X90g5rsB
122SOtjHC3676p0Csn+W1ZBx8Vn3/EwDAobt7hOlR/kYhmmLRp0+590Aq/j0lZ5/
6B14Q8Sp3xMQUfWW2BdVHqLfEU8exzOEhkZ23ksIQH5JnGgYHMAt++PVOZ8ZSYfp
9BxmBWn93ssVb8mXX/HL6M+lX9ijGIJHHBw35wpuEPy8x+jKsbKIG0I2JIhLxs5A
Dnl2wB5QuflhX3LYZBgh+MmrhdRWPnyizETIbVere5CjN1Sf8ke9BbC7GuZ7CNp4
lnaUBhKKV0M0v1zdb9Xo0M/UKGU9N5JirUTiNPJ9cSH243OwXhxoU/CUsts+pnIh
i1pykPg/K/H4BWtko2Uby0gvJmRYZljrLHYS6W3/+THIxyHXCUWmw1YchYBXH0PE
au1m1/M1qxrUXvN2pDfYVREIZuQNZaQEKCy/SioD0YruJ26Yj2NLIu+OrROI6BAU
0LSnhKUGs3r22bx4GqG5M5M//VYMFx6mpkVoqK8KsW2tMSWNTVQvsV2or3l7UVD4
qSdNh7CIFlD6tFwIpgQ8DJdJNEb7w0uFzIbEGHbZdkTWJUU5Y9TXDcpF3fCNcO6V
fL80ltciJU4K55fcLHjtDofnYjp7y+qaE5dzY8FZ2Na9CkQU4mMAkFr/veEwCZi6
jMKBRYf+LF7uW9Nuh0/mPuivQlPeq3v/CsFfTRR90XBvncTy0vc/HLq4HIoklHNR
oQFgGEDQ/VD6jz+Sj6JXK+vtSzKk+Ic6dO48bZepMuj0tpXlEH/hfpE5K24ALLf6
CF4wkQIyyrAm5TIm/0qxnY1kXGyRYYj60bKw6zg8KOouPAHaZ704FGdyT2aPsqKV
Bqncprqcffflv/JR39ly5LGIR13bkvEgaV8IwyhGjnv3J/Teqf4rZkW+1zpv1XxC
J/skOWd7gzC83XdjGiiiJJlHp9Zgxj9BBsv3bWJ7PNWreQ8EiXQKD2JPzCU3f3HX
Qj5fwFBlVP2qE0lSBVPhkjV/hZEThI4Ej5ftgPlQ0RvAXTGPtc/O9lUBmStnY415
fAOiFVnJMmRjd77QEFTwWdklslSXlk9RCyHK9v6CDSdu8IU7yPeyNMmJ7OvzLbfS
lPJ7IVAd0pkX3MupZNXy0/+s2unWz2Rmy0nDIjH7W8K54l86OBv4RAcAjw5x0gbo
Xx/r6vRIxI6AoNmTBjjcbH2nOOEoSFg3lp0P1mVGf23bHIUlNh+tMx5jlGduyDzN
Qht1XZUsQoXDDxZtsO7FgmFZvwJJRbtCpDbPgcb73D4wYN++0i5kbpYgTYwos3y7
H7C2XVbXIa1/2guUcT9p73Khy2MUrKfc4cteF5mwtZKuQ98hrUH12nM2OMc0qJyM
Mf2ntfd/JwJGA0plgqk+u3F2r2QahnkObBbF0g16VqhzPUnDZwrPzYpybPz510+8
iUFSxfOZ2PgZYA4itnKjLbexE/DmpXce/TZKgnpQPhL4BII1gYVNffpoIC02Mq2K
KS+hvZxWS/IQlZFVDNRWpQRbDPpf3VQTiQfLUVQm2rk0TnFd99zechv4AXX5MQeV
zZBhFcsl8UI6CO9hvkqvujX3SCeyNPshaDFc2PlOdSWs5aVHDXQVlECQ4CKEFlsC
ULoZO++6JLdg3tqR4GVi+C1PqzZiU424btpiAAQG+9O75/n86hw418EudrTreQB4
ZDNn9DbSIqmN9R086LWgkX1BRvMDKq+SrZJrmLYg4grfhAAPtrzg7m/JoDhBEn5z
mUrILPOUdsGgnpcvguF2iqtYS0b8CvCwAFo4n7E/lW+kR8S8xxphC9GtyLCAw2Iv
Ui5btbdBzghXn5VLSdA5CZ8CRlpcpFzcAwBQFh9OVIqgNeDprVe5eGkRwSCas2ui
b8JerOOGc+44XcBko+qWtbWfB7zA2MreDvJgLonyS9JJd7Fze0FLcb+WtBZ4L/Cs
0mmOVR8STpPAazerzKVfxcv8oQGMJLsH33Qz0A+09ribllZP0HR3UnT0eixh2ftB
vEfnA/lpl9W/qWzeSpG2zhuPRjvA7gajthqYaMScdUrMF38XvAr91+Q7hS4RSwJ+
yJecq1iW6PYn1TNeRmfetX+fThAIiG4YbfXS9U0kyZdKAp005iPCFUqyBeIRH79g
tV3WlCEJi3SulZylxxgEAOcnCBuWEiG2oj+ue2ATjgYwUTTOvX5yWHfc+8q2jpUT
Dd/TNdTLp1vE6mHBWCDz1zCFpa/3o+LF2jpNiw8m6tchYG0cvJSthyYxpt7O4o8C
6ZILDj3assIDrsqnSzrlMv/XpFyWErw0EsbtVD+ClHKT3lHAQLKKW9AIFfXzlDLw
VEubvNUXGuXF6V9QDZLhhugrPmvpz8LPw6AA0lJebHtXiy0cMOBttVMhTMdrimxs
9/ZNDNtmZ4iQ8G68x/C1nMvIB8lNsjHcSnJlIcVB5VBJYtNksMalPhOnzmmbczOF
gGTj9PqqJx7nNpvcdbswthUQc2c/QCzZk8QgoVF0F5xApa0PDjJgP7O7ew9/hnMy
WUgTlha/GGkIbozwyt+KrGYmwRcr5Z2V2UKgI2ZPQ8T/Z7A9AQHoiNLpV+w4exhw
XI2MRziK2Ccix0I3BmszbPcJEAmTvMlBO6HVpNkc5/rs2N4ZKlxJ5CZYaKnXMftq
OhWrUqjiDL5EcX41Oz45r3HPxidmfvGD7Y2eamGqRnHDxGhH1kGnmbZRsh37uhWI
ORhp2m/VXn3XdYUOOLyPwGv6XgCqUS6NcChNdp5/+gv5hIqgnodRKKwGpO5GxgCF
mNBAKYPxl3+4suI/UHX5OU0rW8yFmUZPNxOhelQEWuQEtVGCN9kg2K2yGj0Zqt7N
O8BBRkvV1G9Uz3hJqwixuFUs2vgDkdCT++WyYSdy8l0zjE4AHpBlCsaDlXN0K6aF
MB35YkK0Ei+dPW5PaUzXY6iS1CEsUplrt0bIBqkpWM/vkaYqVqnvsy3/T7HfRl9m
20a9Pav5hUyM15Zv3qVqsHV09KPLIePvNMZ/bGzlkzO9RcBAqUJQ5Rf9o/y1wE94
rCUunoT7cB+dIw3WwNBahmCLILk9700AwTSX2KdzxTS8L2BKwVJ55LWpcuBXhf33
MeP6GAJhXiOiM4Oa3G0pXzG1+4OfxeE/zovScVOXv40zrSILQhXtn+VTJI/7WRD0
Hjrhz1cZLpI1fkNvyziETzPhClYG32fo1yuJYoP7kQvIPn7vjT2X81oMaO2Hc8J3
RoEot4sI+9hNoBNvsCmRRC/i3TEkmeKF8epo9tyI6N4bGWHi3G2bXbbepRY9RLAN
Y28OwVlGdxxHgxmgsH8qlSPsbk4uWiB4LBVrT24JymaoesVu/RB4vnUO6IfpzLWf
yaODonyx51f5llj3PmiTjbwHzZfpTPK9vD1QPXkw6A7VzoVVTL6XrOOXN5Tgfm4y
LXZif6o9mhBi32goXvG24HIK9D7yCmFoDaCkN5gEOWzwaVbawkrbOcJ5onnaElQa
LXT0MXtVby9eTIZbdSj3JE56v4HVGKgNO0muLIfw2pLGeBOuxEHd7hNFGhysuO7f
7ShLl4KojfPtEoPyQsPjuJhbb20M+Fa4NEdAI8iAoslT6Bg3Ws9rbquRS2Og7Lsl
rA2YnC2HxaLZg8F3PnsAU9TwIttxk7Zfani1Zz3evp2dzGxzIPB5cS9y6Xb7aytY
6LjNJt/E0KP8Nd4w1IQGzb22nFkS9xD7BmGbhigz9AJ4Bt4c/cKqTFRNJWx2rLpd
8Q5B376m4Uq3+c3YZFxSEYj1g+GgypO5YiqXcdt9P/OH6FEdctudv7bKaptX3APC
telwp2zm1Mz2Z5QAHx2LkeVOM8XvqEfg9kTUtuCGyv8jY5oS3gGufYmPJ+sp+gIc
Jv6HZlIyNJgwcFKJ8Off6Bfw2ZRDUQ5kUJWXUFW2xhLSHhFqvA9PlZ/4daSwHhRt
hKndkeUVoZkcppC4wati5fp2CEqNiRQpzrT0fOxfQ69zHyBfgebVbYD/mcObn1Ml
CSPAHQe7xJRkc8leyfKg2wNXfAuZvWYZ3LvpXaG2qSjn/V9Ehf3Kn+0y6o3VX1Hf
a5iNmVMfpydDBFJH6h6oCnwxypitVgt9QLLOBKb2YoMdJhKNnbrZM60gv039E6kG
kyA2umeBbBiq3rBjSgo4PkkmRSk0cZmp3IjzEECGLUbtGeiTrjCaaXFujqDh+2ug
TnnwhO5XdVyDxKD3p/jXRla+kMAa6cJgqL55DVFPRcHyYf+yuwylK/zVetc9GiwV
Ym8NwMXu2PYewRRA5EuGFdZJdz4uqC1ea+zbAXhlgcOJ7nZohWKdUqD9STg/1zhW
205m3D4QR3l9dMAqgUpLXgGrf20ylXzRkzjhCqvQWBvqf69eljw7YdIiUOMYGcEB
Y2X+fIgM3GD3Zu3PQEGcx8irGWz+cN3mzu35JJ3dj8rG2dv9axUTFqeApHRw9mBE
MaoPZfrHQFyD/WfCmNYwDCxJOgcYXVF8Mk+cDKTGpU9jKdNnPZOKWglnNo0xPIsv
hLgvb/dH+EQ+jM74MvLutmnT8lkvXC7t9+bNBlQxNe++IFKUDGp3+vZmmuPqoTKo
sg8g47sGI7lI/8X6Q7gc2NL1b4GpQwnuaC2Lck85/MZTIxyp8la64we1XK+G4IoF
b+xm7iOAly4Ot5W51tTcgicj0OVklZY43qTE27IMMGR4eptxWMUU5D8V+jTNzHiS
L3EkrKY9IY2hy8eGme0lZgGEFkhNAO1elANEy+AaCHl/szO2A67GNx2BeHsSjg1k
I8syeUR1qh7GksfpXFl6n5SFAZGY0R7a3gfLbY7EXmTtcvwYrn9uDhkfMqfSKjDT
s28mp4gRCoUOQQojwFwPD4kaKngHVAa12ojVuxdNy0jMGtDc1Ft1DlZw+3chNdjP
foDcjbWMBK/1DYtmbz8ua8NtOY71itloGmf98H7NjC2rkBr/VyWhGFJsXicV/h1R
Dw2AD5exb8wnX6k5aLhiY7CiVEl5peYzHU6fkdsWIE6SM1w5kd+JK37NUjAK/R62
yhzIgJDOKze3rjdtrIY2QHPPfJnM7PpIn0EAMKae+fgCANpaKWX/njHqiZIBJzKA
LxQYD+f7UslS6mT5iYAOKq+2oIjzsIpsodeM+SZL0NMUpR4l7D3aW5FJKk57SIT9
iIinUYOWsY13lPTDipxOPVfFwPJom50uteNAXf13YdXozV6T+5l1i2hk/KDJ+yz7
VLJeJ2VCFaw9KQBF6d8oq6Z6ffVjiyCR8SiMURpsJLy6gmd9bhqjR6qz3AM0mPbv
2I5HFgqJUHa+eSbLAuH9PMi1EUpPhTuDTcBKPUW1v1Xcd6r+9gRfm9OHY5trulsk
kyWD6GqVxjcVgY5CfAw5qVlRR+E0TnNvcSvt0RUBX8xC0tVA+UwkL6S5WScAPs6D
klQBi8+2w4S4quEqJaKMO1pncvORnuGmEdN4YI1BgL4f0/w+69bDH7mjXJBVeK13
j8dH52cbGQc7fLPo5CsF5BUi7h4PpFHp1FQzbVtXHGin1oNoJrhCzxY7LXQlcH/i
AXlCUIbIsHJ8yXIfn5KP//ZXcGxfubSyo8sfGvQ5CZE2VIsqKi9u/8FUCxTacZme
WNujTihs6rXrJmirOM1Dl/Tv4Zf7vRkQD8IKdZ2rBM6+7uTkYaJHRFZl4iV0qUjh
HVBFLkmk+KXPuCU9QOCIIKI4IAwBJ+dil/mjlr8E7sRnRZddvAyfNhxUyZg1coYZ
owFERYGd9QdN2zaLgcz6nsDC0nKOI/LxywJwtk4sHe7RlX0Cvi01IYgtIuCWarMD
Vqf1cv4eB0Pr7b1uHK/gX+Y8stMZmo7jCvKW1p8jJIx+4PziV0dJp+LW9IfEklTE
5roff01TVgS0G8T0QGo5h8GRea+HUzNcBLeMnAvl6bXdUd7jBRkmg+ge/7ZsPjIZ
XK7FDssgu0FzPiA7X3BccvDzGUogShVvGGqD8K9d36BP+qeaginH08a70Dhn77cR
vDTccUlLKdWQrKCc4FwHPle459MGXOJaWQ6vbwbzi2CPePBqcN5JYvjN8te+kGyq
4PadbCeQiUYD9DquoZoLbwzFOXCJ+9b1zdo6G7YBmCQI2cIvrOMyWErmGVFrQ68q
3lfJJ8OEvCdZleY3+Ob+oipXdaq6PynB8V0v30/sCSkFBCWLTQDaoWzA2McXK6+p
VAuc+p5aQxungo0Qa/Frz3k5CTI6pfSMEnCwAaAfAg+CAhoFXU3wcO0uU2eH9+Pu
V1OpA1d/4R001jIuUn1RVOVkIrNhbVs1FaMHgD90yq9G6T+TN5MzaPYZZCPHrnTa
SaQ2VMV+xKyOAl3pryRREta6jaqTcjnDKvExlbJPc/fdOFz/TwddSu508jeXDQJm
jhp+tJbxV5BAOtTr7lgq0CtHY6WwGh4E0uj/A0w0DCFJ9X4zel92kslHXq1jAPaX
6TrVXHHj1lWHUWT8T2uOyWUkONR5Ho0Z6f43MMFpiiuJ3dEysB6r+7kQvYYiuPXE
bp5DKnowm9TWOVpSM2QElerrDi+8UE7Rb/VFZDwGoJ4zcsnj4FfmH3km3ETmvx1V
4iVFCp7i70UUTG6ms0igilxJhh99IbR1bYBaEhY3hWU7HPJGN4Pil2eqiNhnt2UO
kZJ3pBOtVcg5ymD49IPIq0jHcqG5O1BTkEK1Eu8KVtB4vcN+nE6FLB+w3smwhIjI
I9fFaQ0crtFnd7/L1SyZcGD64RPSUch/KTz5zMSc1rQe+kuZPqC620DBrHXGFuOS
ob4ZSjFraydbEpiQHIO1Cf9yWvT7fjyMmzes2bTH2cOKrSAAPg7wPd8nwF8LligY
dxYQs+CM1nh+7w0XJUbqttUzGluG35GRuZTqj62MTJy6NR4sgL0a+DPT4JcbnhJ2
z9vVI7sDAr2J0pROOKkkgNIx86spwsCBxc+1WbtDPH9inZ4fDcwRmMH1rO4Arsd+
xhSnYy+eLBvTnZG7nwwJWJ2xhX/t5Nht7jPuzmqM8Zsze2OfNYWZOrEvNyHXsd4g
JrmqY4LaQb17CpZeXSCC7MqmB+Oq/rrRqxEKMJwJ/F21pYhVoWiSq3vZ6Y6Ujq04
C5TYvMBc/UCsi4ex9D6z3x89Sw6a42pLPKlCO+MABXYozSA67+VUUOjB5sPRhLsC
58i2ilh1dd87gXZpWzz22bxddFmO8dd2YDWYeLEc+MCHe9xcoPDXG2GHn9mJlTQ6
5in++lWGeGV9+yxSVUTSM2CtU6jjzH1V+B8KxL4psxWWDKS1Q++yB/EOeVgRExqG
WYL6EyXUQYbtuQuxzYMmIe1HxVfhUFk523/SJE5M4Kuqp3yfJJiL0tJ7YDE06xbq
RepCuqmdWx8qxZGiVFsQomX1vkNzAsqPgi4nLq+204kTXWkkWCXac4EJBncaGjE4
lGuLg3VUYnHe13whiBgAz5qyvR27VDNCs4EIMS/syZGAZmaUowfWnZVRJihYdxbl
gLpkGoaIQFPHUrcN2q5L2EJ97LzxaVdUq10LPH7DrwMHu69Nmo3UCFq2BhlXLaBH
t8lRmJADHmzy8TV9+N3SA7T9AFvq9MlGaxxUJNqgXaFKAAaIG961oc5MIJ5+aCeC
iw/FYNBqJrK0cQLPes39PHAxggaHz2rpk35XVWbpqlyw63WwJBhXbZSeJ/2MDBxf
Eg9nHtXMioGpJ9CSDNJs1UDS/rf9knPX0j7/U45aMiw8EXKZoK5YZ86oaElimjz+
R561jbUOqbpIUtWrPFPje3qjK8dkyvk/YfGOSi22cZs6ULFTTdQcvglpGuK4I5h8
dtwpHTGhW6IYQKlZNl4C7yZNl9QlqKLAWeAeOT015vGrn4PePkmVWg00TYgaTQ2/
sZJZrgBJUpbHIDpuljx6vJ3AHiiOhj85q6O9PmF5IZuDNdtAmZ7+rjpKIbje7cj4
+z/j6pVTaxil+F6q8DOD+B9qMZBlPuo97XKLqO7EkJmLRNu2+32nX+7q6XhXtXGq
XGIcYyxnC/PhqwP3+GOY9KlxBS0tkKqiVGkWAUwsWHjoo9B5j20St6gx4ZgNGHGF
/LgzNa0DSeLBaz59FvY6z2Tg5gTprz621kazyazWeQeq6sBLSi36dHc6Z5ROB+OI
3m/PriY+2vBCeE2ibCNw2KkyMZ5sVfwGRuWp59KdKL3CE0XmrKqsiL64iIAOlCMV
inZTfU+1bQivcGUkDK87GH4tFivXLuI96O1dq9WKDD9uq3E338mulDKUS0zt55TM
zvKn5HUhYP+yw6+DErzHq+tJFXu27NBjreRguzd+TbKIHw/nTD5gZSA/udKrK9gW
P7H/MMxsWi0AKsKk3Fwn+LjHz/48L78eRwj22KhWTa8LHAo8xLP0Q8wpMcIt57nT
Ah8g0a49FOGNxsS8KmekzAWuhKdXWB+vCVSQxzEGHOnNkGjZg9SISU70XFw/OIdu
peIIMmPyPBJm7bNn3OcR311qxK6CXYjB7UPu7cK/Q3tz9aKm1P2LiVXngMbQM//c
lZVqdOUylzk8W1WNVtxWPaXyCY1NS3knzdoG9j6EU3IoIytz1cjrMXfn6T5ZHrN5
acKPlcSyGeGWFNkmxiCwb8jX35/CjBSFz2nqi75wOrOr3pNk931Mmq5Qm/ztB5Tk
VKq13DH7ihW9WBJMb8S6U1BVoG30tb7w44t9DwwLXc3hMmm1Hz4D7RO6zCIXgvQC
Kq/0S3WO9xZaTAAjC3dv0k4QPIDPZn3ARHRz474wI1uI069I6mvLrQoCQGHGLSyu
vu+KIlIHskOQ2Y3QPcVHYOBuwRNAU8qsoc28gfJ1TD4uCqwknInJahnM4W7wd6JV
PEJyhlIjaqU/zN0nrnSw3VA5sAfUO65jZCARYIJUCbwil8F06setysnlYF1TjQ3+
EKfLfshps3PEd0lFo1z2keA39/1VVrQMzIuiLuHFNoNepv4yqyMOLVluTSkL2KiF
BbPuYP7M3CyHstykKcx+/PCv2Udj47VdXqquQmFSOrZy4eG04RrR2LZloqP79M43
tT0o9XIk5XIF2q1uedpijnpxXzyOB/ljfgkdBfCmyHuN3kULQ0/WLYk/QfdbMfPN
Cegu/TpgAVgcWgKyN//1WinfMc4pBI5cmw9sJwAbqAIpvwRQb6kuZLw7GJ2Zyhk2
w4HiDPsgDI358Ivha1dl2cKQV/fXkNLzfp7XzdEbltpXTdJ2/3EaE8LJ4fKcFivV
kT2qPImDSEfiXNiTS/oqN2A6aWJNQStyFwLoU8iPO+m2LI96RNYT2R0SkDlFwoa+
TJp04v2vSt3XRU89Kwj1uKHpXpcjTM5vVquz7aeZQhXBe6RyQqvaDq9duVR1hRP7
86KU7Iekb9H3ZZYRKhvwttN6QIkQo3nh+vew0499/jplLnf+LwY0yG2HNGO7qMS2
h4EfMvM3kjKHEIuI75IRNUrhQa9oA/w7gnmfgxHgSA1wubfcVp+HgleKebAjtw/p
nzuW3Cl+9/dFOIkJ75B5MzaHYZAkLzxyw7vKuKYfsjBS6FIiPtftwlhlHOJAGpJZ
0H0S1xq31HWrskhJsHvYQkqAeRNArYGn+XpxLHYwwZZkZQsMfyBdeGQYGZfd/qAO
MgbQYQDIZ+GZiychLIyENULENUgLjACKekJvKKeHpqp+sszp0rxp/v6cjmPAy0hG
lEj234epcs0yp6NStTxQNGwYexnITUHsPNqxg6xNeqdrDWoPMPNX9+NdDOdcO4Qc
WpizYzgSXHNXvBrFcxZ2KyODReVc9X/KkOnOBaTj4yXGgZ4TsH9tQu0YM9C00CGt
mfaGP3u/Lg9KPemLa4mj74jxdE89u62j1PN/FG75pP/sw5CLDlVCAC1TaNoaw9RI
snU/uKMntJ4CcEPad++x02tnUA/5uk67YLHQMQxtMgNq27Yuoz63AvgQNXkk8EH+
WhqAcGuvRnz38PEt42xN77k8SM7Lj6kkHHykahmc/8QlY79XwaFnZeX2NVofMUAp
aXcXg1B9b5FrnjF8dCY6/dnVZfb8R9nv+jd0KDN8lSZxXAdCQa9JpvmUHEoYBYa+
YkQFnw+1MYfs0CFr+wPEtxLFJlIftxRcLblxnJOBtgG85ui3Ws8g+mkZ2i0vIRFW
rty4l6uabl4x89nYfj2CI30zb07LepcUYys6lT3z+5PqbP6SSTQ7+qTi8bYQKZUN
KEmRscaYtBWuKwXfSq/N+v92sx53THIp9BEwxC+pQZVI590Gcsv+BcTvM+gu6eVw
+t/veJg8Ejnhp8kGEcLRp4paNrM1kyYCBm4PMOoVZfUmaTouKFVHh1IjJSKv9r8T
J7PLF9XqAgyoVcW6yFAtNdHjnPrCtr/X0ppqW/TEzsK0unfkeKGFuup0S6GwGJjI
XhZJ+hvfonYOZgvjJyE1CdZaNT46PQg3NpOtcMmC48DTBsgsI6klEc9BfWHsCYMI
VXfT6FilYBjHwk31ROtacPA+M6b9/j9qsIe9Ow2cDko3W6gA5JXHXHF1avAbz2mD
WfSjavsnCM0vKk5/9kzzE0j1yOrd/cqSJ2/X00tD9MCdEKBjPwucEOg6ejG9wJS/
JfivfcJd6JMkdXXxHe/RHY2XPP556upx5iXd7mAKq/hjCwhXFVKPm/78NEzESYhh
Clufh1vzmT42BHnPOJLtq3vpO1C7/sPbicx4AGupAU/F1Hq6nIxoi5eWgmI0VNtv
SlBk45nOrsyVk7BlwxnhKry5aFu+cK8vsfEa0R45FWw5f2dLjogka1BZ0yX488wG
1EDIWxTDG4rKWBQQcQdBbSnfEmISjsd/ZXIZPpIqTuiCNwKGuVIGdsQnqIzIrgZG
y46bNuLPaRhVq3+0Xc+X1eID1vUY/Dc1Wn364pG+JvJfpV/HMgJOldNgqZNBW6AP
B2y6DbnCGSkbQfNhAVv+Rc2f6VttW2eiSbhW38DPgvu3LLt2WBEHeT6PGbRgmFvU
P/7T5MmA+R8MY9jXNDw33uh90Gk1NcKxHzydIzmb/1b1rESpZkECit9V9q+pSTk8
02AzuoNA8jBKX5rEMhRyCsdrw8DLsFNHNuz+t6/gu7QtdhOh0qdelZozOQcC2E/M
/FpfABk3+MmGVF8HQYM7pUYxmyZCEIs7zaxzis/nrCTkigVGKKYAImaYC04Y/yl1
LU5hb30C3M2ykYKi/ocgXbSMaazvmRqOhEA2EojfwgGzYEFo3CLTzxK8v5JgiTT6
pCl0xMiLPjRZAjSjL7SOd23bqVLKHas8E9V4N9zwaRoxUaCNd+D4fH6Di3PLViN9
fWc18DwqMfvrvxpC2vUOHCYKWwd1cw3yMScovqB6UqfBsaXHBB2ZfhUCkDeAZMEw
66qkL8xpAEEqcPU3pJP+miOlCUUKqbDBU/lT26AFNliXvXmRoZKLANeSyc9CEe4x
4IuTCUkCQwpBYWM4gFaWYzI+Rs9+kdjkJAoK0Bu/HxTVUD+xf8jaYcIvoFg1E0QV
Z+fMnQIDee5vd4xxBBrxnubc80+dDCw6A3HGLE5/u8i074Z1xn8PYhWBrruiyLVP
6pVRmFrxZXawfPBJIIbbp1tQ6ahzVEYrHAqRu9rIkqZOibWa4KQNgImAfBCGc4mo
Owp1TaJ9Rzv46zMvCqm2y9H2Mg7bkVihW1XqJIzfTeWjt4ZPchp4sjPGuQrMnDwF
Iv1TQ9Es2mJ8GxcXI3TmJQn1KAmdPZpTIEjbkH2xYP0bVvj2/+Pcu90V4s6ikUaJ
H/BYr8zgR0cOHN3NdNprCBXuyOVUas2ro3VLCoQr2uWsRCYTgAjDTZvoaEn5xSqE
apHs4DyGrtr45mnY/55W2VnHSA1BAdzbiFG10W5FUYNxfvUrtei0d72WNr+KhhBQ
vc1zRWhRMas+fgeq0bqE38elSrzexQwD+bRQ9ZK5aGkpOXfc0aZ9q3VpO/HkvQB/
Q+Bz9uHlSA73lpisCBwBtwDXbsmSYttegcUTG1GbcBUdSThL5K8uFGQia5Ta0WzI
durX2gMF6BjfowkEfsdtlziAA+kChtosRLFK11U1AW1ATugcRpQ8kuHFtROa03sc
ft3EWJixZAxhGyU1oIxskdZCZiEuENuK19w8RAxZKPhDWTSRmJlx4boBsz9mMLH6
F0wdGGzyTG6THsoxxQN6ev5ty3tX3pM5liFkxo909P4di+M/vkUYAIF66yC9Iku6
A3IskNOsD+IYh+wsjUC2E/mQc5rCNkayDR/kMDysYCkC7JKLrDpy8FrsZaZ5xesO
Y2LhleruLm3fiaSlAdcy3/hcYvMFKJKuWpswDXH57mzoRmm7Y8VDnii9VaVxUeNn
epU1RC9YoV8Q+y1YcJ9b5f7MLFmurnmGnhXix4UKOOXfNLpkBmWsAUts/8c90F0p
UAuTWyTLbuWkk5W6G7ydNRFOVf2/dxWGvIr+M/Yl8xX+xxsYpT6V2cN7TwMJG6Zl
GYNO9Of+mqfV2gP4VIUr0V9v44aDYJSYuUR4guidp6alzwXJ1YYQW2muAdHngVjz
jL6lPx3EQF2Z9F88VVbcsZ5VSdcb3xXuDLx8AZAIoAizmfI0nPsL2yTUM3ltV3Rl
iCZWfgylEq25FmGP2U3SlW0V+FIBu/XzKajAqvM7h3cGj0VJP2d2vOlodQGnmR2n
gszuZ1N8KRxZoVamtMVjwV6W2J3hQ+/lQUMNCWzuEc1aZOWTJjA1gGKZ9RMcP5es
yofQM4ksxBs/akZYyLy2cZn/4Nj8zrwP5jGR/Ssae5Yc0/zqIc43Fgr86dvkt0Dj
N765emqQxH61/lijOgsOwn0/+N7ejvELKQnJs+4RKIFai7gSesD1V9itlH0Q1CqY
6RGymehRVQ5IrP62Tusxo8UDGkc3GNBs1klNJzYZVyEXSodHRnYvbAs55jcqJZp2
iydLEuDKGT5ZlZ8skQi0TT5k31IM8vV4aSnjDZzjN2HmMaKT/ndooTLwXrWn6JR8
6g/ntJb6sS8TeY8lAFrOeIlhh5jeR9SX4ST9mH6HG40SjGEJ7vy495kSmC7EyQDB
jVoxlZRNoPxzJQxt3+v2SqGriALc1dh5dlx9ThpCqsZvpqZsoy9W5aHPgXhDUVNV
4uwohlY2LLjc4tWWlsi04oZPzartB2qnvVNtcHSw5sVRc35RLYZAV+o9OOxiEXtg
zYdYrxP1Mog8nNwSlIQ4NT0wHVuue79yr+iXEtTtSvD4tJ08mAJgHJNVyGuXyhcK
7wYY5OeeM9BG/KXOT0jMQ1++2CyrPTN5RmDm0lr9G2hE1jL/Bf+ccsUr2C2ftJjR
VhSWNn1ynkRBVm9gfXIWN2dw6zYnCsTjHbTa8rlNKywhBARCgKQ0k4V/B6tSWouE
x8tj3PlumPF3GN6afzBLrKq13GKvHv06x7RrwNntmcm5Z+YScaGq4QEe1+xo6+Bd
DlGPdnH+yydD6ep2L+HyIa9KXfT+p9wOsIoCGv7QrdemLhuzkizlkdRGWyeiobIb
3xs47GYWfxIGTAISLssWivAHGul5WJsa5IBGR8H9UaGMArJDvuAw9oCqnoq+NeHj
uLzPYLxa+L6GCqT6Q3bYqZxPW0oSvAPVdLwIxrKGBlGSCwqMv7LVW8TDwW37ujjL
yE5txKL5yqmT5WrSIii2AVRdOFJ2ao/LChVrqGv2+8FJGysbbGUx06WDLkQv/Gc0
GT0uV0UMNymT02lpJ1MQ1R2G+ln0CNdvkNiGDOC5XLzJ0agSjX+ajsbdatZ8RW4a
oWwyEMh19fgV9L2oSatvWA1NoNUbneEeYmPklPQ8zQHd3zAkQiWAzKKgQmr1rByd
xWbSIRTTff8eDGhVrXRIYtCLYHI0W/RChtX77eeDugZWCZiBjHEqQZkloN5xJZNm
Nlffa6z36iJxPm2Fc2l0tlBA2SIZY0GYastaRqYXdrHHXcxOKuZStgjih1QdH6EQ
ZPKw0d0yyBz6si6M9O8RlUPxqHN3nIhlyXfVoZRS+HVYzbH1DIOOF3bgNYCnND+4
VJFrdEJbS0JgKjUgqN+i1aNY9EwDZthuCl5/+3oHwrAHMIEtJHLqI9peDFzWoWt0
SGsfd7Q8wX0G0vH9Rx7RNpIhzzbKirkYrD1tst0yYY0jH2b+MnvnBOvzDcIw852A
/2VqM60mxdxjt8SPcTDgFZkuyyqnMAO3XRFkW5Z99pSs01oXWHr0CmaTFY4ykyXK
FfTPM0JcIR3wv6p3qLkssybhsVRHa6veaq9iiSWJvXp6kRDSLXQ9Ydq3VzczkGRL
uy8/O3x+Rs0217cjiCzO/cjcC5KoJnM7GNB6zc2zO06G/1lzFJXO31lSktRHFR+P
k/MR3KKQknFnW0A7KJ80S7nQcn0DKj1x0ffGRAS7lodJHvdpqbbRocCD6XW1GkkK
unyohvI92iX8LOb2IVWoACbnElbqJDlhbPdDgCqUOkWsLhK2U6DJ3Xb0Kt8mNKBn
wA9KlaYS7hm/x5LjTGH/M5WKK475VVs165Zbw/G0NJ55V7SXJgQX2of3gtZnZA7u
a6rlnhYbFqYnzwY3iSC/VdBhbnYrA31KOo4ji0JvAlKaRhaFzVygmYG9s4/84kC7
VJzMnh5GjCAcyald0sjabqafJdNSN3qgJ/x8svkm2ZpIShdcN6slYR+rFP+j3qXK
BqYm9GhwY1awptRY798gVb5PdM08M2w7owSdYopND96y3x+DtPPH57jkteu5yS09
woN/Ex8iVRX9Ui3Nivyh0HuL1sMT5Mn6qcTFzKlMJtfJLYET0YFIJnEnCv0H805M
EGwfnX9MARdBAr6H1U++jfOx/HnqH4OCeSWJQm1tH148GV5jcdQv16KMv7rnUJ79
t3ateceQOoV+Ki5y25BfvQMokRddMIlHsP1cChzjz62Hb5qsU7HQSTfsVBmkE0xM
nXL5R4Nbj9EOpTLWSw8UfjUoa1joR0wgzKiLyYOlwNocdEbDiII0M9ioNBFO3K+P
ANjVn8LCpSHe1PJkB24Yt3J2UhBCUREJoGS9tp5bDZzYTrGGJHp7gh28ni6ab+Mr
2lDPyjdfZloQiRk7+FytX/2PdsKh3+AOHpPkfNpafPnOhRfdmh4ZXT+oEhNheviq
LG3RJVV7HXlNoIcfY3Okty8W96E4rPoqsnExenhLCb9PgbOxKSAM7UaueXcnRb10
U8L1DjMPnToAnYVzR31lJ5733oD6iGpcsGtgDFq88aEETV4cdbWs5mOP6zN1BGnu
GTVCA11lxbNFDyv5uAi6ArC8G1gWdvq0wFKZlyp6sPcDvgI15XySGUP9PY8+Z2i5
mACES11cQYvVo9ALs2F0qa9zzBXFLKPM0q8oH6m9dsHFYtm4htLJhV/kPaguZDhU
kJAAJ0U5kJwgymmEHRFe9THzxG5Jv1r8xwdyofFA2DPAx/hVcIft0h7hV+M2rGEU
myfYVvlgyMBvXRRoHbla6jg25CEicphLt4ah1ReIN9ffhHy1M+bTShJAVHzNCcrb
dhQd2oK4Zuw/BGU/6wB4lYo/1FHNF0CXmtu8R3lN1/1FghaGw6whDYilM70DEljw
RwmjwV0dRUqL+2pbxW624afwsG2jYQszwUmpv090sFkU3jwyONk07mC0MSFXDKBC
1Gr1rBAi419IY8dlUNFne3OvClw9R0IFfDWPBs0kO5GJDTTX1Il+NZ2UnSgjJtup
H9n0EX2SwlADBVHUno8e/5Krd1fGyub8pFiPp/LI8LtZBRf/QJ941ojNHM11TlOv
7pleTMPQywfy+3w2X9rVZkV40dyssW0WM/jmnvPuTCyalU3a1E++mXy27v0qhOSL
hatvLl+/LloZNFthXpa+BqT7oPIDVwQUXLUBcpJifvGdTH23N4wSmoe3pbXotVZv
4vOtik3f1XiJOfZi3PplbrznPERN9PSo18lTRYt7BydIo4/+oRpdua77nXXa+ml2
5dWtAfCWcaOHIt8gkJpMhAqC5HZ/u4oa0WFQkz7MEPua4OjiNh/2uNe7yWW2By5A
14YxSRUhU7XcM37hMQl4rmmbuLRGvJnwG2I/aCcDAv9iHSJ0tTAH/RgKrACgtgs9
nOrn1nV98fg9GKQNDIKAdTrBHpETvl6Trg8FyBB4Y8uSio2/sD0h3hoGmOes04IG
tanqSGLqozeG3f3ro7h9FU1tfcTmGZWci1zABfyVY4MMxXS56G0x6jtEwPxKJBTy
PRnK9VSRG7my2vptBi00M1cKFX3WpHpsCpYveUR4CotKNxssGYGxYtlLBrc8e9lp
/q3EGP42SPf3L5P8vBsnqpaIgpOkGcfLFKjMyfa6IxclJJ7Z5sSi2c+33PnpbN20
Wo13B4tXzbaRIIvXE4y88jXRMeR6GJMOvvmvjt3PYmy7W2VaEhP1YUlBCIv6I1Qm
tXLZh94Gx8p9dUB+s50zdxfq97UEfnTqkEkYoIHbzRqD+Pz+HShCFL/28bFStc1y
HLvUH2fR9NdbfsIgKm6utZCcNp4Du6IdZI+LHkPDzq8AHiB2f1mZJcXKuiDLiTf5
u53sEofJCADkNy29ORMn4S0MGZr70UXkR1xliJlaawZyQ38LZTxMaEYdodX6KMcU
rtk66PRY9yGl1Pq0Ns5b9VsoNpBGxoVd8C3euJnkJ/elXhf/6M1Aa8ObOh3k8IFD
nFhoLC11CxumIIG1Z3QB3YO8X5obGHV27Pl4om/ZkNxEmVyA66i9Shb8Lavxax/h
iAVVYys94yXRgj/vQ6zE7t3IMj6h1k/VT4VhPDwAnk15vQX7hcZLUyyOi+m64MKj
RNxmwzgjwyw8OXD1MdYplZ5AFd9aHQ2KYqcJROJUGw2L2yLnIJWu5nkQzIzFjbIj
vKtruyzsTEY3sxH8GOhoIX4XfEUg61018t3d3u5UwHyT56ZW6Kmik+NyDP0RTdL5
Uy9+LVF4MI1dUXMlxubxHv7JiZUKVUak78IPXPi/1qDYH5o3AsVq3YA918BHgJIC
261pQuOq0G1dqo9MzbC3+orSOXqnxoQTvJUcCX/rtFm5eJT8n55x1srN4AzTbaNy
VoBWhVvGqRZYwy+WW31YZdjGhl28aViAAZtra1H0sCdU6pJve04vdWZ/I6dG5N8J
4Je0k3dMnIAoVSi0Uux2UBsIZaUdtTbVZOcz294YbaSeXPDcA5ZHbS7CJ/m4M/MK
fJ3nzWwj+sb+F6LIl6hRiXLfg9DvIcUVPB8IxIgYwEB2Mlz/rybocaJLrwAkTliR
kjPaTwEopuoseswh5iODoHNDReUvHWSrMnf3fKY9i2Kx9uqh2vYm9QBQJS7MRs1W
pseHZXqhsYh+dQqy+QFLCBGxK0yn1OkhJkVnHSWURHoVpR2zVrBKctBhePWTkpDV
m8xFGDbBsHhM+d9jdoNnpXfz5tzwDTHh5QNsCwgPoq73a1ABLhzajvVb4otH2Y7E
vI0QrxH71ratpcNP/12iMyUCgY2/X7vyOev427AY/pwwVbfMD40lfH88hlLKTjNS
K3sIsrPGy8PEpuw3HG9yw3Jw3homSaj9idgnlK9TBgeaIaPUp58TBZfA2qy3dVT+
IXA2X+3xbuOQnNwvTCaO1YSfGD8vZtIjSY/Pv2I1Ap6P0o8guN0r6BI7KnQd9BH6
9wbdiirO7VJqIbBj0qreTCxP7c+1Ridz4Z+rFPua7MCDXx3/yEhpr7eXxslg67Zo
3i1sQaI30Di+dvthksE2lLRjSuLH8+0rNNn8zH6DXyCXSE9kQ8i3BbhqPJMKgphI
IojbVFGxcjW9cRsjf29Dznq4SWLwuY07ZU68GgqEoaob4Xexf4KvARn1lL7n+eWU
sTr64wMC+BS6IqHzLIou3xgzhVWZzoOXtpHCDAq8ulCdT6bDG8b5fjB9ANu4KghN
9Dl4l/PdMKZ1v0UeIWkHlCVKPhjcM23YQ0TA2S61RnrVqVHFwbmiws0nVNuX8m/k
SglZ5VhMWb/qHXyzLJvcWf3ZcwP3Jo0RQa1hqW5ktZOh1KlkIT3S9LDTyDCsbUmd
8Pf6gmOdx5cd7beqNPbPT2XJEDTtmg3Dv7xX2OjklOcJriO1cPdmWAgxCP+QqiGL
2mojL1TdgdnoPWGslDlWHUTaGXSAu+j06RegYb5Cq9mUiI3eiFaKOweCI4WywfKs
HL+iMF1a9u6C9J1WJpE1C43aeU5iazEu/wU5YL5FTBHU/xRoSbKEA31LG0+7L0Ed
yaL9/6HINhOPM4HRk4jnxSCo8i4kLvQpJ1wusMpMBVBWA8w7DHtzycJ30eu5ff3c
XyopzuedG4KYR1VvOGZY26no3rQgtihmyrQfWV/HnGZUn8W3PS3rNk9i5VqFc297
m0+0S2ieA88r88UC/3aI24//zBpRcUO+kiqkwJ++6xZOWo+mjn/SNDLg3PfdoQHU
AVwCYFNo+PnMmV2R+nVtfxJTQ0Gozq6JQKncED+S1aZO/m4nyt5WWuJEKP7/Iliq
t/c4ADGa7shdnk5PXHzWsBD/zK5a2N/z4t/SAiruYB/t3/s1MrU0WFzPwmzySQrs
bzrMz+GKRzKTZdEfwGH1+9vba/WVzyCoBNhX1G1GLhg++NyTQXA4klZI678FARZ+
uS6LLiuxyfr1k0ygS8F0OM8oTkPF7gqijrCtbujqzt5cv/Kh7ctayBuRc0nSBEDF
wobi4PLBCtHQSFUWg5eI61eaLkZLF+aV33jncfN3V/vCuxwOyo8I3NQXTK+Ef5Qq
qGSs2Os6clI1KF+1+snU6X8lbieaHJBoiq02/EC4XzeSJ/5TokyhYe2UR+QG/iQB
blV6999ov+lhbyo9Vw/Er8DycqNWBj82TByhtm+eyxtC2uOPSZnCGiUe5gHXUMoP
dx5oriouHnizTeOVZaRnVqweVhSzuhQS9pmw4pYg9pQ/KzzczEQyOYZo+wA7YMNC
1wAk+iMvr8tz8haOPhu4hguhxnS7tkXZQdg9+aw8rPQRJwcd0RDOqOY1MK8Ggi7G
JcrzkuISDXsh8jOS7DheGJcaAbAG2vjvlfpyFazTn5SSl2Edzkj00e3zCTXMviHU
r3VMgcr1iTGSWKxCsQq5KgD5uOYr93BfNwGtFsCdlXWY5oCYIzDrpd8IMxKvqvsT
rcNscC/E9ZHFxXEJOyU+2AvpQ9jKJSP+0Oxur71fmXO7Tx7prqFihqX9CTBMScnd
vORxMxJm8BWnSoci6iA05vKQ8v/dZ9c0VJ17J2MfnWalweXhxzlCp1rBAevp9uET
1t4zClbu6Kox1HeUnC3sI9UMEyl1HmhISt1z/jfbzuroICUX+WOl+XU1f90J68Vb
wRGD5P1fNdd8f3qEhWLOWM+BiMR2ANvhVgPLySBRs+cYmT37JoWmUlDo48c8FYkw
v+8vdLtPLcjK4rM41rm7igyZlt7kwuz5rOhckCglMn0tTmbcBZN2jcHfdWw8SqVW
tDWaxDd3LtMclyZOMB5y+/PlGmrREDCJBzWq0bCPfRTECZMvNBKWqYzoxeP72FBu
Vh7K7On3l+DBKymuWeF6szeoZQyGheENn4OVB6z+hYL89NNJWzRehWAgO2Snwd/x
xy0InbIpWTGx/3nz9kKGrxVanbYEC93cz5oUwPmRf9MeuNz/lojElvI1wycIvs0m
nZ/RUeFUqWUjqJg929Jxx+kICuTv9HwLrDhvMnkkFXQgogqTXQDJeA5+J1k0nVi6
+DmR4iqRzKmeAwwnr3SnqbccRPRtF/h4UB5UgT8s/pa9g29451iwpskmvmpWdiTb
onuROCWAjGCyEdH1oPw1JYUUMWiAIvyU0QDJsjfCKGOeX2xFh/oYLdxM1oBB70i+
ZPBK4DJ2VOWPF53Sqm3fU2xpgW8/XXq37HYVwOZaSLkEcfNXrcgsGeUINcGwyZ+/
onENdfgsSoo0bspndv7SndSFSfMtrt42hRSQNAoiYIrVdUIojs6eG777JeemcHvd
t9d5P/3izhMB470wJeJbU05GT9ChUf2g9C+H42CaiY+Ic0Hrppevu980U9Ehg6GS
R4qELQXwAV5MRsBMETYgAF5RR/nM/ZFgq8taCuic8+495nXoaQ8lv2Ux8a3ktSmi
6LoDcsOS3IgNEo9jp2jiQ14DFBdh/t6W6xTxS1FOEoRB+KSHC05CEaybkYtyfoxo
+7WFS/VEUHsIiwtWHCQ8DOlf5vjpxNsW9nSZKk1c4jcuQBpBl0ygTKN2dVu8F+bG
CiAsH9LPJfG+YiOZjnExv03EHu6ww6AKmVpCjVyR6U4fxNTYyDQzsxKr2Ff5+WG+
TfvODCpzCHGd+THh60Fzit1Lg02hJFi+WqgkTC+tjzvKbzEgrHn04XVvkat5qAqk
I/b26xh7PpoAhep1FaQSwpL5itR6G9Zf5vsIr4GzFS+ItbHwuyBNiUazYoVR06hP
YrGp72FaVtBIYY7DevDuTlfvXnGsyQ1mqeOUzXeVr63M9AjecOjFJSsLQMgxgJTz
Cuz5P3f+6NSLHsAgzPLeF5l2E6J17LanvJHb5/mYruJww49O0hNCCb7cboJZ9pG3
BADz36+RoX1XsqVn+d7QpbfLexJKSsQk2sC8MX3Ps0Sj+gOOCUsqiTtOkul787De
MCksxUSFpv9AWgBnWaDRHuq+cNLPniukqwQb4XrDsItkas7fedsHlv3Y0jnhmq0Z
A6levTwxUIkrldWFL15xTvibO6Wb+p83fUoH2cv5QDF9B/2fjn7O+hvL48iGzOCg
8+24MkqQPFye9GNWV7uxN1/wBqb0wp2HpJHpnA4MbcjxEjr6bmbUfq6owrXn4g6h
9+7Yh7fF371WdCSp1OBmX6EbPri2bEQK6AGrtoTcCQXflrEyQzRxahbwaa37GNf4
MqJcW7VVWEpXbX4zxOZvOS408SCwMs5Ty/frBppsOe5hsOUlIXY96TltkINgMs5A
7Y7XHsqX5MBrU36E5Ajx6yY1ow3L8sohHfvel3+CPNsxtCBnoKoYJdmsUz0DDKnC
ZYuIpqK6yIxXLkxGTTXsMZPPqN3C1yFN2FasGsutESJ2eOawcoDnJb2eGfC/kbCy
b3GJybulQY18rDe5JCoX6iqsSHIr/882qaM9Z+euxueptE4pQ2Lx9587RNfwMsQ5
uE/TQJOAjPOozbUGlb7u1b3fBWKPRLdeLKT09lAxKi6GS6RfkbWOX0OKy4ex0yjU
QDe8zQaWrHEtzxxdqMbmGLsEAtorFixImeIY5jYpPMqaUrqrw6k6682IXXP9VP9o
kxAz6jTcwj7XtKvzM1Qg43UKi8Hg8KoqT1LmWzdGwwit6xP909+XRuI/H4cifMmM
7UtMRbjP+gM+ZAEJ3GulSvaKuqOIjEE1lb8QGQOr2U8Ui4TKvcJ3Tf333ELM+Q63
yfvCXyTSXBOsbcXTcb+bHY4gd0i7xcXXOiji5wm+kSg7IwCiAhNNvEHHPw424m33
dEnyylIsLpyAYjfr1RA/7rBbIPKOdK+EsLoFD2ItkrWDuBUuXiuoaRA4T7yRjLQb
3AombhsBDcGx+fpR6L4CPMquhUlsQTk5o7B9NoRfm1ALzE+TJtI9Rp6NMWqVT+uK
1NXEK3PqDbyyBJn+VNjw881MlnokQlIPKzXnFDz0AKM/fUswTh8k3HjjTRGyFKgj
q9kt6exynpiyDzKghVcJTfeo2H96PRT1gaMx+147kruD26tkSzxmUMFsf0V31kAL
+0vpVmS/bKYZsH8ALt7MkzQb9fH45tz4fgK2XRN1HdgsDdi6S8hZftaEAJoDiOEv
q5Kqnvj7zUSfoUy1u/Z8gGmzqGZzwA3IXKLEfXt3QZk3PDhDcpMvQtEWsa1IjuJ9
ra+7Q5uXRwo3Ny1rV+RCNTVvTHXIzCpLcdclPy22xXqgY5GZ3spk6UAut4yrqIvO
24uUCQnKeLT6idVn24atos1elMNeo2kitJLgAwLXK5N4q4B1PiIxY6NzVtdFbPHP
Oqak0+0gxxEyA4roLderuuzRHznOIwHEZhKKk94oukH/lH3H2IcxBUxAbN9ayKXD
p6j9As/Y8IAqoMQtTy392yS4gGuPG2IhUkKMGZtGkZ9caTLL0BwuT4f02a6mCkth
2Ip1HfEFaXwJvPzELbx+043325CQClKg8wrVZigwcHlKiwvsnNY7QjKjlzvTDwCB
FVc2Ow6WWCvcvwZl0Qt4fSwEno3az8isbFJ8z6PLpdBwvNKsiicEoUX+XEJrpflR
UMRjovJYEMkb9XkgPR5qvX3AukP80VHqrNQLHeUQ2fH+R2SYN29Y80Tf6vViEXhK
KoKTN3gRJkPBx+Z5Z2fx6e1CCmIH5KPKsUOXRCzBJ6PfRlh/XsBwiz9+U1H2Lg3Q
0izd4fiPMl6emgwy4m/rd5uqCDenbWZMx+cGtu0ooNKbmuFqMhpqcURn+zYW2zyy
TzZrxtzSTq7ThSK8PaExB77VXeTIpMMlJiyr3/j8VcZtQ8S0K8aIuDszUh+hQNn4
JAUH8I2GVTn+M6nsGuIaGe8ALP/32v6+lym6pNQb0obbS+59Zte1/tX67zRBAiob
DpSiSGBGEgSPON96XOKBlcbHkGRSc9F81ZsEJ4/2G5Zni4500pS+f07ZXhy8IcG3
vL5riJXJX9bfvQuNQQDKO8a8qYpumXBbcMjQdkq69oqdEBPeuwiUbpQgpkhxlfo6
2tHcw1lSOMGXEgDVqymZequv9H53HxGrHIeiaUXg6rlLDOD2JezP68bW5ck6DT3P
ayJAeSNC9NQlMnl4B8ZgtD10k0pjtEx3G4wVINMp5Qk7zNAzj2+wA/cOCgQLnr3F
lRSOajTaC1QnvEpNeRJmEcuzahLnLZ5x9+IsshcRWmGSzzOhk6yGFb7Oegf6Uh91
U/TMxoFd1hjyf1WRJ0kFiA+XPRAFhA+hztHLPDF2vI3cuphg96lR141/2+GuNHyR
1TtcPWJuECuGG0BhAqRDv4rfb60PcGOVTw5vOMI62c9ex55hydgFtTIuWkfkPXCT
UhvJlRxG8Zgb2TUJPLgwqdfgMTI//G7m8E1Mem11IAaeGDRKwRN8p53CO1gNC4bd
tiK6sCUrf+qnGOe8jalupe3hd588GB41aF6wfmeWGkl84Csuv/0PpvG8duY+p+Uv
Tzki0Nms8kspGzUBz6Bvx3w/0Hfxkf2Y6pDXskAgZbM/dIz7hFaJRIwOEH8hgPyS
YPzMF9nd5osfq+Pg4jSubUfH4UJffQatGwevTTv4GTZUwU9jEmCcCdHv6SEVXydP
aRBM1FSEE+bQdG0Y75SmOSAIBfWX0LR+hfYYqUzQsqG3O5qSbk98JzGNdaPZWjgU
qemztY5spHIS/faCpZg21Q+gRVInNAoGtM0q/j3HHunnqexk2nP/GOHsRLldDyIR
MHaZAxhepJ62LHyCVOcMhJ1Ne3nmqdhKnPQB1m+e1r0PFrjsBOysdNn9QYiePwXj
6+6Fn4F2YcF4cZddsmh9Eem0C9KllRo/GH9sxEoFicrOS9GGP4svpQwHy+MVDFkV
Db/2uRvwrsqDjKa9+Du35MiaxxRndVk+fqYerLMrPtKT98i582TohxqSCQI1wzW2
PlmNAoJirPIS6aOt73JD8bsCZPkfx7aKNuFPjFSE3j72HZ7XkyDhOt5awBr2cEgp
NgAPpDRC95dYv/h7AULnkptIsP1rzSXTOubsGOyHKdgIGJTlvuIOMYVm44B2Y9v4
3VzqvsbQ4kkIfMPSMGveb4o6JXrocxPHm0at/xv/fsLuCbjTLFyUWfW1wOIcSUvR
A7BjeRpLP8gwjufeddS/4rJa7cRVSGA25/7De2oyiwJG7pgnnJTfJ8fAQDr25aEg
V6DD66HyDnvKwP9jiG6iwaAJ9n6yzlRB+bZqx/B6YntAygp+fD++EDSzYIJsGKHD
eO9tYKX+97kcFpFIyleN+3HAnvU9mEbc9QZT84K664sXn+z86lJnxNKjL/KozPDD
MRYUiJdW1x1TrNFYNsraMe/U5TrgAts0tf35k0FbtFY/X307V0LHMAM1+XA/uxfI
G4MRRENRypYQ9QlSSuhPC/7Q8McxjkI3+0uHR1OlAdYFYeD6tLH/yJ7WucHiS25S
SE2OGY+Q8tTNJiDTtPjWV4TJmiY4gBoARuTOK8vDhZBmIVgNLtG6cyPOXAXLmIN5
pDEUv9/+d2hvT8vbKet/8Z9BQrQn+MxgpPqbKbUsopnF/TyaVv41eGsLBE60c+bQ
kXIgrTD1Yl+plika7TZZVrGGc3LaiKGqC16gS/VcWNUiWnBP1evrD+Ow1YU+pr/r
vhk9/JaMLuNHe4jidlA0c3qO7vtDrrBQTq28wTc7R+p4SJyEso52m7ITIGmHgAZM
hUnflxcPhZXdLHNCWzF1e77ksARW2WsaZMxlNC7nLvjxBiqR2zumDYQOK6IgN9BV
RuigvjP1YDmTWxIcBbWEA4u3vl7oc2ZKfMj9Ycbr6ZmksPlJZ+BghC17e40femfH
DJKQjTbcVG8FDp+tCegC8coNk3rv9cEEW2bK9bOGwHmSjR7ptcgswysnUEPIvyUs
81hVox2dSieGFP7JBz9c8U9IAwLsigih81CcmGUnXlWGElla35M15YmjfFEpJVl7
vnoliI9/EM5RnvhHqeThfSLiEVc3qVMn0eNjvxe5cg1sHETQP6c5HX5IfDqwAJJH
iiD+3AMbXoliHixs3SNu3mQ00XXrUD8HTqhTRiBkGCu5wyPlL3POAnO36Ez1p940
hfBk79Wn0qtJyZm1FvXOI6YRL6sk1X6FMbSKRIF+KRRmRJLc16Pva9pNG5/putWN
j+aXwJwanA6sge8BpdugKBpqcUc2qQK1vE5n2tX2pnSBk2fzOP/q4kRUSG9slKWA
wybWzVSlR+NcuP/d1OdL8iPiM+6wDkoCDPEnrbJF/2k5FKR9JSJOi/Le4PDC0bh6
DWBi4itjIjQ8Bfjz32/b56Ib1lyNOVuP720HdDDGJC3RjGMFSQyP/kRXjI1acdUI
TS4xIbBAfi1WyBTUIrvl7sVbGT9vwUC/JcNFOxfIhOqjVd6fARXFKuLkGHcC0wby
Q0w/kDpdF2GvlfQ+rX4NWmediRry1QIqHptRhYrKRDohJeGjT9fmSTXOHOcYl+Q6
4PUPW3nSoFsCTgQF7CzW9pDrlgIjlj8bS58MZKhHS/7OgIyfBzfHG9bryu70zNeL
S3koYfsHK5KPE4YvkUqnS8lXAL7C/J6A7V0lphyBahn5a5LXmPMGKmyJFnxRgKrM
Z60eNiLdKjj06B6mpyHD4sDdumAW49uhWpLlxXar0/3hUbIxwfs3diEeIhtKbDQe
grfSpkxnKs8jwODFiLWD3EDINdcj/9Sb9NnRsS06SkMkZqtwzZcndqZpMDOdG9Gi
adWWmxJIAlJ92+xC3UQ+UFrZFc5X+ZjGlldLmDZ1245MpxzuBYq+qkEzBb+IX7LQ
1YBFJIOqRtzDeiQxEJbSHOaWPJ6InjDjY/kaczFGYpe5GKDUCAU9dChCIBq+xNoN
6RDHIqsQWMUMfkRf57a1pusWTnDLbfR24pqN5BMt7+eKsiRmHwiztQi84UswinKr
LFw1+V6DRTc8mxLESwjzjM2cVaUOjTdLgO3k8FtgETjt4uGYbVGApOQTy4ZZTaQ/
69ZW/AmJsm2gL06UKN0unO9Ug7HO3ngbVT9alTmV7syTTEI/8WlQpyecVVsUpi97
CZqRSe1vY3a/zjT2zQjTY6VWhglnL/R7/jr+ZBBNSbRGkNgVt/faHdD7bSZis2Ws
qMDCaNqnOly+B+atCjkgVcwj6g4SFR4fiQI76XRY9Mpza+4tjnf2w3vO8I0Dc3tk
FyE6YajiBqxkxwt7L9jLhuZ50IVyjQDl2SYmxWzPrxM7hKKvOP7enMaxVTbxDcJx
bDkNBJr7E+1T6hJqCaNTHfaG2wduVe/LoVNpSmug9quS/Ulpdh4NeZDCjz+Le6lT
WeQ8XkMU6r+Rr4baRDYVOf6KrwOQzXicJ/p/+FlrwgtXc8qCGyieA5WVaqbpANpq
fVcXrp+kfoM1F9f+akY4BH1H71XdxIsYrsHdXoBNOT2YOIo3vu4nHu5w4tEMgrXN
jwGPw/gdo5tnz3Qq4bH/g69tr3hp0A6noZd7IyYy8EHb1AkuuTBiOBcklt122x38
JbAqXG6ETmk3ZxYyuIsnOQl+B4LWWZ3qnzGO/xd7Db0x0SLgST7n2BAMK/NBiDod
sO2Y4EA7vVFaq1w0PFVdJXYLmyPOy1c87k0alW483baPJmi4X5F0w0xKlDpjjuAg
EJe8sgRd8d+BDHXkqC6F4S+ucnAfB0scN70//G42tBur+IvOHvJkc5tSVGqBO5pC
XPNZiYFLqA5ME8F+N0I1/317N34XJelhLxtIpqmiy2/q2bKcOiMhr6T7sc5+qIBE
mWS/ex+HFJsvGNR4aVYDO+LHyUJsQNz+lXjmuY1HBwX64XCwaohXYgylWinsMoqY
FbMBuugRJ+quYejiiz1JuiS1hWv1BNMkRPZjJNQdhVb5UQji8hZ0t6qw3XBqOmIa
GZBeteU4AkzndzbRyAiII0Mr9gDrIyJ/z17FYjZKc+b4Ktm0Ufp6DtDKaIRsxyhE
tLVKbnooTjxrfrAFxQ8bXhtSyPOCuHlsOFfybieYPkDaIOHcGa9c2jE4gFFXqXYG
+Fx0CqxTlNwQWLGGzTp2K0BhgURL+TdKbIQsYcpdiEaxBLEK9NQbDT5FE01RmE3Z
Fw8pqLEpwNBmGzg0yZJ5l+dtDcljhN2Nxvnm4i+YXXvoDgSAIP1NFmJC9/UNwlW7
0Pa6cmU9ZJ/vUUi3qWMU5EyxLrsxzvh/kYEcVWdqLrJxVpySp6YXv8HTIt77GD/Q
nGgydEAZU8xroyhVAn0TtESfzXAW5awJ4IhBFQQraf+3D8zpKgOfMIGBxqxk78nc
xz39uiiMVWKA2joqgcQxnspsN01w3lyU9xD08kba6lsgbDpWy0XKrKkrXR7gOb57
nQRk72QRNCRBk2SCrVhswSui/S89dkvkJVz8HLmNdBX4dfIZXsvnKWxYIrOjygvh
KNJyh8L/zatD0adk4vmwFj9ye6zpXKG8CvGAgkKWQg2TbwSIC3Xq6hSFYJlFu9m6
eCxZ+raHAp5gpVRO68unA3z6jC+s5mQA9I26fz4lKJlasbSv3UxYFkJAy0rIcmS1
k+vw+/U3mlmr1J0M9XDbPLpU1VUN/5KDuvsxJzKsozkQitK9Oy/z2L/8GggiC4wp
xinAxHJ5GDg4JYQJz2WIxd7WRncxNkK1dzDNLAQNMCvB/NxZeN4AV0TF36IQn/Ed
nUlMeaDEYixnKBVYHGcwZVkNCXj9ie1YfSnRcQrKGQsTTluRC9gYeRfZKbXXSLGC
bGNfDZ7M2gk4pS7M/I+KCJF1gbME3G0+J5SiTmqM7lWTGO2YyrBLkhl4oNhYOMM+
Wbe3E3/FyE0Il1+Bmz/cpwG3gFbxDoUFhJGpDv1ktWbK70QJOpfqBNpZUETi3bma
5kuQ9tTaPtJmlKFjCAZRAaICsKi4g40bgdl9L024oIxLu8IBVW5JSwn2InFioU3T
dMxM+/fTWDokib38UnrOG4Uu9pRz15XNEKBFmTW0BeTrWLyBaxyR3TJMsKI5z/Ri
pHWGVTV/ZnEshfLrlXeBDOE9pH6kPsw6gyyipM68iALmg9fnvAemoUioQMznwv3d
Z/12eKzIMWcBjxLwGD+mVY9ruhIw+ew+zY04imcKw7hlJrnHSxqkuq8Sopmfyzdj
2DC5cIFxMPA6OKy2GzI6C73ibfS6RY/iJrazhXY/EmOHCrvrvH88bu73OCmJp+VX
RaL6dsALGyh3GTnz+Gj8r3aVjYXJtNWG+npHLWcC8RBblTQokzCdtrVI5Ra5yInH
umMTjJvpuYkeyhRMCWpMlwTnWL+OWdQfA62ottJKgKm5iXcZ0bboJEkaoFMt/170
zZBEgRaJcY+ccGnxzBpv8MLeURSaDclmidhrSbFVSC+sdklVBGHII8GUf+KjVdz0
xSO9fACVJVyqE/B8TFgkXBCHZ5QBillE84QfujbGF7gBAXooZWshzx1fnMG+a8ie
tWM+gCrVTPtWM+vOGjfdbybfScPTeVBZ5XMfd4yQKe1GTy1eWHF9ALi76eYtoFER
/p7uAl8vSgsBAxbQSvUu+FRMolVzzPgH6lCIFnQPxcywcPFE0/J0jrrGzX2Rd7Vu
RDz9qUs0tKBOFVCtWE3X6FVkpOGLYrb28JLji9gPD3zuGwFuZSDRp13NFE22btk6
4qsWmIoCEhZD91hIImJqh+u9HC4j8js2CFkV4tcZ/frxBVN+lccBO60QJDWcNdNb
AdM9b72/PDeVecSgq/a7NgddUwFsDOqutwtPK9icvtTny3SMoWCskzGdkP1Zxddz
Xiu4P+iIQnKuz2A9gDlnsMRp9c/lDncsfZmnF0uTJUDpphhHcd9XBl0XUwk3/Sv8
y+hjg1zE/Bg1GEnelfr7VP7bi8++O+yMdeSI8ZhmlmvoqMZP9Q+PkPlzsJOBVXhG
XFam+64LA04Q5Q5Vc6eKc4BUVIn22ofu8WnPRsVAW2kQ1HfekMoUGn9MNQCatxG/
m3ZE63ndvqsaa9daYTqOKaTOaSIFMTAf9wFdQ3fT/5rvL7Zx5WPx5YoriSRRfxOn
3WGeQIvZg2fu40bDVuhPy4sGTXXVBnwRvokoP2vY6T9Omnx/tBiqH0wtlMOdN0It
a81Q4Z3ROFTl11mwNvKyWWE2N2DsRpL4tDtIziULNZoyZPo0zY0h8sKi81rxRnoZ
PsFHkJ8s4M0RZV8bdUUO6NSGo6kLwQeXr1LwzAtjsFCOt5y2arVdUXb3c8uycQh4
oGJ5NyjNfaNl1L9nuuKbCEbZBDcB7ML5ivHAqbdMtlZLOWeZxQIDH2owaSl5pGni
Dk5au6K4Dx2hcLoCKcAUGx5JY+sJVGbF+yoIeiPjqcXcR7RZO2AZKK1qjtmJ+NhG
TNU3iBEGcUHVGg5ndNT9rTP2+cLHa8wFSfdnceiD29MG2kGQ05FZz16leGsBzXLW
mH4VHxxmQE+aCAgWj8lwrWt68b3APVBjWvJLhSwgkp3aGdN4UqjdfDeIkivdEVZg
tElKGUC/uuhzknV3AAhtL2bqtpoyToFhBw//FDH0aTQtN6J10m68KxomZTK7fTOZ
+yYQeF7Qws9mv2/ebHB0z7zsEoIwRfxlHOH5Do/9lU7L/QzgNF1Qw67n3hU+sSGg
oR65AdTQonOIaTTzIV6JnxwmKFue/m2oKlGbWT1OQz5lwGaxioY5QiL7YAT9HNGh
4Z8iTQhjO3JErvQxLI2fYLlGPEiKCjOsKtyXN2gMLNR3iUUatVKl9FCl96Mn+QUH
IDOOAnbq0v9XhbAJxw5faOheK3/huqDb+N8j5CVS1l3A0iPvRCzJfoTguOZuSec7
lzGn+lG61gJHJqV081o5xB9iF/btS+TO2nOQHXO2mKM4cV+4oYp7vwemU7bTkdBw
fArluqg8EQF/PQBkW3Gdb8K4M/MssGifNUT0xsiFbkLYLvhLWbAf1o8LR37bt/+O
0ZWpqiMA6A0qxG0ZjykHYgAnD26+4VLto33PKPG63KkEBTFtv3WYM9owe2cRbxCK
EiWETxLv6IqgdEErTIUUwLn6B+FwgNfuaZt33XI+f0XuzqK2VlPkOMqV/H3b1r6H
O69FunmJr35HQFI75oV9T8YTecrpcYgJkInEdWlTZa51Qe3h0fUWKcTIUkQr7Ghz
64vS76yIT5mz8XGXULH1rjZ/nWYZcZjGNPgPd1zx5Ldnk9hoQg3Fo9erfCY8w1Zo
yh7AMFe/qRvQRjp+Zl+ycD7TQcr8V/n7cGu4SJZudM5NHGxnAXSunjCGDYq190KV
pYryY/xhOG6U2qy0v2Z1r4lNIDLir5+3r93ohPTxS3I0RzSZFkQZbRSqEjgzcrIc
8TMw0GBDGcKZlAy2OW4ffnW8i6L3rnnbgj46BuUAYzfNYGOaSLzn/J9foBTWoZZL
h0foQehEfUe0kZrCcEweiKkyAviqvsAjpbGw0+OYpuQj7C8awj5oJBoaKDrfIFG9
aynhnhOCwiJcMvXzuw21Vm0JPxGoKWYIBwf+IGAtWQJwk7JONywHWqVCIfxtoXCq
PGndGPRVKQ/0uJw2Pk+m6v3SfRDZVFXeQz3XEaeb0fPlColqMRS6EbTu/1ILek4U
lel9ptU4zOSqfhbtGUrc2kwfKRKCKaq2H/K6cWp5hp1c1fPlZUYF/PqiA0o9UvIk
9oJS5D1O58+60X/3EsY2arWM/KjFPWkDx10QAi9DuNx+1EeQhFAV38eNqLT5NfZ9
tNmXp/W40pQEElppnUOszrrq1ai48vq28pbyjawPe7LRHx/sjcQZDT/yKhm2pwGZ
gEUctDKtpmPkDaos79pMRYw60JHeGKybe2qJAT4jMRwAV5agchR4C/MNYl7fa+y5
dt3zSDforUq/IKc8ujp9bNSJ4DQaKH0c2/QwGikp9gNkTSWOoe/ZqzDmV6ndGbSS
zmiIFnFFxk/8Fnxd5yJTMv+lTcnF85WT4YkNC0SwBQsKIZLlzhDkQunZfuQYOKnj
5zlQEuGE0eaT2Aq/Zsg3dnUn+Mt7FRoWgvaeWL+BuU/HQfON7U1MfTTlFN96M3dv
bWMuwuZyRpd6ucAg8fNdRmlYDHYa6a4q+5qvNnSLx33/5InyqdZr+dpuAnUSrC4Z
Q55jS6L7dniKfHMDFjvQdVoSWpFtY6rM5WQqX7ngKLocNmn0kCGKMgFHhQ53YMnc
q5d8Eu9UppS61Cd/FNRiWiZc4dpuBpHde+1JolGB3oNnP7cd7VrUvzC3nl82M80Q
srCN3jK6cvnkwSvssYW+SsG+upl0aAsaWdgvaZbORjesxNAjrwX47T10qJaafqEq
8iBwzLq3faXLavnH/Fml2++w6mLbX2DjTkDb/XxH1xrYfoVwcIYGO/68NsT8Kbay
5AKh3ycagSZAYwj8GFsyEwMviDvb79DCREiFl0pTBF0qr/fjfRTccRcw+hqdrVRt
3AV+l1OkoDYLGGWVvmV6KK6rbbCsxJ5qlFGdjN/CPIkeN1otNoebwCgSyN+aCRku
VRkOPS/HLKMu6fZrEYHgK/ATFOBe0KocZMVgrwqvTZSSzPHRjcwfLmoan06XdXwI
Xt3gr6Q5BBuvep2/P0SUpEr6j1tM6MLpsRyOKltaA3of53j5gSWf75UVi1asPS7s
vtGoYRAnVr41qI36W6mrbedh3Q43HCnWpWOg/5zlDYjunVKGMxMQ+bNuy17m6NS8
Hdsdn9EB4xo9h68nRR5m8Z7TKfVn//SQ56IsUucIvWuDbvbwM8Yp4Cg+bBjsDQHD
F6PGuYTvJGnOb9dV2xuJv2Q6r8n1crFGA3IvtzfKEvlekbF00kGuW872jclVkP5R
SzNHJc06duoNKP9J5xx1wujdwFHJnACF1kY9wIUJrHF89N62f8twSAsm4cfjYsjB
g6b+WpO5oMFuQdCtNJajqcrJtwjaD9uzlx5GVG6pWgi/PfXWezM6JBAdPHCuGxQo
wEWBfPTFyUXVe7wFF9O98XK6TZv4AtunfaPIOHrQ0p42aXTN9kMvnXpntNVZo1cT
KCNozVMQzc993qQXiQ48MGx8ofQoDsyXaG7ZPYYVeamOMnjLBQUMTH2dETiymoOP
sYPtK8ZXW2s0fWRvbBblECDpI+7DhxRDlbWx7w0Uw8HgCM8dmUtRGSxB+2cg2yid
7Blkg5bxDETBDUP+J/0MkcTO2kTc5Br0lBzLTVa8Ua4+CyoUKu1fg9v5LXAUtAqZ
xCJv2eqyW5Xp+OMlPRcslDGI/w6vubcaP5qcQNu6Jy+NBCY2dbme0jInX9XUbs9o
phQDVTf5DNts6yajS8yuT3bEbuNdkeMSZxd5yY7Jb4rIdcdg9Z+TAqTfRdYG1TCV
vv8+4fOIWG2Xi8FqbYAOrtiqHNGYIKBcir7tcBOU3tmB1Zm0Ld5obi94KWdz/t9o
vf8td5OAHQEWrpGCAT/VLd6GO0bAFRBLWvT9XDP9yVOsZIzvp3LndYHF7Q+DqD7h
AdvyMi1Fj0PIFXwSmsjG+UjYZgSJXyUTxLtHvIt70+YUapzhoJVG4AYquXBSBKUc
KqXCwv+Cs4suTO5AB+tjeYwQkNG76rZBK9crdv/JLpVqTsw9ra4Qjq5FpSdLaFji
FLGAovYF18VFWbpkrq8BMomOOaP70cYgm8jWPOcc4HAddcOiq3hHtxNkVIJBTWjc
03JlmMS4f7s4HqN89yhCKckYZkiLmXIEeEczblSRUbM6pid9nj6DK2nKTU8Qlptf
ta5EuulnxE4KdtN7TbBeaK0r/DZyDXtNjt/3/V/YKsPBmDw1hJIGNbrKDo4IJG8S
AC6XIkcVsKcuynclBKHpejHCfYGuHNEWuZnS8FdZiAjOmHHIMQE99u9EsNnyY204
v/5dsMa3+I61St6j89y6k4o5yBx2GkQD6ozCFZf3qX9dzsjjC7JRJ05OTD76a1eN
nFlnliDMEqZXuaWranFTiDKrJ41prvSATOHXZugewB5fPGkcIY1C1gq/sY40lSaQ
mKP/lkhw1y7jfR8+piahAb2BS4eKUO0EyFxk4NNactDfqsSmallNj08a3WySw0QG
dghXbTT6AkjSnaRl5urq8v2Ugt+7BhyOh1YP9k/qvNYJdoWNzU5zY32dNrlO89z+
oQHzrpCBuseaXPIbKk7XJrXPjqsEhmHn8Evmm/iS4NK/0CIuzY4+eTBcWhMa0tA4
4URb2is7VNMPmoIVFDec4jZq00opm9Wmxj/WS5vyiuKqqgce7/gdf8JWci0TCdmA
UJnTMNDwZ4p0PrcV7qVODHHfVK9UQHnj/2H0/E41QFhb26vu+PaxC5PYR8S+cJHl
xAIpwyAL58n8E+GYTiOPC4670fJjt0iOBp7Db58GykveCxiPWOeQGo0Jd+jcY2mH
DL49r+6PL9w0/bn37VcF5WahsDoLsVs9gOELteRRzC6gncT0kh6gEEG7Kf/+LwON
t9NeaRVUeEFgjAf+la4DS7wFmEt56+xVF10bDdNgz5HvTRanL0j2zhx8t2cxOi1V
iXiLpJtByLxlVOLfAJVBq1reYEterGpWwt4pz2gQLpHiRWb0dA0fn10JmMKmaz7i
3Tkm+yBCEuSUKg3yybgjkPBCSiryQGUGZXCvn/Wc2YgLEcjjuUoTXn4P16kcNctw
AbwXiaoRX1JrsXpVSyCXbk8Qbkk+QQG73iVSHRFWkiqjx62C9ohswp2FKgIkYaUe
IJ+jCRnyM5vC1e1rwE20tGnDbIfxoIXaaHyZsfAZbELIJpEI1Ttes12DlGPGSunT
nJAHw2XlFZCvBi3Y6NwmNh83jDZlodCjwOltNAJjyUDPvE3StYIlx563lBUEp3mm
Lrh3z1fvLddUj2lnqBPR9bH++KQhn4DV6VJk1Yv91BuO/UQFFBXrbMnws1CqutbA
lr6yZ0y48Rnhw26ehf5cFY/vXDU7q6IY3qGTJGlOQ/Db9SyUwQUqDtMro1OH0nCy
lRszmZtxJV+PeQPdMCmCcRD0fk/KTokJtiQ+CXDNLWRRwa6IYqptXFeuGsoGtbEq
uH/vVf3FMUDMUnOAiM+X6z9NCgh9eCuWPwlKB1moXJv1QuZMKkuqKIpIhmWorKsr
j/l/sErTgTqlujS9G0nwcXP4cZThD1xTSafZdE6mUZiGsDBbbuL0t9viUrhzQzoL
R1iTXsZ3qrGdc6rYrnpWboYo26TdpvaKkjbjkaKbFu4PLJZ4NFSHZAp7kxVmSKHJ
U2aAebyY3zL5oDrizwqCvOA/jcwkSVQzjrsRb+MneUqPph8pDBovFmQpd3PDDHuK
SFtfOenGFmbYBUigEM8TORFEekZ8a8TjSvUn1Vcm0G9zwi2RV0m7OOCsx3zYtagt
tYE3/M60bb/m3BjJP5h3+kGgIWwE2461k+nUWH3YWpC0wqaQqXPmhY96fLtS7Nm+
w93I6WpVaAu8/GnY7erd9uierV+xpXZ2hCvLOBmCX0ZKCxUt9OKkew9Yc0qIgApa
gfXx61ivYH5pPvyrj6zA86MgT4vez0tilMwqviSMuctZULLCE2PglDm/pUskF4VU
2k9Rt+YfVawsqvzM3ccBlUkMoBdJPwkq7zjBscLXkm5g1jghjpzlZQzNHgJvAsu3
6XUmvYBMkjgA7TEFDhnml84ExUqLjH67TGXhuoJvCaa0fs6E29kKxvqtrRmsZIoa
TskWWRiFAVlUYLQKBVlublSyEYT/NQMwnIRGrOIGIR/BsAqT474TEfFwS+x8uB/w
6pK6HCNeSrXqxRZEaA++r//NBT00G5hYwEHI3BjFMD1gbCeAukiTWTGq7Jxt9OX0
iqroiAJPPr0FqjrOhtPM7smKx12lp+tiI9VVgZh0OD7ypnSxB670yHOlna4zx3Ly
wqZAG1Y7EgcQCE6Q3APJmmVSEW3faU7dBT4xuYS1G05GRH8VwmxPi1FGdmZuHPfg
oJwquQClC8jcIgwLDEkYXlnHcpZ8hc/wsCjF4LQXZuKFeOdbE05DRNqYU1rq4UhK
Uitg/tveXnJcmkwB85UI6lJv5msE6Ws8yESYjYcuEW8XWSxNnsYud+1q1uBfBW9N
rJ7HHUIpYx0UJzv38eHn4TROp6VLcexUBW6qyK5Q1Z3ef9j/8W/MXEajqvUWdYTD
bGFYF+UZwwJg7/RsFQb/JgwPuxbXLvZG0am/euT5OX85hI2a1KfgfFaE3rUSIYPY
vW634lUjLaIQFz8AGzljMYLBMuyalpeXfXI2568ZUGjm7eMt5uaBwXXnuaHmbwoc
ZqcDzcVx41mUxln21g0aJeNbf6ioZV3ug3Cppx3kAvqfsWT6A4ahhS65v5aeRnle
L3QRWzVMMX4Fa3UwlAuxbME4JZ7DiIkPV8T/mjgDmxrDtY6UQEZX2povta1ClVRt
gPD5aAbugbwlZRZLNrwUnMb+yEqL5nsu/89nf57jpB08/62qNa9RvJKNAGRjP0M/
a0jFKjj1U+m3k8A6jw6Ku6btOaT75fzIhS1dBi5HN5HXxtS3OEPyWVCdh2vYQssW
Im66xQ6AMlTvGMBQehLu8S/teiUFvn408cCgXrtdG2xllcgu3Axz+42mX+BSy9OL
gARy1YNq/p/ok8xibohOrQ3ZX5MNerU5DPBYzYb47yR8zFUFLfa413kAWnJnveWN
nyrn2t58kvzD6kUfkoKflPxsII1BtkITRaT1cO3nLvwaiMbdPry9Zxnqd8MXHt/V
Cl0fcS4qSGX2gtKuPtw9Fc2TU9lVShaQOZ0mG7e97woy9qH5tWN4IaVpxTVlRH0+
1ZuxeEVy3YlvUlBKufFw25zc2AwcMcj4QYxvfHFKJWKOP+iTLawqomf1FVPpZ0iI
qTwzJz80I2Uh86Pm9/dg+14qbigNDRljc93zcvZ6zaIdje9CYyzH3QsPjmZWLAEk
308X0JJ7RfKw32tHmSk6RLbwP3lYWQjtPswij1Pc7CDt4c12ad73D4TV+NM/R3yb
g70rzQz7uIh6r+Uft0u5W8rG2+6lnin47UE/5BCFuW5f0Zur2g5jSFyBkx4U5wI4
wpl9oMxYZ+PZShtGrcu7UBgVRcQOEQxCrLji6Ew83aL+ucgiU7o3JqZnVd0s9U9d
L063ZH1EAMiDre0LCC1Atf7dMy5Obj8XmO042ZNbG22unLO36GG/elNy4yPJoBND
MXb3STrGbn4N9ZXb+0ICNqxHkG7oFBCBk4CETQEGu9SeIKWLOlmvDCaTQMU5qYYI
NXmm/XEcaJi1/wondhjFBmr1JTFdWupKdglAA1A95bsKmL1qqX8J+/g+txxUlr3C
BNof5+8++5yDIgCNFUu/GECPxlf5+YXlaixMSh0THb3rAGaQRzqVRggHIq/uUveU
PlJP0iZ2TTQTyFJMeZF6iQQNv0/dcxjAutFypS3vfQnwaprhXojfCe+rNjUv0KpO
6nBG6IfHIx5IdskTFd4kAdhIoCBXI73S4sdRTHTjqBT8PMVycVTviIjqBp+lA25k
jXhZDemSQN1cEJwOuj3hAJCSx+hDRO40F6OIzRVIFdV2mfRATlV/GXfaNW2Sehi2
hXwLjb5IWd9umBEhgX1a8SjsuOwZme2zTrfVAmUBw2iCCE6cymYhpighAJ5ofxa7
StXUaMXXt3n7en79nnDlrSkIseIF4zSZxlCB1tkTjP/dvBrDBFMzPnkl05URYQEd
AuObTK+9D1QGZCwvOgITZ/sOL62B8gjJcZ24ub3SfSoJRzR5SqublvAcuPlP6yWt
k5fanIoh/7UKGv74LLVQ/JoS+RqLlwkKDqOETi/dxZJMHu2Mn95KwJo4D3gBOe6v
J7h76XU21JNAKk9p8wmTqxfbX6ct//Mlzmz2YpQK2PyclHqESzwjK2KfEtAx6H4p
IcnlmABIqNYYMsnOZOjAJ6TLkO6y1mJyd8AULJokLDjfiGfbpyDbtKJiFmiky3pS
dMB8SLuahEu93T8HtQ38HHtSMcUvJaF5e3Aen9Pvyltb8xsV12eEKQoXOq8dfVKi
o3jYpiwKN2U/wluPI3WhYREOIGks9Dgnc1HmA9jHFTjx4dL+7T/sWxXhmEj61M2Z
uYQEhjTKV/wxktJk808xNSoksVcaC4zkcC+4iPr/HT7F9td7d7J1PaaiQxJZ44vT
Fe8S/Ndb2Ts7HbIWqxSu0EP9Tux6yUKlc/EgL3+lee8u+0ENwIAkWWbgz4NlkuF3
kYqH/WXEH6UbqOaHjx29nn1+OeMa/drWsi/JlRmF1J8XJ2k6DZCH9Rpc+hjEYvw+
NbKZh0NhrBQX0EqRetvfEpUJ7RF/Po9QtmmtIvq6wA/slU6r3ZCKECH8TjpVrTRR
z+MLeGapWuI2RwedNhzJS0vzPt1xkBjwwe/M+9dTL45yUWn0rpTfFLsu0cnGOiCA
h64zSIKZz6sW5lGyk3PEBW66OKgVt5XNPefV2ODmcJ2+GX2VcSdvJojkrpZCwbzD
/P3ZSwAOzK0GtWQUT9nC2Ghvy8AMGAFQrTYWzQdwRSQxxe4zq9KRxXHxxPMPvzK1
RVSErYPayXWTuVfob3KwgdZa9q/5Unaewd9U+AY0OI4O60eaVgS3TiCAUbvHLM1s
3tSsYLMo6rckzJiUTOsUjlAwoIUD7qzTkAPEXn881eV8iMpfwXAUknjv35FyzgLx
ykVoFf9Ap9Gzk5FkZsZA7oYOa/ucXFgFSn03mnTYZLEv2BrRxNoB1irQ7WqDj6YZ
kwkvmDl/C0eJaRrMY0Gw79bUV2ulaZwELI4SMoC48C5TwqUZSPbrmfgmk7hnG+5z
b51QmtiF3uSZv92RsxhE6XsHrY9TrcC+K/pffPUUrxXsuixQrrPjcALr9PCY88Az
jKgoxPG3X15GWrmanKkAGcUMQfU3944K55sR/jGfgn2zRs9X7r3vmeDYbqxwGl6S
CynsLceAz4Id9nzErOVGFsejXIyMZFofFs+X4o/EN9fO33e+AzpUy53c/XJv5OuK
1QpqxGvBYxXzYHIfdRxPNmrFcgdG1eOZYIX/OauXNKCCA2QoYnSnJJe+vWdS0h1Q
5F2RF9GKXOdL1yuNc9Q0KmmAkROaD7m0Zp61ZEXiV10EBxQ7d0R9CFPmVeiShlfh
N0Gu3kZWdgriRvnkcVP02ca7CE5yHineT/5qPqdFCB1tacfQWyhDrZN07Ks4ZVUR
bLRgycqZ0LUfU0H/NYulq9QyAHzuJxCCx7jJ7PZBLov2TiADOOw1icUkMEfgWoSN
AqWDo5/DLJo6lJZBciTeJfA94qa9eQFFhDmbPwOJFK7X+nZaizSe+7KNGsYd2D4t
sh2qAMncG5LAWKo3KuP2V6j2Sgxt8hQ2RLXIGEbSGlnip8tmJCZSSJM75/4VtMDg
75aAA5hEH5IF29mCype4hjqLmlCDRO41LJ8XtbOS2GvO3SwVrELDaEWHblJgzGmM
B1xYGMvT3OZWrrnXcDTm/CVqycqZ2LBKUnrahZdTUVKxtFPSrzMaxgUpg1KziqnE
QwHO44J+LJom2bZS8dW2Q/ykPZs92xujQngOyt2s27qLzvHm8xqn//gx6LzHw19l
rtygdS0PYSd+sPYsKCY5TOx7JZmMZiB5NFhV2iw9A5ZuKDttXwTLO96sNCRArR6f
HIvT4lcsY5jIJEFty4UcAGYWkHkt8/NIXZ4rpJ42ShHR2nmdFunkPu+3JEPB+iky
iZ7NYE4OTCZh1Wr2/aDsLqKA7vx/qq5okKcVBrds/G3Fv57tqjngViAwlH77o7rV
HzGeUVXo52Pvb3kYPo+gEDwVbnQ1t9PXGBc0iMCYB2ev4wdtSwfz8UCQg3ey4a46
z4mMYNl+IOE5O2bRPf/VDU1VldhaBHtlY5WJaNVvB7WcrxWSrIdc/901Vvov9/Bw
2Yifjmut63/1Df9zSi/zostm+cYWT2va8VD+xYr+MmjWDhJndcQT49VrJl6vLqNc
cWiGPUO7a+eTX3pzfEaOLvW7Wczm0CFftwyhQBFFBKcHP8xbhOO4XxCSosNgaFDq
jXSgjl0XTBh9CULvjRUud99196R8PVhNCgpr6+RME9N0GK64kBNhzBsFi1j96rjR
3V5HgOAxd9LkFfPgTEYAlnDiBVbGlyR+3oVvL1wLAFcn6ovw5vmRHzCR99u77kkH
1n0bQxFQNyGA4s8Ix5Qi6eOKr9KE/t/Z4B3vZrUkUOaP61K9uWLNp8RA0Ukqcwyc
PxL17sBuPfuTv/hV+w99Bzn8O7onTgez3Ox3JlHjfe2gDlyAHB0i4P0DL9PRTQQh
6X8YlBACEBiDoc5f/EHTReHeUiC6oQGmsA5bKJY+GqmMbwRml+EFHEcAl2Ub6mV0
twF+qAdSjUiaSNUpGDn7PjoXzk9dgO5r8/99mtFIQklVTVjXIxyEbUpAgJA2ASWp
Ga6er6gyL/TNeFtJDWGauW+SCJPSQq9/2IQwaurdmyeSnn/cebF2Hk+YxsU+irwi
snJ38qwUvRcC0sFOFYqCmRpjvzB2EbG0mosQHoJqMiKgGo6DzRRkHpPWa5ttWYg7
MLjmQm+uudk8W9uV6oJaKuAYWt73a3uxEEyXn9v0DKjw2cP+Llta53VDu3Y/ar9u
sQKI6sfGYgR1qHDml0jNzPZglaGqGiAkKGSnbntlLt39sF9QphvINA0w7wbHpzsb
neKq26Tkf9UMoCY9io8f+vBCauKmNP9KJAn+ezd3piVYdSTFZ+8ayFBZLGkK90ht
sns5B08CSUILeshdpH8Rt51HJeCgxxaTza+t/Wi23RWiBfx284Jt/1Vj+Rqp0gvx
4F+Q2n8lQUhC5V7QS+VwUPhTaGf0r0kLvLArx2SwQ9FmCwwtb8UBm1ViKtO5stUA
01SLAHjx25/Q5WXPDOav4JLXy4za4WqjXd/pV3zSRfoxYuhCMfZROipweEXoF8r3
6+gWaRnkZL/S2C6LEvD/UL+sFgFxiNCGIkqA3OQQyxOiTs7yWhXjywT4k7BRPgGd
Lc9tp5N5KqeyOWUS+yIGL+ELrq6TnSn8aemQNC5G87EDywDtaUz6qF1V5LxA2sET
PWw7lKEzz4AEwhN8TqBfMB1cHg6PeidF32M8+HqeDYn4Mv5nFJCU9DMKBR0y/iDQ
u7rMf4lODy3BhSa2v7SBDK59oVgbZGW9nt7NBmZ5h7KJ+K6JPmv4m5clp5Ut1v6v
D9g77BjYB0TNwiKnwrf0AvWDdyc2OLi/IHXBY1YA9DZrHYAa3qvpuGWJDINJWGP8
YJIYYOXE3maF04WbiRsi5DjqN4e25icFNWi1s3GY4JV976F+9kkwGDceYqplNpiK
sMOTjo9fh4nMrbOkrgq/dE/qAArb4sMEE2AyZUNcoyf0d2hXwiRF9WgPmCH6JbdM
CqG77rg4gxeJAdlbxUeRfeuEYUpp3rCDFFQsIoTrFZgserSwqW9t/gQeO1zQYq1D
QFAL08v3VYvMAv/rXESY1dEOMDOyizXwPgDwbiAi4v1egJgCc5DNV/531ONRd7ou
ZNx8lKv4iTR4VjoDYlzZ2Wp8uXhzJLVTzQkus20bL/Vo/uePpCL7OJgYFm8k7pTA
kj0cBNxoWfDyhQ5a7GDa5cM8XmNtqKrxQ//5bksrlYoUv+oa2hKhaKhyu3a9ENqo
uwdudvSCRW1mDCnGEbqrYIjvBKjh3xrDw6k2/KWHb41Bzog0DGiHXI9+gCdx/5wK
ONlc8SwmX492r5egHJHj3lWGc5y/VR3/99XC+VWjketswPKwXrEFqjUGMCKtTVpy
2Q5aTwlU/oJbNZI3DQKfMaCh7YQ8MCdDk32AW3+/jPPuXmuMD3TCQ+K37s9RC7WT
kvWqV6lfQmjd6kacbhPySo5ND8nk8KjtygYIyMEMlQXqGFtJTDK+A6gBLKm6Sp2k
UmSflHjt+FzOs5p2z7Ey/oc7Y/c2WyI20W/9MxhENfFBm0xcIPW8jj5slaowNtsY
Ev8TL+FpiTDwiZEZCuSttbCud8O+hcmx24+RmT85Kf+B+0pqQVEGjiGbgsoJxkPE
34+J1E91gWlwOdPcmZLNwRPaGSMHnlXi8xpBuL+FVbbukWXe+04pZFhZtLN74iBd
olEGamcu4pNJ+p/KxXJdXsTebskZD7JmzWxq++wMe7+K7uHWA7F+dZsv9+UvLCWw
Ic918blD5eTTjPLvOf9bDIaXptDzKEwHWWRRapDgTzaeufp0YjISNzjFDeKVtJ18
8hR/zpsXmf5NcH469x9sVtdBQwLBdNb4eVYBVQ7E1wV0PmtTPv/Wlj2229oYlrgi
o76Sb7922noDt2f0TVNM+aq4ffm3LbCdb9nT+O46AVX2+zH0klTACNNkGIHvNuIC
/2wEWfbZdGcbjDwCT2PaWFLBxIEpL2NPQ9v0m94sVxur93SWA8g06dfHCTBpNQva
8U4VgjeiTPffebQ+sXq1EOP+WSgElAlZloGiPUAC0Dxb011j8sN17ai+tD8ZqKfP
BT4fwL0h4DQxPIUv5w8uYG6XRDKb4mwznNPUyp6FsopLWkC0024AN4Bqbhk8KVAF
h2zfSfd2BEVJA6WeGza2PqvNyGNBatnuYipJT3wBLEIcMIJ9D+DfuXYpTV+TTtM2
Whel36AA1P7mZ1xAfN4ZN3e48GVvhDdjUwfie8jZCXxJ53FBZAb0q/C/+rNYPgbA
NrYTMs6aKKsHjpICef1NDrpNJuiPllL9grxlozRL4DoYCL6GG9ngIj45Rlc3H7Gf
VNzU8HQldl/04svFHj3A1aSN43YPWkDok+HOs8UfLex+7EF66MTCcQtXPy8/05Xc
YYOo2Xs/WAQhCNJMAqaD9fCtYfp3IDnUSYpHbUouJqCq2Fsizodfqh7qWXqBkDeP
5iuDO2DIwHsVHmwGJ96GcLlvMXRL1ogN0G2715Z05pdNqHCL+V9BgXI+KMhfSsiy
oXLFeRlDn3ZSzmRPrgTBlNWgibqyRAXlIDA78eR2wAFXKP0UxNnhI+s2+9Hz6Ij5
qTXVj+FK/tlorifdWiQ53ImBH6EFbkgM4NvN/8JuG6SsTqI2FmBcx4qpT+jZZcfH
yivdbT68ONGCy90r+E3AdRSQOxlOVj6eHr+NxUyaNybqV/Th/itXFep5VNjiz2D5
4NfQmvI0OAo0FOn2YMBWcClguREPD/AChNo5eulWeQlEBul3GaSLIXTztIiQS69j
Nf91Ys5LbWuqLWaoBWvz02P3UtNslTag5oMKkPWQzqln8acwOF6cJPlff0AP/72P
cPY2sjAgJxBaHW2gCwtU+wTn2uc3+4IeZndeOIre2w9RXCoer5pzzrJ/HWJyKxru
yZIIGGdX1NyfR/VLyiFCknWPXXupd/Q438HC1eRE+T1TQbqqp/0foVQ1LpTtUwr/
EJ+uKlgHPlnEkXcNw3zRyXhRUL0GJOoC19FbHC6layao8as8kfEVhk4U7zDYUR2w
dBuDPnLcJGAo0iOkcOk5kDkVbAP8iux5lXec1XT7xJWch1MbGiAzWA7Zbn9GactE
YXaFLdwbYSMphkJjLA/LCgrT9qnlF8H9FncAZzXzPGkrCfpbJMUXLjywu9rrrCqc
H4LkwK/xdtqwNSQNSNUhfGlmyulRecNE3b55lyBtOPRjMeTGNKPSRkMmaaRhFiLp
BmisIjux702ieWXHubqZ65QC+WE7sC/2BQhDHfBa4KE5SI5NY5QfVuB0xidk7Mud
eveePo6yVFVYrxj0fGPHWdzoCkQK8Rm6Pq4zA9PuuMubD5ReCj5HQzJJNeWQW/ca
aIzKEmvW+2zEw437nIN4Hj9AFruSdaOyXEP/EjmigzD8hX7tcmI67i44uvPfyD6i
sq5imiC3QcYCrAP3+IODDN9DqIbc62EltB5kTPyqxsALi4KY4/saKl/WW2mQ+Thn
k1KPVnhdx5V2GlT3bi3EtndHVEvzPRkQv8zpXB+O7MSRvjBCAfCnbuJ0UfhO52OQ
B28CES+K4HzTGvSyyAy9ym4emEoj+1JO64JXeHUwPBZYcSWkm/eOmR8gXKMnMc3B
JkxepI2WIkoW6aRa1uF9UzeQEczVzfLFv4how8BVYx0zSXBtcqMN+OH1TViTC75m
/Y9u/KAjw60Qah8D5GivrIa1wC0LdwTJ3TEDaJwEHJKWbJclbzUd1JJnL4soHNB3
JdHx7BW9dXVUSiXW2X6cfzAuTGpPvxGiMeYYZuvonZTIN8dE1GryaT28IjlwBWts
FRNvj/zUzC04AbFaQzcKd9CZAQDUr6KcJX0wWZtwubsPX5lf70jEh+t+Df3zRIiX
ifYwNWX/8Yn4pc+xiTNb6MBNov1bwMFq9Vl2uqODDZ22isiP268HKmqXcEs+oRHy
p1dEUd5uEtU3XMeoVU89IFfDy194VDp8Xu7pqWEnYIEXOyrbfm34zbOz3AULRZon
UdDnKrrF24i16FeoDJjWf83ZGDM8JfPoe8zd79s5knTiC2F38uxOqvO9Q2mXddzQ
mtiHOqqAgLpfnwJeM5WplnFU71zamygnkvOuDW/ITnsKmxjmVkq2xkpnyd8vpj15
1V6xL8DJcAzbtOT9KxpApWxHdQMHIEBOOnBqWYgwVcJKkJMt3NdC5p6ALhlYeaJI
xLo8XcAzVHirFvFMcBuqrpD7KnVKSTiIPNZqPD30HoJt0kqGnhv4z8MQnBAwGK5R
uAeKsXc+Fn84q6TWhWyVUwrFMH49D/D+qNnarpQBxyNXbT+v5xOSbkb2g+/2vKIx
Ma3ED1OFetsJ0jbRU5E+2Gjzk7zbJUH+7ypd2hIs+Gk98e6arILf5MM8VGg+jgH6
vgh+SilTRXC/eS3o9TulwodIHx2ibBxGWaanqZFEFlsrVwaK+p5Yn/0rDgz+QXZO
ei9Mpv0tNejLjSby26qfSljktaBQMugzs2KBD+gcn4+b9SXv7JkpiyM/EYDmDSmk
m0rRQAvAIl/qAB8ced70h6VYVsb0irCRk8SzueeLOIg5Pyh3p+c6gwnFMOXYrU8/
Hnu0o0xtAUccwueboD/iVciIS8dfD7HhzoC5E6ynNxMfWYqYX7Gm31Un/vzkMNCP
G5UJq6I9mAFNKYYK+AwJC0KRAJ1tyrn1h4laP7+Lbwo9GcDzU4FkEttqPdN1nA0K
DaZZzyRsyN6ETnnVOPKtHYHWCxb2fZY1ydkAXkllYA8rz5VXkCXU8m4IJi9UhNah
GKSYD7xFKxae/rGHB6AsZDnMUgzd1uyutvzA3re4HBiRJYIlr2N1jzx6SCZnm1xo
r7Fw0fUoAEGzJhBIOCxhIMdbi+L695kGhOGfhVCitp2Cql5XNLebsqa2x2D84R5f
OeU7yyqryaLfaXg97itp8OrLcJpXka3k6ql/btVZmHFvT//ctelmZyoerPOlDEWi
KrTil2/ACNUHEhb35YLUrV4V1+KeBeoZvpYRAX3ONaHw2l7C4tTtUud8NVyhkHhJ
HTgvnmXTdanuJCeYBmr4SDpUgmQcB/i8IpQMMDWiA73Iyg7bIlNKCiCQT7ofwjAJ
HGjHOf3cXcMCyvuOw+tJY/z9RbhAsOoFXz5guwOpLocIZGMyHWGmaYtqVf9no6O4
H3VOu2jS9u4BEizZotvoUBLpx475JPX5t8q/KzxyebOXghJnCNBNeXNqs3FGVuzY
k0vprEjrNio2iIxmxOq3ynl4m7O7HkiznL/tO64HLCtMfCHuTS9iSyquAb4WVQT7
XvXp7p0TVWjC0/f754Rqrxi51rJBgiHLbOTQkvKkRYBzazBjO+vThXkcIXTXiYxJ
RXA3j2S86Zi8UgstMlAud/6ml5ruPldPhNTLDwcT8kgi/yje/CznRJPwzzDPvpeV
9uXpMI1GSVbDvSkl+JH5Nd6oGaUlpnE/26pgkQ2WDd1xIBtT9pkWquMPJ1qIMvi8
b4hGZ7IQCKRB+Rr/kp8ulFmTHhzC0EGRk2ihtpDV3nNWW3QVsyEHk1uF9vGfgc85
95dPUF7lO0ARJuyFKWEqufIzWp2+7gxDqWqtfSnWtkZ7aV8AoHSMfDJgIyGvoLcF
Znj8ahBQVoPHwaVdOQeL2HEM9H+W00pg09so9kVTKf9wiDY9bJwFikVFjfzW+eVP
j0XowgqQhYeRQluYt/hlt//gsAUcrG4NroL1i3VPWSan1xMYiATThVLYx4dP14Uz
5GEiHxnxf23W0zti1tvtla2BvJ070sQvm6OdNyJKk0wLCLsQSoKtnyKHtOhPC3MR
qNRf4K5COqJFFEZA+a4WrHTf6OzYayBRQsL9om/waXBPP6ufkhd1VFSyrWXOZP6S
5BKLMlQI0CZ9H3JkBzojtQI3UwhWlRsazwY3dd1iaUF1brBn1dG1/ec/OE20lXct
PYotKju/sozg9Law3j57IgeDXYjTOnrDpGtxzxbE9AjP58xKYpRTZQwYmBytT2Df
b1QUx7soQNGObEoDMlqQ7RbjPiYJQ5mgxoRMCQqHylo1w38YRhlhJlCX+LySA+Ae
j+hwaqf0nU8MbzEuRUzGIj4Dn27Ex9DqZg14JcgXLHCvmJxQUuX98kAsx/pc0VVR
jXszz8/43QKGWdsyCGyJqfq1/1thHPpMSzkU3rHmTUORS+lEXgrRNgHwN+dUyesW
9ULcG3CjUaalFA6vSLF1I80OsdTtG6Jenmj0SjUJ4RLdl60K56SKu0DibzLJub93
WjbxJw3YBywML19eTd6t5o30vbwt56Lax8my+nREuLd1/nV2jdtCRQW1B4UQnRIn
N5SD5oIs1EI58nuGOD810mEkvxN3sklEzMNWDnjaRAXTnxmIwGZxbssPsfVN4WoX
NiJcwoZwdVnHxpV4zINAx2p1ELBq3NE67OHZhtvLK7SXzfMcZnNHvN6XeUZQ2NEI
DpZylvgbp/juxSPG+rMXdNqyvVtGx1wXWkcOYPp5YIAJky2QOQu9GrLPzDny2W3t
VeFN38vLPVssO2Sm8v8Dz9bTuEtVrcN1ttpBa2/V3mK5jqRUWqWibAvY9ueqIw4R
qoN8bYLeQaIfi8rwq/tjoaMTHHRt1LSBtILHYqCIhy44uM3rGQskpNj1aILhL+bX
Nmi/DcDl0t6jljWKdaNmvXXA27KvPoE13T/NUqO3Kq7AstUSD2RzlvNDtS3E5qUx
wYFNdsFnN9/cr7xxPBGJ6IpT2VAQSnoWbYIXiGipn6slkQD436tX2BCVQCxeTpVE
DkD+HaL18/ajlum59G1w+AcJXuw7sVoG02b1EC1YKu5ULusr/m0MN9DR4lgDAlEt
QOP/fY0pEHgwoWa6azSZpFbwPYjYEIgmq6/AiiY09jO9jisPOx+xLbnobKxzwrEn
SPHvl+O9OcvqOu/sWIRTOnmeXnwzZv5nyVidoQ6B02VgSe8zrAI9FqgQtk9719g1
YvH2vMUfC+ePGg+iIQvyQM6MTSPTAIW7WTxB/RVFtkG6354SjgqpjSoLKcLLlg6h
uKim7NbcUhkFTV9a9L1lOlJiueiOzd1YUJbnpBpn1LgDFFKqsB2ol9AbgArdljVA
d797XRst3yyJ0i1vKUBKI6CE+CVmUfk/I3FLbnbVAWT+vZUUqjaSdxSdPVSeArZv
Duah5+vd/W0JipLapwzY1PkBiB6OrwX9svTiQoo6HlQ4mhZ6ZbqH9VhylOdVlCxI
OXAWyX8y2oFGNtPA81vbHtosgYmjDeq3KOG8Fh2EmYKJl6fzo6SVura+r/O/alXr
Tqazp8S7b3GnkZKq6E1LAx4keSj+ThPV3GIgrwe1WKWj0Bcj/kYObnwOH7k455jY
qPSAmNdVaOhXnPMeyNhTK0g/RecnrN9nPy53ZhhqqaKW2KM+4rbNRwqKxq6f0QR0
psNmxSbXufmNSZlwODAz0Biztj1g0eu0N76j+HPVSTOEclpK+fDIHQNmZ9xvnpTh
Ht2Lp29cFPr7924aQ+GF8N3dQwiko87W2hXvwBE5qGZyzWhRdYQEPdCoEDHayfUd
UO1pYAdzhsro/MYw7aXVFhBEiiaYn7LdmGrmHUpDtj1D8O3gPEEYoJt6vifuc1K6
ewW7oNXR9Yy5A9WE99x6TQ+4Lf31kKVu0gj9iTAWiRdRpeWW/UzYYPi23VrZdbze
ro0/VM1BRbyqIu+O8R/lUoJbB52TizlQkdDRlvBNJLrXF8BB716aWhg6JO30sq64
7hFhYSisOfnoW2Hwevdd53+6DYKLF1J2IHEkiwxnRy/s5jBmkCjAr+r3Zi37YMir
fJOKPBCRbRQufHqRXKIuGw6x9cAaAPu7IbYl42mzVk9gs4kh0bV9M9W16w95KySg
QAgea+bzj+HxoadMuhP4c492Cdz+mSO9EX/mGZQ8/I1rqlhe12Hjoq6QFO4+n8L2
0sl4LDI/RON74Hij30NBiqYOvgFhYLJUidsUsh4XA457vumjghXzjstv2AU0yi0N
5UN4sTQLZWALGX5Tiz8F5OyfPzXCxJ0+f4OD1U74mnd6GCl8g9ihEGqbCqHMjG98
CwTZhvpv37z2XccZoYPIb9wnGi5upII1dpVCtnOVNv5nRTD5DbONl+y4EyUKXZww
k6a1B72LkUB3ddWw9F3YMy9SuQJtiskhDP1tKN/A3boX2T9lTHSHZUiLyfZYtsdR
ohkZ92aYbY7Xtn3ISBgXI4yazYRD7Y2P6ilFG+NT5vdXh93GcYV5QBhrb3/pqEdB
BlCGw4F53G+kFf+qsjE3ueBm2kpR8hddCxbppm3pHg9qGTaA9jqdL0no1/LBTabk
af1e5K483Wa1UI9wDhXEQzIr+Oj9Z8yGAm5x2zMt5amm06BkXt5k+8Z3F6L/7PUG
xffXzfxf/atQt0gpsCCwGjQbtqw6qr4dJWyqD4qrZd6YRmiSJu+ZGDkOBDHXyM47
+S1t+JQ/XrLYbbOI+lpCQGbCBWNEN8RMHbx/ZITEexkur4bxTlNb5aC+Xn6ZxxU5
Xm7fo39ZzpmGxyLyh7mWhMtaQKiH0gV6fuVaadfOIk0W07rKx80+tYmJ2f9P/0H9
l3z5i2KxbnwwKSJfiHpImx0nLg+RzLafODbAsRGmoQWYXlHxFEeYuOZAjrIMn3Iv
ldZV3QtLNzn3ag9Cjphu8XHtqG5NJzfcRsnUWl+A/DgyX4QM2Fe60rynv88fdYAp
vGDSDf+44u2RHKDRuLJsQEwHjqWZEtEIqBp+rfkVGLb0RlmN8feA9R7VVEuo8F3n
J/C3e4IP9uq8Znl1aD5JFPapQG7h0FaA1Vs1qgPYYIBh6DZSg3UyC0Xky13S6Adq
as+OAPMRJI+pauF/CHi4TNC0CqJiejAks1NRyd789WzudAxEEDJDZMjYERNbtYvr
wuVRgSUfbmQjyN50XHr7gVjAIdU3ieDmvTxcKv+77g/hWpz/6cZueHQjDSFJPiDg
Hg+wJPO8ct+NX/jGJhIh2Nx0KyKGS5yUyE+I0tvyS+zxkqU6mFbabTGlCAI9WVHD
k0/Nrv6IceTk0og70TW4hAIoSUXWZB4I5zvE1hk1BJ8vWJgYJHaWzxRu5G4MTj/W
y7ahv7P6A+XQrjAHRRDsWwjOObrmp4pxNRm4CPp17/HFIQ56fZrWx0uCA8l2N23C
1Fs1czrtRRMcI2wob46no9HPRxRuz8SVxqX2C7xaX+fPoLDimaf8qfmC1KdpLP60
864Grni57HkanlZQI//IoeddiEN0CWIyOKwHOfMLZk4zIMcMyZU3tfcnonD8SCLq
8x8D1MbOip2fKlre7UqX8IzBmASCS2T3GFxfBPHHAxv94UBRemwBzYLdv+lmqHb5
UvQg7iVw2qG1XOytKjcn0R2aincgU9D+HRyNxm4BTQQuRf3ngyfeKR/dPSfyvl6E
4FF7tS9GNxSyi+7zwwpomZYMtV64tNeZgrv6pGUVFvs+/Wf8+HgsiVCp3vOPsTx4
CRCodrEYWTP2wG9a7r+zHaQxN04lvMfFAftLOhS4kA6m0iaobZaffH8Wbf02gsqo
r72i09yyOglQioWM+18rpEIW0eOzakg40H0R4y7nsTFrGgIXJsFSAC5Gv3O8vqLh
TqjBGjy/rrVZQ8X+NXxBnt5nasLfpzoSFnoDWS5/sP+sSNA1lpM4tMYamVcXVWHe
b0DbCPIB9pb3G/K8EsSy1ixrv0clLlwEpn8CSJ3qVzfs5RqV8lTpG4wdjutDEJhO
Qo+/ZkBLtobHNhiupB7YdR3TxdjXrwMLHstfIftm1ggm/cclOchevMqLnIfuApgU
TWdJ52S1N5AjrmqWZOSCXRY3JLDxs0odu1XKFsca32OUYCBWOH6tVBgjmiWnPh7E
wCte7+jYuNsK6rwLWv0jq7Aw328Y32Hthe4rwXKnWG2gOlw/9L9lYs8eMATSlvP0
yuCFiab3AMjf9ZkysEqT3SlvZDh7hIF+EucbEugRxwanqJAzXsatBQ+zjZKaUn5B
vys3oT5wdrMseRqqz0AU4fAv1NZwNgzAQvDpDKgMfE7q5ucr/wDRrMBqmfxqepzx
h4cKDmC8M0lYUlJOHI4VaUldwyQ65Ul8czpf1joYcz0uRmmdn7nEPYa207M4zxZF
Lpvr2QMxBI0ayf8LlKMxCS446bVRQSrcbaetoauraM4T9uvLEOEh36yu942A4nol
nnltfcnOsYWG+U5oQM/Irr+etom7WjktDUlAePo5uEdVK/ZWXX8ga4LWQy50r6iT
/sqZxnB49NObdQ7/t78hfzQd0faVNduPXUkkjCtVyF0/FmMVW5nwtZYP74n0sPz8
KGTtvi76nrEQfYEvglWvN5spiwNrvrq8y86CWfK9MUZSikiup1mc9FrL6qKHHZRS
8bFwxgIRMa4k6p3ZXczNpltL1BDjwN/yPThgu3QRKEQJUhRXw6q3NixGGgWm0aO4
9Ak4HCm+VZvtjOVd2EDK6osKglUyUoZ1WDU1N/s/JTkN4GXRIu8St9NrKxoeKNhK
trQh8GaxDUnGtMBOZ5AfikPxLgEn5cedzsEnwQpH5z2tYxh7WdNRZOSzkeFoku8r
EQVOaVIr2t9iepBgx8n6mMKFapnGH9qvCYSKb8EjO3ONMcc35XsAA+K5bzcpWMWI
TjB1c9GlAoQ/73aLifboe2JggkZZqbickB5zcz/c/UWu8qBrOA5tWsipp6hHNLqc
VCQbRe9F4TM3JQIZG2CDsoRcdqNEsYXhFZ8vTDVWizNfmXYLjwkrTNQiupkyQIFT
its05KERbGmKu4hDPQPpuC3mCyYvF7pnwvmNIdmJXtvkKYaVr+OQvN+Ll1ERauhH
4c+E39j/v1SEVHsgLVQiKM0mBTcAErNOTdXk/EBEuAS4idtR9JpMnR+x/GDMx3ba
RE7izGJHmbh+7IfJul92el17qJ9tt9Ms3GS0BSELz878bK6M5xijmYBxGA/HjE6R
KPE+8f7t0DSq4+VWFwDqq9gIt0hwKy95WFCCOXYeh2gYW6rUT9e+qEk2bqFyhsvt
s3igwAbcMzo/qWGBk7zp7kReAL5+R1XQU3yqjyXSHTgwh1Sjd5X++vcnLYfqDuFr
3afYMKddV4j0ZQj10lUJrqf5pL+H/CN6IOQsfqKDoeqXtlJf2NcLdiFhDBxLdQ5f
RNQ0MrTZcNMWBDsJO4WOrDh0KQQcrrDT/kK4AYmSkUPqfd1bHcj6lipOckPN59Lg
mnMctyxzfL1Sdg1/UC43EFGhyxcKvGUsVOe64GsyOSH/bp4jJfmVtng2V8nXivuj
9HQtuXLx/nsuAEIRMcpF80LLXWinyZmf0XTdZ6b6a1gvIPkRx2wJpW744nFWfjIu
O77pk2qbK4vB06LCdWFVn1TCIg+YnHxomcATx3dnfENexvVx8T7HCvSCH3HVP3I0
M3mYA7TX234OAfqhWcTo2+QfKAtG4qMixiSqzalJSECSjcGESEQOuMTBcrYG5529
QssLxNYbNX6D1yL2weU33tRgXLDfGZJZMpdlF4mxkQ/cqgj8ayAhW/81zpjYRzkm
ULLfvvyS7ayxL19O41VPTy2pugO6Pohq04Pw6zEEr5x2kPLuKeYHr6jTfeTytFns
PoBu7Cc1bI2W6HhYWOZOBs0JHqLTOqhb8G/M3f7on4zK0wD0yPt+lwKThyylHmUB
WWLZss/2bhuRPGcVhxGDEhVp9hHkBaIbQhaC5X9/IlhGIfK8wRAfuq19UMW8EmAi
XwoFQwXge3xwnMdlwpAtwj7rjQXxd4uqk8soIR6bl5neXVrVeZ7gDJHHltyfulpa
2Gupwz5qBybsipYTmhdO3c5HKcSpRx6Wjw2VAVSXB2UzIdMzySyJBKBf2yE5DI59
XwZuF3HbxsAaRXWld2g8fHhNnyDwvhFhz7AuFaa+xycDdPMwIPzmY/Bl6qqchhmv
7T9jqDzZu0XiZoZPhNUd6XZ1iLxvPXdDIoZerNKVE732GPwx6WuXG2CV+Y+HIm+y
7XH5tRh8EwDvFQuUzCOpgjWoUpN/jcvuYnOV2DkY+GbMeR8Un59eesoUo8Ap9VjS
TON5rOLn8QmZUW121kA9XOzAo2FcYuII+4xZ8f6greJXRRCrUTrjedSOyyQT+Ql+
dnY/75pu2smca8HKcfsuo2Ncx5wm01EtmCOw6MK+xexn7HKP1ueqIyF9PmRU2MJR
Ax2FRTS3DkayJL4zXfjI8eMGjDEhU3PO+vFBgvD3YYp1eRbwq66K8qGt3A68wlZ7
Kx4j5xL3fbY5oRjJjfHmBY+/qVcHesH/zGrbRWLinu8VJF3lJ8YTc+jCir1DQlvW
BVyRPs1HWRRG8cVC6naVUyVold74TyIT49kpb0t0ken54b9Pr9XeFZLLMZHFqGIc
beU9RvyOOVWA6iT32FKmk4T18KoUchOzAZxBjaD41eV/h9fFBxtrxJl1c0mYZeZ2
YITSvhFlu0kLJYSzr2e/HeQTqh2BR8tmasbpnCOzd/EJMOPAUskEEDUcQIqFHnub
AXs88OuZ+QzUhezkVjNqqhUIaoY0TV8hRkQ9+T6KwrQTzO7GDCykXDFS/Jcq8cCt
Bqp0bE0luUq0q8bhDdGFexCMcXs+xFBVGR66T13Nv06E0dv1MZ3xDo24DnWxkxkm
Z/72larFFcTKS39buFhttof2g1Ca2WZoeD2jeWGIwD84BpRqb65EENsz1VE1isiH
rGkgnFsKb+dWD2uuHHv4dcUMHxPQqmztYuDWog0A7prVaT+3OM3Wgfn3mPRPGOB4
3huGwboEJXWRFpRoeDcDvYTOPS/DFmKVHddnlaSU/QhSqS+T1Zgz1epVPm4mlkl+
Up5OiQ97O8JyAQRMuh4qf8nuYbrjP9CngFeKBXFgeMvxQ4WYWa3waCh1N0S+rM/f
LjLbhpz2AbhNy8KPfmQ7Iw/AqCF9IOX1TwMbekRD18LBFrxJoKt8+qhMBmvKjWVk
+TXRT+tJNkWrc/xMg361WMyh5id1DPA1hCmVvnZ42ew9+UZMJhqP3+nmiU6XW6Ov
vtynANixfTCGRSa/jHWecDs9sZVCAbUecHpajf6TZixQRN9/gk4fsLbbb9zUJaiH
HJqC/aOnNSNBK0keuvNq8fYIKWmdIoL19D4nI9b3FY/jm4IpV/bd3z1OVMP35F7Z
HLXsK3GpU7JMUww9tYl6h9vUzzP3JEkgCaYOj94V18dNGscC9YsANGCr+x8SIXlc
9bxSnCPw90XgziNMtGZPT4SliIxiTq5kD5J0n6BP0qG6qH+ibEx0oqXaMQ/xdrgt
p5sZglGiOMWeqLtZvuHP9SBT/ryp1s26zNHOJ01q2u12ykdoY0muRln6oIHpbU+4
AhXQo8PYjgEYlVtwj8wAPvV2WZ86hdmWDOx/4gaNIXgT9et7RpUUBFfuh7Hn3FZu
n1PXXlPnyH7MBS/cP8pOkOJH3EEvtczdMGIiLt16hpQI55GDQZh/GETPZfSnBQhy
goauzvRzmZ1YjSgk47VmWCHRj9LhAh1MRWevqcSZFGeru3U66K84c7uOMn8IIaDu
leeQHpqYkhfw2dUJDjIstd4eukn7v/a1Tr+8zV5lfxLFztZXmg3lP9bB19BjiV6h
Z6l8taXGmYi6h4iePXYIWElGZ3Ids7XsOVDekZL8oz6Kqd2ZCkaOZy7o7sNWZxbm
YIn7HyUa5OtaMqq/3Cg2Ig9o2Ncomu52DXHepQnSQPkQv85RtN2x9DFK0McO9/n3
PHPcWO/Ke3jSJNRT8Jj//BT3T8r6U9UveTrYY4uyOFq8t/h8PZftNrhRVYBFkY23
yfCG4OC7zYfWnPFF8oPBnOIe0X8q6io/TDP6SraM23wD9+8QP8CEKR7IeP4mAmcE
L6uwKPVol2Y/t51U/mI3/WwGIpb0fsf+N2mTGuo4OIR52+gTxRLf8Q7LwcB/6QwI
FWolbe7I+T5hspsbmJXBMZdgnHKGcc6Tp6r0VKKPu1BF0qQSLy+cCjTsMpjENlSO
i3nb69yS0S1Cg4QQeudon6GhNeS+RHZRvgJtaYIZyQSTzDUQ0EaCMF7pNU5rOoA/
uW8CI3YAnP52gglzezbf8TNyfUsCi1/SSsjZI+wgEsJ94GS3H/KzEQIvW+48RiVP
gddoDqUJcAiJEUWyzjo+aAhdbB/5ZDQcTdl4308IVvEEND4vmlPAlG+xSMxLUOrp
aMOiaT+AXVMAAhGZM49t9/9XC0RLfa/GX5oqQGvZR+O0mrLQ0R5LyHVuYiY5l5oo
zCUfDHfCs/FPiAD0KjpIW8Hf8SgjdVv9KccFknUmVcCypOG/8xpR/Rgzq5hXQW0k
MS5He4V5ytaMgc6tlweB1LEm+s4eahhrGezeodc6hTyA+oGlobyHsbmvSmuwtD2u
1qP4bKEYP1wctKxDct528H+lb/vNq4bN74ZImQLrshHMkyCY3lVzypf9QKweYBjg
3gPxxn451UfkUiDVXmJPE18KueVkQrXD0DbdGgYENAzz026rSg0fK1Ra58KX/FaV
E8AWlsQguSKyQ9tAXUTl+ltjoS0t5DhDxM3SvT6C+TohqMuZK7jsfax2dkVgTpiF
ge96CzU6c9KhwAvUrhusBmvl/9N6giUSuq/yUDeu1JPmD80IXW8UMZ+KJisABvF3
S/C66rPASFf+332H0A/X8hY5Da1Yo2P/8TFnBIj1VMYnWzoCtU5uZVM1C13jivvj
hHT5Vn6R87TZrv0JorxN9xTSb4+SwpEWZyfhCgl2Ly9rHLnqbewXqbuUX7pyiysp
dzFE9e664RAu/ot0SlJ6MMi2bOyJmJ4V2ux9WwMt1jnvCEFiG+Tw6zMAPnyxGi/J
dQBViAXigF1dHKceL+KAwVO9ouSvWYGNzizKUfi0ZuD0KdQJ+8P97GzrQD4gkF+p
aRai00+uyM9D0D8WpdG0v0fMExOZt/n1ZcRKEFnhIl5gpuTJTISZUqr5fzbsCTQZ
wxU1iQbG12xNQyi+7bDwJ7Y1D6XzGZ87zZCivHsQFa5iSP4Rhc3vmHjVi23MuyoT
aWnOUVDDw5KcSguU6pdPpaZ6uUYAQF/Pwui7f6qd4nSzBrKImyu/uV/XzJZMtOcy
+Fza528o/sZIg4KaBlJMXpP5nUm7aPr0lEVu2Poz4udKP1pEgPfNXYXpfjG6MFw0
dvtS43yElhXT8+EAl3Teoh9RrdeSvwNkabEBYF3XfVbxhngwasAXcyFldRjNh1C8
gxKsSqK1JKtRB8rmzWTvzVCMJBxM9ipK+7VawIcBT/ZHA5PBcQ/9CyfS9V4WPx+A
GPluR07ndWoIna/GOq7bu7CFjeyiW+/P5UZJEEY6v2C+DkG1DrQizEn3wzCo5eQE
vjZG7XZfrBCSSebmhqm53mvsQ4cxZ5EZcBDNJmgjwah7rHL0WAe6iL0XXeERJAXs
pApc75iNRrF8XaCQPWQrSoxkmKRnR6yoVvcJpfYx1MOzgozikbedBz/p+wySF2F0
GtAlup3EqCktle3gaggkLUioIjlBOnrz7aOSdAJT6ve8OQHTmqaflDn6l0esZVKy
kdVNadoN0kYiXTA2r/snkk8yIBeAGJmU67/jNTFBxYUzNC5m/GUfEsVf/cXiHYXW
SXzFgVahyFZoK5RFuJtxDMSLXW51FkkDI+gmzH1P4zGjzVdogZH1ksjx0yR3QVTN
2JoX4z2pX+1C20G9+W5YK6+oIumUWrefwQTRWiq5EiSgREKT8v4W00JNJUwNZOdM
mAsxKjDzv94zWFmDmzb7ira1G72nVUqUqbhGUyk9gfv1YyZ/LQNPG1A/qzDUNXiO
YSUlpAHFiDfEons01venY2fka8BRTOTI5elS9hi9biE/jDp1zQgvRvdaobRacNu6
QYJZS5sSjPCVXf60h9KbKkE01u5TfTHFFKQZzGJ3TcAvt8CKCM7nmmyM5QJGXBhm
YufBRARWpoxf6MSu84T3NoAE3ApslY2gElF46ahnpv20A3ddxoEs+q+bjvHXNN4b
OF+DtpRKFj4BMscZtAnuUuNEIMrILBpQcCpTe9bvvM3N50dRLvLfvq4djMsRAZNP
Mg9rSMFBzSof+KkpamD3GC3rv+Z5WUuTcNDUttGU5RfimRyPYhQHYkblE30OIN0l
c3jOizRzbAtRbUqkScup4MQT1jRCzNsliAt7qw+9N+9zndB1/Hf8n9VsNZl2XklN
jYiVw8J38JRcm9AVA1fGC0nO2ipTbBrfabPbUXGhIHaDHTOjrVJSrqQ6xLPVprz/
aS466eL0JBkuK5LxNukLu+yG4SyzJlxhXpiXUOaj//cM8rM9qN8/SQtD+796OCH6
yJgUL6SG0RKMj6ErmBZRKeZUkEj3i+4k/4waeoPlUdYQUmq1ljxdGXmx62/3HszV
x0kFMr4PaoaRSzy5uGYi5z4X2WCewqKAh3PFpgI9AS0XyJIetVyTIsUp0jGxl0nb
NBxXzVR725GcPYxaTG/eICCGdi8VxqbY3Ak4GqqdFTJUBHgSJ1cBcCQpHgO9+wCm
wgOmW+ju2w72jZ1Ndjc+OOorV3F89bYZSj+iIz9jW+L96COkyaKSUEp6nASaKwoJ
SkWRJ0YN+qba1umXdfzAnv+/CsUYoizpGCYlf5MpyQdNIXt11kQU/+c9qNnF4czi
8dpjKIRTn8chmK50TVXx8uuvzZX88HED5V8ADdOtvbyQbRowzPcpU0PqvCjaz83V
QVKpyFHH2Jyh622tVPU1XX0HphBj9wHsO/kFstOInC8oFmVFnqZuCoTf/Jwd6BM9
9YSwrsasNdxmrFGaed4fxz+pwAb/QexH3rqrnT1SQ/pi1xkIWLPzFvNyDfN36ihp
pGJ9PjWQIfRfpIE/zXt0i4UTFsYrRXr+6RiJ+v2/1xKJVsvn/TL8jvFX9f8kpGTL
GZDiWTI8Sesq588L+iJZHc/khtMOnLZ7Mc0m4DAbtcnRAU9itr4J+gGaS0lvOsnn
mk4mCE7uEBiOGWtuo8k+WjZhIfDGsnuoOhrK9pRhXBP0mjW8JkAPTWLsmcVNmiOe
A8cUZHg4IOJzStNF8ID0j8g+YJpdFrsmL+GzKWQW4fu8FnJFOsjkldkiEqcGfnjt
Wsb7xCD83xnng+NepJcswfQfN0HadxhDKBuudTq0LbCpASFXIi4QPGfh1a9XYTMj
njT1vYJrAXb8znNZv8Yis4kTRoFj3gnAokr7nVjy99/i3yQMYt3KRKjN6BOJTFt8
x4PQ7TGdlL2o45GOE1yHm9YMfbETN3SIyL5MuRf4gHBbYVcKTgp1CXLfdaVmeTR1
CqUL4/BwYUISmxAk7Coe1iEJDiIIP6cXlQhDkGaBk2Bh+PfK4rvEABXnSAAXjAEF
Q1zZppndi7ckeOsnRxPqdPsBSonxvvcfi+b20Gv73Gr7FDFS+B3GSkb4FYZR7oiq
w/kRRHAjzMIRzgZzXBBS2SPYvC826dDMFxa9MoONCPJYeFfcTSoGzM9ojh0+v8hf
8CO7NQmr9UjBSb+sq9gbroIlbTkoTFSzGaYLankCQkLIg9c2XN0M7XJO7v4Dcwy4
z6jGmL1msPx04nmZRbD7ULO0uMEgGJ8WJSSVBydjx2aAn+t5Xrev69L3jgygg1qQ
9851gaI1JzqOMlIROipuD6xYaLuAo92MY6M+OZvVXQUL1hupky+tJFFLtg/KRS78
UIT4Zy0545znYlGV2bWuMBPGS51ArD5Ujf+gBZCGw8lRp1NU+wNpJ7faFTDF36sn
IST6o1SRhRtDu515u0R7RlcUI20bMFIE82QR2jWg2PwLwZbZNO4TQIz9Ji/Oa7z0
z1jnYNHyTdvLxm2wwcgeZDstU6Js1yiiBfBakS85GrLzfq15dnEfut8il9//rC2l
TXjkWFg0nPsZ/YxfLbyuCvYmnjI7TH9J2fnAm/REexfgb9qwZuDnF5DtY20xk9vh
gTcI6+v7NlJe4QNyVGqOnjIp2NeZOOnzo1BSN4uaGJCF1LJnBff8eV0L8+gVGREk
Vouj1GX6imOvWBjy9qhYoVKsm6P9q+I+8n/5TFW+d3x3qYJ5gU3AFihCcKsezQP2
oqTcH//uMWk3kwn9GEQ6rJlr8rjVnEWSxL9Ont36C4zu57n3AL52T4nlFLUSTBFV
gwZoZnB3fzqttzovOAf6KdD3JGBweTsI/fY3CSJaarV+kC2fMEjm89VcmosxFy0c
3jTLw+D1b+B5jxnb4NP2ktkTtPlV7mtiDHIPL9KNoIJtS8EPlshr63wpS6x0/zd/
ZObwG3VK3hbyQqTiwrGsQRehNuh3ORM4LZzbwfsdEi43nMoWQmsmTiFyKnJfv3X/
2N2TWc3HnT9M4EXdC5WqH15FIfK8P+WFLYrelMnSjceUpO1XHxjDnIJOJQ1uGyHQ
DuqDUVX1otVzVJPcKigWkQMz8J25Qze7ugVtfjKXdG9/xw1Og92pgeMtFJs42nnr
F4VjOg1V7IH8U4MZUP4jVgacaG8B4bRvwi2F8MqYWC0jkKu5ZDQ0IukZqUXiK5aF
yiLF5GIcCz4MDwfTu38FmBnUvpBMVu7aajpoD8ldvmq/n69l2FCAwOsGe3h+wCVM
vc40fNAsvSthsub0DY8H/4NZi52avYjC8PwyKkKOkesJT6zaAlwaIu+WsYsZIIck
3dNITUI9RouUGcP0rv8Z747Pe/fsV46gWaQjVE6k35Fj7FOVDj3pU9G4X85qz6JD
2npFVXimkad3XKfSA5sVRmeJ1APS96SHQ1FOQmfEadzGNAbpcRsiIEXOTo1jqNHC
+vRkFk1ql2VgCixXgH1ARQqo43/mFPyPDmmj6PWdRvOM3rW31K5TFkd6VP0rBAmo
PAl1BgyVCUYae42x/sVDDycigokbJgx01wPnB9jRGlyuDjLewvUm4i+jK81Gnbww
fNnpNSrArOqsuAGYuBfbUvjUweEKs4ri26JuovLDj77mdcBXYZcC/C17GNeC0fdM
jfBET0R6awIg2bW138SWTnDvWOzAcIzQ31QWkTQk8FMn8gFhe+3+b4WhGTT4fHqd
KLwIhiVKImBF61AqQClg1dZvQhfcYBQ0b/9hML7IMWe/kN5IAeEV8XjArCt9vLx7
/+qpWFu2YUcnNy4Ggi/WwblycCkexdtCS4nggkfntUJqL+LoqV+o18W8x2eZl12X
2nstj26wPTBN6rkNqhHX9TrNT2597QPE5ZwX9EvlKNAYgKu9wyiV3YVIysRqzveT
kP3c4umTntsfS/hv9xh5jVnYfe4dBLBVoc5x1Ks+oqodbjNHPFG58cZH6P9+0Hfm
+MMZ0FYLSanQRS4c6bAd1cbdnbieAiBKUxNQXL5BxxSVuvAQ913gMkA2ppF9Twj6
U4rIVkLfApCMsjWSQi6kNd6pb041ZJbv6GigGKIn9yU2Q9YO4xDXVHtLtZhR7RlE
imr6uyFziwvn1mFRvGgGvrafIWYtP/GWAGPidf9b/PJvc3PTaKRC7O+ZV0tcrNuN
YtoxfICySCHBpsxxU+MSsYZAQkEtTjrKc803Ri8CMZ0jvF/8xLpjb3AVUg9leBhE
AOKSt5jzlNK360h0PVny6zijoD7g2fuMsEXBVn+qjigBmVh6/2ciXN02XyBWDm39
Ax95Doeoh4Sz7OH5QRPl7GQEQR8HwobbCdIxru727/084+IGKxc/hbg6H4FsvPaJ
vXueLylZu9aasUUfaF/z+VsHHvbTjA56zzETOWeyKzRISGvgQ6caU+RRq43ZtWsK
ObYd/SaBKTn7YRPOatctyck7zbedrNN5BO4L89mZ/R+NbGI5TGUfsAdef62/ocAf
2YI/KmCMOLGSk6yQ6j+ZQxe60hgNRFA7ba83UFFFLyTXwmg6r5Ga785YNzLHKtrW
OYrA8tt4gC5zS6Lp8UHupox9JnxyL00G8jd2/tqLl4ZwPzrtndcKBJEVeGwg1N8K
Jqw5iy+l83B4AxTAG7Jq0qjqnSLuYmRzXZ4wdPzwCV+Qgs1t2I7REUQ37BKrFu4y
dM+WLKBl1NHVHVYgrrfmchpS9Rpi9Icg4ZbgDcuKFEi/Kte3TwM+c/jSCiVfVPZB
xG9O90X1eLASrNdKUJXDBk5KVtRZnPCR441+MwE5+r9r4JTArFEC1GfLygx5UPOH
Q7EF9kA6ismPNdvhIWBjxkdK9mnWPYO+4ilTqXGGNVYsxOrkGefThdgjC+VB8sc9
mjxcL/He8qpZviv6hU09JUkQvKunxTsc14E+jlxiIJxZMybwMT/bPHAb2cJXNEmB
hS8x1h6clnFEM50vdXW2/6SY49Y+JSCvdfXJ6wP7FuNbkVrwsWRcnb2NwT0Xt1cx
SpwdZc7j+Rf7/wrp7Mg1uliaUMm2X4YlQ4ICUJ7QyEIYJSA6rh2DsNqJdBUuCPVh
MS3tr684u4o9OPH1JzSIayZCDC00BiSY+cBQQEJvqdFnKsIrYF3BmyOcqdA1/yWP
PpYIJklFifSbagnMf/nqOh92we1s2QgXkze2H+SIHH65lEs6wFt6QZjPSJPo9dvN
uSE/Ls3KjUUQA7c+G+sa2Jm9DIAau58HW31K41aAkyEkSwN7OJ+ipXFAg6uXbLqO
klmFTjn3db8Vuh2PB3LV3hUXYxyoo1MdF3oukie7xTBGIjnW+NTasE1vrOi1I9SR
ilBt7K1xJs9nTiUVPoV5+27UeRJm5XXyy7r/ISQoQOctwj7eVnQ3lDOLYURyVgtk
lv7QSzEOx2HxzGI9xeBsm1EfdIRhgz/iuP/ICE48TZC/b+uPhS39M/cPqRPzO1AL
bKhSLwfDL6sPBKEtyueRInjWkQzbGRwYbXfdjIutHqqp7jTtlh6rxk9TwSSJmEMl
JFEs6iaRSrYs4cqBJwgd4JznlsKczV3YCKi1zkF/EAM+omWmnlpRP4eQGBDsIEz2
wTxhdZ5MpbaqWOzfheEAyYq8zaChKumMAc2Y/4ee/KEoYdmkCnJCFHtK0hkutybW
cxeHSdJ6Vepe23YdiHU2XvNgvHYOjaelBK8x9XsG8Jl6GRsAMaJ5LlVrmvvea6MZ
BsEoQdrFny8/uHOOCaCCjJmAtxuxQte0oCbGH+rJbxR6hqtL3eSSHhNp/7KEGRdC
IKUkjpT26GoS+uD7CpCh3H3mCOVJGphv88jllptSjSI8J2QmEIXVbiwVHKgXg+TN
Bg6H7AiuHtCu2nmzFglTSBevHDF9pB/K/p7qzTc60A/BHjIT4MBSNVHH4MaPPY1M
qodpcsAKF2BEpkrKfQ7zRtrZ95x35lrYnTXWFFuOlGQPBuwEGtzFGkBdztkkQvGU
7DYDicTYv6+da4RySTcrtOXKT+w52cAxOu3jQfVoqo/PeweF6W+k+WMMMHlEiPGw
doqjv1wbVkBrrM8MjBy5WwIjFXCx0rmVjdrroaHeKixE+1hcNKp2QTnLvbAsuA7Z
be32P8Yf+TuDy7Pq9gklHujjPTFviLo1Y7MGDoAw2zclscQyjy5EHqWcwsWn4mCr
Fl/0wfWVokFMN1sVJjO8qnbSED/jRspmCFORX+EG3qBdwI8duEALBwHW50i3LViP
xyGU2w5DBOun/gMSagOeB23gVToanJGIRYCXpru/Dl0N6mJ5QzIRXYj/yG4/56Fl
PD9o10kWVX2JNsrVr7CRVDwzn9XxFQde7dS+0nArH/7RsqZKNCgd1Vvh2XxXqu1M
0BT11T+rEQjKdXIjIMovcAsUGZJMMGhZivXjjOg8Cc8gCR3BeqUYAfYzhVwgeWiw
5qFN0b2CxVw/JbRa2Y8dMoTw/iv62GeGgPpueS+BgB9xcmOU7Ruc+X28RkhF6efs
93QcvufMG2/3ukd1gkLDA4IYp/2+HHzcBkULQiI9ue3mQAcEUrgrzJabZMUyw4X5
uma7wHiab359UjbbId6B4DhSrKoKLbIv4d8U9+6JVtT8vnh7n1eHmktXz6q5NlXq
XLKahv+hfv5qpBLvfCktYgdM9FgXW+a/Nu8r6mV2Yorxl89ARA9Erd39APAyjOZx
iLVKWo8Gw7zXe+QcKmj+02atmarHgkMW93vkoX32qkTfUexOXob0Mb9VxZk2laqE
w7GgTgW6E7RWStDaMcc7OUTW3lCD41CNloNgjQ1xfeKMQFMc9x3OJxo747JZzYSZ
G5S4q/WZlpD9Pw5Rirbs1BVLR6Q7VPKPHX/Pfm70koI2QR++9+gkzuKtk5qOWmSv
K16kJDL1YfTj/AVr6BVa0oqgtMlkCZlYiALH8Uq2+Y3XZdOypwXzZ8JnOoKjGeIl
UFcJdVtAUxedV/RdjAeI2govdd6i0ZizG8YMb+GA17lEOOfnAGjnBNh1MgAcjHc/
cs6cgv363nR0FtneiD78t2jcI4OplSDK5dUfJXApS6kQF7X+vP5qtWSpo8n0oHXj
tQ7SnfMjCsmR1o+QaR9RZDYxHC6EHfjE2Lub+ewrR3RckURXtjhxxUwGkGWaSd3h
XxxRYFKvlT/ELRlx1uBkPSxC0aVze4H1/9soos97ru9x+Yj9MYlX9LLYQB4nofcQ
GvvzeBgLtsWi+BMSWfDtBkiSSP+pXDtm2aSw1Rd6FpRJCejPCFblwUe5NTBhiI4I
Tdwlb5A+k7alSIjWhhh5s2j1uXot1uB7/MIdmQ2q9uLwLIKA55G1bUUg3e3erFkp
dlmQZRG7KooMNyPaTxzs1gETFEX9O9bXL1oL2fZ0CwlPEakugFiHOVtjub7mUUoc
t0aEJtLvglWUo4Lp2Bn78Ym39GodaCD61dlmWMxee93sRnZ27BwswpRLQteFq3/x
NPQFa8mbRpURFT5D4mXVMi9cEgDaC7vzNIHS556Cytjsp7cuG3+1y+p7RH0RCA75
ZE0Kmpw3gHa3yIuND79lXSoOv1lfJ7BdmJXBhYJzNV2YiSpWN6oolUFAdyhc2CRp
tR9qol0R0Bp9mNC3TsFXF483bMMnryFP6Dkw2OD9VtBY3QZl+WQMP1K0gPX1URN4
OVsDlQy2a5sj1xPaogmxoSxItMamCYg/W5exgSRxGjbx9zw+MpEfsBLaaNXeBW9M
rCpHCLG3Q78PbFhzI1ksIa8EcHbifJy1P1RfcFHaFJRfWtgS89MZf0siRcjNlCnA
m7SjNcLU3oXFBLhhHrLq4Dr2k2cmBGGvie2J2Fx6GbW0w9uKiHHvBxQSJnGZVwh6
5VRMSmfZHVxWNLtmTFxoS3/JXACiFTTv+UH1K06tol7UsWSpWe3rVxyeqTiIDrVM
gqGcX7U6L2quBDUvAhwlDZeafjd7VwDycmjaZAtgmBVDekSk22DVaxY3HquVOD4p
xYl3mER8J+0MmeUAQiXxRecSGMom9LaC7oX4LMm6143ENSdlONJ7uEJgE5ZuwiCG
0qfXwLJxJUb2P2xBXe5TaSDDLlWz96dh/2ofQ6s44h0ygzX3oFrIjcTngZOg5PVc
h86sxm/Dm8YVns8eOL76aJZzy7bRimyCBuksOCdr6PVPZjdTRYpfal+V2yvkhX+n
Yh2n/9dIiuQTdM91ybQKgOsjPsrdhDtMX+TYv81uewbiXHtpP7rvq11lns5dOeLa
bFOkoGAunxurca3o0tNPWfsUKANtK5hniA8Ic8H2pB1pMUTI/wNUfLNzdP+DaKMW
XVF+HjggGGVmMfsl02e5E5SfkYuyk4bxOw7jVOr/YxHff7onmvVQJFS9AC4oHCld
Ce3uoqLUdCzsf5MVdQUZTEICOyc3ss8R/fhFUFEUcHXQyBH/BkbI0ucWSlUEdJgx
VYXVWdbqKPh1i66yprc9csuk+iDXk37om+sR+9KxP8WiJcQ08z4vlqy9ySXUO3Q8
9JP8cFAVIMPAEM0sYCqsxS2kVh5S2BOe5UERxaHVGdUV+zQioxylJ5eOIK1rNsLY
H1HiZV4Vjpdduj/BETMgffn/TLBDqxxR6feo+9EGeeTzTr+xe4GPSU4zWfdkgMJA
y5wyjRMHFU4Z17G+H2GNuRakwX2Nm3ru1wUJm2v6TIegL6Nf7nqJbGHHNyHkIlpd
mlDZ/FDn2DZtBqqnCqM9n2grlXoQxahxmmKCEYjwhlGTtvg/LlwgMdydqH8bWnjU
VciZQTqMQAo7SujTeD2pJrz8sh6Ek0+WrBSD1usSVCzMFkySe5sgrXqD4z1+ndnO
/nnftXa9Wo3b4jG4ximHyMVhzv1q2OkwrKoHeMypeDDQLlAk0ynkDzRcL9NtQ/qF
i2Y80o0x+JF1MbhlXePuuBM3i9T5s/KF3Q1BuF7oZjOjdb0HUTiBGkUOV0qKq25d
LPX3/pcjVCddDoIsYzLnP4uifzpY0yjGnn9WV2aA8u4IwRxO3AhXbazqF5aH+iNI
NrCEDfMSenIrTJ7mAbUlY8r0bLkIVEocVipBIhdlEEsJoIGmMZhxYkTNqZLBrpLE
wl4EaPYtSG8zakHmaHJKZmI6/R6IRn1Eismi+9jEjZcgbSfRe4FBkcyqHvakfDfX
8D8qk4NpqLatiUQJfswH0TqoePD88ogs1XGr1AVel+Y7dAOCy4BZ19r0YenzAflN
HZ4mksKxT71nB5xZOi0U0rqKnj9z0ClW7/P0REpf84lynudAo2+oAaJmPTzlUE2f
7JfwiYzz9O2a//G3JUXov1cS0oUKWailDbzkd6+nbUu5nlYP1CagJmyi1RXd9Tkq
Ozrxsig5C18I7gjqQ4lyAUkAzP8Wyfff91Bf7YelHZNAsHs0+LEnfXTOwtMf34LI
z0HTjmFq9PNT07XYI5Kt4XtKwpJIPipipGF/R/DWU46024TxLPfTHt4BYLAa/7J2
TwhV//SQ+ZaY9SsSblMO+GRfttMcpevNKPOaZrVZsGQfBcc6Y0z5KR2oCqVNOyxn
rQKmi9ar4TW9Ybl9RxhJqeVnX+STXGIukKrOw0+0DLhM2lm2QLPa2ejUNyzV2VbG
OUThiR7jH1mtrfIxnlWTG9LBeQXO02jFNXL4c1a3oYYnwQFSJZj0mKATQsDRx2VE
icibWQoNXjGzJtLMeuGI8ymvByRmFgc31uO09cnBzbOkuDUXu1nOA6X86eYrEX+Q
pqMgw4uTMOFFbsR+dk7qtVdEb/ers21BPYpuhYRMRxpGcWrKBXzAzwutENixXgLP
aB2lKgNcOgB3xbU1PQlJqwX+frj5qZjzRHYPUW+AZL2DyYyI3e2gq79pQDnpGEQ3
bKXO5H1ha4wpx1mF2BHpWBHcYbP1L2kBL+Eb1be1xWNiSseA0XkgHAI5syyvPjq2
rNRO1vpeTnQy67WdhlHcs58kHY4bAYSKe1Pk2sl7oVgEMDEJou4lsDg37EYTpFOv
USJd0qlmYHfY3pfaa9kfLSW74Z3REZaHMaZaZHSq3BWZVhMHNucxmD04LyJRj3+1
4fhzf86UjNgEd+BclaU5sVdQyMbMFdUIEnUdfV2jyCc8oNlDlEpJzuEVX7Xm+MUT
HJEHffIhjirxGqmtY1Kv4xZQjbwNvF1r8f4WLHgrP9J0Zmkcc/CcE8HFGWU1Jt9J
kI2cT8/efLvzgprVajfELaKDA1elWy6BXi8dTHOy4f6OrXz1idwUTneyHUS04kE3
IUFlkTZ1AJ/tBy9i2z/ObWZedGBKjkL9G9xISaU3EXwQJscueCj3oBcGuE71Y+QF
xgFkBAnw40UdLwsOlqcjN5CPIXhHhTdDd+1Bpo63aL1dHSPm1CfMYSvdbSC3sNMw
b+pZmoKf5i2KiGD1WKdxV1zjq1QF747OIi78djdxd60foMCxm0AG2Csc0Fh2yejp
ufkgVHszdP0vAuhMhAQFQa8HHs9Nt4RGuXE0RvKQa7xkUp6HPR2GJAC1u/2r6i4p
bPpWNsrqHlWlhxlBw3KB/98IqP9Ha9qhXEOuv9fcpCoGHdVRcNfv4WUFETfTvqvb
p9ovmMePhc4OWlCulGHSVzHfLB/shii0pzLvvv/6zj4aGlDUl+H89vf/vlSONToq
MlGiK4IQHgHdNkDWm1Y73KcC8nyDLfqEJrxPgf2Z4FM/MvjpWF1fY/L5qWXmnTd9
yrWR88q/UgfmitKKLLZmCD8oaiQjbrCepgoIiW1VJ6qrv/jpe0A+RabBUSvTTm3c
sJDV4agNFrlYnAURpKObhNVym+8PpYKuMtY5ySIes/u+J0NQLUHoBoHaNRVHCbBv
RLk6+uc1NuPWrI7+yRjfl0GS/p5FVkySZTyRXznsjjCpFLE2zbqngvnPgEZQTpTy
dolCjUtUGoiqpco5NHJU9lgiW20hseCmF43kE0NkLW3tVSma3ifs52qaie7/wKf4
XFFYZOl1sbl7pVb9E0kVRfSKHUG0gCVx5A2CE+PQ+uo0Trjq7GIp2pnR+Uzedn0n
+7iIqw6UXIgt8jRC3SDtH0ZvYDwovOgVQ2OwjZI98zWlQgDKyV/UjOVHINIiM1Qr
fxkUrmv0H/hSTD6zABDLiXNxaRoCYRH9P/wJkpt7UUrCCYMinv8MORpM9GGABWSq
fBgo1OaevMUJnO2yZ+YU5RFSKoCyoAwYLIogNMKnidpgVolCpL2bSYVEUTNbgzZL
kUZtVv91GXgOvoWMkuss0N9y1ZHskkwD9JdUxejBPiMMCpSEAMGgF1iaLUCKg/qg
gLVySU+GnOSQIDiqckkCBmmsFZml3m5w+cDNzr2D66uuBSjLeLoXnIehUEedHOO1
+ruMXxPL+LMAE3DAwVSqYhzn750SV6gy2D/tSZsnRMiElRjk4yi0SawaKTZ8WjPS
1YH8S99rg5Ew1XE/1vXDMJRsdLjBv6Jas3CrbsLWtoKacjkBfLU61QLbqWWBNcZf
VNQ4nKALCRC8E52DNKEBOIlYjANOzgcN+vBOSeClc4vUh6cbeYt3mEOjMrlSW1Z4
4gOJ0R5/MEAVGfVeEqONbmBLHVP2Iu9ybF4BvhV9r4HwGbGygX6d6SOrLhvbEwVV
KcVy/5qUVCwWP54f7QkZhRoH03cg1FAnaEU5QkHRABej2MQWjO865HoTozIuZozI
FpMs2zV18PpWZMiA0o29+LzOMIVpQrrkz7kPvTBmGKGD7IYBQKNI9LthTi5mAef8
2qnnrlCc5+wViO1r4smvtSN28C7oRp8f8/tq9IZvRyuRUtsw33A0q1qjixUO56pj
V+zfrHTcNCTrOGD50/FCjIyDcflgbWXpFUdVsGcNDbmHUepqqN+1B20PgNGLGXdK
fWOvp8rhElAfEOTZNdj8lSn1McErqfCNmFIqo+Y9SdVrc1NaeEjxe8k+wE0rFzDG
fVAqDYSjn8RxI9OQLRYLK3//hv+qqVNZBzrjFe3GuJWCgiopt2i41PIUQiN4ZGPl
I1wvB9lMKwxNVIZ5ftsfIVhVs7dNxukr9Frnz+ZckZC6DsVOJ9sQ/4I0cMHXnXiz
5hi2K3RZ56geNEDZ4Oe3owrvh7Dw2Y6CoUeZfbmPIy2IV+X55CKvtUdDCbKM7fB/
LpevHbSv34JHUtsJs3FjPIToPo+GCvbcTUJfp7flMJ+P9HABh+rRh4eLTXrD2vXj
aWIJ1hz24HumiBIkoSMQV0AKa/s+sfKDLLe+HWyg0WtCVQ/4gAc/i24Ff2/1No1b
wmbgIqJ7IiNTr9B2bzyIj0zFvRxCgeXTOMyle4lLNUjbepFhBa+QkSUch63T7P72
z/Bnt6GnwnKdVDrNfF1cwgDbN9BrkiX/pf+pi2T6/p5MbrblXBaqH2KOJJKudFgG
y+Oy9esWRvuLH1Um7Q3oAWC65L+vaFX1i4AYc4D4ncyHPTeAtDIty7t0w4rSnnCX
WoLhS7F8XXZ0+WdVYZ6RxjVi9E8q+9M6xCIS+4zcxuRg46CFwoGYmWB93BqFwFhR
r60R9AktK+BOwYAWpCX5cy2qYIzvr0qBJ3YFckj9KOq0nC7TANeM4kAt6nD7UKYV
2vwquu/qtZn6WTn14LfidmhvV99PyKBdkqqrqwwpkWk2TcdOJPrH4Yr9Gzjmj2Jh
GqgRfq1BJPj8oAFTHwmrP4QzOBuyJXj1qFw+rpobKSrVuf385pqWRFLcOoyX7NXl
MlBxmySQ8NENODMmalhKzeg+gdrFzMdHPix4sxogvC5qH6ZOcDCUcUh8o3zcz3jD
csa5UdRafo/VG+KSJ8c66EwFW4oH7gQMaV8PpaylM4fFt03croNSZiU7jInslLKS
pKt4w6TVIkphILq67dmDh+KQ2zJsYLB/JTtb3YVvPg7LGQVW8wYgwzXwX5aZPitn
VeFQPPmzYkVeELgtDggYhmkjkOolyI71rQOMj+QvO+LKxsVXhHAf+TYBISqBQfCx
sxRfsIaPaDY7Y53qETTp++/yQuLskegaQRAyzHY4sleXloqRSGxmZ4p2s6CL/wqb
HqKvyf5qKgSBhjnR/s8vesw3PVYJoJ/gIGxiD8XUzVsVPbGaxoNjltJBe7tuz4+f
drXy3km/DqohziR/pOWY3KNmTIrL+xCwjGLXXkmdx7qHTH+QNSIpeGHDskD0jXjh
HG1TgADjiTJCaJp6Lvc+uPfnsHc3xIpf3jh83MjBaNrjYTiztllrppKPx767tY0z
D3uybSo/8hJlUgvukFFMHeaIBMYhNRr7BbzD4gsLAhsFupYEXDwEsB/EFa2ORjxf
jIDPlmngstWUchqtAnJbg88O2nDkhJe6ulXgJc4SwVu3nxBfWDUy4AJeCIhuXAF7
T9B9TCwRV6IedRjy/HxQxDJpsipaXV3ff+vNn4Lma0QmmuWhj1kvA/Tt5dgSJKsL
Z1G8R/rGQ9a3OWW4hsK4N1VjdwX3A3ZQKHWvctfysO42F2T7rvFIDFS5lWmhxcAN
uqCDygr+SyptbbGiLhEXU0MULF5kSbatSKIuYIOr3vLTHV5PSrF+pExpcOb0tBRT
HndwIwXKLn6rAZFpiYpzd8TJ82o4iU3d1lBCyuEL8G5M7JfsKGebEhQMKog5va5o
j+RwbSQBv25hlO9iF6bRbYg8UYaukTz5zloGJVeRKkrDjmA3lOgQQSsdxozeYqwB
tnspJvMWi5RxTbErgEuCnlI+9A4I7n30PrTQTHfcoPdcxL+tXcF8WauSV5DluJ/J
Uo1DCwB71br663ybNTAeZtb0B9MFySF6fe3GuB8iAI+rPKPEv2Oj1CeaA5c4mbh+
Xv381uPrkHwzDciDIWDvouLD9FYh1Vyt/6PQGYYeHT4Vq4dVIskpZ9jBpdqZ8J6c
D7y5/uiINwa319PV1qi+lFqWZqgr/S+SHjS1s2tHNw5R0+kEAuvjR2CiQPzv+5ds
TdZ5w6XrHkrVUXwhFatls6BtdQ6KFYnUgcwgAxgEs1zfqO5PK47PwmkA/+ly1mT+
Jg72/hjDN24I8/RBN719UoX2mJCK7D0Kw9atYRlTXuGZtMQa7+u3I/yebESfzn6m
eRpj0AGiv/4xPXDvCuMNLxfmvAdc5g6813aF3K7Df/0Dh62yTREElvUy2kC2jPZL
EIJIKPxiaCM1mPIBZqWG61KTIzHGm23jcg2qRu/GNlq9jloT21l3barB/ANZxHi7
TEf4FDRytFt2CWK0NqWl5NrpzlK4UIyeV9nrA8VWbQW4fq9AF8kWochZR4X9k/QQ
nnlTJ4dnGTlQeSWqDy2BSG7fUUGp574cyLbKnUWDWclPdIZbdjR7JEH8tnsJuqhF
qge4tbgNRbLNclHn+w3lWfCKLi0XjY7/eY3g0otbsS/5CNwxAekf+DvSl8yvXkxY
7clJ5m/quKG8RfY6+NI6tptxpUAc53kv3y5Mb2OVIQzVePJKrsbEkx4U5DK41Z6r
fgwAxoJZUp9b4EBto8wRSdhmgWWnN/r7aykLnD99AYn3izfUbAtrpbTkVOW7yhDj
LME+dYLSRqAdxYfyJ5e74vHiLJdaK77m1BcBbJ97pDm7pdfIAI6P7IEhZMabQs/f
5S+2BYpbMT2qsG/zmAVgJOLPI1/Z7d4EqwzNfoqttqE3vt6Dzk43ghJqlP/EYmKn
Dz2z2Q8OFaaf3lpynVdEw3oIR1JN9oqH1phumT0JpxW5DyAFqCuQtdzBFa9NV2Nh
ARAYUStjI81c5nwZ2whCZ7wy0NEYcEZdVvIo0QfhXCDyf+32377YgBZszl3czALh
ccwmRXY7mZ6xLQNvob/53RgPfqijEEiWfgr2gc8iwVpKCaE6Nq7akCbMxYgQvS+S
k8kpebmWRYGs4pYahOSgn1gZkCfrY1NGQOZUAfqvkw8JmTjMuwDzSBsXYQFJZtJ3
QODgZRk4RvTzsYQrgKict3vZBRjfXtAtebuxe5+3IPVDU+uvWarTZH7vC5DrOYS6
3Il80KBe+E9fuMBrfcQjoFm3Ig16dNUa4HMG2Kul7ihe9T3KJ6jxa9EP5IFoNNqk
mG4NSVP0nnVJktfrKuNkvTkiF6ooaS5bspXUM5chNOP5lOIlKlwxNySG/GslG77w
TKB92RUyMqHcNjSAxk7w+Dmma+FkyJJwgzpiNKlp1ptrIchUqRgpPfCLdS8UJHAP
rMRcnDCRKLIVA4XKvlcv2E5fk4eVQDDeqC90kibJ0zDreSBkBSiTMLofETJ2qhXL
COuN33kRUD7JxHpb3Un6lfiDRmj3xpC8hR18A9in5HKL4358UUP8b3I8VeZOeQ2J
l4EUsPetzIyrhT9u44iYDJdIVZQZxn8dg7lEUW0B1kgc+5UqYZeofsg1p6N1iu+8
t1QV8i+KsrCxHjAFP7v+ABxQWPRc4ccb3U2c7yNAgCg/QZZxITx8I5h0t21xtTiO
H+3R8NadEsVZ5n8yvZ0nuqAUI10JP5oowJ8yM9tbkU2NUKUGg+WA5Z/oY6cadvfH
ubblA2qThEHm0C/9ifiCNNdukdSirwPm0bbX5ry2ag6EuPnaYU/nGwvCsLZ/eJLq
AMeJ/qSvOgmtwHEyPcBPE3SYLRYg1uqRAuAnn47/WTFkwThQkpBWudjyO/PW5NfE
dMQvBAgCNd2o9H+IiMsw7qWL6DEQS4e4+7qWnejEaL9rrU+7JZowInXunniVxK3M
gOFcxUyWF8QD79px6TRqmWzjFlFxWDFdyscEdzDLYQZxNSdB+nMSKYock6pXY8FF
jyJPLzr/MHr5IkofQ+HJWcoSszhicwOG6NKVo18WyMegHatwKFazShQerqCO94h8
H0+1zOwwXlDhwWenIhje8ThmdOW+fw62xpBYKe0aU1iZ3S6v2POa/etnFdmTlfhU
mkRIWoaPYuMEkV7UBSb8ezQbTxzQeQ7uoVZVXBzQiIF+oq5yoXTR0MHvzGoZzG1n
dfC2YKSjZ3E8oJ+WL6X7BlslJ6FaDE+H5I9CZytAQ+pub0ApS+FzPPQ+E5AwnUzN
6RxU/Z/4tglSntPWSwkLbpT0zUhZPdTPmVxDb/GwZSfxDVnJFuxt/h1otWYMjsMn
w9dhvgRhzMlpFIp+dhdCFZnWfjCZT1n1rZXEA/8UjI6lD0ADlhSyaPf6CEMjz3bN
TmJSJVrtRmz334Zzafyb60PnBEwen0qs+9fKSeL+haAqu+I+mrdU/3w/tfq8mY+u
DgnF5xXKkOfb+PwDVb37lYOw5HIGBwvKKWKNoIfNByTE/FRj82yu4iXxfyhEeHCg
6uRhyDQ3He/H15WKfDP2WfjWNcmjxM8yi1lLWOo+/Vn3QcnlL1Z90iNdOYeU1Art
mNrP7shHn5gr8KjR7wQKVw3EsMN4crCtPQut3CWe3fKEPnMIrFY+d8wz9DfVMOO+
N7nYuqwWSlQ88tTd40GhnWOMhOPE49J8Q578FwEaar5AwJY/DcsgZdaoINm/00Uj
y5wvgBbqor63eY8R985ibS0K4dnn3nTxuVHOl6zkImMbaxkiZH9e99t3L1AJ+pPu
+m0P0opoCqFfA6SG+3dkVxYB1NlDViMf5/7WUvmQRPBqWB73R67QgHSG17ckK8wS
BZ2BlqM5KG65ccLKTGSeLYIy0cpms9rCqmxWGaeJqpG0z8cTIdqBuhjcwmcEs3BF
5a3LiEvRkgc27IowFrmZmBLsJHwD11IVaLUs8rsyvgyF6LUU9Svm54AoqepTTKYs
lH6dOpdNwIvOUl2na9dT07bCsfJGiLzuewnXmDMWJVN/fp0RNBQyqDkOw3Q9O9Xl
pIKWbA4WKVTPhlyxPTwnMh+L822TfFbbZ8i/yH3vbWEFOwX5RyyUuJaVcTjpacM/
JoXBvUO9UlAQnoS6m+FtXpDHW61HVtXjXVBbl7E2xnKrZ/Uca3mBLZKPrfddbDAP
bqSO97Y3TSjzHE/S+Z94VRSsb7R4fdosW+gHAW8cD3Apu9K2YQlKbE6Q4s9RD0Hi
5oCAWzoUmF/qonCIiQGTkfle3tr/ENIMFzzFcRli5dllEmml9YJeOe5FNOTgbT7l
klsbaK6uiGNwq+9tvL/Vh5StbXsvc8v0QUMUdJnYsmw7ru6U0tOCekH5CKpgCnfF
hne2jxSc5HLVhKqZ64kkR8yCMtOcFDRutTsKk9i7HdeoLKsJS5kCaOotflxYZfdR
X2dolrNZaMtwWc7XmS8XC1BZQhsfdohRxiFqKeZKEdnR9WCGgl7LlC8rcacGMEWt
ZCD07PnpCRQ8mZLqhPz7eTpoZG3/OYIozm+Y/7ExFOZvR/J4EOj04Q6hT/ZC2dkd
XcLoYlscLrNFTFF3A6g4wPgWWMS8XJfCow6ndzY//2nupw8ATQpFNzeVIXADRBKY
nE3mQ4SYetMO/RGwcgY1my9hhSVGk/L2sKF2ynWxmYf6JTgfrsafBJumDjK10r7O
y687X4rpYQl6fzD+QWuLkXuROPH6RVkGpH7EQlygD/7KYi8M5pXeozEYlxE4yUbg
JyYl/tFD8BxoxGhBXcCmab6cTQZe4Z2m1FaywkTV8/E6a2o9OaN4TR0Ywayiblu4
xQfBUFnfrVq20BBCUDS4qyFMZ53b8at2em5dt1yVX5QZtMIqcseRgZi37bKDkcG3
g2nm2hPe7E6Ofpqis7rtvsomf1AKSZzRa7oyY0OJJp0t5YnQ3iMSKDo9hu4haTKQ
7rBQAniCIBoqbuqqlnk70AsiTCcXZncCOsEl+3KdxoEtyE0XALJ87pSnanAlVZcZ
FyRg9jJMo3Kk6LMwg6tqscuMjsHt8/r6WT2vOCcByFJKAEO6D8Cks7GLnZrZkEqu
InlYRDT83+lAcAA9kNmcVxn2H5RD2E7eL6XbsHGiiSuy4F9LhcaGZOQI4XSice/u
JcXVkuaRKZ6KPqnNNz+yTaixIt35P2uSKVirsksshYPd/9hv8O2rnUSC+sGNTeMC
ZgWiz8/6PEJEc2m9hKoWduH3Ln0ZPKnnkkdUYvwdz09HX9AvFgFAAUIEzJ9Df74e
mcN17xJQmSgtRResITdShUhody01i0BgwwTNr7qiYtaygIgEdSuvDf3BpVG4v8p+
KL05ig8u+ZkV4ustMHikPqtRpytxk2hV8WnzoMdc8NcP5jssNpycvMMf7fEYhYU5
2Gdlc5GMJA8Dq6VWvVRCy+QBQUUrz0kYcu8IKMB8RSompasTjQ0l9iqWjbDkk5ua
C45sVyYwRxTHBPWsyxohAUkI8nunKQIn5KCGZ1f75kJv5xoiLYc0JItp7qfbNQq7
6PV0dnTYHGrx3c0BjUI2lfO/A6Gjs9DTuQ4iHLAvxG1EFvNgry632dRp26XUNENp
hTHq8p8if7j0rAlEYDWI28qKr0pezIpMFuqKVZL4Cf9tSpIqKyQFqwWI/3HLWuqk
qR9wrN9JQSxApMMa1GWofTq5k9ERcip8oFKeByrM/jsPcLnh20jV75VQG1PhDSiK
TvosHMo/kBvEkR8uYeCzU46OYUyzAX2Cdq7j7rxi4Gbd2ieEBTEahc+2DBpRFfiH
H2dw1PNQYj3PSchzy+Ciqsh28RVVYXLTIkh0eTO3EN2g+j2UJ7GdUnb5TTM01rjG
oDs1lH0HmQqyQeIkWS5GOOckQIIogFlVtDIE2DsPOkN3d9NnlwNOU4DNj1T5H0n5
gLkwRYd9e8DwmRKzOzYeexfhYjh20z6ecp5mGGQEGQpod31wb2GNAEDfv0nvb2lo
boYRsn1fweX9SQyfyeo1+Ju/PRlvV2s1IFg/dLzYm1y/iQ8xSg2koRnWPgfL2Dfo
ALXqmxPvtDNG5KpNNtx7TR0OGzK9513I5b4SJB17DZfyzQE6igF5frJsYemfnCu0
lY476dmTM7b7M/+/rVDdi6cFKlIEVrLl7FtgV0kQ5Y8ZAZfrwKpFFisOatzp/qDl
mW5Eh/WAH3xE7GJQRmz+S0s6EN/TtkLKn84b9ND7Xh9IQE47/rZwcT3Ps4JwYW9r
rcYkBozuBd6ZuA8GV9gfahNO6qunxlyBxDI6f4LWvkLdMp8WkRCg9iob5MCBOK74
h49H/hWRRMGpOOHZl1WFjCsimRXYsT1IwNOXdPXvIW+e/LPXCyeVYcwyYaDbmYSF
RKcLQwo0rTTPF5MSiDGL9Ym+zS4I1QYR9/l2xyFVct1DlipraGhjqyrPppFbskBo
32M/4rzN1lsonBSQ2ukq2RX3rIRtFjWzTqdck6Qno3zyN3uxJAo7CAXVVEv9ETYx
E/2rE7ugPQItxAzYo2cDYdeNQrJgg+8DqbbMOff9KR9nUsXyBfkUlWayWFhkExEZ
E+52YDv7diPQ7r1pE9s9l1tFYHNmgXOKsbUyWvxzU5lfd8nWZwU5wZ6E0MUNiLTQ
IzRLv1Y+ygHnvynK21sOa7rC9/yPf27JYw82EOwTXm87HNLWV7YlstA0/8vaBOVn
ShuAdqvolUwNCM9q9xa3qR+v5Z668Vk3cbeU8XrXRCN7bGbz9LugKcA+HkxCIJZ0
qdqh5yck+sKcHWh7VszsSPtuPlUp3GUtYnsy2Yde+zkCGKyQpJA0UrHNj0BdaBRb
qgQa7iBBzBGwLsqvgYRyFfawj3Y3OXt7h9p+finrXhfH7q+rkuXj28ynWWIl+w1i
qdFqtd/G8N+6GN0eA/Z/U+sYJ/2nkNEfx59pq8aE6BqyGT1PemaJZrifaUjKpv2l
DD0guwskLcbcrS0a3z4BnKZy6nv7hL7ivxBkJhQqOJASZHRAnrA8PGtAziu4qJZa
//A3J0LgolMYyG2+Hp3k3zFkIMsJxq5tvLHqSxYnJxOtft3GGszYbb34B4JTCsF2
+xvjJfR3c7vofjK9twjFR8Py4fhMh3k5R9pGr961NRWMky+WgOVYPal1/qVzUfKV
+e0MkqLfctqSCYg9XIBaGs3zIbKKkd2Sg5Vw5ZT4czU8IqJT35PJi59uMWix9872
N5nzrGhGoL/ZuFmxgPrSbwwFTtiYPUU5h9w42Vi8fwrRTbXgnroHjAqdAg8lD2oO
rlszNSFJQYbfeNFfHZKCuXxIdUHpC5C0yLDWrGb/pJ44g72dittC1Sfhv/0/q08D
ndAgTbuKZC1sfMrsyWD9BQE1n/UMDgCYvpkrJlCVHtnBw0u+LK41A6M8sCE8DHjH
5SWTqGGHPBDMsQ2J+hf39+l1xDTMPRu/aRWXKybO35M9sqKYrorcBSw7Jc/5V77y
11GnPXSii0mNDGoI6mPQtSKFIF8X+BFhxghqa9o6pMJIdj6AfpvJ35pDjhyomdrV
cD8FPcuksQrmfrfO0w4doPtBzaoRaJnPQfBU8RbiMHZwx1Lv5BwL5mSO6xIDMkp+
oMpfRLrnm6u4rZw+IZtGL+MnbfU2FWw487sTLQgPHzwSHml7JXaoWsRCU/G/x8z7
nm7+tjNqixw6Q6q/HGsziIKS90UbinuTbq2cUBRr0YwEtX8MHklXaISsXa4qMKZS
gs3QmqqvwgoE3ziqhbMA6IsoLdIQ0nE5Gy8dwT2f1iIq9ywl/DUTQrAXbM98CjjT
rlhxcnxwLVsQo+6gqp0MV+JaAW9m6R6Ibamk18biy0Q4bZYxr4v3Ol/yrM7Jtv9S
wk7N7vIjzhvYw3Hlcn80gtkwAJvQVlJiSCHoO2BJFc0im8eUiaQvsXcZxPZwkk7V
pTTTHhCV8hzreCAcMMKgI1oHvMSJ++6udwe5rcDhQ49zPMHqoaHXXsob+2tb04C+
g2ce8ZwNF58UKrmM7/oRPXJDdnK4pMY2D83bgkqEiURr4R7PYzwHATC34TzezVmP
aEOlLxcWka8Sw58DFiwtc07ZC/j23WZ2wPCNa+nHIvXh5ApyAW8QinM4c56kbBAt
OoTKkCdvaRHqvWjTk2cyljDuC9y7uk1WZ9kdrvJwMMjyCgyRzoO1RpkryIa5+1pe
7XF1LfIKKjEJl6pbW0K/IVfpQTK+HWkt38SCXHnB0+bjOMs8rwKc38OLf7r6GZHA
ry8I3peOh+BAosubgsCOJtMoHIHehgpTg1fr1Gh+wg2q/e/pi3beE4duAPY9lEig
EJMpQRis5mDY7MhhCGJoJPhJv3xc3QBopMrCU9EtLwDIKAGEyWs/kX+zhcUdg8h2
SYrolEPitB0nLZn61kGhBpszqbG58r2ErH3yLOeMdke/XLWRp9rnHhoYhwEjceEs
rPJkpT9WcBePX6Lc1W6tJ+XgrtPYtgs2y1/Jv4arTOg104ZpKuQGeKrFu/vlezLi
7p1/vhyr7T2sAAuJkN6L+rPp/cjgJQPc2Qa+x5kznUv6mynt2K5mfVF/QFsPCK7C
wLmgGy8PCNuG/inyfOCnHLbtQBUztGSMwGi2lt09onK5lzCZXBlcpmcz84BicdFb
/ek7tEWHn8RvVWN4rR0KBPFvRiYdFyA/2GY9fjE/HXEtPFTwVOzl1PXwTgWngKtL
Zr0kH8PbxZ50xh2uWS+Ze0/HwIWGiJNHMgIDByKKmoejujhU8BHhtOwi+MdSkWGc
RksOBR87c6TWIFyVId3ZMQSd3SogESUB9h+RfzjxORl9wcQhUtcSm2KEoAqwrXOH
klvlI5Ox3U/FSZXqovW5yV7RZxRZoOIYqS9SjiXFsneBTPT7CIi5lFzdxBZxPV4W
Q5BweMth6Ws8Eux89Pvg7qItxAOGjg1hP9KBvUt7bgkMnxwKlOmIIk2K5UT/7YxN
5d1IFavILR8KYqj5C9f45DrXXbTfsIwZOQBLBbMiNGi11xFdz0+GJyGdRBI7Vmqb
i/5ZTGLSDdY+RdMDPkrWpB0EFbiVu35mRclQqQiex6fsPlsPoPIEUYhwenKf7I3W
PUeKK4tBKWCTxxX2lkfh+/i9RYIAkg70Gnq7ZaO3TOmPZga2aciy1wywPspm6jX+
p4JJXyB4P3n/7lG+EnjW77wo+zR6YvqjbFqV16ng8Rc0NSjjVbTVuN9SAUqcWOuC
SnhhM8lPhV69H8tmD+5ZZ5L8jIJQOijuFOWSvO1TizhI6pO0YNtIFlJvdzvqBd99
S6CQQLd7cfSkKxkOrhefkdycJHlUPfuWXYRABboWBIwV33NUVpORswh+ulge1GdF
N1yH6MdBRS8nyoiBHXwiwBv91CDpDMurjUlIPQhkkO6zJite2zkoN0lnDTr4V7V+
jvogzjN/Zpn92up8LIwtWqY1a48YkWfmANxut+rTEg7epA/uKFbSQVTdmkH82W90
SATHABQ+NB+2ibhioyLvDTd2GplmX33JDq7og2H32H6n4BRVWlK2U9ct6iyTshd2
hiL1baoFs5r4Om9uQw/HECpgjK3A7sq6rPMFWvc5ki3qYdagAB+f7gFuESkGG0q3
HYlLG2hped2ttM/7A9XseJfZRJ49CnMzNr+Ust+lBPCoG9OlaF9Sul9DftBfTGJi
7PixSEm5Di7J84ffKUzEwXdM+p+/MZTWu3dK32D6l5DWguUP4SUszUzMmoJIK9m3
RKkgN+pUdzcTD+sTBwq5kzxB09QkhG7viDW/orbOF4cJwn5CyLQs/y4pEMtgyyBu
9o0RzdXcwVMv7eeiUwB1bHsmPOMgYjhfP1NuF5fmcdZYVIg9Rk8ysJx8qJcVsVz5
xzPZhcAVO/bhOJAQgL89OzobKzmSicWqFE/f3np5hJa2Xc2eldzoREOL1lAV4joQ
x1e4kP832ShFVKIow+d3g9m7ypInjdBkpY51ubiEKHO/nwIuBljxPYJbxUr2MBAR
9x+8El8IIVM0oMLoZJRzkTUxE+1U5P08QJL8Uba2PSIKB/15bVhGBWmAgjrXyKxr
VN1Ax8PliG11RgHyT0I1Mp6f5dA7m2ZFwUFmR6RXB3rfH5tB0ThwlyMvEaZokic7
fyAji2O3LXXUqIaVEereFF/P1UCvtax6opAQ5uPZFcCWJAiV0GxQOrJqDAlgQ+Sn
n5DBdyvLX0mXYIs5CgcEyOeli/CNU68PgvA7hUZYFKZ8q5NgUhNgTekM1OOeTt3s
50K1bdeZL8Xc036IO/h2HL+kPQW2HrGGf7o7w5ivqLSClcvy/p/C/8dXmPfr/Fnd
Xip6sXW6y8SqMnC93G4ttqJWHKrk+SRTNejdwjX7AZG1EQAe2UCzIJ2M+L1rda3h
SmBi7FsUUiRZssfdRPZ6IreyP6ccpQMxUAbE5nRvMF8ODZbeGdWLiMvDWLU69Oeu
7mTvIKuDt8UzaQGwW/dsPnYEUHh9GfWOpXLCLp6fuyUY1k8cEBzUJQhbCtUeW0gE
Y18Wu8rbFkrnc3gymwzsxuEn/No3vHtmvZi7r42Vkd4h0gHyvBNR3jotI9Z2AG2w
4W3EZauR7xrpzu5YJoKQXTlL+N1zJgytMiIFq9sN+5Jm72IgWiepM6Q6HDeVJ2ze
GPnTL/56BDPeKK/XTcuwKUZkFohfdal/YxMbyVDWcJthR95o5P5taQpZ+RYp7QGr
U8NM/GfyagnjXEkX2cuwP1T9XDRvG7fOaMpJeTt99tOaIq7NAflBdUlJJg//dEif
vW7342OKkmyv1yYr1tp04havG/j8WI51EnRkqdZ93VUlm/fdF0aDNp2CsptTHPFV
oDLkeDfR0P2do7uSCHQh8QfZyPWjE8vDExYErB1Q3stqAdR9QTF/7Znesg94UBry
ddvEL1Gb4+5zPxhkl+ouB75A/D+5XiPOVuN2xA6BHm8DD6DlILZu4kw3zvjJAqgi
dqGk5WpY3yh74tV10SCniwHXv9ESMeumBRtnaKqNk+cYQUIHGeC6gTzMRc0xiUx1
N2Z7SCdBqc7beYShDL/9prTyXLF18uVgy3faV1BeX+k2ojO5+mR2GL1bEkGE/8xS
zqKF+Hw3AT4gD6Sp8HVGIMhLveHtBJeL6e5VWMBjgbCd2ny+v5LNlSVppttYfOyT
eSBw6Bb778NxXBY4cphKqPX4ri9b8YJFlweny9VwOtEuekekgikz9ahChhflGDPC
74bwAbxvGwDBm3dBKlrqncHm7cejml/jaL+kbyqszNzunRWgrGfS26JUWw47rrPm
Vh5rC6NDfWQJyUwkox+FdebbFOiQ2/ZlEq6dKzQH8lW2V+BiQNGZT6hb3aWshQCt
uNdNpku2FW9DSsgvrjIBw74Cljjz3DrOQWD53l04DleQJF8FIARPtqg8HnnNQNbp
WbN4Tyv+LDSoiGXTJwcFVyevWv2xA9Oydc5n5HRneJq5U1H8OhvnX0fVa3Z0eXhS
rJtJXrQM4LOluSktZ6R8x3kLGH41whoTyLZ3ILnaJnvbUeZXyaNSNSya+H/vG/5E
XUoGIG3lPdpKEm2t61SVxRixbcE0m4IyBvUllsQwt9uuLGbvUB6dP7ITD4cXV7oF
U078XNI/XYuBFkMaahJBP1ubCtc42vO6USA36ZqFMNuw9rgqlrkgrHMhUhzJZZ6E
6B4bB0rngnj8zkPuh0yNU0nhxisU99tDD+h32TzlVf99YtBrHI4ccPz0WcNek2F9
tJNsdBQ9E8wQWXzf70R1Hs22Na638lAGGxXs+YU1h+a5YCQOVdXMfEv0OgDblIhT
Q9kXWgZX3kuH4wGIqFNHaUzjoVhPW61bpjzZJ+In1L//iyGrauP7q8pXwHKiXpml
jg1TjhNlq5Pw5gqlqnuOHcYljd72tUTDwv99M7XdtXWDWpsTSnT2EyBJhyiSDTKT
1LkBC3prghu4IeFrJGTFy+mYnmrZ699SVF/QDWQBjEGh2ELI5im/VdYgRZC8etaD
3wJnzc9Owj4LGMUjdqFuB6Rpj6CJrkqzJnv3xCxJaKCjacQgB3i1ej3+FXq8pZT0
6bBVFMk0n1quY+9jeGG4dmBIzMuw32NouSB+/ccKREY+YlpbwfCuMLfs9FC07Wam
XN2jCX4KDdHJPjdO3rovLTsWyJnDZlAnLx4XCg3pUHBO54z4raHzVWJ1iTCfmpFW
DW5qCBFZ8dad3azYQJn+y8Ffg/TW0iTWNcDwAJzHmL2RKTSISazk2TPKYKwXluQI
4sWv02yvwABjF12a3m1qtmcSzxsLNtF86SOr+5VT43T3iD+wmZgS2VQ8fHkYpJqX
qN8mKa0/5ma2Pp3EUJnslX+Sd/zYC83zySGqlu6sD1kYrFIv8yAYA2Y2v+GoYhAI
79BLmKYPd4TE7VYhAtZzymgWX5XIgOvAlhsT6b+JQLwbXP0A3WHrdpo4iwqmt/UD
BI+wHrxjbyab+POe+Bz8TqDlZsqrU4O1NNtV7jpKIo24pGA7gAcFLv6ijSUWjzR+
sca0sT8D+56xDMrqw7xssK9v/Ue0sjVYwaWvhrmjZRXGnJAja691IYg5QdXS+/b+
GzooECtBqW6sJCBh2RHtsfndIZ6qhvWdEKUIRO7YirOTvVZ4zJQF2znkyXgPh2UK
++xCpzMAfxXRQ3FhTI6fi/jB2/WWt86slohKO/5s7hrnHfwFM/cT+Wf4pffuH4U7
2TZY5CVsdonz+gMtBreYeug7SQMrp8gbFiWK/Drj35uR3DIwwGEY4fthnVb3Bx/c
OGQmnjrW4ewpXCOUqVv7xnDI3JDyDexbQxq6CkEHjXbGda82DtHGnT9nsAFsLVlb
Ukh/AjVpsz6ixh4zg0HV5EBlVUonaGSEOZ4rO5BiB94gQDpXSAj77Q2J65RXwcAA
j3vIMaMB4EB8B++cDHXYNJmuMGU+k6cxCsw9wvyeDditINLdzqpPkGFs/eWlqslg
jcLtIkVDR4vVOmSfcWKILTxabNoBrrUju9KFkjPmx3cU+lDyq7AbWaB+GOOAn0CH
kF3ePkmCL8SwOQRviy042fp/Y0uWULc4TFsGYN4pLeRZ6l3lYSxR3enzs0O6WBix
8p3xhYKnJseoQwK+IANghVDNDfNI5uW6oSq9SGY/gOKEQ4Tgzy4W0e7/0anKvMOC
aysuyrwn9597CO3nUCMgMdaVtkumfZCtRArA+8QwZ87E/Tm68r0AFTCFnewHzvHf
Lfr7Zk3995qt7Ao40QjzD4sci2qFHSJ3EkKQVrQIDmkcSBNG4/lnRp/2SFEqczvy
XSlAlZkVdNYpw2LSYeAqVDzoiQDwGdJgLzOUVIBP3fnCJ3i/xipxzFB4N41GGriQ
O2zqDkSHLIx0LR2lxy14wc8SPYVVal5eI4EYTSq4bjmM1XovuG2+C3OiYDhsvlru
X4JOgyK89UrMtbwZPHkG/BPIQ2+s95X0fiNq5FsGqdylQV8XB9ofJEPoCfcLZUnN
wFlzoLajGZh1gzwmVBu4OSuJDDKBFIu5HNhgfM+IGYwGsoZedSEHPC0y0/RVbZQC
LWLqG5kmdxHfhlSY6bMrRaOOV5MwMM2Y3ZcSiYsu7mOp6ERz2A/vA0WfjxCl0SBX
e2jnKNV1nCZroue8OQWc5SHZM+hZxrJ4BmgQO0a/O0Juh3+romrrCA3W6G68sd33
HbaQA9eRgxermF5a6d9ZaAFqbHUjVHqf79y4jEa9OToVFEOFdw66/WKaTYY+j73e
VhtikRnCcrNY8BzacG9X8F85BFNTaJv7ZIUrU2OWN67fhYtMiTrogwGHD/4dhHtv
EKQ3yJPapNafkYFYDnQDsUKlGRj/cw8ssyB7gw3yKwY4cNC5G7qjH5guXXrt7xFu
QUX4MmyFTsb+zsJw8CzwVmlZQDs4/iH+p1sUAI6lpGOzZX19DnIJeYzKndSokpeY
z6GHhsJCVip4/YSI2OOpgI6MeQKS6qvjp33IPUD6+Di+rvt8lU/IqZEDJ4/Rq01z
052G0TMscRHPJU7PQj3OjTkssh7+lml2PXUwwFIPRJws1eKacLL5RUh5HWpwQ9rG
8BH1lIxxuPsLOlyc/+uUA9t0FMb8Xmn2fgjuN0VSFMJrcn126nIsaqdpkpUhZrYz
XXhLWHhFk/fO9TPEhZqV/DHvp9Tr4QGhB0WA88X2ulh36XJOb+hl3peDwhVlIm8U
eQuE/5vB95M8eCQNONRQIdaksWLKsz3wlxd4F0GldOeuI0h5j+z9oYjbno8mKpzn
mlt10VX6inbkg4FbnwnXNtD2dgcguELCKs02pb752EOf0wHl7JEBeJO+ue1R8lG6
6t21fiaTGmSDArKf9pCel7IA1jsZNFmD0RD6iq5OfWf39Szf5JAp2805pq14wll1
OgGg9kYSgW0288ajBIr8X7XWw94EFVzgO+6v7DSHma7A2qs98eNkbdk16/DPl3Vf
c8HjJSEi6VvjJtzPxOB9a6G2CvwXEDV5WhKLmQiK2GjONzDYLL3P1z8dgVRyQ+wP
6ZupmWDmA4KXn4qRl4T27NXSB03q0TH2jNoxBQ/8q2wDp5XTA+amId/FXV24clhd
NpWQ5hao71TZwTKWGkRIHR1y3/uP3OP0YL652549nvHHRuExShYgXZcfHp41Qv8A
INRnczxSJEdI+sf3cnzi8mCJF3+ZQvatoCcYCgpyZddoyLy6hPpl65nazhCRFNmT
iYmk9wD79Q8gztITCZG6z6sdaVRLC0REMaD1bGNXvwXeb0shHGJq5SN/3ZWLHzp3
LJOnB84hmcCBYxhxXyZXB5MVi/s3XsF9YKD8K0JjfOqsV8jiPGKd3od84r1ingK/
e+nbNmGTJcnCeJU8W3gss5wJ7LKoPujL1zC80qTsYDLTpBrXZdTXaU/DeKfQDBX8
qm01tYqV5ctwB1BEisD32ot0SZUQFhwYUx9mtLAIC02r1Uzr1FTu7t8lJcFktW/c
+/nNmwJenFLj+N91VaI192JWKYuoTw6KVucUtHJgEeJ7d4+ZS/z/l/RP0f8Ibjlt
7kT9nRM+Ve0avUz4xLnUatB9jWgWaJYWh3zt+Ps0PwGB4hYNRvKlcpKhV4kOHgNI
Sfnp9t5AwJ7SlzykNTtU0g218lrttNHoN3H96ZcfZ2uthkT5pvCtxwpNRm/R53DK
Viuy+HssiPJuuiUN9Ygw9kAjzhJ/cv9n7V9AMwj6R5tdeYJI7cOq7z7oCZdk60t9
29JtlOf59WFWWjaKSyyx32tNd+jkXZhi98YdESio8qYSliYQRtdekx1D3fz9gIzy
Wx3Ccp2dttdM2JSZbqPf9gUUICazY0BxD8eoho3xSyMUip6xP5KC0Im+XyiOXzzA
eyU3FXuwYA/hBV/2lBxYHkUY/KT83kZmMj7k2weJXPtX/U3Vp6G/eCUCek33UMrn
a4S/Sk+6zBPgt0ts68nJa1bed50hZNfcQLUtfi+WStrea9gELKsnk9fkasbefehs
qgxnFtJbXDUxN4+U/Vzc82ytqZrGUImEAsRWl6R0XJSETan44mqGu5pNiCzIdO4x
CKMSUpimoKViZ1ZvLMxE1/fN3DbMNoN+xAcUusjKZ8jKo0UTH2NaX+eLGLwHdo3g
ef/9od1jXCCN9dtizOxloL7es8qGDzU/dAl1xrPrIwOqr6A3v2NhFw9SjzJZ61cS
s0tOQzAuFpmVRBz96znvOUDZKlBkRoPKwH/+s+TCpmG/OWAmMZfYSiSvy42x8dMr
eVd93Mei8x76ZglZ3dchyiwN0FvnUirHje6W/r1RThQRdpn6L31DI2wsDz+iIbK3
+5oRpyL49XtvWwYnvO0KVNxZC3hrXkjKc7qvKLCzG1IEjsnTP1rDOtyNVHN3EzFA
BTg/GDV6kE+43IbA3lo1wyMbDsGVweIQ0Zfnm2eEEy2krsZbupnzCcqf/dlSRrXK
hny/AZnSA8Dvf/SZZK4Lmhi/ScRxET4kfF5YXpDEcZq011+a/4pwOkYsN0zfKOqW
R35P/CRc/4U1uf7vJfd9NtPvPM6sV8TqKuy5ZtasFZqLJuunu0T1o6eSQUwx+hWn
SUXSIvMs9yLOcyQ61IonJSqWYgMEUnoaE/p2EU9PGsAzHqGiucr4cai36zkjFjFY
M014KRGFw/gqOoTxaXmkIr+RuMcw1nuSKaswouGxMmWlAykvm09HtlycalLCaISw
nf/UbRi1m3pnj5Ti5cwhcXr9SE3jk95m47EOHdtapEGnhJsnkZNszQkf5On/WXop
9LaLi/+2i214qrLTbgEJvN/jA6/2Af4wFkrBPyTgBva5eARX0QCuuBCnzdX4yUlH
LDE33OOMaah/9Z93fs7pYmWyvJMufXqVsfw/0SyLhB9YY48avTJeWdSKw94NI8kF
ryBd+BJXeqb+VTN/FipZkAb9uoqqW3+RuVvjckl1mUfK4E3hvrEdmbDhsHTAvKHz
7HZXdERxMqzS4eMftN/xO0PDw0FOYxXnHpqtYs3G3qxhcZRY9OWDUgaYVUjFPvGN
8e6JDqUUt9H/Gmn9GoB3SfX3EEgIGDc8jnF4CqlAYTUGph74ja6E+CBIVny3O6Pp
3eeUjUE4bttWU7wStnYvcSwzwk1fSaX0vjiJC9xWcaXrICBwX/sOtKnp+rl/T+IK
kDFe4ZSMFQtRfCvO0PhVTPTEBJEL2LPGihP+MJjA4dcfz+YJBjlSSicYMIaTSant
RcKOT3jrnoz/8ln6zoh75Sj8A7up8X+dO5IlEfZLt5Ueow7kdf01cAHrto+ui9to
B5bcepKxlbBOI8E/WTF9cPpyayrt6zhgVyOxZguPci2scHli25eS+VVfW/ybMBAO
/r0iCHkRukTkkCQwCbhENbNMGVe0uYEEjE5kEdEt1BqeTqSlREKigs71beCdLiHO
lPIdXcu+lkod98SE0jminea2c+VrPn5o+uFPQutYvoewNXU9kv7OhzyJdkJLM2Ps
9zlap/NqJWdxmiZA9RdDrRMDTgagwzBtzH4KwpLtvn35C5/85kbylLYG9bOpDKuF
Z6d6ZywsusHdH0wfE6BsoJWEf7YkUQUNs6uuH48KmJX8ujb5+pJGYd5BgiPqrDTh
vBVYEXpcL1Kzb8G5e81QcPFFCZlDyOabbe3ifpjd+283bBmVbU1exlecX69Y/0EG
ppszPe2UdDabCwz+NJSnQdPfpn2kYf2m0AwHDv2cEq8lXChsj+vbOW15K5n0c4o5
hRSIsNQWwhJcJWZAmIDBvtOkSVDcWJYx3MYvdG+eHhVq3l1edsipu0WcJpudKvV3
jrp9WWrTH6zWD6IH2BfqDFk61SbCQ5fZi2JkAKh5FIJ4xXKc8DRAjTsDiaSB5CF0
lANYjMnXWXon6FqdCrsQTa6A5/6lMHWFKJaIgWW2NN8GnB8fQdnRV4boXC1RENQk
GHHAFn9ylHW6GxmU9Rv93HUuLmIoFJh4XSBCM7MBxTLhio/WbE80GLum7MLVFhcF
asUFGFAnkVVtZk2dIMhiUnAVuXq06MQtbPBXb5ei1wNk3FrYpzp2WnNJY3HBVvwP
GhOkGrIOA/fkasFpUn16ZgNPadc/tI1uRB/kjzhcQSRapTdBjH8PcKaQIFnWPWTN
E/uK9UKO2+Q1mfdQPhi5zf2sOAgsYtSxjbUowCTKy1pXPBsRWOiHHFBQnl/eohSo
LdplM4atYsf3gsXINgrTl7nucE2s0YmlxYD7xpm7AR5h28sbOm/5tqKfXUgQF/7L
DVK9XTjdyCFLvUCHcVrEEubmwS3aNHB7CascxNDdtSxQLw+qUxpLcpugqkhFZE6b
IzrYJ5iSOIgeuStbJTMQM7QyLwQbYaks4R5bVkVOR7yuyGUU2cGQSSY9+p1gsJ9M
QqZgaeegfqwatWI4HeaZgKKCLwIlO+Uj17z0ceHIojtB8ohDORAIlJxtipCUQvWN
hJ6+OzvqwRnqr0e6qZ1fGSPSk7JH6pMMmEbXCNDja0YhiYWAKNj2pT6fMec5m3q6
rFsuScFFOEbQwVqlKte7l2iLhjy5E3pLUdp+pGYOwUgA9umENm/uEFds+rbtrJXD
sDMR627V3nyLECngJ8UF9C10NhLqL5qsUw/u1aA/5T68TS6zgtUwGXVEf0T5BFu7
beJfazf2+FE0MIsMYAc+JU+9BscxNWeg6sqmOp7cdxbmS91D7RxRwQrQ0qFBI1m5
lJn8EJ8+/vAvkCVNAueH6KKF5xQ/idLIm+xynH+Fgn/gq3nKlw0+bOyaeHeno8uk
xeasBUz8IQ20JwGIgZjI+dbCuBgbae7M5FPpu2nMAPArkIe9TBWl7gyuxlSSUkeX
/iiozx23hEOug3zN9haBVva1rR1FqDg6yY42cZBAynU2hNyBvnBgFYC8bgY1gBcm
yCjHowkrvkLfhM/YokNLL+8w1MldlSubho96F6L7J3nNL9FdUzKA1jBWk6tyCzWh
064wdMaQXLq2IYx/jll/ecro+DkYnjijUmjxiWMdI1zCpqL+tR3+kAB1OKNm8kbw
UwMwkR6n5BrxjV1wrG7vsqfcto/+Babt3o1KMC9YAeVatfaxqn+IHfgjiMhn5psr
V+8pBU9xnUGiREmfIva/+kg9lD3MhqCyGVV7dXuRgBGbCVgUzlcjevev5W4TehjL
mMhqxKVyIaPQt7AGbAdZE8N1lECFpMzMiApJdr7JHZaEP+mTqJzNlmk50u37/JvY
Gv9LBf2lNmgCAW2SpxARWqtSBokSCsYFFHf3dB65gDTM0oInZcwgb3gIllVPgrOo
VPZkG/aP8x1bUYrBbSAHTO/e/OGPWuNjppEU0dqMkHIw8gg0wnUFN6BcwG1eLYot
6+ps+Cb2+Jfuy/fPmV4VUxuh2uOiI4/P5UN+cMDS0HMkiykgEll8Dn7sFoOAWBDG
hydeY4MYZSvn5WDUMiYH6/UNfm9L817D4Ox0YqCwmEVI+USwWbuiOkggYcs4vei5
fx65kTtpyafWT5L/6Z6vFw4zMq/4uPSsSHWxySGT/I0pCwoMAqQ+8cSLWCqPu5sy
qBTc8AIbBuzbBBLCrMJRolbwK6nlamXXwZBEwbiOkTd0R1f7W2ktd5ZAK6iI8qLm
sliDpINLS/WUiMzHXy59Udpb3KH4Xzl4FDayfjQ/7Rt010OPGmho8UD37no7exWY
tCfR37e/7g//3bZ9mM32OWhqHz8rf8PcmRzJjhFgS8/1lu06So8hvvIsHFjKG73Q
Gjv6d3rsgGKPQqqIolkRmv5G7Yq7JX9/7tbLyaVqt+FCraKNuxDXmL2oejHeiAhl
kMt033Q0eaOkdhBkFdw20JtW87DfBypY7RQ/46Tjq2IKxMVwerdM1MyiWs4Of5Yn
rdV6//cnp7ZN9r6JcXH3Xk46lyKP4OdIj9PnDIggz4w7JbD5AanDdc1mG2ReGkLB
8/v6mW+tAifh6unoQoq+QX0NzQlGJRiE17MoyLc5WQbcvQDMWShEfvJwxE4JxDzY
4bFsXL0STWX0EmATJ486sUNOLuXd0dUEZOWLupRgNsA0SRv3k4UsdnRGm9d/wmeg
PJ35b5BuDQ1sb9k170jpD0S6fkIS26H/VQtcEwCeCvbx72n0ccwbyAMmcvvh+Wiv
2zxUpxaj0/Fnm7wQM2P7tbqJEPNBuO1A38YHsi7k+o8Y4QahBqnzddAK9MgjjGZB
Q2w7caq6tapDx0KeQ11Q/887+5LOdy687qGRqLrsBE0Rev/DnLK2G5P4hNQAhUvH
8Fq4Dd7wqEjSLErEexTdlZlF+mec07KJHJSJ4JRflHSyPuzOOTrIMNTGCLGmdJhy
lnNB9ihAL4F+jqTvxqNMsaFm5kp5tbjzzwmOw4QqrfDnvuUn7I6dnrGRV5RO/Uzz
XEpGr1HOYwB5h4mc0vBZYUPxVQUC0SlIh3CfpsvKPYXgUDkckZOyLiYQtK3OY4qH
qSAEEoE744x8AgXdkPkpMqZTjFveHZYFr0jwzyFAN+aj/pux9D41NYGprtKqFhLO
jo2z7vwHamvxwzRpdCoJDGf8lYffRerDdraJxPjMTk06myphvdHgfsf7flJx59VX
+T05hYSOayvF4COdITpZQZXcqKRpFM6+0WramItRk6ETUC6mr8Oia0KUdcX6Ja2Y
3yFFgny3AzpZ7n5aSe3sK6k4MPWylYUYrXlFE9mmA/eajKn+awVT46GCbHCFnHMo
Hoh8CohDBnf/0viNbhLavuzb37mCs3FkizTBQ4j2i5d9VKTW5cT5+PM+uM2yCtBV
4Cgu6spmlQTm7azd+K3A7TFG4CS0hOMGjahPm6VduK5+ojtRdMJ6UKPjlgUu02g0
Jwjk0iJFWX9IxhnCL5kIXFHFv8eKTTmJHhCQrtEtpDMT3e44rbP3tZChljeNSf7z
KCBwsnt+XnaGgLlleOvhTYhFf0ahqk7SKVYuWvqZjH/01UoWK+JIpnYHa7MUynd1
mJkPFg6qBIOrlZbmjp5sG1Y36bU1Dahfl6wxs/iCSzAdLvVRzVlmMvWjxnxIBZ41
EC73dC5+u/aKpNgMTp08oXDdVk/q1bkA4+/ceMDQHjswmM2MHPMSlmvMCDajPMU2
v1U5nAZ2FLuQrszkOPFbU1B6xoEkqvg6hjRGihShTeqCDyG5WddYjyp2sANGqIbL
LCrHqJSW3rMNBCEbm3RFvyzPDml+pugo6PCf62BRx9Fet3Yrev71yjPf8iAxALBZ
8uFFASE8RrRkoYlHN1fuHjyLJvJ7GwElxxi8E45u9j/40wyVKIOQhunElujIwcp5
/1HVBhZJis76zCAd7iSqQTcfnW0DyzIA607bBkzPJILtxWVXbXFtmKkVmNi2GC5+
XSr/BJ0wT9XGIvsanoX4W/V+CCIWgwYRSis0TTahPm8k5SuFDzyj+8jMSRJTv3v+
DRc5crPBsoKwGC61Gw/vHrOdffoA50xNXH7fOEwvFRO+jhst/dRluNpp7n06XDZI
oWG/VwvE+ZNA/wmqrFnKZmC3vVA7SbkMnbYQFHvkvOQgykScxqcD+DR4YF0ZhnKm
IsYtXrRgG/YvdAaWv5L/DHOStTpXNz0NSxnZXTLTJ+wy5WnZmb+SWLo3fWQlazln
EibpgrePcJ0RRQCLCIUHjZwcAuvRKCP/i0Y0ZrlqfAVk3nqV+vHgOCS5joOVI7+U
jxGSxZXPWNlkkIP/gYgwkzTovkYPKllQ3Zsr5qIj4GIqn51/bAf8ROFA/MpRQwwM
XjDBLmRFIc81alugKu2jTGgy2Lw6WkljFeZw2OUfv/hVADHHfK6tpk0Jbcc8vulX
yxhIPDWnsjmi7BXbSYeIzoZR3TsYy+MxZAU1PUa6qkkXPFyXiAUNqCDut+zQL5zh
fOWzbGqGYyfYvY6WkDXGzW6gApCze/6NWJK7rfops0WIEFCn30x5oLG7ISn1hxte
1pzYU0cB4tYL3ogIzHtNrzGhX42RkaFv8wWj0bxkshZu0EJeLzfe+XtZU3CuS6Xl
olV0xiwEgG1MH8peJQEiIW81Xhusy8xOd2Z45iAWck8t9Twlqm6n8EoSj5Ymztpt
mUMCa2bjaVdYsocp10sYr0xxOdlUZaUkgyLWHZpWwZ7ltc2yDJOKD64gTjuPpIZ+
cPSXwr6E8I6WEI6CUUQIxNgBe18Eahk+oR/jDj7R6+jYMWiOzg2cl4YLZZKzpTjj
qh7C7QIxxaQQ3oKjuDhQkrf9x9O2sk4q1rHUaVM6sYxMSEsnPbx1lp/brFkFg1XM
H3xuOZCi2FErycicqlU/1+zH+/GTp2nROQCKJO1EVGT4VN+WSqLoHzuO7N6Sis3P
ndka24Lfz1GCLA8akGp5/yFGmMer7vWRw0gvLTeWqbLe+ETmVVULxNaX04pR0KJW
A263DVLnpQNYNCdt7htvIdhV2XE2xmEukhqS0dtrd+puJkSbRVYDU8hTFJSV+L+Q
ThK+k76qCecQAIXnM/jVzzj84KlWn2MEDdZTLowmQxSyng0y3DkwN+8a1GWeYEeq
6ZyR4A2lUQdtbhhcCPTqETDGapCjmehXHhPGgpEcK2lwIyvTAIus6k9FIb65HpP1
F9lrPEgh7jjpRfB9aOATTXvMHR7K5QOzMesBtMnjPM7KGj7iKtZ37DSehjoivjdZ
Pm+Rn0/d1AYGXjYhc3d6NjZjHyogKJfSvz79hrOzUd1Kwm4DNUarAzkA1j3m9KML
W5Eb8qh5T88pTnetsQCp9tmrX/B+MAIp3CZzKJvUyzK4SK5mOBsXykGXzZqmPRiT
M2OnKpe4LB26ampJQ4z4KaH2onL6BZXRxgAlgqXjNF5X+lz4rkWgTC45Nti+Kguq
WEgTlh2oJjnlIOfKA+ktxqe3fFxNMa3PamV746B7Lmd9ZBvcrdzrlm271t+4sCNG
EN9ws1v4/Q4mggcFPtLFgAMXj0rFGnkR1CoLNSKMam+hVIr344zvRVr2v6wJMBkP
J/1Xb382wsDVl/DJzz4Crqg3MHRWwIsDQgQAvXP1S1BbjvfiWasesTmRH9guoW+u
WcrJjKUm0nUyF2KD1HCSzr/VpITIi7o9qfip1WMd1mMCg5zFuER457WcID1f1VTm
PJIFiMr2L5s0GY7yk1n3iF32tlPp4OnwOtKtFhPhcrnROJs1hffcSCkK/COi0KMU
yO9rwj5x00vbDO9L9nHepAC6gPAhCvtm5R17n5i5nky3ejkNQQ1C6raIWNQ/MsXA
GuW+lAMFoU3LBuHJWhjAl10qxHrqGkdhNVpQixQCUb/oGzVK+qlVCwv8cKcF0TSH
3vhQQ0ZGtdiRLFv9b9PiHCzV0R0rOZvdF4kVeVAjjdD5bnMGWTe42pgvYCeLWnvH
xw3BtJjvNIBE9dlsNwJePKYExv2pe2sW1sMQOcc1foiwF+pP1IyLC0qRGnrNw0qD
eHtHMErA2unJwuOEYIPE7Y9Ov5fs0fmSbDrwLRn0naF/Pyhh+R5HthCvEHPv4y2T
62K9x3l/Tt2XMa7JPgPAiOzsz3IqbZm3brhuSrMJAsKZ9U0lBvnspRpD13uqWMeE
uOwlBDjCax6mpzyfPrzNtEfyn37mXEOhhuqXBQHbD0yaayh5J826sZ1HUW81mi+A
fKSTZi9N5o9VaXENkFZSfbNmcn8A0cceb3AEX0VA1CAVoBjSWHRV4voafpO5CeTt
0RtRgonS4vfpmBoLMcuS4uyXqLiJd2krCSHSGbN/KsyXP3NvrROE+/fEIOpEHIFU
vhNdiUoGh2DojDdUf4NQyfFWJpkEKlaF9mBJNrQnw5jixzYqPxokvV+HRgQkYO8n
Ig/cisYRNJqAWind7fmMYrCrIJiZLH1Iotgy+TTUKmm67dRWK7eUgXNi41zrTH1g
WZJR2gLbwUZA/Pc2l16wXRrf53+Xgj5pG5S/9ffj/cSShj9gTODwViY/mXzpdKeP
LKz1/KfXcUp32vRwinwD/c8oVGqifK02zUnnJTuilFwDVD5495b2KYwxGfWU4PRa
uLAEKaD08xK0eYp4hB35YPO8DuDRIApHpXv2odZHzGCtBGS1tjtpYCNlVWCu6Tyv
vnRWYBjeaF+zmhFKdJRBEqxiKhJns9XdWnrgwq/T6EWqHgXTZcDxD4P8zuokJSFp
CyvSqrbq9ozG3NZ3Ha+Ol/2UfUM0wyyWvOZDhNfVfasudIwx/CaRiL9SVlqbPDIH
cyq95MbqH87oKw4GXVvT+BLzYvzH6bpkFySf0Uwbu6SpsOXUINQ/cZzssUQtFnWa
keas9Miw8+lefBjA6i/hDwX6B43Kgnc2TvT+KZNBUtw9ohq4jQzP6TtNqTT9S7pS
vXDG4BTSWQItIVqEBQRGhBU40+fduahTNpz4AdJ6MFYvatukYGmznLHCEZ/wk0rz
70TwQgMw1jtBK48iZ9vyCEBph2QYCAp9KKngn/fg/qcCdaXY7EDhmUfvMHjvNZTc
2caI1UPRorHgOuiSV1bgxIx2nZOHjVBJk6vtIICqF3opdO/QzXG8UR/Ajexuj/xw
U95JKqamkgSh++2t1E/3b1TXLbEhYwBVFRLvnWCEW3KikqHy/tlWKDXdcsxL3Ybh
ILWHglJM1WIo/QZbbwWebLNYHvv4CXx8xGy68iRqd+IA57Z5bQsV4rlVUICC/UVd
SPEvnlT2tEKZJM/N3W/xFqshwTEuAlHiMRiMO5PBcERn53Jg6IhOVe/4PI85Y/nd
LJo1SelfmNqggMqs4zRXvNfiPfmDPILKu6NDSR/pqZGxPynCiPQdwOYD0MxX+aVv
I7snn74zRy5zTp3qNLVSZktLEa3fLrTt9NMAPVvkprtGgn+qhrhYy9cNzF4zSO8P
tZjLgEFdEcO1WNzBztxARaSEAdBc75t5uRENWfw4owhC45T/VvryGjheWCQZjXMH
fyrKh+TaU9dOtsCTj0Z/euMUXmXaaJN4vN11f6ihP21FzXxo6abTRB1JVdsou3lX
jN0E2HQ7iBnACWhEGdupGzgojXb3IgTdpTOY014OIH2NesO3/akXYol0gmsHliOe
2nV5jxvS3U91rQB1G4WaypSYiOjvc3LAKjYMUS6uVYHR7MN7NHtQxtl1DFe5a3uI
sf6iNYkmagdDRD3QcCj+QQJ4IlbC40CMwTVNCQWb8Ob0iv8ILI9pyXYHVTd0qshV
NP/NTDr9L1ytvg8pV1RoyGU2+irFuOmZSXLDCPARkH9FMde4NCo+Ahi0VmQauxTb
ONoPJKF+K+kl4qjvMfJ7CtPBC/dw2+Uy3blbKExtzjf5NVAUNfX/AywTLAJWZ3w/
V4IwLMX4kK8nlnEtp7ENb6C95SEE45jBeZtmErlwYBewU9dBjSCXoaot4pom5vko
zC6qiqBp8bEuCWCbT3+G9Iw8K4PlP1vMpkjGkDtEI0ViBk40XLrGxJgCewnzNMPV
5xqE5Lb4uDMtAiJqPe7HYb49LwlWR5svrOhMnMqTNFJ6tHEBm65wdUEfUTPoNd3b
5dorprFXjsu3PTXoEqLBzTPTW6Hw8rfXwlvTLmsKQ31ehtBmLyRYCmmkbkrokHoh
B52v8ncI14emqOKNe2HA8l12HL/fmz1ymml877wH81h+rKRt4foeY5hvqFYxJRGf
2CLis/WWu6yheM7fAh8t34na75YgAMfnVS6mkh44chRNYw3wVk88vRP2ijMqTxnv
eXE1Q/UWy2D1fDsmvoKFVsYl1qmhq8ecz6BLMhrn29MOONmQSuJPQ5wp0HNCCJH6
dJuLrOPw/+cmX7q35eKxd/2N23oRnfMseUnEYlzBjb5Nu9s6wHGi7umMPatSQQ3V
o7Ged/HL0PXp+SBJgJAWa54xuYnRlLg7BRzCSfCsXlCwHqkhA2920f1g/IOVCPqh
Y5DFzHuUioe44Ufp9mzehhzgn9pMfXW8Jxspl8baW0BSvF3ligVETHhvlFQIuGmQ
KJFS+5sX6/wsBAO5azOvgQHrAHYeGhXvx8JCi1+0oMsbEWlAL2gGnJdz50QuPcgS
E/AXKjJ4GjRXdOf0paHAOA6hz3XVt6znxWuS5/Ej9yVM3FJF4k7N4f3lfPoo3xQt
FaCHrnq6qNyoodlDvoAvNVIAnWc2Fkfv9YAuUahr/MiMlhwObeEEazjeCYFdwpe8
UqRAMW5XjL1+Hrr0dzhvZu3zoJfXiTpKklAiKq3MmXOSg4h31IhFhR0xlLQoVziB
8IvDotayXrzl9xT0SAvztv3ghpiqBz76Sg8MjP7OR0WPvfV01fXHWkr71aLO4v6V
R+Puri9xHWYerVjCUxcVFJy1ldRRKDupkFZ/KQfxHwGQcfVLtHqC033epplvuXaU
Z/Cy8LGyPllk1jTZB4Np450iJnfihy3UcXJmALLXAxWXs2ZczSD0UiTHUmXM6YQ3
MTHasFqAlx7zA2XN7Se+yO4HdxjE3k0NkOQf3cDuRDM8pOfBz71NUEzdNPEljghV
4b8i4Sbl8tM1WZBtuml7UKqNJkkQOWopgUSMJgP9jxImOXFa38jaajny75CZ6ujH
nX1/AzhpeyLFu5m3Zc0ekc+coVWRct09GFOnFdfbpw0kFnvfpNyUNxkNCgNYbuLB
MUZiBRlwhv+zD2YID6BdtLeJesNuVVLYBOG69SQJoNptQJelIWRLWldAXBkfGvnb
ps40L09YPbg+DZ8daUA6Lsq9aZXgQwIiH2MuxibMYFljkcsJWh3nfJqgfmz6oNNP
cDT74r4DswJXgnX0Yy8OKYGyhQ21wWDjiSp7YXnJ71Qys3qLeQ73J1vYH02zqgce
DaQ7x0MbFtkpNuoKWeJTfDobc1+AwwDwuWo6nx7SD+iIKOEuH+9JD4ZPS+0oJVS6
CZX/Fu2HklzLDAgdhPvJxfK9DVKyPDglkMUWUqSNQ9/IMPsSwAOB9ejPX+0CyQe+
wjGLMBfYJ79lRKdKUf0KJhLvXEzSiBUEXgttoPcIeC6Js2BfsMVAgdZ3lycGOfr/
I7ZnoZvm9ZVB3a038QEUQOnZkkRkWsysn+kQ81P4vfYuibCGeJ76mIxTAmV5xcIZ
z843XlpfH2la6MFpVcWQbAuSZ1os1CsHPiHD7pyCaISODEOTvZQJi/v+uS4Ks7Vk
Tp0yfkIWCPId5w9tBx/9wcAYf4FGhzAM8CI9kxf3edYaI3l8440Iz+9hHCbKlEt/
albeYB/wHzxurzCO02Yclna+WjpbgOQEugb2aEllPdk01oWbPEmmbI2KyjMJdnkp
PwZecdpSNN/Y9oCNtCZVnr6m+BzGvliwT5ITxSXOQESGK2COlNaSk63t9eJSw3hQ
70Fhza0w09R28jrWif8qJCMc7cZI0NMOO6c2lsuhsLbVSBJARD1syotzqRKoyVAY
HTK62Uzbcon63FzvRefybpzdUEbLCUwOWtCyfM8pfDmOGUJ5UhAOFwF8Lw3HS5o4
8o1YHYb4Hycg/OkaHF8NfGaUs+If9FoxKJnDDadBFtvU/lZhyQS+lZedKLnpJQ48
Znnk6a/4Ko+vimMSSVFioNG8/gjZNHDNU7d+jzrDNkNLclAyYQYzOl5nbg92Lix8
upQI8xyeW5+p1Hj0SiIdoXl+U/9gnC81sJ+45LIrTMtFfMpL6oTQO7ewxJHrkbNN
6UpyFfN6CMh6UOEFOVC9Y3D0OPbt5J2W/Wl7EXnUVYH1/1Ogb9EzvX9ZAmTQ5aPk
UwLb1LlHJ4hwFOMHxIpIum+rOkywbr4KnGpLZfOpeoet/7V/AZpkbnvdE0PWXkvP
MLqtRmDBGKVFWE9BE/dBgFf9GxaVS7R4D5xJRmGgdLgDx/7xggM1Zgy9Um14hSdM
h409Hj/KQqxqdDylYbt4UhWSLmesPP8OoRpMjptMt0TfVeejxrrhQdoyOAt2B+wn
ilsainLLRSsU014Z3zqPkxCl/chPchv549sBBCUQfl7rVNVL5crsp1y3BkioAEfe
vUwOuPa60s7hlki2UdxaEin0Zv6aoSJ33P+dvIddjkyPQ4iuW9PVYzuMpftpG3xO
6aQ3UA/2ekyRWpNcQ0o+IWje+mBDnLn0Yd1hggfAL5wmyjzb/MszmGHdC1nvRmE9
k9D3fSRETca0KBFSW+vV610dwTHJXi16Ad/12HZkFLiOcVRNkf3Nxe0pmOmxBUAm
TmV0dl12PhFyC5oPNpjIXE8CNdTSxfjN0X/bVl00yqTJpEdpXMjqdbGBSWBBLcCe
uuuL+dYSx5CB0KE50sxEU7P0cMd959mKpFB0SOdWdXxeSwb6N2wO+xIr91C4Knvd
b026ROvfAgvXumtfB8xj2CD/WMOOUWxG5qIchQ/9GB5tfym5dM7wUYVvqyBmlJFD
7zk6hY4uXwk5qzR1ihoEXdmt8toY+M76cMKYB/LXfLAnnAz4n/JvkrQOCq4cVRgm
2K0OkYpQOGHemENUsjJ/8H+FglalNmNh0245p9DITo3ICKjfoZ3YJ96Egp94yDo0
WqX131iQScwQPLjthkQ5GGzoElOPYRoKp49IgVPe9fj1+/Canqo4+4iE7uxX7QgP
u3B99CRvbS9r6v8dOWLa+uTtX3abRc9NGd5XQ/Ll1PGFnwSB9oTAmyp5FX5SLLXv
YBEqUESGTxwd8Dml0dUtCWFNPDcIZEccmDVKKLEJnXzPIKCv/HA6+84S8GiqZEZd
VrdpwkoPxtyJOEQXil+IUOwd/b1nl5RR6XIjd8sfjlx1COdN/QwRo4N1CbraS7r0
bgX3OjqVQWPJbPimKth+1OJion5YeLlR7qK1RV4arE3JwwophpDAq2DIz2XqfEpv
2/ygFSGy2TLoVGsn22UIf0wGuLT4bJozX1+N7YfsznFTC8yZnZRiN6amY9Uf3orf
WpFeXeHxl9J8LYJS+YLRP6Wwp4DIUysO3Bhk/KbLbIlSo9Bd/LwKlnyxEIAKMMsd
KTT5p7k/N3pHy8uK6n0Krx3quiMp8z7jOTFtHkw4JU8cmhFn85Z3QYzbkah9Azn4
Iyj0n5Ic52R/Ngv2aSc76D7r54o4Lihurp40oZFMmrCr55BpGHNvJCKdi5AK/a9/
rbGZNqZgVeUeWCL85Zj12SrOzP5N687zkqbBOSVJPxq/8NPnwDxeGA0GgQuldBfp
cyUxn2n3TsL9HtnOHBFo1fStjxmVkLbRDzay1IydJwYHsgiCNmMU8/wSXWDCVvdw
jGwWQxd4NJrRbo7h2HgBzZ+8Qel+fKQCKi86fA8/udyauFXBboeNDl4R1QJZADg1
r4sYAhxp5cj7HDHriM5V17eTQ9TVz/ApfJboQnhmFnOe985B7Al/WcvPCVqG8VxR
SrSxLWjX8AIvzyR1m2FczrAQaTRHwmJqU2Njth00xw+DT6sojuislzoEmiNWrdah
CWUC21NX5VyNh0kO/Y9QIMAtFtpdSD5iPr9UyJSfXwXEFdH4pOgj6v9djOMsqMrM
FOgxt5Vg0Ts0QkfiIPxoS+FgQjK+EMMsH6lmViIK7EUq4FHdzE5dTNC8cIeOxTfU
mdSAzG8UhkcaWy4rm5uKW00YWknz5fBBX+cEqYjHNHelA3nd/TPXDHorA8Yem5KY
9iJK+qAGxSLivKVoEqYBYKrYDZ7oE0bOMMDJSZ4uOd96RWx6by1JCIOaJSTmqFRM
aFhksL5wd4Pk7bnwD7mdgy7pAEeS3ZKHBHVRFlci1/GPJw8ThO4lXl5gcyXvgKGh
7/4R2+ht1/a33esUunB4PH2OLZV1UVXy3+2onvC76lxjj69ObGr2jREvPd9KV+ph
jRot2dru2TVeIXgPdo1R6YahLaz3nBrUtMX4C9KqyxbmKJ9ZiXBldIE5KsBayEVr
jVoZ5RGrnuJ6/FOsnVpdcd/PooV3Ud5F2FmRZbAI0nwcasQaIK7csDHqCFXoB1CA
oLr8nWYOldaU3V+bgPfvb9bk0HZ4UfkQCJUNSXKSf7YVQMiyEC/vi8csTep2sMTi
/TLPkaHqoFkTSnspexJpHrWl1r7sUa51uzl5aYE4ipyqsKEIAGWSPS1F7sJjectV
9mW/KcP9caMSou90v2SBy3QGDCimzRP6eOl7r9pgIzmRzyIUM1340oG6dbsBXxDt
h6yfFYqj/zfzG5ksWEFp2Qp6auqFN6f5yCrU5m9h8GWsU3+K/N4eILxC+/HlXlFt
ONtL05/BurPz5qcmhjd96W/eHZg/buScC5G+G714f5qsSLyE9Z2Bqqu+Zwj91Oi9
xOioKssM7ZWv5cKjnwjIkWmkjrTsp64BUkzxgKyQVaWL3/kk0bReFqcuUpPc4hXD
0d0ne/AIUYfMWe8siMk5oMflHPGyo3A2PdLZhsWkWB13duydvPFeuBQX5VgB3sKs
o177iEn214U6LS4bo08y2iCRYJsgCVojifgRBESb5W8b87Jxs5xwyhZBZWYBEEn0
vNUXhJotYL0+mUpMjZsTWXNrvunM+m4HXPd5HAZ5Qq7oUFeNM4lhTj6fgYDXaG6f
V3LLMcoECnWyXNMlTn8W59tBjWzDBYXTotnkL9FpcB20EIwS9msTNMwNL98dSlzB
YtVR1asqWEaSP7FdojLPMS0nZPtazi4iwKfF/6XyTKA470Wey36j6f7A3KednAWY
EYeiDJXuvi/GBXyYU9/1ND0KFZEnNi8QIy7vTFfdCp0XVpJak6+xd40w27VL/PMs
JrrKx+e/Q5kq80yr3NOWY2Nr2Jga7RPMnVJI7UMe+gxDbXnGNoK3H3RGmX1rEUNB
GvxBTn6ctUsxC9bmPVMhq6XuwN1dNAcIlFIveNiWfUciqoA8pu9pFLYGp0WoaMbz
EQataTCKw0D58YQW28V2arf94AJDbNlmeinuxxhXeWRX8WQSPVr482i/hOUqjE5l
nb6zzjtFk8Mom5gZyqnpiPL5jebtFicGv2ikyI9qITU5Jil/yx5r03hozG8cOh8j
LAFW1JAAs4sSgf4tjfHFVlydc4L7o8QEfkGLyDwE8lXPeNdkTY+zTcb+l+kywppR
w8Q857+pXsGsFpRGlO4EXFvlZhwWVE5ddVv8XiDZdAkhuAlwGV+alB/c2QD+Jzqb
7wVphLOiYAH7uA9pD07uJPcmYKJkIBVLDmDdHaKIRYzAIobBQmVs0VOQS+V2dm8k
jkriAzrcu/QB2KhNb/G3gZHDNhE+7ss1URiMX7o3a1eQiijq8WH/nbgc81DGfxJd
Y3cHFE0vI6eirs4L1XdQAiDLu6S+140NwR6bKj1DylgSR64Fsw9V0Tplswd4b6x+
nPuGqtmuN18pxl8yNV6lsCvRS+JDF6O/kH+9INbV394hUsRRER+15GmrVn0Ijuzk
Ou4sH76XXk38BMhEXpddv6B1j0V4XXCOOlpezfXETQjeQ+4hl/K0ir/tNz2GXTwz
0QlyzvTNVlLCu939dO8KHOoiEvxEG27JaOFQb7p0EyPokLBdLLtfl+/MQdD5M3A4
Pa6zErENIjD5+mWWN73YeVbGiPVN1XNqy2fkRlcpLncQr58o+uX06ypr+IYHbXeS
hq73/JG6dsIt3pBVyFmSFBfjWWlaGXZLdGEHPcFnaVdYVCa42RcPjp+RBUs6VIdC
kj+Dyti/2FJeAKb8e+vqcCsiUgPfDqZPTePKG8HwCBFit/dkbtaMJULuq6Ck9T+U
4xGEI7VNxN1byboalwX9WQlWztyjrctFxIalwAM3L1WnM6IM661jDRxeCoSkAVyQ
HoB5pleFGj4SZK2W0OMI4vjP5UpjqP37E14jzrmXuUJBu8gQ5zvj4HPAY/dzUtcU
RPnX+6az/jhNherwo2bCuHIhKmy4OfKsLJ17caXBUp1IiKUfGUBU7OkyA5K6PL1Q
QhUKc0MyyKhX8n0VfolmAHfLS3weHxk5NLVFkM6mm3gIVStNbSuD4AnJIub+BAxq
SYRWfnOBzRfy5s9+pZkrsTFZzPfyV1Pj4LDcYTuv1zNNamCs6pvSFFSBYPhHRoZj
c5FWsxJFhdHgP4K5hs/rWgUZZR+79rpbG9f5UNwo89UJ3q61mxBsTQIp6zZqM34U
aW1i6XTiN7ywzL2qSrIHt3AlOuqMrxUgdpP8iSXWCcZin9E0i5VQxL8MzPeWK1FJ
l0m9c7PT4T1ptUWgMaZ0UEPLgn0hfPmWqpfA5l2ZMaU5l4YD6LXuHpn8OFPKvTxt
dRmis1+V0fc60x96NbvKwZ6QvAK2SPxq9yr1xlkzdBCN7KjxjbMlONqte85UmdJN
ZTC7TYDJEQEYefkc74JVlreBDmmx2UVXSZ7jTm9t8R33pGQ6bIicemu9gyH7W9+b
CwpyNvbTKIMzYT3XsLNmZsNT2YeHFMW7xP7o2iHqF6pDN5mPPP8YELeE2Z8PRAdb
5g0clfDeUjTo6vrvq+tvp2RnO6dinwmiOEM494Cf/B6k8eceMeBRs6UxVHp+QbIK
y5fJ4McDkaUhY51oXYAdbD0rGzH/LVHa/9nF+hyC1QtJWgmCvvV2RnlNXYeONcXc
3GV1XR05rfJk2hU84IO66HgvILnx8fTYg90fE8vu7i8xX/cOUv8RzJ0txX3f0z0+
dgWrjiHcn80H2PtfTS7ifQlXuZ2GbX9ZVMQb5pq8Fn3/s5zZ3QbJTO59glaCWfEh
sUBWqevD9jH/s82pC3ifND8BbJBOI+V08/nIBlcg8sG+bWeoi5lclHNfLlSn1JL6
vmiNxHmgNNb+NSUSpyz5DLCw6g3bIYfNlEiHM08LA/vlKXrUYXA1rE4go1CyoBc+
rAHi3249IkpWsow7UTu/oXCLXtxGmP32z+1heKbO5nqxt6X+J0HShG+FyCScOJb8
3+/4Q8lJMYFppsA8O2dkNTlenHeEp0dArOTmZTjqu5K0A1t99HypNUNfNKxlkl3z
pDXcBqt+l7ONYtZcDrSUs5Oqv3ZqkfcI/XHPUE6vhlH1pFX1Hzl0tLaQ7D5AHqWy
ctFuO1Zmo61ApigYNjo83bRicrCduIF+m/RkdvchcDspSII1HZZ5ehvXuYtnHZw0
ePnWrvwFuU7UYyCpUpeSGdp7kw4GX2fryGMUS4r518HBPYMQn3pRF3GCUAq7inf0
G9YfzPKwc1jR4vu0usYRtfA4aiyoV3xtCmxTHYx8KF9JCHT7JY2lSsbZjUO3JLlO
WanRKhGc9ruOaicgbnEvJSYxF5YDMJMuJcpAebilt7KcuARiXy1cJsg+7ZQA6vQT
RNRmlBzGJ2jrwr7ZucPJorrKII3Ptarh9dwYTsa+cSg8iPi2HJy4JEkb1OJDwVL7
3sgbexlpwMYj0UZNj0RrmG52T57qbSMAOUYh5YxHv81e0x8UFjkgqhzzydcA9a9F
DoMLBxlibK2PbaJ0L6V9hzvYItmz68MZbq64fowSam180TuzxdN/lG76FJk7A8Bj
H8eeSHDsS/vJGXIwFculNd13SevmIF1ki3mz+cDX+JMklil4cpRRwEUpmW94U1qK
P1cZoqhPflGwRNIX9wVttJW2Vt/fMU962QxxNIdTR+EselQa5ZPiXEhRzebXE8P0
zBfTei3dem+TIOIqC0To5NU71YufQZd9AX2tFKOp56Uj2Azc5Egix0yyLG35305p
+5wPcRNpp+60agEDLapgEXkgUfY8R9COJQLFulJr5/8HEpyZhj8MdHeCK6NWl3MI
ZC9mJq7AQXir3f49Pfoh3RMa/Dk5F/IhqVfGH9QrYGpCQFeUNbSY3Cv1pndWlDTJ
DspZf4oeiKZ3+LNWpcrj2YGTdz4CC35QlttDIsYg0bZvomBdKWs8+cHfTqxOumqX
95LCL6L8TcatZgsxTtRShzcchq2nD16+XoXCigHKUxO8rrch+n6e+52mpeoFg/Ih
/9OSEjPO1vpbZLW6Zrh0+5BsBlUqEonpAYnRNTGAqkUtulMF861rK6UkIuiyg5TR
BhcPAvwG1LXi4rZFwKtSU4lroVTZRptYfruwIQTGJR2S5Ld+PHp0Wrl5oijTLPYn
Y4vnu7viNC5vLJjTyZ6oJaVxHa42DP2xu8g59RZZI6os1kBqwr81AoJa377RS53y
cQGZznf/YZ5j1MfS6FaNwqUCdi4H/QVBMAPNbpOt2eZBOEQeBxXE8jkCzm0l9HWd
alafkfaTEG3+fen7mFKO5SKd5yzlz4/LvQy10UeMjfTsJ+3Voq08WcWOCTr+FhE8
QBBD7bL8xRQpYr1sK0vKb9ZgUXCBPiEIhWxYgeRMyTOLH0F5Gnr0fCZs8yapCudL
qz6oEor9tyDJBkMAQVZS/MuQlnWcftkJznoI1BFwGRIjwAtAeHGAFbuqtvNlYQpe
RzCXRrAQoVv7V9rDGcNLVNtbapoeOp4a7mPlA1mTOp2l5P3oMKSgIUhxFJqQz+nn
wbwRpukq99dlK5xfQ0A5xlBr75rfOvfh4Vtqmh/0wHL2lHUTrScqpb+x06gaJ+y1
XV3EsGAg1zNhHU1ZTKQqsRW8ugcgr8EhSz/4fsMUwheD83RfmcQzwCHcQ+lr+ihn
Naq97JBd5yT2eXdyvA/dZq+sbvk5JicvgHH6gfq3txqE0zSCCmKkZCsCy4dPfPE9
m0M+KddubZ6J2yy5tb0UFBYdAhl+AkR8ygP5V4pUppk7W6su0Lqo63nc+lswEDR6
Hj//Bk3RWlmBHQhKZyVD21u6Uam8yS2JeLsjZrwhAg4JG1lPQMZkX1Rksy65rmAG
HwrWL+hm+M8UiCZfFHoO1phyLu9OWZv0lgmSaHs583o0QJDx+CKhSoKlK+q+/Jgh
h/1VhO+8RNyR4RIrt5spUtqulNutb32TJ3lpDieFVY91oKXobJcxc4ygCkaRodgh
dB3Ue9Gl5JgjB20Aq1W5bMw+CBJSjtcDliMiv4Fjbedxlyg932DEfbZwg69k1ndA
H831VKoFYN6BE9/rIuF61yXxDsyQo7wAmRGN4aeb4/VAXbWoarVMyLLLQ8/2eJHA
otPwWpxEkDOdqq498H3/T5mQEhvzobdr7Me/XhG9i3hkSZnXWadUO6+aDBJGH9y/
UNmH++assMO0Cp2K3H8tk5GFItK+fGDPuerE3MKAIg5nmea/rXV2mdS89t0D66nf
2YaPXFNnt9rQkpmSOcv+7xkC6p/Dna8I5+sUxKA17tOKJf32VUDuUOmohaDGloEb
VVdFcgVJRyS6uW2MI0Ju7rNZx68Zarlt3h99l4ksanithUISLVPDycF5JJbACC7P
gon3R9iy5eNyT2iGAY3judarn8LnC2gZuZAtqeP1oYwzgRT3d/h5OiXbvtK+wmOX
p897gqkPrZR2mjH1QECaiIKzseqGLW1IFAW7Hdv/1u8N5XJBtSGwvUkO+0A6s3Rf
tgATE2quMHznXJu+93FBYkuCR4iFRN3epERHYc8x1hFaZsbiAfq34A1fXUdUnrrF
fKr+qWuA46xtT8OOg558mGCPCgb63EuKi8RpM21qXMOV02qsepqwEfR6hNAQNQzD
MsPnCpfgnKaxq4gSMDUAGtPCkT6e65vphnGSLsf46asQ9OgaIlfshaTBYAtxg5vU
Y1Q13WpJl9IrV2V7bLNJKmIBO33OzjWzODYfNKY6QA8Icd/x7y8XcoqyLxGIO1/V
4rkY/zNe2vhaI7mIs7YwRSotzuh5Sd5Qedufha50UViN1MzmfJrq+mjj2HCUt47x
G8lMp/R3NVRWWcEU8TPX+TndvKVucoGw2pGNfWDJTsAXfHAJBTHbsrqC4sJHN7Fb
guP/mkVr8cGo4JSztvYBNfiVllGUKAqtiF0hwUkMC7kGpVqyXw7u1spqUHaLhW5k
uw491VE1tG0Gd0OCyqFxsP4dSfb83WdPAjIKy10U9vCGRFtTHG+vUmgLc5thWIku
epBOua5MKaBmB+Pm/2IbyikIRrS6TrZ53mwAc2vG/hL3ODhwkFPF58yXu9u74UnL
rybkXY1xYTiKwDYnFdZ0h9edllJlFI2TMXXcmvG9If1St9CNs/GMBzNABu48gRUg
2R2C3xeI7Ofc2bSd2yyIG3ajppt9Vw+C7de6XX7lMuYgowvuZQ+uNmdHqp+0t0Ab
5Nx+NzspiE4OuyJyfjzzbOsEFgjBQ6vhV6gZoQ2y6XKHpr6FLy12mDCnDEKCiy02
mDAch45ZFrIXWcwgzr7iPKhnjHivE6or7yYHyGg+KyR/LqMUGxcY/xZvN84KOrmU
o/NJ8hKLhz15u1knROOzp6jX3c8v3DylyBfwduPgZfYXf2HK4GPazPp9PbxmaIkC
Y2OMLM6chJG5tJcvNpIKku5eyqg1GG47Asuu5bSwYfPEJPRua7VwrI9V3vWvMu9u
r7BL8DzKw3bpqJ5jeNO2VPIiv/iIkWHD1MO9d69vsZZGk2I8kqY813Jtf1+Q9qhL
BAgld88830vmPcfCLRstm3FWwCVaDAGhxBHHDqWHdhpytj9LoL3UgPosteTfpMKI
3WjMPb+x5jL1Br9tVvn86+jX/QCNdKCFSH7fV+Ibc3J05lQ5P0CJghgaJFlQhf/z
Itm3jJPSLQFljMKSuq8xc6XnaoOMWhtOuHfvpejqLSfjoyo+3M9Y7R9pzlO1HkaC
MxvAIU7l6cajOCJPotwVGM6L2oUhTyxfzFD/JQ+S/WgRfp8xRXsVZHWUAFPAWhvr
slqarTaFzXy+91LgAQFxZ+eMLYpkN/gADOmWoklpMgC/91DF+HQ+mdqsH/iHexfU
2Ee5uA5G6N4l/+/c+FPov1Ocr127NDV1uf5dYKLK2edUDksx6wvzsS0/Mk69b2rf
lprDu2hK7NrrNC0SiJ0aE/nnw7v/zSwYxoV1sazuzPSCP5PG/4YzyahEt3YsU0Oh
lmRDcgGw+SKo3cPFsaSpdamzkV1lJw45XYCAMkFnYpI70Jyg62UbdFf2E0iz9f8S
1ZTv0eHfgXLGkWel3eI6/kJereZwd0QCmalvLXK1Ipp615jyehpIlw2buZ6QHgDG
A/9Cd8oQcYrVnZzBHOlh0MycLPCN5ws2ogLHewkWoRD+48FOxDecMalv+fkd+TlD
Gf4tZtpb22y4Fep/y4Q83O2PNHK3VaxUjUWcQUp9EezHLXaNMjhRslz+kLXR0tZ6
PwtQUmHZL7l54OYwl5Lj861tdM4GlPuY78L0jW+h6VZ78YsEs1yxjJ5kmn46X/jr
b/0i8W5EH3unB5KFr/ay4lpRen2dg+iN+WditT+SIWR1fXGRX5iKhjlp5ngtikC/
GCoMbQx5T7bsA8xQMhUkauRQGqmgW8Ty3bh1kzFUENfCgf0T0KSZGuFupsbKd9mQ
kje/Ms+3/yhrN9+TDKEeg8p8axNczt87tmaBWABZF4kHny0alZOB9R8Brcx+xRE3
EBNw/kqBOlSYopcnU6CoyDWQaA+SUsEN4sAz4SO0smpKgA9nCtHWXYgr7TR0gkpC
+Ap3wIeRCiHdjO3lId2sY5916vj7/l26aeF0cIRZ4uIIwmldKuKzQPua4xecuKDY
YUFaWd4be3xh7gUjVYsTzJSzuk7YSi3PBAkzJ+9xbvovbHiDyM9oUwVQW3hw1V9Q
c+lxykvijzJVSn1Ng6XLjv2CPjKKNBL6wat0JBLqt6AIdorMm5Ac8K70fTiKUzDs
46Ihw2a/WbI/VzNaZC/3TZLok2CicHZAoMMDhGJXY217TZZLhVUyubULmcG5D2gC
qBxlAln+KCPuiAQxJEQLwpv9Ru4pGBHI4B/Lqa8b9FCM9iIe3P0TZLXOpaB6XhNh
6rEQDkqTbpkb4kU4qOaOmoyEB4aoUJVahKxICmATCkVi4w4GesKHzq6yN98mhZJH
pw2ZOzsb1el72VEAFVNrJdfq9vbzE8tOGa3WbsmH3oMRY97LfrJOzblYhADvOwza
8/1SdTex2uVAKIcaFnQPzvP0jwZlYi7hA5iRih3o17431pJUQW0du8f+m7/vHVdJ
sGm0VziHGxbaL4QxztNvXT7LP3s8f7zQu6GaYSinJVmHekI2mtlbNqIIN1P7Vq/h
F7L9WJ57rttde67gJKQHsl/j6uAZGqXfeCEEISWnhcxs8moxDGqXI0M+uOWuZ+RH
HmNI2txytob/gsnechF4HwU/oP377EkvLAV3Y7qkzYR4Nz0+eWSA0haGV0rT4cx3
hakOR8lPO/0imCtgf31zi3fowz3LguPhX2VpGRORzFvw2LXR/bHkuqvR63ZgIN1R
ue5PMvNeOAI60Qq+7eRsdjarMoRcNBydYMDsM+EaSG2VZu2dFgaiB8CBqiJ35JtO
XyrfJaZ04nY8vv4cKqoP8NJ0s94AriQ94yewpGCXB4Rp8xrGSZd6q4w9zvR58ltf
LgEm342JbKxEiq1nWRC6RvzPzd8TMga5we3LFFy0Zq8l1TmPkvWeWm+N7bgiro7w
ufZe/2QQOR2JEwDvbXGZ6coVM1Qul0RL/jZqHPGK9XhdC8FunepnoMxtbFSmIg+u
cBHQECelO+TaRHUP+EDAggPDcUXDmdGzn+3lD2QHhYtcH58GjQqMDv/WWVK+92KX
vXbV0nBiz4Y9jThIckhFgNwIp0n0SvYfTzNgtPgJgDn+TcZjETw0aJfqzqbvZARV
L7KMqobYFmd0EwzM8C0ZzZERcJdbcAb1l4NN+j671MUnIvnO0j2+Yj4Ex2TcnMdr
DzOs0Tlv+gqdC5Rb96ot4vijxygD6acMcNeZRVuBNV2e5tup4yxZjVlRMjmfNPSr
d8U/DNcRgYZ173bn/iKXYCG3v/3PUi8/zEyXYn2PkfESLNcjb76NkbPHwqqU6B/x
TS8hBXiqgZMrPHXgpcV/CFiFbr3X+2Y9VAQGDs6pFIDB4ieVhbmBskOBIw/qO1Jw
HeVqsufltmhiNiScp22E+hATnTjygMEzDBcNNwuqZj94WQKVqeick7U6HCIHPwrQ
JOS3tAZi8CqgAXn1+1K29itmTVgzlfvEtd+VfFKOu75PIrxQKMQwQ0QTJP6M52oB
/I6IhM/yXMrErs1UJZ0i+IYhy/JC3zXbpss2iuh5+eaHgmemQpHlXRBULLqNA44G
r7sjGOudGuX6oeuUegbN5HhfxQd2U9Ok73ePnxsSsdTsPkg5TYQKzv6xd7nJbA/z
CmlcDaE8IpOfcD0GBFAQqNp2xfoX51P8d87XkBBcK4xXM2IOJt60i1NP5EuTwuRA
pT7PGUFPnIPlX3beSL/e7JsuUR9OqMnHxq2cSj7bz8Q1b1lSfG+tZeLfGZjb28Uc
lSIc3JQGUTa693VeDBELG8lt9ui4qvtZtfJ/mwfQRs6ZWVs3ycNCzO91AlNrrvob
ul+naXnUT4/NMxg3i34kKBl6J2tTz+475ATvy8w78Iaxb6F9ibioBEy17p42tSGK
GyQEV+Q3QksMeHsQMfBnaUSaay3WqG+ABySNRbz4/ZJkINY0PwWF2Jub0R2cRaNb
Ti2Rk02Fd39IjN83iq1+WH2B36AGZychVN6cKwt8V02KTfQoZGxd1fcRvnYHSxr6
nXU3TDBkoesKcirjYHQGOoWH7/SYffyRGUEDsH7kanUuuybLlbYpSXUdwRpZs36r
TEE6AsrJLLAcka+/tatn9BlQfP35bGRACWRzEfnN5QoCtWdNSHqnZQSPOav01PTt
DrJiKRa9cWzW1a0l4gIpAy4tj2Z65LF/HUdbD7A0ZXpkSp1P8uAdSWbQdwYoG4Jy
xE/F9qamnkjM7X5X8K9LOAG2fOIT0PyVuW6aDCKRvRJMMy3Qd78uSQ/NevGdKug/
pJ4nsZbq07F/WA/DM+ZKqzn/lkh0wkXjmIa9kEXYPizsP+sc99fTNfORiffTRYcj
4JdXHraNTgS/9iJI2BYC+zcPJq+IP2sgj98p+RM5FKWtgZOJSed93SRRjdBT/oKp
j1IdCO1qiinrvLYjjNviW8z5Pv0Vs8CR1oi7d9XyZpQx8vGsDyl/PwRehVEqZvcb
tHjk2PxDykzHgRKew8K8NcvEIOaSFAHpkTuJtQ5n05dK3/fRS2d7WHeR4SNEJ1Pm
jYrA5fKIsh7ZgnoGeDL+F8tjNGowH/LSUYSrcgFyT1Af4dB6hM1sTPJHLvHizr+W
P+xH/GB5465/2w/zqOpx8fNmkKtMTfZM8qkE1oLjduMkXfxBtwFAEGLCeffQgb16
o4Cdgp3R50pSQ3dQf8okwgC+YFilQ2cDWb58BTomLdYt0eDRqRVyuGbTWZ/O7IuF
i5ZgCFMxNQjhm/F4K4fuD/VHbm5MBFcOgoKWQaCffSL7cnSAJS4uvD/pKI5vDOe2
086hJG5TH/2Z06IBwS0ol60ryCg62U497DpepMlA/GQXGoM7ockTximcNKYkWRke
YxcyQN9WJRDFDvqNdbGx+as7/nTm+ncs5a6ih0oS9lvSlhsVKvXV31q42q4JbpQg
lQNnJg9BBlvV7SsVlOZAWkc2yoTtGg3Tu2nX3lgLXE/QaGzUxzJzxhedtqt1suCu
hEOI98rhQhSVC7RRZw8wnh9LvCuAS7wETbpylY/OqN2Ji3P60hFnFIc305DfJtmo
/sG7alOikh5WOodWtR+Q+NW2DFtye01ITC1xmIM48+tstFP0NgyWxlXCVbQ6i5CC
PJqJCaTXcHqMJXq869SqImIi7loX8L0pHZ+TjjP8DgbHjdBBoPZqYcF4xhx0d34R
aKtixb3kYroaK1lb58eQnIWxPbIkuirs50/ea2eK/DNxffB2aZ+qsmURlQNMzcDN
Mk3mar9fp+4S2v0ljaW/OIMC0HgD42YgmcWdJiad7+he0UjH8jCk4isfuTt6+kHp
9GubQJgCB6G6PtLI5vQyBnLdx8K2LQH+JHuNt6FGWczb8J1FNoVgsWJTCKyHFsc7
Hq5pnw78orY3R4koLRFCD99AHpTFvxWgats0qn/HXW4PhOAO2rbaJwOt9/eYP4hf
uv01Ay4dytPbGZWp7bq2A3Fke8Md8W+aB2OyP65p9eNi6r21V9i+gxe3C0GH4jW0
qgT886S2m/GQQjM+6hjJkI8y8wGUWowBp9Vyvpo5+eZPUjv4PAqeLN7xed6mwiCA
hmwyk8jpKHM40aDtza0DMtQ8TAJYGD/Y5xbfxzjj6A+MZfNPwKaypPMHga0UBnPl
hKt2xQyAgSvilqlCP/LUUQADZ+YXXRQY40Tswq21YS1B0Zyy8C87JihOvwQjNLJ0
1vYDDGoCsP8tisJx1K6QkPh2v5sg+i9FipJxywamR3ciJTw5u/04X/qf4HS1CLLd
HDjKLAZotxEOmhy4/vQmN8o4/Ekvi5RvLhqW3HVIeKlYpcCWZZpGYW9tISRMxdPC
7nccKfL03dJag5mwdreGWTmANoq76XxayVBwsNQcyWMfwH3vLtko2zLbFJ5yGhR6
MhOCZH28TmLtRSQ664vE92MBy+ewcmzqwChJMHxaV/cfXVlEncFzrFrNX1Y+0rlJ
TtLP5QkBui6wH/K+8emJLElATq3e2dinOEEfH0+EO3YUfgRFjSO7ouYk51P7sLCs
oL+X9mPw3wzyIdfkRA4O7OMxvW7+sGJ65yEEQPO2gGDr83YGNximM5rtaMaqTBWi
CpPhNL1q9lvxyBUdmTXVwI6pxpkf+E4rt3C1lokK+l9tdwGhZb0/rf6rEHW7dYX8
xEdOzJ2TUQ0t0q/qYGdwg/IXuPV3pv6cvFKdLwZkk2ns0zkrLEssnf0Wm/ILadTE
K1GOU8pE9aJHizUJ6ioN5mpIaFoU06a5fvgEVxTTYFzATd+lDpwewPMpLPBxw2uR
t0+tE/TQ/F4wYY6Ij1Fpn6b37jksHiEGIuXkKkC6AXkgKUGdq3PRZgk0+kJiCq7D
4gSWa8mXpnXtxLrDKAL6ukgwaZGJJiKQ5y9+P+elY0bjKxFGqV+e6E57imgy+xUl
kOWj/IgZT9HvmAdJTQzyJf5xCJ21GHxCJ/NTbr/QGp+kAkNmlJaKDIN0VTXF270q
l1QFfmmRBcUPqSttBx5isKFyXzjSnFeqT159oD9rnbLSsDcRigW6/8FZOxMaJEez
+Goii+tQKAOyVKLhlwkTLZApXvzXplgihG9rv1WeQCo0mb+17WeLEH2GT6hSt2gK
Zz0Oo8UflDpP3oXmfuglfW/g9RELrypyN+LO6B2ClPkgXlBIvKiIx1oV3tf/NWTB
mkv6JqlNQNZz3SxgIUmICgtGfkURkkbpWBaSCu83wNaKCMPjbix3oRXr+MFHnyQv
znhBq2bKmQ4+q13rHdR1krwTGNMB+zjKP22sqrDqx9V0h98cNIYuLhIBhA7hxKuB
Z9iA7e2TbB3VugDnK/bcW6qW4xMCkL1sH7KGVlhNyagz3WpQXwplPbcLgIJ+CaV8
eJhyokn50xP1E5QH+xG5UdGK8qabkFEElsbmti4flHfbJv+u538M5u9V4i2pjFmu
OoyGqPCitRBarZCoXDF5rakKMwM+U9R0H3BtrWYy/37Ob0w9T0NmbkzxhkdYgUfJ
A9ZUfqV2ntueyYNspfnrfE1PxWnLOaozPFxmiSNJn2ik542qR0sQqoxYipPwGcsd
TRnMppRbHztEJ5EdoPL/R5K1kSjWaFvOdiCxZ5pR75t1zyuVLQzpUr95G66xy0Z8
Qs3KlXyAZH0hjg2Coz7yelDA4lMEP178v0yRNMAxJgTze0b21JXZFGFOtXyOJiyq
rp+VurSL3RURE3zbwml7Wl1woRTvDTZCqnjHXM8eG0KX/IujmcWI/dAx+VNLyUCv
dJuGyyTZWP5SxGZFxkJXUHZJK9HovoqkgFtoNdyMGUBpuZQjwWmvDuDTQ+3858Bp
+Gh9GN3dvp4Lhs7KsmO2bH/2xT9seb9LW9DN3wen78q0lRL36Ano5rTT9ACvPoG2
W8U2gcy/exgWJjQr+1sJniVqh/ynb0hiJ5YIL8Lc1o1jXwPD+muOOAmWQ0WA11h8
kG/OklFYrmW0fEL/PFMX/cdQYK+8FdbpTrDPyRJHqZkIDQ47HGKNcw0KcgjkojJt
5trj/o0MXeFdnwYG1G/ilpOB5QiH11NIvqqs9q/1oPs+whjvWqDtmw1RAwJvToQT
4RdPjh57zzw2XuFCtY/L2FmmLVwYbXYZ2C/cj76i6yrilorB549EQ0qZ7GCyZmk0
cWpZ3rnKhq/GmA7XETP2FjeVcXSQ+AoYMjneW7N8DCS6JcdfnRX7umSS3ZwBxUfu
ji974Vau6k3z0NEEPD/QMtfVS2+m0w98Bc4iTmic48X1pMtpqCn9XSLXTVPi+iLo
i6cGoDgo0G0Fk7rYVpOeQ5HEmIGfloh2KsE7Xu1g7xTa1TybBmkgBAEZEJ7ScRjm
BPGAjfStDyT1a9witpI04dksRbieUM9TCwSCZzeGM+fy9YW3EiPPfWALGMtpyQkt
LIeBXskmArQb0kvwb/66kv8iv7A+pXeDTNYnhSIg55dfegbcZdI9U/bgaa5s9h8X
0/OMKetmN5vUMfV84Gtw4X8tC8AmhystbHDL9kmGHUYxK0czAiliThNqIp8ItcMD
WmDTGE5X/mvAUpnjbCjBU/ufKaMp9eG1FZRD5dZ0qZ8JcQvY/11o2f/zJW8R9pip
6JQVaaDDHEpZ8kAYIxsHLFZHhDMTBtvUlN78OxcfkaQpPGQRW0xQS2dZD+5jc2Xn
VVHZW4y9qBrt3FEcKqv6lMn0EkBdR5qxPtlxSmCMCh2BIWhv3ZbRf21PQn6NuPPr
K4fMM9q45PFAXh39Ya/utT7cJqd3K1+NJi16xLsWKhqhkxx2YkgBFxejGtFJNhwW
U1vs5cMd7OduA/qBHhFc6VAV96vklw88PaW+bdsb0ad4z4/XvcY5cZmt6TIEfd/5
AA4j/CrsTEaD4YAmkv32ObtTYMPg0rByMXRgXN9YWHRUUOP9LOuULbcgddlbKh7q
XMVRrt+FjglBdXwa26EM45oZs9uiEMCifsc5rp/hPTwxz5fF3GlQOew4VHIx+1GT
Ahw27PPm1nnvHLSmzUB1nHyZfpcORlCURPyPUodX+i6HsmA3/hUdcXPaOuUn9IZZ
WxigTfz9NHy/bKikeVGY1JRZzeIE1ib2DXun0H9Xt4nOAhQz9ZPyX8t6aPNkYuVw
aWu9eLsoy8JN1qZi7KJe50o1Q5m7i087wv4QZNscN8Hv6882i/Emsjy8lOIOKusu
vuhadN6LvnWfW0ZUZKLbZLOoW2z5NEPgsl+bC9bXdLHIvXT3sEVrwfGeC93n/QOw
SmSNMMKfEFacLvymO26EAwP5uuZpotBokZsqEMw5XZfG81y/hznZH990mnyHPDpp
urn/Mlv1SAvhQXPCVH3YCvRYq73RA8lTHxkuOUUokSYFuAcERkXvTmPWkUR9dRux
7tZn9cFJXD29TSzC+P8G8bkX4dTbghCHXCAVDXyLNOkhuleowJDNNYf/2pJAs4Fb
A/qq2kZmtetZGeTacn+Y7DPAXX4SxKC5ZNBsUbtRbHw123l7eg+Ab2nx3VJKkM3t
XsupkUtc2Aughdu4wWUU8eQQXdwwLh4ZMa1/hDcr5B6sC1pVVRxyBFbJ6zXNG6bY
RKDFuZAFFGA5q6KpwSrhhicUOA+/TPIu1kDv5B2jPnKzJP6ceheYQRfIorp/YT49
EeJNvzZB6CGrhBcuEin+aSCLvkvEwzsjiqCx0wTf9yFeKU1tBhbufyIC0K84mx9g
QDkvcohcW8ncFZ14BvmffACIuSCkMNWfSojFx37zWY3StsFeksaMuj2/8MsBioZ2
aHVrmia8Pr3cCcVUQBHBUgv7YrPGXtIPhyG9Ec3FrgkfsKR4XznP609gvDU+xWeP
je4mC4wA81Zsr0+F3W3FcF5Za1zNk4hZ0AtyI8zxYGAEVbbyGtzKz7Dvgq8yVYXW
DQ3WznW4/Q/hHv3aWs7Vha2So5Y7lNtM6zCp36q7jwCITZYcS3KyEKuLwg1zsrSg
1oDtsASyywTlpCuUBD+8Xmx2D8I8U0YSAH72EgEVXS9WybDqob+IvHXh6WcbXas2
QEuSVylAW+q89Ab/1Qzxd7VEpCAMLfxKKAE/jbGIU2Ih5NqYHWhsC0KnJdiIZ+Fx
+rib5xPnouxRcub3h70eVq8l0EG0jff41I9nYKpShsOI6/36ohpnEfOqjgjGBL/d
RDPFh+DUqvH4Yi9bTxVCn4ndR0gTTFTvCBHKxiJzVJC5bljLgi69841aBM4gt2u+
eTxV0M2yv8jAB3av2At7JJA9dEsuEXnODammGSZLzo9mAbLqzFmgDMeeTCanmyC3
+FMRCLxsqEMYrFs5+m2MP9Y5KzXkFaXpTDMaU/6J+vUUSl693Zl/8qFIK4+Wq4OC
qCOljWTLbpMC+7GRJbV3S1WkDiKiD/i3GaFL1BfVcS4Xv8hesqsrcbpgH1njqgJb
87/ADgx7o3E77optbyyfI/JzYJ3OoW6IvYX9XFwtjRYXnhX6JmkOEAjRqLvwzqtP
Z6z4Sy3UWmHuRBoF8ltxMG67FvJbhMFiN5Ebl2JIu1DE0dG7jFbZaehrRanQA/Vi
JoPJPU8OplNulju+WWDry4iPw/cUgN7RnBccL+zePI9YvgukCgAdI0zqgDYG1T0I
ud+CSG4b5SKFcOyjXhRem1SnofzOEKeCzmmlxZzKVvmclQ93qbkFLa32FgWmvZIx
TC5eHHrKtzvGb9V00du4npThoDH/zgEuXyCfZlsh/8+F9oGY6W6x9T5EIzHjY0Cn
imhqfcBDRhfPp3j44XYHf6SrRdUYX08UQnd167Fu0m2JdDXVoEJrVtLMu6YCnGiX
2CrrG3AKMxtAOejmf/PAAR9MMkgu5WlFwvbYXqKBwuYA+hqNlAF06CKp9opx95ON
hOsgNpYx8h8c5EzimWb4l0swXeKQdORd4J8WR789Vbp71NSxOeR7K7gR7XFfQhy3
9RyEClZpuwxjQWtESjWY7gbc6ggXRBZGzpT5EWhsdVE4KGWswxDa0bMbuHble9d4
o2o7ECj2carqRLANeFgDHfJBWaoauUdrtjsM6chtj53U3TEhmVz0sFz2o7JWuS+i
BsWdyJteXM++bMyW8Pdy/05NLyIFdCaTc6i9Zo1gIzwGKxHI3ht9V3rtMsPn2Xez
CD5yTof4SHqS23TY0E0GZTAWEhkbPCMDdWUFPGPF9lbPAUFU8UCJ3N1FzVMenQJg
kJSblfbxe8iVUtwTaFmyPbpSJvCCwoQivI0+93sxOYRFgL8BUVxyJ8MS6D7tbNcO
LCmHkOlHeIzMCg9apFqMBYCHgTHOToQ3h5SloWm5HnBERJFGb+ElQCiGc1scl4Vj
tVJk4vv21z7gACyDDLG0J3CioAD4FEPJN7w2nXYmgV9uQTf8BPqI1iHEorbmXvmP
UGkyTNdI+7yrUqIotfDyMpkfBsX1TKcDwEenTVB3os1jvpMOvgCgU9ou9y0q69NP
Bs0PA2niuLWainISpYVowSMDPRiu7Yq6ROegdYuO31JPrpzWm9MxmGvi0xa93Ygn
C+6tfrBjK3FR7tUBzC2G3GYb6+P19bxXS3WaW2G5QjCyI0hI1CPcMIlXiGP5Vuar
wHIbRYPOm/Lxh7BNttaH8RccCjosiY0l04uKXiWwFbeZcH1q2STQ+/SjxK1e96Vj
i1Q1Y1rxgqbev0I4Q9mvLHLfAm8wV4dmppMMOLGTIfWJDBaaAWFH177u7fU9eiG8
HF4X6RrTrHkQXST7OgrimdHtHUEqEZB+LLGZL+UkZo4EXhAgQIjZ69Fg6jzsK9hK
+pQtZTR3MJkAdTo+h1iH34hyzjElTCFjci77qQb5cGo4v39DlSWbKoI5HsFcqcu1
FvRvn64K+ewOJDCF9gWJHf4mLh9n4uvJ1QFBpMk3PjPiZpHxEhU7wtRfKtomUx4s
NpX5vh+EZssms3f/7RixhZfkBPjZekMfuBBrAdFsJR+k1qQTcuvcYNKYOt/HiWVx
PWegLe7RfOM9WmRaVU3UkoydVEY7wx3p2Q1g2Wvq3WDMI2evG0upE5y8e6u6koVX
mygq74mO9vQWDLDIS3LMUOEUWUCi8ja9qANJeFqoDXVSZ+QeOsRXnBwvBkCAKQJh
xxd5LSu2mmMC1Yk7cx9E3tREtpYgFAKGS0kG74GYSNtNqQyrQ4MVoimKOyydYFow
Owzq+XvQvSnSlwYsfV5kDW24LA5HyVG5pv2YyE/e0r0BF0m7SpwIHpOCwsn2xi/c
PF9r5jF4nJCdHt53Mv227kO6Jh+1JPgTqrQMKixhdkpZ0LZJzlGcQ9NObqWTKybj
9gPXQstEGYu1JvFte2xvelIHEoS7pEhIbZgcPic0tjURyVphRNT4cSGhF+umWHCb
RfyfVUDI7xZ9rrf/cpfeuam3udkmL1ESwvkp/d4vebgDB8/lfRxxzCbyW/KAUT1B
lxjewLXSfNzPecZ87+TeH82OGZT2w5l52IlkjP8JZYogLafU96q/UNH0x69JM3+q
qhm49JQvOJ5map226uaZYb9gu5H1IwLSVH75xMU9vOhNdl2ZQQTgpf3YXEhFO1d4
4hZ9YT3AX3riqmoLXjd7A0hhiuraSZLyvNpZlaRTf54CAouEhJa/2tz+FGFaoCXb
sMHO7rmMU1vmTuVnDZimxOSSod6L6K/wugU/j1I+D0SaVVNWgrxdJ8wB7JAsl3h2
l78ZfoJutgb44ys33kS+RFifdNqXQCwICCguDGpCsM0TG+jLLY1QLOcmahTfH5ob
njPPRelpzYcxBm0yUnXrCbzeGsRqFzk7zWUL+UKXRm6la4ty1vwMETLnELHZw67p
f3aoo+NKcrDkslvD2rKYc5xmyMxYjfz65zwjQ39ZDO/x6a8AwzNZ32RmVjDgo97F
Kd2GOkvYAnP3VCFMOeM1oZRQEyTmb3/7DBcQvsDKBWayZ1Za+tjgN0gjNiLrOBZy
5bhaqcf2P7cricQdRbOiWkDO2+e/lVwL8L7xQRN4Ef9z4H7CdgKGD7SNjYnBJ0+L
0ucV0893UxVYHkKESGlorxQYYVXr/61yBfTQr1Dcxfzht6HxxOWVSewrd0dSZgau
pKRA3BacQzQ/l2RxXCQbGGHxow2jils6rY4vs60havq+IIbSzNDn9ezNaCIe0kgo
kM6w9dpX0mZ6VscF4zMnyd/cud+iTEHas9VQpCqzE6Qp80QBpksHCnjQAnpG9gmk
aLbknadJI/YFhDnSrSv5rryAGF/kDCf1rkDO2WqvTLOrnjLp2QBQ/dOXk2ZERUCU
X6MlS5CzViyvDbew2URtQ8uMmeDlSngf+huLOWrVtREfepCa30M8PVT7fwWlmM+l
cPO7SpaAPv9Lt/DYLJUSm8leeFDrRKXBzHNEVc28QDB8xmBldUnd3hLhhow/qwLu
ZkVRu1sg59o5gzi+A/fQFKU/RJSuP31wxhbLJ0O/5LndXjBZJ/J3/piG+DmeNHb7
TBfVUg1AxG435DFL5yQ637d6pPnkByg1QtqhifuImmjvfhjJN7QwAy2yGuLXMxUn
sWUeqLDbav8Xp1OxI+Xu2ohrR5c93R7nuQfnv9S0uD+9diIMYGBPrNsXj2libUvp
N+MR+j8NXPt193XtEHpq4VFWfMrfsqYMp7EM34tFCTcKAx5Nt9PsNME7S0oSGFoq
p0N/Ra6LmR81TEn54LImSOA/v/sr/hhTgNVr/+roSMP277y7NIKHy/CIgJ+eyu8Z
62QJmGZmEg0ges2T5LbuYRPt1MMk8CK8oWOXq6pVHKy9G7aqegKUocA6j6Knx07R
/eVWfOuS3/q4hktD1Izu7dzNXl/4qTqgfXte2dlyJL9UcXEIRI/HCDmw94U3LSVY
5kiVN0nMLiJMeIUlLGNgjkcliwbSUOGGrvM0MbD+quXlH8OhmGGcwPDLJbNmdK6H
KjE7lxUD+O1ExWPuGVB8RLTdAqzOpJiptxlGXksrB1VsPxwmGMljhGOpRZWLvrHy
oDqWdrSXNIgwfCxzZ8F936gfVJOQt5bpgerAhxF9bAWHfDTp41MJKOnZ8F1OGH4/
QfAu4hfUCLKqzG54wajf8Orq/d8TiTxgfmqcnybeDICbbyCDOYQ3ypo2JucPpQrj
3c9l6fIjd8tfo+2ax/HSp4mkFBAtRfetgiHvpkRpQpLVtFE/gEzdjqJs2iS48ZTO
QOaRk+UxKMuQSNeb+jzVacS58Fy1Et4GUux+J5jhuIICSxktLCr3bRF4qaN/3Gpt
aIBC6BXr4a2hvtWdGx6SFoc+YphSS/tafoRa2p+IyX2KmRRcCPjxKn+haQIy+AKL
bo3rreTrwnB3iytrL3C1fYUVGEwcL9waWxZ2NCjry2TdkywTd7UDI7vrPMKzjGUv
y4lHwH/ujWZuHXIeXud8uCjE67VXo6lCF7z3DEdIbnNaPt7+SeYucOn28OojFKIc
QULKtaMQeUq0EXU1VtEfBaZQ7TbfCe6CrZjBehv0Svq6xyA5pgSM8BEMBu987fgr
V9YoZ4goXneuFguineDIVpwMKk1nutk1zggKLGgtc7uPMdfZ6SRuK807DmLwJMxx
uy/sd0d12mLzIo3OzBzkPCpDarcfLe/sve/T6xQTDd6Ti7s3zujeVw8PfRpSgP3u
KKf9nmENJiKyjDBYmwrQLVCY03j/NlhmVnDQbGvsANX3BkyUMhCZ89gMJUqgYiQm
S/A1zGXrqB8UktmITkf9osed0BXLfCsunoSuQO5pbn7mqyrMlV7lBmwkS8f+pFun
LZifmK/pdYiUu0biUkywd1fY7gVDUBE9k8i2tfMrHzrFCU/yMFm8k4ismxpuYNQ9
4JdQkxBV5g6oXHWoLP1ZC+UzXAp0LfJbAp54NxXpYUlAKU9A1cCd/HnNrm46A+ms
EvHSfCP8nPItoLkw3nZ5aGzBSZcISMIu9qyjXx2yywXf3ArVBh7jRzx6+R2i+gQu
BI2cevbxomkkqp9cMo1KfwXRWCyL1uT0Ybjm3yM8nf4jb0jY5tmxckskQ+scqIEC
dUTn6davIqCZW1g4clIqUxw9mOOnz4S/xoMVtMeKFfKEKZ9oSoVkUJJJtw6sfK36
LKfmN1j5yidKzjxMPhAE3XQrNMq/HVrSA8Wr5EjcdV58BBT+Wwz2JWqEMY/qsBNT
Tgo0vJiENnF/MMdETBooGFOvuWJeUwhdDBfCnZYqYru91iKM5V1A7ib3wPG8RiSe
sHHHgaBe/v059U8+y+da6tlvLfQRH/x4Ihy95sBXeJbBsX9b/dvCuTVDGZui2Pa/
s49gp6d9EG1MBrIrtf2sf6q8bcaTXWpCZnnO1SaUGAry9k0gTEDc39oh8nHEk+k4
+4Id5JvDBj2WhcIC0J5b5zgrJKIeQd5DxHDoZwzFeQO+jmKOl7nwvWvYEq7ITzcv
xRaRIzi4W+TCcWTdoOT+Ynx2RPoQuNkVn0Lq/1cpk8WA80PbaGDdhnEw2a/moudU
ig833WGM1Bu0AgGkSdLDONtm4uDEiD6tujnFKatemu9eSs7gr/65CHBHlvhkmrzK
irYuQNzFw4vUNyMX8ounF4lEwe4HCureWDgCX+QA+ltFrJXgbRsdoNq2MXDvDrYS
AyUKArusyPT6m7Ov7R+49LZjNIb9I+u1Bp0O0I9tj6J59uiitl4gw6OD0tTRxgbY
pgOI4vhJ9/vNF2WdYBkCzXNcfONiyZsFkKzn5kwMfR0DzLuNOpTuNym94/d9ttV7
tfOkUWGhmDvGwsDK5VCD1RcE4hbxRhIROTL92ommFA0NGtdMEGIVANzjHD2Gua6+
Fkqljdu39AbM6TrdRHRBWTyi2mpP6NezelJ6yr+eNIAMYQCY59DCj7aKb2Ep5fJH
yr7VFDOku47OnB2zgndkV/1cvJWcV8BnAKE0bYr0yRM4VJxCRya+LHOV+7XQqZ5M
QcNOJXKTrr4ucSgvDrifVvDG664FIbGO1PrP/JfzOcKPydS5cZEtkeQL6196EcPh
8GJ9TYZngoHsmDiV0BXHymXNrtySde7bzsBuHZKjK95fuN51gzfP0+5ZXpWKyiuq
HUVBGAtA5r3OFKU60QBBsj3sBOk198NGA73m1TtjQJBQ0VIUKoApQycfOdMQKdrM
msBoOjapdqzdtuneIi1uFuESbh9QZ8G9GgXzjPK7To8XwJHD7wZkTSlnU/2/hrT0
S9dStgMds8hEiPLUds52a2Dx5hPcL3ReByFx9+DhRJyC5hNvYOP8hG4+jzfX743/
2uTZeneyl64PRgROGE5Bt03FxiHUmRBmFf9EBpEe7dl2aWPo9lQzeIHuFKkebuVV
lfUbFDHZP8/wbMjBAuFClc3JlK/gSMZErVhT3FeEZPKrxsbHKRxtU7ayY3nBwmCl
Neg2orbQh/u/cbCRQxjbpG16eE8Rb5ROiraz3F4WNYI8oUrYYdRMD18gufECjeSd
5YB9rMuQejnJ1N0kAKHJtFbIvqR0dt6R8H4bQLXyqNl77TjPzbnYGY+taeYYVr1r
OLsb6mDAnAd0CeDpXqbQ4xCuJ0JaCWQtOV9a1QSg+cu/AVUT7KIA1d1cHyhK8MBq
DXE5kP3E6VcaQj4ZAXabrpgHe+WeltukfMqD0oPUemH4t102WPHJ8LTOBzbS7u1c
DFLD1nHr2hqfFdQajWXZvj11Z8VDOj8eIJoGwpUDUl7CoYVoxGVlluzDTXukBo8p
OCqVKyKG00LlatmXmHylvAjQqg4XJcEH10H0orieGuQEE8379m3dtWDU2SZk+0I4
M5PeGBbwDX+QQx0rLC9NTFopXOsRZQ1LpuCLtt5KN8zASl4h1n8gOrxI8LJk0x0t
5S5GwLq5hDhlH+TzbibJdOpN+9PGSJW4sQb4s2fm2QmzbKc+tVLqdl8RqqRckDkz
6B0pw4tSzJg9vit/62Fzrvs5N0EJ861nsOjs+7okByDJATw5qkY7oQYXFymZCGWi
YtbGLY54IwlA7SMbj2KfkfDqUk0y/Z94jWjbTDTsQcOO+Pis9h4wFyykHlBwAtlW
UeH6u7KnLAhWuPGf5eICtpAaEZVTsHr3me6W1cXP6NeHYvCtGHs3g7iIx06c67EM
l0TzI4LaGrvyAaFNdTsoJULTjE8tPG2U+f0g/mSG8U/TvfeQ3IzLDiwB/IlaTWwu
HkivYcwppk5sG0g+zwH/rAbxMhhBEOs4XtAQlqo0/2IYTzcEzAvhkSGn2TuvsoNw
1NJrXusU4CqzxVBANtXbSgm6Oupd4rtwi+swg1GC5pVzAB5zhswyzi4C7SIix5/A
FF6BupU0W5SFFc0GqfqJysn9ya9fAM0ZmzoNeCZeUNY8iYSG6DBcfGnSqyT4RVLr
AZjyOE/9UQN/nVc3xQgH8Gn4jQ7ri+yT8/aBRypPUvbo7KbWo3fbj2V7PZblSxsy
XbRoT1v+Y9ZgNEw207RiFjTvcYJgDcA7IBfzXH0D+Z2uDCJl0bAis1GdI/dvklou
l2v1SNN29i26Ybl289TCnkducun/UnEwJHYzFmN93nvijCpduLfhQJZZD/wQVtIJ
nKnhM/RTNW+edsVvWc8WqXukVoKY8ExdlwnXZaxQWqzA8dqoN09OwaZ7Ff02c1dJ
HSFu9URGOD+lZyYnzgntzmNJkhSfETvRpCDh+XW4wOE3dCrkJGCYGxJx4kTecT9l
BFtW2ys4ZU1G6+IKF4WYZzhh1vEdNm7ru/JPqiyDQen7Auo1E2DYt+VRKuZFtooR
krwqwXFI4SlHHHPYQn5m68n2HGQMPfQvwY324V95CATR4o941zuUfFjDfjiILg3x
TypALziN+jIApUJbyK/gVV86wLS39Ba5TuATPk8On+1r6249TzoAqrweuqwkNTBe
qGCoolthHjhnb0qse+QuCTOGSFZsFrVBjgHuRwLzMO1KYum4UnzjOsY+gK69YkC6
x4Od9VxVihKO6jTN/pH2A+WTbgFNBPCi86mxQY0LXFDOtpDIVfrupq4f17rZOnD/
+SBY7EqftGIecDoE+XQWRNaSquQ4rUhhiHBDVhDytnUtH2LvKv6QknuFql3tEdAm
0IK6hNEW0U1lxOJs+lHvofj9wtj1i9bK6ktyzInKjMCW1zNdoR8zmCaM91bmqmsv
HSxyzMpzO4ItbsKCSLPDar2ajWu26OoTQowJLLP1xoPJ1cteqnVlOtOTxOs+1ws4
MYyTb4I8lPTotAVw2hYiZlrp9ethiQuV8Pn6A7wuo6Vt4X0jvtril4RfZFI2fPq7
loteYIjntz5wGjumZxs2YNZ+HS+8lijvFWYl4h7s4iyX89rzS/lLi3v3v07wiXXf
SmAhJ8/NmQo/05+cHJ/D8QIPK1gF9V8KY9UIXJJFZzs0v2Z5puONo9mY9T01EYiL
Q4Q1hOqEfiL+wXz0ZSAXYbcYsUSPn2PYSLwlJ85/zkROfJ84NgsrFeSIaqJOzaLn
owbvfE2E5t68BItTc6lF7yqZ+gBLTTP+c9saLI4npVve81c1e9ZeU9zCLd5SdjlW
3XmCfWk4gQb+vl85IraJviTzzdHcnwRHnC3fDmugN8CtGKywruxOFoBMRmgglqQu
7Qy5qQrQr6FudCAGec6BOCzRXJtoHi8+nhmHVVmx7ZROmOT83tKcNc9E5PtAahYZ
h1L5/nzrr58mmLH9G0Ktte+Gv3pC7YaZ+aI+fmwwveJFwDd/Vk9zjeS+LUavomyt
MGaD0Mu+rEg2pimk7ryddvVRVSMgYGFLikTgQnkDvlaKZIwMuajj2qou6pLQ54ND
TeWsHieLDt65Dcr4OVvJdNtTwNgT0umjOA4xrxAQMtWQztH7+h8VlnPbr0BWgEBs
BR4UJFlVBE1MahOYsx4R8JzsozEeElZGUdlAx/AF9P7Esi6DYmnO1CxgPUAcyTP3
jwMssHI52tEdJafoDvT81WtDqU0hFdl+PNi7zMmYqeWXAoRYHKD10Jqdt32IBJg7
mZ0a8A4gpcX5SK+69GRp8Ol4qT8GdfX++178W8O5GOFxlSnceXfLAQJQwuZGimHV
18z8U06OvX9Q4C6kAl4AvtqoGK8xhrB0OOmSKoSlNYh0Lv0EvKsmw+fSCyU/PgYU
NT7UvWUyzCzuH8LPRjXhJgEtgtdOykJD+8JE8hDT/Rq0lg3xzDoWb3bOXWpuhpwp
+r1X89oukAwdLA1/u3J1wC7+vkzcLwgtWS4FWUX7jYzLglofsggAzGX7K/fJ6Mgd
ukEH3+8hZNLKEqexaes8JqCZn3TNTY88YyMJKsHZ7MybFzdmVih0TZwCHxGI974o
gj2ZxHluJbnGlev88ikV8mUw12HrRvWPr9w6Vz+3iVX07Lu8dVA8MejUkIweid+e
Jo0tFu5mq+hYXMRAjY0Vhus7s6OW6v34ONYX8G7x3UgeJN39kGeRWtbLZ9aAdJCR
M32ComcDAzvC4dOv+FW+vSOsCOjj8cmpkriqrRFKRrGQ1Cj9ZfZwF7bK2lTpJTgK
bWFXqofTEoZr4dI9QK/LfIFAGcAk2JkzQcye1E7xPiIf90w757az0BtYe+wanY7l
1o78jPLpZs7g7wL6x4GqtmzXm054yUVhETkQKxFiAHnZ7eKWtsaJjsBeS/bKBQeo
cfNc7NZ0emEJMICdjT47AWy3V+kXy3PZllyu6wnZkTdoWpuCkhnHeaMJY4apZpKB
z6try2Dj5P0pFwOquBXav7vLTFCM+mRUu9i1qs/zR3daQcGUZkyhswQibBm30aZW
Ryg9ux/poZcqQh3MJ2f8kSJtWXl1z0PQWwMDtwf4WGCS12yC4rb6DemIZj18nLV6
vWiDi2ePkjffqKoXdpsQdCj0BQLXn0QHZ3rDsEDJKNZ4qGk9+xpS9gyKZV7JtMN6
ylRF+EwV6G+9/loExXUDpdcovbRBEbw+f7zyqBb3yK7UWXEAYNb6Z73dYUE6eCW3
oClu1A9W4e2WeD2xolkqNtVFfFqKDBG6X/7ImpHCdPL1IaLa2NZk98leV7hCYbIZ
k4Z3YUG1h7ggwyEmKQ/znpnuswfIYfCcqk9umTqTtQ9C67cLGHgWbhgz1NjNvTT1
xbJSDYu2+pfGvUPdS11dQpdWlNo9qE2BegjwYOtoxW8eJSYVdWZfETDwQvJiHHjS
58oIU5+Lhbig/0Pr21ljqqymnIx3zQYNeBvZQc5UT4aeymyUzjfhFID4UzBnYHLl
anOl2bcHzJIouChXIgEhBNlqkpmSMJBdG/1//b4xJXDcF82Zu7Jh7C86DoM29zxR
Sp4zXhixkj9V4cE9pH3n9A1euYT3Azd0Qz7dDj2yqRg1dbbVvDJSMCi6rUKU1VMZ
FIqYvvsrFYiGDBlg9i8W6kkQoxRN8ZaVL3fMubFsVH+ToxYH+8u4z4resETCqEoJ
tbJQrbltYA/Ti3/P1L4yqJlnqU7goUFraWeyvn0Wse1LjpWuKcom2rTr/fwmns1O
wv05hMRoTtkeBGyntTSW/8t+INKoSR8D4qtX5ksI3yVVYyrgAO0EWa9ApMdE0bYh
90/jU5avh9sD9fAOHseCY/PnI4qhr0O75ciuYTgRRWBGwKfOjUYVr80j3NQpkfyi
Je184mxyWf9Gom3dewrzkkZ2dbHe/rzbka95YOl9w67gjmx7vwg7gld/omYdzADH
1UIakrh3933uiKKwzZMe9Dozp01pWT28wLFixjkSCd9nXlZqhlfKSuHVXyg2Obpb
SCJm8EZ3anCogiiaBTe56dqmk3Cnno2H29h+/xihNOnIfLE66Q6K7iltzhgMnsHZ
oJRd+Po/B7AJVZwL6nZQC/uvg+jJ76Y1EgBEgUcyTcP28sqztULYOjOqSNsT0hvL
nrxF9NQlN4g4X5ISQcWC89/N9ze46HrSZcwJA7DX6SA1VwJMcgsoteiSL6oF86Wj
P2FHc/2fnqGAjpvTSDp9E6b3X69mvSm+RXylidWcMWhNuKw6NvovO408hllnm+cj
00Fib2mEByRX06oVvnRCyuR5RBZow6wZzPiuNApqtgknk21lUeFb9acxkI7L0umu
6Y4iSmrAoiih6UCsrfMpVZdCHWr+0ZVRUHufpcdwHVVdY+B+NU621x0RMj+eDxB3
LXlfkri5469wpTkYfTdwOYxtmGt8lksO+9EHj883mHSuLMSAAAD7iWsG+eHOpB6x
MtKR5KG0RZPJHl3R1xv3FFAc+GyhkMY8INdGBAXAe64r9Pdn4GxWykiAA2EPhW6E
jjVVzBajjdss7hfnbeHvR+gEXVe9V57tZLnbZ+wPzeqmF0D0DFFxBiNu0eiYP1uG
8WGyOakkyPQevfb87Y0OuUwQl89X57dOXcnktpicG2Vs4GITiikALSyQTQYNgngV
CgQGOtD6hsMyArgwrBwKs91sCLil7AKqrWc93CT7TdKZ0Ii2cQJcg61073VGdusF
tc6jt7uMWeFirhfnwjuBZ7Hl+k8dDy1f+6wVLl7HcxK7DL+lRd936A4UUdH/SvjF
AvDfQnPVeu73I0r2Z14P0KXg6rsdqbVh738OQlJ7eR/nqiwfukYO7kE8aYznEUC0
Dp1DVsYgjdMe4bA3aonG2VmXMfMDkbrveGa3WUqGGoAWLvHiP9k4U/ACIYNHLCrf
opAsKGYiD5Roa/5Q0fx0aOiuRS2oGWhACC8/w6iIa/AepWlU1UBPNaXtvYKUyPaj
PEXDkV9PW75jzwWlfCTAmE4KA27sOJ5japThBd36jCJuSvpLXAHgszkl0s14O04k
J5x3tm3zmdzPMxop6iL5qof5FkUBhZc5G32oYvpaPvO1pWUhl3XNhZ2fJn5jnQHZ
Bf0dKs5L25LcNLKhHK/MMExI7FMA4XXTaLfu0QUUv0qOiOmeUfrHBAuadSOxSjek
HmaZHvx06GncdoQyKK4bvTqIlnVykQtpJwPW3xntiygb2hwQvh7mi5sqFgQWTvGa
3w/QsmwwY56tB/Ax8bPpb2a2Ww83yh/UQ6La6a3ir0oKLWbhiw1mis/HG25EQRbp
qyG+AIDWUutJBtw8G1TWsOpmr3gVyWiUOSxY2cYa/Z1++zikbohWr8TLEP8PvSRS
rL3wdREOXY+RwzJYtyfN9ysI9r29kAv+DlF8JVX6IsiXQPlaEHwA3vpYdCPcjg8j
NHmsnZvoU/th88f1Xd+x6RFpTaKi2JTaYRqw0Q7MO7uABlGDc6lmRgeo80RcPuQP
X84E/P55u7yJRu1Ce5EzwtY+z83d4b3KbnCYKZhEMkLW9b/oqKkAtaEKYdstg8io
uSMlCHifFb135ZF994OMeu/2WxE8xR61mfljrFnrDRKCSZvsxa+JL8YpTpgOseFp
cjj3YdUo18bDPTPpqEYf4q+uYbTXmziWkWksWtuit2bmYyxXGd+UY13Hl2qpQqlF
F0urGoHtPQdo2AvUj9YSZjh0bMdLKs7C752Tjez7yJhzhF5ToKeLqmbAvnXgf0qc
KJm2FYxmlhPX/v2Ug4Bu57UXZ2/Jpu87BNC7X84fU5Tf+ohQeb4FJ8u6pxGmnM65
+PycJKWyF7x8M3SCU5GyDeUSyesV1uCKflCK0qeMnGOlmw3TWQzZHbBDkuNrk33R
UT5OZNuOqmATmm743KfRsh7K9QLeh+oeNegp6b//WIBJq/zRj7T8ugViamNMWf1s
FtRWRAOH2i3gHuU0/R2EMzN8e0s/1dKrRA8cb5NI1NQUyKWzcs0D5mm6FsE3NoYr
Ki/ixFjwQhiEq/IjCj54wRusZX3yWJAN4di3soExnHSyp0VGhN3+/7mr+4piZf8J
JGXr/nxy2tV9tkN1tx3KZ5OMrFsir1LgvSHQDO+vtxQLarO9qDEaQZF8S73Pshuf
89JrxHMowLJ2t9ehz/lf1AFYwZBMmCLVmLIYE1nQ5BbbgBFGJ/HhNXsZ8VKnwPsW
M8vbmFTIRQW7x1weddsglr8olbPLW7sOyHkPKLKsYtXXlYsnK4IZLAMvpy1lcuKJ
zl81jK3JNIEOB/zt65MXw7KSXMyU9+sIS8/MLE7f0Xasxuuy9iLYTPqc2TSWB1GO
zbTOiukjGvQ1I/0be49Ib13De25xAtC/etO5nhlpw9GPRI9t9X3ygqum6urHc56Q
yUMuwXuHeASTf0RHOB26dmSG0pyCsAQQ2741nJuSlW0q2TXpk0fMyXxaMKr5OuK9
AVY5NFGTjnbHFUzz++QslIK2OHms0qqBwb6baT7vI0d2Gzl9vYrJOr5UUS5m4FmP
kJe3iObyrgd0qfn36L0pLarJUrvTxLjUE+7KdQvvJrb9ycQlH7ycGFRmL3/Fhen5
cnChJ7rDGRTVe0ww8ogg86zT+aUHkbFYP2Brl584PPBVmso48tKGwSXCqZPO3NXT
Rxr6fRp7oBdSJ1u3+QOWogwo/SKagq5Qqyv4E+xpcQC5bGSBD7OzT03OPDl153Hi
OSLN/qt0KL/QTpuvLzsVgeNz8pzxcRSbhT4iwT43SXYLkIpLs3UPFeNqzGZu7fZ9
j47pKFUdT99WNKqQS8Bdzz2OY8YrPMtZDPMHSZ73Zz9hHZj93SGF/P/G5q74InuL
GQK7GgZDKD3exVJtknHep/tJijNaNfCDBLO3MpThtOZHIV7z/KRtFJuiXT2qcB39
6aXY/lY7g1WFdDoheFRXzRpGW+1Tq3EQBioq0sg9ZoT39eyvNlFcJ7TfVg0TH139
cfXmOcNcLb/JKZQI/kXEcugn1eURDJaxSZ6AualOtXZv6D7GTl9raA32pU//pQbZ
WoIyLQg3HDmT6fLEXep1Sron3I3TJLQj4mPGv1tgD/uswmOJwdbHSBgVI8MeF58Y
p/XjITAzkUgsXlV2KO/wx2AVQEPZa3aKpA98nSZpK9IgxCN2H2sJpkvIr2hXPQPB
IyWYZDu6a5BBN3AXnPqmyvbRJ9T2tlRS/RRik5EMsT1PBr7RUt7bs+QQXW21ycvw
ltO2R/YbRbMkR7+vMNzyu5IZ+Vvwdc4KzcYWGU3kLpmL9SrzIhva18tiCkzOc4Qj
WbsXvL3wQhxSxQ9kgVTLxJJdj2urYae9w5HNFzq0Qc1NN0m9tM0emQAOaoysp4Sg
hp9RWfOqdE58DSvqb/1exNx7HQFVsGFd7NpoH5eDxIJo++TNLvHWC20OsaUwrlmZ
REOfni12pGNEX/VBRXcZ2gFceWCc7hU9ovTR24AIQDwj149kBEXBLgvcKacRjOYh
d+GfNZC1KOVYtZfzGd6zXG5vopk2GPH9d7SoQC4uUci/Ys3io34HcezPrJxbY4gI
fKoDtpkKX0+Qtqc8HL/SHniCavZiFlfXkoybk2hJSMwueMRbfCWcyhVTP0YTe6LD
Jp4nwQT9/0RL4sR5Ej72mruqTzC0ltb7aaNM4UrEX/ukFfKqXQpkywN+3se6NcUc
DBwdNdvSmw64+Jn3xA60qn4Q2pPMNvwBDrADGQFdWx+g6/Yr9u1L2qitTKez/XD3
/zMYdy7zpDuWVPJS/9HSivcgTUpSQz9+mcpTnIhNSmAih1cM7GTmzFSwiVhoV/6R
y7HPLpmKwvIeCu+xlf4HYUt6JIr1JlgzhBrkiKT1JxNvojHnLsEbzJFxguEK2jKD
mkw7aBzP5MaCuwzYQ4MeBKIaCLxWJLO3Uu2qprvbAbRMFaGEOv8V7uO23h+kMyD2
rPjCHotGUZEt6gX1lSBE4Wxj7kzRmMSGwKTDPyOBHwGJhMXjuU6czp9NSEh58Sgk
AqeeM7HqdVp4OjS/bUeKsz6OAltXAvjuKPaHPhwZhfMZ+22s9hfl4euOWXs6pcDT
4w1lyrkAx8drEZKcG27m53oXEl00Rmqr6+LnQPsA9xLxBzN+wrlg0ZjJs7KHSkl7
GwrR0qCmHYWvzXsN+LmnoZ/MLLQe1P8Fa4RZi5cr08WtlZJLiJOy8rqGUVp57inc
n1P3syC4ZnDd5k3/xwCRPlgBonilWMHY0XwpcwbJy01bBLxpNlwGEb6SaTCDthzW
QbzTxM3ujYppLBResQjxXD0FfI1pPZKJnZQSVk2HWnn8vHoRfcOFJJpHvzjmM2cQ
fW7Zz2ZuN+vIevbJs3L8l9mAlpR0gn7kmk54QLYo02V1+2wu2ZN91bGEq9vYIYbS
RaaGCtSKNHz0pLnu2AdT4OqHwY9SyvYHiNNbWkNSsSszqolo/5iGnEgOx+zQ65yz
jkcL9Uv4r5zwuojAbwxuu1NYJ4hMgKHVjJSVvqR+BouieGLKDmbpQ1Pn0TyFfSwn
GdimIJsoZ+pxAEMJT5kgH9HGjYnmtFpFaqQ5r8lV6Ddtmi3/YpzThKKbfcCC/+B5
N1Xi8Oa9k/JNg5RYKFOmHV3PhxHKrztUEOns7K3ugs9GLAuiDbURCZJXS4a3XMPh
2xj7iLozLb9oyHbVnMZDO0WgRnT+yZmAHJAe/5p/dB4VlQzpb7rbpGDvS3dnYtZv
a+d7Xw1OC2aVYlcJ8hpsCA6ki2Bw9QxWvAIDI49J4a32oT1LyPtwqHJmlfZd9y7p
3U/1Hcn1RT8O3106ZlFXMnhGwCCwjrBbNMIjoU2Luae//Wd39zTP1b0FFVb1TFdX
hLQ2I/Fh4ct76TNd0dUWzla+p288iKK5KO86NJVgZCcjxRXdhrR/uLFv/tb3Hu9X
WrMcUcLxeNXpsMAln3EJ/mtY0A8/uNBPzANgkG6yKxBiT/R4XyOJQmMtFS2k5fnb
xbLFYL9iN22a4yWlXk23c2T2l57ADmuN+dTVVCkEzdWLihkYqHbO6oPn2k/14V2l
5sEkG3aLMD9DnmzShskrpn/I218zCia+MXhhrJTa2ZxPkoLMFAIv0eEcF8EDwMjg
DNatsWL57ollfZ5c93K5YhwaA1Radh76Ui46STuO484xpO7LGjCesKkj5rFA4KzE
7koaImDPGExWNufT2hhQEPunC44WqL7qXOU0DBYZYeG6/l7Fz3UdVqJUbdvkKqA3
jtJ1VCm+aHYtG0iUmnZ8gedJAHHUsLOmgrW0KPnaCrjswFSanvR7uE0hd3X1rkUp
Dg40T1JP8L7A3SqLbYoiz6c1QoR4QRx/yasQX2VgR1Nz7Klxr4zZDEX4bx2NVKeg
mtOQToBZ/vxBdOV/+XqKce2hrjlL3RUDXsBZQgq1lGTNjHcN+rRsHeI6snJGeHil
2MOBGGgBw0N7/6M+JUKOGg2DZYn0DwLfKJZmpeLMIkZDreP+KxOwZ3SD6R/r2jsh
tE1jCb8EPjgutkJjd9zJdaRSN7TLIACN28sazSD5KWX8Xe38AF/fPK4LLcYT6AmQ
JKesy026YoATri3tOrZECaTX1hzMtSUsoyB8UoP7dKSTfP0xy26n5QbBDDfJD6yJ
57mvAGK61BhRR1OXu2xYMOCTQZMVw/dhfZdVzutctDbxSMvGYJOcf4u3IAU5LNfo
t7aGgm00zMXvaRsE7G0BxnkEQal1c3MPPH09So8eQcKIKnNdL9/kJo5+HaeOAPNU
y/zGXg63eB1ikGcWQ2x/gPOXa9TsxyuBUx89SdkHbn3gCx4fGH8dDtGXLRuXqtI5
FhJrpZ7N1rlTa05GQx79TtgyKDKlfzG1RmMZJlO9cZJdNFj00fPQc9t/6ZUBGcEW
jv3jSOrENsSxDRQWLtGv+Z+T/yOIha6+JozKEE35zSzqz3WBsebuvIWsmRUMco1l
FJMZGZLV2OVr0ctebTHEVToyjkNEncOIGfw2pFC1fWl7c+eQc56+7IKQQ8LSIGt3
bw9Gt89kcV2oo+Olj14e0rqNnXKrdX61zvTzLjCMT44wRdeoGs0ppCnk9F3dT1p9
eWZi/cWHJ/GHItFTsjQlK5eVO6TIjOShnDk8aQQXoDI9wCT6R0qKVaWepIBVN0Qn
UKGjBepLMHHgR/htvIokayTTkeEbhwzexCignWuzNYFOyH8APYdBImQh9PbagCiv
NGC6fBykagTF26/5yiyJWHeqXq2ZC8fpZsA5rifXFPcP6NFhwt5uA+ZzZeOyxnfe
XrDvwJeeJfKsSClTzrkIzZmcwQBeCDp0FmfG/ISdhF1vFHWCUvAMf2Rf7twkxqAf
H9uTEX+izwlEL/bna5IYCz3emgUfOqH+fVU3GWJ4PAJnFSLntMtuhzdHdircDmJw
IxdY2mxbTZDC3ba6L0lTrFWFLbWmhbHx1LNOrs6Sri30kGNgi9iJ3OrfasV5JR/C
GTuC5L3zew4APj09t+wyq7Z2RRlBS9rAMu8JsOi9H34LHTD59yjYv/0T9WCijWbm
167KGwZ0OF9E+uNM00WF4LbfkE8JTeEKB28rn7Ts4wq4o+nPI3d1uYVjxhzqczGh
BrI5xiIKcnk3yZhut6KgQ8i0PAnewX8bj5ahLzvuyRNqvPYJD3yqd8s4PM4zNvZY
oGT0+eSqd8BSdbTKMgkiZFcLSIRAH05Pr42K+KsE+3Ufs0ADIjcSWZNLQ30paMLs
MjMcK0mlKM7qUZa+MgUHNhGWISj4ufe1k+J+ho+ZINRcKv1NvkCIAecNTkU8PCHX
4UNS8dHMYcwzr6EjQeGRrWbNGy882eXQIIlBXFUeR+vPTX/arq8CB6mxKSm0BEqQ
XbgmMq1bJQ+y0zHpfsqMbo3qwkAzClRJrAz8gLWP8VEtTGuhKpKVfFD4b0sOIAU/
AuPJDMrFmkXdyW1vdvuEYH7UCRHSW9jFCmR6XNcOlXEtCMHWWFUSrd+ETMYQaYhK
Bl/lWw36H2EEHv22iYooc3O6l0SNnhh3ML4TUel7snU4IO2JdmbJqNKiJGEb1d0K
L3CcqCMVb6COHTx2S7nJLPv/unxEM3zpFdBHxFKZzMKOt3Q8cVMLmJfk9Wv4Begr
6xPwY0j7BAvc3Ho1NK0yCA7xFzK8u6Q53jwJCXsqdgmlWTY0BjZPDViRps0w8GuQ
8F/bhWBNdG3uw/cZXgn4U5ms1oEND8/SVeyIGCBkraUJS+kUgl1r3ii6QBAAbFb9
MWo39VC/e7XvvnfCYiDgk4UXxSqfOy9FYHJ1i2JOlIP/n2rJAE8ykHpJThy9UYLk
JM1pvSm51zbTDFSsZPrEeX44LWvqaZZUaHkRpOrrJ8r5tUa/lA9CojGncVgXt7hO
LXlJt7Ho4+D4S6IYuemFPU3aK0JLFCnxOxgq9jdN9X8pitz6N3ZP/ckkjE2ALUDr
8DUAVaWT/RhK3fcVskt9eHoqwvw3gIO8apiEYFc+NxuUuzeGcOf5W1If/L4Hp3Ev
qTc9gtUPQPUNkgdqKTVx70vS20pGLVUNRt96atuowOjwMn7ZlE5S027s4y4p9m4b
0RQxTxb4p7lbxt103O3JfE24rAe/8dqGDLUFn+IELqljYvgGnQc3UsRlVLo9XkeB
+k2dUubQDKzzdd9H+RvVHMgh/rHeFm6TSd1yrgfWetfLa2dkS6qtzkAtSJ9FS+vY
o181BGHreQ2IhmWlpiZlYyzPgxFfHzDfwuT80eorNagqBFg+Dhy3VYrAcgOfSpnS
9w8DQRKO7G7WQQZgsMwGwTOycWtcv6qG4BlD5CgLWGo5LwNhQWs5kadKvFOponBf
E8/pj5p0jwTnCU3nTd55yqgNWtD5UsYgLM25Vq6X4/XZ1go/oeIGYON3W7QIycPb
oQM9PJG0jskKbsu+L05F67KjBQPlXiijAf3kBicGcNM5kTMFjAGZB5uTZ+sbdL2Y
lgdDnx8bbzF5qcIUxbRRIGjSL8NOPmQaYedX034nHqIv3CSaGwIxLkZXRwRQaIuR
F+FNP6qSh8lxobFR2Z7jOXLLmSw7cFqGljWB+eHJXI62AYKE+za0cIxnBGuYR5vX
Yy6IRJv+IMQ5ysB/H6MPoRrTQskdc7piZ1cTGlOLQIJMLPDOL69j0tSKTKndpCQa
N4A/spr4SjA4RK3uQ+fgIe7rlpWo27QrWTLLr6HaSmJ9fYA2YKRkzXtGO08nnsr1
0rv+er0r/j8lyGikl8zXEY6NlUZZBOQug2MTU+YoameJ52fwJMwJgYlTBtxydC+d
shzpdwDSliNVLqi3tlGx0PJJ+SSbz+JZa96zVIKHQRzDO/VGXBxD6Byb1wyC/G2p
lZvd9J/Gt8iPxMMYDVq3stjCtIGjjTPaxiY4WAY0FpETWHS2I+IOoTMaDgdULpqh
aehXjpaPVyGUXKKK9+mDzMW2Ek7QI+9+RLbaJLAxS62OZoLpSBBbz07aw+OwHstb
pK/2AxEI7P2rXVc4AskllR5ISFRVo4WtVkEq0V5hHJ5H4CLnBSSbzuWdJFZYnLN0
1V6oAGiWU0VhCvlG5vfm1gtpfLyzx+rBdFcpCMrIm2ZLdZmk/AD7YhKfY7qYg93a
B/CEf6wGt5JDZgoS4FWY3sgxgoC63mnZtQBBtZjOUos2ZGaveg/0prle9bePL0Bg
pQSkeTSOvGuY0dqts/lZGibihj7AhFJDi6Juxwa6G5i2BZvkEn+R1TtaqbaecOuu
Jp8qim6lXi3RXEVP1j7hrIEyA3lN8Zfm9MoNTKVIwGJ28A9mOoLwC+GfSW+09i5/
HBbRHNDhijxu92K/2lcYfmx5tYblDZ58343lnwkw+Ob2zZoVuih/Mx6ZAiwO4mrr
KdPmYj9jj/YEI/K98URissh2x63W4eCHOHYKWkxfHGTmntEbPs7BhZHyONtlm4Ph
gyGzy44hOhajQ44kl2hm6GTp+hSJJj6pZxdvxiqsD3eDQBW9F1HqPh0nvmNhhgIk
oDZc+d8ctYHGuYmIcoixz1TgY4dxPQjVX+SjggnFiXNspL3qAVEIP24+vmwajj6y
8hz1hdWz1oCyyC3A9sI8qJB4zkJt67zINjxrfWPTh7MWK55eBR6cSdaFDQ18S5Rq
2iyuvL2EvwF4sJasjDiPuy1gMDlcJTe825cnDGX8XsXS9njYnA7EB4M0KR3AzbpA
o0B/5u1PgEGwoasmUc1BoFwpVPTyIqLcB7GwQei900k4wGjKIbTlQIFiMTciAwqv
QSYv7Irn9P8iliHiV2+TAf12OAk6oOK43srk30OM1r4XYLLdwd674Epa+kQcNlBz
EGMc5nNZ4Adtvs1L6BwRi0GRD5O5abnfSKRokw3lSWvE0Jmakx2hDnV0yw5BSXdY
2+FnjQrDZkyQpCQKtM0VIMSBmO7o1onGIJo0KMrOGSCSy7fXUP7kiO8ThHSrHTX0
Aqj3+cnEbWH/kqa9mk/T3ZKDLZfpLjhGxAdaLdiDCER5KEq0rvTEAY+dgW8dxL8p
kfFEZec6hpvPsuHTZfwQyrTEsqUvgpwBfd32VTpMKwyBjZ8uf53n+pUDLm4DPtVW
kD97Awjx9hlAPVFnbi2K4hni0+NrK9ZwTSfXCuNjmJmI/zO71E9D63vYyKW5nadJ
kvFzyjdY6NADU3Dhw3iDHMgxmDREUt3m0B5tbIs4DRpEtyenOvFTAxtsVeeWHG7V
uE557RMriyJVOIV2liPpUd+bvE6HOf/N5WZ7o5i6h3DsGFGSpQHmrGbvPoGtiU0/
B9iNNbgmeg0X+OkruYE1SQpSkWqB/UCoU8wGS+Bco73yHjO+SsS0Z/lC4gAZGm6V
8OQQNFTmLRV1pKIZponCE1Q55Fp/Cx3ORN1Dl3Ey5EPAY7KN1DAVfirCmEyMz53u
zNjKK1MnUPXt9Dz9pSAynZHGuWgNFO+sC7RHf4pvTVCHz/+STWmbdQ64PLcYP+a6
uoWwUeL0ubA72fGn01T3eO7JTZoQoJKaGNdMoYERN/815kdCXiXsfeuK3Pdq/5Fk
o/mPy7zefc2ab6/7RCf3vs81dzODWmpYnYTX6xVdi7X3XFlzp/4hIq0G0FBYnubO
0q+Qo6uUoLSrIjj36ZC3HZzbjgCfPFR6y38DTEQoeeHdctnNtpY+uxMd+BgCeQ4N
U7yCgJGMBy/4CTIBbZD261UpKa3X78dREd/Qe7vL34n2B2YyNT+uRjdgV1n2dku9
1mIHqtMzqM/Q4r34mzvO4tw5u1QJLs3Ipy46aI4OQkd9TreKTSYVeAvdq/iv/BPh
C6giFz6pHPMxWMYi7elZCBv07K8zqLHWBYb3op5js6L3kEg4Su5h0kemFZ1BKdnU
VM4iUs2WQxe9oima8cAdsjSCks9b1r6OfwC/vrbiHTy6scyT9OselcaZd+u26ARo
ZUNqdL+bYBb6Fs9MUzavPv+5wBWKQb0w2JnXO+y9YCyCMZbrbK1axS5FU1UqHkjp
a2tL7d127QF1wk99EdFES26dtvQOZwZV4aHlqpb5SRlXgmS0iF8THXSsV9IlLnQt
VCREvts0R+wg7Th2L2WIshwUyz/2F/WC8pOV2o5NvZeHsK/s3t66k5BPBqFO4eMz
pQiTJnpj6A6vQZ3qasraNXVKxccTk4cqnd3IRolhR6WRQ06DQOJyPSOCrC4OcAO9
Q+oRCjNS3remqxZEdRg4+XHreIw1KsOhwKJz5qaCKGo4ghHN0Kr5n918ut+PHmZR
M666GoJJqVzBUVG+uRukiWoZ+KFWUzDfYYWrMxTF44s5mQu0ul7pavfCW541THf9
Dqq2pmzb2RaLCHNMa8rKpgqdpcwWIN5Mz1Ve/5xUqg7wOzncUZFJZLCKeutDKH9i
CrmlOfYiwyKL1MC9Zb9Rnk3/+w7YbkBlHUjrvxs6h1Gm14UWLko/I6QSHIO+L4ya
9ygeONL5MVVBTkw58AnDVrPHk6wZgZym7fVr45rUHoDtYYY/60hbJEIbD0dYewhm
ovFm8aVSp33qEopd983TDCk+XLZ8ei0dZfoznHh0l57ly7KWWXYdYG1B04v6Fe0S
cYGig7l6DvHN7T1v5XXQ45TuYUndAtIlLh/ZolExkmbym4PazjjSxw9j8EFRwkph
lr/mizPl4eXxRTzq5XXs755UGfOfh5hI4+98Tcg9ioiYUL5kI8dDcwDARVK9uKF5
+vLJjaxmT/AMRwzxS5mWnC3p31NKp6rcv7rOVb57bpYcinGzDPm4G9FG27llGiqH
p4vZtgvUOGX5WYgsUs7CShOhfkSKyQ9NjmL5JMcX7zDGM4V4VMFXjoRrfUpZHmNf
KqEo6SudOe2MXGvX+cvshGsQ5JgvzdIa+AreJCbQRWhRbdjSkSMOTDl9XJs16tiW
GiTbY0l5wsx1VLfB/OeiQNKrboKwdMthZ/kF6llDkIUQBZus4+x3o/bblGTSVbTG
escCdBBq/06jjXreZ12K0qUIZPe+VvgIP16Bit4q8r/TIahJUQ0sud3yiCmSd9z5
93BdHGSR/I43LuybdBR+XuVOF+FXb0mik5jK9l/YIEF2lutdb6DARovKvdefZVTq
6cm1vHhe5qK8bYa1hV058RpGc5ZG8ckXtT3qYAAHWR8/CI8mWAE0no0uZ632clBt
PhaQPXgXS2IpZVs/15dLJthq7iYdDRS2MJ05+GVSJjlM+w67rnMKBTwJ208FR67F
T8XLiByo9MAmuYJAQy9z63TVWzRv975qAqA5DJVxkaM+YORKNAz0KJO4HQNMFaWJ
NLKXsGZudT8zit7RjRoSjoyYOD+QIXMg9jpx6ZgrOtUyxnf4SReDd01H9iEG2CoQ
7Eyll8U1zhQpiN7Q7LzsolMDNafaZl8kUmIQp2rc9+z8N6/DrAiclqRszl51zam3
v9ZxYSQECcEqOW7/WfOQoUp4T+S0cOqsJaiEqTl0iE4+zKbDYrU+7BRIF9x12CkR
+EsqTOa4BwRaInwUxaxzPWvteevgGgUtZ2QF177L+6ep5MG81cY2ncGa5/st9lRL
1lUsejNG2nptxENzsIGcKzU+/wpbMpAQASBx3ofhQKTfdRYdLqwn1xx3gFcitxha
x1ai7TX83e3LWNopPBJyXveBo9UPFYF3ZlEMFX7WZWjRwhEdyBu0RZlgwjA4QOnu
TO7/iTUnPx5y0mBKxtsXEGZStbZu11Xsy5f0r20diXrpNG/d8JgwepBoPp6o0fDN
I5O96uT0SSb9Yf3rsXksA2Sf65qksos3G2LssIfCZwPceduXRwIrto0LCeZ9llUr
BG11RO4EvnLx+2ZK4SGHvjuPyzHUwF4vM7DaxMFvC+MMMoFqciHaNt//q8Gbs+Zp
nKhk8JSmnct7hHYTvkSQ0cf1wokSyVQteqtwVa1VvR9dk3x5byISmRXkP/AiQr+4
R4C6ZTTxSRq3m9VqEBC+EtxrjMb7FeAK6ceB9/+WRYPv04g/jGcjMMrN4cU6WZWe
H1SJKi9kvghH63SL39k1qw5bBFEHA4QSmWgtC6yIrwXzknVt/DJyEvPgEMo8U7Yh
tK6A/NtlqEXWbHeZ9cwHlX9kX85eGU0KLCVMnlcKLT5v2+2jkCUlKNK6bFYBWBUX
5h1OFRyTndqtXx/3VWXgVLGjPjpLNKtSV/Oei9Em5SkVWkf6H7iaFq92L6kTK0kI
f8EC6yiduFBwe0wALi0F4xshNCiUMBDRJPWXA2/hatwpvtTMAZWJ23WWSaNuPqCO
rc7F8LzdyENqFLLKrAobcXA+vLr0z+6wudVXy9ZJbKy9BXgw0IsZlEGBdcNUGF8k
3lhEyvuiR+jWClH4f+SKjJRwFv/0OluDBi9QrBxg828hDpTdlPG6pDAM1GAdDjcm
OtnevdL8PJSSUpWH8LCPzboJl4Qqj90zbzrNeoGNu6y/7bxdCc27h8vlVpvFVJko
GUFPvsVTeWTJqBEwLDYEdwkDrdDD0tz3SO05uLZaYBn8kBlfi09mkX4mesdjRxIV
lb/Z5i9NE/sa3Oc9NnoiP9ykpmOmowX/f4xjZxtnQ/YYrkemAHuKfoVibYoqQzq0
5lxNLRfHnKAduhNoxEKy0dgmIx8icr+BsHgRQXAGsmCj/35r/OBl8uemPIUoFXiH
9ayI0QsoEv6iYjA5bGxW8kNuydcqDq2fWSLJXTEF7UzNKvr4EuQTpvurCL9TRXd1
j1e42quPh7i2WPiqxCDLVGtcLQ9BlMlczL+x6U0BOUFSscBR8koeWx7UG4vSH+tW
gH5AhoSZ+Cn7gItT0Mw3+mBnLCEM1LcbpFHqtM1S962xZVDz5DgxLzoNrNPzDNGy
B/SyJmjM8UpPS+kzkZ7qzh12QwdMJr5mvM6kvFZRG27185W4vnAvq/Mlbv1DRDoq
MAP24bzy5a5DtQnmTIk7O7pcd0tZzZLO5b0NVzxXcjEQ4MP3/9CS5SgVoytqDrkh
SCEM7FZidTm8QukR18U3E69OunpHRJpjP8OLJk27hb3Gu1UYY/sCDLrocjdoLc/j
El/I3YMeYZt1wXbWRbi0+fFyDy7oYGCIuxRW040OCSXgHqmJFNPSiqdfIQsrgryr
iBSbBdK3fbzV8PyFU+bp5wBKbfnRulsfoeDM1cv6auJN6X9aw3G6t4PraHeQO6bM
sUtg3/Zdh2pl9R4dVXWBBeLLKYJG3UrPA5KYuo3UiWfS7pVunnkqR2pR2gwmfRAh
xrkKMbNz8qwnpyKSSTJVYC4FtA9MI6aXuNJKjnJJI/f/jd45RGm4iZgAxgE76MZP
yIveOCi+ZeBGs2AUqLwP9XNSq4WyCk4d6iorhImPmCGIqQg6zdvww4HDQvqkK1aD
DhkuCAaKAts1BhgQ/iU51oVawtDIU1YxmBBLblbJ3oMzNK/HzOy36NI2ygQpt9o0
/E+Q+pMe4EXHfnpBVH0ttnnSAIV1/F/RZ8Tou6Om59bGnMphhtIkSWrjWiH3iDG4
nniW8q2zH8uhjovZ9sZd2hD5JorqmpAQiZcgwtU43vkVzIN466DHCgW9Mc5+JPp0
uSnsVfkheDtEvljY6Pkf204YNWcjnsBPOCxOrK8rO3HfauXgAbScd0kOTHcoKPZL
ifEEyOlQugEY1PrmUFni/dUZY85bQfmA1rU1Zq99QSLbvMZaSU9niYeeIrz+Xfuy
JxQ4kkcIYDgkIa2L/e+RwSlHElR8kAP8kGh/fXH2GYZljVCj4rgfHBNU3RMGiizY
qwtrbrG/j0S+us8vyTbLW4oYRYQLNP4qqSVQU0E1vumKLdbMF0XRtVu0mSBdpSdS
ED8IAUa5uH55byzBsOwcfqkilvPrOUGCNEcaECZ5siPFMkcX3RiCGux2Sc3A63Yc
7Z7vq0heX9mZlgVWzQ2A0Iai/RXf0Qv0HP/S4DzAOB2YQGhx75xDpxCB0tlEOs2+
IEqoHD2S1KL0ZPjlAq057COe2u9rIHSDky6KrXINvfTOLOfBeDlhnitO7h67gMe1
tE61+IPTzc9fBj3mIG78Uj0ReUAC5Yv23R1er2F3phlIAvOuJFE5VGlmkyMRfWVJ
TQ0HJ6s6RoxFevDWPzfnWPH65N1ahK8VYhrfdzryvQdlkvWvI4pxMiNAzEBiheS5
y2DH11pY+SUzSn4Tg+3cIRSx7Q97ABpw9z6f3c/YLYPJMY2WNg94qb7K+QJOL/+Y
Ty1BC0ivTz+LwPlCModstQCDWp3D8Q6+Sp7BOakxvQh9pzQeFgmfrKUZBRvZfD0r
wvJh6dZvUGS8qNG5IucZCsj29cQ6m0Sv8Fo6GllgDBjFNg/LU/1QFwOJdxvVS4HV
NnBsnjG8Yj8oOEPMFkkvJGCmaczxKwU21JHnQ46G0D4GlxsBrbHmkw8+Za4WQzZ5
X/MbNwAU26vlzAWvp9RbNgEskjxSMw15swsL2FpKaU3IHo8t7AHQc5yvaVWMcgsq
seYOKX+DjBg1FVRQVISN87Fi2HII47Ql0GQUXWBboADfOZZrGw4/G7+BH0RolpQj
V+FTkxl2HJGozJvHQuW44UqP1YXUbaTINmRf4qLlzzFAcn2V+n614OHGBOUkpZ1z
5OpNsbmlotlHf2u3ieW/tI8MSo21Vaj6/4xtN8e4J9Q+PvZkZFeyAXDbvoVRX9i8
osZAuIAUWCPtQ77IAuGHpPuRT83nWvbuQBVsYvM2fXdU4CVJjtv7xCS9tbtiYvcm
h9Xu7qDAFc9asufk4j668RKQEqfvFdRl9pHJfRXK3usxFpMq+hVKePLbAYHO51G9
06LAnQxKaIEyrTAMKrcLvb2xFZsTlvCY/N2i4j75xXrmrEUv9DAA0nqrkmnMnm5K
+KHxdVxhUGeVvSOjD8tet7z4K0aT9j8iYtwOqIBUMhL+pOPMO12ySNRcULnCqxp2
/l9osruwUnFJfZwEew2D/u1krWXInv9a41+0oRk96YRETpStZnCgf/YcGC1lQuUU
IWqmpDsEvet9rSmjMbYOS+w1c/ITNZKta8w8H7NlG4DffS3dWxkgS4PWMiQiYwuU
XtRfn5Ru/RErJ6mZVhASrTPoUabxO7ASlWUsihPvuIOz3CQIjNeZSy2pLXsmOBvA
kBb4Pf3yr0Gj1pzjNNaoweGTcz5ik0wJ/eOIQcdaZJShxEm4TzgRh4wu5WpPfi/3
MAiHQj2EjzGWLNerfC7ltWnBCQhmzhywKhUgjTxsiUvsaqaS8WF0zNzYrKO/Gr9w
c5nO9uBZ59pUU1P2bTgtxDW1sRvcLFDNXuPZTtooFB+6o6Ur2r4O98++EdZlDn56
2NJCLpWPK/vjqigamOiNols718hdh9yp0RKjsmY6DJ8MoPc34RBi2FoWWFGHfieM
agMpcZ7YSCjCjQJ88ICP3VbtZb/fUN28SKwvB09X4DOMs+F0nR2rygggpHdtshU+
1v+2L5ofDBzl/0tF1uel1S9T3r5etPZBcV1SX1tNanTAO+/wfDgiz9VTO29BWSki
yKSzrvIbQHg/4HYIAi2HqlDYsZbDvl6RViK11YBtWfzg9OOfIX/NEveYLZM72ZRJ
78WAV8kLIaHPJ32uemzNsn0uDzaJ98HuwfeqOcLuaOSnZB7toNEuQSlGv4/92vvw
eUKDMsXNcHHJg52442LiR/yJGLBuE2xSLT+rZ+o1pheHSE0tCKWaMGvzSeGHRpNy
Yr8nqjJstcTCsqCTa97MIr/48qaC034P2o1kGgjBI/smfHyYG8F8cy7pNWd+Rr73
LL5IlJDKqmxF4GzGnPrkOtUxWrEXp1neDEyQjVftNaKgI4HdjznTAQq7FaF0PALv
2KbvqRjotqyPfDMSuX+l51GcA2c3t+jIO8efyBXlkmTHaFb/gua41yDWQPe68MFW
JzRrK/6ILRuQbfxObZIK9vwkPWQ0qIG5YWoAPr9AI9GtjhEaoXhHnl/ll4Ct5Jxn
WRyfHkfgkG9CblZlr9bWY0RuUPJv3+Z2q5tFT3LgDmqzxknAy0eWKmcOFup3L+1J
7T+PpMDg26SblKJlD2eUdgPOrJi/HWLsLyORiZrg1pfE6hGmekrqBEF3pOHpsltu
yLa+NYYHozPYWVSYDc4YABbHzmjG8YYGusc1N1ZtE0aS6QELZhLm3/yBWrj2EtrE
AQFv7NLqFEHO3ZUWp6fzRlMsKjpR6m1nZ9rXau7f0ackFk2tpfDbIpS/Vqz0sKGY
utPnJwjMfjKTpp0VnbRZ9nFIOexs3Zy2gn9PNal/ACAxyBNK7r4jVwPL5X22FpZ2
duW0bFa5q3OYcElrx1ZZldcgpNM7kfftXmhrZeBxtFaLY2mfoIrrxM7BXrF8325S
cVDEygSg/NOT4SgezOAR2uCH3lOIB/H4uje5F+3qMsGdwAVoT26UB5ktCq1MSFpC
FrFkon8pxAeGSoDU5f80XCjiJJhDs72M7Uqb+JGsJicF+1bS0IP7wNNaklrQh9Is
BrvV+haOVL3KK/JDmRg8lGq09jQfTm6XnYNl4X/k5xrVHbptJGMws2YX1aqWHxeo
WShFCMmgmn/oyt0LVIl996AXD+azzfzrilm3raqwLALBLyxcvj+oB1Llv5GuhoDe
vLCkOUa3r/smBe3sYVlILiUkzblZfpdxbAe5ZAiigzzoOd1EDk3fwdxWizAJ16s+
ken0iQrErgj5qdhPFQa3R2d00Syyy9+CqAilFjQz+SwqQA4P9QC20vag1eRv40ZZ
AHttM4jlQ5jFG3lAVdJMHASVD/CTEzKPSU/Otzcp8oNcNVwHA0ZW8HSr7rXFMZDQ
xtoEJWzQqpruz1TroHLgnIkOA/o10FFrUNXOIvwOQKEmp8oie/DySHuUziaOjG9L
1jhppqCznHAZ8gCoiw3iUUBls+uzrL5cXrr7wW6NyYGB5sfL21v9eKirlWj9IG5a
2vDCI6O9j+U+0pZFQE+DjM8xaHCP0Y04wffML25OWNekvLUiAV79yZzsbw/gE73z
8p913vwoMsR9rdjrGjDNytqaTT14IpFrQgQndceaiRYeOB2lEAOv198A+6Qp/rwq
Otj/mAHTCeCR9d+4R9jdGvPuQ0BSKMZ/yN/YGH+PEQESwhPOvZepGhIRxG385AeZ
nsNiWF3mUnZwIZxibcy+xuyGYLbqagw11Y/n9CAE84Ryt03/348gTAfROiCCmhc3
bQ/hbTjF8W0w7hCEA1FQNx6CN/MRUsVhMOj2n5sCoxZb7bAErxmhU7qNIxKxdSDq
pxbk/XFJlsJvYFF0jIdKw6BhECfPvxGRssw8R8+SXgdlig/rTCDKwVrtkV78wVqp
HWScvYfASI2nMlV8MMKFGEE+++YaiE+DC8g4fjQMt2XYimtzaNI03A2eU16gEDeP
VkFdtty61tgrNrEVk9NebFIa5aDhECUoEXn/4lTJSVi/QafpYhhi4sHFitwajO0O
Bl7eVjzoAnuYzSpE1GP+TzS/FRMB8HbWUYygku4l4MPvWb8d3KA6sSlouQY0DoNd
asXJSYD1ELjBy9I+4tQoVzK8+TU/7UXhEhy0hJXLPsjTE28tRKbQmKhYkccQdbhK
3OCBwrsg6KYKL5XKoczyaed1wAv0QoWOvjkOyqQerF629LO27B/is4xmF/MMasEL
esEzr+yA629aFCxOjs5u4xe1qzi4/WVFYWGOPDgrk/dwUGYcxX9TuE99pkD8AaPk
cIOslBrW246L+1MMBziV3jb8yPh1grBn+wTBoLlhHYGKkAHD0Ee95is0FvOgrnN1
J5QBFDlpUiAM7Q04Ly8J148J56fH4A435UMgDVP+55vEOYWE8MRp4ELcFGaYJcMf
fffJa5FTCqTb9jITKF1cD6Q7IBcWh0KgbqaMJqz6tjKQ8j4MLq5itTSnQsvbJOEv
/8fCGjYqrJVHnS3yInL4X52l4bHi/5dkh8EA6Y5IdIUNI9JfdyKmWkX9myD7NCvP
/9MwTwDyA6uZMiH2sNSMbSCOnZYCUpOkoALngPXc0h2d/TaBoXb0LgMs1EOl3ApH
/oNb5ZIC1YYIxgltCgb+zUNQpva4PBPs4h8+j2/T8LBr/G9m+5AdQazEG72q4d4c
CbLsOjM+V9VHa0l8vQgUA3R8eOTd3gt7WKdd1iyZe4U4cIWeDnlom9iVGZbVn4ty
H8Y47Asorl2CpOlgHNqK/R8I74cJnorwWd1NsUz39k4NbD8hOn4P8nFMU7EXDfK5
4aybQjMGOh5BD0p4uUas/XUFeo6RHnxhLQjgvmIXXrBaJXcEbdSDVB3dPDGt2RD9
C1usYgUixkrsDXYEoPzn4Cm2Re5W3eFAUsY5uM9BwZpBr0pusDwy5tlHbEE4a6X1
kwwPZfSFVMOTP940YnlUHqGtj/FkBVZkgEiS2BDRtVhn4j7cDP5XkVO5uUc8huzu
PoNIrfbM0iZxG5iFc2h4cnvZ7KWz3LEXib2HoA+h/Hd8gGESiDuXLdv78MxxiWgK
FGc4wPvyaAZ8R4f58piqxJv+ZtsAotVYdXCEnmQYOHlhOTkv3w6+a5XIayYxIBWm
fmzysnfr1xOUG0nVs3lb0DoQKEdJwVCF6Os4OYEOQjz48fhYFtg3K6K0tTFyuP4q
1lF+kZZsaQSCM3SLCBLZDl2VCEpNShMgCNoPFeymSVCor0GraYhiPChizqQn8hDf
MKqZffCOTF4xk3SrFx+EmyuVwuukUyAGp9IoUFmRa6CmL1rgPjquK02MNPm89GG5
4LbnrZ7jaoGOPukse3yzOK4QvbWulxCspf2lgl/rrfrj58FIcecx+MLa+/caxyuy
IBv8o3CEVVHtxsKTqafR+Y19Cw+vWbYLczNzOfqCG/A9YZHUvTf2erO5biCGDfB/
iyL6P5nOgitQcBjxbG1OFboST4iuS5MLarVsVnSr0XCPlNsTcG6noKY8shhOPPxJ
1OA11nH5ceizwPJebGfuWMZf1vfyQSrckm5U+rPK02pyv+SNaevRtThbkpRqrxap
rn9teucG2WcBbi4FPkHPJsykYzrbR9pMAVM5PEHOur8MCenTBIZ+9RsIPO9t9ijA
Z/0xnlFKqJ07vLufNT4YQsuZc4nUP6uvFmSThME7O2mA712qg7I+BZGxhuaLj8D3
Ub54HMDIRHtKGVRgBIZ1UV4MjT36qHVAKUo6i7fJOb1Za24igaG4mQaX7+TQ7XEh
Lah7FQAz0UGZXJwqPOb8f3CZlS8MU4zDv3rAX5c1bvyeS/CGPc5kVw7E2RTWycR8
2ikN+jz5b2DuMe4aHn8zCkFtr9+dhPQrzButupTgVbATkzf09VchQuLoo49L3DCs
vfd7fHEUVYptFBLlnDu429+SIfHN5AN2LovEAeA8fiBi3ju4aYSyspQY55ySEfZL
3+02Io7R9u7I3EUJKjm3K4bXu2H4VP4fvlAzmZ/9eV/3RgUZJvCRZK/cIfbdjAgA
rXycqqyiJbcxxe9GVePikRmH+MRsJoTgzHuLl50pQwAsNuAceXtyJmo6DX2iOPxI
KpgPcENVX4hqq/OjDCC8uZJxfVs2H171Lqr1ZWuWBIJ72QA7rmhPVAkIx1WCLY9h
+D2qPdJmf9NByRK8GCVLQsdbCyxbu5OB8BSx8hqpDYAtNK8imKGgvo9AvRpMQ2E1
dH12mmRAtRvu7ueWOfFwIfMGxAbCFrGwoggm9TxdhrYbtv1lkzo58rT7/fJeeJIC
NkfgQU0m43tMeA/zaQKJhjK0vH8RgOAGEJA0xfXRjEUsFPkJc0FrSq2MlYDL44En
fds+5JOkCpreN7dVMI/Mbjcu38vbvhXnMDlAqMulTjruLlOVXN2oW6NFmUEsJBs2
hGNVQBXUw3GImtyAx43nymr5ZZ7H49hKzZmf/q4//2hCZbsopOE0s7CuPAqGEQNt
XXKvWEpmznZWqzTDNXr0mxAcLk9qgAPpqXXYfQ29Z8yCSI15Yqz1JT/LfDKh4Fpk
TaKLC2WNBxAL5k9QA1ChCxMYHd5OXaSNnWeW4Pip94M4Hb7jz3AktBtd60Qn2FB5
wVJpSzevQKbOZ6PoCsJuVqhnFczIQsPfAmkWoht68Zy6+I4Km3tcalSfC/BiRiCh
9CjsQCV9/eNUAw58vRlQglRWpqm6Nr3kNvmDXKgthqgqBFwUHkDD+c9GEhRlXeXY
sX4NOhESr6oflfjGAvbV632iquzTu0kxRJy5Rfw/v2tuWapcxKcW6xaYY488vmLS
sfquLnU+Fb6vzDL0AAOI9J2SSM1ytnYdA3T9vCm+6ppPa+X5U5sRrVfDSXBlm3uj
krDywyhlGlTu78R28oshcEFxGBYAViCAKsYQyTdyISJaoIqojh2dTzf9oV8L4Ywc
bKczxBeBrOsHa/yNrSdpYb4CuwGjBwQ5t7rTvcAYiGt7QH3H8EB6KNLETEPdsWUc
Bma0pBlcbSiSeJfTFl9+pE58Yiap/pRScLsywCqyHCL5XQ5BaP2pcpgwaolWfoD2
u6DEisNrl7+vJzcRN/umN4Nmhjseg451ULhO3Y9oI+/SKSCXy3OE5BfC5ak4v8eQ
KNSne2wOo9J7azYS8xFGFgC/0r+cfCxpaCdFWZ3nOJSKr4QbcOi0x3TN2MzlTEpi
DtfCraOQu2ELnLfMBrobFenUuEfNgsaicBDTGhRvVmKbAsL2iUYMa323YHnqqUJf
rBPjLJ+pCF4590qA2P3MqUIEtnEU+MbVkapJHuTMEnDqt8be9sFBIu3u92BVbMwt
9tm3YH3dDgRpjVKjn0O8yhqaLAMRW46MJ7GmhpxqXjaoN9VGCmsISgcoPXeF2CBm
8EugTNBu1OOHn9lnstyas7m8vcHMjaWt+o4lFDilDnSg5xM7AzMQEaz4iy+DdNBx
fIQOKmkNk0XqLlnsgzhoSVXfEjj6jpHdcu9YhiZr0UsdborYGkYNSOTG9cqJ2Zl8
pf67GOmsEzFJ6foiSLJFNGnnzNZ9nBe+OSRkBylfDvEHJ/d4TjrzK+sh96FmxzMT
iht4pijBhpHB9pmGJH14Xvrqql+kJqrVhQTlUbcWARPqSUcvdJqlNNjmdaJO+bFz
0q4QNcQbgYb66+B48jMSTmvUAmPfAg7gi8HKmgoUikiKrcFiL7eoql7E+dnxia8o
nGO+kcV14QZlhTXV4+hBW/DuKWZb0a5rknkuhVQTOWdrWXdOkVTx+50f38o//giL
Y39Py4wo+q+4Jqsqu0STyPShHOlEu8u9w6x3Vz2xNsjYPJtZa9FznsByOPx1BSTL
ZE+JXYcwLAb/4OFH4i24O1B9w1WZE6UspSBDWmBPOHR/ooMewsLd7REthqOA5HCQ
ukiYof19GhLGkgkdJAV9t5PhsnmdX6hjuR2ftcw/2N5X81LiQ+u9gecZ5PXEsG/5
0PEZ7wnBAYWPM8SAURI7569CYEZsbfkPWpiLJGbPEwsTgJeYGHKFuApK73vDyBWX
KGI/rfz2q6AgLzX13utOt9pEYanxD2XWLoezljpdg0M/UODASKLQxJkGlTa18xfo
lhPfhVyXZbj/e3/f9Wr6y0Y4u70ZNe7kk2zJ4g6YKwAKDhT7idJSPrVv7AP44s0X
RFZ+NTfWexjzwqHafLRRJZx0OqHoRQD+kxFkGZ6Rv8JE/k4FIPH7i88DTWWg3Npy
LErqZBfeAHeXmc8h5yd/4jHV0UsgYld9ZfPfG4p4O1oI+Mo0+fQiZ0sAkCmd+amc
2vN+piEsXLmlr9VvD1fLrHUNSRTbPGxJnYIGNttQnQyYbZ3OyBLbYFwjM+jvYLHP
w72W0Q8jpLbromJGfc4CmtenqWR11e83GamMXDDv3licEYkxe7z9jSJlt8CqlVDY
JF4bpSu/T1RGzPf98zhmwASSLSIQo18Tf9584NJJnBL/r6NEjIbwJyOjBJZnWYzf
hIScv7ZNiDpdY54abu5AtcFZoWaNeicYtVqQ5i6Np0VUx3xzGVApAv1F/6XTaNOl
hW3mc5eEZl8wCoUKQintXk4AsKKglQfTJRNDlnBk++xRkaF8PAxNqAIlnDiftqAI
pA+gwlWzP5pQCuH1ALVwI+kcXScuw9H499NMHOL+jqu5g+KrdRuwap1XeV015m8Q
J1XeM1+tRUwLdn2qaxvGlQyssMgcGyJHhjQWbW5FqhlRIKyVs9DxQfmW+oBzR8BG
EHmrLjbZ26kSX98G4xgLL2ECfHl21/yQu5kI3C81j7HoxTICtX21HGJDyugq8rNr
6iJimYQChxxUfUKQ3XyIyp+swKXWvZBY9gs9F/wIlhQV1OLpyRgn9Ky0Qtzw3geG
YDxt9hZGhU3Q0GuUzUX0EiyzbRvjkxuAqd+8w7AoGE6M/AXx1iCohM2LC5K+iJjD
RCofaMwP2Qwq7YZ/tfYjfAn+jWFY4UBzOLKj+H8Qj+9iNJcEhkK0/9e9sYnlH77/
0978QZdzPMQshmrXvkbwcj34x8/ocDzumU0QZr0lRnQymWcGykxCx69TE0Pz8KD0
IWVFWyJEa79CQMWBYPqc0qeDDnEieZHvgfoiQwkTy435jZpjjGmwzfMFCg3+FJ25
wrgUghYd322ZMdsarjscXPRxrSUTtXWM+o2QxOiw5gdFcMVebySlja5ILDtjcUpD
QtWxva31CXJ1qylQ+OzOAyc6CjjD6aTEyO5cg2Pqyj9f836zb3HH20m+gRTzmIfi
VDCA8Ya5cH6L/034yohlOb/3/MGIs56jg59XGhbRyMsG27T3JEYz79II/d0fksNz
1eUph/AbgEXmwPlftiqGf2u9g8AYGhzjaLM20KMqhOZv9F0awwW17DKuSQHDfmkk
hA8CvDhsovOOyfA/mNkZGiTHu3ga2YOoVFGhqhHJ2JDZsb+sFoTqYh4bqELVqg1b
bYRLIKQpS5bqemLLP+/vxIUmN9GrNyylZkQb9fJeRMnt7oj1AagkewZ6nIPXa3/N
TGXfRk8p7ZmWusHWTyFwwIU+Rc7H+xIEGUH38TzqcT1VL9UK4Kg0zqIvhemdAZcZ
LfTqqUUmrU80k8Nfr4+LD/iJy1jgD5vYs4+L6TwcEGi7F3RLRW8aTah/ZfRJPq/Y
4aFtsGswDtwhdJ6epfW+G+TL91jl97lN39bj2R1ZBPV1AfiVTo/SXAjxoAgThzM2
cDFqdOx5ne6NabjH6QDU4ztIDhSeaox6SFfgC6kqMqSL8Z4YU/fPw1d9Ijtv25mG
QdIcnMZnZ5uemozV1CJxKjy1sVIpYrtJOjmm6p8F7/CQX4MLPJCktHKuI4WmtLDn
xHgev+utv4FyeK3H7TRrUNPfvFvMJWwzRLQBgJ94dwG2G12g6WehZ5mIEzzmck5D
AP/J00CEXwHc1sVXWde0dbBpppnR0MwjRUC1O7MaQ+Wle1qoiW3bylb+W+gV8xC/
Tv4d6aproQ1u0R0Pp+VBdJMFeem5abXL2fDApZCiJH46XeZP5FgR3kKB9ooqhaB9
m0fIQlYcPWWWJ5TXluij76R6VU+7jXuJHjWSnSIkYyzGWVvmouDp9ErB4GnZHajk
WElrN7BSyuytKGiK6LCXAJ40d931J5bnXvuo29n9OHDGgvbR6HzRcM7/Cl1R5BfM
ttt9YPzEFZcAGVvdah1mkLl0mOwsnmaVfU5F29uG/z3oYfjC61ofqvplwIyyX9ch
1UmSJwmKNNd+OqJRl433E+KsGYBhCBXZ87eRIkiYf6htIaw20pgtZ0DJHT4qeHQJ
6RhonlBQTUqzXSpeWMvwPUgkXQbxJux2M9Wea6wng2C4SAibc/bwRIWxWfgQ5gRB
y5egra6PGQH0lmOHDFxXww8eVSvyeXo+rFU7BhA0opRq7ed6jKNyfZ/xrKIDly2b
1jPmuUCZ7Eo2jVUiRZjqNPV5A+srVZqpF//vkNPTLV+xl7WspxcaAplNJVxZAQ0H
17aIlq4AYcW23B/+p4PN8r7QzsaTkI8jZOOCibIhBmsnAEqLEoKOnWtKSuvYAbDT
3gOAEIJG3aPVdiieBIS1f0FNmv1Ryzvu9nlxTBEThBG3rAWUuuEwsoI+1GSpxdFx
ZJYy/qeUOFl+OhGa6+eMXcZiHa65PvpmmwtUSu9MHbBoxnLlhdx5OpDdqko/AiMC
Pld8ih5NdkDYJeiYMIWE11sNpgPnvG3kO+ZcNC+aiyIpTtrJ0zZ177ZM8ch7HuxH
66WGbiVEp3UNlQ12LT6Ay9BhoILk+OVcNN7oOS2jmIXGBaDRaFsWn9ezmwCds4Ul
3HWeUGqlJIaIWScZ6dGrqo8SXn5Nnv6gZgwiBupOHJ9YyR6O70b3BQsbHZcRB4/9
1iN7EscQ+fvK5RXKnOVHYk73MYAIrIzYMly1gXT34QuF0KH7rBBC810UxfNKwKLQ
5El+VvJUpaZcsuktlGm/fUMqe2+xxA4FJWg6f4YG/5/zrpcRdWu9HtLsv++9cR5u
6m+lV3LGtUg8v7rnsHjj7SGtFe2HLrwffpQnpGSt1G8KMizHqqSK9NS6JlKLBTKs
p30p6/RaH7ubZ2Z2k5wBFuar1hjK174UM+TxbEmtddljkt6W4HxQU246b2mWp8H4
yMGsn25lizT9CyFc1CfgK2VIT49+5plTlUQVEZnlqBbQVJRbOXZrEtTElLOz1Der
yLVWCKWaMkuXoPk/u1Hz4yHlxo3g4+9S5X67Ni8lGLMgkrqApk7Yb4jakmSWTgzc
kqfP62P/6Cqay6bg+gzhkye0LaZiuW8wqmkOhOEKC/HsYAlJ2G0jlYq2wUw2pEo8
TYIMwKjAUSva56MkceQzqhwtI9zbuJdXzEt/uuPWvXfqJzXHvOYsdoZtV44rC7yV
e2KnaEuE8bNeJdb4QImMTc+T+14ZDZdN/VhPvDvQg4UjMYQ182RdYEqqolcYTj0t
1TbaYNdP2jfOz7YCI9XxydRTwOEbrChuHrLqlPDoz1hqxtI1CIilMQJC4mpF/pgG
SbaU2FBVRrWLlGD0/6l2ioUl7d1SjfXINXwopyZg96WYidlI4ZjrA6r2pBYvabfp
M1Ziu7XPinAdVe0Ynmt39YquOKCQJTzX1rWGlj7yOoKjqgAYY8T+kDJAXYXB8O9X
rSwHt/RhVBc2brLnvHLcL+LhFvEeQWF3u6DLujAjNVIZFLvJuMdyIFGIUTXbbklq
NSrtyXrraTA21koJx/kN/3V2DmBMmEPaBhzZS2pKgnLM+NIK943hoZhNLPX/OcCC
ruXwuQFfHHlcpFErcxYG6zfItEgv/51AmOOkjsnB+aEaiFmLwVAtzWfyP06X6Ji+
vKXP+DwcwLNqnntJ2llk8nbh1h+Dj/RO7F1Y4PCWPrt2vXebv6idmzx7eAjevgvn
G2iQq06i/Lufnv2EYn6IX8/XNNOpoJmDT70KnbqZr9t4yAqU5r44lEftQdxb+QGC
tjD2zM/DJSFmTdiXOwjDQrVWrTVYtbYVBa+U5NyXcBYGVFQoVIYcsb2v5Jdhp9aa
EOWWw+AREXRI0OEE+YipTdr9tUO2g4Fn0C1AQjR0o734bQqZsywGIR2ZKA/j7UKd
D3HT5zDk0rX2Oib+/BbIdJ818lIu0qJydtb0+XLa8/+Uf+Jt2ASjb0mXwxqLWcYZ
dL0kSks3NQIgrqYeRVr+dngG8dIecnvlMP8e1/O5wZjMpfZFTHI+joju5tvwvfEB
0VQPXZxpeC34urbLyj+lZJhEiRCIOaBIUz7TEs3yYaF8bweWZJKsBMmrqithUuaa
HyaHhPh/CGukDGlPMP/Grc2uvMsKoFnRchXSYgkFzhoh3J3xaJmoOZV8U388+1RB
gW0aCRmSaIHlamK6jxCUO58R4LRvX0Eidb5b7/A4cowotRZGjpjuOB47hp3PO1fz
q4ue/JjT85+2euDzzZFl2pApz7G8dMml/qEUc1ZdPmpRUfGFSdzPvFyLZryIUrTI
CoJ4icY9cV8wu7Mbw2kVQQepC1mGZnkgpjlaXlHG7clcxOxAZONFwzBbImFhJ7B5
n2KfHaDFQwYxlVeQUQpn+E7e2ULMBuYUau1eltfVqUXboKxDD06FWUhluPsSkBEo
yagIE3V0R9O2/ytndSDSyAP551+NWrO2olg4r5yExa9R3VGeDcbm2hDAYzX+Vc9j
rcc3ds/QKyps3YOKPnVjDaxu63ZiUkHNBCHVEMDrf28L/ZfuqyaBorbaLA/REnBP
QuvKQxvgspvD0l4sn22LvLmjv0GxRsT1iCbkP6U50NKN3pgPhMt3j7zzy9itGIl9
P3//nI/VrcZ9x4IgW9jAoGGrNGIrEan7zCdnbkeUVGeINfrXVMGg121DBslKKO+8
PfSeBMegvWnYAJMWWAh3olrsZg61DFdbVYOBhDt7Y5lleVbirBk2Dc0MZwOnRNEj
haKfjfZKian7cbx/9cTntJXwklUx1prg2g9+2IJKUZdOAhumZ4toEvCc0oes30pJ
V2mFt71wzapjOSRfu+uvqzxMp3ZmSFWR8i2xeQU0R3hsQqu0QEE/uWwxDf2+dJOY
nnVjHfIO4RRhCLl39TP/pFyNO6L/8+j3z1Ypb9rqu90+QinrQmViNs13N9EXqWEh
N9DaXWCCxbC8LCmm2mHcbdtw3+SgLsESSC9jHeGZ5LH7a+TMJkPJ/ZSJfZzCqmof
NOOLysCSo2bW2akrCkPGf2jYh/bjc9e8uM2r/6N+7NBe8urIJIc63d17N8IcC7LN
gaTP+tmkuPjCn7F5sdz7xYIZ9WBDD9xbNWDnH6XJSZ8j4q3yVHqq2MkWJWign4L5
Kkyxtp2L3qX/UspwDknRqFB4zGX18ragzcqdGjem1UFQef2AYQU85u6hw9/S11Ls
ut4IuqWs5ZfYqzg1eSwsHDLtuWJAP7goVK66iksD826hhfP5qO3R6gomaoo1eefQ
8JG9OkyDGxoeoGbA2SgWYRIItmkv0knmKp2an3eo9S58hio8HSZUR/OlkhR6zNfB
YAfgSFQ5mLefEBPkS+I8KutjQo6Yw4gARiaz4s+E2lDlo1+G8Hszp5KyRoUr6xEO
/VGm0/wglu916INUojqDxxx6sVH2iGmqeaxlNJoSLwaGxImhC9Xu9b+yAjnN3+Vh
CVKCElIrG94Cio4xObine3UAdSFwjXO9J9TMFxawq9ewujXLUTKMwDgm+jvbTfEG
LlHksk6gzsXnUI74R4nkhdJHXjRbQRM3q4KAZdh2BiR8i/t7uwl2Ijqga3UcfrCP
gLTDFwUDuMKZj1elhdjPgKz2MToUVtZvMFi0yhF4f6gy7Tso6WMM/pJwnSpazE60
RkBFVayV43DiwrerTbAEGt82iy1VM2E69HsrUEni5boJcetedg3uu3w5oXyRt5zf
wVDth7KqBuwC4Ijc7ijpm5Yv210sIo4lkzNHDzlr9d5GRPQ6A1QWP6Mx07se7HUz
Qye/LJ1A98/wEIiZPUMPM208HHk84rXcPBkMCKnXO4d77cOGNKz4qxeXGgTOZrbl
L0pDHAbrs0prG7/22En2fw8efsrAdD1hvCybtD29VfHq/GWpJjGe4OzpiknFFtM5
ksov/Wm/R68nIG1mx2+WHycbWpOTCxjwRZzMYyiMhnpPhY3Tb3U4D/TmzNsrVN7g
O2L2e4w/g/Kyx5rmXIs/KqsethnJ6mGCE8evl7QjdVH2AlwCXSgmJEPVhlsEQi9z
P1qUNwXA3lJhhp4SV1yuctWN7kZ+eEEe1OXbXVQGeNVIFJDF77WQl65NPmeI+Zkj
h6iJciztX/CzSRaZN1y7WWZca1HRG+z4MfyV6Zf8WvI5vZQkW5RsU/xryqe9H2VA
v8Hiy0Qb+Rp5OZLxOiX9uUcmUBk3SXsXS+1KJJoL3kobU+BKaI5NjAbwi04nG99Z
V6sAgxSM4ZhvAAz9Dgrd0IFEbQDlbStvWT7Q3ZewwFy/z0rUnrRi4g+b2NHlx7eo
bBwF8Uv2TYk6/8FiuAHC3WXplJiYceDIoSCA2zI+VIG02zOMqSXeKe+bNkjL2Baa
QeQnGZobh11P2ao+dblReivMq+XTz7XAhB9Y9KXdV6E2bCqhFYpqiVOzJFVR5QyF
k26aYI0YOKSBA3dfFlvQVqWRA+ni9byLJKl4fZVJB5rALRrx4/UF8XN4xUr+ZGJH
UK6v3ReaVCdXigTv5pDru/eiuMDZ6LcjQYKpdWaD7YYZJD4z5I1UT/7pv64vtXSU
30YEVc4HTHhntHbmvCgNcRUeGtb1pkFtLnOSz/+//84RySTvmpuN0IGuLLY1kyFz
zo83hWWmv9TmEKa5HyV6+64RCAQha6JeBPguob9VieL9YXSUxo8LlAWPz12tGTJ9
R76F4Bpor3BCspJoij677ql2ioFtHk2dqrZ+wP3+uKsleASXppJ3+wrlCbEO/hLt
GVA+TdsM6/1ZCDtFwtlUZggIqrPMMhFvJELHErHvqDIxkfNhb1FMusMTAYFZP6PO
uNSd03T2tQkfmnJ0fsTT/GJiVtygbUWRtQ19EIaAAYPDBSGzqdkQMs6t9BEsGoqF
Z4Jg9WUKC07VfYjRaU5k9omwOt5hzKdiB56/yfQt+KHeVM1jTg7r6OcAMCaR6pr8
NfDZhs5m+VOEl50ApT9ATmv3kfadoQT1Dk18uQapcinyIrPWTeBsiCDIM8Oy93wb
4TBVE6i12YBn3FTRWZ/nDpaBbn89b0xlcvVjOBgCcPfFXOmWcghZr/KqYHs535MK
UjPRxK712YpQLw5CLP4WaJ8k9xGDCMMNwjQdXH+sSHd6C5SAq5v+tsFLXmPSBcvn
VGORK8c0EAseRUoO76fqRRYCT+aNfvL1Wb9yYTtGsGwhzbBdHrQcNnGfsIszm73a
bS+2MAVCYCtPXT4aPcDthqZjUS6ugACjKZ9gJ8U5cQhTQOqOATz0LBmblheMcOyz
HhaZHIMM2e1tIjETR38GId3UDD4kICI1WiN6JAOoqxgVXL/wGGzOoY1G3TJ0YvgP
dv42A7tyEa2Mf+7KFxNcpXpplMXEjefZzz8egRXyl/FRzGeQ9ZJrWmviilzhPCzO
kATqKqWkOBVhX1YWKrhlfegP6O9riiO9ttSwEoUmmTm3sXaqPwUnq71Pj5CFE+DN
pryAs+bJE5CxtwFMIZJ0wvSLsK+L9FF2ynW/wnnM8Leg+UXU76TaWSrr27tqIGD2
lnAftnhd3xYTO2DFneQ0sXZUt6+QJn6dgEECb/GjPg/1P5ZAsEI+rYkMKpaSK52Q
yfYZFPvAHxpNqHVWob16P3191aDe1fjUGwswN9hCn6xCN4zg7er1QjUJu/K40Gyv
CpQQjMIaP10AMhguhlQZal1hy7olpBgzFSftftcqc056SHAf0r3w9hoShGVgu0XN
yptNFaBox48cbggySatIpB50kaqj9ttntA05oDEp9PClMuQvHtbeYJ5LSZh+h0tl
2n4RSdMvePtr/u9rFkgCoAZMjEQbErwHhiQx44fdCUJACsZ1F0DasNToOk+oi5a7
/N1A+wfsXFsbDMPntolXPPl68cRPTKPeoGZP74RGKVe/pQLozCdOE2SBs4cX6Z18
PRnZVNWmPWnUztmT12vI/t1KB7Ackqpq9BwbmTgBuLipgNrT0JrlM0GdzMUnJb/8
Wg0/hQY3M2VpcroxFshEfyjaj1R3/3iCGOAkPXyEoFRSDh4I2JqhycGeRtJZpDLE
WG/JMiejQPdgm/5vQjznby5eVRIWkZKa2BzmaqXkTe+M1yyl6LMVAyBqNDTJvzGL
mFrHfsxZMxJNUW6YVp5coOeUoBj2LleoRSq3hmAlQ2fJlj9Va1dec4Mg0eFiAxke
57LcOwfX6X+UjEHB9/KPYtKCZTO3VHRCJFpSyb7dHdjua0J9uSU+0qsMh9+44Tks
RNfP62FoNmsYj4ljJCPiOhbBRx8e+dgFeMpYb774H/b5jRGvjbCLniWfrIJZzEhh
674tZzDPUMP34AGypKdWKLFQKf/yPEW6UKsGQiumqgkkU/+l2OAVHptMZPInjs4H
MFEQc9YWQqYuIUqNH6Giahv6ysEuwnK9IigXGbZmxJb3BrUW5ifCsMMkBgoecFmq
3HYVE4KUlIMxHwLaSgGioHcOA3Q8WR4BoP9tmTMuP2JID24IQb2Lm+o3t3u6PWhd
gBvRE/LUDoEaIMNnJERXhAj2lemMh7iMxeiSsSPToW7e7sTSKgrkUdqsS5d1CMQh
w4z3FCQFqgi08dE96f3iBWPckaDIRsRKd8ImfuAasmf555Sq7mlt5uy+SEKJmrab
KgSabMURGZO/jVRIM7bZFsGMF20Z71FCgVEKQC42NKL903ZILMBtVthe5DBpPm6z
n+yJt/KUdlyoWzdIsYW2GQsB7GNuDcUCpoAg56yQO/IsqOvYC6GDvhV2TF58gx6G
kgvA4+OFwEDwMNrafZZuuuF1cCc6URtr3CHOVRbcynk+NxyQ9c8rdm27R4K4YzRn
s0bTq+Yv9t44ACgT5KF5vK6KgFfsM4F5HWXsdCHTjeK29irjElzDB4MEY1iEaGx2
6DPlHlpvswyq2M2nI2uHECDh7SdXQr2R9aY2HkpFLe/70bX2YMoViN+Jf2lxzExs
ekxzM89JwRRXzRNtDuVZ9UhHkm1Ke9FG4x0URbXuisXcXsL58fBcV9nz6NTWq1O1
25ekgKk+c4a8RdDLExPTLvYpKfd8abp6VDJOk2Sa4mSC2ojkKj/AAoSDNrOuyLGH
gmcVxVDujnfSWUSDE4x/ky1UHrXMKtSZQ7d8SAeH6BvIT+M8MLSdIBGZWRwNGv83
Vuak7SSeQiEZR60qZKaoMXIPxumDj+HCT384JoRV0PWP0e84St4/xwhYQRFVoTgU
Zkj80+EcOjxv7a+LKN+GNZrtBb1ttwDlwod4cmXqczx73z+/fFGAfoxYfq2cvTc7
vEgWDVZwLPJKeqonQlYqDIamx3CDDQyMJADNa/9+GxU7kMC7RXXL06z//7E4jhDM
lp3aohzxNcIUdbNpFR1wnOCg7cRfoyLhJqKlzUWmA6D3y380DbOYmOvfpg59ttkq
QFqD1m/nn6SsmmKYfkuSrlSYkc/rnLetESjhXNZftmlboIQ6+G3Zt1C8Cbkeokx+
T7tgwFCmXrqAeDb06mvH2eRKPTLyORgxb9eaeuTYc8RgDIBu7RI/VSOP+y+lkhGg
1v4+81PsvaxGUtA0xt3YV5zAM5RFA2oTfiFKTch2sVbNFSUcm11yHITXAb6Avkut
SwBww4eRxp+F/padaImi2XP7qOXzskdaKCj1gwBcP9mCxOHxkgyFa3wIA0a+ZvXt
WYiPZ5FWwSZxBkrklqe0XkvvlhqIejOnGCh+zHACRXajT+A3o0+SZzjCqSGgw7sZ
U8bFl1udqjaYqBXECn3Sfg+2IuxBq5LQTgno+vjeYj8/ShSKKG0eccNNPnHbspLW
qgStlhPpIpbwcI/RF1dMOrNUkU+WSFb2tSGtqz7YZhJ6A5JiWmNG8I5OxZ0EIj/v
Z+cjFxbKlQzHzGefZ2eZ+Rm7orLjyH6MXH1baGp3MjgaYgh3swVtR56WSVJS/AgT
Ulfn+O4h7uanYqw1RK5efdGid20K5WI27vQDzQk0xensESa80FuH7+I9jj6c04bP
TtOEsQVVU5SvDd0TsarsiyAffHFJkQgX5/E6TAFWjwWoYdXVVX9cT0jzA7gMKZUu
GwHKJFylfu3bhgWMCdp6aR62PS4/AUyDsu/jNUBiNMAlEC04g9x+ZbUszMdMSl76
aH63Sy+zfc8m8pJY8Gz0mV+n/EEHySSTZamk18qX1A4ycOZwdUSeBKMFh81nzbed
u+ZF82/xZYqaP0keBP+OC/dSYenUVCMoazocZ0SnyhcCjD1e0z9E+sgCoWY0woUd
ndHvx3T214uyqR/7WKf50IqbUY73F5o2Qh3XmeQym3Kwm8vS0ohVBDZ6Ruck4m4I
N0Jsxo/fC+CGUC0GKV2DEgbKlKp0U8hzfNvs+Miycechs5XR0TGbbDHLAWsLFzkC
MB8Cp6FiBbrnPZ6LyPKWRMbMlrF8E3IA5IC0gWZ6/mZkl7+3/Lxh+rsVFHaaE9Dy
7lKM2sr0n+DdDDN1+ioHqLb7TIurp+EU8jX6MeZ6bAJsZRAS5i8ipNmgJ1FP+DTY
G/4j0WkYggN7ehqnKn+Tq6Ye/5QJK9PUje1ZA0ZJr1R5iinGKQpo7kc2AsY82C6z
n0hjE102Xrb0M7+DGPtMRPmEreVT79Cr9q6MBI5i5p3Tkak95jQ4kp3LasE9Yov5
m9NfYW2gZPbPSE1C7YhiLukBEqRDrTX9LpfOd6ANjz8Wd8D/3HfK1ZdcxW7Kows9
QKvoUwteYO3jRx1Jojem1JsoEA2Hk4X4b+LTLPA4VO8xZeT9h1VgotY3B3z7U4In
utWUSCJ5pn0fhSpXDIkl4DxiUuK0wW/qh4etkSWjZcQo/0AiEgsbhVLFjTQBPnEp
JKWWyloyz0XbCREZRrbESceJ8xsL5BhWlI5QxLmo6tDUdHCjuIpgwZ1LRUQKi0G+
FzywL1toUfpRn6DB1A3gwyxvq231wj+BJT7Ru47b1V1POXf+SRJNJwtLqFI9aCck
PnoVhu3ku2N7WdN0LlTcA2sQkepv9Azc7HF/nx5oBqjVC/2QIu0jiCngvZrMrWFu
g0q3pQEwH7DOWeK+jhARrWXyAFjvzyLS5dKweGMfJOJ08uKq0GCbIF4bAbmT3Bdq
WsC+1uinpz6Rmx7Xdjh/WhQCtqi+nF3EWNfUomL7JNqcrVcgi2jgARC9rUl9WRRE
MpRBe7ceD1A79zy8WLv2r+shc32uK82Xp7NvbLOj6OqIvx2ZqZeUjgmZlVkmWtwM
2Dno+0i4WEs/A3oNcBPtPaWHtPjd0m+Jf4MlgAjIOD2g1N8WzxwGOm5Ye/5aU7FT
HESy4Jy3BmhOWEimuc8gRgE0efjewWQW0dUOc/eosCCWMOFuuQ5mhkzPOKsuFIKQ
BT6wC5onT2tCYaQKI3IMjQTvwBs1vrf4PlayLxF4k9XIayThPp1lXhLsocsQXU6O
3hchFJ4bq1u+yx3CT3u6KBOxZVffu1qaiTByaoaMF5lJ5zwSnEdStV3heg+Pe6hK
bUlsPk43atcXTlciXAJr3Wt9oXOOWjYgeyErQQNHyNEWCHcAx2qIK2Pa0VVbphhx
l/G+OjFRDu5XCLftf4FXOdo66In4VIuMAnoL4Wx9nbI7iUtZ2topyExeVz03DyBN
tiGdumdCu+6+Nb/9WL3rzN27dCUF0Qsjx+eIsJD0ngUUzQaiwOhfY/QMSOkNFT4U
V17wuREF1HFUf8Fzb0ykUfLKt/oy9W4/36LgjzKaK1fNAFq6XkThsEe1VMikE33y
DqbXlJiNMUFtEO5hxAWXDZcyvuJRKBj+eXheAldJKidgP/h+c/YzdMR0i2XNTZPw
nGKkKtPmJobKFWCkOO303T5C8zDZ9AdYbghOJZnSLPw/tbPk8UjQx11N5cGaTS4I
FBJNw4ywBsCt8MUnTJK/39ENQRzZDj0k/6+qmpLZk5Yrzgf/WdJeWQtphyMfbYor
Alhqynl/T5jc09cOTEKpkZ6BMiPd4xdcm6mn/tOycwEb/GuoG81RwvNT9rqb2Ard
SqFs2HndvVuk1HwbErRo6o1kFHc0lR+MrqIdOlgLt7Fn35KojFkBFN/3ueI2OD6L
RGEVNGLEaJEohOeSk0r71G3ChQQmSr1BY3mHF1DEGv1BrJG7yR21RGUT8PlO19CU
comwXPYie2/bJOah5pK/CBx7nuF4dQp+H5ZMtIYJHqN0L0JVPU+tVE/JUKa6Nz/S
o/Be7EsRE3ulAdYrn8J6vr1teC7pzNmGNMWlDq+/hdm+Da0VpP3XQ3TDX1Wl9vtK
D+LKkNJyEiDugZY5U/xvJNi+M1EI868f6oLis9LEXUWpeDL9QPscN5nEQczJvRX5
v+Go9BWbE7W+QzqnnKNREcVB63eaiZ5kZ9RhvzW+NIwVK45RnKJGSpdC6sS3f7/g
oo3kRycQagLoAQCvX1oBCiM5O3PfqFQ270LTAOV/NB/r/UoadbxoYIQjT9gzOv5T
EpSsoLKk0fx78JJ0pK46RIgG/AOSG2+8rCx2wfTKk8L3YBgyYDj/I2GSKbBhpyoT
uWcFEpFNf9tFGNeY4DaEhlndPo46D9ieCGbSwus4rrBou8PKJwkwFQ9ol5v2YdEM
nFvNT5NxXAx3zvCpOY2JjszbRm6iHIin3t1azwoSxPZJflxwK4N7e5xNG135potQ
U4Ba5litWlkw84h7fm7vr5jjM6FDCEdt3Ar6/DHAspni6CM+W7F/83N8gtZYyxUO
biIUxhagOMhKilY/rmoUUAO+9TFcmy/CcQlX7IdT7bTxOkbo5Hln9apBoN6So8oV
37+d7AXj81d6q9FtjYgqVD/98sc0cEfGvwjY62h6pBYXKEZjT236TY32U8//1iay
DEIuZBqnfCsug4hPXLAW10GTTn3vOHwQSkA1fOmq/6NGTzZRNWyDqd9k+JT/D7Vk
XOtSlLWzHjYPr154K1+Nd0mGz0i5/b6CDjVnqIc2es3isvIzXUKSI7UPC4mX0tFV
mMdrNmkOKKwjYz2BkmUnuvYQn0MhpXTKNX9AUu/98DHv2Tr0vq0Z9WBodAwnFMSu
iLiZB4xyzVjJLV1iq9/whBdOOqLxSbuLaYeKlV87qkQnb7f6npKmcS/wlGgdIOY1
/KFOWuWCpXEduWsWsYnSqEBdC65/h9lDW0oTVrl8m652QRYmxkj5w11oHux0ILTa
SZPbyP/jysC345yR5nWvR6Pk/IsIODguNVB4C3/Fzgdw9GxZ8NcaNOcfFqJJKGVE
7DTK05FcKz615xO6skI67GD+2uYoNSk4XaqiaoMM+6Q2Gx5ZiFxTNj4TgW2lYqWz
KcH74KwN1ZH8uzU3soJhcNcBgqKAjyTW9oE5WrwgvQwbumxqq1brxy0+Y3v4E/+6
jj0BGxxBVIaf9vLMsuWhstol27jYnuoWB1IPNRgu5048weqkfegmrmuY6wfUu2Op
Sxim7zxCrGWzL9r39rF8C4KTt6SL9y2dMkN6h9K7CkM8qY8XwjRkruZkRrqXgC9n
QEDyE5+fVXvqws8qgNJb8BhcvC7fhwnwz2UQEBKWBJ02zbzpLfeykwEU6dam49no
OUAdGYBEG3LqW3N0ckjRiUTq3TMzlLzyojBq7wIRQ1EOQP7A0TQ736UQcOoF4Y4J
ZxIm2z1CavwvVkeXmbzDeJx0qR7irjl1wvmmrAdhKUH0IqOka/Pt96t6KCflEmDe
zQHRB4yd8gQNTY39qrO23srJRffUffyljqfyDQabVEu1zHcJhIlqlXTemk/yrgCe
l3oElTKgMa45JYm3PJTBtItUWsQcq+W/c0nsr19Ul4pTgvuQ2msWnbCxy2QXZEn+
R3RumQvWu5A7wOUBtCUiMukXlmM/qYt9X2Fjv5ONvHndfiZCeof2R2yFJsx4yDvL
Mztqk+ZXszFVOCEZBx7Z/eOse6A6Ir85QAC2qzNdm2vRcf2a2moMpfe4NuGhjPwV
MLEQ3q1BJjGPqSdd3xA8znMCNctoLxWaOWBWia5el4eo6t5kIGn34QI/PpgMGKPL
FUTAPWjCL1APYMPyofJxkQ3TQ8MpV/TKVIlrfjZFHBIVC2D8QTTpHPIP0M+XpcIW
mB6OG3TgBfnwml+8Df8Qq6phSFccl784CtZOhrIBihtk0lmoSTD7xS0T0kKtr5nR
6faKW/16t9KRGds26+xGTFJ/mpr1+GJVoX+vYjzVfv87OkOFqEnj+plIZuE0E1pp
W7bJI1yzPhHCWPEe9foMtSRglnIU+75FKoPlwykIhK3a751jssfErSXknuUsTwFE
SoGJxaJsn+OI48qoV9kNS6OzdgrtyI2MSPr8ptvjH1pQGQzqMhOfiGD5kZS/f2dX
ZuVoPDSwt7x3qUkk6Dfzt8JzGRTcsKYDgk5PCEmVN9TpVBZzX/Lv9eE7JlQzzsf5
Gjnum4vHHcxZB/eFYtxLsM8aDZlNTPFXi6Rcwsm1j+XsjWPxaP+O8rwHB+6KvlSq
vnQRkSMXmpprq1zrWlx3GcI4f5tSX/fESuE2Nh0V+bsxo03Phjrqyo5wOI5D1Fff
Uaqb0YID0PR8VNuOmBKoF4ZLfNmbRCpb1OzV33ZWbOf4gZCoiZ6cbcfWZPqmze4P
cyZsXirVbraNbG3OfaW8IhY3ytOvHoNKpcM5PWqCuN6pn0J7N3b/K8uqhZuwpNh3
T5OwZKyxqtwUUSly8UH8SJWzqVlnztgzr2XsYtddJq2GRX3SkeKUona5JYA0NJQu
/tzh5SAOoiUGMIPeQ7fkPJv6ahVCze1ZbGT5yvXZFxmeRv2J07+ePdChMSadWqsJ
dcu/g4XLRZBSSV5Oayh3cKM81Ok6PRBKkr5zUdJZNfemoXQPA/zRe5Wk4+lrJnZY
f2oEKYaFQBWdWPsPHbj/fzhqcIMhT5Jc4FwXqjT6XhehuZ4nqoKsLt5fXMnmuRdI
rcycU5wO1tcRnwRi0ahs2PT7KSbmL1zsZmhLyXMzE+yH44RBp6+iDZ3v9LkOaSgy
Qrnfd3QixA6cN7ey6yRNK7CcKqNWu0SVBFn0C3xfKsBHFS+GFqQkrB8R0o3MO1BC
AaAt+L0y4I7iOmSNUbrw4ALVpysEEM58Pz0GBC/6eNG+Nwu2swHt/9t5Yo8ZLkyE
YhjSU9eepkwBbn2EYfd0mbtFf/cBBhU2TBXgiiVjwSlyDrBpIE6LlCvhB9JqBpIs
sHycQL0OpP11mK05xQ5OveZ+EmXD3C3VX6/6k5xwKI7D8Djff3M9CMWI3g/VGhsy
Eay+PvET/qmLYmsy0ygy7mb8zlTG5bXsjQBfDRIsHdKMKJANC1ForTWLsR8LAlud
zLk/YUQUbOaKjoq+9cQv9NuUrLYAMtQ1TG75c/e+AkK/ehy4dLTejJUx6POyknuJ
JSabqIc0eEMuKxZZ4CH6upjGYyAfa3Mm2R+arpMOYfBFX92ZvqmU+P4QjKBl5891
5t3mTAFrtIKGWVk2yF9jwQvlch81ToQ0a7NVrYr1oLOWo7nLu/4OZckh2N6qMOJO
ySr0P4TxLEmVItv22cL5c1lx0dNMgOhVmzPPBQ+VkB/2cT1Y0WwGIv//4hNqfG80
Sf1S34S1ogaUDURIMCLxOf7aRkxfuDsfTzS0B2UfDE4Akpa26fZ6SnCQ7xW1Ab1z
kSLbpmRoAne64nOVPJVArl9PeZi2b4N9sXo8nz0KWreIFvWqPpkJSxInidNnbUc7
InZWS1aeQgar5qPeXHypKw4UzpFYU0Yit9j1HBFHoH8DOSTkOLcSjjwd18TtPNl1
YEGOBWvG0WxdYnvgKpUup99NxXZa5UlVAfdDTdNXsrVRsrqy/QxnDSBSFGuFjUyI
28xm42qbPR7n3LYKcnsZlwjWE9SLl+mM/EeOjwNg4TdlEoGVEcOqZIHKjCS6uSFD
QLc/HX4ggZjVct86X1Q9OEmiYceEjSqDa+hImt32wr412yWWj7JK1+cABKY8As81
/F8sl49yDrUWdrhT+jxPjaf0/xeDNSO07DX9RGSesYcz9ve3KqyJ9zt1t6Iohpan
mlebGiHXSU+7bnaW1wKRKP+K5/+ri5R58aAGNKU/Xdkd104LUehYtrY6yDu+iwdf
Gb5jEIraxAXTY+ucjWPL+GldPCzn4l3MkWxitj8bRPmLc51JS+lfhF3wWi6rLSHV
a/O6ESC2Ga3Ksie+SQH9rqjF9ByV0IZkhh01GIRixx+G57J6UIzMW0W8wBLsTTop
jVlMl+w1B5HxUyqsabKr+hzUSyJEzKDn6GbQQaZgRnkjIoG8lKSi+PwUikfLCYVv
jRTPvp0JEYrZcwt+PZfkwrV4hIIm+ifawb6A4WwdHb3gwU8gEeDyZJ4lBkK2hG+k
NaWpB3vUL0iB8xCxrJYBmgGuLf+zPrZECkoh1/TxyXBIjMJfoGsLPDQx5TJbIfcg
ewZqe0qOLWibB3iXDMxipqUtz08K6CDVNHfYRPXOZpk8HisekW+RjMxq9AwXmcOR
Wf0oAEm/Ivducag0tbeMJYN+VGQufjCQh04HI40Zby5wvPs71OGzMDgTvni3Woat
QPu2KBEr50foK2R7mkZRZGsxsSE337A2ikV/ktYlgVd2AtO2FUZJLWFMOPZ9jse7
LloptlxLSiCO45sDmecoS5PNtdyQXFDj6nrW7E3pKmlfE90o3VSsQ64EVFPcJ9bp
bG9Kg5nmU9x+KS4af1IAIlFu6ecYpvahb8iMnDfnwUi6bfOUA52CcGPGi78MX2CZ
WZoezW3OtzisMOZ85jkH0n/ez/dJxueTtFlHmpDExt6ePo5IfaFNSmolAdER7moO
iEs0gPae8GjwxpbrlVG9PSYzLeUoZFjUoTWfolRwY3SveZf1z3/HPuMjaF2xWZ/F
mHM2btQolT1kXvlVV9BqvqK/SZRo7r+9OobqvXIRpmnL+3Ig7rxdWU51/BQrwJRb
TQWBOd6ojjea9tZcowVfUdaDJKIzwTtFMZH3bKpfo1qc+8iTFtOv7NKDhbMIurgT
rVWw7y/xToxXaiZCg5FI+V/kBrdobAXlGnzquGGysFHeJqYMMZ1j/avmZasmVUq6
L3alFSd1AAn+0r9wYGebwem9cD53738klUbQNlAIA4dEWXgHV3uXYAfXsCC9NozT
6sQrRAPI6qifWy3JJVakn6diW4GgVRgn/EsIgJr86ioM7viye8LbErK24uOaGWPy
UL4v6D6imJX3oNVsPR1+Jc6+4XGvd/Hu2ZAYZpO1LuSMPNmlAIq5SeOAaE8IyQr3
nExGW5wTmHw+N5CfabeI+LdX/mBJB1WbFXTB6cDjfUGlg9xyPtVvtKX7uK9wmF0U
gkUSLNkVENwbELX2Y7y6jVQ8YbnEV1JUorMVkZm9y6fIeM+aWqD0MbNtYy+M7I4B
GhuKJ8pFfHPDy8GFojKwNWSPDpfbbZBHCMg8vGLQ0QV1ylH3flpg2fD47yoHk5Qv
yCqX+o/6sMRXrogE1uWUhtMf2gZ+NxpJGjOSYTBD4S6FoTfvUS2qflq6vhYrXZuy
JlLwCyoSL80OGfSvulOplA9TsV8QgV2+yf5T8a1GsdoIq38Fi4nyt3ZiRpDVhEw1
NERRJa3QJve/BpNWUHYX7/zTgIqJg0EZiIjJ11AWjGLbLpfyJey8L9qZ8X0QtgOO
fflYG1hQ2+8pDNONlnlp8+k3/ovxVIoHof84YqlVFsFwu6983tVeuuDFxkKa7+sw
d9xR9viPN4yadFTDrinlD+QugwVGnxDoslpub9mxWK3GH8GtZHpkebz+540WmxR7
JYfCve+hrqcDYPJsujAJVejuopcnTqbQW7FWR3MmX6U/0pOg+DDOYYbpDUNFS5ud
a6iXCQCcKi/5FH2irt91ePXSOxoM1O/wOBGyU0ttrhliDNDs1UPxrJzSvdqlrZ4j
v8q4FeH7OVoEZRp1M9nTBrAGdBgutPAm/jFy2hGntNvXrj+2CWCHOOJYXmnltAgw
nEBF7+usjcsdUobXUQVfDNGkMkecp2BfQtgPOzC7CXYBhC5QusLOA9+yRC8meBBO
aJB8E3V6/1lE6cdLPcn1JYSE/227lGQeuGn769SWPvzc9syWE4+KB8E9BLzOBgYZ
wI2JKmowu/7u4Vdxy51niiOk1IrW7CsV/V/XowAAEFV36A2vTLEvQgeJMq/Yu2M1
ydAfm6Pg7KVPQBVv5FjUq0XBM0r/DXduoVmDnbJhj8/8IYbszToNwQgW8SSPNUCp
TfIhItesgi9Iv6FcqbWfI0MHh1WbasvRgsSodMGUDeE4wZPmmIFCBmvFxCUbN/b+
dbda6zwrqzdDaF20CUGCkK06ogFGKM1qasKJMqD0WBU6c+sXzupYXSjbGwhVJIZk
wmioojZtt6cuKxFy3IBQlnd+NqcQpRQrKMu73sEwnn/NJTbDFxDZgE2TWNJ9Yr7A
7dGKQB/FGtgaaS//hJeyDCYczhFpVrKSjGjcOqTkUx/V1MHWMYGiUtmSFBQNHRV3
xQvA6pCGCnzRANRpRcZ5H+TEuzNwGg1nolpwQ+53QJApMdnbTOjTc/4bxkYVcoNj
hKYsmMN7oo3iYT7nm4Q/JRT9amubE9K1sUYx+zLj18rs6j6ZSMdQWsSgXqxfxy4E
bmt/i1D2J+51IEIzfQD21NZEKwG01sawJptjD511wH88O1DI+hWUaibAbaAUlFps
+53fJoRV7x+/ILME7v461rstwIfmGDo8hu5puzyYSBQuNh6JDAVExaRtyaxVySJq
QsAL9TG6dXX4g2skUfd87agsWj9dCbsXErdFxcN1A7DbhBbmGlUkdw1bvne9y+O0
i7dd+lLaGq7rOE9cediVs9UqcTvktFJFTVaGo2a6z9gm2pZVf6NX8Xxk16XNSqGE
5ufcRucEFB6bpmfTS+YYMz4UKVSuLFRsQOD1AVbJv8GKFiDoup7Zad10af1j9Juw
ZdZGQmbNfSUJ347vX5TlXZWk1Rn7oqvxGmnHodwbX3oghE9v5zz25vB3B+KUtQtR
3+FQzqxIoKzDubcgf+kiGOS1mcA1geAJsX1cqD+HxzCL7hI76yu6ZqZNpQqWKYYJ
dMwCGfhm/xnLqP0uaFy5zuPxs22mHU2EFa5McNanQDycr5uup2DJjsPtYzKBDNia
3Y8a7MEaeI3KM+aNHRBHXgNyJDtFdmsf2jRAdu6SJbz5Dc2GzvqpJj0Fbx65BWH0
YXpe9nWIJcNKUqbLUv9vHt27rXlSWRW8ctvOu5hv4cnd1CpzkHXpJsm7cMQjBl33
2eZFdTMGX/i+yTfKjE0/Q+dzFdDhSXNV8KU5KRMxO/lKrM1Qa1ksEiun/m2+Fq7Q
Jrv4yAQlVTqb22bdutsK/KAhIKYhQZNKFKgLdwoIUxqr1hb+b/1zmPHeF1oXKCl4
NaC9+kRT3XGIQT1ILuLLP8VDxvtGBHCynXXq7lzxYK6xWK8iDt39cLgVSFbFPWpA
mUlz1M0oR0kw8AYHqnMQXbzeVj6kJjCgcNxt6VV/eB8DMYhfwQtWDcCZAU3Dn7/d
XWy+FesXiEiZOlN4dsZ1ym2JeHKFi1Uu0sZoHNO0KAt6Wa7WJkT4wwnMLZ1yLRML
40WUUAyNOhtmpMMswzfiJ55kEwick4FbWZ2+a72LComlohvfFbOeaP/orqBpO1bu
gbluefPnbi+jB2lQHWkYEnFljQYsv/Ffa2rPI6P1RTkWzziijAeohih79Hw7/5gE
4Q/3wf7j9RCoWUdlHn6CUhiT8dC01iZEISfUPHzUiCq6h3rWKafkqBAWvd3UCJVh
QWjpYgUwBH78/94bCRatmsrP8cq1U7RcAYRbTZiCvqOkZMSOK5PETKomB9bynqYd
A78mYlGalY1eIEEOz5lxw4jJoYw+K24f0BRIEVlmWKBbh4iSBdPGf9SUzEUeJuib
vzp7jqDpxSxl0u9ZDzjxH2PzpccJqmjtkM+x1mVTXz4pmx3qXBnCteY/QxbBUwjl
7tlrWFOs61GCNSc0PQqwLn3qcPwjT+/eLdP4FgC0nW1GkeIFtyK9cJwDmZyn93MJ
XOx8dAmxJS82ONoUcwJxcnnZPWjkIvcbK+AGxdaWnBuI2oXFaUkn4yIQ9/l99RkP
GrSGgolTXgVUuotOAUmDE3sX0+fALXWPlH4AnP1XEy9UIh4xWi8jiuFzXGuofk13
M8WxkzN9T8vjgXx21F0NDTnxrqG9jtBTTF1xLuzdps4v9qhjC1zZZedSSwqzxXpv
DCTOSZ8ConTctfZUSD+3IpNpAngMRjhl5ICMuT+/8wSXspOdFtesfVJ5u/b9jo3h
u0k7a+9N+/zx6mPN55JCP30uetZbg9gDd9iktOu6AQrlrr4oINlTj/o1VVbYDwQH
t/IEEw4a/KgBgTwvb/r83gYpkOvvSR4zbQY/L9R14Y6p1airaT6pqNaGCDD+xYOH
Yj4dZDZJV2qGa5767Bat7bAGcI2Sd8I6lUJaH6VYmp6728Uv0NWOIwgr8aHnqRXB
vLryPGWV9drhnPI9NyaB6mLO5EHs7wzmSiT9B22hPhitb0r1BOEv+fX5LKfaahX/
g/lefdgTPg6EpBF6tmt9aU2kyqpfD3GqO27zhcCMM6VKb83cGI0uzhPsIp+m1OJz
AHjemjPkZclRbHAsQY1mI0vL+HmhvO03x8vwiicwQu5zek+cLHR7Zk1Psr7uGe/P
TT+L5+syLHRDl+fXomn/oZo7UrQ4/Jd1BwxSq3tkYdOez4HxBBGz1/rRx5atnyeC
aM9x5ByCbxOH68/b+fv10yUvUSBpmboM/N/oMVQOacYDqBDeV1wkIToEIO3tHYOy
aluES/AGpshgew7nuky6hFm6OiU/JTT0VxKfiVF2USstz/IUTYVOrgtO3jn0nSE/
8e4jn275KfcRUiCl19GZykv2zesLj7rq+i6eYIbSjNcjEQYAVJ6eN3d63ay3w9KD
JzaCuvpLhol7Jun46niRqfjMo4VD/832c5j4yj8XlO0HB7kfla8uybbk4eubENNF
h74YGUjoiacHQZzN0HTZbWXFULkHTAml4HuaCGZSxcgC5ys+wotYJGRYejGj20iu
20rPpEAEnHcYuSaCgxlDVLOEFfuPjDzazNpp+v5o+s8Xg8yvk3Ix5aMor1mjc1pR
9tcg0Nt3uJSTCL5sm9CAVa6dy5NoFgvVKJg/4md7nLLjqLYEYuryVv7xTasxVf1h
Qk3dE7L2sdceNtItRAdL4gDbk8nuXn3+lket757Hu93GQ2TUyryCTwYTTMO1q8NE
s/zLztE48uJQPP9l24YCa+sNCY1cfhIeA3InR1nyMEqdzTZT7cI5AnfOMJ0gcwn1
BAmL7WnCUTUSFhBKvzoRCKtxqCUO8aLaLk8ABEmfXoI02qAhJsLqLaPiln6B5jdf
Z5mYlGJc55Tr89mkJzFC4EYGULDPwWHgzBgZ943TE2AFJklf1IW18+WCZXKkGgEd
HRFGHQ6/0M1na4RGp8TEj7D/DC0fuAy9F596oF3Mr0wQigrzzXp8bZ2bNHTGboX9
FjRz09jIDgq0PI+uaRmwWkhZTyZKyLy9MmpWkk4vUC9LMs2g+aLPx67VPpFc0hDu
u8TFuQ3d1cKKsXSdlG45NcjHVmDCPt6ZHTIssWNovw6HVoXO8MlE5dIsbiFQ3lKz
fpzM3oGQs2gu7sFnIArzAoaxn0DTMMMeDyjaDlkCLbTDy69hh5A7qUNOSHXuD98X
h2R2sbBFci0BJz1Bw38VizlUtL8F4VlGbkT7xYEXOJDjHVgx8oM0xdSo5UC304Hp
PIHspKDkWSfkguGxJmF4MVeuIIUQVL8Dyatg7Iqv+anp6LS7dIZjaOcgaedZTmHS
QlmYFcs0M72IHGEvRWyuv6gxGSsfLnLMolGmB2u7jHs+6234QWhjzAG8EJbqs//d
e8C2HAHEF2JoSxkCuFUaNzjp+vWCloSjFGOk1Fi8rEWmQLtoa237QuSYwuoQqZ+0
fqPYMBiJ+xHCBc8tCjWKcxnWaV8mwGmO4vV8dlH1ZFF/Wcely4hzjg/9Kpf2+WmQ
tOaSZN6mIQ6ksjcLQgoJRdO8JuiHxMMg2G8xpuIl0Vu5Z39aiznOrrZYWAIeOu7L
uOKc1PIVbHnQQ9ir0Or5I1sFhBsR7kAyARphQ/3Qtx5Vr+jj+i3BOeswHzSq6ZPH
arRg1Y0UzywKM7EwoHD2qGJRmkOl6Bb1mSj9SNz7YtTv9g7jfeExHtSFrUQDOK09
MNVTJiCQfGgX2ns09XKhRKI48GmjI2dd/EWqRQvo5msiGfpRGq22cYD+JajLWNRA
T3HhmlbTHJf944nFXsP7iD5QVnVx1wgt8d59CPchhKoLEc06XZ39slj4mmvc4lgA
HvGw6VBW487N9oingSDb4ZaLPMY4bN/6Il9vwfxja0dM8Un8PUuhQC0AZfFqS6ju
NolQ1dkBOJ3R2vd6XzExACNXkWPDvv8ohpD6YcAAkiwEqN67ZDWkPcW+kE2A92kj
mLxm4UZ8rKeNasbn4VEWhdaRzyLXfuHth6cIK2spw6VoQ03/4DxYE5hsKgPcHpHr
smD0Ib+ws1NngNob1nz8Hz3kOMvY/iKAHsidTXzrJ6RsiMZvKS5Vf7lQIf8u72mW
VV8Kz1BierVY4G0lEbqZiBIdNnqQeVnnaPE0UajbF6TRr1ycqgk2jSPY7snosn/k
d3Rv8K7jFvICjATC4prOm2nPyAy+ez59Ys0W6MPeuzb8DQYWPPSK9YebIAuyRW1w
YxvC14kuM7H6a/njlX/2FOH/YoHf/JdMtSLBq01uRmIe37kVzdJWwh+0RmPP2iU4
0WBRsTB4H7fHrvk4J5FhUkyod3GgdQszF23d5Fu5Q2R9HQ7VS0aep2bkFlTnSufG
fFrFqFSPHP+Cow9symoeOkZG60InfMCFRFDtQsvrtmnkvqEj/EkbhDNCW/Sjc5Ou
XW5TBF1f6EnIPY78P9hJ+cELpjTHtdsfVuG3T0v/c1TlqflU3HcsxbTfR8R3p10X
V+Izbcwnfpw4q30vCAh8MuvQVERu9jYeB8hItHd/DkJKLRAkW0rKEFWwojQRaJZF
AtrbYsAya/f/3kCFVJAHxVzWpcsZ006Kar3FQdvj3MzkeNuNF5zdVdqBSVT0Scjl
9e9t/pQwfaCe1ff5eR13RyBtoRvJIQpHu3Q+5Pa0Wl6SnVRMgMjh1iTlEx+EZxtn
GoBOmle3Lur3XVT88gSG6GhM+qFYwoteIeWYIQR/1UmmFgKMwavYrFclKK1DAzHd
xH4nhw7+MANrm7w69kJ+r3RA4nKG59gcpdqcFFbbNVEpLoNJDqI2d6EnpP3+WwwH
MV8S69mFYXJUASBcR+Ec2qAA/M3tapToLN2Gj3W+7UtZgW8Koq40JV9gKytUxeuF
FKGKbpW2xF1C+yv6qhcHd2XLoEjuEbxaDmezV7xSWXx+aEevOPBOSHZNhYMKnrfq
eA71oWaY53PpY2k5LWzHnzgdOMz1wOF87xF5pQA6Qkpj4EjAO5TyUreiALCksfpL
mYs0ehVHMekKnEyYOtwaiL/LkTPyWKZRyRGkKYJc/u6Q2zU5impNnYZrMa++0Pj0
+uvxsLfnNerBxsIKxw2/OtPJKNfyIq6MflEDwXSxm1/kYeZC4s8Ay5Yw/q4Z96Pf
g/X5QnSeqH3UCOMsXNweNv4Edbi/JVVBUSov3NuBhshw/iKc9d4kNZMm1wWBy34t
czweT10P1Sax1eXuOSFwV68R138bAMCEFwQbfNasiOyYu9r59b/3wM1UGqjFXR+e
Cql7kT1ib7/wHNLq5XCw0u67jJczS1YzQ6zBLVCVh2j4h+PbiBM6fzfkrPlT9lYu
eU8xPgejmwAvqoniejzN7ORQ9XyA7B5cNb4iAk2aUzEJeolHXuAa2X3GhDdpXbha
ST1vlmWWJ67kfrPcVh3sxvinmuMErNQwk+msiwFWPjiG2TzetEX67qA8ayPS/P2K
USIATvl0pwlJ1sgyb7Bm94C3IjbG1M3hUwe3k7SOFOXLZQdrlGLMQmNl6nFRzFeC
8q0jJVaP0x3GwAnnPNXjK7vNZxO2t0fkCn8wytQhfCvNGCuFntxAAKnV1NT7Xuyi
HZ9t/178yEO6wD4OeweDo4LvohIrmp8kZueJ+NhOnokO2tyl8s7CVqYCHgbfqXja
LCKBBTu9XqWlQ+m9ulL8WUUP96bGk+7vFCO/OAN0EYBbZaSuB4e741CDkGxtUgPu
pIN9l+Bh1zWHgehGlPkbH02PXJqp95fLx5pg7aW1fJ36lnXr9YpfBZpQTr+dk31C
phsPhPbVjQE63VUWDfvoysZRDvDu98Tt6+O0ZeKVCmUOjC4eUDIdrmRfjhbhrWlx
JYTuZJnw3xNAGLgqdYMva5Joscy1lstStbxZdSJLkf6zB5ibXl6mH2zHWKJWiOVA
tS8ENDLSXTtwBS5SXCAgfiOvKxhw1qZG81qX/I2wKgDFN0CF+aSZt3cykFkQBbQu
b7FBgD7SWHXtlkEGH2m6v4ZBhY6vRP7ds1Otuq19zzsLpAy6ovE4BsNtXtgPGBNl
dhToEVKk/LYcSY9DsEJtYjyE874x91WnsHSvbwWafYJl9Tj66ZAA/iitdXeP7mBF
PjYwxP4hcPDLXlU7q8XrKyi4yBnYVh6g7b2X3ip31BFdy0EMn5MhO59XkRHsBOMb
JX4AuHpfUbuTpBbqFpj/FldGt+ZAxH8ZBJ430BrNyqdIZnn+ziX1ELjdJNKMQmYb
E760GRlGTx8Llkp4JLEuuEONcXurCn7yGcQ959QHprhZgjYFSlUufdN1sNu2FE00
JGyKoxxfttt3fg/yuT4TVNascLS/fKRmDKh8TYkJRoIR5XVTksKjEGdSZQgIGBpV
GpXFM1h/DMaW7jRn2ppbh3wVtBELuv5N3txOdzEiAcjiPoM0Rn2D/ZOQcTSoSxDF
AnQn/B3Kh2IsYrEssASK2Hz/QHY5G8Pe1fsPO1jN3pN4gcejl24yJgUJvS1NLmrr
Yub1DAEz9Evumz4Fz/WXouFLQ3sHEcKnG6ax0IglFoRp6gUvL+shEKmvZXAah2Cz
TKBfo4pNs3/jO7RyIqF5jaRSd7bpBG2cDN8O2Q6n80ipYbC573OYKxXrzAA2nrEu
L/nedF0T8iIKwp9JpN27qTqEqUKSrA2BYeW9SUiswSS6AkCYUSUFlDJOgorUqR+A
BTqpoSodeXHYeAkloXue9PHzAwZ+gSe2ZnjFichCx3VkMHs0rwb4GLHP6IiyR+36
yzXhDvv5hjV5JUFLtyqhCbKrPG0+Pv/rivhpv8xwfJqbhu2mbB9gTw4mi07OZtl0
6xeODCUG6l3RXH1vsrGVqPuVoeVFlhQ+hLSb1rStKD2xV80ivPp7yAXlgTUXhJZC
DnBB6CtkNcKIXJm0UdSwGOHQRJuqcWQc5BPE3Jf1LAZbUF2OcT0IUWHL+7jif/L5
a8Izfz6DxnrzIwpZkYLVST64bCUnyXar5jAEf4OlIirENZm7GHMe5XaxNoTGsysi
taVwVOdhvnob2v/6/ye1XCDB6ea1mKh66+VS2Uku8rR6N/0YhY3XGEdGW7IPAQCA
3TD7SbNjCEWE4ymvWrOR5CtBNFS0bYPWtJ3DtYyzXTT6nxnm1yHoGdgiODTHN8tM
ysRz7UpVB7u3DJy0xjYWqkzvZx+Fa6kcBmTmSJ5ET8OTwTCJI4X9glJ7ZoCYZM/l
xzXdrRQ8dMQpaffydZOky9A2JH/FjtbNVbetHt3yfg8nG8pr1Gtvd/v7J3Zw2Fur
keDiOG48F87UEk2ZXapr32ijo0KWvf5Dp53VzKYdqxiDVnIPEaK7fszUicXSSIox
OsNymK3sLDFGnsnJ2o28rS5Johzej67ISBnrnD5H7eqBWDWdOZn1pNcupXnULNu8
b8yDxCvigU4KC1faK2Gil/7Uz+S00cxpGTZ+w8zP7BxvHsICpWH9cBCyWdeWixQu
jLx3BeeJ9jCUQp7+LM9QV5HSRuq0GB9NHKYYhKMd0shDXZm3dQ6hP8WxbCqzdbbk
s5lpPdSeQB3jycBGMqPSNdmxB2osDaDrHhBrTY8RLsfvjFfOov2ZJ2lLFgXe8jIY
39DlCktOgoH7EyB2XplcNzHRB6JAh90VeurPire9n6gHfi9dUaIQiBkaEuAm9ThV
k6dDecF3+Z2H7TUSDq7s58dJR28T2xr4EOFLMrVV4Zd6gFhNIfMhcb6DSNYM/yvH
wIrqrsMpKf89n1rAfhFTFaCf/w9g/po7hIcNBIVbeFY54jxDT1UquI5QhZU1F5g0
Q90Va6//G6zlRdQ2T2x8mYkGOYWxH9ACuPsI2NtYylkOkjYx62NA28PRD9D7de9p
e0Xji4qZnO+SEAqYi6OwMqToSu9XwYpGhGFFfTzI6FwFy5iclyK6hXNW+JpUaz/n
NZEg++QdYozXBIZ9bMepKFi3jx2tJbfx7OTbBA1R/gvQIZ6N4e7QnK88aFC277zd
RZ0t9MXabiNF+SMiJpH6ZMj8/F+l64B5UE2kjd0FOIEiOCWgEd01+9xVFI0xCdGz
QZW/m+Kd+MJ9IJLmupvzX5GJQ/Pj7mUjk/JtpVtejRA4feCSME9wRsDsedexA2ve
btInBmQFbpYcnrET1T0hAagmaVKeNSwRXrFligc+WQb+YMFmbEOfH0h8K7m6k0fs
rerPP+wGooxa6gPaBtO/bKWp67qthk3qQW12KNYa6NIN1HKaPuyVAtUlwciPSOtn
Cj2WdVLiMH+mTVAFKXrZEp6urSLPowlZ1gKur25egsaDwK8gl0bqeOS+H7j8+ZGT
PIGhcwfONfZGYQjmOeZUfPzPTgzARpvtoxqJejQ5CEZ+D50TF+/YVSDtraz+4MQN
Wkt+xNBEPERJzddkgOkEujLJPhWh+50hhuwrbmIMhmVCe5UA7Ktq2mZztq8vsbDV
QOZHE9fiCfzbw8F+DF8rPeT7Udht/hnmk86tRM2huNkXbssPeGjkQd3hV1v1TDfa
6kuABozFfDKVpYnE6hCXzRG64tP1nt/y1bgq1mtSNTKnN02/J+T34LnClHb9NQdO
UWmuCVVJmcQ6ypiEJQrk2Neof4qtAy5S44TJU3YkV5jRyHezmpgXzEF911BMJYzx
vvoVH/yMV62B9vJEoaahqZg5tfkE7P1qb4/HKODdv//ys/Dp9H33xIyw84zPxuBK
4mv2FXFNsZrnV7Zp6JKsYWX7K18z8Pd9qqVBNPBY9Urir3X+gREDYdt8M5JFoil3
curQnyko1Yon6U/8PXyiQAUgt1voPQ3d5pk1dwlzNtTHyFATjyPYdOL9mr6DpTBz
HG3yJMR6s54r9EnM8HaJbuGywgymVwBCMb6luqJ5SBVZW/+ScWlNtteSsqj2C6Lg
dBvc/w5i0PWbWPqKK+RdpIffG1n54U+LUVUEqkWcAov5/ENeBA9lX7XE91RtGiU1
6yZq1ytC5S62cxiXBF2xv57L1ooeAl7BtKDgmzOZy0UONpAt0gg0ZoKELSK5q1jT
4tY5tXDNyyorXB5k/rdyzg6SxvFKP+moznXyPVeIHvXYxmJfT1X0IHvQhbMwxZkx
cNeLtCLJY228EGi58Wji/wwoA+QRW0RfLvzfW2vebeQlG9hl4G0m0H1GhRz8GL2e
6o1lU8nfL8Jmry3r/z3qMiTMXDPUoZi/ri2Tje8Xi0e/tu+pcchO0I/YoeKx6X/5
wk1muDW9/KVWEvqwSjy4orscO2hNAXchSLl7L+3mIM4MqMzT/ZQm+mt38oeq2lru
8hYlNyDfc6anIFkbhPNNURgqzkm98mCerlh5zHZPgAPIVqrq4syZjZvrE8IS9iBa
QuoKsOF40ZsXZdClLkDrElXGQ2HAmYvu5UzbfcxSxxzVfZysg/UDJMpkLYp/wg0v
8q7GPxfuS3pNcl6rLgt0c2R2vIR6H4qxFGZJZEX9eIOciHDmOpSFoOplcreRHiKn
sTnj2oxhEL2eK5cNPx2n23eYWTAK99c2AYLMHqIT8yjpQlydHb1znW8MI2SwWPgd
2E+/4on896pryBq0eN2ofwWfLays7bydXDD9k6Fhpu/FiTw9d8Kw0m+m5ZU+HMPD
FW7/1ZCZPTrRspkraR5mtM7KoWnkNueCZ5BO4G3y6j4N+cYZgTTP6hEgDo/ExWHb
NOu8xBliGJJ1J2HknlhqpLEC46p2a0rvpnOqb49UjK4wWFX/N7P7AuNCygcjT0Sp
VW6J7mfRIskU0g9xPFKLVx7fv7cuxSf2NjK21hcVHdkLqzA3oeRYHtXsaE/iOIlZ
nfCY3pI2BJraZiAjB+Og06nsvV5m6LkmUPTTmBdjJyKLu8iMRlZ6mCB29eWdgQwI
VOvWfA8q5kJVHrLq7K5Nv8pZHMhJ2STvnqN7EhIrRZoICIb4lyBu95kkNh5N/Uzj
e5FR7iYjIYJ6VVonyqAzqTAHX3jOowep5YnFGEEzRs6IkvtUfSPTa8wHsp0/zY7t
FvTQjAv8wGASEuPNtqdAbqfpsYkvOhq3pwDkCF8j0kjRGTel/74q7YbUZmn9ULA6
lB2uUsyNp0WZDhRjm/WdUbYG7172+gMPNgUvkj5rI92FZyp6qf5njMbh97CGI2/D
xZWLmgQDOCpj27YGa2QvkE1cOsrD0FoiDWxpo+CcFAvT9RIIcWOkBPsC1W29gJhN
pmlVcRG6KX/g3yJ6VX0RKn34lJ80A871ki3EQ1g+k9suByHMCVPWOte/f4STo9TO
M7S2iig5h5ZPrry9zIU7hpPeJIu51r4MB06TBi+kGP7hD+222JUgK5qbAk7kLEVY
6dQhLzd/bI261bZMwhNCI5cZulPDhFNXqc5Oh2iFFIggvfx72y//sHdn5UmHaMZm
iCdaWKsujs2ANBOsY0Jq+ie75K3gJfsGEE7RU1dV3sLP+flLQsa41TKLcMWTiUxh
t9+5X21lsZr3KnN4dDvrLQxCp38VOBZHhykYA4BfGOe5px/ItQmqGwvQwCHBR6G6
iJocRY8C4spEbSmfihXMNJZFJT2efA/Po/lC6yMqQg+pftdktb7eGs44C/kDySLy
QC//wBOsIub0bDaKetiClUQujDociuMPmmvW91H09C3A200wl11dG24W9v+Ta/xU
PPlE9rQN/boWXva4vVWjHgqcAhRNGMlZLUtK6d8KxrR8oN8CSGj+zNFvl4JKDehg
ZPOwUH1urHksIySqrEZEhrHcYJj1WFOXXiEcpzM9mczVieGoqbSfFbr5cysbnumG
nmBTR6Kgi9umE0+zkeGrQxqf3gJ7V2/Qmv2+yxqi8xQAGlMCd7v4xYBxorOtQ4Ov
AB9JGBhjpEKNrXG26XOhg1HLZsGXOalLS2+06csEsQrkEHdiUWzv4wxbtoNbC8zh
IRC03DK7ZEo18BuUPrLMLIwyQYh+DPj2HCV+ab38+D/Y8nmuTGgnYfgia8qd1jA0
JfYAkLWNa1/kK5Dll7H1J3RB9o51mlLECW/6RMmLUblr2tWv00LGcqu0MPE9Dr8J
5eih/uaGT1Dt87Iooz38zz71gEf+BXnDAmllHb++NIIctKwDg34Fpf5ECxr7QJPd
SQqWisNRVP7btm6ZJZOzvcaVDyRKRv0DUaGkCHimL4Ok25YYWqS08ppTRn+W6Ov0
NnZ1aJ9+8EV1Nipb0BjSGnt9CBKGkqTWTvkgGNBZQam5zkEpvDK2k9D+JsOWEDYn
c1fmDOFREfonf0FXHQtLTL+J53dVjsa2kGnDUMmrZcUxOHPZ1mBS/PuMCMQyN4df
JgirJtC9+f0amnBl2n85g+nXmI1R7czxTE/cqCFIzgn/j8HnRZrhKRX0wXjR+FXf
4XYkj/hv2b2X22+CzZIJr9xeyYKVLqpteKiH8klk4Fp/sSbbZBbZ8XOGKw/OnhuY
xQI7GVaVm4mqNh4rK4nQSWVIS8uXuBlp9WOk2cirJxAqKMjQtBqBQiQR6KA1KijZ
Ulgb4aYse2H4gGoO9SWl2MklBEAU4EJOmuzUN9FvkCxrwyfgKVsTcUJaGL+Y5+mE
JDP1jcQ57pDPs4N4a/txxGkpZGgVS7JOq31c0QDtGtS6+YzeVZAkfr/0TcXfu5QD
uOV7ygR6lrzp/x3E8idbWuvRMKUBiy0b8M5LR2STcvvpYqQUBaQsxZRNE01USYXu
+C9ixP17jvcPT0Yyr97y65M8w4CDuDK4uE+WWVUK4Kp796B60wOLYx4YD44liC7G
d4h5FfC8WKo3pEg6Ud7XLIsJMv8BMBuZStIV0tsnveTHFYxbSytgh0O6XSzQEG0A
RU56WF7I5FyHhrWSoaHo9v/3cO6JxAu1nQkEuLRJnfEF7EnqzWG3B+tgaFUWAj/g
DY9WnHQv5HzubPNtu2j446NUGvaifAN0WMEhr4Rm0wFk5HCJgRc/ztYyIrBXgtxr
pMc6b1udDKb9Ew3xQvOSma9G14tcQ+BMXJ3/bOOYCNx9UDL6Or56X0EeoukUrcWv
hxAlO2yQRelteb1AKKuN/tFfJZCkoMG9Rud8ywDzko4bjNp7amCnQdCU1CU5hnY0
Snzw3iapgC60HCoKRe2snaCQjyxHxA5yWZ7AdJz1AJ8WeLfMzhhb1OWYkB6lcqYw
D/0yGbU01yk3jWdJ8WtOBwHYFVGafdhly0R2Q3oetvHX1itfFe22WQqVxmggQ7BO
dOSSLtSHg6NEVEnxLu4+nz4U/bzNkTdTKBjePV3Z/C4dlUNPzVXG+D2RlvJSGUcM
K1xlaujWYzy5AZNUMkdIqlitD4DRU2zSNt9gkS5z3V2yIZhVyLX6KFilX5I5btWE
TvDpaxkPrEzZg8sqpMe/NfUfHvqUtc5fEcvCTIONMS1jgZyclvwQ1BKzviHHh3XD
NAoUYwFln/+BSe37kkIFwhskaNb6WfDLVFtiseAQsRg1G44j3WC2bkQddN+CQc2f
j3tLvMx+VgNADpbSzglDnmwbJT5jN8aqjBqhjWzG/7tZs2kryXlI8cm8EGMcwe4g
DwpOdw4uQLXgT+9QYcX156yttW2HHbHukUPTnSo22pyDdOKhbvT021n8t14s3fwJ
N4kxO2veTBfCOviJfisVQaciUDgmnYcFPs0N0I/5Nq8n8TAmUFDvbdHPNvgjCCJr
cmM747OMXUDGRdz8jbTg4mTN7C+QpvRNLAX1awSSycbQ1KCPQ1cS3wTArs2LFJzV
cXzwJErbHQZTbpU1JDx0U7auOcdrlOq9XUfEHYFo0S4ZTqw/jwgXDiNJqw4lveEO
v3sMwO3N5BmKh+2cY6GFN9ub6hfz6ouOASV12K1t5mlFIitJ0i6V0Zw0utVO6gxu
dOTZHCHWIHkotia48UPIEeyBRRHPwgc6Ou9Ah57/7qAiFhdyM9mt0wMq/9ItJYck
iKbGuexX9OMi8IxOjj9l8RwItn04pbIj8doJNdMk+g0CWotGmEaP41dgDVqrjwVC
qzPrnEkwJyX/JYLQowRnjmKRj+j3EEYYc41F1IUV16AohB+0+7dTglMUS9zkWx4q
c1+HbUMwvydb6+TtiqeMlxSXD9YHh4PdragZ9GX7Ln9qmwO3VAPNN3ZvO/6L7H1i
c+phjJyLaUnGIzQ7despW4ZXFcXgS83Qwp0Zr2ds+T9o8851ZJnAH6nGNjw3OMNl
u1N4Ak4BxnV/xAazUMS33L0CyPnKxtrWA5NPTrCiYWy4AlfNnayIdU+hiHRx9RuB
PzGPBDtEDx6B8kStkujbuD+Qzy8kwQ0tAskWxi2LHuKjoO0E+vNJKnoIuytyZTQZ
QGnuWxL6TR5KhJgbpRY5tMx8vDcR6daRPWskxYbMcxzsgDjR2WrW3ZSxSkapPwVC
cQCVuhZTH6mJD3xMXXzJwpwQeKCxaHy5l7NWh0/8NwEMKynXla+Ts+jIooB4He30
EL1Ihner+H6S8m1NSNNSbjsajcZXrgVq23MiPLv5luzUEDyMicKWzOdxIoJ2/FDo
fAUS9hK0a2ZfVtAp5B4wlHWO0r26i3XRsPaEEzraulqaEsWhf4DWWF+A29kDjA/N
8jRIw4jehSbhZLv+Ew47YKm3DGJAaW2O7c1TO5qPlvgrFehikZudqpwn7RqXXSkD
qRZMlWVkHwhAybM/hRTpoi6YpElgCLKjuZW6+RhmrfQcxcsopWFYMMaCSqr0+OJy
Hn3StE26DXtyzUM2UebNrPq3J6z6NFOO68NELnyA9T/pIgo9CnxnPKHp5IXejvpI
8qjUAPfxiHKeCSbsxFI9P1jTIF2QuLKHZSZ7yDMv+wA+kSDforpvY9rEk9FVJgkM
fKRlJglD++U3XIOhPPnufshGILsgpVgdcd10VEwFEGcTfOMQhZPIg9CANPvdVAyL
rxyhEIs+g7HP8x31NGCYal95bq0pkIW5hOR+vkTiB5Laeeus6uSiYvKpCR2mTnWp
Wlcq0LQENQngTbYGuJL+t5FFFgoKNQS66P4IeCNNoI3w+icG/euHeVjaLprlLQgy
4wg5P3cveW1Wssg6RLSlcU7nKjHNNyKFevqyru8QhlD2gRyhtu69bmZgeMlHudFn
2EyHnUGZL+F9EkWRJZl7sXLCnQJeYDP9HCcRbqZYSf/xkJV+qtKjfKtr7CgZQNR3
xgcJS0Ge9Lpwr9BXncUuFtQp3VXL/BQgXE/XFUevJApXf4szX5mD8oCZE/pgUxGi
liETQ7z6WFo4x2R5P3AetnNRfnVSSb6pmsY5ZkK5wFdqVJTSlxKfS3g7comuGZMz
gWECM6Nyj9ULJ2/g4ZD9pJeRHq/7rMp9JwmbDwq9/BBLNmJPnbW1r4yZn7XMQrrd
KbO7UJTbTSWmCvHLhQcS9AvEVe8l6jdsFMUeqk4DFEi8BosicV2WAXESBJm29t+o
aJfSqnxUVD6/B8aWihqKTQYTheMrpy/eKlF2yB4f5eBpnSTPM8H3W9ztXEfAwtRv
lRpVmSSTUjlWJUtHdA1G8umJB6S/Jdu60oP+WBtsgnaUUzNkPQGRECgM6ZHCSZEn
87Ys5QLRCJdn7ULziSEPXSkkzfLGOM7mlhPWzZctY9pPT3vZZl0Q7wgUqpZY3/iM
7xB6JOn4GEBN5YDyGTPIQcuXBS6eOtDh4iJGE2h8c2jKD/ucQ48y8SjnBcwL10vZ
fDfLWk5XJn7Cr52wIRrl4aulzneG39BVUthHXM81cE8gW3tIEVOBaWYHuWoZdUGM
vvotYetkADqO7kAWsQ5PNhQ8l8dbuWxtN+7MUTzYZYRs1OiNgzUglJF8hjocZGci
FxmQCfpHeRVk0WvPxHNi0i+r+XzUx8sBs3LjYvfP3qjnbX4xN3jmk9q2FBfZ+HyL
SrLem546+o8hYfhPyRrPFnHdmPfeC8j8dGVAIFCZO7PXF3vVfCHPZPPmm3sXx6Gu
WERqI/Spm2/fUs3tJHYEPG5zbnzO9M0yfpOBbR6fceY3wWabQ3HRd79GBwr345XT
TI5bnJECxmND9epdwxtV81aM/2lF4NDqSBSCWbd+joPAlpgby3L/mIxNONXWL97b
48mCtCi1ea6IOrR37RnoFoBeh0C2jtFzm+9GOJYH9MmOz/041/0vUYKyvIvOFtsN
1/5pwrzEZuatzQ+YhB8hZssitF/9LYkJQNy1SjzTfoCZhDKGUKZGaV+oX2J43gET
BTI2te8unhliNGJp3QEGZJ77msnwjiPAY5GWzjo9RH9XH+R9QP2RfBJpESUF/7qj
9ZWWTLiJuoYuYEWF2TEi+R92Yl683qYuiEMkQXFpL0MhasJkHBBkUHJ89PakwuHM
8aL2BTpn0WsUjWCktdiwYCjrXJn1aqe8ykqI0OejsXaMkLWSC1M875H0ydreHHiB
+790V1ucIT3QHtY4tELMLVGRqxuv0/q2wQA6InectG9x3BQEUkhBQRaQKtWzF0fZ
VccsTti1zr3pcZv+cg1bMiUwptXXoH8Ogjapiijxtfl/IcH2I9ZfOYIqrbNIR+He
xlcqQe3V8q3IUhgRz/KDTpEBvTdmTWo8uVYkwgoQx9EAYcarylk9pPO4qqDcIqXs
Z21uxdEOipFPGQFeLZKwYhzX2AdFQI3A89tQVeARfczChQ64CaAvWMTL9TiP0UPJ
FAYY32d4HjMaub6tUsY00d+tTVBiblQSq1/pPQCyEqf8lENFuaoPAAGnzBcHT9Uc
B/uTULyilRsbksSg+hFry3OuUedkN34J4987hih7rD2QcvP6JsD+4WJbtIHi2CDU
rgB9wsV7CVuKv1Koh779cjN8gHfq9lt/an3ZKfRzz91iIjpOPTW9+wU8KgASxGJd
xp5u2oYD9a7XkzoObTGoJ71JAc/NFsdFPw56yJkMNupjVj5EQlLupqLT6VuO4hLa
ql6URDa2FN6UXQBrgXH0v2Vn/0uPgL4ZXqtEynrrJNMdE85QqRs8kgCjthtYviWO
rS7W3tLvA7rG00YFv07pQvkp21UvXHuJxp9yhuSZdc0s+PtJoiFZpeGrWwAt9ogh
q9UpBYbdXAnpIL33bV49wrMd1NpqRIqIyIvUyymvRsrBIvPKFL/rYRlDCMQHs83/
zTrIKrNQLMGA24J9tI2NUtK+Ous2DPIIEytk9eAc7K+Uh7CJDk6uuw6uywaiFQqE
SvIN5k2Co3nF092yH8htyjs3Ib3SPlx6s6a8ASfD26GL3ngtTVq9fa/GFepxQll5
gQnxxeKOER8h/MhaiHhsWxyIK/RzVqlqwmaEQEyQvAGMoYVpcg4F8U6TxeDWsZUo
dDZOEO9dyvZjEiQW3deXdCLjj9y9Ae7/hd2vLn/eOmge/X5Oz1SN7OsoX8Bl0259
hllqYcBx3zMVMvVeOx3WBYThEnqf506NsYc4hCgiUvefw8U534eoO/RBcfldkbV3
pZI/FzpGofwYsuEjfVH41UiU0M3ApydQp7TSQqHX7gojptwkbP7ZE8PCr3je5604
ShUwlUUE4kOnlkI+K9py1saIBxZvgHriH6RUgnSHMim6kPsu/zpk0Po2SdPtiB8Z
tiQPj4eCFPJ24kyU90Mjk81yEZjgw5fJRVtlvpnk6NbbxYDOSMNEAiEOwHWQTa8h
LNxqmbsWHZW2sJ5U5zj1LwCXrRUz1WOGxctHLdTbMI6D8oud6zrR21/Up9t0BqAq
bzSaIfQ+LkGCYNnWQgSCegJuzkcK+gtZbcBvNqJ5EwvY0NFFA3mDUrxkvFtSeblz
iCbM+21cb0VLO4JrQ9OeUBA7OBpYmUtDV9BYV0aSZcJk+NwE9QjbGt0JxlQaaQLk
jsAoVy1PQOhn07FmJuMj2KsJRE4ZpvanJMEm0HABMjY+LS2wkpSPzRyfSGRK/WkK
hpPjxmSZKb2Pu5nhS4suewaeZmRrCvT6IfIW4x3jJgVvN+6x37jZeZ0NRLD3BzO8
Gpc+qbGhDAk1Dn4z2WUlusWT9UElR3Z6Q1qsfijVjrqbUEWeyGB6ZkId2qFn6/Zw
qtFknW0qJ6dsEhQ04tn2WbPt/7GZixYtV543FQfcZL8letWKWK+FDW4Lwb5zl1aw
Vf5ypOUrDHs/ZIMjEEhY5zc9+9HdTNS9LmA4CNv33J9qUZw2kLw4tZH3iEOUZJ1v
zzPRDk4vdwRtfBRpMxp9HDzBVaOJNr6YUOgFP3bEx0mgldY34m9yWLputbmULqA+
QUIHUWQNa78UUDQtx+5t3G61ih7YpoFwWU2f6q2kyXG+0xwedqt8UBh3dbzXcZzX
YJeMBwMTjQTae7WLajoZtOtzMX0zSwreFSVmK/RZUxceOx/9Bj2lTmGJhrlsNyW+
YddtM8kUJVXtJVnLUWnP+t7kVOVVyORZfL8FoYX+sqvsB4IdNSglh6zpJ3exS3ZV
llmhYh6YltQflW7Psl/drvdN1M5OdtP08dedmCsTffsQKWChOMIUV2/f6w/7pG4O
zfpMRf8pE/iD1jZEzK365pkmBJB5yK+wNQUL4UoaWqSHKtKhLQLQvy7zE2mU3DuX
s2uOxgHA/1C53lPa2MvjdWR5GRtPST6+UuYVpJeK4hAXQF4IuUAMkNGFEiGiTpjk
QQqGBmJO9iuZfLVDFa0gDU759f8dojQJd7XD3uM6CV72XsIN6xoDknE4geh0sO3l
9Qn2CqNaapS43kE8JzcK3O/pIDA6HJhSs8xJOHcZ5sw6KRGCp1f7wZhUIdRaMi4X
BRXJFgKYR6l5su0QpIOpXbYuCao08KtwZFPO9ZXWI9gDmRmMeB8ufevLTp26S7sS
hfKDUuX7GeZY5n+bhFmq5xoQfGiEyOXNYEqqmXiPllUvLDyfw6fVmIXz3OMyttG4
qXOITKiqat2QleKpPA4MbXkkAFDeGBDSybeZsh8pvPzWOLLQgqSpI5NfZ15PaHbu
x2EviG1Ka02uNxxSI7fKzIziQGqpgV8n2hkTxDUSmuJPMKjT1rLehruQFlHxGmXd
WDQMtfZK77/S2aKZv12RpK9zSz33fOcPRPU3MylDbYv+n7mjeTUSdJ3RdWqzGaY6
q9UONDEbOh7Nm2ez/mOPQBFE1ysSJuxG918l12/Bn14JsCDsFAQ7niU0leC6LVxJ
2J0L4+xD00GY5wwcYkCFiv75fX7XVGdeBZOefwhxYn02EuQlHSBrQZPlTLTLp/Wg
IJenYepq51bbOqSwHCXs7TpNnl7bNBU2Gkt3Xxi/LBb/tw9nciuXVu/OwbIwz6KK
HZxRwNup1F626FBg46EiXq+1bMa5AN/krIRB7v0Vy8Cjv/2oGTMkzuZe2qCNGGxG
+d1kgNPLd26ULofVCPdE571SQhnjTrQlxYoIyZ3S4/wBh24AnKSORwM4NmgnC4V2
aiWO+RxJyjiEDVZo+rTS6smK8QsBb8ShXr/IyD4+0U0pEoPLlfsC2tPHDXrz9GoC
8lN1knsLtEyQwIN+B/v328URblr6n3CZ6SyV7w7GuKRRfNlPMCOqrdC8gccmE+ox
SDDnNAoLcIjroUBlVixDm5EhzPHHLP8G3+9dJGG4/fjII2fw+TFRWDj9Szr9fYC4
EF0UeHQjL5btCQy941U/K8LySuRgUczaY0MAq+exCEpPp5vwjUA4G1Y4A2HYnb2l
JBvABYsFxogI094hoYL/N/jXIfelnusdQFSrhNe9WIghz07IdV0yNHCZ93DVA3Ga
iqz5iuljgtfy/6UYEvA71Q0RiW2UKWeSQ6YADZ5JiACTs7Om23+RSMifY5tpIekM
sIX4bkdJzZveURmklLB+4kd6pw007H6BuooWiNydGarDaWU4aD/aB978sbgM8zGc
R5Wkqk/PLhWDX1lQjdyyQ4kc/yb81SHD1+XoRm1XrSqa0XHSF8zmsCX9HqHZGbbB
J9rOfKJxLKn88Gaf4MzJCs+76hLu8J1DW46MOezPV9VTwtYTD8dmP3w6GMpbH0DN
/fUsemJ9KODGxWJ4UJ6jZJyZT3uVwQxZdhGLEDM3JNm3WO5ej6CeON09HK1Dijza
UpjtTt81GtXaBWRcnHQyJZEU7Ofvtq4dXOfD7d1lxmKVL5qvr7l53iL3dgyoV98g
nhgPkSAyx9YMvQa6H3ZvH30z0NbVvhea5VQFRlpD/VKmlGIFXFlScNf852E9c+qM
T44wrxT8xyPdaPg3EGNKDE7MDmLaA8ldPO6UwGcIiz1GUzK5k5xv6mTlTGosHzvG
gSDuxx1YeE+cFxgnUvxp6GB3YH5fEHIUQj00t+8u3w707ANHlYUE0Kr3CcsJGIhT
MLRF9CZAn44l1qU+8kj1bJ4dHU29L/8W1yiHlcZuAdcI9fHxZ/wpKhyIKSGr35Z5
K5OKpPVRnP+ZCvoT8QsY5jIncRs2zDpwb/nlwXeeVLkG+REgvZ3jhyG+mF4+oc+A
AJyz44hZS5m0ESMSS9Wx0qfvqBjF3dZDdSQzR9hmq36uSjVltFlVfqLvignJOfXA
cGHaH+KOJmn4uxPx/TA9qIWSDEEzLGDY3BoT86t32RU314MpUAhGPWXU7hcZXnrd
e9pY0fTcLpYtCobCT0OUPgxGeNZz3OykwVXn7MEicEuwv0QyDUoxY3O4BzjSVpFp
8bKxqb/IQy0cHhzvnitTTI39ftJfE3jXxjBpv9wvlApI0ZJ752/0NgrsLz96gQUh
GpK4CQ9WETnHAn4GrYHgIP89wsEU+agkKggA5IXT18Fc1SIKFi3RqryDgf0owKUz
a6MSTe2cZE9pgONfM17BbLtN89EBm1oO/mwNNEM9kfM0Kp3BXcBCobVyZX4wiKWA
U7WuzKATgHZvamdsGrKN9JAw/5AHCmaVAXALj2N/PxSRK/jr6l2DVM/DlL1Gd3Do
SRlLUdkChsnprQXbfeMtoj4BWRWzrKgbpO++RqM9q/WaRUni3JJBQcAcqE6fl7u6
/1FETiewODlFES4/XdneBAgrTFeHUW3/PRlJp/aWgeNiEupKN9O46qvF7OR61CRN
dtZtK/ERxGJj15pLN2f/i8wEdwfgbZFjQ43zWZ8yMGWeJ3OeBDbAsDveDWy5bLX4
SNpbrbgira0+cKvmnWOSXtwDH9LG2p6ydg79uSqioKgezjsM2Zr14s4WYGxoOPv7
bMg8eUkAGtXwB5/faLU3obfGTWVPZ7HZrgblP+nmlQ+ddYBGJhsC7k+QGxEe43IV
eK0qipXmupgNbYdBxE2kQjf1kTWpFncT0CCPN/EWBLi3ZID0+4Dv2B8+DSoQ4yD5
UdwRjJx2npfPh93j7iBbN1NzBkASglG/63YQL4XmTFHXPcXlEOOs4qiYmzB+4hV1
En72bWN1baiQgQBgF1ZCqma1B9IJoeDh4mFR5M/jPnino+3Hb0C0fL9g7rcBe2YI
j+YZi92KtcKKiiA5oXMn6bdhuQOcKZ/J+7kGbfLX06jeigyeRHTnlJcngPh/BiMp
6lLlJh+xDvlZ8ohEUL2PcL2yIs4TaVugQvh6dGfE3ivQaoajCh5GJ+tbHUp+3va3
rYdKWSqbqnIbp/xCUdoTCKir9SKO/KsUsjwfSqOi0+vMAFR6h6uI1SfHV+G1am4L
WFmnJFRYq25REGBN1c5kVMBFjsB2T2GFoU6H0NPwoCWm3XXNj3D0oQrMJY5vh64f
+fAQ1Fi9C+qArz69TT5zeT9WABRr2KsXH3KEMM4VzU6sysKQL76EGIY3TV80j8bL
3zv46+aJ92EqQqbBneR4GNQzvydLI0z1ulFf83PniFfbMRHNLMHwfIFz1EqZo7+o
NWdrilNIkPL94A0CIe9uZywj8GJL1Rg5g+ov0Omgnh+lwnM2ww0bepheeBF6isGU
rCvODi77jaACXDrBZKyeIQLMEzd+v2cEvj38SkQjUtWN1uQHs/bqf+zQklaxQTRP
tAzkX4b47j85ndEcn03047Bex/4ZYvgWu2n59FyKlpU+W2CyIwfUT4qTOOss6R3P
lP2E9hoy+GwAqgCFLw2D9F6Jgcg8Jqam9suEvQh0VXT4S/LjI7fAY5UgcovA9rMD
BBMW0gpEpDndwa9NqgYjbUTTwN1Bl2VYdiz04gfm3iFFMbGr6qrXrvAZT56098Tf
UGsAIt5yBkUlzgAlH56SYRKQSqN/vb8CHOXHh3F7FBrQCDid3MHrZMzjCL//NRZ+
OlPJwX9AQKEnD4z7ADIgEm0qPNstLw6Jgpgn/rEtSaCWGty+gnKIeTUuK2TOCve7
xyXOEAWg9dDwT0mnwe+PX+SZr/VVCMi8kHv9qk3vFmOrSFBVpq0evkl4Pgqb25KM
fJqO9KUG8J+qGJMofY1ZM8Eec9DDfd2KwXaPDitgUw9Tkn3r5QAnqTBRq0T5afZu
VV6gzNEMP7MuHzqlLScYdjt1BPs0aQx6GZnqvI1N3M4PlGOGr/k6wBspyov6hhvs
9XakO5r5IL+22dSy4nVCsjE8NWL7mT+gVOnZ6rvDoROveS0PLM9n62b/vc0+SCdh
s9XdrP/s21Knxa232V/e20XZAP5BvSY3bXa+LJVk4b2qTTGIz4gCk40ia3SmSRbO
uRPvUD3aYcEwzMny2mHxoUjoyd9aLadSezr7NIPjCzohjy5rIUjXA8kKD36dYwtI
vwK7b52+Q+poxqZlVvIaE2ALQzNA06yFhynnCQW98312BsHCql8mGtOXVRuSvmZw
wANrDIWS/JMIGkBzr544VhqXruLZbnrX9G43pdnvagVV0rIV7d2dAfOZ63hZ6Moi
H8rTNly+vKDCOWZET8i2xNMzTF8xxKlft6jZM+HPytAVVGSIQ53S9rdWQEjV8Ehf
fta4wOrl8ruhhbLKKh5NrioSmqIkXytAtpJAInLunpY+HtN9vLKnoDOMwCZRdQJn
/9fB8bhp+Z1wZsHgohW2ovppRBlPX8eekmttxl+4M44eiiU9pPbwYMyIdGszDkqY
z2Js6pd644iggjRxmcAccq/1c1vR4TDvkaR1jOqZk6O5lcLSE8SN9ODeX+Syz87p
DvSrmdSwcUrxWcKiCBoz5pNnjkz9sHzUKZh/ZKxalWSI/Iya1/69ltPqkdhA4p3I
tctbbEn0lZcy36VC2HwDXfYDK8liv9S6KNfTdKRVdfmMKThBrR3EF7t6OMk43xbr
C7dy8yrvR8bzkWtfkEYXSDc3YfK0mskeRbDn1J7h/RnB+TcUOUUM+Y8v3q/9CPRU
4dGIa1kBpWvYR3PR5dIxv7RdHkYDWSIyL8vx68D3MjEQG5PmCVOe+a4/SadvLItd
VRq3KD+zuu1mnnnXT/BB1/LjeM8XdOFy3hZ1X0sPUThw6qUaFrU6cGapie5Kh+Cq
U+BOqhZUcN9eGdmNym3xqGrm6u285JKMpSHCgqCnkpOPtro5PB2FIJH1NPgjtb7X
Sum3A61wKsShgb+TBGips4tGk/C/mlSzuXXKAPIfda3X6MzWHv3joy0K6qtQmgN3
ssNg4kP1xasJuai4iAXS1elEVWf1PaMEcb1w1Tp0Iln9JzsbuxRxdAdSMGyuozfS
8tn7qpC0oaSTFbwZfqCbm3ZT3u4jT0hKEMZWJ4OPqPt0BL6B2eYT/15io27pChu+
F7/kkmj3aUFIMPj9+iV2S9n7teKEQ8h76qssm8Oh50qp12/zG3vitxIFEDZDAeah
3tYvAPgp5BXq3jNwAlWSMYYs+bgSVwUcOv7a24TQmEWUQmGjH/ptqhBmDM6q16I3
1mcu3z/snaCYFyMNAz2tdDMpeLFBVqFCWDhc/yIVuEDiYDgu/v4YTNsQlfMyZG6F
A0H+np4m9/jKr/m3k5D0iiIfLPwrOLp8exsuBDz9ge42IaOCEhtHReTaIYRIyH7c
U6Amy3/EepsJVOJbYDxt3FTdiqLPuXfD9HVhYEl3HQSys8ulXsRogVvU9EYHNhEL
B4BHEqjfYzbLQNkDtj5OjYWIxJaoo/yPq/dCkREJlUtENr0EqxUrxANW9JlpQ1So
O8iXWSs+sM8Ofc3MibRF/RpQJIdA5ul7kA/e46Vq7jYufNn5aUnLZXbdeyib+8kO
QFGp31SAjh9HhwtTFrS8iXZZ92PDInq51MRmepWm7vj/kzhxLEGVoOY5Tv8owiS8
qnQCQaOiSXFPQY4VdXOBhFCuPo1GzrMh7Xg5j7iA4v4n3A7yJs+6nM4ixviUvcEJ
WFP8GVKuB2vMp9AQvmDp7JU9FMJ22GqGlZN3eSU/veqG7Jful+DPo7M00OARUtBr
CihWYqDl3D5v7C9xWNyIGo2C5F/5l91qvJQ3i/YF/oTEgsQYCZR+0DN8DUncpIDy
XyBY1GakTiF4rhJVf9d1Bdg4f5LOqYbD9ZOfBzsTA4EiG0vMbDLDj/1K8SRlKTp6
7m0YwWOmHzQSoK5jBf6f/of147t/1/6zo6ZcFdhBcmTvVES7KLUrs1/WK8iBq/BH
bt8uUvOcFrb4BXmGXExUUPsAAS8DMl/nnjD32ichRdDjtnjC8+wDsaNPlxzqeIYK
KC6OAoLGZLyYAROfKUUvMRbVe/btse5g0HQNMBWkhnl3h70yDKfzq8w7OwQY/kG+
YidM0lq7yZsqueCms7R8SUeLFjT7OsZHC9JoXRGbDCI9n21kZWQeEGTPg6NyKenA
p9hKnzF2bGNV46g6wGE4Euqo84WJt8/nmo2xcULqjIcCmzEBCZaASs7GTXFwbIDA
8XpJxEj76PY6D8wXb8926Cj0ztFyyIqPZ61sP2m3Daa3eYw0e+9ZovNLowHm/1Gl
r26SuDnplCXUNnzEdRtLAVQ094vDTLERDqpASilfInEucMz7pXNdJaNBsd/SKrop
2PcoqD5ZezDkngbSLSymmQ5viCj8gSbRIrBCwe4FT5e84d9WDJf3NqaTguseXd+U
jgOdInNvKVZyVLM1BOpmTDF+6zzveww4nWflKB46Oa5RYGRU+axTSaC1d05VBNvB
mJe9AICDe2JZIlL5dOX8yHvX1SoPGOsOlisBsAKjjBED4ppDuGZV8t+ELJiRc0+J
d8wQMMzEB7ILoZlMxhL2Nqfz6IjOUgqasEZ6KNs8mHgrrblONnlBqQ0Uhie+70Rl
NDkSdzKM4SAannPOqBLIoH23VOms0QYxpY5ijZ4pVXAHL68yvLXHgX2BAc0mbDV3
jR06UC7rQOoHMcCNrksKSZQ1q6s0+WFKEaXw6dEHtZR3a3qE8bdeJizbY0JmHLnd
h77Qv2XFrQ3nAaAmLhnnXOQIYtIhM0MuTOvI3YYwNWr3WhB4o+quk8D3d8EmOk9V
4FwBV2aKC8tQ4HrtNeS6SWFvXGXa2XGQkGF/7Oqns0hj5/os/mCUd1lKkd37z2nj
0wh8zKZpymsxSVOHKJnLbwxfK7N1lS+LyMFGVR9rCoCsXFvHZpGbyl6Tp6x1PF2O
xeqgu/tge6DOSfTxGWpJcSTBVwB2A1aFlLPUVV0xP2f/vblpYt9SCxw2pbaQEUO5
imc/r1M2dsFzE6wvHxpVTKoJGQtE9uVTXghxxNS6dQE3JM+4iQo/ct7x77Nrbr7l
CVpXzwhV0kJbDnOfId6Jkv9sME/ejyJ4e2RQUdgRqYeSIY2dgcdh5oHZN4MMejaP
safnBRxBJHqEbU1eamwl7brRE/dJPqruzT0Vi6/zUeOO5/V91IEV2ZGLNWNPxs+7
rSz9DRMCXMdda5NNKhK6NjCgEq6cENdm4a+A+vwszWNshZjOZzoS2619ZHzLPPVk
hnAkkfJIHegyIjmlWPomj1RiaGurvRlE564W36ljU10QmqtpWGqoG7eNUI1gYZmI
nXv3gn+hEmZHc0fwa8b5wF1Z+EbyDCZxn3YHjgi8pw/i/4QL3mOojIMq1fN89qOA
HE0gpE4io3MqzBbnNk+gqWiOcMZsQV+w739vmlSwlO7b1Iy7ahIeeH9iWHCEWNSQ
XYlNksKu40HD4ZRgP1SkRwOHwIbwARRDzGiZ00tIvTcluGo0RlLTlF/+4VSRkBAQ
hsGbR/NaL7umvnCCtzQPZT8MQ9AhLRPO76mqgrWBp1ceOobZfWtesUKVQpPhPBfd
uHAdCYnyt0e6XstWRMKlbLDhyJvxvQx6dHlgY0aJKfQSxy6SSOkS1UOwwV+u9s2B
rBLgLE/5kfSvlYD8oCC2iQLdBMrEDj2iXkMEzHmv3Us6ee9HVEXtXe7Jku0SIIzf
a8Gqa0p2WvQwdJoCe+eke8s1ARmC8Two9tv5nC7meU6boA9nmv3m59fPC5cJ+ogo
6C04tX9aLOhCOF1j399+Pma5O4iP48sjiHwqgEO24q4cvtnIiJCtrJwtnjSCXIbg
jSSN7aXUd21EyPQEVxInmbueqRZIA4BghAyiviNsUMT3Nm87q1P0JC9RN5i0Qt5X
6xTfWsu8lRfjMSgqZEK9D90Im7Z913qquny9DsAGo6ZOrLfo4FFmPo9OB5viFZ34
zZDkpxyoTVTvmOV4HzuhCjA5BWxxDycEcmkG/c2wlh5nPfQA2m84L2WyPqGp0oco
EQwnyu8nPtLk6i8azyQs6mBgYDx6VN4iuc1nu/R8vXPJVFgq12oq4Cvhku30xNx6
1SZUBKB74actcDrwfIu5qsnQt2zWAVpQ5sUS8smF4vEJdJ2gD+/1t6d/rDQKD+Ru
DvMSCOF+uyKGh8BxZGxwMncUBKmtkn2NKGW/EI7AjG92NS/ERJS6EWMPbLFSErVF
PskW47DAp8gXFqFFzZbO0TXJ+DqxNdpnjlToi1j4BghzS/jLFtIzQx0zk3m+fCzi
A6m46RoAN1FSWGRM7qfN5Zto3K+6yYOyhhliFv+lGCrtOTZPZq3nXE6oG4691XCT
3A04p2LupZyZx4FweuC3v6EdZaStopOTjieEwhCo7hXW0K9VnW9C9RtWMN062M2G
hsT2R/ajq42fU7ef9Cq+qFFQtynArPMK7mdgB07frJDpYrxv58tRVF3/+3GH0HS3
CvmYpIOQjDZhEGDnF7kddjpdJ2ZOE7Q5MDs2UnDLVn+eZzduyhldwaZl9MSTlfoV
HzMCjV4Ul7Xh0URgQcGul2+MUO5Lh6TgOL+zAmb+1bBCaa0sZFzgxEP5b72dwNDR
z1X6xmIfUXHSqi/q9n/C5ZhzpTO/iYVTb6btVaz+UclFcNo+1sWF5umPCU3ylVk5
CpROZqBL6AB1YXJtP8kSxsismr6qij/VYi93Qds5yRha2uGZmPLuGO0kcMnZTPG/
uyMl6dENZQBcRV5G4HC8VT7x3Tw5Sr104IkKuOSvORkfs/+1sGO4aoMyPm72W4X7
6Gaw6fD6/AakkldXwIEDKDUJ6T+4UtUUnUts3v6ABI40Qmb3VtZrAnaITtTQ5vey
bcPAF5VMBx+CAaoLtx0kn1AnMsH9Kf+5Gpi968sbWo6qFrYz7fB5TEAWf6yTQzNO
3+UPr0dRAHcPIp9svcLsojIr25PmnoES1+7dx8l4AT7zDGxWtUGbYrU4jdrffEGy
0mMkmhGGcGCCCqwmUm/ty20vI3rKimgEbg82QNgxALkTlm3WBU8zJxATKjwieqZl
g1gaS2etmOvWlOa5JiWZrNiSNlshyhTlO7W+6D5gA0phOHrEBi636SDa8GTi/gZv
5JP1s4ePO6hkoPHOIJTDf6YHOfnvGym9uiTcruTsCxsejrwLuuN3PBClQNfTOebb
JGf1MdG1cdKxGfIrlHVzDrhADJ6jwotuAOQgO9wadcEdJlebYoA5tUTSdNSxiyvd
uAsgaqp25DhE5znfhXjj2JINh/DqoH/KOZbz6K4nGKcZ+VpwQKpfgtn0ddUnQlFZ
5ND6z8Ero8Q+RRtYCm7Y73waikWiBOoesYrMnedn/JoZ7AfG/Xe21LTcXsjmH89u
k6kogKkR7ot3YPtvca3IPJBDAGK78iCM6bb1DQNQUiiIK3O3UhlGZvZvlLDQuiCU
ibQdCvjO7LBOrwNb1wZrzCIqQUuldp9xWvWUj5HNuh7GEfAQvy8PI0UFjePi8hH8
AbG3TeNmoRxAEK7FopMFWyKMxMj8ZWn/Z9wk9SXg75uErh84nca7CnHp/ozhKHjZ
J239OwnT+NP/fWNgWMCft+EKkhrJIc0p07j1m8PthCBBU4maYgv5brej3l6PoQAU
9/RmXSV+g7b5nKoHWZ5+Fbi2hvX9xuMs1Uqk+hTk2BvBpX0XME7uoNUHEFSxSX2X
i26NDbHqE+NdFXpgvwzjVGvpR3dgyxOjRj6z8CqF9JbEjNY0nsOVRjthgbFN0Em7
F1r1O78+hMxgk9ebea80pM11Egx6NmO7H0VUsxNUTpjseEyE/1iyUfBxeWhrLaZ+
KfmK3xUrXXOUyZYn5GYKskAsKBwaJjSYa9YrEhEGdlhcMMBibdYlNPHWYXWq+pYH
gD5zjqYmWr8/MoJDm5IsTJibjchOTltoNUMAf3FxNiTOjouuO7hd8Sr/IoID5qz+
vtbQW1/8RqMczMiEJAJ32o58q5TUXYKGvM3OVmgMTkpU/opSCIloYEVvCEXlJGLf
bggULPaMCI8TzH7PoqHbECuDKw+S+StC0GTRZtix1e2ljVTAvUldV1wVujt3a1bZ
2yuAI78krRmMzWwxYfi5umLw4bIIXk4vjI/la3qK52HEOquN9sAdAucmIfsyui1E
UsRxc9qaty1tLMN2/v9P5/ljHzXh2h0kZkGWs1AM/d4EJrY44dHA8xz0vSF9APud
YRv3qfjOPYe4fAp4+K2byb2qnJxTFqyVanxhMQf6ifqB4J+PILyxHR9e0CZbwfu+
CVr1eyi1HUg0LV+978s/2JMlndHvyeoIdU2g+NDTibXNNnmATUHcTXk7BqP5rp7V
CYQqdioUVzQJBRQPlZUf7be89IBtl58gqZX3ZejBBxLeDxOAC2Zcd+cV4gXsHZM8
ieqDdQPQzeHqXSKVPT88ARmBPkQQirfnaoHcuEjiEUwTf0r9R+ceowPbpokmnha3
WQRs27ad3NnOiqt9lyQJxFyUoPlfN4tKVYlf8WIoPp2Zere7tjvF+aPWLsMWKHk8
wd15IpFxEY8gwaG3YMd5vmqtV+u84Dx32IUgEz8Bme4VOZut6Izee7Kw0uvZX9FC
/qWgxO61vQ5aovIzbTqVb4LZSB+i0swdn5UkACBthk41A/8fRIgPxsH5/SnzfcFf
iDIpZaykdxeHiFlc5tHYnemq3Cgg5bC2UcOKK1SXdI8wOvhe1fVdKFQWOph7ebwt
lOp35yS8D67zi3phC3YK7diWAOAVOJbqaSC1e8fc35rYkx/iImiM+wwBKttqWrx0
koxhZiyfxkpn8+m51J+P3Y7+wzTDDu67ZDd3APvYwanXZCdeZpG4J+cYeEFfin5t
6ltFn6JOtHvdMWEPLAzh/xtfpz0pVBFYU+NIFjSBP6V/K7MuZ2uIsRfJdUn45m8h
/2f35i3iRRfQGtSGz+b886zzG5KjAOttDxRFUVDqP49Mzj6aKuKwpr8QOsnQn6M6
1cQFnmRbt3mkJbSlHHHEgsmyi4KMpmMh/WkrBrXItSHanfWR44aqaqxjNak/+kMZ
8H4VVok4oYqNodglW0MR27r6HpcOEigQFAD5i0h8W93ZbXIu30XOY94JghC3DkU/
KgMBWba6De1jMKyFKny4rYPsM/Bg9TSkpVIYfchhrct3d7J8kZ416rnF1QL8XIk9
uVultV17hRxL2YRhaXKa3aXismbS6V7FtCI7q0H8h5wKekR4Pj2hMRAlo/pImR6n
R274gKU6T6FlPQZZIQJCW7ZzQxPEvmpZfWKFcQQlMMVKjR8QyqWEZ/xcs240/B+9
k4sjuzQHbOyGOk3ABwlcMdEeG9FyeURjwg5xlVcS7Oj9b7GS15ka9DfDoZlthf2e
U2dcbMsifOprZ1mA6vgXxlSJPO4xRroAhzHdPUo6/vycMg+qDX8GObHSss7cL1OI
p76LAEJu/iClKsm5wlKmekkWDf+xxW2fejKtq2j1w1/NWSzTO0hSro2MUogM7+q9
dT9eQlJStr1gc3Pezox7LXIuthGwa7a7f9Rhy7mMfKOukJ00xdM5erOGGPAhAbOu
/qJAanxNNfmN6+E7ggsXjesGxNEYgDDAWUGCWlMjvP/q490hvUIlOCz72/KXTjVU
I7EfwKqHJpzPylEnlV+xwSY0BBeCNZok/h7cot3tCuITWgJEn/vU9IV+W52r0ehr
STKU+0lwVfCxqxc0A2isKRurjpW3HaKsDtXwUjO8IxGlK3BdqKyfi0YLufv83eFH
BGY9297D2fYefKBOj/nk2MePQ+yz+ysg/I4n1Jqs3O/IJ3AeNhMHDNlPTkTNz0kH
kPbgw14JU/8yDwZ7BMiADxTW0Iqvsz9XaKsn9W+gYMGjiI8lyjEMz9LJ504HZHSo
w06WW82eCPmlZB1k5SgasQE4Il7nLr53GgSoveAeEG/WZdZYMOb9mvstgBf+TJTK
ZL0dLGdR6DDBQ9oVvvZQGJrIjxBI/rCgPqeG5O6VcxXohnQ4KvPiwv+bI+dk7bwt
ynAwZ5yyIXVIns/ME4uL9n1G702lq5z/cRqzRk7BHx+uj0Kfxsy4Tg1DVKI5IJk0
DXSwoyVKkDCn28WBYz88hgYYgxn92s6Zcu4wokq6wTNDE0mLo1flXaHK+/1vVQMh
2ot1oeIhFa5O9luKI2kcqtBId09TDJXRRSgEkFIsBT/s645bMQH3S6tQvpSv0xYh
/0LeJVx+m9ZILUSAbYAf3vpgAX9fP7QAOHQ/5qXRYK27CStZ3MhV2uJCCtt3Iq1F
bemuec8rLP7Cu12UvvwLGtJTZ1JRunUuNRRmPVrH5x2oRsvRfzpp9ewRp8T8Uspx
ef93W4kE1HFkqLZcfD5rRxLSXQXlrvrmEW8ePlxf6BHADXYUPSJ2cte+prUVYoCA
Mr8d26T4rCsw3Q7iowGsKBOxvsTG7vqIS3CcmLN6CJw2G2N7oNBOwBEvOszjBqLB
l8dt2iVkyZp5YxApWAtKT4mqEyMaWd12llIBBXhNmmv36enXU7vdQ/iAo/btkXTl
HLpGTl2aaCkR00VYfRcQbjmzt985ECGKytTiIF6mH6yDdqirj+ElXEzfB/NDvunJ
kbHfnOtoeYl+/+qKvr5D8Y7NUE0J3wLniU8z+PkWEVeRoZ5kdA8XlcV7MF4km91E
DnmZWF2SBUwlUV6UbJC5w2Dv2g9sDPbnhIol4MjDq2NMuSDjYPwmZV19ZjVp9MVb
RMNLkSIKZ61OSJ/ghpGoFPE+xHw0RIBrjtlTeqC2Tmi7JJPCeJ0urnlFk4ZjPOAy
a7VVxOzE7iXAM/zLcFMcULP5LOenD9qyhT6Z+nHMWvWKdfua1lYiyld+/P9LC6GF
2QNgx24zEDdf2oNX1m3T97ex29reOVh+p1WZnRYMXiwewWVe5o4VQ0XPDDDYPkbU
r33yH2bLb5HpM3kMCeldSuID9YApo9EOI2MRMu+YgLKqfqDH87wTjBVWnKuQf9wh
8mx7yWWPV3E1y53dgGPu2ov1PdLfL7pGbTIkfjTcynLMzz9A2E8xSWc3EofHAgfP
Q4aONI8NQ7uEj2TUB5QxymFNCZ47kGy0r4dMOeTrfboOaoXItWi+Sqa4hyVWy65B
zCY1fs8Y7fH0HEEGeBT9e2pQ+b3k4otgHXhLuJqRbyBNRftknKf80CjSM+up1Zo7
axahUdkMF43nR1VQkJWZ+qm6WTT0DOHiJ1FJ6HC8gyPwkeB2H9ziKToMUC+QdCZi
oLbXMPv2OMDZO+l/eUWfWPRitwITf9BLdB8uaTJ281KzBrDx40cEtTUdLQJIKfHI
QARQLs5Ysuv5nc5qQbFyvoMWTDEls99B491ObVf0iKt5BvpWxmDqjwZDVq1i3Tqm
OqN2SLFw4jPKJtY1141+ZttGSxIOm8VxvyCBt/DUWWxQgoDy6iWzK0Tp4jB7jgxU
WJiFoD1kifue+Qk5IEyIMAtZxPs2lGRY4tnvDxlRWbgHiaVrudQg7yVHPAwQx3o2
FY7YlJqQObL6QUrZOpPTH/MmtP35JYjarVRoyDyb89M8Y5FOTB/JTCFyAk0K8ZrR
arVlN+Lv/ZKBMSOVr9XXT+w4hkhCOsKAfNqZvbrQ7JvRZn+mdRsLZ/2699yLz7sY
OK/d4QgDEdY+RCZAnmcgfbaSZRJCTb3yGtFeBIACf1qeGk/ob23w1ZOFfNWAx5XW
x9kwuKl8zdLw0kQ2Mfj94aBY8y4agoeQcHyeO5jB2dEFF1aO5FGd1iL4h1EATQoI
ptVG6ChjgrEpHV5tVjFuvxFd8rRvRXt/6oCdUk8q231Gl1bW9n90bWwFV3hn0rbB
1xP1T+QLzEgPa8ho9H+V/OaoQfeP1vnl66hrH65zGpTIvZPcmmKtZeZvPR2vtsp6
u/JeLqvDirkNzdvk5My2xUAKxyTFaVimszowgjZFtpT/aFx8VROoxV31UZnjAle1
0zvjl56D7uLEj8eCbAIVYz0+6g7UNgdu8w+iUrUwiFkyUxQzPZ+/j5kzg0tD4nvg
OuXRm7A3yr0yS0ErwwOJkiGJlRnUilwSSDJkG4HR7wW0ecUJd/Bx1nOBhTeJqvIm
xNjVlJix1aWq7Soj/k5yRrIg7bHBWb5xbhTpeVZwaooWZ4XClM0yR8FGPQZjMQtt
blWmowGhaiL1J3Rcpa+NMdqsCD1JAPKCAltuXg4y8ErRkl9ppsymGd4OoEmgP0YB
bEyV6d1FDI22gjo/U7xYEyr221GC40066TUpcrCpaMIddwK3rf1OMrQmOA6ypb7B
Ezuff8+MGQbtpOLhMNlKi3PJIKSbXdxQSFlV+j01JBA5/yjssZuK3G4iE5jCBa/I
U2pEokKMygHTO+cf1rvtK86m109tl2d8uiSdQe6Ig9a3cMRnVufZjSUnZ+YRHOqO
01NhNKDLKull17qx2S0KcpwQXDfLQubaaBN5L6l3VBo/bfAoqN9SKO18IWShJHUp
xeTnMloL9nGsglNUS10aIXzcwk2RF09tneAQ7E5e4Vg/t3wbllCyl2lAqwKqtNEx
y3QCERek+t3RZ70H2zACbDIbRVs89NGVM1jC30mbPGS79Sxh0hLOETIwAsJtP9S2
4vrv28fyQDo6dm09g59brCDY2saZc59GcVrCtuSkQfaDeEuD7nRxb4GYKSAL6JN2
Lka/Btf4ISa2JzOSQxKp1LILVQSxN+vWhxj8eI8JdQUcRbfCCpKWOhzNj4Cr8Evs
PrqCmFzVQN9pfhFLjE2YBC8eB/1ijh7S5DUKki5XmkOmmF5RfoOzFr0sUxv59j18
+2umIRHa+EB+H4Dhc1eNiLfkM7HkVTTx+OWZ75nB6GUrD7iawRRXcWcY717R1yP/
Nb1wDo2cF+wqt+8CpF7yWEihaR8+IfO+Na+k4eC8fYQTn7pCm6kYLNshkKw0w2SW
zgbX32gYsiPD94Wn5kDquIp+SLzKEstvYpOncH0p5p5dArmaBKtN6ccKbyxPOH34
mySeXqE23ytPrh2FVa9JgmuX5d2uG0/LKb8lKf7ttZMta8o4R6luid2ZraSQx14W
i9rjzcnA2gfwit7YpkoJMOnuJ2HatFxcxrZLi4yBL9XFncu3TSQYC5Jf0KDGVbC9
j6ZYy/3J9mxyDAdo3Zh2j2Fr5e1SjA9D7AoMEEB++2g3DMCGLadxxUBw/O/9kcEq
pvFu7aM9Tm65ymeNxk96UYUwgks5l7XdFLsT0PM9e6PlhEhm1dz9lSvBJhOrdNtG
MmQcvN6YEpvr5wrDQbmHOoQ7qD2p5ODdkyWrWpsRgZlxxpLOp8617wS7S1G/aU7d
tm0CTDazBTnxCCB0woXuZ5t4TKiq65lR50l9ar5FBIFrkYabiLmfE9TuHFH9yZG4
TzEl/CPS5Nffa45CJiWwT5T3NKNcVD2hJ12xD95yhCpQkgYd2DkEaxU0o3o5IYj5
C/95owhuNzXYOKmMkNyrsyoDMLkmQ+kTPmFfGl0SNHyqK+SPtGHP9FxfP/1x/QwT
hd929cN0Kd30oz7MJqPScHctIMKY8PeOVfWhyJhP8joweOeyfsQeiwfSSBLXwraP
txgSGuKwXCjesb1ZVF1XrfIs4+zsdXiBGOl/4Kktfb/nEVGtbDjoVlNDf33Km+Tf
yPBjN94dsDuYys/tIZuxq2Jk0BpKRJqTwAFt06oiU6JN1WK45LvVepJhIPmKgmXD
Yb78j0nb6pf0AecE+LLDbbug07p6vp5x47QuiRpCuKw8/aiYwELEprpkD0mVaf2R
9diNvCQj6r95aU6LWOOwiPw6/sKbQ6KhKqe5IdIu9nBkDFHBGv801ql5Rj4AuMNa
K3u5B0ceykzRfnZNpocrEaHAE/J94CUuTBnopFn75n0RXXTVQXvZOojgS2j4mUkK
r0Kzj0JRMD6Bz8MPvSd4zjF0EgQvMPITT+nTqrg+SnG/o13ZK1i+SpdjjcU7Q0oJ
MgDhQRIxUg5UOMfznHsD/QYeiPP9x8naZN+2QQcj5qgtfsTTblrwF4x+m4j0WIJg
murHtv7Gblyyu15KEg9iZDXeIsBUMreKw/WotF+B/9rxDFOxuUo0IuV9C34AFMt8
LDFNzAiCh6ZBNXpZBBEDQppb2zhtxcHappQRYiT3eSCx8yBGPJEvURiwXPhEM6kQ
TmXsRmxVhSJalLb9ktU1TGxwge94pvY2vdjnRZGXOJQUtS0U5lbOpCQ/Hs+kPurG
KTqZwPBmXW6R5e+TWX4o/hHVejY+Avv8nmBz73JFE665xy9FNCWGtdBZOb4YV20H
tOu01w0mEEnXUdqIwV0QgkQ58McJ6U0zwVv950rX0TwDxFAy2/5oTNV7k9gXHIN9
e4Ic51ewg6p0bH9uBnjxCJSZXPVp0IPdNIjyVR6ilELFULvcr651ThG2cwPU3+ZP
7FzlTYgPQjPFxlinRodQkPfz8MBJn+qOG7nMqLoeN+5INuupNkHb4lUSr4MsAdmz
ByNFnC60UaUdXwMg5gmCd9LxSZ43BH2298ZMQlgFKqL8vWGvZxh6HVxmGg06BrSl
AwJTirBuGK4d1u8pG/CCIfWgqY+KBEP0ZMz0w+OfpBZ9+xW4Yao+n6Sa2QzmQxcX
2tujfE4HRo2Mf6lK0RQU7EmlzRlok8u4UdM6gGU/Zlz0ztgVkK328L+cWAeohKId
he0GX+0M4YKpOWvpjjrSZLLaO8JkeD7AuaBoJtmJqHhI2eJLtRTc3eMZtcmzKccM
ymiEOITC7k8v6UOgTJwUAlo4j5+c+fKLxqsR1yfwDFpPjX5ZkaUqXFHpe+pXPNc8
hrdyWmEpP62INPuY9818tzsPEMpBXbAaPPA0wNid4g2FCu+8Qays8afZDhLu0nee
+V6bsu6DNkwGDen9Aja8TZaVSWVeAkMFw4E5DwNhWg6vQuyvG4TNe5FOU2rjspkO
j+1ha3wJPP+bTo9jn/kqyeFSHiy3iDc/l0FbseklF+txUh+GMILn+OPkllbj0uRf
tkjeCNw3FRDbDp4fdfSpSRR76UAvO/uah/ijaBIaSvstAzRBMxIkrOs6jZ+4gUMF
kmOZF0PV4nYfehZSh/HBtC8tnB2Nhb2bdhkqwm7ax4Wd4564O7D3+MFEr3yYD7LG
kL535/KU9weMaMYfGFhCi1lTEBaAqwaUrty5Mry0rqBgUvneO7Gn0l/Fnzeml5wf
kqPJjAneLw4Sln+q3V58dHkk3WiKAnM4fAqlRZ1hZfQ99dMGs9kuPChmuXoL1GQA
ueiR9QB6Xfa6NJGiH5k/gDTAW8GuqQBXq90hk2quQdgIcgvXQ1riCZaX3MZ7SH7A
9Ls6kX1ZImDsAWpSrsYA173xhCJwEDuwZIIXZ6Y3O6MkltyJPa5wL45KPoCUsuLb
LZT01KNl+zlEwF3UfrPLpiQ+bq65urhZTu/zXi9LnXjRi5oNLBPTaGGLtONv1WT5
e3anbihmJTQ6aP7N+WRnmNvcHRA2aQMLok/D0e9tlDA113qsGzY1IFqoLEnpFh18
Rc2JrAdCSKb+VWvqSPColg+x4JgfOIYd8+P5BFY831fOsQVG5+bJHLEFyqzXAzev
QwmPRKayKoFK2+z/KlTTQ334O53EQVJn6+0O4NqHf4zVQ48F2RU83w5Hs9yls6Iy
kbCB/KlQKatijlrLYhPy8VznSCLmoIh1PPMIs4Vei+tLQUZqkIoQnepSvzUTJERK
RtXFuPEdIf0wL/X1f+i5UHs14xM058TgVe76vssG6jiNciL0IXtwICJJ/nhTx+/9
B5ijvpOCq7QjSGRXxT/Pa/MgWNr0WoaTQ8j+i3PCG+SyycXqsqcgeKsxU2qWupGj
AmXhsAuQavc4XIv1GwJ6OczNT1zHuIp77lKxDL9EtH2Rhe9NSzgx72eo89SKgly5
/u7XOhTGA9e5JF+3+6OXWly5sSFPJrxAZn0nMY+rQh4d9/s/vWPcj4upIZVqlhCd
zX/o+lhvwd4sIt6BL4RBVKYY7bPxdCbXNJ3qUOoKwHHByFcWKZv9TX5C9hr1ASat
PM2NNXdkbZ4TfPgXXTvImR63AO5va2YWKcPYOU0Bon7ytO/mofgDtbWnJrkCKhGt
S0i6kuDGlCFQR5RQsuH8ZG6JQljszmAhGF1c9QOBiauVGs//FmDHb5CB02l8rg0U
sX4DiB70QX+v0zIf6hy4Atpk4/nePN1AtMui5ZANBCiLNJ3UZqrQlnkIGbfHzksK
ZC1QkrH569DRFakzVPNroJ81xaBpL7z9/H3iWEXUHJ0467iNMhn+EabOsBy1R6z3
c2FUI0uFs8am8kilm73KbGHmk4mqQ1P4HvfDLCA298zpcSWJAXyaWG0xzj2lo+gp
MlrsfemkGnOLwTvv8ykphzZbasEqj0v7ofkRMgr3GtxeWmn1zS4l85dzCI1Vmhtg
OGAIwiyoFeis5qjtyDWf5b0PwQxEZEVOlMXefCYpnF48Ez/gFEzRDSPabwg2n+UQ
hrUYSPW4pmoZorDCImmBOtH7Ic5+PdsUYUsYBllsuSEhpxpp9L1ziFGxFxHboN/2
uWmUqX6+7lpfO8PQrLNSmf3GVH4S+EUcKulrMLglBhdhkb6kB5v3atcCv6FVeCgV
Qxk4NrEWHVF0jeJ/uVMD4WkmJG29FDzGESHx/7iT3Hr8mxXiN+0grNADDtSF1Lbd
gp7DcF4W8Ezu5VVW7PtV9q4OFdLNU9mmcfUk2MO+T7Hc0tytToh/e8R9IE1rxvER
OwyLc26D0r3uRG+g3zWFmDqzcbxjhE3Ao1P8t1ZSWUCyIxHEVFHGheaFKn1hFkxz
gQxy77XGnKwmGYSmKyjlrOtazXFdrE4PePV3Vo4kj5lj0C5FqUM9AyAGGgjiMyzy
zSCbtI8Mmml9vB7hJ6YSWclGg/Iueo4S/iSymF5FVy0awJL76+eEYdoVImENftj6
zRTeQy7x9K+h7R1Hfz5p2RpHy27gQREADnNqFQuU5C1R9GWH6d2UpSan1oAgIR4x
6Cmox6/jKXKxZUzQu/xYauPuGu1D5NpW+/fyxZXmY2td9iB2PNcGT734pUFp8max
YWvE/pTjgLex1Bk5duyp7lrHvJKXI/9zbSdrM7JlcfDQ0n8Q6AUoJ3NODtZcNj+v
s4uEYhQ80fbwdmUppavznVa8S15MdZuwjj+4y/fdWBjh+lf//X6DzhJH1f4vWTfa
9gesE8NN4zOrSAa7e50T1w0vRzRLmVqBmqUTeC0dyEAsXH6ySsi3nZ6sYmzbuBD0
EoezBJcOZUPyGs/QfUwyyCo/aWQwfMuYFGHeI1LVbXeYaaHClAf0pC9x4Q14uNar
aDMpTu9px3bXSeMcS6f7kXRrXxUoA5POS9yvMFV5L/sxaWaGB/P5J2XlPUHKeSOb
tmmDRpbtlHWysZjBu9G+eXOGZRjr8AAMJvI5dcoYkzw8zbutIUkOZpSv9BUrVHcR
aYCXTy5ljNCrIfRAelosakJbBgm7WqSeF6XDNBU779+E8ssnqZBGIonry1GZgA8g
mLXdY7R2uwrSs6ONY2uf+x4ni4OJz8Hf9mQAfo2AAtNyyUe7J9hzzO3WHxSalQVb
PEYifBAJJ9cvc0B1PitsSGE47x5aKK1SJ/pi7UbXGpIBemsGenmrMxwoebzt/Q6n
Y95lm7Wd6OicU8iNpiaCbo0FhX2HR5yd2iVOrAZsd8UHMksWMg//fcW0kCvtxbLp
VewvzL2FyNFi0fZ4fKEhZDYswK3gaYNZiVwId/bDRcJo7bUfzfgWRAxmR4/PbD3e
zRZ3FE0DY2wfY7TwUwW7wqOEBIxgOQF8vmH34u19gLmordQbuNVX+AEIu1i/SSTQ
WruaFQnTfbx2Ax5qUwvb42+5SceOPqQCzYIQ9JHd9Ji2Qs5TM9s3zbfOiMFiU7k/
3d7fGCTDKl5K/+vAsWgMLva7I7rp+hy9znRjdlLLrTpDlYqwim6N0qeUFQCNJ6oo
qos3/wWg7b519RHgRBuU6CJfMl/7ErEMvWRfKnCB0EGYOWEtuWJLfh82Ffnog866
NlmowElTK1gIzdou+ggxEhmWFaEGBWYA4wbdLFJTf2eeESFQSJW9SOG//N6hDPUa
f675OkhAuuXwZyXfSNgyJsS1sPln30AW2pu27LpRrPsUrqVYlc5scrUUS2W1cBJM
m2h6M4K22wryPdnNr+gV35YxcguHcdFqfuOKLSupSbNUDNk15mb8OCpusHI+dcnP
p0OuzL5nuQzurViyRCbOmglpY9Ksf92DwtgBm76tMtRFeDAmd4w/s4PpY3MlLMe6
pUuaCgJtzvgIyU+3ibJsIhv8d1dxilonRiymh3LLL1zQjn4lVp9NALMYXxCjgOxI
9yENFHkDYyYvkqf7S2GRma5teBbaYE5RFp6XixF2DjYk3kCsh04eBlIQ0rn6CRRt
BdjCMffkxIqX5S6bznzqWD063MhBeHDWfEdW432TgSzXNZiBe2aGeNA0FQdbl6qE
QIsUZrJn0jGazi3XlW0+NopwSVPGkY6bXdnSmct2oslDq+KV53ZOBIrrpczkZ/Xg
UXZnVCCymwQWtEoQebKvfv8oeQiCUEaCC4R6NmlvEQUao0Wozfo9irF0TP4i7Kcj
4+fjQ90+bPe2dDS5D8VoG1DnCY2ZCIxpA4ktOLG7i3266hcf+RgyvKt2tsHn4yui
nvs2IOMqlg2ZX/npojbcgG6eo08ccCqeIbyr2LkiODUSSa1FTd8owR8KmUpiPCCC
DPjxFrvLxi567rE9m7qImjYilhxJPYruoaG4J1bX4+8+TmLvWklrqqQkt/HzDAO6
v4EGAigqu7l8uyTKECjFMqiOFn8ns7mdPYP5LFgV79E5KZnNGnlHFtqSiiSU9XZ/
qcNE5G5TkXxA4Sp93TXjDHHqUeaUfC162nO7IcqsZKOYmARliLfT9e7vAy18OONh
+q481aNKBdATWsafZiMa18rmwAZ/ke6VlW16ZduP5djghKFLRDdPAUbCz+JnD9c2
R0W7VylSmfrpwer9Oy7yj5NDmgF/+/DqrdGIq533N3Ln3+phzCSnOJ+UANgUKJwU
36IZP+CvoPs7RLvHg61phLAGfJ5KKidJDi+ZQ+XfhquFIscDIW1hacyfxHsk/U+h
XenVfXjT9m6LbmJkiKQzv3hLVeogA4iURMVIxtNQb3x0JIo+hTfaPAEiy+T034vS
SclhC9Aotg6bQo1tyaz9zkDj1gY5nO+eflvO2F8yANj8lzTcJCXDGuQaqpV2NYXc
0WN9kgDsKJHLH/D3FyE+t4Ouw+3EnsjD6Hx8hpmEb3veuQJKYVbFlcZ79aoGlFiB
vlA0CrK352UGQshFO056HF7mVQKMzNuczZkrHX/ezlr+cvXoLEhtvisvkqDmPBAC
orzjWzDgZAM1hjk6KX5ze5qRdL72FOVey8stRTLr0nKe8pnH9X7g+pb4KbNcivVz
IgZwdoZ+tqQC30GBZr9RiQAacTwiEq8AHAvAfqvEqyWCeZBPumfDx39TaTWxYZes
yKsgmBs4TnWQQ9YZ0ZzX2LvHdjG7AmS2GDQ++DET4cVSAFPLEEEGdOnIrIT9Q2xZ
1/fqsTCuDP5i7NLpKBb7jma5HzAcgwh7qx+uTppvJLtLbOc06boBGdOAYf8c/Il2
yX3NS7GdumXAHvSRRdZvcjjQ8tRSlwsoI/+SFu3o4YE6sa6eZ55yNDINd2cCX64x
56L4HHfTHH3sSy80k6pKfbtcEB8YRYlt/4OlJ3vaY/ZonOJBx5o+Qo5FXes792RY
jACx85PkyK8bAq8gs6ZF1Z33NLusYpn2+mqwaky5HVbX/334em29X7Ziocves8ga
H8EbttbZcO3KI3qEJYNilakUQXXzq5ENoS5ySuJN5TgIXz+vXQ+p6cD0ynDLuk0Q
AGySwXoZcJ57UzB8pccQBGrir/tWh46x0MxkDKmgrCe4fvJLRXzBFqF1m+nL3w8s
arRXQMP8/9LhefPL/egM/x8DZ9EYFBzhxIx1fxMl+RbVF3IZ+fUVnAyJgLcyrp5L
hLc9OQbFyrwc6vzp79FP9SZDSb7tLYjbk31nKp4atdAmqi/tLtveH/EoGELo/tIq
Zqrt9UnJWtshDhdSv7V3HL2wet4rZQPqi3iNiTjxjnaKHAtY1pfTP9FJEEYorh7J
b+Q6qltI58Tyk9Sd8BZDvd1DVevjDMBEfFNgE7TjPdTqnRE1Eo7S1FEkrbEUbrxP
2NjnvxA7f/vxkRuHjvpD5AZTGW93s2kweWfwquTxprQxVuruYAeuRWLIgjsNnJFI
h4fObID4t9xtRCtsESaQuAyc+Hh3OcF3zNXe5umOO4kGLhk67SLNX3fosdfI984b
5vbCmmOlt5MrojhIaqAAgJVIfsKL9NHcn8LD1deonkKna7UPOYDbX05YdRhVqwFo
WzbCz6UgNSSvs/uqWfHOVNIF3ToAGbV+x04RTa57d7ga/grEtJGNv58P2lFb5dWM
qXl53lUtPKJPU0Y7m1gsBe+yy+iI+dOKeuug80XZLYJkvGpfXgbEYsXCwFzq88b9
a0fvTCNuthNbvFqgrlw92QleBfNbURDbicQu6LXpWylcoULBleFlOnk/7stoaP2n
PYpMu8Ztw7QO80+4pUpAapUwR/ECigLEwAqs3CgSuSpUIHTNG6+ny03gZsO4oH9S
LoAOzSdBni8eti7kcVxIcT3SKoRLDYx7G8E0Mn6W/Mj67a4KoEV9hn3oBpkr+XQS
gajak1kH5sg4BW3kTEAeI+ruxoakIrJYdXZqMhqmEH8txFirUyZdiopFMc+mBAnI
iqRqVxyHqIM3y36sGO6rjPijmKQp7/lH3wncduriFWcL9RAmHQW82yl6Heu5H0Uh
/6SeupH0tT/UokqegsNbysD7weEj6AMmgnudqnTmjdXwJmT8sFQLda/pXV4UIDAm
RSdW40KGkXq1OCqbvDjd43UiGpBWzamvyyP3QpICPYTIb4KG8kxozm/xENzRnsxT
MmSjQc/5Iy8LwkNUeVRgfmQnkvdUlHMBA2m8hq99ZhBcGKpOd6up4R8Hj/g/TYeh
zyTKs8xaxsgn09rY7+WjVwHmkjYmjaevIB+U0Z8MRsUGeRc9jtEA+XX7DEUXIyEY
dEIQ3RPh1SxmKndWEnhxsBrfJILpJh+75wGAw/G2eNlQUDRSmVmvR+Ez4qQey0N6
MD50xdWon7t2ypDcXF7BX1K17GXO7dvD2z1vqOWp5A+2RQJUzka4LNoX1giejwuY
UAbI6CdKSdszpaf2VtTyMlkHD+qXnGkZKchJg5FRaROXzvwevdIZ4Cc6RcTpM1Dd
75sWFXQ4CDJVqwkjEU+iBf/i6IHnAPhWdh8nvTjOj66qwPBvWwylFYhDgVQdRxtt
ivZhowQ5D08OHVE86mlfFvAjIpoGcHQ/uR9nX1Or3UI1zRatcC/KVVSpO9S4PPyx
QoFsU2YVBE0kP9yciWlLcITSPC8dbIYO5jIpAqR5S1Gpz+hDkLU0wvvbZRycG0Ee
HU7eKeW46KrvENGlkFagWQULM/mU3nUcSdSltjRJv+Otli2wNDB3KTM1bHxBNGWm
ugMO9uFklz5UFEpg4laqysly4Z+g5kXluPB4+FOkpjf44tv1Sm2TtQOpqt+Yu1de
GJOMNw/NrGSFaxIBzTpVXwJRYxdtTPkAUw4R5vk49F8vQn40dIJCOM9k1cbribxM
Kuw6KlTajl64wqenQQQRf2dXRSdmXDAQu5T0g2sdr5Qh0OZYHmL7R7Wpni90+PNU
tUgYxpHf1qxzJo7t2e0hkJl2rykvsgN/SC0Z/EmhJlqgh0idd47e8B8KyJw1XgL3
MprYgIvUo04CRBfd1DBf/KUMAw11pF3Sqq7s4sBxmHBssYfmk2wvCgo4GJJEUw87
eOFWcxmMGyFPrWJE91VYqdBKoLAzc0QLcaCsIVci9uWGi9weOTHwPJO3VrKkehsu
o5d6N4ywAJ/TMbGVlV//XJ+AsqYWRmFXhQ4DLxPIg1IFbx2Ae6G4MyS5N5ZGpC5u
P4pEIkOolvYg6neIQHrnZqLwZlqtrUbBEHjjY1WLwuULr9qy38FEu0vjERBlZZcX
zKPBWAe26HCjZWJ3+xSfeWtpABZAagjigK+gKFmNcEJ5ulf2FSYiPMrtzuDeZBQe
tIa1IqCHxp/Wxpnwr9wRiRsG2OU7NMXdqdJEp0Cco1R3gcBjznT8FmdK8jqj0E/V
R9YJroM9YlVQ/tX4IlwlbkHkcJyqUS5k/MOB/eujhaWTlC0NDmba5BcY6QcF8QNS
DvAe8n8pSKJv9r/FUZS2AWvIL4RpmwwjD48OGTrkZK0dOWETZlRarLdTSEZMeLw5
hecNReq4Rl+36Bh6Sqw4SakhiVvyeqGylhzQBhhrcVebzq6SBbut3YuJ7/IlVr3+
UhEScz7EPTT/5Vm4yuLFZTaFRF3JSmXwWfMIqLsPZFWgMm+795NXEhEkzsMTeOYa
HeaB1LyM7NU7ppMrWHRQk3DsFLsT3uW0v7FQ0gQvr87r0fu4Ohad8sR3M4T33Mv6
S8+wGz6EAUJ/qFgT2i0lyCtlS1zdmfjBesqpvGWZBw4n8TQTMdfhu+GiCPLc56RQ
/TKqOnvcUTuLovuNvzFJoOXoOOo17N2woRBjfd1wiTbPq6q7MfSQY4VqeuHhSpMw
UQ8Tu90f4Y7Cf58LTtnKoi4RX6d0TYd6QbVd842nqvw2uU7+D0VAVR7P+29q/tGk
elS4L6m3o6yf0Fvl9uxPap+hUhGZL6tJiKNis5rMXW47KlwYcr4kbTiGjycrB4tX
79Rfjt6plk0/EtIw1cUnrwnkgMFGBrcJYrTWVTJpWrFUxoe3RsRJSnovD50f3/Hg
p901Oc/iCGQ1aKAQ6aTJ7O3q9ng0RqcnK4/jhnTR1bWfNyD5pv7sz5lRnGrmUHYt
1BmF8WD6Jsvjc1fxW9gYVLUFn4KJDiKHqMWFDjBX9G5RUnT+e624MabTnOPkglqf
3DKZQyQioOpU+PSZyGnz+/ZO8WKXEUdtA/po3Zvp4PUV6nMMZv3z5ihaKAjuMNsT
Fs+i2ht+fiXiQ5WZ1rgvsG1IDoMfIdOw0Lq3Bp0ytEReI9PeQh1aKG16UN1UcaGi
2LT7UYTCO/yGqaKUeYYEQq6fKmvQ/tiGUjxsxCkPCVn8qYijTTB+Tws8qLfiZTQc
1rw9W7efoS/smPp9sPjMx+Ho6FNXmsAiyCIGWu8mwrlt1ZSowLhDGsYFk6VEMSo2
ywppKqBLwB9ETgJjWjNGhzjl1/nkTENbr8lOtydQyCCGxFIwt5sY2a3TeiTlrygK
uFvW91egrGlH/tRKGtsSD8ybAr714jzR5vXPX8JaSa8LcH/sYSvwTuBgiBKqiEOF
SK3QUUuJEPmkwY29hN7R7EkhmVE1b4E57zRWXG83ZfZMTn6/jfu8UfATHmrYxYxz
m0HO0uqPbLlz7Rji6nkSw0qKwL8LxURuN7hjJX9Oeaf8iz9a6UK2ZTTlW9eBtHal
RIKggojP76L7bduMWBXbzpHh5DUkDZ1/4mQW3/AYl2D30yEm5tt+T9228WXfc8+l
ZCQptuOb1gXNCbv90WJ8D8zEnCZps7n3jNYW65j9Uv07pZZYCl0RzHBUGrvV+DCV
9BvPRz+gMYWY9Jr8nuU4h+ORyxbK46Z/5t9PO20sb0bWf1es1x1V0G8uL3dkqA0y
LoxUC8aA+VaP9kmGaVYwBsXhJaShxP7n96f5Umh7D6TN3ix+l5cZMcAQic5XofRx
oKibsOx3Ks2oWTb0hqbJuSUjUldSpn+2kV4J6CwkD/95cB5hZWR2bRRmFyoyEq/C
LPbiRgF+pQv+o3gjgqX5itGt9BcIj+wWWiRPqU4RrVMTMJpneb1HDoPwcqUGtap5
DgPeQqPFkCfIY4+ijTNrTVPBJ3qMutvqYONU++Mf1zvZBDDFd9sAxHQzttsGu3PI
H3ZXTEpso9AFbpGzNowoZLH6uvTlg5INi60HRjqvAB7VGiKdlLxZ/lIAd7c96FPZ
a9dUNlAz/qabTlwNAY28Z9NKNG8Ywpf9HT641v0FQE4/py8WfdZWHan1nZEloZsH
qc2MT7HIFIXP96u2I4gLSXrd4MQto7m1t3sx7rKD09xlHJwHPzBPTZaaFwr91Ugm
Aq3Y21O1CKZ+y9zpchVhfcFGrzmMCDCESkhp2zgRJ+7D4tGWIuTqIPtVKRtR8SwM
qdmezbrzjezAIRYXIS3gm1R6vKmqkK+6/6ervz0S4oYZj31dt2iLoJOkY33uckPv
5yS5olFx0FNJomR24uyCGnh0yRZxNC2mNtWxibBDxFRlotBZsI3gpMe9k1h8k/PF
+O+c+NmH+m0aQebAVx6qY8Ng60K93UJ2lFFqQG1gwmx48giYGITsaRE4A4Mb0dvl
NiwGNGcN6l84nC/U6SSk9NG574icyND5wBaSMwx0lI3iYKu44xLlEJyB/xzA32Tz
qFdPOl7mNF3gm/yz73cXubitXrXYanPXYza4iaoC2TXVcsFeGrxDriM3HhAGEdtk
q+HSpcyzyZDjs0dMP5M6V3bdTCNzWikAUJ7eU+YWXg1X2Y3bx6x0bBU0yNZGNACQ
cSV3K1PS7bTHabY19k3TfGyFIuJMVDLzsjhliFkhZMnHqAB+6uBnklKFsY4K1Gcz
Hn4Tyu0zXO6FwtxBHFTHVTBB5BRGD/jvtDfqLRFQFu3WdXW4GYGA+r5SOe3lQf0N
D9CV6WjGwdCVyLpXxVgMsAJvPAt90GynV5wTwIAHmR5bH1pfGbPlJevP+TqrVjX1
sWFHp4fmdv87C21tbvJdLZ7HSzc61d6PzuusvYVqc+E2gq962oY0OYY9uXiMvmg6
9RAFJXbfPyDHbqFcW4a2ipM3Y5SFO9W8+RceQ0RB5ocIop9OOouTfCBkNv/anFhq
xAMwctq6pvte/vvO7DpM7+sz/dRKBhqUd+mPINBz8/gq2//38Zk/PkJSD+EecXc1
CrzLhODbMXQLfOVaJVBMozk1tQA3tBTxyLrvQ0Tun92/fHpCqsUxnY3y4K2r7UHR
ezrE5y1La8wqQ39g9SmAkSsFVWYA1F99oPZm80LvyD/rcndDR7+KlIR/p3/W26oU
m7USsyOS/QBBoq4ED/CmF0WeX6e/e75qN00FpJ707vTYFoOjVdjZkLwO8dv9WaCE
zrpTdR5AMyFEQ2unMyK9lDNz9d0GhZ8wUcXBXYUSJYC+mcY9eoyMBkKkLThfREfU
Q+eBFZvAGGvJ0/dL09S0J/FLo6rTQqzfCgtxWL6oA8QsjAfsZVOqBadqdI0dwN82
xMDEVbPLxNR9ZoMFOHVfMv8wS7bV3QlHHPz1aAqpNjiJ8hGr6gqdGofJwVTGNgT4
lo7M28pnLVs7vx6jrzeuWNXFFWNH/2Cb8q8RBfJqvNT7GxwA4czKkdE8LzQPdA8l
4fg6pmw0Qp1XGvbRphyRFDMKlqnfiILMVWRrVlG+LsYtz9iSSDXZ4Ufl2EfqWuSr
9kFJEV5sb8frAzfiDRD0Q0+/gA+8RmyrA5NampSiJagwr0Zo8T7Ual7S1V+s3v+d
EEw7j4ua+JghrnNHxFfdJgOAKsXN3XBuVcskrf9YaKLfriyTfS7KJPfpR7WdIDfO
xJpasvJsK7zVZtLrzYCM8MGNjFTAY8eLoQF642sdkAtRGzam311Vs/3cQhno6Cfy
lopF/lFOc3dOuXn8XKqLfh2oGQKoTCZVDBFee9Wu/pGOVKmef3AoMZp/FbTqK4qx
HnfwHE7Ltt18R5AY4i45nXjm2SzE2YRvFk29/eWWPF6LQ4Ram4p/r0CyMuVzgSDa
dd18dPRr9qjeoy4r7dthhDMFHuDivDRsGfC6ZI3WTQkLuNbZJvXwK8Sp6VtNEEHr
OzmTCA/AUxreT38tPW6qTF/qOnTIqfC91Rx+GjpOH7MKXQ2X87hOL7S+THlyZujK
dIJMKoT3e9ynyXynuMAwqDd2gOKywy6nPM97O8ctH70QCkI8avOliM8+deaQpQ2A
OPHf63KIvQ2E59v1nIYalQPtnuCLBZ1OyBqhrF3GNv56Ed2AYki+D6MPFApKb6Ad
b5OnVa6WAqXE9U7wKaXJiXo6TUpcilF6O9J37FljH5V3GeIwYAN9lOrtxBMoIRj4
urwQM1Te60DXAWcc/pL3P+Qq5Os9K4bjvhF1sSxwIhw5fwRj8umXGk+D/3y4gJbU
Wk9mTeicPvq9gprz7X+vFrGmK275EnHECcJX1hoomTEiTuHWkzxG2zpITrcA56B2
NwzKbOmp6ZWO7df8Xsm1mS+B0Pepy+1queGLYPmcQUJo9a22H2D1H+8hOR9Rx9Z8
EasLPIndJgpIXZuOcB2YTQ7nIUWBc68N4wjmqkUN9Sl4LUBT2J7BvkhZ+nNnsS70
TsFaThi0rIYHSyEr0+Q13pfV8sr4+CqrTbqlACPsQqTxUjFVbq8WD3lFcZ7z4uij
2OiurgET3nAzn03VaNKIPtmHMSWTS9qKFyj4WOErGl15mpv2IretsyCoieBJHjuZ
b+331mqzVzdKmpeekvkiJH1p/YF/DjQGjIsUBfjWzxlGj3bMk+hVEDqVtyJ2SJ80
R4U+OeCQriBno4Pu0n1Gtg4Qn6304PZIJiSnKgMnAXOGLrvydA0SCPyNwEAWqxZy
FqXWR1/GDlMQ9LBOwTrvrrJP7AP5CRsreP2HAgT+6rEsP1NmCsrh5XBHAPncYgur
nM2SFjEUCDBnmDSr4fT1M2YXe9d4R8+FwcoVMHe6xOZ5afXHuFwZGGQWF8CrKkKZ
ObzuTaIeTh1aid+gvH0YE8h5mFkffHnyr87N3Dy8KjXOeJMNQcXFQCwSYOQIKGlb
/7BmbGzV1sIkdPA/2XEA2L6pdFtoZza83+0Ki2h9ATI4carbrLypAmk1NAGyjQjj
zFGwn4jwoulSNJFkrCnM9TWUFgcQvYDo5i2DttVOZJSYuBdRiCvB09CTcCdb8w8b
0z4Nef7+Se0iDgyd5KcLKbAmL8i+VUOy47rKvAzVrkgPbLRID4evSXMQHnIh7vOq
YgypS3kG6+oRER/uub5z7dqTxlAzuQvT6ZtHDTTo3o/Z4g95ZGLl3bSZ1tZ/C6lz
847TDXdmV7bplNvKRPJiA+OVOAn4oIhTu8SIurDRowKx8LeBUM6eQasUrMeGOOZj
cC2LTDlZzY0kCQGAr+sdb69a7LGz1FkaiskZ+9EHN7BQdlYoAPm+L7OHm+t7fKrp
CaWARwuZnOCiV3Yg8r1jNZZ+PIHlDGW3XOn3Or2kWtIAbI3EceXbo39NV5iFsKMY
mBzz2HIjUoqv2WxQdczA6fehyXLAIU6AyNHOSvZ5k1UxCKa9uX1cBaBGhPEJmmC/
4Yvp9cq1KSvKNgSOOhm0qWyNQ1Oh48eu1J4VxdsLRl0uzhj76mmF68LzEsUHyCOq
nHjC/Uxh+A7GdJwq83ci035JBjiQJD7rlekhyxpahGNjvFGSBsznmtl7uEXGPiH3
0pa3Y+Uhh/o3dRnkHtDYx1wSu8ma2Bemeax5LUtbutQF0BXJUBtpCXZFg/lSCumt
7e+s6ARNrWbXj4WRZQFqEGwD4SRk6N7UFBpT0xBRezgKvnRyzKq8W1VaibtJX+9g
yzDoi6yUB99PxTuy5EokY8uoaoZmjiC3e5S8rlSD8Nd9VNpZuZFnnIdOSZG1FKMj
x3sjAFAxO2YbArLvt/VkHKo7HLWi+H5mJv/1xEuihcAo5YKMonUSzQqvFdF1lkFV
en2Tf6iWkErwD2120Q73u4FEPYis/f3xMba5jtqM7vdEAgzPJ4fkHjHkIeGran5j
pVFIoGXurO7HXOQ26iiy5zwZ0gCs0tNNo0y5jv8lziK4z9XxfQNAKMnC4X17Y2d/
VfSLGq4bb0LydP2c4bZgsWWjZ9S3ddDVnXsLGSXEaRzGX3AcB5Bn0s8Vn/s59oPU
/0BuuKQmF8mtfglneujNG9jOxr4l8pNukok30CFN8wAo7BSHODHtxy+QViUMp9Dz
2+ksPLeSDRC/oKg3yVuv3t7gBV9UhNwYcXq2igd6xF0dQ0eh918/22PL31Xt5tOf
cEBsM95pBVzPPho3dlh6Uppw9BqDNMdvncd0PHrjb8JrGuDwtwR/eRjMf+l9y/hY
o7L7eHhiSVqVBF9uuO8aCQ2E7PvgvQ5LSYSvF3Zy04PTMfjxICROMKVnaWD9P5bl
AloRgadWaRLiuXMCJJWsZ3X9qZ/Be2kCaZUKGFTrMSHdbzI3NZ/ABXKt89g8Kctv
Q2FXuSif81zIt+QvoRB/nXwuyJd7JkNaF71yj5iNKTbMzi/0ukYXOghwYbV/mdRw
PPrur5K2ZFI9JypM+BlpV0NxHzNNgkQLdfiZdB6bE5lI+hTIrVA33VR2yp7duFW7
nlqnKQPoPA9tI3/3Up9akDc7CNfNMhncQDAMbfW8Sde/wM9DhmlIYlQb7C5IoTPU
14DLvhr1i948ZdXunUsV2icLZu7wUlSf9HAj6dVnFqAHMvwqzU8gBX5lR4US1yNF
/6QZudO0r6dR1g5CPKh0fkPJ9CXeEubsDxKcE+sy89SYfhpmp2my+L9GVg88e6zM
sz9VleQDU+hP4RYhXqDF2Da/GauGZJGMuDKuQzHDEigArbhtrlUmxc96fh4ZuI0D
738HjOth3TKxezx45Z8L2MdNKGZPubolhVVvaInRqRbsWwYxGU28GwjPLdiKNfzd
FbRTxMusqyat5zHVK395Yh7gyoCcw0XkcxKybNsnVWSHD1cpgY22abEv9RIcwCuP
SYb6JwCzLbasy6cdHnUqRFsQ15giQ6d//CUFcsNqUBReZwrVUb8UWGBCSopDAbE0
RVmzL3d5ToX4dfXJRkr9MdLgPyrKFEumU0fhYectwBV2zTE8PC0+5fbeksmcOSjV
VlVKvVCi4OA8H0wVbgueNwbPBqPXB1NwE7W/cne77Ivii+bifO9ttnpruVHiYJOm
qMKBGmLd1L6O7MXB+rRIYDOSkFLqiwnGn+PyG72/zGZPioN2SSvBUTGr/Ns8qzAD
ZYQcE6zNhdw7b+gryliioGCDzJlc8drOEsWZQSHz8Jcll0mIjYAWS4wr3yoBNoXE
5mk6OWUO4OMDkKLcHPMcGvXeyo+WMe1owICtedjBmjyilK/jXajMt2N2cdK6htS7
Bcpreywqf2XTandha3IDeE5D423OxDB/FX8KkxUgqORRjQmKUE0/ccQ6bQeACAAF
Xbn7l5+jFk2eKvJLkURVYADHcEGb9ASZus3NflwFVNIlqFjppT8yKPTpdrPBHdnG
fFd95KKDJMdZBHl6r4uDzWRPY08do8zeaSqBMUTKQgZpSRM7OpD4864OxzrFKGn3
WaS5h4KHHSuAcx5dT2uhB3Bi8IkPDnmDj1OOVcfVeTwO7i5JIWSvhDz5orxTEZZv
ToXfOrVnVyMzkq3MSrptXtm22zmBqRxkyGNoPCWnb7X0XjAtVhH2tV/S5dx2n6Vg
KBCWyDZKXZRj86zMZ9SSz7uRc4b7aMQ4pnUx7FU6wwqWYO1nQ/Dth223tKr6m0nw
tz6141LGTnzoOYMDukjvKqyIsMbHN5GUkntQOpxo8qHdr0Kn5o8GXnuqLlopAYxv
GOCC6pgl6zjNXRdohjRertitIAuCePFmxUUtCtciCTZurD+3Q4jLf+iY7z8p41jv
P5FkhfkObd6Lw66ueS8rMlyyZ2KConHDT19wOxkAwaQrccYLynQkHue0xDjCGIu6
O61oPlYq3qCl9lH3D4bPOjgn4k2lTjkt8TmTaYi66J+MQ9ehKt7dqTAEa2w3CqAs
lw5KnKpfhPnYmV5Qxfn84qYpmGk2P7muwmpeMsZNR+XJ5SWyVFi7XWoxPtcWSL+A
luXPoi48C3QvcJsSDh1x5jRI5hgpEBO0Js4adf5RVyF01AEiLfE3N+yg5YZhyWlT
dH/nFUqfy84294r5N8zt4CSvd6SUteqm0KbcEWAUz+F+eMur6EbCVipFi0xiBKng
BExKCgAN4D3YP/D10JoSo+eb7Upi68QKTnVAaAZG1m7TQcj6uHVHB2skWed8P+Cx
pzdmELFuKJHkXxIyGgA1odWGlNYBbRMkO7+CxCU4wnMCDmke0cL/uTVhUVS/uHBf
PerMB5vPdnAdFOqVCFjWlQA6fdF61Iu0BUcp68DEIOUJfEe8F+uJsO/FjRkLnUSC
qHkn0tjkFdQZHvNgM4kWch47LsXLe9y29R1xODbDZ74OmN1COUmhj/uE3mZ1IvAr
HNFDRBHZcGkvlqKVU9hS91ryM5hT0D6H0Af7pLJCQgzDE+RtuP7c9cx7Ot6tJSyb
DFIFphHXDUliMHdW2t08jhuA4nWHKKsXHOu1i99OFmgiHeuCQlAlOuH/4pfNLz+4
TEzjChZ2eivKp6eMgk5du4yAQ8jTNxze3a9nwbT3e6a4EyIvShiyEhmg3qF12P1C
sCvHQVoq//a1Bw71rmGnSpgVqQ1kFDkAPNx7V/xtxJj09MhIFJuUjGkINvUsUFWH
0wp55TJ2WZLWZX+U6yM/byz8hd7zGG0t7mtr5CgRNHRfcn4ew8JZTBCsrMeJCwU0
+jvFSK6DFQlCgFbzRbVAlcwiu8AKv2CzwM3n+KlOR55Edx9QJB2px8sCt4eOF2xd
hZazZvOx0IHUPqH5hnfo3/ZP0ZDnSyXIDbjYmXxcAlm1LLsNstQLLEMwQHsG2ZiE
w3eFTrchQSp/Wpwl+LNaCk48hx3nhqfVEki8qDnmmZjD7PX1WI0si1At9sWisX1t
arexbdV9HEd8jRQbUhQc4sgNPDVFmmy4LhcuxeD2zgnMFJ3vkP3omxPs8pncXIJP
OXEcgvU059W6QjNrCA0nYmCjYl0ZPgTQ71EckzqHKV4TQ1ftBl8j8pUpnopyDmPy
DHvJtyvBEi9mrazm1KKuRANzg0OK0AKBSFTPwVuZ3t4oOUbaGniOtb3n+norL58+
rFbeSLi67C7KY49bqOjeIrOgqTpYU2OX/+JWd9SSEeWE/P07ZkXjoAgO/A7wWf0v
Vn/w8LpZzBNry4I7G7dyrfiUJJmxnftRnzXeS/vSqzBwNywVtncfwlXYjuiuzdGW
tbk5/DOOKAuyQFrFhkBUDnu1LCyKFcrz42WQ1/+jpB5NBCtQa9OUfJzoL2Uu/jH1
ScB5pXoQn68Z22CbOVuwZoJ1S516khO6lCX53rf9J41qzAm6+4sQUKwJ7fprd2tY
18Ub9YzpvVTMehqekvh7KIzddDCVC54T3H0iHvV1t39BnmIzqUya5tGyhpHWeK17
MM7rrtKiej8HSqYEAckCGhLO7nLxuRo84pd9d1eVfram0nWBn+/kVwZIvA+qG+C4
GbOsQq2sxb61eVGYBMtTz0UAzMaBFjdDB8+zxSp4fDG+R9RnOzHypyu4yXCrneOz
pUaUwmEOFlsS02bLb0MN9ke6q02Y9+BDIdl4O1AeBW0N+d+weB68PV7cGdPQamaQ
5V04da5dioeKwK9wnccl7nGaVaQ5D/GmAl3w8fhUwsivRxe013utULiY1Ieuv2mN
mGEL8S0VURcVyPQWu1wM+xCj3GAuwMpTyLISdBoV6nB09VT6D1qd+ruxwMUb1w42
oDrX3P4BJhtRgiYo9sSivrAPSOn1ZPIcSQBo7TLdqFangAGLenj7xqb8xeD9jqg3
n+zbsxhy3g43E0J4gFM9jDzha1bSHT99cuyEeyQVjn8JtWKremjx+0nX8FVlPuUm
P8I9hDODGUNewKNPb5HwRWyjUk4KjzXRG4Tm03wQoLNAa7tpwuZU7pjtXlGg353Y
Fod26aRGa1fYzpgZ+/yRe4cmcBIGnPVLX7FaFh68DjcZUZ9R5wYfJYnFDSm7dJE1
4oB3/8ISxLSaGdgtdLMWohhsM5Wx0KR+db74irCeiq0BJKok859bY8WUIW1Hap9E
3DvtGxxdJ9MbHONB6U+d89SiyckR2IfBK+Sj0cf2VqL78mwMeMZZ/i65Yj8n3kdg
HWhlQbyi9x/pY3RiHgVoqI1uPJq5Q0elhxKGQlJLAHMzcyoeMfqFTlbcQeiMds0l
3zDlFOG1yorInA264yc29oys0jIrYNitnX/xIZ8pCJOvVBCx1PjU+JDQamnsgudP
jNEi4Lr4qnG7Md7F9NpehPTgESevUZV4Pna4/JlIfF2Qj0qqxI5R++kXordb+VKy
IndWWZThKIws15DH4MqyG81jr/xypcXAcaaDzOp9Mh+ehUT9FNK++iBThUqeDkg2
qlqJzs3qLVbOmyQVXTUTQriGdO+Gk+4HcMtSKLuBNxt93bjtCG960HwqG0f8sTNK
xzsWjj+RJT4WZzh1Hom675/B5Ub1uQT4eKZMcxqBAc3AvDkaId1nF/TfjalEUfTf
/z6MtCXNjiScbKPRfkbNnJqhZlRIo0RaC7Z1Fmy1kuVKPwd0HmHy8mQR4G8hWQed
uIqyhwbDXqZ5ApQ3sk9ve/gSyl04n5Vz+ckzqbLSrwqKdN34Kz+mcLQ0MFoaqF49
8MRHS8FgxJkhlPfYu8zr8H3Ur4s1eTZnJ5+PzMC+H4CHfPsR0ON7vn02NFW5LG8q
fx5R5S7LE1Bq3FN07ogblU/zPKsLMqxAMQsjTFMlE3fZTCcke5aIW99IxD3IQ+M8
io0HgJ0FiIatStrm//rzCMrE9tmzpGlrsSUnjNxhlyT3/aeNTdyn64pGFKkq5Zo4
q057s6AmBKBiXsaSBYIPaBEidceX9zSp3yq4SYTrgzb1FJMIrOlHuYscpm1Xd9qG
HAsrvbbPGQZX2QWmIJ6LvtsG79TGDdIVHz1FwR8r3vUvtn4gEs3eboQTBmGjFMpx
cO438QUggecPm7qBMs4tRNykBT65Gg+2x59wxmHYeYxigTjlmjeNEevbBUhjgKCo
X8pikWSKUjIdj7BP482nBp9bmJxS3NtQiAelPK11oSvuPJTe8wppmCDWJa2ziKU6
64aY7P2+Ip+mW7rzNGs4iYXOb+f9Mg+aCpfG4SWTdTWOrT3HgoFKiQuUnAD539B2
601LinWX1imbW7ZoFp+8YNWdreP80apfJPK/zikouOD+w2sxXhp41IT7hzoBBXC8
aTczD7lFsvPazT5PcDIu93Kh1MabyMNEtcKP1suB2CibvGsVeJltGDfo+MBZausc
oxN5DvqKsRJN1cv3vzgbqacN/hMJDygZkj9wZ7Id1IMuBl10uOMcmX2wktyLWwGu
Vr5FTvCJuR44xnDE1FIC8iZf+PB+xfhyqO2Ep6AFKjAkSzVtjNHKuQseZf3/PRpR
bI9ImcFbiyLz5OLqeOJ3Nsq6edXr4mYiFDOlR0Z5NQJJlz4kBPVGkq0PCOEK6OmW
U1TinzdMMPWC8VtPILYI4sVLrqvf2ZJDDjKqTOkkCGEXxxTudMDJCfQFIApqiX/+
B4WvQY0679g8/epDVZirZRavTjj8189O7fU2ylfcqUC9pwWGYVuPPyJlUU9i/cLM
J/hFb1rrdoTsbgU1Q6hIiCkQwIeyrGlTyJpO/6zTEUKnaoWpXWL9Eh1Gt0oUmjnt
NNMrm19kKLM5NK5NrXfVvVcCyKm2PFmjkxTkC8wVshNRhMdhozqz7UM6LiFOQM5Y
NcFj933TAnIhhKrMOw6w70E0m6ycEGDLjZYYRa9Uo0NnAGNcIsdfGVh5ePHUR4fo
gf6TbWYtCZN7Bki9ax5rUf1YV3K+sK0ra3PBrqJaG1Ur3LoIaNnEjlQGBmi7fe9k
1qRXbGrbOIAFL9lXBVXUjZkrEhbkiSxQcMtIvGkBLsBQrvQ4FnBlOnesuhx48Sgq
6809DrxHmsv6u02EESW0RU1Q2pkG5eoicYt8X3+1gDXHhxStFudXf2NWFy3OIVVw
4C6qmY3wLiJt4oft8kqMELgTSpJj1lCHLwP+mg0ZtrHHx+dqnNZBMhCUDovnVqpB
8IFGqvz+6uW5X1oxI6ltbbG3csqmQUkI5CuIi97tPvaBLzO4VKzKaFAKYtc7l0sU
Q+PGYpLpwd2mYG+Cofmv6yk+8A4KExhoxLGb86ITn+qnVJogdbfq0bJVOvqe/tIw
nRNLI5uDkhoaESUqCSr9wATv82POpRhj2ZRsWj+STkooNs5W3ntxPDG2YdVt68Cu
j5fufFQkd0OW3/COSYTq3+1EIIz3y7N6uY1Vu2DiWLeejy/5HTeetAJDL3H9Kutx
VV2qKtLw9yTUoLvI5l579ELeb3A3OH5/0klrwXiVCyh7PjpXLornfsokODJnKQnl
wkH6zKAGJG5qt8V6avv5fhuB2eBKdRDUM8W3iliAoc3pJv4cF2hUwCGTvDZhnVz7
07c9bWW55xRxMvOSJKOsCp3zVI+HLnBQ3Y7r6wzcFn6C5FlcI4eRKb+BBZSb9Xa+
KsAuV6EZx79F7bNvPF/p7B170P2UYL6DjTTnck4Yo1ZkpK1+tzUTiYg5WOuL7r2o
rc6HGvJwcVX3hpuvFB+IERB8gnD2NecmZeG0wTm+rbpDe3qLkZLkEEIYUKuOiyVT
iJyYJOsLZTGatndAt8eys5/cDsDrJYeXpgIi2ifkqSxIIUmUcqLdSfLQ3UBO/yxS
oQw0IR4DhOH8TOwIAYLu6oHWpVkFgsZCJ8TgV8zYXtz4vEcVCiT6x+rRBlY0Kqbx
vLcOUgFW6fx1oih+MmHyR3xA6Bk8AGUQXOpybpGZ3nTmYP6rCTr/kVhurrLb51/K
XyrUIYbVbBfMtPNbVoydHa/CPlkxluBYooX27ObyR6XJgIs6VTlwmZS7yVmdt1YR
yeQIOekF3Dcpo/bAYKCt5SbvkodHJ9gWprANvs6aflgofKCKnQSKMvhTFnG9KsqM
RzVTa+EqEiCUWBnVqgjxbFvwvseRNUd6b7xCaISc/Mn7QoHqIFW86C/vyaJoe6Dx
bIdp4NVym6ni9WDswrSVduZgKRq1Ea670bJaoqEcozpLIcnZSAt9bR8Bd46qifws
ESXH1/5Jmeb+IpBmxOWbwqbz8GF9mHEGbRr3PL5VJfvhoBOvlM9ZAoI3AycxrOph
xdNERxXjBS180nNVol2Te/rb2XZKMnBSyHDCC+R/GexrEz/0t+vAwpgpxsBRCKd7
wZk/UjXKL0jyVtcJS1/CKtLH+6IXFKojb1gN1UH5RKyI3Dh7UJoEE2uCk4uHqVxY
4wcD9cfi3VKDCXkOvXUW9vjvAuKVB0p96paM/bjcRAnVYFvPEv/VMMaUvrnJlhLB
qr/E8fWe2qa9jztpxeRkpQtqUZS/qmRTL1bx30qH+FfzYI5rC1wBHEZ6m2Wz19Qu
Yw1en2DpK58M4PKKwescpSt0Mg3flWo2+uB1sWNEn6NEMT3WsYUQs6x5UVBMVKmr
Msanwdf4DEEnyQ1F4RwvZZ4hEFV9ORoCWx0AU/m5NKw6Chi0SBSLQCxhkePALqLF
TbxpXKGWjZsE4nY0fHedugx4uGynTXuqZ+pK+hffF90Dnc/QcfbvZlZ9mybCC05a
dfD8HN7ADye7PtD+sPyM1Cre6wlU7HLMXGbRBg9zzByA1saLX48sVvUhRTsCDUm8
5dQvaw23TpiZ+I75osUfzrwrcXVrRcp7gpQaxXRGRryh5p73QRiANqGT8Kt0sNBr
xiFCZk7fe7VH03F5iS48hNlHqrr3D00354QhRZU/3N77OyTTSkOtPAjfc2kLNbov
umduzfZvXgHjcKAxvmrVLsc2fBupLHtJonzIj9IVCTVypvsGz9oN2qnXw0uL3uTt
sQ7mH6V8LOsmLUlOysJGYi01f8whOOiWEKZH5YNaR0Oo0DFkW1hZszt1KWkh5R44
dY+HjFrFpay9edPlzAAwysedE7D/NZTChl5JFIFKFc3TZKA3QfUrKdY5HeoiplN7
CK3CO+sgvFUwgAr2ZQv8n3rjNP/VPUUbj/kKkYGFutIfLWI1knx4fdwnJ62RsXlH
nkm7sqFefxd261aBLoVMkppm+0LHZB2Tk3XRkXPh2WluF/OAYRD56Pp/aORuNeZY
/Bnruf8s+23QvTbhLrwK2KtkIyIwEPrDXSyuOi6QnzNGopcp9j6ntKTCUQTujl8D
72NVP32ruh8cQukJ55IXhB9PwNdZsaF4kOV/I73H/RShx1QYfRomuZaY0fBpkG/e
g3TQTAhEn3qjKEyzOtzeyM9BWBZ7zpwWkqQqZqsxXfLGL+RALgxfX5ijEPsTKc4t
+HmFoTMaw7FmD8jeNwxwqgpRz4rp6mlmQvhQpXUiSSP7tNaER96OlLRZ4B0s7p9R
ypI5hEgBH6G6iWi/q3qI6+naSUn9iMvm5MieLakRlolyaapTNswFS58F0vll8gek
LIFzB2FaXi6CETgJyOwaw9o6XZRoiF101DsBTpmCjI9A6my1i6j1T6mGmxRRSA2d
LfYOxJIPD6M/XEh0K5Eud7Lom6raUH558WXotSFhyvy42cGzaarUerOBQVhuKIT9
zHuV71Ehis5exp4TltIwQdClQfbYRTd0Zr+j4bRGl908RU+sDLOwFxaXBbW7Q1eA
F+xplKa3lMf3Pn2kz41x0Lm1GbHApibD0OEji+tb7cfuV+toA/IURSovaG3VMXHH
mejr0vQY6UjyjWohGwJv84v2t9l/MKOcbGrmE0M7IzQ0HuApwb9qXJ7iqmqRHvvf
D57rtq1DNr3L0uPMKTTDrN8Uidgfl7YYnXLNrr8LcBL5Ka7GTNjv37qkROMnmPKR
zCI44Xn+KhXVop3DrOCOSgR3DkbrTe/H8LEJeIlJqDRdgyYfSUHZqGj73No5bgG3
csBSxSqwl472PVMgaJelXdrs7Ypbm36O8vKyCp6NiyyQqWzwL3BKe9ZEQCGmqDfj
gH3OlCJjIO8Qvdq01tv+kb8hPPrytxxj9rkc8hD2SC8on1Vw+lw1dZZ36ycxGOMN
8AT9Ta7gBqV45pRVnxIor8OR+tEhmciYzymJro9odBXHZdm479u1AjuST++dTg5K
iaA7rGS63fK6CfdI4UrlerPGXEtFWRYzUYZ5YJN2V0te24m/NXb5Va8OcBi79cWk
JpivOP8PH0pNuuVQZsWiqvTRpqtEIrL13cg7uY39DmuIsFMPY0NBFFuYnqFUZDAa
fQsQjJZx3iq6/16GYto2UrUnJwqeFKQImYcbe7R8a9ALYrPDyLgaKgqx8RKYD5kp
1j+12LKGBu3w/NrazcmbaE/PymxdpuSmJ8pBQ9R630WAooj+XZWJQWJVzivVjplW
kf9q3am3JJGtQUsHCcAnOEdvfJQcLmX2M8fO8dtDfCcMsEj+Ipvl9Od+vhG6nwLw
QPLAPaCfiT2q+KEg2ina2isozf/mqrKOG/CPqfTL7wG2643AkF5nQmhPEvwQuZWz
/j53xdQdH4YEqf9RjZAolxnFqVnyGrlziX/bRAMLzIK8PnoiWJU3VlW6m0zAZc5B
M3LstkmbUsbyBqIN817gQrHQHzwqgM0m+624Zs7Zan4DHSHFIQloCzi6q2EiijIm
p5uiAd1hXFSqlHj6ELQZKc2JeYxZO7m/cZuCxJgv5qPvP0g/ZWrFhfX8IVgQOib7
obKg3FUSFGRz2A9DJqXoEO1uRWTujZhp/UI9MKSJl0ahr2NMN3o/U50x/4J2tKge
jPEI/V8OcCNHtj3kA4fF851swTqoXU4AekWNf2DdrmfBSPT4HPR4k9EeTZJFDyR7
cGwVBCAD50+UK7z1jxg35tVuTpasBYgJr1YnBZG6KZDNOkmRGroy4rPs9vURb5yR
/Te4ufAe9NFc4OgeZp/wOcpRKJlynKNFqkWZk4AREsB4dJ60z2hLv8BZK1j9ttG3
5vJcnRVSVpZFi9rGstPuoil83CauImpYOjVMi+D82FkjbC06ztQosyy3fhWYPaNk
3clGpIVQFoJ4xAyeiW0TEBU5LWtpAATzQ1n524+DpmSgKsCYDVr2zzk5ualwx/5f
Mv92ca5BGuMfwQixSJefxoaC67/eXiwgjoYpzv0Ia+3iZnWLtws3sIR736a4MVgR
GUJXKWL2yYpBAOMcvALNIwrqPQPhb+lfLvXF4I3ReGk7cJzx+XCnOoD5DEeJF5qk
78QotazFPPZc6M9mlqLsnHStworo9f64d5VS+LkWN8nIkL/tpikxV35Jl7Y6XAI4
a0K41LUkQXH3MWQqBg14UHYnFAtZ2t/wUcvhRfFT6TnVQgPq4O2AZnHYL2qQ4pac
vEogCYd3XEtqLBj6fQATwKXffHnQJQ4UkkEkP0pPaQzHgnnwskjimxf0NURi3Rz5
VdRGv6MxctC6knDUxkYJz+u7qJxGd0coNOfOyA/zJCiwEoY2vyisXKCYGHpIUB93
0tWNJg+LWlkHQUg9qN9u2jxDRbw4Rh9OwfMint5rLJ0T07YqEYq1tVXxDO9izogX
OaSUUzUqoT0TfSs6sto1nQ4qpqg5XzbhFeRAI1eXCQS2xoz3tgVzOQVj13ctWtBO
ZBJixze57nYxqNsXU6zqA1ytujAxvpeyswhTtwvzvWNYT/xZELFV2kko6V6QH4nX
Zxa/OI1Atrt8bxL3l4hk76WDWr1I7iN2kANFEugmU9EHQ9VfvdLYEw7HLeKiMvTi
PCJ14EYib4wDmMiSJNlhrGH0+ZdTzPV+bPj1RNRISKb9GKbRrv8qDkjoBwsm6uA6
C8TbAPZvuLQBnDQKJ1JMFjQSbB8hUNZ52AKAs0kmi32XKPhLRF39Wyx1efGRub1A
VX9kIHE2yoGF20UE9v7c6VsIRjtFsvzj6YHmqtrGgu912KQBNnmAzYvG7qvAhH4e
1/LgOaBTT88DoKiOybCOEk8hzZ0BlP6Pk8QG+I9gbUjqy2qBaKH9TuIMFiMgcumY
9QJgEHYSZoc2E7jr9HA7AOuJ/SJnfXeUdaKNHYaiZ0ajnE0/3JoYUYYseDj4WCTJ
Qdc/JrxWDczWdZm+/ve0NZmG0jQZUfs2TddQPrDdMPN0+llLAyUY7agsbT3vmml8
qBFfy/gXJOwct7jJ6MKE8wi99xsBadsvY595VAlFzXZ/KlOTXnC4wILUvQRzmqKZ
n2Pm16SOHKNqondll3NSkpp7wrNUF1yfEQMWfvzU3JOjt9oQbXX1WhJQND+Tqxnh
IHW2k3wnDBLBowXodfpMMeyOPjmtEnczncpO+xgMvaq+YXxh4yiKgiLKe3ZKxia4
8i5EDxYTZuCRapsoow2V6EJ4sUzXZmaimOOFbApJdQgS42xobCgWaBCu671/B8iH
RbzFEQwPYwO1TThy+LcqVx+MlBC2LkHZFcpe7hU3PmedzE3d/f1DIvuc/z6CMIC+
j9/APWu19H8wue5k4MjAJSGQrWE4Zd/pkln2eayHvApzolU2BU5z8YNruJDeKA5m
M7IV3eKqVUX6+vbHH54zczeyIZ2f0aOecLGTdJV/Ng+/KEdMinmQ/Wljj8prMis4
sh/PsGgimyVqGZw766zUxYFAnZ6zngGvRQMr8Zj+i2NN/RL7EbylPrYX9Gn76psa
WvRaRmfmLV70HwDf2F86NTkGJ7oexztg6++dtFj7pmD6+/ikDrQtNV43DO7msf38
kjaw9F/AP1VDWgMqyysNCHTqlse6ue4Zz2aaHIVVf3fDQzBpWbRzNW7jLo+uLzgP
nnklrBNnHUBuavH23lJooI5SRl3wOPGCfqgQCCREneZjLHqBcfbatJsQHbYRLWyw
bLBs1e4ggP/XcmF19eqbYgS/nTQs3agn3Kigv/8Rka6tghzcbP1ZMGed6zM74BFb
2wXcb6+4wKos1OTQZsxcvEkEjsV8JQDdt4eaOm1HUo2pRb3qc7qKjiqUCK7T0m1O
d7XuIvXGhByOYtw6XflFxDHqb5t8V/2qqgv2RmNcSJxW/FsMZS6FjQa5xc8mtwYd
o3kS6JqYLN0gEAkKuRx3TKyDqI39MyKlF/ag8j3/S/q3qyfqI1Eip7Qcm3fx54o4
zVZCKZV8H78+oQCjpig/0Xx4AgyZJzqNm9F4plvfWp/vAmzG4QwJ9G2dW/T8OtlS
ufBpxAqpFq3mTOzRDd5WSaTEy8JKObsHQ8oojq/UBSACzqhWnEvMZKfCDkRylKCv
vYTZOBC3cDucDiwppL42ZQbw7e+R0cydF0gjfFohT20Gxet9ZyGkgwvwnQHroZRB
4qGFnckO9ExY8Eyhtkb4tZ8Xhz3DM8J+YMbLDfXl2pKXUE9qOG41CRsi1WrRIODx
GMlb79Zsd75djRGtwwMUmspEEq+MsVII0/fTzhxprhMHEP3QoTA/f8wCI2OgWD8W
pYcVNQAaOa1fUxZy616Abrwz/RActlZ7xnzUUkQ93Vgb/jLUUuTPK+/THAxvNSJx
6BM+q7emwCU9JFT0Y7AjIOfm1cxx3yUEbkn4oxJyCTQ517cAtHcUdzYs0YYpKXze
Ik3caIMG7OB1+k4RNVTnj/udixyZjSvrU0BUIJ4ezPwfbxVYI9xGFo4Bh4pegyew
Irbe/LK8LCDDMOuOakJgEaYQGouIQzLFetYcpkZkWR1DZIiUr2fNqSPc9DEIj9Zv
hw5z8zfLQhE1mlOZ9MGu728q6Cnhuir3g7yl//Paywhs9+WJIj8BdTTuDTCqi8BS
bkhnHxlT0I2fUr4p4pQ8KKqAQZJnpiVfetAK5av3c3QpuR7gPfVwYNjoDoDeweux
JTLCUNQfI8+556wcqTMU9XgStkyNv1YlIRpBS38J/YRyCFrrxDxVH8ODaJEKbN9x
A5MOvgxsrWSeMhIFCaa+AtsiSk97cFfCz797IvyThxMzxsJi71bDvE1SWqBHgswA
6I6M5p1G4+SojW8KcknM1Rl8mENuNa1Ez8tM0PEeRYGv9XtSIANWNKnLJ2kGEr0N
8EtQeqIwHuW9WMYiT07Y33ILmmEtAZ/NCyOrXSTGq05/J+9H7U0XrV4ZxtNoaSGP
tvWxBGwxC2K9/WLetMOfjIhgL8sQHWiaLXN/orNr5dGTqT5NrDazx1HdCsHoMzvx
yaC33/ROOyfw6hG6hfjgVYtzt2/u08ISWr8Tr1uX664fW5i/kXqzssJBfAadzakm
5M1OGAokGV3Z8WIVKxC2QVscBVob3dqwI2OaU5aVQJ6s7eHkGB7kS2HOLP0xJ1ol
mgUVSPG1tr5aguYtDXQcV0bJq5uC+ySespaiW/iowEt/tAR3s+VV31luYaY5gPol
Rv5+nS6xeD/KimBmM16j9A4j1IPqffbePLdG9b2LYgeo7e86+QWvKxQmuSyVZb4Z
+uA7uQCe4BOPf/+XqnhnjFzHUXgBfagBRqjZZLseuRpQKl7NePATt+4yEy8PcjN9
NvISc0T1XOIaT0XrbnQQ2T0QCxK9KDvP3veaaIoY6LD3mUHRlGj9ZSZhSdMZzJXQ
S0jZg3+5sbYPz9VFm+JVZ9kBOotmDOlqUkVTjFB0TEpNhbm+qhV/Jrq5t5rnxgJM
xD/7flVAGVzZJAn/nwzTKRexWqFwDp2fSEZIONmjMCjGFQ8hqk9ow73Q3q0Y6YZk
unmvERSWsmI6LMYqFtsQfszXtp4JeXWpgIZ07IwqqFxwMIXGk6EJMSFQ5Qic1fEx
0NMDoPQr/bRZ17YzVWgveS7HC3TEI8P2Bu6zX16QLoBZEjj0eEnlOIl8XUhM62p7
IrzhnKdZgzmBtGQFcaZK6dOiPsBAP5Tea87GNDhSM6W42VP6qjJCzvzc9qlIopGS
vezQcBDs5w+QGS29v+UOt7m311v+nowDjvEs85hffEiHeZaYUAF2geMnr4JruhWH
2YfHRu950bGiGGBAFAkl2FoEMHXENiU3l2dFiPQF9p9QGocHyIubeKc/u9GD/bS6
7TVUqVJ0bCo2DOXhlSFI17MoqIs+e7RCRy8EypD9ofNCzKivpdcw7Y8kBSyPER5s
fbl2YP8cjZtGexEIewpDHfScVx2jXLE4c8d0umKFYBkHwn9ofDFHt6jEQetjGGC/
It063lyXXN/+UhJB3BtkYbQJatT3hnh389Xhyqxs0P2dIgxX9yKuAof3bgrw8XrI
1CKNU6rYi7sLDoAEbJodpWZmp4NTAgb9B+Uaz3/mRbUR0if9Z2G1SqB3pfdBHPwA
yw+qP9Xw5jbDiDvq5ApRoAAe511aT4T/tx7xxAJnVxxywZ1npOS5ccBnaOtJTFPd
MtX7NolkEdnPIyPTNK/OwH+h94HsTSry+ZrfGFThXE1I35DHwLc2z5Xpp1YPYG1y
nFv8zqoORHcVzCrmN8QjhLPeEzWfIOemS8whQkgJyU08+5XL50/t3JMAUsRZIYrc
67mcWiAiyl8iRoUGWlXj9cStchOjSFljYjf5Gtz/g/y3yeZDVv4osLIiK6GW94K+
qDBwhG8XS0YMvS+kUbJ88frzvuIuumtB+5VpZw4PvYDvOvyKtfNKVay+L7WV8cnJ
PEVChTo5cNOPaHiElpvr5G1goGYPam5ZDZu+0OZdJn95skm47Olzg7x7o09ZrGXi
s1VdnI0TRzyaPBjn4n6JmEeGDECc3e5As5R60jRu3xJGYwDyVTvn5wXpZvizObgn
FAF3KHZWKha0HPmVwr6pJSAv0fAZZjO4xmCfsFbX02ZKVPd0gB+G54Wg6nqc68z1
uu9+XPRgfg1KuCpvumc1Cr8rqyR2vcIkJ88hZzWNrTZzJ85+WwgANIrGU4F39Xlv
LvdelVWbl4FhMs+bm53lM+cEAeVBV1YHt+9XGucY8z4QJBZkrg9s1Eb/DwAD92WI
6qvT6UulJfwUVm/8B0CxxuvC/LkYBsskjIV9sG7ywaqGBpwu1puVUDRZPaTH87Jb
tpBjVBzNJ1Je2JWVw9Opih7nJE1BQMfSKNTJ/8M/MfNvrlXucHLrM3cIsHnvoYox
29o7Qrs1ebKPMF9xWFmuQkryERlv7oF00ni6S5+4lk+X5gCfzy6mf1cyp5PT/0xe
4tzuLfGgMGQlAso3a9YcUG/fok8LWEXQ1qhpT97rONdJsO//iN9AyEsflfvLqRhp
80NFtd7SLyW8EIUNgg4z84vCbFCP7mcLbRppisrLu+auKlm1/ZDyE1pANfxZ0mRM
4LayJYCknvt4HYRQkkeI4fFk17ZqEJ0IYha1DujktLfnnKT1lMeuyo5RFWcOd+Cg
nWc66PajsH8cvgQfZdGCNF64DOrmrxjGNLqU7r7/TpnAIMapLVIHmH5i8S6hq/Sm
j4oEXE9Byn3Zve4EAG13xgFSBytTbV5cAIgMCJl+A5YQm1tG1wVCit5pe+6geDRY
Y0J9RXBY0Smcl11xYDzR6LAk0EGveHi5R5Psk1/kfAYvyLgpJ7mFL+Dv1WkHlXnF
VilwneurwEQqjIu5+ShEotRXG69WfymieVp6gzeO5fDspgGRTVzYsNoqYpm8wuS8
8IVAQbP3MQ3o3NDgrlGMs7pQqw8xDic1pSTflIMSpycHapS8DxswulffYKPvHleE
Y4Fdk1EhZsMocnxyHL/y5AIJxA0WzyI891a0yuTrdEYUH/IpmztgjHukgHgFVqwG
GB8/bt3g66fowLIKppzYqSKIv6urJMVXv/60yI1MGhrQL4u9meiR/8bVjqsKiZzy
9cbxLgoSql7m0GywWctTbexjqMIN2hlp3CzSCO0bg8V7/87PaXLaivQ1V6nPlpAc
+/+rKj6WY8d0r7p8Tq7JIrTQhdttOlU3TWNRdus3d1wkZ485XYT9gxKlolvALLrN
qRhkm5nl3axK+rqvWBBFjPqYFjuRR0SXOKLy8qQ7Gl1b8SmepJ/OIoOLKSeKK7ip
qskbrotjqdV1uLYOC7bUA1/uASLMvlXBgGq4hObqXEhGC8FVkHcwJggPz4aPHm84
uqWVfSGS2U2IwTDqxXsMyhEz6WSNL1uHk59zBuRP0uyRSs0pWSNvCulAcqk/PeTo
X7s3SSvA70LWwcrBzBjPMzdcK+qfoq6pSICGu3naWWR70+JJnvyYqijDaQvj399C
IDtFFaUWtSviQ17dbTrJewJPGYrezKMfMbzf9u4oQtt22a+VFXXMeaJMJEKN9wj2
UW82bXv69w/ywkxVIkIhtwIpIyk5PmmBBUHQ6v7QgVVdjLAZ6OQdtDUFdYgleVsM
PIKziQSAEd1txh2TTlNciQZL29Yz3YFhI2qEaP2kf41Ak5TH7kdpBezsJ6m2tl7l
YZwB2uh4aqcSZvFr5dLOj2gDx2dh8jeFB7pOAY/M+rHAlwYM6uQluQs2bsQFlcUh
oX2dLMBlc56SCQrBXPIBhrDgdSsDl1yQ23fX1hNwJzd9gi1jse+h9XT3j11H2myv
JPumOiDfO3ZqSpOyNwpWaDQ06/Q4s3HQiIyU3hGuBN9VFVFS1YsLu7e0qRE2H4S/
/j9zUZOQE9jRr+nHdg79py7wnLGx9Tmpe3bISVgTypZQm/oVobJ4dBQPkqioP9cl
tFZVyJRUUOeGCDfVueNBHSzXECqTVjbSpwS+64rFVm6gj+GpHBTgviGJRxESpapF
phT40bmPUUmY7++0nXBrZ8MismqYBZwe/OihP4D573hYJHCZtBTSYu7fJwrtQ7E0
QRf9LTR4AW7gKv0bbhPnNlFqJc5HmxtUmvwEyszhg6DQ3oBX6bKH7Uk9bt+7tC+c
EAqpb7zCQIFa5rUTjY9okMEnTREbiwHQf91ZDG8QIZnRCtYJf7ighVgxkxmQJRTL
TKsz88rLYCYtFGzz1wIEXcIW4JNVSR8yIdOEe2Fds0uiGbmVP6zKyUQpzwT0+FHB
dfrOo3LIVT/d9f5G8DN+Z8zvSawFehGdKJpNxG3bgTmbEQT4NMwY7N1XUYN2tHRd
Y4S9/f2mzkhhpGydueVmvyrbGIGfBWVrJtKvxujGBDMWlvf/TKawEUjEcuL/lDE9
inACenoBC9aQ8t32aUsfnoXgV4LaIl4LFwo7Njm2rQ5oghyVxAuJw8OAVPo9h2w4
OwLiFW+FjeEw0ktC5t6OV7hS8L3QDbbLYbrNXBRVSoh748taqvutUE3ASyw0JoDN
N4Xl4o05nA5PC1zZduNLk5LxTTU2L+ClcTUpT/LdVA30xvfw5/viPl7B8ab8MK3k
dWDUFBzOopUN9RPbRdMNclxBKfu6B+pk9/kWIer4A0/AM9n78rAKeXTpxwmF1dqh
E/frAC//3A5deyt+BwnnyoOEqp/tT534TieDfiiFyg+3YPW+cX/xmlAjMw/UPOyA
o/btvyepcbJ7lc0fUGy0BJOyaKjaDVRdQxwJ25X8vSoAxBStTdGt9uim35dHqgQn
lJo+5K4G7Z6ngLYG5+4wlkMJwz6kb//qgjs1hNxRtABEkvuGhl2r9bxT25blNPYu
RK94xHVdyhI7pqWdUJ5Wo+L792j94FVRac/xL5dDPgWlp3cG0GaL8NSDWqXMI4J+
Axv2uNl+2bDd45sNwwUmf55qByEZ8grQsLyvV+rPmsHDEZQtkuzDdmAm0rpIdvwI
HT2g9X9Mt9g5b8U9Qm/6PvL81RHLE3X8btqU5MjclzeYNYZ/GtsEOlPLVOAsNUHF
ZwLikRTznn0cu8HMf9DPaT5XFdSHNlqeSiBKIdZ40AeXal4ESgk+HTy0Xc61MpWn
7tXv9Jvr/vjBYhFja/T2yNYzJbev9QQJ2X8ycWl05nH6StxGZLfR24M1ZYfuB6Qx
WHkXK7HzslAURma4gDIbE65NrcBGVDx8H0j25GeZL+xkkatdB9Uo20uydqIFB1WT
RL8FYTSGy/VN9WHET60heiQt+ozD7gR30mAekoGRlxNOwHRizzBdHaFsTVhBXQ+N
0R2CKQxdviYgbvhaiWPSt3qCbVbSU+Vrrg0ussNvsmc3qOEZfNuTMeTodl0xwK2r
4FpCaQCDHjKU/eCsI7IC5BgQjWXHZCi7jN7LsENc9joK4LIBkOdMGWnteACUrgby
VRcGUKrtKSXrjzLf7qxGHGtowrGNNUjmGT0LrcUKMmUdFljPvSeZbXG13YiEjlAk
ainuEZ7BVXVB04CLukzwSwvhI+e0rjKNsNK9OJ9+cCkGoTgfZAF8noNiVu5KhPFf
Wtav5Y7ZcQwqezYkRtQ7WSDRVTlZTJRfgUISRXUscQQ8jtrw3kjOzpgbpTZ1Xh7a
kvYHOEbwz6U8WKmJi6FUqpZSbNb/P7YuCQifTMqL0+HfcPd4Pc+ufHlk3IknWnUG
qmLRNmYSblRF6HHCYfqaCy6X9VWe+P7wpLerTLK6qzy+SmnmYkYmU/MnVpqSYWMO
lE0Q9uNap5JHiNLOh/XsEMLPROtljYuU/5MwuC1MKuljVWvXQi4/5PGm6+lFN1G2
xo64VuHjMmjxDCMSpX/svsLzfIRefr7mZ8+9l1LczVK0UJZQGh6s6BshUOY/5vQE
jtdMHG/aesngaKQJVU2waz5ohLdnfKWgi5KVXiaIGB6LvD6A6dFLC9wnzRtlVq+A
pw1iN8U2kDuZOl7j1NZ9HKRdvgC0rZp3pBjo88qq69KMUq0q16TXfGrofEnVK2+K
udoV4KBk1oxJRLh/Ozdi/yAd/UDTnRMNyFVa1zXs0cYQD6+MhVwwcqoXZOhf4pge
7nXfySJ432pfYTTk2j6nsbzroUH2fjqRfBiXKA3eOZR5f7l2YLce1IdzmMcttHiK
bo9LE+vZTgJFheCM9+cD7h76uKKdex2R9gdq69JbzBSzQa7czYA9+WtdWYDil7If
Xe6/SbzFUp1V3+xUieupncRSJDo8RE4h6oMi2cDfsSDBXarhdDuGPMB4dxDxJ3v0
Fvki3SCiqgErE41c7RHdtt8s6ZeSZCKg3wm3hum0vSOa1pvHwTniG8j0c8h3pE7X
jOqZKuSDbvnuDUTHHPqpJDgeTTNf72YkBAuv5Flt1/i0yS6Yixx6k9RX7MLRPJhP
/NVnIbKMWNzlBSlv6tPyp84ukOrtY9RcLR5ST0FVdiYOTIpD9f1yT8eDLt0qyLpL
OZLbc4Geli5X3fJ6fdm2gjxoStZSMbpMqAw1bdy2pUSybZNEq9W42RE0/MZP54AU
KJBjCKM+i9BL+DtHKepq1gtDcI69a6nKlUaG30V5Z9SB+VLLrzy916oNMB6ANyEK
AZEk30klz/E8uuEN2R4t7D+F26tZMj/rAqiudt5Tx7yfN3s9UMWthEG81YTzQHlQ
Mx6r5C4Kf+vGcbiSw0B5MqCy0oWYkSNt0QJ5v2/39exPcRjZn7guW5XRJlZCMDx6
v4GYQjxL5tf6ya+sxplA/pYLHAp70qu4m5rHLVchxHA6ph95e1sv++OQqA4j8kv0
G9LQbcJ6vM8ro51WmRZeqXVYfiJFzH6340LWZAZFEcmFXk83ATQiISqL4RGLk4+l
ldKyKe3bZf9SoN48oUNbkNL/G51TEMXq5YCJKYTzOkrXTsbjSCjTKgC2xKnwl0R0
vTrMhwoWWPRnaV+17BBq+WRN1s6eXzEzzToOs1LO2kz0NIaf2L+3hov6vICZSBd6
UOS3+s33uXEE5jNJ6Kim6rW7sJnOfxtXT7vG6QlqrpayLCup3bBD+40OzXl2mxnT
KUiBQN85KMz6SCIGBhb/SUsPAGIIaG+mNxmZfz6emCztZNtcEc0myZTdaJzg6lRk
yKNs4a8uArsa/CmwXnNI241nUWACpz1HSQ+9gUbw78DjWwt5a3pw+rvoEC66gV2t
NYzeQd4eyMJfNWq7ZHG+i56XJ83mDiI8COrag9K7UkCKuQ2cWlwSkHk/JxlkuYSW
n7ojkAtUT3DBey3nXqj78ioSX3xL/jpEbSoFfs+ElgHA8zjFc2ykNfecpintAogT
bla1DUlDEORWelMks7amktHclh6JcOrBpw6/oGp/ATH5pn6Syf+9+tyusCMk/9WY
Pi39ey8C4ESjoA95Iyno5qyxdHZdFTowM89TvIpay1tsrc8n7VplLZnU4/o+kiP8
k3R3MT0t0zN+CDMmCyKcyTYcutbjf4FbhrHEPhKl++1NSx//4mUzvAsM+mrzgePW
UCnjMt2LWyPnzHxq++tA4yxEVOFgvq0/VILbA6oeRUGU8azM0XlOUV1i3tOGrjFm
g2IEfjJlXdXW8KvnUaVFz/8VArewA65ZvsBW10KM0mde9SWsyyVSh4nZBWFww3to
4m0QHRdZYuH5tYo2fAWjNbYYgQ1MohM1Y9Z5eGmVjTXZjevqS94M8aZ2tPJasEKM
PDoa2czYwKyDJSLThT0KP6ZHBtW6RygmlcAuCGsy9cF6xHFjyViSouJ8+3Lm+OHl
zT8yVQ1WVhTIfojyYgYq/ivsTY93Joxnbx70ZA6Is0gQohAJkOmIFpa9WRYajj/a
G77h8Ptn/9kSObw2HBxIFudKMHc1NXBZGS13bG5dgA6DqhBMeTVSFyQBqPJYaOWc
5ZRdzgqJ1ir6ZVqQkJo2NPMF8haCTRrStwK6hXDSSKXqzP1rtin6zC4/9rmOZo1l
eLcg7FtkaOmg3kTzTRbhSHeABhnwUUFsnw9K/tryC/j8PMHIzRvBU5+ZL9LbPRlb
/pJCWvCpHt25nxyAXtyjVO4RuNHfNHoTKGenZsm4c5BguVFlblAeUNFV6AGSnO9u
e6bAZLheTCLY6Bb6Mu0xccnYhrV/HOBPtS3R5sR600AuXl7cAEguhGbDjJolkDlb
Fv7NjRQziHQ/6j3EAhgmCxMxGgvv+nvlCNRp6lZF/3Ar9mVukQY48Ro5dBKHogT9
hUdvKU0z00evZkMKDPx6CHLavlOMhSq47iLmKRuy8J5lcPev7x8NzgNZJxFezyOb
+1U9DHrMLHZlS9rBX1A2Wd7aWJ2FknmTgE0k/AYP/zQP80zYCaLAmPBxHkkHjJ6h
D5QBP59D/iJeT11Zg3JsUQ5t3I5/NoREsjKV4zB3mxq19OtLxJkSZuvWWxtbiGin
jUJgaybPQ3OlVGB5atvcCfcDf+ap24jcvLT/5JMV9dC6jNL4x+fjPUj621yPblYE
JKWxK0DedlMhyhL20koFq54xBj9p0i12sWvpgb7aosqeiATSVDWST8M84DNLaTvS
uaxEo9Lc5ox2p7towPNZMUK5ytVjo39Hln0XVeokY4w7cWuJNbm0ct+pGfLkQTJb
kYS1Sn9OIJ2L9U+XU4iijUstbHrBPgnxCAMcfbxqJro1H4Phpaw3K/sI1I4+R7Fm
ZRUQFF66PjEe3lvqgVmT1wbroZ2Wgccw+uJOca1KWO3LHZajzEO5ICbhVA5kj7RS
L1z2PTAOZwGlhmHqqWazDH9zExUzyp+qExMG3B0pmNp03hUkUolsb/q2HhU9URpM
eSrh9eMaIZwhsDAnttZp6XlDnHIttVua6sT8/mBpUVfDV67o7gBVbJuqxNJiNC32
itbTYzYNREMQ0jtUCtsMq3zKZtY2u8szUTMeNXkjrg+3BDYs2FbTI8S4uvO4SX9O
HOoN+QoyNLMARko7uNoJePnvPtnim++lWDOuAgb1gNKXfVmrA/pjfQKy/wSbJaZm
27ZckgebMmaSEcTgo/oienI4ZPwMDFago/SLQxnr95oMrrIF9ptApJZABBWRpU7r
FgJ3tvcgwOaUpqQNTW4dljAvsLWAMux+iUsZ4eUyI2nqGahqRIg2YJkiEnTsgrqK
7P6vOT+Lzz2A5kqOu4u1maNv42rt/bi2DoZ0paA/k6lbYld8ISFtWiAzhLZL8oJM
N5fJt0QCJJ00cuHcKS7bOCfckeuKWE3/BPezBQr9gRQa7ZUknzs5xpOXdYbSJ79b
362EsWIq4R3Gl0k3BBx2kz4vYg7PnsM+ObOJDQCyblJRIpSKYCay1b9DqSLofua8
TyGj7WHEQ92GW4SlhpnVBzNjhrPex0lRHlXKRuL0FrKrnXIZPpCbtUNaj188lVk+
LAtV2pKjIQtet3XQpO/wdnEcYtX7FnfJXvru4xB70/3rccFF+n5bYlEhCjmVLtnX
RjYAiIRKwqrJmDpwTZURxgT8R49Du9ggCTnq+/cSe9pTC/pJUYC/AFb+THIMiASM
KAr73Sq4NYt2VE0JuQ5cMCa6wZherF/UxHIPONxT6cORdBDcs6SKwAkVkxiNuYaq
nVt1tn2KMYEykrT76AJ57cAo7Zdf5hdYzB2Pg8RgqyPbAh351HTOYlviVHmX+vai
+dX1Z8HAzGuXxOrsyAsffajFKNGJTjbqdGwRdhTetaaDGKEwqfiK4AnKaI9sctao
pfqITFeZg2qObGq0KWLbi22kQea2oOE8p0A+guolHU6nV+MUOmJumYCaMOV48lxX
QzKnXs0Zj0T6cqQGp0cnqLjgRXTzUoH8Y7/9cAV1kNbSbqP4VV668lbtPhAjG2Mq
NsrMFft5SkIkUL7ToecZEqNHbQpdCw/6IgM5edMEuYkXQhBMje+99T1UR2LIcmMi
jmJNmHiiZzOrEf4Lg9X/LCfnJVnD44xHK3Ih9nEf8Rn1xsOolj0hdQpjRW15rPxM
7/DaureM1Za2dZ5ZRTULr/gl9Ja1UWJ96ux+pzKwwjlQQS2su7fjcGB0oTFbnUZr
B2vMMNVrfDpyZ6SnDLFkGlBNw4RY5/m2bvnU8zmcqQ4TxBSMy+rnDWerpm/hBfIp
waafo8RuE/Ta6YIPONgm3TWyivC8jcLvRWN4IjRqVd8uDyR7l2LCFVyy+vZVLh5R
agFWV7gAC3dENRt9RA1Ja7qUxgPV2E/pdHTcx0Wg/oxeosEyF7r6nBC88KF1OxUS
Df5vnbdWftoxRIgwrJzcrnoAtghaxvVkJY6yZKO+pP/YC+XFUT6gRE/BkVBwU+9q
lmSQpLSzM8r7HPdC0FpIS9oUe+smXpSNYpT3f7R8OioMVd1GPHgSEMh+3iWSCV+c
DEgBIyWCRqj7pMJBLT63rw74hxeEzem+OmKEs+nDHJP9ZAS9W1hc6OLRmxe+VZZo
rrMpBuNI9+MlVCt3RL/Tw7ATBaVLkLwv3tMT+HYyIdzjtsChUkW/xTr+btTUXsqY
AzwppkNzgJS7VkVmZyFfzko980vp1mI5foHfMSrYONbPdfUyd9ZJ2APkP5j+vA46
wsHn+UnG5NigF6+fcO7l4mjQ5gCs1j+eKEahBSCbcMWs0Vpe8lJ39er1OgpNW5al
awc0LeQss/SKnyaHQEim/DzxTflu/8aMdk4XuaBbJHDVEsm+nZXiaEJl3hlLdWa/
bfkJqzfxmiU7dOQ5XN8xG92+iQ+RDRgU6RGS0Aw4JjmB+9iZKGg/cJJS0Xtts0tc
PPFAE2sF7PwWEvkec7SRs8V/YKq8G7Mix1izchoN0hX6VbSlXxDFAYKA35HaPwqQ
DSD+jB+UlzD5rXDbLTbfIaSvHskwnp1j/2gaZh2TNHm0MMDYdeqbriUh4y413K5+
zosnq0WHp+An7uyFLFvWEdeDx/Vsnh24NHJAdqgiDcBEof9rL0Yp205oI4T7Myid
2bM60B24m4LlhEQZilpChKRuw2VzSbBVM5qocDFawySQym+hhroYddsUTj/jvaWB
gP0J0LlbBGMu5LFhZBjeyereT7UXmT3Jzfv1iDyOS34+xKMVtyp4FoSYjdk/3eTH
Dz+1c216XDLYpoZvl9QkfNbj3u4WYALbJFxeHPV6YVno0M3gm6EEMgYXzVjBeWkh
oHldj4HZza4qsx21EybWHZYIk0TyH1ZqU5/USD+zvD6P831DfoxFAmKe/oq9YsyS
JKl/TPXqAeKbfPWrazaWmH7Mq2rSi1ax7NrEuufgaxHxRBJoisQn59ZjtX/svACa
RFLxna903FcM5ZzkimMup8f7qafg5ax7qVz+z7VFnVRF9/WH/fdKaF1YvI4ArpF2
38pYr9KBrL9YQHJ8Lz0BwUx78dl9SozdD2otyNw4/7juPEgm+BmoGfXkZ5s+cZRv
fXZdcpAsf6eN+1D1MR/tjoIh5OGP/35dpBRmFTNwkJoZ4nhRZKx6gTl5nSB6kPND
UP5xyf6QxrsJQFd2tua1I4JDbGS5k7T20Xmvml7BmKWzn3rHmkhJb0vQsbEtiXlt
RJjz5FvIZ9s7acieVBshnU4kZ1wUcQj1S5AhricUO24rKdecXZ/XbV+LrHr0T5q6
rGsvFPLlohXvI+XgZ9kdtq3BtlaPlqpTdkL9GBBRMM9EatY8yrmxhymz27POATs5
W50K86sfOwcd2GZO/3pcxbSH17z+RYtL5apRZvNvhXbuCsmICABHEBjSsvkopfVE
SU9ZaOV8TY+i3BGoC8crGwxLoq+U67s8/mzm9dkesi9+HJAW8AnE+a0L/6dh+r+g
7//wzwLQknMBonYJKV5Ep+iTCjoM2Ir+5eqcrcMl0vMPpkJHdmh+3qW8CzqhTDMA
vNlrPWxsFD5bgIIbQlaWW5oNy4IPGRoVK89G+ySSFYQOtkcVIz6ggW4rrz0M6l0+
jpmQrOm3xzk0byNy3N8kIhYP0tgH9S4/UcGqlXehyD4+Eky0ZHom+hKxpoymkUZM
ThIkE9FKnNwl7v6Wp8+Bsa9ysp+/RWk9XqlAwQiRpP5HGKNw2TIgyNXblaN66z97
9d6YHP1m3UqIcfBSinlGuW0zooDHwa3cNYgj4UMS7UYLbYNs+9yuDRsEXa0g6+Dq
06jKzy8gXOyNZf3fOte1HORAzbZ+o29uo+4uKUDQAFhWs6nQMhapFcoOfuMyxSRL
yXQSyf3DQap8v0zeEZweG2f0OAf96WF7bc+hQO7Wmg77HuOaa6XWgG80ZqMtl5DL
pvP8jeWXy5PVDhKEkr6h9Y4yC1E9DZdaoOMMf2tIyX13kcL6at5DqVs0/uPICjND
KhRHvrZ3Nuhs6oRlW49AINwTXOpNajyc6A7h/09HOFdPsvUzTEm4ifba54A6D+DD
ctiXM1l5kSCnJD3O+GKTtK/fnlqbpUmQg+I0LtubaBbxuikCgTtFxUdCpXpbF8AO
GvRExtGNx8crQlxlqYAUiy2e5rudx/q0dLj7t+pSFMpQlt2qlPEz2D8PVwCUSRIm
Y6Vjo3cwi9uoAAjF4tRdh6pKuPAvPO/pdkJhe/hscJ7v+GBo+c013IHbRjvbjOTj
hCftHDQxgldf+HevdUFfH4ihZJsmC+tQ1mY7mnEAXpv7oIOyTEMkSlQi9QjzO6Im
aOtnxPEJuZmXy+OCeejUssBl2MZIxxaV+YnmlQtkpJ1m5q74gwicbVkkdB8csJ40
bobdhnmJwTJWcSxb8/zou2nsbMK/RVeCluqJ6zj0kN8viMvZqqz+3RD9qm/42oRN
8XDMDwnCkeqJOoaUOEmp0Y7k7o8BIVnOG85iZPAPaYR+RTGJ9INm2imxwCOl4R/v
bFz8mj1F83KgY7sgXULE9t5iXhcuxZhMvavkh1PUkCNCiVSzDg3myO470OgRKUYK
RRUuRpzDbz+EK2dByVCgA+eH1zSx2GexOHJAfHwlH4Iey6PImvZjQizTuqMs4fnL
RXPml3djWPlroe+EFw+AfU07vY3YyrULYbljMA0Rd/OtVRxkgegbk/H+1KQ1e1Df
AqQD1iNnaTUqcwkLeaad4IfcSmCrl1KdkJhRszR2+8zWOAVao3oBu2jYszlPe3im
knfy69Ba/D2D9mHq1iSvN2mMhlcuUE+24zNzI75oNZCsX9cdHlSENkE4ukRUSjdU
AWCqpkRnjq4B04QSKAjToVW/VtE4cXlbkA9SxRBH4iwhNmX2k7xSQhLc6juPpO2d
fPm3GHtMzHKWCn6nl328DZi1afkpPjaakUE8PBYh9EfJ2oa/RRdeEqKL0Aa4ro2l
w0CweOYvjNzPn/I6Ytw/gjlIMsh/gI8EPqq0SINrS/+iK0Qv2JbmjzAKKNZW+oRd
oCD8RwKBkMESjANCGFO9SaHMYhyw4efrwn+O+l4evJ1lML1EUXiTVebnJtjZQb2v
I9HUzKESatk8CT16Cs8pGdYSVZU9hj6TPt5tKb0mQ19Xaa+OFFFolhdGHas4S1aw
9aTtPtiajZW9BD9Y8kjsBNbUHQJ6khGwqct7gSO1kTdbeBD6fbjXeNAEgvbIIZHr
L8f1icbJBOC45G9kkcc8wyrkYDZrwJ3+b6EWAVoBQRZb9GfheHnbuycqR+8WJlPW
XXKJtf7HLPcVPOx1O2mplYmbSf7PAwifrOrlrDOvHfUCwo/KEbdTQPw577K0SbGQ
vg6NrzJsiFy+7uKHPS6H+kyThN/3hC60paQYCc0NdYbUL2TyG9LqTGx3nqAqnbsB
jRaT73/2xdLVmlXc/9up9KYpGQsowJeWsUsBbDzbsYAav04/L2Crav/qWe/K81OG
wSrdIw1zeS7q4zg35dXpQ9IIGRoAQR20WWtyMeA3r9jw6P939pZuV5LPfvC6Atmw
gWbgdS732kkf+tN1/NpYV0fRy79jqP2uZP9wijAbVMuxUR3pq6z/cTlhQwzToUgp
JX9tVa01o5clV2AbuqTweHfPqfOTb/4WbPKZN5+Wr2KjKl292kHdaP0zvM1N27AY
0/JPSnK8f1c9QJwVbDCl8FWxU3CHvfUV9WbvonZ4sWFqbiHOJTPHDvIXLchLGx/W
qmq+E9Zr9EhYcnwguwCkeDacNa0hmvAnGwyhEt8Acqveyf8G1iJSta7qM/IpKXVy
x9UoY5MG8GL0007kiZx5Qq4u7hT/23nQsHPgqSyPsvaDXhBgMwBrnXy1UG1/PDed
Sto+vROiBaOsFTO/13uS9F7rlU7b1lVs6DaoWRoT9FoFcwm0Q+Zt61CrsY6OJKMi
etMac60IgzdYGKgyxcQudITIKgWKRYImq90VKpUzJwqaJdpfwGjKB6RGeW7mGnx6
QbbzTKdpKJZkS1y4+4k3nHMCJn4GcT27IftP71k3P2weRraZnQe7A4FUgBWh16ud
K0T5UfD908FlMIf/MhkxFvgAU4hjPYnEIMpt3wTKsl+ghItDdydlzJC3Bw2JEGIj
Fbx9buUEHBBp0ei19nqmXlTwq2GTBr6Kkl/jK29GDFVCLgaFThDV0bgQQFYPYufO
WOgcbs5cZZg7q8uXuLAdCilVMxGGmhj5FUE9EZM7wOnpPdcqSKuWN5zkRnA/JGAx
QpFxlisJWURu29wt+c3jav3LuS+mEsIxCESrZdjqS13G6n8UJPv7QOdugYAoZWQU
YafBXBQhO6lvqBjMjT86WQvi/Wh9wKWS5NwWlYBXuwE4vpl+59SNCULmFMm0/uGM
9+eunlm44sr8Msykdho/oI99ZgnZotzdkuJviVjqf/1IM3MQZavs80f1z4vDqWW3
zH9X6Ya6/5z1yxMtD1LLjCaymV5HKz05XxPSydYczY9OPrJX1xbXJILjTYTvv31E
w18fArmhYbGEIGCEWNWI7FC5glaZ1Xn4bJ/UmZqMXpMwx0jd6Z1FUw3EupVVQzay
UlMcAtdkFTRmW9vjK+QGByNgo4mXnBDjvvpXwgw5YTboGeGUMkgjUmwaPbQwHQYS
Tzcw9NjVTrEAKIUpoeNXOpm5ActVLfMo64uh0xRaOKfhlyzEQWRCs4QPsJq8pxl3
2BjixBBWqJr2N7VuqnMg/zlB3EYvJLNbhL8flQXVZP8Epw8oyb4APce9qlEwtfXO
s/i83ZYWGx0InIAPmx9xtCgfwciysybHrzkMSz30ED4J2kT7awno/KcMRZwDcY8J
vbN9iT5C2DvgbsYBrLwGY7qie9ZGyUCT9nvfrwCIt3saoM/mwLjhPKPDtrsKAmyE
qpLJZ1JrceTzgXgGKprVUe5nhH/oD0zPcM2gvkfMNy7oA9FR5wt4r8o8Uzi19QQ0
Tjf1ydC7hecfcES57zVZabvAB36ZwzWO4CGWxIWlWfQivKtVEPd4u6YEfqlYAOkJ
phgRKt10/wrhgFr5wH+nBGXor/XoSv8ILRC106bDZd8IXGGSKrEw8QiTICksC6/i
BKbdVKKdFyBDwtxgCI3yFtWQpeL0yrmmhFZ5nH1l7KDHr+GBbCwe9Lw2EvCsDuV5
Uw92k1tQO37ge/G3aQHv7c7jXTEvq3EA5K7VYiCFQ1uXyGMNLFgrk6p3solKRXUt
Dgzewzqs03rHQseA0I1VsouWIiKXna8hajnUOBnOIGf0tJyQF1FI9AUcg3vwt58K
qpIWQYlFJTN/K34pnwH6X2bprLciwPV5zsTbblw0PPxCFKg4TETZRnagy2D70xrG
ACNyuKcK921+Gt2Y48bNCS+Hc+kpnYT43l4ByUfazus/EaY2FTZjCUf0AkFiKDZp
xWRKhWNRaFfbhMXMpXb0FKbaVeT5lr5GWfXrereFXxvG0JRLLjah1FD8lt1b2lqZ
jXFoU0DMzQI75SsG5PQYKdQPeY141OjvgUZbNi0wNgUknGOZpsm0MPvYe5DGLkec
IcYPaptfbJjtEht0XTvulldzBNdyZVUqElxcfb6YELWeM8lLH+T7NH8itNDTENJ2
iLrWtknb+dXcgSDS+eVquk/5r/Ihzqvxn1tyRsnv6b+QhsKnkBweerjRHefCWQXX
BxaGa4LBandOzoIzrzfBYvtnR4BnJokcrDnDLf5dsHtD2qpDkXIeg3BEf0qxEoiw
N6OjWWxjnk/I2PGp/sklrKwSMk/z9IDaM/f7JCVV3tzPWxR1XpiESVNMecX1n3Km
9gr3whcL01IAJMGD/DmoJQS3Ar3hzHIUlzLZV4LujkGnHk4VTJTh/8kdkfZADf1k
tEcbJdx0NeOVQo450DkMzZtdq7CBnrn5VUuep4TZfpC77CEFzfPwN8dK4htXF+Yg
HxKcXoOw/H6j8a7LIl3srfVDGJHjMiSiCM2VMZB8VJ+nUpou5i0jr1ywKuE0rIwv
Pk4Bgo9OXtkfc0ANiibOxPZir0qiYK3kQhp6D8ywA+rSw/B5ZMQhqQS3tY1P8K0p
RV3sdU2AfgFmhSAS4BuFFLiN8xMGUTUK842ZXYhglrW6vWy83AE83lC6eIQQq0pi
n9M216qtQL48hiS+pMkmBK2k9TLaEbNfBQnoUbsW3ZHbLPqgxkAHXIyvyY03BqkE
upjsGMZiPxeUR5RR//CIKtJl9Z43eAJj7glKl7dzTINjvjkVbfep9b4dparKu9sJ
cYAaFZ9S9vN30+IgvQJBr5cAdIL3wvL/QA2QKfS5F0bd16w97g3W65gX4do6/VqR
VbK4vit64b+RNjn9JpbG0KBi1hYuVtgToajtz8nc9eEpl/xFPMYe6hYp9ctvzzk2
2ppkSM0LTaQui++XZ7HUeFsmfsH/Yj1I+e/j/pc8tvakllJfVLu/ohDx76AYme2h
rVqw96W9+G1OSQ4pyxkDQmqQl0GrjKZk+F1X1HvXr6LVSDgVebkExBgc2pb3lYJ1
7so7ps0+4PJh9wG4nph8voLgiqHZQhJQLvGu1AysblRtd7l7N3Y7ErPSci0qAFUF
S3YyfVqTDKx5XODZOMVd3Zgmi41ZJdQyj6aycH6koUUX1hEDXhxzO6eTHy7eSXmI
LltQDb8CzAamOf52aCVEhV4KUtOMZ0fvOGXCPGaU/yf9YBhneWvJ88tEVqOZ/UE5
NcUfRBUtzSrBI3mmTPiFLhlntpv0zNrcwYRGhRs6vDAYuPCvXv8BWsX2Uj37ELr2
WGWXNQchxPoLjsD3RevVwjcio58ZcN+NV4VjRrbBjNRyyK93o837XmEN7VcioqTY
scvDFJ5Pxd38aMfUe+3kGKi4V7xISNUqBbLRbFehHZL0ER52alsW8yb6xs0uKMF0
bBoo5oL2Vbm1Jt5RDt/8hSLxsmN6m3PuUIF4HoPyhviBeeqFSxKd8yQ4MPwfj1WS
AotWtwLj9s5NR/mnMEny7ue/N6v1o21tvLWTX6bAMKxYEWBKG0l4h36fQCT/ePGb
tSQTxp70XIilpUPNsllpO+TI+hikQ94zKBL+6/JDKZjLwxyVh68Z8LGzoN3s5qRk
CCitDT6rsL215NRNuVNJ/ZCQji9BmMOnjoE2im/BznfN2wxfH7jnHBHeCDGDh1my
T1aPPvLjQer0EX5CKVsbjEIBhZWtxDN8o1W3ZobZU1mEiPQs7DPEAMOJTUxI7NB2
mXDySc4JnM65sEzG5xkMZoIrfDNeIOcMYS06BhmDvN8Y6k4g6P5drOQ4nki9cjXv
M8TFAEW2tO4Ap+YxCzhOL8VOkVcPjXSRY2G5oDK9kCQh/aOwjkPq+2n/llJE+Kfs
3h/Qb01t9GVb7PQRm/4wSQgFAFggv462TJYar7w6OccIvkU4gBsSE1pFXjMllAaM
aFBvHd9neb6RpWiFOAo8KKeK1JCzvjDLFRg6QVma2p80tx0FoNJsjur12Sk1gSEU
oOxODJTapUQJds1csycJh5blm0wJVNzdAzLjzR0A/V16pcsaqxJdZXE4kwBCgaoB
OXEiqa4+P7148LR1F4VnFKQrDzNdV71BU2uIAO9rMneJoJ+k4DVuIzJrmiVbdigj
Ru4QdycCDqRwPRPd0TNttbxU+g7KVomxfm1rG9K768i3Y324Q1j5W6UIyTSLJjZW
eNv3fnH7D4y1CpUvbzXQnAMCAhwFFTzJ4rCMmfo6yXYOLK0SHkr3S9NDJSlwovli
cHQr3py/EN0GbW8VnE6Q6BJzKK/0e7RsJ/PvB1k8lLGnmSQN6Ve+xhyv/57hNyIS
/c74+pONf+R0tOXzcj97iKcbfL5IaAw72RQARvwkIINMNEKc4PfHwgcG9xnihsBi
lwEz76kq2NSaLCpqNZ3KWFl7nmK6/2oMYPQQmH7PDAmichQxa1R5XfSf4YAhIj8+
+0YBaHWN0bjoJfjFW8XkDw8f8Jgk5Upuyzhc/VEGZed5Y4EJvgyslvXMWIdzLABB
mi1O6A3gdtsuK2TQQ8YJRUinPrnXsW6dfpMNAdKXvaxOtaJq3BH4X/P12xx8GdqQ
XAUj/tvPQ/JjspgPCyoxrga3M8eMckgi74mowlxFgroromkZ1E+Kjc+2uaill7tb
fEg1DsGow4GfvKgddd8VQ5ewFKcbPbJUQZW6u4PAQJiXjmpJCtZHE2PttyM5P8rg
VpWDOeSzX5t9GbcjYenHy1GEmwTt8qUEMxvgLr/IjTWESggwBi1Rquap7EcYZP32
F7ZB7EjA62hiDzNEAVexrqQvmNhryzfprY9xfZ6phPdlVOIh3ynENAYd29KmV8CP
GMD7/X66q1gmWPVwei++kah6KiyvrlH8uBY9l4vN5P6fVyuslagUJwD8hv2x0Lpy
NUyq15W8OhZbCn/VLlXzSBco4uQAA+4SEZulREwbHQUSefqW29FEkumm1BCRnxYG
y5xrgC7CW5+MKkj8+HG82EEQZI0hwJzvkbiFitWkXvAGTBhUSiEqaDWjr64hbi1g
iIRSqd7x2LzbcJ1/LtWN3z/5L7w2YLbT7cLTj1G6Acy8PZsZ/C+ufduCplsGNj1G
bqmTcUhJSfWEMru8r19gxJbVQlecetCowo2mcII2brRziOo465+RSHUr61M/J1g7
tKPc0R6HvTDaO71slnwfHsyyouqgUIrYQTn2eLiLasB4+XwYTGG/uImMcSQZT2u1
xQcSGxUy2W3KGsX9i6lQJAZogOIvbWtbGCfHrxZUG/fTajcDbIpVK+zCIURwYw7C
qya496zbJztMAYsEOoZpHoJcO36gfhMwHxPYKqxqa98rDPuLAjC0T1GwUlHFxbfZ
P6jBv994lFfE3WBIEO2TbZfuAZa2036565f0IY3KcbrrXejHsjWKnBdiVnmiQtCz
fGCNPvNsH36w47GKqxn/CCmTTGbA5yjB5OM7OPFtbAGcw7WwWpeid8ftoEdmIv08
i0T/mUZB8/DCQZouJPDDY670utEDwcg9gnYzP+Q1SEfw/LqCzY7KvTe/a9rogutQ
Tjz+ONG4WbONZmXgl9NhpW3wf3c9ZrCV9nNfIYBy0d98raGXxl525nO6NzVkPCVA
Oy5ThITdIOrl9plOa2iniWj/A1EW/Chv7gN6wHKDWlrFlEjbUiWnZBSPBIpbnGmN
zgu31WDTG+ey1NWHCW14lxiBFoUlvmIONA5sxMRzgw6i2K+EQJkSg4pZfAddLqFc
u9lA05l3EGuQ0c3DOgeRioKHjFTut+qIqvSsm3JJ8aBBWN+T+czygZZ3KAOb0FY2
8eLUOhZOHl7bzZRCKyS66CnQb+noMp4k3905HDww8gEdSSApXEkve9TobJHAPZXN
B06WCjnK8DfuD07k5+VboqlC7PcIgyvTdU5gQsmSM1LQDFW61EqbfG2U39bGBHrj
rOpoUA30hVXv7eC2OMDoIeIbzlammB6/8OBV72ByY5+Trt/osv/NROAjGd3J+9Qv
+yGh0kYVbGf0GN5Fjpe9yd0lTlhesbPMOa3qcozQnhrDHr6aFeM/MDnUb/AytbmN
cmwq1FdVJIQMsUbLXmP/RDPn6YFhbReEgjJ2aGljz8cv+8dZNKhC0ZiSzy8r8n6M
ht67/OzbOqek7MKn9AK/RYMAfLb1eV/wfLN04nu35Gcsi8iClyEqTA5NUWeuKG2q
0De3KWCWi+3F9qKFb3Esw9REm2hLLjKpYYFnyh+d+jCsPqJUDOC1Wp4u/4oZaUb4
jaoCbJM3LOecd3sCZSEaQ+mCIxjDVdeawPDabXSfMitqXnc+5BUUP+xr5F1ugvY+
Jv9lxTstz/9cBR4P3M4EBAyQdEUwyBmOiKXTmvrkE0QDHSmYHbEU3N0Yj2qzTvCk
8hzWAgw/5PNIic/dtTUclQStM4TAd4Mer6f/3942z7BRp26wvGcaDgLi9YV5OlLH
fqIeiURG/L1aAjX0HeJ9N1zYOp788brxiMcKAsI112OMm4seT5ahf1pVd/bRV1Jp
7fPTwraOw1KQ+DOtCgWqB7aEbC+TOz3tZSE9FAq18Co6Ga0XF0W5Kx33L5q4ZKbn
+Ig/tTYl0DGVLivR9rgIyDbVEKhsaNF0xSARKAcqCUxssHniK/b/b48FZGpPfXeI
UG7TPCp6PwZwDWh21eUVA6B6od+5pscuQ3AMhjcxeZd3+jJgWXhyUtf/u2maEX6o
gNCRAWbMisyOD32+B1W9KsMKvFYmiow7I42gfHMxxmdhFqyO49Y5DABjL07LdvRc
+WS3Kr7OV2YD0VB5BVRIE8aoJNADpbzZrFyLDNiTc/L5eKs/YtPNpYWQwV1juX1H
Xzk9y5d+4GkcSUs4qTbvhc41jaFZkPXJab8sJYJaOPcXDURWXhFlbtmgB6pYbPkw
vmeMUcT1Gnce2M4KXJHxs39pqqwrZZPPIic8HWhQsNCl6tA7vliAgN/vrLyK+IX0
HsPyphrAZPjCcHjn3d5Z6YiK/OdOOipmkC+dXtX4dXYD3Ww6wPEwjfucc0ZhqHUQ
He++t3He5jngetjc53S0COYcTbYzTZtGUns/p+AMZpLVbNuZtb2lcNDzW1gTxoT+
W/3FJKDBftmQnC59F8Hglua03EtyDB75pzR7o76FbxFWLoAlrD5CCMbJfeA8Boni
4RRZwmY+qhTnWK9jB6cLmUA2G2iI/gidGMRgaB/R87UE8AU9A97uu80rgPVmI7/W
3P8aVd9noMoK5S7qak7oicf/lprCZ8kroocOA/9uaz/yu82pX0P4lJqmeWDc9ICw
vT+E+qnMZ+3PegAUjudf0ZfQOH/+9X5VEBksY6lCB3B4gook5AnGbYQO4u8VSnRr
Shqq87OtP62iMVd6eFuG3rLGwQfWXIHP4l27UgBfY/wIITZB3cBN9Ax66ASqg2jp
xmdtj6GwhBUXrUYq/e5nLUpfdwo/Qp4jj1LBZN3TndonOLfpod6aoxInwwuPM6O+
GCd2oRjBeJ3gt1zaMGSG+jOKvqlUvG+z2EhIFsxMG4JtnhmqOT5sQFaOVxCcSRIf
6XUyqwD5ajAL4qhlN4jZ6frBbXOrFncoLggi5TdNdoA2P14kyLloI02nkSxtBRfw
CoofvPlSS2f84t31XOWk/uYjNqxi0unSVamAdaQIiHSOcyWCYLZQuSA7BAxiZgjm
nqyJ5yyFkhaCqV8MH9kHpGr61KkRz5EM4D3AiyOqx+dslLYEGADQCI2ANYLgG2Tm
36c4ZvEQRbWAtt/aLfC8od7q1m7wmInz7xV64BEpDc/CXgn2VBFdQbfazg8vLour
dR/cmHcqyql0HMpg31pv1hr8Zhb4PnYaqHj6ij/mC+2SIyL8pcHr6ZeysLw19760
hablGjWXM143mpEvSzyNO6hJC8TMvNtQMl46InzVn4Co1fLiorxd53XHmWYWu7lp
2bbnaWXRvBXRGMyWJjhAwwAg4TVaUVRKBk34sgDn8SAAOePR/AIT0ec6MFqpVcF2
IqLqGSf4KzPTKG2GMFgj/wx3oR/Y3aV/SxwleSdDuuMATKh/rzPkrAxvDtv1WxTi
0Lebwoes1b4IQrzUwjs4GR3+NaMnzh9WF44833OWUgPvG5E60IUKkW4yZ6+4E0VZ
T7BSuDnbG2vNOE+LO1PCK/zZMAd/IU+QbcChDtPbcgZHv1l0osuswSX1KyaDBtgZ
batHOH4sJDd091e63WVk/U5+dSW0uUK3tH3b+N++Qnri8PUNJ7B+w8olEJulfVED
oec5KDqNV2R2kHJJGaJVCA/WXQtNcPzP2UShvVcmnR6zZcXp/rdeutdtPFyeCA7b
dPDnXMg4ZlGTN4hxrH/IZzbC9UIBKPTl3V2DOPFnjBJVLdVW19ouQ1uNwbo5R/+L
9gYLJwFdjzwNlqt7X1hvGBYIwIMRTXnf+R2W1WxMaOobXMbYJdtZnBeUlFrHs6fL
BqPXqIRbHc2yT5PL6Si09XyWw5xWYtnPeWfgaiWNMVcDN9w46uJbgLVGT0KThkpA
nN+Ypjppw2b8EPbEp1lO/x53P0YcT4D5NGcYBu4/oQLvkURQ84vTwQu8uE9K0GQA
pUINREcObg8opQprTePm/jxOaX7ShJMLsWBMl97rQlchX3xCuJbbNaUX/SsEXFeJ
3OLL37lBdGqvkjANJvUNuWagTRERORQ1Op5ha3osmuKqCrvu53CW9uSnALUNIxAu
GAHqhXdX3N2rgYMzmXBoMr+mfEh0NUVS3VSD3zgrDf0EOGjCh+s9UvMfiFm/yxsY
P+kNmFTTCAEDZmTtXHHHIHIGDev4+snkK33nDjO4WCGdNXpVIhDcI2DSoMVV3tat
/8G4J1XZaSuyrwXmXpo8yE9z/U7sY7WAwVhmi+t7ircmzbfUFvgOIXNLr19ZVfw3
OLyyaRaZ3VdXd9sakdB6A4jzDjqFLpi4wvvllBUWrtUoH+kLZQezcnkOxYWULzrv
pxFMVnQsWB3JlaBOKnClDthe2YsL2MNOnMe3g95ePeh/UodXP59C7XRQb/s9q8eB
IO7JCTWBdvUgX40oAaaUAbkUdeotm+PIQUEuZ4WgC3o6CDCCEXeLSRTvP+Aq9mgv
sK3iJmmazE41oGuRqpzHqrvbFItEvJSm3dDybpap6sB97ukX/9RPxUl1UliARtT6
fPOZh+Xjypjkd7RJWhDNxXvlC1JbJsQ8YOiHl53CdSPYyuJmSJIOWXPFFWuuCUaQ
YHXlCZzXpki/vF5WEKqExS77myOlwBBjC/ZfQqvgN6DawNzoHSxxJU7kmbvpxkA7
7MBR5LEHOBWIcWEL3HhV79DlUjzFOYY+P27Af4iGpEpI57CzDeyW7H5I/qgfCjFx
0Vj2L7noEhUqLKL0PjEq1piFh7O5OlbBSpZZOVhfGoTgZGtAs/OcZHfIxwohVBF8
OVNGGTJjOfm485FV6DOubHLD+xslJVCoCEl1ydebA4CTIV5dcOhImY2WKP3igXgH
FjyEh3dF/0FStuOiaz0iwOI7BfG2KJkoWfP0fjxJWlxtd7TCYTUF4ai/9PO5qqPJ
ChksKtvgi3kzCuKitPwOuQSddJjd7s+5PFHxM5eVp67xZqYoXY48q88z+L+DHMpK
MOGkMumW/iVGIAdYyMD4Mocvgz5Rp4kX9sArCjxwW+bAb9jNvv5n8Igv8CEr4mf3
vIinn1+Fh0jxTOnlDwPZz+MeJM5R8PPL/P+9nPc8ZGDmrlZdo8NeMZztvRM8b2vX
qPTTSi9gRb3TTDC7LHIs+apTXIxwbMotoiprYjjanP5bj3MnEKkR2fLOCVC5dQ84
DdtiGXoOLpP3JuR/7hb/cLTYK8QB9dqoLiGMX+8eFYo++P0v0+5Gq8kKQcILcIaF
ay6W/l1JXARPenlN5znVKRIXWbALzAUy3x/Z+RY0D5wnnVo/B6py2rzjQAEoYGwE
0h8eQEo/CvOoZPOoiXpnOyWFjxOEjLSY8geW96L0wMHsc3PSDxNInYPX1b6xXPBp
iiUcYIGuOPesJp2zyThfkGhbbPVP+MDG6sGENyxnDn+6cau7qDA7qmdZwIIwmMjD
t2vNNCPqHYpIVWH3wqBN9md0q587RLCzzMlKO3UQrr/C2ULvtgOwB7BNWLVBaama
gxBBJGiyQVALuwtej9sRASPPFbobXOmrrqZHgGt1EGh1J/nlVjVTZaU5QXrgeeXF
CqdgLYwtWx9iRVtWgzllzsY8ol7Bm0QEV8jmy3D7NzOoqIuDrAf25QfO2eoxQDEd
ckzhhbJdq8OdP9sdDQ0ha/ynv/xFFcFtfNwLUs+6Z0JS3Y/fNqvvl7ZvWFFZPtw3
JKarEiRSsyUdhNbDaKhmuFpgcMeEBDAqOiAv/yHQKbNszeuQvmJf8vyCiOPwmlxQ
ysYKK59/WJNKUQ918G8gWrjQN1Ey0DFF79aj+rawu+1SuywkUoQsBqTdNEqxjyAC
b38Z9cPfgsOSL+E1C8d68HXgDZD4gqJOBtBZc7jrMNKQDBaA7wnEWd7P9Xiid0m1
jrtHR4mjWsXtSyYxCEBGNXsutop71Efmxz7FPUBmH1hP3gyFBAqifX94ocJByOMc
JJY5k4AAzK+kWs6NDTRmDFuj+V/I0iY42gGkHMJBqz/tgC6j6a7dHGKhQ9a0J46h
HXrC9oCXEJmeEw0fiQ6It0jDA8GrSzSVgU4GQGAZrsXpXE16wqZR+ahOdcp1J5td
rgQ0SvQNLv0qAl1kPREv4F/B55+LiNtrDrgK6XfOTh5m/4YEU+bNchDtryMqXSUY
ZulsObmhn0LLv9dSObfCyTQxRyfLBTHO/d//TwC05C+RmqGv0rkId/BJ09NdsfxE
DZb9pXejB+3RAcJ12jt1UrisTVNvOfnrYJZvEtl11ZEVSBbHjYbQvkGkxCsFo3C8
R27e6YBdTSY5TCEkS3zp01p9jP6OuARaPlrOjaePtudhthRqliRI8SG41jHlZ7AR
FKkvTSg6GgMyxTy3PllLD/83rk75G9LvzY4WmO0VlKBbG9lQYWPOapq5Z6KteTgT
y6H+LTRnsL2dhRObrEyyj0xGAfEeNwZs7xYwdaEBfgqBkE/vyDldTTvbMTcuawbZ
+X5dxINfKjCeuKC+auoLXhB7aHNdnfP0t7GJ6qx41j6PuzYVg9iztb8DE0POzTzi
TDDD8URdLUp0X7flZhXr7EQrVsemXZMZgieSDWqnazsfhzXVBQad15Omze3G66Aw
qG7oA7UtEkMZ43ZGLsy99RDRAzGqAnn+YKr/Pcpzv6nYXzVFM+N3QgU75eOP89YF
ZjKVgQ8ZRyOxTvQR5zGerlovvWkGM5NYlzViwkCsHZBmIrk0MAU0FsPv9q3bvOK+
lbNWvfmYgYmoifCULtkON5JTyXEQQowZmDqJFWjfcewpVGuj7UmhpaD2Z2rcvwUm
Tu3FKOnZu5XqSAsdZzAuU+DKbw8hzw0VSVi59Z4hIiSA9EqZvuX6WvoVuDM8PO1t
qlfssPebw9NQEuWaPKxg0xDEXpXT7BaCTPObsbPuEXrhU8yJL1R+5HS3qFqmPvX5
cNEjwdFT6qLpnIasJXMATR31NaAvk0CAWJw5HjBQ4r1DlfKKKNsEgfEYKijzqJXF
2qkFdNpwpTEjrjvaFXzEzlQ4SwM1UrDIVr3uLDKRlAkdgvfWiigPN1XDhHEQm16J
xMMzCNBV1a8F5eFHjyw77ayARTZ8S1/KWa9otFfZzzsg9g5nh3tz8teORfvhKR18
GNNlU1oVlW4RuAIhDdF9nIX1kZTxCAbxW5zHtQasZ1nPasCDuG6SQ8KjHBn2giaD
GM1i1LYqaHaHdn6fFE2HtQz5U+WxzrYy/7dPwbK5pkj6qUiw/I1k1My8WSr6MLFW
AkbcK+6LgwTHJU8+5H3NibesxhJGjYNjDlUhVOhs8aRYmgThhHBjQhvVJJUaf0nJ
r/M6qBh0G3ZL+Q450KWh3rAHZuxmjtagoYRJm1mT7q3JLMHXS+NRKTqN4TrC3RWt
seznzHfh37fV0L5TCEevJcO6rHnHLDaOdpgl7fs7EKAeh9FJ+0nzHMWbI+JPDApX
kJPbhAJEq/cel95xWyE0Mm064fQTDrL6ZKGqNr4pi1wV7K5WQScPhcUtxHJN/tvX
OXxDPJzcl1Z3QUSdKgckot/Dk5OklLeaF46/YGrU/ZBOHb1ugrHNjofO7Yb8DT8L
gL6N0S+JiazugDoIq61fM8jysgH/O9qbv5IfyKaPtp5IvDpvElyKim1A0Lt5dQPP
EblexE9WLiR1zHIdcSwSypcbkNM1QPufvmwbiTDv067WB3FrqF1Q0HGBj484+d8c
4yTYqa52LzaPReAG69CW9k5RAVm+9SkS/z2WW+bhn1SjBli7lf2kdGrMTzXhU1Al
foxJCVS/n3K8VEWZmmxIO+MwrkOz7O5tRNn7D08y0d8+k7CFfcTAFs1PWB8p9cLF
BhdzRehVOueRqFNtW/Udabjm0I/WD7aL2cEk2/A74Kr8L9CNyCaCDPgqO9IckaLl
jHYPVvdRuMKT6cerJFlNp3TTqMQDFcLkR1LZm0mm1ptpRwuSQu/wyFgphMcwx7gz
ia25svKchTq4pQOFeXKodXZS7kmQsmZNAwJZxA2e7wlMbmryBeghj3AdzfXqkCZD
t3qif5OzBjGI6rO0CfyUMnd02mdwUyZFEfNy7xOg3K9h2x+QHO3P3MKAhf4bgI9F
d+Irr2Od9R1BLazukgm8Nb+9yilcHiqg2Bt3jvbe/NHLb1oN7bb9z5uSRoVQQdeQ
GcksBuusPeteF/Xyfz4ZOKVm/JrjIzE1OE39OSqDpwKVtSYS1YoLV1g/TKSWh6CW
G5nFOcHBkdr+JlCNqoa+fWRldfj7uQlf/otG749T4MHFSrZvtWVJcg8bl82HJ30J
iqSZYXoeERGvUHsZNi49LLoVSEm7WBkbawkEggpCwKDvvxSHSeWlpjJZalgA4V5a
ZqvpiIL3RO1NXiHQoSL73xotDf01qHOlyJZdrfBZGDscMRVg+zHr7T655o/1C4KA
5o1ZLi/waB9fGhquUyP6EJlwXI+/nk067KXiFwb1r8h9sPXiOh5toMkp9Wrj6UbE
Ni/ygJcAoveH/ubc03ZqyjA96gUCLERWOHkD3XRFS0AARUBhrYPV8K4QKk6Zffer
4RGu8PQ27EjHOZ1D0Lg/1EOb9qZTFcWMHWePyP5t43YwW9uba7Hi7wIVDRA5wGac
+sn58wQWTQld+HFh3HVg7MUQakx93a5qAjpWOZeLHZaMOscI78ME9Hqdn/y5euTU
Oiw0tqkIXox+L0Q17jAh4h1iETQmzdgMnXVu/OmDmdtuEpfqCNJtazsR2zPbGD9M
3N/YyIKl9girU1IanMdnuihaOn55MwEkjdTerv2WbAyWfyVJE8Y836SXDVWpnhh/
xPGOipAw4t5sEt5x61Ny3i8D7kHmdtPydxyLJPKlcPCconRHI/mCqqYY6wwmCZ0W
FVzQ7rbO0BOlYZN3TikgIJE4iyZsSFF6bYEFcOWT1MO1qzJy3vVmLexKgW62lLtz
v7oTpKZuEydmd6d3K0iHpYuhqYjKsgVnsK5pfQ2HF/CtwBEtr5grvN7bgx8SYJCc
F/CuYtv8bS6xUuDzTSq/C+ejLT0zoLz2SED2z4aOqL4ExK3win5ro7YEvqfMbzPz
3ZuTVCdrNBlG+cwVWkEsRY0tkn3awTEjdwZWxThP2HFE1zMbSAocPWkAx4Yti+eL
KXumydR9ydKEYY+egU5gLv9+T1cUGkQAJg4fc1w4vRQVoRExkDc1XcAHFwm0mq8z
SpEvi/c+RurbGO0Jqik5dEYTQYhK8yFfRMXHofgS7c4GjwgyAImL1LqHjFc9yNfa
vlg6k3TbcQJhIzZ+1z2efTOGEEoKajHxDLHr3m6sU/3gw6kesKASbBPg4LOeEbBp
l14IVDc7Giyutltlt6kBoPtqycjCjWlYrYDwlMVamOas1orZ776LMyc4wKChkfMK
mpdV8q+vStA9MJ6KFPuV0NSYA93fG0FrsS4CEqKWJgtH9wizNfQpftgYd5cYRVyu
rAJ1qJDa1iRzdWkGnBFlSgsAXdBC6RoUzvJ+6hV/j4A/cwJvmkPMcllk1NJGJ4pb
7AX9ABcy9lvxGfb1HcWqb557x+Dmoqwlc/pvyXNFelzH36A31QcgzgHmhKHgHJ+C
m5UBYTQAb5hK6i9MQVR2gocDPY0p7FAE7wcipTlSGhGJSR7jtIszPTy3BSw2lW2p
SKoG9r6SQlI7ycQwoxFeivGCn/9PK9MTBlhIAVUpabqGvXHSyF67lSLl24Z0uh3B
yrUXv/H9EjEPTfMV8wgLaICJK2+H5bHilyLuPcUZ2bc6KJ+UYE7oD05uR+VhIyjQ
WYmNJPkCDZKuYH0gPqiTHoER4EriysfPA3KjG1cqDiGotNupH6Jg6brXJns/oN12
wvQeF37gn1mSXtBHLGiFY6ttMeAiMHufHvqXIbEcK6PJicTvX76py0FNs9Lfojzo
sacfDD1hSCdlZvMuB8FxJ5b3uTh5VYy+XtwlNP21OqYNsaSIHUj7MwwBzDSbS08o
xJsrk9OyPmpM7g93LxBIkymArqMv+BGxqOFkm8bjKxESQLQiZ39tyj6ipN97four
SrH/qG67D6WAfcH0hFl9HZJ83glHWDNlDQ12N1m9+FVPLIQ6DMoj89MC8hfh0QKs
osw0TMEB0vUOE78bzM8u3RoDMUjkmfMDF1SsrtpDQXGwl3AQAGlV5FfZMhTjuC2n
SfqvqYwA1rP75s+AUlsCnMz1t6FNluOmFilnLxh32IlVKwo6lq93WeE9Bh07Li6y
677T4hX/ZdrkrsciXaxFUhmR+EEwuJo4IVSaOU5kTu0aIl+nOc4f7TF6MVJw/hUG
gEG7IOF8oUvQ58FdEoIVdrI9DAvfgsJl3ZBznQz7BfxiyFZlWDcSjsvTusFydZf1
4KjJrSSuuZK86KCnNJZ3JgdUEN3HzaFL0MG4xhBFlX3BH9oPVUKlyt6LyZnYmU3E
z5JMr/Z6QAB1v7IqiYkPurrJdkFxwjvF1gaMn/G0lr5MlnS+y3iFgxoIsLmkzkpv
ppIeBsBz8JJu5AeTSOATlmAsDEXFrZrdjOz/Zjwp7tPjkRZbC71hJzwGfwoPb9fD
7Vm9EDa3VFgC1v659izTO13IhwP7BE3xhQanLwex4bL5Xw46HsYCEHYe3KFUvBB+
zXXLM712QbWCI0MU+llIS3509rjDV/RhaFNJYniJ0MrUuK6TwnB6yvYmVSeqsXQI
NkSP3aM4sBP/ftz0IlWRVJS+lUt4OWgXot98O8RDRvsq2ci9q0YoJW+sZHimC1Pt
zGHwsDr8Cjh5cHXcpVEKWS+4rSCjpQZ19VQY7eZslR80hwmE8cIQgQwTI7H8fC22
zDMKWsQ7Ixk2gRQDU1BtQ13dO9I5R5hLpJgbD9FRZexfknDlu4hFSUBKMYmJUnAA
sihIthwQOZ1CHsyfccYXBAC8OGhT95dIYPfEZ/4OkMpfuC05eA6VhHSx4NoNIg41
jUDyLdNh+q5h/0grgq1Tk3hrLzu6g52cpzxwGLB34r2HlvAt0zg4Hy6S27/FGYdw
cdRDPsjuoulJK6WOTgeWF4RC7q3TlUaKyo5ajSE6q03QcYca1dj68Ne2ERklqO7A
PKcBSZcJXiSnnlplaK7k1xPwgW6Vv80JZ5HAqRfJlcI1Z+duTtIxqZ9IhjnnV9Aj
Mf0CKysilxsTBfixktLQnrag3pzReW8PCPBPW4GrH+b3LpriykJQN5/oPDaItINu
PTLfD33rih0ictNU05OLajoCvFXtmxOcSQ2OBqqYOjfpQcfpN8EOT7uV72PSuljW
SQ8va5r+p4is0dGHkJYzNJ7yoG2P3nhclL/YxawReXGZSn0xXFkj32PDv2zB+z/p
Ldo/7DkXqrT6MlCk3wjT9yas1E6Q6Kq20GmZY/A7vGkHp8tE9fGWozjgQGk6GCHY
edgeWyVv/jH0FkikOnWn1fDwnJjaawYlIwFcG3h3ghEv7R4a3vKEYUsgGs8tH7fF
V1nOlPTQ40ZTQrtCuulDe3gYWzD9MFJXxDIh+jbNIDV9+ubyCKZtHcg2g2bZkhcy
612QO12kkn+L+bvod5SuIJIsr52HncrLjqoe1g7wBuUaYVP45j1C5h9VE8/v2z2R
eFtsQ0vzgMzKc/WKAZz+H6+3O9B9Wa9XsTU2kp2JCVIevImcA3m+WW67U/+ZPs1k
FZIgAx39sVbKO9aGwVEuZmsdyWXk5V+hJ3oDTOruttwt8DzNl+x4RcUMtJLfRxNd
Xf6MVg0sWcDxCIZoUOt7jgPmgrBoZCtYA1IlUmPjPQKh9aDgxEyv8dZ4TZTXbPR3
Z3mqehaeMtXWxt5SVFz7KwI4/5JiW8iFCSeMpKrOruQUuR4MDTFfEpZfNQm54Rp1
bgpspOzCIUylkCd+A1ihdE4yF27uh4REbq55t3N7dytv8V2A+m6z+/AHeGpgN0Ju
80xMMskj5KJt2vTVAHxs2aiKSE7p9TCB17fZOqppMhWT9fgUF02Ko5snrEG2hr3H
j6sF6Tn6rRI90RyMj5chl+dV7g+i3/jZ3+HXq10u2L8SmvD3MQXSpYZPnWtbr6X3
LnuuJn/A0Qf4rXP+YCkGj6LGcKU21mqN2FgnI/Z6lSBr1oj9FF9LsVpn+7nMd82I
sI8i1izRk6DnzbfWVmE5SX2Vmu+Llr7ZfeBB+dJKxERNPvSVWFO6NKnuy5lKbhie
Nafr+GS8/HDi81RYquyKDhdCjvaCuSbK85Vfp99EcXuJ3aGWb1yAJhfEGKFcx4o4
aV//aLFNtKcfIoqEGFY4DqKOCxULVxxFbAchh4ZGU9SaUf+H4UYjHpAdiP8CjKLL
2p4531DpiH+OYSLIkSNX0KkAZbf4pUDz21Jf2BYj7sIhCjIYe0MGvecJFUnELuvr
nEjEJ23fY/ACUAXRka8CSwMTcPbcGSZisFJ0U+iHX3Tk/KUSK19vFu3kN5mxN/qw
dH/sE0TZ0L5WO7eXB+H96B0fkHDlZ/AuxILv2PL8p0rqEldVt5yZf9nBp3KQR8KC
J2VaiB9cvVyu0hARDb2TCYOgk12+QR6PjYiS5A1A2TcDq3pxylgC8X46aNJeR2iE
1cm2m6x31OjVqJjRMCSAwiLTHLZR6t53jfnEyvfNi46Bt7UJlLahQXptGKhyPVyS
KjVPfSs6uc8xj2kdplLAChyMtYbDPoJGf3eGm2c4JxhvnQYg9Y5Ckso/aWRb3v3w
SUfZkT3oQon8TXmKgAosxBuPYGyqcB4PjQ+zOdErau14Y4ajBZwGMtttBBjvjyg7
K4YnqDOo5UCytRFIsdug/89OEmumcXptUY1ytsDLmjTCoEJVjuaseytOyiptAHiJ
yM5auxSVY9vjfGfAffJsp8FTBNgfmFZoffCyKsGazcNsZVeDPQPcacoSAdrW+zuy
OOQCPuvyinO/64rQnznU0cdYTLDbaTtmediVic5P3jvGAfr95q9NDvQ6SWgOKocq
Ha3CCqx7W/0dIXzQ7UvK9dFzMbi/qqmEKIVvB6Oe38zvacgiW61CIIug2VCuqR0e
jwQafE+ClawDv42CNawOZfsnS06QeMpnl3fKBfk1KvWU0X3LE2yJIyIAefouX/Ds
sk/+K07drV1E++usYZaR5ZyeUygoUfEIHDVBLvLEJfru4GBNAV7BePPjlnV9RxRF
764xqxZuDk2o37fTH9p519irASWHI6a3a+biGtprzdF0usY+dV22B/CnQbEytFkt
3rI0M8c5JKiemWRzhm2q6wXuPZLV6l4C9Vo5STAsUUd4U/f79a8A+nUDkio39qWr
sglz6oomyjjIPDZeZ9Txw22vuujBATu8jrLt6SPH+EgEnwx9IMtWHIealHkYIMWX
8lFLJe9+zehGffASXheSrtqgWwnNHeppo61eHEH6uEm2WbootHnbZtZuQO7aJ0Xk
1KErPREUMAVT6VyGFINK1BPB4hhKjUu7qdr7bnkTSN2Phn1acQW4a6zVkDxvSw9i
KsQuOYTps13U+r9Qc1MidP7qz6bidXGCFP9wR05g5OedjUapWIY4LOiQoVzfIkjY
IqIGUd7Wjk5Ynx1qRzYcFlH+kyykhsmnDe7MEiG+hfhvUDdyQHOcickITSwd8lPV
6c0lPgfDY4nPEyUZ6kekk1TN4NFuyIuQOFgYJNEyZs0Y5oji8MIdzEoysr70iR9f
/LBRqT9RvFR9hyJ2oT7OroVHIjiEZNHmyYMTM37ca1KfLGkFmZ0JgapMQmNR5KXP
Ny/lS6tBKJe8/g4S/KpWI1SOuiDiYGCrnjbYusreGvVEHIyRdIrkh4wn2xwAeDo7
KYMyd4xf8YyGVp3auvMisvwlG+5Nubx9E7/WRHboaBKOCh7yhIm9aX+dNM9e3xvZ
3TIouG50l4dQM4pxqox23CNwPtinMDe/eTp63HyHyMMfK7bfsHtiUF2c4J24izWS
eZ+vYviDIOmnJR5/55JN01MZo6mbRB3/0IDmngCDEn4dQznUJngXaAkjOpCaQ4Nz
yYjPi4sENvGBi2hQiXpI/KnfUHNOaHXjVW79bf9/4MFruD+sfZqFmWOibihi4LZL
daPFXVDDNi7gCAQdPrxd/cyyI13cUSlbLmXZVcchtFC0kAi4+HLtIyCUro5mCAns
E+WJmDbsuKdePd4QP5+ncghOoJMpwnvz7s4oxlKQD4mLS4iOwZtJ/vzqCt/kqPY4
EekZmSLvzeJkP/afUaS7t8kAXhkmcJcFUFZOySM3qd9jqPVDepPIKyHZXci/m+6k
Xf2yVsLfNR7/Q4OPdcGtn3k0TGCwv2DCNjm3T+SJEhRQyVN+HEORG94bZPLfFsWM
u4SVwTgdOSRAdHf0fSY14h6HJllXtV2OcY1QKjzZKnupebB/0LJibTL1rZlOHHz1
FYV/gpdPfMbJ2RmBhRkakZxm4LBY8mqj0kGDusldN5UjoU9XPF3mryUncX8cMvr5
w0Th8r202O6taAMyConAQTQuf6xj6PwJ+aFYaKGb7M4OLyMGad8YESeiCBaIbGdW
pZtL3xRS6ZkjvL0NjEnlJNlXfuufaOoslAkZJuuhz227Xir2Qj9wntXvfDZlmNMk
xs3BgmBneIs+9zqHF0suPVcr8U7BsVzIT8Gu2d2rDXEGMFYOz5LtsK1vybRjS5Xy
iZ8hkxI/60Xu/OJkWPTuLteWaJId7FeXuWYg7hL3vLobA5539ZZLgWx78C8bbbp/
x4A7osBZVwDbH7iogdOUxB+sEkf2Hr7XJmOsMUPQuUChM24mLlFm181yuWqJwjYa
QcKZ1n8oLkIkOerke/voxAa6BAxK8HcSLc7XTknfu64GBIItA+PLilADWgw3tEGJ
ovXt2GC1404ZnwPJCNcU1AHB75/PmO0/nY/l0DIzcwv9S+puD4Wfs9UcSL/6XfqG
ScWackCpjdy0H9GH036dxpAwZiBHXINU1q5CHR5tlt3rTnQ7fKjEo5WBKUi9C5By
xxr7lY7vVcrF9CIMuqaifVN0gdXAt2GDJilIzmhrWc2iMml9DADZOd8tyHL4U/Ff
eP9NW5vi+RUnTy0+Q3+d7/qJiDQHpOXYEQZB3Inx+i3OUkxBO1U4NGls5YaZA4DE
pBliJkg/R0WfofAxJxLjkoquCF+OccMZGy9sXG7CC3cUIDwFeeAb30qb9LcfkNrh
M56apTkrE0ezx9UvsWYBb/ubAYgEctSPqkZ3SGD1vNvHtXSyWm26r1Kr9mJCqawM
9NGSZ4OF/TrW718jErCZkAcPpmzxOXH+BspiUeUNOUXJxpg69C/cqwtwtA0Y+VJp
IpsWtdGWlOAUOy61PF8JqmVbDM9dM9a3AuoutCvHOZP3WM4CtTLyDh71n86eElGL
BVjeuOSQdd11TIMcYGoEvND4BR3N3MkAhDKdK1dl2WJZGPsLFOeQQpOD+5h/jC0s
AqGjzoxU7SmEJYvtJZEkZpfio3g/ok0Vy+o3ld31p3rsw6Wk0yGkkfO2mvc2t39Q
+h0naV9unVHLHZ5a819ytE31JLUGEX3ASEXQde6/49gQor2CRcw08pn7Pvp9OAb3
NUvy+XJdd+9Eazi3HL79DJ57CwieThjmzT5bIvM04GyWW5636tGCkq0Eln1AkNCt
0WdjuurQrWazLSZWToB/PBqI59LrGBv/9mP+GWY/+HKd3unjx9r+SPiQhpCl0H3P
3vFOdn+kcjYtjntZyWfYfftKxbYYUNm4lVfTwttdqOMJSssj/H+h0fAeQjC8ojFS
r8HuaHKeUF3zKdL+veuRrs7sWHeiexBO44CdbGOmTpH0QUFCV7jCckqD6aJrLJni
TE7UWf7f3UHHpK3TqGPLgpvmjRQKktDPbrSkb4xodWDdwTLVrcqu/GRiGjrkDdIw
kJGJ4my7Rniyci39QGDukslrNrh2lg/541xLLNow2YA2aDBgZa8wU4jbAt/AvLU2
X5XCpPjnt/Yz/Ie83dFSL0XlERdeuhL3tlJ0Y0ou8tIYrCFvTagXcmASHLEkuATV
K+etFf4Y+0K9QLtnd1tAgRUNs8weKDpTgNit73t/OHWGNZD7QRB1p8j/xXWEalVQ
ycTIMB/W02YTXK1edV1JazQm1ji0RqO5365NxN6HSLzII9L7vEptSfQ+H9fujW0y
ddQEZ1kq6LJsdvoWQpSPfUV0EHffs8+mOeGRs8AYdnaSKdHYDzzj+d/wY0RCY0Nb
MFmk+myE2OyOWH8Y4SvCbkdb4sMDHxggRrJfYWggXNXPQmfAX2Ta2ZJMh8JrAvmP
Rk/jPawmuRSZs0Xe1+U7qTLzn1na1Q6sXnIfq+GmUlj/zN4NWrnPYtCDUv5Uenub
QZxc+nPH4pLJEziLPyC3UcpgHqio3ErAv+2Od9vTqSNJyRwBGn+xa0lzU+kLHfQa
DBGZ4a5YSLJ5URUWkEx1oJGOsCk/UTYaioJd59267eSRec2hPUYsVfpNy7R2I/3G
smiYEXNteAmNhr9bL0XITupcfNfPS+pyF775k2vXGNHy/Ug6jZDd91IMn7VWfanY
k1o9X/H2JfW0UfGksUyp8kTeli7Uhz9TnJZHJnNXKotGp+AfWeadwfx24HOKnwH1
LXcOScLBeCwun3FkRehG1YDP50oiv+S853m9sw1XHXyPsftHNkucJBZ6ZBz9fmsZ
ZTO5aQH4423xKTRwI79X/0j+5Rd6/P1kCCp3Bp0djMhjoL7WaBGLJo3Pi53P9iYP
4E75O32uYJ7Ou+RzyarrZDChdvCn8d2+8enIZGqRu+IiZMY6BRNi6l+kZDjQ2Lqx
Bpbzw74kDxz9hK77aWP7em5aFORNrDCLA+1iUDIehatVHTzxqgvCxamkQTb1tbE6
iAP7M5HHqCU3X3XwZAJUp9cp8dNHkbZpDx5b6e78XQjfT2EKKMVFureYGCABKz3U
qwzuDxePUMiMix/1O15H4qs7+SYdduOe+rM55IVgCfDWhC9dTJKK8Bq0MONOeIVF
xh1E3Y82CQHMv0toZ8RbH+MbBleET6Z5ZOEtmDUDPwsDNWbYwGzEVOf8S1Ff9HVi
X2exGTkEBm6WDpucHgAU9KFfHNf0+GbeKfCxGQeupf/QedPFFYK9wNILb0P51Ubw
uDfs1tWAF7bU01X0WOf8Dk22PtzqF/At8g7q5q45M9mvsLzXDMnp+ZezY7dooxH3
4HLRPBkbE8ZLYlPUy4TkW6yP1JUcHHCHtvCFRGk8ICU30S219e9zUjo+nQVvQiDD
oFw7LNuNMAgmdYxaiT1tMDX7/yUnF1H1NYi68dC30te3oNykWSUoxMUMqCJmLoob
TLmcKGAhrDc1YE1x8kWYT8NRNgrGR9EJvXKg+bpO8tOjGmTo4ACtF0oElMXkT3UH
8BM/iTPE0yVeZ5iE/sgj7N7dXecHurKZq5I54OBe8AZfP7e/Un0vX3Dq7cRfjVGb
1wynnSVh0rs+Ds2RDKeme78iUDUJkyh4DP5V+JFluWyzqD06y0V45jZyL2jey7y6
x3vV5bi+WC4rF8he/F80W7F9K4EOs9vvqLqiJuhAMvMVu78hit04YfKvF9K4KDC2
5LN3sRI1K5hiQeXHY8Xa/jDGeMD8OfUZBj58NAum/d0UUkSE0daTc/LXJhg4QlGB
3sdUWoFyHxomG20Qb3RYBZ6F7ha0+RGOs6Ve5zEGFdj2wWfCSMpJ7+F5YtbW5i4l
hNCjg8UbIEzbHcMDZch3xjqGQki4Q03uVq+ExCBwi5YJdLZLBEIwINZJ7ApIEQsE
+Bxp6ff2Y4byf4HbvMBjCKE8ZuGAsK4X4TxKtqfqtR8brTUhY/kH24W0Jl6I00oK
qjY24W7gVQpmSYAc9b07bSe30OEKGq4fUdIxs58hi4uH4rEzTxqZCF7j7/yDmicA
z6krk+XhPsS5kqrTnvD1kM3B5HMJLKsjMAMkU7Up90lmQDaGDyViz6rO+AIrFF9K
PWAJ8EUy5tuJ9ANlBH6IlzYmVQ/8yt9n/j8IiLmxl6xTeXvTwqBp5q3O3sdYy3CC
wdEfabXmP7h9uwzX8biilagxh6axydHO0gSJngqcn8FT1eHhyeQECEYuUUmHiBgL
TYY3HZjD1d7kThvlibrbxE1SslI6bbo85j4hLh3XWVmNC40FRvAQ8Qd7ZfhosJnt
76TVI+iYrn2o/f67IubFsbLw0kr5nfnNMeRyEbHIUeKRNhXoX1Qa9S/TKCRUMa0N
QzZpXoQ3kcgj7rW9jZxBRCsDeJojWBqjkIOO2eQ9Qvvly97TJiLzUZPxKk0Kfc+H
VkjWzA2zL4kv00HqHgxGz1NCFzWQga5N6IjY06QAoIXupvJHeB7086urnT+S5zM5
hHYe9F4C7xDo48J/TqjeS0BBTGGSajRiBLAoHKx3pt2aOIcP2jyRcQQX7n7/AygB
CkNS7cw+Cbkv6vdNCrNFs4qPBaBaBxrnEyuWe083LXiRQ9oOnzCfIy/3OAsE60P5
KE3oGkQUxLSdvxE0YA5Bh8DJjw50m5E1M8Y8cxcmbJKTwyng/pdqt2U5GV2wimfl
duZW27Dr5CjcI6hErWVGuLdDRf4QfEJSZKUbdZko2kx0HRkxUfRaPsNc73sDDaVB
N28+5sTpUg1WVXUcqWagDCb9aElJfObMwTBIufNHNO7MFj0nUlFALti68EEvL4gk
oRr5v7ZG+SRJ3fJM8N0OFRHlq85B+w0iti3Y407frYrU1UJcUbVI51rC2dmf08Cn
e2ZvwwlxWKLsjuwBcNTzEeJmY3EYejuOXvMY3FGic1jbKQ4cLVJYoyxyijXcELGH
ejv5+I9JbgvXwF8+bQD9royHaQg+S+FuAEKwkJ9QsLi4zDtWpNme+p+aECm+pHyO
5YopnNZXixDunsqM+uySXK8s4P7NyDuUKF3ae7WXIEc243eVPMu104MK8HZgEAa6
3eky+P/SxmfZbvYrS0p2UqV4kvJokL9DEWjmemGGEEBL86Ut3IIHKH9CgJvETaed
BBK4LHxWiiJdEDdTo7nUVJTaHfqWbGNZAqNshPBY3enB29qiiI5c5LEh/cWz7035
pGsMz6C9gQ2x0/HiN3XuXOpaUwZVbC02nMBjGNmKNreSZyWZKNp1GStgFDEd6XT8
892356rTHh8wpzMRx57ANm243eyNc4rhfSG9ywdqU4qDtnEgkAyovF5YlZhc5Xy7
Z1zNbpSojf2jMTEXpvB+BpBrn3LwG2mi7NDZY8Zc5vdlrISLx48zRri0Yne2rKxr
HRIVNDXKXHl+mLxRiqL4ysOdwZ7Rszzi1S6A89drjR085m7CW3CPpSGsAheWY3Vu
Gwq3ZlxmuR8mLJiChyfEmW/QCDHaDtzn7QDGKJ1SQ/JBqCuyqLuOrjUc0K2FIUgp
xr0+fg9wfY713JXxtW0iK3jNR/BbpIjBtS7/mAQerTm0xiZSAZtoDgf4u2Rni2Js
uzw9Z86eiZeUh5VmpY8U17fmIjXLO2Wvx5K7nAHShlvrVLKXohqTyEgy3mXzHxl3
5Mtbn1UBRdtCzVM7EnlaRCEy01YouqoD4aCoissKiV4fMFlnuEFaxyDjRHZ7MnnB
iOhOZghHeIRQr2TIXP/ldRoFsCk+M1LRpp+R83PZ/pdNQdy3KBuOCZFh9LoA22AY
jj3vF4xq9kTXBDChIEj21x4n3ciyf1tYrm/7+o9Wy4lLSky4EGjYoxMibPv01vfm
it79Je+QCSMzkNoDdM+p2Gyy/wMtVTmehF1RJEuxLHLseS0qBug0OmAWXUuy8AxK
1Oyl8iQPFjm1je7hAWKhhUpfpZUdrQuAxq362QhA9Ec7UzDNpm4t1EyXVh+0kunt
t2YXjg5FyA3yZaKajHYx02VdofVdCS8aMmnOYIZHgMSMLKLQUR2W1sKCFmHEYAiz
obEZWr5RKsPM9nFLc7NpNjrRxU4QcggcQvOiW7vo1Qsg0D7NPWo0UqrLrBwnFT6P
smkbYEA0QNi6eQSi5HuLWABQO9T5Xu/YUc1Z6iW19S0QIjATj4obNhzzscTFN7gH
/5geU9IX7EZ+4sPhrunfD93/QlWAxrrAi42i36Dw+OunsK6Y2mEsrgAuz4RJaMLR
gR5nmM6fU52JYxVsCRnrIV80D2DTDpLXcL4ZmoZ/Syk+1lNda/zFQ6yVpn/oGho1
wgYdhsGzDQMlxjgM2KMXWJNFK2NJRia9flDutMn6ruZg9St7vDbNUpJ3qLUG1LWc
8CxnliQbVw0h7hoSFRihpMIeEXNdX9dhKQukhMeaWrrO7GMBJXrSgoLkQvyoZJjk
LOc/0Sp3MO1LoR3VdYmCBENV+iH/XRL/o401xOvP6LDS4HmLYc93DAhAgUvPIdwb
N80ui7tNs4xD0DhoS2k0NDH/Pf5rGXBaqVYWdXBmON8EMs6HiH0CkBFt6mJtyJyG
hc5qIi7xJXkggurx4Rh8/YYQAqeeECtRR+i5/tQLowdrbIYAfxSN5gS0zOcBJMLa
fUZklS3pGF4cDQvKX/3hdTk3rYhRX2cNoDpTP2j0GEKCFC9juvdvNYrSSsVhItAW
dXYtf6kSnCfq6HISolM9uuLVxV5pFYXpkgTXOuFnr8jHDjiqvvC9vJDjlmTUUawe
85S0C4yI4NurfYVUdAufBQM3a4+2R3RYcyqWxTdtBygUMPiHjAyc3KkUgSfQv8h8
hiZSy+D4elnG8XOhD9pPgqoHTCmcCcYmZ1+2H5nfBlaXDEvxGNEIFOHlKNHxIYlN
PsVjPJqJaKAO0xvkT/vm15JWJvU+E/defYn2oacLqZfYLcz0RAo/OpoRDdtcijIC
XEgaugHmjuLB4m+uplBCn6EODD6Q+V3z9xQFbbNAi76bzy+FQDfq6WhMqnDS4r5v
UgMf8Cg9nI3GGfQPFuH7d7DMBR1GFfEc5dSuT/WieMfHZL4ilznDGdXH51AH/HRR
+VXRJnmIsAfIPg3vCOFsTbi5V8YN7YWijHqo+t7JlpLob+xc5EoHRj/95do4H/Pe
ux515sYkWPdTDSsC6jZXO8zjcwOFMRad9lJ5h0N7W74PNZiyU5cFwHv7wyyRLITs
lSxbeodrjpxQBlNj9DMQ+W7Jf9Q+dWSf3lEBMGOjlTa+Isy4Fu/BHMgoN3rsIuP4
C0SwGap00xaQ+a4qig5bc1P4JRq7A8saSkSNhqIn4d4dr+J+CafHRxNlMDu7Di27
JaOiiFa2vG2/TYMD/kzUpMbU/Sjp8zt0XDGPTeqW1rrEBxOmVgIUX7bKP2vOiURk
YQikA5MsMZ+kZIHv1JFNLHCgR+HjvbSHRIOfnL2ngZBmwcNFS9SuO20GCV4qdSSJ
IUN4Mtdcpc9G8U4GhoVIL6Ymn7omfMSoowhNELRc7s7gysbcW4FF2OYmyEA3tVt4
FijefhAbOegLLjm4dhGW6XPns2lD3Y07OGxy27jHAQIHVn5rO8BJXcglV7tbizLW
kdGn553xtEvGx0ghLxH0gjS5OSddY9Z1lyTLkZB//FacQ4l4AG6/atSAJqc9jQLL
LkU+M7QFELOWzDfJ6WrZIUhESa0CweEsUrTb3jmGIA2NGEu46naDvjLyO+ORVmzc
shNmfI3lqfchI2GUkjna2ue13l5yd5icFpPNBxA6clDmHX6VFcMNkmRtqOicXSXC
ddIDE+LF7Y3CLcO/vA/4nwLNs3p28Ozyqqilfs50Yx7b9lKjz0/Qo4EX647r9eGX
FviNiZ9DLyKmdyTSa2Qd1/7EJ6NzxvTsyACjYBVMk+x3Kxq6f9wvv9PMEuHaDmUT
ShZJebZ0utVDEy7+v2WDJkJPfEc/BW+lZrUma5Ve5DJ3NU8EKMo6ypxTj5hdlB58
00qrHloSCe1UH2Y9F+4+Hhs0bJDdyCCZNkOF2gzYZqHVsBrqnhmH/2QzTXCLNK12
GtSOnp9m60aZf5GQarJvDRXuxdAZsEvPTyIeMuWceIl2yUH5vCwa5tQDvrMwpPf+
Moe8KTI/prcrqJtNg/9cNvc6Aje/W9X/g0RJY5tMUhua2a868VEhx6gJcrV11ztW
b9D1sE7LjYOJzgplpN1gK2ElJayhsfrL739fIq3qsZEE4IomhymAMrFAkfplDYrk
yOjwR5vLvXYjNc6MDqfsoP3Z+A4V1gNqm6v9QMhER9rkApP6yvDhjRhwWhwc9GN/
CuU5WdX76YA6w18xxkBBGAKebMb1ZuzwJJutNH3q3ZONPXqU6TfLIQvWfLgD5IrK
zGtJxi+OU6vU3hxykrAxszgVJOt7enPUFcf+wDK1R3DJfVVY7lhAVjN6rIOPr3Ey
0/w2KAJRLPojEyzfAbKc+MXbNVcl4lViuxHaz2RsVgnMkiAhbMI/CwBf7LqMYmn8
FOonEQMv5lhSwmTgQg58gr/ilzbTREzLl24tIza6NZlkoa5GX9SGyBdgIerozr+Y
YqT0ylRMeQRbPqPYLpR1S69HM/zLbbOzcgHoUoWogby22DaetNlicUDZx0wloAn1
JirzsRleyKsBcbPbmcMstgFoC+TEQ+OGZzGJ33O5ydBrEFrWMi4rdUo5HWkZY7FA
D3yYMVUT9ixmj0PVFbFxcf8PjTkyGfvQvI77rSnDCkxjxMxGJXC8e097vCDFHoRV
YMR2pzP0UQthbEw5+hCBxlkJjAuoXIGooQ7CxxN7tzZMDu3dztp04Ld5tu3b0KxV
FFCtZib31t975uPzJRIfDdbpPfX0CQnG2kdlQv+nF5FAP+gdfjmDVJbNFb7nN733
74IdUZqspeRkq4q0OENvbRMqanwf1ShrQLb2HvMyrf1nE5SBbSFSwZ5SPMSm+Ghn
S5sn7LaljoRd/FD0kwGwGMcXowSJDIFisnxmKKl8UXVqVd/VXJc7eIV3ifxAwRBX
4mkV8nwqG+DnJz9pLn9Yd9QOiJ/MyAW0wCpKvuNrPUuDmw5tVnrIDStHJySODa9X
hmPlr03oaRU5Mq/np357w67CGQPFKWuHTJGFzNtJXBYW8bHxJmeruvY8+uFWlt48
neuapVIDcYhnp+Xn/RaLHJ2fViNKTLBJmsrhbCJZdmSG5pOjJqtbFpvPAx/cCZHg
TbJLF41WVJFr+tJUi7Hj7ZMAnoqv448yymQd1FeYRC1s0SjPdhhsGz67N45nsBQ0
XTBeALbjve3/CSLOzIjCMhWtKiNIBnM+2Rn+PvRlD6PhJhodr8K9XX1FFgFG/o6Q
ryX6QnYYdFK4RjYbc+guZs1ktTrvTOctzv3z/aDo0jE49F5F+BB1NJ2iOYsAwJmy
jN4OyEuyDMEliOBpOxHEGpKIrZAEgPShAUvo31DAkVwAl1jOWwKZfqB8BqhH0Skt
5u9bJunK4aC4QCtBUxNKm6LdLYJoIJxE7tyvxbERPUzehvxStdLKeuDgyJKUKpQU
Krth1D/dySNnT7GRjKOPPifPoAzWHlN8RCDfM2VgG+K1da4mrFDmaYPq2m/Nu461
3Fmlymt/c2DHcF+48fjAV9PP8NE5Y6566l00bjnIHzB3yJkUYKIvK0t5BApEiDdE
rJNmrw6tDAyiazM2BILHKoy8okA438WZ86JUHSX62xaMCUpJs7dWhEafh+6nU4d2
RYU5oCH2F9QGZR+VkFNyzhHNUxkLL98HvoTGet59xoD6PWZpAG07QHy5N1RfZb2D
iOgoE9ni7v+VzRZBc93sK6UPE4XMFjWGyiqMwWCkP4ajAEOdiz9tEjL4KAXlbdyU
jRs8uOd/64GRv2kYxkehLb+t4lHcAQuU3/m4kMdzAOe5K2vQAzbl/MLzgnJIMpa+
ykonK5iDx6BvQcCLWDhJvaby4sMJEULKnrENFPi/kfBMzKR76sTm9c0Oj1LRzFOw
gg7wmFmwbbX4M9hY1rALhLUjEVrFrfVe6i/AJ7VvlXPpxPaczUw70KO12iKqSGcp
XEoABS0wYbt/WJGeHnEMuVcrPyN0ktg7EvyCdAx8ioO4nMG2A5SXWZvMcI4Fvt3g
41Oi65mppLZAQk9aLl9xlQdGXgkU+oUTf8yKcQwrBZPyQaO7p8MauWVfJrc39bfQ
ProIbgp55MNq4JlFCz707+X1uw4grlbiuyPzBS7MpPjNqQ8BsuIeFB0h3PCQSKTZ
DsIFSeTvT+HGl3Bzj/JS1P4z7rVCxfGF5PqL4svisqWYV5RM10NrWmbgJin0y9vv
8X8xEZ1/heHaqg2P62wbSvVqx3yjM7f5X74VwCitkpGS7uSbmOku9ckS7YYyPXAt
lT6vE2W3TcaAlTHPLPtolGuhv3Nrb3G6dBhHs5yMnHJ0TytvmTFKAdtJ4Bg7yMae
DfPUKSZPWG3JMKa2WA/kL0rEQjZM9eUtQDy1ZBnTUXPPeOyjGaGkmf3gk+asDyII
Y1z/Zca5XikqUukLoqDxwBbnGvSEsyKq0kzvVQDSny9VCzDZGaqWj8UIAZRucJNC
SOVgP3AcZhoF8v4IquroY7ABVXjFRVescR4wDSNaoqHXO1QrYr58bF2KrKot4wig
U9PijYhBqzCq96dyC83jNadE1hbkhQj5AaqJvhV7gYiFM35fjGqwVuP2Z0S/pUKH
S0nGPh5Ig3Hq7UGwDnMLTOvTBSx6/1X68r/z1sqEP4oLxbnkp6n1wQAjsaXF8h8R
xJvmYJEfdkkA4Xne/rCNbwwVNteDLFP5Crao5JbyxqsCHRaIChnkfR0KCKRmSCew
HTn6DoN5cYBU5qI+UrSlV9bsQCrAK9IpVhDVTaFOcTZX6IcWe4fk6oGDp9OjHTZQ
0lDR/WEPEisYidVZhCg+2AocBZPgvSOUl6tfeuS5pZjFSFc5PF7HiY/bW0KrltkJ
ZlNXK+fJquy7j6rVQgJ483na/nzmbotzeTGVwsiXHpjcDtt9wQ+Z4foUPsFazY2f
IU6W5aXf2FCx3rH7Xv5kLrPQ3AUgBSIi0tr+Fu3c6UmiSUXCIg3IGnFKqxxsTFvU
KA9JP/qR3vQ7PX6qZC0gDReWQjuvS7JjSe7pRFRxCWZpldltGmZIhEIJGV6i/ImU
+wyxW0gXOxNc5m662gYB4HLvvj0T2HQdxX1yE+yIbDe/iif87Xq0ILfweQ1udtDO
iMtmBffxjVuwcwPrfSP5VlBnv2gYGBGU7aricwRlDEUAsV4KtEzPdsrrdsg4cRc8
KeD6x8D/lLcUuTgyaw5It9q7YCr4r/4X1XT4WcEtsWGSLV3YNnaQxfxXVeNxFfsV
CARwzogeVJ9Zkjw8R52Miib2mWK/Sps3/lH+hAGVi2gouKAhEoLwrbuPHr+oM8Mx
TGLn8gC72Pgh0/OlJ7rmQc94x24/QRfJENiIGk4Z5MQBofLLPfIIHY1nmyK8hWIp
vGIIxUlfC1v2bKNke16+2MQ6fXAa/HsrDgYMjh8C/gVRbrzwY+rd8D0RQf2gxt+f
QIzAObf/kIRmeiwtSObN/NF2gunJjVncWVfUCR9kl6m1TV2fmN62Hzwp/k5aBwmt
xkHz875tzSDHU+/JMS/73XAPlCtnIRXSKTjw2bvxDgNVkMn2Sx6qs03g6LdhJiFl
59Hn80OJCZv5N9Rfvrx+ZBv+p7ukryMrlFf+wWXH2zUqBlixl5Y7yh4dYQHuiN+I
Vp2s5yzKWpWtWI7kASFJqtMtyTlT9D8yy0WcDM3fBzX+RBCax0A5+Uy8dtQ8iMxl
Z+AHSHbjGrlvhXboriwB2E/q/4ZQLzj1jrdfXuMr2qB33S8JVpArOpScqhwjUmJB
M22GPbBogB3tZ7KW4ng9NNv+dwj+2fL6aexVfGybGXaY/BKEapvzIfcFU4+ei8bl
qfLimRW5oScOD4TqFBHfY6FATtH1wgjXIZ/P7KN9hqRZlolxTcSAxH4qVUCMwTFS
EQUjV1XToWVEZJgTGgdPg0HI5shkYI12WzGF4F9cea5ifhA8cCdDoRPFlGuKrZ9w
H8jcDSlsv0t5SpOuPzJiMg18F01RFP73nwZxobsUXcbz16CxjPf5ItijirQ8Hz/R
jmuZAZSDiorchfswo5eLTZGHg8SCEjeoFNqq/hQyu/FNKykfphpTs5tm9wUtF89h
ut6pSQeYTfFNBcOOb6U+8Eb8yfvIiBVeYW5ya6bNZmK+xon9iWm0sem3QmujUQGP
buONtVga0Q5i4F/mhLo5t1SnsDYiuBZ+geuVRLyTh/exP5Gkf5PhLn1nI7H/Miag
H7OfS5ZZAM/Igfg0fH2h06qUYeD9kQvbDLkS/PQyx5NlDy8L8Qc/eY/QqDY3GVFG
G938pRnUANh8JW8ZQ17eRmVHLrC0lyCtse81hlxjbfW+OavA61lvhOlrS5R5XN6+
nhmvZvhglKKFKEY+e85NybU+n01r2XMei34na9UIgYG360LwRi7dkgaI41h9YH5J
+wBqCe72Esikv6LOrJsirv72YDcCdOStYVJHrYxod5gP5ua5VPhYavTe+MBFhOWI
gEvKkt/3fEBQXV0iIVNDOSFUBG7GFsSy5z8V87QgndJjEZhdVFBmCdLFUzbTOggB
+NdA6JFJqG4sHhrJpBpvn66izzu/PX6XfLmuEf5Z0uBXk4lOSg1/IRutDuGcUPEd
mINV2i7dt6wc8f+/S7yQNu3wxvuZIgjOc8zI4UeAZfDNJzDUgOpbv5Ut9xdRzb2i
9iwVQC0qbWCbFMYnNZRqazX3G0aVhcQdrS7CzFRXMC6ZEjC8mrTu8/AASQBygfSW
Ofb7MzfAwQKpYYt+ob2vCP03z7AX9yTY/6fj6MTc0NQb1DVD/ZHhpYUkHdYOItjj
h0mtbyxsCUo+eOTrH0J6QYprHH8qVkzAk5wnRisguVbcQ2yh1nXNMvSa7Q6QMTNM
+rJbusQAHV2Rd/bVSbnMdRVmbVmtRDDWLVUkCLIECy8flmWb6oJnSYt/j9rFTQgR
ffGJIlM7MGGv6UshBsEJ6n85bsribDg8byEgWWbOGbpaRMbwvj1D4gHODr4yvL7q
iA7wDMu1y6rJeTwKPcHm9oubfIuAoqPVHTUtdDEccq/G1+oY73Ycp83b7zuXZUmR
78Ukpv5YveyznmOaThuwOrcRyvcQrhBC4YYIRFrVyYvhQT9jlZPg0eoT0JeHAvxH
E6/3x1E5g6UBTdriwgrZwmLDhbVvG9igszq5jDaf9A3duBekfEWi151MVsW3bvBv
Yk5C28usmZXDprzDEuC/w233zv2JnLn99d7jhVhHstuECkMKnN9wuvSUeVtSKaKG
psUgokyvhPz5LhX7weNJ+9cHfbbPTTE1xYkH79yQszeV7+b93Ms2KMVrnK5LsSWT
Tqux+4QAMMpMSDdTNSil9Y8RIZiG93ITJmjHApKAgt88ccGqa9C2pLc7igxzBprT
FwR1x+DdZYnH33RMItwMvyn57x8CnMY9Ray1Q3orgeFQU7TqaClwOkmBGwUfPLSU
IOsz7ihrWNQ6/HeC2mYLGQFAl2+bJZOSL1A4GfmwN53VbpHR9viTQaJWyICrYOss
ZFClxZFDl4bLO4VFhngVhm7Hwx4AdCWikLg9SWFM9k/ysW6b1NFLmK2AhDG16zLK
3vELgM33ysl6GNDYKwA30g9uU0LX57OT/g64V0TWXzOm8ww+0W/ZNe7dUoGdOuE3
c23p7NRpijt+kOzES8G1ke35n4bROyFRGx0HnvNeCI0KuR/J5u5uv40wIWpfg/fh
sPpx7S+tIAUm+6916799nwB00eHKvUdsueIm+QiPdyn6M4poaZl21jgmvaBeQZBi
Wp/vjIWM4+KbGBf3FPJNirSE1cKkbqPGUBAfq/4XG+g1BTMJgYcNrWl5AJqKNH8C
Vcz2AXy4qe3BfQPObWwlvEjX8i8iApCMtSnwAs/yIpzzZmgpR6O33LTFAbKpnFeN
KBuhBPm9irXGPL2uqIN76isFPFjZoXZg+Npcm+yoN3Lu2S5ODyabEviHNqIzZNRA
RGbj4IoI9k/gy6Qn1HDfELSQG53N7Y/6YflcJLKQaNH73QJwfC4VQCVtz7I+jqtr
8TU84dmfoe2lOHlcgIO/irNKaPOEDOy9inYLfgSSi6fXj5Nd2TMyMQSv2l4GsYpx
5PgNSeyYJqi0irSrochooL4X80YX0CM9mTRrmEK0dZqs/UAD6CGKoWjpTgSVH9Ux
kcwSntj47uT45vDOCHqjJr4Cv7Log5NotcUsIoNFbGmbuhYvnpKNXTqXd3B8EFY/
3sRmkeW2u0UiloKcsbY0MfXeAcQxznrNwPghi6PBPJ7mmAWQOEiQF07hJ3h+9ZKA
L3Nhsov4cQkA3YNZ7V5lJTDUHgv2QwleGQB/nj00cULcGz3dxuXhZlfJo+LRFLsB
38GJUcXHtQHG+Uz+YQdSS9tI9nTJpFItS4/NlLiQQyIrLZ6llQhFDyLmWFtgSB3p
V+JB06PEa1sgP7o72dYLBNyDrdqTrulOZbQh0flH/7wrHqQFW/7kSFACkzZdyd3c
QBCoR2dGrF6Omi+UXjqvRJm95EE18IP9D6b2igw9blJyO1VX3BE5MJTWb06T57Np
Sw8CbujbR0tU7y2buyAj7Yliqdhd8QtVYBOJC5iFiV7eqGgz4X2cOqam1V2osQH3
8CURhGVoh4Y7wPZq80t+8uqarh/lgBJPLiAfn/XPEVOsX7XFKjtfJSxEKYSLbZkr
ujKwMLpouvHh1LdtEfwXL/KDsEcKefYmCiS2vid8PTa0m6FJ2FKjt4HvznzCtf+M
EmGzw54hzhoI2B8LhFyHjjof9bkdUlGXU2ghIJIZOMEJixHu5XYAGq6XGTjUfTIP
zxOPHhWVZ4sHTFs+vstVyOYFElTxFVlK1gaVeQo37krpml0K2THOsGusxzBFHLVY
JPeFslg0yrs+HprN5PlXr3ipQ3yekFeMSUwYM1vcgraESqkN8HeOZOwhonKZ0mVu
18W6Zmq6fO4u58Lrqj8V7b4/7U6uGQF9r++YXCizTsHWGqYQF8yms5imL64GhOhG
4kzCMfztla8gf6+7I5CQTO5QeAkzPXYDjbGT1Fx2FWl6UF/XsUmIIoaiVMySSay+
J5KDzJWnM6Px14tvBl8pA4GqdrdtoxkgAhZNzvzSw/Rfq4oO7wvliJLn4/pI2gkQ
loB87mpxDQaBAHfqCAzCTohQaZjSU6ZjT5NPbxqc2eYeuwR7QtXjQRjOneZARYe5
6ggY/Fn0hcirVuJ3UR69bwHVefI/PDWcJHkviDMDada6fppH+Vdqg1VhnuzqO+/3
qYffiUbl/M2uwn3dciaSC/2U8J1OT0HOuBW42e8LPTOS+5yzsU2C0RcWbByffrWL
J7z1u/ff2ntlbevmrKhvvF/R0g+3NF/WD5G9hJ4gpRb0sf4nl5esKMo6p811NGmw
J7i19FOIjTDKYHPMWaSrARfNYcZP8T1mRjXNJ9XS6SGdAW5uKBUmXv5V0oEh0iSh
Xxh89wQXv0KK9Uj/X3gqQlnK4PddPQw/wpA6oaBxbmP50IeSTHmrtJr9KDdcwQMe
YAJfKEHa1ESWE9t0HuCGkHfHYO+ZhE4pei4AhxxrF6uF1ADVhew/nc5J2GJJVdSU
lhYT848Cs6vSfg0AASvwKcTPWHYz9pwFrgoUqU5nJIc+PhPiKsI45f1axKKYMWCo
lC+bf/nPtw5Gxg0Pg5hcqh0/Dr5nC4xee+TDR5/bwc76i/qblnieXvU8SG8APNPf
jjXtVvnLectbZhuspPlODOSOg4U3YH3A5owXG9vrP/TrnlhEUehDdlgvw58jIZzt
bC6mhiGzwT2SueRnokLPAByk+g/r+ZPy3N5s7zV2noiAN4HBph4r2Sgh6ZTOJ6Jh
4oBRLgKPWpSvwLJsUoMovcndv736pwZO5KC5OmUKjsEDVc+Bp2iE22S3f9aDjNCP
f4EymADfgV1gPaUS84jHj6+KHGpOswaoV+Et0lWUmc8BDSbMD/1eU7MPv8sicyo1
D281P8GwT2a206BV/e9zuFH2uMqlAKPJircFHTlBsQDZoQ5ndQVwl3VOZ21yk3mf
S32v9M9VAWT2ixl0h1DbtaxxUsZE+m1D3PN3TuTIglJJ+TvJX7AThfXo0THEdj/d
y/3KiiJfWtFLjcDQrz9GcwIkFXix0WBJO9gwbxDjs2gjLW6B+D/NTuJlEbfN3pHr
1SZVoB31nTP1VQkK3Mku+S4CHYnHvxh8CfE8lXXxcr9vfJcrU/IoZinHFqV3NPUs
yVQpfgb/9Czek+6/v6goXMbqWFNM+7lRAAuCS4r74wPxRLRfsxXFtxOQdLSqRbBI
0pUG1/pVQFjlJOYnwjDQ8/PRIDmCHRzWDLNbOrHS5INdUJQ+6T+INuxLtluPtPv3
KifUCukHrIsiwbuMkpHqaRPIsvbdCyT1J/uit1qsMlgEqbDVmKLSnmoRVFvNsyK4
gidV0Et/v/EczGiSQSEyFuUK5pkx9rsh4g3BEoyVOqIReKTIdn1s1FZQACFICpMr
mPtlcd5lDuPUWuw3i3J5jOa9R164SPDl8nKwqYqUYeO0BRER1NvUTjiX7H30CWc/
MuvOQyroey5o+hsaG0EJYiHzJlHJW4WPwl7EPCJMLCZF8aH8C7qCFQYgDv5d+SHi
xaQph/hrBsT0PuuYQfw19EPZmdncFDDszZxA1YsonAG/gktfPo0DUejjEfKkXqoy
YaWH+MQhbRdBg+G6zqoFKiaZ8RLYGKX1ZVjK3zRFtQD6DXyzNUwMUk2MCYgKGsZ/
ey0+GSei+45P+2GCobe+t0EEO7nESL6Zo87nDH3KTXb0+TBKqiA+p3mHTOCH59l9
0rLGVrQQNssv73HB134OAmclnNJrZVKdRNilNs/qaD9pW3+ra1fZXUBSK1Lk1OQP
2FxaEZgRJnlzNHoCYp5OKO4zVkrTVB/dr6fYnfN61Og2KsgJ9ew+uIosRsGDMpL3
zFanAE8dzPrGhhDf7tETE0nVWYOYKlG5rYpi+uDp2I5DAOdI3oun5+SIhrp4gaKY
ICB/s6w7A0hkvasKGvcE8y4z2wDbor2zna2eHy7SoQVhPSiyNAGRhnwcKq+6JHuM
st8JIcO/AbOSHzLEmrMmujcEFBFqdOtixfuho3r9VdCcY/vGw8sDg2VQw6ougDJg
KWdPpxz1c9D0FGUnW3cn0ByTqU0WWAnHZuxo2tuL3oN6gs2fQARle09WJzCht863
yr5g89cT/fXWkkiPKSfNAQzOv1fGfqykqWhu0lH0VlJmGTghVVg/YOvDE5CR5vaJ
g6OKqJMa0xvoWgfM1IrUrKvurbXzr82zM+PL6mpsgkkQ7EWmudmm4nRKlywwPOAs
V6J4ykkoHFmJh3V0L6EJHRWKR8gjoCxpwG0kHJqRnTs44RI+ZnrAoqOfsjcgDvuR
iCyKCCJuErSejaswVanIESasVwn6BL/pQbBEBNfpGttHIiDN581WOcE+uVzJzBwh
Vf+cKSTt2139XE/CQOeN+3T4M5/pbLjhUKaR8IEHHbi7dVjF7etGlLTiJvUWkaVw
xezvo2uI/KXG2MWJWi/buwj+GIAB05Lt2ApVYcf7g3yDcWR+rS07MyLXCSu2sDeE
iQ+i+cJvNosUWvC5e2JosCuql74sQLvGr2WQrcRAXbI1e1tO2+/fE8C5Tk4MUV3b
XpxDTTazfKlD/OktpoTigM/dYS0d+v0e5X940lSPzU2fJ6NGkw1BWGLil/svzr47
oGVN2A/wmUOsj3bV2waLjGZIlTtDn8GD7I6vbohIQZnzIUeBzmOLElW0JJjnWZ31
CeB303U5fBBQvcfIGdIkN1zQedyYLoqRV8fQ4ypzn+dhE3rDRjUNe03axqtPGdnX
fU2OaAh78HlVq9q5UaVb6eONIh9Pr7WufPZxNzWpoo4Vz6+jfq/PjpAO0bF0gXQR
ynaHc0f1QRQlPXx8gFv3DkSptRBAcnOmnyrGQ0Na/+ysMttVLkxGVvvPTTsjisDI
bnG1Em3NVuSi+nJYWV16naH/we30jzhQaONZG3BHrjCksK+axidr9LK/KHKRKDQH
zjUlxv7q47HgBCJUS+heRGN2+6Kspyvx1QdHAovqHjsE2YxjGSJ1yr+kx2s9quOE
i41r1aDgiS/xbBFubzT2R8QZyFA0JtXd1E9+p0b/PEcOgKybMoWTXGlMWhffPxMv
pHoSgy5EdcgNJe9UmabJ419qHCOdAO3aDb6gZW51m9+5QWUWuYrisSepZlp4Uhq/
vAsKDZCcwKwq26045o17+sWnRlNOBB1elJwFP0VIYgBIbjcDyRVnnSd+0Toizwdw
e6VTBr6pMCTmMRGpr4bv0rUpxQQq0Qp++ixhvzrijhz9suPXXSrFxb3gDIMZTjg4
6VWzV7OCbZfsJ0YKyIeN+aSdbmLkeB8aaTt8GP7kuZu8UlsfPivtXWotIypvKwz/
XTqa9S5wp+aRNrtKSQ89j0wSxCu+E94bOcPyKGB1AuxF/NT4FZ2gq7x/DbNC6+ky
gHHQJg51EDV3hVexsLWAr9lboG+pCsyQNQTZaLigu1whIxmbA8I9pI71s9cwsorY
S3FLcMYiM2DuIHkV7a0qc4UqabkhjmAlFO5cj3kDdKnSJCIReS59W/QeJXJne26B
/BAis78IJNg84HgO2+hAL5nW3sz5NsVR0Nygp+/6+7g6MD0jAqpdMOcWkPbf8tfp
yDBs/cq8U+QbFAPoaD1Ean9NEJOOvvzPx4PbM0zWzeBv/jLv5XyXLfaPoLuDEd+q
H/95Ilqi7Cjuxxxhwi57itNaiajy9K23JfWxLMFcV7Q+AFYPPSZwifVkJZ2VuOIt
OSbCXm+IAYlzQL7zPuihzIl9WCb/9Y8lh07zCaBfcycI0mVlba2U4ULyOHQzOvym
zfaCkKkkkfvp2xaOI1JGU4GSUr6AOiKOjYzK6uBJW8lOg/0DP8TNLwTkcIIWoPul
idTqvaGgECUifZi9PPTwLR0x86fU8CXw0KIGdypnXaG6PEMQmFuERAxdyvVCWMip
KEptXTpZMyA2BiyE9dgV3kbB3c5WaP8Y5kdzclfMMrxtfxKJdkfrV/IqT2ZLKoFF
qh01uErHplV6saxn2bhcn28n1T+Msd40KYANYSXoVDOI6/TeLODT+uoGYoVKvpcZ
H0mMeHGcTnbe4pWKzuy427q6+6GtGi+oD0yj5JYPwvlJxPE5PMPMUofw1cshZPKj
1BYtBhC+NArBM0M+2b+0uJyVQmGsP3eF9x5v9eTkNxkA8VnEysuxImgwC30pD4pb
ViE9EFf5us0Zi7nGUjwhvw6RacjELZC5JZA7s1GNyNR6vpvtnlb2dFPT/hXolkE+
nSZg5cL0s7+JKq4uKpx3HILVvU2D1psgKbvqLdGl6QxE9xQAxQmCKYesYVOMNoCn
yiTzYxbTGe8vt9wpiGggvfWjp+QdAbnx9gkzfaXTPCDNlLNsV7O0UxcFeP59v4K2
FKoWqn97jRED/Kjj+Pj6lIVMM1jtqiUrDUKgzO4Yuq2kBfNyZd3VdCt9fJJ/UtXR
obDoYFpq09k5E1lcLb6w0pvkLkJThoTCFbBJHnDMlLW5VdPJbcomIbxSEJKQwaqt
TMK2A6ZqE/4E0eiVX/67H7NGfNawGJJVXJJbaG1kTf4nYTMD9NCtC+RcTHtHUTmE
OH7yM1tg8MrC43fUupoF77ykyWHnSOIy96Dq7PLkatqj0o6K2ZcBMsa8ghSVUIuS
anWgEQIb65SKtaLIP7aaUpHH4pC8SPxfi3lmEWfEGlAm/u2BxiSfIyabdAQ9ApiM
Bgs5Fq3rgTNa9yPi2MHvFlGgQ13l89qqqwcMH0a12xpf9SfICXwH31taZC8VTcCf
8Sw/z2FIbmfHrmSoQLJ5D/eJTCFo0J4Cq07kmreD0d53AixR4ODNAVTr2iZoK8/+
BM2ejDTD39Vkc39g48GDUt/Hj+Or+no3571vAdxLohXH/KvfmnbZCJlLfDn4W0eZ
NphKN5A2txE68N9qZzeSM/KJxJ6CznESYfQi0GCbYGVCfvHK62pBG+eNqkrIXv1T
/b0Gq2EI1JqXWTOAaOIqDhgveXnzw/IFe55bWDchbiEAIZMA6O6kG8/4veXgXlyT
piy/5R5qnHAt8AU3xIcajGzmMec0jMZKz8Lt9paACHCCKn8MSueTZOCTFTpHhR0j
YzuIX28uTHwQG5aCSDTuKgVdZLR8HxcK8RgnnYH//Jdxi+NNModwobbes29AnckE
odz05mPpRW+nebOzL6ukGDSZlhXngsd7ixOGct2xE+kJCliG7MWcm1Ud0709JIzm
TRRP7QajPhSillGxP9bdYRghZBp85CFfIUHWREpSCNDiEpQiHey1+7FUd/9AwqL5
ENGiRoKnkUphbocAsI5cV/prfKsu5j/iOB12IP9A4UsvAKJTvGwfQ+f3tOk4X6JQ
uw72LmR2Sm7n57WtxZ3F0OnqfAPCKHE6MQs5XfsqHU4LudsEBuIjoXhv3AdDJwAW
dSJsm+PA6o7j5rYD51ZoZ5CTSMvDlt8PMKGxSOnLO941oeRPelf/+ZsRtdOJEIIK
DQDP/DmYpwoT4PCvMNyWEC9F3IsYpyLLMq/rNpg+rqMZDYWm0N/BbVCrL88WvWpJ
LovEjjHLpcl7EMrDvRNlOotWSmFtgZfc21ENulvHCO44Qkn2jbI4fV9/+dU96SgF
Ft32Fgca53Pf/rB5ImSgkcX/khdL4swguxnJW64NkXvTjL6m71kv5Tz/T7H7Zo1v
9ZgA6lm9g+t9fzU5zAHDsYVZ2Izh7qoUJ/9Ygslrfqtodbj5nH5dh/mq1PzecwtQ
2fOR6RrK2XIcl1zFUb9yoN0qrs4U9N3V2fckN+Oige39cQxK8rydWlJXhVrni4L1
YAfIsPGANu1Cm3K5BQ8eKch4qKw8fnUo5omWCas+NaGxGSwlxqdPkX5wPajibTLB
RmEd/MfK+4iqh3g2go2fmgn50nGaC4UnyF8JC7O9rrh3NM1PXYDgO9qS65p7BvBA
KkRooHFvS5l0ytEBMQNuOT67Q1U+PmCDq35BMU2ViUYh1sFHl+/Cr/W/DAS/4Hm6
4zH9Ot0UAa+7915ujQjxB88R+Oodqxz4mvvyb7MEWe7AilYa9Ef7/3MOqDzPQikm
QafAeACoLOgbuOC8Yk0BzXIoBUHKyyZ8MTCdZhL6iLNL6+FODe7jgZQoIW3EHnSM
p67t5aq1y1110sRf/QYvKezoksgT1vLr4AmB5wpVruizuvfnc+w8p6QAbWRsevpi
OphRby+HvYJBq0O875tzvZp9XBmKlBcamdwpFlYs7OzpA6t5W+cZrHvCU0uhSbuj
hELrIefsv9psnZIgpr0/zjj4K8NRJtHu0tUOYD5d95/hb5G32gO4s2FcTB3tV1Bd
ovJh9QeIHPAH5Lwkk247uTvGgS6ShYIroIfY7q6NNBMdAzcxc/RoDO7J+5sQQYDa
ecXTLyNYEUZfKaCBXT4D0YZjD5M3/Exl3RQp1r24p52gCqCjyuhncN1wLIjcOFwU
c4Opnt0InuAlojLeUorZMmIz0YD2u0aJy3JFZ/fqYJH1JmuDuCYlaD7GZs6VSVcn
pyguRu2jxKG7UA+3u9Hcf6lDtN7P4h3xdMdA1Ccz4XL+mWiiuduHTzmY/a8RDwj4
tnpZdZVcMRzXjeZbuSPU6GI3kC89PVaBq2sVjeQLvpRUQiEbqLQbSRz8iFqD4+s5
H99twyqKFQ63dTETu5ee0F+q+hG7CLYDyGbrg0NcUPmNPwKVP0pXwc+Nz6+VhSJV
3+AmOtxXSGWd9Zjb/Xexj2zoGlcgTkruT0WMAkApCy7JcFb7piQx/3WHeJEiUWHf
rjwUKJORgg42uqfd638cEKD18IThzNHlEQwNrJd7tqwVgEIFUDNT4X7EFESFsrtr
p2bKwM4Ln2AMdP+vEswoDVbo/3lOmeJYf9oaKNLC8Vkiv8nElG+z6VgOuWD+8Wtd
2a/goIDgkDNJlOnpQQ+9zVlB0lU4uXl1J/zBKf2F3orL8Rub3bavBWswUc/NGL8p
IzWBsJKOiboZxfgSdJmMjmBv0GljIrAKKFRo1kDe7i3GkqTz0ld/C6BABkg8HQCS
nbyNGj+7/XDEvSbmFUoZAGziq5il/R/8fWo+xNBiSGqe2mD+6OWlO5owPsgnLu5f
Yfotk0UvaMFDEy+5FyQNq5V6NyBn/eQIfsuOMxMuoSPN4w79U09RuKUkoMmnfrar
keTHZgMKAqtHjsh3WVogBNepiUJe6PDYqo55vbn3URzlqMXB3YV1fMxUhR+03R7z
7MWlgm4wWhk3jVCNxwWuOZdrWIzEO5ZPCjhKCir0GlDvs9Ev1x21zzXIl/KJiotl
CvWiPem9ZssJi/Yz0md0zbFN7AB3FOefLqxJIaljnbAxcQK9Tsv5jv9ok9SsM8k6
S7U8W35ZpfjC/9v6La7qvSQb2JuSpUrjYtb1G+QjueV+B5sszLnx8IKlR8QKaPIV
vgH+loTAp4CjdVR6X7s0XDu0TlOGLKkkRNJK1Jm7+16jxF9O1Uhsvi80JXDvGH3f
qhW0UGIfEwa+dzWb+pWYJ1xFL49kaqMT1uXoc90pqOGEfOrt1ydgbE0em0WANEja
VLIDLHYKe5Cetn9Bly8+n/NQNVJD89TNC6ivtne2KjhyCBbfMxjYcBeS8L/lwLLw
erbw9Fe6H8evISwy36DH94kF06W02b2Y7Rh55HIGgZXZgAUM8zSSMRkKRGHUl4j2
Qfr9XNLOM/BHCtjL9W6eRWrjDPBrNDkos9FPPmjq/kG9YHexGud8fJyi8ZG8DCxi
vlXp9rJj/oC3zeur5J0aQOnMnUoYKaZ2yKaLbsAvYJtngk7EVesLCfK4x9yISvtm
Q/66SkYq6ek7vAW4s9tCF5YRy//iEh43bwvIS8eWpSsx9ZBVeck5emCTefnOJOMg
ryHe/QURXqO/k8nkSXap5AkXjRqTj/gdIqcgi1y8HluWzCz7SRLGP5uyzNhW56mC
MBtdYNVp809CttFz+MNctGhzR4rTSL1dr/5lWcQ/7ALXd3DEUvB3aRF7RQO4UUCa
gs24Njis/KaPdCGuU9OGHdMMATRJihHWjyPNJ+AEkRibidofbH4rqNW7vQUSV7f0
77pdLCbTUBApiHqK/8jQHhn+u3ufdz+JbcmqGzN7iDvGQCJw3TGq/MXFVc3nqE9g
fJtL0c7tqsXuO8h3IBb27GjKixDzFDp3/PgwC6kNrlfgnm1yBZju/r8Vn+Q5LmMg
AlfYCTsdnRCHbMDt6CRAXO5fkuq25s2i3iYgG0yL9XtKjp/jwa+e9aQPN7huJXQ0
VPatC7ud95lGj6AyJgWYIIjYpoS9T2s4W3caFgvt+ky4rDWFN7SAjy5+LZADoC6U
3QCCLFCMlFCYIvlvAUcBbg/87Yw4KodfthYxlcOOQHS1ZrFeOV4U2ZFOoinvjji1
hPnaCnm9j4a30NjtM/19xglrnRiaW2+Q6AL8oc6pKWGopHJLmUbbrj4lAW2H+uug
CqkWrjz61EZtfVqsuFgN66DlCItaAgvhqmjijedo1FY1COUwLLhn6D3xl0u9S+QB
7+j0ryK/2IcSFo53cEqZWvgk+YLmK/NgM2UoH89meAAfaaIrHkm7ejxmLaFIJJHH
7XJNQJ0noR2CvKtNGwdX0m8UWkd0giY5MV/4gGqotzkSkRZLpn4fA4IEGAKXrqd8
l7eCK84pOF82wogTf/fuN4+bzai1qz5U1SV+YAn1CsoQKS3gb4sTwAUfWDbxWo6N
+X1P9zoDje5S2Jt6AHgiCQNQb2fGvC9AR1hMl3uKHMFBroGYQT8C3W1uFlGG11LF
7qdgyZAZFcXTobC1E9BHgKrg8G3MadBf1ne9umqUq5BEsKIlHkbq/Hfu/BxpWXnn
EqYlVFnquAizYrYaWWqw5jqKO/CCNbV1//neV9w+U+MyfM3jq332AEoKRV6zOypV
aCTuf98CD01F/wHm9fk1ACukYHStShZAletahivtw40NhFSpiaKdjktFHUsqyniq
t+M15emVf9h+yzV5WivhpSLp3KnQUqKXw1TkAqZBhhA2NFjiDlrgiBusrmUNUyXp
xBFzaSyVsEGAkcKiNde2sXI9lI95Reby+CojKDAvDby/rwA3VzEj/xTUgegHCKaf
7iwj1YcSC2G6gSB22OausNShbV+uXyx7Zay87iaLSVPPEEtvPUSmEIB6eS6px5Mw
NE9ZvIM5NXLxOk3ndiUlp1JpmDUM0nVfR466tP8dKdLTJebucjmDSA9dKrBFhcHQ
f9fJN8WODjscqWUkdhjQbTlTV5BwL9b/oToGEwyjj2b2EKRwDeZ0oA9RZgVzRKkG
8Bs3047RFu0pDSQIpDCFwTFUhpguTk2L/72JY5AjHA/NSaoVz4U2AAEbgMz90iLQ
wPsGC+J98BzUD8SyFxll0VhmJHZJd1IooFHmortbJoG3CHUGbkWKSDf2bqRfKkGr
wFJA6r9gZYpXnPDTvsnVM1Lp/PkQF5aNjpD5HYb10JGPfJcgcSL2BSSaZaHpBwZL
JUK0fYC69FyjDT1arGso+2UedN6nOhC01sGZoYEhcvjAvU21p5m3ykcfGVg6hjll
QybB5cOZr0s3eLG0Zoo/vK9QHMzMyBYdpHVIIGkT200cbHwJtY8qqsI4Xtyp0Cgp
wJ+A0ByWt+Tz/p6zKo6c769s8OXW4aDyQoLUDm0ZXME38gWuwS5rRMOLrnEH8CiW
JYhEl9k7B0F9Ks8B3n+iJ9TEyNzsT7m9mhgX/sekC5e+EzH7pD6ifrXS72N4jBch
R84TeoOcmXVNKHdW5EFTHwrOiF0LhKOMN6jLLv7xVGtZKqQ6wU874oXCigji+ruj
n5NN6gSHgI2TGpNaSbeE9bcTE6xRqtD+qbWdo6yGedRrruNrqoIYpRevzvpp/b4L
0LaFkeg40/EkAItx0E/TPZjEH/fedJSjRew8ZbDFORjK4i20tasWsWudlVNtPnPe
2X3r4GBfSO7rxNrhppNJ7Fs1UB0Q6zRr266X13scXJJbRx1nRIrKGYMB//8Di1u0
tuahcjqPhKaspBOAZJJCYzQ7sRzXlLZb0qdNgzLgrIc4qJD1JvOlGW5kjlIw765T
6qR6mkKaPKs01/4jyzyOy76/zExLqQezka7XvwJYh1xaeXkGoChbIV1IB5fYTc4K
8/GpeO+XcXFY6Id/bXUDa37yu4sWJ1uCCXuzVNeAC7fSvJd2K8Isi63tsm0cKN0K
jcPp+rRd/1nD+zNZnXwnUET0EioxsZgBZyKs02b7m9z6hc1RqgGIGCGUDxeYcJ79
RaO5i2XeHBH1mC75O+0wREkpwL7HzjhZL93hhYJHVCDSVQFc1eo2CXkHfe4/kPO+
tvMNLYFNLkRbA/ox9Hc2w2pAXRPM+hcfvEnfGpSEeOHU5/Jo60kQHZHNcB0QB+jp
WmmtdcXtTnhlyqcFC7U+qa2iuDL+VD7TL3mKl2iIvaK6IG3QE6ehkLLU+Amic5aJ
6BO3eRUVeiFfJ105ojV+uPxX+F7xLlpiqnfMnth20KuCFzZqp7PEZN5K8EjvpinO
23hvESF2sSm73ZCKGvdE7qtjpSqRorPWZcZTs77kVpE7bsRq+r1X34dd4f3j3lgz
v/98tlzpd1DSqECyxcOJA02LIWe14RtgfzAivf876j1fHvWEw+tLPh69hPY6d2+y
PvYzyodl9Ov/Wsqr0+p5cK4tEQAomaOiCpobO6AXEO+oxccJa/jucYvoQh6kC3uV
KZ/qJ0cglIlbsWQEkaHflXdghLvnS+cmx7hHPRhfJePFopOUih0NmVO9DqqLkb66
K7Ryt8fMrKiMWMyBvGl3pnlSzCvbqIai9e+hcyc9JF0sOlFZWXhOw4NpETspgE/d
O4CzV7OSAhauON5FGRu2EUkgSM2l4gX/YafxDJhMYA0hpgQ7rkovUv9qCPW+MCHJ
eJkXt1GiWi6lO65PTDQWCK5tmlCkyb+owvskkTJFKXTqlYcIcIJCsw9jb7Oddoae
Bg9iLTestykKeQ+HurWs+07wxb8xMAXPp5yjtn8Sc84EfOMeQw+VyuW+aS2hE1j2
H5csZNuo/tk1o7f87hSs6ePLvAbrQCMMzD0A/K9e5ijxcEwLT3rkP/hEa+IjbI1m
U0iRxU1pJ2WUUkwcDM9VrTO2QoE/hLxKRP8ZSQPITAtg0rbV8a0vVyz93Oq1BKO7
ADGFZZKxsySWa4HYarSl/+75V4kWQClIIwvA3C3Vht312m6gZOqDZbdo5pyKcj38
Z5oNaGd8jWJaflNRkiTPIsShgnEUvOW0K+R5N7kDISEBj7C382g4p80Ab9Sw5INn
DoG4WmSiZB+RoJH8d3lYyp6jVVeVdmCyhzEJEFxyD2YaKH+YpaY9zYJ72kP4gqx3
M/xHt8S7piBnY5VlRYzLC8z/c7APxgPDPfKB9Vr8mjkGGM3svLOYfABBNVliQ4JV
KvLu6DGbLXA/WUPYinTwhtScsy8s4OK9xqJtW8ED8QQEqXrienB4ibVaqvqFYFOi
3qykwY4LrXRGs74g3A3VO925sGfIYTDgNhKps6Kf9j8rcra/bVBa/SDRJiNGtg1u
/AMaefGGDQxvFjDhjytFcgT/+TD8oUgzyxcxsRM7InEX32+oB3Uwcs48IxsGdEoo
T5h9E0fQ23GPPNq0gJ51mvRrxxt6FS5nWW6X0vziKYjDSsd3zrzk1wzi4wjXnnUi
kKY3D6J4ZsBj4SpKs9QhOpGgBi9JYX7Z6CZ/5FvHs3epCD7wRWW97Gac4AZtpv3r
WIExYa0i50F4xxEXDEA8Qp5yFNrTj90rHRyUknPU9vDkM4UIyrNiWMWbozVv6SUi
PlYK7mYeXFBVNMHg/OrMdborLS4XZD05L0zuilkKQ6ZeTG27vrxQQDs66RQVikoc
6St1iltmGP3TeMZA0MfCOG4OixAhWxFi7D06xJcoDE23fpcoplwIrSOKeGKZhv7t
WVZXazXXFA2MfymD/QGDc4VDUOIqtapIxLYbcDLBWchisMFe/eEPOteT2CaRXQHI
xYKDKJA7X0C2ePV77NdnjiKOuxVZH2ZkPww7saES4ABOW6RN05fLcKled5H9dEX3
OmawGCggi52mIaUYk5fm9lTFHWPgyRiPGyuh71TWKhjdQWL4cPcggtCzyONlNkCx
/+wTKsVuzAom5RrEvBOprKjZZdJA5Ge2VO9g+BHHzt6LvLduNMQeOxaYZkLKxk7I
4kdVvpOf2J1irmZIRXi7zvGi3uYrdUeU3beHeJhtnKgVmL7LdrET9oOyMpjHsot9
37DkweL1Eb4G3zanI7Awkw9vMQV1ofVnSbvzCS1Hnr7IYOXfXpUJD+rYuFFUeVFI
8L6t8aq8wCR5Xc9njy+PaOeGgLAGhnUlOgWOnyFhKBSSFSOVOrRCWFg0iG84yCAD
E+ZwlvRetc1ZMLawTIWPnwzlgWxQsjmaKQhlX8DiRfAGhOM0IwLOthW2Ls10ne4U
AG7BbfksXFFpYmBlOaevgw7cwEMJKbbk4QafZPOh3mYo3aRi+wfhJwtBNQuy8oA5
jdUopFfyRBxHLeSpfgZHQv1gE9hYl5TR1sZbCKFVBqP9hOfO1BFXFpwf6BqrS9xE
GGLuJYFnXM3M6voy+IAy8zrJ6b6yRyQ9h/5yVlElvHKHKBy+bgaxdFErVvMi0wk/
rIDgwxP2n8DQzsFyrydjgXds1OG0bZwV/VOGbFIETUPZF2RV2O7Yjxh+Z3GLl0HG
vBZ43rm5h+SaIvqDrSzH+rMPzfqtxK9AIFvlYQdmjA0wfvHoYZ1W9pi2mI/c73tX
x3zh/pYNDssZGXs05o/n0yBY1sCKDbjvIN4eXtY3NXX3DyM9ne3mfO/8wW2xyHh3
+Hb/sQ39VG54UKO4ogO6nLTejZFwG8UUlTu9nsbTQj3+JaqDpYvOqMC130++tmAN
svuliHuRG3MVDUX3erLkOAOQduI/ZmskbdWeAf/A5R0fK71I32E1WwDsQPsI7Yba
an7mvigU0WgFCPyMYo+BDDtT1ac8a3ClL9naYxWEnRSw85QIXu6t37/Gee338F/2
xDGACApKQFSiqcZRNqXRUpBYdodK2FeNYRepp0NcS0b5jOUZqbxZG1mU3IF4n88K
IahoAiWbYNsJXpSdgo71AWxWjvOQAvVsWoZzl6xq3rxlo5BDylS9jbOOrR5FrzIq
NkLREkEnT6vvF5fIqV9PX7XRWT58J80jGH46ssLm3yglb2J0qHPhHbjklKUfewMx
SoMYORyxR5MH3/pTuHxyBC6now3cws2nD0uAN+N28wriWO6Gm6cgP9RJE2LO3u4b
9hTzzFD2nXgW73Qzsg3PkzE2A/7eH/RpYaF7MSk6ikfZt+q320btdndATdEh0Ebf
FeCGGozT6PWaPyfvgj5YRLcNeF4DLwbULyKmVU/un367FcX3ytXy/nliRs75ptr7
+9K/5WT3a4BVOZWzeTdQhmXfecJeCTvuzdj6FZNQaZkFXfAXaaozT/YmVqmx2nCt
kT5ucLdPpdiZHBs4ekNluvcCipu6alaF2uGDcH3PY8+w8KGhwTxK21pwjv3NqHbQ
1oAH+B4ao6jdzzHMhS/YzsJHgbg9AIql2/iBiQhFSdLiZiTPkW/VHWVmmcwF69on
T3ZnMZDHDhkHVs9T/QTSX9FCTCooqYrAPY44LhLRByOBnZmZabcfLA9O0nqCUUez
o+ctNhrU8MB5l9qt2aeAq01IeBOv0+bSl26e8wLMQnlEXaYmJ2BpgeGte7XBMT6g
ygsZUpAOHvd45tumWy56gEfGTmOvg7eAcAiyFNitpQgd8EPY2NMudWGstTz7ZAzD
UScKzXJvbrJOQplgWoL1oLfaSdqaAqyhrJX/pmzvlq25DXhdr4/AsaVvUiCvCgiU
HNtLinNM/95BqogfvjjbgtKphXhLToUXRK2/s0D232VvMX528XisdxLdKAEWN+rZ
IUkhJX3+bEOzy2PHPsp6hwlcfd6fgLNYIodZ4CQc+t91vGE/g7SZUbapgOvK6yYH
rhg7LBevPQvbcChR0te2gjSdwprxiADZdkZYW36+cU6iZOlWyMU1P9mt8i0R3cD5
JU7DEF4EmV2Pu59USBto0FjA2Z1PCvMElXy4EkIA8DR5+hrGuiAo5YmDakkwrF1w
rtgdCTx9DvNeLoOMj+DnH1zfL3KSoyO5wXipgyn8AMdrKgetHbrsYBTmCoKPUuUl
Vz6sSkRoW8BFBUCXxtTeN1mqTw7iEwvIACLZGaggNvvzlJz/u2vjzYOQx/ZAVnr9
0W5wxOv84VPa1J9GLBMYDnliPLLn7lXwGuN3yPXNSQibyPlbbdwlEzmmUUnhMyVc
XChFO53fin8QOnzQKZKsk3NgNRYx+1Ydm8+385DI8IsKVS0ohklU8NkI8CCMpm6H
P6fKakbNaK4Yle8w0CiGsokhVb/CgjHPBsahXjdi83TVj7zez6tKAhOwUfz2rD/+
Vr3tsA9G4b7nKUpByJjnBrl3jZ1bCV6u5kS7WEOpLDuIFCZuhFzjkiXzABBLA6jA
gUS1K4wZW6Qnk54iL5cAHyU8y9jI2mFXPSRZD4qetkW6tE69gISjXfYG6x9rc8JW
kKI1Vgo2fLtZUdaQVwUAx2raL3b5fT1nYRmAFAChmycPQeaf87uLI+qUuyomST8c
Hu5Qmf3Wrc++gwq0wsLKiqp98Qc8047mMF9UghGnz33miiZsEBIJXCBYg4kkAEkG
cSSQ4pTNlwdJKdLZLjdNKnXScjDobLJZ6JOiHTpUH/w8WDHDm7lqEumjOF94orXk
v0kyFVm6tm3DPEuTiKVcRstsSGrqM1NUkUc3fRDNvbTf12zwVM7fL/Q5HgGyyaTU
1ogB9K6tbVi3OVCmAAJvOwhRKFDB9rymZ+pD0eciQGc24WSlewO9nIXB+hQnAbZT
xOaGAal1TepkfHA4QteSYt24BVI2KJwDt9x/5oNBX0H2Xdw4XABiG5ojGnOnm9Mo
nzQtyp+5x5XyBP8mwgn7+S7lykSQwSWUIw4puXCjSorp55wTvnqk7i1YukQyVrf+
8rOyZfK7/EoRbKdHdpQU1bDJEOUhhYlkiXtNm14RjThcZdLLZ01V/ZURT/ggNgGB
Ngk3uz6Vm0y3+wNDu/quNX1+mg27GEGwyg+g0EzQx6tp5qjVRxULPsX+uPsZywnA
SoHLuhvWa7+jzclNGDQUwnG2olMTZe6Moa5q+PrV65IfhFgpwvGpvH7MKWmptBDx
bOeEKlYg1Q1vvIUGcHYQrcUKxwbFMldGHkjur9Q5VHhjJzsPvZFlQi166Ka3q+wL
kIV84bFMjokyND7IBxSuYFYM0yUocfStC+54iCmgSEUyUuqPavPrey9WmBpSCYQV
8hofR4SuUuZMrew7zRi/pQOZ37fr0RXGZFJbhSGfsMnHuMcbXlxz7Qw43TxmGs/f
0ZEZvf8OTZFsDjURdp94lySqLt0Q5BKh1mniWjfoCd8DcBk8xYNzX+lSoRE61/21
5OLmyZdPU9DMsR1d1Qx4KIwy1yy4ydGA3AlZaRP4urAGSTvYZXD0abP9qWU1zqSN
1xHldmc97/feFz9+IpsVTH3OYmN2zzMKoNLcNNnKE2L3lc3x9uE1F1XBQ3FfE4CS
A+4OB2yNTiufYQZ9NGwUUlXPKeCKlD+uLR48fP9QEy5o558hPVnoOGwDV/7MRJzh
qghUDiEfMhX81PslQR8zHh5AC49pyKoJYymrI/eXNnLJAyKpq5a9gGjSfKG2+s6M
lo5VYqcJZNQZVN1mWV88dQEc+VBnFCvxns4sRMR8ItfW210RNhIoiHOsGNa75YFO
q95CRu4xQCTlnJ1N+X8tXueAouNalYDozE93DK6yaVYHqejJDOF61NuLZfdCj04T
7HJx1gQnW2JJlqAVXxaKtHzcxJE0yvlXbPsHhcwBIPp6AmHPwlTf1D1A7bnt6wfA
zCe1CAQvUlFKns2vs6W1CRAdLQZFtswWaJq4b2pi3TRa1IxHF2Amki131O6XEDEz
VHHAnXqhdWPW6t8lHKlAVOHoC5pxNmr+Gd78DlW4tW02FHqToa0ki7h1pg+jauE4
1xRDl2PCvy8Efu9B7SD/JaRowwL0QA7Wc2nJs7A2S8Cv3twSUCg6dtXxNMmxJFkV
Mx1DUbhDRERQQ7iJhbNwDgKW9JF56yi/au+5b2AL0j7YOe4eJAqSF4gPIdDSulqe
W2NuGpCRLjvh3o9ckQLesRPrK39I3OCchzEAs7wWyZyL4dr1UnP+Szz+wb+u/fmd
xvFWw5dKnKb84x0puBQv2Lx2tXcDZIqQJ1uqBfpQjskaw/AnnAvNS9BXPHV5W4OJ
ph7pfIEcZH+S8OmpjHwr+7igPGRMfN8dvnQeICjFO4gTtDn4rMgoLc12/Mcj7QA5
f315h1kVssEAeEuxB5O1rnpkCKtK752Taoc4kagRUSSDEg1Dixtzpori2IqHGC2X
AwvHQgqcjEVbjcvoeOpiGhtn+61f5cedvKwi1QWImqL5RB55H8pQi73XGp4LZo1T
zUPsDfvT4nbpr1zdggXuSRYGqXakB0SVe7YnZH0/kS6yKJKQFegfLNzLRBtZEqAG
BgiVqOJ5f0VAEHQrc/8LZPueVZDfrE8XUjrJE0gIQjbAo1bMDzrNEAnzXmKdYgcX
e2BfJAKr8OuRVWz9HqJsBgUGKIAmh0UPO64DWRcZTBu7raeZB56B4Pd9IJstsof1
P3P3W7IPfWvEqURelepwg4DJNqqooxxWQYs6WbhcEZewAxSZ48Rq/cGpznVY5lsv
rO5jjWTVrqubZxnG0ptb+PqOFe332NeqvgEOw6mh2kutO/lnqXbFKWVb3ZK8nspj
sWdKYvIMxnE/9TIt2xxvG8X8+c2WmxhMFRf4IglKb7BXzhvGW2gHmfAQNtJ7q0AQ
dVh2ucDvONXYIeolwICpSxIV5JhaUauNZzWRjVrDbXysXz/UBD3GAJFfSqUcjQ2k
Ec5zJ6QCi6ETR+HIw9Uee2HM++KGBjD9dxYV+yIEBHzhAjyCmwaXa403ovar5IJO
OkeCU1x3r3uQGHzQ2a5E4NsM8mf3o+gax562MM57YJQI7aCm/brT3L/USSHsPxm/
otRkrH53uQ5NQqMx60uCBxCf4IDxOvkFMnNIYazCJQPHMuwhsZH3pMKuEtZD0Cci
Zm71hjvKYT3+6JHgNidwnKpnFlqwugkvMwCgHSqJ2cSGn0+Qlu1OuB7mJrCx+6w4
ut+1R9p21Tfn572YRelcLWoBuM9J8UHaNcKiS1MZMNgzFqcs6+f+6IqjtqP/qQau
qn4hKxK/yuq61KeOLHNxmMX1cTMpySu6qZN7Oe4YAaZyqxtuLQgFGeBVdTMydE0O
dQI1f8GF4WFqKRWUp7lQXGoAjRU8xrxyL4Jf2zec7mtyusfqzmUP7vLuawPPP19d
scZBfb/DMeJ5aR0UTYBwjH1bx8S59Fah5LuoIO8ZD0RucsYdGo9VKl8ebJUhaSiu
jcyy42XuKR1XG5U+VHVzqHkEPRMh7lVCRujpzP9OPpQhySMiYCDUkIPDZdQHkPD0
EaSUzqqxqvNc66n0S4xICXXxBuq5bvcmlfewoJO5vqDICaXspZpnZHrQjUr1yYZe
rYTX6j6pq9+j3YZcwJzHx1TOErqaG3tNozVhllUSZ3fWx//YDBxCG7DZjgyCUjxb
A4vEW801BHqy/u2DAj3RzCC4H0w/i7qpvg6KkjdHPqEzz87jEldOIEwteGqOwmv9
om0dTbHQ0pOSezXB+g4qs7Xhd3y0tLFGM2It3gyt8gUIKYLVBXq3ayMSZvQHlTW1
rt2qhJC6EhMlmvKwJi6VnOXKW+fY3f8RcDKKDKbP6H1rNB1seXbP9iLYNFRgQQot
1xrC4kkKdkkg31tw2/oBPR5S4ae+R0T7MLX3xc+NYCoSZ6VyYRutjgw2ss5JTG7f
+90T1urDfIH/cG4VY9Lj6v4Hl0kO5fbpYsGlGtdjVVukyvzpJoWBgFU8t/viQPqO
acFPBxBF8PMax7gDHFAvFs/VR/5xhBP337C8bLvQRO03VIyzooJvB4CS+VevsB6t
hgtGyjoLc1DsBZMaiD/MDRlDSSAaT9ZOakRBGMhESWNEeK46QuXFbBTvbvzucooW
pPzyqxLnwQtggAkFo7M12/MnzriSCqqC2kgptgnlg7PiNbda3LvLi1zhxuafjfZR
zGSm7GkU2EyvgKCmO5x8+jL2b/KtQSg5p1qaLZzwy8mc4FeAa9Yrw32+n0KNjDQz
XbQHsXwzZoHHj6cj6GoDXRV9CTAHusIRXSbQQg/5IqyBaZMg8pXOEtWvU9KfImjR
2mIdp3jp/T6T7VH7yBEvK8KCZ7ZmiyfJgzMpUtAeJ5NwW4CITXdRTYLLmSQOw+A1
9rpFMUJct6teTZbCwmIYyA7WmlWY1ZLLb2pu7CKSkFTEaA/BCS0OGNrfE1N4vMfn
pFbyg/U9y5BG5464KCtEShNRNHofsHwc+h/Tq0a/IRV0wFucI6OD7D2YMWBKHC2/
mLX/SL9qHnh61oovL5iraoWgA4nRm8NSZkLwOdlZwbVgDLqJP7Duep06DEnl2M1S
/vV7Dtch0QudnutCSMU4labQETbVx6LJZPbwCwAlgK+a+DT2cR8fk8I2HSSYiAkN
d0sBYPId9M3FTbfK+YgOf4qDuFh4D1pYeTLkp/MsCa+DkAyqAzyE5J8iipp0JW/v
7bcfV1vNsmp8o7V/Y2rTEqvqKafGlwjFWficfI5dbozCPAyZGo1w6acwwnuQ4QNR
Is++MPTmJl1867/uvQ7szO0moNOuO5KGGToxIb7y7o5hpGVW1xK9P2Km+HOGHPWO
mtsWqdHcUZvwYmKhhEHB9ivAJdv0CTjG47ZSnXihlT3E7bftfsEwJRlIe7r/b3tt
SNBe9dBGVo+uXjgaBCZMSPsgabJ70hRFuTDQKVFawn7HALnuBoJCw+eJbQGK3Q47
aN9n2zvcwagdOjnTEGIiDt+rfTWELLMSTZvyMuiP1XWLgU+46a+R+hj0hzQ9kkKE
PF5Hz80K65F0yHqa6Ja79msVRnqjdZNKKz4yF7SWEMPe9bzOTSjmE1WpnyIN79GR
okixjJJbPz33hJ687aOSY4v9Dmys+2Gnfaq3zxomp8O4LsEbkklwM/LokaOIat08
xAnIucIrS5Seb2Zbw3hQKGmPyIBnQjwS9w39TvkDBkggpKahJnlsuvitijfZGnpR
do4hnw6XY5DCJTsCPgpsKjJWp8MqiPH6FRGYc1pnibO12c250GKPlxD+ESiYecgu
XuO65HcsBlTgAC2mUBnWXqXsjHS/DA+of/532pE2qyjKrI5OxHLX3+q0ObaeBj8N
l+PCLWRxNC+dNwIyir6gKXsDBCJZEK+xhSug3WE2P/Emad5sZV3SdMYu/kYl6PVi
0OOwoR01YJeH287FVtBXCZ7HqLrFHVxLeTjkXdGCt+mmQ2N2NYZVm0v0m0ebj1C7
PSBE1iUSDn3rUjsOAQvg5iu9+YAB6Uwi//8D6HamuVeKsAY+Mz0Iilp87EJra3Tl
JjvzFUrWduNDMOx3o2AdwANUOTzCLS+Q9vFZEUBHsZPxyNR2lMXpuAIv0Ys6SFUD
qZzx4IcMwMhoCET54Spjv82kQbSIX5tOBVSnjtBm/p1QoMSLgXY6xgV/+b9TCRJN
gDNftQGHjZbb8mz9gjRoNtnFUxYH3FHuUPSkT+FeCroyCjMcM2ZQp63f9mgIV5aL
gPMCKUWWzNVS1YO1u9VBnrc/GD114D25KurXFEMLTqHM5DYTSmeFbacFe8sa+RaC
VeIgSfeoCaDtkZUz+C7FTLhUXG5THomcZFW2mifOfCee4qumTagzJMpQFvhv/rkd
WBXjl2jWREKaHkTXf72rKlyq23p2uS41PN5eo6KoaruomNtTr6uSJ5P75QSWL2Fy
rjPxjiGrL402gPPWo9DAzSzgUKv74tUlGeYkQP0Jwd1A23dY9JE+DnA5JteFOGTA
wbKUAnx77PqIC55NUxYmZgXxtb+pUreYxqiydaf5Ax051qeFmWGzgDAO/YMPIMNL
xWh9VfhwU7HbF0Xk35yh6eDlZUDEh421KPjUgsGMztys6zAdPHatXOA/npDDf3X2
RTHF6KSHJTYZJUMd1dn0zDA4HOrvE6Yvf+sVwv+OHDXPCV1puQO6EWwKnZ8Hva+i
SDCltF+5mfpxE6VoQl57ZPl9ukklMuZD8hoW4OJ7GYKR+EwUFOMSovbDgJ7gg940
80uFenhLQNH8NL5zGzLuwFyIUdqB655QiyVoMfQFzvtHLa38e4A5JsNGjyH7Hpx3
J5YtcaA0+MgJBjLghxYwXDVB9KMiU9/ADcE+HlVSolc0wZSdmAMb4T0ne4a2lIzY
+wYFJbKUDJ18X7T4KFyjHuJBv5wkyogXFa24Bx5d+StpKES9MYQ3gl1v+U6vYcts
UesFFBlRetpRU6kCCplNAF4Fgn/vry2eJn8dtMADFZL7HDpMIjcNtrlV3bsOhVN0
SwnsXXKaOqsmac1d02TphkYk9oJoxoTqwNXOQSvw1PjGVeOPtUvyhjDKk0kNdBMC
mYa9vMPzaV3Mx+J3G7c6fK44A4zocrIyz+G58853IeaW+8Z2lG728YLQ8hIdnqB+
qwPh3Ppb2LVMGkqoIE+U96odcUVJPWwgGHcZWnne9LwiyBFx15xRw9UnBzVIEmQp
TIWlBQgm03AbeXZgDGpaST6gTNyz89IRatRVfo+XFLTIL4gsuL41Ypb+1QTBOg0q
XhjovWGLlrGjZoz5v1uDLjHXOdf3gpcVJtuzlb4OUiyP0gfjU3Hwp/4io/f7PZ7M
BKZle/gtiBWLRCPz4tCbwE7B3MakMoVxxnD9fbT6TaSj//M0kScn60jfDnXE0ujc
Avqe5SNGlVKW/lYgdoNyC3hSskouzgr6phprLmKSSiqzxsWfsBDjFLBMaGSx4e5g
/WJCPyyXGVuo1LOEg8W5hUqviqFsVTdE4EdVLJw/gZ1bgMqG8SqRui0X0GKrHTwd
to2Qi3pMjyZ+LT0615WfXJsSpgp3D2Bu/tKXqCdtGH/TNdZ9IWTaZQX6qtrj6El/
D8IaBUO1kH6s5UEwqCLZAutA1PLSW2QOYL91yC3pUVluJ02HFiYfspo1rdgIdHEP
yJzYeWzGKOXQ/eh4IVu8WmBhQhCWJpAqVrJ5v6GxFMrqjCAKJK7B+5whMwK+pqMg
e2cqQypVhT9W47zdKqluVMaXUx3j/NK2QaT+4B7DhvwJdWP4h0d81tU7akSCpvxg
1M8Hvbdwg4vePWCvu0oEUysomWK1NMaaxelrGUrDu56oddVs7HLvugGAIWQyUaPS
y0N+QF079blnHxjGOCVuW6VPX7M2mf49po2PrPz5lhFUvMe6FmtI0I9oTb8ZEgjX
TtGxqErqoLXlWCj5KqKSrMdv/8sUktK9QiUFOQI/kf4C+fDMpU2W+EByqFlSPB4J
OL3R53UN1LxMG6vpQJaZAqZtvO+TKFwkfU8BsVhrPqq2ku9N4E1Fe8SHZNyk9djC
67ipq+6HbL/Vsi+qz+weebwSggn7/YggQ3HQbeNlrYyuDEy1gz/ix+2GtC5f4XnS
loQZ+e+o/cnRd+BLICzFg9OKpfhuZuPqmuzGf+bMqqn75RIxgZtPZLx9Ct8kLMT6
S2iL3q4Pr7f2up5HUqg2qGXygh4SeOyg4/v7C2+Meo+YZG9kXcYbgSEku8jbUh3D
Xn0lHHIFTC4ueBZjR05MgRlSVpP15R2hfp+DzrhoF6rFmILLZLYnNzqUHrevqhF4
O0aSSOH06ds/OxVXE56WEddQ0+0U8DiA41zK8jGSXDYGD6D2hGhmaWYKTT2YJkcJ
UP35AAP61nnFMhZYpoHpcbBqLfOB07hw1E0+kX88It0Bgv4zY3tbQycQpQjbj+8i
7LQ36VdbAFAWjqDb+ZIUJzF0T5GyVEok5GH7nU8M4vdveQ0vd/jyJTg48LKriPKv
3a5cWi2jrNhCje1ZYg8iOxMdt/S06xfc4lYmdN/DCvO97MpfC+wflF+MLNKF5KsD
JicqwY63mlP2WrFTDRr72p8rhwbdw43WZEOiUTfQ8mzc/LNTRJM7SHgRw9s7JpVz
Gs3BX9YqSTi1X5FdAf1WSRCv01JpY/TWMe+ausCqBWNPLDayBkHpZ9BSm/IuG/b9
zWBJT/WSG/raGnv8M1lk5Qx5dQREdqiYMPywSt+4YXTtQGleS+hjXEhaxeFTlHpr
V7ZnQfLRCYCFnnkWj3l2MdDGMuaSr1ExKHA2H670okYlLVJnTAz+RfzmbI+avj5o
JV+z7JLGRE07h3RQK0T27CEZmGxXxkNzP/7RNd0/k2fAD5z0Cc6mTKytWroxzLdw
Ar1jCTXtMgp8xypUsGGpY/S9sSTmrtwCX8uU3TP86Rza/nVKiSviCw4uK2cfXtMH
2fQFLHx46Yn/z5ZBBeWHDXFfbLIr5IkgGOWhpKJzARqnf83IpvGFCDBEb+sWp4co
fxYCZ481q9uA/Cf8Y4i+fGIU0oPf2/E8xKiP5JjYp/jJExmtjicOg8LTfSRijfAh
2XLsmsxXleB2WijQachjRbULfT3rfs0lx9N1ftXFb++rKo/WBVfSXAYbfz8cKJWk
X/OBhK2StI13dCuYHzLNQ912purRmZ+2SxigDZN6n92YqwDZ7pGt5xm0vlmcWFRk
R2xCPiaN1NsfUwtQEdwGSDSk+U2Szc1Q11q/oOHKaByGkxstgqMf6JekAXRljRFi
tv/W75s3eWuz2KWyQSaar7Pu//6Ya3bHNien98/PfDtN9X+jCiNi/lQUuDMp1owQ
2APFGkuB7EnPbwwinjWGmncs2QUXW1nOSwEvGtGPJUjW+nQySrr4FeFRSuTl+KW7
H0daAM9Gy1GIc+I8WaffCOFN628rGb7UqWZdalNqTzE0apeCzqelhW94xnYLWMA4
q1F56akvZIctY8i2U+w6vE7htOsq4bLBvUT+1Tn4g114Hdfuu0tzmAvLUQyX4rOd
oHTkhX8chhb8xK/PgGHza9s98MAVjoCLVtcuDfg+q8HA2/o7fbW7q+RWqNRs04cx
QiIRhE98r6OvOqBoAtIXaS4R5eRjZ36DCQmenOE44ip5IrcP9mglpH/Od280SL6m
GKJkwSALtanySJepTrpHRM86/rvYpkTibxj8Ad9RXwCUEdpxEMeHpkr5TjBq9U11
ZT7QsviW2ynYdU2oTwkBLVW9em2p9Xipocun+zyIoEKWyV1NhrCzQd6Xpan475f8
9+UauuStW7owkVAE2KqX4IgB0wnLUQnD4rMWBB2IOkUiR1rEliV2Qvhm+4BXhjy3
YtCsxhineYLYoN6cgfhElvs2iAVPib3M4UyZ5Wm6mH5k0L3Jd5GJWtu18KnusiQe
99KDBC+xtsn5WYnBWCWCwPzGT2nD6gzuWuKdFgwQ0NobteU9y25fstKbtQ00h8B7
2/Uz+uQmfSz/cVAynfiKC11ykUdwzoa406tKBZ79xPMpN7TJEV0G/0eoJs8nsueV
pQX5ODaDagQX9O5oYfC4w4H5cj6hTnkWCjwpdRQLfoEbWq68rAaxafRVWz6qLX75
//qAI3rwXiGvyujmh6jO/tOgBWspLi5JXrDZBC9rIe1g35VlATnaa1x1ClM4PHu3
sUP0xsDOPIbLZIrOYkROFgpznvert46jS1eRcOdFHsaFXuIAiOD96lsejsjNKwEG
cTBjcYxKAyRpsShMYKuq1HU5J6woEXk9xo/ik8WlHF+voRZugdXXBJUPSQfNpMLo
Z1M2G1BQpP0t3oC1zMsyl6+RghyWMlRBdWda32dneTJCo5Kj32qBphj682gYVga4
Pr0KRXQXlzaMrYn5Qa8nP0caQESLjNbwt/2CyV4FilcY2cBEWyg05T0hqgBdqhr7
am3wyEGePnzifreMorjuC5JKwrDsrYObUKQfitnO0JhG0+bFpBfiWec+n8CSJiCF
h0KONQ9Luhu4kSj4XTBkKSuCedl2gjM/ivaoUg9i+WxFEOzbcft0yNe2oDjQvowx
WcMFTZBDQaTwA8HfXCL+H3ZhDxDoNteOqPI7JaGD4fEXuQSd3aLHbY55Yc0ZXkJn
qoR8vZ9DGnJ8k/WmcKheM6UNOUw7R7J8Q9Mj5v7Hu4CQLWhzcUqitsnVcO3ADNIA
7o1re3CnfKjsPexxpUIDyqMSk4kTz4IoM0d7ZTtc8EIos1Lvs+vJ1ik8tm9JxMT0
MZoXGuYCgdTEnhaIBTaR00QhhdOZp5VSflRNBTVXjITET6Z3o7ixj2nbE+m6T/h6
P2qhSh7RcYgXKAB82Krzh1uP6bmd9ebs26n7COUnNaMmP6cevYBLOU3BuKvDTNok
n7qJ3p6FaLA4T3iabJ0VAOrsfkSFCZiWUCZDFGEt6Soy8fBxjJ5+/pvabiTHK6sM
Oa6CIXhKSr3fDCN1cYFw1NJz1I0zu9Vzfwlf2/wir5i2QpxrWZRH8gvivtmJLu6f
bsOU9+Eoi4J7w1gif926dI4oVkYGU0LWjtMBC8+qoGKa4n+7amjnGcgzcMG7q7ey
iv1/Gec58+LYRl+CvGK2URTclwB+LD+pa6ZgJP1xuuEIIpz6n5skrvR/78kFy3zd
eQEmn9xCm8HB15rGlK/w03DsArdItpzHTKmeSb/15DiN6YnGD3orjKj9a6dqVtcE
AtJKOODEd6bVzqHZNMkHRGhgX4xGQmpXvOHEI6g/1SRRcvxegjvRPfHvksUiejp4
4mPNpDHTWEbh43V8kjOS4fOXnmrQp/jp7sdsmSahJsWp6DYculL94EQOL9dprzXD
tcXGgct/i6hXjyO8jNN+zuG5gzv1LntK63TRgKxqVbjP1QyS39iU1L5v+aP6OgsJ
HCA4ASRzMNS9GJT6U9z0waRn3GF5EJRIaIhLPf10oRWZUgm2QEEDQ7LBs05LRx1W
II354OatG8EVnFMf4BdBMUeRCoft23GrqGrNiEdQnrBdfN2OB3DMCjXAu95k+CDd
eB+uMgcUFxxSOsRlpdg2KHB7yYhhPfK0S/rPVzYisoAuU9wRtLJy3Z0kr2VgWvpZ
TEDrZpIwmyNoci9OwiT8e92Mn/kA/pxECpnjR+Zo58onkK8UfJnprvXUM87kUyBm
NYCpdrojkykaU7o5yatII8cwKTeobepShE43VczkXEoLtdH0zoxvwYNZtq+GGc1L
rT2x+xLMWDcVZXkN+aE/W9EIAY7whgwqPtKwNfL9GARVj8v33kOzlLaL/egGn98J
pWfwTVpbrfrwZlmkJEecMzLl7DCJxnnoAAiQpiX9pI/rd5XnehllOCZ3GByJpplu
owEjHrcyNoksY2daDhIBYsZBk5xBAcetKQKEbMeWtBSdW4i96Z7q1SBWo/DosLHX
2kQKV9+yXhoCXCjRAVFu7aZkXNekwS5yGMrMpXtV8wuezWtBzL1l2xf7U2L9OMFB
Vg+LylQTVSaNIaIFj9H7JCokXSrLO3grwkpTs5XZuHwduCiqoQ+iWj35uZelO46w
Yda5cglhwnBXLy3GFs/raLHdVNm8sd5Jtqg41/j7VFMdBtkRXifqNUp2pveaVK1t
wQGuFaRhlF2unw/v6PWJYSEO1UTeMH/kzgiIpmBGdJOPiQGuOA03kFTSTc7DnHmh
HcUYJXbPQBywpMunfMcvKSfj6nMrrPv0PlShDWpVOJQ5pcV4StLL9hPnrGT0Z6ON
uHvpg7CMxYu7kx0+A1dhQ0CQwEvQ5oUh4VE4rqLnpSielfuV8O7qdX8siGhJ5XMm
RRDUWaiMhSzN6k377NQO+yiKyTBoC7G6k7DLMVA+GXF5oUjHcXjNF2G6kPCAyykt
OwKJzyIXwpJBDqN+G0UJO11uRtjli5DZAi8JsxgDO0RY9P6u60pWMATK0DWhGdO5
QyYqYo0rYZgXzr6XwGCqCJlyRH/e5e4pWtc8s/3vkxaiSyxsN9ybGfc+c0rQ8Nis
hWhIbtdk4ADIc9L3AH8UuoEgtLPR3FkFcil/2nMQ2VTZivVxSmP3h6auTUwmBQhq
77PGbiHth548R/pmI1EM+s/A9gPihxIeTxwbjOomYnhq2/MpKgSLeqC6d99SjsCo
rbTKgVa74HxSDd/FTEgReZAyKW70EFrpR6v3Ei0aAGzSlsbfcpqW3TkzHgBgn1p5
z7gkeYuKimDbANfzbUtuvlo1wpcEY8IGf5i+Nab5oipH9IToyua6p6FZp9Rf9zuE
bJV5Ic4H0jmYCphj1kthzNDWcclPzqJBPJ8p5RF0DGCCOhzvtR8C+KaAAdJqkabW
o8DtiRcrlarOVAGdarzWOn90oDkoYMi2Ug7evOxBF/vnWDo3fNafYu9+WGgzkeSW
Q3AwdMLL7qE0sccKhVaZz8cvDA757ejInNNBIs9ICu3YLDbWMNTOroJczCLYM1Ea
B8xC9jOP9h/fE1jvmIGiPw3Gu7EkzZwFSCFdLhYMfnyrgdyI0ApaFu1Hx58B3pKA
2agnVTtQ4iF4mdADkYv/cbjaCmNkr6kGqMkIbZxnd3xnmjra5VSRlKLln97UxQD8
UfnFXQ1aMqx23ad2Fol8AB9+aqiso0M1hzmDqYKGQlY2hvLyBiWESZLZ5mYG7KxV
riQY3ZeKVryg51vIEepSO4CSbo4QG4S9GuWFtIHYX0gBdJ7pJdkSYRyurpGDqPFL
PXjyjXnJ3y2Cg3tyeTlveOoxfA+l7J5IQbs/HmIYMOzJIHik2gRJz734N+S9J305
9x7knHi85q1o+h5PoKePlGq15SB1v+PE12xs8vWJ4kxvAtznmAebN4UYU7dk6ebk
de2DBtRgpk+rPDEW9ptc51i9FUXES4Opvn5tsT93StQondBRk+UR4kJyu6xbiDWY
98ZXtzxP2OY3lNXRGzprVFnBg2A8ORDXXif5hFbp4ccH+gVBMUpa9DENd7zLw2OW
Zqts+jveU1SFqUNGfvr0qE9MII+T0zpgLHbdunKKOIIeP/TRzPvZSw1aM/U9EgRe
tVpCV/oDcoc/V5FCffycr2IgFDryMblKRrwri/KxEhFtboIYTxMZDPGLSarHEFeb
afn+gqAlL8R+7eD7fshe+5bpp4JPAUcusmWUJ/cJXGW2XLYsEnj4RNjM57SVSLBg
fQw88JqzsOyN/N/SfBiYWE3nLzm1xkh+H6gTssG8Ksq0TyqN/mF7koaFqa3dB6D2
C/SniMYUJ0LU6Ner7bzp2X0SjHYLr3Jueb/+ixoVykNnUOa4nueiAICv87sRud2f
CwCN+HdVtjuifAa1skQS0kFAWV8PfublcnrRXS0hp/Mf9BTFuNzPdf+nzmoVQeUN
qgz3lSzuhSxPqbINHqqGXl0/9rUOCVEPRDa/oyAiSNshzf3tr4R+q1/pU8z4qw1c
pJPAONopvriIiq99rrvEb6flfHiNTydV/JfJ+G+N5i9Mlc6PD7qj8/GnDld19Mh4
AktCuRXtuCVqWd4WR70glMb4V/npjacvfDjJYfAEP/izXQbv8K4PnbN5ifo2TrGM
vdTRCi0oZzU2gHN1qDiZ3ptiMJ0bvZb0n1+9Njh2QhXUVZD7ld6DZ8kZs7mKYv3Y
X+F/uNvnqE2Qak8BwoQuFh6MXd0jjU+jK9bGur/zPee3rQ7WQWyg864aZYK4UrHI
jS1lMovB4kWAUH/itV+KDUeEFYVGIb4SrRx4Z/0X5pmYyDg2833SutVAbyLJFPg1
ObxX77/FeZ1JC8bEBkY+ey/R2vKtw0WODgiTYqYpdmlWAox3aCnQLdzLSwPSbQMj
eiQMdKsZalrRQhpB5Vo8Hsftvzvx2hNtk6lZGsvAWflhAGxCqV7P9uC12zgwE6aj
YIT8QSEzytiaQOBW0WPER9DIZ+FJE4uY4jely2bncK7H+j+IjMLL+P9LgsJM1Cme
54bj6FLybpVpoHjmIcYeqTdOtgqhA4tWKw2DvONr490akH3npuDbQWPgMW9R6pT5
zZEkLNxaHkSZw8oAdeyZuxJOpsSnuCdk+EOVAhv4cfqOaPBKv4loc2EWGhQvCgej
uR67aPaR6BdmztLqxPJksVJCUzQlHrAo4oPnOR89AXf/BWLy4P/rXgaoIUOfkpc8
eoID+rJtcdimVr5j4ErWtct8p9ROj92rvAaCC6QYBKtTXtrxbYwMeKldFZrhz20t
40Hz6ZkWujCTqoNukCjAiK/55LVjfTP3tKq3oU1uHBMsqF5IDkRRgRwNjl6fjYZy
wFp1oVRjyCVocfI6PGI3qR7ka34Oxcsr//F+etGZcRtD3OJGDr/O2CTN8YwZUx4y
9nITJ9UD9vBHLmjy7gaQWCe+gUhTTCmE7pSCq37t01CCrFbPc809loeY4RevHfEz
0/dvEZh4zNfOEUXWOlXUT/pUjLpHhFWMFR8BGc1JRYUAL+/yTECQoKJGb/Olc7qM
6x19IwBFrNRXh9+3RFsi0G/gxwPLb5a9omSZVwvWw/aMofS5VVkZlIhP6KFStpvP
T5O4hKViHu3Bc7ysSRaKDE0J5aXiP2uKdxf/2olkfpCeEVIgKXrzHJ87vdVNrsN6
ccbUPP46bSIOqOlvGo19oA5XsITffO9C1Sjto1VWiBG1CFw6sNnHZIGZAg35saDv
XvST35RDBXFDAQa/iFmKNsB7IAPnq9CwgHd3C68HOhGBCeJa95ZdWdMnxDc1cq7t
jQ2a3hdoKjH8NyTbt9nNfmVaGnG1MU7jvKFIJl/9T80FlCZ1bRZcMH8bwSUmBCq3
BgvZ3vVuu3uvdijwFMHTPU4qDEsBXBWr7qYY00kfg74KHUlbloik2rmpLxYc9N9l
ktdaAOQkOQwEbAWpM0BvFRQbFKQvQVK6x/1Fh4mqNh6Cv3Sucfb7tluD8E14XOy7
trBm0sbH0ns/JH93qvK4/BG3o4asZ7DTEwDhGps9nB4tM8y1QeFK2ZiFWmvNig9X
HhnbmljRhNPiubgaRrwFSly9/2BS7rl6AQyYayd5RVtY3DbiyA3zsEtU9Vg10Hu9
DKTzWRCn5jm0x+KWcb5quP9q/D6dNqTQcntpazgX9qsNtK9wvnBqvX+nVhkFpRl/
CHR1pjJ8ZPt3cLVf87dVcHfX90Zgg5GrbZZjWo2IGqLn+BRhBDJaHWAGr/3lTRlf
k2Tg9NgEKiMvbklWmcSEBmnOrdfJkCEYCtjxOLdHpBLd0Kwe7P/rafCmUhTSAT6r
7p3Jx96iQllol6E0atTt1fZr/zR667YIsEcjzqXo+nR7pVF0pVCcQnrBIXZ3BCiZ
VHPiaKt8lYa6DvSNwHPvTKr7OD5flgQchTScMjB2gBRS72d1vgLBZDaQNz2kU6hO
SLC5130R6RkfEnz5OpZSqquXo0E4S92ep5903EwgkyzmY7tZwvp170kL4lefVkMR
c03oBo6IKitZPfY0EpgWripyZQjSrRb24IYppgObSGcpP5kxNhBMJLguDq6S15zS
kY5+wuny2BBr1UElWFv5Et+CO1NoLHo7fbikCfNpfv0dmCCIZGUI61HHydMj0nUi
5c7gnJFKacQrgIdHPlygvWkgAlQH3kg3kQlIJkWYbnKBYvNuIhZ65ZANVk+W9iGb
lj3uKkuKJSnY11H1bQauQf+k4Kf9G/DAOPdZW/6ciWSErJvrtlUuiM8yfNm+TXJ7
Ic5RDaFyycoPSHoBI3EwHCYsFHjCcmmoOAnOBx/IO+ssHGh24E8X7vd6mCPt98np
zHwbYMZbYXtOY6KCiea82oQ+cc3cqE9thimV1TNRRx48ar4orKlAJrpTgwiI0Fzz
S/N04Wbzd32RuYZWO+7Zxp3FXCBMvJLU3HCmrPLYE+LE1NMHrBHqLY+U7xvbOXvI
WEL2jbI6abdyy42zQy4cbc+gLQSmlWw0mME4Ln44Luu/nBWkUXV+TIrylW31mC31
+d8NUqBKtdtK9SgB308/O1HXUTCSEqJLTFF1W3O0g/j9UDe2q2GcTXsB0nAmX+Xr
tHr8QmlAf2hI0KKySm4Emg2BI0DJVBF+RZYes2DkT2HcGJJKMXMqt+oYrd7G1SmX
bHn8tZEp1sOP2X97O5RG0QMMPvCugL10ZecpDsxhFnLYVuAfibg7GoJWWWPe9ndZ
HYErVKOzhkdkJYZ6ZJjOuCoEJNnLni1m1biGa9/CTKDfbJLapAJ1/mrKFTfEIxfD
auxZZcr6YFNAtZhpI2g4j4yBqXNrTDea3+c4pnOkyIiL17b/YHwHHcw5e+yW5vwD
sNLzHbIF02HKOJurApX3X0coZGRx/2dtGit1MUGaOl3RltmTFCBLJNXut/UsWzRZ
QpX9IzWeddcQ6nnYAgCIWbV71ChvGJerRTzkIjhs0AXcuEFBCBGidvauQcr6lM3V
o0o9Bx8qmCRfwhLXTPhOB2RYWY66ldBxwz1c2c48syTGD/M3dxdhJXOogfQbvTJi
WaDI2t1usFzcHCya+Ke8YcRWqNCbO0PBmIUTKt18Cbdwd6+tSoGsKIlIw7a2oMpz
R0YtMozeiw7goBglU7cHdu/O3O9wHawkDfLfhUVm9Jydpk0DH79IssgNm/SN5qin
iT4gKn4x5B4VB9LuM6SuTckJ6D+Frw0o0INY0/BFIlWAvxZRmO6bFSaeDU1vJc7s
v0Agoml9y9U1jdB2Ecs0HL3bdwQ5Jmo8ntCpZKqC6pi2TxTyvI/7MrYOSM79W8Q2
g4wYG5cB6GSDam4rwGi7erhYZOMVOwr7rrPluKDvi9W6XxX7CcODvHjJCfOv+ZbH
VImUGYr2MelIWwW7QYhDsUovF5hweKAjG3TrTn5y4TysberB+MHJyw2apldBa+Mu
N4JawlsOV3gJEuX8RD7bw/9KM3gtxLxcMblKowsa0lBg8Jr/+1XLgRxuynYwHKhg
eHTluKmpv1kcyqo7/y7ujxuhOyhyckw6Ot+gDnlF5buolyMH2DzJWgsstrQ9P1Tg
p8W8zow7Px84JwwgMLlZQQiJbrGL0ZiKi1W4700XTEQtTgt7kq13AgUAsxA7PDbr
M/x9EKeCCtaBiXSoi9kNXrB9CylnTPLq1i1XM6e7AalCTRWbko1eVgAyhpECUqH8
KhZL1r8naBQ+GssroSWxuUY1zxY/ICWkX0qN+xwEOo3aNVlF0BpjeYbexQCUpjPo
X28h1GUgwIusctkqMnezYl6dDhA4lv5yYTOArTZYaXSnm2m6AkTOUXOsDpbFBvjx
Sn7pFeTSCQFBh0DqOqH9aTOomLzEdey7Vz4uPcaIA/HvTHNOdqSgxIf2lEafjI6W
AQSVhV4g5iqL2QGT/y7U+cN/G8AUbxFR67m97AKHWm1uebFlvIyTsmCR8VFXaQ+o
SgGqUKsFPMaQkNcUWMZn1sUYNvNF9m87dEYbHGL46uq9+IG5zgmf5a0L51gguPCF
VrA242XfFwkjW20jVi//4WoVy3qHGI2TEyCNZyS0qgD/wCkMRmKTNDfehCSfuGwh
YVoU7GxYvXkA2sMiycibzckex+4XmIPeKphpknm6jlT2jaTZYCm4q9BxtQVWH7si
lH7pCKoAV8Qs/iRMyoV6dUv97EQIXOVLrxHEcr2QPXC3c7tJqZKxhxFl4tMjsuC5
qq3wnYHz/0mWCgLlRq2neB/nZkwAhfbx6fwHy1/Pby6ecanQ2j8XsNIHNtN3zpUw
IGHe8a3/b3EL6SuqgllOIAbPNvb3xD2BEaJVU7Eh90qhvhruodssUmt8fx00BeBd
yrput4jousEymvnIhHM3XxaMDcu7s2+IyVH5MPprZhoogfWAFquJaek7ISUGGKW2
QIAB/fZJOENUfyJqvms+IJYyGxTyx5wM0MZBXppm+ur1wwMF9JbbFkMHVZtRMvV0
iR9cgViRhJNT7QOWDdw837qUatvzny4whokUTh63T+7ccs9zRimcliclMPw7IqMy
sl3dSOLT5Y0R9QdC2d0/KP/a9iDwr0Savs11bsE/ccRKufpMFNiRkcVlkxUgO21e
woL4tZzEbJeHzvt0IALgEsoKIIExL5ovDgsoscF5EUGh4b+tGIuZytCIJ1kYTky4
xnOx1y7KPwDsscea26dLqFg8yPt7/m0tmlC1sAQdkg12gg6lSr5dwuDLGaibhVwM
9dlYxBbBAOPVnlCiLaMC7VjUYrU0RDiVLaInDfGeGRPBzGv0bhzeRQDuui0N6dYx
OUqPlaCSkPIqVFTWir3RuLGUj3wLo8mXoLernKreOj43MIOD0163TI4aL0SyN7Yi
yPhQLpE4lzOd8vTGgleHbU1yd3lUiqdFcGJFYdbHRtZQS5QLGlYb0W8CmYuYCLB8
uI77VT3xkXg/S0VmjYUfj3hCqa01qYJ3++p6QqAOrmtKkcEBIcYfZMT73+vqe6+/
4V13aY/FemOfAYR0FQEUdhbms67RJjEAnwQfW30521l6xJbOSIE1Dp/TcdLn4a6R
5z9RpFkVyhKEfxcWnrQJ61t9C2lzR9JSFkVR0jIx0QP37MRAk++0Wi4bS9dBMeuJ
oUwN3DQnTHWcvdkDy1G8NME+tTTrE//r+0OxIdPm/UcvBvrEAzWbRNRGxXHkC54y
aOe+IPTFV1QjGJb/VdELPljpOmyCSKBKuAAefONJZu9pbsHwsNk+f+RGYRjp0vZ8
aYnp30QQpQfLK9N6mFcL9jxge+rTgnmIAxYVH+X21ctMFsIg5Me692mQj7FO3nlV
EQ8wEh2QxdLZJbh5T2X5NxQePClaN3M+Y2u3SE2Svt3INU7+HwOwgPJblLyF0yKs
uPjWwigwC8Fa3nAszM9DKzcJHLML8fzXshXEXWz5NaEE89Myy82zUqaTR3Pdqfir
sGDG0ZFRDx7yTu1mhm/x2VYhbd1y7vB0DNkD7K+q6kN64lYg5uu9NRysNpXOynlH
tU9y39HImWPvsA1xH5YkhV8RBGsrlRtzZ02u6vyHXSdIdTZ5M7FsN37+2Bbwpi1Y
VI1qshtwhbblV/TIl7AC4TIRAF0stqrmaZz9j9gVyKbD0EChcomgNxENEh5ChyIJ
SJXIhips4Zw9qP/pXodxNVc1VhoILsQ3i9ht6Vt2DxoGRQAGBNe6mYtt6nTVNZT4
mBV2SVwmyKHsGB0GFo/Bfo4rI662SUXoxRJIh2lhvYFaB1sTl3AcI00HkCiRuoDu
1TLJIAIWo5YMI7H/AhFJ3tbwS9D0zv6BagrqOdiq3Y6zlXd4WZ2Qk8WDUeW5bM16
thVH9CvqvkUX5CQYRsLrnJb5y5FbbMi/Dugo56y47PJI0ekMoGQ+LslvapSjNUPp
GRA+RN6LM68K1FpW8Adto4r1Z4S9oM6+gtuEAAFCY4Og1zUFVDWhntCmm8n2dV0Z
2AJjL3tpiNhcdj/r9SKfbvgav3x7sWXrviexCvm6DzbrISQHW4mmyNDDvT78TQn5
n2ZgjfngJ1kyMLaB+EAcoxihzd3T7mr3kL8txTquhxVSngZCCgaLHdgpp/yxNUMA
p9++A8/7H55/PgxGSgMBKn+3ZHYCKWHFIowugfHNCzO1WYhrITrEql3aYYAWFu1T
XLek03iIn3bEzEMEVNvE9Xc1tLVlupytvVnyGY8MZIi+TzgQ7W5uguHbuYh3iWiS
KTK2T800JW43iK7o2ekgpGKsSScmLIhfEdk8u7/e87wba3G/mdGmohYkZ+uK90DO
/KrnP0fWKmchVbT5Uxgmw0RFoKdBFsD8j3tD9mM7JU0cXjlYKJ4ZNqO+odnvR+yO
HBBFP2n4nHEgQmgvrI9PPMefmQBn1pOW4QQCVHF+aR7+ZbK9MGxzbjLvG1Fyw8di
pVzEw8RDYaPqLGhmEVDGDGKW+sQ8g31MZKaCtfzQnabNXiumRaavH0NCVAHyMoN6
y26aG/+n+2mqZPvo0kIlMH3wCnmshe1g32YcNoxmD/5MU8updSHQak6SthJ941kl
zHwVhtstK7AZ+OQHZBR7hy6yzxp7M7Tz1ZYzz4q0u5JCiWEOTHGwCtKAH8TbKh21
COeMPRmscGAthxDvhqcdRVNdBcCyn24gwMbs5eXd0lIrg09hjH4b7G3yLNgyGW1r
1HNrU7RaYrkgXzCbkGcNFqSCgy8kZhcMK12pzHQseUTSUlckEZrMr5moaQ0XIZNH
OmL+GVP0BJDhycRyFOu+kBWoP7G6fRkx7auGSkICFp8x52KAJsHBQ6itDUU9Ex9a
kyaARv+9Ldo3vd7L6CU51CAK56xaifvhBbWxbsPiOWvTwz/4wmD/ERyw/tTdyNGX
pSOSv75vouDThOF1mCsPZ0riXK+8X6mRcSnM9eQo7kUPVuNlZ+ODo4M9Vy3871BV
lRTkr2t7OQyntaJXMZLMXsWzAJ2pzoc5s8gPeKgM/AUj3qQNGScUzHin85rKzVio
Khde3il9zDhM3g1Q8xLWuxXMCZH596YLYVRPQIFkMLogtjnm+tysEmpfrdkqpJw0
dOpNWJyl2k0Yr+7yJmeCDuiIozU7K2qANxbCenm0upK4DG6WkK/Y87ig4r3JQYcm
vQa4YcSDND1WCA5iU5mia4Xq6r7q/iENQLgCydH5XAn2rt71TxeTyqP2hHmIoQO8
hq6Nt0dMnbtaUdScvHoZaJUWJXReqteVCsnI+71iuMCeCPHEzToCTnQrbP39vGlV
/IVwiSO/ZsJ6aTaSIPmsm19N1Cd6ndjMwE28l+0whucj/fXPCu1/qbg0pHDiqsuW
Cccl4R+cA43IhlzmN8C8GU2yK5TKJcjamwJfETiCR7tjsO2XneimxVyr63ZKzBeC
tIX9UCNVgoGyVucbTjIayLJJKjpI3k8E5UeWSSKQ3UnmCpqDjulcEBhNjN+lEGlM
JVJnM94bZ0p40/ieUzqwEAIYskK4TYTkZKiPkM2HyCMB7/GVvpxm2QRqJgaDRNwU
8xGWiTgHFo3CfCVMivHj7FmYHWAlaUmwLMnCBd+FAOWKC3nehwNbF1+RLG8tEfQ8
50yXWMf2wFE/y0YelrWzNgCJanmskWj7FPICmoIZhsGHiMk4lg/fD7+6Z4uIapNl
5FSA1/afbmw5FC1xRmegd6EKDZrRe82Ouyt+tPZIjYv0uQPpsXOWonu+FGcw9JHa
cijOWdT444TP4Zq1l7dhyG77xj2XkI+9dL46Ii8SxMZ9bNTC6sLmll3e5DMvRBSJ
x7UtJxTmEV3rQoIFVRq/yCrhpkd1O6UKDkFTL6B/LVm7P6Bii1hmW+OgzM7eJWB6
dtqNhiD0p+Tg6WRU6l3fso+4UdQ/S8aUOr5E91WiubGREbe7mFM6qttbgMDbTy5c
enlVpdAHHM8uUPovD9jvPNv4iZVRNgHIRQi+cxrBP1tedkKr/WMwHboXbLQ3G+wV
HByeHBlZupfIAOK7NU1ErotogLZhiQ7SZ400mVGX+5PPQWWhm6LiJ0MXJJjp9pXa
f4029nf0SDMsUHUjEvfq+CGB6vgLB1MS2izVS6WfIzq3gwsDssCQmdeBddXd3Dv0
2B59veyUUqvddgeI5w9Xf1J8M8VkYkBhO8x/0yfyZwA1rzouuLsQ8TbP3bwQR7XN
OHlthzzvywPOMwkgc1oD8GWM03J4j4ntlIEgQBVB4Vgs8CwPCtDowylHJ44jyWd5
osntEeYhWueSRsoSinPBVLN0ntY0h+MWRKOJk+Y239pxNpdvYusuO486TPuaCwYo
0fPPxRistUtb6Azg0ViiBtLf5hLSn2IjvB3KXulAI1n5rH0M/F7hVRMc48ZTE+10
Jjm5AJA8R/2iipFKpjTWi+lZbFImfbwTcxEd6bDq8ezx7je1Rm/iIT5HK1X1xeW9
qyIjorGgyKy7pvqBhgP3WItkD3YOAB3i/J+PwWKeDP7fPej1zRZ7XGM6J3vjuvzd
tGwS/xFaoxJHzM+bFhUwQj6XFIMgIYOYYwgU7GcjD/hMztzw+DiMAQUk91sIWbBz
8Pjo9EmVjOHYtCcsBV526P0knZdA/ae9evgS/3E3Su0T5qR0BfaoQA8/CU1qmJ71
ZSdaU3Bvk404bBd/ORAWaTCL/bIO4jrllGGZmu2I4NT8wqr9fsyHeFP7X3TRmsJk
hzPZSAfXOEI7pVL7tA2chwAB3A5Wa7D+3PKwdtZm+60vDrTtAHNacv96xH0mS3mN
xEVLjd28+jcLy3r07n8LFfDdWPcZ0zS28L0HNfUiD7EPZBaXFI1K5oe0jnpj2ZfM
R0uquAnOrbWAgxFhw1UACzhfpdOMNOsBehd27ly/YDi9bdHHJKTMMgp+1p/RbECl
ilmcCBOGgeE/wka1r7qOs/GJaXheSZM4xPKxsnXPkHxU0yQSYD3Pnv+aJHxIdxMk
JFHnUAJtlTBPEFJ9bmkA0aZvIq1ou1DHXpTE4uvipzfeuSxZqjMxr2DHoUP8fI96
taiCUsu0oUyiVYrybxk35lo1PHGeef8s04zHrgG8rxRQkp4Hzx7I01HUPJ/7ygN7
pSLj/5j/4vanX8Uxe3fF/mEcctu2ctdzZvJ72/yraAPchwE6ccxXQWaYtxTp5EXj
B9XcTVl8f7rCWT6NbqlhHAfaFFgKK454YGCE3EAKh5KQCiWV/JU8+5DvQ0KN1KMg
79l35cn+S0kfoXl2hjPBcb9kXWUone/cU3W/HwjlqgPFfGr9CRXsQnmFm3XpWf0V
mt4KRUGVgYH20E1he18EqEVZpRBzFHHUebX16hxR3gsnOsjO3Q6lRGoFdT3RQ62w
gDHskKMoKpqaPfBofs+oT2pVzO6tskRDji44oal2FsU6MRFaBo/z1VFMHZ/EWVNf
Jciq2S5BXYTEO5yLzBjFP05sgizZjGkMO/tgwyOIk8oiirM6Ez+G0YSJxmSr9iqq
4ykCsswaik3Ym7/EHhLLF0eMLwOB9/9cV2uYvi5RTthD81vUgQI9IOh//Rk3Za1r
q6RePYcKxcWVZ2Dc3F7krlVFEcY5EZuksesIsDrhkTUcjMbLy2Vgxzp9nXnz6CXD
2JqPLofBqO7ftMrkwLC5fBkN1dXYM4k2rIpJy78pYw/OuVodzYY3SizfKG7mJhx4
orKsQn1AfuHjHeks9y0pTAcZXGpravm2A7dCbqfMktqh2MW6yDZcqsGJrep3nKJv
f6Ya9AC5y7M3RTThxJ7zKeSx+pjcnCkqcdC/jsX69ELBjWnKiiY1vmPVNLe49F6V
oUhxjfYW2qOd14+L3QOsMt81sYt/wIcKfWvyK5UD4sp0UHzHh77J00d4ZXFAB5C6
IoTP2Vv4PSWYGx06WlPcgeOJ+gkCUomgPhB2NIKhB3isJ4KXT20pcfnZj3Vo/ZQu
1DVhl5tVd0N2vG7SdKa3FnzcD03gLKr2g1owxvX/a0VrpL24jHhufVEIvD9/JvOe
lXAQT8dpqIgEspds28B6ODvJ7rk8V41y7zWLlRb/RSX/kFUEQBga1nVomb8fUZx4
0Df5HajJj3a9F2S8Aj07soChqd/cLnohiIzjGe8CmhYgp4pWKWUf65bPkqS3gZCj
4RD0RSWczIDjwZZIhslRkssnaZ+P3AQPzyTurV/2S8bifTbEAXvht+A/RoUk0vOL
UEWFAw/djiw15YL+A0NIIdhvirXCIJHSRKga/Bt8gX0YiZK6FtbZnPDQpGRK/B+t
DSIF9PA2KsmFnxR2MI7Epd4nOaX4EuAQP6RTyIFwuU8dEFTfW7h3YtPKGg8a6IgK
zSEm4taZzIgJGyYRMOeuKZVNRzPxEnZ2aAZUM7+hut5YhreVHHvZ5nn6NidzH26N
jBHyhFI723qWWUkvxIj3fmNfUOmMLAW0bw6BmgGY15nzJ81MQRpXT+2rJNuv+ZBr
nU8NynbfFyufViDZMiwQbwPjr+NG0Gxo8xucCn063a7U+ax5j88B9x7zzgbjvOgh
NonxfmG0aOQ7IYVgBUtGv+oqNWD2Z/oX6OtClASVkr0BIC+E76AIpMsX5Cmhn4i9
LinYn93eBB4QaaEQOxkiywNGI2SqSEWuwpRJDrkcaQjs69gqCKWq9oKAIzJOwYzE
I+UsMBUPCkBMmLNxftGcfdeiZkTH91GrvGn4DOj+/QyFs6tfmQUGKOBSz0zy4CEO
wgeicJzScnmE1f6qq/qhScVSNgsptIsXtqdSU+KPVOi5of+4Z9twE/pgWFcK5L9d
331ZyuwjH14tZej98VO6dGsc0Fs0achUUboARk9ZW4jTH5B38+Iy/1Z39MQSL1Q8
GJiZrwepsCeXW/wNWVk+E2nbdq8J8ei7vF3eiI72O1LgtQ7Kg+bzt29MZIEXVaIT
fVOHMdiy7NyDz7M3pqjSwyoFa/ATvaZz8buYzbcqtvaNM7CCvB9c9zCuzexkXQYW
0udCH9Zc+2HraL82K9H5ihfarEr/pk8kxa+vqWpnz5LzbtLAd4mgG7dxAeZtQwi4
kc0b6ftWqadC8niruI08pNfEV1zJ0iuj73L5X1LQVWevxH42Sg+9e7d4PdICFl5h
fLzhsMFBtiSRddWXyixFHsZQgnWNLPLmu+gKF47Mg1Q3IweinrvU2CgWK6FqmZIc
csWjB57yb4S858JzSiTGNQ8Eruhrubeh8HiA9bPJ7ORjnovzbIarA3poBumebbjb
ZLTOniSOgRj1RZqOnCc4DsxtvCB9cjJky8E2w+PEB1Z4glm9vXtP2bteJZd8hlcB
EbwM0Guf6hK+QCMZCh33SgnIoP9JFHr01sCo85CfPCfRWbz5FM8kcIYXwJ+OTAQx
dJU5NSxbfaQuuYJfrvvPWy36/2J4aBN/cUmP4H5YIoXTBlVoj8fshSYRCpvW2fz6
WeOmbW03BtjPR4MRSjfbtAZ4vmR8+rozvhDrdFufYQ0Rr0vaWdn3o1+cCI1FgkWz
mTg0sGpYqw94+U+4Z+8XaZePIY1hQ03CWx4gVDo/jqfkZ7XVdoX7f42Cb/FxLeou
znGyMxo3MbYHE8+jcDdgt7Y4JxmP1iLygXXv/lIwRUq7wbMsF9WS/GwdwAq4Ql7G
qVjPnuHhNd/VBGN/6L5aJDPS7LoBfkdtlpu1IXjiHDtscR+57C7WL3m9AJyfgVtw
XVBWqNyZnlmkoT7hV9hSbliV9MBcCnXOO7rpV4CwFyp6OOYwCF3LqAOXZxbDNzf7
TmtPSkdV0yxDCXuzgFkMtq7HM9R1VUe9Lr5RcyZtAo48evt4IEi57IKhzJe3T2gY
Oxa8ObH36GcpFuSawFiAN9FhfL3hx4A0yLi9RHyqonYCYVgKs38XKRq2mnsxvnc/
2Vrh3gSYnfuGwWv24ohcmnBu3g5C3pSjlLOH0OilBEXIRlF7pP3JbLKV4E/1OkzW
kwz7IIPkclKEPeVwO2mUMcFSnOF+WGB30+WOSVv84Ki9FMKbn4lbBAruBfzRPEGc
bxptFOq6nlL/1/fyM9af1ffTx6yUO0sTNgbWb7+v5gxCJrF/xtBSDpvJVWTPRujB
C2RSjqQP2lMySECy1zwSq/mkikJQHfr+6kNQz+qlJEQQBtwkyDitWRXQFVJ0vtbP
M325XUbX/VFizEClE3en8V8Caj/WJiDSeDMnfBUHBXCzpGmbOPDKgIQcPVWe7fA2
oqPlCTC3cFHzc7uIzo6u+TQYYKDgI1jwipNnmkNDVaFTMuVrHm7NRa+Llim8xYtR
PrNuAh8eoesVgDHb8C9JZ+jRX+Q8XFpoQyocCkt2WdcJ8c1Wp4Byp00dly/k454m
uiE4iGsAwc+32jm32Vorl3rxa+Jj4J4gt4k0ksAtQojmtoKxo/YnkSg4oL4FVpT6
kqX7wehBGuR9vRWln/nmkE9/aYpvWUQnMwWZYEt9pYtYxIRiQXNIEogKehb2zakq
WlA+461P8CAZjHDx4zWJdCF+jPYRFjrsb125FCgjs/gPGW+tAYlB06SyqbNHm6jI
hHkEkbPO8vChqbhOuQhpE+UbvdQxFUdNoA9cmd6b1Gh4+0WdLZtZUCvocyILHpyi
nP8bDjcJ5FSQOI4847GGYuqdYb4sPiqsFG4q9POeZbjWhJkIPwfcJkX5G/g72zpn
dTDtzgbkVMX0nGRk4UVj1/S0REVZG/mnil/9RxiiAqJrZCs7Vou1g6DmNaolTtR2
nt3poZJDGxVUy23qvezgU3vhos1D4X2mOzy/yJ8WU4MXz38akVt2liBJ+CwoucEB
er7cXUP0gAB3MoUiOxmUZyB2blmTw+wfiPZ04U0SUxNqPJ2CgdeiTrHbnnJHrnEA
v77JkorhM20npLqmlJAhZz9BbPJBeas9PSbS9xYM8NBwU9lGecm8PMhYx+IbRg9i
0hBhmaCySS/yMWPMswgpX+EBe38zgYeEhGfhWprEVfefWKFeDk8l/bRtT8bw+OyG
khS8XsMJGetGe5Ocfgw56rHrC8v7Ls2j9ynTVxr+g9YRFkIFkCGyBq3JXI27QyLa
Yl9ZmNb2OeA0Cc/HnVkcmKcJCjsJIX99tCqM9zp/XdUSGNVgghebDy397vnrQiFs
i4uH6mINe7UhO/xazozhn5292Jt9FJMYahs/XFFLNd3r+pA/X9RVgAV9VnZ9ba0O
I3St5mJmDhLt4KmziApB50h390nH9OIaGcpgao3+5s52H9ZwmFz49JaH8wiNf/vu
TYPClawuoqpZAq1F7O3mCUjTX9pH/NrM4vNm3QO4ioVz0291zyGNlIcfejle9bOv
5WgOQrX+CLuSBXFicshPMtBNJYT98oHsrKcJ8Vq4+HM9OEjt80VpLWSgJiu6BVWh
2Lwr+h5tt2wP8EZtHAFVVv5bP/OIiCnClMiFmyZ7Q130VBHVI/1/l7Q0+034JNY2
R39bCLODsYho8tvfi4v8TkSB7wiLkfKkkkUDUoGa/GR2wxG2b4ynUs5K69owLLST
11ltF4R88pIM78vTkI7CJNo3qXgAwG1JWjH3MeC7qVa2hsgs1yzGDKiIx+6T6SUX
qA6oQNc93Rb/rkZVN2q5IvRN7Hk/T7zXd8eYUoBskplWgXgJdV+QE0Qpc7QMhDrm
g6RbY7GvHINbp984nQrTsy6jRBvpPAXOuLCIUvI1pzIbCNrab0m+yLXubNigrMFW
WmQl7VRs+vYhBGEDBnnfH+flNJi4u8nprUm5uAKVychakO5Vox+Z3NqirXa6PJSD
qpsor19hpSKXrxLz5OVG0cI38Cl2wQnMTxQlqr5YONbl5RSWcekREn0WNphQTxc/
OXAu9+XqlIuM5LlkEYCa9AVhYfvJBJ/yNVbhDuYR3XW4kj22/hxiUi/VS/W0yM5Z
TnHIJ6KdQbHQ6SXJTKTkczyvSA3BbALBqq5IhEw8L04Jb1szKkZugiF1V1TgHIV5
s8tcg42Prt9kGGxX84bzzzFHRS28+htNaAg5BVmul7PatfZkBHL15/aM9ZSHgwR+
RgI0v4oFh2HZJs+imDoW1bDO+FD0Gt/B52R139Loz0t1e1Of33BfazGwgseytMdS
YiIGN/Q25ptycZ8Y4vSNFsmutiDhvdnissNolN5BxUibi3YkWQpCwz92+YQe5ht9
r6sQxAka4AkICUDWhWvPOyDEFWfgrLeaGX52jrYJQGv15R12AhObPa/tSyUQtPEb
RR0tfIc7NOqo7isLN/fRjKzAzgp09973NWK8dR4zZuq+Q8adTagnydB2pKdjZ25s
0N7Ze/Q1B4fLlcaKm5JnkMesYs2G7wbf7wqZ0HijD2TgAwl2JVCjrOqEQaWdtJKg
xkI3z0N8fMHpgR1zMWpjbzvd737KHPL3EiGTZDORfl0gjyBJJoBG+5FKuaOqIc/H
/y6hPIZ9E9ctziTbTkvARCCQU+sy9ADbjPMR+8U06Wgjd0hK/BsbKyUqv40DZN55
FfkffkzN4W/RSJL89ktTkt1CfBB0Qgu25YLmjYwjYyG3R2eRlsij6nooswa8an47
TijMj77XfsvVkeva3Oi0th7eAK747/4PhrgnWuHgn4KZV79FXZaXHVtL+04+N3HB
ZjAsI020pJaerzdLSCv1yVyot3D3Tc6dsB0wV3XQTEDFQ1M8uT9PMwYCQA/UGn6W
sC2SaljFe8QcQYC1nOuNRw5iZzL6ugy2sPTr+Moa/p2lMP544IaIR9v9U397sNoq
LGt9F9z0HsVfWabxGbjs8J5qUJgqolpi5r7cP5al7d3iF7PzPQa87N9i5k6m7wi5
DRqh4u6ElzqOjdh8lOjazYuzKiqKOZkDcVHp13WozJcYnvyrzLI5CWl0qkZHDy0A
SsnonopfkfwX4AG2hAqypdBEcenB+dyiDwMVtTJcptmoB83C7fPfLX8APyBFOcsS
l+nxqZLqP+8an/nvoxLvW/aMT5sG8gu9R74V1HlrDEhY24MEd0Y6IR7AIZJvb4Kk
WZ6+jhxw7/MoXPL5nM6KMwjzq4ggb/g3ZDOZWYjBqSWNAp2YJaEyI0FzgCUNbtmT
R8sAkqN428oO8yx4/onaT5siUthaw8Pjp43L+Ne1lmT6s92d6hde7hxHL1i/y+O+
zeKXo2WiiGiTJKf6v4PaMPbUrBlBAbwEwWNAM2S2Qq+bUOE+lboEQIGS8RjEKVyM
s0JgCj1dfLYwJBjG6fguAVBSl0iUKgdA6hgC6qmfiff5VdEeOKNfyoROt4HLXSPz
qA2xBprL3Mdr/0Hu8ttEniIwGIRW2uSP6MXL8nwWFjEqNWcLl46kAF/JKnBsNV3w
SAth+vDJh9TjuDt73mTgVNweX6/TQzD7a7TJZ6OKdbvMNKEFDFhQXz2qnJB5q30E
oz4IHVPMIAt5wt8leRkoCA7d5SZMj9RChhQX0f+DU7rC3qm5xfjzDgLzTjzLAyl9
AM4cHBbNKH+QoXHS+kZSEu1Edqsqn2rWuyaHSXQrewoqwqyM3pOEgoptH4al9qtG
LLwBI0yV+lEaJtyne1Sh4oYwFaEwwJZHuB6MhEOIPbp/qffFPm88Bqn8+cphG+kM
n9B1PCkaCwahdxNgHzC/RKwsAnDTy2GmeJtKTTYYHzqextbDFum0IYq2IZI0LxPS
HyS/wOgwnirprm44TP+4GVGm3tiMVv+TAWe7mF5xwJkS9h1wMgYCExUHqTkBD3El
r6BvcOuQRsBv1O5qh3Ww6WxvXORBHHdal/vMS3jSyvof50GWwDSG6tnenpDJA6oC
7Ln8UQyLpbEH5GeznbddslixmPaPY0MQQr1WbJtvrAowVNFsMErcVOEi+ZdlMP4v
wJ5QopJSyBtA4yLRqN8Adk0GCyw9HXrzGVKj63+DP3A3hHSAi7Hr0bC2OvK7ARKU
JxMA/je3yEukVrT9XfurCJN7CeUoAmr6PJmKULxgb3diSE1ujZp/jgSbxg842h5f
lg/lMSuhbspY6rMwUCwbbFtHC3R7RHRcSdX5Pue5paUmJAMttEtHIG/ZoOYNYLRM
HGRrKeHGmIKDFZnPEGwpAfAaL6RAm05lsI+AkYeg/Ve/o/4KAYtHAKMcWKfKBWAX
VvYSUrojVqJdvETpKskF53ZmjTrpYOi69p4HG+/5lOlZAB6Eu2YlaaLmjFgot2lv
487s/fCz5cS3EGdQfSHlBL0ViGKiYTHSgzMKJXszOV2KIRMS2IQwsPInZGIIXbvc
+0uzcvlHIptHlr5si0o4HPKgdSkOz21rdDWMn8AAlM71ICPOR72+YMwAUxy2Bh1i
8O8nLqtbEQymdFz/E4F0hUQmvx2Y7G9BM8DUB74AiwQG3UQqiEeQHzSAO3Q+NiIV
fFzMToZ4cN43dTj32J3W1m9GuUtXbvTYUif9YnCsyLD9TYUntD1jLiNZLcuf1JT9
3rnFKTPJYvb25sYR7E8ZxTzwGFMEpikvmOIKFSAKxLu9gCXlb1MIj+EotUh4yfb9
Q0vT/luXRIZDthndA48GL0dBmKTDPJeMG+JGvPKC5S9EQ/07LvmSYrJOFycFQ32i
HlxZ57QZ3R/cBbZgJGECghiGHDCRm3rftsjH7IwI1CpgPXcs0EkreZZ2cTJ5SrwD
9tCjH4688DWDnZfXYOlagLBl8o538IORCBSxCRkVnNVaUfcoD6TscPcVGROxO/25
+y8WRA4qCd6v5da6nugTPLdW+8Lk4/aNQtevr9/CCsn6lk2JX5Ax5GvoXgATBa8N
T+NT+MIngW3WMnN0tJqNAUE9et+gxMxqAkh+Xy4Ga732w1H0gHY3R6p8f4Glt7jD
jjTscXad1iukK3squv7dABdWLWYZHyjnP1q9MQfa5H8vDv5bSOJspIsuHon3rx/C
+vQWC4NhsPsccgTlhXatlg1dSCifN8T0Q3DvG73wd1FCGxokctXuqiRI0Z5jK4e9
WZOGcYFKQa2NjVWQNiDJA4Pib2QdgiaItSnlPrwElmX4/hnR02jq/l28s6VW6TGk
tlP9vZVcH5CupB9lwW5h/6nZtM9OXIOye6V9yfWFMhdXLjQeJ5zryywx6dTdK62v
Y/UyLnyM4g8bCfY9gZ1vNwyKO8pjl/n7eQYNyh7zvemPw9zPf7XY5Wph8eIy39da
IbBrtlgOkzr3L0cZGsei8N3lvs7pB+NsAvzxno/L1y/EB/ws1EJG6eqvsUhkYOyt
zLHxyQEu03rRUXqJ2Nyg3hWe/lMjcCRvhrGHyu+gNvwM9Z9CD8pm/kwsnBed2InZ
WKTdOIqlvy21xib9rjU54plP6+2msgxwtTNTd9n5NqFaH3wNd846aTuUEaZQEgLM
vmFh+3w0W7COJ8LgXZrNPMF+deV9iE8JZF/UiGBDRiSjiq4sPC57relTAJIcGBoa
C12TH5Id4WJV9hl+jvAOTv7OwqdRf14s4E0lwY8NG/g5tQxRE9M3VWbRu4BejNOX
VN29l39d13kBlKOgFg6tqP6Jfsatpg3DLNB2lje9AoamuVSpsCtHlA1VT07/euP6
ct72q+OaCXhbM4G5ZWz92G8o4BA71ox9cpyNxM5rBHukI/r1MWZv/K7AbAfL0kD1
xdPJLV1/E+7UCdkZ5rJQu+5fR8BNXzQXldjjwdF1Forsx2Q6ycPPxXdD53ZPF0kN
I4RSiMOa6eHHbVD8Bi/QYNB7EXf7l6fO4VFea+CTUFUlmUBJ01L9Op7i3XFRgWvw
HNhV5VXtK5nMZ9tuGaa/WuyG95UttTz56d9SUqHwP2AIkOWU4TOjLLv3Z1+vTCCw
8dgOg/H79pah0fMz5aIdAz6IUdFlGH2OvGirmucpCwlZG0vwRbs/a93I4dadTx4D
f0Hvfe6M+VtXFog8WRLFaTo7G/xmPk9T9SqY4+a2oV2+GtIsmUDq9HjTUnjf6aJY
szUGP8RIKIrjajrbfwwLURAN2TcusN8GyXd3XhnDw84t2HDhPU+Hk5wN6LMsn6hG
yZd9bmfewxQJwDaI1OZliIbuVovj1GEeg5Krh6ZixCZxpLyBLp8yRxBzxN86Widc
vYctDowdpzthsGAPQGpEx0QrX8y8dl309Vlujv8QtNR1ArkPq78x1KnEbrsTIq2z
UhlTJ+XCBMiS50tKPizTsE6vMUDiTkFuTU7+Zc8i9RbeTc35ovjwv1F4IvyK+8l7
jFxREmchi2TcsGyTN12c9YADX9Fwl49MAPXOu6yYJkVD0G4J35HkAurr2XyDATKL
+tfe6d1TCMOpRF6WYOks6m3oCW8xVdFV64jl3w5pvdjgHOjw0HPwbP0P5+qQUPfG
K28D4kKL19G/wz6Kv1L64tnY4dttrS1Njl4TygwATPW8kmF+oimh8+igzJOk/G0x
Me9BweZQ10SXWod3rCHIt1MYyIvEGKRIPB99Sf+VqyBadDudUe0JF8gvDyJYISsO
zrdJCH7Ec/5QxAhxY6o3qLYP7yLg8ersOdmX6EVdq+9SsoZkHARdYY3BITjr+Ie0
1XKYo+NUmCAeSHnOERniqhHU7Vm32FpbIjEoXZB/A3EdZi/Uq90HXmg11J2sHhv6
5j1iWMS8tvLgHV9POHZ7omFgKqgZSTHHHXfI+MctaG+TdeDmrB6K2OCDQDIHkLht
QaMK/1Z7xuwwCXHXMeUerODNFDT9NZTmGvihdTUEtswHcCi06cUolqEvk9eot/Mj
74u+nZ3SqQNG11j1XOqVvqHid3c7YaDtEZ5YMPDl79VbJmhJRs79RZBYI6ZStqXF
zW0cRitlz8bfDrZoJKiLg2ZR2FtTwYWZhi+S6qSv/1gZ79EYK7v3XVIk+FccgebI
KA3lJt/hUg8KfICb6Ntbij3Q8zccOSMffjl0yLBWd6E+Ips05Z9wzJEl6eCIXP90
PCBYvWzpwCPJu7USLMK3aHQvQUGpeQYFEydrI610KHzBcFREVQqRsQnVtGT97/Ix
vigBB6yaVP1R4wEAat+Reuahtu0pJTzgsE+YETtV6nF4uvDimfdQvZ9LssM1AU42
g1WGy6Ft8WDGaPl/JXAu7WnHMEKbjZ6qBnki709lG87vbze6qonc0qLJwnfmkIUR
y2Fy2wuZx+UznUuWPxnXvDWHULqj2gPyhoOldW2ejTVV811M6naKpcRW/0ZsOSR5
1Hg8l4QYGQl3sgKZue0FMCFhTS19CU2qzfqyuVCOaU8fxc0d9BdCFgIctdwafVW5
NXmi9zPsmCITedy8T9oZKk8swYZjd+JSxQRlnNTENfSh0Y3rvGtNfNCCmhcuODTq
GQBmL3TIjUdYUH2KzCXVda7aCL2VE8clnngIL2iPMUcdy7U4Gp9YAvhS/CdWWzqO
HYxaPfMRRGOBXfzsmz05z1FU4lN96RSMGOgXOXzW4fTANqHQ6O74pPagNLiWp67v
q3STRyfQsbCbrfx6n+p5z8k9dEuRkNEayg+N8Ln17Han3oWcG6+hPz6fmfFTkjfH
OPk7p+LGtTwfr8DP1Ts6ylCEtEryS9Ps/hq8HulKC1jjm+37/Lt4Q82tHyKsTobV
q8D2kJogiR8rx28YF9rm0BfLmupeo1X5i+ZpOWIHbRXby4s10CV1JuGeSecWovwF
v3RXPtTpPZUQZDlb7nxzvv8TnuKERaCE4cS7POKgX6Pvaj6GrpVc+FXe4IdsSnqH
ovEdXZEUJieF8rIYAg3ITYXvac7laWmz5BLS5ytDOlHzRYkcptoUw5K4fRZjgkp0
hZhfmnzHHNyv/toYdiMLNwW3TBcudsG3dMlrv9xm+6phmU9biXtknR8L3/pAp0WW
eRKXWo0PMQ3O78VN4aONNsXP0aCjUbvU6+/m6xzdRMmJB3z8b8AH1YU2vwgHykfY
iUoRjkssVi86cu1POQtII5xQWu+LKCOcvDc6JcJoHBqAljSJUBCU6XsKMDnYmBWQ
+w9WCVr7wb2XZMJXC53VupAfgpZFmcmFgMStZmg3NudBCPsW/Ag9b18rESiWm9uT
YEPIVT8mgHkXODKYITxxVvP7fAKLngzoVUz6cgaSpPWDf/acfoR5nJQFedQ7X7HZ
wVQdhmQX5SMWojFYGu01YxsubRQ23qjXD2GrLilVjQkyQgrQu/9GV4/WRhfbR1vm
RIm+WUw9xW/sxfjZXN7D/B2WVpd4qK89PW376q3FGJL+LREKTfSIlROXTKjLg+Jn
Z6hvfXEw2jxmHTUyENSBWadY8xrEsRdriP3U+rL0cfz9G44qqVRr6PtO69Fs1nkv
eIiSP0/KTFWlr4ygoJa6V2NGNWOowakRQUebXHkhZjzn81XojnIgMzrwGi9qalUD
vD6yBFpRTQFIOJ6ig+YITOVxNsbq8i9Y88VpDFwnKJWBkLA6mdnKk+scjf+em5EV
3sXtNxzju9SlEV82QdT9eC5DQizDPMaRLH/SnZve1k6jYZdmz27vz/0RYI/p19P2
MDAVWYjvzvlacPRuv7p58ddVnG3+lJ4RH2vy/e6biMI1egurRAx86y13R6Ku+TQJ
PtcPbss26dphFfmybAQ3KFbB+MIrzN2P38ctSy1f3C0lb2CMxOvaus0z6m+2Pdhj
AYSoHk5vGoouYWGKNYblyhV7x8Nbdau5RN8gaZwa9ZmGUUIjpFckflpb+bwygBA8
7lol3opGiDeKeWNEk5xI08mYQ+otdt/bpb0+S3EKx7coiCVQ7bcxrcU2WMGZ5Sd8
5YFKa4EZcTqHXw0yzwBAAuqwGWVHqq6tQbpuaf1QSJO30PJldWWm6SQ0iOzbSuca
OTDE1mlBu0Z82hoCRbvfpaxAImBLWHzFrd3rN4KmwVwEWjYfweH+tEySPWruahCo
c4xBzQM+dTuU4BkICryN+IP6KPhQfNb3rCaBnaMmljkkXEWN08aIClctsjJiDIiy
l7N2wi0Ak+MECajqG3CdNkbzhOcoXkq8vi3sl6p8hLZIcBee7yymFdE1gjJW4UuY
t6sPcTEIxYasMgauUGc7/i7fpXjMFY06+YxLYWL3MuZFBDTL1RIEcn5fM4CSytJ3
zwXHeckHf7ssQveDWhc5iSnVNa12XoEGsmgHb6KUOxHJ4FHhLE9SLJJFmCJ3nibm
Ax/tsTF8MRBer+xunkITnScqzQWJTWgbwOGQAvXL7xSM2kqHibBBGtK45YkGvXB4
mIJGmK+Q+TvP6SZMoFNbDLTAqhgOEHkOKZ+4/BFUfbDCo9Xyhdb/HS4jJaOrpoJo
HAp/7t82Eo/sNLN6/ZWzqyY/ftvIIYw9uUQKXiGPTLo89zjNtknW6ps31G0mCrh+
MovwHRqMIgEA6DEMHCfMcH9BFl7Z1M4YxPWALQCx4qQEvfjp/lYzKzNFHSIci09e
NsT6YIAfWo9ZPF1cD38VIvWgM/a5+ekuMoE6rI3jlfB3moqWpa28VS4SpqxLMzab
EHEFbW1dVjxYAP1M+t7q3ZN1Gz7n6CIFspM116HiC2O8yx7gR+JqT3PrVd/URmSV
hGyfjxLOYBS6+XDVM5V+Is7/le7RPIsiKdFzEHBLCciCAZKImg3o0i2kz4iyjkwI
HfjU/O6eMg0tCgYsBCbcg40ms1D2pUTEpX3wVVip7oewg792+o2rZdsBxVpgtXVv
l0Dbys20IUsWgsi2S+wrmtzw2w/UbGjV9XlauBOG4V7o4qAy0QlnWggIkqovR86H
y9SRZIYVWPRElIwRDghIvnTmnhB4tjSjVe/GlAqyj8xrjsxnK9bzaayGvwz8eMo7
dje9CJfayFkMi1bvS3A5ly9j0bLSS8JMq9KBdIHp4NZ5f6wSDeA+3gJe1krpvdkr
pmaAYRlVOcz/QU9ZoML2L0dYP3uUWJOPpUvqZTTHj0/smzfQsmYRwpDJvuhjgmx3
P1c2Uk31bVFRuq4ymXXxdrgoFLbPA7XwkPzo+fBX8hy4/8zxnfPL8MaYUiIK3/+U
R4jsqO9rtDZOyDcmIe7sXeg2Fx5DJ14H1anJeSXXu8rNu7wAKhRnf6YnV7FweKoC
2UnubdipD2NsHBquDMHCgmPuOzfvb6CT0N8oHOoBg7zaMbWb1S+TUD9ooT2Z/PPh
SXK6eE0JkPhdX/mDIWl6z064v1YHXcyHZemIi6ZaZTJA+p+lqFiHWF7ULYzX3/n7
wpSoqFPwadj+YFaQkVUkcax6dnCpDzp3vg9Ya3jdSqDXymuABOB6tFgQmMipl6QU
LP97XoyTvr89+cX6xi8nOiR6wDKrPRK65jCLOlg8o0Nq8i9SjKTdifu764ZIBtoG
6Ee8DF9A1oENQCIaJYVxV7Yao/VKcy7WSiylu743ySdCaVz2eH1xnjVCHNuxxm1x
6DlJVMsj1Wviw3hjquk18eqou3RSdId5/1jj0Xi8XR1YU2MxI+dGy142tMa6ljtt
Pp+BmP4JhV6sjv0xUJu1TbdFOF4h/Ppi05FQhHRAw2PkUZzM6ezZIRRS6aEXHv0S
tJer6/hPTgdg2u1womneGcZ0WXLCX8R5spmMVur3E4VVzJDHTL+lfZ5TiYDXI+Bg
pnz9bIqBuiEC0zEUf/L2xgEYTh+ytxvkj32JArboLEFHKHDWxITsjcxIh+mK4Sww
7blmmRV0u8biNnopjoLqnEtaJY+oLBZ2MG3MlQg/Q1IyQmxZDfYazYfdmxUtSumB
k9ts4GjE9YzA3qIqic0TtZ68JS5AbOSqF7irO2jMlilFHgOQHqLOmtaRstJsYgX/
UyrHstWQnn5kS/EsnnqjERk4uxtytIHEyxkLyiXpA9OE5b4v1ET5RevDTv/7NhO8
ncMxBexOK1vyO3c+RqEpea3hZqXlnzqeEEnAFdheTPOtU/eM/fSFzUGD4YsaFUfI
NIOozfJYYJvlHcfETmQJWW2FEXvj4yVwwX7XGt75P6KeqXpg+0kkaV0cmOQRSo4T
KHFPWPxIYFo39oIvlfKrhZEuKtljIQWpOhk5L+EtDdMSlQN9ncQeoGnMH90Oapeb
XzXaNZXAJdF/UYGf7FhE6gKOcg3HUslwYx7xRqwbUKNq4NIpd4m7gyaasO20rwFI
BsL9nHFAcL6aVhq00pO9d/xh5os4rA+BmhItIj7vd2XEw+lRqqoYRY0w8HcC7+XJ
1JMnznv7YPmXcTCzo54ec/D5Xa74vmnPQDbpTrvCLHOah7H0r6sz3cwPcSoJUcYs
DHw6Q4jSmDu80X0ZhdTk47Z5yjjN0x1aieQ/q4cPlN9RfWATZB2hwbFKPsxeeec+
GnG27uzUXBaRrV2vett7pB3rtUFemVtif4x1stICBOqx2B8siwHIokaLhewTMZHg
rQBLnwz8hjVmUUf6iu73s29DnnFEhCVk7nIoUCcck4ruNUkEVEb/jmRlRXR9L0m8
zl4PNH7NG+/abzu3+Mm/N8NCteRCika0a7+qPc51ImdpCyv1t6kpgdvMnDZdHrrP
GK00wpdvpZF8qR6nUpJph9+61C3LkuLuXYKwtkin1mCII+ReMvXxfPR2XDlu+SQJ
qkxGDXRYIvS60cxJpEtSJ/3PBLFaKsw6wRYgMpGEyWHnSj6Ph7uVuGbVInvgtNV2
QQGeGfPhg5YneDqDHpQpBFDJmftTTjve7Cu+GsNJxGDgOF/vnHWf6hs2DEflybOB
Jvxsx1ZOX9Ca7pmcn+KMXTY8gjTyB3wJGB8MTm7hFDZ/yAd48Hgw28Uycjzcw7zH
65C8PSQP3RL4LWrB3E5GvGMWYZEgMpXMW37vJC6ZZUFEPlrGDgcGDYBozyLUFXxu
ddpIaXmlxYdZvfjsHGKrmqqg4xMJYwcD6ePQ78L6c7qhctUV3elEOqumBlOa5GMr
odC7t5vmyt0IyUWVougy6SdX1SaBJqNPHx8pQc/HDm0YEMBGq7zp5L2cviCF+1d0
Pi5zoNPmt6zLxJfrAREmjMGdtNyxfN9rLNaToynf//BydyKj1tnen1Bslg5QJ9xm
n2Gn1zk5jmMKRJO/SPLGZ8LnR8ye9jcpKYtQa4Bs6Y4fpsLyXV1MVkdfIr4ZKvAE
fjb3B10If136mX70Toe/Dor8JvQx6VAQJneTJyAugADHl/GBO5JgciEN4akla3c0
sKce0iGJNfnT66jVf7XU57OJD91BxbPAdNrjk8qe0Oi/goDTrwCviiLSBeFWh2bP
TfnlsT72PilccYtaHv0zQoA1bD4pCkOzRzwxAh8uYDtHn4NneQVg0QZ89Cd7sboS
qRnJsjTvbgr+9aj8VrBLSzKLnw3d2L05KwBZXZ1sv13tRtChsqjrIYP27o7fSqO8
bQ2of7AW1dO7W80/JtqyeMAkOWJ6QKe6n+tkgMPXpvUE26kLu3KqXDStMHnuwAeX
XJ6iSToj5TwkVRc/0Jo0OQpOjzVOC4yFwFBtgCFTOlkBhvA+EjfBbtERs1OuTrV6
ijUuEp7vP1I9RT9/V5YWzu2PVWmqGN5dwfkSaGcBVeLIy3pcOPROTU2CBhLst5rV
6U651ATK6CvfnOLKfmiJ69ND++YU6fyATIPueRqSU11Dp4iuH6ZOg3VmZlP0/0PW
QGhjIRWfT6AfwEiVAFu9nsPjlBTszhjzd8RD5bMCf+xJchUR6Q1nWeckD98iRiUS
awV2R/R69l+5KySIa36RqiEZw68WUnzevyiV7dYzv2KfH2h3qVUJQCawdIE2u4cy
zfsVocGkteRaSgo+0rZPOp+38qv09Qv7buPkgArJuKSPmxrShWW3icj61OxId1g6
/drJ668JwXeJomtcQRTYf4B+AmWOIq5BKn8dDwxl9VbcG4rjeVess25kAUVzgaCq
0G9FpWej+E85kfKGpUZCqFWqZCOXgS3w90weK46iciMCkhjVvGFyU6ZXJRlqQLIu
9x5dBKqPu2NR8Smx2pZycvOi+tCsZOsUvCW76NdO2b2MLHDeCnZUaNRCZzX4QKT4
3/U9Ho+enfAFRAxAHeh+N2UB1xPrhTMpzY4ga61ZXWeuqsPsJztwvQgSLeWXE8Y3
Gu1m7Srvp5TLDRXZn6PGVytEVuxh410+SoYamM7MlIQ3wmw3o8GdJAU39BeDWxNz
npCvA/nk/vk4f062V+3jGvGdmzYXvK/sLHTvJhwcRMHyDejJpqMyVjMg5aRrhgcG
RVW8fAYxcZPpJTl5QlwX2Q462FkZwDD4YA1KzeOJrL4ya3/QYMMqINg+oJFrCUB4
pH/PCld4a0nvTkVrxo83KosR8NVTRrrWUgtlxErTjWMTsIyc5WkseXg6NW0qIMBI
4cRLgUChW/gUjeqZ+phLzm1Fl7JK0FAdCHQuH7hofAxzN96FW3fuYC2r2YPeWhRM
T/8vygfM5Yay5vdRzdfPeTbGgO/0hHMFXTf+Ma/WNCK0ISsJa4XLCnF4SqFnamEU
w0AupNrFK54jkO+/gQVKrDqgAIH8enmI5CCLYiPfrsct1focu2fsmhT72Y8sHlee
TP5zKnmpuOMXHnOb51Jcd3lihotPSuMgBFdUCY5G00ZorB3aC3//zhXIw4HX7IEL
vCVcmo+Md2ht/evbR93A7unxUg4EE0DETXxQfi97A9zTLSAl66HXh5mOxJPffhXG
UxRkGoEqzGJLANKUjoJUD5tWg0lvnnAqCiyLDnYtJYJiGKABFugwo8wqaY9SKIzb
kJhgF8ANBcPMD11g2NOQSxml6BRAhaqZbrb8fIudqtPBTHnzu+v5ioLkHmih4CKq
WYqycQvxplc/ij3E1u3U6aFCvZ6TX2LCr/lGbrLkP0Lcm1n4cSc4pB/t91Qy3w8K
w3JfgJTMkRNJUJ4XtFsi3Q8WKTFsYGfpWyDX8VCkkDbBT5V97QipoaDEOE57E93B
tXu2LfjioBC2lqnYVO/ZCNL4i9dOXpweeuQSEwkYlbkivweJsPsZHS7pizdqkHmL
1apaivB6qilI3Jx97THbxX45lai+tTAom5wbyp96gBn7hfwmqRVFmkRekBikGFXj
2r1DGe/17KlK5xymSSouFd7EhIqVdVkXWOQVljPfQWgDY5IPbEUm/a6Czd/6Am3m
UiLXiCb/47E7dFnAgBopfYh68fVelHljhNCZkLr4TEh9NBjEfc9oYgCFN8zocQt1
k3eVZTt5b/SVJHzPSr3XzWzSAFIAYUKQtNInWYuSnjrY+L/onCuJBD5F/9YRiWAi
DQLdiEG5LwDf4by8kwLxyjAO+LSzgw6AlyhUqdlSPj5JcIihfninEEitEB0rKHAM
56JsaCt4E02I+LyZVWI2sfaEX+vXNAnUydIpqKbQ6YtIfbWiG1m6PxEQQbeyo9hf
fcRUXi8FdTuh9FPnn1nGnBpjznPpML6okJ3293sSFZdOWYj2Ad/SKmBnAcOZv/sF
L9nvbyutmB4cMC1zJpedIo91B7NqS5sAaC3+/+DS3N41WC2FOQEbuzJXibYP/zlH
2AFQAzgLLg2h+9pxAWgUBO1gSAfNlI3T6XvvSGr6gnHOZ7vY2xOiKuGAaTV97iUb
jxuNVP2fhBmMl6NCf7Z204UI94DQDjG/z6gLl7vOzvpEBO3juWawDccw6nk6yei+
9tYChmyTm/1Ne8oypcIYmsKrPxOIqHIF39l9qZWrPUCkprIu9Qa9Drm7AEwi3nx7
qgZaXF7r5O7LfTqNJYY++LVx9flDK6L5peRpDrj0GR+XhYkomQdkV0ZQzBPVxC4r
0jGfkN51sVqaHQ7J4O5xMB4Vs3/7UkYkiQKupXLUN/FP7Dh2JHFYV6+r7v8uRVgh
RMHgxOpEGS4ynDFrZ5tct205X7mL8KLw4xeszBmOZa9yNzB7vSgdXDVNaJLE3NcW
2tvP4YWLn+caUfvKPRBf4zEB+jYnOQCGYujD6nMXeiIWuQ493igg3vrn6vR479KX
cIOpQDsG+zrrgwR/HFwYlB32lOHW2WWjG4ZwpscJ7tyZYo2HKuyXX82OV+v37rot
CX/hsIrg787N1v9dfYeswFrwHxPMAVkBEkvLTKdN5UiQT9z+uZS6jPVtla3ztFnU
toGED1O5SE2QzPKGhTYuETHt57JP27Xy0Q51+oPsJtKM/MVw92A92brdwIAIW9hF
fl5TGv/tqU30tjoqtXCYmzubOxv3vqXyG65w3Le/PQw5qTbzpcj75EiGba9tVQg2
Jve+TGSgQfXTk3H3/6mHHEFE4j+0Z2i/jE7XWYW1jnBdFANPl2SyP0w/fX1odJvk
92IowiBdBfiK+0lKS8r6QVVNOrACz/ZB3B6d2dcxyRT5o9fz8IBu5QE6HPO/x9jZ
CGvioWX0Uq978UvTvfQgsjRil1TD8OQLDULt3aSjPop5qUsCcJnUi/KksRnQZFkl
/iqNOe6jynadtVVKiMCe8/9/GGFBk0JosDt0T4mrj93SrxwdoXlSc5Fta6uMv70G
QBg3XQZkUX1+/2KwjlDnPxg9y85bfQ3hYA8Oqo4PacIopo/bjhjWXfdAi5KzTNLx
dcglyU74Sk5js/f0aDEP64UeQHgrdSFXm6axzPatadnk8qW/AHGHSnGVI2lH6aqC
MvZD/JdwUDYvibiTeZQDLyauFfzKM8fIg9ZOsXzH+Dt5FDVCRchH8apotjlkSzft
TiXCqdij4pcOitwwyCOnPSAQ7faSL/1ZKx8+wqnwSfKqNJhL7/Urqpt9yCBBGrnI
mf3WdfbfhJqLlinbCDFDQG/+1jdm4mRMlzEUzmkXW1/mIG4fj9BxOUhEnL1klijB
U3TIxt64rwMVGDpFL9M4MIZtsXzKcOi/3MCjfqKcv7KkwqUi+2lLa7Eu/vg0OTX+
T/s6cArIXVesJM68ImtaPG4rQJTENz1xjWi8WmT+4qkb9MBOHQIqyTZHMf1nXTMQ
4Rxak62iVnRKAJjYqITHHVO7xJTUyjv9/RrnFTHxwQEGY8J4gfqEVKqE52XC2d9q
5zMxgG/zAMKBp2TgwNQA/iGdpldCv3BYo+B6vt2QywFDCT/fRkWyCPtHIql8qk8o
4xhra0q+vR1H18VydrdveGtEFxembge0NibX6IQMfQD46vL9GJwmeBskt6yav8iD
LeEuzo90ZFxwx0XcGeJ7MJezxc4omFpGmdZW5sSTKu8MI88KR5Iq4tVwp5mkqrxv
ihl6M0SBmvQvrupujrvdbqLaqegmjcxtsCoV3SOrzyIFAmMPdUChkkDMHPvMTAF2
NHwBHs/6NOmekqiz6AZfkCrfm8Rakaa6eiDTnM4uZlBc63kheHm2+jzqo8CKhpn3
DikQzPNM8jQG6b286VP5MSCd8uyTT4WL/9EGgQIp8dru/At25RmOtFqpk0UaQUYK
/OWBLol06x6gi/ZWs6BM9grgG6FbGUuj3o+4EI3SKuVUF5bHzhlaJdWiQKvnDUKI
k6WKOi80t1qMkrbR/2vwe/ENzK08EWNO0ksIwbPiacAoomuumZ7LNTwEDD/ZVSCn
/7addx9k2fqGLyEqbW3yNmB3s6BXkrYLtaFRw52HH8LpPt36SiYrJYjfMpK3knYC
dtOJ53f170Muq4SqipnebNtHgbHXVZCrD4bP1nG6wYVPjHZArG1Di1voPDMrMy5H
tz5/Q/WYnUxz46iLnruIbajpMEL7MjRxbdcll/iJbK4i1aZtzJuVySyCzJATipss
Daie/jZGq/a7tkJnbQsqR47MUZF22NUdxCMnaik7gdI6pEGzjJQ4cnBgZpHWHPYs
ZwZ8GgbB+N6+/s70aG1vbfH54Txla33rcmso5mZC879iWQN2gKnalSELBIxaj2GG
RKSAK1hm0mOiplVIyq2yjVk40+Tl4lbc93ztsxFeNsTbWLGcAU3J82o9mzLgjiwr
ENO5NpyXONmMw2ovv2RIkC84uY36REtgti2o9QTNVOjZQdJwQcx6ky5om4dXbhyO
HduxMeHoxGway2gfcZir4GP4NlRpzdqx58r9w+UhxTaqkkQi9IN+fS6UZIaeHfK3
lzPWoJvP+R/X+4jNjkmZszpPtueu1n1VcVvA0jsabWKd5t6b2EHnaCB5ljMa8UN2
AU/MWuwACToXs5UEv7du238fEftfUaLkQk0U8rbHrDpH2et8lxu2I4uO3WXPZZ4V
AhQtyDMxPKjhZXljd+Ro9aunwinFR879z9izAfYIfuUZmYnfTr/qWRrDrPEQgwBW
B/Xx0GzjC8ZYJwJuvhDTvKdZRTgPdoNm8gKnXCxo2Da084PHUqlnoWrj3w2WMHdi
PWuCe5qqQLyoEFhv+Ip6eVu3Bc25MxY/uPJxrHUZtXHNiSY94z+X3W0JYbbgFtWw
r1r7B5qjbJOcVXdDCFpNoWBT9PaoLk4hVDuuyjG96jYNZ4pGFY7AZYIrU4oOiQzq
oc/eOgC7G/9z1FYiBmrroHRUcMFlvWmaGV38O7k/Vv1vJNoDTmRT73M+BQ1yI90q
IHl/hsAKYq4/u2p0t5s2cH5kKI3FgvSuroYsaJG7lGfI8P5HoF6JP4XEZnWxrphC
fU973WiKVPqz6egDilL/Nyvt6mhBlxraSu3iFxiK9t097c0YtWDDhbbQWGlxWBlB
c9jg15Ng030rZLKsbPHuPpOtG53Pw0QMoGzx5+LOkD1jLN6vsbsyEHxExUHXQnbJ
Fiv6XtxHlgQY1oWxH4b3foH+q0uWZcUVRLmNoMBF4Mu1ERSy31CdnB51PxXLZMDf
+gZ3mzkR3fPlzPpgq6TT2Lt+4QJrpAo2lPsWkDQWNcZyiPwwIbp4hQb50ZjrIiRR
RJmoJLffwNacJygNtunA++6nSwljC2iADWbZ0dfeEJ0k7fB5hj7svnEPy+IPMVeW
XeRFlJzS6057/GOIID1kxPqOFpPevAK/OeWmuaf0SIUbRv8iqL6yxC6ER+WXk1Uf
wkSjo0MqH4wHT5dHHN23QyCbOhCZ2aiVW9Chcq1KQ4oqlI8KrISzDNn0ouz3OMyp
9Bcar4SlhsfLN625ATLnMOQ42EycTrsJwqYb44XSUy/rYpfpeRuoEvM/I6GVkZkF
3PVXDf8vSCtJwAgREEhrzFeNVQjdbbU19sXhSaBurofe5fo1pgeB9BF1bpwf/Ohh
xBdxJL/NsJlJ3pRmRS8vQHjo60l+ILfrIoBT5I+OSKzeLA5wN7r23nJoZZaG1MsV
44xskZItSjiaBL9+Z6ZJR/8f9zCsksbgqWipZHJ8QCM7wfoIm1/xcS6jlwHXIukb
uE+393QuHu/aXNuMD3AriAl5ptwKzJ7L45cl74XAnW8+RxYomShAp5BxgzIXNZoW
/cIhis/QvoqOBecMeXknOxjOHbSIvS65bbUdQ3o/LaRyZfguzrpgH/o0PmhBnIOI
FgrUHhn589jL9wFVQqxW/AkMhb5A8N1yh8JRIJX9JVw8Oe4E388WyYa6of3yjZuP
0Cc2tufd1+ZmjdTXViCZZLVZRiop2k2eOI/k6JSH5Qq9VuBb6qQkI7+AqmBeYETn
0SN5ETs4mJl6nX4zJ9bvJ1OFfSTUpx4cErDJ4iJiWwMysHQv50yq//WKq3H3YwVp
ZsMHbu3zaYpBsompT7piBys1n4XY8slqRzNRhUwsiq421zkWNsen6/H0rvfnFSOj
1Oxk1gAYK/FXD8KqnRND0q5mFB2Wlw6nBEzycFRnAPXrHDDXJHOQb7JeihLGFpuF
VQFgZDxJjAbJHvSeHthRn77SJ/PgaE7kNLXqSO0E7oy8ezNeJN4rdFIrGCQGLzM3
xNvCKJyqjPPjVfVFq9QbE1Lp6pVj74hYRgkNeC2jmHo0s7lybG3Bt2GZpliYGdUs
HCWLT8UxaA796kXMRva1ZxC/6HeK6o+WbWyVaw6Qiw0qgn4k5F+x4nD4yrVTHGah
ngJzohvuN0ihwpp8N9mlEOu0aKh8vc4yVr4LwB/bcMf2Xyb2AO0lP3fqtdhdD1zm
DzrtRkQdn2ukMIx3fHa0BvmcDLbtQ/Qmqy8QF03hxrobobSlKd3oxdzt8ucbMMTX
nKO/MSuCZmVXJfr6mTM/TFibIAao9N1Vr8zi+jfSUL0ud2ZfVQ2imRQI+I338wgK
SvHtGsNM5oWGXl90kwPnY8nH+9Wghi3RoXaG3JJBCnaDTKx929i1cGOofQScO1n3
nWVdHcX3pFWjbDg9P2ELFo0oDVCqb/fsT1S1xmJOjHCKxgn/MCVyFIXy2c9fIEGR
0N1+CrQiKnu43mLHSf0xq+wsdbH/NkwdNOUkjeCNHkJWrdRYaR/pkXWz0ph/zIe+
BFLTLg3m7DjuFvTPlx/6qnV4jytb/u+oJIRSFVnBdUo8haFvrPbyLDZudmEq6F5r
9JV+ObN/D6kWQlb8SreJTFynmWLGxxADePinVofj/dw5BtZf5e47H/FGwY7i5eho
Xvzi7+Pe5yCoSQYzj1h13A7N+PfvGiUn9NtnNqHxwN0RoqYMWaWRozzkoqJaZ/IY
syhdPKMAnU/pzI4esw1dsgkdl3turAeXS4XFek6CdYuDh9AGwikC0XxfNzBzYUnD
wmWwt7Ux5Ree/MRcL1A9T/zXyac35rFZSHAQv5xF17DRZRkpRvJ+y2zk3MUJksXs
L2VPZhLiHjjWNuaBdWQQtGPO/OBCJOHCwhRT17kJoaWFCmvxZsb/QvPbQkLRJw6x
VrlrJsmdS1B5DzGsVuKh1L8EiqSGQWCgsW1guUEI1cBX21cOXMWNVMdnLkuM4q5S
tnTggkLJZMPNHLbR8avz80b3BkhVgO59G7c3GWDmjnhjZSqO6tB+2WqrV81WCH+0
3RHFug7teP89qvNgFV+vAK/j9rNo+zG/AUUO3QLUDsJEkDEcO5MGOjmbfkwkMNWN
CLs0WUWfGZ4ONQB/bAPYUte3qrZKT/U4V9aUpTVDxq1KL9Ls4SG5cFmh7xkVUSD5
xS0Pob4pcJfy6qS08oqWot/ClU0npnMWYBqnusRr5wutkgraNAosKp5YlDswYZ+H
f00Oqa1e5H/udewI5Rw7sa40q2ODDD+ajn1sdr0PogFeRiH7zSNuZ/Op3iH9jHeh
ImVspWckp5Ktw8f8bhi+D02ix2x80zgWgcpGnNauNsXBPZ8WquxVloVtVShmGrKV
BWMCRnZHl6Sozlo55tZEOzwtFcQm9UN1SoPFcDQkB+OCyecuA4Sf62sVOOwkoSLx
JmIXmkA5rydN7NyZUlyt7Pqg3d5vv4sPJclmOwwuOs1wiIf40jzvOStFwveXnue+
7BufD/i6YIc5x2fdM8nbaZ5Mpmwed76Hrd7/ouGuS3qW2xRs+K8rRdco8iNzgXbf
rowu0GXohac+RMpwf1PhAL9TToilVWFUTXcL6fAQfikfLYZgbwFp3fFsIpxZfvNr
z8cWD7e6HuKTrji4vVCKwB70hHRcYKYJtVeFShNH2x/37uYWQTlnKEtGhjg5RRaW
V+1YqUUMqg2Hrgax7cqaJz1TnnHQRM+oQvWyfeH9wRRz/KjDAQwRQiOFSX6zjfrb
dmOCrzjYomC1dXtVR9jodV+cOrFJW+xymakfUJA1woTa0jOF+vgkcyeDJr9tIXrv
U+CGRdqWBPzOre7tUDTG97VPKTh3CmD1jpq1U3Go4j0P/PXFL08tM8e85iT1nGWb
MOkhRAwXAMq1tIC6KVkdXIa3WMYirkPflAU8BL1rzosDw7qsPqGsh94zT9eY/jNk
x+64B3iRvUAi3dLQBkahuFCXyg25Y530O57ulY+nHLExGVXaLqxY0hynrGHNk3HN
vksCwpkqhnKW23u2DSd7u48XYStntcXLIL4twu/fd0FJtbrjQ7JXZwrTqej+LY9S
zDpwq/DnUWA1zLJuzqahTEQhyiC0cPcnSAbUKZLMGGwnskA0Pblfeqyxnj0sspyG
UmQMp4spdFD8+yLAEWsyrL/rn26okuwwnRB8J2qjFz5cto5ZvrARPNm4pf7Gw0Q1
xVnkaFESAWEjg9rOdiXnFM6nPVvelhXBfXfinrO5QurOQJCso64YNwDrdR63nAv6
bcRqMegrPcCn7u4qsqwcTzjrjFmP034BrHA7sug83QrG8o/zus2OCAsf85nyfuaT
3DTSVTjVoriQmj6g9i8bZg4XFCEP/3sEj4x6Fl+C3AIbJcdBSrMVA++VpFSInS5h
Kma+kzMAyjHXNMnR1hEU5alHUA/TuHtAuQmoiLaUiN5Umm2eYpAve9ym6PK/tTzu
MAdLclIKoyagcAIduip1gS3Q6QdQpWTf74Lm/XtdGQptPXraZvy+xxEzBPIn0PVM
HtckJQIbGN++N+XE0tuqxW3O4tTIDR5xI/otN/6twmshDmmjJKskc+PlGtzwZxxR
UfPSD5VC8wL7DhHG2BD3v2Bl0Cy/Ui6EQQob6p4KDyRNVWR2lAT7y5xDW3hJVJWB
oYdz84XDmzyXpyUCRiVtEyx4IS+xf2TK9oPsCis3Jp8MA1DVn8u2NBuHq8EPC0gn
DACxYZgX2Z+vRmlIheC5XtJRuQbO2I0vHClQZClsz0Gu4Y2TH8Zxzar0m5Hlfe7g
8KtaR2ztlXrhYtmxV1EtktfFMK5XQA+mu1ni8Ikvj8uxw8ijArCoPPq/H7xHHtDM
Rq3/2fOunccVKGaX0razVnGNqFz5dhYG5weJtvlt8RvP8ZeTqQ2o1bXbbW7uCrqv
90EUdjmgUQIbraO7P0wz1IuB9Qh5JagCSBt8jDpPFQwM3c4lOeGFtZoys6K4OtlB
02flJJocmyMui3gs2DerA9k8dXWTM4Hkh7kHtFm23MkqyZ88ZUQ6BkHyP2qTMWgQ
fq2h9+qqiElJjaRCc1iYCQJOjrLTeJALupeY6mT29jOwxxxEZvfvdmEgJd2gNqow
3wwIeVxdpGBDyOVvNo//hGwXGqr+fRKygYS4S1rFiqB2zKI/m65CjEDDh7jNzaoJ
wSRRvH8YuluZJTDKycPf/DqedoxDGQTLqy7OBwUYRh2GDqwo4K4o4aDdLllzdWJI
eLxYoM4P/3u1FUD7Z6ylT577E0T+hBGV5ZYxDt5nWmWMoLIXxlqbS5vayloPmqXZ
+cV8Seans9hRRSFc9z/HtfrYBQxqmX/JYBVHMZjJM/7lCzz6ZlTyQ23MEFJpV3pZ
ADtqmC+9VFVzLzlJHbSss+/EfcCYyh0PKHoGEnewbx/WCVCHgY1wXRAsQpFNjY5C
IpjerDzUBbPPIwbwkOKz+TNVJWLGX4rWCVW+n7nJqCb4S/j6iumAmNlo/vLNbuJ1
bzlFTOWZPGIydaDZlJwcjmo4JMnbVYsToHFgXYhfxs+lYWmXdMppSWDPc5Lt7jSC
hDMAOfylsCPkDnM8cvKuW9WNV4jxHYWiSOFxTnPXClPiPaNEgm3AyjcaOkNbfh0Z
f8Bwhn98BvMjN3y73AWSbKqzFK0sUHslZfKlaQ1T9eMjB7VB4BZCRZwjPLVRnUzI
9wB87t32NdL84cpBAA6FAG0RypQNyuAfoKwwaAhYzQCI7gUKWBUaTMPC2qaXOcly
fCxpaS7Mi0MCUXiPn7NBLWkrwAAumSqe012ZGD1/qLjKpSS3HcQFHglF7Pqembjo
fxdqkP2zjOHB6D9ArE0v8zhemm113NqWR6EUvU4R6MXcdNE83kzwK77vVeTbkWfN
FWNyznbdT7J5tIsedEgWfRQuC1Ewwf4sVJJAsBu9VsEJDYcVT9KTvTuhOnmCbipF
nPiajJHsXxue1Zlfy6T2gARlz1m9qKW7zEedyZ9l9DFnPrQBkno7PqfbAKbvjg27
oh7fR+pa/+X6GC81tmwJIz5GRxuV4o8cZ5mU1i8uKwAHc5X1SKtp3VSkxTG9A2/4
Yap4O44skOktnxfjt1ewZbsENfimXRcOJf5twwosvN2ao4JgYJV/+xoC7VQK5oTc
P09cr9BBzA/oKH1C6iye+vhF9idQ28xExDJsmSQOgrC/+PiExMc0v0uDHdVqePT7
f2nMYPfOXnS9OVMDt4aUAANXtjHOBX0ZGU0hYRfmD6npe3zQ15e0gENghkdiiCyZ
h9PCk23bLHKenpPQ5E0b6hEuSwtaMp+P6yuvK+UHJh91nII74gaE2kEALqAyS4j9
XV5WhJm9AfoWLM33ele8FKiSMuJAjGrHGqRhTydtXGWwRZYL83ziwLYuwLzOSdWp
L6Peej14+I/V6ll9zsQ1Bjuy1/DSWjXNDgFjLVLBZgddwaGXamPgr/aVqyR6Q9hn
pSlBkf7VGZsJwmHeDmopDdfAlISJav6pBWOxf8y5bM+HyvZVi1PquR80pToPDKyV
GxfAvWy6R1y2ioBoXyPG6KgoTKvuk+ETsodJwMod+e34X3+i9B488ilcBkFolb5h
ms5Aq1FOnC1P09sjIUkJiYeQGsIKxNzGM3a3CXznOC4FurDau3qbwN68rDn+MMH+
obozc95Mr6jESKxpYpPPKjMcqI5z8wQlib1tlagVngtHcZ81FjQrBvsHyjmoWn5V
RTFl2GPdpn+Bz+9uE9W398EI9pynM3+zXdXeND/xzGQ5Jk8y4Pw84oQZ4QWkEPNA
f0igdUOBQDYnUjNH2VWtTygKFpkrzT0G8ElVkWgdpqXO1iJx0laY0zZeR6obTf9I
l8y3xMa4PFU86V+BFSIDfue0uO5iqtCtk9RscyA5ILSdrtTOokjG+d2GydQG6GkK
9jAONqQXxZqLVgbf1mk5/t107jsQbijOLk/+YxrYNIZhCJxjDKs18mBtHBdWd1P4
BEnVpg3hhLfYA/FNetd3fivQ/QIPomuk7+54jWaCsZa72RaF5Kd7wnICu1P6ceT/
9UhPgRIAmMRRbiCnBp/xUehvcTUw3e44hDWlN8+7YDnJakZypqJNWwPUzR+m8wNb
yDk3BAGp38/Yg43Bz1pXuWroGaLm0PF3BfwDQaW0ayD+YbCCGEo4KaoLwnXe7zZd
MhQiXu3TusSlWx35avnMddpyvafiMPuEBsZ9TZZekcG3XGi1eJapWVtO65wfdZYn
DT3m1HREm++bspoW69TN11vo9ITmO4m5qikI2pSiIjbdKtivgXC03ZZvpUUMgx2H
LQf84kLoVzfafv3G3oAhzmkrOcKqODBWciLbWOIE404f9Xah8CFj5v69kXQlYygC
jPEMQWRtiPQwYmRPfduca11j6ZZrPWNhCRkeOjg/8VPNMCqcQnYamJ6u0PHxo3mt
bU/jwhuGon+mtKrjsS1jhHG8EGl5aNJzWGRO8USI7W+H9D3REhY4US054HJbCuSC
RsAPsyhLd2Yp+e8QUvJWxVYXqiOStVO0DkIBvcLvBx0ImHO101DmP3KIpPOMJ5FY
N+zZRfMXNPZuewrUULSu9M3NHxaICEb0GCtAaCHt+UKo+dDVMUjVYLkJipJfIPWA
XPwn4c+ZVA/ofrXtUSc24+0PaDXdt8WqeGV5cWZwJPKtFxlvSdMwrQr+qoGpi+ql
aJSr9dq9voLTf88me0/HPzdvSngfNERyD2kwUIg0Btv9xpdFmkodYXL69xp/mxLj
C/ArbGuumYqWkFqnXnNJzjDWvQLuvlG69w3E7PcyDvYp1R+ew+NsdX4dNkf7jaDI
462oK1499otffsOhe7Zuo2csxIpkPpK0sbNGUskX96YAhapiYdFth4gSJPIvO2xo
ypmF/QOAR6ZlQ+QkxmN4J+7K2v5VNQWTe0Xvg1Ij2rOw+5JMKcggRJdJU2wTKZB8
HFpy7lYWC4YShf9oGKk8eSe4ZiDjXCq+kAEkMnahS0DHwTo0hZ2rj/FeeM8o7FIO
eWs7Y/aoyuSdv+erOu1vLZagUtObFWQ5I+7mCZjDb7g94hWkoQQM3UzocwRPBgew
R2u27mpJ1OFRi+jlWsT0jHzBKKHsEAZc2PDf1w/2bTF7IuPVP1yr62+OMkPi63nb
jn/xmLz6hEewXVysrkqo6IvAU013075qnZbgPZTPxvUstbyQuxYC8z60OOhXwTgg
ULQDmpwFb6kq+selwNDOeBd72qddYjp3Dp+YQnu2KQrc+p5d8veBab9BNNnSkWLK
vE/j+zzJA5dCPDj7LYETr9s45IIc4Ct0rpLWqWQ/5QDEI2hdAbmf0ncqoaSRkzOF
2YYbG4Yan06p3p0CAxGMzL4UqlpVz4KBo3SboJFyEioFi1qt3Qpa9HcalVgixvqB
k3N4okXGRuhrV78dz2EqYCiXq2SWUmwrTNXUzIWHld13i/wkjBzKTCQKRdh/WcUV
sgDtWiG0pSjFbMeZl3yLzYWiHC41AT/5fbj/cSfUEWJpRWxuZEq7O8GzypYUYzLR
/SPan2EwRS3AxxjGfZUSieMScBh0d3+RbBkorAEMWs+xs15X6/eS0TQYHaFBk2cA
HIVYXd+uVn0l8idjF8WM+P/QQ4Jz4pkn4/SlBtFhWnZUjVxGfOfjQEAITnTqJgOb
JhjbcGe3XGHdUoo+tCUD2oWS1D0MtQxq/VvldrX2d/SUpYGGHqsWgbYqhhKuSJuB
NfKEwn/dI9XoV0pD7hmz/KQLSYr7xjx4Z9TgeOO/gbwxWmDBmVsPQMBd3Tgp6uBO
gAGbbHNUCMsv+irNnaAP/Hnvc9Zzp+WXvYqO/Df5h6yZfI24ci26m3B6MV/v1aH6
nYKiiSoIMzKKvBt2saUTmb3zJ5kdcdwTzjWQ2QkQA+NkhtBtDvWm2SqU69O3Rmkr
VJSYlFC/Tcq+Z7ElNE+B1ZsJfZYH2GMHbHh7bpUVCoPxult+lrAE7VGmjKTDNKtY
kxyfy+XgLND86kNevdqk8/MpafM+0Gi0aNG/fZTPk3wEz12DNAR3outZRADLCDI8
28wjPepJgfpr6uQQGvsWPJQewwj39S715r4WPk7NuN/9s0ieMh2Gv3b+JeV3ivM3
thhyH4nLXFcBTlyil5cU8fUmMrwQ5byY859/p6pSonvGdxagnSWi18fDeRHO2pW/
s0yxXt2rq5julnSNZ/Zp6G+ib6tyYPCje5wuts7o7rx3UTMk/bMLTP5gB9TOISib
q1dwUaFz3In2UyvAaBMynaNTbI1pNImcR2TItaDrRX9kLut2JQo7haWGio2xFn58
b4GEqO4Ux/TdKTjer/Kg+0575T/GG22BCVqJaaegLt5VqWNKq9HjcedLLwvaF73T
oGcDSwjJDjeXg3EVk/vgwYcI0akYR0Qnw3IEuWVnSoz92+kRAGCCObOXTlUwACfJ
RrEStkRmd7upF5RbFTljwVeICxubY6+kgunrthqvzKFT2AEf+q6IpDHu3sSzw6ln
0nUr+8wxBwWpTVDFuJErsWjWeoegIbuLbSmay1D/tHrN7J7/N5gwfvFl8I36QCgt
JtTBqAZeLoZhV1g+UNzE13Plic4k4m3wHul/RvnPreJV9Gw6ZtiKkWp+jLUUuQKD
V38YJSrbCNPbHNSFPhBxaQXfuHG9IjYBA4NBbdJuPOuUSqFSTa/iVgih8q8KjLoP
8SKijV7DaXjuzpMi+tW6TERWGGznD6QhInuIK820c5cXLBvXx57Ue2zpwrRaZ5jV
oHAWbXyKoHwF1c9HG+/KQw5okGKnZMfKBcP+RA5Zi/xUPvpJiCse/RbW88R0R0Tp
NVjs6eliol8e3OIlAlpnv92MxZZvPCT3azTfv+/L012E0elmyFXVBN9abs9EMUKM
5TA57h08UbxZW94p56DHrjeMbWmqE21eEKzUIvrK/pzPARJ9Kqi9U8F8sXXQ9cAY
whuOXgwTZ2uO2sm4L4B6W6GNgOO6/s8KvbHNdr8E+mXrY7y+/m4QQBywysK8d9yu
nhQTV9nyYS+A3N+B0crob+KRyjO/5iskgZwqB91AnQ59vPSVMxocEshcL9EWx/t2
1kiCrcJfFGDtb6gU/ZciykVAFFErmJuCua+WvxmUWAXFE2D42EgNvmm/pJt8tSmA
JU3uogMU7z/IwItUGMqSNifM2MCqZeR+R7rJ7XAkKYiCJTl7CF5JcguIs0AAK+Bl
DEDgLhSoTu7mOhgLuGLPdktz+x0Sy5FKQwsiP0nGST27lWcO7fce1TwVG8MrXaVi
+/a2ZKGWKjpLMlzN5T7Y+d3NoSpwNCSZMeyoeqpLC3rdeva1nMJfYT1mxZVMk2DU
XfI+0ysIFUENMjHwWr4M/Mzgr89g2GedYEiIJ0X4kICuFZYyelX6NRfin3NzH90V
bulwCXkhNc88+/an4dfP9fNbHEw1CQGOWqVQRwJJPobDx4ydTdWr3iJN0GhIrtKV
CWx1dfmscOooJ4kJm1PqOH+AE44GCofSqgLWM754kTEBdYpy0btJGfTEBbzh/XPi
js0AfgbufriAgs57374p3pjlxG+8hi4GGWflishRm49NHjd0eei7bBi/ZfVMFZk9
bUE3RGYXnV1YkGx9SCjrP3Ha+bGDH9V4ImbfzvdglUTbRJtcdgjwKVXo5yToTcOd
Q5fAN2MK4JW9K+YfoPM3GsASXuSECjvcmk2NS3JlJFdtTZSX/2CR5iRpDjHWmd0d
PgZgC5gJKrWBl0GUfYw12ilxLuNAgIrSYFSNxREwcoGEVPdqozOeFsPHrKLZlYpE
JQdFZ2iBWLC0jROS5RDYGgRsBZEhHsTEKi0864rAQKkpg0a+i7U8PLSAenJqsdB6
x28ZiE29hmSBRX82/O/1cUngVPXNuUY1Kolb1WcJBzfuWc74Zd8RrHoTTMAlKHPg
rKZCM/KGQVv4F0oJnmLwksgNMDDEDDlu8AvN9TSdC9mfQCD3WEftKggd/IjuWeen
wA636Tg7eNs/a6LQwwGEQtp44e7Ol6SGwUds4D6wwcKC52MNighQrkdHZbX1YBZ3
3IzTByJFQs2/pE6cKyhfznJBACkLMD7GNz9Bzm/98nmIoiPSvBS79xipByiUcdre
FxPiECqN2FdJGm8OlH/76htN+n18wNx9QV32ugjR29P6+WXevkvXxoFDh5wxpmFT
I+lcMdOCNXiiNYvZkAvFu6M1Lg+lyeU0h9TRFjQCNEh/SRoVnO6bYMnXXkXhJPsp
ckwnEHyi7IAVVk9HxypiG+ONgkLuzmxZ68xkNr04xlUQVhLE61N0pn1Ia6kiR0sb
B1Pq6E+1XnU8hFjG5J9R2Lj1dJB6CH5pl3AvwLat/mwm9XegBn+nZoSlAKD6Jorc
7+sGfU629p+EEGXM29q8lliB1sTm7MLhTkLpQwdEVv2fE4VHn7j3766/hhdlTmd3
6GldmITQS+yE+ybQ1MSb8bCqX4ulQwnOL6EM4ED1ys9gLLKzIKd0b0oM1qFEwMTV
mwXFLpdxLdAqGVtqp1VlFs2nwHdlW5lldJ9m0sioQKR6FR56ZnGuE8t+15hZmJGy
RNaLQGqfz3RTaqQfPUHAPYj2oTqA57wy4ESZdFJg5bkLXLgPf/0QFRTH9lRrgINV
QneDZrR1OhsMDldv/4/WsN70bXul8ZPP3KqNQeWwl2sq4VwNLCpxVv1g0VIkAO0X
1uzv9Pogtxv3QliaufvIkV5V/O8dPArm06B6HO2XioVHHFYHCF7R9tHn+je7XfTd
20mILvIY6374Y+4pAlTm6HM78ogRt89iEJdYC5BkTK+AopAjv9+gD+X30aJwCM7t
ROzzYdPDpAd6VosEfBgxKqmSL/0V3md6a5m5BIkRNdvjETUP7faqsb4qPtFFNJUu
ekwy/E8+xvZ6rvPimTYYBoWfiVv3PGNWeeeZsn7zlj96qffmdDrttAm2KQqTqyYo
BO5e4Ptof/IQk4ywKZXwXjRwtMonGdSbDYMoRCk+EyXy2KgKBk83miu9EhTrAbFM
pL8At9HDSBNqxa3/KdLlYxYbNrW7VrLa3UNyDekKQYA14ANobIMebetactedNxfR
hlfJigu0iHVN93P430JyphpJsr0DSE9FTdVfuS6WrPNIsASQ5fCe82CoNe/sZpPD
WjnWGmxW0yNC6Eo97cwz8tZn/7cszBU8H2WyjBUNO2uyFJv/5v0d03Ym+CHKZauq
1hpgizUF0tFa1ITBzB2bxOSy1iaK4gbK3TpYI4cI/gyyFBqlctwCjCdFbLqJTIc5
gh1tN/GTufj6m3Rullx7QFvEqbR8okBeoD9nnGSw0FER2k6d26ILcoD1iNuDPBkg
zY5kUJUpfpiRoKlZWaUUf8Fk7qUljQcr8s+xNjz6fsLhEgoUcM+073DGLpiVnNiv
1GjE0tlMHr4z11ae5ELmvWKDWBzU5Ln6SxQQqVwo0LjNO3+hoy0b8PZ9gQT/BFXO
aGwCe1KUhym4jPAvv3R33fpGYuo1TK3YUgxlcWg3sx1+XtqVz0ZBrci0NHn38eV8
xQ6Zqi4xigPkuTbDY6sW4S6xpq0ULJxMnWa/k/Xv5ft1UFikyv+X2/lf61PeXcnT
zFv/uLnaXrb0KwVpiSMPFfORZej8wh7U9NaS+HDGObu+7BDEP0uAd85E3ALzfVg9
vv/XBZajBPCN2CP2FKO7BHYWhSbmWWzXHtTwGJ2bs2xNkemjuBxyGTe9TE9DM97b
eWbkSIsUrFI5ooyW3VKz0URsR0cc9Px6olVypqgXueDRdXOYMiuTMUXxeE/uUKe/
7eoCNoXDowGnhjnnqB2nNam5L+hO3KidvsVYf8mHkEPltYJOy7Z0PwBAaMQh2UC9
+L5Ekf9bfZxRcCUGXxuARf0fSRXxGj4bvFwF/vQUE0cqo9YFZTJv2j6uiFLG6VCD
z/X+4VTnptiVJSXoWf/MkZpz/90ml6oOrqRCtpK3WCJLvyg121XE2vKTAA9ewjgJ
o2li5AmW9qa8+xLNGqnZacrRnAlkuBrV8+i+Jb0VRnQfW1q0iJ1X1UKjA3q+fjcQ
KykJ6F7c7WZ+c6QE+lZLWU6YNVJwzSAkGVu94PIFzO1Lh8PnUC4TxBacVDR8rfMw
cOl7MeRgu2qdf1/2wMKcqGMmydr7hol2CEkgDbPt+3o8qSGXgRDytGbk0xy+DOMN
JEoTqErW+TEF54FY6oAG3NN16nFY/bYT/uzZvp8gfROqw6aP2sCbiNS9h+KGAMAv
9MlX2gRObh1xqQpdEu6hozImid83/Px2dFjozLBEXHwq9/gPrsZK1qN+SwP8B1hh
LrbXou2ELYp2C75zCQF2pYtT08xhrSbmX3wnZKbyvCt1EimkqAOuayEqDP0p+Bg4
Nf+0GbOYMMYJx7dapSWSut4Ngmajrn/ZgeTiWRrJPiIkEgzdxKHsbnKq4mba/umv
YHJxUVKjL853j/1FbZDqs61RNjrypKgrFO3N41lnsZ2Yl2MvX2U4uHxvpJ2pPnAK
CHWSPiNKi7dBGqHK8A/ulLHh/ezJNEUvuv7fk+zjWDrZNA+ExazJPG7BOfSdl+Vo
XOpt2IIZD2isbZqSkrkPcuo2ENsa2ZlBREuItga921G6gIkxLbmCcOROyz7Izpti
PkAe9va2wLSTum57Mnpj7w6ym6pqo5w5pykN56bJGczfZ7/cKgREqktXFsQt0mUA
BkuwRjXc8zMBXCM9qh46mo8dJcj6xV9GDXCNjKQaXlv/OiS9jiEUuCeme9bvd5L1
5G6LGjNCLl1cwQkxBwS9mxRMfsMBwub1hK3izWJcF8+/YpkgxeodVDV1SwdXv5Xv
EFstKChDmVrtB7DqOWVq5LsaDLIPvZKAxM6Cwdod5aD4FQm8GNWUhLtS5cQhW4Iy
u9xJmJ+aIv3XFJybgMpS6wrb6z+Q4mjbtjwNrnl/DfqWbgv9pQQWUQ5vKOA0uNv+
NGlwMAeTf0padRe8YOSHuLcYPgT33bxKPBOSG25jFcMmIiZtRxqXSLDOKXOt9OgJ
Qg9Co62d+0FzU72bHzWN8jY0ya7Fw24Bf+84bla06hGDhSiKAigrwBXx/WoCXOZO
D2cY7Q8/CubGsxzcuyrV8oUNqEwAWLE5IhNkPrxE9PMnCm5+yHUy9r5Feg5f7wUh
5pDQSLp2n7dX2xJrV7Jo7+1M8zC8FZlVFm6p4oouro8kQOn0F81t3q7Bi9gCkyJT
0pny4KfoAkM+IVMKp0GC5RoNHFLISZ5jy90VTMVQ6yn108QMDfVaTdHws6zucTgb
mBxqMH/BulGc1AS/Z5CIEM26XSyhQ6NDi0p73bzyXlgu6teuiAEr7HmaZUWPNBBc
gj4r8sQo/q+eM++4xsPyW0fGnx+QI3ser/8qRlii0X+DEdrUamvaKyF0HX2get/l
5ilcU+3q7fz8roYBoqaFOwQb+iOpCjDdnryNzEu+lILhsiznhKAIbgGUZS6mTJSJ
qpTD4+QNGN10D/fmGax8Sb3jQaUqCLpY4upo9B3iHK6YuDIuHZitTNpL9E90sChm
S2y0CtxZgUtM8tYRewdDfoAvhiCNrgv2UMu906MMh06ONpHT5VsoNhgamOfoFZrt
Kv4mZPhAJ7fBJoXflQ/3mgYif6cnGmW2nDZyOlLdLYKYdk0LBIH1/+Ai3U6F+a0C
9joPC8cZUx/v5nwQBxA6e5hpstLPTA/ZLOMOzTffuWWrhrjqw1w40KfqKEy5VvLe
PHihNgVj9XxMxTM1SSztaHtHLTPT3dOp2M9qLGEPWDBrTX3UrsEFlCVnsrloipjP
sNblXy7RkRDXoTmYYMhqGKMDCwE9C3Q2YSTbT9LTForn4npjKPeWfBjXm2KokhA1
fE0eqodJftdpdUFpG12rAql068KxVr4T7e7n9yXTtY8QS6fPkzASeO5JN52f2DHe
ptdzHqV1/KMkpFx3QLFBjqLHnpzxipbyFz2LMHwihQCqyEQtURLOor7D6LnVzywu
SZ3nz7unQJ5k3UVAORxTrqqFYj+aKkPo55qe0PYQixejEGMHb5dMdEwK+/FayZYV
SL7p12ORtxTclS1ZYnZc1mgps1/ALGitK73+lRETXVwy5s9clQWcJwLUt6uj7UJO
XHnWeNIIAWf4Go+Axd68vA6eVrf/LIRTkhcXWsBt0CMhPA1EgFwH4nGG9kMk0yr0
vCv2ua7yPJsMJmdehLUV6yIyebWe7nFagcOBR320Nez/uy9W6IDHSh2UdTqXJ4ky
gLCB8c5j7LXndA87V3A84GWMo8PDkKtqSiilDFbrKplX+mevUeAJsRgGq+TidN/Z
gWm68xI9NW10J/Z8dE9UjNwtCcDNQ1gV8haDKEQ2hCeuNHV1zTIyh/KYG5GwVXTi
a8d9hB9zSiahQWLNgvppZPIrHyFEIkL7GYWCjEMMrvdT2pK18wVrnVik23Np/aeU
VjKY6zpVBYnSkk6fiHPCmpPe+AeX+lV/wl0vxwsP/7m9Azd1etJteqPKomSejp+y
MOmLlmW3PE2ymNJZs/sStKrWO6H/RWtQMH8Gs5aOugi2luaXUk5+vGaNtdAxHWyg
O4e65gDR5fCyL28i3yGhqJLy6gkQN7TCeUzd7sL/ZaMAYo4y9+Ng55OUlIbKbmK5
gx/jtsrZo95kdmbvGZx0mU8aWjVosxxrK+MoBrGcuwG/2jgTwQ86Qg968F5GuJk7
XBMSMyVYRL51AIY3appXmgY8Uk1Gfkt97qo/eAg3fJLKQclOUOiRCLHioc8ht4Q9
Q9wphfQP/jYtsIX/1Ek52jsxTg4WUC6ImzSoCVuN7WhK4qU9JuHLw7a0pxZ/01M1
ldO59XKiMJ+RRMuuCGGSoOb8B3e//RWhZgueGg5+EXYB86n4Oww9RGJNZivgSE8I
seuM24XgTA24y4xYWqFIVibkbTrDhU7XPmpGuGKpOq2axUPMZyQu7g5mN3YN12Ck
1dLEF42+86VIMSCRhriT0ilbVUunX4GkBBQDtLLEFmvfjxkRGrN0Smv2ZVHppFf3
E+Ipt05/XeoZY3XAGSFYFlyH7c6xKoexgxwlT8kvSOEvNg88Z7K+2ggqqRBW6LFH
RjsimehrHF51VApLm3opPr0Ts5rJ0AMTv641K3oRk09JK3qxgFQ5+ua6bZFGFKl1
AS4Q1UNgWSfua/8wdgTG/Eext/Vz00Z8rztDSt9QYLP1NKyjPAXfmGngp71NQbXp
fJEDFoe37RgMh95pvp0oP9nWbf4cKYRyYKXGGPi3iUDSyp2OKtKWUiYI5NNKuH5O
ra+GfWW5yOy5w+DlB1XOc+ovpw/XQ0ItApYcJsW/gQL4iVLCTKfTC05nxZ8I0Xhq
4xqmNil++8D5stdtzibLRNgSYIhP5Gu8Cb3K8Vlh7l8qpOfuQnmunzLL+zGKFtI/
uOOVY246cQbAz1u9iWx4qmIKeYHJ3peF/bT8KVuD74P9cywhmdOEsjYY5IFyNqeh
yEUPcqfO88txZH5WJRcNV4+iPZQW+VvF0738N4KOh9xUdSuf2/91GJglChzkTcr+
c8Voely0yJAHnL21EbaNS57QE5FZrJs8Jc1LLwMpPeWr1mad1T0E8MGqDqyPnppk
n4yFWJZu77DUiF93/BXQP3/9aC6qKkSG8Eh4huY0qEYi2KXxdItnjuOwMhoK6Qox
U13bwz+6RPlJpIFaB9rZbUPIcQ2zgBlVsoBvtJvTvHJYMIiHflbYvNf+Zw9bfN1K
E3a36/g796icXmQSGbUwLSxuZdNruSbcPY3QFFQsDRMuSVZF2e2YkOjFtp3YYfUX
x1GbpASkisRp+dlF8w3pkpzX8dZJ+v4KyO0xCWjwiQ6MNZoUTLEaGMHCHqP/7fd2
qSV911HCIfbFu+tQQZdTLDmL+CgrAES7Lmm5k9X3c7ipPrBl1J4+wX3LjveleKKb
Atqb500Tszj24ihc8fwhFR07on0pN912751xN857rIXRpnfpMRwg6EwvwO0VXFwU
vxWCZrNoyilFxnpKrTuKAX8V7uKxo+krwhkTZKuRgvFgwMIeWp1w88gm+eOOSTG0
Pg5E4e8YU9FxJIBHVEax0FvDwUcH3sF8XzIn31zrc4TrBps5fkr0Ik0mScYMn++v
ZSAbEgudZuLCGd28GIkAc4asev6sTbaJ7yOQGxykrh/EXHdW9HVov1yMBBXHsCCJ
QwlgIWlQ+p+1rVbla2bYoXQKZWtKyscGCWbvSUpW09Wl6Wz/mg+wmcfguIn1N/ZU
5ATLMsD7Yj95pnNkJhH+jGzcszJgkwQ0r5TgFvwstJmlugXM/gRuSND1JSoeToGF
Vci1N6YNbZG02E1t2L66fyvLFLVapSf93eHAPXesbx1BRYty00XeNX9NgxKKn7C7
Q+n0t4l2m7mBXary6mI0bT6q6kZ6goMy93OhGIzO9nUcz6paU+97v8Aj06Cs6oGr
OGNj0OIqiE1znyW2suSicug69D7b9Xk3axWS42fhyo37NuNdlOe+PQRYegSTnWfx
TgCm/viMZsQfUFoNcvI6JTssD7lk1oGirjXU2eTXffI2ONQbvuyCpLqsfHNXF7pN
Ux8J2Sol9xlT54TmLdjOqTTBvYaPYLdXcQeokd680l836JHoO9vutHdZTPkyJowp
5cIo7iqjnf45cVFEpO0Yy2HehfyktkY8uuYtE4K28Ag/H6WWp63nwIM+wXeYlZHC
UzxEZeueLmtg2k/dcuKSz1awzzk29cKNaXib5nu5KGgV94kJCpbWLE3/TM+vrK36
gO73CapEyde0KjWX3nnodb6mjXNWhemE0e8r7PWuP3i58bcoOLrdAmpPeUzl81Y1
uJAednzqXhTOf31QtlxAQyOoE5YsiIEWHVGPAlnbq64zwBw/IpsdYaA1PvfVd/dT
yMAsRFQaKwpFDbT3fgfHSWqNY8ffjFRWUapekoKR4zicfRHlvpslR3NPSov7smWW
lB+ixYJFHba1ADtOSHpgyPdO0VjLNtQ5paCBa4ntyl2ZIYvgsuxtT+WEepo2oCKl
wAErNui+AgaIreHkq9igop1avs105z65m+Y7h47dtR4XNJTBZIrHCRpWTytHMvTb
WcvNt2/wNk/Vxdeehcw62k2tyrcMIkFOgN0ZGu9YgEsI73yWKf5ABMO4h1Y3Kfcy
MqBmDmkDh6RQWB2cXU5qSW/mQg6f6A5kRnNKuUTRQtW4usQHtLzufYW8RCjdys9u
InmqS+qO5eaTPlqLykuwb2n405/LkARrydVYBr0CGjDAWSES7qprtKYZdZf7pF2y
muuitrGu2Jbr4DNxmOvPlv1cjof1M+4cH4Z7EqkT+/dN9BLbRKpc3PTR7PiTozca
cMATk+WVAaxv17HGZL5EsFJ1olhLjVnInYzp0VK88Pjfiztpuy/MXTR+yLplPidC
A41J9+UOKeEwgb7trFf2JVS4ArBAtZ4bLR8hP4zgshltDokA9qVSTx20WbxCaxc1
ymvlICwT0hW/Zg+Ro23kiiAZsVeT+/yP1x2yg65FnPwgpDI+lCSudu6CCPNww8zz
JBnmdzJusE4LsDRUltYM2zARK8mT6JfqfTWIzU0k48IgdFAfb6Eg3pRuOKWtf1c5
f9bp+QQ+mVDJkgj53D6//AbKOYup9uXvWUZiwHqLSJfZGn7rMk3yDlrjLNWn0uhB
oQ3UlRyiyfLLDCF7tQGR7MtnNV5UbXwTRtOmvxaUsnv134PetztSfbIv8lJBIaHE
acGK3ujlE6wr0nEqoLWH0e6mE9sQylmQbCL71vvJfP9OHUvK/72MEZzCjhKJObL/
bQnHvPyoYRjDzIG9tMf/PeDfs81+npaIomqiciM1P/cVPu2QBT5FGCU1sPcGL1in
L/2b9bYCeoLaTYWTC/EIeI612zChzKkricCbPzlenTOooN2Ato037bUBNfziXftL
CqoJ6GR8WOVRq1NOvmWqKGjVCADDQxuTGcy/luQ+0i2Evfs62NI79eFYu3OFCHYX
Vb/s5PMKxPRaudnmusySruR7eatoTwFGJhmy1+ySnpYuMR+N6IjUIwG/wofPykDd
NGYo6tvDBsq7dVvWldM6VDb/rHHySiygk/EYwpvXcUx+3JSH5B45zRzFP9OYtC0D
EzND8NOfZdobaOrIbmq3WwIBkTAlDaLmOxu750s4jcbqoLa/M3lpHuUjeDXEbp3K
JmhaKQWmf0z+AsyR3IN14ILlF1OuRpTN/XzgnUtwTIwf3/unctYR5CqXEzGcwNUl
2c0WMLCon32ZMMjNLNphguH2OiybT5UBSDjn4/gKIPENL5+4YON5G9gWHKknsgTo
kCqhpsuxI5+RpgQRUFKzXnNl4AUu7KioRR+84XyT5/QzoLmjR3VOrE4WtgzhmvWk
nhJkFBER0T+Ii4pLqDy0IJtQOW9TI2mqZ9jsuVvBexrjfVRNf/jfyn2LFnaVHYbN
laqBtlQA29vEceROLpE8r+Pk3qlFdH3PbDXP/9t8Kejpw2lYkfWUxEsrxR5eUcm9
54fL1qRMkMdn8p/GqsAKT8kTRF0mG15n9UEyk1whDtQO57vXXM7JSwumIkFE2/I/
GIz3ckBfj4r8hfVWqXCqg216X5YnyB8sGRvX09StwAKkVFvvVCF3qaOabQV8ixNY
UW5sycNWoud199xWC5WKv/1tcb5xs8Dd7tRKv7Xdf2vRJm4lji5dDzSzy5hub1XE
gNVB23bxsoe8mIsJGif4hojU/z+pDIlSQIxeFduiFmSfSjY5f2SeOK/Wdt0COPz7
URsrAlHV/idJPdfIjeaMPLCpnjRqb3j+cj13pj6quDUGyqcTx/PDrBZ/IY2VS72c
sI9spFraf6eEs2EVoBS1Kykxy7j8P4LbbfCaM2JPXVxbEBm9ewgh5AcGEwjo7LcU
MNG5rKTa50qBijzwPjG7EGRSVxFmIB0MqWgDHOHgq1EsfIajR7JGGVeLSLam6MrN
s3YmcL0dbGdRb+CW7fA484DJXKLTgxPGMBAm4rRfX8Prf1fMh9t8y+JF6wwF4nFD
dCe2gpMnB+VVzW6lF0bZYpN3FZVuHneE5Yur83pJ4fNsk8mMUW0ilW8TYVHZ8H8H
ZK+F7FfDbw2hYaMYUp0VPe7vBW8/fseCrvrs82adVHpOM9Vgwvq+yhUQx/bBwmE1
8/XsxA/dXQLzZeflDDkMgyHpXPIQ2D4WikXzS276UVdw/QkIz381mOEW6r/8dXyr
1W/R3tng/xFSLPTcZwE/wqH4RLzCB9QVMVg/X7txsqwW25XJvtlAdaabBMyKlJJg
p3weA2S4CI0PhA4ngs12XueMpL0CzxolX9jfe5gclAXCNNY7Wu1jKmNuYnE2CRiu
meICDJaWr2flFvCf5iOCcKjEPLebe1R1xgYJvGZGo37kIw/XkpQ58NS0Moigfa6t
4d0zrvxkvEY3HcKCjfDz7qmAxxpAVYq60wXEN2ky6aaGBR5AjdUbPOjwfHesoD1i
5EIjYysq1kvEs393TAczxIVXE61jTYSCRjyCyu546KtVVJegj620IAsm1AgEGGWE
lsIVL70C8W22yXRGr9HemfpSGCbFh8V5u0tN/BKRXbQK/NpMJeMa21zV+uixGiMc
JPaM98JXv+vhB50L8G5H5XcL0hyWM5gfsHVrO0EV62lNj7O3xD9ZIrCzTj1CbsKv
NG2tY3SxiJ09x3v2vv3/I985M3hRu12t9ybEXD/cC9dL9xzdbDWmvTNi8jPMJY11
YeFpbMS4QzsZ/7IdENwMful3+6pG34kNRNtUXT3lZ8iOdeKo8FamS5bBUSQaj3uk
UAnc9td8AOKGL6jK5YgGTiF5NFaokKRFV5XcMPVt+ujXLTRfqN39WPFWS7xoXuG7
whmVAjGf1Hve87oKIN0/p0oJpPD6DgtPtIfgLT4OQEzd6++9MaeTAO6I1q2Ur8wQ
+i3E4kwhRG9QnkLYTmkQnJJKGAycVmwrIIzPVbH8bF6tpxTs72vIxCQmbRJfO4E1
LW7oOQ+uqKcKsoKyo2oI3jKRkyJclVtT0k+A/jEja8WvO3Dkenz+rPmKAE1a/7Kz
TicJ7TrtTFXgGpTvl9bRk7by1Sif26p9qbtNjJxECxQ6U1XSc6TZnuISljJyDBdT
NmywRtcrV1ZhLWCT1AIMCrI6PFhb7DeAjtWBWB99POAQzmfSD8XEPLSsu9/BDnOo
JzHop10CqlwaxKJ/QeG1dJZFdFxJicVCcLVtYIDTSlYjEGWbfRlxGNn++bik0TOZ
Jc9xcAogxuxXYPaLuB2xOXqH0kmqBNFLJAVkONubApfisdZNorLuoo7k3YItadWA
hqITBKvzdyNsVThw6ffEMy/p5TpMR64+QanVgeQWK1jlX3NRBfn3GGUchRhl6tHK
ZivJIL0UeHFxAGv//YazgGUwnqBMMfGMU+khH9RdGi6UEd/cSBM0J7vdFLVqeqHU
Y3d0pCA63jfgLZqjC4tKSxcThmXv4V/wLTOq3qtAKoTx3wWkqc8XpP2QlHwpl/mX
o6YRDbOQd9EofeHZliz1FlcCLGwPQENx6Lui2bUX23rZy+ZX5u2FIvV8mhxwgXPW
kQZyUf2rU8ix1CEKymh51prquorUu69PP4xQQK6wrx16HvYxvqt9v4peio8tPdc/
DF3F/veJQ6i2yeRYdyJeHOAZx5fI/K6AgEG4hZ6jKZMJJEcNP2EyWtZ2/tHlI4rZ
m4Iy18Lj96y64SEtuVmWeJfS54DkwhQyMEmf5jTb/6mzUZUJlSW+lv8tgeHxld5I
fmvMCIDZ8c00oYzFfZ3uBpVgC8zSO4nfy9BWIdLANRdLw9x7VNFI7flUNGOCYmuK
Jx3Hh+WxdTYHGLkusI7p7JLfFKYXVByJfllm58KIvwcgZg+pMFUYsWnahqwzmQNt
9zu9sxSBJuXv8911ALcxAdSGepNw++5JdRqV+0vlDyMAoaGycMbPZJP8EXXGRwvM
DVx4ThzOPiBe6KDchknxOhCzN5T/sSG07frgTenZ4oSPZt1l7y0yLAnc3J9Whp2+
tqIbKZQSnL0fSO+fN5pCgII9hCWCv4rzO4JE6idKOUQtjHaMKO4Y4EL8JVcVImBc
q8Y3fYXVnhhZSF9fWBg+Kb726PMLnJ+m5uZs48Joa0qtUfLFc7CwmL1fHEzwOx3O
GXqlFt+AS3o1vJjKforKHZP8Hi00GtnBDSibez0GvpGOYSHPZqKwVKnx4TOJ/GFs
wFGKRWUZY+jD1zf6NqqgUHZ7SIOkiJJydLPalldjM/SOfLJUNftPvOnsZ1AYSAE1
8AgiX9BYCLZOv4eaN0kyhNM6TGzkbfsuMWIzVsFzy2TxKNaZJppvfj0gPp9aCxSk
8Z7+kvg8V5rYFWlHhZYOB7KbG/jy2qfQsn7h/OJFVbUu3OvneeYcCJ7MIPVBW96q
4bndfSDmgT4lmOwBM/sjzpzxfTiP5B8x2ucopWVb6WfoJlJfSylTG6P/X8msV6Ne
IpTYaSLmrv5yJmIkHfEWV2TivAbzs4rZRbSEYde82ajcOR2O2wUFWRYpEslCqr3b
AO6/RfoogyQrfb8xRW/JVtiek2GPMbifEgcO/Ds7lUOjypqM4YOPD1YEcOgdNhAi
X7Y0i/rWSW8eKocG7VCA00O5W3XJsm+S35EjFf+q3BcNDv7sbiicioCjVUZSSRh5
0rqYBOLgajUIYurhQX+VpUNgM4qBwab9QSE3HNJLCLZfJ09ulrKbog5gP9Dcl/IR
v4b1rYE2so4M/a8mVc+B3+BniIQnzrE/zGRNwbjXdzorZZIS8E5cpCShg37F6W0j
pYFarkmwBeZNXVwBR+8cA6JvlNbdIhbEog2REt0pFFbSDTQKGm9TnCVR6/aayJhk
t+LOvQYtU1SPXMyj11+T0zPzQUw5MwXl+oFfQwX65k9JF31bNeDlxh8da10pbi6M
TtIlA0X0FP5cFZleOf2MQq1VCdRvZ5zfw1iWUuESsJbXGc2yzUEDhcth3Wr+Vw4b
x43FrJ9LbDSBIl5eN+GAomIrrgTSqz/vXbvblhsWg8VchEG94u7a5TRx5su47H7O
gi8hcictC0Dwf985tkOxDIt/0wL9PD3MzzMtsjnQ0uSSOj4HYpJQFXVakpTAbI1I
lP07ELKGIvTe6RjX5nKT8yLbtV72RayTRx+9rzNqYzhRKE3lOAqIZPmRDW6lZSZt
M3DUq4/PUhSvStq7v6u/uGRPiIOfPv2FAemarGOUGCAGDoqJDkqqi64GhM72/AJw
f0bBBoDfxFLyC2wWy85V4WuuJqytsSCvoJYh+/+IRF9Vr5Fv7z/TXIAnHvaqO0Qp
D7C0iMJEL8v4d5KhnfuO6voMGjp+KGR/GpzYq86wM2YCDGEfir8Vn7njPBqlfS92
4TGimrb8TucHN2DjPlX1hQnhepEGrDv7uXiZrF6O1dLkEQ1UMbEySJacsGgJsYUM
VSMZZknBXk2/ucU4O+2PGFixvJw6TYONQQwVwN8tOUfW01eheSRA9B2KjnGoPtRL
+n9xnZ9ehibmyXkWUOWAtHhfFuwOzrt21T15N9pXwBfY31oBrBDPgM3cVeFm/Vpg
bbI2RZoLYK09sMJCjBYSm8ksiuZsoOKNKTfweXGtuaEnzmImmeea1p4Rv9nFvIzG
fQQiTd/BHJqPc483fGQxZrcpCN6f3r9/CiS82RiwIyc2h9dqAwj8A49W7abGTdoC
GQyVIdhSxRrkNbH8pFDFjU+Rev2ZbEMT9wDxcnOeaclguvPkkG7GnANpma8IbRka
prEOScB/T7qlnafM3Mcj7B9g92Ni9/M1DT31IIUY7JRNctjoyDU+7fAZWZ4vhtfN
nqrqfilqB+EE5mN3XAY8gFnKgnzZmDcY8XFvIgku+7nK08m10dHACJGPILXPyRq2
HwkRJMmE6TOdWHXjhpen9iWhzBej5do69FUGjqg8fw8WxHcy2wgm3XpZwoHKA1JO
qAqKKtwJHfjNQ6YXwcldBMGCUtwfe7fKXxLvUm73jTCbCZFBU0AY8T/ozKTzteBn
DayHSfqaR0mSB0MO5scX1l1w5mQ1NVxjLg6+Oz1YqsJ9M98ClIgTjfN2/hP88NA3
ZY436uRt+bEmC10HVM6EgXdFecUBRSDMtCoFPbPt1zM4lFMtMg21QGN1iJqsVBNi
dLDDNijB+WDoZKoAvxxCIFe0GWrseJzMf638VR57pIsNIkVD4gJlhuqCkJgu3Jix
bGYwTCI0BYc1wyjUU9eXYWbFO3fID2mo+cAV88zeHctzVw4tS5uNg+SvjE+Y6R3A
dH1pGGj6VXQDtCqUhORY4406SF5puFUtS9hGqtCvUtqKrlR/aIMqXTmuBzTqZK1y
jko5/vR2VKeHhgAchk77VotdmuCEzaVYNyFbE92h32UcaORJzU4dsr3RFUW/1dAw
5A7011k+upimBfozMJV4Qhu8OKGW5JDZf+BRhX0B49gJdmmyE0LWuoW2zobZvgnW
FbVeRgG3tRJsHhQNuuXmRuKTArx12kq2M/MyJaOGVGt/G2uFeiCIUE3Xd5hDb7Is
SycA2PuHCGMUeiNTf9ZKDX2j07lhfrS1/aJJj04TZO0lt6DElpl7sy6p34JCCuO0
ETV1i6GjUf5sUbToCv3mgVFCfGGQkxpMBoJEH7n0vGxLJOllbcivG2qV4yXirMYs
ZMBpUHbEaXnOAEaGxEXSFd7tJzBbzkRRlOr40YFtUD1G5TdYYTWSdGTIBUtGBpT8
iELaJOCJ+NZL8Fa3X8c63leAPges4ivCPDJzoc8FzHl7wW9AfI3fMIAeSVw3Z5GT
gDrAr3BZN2cGVQxf87CQYplzYch6FYXwuplEeW+pSUFajBNaj9FMU3NK7DHn/e87
PdRdw0MjiwLN8imG7pKBJcRFvti5p3r2zrR19iYNHKPgxLjPzKGmeRavIlR3ypAF
Csfr2znzsPJLP5zdWWQC9Xj+cTvJMZMifQJhIelWi8scvr7soH9BrHgyEouuXyIm
UNGUK8lr4oGAP+iafSmSNJy436Q65mzFzvN/rppJ5D3RXVsAOMj/ybAdBxy7a1eH
W79j2MiGeO/WApCVLWkzPA0LI8TPHWfT6Cc8JrQOeUbxwdbQ3cx2yx7hHCtyWEOv
qDCMVkh6UzDL1cMNdCvDwjtdh08qvULDJR7Sj1GYDDASqj1QZgZ/we1Wp99ozVko
axxieY+kdPR/nwcWSVFP+GXz6HMHPDAh3j2rAHCEMBAVq2ozhFeNEEUfRKowShC6
bLNHdQMSAFIkI6gWnS/UWJbJ8mtg6Tn3hhcXfzfUltC1qYjhTmsZ8KlF7Nw6iC1N
0nFnKtEKMznw54kiWiIbtj7+pmEysA5/ePYiT/0klVXxyfOiOU7KX1F3LTdkFLu0
hRowDhlkEFd9ckXx0XWVtpD4sVhx/dBmdhWd5uFZwifY+/ODcekqy3QNGIUG2wr0
aCwCRSfBvYs69u/O8S3CAvr1V6Q36ODQ5V7+/Tbsgg2NNhf6v1WcBs3DGDN7FT3a
+ZwVk4EXqdQx+aplEjd/yb0x5cU3IM/n3E92iAej4aOqHC5Jo3UZMzR141pHnhAX
rU6lp6FTmth8lQLyDeikpG8RK+9zME8G8IuFos49nE5COFaej3X44Lw5ugnNT60S
i3iYEoIoyCSUT2NH9GxR1nRVZISNf8vNGfs2/2L/HQ7uHnLwjxhov3vBCDyKXDJw
AQsGme09zlRS6KeAoCz59D0SBBNoc541qrKqv3hwn5FAfIHoKsfEXCFggMLmbplF
HcpTijtePW140FoCIIvUAo3+LeoDKcz08keJAW3cD/mwaEA9B3vE28RNNQJVxN07
8iM7bRNSB6kLC1422hjvsYNvfqjW9eBumRqZbrZhwHb1EQMY0b75217KmTZtzi6j
kCclFKO9PUD0xLQPgcwDKpqtn9GldxxSI4K86dyJtY4ccryXQDibtNiv5RhGEPs+
FCl+NHcEVyXSFTbNgLjmtPAVolXHqesKZP/neeS9Yz/8C+zMhFt+9U4/dw1Ej1gD
+RU8YSZZGAYINKGzkw8DlgzkSAWN9vqDoelOqD7/JQLInXXwlz6DqZj5nXtIB0wm
YR9U+3hbPIrie4qPVCksgkq75b4Nis13JTgHgZwBHvW4N/0QaEL7hkffrBad4yJW
bN9jBthpPrVsThhbgE+9PIRkPLXgjD5yEaa9jCVQB6UKf9z07aRJBsGIeEUGjx5J
NMKJnlgH7e/mN3YtfDS8coEaB0dQ1NgkIgksa+M3L5u+6by1+QkmdKYNabbhMIsM
r7l6oj+dWZEEQIYN+4yl69EZ24+fqjr0yKKDgfiUffBYCx3gotseoGlaHaLeFT3u
orLAAN66SEyDbMSldVSvHR0zMc4hl8O3E7ODJnFslBfzxZCkurZBTNk3XxsSd5kq
ebBRuyLaeCjJHf6ATzP8RdLorbVwfZ1Y5i85qNL6qXjnt+74A8rjGFAV5EzErRCS
w1BsW4MViTqmUY/mg9zJZvtj5EvZKz0eJ6wmh/X5ey1D3fypr3KuzJtKso8Uz+Yu
SVcab9EBb/yLyV1iMJypq2MtL8jVVneSW0DT0mgD/phG9mJVqi+OlevihG6JgR0E
lCVbawUy8I3DAWDVyz6P1bX3AtC8KJvh1Tt4WA07QP4He+nOHu9B5RF2K734dfmv
uS1aXrKefnDCuI0NYM5sRXtccbf+GvZqlrlvH4OS3mpqBo5ASAiJbGLYDzRlHbJe
rXPnFLzbzYHaHpyi4jEBq8fQcWMD0hvBLi+VfVECGG20IGUDoIfNMkBRUohvoUUp
YIVXcervXS7mclogQ1DGuwuPORmWfEd9YLV+OFovv8JhzdsFIHEJFQsKF5D2sERy
eip1x76/lkyVUTNfYTNfr6vwOSf/1F1e4Wq9XHanOf9RLFB6EUoHrABwscEZF4hz
p6l++voAX4dfykWw7a77+WPYRSHeIhoRv5wH4gtmxQDSFh0PjOrx0KzAA9tcHYee
vDdvq3XA0rH3IrCbxVnU/WU8J37dtOzStWIOM4BGADJjxWu1GljDxIp1rII00iNM
J+FkOMYqG501EsgVAybq2n5KC9gsJxdbDaIHBYwnr8L13YR9vBM6ntJyoZCnMzMt
5FN+SAiw5B3Qvxo5Ne7LtQl9pCJ0ne9EpVRRb8KZkf65+TbeC8WoW3rX6/1nldR3
WNS3DRS1y5hcWF5G2XPhXbiqdnYUdnpwWlKQfq52U6Xf72NyZSGcR9A53XyP8J/H
k0z8m8fWvtKwKvU7k0IxVG1wjDXaNdwNbRo4oa9c2fUJv7mzpoWibaAA0T7MUAE3
uQWIamCaEYvWcTv5VcnARXhCyGePEtv4pQZtQWpar8ISa3yW4COFkU6T+vM4uXvx
h5boOZq+F7Kw/P4EhGxHvx7aGZmHBXhAeD/MhoSQAd6+FgmzEymt25cg1tliLsjL
SLX+XL6tgX2AwXrcjEWH0hb/DATxT8aXlUGyUXrabWCWqm1bXFPdxTEDe0RSDX93
hmIMqSBHS1UmMKB+/l4RUYa+NmuhOglPBYzYxq6xPyVNkoiAaoCXCZ5CBAQCrpu5
hU9O7DLEsShaaKrtAlQ5eJRS8T0elOMKUVyt4AOa4ZLZXqzVXmCg0W/ztQgfLy6L
rIUUbzk8HbDFqAsKZxc9nftECF4yAJhZu15izXGJTJdkh4F+tfVBu0LTv/sCDDpi
VBrAxO0i47s0hgiywkPwIb5p2O4xEBk1BDCx2IEqkouMRxmsaaS/SW4iUejtFoOO
LgOme5if61DtkOV2a3jq5b0DAgckXdas6vAy1VsN/7HJrUnRnjaClCbUtXCG8WF1
/EfLGqgFYm6BG22xGtMvRVv9e7rnp43lct2tzryWu3cV6jwWcc1mzhHrn2zRluL1
jIqGJ442MBwy4ByTCwD2jSUys00eamHk5aiMdbQSKMUM56uA08kFsZRfIEdb4L+J
I3klso6ZB+y/YU2IdBiEvxlq8BzLtLHS1JkYyDl6R0V+nI7n8IfuqXhNJrYnIyJv
Dlr3BNiLumE/3B0IrBuTTww0xi6BoY8llWPyCMGlVvHn5Js0VwFAP3QDVOMT3NOc
KmIY6MU2xV0X8zR0OCvkS9G8FmmJEgq9GlBrVm74jOymIr6wEfdyXE2oVkSvkaVY
av9sNIcslDwf6KcUDESgdZt5Z9R5Uh4V7VovIES3szSUpYFqySygFIm/a8PP0GF7
TvRWwAQlTQDd0Q5N+mgoY0VdO8AHgWYcUVjmjqksp4fXu/OfuJ62wXwNktDFMkea
EXE6fSHwOcdYqwYRuTUxB/PlX7OvmfC7kB6fiSdEPzjes5hIXo7bBYSL6amI5VOm
dEpp2dfC3xDiFHDVzdJJt0HaVIOV5qER8JEGXLC5Oq30cB5FcUHWiesk+y6gUF/Q
yKMZZDGRFjWzjxEQv0culscQ+LhX/7UpIXPmOiN8nH6bI02wXCpMgGSjQv5c6xYX
BqPLKd0PYdjlv0FZDuu62yRZ8ygAaaU2yMNSKD0XUX0xm7p+VByyXolyNco09fTA
F+yDXW4WDRrLhSMClavJRnPNPMbJv8esPHAQ6e5PqULZOKHaU632NhoIeWY794dF
IU9aB/zpyROUVxRILZ47+bA84ArvJBq1Ix0EHn1E8LFgdrW1t72QtPvq0xz5r4/p
oPkIn5YjlVoMKDCwi1XQXEpf9jJzqUIGR003+ztlKtVp3Md0rTUy24m7mkvK09Gc
5nFhxrjhHT52EuNtFaGAOzBxeisK7zpB9I+6fPkiyrv27yFzDfXsHQCHIZSz0SUA
n2yUr3KJIBOHasOvSNynHD9uY/ZzEw5hVkpZgIq2MrOsYKrGND8FdidEj90K0PRf
T+R+eMkEObjIrWKKmX8WPGp89KET4OajLYRajZ0jx8vQvOlFbdbLjCKXTIA1MP7p
RtaxbfeQpLKDDz6SwV6k/C82xlULq3Lyh/OiUd7pwkcGWPEyFd1PWePzAKniwKPQ
rJTgqCNqkP5x8EhEwLSrpZX0Bmn3EZ//1edjdDZJsGzD0eGVWDybq6+6DnmCo66P
kQhwMmm/MXkIJW9pj4bR5TzQWbZEaXRdCVuFX6TKcZArbrwCKZZjEtzkoeJyNMn5
BjuQiHSJkLTLuCv9X6EC8C1vNQUBDZcAho5QOgjrDJaYJe7VHrtnJT8Ppcqf6NI8
arVnUmln82bKSB7dCqrIoefbfZXKzfIALyK0b9eG9jkoz8LKraYpC7M814z39RyD
QsQ2VmI1AkzP8npyKZ5y2nGtRsNAcNq/QH2t64gSSzGKgn0PHMxM+ekJ0fPDYdBv
3wElJ9Fa30PDZznv+D2TeeOQg/tXc83lJZwApRbosAHcZu87XcJS4nY7yWlkONx5
5Pd+lDNJYSPu15stgVKf3ZTc1WWp01un2DzxpmFZEho+aPZWZ7DO0qlfceHk8LV/
ASh9e2uoDzsET4FPxIzo3U0Jav7qn4TBwSV595JxlnQUjj3KK+npjfehaASj1ixN
VQXaSIth0tMpqwSu4b7xCN+84ZJn+e8xSCQ+mel98Ow8aoJ6jhsONJ7Migz4YHJA
EQNYIBBwV5k/BKISxSIqIG3LuvIWjO7l7Ux1/I48a/M8/Pj/dZ8YX0+uMW5n1NeY
dCliC9zNGJ2Gf8x+gjFX6TkhS+UsGT3TGH/f0lULb+/GHOx3glH2rHv6EI6Tem2p
T6roDvc0Q5XxOH6eTwtcZSrxmG6THUeV1DGSWd6yuHz2aKnv0kPaZ0Y+1Oeq9pEz
2imQMIdjsEJojiIO4/Qoejki6uMa3ca55fvMYVM1MY8pa7hfsz3R4nYCgdkC8uqB
StaDmixH+mtMciOrqrk72pEvDhnZFHLGbP+5MTYjEkM1Vg0QBPki8eaCILAxG4Hn
IVqU3z1o5IpvgM7Pmpd86rKO/AsLaK1iyagYohWPP1FGce3KNqX8u0tV8YbeeCLX
CXW7Mw7YBqD+0h6ZDz8yAdzhNq2iJMt7Z+0wxo9FzhyfjhcZewWeehmH8CwGHokm
a9ECBnmsM8eqixLTfxoGMEQPL1afriAe35uNrNu6OYv8qmNLLxD8Csy3AFORI/DU
h6nzDsysW5Co1GxgUQshaxUFnqTgOfRpV+uPtWDECNczrepzLK8cGiTRMw8wSe9m
QHzk75kRnclPeR2ZAGa72Uia/p7+p4f4Zx5bqfbMKaEC5zjAUAUDGDT6XVxZwMq8
RTLXGqcST9wLkv1Y9BOVw4B9DVT2IeDsSjrsfR+ti+jRBUta1W0kpyRZImCfTxXh
f8PR0akQc6bakm2sHK9ZtcRfs1ih7q7SmFYcLAfIZmOmXWCjNOH4DW3oZ5mHFrIg
Q1MCk95nfP5biM9Sra2o33zF+ELShMi3C7U+BHqPYh92mysHsIxHtUuS0vsPNPic
/2zHT3evHn9Sf1Uzcv5TTd6pEASurtFuO1u6ciQDJhMBE/DdgvN2wKXHoWLhBtKI
mAxaqJ0wCH+3CkExLicPA++eUhVwVP2aw3mCIURl8rQeocPaEZxadziyRMU3u+fN
yk6uO+hv7mAU3dAzAL8DTquLCr3NyqWxloiCCPrfjOpUbPAZsc61A/wF/a9TzkcK
tGha1nmOU3zfmgFl97xFN/xSgDm/YtFE7P3ByIpzOO/97SqH4nhOXTEnCxrCdn0Q
KFaXne0LYvUsyQp404QVN002p+5HUY/NMbIoCJPoXwMBmZPklqxXPnnIih0r4F7k
04bPZ/EBSIrwnp2rtjizyuHfaGj615luUN4Z19IjDEOy8BFAzvziFvfq/X3F5ZR8
Cc7chzKBwOID3tj9VGvlcJiYn9ghgkF4McTrWuOB2sO9SRgGAnK6idjJhz4BsGKV
lavgaKxUPHwsPCD9nt6LNz6nOYR+6Sv2xINGRnfIue6TUoETUGwoKIvvn0MGshWZ
r0fRVOMts2Jev0SPjFV0M9IsSjcPfoFjt9HJSvtQqPL+JOhE836m/BfS2WpuIZUu
wQs5k0EqPEr7qIxxMhSEbzCG5SfIkgO1iuzXm9KqQ7yZEyVHSOqNqBn8ZE2he8V2
G5UIDvdrziCJvPEwk1tjjnGo/RqnvK9Q+vZrVCpSXyx+yRGehJh4tFpiS/eQzjOs
Bqk1NjnzqDVtkPLHIQreYnbJ1WcZQjBLCKG+VmCfDfejnTroBZJbw9exmzH1dau1
nqHoxabjkYljVHUjghnJ6IyGIsFOx1y5aBgoElEhDjdlTmaCEAT+J8DJd3BO3joC
s5liC5PiWWxAtBU2InV4p9bJJjsOgwLOCO30ZpuFaAIRvoR0orVe2d29dr0pyTsG
XFZzPbXmmJWBnorMxU01Y1tTdZNuQ4ES092PtSWlchBBX/X8j0GUs/sNzEEdRPMB
fCKAFaHW93+95KdquMMueO9BtSBIdb2QwOnxFL20JSiUkC24lz9olj7HFEN4nXR9
/tGhkcEjWhLuOuBBBCMHTx56ZsPeGxk2uJH5LHXqzG1d3QlFBA6LMObsEiMnhMTC
7Xu6enNo90a/CyFBqYBxkzthZTFT0x+Cld5EZrGRUzd1Qg3DQl1gQt46B9KiTSsL
1tdSjz6sWsndTPa5IqgGKISnFFErRllfkyj8NM1LjZETZvUq7TZ/LKUFK2YMsQAC
7dwd+TVYs1f2Ef7l3f8FzPUmNOljAIVQ9Xn1EGU38fZc7Dhsmwfu8jEXqiv+dwFm
tlsS3Img0GpFUB7gFKqaADgKiVXmwBbOE+CDIIt3Qeksp8qW+BDMg4HE4m/inv3j
/isz0cQuX6D6Y0iZgpGjQ2xOuNYW8jm2kv8KPqDTP0BSI1YvYCDZxf01ev511/K+
baITu4hJWeidp3jt6uAw9CwMxPhqJoP1CrgKYfo2ErDUxsMPIYQe8z0G4xBPTvHE
SZyNn/99RTC/67uok74XZ2j+keV+hhQYucV0EHdgrKO2HPTHud11bWdAFucVjdYZ
5zWlZlE6UC683+Hodp2j+ByfGJ+gd9aUcM/2omT63TA5Q0m6L9UB0y2WTqkoVHXY
5bq9sAwId4QFD+ANU1PJAkoYv6mWxd6ni13V9pYrp/UMZ9kKuuTZcuYuxp6md+WL
PSKDYj9yNNHqmUna15arApsg/wDBuv3QRvsh6N+zSU6DQtZkb9LA44vN5pnpczsq
d6kacHgwvnxJ1x1f4bllnhSarQ335wv60NpgJojzGZEuy316+z1bgbMHoulttAT7
ThPTIL4an2SdU0dnfRLk+rrbX7dQm4EEG8gNLhPi/bJEsb8Cq3LQrXF3cAD3sC+6
tuXxaiksizaNtp8YEljs44rpxqZMfds+VqX2SGXGzE65N6zE82f+5RKfno4vAqKY
6WznbfnnuvrwSJsr+mc/8PlU3BQLg4DLlevL/isi4JCrxEdoi6L6wpEG2XKlS3b6
8u7bE3rhjPjfMbnvgkCB8TU9RME6xNoZem219LQmD8BfWXu0lWBodH2qPkIqH3GX
OJorolK2vOIoh4PZ4zHb/0Dr2usvMnSDkHxQ/DBVUp5BS3q2IH4GtD/UxNp0UnsA
ebrhDNi5qi1iNuzsrLncK9jRorS5HKbO5ShoUmYhWaNev1qZo8GkI+Xa4B6oWpo5
FkJoGglEF1hl7+jBZqkLEbblBxQ8KCShGMBYl+zQmEr8xoPYNfF47uMu7UC7bSKA
YEURCFHdAVvu7/GqguNXfDWM1AFZgDFlw1VznROJ54E6iAAF2vZLXcMBV7I7LuUO
dN6vPPa2tr/iqtvPKIiyNG1aF03FTSsX4ReK6mM3k0NGH17+e7Byn7018iZ644pw
mQMOfu3SbNEclzDDBkpPqEQggCSwSZdL7hRuVIGgsZ7Ww02a9JFGW70hBcpxvK5m
z16jb3nGuRYyUR8EqxgH9cwSV8BmC5XvJl18a2PHYsny1GXejpmCJnaD2KYnkcXq
IC4kDDrdvoQ1U9Lkk9zuVMwaJC+aFUAAnJEijNS4JpjGrRWL3N2xavWKFV9OqjjH
ehHcfj1S4CQ5cLgO/hHWjCQf7rXWcUNg64j29EgFJZNrQ5AhPCJQo3MxbM18uAsT
cMjQhQmHRAO+L8SyMIaJBxQdUlQMULZBaZ7gYDJ739tp3YqlNN3A1lamhL0SaxIe
M4/cMaimZX29jtPcca3U3ETV51Ixo2ygyuTfRsJwvBOqUdBb0Amur/jjf4qOZVNA
RJ1H60sXFvb8yj/LTI3ZdItm+F+NCtJQpGOZgxYeKpN4QPbv96OXxXkWTQSQLe2I
YJrVX1MLm50R1EBxM7qtCZBABI7CWj+pYfH5DeRryDo4bxV6gQ5A19K7YqELP2dI
nSgc93tdoKgZR/MGh/sej3Dt6KiReM7A7grU+Ls6Pfst09T7ppFknx/9O1M1alUx
KbgjjblWKJWVxQ8fuMHu7Fgu61aLprEdWwELNkmfcbqKRdoeqQzE+MglclrrEGxX
ix+dYxTO2eEx99pR32K+6Zw7xhtqc1HsiE+ph30KhlCTpOpkJYMuqfK0eohjccDw
+EhITOvOTmyji+e1j/ievjyr7PLQ2CbncsL4adAd7/oMsrdCv3IWNmOr/YLSPX4/
GBvttNv1/HfvZY5O+P0RHOUkYv6X4mGgaOyR17FuUryR3zd4lgIDjJweVZXCwJFE
zBorz7IxA6jFFnlPAyr423HbtG7ewRRXZJWvW3/IxJJoW4udYcQMi/4C7kiprwC7
pdvxKK55exk9FDRqoFdnvWnnh/tEh55kkzYfTtVkMsXvIT6NfWC+52T/6JDbj8B6
bUmjKnymVMN1KNF/DNh8EBcpDUWF0vC5Ztyp+2ASFmPr3i6N/k3IdE+Yw/AENmcU
hcXEbumRtEBBVfjL8813Ra2ykDM5dzB14rjhlO6uMU74w19BowBYH1o8U3OIdx2g
gh3PrX+nMEbLjlMMIPhOXbi+uoIZg5wXx9Hn2MNBOoLqCAk/6oGiqvwH063NjkM+
d6u74WQEEDccSvFBy/sLIUN6sXLnT5yT6DFgjrUXFr6EyHtGQj43m9r+XQkmCkBo
F3SEbDJ8s4GPfnxHkqvAVHH5qSkSRcAgmjWMX6+fw8CwLnUu743hSwqnHtLRzLWT
YqZD3iEs0QVopDey3y0MnFjL0wVPXQ8yy15zquxDWvjGgzrRZgLLQh6JsIDndtGS
ax5x95HviFoFG5wKb7nRsSUN8mLVI2xW+JgKfUJAWBrcSLc5U18oCGnOiRmw9Bbc
E8Z6A1dqN3veYd9vOl54FPp/zDAAwQ4qTsKf74IQ3EdDdo218gIBwqYsMXTpyqyk
TuEMlD+fjIqfWTxMxygm2UmNR0iTY9k30lzx6zjOaPVm2VlbtllM6nhP7bFWCIf8
eBnKjy68rdZ8II//G9UXIJnTl/52dEaQXBRhgk27YOlP90xCHN15XELQD3PvKh0a
zPUh2e+qp9AHZY1biD2sPw5p3aUYZH4rS6k8s/khvxb8897jCFw26qpANfqp/ly/
OFB5mcy/+EorY2ZzDV/rO3GN45hytwpL2Ah8pFGx1PVk5tF64Dpt6Q662Je6CMEi
XHseqjnhGuDkKAE0h45cvAI2qid0Af0PAtZdikIFVGj5QJ/X2y/vePj7ljRnL0JQ
XHTzVpeWJTe/Xe7MjA0qqGWiRCzYVOuUT2bPTa/sClHd3avxyHmToSHhr6VBEfC9
K2Q+79eJPxp7uaMraHJe8sBu8igtt53fnwLXPae7DS4M9whBj4x3iDOBH2CoXE1t
nEh6HwUZAtoPgssbt4xquNU88UGHY/kFdMkgo6kPHSW9ozhHWLoD6pG1EMaKml9n
YDB+iTV+PYUtCELY6EmXJjjCbBuoytCZcUburd7QDlVEBbXIvzq0n0ZGiFbeCnnT
c64gGU4pAPDTTB3DByD2Be0Y/l2KQWuWix/eCym7uMZCWQdX+Lvp8MCpCd0JW8Es
OmMweVl+KW2ATVS5uxhxl5f5sOZeL6rZmwcHbV0YBcKSi6GRUGvoLsEC3J1FaTU1
dsHbHvRuHnqKgUYP1t3IoF6QHorVzn3oRPwY+edFy+XFJUac4qvANP5pL8gWqdC4
OqcJp0St27nrJJQQI7s07IgeFAtrKisnONk7sCaINZ09X+l37cXicrJYZRC6iqt5
3n7GyLnC2hZizqJhT379dem4lzVf/MN/XMaZ4j4TrQW3QgS+3IoaM5Uh1S5PCZF/
4LkIQrXDLDgvgmU2oCRpTPGaconhCmFM9k25SEz89bEUR8LNOT7YeKsmNBwADSvU
2yLkLS/QSEbHBlO8IsZ2JXvR5yQSA4+aD4y0WINnp3LnuLms5IqBT4dhyLnjrYZP
U8Q7zIPUB7QsYkDkxhBZh1PgQRC2eUj8dBZY2cxy5+cU4Bw2ogeJ/OneXawvn2lT
xXRA2qoizWX9viPa+LRO1ekTD5jCilR0icWmfBc+2P3406VQTcZPXnuUpUqRiRTK
WvAWON8QpWT2PaEQW2fQgCPb/OgnekNwVEVmWJXtFJc0qKHHs4M7gAAhUQ//80FX
LuncYDYWBIip3aJ6o5Bd/bjQOB8a2FvxN9RoSkNc/PweN5EiRo5CjYOvTn7OlWqb
FbB5PxC0xIZvAiOdkKTUtsVdJ57tp7v+iCIBj3+L1T+r4ezEOKQx9cVC8FwcMYwn
icTS3E8HcTkE67ljVsDVBwzrorgDHy3cC5AEhgM20ETgwU9VnR9sGnAAbtN4ITQT
oNbAOhc9fDbyJNWx/2L3VR21VMDRNVZ46uenTyMMQ76HvDU67mOHqUFHJ4dVa8dO
idurMda+OYrHJQc2ssLVEJyS+4vj4pGYmx7Fp2maHxxOUf97dP5G9+gLrMaJxjcV
J6fKTlrj+8AOA4VvvL6c0yaAWgceOgq9/8DpUVkEwv9kJGBAIjiayTinhhz+Kpj6
ocI01afU+6G7EHU+XtTFz/46C+PogTfZHLN1rvAbmyU+7AYu9uWEMID7AYdgXndX
gIWmSonbVwV229ffJo+pmuXX/ytYCA5tE7DclAq6+u5/Yw+gy/7slSKrO38g/GIq
xuymOFEyjVt3B8dYJykwFscj13ZwVu+s2pIXTmn1S3wxf3Sy7TrajIfxNgTYxvrS
nMAcZWSMDjyX18gZkf9p1JLBszaAGNvmG+QQBfAd450O3jXYJU3xnq47U5HU/cZJ
qxsEhfwxL/fkvl3o3gPyWMrg/3Rg5jZFVqyI7ypz/NxiISvqxFXgk3V8X6l55TYo
hPnAq0eKY4Ei1cqyG54MNNWio18wzmHhhxHMcT66WNh4zEBgVaTlbG6xpHtRgfZj
xrawUVBoddqAgBV3KEqTVEdck+xGV9Z+CuJLM2VDl5hAixiGWo2YFdQxWaQs13e6
TalPDQlRiM7dyWuLxy4dyr0H3Ybz8qPDDmEGBll+PYGrM65XHhmnU+tTR+pKOHqy
X2z27Dw2VylH0yraKinZ6wsvnWAoKk15E7H+X1Ui941Mouf513OEyepqOzsk5XsD
rQPvFshBKRpL5zoE2iqfkFzg1eeT6zkNuaBVbkxlUjsWDUcFDwHbqGWRSPE0Rl3B
pfxkEZvxX7Wwqwa4oxQKXAzYfgcvXNq6FZTMWDOYh540UqdV2bcAfqY7X+MnTmSi
QV3L5RkVBmZ3qaM8Kwsbrjn1h+LvcDmgtAZvZDUNiQ8WTxE20lGQxirJwaYPOFAc
OphaQl85ui94q1fgvJBQa4DNGJgpa8rt79OPQC/wzEuBt6AdgdhMCg+n6A9NWGHT
q05cFjdNQggQ1P5KcGRAKFBJj/QREtP/VMH2YAJTi4iU3eKWbp2iUEztJJrDlR8K
LLJN1mItyvRNvnOBnzwS3+TVKYNjbO7i+kEDdplaYE4dNqumYmBQxw/7aQxGmfmR
kXGr5WiuHkSfin30HDtKvq6VuAehXjwukRlcFjfNavuyKfwIbS7tTI56YaNfmH9F
rsmBrEfw5LHTtR8jO/6dTzgtGXo749zqHqr4kyV/VsfbKPjBQ76O8DJ4aEIL3Z6e
n/uByetSTYoyqqWfmsv0PZ7F7VygZHEBFvHKZJUiUpsoJuhTCu1roJs6v0p1d3zY
dp4EE6Hcy+zsujzOsbSCO/Z3Hc+okFFUKJrcUobqFrU52BL88HPg9EUR3tHAYtIE
C0WilrQcdJAK5wtC2ylcZIAR1vlGRuzOoeaoskKlBAX01hDOUkrzXTNpR7+mXcT0
O3lrn1fWIQ4OwICjr0s11zBCUEmq5mefB34jHrcydYwFMFCKtIN8gfdUdR1gsCah
CbEPpK61MkHa1DgvdTQESNcAjBrAm3+WxB6ibK03NXjpifYteSIBt2ykqvalXvgr
FLecI8GVDNQyBRIbvPLuow/mOuOtkp02ak9xO/jYIHUZU7BEuDBpWO13y44jrdld
azNuIXIP2LL/tkhJn169llmLT45Q7boP/lLAJoK3Z3/SntFYw+8aOs62tCUycRhg
QVDJr1saRIwANAOOGRKE5qhrFiJaWtHn+TjEAJ2FV29b/2coWCjxxjcmAyqURHH1
1s3Gk574nj3q0+8EGycIjo5Rg98xD6/gAL5zM1eHR4dCTWvKNkh7lIdBN06fbSTD
J5OFfLdfI83It8fnNq8jO56awoIxO8w5FvihATk81OYrijF0l436d5Wm3r1cuN3F
kJfSQdlaE6llVmF3nDOMSTnBVyc1QhZ31mX28D0VvR61XwBFY3Dqf1BuN+Y0XWuR
w0RUfw3Mw85sVh/a6ZxpMxWfl3N+QfkvJru7Ve10VvkSP4N/YKW9Hi2T+jhWaWRk
3A4YEuhAD7BV+HFWlUJmPW49lliMAJaXxnWVxdmmlWUV0DZ8CXEuc4+z9d68+n2d
/By3d6905edaD9oDE0s/fZsLgjVEwQZHBrO4ngVpAzTkHhNij5tEavDqOcCUnC9w
UXYCBuNsX96+ploP5BIaoHgXuCGZVowd7L4i1rmraPq8NkYbJge+9Kco0WFR2Euz
lJlOZcHEcmqTYS1pHrap1C8sE9UDanaHEBN5S8LmZE9Jt1fXXDXKs3Mtr6VBa4sy
YI4dgwLi/zq/SmOzly8Bvx0uhP6mfJ57yqTosFHFdfJZBUrt8yTEELJF0L2YcQEN
ABv9LexK608oJGZ8jm+A5YHkXmqZ8FbV49MijEfKZuAmez6L3vy7VznY3w9XcSss
T/drX5rxX39YqAdfsYOkHPFEJvo7g3vAVLW2YsbIwDnR2jVJIOkWUKn3fBOPQaCU
0vLMgI63TC3bH+cpMtw5SEwUWCc8V5OasmYawWgn2xkjf1yCaGZzW2qYWcoIp0Sh
zMY0B+DpkfLZ9qjXhXd98l+4IPMCXdURJIFg8WSoGPAp0+sMMRHNFT+IwRT8SVpK
XX8apT40d4PG0d6xe4LHO6zxA1loeUh+n/37hRQsm7HnHIGTGOn79Q8IzPVw05D0
O0+511WVISC6FLBCmMLm6qlCCFd1HqDjR7mIpqozyrHaGE680wYrPhbEuzATu+Dg
wjrOLhEj50c2YeQfUdzjwAinPZ5pHfgdGeqe0iSVLEMqjvuZ4w0vyoBOzsPVwM7K
OjjvnkutXJa8AcyCDO1SRQuOZoD5SjhIrncQ70xGWe/5D+zyybBNaze0gXPPhssb
Dkyqe+5oPljBLnamzLBdUgcLGS42yVLzW8Nf3LXSEtRhw4Fu/XKEUMOeS2wkc9pT
+h1m6XjEHgoY1mir58b5GfHODWMQYK4SCl1tDPANXqyqm8EG9FHDKxk0+5OfdFPC
Cb8p4qecW6y8loWZ+XANJdFJKFQyfNG8jOilGTrJaqamC1vtdI4MeLEPFd0x/Vgs
mVRJ3uezW6IIdKc2f25ARQIz+PQ7HdRs1uIn5u2FD8DkgpqlhuwjCOkCYy2HfFIo
B6O2AWkqhau/ycCPoNx0bzj8hJIpNclpctOHmOhnKqR9uFaczPKki85xDimiGN5S
fPfG+7pH1Aqc2ft+k+D03t29wVAl9enLkL0n1303zkeMG6m01+qsuP72EnY1ZZuS
T8nJuiFlJil/44MBNazlFsaxbY+sMuX2jsiRgXN2xhHqYNA2K1kkRY5utBOawkkd
/4FR7AAB86iVcdlyOq5CHpkkSF2bBR60am0A0cX4hhZHAOiEW6JH8AmN0JJ6LBRr
gP3migMsSazttYfFek/cMrjoX1aC6JG9RkqMUgPVOFXAas65EjRnQgq7vEp5kc+W
uDhj98QOmEVxDTb2MKn1rkeTsHInuVQj51U68oVmIgnE6NmpUhGA7Gab5f0yOdOh
JundUfH1i7SqIqsXSuW/vffU8mKmiJkgoFHScewIMKxWCWpD5dQWPPsV+d5GoKDd
I0+AjtNl4sA2Du1/jA3IB2zb8NhFsw7ql1jMyUph1b3ra5SH6z3MS7ZptEXfcgIK
WNPaQfHZp+FZuqyEzvNff8OUjTJPRJBb2UMuXUe6W2zJt9dxTcaYu/Z9MF4U4bgS
SWXBE5WU0s9M7xFip8GOMn+jzwq7lsTMZteTcq9J+0hcxTXeVgAKI9z2i5U4GdpY
ZZxi1LIgOetwD106DBXrEI045fyiE89gunan4UmvL4aHIeKbWmf+BY9qUwVyLUWu
LN9IevCfjvoTzrDIERKOviOtZhZAVjfZKiqGiYqHE58ju1TLl9UGHxKKiNLo/N9T
gKLGJe071RD2pNUH+dDm9VrPqhe17HNKB4hbxJtA8oHCNo70Wvrt2vHoNHsVoJxw
8ESxBhbZ2b9hg2RH+w0ACJOxvgTidln97jWDy937zPnvhruibBiBIWGSriz+nFZ5
ePmdAXBNKLwSOZAaxK/ou8SdteEI29vOvb87+sMD2Sh9RUr9pzRbIa6reJA4x9pZ
3tot1IwEoY949ODs9HhgE7dbv9Mx+jB8TtiRkxs0Ey8EZnuBNvNjVKI2ZrelI2n2
A50k6GFzVkT73vxaTk13vq0IMxl4aiwC7wPLttNISfVHV0Gd6DaPvK6jFYSwWOVI
mCBgWGClCyvF3fR2yJaXTcEeLc1QG9OtyjrSjfZZwJkxWh6bCFMkTf7/V827EDn6
kxf++YE8QygriAQkjucxWn8HzUUObgV8zITbf/dB6GL07XOWz5jiGSB+Wrh6mbAG
YXZPlO5n/wfoNFf2khC/OqI7JbyleeNWEepLDBZnvRuFvGkk08IggEv8Mi2+fMJ1
5N8BfkfCu2B6OAoIuMclBozOa23D8uzcQHdMaQlxrJLmh/T24vmpdpSnH5acmzkc
ky6VwYTybBLFcAy7azokHBy2JvVk5Z2tVVpR90ejCkqecVCyG+Emilza7d8wpLHk
TYezQXLm0+MRm/VjOhjskD5/ju6dsm4Ayg6cFNmiKzjuR1jp8t5tHlrAiljOymnc
5R2vhULwlNin8dzCzefLjjmcQsTHeolJSFotkXScvEyVleUq8ODDieTEKDTh+AsS
29BwTt7wGgxePowfaFLSHH7WuqvyIyC8l7IAZeIIgzRmGGJulMu6zJogYIx00FZ0
NxXRjQTo8TTIl9wrJkUOHfpK9KMASgP85zzEa2eaqh8rDiVR5rphqgqX/1ao7gJM
imUkN/WTg7VbHzmtde64bUzfOUe6CVdnq3c6bdPU053XsgY+sPjehRZrr+ierlo6
GepkK3bdoX/HmKY5T85xK5sJljcN3RngOA1iXHiglWdPpJjpfFXlni82H5GLEt4e
DQAmnHl+1eEUSMTvv9cChTcoAoA89a04pV6Zv8zy3soP+FAK9RBAzI/utvWaGI0O
Sa1YmSTW6smhhRVPBzqRltLFK7wKUD3Eb+r5qe/g5NC2Og20YbD2AGQmJeoCL/fU
gXKPuRee3J7utCNzDkHwYLAsrCN0ZEbLIagmJIwdJt0LCWWrqSADT5LvkBqMxf8p
1O+pD5BI6ZcUcQxt8PMLchoTSuE1O2Zffc8lRPGDP/RypfsT6qqGFxfnR1DgIRwb
mzwiq41DvewHPe9CDO+gP4+TZ2AtWLjImsjHyRHR9D2QKfZSEFqmTkgj2+0q3ymf
Jd7xvYOAZ6BAdCLiwdcFmLTWRK2rJkI413X6YUU2DQySd9D0iE+WFdgtLMHXMbbo
I6K8J+lgiKEPYH+LO6uZEiDxmng2GVgfCVA0v9sq8nQ9ce1VjGHE/nXOBHza9tJ7
Zbk5WoNd2pZr/72CBL0w6yZIA5Z7GfEZSPCVeMErkc8+ltScMmi81BQiiU67u+IK
+pLlU5bMYfP+dqVtqsP8UYxgCk8xVi5U2SN20T2d4/jqdogMl6heqrwINiy7sKTk
N3W/IYA7iYzpgz5uQHDXze5Jz9I2n8z3WbDCrU0robKtaoac6Etfw36qW9bZxTka
Yfs6Y4keTfDu3aK0aa9AqBfUyvEnlZdraOSeZ5L320NVbvpRAMEdANza2IE8cFOW
xuJJ09JY+vCLNszVS5JWsiIrkMYM2fJ7q0DS5tAIklnQtJLmdWMsoJ/dw1mWPsyV
itWHFc2Yj8l0mOlgMelqflPzkc+c++4IMgCGUFekyEqwHL9fkKUj/pt4M6vVm/aY
mOJyl/6naqxSTmXug5LfXv4DVS4iPKiFQFozGu4pZ4zaYQa4+6RH0gDs2WzxKUAH
E9y9NbAG6d665BDYsT5+7XLYdrdviEI7TwY7Dqn+ZuEQppunIdQNbcpXgNqE2noi
S7oitDkrOiNLn/rRymvSyXSp1g8+0ZZBk/T0byYq36bKql+RdRCqNXsSqxv5N02v
K8cvnY/QmltHgmBl8/dvz26AiixAymhCkwM45+o7f0uIkV48fkVOE6gv/zA0ERRy
wml0tvCAESY7P8nnIYnlamBxjLpmizk+84s39MCaIa27Q4Kwz9M+VSfv9tuD7oS7
gA9NoSgolYVuiYlt6/rz92Qob8ukjOepadoSf6Lqw8RQsKOuhx33nDxHoxkJoqcZ
rbcwlOS1Q7vIAVamdJpxAQsEGbceEQ4cPU0mdzxWaOKVAcXvQSz0ocRHOKieEznM
cgVg9SXcg8PYp2t4eB2Lm6wwGffofJSk/c5KN1M9MJ1kRertfHj7skU1N7QSr4cZ
D9viYO+LH7/0xmLI0cIzipOUkgZtNu+eFePk4tTTVkrVrZsA6wBIHp2u2LgEIswD
ldcatZTTnRCbFT3kGn73JUhpXKUhcIkhg5PB+BsYFvQro4ieE9udgdF2B9PIFBuo
tjCAiflcE4Vv0UCkkqjT3ykvtL1NAV7IfmAo0i9/1Y/P2ZFgB6kPmbmspxkzixJY
vkocZ7ZvmKL3W9h3KpMmegqLvzwzspDl9ifPPxbg5dh6GU/ZSJagvUPR4+3ptE/m
grgOfabpKzXsmabkSwSYSOohbObhvKifPwPLgC3s0H2HfC2/wf3Ij6IUJc+EOSPu
7V5/MeG+aRMWPudrqWgpCaDoHhj7MpBFJqPF6775XeiJ3Ns9KW7NR0brRd30S/nJ
IlrKiTUXPgAswr9WMlHC9nehbrlpvrzqUdoNk900wstbc5Jtiu6oQJXqcD2mKriz
oq0E1JS5qluTp02Fg03VxYmWl5NeSqjhDCcQV/LRYAhECcxbNWPRJXiDT/vVfX7z
TY7BmFixeXsz3hd1YAXYfUIGhD3bMKg8XH5Z+F+uzRfmG10khm02CWvqcpXkNT9A
+pZUxTLo3ZSzY4xGDhvNjJBRUQo7YuqF4tystWUosT8wBWJYAuxbcuYAUvSi/PPc
iUiGReeW0oM0GseV135MO5wEWGWsFTt9tGal+Zv227u29RdFtjZbYlO3XqeeKGiv
0IcNvzNWPoiJLYqOC+OkfKK8NgWQa2VABRTQByGqokdNzZeDSlrxjG3bJGYMz616
T+2rB8qAhdnnRifqYY8CaNcmeiR5PFMbS57EbTI5qWYKbmZnofNEBRLR+pTbnfqC
kLd/YxTMvfy3KZC9cBltEQVrheD9DOLGmny5ongTpLOViWPMO85VCFG8XFaEwJXh
KKv/jzFvm6/n2wP1GCaDLfCeKlHlQqqPZWrxwBySem2LPSZK9mSVs0+oALb+wGBg
wP/6nI68Tz3vfmw+0jnQVGyVEVxzlYVu+ehVniQFEU4IGBhQyCvAzBsS6D3lItHR
2DVh0JRfF9jhQ/zuMV+ii+7gl4ewUJ4EDlWjLQ56oMhVovKcZJ7FOhxG728zB+34
+Z4Qq6cinl8CnSM6XSvknU0AqHzqH1NhgC4YxFYH6JMLpj7Y/Ze02519O6061MRZ
RDNdanq+/3UBdueBvlHdcqSOIqR6kmbe3B5o0fq0h50v5F2ndI7XwwHdqi8cLeZc
gWPl5+Hdw6OGcwv2DFEn/ydVZ0TmzwXveVU3JOVIB6ZNmd3FbfBc6Jjr34z9zvLl
+URQNtF7P80xwGsKwgnvmfLTF/KvJt1R6pGdO9MkOmXo8jR+gAWPukhFgkax9orf
Xxb2kIVjN776JuvzJywSDm1Ugcj0m9L0QhbOPLsI0sUmzEn6Z/O3X7HFr+plLLA/
9PtmXnUEEK535/F0GbYeBXBGbAZiOgK0+Ea3xhUXf/ynZCbOC+EEmfBFiEPrZ59N
I034uVWql5rDHLHzgac9T1nvAQZvWjt3f8xDMt5K07rNQAupcq3nWqgTvKd6lYr/
sOi58NYLXCkVBB6XgTLYBLul08tnLI856uFBclohcvIKGS3ED3htVai0HLX+l9gz
QaRii5BlTl91EGdQjSvjhhCRVSi4/wptw+Mf5mS7IXD3mWYMDIO0mPyQLO/TsLrF
EHpTI5zd8GvUwuqKoq1iC7GqyVaNaLGeQO0Mp4p4+344dE4wfvHZdiOq09FM0Hq+
DStPdpSZQxW42QfpqV6s0Ei7hX9NSeA9Ew8GhwV4Gou4Ei879hdHxbL4bF6SC6hM
W9cIq3f5inXAcDKx100RfF6qdzAwGprhtZWBlRJASq1ZJQP9BJemRc3qcDSSBfS+
JuqEOUMm1dRwQ0gYt2wUZfVzo38Q11PQjCP56+hEjYZdF+ZIQbYacKKHrAL6X4WJ
xtk+Q9l23xKybWf2c6iFymaYzIQTmV2uNIJYpMMSCA9XmZtd0CVsOOHTC7QKRUrm
d9B7yetBCRzH6ksvw+DzM4ul0CKYmJ/UzvhfL2Ktj8tb9hUODmsneUD0gPBuVOyD
ixAPQgYJ2RChGosLmxR/FfjoELuoI75Qxj9ng6PwDtvolYREsquyitUQXdv7yXYm
9UPltmy4j+YUNyqQGq15E4QvN41t6XLm31YKGmh1qsL3Qw0KEqle3y7mi/V/9CkA
qsEL8D9X8qDUAjSG5O7Bk7DEX0Y6jynnRzOIgHU+35FZEC+LWn5jFvM9CgeTDQ9d
+P6P/kQH1gST7zsAi8+bbboXjnLVO57Q20Py0hzymupvXJmdMvCeB920cZBv7/48
BvABmK5E30Ns0B5ovzwL1xccOh+uugBwpT95wYq8TH7H29PSk1MyuqAVBgX+rZ38
+dkvLRk8gYjP5YDEEefnDZx+2IzMRKXCo4Yg6DWhZJ8zheeYg8yIyZgtVrv7bC0a
6wv5hepDGsrArG0bnV8Bpo9H7J6zGgSADm6bP5tEmuhyK6lqCIjwJkC4n+MUPinF
y2OyKevHbHO39xeBHSVgh+lmo4qZBC29QLMhjad85kbPQGqOhgO7ZrDeihZIr6Mo
7ZYnzJ1qWLqajyzGenx4+Pu1gzlLrN64zuGCE1Nf9i9cSKekx9IgB5QG88CmDj/1
wP63Yjr1FrEv/deg+3hiNklJFa9rJwQJIcsA2CgMfQQe0hNHpRFmUozezEZY3Ohc
Dbef8jiLcsS9Lg4wAt3VhLoETFmCxGkzl98AE3kKxKx3Z8LU12lzMSXOVUVdnvHt
pkhY63FnN/FsMN5oaZNWWu0NEbKbdbPdExO8U5eFV2kJxvdBB8MTzthCN6+VQIBC
Zg87QIrupZEgNPN/32EpFtoLcX2OYRjbZF1QeNhyI3Q8o5JIHsT1IexNABrJQsbL
eTBW4egUGP5bsciFM1jrlxjm06bEnqPk8UQw7zsuAnr3ptbxpkBuAK5UnAtfL4VY
NBIIJ6ZOpAGwuMu3DzXBp5CNsGtYdvf2FEz3UM3Sy7xei8uKm1ASF2r5MB1vmqcb
2mZc/Ih81x26gb5YcTPzeVuoCgu4Sav61rURpInlW/WMVunBCvn4yyHce1LIlTtt
pUTSA2vjba4S7e2EhFG4Gsj/0BN04UvgBSD1RcKz1GstvDEhOv8IhY7vnmhS+uN+
na9XKL/HvOFClJWmhXeX0py5eLBzPhlLQ79Sssl7MsFxY7rs3DE3PGd/XL8HB9YG
bfZUJpvpQZHbyAC+XTNAjgr/tbca/P/t51KPzVTNlFUGOo4tP36U8e02wdyBOuU4
rWNgLvhPhvju81xwRHdKbExH9sn17k5t6YKlhaKB+Ddfol5dy4L4tm9OXGcxrOm+
x9oUSNIpRa7GBm1qreobOJ05UKNJ+Hu2Nt3m1m6iCwwDDA2z/tOlLIY0zaz7EYkh
nvVwFipfYL8lbiOaCEn0lI1ktXH+eAxzPc/wV5Vz6CoQ0MDKOCcLp16Ek0vN7Fty
UcXrYlIzAlaqt59a9skIRvliOEZMmcLDNMoItIZONvGlWHVHoZ3b8/1LXN7ixsnd
riSCGy8z1mvVO7HhglM2vB46DwrZOeTz0HR1mWQmj1Tz3xJFhsrc2YeL48PZRDN/
hBkBBW/0B8+wxAwribSO1gvNSF+AWIBtgLDlHYF7NJPkJXRjt65N7VisNzUP2qkH
z3ZsiNcVuKx4BD/hG+exWEX9mki+jn/whFSPVBKxxg4GqbcS4lL6NaJoiEcjB3Gr
90FK1ReDHltRoR4T36V/Ep6/o5v9s0FB4iTmuJRHM9KQSd2L8noHSyCVH9uGwMqM
lrE+WxbkRdWh9r4RU85L4IHpmaeZqcWBVQ3W3SqskKBHkpqd+efkAdvomHrDBemd
4Fp+FtCNmboE/ibjic16qEp11/IY5IyQMVvvfl2wJYRwtmLldIkATPsy6sMdt+ej
CBDhn7ixtS5kaA3wmgU3fKie8ByyTbarJgCbSuX/jO/T7eKdb3REnm1WVUwOE+p6
wbBkwB6PNnkQa8gYZOr6P34fTnIrrr0xZQr5v3eWfPhAtprZnCyG42A3+/eTCCD7
9Hc1N5qxrkbOn5zTsQsRhFYf9CkoNZ62cAEw2rB2lwD+wDQvzn4UNnZuzb5+F4av
QEE5Td9n5X+Jdqz+Dbvg8zdWqsp6yBNcNccpbPvoHsvGzTWZAIr12nTIUfu8ZL1d
1BrDZgo9CoZstKj5XzYLpflp/gZPtDTzcRMZOpHj62RLFByMII6o1j5gFcfXRwQI
oNSkm1l2L8ONZbYcY/Hzr6ncH1LVv+EnThUTZOHCQzwvSLA/exiTdhLrTjgV/ikU
2mAyOaJV7NYf4KEFwQfTK2IYOP36opQ/1gauwiNnJEq33sw8hhejOd0eu4Crnlch
zn0Uehc4gEtXrBwOqWSXWCJikbx/FAByjImq6UChSk0fNbfK08fnOdJQ9YW/f3eO
I+EcGd21JWa5KTbQfoTGM5D6demZk/WD4kzvZ7oLqrgmBjI5hRsSBeIojXvaqjtu
hw3Lu/05kX0F5hkE/qiUDcjH23A7V4h35vRfMJlMEag6uPauztycsDFvehVxF7J1
2NquPw9vT2lVqiJKiO4bo01mcFzfckaMuboN2NYT99IzM+exX4wvczqAdhVnM/t5
lG2dQwsqe4w/LzanNMcVS4tcj1Xjq9GTHAaKn4rXBUZkEsJzM9d+98puXRpRQt1p
E7XVq9Slxl8vYy0FY8iNzPPpX6SfDvtuIgkG1risGAJVXRYmxx0n/5dfAviHLkdd
8ejhDNj67XMJvXyEvIHCCeiPJTA2q3d/SXHY7XxXEbSzA/L/KapZvAi+6ejTSMdV
MUAzk/6Bi9wKmfGpxixE9hwOoHI7QuK6/e3gU69RquDhjQRfkQq63YNqTWry6Qmm
9k3mEuQ+pU9sbXU2gXer7JQB+M3y7/aEXx0u5fzYskY7429wB3dSSuB+iPNMFmoz
058YHPN+pAgr5fENbJQefVtqzomu7Eh0jU0hItiSESTKp0Q8XbZ0BkDbpSC9dhBy
IHai3h7lewVhda0Nzjq6AIpYHLIQIcU3OmQcNSmZqo4tmmbTLtJeUL/8e5Pnfm8f
lkqF1PCFzlS0VXgdSRVoJlIto5wOXeRBUNKv+yOpMaIE6/lXL3Otzyj/qt68nK5k
LaYt7ry0Ddai3upa9/sENPeiWTnDrJVqnVsgajQolVJrWVMvx4vPmzG4hsbeC/eL
NQgUHNeviJP9/goa4B5TN8H4Y31Oi9S9zFcCy+sctpZhGAtsEwd6OYwBNfTWA7gm
8kmyJQ0ObkfbELGXdXEyHke5cZ2tPuzKLwlpg7+Mr9zP99oJC4+rQ7DCx7nh+cNY
99OZ9/CV3VVoOJ4NLJOVkWgCumcJibV9tbAeVfRvvdAlXWjNw6lpl4eni9jFai4I
gd6ndI0Isli/Duje4vMvm+19xEW74MD+DPf/23y5aViIRuSOj6Za5KVuCBDq6S3K
kNRMP//TgLbFmqW0JFyqLRqIFvohkVtwjxq+YCkCHmh1omyaYbQlHagec/toBUt8
8thQyohn/LDrnLEHh/DyuctPlesrdAvID4kB/JO41Ll9cCOUvAosvnx45j0RUMbn
5t6gFGdmh1PDRQBevBDDlvMqwzLf1ng2feZngQKmbuXhcb70te7doOT3i/r6ofhZ
LbbqvYrc2n7V2RYB631MW15olHnNNV0pERKLQEzrG+Fwhrd6IwdQ4XeZACXMG2/r
9Knfe9NqCy0RU+yUsEpwMai6D6Vc43vM5RlRDCaxtOLRorabO2iF8ojPCwEkrWeJ
n186AXhaVz9Q1u6TX6yFrImXtDE94oZBydPtfwYbHQfB08BjoxL+LiN2PaXm/2lf
9qxAwkxCN7meAF4OKSsrY9R3GeZTW5GmHcC9lPBSdNEM2UuH7mEGZr9/cJkFX8tT
Slkwr/mdWHNrEpjORzDpzFadiXCnVLTAJLFXx7UJ9e9B52+9XnC1JWI0F+XEwZk5
4/O4yamlMUeXtGSTN0EcIESvM5pncucM0CRxD0LkDylnphR7a47QSDmGqgsGHGGC
/233DYhaXUrdsAX5JkCb1EGsf2iIxRtC7jnvgV/7jh6ejNmiCnNLdv4uu5Hjg1Mk
saFYTGOd5iQ8juLgg6v0LtwbF5BGaX+6RlN0qCqZW9gjQXETsOA4L8Ge+9xVJztl
kcTgZMzMxTyECMWWp6DoUr368V50tCehBqrLxVQma0cwlhtRdHBb5HkN6022GkWA
6i4+5jueFOsAufXYXmAchi9SA1HoRTP7BEPt2fbZXWR9myvwCAycut4fCPLfYLi/
RUkv+9bBE9MwkKHCe4hKLZe/Yx846Nk/eTO8pVLkkuPx+BfuBjuYluRRq8bANEpG
PFby9ii173kbDX51Jl2LKztOt+gk8Fg16s/Ol3lbLXNI6hoveBRogEtYBHdajl5I
BIDx2X3HoufTW/JdU9aVnJ0vXtZy9fFusbFZn0pe9DzEG7Xa5e6/7lLRpDfH1cMf
8hO9eauQp+iFrY7rtBIR+WKNAfxmFSgOh0qfMvnWZBBesmIOLzr5sk5tMYLuZ4nL
u14AqZuaFmlA9VE5BjnZ0PU9Hgwjw7boVhy/MFvNNpoP5pO6w2LEBM8fMZaVkFiP
I0K5becfuX4TcTMJ2mSdML2hRWfT76oBjaI6qdY5jKaCtNDMu6B1qNymPmAkvhk4
qGWrURdj41/qLomQ8NKynMSCP6MSaD8HkGXvElKTuMXrYmKD3c1+Ho4HekpEW6sZ
6qTjFvaRprL+ifrAzRDDzK2afzJ4ozzHWnJ/eKBZxCeyMm/3htkZQaNMZ693FVlm
k9uA64WrG+vDEs31CddwglXwUmavB9voD/OWiEx+iti5zl4fxO8ahkzzYHJFNvWS
xtgE3LL5ffpLALi6k+i9cXJ3fp2ePPaciNz/VQVEvEs7CCcPLKE9Jy1tu14Flfh4
5i+TT8YhEkQH1YFDMmx+RMih2Jm/VluPv4yTAsnFdWkDWi8fJFXz3t0gaAi2lMwf
XyKZOTNRp5bfM8agpvG7ITv3iY6g5NAZr7pGHsBID7lSIIL/xCv/+0+7yx9UE+J9
mfj60o4fdlCtL6Jo1Nd3srO4Lm2c1GJ6e7fKGtbz9FtjpjTxikqSujOiyTh5a3Vo
P/MzdDLrCFBXzOweFyXWUO3N9Hl0JyEvyUS9g2ubw5GCR2t8EVcxrtukWuKG0XCe
DffJAmZc95MppYAfVvsTWUhPw9w4VXoDlx3GnJyQ7VwQSMGfzwcOyh09WNXICG2z
I1VVSARRHk3Gkft2t1HAhbxvxbaIHBb88sTF36CdcfckdQTe1eKlRTTmgIr6fD3g
XO1VlccpH73pXsAWfwN30RuSSbh3OaC5aq8APuMUCrDE56LqODhOm3zEJ07pgyQy
fmiNtjr5g3hrpUyFw3FzroIMH6NpFHfwdy29fcqC6Yu/CEMPv7hUBZj1YWe1GdOu
gT5ttJRtf0Xki9+cKtzwWQUFNC43dg/PXciGsRzrXWUZPIw6HoygJ8wYv4aKmGvv
aaISdIkAJmohXUjJ4yHpxTHYBgBfS7xKqL64f1wJBZUiRucONDnMSXZpyQafRuDb
5MCDEAlczBjpEKjsKyA0FfpCiYPL8m+cu1Xpzg+7NrPYTv1ejHSbZsEfUWkwiHDq
XEWj58VKqwbsISw/zNJc7hB3VIVcq+bzZvEwfQwAjZ8Oj9SJKp9j9VlonCl3HRXG
GiReCCgDy0NQ7CpTO7+bxdjoP1U8J93V5q+Dc+272B9ntXs9RopWr898FvvnpJwm
Lg+qhLtVeOvSlWHp2Mvv5awZq0VZP0EGchFzLJo/MD0CUhhzaVXxHwaGs37OGpcB
spsEn3OjjdLGhtpU3A92skYglED3rnY9VfLSJ/X2gMGAh15VzpCLbIbaCdwfZctF
S/6C5xQ3iy4+CW1c280z2MsKdD/JA2+rZl0O3RzttOe3MOVCeD/l91MDgxZ9iLY6
N459EgWj9EuP2Yc5VsCiF9jJleScIKDg3pywzFSlgdzy53DNjBosZvIhx3ZJjbSG
lIJMncKrUx2r8ukXlB3DbrMCSznxoMA0z1AXP5qLIKw6bV877ygZd4uHYo+9z7c0
hmZlh4fHg77KS8YABEaKvT9PdG7NV9e61VWuFSTSiIBdzyZ+M1acOeYMrNE/sK76
Oum7m9lqsgStxkwXNLWyj9c1iF0CwSLLTAfYJ2+/JkD7MwrsMLpE6bCe+U8BBeAk
/ktiuFMxmU7Hns5Q6MyHkN3Y/G/6J/EUhyK1mOrupX72hJN0gWRYqeDnH8iv048W
zyYZpqkf47OwvzICgZNWcLx5sY7/+TnjMDI1Fwn+S8wvQ4/WfEsCNdfyxtt6u27M
jDTXrqfjN53w+MIVRMvyofAKy99j75pYZBZj7oNY7ZHzK1OmRBTeJFBeAF8w4jrT
lA7yJRqFuW5DMXVS31UE1u7cFpv4ozbHq4vLqI9/hNkzLoLvcO3GeGUgX2d1UY0G
gKEmPai32OB/1E0DoG78yOqUlzzCPzJAeW1yR8AVq22IZOK3Sywr/pnTwojwMXCM
FrodgoA0BUy0ib+qrC/cXga0HpIUMeazRbkGX8U+ea7sjOa9te3WBsyquzfQVRQM
w5R4plAIiis1Qj20Nlnz99W7hgU2mlKHabAeUrm/uuGJVuKHwQg58KLxOV2qBWo6
1N5D8YehVDQbtfLlvKcP4CQOR8iPtc0m5F9okOwM+PpYxzHXxskGiVJA+mmsS6cE
PCZq50WDI5jBXam64AoGqLK4N6lCYjv+bW6bvKBV+HWuFXzFB1x/f0nvyNz7F0Qx
BtgPMd7TrkXTuiG1WLgQe3Ix8R3qF95gaeJLJuLxl4xJbibPCX9TNs7FD5/1/cHB
savjvBMEgVqN05Uoi4OxS7JvbvPaEer6cFQjFPeuhKAusPTvG7dwOh9YByAk2zMY
cXQyrM5LGOXc/75BbJMA7zJWY2SoA78J/xjm5dfKkmIW37VfTTAFtp7Aj1PHLx1+
CUMbnwE+d0r5e9+tFZShPCYBdnwfFZirTwkgTahRRdAAryUZjsdq5N/RCmtVbnBU
iH2Nhs1Uy9C0fjzeHE1eLHg6kfOLmEDOFm8DpG29tbBTMUgIVzrEFlxkC9F2jegy
xw53FKkoXDQGtDlzFrHG/SqKO+MFF5K920kgic/c8M6Ru0qkR0yLNyUBKG5JO0QX
Awn0wVQo+RraqsF70kRAW7xN0XitKKfkDNNtZbT3cpmK67WxJF8iAR4o1ylGtD2h
JIXm/j+GohvlpEk3nv7hlchkfCFZ7Sif98TOOMpeyWQcX8x9qqSzLNVHdxn9Ixek
cKedyu6LFc3Pl4Y+QeqG/ry8Q9Qso8MEKXE3KkkW3dH8E85MvwY8QuDeBlA742Ha
+0TukDZtWhrtqY77iHiJeV2vG4bhxfQE/uF7jWTwcuynqXCtZJnCY2SfL48LPodk
eUmry0l+j2JU0XLxgGPexE+6szR34g+V2jbIBWcrFn+I3v2yMzF9EbjV4rcBBOxi
3+nQ/7WkaWH6QQk85PSS1cDiCXkFtDs5SbeC1x4f0fAnwa0znAxPcg4Erzeax2R+
976oTlOKlOnjwSUR0SVtgdT5YPNDdB7Mf/ePOmFaefGf40yze853jxncH/3q9CH1
oOUCuReJpgXhk3AyhOelqdc3NtWaoFCKhka7yvMRDARfOElvstJjl7WQ0PettfmG
1JrlqraKEdrdOINOIFDJdKukdJDIS0J5ER35XhenFps66mkL16FhKD2TFaAa4oCc
6Ll5lQ6FW7JfWzH65eHqTmb1+FcTgXtkv6C26y/y9qiVxS06Ei1YrPBbC8Y4FSlO
WgipXXVOQBPwELHvKotMkKmMFA4mG30BU3369RuG05zOXfg3ICoDwma8ghOXUNKG
NyjQrrLIkVlkSFXdyZEirbX4Xu1e2RpMdrbZ0yV+7NgwxzLjIfOMgIoLZ621ray0
0dBd6t5WhDiHWZFgu9JjUSVQam1PINQL1AnHjWeFIfUAOMkZPswCRKRegAsxukI9
U4PCP5MQ8RNu5AJ8JL0xXdq8UUA2tyk9OIltEbWBli/BLvBhVYJ8redGNcHSc/v0
lFw2FXnnApsjxNUzxqYc7qGEk3keYG9eOrgMnvPu+aA91bCmHG0Ps9GAqmRvTKT7
QBBHHy1yhAfPsqViagHsLOmDv1PaNGmcg1LnliTP99Mtmd5FD0ynpFyIKUDJnAkS
zUNGvBXjyhTHByBGqRtwo8pR1cJrZTTvtmjSmivj0NwqmSJEnaqxcrkmvDABezZV
Sxzvv1BO1vIannQplFCP1RZeCfNQXzxMuvGCvoiNYdOkTg2OV0pjqhB7AY6sOSmq
HaPHKEqRUzBZv9j5/wW8jc2nyPFs9SwPVSD79osUU0eyiGajHvxNGHo95l21VKHE
+8dSGOHUncphLo2KndE6MpXJ/wRRA3w4E4XgPoCE0K+dmsleFbb9Gmd9MZCLYqg7
vSK15f6c50Rniv4/DIuv0Ag9veM9UrTT70p47N0W7ezY9LAvl9xuoJjBRWNsKq95
h6+MhT7b0aNNzc+Oenq9n4mjbhHNVtHBVoO11bKpT6tC9WQYcPE0Ql34gmHcavMJ
+C8NENGtD36IipzWEwzPduqpGUn/lISzuM1EEdTe0+EPdNidomri11rmY8Uw5r5L
PIp0K2nkV9XIGqWA4CH6osB9QQZ+2rPYnZ47budyLpHy9g8qejnr7N++LLLE3yK6
yEVseMts8JW8T6hwfekuP5NiqGXwBNHpsD6iH5LLsSHAcOUncGTxVb635jsMyaL6
yww7UZBHTOX02p9rtxK45wyR9adeGt0X/UmN8CfRD4SkH+j7wuj5ug65rHcOFIGw
8CkvI1hsH0BAvYHA0GUkUcOEfG9yEJ9AM/wbScFHniTVace2TPOlq0iDCLE2RZ6k
I+lDQSLbZbR3irFZ++gl4t8FCY0RDDfOAHmHJwqWrZXZTdz5QVjMGFTnhTPotqrp
wRJpPcrCkLi1eJgmQqfYRwCSz6h+BN69aIf2s4AQEZfxPFswYXeEaqwaUaQ8MF/H
b/pckdUNY/SHi/ejvg2Mf6Z9drPl3+3CC+2pvprQe477kSvzQJuGsMhZmeVnPvLf
3ofWI0WNDU7Tij0rEB1QDm/WrsFAJ9yq2Tldtdw53Njn40O3a5+ycmig67CZSBio
7CeqVfUwFvpYiK5ttZw78SkgElK0zNZgLTGElu2rUh6lslXZ1qG1SfIQWhWZ9q/1
GP7A+6RdkglWs1kvOkvjTp23875gXDKey4QCnBjCmXu8IOTSUXcBMP073TrFBeQa
7Km2+YK4MNovxb31daYkodtA16mndPlR23j/Gd9e9WhzJNrffCe+Vk+Swjj4PnhW
u9bnpZDKLPihhT44Ry13AFaQQ7LTliU9PUX6E1R6+N150kgL3FFciTg4wEZsNuBU
MAeNgl8ikSRX4JVKbMxqC1t85Cp1Eu8tEFVvl5PhElUHtRPSKVo2y6/bDWZj8PSn
WFVjzioWis3bPGeynm642qWFlEoQU16AHDW9viN13q02TGK6lZ0JVmwhjY4lco58
ubMP+SAfDTn0iZwbARNaSIJp5UojyF4l8WxFp9wWH2JbjQtR2I6IGEtf+y+zlfgw
hbCZ5Oq8VB/rOrp4IwalBWbyn5IuL67GBJzJyWwFqLdShHUNXblotY0esfowJ/6a
o6x2uGdp5hA17IDceAvbMvkq25k+PRxG7pNh/xmC/xy3tpzbc5E5H1egVhR2hLLr
YSc7dyppkouiRGq35grfex+A3Ey2VduVJIYWNwV/pnMv6OXvvGk3dwWGakasBtSB
UR/PIBDqWFZ9fLb85PEhRhrBQRvHSc953exJC1t5kfVFIOmp3R0d65Wxgqp47A8a
tpsfVzpVsBqPpjj5y/ks0XtovFhgdBbbjkr/StbNqyQcKnto1abh1QPFW+PfTTSe
V2+BE31jbTbI4Y6Fz6J5FOoM4XFrIG90kKDqWR0IxvEEioJmA2R/h+Cmq/9iW33Y
SlbD6ndhiR3zaqaZIpXAJf+jks6+4p5GUDJ5FWlty3Cavv6IH2cykQzH5LKgRBY+
Jkn2cP8NwORD//buUaJG01F0Ijr/tEuFCukHXoYApdtDGlVphhuq2zGf+Wnkj+vN
FkrM9KTYu/FM7QQj0eIwa0UrzWgwGGLw1pdvE2G4Grl1xR82NSu6iKGZJa4Azg0/
6KKj6LnMogReQsoDWQ2eAn48YNVBaV6RcPmGzLi6ldXqxWC8sUDtQ1NcP6tWhVc8
ERcZf6ksWdrlLZSt2dWTNSIMsjLmX2s2o5zcTMQ8VFn3RgO1zV/N7aMkuT8rS2wK
yQtYmKr5TcJ6hHr9kGx0uuOLZa0xqxdhNXyx88fWxvB3takz1+XT15AjzZ0lmQAO
o3wzOKWbSBmSZckRmrWvVNbkdHm0Nhjfuj/20urE5Y3T9Da0vcXJrkb18+tTt006
kWKAy8KqRyPoJ1LrAPXpIA+RlcywGXI2EjVGgvvqa+8inHm8aVM2KATtOiDIL4S1
KD1Dqo40QZ7pQJ5u/8eiffsxhm3q404E1xvN9jAsej7i6Q2pfcHuiJ1uILY8Jtdc
aciVodH8HGFIPFAwAPFwqzjEqq4vswnvd0GAvI5mlx4WTgn1RacOENFD6jULidZZ
iceX0zBhP5lqn3Pc4WQpSAaTnXFsjdZAwqLj8YZIcGRypkKbJtTU4TjcrzBL3fgL
niUm9vGCelUbhg3b8NWZV7q9+8YMpeTZKdYicNV7JzefhK+t6Crg3K80wzRoU8Ee
3PgKbtNsLj0SVzmpEC67Yd3k+QS4Aj9pIG1/8uNLBNBxMqi4fQcvJlrNLAP805hi
UMS6PwSYTuZyRmbVPzPSZ0jyzmd6Vg32dWLzfmziu56D1sd3zKG/Iwxkexv8eyeD
9lrczZdD1VTWj/kucQvx+TA0bGRe0ihvC43WpwiOKCI8t3mri28qUtUAXea8Yowb
jbm3PWxrW3rpXMIJIjtus3mfntztn38KAe3og7mDZnIP5h+MBWFUpPEoad8iRpZv
WEjwqjbyQzVFH0VnqlNJ3Uz9cEPACnP1nkXnBfQ5nmlka4eanoRg8WFSQq81pVKi
BWxp3wV8L7y2ryAQ4CPbJYJx0RxjP2W0l1+PodxsrjcwYYoygi2LzwnALYiYBD6I
P8V2d6FoNwwj9rutz8lhreGLzLY4/m9r/QZrifdfpAaKCVxcaWsPqqxdUo0/cCHE
+RT1Gply6GoQuYnB0Wf3U8LoY5von5xMI/jO7o9tc98tu5V9a9IAYlqz8BeABjTj
OaNgqfmdI3FiV7ve0TygEq8wfrJJkunXMZQ16VIA/RT4loMsUCqoipcp8/UdVTYr
zMxhE+Mf2E2MdanMIq9gERuyc19NAVkqAIgkAsclRAoeIsMZaXeMRhILzeFH1GZ0
EDmo3Dlc5r7Smy2QIqU6CdmSP6Xylm6IVcUhhxJ+wYGrPO5Z4NOgmpndmkmWzW/J
ba3id07Tl+AR/VKCvQW6U1dhv+Ba5spcjnoDo3QoZkjQ2bpFY5xOKd+kuyQz2RWP
X5pL7xkeZIjtq1NuyX2vDobLHvR0ZEz7u3YZ1SeQV8nf25TH6Q/2ClUJOt2fjdAi
M8XpOLq4EFHUntCJ4iuAKt9eUkbOW6sKXzDq71VWcZB3qEVAiEeZi7xGojyGhB5c
irjMBrAmFbVL1CBavurFb6GQ7duD7roPZrS7eG7grUPd888rt/sslY4z1O3Wwg+6
ikW7Iyh1E2LaBaqORVHs3ZM2P7itcBqjskIr7rWDowUwUP3g6EOYmWI5FhhLyQJ/
RCiBnWBVG+2hXKV3xOHnOMkl1r8DyIeNoywwzAEjipoJFPogF3zJIR7QdwGmSi6s
/Zy+RXTVcuFBVJ702dcg7AAF9l9Y/2kFMuWDz5ijgn0mr24wsGKH/3PPS8A0Kh6j
e91HP9MgeBXqliJ/gT4mrrpH4IYUgMBJ6NtMe5FdjoMQkFvbj63kh1XzEWJdJ/H3
XgIeKKpYMI6xHC0ZWuG/d/0gDts6X1Jy6IV5M1SwyQVaYOiKaUZZsBnk2jS3g048
T5AJLp2KboKzL92gdhm59Ri48UPnrbvmlsHF+RR5o58d/2Fcl2s5+ogNFiqoXfK3
OfZ1+bM6UW/g3w5q0SIh8XxKwBptM/q3xi4pmN6a1LMXC04e7yPofvNE6+I+C2nX
Nwg2sEAoCNCPObnyw8jLIryjxXnr5gN0ZRy/Qg07xAj86KP04EobE4hFzfJ7yNT4
b9qgQoyRXUdk+i8Qnk9TnohNIjRpCs1geawdg5U0TTuEgz6mCOkmvJ7Um13HhI+j
lxQ4r6mWPtpo3G1x/1Tbebo6u4PrTMhjsqOZhODCvkFsLfVUn09oGhhvgLawRbg5
UEljbhKp7b1YwEgKmb3sQc6bIanspgZDOBzvU2RwtAXzvf8WR+HXVcGBga4L/3ic
897KrT4msUWKHcN/uzgO9yoBIk9/CQjXTPG5gEmkcQJFXSqr71keiytgjN6MR98t
uEIAbuCI/2XT/oNceGUFA/UUWIlHc5WxXSaSkvYhA7J+1WoKLjaFZsKJiipNpdbd
BOr3y5F8CZtA6bhhZ5QopSd2+Ghz0MNn1GNEZaOTyz3/hRsKpmfn8Ku7T50Wv6ED
bMpJz3VnC1ZNHyRLweAvetvaioruQscxnkYVjvFL4EBNcQ5+EhtbKWkOGxMKnT6Z
gozDu95MlPSwpWKKCp+sh6BCahm4P7GTFYq4Vfdvxa4iUAccEQcPa4nWvwgKR64U
533dBuZtJjDA6i94LEVYtFi6qkWuLp6rJJLG2RNK2Rk5VWs9+R9wwVgy9s9dydpC
91vUrjiOr+En194XK7GNXmwWu9keK3zF+/8gpCwnRQCKg8i2Cqh+SDrZIA9o2WiD
Chdcd5XJl1HGaXhmVcagCWU3ACtSZ2afEnMfTu6KlzmwZB3AwrKUDLIDyqJkwOFi
+Kppx13bGRxcYw1P7GhZG9F8fYo+rXQEHw7EBmiUXyCSAgmLJKetEY21GZ9/Oqmr
6XjGepqkgXdmsPCC14S84WAvo+l0nHiug6Wi8f0Py89oxaJSjnhmhSuh/ewWNUE7
lN6waRHyU7NdoI9ePMl88HmFqYhp/hR2eeqcpGFs8O1NcqLyup0Q4EN94O3oAf7S
d8gza6xoAKau7s2iOnwBAlq1NQSUkB9NPhB0WzjkZymDwWFE82W8RHZt0RjKW3VU
554F676pT6TRKMmaise6oOj4KNTsvCU7As/40WSjApXD0a8gENeOkCdKV+uXVAaR
S4oA5ndgFl56hGIh385EgW5BbUtZK/+YwWgONbkxjZjefvD+MZnvKMhsgB6VjmAx
mxhc52IB6EXr43qcGb7npClhl1VohuoIlQYuTXQURdWuDMT0U5/0z8VDM6HRwcgH
ZrXhzn090EwcBUWyJfK8uKkljcFHhN13bhtm86Ad0eumn96yzyYwXBfWfJUtiX2Z
8i6MN4IZEooukQtjVXQnJF1JR73B2eUiE2vMJhBL2TlPKWlzhozI72dUmtGPanQx
i56w1ZjW1TbFgGez3bAXikFr7pjY8g/kJmncfc0zrWXv8PcSsGmdbDo/n78YddLu
4PhMbfauUGed7UCHhlsvdQKA789t3zQ6lVEt2Rtuk5HfGJPRQVRzAdzTKqC8Vpb8
1y4WKItYWhNqgXV8V+3lbXgQzLltRYf48Q6grLgb4MnLi2hA+3edzfSxD/zF5sO7
4/qRHNqfzR9aW6TY86S5ST4WJFJL3bLiMLrMLuGR/l1CxYliTf09xcVKo//6Mowq
wm1R2J6+H08RsZJvqUV6SM4ipQ+YZkNlch+UwrVChGlHkoEQhMj92S645NTxS25j
eoIq/dqK7nqBM7Mvk1FMU5+vJCxk1118eL3ClioDlErIl5y1MzVzXHGITN+60mIn
0F71KrEmbkmEnlKT/jSejSlvz9D7tUL06i1dbWp5C4E96DW2MB8zShghNPvYpzUZ
Wj26co+1XrlnvccD6E4JzxlXAjbCSCxnRZ3ghsfTyrlqKw3FZ72TWdW8EGovQinC
G1hRq/iBXYy9+6XpLc6VSFzIXsgnE9K/fQ+zdF3h5NWgaCIuHn+oxJLk7wEowC7z
9Lf7cOxzi/USVB/6qCasQJJqPJPF8UEzNKxyxQwTpnGRUH5z9Y2RL2PedFEkwFdI
lxEIp0kWLjR5yRSIjoZINvoTYaZ7TejE7XEw+3W693RhhC2rOKUHuqTmW+xpXNDK
4xLPTMWIOGVkLHsOaDbalvcpSi4Sas61fZFDZE5nV5mTJDyAEsE4bGnmI1W3vS1z
SFDC+Ng0dWY4Tyga5bXUnA1qJ7pFECN2SpSm5oChLKD4qhaQaOimdkFHboUKXHsH
3Sl5QgVNgMqLRcPGYhTPXP6lCCgjPTS54hVsW4t96OJhZOqlU2vM0DSHeiwaYKIU
vkA0R2wDLdA3cxpFEZ2AY9sYxpH3I1XXNmMkyYIJ/+VciPPySmBOeWuTW6KQcfw9
s3CtuRZAiD6/6CHNWwDhHee8zzKbEK8fa9PSP0CZ1BOOUkH12GeZ9ov18n+fILCK
x9xd1ar5wsZZIOSIvdk/rehokZCP2IzKqqv97XSomx0BLwzUJQ9SXrQ3R4nTlFQJ
OftbFVsxrfKA8OAC+Q4K+wNzkgW2Goo9ut4LgdrOFse6O4V6kIZo/xhzRCUO/b/5
gMm8+psBdARuG6dwuxHG+Jw1iyvHRooOKJGcTIcvf+wX2Sb9In4BkcQjvyAz9QK1
xLasw15XHgSiqFblek6gGWHVPX2ogiPtYY50U7gjp3yIOlFx2t7Z7hJqBTn2f398
OkDFhIYnF1EkljRa9NoKvimM6psUzcIfC/d614l/lQwN41YSHspZYbflad3IzrtP
9voIJ6Hc2xFewHuVjgN8tf+VNvzBXfeGO2jUy6h+HKtqHnvodJYMfJttcGUeZk2O
P3D9FZ8gf+9cGktEg1V+hgNjpuBLTh6f37UyPF29np01PfcGXqdRJEdmOcGUOZmQ
bMCbIpCSsKMrZadekENnrEItBy99iCAXtratUmiXYQ88tCb+pVX0RqI35ntd2Jyf
coK2BQxk/KyDKkV6e5yPR8v3dvhrqXudFcAN3wvYw/4xkY/BQtPqcA2RfL8w4tw/
BR5eUtB7u3o+Du9ol+VKjyBYHhnHJN8sa3HxtMudrdtrBwzePIDx9/eK2+rtXAJ2
yonZeqAvvpkamcKzQDaVRfUkXwYuHbzuOGnucQt7F0HO4yU1x3zb083KCKWFp8hl
7xcLzJAiXl2o0Q2cYVW7eoPjG07fbcr7hey+xdYpg09+ov5S6gdRUKZAFb/9pBhC
Pi3EXUNMZysilbyFXB8b47qYB8X2syZ5KdBwwN8249Ilycc3OnGHOWQm4nUBMgHl
1tmaYoCvNPP2U5v3KsIlihfoOJ1J1rkAnVMcoSRvz7YF4xvNdxrNR3Gh8Mmn9UaL
2TyYmF7JmQeplWYHt9DjNhCbS4gNvT3wLeHIa62U8w82c2iyTc8kQYgTvVRtGcKM
bq/RbGteMiUps+tWFp3hucGPJRCn0cmwEtz9oJUAiD+faAU7Fo6Sawy7wZdbqjkD
cvv3QHgEzYg4sXTYczsdPi8b1pJk3n9G35FylHdohcNfXisLupFoxNci2iVLy/7R
Zl2xM9Arr9NAwL/czyrgFApEz64iGDM7MAiUs/unmz/LS3zOQk8lsEuTF5GA1V5W
XNWd9aH0yHT7UVRjSI+qkv54I+usQoAFHeQVdgVP6sl3zM21n75hzGftcV6lSSlK
NBiF8ZQEfufNAWwktWX9H+JDkhcqP+StCvlIbJOexHGACXwWgbLXM7dBuf1hQeNC
ZUTE/iAq+xubutzvDs39HG2v5oX523pzprTdK1TG/WvvmclLbrGIK9Nxo9rs5svP
U8SLZtZ97I6cBW0y1L+H7+x/6IWIDcMqufHpHa4U4UYD7kCUt6v8Dk/ETSAMlO5v
Wz9R9Ppw3lVGH8OV4w8IzqycpP24l9WHsNMwlkTlGpY01DJMQWx4CmtL4Zc7UPbi
R087GBt7hjRhZUUoGXNq43/cwBhblnbn1S8wXe490Pnip4iHRGL04GwcZhJNaGRf
Gays0sh4iIHyOjGEnuhmzZDsjIRdjvH3Mb2EMDDAGGDboKKuNSK1UI5Vci0UGJvS
gbN4BonXx4q0qRgznKHEZELkCVQ82FOFKwCfwWyzfg6McH5mrmgggtLEPWSCaSTL
mS+s6aSs7tJsGUuhDwVUFBLEFIdeBthSe9tnp+4ptym6pzPM1IG8fgYKPnnbwQWS
9BxVORfFSEhmXFNmLHOufUSWQaW45lImqfv4EMTnei8rrJuhjQ2S6W7lXRqG/HBU
Rx9XOYe95wLo4IWNhOnTjzrmfwgWEcaIe5In8gGOUvaBk9cIKKPgD2CoyiAz/qqM
9zP1qDC34+GBAnxVkXK5W9iw6zEwdGSdBxSO9GK9t71I13d/8Ilge3ri3H51tAYA
bgRMtSaNT3UsURLPv3gWlrv+MNdRv3M0kQb/dxWqnkPTE+q8N8zOB8qQha3ozys1
QgfTwukJsfyo40K1/dvRLY3x0/dZjYfCZYZl5Um7AA6CuJPYbirX5n6eZshq8mch
wc+hCBbjMHjYl0VEvqluoy+sciKGf+cIzdTpTudiPUDZsICndv7t0VPP6y6U0KJP
YvTtgEloZisa7j2kEl71WBhu/gT6V5VCgrV6vIIiqfrwfiYoveaNeul2w+M0HN34
KdivS5nnwOv0kUPD2tbg5YPKjgBennYvyeAJTQs7/8d1RIFx6lyWIEh3oeNrePBY
MtstHDGmYtWogFf43mqL/j5j/I07wn9bpAUdTN1Fj8OfBngAf/i3PeZBoCOe4nXb
65EBWzXLQ2w6A/tb6O8XLdApcJdpdhSHWye3RGoyepNVVnJFxKTLsTy04R3167f1
V27YF5dG/1nImtUGZtgiF8ODlAlYE/xPNSIthzz+2Ar3pkqKp0Pa7Tow5BiPADPd
FzC4W03qU+xwQcMVSOf/EbQAht1+Is+wg22x9WEsiWkwyuV5WkyeGiNoqF3832UX
b5Qhw3vUjUYLI+RD3o6Sq0NIqiMnb4fT8sGyDmV8ARzFIIMKBk15YVn7ws4wBJgq
JMthZiZq7YOE7drlTbRoLYLw7g1CTyKYQ28AG5oVZX6NRUSQ8SzY3K58LjAFJo2a
bap5hnavzuJcEWLbrstA2GxTnDDAGoVj+oQy2wPmbtT07tsMUh2YLxojDFbTT6Hw
9TIJSED6MtLX8bR1kjSvly/kkVdNNZcBph3NQLWY1VuUej0qSoEvVrZZ1EypW0lH
GgSbdfKCNGEEnmM0GRUrnLA22KjJhWQRyMBpcMfbiqGp2HKlu9upSdP6TJMF1lje
/5vYOkcFNg7OWaTHGcC1wzavRejwID2S2rOQkLVjES9630fQgf9p+4ly1c8KnMxf
erhFpFUIJUVg5NyRLE+9HFnafG6jI2Z/+18Byis7aHe1sLmMFAHLjU7qMA7+Y/fd
ovJButxvVSHGo1+Rvs1t6JDZUdCNiqhPuvltNfOVhPTJuu2ftQCg/CwrrrZ3fhjd
XPZIAbUH9QVnGR+CwgZICQaROU5mxNLgMd/RvhQrG5Brk+TUVP7AJrgRDY5UXq91
bPp5RyabxL/Jp8X/p9/D66CyRYqGp3nQVG/Y5jpmqkIs7NFbr2g8x50EPDlmu82r
ERgJE/Puqj7zuAgJZRvlJkSKwvnCfnelMfxsz1sLp6xjjd5jOdN4Q22w0bMM4oqu
EmdbV8+MUzg+N2uoeXU2aNQqxDMue1sB1sQZOJ80OIDMKtAqBHcmEbqJiP08BO5+
lyahdn9NFK7maLDaeNXHcm2c3D8ZMpbPRgn4iTWAS0Hoia7+A4OxhjozPpq8PNE/
ZD+cDKqHLEEADy8ua5UqxLUS2T0r/MAEZaSKtrkHAQmOwoA48TiIbH/Ow5bIEHCP
93PRA+eR+D4hrWdsucCfUNhUAvyMCVm6gaOrRH1sO9KHE3TIDVIIYiIEOdxceVg7
A64/wUmqQACvJmzwMr1xzHSve2wvxF55ZGbQjYgLPVC0N0OGr5WQajZL/lHPPR52
j7nq9K/wtS+U1rYXzdt9bKUDkXjyyrUtR5UviTMBq56AE8zbgD1mh8egzYzkfS3R
xOQHyK+wiFHGnsXy2LF9llfpKrOSAUPOgCHr7paDnfi86T6r+9NXR2octgZv8zbO
I6/bVF6mDYfY4Oet4kfKAnehRUkV99C2Ws62mz54XejxYjlNycJksjPloBIPKT3s
fezqv1oRapcP9kPJsSCMXnvyiY6R5p/w7zmL7096Q4VbtrwT39dYB4DU5z5zdbVM
6udhd+sifOftyDNvJ2DmxeIRF/nfk2DZ4O0JIQeoZURo06VxCesdwtYuATqLCQio
5W2z+5quW+WoP9M05L9oVgzeRfNeH1zZ8jNLDk81hS1etQW/8R5pUNfMahen/NJp
spkJvhaIW01ZOh5cSyaAByW7I9yGwIVNs1GERqM7etIUbNAZomOnxGIVIR8JzuUw
tXLlzAnSAlD08Rc5kmWT0uFk+4oL/my6aMS//TmYwddVv4NS0zYqL1JWGlgUEyQO
YfGvWVj6fc98/peaEe9Xr8JQjIig8RlmShuBFcS9h/KD6Aq0RmfYSK686sHbsoGO
KVEH6MoFt6EX9jj8MmCr6HxooSFnotSaD7N3wO2fv1KXxlkhlxfe92pXj5jLxYM4
RL9FzfseGXZu3WDtEte5b17DpPu0ockcGeApwAyJ6WMQ39atmh10RRp91D0FB3pP
Ak7bOJMrd7cxX2/XWlkvEM6PgMcD0zlnYz1dSBtpOCbhfno8lReJ3f/zF6poOo2F
qtdtqFiNCJyT/ZJejGQl2njLarWWxFNoPxy7KeR1SaXm0ZoAqOsDbLdhzA1racuA
Iw6jjOh8B5tJE+uN253umkoUlu47T+TITtzcV0JSmspdr+v7McnUBhEOW3laRXXj
ZKrGZujYF+N/d82OdFsj9szyoFw9I29nGNPZMa8MYS1wbnivorEhh2J/Sv7hnm8g
S6VvEja+zNHSjQCNJXLfZQzw1ZyVOODJG8iUc0THZEXgG5+AFz6w9buaiV+XbA+z
Y2KM55m+bFpt450acPTalNubIyka5/FGC12btUYFlZnUhLTawYmvzs++usiv0CLC
7MRjI0hRsBb1pNs4N5R+Q5X+875I23TPOrAcMvIDFlIuFRc0yNLjar6PKaSd152r
GMi8nmF3m3+sp9Sephee08+DR/puNfEOLNirz5ElvBflLu2NImtCAcLQW2p3RWGf
gmJ31UNax09sIqT90HX1bnyYNkSuy5WWbicR2TshQMICoCk6Enil7kp7749Q5gP/
a5a17SSZPRIAFf9bGpEfJK8sM+kVx7kAnPaqWCkS0mCCgAFoYPRzJvwH2T3EF1Ih
0vlgHZdJ1KIbFWkeomvTLZbHH1niGgcT7l/II/n7DzukBucWTIgUL6xi0NWN+8Mh
1P5vmxUIyCToIKkSrbyxnj+s0kbZzYVCh1/XgLiENf4GEDfO6vuVt9DoOh6xd6IW
Ww01Mv7XwcpueNzm07a+KyK/+8VoQAUv0vDhjrGiymwhMGlHczky3VBr+DrDBBCU
qJzMiGDpVJgniUEDTE1dn+XNUcMNeA2jc5ckzb6+bmzDpFWFAWu9HwvpQWFCB73O
4yieisB/Sg3XmkRpatBkGsCqYHKqYL5fC3faF56Y6sCeY8K3EzdkJuadIEwXaUyi
M1S/WdlXV4veGtpM5MXITciBbfm6VJeNRAoF+aONVnDyOUPmXhn9dMmkk53rT3XP
RolkL0V0q5ODQX6MBmRek96Sa//aHIMdHVGiVfQB8EYXItQVy23zjg80DFgELpsb
HZQPqqL5cRMbg9RvcJG0TzZvwtccpNm8RNFfrjJhiXzOKLzoWBsIIvC3mVAJ6vEl
bxGXFphOV0xbewNxoesGtp4yqEj39yH6He/KqWC5HrmjsYMbRHP1D/H46EYrm56j
M+CJoHzkMYS16py8QNKzWVKfsWww2nxypmRcX0vHXbnbiyQrUeAbwu8SNkOgc8FZ
DFMmga7+TTyLZCDm7D/HBKi5PWLyK+oEngb1gmfwhBX4twxQoqlEePPnjkWpn/Pc
pppWWcms4ERNEJWBNlRgH8UuJxXzmxj5ZNgLvXcxdHCBJ45RIxY3kX3MGPiBc16a
shsUgb8MOgNzfPrvUDvvhL7ViqALosOpyvxwvd/PhXH+VNgGF+I9d2uo3HrrQ5KM
3tarXCB3vZghYZ2yd14jXkrB8JYQmArlSMLoiqz6yAKtyRyaF7yJryYxkIiNSC3A
a/opr1tGy2AH6YqlMo/LXotA62Jmsa9ZgaytspBCLotyRiMC4tNm31nJwtL0x/us
nObVf8ZLSuitS7u2qJ5IN9LTVIzejsmNtE1T6qEn4TIG3FdfEZu8Z26IzV19rKaD
CaK8JCBHfymHk5zdCr9VvSyqIgAhlWhw9FwX3mOS6KYIz/D0+m2v8mQ97GjXG84r
F54PqUyNeLvcq2tkO6jEtQHSHgXUh4pQQHXWbMabNtR91vMlQiuvCPU3THbiCfP9
8n1TjmkI2l4qglV6eZl97FR0d3+BRrgZSRMwYd6ZY61h3/9sWaPC44bVNVjAR3mB
1jb0gizgA0YPb8ECqSLjK1HSsYVLsg2P65p48prax2jhq2Ist2HVXLq5TkKZL/qg
U5dVVD+86wBjk7ePA4jd+3CpinS/+Yp5swFLsJE/7ZAvGzns2romNjnbX5SX+xGG
78S7Q8U5XZMpfBnuy3pc82T6WcKkj6/4jZQFUyw5/azffhSIizz8LvwKj0ozIjVW
xO7NtO5rlxUdCLd2b4kWUUs/4SDIuyu5oJise6r4wMvph/SACGOPJsto6gJQHCLr
bcowBJ3m0eHi2txhsFb9+NVxffEBa7lc/l+5TLxLP981B+tHJQzXsE/GpQevhuF5
anBe+j57+E9nsMua2Yswavoaf7XSdgVIcF4LkUPXOf+0+O81uBW3MWiiXGcwiX/K
kaXsnQS3HQhkqlqRi5ecLE9PZZXpzkSAVoWTcCAz2vlQ2rjNuhldf29+18ScSwqh
WuowK/zWgu1DaleBoBOlOKy3ZKbMKrF6EFqk5Xu1+FcTxye02z5x20Dj0zsloZgv
G9FKMJFLPR9XgboRER3mbv/7T2c5BUW/E5pt8CaLj5cc6sakIbAHOd6smVgQKDrK
UWScKaezQrN1Z5Ohk74my/EmxB8tRaAB6WZG9VsD1akJtZuxu8dW4qPYfh4UHXHN
CaOWizbcPIYdpPQ7H9Ce99FzBUAZjrWeik+i6U1Oa1KgLim4Yv2+EN+zoA7WkCBn
CnrrAyVVnj2/DqJey1eeePb7vlhmGjW11nVzdhXfzQH6r+c2bQgbry1BPCWkNL60
DFF9AZM23PmKYF3wh2wbEpwOQ9r6CartHuyiuxoK6uNzWnS+AvXqY/J4UEaxWXk9
jyAnVoVYoazpOnr24G9XP/jOajWx+QAO+SbB2Pd4oqb6MPlA5xZBEgvte3thqLQ5
N1gp1RwhcboA0rN3yGTrtrSpFonY8YPLbZlNKyT0qh/Vjujxtdny9+efXVRcQZcd
pEZfp+T084DI3MV9NTlmSaMRLtSPZacDDx3+Jc1+Ba1ZiqJgEOwvP64Cjz0IEmo9
uVVZBo7IeR+lNlRsxBZedJyVlVkSK9py7RRyXD2p4BaxsT4+RDXk23R8F87Pf9Zm
oOuZR3cs/FNsW6Z9vlhtU1jRcyvR008YNhO1PzTtSKS0h+dBQcMaHQBfJYmmUCk6
sGc9G7O9kJhKAolruLNKHfoT26AxmdrEfYtF8VhlBPU05XPgaP7vFfa5mvvYSskX
xTdwYC12JnHx3dTJDoTOsSsN+YdeNKGYWrgQJ/dGAEcPFV7fEF6AVxX0cai1t6B1
82+BbXYH44y7cTR0Vo8WCtC23E7wnoytsQJLI68xVPBVu2ag1Ts2ekhkWgMPy5yC
MJXWxJoaT4a3PU0OKHS1G3fgp454BzyOtQ5WeEKu1HN5T19sAKLsGIYf1YPY3vK8
quT+882AKi+iHjKyrWRsVnec2MgcwJPotsf+/76wvMWXXEBsnaa0/dDitpllPXU6
KRAXiex5e8pXTZMZDYeZd/406axrROK8cqDh/b4ihN3bgQF8oSz7bH0sU+pHsdHG
+psiKWOWJ8wkJNELgNqAkLVKCD0hkjRpRLxhH26mDHtuRto4iHLHUTFMUobN1CS7
oQ5Ts1ILGv3ukybMDBLs++bHg6+gasuxC8sKZf2hHFS/wklJr5UhpW6MgAoHlzpj
cBKEfQP8ljjt3TZxwl8H7nZXdromUlMDO5jnbnvDGhco8FoAl8TS9qM3cMJIF9+w
2FtcyOzoezi7HPiyK/LTvwDVqmCoQVk4xooiN/ZzuricADXoUpPnhg4ovk44eOSH
g6uJA1Y7uxOTw84Zo1t5IFg1QfjCdh8/Lboyv1pFh0A1goVkCl8VgWp++z6CfE6g
oqDKTQ0eDeEOxUh+mwRh1lNgws1qIVXwRcksgZSDGt4gOIIcKouJ+B/b0ojObRmi
IXhsc5qQlRW56e4/T6GoeL+2WEJy9IFZ3pnbTrNebKcrwoyfpIyel9RW9sVO34jV
C3EG21aFDXH7ENRVdOgVCZjvPNMuWmBgmiecmiG04SSP7jyWLmG5U4GAq47ah3Ni
Q+gjNsQovdaH2Wil/n0i1fhLHoncR1VAnYjw3reOz/qYajS/srVOSst5fAJ2cK2b
rtLtTmtjNEvt2udYNuoyIfW3C8Yt9nHpJQ0Bug/I/wQ/xaXSbB4fc9Kyec+SRU7t
ScTP2kFRtf4H5yrl/TdgBUKRO4qVoGIe6RysuV28xtQUdT8Vn0W4TGihoNUxIexB
WQEaSu+IteaWjG8T8dnSvM+jqFzWyvV6D++kGCXhZGjBiSsOHZyc2j6dqgrLWUTa
p4o6t/ZtKvHOjauuBFHnnkqBAdFXUgvRghzScYhvAxrt66BKTtcfGuMtyuECdcPG
xZfsewIfuWaxBb6KquGcIphCRw1NAFj5Sv20+cE+4gQz5kgoHI53B/won+NQ28Xt
FmrL21XoFFvIGjI+YfGqKctGqhs1hWZxsh1mBWFsvtn/QHhvO4Y4FVzKejdmKnnm
jmWjNlLi6aL643gQCyLVeuPzacWrptwPeoVep8ryr1WZS3ZFf8FMGq8Mg8HpOHfm
gSB3XMckrjZPSmpxeOMg3A37fWVOQxnr2unn2CvsIuwiQat0dP7EQ97dkhmZ1ScW
74yNqJ63kmjVtJLBOMlX1vGoqGXbyGcKlmgi57Q2Mmiq33dqxvoVWBx7Q9txYAmx
GovehdYp0FEqrxKNPT8BFoltvS3Tqdf0GiGQkaaUbgxp4IfxW0T3lbBiVCan4qKr
JbYy7iSgObD3SkZIvS9ZBFbWLEHhD2b7BsjQZC0LF9+2/EE3CK/bZSzhaE4qo/u1
QW8EMlY1JYKkvH2HHXUmUYMt2yyWzzZ95VydMvfGtB7hiJnJx+RAOiYLraABuHuy
cGa4t6ApAO5XVjDRZr64tdtnXUzpuUDkgYFlJ3ACczJcAAVEwZhCuqwwl5XHdq8v
exauAbu0QssapOqAUODry9dSl3xgi9CD+sb0CdHHXb7lxE827ujae+DxMP0H+rnM
su+KKg6iVoVTNn5uCrK6+zk+NqjK+9m9QOAcZW1bz7HJb4iYmnqSWBMoqU5B5AF2
O4Cj7lz45JbfDWkY9hHb8cHTcfniguO4s9Xod7BDVobsenGVqKc91lXNTz0RrQL1
XpoBQ1XMjyO/9WWeDdkl+v1BKktWQSnr3q0D/lHBPcHF7cA5KXhrHrp+c0JicfRc
zT2X+gSIMOMss01Yp6e3it7yrZ/wOV2wZsvbzoPTqEsh+6ye630JG96ty1fvvVfs
4U/t1ZMtVny7nmF8hTX2uMw5vcDtiv2vkeYAAdzABgGJ7R9BSnxsGEAmu7937Ia6
5oxFgxIED1P0x8Qet1aMSz+YjT8TT0lwEFTKT6E5pCxR4g4BB1ywerf49skUEblO
m9gsisaxH8L7BbQYjmXOF/c18idrNk9mx3JbkcsNJ+6wvMswkvSX/EN/NaRTaVVg
MBPezMXsSxQo5S1xWyg8IS6xr6kPgeLBnXb+yUzOF4hlCVjZa5So37zmr8ed7/Sp
FORw/N7FddpvsZikc00SpCmROW/bXlR5HU9pn/MtXDCrlNKaoGCXwu6g2sZ8uvbM
ofKvNUTE/B6w+vqrZL7F2K/Xew+/xLi9gzm86CNNRY7WFSq5iMGi5MJYPp7b8q7Q
9DEvopr/OVIPEWrV35BfPmZQL7fK0GQC+UX+0EnvnU7eRf1653yRDlt96e8IJbfq
KQLzWoX9xnZr6Qg+mLw8waI1frv3VmLp7IFsvzhi/i5DYi5vAUe0rtf/0CQhWe0P
m+2uoR83SoT8MsIvdED4scfEskwvI0o7ndQx5EZVCkfOa56Ojqr1X3xwWF0P6juh
r6dlEo/WrZxVbMx24hu3Hxp375PfIOfTahXqWILqp8yNZRxO+ykRQ/nTwBZd/7GW
LhfO2K0urUNDmr58WIs3K1FFdGeEqhVzvSGIVLtVV7jECK8+DCnqBUVxiXctifCK
npPfSeKHG22QqPbbz0nlqc/DBeTyL83CPh2YRzcgHVmsZs0jshbya1p26WAH4Kkb
4U8lMWs+C9YI482webYfEmDSlANT957pyW3OOJbfKdRMxmjHAwqad0XjP+XgBLhL
UP8MzIxxQAsHBYyLgi687+owh4LfLeJNapfbKnVbX3vs6ClKRjLCMR4EiNRfhgpL
0NzSsbJfcfeQE8wIOKdX/KMNPL+IkQkITaUNYmywpXpTskyn5ivpAd/6FsDph6pK
2uMWJupld92UTwTXuCL9rmT2JamW3eBq9jFVqQTqhQ5kHMFjO9pxIvADuTIA/cTW
m40Eb+mDblPZ0Pyplnqdv8o94UEqfVxqIsuyRCXWm+VElKGiddgPB9AgoXkllml0
MgmmSkBGxghB7kXhJjxC6h59C6jH2KYtimB9V4Kl5miBaTi6PewVHdolr4+FibYp
/WOjyNQAQ6L8CX2s9/gkcUlvdiH7iU5EoHBOIP71rb7HDyuBQ8KIPSWCETnyAXf7
RjL1/CDlBmf7Fdy7lmf4i6DJdwnsDIhFJOrTkV7MWE0/0Umb12JJZyIXABDj2o9M
pFvti2a04HCdU0ITOTp/ezRYmwwp8SPMzfvFgOiilkeeQpGQM80xqT8huGlWzNmv
F6FJ0uzGdm0Kn7MB2pJ+fD0YygKhs6QD16rg0+AOkicdtLJ1qkblH8t1EekdYYwz
Cou1CchH295hrBM4tTCwq2DCra1Cn16Gil5EP0B6LyWhQofZXLdulf1yGwncp80k
Tfz8GMDO14Ca5tWnG2OGUHL+rpW+VtMTUbn24J6zH7VrIAN5PGXsPIhK8uj5vWlF
jdFHaZsHTO+/jeZGRavJaLfyimsi8ze0Ao7sJvPNlj3x2M9M1ol4w6mP0G8VIdp5
wIZHKfDQ0SNyDYx78EWx75ugN3QCtZ4KairMIluAVMCt51bj2BxScyj6bRtSbzaV
hPQJC7yrr+hJ1ABWwfUwDz+uVaunbv8beqmxWX5EUmyELkVLUmQ5qtuDSj6NSZxC
FTcos28Ye01uNG1i6bMzhaMKf9SXOzeL/oRR6cihDzFB+WbLh3OB+RHnBIm5KfYR
j6oscjbPoJJ8AMF3w60NFS7BTO5fIb2SQ2qghWHpzL1/ZgbovAX4l5HmWEnFSRAZ
vbRcA7be3xH9gdlXuEirUA4+Z1cSMh4OYEtBfr0llK/ofmjjJY1lbbHlSye9tKj4
ZHOID+I+TaMACFBj2NXPWyJqqvQbkYAybIxRCFCwFuhXKxRlvKV1tO6eMUfXZPxO
6sr0RIhDVLHiOsWs5XhNHvP8mlAehAs+N5LaWU5g3fuHBQM1Zh/Bv9JTPZT7ZrYR
2wiTAP2f2Wi3RdVMIs+/UxLGZCfq0fd4m6KvQKIAnRGSoqoqsqSDb+1CdnrOKePA
/FCf7GpbxTQUbNu57vA50gl0Xf5x3ZO0gZIztdYATE3XFD5xM/I6LgiATjmVsrqg
oUWUVUnFs9/l5k6zR2xj50ObXuMtE3vmUhUzBjd7VJfmijv+Jb9WVV53560CWzuA
r1nVL1Iz8VsFUcsfw6u4mGI5GzqnqkdMwaEomBCUWrlN4kzcOvGUySR7UJ4lMKiL
X6bPtrFu/KWkrHFaY41q7M8/kkxPHbWqHlQilwGWbB0k6onyN2zDDoOIjWtjtKVn
AcWQr1p+dtovflSy+U4wRO71cNLD6Y6OyFSdBJGNHjTFQ9WhiWjX7pwNU0RQ8tys
wGPX0Vl2/gHUlCaImQ1bMH8heR0b7K80Nk1sE1C7S+03ETPw9zoV9tsj26/819hv
bosLzn3It9nvwUbY0u6p7CZhxoFlOHAv5ZnfZh4ixY/cI2p+jcd3sHk90sa7+Xpg
n4royJ0lodZkNt2xLjqZsoT04IaO47Jv4ay9+d8jpfWvbw5McI4JB0oCo08rugB1
msi3aHilyAcQmZuXVELkoYAq/vF2/8pBgqwfvOOqXFK1XEcmxKnyXgTT1JLVK2o/
IbL3G51ZILsWhKjlFZjWo4+sYZLiA7QNiYCJz61NwJKZnJjDT7cKSjLGqJeCsFdo
k1yYu48r1KrDdgVxxUSFnTpBC6c4zTiXi2ITSS0L5kb5f8yAfYcnOy+AdJzoiUwR
Q02gKe9jCMEbtb7eENCFFb8m7cUsLTGsztS0PURdIx7pCXS1W/26Vme/tLa/qZBO
Rf6ZJPUj5BO71KchWKt15B9oGOcVFqglCkWQDFBLkWvCTFjezm2WqjDJMenJ238v
YlHCveUpdWtJhsH8TFz23cbngQHgFigZGAbx8LbPF51jA+MH9DvkGnmy4LhzBolU
/l7RLJyPo4wgbPgFB2IB0n3OaPH+sKMJNSMCUoS7QqWR6IozV/ZbKh7ImTTQ0zxr
psS8Qch9OGwnCXPl2drxiSdM/FeuoIGXX1hc8LDpzcIpSDSK/4NM4d/3xyeeGAh3
UqTZGod+MYQcnd8c1sF/ZjxAEFKjfeSLVDqVAWlIq32mBJGGp9XzYkIYo5KVB0d2
I2YNpwxldJsgCYmCIPkNBmhtgyhUUzzfhwna5gdSTPRsKKm9sXtwjDXGSct86Nua
BEG9VBHjlPSrKuN0IezI3Q6JHd1wLJvgV1TY7bgG8yRx3wVyCwVkGZNTUSuMNUp5
fnBou6vnAWuxkDFGeTUrWS9T2plMBjb8AJLs3d8QStdeHf/xdSmR5F6GialF2uTU
6PfpvbEVB/2me8tU5Uj0UPB9LPc/ODZ7jdtp06FUP9LBchy2tMQtD/CHRQvIT9hU
Ep6cj4hFZAN7tslHfHqyoabw4bPJiAnw9pdiGL/dxW0ya/ekbYhfug7DAtzt5LZ4
/y4L1gkGENNO1A+y+v0PC9aM647UkWPLiaEKNHU2XipfwspdbeD3nnjfEjJtwUJg
7ElkHkUT8PIVAVQ823N4zWvrrRdrW+yht+kFAyapfzWXQX4LTZrFsXRK+hmwcvAV
//poB+gctagzo8yrCVjoEPRFp4hIIPNEatJlKoIJyshxWSvDEmJj6j3x2EWA02+6
1Dr+vkHK7fYffPh/FvEmTQzt71qDtwyRMW9FHa7EaSE2MrQq9rl/U/9SnFLbe/Pf
oosPLPz/W5gz94GUZ/RA2DTYQBuRMdmU8VoVnY8krkV67sIGwvEBWYWcR1VsimYC
HaJmtMTuIrhzJdravzoiANS6Hoczh9vZ66G1b1WWjYWsuCAojKSLbhF16iP7nzIF
Mq+RIpXb13Wbx9AXW6lKoc3nATxKECIviNGc5t2OfKvF9tXRtbUOmHiCLjYQAt3Q
tzzg4RhEVhmDiZGom+1Cv8nc+YK6El8jNvuz8RoXRErJpEIxsai4u9lFQT6i4MUB
5/zgqRyewoVJIwZJqRNYU+UWgUx8OgH/E3GY2FdeJeZj/GYRWzfgssyfZy5pw+BZ
mNW1DZE6ErAW5oPIWk360CA3DFQ0PB80HHEzhbVgxCzF1RA4nBgg2zZ+KsmcCoA4
w+CxlZQrbS5GsNdjYLz/Lneb+lVQHTVi+zFkHzKCgQhZZhzg6dTzWqTxTVBawjQ8
CfzLkwebxN71PXYpttTQWVHDzbJH43eqt3rv2aut8Y9GIQk+npCLBHv0tXci2Fd1
1TtJyqedgE6ARGoZ7/WQo9lQ5twGlbSKKeYMaUYGHIxuJmwd95zkjPXmDHoiLldd
k7/8MZw1CF9qb4Tww/Z8Oz3gone33bXXPdaKuCHrGmriV5r8jVq6AWij9oaFcvr8
Ye1DQz54WcEprhDDs/zpov3NL/0gyZqU+7x2EBw12s732voKzGSLQfq9uam5NoW+
2goVG5XoYLtTcihnjB0m6A2xpcKkSAI/XxqOozR5NfAal9XPKW8GZHdpGZAyAsxv
IbXxN7zI8TGcvB3lim74QKTFbdFrVLYoFeM7msekWNzuypNnDGl6uL0PbUbis7jc
XyvFbPHYX/P+tHEgWP7s5WDEnBHO1+pvZWPjG1xsIWMQI464nko5G+2tBYmMlJAq
p2BIYrpOgRK3rPKE73J4vyMGVsIjfLumEdU04ZLvryuhNFZObYLg5xBRzbg/I3Kb
Boobp60Mi/b0T6QkXhToryBDwrvrDPmoP6hXdKKHZzVtUdooHgtyUKYzBswlj6kA
fyEEMl7MxPcTJlAUstLwuODzEIwFhsnRvbLuPfVCd1vIdAXpe7LXLor5Yh6JEjof
vz8ATHcxkun9yWGNN6gzijRvUwml2sA9Ayl5WLwnrleXqDgKahuS65DXNcZFAyMA
6Z+6DsTZJ/yhAiX1WzzF1cKWL9kvEeUpw2O/+5Z3xeF3wWuIvG6bRJQfjRS6Ig5w
8jSaighjH1K8DsUyLag7cO0cpUhtaVyWeGV4OH56UWI+DmgT83Maw3zUOIrqxrYw
7OQS0fO212s4ULe1JYrfizD0o0dkmYZrfWZ62PnuiC22BHPRigCCwWAUavFhBRuT
7yZmUlGK7QFeVLnsjrly939vkMWtYENfdZoxjn2KlbCA3RfoGmHUs/Im/jNtF4hP
XTE6Yhp5onUIO6wotJ/P0jSK99Tbec3mnghDaCt1uaRXCHUSi0MHq1AQGx6zPDCY
XXRcP6hWD2K2fjxEGdD477ut3uazfO8VmTgpahFQ25EWnS8zmHoW4sgiQLkpiQzQ
OXFKd60hfzhIcSvhGNpBW/29poVEpKuBGT+YnL1rYlQjwuKdQTqocdEjMvcaqGed
2XDlEIuDNcET+vyTWw/bCY7K+R0VW8uNW6T0LEkC1BdQKkdImD58M8EUL9FtzACo
GhduCvtRRPw4/cfhQDLXCsTSyOtI5/GBDEU5PmmpITeY1uNrOOGmISbkGOVMsVHj
XBqiAbWgQ4XIm57Mg1J4mV1KZfzBZXw/I/950cIbkxqMEu288krxv27G5ZPf5pYC
cKcRe/d1sF9kr9+xDpJ6JqNhRbjUeoDcScH2F4OXnDRXglCUR5zCmxjtdB+zZYKn
r7Sz2FZQIGBI54hlpBufUq23J0bT8kRUyfju2Katp9LfBsVxCwxoM62GHIGaTX6n
MD1wBeChZpLSfKM8ast7nNrTXu8FJ7ODnzgXG/eWbrWECd14vQJuCas47e1UVwZF
bMiw/vhIrhAU9GModhrS8hYFowK7Sbj9DTjobsWyFMxZW9drvk19R9mZXuqJl2mw
NqBQX9uMB8FRx9zpG2k7nv2XU0Cq/5ae1LQ6Vu2dZ6f+JYqFEkHRDpkXv51igpI2
UfBLkDTSuX9GNoSvsS2PHJ7CRl26OCUEqfckt9ZsK+51UDaUTKuw0NLU0YMWizYn
eGTJ4e8J4PG2LkBDoMZ+DoKvrROh+WdUCGrzeZHBS+jotxwtuv2u49FPAM0Vg+Yq
ej6YrA09dV4O/RnD/cXSEpPf5cfGwaaQicrKlkLOeDYmq04caIHyK74QJUPvtJVE
yy/9/pDEAz8FUspqHVnDuD1tY/e+46pW0s3hPAFS3/RyllstuWMP8mLg6N7aKUyH
oTHuTz9uKZidnnvRRlJyPQda10cLllZFvPzTsPzXjssl7LPaHS57GCUcQzoMO1iQ
CLP2SknXeNHl2hPJEMifBVFAXKhzonMxrDY/NVJdArQ/Dofw2qgaUUsOiubT0WYB
iwGqvSJiGk3uIrKyOnV0IfRonhNZYGUQVn1ja/nUxCElU0mgwKbPP7RpkfkvMvVV
C0tXBT4KpqaQ/Uy+IUmrVG0Cs2H07oMBFUysXhX0sWqhpd9vgZ1d1RUnNWh3/jaZ
JaBD4hfiWF6bsL15P3zFjs+CWDwyX7Chl3qzNlGOIqU0VS0TtTiTR+KN7nccJmHQ
oeDGO86HGfrWS9V3j4zmnLMUtYPguJzTBkWaBc8eOx9mtuDbnhVuncuuHccqXw67
t8XIzX84sKgVtOsoCc19QixoIBS8TetjGdFkR01Wk5BhUnauIgQ6a8dNhVoiKC81
DFUpZ+j8U9smikn01v3dY6BTm7nIJ0xbB/XzU7oI81N3FU1zafx2iDPt4YKUTr2M
3JHa6aLvz6XfD+CuySlt6kFcEFNTNJinEwEImr60R356A0TNya1gnuDKt2damSeG
lAzdDNFU0ATDK/DV+k4RRgq5XTUTbo2QT2myTrKN1hHcqUo70z/Ps3OlmVCAcJmp
Tip9LMMnRVw9Hc/meTXst5zA4STiazHFrjNYQZhzYHYYN/0F4NCMPbBA7ZLxx9nn
ImMuuvwP6FDF/Mp/MaaKrje3YxAG2kh35cHDTHT31ITuj4Oyrwb4FvAYNybP9EUj
0XGgAeKDa5klpe9K9yvampcK/zrn5c1HpUtoPuBWhQm+Wmu+KEzzxBVyCtDg2zqc
ENDqDH2xqrKT3/IzSZoZPCc/78wo6ZFuH3dwssaNP+PT1/RMyFQejk+SsdVBjw83
Cq+Mq5MWvNe6FyK9V9oEQgId5ks5L7aKBEmw/5c/nxenAiWoMcMP7faprU7boJJp
anmxp3VkI1xmmRbzjjW4A7GqfhTtIdoxDhMfa+X5+rAtE5NUlS8IKGGbvZp/vXkZ
GCoLGqTeSVVXe64Er39b7vkCJn+1aCCcNytx62ubddPNVEH6HU6hGRFaK1+mQaI/
7Bm9Qcs5IP/3nU55wG914h/LigHXv+kYrg3sj8VkIWgf24KhCGjE8OtCS2JFX4Ow
r7u41/umx333VYKwEWx3AXzhY/0MSQzGWrdcWFcPw0zNrO39SbsXYFc325wriYJe
I3JR4EgmuTStae+/0z4b4AE/67UX6GvYNfCo2lG0xNWhPrZyeawt/acUAR8+bpI3
weeTQ5UD7yxPVCb5U9t6VZih+otD4UiYNbwDN7l4qGWF0jMBXnO5qrXsrzbJI5ZC
5HGuw1VQsflnKHWbD8PyxR3BKrYlPFPSXX6FqcLeLIOBiUDpE8uuwu6MGcQ8dNHI
i7N+xv3RaFiCxdV169RA88acKV7WB2NFBlq7vEedIVLJh/oi43o9+Z+Vg36igrQL
YamlJXMecxVB1GoIMEqCo+FGBuC1KwvRQZpYZe+E/auW1IcmsT/C/4yLHGbfzblJ
jy58KT2ysxdnBoYePHPIm9JoUYBI15ZsdQBw42lx10iYqGSW8L2eobaVR++bYq7q
z+Eepam/56xYAu3wA1cVa1w9QC5kjJnjnkGSch2ABrCVfxvvkjol/sl1S0vKWsF1
7QWtcD9/toneyojXGvXS6HEyqumtxPhVu0A7Fp1nVXPd3y9yyWwM2+34w7csB1SW
3wTIcpqibdcPJZ5BYyb4byk2PpT/prpYmEKl2C5LvyDatLd85S4THoqau1NjT8r6
CgO6xIel6JX/x2IWWeWPhN58Rqd5eTeYXPgdgcC3xuZv8LtS8b9PfUfAkzOg+SW5
e1T+HRJoBrQO0Fd/8CGJs1Wqq/WrOQ6KoY/Xl0DIw1QkbB5Mqs59oJqnq9SdvvtU
uk46ZlMAEJiNkQjiTGFZUD1BYRBWnpJZQe/RtzweNEpwJ3pM5Puj1x5wYCEHStwx
BBY8bzn0TcOKvZC4qi1iYugBBNWjhYZw8AFfqOtrRl3mgKsIHZZTH/iXC8HeXGO2
Lnh60ym+6hWPR0y+5o0cfcI4NRtMThxTKd1CwEt7Fl1jSVVnHpO0PdX9SgmOSf7z
4xIFCuf+OP96519vjphl2tRKESXIbIWfhd2k6xzmkaz3/iSGnmMD1Q5am3uvBlR1
Ig7DGvM/MhMrpywIeoX+NRoM+LplShqiZ5BkFmgP5zQNkWwB5fNS4iXrjM/uvVT3
WUJYOVuTl9SoqZ1ykUwzP7oIhcnig1zwvFyuiRyfgqsHPMRqGcYqNbDlPyPcQos4
Y6L80sjxiF4qOPZCaZWumz+phjrF6FcJ7jsoebcHB2p4H5W34WJyArv+zU4DtanR
tPYJkD34RShSkXotJb7zjAz2OfyNc7fqmgWIYa1oKgU23L09vh5IKmI54OE5cv6P
qfrASoxHTbn2phxwLQ1oL0VjMxAyhU2PzFMIlfIfGNevfjF00LPZj6+3oC04ue6i
GErTj3sOjZuODbfSrv7ut8BIZu67+K+UeTX2GHf+mI9QKslxMBtoRQRiuvgj/q1v
ypP/qlcRMsrPwqPnV4GPPrTOoD4zhnIbxkPKPpSM/TSnaxTLvRZNoZJT3pMXCuvJ
kDpfULMlwt+mopKujbzWP1rkHCMxBq2NiC1rEB19G+lttUrPfUc379yCsDNGNDUj
iHMM0373e0mLSXMROuV3UpuVGVjq0i+jy8R2t4WEYrrOEsHsBINl3ZU9hG2D0J7b
v2MYoNXbJYGmsyI+QolFvqZR/0MBkb30Su8Jqaq9IAdInPwYcxMQTwsNsMeBaa4x
gE/qix0chewffaPHNfcLM+iZrKOQ4FGhzj8kJkSFc23RsQG08fe8zNy15TUaHfSg
X7iLlDbwGREypoTmyJETzq9AnEBbYljQCRebdjatZJjRj6jK8D+h+eYA5+amA4So
2kakH2KzX7C71+5cnY43ZpwrJY6zr/A18ooHNNs5IswYx3NBYvLfnjhDhK+aQmiz
2J1iu/v5P6eufWdSzL0l0CyOkcK2oRyEX1e+bHI7wclRJlUuR300IOlAj1bmPzla
j5Piv+7u2hgPHSwuk+wbYqlEtof4gP2Dj32XQDp5bFSb6bTJMC2QJ7A15J631G9D
SfHDp9Yl06unQq74tAyYQ+t0hFwAOZQV93Jky7lKwEg+VF4aR6/O8bTccYGOSmqB
au/oY1AG7u4Rn5jTrxHLAtLLuHcLYT3NofWS8lTmxP3tRCsLPKYH90+rGjHUoQFj
SgV13Ra2dbe6Re9NuY3e+0Jm+vMJWhtxLRlGmCNngrmtQpkervZClfkPNEifSlin
AQSY0SJmZ5umXaoXZ7j0sXfpo13xQnbApbCnu/vfq3Kgb3JlC3djqWmFYBEzzUWD
pPnodLHsg3fQciSoWXY7bAWfY5lbDuEc33gpGfM2RFOnV/mxTrjR/gvuZd9dNY1s
2AViKpO8+x2kobfXqUtlyxHdFzMq+pSCFfFh1luGQLiAVeiaGBEbhSEaJtlC+RWM
nfVkN6qVxGyDvEzsvBFsek+JcdHEQY7+ldpqkxlr/snlnmZfRtuXMbDVYYv/9rav
kOmZkeTAZLLNDncHSDu4I4uPHIGwS0D4P+KKnf44PU6i9glJ6eBNwkS0sDvJbxAG
smxmkK+M9c2Vb8FApjH5e6zboW4BNvesiAOIJCYDXn1ST3ckC/ocKroT+dyUtp5X
WoA0tXHrsc/B2rdf3Lzbm/aHKRcFuETBuRk5qDVjSgBYsd498+d8V0waUNgRThOS
mjVEsfEd0gU0IhKdutRJG/TPywgqE121678HNVyPObJd/Z6HHEbwzdNTqpLDIFwg
RkSEEcd2n8kAr+WLtfsiwddrpmKwzMuzfM1AYm/Tmzp0RNjPQe0m6F4VvQieSpBP
YfCEGZgCWzYolf6IErdjwyH8emaslVFwcVOoBYBe5fdOMV9rMr+Uyc1jHP1d9ZhC
66aEQNdTUDacqS47vY4hpPUOOgqSHghRCgVc8y79zQKt3hiYHA/7vEaUUzs+jlnT
QlbcV0G8MPPV3AK5EWzOf1QDgciGsX3F7wy198Zj6Tq894CssxvoPNvW5feVG/8v
wEJKsvWZFcTRq/ssiQoQtO+O2Cj47W7H20Fk2HrANGi5rbxe8lHjVcgzoL0j5vCK
iBVUBDn//+Y5nMbsN3eQSdciweVVvCNXh33es8NWvfMT8uiK9mWbI4xwBsNp5ro8
eai77paO2hlbtyzLQcAEQTzrrELzaKqfb6EP3r8RcFsReJhsxOBW0hTwR7tu1qqw
ugolYCym7SlDOaQ0PvlRMHiWcO2gqssqT/9HcuieqorRPQQH3GznNkReYg58Calv
Kwyyn1eA47UpKcLtOSfkZXfKG6tRUd++/Ii6Fs88pWRSsGhZcrz+Uuqt0zoIQq3P
cjKqYKh7Ex4R6P2x9G+9dvERuMHeSwbt9URinNJaFNVC+yWcXu6wsjq080mMlFIf
2c9WZZevBckehyd8oJtMqfQ4r3dRpVEMrhphDDEpPTnInfTcDs4mLkjg/Yi7wDNx
Lm1sYqKP2jZviGbQWAZGsAbCbaerP+wgC66GzvBVkpBzwrTmSbVrH5EOf76+sBAX
5VxVrN9C5MSyvASrJZsTUx0Yy/0CZso7ggxmVn9Ay+/cEZgFpX+zPMqzcTAGU6RF
Q7UYlUn8UaSHYnpEDuOY2NVBpEqT8bWvTA9cw0XkxJj8EA+XiyoU/TFhKzONYlL7
uZv7FMxEwSZ6otwVPjrMEKDa65+B/vVncbzU8FG6aQtECU9q4X12PE/+dtZcbHAC
kSwFDgoh4c5S57uekKbLmWWiqYQ76Sm31F6YDIeTs2H4V1ovG2JQFK9KbSORyCDq
7j3x25GjfC/uS5y/5Jxg+kB9INeR/o9ck1WWhBv13iKGYfMUdTvfmwl/nk0QE8bS
jOzIRCyYo8F0mvIL+Y4T4jP/5VSc4y89b5qjazaKZk8SVUfDIDa+Z4rKZ9P31359
iH48NPDKq4yfVPhkv8Nd7BMvYVF3bN18A/pJ0WakEC25lhyxFidj8+FdxbuBsajJ
NHPuxtvdWijDikQ/S/lAslonccJIYPVRLL7CGOfs+I9fc7ScUwB4F4eXBjGs0Gb7
Ri9FhI+EPMxIZrjuaor03niXa4H4T9hqb2KXlaKkxiA9qQSrUbiWtXuBxwxcWNlD
idcPYQD8PJ44w/sjGAv7dqklxO8Stt+8LqYx8XCL+xZdQKH1qgOEoom4KuOmuGDw
YFHJXySS3e6cawm+8OoB0kAHG57i92B1np7LP3j41J4RYyGf42bUhTp5nH173D/s
hu0XmpiASvdxHfDxERVjdSHMHuoT1GAXg2XriGzgbjL/WZuAE9Bp2Lv1DOrjSRPa
QZlFG5hCShdDOQtrKnuNXOI75AxjW3EqxtSj+tYk2ytQlyjNUiGI66zpZ3ghXtMj
Uk5H9ej3EBVkE1IztIgrOvk8l/VwUAYqI55hjuOoSPeY0eV0PAIF4hE61AQi4Np7
V10nnfhc+fAI5xsUvskmzWQu7SLVUDZpo7xv3yNcsBlJe3e8YMx34KDXeLX5thsI
XBcc0AsPhPTBqypItE04kqcWz96IcivFAZ8h1cTZKfJI8Hjpe6dROuJsAd+nJLxC
Q3k32Jv1erdvYbbFPqfVeKCt1MqJxlmoK7wwn4kKt0ZF/xf4whboa+qvU7JCGosf
h8L+AqH/4xeO7Z5xDW09bwn0G9B5RHO2u//Aiv+23thY4a3npadoMFI2bOWfOSRD
RiLQ9WOKpKvLPTDE20uyrKXc2B/2C3vlUmJldWM8H0NjVRj4DuvpI+6zf9xwnKOG
pFFyNAyH/sWGjS54C+lrWZUZhemHkc5C9LWcUoQhJ7nVXmlOrycjUcWTTEHRcDmn
+ykTN5x7fqdqXEdmPv2pYMUvlwSwkhYfuzWxTZg5o9WbI6GQXaSVRZKq2FxLDScm
Krkj6uFYOJe8WzxZxylDsOS/9VIzrHtPbrHCx1aNNm3NSGSmP5eStK8+u7iop/lC
ePeksDsuyYLSUwTy8qHUN/9F3o7TXpbr6mg9371eijdhmh79SvIAXAm+5x0bixRm
ZK7L4brPEmI/2j4itcXajwZ1YsyABQEA8RI/Brvi/7iO+LE5dHVGJyxMjQy4POVg
lur5UfFezxAreDLXkJ5ezIHqXwAk4XDdTyCN/tojO7arVTSLLhtOvzn/9Y8/bIGu
oW/en2hFLVoCRtLJ5CwTYHsPggtCsSB0GQJ2YBy9uptXMUUJOCtz1veBFAURoInz
HdlnFkS2ihBRIKZLc/9OhjXats5G/MxYBQuZwZ63st1BeQJ67NzOgb7VpK4zYhQ2
26xfHRzjSp8UMPrLeqMmrialDJVJ0+xM9RUS8O+Gscwxndan5pQ4F9pVpZicz3Rj
BHrmoCEJ4Pye0ACnhLrLqcNbAl7KhbCRKQkR0Ox4whjXkpKzXL79XnWMsFHdW85l
KVsmj0Ght949NJSKGWpjEh5DOQkD8Sn6i69FOEQFM0Wg4+OyshdH9Kb7a3xU+xlP
6gPHNAHhPJnXKnjC5R8LsB2nPpECLqnchqyYR9wRPBs4RF1P3smAMPaRCZ06EWBI
RsD/+oEjBZejAfU6EZ8ydFQlfRLDIYJRt2x48jjLDcY8o8NWD0gEjR9UN2p9cooy
nACyb/wZyoRWqrg5YEaV7pXNtMv38gk7J6Wnt3PkftRV32rnYokWYBJOfYY0V7Yr
n2K/DVsLk8elAAPvqgtZ7/7CnG9Lv0yNW+BHltIwZLX1LttfqgWnwLKeJkhUaP9M
hY2UyvvN3zvKVYF/Y4Omuj2bjexcXOv+uI0PHlLZb7DfjKAVEGD+BIm86iYsfEcx
0supBGjsOQP7piE1eVOCNsgfRVijacY8gr3n6lsAsKnbLhDvdoPHr/uvLpq29p5c
1jn7IqJB+I/HC7nQH1TMjkmq94Y70VM2ynhX5BNdbeiXGxC+ssHZl+LxJYhTrscB
0oTS3feuRe/voebbMPmqhF6awJHBGAMAf8X1IST4emrh1sdghAznTKXpbBtBjGVZ
wO20JIMY2772yh4EZnciW47NK6Ai0IKH53CU+rzEl1TkXieyEp+XNC0d5tg0GfVO
DAtzExm/zL8AeYljfqQJCqGjDTf96FAFRBI2H/yb2nqh2b7WVmUos7wxz7M9orUc
6AWqaQ2+PQNCWTx4Eg7kYp8NII4SwCboDZKgoB8F4xb9xfxogcU0mI/fzWux6oN9
9pGkOHiSlLL4z76ixuxLEcaN66cmRw2+DmdCcQZOLKtZxKRFvqYNi41mGV6GUmRo
faynCgexMPdJQfSLbzDCcMMc7HcIttKUY2NUuUJZZMDawZoXwh2ZfIVy7UraqhXc
Yo1y6sMJM4L80tc6jMY3kQ1wK33I3V9TxJsy31i+NiBEWKDyPUJTMdT4+tHBjO+f
2x1mofWPmWXRLo3qtLMNR6L1u15eQcqWy10a4CWxbnEqIpXeIT6pElmoz2hWJPkj
Z9404w5oePS6KaDfu7UpTIkKYJyFQKOKhX+W9nfiWg1ZINQ1vOl0u7DbU/jPnEZj
rSDlFs0HwzO2NkkTHJ+Cf0wRDSJuPHWzdFNFB923/HaL/TtprFrNGSFtTrTxJvv3
LYoBHt1oWOxBkDk3MbHKn2R/7utrdNBLoCt8PMAdNmkm2NqhkphOL7B+rh4XEnH9
rjx2K33gAdrHPhfoR4MlHSkMB7b/JxLqDfY5KtL/Fott6745N1Z4YDVeTgkZL0Bf
e1HWvOWCVvJn35O0Ntr75U8CVGBq5s7nITNAMb+i3duJElKmx/kNKQ9J7w/vI/ZV
FATAvGzS1jEpfyrSV08eI2Nnflj6h9gbx3uxDb1Zf0H8Z24vOpidv5/1UWve0y9v
Eic3t655UhPwpHQFHV4Fjl59RSvdp9ASDriqBm8a03mLwOnsow/PRazB77ERZijs
uBs5KWnDx7R0MDRVxHiAg9UInlhq6AT55pV4u3zrt/EH2PhmUhUClG01GBuBCE7W
LLM3RcnQISJMudqHxy81Kuc5ImkKghFseMutmiWIOEFirlJzwF4AJKcVNpek1WEj
T4cGWCP3lWejm/ZqwT7sno0MHepQ2C8WkqgycW6Jt4pV052hfFRMEMY3lOWPRW52
k7FgMvKgFOV2WZb/Xlr4NVisfTi+uZWP9GbkAdQC2cJOXSuocYsllq47JwBEaj7M
Jkz20/7RCipB61tZm0O1HoEQiJyrsT2/7hYWmfIC47HgV+hT2cz65toAbq+uz2sC
9srmCDYvbOUmg1tTE8nP/ypf0xS9yevxjZzgS6O7nHcZVpNbtw9xe71ae6k62KFd
TXIyr9F1V63GRnsUidrNkHz/w6sL1KRBdFiw3VnU4ys0OtlLrtD9Cd+8g7jeklKr
eSFwbcJq3hLlSMA3mV5PZUyGCbrs8vWBKQ+KI1/aEa5VYdZbjOlyQ2Lek+qHhNTD
xD53iX4VzxIGHSAbBWMg8Yy87nASi2THLZGpy3WJheNs8PRvp/5bwoBvHaSe+E9Z
cwlz6dwShjohfkuhxA5MpXPemTNbyJVzSwk4StSdNoS3WTBdwrtVJDLSynO3L6Z4
v8tRkh4By6mitFRe2hXrUsm9Tija+TaQwlIwyXFeLR+uDytVjUiy9UZ+MRtZOGSH
aoBUXh/LgEOgRjtWvU+bBmV6sQZrrYj3YNBiiOPtb+kwdVlj+a5ODmFBvo7LB9GH
AunvPx3dIVKVAAD3aHDwSCvFDjEia2oI2TeQZ4D0rZOpktoEPAxBqmhtsylVSwJR
Eb8nsG0khZcLvvWpkFZi5e3og0fhwqvjPCZhsVNKasNYt5dfb+z3NYuBPsXDZVoV
W3Rfx6A3ClqlehelOBLw/4xXK4p0ZvDeykeEP4KTbZ2dGrXpA0uxcuJGaSkW3e6N
Ifd4XNQ0FphZbgTDvB7wqIDZsv7Zgu1k9GgoOo+gA4s5LvBLjAijSkmIb6cCnGmT
Fi/yyHRNSdcF8j3kRdNPAegOXLHy6wBeXN+s33JST0Pg0xpIonfEPLHzJgAd+XyB
78fSup+grYH3JZPOGE8sJv4iGpFgpJuogDc8xomZG21MUuHd2CIGUWBmUdsN6KqU
yLuU4ICfXVHgMINitvS41dNGhU73fzpQGAQh+dFfSpSUc+elyPQBPVdBmeJOHgya
td6sbFGA+ysTDGiq7RKz5dOAI/3PzcaHzdzvnxapzSeBsa6/YG7yADUdYCxMaknt
4As2FxUT+vPWifKHQK/QQo4WKTb83Wo5j7npRNTXA1n1SrzeMlDLtLdRkpJf1nPa
k9iJyi7i/X7n0R/VQcJZfzbrJliYCkAQwTSPNBj9UHKXis6pXDQsbYrDfvjvbIDq
zeN5ZHdo7xbqT2Tupd6nDWvADkD9x0hUTxOHd3ZeNizDzt2eLY63kkO3Vmni1Yc+
dmgVAmW2LXPlx+outgD+VkmXn//FromLFyK22dPJLPY4JGUJlpa1EePvt/JRtKR+
Of+9KcHH0C7vmls2DUeR0bhzWmiSlSwlnBWsdOY/ndq6YZ3BWaIdrey2aNcqcXbL
zZhQQyeSIDg7Q2a/6a63GsJx1Og5djB6onWszOmZJ5dDNt2DXz35RUkXZFCnGiPh
6FcausWyI8bQWtQbKDCBX3966oZ2o7Swlr3sWYlTecql/d+PZmXFUWmq94GbaYRB
8GkB/SRFx+0fFcTYVw+GYykFQa9AUW/CgnYkhSl4KEZyn12vyyh2BxUeLRzPez3s
nSYjE1Qls836rfpoMHKOBck5+56Vu8ZNrLpFFQWcKiSO/RjCKPGfPJtStP+fFLOo
bMaDY6wRV9RlpXtWrOLL+AViqXJbfIGCZrcmJSH3YtHeL8+Jhb2s57Fc0F/ZKB2g
RJ805G6ay2SqszUNmFROD4Qqrc74pmSZDk8S3nNFvP0lNkSUKsnRZOkqtpWawpLM
hOtM45WSHHiO2Fhkn3TkXOht2IERR8uwvsT9D0Nog1LYbsmqZd0vUFZ64N7Nw+CS
vYIHu6pVe34CWyIRFE4P8fDiy0F2O8vz7w7rtb4zBX3es8XtNNjbYuXBbD4i8zkM
bvdw0/F7WdjLvyaib+7jGgB7aiIHxczY2ApzKwgH5WTvUsC7qLMhNnSXfRkQVBxN
XizK5zFsxLOwP1913oAJXXqLUukBkUCgxyqCEbcqYDPinyF6ZPh0ZZWLPZMz4UXk
xFeH+IWCoifWMi/NC+a8j+f2l5wZL3QhYr/npmGrNRB0ZCdxqgXM5zrn6tuK6T+F
sQ9x17JaXsDdStr7qkv9GF7oSke8lY3IRN9bCzK35M5vXsi7bRVLGCF1iqXgSx2d
hc+ldIv4zzUnIzdVyj+g/4vX3dmalGWqFTd6l7SM/KzWn3xih/0mfEmkzm+lcJVi
C/X56qkVe4Dwyc1PR5MAj9Q8CZUXo0Rulyoqi+lSbq0YqfQHVtNfl7k1ZnaYaKBj
ld+LjBJHOGfHnmOtQjE7x45XxfBL14On/HJijX6LRR1ZrvzMBXqZvMePwyKsGrTT
Sf0gAFCzHNk9jFyxMADfPZBVM+9vCCjTiB0v2HE9v/Pq91OdsJ6Y4Rr9/sUow77M
SCnrFizWeVz+EZxDsvOi8JZ1XDFw6eQWRKAJi+OTdlhcpvdvZxEjH/I3uh14hE8m
0yiy53FR1c8UKa4AnB8LBICekooahhzrvuqCbVghsjY6jYdaZFWdeWtI3m2TduOT
MzpUKaCX03cgGHnG6a9j4+p/EZQY7/V2FiWYhvxJCxtkQ87DSsMRBg0vsEnJtjhF
gAgoIuDyZrOXUEPcSmJOh9bhFBrVWtgLRlk7WQofg+KKFxCvi1cDZnM+JXPNY0Mp
9kvZAs0YXGaHRceELTc+LBXaKNcBO3xtpVANZisSiRURiJrEKVi4rPjX0YYw0Myl
EHEW1j+i1lJXqgNoZ81B6UiQOtDegdIxQjqxN2wq5SpL5etZ6wN88gBo+dvlpOJS
AssdrNH3HK9j34HQHyE4WznrRLnz2MNHo8If5AzO0xMROX1aNto2/mkzYVN+KSkD
vxYBWmebkzQtHvvFPmvzJ4v1KNHvB61m6B+n4d0XvLq0dnLUp2cGvurrqZR4ttQv
KGuF76URqMUCzj1r3G4oMhvhz6wYYxkr4tfjTZpJYuB90L9p7xL3hsodd3A+uu0b
m/HIMwDALLOyk5q0sD3vSXd2pGeDB9S5S/TVEOJj+3929k8a5tKgGLXEnHyJ3a3+
sAHeM1qqmlrX0tMIKINH+HoTf6Y5Ou8bXXkX6upF5mJTr6BY8NpTLczMtNZw3g9r
Ydja92cyJPLSPOENbK1E+pe99xdhEdw312a4sp/zuthloZ6TEuUwwMajlV/ml8G+
7LquXtmPm+C/JjXb9Bb161MZKfr+Scp+r6YXWc5si+E/R+xs1PpgHFQ8trXrqtpU
DPJZHykQwx7e6To8iF0hgWriFYn+Cle5cBEsbmp26v3IxjZRaLP1py3PjGNus8Ff
Amhz9ckEKmNErayO46Kfc+Xhgh8eBoWjccWx09MDhSVFijYSoQ6iyvY01Z4FPumK
YXYcHprtryNyjtD1jrP7VUhEdZFSSoqHjRI+uO88I7GPRX5S8VT3X1jZcncN2yZo
Wk6Nah9fKIiGYOkjvQ3/3DrEVqnrt/f6DE8ZIkgTJPv/48OGDiRW58gOEcqw2IVb
L/IajT8PH8p/DK7Y3apn03JPzDd9pyaU/1eY1W8mWkipsKmeU083VWqlgU8mjuQ+
3mhV8mFo7AKnwl+i2KpWB5b3B0TEREJ8J+B+n/i1P1q9BcrLEFg+7WiIdWv04xvC
ObmeiIceAFsGiTMYfQfEAfgexhK8xJXmjPInPcVswPCj4hNlnklRg9Rp14/hyXHQ
gKrOTY34zuf9AEQdaCKQgAlHGEvKDkUbD67ZhebX2+4fuJsvOS+tDdxTBsgSTPcP
fSkwfTz+cqhfI0Q90jeeBTpMZ1VwMJfMQEl8cm1DsW+dmemIh2Ue0a6jlp2doyZ9
fMCI8ciM2CztfW1yVjqncFM20siewMQQAV8eCnzWS19Vc0glTd09INUPChLigUbV
UKe4OeH2vTuqetEQNsP1T4R7iCb0kXpzc7zAlVABp4afinmWS93T9MgReTmxJQRm
g4K+xJrTrK132AUZjwwsER3wwq6ErO8LxmUsebStuJLI8/PNozvADsOBPug8PS8D
ZXgsGGnZkttBcdYU6ifzJReDGkUtpgGiQxCweJH//YHjrIc0PGPQJF6M+jdZ2dhb
6Ng0UhBzDpCd57FDZx4q2JXmoa54I/dwtJ1ISzUOKfkQGUAdp/K/4VdMYzQMQxIX
TVuzZ1ZRLpsPYVkzDnO43RLKqHERkfp335RsGC0csQfETGGenVZeU5h5HdREFbVe
CS553HQD/oAbRc/xOhDz2nrCrG//ZDyQPxBgQyykw8YohCr71Uy9gRQmSkWW10tB
Cf0zuPsiVVt3OgM0ONRmBGjnZToyfYk7KxWzc3RfQy/VWtWN5OV+1MFxIIjQCtG/
/tTm9G9EmgFTfHu8qB0FLo8V1QDaCTO/o5ZcOjkDCYdbKqx818HRa0oIBWmXMQ/r
y0iWeiukBDBtfEUms4R7C3c/9ej/8YT+hUp5a01vPoDlT+xxrWsPy6PXsbqBFc5l
cLp2kK12CMgFna3sI3DLWxkt7KiEL9kEDut70She7G/r9Cm/dkXw5iKJMt6cvUx4
WkOgs1oZ5yKKlGkQm8ZPPiJMdh4xLZrz1QiLYYGJZeLwSGNfcnGGQKe/NR2xP14m
qAluWN579Y7kTceKH3CW42CENb1+JVuOdcEMscRMo/pG684G6iIY055tqKc3Y+bM
oU/5wfScWHquhgSAeepMLUBF9C8gOMwwnuxbMxwNFX5miuZMmiAKgkCxil7APbB3
4GjoBbN0UZ3qfOog2ROpQuhAiPaXyZ8FP1FHdl4ll5ySdtWKG23K8tCwzGLkjvp3
aoLzLbHYvY929txcB/SqRs4l4dtLgZFq7pOoAnFH6hpsG6qZt9GjRF77BTcEIfYP
yQx96zsMea6BTp7vwMk0uDdWXQePNfzDw1NV40uiNG6BoNgC3Sjb0vbeNLqcIkq4
PleT1V+0NFsdMtUUAkgbMTe1weEh4tnjejsN9lYakeZHCNgaVVXI8lRCTdO25D1A
DQU/xM4neAJq3UedX4YTIzEfyzer06xGGJrsQv/tQymPdVnAG3GY+mzl28pOYQTl
r2tuYAydd5EYZ0uX53bPBwTkCq6rwudZZsmtjyr/nYh7H2WaqiWk3nlhch4gnpNj
ogazU5gK2kg7tC3GDBqF9QtUQcjuGQwArbCiK4jm9403hMAjQZ8QSp81pAD7Seji
Uhb99VCAP/5sXp3I0qfUyvhjkuI3fV4omE+LWe5UauCTOh0pAcm8i7l+kQtYNUGM
0xsPKkFqwP/3EvS2xu7waD6ZN1Wm5TQqbHw/qTvWNxJxVO2yU23/8wWJiifthZdu
u/rIDqiQLOocAwf7sfyQR6TIXmncURq4tTH0QoDPT7giszy0HA29S5IpmhshPNLP
8QfN2bu01pzn430W/qbavXsNpHU0k7I5C7TXdZx/ceo8x+hErPUFlSNxO2AdMypi
t6yxX89CxXIus7evfj4TTlQrSy+COPYStxU7P5W7bzcQYETw69ZiUfHPqKbP5+JP
KDhcB7eQlk88SYb06Il33/y1Zp2B7XxCr8aQTFxm7WMCqOsmW1aazkcm2WWDyfC3
KcLKyVC1za2Y6RMSiAdtf72l/NzDQMNJrAOOA6JA3I45b0Mt+EU6ZCFnrf6/BB5i
2P7jnIcFTt4/4yDfI6nRbeG+Co5m53RyLcv0XpVYdNjuAoRWpvGrXeepGo/gKzPm
xklInZC/eWbM9/t4MbkDG83ylXFYW+O+D0gDbg0UMyNM7eh/kIhl9WSk9Y2zfJWB
4n/UO2gP8pQnQtmXA5x4nJ8+auwGgGxyAMyVwjYjCV64n23AJJiOTZPD8uBUt79y
2h92En8RIkmSkqpdIXCUTD2Zf+UD2ANcksv9+5SZz0WkE4AA8XxqPNFiXWhVEfnf
mFQzJkum2yx+8iqY2ZAcs7YVqfXSqX8dsdwcIO8qdU5WQeiVIHiHaMI//Q0PcDEi
Okc32aIKLbwMci/Hya5RpR2knj+zziZCY9EtyF0OzUlkEVaCmN1Wgqab8JraWv20
Yhdm7JmlGBmkp3zTTJZJktEro1aq6SBJBxI1TIweMmkXn4R92NanoD0h3Nge5fy8
ShaIaH8N+0mYeNn4huLRuf02vJUsuQzjcMFhRYDjVmL6xOxtFDHiV0u7MGNF2+GP
EAKPZjR7IpeVy5O0f66UerAZgpN31AbRYEpm49lxS8L4puRD9QYmKlksoQEjwUN+
jd5uQfNK2l3EauygFyIkuDGS8TNIq3ub2yLFSPJcqlg0b5QNDjlzFotNqR9a/gdc
MHSfnkz87Jf/O7mUYTRURj6IjGtVIHy5PT7Kjc4uVYf1PtFwbU/HCM+raokqQTqG
B9szRZKf2T3HsvyYym0vP2RTjHZ5B+hakvHioVw6gZzmu2UtNHC88sNte604zlSu
dPMkHW+cBtI8+1+85E7yWP7kTByDCyM7MsEoPrtpiqLoEjWGgvHO4lyDm9HFgasE
zHgJcw0ike246n6MOg4MP2fLZaEkBir0z+oQnfT7yOyad3h2cRyPMaD9gMiDkl6V
i3htmMwHXvLbjpg/PpwDwfKle+l3ccCBGoURrn8pS1yTDglal1fN+UCUdfeGHt/b
kEcFn/aBWRIhvd3nYVaEspRpvlRBHgffpONmXFCxnWGwUbP0THb8+m6AFXOZM7c3
TcaqqG/IqHn9hRSAib3muORAj92dnTqUtbNnxfzW32iaaM9T2DMhODIsN9pGHR7T
LFtxrdGvJ/Cqp/vT177SsBPS5eX/VA+OixBTbG0/lqNJqWDJVE6GfT+OSjDU5FPW
NnxHTtOoSwLU3m5aHhCvnZhyA0IKNNOxh0+G+HXO5Sm9wlFPtjlZ6rcfX9xkOzOh
06o95TZHe5WNM8jQiVhN0uZkSCMFO/8klI+Wjy2BV3iX1S2Isg8boMttZmOhRh7+
wLKhxVs9tN6tLCvFg8/AfrMgeR/hwOV5qDm5zhLZj2mr5d9fdDdFYcOsSX6cUvAM
oQpx/4leRYFnRxjXDdSrY55HlJJYEykKqSIW/CO+xLPXIhybg/Mmh9QqPczMkW/q
n+0sinVtmrVioPALEIZ9fSvgOy3al6M5rkghGAjGOrNFYsu2M1Fj9xECkQ2Acf9j
j/IMMMpimBV1VmJgJIClJNU+8yZU38j+FpzQAm9heqZcpe0hHpEC4fJ1PWbM9r/K
i0jrn22HlRZQBv2LGnuKAxhvjlco5M+OBxTqMw/nYTtKYMoOA+HQWJQ//vUR4DsD
e2i3vvCc30E+AZ0sO2dlNo+6MRSCxL/2b6kl6UyiQlR5sGi9e5XiqB1qLJ7e9yG3
rMmnJ/Y6fPStPJYAnO0W9bP2gStFoaEqBAwzIQO6rZCnXTvZweIIbhNtR+h7jWc5
TYfl1qdUL64Bj1nPekCXGYYt3zlokh/q77Dgvj6YzFO/PZT7GML9ubgV9Fe2OUOa
wX1W4cm3NKcUsT7ctDqcIX9mH3NLrVcgio3piM4hiWfJWrQNodfO/YK761+2f5QT
/m5XgirGe7D+Nbj7jlFZzcFlEecn1avdDqiKZfFEfKxzHuQftou/fX1rURNmh0oV
cH7r/4Rm0pYbEr4qD9rhfYbxrKtqls17oBSuzI0MN1CAqqpdGnU+NTkd0kzxGcVs
gdRyxbW8XNLLa0+X96Zo9JbKQPzXlHUXurv+jK9lEpaIZLHfBYvakSzR6pnGVEwm
T1GIlkloZcNP0ZViwiBXg2BbVtm1M0gXzqnajGlneBZMU8RnZU8mIDrLZXNRtJzh
04K4RICLT4nZL08H7dnEpLrblrXVExqyikD7xtQcxLuoR9ocIwnhqtHDTyTuIKxa
yfEJB3i12bWNMDTSlWjczlHjREWcZ3b8W9M/qh49szyFNpM5YHS1n6xcuPNLeL7+
l3naLznpNHtyUhNhnMUE/FO9gNHttWsl+ylP0AIijUsoFcjFfU33Id5nnswSm4TO
zvx4RAjrziYHndfFJ15fIwUIgEXGyrSz/P3g43fONqnBe0Qoelel93mq+NDzcMmx
iZakt08E+5asiqFFq2mmJl+mi9JX3Qke6KQNCFZKwLVhTwtWuspIhUzuZoTMt3Qt
kZ+VQaHHBguzIcwEA+di/MDq4CaOlz4aYHGGoQtKR/NvlILjHQ4FqfyjrVK/l563
5I/1uTDkN2NHtf+rJ/FEBSBKzgfsVjaXEEgSW4MIEGOmo4wJk0VCC/Feq+IOODJh
VEgmfviN1PNCvGkGJuU+KHOcyCIV5qdN/3DYQfx2p98+TyM3MHb27eeUIpk+bCoB
ORz5WiTSgSISN1HwIArtLfPsUc3Sfz4EmPlgtChusvU/GSPqoogERTA5nLrU29VV
UBR94Oxfw1N1LG27uQBUqgFRynj0H8xQiChtB1B01EQketYlh47U8OhFgS7mY8Zd
7qFPdY76qoUD5CjKkkBwK4KdXPNSEQdYoSODGsPJl4jvk0OQRI7+bpkZdfJRefnH
jdTovCg7Xv8pp9DUgYN857Vjk6ftLTAZsbUwrEPyixQSyoPkwAOEhDBuZDnVrtUr
7C8iBnFenSVHlwm/Gdq8KXNzyCmR/j4Utm32NEAb+06dYqqXkAGJBJ8M8oGZnED5
SaLY7yOa5Msnq9yjKYdM371+LZjp55Av7Jlo6CJJ898L83r5efz6Tyxp9xJBfAcT
pMPv9Bw7y0OTT6an0CUzO0Lp+f+2xkBoUNFtftXkckU9lE1T7C0r7ha0fofg2qDN
FqTD3B91f0gUWfzO7ncADkfGvR08vwCJQvyknNT2oyhziT2oNaTaDHyOFzl1rKz+
8i2n2+cBh56aUV8QZQPIvg93xbZOyGzcBJDsn2FK3D1g/rbgS1tmy4J6q1DE35NA
ZuM9TYTHbwYKvhlLaB8CnfJZuADp6t4pWQQG2c2jkHBzR3zcJckOFSoafvkcM1hv
lJFJYs6LU5oLn1pMo8a0Tz+ml8ffpC5qUvxHHHYNFTYHMlTxZ1Il2wObLyuN5vwj
uFyOFoTlClNZRcwwCp570F2sz//QSHLpkoeFhnIaz6yuElOXoPpsEeJQHZKfuY2A
oDBppxmg3VzalLxoLP2DVeXGiNAHQlquoVr5FabO/OAkhys6MGekJKsumIXBPd8b
MrbPKEgqmAvWlU8v0Gaf9mdsL7lcIfUnPtmy4++qx/yccHt/A2KOFYEQWSWBZrqU
ZI0ExmGGZPc3JJm2xnxLYAhcaK+EnDWSyN+nSLen42znsbPxYdJ6+uqIMIVas0+/
kjRsjdO+a8K72QqZxSISGXZLvr1C67nzbLGUM4c6JuD2KuIdupAjLt1N3oCfnxeW
p7aH65GCEf0au5H2s7PsVZ0IKDD2xPJWiyinDd72CJtAjytKPshjIY6JnVNARe3e
847uThyNajLClghZTDOgbLKQyMwCnhiQVFzxhlWcSxiC8zA0b8d6b2iv8nzGnjX/
egKKmD+GM/YjGEcMugYHRlQ8CDlUbav+WzMdszg4cj6cwY4MarbTW8WIM31OOs3K
Hr1TSOGmb65cPHkTcOfNVR5+HkShviWMvHpvrqu2X7OpizMCltZ0OdC3sgcXM006
fbW9baqzuqDK+xW2TrVR5wysBuVVnDlNocX03IreC3KuQ2ZW9/Znn8cObMA46qyc
0qh0jW4NynADnYmH9pm8e1Jyq217clwdydy+S+hXqbK+SuTObANVG1tO5wt2ChDK
G0IihmdQv/tIDvmIYTPzjlXfJ+RUX0mT6MzMc1wp2EfWX1Hpo2p43S/W6w24JyMQ
MctxVt8rWXlFqQbssFpvSKIjMhGb2W4dLTBc9x2njmr47pkT1IJs4mHH+mqgWeHq
0Sy+sr81oz2Sajg/vxx+3PreTweWKH4e60m8/zvKUx9/oa/7uIjaMvcjx4hVtuxy
GA7AGvLzwK5vIXGUb0YHxB+qlSEtbkn4eL0V9FBoAQQZXjrStgG+MaELd6wrSrVi
lN/nAMyNJBA8fxIJljnNX+wt1MkZvZo8MckLjVN2rK248LszeK3DKl/N3a14K+ij
J2lG8tLY7eTTEPgqWsx3LZ1sLHrEO83ufl1UbG4yBEz7DuvLX253bcxJfnOuWMkB
L1KpaC2zOvd53ucklGxArTZXsWpK5rCqCIPwgp68+oeMNqhnr3Ok4aPub/9a0WX/
GNxwRfQAXDCEEjkV6CIQRX2BNif8015ur1ez65b/HQpx//NDUus0eioKQraN7X9L
jrW+MTjBVhl7XFAdWEX3STK2ShSu9XENkJGJLjOInf6iBCNBtFwaN3CMWfvAM8gI
Rbw9DtQeiLzO5fL97ZEW+RNYGxcsqH7xcO0qiiZ2z49HGzTbiwv0sVFjoTtHMK8+
UGaUdCxpRLisOK9hQ2KbNvMIwVR9OfPyp29+Xpl3A3oNU2spVuNulxZSFp4YDdgc
Rb31v+fp0GN1Marqv3wM7h6+0dMyn9NwcNsRDtM7RtO+KiDS3mHVYuL6cNsTLQvb
k9vvL8yYQezbdeoQUTGq8rMHAT9G5Uf6LkbFzpR6iFFouGt5q2ObOa5jGjxeR3KD
KKrbdIXIi9a5zJehTnCEzKCLBCckRWPUFwxI9Ji2VSYIbQrC5S7YDBExAOxNdsT4
MLIhMXU+nml4QgVOwFZV5fIRb3cvjL89hEWjY5aIFkmQt5KFjuDhkaGQkMZh1hVD
VkdL5hRRQkypWXVclVX1KdWg68XLjhNH0wZWkh75jvXsHeTKpkj9u98XrTCl+vLF
RxIRzWW5CMBFqsLJ4I1sNXfcP9BH1Y1TaQ3IcdGrSx2Mk3S0+XMxdSZW8Q7EtyFi
+p4YB+i4zl0OxA0T9Qn59zk9v2Do5r808Q1IzH3ZX30fdHAdSUjBGs45pku3QlgF
MJlnjTKo2zK46EjqO3ShRdPL6TKYwT7OH51N5Q8lDCaqbYPHgkwFlEqJwRqibCJl
sxQiaRYc6DiJYzVMG2APUZSVCS1frIHDN777dYTzg0r5v9mBRi7TXCBbyGMU71/5
hpgJAU81Rgj4h5xILOCaXGWcFejdnXGbX5j/CjwP/hBssXWXKFT7TZGFLNdJKTCI
fEYIVlFIXetK6GjicTZdpv3trBzrJWvILB6sdot05rQIOpY41nYQXYwW6wEp9Af3
C2hoa3nEC3KTwxD7hOnbkQQgzNn1fbQa1HIl14EuCYJZQfCruAWuwS6BCXkP5Bx2
VgjUNzFEuHe9oOrrmejwN/JYEIFFMyYT2bVbskW4nrUe6dF4RLhZQHYKS0iSawng
aymD2t9ep04m/OmpXk810udwDDakkYNk858FBhVty23yDPhbZvRT4mOPrGHTb9in
Ix/KAQaUCE6SEGECsyPsJs2V0lO6WI2oqdbKKXBEAVgAI/iKR6BVIBBL+earz1go
+BE4XwVKYVkNigQ/O42Vvgj7wTnE4P36ArjVyIHqMPOeADVBuwslgMf9XDdm/a1C
RocWr5FbPj47a1ceNaN6aylTfCrtr/giVkNp1hbNA5ybBaz0EC2X+nMFQol2w3KC
54T1uQK7NeLpo3leqCFrluZyZR4B6+RzEXl/lZoKdcD15XwzcC+3QVCie89NniOs
QSu5KvLiQkPDEgpVzsADYO6fNhF+iy7A9uKUE831gMLVOQd5CwaBFFD9eC3zuVjq
dYbPPaY1N9mk9hczWkWTSGXdn/jhJ4ygYJ4dzfTy6iMUfdHOB5yIyu04Tp57BvM2
Dxfv89p5ZW89crOKbK9Ockrg1uELtOsIJ7XqqoJfbmeLfhm4OPvJN3dJGdhMw+Po
sPpBjoRhW+BGuDKTa0J6zT0fJvBEpbmc16pLSxTRcGv3wTLNF7gNJSCy1l0Z6sbj
FmAiLi/5wm/mmaonQyDymkEBPVFDcaUAsDzGomcCMa6+sFV+3faoMF073YpV+6vB
SlFCqEc40h0mQMO39pxNsQ0ijAZjbyPviiLSsZwpDxqcQRRWW/lwKep9pe77+38U
UbrxrxOan1WOCGIa9HSY1zR2dzppgFo7PXjm8r+VVlYaxu5Dqof3MECclVoVk40F
9dHXnLbMxciz01S5inCS72iy8qtjSCIXxLx4W7JD51aT00tqdKvshRJA4iqNhB9k
uWS8BylDhqZIOJDJpGIVIOvZLbi8TLV2gZnsNXFnj4carSSD5dcacihvm/FkpO4A
CL60q2ljgibZeFzd5iclTScUjJ5yO01pxbaC4i96yI7E2RguqBWLfN2/iYPMaZ5U
EVy4Uz8QcOJkiTcb02MTLBVeJ02+p20pteVNPmnbGAbVntXvbumRZa0VHjW5oyU2
H5IfKea0KG1pe0pOq1tGgeZybBMvR0dtqs5DIvoblQeDyQwseitDBx0BHlBLVGYz
cJW9th44ZENIXYksHJ/DFTaNsiE2iUSbW/4OmZi/gnQEvIKKFG5sl9pBocLNujwq
l+yh26AicF5On2M9BYOa6t4dGpaXByUy/vUj+a9R5fc+85dokBQD4gdcK3jsYfNc
/BBHpsIDPdQjAfhmR7TnaJf7aJAjbUF9brZO4AewnFvCyyEm8EyD1gFI8BSU6NXp
qcV/TBA6wIJvY6a+wJe+5E5L0ijfE5xm8tJ60J47tvaqx+ZmfkexPXJa5cOHWzK1
1FyvbIexvEODjIkEJ+DLsz9gPc4BPZFZL0GISSdYPWwqNSKZe40m9EHUBMH+5Tf6
YG9WaAInU/1HAqxcg83Y4bw4xqRQl/r9UuHh6R4HC03igASVq9H6s/NVL//i9h+N
zTc1nfbvYWGj1bggAER5YO2Nx7vNheLvqUFJ7uh+6H5fbumLwqplV8oV9fCoj3fg
w3ofnmzpGbYMXd3uk3Uai9gKTNnxlDrEB60ysiEHjjb+uju1uuFjxeBfCD4JeVQL
9NCAyZe+gh2QaQu0O+yzh21vaNtNVcljIlbyjv6DqGZ+7HCWRVtQPYm3OTsg47Br
S6rgXtUkj/ndJfrlmkDN+cgzMvA9OX3Oz7adkdZXofVfvOVuzrn04BerOHrRKppS
XpdGfntiojSByDtxxzfM1GYShAXXg6xJ6IGzixSmABgp+vXmJfb94JBmJ91IbD6S
ZfuWneaeytlxreujD/vqm51Q8JjPA21n/ZpFtyKSWdJMloO1obE3xlDK/VCAlra7
sMbxSN45m5psz/8WPHVNV7MgNxdFy/DQTEZzLGGoqAa40X4EUhfA94dvrv0Vm0aS
QfhWwpAR/xijVGooBv2AzPHx18Q1kbmbHPPgHVFArS1fIdF9jQ0YoLVSRrFtIYX4
r/m4LRvqELC4QC36D45i51FBmJydYIdMzkAt2bQ8QKMcXrv2a8A1+CQTO3LxvuW4
/0hRj+bA+dBX+C5tWwM9QH1Q3kaXXB0W9DFX3/Cjv8QFeGROsS1J/eqKPD0uy1e5
VzGm1emfAhp9APClFMQTXMFnkeQ9iP2Oc6iacbPm74cTMQdiQwTGwE3PEES+gvZU
u5z7HHlnswYcgPDsxIiyGkW+QMaA2paWYNZVapnCUFzjEiPJK2i1DKNEC2EWZly0
GxlfgjXZjtnUW0ul2Mc6TSF0pCE6JdH9QLx5MT+g0RQdORiX/BBknK9a/+Dk66lH
CrKtZbrmEgKbRHn1InLGeVh3UJh/3lzkTBWAMkyppy3GBapaX030rQBbqWuhh4LC
Ghn+Z1wHQ3g6rBCJjZ7s0apOA0tqqd6xKsXPYMmS27mNsUCxFTpSdikgBZpq+5tK
v2tFkFkozuOrv4MX95et9aOKxq9KU7MmPwPJcv7Qse2WY27LVKYXqiJuEtf1AB7o
f7LpGNY4otD6I1TglYKtxZcWYB9+xd2ez7p8WmWgsw8GDpgj2bjW+ItcgL1j8Y+y
NN25XOjC8Hv4bTbRyYs3PwhUWl9RXPFeNn87kZ8kkZb9kaRw02/ws6BJ8Jqq/U7X
1JnfxTvSkJOwawMn10tqf1IHi3ZvsvMr5O+aCRqkf3QaJSrXQfo7TtftSfSKzPyy
xHHOrZg7Fo31pL2RucsjZX7jxkZinaETVqCmEjpvgr05trtkGmJ4zujxrJumRphg
Mx97nTLTp76h8fN2MFTyvgqk9pcVXvtJqCA1FAZMdbxosnIR/t2Crpr3LlxMMcBB
8qD4/W4FNCvJjU4qfCrHEt4KQm8Qmfxs4g9deb+ALsFTCh8UdeMCEvQio72Hwi3Z
sLA9ZzAtL4I6r7kGViU9FY1BDJdJnnFzajTyNFgwSOpW6enw6aT1qicCw+QpvxLf
RuA8l4RWJFjKehO92rCH0Ej7knhpdzXXPNLAXJV2JvPX5FahVMb4JAqHwoB4OLSM
qb2FVYKlTssl2mk5fYipmbuQIZyI/pjP5UtlHSPGSFc44FzXqx6TL9oqw2NtVuBQ
sWNIYBZJ0ePrOT+8RD7/M9qzR4rj4pAxKhTvrlSRIh/SBp+pH1+5ivS23mfnOvfw
+sU9p4ZDp6KUj4TiY/AUrnFQCvjJRVSk8DNyxUgSj6I7UtXjojA2y0pvhCtLjnNU
G2p7TZGto7P4XnfDwNNbpt1FArXAG+Rr1uRVtJLcbMRZIYrXMED4xYD2m3oSCy6r
GC2cr+b0MLo1Opo5FdzHdWzLxfupvdLXXuDV3nODbEiLFpz2h4kvbRoDYZN5tb44
gAEckaAPhGHhJnqU43L/5wCGZpbWBvuWz9NhdtH7iOlCNvmRyLDwLLy3TW3jgUiv
hBvLn9SK0yqV7FV7r5uYYro+0lhR0QsVB8SMNCced4WSlp2f/qNjb3xXlcP1qZxY
OO9sgMeLR1acsVAK/rXU2Sy6/MHomrMhhKOwU+nanMaAKfkAlS5hCvcw/zqWfz6V
37XQalrPrXyXREHvJT3+SHSM0GWuULx0d4q/o+IUXGvQQozx32WxeOA6/2eNA3tz
4YXnVHOeIgJ2i6JbBMAY8iuQjeKafUXxGgAJ4ZW4TDESUwz5+seOa3LdhGDOxQql
SA6LXyJIw9Ge/zan9uI2dWammPAm3I6+3rElGRlRDpBXqNenoA190JDU9GrRBDIM
MMPeeZJfYCwBT+O8cDWDGPwjxzDgrzOJ5uYXXSFcHTmv1yRfHD7Hbb3lwQ00Ukrd
4bjIxKWlMlU9HzFgGrjXSEULIrVR2enNlhunkSScoZG3EJbXi/DoD/+g4McUdpLx
fif4jKwigVuxlIaZopDvKP9K+BAax7osae4LDbbGpeCtNgHwES7bI2QLwxQlea1W
I2KTkCQm8VSBveGLvp7DYbGoFarQ5YMTaRJNdd5YyLCR/bJI+JYCdtSCbesL4vaE
rsA6qfPS8q2Z0raM8PBl1AzGPU1GgvIuX6RTh8yNsL1oq2n/xq0AKEpdBiFMxzAc
AKaHkli7379exDtv3TI1evvkKJVe6sbd+gZ+kE7mNKxsdvZjWDpXuuwk7bkK7E2U
HDIT9ls8Bp2K1yO7qPP0UawFE1+xbfo00vPPq0IAP8uXhTHuH5hcrqrqSDoL4bnG
LZoxLiVIFh/u5BMzidLGXe829ixQa1WKDb/VsmaXemjIWpN36AaYRNRLDmtWQhGM
zFRGWfoLMJoSGMh9a5F2wJbRc0HBrq9luyvZ3LlNjdNqLv0Epjiw1CbaqnmR4M5f
SC51syPcq4191A43aJe7hld53rJNgUua0Ix1sntOthF6w9w2SLS3vDAML0Mah5tK
+zOb+nZIQF1Rv2T6FXixoCVtjX5Xv4gJ0yEpTffKINkd3r6oXVdM1VmyEO5VNm9f
RT5hQ+sK4jDUSL9h6l7vAlysgZQlhxSQSgbiQKb/zF5PbrMzIHCp2zplB1aJihkU
Yeku/6EWgV7EmBCq5HJjYppT8u3x3mGVNe5oBeUDjWkpfbt8MUe7JR012bL2u7Vn
RRsak+XQ+sz7UUvCM/Bwapdq/b1g2zNFT4SyVh9KiLmFbtQ/0MqK0L8SVIBy5ndB
998xoZ3Tq0YsOYByBm565W2vmytSyGRA/F9VgA/1UYVnHlVv0YlQ8xPA097qccNO
DytaEkSobdlTQemDrig8c3IPOKNkudm1XU6xngYy5O1coWHNoFlb2cIFL8a/20xm
rICWBqosV+JSUN16SAtDcjF+F6NtL33RbBhrvd2dgqlYH41de5zsOZZbi4ja6pdJ
A6cvErc5A/ngi4xJJ+DkKZdqxt+BNnLLAsFqZDgx4AlMlMznZC3NGsRBGIwtMmlw
8YDaJNOwN0CP0zOT+ayGLRiD9b7RWDVhoyFN3G150dpB8MHe0HYwNCDnsIiFZVdX
coDt8Fzn3yq1aZOcArc+m/47XO/J5mgw1D77ZW10pqOgDv7eF39NeL/oq/RLjyML
B7ICrLUjF3vxWEuwA6XmHQTR1C1/yOVv/zR+tDqcOR3eWxHRMZLztvZ4S1HhHBG4
SvHEHAlsfKzXwBhkYwkRtDauJznt+RDiH0kSnDfK8RKo6AyycBMbRDAECih4Mkbo
sgy3IRqaQvlskFz5cm7G+Ms/mV4qKYnsw5zWhWCInm+3j06EzVjJSIjYqakk0Krw
Erhf+xYixn0S37VrLMQPvC8WuyS/4Og5YmuAUd4hrV22CFzNe8XO2uM9uaZwoGy5
Wsxwh1rfb9/a2Yo+We3cALScAyyVqZ4AN13vFuKVkyHQb6Oo6fGxJ9760XqJdWet
NAIeGOJi0oFRq0riPmb3H17Tk7TSuhxdcMHLTFd5K39Mh/7nmPZ+mh0zlmJfvRUd
6t+jkt/HhbIBvgnVBOoqvyG8VMJCUThQc9w96IwdfHlBZrjZ0ChCNaawkIxGxFjO
hJJTtJHnheVTBfwtV1pWqyt8nWEDfGyB34vOdJ9lrh5sFLt5t2phRyW4IGHudZOJ
1cIaKvZQqizAgVgO4d6qUbezJnjRqXGVK85CrTmZXsnKE/HtKA9qYxCAhfyuo3i+
q4smpy5Sg+gYQWIZeBWj2e3tZsW3Ctb8lif988X98M/iNm716ndp28R2zAhIWnAS
0uXtLIC3tKFqp769D83Jgj9/zqsfweBM7WzCxOK93j4wIvzfGE4i2lohKZeAK/Ww
U+l32LVjgtOYTjAcV1GlKw+0MVWDOGIdsP5kikZGK6JC61PoEUJGAvpZtH02ANdj
QIYiD6oQAWOXZifg1p+kFO4bE8TuOdgBTxC3DHI5A8ThyWIMYQzEc8J9cfpFkWAc
oCajjq/hmwyxRfdjMC6dITmajCyxoVZdLQT/2l+Q1YNZZC5naSUN0bBFbPJkplGW
JmIMzTkndgVSRIap4s5OzRJnvgrlXSbkMa1TkulK4S2I2hFqDmO/HUakpAa3k83f
PRNQbH/AzpUE3NYq1awNfACzNo7u8m6dUouwLQFNm28UYJeSoalHe7msYc87AB/Q
8y6wvVJ3MD4IuAey706cm8roR7GYOmVK1nem6BAVezUAptkTYW3Gc9uGUmR9ySNJ
pbbL4mM8JBeMHwst3SN+hJlbTQ4EhFEcTYPTgD5QHxxWKMWXO46Is/IcF3oWcWRD
BOPN7xHQ3yU0RiTq2tfh+cOFVF8t7wM9IS4h+l8CGhheHHV578f9GCrRwLgS0aEH
6wuGNYjUpPLoeB2Vqt7pDWiT0dcRfBbfxtOYDBvXXWsEq0RuK2/C3gIMFeK8lp//
OqxT+PfDEjO5eZ4FNBKLUWJNcUUp139BD8KNaDZfpC3394ryE8bHuUTKliUbzR2d
J85VETrqC1O8MCtg8syNa8Tl8typzEIYUSdStBZp+sZ9qfB6LXo+qlji8wMyo9gL
/zKaZbRDUTvZqDe4H/x7trsGcw2SpYETEhShG7k1DRtWAoZnvCrLQtAV2ELELzmO
OSPcyV3vOlRjRBldGwq9S1pnYjgApRhVAmj7+fKLJw6Uh7LUQQ5qjSQadmRAkZlJ
gJW3pZSFzKpzmahhKkm3UKX34lE+1VQm9oakvx97fn5TUo0ldCCsp0Hxc6uFNpfr
E1jTrZLKNlwm8B5tt2Gv1D9h6d106Xqyqc7qc05Z8iWPzbPKaZSaH0ozF41IinF0
WPJcjm4OGmE7oZGl15TyGUlsr7DEiYnaZ6XMBk91B0kYExHIJnAxFu7NABw3nTDL
SDRHFBbMu0ik6BZ01+4W+TgRDQBuhXkvChfQNEWpGZvrSTIqZL9JceTIJQR/HwVK
JocpzJOXxedzzTFj7HJnqIkw8B+y6i5thhVvsxseWKzZCHQXBgAcsoMdFKcq9Rxj
Gyo4bnaswKZUHw2ZN/vx3n43wrX7vKcX+5bgEredfl+x4lyz40xn5IeqDVOE1GBp
2nOQO+Cgz70icghMFYsUhJFbiKztxPpXM8Fuc/zaVrfcYSCV3iBdFqPjpuAa8+6X
AGuo/HYo1k7rL/vM/y7gOArwxhCCEBtrstq0HQk928sr/Laix4ph5fzFzkeSQzXR
PqkIACmLYnl2sNCsY5rN4wdPDSijGa34X5+DcugydU5CJNsgCdm24QMy4v/2OD5R
Vlea6hRB9t/A+MSC2sOTy+mfEziXi8JZGkB2CgSli6BxRvtzqeI1BwJl8W7+PWwx
oSIh8VmJoCfFmjZqIsYwUWuI9BnY3wYuDK5YCMlv4s+RVjvpqTLlr9UTsZFUhTMt
uLkQ4N42MjdAvdr+9xWVvDgdVTl+JVhnC63h7eQsnFPFaJIB3MZUAHPvqTQZ6gH2
moe2zQlwzpok/9531okqzAn9YqI7oqg6dgC9NYtrIVm8SE3k1R28dZVs1+O4G3gR
98KXMZQsZdxKr9/KOmnxx+IjtVJ5aDw9yLPZLUkbSNSlIQLS9oAc5pL52CCQjmw5
XDZyGwkvUILda27dCh7nDc2ZV+EsfceBgVOnxex3D3IjNAYpG1pB9qBAMNuZnyoQ
ObubEoJcRT01Q3p8mGXbsaJNp5MzfF9ou0aXcxITgKITa97gyD8Xp5zRE/u7CLFG
5fNpubC8fDYI7mnH9sVKAOhyrnCSsWS8SOKeZ2naEXyd0zJyIKxSZPNaum8c5sx4
aTb4O757Ac658r3LRNi+HaS7Fp0ldBKgy5OVphoPmYzeQYNKaFQXv8JkIt+5CNml
1+eYqev+Vq/OaxZ7QoKhwfKi+kxgosJE2/D/mRuAKA/9rIcLZskMTBcZI/3JTojq
ev93ZZaw1QPbF7cCl5uId4CAMoktG4aToHx3WFmcFl7MIpTpkjGSE4y1yeczEGeS
z32njHT3gqscWoO99MaKxcF/04tT7UPNxwc59Xu1TBHQInldwF0qxuPPpGCcAbz5
39B9Gv4YR7UHUmFnTCU39Fflep4XQsssyp9MC664hDz+BTVoTZXFb2325whWfgXK
xNeWt2bC7C0osJcP7vdQJcMDsOsq529KcRUscSqWMDtvOFstKRAyu/D4oWATlYdo
ImaPlLEi+cEL8IMNQqVbV3H52/pZAYDI94kRTiOj/9mvVHfqmlLb0jtTZ5rSQmV6
2IsLlFDYHVYb+CTa2W5noZuM9hALqxrqCCvO7MN1RkZCWWcQOiXIfqSZ+9yeqVOt
z4T++C01G+6RqG8dXH1FDokEWzCNXj54L7ZSe4KQcEo+2XZqM7aCQ6Ee6yGcEbmf
3+IBV20h/R+DCki0fET6U29p2vqz2MMV5GaVrEs2EsWVhmgsv41e9szqEcnFSc+C
a2YOfAeNJ+ZoYkp74e/WW+4eEsmOCfPIBuDJZO6aQZsa3nofU0Hd4Q9x6SDWyZc5
54iSEFd9pKkyW4qR7xBBrL8dY5Pwn7cnPU1XY50/oMeFKan8EM7Wr/o6y8H0PEd1
m7NPYAsJnc1kHh7um9tHyYdoM5RjS3aro7LQfR0fGFO8BFPcksAG6alWhzvEBeMc
rATwbAkGV3ekTLVta/C8cuiQJ9agGqJDchHK7oA76jn5s2MuyMdi+hWigEh7fwVN
m+etdA6bs2VrPpzmRm9oV7nIO/zif69nnqCJ2SVQI16CZdxotCcpLk32udS3U2/8
zTtjqLd8T0GzooH4FYLEzIC3PPF0dCUpmQ+vQHotCilGjIfkzu72djygapqFrPvE
f4Vsu7BMAND3sXv18quxEeBQXVRTm7a6J4EPCgT4bAG1GGPPBAQ6LLj5h8HJn+rL
/Shdlz/ol0PRdcM4ESpmAzxAWB2V4SyeTGIg6bbq/wIrEwGCsz6If+LEpF/hEm3E
P+GbuaF3q5LDRpr40UcWWepptkXa3SHzUH+puIi2TjBHCZzWZYBpxXzd/JcC22Rr
f/58QuFPv5rGqvLgjQy5KXyR/2wPkrOhkiHzgwZeFL7K0EnFKmMi0fKzi2arOq0t
P8F1rVK03ShMlZ96wPehvQ7Xz2DnQmvC4AuwBMlC14UxjG/wps0GHmistHLUS/g4
KtgSFcydr1yA3pa5Io4OYWMAilUB0MMEIy5Pbc840e+7TzWhaUfOIzZiQsR2mnwB
Sp/frT/kGFRC91PWQJKeCPFXfJs6chZF+DQ1TkB6F1M9Vi/JH9pm41Gn8t/QMAdc
qHVeZ719a12v6pZ4ORsOphj1VkD2LEvskYlPV7GVamVWfMNnrDiGeBdOvZ7ueub/
eAY/+qgHlabJ0/POHgKZetNHszB942rEnQuJUcmrtjMmEfvyHey8d3551RKxIjps
OEaWF1nn0Lk6jpFtABPf2QRZlHbh7+fVt7sbZQ6XwreOEpTIeUNWwu8I8wwgQV9x
pGKbhey3NStbN3HLJRjmYgcTC4oMo7zRQ1nYRsSR1e0P/Kw0omR1xxb9GuwYDsgl
VVRm1yRcyHZkSjGYoeHCvQJWCgPNHtVQs1T3M6T1QhIWQpogo8wftCzCOei75tyj
QHUOyNhKICUVMZFqMozHjGJNEDTILV3nOYB6WsrLXxxAvCcJFUNlYffmeJiIPTDh
4pmLOTRJrkCGidPQvPglhEAFK55apIcphYtkTtKq48qDqgcZr0QB9ga2EtPfhSVC
r4Rc/14YYwLaw2GDtXIZEIGebfSpMYoiQYdPetIWleltAi8n/x3B/1sAdgnZj3Nf
VXXgDl1h6JWyx4QVgGD+o6qCYbhGooUsp4ILmCF/wBM20MdZ7xY3nLM864+nE2DJ
NDIb6ee6r2IeRlj4oSt7L72sIGMOVfc8hUpyJ8nTr+ku0cVRnGRN/QsnawThoK2c
3CqV6YQJPAJxAcDNgG5utvV9k0H5Aj99znwYY0qmW3QkxHW/NfyLDM9lptHbborE
11aX9gy4ui05JQsutBv58EAchlEX36i6J94t0wyKWoSHivS+exAVNxfq2riFbkUM
yNMQZBuwVl1ZTdNFTC/pdh8rELwY8URnhgFFqNBexHnJ3iVu7WQWfx2czaZWDk2I
xvE5G3I73557YdcVKn9lNqvXO01o4jrS0SbbdtPQWn5vTMs425UHGI0xJyG1NUra
DzuOOcdiCQkwuMq+YCFc4t9z0x1kPLHwu/cHEfQfGOcIV7lkf2x8iiQp2Z+DHR5S
/+TLtALA+bQure1enyRaeEucY8UgdzMIBjf6mTDh+5CjATxDT/iQ3FiCMBXYBFQE
SHyR47TebZVX8hjvvJtljmhGA+lb0MasyzjASzkdgUv+tFlslsjpWECM4WAvtf1P
G2EgNrC4EuAySz0KOfopeUD4zC+2lz2O3eJmcvKiufl+G1Or58xwc23RqDxqjE9A
zZyA3NS8XDq/iaTWlIHol2tCcWcWF4g9EIoXntid+5B7gWIcNma1WENRtiNVTt/y
6magBvf9XeGoYJp7K/cXNHs0IjjI2Xxz7FnRbmrTesE9JXOamO7v4AaXv8o+m6Vg
IXj/5/uYbJMy01QM7exX6idoPMeUyW5dVKb2qcxG/LjlTb81Zv3ntoaM542/0QUl
SKx2XrsR62WDLZQ/qiw1I5eK9lonHTe9QfYcud2uT4K3WBaUSK0Fy5+k0BS3lsAD
h7BMQ+8zkpTS80vRR8bI3tV3Y08lWIR5SGNNS5P0OJnfEE+KwW0IuCw8HvgLnfS+
NnYmwd0dISCmBVQxij30hXXtzllz4qXJym2FApUTbivzD963yLfvfFgzEDg9DwQC
sIqw0J9D1Gud26qRx1M+X8wT4PPMLcSn8cIQw6Euj+A/qgRahnSk5jHNKlxb6w4W
RpD6OySORLiqQ1FyYs6BW1Ln4HDnzmjR7VXJH2jqy02+KjYCaL0j/m5nA4I9KJqc
XhVMa6AJ5E+30lDm6JKs8Uq4+NvO75crBLFQJBTEKgK0xcbp7r6sYdWhb0/GhY0m
QYUA2vLrz8Yno5NDFBwBI49bdlr3dieui1DHP9k6LzRDN5Nt4oA9/f3gB+MhmYEC
+OhPmAQK+khCLr5PuLr0vQUWc5g/bhvQ75BuLAlPujWHmArfIgi8BDefQ5q2bi2h
7C69/eo6PAkZ1uMrYYnOBYGa5IqBdWGeCCFow1bZptaWsG2SmN2g7/YvbNozVJZR
XZL+Qr2j6/QK7lAdvTKkbkUIIl8mvbXQ4/Uu+UMBr5bkKj2Xrqj04GnLmfs/XmDc
SaqQfHi+/ugDaU1g4a63S7l1Je/Uuc35WrOyjtpLgfcNfse42Q25ZEcarwGlTIKU
KLXb4SVRi5c/4j6d57R1l+EPsjX+Xb1vwKu4sPwdueFfVL4G5gR6munhQWbuvab3
L3IpSw1wVY2FmK8Ei961fN/vaBx26przOoOCCHdz6GTLjybMZ+wQgxUa1z3WUU4q
m4vefxP1GvicyItbb/EsXB8FxS3u6E84fKIgyda2vGyFapX6GBtEQfCM++XkWo+O
T+QrjDu/spZ/6g1e59qdAGE73n6b0vdiKUY0TJ3LWoBF5LveFbfd40q2n9bxiima
JeRSyAm97LXDMXR8cFFyUAhKzA4kpM4gWer9l45z4NC58ITojNDFq+flcT2tm3mJ
7ynId7uYGfV91pzSBfCSDEpcgwVZ9aVL+H2xsemZ2POoUpR76DjATAd1YN99zHYW
BQ8fnFzXUj0eOeKQOahRlPphPoL03vZyktMiduXfRleJMKZwzParBIk31k0rGSPo
er+FbG9pT3RL6XDSLaQz1tx9iZmiAIbooXr5ekdGJ56909vUwVGn2mrzjswbWmJu
UtLDCX6rJzEDVYqHjQDiA1vyiewsnuFD6YeEztIZNd2z79DAGVyj6S7NqP9GHT8U
Vfp7AqRbX4y4pYt9mczUwkoDTRITBbC51VoDqaRLMMU2Gx3Kg5wdgdzE/bJwf3Qg
9Pdr9rrgUeht+doRw/IiRp29J6fycmvI5zo34ZjHvNCu2+GxJjzb1zIOIMy1hWPV
zT2dvIPwdX/ffaF+fxZLMhgNw8gkOZmXCKRnzXmQ9cBOeaVdsqVICnKVHRHTmoTw
XM8ulzrHq304gYZQTvnqGz4CHrBxLSfSDKEX/HItsuO8RUFwzP4VdGffxieNURjs
0EVURJ7pyHxE9ZA1HO/ASNpAs+SrY10UuHShV+Z8oQjfeC9a9y/1W1tX8Dk7aUL2
p+Hoap4OOgPpbMb6ZiHvWk4SVi09XPeQdhMAr7uBU3+hR2uiTZe1ixbbrllM0zKi
7YqQcciUypc05o2sKqRpCThdju5NZnmtzpdUhYG4X5KD1YIeouLTDVbGloICtYfP
SSPTk/ytcMHO5XEdYo5dvMPXde1PGV0TqUREArPG/TC4bYiwHdXHMJQUxRKZYROb
a7vlJzf2srBqSB5v0tQFMxykFSPdDeeoA6xRMu5YssELXLHFCGISTI296TnFmjz6
W3EPDDPxF6hMwRxPbXiZZ2A7F9mwpnJjHTIQhIL34FQ83ILv6uS7DVS9HGIEoz3t
hd5qxg/AJ7ZKv3GxmcrXbLoAp/r7i5JhsiZnuxMbUHKKaoNwl5hm2W4gjAKBDl9P
j0HtoFQTvbBc3n3bEtx5kyzOWDZANWVtjqvOftyGjA+sPpPdWDpCR1CHJphrXTDG
jJ19yebWmfRlU2c/oyCe2NfsP4WoIZ+Px4r5l37DXBI8ToMSqknsvwyFNMmgXxiN
4e51YIDf/Uwxvz0unbm/tiPLfv9bkUyJyvE4HyWGkfBhFCKPYizVzdboYBREZhsw
yZLxwiCthvmKpYlUZ6I8jyEiAaNjXx1lDhipalO+gZk9++rP8QaNPFMn4DoU3FfR
0Ut2Kmx/Tih+BSsmNrXNT1ea/tGXPSs3whGX4SwAmCiAERABF2RI5cTuqlqGdxul
5XgtQzCK40g/afuO0aw0z+rlVCDnjv7Lcr2+XDC078L5v0xHdpWVSb3HMpVAcDBv
EwdqNcqGBgNJyFRZZSAc2DP8Vy4Qza1fCSJ3XPPwY8wasmcx+tWDub8nSVl8FY6i
SCwZZdOXRHKIYVwALX1kGAjZGvEKYBkuejGqFfTlLJB2i5K07ifP0HP1GUAewDyW
opB62023Rhw5Q9HZUDU65sd0imwrqYfGFLdk5KGrv9T0Ee0Up2OR+m0wFE+CTJPs
IqZiGS5uyhONu6pa9ijau4Iscw6iAWQY5I5l5wcGZaw/c1s+LNb4rUwZ7z4vJx9D
EJUaeVlX5EKdslPAyZ+yNz0vR/TQ3LQIWYO1rt8wVUqQny9PYv7mdlRzx12G6+fA
k580hfWOsFZVPEKwGjLkUzOCIHOarI45DvscnnT7rcB24yuuUC1Be+3NnPGYI09/
OwvFOvSgfHaTm4cfdOIUKQQkViohKi52nnUZ8C2yASXfnr74J040Kb9TzAEcalbj
i8M+h7wXpZ/ZS+jY16odQvBNeR/nrkuoFF6g75oD/MHM1TPExE/PrDZG8wAxaK8K
HfwxeOse1ArUZm4uGmWtFRoFEifPFZMdWC/2HVGMHlF3M4/QTu96oSkDFbOt+kjV
v9KlnrT2lVRf3b/EvhHq5waentCeHxLMFnn/0dZOekSE/t01g82FXVY8M8MKAiR9
oYWUlfsVaA93jsmmzkVe/jghItcBGLvyLQK86KbU4ZZ6Mk2Ogn4+KyQn7UhBDqax
W5BP+12pT1Wjy5v+0Xraok5Vq5MbS3lAMJwZbghqMwSnpjcyo8k3n+feLWA8RsmR
mfEQU+17+dLYJls6SwhjFN8rvAwhw0e33FejGIBZ33ziAhwR0VqsWl6H4884pbN4
G+TW73Dou+a+8Zuwa+Ra2ohmGUY4tbUO4r1zXdgj6ec0bYDDe6ZXEKPd9pikD/QK
3wpE6or2he9WBgbaRyaUGVpfl7ve/4VcjdSXUAiLmBtnJ1eWa3iLB6mSVmr5fvhb
k+K2D5Qj7PvTzaH18bWLisLEOYTl2RmGKwb2BmZ/ghtvUwYP5avrudBnvuBrm1Sv
PQLH9NSjY+c5gWBPXi8pniKKck1dm38SAlj5n1vq73pd2vBifsqMV29NrTv8Pvg2
ekjFGvKirPphDnl2G62jtvNUYGwKa6UAyx4OaQWLKoWI1C7izQ1HW0mCf2I7NwtP
0k6BEE4d+WxqlUsr73oQjNij9LgUa5YViZuJ4u5AxecoVZ6BHmoqlUPFIjGfd9G0
3Z4tqgM69QDY81r9/dvPWL78Rc8sIwKY3mFtx97gOwK7MsGoprI7YElmt/ypd3ha
Ny62/aHKdff34JYmaG5ieNxFLctF3qoTJUMVylJtPOeloRqWnYfmnWlxiYkumqv8
4RE7twtvvliQMqHW57nwHqEip3iewE8rrpWxcZnXcFdxi/KuPwts9DQGIeYpe7IV
OIwYSefF0XAFlrg+OamcCTHm5QJ209Vn6EXFBaUVV/H8NXhOzkKKedblp8XQmtb+
Ve0ThCSpPFe0gdPSGawZxJy10ZgwZ5dtU1XVmIZZpV3dD7bbE3EHKySvXDpNKacO
q6qwK3lr538sV/+p2U9KjxzJekwNtBoY/eDPSPpak9kFpGmNhlvyxpSNZoqx4WvA
sRiccP0Gqu48wFX+vBRUM2n1NDErM4M6PsrHkUCZLLvRidQOT53MDJHdJIASbfeg
Zo0fMcRFBmKF0HsLQzB47DEW9VewzM/Jp5WTyAwBJezhRVtfmuxEBI5hZyS26N2D
VhRNpPqBsgaaC8M+M9smqcleiaCgD/jpmpJs4O6cSN/hie/QDq1lkF8oHofUIJhN
phR98krTSU8bZQxnsqYGc8DPhO6IPqJsoURLeJuTQ2KMsYK8Jtro/yzV0XkiQ3fM
aFaIkCMzDkJ1kS+Yxk/8X196lsAoilk0F+um7Ler4bY97HQmcodDBWusWV6zLkPd
Z0WEIY4fP1XJiLMzTbiu0nwdeTUDtUl15a6auxAhOYcDFUv35BBAzwIoHiw60fbh
LaBG6m+wWvbqOoeVghOl2NcIVjBUDKxNdLae9vnH/+I34HRYBclpvW5XqL66aCuG
SwkLCnnYp1eGtxzMWCcKt6LviXuqrLXiYXHUQ8CRhsay/lKp+y72PeAaCxiA0NbS
k1uSTvjVWdDgH86olyYw8WvwbINZgqh/6s4ifURSLVDHeOKbH7LyHwZOeM7fTazk
XJKaOOsLIS2FQWPgaoa1YmY4LbLV1gFrZek0hbIX6FF6172rYA/Ui1kK7ARCFxfU
KLy6racu+RqoazoMlXCIYiuXQqHgptbcPwJZU000S9rpMlN5OXZjzKtbgMIRsOrR
PWH1eVJte4J3NKymp6cvItvWLgvpr4Q2vrb6Yur1YZfRRQan3199tq+oI8pPOxLn
u4e/PfalDM1oHEt0J4lUbuOpCL9otqDWHrT2ifyB7fGcJ6T0duJ70LPMgViN2mH2
dqP7//2jB7VpZzYcqfQPJWifTl7xy/bph4xvqH2Td1EJnwvCZIcSrhDF1U8RbiZh
ChUaYu8XsdigmE76sXAVu07IgPPdWzWo1j5l123x7ayzVaJiNQvRhlFg0EphP1US
8yCTahmRYKG9iO154Wh1/IAYD01iZJGlCiyph5dXhbuwG+rK4Obcp9Q9o3ohwmkQ
62ihorLvS9HQB7ZZNCFqa8eJYqfjtmqYE7A7TdSV9tv7tg/4MnFalV+jivHwhT+Y
DYoRKH3vIUQTFl6hweiEppWmTlVFZoNua8u23TTu/yVq/LT02Jwm2QTSNwGLxOt8
PGZM68KlMAFol7mGs6Ply1cBUz1fGv65mN+xZDe/FTJAe9j2vQacwxq56CXcSLZz
9PtFIpaCb3vP/H35XQbUsIgnBBinifVOHb6b0yzTQKFYtXH6Khw3dDavvSPENC6f
8gkHEdRfk/My2VgaqDT1Prevc/IhSI8JaaCvn7+DlzyUBuqu380nuP4M57vDpjkh
2pZ7+UsW5KHPCxA8M9rwTWC8/FCBTF1hX5CspZv1Qx1SapjfyvgFGGgIu/gEVfun
7TdYrLXv7YzJmmLiv5l/GEeBP+Y7o41S6qAwXUITSJJ5LH5EVZpfQjK7Kw04wl68
zXabpodRyg4dKuqtpGZXX28/keskT1YZDBDwI1lh5oyoojL21Gf+YcBDOQ74Kyck
MmfA0E8ivoiqpaKv7AioGn5rj+XBl2T/vYKm+F/aNsxtWfTS1ibKu9R9z22Np1Sf
3+M6+A/HlxocxQXbCnq296YFxLCNjyt/OY9kcE/7uwfkSp96jF2X7Q2doZUu8wjW
ug8Iqq+ANq6tjyECdWESJrK3KSDkKCMTI2vi3LwUWX4hKrfzNi32BKeknzuhuD7Z
TL4Qm3d0oZwqz+x8niOHCvNkralkC91bqN3LNDbxVitCsFNyRpXw56qOn/HFJ10L
JoUdfXcA5v6WgXUog71HfdjNt7wlCyrvxYO6aHkxvNRiGrYZw8D9C2HguBx6YHsg
qLiHkzxCA4NoTi4MFIk6F6UybKO4vL/+DMOl7OQ6ZhaPaNEgeDUXh8K/HGTVx1tr
uuajtT1H8YkVIW/LJO+hdNyK/6vglB8H0oupQTpZirmN+LCbeACMtmJEKeYVxktM
WOUlBkFugB2XqQGzk9Cpw6S/kS0Z+7AKUiI4JDZGz/+AU3Giyn59ZPqSmOBde/9V
jX2hlEjgH/O9nhPPiME25YPds6r3+AgtM+kGEnR2OAuLAMFOZ4QeYOSYVHI7n5/V
xxed0eD2c5HDibcyO/dsurD2U3DadJ2ZmPupmrwn3m2JNZimwGDthna/vX5jqp4Q
stMASVAHblLcu9/bHLL/agA/eC+yVHmECylYT20PtcOCdhK34VKB0VZZbaa6OBiK
cPHDexd4c8vdYA+nqS/ARW/3VXNMiupAvjy+L/5PF7+r2OhiS04oLl55MGC+eNSP
8iwsYSnVqjIzjll0/8FxTziki9JGgcvf0MDAryFVefIUYBcwQ2hA+NCMpafz4l+A
ozIF6eW7aMqKE8rEjRWQG88aM366GuIWcYh8rSNMHrscjeyz7gPAIE7l5DyAbSnw
N11hSJ5U8au2yikRZRJi8sL2M11Sv4n9mQt1YOiIf+Bgw5Xii/pItHlqcdmDTdZq
EAzvGp6EB2gXpgpf3tyepU12TN6TXOxgn/I7p96xcLH1poT/KcqJ2v7h4SchlD3q
0U3DqGh13clwUXE0sq4VxlYtlhIcrfk5sVyJ34ZGfMZmdb5oRDkPy79OlHHwZnJV
6cddwsOftLuahgevMX3SSdoxPlgStQ0Hr0qMHmMwxWgUWM9BhUP1cI81GFSeF5He
BCS+qYIrQgyyAhgLyjIR9VKTNWw4aepkunCDg1gWB+C+i2kovZOEui4iHHSlyU2+
/9BK97ktcrryub0wTa1nkfhzrTNyu5rHnM8k4+fA8k45a6W6HtkU30zWGfPSj7Tq
Ve4fUN+FWM1jdfns8aLcnx7ZBLaDNyHTPvvIBmzNbIQxkYPGxen4m/Qaq8YCL3hi
SucMiuM3QuBcZT6vaC4tN9zAQ/vpzVLbIU1L7BW2u2CuOSsicISEd2eTj49XmLHZ
iZnCC5ppfEUcEH+GkeJNtrc3LXHHB5uKe3Dmt/mXQZct54asAyKsXSM01zNLtzIJ
/Yv/jLgYxqKPh0WEUYpLKog+bW+7N83DJkqDn5+hgEx7HKS8yVUeq7RjiLqKmgID
vnUfs5O95L0e1ZNVlhrdQM9iBjkKpmmq8AMDKokqSOD4mNWdb2cgD3Rnx4mwTvHq
cCeMVTz8LPp1R3a33oEm+vmSIpyeNoA5/HJFPQIn7RXFOuDQW1CbPzZOcnZM8VMD
VluO3xvY0qgGVeNzCBtYRJ/Y76F8GWeGYNi4HdMs0Q19xfBKLl8rtKlcCDwk0LEt
X3MvZC29cIDyuzaBD4eq3RDSAqGRrhDr/sCr770XE00Yr6+ADCSlYOPgJeDb1NhI
AnX4a9zyCgnEK/CNr230Gf3FXqC6SZGpUt9nJD+Uw2wr/lJsx9Msi0vLEBJIP4o2
5MFc7ZkvZgl/w+Re+R+QCuDzIFXXojPMOqys0lRT1QiqBAW/pPKdhEYtwWV/2J3S
zTvckk47ezdVlaIKQ8CzIyWzF8HWBfRHVi3DFNQPfTtXgMSEmq70QSSYxH3hIOoS
QX6S137TbSvD5NhDtcTMbGY0JzWaOYLAAxVNZdSCB3Ndf7vwi5Rmu7aETKeiDS+e
d0jNx4EgI9Hlbf+0gRWNcFSwTaIFRge5ZSqp0CdEt9TQBrx6A4M2gNkwLKcJuTOI
THjk4hKIGXs01AzeFOMMBpZpaGIhqSZbLz95GhaR1QCGnYFOPrTztslo8KDFKMWU
mcc8lMAWgKW0Ra0vlYLCQuM7Lk3tzQjP03i2catE4iLj/FqE4w5yFSgULxQW0ULh
5bqppU1C4s6qzjwToL31eGhN61hoGVuq8ZLBUiwPIxTm4/2mutGruRilyfX4QHZJ
LiHOE73rEGqu0IWdA4FfF+5HLOPoziVfmBljlru8vMgWsUGXOMAOD1a8mmDxTVBP
J/TKhJ3AYWsC0RUIKOx8Rw4nTuiIF2nQOidnlMiHWbfLwr7PxxzvH6Nsywk7qRA9
be0DoYth0KnxeJf7FaKXDo4EDj6WDThx0r1D8CgL0n8GFJ5YmqG89TlixKk6kTA4
7eFB4HT5Ho4y7PmATDk4Eqvn8Q9q4v8KG+YXEIjfcrQvSQ1Ujw3dH0tSb/mwv2P7
hyEt+LnQlmez1iXrs5o0N43ZTqz324UeJdJGDlAb7rN/sf/IV3lOfLJlSFs0s4xQ
NrmgIoKmbFsUKUCCBy0AuD3mC2y8m+1+xgqOzmk+ZyqMeYkftkIj+BupS07yYq4T
R2IDGnlNBwHxsLrD+EcKrGaYhwEZO85G6h096KUGEvXxJnGBOPeImCOhETH2kMQh
QNPHFmjMqnHeB8K+lwx/fj+WIjyVvLoJYPynRgopw7vYZqbxddaO3RwzyL0uKJci
oUYOfM+nm9/GWh7MM1kFAvfExrZ+8vfjSkLHFo5ER4p9JgI1O2BZShhPbDECZiYm
WoQ7j2AWSYGrlK1gNJpt4q0KfwZm0FOcMVlDERm6ipxCDpXWvQ1aJc47yjGHWXdo
EuOpU7j/jQHUlgVVh4pVaBgmvbbIvUiXT/8UmCdX8HAbw0zmwC9mOuAK+fMP+/z6
NGBya4BUgy59uhHr1vaDyKvhZIMDwuEjNcNzv6MUqGDby2YBsxQYOAzSCL9P1odl
YUUarbx05avO89FtHABheRuqjqSH/FSx5vOfd71RNGJopawSGMdB9Jl95EAdNDCp
4qIQUwWoZno6Ny8tag064NRUDapVDfV+LD7ChQbujMseEN7WNWz+DkA7QpdB9wQj
0mLyGlJx+E8RAGGghSTD0xMk3IKQ/HkfVKTugfiFSaEJLu4DVfTuExwPIUkL38JV
V6KdhnikRu/wHhECbZ9PrJLUTnon4u3vFJw+nMzZwQg+p4zAfJJ7HsBEd5rds+6S
RDXte5+KFdogSMv2dkgkQo1WP5063YOOwlriHr43jlM5vJsVGqmDOUxGAq0kweJd
zGyoQVaobJGXITuO7sgfR7D9gmFELszbO5+9b1mSWNhsWIBZ+NvEz+nkooxx1bzv
Wt0277e9CRVl5EdkJDwImm4eocIcsAaq2qhdSvZg13sA/fId3tZVT3PlxPFr7PMf
2tTx3hWcwDWLRTb1ZPkoDTGssT6tNtKj01dhOTz709B26Zp7fUhNgU4IUBe4feZM
4N8uTd6susi7FUvVumrD+Ad/cPLnGZ6ZRH9Y0s/xCV0qiMrKQI965Bux5779WO0f
AOaIpPBfgdW1aysEjJSANXj0UNOImbwm3V9XDfIRIcRdcdbV3TFBiqPwFRxWRLQR
19T4BWs9E0dTsy7nk/H0nyYrUG5j+hwJlsQWxpUKDlz9i3sZRrs5zMQlO82uQuYv
1xAEl2KKDRccrAFLyuAvT5DO7Qxyfi4YNmoZIAgiU0H4zsiKvwyoCFeBGHyW+xkr
xVnJHcp4Ix/VIpOoAJaZT9vd/bPNwuA7zSqNJt9Yr/87tEGtc7DqsW+Y0vEWxHsA
BOYIqXA0X4MjUJTxKeXf6XeinTUFMTcMvIJbdzWrFiDFDjymJ6pqaJAWJHqNBdOe
TsZJezvbHj/KEn3cEvCXFENTe6JAKVXC+0EsFZfqqhdSijp2q/NdTHwazSzgx7Uq
6FwCXrKfzX5lDnMaB2yjAA4PnECb/oCH/RmmCsfo2UKGWkVdETtWqpX+gBo7ID5b
I+eYFQIwurPNxX/bD0PbNGb/hcgkEzi5oalh3aZMDDEJEWqPaJ2q317XPxFtd08k
61zgjQyhIHNj4je/J6MtTP+/N4bEnBHOCG48cyXkwqQNnYJD8VV2xOjN93uolq7l
zudEk0DIyW2R1vgQmMjDo/aSfXKARDdBi0eAGREcfLorWnAHx1Aqe8PDIjLufnbJ
56yBhjjL4aeCBb2+HJdOaLFNSNH4m6WeBxlSIIb1EdYja0puwP8d6dKMlbLOjbOs
JQKS8nVRKqH2cL5V35k72NjaT+rIFZgZvtU4iFwGXWQrqE9271kBBqfDZ/YPJZHH
D3sGm1Zq1iz+1hsNW5oUmxvSUC5Xbrmartr7hUyVasFGW10osgmT5sB1SkZw8POj
MIt1dLaDeVntCu4LC3QzgTVwyj6//KIdL4ZKD3LjuH7AaPaxHEXW2SE70MuGVf8L
y+JsksuofkoqZfHQKtmbBX9htWLLaVcRbINnY9CGzzR9QfiZH5OjTjOpkhOnaVex
SwB3Mg4Zzy+8H3Ppl4DLIknhJOff+e1meIRJ1H1f9ij+nd0sRuSvBjB+AmpMsyu/
EcSEIPleiPkVI0yV0909xCDTvJU2wruRtaG1VkJoWdXbu4IYsu8pPqkQjXvBdctY
+E2GuRk2O6OxZKNAp03KZ4UBFVQzg+O6ZGuy7uhySolO2Rv/T/WMJ6oS4sjV2Qby
B3a07ps1SxEZnZNyltZKqgJkWLHa6aVFH8A9dxNeNiCUy4FGtDSkaJ82O3iVlrfV
w+55VspkKwNs+eHIx8PSIevbs/JBm6rT9GPlsbc91D50LzSl9IHsKkqDbMp32pHM
6HU4zs5qlnG64kPWUj0QslyYETjb66icskub0rwRJJzNM9DyLBVq4pkAyznxoWlm
aJFwaNfYXMyafsK5ejeLZ0LdGadMVZelaRfWWSfZ0zSKeqOySMvZ0CLotQJ5/il9
jqsbCJunvJXtPAY8QxiZClaDOy+PArYufhtl5fTW2KHM2qUe9b9nKc9FxgQJi8oO
NDPC/JqOcp0ngzDg+kIWafVPRN4Ga9ob8U9fEYvKcwLRdReI0VfNUYDTCz4HCbCG
y6nx5zqturZaL/lTXBu4mV+UrEFvFbn5BaoBxC+VQZ1xkQu+Tl3c6wqJlBd8G1nc
QqLCSpB4SAaPxnKSmIm+oIF4UbpWHzcZXg49f4cv9HBOR+2mS0cYijGxLu8geShQ
tqPXXF0aedAWpswc24HLQqKAyPLf6UxIVR1lfY2LSHq/10LJkZNmA8VvINFMBADU
1iDRzIXH8OybREG+5dUe4tzi7JWhQiAmeNsVrG38mU+mj2oPrzfGiN3EOSqdSiF0
b/wXEXJ2ixkUQHJfPXIYw597r/meF4o0JOd3SxhYBcSMTd0KMzwfkjH67O/hq556
NJAbc+o7k5GBgJqjNTxZDVk/3P2vho0pQO6EPtmjHVf6U6JN2MybUTz1UIv6rSWp
jaRH1BTGCOfKnYT/CACx9gbJFxpsJhO4G0gQTXr51IIjR7R5PIwS8ulEHft1a/Ns
/sEMeh1NLK4VisX+4wn7LIL2hg7/NK0/rT4R3cGCi5qKAW848+9TLo1lNs9rSedX
LzmaNX77013bqD4ZdXHP/8vZT2wDtg5PMsyI6WRajRFDojd6pv0NaLolldeNUuZb
2iZYiXqDFkOwHUqsfYGUP1/dR/UVOoG90KoDStaHW8e+UX+Oo9cHlpDc/fPIlVbd
/WPDV2TKP9wCm85jyeJicRX5RljHuQUztDptHsWIcf0WgLbY9eJIlW3WBfQ2mMov
JdwRHkEf4qHRGQet8y0pDKGOI0KqohEiJ+RmSBEhsFWdQ7ATVdlyaiHr7uAPLD54
DkGzWWkH3zNTynNN585Wv55lnerKeLoalHzGH2ow7NPk6sdq7X/Jbd55VfVYqSCq
iRbAKIztlkDfssNxrzlzl4WNI23RtnIjKUp1bjwQNQw/L2rvHkLzCOY+Jtztzfge
FwKRXQrxKULOaBLd8atsYJnxNQIt3FIpKjTiBKtVs7ONl//whEnCCPaKYRbuNsHP
E0+V86tQgC6KLzQNtKWB+zBPB2RsKJHyRwJCAQSTZ7eM6c+yk+faBXldI36Ylj04
nKUSRrmnfPxFAD6QhjH6w+B9BoPaHu8Y53/lMV8LOgE/7gJx4cszw389Y+hzcP8t
faiUddQlqLUEmFdMueIecE2a+Y5MzRk1+x4rlIzAA0Jj1xWaqc07dTx7StZ95joZ
ehShC/QkMbjatmQYdkXskWv3Ex1j/kU0phPY1s5+e1meYx1Q48Aawg073F6Ytnrp
Et5A+z96ohFKCJRLRJusdPvVJO/PqBnctDfmqIaoOJNIOF1gyFcoPam/urP4wB56
8jUCy7247mPIQ3BflxukDsXb41qERHn2adGCMAyvRnGKmiBcVYdOMssCHg1Sj1hO
t4vn4R61pKwSvCLVAtKS+9pAHfAvIDZIPthkmQo6W+FKe3T1sg3NAotaG3H2MNZS
M+n6STXBYn4XfjY8O86whMbLIBk6lYJc17U37k/qekt1KXMLIVggV13f6yeglaUf
oKzPx5GiyL+68WCMjXTC4iZ8Yt8dPbl5yopUSG5C04Zg3EcCPn0sk1Jda2dmVkLR
Ma91yqyLoLtWBOgnegC9s5Iwixpf7BHOUp8qXQs10LYebATPlouzMIUqPqduEvXH
PI2S54F5bh0zPm0hINlsDtfAQb7iRRky9j9mm55FogXPIqpm3bMdtqqdzVG5rIvy
cmJUPA3vlpowazBFaCfH21iupJ1e1XvKJD5eYwpipASA7m1dxSRWu0JKCw3M9W6A
0+z0Ui+UrLT+EhfCAOA/cZLeBeV0DKOb5xrjUhZTn72RHhZH7dOnnMtill++LmD8
kbUI54Ga/DpziWJyBkmdJxsFYNjxmFWOKeUOYfllwILZDsDFQPqiXPnjFi9lkh6r
1E/2DAz92Vg/JLLztzQg40SnfrJox6TZLxw3yEmF7utbr6yJVELrcVxiKxihoLfG
QV95FDoiwojsWZvAzKsxRhtexhJrSj2zJV6mMmGDeDp/D9dkljsnkaaloBxPafBT
l8DARyUA1Ab+mR7K5zrNDeqie8PslO+1tZBm5B9KFiGD94FzmU8fezouXj+QelPt
67nGdxf9gzEN5fnG863NH74giLER6pfx6/YavIsw2it6aKkC1jLyI4sxeijvKKCj
fBVwBR7n7xtQp3g6zDjEBUQzWoOtPtqvAyoByRDsWJljTFne65GcGwvYmPdS2gbg
Y24lXygkT/wqz5DZy/EmCRrJPwB0IDDgSsvNt9t9n28d/k/EKPmAqefJDc3kk5tU
89N2uAD2bk4XCAU/KzYkX7Oacsn9fqfqZMrsO+ewb/2nISlyy8/lQUQM+S2O5lYo
TrdUh1Scc+dojYltJ4dk6QLv0zjn+TWFGlUvgos38k6PED0N4QaT6z/u0bYx3vfX
AUE7DIA23nkyxl6n0HK9Mq0O7JyegoOgGt2GWLULIIb3OZNjX/S9u1hW96h4Aa9u
Xa5pdppQg51A/yExsqrcEoub04XmvTchPXd8Nnamn40PskaKTC0wwGUXD1Qxyh8m
kTUh7KDwcqEYBo7bbOIybSPMndTT+YgsF0IuDJE/eErboRIvQaaIDokI6WWulko8
UGKB9/ASj7YdPOEALKrevw4rMYtDY1M54bwFjt4E2FIWWviFzFGVZUl3JWX2RGKh
/DczBreQxvWRSszvih3D/IY+/vHBdbNjPldSvB8GCXvGGVuzN19eeAlD5sj8PYpm
uWgB+xBkWNxPWPYrPm2rE45rxuTl160nOFKpFMjJw/Txn2WQI9w2bu2Rk0+HlWr6
nl3LE2JCC5/TAAyp9juwDk4l1WHvXsce3Y2aHho2rgjbBRFEJfj6KZLkAewCIbz9
oHCd5Vxmny3oVf5rFsNEfvQzK5ooIY32ta97nC19nY3Dy56AAQ4Q3fc+ltVN0uPe
OEv7BhBiT7BEv96EH+XyiyobA4JvRhgEKWks7LVWsHVVMVclX0UuC0TG4hdJC/+O
KNN3ZZV9CytjUhao5f5WLimz2mr4Dywr7KUPrGsHeGSsO9b+5q7vuU6UHdaAwRd1
HDSwjT61CSThChjD+8sc9lJ5SYy5eUrWBbJXV6qoMubyqqSyVGIfHt929D6s995Z
XrZuP9srXtVUP9FCdqX+1Wfz9qALyInku5tKYlkMXOlF6nnYgsjHyyo9roMd7C3W
LxUe4umJfmyry28DaCQtxyWABSn+DA25GRAHKYYwlS2iIMHj0rTSgqmzfgoyoJ4k
H3IZD7py2vvmzvxcob1CeLd7666O3wpvAFkUmq4v3DPW8s050pgSMSo4YOLx7Iqu
iiRcrOh30df9227DGUgLn+Wethdp0l2vbjZw8hhoCe7XBNQhftZ1apDZgGUwkUgE
tEUpbN/dxusYNMBxtavnHQ0JddJVbXeq147o4Yro4XRomxBnGN5rVTLtOdQp7IMS
5YzN335yD7fXVswZN7r7WaC9Gy/MG0GLeZcLgp4sw6mPz+mCiHoc9v1wORR7cK3k
4zuES/EeblLv2cV156xqKN7UQhmfrhkM1wA/6d9nlf8TUGooCtoM0sMTMtyajWtD
AfS1VvDezr/1yBH5lHFoc/dZ4AqyKMGgA6P07zGCeOwrvzBQC+EKEAQry9O8IYIN
xyLHqDKQg0ndeIN8HIkzJsWXD4ErfEINzcD9XOkjHko9xgv1qUgTVNkLhZdUdGsY
8M5w5uRZqnA3Ze7Sxd1gcREXAq/uG07HfJLcMyZ3d2otWD/vMvxIGGoqUBIT98fO
0Ba9nPva1BLVnFJsxmxYvw1U7DedgNdwErZSgra3N7RJDGAeljJ6ro9wvHl3KFZ7
UAKytsHlWo4AAxQ+ks8K+FQRYiGnFLISwneGO6+KaaiTBkkNZgNzAMhhFK+AfPdg
bY4ZxP4uJlXL+3sHsWu/eT0l4t8O1C5dYvRUGf4kB44eVmRmE40nHyv3rAwdZPvA
X6tJXBAKuWkricBecOTbRSAbhjIjUTjQO7DvKsAMa6s6Kep9DOeGW1uK2w7GDOXy
npFlD2HaPsKzgPAJM7k4ln8+ulmyME3kmfQAaK12yVNCxrirtZA+ELGEMsMci5t+
EXBI6pH61a1KYZBXiIm0OgFP9uwQ3kiMYTt0IjN0CwqtoXgf4xQwRa9Pv25wNGvS
dOlyNPW1Kwe0u7NYhtGGRjjzHAokiMu7goMlAbM+AbbyZVUCq2LepXuK5XnyE/m0
rUG/IAjE0hfbJyLl7QOVvgzvE6dZYlUDzq2C8x5UXAIr9jaWlLFZrTO1uQleXv9P
tScZl6EpdD12wR0LaBIFcw51ZpIPKZ5xandCQQiaw6+2/w5f8DipOiz1mwFDKGaI
COttlR7oAjRaTI05/a7lTlKQ3uIInH+lfLsGIbF/bmFx2Pt6X4DkdfXceISriNnT
9WSCB8EIr+m7JFYXY6KG/MLbiEMUjNCvY0lPaYRxQoJM8IbJHx6fnuXP9C+XqENY
5kpV2LFCwyKBTIjHdcU+k5GgolAi6Ds1ikajSTFnVuMVzbdIDTjKB7whuqITdJ8I
G0k6u1XVobb9wnrJJK1kRGbyvunyJ51SccB3he2fOVskzU4YiNFq8lGEdiVzxe0u
6mX9SY2HwIOKJmItCTd5OnOoyNtBdvsM0cRcyTKrSAhidD1IhJouK8e/FrwrZ2/G
/CfQ6jwyrdu7AUZzYY9iQKKo23TjlNQLEWnmgyW5K2CJ/4hC4KnDemancKrlX3EF
rCgID+8SUD3At6/yIu6qCL+GHegKIipqPztrS7ITgwvCj5w0201BlQF1kHLXBXzf
r+qJ6FVYS0oGzxOvH6fQ8xBzqholtEsd3hJFKjGOvUlnclnrb9+W9pVt+jSDAqj/
l1ism6dvHX6r8QZBtSrCSJNh1Rg5aPBkcE5z0yHwtY3IQhepgjbZWgs5zOwNIEln
ZeXuVWi2ZVATNam1P3s7jkIAUcT/G66jsPr+CM2WDCwXwxPdRwPNNdkZtJhCadRw
wf0z4h0/seZScVljHnCW2axb+t/crYILT8t3COMyAEobMLjBYF0hNhJGoGpLQxht
HSA0uwRWjqyJPimiE2R7hVznbAx61ee9sHkR+rRE2EbXhwK4bjtQhE2bxAfdQOmn
pTrYXDSe2fp+mKCYanxtlOlCGO7xFuXX9qUBpkdAKm6WSBYQQyQdy7lMtrkitaWJ
4/68WsHnv2YhqJRlrgIfTMxHgjk0P3+yufRJSNa8piwhrbwA1KXSuTrNNRSkjWzF
Kjal/fojMBZi7ZpWghJZhYEYuP6rBflG0jYIqXUa0oF5EIECYgpHjsoix94lruL4
bdmV7ACqBuJdmaNoJWiAnyNuBOHSYKvnnN0eHMsl5ceV2Go98CoUcMKIgvE4qywf
Zxh/vGaoO4OBYQGU9eg1feC5h5ZxytOIJauK7IccRKkK9QcPj9sgI6kAFtFSd0YU
vkwCSvcL6VPZ2aWaZLSBVIy7qa5dE+Zc0dpZtNw8r6ApXmTGC/M/Lj9L8DI2t6Ch
GRrsIipgsiUFLb6qbVx86qewymOHEdp7FSGF5CmhxFnkJnPAeZgsXUraGR4q6EES
mWQBN8SiLklkd+s/5/ALSUqf3QiQfGTwpSjUjCRU5cmkE/cFdZkwf5HubJuewuNT
ZsDu59ohfVHcYdAL1BVRnV6iScL1fueooee5DXQ/lOO3CDUt2rkVxDluxmCjAUQP
EWwDNoUIhS++YRgbGJENq3vh4iSq0WZLu7guv2AJeAK5+HQdfSm8j38XSQIvrk1V
nEPPwUJiFdM10DeH1/qMZZ6YDPK+o0+brZIVlaHqIt59vi8nBlMPKeN8hjVCF+SH
Nwn8Jp4i7G50CXniPA+bUKRkkOVhiCgmyg+ZE5uhhIJJxG0GTuvOwiJ8YpaNSyVc
Fu9GR2dVLeSPu/YD8t8Y1Om9pS/ygc7k4pS59C5XADBIgyX51A3vWTWHlTvY8zFa
mF2g0/QJn9nKqzy6LuEIREgwYU8XFTqlKDSwFhKTFzTjDnuAq0y+1HnZs6mG01JC
W2w9MKyUsi/SdyOqMLO5fruQMdULYFBJji1hilaK/KQ6IhKBBiRYwF3TK2D8JOwr
h/NTYSv0jGPCXtHoPzR1P+YdV1Gjse9bybHa/pCxz6Dgbuvyx1/7bOSTkUf4wdv7
yzLvyFmZ8l11xcZ/YwaifCVxMeBcDKllx86HITKoU4zm38UsBUeSch41kzHEixAM
aQuopc/l17fMImfn4/39pbF8Pn2SWjErXlet2WgPvDZSoiW+FwApAhLIt1kthR8J
r5exS3WfxDMxConZqqNxnuC7PhJfwJByIkGSwnaotUw/TzC2JKPifU1Fo5JDqQtz
QWlT4jH3CpE4exyiUlql87S8uIYp2PrmnLuTvMJDN/B8yLtr4qRO3P70Qji2Ga7i
5rQWvArsJYWmSA980r4W/HHA4WG345F1slM/d8nA7u5U602GPiUsPFVxfvjGKCWc
IyYpSJS5hnq7Q+oz5OemJekqty3OVR39mv0TU5hz5Kbr/1DcRXj6Ck4tSHW23TOG
zFI1TRcSQopUpAZQ/wG1vncmxmHSHueHDAMsd3ZT1hMNjHNsRbNjWQHU9p/mV7jz
PliW2ZDkpm4WcRe5qH2Dds1Q3w0w5ZppXrYCdPjOYo/KTxV2CG/5eqwUiuCHaGcX
uMG9c7sp5S6zQNMWTIJr1sOqlkWtr5dvcUlR1rXNbACaMeJifQZpD2CouNjjd7Tx
5YwEQKC/OKZXcdm/anxOkKFCT6M5ARBJRDdERMdKceFZ2pBRLf74Om15INOLv+TN
7BN7wt74E/RInWYyWyslVKEbqyrWqkrrkQgE72AoStX7SrbFD4ER5hHWtoZ5ZGfI
sGobGB++H/6VsUCMq5HjpYCf72pj+i1fHuQXfyqjMbVjt5QiK/cDIFQ7Qri9k+BC
GrDox8VPMA/HZZw7CZi0/4OWl7nDwzQGE8SEqnJUgIOw3BrchlgGPA64uyCGPbEr
PwTYyHnkOQaX/nE8GEB9e0OJSUHNfvkJGmuHl3YayfLCokeWl4TG9ytAXLgO3+lP
bvq8uyiWxsyjbRPePhqrUSJuWgtPYliDdg9BFZXxo7NghSybG1zrz2tE5MRZKYxm
SsF5Sk++EvCdBOaPh+jrT+ZwLOAeM7ObMIUndmijHM3FnwW8x/UzPV2nSNNObwNA
VaE37ZE6iqdG+LZb83nDwCgiuKR7+JS1d7AaTf/zbl6svkKvh5+Y/xbtbbtxO8Ln
qBMA8b5vokCnDeM6UyMbFsgqiHj3UWHFlZlTn9MeNg7PeDNeBzlACdR6dcdZxfdG
g5oiu22RWD2Iw7kEoQJrvW57Z73IQ0xY1wVpI5ZwOjT/zgejQfbx94QYG5Eq5VLm
UWHBFbNsDs1VWeJhSmtmoD5CBxZjfgprOnrd8o9ef8Qol3S3G3N4k/jHgzeKDYq+
iDe+o6OJsW8jFmirHFMa3QP4kKVpbdvJmm7zbrdqJhBnvJo88FnvEbQCV84ImRrO
llvGL97iB/D670w/paZnPe2hos5N044k+GSNmqH9XXGBf8V8Oa+wNv/L++Z1IoVr
ZlQ+nr/GCs9bBTe7g/1sQxcOKWOLKqfPHxGr2iOFEWvNhSgaMdHjxv/aj4INqnPc
rm6OPssEUyeJ7kA/6YP5GWB85hjAOU+1VY3PxPiAyMGoAzHBUkGAk4GKaSu7lrr4
h+AfKlFgnc/ltussNcbzd6WIcl8hvKI6gvhQltWQ0yU9Z1QYR2b46oimgk4fJqLI
xR9Z3rGeq4lc+L/hvC5GIFzKL6+ZmYf5ea8nReMFjMXwS5xtWCcaiTxTMGF+xYe5
xQxXr3MZqAVa1XJGujqfdf53WkaHmIuoq3vYJEFS/yRTXPgkCx2K2nlDWIGwPArS
26GSTGuyGh7YS8llUSHCRg8UyJykkitmVFKiSK8s5cPbS3ntdIsliQQo7S15HwCf
B73IycMUaIjrE9G9JZkb3VsTGt2bqvjhoG20OQWxR6gmchzebF81TOR/HQX0A+wc
dEA0bibXiZhIb0Amg7zJHMcgKNds9Qj2Iy/+8kVguh4z698i7EToOOILxFwhhclR
VKsagCnyNNf9JQ3fm6bbXE0UmcevuR/dq/fX4hdVu0tHwoBQ/7tX0j2pt2W8x3G4
nD9aioAjzQt6mCKsKOpESxUJ3BNMj9W2CpojAm974R/BlAHU2yvnRdj4c0crCvh9
7uk2LTtFkMpUWzceE8/ERoVcgDvxuh245dQfsJsnm5fk3X3SuTTGvpj8rIiDYyVA
MXMIrkgK+27j36qVat0I0/r5R1SEKppdHU4lQBqvMIe2KqN9edwEzGXiNRYK/rKA
Tm+ZAmuyit0KFsiQd/6VMuYrAaLUGnl8vS4JSXsA+tQfjk88Bvy0taQ53gjGsEuQ
Uqf18GLe52HOd6Jrz7c9zzwPZKPp2at6INJI13+PRU7sXFdvdIy6Qa55zxz9uz0c
K/pae9su4BRwmWja7Ty6GAo2v22qQoNlNfHb1GLSB5ekEt6h4R9dAoR8T888BR9p
crtsug6CmwKISIFzfbvmnAKwUufJAxnCHZMeCT48nhLoBB9wRQxcige9lpKmwTFO
opt4yzjFGUR9thxrNTyHRYvKNgKccIl/yIr62sf3QRwaJu9dSYLdoyOMhkqdchwB
z1Vioshxgwa6Qh1SoR6rtIU+toJCm+TYthQuqpFHGP6lsd4KSz01Gp7UAgBylvCy
AzhcN8cbN5Mrgc35C224I6o9w8eTmRDK29BGGXWs5LtwkuBBpD7UucS7QmJ9kkss
0fivuV+1ops6zpGiDuSXtqjdtLuaVcwtIbqPndf9DAfN0eqcU0fsL4AaUXYZ4pWH
icquEES42L3m8+Uw5ZGhLJpAT7/GoHXvxcxNIITJuvQ0z5Ilzt7kP9lbxXttL07c
yMgpsaQ6Jk5L5dzSsBpuimulRLb3YFv2prGuynKGc0QgLff3+e8VELIGPQvYay7f
pIXGr+3Qmnk9Dqt8heTUcVV/HtuD2keVD3tmpgJspDpucGUJ9YVpuc2tDULWWOk4
a217LeMtHF8XZhR/0HrW5m1ieWjY8oZP8jlArthpwSzw2dZvrAB4/d2GrZSfScy0
11nLdXqyo5VWdHPmNzuXR2BuJKxO05mwe6X4at+SerDSYQcht+4aw5YNepiSRmB3
YiRlniWOQukwPVwbdicSjdhiELNqpQtjBf2S7livczrOmXV046de832vOhJTBwrC
OeWF9uAcVNSsPCQwednwJAcDWDz/0aOtZFPVPVMrdOC0Vu2LDN2gBouB5iV967Ss
ltKFqgLtBrnd18kzkysWmQXxJRDEzso2JMEyxDRjV6R4/fmcyGQTE8ALxheh8R+t
48FVAnwTYLkexP9/oT4Drr5h6sNPqCR75VSOL7K4cjXXKFXtFhBfRCkqw6aRhI5S
WHcX2mRB9bpMnhU3Y1YrOXYXxQuLNqIGfJwW99z+meGTXp8fmEY9Z60UxBxhebfU
cY+DSkGxEygEU6Krm4aMMMaBBlJmRpNif9DU4Dr9G9AeH//57lqYDqfB+7y5GY/0
SLVQnMlxxVPo+pSL7TBxjpIILCgwGYWX5lqn/3Z9fvN5XIDaQQWZgNVUYXKDMtsy
ztYfj8IHHkqXm5+WF9b1w2rQQV5dKSDQWRNWSRVN/Hf8b9xBF/dI1LML/YFLn+Rs
hmRpyIaVfnfGUkaVhn85AKriRfCj8rEbojWDRisqpErnwW5PlQZZ1TAMw+WL3hws
tbFlc6N5CWHLDmwNR7HoCNE/1jfNMYT+1fr0+laDPGNdlr9pU/UhmAtGQQBclC3L
NtVf6mJWoeDKHb8JG33aVDnci7iSeRsa8H3LCx3k+V53T7WT4BinaylLDZ1pMRdc
r7LDq3fKUH//80UxCkSRqbVu07sC0dKhjA8E9JRutRy2J7X1b2J2DsRqMYGk/FNL
4EyLCNa/5p6UvJiND2W2g/uuFB4BRxv+M8CVSkMYhKzbb5ol8MUvFC4TVYb7FyVG
fZgFM9MsV+bI5k9Unge2DjLMEploJnpL8yg2QnvpknQ6JVHqft3dLRBSz6JQrqsZ
aOwLf+hUIzi1PnJGUHZ/jNqR4lSVe+4zWvms5wcDsmNkugaeMS5Wt3+hlX93S4UO
/GlRvl1BZuoMDx4fWxKblro6CmFTaGgQF372a6w1G8YuvRkJmUA5ggl538hptEcb
eRjH8MWc2ruTIfcq+2XE3mJZ4AwJR4ux4YIKCKy7xw4d7dZGPFkhz4mh90gmIItl
vpO4KP7Fa4t+/bPZGJLzlU4qurB7bEJf8GXmq9b2pFXL3lhe7Ydzs0sufOHMJg4K
IPMoJQzVAqVTGZ8rXgHm/hChdt7qDMbwRsu6y6qeW5QRM0DxfEVDRWkVu0ZS0syW
IG9Adt3PpMoHRtqYu9UhkFWomc561RpTGzLLJ7ck1AUFgl1CAMRrmG78gY7aK2yC
s90GbgDY0oATe1vdAM0r1KmBHYan78PfXbGBdIOyujhN+vrZPsV6LA371UoVft7T
6D7mN5Ok5poDbnkMcHbbmgc7rSrNLY+es4tjUiiAghpLkuhBr9MMT8UXYCbPw2nr
xv1x7Jey+BRCRyW64eiHAL2AXn0GN8j72reamj/pLJ7RtbR9dJIgFnflZR6Q+GlN
R6LODM1OeiLKdMUCSi2HZUsucZieZb3QY0ADHLZpR7QH9mAwHPz3bQDijHfUjgdz
N0YzlTK9w9rNAzUELDlxHytif5A+cNQpVIP7BuFozmGpOvFQa6l7s/3rVRYOESks
8JDDG6J11YOnGZmczeB2mXUHBQZXDUBBFh/dzVoLFS5PHApnmICYhO+lkwr1+33o
K4nTs8QTu5ud1l9trEFxPnEinj+trksxiuxF9VKNYlO33STPGPxTjAsrAw9iyggp
WkXj/20goBy879rUlFeCsD5h5j650S89vTj8U6Q4nF0IKwc8O6+5AORliGZZhbVd
9JLTCO2p3GPhF0zCnHsWgek+m95m7M9ae3mFxyPWnn25u0Dvf7O4qJrwarLXp07u
I9K4b6dugXXbyj/iqnHPTJSweaDHtfOkKxs5kPdxeE7NnQZ1ACVJ7++iUuDChHW6
bdOUWvEId8WBN0mQXL7bQwhDB7f0VdPr4vnhxGDwyCtpRS/jOzDgqxcY1CTDh55r
w/e1fMZA9J9XS8O8jPitafMrGHrWA4MUtgCXgS50s1N8gE2wydldyPIRSGmC4VDr
ILob/4FCohb5vqSjpjf1NTvYpkQbQjLuyq8VtFsqjGSbLxxvwMnBLEriKyyEvrJj
D+HHFbieP1J3K7F6dEdCKBNHXzj8St6GO28/6vPERmXGcm1iJxMGyFH1d3FDT1ll
bfv5ksi+qLYEkQ1q0mV30Rb5wqzKR+cnKfQFOae+j4mp87m4C0YPedVFmGWPPooj
XaYU/qCwuFNj4CEtBlYWMnxJAZGVyLz91LWS+B5vYI3deRtpSBdEioMoiJA181su
f09G3giSRbLDjC9d1Bn52RFgIqYRujzhd7WvE+5jH57qA4R4IgrXkBB/P3apajUH
Q8B7jeDaDGs4/pVCTcHZp3RvHKWQyst7romTpTYvdIuokfNvcqRklReet+G7dgiP
BxVth7vch8UXhG3St6jBAG5n3pmYYiQihRjCEO8JMlqDwUP9P1y7912hjXWTFZkE
e1FJFSgYaiFrif4u4EfqDg7Sz4YgBH2RNmfR1G+mhB5z2kLZGwiNYFSuphDNUUWR
mwqZywBX1wsllQ5IjuqsR8i9BUiQgoQr0TAg8LX5dQo0c3WpCc4JyQsJyeUkR28P
1fG4smRUlAa005qif9pkGfJTL2iBCYFC6u6pMDemU1c3ifRe7c08VqThvWsTtc+5
qChcCzsEknntG9gMyLiGDvYZNkaUFD9pLf1TX09Qxk6AhQCbZrThT5LjvYDMTOHi
uW4lA1l2Qjvv3A1MhoYrBxzJOEDbfqOAI3LgL74fz+ttkdjx60mCPzokANL/Jgs4
9O9MKBnJpL4UmHwTvmYPli4Kp/ZoQWyJLDp3knc+HqDXV8Ho3fKutMFgKVZso187
eL5H537CE9tZB+HQPZ4gSeFp55OKypqE8TpkOUJpm/HFdmSViA8oBeMYCBuJHPNH
W84j7vhHJ116zZ0Vdhl58reqo8Q6AZljnuuINf1WCXJWa6Xoa+wuzccM+528ti/7
erNRzAacx9ykwTg8jd4YdvfY7NIqCxU/6RXZvniXmRs1uuTGxS/f0SBTsxpnFT1j
dCbeRZ4Xs3X1VZ6B/UnX21C0V9dTcCLs4IVQIfK04QLlpHCP2QfUZmI1n8xw3M6l
sw3dBQD9STot6sjT5fm+3uRxqiJA6L+75RGQ50jJw11d7LRbTY+qxoVvA4Im5/Nc
190Ipa7iNHrlNS3XRfFCK5GVXyWjs5GvM9MonXraeXcrhiKe1+1ZqnUsMq/XLOXk
Ra5+3NJ2fIn6LWcwYYJh8kjbmWNJhaV5SyjgaAHJeXQ840LJaHnVMkbFa6D8g5y4
Pryv4lgQfdNvWNWQJ7sCNzZjdBfDBnzSZ0z2i/psE3T/OVyd05T109DCPxGA1WO1
HgiFwZ67ixKCH6HWA6FQpWa8GEOlQa4E7NEQX9WbNx+AhDVXgsEZXuAe5vKz2rZR
WMTpJa/F1DMR93HH50Kky7P9m5/f1IPfDrmyT7308vjgGJ8zcR/VdmKUvsCNkc1K
UNl0TKKfHirtKDOCdMVNo3Dk0yuyAaLkPVllQzK9e2JYo8/3mM5dBHqNiyO8USJP
1GOIcOKzHoBqGb+xhlhogTFnU/HR+k1/R7yRMVzok7jxNOsyqgy7ikRKyrcsyqAE
GLBZ9RcKfxDsEEqHWnX7VaeoCkaY7T6Qmqxtd/hRQy34oTl4YtE/75HYQMVP5s0v
usqBDnPZhJVh1D3D6rcCelU3jcP/O9N5ZuHP1dfdD43nIsM0X7WKJWOW6N0/Z5xK
i6d7hm39WLt+Og5gsLsAD/iQEmO1uSgQHmhdODiuoB21/kGxVWnN+TCz7u2TX/S4
NrYx7PCypGz9LfFMQdwH3cdqeVaf5HPpUiChbWXPuG4j+xPG2EW8FObZJFfCd0mp
qLimcz7/7qJV7Yx9Uu3fCWj86UpZJcowvIGslWs6YawMjyjbnRdbS1mjtFA0OFf3
XJFc8lTHqi9jNw789c02lrlk4AsqDg1NSeDBJLjJLUxPP6WYnXl9GK5i8DNvCINl
D6QMgFOtMHrGvsL9prYK4bRWFiJs4jaBlQKV8IK8NtV9SkM/EVIsEm5OZymJntZ3
ONi8CXw/f8Q0bHzhKW367sY4HIh8thureNdLK1pZ/wsqrIWPcY+dkhQY9Q+GsvY7
MjiELjEvNjCLGwl2ooLSpa0VFvIC4wCPPYkRTXuagH/tac1BOQ4zMfKtTB3k5upt
rtzYR4pRhDHWQa4gld5LkH/0CYssEof0FavyhVlZe+eu5Mpvl7KR6E0xaJnAGdmA
sKdVUTRfF56xLYYZ9B88L7G52ZR5G4z+qIRIKahb3eghNUdtSjs+OVZCauEk3GE/
81t151oLFlfASsPXOeGGV/IE3Iw3EEyixoFvKgG6+efO+vLC22sZl9Av3dqVWAQY
oavHYBnqMEu2YwiPv+w+2Xq0TUk2JxiIY9hlD70Sytx5Z+/YgYBimdrdkJPXCH4M
HeXdM+ylYbuJsRq6Jdy2r2hkSJ4+/d0d+ChS0zpj/bOVwncrm/xcAjF24NnKJC+3
CJisgdnSVrS6zRvbpqz+eumHCYYKJgTmvwfF7shKZheVyuIMCopxeuU8bypEp8Ty
MtxDw9KJxQv64123KkRwTWhWZtuK8QBKlljZclNvYSj0350tX7oeHCOC3Igrfrx8
WvTe2pxuoDjKwzOm2eJrEDrkN/sW+vXdtPN0s6gMlBRZ4TZM70pKZqWpGDKvFpAc
oy8redfR335N41eb/vDDRdAmIKO2EkGOiP7C7V86EJiINYEEVvQvYA1UrmxZ4YCf
N4u5eOPmab87M+MiirWiQ0VjWJo5kgvZctqnQF0LsLKzACtZ2RYfh3g5+fFLLd42
XuQVI3TwTkuKC7Sa6M03thxeqjKKCqMtxCUOK2mUmdCrjmtaSbx81WilkY0ri7lR
PsPLL6eN8nT129tFcc0u/4kMnfwNb79viUiEQw7U2QqmRMVmydix5+nGb6di8UyQ
29jQbdyqzuzNQ3kYH8GsrHTql6XbCFh48xA30GMwJAytwJ6hCV/sLR0ge9Nxp1fa
RUYfY0XyUmL92ebHAvNSKBNijJdWa4w5s7UFjXhkJaWaRGybSlE7S7O2cWSn6Id2
CEPppwHtjn1H3IX4lqIhaWQfx3ZlxuKlFBUhiMQ+zyxE05txdDgXJrYi1Ipvlxnp
bTkh6rSvN/8K1fL4xliJLVr/ACBs6/zJ/t122fIsTbjqCAcoDbRsfK1FZF1y6UmD
HAdxj1b+gLBK5dYHerzPIshs8tbCpNnOruT2xr/NXKpoeAPKPsGUVaVZLuDmBFjq
zctxZHh5pMA0bOXj3xBsjk4GoKNP/8s56vaaILm+O+JaSu55TLoFKnPYDNPt/eHK
UO7h88cL6xvoQC+w8dhQz3wS/wOvJ/8S0dPwigVBO5vRMvMkCZRtgzJm0SoeSUSW
E/T6sadnujjl6DwQ0Z1IrpMitJ+hxIVzzaHvLuy/FSlAAZP9fub3CWnU8UTf3rx4
hn4F8rKlDfzAtWy4J+cHED8xb3stwr1IbwjTyOPkdWenvw7TpiA+K8Mgqrk/CPUb
f/ILgCisU6vcgkRGjNQ+NwePAUfm1mY/zxhvArqMttKXOMoFrW8byexoOWVZsqBX
Yyo0aSWd9WbtIyPeN2FKNB3s5wVmHsR5g+Hho8n2BLDDVmZs8au6+zZXFUY5jB0y
9gbIGaZv8TVRnmDIRo8HmFuyB1pX02X/nokY5hDTvFOgeeJRm3ut698BmuB9dnAZ
zPxfbXSWmnY6/d5XKkbbaZkKuhUz+vfF2bU2lUmpjdxzYMuqxZDm7zcbwpjgQ2AX
5+OIFttRU6hr8Scs2DMAmIwCH18VVmp1CKTBRiMe9IYKpExSVWAHMLnfNh10soic
1O+tITBTTGzNb6siWvTyCvVu1tXcMiK+lWtK4zFxOYwZ8L80hDgya7N8G7EqKf3u
o4BgiGw0crRqmtzGDQ1EtjAEOL5Qr6oQu7WqOo44te7wpt/ntYgZQRZ69d1Zr+q1
Y5q7hYhf8mSMAvcZwvB2OsIB2T1oCGMWcM87ZNbq2YBuK89bQhWDr8vSBdg59QvF
ZIC+u1+pNbWjr6GaEqzncgJokahHecpYwXjcbG32xYCc1iMwV8Pj1A43LSSKc0Sj
O4nZGa4SFnmvriNlt5q780pA6cyIohiwlhHb7whOZ5XXaqMrkG9NI/WHxtuPiNnf
6ec97QYhhXQfTDQDvTFicgia8a7NFja3BTUnOap2o4zKUtvbzoXd2/2vifOVUfwu
B1WBj0kjhVYSem+uBik4HKP0JBNbqOYcHWqCgMFRegLxiJ/0odriIVsjrwMfLzeB
nAaGIfwARh7eeSicP94+YeIUlI1BDZtUnWka91UhrWC/Wt2ff14poM4OYElIoLWl
3ub0cdLpdNErxFMlAs8Zim5PKRDM4SNwRa6QwtZKtBRbuwPEns/G3moGXLC+K+XM
32mejajOpYuTLSiCMmAOu9EoXflXyUUO6HNU2f/Ahe2Ln3fKz1WN5bIJ9qUsasLU
lPAfDcO+oJftZ+roLtWKEhVOvm/G3N5lWkx9nItSNlQ+zur3Orry49lkDuUC3Y3p
Mb54YXeoOfUG6Mpo2Wo5Hqg/ZLX+Wd2xuJsoXXpEghOdEjk6aBVfCT/9eaXuwot6
Q6CT1sPm+lvRu7Iwv872wD7nB2HrsD4btBWh35TEDGCe2Y0BaybZbkOiPOMDlAPu
PaMntaHXKx4Se99zectOn0wK1BB5NVTIBS+FdXuQa++AUpBhVirr2oWyF6zfkJ5x
/Fp0FcHalD/s7aX8KqeIxxTPGu1vYoYnkLbt1w9JbYI4Mii2msRn03nUkn/9L+6L
rmRLSSzocfzT5N1Gs1FJc7xo6DKSXQGngeIO6I/fSuKX1hPjoP9CYf7Yckr1FZ8b
388BJCFA7+Vvg5ptTsTpNrcqloEnwxOxxuT5QAFN2/9s6C9wPGacsNDpamprFdky
fJ1scYr/jQwFnukeFxEwdUOqXjUNkL6Eva0SBn690zxjuFmTB8/YuHg6bxh+2/dX
kYcJBDF+PBhXiWQUMvhn5Q3eSa1PXuJpI7C9BVGyqwPewghp5SoOv+NK7aeefy/B
l2FKYNqxHKGIobh9NpKHRh89GEis+NjXt/QMxWCB0uIqs7Hh4LRmm+R/11ULYaix
dskVuETMsJ1P/thkojPECi9ruZebEKW51unZGTkc1dvv/4AD841LfkOt+h/J507g
CtK9RfUGpvIEnBiYJH7FbhxHyb/JqvpSUsWEpb1er2gh8g2bpaYr9SnKv7W5iPQy
mFkTIZSz8k7toD0ZGxoCpPfJ6zbcfUAgHTyKvIaENQ8e7Ic0LGpXCkh6H1VeYTy8
b8LLl0ozJ0kuI6ZMJjWJii/9uNPYR1jtDl9Gm+dI1TPO2YhAVPGhal0eAeBTqdo7
L+pjwwfwK4/pxY9/xb909bSrytCKBXWmaP6e2C8jsEVtPYI4CP0JA7TiNtnjXs94
5xfCtRsbIPe4cHwepAUaetiDd5Lp+57a26Yl+n9p+NL8wJmWrhyjePNnk5d3jNAk
hItVw9UPDPeIFHxEgO1N+LaLWDKhMEh3spCKAL/Etor+IZN9dHZZJou/aUGxd9NV
UHlAKRdcNCNnyTpw2Y/ZBc+/lXnkMRQt9plf5bMAEqvztC6npWmKBaAlaWPtadTY
x9Of9uZrYIadI9dktwf+0KesEFKG9VY5py4hOFIR51B1KJgb8NmX9ZHlha8Hknjf
gFpiyXz1dyjs199tWNU9RXj3yQznc5N8wkv/2eaSFkrdh31mXP8IMWRC9YF8iWcB
KuICEdyNu3IZW017qQFU0XF/zJW179S504wcgcxNHxsb8getUp4Qj5XD7YTUcJtj
28s39BAcrnIv2y2FmDL4shMB0ZWQQjuduyFshWWq6X0xiNkH5LqsUZW9z8yex+F9
06gVvXCW39wkvaUpPHc3RVlJ3PzSonvwqYJf1MyFlazBX3B1avyDVUYt8FM1eupa
rIcWlwSsQuzrlnZK+jEIk1/DCc11MSYTlbVja7fQNdlR6faAXoIjorSmmrupHFhW
9OEERu46mNz8m4mh6g1AsR3tgV0xVwE8Vl+kPXvcaaBE+6PEVGlsWz+nE1IwzJbJ
nZPP/wggBLipY1FWOqd5fEXOQt8wW4r7QxEO+e2PjH1qN5MDty74DmyD57aDVL8X
rvgibxwVXvvRSv2HFfBtPVlW6jM3mogXtHVy1HvTEPcdfYgHLmaD+TghHQA9INAE
kJ5hvPgKMSW/IU2qmz8oobmeOeyMj2/SpTjDBossT7mYPXXR58a2fUeoEQtIBCAo
Jl9AhMUHDUtomMdltjwoZLcbqXVX5FUlE6FO0D+OwTottZj+sAHZ8Gg46pg09CZe
Xu/D9coJEje2b9lyjmO2PRdYWRr7wBMwCq0xH3SP/OjDACeTdi5EBus1G9gJpLbP
+HzgSiinhprrpz//4Qw4mRqokWa5XxUpsBZg96yr098W4As15AO+6J9Q2qiYJzTe
jmTAi/bGtVv7fcEQp4V3T5H34KEFhbtH3HHKzU4KQllpBKb7oYtFLFrs5oXZ3Y4T
DDQAR5HpKcme+hD0EpuTgFNI5IbsKPIyoIjO31XrNdWjrBx7d+3kKeJONCANwUcZ
WY58vPDr4IgvzmALQoSG8DupehKxUtoHZohSx8Ulx8R7qDnjp35lUHYS7BVJ+l0Q
JE1yLkX7/OhLKdtaAWNIvdGNTv3lhCzka4G1krIj5A/j90Itqp2HKF9/nmuAht35
JQ/czBbecJ5pqdv7xpX+kdTv/6SlOVL+pW/iden8HHrD6zMC7t2b1WUqNJKJJUg3
ZukqKrnPUrn4rFL0I3Arf08cDqDJAAPPjuAXa1b/XFCN0wZeVeXjYL5ueL1V831t
IpIVtUNLsrRubk+eIiXDeR9NNT4XGPsugyaX3T+iE1sPSuybaBfGrD4gG1gqmerX
B8/vWx/aryCwduBmbXLx1UjzhS7xVme+yvSzkDaJ1fCOXXHRWGvVA0e7MecRjp4J
OScPmEweQUWvypdH9YeU2jpDaF9XHqC3RJaCuifdHGA6fYHtjWnvg+/O2duZ4QBp
TO75pmTBgq8d11uKA3a+M8fV/Kmj2NDt/ui3lIxgtztxDL0qFOTTzg/fDywTLXgQ
BQyzn3A+SuEVM8Kzo/bcxNl3f572X4LcXS9o7Wh5yOz1qSXEg/75gXRU9O3cVC22
RyyjAjtRxQFACRmSUrTqOmj1qnklZIHcF/7QgQL8/OgzJpK7VSKN92p70JD0/4eI
ECvNd/r/KywUe/UbzoLLeLfcrCBvGrXDlivcMuYr1LgtkFZGz8/8TChNSW4bkk7r
ldGL+BvbWP12tF+27rHo8keOQLVGiJOOS25Y7XUy5ezDn6qyblY4pYqiA2I2iQuq
MQznKsbO0Kh/YLFwAM/vE8ODRN134ovWVutU0dN+krKC20MBll9DtjokB48xtnFP
mrpRdIW1EZ+JJ02EHHYsV0rdkvLJDF7Y3yKED8FnFp/rbLYhlaNR+J8nbXmFIqHk
c4EN3iS9Zs0RfJSDgvkeDUd8aYOqeY/4bXiMeN+tLkSQAFFBg/8kC85vhWo0lx8P
6sxdVaOldMOhu70B+q2Go5KVzwO0Bln8WIbkgCGl+PbDoeoYZ+qjbX3oNaHyg16U
GQc+SWTXxcltUoktx63jAEDgxgSq9VtdZ79blKi5fAmUgtuOv5CtgExDzHdijQXG
IH00wPwS+Rhg2bAL0pFZBMQ6o5lk58ShARVVs8c/DLv1L/SN3TlJ8vdjhLhwoGT2
+LIofId2n+zkWXU2JCHJkcKyswrIw5aCuVpfNTdjJjQ3IcoGLEMRA6/hIv5pbEiJ
/7+9Bks2nwxrSPb8eRiOsXPiXLLYnS5lk+bIXqGsrXIeLGmkKoRxMMjmo1FMmEqS
ClDbL0TTXK3/fvnBcPvXAt3PUfPKCVPou3+G8AEdNNKignNSaYa0U6LG6hKSC6od
QLSjq2tRYsMOFyB7LdB4n+DqhwQsm8fBAD5lPWsfV1TGtyICmSuptDdOznfLrr/J
bRXD5QN9rMmuxQYdxgmljkCXWNiK2U/jW0/kX0H/u9aH8eYHgE0dkogDMsVSiVNB
8ll56Ihqw3lwottNgPenf4PZb8wBNUQ41sfgRtv1FakqTyJ7e3o3wtvK0cstnSiy
p3eZpaX21w+Ikgm2A957ByhDOhXfIwKMbjZaLNKBKXOAUhaxnZNsl1XnaLVKVJj8
IJ8BzmqEJRclCqwyVDgVyACKEMHAFyONV88XFjJRjr+9s7UV24l4KDNF6JxRNF8r
rCseCfrBgEzvcbK9nf1TKeBAwwGzGKm8ToSzT/rARUiZ9hCH1C2PtcXWvs2gYJ0q
HRi7nWQsxqIIcIvG93119+oFn9l0ko2UDoM0fyzyuiXdvDM6p6Q5Z2jzegqPSK3D
sJMkPXRGg8G/FVZSYiH3vIKaE0YG/dQAspVRuLdx0Y2AD5zpym4IskwqatlYu2AS
vWC6XoBBkQptp8yVbRDhwoEB4yZYX/aC+Am+2P0mTIqzYOBsXjLaAknzXVhwQoZM
eJPMTReeiGan1ge1kwcAFH3Epche5j/qWdZTlx4WD3HwdL0uHW3HTyH4p9lSCbLe
SVpDV31A3l8GZkmtDlR9H8iPbZHRXiLs9ucUjlnH+MiyPKNi1NZpzPB8myJYXVrz
AFWcMKMCwYOr0RqqsVbhPXg9XMGpQFFmsLbeO4puY2upHYSFyUUv9cKEOj4dZ+Hx
C7djnK0WQTjztyEEvIaUXZdFdcQ21jR1I/IbpdmJ7wxRGFUKYakyY+om6PxwuK1K
EMJU31QZT/0R0K8Z6f8Rwf3Fsp5DQK05EqouDsCLDGvLnxDy/PMzlZ1vI1Y0+SJ+
Dzp3egojAXqL9VhYbGXr1dZrguz/8LSmLtF0pu0qGckc0WzmckgPui2pk/z9Yr5J
RgMJVYBIyzxYmpnRlMEd2KqNMXK87PsNO2pL7LUQNQV127bihTttHJyCsAuCuQKj
6B3LJeMox2hrR9F6eYnXfwd9CAYdpLZY3cWITGgvAWNiKWGJ1sbZPnp+pLwRZeSo
iD3ZOJQW/i3m2HgQDM2H4tvzIa+JMt7DW0Sg5AAhxYcuF7Ypt2Q2Fgy4h8LrL8SX
b1NDi+P3OYlKoq6BgHG1kNWkMQmkvqqCxt7okM7DfgB84eud421ag9gwK0nbMSg5
8f53fBej2HPDAPM4Xhvf9uUUbVGzQuLq5Y0b/kB4WYj/sI1V76tnYxkJ/m0lRsz9
dgaaWr3wrIvZc1ID0GjyLpSEmx47YEqypOZghDMufkHpXh/X7kjGsfJTp7wVUw+N
dQraBH+96JLZ9OgEar3vz4yhNWIJBKnnTOrY26g8HPbBKJ5LApcBmlzy9zj480ll
+WOtIMwIvuTb2oUrcJu94a5A2K2EZf4ymxxqSXgZiGuyAIx10wDcJQfbuKmTq+pZ
gJuHF7dalfceVybeWiedhufdbvUCDUq1gmLfqeYjcWxFIWYcLseMgyuhUI41hM1Q
YQMU/ITtgHBvN9BlSvs2VrPnMuoowveN0nx0LXqQ9nNNfUmInQyNExcbUEsMYquA
ICi2T66ywpVtjPFk9FDhL3sYKGq4Y+HQQ5/kPhEQf4VhWtC4/HL87CHktVItzRH8
OvmfkWi3TOHk2G+K6y3J6YxQh46JxHIn4cZnK8Q0vcqNZwEy5eeGSdDL66+yMz3r
1FKEOK3QTL6HSsksZSpMu22CjPnx9p//n/NcWUcAzS3rCsTJKJBQ+lTEjuHhf9t2
2aqT7VowTVT44H/Dvx3uqGz1Bdbb8/jDRRwO2g0VbR1qZ4PpDf7vT1b9Qu1YN+TC
f1ElfB7K7yeazpql+IwbD/P30F/rcsj3eNsq+LESQWfmY5vYmdcW0sJJVk/YYDjM
S39vf6yJm1gTL5fhZrfmEMLlZiX61ocMZVKLbO7jLoLwuzka+ZrGXujhTTnbWaMJ
0GXaCUrP9heIzYNajrtmIIRrBBaMSeNgXIAzj7yCT4BBoirAaiejftcePha2rHVD
PPIx8ImGhSN50nMA/9Tf6zaY3PpB0V35WiMEoJNjU1HY9f9TNGc9rH3ro591N8+d
lDbsOpgjKh6oh8psUmpcDtep7q6sorgXXiMKmBk+E5njtIStaYFnQWXHF3IvSiZU
dCGUkNid4jEQs2fr5tOMbpsS0dlVOOjahiX64TUgknSK22StCUEuEPfuU+nQzRV9
2SFGjH2gSdRy0LCDs4p0pgJTwfc9Uw3AwEs+L+IB2mHZ1psvirAraJGChkAygN/9
l4n2clDIX/Kg1hH7MtzsC3hrcWuY5pXJXxcK7349QVYNtLbrEc6wfHNYrpf42lGi
EWcHyoJX/KExaQS6gu2kk/RVp5naK9SwXad4Ps60dlbqBk9cV9cqIX2hMWEoYqFy
CrHjZ31yAZLAahKMlGB2bSEfsDn2Oq4Mq4I0zeifyLpxM9b/ULFDTuW/6jfy91dR
iWfnLVvDOzVZxi3dEKDjCid6rbl+lBkxMxpm7opemIEfgrIZPajCT3j7Qrk2mS8a
XMVNGgC1qDTBxLDSFaz27GZH5NNT7TijQEh+eSEEXg53j2SwO6WpNVzWAhGHyZ6W
277kXkbeJvCEQdyhQOjidUd2z9hF0ipieKYWNAa8Jb0ChAtN0EI8H7tz2sBd/LkD
+iTeAqvIR4FlKdEgklVvsqvRnTGGKzMT2Z91uAfSFH8sZoezYF64HDG0amnFHPk5
L7Q1S32CgXqQ8xIEHr6NfXV6q2/pnpYn3hrdpMLJSA28Db6RfixlmCB3Kg84rNyX
4b+0KcdaUv/aGj6jS2JExJ++9Ibd/0sEUdQprYp4b8fFLvN8SWKTfdI4WOdkew48
cSnV1QcKqRIf7JpUFE63H8ltCBaMwiqbrnmG84ZQb3W6YzCk8KkKyy2v5sd2ALdI
7JATix+qduef5ntPhdlaqJbWl2uEX+1LmWKpC43iMlezNYCLwMbCM/j2Fq6HNzRn
CKZqmO7yJ9xpGO+LN+I3t4m14O+zMaEPCgbKu7PPRYzC+ZB6VnF6qyxbSw4jNZJU
y9dXBQv1UUSaZt06OOHnOcsXadl/wsLachMW3yzX2igTGW66gdoxyZBsiOsbqHhD
39ClqbVcWxMrU/TgqMtF0alLDgw4H1ItpzlZj72ZsUCB+Xq6aSEiA6jWEOdA3Qnw
HzG9jpS3gHefWide7jxitkDc9w7W2gwB3UE7WHWhqz2uPx9c1vdVZkWM1ehQkAhi
aybZtx047UFMSXArELpwMTv+CWfR/q8hH+pjNaLLH2NRTIuotUbPLpQhSHJFZnAi
eorI3YZuKnujy/njXdR45RxaHu3z7YtdIun++LCkAZlCjNj1Ib90zTxOj3Qu9y/C
gZRFabHulD0npbsgVtHvQADs+9Xt1nI+5whpwMJwgYcyBtOcLHJJk65YN9naD+bi
/c7xkWRuGK4e/zUH5Fh8Q0+IVv7RnW+vRb4qJPjXM05ycHnbqw84VSQhjQTRDftr
M/7jq9IVEW27w0PA2gRQWSuoGnBSmPHhOlO2omoRRu2EtF3fEoV9f/rQav2AmEEI
NY9wexAytZ7KAXk0RcXXCRrW4YKK8QaYMko25bD03iupSqRGvPNKBa4hPZU16ciD
Cq7gDkoM+JucSZ6Je8gG2RJRiQ0kg3CCD10svalk3t5o9ybSvjHi0prS7f05DQph
akM4nw5MxBWdVcXg+3hg1gArWnhcf858yfhB6h2bJcRRx3M4I2ruKTuGXjgeb0jS
Sdt/1Q+VIFX1G1gE83eoy50rGnh8JTEcU20n0liiydub8FOLd4dssCFKfhhuCTBX
ySbnee7rx3dzyzbkPIVRZJGE7GLa1fPxk+KHQlm2UV1CMVTRI9pk1sEi1GxXx6eq
agKeoQC8jeFM/HLceA2ioG1Wk+eUioG1+mWrGboOG8YGyu/lEeaPBt447sdqldLy
kHyMB7WRIbshzog8Qx+/lPje6tbN8h/yc05pN6Ra3vng1C0zQhzqC78Y15zbnlbH
MQz8RiPKRZtTtGE1QU0RFpGDDPA8vo8IogtLkvOjjJzFxMsBy5oLvXRmJ9FbjByJ
9Lx3aT3G+DEhR6HXpgNeY7SnQzJaWoKAq98CVrGgiXnusjCSk9DL/rTo/OmsoXhz
JACS//GB4AWe+hyRklUubeogeSZdY7rkNOG4EyXpAqGBFbwEWj+6s/c15HVd8SyQ
SRQyMTjNjlB+4jGSyd9fbZUnkO1f8Tdde+f0PrFicaBk019K+gxS5nIwxhXLl+O+
3sxnNkZm/SfMFAHMnPXsl2vkxYdj4sfOJgi1iI9cpv9HLLiqtljVnWl+urSF+M+S
BA6JtzYkLEXr5iGp3t4iwAPfVaUGZ8CfB1eoQkqmTvL6QPFukpX5axP2xXQ5vHJu
SBiqqpkZ72fod84vfVHErYqsCPEqO2niT/pmkGudlc+fbO5b2g/w4yx3sUUu6mbz
kfci/8XX72hXwbGGCO6BiG3oh3gAVgG0UNqBCtedCrVXde1SI1LGQb1T0pyt3xD3
7Fy2FRE+CYQWX28kMCuCV5Zg1R5HQ2d5c7aiSEbV6uZauvl8Wgw/8cAZ2JqnmlCP
uYPHPr+Dba2Uff/PvGl736nwaeMwck7AV3JTGh704xAdGzgT+2ej7dLdQElpGR+P
M9mNAv8FBmJxauJZm2U5y5K0D9AegbL2ExqImSK4blbHXSE5KPZM4BJ7ei3MyVeu
b4WkZ1bL8gx5a+7qWtZ3RmDtc+UZo2Q8b4paoIMjON2C0nViloAaKMKsCOCP/CBf
WriiJrT50eGz0Ezm4/lgL1H1zJQYW7UszUBJ5WOHwmFeXIVWuegtzdin2l/HQ1vK
7kWkwWg+/LXBQCZc97HM+0XeojZNJZYrKSelFpIiMg3ZefWFw3bD65SgFA+2aTCn
zl6E3YGOQKjAR8HXuDa/gy5Si97ug7JaCpGxjN8r5WYet5+QL/Hrb1F8/ta06qjj
o7PuHVGr7OHfCjbDW5wZVH2tUc5pbDlDqrXa3RUcYt8twAgxw5VBIsen3BNfinSL
UgScm9uCo33VjnSMy0kEKl+EixpnN68BXx3jrt9miHd/sXNiL0/U6X5AFZywwp87
t6ULuwUJmCpWGr81zJx6LQ1L2kwVBv69BRbiVP6O8FpUBRhOhHBdiACQ12jnJ7E2
Y5VcxBGRbza8scG/MgkqIX6c01C7XiPSshxIQGj3pleK9llSPcWRKTgkbs363kk4
NSUQVrjjpjHO23GCnYgUVg7Fby8QElZBxw+ih0/Z65BStZkG9k/QbwMRkeDbF5Pr
jyRScbpimOJq717iJZdL9kblo7JOQ+DSRP32As+1HYhH2cwRotRXjK0gl2QQwqdM
A9DSKbi+fLbgu217DpH/pPuQVLcaA72WOs4CnnqYt9zN0yissanvQJGszS+Px1TL
oZWJ5sQy2TnyxBbZukBXg3cMWKFf3DAU9HMDUxz/RvOHoHXnwjdCflpfg63uLQbE
JZJKNczefMQsUiNQuiPZxzcG60zCzLnJVh4YEJUt088wQvHP1kl5uADQyEzBqKnr
G7o/ljIfAPUKa0ahZBRY257O5nVyE/beu/OPxm6EAoNX5+FRJzEUADr3JOWkZIFM
W6bcWGz6OodWyjupm2rLvYmSvTcnuj8Eu2SqqL8vWK0zyQYnnvTMqv50ZzL2RniC
xObNF4n3Kub+3VrCPHgUSzJ+J3xwEN4Y70t07r7wNfsupvfvdAVhWxI8PCSFdgYa
J+CQa0tmDqE1OGwHTtdzHbAjTFSPISIJohqcHsfXHFNs+DNSn8fUCejHfsLbmoZ5
PLIHfbbIHY1reW5sez2V+nP9r6EnC9VP8vdIjlzFouK9BKk5Mzsd4MJIDwv3mtgK
wJRsdKw3uTjr4ThspyPFVo+xffvf2AZ904tXKx9CwPv3XfhhITTBRB6mdu3qV5iA
w+OBSmv4u+qEUB1C/8jQa7bLYDeAm4ur9hI6H5+cP3mXXqKZHvg8xV6Mz9MZSztU
KvSC8D/QBsy4iPn6Rx1oMYBCDuQrDmlGar2L3hb7WvKrqG2n2MjsEnv4x+vCkyhE
guhzd4IvXJg/Aq94cSphYcPOBp3H8KAB7SszGtnykS2qAXnD9Vw4+Mb20Qco9jRf
RowQALaY1gu0zmFnT2/kZW+vDGE6TePN2AsA6pw+32MwcdXQmjtJdew70y419off
rnRV0W5MutKzCX/DE5c4RIHDrlqbSpgDvqQh26fTzmhTNXm1WYMI5a7YJfD+QM4M
YjBcBIKvYkzC3P+1EhZPswjn+/0DdEemNSuRvNqF93SRcL5RLRJH6eVBhdKaKu6M
oXVgyc0Dkr6Prr7DKWKPSs1sB/aHjpxTUpCBioOVUUx5lAhuXjVXT+Nd8/5bnLoH
iw5B+UmBU444zO5AW2imHW9KO43sL1DYE+t5QCZaEzayfSejAiNoRF/zEMNXdE6/
SOEZKxtACBtSUWD/whLZjxSqNT1QPgVk8vfbKZn3kGiP8dwl//7W/eNQax3Nni/h
s5UMsIAJE+D4i8WAtEPTYdqFYmmHdTQkSP5zqTfM6917gjRcZUhIeAG86ZUHVduL
kAMIhYfdfQVdkmgWstTcrBVG7GzTHFkKLVrtm1R1i5OJDQdsxUV2aJEsOgDGJdOp
Lk3Q5KGz0QXUOoKU1S4vSnyJoNx9vXI07MJQQGAZaqpEmfAg27CNvI6IvMAzdClt
JfBylYwjSmjQTFQDAxrhvYwGor8f4IxfOFXyMvEXEEl8lTYfhMIgO7uohvGCI0d8
Ug3MRLj9KuWmoq22SN8s4zmRCzotgbDDAZQbmaKaDXWXb5MhGcKAKg6be/vTKq9p
scRYmS2If7o/oCDebwnY63hojBXYgblUgDEpP+VvWzJUOfeqa86l+JRzLuzVvLAr
ym516TU1wY/VA/v9GMvT4vEyUxySY9dZde/s+rtYfgtPgmflBN6yuTREn9bmyXDz
dlfF5afixV67FS1BSEDtu/oL+g4BqduTLQZ93wMBmWpv4XcIcDQzUC41A1VVQoW9
gIs7qNQciFkIpXrk1WeZo8a0J8GYqUigkmynXt0CCUTAJA4Fas2nGAu24gzWBRM9
iPJWpX5xAto0xuy+cxaXvGKG+HBnaMH4PLEOkiRKSWZshhuzi3b1jzXFNWTm2xJJ
N6MDzqndxrDTy2VFPZ3AHGkXrHTGbX9t3JXaFGRU00ypijV8qRF5zvjlQ95x54p+
NyPY+PaMVOzJZRLjPX3wjOm/QwzlrOowtlv7Nk0MUgPOV7ev+FE1Op5mrucZ7ehI
dGtKc1bdYwkl2/O+iurN/c1LNwOUczyk5FhF3XcoS2vkEfoTpZb+Vjvbl6GJrUpf
H/hAAO3DtDTePkfMfElBGhTgHOBUazgUi0GX5ZoMEs3DcFo5e6AagPVTtRK0y1B5
mww7IDJXbN0Q4uk06xah+7BNc6OJT6Ra9oxsFiYyrs1S2AI1KdpcGpztkZZJuJKJ
7zGYJ//iQSv20PyeN9RQsqx+SqrD8UeeX+Wy0XRZXB0i0I3H2HR8OeOvTb0b8zB2
dMF+MBSPVQhsW02ufM1JaE+ZtDfDkefhSwvKaogJMu0TiLmhaDyKHxmvo867jYoW
ueyVZdSDqI+r5MEjoF044CukYuKHD1k07dFwpqBMrqnStiQsUmms8EHXX4bu+7Al
iyPn/H5FVvKaEgn7JDhBxsED1E9BK9tG/qPOtTcZ04s3OdMBSgd6xj9dRNjub8sJ
/9kNcNF1YxjisXbh9lqod2pYCqqb/JpKDQmkKs7ycB+cUoA4Gabt886FqLbjTpdd
UtguLjdV/GolOc1JryQwgoegmoAvHR3Hj0fkLsJxZ5K+vwTG1yzBUbvEiJCL6YF9
41vIbGZwyBc9BivgNaA/WHVESqNdjcHIEX02HLOeAPDJnkdA+nPrz2edJleVmXXs
EB4pNlrMylMwLSuhYBJFitFYhiPELWlJ2R8bHpNzt98C4UWWhKfOSeEUajyAZcnl
6IrPGBPGajgvI/6e76uE0l2/WdYJlsYMc41nayyh85fXY5MVGoZB7mgWrZjL6L90
8sA3wdrLH1mp880bcveubADgM+ttPaaA7nVWE59ZwKujsaylL2rDADIJ8Y63iLIG
Q/VES4FVBmKJ1/JWhUVwNIwI+BVfFVcXAZ0DhPsrN3SPeF8nf9K8TWwd4GK21OR6
GwUuyBeEKBfw7m26EIl1XTb8LLU0SRCdDZDURHKagwuTcn5pasW4HyPNn76NdPJ+
S2JtpACJX46Y37F00NZv8ZLH/Ecp1Kz+b4xJxS/avpw8DPGKaOYUoYCbX7VuP8Py
QEWniFzwulAWXTn0C01qpKoT/xVIyi7s5M6po0z2uI4G05mg3sWRv61Hilt13d1/
liRWL1rr6ULCTC3a+W6zeHjRUKD/uAEUpJedUTpFZLJekA9Ao/nOR9ROG10fm5eL
rZXIaVnXOi/DlQ7Y+iJYt35R4CL/k/Kscrz8DSApngAikShEPTDdK/xZVupXn6Q9
HuMMnGpVXSZCPyVfQoiiSM/ennvenuvqlgGcmfCXh5ErJns1s5DzjynIP3p5FmHg
sSrzS6ffZKn6lno73/ddYZPL8OlHEaqVyhJnBW+qa6oM6cW1n9xIB6OnSdpQnkzH
AeDTXAPl20eQkV2gR+jMdn+oQwEcZ5unPfQqD7ogOfNKCMj0WPsnEoZQatUxAqs1
3d/Q0+WC+0XsaPJGm7UdBUD08TKTgiv2dLuiFz2ZmEdx3YHT/Qat7Z7MFdCNi7mD
gSm8tI9jaU/BUqRIWwARbVduvvoGvt3Fo2S5ZO05eug2QPbO+35ccvUaJcE5SsG7
CMHBblPtLidWkwMG4iruKS90s+lmjh4b9j1EqQxHnvFhMjbaZIc5R+NIlDaQtwjJ
mZP+afjmsFkAJ5dEjrFiLHKPZ2YwLoqMJ5iSmbDLS11zOBI5pkKbEwUkkjBmIkNY
qmHlUIpqKl2wkrQVwC3wEXJeUWrNteAucbAQcMYPXQZn/tD/3cvhhx7gpVEWbA11
wJjaR286pIV4+qnIkNCIpOEQ4ydIVWlENELh+eKs6aiO/2HHd+7FiMOZF3yW2wnz
3AwUNwdMLfOZmT3ZfXBFp53kgHl71ds97hnq4b8rANjfgFFFR1fSRvrKnvZKi9ZZ
n8Ehm8FFSIYv4D2oaYYhGztZhH0lyaTrKB2c8ODOoslgykTMixUdoVlWct+YlAJS
4BAnxORvi+K5zKSSwew2emTKuUP05G0zpShA8+wBPKxj7C9DJjzcklcDgRd6PQFa
kCcZ91XqOgP8dwq9ERwP6RfHLUExIiXYNjzgCH0Dfr18o82LFq7fOV8UwFxr8EF3
tL/Ivnk2k1JcoUpg93TDWM/zrC4J4k/ZsYEIK2j/s37anc+Mr5vwnXAVS2q88Tgl
rgusIKDZc+2SEUxJkHYQ4rnlOxviRS8fopcAFnaiRlCQe1+1S9jMy/e9J2XHt6zH
Is3IpL5IRFw7PaSMwBhbRtiISiUxopH4VVtS+pEP2zE+Qs62SaDDc39RY62CyAGj
okF4HzpDTmigCqvu6yukFwlgO33KC+u0fjh81AUz/y0/uoJqBodtCxJt4N5gepgy
27PCWAaNbwrWOgdV9pMTdzcKxNY8seCnwOXzi1CCuU76CcgxOdf1uXdnYPmf32A8
gLZCk2+boIuedxHUCqfY5uUswCBcEd1KriQo9OuAYW8y1zvRIN3rM1+4YKq8DFIK
ozchHc8F7mDLJ1nPR9+ixaR5YsIu2EQzI/Ugr8BcWBzoNeNIkxtrXdtF4hKD3jEp
d3SF7ig6lUyEUR/YLgBqYep4yLiAca0SDhtTCUAP1kWj3BGbsgSD+v+eI0/39Zs2
C4q6zKj+Lus2rF2i5GQc7H6rLPnm84paHlUjiqBaDSG4hvDGEtbaAuYMiTG0B85e
DKgFhos/JC3YJU9oHF18cucIGOx4q9I6pJZd2dCgBNm0gngnpEtA8t4p/jAfziRy
QNRS9cRBSVPg8tBBRLjwqaR1nsFWjpvZ6lMdj459PgQ0bFZPlB+ighdNEEP6NIHX
kUFoy29yBrNpL9sqmfdDvPi4QkTcQA+kDN1pReyrnDVfwPPitMl7s55iP4RrI0Lg
ha201+/DgAIHym7yvInpqYvoPaQtMyaIFQHC52drkSPTfVCm+wJWyRYzDPGlainD
ouPk3PGAjrul13LJV0QxqXYRUyxCa/OlfuoRg3H9NPI6iCe4u3Lco3pUlb5InT/X
4iH2OCs1+6e/uwJbKyV4gLmIe/CZ5sNCZDUKObMGQyg8HMtsnF/AORCxOZUntqiZ
URStN4VqN1S1n6bvGV7Kc5iiKqGKQtrjEo3ZIkwD4yp8bDOPGKBjlX3qTo0wVESp
dNn/tnUod/FPNHuzBfovyISilyBuynAT9eAus+F8zhZa4Wl4lVHS22hQ7VJYjkbk
CnXt3HtttD3cxYMsfpHzN4iP4Bh/TX4VUpPghsChITItXlykF75pr8NESI7SSgxe
pmrzRwaXsElF/+kC63hUOfTr9KGTqkl/waHooSduEcmfGC5W6OFvxfzp9YqDXjCP
7iYLY7tUXK7qOq7jANhHs3qZisdrrUmjEDy+Tm/KOeDqkiqbbyxo2TpxJxQ7BG6M
IcPSbWJJp2LlsvC6P4WyZXy1CSJMzGw4iHGwT9PYIfrrD413/LWCp8sm7uuFwFrO
0R0FVmW9LXIOSs2pfRf1n3RGj/sHVtWM+K7g+SD1edE5/iQdMmKZV6KmIMT97vuQ
UWbIGDEXF9W9mV6xfFMf/CZsxv7QREWJa8tPKBYAuQUaj+L4jaL6he+G3dbJyTmu
Yp9IMR9h7WD0NzQflBlxu06jtkf67iAIb+7aMP0pX1gCFEt2/OoMhUrLqvkUnYDr
XpQ86mvsEeI7Yo9SlFv+sB0SPGT53KN5ss+lEMkSJdGjqcL/eCJn3Dl4Q/qMH4aJ
kfI10/XljjxbbuzJ5wWKE2UamE8n9exLa+/Pen0EH2QvfX/qIdMkxwdpDxQNgUZs
w2ZdoblWNdis1t3Tk7y6SqKtl1E8dbvi6Xl9rg0qifx3k/TmUAtl0ohOSyObPcLP
XUXFeJ9gaKwSyXiqwsOr+SAY86/Oitp09WcX2Aqzaxrm98Jn7TSv8SZP2u7ZrmSq
TcxhjYQhPmwrUCM6f5t6RaJqj1ruyMwlIxX/jGoLWPeNnOUhEj2/PGu6d3UeCVHW
ZfQkBGLgjZy7e0B2IHu9y7XyVBhDwpFtGblbYUQiWsb5oUTL06qFtLZGAhZodirU
By4WBNfbAiaJb9pJN0Q9YAuNbSgj9BGbqD5vAXqABR1LUlBsF9Uo1b3vhjEZteBh
YP+n5SsmEJP1hFdQR3cROd6nTD9sdtGxroKGvgaP2f+AfJffFG1la1cDDP7jhsIX
uBBeSh1zu9L2BoVr8t8HxJe1GgqYwVzjDzLEf9P/dAasADuaVvlRLNvdLJ/EwH7d
5h9E93KYvSQybTNQxp3o8qq+EYdGG+Dzsw+uUJvBt7o62GfwfaLckf+RqWLCH2o7
mtUc7C1e3sjzUMWSQbZYJe7V/z+QU5hMc+5Y6TEMpxYsEZHlPswXcZAnpKCIA83F
WrZ9uOjrRT8i504VZEU759R8vl3oXJi31t3jr1VSz0w0c5wGVeqb5TBiJjdUWw6X
hkRvrR6CZ7/0fe8zY2Z2nB0IelynDC98C+jUn4UxFxufsZdAsuQViPQdz2wDWH+G
IMIFOlRwVoSFxR4ZCEJsDWeq613qcG41w9zHGXg4tHSeMda6CfqSbS1rB1HIZuN6
+YWU6s8z1ZxvC+aCXaryEyrwQpA6xakwbdCnwiuIpbJpgfmGxEVmMlifmmCGIyNx
MsKmXT8Ys6wCSX1ons4UYwOFUvn3n5frxK3sDzNyNcZ0XfbF9HvI4SYvqms8ahcC
YFVX6Fqwk2PK3TMW/KCK2g00IQmZ1oaKLLyXV25pnlyp3eWokc+e6mwCDZxv90k3
XzllOKStWqfzWdQVXmygULjRJ3prxTlKs3SG0OiaKg43W4Ix43asji0Qh+sn7zee
/YDoBjJnymkLzYwLDydzH/M91pnrGRAlesZXF35dTPRn3m1rjPLQJRK6HmdC1l6E
nKwGZH/9Ep73gieeJNofOdOrKinr9zV9oK89hsGxUkz6jQw20Lh9eFXa3cqMTN+c
NCN/g7K/BCH2jf9C/bG/CaPCf94m1/RKmsDTdmuOxLqgmV2ukKubioEMTiEq04dy
BmagX+PNVaN54KIkkb6Ad7m4PJllMN9WKHE3hSx5iBgM4uyECDuCKkHs/stYznp3
LYObzvROMmOjcqq0DQrMTYPqtDSM4GPWFJ4n0em62tm0/p8pDYx+zoF0fcB8W/UM
Z2hK425DqaotkacvQTFAnmqnSftW0Wu1vuS3BSeJIlbFo8ChyemD8sgZGxdc7LIS
7mVfb3MPpQkyjMbEO7C7eyRTAHaGy3+7KLQO/0OJ/WEZ97neqpSBXZW+ZNGIQEEs
DTy6tBvG1gIVaa3z27SDW8Cfwdv45BXTbxdn0/jOfuzz9/HR7um8Kcm04/dulUzC
mjbjdDEW4T9DXdVHMfxCnNbqopGCes+gQbmlqKUUaiJOZ2+Pu/bCzZh6rMg8O48r
AhzKgBH0vRFFo6oHLzNdV1QNzX6x+C2DE89x3OHLQbwx7gZD5vOMLxlWpt6pHSVM
qIOPwXPqHJhwmCRXKgEjrFzrMGGuSI5MKA7PcNvkCv3hOvjsptBHios4ud1/PjVD
ZqsIt1C+4UMvf10Ukq1ebwupieuxy/CWb82osYu1PNsl8c7AZmZtyC3IONkHou2+
lqiO5hncepyVhFzer+iI1wBbj8PCILb92xuxSvdX3UTIpXfSaf46HqWKg2kwZIYS
6/dpYCzpKzzrZnS0zeCgGYTZAyTcpwQKAgcYBDCTirdqx3eyomeCsrWIJ4XcBYzY
ZNPniQcRoE50PjW+GEwbCDwi4J/hANufvhYENXWwN3+RPjtPcR53gnxRdA9bSYiG
ViiLqcQuNrQ7S+lInnWG+lE/WYyVz+1pFz1ktUx7w1uqzM4F/nFfNdGG7RmHU44p
5a3g+juTJ4/vzAN3mKZPbKmMH1PUzyrwYklLV08NRGDkEapGVRaayEfNiRoozGU4
BDIJN5ngXOfqvOXBoRf1VuXpy7POGcJQy9e9sgZP9P4R83W/gHIqcPjRYjvAxK5n
9jktPyXRbPpO1ZfZEkVX5JXCDAhVDhXjSiTl6SBC0zI7JS5u/boyWcRZScN8D1EF
j1ts/Ubj2y0Ld38hHLx9DAKF1E9vUI01QaXwYxui/gIT5ico2KnEvuI0CZJAyG0T
N5+igsWELocfG+0UPDwUVNpVlizUCYy5IEmnrq1+plHOcxp1/ldO1a1nn6jQHf+F
cmHXJjX/7L2Y9Q8MCtYEHgaKraYI4I3iVk0i4i27OoxqkHFkxnSb0AN7fHcCaK3T
BcX68i0sohTkkDuCBgOf6OsRveQg+gaJKipDbdqGTU4YAzxO8AFEGIHQ+sMAVLNJ
RDKZw/QqtiLYNVal7vMGZ3xfzQfHgE/ftOB+OvUWearD+dLf5xyAKGwNs3VTBodE
xH0IIll9C9QirPhr040yhNRXkEBYeTEf8l1EoQEBOwuOOvuTASfHgnTB/A350pRJ
r3R6KRTIs9k3Dfph6BDSOY2oBYwCCpTYmYiP6+dMgVf1uBq44YK2GYZWefQlqlDX
l10avIoQOzDG90Qw2jlNVjnsHmYwPa76YTZUPvyjJ2rZP38vG3Ct6sldlSScoWIC
ZYkn7FJvXmwUER6Ro3mDoPN4drsfRgfyQfljQClRtqT8IK9nJtvgQLX76WwnNJ0C
r7wrb9+oHYThl2QjO85qLJn8e/BF6x14aqYc+TaqdBWjVGHOpbnxeomqNhCtIS9b
Jrgkl1lA5fm3bRbAeTz4dISj8mJ2ToJF49fQgrR+ZYAKwio7qvnYDnSFOsnDl79r
Vyv+o7INiES+KTYx3yUPggD48jh+pXgvU3Uj0SNqSFNzMJjAu2SrlO0uUNpEP4VK
U7h8eQxnup9I7K+gG0lTyJcDSw1x2qzwfeEtQBMj/ZtWTdTbYgxC94lSGeDASJHG
tt41cI4gMwkuGXqSSLNRhL9yXFw2zr+AGY4uK/DQVyTd0tYUEHEV/jIw314Dv/U1
5dkcrk3VSaPvtsktnMPamhYvbXWcuxNIDky+meJNcZgd2wUZRajo3959Gq1qyYbU
6trFNkJUS07Skj0QhQP1rawEWpIaAhYHLp5G3k0RMUbxoR38grVm0sH3tJ2MWClw
0R0zccNeh43uNhM8i0CiEUtvjmj1501jjNfHwawm5GEX18bljvCiwdAn0pj9jKEm
dZxmPNRf46hawK2MYcQhJwwhg1sAuF1rpVFUrdkPZX2nQKleafWfLZEj2GVtGF0Q
YgiImFEXY4ARpffiW57F2+Q58780CLRhe3xcLT7UX6OgTXK/xe6yUwhi7pk7M5RQ
aMaCbwFHginD5GML6YeVqueU7wkECS+N3FlFegd/5M7PfTGz6/vzMS7F6/bMSdJ5
wkuh6PU0QKFH7rI2YXXP+hIIRMPO/qmRA1pEMZUV1zlbu1wE1I91U107k+NwP0w9
jmkmaUB6AR1DGw53JFSWDRKCuJz1Pl9NkQKVrB7EqtLPIBD8OeyOjGfV+DLiht6v
7fyzZpvZcrPeLcEV/WO8ldGgAUkCirKXNzRfKNMwU+vZHya7Wk212glpNaqLvAp5
wAqrsYthCsQ0wAojEnLdAn0xeXx7xwKLMUoVPDOUO3zspEXnJOu2HgvXHN2xABHp
dKD7O+3RQnUrght1pkZ+Pr45Kz/7HNBIJ6rNtsNHewe5N4bZgFdHoLzJxumYL5O0
8MLW5ELB8KvifHQAbyjH8w45FsNho80A5ZUBEbisQBf5LqoqnOJ96PWPqto8oah7
b3KpCt6bDXiBTFzg7UQdoxu6BembfE8vrobEjqz9gqR48WfdXB2+A/xZryTEO/Pj
7gmi56lYVx+8VQSkKMSRpAqKnwAaH+3sgFsVr14zSBmBnVe0CWT5LLglnPYNp4Gh
KY9xMafHyxltjKyj10kqASu9ijRQYBRM5nkgqgFeQmCMRmbYlQHRfBJmjOJ5cZ43
nUganEfsBM0NL7mu+JTVynQ23pC8k9zWHRP6dxdrexf/CqBtgnbQvWg9M2F6xHah
DnRd1GhiHoZ13g8DhKjzOnyt/8O4DHNzd/eOQNxFu6Z8NSDMxMXPDp8mD72CDBK8
WmCyr8Z00Bn3TZMAaIh3Im0FeSUjLiOdRHXnwdO/aJ+jApkI0fie469Z+8ZxG+hO
ZRp9ie5yQ2nD2vw3uAMMV7Wj5u561z4mf+GAlPeZljQJV2bqPFXn3M3/bCvdugiK
4KcbA8mR/OyYyp1aT4FFUIvxgsgjb+aPEGvXP/Ubv0vqUwihH1H5vd2+5KIoH7t1
gFEgKXyoD0a58MLlGLJBW+2/5XLr7J3RMMUm2m8ofTV3f0MKU7A8K73UIiHLAdX7
uP0VsEUvl8vfd7n8sbI3X2y00wkkI19oyd8nKknhx6ihRdykbx9Tfx5bY1OPVdTG
EBYbb8wxk0H4DVBMvFRFLw05BJwbAuSIhl1CDM66/6F01IP9mFpIwUcZvdIOzfPJ
jVJhxGwp4Ufncy04p77c52FIpwxNOFEtouOxShmdkll4+6e+S+B5AGbR7QPPN0Y+
ekOyR/bkxQ3HyDRiKugK02KMN/LtboT+wxLfFJ2IxahJc/jJ8qOSAJDc2Xg5WS9F
MQIzNya5y+62nLIxl8TuptF8N1C4TwB9RUvs/ncL27LxHODBnOIntyq4IX52OYfR
fJtb4ZsOc0OT01Ufcs+jG6PgD3M1JEHSKd7WDdlF7YoRectA6NkdeDbzab41eoVv
ROAxzEY/ceiaWkxvmT3lu4gWPP7v6Ig9rZJtj+zeUOrv9r8FKQR4EQDyIOp59kA1
2KT4DCd20y8WMgPZMZgPS1Vu7TPdlVwyXe+2y7g5q5Kjs8UIPzXd5n0deYdPLSgh
bub9rLXw9/Sp77yEphh4kc6LmVELh12pPBC074LVnUIkYjxMvgPhGjjcHhzeBx8U
7sEW/JKvMZqs8USW7JfKbj0UMzGD8ZQVPIoSFpDLpyRnoboGgmGMySUuRMG9k7ew
lUxoQ36dO1cQIqnULB/C+sncfrzjOYov/k5CfVOCJw0QX8HkJ00pdVcLltP/MHTJ
epbbmVHhXV+q/fV75osMRuV4XMBCLPwaFLcNpvGk3Z8BgWBdcAKGoZFjoUt5K481
51CbJcto3LZwBRbLsAPQwb46XwyVGcilg8dOYhMD8RZ5D9TEz67bmiVV166IrI7m
T22I9r/hBypUmY1JQBOKWGA7gZuiFVE4fqz6eiqT+Euu6Oj/35jzH0yOiDWN2TVf
49Z0X8x9v95YRfLk9vObo5QBb0atYO+nZP6hy0qTt7uzzMJKuQKsQIYRWljjmIHF
lRCxegvrvuTPxvhpaD5vUIg0Jjt/uM/5rqTFRSAIgclkK3f3hjS0RUjhuR5AYB0D
j76X4tVEZ6TPBME8lX0iHDuAgdrPrAAx6uVd88ZzXrZ0j2ilY2dlqj95XDa44oOd
nBD7ejHeeD5TXULHFFUFRIUZh8VuVNSKtaZzZ+Vs96vMRsyc7C8AObPK8+PzncVf
6xflXALo8I7gfxdAwQg4P2kzati6/2vZ4XNBenTHA4NL99SWeeHy/6OhdhMQS4Nd
PRpW79zHfNl+9yzAV2G5pHzokNYMCL4q8j2SnzYpWmBuOnkyY+yha7RsPdkzR34c
KPxjc1JjyVf/mLB0ORVjZzeQWhZ9U3tPgKC3HAobfl2NAPxYkXcnvFqBhZhBw1iJ
oJOgWeC6VYI81tfM+1lL/lybkRFHpKd62uxs2i5f38Z/F0X6u3aEnNSBDGP5ojd6
9me7lvI9LnPGCZ9PAEQ9YcLlqLQgofMH7mhN2QltPxKu5YnYgt8mL/gvwUSjoBji
Vw3dVEtTnePRK1z0Skvr0sWST5bxdDMtjN/vUGmop8BqpgAX38BVsN/PxDpDk7gU
qEQhllczzsD+H+mNKRSVCgGClJnjKnzg8a0bfi7Z+kPdU+6etOPxlZGsC3Y74fiU
WRM56luVFvetHAX/DEuEeL71JMB7bs8vxlmFwyaMSl5cIaEJ+FghPZRudFdA2yRz
cFn1nixqzXCR6GU+uR+WS4PfKBfBpxZ+7OCQnExVOHPCBO5j7CveIUfcKoRykwqO
Fgh8tNsqEvP8DOCf+9lCd097W2LJOoLCk3CMxTSLx4p3NQciVLQRxx5lMBw8DwUA
NmrWHwGqGdYMpTEgjDPfNjbXyJyPgFWBlKEpRcYkP+CmxqHlLtv6SLyYUqDFkYxd
3UQM0hOtryCz+vOIX29yN8qduH/jPy8szC7AG8yX9EUswKoAciECwjCUisahfhPf
d/UbmmuNf0tPFrhOxz2NlN6/hEzOGZ0A9Fn2X2cvvWAJy/lQvZtzvGi4Gaxryf+F
TiEomsEYHooNnk0P1seZkmBxl3GKXn9Y50VJopK2aM2NPl/Zg/belA73I3kLNlwI
BULF2xmplWjbYfV2B4RXnQL+O5fAsXa1zR4CKXP+Y5lygwRGshjAOaakzu5kfxJh
zLhTUxUCbVsTFJefFOEojUo/6qw6ywntVbntt76Ig4e1exrZtBFeaLIZXGqEucTb
v3fK6E+9UoTlfYy7CwcmcSRWynKNZSsL7ATS5NPIGk5TbSWnC2oxPMULsNJQSAAv
KkNSpifX5zTAqeNcLSIppuCALsj0Ry0j5NOyCYXabaYcDStGMdpSHSrGfkFE+5tl
y4P7p2CCFs+UWyT9GXkFHBpy73sYaGgqMRpZkJRkpV+wdQzWl7wjZZINgRrj3DLN
QcHu7h/ZXUbkP74jOrynfUbS3i1c2iYVkUaCno4zYL3BaUt0mAdBeYhqH0X+sYWl
n6Y43fvPJ84y6IYOt9uLBJ4UfEmnk03Fz3PwdtJiivIsvBZYEYMdva9zJrBzai+U
H0LwSOFK87wXgoj92e1Gx8XN+AQ2tELKo274kFTRKpRfiAFjrOldLlS2ZWIyUW8t
B4dpr735QmT2TB2EzYQcD9noH/80k/3s0YTIw3/j+F+bklFQaGOh5aFK2EKovKbm
a69DgGiR5Xzjh9Y9vOUIbVGcC6ObecS/E8nSeXAzZ8k29GShMME+WNfc+pv3bGUr
Nyvt5RUwKDsSNdgnkzPzmq4T9nYJvM2uGIykNG/8aQ1pj+uI6KWEHzoWU/gNCoXQ
UHKiAJXOt80ofxtJqjJWw60ia+b4UME/DHwcNZK6cOZJ0DajC4ssvy0NE2rZiVmH
GmcGcvq2SaqhmvHe+ipzxcgNQCSaKWLOMzB9BTnSA5O8e+36r8TV/jRCtnJdVE2i
IXKjqqyy3cCOsXupJG1lD/RaK294SyGZdEcWfFFrktBF/0zkVV8wBYghyvEF3WbY
SYFkC/asVQcZ6yaO+mMOQQIqDDs3VzkWSqRZnfV7KqBJ5eVh6fJ+YATCDIYrFbRb
LfrNw7/Iz/cukbwl7kczTZT7OJndkGrQsa+vg98uwEvNAgEOKXPtGwVgN07cDSDb
j+kZx5tjOLTWvRgVZe5jYx7pURfk9GaTd1wSgokIT5/SgxAfWuq38IO6lkwyC2uu
qIbSWzEFC5Z5tb56gB6yrgHhPHvI6afObijpCJrqrMVmgEcsvly/fUWWnAastkG3
ljWdeQ9rDQwhd8DjGESjeYg1SEltwwP4ZMBKynyC+kkKe6bc/Cty0N+0LEhqlidx
CKb8Iu8tJTtfPWBDurr1Iu5z/7RFAK5ZhuSQfYiF4/6O4+R0NYHpkLNPftHEPlfh
zhyC+7qGqeRfDFa4eSdW+1sl1bQhWvgLNv0/PPnupKKifh2r+tXEebMyxs7WbOon
F6U2I2L8NIWAi8YoZ2xs84Z3lNbbPfNdEzdVyff9QTJtCsHn3Y5N49vanIBYdImW
xDFNdos1jfDFKUAIA32FF9frZAAFmeXcGjx902oiUWJEwr5QI2jiC5Iarokd8jg5
j7YjhXM+vD6R6UZyH3kUfG5lASMoxPDodOlGZJpU8BHCZZR6SglCn4nmoH4QIrK4
70xDm+MGeqzU4gWKnbnnlXgYYb/pObcvRzvFBBGBCjHCF15m6w79pPcclkyRx63d
qDY6t2y6s7ltebEHfuSg77CvxmC8HxxIJxEeb0FEiTeinUsJLH/qq3NYZax7E37t
cKhrwcLkWmOy6AxvaTRL5hdiITp1ZQKqM2EUulK5AOpIWMAR9FNHgUVpf1EzxDm9
pn6Fxtv6UCL5hWTjlPNtWMRnsgad/HXQPL9NgCsHOgBIkCz1MROz512Cw7SbFSNB
2LUVdrx443qJXHz5wL7qurQKlehxmb47PkOfZFapsdI8RLSMYWRsWEfRgrg5ZIeL
UcgqAIQcfPLOqMS02crpsCTt/PCoJTrSjKOMzizlw2hNFiBFOsv7eoNP+2sk3XWI
bxug1JEEmxaIR2KVfSvVAPVBbDKcCFgU0NcWjPeWG/R3TprVSdNofmw+ag3zV26S
yizHwAOy5pyrIi53bDMRneehvChyOgp4Hdhsx8GEYrmfB/Yj7RY/J6cO1eo3kcNL
7GSD+qBaqnsxxpiYQf+gfSj1IT346ZvT0JoUdhfXJb7SuRlVxIyGSBfhF8I4L/cx
+ejCErd4UgVD1YeN5qNUvHPCXxRcE+6AT9rlrduKP/DyGBdpOwAWW2M7ZnqdC1hg
zj66YjC9GxlL1hDpE41Vx5u2/lkD1J7PLSx/nHirckyo4ARDZ7FuchYj0wKH5Kcs
DlIjnWjJpSs8yTKuYib1xa3huiMDTVolxIU1id4M4T/mcINtsTQbcQyQKiWow9KL
PbCJqhi2KSUfHPuU9LuRvn24mRJz3bA9r7nOvju6bvIsx2QPmMKHJ2UAYywyylRi
0MrX8ReAgwIJFo0qbeqcS6Qd8ATmyOPnvXX4C9Y0vZU4TqnmcUYq2qAdryUUiPyQ
GMSvpkrfn9mfWrzkFAIxj+D3UM+s8CjKJa+fuaSlxexCimCP3W+QpXiC/km9SSq/
3scX7lpzt5rIOQOOU6pxSQtH3EifOCVgRsEN1EoSa2KwmNUJmhTBsLSxzjBfYuNx
8V7Uzv4RvfM1tR/oq590u8pjrCfeBsVgPaLNUTwt6JKYZLv1S4KvO9PNcRuqVsQi
OI0CKTWMgO6h7lPYRmngkJWXx8sGt8kjIXjAOHOCRh+0U2iIaEFscJkzLymcFriG
NUEvEEyiJ3L4hYp9NtMpw0H9y5/w19I7m3sawkNLBe5rQ2J8krGisupMb+Ni3YGd
nMcb/DjJqYPgQd0Z67d76JXwzRlwKVKdgr69xF4cwTWeMO2BbgFDuVljUHDJ7kS3
bQj3km4tdPLU5SIVjDFh+6Kr8bhYnXe4B2GUP/u5l22kjWgRAbUpTGHiWvBTBY0J
FG6HJr+yqeglp8a2DgFCg7yIk5GtGw2aMonHJ2sZn8b+U+/JO9cuGqdoDUGMmiGv
YfBV3XKocNHZpC7CNpNBBqap/1UR0ke7E1xZBX9AZ4FCeCYFfCEoMBow+tMTAzde
HTQKiC/ZSF0Uxvb/skDMSPWOL8A3/2Na6a0Nz1QnGDstnehuUDyThx/YnAg4KljI
Iow5+zS2SUSrxqfOnuU0hC0HmvrpK4iUCHkmEaqdELsRq9aE2mfraRrFn7FzGca3
9t+Yei+M0D9AlZInSWaDbjAFZ4yzz1IZio1CdZaJk9GJfRoN9XrXRp6ApO2vcMn6
L5TQBK3e05e3j5+Ebggm6Y8bOp3j9oUrm6N9e2oBPB4n497k+agVENiN0BVvCrMT
YTxfEnyJ2xYro4aUsbqZ8j+Wpd+AnO/irXw8mYPQqUrYvsEcRw2tLvae8L7SXFU4
Es3CHURTL9jJ4/XaIfGPQFCiCOWQSwFbmNohBv3t/gItU0qXqoIAcv6FHmxaoK0l
qtUQ5eTOMAF0SAMSgLIew1qPsBgeYasx/MKzwqkAMy3rtI33hlossTD30cHVCKOp
uR7bfuBjxB4KZPDPbHofxDrm/lBSn3XF/Fny73Yz6aCgxYtpHmLLKoX6Aqnj7vNF
4SOSUfVIovRL4Mi0jH0FBzR/wasgmzP5bh3szEMEBcrp8X2GbFvLZyHvmI8r2hDe
GYPvynxvs1MrCr3ccWhxU8zV8KFHKiUgCELHmMTlQy0JQIB0jiebi0Wlh+8Us8/U
H1oeR464YICr/F0SGyjAKLIsGK1VX2ED8C6ZHoXaZdZrghow++1djEhhEWOvubPV
+u3XT8jwG3incDatO5FU9xBc/IInJWkUKTTvbHepmu7XWVLWL5tAWohu86pSCmjy
DfnxPHyTdmh1eIojA+iErNcb+efKdkmX3EX5n/yyCLzYQqy962FCRUW62ASnvfJy
/d3P5aWZS1bmtF8E4O8BQj14lqE5mw9yAIdZUfKoBl1ncDU9YxD2dtsbWK5mNsyS
YiUk/C4G9yGThjzW/iCQMZH95AQwt/J/14HfUkZDkqvQDlftToisZHEbMkDbDNfC
T1IfT6LRFCeJgf6tUGSFIBkhRodub+2KosINpqCPkwCNhjypM338vm9imDOXctTC
qNRMomoB2ath9zQF5EFNFWJkk76iyTIuVE4iXAb2xyNbNQYNb1vFOMF2rCzklx3d
RSl5OOetjfFVKlroNRsxqxNsObmpqljntT8QVQGV6c5/4ic5qSOsxZYSC3VLjo+Q
jLK7ZXQ2DpyYZaPfP5xDzXQEIj236l2JS/m5Z8ThyknxhCgHCEkOVPsKERvFHtRf
uXz3ouDxl8/JI45CinPO8Uk58H6FYkFdyymh476449RQe2Z1llH/wzLTX82VGJHF
/Sn7VXAjvmE6Bwe3ZdqtMPaQAhgf/0nazni+G+9u3KY6krqX1Xu/Dj3R5kTP3COx
M29w4DGySxYv8iSaGcJ7AjfTwHgk24Oy9rKbzy1akkgAcDClCfAozgq3fRNGzy0e
5tUJp/gkNXeMjDln7aX0BxnDWPvVzFsmf6e1iSoM/Zu3PTqDb30Q3eGmYv3DzuAN
9It4BtyIu1p2j1ZQ0w/FYm+s2aP2Z6lexeNfVwaYmw7UH3mML6nP9Po4eUbJTFHz
BkV6ItCRWtl2wes6QqVjFsmsSwNRCcKCM2UYWbiAJRaRohfbt0Aq6sWiOh32ZjH5
vStHecG/u0VMJuceecFPp8ebL5Ud6GvMxiBVX+1fQ3sQZszGIFjvUv8K5UCR8376
/xPEibNKrIN5g58HgFstkgxLgEBChvOzbQtCzKNKr6nOpGDFk0cqEq2ZtT0vkroM
wxn11j96t5nvrTS9/ngEKkGjt4HknujVuRsTxen5UGxqLkxh9rurun1aEhBE5bbE
zS4sNiRi96LR4AUSRl6ZMUg0tTnpWzHS3zE3gA/+zaVHRfXf9xuqU5dux4llFJhb
C4CTNmTMlnEkyOQE5LxBe9FD943oKLFhZSS0fUkCNDnngNAhg0ktCaixLBfk2XHz
UkinJ+PE/l3zYq4ntJmHMbPXPq0eIyYqDlfLJVdnvagwmElbj0W6PJFXDsj2M3Xz
A7EnSiT74/wpXftQ5rvy1sz/itcH//FWGePP1e6hI7Rg6Daw4AZsBuVId1mXsABi
uQO1m0jL/FnSVF0FWxG9W3GQCPX0eVCHo0zo60Z+O73ZbU2mZ5XD2Nmnumjx+ejj
4AB9bexg4JDNyQ/3jKVUMMrV0wc0PM7U3YWwc8DmG6a0JQqrrMsdm5q5isIcm+aJ
g5W8SiMO0Oo0ZIBg8wIn3dGzL1CTXhiiCMGWxjYBrPbO0nVsPLu6Fdr3D4eT66Rw
4Cwl9c6iJpLA4ykefyizrLR7cT2IrOQCc+9+W/zmWa7mR1uB9O9BqWp994uuD6XR
lASfT/ZzaVKR0IcT30aEb+0vjTmRONCkzBe/KXVtEoWz4TGz3VwxYNYFN+gxg8ed
7JewPQteFpf4ShxOD5AGgr2qkj0lomvBvjkuMfBlOmfoCx/f13YQCNq80kQbLcgw
mcJGcySkTcwgJhN56rg3o1UXZZIuDSWN30OLi1fGPoFBKyVdzcHwRZVM74O2nLNm
zDvyfjZZ81RaGKGAmE0sZY25fQgO4ofIgcSm6eFGPRRjJMABrYbE5xeN2jOiI5Cw
4Ryi/J9GN6PzSJq8DSiuBZJtclbxO70EyqLMyacO5APpm494WBBA189bdv0u7yvk
g+mSrK6GQDWrqGF00Z8RgL/bw5GTzZmtj2J6r4cIbHKVJmAUP3QzJnVZHveMaRfK
ITHZ7JejGPtayT9hBlFzjSXXp5XRy33e0ptvfkLXBbC9ICTkip2gJmeS6SfEdCxZ
nw9YATkWvwpL1bB2JIU+ohIECWbCNz+UWHlgCn147Gl9YX1a8p90ifZ8WFNkDPjd
dRmt+nEO8fT0FN5JAocWaNn1R5lgLR2N/PN4vHwEigwAIyPMdFpJ3fJodTuU7ZF/
MrjeJcQZofeiAeMVNPASiR5jDfnHdKdCDOp/cbr8B3yLVTKLQvDyljKmoZqNIrRI
4J2speV+BLHhEZg8vkqOA/XgusZI2EDcv2L8kzBpK8aqFrbckT4Ax+ZldAhEwnLw
TBZbgdxikneyOgoo9xVkVn4FgHtsmqXabktvAuKcxrt+ZGPNVU/TmxQmYrSJv0PN
jvKRXys2eMC1acY4dSCWoS1sRp8Uzm1H4yzXszkEAlCp+8jpbajtUY5fJEN28FPd
Lsep3QRVOBgvJnqdO8iQjFVKBYd2u4Ya4cMgC/oIUioenmaw6Wd0FOp2fNn7OKIm
yirpWuPXavtTHlHA34Q1q57f1ql4+X6Y7u9CQ6oFsPNcHOK8Uf8b3X517NaIaxpb
a4NZxZklauhwcDBzCkSbCRiXWFMl/ryQwrR5z4GXgyK4HgVkmhmCkj8LaH8YiY9u
TSxwHneOyOI4fNTnWGDTh/z6Dd4/LtLQ6GF+5UjOygpAZLFxYOkztUTDn1S7To/O
bJJgHtAScdXIMTeLMbN0cRrshpdgK57AZa7Gj5ykmgLIjMm1o4No9MvDyMeQzb/S
oOpFMSHq+tnDxLkKRYoDpS1E/toLfppFrLrNDWnJoVUvxQUupULHqab0kDu3bq8K
CRKcFqrOhckPmRmGjgBrhoHucMlnRjG2djKlzsqE2ni6lEWlVN4vId7eZydLfewo
NuBT+kXKb42p0D9xulNB9GLCRrlTmwEO+t8ToCQZKudWA6VZkzCmoiaPwW6jG/Td
oeyTzNPi2Nwq1GYO5xTJ57f1idB2xCP5eHvEMm0rtrFdDJpMoE2HYgya1sOZNxzN
cTM03+zQkP58Uzlwu8bhQDUpELZU9X4681QArtaTGVd68HmtngLQ2WmV2necDosM
2PmVLucRg4zyvqS7ASIPCXyPBMbWHpJTcTt7AL31iLAO1tOVv7ZM48gFylgABBDk
7j63SDERLxTJHxF1Sq2f7JRN2LEOS0utafEkt7YDke15M6YD4YwnLZ6Ly/JrjLRG
clhTK0W07HaqhdBKXe4N5ItMcZSJkO0nZ+82CEGNkVCwzo8EvVYutH1u1QR9cY/E
5cJksH5Um7OYereluNHbfaV2FfG7bDuc1yG/cVg+248cWLqMRsbSnEMCotLoxOTN
bDGO95kWUAoBv24r8KzewGJLNESdL+L4q86MNuwV1zlZaLX5qWMs9C13yNqruT3k
oX5L3TnhEDW4Z4hdIMb9LQeY5kL64yp/OQEK318NC1MVSUyZxviXhxOis+gqoaJo
CdxnZOXnIxL9oZ6e3xnB3bSMgstYmzVUdH1w/hNEvOJReQTwxZCgOd+CDDQsvgFG
/HT6pJvE8wIyFPv05qIS9VKlZCIU1JUhch6SFZqaI6Oqa/dRC5vbKueQJtJtvbmR
DtNsXAcYDkRfgwJVaR+wFpadq9mXBPfsr4M5ItG5HEqCOAncOJPMJePUBlsQ9Z8F
uxSfEX36L8KlY0t7/37+AN3nz1zNG9Xadcvlme5Z4rZO4YAtzFIju0m1cxX5Lzsy
Po4D8kDz6mNyE5LSk8C04OcHT6HGm1RJIEqYfohWBb58o/IAWUN87CQUQHHDjwQB
WR0jcn2V6KWpN2XyzwvPIHLzVm5C9XtpTe9K2ZBfczDCovWFmEXhQ8xc/piVHMTT
3nCR1XtJqrEtUrXHIoLCtTkuGulhwqX/pmEXBoxsE9VlNQ4WKmuzDByK0vV8OGwO
JIxpmAIqS+P+qi6kvm/F33qT26JzR8UBK1636E+tC8EHTdMSE1iJm3vgXAhqsTIZ
3CY92qVxoXFE0xkdmCsB7S8PhNiIINk2q5CafkKzzPapRXkvHh8NS6tqpQfXPpcC
uAgt+dfFaRcTxexwMWWpfujhNm9IyOwd0m3GQ6NK28i2v1BRx3q4k+5x6+V7eB4n
UGXaQUAqcAMrG/0Z56GhGzB0kaZc3u+roucozhBorHR7jkb2huU9gpPMnNmkQQr4
5m6gOvaCh5pgwA+i1tMo+32iLewzi7PMzKQeGisNVro75PXRayUmDirL6ghKEvyE
8rBcGrrpWGE2NQF0ilqy4rnrNxH8yYIONXHKjwZSd2QjmE2CfjcSYlnEFUwM6txj
+9LoxIvZjyD5kVi+uSqhfwewsehEppYAVQr6vGxs0bEr5M3Nz2jwacOFe9MWdtV7
JPELgov/u5p3OG9+wr8vLBOh8yFN6Yp1IDZz2Jt00XEF/1IiW7EviXP7fIIItx22
dWOcg6nAeKy6bApoU3b2VCmpZ+fSeINAc2gwLQcu1GfhbTK4Hyf+bD0sF4PpF6IN
NwD0IkcPoTRHrvaUe9baRvSdLZzw3KFsolhevgKOqlpgEU1sRZrl4gFrnQbmRJKp
hldGway6oy74Q7oHgCHuZU+g4ppQ1hPuB4fbgIoqBLQMjUqKF7Un+tyTtynrTqEv
nYCqUFqkck+WjYKLZGtLIfUf691n8EzwIsOA29ge2thJYXrJgUzpIvhORXPFoFf2
/4lQ7d8vS95933Orj76gqEeRdwKV+g+NO1DtQgOWOT7aEyhJK8+R7xZVYxJOUIHj
4I9L+TjQgOimcK5Qh+NpBT6/AYvrXVzCaNtXrvhXAdUZUrWrxle4ckgqw5VJQ0eO
tmTF4z6fnCxD+yDhCbTqoOyDjvDJvdEiIbI5OITXPSLeLHtMUVFybqkSVrhzjEhX
IQ7oluu7jJAEw6QoM+W8mHxmHT8ExVU9rtmPwRF1fKyPpVP/D+BDC/yCOogk1ywM
2tcYJXJkaQxM/rMHDd49NFf81EI+BSeoV5GMujYh/gzmWEkUrm35gl51+KUmj3/9
O2ZHwxWDeAEcmMPhsDcIWHODAl0v99I3lAQCYKkq31CxGkcDJr49sfQqTZms0Wwx
XJ8do/5tWRnEr14P9qCNy3ajHhJGiFJeysBEWUuFKXwvXCQobkVb1iomgK4TZKZz
yFtndf5zVCwX93wzXfA0LGgfnBoTf6honjyA6L6mnmbBUvgqwiZSSAOWobKAiUvq
U0AbU6aiIFpce1XbAXb+9wjaiJs12gW0/Rj0/g17hiK/BbntqZovnJbESzNDitcR
NvMAl9O1BczRWs/Gyc0ouT10HN0MTMIDZzgwubcyabHfvwXCjevft7oqpQ5D37bM
jdYV88zez8cqcEZmemaPrYsrl8e0PkPfkIgkG/C/TZdAGKRNM38tND9Ef+jjWn8h
m0JU+sOQW1HQV0Yx01nm5gir9Nm60QsBPR+mPXVypQqiTRkc1CAks4dSFysR89vx
XAZZ3dUNDD71H1Aqrz8JDGa2PvnTwsVv7QiDgD4YfD8LItexuTDoBPoxxNdIaAm2
aHs47tJxy8qydqSMtqV2+cXilePP97WEfi5YamLUltmDsvI9EfwsJd8V+kKMtib2
z1vuWSoc/DhOtV0CAECSZLhYZJQv4WvC+yZBXnE2Xd7ctdtIp+DRmXr4Dkb4BdQf
a1HhnSRQAO7osBQFDBRCmLc98ZeF5wJVKTm/iq17bj9dBJqiPKjb8740Y9whhSBn
4knq1QaNfvrHiU8AAbJoUJ+X2q7jlbNXDJWBczusWCOkc6NHUrAYtG09jwGFkE3O
3FgoyHa/y/kTpucnBTm7WRHGpp4WH7f9S8WYDJ0uFxZFa60kJJEIkxhZPdaI9OJZ
OSdAhPYlRaxprxXJxylqDTYm41HGzmAsrLZSFSvLuBjCRqMFda/wkZDwqkqguL4j
3uKd9yq7UXtX6YBVMuy7ycUlwIp94Awyt7+qXJ+kbTV0Wel8+TRO6sgPXjkwQ7XJ
3uUi7mzikueqwiCdxD59L8h7xT9qYw++bPTQ/MJX21lc1B1Qpjg4w1leQ/t+MkYI
Y4kxjdvJUpQutLF4Phkg4xpOYS3L7j/AlISwCTrkVdvdBTUM9tdkV3Q27WVL+NR+
fKPtiQF9mEOsKUs6AJwhOPfSTh9aKQBQoJh135rBIZEHlqbqCOzP+j4UL8HEONLW
7NxgOD1bN9OVT+pQndfldF9ElsSbyTvsjGff76BBvMc+MUew7s/uQp5aK4hmZom2
cZ2czN4RACHNCOJ5H9VxMDWWnX3nWsr3pkRyeKBwjslj+5wBEQ8UjL5IC7HjV5+V
lj1/Mh/Vo6stMRLrtKBl5DkJ/hgqoDRhc6X36hQmYaKiX0fdeHhpLExJCEvpbPi0
Fp0uH9I9GtiFP3gQN5gP5i/bZTDwvcJWjGgcXcilNCq+rydWZ5oTETjX2q+EoPo9
hrWW/qYt0qgA2wpiTTt1VEr7ED7i6KWihC3oqAtI99n7O9c5lftvyoBLkKu5gU13
F8lnA/G/znPQwwYNA3ZM2SbqbxGOsbangjGC325sXMh5XHIEOqEEDYGlYHb3BuJg
qjIE6woUznkjq5jtSyaHk0pvY7hxpgXKaN3SKG1B2A+XnNi+X7BffrjGR3hCtzCF
jniIqgshSJptcSmM57nw8iqIzbt7qMBzbayvaCVQdL0PeOA9L4OYQe5Z4MJqtVV1
hNvvavy0F/lcoJVoUGumowHCpQVtWuK9wSI4ai0/3xBPCfBROmRxYBNkiEI3VEKw
X/H8E1ZUgi7bc19H+ogNml9sGWegSiEyTCxQq+8i5SYuo4FDNp5TNuqM32XLtTKE
+2UK72KotHygXVoXsA7ueNcEyYdMr0EgzZ5m8Qz9Ecsqg6O5qUCH5cMvXiPVW5zA
B3mHsPQOWX1cw9xfa0PFfMJPh8AQ+yl11Vi/0mwAz119xQEeTECenfpx40aA90PI
ks5W5cowVqdbQKBoFmPJkif1n01ypvWuPPYJQGTiPLlBW73LUq+VXOkAKzMAPxch
ht9/QW5tPEAqtnye5YQprmeqwGaq8n7GlQZgu2HxYPnGMBW/XArdiSeQTZB6WWDj
3iNvXxSAOsPuYJIJpFBKYTpTvd8u/uF1l2DIqn5VmJFYK8iypUYM+zlldc9ggW6l
tHTwniwbgwPSoQO7Aal5ZJ7sxcOndSEcsVb4GVnLP4uSuBnrmyouEMvLbFJV/zFI
MshA+s350VOhXPk3udj8SatfD6M9VwS5C4ZhV62ou9P66FEEepnZQvSt4rEh9N65
eaOgX7ZofvxygiXh1SLw01GkE9qejKj+DMswCq4Nk0iJ522j88eonZlvcwZqOdNY
i8vESt4Fdv/iIfTH2o7+CSzvSRFNgvu7PgEj/fgV9LhghRQl9GMLxQg6Rf5n0lSy
eAr+fFrn0LYsns5+nR97tQWqmviphHP7thRrMbCsDzf92JZ7r6E3T1XjFCnftS7L
1Ic/rnEOJiAoEoHwDdGnFhuDmPgfnl1pLg4T8aAjO923yAd5zsq1nXbFmOGlK+MI
/zOJ8+C7WX9oCwWOW/mHEsRyYJrghrCyIhuvItCaYMTeT7BSTedGempshZIgAW00
BS5OXMKl9G3s0vfm+7vhk6vgJ+iKtWr36g3pOtHjwBJRBBCmCI6G6dqMu0i5dWwn
3ptt86hwEdFtHqJlG8qKhea6/hULpt7ZMG7Zb1gOY4+RoflfWC64wBfnsXOd5Hb0
ykONjFN3gWZWbXloGZ/o3tMFajdCFd3i8mLJkt7yWHYoayIHqkdfKL3+KcMjSrjZ
Dm3IoCqACK8ZtAYr4sXyPCd1CkBDkTI15YOJYYRI76OmQs5/uB5jjWTufS+3SzYG
NVcByOR2ewVvk2Q66rO/gVmEf7i5FwReoQhDrSStw6ZtjVHftq3TQ0I1PalwPhW/
yov40STrfa7E2PGVKtDj/nI0qp40vPaPKpS/hohjg33ZkYssh1CpvoPBAdbgvQJ/
t12UiSjEUuvfiqJthL4/bti61+YJMrGRDi5BIFUWSpibaU0hYA8A3oVanGY+CNMM
fhQi+gAvRgv79jq3ZGVKqsQo96RgjWn9hJqSmyG1kelYjZXAi5/r68AgybH0nfYR
AUwUMFjwRaShxcq17RVzh5fKU0Lth14uwGhqxfq99zinX18LBafi1uxLXKc+F1sr
YfG95krZAZZwbMaLrzRAI4uJ0t4rBIGITt+rlfjE1lejzKzFm8S0JwPT29oydd3K
cSqCnrhC6NOCT9QmvgSgRtl0n6JxuCObUKCoj+X1fQv9P++dIHklkrgn+lqYEaYI
AMcGDA1gxYfx5SEBNxUJ5tzCHwc4ERygBDhv9sZNeaXySYgCcsceqnGavx1w2cxL
7rRNAC62gAftbg15q+vRRL795l1De+IhSpFZ3c6alpb6KXr+DwiPtm6XsPkGjvcZ
05DwXOtMWdGte7tw4S4R2o0DrLkprwp9s4umm+LbwC8prgsX8rcaeriJXM6kTv36
53XIpHWeoxNJGDYHluExGu6/v4IUxcpmJZTr3Fpwbv7FLI9PhV3p/shDYx0+oOYs
b2F5RSAubp4sEpgvBAiitA43tLOEKFtZmJFaiuUE6BEsMbI7uu6eh2xH0y7qmHJW
upDUwLOZrdiACnAusM8A5V8CbUoMkYfgDuFPfQ7vJ4honf8M5ufPD3NWQXyJ/RP3
L+GVUT4DRSBXdPkRTZuDaStZYZiPucLedDhD20gCzG0Zqu26fRPy03rIthlerfAG
3f8aF0K3zcskriTqIFyMKAFabwd8etEozEsi+WwajYohBqQRMlKeVzBPxTkIJ0UJ
9JXQnBFSe7Rspj4pVoId5Did3W+SXx9DliPao19xC/nyiyStT/RUSz5UZ3XQjsxs
zW1qfwOizfSMhQi9G4IpX1Mh7fHYaI4+PZz98CSpxk0Cj0536+hUb4ehiZuxGYrL
vAeYE7t5Ef87ctNnALaWiVrrsEeYiclwZQZIiOFeV9qpY1CXQSfrXc6zOVkwV4EH
qgMIuJwHhfoF44PNI+lZuTnxQq4d6+dxbCrVurIE/hNmoOz/7CNtEouaXurqH9Ys
3OBhLl5wQ2k4PIkHXegJ06//oY5z7pXA2HeTGcJKlHfS3IjjD/Hx0odyXxntpu35
0+PZoVJU7a/qpyM4KX/FQGZviZjk7KthgsDQUdFt/Cd45yOVBoOWPFA3HyutukEE
OfoCXHT0b331gG1KooIdXqY+QghhxOtVNBCAVF70GMboaKyEYR9x9Sg1x930tWih
ik3Oi0lLtxT13+Mo9irpkEQ9azGKl+UdhKUTC8cGG8+qI0z1xrjtyabV8dStgIuD
dZR3A5II4ssmOJDtp+ZUC40teOASafORTLP4jFSxzLwBwQebAWZ/vgD+WpD2ON6V
mL3kATycg5G9DSHxMW/crPccHEX87/6dpKra0ywCB0M6p6m1d7Vd1YCdqSU9+E4K
cnAlZpq9eVQgaxwiOvrpLq4ckmV3l9+GYW+HJRbAJ3n9kDf4Zf6sL3pDYDRrx1Ur
Qzy8Q/EJXrHRsh3SL47RDLTLv7uLLG8XZ4GzQmsFjBOxm55GwR5woWSCbF7lQdX5
yYib/tgliKiicX+QrgX+Zxltd0qIfOFPnJx+XtjNCJZtbq4+oHZNNX64JT/DBfFu
EgPXzVzN+QIoy+GrY2/ZBpbOC0KrPJyiyyehJv3d3VEZF535SzeWTk0H77Zx9vKL
GNFi5fxoZQN43bfRjEJVvz/diMk1wjkvkQT6zb6PFDei1KFXdooqD+ChppkPKQdH
iP6FPQ8MGsWu7al9UVUrI9SqQlxpTcgVduEbWm+Xlj6kniyBf8PJ+yLUFL2hAqOC
ARzVnx8rQHEfd2/qATJWNOOcLwQTdikGX69ZTuXv/sVtog/ZIbgd5Q1Rr81W9CPn
25hJ67vsNA/2y2gUZAaQfhZ0LQ8uIuvmbvdrUy00G4P48acJRIpMRBStbPJrI6Wm
EWei4v6MfSj69fcKPRiFTh/lUQYyUaPyhdc11xPDPWfugS+OGnRXxwUiRrW1SPir
m+3jgXTTH5/9BOgVKvQ+cMI7MI2p3a7vfhOPJEDP2qMcNGj3rcNLwPBfKoge8sKO
4IMTO+R4CtSLAZg0C1p5jUElmmUpgC7BEyfO0ZLJC2dAF8RqjIYF4ViSXw+e7+Fk
Ji+5/awkVzAhdjw2UgoK6cOX4/kDaa0/QcTwluup+GoxS4AiEJAJipB71261K8W2
pjCpjEGMH+y2wNbnTL5gQ98Ucr4bBqtvVCgOgH6eFCrZzlNGMjwRaM+PveYbe6Of
GlTf9Q86IUNEJUu13Z5i5kkInCl9h34kyAwqyoJrfUe55pCBYV6QBXG9hrA1RJBd
TGLyb1eULG9wSK0UBeVS6DpaIF5s+eP+WRMurRqt1YUsNRkdO9NCoHfuoanDBikg
CHJGD41RFPDs3VJmmI/bm4CpAXMew5B9eELRX+D18GRhS5n81K36b8fVYdnbkH4Z
2UPe2z25MVyQv57WFaL/ZCNuS9OewfCSPvWGblmQMrvwbnKYji9X6oSZkEfcgL+c
votntbcZaKo3Ee8NyEIgrKg23cmvGLxStAu3B/RN75fWajb9W5JiKp7DfoSnBynB
o50nhPzngIGivWoSHfv6kp24N+nqZtCz9yS2utH0Tw14alNhHmnD5oXlrXaeDf1+
es73hpcm58h0VUvJPZf0CQCN086trtyJZA+48F1fpedeEUPpE8RHm2O4zmkdgiMA
AQGZnDSUlijbbx4G/dPWnf+C+3YyQNO8+8jWy/V6gIZOJtDkWzZ0wXfasXjKHOSQ
scE5iYRiUboEv2O70Xk20U7oH6+a60frVMjorU6oajc0c7apJfpejy5nAVVQeyMk
Dt7td8c7QhPv7C28ldQfe63hjLsGdGMWrygT/BUKdYlwpudFhXVCKstpm0Rbh9Xy
v2pUycUPme+GiQU6mut80wWNfdpgH2WXYum3NevXgwt3pS+Bi6MsXqtlclHnARPn
CD3E7FrCbdD9JgDzpkCvEsshLM3NkmcXX39wiyDYQUjfjEV6rQdXniAgOxNZ2Y9d
60fkWFfEFgNhz/hpfusktag4aPw/yXJplGJ8F1yX0BGruKzkvCPoEldEm/ct+K/8
Oq7W2zOEV4VEocPVtNt1XCMO5z9Emu2DHdhm7S0gABYxdB7WeuzgbnQp0pSskFHR
oJlqXQMnv71hV0CaW9X7O4e8akYJLtMjbCKonfCLXf2z+fnmcnna5N2VnawOvx4S
2mLc6rvw+B6du75NC7TjPkxsaZH1tnRhbwLJtwD2NtAMqj3y704JY4234KFt6ywB
qInr+LVGfHwylU+AmQMKOIOoTm10cQFQ7M4BDqyuPHn2OIxPkh2nJkh1QARTTOLT
3rIKUj4CfGp5y74803RhskXTF2qAZnqUzWPQTM+gCf7l3uQQjDnvOoEvxbrhwd1E
8Vbrwgvzo5GZxEKWTDyfk5RIkeF6JaDHNaFwRkcbV7bdxGoX2tbpz5q0km0tDvq2
k845FnRoDaG+BTaFhSbS731Li8UGcyDxdIxIKKgTam3d24bzqHYBeC2Q/fOAyeIU
3ZHBB4V0EbzF7c6Cr9qNbxpgtS0WMWNYLow1zHSbeHEcLaQG4u/xYdzBfhVPFnCm
PF8XMtVa6Vwo78gn0jpsnJUhmwmDdJkqIhF6TCSYrVdp521xRvquyruoLDUtMyk4
0qPp8HzryYHjrUJTdIN77ryiuOVaG1KVH7J4736x7y0qUAzeu44gUGEyXsJeTQEj
rhcJG6BOBSZPWB1/ePuW45+FuryL6CtpZP+uAPhx3gR3wQgady3JWAy/Oj2369Kf
482EfyhYMvzOayEw8LKyB71Dm+YGfx+pnKuEGr9It6kFBnW7NrjsZfLet//Zj5i/
b+S5KS+wn5SOed0+1A3v7fkm4sxhDFbcU7DyzayR6L2pJyHIVCsCG5AWZ3FF77kv
yavVEm+Oe+HCbgjBPJV0a+O3cX1yzDRowCNXrABStuOGTlL3FHs004Q51W2Xi/vs
qCHjV6t33MHEBsI6xzcqlNn8KQ2r/2FRhREAUAlkB39ljOm2rGvwp8knAcTQD3jc
a8bKcdpjGrLzQFdaG+BFomYXydugV1tzNqLpSCorK1jgdtW3W2yhCHcWf3bD5ocA
LEAnJiX63WDBzr+geTPlvBwT7k0grZYhYzcUp62bq/cFUKIIW2o7g9b/N614OSRU
/6fnWzFAPTTCq+dHzXJLitrhhZCY8p08X+87z8UjW3iztK4zM/oO46dGlhHdtjU9
pc3kfve99/pz6rJfH3NnMz2mfjxgTGuVegFGbC9i7hn60WKoNz3NMP+W6Nx/TC87
Ggky1qBbuKVR5uuMCdKwitCeHUVTtzqUCGsJOIaFVKDozWM27lD44JVRl3Vs2xO/
sZHD4n0y+4U1MeBnxrEzhEC39mHlaloPv3aTqaO2+s87yR0jypkIW9HerHlgc7JX
0qIdYUxG+G3QetJvZ/UFSafGPJJIux5FaRkdFjoXwRyzbqOJLTf9dnhy0/EI0V91
5y5QdFXE7fazUbI24C84d+5MWpYsmgC2ZsPZbI1FQiUl61pawg9OOqnHF/CJSbI/
j+roKSL/xQM6YRIwMa39Oyfn1iO5UOTLjQn1eEXlosMPirN8iQX/iFN+Fn+leZ0x
48SdOWhEsYJ5H7c3cAR4ORByffTG4r+lVtKznG5QJ5G2YWDV/SKlC0iHgDH80rN0
ffONjKGS6l/1dsYMqFDN2GP79pOeZ5UT7yR4FWNwze+O64aVfW6PvQ0GRU780X7+
6//UgjrhHjb8b6rCvaV13PGMYSCugp2UGMs9nhEqpThCRIIWvKBWdAJflX5IUQaq
mCuUdxJJCJBpPCj2OV9F3G0jirxuelhQ1lSiaRMnl5jDRmVVO8oPpcGB48TCZXyk
eQk4yf0dyh5GS6SU7+o2xYlzvuKehc6xcS48/cBgGaHmdX1SSGfnXuMyMUffce20
LSd4AcvBGlX1Lq2WN8dsBPZHei/OUiixi9Qb/YXQjXPEBKHbKlUjfzZDwOHno+Uh
D0/HcmeByPR5/LJ3W5AjbaRwFC38OL1lqbR49utCgAlUJ+++9ZprpdNbkccA4lyg
u6gPz72fG3eY51kaEd+GLNafvKHkodtJYEh8wC02axzUzbrSCh0+jfk16SRc60DF
JrHXeVeQiXQWZZCvAN9LMIEpON6QrWFFynOLk8WZ2zSjksAt5fD2LaX8R/M4DgmE
uSCwVr8MtqJgeYGByd0/s6tN0q2xmoMiqTMCoyoTcS9jFjZEXwBpSnQsTkvSnfEU
s1e/E2dbrd/YZUChA4XlzBdSURQuoeL3/LwFbsUHcwwGUp9Gbmw9jNykDht4eKO3
U6eLm+dZLOUqQu/HAo69QRnZO5KB0l/NGgj8uNaoeRK5c/xBTp88yMDySIE1vJzD
sf+c6UYnw3dBJkMpOo5bNMM6VoJCWjFyddUyAVOrRKJ1D9ByFPJ49A1e6N1VmFUD
u1ti6mR1id37T0ky2Di8VwyD/d82Rlq9rIQ67dc7be0RH4k0oV+EpI8GT3VOaBfP
UnBfQcT7riPaSsK5ZkuQjOP75iTsayTwiCsODB1ZP8WHHh5p0Zl/3ojj64qEFmKz
8xR0cWWHMjHgj6F+wsG2M8m6Wcf/HtT3FavqXegjr8zHn9PGniPzkhOBNp6HjmRj
m+rppJnhA3/VqBEW+gKtbPygAd+dtRKybM/QbSwXOmGUK6Uvk41NXv5iBmxPW8mA
/kn1gsadg++mXcr8cy/19BBtPM/s77zunVFSckJSLMXN2NQm1AlvF7D3EeCt4Hz6
Mc4EfU9msV0PkAYTDyRnwo+yRG0PwA7xTqoZkkn1M0Ik//KO3LR9YHnXmpcVWjv7
r50jmB4WbguvRbevTEjChXrXXUOVsBhrp3N5rr07VaQm+qMLqaSW4jfeuB+LJbvN
cpiHz6AMrmRG0ueJGlMNA/zWNqLLniTirTYfrFvLHLDBLwWErYeS8skgnzOv86lz
Q9lyj4tU520MI78dK+Ynllucndr0keV7WeLU/xl1A7MUs12W7CnYC/jWoeWB75rn
2A54nJRB94ZTXUZxKOeNDqyeLROW/7vkcaZ5EhkcePUC0AQ8l5kI4OgIhdPTRFwa
eYsNuohas2Y8axfbTp6W4Z6gmcZvfE0Jk90ZI4RoCZFXroCNPXo0cEmYF1vR8shM
deXVNpt/OWcwNiBKbWMBTDKt8D9ZMT8KnCkqUKqA5zurkR1/8A6Xs2vg+PE7+b72
yDzV94QDjYulA4+J7Xv4X4hYqnRF40UwLJME4XjPBgM/7LBKZK0h/fmyv5qq0WRX
8Q4fVzvKHr6AfIi3mVJLsrPOfmONY2WVBnoElm7ujW5U6P5a99xtenXTh36QbL//
LnW73a0DoIjjKwj3xg6SGLboyfOlhGK09U0tu/eug5yamLQ/m4CSXnYWA7M2+D9p
apCq/JnfLJ5YHz66F5pxQSg1MYT8AivB7ChEOQrd+8H84g8oQ3elBbO8GbjPWRGv
jpQPgbqpu+EUxDbRsMwh4sWfkwYtf+NupTadWfNj/pxNkLrmUz9RUndGyUzW8UHD
K01PA+u7Tx5mUwBpzMjLvQ2lZ7Dr7XWDla+2oiS+9XyYhfqWh8qOc6JwVOtFOeZ1
ZwOCiysKKSl2PFk4ErFnNIOi8vS17kFZ769Up3NWIBBSVYGs64oLn+0dkLioFwvn
bAmUg86Zy5TwUUSHd6a5f+Q2x6mXzGNJFMWUSoNIeU+9FtDQA4zTVEX4OMC89gDD
dfuGq9L2iDF8Jb3pHsj6yrbEDZ8eiZbPgGLZnWdz8KTGF3K03cKxgqFzpaOGYP8U
J2co6PgHUDJfjrDW3NHcMlnAle1TRUXGSP/wvEYjqpX/ELDp9cTGUlES1iFJBBT7
o5/zYAhta1bxkYcLR8uR2lj/h11XFMXFjTZB+8KiDD8I52GIlw0fzjyMZy9sZHlp
VK+zyCvLeyNUH5TjhU8D9JPBfe+u+t1vf9gE1+6KkUNZbk6B4MXa9gQ6L7pbcPpr
PYgtyjSqd0ChJz+SkC9O/VAwOy1WcJZS2XnNqE5HTM772CuU+LaOkw4dL19FsHmd
pUKGrxweOKRRBf06aNSHiJCNQ+GmGhv7Spq0i0WW4U5uzm9NhAYd3oidfJVvvSfZ
Akszt6D7Xb+RqhR68HWTLkPD83uNdO3yN9bdU8iAweIWq36a1PkToB+qTLUUHKFO
p++mj7lx6f56gRUKKBfS4fyNwabV6vxD0tEeg6ktCA8Tp4tt5tkYaJ4MveJXqvnV
PKrBJ/ZwSdNmnBWDfmuGMZ41xn6QkfKM0TJhkcTAfeA3FaLLMqhN0vCGoxaG80X/
tFEAuzFn0vAozMeE3xZ0k/bTMyH0A3g3swp/61R1yp7o4O5fpodzFH1BvQo7oPUK
s78LxJxrckFNbKMzqckheeGo82kvnhP542ijug/jHjcUVuaNXvgQSoteLgvfHnji
OpXRfE8wbaAFh4q+jUuvuF9NknCY7FRFMR5hIflq70Zhk2eIhywIWWaQ43DjXZWU
jCWJz8smBkNyvyKK4v217Fu09Sgcpt6O0XIYeaGnS2FgJGQLGTimk25H2CH925KE
SpEYz+A55pXnRffEEmWngXd4scWZaThpmNvqUS0LYEfDQKVc9Uaw5MiZd+RiVZ06
f1ydOFeFVl1VBAMuQsX0hZfRHHJ6oH67s5Jf/drI6cHwXFIamDFc4dJjBFx5AxNs
B1reUaJX7rp/YQmrkLSjYj/qbIE9RehBV7L91VwYkToT5DUM50YYuyTObqZr9nZf
VJ3EUh7euRxlG7i5VwOGB8iQ3yJ/nzJU4VBwDOCyB1EAxpcpfqBLdUEamY3OkOE/
l1ZLrPPvzfFADXigoj1pDpY4FP4Vo2xZCEGm+ifpZiAfvaZ9Cfq8MVv9/uS7/7VC
YiMFmf+gz+DsnCjqiUC9BGY/Y6YiVWnWNjCZjzGJ9jDE1TR7on1GZr4+rttDEUYK
to1AEMT9dx8V6qtOjoekeCKKzcbJImVrJMa36cCRr0UvjHucAQk0FDyAgwLJQm3Y
Prg0cR0nVkdV8SjdXbLMEx/e3bxIasuCJth4zzamD2mqe3r+fqI9AuC5VmlAmZgb
nAVqXpXFEKMPDOW5rxrftW+G4NWKVvbqqkBAliUq1rkkXM6q5DWYWpP9GWeeBh5B
n8AjGTQVumvYwL0GsyIZQ1KlwS1OSVydA8fnlPQG5EzM3kAkYnU5Ufo7pXdWG8Z5
nItLie+u/BOX5sOrVK4GnAE/rcZ7pSlTCLXZqEV599Fw0r+aSWyres5UAp66Li6+
ImZ/QMIQKCWqrH3YTFwHPvjAajU5NSgjhgVJgGAI1kI5d7SOCbWNdX6GdYpczAw4
EfSd2JMiUrUEKjkPhyeH48AoFX9XPhC+n+dVly+C970hdO3fKZ5GErjt3EtzMd07
3MkqjfI+1zMZbKuNFPZJE7WA6nyolJKnoSVEPSXFayXNc/SdppBDdUpp4nAK3cCf
R8ClEPcgbxv+nKRwltRvc+/wNcd2O7Vp7K8p6aVeZi6dMvW/kodWin/5XjkpbC/F
kvG6SYxeR289vbG/j1SCOEujCznBISYhRira/cYlBkhP2SucAeOKr2O5wHq2wXWN
pyQzjwnR3aRIJTjLlRSBcb0JCQ/bIieo7AIaP+BZ0pnu5w4Qp46C591Y2UYRara6
2FzGy40zjoba0YTwyLmZGVdq4r6mlPJSkmPAajoRoqyGp/8RMQ7LWSN53sv8wbUg
hZC2Pp4zGdF2c8i7uwwrvfzTcCX8fMXOmscozMWAiv3NITLXAm3ayB+jgQ8CR3Kv
rPcXBRmZJXQDk3nnK7r+b4uxYX/OJCjbWpuuqoNLfTTNCtB2SF1ccrG6/uuM+W0a
rTsZWt502WzVBeN26uWF5jBlIFgXUIHgbzgMBwTplCsV/aqm0p/ArAKLsmv1+Mcs
tBcuih6UZ9e8RLaBlEld7P8Ox5Qcqa+OBNF1IFyK/MBJjF7m4id0dl/ke5anhQlg
PzCkIEVsDluc4pAGvEc/LBBDPNlmGO+/Stzt1kUJNHYedO+v43FVQmLEiHQPsypX
u1d4j5EPI9KSgXOyGlkJsg2dAPQzLRSrj0XqczWsRHJofTl1/tQITRCXYG1aWx70
iGij49dQcnEZRSkclMEUK59AmBLALmljjarbI/8QEgx+8IofsI18zKaXzVqrRr7s
LLnYf/sPizc548O2qHrlMgWlf9OqRSMhKRaP8sNRLSE5tizvyS+sKjjq6v4MLHMg
4hpCff5wJyZ5DaJJJcMssMke13UwrZYljc4/YXFSzfIWCV3s/4Y2kCE0dA6tIOek
bO9tGDoCJazzaeXRHOVE5M55TEmN5mNWu+6BTIhuIwW9Syq3A34RUxxoTvnMVqqA
wP+TWy+SSwoMeMjBUwjXF6XJQbb6Rk4fA38dJ/liItLCj9zWfkQDQ8tNZGN1Xvuh
t/WWyUE/9bql+k42gMPk8UnSOiw8djt8z0ouqupKBsHTd4mN+JpAOEFZVzsYsvzh
KZi8bUwwg9yMTs5bAEAuHP9ZWHHDbMdiRAUeoLW4P91CEr/omZ/b6aR7YlTeQtpz
3PhgIixd/GiytQTHZhpj7iaJ9x383ZJAKZCTCVsmNcxX5KejYrFxkETqcxHF6Feq
P095JBRr+TcAg2Bii2hi1ua5myiYjNFIxc4r23qqOgCuPac4SH0gD+2BmqzNMHIT
LSrDJF+5wIka2+y61h1RHHUsjF4UFwO32dBo83LCRQq+8yg1qn3l0OpTSlvcTpDY
o5IIQTKY1Px5bVck3LVdmj4uKdGmgEdqd4LNuFjxoyD6GOnDwhcC+7WfvJ1NY+4J
ieLPVEAkCS1UW/MCv6siJNqBLF8fDiHsjEx7oqDlqvWlK/EpI18p63SgTOExlj44
ryyDGvRmgcpY/mEzGwGWGmOnkwSCFCxz6fK8Lva6D9KLO/cxFxPeX/We6BcD8fl0
Ir5kUbFyPA3m5uaB9XxMyFNNxKD9MqZDzlOuHPz1CX5LgNJ2dpONoSku/U2FYkcC
Pru1tT9FziKvFSDsizEO2Y9DsvOU2G+vENwlKCC6As8NUEAwXS5zfSOsLyC8Q8FA
/w6hizCNT9j+WxyHxJuRYMOd1Cfvvdczt23kKXbJDxoMsSo28YhLfBqM91cKswOV
IdwgnFxwMB1C4CW1img+Z+KZObn/rkcxHmmnGANKTAC0lx6ZCHMWfEEJDLSG5AcR
q773BZmaLFUxpu58AekR4PwXydibEtkML4rp6U78XGA0j9Im9B+T7gjLHx4bJzmo
JZa4RVkMAHVbK/HBzNbnbOotsdzaLDJxPV3Frw3vLuOhfRUAAWnQ0b978L1lk6Q0
TTldIXwSi53g/qoDsqPLobXnc3GZcsmGUpRxuJHR3MQ9w4j5/PhVojxy03nKRZJx
rgOVv1yPRgHYOG90ToC+G0d/ar4TL8Z4s3ERRqesJtMebdtade6CLlg+9+hK7lVB
3clRULARC4i//+WKYsCLojs7Ih9WrX2FV+DpncKRYOwGOYfVc5+IYqzu5xou6dIS
cq5FEa3NY6FLnzMSHwa4TsH7eDQgtmck2h6erum6xl++zhwaZImdiQnMFkjSFoYZ
CFwqU+5UG0vs9ZmOMbzi8Mll91Hpq8s2pOLHE8TAZhi07d0pIpzfTrQ2kF0ClGYE
0cZ4GZPEy0NYkVjMdxtosxC5+usC5oBVZPt+rJaTuNOMeHf6ENqQnLMaQRtF4a41
s8gpOYFSOtcMcelL78/01DHWVkUcTjt/QHXgkzBiEWuC7n+4eOFdT7Rf5swPB1kr
DVkWLvuf09+7tr9ZgTEJC/NDBeZdVd69yShncSIVjxZHU226Ot9msahqyfl4B1lD
U+54qYblDi2svAuGqeRAn7oq1jgdISj85qtBuC6b0NcVD1eKF2S389IaiLbtybl4
/Og/iDH83GeGE0MoiUx3GQmoATanjOXSvSWidT4tMzIKnJOWV9jPL9RKt6LHIabZ
FTxuG4Po0KnzaP4WAxnvLK8f0x7tElHhop23mjwMQ/PCE6a5TNash9LPgaYKraDf
BIn9TcE382xSnp0Sa8lsidOGQK63AZrMWomMlALNDEahn5LtCQpy6CbXzo7o7d/R
WyJwuL/qXCebDU/Qz7z1lzW9s8fIDi/Nz6yaC4ORyQEGIC9zKFkeRf8uAfgbHvSe
oyYG/rEcijoRFtYfykHELD5Yp/WsrOenoLelhwjHPmxyz+eXJmndNhPIrTI1HKGD
rcy5SzxBrSIvAfLYxIFy216eKXM/Y7JbsItIPKXEAIjzUAlsRuFNq/RuCe8vOYeW
K8t8erMH62WHLt0Jr5YmvQqVFItafchSpBYJD7ok5qKdObN4vMiQaafolnrlGDPI
+wDfSij0q6XDPQgkQ1nK+vhOndfcKwIPiR1Qf7Dh3MsOpgCcyuv94IN2cedlJpJk
ZBYUyHGXmgX5daAmeLL/uzPsYnkYF0LZLpYcXpquoOrZn5QvCgkXEFOeEZPdU867
7E8fnt1muoMWUKJ8Ls305iUJFE1UmuBYbDVIBJPTfMA8yaAT4zSs7snV77nW1WMd
yE2/w+rxUMw/6Fj7O/NtFwA8W+RMi1CK6k+ehB9tUuy8Iq6G3NmDSlxDnxGlHyGa
tgMPsimtfA4jTYWa+pxrYTpYNfUeIXUoVvZNgqDVdSo1mVfMFQhmljcGKLGlQ+9N
TDwBIPKp6NPuYSfueP8ItgFul7uEi4SrpuWKX2rYJGtlwtA0XTRBVGkreZg86MP5
vk2pazadk8BenhHY5//r0zyyF823uqc4Xr3QbWNx31vjFJY65VsrMpqdNtE9Aicp
0PJIj3m6RV8P6bdZj1Sy67eBwibG+Gzg+fpqWsMZFwMyT7VoJT8N5M+Zw6Ffszyi
m9GVN6Us4/CNV/0ZnoMZNjtfzjd7lE8QTvOD1tD/g4aDXG0UetLodAZUdLwB8okC
iMo9oJPnkmuPEMYLiS+xvqUUwmvRXWo3IYhG/ZcGCXeSCLQ2PsITvqVY7YWrt500
loLfxKyddmKndBVErRvBpQ4DesftOdNmOgqH+Qx9rBFiRdusxJi99ByMFSQB3Z62
4Zb/IsL+8zqrXTRatjsjaOeSddylflO0nRLWmjsvShB71t7qcRNIZ3RZb0dNi6lL
keA5jRa+vLQLyaZ5fQOch0kk35CIF4PFQfB7Ub8tRWOh0Ke7szRPkjrAsIx50V3e
HZRrisY7apMniHt3L3r0q+gXGk1XrCocbq2sbf6OtHdm+AZEtJK2iGhNzgRdF6Ar
mtSrDOk3gl7MLQdNpGpQXAOPXnj2agsgvxVTBHUdfvPDBSLU/qu/QvtL+BqnEo6F
Kr6QHaZV5VMOrfB/z/OnylFPrUl8L4pj9YA/thja+lBYKasbphucHvkWSGcFbBDA
r3AnC3mkmkukXvNLcAv+ct9KxppQVTQKQyuTf1PT+NJaDf0f8VgJoyyGhY/FymbG
+AfUpbnPb8b8NjmorW54chPrKnCT8AxtAW9qpGzAQk8c0ZeVT9J6CywmZJZtwsS8
HPfMtRUx2SUDvra2mzqL6CqUKPXgf80bVkoweG+SRuT0iUA8yWbcER7ztbozsguP
LXj36uSdLRGOedwvjapzswQTRWi+UNzQs0q1pL2tPKEPW80dJE02Fb+qmS7XIh+K
pvKslUepGolgJA1NbAUXhohPryY0ZSSrPR4kDIbmv5BRS5mDuY3zWsBcVUf/NvBU
/212pckXDRNYu1nFKgLJkwSpJ+R236AoMNIhd/eeq0iYBw9FtpN48AtTYhRjeFIa
XjkqpI36OGzRo1VAnUYRcBGVE4CvcAY0HB+tkoVaaHtl4yL8VAXvImjuShxlFIGE
F3JySwCD7jhzYppDfaa91IpAbzk0KojSJ/rClx3QTUe9N0F46QYf1R7MzbwhfInc
27pPJZvSjJnGYSPeYKzpJHdW5AsxqbuJ0N2inUuX4uTLbbeoTtJoNL8IHJuNJI/H
iRusthSBXWNdjp4JyUKECGpV5YlNYAFLNZTH8s0NlGFMOF1bOko/vwAx8RW5UPme
oZVWes/A8fKvz66FMv9br4YlWwschqQPp7N+QhpO1ZzlP2qFW/fPsaKSwaB39PJD
kZp6YHxNITMrOx3YzSPf8dCvH0BWuk0pFvqOsbGqeeYK3J6RmeBih4m33yv1ZENH
qH7VqnV6SLyKxZtAh/ydBTA4WS5Orp4F+vczALnfJ5Klzk1Ntp91XGJKNViBJiP0
Nch4FCr9BZAMZyEQzfhNU25gYA3oPd0l+OhNz2kj1Ahm6cwkFjdrgjyxgDqoFk9m
6JmIEI/b57hkqukBd2BxPC+InWq1/AMk7oi/sHf/ELYc9/44HjVe939oIzR5Kg0i
chw/tFBPYLErva/zwbOgz4R+hEp77eZ/32gsZ7p3VV6fRTm7ErbWmMj9WneaUb13
HOk8QCvC915y4wC+a/p/jfYI2Z5u/a+46e26fgu2lnU9Xk0vtJHCUnJaOfmkyudE
WMpsO8D4Z/bVlB1u3WD66dpOexQdx9JL9HdXJb64phphj4uc7X3odiNiKmktKhf9
ItsGSEkjk9jvMWL6FzQ2BYkCEMqJvrgCQvbmzZtY1TfdXbgu9487ounJ/3rtpKDp
bJzWzDJ9MRKCeyUfxnGXB1R9n6zs8yNeAvzxC9g6k3wJqWXM0Z0OPqN3Y1PadrzW
VuXS88m4t7nh1DRfOe6r7t+GGQqmPUSp/7fN1hAMnzso+Nk8mXAgxBVs1RCeTfiq
bhXTiJ/vWyGsmn/qPFUP+YKdnUNgb8DvlQURuTe3QFacNQgvtrhIOeye10dWfpr0
1ONnsAFldxvb7I2fNTzPR/EB1FeD2t5baMxc2tqlL0BmIXXVMB+Rl4ro6CZ7NIt1
X9d7GGrwitpCeKRDi0utO9PblE8nqrDnZR56jiggudI3SWdgehCQEvOJcIiBCzKn
6GXx7A9+2GmmO1kT3bBsab+BfBLJoVCP4sPEPPKU7nfjgxPcqpvM5Nu8zKoKuiwH
DJRmQud5q1z/kENNYLnXdzfNY1mSVzG7XZCySYerhpgYbt3XD4tTbvrMsz0zm48E
ZaxJ3+3fqf3cYcrXr4h7iNhaNWshUNmzCpVvXymAxx09O97LDNSaFHX2S3CVPODM
OVxtf1HXuzTrvM0tK6WBsqIznRZY5228atR5gFeobaVqJBFo6sh2tpN+tJHcAdcn
wvGutvLY1Rd+1GxQNnsH12geSXj2DWBLG6e7gaKnaItyUy/L+zw2VDq8KTyKJcJp
yZD5tXCu5WoyJkf+4nTDEVBQJGUrf+IvySPLj7sbFVX+nUEVB1bruElmAXf/ZqNy
VCxa+Q5xJ8x4E32mzZAXZZVoy7QucQZef95CQ05PAHDLgeWgtAILOTSKf1sEGGPK
wh3IoiWI1GqeQSW48RcGOVNfrdo5wbI5ZiJoHLKxdvCy7fS2VwktYK7OxhtV5/WZ
Y54e2ZW2yfFsGa0Pu0GG31ps0AdH3keKS8yhudxCba4bdkr7L0dvxW45NvdQINgq
F1WUWzn6H9vX4d94h0wpiM58rSEHAe75SDi/z1fMNePZywqY2goIW+WaC2jFjc9K
IqVz897DwBG27CxwWOzZoe+IEi3EeRNX1S+9UVkeIbEftaD7xtF6LvCU2dOHNQCu
YAM1TXz8YKtEdhNDOXRWD8QwGZREUlm0MF8birftYDixFHs4JlRK3RKcOHSFXM5i
bb/w+RTonBI2quEfxIfLYzHLDHGPTG+4WSQWmQ2g2g2Qtto88Uu7aRcvetAELTrN
6AuCoyEehn5YTxVAN9QtLfwWgcGReInPbz62jSpAFw8mytfaA9U+Syr3J3jWOfoU
LUVzhBzDdfo+a4dcoj+Q8tM8gZ4hJ4oIg0Mh/EDlil/xqJKTnSdj8Qw97xizb+yY
q903uN8uYD/rOeDTAs10tHDeuDfG7nKhkUrEvXm3A4nk/IOftXQzSNFqt2xPgINy
/78KnFkA3D3JhEHO9QmmEU34bNE2H21ZejMK53loVcyvVQZUk1/5BsasFmPByo/N
na3HfrurfRiZYyTJYNkLTCf+o8mpARxB4zUhHoel4NBgskKw3rXaoeOFqP1KjLUF
Wc3P6UftqSMHRY7iDa2LVIlnChO6XcUC0ztNwi6vXtull4yTOUasPM1B2cMK5Lp2
TeQU/G2a/MupIrbEtMpHdMsNgknGZIYgxlfbbE5mFfpCi+24FF7Hiyi6NZQ8rNRz
UBK+gL6AzHGX83S5k2G+Gt2Szxwgkh36eS5QvCpFoVfstQwquJ6ufKjDLONu2S/u
ueBn/e8iAuMx3N01Hhd9ePVW2ZljdKRD10ysWsKXyr5YG9XFXUz/QU2dorzV21W4
GVjNLTjWF9agaTV8k9YKpsmJXp61cIjo24kYKlP2awh2RTmNcit83THFXqgCANES
ydjfKkILVMfgpRp8q68AWHIhm3LMRF3bEsuZEJOh0zDoT/Ky89cSsEl6AcIrcNn7
xkJq6iFZgmerxZYWnGTNcSUr793MSix9RFFQOVFGo7nZlLZOzn1KaqKS5pvItnbt
lI4sDDw33VOCc9Ik7tohf0OQvIlouBya7ShVOUNyjYfa1F/LfCb2o2q27PJXk7hP
Ypk+n6lSsgO/XPYmlO0VkhT/wviiqOigTVpzsgrNKedoEkFmeJ6GwIOIVL5yeIRe
ruD99aa23WEog8vV4LqiF0L6DZPK+iuSZgxMsv93pemt9R0IsKCuVXjsNesYuSf4
pF5vH5FprYhQ18Yh8zO1hop6B7mACJ7vFod/VGgkbWnqFdTZ57YM+3jqmFvRVJb6
026dYXIxsDldUbouIpHMXMowpovtZxK4oD24ip/3MMMHySdjzZEX6KiJihJ7V9cE
VWwUtzBYTZjzBzcnr5yJBx0Mq+GZjwU3W/vfT/jlxfWESKBD2uwybZST8mF+7kxJ
4YNKsnxCGn++1voU2yqxz8/E4gLLNve42LXLHCEd6jCN1/kIYPpXYRN6B0M8yDbH
bATCXig2VvJOz4IH213Orhn/CdVYTLHuYciSnv0BbeYR8ykpNf+XjZ4n6ciYlmtT
0GAxpOkuQrez0c9L4UaYcICHZmqR3qw/SVdf6EuX4mFIftJI7Csoafped/RYiX0M
7vt2AeoaWayseQLWlXQFIvrx3+eKrftSBvdYKxlaW2vtXzX4UPOuEJwaVuEO2+ec
gefB6+AaivWOkW2K3tMzHDFOQMqzj/2mvabs/d+iTJredzXZxNJFWDTy62siIn/C
O4UVdvDTomDFwahuL0mo3kue19/KuRcNvNGABceEcPJZENuQIrgG7UebaVT2deQc
fp90lCa23sd1CsrMqCViH7icFYUVZkARyid7pKMC7hALnCfFa1ACCIfPUaQz3xSm
OtSYE1BKdPqKjR9pTZOMljmB7RJ/frknr/GGNTkC4qph8fiC0kyuKGKXvssAzvEb
Nb8EVjxyyTKNX7HSOYnIrdzilmwo5rE/WwjWt6oEt/On0YfvidaqMjqR/uJbh0Sv
SZytFSZN8+QpgEl8c9C/zFAJZBuNxPo+5VttAeATvJ3CFxYjk1nVJ4KOGMqcWhI5
fLpj4Q2z3OLcezUzmgVfMSghnuI9+P82i6V1f04ZodERaIpyEZsFA1dLZm8FREQp
5Q5KzjyWzIRG2QU/oXEs0UmCMFduXAzyIAkzwvnc9JXpA0uFP9PGDiVtoAXw6wWK
evHKfQIvoD2AkYSTVerHEA94VVupoxMrgHBU8xUCTF6z2sVNoIZw4i6lhI+Ylbtg
qu7JSVREpXnKAshq4MHwV8+4ank/m27s8ut1FhKbNEiu6LvG8BGx4CtFDK12Lk2I
8Byhn4PiXJ6ZjGP9xXOp2d2CPikvvZNt84HUk2vd/F0Mnqb2GyAjlva6iEbGgn7b
1xGMFWGRXqkrJkBmHVqv0Uuy8W5l69sf5ptgyXm4DXFctDIdTMT2NpmKDQ+Sg4qd
rDwjyoZmK/TI06l22a6afmWg6Uyd/bZiN0/verpbEh0i4GNPuK78pwO/B0InNcG9
llTfBWX62wB8IoUFBIEprHiWCRl/3fKLvkIB7QVOhdYgZGVdpS7Px6Qs5UD6Vonm
FllkX8xmNuiRARGXJF6pffm0Nux9sTyI6BBwBA4T3bvPPM4s8dYWFYGiP+USHppl
23DGZqER7lBUnvQJxBMb37ZSY/snMyAAGQWEJ4UYiK/kcdhoMHgoJqS28/c6Xh1n
RlaNcQeDa/0YSvvddEyEcJ5PKWoX5pszUlso4THs6kgbcw8zr1zEU0Qb8eiYl/rz
Vk2kJFX9LNuDGmxLoD9Jix1tI7f7o+KcXc+K8i/O8bLhNVEFiLqaGlJr+LPMu29y
ssoQz1/yoU8lLlS2gsRLQMg2hke/lymvpw6isU8kYmPzqwrGPfUzNcX3xS0sm01M
YQ3ndQhLU7klnrG/IN2x2iVSuvkhS7sg/Q6nWnRoIqYbms4psSUMW/DJGAdIrKTp
n0MSth7volBZDr1ASXY7jplgDDHGl6t88uW1D/iYVf+ecxFxowrHdYpBPrnUd/qY
nCh6euTb91soCZdOiuju3EYfLOitQIwTlm308UAw0+O8ywlCIqBKLXg85L4lKiR+
lzuVrSIZhzZHzy5jsFdlzD+DIxDVoCJXkb/+5eLoY6u8gRvf4yIIZAMfr5CwgTps
w/hNDi6zbKtxlgYG1kSN2Itkfke9FiOF3IYYHHnKW53e0jwA/wbeWGTwM8A7AP6O
IiQT6w159pqx4gN0KBJNDh7Xxi/cIjED0KCIiPCp6UnL/G2GASBEyf1zEUhKZ4ps
itt5wkjyEcPliy+JHk9MVV8Dn7rIRIHzye5cFaugqsm23NNsRCOFnxNjhQsd/SVA
IZYUT8KrqdJb72hTlOFX/vvdVPmfoCGVNAC68Y5PFAJV0urP5T847p5pRYDz2w4i
1kmu/FndAsfarDKQnqCFlif8bM5y24qa3lZ9F7VvxDvGWcNoV2NyctWyZVoJIOwB
SptJwXaxJFFeANI4ofirnIigWj8gK4wlH1aGxMZQDwJLu8JUzgVOqrQ++dp7nbpP
q0agNV5sQUP7nMkrtBRvowFg3wQnOAwrkR97AgmJcZwymQd7yqXPNkKqeC+lxfhu
FlDEJDx0mnzHVHS+Jts+MFuXp0Ywfj0S0dSwpv71RzbeH9nfHKmz3AhsAfcl38uu
6TjKe0OTsccfPvmBS8e+Y1ngNPc4nvmNBCFABUyfrxv6WBsy4JkVAs00wuS8EASC
RCY3jVYfrMpa5reGEUb9B+LoWEcWJChezrtVAPDh4xw2RWwy1SpZcH4ydai8omFj
K2uBPAPKpCWZS8Uu/Nh/LwXcDHMqQl3ZTpSOmrgUPrqckbt+5nZ491RFJDJxNhRu
geSF0ICNaXdIdfRGRhX/0/wgAi2ZbQcNZX/fyK6lKN1zuKbhYjQI9j4eaLMHnL48
qB3eVE3OGZRFli+w4exqDzGNdli1tUETuMViLbNG1/dukvifvCaUuOnM5MmY0C1N
N+q4utJSET6nAVVhap8oq3qJyq6+KTv4O8IQI433WghLcFlmyzbgsFi+3utOjAh1
9AxiEMgBNBR+mX2zAN711nz8HRN9/1usk59PKsKql9J+y0YjrH+cwpl1J7k68Vt/
CztR+qvlWmoes3TLMul+b/uXTp3QHHhmCwMXNSoglVNsDshkj1aaD2PWsmSkXygK
s0t3XdQfLt938D8w/xjP1bikglFan+cXNl7Jkj+orgLhBJW0F2M09BTd11vv1IhB
KJ7yJ7UOJCeGAicgZREIcP4Zr4N5PyJn78GzooKV4ZF3HsTfDA0IuzgiSjNvHEEp
m0xXUg3IwHNqGG9t174bdlk6OpxjkXFRKk6FZ5aRzPbjp0Ji97cuiacw89CnuRTF
Sdhw2z6NbkonWWIDRbAGvxg4SI5/en5sElRNjYr1cvJ1XER7KtBD5SfBStZMxbyb
Y0UuZJUB6TwEvAAKpL2IRWl9v41LISK+/TkcUJQVlVEAWjyxXC3trOenlyDkD7x/
oM/PnYlff8wngkUGM85lzl01J1vYmF4Z0vu3wm60/65mKTTXCezJ8105uCh8U+BR
1mZoBX5vO4HdD0c5CHdXLBztb2EfHnJV8Cc/KnYrszjqpKQTeD89yhldJKoGYRtV
mjNU1tYEbvUN7CcBJCguUU6qc8moOvMIaIK1J9H9h25QNoSvwqfAQhKAfMMR9T22
tTWGTZrae1LItVMHPKJ5+29/x/l5XHOn732JB7es++BDMM5vdRLwH9AofpvSgEy/
J617OEbSmQyY1fu4lFfN2WTtHu6DC1uonBYCi5ovUk0Oqn1cR7CLoIsb8ea7eXU8
6GrE5Lr/n2xdKdRAsGKwehH0rsdI+hujefUe6nhbRW6D/MPcAjOB7Pk8XxeUu090
Wj7y4V3qtHr3O+w0YmNTu8yQCADE+5TDBmurbC3pE0Pdd5YjOCMfvsKZJelo1nv4
XGgve+RiAHsdZL8lgq4N+VCVPEHkqZaPBEJT2hkR4e2/hGPTWFWvScQVqjoQ0Cap
KBB7pElyeLRCxK8kdDogG5b/CLNEtCOT03pYr8zI0s7f/dXcs3ccIbCAIjkMs9Or
/4qkGJAWr0rEx+p7FAGiUXeQTwJIFKcWnthwB6zm0yycRaLqkvE9kevSNTsx5V/2
bi+6ERlWFRe/0wza9iaAbxutASwfqaycv7iqPSaiv9nvXxum9i6u2IUtinhnxg8t
3KrLNW4fIrN9hXVxIxoz42AbMXoL+grwBASQZlf6Rb/GNjPFUJd6V574XAL8S/8+
zUGXCuvPH/qGyGbTANZxPy1q1T4ZiFr8egPMspq6W9F8eahktxRzCyHlhre8sV7B
UbywZb1CHGD4yiZnB60+cCPbKpiBd6SI70BJHiEBqtEcMoXmvVysrAbTZEvs2YPw
KygFE4opJsaL0OUT3eFnDOjufi85d18RLz370UUvgUG5lXJC0RjTjKsVnitqR95v
BvDbwhMIZ/Izvudf7oYYVUg/mWAXwjkIy/W+t4amFTek9wjI7oG1WjaKUZ+Dth93
v73ozSBMTxFiabr/5EKXu30BMsnUeIbrnzPI6W8qvH6PTe7XcdFEfKJlRbZ5za4M
kKFcvwVJNnjDXk5OCsEPCSQoQTCH3B10huS7rU9W1VnEopPLf0olXxOJT/Xjry/B
4ZaTbfeMt3DB+OIlnEOWkGqmIv5e7svcHwTfZfNW2kHxoWaWM8IR/RexIHlYdCuF
cmzr9qXaQlX351uxr8wQFZ9FFgU2lPGzI26MPme43/IkPuLNSngDHmjC2bE2yz8Q
s8Ap0tn+o25kmcxWtXb05EVLhqS7IwcZF3Yr4qEYoNBy8M012Rox/TB7tGqW6ZqG
eO1ExO+zu93LrgsHXx9psVoQdyF/PXRVZD/gJBM721fIPoaVo/KyJjrLjqid8chT
SINRGjbu6ptDViiqDIbIPQYAcM6L1gPGK/6atQO06kp/w9Rbv9+QyFqUpXewssqM
ehHw9cZa/Lg5R77W2w/pxf3U0Qr9F+crHC8FslXX5rHYOmpjv+K54b0NOHFobO0+
uPbKptG9SZuA6A8rAcY1XhMRsYG+gjK1tuew64whq532gWoFyNeEwTPev2PkORZ0
SRrNRGGJEuVU69HhjGQqDnt7lna6q1gSP+/ZW86F4zPgry2RLJ+QVFSEj4PW/+zg
RLC9aBUzv30odoCtszxhGNoX8JAp2MX043BsgwOWBIBDyoVbwIC7X3cZPRPkck9i
W7QCl8/6fwaWRpKW4Tj+TyO0uhx3jZa3gs8ykbN6klXR62UcsCZ8Ik5lb+8lZr+B
sGClrw+TZwxjWnJkacnf8K0yLuS/mrXwcW0q/0rauGHOTZEuUMK1xO0WI8f+fOUf
PYGwqSr5qBxk7aykwpUkCHyhgiYVYuYaNER+mTKkKcOVh8eaVupytYZJezA9riS4
htwAZelYL/xV+Pw2maDPDJdt0I9CbzeAgni9yaZlsloOb0fW+JBUXqptCDoKuw81
qIfCH0wKtuCbVQfJKkaUXnOuFneq4AoFyd2FLF6CFKn9jy6MH+P1yUtY/Q9lWgyf
8gQQH4k25+K+3k1wf/JkyrhT3vwXEjyUGtUWlNeJsydJ2BP0YA518f3CN+3a/q2D
jPyUihJBJlckjwcxsuUdaaZ5Je0sqwWBhrKEGZUoiifXjPUYsd3wuwtfCWvbHaBl
RxrpCzOEGtbjTBcX3LLMiEzWpzqNxLxzxLySV0QNAvLgGimnhpxpNtDpDsysBvjQ
9y7+xxZQbEnk7vg2peXDq+dzKLPVWTlEqbSiCK2A2Pi8ji3EBLMKDugiLtT5xa4D
YV+YuqgcFVCXv/NPmIyQ6iOSRXwBtbKTZ5cxGvbcemBORTYgQvl+HXCvYVsbsLLh
9nxPR3s75Ip8EE6mJDU+R74av9AlRrLLIrcWnBbVui823+Kdk7dquD1d3u0njtJD
g4UcDtA2zGrLcOhibB3SuTcBfjrWItr5RPRzZgwcxMpe8KG9Ifw8KefQrYU6g/oj
Nuok7HMCRlGx8YOYENqgvFkCLrecEnSYMw8lxsuj7g3IQu+DLkas2OHCsV+bjewE
kHcz3H9I1EXHVt0E65UIRvNv7BQlF2Gz6mC+KQzFjHg10L4Gs008f4faBD8lJNMl
Qkl+HrT6Aiyi46RanA41l+bT46R2hLx/REV5cClNkmAJQ8ziu3jbrrP3ovwMDvqM
1YSGCdzkz4fDHy0LSmyO72Q2YCIIei4iKXNrmwlG9htMWBh1UD4/utpHV4usMi6H
5Z2uxmZNx4OGKHP6hr6mzBoUPDho2UQe1Ir3RlLXo2WIHNDOb8xHihoq7nBK6v7a
ALmTs9Ogl+OTSo2WiAU8luWyzs0Fa3S9li4FD2KVt4t1djmknqP543/dQPWrK1sD
zJC0PyucPVLvXX3rj3WKrg1IS5gcdf0QhPpRZaUhWNGvSevD+5+AuqiQNpfDg5VW
oY1nDzK+J+zqIAfI2BhDQpYnLo+Pbwg0spW/GiaY2HtEFN2VuBFpq/S4jPMlX5jh
3hNBCi0W6eQXfukH5TfpnSDH8nnEBa9IWiHNlA0bZGY9Qc2NX+XPXHjP2EQsvq5x
6WmUsFg+iTaDakp4ImD51pU5uNJg3V2pQR3XcSXUIThv7waZ5tQc4dBKat4Xb6r6
+Ri6FH9hpH7daoCEdFVo152z6VHUuROi33RSw7l/bE2gUTI9x3z6IDjACw3F94fe
WBsuHmpevSpRANzOgdhbqHfGlVM1UU1dw9189+2k4V4ropBaAhBgIxT9U3LZdjz8
TBDMQcyjYHAn2469gEvDoTXOomKpE0nX9tKE7HmN1PW/0ZWGjEuexyU+SX5Kw+03
ozKA2mhHJz9nesrsCibe8pIDjSJb+v9+zdRZZe2lVPXvWjJoZYaZmcsLDHolbUa4
jXhx7vTr4nwc8Y5m30ow4Q5r0/OsSNL/lGLARjMYMOqCkVCct4f99ByOrf2XMUGa
qXTdpRcdM4/C2mA0ifFiyyFdWE/vtlVhLoIOI4Y5in/VRX75Mh2ZWh3uKc1CtOpz
Xfwp1n8tVCNye853d26gtskN803AY7Od+z00g221z3vDM/bxou1YUyf/3H4INNY7
1aNRBGoriDU6Ry9mzXOquCyGibATHk3n+ATzfV1YenOK7k2Z5loErr+HqLx/uWWu
OeykJA20d68T/Bmjyu4/EA06dKB51/fomNb59+uGVdxvExyvsSM+IYAmQ7BK8i6N
oGWl6sMRSRE+QE7haAeDCAnLQqZoGRITnCNp2Lr3ujtsCbgiUCQ6v+9dzBY14cRJ
XySYCeEEM/9WRGxMiumU57WkXjTA2d5YXbDeQDqFxcQP4NLxn5VATVeH3/LTHPYd
jOVjXYG4XYOVpP5s6qVUzC8Ayv/aPEP9Ku8AFJED+6xK7KylQS67QO+F3IJ+ziWt
BFEI88CCX14nmRpy01jeUvFd8brsafzT+K8A+mUzl5PikB72Q3IEkPOvaXimIVYq
DIVo1NZlDDTgjfQwivGXHm+LXSVaUBJ663GVwyeZqCAyAvN86mq9HpomJ46oMWZS
xt3mo70xieLyNXi03wEHju3b/1yu3OuNpyEZfmKouPXyd0OM0aDbSogPtoqoSpRK
5rwJnD65a6STcthMLPnQVYLVQb63412uRYqYb59iusD0lQdseyl2gYjrhy8/FfgV
D9LxLnz6G5iTR1I0yGuIUubtw/kW3p15WorAe5RqaNL+0uyXR9m24CkKJKmSipIa
nO0kmwqK+EqdKYlpHKC704Rwqe6ynP2rJtX1AFqc5ptyesbxj8GxI77MB1Y9ITtG
eWOezQo/amOVgPZXWPJKfNEvGg+rVSgCGvdrNScIMAk7tj9ouyBxINOF/WiCa+VF
ses2ZtPfU9svKh7mRfhnV9rADVwblI4rmzrmpzm/NstTfxdimXthXFfQ0q6qDFcF
rppW9CzkO7Wq2Rbj/K690Xvbvmg1gcUeUD5eK+AFzB4cb92INyBkKiVFqy2a61w+
fHLYdSQrtfM/fNt4qz9aixRSOy4lF8dzOq2ZvYDk8X+iAiVW1LG/W8uVOI/ovsAS
32A0suB5SrkkICIfxAdkx1i8TGk5HAv2IjseYRlHgA3YWE26ys8i88HwU/25zirA
0sqiM7FEOr+iTtgdEVfEdoRSRbx6GJQzT0iClISIRHnTv9kj7WTKTREMrx/MKlhX
A8hOSQfMl9uZkMPh6K0xJoWiNjBaueixINL1HevKteIdKvzZbXsekl+YbaIURkB3
Vfo8k0f3AtCNADj15gaqpzs3k7uGRGsu0IGysJvPA0Vk7WudiKaRyy4GqNP1+2Bg
1529aJ87hbDXmwDJa5yGNeNaJV+3GDO4CNt45M7hvyktzlrsWetjCFR7WwqV230x
NA5I5XzebFv/0xA326Lm3p3vsyDGvYMWWfvkj+tlYi7O++4+uTEJpyaYgLyEDCwA
MTXx+BFtiYECzdic25DzQH4wjpDlz4wma8gIgQnx1JsshHkYsi7Tkfw0Tiv4/G3q
0bIphUPw5iP0yPOfPLLf7HIIOtBCHnmgtZgYmo79nETK56fAWIOcQLg0fqQbZvHs
4z0O2gAjj9Rk1nDdQqWpOHsrwZZJhu+V313rqfF8bjbeyk/N78R9ihjdwCgkEBKY
QpIz1z9QTVg3WUO+BPgglKElNLrMO7+F8OHSFrahLwylGGMD9jeouG3SrCE6WwE+
EydcrDtExpVhu9LPKXjd7KiJwF9iyFqxhiETGEAOd7qbRoSV16J8BZeU1P/vH3nV
xXKo3nbu5vENlpatEMLbbyiTd/+PoLhmLbJES4LUxmfMqevzPwrHI1jWHo7h71Lb
qHF7xDYAYzBYl7kd1fGML3dx/phLHr/LFygkoYsI79Ra3f8ZraGnX7i+IlhiMKH+
V89hk5PCyxZ9ppimrIpL/HWe5fXywvg3V/0nee0UfWife1QZVCLZKeChnhPrJ6AU
ntejNO48wG/y+2j1qkBfKtjJWaWZHi4sqveSdTxFH0NIeTl2y/8EpNaeZJgGonG0
r9QibZCPYWSZ/vxDLyRgHfH+JkRsU+2xhmclceLE/982q6zCYCeiV505A6tqGwa5
da3cddoqmqufp2jxS/b22kUTc6s0i34q0Oa4CLlvBCc4F/14DNEc0JRmtKDhTM42
aHFAH0zXAINxwzASNXuaKKEiCd0FH1Asct3MHE6e3cXIs7XPBPywIIHOlzv1RULA
TFf7dqtbp4UW6KBfZE0uVsXjZnh4psrXWaERIGBIokoA0C+V/S4vBbZ6mnlLuu4V
f2ndW6A7k0vBw/KXD7CimgLRX2kL0zI3+Q7KmZj7GBYUNBEwDoJAIgp+4xysmUbI
Pj7y2uC0kIa1burO5oj8lKnxPad7IRIRYJ5OTpx0LlQtZdwkFjHNt1b59AeRcuOy
I7rzAOo/a0dbFh8MnHmp/l5zyUjc/GV46W9rj3+l/IvOILJj3tFmmG0YVf6K+8il
JPdmF+8At8sA73wojEJcerXeyGwUDViHYNxN6etFYdbc8aEXdGjbSJEXbvgcYleY
6QsC8DXQl9E7zyX/J/nlFSz94O77fnFP4uQabf8QByMsLq8v4MwW2l3B98YYiU3n
haDIf3fjKbibKCo3a71I+eE8LqeBx93ECbn07tnyuAHXTATa0TwSRq3LtWLO/E09
nkuyeJSiMAfTqP0dI4AD1GTO1aWwjHUxBssoe4J2PJCwJaHl47Y0AuUZukOfjUre
8u1T6sD/kMrS+a+cP/3tdZtsxEhbxrM43tXSE51yt8Y3vQla1OXpAOsjp91sRIkx
/cdlqaovJ+Eh14dFGYJaJmWn4Fc79saweyG/hGYbRd/YDcRjJNaG+u7qxYxF+dtw
VN+A5dtXe/RmYbCAL7etyngJxO3cnBKyWaUIqu20H0kLR7yMc4lYP6/cug6ajfE8
/zKrv7RWMDxYlTEnWQwpMJI/f8x3/lK32Rf2c8IQRGe0TCjAFAJ2yx5EHWkp5nbC
Tz7+9WK1xX3NfffDJi8pxZ857n/mqNqsstaqwJ+Yv86kxA8aQr0CjKjk+TcDAt0y
+BMH1oGc2r26xxdh12nBuuhGJ25X+A2GLpxNaw2qLsKAY4EbvuO+6Sk8/maIn9ea
xFp3cZIjGv3DRtZaq+Ve6IuafFkfII0iE32zjN9PK41XkFb0proeUCcBNFC3HvJm
ypjBsLKlpPrGNgoSspV2ApFZy8JEzwm/WN9F3TZdLQoDTs3znekhalbqNPCozwJj
/0GCvt5tV2ZQu9ZB06USXQKsfI17vKpUyr0jsqoPj14koEls6KlPOIYeN0vqaZKh
6qQb4ykb4iwEXSL3oFhLkEwJMyDCUIkXFfrw41XCgImTZRX7Cc6t6cpBIuUnsB83
lMRJuMy1X0DfulkeK2iZySAx0VjqysQrz8iHfE8hqtUGDYBXlVO6fO0b5wl0rz7B
fGlyfeb7Pzeeg3R2fSqbLIg2meC/hijuJfX7UEylgV7GgWZPWXWUmwcGihJSlhMV
h9/ld5zn1k9NeWjCzJGnxbTnlaOSzbgIXT9+przblKlTYr5aPI6QPfVx45h2yyNR
i49CFnw9Jj3tde/PzN7RQ3qgV8lJjoWSzr7fUj40G4zu00BJDJL8w/geaNgax/Mt
ltfzmCvRqowr6/cdnl24RZUb1wU1YqEl+k2h+VAxj83nW2qbRQMcNzEZ1+avGlUf
90BIlL0jjR+ZuxevjubVy1rVBtNhEPzOAUmtI73ypxiuB688TtQmlnEldwVM5CgY
NbMxKUdTDvW2jnB1TBDwGadPy/VZHdPd5PohiksRu9WhRlIrvFWwL7RyJlfED4GO
wfNZDSicEcbcvJyifFU35pmulLkSymlInApfKn1zG6I5B0K7PE3MKt5CyatBNmGC
w3w4tK5obA/7yQidj3xV2svaPZ9dkUIB6AK0Wc4olGuZKRF4bi4swoO5X72SUkBT
2LNrplXxqvD3HhnsWmLp6OGdAZ6qG508YDBmxPKRAXJhPPQrLOO20SUQxBx3rTzR
JCrzNEQZWxH2O5e3M+QXxrWLp82VMZGhn05BQFyRG/DoC9qw/K2ypV1c2Cpv3ROQ
AyqWacTxw0+IV4W0U7uIU8VEqZdNbPt04rWI0VO6e0CAB17r/gVW7xuld/vo4057
xLmBszN9TNwVRzTAAM68spncfduQEbqT12eWr9zvO5z+4vrxYNo0AgBk8YMQz9sP
H/IDmWgZKOrmS65AjRr625/dk77nYokMHWqdzKYRvgWgLCmOEDpxGtF2lv1lLJmj
R2i686viyxLaMrK90g7UfqbtuOqRuf9I05Ap5FdL1q/gFvh0dCUDYUpa8LeqWxBf
aSwBS9J5lEoS6GYzjM8BK0B15FujeWfKM6IGeQD1VjYNZOMvrUmVsQaJfazGhC36
KgGk3YLXH1Bx70XJhcCpX6y4ienK5oS7hvSNYV2U1Os6Vr2ZDQjr3UKWrT05HW2H
dFK3ym9Tm23MlY4TJCBVvSJBDuD8L5lO7VzyJlEQE/rN03tPTnQ9kLY8D/W9YIsd
VXZeHBYqVNpsrn1oB67H+/FIyvQ6HhjKo7ySejvF+9eB2laXzZHYs1cI3KlkJ1Zx
w1w1bFBMGs/83Wr0kf1cD3Pa4Z7FvXxhJiMvO8xrQGjHN8R5ieZJl316eJFZwiY/
mmRd/QZXGsqAa3nQPc0iH3CpG5KgaKVLp5p1iWugbdQDtg35vbLbM9AHrGYBQixr
t8nrMWRTudxMsKlTTc/Bjr4rv6iI07GMaXIAOpI5VS1a69aLfX2dyvTHBEMDzA7u
2UiFbsmBMxuaVawPOuNF7/D9IINNuWJQ0T1iDtDB66S45CNdeRzAyM79YJBVDYY3
Yp4TBSkMg5G34xc6NO/zE3N/s2YkzybAcYoClUx+sHUyDvxFt+3MVDMO+cj1FS1z
81veCaeZNXcjH6wYwazS45QDn9Nxfc609EG1xlo7MwJWYaLz3o6e6h+gRtFBM7xm
oLhMGYmjusEvPsKbdmwCLTaPuspSNakZy4FWGC5vhUwgHh/dOWxbqYb52ZHzZjlA
JnFQJObJ8FkVyfEKD9LJKLpdzUZAL0D4n2puKLmXLeKM8PTojriKO6X8SETEHGao
AHKzJo2PhCILQtYRHaPmcMQZS2D4qXDTc53g7KqNRt33Y3Xg2SRXcQ+2erG2x1tq
6caivfAln7Nq/Ng+5P74k4vdMVv2zsROZGVsoKnzThPidOJSJhSbKXFkUIIdovEf
ZEt9tf7pmQl7HbV7ooeAtmXvFgxAycRBH6CyUUzigyPd8VgbMAAko8+0TAkCBoT0
2QA2RfSpRTawmg41yijUT0S54XLtDJcj6AWzaBWuqbxeRGd+SoZ3c8viaR14y71K
SFbLobHbvVXmVt9ILVegJsyp18AKREFJROGbF+W5DzlQRdGl/bML6ZhKetM6KeWh
fMugFyCUviQPz+jdEhvlKVV8DhKq9uTXf+axcYng7rCxEuyOh7j+BQ8qb7mp3dda
NV3LnqeNgegrEqyTHy8Cf8gMSVFncj4y8NYT2idU2mllR8evZpFWf0S3XPF7xzr8
Gsc62NBpaJc5t7cbzBO2Z3TyLyLY95OWkF/D8BtRbB+l2u39OJAYIK8AyFIl6fy9
5E1oWTR6IIYfz3E3jU0YRYDvNjufywrfJn8q5CBeiMGIuWL5ibZh+zj8i9QI+/YX
ugT1cuadyOtWKriRHj5oR6TEldE/Wkzc2yKi/PcXamkT0h91wtrSQU6AQaneRnoV
aLyhPFAM/1By99MXmK2SNxx3RD8YLnQAjfCERok3V5E03inkANOElRZSSoATR0ZP
Y3ZOUxAltxOs9gVnPuSsaEmivvXAfPrULotW9n9BtwHVaMp6m1n6bOfzklErrYJh
i3vLpehibd0On1gxv7KbA5PQrFlQgfN/qCKN36i8/YVkMsd7DEz5si/7UqBwHiDm
b+7BXz3J7LoungUvCnQl83Q4dwTjDmR90QWOeo9IYuLL8TuwvCvqe0AEqzWxU7bv
Kqb9Di2Fm8yQIIPKp2igw9hLh2PO/fF9HILgOV/k67V3Nw7w1tgFXMcubAa2yIvU
UgGnCGNJy/cx1I1jLDKse1eycg5M5afPnnLT/Mb5Q5OHWie9jSDBuvCGLGutreGe
rtWy0Slm+IMLhJGQTiPmfIZgUHb6ltfSOzYZOtY2rzagCt0c3W+SYHRAr/FGQcDf
StwnXLVgQXhddysKyMKOpZzglL/8TtCBbcEZhMdLudepylNN1MEyhuhy9bHfFTpn
ibD+LlNzSHCxbNekVdGFrBlTPvVcV+6jDUKCNSpTbohBxxSuNaX4W+RxJPc04RRL
zxQwX2O77SguoekqA+Eyl+EMv/Gdiq8A5OC8rSR+VTbb3SVZaWBv7P9xHTzYb5J+
VnbQ6s0PKyxp5uQxBuW9N9fKHTMLlIThpo3wEt1GfzvxzFJRFCl/+UtU2UWI2If1
YtF+kXb+TVAadv+LlDRM/NbkLP/Kj+2j2odQPAUMghm9JUR+9cDkYIZk8SlSQc/w
RtTApBTGjLFQJPIKSh5P+wFVJIbyA1F5Ckzx7skRlcH21UE2gI5uqGkYSc4y0PTe
w4zh+VpPt5CELZZKTnH/KXNKdbPD7ZH8L4N9UBKhGQA53yCqp0uSqFMBSbwBX1sa
RhT/S1AbqMu9YtrYB3EaRo9oXAzxtI3FPyUfYO1k7RFHXEYQQTkhTkE+avhgmWKi
yKFl8Wj7fsYo+Up/kl+2W4fm/h+eEQSYTJLd4CWTn3uRcT0+n/5J+KvdpuxTu9lE
L2EN+QUvf18qITTEZukf8lJE/hg/Rtrsggyq21piQFhtXd57qne1Uy8Dl7IVZm5h
52kqLvYkmoS6I6GKL0qtQw/y1TbLB9ujBs+r2n62nS0T8ifVXyEbofq8p7KxQsUw
1/Gd2FJxAqpxi87fBesk4wYErpAO6RyXxo++1+6mPexCQLZCfinwcIiTYZ4kf2je
dVdKiOYzgQxs1DpSCQ+HMMfapU++BTObRIis8jp2FNVO77ndyAQXbQzn4ZEUYhd1
Tk81n60TOtkEypM8nwR3Kvd5mtFQ8s5C8ALxJ25JTPsEzUCbbOAcmIBjKLTAHcT/
HvT2J26RBLc0FmycLFl4U/iTg3If+dMD3p9hqjH6uLIJxrvo4RdGT8lleEPSdB+f
NIt/sjb10rpScMj+J28qPpYOIldDSGacG/81DTdFbRmPMWHT/bj0YqriltiURJck
/91fvdivgM1aY/JFBFwodOa6MYvJKM2HHRNkHecOShM6z13nOA4XZ/QGNP7Z+YwR
CJjIxjCpUKlGojsGSMgtCde4ipznDUnggWlbZTeG+gbYJfoxAZNnhmo2GLOxvQQ4
azBN0y4q1ZzmQ4+C9C3uRk42nzEciiOW7g3d+lG/u5z1yWu+Da9VDxQAMFY81mxg
2DnuoCWWNf2NZVnDb9Y1/+2bqll0VpZiPl9JMxLafpxYe6WnoX4X7amsWDqUkRnk
eKEBDgoKiDfbk5NETckYnuewNMmLbDfDuHebRmDamiLq5JJbWY8aFpgHo76wUZXY
kGX3u+vzCAGaU323xD2nOqkOEjoE/BIHsbLwVxz0ylEtbv+TcCNy3UwM+3JsNd8i
mz8yeCsPI6m45ndbG1+6Bq75w/I+1E1/4w+ntlUV3JIwr+YKziP9451sjUL0LnqO
v+NWv+PwGC1OQd+57HrMNAN0zJBMmN3m3z4+IEp68LfTNMjN3f5Zt818DVogtDRf
IuLPRqwzK7xJatYD51VGvoH4m/wUrho6pORrC+/cVMFWj/oOz9CR4iMDXlrv3XWg
6NhtH7QJ/Zy5yxzbKKvvYqLj9pwjD2lXzFqlvEHkaf6SF9j9HzIi/NzBvOF3jCuR
PzTsiOfMsRAFzVJMWGuzsU+lA0xI/XhbFX5twSQ0rqMZltY9VzxSqDHJVjHS6JZp
rYfcC84YtXsJ7CxPVFAs1ZwQ6Ngt9Vi3LLool4ERT58xRbkAZ+W39ucj2wso3a30
2V6ynJozKUX69BQFaXJzJDNtEBzgTneKgkw5LNGjPrpy7rQGxi4EevWagF408mzA
OkZ3tG/ATaDaFFjOCiTDrM4MSew22wzBi/8jFtVejMGhFc8612COkTn0LJ2w4FCW
pJF7bNN5VE0HFy21w4O3m8CVL0rI/kc9rokly5xFkLc8JvOFNP7+uFgqWuJiuSSv
oXevkeTCr9Z5BBg/Md7IGrq8j0EOqiLWUluncZnwwbe3QJM2z22waAH16yaBvKeI
MFsxURqf6whldYD6HIxbC1barBfQeLnHOqSPTqbXg48zQEmApeGXW41QmC8NwKlj
YK22jOmE+Pe3T5h8TW7BB7f9RtGAWy/lx9T9nHy08wHFS+tD8puwEQ1w55zEJyuA
yByNq1dsQHtpS7y2iwPdT35o8HCImFln+SjGer/OLPFeCp+1Ky3MfkuMmAT/wT01
Rb3j45b1TU/TrbTJiWUhU/Umi0V0gTsp6H3ohVa3/2rklLWRe8fIamfd/CreODNG
wGD9ftBBmTRdexUfhUjxXsj6h/XmP5ri7kuZK6GKF2B8760xxbfxKyABmZFSytAX
Z6Sq/JvJHHrUEVz9YHK8QLG0aZk70GmWRObLMAp1gZ+FWm3frOstFdW0N5V2gGlA
N5QtnJSnwOI6em7DbsC4HVsyguxOiUZu3g/b1YeykFJwDk7YGOp6BBfi4j2NJiPI
Y5dJP+86TXwsiUfATG+sSrw4R33Z6FANeCJw2lqvUhNxwKKkzLC8IqKNanjY2IM5
pt3wGpV/wlukHeVlYPHMkJrQIgloMXM2OT2TLx7Jb1MPntvL/Nt/x6o4A/JweLK/
0AiMEKxbdBPbtuXeLUJzjpCScecb6N9zHLXF7mkHuM87kS1eXucRnIy5vi9sBoc0
Oo2atWnFjxihMXlfAEebI+BhJbsHLw9B0Su6Dj17aPsSepTkdif3NS6guOXmDUMS
z+B8Ir1nSjKu+7QPAsWhsZmHJy4qI4ePH+Qyw/HFPdm6z/+ayx3oZpoYNweb4JRx
/Tbb4Muac+IDVlB3k8vkutD/BPSkWXxjeD2wZ4fGRXV2HLISsGxnrctguAer6QCe
HGDW2doLvPKJH1joYBl9AUD2ULQYK+Ho4HMRDwif4/uf+7eaZ5AJiRLtudowdQ2Z
c5/1DHw6I2q+GczkMpMaZhlJjKstqK9+FqoMQa8AP3+89UGUi9+aS3FH+qaBMgHi
4IgVHjCh4Vq++qtONZbplEjmwb3XSUP/T17Hky11LTa2qZOSenAJl6NaaSmS3q5X
SXQ9S/0UQi12L0P3juN0sPMuPV/Uz4rQxdJ45kP4ATw5ZXsI8Vm8Wg4xRnKdYbLL
1GK4MxxrFIrXsJMjl9qE1b305QkAel68xi5Z0XuFQLBBGNOCUKQ2AYNM6Q4OHyZ4
d1/prnpz8TaD3j2UvhDlVK3vvsN8IwWM4XoPER9VFW4yUZ5rpoMWzlsnB5thoFoh
gUjAvKy3LUJuKTyA2gH6s8kuHEeC1cNGcxPzfMCYjXaEaueqkA4BbYV08c2MCig1
GDH5SYbyeOaXjWCYpCIoeQH7Pvopc+6bBw4+xG6TsOGnUrg/Ht+g7+o2DRjr6E82
OTrkXX9oh7sa5ODu6+8/B0SFf0eODLjriNk3iP8YThNMILfwHxVbBnBB9gLf8Jh0
eRTl/1OWyQhWhl26Vm8hkFw8j31U/moIHG8Q1DWLE6oclwyytxMUodtzacPjTiEM
TUVUuVhlvuJaDVcZbmsyr9Ng6ubiiEjw/2/l+fUgG/ff1yl2z6917uyDgaDqshvl
1rQv9fN02Xbffjf/3zxRp3f3l+acRAh7c2DDSzGLDnRNP7910zcRpU6qsoPUPb3t
9WqoS6WMRq9oymRnykZn7Sbg6kj0Kvmx1H/spvJr97+h+pKFsxK0606CPLM6j6MG
tFLAQ4kTtBApUe6644TosVZRdH9BuXFsF6jLTrW+0MtujVxuifUI7Lo3dFz2+rcO
uulcRfLks9nWw3XgZlvYLooPdMmKAgTLcdtpjkWVUGR7O81Pilegnpu8t1o+GQRd
trXWap05DIvWegnL24RhGB7tj0KACkpKP4+fnK3ARFBfC9ysvJGdRlG8EZkRao+l
dQJZ36ieF1wM0ga9AjWTTVpb3u3jJlZQ7QK6HiLPUI8NP3MVBKASmwKbnyEITRgx
5W5JWd933JiC/ArWiNrgeSKe6x0VVp4V6OfyRuOn2dlIBxoUD7r2JAySwBpkHWQr
Daud3lAbZotOqBDJC6feXAezHKggPd36KLOfVbSq9euMQrZfufBekUhII1kVzEsu
iqv5Wog6czQkn+F3R7gP9sMMNA2EhneB6cDyQL6c2BvQJBUOlztbAxZvKLOjoug0
Ii0z67HniW06HV9m77LJcf7pbnx78bR2KK+tNWlROYTq+lRPA4zlCoKYWy8h2Q+c
RcON9BGc6hl4kBA4ot1O9H+S/ExshJSWNtNSTDs5gzPp33T2pU42toPWFBgE548i
JiegUOWFGH+G/4/gGPXN4nxen0tOto5jfIUFXXdTpWEojt11ZiDUAD3/gwOcbBof
yjsJegkf7DU/mJITiwOHuDw+++z7ggr9tC9jcoGi3ECVCl4sZg3ZhHf4JI9aramK
YKKuvahO3q2iQA5kbJdB4S08MibsEQ/Ii4P4E++/rnXsGSPHpIc/7CO/u2qVp+BU
XfnMFEoKaQwHiuhiGJLwwe759aW2xtJh0mTsXFkYIFqdJkGn526xAdiIZUswLcpc
M3SUCdo9oQBN3xeqQ8fJd0O3go6UcJf/rQV1xZE54cT6EfsDSJqmRfkV1cSxlt8i
C1zZf5pyxhwSI7JudBfrP0N31vZCGMr0tw/2bnREgmMU+UfzQK3/26lor1vJy55/
WiO3uBiw1vI905CElUK2pLAW6JLcWrXtyIcCf6kpW0zXtr3m7cy/a/1LHgqC/hHC
VsU3YoQhN2spwYf3w+dBO0kIYph6ygL22iMhqxalAUzRynmH0ttnMevzwdzyrxdO
rQElOXfPYMGyxcaiG5QvUStNvIv3PNoYQvsOA4vT47XZa4e7y7OBaVnfloy5+aBh
ZYOZ+Ttj+BGw2+g4SGSET48kcOm6VxlW6KWNYiRL/JmIcRNKet8J+pLMkqPFdvlO
hvlDPATEiJ2Xb2uMVQM3wpVPp0t4u/YKbaIPRuCvVABDoileqqLYhso5spqwwROM
/yQ1IvFi5mrFpDjsHaHh9fY8XhTp3wOMejYU6Wbl6VfP4zyCTAO54TJgi0jHWKaw
+TMuQKAK3M1lXfNyuWsDXNWs+uc11BhbYibOs42DJNFrc7hPiGWUzk9ToHZJ6C4o
RzxXl9mwHSOkVstStzJlf2Tj6jezscJLvPWtESPkePiWXfWX3ggdu7od1gD0E1tT
bzb8bAJAA2x+sz2VB5ScUQ1LO/TFr8jxCIXrvv777VKEjMTwk3JmAwMR+pQutJC+
wpaegutuDa0Un34A9J2SVcVeA6d+99stQcFX8QEgAKauMEHaGFcVJM0KqH4YTjaD
/1LOCA6B2Zaq6ElyBDZdDRBV7IE6QfBdAQg0i8e8WYdvRZFuTbFzPZ4Q/qZQRw/7
CdAMDz3et/ZwkURjP8wsrTUWm3hZy0IOCnbuXir1vdoakewEVRjkh4RnZ392l61N
D+h6ksgDzPrIe98f5NG7cetAHKoExAPF1E3gINqXr/m/+J7NfHapQEwMUeJLtchy
pDKRKfHMzcqKbHsCmBKdXXybARfI4TvxhWjT+JrRf08BlRSDYNr1OfOxmW/5e0kq
jl3Il1AuLFX0FamqXPEDgbhDWn9nSW23I1MzMejyahl/0adPIdARAwt9VXKeXbZE
t9ZmxsGCLiHFEc4RVvQkC5wuAmbqTzypz1WypzPxOdIpdJnuPQ+A+mjeJjD2TlfF
GP8f4blpPfkZtpsaynN/IwP1pu3WfTKgt0xacmw72DFipd75lxpFw0OyD3+IIpZg
QNlvjLiPMlWrWgjl288phxPvShDBaDbfZRq/jJXhiH+wRFdvthh+u+QXerH/mMGs
4Y/WNQwv3+RhqMP7qdRD3IguCtQx0oA2aQ5U0DvPYbij2WHIOaqT8sy5hMHc51X4
h9VxoALJXjpQnWWJ6ck2xl+o+7KqkH1mffDQ3W4zxcJ6nvbkAtTvgajbIXUKEPKf
r57smFulo7fAQw8jOJX9WaD/9EOGgWqkaWD3nAZffXZ9B2vnCOGHKViY315NpSVX
JI5TrIS8rdj3MI8WCGeWwYG1UO0U1zrEhdBdiiSNF328QaCKW4/BmqsxUC/Yo1U9
XuYf8nor0ZJECviYLelZ+otiwvGe9EEanWZbXn5iDoWcr94PCstgpGUUfSemCWwd
KZK/qW59s3QEliRxI4O3tZlY2eORnBiq7ehQPRJQWHtL+AK/dXI2M3Tvc3+dbv7b
aQblKNBs7ZhRGSLFDq/x2WC//vJEtP6hZsf3d+m+pQlsmt48WwyK/x0rYJgw7rG8
tzpo8Xue07aIv7NQqedqI4gWPdxJWlhSFH9atsqw7m3IjFVlLe9V3CmOUURjhWsO
RgtvHnmF+QgIWCMwQDIZ29L9QN+qtYoi6z6/TyvNn7/O1YEHmBZo7bSGWTF27Hqi
0tdEEMK/yMvDdB/6B5BloO7Q28ogqPBlRfli8Rq9zJu2m4/M41iXxbogyDl2zjhF
gBZ3VaZExyJY2a2gpecJ9Cz6F3/Zzqj/+jNxQYH4mvdUygnpkcXhy3rxU+gx/Frr
fyy7RTb9cqQ7gWJ0+we3bXgBrExCcqCsvqm97zT2+fPqHN3EIhXjyhLHYefltCYm
LMiyziK559r6t8/gz4pPnrUd4apD1sutJII4yxtonVQET/P1QGPwt4Zpa1rdmley
LoPsUo2vpe7e1B1PuN4qBq9J2hQT12s8dJ37CK5nDYnYSP3dPq2XUhpArZRupIdJ
YIF2JBUo8LxRth5bxvqJWfCIMlKDuUict4V71KKrpp/5jIZZKRptbZYSRWS6O9Rc
EFeV41ZMCotwkiWK7dH/77BnIxIrh+r+l5DSJ2ANIbWdTMuQKOsKByUqadVoMUaZ
/G4uOqFtp6gFTs5j1xmZqRpGPgrLVpyYK/4whZoTI9Jz6BAzFJMAniMpXHYmB5Ko
BHbenDoQkDoQOfyiNlZ8/0vxRUNBdIy4sgy6olkA6oLOdXM8k+x2mLQR647Y0hBc
Z19I3uO8Tp7HSb/7ZlFIbd+SGmlKmF6Dccmf4L0atYR7Iufwi7qU27MCBmDRVrxN
PqqIZ5Tpt22FzvrirOVRceb1XEUzaEeuQWnJFImu3ADHhFX9jatS1sL8WDvbfwCd
x+8jNx2As1ooGPD8c1sbPpLpcGQ/qUAYGADfB8kZe/KbSBJVaR09jCWBzpEE4qm9
1b1Ti1KMXql/9S1qfxeIP9k14IevzxpeGF2z/XYptzLRssTU+OmF6Kz1zbdO6VJ+
9JVq6ECfoWLlzWhpbi8U4FEBA2Jdn7wEfMJ08jEHjAYkclR9f3vwIaP5IJvsDw/j
fzZcPThhl1cUQKJPVvsRPvRLDnwgeyzLLxvPUjNw+Q55StiSAO8uao5nYwjr7Zni
1lYEogy2k8f4y2IyeMwSygEZPCB4h56jyIScXSIdYH59dXysNV8AE/anq1UODLMR
+7HsBwd4hHwK+CQDiS7a3ABvoj6sIGX1oEKU/RcsWBaOBpZtCv47sI0CvMQWEI5U
/QcpM7CZvkYkCalsrnLuGdQ82SohiNVCZKEIqFkoLigbL6wFUzxGrKGVAACWGK/5
pErw4MpA3wsoV11NvZ5f0BvArc7q6QmzCM/swRl5WT76tHKdEu05k+5iPGIxPM6s
T7sX+qUQ6bocZV3s9F7VqnYPzz3l+fU9cWVKiDhh9bhTP3qr/LLBucCRpMyukvdS
63S3iSNwoHCREO5eUhyX18+u6gWJQpm6OJCtisQ/0s+7k4ZpUHNXEGsENK5dv01e
FUtm+B1rBQFPSGB0jdtAVVli/965zJQhOqx84E50A4re02+xAceNFNIAwyUUSV7F
WLzSFlaUgVSVH7//PtYJaw75xlIJEye0N1gR/h+ULpAqhCbekJ+MxvLNCoE+oKPh
sut21oXLhPSyULJvMDT1xJm9Bbkbdt1o6WizHZIIYqrd99W2P/b1e3Gouq4c/isI
R187SsBvM/bQmxyzanrXMeTNkWcuNeolOOYeT6mUloXu1cRGMy9EcQtBe9C8IeiT
GMotUGXExo4ZxeSDuA8QzD4ljtNNI/yDF2lituOkFRB5xLxlfpCgJyjSxM6ImtQa
z8uMu5t/3gI0HSBjvhWO8mhZssHMVv/uMRyQGEf7GTBHu6ccWYVxOtCKuHw1ExBX
lvoNiGnafZNzF52oDNt3oWyRQ32rds1XUz8rttxr4J0Ewf/Vs2UNdZJqCXGPZ6bc
1a5n6RJ6lywCYF4M7SsqFOudmASvGY1/jYkC+UTDPs7S2PF05WqaJd95xHqSpYdK
se0H7M/ofJjDAE1x1GFZSRdbE34b1nbieA7pu77lNjv0BIRwkCBSlQdLJAI8mzGz
OXve7Bwd630uE2MN8Kf+Fnn/bCTPC+PBvfjLpzdO5Q2nP7DyalYlXRgQevrmeH/v
YoWZIZbYrmHI8LorT1dI0TrCglHyaD7RmWe87lz+2NRiszK8FPAxmPfMWuFWRSOS
8C4t+8P5JbrgwvkmEcHSObXQd4M+ESfs0djxgNt6/ggIPEDuF65xf2DF/0/SJ9q4
n6uXau8fhXsJt+sATFMioT4tuf8uk7maUwjrpMjONA7SKgvGlWhZF15RDhBTf2BZ
2ErVOtzj800out5U0ScUWlbpuTg6uuH4lZLYU/eKBhYKob8QntL5Ykqxlfcwn6Mn
SFg7/VV6+wIUtleYHlck5R1IqYIADLYhDFJ6mKjq5nk0Q17NJl3WmzLYUOEgqpPb
SvCqqY3RkHfZJ1DQDExuAY98bZZdgLJV6+jK2CDNx8WkelHwA6WPiqPhbyGeTwFH
/Dqn4hY7X4WV53gDFQX5JcOCZmqKy6ECGzKQFJOxglenw4HMET0Z72QgMv3LPaPA
R+Bj4WCB2LPRUNqnxIGAO4wO5NnA/7MLJTZvrtZJPv8O2F+o2EGlHE87WGvSm+2w
cNBTBCjPiobGtFCl59husE+Oe34BqYL1XWPGdplrGFL/Wsz0DF1lpgkpAicYGDnf
mYPnfMFGYCJ3fFLtxBFpbz7kSYiROXt25zGo681Tr6A6h+x4RvMUarm4tAmmh4t7
yzrzmtt6qBBlPf5ZGGqnzEUP3Mjl19IQW14AiJZpjbwqmL53X1Iv0hHSfodgm0IH
mxLAZ+55eQFBEvHxyhfiTlJWOw5xmn7WfeB5F+gtlh7T1PPliEGnLAh49MT0s/cZ
qbjdb/Mk6rOP/DZOztimzf8e8ACZzEfXyB97R9FwJGds+MMmFnK0S+e1igDGQqH1
/+ouGxgdTT51MAVwdOP1T2RCdTsfbwCaaMdymeD4S3WDGS7Qbeg+YR4B6a73SJ9O
d6QGJVuTd9jjsX6CwMPQiOD1M0wpfUby3MSfOugxSxImTWQBBry5aO0/GKmRl/tY
B6wN3GYZibXEJTxiBUoO5vhbvwCOT3GXdTLDXJbFLF8ydhjuSZPNc4SsgKQFfnAm
1cZD9YfO/nwcdxN2qJgk/IQnh2GAd56f6KKfsj7Sq8H/MEGAGgssi1VHboATXY/r
iav+8QuUhETrTyvXMvusEzDO7SpRN8ILJeo7MXtfEp8SSF4IzE/taZpYMZfBPXxu
LX4pKP/B4aYuIlymFn9fEOo2F+Q5IM8oK2Rm/X4iqwFzkT0rH4G+gEJSpjwUfy3J
laHvc9vLMpCX2SReJpIit0I/xBZ5v5h2cC1D+UdhuHPOySh03yc1RBujbELJ0n0C
CU3M5AoGz/h2s/2IK8i/k+/ScCC+pYTNJ+/nqpvnKMAoiBZvfPq+4/llR9sVpbt7
ejAXDuGFW6uhuiJaxdhdxZp3drRq1pCuQoqXpQmXa338X2nuEL+nPrWMNW86w6U9
oiyvB+4II2Cjyy+BYpCVjvAv3L5n/+kjrx/Z4PMvfSMbTQAbs4BNosmPfn63VrQm
FrRS4orY9AQ8YcAUPar6/8No4YLOnO0bk1Vpoa/7ior6yZmjGh0by6v1TtAeYliX
VOosMgJC1qYLUdQIQ7bQ5pMVEnoSKpUq4fZbqo7Xh/ccUwtu0UceUEmT3K9/q9Ze
akJ2R6SnTz+6NbLwC7+Q31nGGEHnr2WwlRSTxjWWH/Pv5Vy7IR+dej79hzJaCVv6
yIYNnE39RIvMsm0fN+lHHvm0B7+wc6cx10VdjWkaeWiK2E2zqW6lz+MnugO3Oidq
b7WBT7PDJV/N3zfgVeCI8Kwp6eNf49FzgCOYt+aFQufOGd4MBBmhnyI/3pzxE390
hhgjmzPxxXnuKlJhcfOUpjWel6BLQGT3YJTP+bSy7VqYBpQRYj+uGO9kgIOWtjtW
s+EL7jHqMsHbM6estwWv6sALGhmN8BRESOf9T1lnK4NE1gL/UAtsXgowL9Pkgr6P
rM+1dY9L/P4EZmTFeC96uMKqzax9YrpwXbw215QiUjSC93VLhoutXdbKvunNU/YH
sWaJbIcnrj76Trz+qUz/Gjuk6REhl08MuTTlJ19AAPbqyjuNXHRLbS3V1qM4kK70
aAxsjSGIgVWYAQai+6BCyZ0nkVZ+6NI1CxQiVzu18z+0Ztohkz6NyP62LmNdkhrV
hiYqiexzlqPquJRzfu77Pq+qIsDfwWdE3qf5D2OR4YBdV2ZtLbg78PlSSrbtrtUG
V13r1i/Ia6jFn3rTQmmpcWEYvwEdzLgnPqC6pV58kH8SXLRejILuqvx/nUVKVoZy
Z9Y2nuZqnINFUc8uCeRUgUEnDcLLHSbXksZybuB4ai8IyUGwqvow6FLLLzkTt3dI
PP1juIsPr4TuuvbXksndlaKZeDDU345gAoCppLlOWX+JyVcVhx9OGNfDaes49G/G
x/ybNm/G1ZAs08DMbQHvF7BUguG+Z19ZX9IioK431NVGw4ooM25CWYi8WIPoLgqP
IEytNWTBC+25hXf8pyLaNKZh11gw8XkEDb0mmHJpAX/s5F95ypJh8qTUrV1jcw5g
sUcMDfHOK5EkQn7Gq4ULLqJ1LY/9hh76gX37mO8JDbPrBxRXEceZLBkQRm77nLC2
dhfzjQuVm1iF7o52D/o/mE9XDbggYypGQ9CHSa7u0fh3m31VZRLtLRqxnzvTZlJg
jhwtxhmyON1V1fYQklQ5s17wtvydAbPL38/rL1Cl+v8nIDWCj+5cFWT9EyF1DX1o
s8yPnA6OsxNTCYRZGwhpNDTXRv0rSXccZwXawlpiL4nnBqqlVsEV8ZRHJIgtIDh3
gGyV5391BZkFtd1H1M49lHLr2w24rl9MFaKql/DI5Vz68aOgAJIfHxiwTPTMeP+K
M47jtSG6EeGLpTn/D4/y2qUifjeNEENNdkS2xRjjufUEdKQ+38b9KS5Qsfs9iIUu
74TQo2uH2xE2K9PBcG9emHaTJWz2gr7OYhNuAFk9jytbt/1CSCLlkeYLnBzmfQdE
BO7TlpSdcsP3vhpIoBInUOkTzSB+BjwSPWNbH2cf6PgRoHosNhqWwOayKmBL/oy2
IL5HYzNcgyiY5QvCpo1XbsJqTaLcFW9j3T7FCQPwfhM9Sl50Pupk0sUIUUxgl1SI
GR6IhtrZ/ypXE5KYwT2JBNvgBj2My4FHJqiwsDYcICDKP713kJEkMK85K2P/OLp8
DAKX0X1FhNG5mpg0ivObZGq58LiWaxbBmz8A6nKhHOYZ7sClEDCE+/g+xHnWT6ZD
xTCVKXoq5Q6tuhjpr6vCATi+4uAcUs8jT4mWIgii8cNfsBHdOoj2W49+JwFvF1Ae
XGel0ZRPIkFTrxbMEtwpbJ2ub2NxsxK/lLtkx9myZDgxKcllT/jkwonOrSu0wo9t
9YWj58jZBdLV9RkWDf9242wLbi1VE2XGVvOT1lKkZA3V/rKRWeiPmL0K0MaDSFGL
y0FleWNR5PO+/UwmIzUrD7H4hBHq/hmbXLTAAfR3BgMsidOWAdH5hKBzHqQhtFTg
9GCAYBZXwJrgOCAapfMv1hB3m3pgnIf6SUQlGYi6c5FUT9WvdiXYIfs1IcICrPWC
ocEuWKcrR1BM8//TTir502dEA8QlMgJ/FQSdj8MykCeRDDDWnY1TZYJsnRPQi8ER
O+EgcQ4A9HWQq9AuNmZwznR105s+Vfkjf0gKyx2bRCiI/Vmrek5zzYE7YAnJO7XW
/aOXR7+5C+CZHlm3QIamPD056TAZsNSsw0araNR6GfkI+YI5kikPX266SrijKLQL
FobKNL0KxQVQtEpv8AoCsa480E5oW/B6m736ML8tAP8w9719pv4UPgdn9VCDibOZ
1HqhZXQxUB5OHFtkACXOLSft3eo+ZCP7tOKaeO9XEhLg+j7gcpsyimsYw+q9ef6e
VNN0UIseyXdeaHZ00hobOa7qdORkBQ6dUdEhgxF5e9p3YhR5jc2mTKxFXHWDStxz
YIncS9IQj09bcoJqRNRSrUzukOa2b4oFv5t1tKmvIpPW7ynv4cjAhp9tSyF66AZF
pm9OMLxVFpFiL/2gq3p6YLmP2Vlhk714s6RrEOyA5PTsEV6qj8TCjk6He6xjeY22
FQIGIwQ34wLc1Wf8YchwnlM1gYIwJfmI2n7lXdK6EhGVVr/1+TFMQN+XcuVPes/S
7BB1o0pUHRk9Wk6LcjTSwK38oeHgCS0909Fh8gBkLOlU1TcRORooqpQjC3522doU
nDKPG5/WgUymHzGSsx1ApNZkga6VF+hHhL7COOU79ARTndBumoAfrq1d5qKMBPDM
bXkxcf0xm6moNV6obg+uI6/rBXtjrrk+dBiASJkOZoA6WdwqYDpojht6Xjj6EF9o
Vwc9NRyk1GFRShen03LGtk2LVGsgoHxA960pCxHDfIuscJPlzgOcqKk41tHGsEl1
8Yu0ddSQaxB5MwRelm3H6+InRAQw0yOeqicbE7T7bG+AlDYjjBZMKvQkx2L1cO2r
6JENvM3kVqL+YyQsvORbEVsCDUJnFfqaXBQtXybFpxb3/fuDvbq5z/rDVyl2q3Ix
wBZ4Ob6OW5zh/zMt2OLye/OrfSr2+TCU7dEUOjL1SdGIMpi2H2XZSIgKp52P0EbT
ru2VwaAZ6AsFDfCuEJah+a/NEO23JMyWfzXsNqURipwuNMxAcv08hV6ig2wMEk/p
jHUIfqk0VeqMeCV4OWQBFC3+JII2Y8o3cpyD1qF6oBGb0zWFNccbwTrjEuc9t3rx
fFgT202hArBjBc4CDvKslXnX9b+Zxrt1EFX/9GRXfQZbucEvcsmOD9401ZjRJldy
+D1bKoCRNwYTD6o3TZWzSRkhMTEpBse+AekJVaQYlzVo3Y4/0QaIGHJJLtMXRDUH
EZPUiGTdrbtTfZ5vwAZg4Gqm6jvvuBn9BBpqH1m30zbLNlVNoTmJGm7V2cWuh0Jr
+UmvIgJGAwomfjgCYbaARNh6CjZYrhgYX3rn9Z/S2gxB4k6kDzwZOXwdj9fVRmD+
47CfrlvzNOdAhiQPiiu4yx5FV58Y9+Jh2cWfhqinPm43ZjfMr58Pp6qeXUkBdk+c
RbOJtUX99JWO7dJcesI4elaBWQxWoAf68TSWvFuGpi3s19nU+Pw+hO+VJzOt6U2m
VYsMqxQmPWaSLa5YQwMSqnqcaZPPPfM1JZaYp+ehxhUT3LUuP45JSZHQ5f0nYnmx
0rwR3npteUncsH1nvOG6J2QPYt1AB4kVC8MSc2UIjAHvHe4HjAGdM9ITVmC3IZbf
R6wZ3gQRK7A9eaV1XI6zVfNAeqhbteBkq/gHkcfM0+nfo53EnRViLQW3476/sQQ4
L7Rh9RrE5L7RqTyPaNJLa0IYp/RSWdkUIyzCL9ENQPXi8VnkRD5vFJrhuRGvFm8a
LDBmZKUtabjGnVEwcl1YnL3GFMTKh5hYHPpK2ksOV1DDSUvLILxuYuozkBXRyZN0
LS+8NGTjL1KmC4/JZ2tsDsjgV96nvRMXaA1cig+asH2cMTYkfxpTOvyaDF7C43G8
EVUJV6KhEUZ5r+RZUqgN7Y6eDFgLAx7EUJ4js8h1EdmDkDzDxYatcBnq83bJKE/e
ljOvWzst1mCIEB/bYKjoyKvXVjEpmpYbzfOaFRubs+cDSIYiaaerhikbDE2e3+74
9hLBfUGRtAfFtOXvAZ8sZkPg8gz96Ptb0ZKN6XqziL1cYI2F/j4dkCJnVTlMdDza
tdsZXmSQsENmWTKuAGy9PFHJuHxukFjizOhQOvrvqK3dHU0+Q+BJaXyJJ51og/Mw
f5DPmOEzC2xbJDgS8XUFvnUqxiGHojt+SnMudccH6uh0bDTba1yp8h9KGcXGzy18
rkO+LC/KHRKLLjuIiM+5HYPDAdcWdNidpOAEngAhHQE6scB8siQAX/bxiUv2AdOj
+o0jvVl2hcI6+bFlCb8BKg0XrRHcLcpWZM9L+FN2Yjax6QGmjMapKCIF8iqmXXOn
Nz/Mwgr9/EF/xYmzMJJuaBJC6xduNQJjFFh2IRAsQd5OFLOHTfBrdUzbrWsyelL9
PKDUGHPWBtHiNmv8jYvcyZezRxAq+70W85yJst3KKOdHLyXZTX3qXW0+HN+etQcG
Hy/1M23NeOeGtz1fO/xkjgIZ/R6saVoRwHxnl93JrbIdNhd9Gvwnx4K5MB+H9xh3
sLIZImVhkGaT9HXvqhShzslEx/35bkYiFHrDJTrPoh6QTUH8n9PNao+nk0JIUkt0
trHNMVg6sOJlte+4USUdDB82f9Ev0p9hT7yp9KcJYL7xYIG3b9obQngeLATraFEI
PwouQUgbZSC1/rqiZIMKNXlifRHaVmw2o5SkxDPWgljxXPQoPnNNRi6sT5vL1yCM
cPyCQfj4gbXy5vOnbAOdMvKFc5d+qW+bJlOHgCpmRrlPZTs/N3DlDOOsaNFmTpPv
LgWaz+zG2R3t5wGwZOb/yxka+e41GPVb2K7Req5pvOpxPkSOlk0hVwGg8uOEPyPo
5QCdxHl19D765FcB6tUYOzz0ICgPWqY8gaOBgYG45p7gDGY8ZVE7ewt7Au2U6q4i
T5Pd8+FdtO8Sip9yEge9JHCK+H0XN7UoDPF+xv0BCIEr4xSD/dTQV8Z3+RHtJSSM
mJ8Lc2HGYLrwMMagMo06cPgB4ulk/yuTnHL5gwxt3o1LND0iayQU2Z9Yhnr5LbcR
7F/dqRDmrGkn5SrO/Ll4YdOJrWIcR8WdrA3GjnV883q3tfYM3ByQqHoewA5wk+o+
oBJtHKhI8Qh+9FmabNSwxdD968hVsQI8FMZN/virYR9//lYL4skhBYj9UucWPh0X
qfQFmUQ8zhACQ8zjMoEeLtM7UlGldgvDKYns294HavRwN+ClEkNOHsIE8gcE/Rl+
SLMuiEfzo42ajrwiNrTx85Tvie/ZTOqos5y3W5Ej5Gdt4RZz/hAc+yD1/zG/ygQc
wjJoS4HvafvamNBeGA7164vNSE8kxKU5gWuBXrhmmU29tCVtz2eWYXnZlkB75d9E
wPO7U+a8t5RZyCTvQWupF5KkPo5y5NIpxdScd74dhaQv1NUXzBzCfa37sc17ceZd
KXFUNoPARdwBLbAtH9ScqHv89Z0QGLPdjkElF0TDoIbiREy3CVFy7c0zTcL8cWrO
zSZrraM/KH3q0wFA//H9O6QQA+8MWR8hTvrsNLMvUAuZEsz4clYpWhu9/rrSEtdo
7AObjRJsECu7gDCcbFur8Fci/P5U0hrwfRn5rOg1M1WVY9bUYH5AcR1M3kPLLFwT
N7mnuVycNZ4LZ0ZXTa9ifDl9DmtsHWgcFf8iAmu3QCPqY0s1ySg47uO/ehT9DsMc
y4eTmY/oZRa8Z+NHVOhil0kdE5YFXwDL12Rh4MuPwr9K61pPHuRCan7KMrpXoIc/
AgzW8CK+ATzMqLZFHmoVaheYK+zZIUkoWOta73nGjv8wv/4m7n482PpDi2AElfeS
iIWDL7gxzeNWHMWruLlWjd1qbLIbZlZFIkIRAu5Kpdzdro6deusUL+CLZOVs1f6z
VuKqWjAHCzIq7+ekR6cp13jaQ50JTd6pUyio6A2M3vCTzgBnJqtOPdOCLaCZS2EC
+N9prhalT9k8keVV/lam8cu5l5JiJtMUkJrLKxg9l3tntrHrWFB8eM12nLWO+Hb8
JNRhYO+IKLqf+rNat3lcqQIUz4Q6FmT0WGYXJdsnD0eyH/XFnPyJs6GgGhcEx9hY
Wn3JtwDn9aNMA+jbiUWpKHicQVJArfw8Vix5yODb2tSu96aXDDCd0gsfNz2mOXSU
Zz+b6xalxslmExrWJja55wNGZt5EH7x3R0rwBSqR7PsZnqK6jUuZ5nUCgQKb8eOX
uPXGA2UuWzLH4wgX3RB9XMjZI8V2ZwNuNR/gfRnY+xcuPtvUEklAo8I5QKC17HF4
7J5tMjIhXOG8lj8zYLGdv3+PMQC/+B9L32N6Tw+X2eEl5j0HfJP6MFyIE9i3O4On
4oJxlHjzYrlAYbk0mMryfmB0rF/xmESVWM40mT+ChI0YnS/8+jV4F5uycvaeKMVl
VvecGtZwBKh0y0kyRGvIPtNPyc8ZyF7Sao/glon4+dM/LGAXili9bYpmJ8Q1WMG+
jSa0xUjlvsaQQx+Trdzc94nqSuad8eu7Xbly6VjVX9ezusCIUSd/733QOEBFc/WG
H2Hf9Ioxic2l5+eK2ds750xDUr+2vN6WtYV4yaCJzCmFOQeJdf6kleEf6kvvKCYd
DF1bBQD67eM1b8JhKxQ7qarWxT8liu6dfHvv5nU/blJP27LA8cz4qtFMXBBWFmDC
IcCWVZUIKR4mJA+wzvsd+6HXb7MmS0MyPH5iJaUFWU+fjaQ3vb86vGG5RrgwhZ5v
p54E05WborwGqkP8BFaveC/etB7nQGc9A6xue3+o2ngBLu26cp/b3e/foMKNSVeE
WQVJtMUQUCoCu+nI/DCelxgeACE8iGK2jueB4jJMSeRnue4RDTuE1In4frgTfIkB
fo4eEygcTEtHuEtnslP0e/QWd6mvAlKUAM2HGYjvTkNH3xLVceSKQe9xMOLs10/U
tB/CPE+b2Q5tkIoz1+M6j/4saE8MOiYmDZMjGFHRDaMtLJhG7DW7dEzgwhqk+yst
4tpL7NuYfpqYVtAVS+tWN6YY4Dy2j90ey6zefIZSKkB727YGzitoeW/DxuXhqAbw
yqYglJhTehE33uLuFmo9+cFYbDnHxxPUvKqTpOdVRgPiHtngGsk7VepDXiFrWGqm
87Lh3tfHVmQG9AEtBVppHbvKFHNT9ayJQVTZ3JFFh4JTHDDwFK5M5jYcSASIJ0DW
ZGVn5eVYZNq3X3Yr3wed5usArN87grPZYgjBCoD1zrqniyjgABKRfYJ1nHkE50WW
A4pkD2KZAcF7Zy8oNUL0DZrtxY1hpDvBkLtkitKWbHckDhIapgi9em4IwlFsx1Ne
+bneDPnjN3R671JVLya6rQw1WCYV0H2nQrkqxcOZkWS7v8vuCoTSMpNQ2MEQaVGQ
LPzrpOw2uRFU8HRMUDDRE7N5EVtWZ2beUos4HYxbqF/6DM/dHTR7ZTWqdOx6VLNW
H928Tw8bXW4HlIt0yRqEmQtBs9FbLuokzkOmZ8pAl3OokKfHH6OuSECjqzCnhx+n
yIvwhufcEDRuFGuAxWQCwD4fFlrXr2dL1lQHFkjDqJG/7QqtQbyToXuyuvJMGDRl
AEEwQyPL2YuHyLTfT4B4MGwNODKeU0P9JxrwYdUfXmdWbWYxLNw2ElaOHSvvhsKy
AsFMFaRIiqYWOIAz5we3kvtpOHJynVz0l8NslO8YQFHdwFUvrJtgvyn8tk4WKuib
wBWCQQHOtaXUftX5xFLceS00qKepRShOAoxrXcXi+NmMqNeRLByPDba+/z0WJcng
Ru205qs5KCgurVdcanfDaP9+qdpB1spRGxaFERRmKcv1KN5roS7gi8798tV53+ck
OKSKb9ANSoOe/9fRhoOFL3YG6Ob46g1sz9dyGuaoAShfuQ20Vo9LV/UqoYqouu1r
ToZ9Gd+ekKAovInGQpL70wkzt5ia226bc+NY+2pDQk2Xk6ziTwZrrPLzF2P8FTpS
BIVq44R3o7nSeNpY58Vg9Z9CEbA1mlfSi1gyCIpw02k5dPztJxCe9zWDxHd58YoA
Aslu/e2w0dudc4xR1pdRrUQvBW3EGI1LGpMc3wl48odb8X5hXEECRPrBH+E5EoCT
+ZJeA9ycSH9FILHc0nstq8+6fHY57VS8WEDYpq4vCjnK+310Ur0CHqs1stl8c3Wj
Tb8EYZ5iFuMM4NxeDez2sX1kKXmBNIIRCXfXeXHNvTLie6IUNWIVuqThZYwdE0lg
fIQJbBNfsXYqlBsVTPdMUliKTis7pv6W+AGpTxQoc0KpKNdb13abMqjjEM/9FnI4
FfIaT+EQ0zajVUiD20Rhm651gMQOPxHohJ7h4Redo2b8RLnENeEMqaB/aVDYN4OQ
C6ErQGWPAjpPOWqv6pUWKpnVDNxlJcTVkQ5F63XvEKU1Hd2uhRS4v8RXz/ucJwra
5d0y1qpjZRJDRjyaCiET06XqfhRlBsb5MUFc12p4nN8PnYFhE+0bvnGTn0X4V+qc
cd8D0mgW+0rFeG195pNrCpnRMdq5st2HTfJ1JeWGpLSpLtL5MEQCzAINMPUq6WXE
XMeRLy50pylaVKWPIL2PAzi0PX2roqHyKqS6CsuqY+hkhfGFmQ9YCe8xtmb2ICJ1
L1kJguXhvFIosyKMd5LG1db/9ARE2t1HnUTvIFkaDlNvp4LjSTqjYwYt4sDc7ZIF
4VH9CAsLnDZcsOU+r3g1Jc9qxN45PmcYbTaEOcGwAGR7sGXNPqAI4JOP5WL0TwiS
c4aAM28WrjNmtP3f+3IYc3SbG2+eD2X5wcUgJhc9ZzhKaJllSfjTcOueC3txOq6+
htRBzf3ye1ShLc9uSxpv6VMJOK1IX9pgPJbjuk4y83gr5P6/T+MsIHz4QFU4EbEO
fJOEFNTSDAYfK/MQ5XBM+UmY3Hdtd56Aah/NioGlGv0zuybMdWt+M2xFkpiFheHw
7vkpakj7IHcZCVGX4TmwqdzSobzTHB1F9ymom6stnJlVWCF7ZIcUotwdqx8zqAKo
no29FAbEoF0OCYiASIcctfgEQkgTtHkQkE4/FjirGT2lyipGAapOfexzbQI51JT1
g1yeUR7jNOoiJeKdh6OveyX2MPEQAX3u4X7SXFTD5Sb6CIThrE0nIh7/TvvtUKs8
OyQuLAP102jVmHuVwM/mMnjY4zDubC1NYaw9zg4yfnimZavbbW7ENlgZuBzkeu/I
UrDI5XMQNjyuXqOtcnGpiBNUIJbB65f7OQ+bFzuVBrvWLsGfXdB4QLCG5AvZRqfn
t1909/d3lhvigD3GAjDMyfnX7qcMcCjZFtbKECZKCQfT27DTYb/qwkDeW5qHlsgk
CmIACSjDIfMeDC5AIB/gKOX+zU9R9wR8SJXbTpNlZm5GAUWyCzbrgX1Lb4CN3MHW
cpKweic/jSLqeJ81xA3Ejuwtn1euxJrw79+zGadpV0xY+oofG95EGReFARSgNZp2
xjE60i7YrXH0sDS04T99fEZ/BWomA9IUnJyZ6km8QYf77UaqiaIkdxUnCkh5hXDz
7DJRgm2wRID2y1ZYvVID0HOs/Kj3Tk8xBgBPGcFR6U8qDWufHojcvzoDLaL1L/aR
qWc222tz/dCAAWHJeeAF+dL94sZHwdC0lp8ipDceHIPNLj8KUD1+eX2Ups2nysOZ
n/r0VLOsJ0dte/W1ya29BSC2eJMPXvdipIAX46lilAEoTfFXJJ7BVKIefTu6nyi8
K4wtWv5jrVlE5hZCG67E/5vWSZfQk++snqO3JnNUw4CubTZ+6K1bePDK9D47Bv/k
ztUYVkWzBF7wOxojoYKrcBTrtbp2f75YKMZERXl1ME0NCuT0G/khGLjoYd2UQQox
yXJLEKt159uBUq11y5uYzxDKC84h9ozyQ8D4kotUyhB6kyOrITTZC7r2EJnLivjp
Moy0pYdjOBfOJ6R3Mnct8KCjnsckTWjoEgJckddNRpzCZz2I4sit5+j2883eWKoi
VMefS4fkFvlXaXQf7wFGR16SaAsZzfxcFcztHU1zJ/RBBSky1GfKUaqa4L1oNbME
2vdD7v6SjqPVXGaGZQa4r2R++jS4JAlwYwxu6ntz0LgGMPxguhX8R0j05pemx5jj
/6DwmcAboKYNKGkOjP6RijaBuNjSKu6TEGuUYvk+RLxCA3tzImXfqjI3OXYZh+Ul
amcKODVkJxNXopghEve4kVhkr0MB4RsDskAlIbqODSyBAihdLlNv4VWgTESq0bdc
yVQHE/Dby3CXaWAuzCcA5lGEJ3ahEOb4rrMzJZ1QQAVrQdqQOqcs8XRX4nsGoZn5
nrlAxpd1dpfz0II2jf3fNa28tUMQ40ZS1mBJiOmKfKWDgf8m0FzfCI9qm41SYTLj
ZQpMrdXoLYriSID85dD1zK7mRDuAKunPyTxSK9sDrELM8yH2L8VnTH9Zh6/FDpmn
0/j9QqifRKXBm/tw1q1FfMOp7JTfqEsWWVXVaLlzP79mnjHX7wnsDagWHrXiBMFd
Oy1kYmID6fwR/bRp+O8TkuEvpwDHxz5v0asy/aqr+s449Uc+bpcF95xdMfyAV5j7
rlHoZF1DPbFwpWPKY3YBmIH7qKh9ZKHtUOjohM8ScGbpXhW17RecbGoBI6cGxJsx
NRMWE3P9FuFkX75ORmu/iazUMVT7HyrtlKADit4T3e05MRNElsgYnaSZGYLV/A54
uEAuL67ygd9XKDfpkm9dwyUSVORbn3OUeITdn632ix34iggJWqLAEmms0a+n2yZN
bRKXb/TkEW7N4pt5nVb4Ps8CFfX0OHUePU/BTMK85auJxcHyRhk73qKSwVLPCXZy
OHlzlZZ5dp6rGSvML8F48A8GkvqHMCPUqzX/XTOVu2nAogCuaK0xiUYfL0nfETVL
Yie8CXNTG4gNrO4Tc7lxwpB9n4KvzCXPAOnLlaeSxvocUTtTG5YaXyQmaoTeTKWW
RhMpWhXS6kL/aQwvpdqgwaJN2AmAWi1tLHSh3Z5WlTu3QlWXXIXxEsLvp8IIcUKv
8/1bU9U3mlaoHo+5gSojh2GbSqDPo36X/tgwqU8ClBPOYua9Q3NhiSYiXxOJZq/T
y+gIbvXIu4jCOmGeIBRqiw7kUvCTg6UXXiTJuVbK3MUZ58M/10Z10izhB+FOvk4l
rwryPwgJefMyRuKbc1WAskz/gnLQXO7MNQMYB5vEhOLxJkAqZyZPwo6fkLIVRIwP
n8t1E5HeAmZA03eoJJVqYc+J0nEZSnDHVz+2c7ikk2yryh83cyyfhu8WyDVxr9Gp
Kd8K1XKuMIXlpLvf8v86HpkT3uEdhaABhtRmp8RpClB9M4yrTtx/YQHvJY0XA/jK
5KXD7TQnsSwjhFC7eK35qms8xDlilRwDMTEJKX/s8qzRnuewtp1dn71d81uKLnHS
nzKJIFQKpLKx8StHMdLN02zJMlzB090FGiJZNUZIZsTtq/JYBNF3YogJ+xn0S063
mDhO0OFw/dYpZR+nevtK5/Gd0+2t/7xmuaRDUymwU71+/qqmaaGXZkjHOqcGgdsr
5VvNYfPenzNXAovrzSjtMS9gEsBE1gw/N0bFWD4wWw4PsqLJ4y8+TdijpAwyAnDe
R4NAYSK239OXHvSe+vX8+ORqiCq91E5AlxhSLXkPdY1UTLiK0yYMvBHE07N01jc0
NBF86bCvEBR/tlFdkodVfeaEqwvhbpS/h88spxyo3h7JUxZTYHrR0Kzvxr+d4Dsd
2HEgwMHiYz/M1PyKHtm7P0vNPIqEv1OdYbg6Jnn6SmD/eT0N+PDtSc0Zr5jmHaGL
2yh9VLKltqE8rhxKsBrKfOAtS3zQDacFW39tqodV3TfXGywYb80pN9e3YFKKiBQ5
5OtW4NeG4zrzGvF3rKtgLprWj2rHvR15xwb4s4VdPAiGF/NKhlMWg258v7fPgy1H
vTEF8GLghiraDNDN6YC9Anh6mA4Ax89/kE37iDJ3ftwLB2JUQBUfUA3HUkdgUzWL
wsmytGh0GHROpj647gTV9pZfvPIcnuc6qDyQCour0nByKHbxV0gJkZykn2FEl8sK
CtSeHqKYG2fXrgXeFesMb8dfx+cwwjkdgYH7cMo8tMHeq4pI82NYIj68HwTB5qxp
sABdV9gusaNek3j5m5aq74FH41ellkv42iAAwTAfr2I80KfeTIqUdHd92UnEBNoL
mHrriwDN+ZOnIv/OE2FNHsKDzYzN8jeUF0T9V2kXwxh+zBMlmY4vofE+r6AjwrNz
MnkfhNWvbgNGHu54/9dnc3H1jFGPqZ6HTjgAP+PSjIRa4yD2936kk3tIag+n+9BK
lo0IoBhORdR+V7XStiRVEUiTaFkmZGWuSTwt3PwAkok406zfYjj6zsIAPBoiHdRf
FvpMdeuh0jbZ8Ea4G4V8kFCUAAec3mmugzLPYvnb7KreAmiAAI6Ix/RiIdrgd4Me
RCsJX209QNyMxmHOIN+hfRJgO7M5hFd2GfzS0htmBwwq7/GHDthAFrCqccsztjgx
sOP5gdwpGFYb3v5S9CW17V9OTE1I8FKFB9fIX+w+hrUznOmVhxIB5jqA666JMCfj
G2AjIG5S1jIh2s8QNgohMwO1+zutAgjW3WWUg66MR0tnz8EiwMKAsA7jyGRY7+j5
hFU9leHiSEuB6xip/Zv6dXS5RWLMQV+LN4R1mYoVnmvxJdR+s/D4HLzClmMmWVHb
MZRbk+acVernRQufIoIh+UdMUtkO1HpHfuBM6wfooe9tbGwZLecxS3MVecBrdJzf
eHnybWQOI1UENftlXKSbqdctDTDB2zZKan0jo8uLYelRafq0gszTNzR/W0Id5J6t
bKS79bW0U/B6wPd3LYyhHnpRH9aQh6/XaR0K8eZb30b4aDFs1/TDgWTQVGOY1/+i
YmNwyPw5SiVpEvuAvdzQHvqhLuec26bD0bVQFXEECIuf7LLFDOh99wYquNRPPJzH
j5pdrkxWN2Amie3Sq1rEOBCUQxzNb9K1BjNceNNaP3AbJhP6dsedOQZU5oW50ooF
7BAemeu5un08/hfDiUvRwmTiQMVZjdPOHOHLjQrNtiXzsI75jJ5ctoxr3bhzctBU
oOzo8WVO3KtsAegFMzudIvddAFn196EL+MBWWCr05us1rCTjtexviIcDY00ZEEmd
4eH+Rg0BMvJqC/K91CHfkYBTJJRps1QHp0zv7jgFkq60oZHzHHOwohDYmnW9JwRF
Z28yCzGK0TpH/sRAyf6o4i4OSmyvSSen1dX8jojXHqi/4aj+PfNWhypDEwIq4OI/
l3LnMAMNjG0JjXJOgWrCNYQWope+aNhUU42jC65OQLkl2lMIN4VtGj2p9g5/TALy
2KLTcfR9es3jYjeHwXLFvY1LPMrOIOVJz/7GZcFvBsZDrTGSTU0C6e8XDNW2ZUcY
FuNOOFtzFoQuo0Z2ZfJ/IJVGe1UhOTj+iPctTWucUcVr4KbZxKBErNzfKAceAMkJ
ODxX2qsPfWZbDMnaoq4N7wR6FWj0Y39i7ar1mYxe4oaDp/3FvwMrl2frIgdnwkyY
EYsJVPZeHk+GMJsCDC41UpEBUkgEbtzifkgs+8AELEtDqCayvCiRXXGo832WENP6
qlmxurdxOXmosySKbIpGMGQczyuf/nhG8xmeP2lhzbtlzLSN5AfKc7pZZjJpp4BD
LLfXbE1P3IU4bRQvDwAzlYcg9bU8ZEjeaA3zP0UGLAcHGTi8Z5DI3c4axmPIXqCA
JaDfO5DnYKnnp0uZvYxlEaDiISG5JlVRfilC7Ls3ivp4NQNqnqchEGpa3OWJ2SBV
ZsI+gkHavOjhYpLkYThNeLjWHIoTDtvBwtpGhdlGWYH7J3TxD5lJQh98W0tFPh00
I/0b6CpuOZW7woeyxZFysxnkDmwNOAcPoAIMbeyWlHW8Jo5ADmkGeziy1nHsD+fv
PSmodvfJ39L9v/BbOMdxDpmw1/bCgqtI/kafBoKVL+2id2ADPq/i6oEixFFEO3fE
xfmXGhZbdhztuihB/sO7b0NWohSa0zJTNBlwIeQenmscXyJMW9Sy2IUMBIDJ8KhC
Na69OTGpzr1Peju/1y8VJaAIDhu6b4Aqi4VMxMvi8nbiEcAhyBKTFCAuuXIC9E8G
Cag5sU2n3bqbSRZBJgZLZKWd3pys6rpKzPUusiz9Yig9aIInvrZ/hhAOeRTj7RIB
SON3bc8E8eHZ+OBEeeboEkkymESLZA180yeeuxtuWz4ZHdl2OaVn4nAZIb8S0ajH
DUMQYD3CWORqYfqXCSa2GM0nxIL1MDeBV261CjSBtNndURpHwZ2BLV5Azw7FLBxj
uIKrVuPlkPrCg5+MwCHHGRJFQUNSC4m+rhD64Q/YKwphLIGiRFof43rP+fKMLLHT
RTj6Boy4d0D+r2Tcz+n92zoKqtpEv+GoJl1zJjRzDomC09/vf6pHEW7UGP+T2VmK
7XtFrvpp2RlkWYe/jumCH6fwzn4TZrfiozz+B8jntoq9q7tJ1nCu+jlg6KpBRi/W
jId/N9maRi4m2ncfRUp8YNDgRDb82SaI87qXW3Il0XCDA8n3UUaeLbhP4ZZLSK3X
V2vWWNEStiofWBHukfDErH41yUIsdl/qRjUVlq3IACHNp+i+gA7r0N8yowR0j5xw
woVpj7ik8gLSmGxFfxhQVOb/LE9uCpxfuMpG0vo0HPqiDtJdhdJkmBaS9Qrw22ga
0uYD4ENXV/uRFZp7W7IiVmIsG7hWshtBaZ1tpjfuLEU48xdoKj7deucnEVRpd1At
lOtB4cRQ2JLaPfhFr05ZhZP7rqf2SK6Hj7ZNeRTeNLMavn/ZKzrcaW+VLMcymVNO
0R7LsckjC4oJ3PFVEMPR0C7i7uQDO9wtFvvC/Eba5jPIkQ8aesP7DXJ/DC47HCPo
6CLFGtLLuSi0bPI6FQ6X4OltgRx7/IDOeHS6R4YJ0sZCto5q2VXNj4GGvbnS4foK
6UrgzqMRCbpk4ZYlDtIdQjuhwJ3tfXjkOrP2C75ELobvXTrDJPP+uy2Ye6Lub8TU
qOlck4IxQ26PYJE+/XhrpSiQisJYO4LUN8SR8zGJpSSrU12AmwQoH8B9N48JsHOi
HdFRQqipaZotnm+nTQ4oTdRzoKvvK9O2JtUaHA7NSmWnDcDMJ8XNfnqiifzkOyry
nME0i1yHO6nkmPqxjpDpAWdLzcEIV3YvznufgUlGRb0mwHNJzWNxms+oJ4RVjW1i
gTEX+ulXnuszjrL4wZ59CuSFevNig96Svj/JJJ2gOVo7ojTorvmFU8JPzuv6SavE
7K9/udDnq8mlbqIeO11PCjUb4bTGiqjiCt8T5ENv2pcGBbHsto8yfnImh8GfGSK3
1dC6rFrYsqWiTRMqTpraQSaCV2Zddy1pWtI8srVNMi9INSoVP0CMgsYJ9YKBfS1S
vLgp982fHbS1dWlDl1AJ4hZAepQ5jMJHwod3DlF1blr36/G6cf6U93BZx/7O1Uj1
mGO2EwZU0lyJmt6M79jbBcy67rVYoJEDGVAepxIVbB9mI6zMRUGNgGIsJjTQ+CM5
+NdfwibsJGkEDyNX0MPhRZFZ6oROepbZoSsvRhbp+4u/BsMCfLH+OIZVQ+XSQcKp
Zq0CLUs2gNUC+vwOLkXwA5ArGVnhe2qe8Trk2x5Tn4PJ35ey1+rb2+weodNlL55k
/+min4uExoIiywUT9ISZkPboStHSSRchvUs4k/ce4GVvz8mhEfO9+gdkNVjMAOry
APCQNzGz7QkACLD6sr1NZIPWrFB6Wk6I+BFgVBrFEWRWCojmhy01KalDkwRoEQpc
VwnPDVZX+O84aUpDe1YucBlo5dLkJdRXDOs0jS4etqQOKmYU1ZU7bTI+xQfHEOUp
2MM/qhBR4fE8KG4A5W8qIa2W0gDKGIapsc1q/MGy+sGJ0m/gZrBdfQWPQ7l2I8Iu
cP4Tj3W+BuoWxGcSDuwHZdnqqh8yPsuMeXj5lBSuxhk9U/89YbT6RjTHOVmsJRti
xsNfrG9X1njCPmtopbHRmWKBtq/x2fJEZHHAPxBGidxX0Dsi/COZGFItNq1VA78M
4EuF9ICUtiRd9h9kzExOelbXj+p1SjffIbZvBKmSgvR95PACe5ihSYyMNWGMIhQp
I4SEGshM1oTEdAKKICQYaA47yZwbvVu2I514Za44mwh8H2Ql61wENz9jHwf2HSM9
7zDMmu9db9aNjSzDAGBZAeBxR2z+aUddgPf8OFYmqNwOxpGDa/Gn67vGG2/4mc+t
QTNzRgC7YqkHsZ3IC1xQ3MIntN6hyWn3DdEmU4GJ0mYm30FlqKVisV862Yo+D7Wv
6ED5vktMtKJXJrpbPnad0TON7enySmN0FKoR1UXPbzhzGqVfaQ1taSsSCeQkEpun
fO4r/dn3nCO61HbvLKocsYzmHyplRIjdTBAYu/sZvizEW7brcYsVIbF0HJ5KCjWb
NosZmLr7/XeiOgU0cTYouEodBMD+G0q03DZJAi3YsYaL5s2bXRsNMwjME2IJb/Gc
6NxGt9Zq4VrYOBbfbxM86uoYrR2CtM3wMXql+a4BClbr60n35kNKsC5bAgGT2BSJ
FgwpawF08FUJJHdFLjkUsVHCeu99Z3ltImSNQaS/pQxDHbAe2rsPGhn55mJwORnt
dVi+Z/t8g7918pXz4K/c+TYwjfD75D3vg0SN4rmDHVRdqLrgQOnOUo6TAzsIAsaH
WAwsBlh+QK5fuwVUAm8eGmSzYSIK9AYn7UmckMYxajXGkBdRNQyqUO/ACzvetAbC
OuISO5pgtqZPo4R7T7QQTabdvRtt5qcCfriEDLoQdzwFOd82kL+UaM1GhujMK+un
BlM0y9Zti9dMCeftibAooMbdsnNQ6oTuUmY8jtcbG1OJfOP7QYTS0KwcDElI8VsS
mnp9rPUjggXQv3je8B/zrQU9g8LZmTDzL2eNVNKpPvebK6CWLE2nMN9NuVC4FxxM
1qsMSYgY4ArkF/LL/fSPXy4J4yzW2sz2serSujokZ2PLUa2rGj583HqXTFGCS1Dj
tXbvlttWANsYGi15ILJlIt0cDrsmzWxx74c8peID2NttRoS3QMcSEkCZqJEj69Uc
NsZUmKKaySfsAacxqKeWcsV3ZYYKXyt6LZ2hKVHdVsRh5PPiyT3f3Keq8/Bnz7jF
FNtsg29+Xfw/eaARG9SWZTxi93sg8JL0m2cjMISSkQjVmvzH5wIVo2aoTDTjG0nk
2/pQ18HSie52LRv4meAhE5RFIiz0QDye96uPd0huD2UCxYBuxz9PPuoY4E+Ic55a
MRcMqMt9jCzDrYyhgobZx3Qs2xaylWbCaPA2mGqgjD4Cb19U/iNw583z3VU18EhQ
xlHfgNGArT+JWTvaXrnPBWE74nFpY20NCHhyXZ0wEI0BnFiqMKGAwqgAG63K76sB
PksYv3ZOFlSIteAV6tAPjkh+99o92ehWxWjgWNq9g4B3JljD8BiP5u07rMEg6hzX
W61+/7gEOu/KUlHM9ILoW/vcfE3bbUrXHdLFV+I/mw36Ck037lBI6x5BgTTF16hH
X5NZLvy5bM895BXDW1SkAPMEOqWj2pCnTPcGZt1c8rb1ugeF5a3zaWxwmnNzZshO
PvOg66zzAqurk1m9/hjUztknba3aO5/2Afs2v2dKAw+p2dz9Ep6zRYOr33pJDsCd
gDJA/K/FoYOJyw3UOCq2dIQBGtXTZkz80m5wCBlhs+/2UvA3SHn2DAYf2lMMNMhd
D8Dp28FLFq+ZEX0OS0iXEwlUc8FAi7viNKT7tI1DKkQmWDOWoObz1XQ8WrCHbHts
uz2DHmCpHtwi0BgpDAYIxUsveludeZbqrA84VlmWrWbYuz5a7Zte480ga7Oiy5he
Kn5kVJy59+mMq9jW9oD/2vsLNluVgJBhx0Mb7MuezDugUmlnJ0Sqg3bet9nG5C2Y
bPRspgbd08mLELH+uGZij7QdCf/QEPUvcNO+n6LBsSuvUAWCci2cSddOOGws7nKC
xHz1yczSqILSlsCPUfdqW9WAYyOEyprwPK2cCMu/7KHOfLM8/MbZhZJvUB3sO9ul
OZRYdT7XJ/VaI00nbV3ggTOms4HuaxwSkr/YeHYKlnSNwwBhAQY+IytJB3KCdyGJ
Lo6yp5WyA9zpZCf1atVGMvBBgueX+gzZPTLAc4+EgTpDR4JFZFPpnCDUY1Spl8Pb
uMmCI82Ga/j5pkpQTevssmFK51Ra7LlpiRq/VxnfzfqqRXaWqpy1Y1JgkdxMM/ip
M7QmJJNcnLYBzhOwNxFAalJX6UA9V2XMj6MuaQpOMtxDdQXjZW0Q9CGm0g/Qj3wP
yBBTTtFM7tXwUvr1jUMly/Fw3WvtmHHzfeR0newjIazvJrvUtOskGMMjperlQzFU
xVgjC8U03TgUsYE80I51MXklSbTw22EuQpt/V3qBhXrj8rowvAraRogW451mtkqv
BFPYoTYKdqoJxXo5NqPV4gCZh/yphZpJXT7gJQ+0RmDFZHqXh/MrlQtL++I5AB0a
JdrV3D/dsHHZOSmuaLT7Fr0PlvaIJ/5RBrGtZ8BBAWGBjPK3aSOTadskYaInmv2Y
PEquUZ8XHyHHDkxtfYTEQq0QzbwNVbtqD0V1tY1mL+D1sfY6GN4pCyWP2/RQ/rd2
+JGKcYtLqLWAuqXVUGMCrnLwIAN9L00VtlB4WGssCp4nrt73BUKp48kzBsprxVfR
tSSVh3df0p67rCzhtiOptTRCFUBEe8Ng+XBykAa7WwhwBGXaai8E2W6DFyQ6BBno
omDGzuKOZGV8Lw2jH0Upr2VUuc3eFJZU9xbWO5/fV3lalii9TYrL5P7pGKFY/hAF
PMe4+epBFfTxFhmwRRqobEjTyZ5j/Mzq/9xKmA1Q6a2vOpzuSEhE67ARbWjIhuWZ
KvtE9eOX9QzGPjWENbenYpDZlgpzvMWjW3yM3z1AHtVMfzaiZ1UUl4XpIt8pO4vO
zuhGWUfdzg9fX9CDSk5ADxeRjHUbdZX+baeg3HAiprbXwzgHy1mMboIUuDp86k8O
HvRB20cjS2XRS1A3EthCWR59TCEJVR8wCAGocbTwaN9Tbyc87UuJefwCcmD8SGmo
xMEhj9CLkRiBGf70bjK5MlfXmm3aVCoBBTT5IXGNCPrQPaICnLIZ6AmlhYTa433r
ZFHMSElV0y+HqpM20U12B14c72Sgb/nRDmdQU5rHnFjFc6wY15oeb3OIfLcG1Jq9
d9SEvWkUECyNQPo/xp5sN4ncACzknZrvrPUYJDCf7zEl1eMU1AxvQgzfhiiz8+2P
xH4Vrg+uYCcOAN9LTohtc1LBQCA3/03mpSlnzh51azJjnFWkef6Phv7naC5fUVZp
ZjMoUPB1JMH4hlttcg3qZfDBvHhUXgZeffMuW1PitVXxbiG/N4jx5Oy2P/AHwoYm
X9em14GwJfxZmlrpXe1WuAQNIX7CYJ27VjHAG16y3Yy2QIfXdiMTcN7adRnNo9Pl
L1ZRsEMjPKk7I7S69329kbFBhBrxZFirUQF2ytoyrART29gM2keOXBqathMWTZkH
hDicMxZZ5kfzt8RN7ZiboqHLNNHYgBI0sI51YLqZAjMt/OA/ZNTEpc42T4him1l/
IeK/965gCaB6QLHSEes3oZossbngPMlnpWw9AiCc+s8aTc/9lfqvKAEX00n4pZWd
Djt79QviJwJ35Th4lIyKMpX7BaM5pTXp1timg64PPNkBQ/sqgpFKSZJIWxKOY2nB
paAKDJMyp2xP65Mwr1/THoLVfFJboJkVFIuwRNdoAImJayzoR01bdWM7aiWECy4q
THGQDlJGdAbKoBjUo8zumhBdVHSikuyljeODjaf8La5Ef/lxSSm3jCfHgZxsdVG9
Fo/b2EaBpvL4VjmJr3+Ii6pPLp6Rr97Bdn0lvEr5BIZOhGpEJtfpthsglgFmEjEe
WjnsxTcrQ6fCbuILbf6EC7lzWXPlG6pXTK3GmRk4VNrvOn6slw9G6vI/22RvXsc/
ckb++GuJBBn3X+fGMzZgbxlRx3JnzeQo/mw4gAIUKHfrdmnbnsIMN8SQAHqkChtY
rxxgm1aCKfVAiD170QO/kBQV45dDIYqufteNdMVggHQVtuJDSzKFYnfM1QCQJJsc
VjDj5nZTlAQ6wZteKBKcw6qCn+Rq+CfJbFN8UvVz9nlklgben8iu/8DunFQhIOw8
kAPNhUaUDtwUGOhKiZI+HqU547L3FsR6/3CBvA8/2T1TAVay3ARO2cG6zQzbRcyc
vbNhnq337NMBlp2LJaQiI3pPnstCLiMHqIFDn8R0/1QZeN3xPmaJ8BcahwFYe6xr
y7BUNY1ZZjSqfFNvuSgiVgpWovoe3vj3R8i4B+6mY/yTzmxZy0U6STGFBuJcyEXv
fcMU6mAGJb9EMFT0AKuMDF/rpW+3K7Vc62N53zuCPGzzarlnuMVeyXK0RbcHljOb
8U0mnFVsJ93UQxYwhJKKlxfQRuKRnHSUllIPrqT+ZzLnDGd5Y90mrrgxcfLcmfVG
KTUknIVXrPlsvjU3k2JmlfzL2YzYZU48hkGNEKBs7hU6uBGnmxqSWpNBR8+Nm2PF
K/3VGWL/nEzC0wCNn0Jy9bPrg5AE7SAZ11kk7zokde386KM85ZLK7D59bTRCcd/r
PfHF6twVlaYx+XBtuc4ZSzy0KBX/fmPvUsTjNimKHS/24IbH9owDb12VBKNkFPm+
WUtsQ3l2Rs0Cv8iOlAm3vffvE2r7AyBFs+hD6puCnqdp22CQRioFI6IAhQut/De1
ndngCeen9iW76ypmw2vjtKMQ+IR6crPbGfSj+YXKQ1YZvUsgeLcxqfDAY+Df88w7
hOio2k1WLWkb7+MQLiqCPm8PJgEclWdjIU2OxE+elPLG15ylR44c/d/XUHX+JX8r
Zw4SSr4AVUCg4cDIBkCZkDi0WEpebaruIGdt7ueiNKkojR/XBWxkb3dEbze4motE
sl/ycjl2XwpxkUxIxtXuUhieW8GMD9wTa2wtw/1Yshk3Q7zP0vBA96TmBx8tSSDW
dCiWPB9k6wPmBTC5a76Hq+dUilYcpON/JAQsRJrtbPIQA9VCHsv9mm857Bl2lIfW
wY8LoICTQlRmAWh5PS3GuLFxjp9ps14bNiRJaNohiQ/j3WqR5kbeKFiq6gUltvPE
aSZvUYnZb717DzVRWcWUb+qU7UuX97Dztz5gdbKQXW5py3pcHckIFwA+O4Eo0E17
LFIGfQknLmx3FULFXlT3uzkqEYR7ZSb651CcBlKEwaEZcI60/rZjB3jgV50SNiIO
v8B4FBwcBWdT5dOKBZhhKIfV08mH5Z7Blx3QSKlaEiJl7Csb1p9XerY1/a0fxRQ+
Stvi78JuHx0Tb/kDHewO+BPGeQCTGCyGwSN6Vnruz+wVed5HIqiC3gvSLqMgVdJk
NhvDSVb7RttzNgy6fRpwnBbDJay6bNrgGCysvkAwITbA6NkQK2rM6ItdOsfou7J9
aukSSOB16THvN4X7URWKDB+2Ux1Yi9bS082UYdG9EU29usfXENmbUCiliaQ8C8Ni
aSQgd45hibrC9P85Shq9NY2o9uxj+QEgKdxpsX8LyFpIO/ed6NbM5tIj5avi3ct+
izmGyN23/cbsXEAzT35ir37GMioMjloGvsFndCWb8vVEHJlWeMG1T3ysNauSESpk
YyP/OdSmjy0KwwDugsjZkvnB8jGhkXiTKjGcDWdWDo0mRV7+mNbVIfEGLUeU0EvQ
ZPftoqRH0OUKJjuH61GgPm0NbZmJbds1DHaxbruElsPgETaQ/sTBMwYrj2SK8g60
DEkICbg/D4P+ATX8P9u5yLkq02wdLywZrxx/aEYXin49u9vax2UVcLn1W5Wa787L
3VyMd3NSMAOsBjVp8DaCMbFpbZ98GhO2CntLp1sXSNjV4XeCP8bAzourFn+/e5BS
4lljW0MTAWhUzJJxpPMpuI/N4JxZ/K4mOqB56hFsLminaiXHLJzBjB5p2ltOG2Y2
gl2Z7SidWRSUioNhasWF3JWcFT2l/oamxdlzYtnPEEegP82NdAI6R44Wg7aRvfh+
D5MpQDJX4NpdYiJONRYC0AaPjiflOYVKvP9JqKTzm0g+OPqfCY6ME80ysuwqfpdk
E9fG1jMCkgVjN4qpQ39i5e9TWaZTEBJ9txuMwOsdW/4omh/84WngMsSXjRb+gkVu
7WLwSORLvtgEQyyF+VMdPldwEEuOjKjWBdGlS/qaGvKtXxT8QK2IT/ziiMb0Px/S
KpyRA61xZT9YqNwtuHLiwMYCh+mF1zmm+1YPeqj6ZzqxtTIWHz7BCGPpUjG7v48r
eeH4VgcY4qbHo9jQ6roMc+XEgxvqJtZmytZjdHC4RjvajfL6+3pzUCqtYslrijWL
AY1V62q7K3wGeT+kwp41kPCM7z2dcrQh7tc4e49vf4omMZZCr6zaDmZ3BRaX6hJ6
rACKD+YpDD5YHfOBQuweq6LI4T5ljCPDkwJqQXMGjnxyzWG0J3xG5Oeb8V4cGkt3
Z3Wiz8DIYQPBvKODUZ/Cmo8ouWHPnmYfKS9sbiAuehVbObanG/u5cTjlZN79Ke+J
e/tjUzAT9uGRD6zaR9wu1ZAJZF4/KDNAjlCU2V/4cBSn7pF3R9Lnf09O801TZ7BS
qXLQWGMft5lULP9vGGyiImwjyzX5NUsqKQoDFjvMJtZrMzlPu2ZgYld0Ne/Ne/1a
nOIEemqplWQNIFBxCDOJsOkDFnafQvC+w9Kw4fQMYWK/7NMvLGDFMkuSvfQNNlrp
N1gkhlzSpXPEQwbUnZkyYAjf0RlsTZelC9kUvibT4UHTc3qOKIm+qpZdgXLUGwRA
AdGOU4iaNyj3XgsXnfpbYyx2XgJmWx656t+sDzcxUMMz4YhJvAsaYCy+k0lCDG5F
gbdC71wGZ8SWmRMsdNhLtG9cOpN8mdSC42hVJ0UruFHMLqoY8+JLN/UmxEF9r3Jk
DySdZBZDWaFeXv4P/2SN8eNsKiT8+5nIGNWqX3xIL2KD+gz/QebDip/s8RVVlnFx
FT+CqH04mxVUjVWaBKfMxA+QZ2JFBxlmwGYr57/hagyY4cVwXauMPRCzStbAjOeq
OHOGhCTisiMbtD/xXLNmARkEyInw13y9yFC7tUYRIk5Yqw0T59yx9w87/NxU2Kzt
CWEa0T5JNGuS8fW2QG2cNTRdCfgHStcW2gGZRgboaRRTYNXpb3fIbi8Ly25Gc5uC
gNxwaXcFJuwpV3OjyU/jQS1vRp1VKq03e9c55XTWAlOJCZFSReiL3/qrliBY85vZ
zAl/tIhCr+5SajAer/SiTt+Ib0+TW6qo0moUiGW5JMK+uxuTjQ08RIPF/8ye0owp
n9MvmTJPTLrCvWOGn/WJku53rDyxaX56jqX03lLbBLWKYJtS+XykhN2CoSRs3y7a
uc1MADchyxE0mjT3CBclgQ99BpkWSi6EUwlW0zXDyeZ9PYL7c+Al35M1A/q8t31Y
JVD+UH69ZEz2789KLGwlzLxwHIPyUeGU5IPark9HzFMfgDzfk5WBVVRKygUV2bPv
D3njQ6J5uQKizZC1+s27vm9do6b11Lm91pODMZFbWoNMGK3ZPsoua2Zzs+VBjsMC
jv0EwYVic2EwZxNwnInAu+2G2rgcurCFc9K0epxTY7iBayk3BCFhtyJwCwiLg/dc
fiC791poYI06Op4UiMgAUXQKTe3tlLSQe6aLWImxFYi5IZMDzQMDACNwWI1c49GP
CJ4gy/COl6n9eJmDV4hvA6BEA01uNwmlpYTt+RoIVCoEx/A4BnmhGjrhxeqJNDiQ
OtgWv2nHiswuxGp/bqYB7XySVbSlR6r1bgWD1oxiwLhWSYd85uHb2M3yL4Lg4yDT
1XRtoaANLhKVlKjeM4r6hPb3obLouWpmGK55LCulP3j6Pgnhfk/FASgG/fqJKKhE
zXk67VR3LyrFfRAyDeADiilcKrvahS6vguN4ZeYd6nd3HK46/nfxGu4+DvOBwgoP
bL3tfm8x5coLyOxJzcS5pEdgib8pTsddRZYAJ46t5Vfan+z0evSVKybeB4ck+sT5
1Y+ymSYi5fd+RuywSPUyX+IQzWGdm7Rv9i7eqJhSVBCrxb76sPy4B/MzO8aAtlQ1
I07Ub8chTIxvdIpdcD0AcnRgAnih8AEQ0PteO441gI3P9rt6SOwVZsHJitDuDC1f
jnl0AL3PXYJaobP47QOAjBafy4forotTcw9EsxSr5U3tz6MCsy8D3CZRNLQMw6j2
B4P9Ljr6jPsDdvmJoAXn2XhneqTaEHcgY6105W9Td9g0iaCkG+BYFStYKWF4q2ge
xGMJ+xd7jvsQH41cB6c9X++y4974Snpj9B24njB6ez8p32dPfQHmoRPn5yksbTXR
ni96UyPniE/5jd21ek8HYc1xHbm6wljO2Wr3Y0xPcnau6ZfN05vFcWuUYB4Jb4Ck
F42uwczuTvbvar8qGVeLerQ/zrwQDqYubvrxlFaOxOrMh3OZpk6g1hdsT1pNdBxh
ukeoxs85fG738Dk/H4gR6aZlYsg8Q/XXD/IfnbpLkY9iUFGfqa+H6ljXvNEO7MGj
BULUGJ3Xcw16MCf5BzPogqf+tU9cIZTd1xD2De24eNnlUyWxCchOOC9y25R1qtM7
ost2b5UwElsC+sPTELSQOvPQOw/Bx+zuXCFBtOtriJ6yKl+jH6Kv5c0TYRDBGO/z
gTX9uX6ymtkc4+fG9M3+mXwbzK4llFSK0IkLoUJLODJqttKCt8P7vKM2Keln+Zsn
Em7+Lw1+8U49hJEgJCwBdgP4MOB22gcENzkDEZbnFG6CdMxaD8cnpqQjsxekfYcg
271nyuweYMYamcj3hek8sOxeqRJnhnIfSwNk8P0DKw3RyfnvJyZxvW0zCVYQc8k2
D61ucsYPos29bQguEhjqBPJNKBcSYEH1hHgGx4kJ+LlVDAuSVfu5uY9CHeE1OTzt
p8BphlHuePcsac8EN2i7mKIKIjX1Ms+NxDiS/SlPr7KqOnCHlxvD9UAs8zhIae8c
JyxCvfoYxmodPgwaA13x85eWxYIExzr0ZruYHVzkO9Pzwl+3CAlwJVHAIxnXjBre
pXjNIJPcydPw/XIuOSEY87jBcD8rEbDn3nYRFFHe9lpWTz6aZVo13xNjJT/tc5an
EVw5EhfGDS8HrD3FOTbT/O0cQo9xAyPLh6zJ5VDOYk5JAGmiHJ59RJRpQGnov6uN
LhSkNt5vchZdnLqF8HuwXZG8GiqPe5joBY6YKl7cKkg04X/fYBLsmSjE68pNYvQx
7+tI8kBibWW6asyqygGZWpRSlgv0OAGvYoMbIRzb9GJOPJ0aS3NeslFBIHOdEN9j
oZ4PPyPYxL3a77mCXjFirRZYHdX5fTKVWZB1p6udnbz6FTJxVmlDZriT+5NAfCTx
kEdM+K0E2pLYdhtGeaJDGU2mpGDiZRn7sY4C+EU4/aBUGQ13gNzDQhVwouExjrtk
wysz2/TX2zzpwx265jOjbRxqIOma/Ws5JNfIovEphQFm/cHGN/7XxFOE8nnAjC9X
Mffc0nQHAund9jH06AaKSRGflu9X+LmlGqA85mVo8dxJK4COalN1KtnhBj+JaD7b
1CoSEqYuunbe4h4+DvbWwLu8vfseTzkydmJvaCVqBe6oMtEasIC4jsmfTpNw+ubA
Jy7SVCWyIso4V45dAJ8fiaGivxzVlGZjjM8T9S0TKUTKKyEieCQNXl/ic7HgLlT5
iW/vWGUrvaDNNWZMKDG3oG689e/kwMmlJwSNKqPcrJZNps/SPxM5OUxGP7oCGrxE
PzXcdp0mc3agzuIegB0NbmrrUWBHXFMRILKRQsu9o7KGTD7n6rXDxmmY6/QoVNpB
PubMbuFwSMrBHA/QUS6Y8vvaOCZ/Z9wOptGs7s+JihYy0soinRIHh7OxAkCW6ANJ
+89aOwQTrNA6MhsY331xqjidERJQaq4xy0VxUR/iaKav2WXhgQc8fY86IHBtaavK
oRgpLNyJHVIVCj3P1DAmIXvoGFVOhCVa4YW/AfcnbkvLFgc8eu42LnOKZf1Spp/U
C6qo4fd8nN5ZeGc00P7303+mxKr78VFJ8A6swZugxybP/fsaVcxMzXg7xpSSzUkK
yZZNglcivuRTE4oxQoFzIXUuZ6fvKI0aA1qDf0HAcxg8spdcZwTERfgYrWVzgyMc
1CuLbs/fY4XPm1/toedU6a2BznaSZqOnbz/SiaTINdqZhX5uJp+7M9gram9Riysu
KPHHRCc3UIYgFulokukFCz2Wx3GHoiCP2LpALsxPutMoG/pXPLU6svGbaJkF7E95
LXpm4rqtRzVIEjESdROstw94e42zm+Xqw7GZha5xl26SfrmXzGhHC6e3Hj1MCFvP
IViX85FPibNsZCOzUAQ5UzQ1j76oq5Tj7SjwXADJKuFsSkl66XbLIT+U2CNI8DED
yI/wVga2mE+R4KTSTG7L97D11rSKbmermLQ2ngbp7rwMKwjGp2Hk9IEYQu6QOb0c
29iN7OlS1yJquTssEk3WQyJ8/LnV61S3l4fg+naADofXUOllYxTTxDIzpu9H4DCd
P+VcDnZHOcxbM0QAvFOCEq8hFGAkVo2ojcGesQND/WiUuMr1oJm3Zu9ZXa+0cnFn
2nT3/Uwdt7TOuyqRGgSxBKtrG5XOF668mXuzyCt44i8YigJvR+r7qQXBzGlTzr1H
zkWwVUqEnsA8SVmuIJg4m+kATdMFUqbDEwYi4NRkV+FDTXV5ZMevLKPkfm44naoh
DsXkwldTna59aYs/mQhDHS0LsHit5eD7Kf7F14AUJZZ7jptFSRzRg5S7EAu9Zx/M
tjbebDmtR9P4QzTFeQARTGhjXQihYkk5VvxU4YTvidPaMRNLAhXKAuUUF/ZFHEjG
3E0TfJnKR6SLfx5w9F7ckAS0qPo9ShCjvQ+KWhWFJTRgF+FghJH4hW5O3Via0GRb
3KIZEBCVOH1mI2EP6euC0Fw6jUqFwhTk1P2TILnV5A9EIp09tks4yF6Qk1WxIOHx
RG8pVO9agUtJHlHpZwXMOvS/Y+QSQJKlqrDbA5dGl6rIhk2aWT0B6VxKkCQ00AsT
0P4UCQp/mPotMtaNEzCTJTAR3xCvYFsz0qMlEtIZPd0Tr9J8x8arLgouPdL9/h99
ysIUwbKST7AcElAFHlerb2f6iN26BiOnV0y9DR9AMhGLZ7Q+bZQd4PAPxUc+o3JL
gPxNhAtgcUSj+en4PJU8QVS9KWfEmVt1fHJmwfVaB5oHx46vatE0PEQgwH0rT1ZO
EtqixnDqdc4ZztI+HVuz94pr7Qq9x0KBZZ91cLPKY83CMxvDpa/OiclyFirqfYOh
V4swLo++69i8cs9P5FTxEM7lzGdoMjEC+qXJkXfzRjAISkYIHRTSSN6rd8Ky3NY3
aueH5RnoZnBnop0guAxVu+hOr6VKLRIJai2+/tQaR88q/LbLbhF/4Xl1DbPQD/wu
Tk1mUIPR3gm+/sGHUk3n6OeJv1zr3sR44nWjvtMbKOfp9AfkhuAAOFWqUvLxukF5
UQRfaIhobJkzTKw9LaevrBpkUS82REPCWcW1uLUT3LD0NW7xwXliv6r/PNvIAEHq
yRAenC1B3F9evZbXgkz1KtfrVLZfhjfQmOeIzrxJ6ZK7xaw1hJ+DqptYczRofZ2c
+/5MxUFwXyLCadrNgDExNBBnODM+qHCg+YaJKghc1t6KodT5Y5LW/TvJeXsAQRs0
e+/s85FBEvIF4dwup3l0HyV6hi1sHETxK1stvn2CEkY3yMdku1coihxdLuSEIgZo
MG4bDa5KYZ2i/4P2w2kBfLAWcGWQAe6+emx8LoblDxyUC+KOKJ2Bjn9EqRdJG+Yh
KKVIjkeLqYcubHLcka7piVSA/xwTVcBaGq4d2q10ZEzTGs1a873UACyPAge4nTej
LeeKPBoO1qoL2l4OFAELRHElF/FbZtqXXY94uxbfh3GhoOUYFHqktN5iywyqtdg0
Xb/Qpt+Ma9pko7U84DuBoWPUsW2eAZsI+lyVq5L/RXdHRqQJ1bDti4XvQTyVsS5q
OO+px8UBYDSQHOsoHZamNGdBmSbrEkRCpLcAdFt1EJ2z8G/iP3g/S/IMaL5L4/n5
PteVvkOyaaAKdJbHgVLb6z+qNw5IpblBZOLGje8orwtO6bSkRYDheONVekBSXSqe
2f9n2K6L6l2Uj4hB60qE4sTO28ku9z4b/Zp4fueDI/ki/BQN+Jc/KVvfjpsYAgt5
yak7zF7WZe5tXW9LOxx0W6hdIho+/XlXIiunSmpOr+lCl/uj2DuhRALGI/TIlodo
pG7Mj+ve4QBUYmAoxXDrhxAJQiubUcrJGkjf06XWNi6bpFXrSLmS72f2CsEusgR4
4Kmhdg8kuuYXZRi4T6iLPigSfvMHHQiUnkH6iTVo2Z0M3s/9TO2c+0+o6xtj+0Sg
HXLwY8lrWkQUp3wcwUABKSzA7G/ifKB53kseypfyjcow4YGr0PIq6QbpW05ZATp9
cBH59ip7yBCXJqfSKsKaayAJ0HWmA2wbtPm/VF7MZU7oli51F4tKwZlXtOA4Eb6G
+zPeaceCsJyCS5QAQr7+3Abq214yN5SwPkxamCpftHXw5YPEvhzAbx/xDrrXhvhZ
50qU/rlZRDR1e6mqaxyiMLiGqt0gXajiJM4K7zmPIsY24J9yqonF4LXl+pP7GqxY
cH1zzZtA1GewXcMaybJXwpL/6exKPr+2Fs7MnVNjpiKo6jHbrwWdJLVhHh4a8HUN
j7kUyyaTTWnejADvncMEur97BdeGsDR7YzNnvQ8KXZa0Z6ISzZCc/MtZDM3IYX22
9vlv/0G8v/FxgN1GW+48cJSJTWpRFYRJTs8NCMNkoyuzY2TiQjdanmoaoAo2B3NG
d1/a2ayk6aAniKfP+f+Ozj+N6Za7ZecYNqe9AM79YCzMRrn3xteG8/wgtbUMMMQo
lxlQQf+YGBh49t9WWoQ26IRnFKUHlhgo/Cs8LwHM8rsZHlTwMsu+MamMJGU/I2Qz
i92u6ORXHlCgssDJTjSUzNQzOaktdf3cwQq+9puWwOBcaHdrhl/bpm155Xu/hEwF
RCL9Y4ZdiVGo1BDXNbxCATasSlBVNphs2Ed20bjE0rULpdpvbgRbFZfATZ1V7cj9
bqgiCKO2oF3D9s+PIaBfijawn98qmLA+nkC184w5kh1wvvPfSenG1vT0/6Bk89M3
CklfmDYaTh8MG7yuGZ5WcMI492/ZaBW3i0ba/m9WvtkrSLdXZk+iyRuVY4a9Us/6
X0FPz3o9IhWu7gYQ5JaJusGfokhu81he4ZUeGasVhfmN8X77MlXJZNOyDwLxTsL3
2hXW8cPfAAZP379RsfshA8KIRHZfO3MIsdy5iIuAZhnyDjkxxnZcZ7TC1+Kx9cWo
oZeuPT3biYWhPfIsX4M68J/GB6LP9u3r6VdeWx6h9te1cyWylPFSiEdCRweylOAO
VsqUDY+KUTYNtH97x+Ax9nDTZG0+ZIaWZvuGenRkOX4e3Nthe5gHI0bKXIWEA7Vh
QIse0f8MkZcFv3UBaVQmCAFdFuQnVZvuJJsPl+oYpaUXqRlwbz7fCTZjqhgd2XbZ
He5SexfloaR6gmAXMcKL+wjFqrmRRuksurOeZ1IHzDOsYwtdE8vcSBrrfTLqmAW1
4tbpMhQUOC+5xKunBG5YN3TcacnRK24rEDh2u3ILdK4DJbVUjC5pRZTZ48rRPW+V
B5s/vHGjxnezJdZipHktgbU3twkFL3NXy3iz2RD+qPrrZjeM6CN69D7Kcfs/lJ1e
QRQawzaWRzwdimDoPL8JLbRcgAARK4okWO0O89SOyfpE1P8vMOIO6NaUw6vsLGBs
ew3qFGhQLZZpmfwYsvJorDKUJ7Tv9Vx4R18mOVxR8aV9TXkPXiFMIIMi+2+iofMg
+o8NTafV1qY6irkQseVNXqBaaVefqc5Kn7r/BMNhd5AlUYQRBgDgHDyIFYuDnbCu
jcRnkuSSUE3JqlPmHSLraKXMqbfEeOoy5Rbr6fkxIwEedvmazdLLH3sgk0MYEvBV
yckxBpnkGzbltges+fDOnU96UthWAsL8I1oomEv/zwVSjw6qeTO/2SUd5usv7Rz0
CwBC58Di2fTrRLdxEgSXR1GLn0IXPKYkMmE6LojjQshkEZENneu5wyfBinJYG30j
kqu2It2iVggr5nrcilDiU/PKbFBVm/1gVlLdBNqw/yssaSxPSHIpBe0RtT5+x54G
yyYbUlk7bQRWcWCM/wO3Hrd6jhrGSpcH6tsXWk176ULrSswnBvsUtfY4wjtbrClS
tNJK7G0Hu/cj4brad56fQ+Qi+7qNVdVGrg29yQPIaUqR83aF8J1lszaye+gw03Tl
O1JrJwkjGtyi9EIiEORPugD/hfIX96PShW7HFNWs1zTpUsiwNOm43sBjSjHJQ/ac
EZ7StcdM9TFKmxqNrPBOyL3Fi/EGXOm24Nk+Mmkbwg+UOnsebJ6Ilah0xTpnth2S
XfarXII4OxpzHpyWqqEDTbXXDBga+x2obA5LsvRobFlXtOLmSid22HaBD22nbQIZ
i9wHaPZhT3ddHjXpfLu9dK2CcothhiRhRsJzt62DEdpaX4q5RwkPy8RHYkzy37Ao
iO3r/JOE3EOrmOyUYj9kjOhC1HEeOh/tr1iU3wF8idGmn1UjoLh/JwBche3X5AXH
5fozYRniLR3D6LHpyiDuDDiX8QGMLjsDjMGgiBve2SYApgcBj3PXhtVgMPnK3FVc
Ux8SwCv6RyzhRxL0Cq+zCqGINaozToCwSPz4fTQuNXBj4EDoWz7RK3E6lXN9oj4F
9xhiSu+F64Ai2B4H8cARPEY4Z3MnnPcuywXi+sJkwiK/zzNLOPpIH20a/NgxX5LA
t3hK31ZzrK8mb+7Jx9jUFTQYdvqN12kNktHn4HmpvlgkwSihzg+bAy9uO1k/3Wwk
776kMCo8vUG8m5howKDFMLgXoRzOWMC2N5QwV2HnQD8SZRnLXkrYTLiyrgcwrowH
IdN1t/nRl4Ev11SYi9Cv2Kdd73Jvs1xLct3zQnbjUGFjX0RitnyDQk+Mdp7tuQ+L
IT7lQnFPcv6YDyGfrFoSf/5M/qFk0iBRsb78icB0pDmTR0R5MbeJ0zzVpVKv05u7
g+W8PzVeun//WDSK5jli8EpvgdXcY1tVrkvUaUhVN5UapvfkU952IyHxcxfC2uEG
ECj07qpyexDD7EP7i1+DNBApnuZEbPFqFO65pj4YmrwQTnmBjgfqmiUjZ50Dt+uG
JjKR+eeam0BVo4BTVL4ddGstpTGaC8KSQg3fkwwf/05auWEBdMSe/m4a3twaw3NE
Y5hEiO6DF8KXLb7JAOHDDKWjNE7S+XKAel5gGGqsNdr6y4RRnjsOY13WfgiblmO+
wEd5pXcUrJV/9BMbyGtnBxKspBISnRc0QSqUR8SIJQrKiYCOMwAZwxiFXRr/s7qX
theNoecC2J4Kptveg8SG+nPy9dkApmQ8aTyU+iSkY764D4Iz/ty1xKk6HPFKjunT
Ed2H9EQrYEfwYOMV82OXalnjBY6FClu7dYfQGziefyPrFDEb2mT9yu4f/McZxaxW
aQQAjice8ryvaykDMCydHWXInwzzC3XKisUGnvLnJAZxswvfa5GW3MBFEejiG+ZJ
mefMpW138msg6EW2dgbNqVikN9OeP+JBakAiuOq8AIFmtQSyTcpwDluKL6Gcz8If
axIQliK8EQ5K5DiKVqpNPyuaIB3+vqZ9FwiWaI4hQm0QpUxKKX2aIplKIWf8o1jz
Sk2zsLAeY2Ym9pig9uTefzV4DeF9J9irkSBF0Z6bwu31q+YtDjzxWH2I6EGFeyV0
UK3QrX0CxKxStYcANRt0ZdAvPN/+MuBbqCvjgal3Q/rA00o0Wn97spsFpikpE2MT
htIoMFhJYs6jCdIJaPMzJZuNAsQf0QEjTRBrKYml+/Jg86WjvNz7iMlWXluic4B1
m+ggzlFAuJ0FoWxX/vJuYnWcRsbWCVfcaWAEzq4AcqrPacpphhEgJXet1+QPtx02
10v5UPfoCvEONPOVmMF5/XCdRO1/CTP//ipTe3UFbfWUN2+XNnPZ0tPgveTyuTSw
cpZGRtXEQxgspQkkOSoJh5zJ+Nv39gCToheOCQcU73+j0GvRWnbjWnIOA2tj68bA
uGpVPHparLmTIZjXG3ycsLVlJQuaOFe/nBDb9DwrOqIo9NL6YNMINkrn62Wd/2dX
y7gRPMsDPh7gMt+6Qk/ooKOGZp9Cx2WervWYpGurvkSo000Q4Z1S1x/nKukK8RBH
obkCHFLHAvgCbEUeIWQJ2Ww8XrnGOtRGWYWMg6D23gJV7jGCNCi43NrnvOeXOKl8
OR57NAP/7PeXUcytLEPHfBaghlZBhD6NhEJZQ2MxQanU3IYBTK3XSMl/WoEi6ijR
pQmBr5TRPAQmNXzpvU1/+2IrXc0UJP8LogiEzd3+CeGlT8yJVVo42QXq5lsUQGI6
jLgusRmOJtlgMo2gWv/dCDb5oaEElhBJGmRYWv2Cp3zA6lPtoivZY2snz89ZZihS
KRROgjX5gAUQ5/fnInwm+3X2zdG2t6gG2Z6G8AlsAveqT7JHFJXBkjNcwcE1E+Bx
xmlckCVkL9XaCCXTR2uzWkXiB6lfG5Szasj8J+LqOJuBuP+U73IzHg2Qs3XE7o96
lTgZ7OM3vAZvjRcM37R9MgzGsCKtCR0iO6naKXQtMCJUt7V3juXlTfFaCHH2iuAp
o4DV5Bov1qAmuHuJ/43Sdz9r1iU/752cWvEy5nhtMT6nqOEH8yDJRr12f9dhL4zm
Q/Y/HP42osNfAaNIDiiLSmlTGeI8HLEwCRW6iosKEoc49TT6CEbCVxGraNQLuybE
atrNg70AQP1opNThGRHK0iN59w2SAXgAbHEq4WLH8w7VEViO36GWKuByuJDB+t3A
QN7sMPmGhad6Bd7hMgof+sDn3gp+h0lJ33FSOa7d7sjUOp5Fnkljk71MAZsjUhfK
Cpi/lqS57+guAxybwWQ9NoOnijmTk1UDoeViJFpB1OCDkaQT5yf+f7ydtWMI2hFs
RBpSev96IDL5UyLtE2s86NcbLJbzadAE7fCWPcKwwBQ9i86XifgZIj0mcntwU1Po
whUBaqWeHWHJOu2SlsOWa3rzW/ni5oc/+vbx0MChpwZqOX8rAxps7rhZtu4eEPZi
do03VQzQ/poCCnDw774wNg5flTOXNox488CYvtbbdN1x6OOJPsX2b0gYNTZFa80c
/eMOsp+8e/iGUwfysXEe4HrcloWAPgQC/NZDn6mghhuznBrqk8dSX4AJPvAQrffz
02cf4EZ059uAc6Fx36107H2OAUS7DYe8wLkL2elV8Gj0MoiRCf+QLsgvJD9cgYfd
65h3G0tVR5GHW57FEPz7hgR+RJev5SAjaJp2Y1qLG6Zhsdr2hy5Oyr8P4aY8ca+Y
hYlbETOQWPK9eWrr45YLB+f22pQTdwYWxj21tNStmd/SiYSgvJ6dlS1owbKqS0Wj
9l31FXrjKBZ6pS3rXRcy9BE5/UXCkKqgBcdyRfD/ffUJrLlV3+CmwcPF8qAcX0r8
MG5GiGZBx6IECMdyaCvN/1yQJEMo5qixYbbGFAfdKUhaqlN0UcT9c2MrTZbPpatH
eThlrr6i9BPdkDUrXE2EUhtO4hN/ZZ+Q62n6eGZMTmwD8dzWmmID0S0VDf6DsYzT
5GQzYewn2IwKHnC6QfRzyTNdxwI3iju934R42vQwCwObtk3PlHi/L2CYB+uapuWq
zZhbenrkhlnEX2qmoRak+uTUOAKLR1U/4dHoydku+C3DUH5TywEHIeMZFVMPK1Gr
DJfv9WDzJbtoImh8FIHZ70D5GcHyTQFtIj3CeWcTZqGv1R9CxiGcrUv4gL3QcJ5E
QzRh6bUGi2PV6LS0/kTdHwzRSkBfWB3YocedcsDhQs+UBBPlr1Mqjl5FgOKtFoMl
SNZ1aaiaWqFnAlyKl6OQAn252+vXnop9OgZewuDIl6QlKw2U2IiWSCYB+tZDUE4W
m/GtccjhJbtl7hQzR/fbSGRwDFJ9966ol3RAU+59UWgecd1GMsAcf40LOt05S2Tw
tn8oXWSgKSdvvRnrBJzGr/lGn/gHXuLPcNS8ULS0xvJl1YQvj/Bf9diSOj6I6ytv
VXcv4MMNgfjekCh/ZSDKVPcfOziXMkPM9s/SeKFaeVjH5eQMqs8PgnyIboVwA/Ps
weH6uanfLa7x3R2NyeeAAJtDOSIp7T+XVLTNYTAyux70F/1JT1q43W1tU6qFBFhL
OF2DHdWAdCUys9Lp6v8TY20i+JfGhilfgKqWTzRmC9VRgKk/pch5sG7Plsv5cUA4
wpaVWy40hxp/rIZx5IGzmzUMPlqiGxzL8Tbm3OmdPyMnkgc688Kv+IOGKDfGo7Ne
BVXA/aw8bJIjID+kicaM2dEGL97Uir/b+PefIS8mBceZl3P2YuO8q3/++sNgLiRY
31Poi7veaKYLa4WP8CzSZfEK/+KCH85gX6NGH8nFpnmanDEALkkCc3Ws4dmtreDL
VLqW63XpNB1lsdLJttnnj5tr6FumBh4zh/5QVsrgW3UWX2fsaP5EZzkjqssaV0XJ
9CWl1dmuHdk/swgn+tRijHVHzP5uq6MtZoR8gZMPaP2m3AxSvypkaFP1z/VCu8Wo
8cj0MwaWKnw0uVlImm1X/F6C005iWQpGlIhDjn8DCIiFFkcjKPxK+Ibmga/lZCUE
IticN2UriDSdDeF57qpr/o5dFb40KE91+ulIQmpmi6hOx9lMDWS6Aa/Ccybo8QmT
EXnBwFrgUSagx2H+TcS2vkXXvFu0psQK8XX0acWQ18MqS3uzMS7IlaBe9m7pMwcQ
62olOJHuqzgk9552hbsu9XlHb6ku42urfmVviPWtzK/hi3V/E8mP+vd3ys3T3f7Z
Ub3CEcUvAIxLt+agM+qATvzKhkE0Wkoqb8XIsfONnDwk2rbtcEATO0thE16a/8YE
ROX0TcvHhGwaeaomTkHDPlDBKoNBTuj4lrZRpmHAIIVCpqwE9ml6SkB/gfrfxguH
FAfkLbbmtRVZFcQc/cpTtNcy++OBKV8pCy2jTQz09odADyUJzTfCKq55GAcwPhky
MmUWUWcdSeb9QDc3JLtYCPXc4vVKrOZJzUKj6UQW2h3m4Y4u8djseYHmxgaCyVpz
nSBShDhOIthfY71YPPtFIR0H8q0zsiY9sGpGhfqRcMDRK0403FYZfS/rABIXcEnN
KvlODRvoIOAWpw+v48dhuSaNhfy0LB6csP0Jiz2Jsh7KAbFlNte/BLi5sfpXvprs
5MmAxjcNx6Jmfr3CSJNnSWahAOcA+OO+N272hDsQgaX6QOiTs/BoapiBKO0HaYCE
BDozNqu9dlP84HP8pZpZV0oOuT5BYn1kXmSUxd2pwQZxC8zXn6fVOcijLT6PhrPY
1CVcZMP5bej8KW1pUGiC0zjruyswAnqH1fZPPewOdY6nI+k7e4hf7SZgveZKVzGD
fypLjkEJQVPXriO4/TVa91uxSLoHZf5z1laNh+zyThf1hmzPvnLCLET5tAKBk7wk
+oWqACwwMlG/LHfryFLnPCzc0rE/dJcNrdQ2StNXMCRy4LmKkTG4lXg1c9yjcG2r
65w17vqV768nb2SrZDPafb/hLeYkrp880pCqY09hjZAuMqR0GBzE0ull+8yr9e+0
DOIp5S22HqLTBPn2q7LUjDNIQ3UDoVh9UCTnDQCwqxEbOtYCvHoz6q/fhlL30HC7
LpRVzxR7M2ZjiiX5PxpR/wXmBpSfqrOHSmSxb2Jz8t33307MNmI2giP3N1r4tRcm
pPjS+2bD2SdBMSgKZ74pHU3YTYrEhOsQHs+UzuZ+BjuRnIbFegiUSp74/JBErPXL
mTk6Z63+kTWoM2h5X/SFxpf9WeDCAdpM+k/cvAR+XBU4c9GZA3Cy8oZaw6amO/Kr
CRq1Gg8dceLfpjkDZlxy1DCwikApiDNq/mP9n9QbEkM8fjZsHIVxK4Gb9BR5O198
LiyZrmZgTBmRUaNO3DOwDJ8FYbvKAqXbRy0CkGKRbsxKdUhkcvHFd8snqDn5lS2H
nqprCWew1N5JIBk/mlKLl555leJi+Asf/VXxyDKYbJ/UUgdkUXzZvcaeWAoQWDyu
9VWFhS57HeFZBs8kf7Y3/xqmucgFD+RJmcaFm0bXyjAL2H+zL2kmfXwXtSNNmv/j
7mNEuzICTCck6HbU6cZej8uVE5xM4xyzTpdhDoUFIGtgCkkOi/CCPl/cix0E3G69
+q9RtiI6zYHlW4w7FVMsnFQXbzghxvRQ7yXZOBLKxGljCE3Whf/l7HxEi65v+VPO
nKwyzL0YAG8Z5ZKcp9O7I0FJHrpqNVYOWi3poqjSd37w4w96kNH8GdVcw2HBsPf4
GmQ0AhbzhW6YrJ1GXh35au8Ssaek6VMXZszzwvQB6PiCWp07k+sJESeFf5xjnyuw
p7Ht4pCT1Jk8aRjXYH3VcqazIITvsUFIGTLAHW1Egiex5zwd8XUpLA2rSsTdMKX0
hHa6Astb1nYVXL2uncMTGA/5LBQsJ9KoDpRCNS2lK5LSdLdM9MrtCHIMXQ8UHkU7
G70QPyLz30H3AAg1rC3y+JtWBHpgpE6bNLl2vr8SW60JPvDXXXI3eHvlXfW9uHMz
O6qpKPFRFML/Gc0XKS4nrXzgAmNL1r5wGGhopls6i+uxrBTWwqO/iGvTTVzUzOy0
vZqFihPzP1R9/5Gvph7ocNHQ5i0BEprRWUGebdYWM77L9yGHELJVT561JWcX+zOy
ShKecR8hZALCQmdQH90L0OZ6VzTlFcqYFYKbfZRchYoaOXI8zWY+A5UOmqQI/hA1
AwOS7gTy3qRU20dg2AemoxMd48tiPFAKSbDZMONqsUyf0fsVWs3Yr4pmIWSu0azT
qrOO0CPQqLSOlzCjbGNBgu3I6q9KWlCBRgpmTS9Sp0BFK56rRCy3s+rLdzffS4l2
CDT567SLBH7/5II8CJpClzA9ojcTgnYDkqPZJkkWyccpA5GgljU++7uEh/55Roam
mh2Kj/Onlzp371uWd5ICQjYjwVKjDogL/ch+oCSK3vnxqtpchz+dV6szHG7YVGmT
/CyhDjTRBXa9VMeK/AQrTkOYQDCCib9UzfYqecrqQHKf3Rbh4JcsUCvLicOsj7LD
bLRFPR0jzJo6/XDrROANK4tsvRSd9G6BN52pBWj9a9YQnKYR+M1nb3TvD0xNiKyj
hsKgTCzREjKH/YrGE8G6B6YBzDPeFima5zMS38IFO/RYdStzwZ7WZeRvjZgjo61Q
yeT9GAQoznRi/HAIH/UVHNiE+atIATmumgERYvDERkCVrPbQ3wSJ/f23yoYsISIw
5EyrpTXuq4hCoThFaA8t6vuamlM/5OkgpX2KLHyZ2ENlA05pFpXxTEo/t8lovUui
yhk/0qoUIHTLISfvxvXdPiNuGSonWcCqUnvAPvKBNSrwgyaoztqsGsqNHwiej2Sl
G6oHrXeByfKwY/LK9gtsZBndrFadVy1H0WFs11VkNQIfa9L1XvRH8FAvyxPI+Ne8
CRRjB+A3HFGTAja/bV9AfwyqB2Ex3Xwpx4wEG0eZVMHhlN8MZNtEM4v0SdJBoxz+
64kfrrcMwL14XOnYQTeM/QrFbJDAp3jhPH4Hva7DXyye32U6DJuXDOiqZJyjWJrI
vXUJw2vwgmejbdrqgBLKwyhjC8/I5C5YAzIdhdF5CcYy5aIo4mgu+zvCYuqd4/ZK
XrPL26gaqC8ABsK2zUNJq2x3zOg/3d0cT/+nKHy+rB2VOLvDctAB8izFuNGrADnh
gS9mL9Eh76E3KOBumoytMOTrP6JVzdOAdhso2FgCQ70ySwrVAWjgtVUcLG34LRB0
cAoICWTr0ftcuaBM91SsdcqTzy9TEfFXf2hsUcXjyTMIFrL7oRILGTBy3uwHF08a
x05dds8rWIip8wxEXYmXY9SA476Ur0/u/1jhkHEwlwn5aBPprKIBbYtYimcTI3+I
KqAkF9N4sou5RngLoTSwH1Oig+kxWPM5xpqkTdhq5U6wbUNPI5BFLKqGtVJbhfy3
G0L5Yv6Wotf5hdP1q1fABmNWBuUxhKkL0DUS+lf5gXgVV6jeYAgdoTPezRPCa/PN
GKatMDjzNZX//YvQocvycCyyds6IBlyJM1zPMlQqZurEgNGux0s2pI47ioda4od6
BIKTaQATz9wgkBDGHylRam/TPzWFIbyR3y/s/owANW789NgWyLKhFIi5/uatPqVw
rNn4QOePvqHy7lB5N9MmxEzRp5708MDIZTp9QhBN9aDFLjlEblBjh5HiPwtjBgKC
YTFoGsiQ1r7OIobpbZO/sPbf1NYn4mK5PsVbV+XPU8yRqXTs/REOeSIZVv17RQnz
tDZ868RsOovPsL72o3lqPd1zpiqpiCh+WFtVZLEPfTNXa8UiglbeyEE7FOJAx92/
4Sff5p58UbySdNN4ctj53cNfipmeAQ2dadlTNZOj3xX8MdgU1x9DmpVyhFtN6rC5
CnyV05YavgquItgSdaCEen9FHhMYtXLcddPc75xYZIlNt0rapto/ZNnhKrOwV+qs
EGdr/dG+6ft+C6cAqs+e24BuQFwKZvZRkCpUg6b015iT+LaxVCltp7rWyHOtM1Jd
7UrwGifd5Bu2OY5whG52qSMOQJ90Jis8ou8T8lCMday41iwlmFxAYyGY9JQbfrwj
IhwzLH63vfYBsDDtglSJP/iePPXbMklQpoLN+f89hh7D7Uvy93Pe+KGXSWhUA6vj
a5Xb8gdFeSXFeSYToey7+kumvcFWNrXOzvxB9yqrilG46gvBmrg6NTWXppfE/d70
GDl3W6sLaiJAqLz5Hv8RGDkKURR9ZPNom36qFcFZFpYuonfWWsgiPDtxMUNMtO7m
ckoFUHqQVaBPedy8m0pw9bonb1GiC/g+y7ci2DfYura9CFeGAmCmj7coFrxRJ78C
1uRiBiizyUoEHgOMm7BvnsBwSHeP15tRCwQrQpFwv5o/T/4T0l4fG4b8YM/TdCgD
JaxNuXYS/blualoOJn71KfuDvVJLJpXLiz+dIB1T8nBpe8yP9tdJDf26Tuwml6tc
HF4KGj6Y+BsqHSBB6v/ACeZ4byYf1r7LX3x3ftIBbXiVf39gDgL52ckPtoPFLtJk
Ic1l7fCuuS6T/LKKgKAuAIcZalofNtnqQpp/pMiPsdfP/4bCW0ZYYNnsL/2Bx03q
1dCQTn7JakHdB4gPX4q2S/sy5lAuw/shejv6AwsqeDcdCr103UJpzmsBDEUVy6il
94DwixlwXnsbCF44gYeWbMl+v2uUVnSwkur5GgdFCL99fnf/NkU2hIaX/5DJZJ5J
PXRQ+9M3ZFSYILlDS6NYmQ19hd1/N4H90o1TUHyhqpwDdGixA1/DiYu6klOa++6v
w8LLCMKMcjBbSfuAGjbv22isCWAwCph3zW3u5Xmo+Iwn+Y5hpL92CfTjeYYH7mlV
B1TbHv8ixmIJMsYtF0dTeVs2l/fkJQEfJe7Jo0rt27tWmNfQlSM0WXl0Bc9c0bF4
aCqTGaxLAXHbHF7F20MIWPXuyTwZbM9V/C15WHYBI/4Zr/Gy791wSiN7uGv2/swp
O5Mgu6B9OveZ6yFvVNtXEogUjXsnCHRg+QRtGtYfypNeAgdEwnpfv6ThzYCoMFWY
CJXP0xLsZvkm1+9CwKvqLXffWZHfsoMUQzFCc6Esd+KRi6Cgu1EWzVxbbblG8tWb
geTjxx7CKyoXb2sM0b5XE6ydTYENCrcSjN/pnK3KAZJ90uG1WEZIP6Ig4/EaXVMJ
oHOpyuiie9DXvMiJfykE2QVaXocTeGBqX5rXFQNzJDkbsX9cW9X+X4/Ar/bGm5PC
J84Q9sN+qwMlDVxKL9GoeISOKjJ+/x/5mYKc5Ak4AEU0fuSxYbPFWjHTyGT1ZHMf
2YcuSws0twlmLjTjbVVuPHr1UPq7f7AJm+FdI0dHA3Sutvxds2CFF9rjKPX4GInh
bD7iAZ/L/TyUimSE6o4Gnv1f/90VBGFWwZg2+vhvA3CAcPhbt3lHcvwITePn0Cs2
JPxZzDC8jkHzSTYHJNBFbkbJWNlpWz26K7aVxmFrENQ/pyy2qCkbGtXhWcGDfBOo
dIFptHyxDdgWSuAMrsk417EuHQlFVQpYQ3kB2HK4Ek/NDEqvf0ub6xUTybCCP+4X
7SILiPB2u4krgeERy/oP0GCbPp5JdrL5reNPfC4hTwVk2Y5StXL1tQiKpp+QhqNn
hIDng8UrcFTEpYAiMuvXEW70oTYJCSFsu74Dx/vS1Tu6mMMaaQTSDeEXZr4C/WMi
+q2wX3bbaqrimDFZqYqq8d0801AUbdO5kf1J7nl+sNl0tmImI0I16h00ISxuN46o
oRyc5WDeOzh+pdG632RP2rgXIy4RFvATU1HNovnRfP5jZYnreX8WE5RXgKrm01to
VYFPBI5FOuq/xlUFQkpd36BvD6RzXS/xWJ4VFizZWckapqRgOUO3FK9EErgISRtd
zD9Pq2+yWTJH4S3qf4K5Ttaf5woAtARvM5NE7mfUWugq9Xd6x20nDl5HwzS4SCri
ydlmFWPFRQmlXfJqxmuq8GdNEtvZnN4HsARhyj9y1NicmwkHYguhSD7pirDeVgIS
ipNNkBi2qNd0dlJGBOFLTQAJLAimhu0SzBknWURODUceBlKYeZUFsBfngONzFoob
mpio6AHc/3ogxP1Y53mp5L/YNXfVwybl0r22rbLGTrvsP8dBdMfH+HY+8NjzrtZ8
L9afHk/jf7lg1MT1tsBNRFF3HKkptP8fJ6X22ZNuTE8FdUwIUFgHCg6LSlxySWEV
UsYWp6vc0V+StywzK5NzlhZ5iHXTwpb0UVRN3BdGDuNigX7/ksR8/8HlmFTjZywo
at8SUQKVhlPA5hBPMPIO1dNpq8BVSdj65LiirTinj4Svy0PEUb4TSlT4VknowIcO
kHhMFTC2r+ri/9jov3vQYobA/cmKmX2xzyGKMjBPQBA3VAU34/Wd+MqLkk96H/2F
rtdRo9vABRn8N4AvNbS8VWqxnPJvStxCkCU7wV+IQRIkOFd7hGsYyEAhVBnvagyZ
LgTqcZhwLL5N1Y54QzOf9m6v7XcWVIIVYuLeTYzTtfMAgBi2hJp9V3zEBFc0102v
XhLexc/+bnGkE6YT/2RN9G8Dw/gxTh6LfnqaUjllXlMBXdmEmfbzbyjF0D0ceLCk
S7FkfanL5eK3FEUkOR7U0WObRu4rpXUWsZWPylJlNjU/hA7g1YxQjtFmgMUPS7OI
Hew0LVwyvLcAfCPSjt83cCHQbIQeNPottMl7jaNE6FqxEHbDBh2YiWiDtowFbL2p
TjQ3r0gxMQgGps2qiGGjfboptKpomaSo7+MjRzBlqMkJZNMKXrKhKn+YIX+njxia
f53RXf0OmrTOARqwGPOI880fCUUG0MrkIB2Cz4syT2HJW8Tudp+DDYfU+dXTE6qp
jzUYugmh7fDX8lS5FGrQkDfzI5xXAmLhYtWkNlKPr+OpR1bDHgyMw5NH677nmY92
peqSd5V5J8j6LxB3lHqCJ5VRqk89NlnsjcwkQeHP1cg+L6aFHX3zUASVOd4nv3gI
K2Pjwy6hGHngoafrFgkcZBesU9/d1rsQM2Zv0zr8GO0bjLD7x8IDCpO+psBgFyRz
TpljL1UTYsVpmWYVHBXkBfQ4BLNSiOLfbA4QUidtuwjOn8AazwRy799PGacnaz+6
gnPuNzxBy1INGlbdFvpmRfVTb4m5hk4nXfVpk8RolFuK+PxquetnnFVgftc6uYB9
SpF3v/XZ0d8x+fjgUMRvCmLyy/ua4uAJf0s55fNrKfyydSI4d8hvftEXHHjlR7x5
YQT+2eIsVKtYowp6Q+uJ6zQk4Bg7hXalwa4cFbEada3N7wHtAx4AcssnqUKRN/qy
4blvl5C85jpGavNNxn5fkQTXEcWNpT+geI+bSMhMTKZHA70h/9SFoOnAxRz0JTSC
m0MVcGBjpGaBDb7s9zrIYClmXI4mQT73ICMMkGdxXBIaj6noK+wWf8BUF6Se8tgB
+l0XTLV+TESGbvNRktve1ijjEjNihniZycf9Bf81hBndPi5eHhI3A+n075popcH5
leyka1unxfKgw2ucBTXyBFRnf6TXewTdzOML1MKUZ8z0VDTxGlyd67Bl7Yvg0U0j
3vpdvMR/Bt1DRnE92ccClT3ekml3D1/ETwp2xw37/cyafQKoaZ2+LuF9iufrqCtU
hwFptH7J1DuvTj9Pc4chuQ1W1EmdIa6D9tZzPKPi/vQo6bG9UBbufzzAC/Su4uhJ
Nvgoar3gMBrq3xgFsFD3nMErDUszv3z2z5vLQoD1r34n1gUEGnJsWv7jRLLbkCup
SEVY361I+LpL69RnCfx9S40/Gtt0YvRvvHSAyjj52c3tDsiGIbWbDF92PcZLb1dr
ElseK3RV8AZsCmfm1X1q82+3mIOH5yCcHHgDqcgZrmoZm2NHdn3bzQxCSN+qvjah
cGEmBY7DDqVymMSHPfJUe9aKqs0i7OqvqGwWZCYuA6rdeJtlJzCPe5SFVPRW3O7x
Rv+LbJS3Kt/FyKtrX5ZrOlLqomHQd7T/O2gCvjAoQyO00/qgtiET0AxDMyGQRUu3
yCP9e0Y83H4PxyeMkZxDmiTsYva0WqJ7Da2acJCzlY1//ngTaBUWUIrNfR6WSfjU
9SVoihnF73EEuoiI4eljfbmCtL5hlPU4RWDoQwOxSWfkzuVEQkW2DYFBuAEOARFR
06dUnu3RzYUiOaXaObKLsAPPDlUoXBCEk8ikAi1l62ZWU79UWoITX2ItjJnQMabS
oNnqF8y9tSs9/VyaN5r8FaytwjgSLX+S7/d7s99iWCSLyqd8v91cOPP9YGxvgpaj
oIhm58zlUIrx9yd392ldKujHhtUSPW3SxIU/2JRUaCyhQSysV/QvQ1grkiF4+tk1
IDRIyLME+xHnGelb0mdDz6EItyLg0nobfxyFaC/S1H0H8yUIlKMCi4mK3YyDPDQS
1yznOXrmsoMj3CcUs6nWhJfGYty7zMJBedkLt/RL4AtuCWcSYOwkDqEOL0mqW4qm
uM1fLaSNPJ/2QaMvMck+l1tudXQKcUgts3K5VX7rhDf8aNZL4639IT3ebe+DhD0C
jDarFMQruTuUMeF5BMyEGfWo53HEFca4Qi8DRupvdNus1BuWM/nWcQQko8bBUwQL
9BAQnOQ0LBcBnfvtspQV22XY8CO9dAOn98JKR8uEgNl5yRk1sktWVYzEp20PLbjD
lhw7e6swpqpU7l7TheG5m0X2U/vXGg2hohRQrSZrcQ1RsLeoZpyxDeCaAL8a52PZ
eNx/zXRWOR5GT9ISkccq/qdoe4v9wn25Vuyl19Vr6viZ42U5KloEdCyPjWzcw7Lt
xOro9RSvQykFOHl6TlpHTbcnYpnDgqycIjd+qXwUct2B+VkCBtjwoeUGk9mj+lM9
oqRkP5RM3nIGNvgQbPm3IfnrL0QdDXmuu7tG8lEkliT4gJueUdDg2ScjPJ6muePa
v6YW+/Iap2txC1PzLuaTpNSPINEpkuugwDusBdoxWU3EfYpxggaz+qPzTz2Xieem
A3jVqVSOpWeo913NtHCPf4DvK6IqfZpBywXAa156QQi5+/DV47Jvja2L/jPiUFj+
mDBC2cSikPvlCSGrDT0mzjaoIuMx2w5HKY12IHHoOx5h/B8Ej0t5DnBlXggfFT6J
tINJ/flyFedQaA2NybVprAoiImC+xqOIcZfzKOWhQiCBxJDRQ2aeGeVOYg357gaA
ZHQImlar+LFofjiIgJYIt/2hma7JwEr4+iZU1m8VOfwOx7S2qLZqgsHyhRMksWpM
DYeGj8HrzoGgyYN+avTRAuL2SmwOcRLM8TNlEto1ORAs8HNWDxthTti+Eg9vFAtF
qY1PL1ZIHf0LOHCrQEkvznoawcYPpYnLnhe0iM7jwqVd5yWwfPvAikflY4K53kZf
vSuSQgdPdC5VpDS1FrBeyHPnMwuPrJi4OCGR4iY+PXkHmQDidxZA+q04lSS5ca+Z
iQl0njugHEwZiNpRB1cY+9oXbnCy7OcqNe7Wsx9o9B0L56gTMauhzJ7OBikajYzp
82MVnHByl2ArUu42o0hL6JSyiRkW0GpTMZLgo3V+s9vGoA5N18l+xTRlQPotufR7
Usw1WK8btRirRoRs1T+1xEtMELTbVYElJdfzIj8+7Ent0mRWtzRX6LpF4ipNoUX7
xaxyIn1lE2NHV0F+vjT9vhEExbSDl0Ybwj3onXU8O1mDyUFQcKywWkrU0pPTxzil
7/caoaJlViKxMPoVEQPBzDRGtfbpEYWNG5pcqLgu0UmshEAJQZhTZRbbRAIWRBVw
xQArtm2Lm4b9+K0yYmfI1hU0pP/ZSsedTPEfGoP3fgRUR+HipR7uyZOW2oUHyhJY
kd/RoUrji6rE5tjxR3HjxmOtLvECsZEBTmbGsRicyHoZAIi/zvNQ/0QAWSNoqdqi
GI2w32wxblWS+ifhjxSLrXivTZ5EI4Y/O4Jc/i99iI+LEq25qknj2Xm/ut5nktyR
Qi1mbihjJNaGH2cQ0KV89NujKFuljFGOHb3FC7kvbdzYpxaS7QubRr6jIxmuBEfO
uoeQIUCV5HmmCoIZiotBLmdEpGnhXe6qaczQ0szK6wa4lK8BGLyHkG9e6RLb6uON
FghA8Q4quCoOBD5Ce1ClNX8NbGgez+rqKDhOKZnZV0ODH2v9BY7YzJm7GPDqgaHN
hvkWoBv4L/ShJP40+4/PNRPlsq9ipiS0WVaIEO4j4G9J0ZVS7q8tOZ8KxLFeXF22
YQ0LxulszsbmXZ+7L6EJT0FqzL/3V6mzQExaAjDd9z9lT1FtQSpZyb4G+Q5SOb7a
b71KC75VPv3Ca1pJ5qBI+nHtJGAjmazt5MUZu+7sQzqWCjtWHvvUDBnHiZq/VE74
9ddWPD540yd4+8UfvYZjWqBPJsaAY6nRUPO1bqFYB1eD0yErh8teIsHM88zpj+1j
r3kz0v4Chj/DFwbAa3X74zBE+LojKkFzxmwxtTOfX4ptlelZKmrB2PQfPEkVnBfM
F9tN+75yMXA+BzWhLmbGP9TvVwbh0LB5BqGO2Bx8FVFPbyZEF+juE04AnIO4ZZwQ
UateJTiGaxZSMNrpiikwV+9ne8aLZhnpsD/HmpgTLyGIFVR86wmvUcZq1LI4hk9v
L4JEtvonl+vxcNkwJfxczxOra30PkYTZR1OChUSA3wd/Hl+Gamx1eUnetRc6YWNN
ayQCY2XjtjN2EvsV4cCo8JaaUniIFkVCV4Wq0vaMXWcq+T8yujbeIAJkrrcU5w/t
H5K9CjZr991lIM6Pc7ROsmWGK5x/fNlOASBZBlevH4sksbYilEPQFJp2PYJ1jwFa
zANWWvDqH3U54ABMUvWE94cUKifkzOc99MYycngF/32NklAJFrf+Rnf62wyXpfLs
yHJIQZS1Yvh9CdlaBGL94tUvvS4MFBQAEbisU6rFNHU6xhzRPWR92nbfq7uikG13
EgTu5ms/Ht8EGEx0C7fvD2s2pW8tupT4tJmEQf3B6Tn6EBfaaXgLKKZF+LNS009Y
EP8/H5IhnzKIcyTjEBuXFJ2vtXyBRMmR0yUiAAJjwbzoguWwPjnD5ozoFBXCd8P/
PZZ3MBXhuP4vsnFBeECxAz8vdrjmnpBryjL4H9g972EDtAiY4Umg9qmUSjLO4NwS
QcLUqHvZGgZnIjrIZll22ol5Sl2/ajKPdFxLJutU38YUZcmuKGzBa8D4MvvE7ZlK
AEaJZ+UJAAsWeAUpQvNEC+KL/eJ7YgF6yj6w4KLMqJ0cIEOt2fIe0KvTYzH2PZxj
/vOp3458da1hAgRx/WKVseS6nBtMVGeuM02HYv1Q8GmVMjVvA13mGhEt4wQx5CRN
UnPc663X3mANGE0BQYV6NJ/Z/xDVgVs8keIxJ6TJvg6nYX9g2boIwPkK8ynzlmQw
X6+VTp8K1BJnZlxFtkX0nQ+U7JL6uGO2bCkWoHpJmMODf0Qtj+PeranYKKMkxVOV
2XXe8C9yqSpJ4mwDpdJLp3aLF+EkqVg+x8AlOKyQ3WDnP8KMhTk1x+7vukho3Jo0
ZZ3HWOC+E+lIICKQZJOJYwS7LVbYnOzZc2S3KV6QTr6LD1bARF7KnI9NdgDjHsv/
7pbIIwUTAiZ/Y5fjKxJbB7lpU7xBIOGNtoeh4svvADll68Iu2OInghUDY3MOD+GX
z4uZW3C9rFsv5pw6R8AJjlrIVpmN8rky6y8ze3hgqLgY5sG3JexmY6Yldik3T9if
FjhuPx55rG8zFOM+CUxgSmpZfc/189RWGYyLnH2nwVI1dHsrt6rIA1bk31DFtTQp
PGqniJ8US3O9hWVXB4PBkZpQ3GBF1Ple0Sxas0lxiVBrpNmKybFebRyDSjne1Z/d
nC+Mva+prLkuuAp47B77jfFc/Nixslrwtmr/edBoxKINi4METNn9U3rc+KCvyBb3
h+nCbguBT9KFQRl9cuEwfr1C1G0s9L9SdkZC2flxiZhl20fbuguzbcQF2YpxlSx5
/qnfrIAhw0GakrRYGHOVzUU9iA7tDsjHguBGsDCpvh1SGEmOmWjIsMk3t5A1bSkd
FX3zBWopvocnAg+hfwXP7uw0LuuBV7laepBtMc5P/UWPTmsWyHhEngz4gU0qlMX5
m7lgE4vqKGG4dZh6086zgVM1iWbwiLJ75q25TrKSNqfIBgdbw3sLgUbctuNQbkqS
cV4q8T9FtAcvYOCU/yoeFBIQM9cvyYk/lxlryktFCWG5W+dHO2dNo7yGwVKZoJLG
v3rggYeYIo5mIwmwBlTNh53r6exkVAAiQzbLIm1H40YZ1yi08uJACwSGopvoFHQ+
iKj8/JbGazkw+/JNhrROosSRikZ0wDMeqHsuc2O/mu2qEXYACoF5u3NRberM3Ygl
U2qpaELMfV4K5mEtDkeSX0U4PJSrsYVZMpqdjj7WuDSRM8dFGzJ6DRucx88On55O
DYlPUXXbA0x6eLQ5dv6rYXZPyxLyxHsefPxmE7oaesxq4yHUEKO7HoehGzZZERYu
ol7YPGMQZp7eT5Kpc0+LCJc3xsRFG//QJ9LW0SnNxETKbmQ+ERMhJnP36lwBJ1MI
/TwVpMJ/sElbzZeQBgVtHgMsPvrIjVT7R5iXBhIHdFBkI4e56Y4lavt18ne6mevk
RwWMSzzCiWwayehJSc+G46ijfqZWfXmeScXS1DPEGq9B5rB7lLQ9DkJ6n5uSY75B
4fbJOlGCkwTl2I0Fihz345ObCZTmnVWgH1GY5OA71ZkQoYmrMet1eO8IBEKXsSDv
EGm37gdxs4C2Y0tFc+OpaTwrpeRXFxZqrTfVIAipGE3vLr+3MlHc9kuRskr3q34U
u3KQkKFNmvEnpsvmvp9SJdZ0ETXrAVSBD/QrzxqMH/Bi1bl2EGxAK6iHFiyNZSpv
/DweUakc4qvZdWyU/RVcLLRuUvgx26lg8qlcQqFj2Fs3KNIXtU/eMWoYCmn8xDfn
iYm2dELtwAkJt7Rrl3sgPsIuAft/lgfAItmvtFwbS3WFhbDyZ20NfocvwnViibxX
UaMoFex/zqfHztQjRYIystNRXhjTu8pro/29GW8dEF7jRFP3yzAKo7SJKGRnKSQS
6PuteU9QMqtFw0eReS0Uf2jPSWfxOeFf5wh1v2v9NffbCz0rs6O3iWQxGTGeV0cO
XLb0r1tnCgNzu/LelWp6Y43AvRKlMnMfE6timtcZVIFkVeH4J0sP9L0Q5ZrnfeVb
FII3k4Cq3Clc8XIM2je/sqdVsEIwvwFrfpTVcdsixlE3WlgQBd/upvpNy7ib1ERF
WQ+rRfZ4tTDL7JJAUNlejzdotT9rU7YffQOYh5UNhxkrNeXN+yHQevt9WKPseHtN
jLchEKUOqep0BBiLFh1mGZkyZhqgSeDAm/q0FmGi7UiBBqe9ROS5rUu33hf+C/Tj
IzwRRROEVz8g+SLP8MY4L1FdSEqx5pZDoKtpy/MbaW6810EcNO+Q4wpILVxcNAli
SC82UPhZ+Krf6xGXJ0uKQRdHDFECXfP9VZ9hDjfx9K4lsJaURaH3Zfe16SGOh7F9
THQQzsmfZRbdMqts14e+1rlU6YEmTqNGtMWKjoJZa7vmUNvN3H0SUyPzPm53wRfi
paNZbBzKYEFq+MFG4BZs4TzYPARghklyGNZcQ8KCEcxxNTsiqbIR/oErNCLCuiU+
1X0vQptgPhTSExD8d7kbUXbC7UlPRbakDAjsrRTMd2hAO0zNsUFJsMB1hRtZVYqK
ZdRqT4j2goqkLqjW3fB2XEpBNeX413mMFRLqyiKrKVRsfZqTUVbxLtsVp1jXY7UJ
GS0/LBz2oc2Tlvj2Odufx7qLw6jAFP8wABIlf/Xl9hDWbCndRVVVNs27QMc/S0IF
ixb3eiV4CDZcOQHcn55A7aboNyLLkdxqwY4nLAEjlToWZUYufIDhjgC1dzf0tZ+5
V0BWDHiXI4UZUtJoZ835bZOz7ah/uLhu+H1eh1nBcAq5LpE0E3eBndC84BWGSdz4
0Q6TTJwvgqQKRmXZSnzQWSI9SWv93KZiKTrMVmDj741mos1kVpQ/5NARo2aIbGK+
AleAH0AOzHRUJK73CE/jyQsCiLz0bieaYg0v0rSFvrjKODkEprtulCEHMFZp9PlM
XbCCTUC0oYHVEwVC12x1IhYLtxQf/zVaU1uYX7r8oBRIk5ZLg9YzTi2/6v43pYJx
Lutc1xhlnGsIk4RTQZfxYyqwb+iQ/GM6MzD5gctFqA7DoWkP6YR68hTB2PwW60Db
GChHXKqOdDyhRpmNCtJp/GXMwgMdJOAXVtl4Cb54zeeqXeU4lYedXvJ8eRzCeCyR
JeBt0AxaRoxF4vvtBnEnPURZwqRs2ZrBWm6z1Ak2fizcIMLpbyPiYt3HfTNR1iyd
j2NdXgB1nTVxPymMDCskEx3tNR4qa3QyPCxkc+Vw00x5La++5+MxIGCh1b+xbasE
FkO6n2kmee0kPp7lbVHLRWaZbq6EQS2BqzG1zNNEk71JMb1C/RLVim9AHDUKm5kg
ElmioDbtIhrdrvzN/l9SCDqR7S8FpgabnizLLdJ4BsmSwMOq7YfqwUJ3Rl32LMUa
KS6XBYKHmR7OlB3wuXLvQJ+0F2wiGVi0DSZizGJmm6TTkTd/e0LhV3VkbCcbqqjZ
svmRlB062A0+8hWAIY4CnClY8oJ7AwVufnThX77cQcYXA8fyNjdSyQGVdcqVyAEo
tZaHC+23MFnprczEMGXWwjCcKfq3MGDqunVVPzusxuyZPQjjWsBvuYIFyZ1hpx2L
URE34oPUfizGIcjG1zGv7PJ7ZZUESRyFDH8Ad+X/bcNDyo+wrGYn1Zb46yLr4oA2
uJ/mkUNFN9H9Zt9YTUuuEHQkP8U1bxlVNqoGm1HwkOXqWPHxw1B2CG77VEjFVpcF
WIqHZDpfujlBTRr3l1mDjGnOiCYFQcWDvPE90yf6QjL7Y+FTU/16oQT11FWmY+Ez
kZeCgbTVCcKwCA9smymskfYBcnHBnhLccHjRiobRWYnrlokFFz8yqBTJPPIlrfZU
Qi7Qe9wVX3e5VhduUbn483mTXLeUXKQ0J1axjcJkZMSAsYO9sVYDCHLtQdJn/z5z
Mk4eSKxe4highSTlg8HPHEUUty+rIgACzK94bEH7Gcs/XWeX2L0xOPR+GQuYifPM
9Qsl4mZqb4bcUkKtNldNoxt3zT1tuZfa0axgkHvqBgyFJcsg7ANgxguLH6EzQJzw
EICbQYOkaIVEL7FUT/gw/xOeKiuI2QWYUu3gW7rhis2zjCTsNRhGgXf4mnzGOxdc
DfsOGhhG3d1qz6DNE755JfNc+S77Np8apOlRW9+DTrTFnhdKf8R86pNddrWmjlgQ
ES6oYsPU0S9zmh3XXYCAx40qVtNczNZjwSE4ORX5qtW72bPba5D7jd1iuZsAw9xl
0yz/sYErS5CrR7uRfPqx1ubJn9t8I/85Ch1Dhm4b0VWhl/EijmBSUWroDpiKzr6o
a70AE+w/60hd5R2GkhBHR8vMetPuDKBQ2qJglUD4zQAvL0N4ROeFHIvU5jvG1gwm
OnGXYH9hp1nH0tHiSN7qEMOSzj0KfGxrH7OHdMt2q/eGVvRipbA0MIwc1eT9TZyk
/lprJVYWxmw7xXwfyzBMt8GXF6Haz4v4vXPX2bzN/fykRMeZ94ZTl8D4sGDi/Wu8
Zwo1VMsbkzvzeFDzoYAK4u++paD0mJZi0TeHePifmpN79HitPS4srzWoHDBju0DT
rQOY2BYgH20yZdn6pRORPfbe6tpschK7F+HWpXwP/75+yzP81hyksc25D12Tynj3
YoRRpsuIO3Iy7IIOFVLtBDl+aV597IJ/es8CqSxdGPWwXBhuhds4UxhAcWG8k32j
AG1dUaBEXDHVKZsOOLncAVMm/vN/JBZtk4h/HZFywZWgDGKqdxBJq9xa/dGi8uRn
jPzkpYYZcu0sP7G2uujZp6mW1skxYdvAVh8jxUAokR2WhsyHnwK6Ynqez+qKTHli
zU7rrDh7lmNPKKH1wDID2n9mwwU2lOi8a/CDi4otihy0K5wIKZyGNLfvovhilzZy
7BEdnhlgxQ7S5n+tuo1b+poio5Fv+Yz4nglwKmHOjEwQxGHOflvuzm5avjyIIjvf
tqj+ys4Ln3KJBSZTS4tv4vLz6oAUQGBBbClieyl0+GFYM0TutfGK5mTuWOkESeFK
bY7W6MbZztzvzGZzC+NcZv0H/s1K043OCdtX33BGPXxE1UTyXvzIXSWzRT1Vbek0
NOQ9tlfdD2kkrxsjM3bZKaE+7xKiXbime9KL2rBa2j9fNizN6G739N2+HH+ovZ00
KzBb7HCdYOkUNzF7z61vmU+8VtUFhgb0GirYhzupFWV4xD4r/TI4+r9tjmkp7up3
rj4a5veK8aQuqM96fc4EWpbQk8F80S9EW/RYhdbRnJCck4sm1aWRMkzbQJN9gPRp
rR9PO4swfmbqD7MHFOqkMh66HQrCqKKtyQfvqjUyM1ZW5Tw8DQ6bTrScR6YC4P0s
4F2Boh/blykcA0TablNuLIOzycdwyI/vVSU8WYKjcwru3O4Izr5TRlmT/zzMCSlg
S+4NQxNgsOyEh8qf0PNI1nEL+/m+83extckK3WvA0vypy1MSWaHzj5w+8mLG4enO
XZcsJUPkR/QBuc04NwXUD54qsmrhmY44I3zZsvN9VzKGsDsQBkuPkk+iLtwYfFGi
Dn3I7zHgLWMNYed/qZAlnBqRjiVnF+DrpnKzHbg4oifCJo0C8uXpzNmG1VX+wNyQ
nysXx+xpOL4JUWkLEvNVu9u2vJwtq2iQ3V7Lg9Fh6vk37Cthj0pa1UOdqhuD+5JG
IsfhDzcSHxhpwjS8DtPorQDyOG44q/3X70Q2gxaUl+7GNAq/dPx6zBafsl6/5xwc
Ro27C5JsInEHYrvq96KbhRCKttSAdFZJ+Nrmt4nxQNfQC4euQtCrR/RLdB5sZtVZ
q07HqympGX7snvG/HfLIiIdO3HhXjGRWTPMZjjTZVmPjnDoKO7pOjZemXp/k1JMN
jv9k8yeo0eG/GRbm+Cs2QgLx/+ug/x4dzz4c8GxOhFNMayVmey9ItnzA2lYnfj31
gWe2tisYcDEK6nftwQUkWW0/rwoDjnn34pZd8VFpg78Hg0EMISzvLo8c8rGb4GxL
62UJVfSlhnZmHTJwXPU5oBd4wlRdZqAVlrRygWup7Rhq4kEdEtoKBY7NQOJDe2eZ
SsJRkyqokIs2T4q/e2MgREKttjIodk8iJnTHsKEjFCIEX/lgNEUXTT1hHdvVMA5S
bgDu3Upr9Ls2qns7B4mk4jB7vH3tWnwotnndyfMqSyvURG921UerRbG8IUxBRFhr
0LU6RwNUoRhkRl0kisSJ9HxXp4rbZOuRUPaIOoqgWEm1LeRyH2YqzWdtT3oXnds3
VBVfIZYLkOql613hP7BWn9uFJ/GDr+lR8sDmEDLuJ2ig/HDRhW+V9x1lwvYi22LB
dGeCetPV5cUhXqO/eUk6f4UioYd9yeS5ahPbUWIpxr1ye625bZyDycabAf8cgRX1
94XiP43B8pqj5zXSO2iRIUJkvHPgBycUqT+Wv996AKdO/dtRSr6fNzOQx1ttIC3W
oFoXjOZrQoNCf2Yxndjx1UF3Aijlkq9Uv4DwVgqXROgkDSg6Wimo+pO2ec2n+xOZ
TSIIjM1REdXYjkDA2DvHLMvxX6DK/eix8f4NqOM+z4yKwAVUeEZfcXaX6xOR6gBP
DQdPgpvJiWMHtNPP1NW2VzdYl2V84iqeIqYB+RH3cprFWMiSPB8GgFTHtN3G7T4B
v6MP3KIW4b8c6LeMl/Adkn6lg3u0mFPEayTlxKciSv04I9cM+B673XWewrwRu8HV
MwQscw0tIQeL5ao1bhuTfKrWUUeLmw3sLTv+oEGN8lCQDpSJcCy6gl5WM/rClJHM
/2m2WQSF5vLqbsaEihQMzJnrDZkns/gaNEZXMe+Ot5lBatc/UfBruPr/eGKe2Lkn
q2G1nTcl0/spqyXaKj541Ys2FG80zAMI6pZM4KqaZhkWJtMuMeXovXtx1g+RsNFf
dNYateDUQhxk3LN7m96T6MkD6akcFq0rS2HULkB6gAHD7yp3oBfsKByNFJ+Rdtxj
6HEwUGugvqOt0x9UwNUskYMskneqBPZmxYUK6HqpR00O0iXqPV3b3Cb0I1VZUE64
sQVo2JKrAsdKznRYID4x6FK9fz8hRqX9N4zZqOP+ilPJREwnjheYz3kQQWopvXou
zhfU4plCN9kLVnd/nQJI3ezdKQWK4iivnewXh+UZVecXTweWXrHfWV3eM5DJOseH
rDEeTFNFaJaG6q/yi4UFhDyTAKh43OvVbfLux2xGdbD/hTjP7BYKg1b2a08Zu4xN
f099yNUahJMAf9jSDCswd6Qvc7tix4mGquveb4lE1TxdmrqG0Gn4XBYndq55Uvhx
NVX8WLXJNn8+jgQmS+i/UygRhD7OiWkLhMWqHssGnkdm+vx36yVA5bPvdl6LMtBu
8KtQC17wl7FU01qFQuiE02T1BZGRjOZbh6BkDY11PRv1yawoTuY4cgYw8HF7E7TZ
5gGERYTulYuuIbsygqetYQRoO+DNTBPjrmuYA3P8RTUbDY01lZcHAKdHhdBS9Thz
78cfd1uEIK62v6fVJRHc38VtrLBscrXsUHac0YDKvSa6t9+MjjtjVGkj65CT5iVz
cf8QGp6mWfdveW1duZaPcPQRIoSOW7DFv26Qs2FASVGAk8N/54OGb0/dOKuPrNGJ
JIS7sd4GLGHxFeSrZ4zadyLmFLaJe5lLWxFkUUFHrWzu8eu8MPE6mekMx4b3BWYE
lPXZX89hE3pTiYW6TjwCw8n8cTZWf1KHWEIBNXd0SU0TW7KtvDPVDiSw5/Sd/Ltn
m0kH/v7M1sOn+TISRvazqfO9vswBk/WSH9maUh/Ub9b6Mf5kxkJ8xcsqLsNGAaOa
5InBxWjYv2gpp2DDdraaAkN0qHKIBT7PnnrWh6gd3uAq+d+lQIMoZFWmdgaooIaJ
1XgXaBXGIhWAuclibIMG1S2qbkpsR1T3R0v1ZdBO+Ggu+Y5jPG2uk/mlkiTAF46Y
DuKt77ToMvpKWElBRcFPM8yi9KE9frRPmb+X0vPU1tHHSTjc23RILWK3Lq0/h60l
WgUcleFDQuIf6cUlC60sSnBSmdLxxVDq4Jg5DY/S+rv1BTksspFNoZUPWMoY1kP+
z8BpxZm/9d9do+zbfvQK9qfmZ1wwQA+eDqeiTGKuQivN+z+zqKgjuFuDC4dBYGHu
QvibBqP1AlUOsGZRdRBIEtKGYbRKC6I/HqLvckD8sRv1OXjdawIFSTnzPJ1wQhOK
Z+vjgmx6u63OeHqvwITxVkQNVerKkAuxykhYU+/rLxg0WKoAf0OKzEGeWVOXBIFf
WxODzp1UwhIWsBAv4UMikmPswARisefflM5hIThHAdhPHoA57G+63DtGlhsE1guz
2GJOb5PDmqqfk3vpxNFjg11nxquQR3nLz+HGEl3C5CrhnKZxUC+d+vJfgtgG/yuh
vbpuQ43LTpznTPGVITulouEP64syr82rpvjy25slmWVfsVCcpZNSGEfbaiHn8kGN
Pk/7PEhem6wVCcrnxH3MvN8Jnr8BpWS+XzzQIZIyMynqmzaPRdhDPr6RsXRnHl/v
iLyWuSShqX6D87jkSTRsrU5p4KIFZ4Jv8jwKdy7dNq/9eqqn3XEj6KT28xCeFoiI
1f2feuHYEWW7Bx197hicy3vG+2kop3jyqAOpgXtlvO8nWE5nRf/n6Y7WNr+cOE9j
KOt5jJjRH4tkO9gkTeHRcpwtV/NBxMiqG2DuvPxcyDcDNKuQ+OrRNPofoBqp3W2R
o10XrJVTh7uSbLpAyDgByUM2mBVSPYbDSm8KLJjfG54t+63OLK3+jCzb7Bt56dJf
pWPNcSgViMgHJemUddmPMYt9KeOhq0MUGmiWF/pON8jZlm7U+dbwKFWV2ulZ3/3x
PAW629fgVLWNqI1xI7CRAuaTSDanhWQ1VAwdz2XqTvwq2PTA+y2D8POAM+apEih+
zlJ/OY9wGC252cZ9AOkIeDra147w+WeMHh+871OWhnXEwpRBSu/Jz/JBUBqPJPVH
1MXSmWVrIeIRk/neXkkfBIMYXh+c/rKGG2wsy4Cj6KA98ELkxezz+TKOrX9UiK2g
UCqLUfNifLZKAdq6RPA1zl+HUizXHd4X6VaT2+owfwR/IHBfb0KJi+tuH1AZPLkh
dC8SiZsNBoR0lqHdVTwIutcHpl+ouQuNtGqk1e1RoohVQqbKcaGPCJJjWAegllGH
pX6tx9BAWncc3pIvxQHsQZ/erQd4wa3XruOFRE+KO+IqnDCVwOg5qswRieoGhPU+
GqiShdG4EEPJtlrgcHQ6ZZj68QyJjyFl6iooiHMe95docXD/s4MDh4T6WfJpoMIq
5zTFA1GQfIWRgGssDIfLGbPx2nLml1cUA/bxY7XuoewI9cO+HeKVsChC6SkjqAtx
QSj8qU3sNITkBn8kVT+6NVZxsjCN1rU0WPuvrU4FDLUKlziHnUY5N5ldBKYD63vL
LgD7aS/ogmpFCe1YApl1lvQJCHIlgO/c4iByHViFXXO7wnizoUmHt04aUJ8QfE44
aW7bGsytt0Hs3Bhh8cZPh9hnUijIHSOy8Odm3ID10gBeTxGwxgVJ9/HFXbmNtUD6
HrP3Q+rDb1EwfLDmIwYmzhdnjLK5iqkEWBlqOogx6uTHGSbMgWPVsUs1dSM+MoLq
x3N2pzLglgmWdTcJokp8A117MjeAFmesl8srkGqqrUVEXTuD6RqAT+AA8npjoARy
80Rpd14ycCWB/3Y+oXsSOnGY0P8w8gxn6rJL4LJHT1n67UGnNn38f1TvqCaR/hug
aategK3BvveDZrNwIXsgmeDsMK+gqAVGUDObCYb7GHl2ZiGQgpVgm0vL/5SANtDh
sWB+nolE3tnFKF+RScSmGR/LiTtGHXnbrq7FDf9z76+Lf+n1wqyRkWGjANhwwlX0
wILgSyq3gedyUZ+y33qpkcQfW2NJJY9nFtfIoyFMzljvq4Z/XQzXPqPXIFNqJh7N
k0zlrJ8RaSJ9lH+93wx7eCn3euErX0Mk/Sot4DOXOtQFNZiLB51AC3cBavT/FhM9
Ww8U+0kHp1OVF76g4XatDVKJwmbQXLLVXkyMfkp090QiXDpDXarmb3SIkciT6gcq
NJSQFnukQFbknIzsMC4BjB8QGyyafWx9Xp5J1CMCATpeL3QLBH6kPziW70LfQORB
HW23NsjReqpBt6rIMqsqVFDz+nqHB2ILMgDCC2FgPrWVtkzsNsLT8qFV51gYkH6+
LzZ71eSA/xs/d50mfPNTapM8hmfpYZhOYQu7bmiI8VExXXOu/AF5CKWjH/KR6LEt
KERKyf2gY8san974ERUV5/MJ8MaJtw1YgaecyM2xC1YRAPRtvqIcSZFfWTPWEhK1
cc8uzyJQ4np0ZU8NzV5x/W0R1kEKmckHltkup5FTDkQ2goeOOyeyQ5cu/mfRskt5
9OgtQK15AjTS88s/SelQT8BVl14gPQ6j1seT43ZRCnc9Wycke7GYqF6myQJZ4NqP
VhQ2olwwhJf62IXzePcKHf/S3At6+sLN3GVZaOwR24nmOPpuX0i3hhkSxja71j76
0Cqv+bTI/CDzvObY1m9PElSAmlYxtyxsKV6Rw3F8pLCkEKwIc3yUom5hbHIa5Luh
dzujfAu8+pDxbvflhS/OiDAIwx+2hMspzB9nsF9wxKYPJUFcADIOSmbALu3le7xG
vp8TlbGTeKaEUHA9Oo9ttiwcsqvHRX4WZtGI7Y3ZLcAe+YLfLSJ8mbACeNDoGb3t
Iarl4+zrRqgsnn6oWzb3b8eXfQRAQ1Uy2K45wCvkJqCwUkQtXuaDEXzly1gitgzM
Gz8xKFemzmAS7JA6z5d2Uvw9g68/b0WCVl3b1iPPWDDkwRKcF1WiCQtdw8ze2sSN
0ljHisArDVXVfOxwv86JBkuL7KgPQSpAyPimLMSFVyMnegJWfhRDCFq6yXtAs/jc
gc29E10b5kgo2afNmotx12Gp6nYDVZKsfcTb4/fR6AoYidavgc9zqYOof1RSa+RI
tGVkOzL6FAR5z70qA7TaN9toapoNqxx/OmYVUY4wCHcIkDSsIyshR/ID+B2AQHNP
i3xoJF8/1XMZYagylcZ+N4of3b+7By9MduJgyhuxXMMIsmOLDOSexgHF3fUJltWp
pdPLaDTkIwVzNfT4GA7T8jfZD8q0rQ82osaFqzxP9vR3P5s91SXk38VHu+gfd1Lu
JTHRaQSmTclavWCNpNbW9/8w4dztzMkLvHCB0SMskJefh3QHWpz0pVfgEtUeGR3t
IShRe3C7HvhyeNvQ+P26yDsm9awmV4SdHsu4HES5h9rrzzgLlTUGb7WQSqeV7csh
rOj3RbmR034tG/GPBGH0NbYPn1+SeN1cH48J6VJzsEE2F1Ml9mZr0bAhQRl6PFJW
YWBfiubqxJrVb4bDSCOZIqrVxG7LAt6BeYwSWRWVZw7GDm5SsOCLTzB2cLM7bgMF
HQB/3rc+YxM2D+7WIinZgicE2gokC1TsRwyUFUjsqT0iqiRV/8oIyzmt+0fhhKfU
ot2WHP4Kw0N4y/PkCX6Y62UYDKbKRLxQU92aqR1z6UBn4RLsAdpPQ21aLO146QhX
n398VERt/PV6h9Kli8cJyma9RiexUBBUOiLegkYLk20HBl9GvdHPK3vo4LhKgwwj
S7zKzGslLHLleXMu7hMpXHHcirmGF8kTHkuS86QSW0YJGKAWWTbDhwZDeUcUV1CA
M9PKqQL04CQZhQvjnwZrV+SXn5bATJKi4d9eowXzGHZZ3EWrn5m5k0GFFf9M4b2D
vATeLa5X5w7KwgMClubQMjVRwMXl0HkdroaBLJA90E3T5EdL9iYpxYDvFG8YEk4o
8+9Qv8E6Q/cViTmCFcmEfnMXieXZBPNJxGe+Jo5DLnypWZpqAHFRov6SP1EtUzoc
KycgzmXpKjuEyg0rbb/zWt9S4+J57yvnnOmaHlCiY3Ekqhtfl9EIsT7o/4m2eXh1
FqDAXO08jfvGf0aiR2iBXT5mAl581tVdcfobjXw0rCZ9UylpNAGstCYWJ3/dg041
Ycg7Ibf+VMlMZl8oDb8zywKsro5rPjmMrvrqibN6UcdunFZ66wT90BbWkGi1yfg3
rO52vXJmniiSy8VaI7lF8tudU2Frxsg9BMwzoi7mL109iHCDmyzC2BEgilJioCU4
31zRDOP5qwqZ/j3x4VJG0suapTZNHUHLGaS4qVThJk0iPZuspQIDqL3bx6e9GeyA
WG/FuHbEzha3BAam/cFRTVZa169QsCeitAPMfGaVPONEZWbPDK2TKniF8VnoL3KV
d2UyOt7RPcuoO8q0FTvSv9Igstg4+LjkPGQxFJOjf4c5AWTqb9OE+BKLFstC06na
VX9yRQTFD2G/gEi5G2ke8mVpqS/gyjX8WxGFYS13MZobZXV5cKxLzfFaldAc1f96
h3VViQr1gOFro22V/B58PZXqzAiRG+eCHmBFTj/VmMdNYfMG8vRvsULY+n90R6TU
WZbJf1wjWdxTDH6wSKbMwRddMir1wPWKb8NNE2MfcsWEKsNWjyj5o4rNy71srO3j
74pgVwAvG+tBYSGnfGU5gLRmN45B/LNKu8pWI7cQahcNw/90Ri0OPTZ1/WoOXBQG
7zC6Fb8TgQff0OxWcogjpzbC0ZVYdqVmfGkv7SCRDYnl28ObNJw/dc5fuf5Nsvsa
wLySRA41kmMDdVO+QMyoZoF3j1ZajA/zXEl095qJZqrS5wsr4EcSazcn0BHpHXP6
Rd/j9otcUr5AmZaDZbtqv6ka8QP2rbXxjx5VYfJImlEYERmZ21tnsAp/uGNxAW3n
v0hFTeC+vqSLSrVVRhGL79S0geTc6dNWuG9xs/Po2qiv0Aaync+ilhNvv5zTzWVA
hls7qqDyaUfKKDoymSMWXAaeBVC2zHD1ORTnseqZgFRI/HeaFued2QFdRV4Nxvmh
Ap7Qe9AJLOaDsDIzyQSN66tokIU1cBHor7QYEL0YrADfCSeNuBdNMqTU2gid0omR
85LHaeykgylOAfzlG+XQovWES1RCsSncO6I6PBzW33BqKt9zSIeIB2IA0FTOrq22
Jo0GEkwlztBeHi0eOF78AHA8xQannuhQHRBR9O5Ft8o4UrZKIIa9FHcVzoyDHczG
DViaJRYXr6rNO12Xu3ul6gc8Z92H3Aah34RqYrWJV75KbYeW0iHl0ToTgMnvCZbh
AdCZ0EhX1Ts27KHLrOwHlbZOD0fdxtLLXiiekSip4oqvOUkssE+Ynd5m2/WBf3F2
RxttN1Hc/8ZdjliQZZFDyS2HDHXN83w//Sr/uLTfHWMMFi8NMf1K9QlitgQt88ug
0BlgGaq4t7DS6RNaQ/puQCT+zFsxTdz/d2qae3HXQERCenqsS7gwPFkygvZM2QLj
uaM6/cu2mT2tksT1FdEH26RsFXI28LIhJGkVWLbdJdkMcWXfvKwIARnsmUqy042u
mZh8DVvpnXejyiz+FB7GAsevOt8VM6+txmuwh4W2bh0evWaSzo3uClXfFTCtixJc
CtGlHm+32H0aEaCuFK4y8a0coGZQE33NL8rRk4DxaYcE2mGY99BkSUCGMm1cE8w2
1RPUi01LpXcww94tzKXfldE+6ENwFBExoixLZ2eF4BpG6otgxjeUBHidauOey9zu
WgW2PL6OyCIvZxceuojhTXLokXoNbsLsC/DHa30qYYg4Ummq8Ql2fhhVtes9sJJa
+h9hKG0Do25mdkvq2u8vADK3kAFw51rtlVXgX1hnvEDkGOdoOGU9rnXgKMiVQGom
pYQBKhNNQsvyUj5HbvrcRW7RS55mYJdbEshZYJTqMX3mMFKO/rpo1LEowyWyTc73
UnSQRCkZu6szOqJP47B2iZdzvlKURUx0FY51qY2gaq/2E8BRBbX/GkJrKpIetj9+
0AAcgTqHvktvvfFkeVIm2AoUQYyuDt5gzmS9vOAZcokomWEyuEsV+tPevDbIVWF4
JNsc6G+p25xGN5H5yE8wb+psouIgVgoSNR212PyZaLwCgguD1WouQNzeeD9WeUiW
/cZD6c9b29OTLgYWe1C76DRjWPphNJn2of0svPbW0JwGgNBm6Zy0xyTwv9UFar2x
nlzQieuWgYhP826zF1kTJXSegh52ZUR/oz/7BnLv6TBn+ZTc3mwwKOyLdLgD5oOi
cWWHZwh+S4VHGvdZ+iJgx6NVpRCXKbwstdQPWGtB6boC50L+F9vzPP6b5aoba6mK
R5D5rAEH1PoIKkgxSFARF4mLEXz/AeqTgsQIvRE+Z9Kgnp3YuYYtIEaolwYbElU3
ONZS5hsInEaU4hqtQ4QWvSDtN0TVUT02s3e2IplMG/27oGMLJWIxgphQ3pSoGKuZ
m2/mZK8HKuFhEMr6Re9nrJJarKh3KEvtUfMfaQCm9hXIY/O2OO2pL5gB/xAha+I2
/fsbaHh/gLMvIVmFkXF7cl1CeremH3l3zuNQp0XpPsHZP7rqTApMbQU2ZADJS++K
DVQrhzvkowaTOY9b2wIlvk2QDUEy2cpT6LaEQ27WhL+F2XGkrq+p9WvUr8B89roq
rAyO22zDwDytjEnYvqJS1fBX7rfMkZu3R1kr5Ia7N2kh/zLAQ2eCwcpSNT74uS17
B8ugVSXhllmRClm/f5+rhu7kJ9502ShXOw0Fs5dRVBJvHDk2nakDeLgsEEXgK1Et
qQLTV2NRSZ6c+JZG6V4oQhCKJwqhEqTC8Us2ewnM712uGghKAYTTE63U4O65XoCg
Y0v5K9pXoNbYXA8+SRMlYe+I5MKmnK0QXyOAJC4zci2ZcGf/lgCkvn0MTlkPsjrb
TO7xtwjmoBUF6nZfVAfp4y/nWDOpsbqXREYJxI1VyRrwOY3WHyJ6Tkyik5lh1+XJ
PruZKrjQ2GDdPoJjPhT3KunKkk/rUg+GPIL4F+GJWIlYQD9C3Uklt1L2Pm/5A6GO
xnJbqUce6XUWSQPsA4OpE0QByr90lCHiULVEL5Y5MJ0R+xoEMTcM0v/NTu3G+RP/
w/z9YJB4Poz7Vb1igrZhbXhcT3MX7tUGqq1BscZ0FGgy30gfwiWIEyIPqyrDH3k4
UjWG1iNM60YpwJz5jPaOH+eHjA0MkJkYbRMJUB6sX2ekhWwCUgITEq1opllrWi03
qMeoMDX5VPET4w/mvLCbHMRifWo1KGyQjZs0A8XIuBxhe/QPgKcYDCmGwqF2LIfi
xa5KAU9Uw/R9CwjgsWlJR/bpHrkFSsixzAdxtfZ4EcnwOiDfJN05cRAHZ6sPLysN
fn+lcTTkVr5TGk9zDbkdatGV+6vU2PEsVZVfLub4FJKtOm2mevjDPXFA5QbcjZ0J
ZV1comoWqNLqrl3uq0XaXu1F6kNuRDuvY8yz1DgpJjaC5RZUvCPKH79Oj8rX2oR8
XLr7IerWDPMhqPmNQi275L7cbAMY7i4aqRn5x8IpRvzmgBBMks0FaJZ4r/uo3ejv
nnkzv3pUgYq97si8Lr03WPHvABqQCvMa1TCx4Vjs2lXQUZlu523RlDoOk8rtr05J
4PNhMBEBvBsiHykKLZjJGBNplAUwyRQCiKuB0WM+bI7FrCcmqqp8Rh7ipcrqqNKq
pslqtjsX4tb4+lwMZSvxx6WdqXHZgsfj2fBCRRvvCjFVlS2z/845g/GWzfsqjFQC
9Ks05DUNsMvh1LyVsfImDYFHAXbTYRmkj+jzWz6+pkBMy2hBPFcoThRSpi0nJoBR
qkFSuSQ6wAoLD8hq6kWgxefNtJ3ELB4bf3wdxhAjzrvCY45ysIHA+jPdkxMXP8lA
nnDzB1g77eRShNbBTjtgfTNSpOt8lnaiQKTvwVLODuwtvSDZ9lqfdvkYapBHm744
Md2ptUWxhdBwJjk2MKb+VRKK7JT4e+1mDQUnBMQdFuI0k3orLHVX6LGnXrXyKsMs
Q6OWlmXTmyr1n02utdUj/5awYgV0qAqzXxEFeQyOPun1Sp9m3qwA9YdOaO/e22wW
j6IRHJToE8abA3Lf3ymCUJc/0QCa+mVMxXPBbirSgM5+c7j57zj+EQzxjMzZVPhG
/wXMLok6hoiONpvS6oOXMKE4UiQJanni+iemXXMW3MKt/x6Q5GxBgINFjDZR21ob
UoVONUw/fH9cq+/6cQH/Jz5WXlEE8qBw8MUoBUWcPDOXFHR/rRUG3Ws7Ph/KHzsF
a0vNM2MHEM7tptDQrk0bBaFvROtNbcvu3Twmx/mRDiu6plvtjKEsNl36uN1PtXyr
zx51knOuyzA9d6i2zo6/z5pJQfCTDTNjQcm0ew5/EvRcRdpyUbTIbmatCRQamh4q
rQaJ3OdTi3QOPHgVkALf095lHVs0XrHfOBcg7DMB82m/Wa4UPHswM0XK0+swi9J5
+iSxqv0dKcmrTpC9+vdIgY8VTI5ndMlkQ049qoS4Y3T49lLAlkYnIoW1SSJ8IMZb
QHdI1a4L7GFkB/VG7d2u7GnOp8ayAaL6z/fFiJZ3/HIV6OWvFy06qRKdPkYkSaxM
qWHnkiIbKFI847M74ITnekL8FzWnmTZCkiNVI0iFwUFVYCdlJQtRATh7HWcYLAa4
OzBTQaMfMnDHA7ZKu+fn6eS97N5PVfTwIfDcgNbZgrGCYu4MUXwYs9xfWmJ/Zi5d
OyGxiJ4FXtvvkrk+jOh1YjyJzSgxkodrpxD6IciE295OAJUsh+9WsHMhLmf7WOZx
WV4gAErjoQlRETKeNCi2jNmHAMbdS091IGUvcOuG/613KD/N2CAp9Bne1BrYNoUf
PiQyQus47ZmagoQMWnm1BoKTtPqh2YGG/WQE6o6OQxMv4xUewO54G2TbLAUYnpl3
sYQQUJ/auWnPBMvIFa8Yd/Bt5fnofMCJ1OlO6EJzTYHt90TYiKzXtX7fwGoZuuVF
yrJtrYeHE1fzBArp5i2Cu55//LIo+HdKjtYU+puBZx2FAiWwYilxkmYx+VJGnlBc
LD6MNzrRCqrJAUVVwt8G60nkziOWJY6aBdsDYrr+4FtYrylmHzjeEvbTm3U2Rmtj
ljkKwoQaDY09UsOVKZKE8oQeRb8ideiW8tnyfXqU27dN2m+bgp4M/bizwpj+d2u2
QvvJWG2CAatLxigVMqxGxZiZV74rqGDREOWjNVPyv/6ilruDZ5fxbHaS/YdIRDxQ
lpEy5z232PzTXQpZQKUbDwRJMy97ETXIchtMUOkcupjp/EtVFJkuflhASj2caMbT
LOq74Of7S2NzPO9VKwmF4mtw7nI45srteL9Ow7ty12J2fleV2DUeRofSXTRpCLjE
DSXo78OvL7BI9DM5y7Ui+P0i2R6uZoKVnHqtGEdiHsjIFLygH0QB3j7vonWqH+58
vT5y1mm/W2miEUqxbaXAriJhbfjpI/JS5mwFkXraDXnjUkfA0gwfaUL2GbkviaLy
vxDEa1g/Jsmr+0WD5K71I0v/nnLmOgnlZQPmIf7EM4o5fG4p+RK5Dzt5vAEgrhGF
xSLOTaajaC2KHjft5qrXPPWoH97qJEE+XKfW/fVtGYNka/dIsjGyPXlxbE8hdexR
+fuEKerH28MWuM5YACB4f4KyaQW1y9/g3ZncGbWXdtQsCDDszompl/uIybjuCEb8
tiUBdHOn0ATNJsZw1yS5nVV6I6yDqXv2Xb0gYEc3sDE6yxhlniJ4Fg6MEdKBOQ9q
FjP1fme7JddHktwUV4phJsrtNogCMr4oFRqi17LqOw5RxEQxpW2Qm0UKV9EPMqpt
Mbj7JOSZOuVGVm2fHHRVE0FpMdwnpSHDkLD8xJBqP1Y+lBtkoD7PA5jqW2Bocj6I
Pm1DA9s9N5J633NGtzJWw75mGFhKllJo4nJVNTC9xeQRJKl9mwXVVUTtwVWsXUCQ
qFIrqRB2JtTaziW2xUI3hyMaYjp5PZrSNJAlIpbWo+9A79GXrxZQI+d8eBgJ+2PH
89J02hIMb9gXEN6u5EuluTDI5Dt84W4hbDP91cVTnBiu85yiP4ShOtx/sPkVLbbr
EefODCsVc1LyRfesAfujsuvvme2D1yckaDvTvMnnA8NhifVw3qOWV8dQnePWZB6M
MASKgR49QmQBWGfwxZdrxRk4fZ+vq211XQCB4+RM2l0zh1Kv+2m4Agcpl8WwGtXu
d4ejwQPm6GxneMHbPA/ga2gav8LGqp6gwmLtHoeWdVC5J3SKu/EQII0DwwbHqFdj
J21FaEbIXB9etZwmpsZ0q2Z1JWPV1Wto0bZATVPHL00Goe2VD/dvVPrjUEQBMa8G
t6RcV32+qwHo2dl0Lpigo4OOFr2v7498zQeGZluEwEaBat+86uiScH6EZZMizU7+
dYw8YeM6B/4WkXaFNIBMIwceitajnaC1uI72AXU57kpt4A/GBExVTRFZn/yNbkwi
ijugWK+A/010JNse6U8ZzCo5xCRrdrzpANkNg1WPQmAPg4mxLMHepizPYLJPwtXf
189o64C8Sz+i+iIyJw44HTmYnQ3OcURYGPLonUrB8PMoIlbXlzAtoSgcE3LXmHZ1
LfLWZS8Xk/R2DZQdkfQmTSPVkAKoov6SWCwpqbAC5cUpRMnFs3GGYs1EbRh9Fk61
o443v9rUSyI/5tfgJmIQfeboTi3fym+GQMVUX+UHQOw1JYiqWA42kRCYIRZitmbp
ImwRoEaxmkeEbxUZ0zeNXE4GLkLTL7jctlStlwtxHLo/LUlY/nN6jnyKoi8kclaL
l53wcTV8QL2DTmIoegStKf+7FkEqIwreGU4TbbJ0PqtqbjmPuwauKZiFgwToMg0p
EU1Qz68g3QYUO4YIm4+Oq2O79TUcKOsugCM2lIxbHU4zpx6nJ8DpVka8Q0nNZ/Bl
EpNXEhK3tPL4oR/ZeWr/tfg7KVbpQblSx3mUWY3WwV3GjwogejhA7WoVtx+EYzgy
0jl7rBg8Rw2ccuHovp6yBrz/kzqzYJ0XHVrtlt1erxEGjpKL/hEDVWCueM9UWz41
ShcWerdAy4pKevKEzPAnQeMR2yszcr+y6CSLKeJvZy0sjaKWiRn6rDA1aX0xEBdk
o1JhFYxDzFeQjDjayN29hAOeiEoYJCUNpqVx4hKtxO0kW1SnXePInVFUEfpH04YW
1XRBWKc9QqBWpUSSV7YrGeca1nykYKox5G3n1oCWe6S4Q/fXnLgQNiqKFB6UYw2T
0mozOn3MnV0DVuLSUUEAKc3NaQcVbcsqEuP8fxYp/7mOenS15GMJ78TpfaEg1/if
FoZ4p/4AqjMi2qhrbStp+DHmMYx+wcvn169IaRmIZEYSZUlWIaz4JsymbrAYySyh
/i2NCaf1I1O076XR0HCudU+xz1l2+EYsfc6aOtEE3l6sPY0+xWmBkGfr3/q77qFM
qCgKRJnTWno+JRSE+H0u3CGEOAIWfBlCXNsRHlb9nJCYKSd8OXD0LubE4VqqEob+
SMI876W/aXxnqXmc1WH5BryIkcp2Q1eOJnf2IsTOujNvmfpt5FoXiDP7NocizPID
AubU+EzF2faSqqZYD3v/aIj8IQI3y6D1yU+/moxsi7A1TwojqeD03JV/CiX6TegM
dXa+2yWXfs+C2EBVXmcjwdwhBOim0ma1pX/YS5I/RUUIF9kDPq9VaAi3WH3xMlI3
D+EcMoL/oURwhTfDM/EeyBFRHbsItZkMrjbKl8o57Cmb7b89kMoUASxFyuwVXXsx
hxfrSa1da/QcJJ9zcwjZSC47v5lNnmqtz7JtFRu666V4FoAj1jCijaDlofc6XjeV
OhM7WHI3lQHCeP8Bp81JOQJwr974FqOv8zMvIDlY/WzYJ4PuHlhVDNcZ1AUoihjq
vLjZ7UOVrmBgaRnigsY6cMUA33XlimOWW6bhDt/OGOuOTeJKaI8KwaWb1+KjMWAg
663x/WkrsLhUE86Pz4uLJH9BDBN2it+0FtjoJnOdb+L+56uza3BfnMYiK8p6DD1c
CN7q6MGoKCkU/jV4pa9VPaftsMzgNT6PVFMNkvvdTpASWmVtAYc9KoyaK2YW9qoI
QfzORuf9L78DVUDlZSGK+jNCt/WAxZB9iHXGNCPm79wgVV5+b76+iuWUBNyresus
aiqJRuJn2WlAE1WOBxTuZmG/tcqq0rpACQrXBs4rGAtf1436iAsOe9SVpDSVLAEF
7mPCz9KIBgpqD9CEPLE54i+oNtQEUjwBBsHW4SlxWwdk6qfchKPpkMhgwABcEZ/W
uETpZ46o9iYF9XP7KXHqQ435dz7nmuI7GiaECxrT9dw1g93UBpRscYxU5F2XjReK
VlMtbre+M+p2kouB0KI32g9nvWgAmDmZyKsWw9LWs4bqn3zbiEYGEQ10dj9D5YsU
+5uUv3MzuW8Qw5F1Cyeapgy3Wqod2bV89+6gWXe5dI7baqzGwGzJYZ1JI0Gg0xiP
K3Ux2xYYqTa4ecdNcSQc2wN+W+IiIfBuzhix64S7pYOkp+FvLBRwGKJaq3E3lckt
pxW+uFFVxagjY3wxbEsO0ld9Ykowui54y9Tygo9CfYPcsNaHyTUpAchBI//MDI/R
jo3cTzzEu7Bop5kGA9LXbGARjn0BuyElF6bHDv9zawJN8ljtFo2s/ZR8zNDtXQs0
wz993xas3LNTaAL+YONBSNa8S6xSXwZHrIKWcw6PeWJ8Ih7HSOqf6myBhKfymmT+
3WmvXAAO7c5tYf3g3h2U5eONy9tfSB/zVL0MAeSokCKE/ZQCKs6/IvCqkKVrBQvZ
MFv1NPQc249tRGi56hg04gBKCcvmrVE1M+LuQ3QzTOReJRGTzDDuPZIbsMBPyZRT
JiDZvT6Os7vJ2Gq3zV9gEKUy2kKHvb4EKZG3DMZMWcelAgNSGdynEpnKatVQmuFb
i1yyFlimpg3uSGRLGb0NIAsj6MfItS43dr2r2Yhs2yEGFH8fpieNyPlfhM1glFri
SVW5ocpEjRJq/QzTJXganJh3Px+sr23ghBX7bbl1K37PqY+/dNWJF7Xd6ZqzSXvZ
/GE/HfrSiT6ZeJhnMhq4/bQ2MuO6bjuLVZLg0YWLl/1VSxptimVaGU7pfGTBzDok
8K2gegVCxJf93pkl8Wm8XHvdiJZGThcdg7XF0yK1z3tRWGgZyMJBiw+Ty9Z6W9pp
axjSgRfvMRBtrGr0F09X5PhO1qmPa+N6Dj0028FD6TDfvkspRFSoXQdVle19nPXH
ge9MQjp1ZZxIkHmI7HG52y2eJ3oqcftzMt4qE9QpthCbywN2yJbTWpqHaAMFqFnD
wGM21rUZIYgXYMy9EkOI9Fvi50WgXOoh/LK0LOJEYYOgjJj+Q+QQLsVFeUIUBhw4
2dBQjZx6lgIzqVArUNvVKBbq7U41oHDtLj5INjWhiB/IXsXTixXmi0rMGPCQcviH
QY0NygrEDmMqj+HOPQuQ+IC7aWwq7Jb7zvluazoTdye9s5jx4kD7bLgC9CHVuHpL
N9sMzhM1yLf6rmNLN2aWjPKgVYs3jvB8TnztfQZlqlbrPkCjMumoDcZ42fb0vlyc
bPlfs3smg75ybLxtAu/59rRuchA/BXxsv4jp+CIIgMU0clDRxEwuUWgWjiAL1zQW
U6fVu4Vx5MNLPfKPVQRhPmhuS2UpiE21Ek6WeI44nAclprT3UDxDboYegEczPeed
sTJQtMfUtq0n0Cty1bYs2k0zrglXvULuukVXNasiaredtgffRprzXeOiPxrLScOt
hTIjikHQM46FAXL/LKgE2+M7KdZ0S5O7IP4R6H9jYtNdPm6SlcUnG3e2WLHfBHgA
ySJtkBbhfth+HMJ2omnLTrArQgmkLHkJBxc8ZPKEeCzib5/1o3mimwd2PBFddxtW
TkkHEM1l2osL1efKM5MRa+qsT8ACQF72dRIiyTHQBzghJd1EgbTQM/jE8hUvw0qj
/g4xm1pY2zMY5fBigWTbD8iRsfYpNR5UULxwZOQ/IaOTgA4Ul7l7Rz1fLx4JqMLf
PoRy3BHi0Q6X2IdqlCaH9X7bZ95Sdf/HZrUh3RXi2b6N62GXDKYG7HQEOnyiAQT2
/8x0NvFleyj1h2cocDOfq8E3Fi1adgYZ+1QrsGY7LCNIXCROhKtTsDe5wJOBcX1D
B95rFsPtQmBi9DadYB7qeaXyvl3tBJAMh1n4UH+ZsylFxK8O3+yQapTVKq7W/BaH
Z0MfstUZuxBXg3iYX99IezCB0A3Z8qdr/5Fr1IkNmRXwU0PqFlcQR9PDooVoAegX
/SuYxh3WA5QtCP4RwT7hTMgHKFf2+TkuGeeKAQ1WavYnOdyQFDDaVuutfp9q6e1p
OTKu/iY+lVRM26BkAzXTjjfTEpxChfUia/Z8S4h+FcvOKDbvrtQARX8/reXPkvGB
jJJT2Q69/dQ8F6wUWHp36lEdR76ODwg0/DTPG3rCyN2yNTv9yZX/GdfKzBHueuAg
iSi7fCBmIf4dQgaw4Igb/fADxwXJLeuHm/AfAoCCkGAFgeda9OaWEZVstjkQjPWd
OodmkppX4TTgvETBBz0OlQMnYMPdJsWg2J7+b2Ye2d2r73G2rOoErvkLRge9wDF7
rlh3LDcpPvP20LguIc2DZjDWXotDL3ux4JNu/KMVwqHS7XJtZUNvrpJaI6ujxspI
uL5ZgUQAHd6XkigP6XUNL+yB5r9sB+3JifOVyISmjXw43ClvZYmbUhqh6Q5oimXF
qLw3YT3x5BNnmy+wFfWcRSF8seb1hciWbktpWRFR5MKOSN75c50c8yENUjhn/BL3
WPX87DctrJj40ssXiXE5qRHs4ipJO5Iu7aulyd07HQLB2gCP4g7fulaR1AswOQDg
+lCd2SJgn4au5ye5789lWTlcQelOkKElD7PvLnFMAE2x5Puq9EHn1yvGHv8Tg6H9
3CzmCQirVpS6B83ZlyTwWXkTbDkYz7L5JJoTUZBhw7MlgwmIzAacpbFwc1OPaYWD
L48ArbN7r4KCGjqEnfujOOzsDH55vioK8cTnt5TpM4tnKJEbFcW3gqFcYsjzdljt
9PlvG4aDJ++6I1ARDzxMM8mpgXWC7lbOs6j36IHR9/qkrTFbLovdVVTmhLC7zLk7
uIux3/fqsW1uQ0mxQ3429fAoGi5grBi/yoWSre7wx05U9xP+7va8fSXXU/TLN9M7
QvBVjhrPiBI/+X7GkspqeFEX8CISOs/+iZxER/ZxIAAbVYrzOwMXEEfAMneepIdj
SBhjakKRJzDwsFDVCOlmOW/IZbq0FvTxsPLpbqAHWyV01MdNJVxc+m6F/U+o28Bg
g+mDmFgRvMZZT+FAxODTV/mNFWIrqopXDjmm3hihj8pIE3rTtQzw482bU7FoB2A4
xG0hS7TKRaZ5XMcRgTHBpdRE7ZFS+cGYvFR4x6HeSmRHp+Y27XQeEC9Os5z2cWdw
esUOk7dyjVH3JDi2clyx8wKMdzVfZCO9it7AAp3pXQAtGiQayF26Hlpg8vLdLPEo
7xo8We4OWyiGD4zOGxFBG8wDYhE4YwZZPSXLm/8Frv5VCfE8rGYN5j52M+OYSvOz
TJMpxJdP/ONm7qCdIXbWFlHSdBoHUKIJFk6mkwt/ZCLKcFFLIZezzBRDDbx6Cg+7
4z4GWNMGBjLK+YFfTEtJv95o/Aaj6BCwfaNzGUmWnNmYhGQFGJcoNhqv06hFDZ9l
W5NwpXuiMmYfXu7ScL1u6gymS4w2KEUwX2Zenyi5K24qyMhAfStbLPLSOkPd14zH
Ew6dSXyEp9F1u9p6y3oEWnA7AGMC0YrCEQtDMYt23BfIXujMtCw1RkifIo8e1reV
WfZ0kqQrQ8HudsHNPwsl5rsLlPp2Izy7gjuLuAXnI9nORfkg4Xr0vW8kTkJvnh8d
Td4gTF2OknlthyuGNpnNKqOKBEFu8uPuLhwRWMCUlcqTKZsnZgcDRaUc48sz3yQ7
kD1KDw81wHYc4uR/n/tfYDskFr2KdB6V3gRR4/V/MEJOVvcLECqGIm3M0SHhraqR
skLN9VUd+6fQCvBJmf7olokfonipURUY7q4ugc7D6V/D6bJhgBcRjAiYMxfCo3LC
VhvedJB291MEXGmrdfszH4g0YmvoNpbm5/nBdLm0puSMZ6Whme1kuKe/QPsdwSjI
P6XqhwzGOMgH+Io+Mgxsu4m6BCkaijnftWzXo3zyKX+WjPJANwo4mmwkexXT0zQk
hmrEtMWjonKmY3KHX45oIjde14futQ5pWyVgns2F2r6A8u9udL8lZSQP5E4UmuTa
Wh9bmjCacEiI/WzxSF/Xm0yZLIbAaQDr7+tKKLZtzIM+HCXcmonXFAbJUo2mjgj4
/0b6AEhbPzUNbVzSSkgEzR2H/2MVmQVHgU2+kzPvPjB5MYockBak6ZHgfTJoP+zm
H8PWPUGa2he5DGyJSof4Wi6YrQ12CLjqfBnu7AGQ8dA0NrycwP6TuNIGY5O+VNP0
A6qEGGdnwhPmhXMVmnYYk9C9heNsOT16+C/uM6SUwe/dbxpoAhbiQqy6wOVjs1KV
TdkvqwvWavjIyLp2oToRiXAfmPTvDhvfKNTbsNVd6np5y/HWwfDbT/77XuOED0U6
PTqv6R5tn5XvzL+MGHzYTCMX4/RGAx65fQZ5M9hvlcliDaCe4Yb4dsRR2pPKj5Sh
zMCZA5S5yw9zbpwsoDNBZkf8XhDowu6gCLoyiLhXzyB+VdVJPRDPk1jgHpsydKHe
vHIVaL7C6/idkgFLBhRn4BCaUKsGHFKwfTbVWQ/wtI/wHPHdFwoyp69eKzgLTM6m
yR8FP18HUzywDF3cTcf+kuNaA3oLeW2LXtZqNCJzmzWmZ2y7mdOEyrvhkSfmSVlD
zUqq7HVpkpyElSKId50N3nNheyPkHgeqJlOJbDM73Z4UY9tRCM3MZwmznNg3Fv48
youZxP13KMNdNz+tK21OPO0R54SoVN8ppsLqIyIw44QO6ZP00UhZ6yBsIhI+0UYs
8dofEX/2ZqnXRfD6X30jwPR43ZpaBYVMtfwBTMa3AfjgyqeBuK0OVvTYqoZMBFu0
RlcycEL41+QG8+2Lz6wKQKVC5q1nZfYvJd3l+A9Nn1Wmpsrd4mig1kLqIAqTK8sh
NfZtQEJh7q9PhXCVBJoAfbgVr0hwAFTyRJwLjSHv2irCu8le/lX8VRS+mD5xbOTn
wBbGEF2AD5a7uCi9KEf0hp8jxE+2r7l7W0r4yHtR3JArK4f5s4xu8k5cmA6A52YA
OHzyTCnct387Cl/lFXeyAHk6jMVYNFe9oVzDrP6Fb2dBm4GufGt6abfTr5NeRshC
//HPUdmLcpSy3Jf88nF/c7rIfC1J88xfex4OB8pM+3xaBSI74AOIlsRSAbvdC6af
+RjnnWZCAMZUMfuZqYS49LEc5oBOtuhpSk1S0itNgd4P5H6yEYIN+b/3XnyHsuwf
t3JLRBd7Dj0eXAteUicQLiBByW//aWOBKdOsBr+btZUyWcbvfYleabJYElvdFtlH
7RmxrYTMr1mmXyR7QuZmsf2rq+sS4csC/cpjcsFUFdeFb7wpEMNX/lTt5gEbeKId
xW1z9mJ5JChdbjczDyImCOfM7yqLIs1gEim03WoW+ZIrrQmURurT3QujSwTD5GDQ
LVkD6XYewB8Sr6pyJ5FtPmEFT0rTd1CPC6u9zLLND7fKIdfyvcUK3XmAKJicrivF
69EnEzzB4UZWQg1HHUMtMhWGh29wcAc3MVF0nc/UEhWgDRx+BrKPxPD29LJO7yO7
1u3DHMumt4HizVf+TkZnLQj2rK7fs7Unx/ea+ug2bY4eSUXhkj7GfGYUqNmiZQX+
jTVEjWvkAU1SvXN3d/cg5DoJfER7r5lpYYRwnh8LMcjOhthTztV1DwsI/SRUvVC1
LFxgbtHBVYEeigjnqKmG5ZW6yYKfe/NGxDB8GTKrUTPN0Sx+nRgqAxkJeLexpWnW
CVhvOfoe2KVdGL92XAreGgLXEam2oQbK3xwrx0SRBVwLdu79HbJz7UKfQJAXqt9p
99R6EqRHUT/RvHNSNG6e6y2VzKxlABKdLlhP8TAQgnW2dUiPhpNXIIELz+ydIi5t
eJmyigO88AnzhfGaxS+zmi9sn9bVb1yKdIiOmNmVJLv5jmN8xaR0R9oKCUX4+0P+
oNjenXPAZd1/nM6UreR/VUjXAo+r9gu02c37a1XbMF7GeVvha4OTorSLGVEczrNV
IR2f5ikSljyqDPlWxQ8cDBmt3yAnp8FmQurL3p2mqfEtROzpjbByU5eKutV48ikD
DXKUqKZnsRjUrM5PfmhC/uqfCcHQwPqFpPqXlOIN4iroEsesPqgwkRxphE+p08PF
7wQKMYlqmtFfwOK43qVuU8d9aFHf4HfQZOVz7q5YUhYL0/GRv/2CUGTR7sOZkmHL
CTsKeJ9ohKGcZaAqHE5Trk8Hc32MyYSJxCdxkKjDPzUVA9GEZ0pEsh1Bcsr65+wi
8iDyacW2lW5Eqb7orEoFczMbsXvcvlC1KXMPpGpDstMdDQZFWzj9JAg/kMpBT2eH
de3wr/+9NxbKR4kdxYNwcnU4ofRxrsbvHyABKf63rK57YxqVEgPT0ZawSLNvsowk
+owFgXP1RzAZV1qpu0PrIIgyaPdKoMRN9ZUuq3fHLEWX3wuQsx3ls0bxJ6eHFLrK
5kzrsrVp/KBs1IgFiaEgWecs1JYDuWDy14VyOuM1Pg/MTuDKNpa91fU7gHH/M9Hi
gmZ+wwrLc/TdVN69jSJduwucPm2ttcCD2x9xXy8gsLf7dLrAg5MvPYftTHlEZ6mA
udYMNqyjbV9in5aDNPg9V61UpfVG7C+xh/w11H4Sc5XMsluPrpxfbbEP22Mf0HIS
kamiF5httSftQmziknMyvVblfGHX2UXzXh2013jxi7qsexbZQ7NHdhc3Li7QDJDA
d1HaSk4Sl2zGBpAJFz0xyeiVWo0/PBqVVGLj3kkSj/W7kkPxPHLv1ztbIr2j09FS
81l2vREbq1TdkW0ugbnsCNhvCk4SZEYQjiKAUl9CHiTdmC261knfTTIY47j+glrB
Z+bb8XPE/ITjthl4iAXKuUPkUP6edgjVNTxmGHe3oTf6QBW9ZVrftKWc2f0F43+Q
ViEmJwi4dZYH+iGsqKLHS0aDI840MK/0a+toY7CmGta9L3eWgVbH+7L9zum2/PoA
p9N5+MQYE0g/7tRINT9fgHESOP9HyR1KFp7tSzd5rOWIk3DiD23wHGAsRp8Eu1qZ
ie93kZXuAxbIQ5nww6h1B42KB1tDZwNzG4hcDnpjPeGMJXhHm29S1JyFqpEmerK7
SaUWd+k2xfQf+oCxtLceu5E2TJPiENklSd/nlf9A+uwBQzD/OC0gbVYpHVWnsVOx
n9GkPwWH4ky6FAfSy0tahcpy0yGYCepCdAv9EyRTMVW8H8WGslzeSi+e0LFRwjCl
IUo/q/zh+xneDsx73+hr5p7arb1VV/ojlW49i9WOoKRr5HHPF7GiHMA7R1ox6uIv
7pIzEroukisgXas4/T7LbuA3zfkiwMHfkemN+1ogZHb2xPYJmMGu4sAI7X0z5A8x
SmBb9wh4C+nc+c8kvNEhJJLddGIF8Id5S2Wwzpnj7G9YHriZShtFQ06vieMSDU8X
ADIIyPvC9cep6/R6xfSW5QIH5WNO2kuWIFyVlLBgwwFL0uUj1vRNY/CzNUGgUq0H
AuxMOFad//Zhrqx2N0Epzg2VYVJFrdcF7tWZ3tUKQEaF5fICcr7sHrCoIm3iEvo9
y3c3ZH5ufj5UAuwlWFnc0icECs2eNMqknfqzS1/tAgqZsksWArPG6QkswwbJQmM7
dl6F+VhfXwCIdOJC9xjaAXM/HVXg/k7pam6PG2GozvQ2a+euR3zTkX9SaBLwiYhd
xTopiYUBeL8MzNBjO2bHZhqtGK75DujPD+Nb+7vSUUo/Xh7MmlpZ/3pu8gUwI+Ui
/A/dzRM4+W5GCbSARD45a0sbaNZMTTxuJN5ekPQtfQOL0N9Uvwrs6kohkso0lv22
/L+A8p99BBLoiuNSxWelrPticId2AQJSGNxyrhXwD2w5VpWhbQQeG7D6ufsLWg9S
JMFqcc0mA3BlFEfuwvs3xPZJVDgQrYK8Lt5p9tTJNrd7ULHpMwPYmn9OVl2vv2t5
d3clLeIMFNR+glwLZOmSWF1fnSisRcqY/mvw6QDXMwZDR/nRGb0vaUFU8Xw/K9bT
9h4CdbBot74eaxNIpZKBtAYqVZQIZcuS2IUSCXmhdAqVjfh4prj3WahfGKKGIdIK
/ESvXMoXekfdCgKjtYwFBXKY1ND+nRu3Kkj1dWpW6tLuNHjyISuOW+sYMsrY3F2L
WvvpE7UopeLND992IVSM8KLkbIlBXKxoekUlEQNXHtxLEQ0DkxxKttnWK1slGWuU
TFiC0ZsFwurZN0J6w/HHmhaUu+2of//XtMGmJcdDLQzWaWOEheY/nv/aMVd7aXg3
JpWKC9VLSfoUAigOFG4FQhg6h5bBXbq4tsZcTsXCseHC7ffXbLdyHroFOHi0txQL
19o3D8s725TjIPkurheSl6HUkxmQF8vkTAwAUB3Mt8oIPk73zeMODjrBYtJxKPkC
Yoq/DCWdrLf/mnAGC8ISbEOgdm4IcSJHzBK1h/HuuTzVOeGqJRJriSuoavVC++Hh
QA5OTp1PitpyXjIOWG0fV9yfR7LUR8UlsvLOdy0evRRPN00ENNLDKfSb8Tk+qYeS
/x5TN6eJDo6zN2YYbjKAwcfZCgL5hLacUdJ4Cdvmj6fwdkPr8jNSmku87llwLJwT
0G98fGfIkCKea5xrc3AMOECCm8LVWIOqklgObbvOtmfgs/UwOWMr3UyNVNQXRHFi
l63gCQpQajI4XK84TskkdC7z50rTmKT0bQvkS8QGcKmhsprKUvQCVob99+KJDQ0C
xpzx4flwtzzs4AKZ0TZB8XBYrvV8KL/V05+HGGm66AxXRAgbQyGImVB07MZEoXgt
prAGEe14HPQj2dIviKX6vVB4UlTMs4M50umKcGrUe7kI0Uy7wmPnJ1TCPH2082DG
M+Inyp+Ofn9E+aYsGdQDvi3npyBpcglNZBm8m1geNe2xuQCDFjl1flQoghNYlU9J
kJgIJZjZ8ShCYOl+9Iz3GQjNorqKiDBlTYQbKHCGHuzQ2ukDNEJtuNODFozLfE1n
VZzOqgUasvXB38vZhAWeKtriH1+vTyjX0JIg/AQH1SBRa1HG6YyDfjXW/wtvuxSV
2HTH3nXx5cfnDC8PYGtSV1aCGOD3Io8IxT/fpQUz0zEoGII40gS2E9oQUucmIkfP
SVwwm+SvjNRYcY9hqbScnfORsnkTggTQRPT71HgVqvel/XM2w3Tpe3ErVQuchXfO
s5Df00lNEC7hz3B8bdhTLEMGF7fZ/61mPWDqyQdOt7Q0QZrTJPFk+m0b+Ayzylmv
+XtELMiZGAHmea2shXeelvtdxO0HM1bjjOVC6RPQOosl1yZO8p6T3KzTL6Y2nhjj
yyJ3A5yWXwN1E0uHw2LgPvGEMoTIL1d+jU9v7tWBaPnYnA9tnyvyDciwKDNtGGMY
2rU7f/deSJuT1TbOHkY055vOXrh+TI1qkr7jOf7b9fnTlat3X25UJcBupPdl3Z8R
j1ujRcDFGKTfrY99Hve5VTOFO47RoOF57ZA/Pu2ZjrMTtlMQlcF41U2EK0ZqLPYe
9ufUlLyAbTgHvSt7CUwaj+63Z1nTuC0Lj9Rq+pvUEt5tgR+KuA8OWzNQ1dVhks1N
zkAZmpB9V7taCYr3QmXjTOvjQrc8Q+8PsYB/QbPUg7ETM8k2JZeLDKr73FZwzaF7
bxX8OiIOiDNZ5MpS2Yu2mjtma7h8yg+MOFoIzUX4uSrCME+qRlPY6t1ndWfJWlks
cWO0JmPk3fOAT+eqaIwI6OAaRHfLW9z2UX0MbYvxfkhXOWMG+KpNFdfDcPzFPkGf
Te1Pxgj/LOOgJN+oWP8yE/85npVz8I8XbTjuGjzg42e7pKun45a3EvFAt5+O6lgv
PuMFOd4UCSs7ktYb2WvuuY539E7L1WUg+2B1345zdAe2e/35206UTGsvKwcIFRG6
ULLejiSjMa/po3sy4sg16xX8SAgINVLcBP5sfVLKfCHblwQTidg68KWaqC1uPA3c
9AyIU1nku26xEBZn0M7Izfur0PNjBeqesZ6Gxy6ibKR8G0i723GnggF2UwYz5Est
uMpBhZJqQzalKrS+58g8cg2LXXc+pMh22JxMcPFiL4RpP+NpDTYKswRFg/s4cBSj
pWe+fo70AJ/R1tu4JjmfbnEk2F/pNOpDYWo9jG1cHOV/O7TJpHnjmwwAya/Uo3Q4
vsX87JTMrI4D9Gb9JqUpnYVfZBhVmuR9dcq3DujLtkQpV2XwvbwYfmQhGe/Ygv11
eTXMCwjDUs5edTpYzqVrHm3NEgzbkcdmcd/T+K6krYVkxCY23bDfpC3EZ+v2FXCF
m7F18zqx8VD+HOerChk5ZXHgDbQljdHt8iO1YqH7O6hEZNCp/vkzUaBWT9RUGDKh
LFKy6M6ea9JEYiaS9fhFLLZVBPMRb+ZRdzMsY99Fn8fPMRtqdx0DHofu7IaamI0P
jG0dxjJwOWLz0eBzvpIllNbqWzObOvNy2yndEHlq/sMov5Zmlwttd9QNCBMIpz2O
86p5LCwQClmn+21dndDq629tQ1+Rx8QOASvlSxyBt143gc27yV3nQnWiYMKZQVbI
ypVj6qtVhBEwJyvKqV08KgNI1TdGuCgdOMUbRehFmHMOKUhGNhwwIWpmPLHGijAS
JuDMpVHq8wFcHxPrZz9EIzzj6FGAT53JlBdXQhUpnhil6XceLL18vV7D9TdqrAz0
F5WeIY29qgZOI5Xv5BisBRkkY55IqOb8XxcEyNcVT1SFg7K+EQAqDBnz8P/el8Vb
QwbQZaoPRxwz10MoNkTB2l295og80ruxyZKnXLpj1jM0tfJQjmEmbEUFmhAvx30Q
kiC4tBlevwvEiFqKucIf2BtNZj4g3wbLk+ocg6mi/XDx6sIk+6uP7XGKfhTQAmEV
kLTgHbYcMT8uYz7Y4GvAE/7YuIENG3La+VFKXYwIm3sGjL+NENbmoWy2b76PLHdZ
+e9bFN0qlvdXcQXbThTxgpiUuuI/3Viqi28F3LAAovlfz8Wunq+6bQrOrfkXGK4g
dUovjW+YMk8XIFW8/x4YBBqOtSzxHPS/VT8dE54S0kFpwUNVDhJhNIQFglhzBbjX
l8gr7xuI4ULmHLE245PKP3gbW1vtt6p6oCEbG+C8uMmzhTFhFA+oH/gHANKvYkcY
ptAQU+a/tHEn7RENKn3Nxsm3oOQNClaXpvjx3PXv42d2o9btmf3Ueb3GyUFMhfMC
6yqQmbAJuzfo/Ze+/YEwax9Bn1DaQ1UHfjd1hBqUMFyLTprShGPkhM8dGoJDiSjs
hwQTkWH1ToHi7k+esEvC4LpVoZLw94Y+pyWZX0SWH6GxSqJgE3wWkqrUMiBD3kzP
Ydu/6peT5Xl5M8JhxTyxIPLiH5yKtmy8YZPjGP2kbleStPlaPtL05ZwT9QYZX5zG
vp1pEPp1PvQpxNa9B6D87b1ODEhtAwyNT+q35tMLgWFEgkCeZarstnaWoHFG6QFu
7GEEPJZ5Ya0nj7+zxiKG3zE9c/Zte+UzLPv6NstzoDm1+/e9xI4ruNmhbPxPNIWL
43h9tpbNIIn+UvisLxEcFcWrMMOlqnO/OSd/pyL/lLSidUgD+qkOwelO7V0/GRTe
hVgOWYe4VYHZpeGNw3CRcMl3TN37MFwUwOLr8qnrE+xblwUsqqIgXPOofjHZpnlP
8CTCkNkOCPyKOZfvLbftdLyM7SlMDD/y9C92N2JmOKRLJT2S7UE7pbrnYmj/Wm6b
B8gGEeABtNF+X8K29x3t+CsXD6OweEvSTCBLxX2Hvf8Q0/Wlr+nkI9h3sBvO8Bh6
cmdd02/HvvPgyGIJaPer2mWBFN50UlxFFlaazOY5fdauZVDEj5v+Agpi/x7CLNIo
7W6QZ36ZrSpHAOgvxI7jQEbFOgMkXP+NKofsSa4ixSJKCoz0s0ogN7yHq05+Gj2/
e7E1b6AFilVRf0aXRYQUF4xG9L6wtYACwwVWkb2zdrl3CCuefyQIwgKdowIKwZer
lB38Ef64QzbH+N1H2NDWvqXf5a11KAv6HG88feEdIOQq9Zmd3GQX9DYk0DubvgVa
kT9nlUFGv/9PgHgzQ8D3tuhIEL/tUaQnNmsXx9pJXM2ev7RlLpGmKWK7PG16BZEB
ntDrTjC4z8RMrsscyMqXxSlqoy0Lq9NlintkxaF+u7yak8XKxXXT6yYpT0XWM84x
U/WcOi5Ajzqq3MRsResyqVr534VhSy6Uu3pyMkKVUcLtYiZyqBREPNOy+Alr65Lm
t67GMvzKNVnTUcpgxgS0dfLF+T84CKqBRPEav4t4JjIt6VJzIFfRagJzEskDP4j+
F/sQ3nBJ1mA7D1avfTLelnVbGumrrmv/Rx/SlcmM+OHOAys6mRpLyaCY30ajYEdk
UDkgBT/raOfLyueGw13xxPsOH7FPuoIbV7F0qgE+wjTHDH9EOgJ7WpkbWSva8xDh
cwjQvANTpTymCyEdUdhQWgP5PzKzU8Ic66vcDTiv9rb24sBm23nX77Yy8DKqXtCT
N9layRHBlWg5SESTPp+MKV3w11wjPDTQpenQ+QCsNeeijUAZ1QFveMidDB2l0Dfx
rmdUWjDN8UV7wZDLpcWuOxxVdGktHCOyY2Eg7xVguo4asR4rkYzsHpYbzQlX6YAK
W7xCJVRErgePbuYTMwsndZpzO8Jh/ls7C696JvEQLKc4kHJW+hHkaLzL61E1Z1Ic
3KX5EXJfhgHCQ7RHXQpdb/9QjepVr/icBaM4GFcvkWUg9XYlMseQYZgjp0tfbJA4
Uvqzk7hSiacv+jNy9DYHjaEAvQIaIZOJ8VsD6zGdHbL+7LyRdpyS7cszFP6Drl2O
tCP8CMHZZJ7BEU5djUwpv3aWe2CePzIbx3qQOY3LuwJPoBSn1fy9/JvNKjLoakx7
EwjgLaSTPE8A4hsg0yUgzZg0vEPL+a6g2lCTNcrK7AVX3WWaZ6wf2qCTv9ZsC5AZ
ohV4OclIhvhToJQUNkGc44oLth8DNTEyhp7hXczI8kVE3vQ1C4gM3ZSezeSwGhCO
tuKJnyma7a6ihNfvxcNP6i8bbIr91TQUpoHFS22Wf0H9yAajXUn5pM1Onaskg/4K
VSGDyY5T+51mwHkfMetpxDVBuMSyuPgJksDWLhRKweQZFZBrY5yq+qU6J0Nv0UHz
secp9bC2KNzMVFMRDb+dN5cm4PmGTnJauhHWX+hmTsk+XzXOmJFDJfVDa65v64lW
bv4H+Z77LtqNANR7Cr5Jodnpx7iMbdnGmHlOmuAn63emN6d+mRHnaileu2Wn84nJ
iqgSUXrTiJH30AZc3MaFars8uoF6A2FOqymJLrIcPfGCgKiQgVTeps31q7UEwgZP
Mt19vdscbtfLH/YIYDKFk28ScEwlrbmSPuZnztnyDqGV52wxL8opCGkx85GsOFU4
05J2RWYDjfogLMlne97KKewF/LrqfoC++OmeaKZWhTOpy6pahCIYdCJohsJcuii3
SBAA7KQBE28PNijCnRcWxWFVdy91iaJDvmNcmq3ipLGdNfUgtuYErDj+0R6KIo+Q
nMm9Thu4LYZtJzp2mKp5h2XX3NOJNA5vzo1ZaKsl1mbwGanxnVJA3sXLzOVIUd+v
pA6UaQXgOnTUcJgo2pvBBJlXIb3SpvzmIiCaJuXi7y0e7LgiiGAPCGND+KrNX7oi
HqQS7g80EvWzlXzX891cvDtmyw78AWIt5H43TQITTutSRjrH8Xkdsqai+qRKG4fz
/AlcORPKcNdTn2U9+CUzqSpjuBmvFH2M6S0GkHWbUXnPgeXgFcydL99VtKwMUG9u
ak6cNgVAD3Vw1Rz4Fx+uCTwq0ym2DUGS0DHdL9k7SgUKvQHVIFz6CD8Ev13RI6yR
aAnAJx/5aBnx1BVxUL3o7DjE6U26n1mMtx6pUxaOnrK8EmozTKLEkkfp8y2ub6P6
dg5qIzL/3XWDN1MgzCjds0fgUjd7RlKXVfoJp1gjeZX+mIC0MckWulCd707W73MB
E0Y4fjWygr9exCIyj9IckYnTRmzbC9lbh/pd95FxxdlSnkFKzxXxwGzDXBv4aReC
p+BsBv8rmLbSSfdAJ96yHAqdVAXLezgUgpqQMNbO1pL2O5bjS2NK/eSSdcGIfVMp
kZiiCvHImr90lRG2jYeWlnONsCvQRmtUM5OX9Et/5ZFqD4GdiIJUlnEW/TB7GEUk
bLGxJyL32wBqMmzlcFolN/xZFYU5xseSmIeRpTZ8WQ/MzF2BOnTwJkrp/3v5g7/O
PM1R72EJag8JMiCvYawM4euLCTHsksxPs29+fuKj4ZAC/kc1f9GyzX/q+7MBtdyl
bF01rbZoGjrzeSe/Od8mgGdtR5YP8afYHkLhlHmmQ7L8yQhN9XmTiO2ITDQrWziW
lB753Tj2oeVAeYvib8dsAHVDqEscDsRe71viTZr+iAHA+4/IHuFjPNidxy4+05FL
BolCmOmIqDaD5oKyuRz+Vvp8K5q9dHPLtXxHCxidLJcoAXbfM/rJ5uzf+TnArs7N
ciCL0eiMeqwFEwwZlsg2IRSfwHI4JREl4p9wUoh7VPl7nFoNugN/IOnAmIyUawkN
ZlHAJ7rCDpWXsehLXpcPsS7C97sTrx9VTYm4u+AwJgZODUS5eQLFVP4DvA4aFAhP
zdPHYZYP1v3X0CqfUWXs6kSECydzwHVTyiVCFMjZYLHf+BaEOqx2GmzRaVVJ4rEJ
yGNudVax/qdWRVasvLLgEGH/IMgYCLbJFtGuorkq1r4fH2U0DVdnUQX6YhN42fZJ
23Kij/qS5OLgo0GJaidTqkd9wWZzWEvYms0YvEgFk7gs3WKQrttK+qKgi2mNNssk
bmHbrVtX6lNdVgwosmEAyxfUtnN6NMS3IC0eSTwsli58T6p20CrCxlG7zkHp1JSX
qzHmmuZZQfBe4w1CTU87NVre4VqIQTHLuAYN9wBVImkOoZFXFB/KzDwyEesGtpFv
IsxyA5zPvxrTQ1U5bUD7MprQX2IzF6HqOPYY80jGUx4ITwEbPQRRfL7APhkTzl6C
aybiMeIDCIFBWF9Re7rSebmRhFQp9mo/3hYKXh7hxRGUwq+djSPmGsrSZbL9mbNj
0/YOKqTj2/kwjb/D43QzTWuViutaKso1FH3zQwoqMXb6QaAAVF9Uor10tHFCjiAJ
wi6okeECH/5tMjJv1WAzQ9rt2hN1pjSaRTw8zd88vh6heIIrohvgjLWUDU116+d+
uPe/q1Inv+Y8gNOm7AW1fxKX3rFHGP1KXpC4b/BzK+7bXipZGyQ3WZDqAzheRg+b
HvJzjlmvrColBiw9ICBa21Uz31kvk5KKI/vPuhaKI19zWYHxjIl9ARlOxhASPeer
z3VqaWHbMbDTAJlrjEOhYCj6pRAU+Q8Rr+Mfmf3ljKHH60qZtLekmmjrwj2RwhLn
T4tqfHuzbzwk1OOKzrBUR2aqEDZD40/U0qmlyStnSQCGlxX9MSaJTvdMeO/7MTk+
oFMB/R2rvWwSfBh6NnnPIqY8BjwutaTBybNTz5sq4aub5mrBE8BEjY0ydjqyLwlD
bXpIlF1YhgwRzTHESzUsOo4KBwTyp3pTjlm9MWUeIVEA/7hYRMGRRPDrBRVGXm6T
cyUC2SSOmKLVDC1jIifv/msxO68GbfHHa5cqPa71Gv8J9cE+Ae79FR9kW2hiiP9M
XnMNrsx6qMFjRlXKYPv+fohhTSovqR/h7iPmsQ/yFZBAn8El9tmwCu74J6Rz0tHG
ZT2pSSyNF0COQ/CgcTjn0XMmCmQ0u3kdhyPlqNz6Ccl0ReGEHVXvvGjGOaXpYOjO
wssNUjXZqh7v/tMBLq5wP7V5JUFzS1B9VDYOYCkPF8roKFk+ZeHebRNMg+8fFAT3
XV5bx5DCIXb4G973hQMhXRhdUJNIMrdUk4i+/n6FNj7LX7BO8j56ziDOPQcBtKfj
HCGhTK3ZeB3m7qlMm9EY1L9L9BPfQ0vvPzy7NPwhcfvLC1D5ExlpXF4bWCA5YRlu
zLKMaQ8YNKSREtxhr3fcecrAHgmB9mvtYVUekHWLmeaHBPhFObPjuUWaQzRl3L9l
UWQncBwmThNHpnGPjPvEVNlNQ0jLvuBiYxfTS1XG2jqFIj26fDWSO3xQz1vDwLeZ
CnA5eU3pzXhdgDCe1BuoOhDM9EkHk124HDR8CPwI7Vn7zD/JxPC1gAGFa9mzcu9e
a6tAYkC2A1jj6VlBYMyTWSgPfpMdJa6Eu64/nXm/2hC+gJNb0BZYvCFU0x8jmlMY
vW6SECg4rJx0DPVHkOBYXhuoLNMQEWQfHPgiAlRLygj7g54n6S967vlVTYerJS03
d35ZZGyUwQBBgUjwgWsukqhUaDZxJZCN91iSKFW+KXv0+SChAcmUhYl5LniRRhnx
kLdWPVf7eduoo+D2qynszYGSCwiSqBn7Q1tI4Vpqlu1k5aHI3AI5nXhVmIhK3Ldc
2EQfUUGN4/k7B7xCT5fSP+75Yn8BP6BbHz/BBS5SqpYZTuQ7TXyFyyk564HpRtOh
JwMEezfo6p7ZHXwzfojHpzTGnax5l1EaSMhSMPAjMg7YU8b+7VE2U7OgK8rci1W0
9Sw86vJnVhVqLMxNYVUIPF/Ll0xME8ZQu4hDWQyDrg7KZ8Ow/HS3TKgKnjdq/ah/
lksA0oiAKCK88AXeQOcIsRNCyIMX5ShmbrHTZ6lu2Bzsq8cia7jLF+GxmKijK0OK
0qnwbergcXgW5iOfFO9pzeu7Wdy1hcMhP4szw67AqynuMhOi/G8BQGkJ0snDRK6Y
lYbiumksAtnTb5XR6txlezkTM945sic8E8YSZJbxkEzJYCeOJSisoSRpBYw0Z2rS
63TR0hSXxVmn4pJubGquDGnIGsIH4njPCWNo8KELGHwOVWlWoUkudLlDweXJZbiZ
U3QMS6mWpUqIAxNR0TdGijuLmBD4hwp5Gbxh+zChPNBDfVm0IGbC55SZKvrACXEh
4j3m+TYaBZR1HEzSwIZgxaNkK2+2qxF49dTnayURzM/3jkFMWES41lkZLNeO+60V
YTXwMzFRQkjkY9dTESy7ElpcBmTgPuNcc4j5LN9BL7BqlpySFraMSyZhu9ME7lr1
eE06H4LhEDTUPWFPBbht5ulZjjfDHqdgdl004pRkuvzB534ma5iMXzrzq41POco2
UFLqakn2+eUHt2M7H2NtTAkvFwmbKYfna6a1j1JQAedMV253xgn/Skexy4xLsfoI
rZbmbMYNZzI2dypwqNKML63Ds+g1phBvwiy2s/XR6fS19LKs8FB4zy3QiMUu2qXl
ublLoP1OVPJKJn7iDLAWHiQZpsD4prkPdARR3N1rsh6VUPwnulmprKJ/DTUuKZIA
Lg6nSqOGYDML7RMuKeF4/28lnk+yufA6O60M9MtTlLSQiWoSzalx4+2uVBBmfSdS
q8lV/qj5aAiUneLjLHGAFsnlCd7fmx6y5kjlFblg5fQEdRAcNcatNWsd4jeN7lUd
UisInJdduxaVg5fpt1Qof5Wa5tQWfrBOS+5W3CqcTZ4BUmTrrbLYzrf9fB54Hnbo
H1TXb51B2ZinpWbjVHpOCb6Wtfo+5cbUhJJ87/ZjthddMHGk55ZhW5CROmmbZd9K
w2Fo++1R1key/c+2ABrnRcFd2hUaDBX6VYLCrFeehhEx/yhq7Iugi2jVCuG9vsq5
z7+9U5/gjpoW3lajRzgCpsy0w8jkJ9DG/80OK4lH7iE0+GoSAP4ciNgzBUpOC/3o
Qg/EGn+9941O0vDW8s4szKonm2ox6DmxtEV+bx2Jz/1W+guAmSQzfteoJoNh3IVl
0enXmDM2v3s4GYS1eYQJ2APqKu3msOCVDGWFTXAmgr4ZHUNenp/wEhWCB2pcFRU1
Bgd/IdA+c3dUW+E/prg1ArNrHblvZwvZbi2qjVPsfMUVGAlacSbwzVuNAwSTyY1b
U6cLp10wPVSeoYqHnyfsu0sYZy9eLrOGEUZqTWH04xcPXTp89PLdZhf4NqqihG4o
bb0YJAKPhfdyjiIGkZT36cLnKx1vCNAhzisSZY+8GzSdGad0MijPc1RBsS8+5YAk
JcUnLJ11QC0IUXWTnxE+7/8IUaNoM/90Q8BxDkSN2Vojl51Y8rwki1HSrDpIirWP
Jwhqw7jioziPsKQoUrpo6IJg1j0xJ44DZtqMoOii+e9IfP+NcnYje7ihIu21JNlT
Ei4rfO3vDmTcKAUJEncp/PJKqZVfhEePQkeUw/q81AIC6eSnAfGZZaIL30/0XlA0
3yJR4Hs1S1Vrx/p3IbmYje125bvm//nXAnjKs5zQX59rxETrWvYZwLtExnTytlcR
3qICbuV9CX+EFBd6g5Dotu9t7WTD0rjv18sUNqL9WtGsIVfDoIlj6KkWLRSkZBCv
xTWtxgQ7G2s1h+KS7BhQdU4D8p8lWRQvV7FlFARgf1kkaFgGbeLJiodQO8Z3GIqh
VBvIDQYqY1FN1TXMSZRgbSknOrFORPTGpN+gtTwoxp2ZPw6oWVNFWluUdt5dhvbl
hgLFrttP4prm3Szt2KXTVBLNqYSElfQUJMvWCVLj9HpVilUT79AnWpdhpgtgijTf
JVDSo7M1IivW8xmR77SWcZR+Vn6uE+yxJZdZcnXFahmmIG3zYv+XIqY8kDHLPhPF
1032ar9oeBy4WShSlIGjZflghhSCs2gIgnEbwFKgB/PNuDT8W0yjXEZJ9eBX2bko
jSQ3ofTelv26S6B18ev8ROx0WLva7kG/4oUxsgZ3Qb5Z5KkF7NGoQL2bKFRspaIo
rn2rUgzyFMlcBRjK6h7E4CjhEuCJu4kODztWnewf8ZBW3jJXFhz5zrum9TavEzJT
sECygg+mkeC1dMK+X1xLDel/IiA0PGA8jU6rP8NDSERLsQ4D8mZFzNmSTSLBiZ4T
aOj+ZOhtIeBjKESc1IWlJ2c9uDyLRBwPpSLSyVaMoDd+zgxzTX1J+jsijDJ6TOKE
qcqer2J9XTVHzPcKOAMOWfqlxEDNnAVKCglDUStm7Qq/Ahzp1ybledxpbuUaEWfW
gkbjv2dBJfj0Ri2lynVIAtLuxUqenSKYsam+3cikwHCrI7wDW1Uyrmk2zZFKQSgB
ulrbyt5/Eb+TbSd+7/DRg5tEpaRmfQND+hWiidEGFh14s56Vzv76II18uMrbv06C
iePU5JC5o9sWtwu/jXtpEWJyLAY+mRntbGP6EwOJSpfvaQ3RbBG3xeNAlc4ApVCC
GYPTH9I/GlLM0UyKquebS2DP+qYOuEyrNzbKNvnLURkkohB7jszWm4VrpWOcKIEM
YzgAceB7nhL9ZB/eueyJnqdEE4LtLUkDo7OzA8SBNFixs+FutZBzh5ZodfuuPv7X
ITh0c0OXbSkzvpKauoYFzL6n96MZCepJ4EkS13qNnp/X6ntp1f8UyPACMNg8gV3V
pj9AQEmeVgVmOjheputTWLddEzMNLjd5HJkLXVkNuAlMSHWkAZm5PrU7xLRLc3dd
OsS5v/jp4ciYvCwrMVeGls8UqmCqdAlVZkH/ZDtDmfXb0LjINCgUVDyHaKWGheKw
eeFeZfsP/zZMAh+5GSRawvpQdppoR1edGjWznhGMIVvgTt78LwtZWFl5pYkw/ErX
aY89IXn6BElV0cNCqkuqWguaGUfsIhcLIQ/iBYe41BJ79ujKFFAtcX3QK7+s2QtU
evsB7GYniF0tzLwDUz3RaE3dUFZODRZjgSg/2TYs8QSNA3N/V56SQX4Jmkxzn8DB
b0fWGhNKu9yIiZUtAE8VRoxeosw4Mn8EZnbaeCBoEYMrRCQRZsc3mqr2V26ZeTe0
advbmnwPCpg7aV0VLQoQMBS7c+Cwfjk0EHEC20vb+kuitkw8wOV5Ke5XsbKcFZwX
BK4KpDvSZy4ODlVP47ZFm49pUixVOMiqutomEq7A5J2x52Y5pD6T4KzPk0J2qvuK
xFHCljVLEtP3bQfLTRdeETVRJg6hbEc3rr35OMhiPSEva3XXCqIY7mc3/D8fOFPY
GAw2Ou/rHj5TjWzrtHY+Mfq+XT4FlmoN44VUcp3nbzlxsFuirSxxOkeQaRgwu9mz
eb3r7cElGTAJxkUJTzv1DCfl4OcEl/qOC4nVZaCC/5LTQqlRWhju3fn2okIG+Xdh
RtGBgOlzj0XXAxmzIUVSUVIDfrLlZ6zUVinad0QL7xwoDF1wQ5xZzFppaVJCTfp2
WtKykwWp5cMV5/aJK6NtG9vqKbf6x6HvmO86TmY9DWI8hzn4Dkc7K7a4iPAqsypQ
skJpTNFRoXb5AwZNKxzYVdp/mhMURcuAhprsFetWBCbPNBA+7RO4vX0oU1EDcIub
aD6V545FCZwVPW9TOmXAbxFQK1GduGLqxQ9vqcC6k9SCfPJg8DeoWAT9u4wmosuD
uLgmxxpwvtL9NhNFMpp+wO5bdQFgcPa4+tMmTZBlhvbjBZph8hWfELWOnZ/MKCPv
tMHTTi3zF9ZWYnx2gz2DhZEbqmfky170oadjLlqeQLR72MiUEc672S+ZVtbMyBoj
i9gyVWU4EufIdYAuAiNhpVy6Oq1ozS805rMA8/Tw5PdHV0pxAegYRV6AOu/ukvJf
KxKlkik/OxdjMqhYYXcxfivkzRs+rX73TPbzCLx1nSoy5HukznrL9AAxCNMnKIVI
yw12kQJBUtBhcAd+BcWs4/PLlbDU9PKyDuROiXDau56gd0/TTBs+DyqyAhAu+E44
dutE/FXswdHr4JE2JJeVSNQYfRlR9I15Lw6UuCGmEsU2Q3oZFKmWw5v74T3K19N9
qK48hCrXBNzl5evvgzuKCglxgkvm0XMvKebdeXphEREnvHwtfY4dH4JUVo+XZ1r9
ZPNxkHjvxPUXoNcsBudfGrkmepdgXB4/Pfq3tkB9LiMKJcj/qzPLSgvaGH8s3QpT
FdXRMbfbXNhtwCec2w9atcUgv3BBqYzbUfIHkvaASn1Cz7PO37LnSwYjJ8BczQJS
0nvnsASJHdxrcxv/qxpym+1GWWKZl+w7u0LSgsDvFgu02ex2409qjt/rC6nzmey8
xj2whbCFUNx2apY8yhPlMJtCUbuDz9IrD7fwpp/DlQavGpHI4LDZDO9oEqTxG1Cz
ItV0MKNarvoeWK1hmJrvZPAcR+rvkSHxXGEQsiQ2y8H4VlJ2IyNytbUXcZJqaXUR
zdZprGztHUo5goYTT7OWS2miHF/SXohGZL8ayy/kLMkz4FO6n6zEGelCeOLdljrr
NBtygT8BiWenjeFL9xdxvKEtC2IK8jgLqjPwflMO2wL+l/LMSFd4l1loyH75NJhc
Jng2gtSoEsT9LYAGK672mR3xhLgGmStcmpdQ3Ql2LIuTjXaJEJD2+UNN++tPQsll
wzFizrE1o3R8EeMIQ7sCbTYd5FyuRKXU8+ozSZVTGyWy2BBTlk8u9hZiTaXs6k1n
x864a+H3XoayuFFclU3Ngd3v/LG6tUNJiAbTJDOJZw+VBUuuNg+213ufOJtK3BaC
8cxDMPYI6SDgT/CmSjeQyYQAE1q5WXi23hMjCwXUQDk3T32ImAIe9a4LTzNJF8WG
iWpAyXCBGswPKp0jVgsSqiPTjx8gJUHa1yDQXubKsoVCKPxAu2tPlfw7Ppc3FyZe
tLWO00w/6HD3u6YX0dkZgkNb9YAO03KEjJ5mumPDYb+uxiA1f9WPBpAorBDns+Qt
Gjz34xa0BlUBbpOs9aBUvkNkAYabCyCkBqy3aHi2AdHGwXtdf8YBTExkJ+Be8NlN
t9SdBr+8k/kYzLllqVZbYWXUbZrVSwJ84fxIHSkx+yT5LimZBhZEuJf5lhPd7iof
e/P5+zWz3tIOAbtx9qWqt04OFVL6ROKQM882+Lvx0danisEK6uXfl6gndAqhUObY
yKdzYr3QJgohOwZcVdJ94FDFTSQdWoWCP7uTADDcnhMZTTGJoJgnQEJ8fqqRwAkU
qedb5UkFib0tG+ugEB5Gy6l2brYuc3ayXDDUcEXStz/eIQcSpB/yyVdWW8/xQYl6
VKJif7snSKx1UXb078lJLnjEWQcpaOGyxv2kA65Kdk7EgYQJEAxQZQG/9ZyMDIvy
u5o4t1HNRRN34QfqnHC2YWSCvQuI2AAbGVLBiQll76xRywbEYg5NVB+heuGDDcOW
8dAN9+6/921YqXxc2G0fjrSIvJJSw6vJSzPOt5jLeHDLAmrni/wQWMZjeurjNz1R
HxGaUJUIeCK/K7UEh17tkxl+/24eIwHCvRG3ZrxE8em2o/nld+L2J7462TZsL6aU
jTGc4Tt32IAD2Z6IqmXhdefnl0n/5kAh4W11na/XrF0XdBcs1yQ9VbWPWTS+x+Qw
95UK05ICwUFXUffiGT+CyisCytYpPsOaFh4y7L6CaTa8sZuGzgZn3GhUOZj9K318
k4Nn3oInVhRbUBCCzQ9HtYdnQKk+gdbELZvTBj6AaeTnMEQwFk3AvOljvylpXqXS
rlFpk8wEjcIlICVEyaqzBNYR1lB+MeUwwW2A5GiqSVrLd0WawSgqYW7IMZuV7jPS
I/hVNiOzTO7mRmTKOzTK5RhGNn1kOeGUY6Vim9UtJO+HsY95Nrv4aBUX2SciBWQr
yFMhwDCZUKxh7d6hFz4aEj/inKxtNDjhRza2qERk/FyiraTLwgmpTCmivoPM2uMC
999vPvpxyaHx1UBRC6STYt6RaUsgQDfmcolJ4JYv1Sa/vSNvrDfsT/Zi0wBRcwZC
He2lKsVmaFPMi7irE7NiSsl+n8/9jw7Bod7BH+kTV5AcZa1OLut4iLuwCwBvC/+3
pC7rDs3pzW0W5ouyKLN3SUijo+L0VL4qKTj+jm6VbqzJQCC9QdSrdvVWV+APRgf2
S7qGxahvm0R73bnMH7W5JqbyZwsyjOo28iv3ZwxUxvRUmZ8oi2mA0bt6fvc3Scto
0xTqNJonUfxY+B123mMuWi6QvPwlkHGvNzmoLH8UhJOTg68lR4YS1ZbDEn1uQb8k
FrC6LooBSGk4XjjiFYkwMPuHWCNdoBPwXDwU+eiMmOmgXelWDQY9bB35tmkD/Vga
E1ZiL0PXO5R+3koKF0OYdw+0m8t/BYkJU06pRkz86aFa187KDO93BfXh+DGmXvTp
rdkc13LO8k+esdlgWF8/J+Ug2yPunKkSPbwhyzf7vR1HmfX5yOJy7rRRW1Nm4bH6
lqNfZG9jsbTi9HbQ5N67vzKC91db3fStG59CzA8KMSYz52bJsIqMUjI8naZJqZRM
XOsiFr5MeW8OnF5ihetLHG5xqdA21xxJDuMzQaxSRqfL4EYLRipsQ8QWUBmiuOa3
WNi8YO9t55LqppMWWqfFz8kWTb/TpwdwThQK1yBuzJwae+kFbXB2/MkYHsJoxV8u
bGOjneW6Xk1HFQUMuMUoO3FOcGsXwKhpOzxehcQZJTYVF9pLOilyTe+PwKLWfadu
gqTQitNmdgAtnroKe7Y1RJcgykR3LMriqqqZ0QgRCUTibsQFS2DzRueRBuJ3S7q3
sJOZ7ZinUI4QbKxNL5TFm8uuX/+tftYJOMkIkSv0Wt8cwpDdUFF0oJFFThCOXnbx
nFvItAiQkmuhpRgR3X4DeYKVrIEgnj62D600LkTgZYuW/akD5lS644+dgen35ksM
5DUSCAbbvb7m/MLaA/ukIMJcj5oStDwg/Eo6/FXlopYrmJwifTxZfDQfHl8C0PJr
Q4kze4ZWmWNJIFvAhW5+HnqigfijyeWI+8B/vSF5LICnim9d4oYz0DZvdiOdJGxA
uu+33RiyZsXbBY7SIfeXTdRVL+dronuF3vn4pJYdfvRYMrdk1VJiqyX6M0x9/CiQ
gDib2UD/d7p4sASV7k0nfCUEn7wncO188DTFm9eziIsXVGnL6/twnXQ8JzglO36R
WKvCEfnfiwy0o5FD3uOhX182jwoEI9btaTbOADxKuw/0kXSi6jZIc1iJrV8CMVis
KI+USNxzcrfEUSxIWTsasxaEqGyR+MgD/0h5NL/Dcnx+2NWeULFU/JTKsAGjeeGz
wDp8QN9Q7Logmf8jpA8sCaA1UxLqLMmkxYgeQYpv3JxalSZb8Grib6EKGGKd5k6l
CnCmzL6bJpnHKJo73rpPWA3CQl3IAksp9925vhhD7eqaWB76tyVpo9aDpJnIjDnS
JoeZ78/GSokQXFZCHrx9z6ucXW9fPwKYpMYRVkO9UFUCX/24z/bB1aVLipOd6ioC
ienUIT8vtt63tmehwQV8rLFVBXeedB4va2LQ0O78OggIRWwswLaZItTDcn+5cYyb
mHio3vTwZlgh8qqxQu+in8eRLQqkYAPBlumqhghJODGkI8RUPtCr86QNepvSTlPR
WBEIGAC+zkXnT44ohBtas7QwP4SsV0+tiMfiIf+/E9TUGU4z27EaLZ7GDntvyZMk
axbsEvTPc7ULqu4BK32Qs1Xz74hOHKEaDcRkwcKjLvbP4zHlZbNbX5xFCmA/lz9Q
MzXDOEfrBpKgugYWgbricVbcdmBUTVKuPXPQ5d6jR4ptnB6guUo4sRo91++ApNwW
/9siHTuMItlmzvdtNQJe3LZQdeRaSGhAKN8YNSGRmAkujXaKXoeNd1rPPhToVQkF
oUlzoVIX4fOfzJYPpgOxf8nlvhJe3EiJ0ksT5uFkNEWcf2X17u2O16Q89e1CttQC
Ixzt7IWi5FqqQOylI942Out4chKAXsFhjsbt5M3rZNs6t1O5KkTCPCtRnY7njU1j
fjja8AbWr+C5b5q2FzfZHHszKQGD9Wq2WMAwlobCNJjgw6Q/zE7/b7U78m85v91A
8ScmmQfZYWeACehxnTBv64NFjjTPk+i5QrPZrkTwn8c0RE4y0brFPs3djOhlJ1jA
gFIlpwBpDme+2FzKeKRzlnQEdKxzB+1GSiV/Kl3/3ZF3QfYwXIdSDH+IIdc7Ecti
Rlvr9i03F4Ytcs7y9wFphW/WoVfAy393C26LU84RRQjGkS47yfC0XdPyWz90Hw1h
cDnYQQFqNNYM95B7UbKplcZtBqwcXQkXxgUvdrpKpkn0jUOgsJiU55TZj9RECa6x
3kaBr5eDJCSS5/e03Winipq1lfU8CYcUgCBlXpcZzXUjzs1szQ1/fbD+00k4rtLI
v1sFIrW+7wrvBTMDv3b22uwFxzLCqNX/as5gGhE2Kq0bE/M5SFD8u9LIi8GJtZ9i
zoGlnKx/H7uTipRSG97u7utnoRKxLOg5uel3Sub5R9DXkubM5rpT7gCHjhUTs99b
7ae9OpAxpHstb9uMyVFPGaz+qlUz1QKUWSMvUy7qPvD7lTQfMn0MYFcERBSHPWCX
3xY/AMPrPSrm442EiVCD+Q4+DqazC5q9MiQXyw7pKplol90R12Z6+zbol1cofj9+
3TuyW0bp00LjfKpcCFPopAc1sc4aBbvG2WYtUMYZYaGL+JoDSP4NVsM2L663qbeQ
J5EN8JZwtfYwiR6ibn3bbaQAEcKgeSlpKF4Vlrw5BpLzqI0Odehg1iZPca/wSGPh
o7Vj0hX7iu1qbgXP8Uf0oY67Ls4FzyXEtYb8H2c6uUCcTNOr2uLJZosFpscGTzW6
hRYM/n3F61f19fM0kfKUvk2o/RXO7A6AUfIlPTL+IduamARpmJulZeLvdKgvx6sB
4xnj7ubVOOZMjK/wSvogmxE1dEdp/E3bmWPukuWMNubOYqenPP8EyzsWnwztaDn6
ewHU5HipFon7p/MhnuAwX0LVIYurEnNbUEyRpsKAO5Z6mNht6hKfQDLueA6btd1q
jzQ57GxfBGXGwBDcqCRrhm/dHWPYANQMJgDaNwN1+lDIks/LzNVkDGnx1uRoHxTI
Ox1bdUNjXPDaQIFGssklGS2lqVJ8q+n65glGDF9o25UgPK/46kf1oqtF4EeKXBnx
pEYJTAjp/+sAdFyul5QU8GpaEcWeEHR22+oUHxHU8K2psR94GhD5mirA7ci3hi93
PBttCMjWUjxlHL4xDXnaL6VIFPHgXqHDUl/CYH5beLn1oP5ScggXWgP50BzKrgmT
9TcxE1MZ7GrGwjGuBJX84c1t8GYunubw4jOauBWHT+Ul+ZQekY1WacujJr0oeHNL
v7/Sdw5SVSmZ/Tp1kW9ZnVuZp3vB/8oRmBT4HG330AcaBmWB/8HqkhoRLqwkptB6
VTcPKyNzc4tfIOXNALsB3Sd7HIpP2aqMnc9KTONyl32ItLaSB6YVbTF32p7zjd+2
KxLXSkbQNUzyuIbeM07Lguu2Z37RTYVPIKfRHKKUQkxbnxbC+ynzfoWgnVevMZdc
k4oIz46i9yV/v7X+pUz/qko/oZeMBx9+bnlP1h3Atq0/YnYUObcpjUsgakfVsRZh
d/Np422La7TlNQ6NeRWe1H1nH1t3TPpz9JC+1a10y1zGxvQuEcCKkq8Zw7n5nfTv
y4NcQu+VftQzViKazjMcerKsgvzyQ3oUE2y0C8Y0pQSCJgJrrknzThsZG6Fhvgl3
H1x/UIcWwKSp9RjtKgbosxcbNDo2Jm3Hyl99bwAI1yFVZlbMKk5wZbWAB3iA2db6
C06tGxQ2mMmvMB7MuK8jTFTo+a+I3GMHmxqUEO4ZPQmpovEGqv/WTB1s/gIUb36f
a97+42PHuliP9G031UhBbN0hYtDlSnb5kSYTgnvuNojzswnJRYo1K3HZO6bEEVDR
2PZJUWYGR2qJ404X0QVZQ5dtctXieq41AmIpB03bHNrPprkkulsHb6ybIF1hcZ4T
TuXp+YD8blAN84kjGrYY5xjmg+BXOiPLi/IjVbaerNnoc6jbQf+JHRR0BjSbtiD0
Ft+fGuef/3zHXUALNRJSS6enuYEgz8HnjHvUBLRRymks68V7+H6vanyirwC0oJoQ
9PNuDo4EWKjF4x1O7mz9UEKw9oVlBJKNRAUHi/BMx/cifR6ogl1dyrw1fldswz+9
NZBVrJx7+RY5UIkxvslJ3VSYLLZm1/hRgIGEw/5GJeTd1tUrrWNwSgFQFAoPKsXv
8E67GMa7qh6Ty27I0tV8sAfeT9MiO3EE26qoN2xIwIkcY9IVpNV0i+V+j2k6Nutk
0XwjpWCPDGPljQhtZKTLS35+LBDMG0ny5buAzFJ+ZLpphALz2JPutVdPYfwlxGOg
ppU0FfSP82ncddSr00kbbtfm/nqsThFgsz3iVOQtnVHMBvQ0TLA8nUHAmfglicxT
Py1kDE9Fp0oaLW0+8gMblG2Bz3lTZVeljzNkK5lWtIlEE+IZRFWdi3j56Y2XVX8K
qzXZ5jZax8KSNPfIQ8tIC2tCDGUp/f2KPWNMxccCKm7O3KGEJdW/Xd2DQ7ec02TW
97UUh5I64uO9GwjQIr970Re/Jzyd3Le5cf5hNDmk9DUQA0GyX9D35PTGzq11VnO7
bScVu/tS7UM4czSmwPpuaqbJWGmxh+AFffSZd/GRIeRBykVusrPH1caEZx/mEH0w
xYlLyMm3Q0Bh1JzPjRZHmMYhiiB4CcX1eDtn40/PTJhGRnjStyMh9f0bdkcILBP6
T4icWNZmsspzQUNO7y4QGYHon+oQiE0hFnSNAsn3KiYwk6El5rgUk5+JRff4wuj4
g2HmgvjpWhy/Abel0PPMUkzBX7YOGPeZGHLYd29cwYONAil7V/MfnWPvBxpoWsMr
jwjHzMR3/rxkMHbVaXpl9z7VOOBAnsI4+CFvz6WbUAiTtjSESi4W0WwrJyFOj0gx
GGUexgFWfYRCvH0xbfFnpdxykzB4Dk8u2ViD0jDsoJtMgmEbxNmbFNgxgPX3jcfO
bzpWdhBDXJm30cbovzVzGvRVxsPagbfPfvD6yFO6vtMdW7P+06wM/8OgcWD7+j4N
81WBSOa7CmwVnKbjtYMjV2seuGiD+QxRp9XoH/WK97w+fWpsKa/G62maTTHn1do8
ZdA6Qecn7nBYxHUMv3NZPmL1ZIqumfTRbzzaDdRG1+hlFLMU+sfpGoTF2wa9g+JR
u2OVSuTYhjqOYi0J+04rLPoMrtYRX4oZE6kdzc8CHyR6vI62WoZo22KjC/A1Vi33
fbMyhVoA6OAVLsiXdz8VfDr13OfpLh9wgbL9ChZiXJuHuARsHditsqhNjK/XYUen
03LrnhNq8hNA+kxn1xu11q2YAwnPZdOR2OKG5vWcNtEbwvIcu92wtf4cDIRMHIRG
+hYJirVVxKeCiKdX1FnrR/0nmBvGxsJgfPPlcwSi3myQaiBjmidNQHZHBYgpEPYg
u8e0WNFlBeEkDq17NdafBYqe9TYIJoXmau9+hCr1mztSwyp+PS7plGj2CruI8DRS
VpVp4RFJQ0ycGcp8e3qYWdFmFgIrDsU9QFKG+bpPkfRqSzjY5l04SkPd9NhQsZav
daanmoYVdPi33knZsHHKOeIbinQ13NK7k8Ph9xM8Zfd5E1HMGBvnNoXPDOU/j3yl
GMPX2ctB/W+XztAY79i2FlvWSsDRlkjjUsiFdyoSq9FlKUSBWQA741s/v5MIPg07
wmo0VsGQ2ujUlqQYZ87SywrSnVxg4YGAuUrtQCWOIQV/tN5fQWPTVb706Fh1twTe
qkOEwsQ76LpfcouvDTqltRBzAPtyDFoyc7dPfU8nkiSV4GHFUeWOXwWro8tYvS6v
2Kb2xtsXhIXiPI3SEhjMzxHirfX6sUpWhg7K4ll9mUEjM5Mt3GYZAcF74yqqJ98A
npT17Pfa1r9MMLEhv7WwnkWIRrLknsdrM1LD4tLYAXrUJs+XEAlwAFqHlBDEkVp8
Fknq3lDf8D53gmY7buJN3dZ0n8IVMxdBPPsLOSzXwlGl0/VrJhIxO59aSue2EJ8u
aTr5MnULNnTshyKTq37Jz3ZCxZ4o6Z+V9w3w3rDnHKMMFORHpo+d0V1DLZzFpjFq
ZSO4UXdSWZIH1l4xyTxq4QrZDki791MugkvQU0OV9kqAKY07tEZDg1l9d153+xZY
FCGKyx2/e2oQiHBNjG7mkhBHDf4JrVMPXnuVSiF2DhtMsZkAbY2nddeXjFnsfSQ5
cgE/3X+VotS90n2QC1TVeQbKJEn5ylFAwm8/dpyeUGr0fnAnjhjL/ThSh3+gFc1E
N4yfDwHTWOVZG1hvBrokEG9T4Z/+po+gYp8pJZ4DEuGdsASScO5FikuD4Y3ktaPY
ucQysLVdbSXaJtt2TgBDXtNF6SdIrkALIYVaHFS71quBWkxU43lkKAhuXlBSD/wm
/Y5GHIeZU3HQOLOMUK/bKi1a/G3Eb3dWp56pIzJspvq7TjwckZdqlAytJ6SgmQ88
5wJryH0to/Bkn1CBDQx5d1uq5AtNkB7H66k9YvqX0TuaEyQpPMocy9jNiuK58rR7
A1m9M4PHg3wFWyM/WM2kYiHD+JyMXdS6nxJ794NHwv1k0xFceCK2v1UJXbETZmmj
99GPiW9Ylu9LC/GzaYL1OpkzQWN6KVIlfI54gCgfVL76WwE9wnljWOGuzl7qxDlg
f5igg0MrzclNFlvGXBrW4FiSxeRjdgCLYrUMEG2q0zsWbaaM1FzuVBVdVjIPc3FE
h/AyZq7hsU/KHaZDv0USV37x68cxBRdzryRCUk6gNpFKvc3BHl5xpo7k9hwYQGBc
eEq8uVpVSqPyloQlZ/zzo/u4bc6q8Z8WGeTLuGwYBfWNXIFKu1H9HycklLzIBsV5
Zn/keYDN9Kwqxm9oVEiDF1GLBKWtgo0F2P9Iss4XPc34U1eE3TO7R8bS9az+hJfs
5ddff/dRcu1T4VkRy3Anb86/vUL2DHqrama3YexUSp2wsy6LB37mm4QPxXm23ixa
nkIvohm9dTq1h5RVxioO1JTeVXx5izmxZ7YF2yFH4dxKUyaSwJRdAPQGWsHKiyQO
4QFjI97Btpcqxt3EG206vcxMi0gshhCsDh6mTtTG12TXqBczLrE0byGzEf9p6/1U
Oh2zvBvIW5nCZhw3k/5mOIM4aIibzVUehWApL+iLvs4BqkHaiA1FnOb1astsbqSi
EDPAYeLJrPauuQc38p9+6akkHZtCwLIJD12Z+tvgSgKsbya2CWpoD7WqNkj6KMVM
7zkeNcUQGYQfot39/HOMIk7x7MbPiMI3TuD7hhlkijkVb3TPo3nU6vV3v3TFneD8
t/CbEDkqslCJp0OYjAhDkkIMCSWKSn0Ki+MJiL2qLrJqiFhKLbwwKd0rYEj8DWOb
yKfNNTdZIbO6F5tlC6qwz1bJm/VE7+lKTKDB5683mPkDq2PVB+ulpwLBVRY1fATC
/Hs9NXmq4pIgqD6CqIIVOd4nJPkgh6pw+waOXulJF49RsMEdJuFoaIhlQWMwhzAm
oga/VpmFTt0Pti7Ls5UoeLD/yrFFUqagaVzPhLKcaeK0UVzMSCt+iGmCNL9RPsL2
lwuazmQ1BfRIh03XRqUboVwSXSb9zkN8T3m0TAkGdYOddYQeaBonqD+O+CSqY6VF
lBQO7wx3Bbokdmx1zGX3eXn42nuFAjUeLIBazgV6iD5lpov4KaBi6pZWRqXBFlzR
gcatLiSSQHzbNPuGTWD424/+QaVqwapKVRO5cduT2coqX5iZOj9d806XZg67SUJV
VWGawKdfRutVpP8NwDJDxA+ysgIOdBkqd/0lkGGu0zt7GSv2JIYrOcGMXXGpa2Mv
Mu2z9jOCpkjzUe9zaAK7IZoovvBtj6PbIUo6e8jigJb5UDwogH/Y2R+IqjFgl67j
+CxpMeKZXEPHUgx5I7eID6Ov9QD8aAHHsVe1NBUZ1dLpV+pMcp0qECh1uZB4ddYK
NBWbrmG1/FQhSlyN/whtwi/cXCq6m6qiSf7bRBM/88TF5KYtXM3Y/NqQA3wSvVq5
e6EcCAHH6H+EJxvqlei7jcMMfbPT2ayDGSgwNaY1B+DM8IoR+rjP+kkdjOxW6zbc
I336yDyOeNcAan3AUChtd3iQyyClqCfAvDWQcvFLOEFRDk9YXMa+B7TWGQCDE+2B
EWUT3Wfn5W3VqzGHzuWrRbuLq38c/+cHZwsOYAyzv0Nlo0Iifilw+VgIi1iImxPB
keg3UiTUUE6fRnQyIfT1bH6FbzqhoecDeEiuFc68UsTl9bK1MCisdAoNN+tWLsXr
xujapGc3C7CBc19L5L/VAPeXQUeS8Dky9h2z64Tuj17uRRAeY0ZlEKaxIdo6y1r2
13/ehAjRaZ/JgBy4swmGWOaOHSGk9F0AdEo1y2ZyntpndlO0tl/3BoRgg2OTC36w
4tGmjdP8mU4Zmobx3Y8k6poNsJW0F2Z5UF8TrmrdiHMBqpOeRA08VbMLMW2EidB7
3bibbZS4UmLChFaS8yeJjOyQ3VyrD6Ts+xoXd0Y02/jJSCg95Mi+tP3VKI0uKzJw
91+TQWYnP1XQhhUVIW5y9tPPQrqMFp36O8/UGUkpq0BfyJrsCXVTt8nB+L8WOVw6
YzI6cRScRF+ThVHV2IAj0v/bE/XHAmEi7UWB2QxMnDhOm+ppsMYEyCQyTgd9umJI
5U7duVo9hyr7siew5J9dzAEXhFIuzrgHdN50zbeJdwEODw6ZKiIJQcRiR6kZoxte
y3Th7s7TdTvZCBdAIpwTNeT1x2m5VGR7bqxA/q05oxf30rgYr9SSx0eSIntFZliA
e6BpdT0bvkn2REif2b63j6z8GXA8h9/8MJ55KynJHnk5uYtlUtyN/64Ud3srgwPc
dLf00adsIiAReCwBtj4ea0FhtPaoshKUDDt6c8HfgjWVFBwYIRhYJmPDFyzS3tES
YXA2xxZu/oqioKfZGW0kFzoAjAk5UxcXBNja4VRkNikf3GCrf1vFdGEtiui7GwrW
6AmXNVyauJxf8SwBJFJkpTJjtk6jD3r1nG+9Esn8ZkM7s9ihh4BHjF4cb2t/zCGE
gX9HDv0AQzfJpVxEp/e14npd8r7WXsCifws9lCL8+EkM1ygRZCPjgD0JdLxUuS5A
LGFWSKPlmgNlN7/zAQQpEVGOh2KbRwtINgTj2+BlvMQDNoVVeZndAFz4H/r5jpRG
LhnT7dm7RBzhymR3Mb41bZJoWwhod8CJAWOHesHnvPyD4yTDdUTeEM3vQ4TAPxzW
YU+gDe1UJLidFVutZPTYVGkc+UZJviNYjv25AnqNSQpqYN+d1UcLUC3nG6WDUsq/
85FuBAJpZCWmrJz4bwL6tbQuL2y3MetteSMFUivjOZUCaOXPyTOdevHcxXaFGW2q
j2rRGqjNf8GRm0PUGNGFHC0gi7R2yfZKSC7YGjW4VKp3XDUxwaKTsXPRZFWPRso9
tm+WO+ah+mxQt/6uDrTPlML1lDE3SDLT4VIclVAJ523py2pLIs41PYsMh3cbTBKV
Q8k9CGr53FCHEMFlF7GK8Yj520Nbqa00DO6DbgJORH72aJQW0rfJ/Bewn3Fuwdvy
ATy+AL8lIVFMTt5MhqsNtRDzXkNuMG8GQoAUSXX7icLze2ccwSKy6+zr2fwHzfjH
bYlCXLTLnQ51sZYgwaAoSBHiF41jaPUjP6ZyIQT4xHPO0z2VpuybadFAcyg6kwNk
WdVR+k2gRnKn6n669TaJ9Fct/1r7TVojrcnLdjaZezBKfvQxWu3ZO4XCH1m3ev2R
sZAzcH4AEsEa/wU0ZnCZDH81Ot6+X/3j3iX0KGkM5+BsRle9IEG+U/DG8f0c9pF1
tf+WKCJakfwCDY3FRKCN8Oaqb7P8og6g/kFnZ4CStZPQRS8SrajqA1oW4PYBmTZ1
UDk/MCqZbmjo0rp/J/gNwxYy8dnPWg4UiQA7GCd6y6joFKSLj/oU7VrQFSoc7zba
BoHWio+MoE7beoTIpJit6xRTcwI4u2nK/wv0yHY+3ptoGbz62CXrKYpMu3XLs33v
U9vHMDc0aZduNahMItZiYEZUuauMOqKU2hUdqBfyG6tA8cQsNRWfCdhxBZurW6Rt
f1vNBKyeWpGrMEf2UjoLY5Io12fvyWDso0YyEGLSp9FCjKdSleW+ETfgXS2Cgpfr
I+JSGHasHctQV0dbXPSAhmNRP2BbqoFYMDQ4zMP8p4jkf08XOaYyHen5mWqc2SdT
FHGH9O4JC4AAdvWS2zBa/xr10MwDwAs357OLtiBQkXEZUeTWSoWEL2hB/grgqe+0
kUGcEAwZkWS6G6ZQL+h8Tgve9AZBFsiO2KH+eukS6sfWoBcDYHhdt2hdCStBCAC9
b4zHDbE/IzWnv2oRJJrHHxlISh94n/U4I1S+89k/8gURIa04Nk2S0W6y332gEV56
jFVc3Aq83i1iNSUkYrR9uBIgdK7YJLpMUiW77R6h328mJmGUZArmzmZAJvNwMGyM
w6b5VOxgJiqR8sZohV0IHmF/chvkmuybTPxXqa9AuZvqmL6ss/hQOy/ScbWqq1vw
sykFlvQbh/xyanY4KJcguidyxdqhFDfF9OTgHysncJG3mnycos5d1TRXUwbZ4lLE
it4cKk3d7boPKocUlODvJ9MrUWfbjg3Whf1SH4czQdtnmXhORWLP8CWsOn2y72O4
PCsh7KVKc+raB4prG1z49XuWkKgLkZi3R20KtUAOq/ZOq9FCcjS8KuHXgAIvqSC5
00pX0z3FZ7AggNkWGzyZQAWqRihVQzZhpSFnG2e6+BQh6FEmbyhZdfWjwNCgAQhj
xKHEnwa150ljjIr1iHxb54q3N8cwCsjhWghLwvNcC1WQ06ZWFBSwshaIZdCL8CYB
SXSgIe4j5gfP87N3vczIvsWiXViMQsbWZ6a6pzYsockbP58FtRMWZ7mTTZsPWGid
4pZMWagmJ0OctgPE8wPlYesd8SJLuhsQ/28a89RNzUBkF8Z7SY10Jpvxtbj8cWqQ
gEZUqkJr8mOE9O+JVtPBBSiJAAUQk7Qht5wvRLrDT3Prt6cqY+pj61ub6zm5f96S
bSlKb/xyMZeC6g78ZxiqQngzcEZDPgEwHfsaQx25mepGazT6ddAxlWKZQRfLwbYE
LCbVn0EF+QGSm9/8qNp0clfrgBJKWWPTbx8p0EqHNcHeO+UNTKPJkMdQMg0A2HR9
j5rl2a6nQxtLGU/Yc9Z1Z6nuCs9viiCYLkhq8KqnvRt5TvmI0Vhqx2JjIE8kN/Q1
VHhRDTCnCPE8+/djv5bc+qRMzkAPPGU17GQX/gRCdP2DKk9/YC32PhvKrqU4SOwX
Ltg4CpzTHb/xk75aOw5JXKp1woNcHaXBRlw+z253RYS+yKiRDWBE04KHhIsMniQQ
Kqx2eT4yUeoeStRPvPCnMb4gR83GB7SWAjVPVvJfJeACS6ga7sU5bCEOd9FoOhRZ
z+WkCydr9ZHlC1KjAup3i3ss3fU1HC7pkiMOB7nizS0u3gjH0B6oqmwDBT0QpZHD
STlby8gXQIWSnF78DY+U1BqVE+ty6UNDuRB9vgqCDyrtvO47G/aQZybNivJtPX3M
fbSQSTr3S1LlQH1bme3JgVqUdMiPA3xv0QGQLc+nDLVFrkwbxfZyURDH+CNn79IM
g+lpfx59VplmkOjnvAcBHDbw7af7QjxtnOFgba0Z9GJ91WSMfX7M7C4t7/aFOY+k
FCnXkHaOywMusUPHlNXPJblyXznsFbSH6/vp0KqWlAWtFnZyku3TZcrmssgk6WfX
UiAfRfx6YVhHTZFoH/DrGdP80ZKlgdgSg7ch443jDHqF+keF6TOWcPlhUvxmvv/j
iM6ABFTFFeTB/1BKW+THVGPTIvmrJFG8fdNQ8Dg5/+CydAaG9A59fGBWBmNhpMAc
nmYFiMivLtr0eall/2jvHCJFKh2+tnLmNdI1tz3h3/BBdTZ+5dHe78yNuXvTcIEH
KAt9WASHKvPwGA3wDXHShvsTkd8zH3mxK0GoWUzuGl4BPi7F9YcYVp86ydxZMy8M
Lg56w7wJlbqQbEUDw8fDQY4Kn45b1K5Oh1ZmhnhlRCTQRaR1XTb6EWc2lcSESV8+
MjDSG4n3UChoYcqAVnIDQ80E8EyR92NfVmuehEtsTn3NKji1o/PBAMPiq2hd6FH/
H82jELWTqFer2MOnjB9Y93SjWZfCbtqbyU0ikwTpI71jjs486isRf6vScIIVMcrg
VY/fVs2KDFnmubjJ8+RUfXVZviR5Mlo94LX/Vy+NZrsDkrb48FRwsP2VmvQx2K/G
OO2wgLtSODQbBNJXy/2YJBRIczR4x7030erimAFT34W9Wuhh3oOL1BcBTPnZAPW1
v6SRVjNjcQsKbB9/3T4WR1VcEl2W4Vm33fNDGqJjlpntPtE+IxeUmvrYqeKSg6Gv
yw7VHqfzmk40UobMBvLOe4StSUdCzS/0Qb/ys/SO836nepLPGDyDd0nvCJiGW8fS
B0Szu7rd/DVaukUVqa3ELpp6+RgSELfnxjgyoGfyU6D26vb4eAPl0PX1C61Jeoyy
xG3qiToE1zuTon7mDSW+OYs5RY+dEugoXABit2Y+S5bmwXNA/mluKsuCLy5vWI8b
DUKGYYIbj+P95BiiamM8cSaMZzCgzbSZRUKg8JFpWEnuZR+SGD7kh52COI2QtHya
xvuW7LwJ9A6BzJHiXUz8b5HZOhLMt5CHknz+kq2P1EfJ7j5PFNYZrK/H7H/DS3wY
v7iHYeb7XJPwNdhMMnBi2gssY1NLKtCB4KSNeihR2lkJz2+S8bKZUwZ4yOkX+5IE
QAflyQzuhCsaT6Fa28R1rDzJLyZdSnVOUgwNp2btbgKkCC6avLYtWNWCwyH1yEUR
2TgraBK2UhXn5DFFXo8S8bmKyJY5a5dq5CZ/JDvbqoAGhfr10GXK0UiuNsaCHD9c
+xFFOvCSYtY/3Q6WMxkvM3g4ibWOgy5o4r55ASLGMzaANnAn8u6WvbzFOcXAcLi9
d2pPRGYhNicDR7fvUoiBo51nuj2lasQMKlS/QtocGiAXbMRArcQLKpClFukLSEiy
8kqJxjR9Bk1LmW2461AK2MKhpimkaZfoz7IelDNcJhEpDFmPmq0k0/2kef2dMj9E
EO7Wr9ZxkTKgmqJORYNRV1X5K7QCMNDg4sFBgSTap92EWXIdoFx4oovEp+9Dg9sq
OxZM1CYMkkhwLiOK+mn3BZLHcr+VsqiBVAb897M+REglNqqa9dBgq8EInEJdzJ4u
TJAs1iTqQjQOU0+GPy+ixCVlyXt4AYMICQbf4zBgQTt1txAvOG2ulOrcwrrHNrXB
JktEYSn3BuUc7OZKSQO8YYvT5jLVnk39mtGRMZ6M2Piq/RkjO/p4hY+4wRUwo1oH
OoneC6UDd8of/qxz+wuV+JeMkreMN8Nh1KWgKB/o0Z0EbxRsHECZhtTyRj5igcZq
rCsjyP7bNrRhuZfhisIQyn7CBnHWJ1mGKOBjLaYYDoAYkz6YK+00LUFIxg+PoFZf
OFzXzjoVk5CgynQD67K4Fi3yplozve4lrOlQNXLhBmDS3PPswx0Z5kJcYkXXrzUo
1vWG0Kt9xz4x+k0/bAF0rtY8Pe0GGe8bOk1xsYY99EAu5Fmf+b64LanOf6PKZ8ur
z8a3SXCPLZnRUF9M3NZ88IdArOBy6wkRjociNmrxoudB0lRJ8kFP5tLRchWsYDpp
HjGIVT88Ftfu3WoFjRbx8sgeaYH/yMqjBeRm9QQIyOZLBLPsOVhKiqtCwAPw4bnS
yJaDxF5QrlOYSQ4XAk9OMyswESYPDfWt9bZp/nSzGWSYmjUOxMewBGJCYuP8datI
cSpMDAkcQEedxJAJHah2OMXXGDuHF1hdNAK2maMZ6q/GG3yDT1Bq/kLZ8AYjoXcA
xXfs8W61BUz5EoltaZpqoohEYNcMKJW1P7jfuaejNO3lyBdpeXnU+TL1cEs1tnCR
FkJScQUtioKGZ4nVTSPlOFxJIqjr3qC1GRyNfggcZoArwUOYG0a+bQnUGfBS2kY+
mK0XSqgqkkeeQiXSOcIEDOzh4E0W9KWmJ+y7sVJwaj0mMCc0R8APLhjBxe3/TKZk
gt3YoMmNDgA8zA/pVA/PzsnVGenwUiU9r8TqMZxHn9pzU1AeULTn6JHIvUF+iFqL
TXWUJN36ZRfjtaFQGMgMLwJLE6twLyChUwAcA4bVZcfu9VKbLVgbbHyyQP99YRHx
xwCDCjwsV3Da0iBxp/QmbtvcOwb1T6tODDfViV70eOpa8HteiSuaLRy83HxC+ma1
E+amkxcdLHPiUY+WNv5YhW+E9zct/3FRrGGptHNRZ78ijYY/h+9U6efWxxQJ1O5a
O7FBbwuDboPSSGhjwsUwRLZn6n+tUd9TnQ8fRvGLg9rG0s3hu6BSv/zIoD7sY7TT
Muaw3/QAUUICOfTxAF4rn6khCBYBTWkqaOm744x0XlvktiI45i6m7pfb8vWbdrYK
N6CGxw/PNUMb4cm6W4+IOlES2IKmgQ24i6XfV5eXOk8kxY+sPrjTIMe+O70zjTGa
5oV0jAyguMk6xQwbFOIMHiOacjeaFYL2FYeuk6HJFkHQfjahqGdFhkOQqiaBNdbM
3XdyHF9ow5XYDka2tiyFPGIflZfRmX7UPeDiHNHXWXomPNs7RyK1yjT4YayCDboe
sHyk07GZmZShEgxz/u9JbfJaVUN50wE8LRgUiE8zeKRthD7ws/GZ8+5cziyPmclN
43udVkPBQ0EGCjOsTNaR+yrXCd+PZGIr4nfUGwT1Oq06M3kt3QrU/h0a9lENP2ia
wSVUNbHIM4at2Clz5i0dU37z8i6ZX0x/UMrkOcCDY40XfjmctPD/1czYCzm32qMZ
zbU6QzNcJ/CEKZTaksrVZnqWtxSf8EVtnXsS9coGrUdGHKo4m0a6sve7OxFFLKRI
KV38cTPSOjoChrtZUEgONZUEvicPIVevTfaybQ82o2i75eLfWPy5yFUyfDUI8GT1
JLCiI/AHezdeKDg+sVQL8aWJI6SLj0j2trDf39s21Jl0jrXxoyfmQhLKih9SELV8
BF7/nXHvP0R/7+oOORpgZCva5CFE2Qli8sY1ssrFbsyts+4Q2xqeDSsLsLjSGk4S
nPE44AyezfCPKOgpAY80kz7If4YcAlFUeB9k2FJXvM5wCixdVzPuftQcIj5ZRgnt
7FIyem2Bo9iJge3vkSFaysOjZgBxWavLJUCF+V9bZztqnmuTK5qXyZCCfmBNWXjs
SnY3bhScO3o587fRhSkwF7quE5bsyBGySkedegalPVG6r/G/i27rnnysdevnD8TZ
TltHV127ALXvWEOiYGlZNUbQeInpgUX4xhwsR31WNUKaSecON5F8rYzX3UzZIwle
q7ZiEgC6rJ+yjcZEkSMr5LGdrPy39JqvbM6qjHDE2+iVyFSazcF/pX2QdMyStMHx
ZLXCittSzkke4rYkQPyrSUylNsRa7DtL4GxTlz7cWUpIB/dAD1EfiJ2I1JQ06sqK
2ymzFDjsC/EMuLANmyQJU6Uh7LtPQlJp6Z2LLV/acDG+QlX+m0ZTOOwV7RXuaToK
01lH1KBinRZHeFacsG4c2RHblv2R6A78GzOgUDckne4VZFFuBGgDij3oZA0/2AYe
LjWCc5RfGCj3Q4NbvrJNuTsKbRUxt/RqZC/Eh+YDFlBmLHfIBQB1LEaogT4E/c58
StGFisIz/y+W5P6/A1WL1ag2xK9kFpUWU+D0brlyhWtWUSymsvD92NHZrVWOIWTl
5LKmIbSRyl3Ew72gf+LPSEo7nWboIzD0NFw/wIanVzVO7dk8bMI8oRMj4h7nCsND
AZbUi3KD9B/UW7FUQxHQE6x6rFZnUrnyu6Iqggpz5XQx559eEbJqmJKAjUlx3qJF
tdbEKngvZv8M9kriWsYRgyb/LCbT9n2D5wZJXkiRP7qAEf4hJhP//8ZbWthQNWgo
FWhuha3Id+OH31cPRs5ASqDwP684H/xm7XaN73VL6T88Vy8lreYNRzqhfBP6pYOv
6tmcym6v2Txa8w4nYnJ5hJioyYjiNHsztgQf70YKGGfDPozLGJ/ETn73vwMcLNGj
iuZt9IULOCWGUEoqeHMv83HSH/AJGSRLEtvi8850xT9jIEpf3iuYbY17mDIFecxr
IPgXGMw9n6o9ByWltj+7w+05Z5Up347RiWe7N8VIDqX47C6YKNMmK943XNflWIGE
pU++uVpwrqbSkxiX4cpxLVijoS+A/st7uD3uXs8vxPkp9oASsknf6I00J901k85s
fLJvAZnXXR2YOOW49riPUFsVIPWUoVr1aL2eqla/mzXKH7cNY+vh8/b3A+JrcDB7
rmrxDDsaxqHdtQG6acDx38oMZ91y29yRgi9YRBxEVooDXDkvMManqHoSrT45YP/l
/cA9nUTddfoKZguTJI/Kfn2Vu5W2HcT+bT/qklrykEWNuX3Zi66C7KJzqNsX1nEe
zyuaDtRpHOWyG3BgSt9B40E8PTHN6bkRjxbzFcXatyZK3SVCSY4PBX8gWOWzJnLn
wXxb1Xx5I9dA9m14oVeZPy2HzaeeZq2S0XKJN6B5eA+iMEWdks3M3KvDmrE5MI2i
ZF5tApE8SeUEN9ICwaSHZCT3XHGqmnlXtpdUmxfXni7/74n3fU5LjOwhUpmR2Ess
WWMqYSPqkKljc+aL48DmFflid9Ilgj2QmC/nliVTKbCJc4wFLA1yfX7zBHJdgPzv
unzNGwaS2Ck7XDjqqz27OASFuDGQJ4/WHNj6yW+rgvbrerv2EFQj7j1Q7fo7Amky
58AdyqnBA/yPl3miKCp/8HcXz6C51oqML5qlUXARHDjwwQM8tNquP+G3uVUlXl0W
CEU9xbdEhr0aO1v0byEcIfhAhyQWHjHEFJoJJitEFZEkDY6A3naw6eAi6C9VEEz4
hitJNYjT2Q8HtB+9qpdmZW6HMqpA73NTYwtsERC5yw7hILNY3m5Z7top2uyJrxUt
tWTLcpDXatLK5/5o8vfIQhKXMm16Jp3D6hY8fIbJhq0wRygAB+9OAsD6wsYDCMhc
hMmQ3/f1jD9iJJwbLJirGlahtwck8MOpbv2xW35cOb8Xi22vUHmt4z5j4Jk5J8as
pa0EThXPBuORWhw03hX40Olq/LCYBaStn/IFMMXhFRcFPagFAsyibaqlJrU2Po5N
HW1j0ouv9oe0xX4qECgtUjnUYa0tkwktbBjLdvBwckgqqZbY8SDpEZtsTr9UJeEL
H+YHkqN/kVrD5pZsgZ3tuXc+OpRSkVvti+u/pvz4bC79zjoHk+NEHK+tVCoYgDuz
V2WHJwn0El7PBecWM0UYjfcPpXFh2oV2ytN/ae5QqZ7W+z7e56N6Ho/h7/S282/i
kO0cPLrIMmlJ5dnvPEn//Khlop8tkW7Cy8VhzOotaLAX0hY+Ani+Rfg4euernrpR
Ic3hzrVvVIi21+/o54GVqITEn4XJH105Q6WJHtOJ+QpHe+18TwU0jNinpaw/OLJJ
+BodUPxfe2DXQiJ7J0aKDib7E1NnsOa9ABZml+05Orl4DdZYqu+CfX/8mHZDY4BX
T+DIvCq86ihLpcvx08SLdgNs7s81wMIPB5fPiYU/yU4h/m0jHcFgU/d6sZLTRxoo
DvTJPgGYj9y+7+4Y3vP7v6FgRWW+FNb7AqITxTn5iLd9rbQ7wEaenLaOKLxcYGSF
U9Xbttq5GKcpcWfUKHPtsG8duczj7sV/xuuu/Dc+CBnsMbUZoorVc4ilccufU8d8
wySgpfus7aZuPAi9hs2ZJ/5pVOFh2NAcbODL8HOaXP6JmuqGtj6WrCEugee8N+1a
F8aThEwPzw9Z65z51fOWUgSNm+IbB5fTxIgUcRT7Q82qA6N3MZX8mKzD8uTG3Yd2
GQJ9MPrmhmJl6lzuo18svFJE8JFIeoFH5heVVkQRXTk/U0clf7Ex9ATYAS52uDr2
TItJUBN49hw1+hrSVAdQdqgIHCYrFxlksDUgCeexnOvsyH9DAQFSTep5n+iV3Z0a
deDdtsqlpgtX/8i9i/uTfQ9txWY5h3qRxPNK0gA78w/J3lUW2d3+MLdBjeyT7aKS
6XSJJL64AAU4ds2hvYJ23MAxeO9eAUMasD1VJk+Jrrf32u+cvm3TjMw1y6jIscUg
PJb1KYKBmHGkaimu10uqplA4nvjlEa+Uneh4ecMh7mpWTJH/QNg2YUjfYq2JQOCq
fVXDxx1QSuFzlhOGxWP8uA4mYNzvB11cksH1C2SE2zsc/fLHrCTANiII0GMYnUFc
D5BzoEKagcjnQkl5V9RwKO8845b1lHb3Lx/tiqRiBFCdZi1nbEQFXgRZb6+GQRmp
DOVNdRXSk4jtBt0mUy1lbd1FUq6g+Q/AyhQZxei07dXHs5zp+xPFtKWUlaOPYIe5
DUh4D0uYz3q0ZMqS4fAImR/Izu4sZErN8ZX4cPnXNPiswHSxWoV9z1y3H/8bZ4T0
aZdGeQXrVy1CPnuXmLpETUL3sxcy2pkk8qlzy5yLvyindhg8cJt8EerOM6djc7Gf
GVxges/q118akDwB7rky6utEjCBWjAIpOTWl3ReDkvMeYGiktaV4SXuzHlXHNvKX
kvIQyWn5MgoHJJ2smbremGSI24HzCzqqZr7V1s9g1hn6xUGmvV8GdDNyDEmcAMWD
A+nCT1jCEcgpmtagkeNyUSxupNc5MQwh60V5L6k0ezz821hf3t2ouMHGAB8pMUiB
VwM1JRcN7H3APRFaUVqRcLyb9Btrlnaufayh1cXNuQkjLHFtFfAqJ6ZjNC4UqueM
L43TrGg0qaM/2qZYrjtkpu6ZNlVlAlHpszj8RnOM3PUsQIxzPd/+rZe7C0mYLMh4
lM0+F9wIuH9aAxb6+y1fQ2uZ/h0JgXerqEdtrS/roAaMVl4orBKDO3twXti3Re+z
RT5hQTPZMXu7WAjXW5Q4Wk+MR0nz7SPR2QR1TUJU1y4G9XfEmgY+MuucrCgcrb4C
wgy0IBw+k9WldA10BgInL38IVf/1YP78ZKf9IkX7FMlH+yzAbx07gsi7Z6x3M7pP
7q9MVDZaYHpx0a8API7XVKuwaqkPfqeFvpp0/6qj5FW765FMy4k34dxv0W7GmlDe
xLkE+K2xOI7GDwex5iHXFc4fycXZUPCmhP0y8H5GVv8Y/rorpsLxqZkc3L2adOMN
9kU63L+5FPX82nu4MziB3tcf7cfgyI/rPmSeIhcVc6ltZmzUksJB7ejgAFkIYbLP
WGjAcG7LX3IGO90AndJ2Yn2isW7B7nqHMKoqN+00BRUD6dJxtI4Qv+DekKwNr0dk
GEcgB4yCbkZqlkB8Eoph2kvuJHJ+ybVW/+TCh4TYQnHODhq6nEyRFx6j2m4oyHPh
nYuvqYre6bNwKFPuwRSanc1gkIqO3P3g0dNX5Mac6RZ/c/xdGpDc0t7bCG/8boAF
VYqdGPQVR3VvzPBZuwjW5LCyGa62ZYyc3ObLUie0/ZSqK3PVty9H8oMqJK+GLBoX
MfT8kZwiEjnsFDKyVrY9AJD5m2mwZxUVu6dMdiShss7X3thkdRCoHgQ0KcbNaxXs
Lfl7/DXhtBGyUQ49rK4QjSNnIKs2gHzkOvhiKGpCq45Jo3aAE9trvp3aLTS6BovW
t2zR1YU9py/ZMbVJbRT7SMfiAYM5h+RSWHgbXxlLMwPytAhnKQcizDruB4lke53L
WIiMODPTFtYpOcSJmr2U8t+4gu/Z29tjMb4NgUpJS/cv2Wx9RnvFQ+jzP4Yq7GAJ
yXB2sBWKMczPOxqznt8fltBahrNC+SaOstJfnUd5AbkxpoyxmKI2LCGJ4dSJ4DMd
aoD3vK4knJ49vvHCq7Bvl+MDw1Um1KdTFz1lyv+aqDGMRm7APNAF96z9adfi5646
F7tjgwsfYceTgJX+qkZ3StKZ8ZU/ZBCIHmIfDBlfZTGdpbaLJPyCf3g4RZeSM8DS
ZxYwTNmZNbEbSe/hhYu6RGuQXDLzdCIITmsATdD4d04OAWqZka7ngZUBfQjgOiBL
85NrHCk/bvc0UHZBQflMZRDS6IOhc+qX7xcBkPa7iIFaucewLix+1UqZgfA6U+Xw
nSoEp0xKYWHa/E15ezx/PuqYpKeJ3KrCeoOHAn6ZaJmPS5Z3077SZSKLJDx963Jl
gHUA1hr6BFUmsOtAIZLUS3V4loWw7ROtcQTgEylD+P0xhJsYXfw94PMo/Zv0sTUK
XJR9eHCSxtug96lh7mItrSWpN80pyrJyTp2uS2Qva5iKsCkKZRb9RXmUUKYtNqhE
VZ6aVmXQU0I3xEV4fJj6hqhK2YOjkt3tvrlR3zavH0Awu9fCacZSEEu0X/UxhUuG
PXWhhiqjwDhlExECnRMnxZ78uDaCSd3ATr55bpNmbSXUmIOJW4XDnFeMvRMA8uiS
gpNRAtQN1yHyGm/nr22PzWyZjjQ7sBKf/ACoOVq+ibvCbZyjVbWsdSn1+lZNjpO4
TQjdgE9tHHx9U+kqbQ83yWTVSje4IvPH1lKLU3jYbBV74rPXeIUowBKJB0/5GdHK
QCfYXaKPnTVJBvvZAvUAKkPl1+2en6il5hzeRnjTK41OdmEKbO6cwU5wDYakEh9p
Q7We2n5OFjoYi7GfueH0l+Iq1oy7n+hmIrECA7pUl0BwFrN9ToRqnGHfVTfcNnul
yKxwQMujZ0EXiKHTpSOsaOeJRVpECAZ9d4CiejCyWH63rL1w9C/XSfo+ESiGUiA7
fzs0biWiceFgKZvfeSyXRbHMHbGNGj7XuPjHLcHBKqEdml6TCrb3oxlk7dWXHHQ/
aF/20pU0MHiWrvXJ4y2xkVXmogusvCwoZwAgVL2X+VNVqcaR82ZPOs9UshCyhore
KyZkxdgqo3b72G9BbK0OICl3TWMZph+HwHadCqnXksx+3GrnVyOKzqqs0Eag9JyK
Q1n55UKsACEcRdQ0Ic7y55O3kzmD4OtOs5W5BggLAtbbSJicFNw1ZN3rdaISxe51
iF2HD+gnLEW6QC9Z3PJ8staga2JTVQoBZNbhRxL7uZiOt2Dl+V8biY0x2ieFFWOh
+XzhXiwj6W2yNNO/JvKkB0OmG5+mCKjrszZs+vGiLoWolzdjUM4zwdCZQxkR8pdx
/r7bJtMbUE2lMWmhGG9hnh5FKmZYKoVLwPQrmjl/9DkdgqDGoY2sEG593btjVRSB
qm63LWFZvzvVjeZ3X/F91NojjAss9UwJtF8PiJ+HTB7vnvAsMUo3ybR8EaPoM45N
16kg0LXW21zfiyoD0aMyqr/rly1Wm/8/kEHW/V8nd1/z4URA85uAtP0OvD20fXEs
RxTI8n8rMld4BUdpk3KQ+KqBUPgCmcNP75kmRC1Zh4SHFsdGz7xKl9d+V9Y9GMps
/DcqYsyCfwCK8ksmnb7Uz3eut0r3eOBXVdm0z0pH3k/Sh3iAvKpjDJrkiu9fTycp
ZEtprhRhfr+I/hmiyHj6e0L0DD6TcSSsUMf7xGSZdSs/zfz9/Dw+LKVAAOFs60bw
VfgOynhAKis741QEasAl7iTG2WpwoSGRpPtyepcAWhqm4yoOryoz6gPtLS4fvYmv
13OJLoiCFNkVmzwaXa94z2R6FRbvPebhqsTF0uoXrWFTzsyenkRuSpYye2N8R5S6
bCyORgpEqdsD7U8ptZZ+eqinQNeFIVtNt9AvcUnlb3JhdLiAoFz2Wv+FQUZQt+0R
lXNsClKxJq/I7QV8vN+FDOiY8iLuQElS244ROpgJabvqjI/NXl4fbw9upKCH21n4
91HYzZ1+14Iru2n9OfAJ9iDU8biMBmaI4Rdu68SdHwdyt2C/NmtS+eKFyB4q5aZ9
mXfCx8auD1vLdp54pqp+26CP3yKD/ylOJ5F5EOd2tMbRdo5D6AOPU5NqDr++dgE3
wiraxl4gAYcFAxgitgxP4y+SMgJuwQD0+Vbb8b1va3SOZpLFNZ4xyd62ytQdRo5y
DGQ9xMR31eGgaxk6EsdGm3vJFnt6+nwv34zposugHGBBLaO6jv6AJIUBVJltn7cW
cEGnrVHPapHkYG3CDaIs/OewJsMtIGyLkWdcIm8j44tvTd08dxnv7WtSwO1lanFs
VNmQwLrDT2G4sTARPdXWQwCmezsTxjjiHVftABJgJEFyQUnMjaKSsaoSTliQgnMU
GD5fXARTTxFlXdiH8GsLSGESzatiwYTn/KyDO0jenX+0G/5hgRPfEhD0EX/87g2L
OJyEZL766EmF9lYMSgRlOE5jSO9rS0wgvSgkthV8xrz3vogMQ1ZUlVLxlegPJEQh
7IqVDkmS8gWafPoAuhy3oXKrAaVm6bwCod+SMdF9PyDNU2tmnGQhMdXriSG8TrOm
n9B4DOHvHlOuz0bte14C5bbzQYvJp4hhtUBphrbvMVTE/qx5gWnre2BPnb0sPhbn
Fej5cs8uDD1IOsWCfjr60gC1bBjcyUA860gEJNzVYOaXdSU0gysAInGtpTkvq5Zd
XaZLfZ5ddIIhzRfzJhMeF+PqUMDHDtebGtWo7/PHUHkGH8z3KCm3/x9iA2n/I/WV
mpv39eIT73x+/Z8Mwo8Kt6agc5w4g8LHxn7rZq4c0WQpocVQCPw1eA2inmHs7PNI
QVSSFIta/x7CrKolTcPfsX7BkXuucnHGd+QwJ0p7L9wU6UnOprovelizVCqiGlPz
QmoinaqLtdjoQmDtghkZis5RDFtQRbiw7p/sMKVlT6UKNbTBODpuSpL2kPMC6Mhg
iVAELA2jYkGuEbNQsT23l2Ofy884i/3EmdWqzsr11abOwIRtPcr1MIiwAGVPUumb
yNcjeml8HGLL54cUtOJhEU/uX2BZJwvcMpD00OjjlcZUrtk+Xyfoy2fBh3Myb4W+
F0flR35h/Pe067m8vUehC+L+aVNYffPc+SkLXz5kIha46JZXnmcIMRuLr31boQKW
yD6yg5xwNDga05O11aHxQO2ng0JP9iexTo/+zwgx6YC6rJYavB1DIwAm2p7FAF8+
vAUfDx1jjpm8OkEYSsCbHg4MSE4/BNED+xGsCPRKev8dk4RM758aTQzdcq2gxli8
wQ/CRxr14bA0MeODD9U8lUYpMUlHpbKsoCVu0QKKU6YOXO+KfmXuV4sz6SmQWnC8
XYeuKTb1fFBOpGZDRWTG28aWQC1h+cnc3Bxr++clgf2swElbKoOIYCOTN1JKFdEJ
thYul9CvHXOgp5XAOWoB4dc6NO5UA0r1SVHa7L3hSlWxOV4DwkQyia14MA5bswKf
DAMZGwFJDVvgEJLTszWAbBapMT4whSihaRiptRY7n9R4oJNZRreyVpowLR7E6OMw
/LZyNLyLS846VMbBcT0xe4cLMFQZiH/5oBgyZis6kpfC9h1bTVQH6fFSh20LZYHg
ojMwJnhAC5hYzuH3egodBIhVVtIWs/Q6GKgW24akOPWgaQVXI8AtqY96PtV60XIQ
N1Dt3I/BqZp0ccvtokbzWbU9Xy/xtD6u4QiITzk8/0IIPxnN0AT/QiX/h/FhzvM0
MSyIPk9vd96dMkOhTS2HlkGao1nMCzsepecAl6tUagnpQ+SEffbzgvNxLxFyolAj
AYyBsXEFHEQSLpinifJptf5lzxMD8s7jbdNZHFvxjeoXC7bOow9OPI2AIjXmouIb
FIZHEqXeNhXET48bfF5XITlScF790S/973XP03bMAz2eLymNtZGiFxaLq7pFffAS
yozGy483m/0bWwNZzlNrmbzsg4u/2OPFyccKVQlTz8OwVLWjk9SKeM3Qr2H/nyhZ
Liyse5NjDJNtJm8g8R3yRQT9KGnMfH8I36zpt7nEDrx/DnNh7WnlbcxmfZUizLTF
abrlEwroxceh2M9frA0zOzEYRp/mzViEBwSEtg9FKEN7v8TImact2hDJtBhht1at
7nq8+geL0HM0jpCm1rVuDDuAw2V/smYK+VoZqwY5wjKLsu59zQhxi+yvjhRrIMDC
hv4dlbupiB6qAntkIYeyLKT3gC8d0CrJkA1UmZOSAcRGOUTfWYwlAkifgWwuf0Uu
yOt8H54/6qdaHiDkswQfnrUEWWGsHUjf9zbEaU7RVO8/SimxDSuwTfcGVowMLHbr
quqYAxcufYAQ1tWnsDnZZcFZETBZ3auc7XRuqkf0Nr984TBNFOn9qkkOiT1FxrV7
9GdN68qMoNCUfbDRD9EDZ/i1M0PZ5l8Cg+4gldkZR0K8UMQKJmp2EHUooQRXqxnj
6vWNyAOOsW1dFmqLgD+2gF9mO7ByvZLpeqlOA1zPTElOn3BcWrdRRBfgFLnfkpe/
X2A2LgmNkue0WcywDfpKN/ydJnxjhPhU9EzXBQYYzCWjysL9qg/i2yXXZHd/Bd7B
WAICj9DEnqdLluZrm9KPefHzjcDydoA+hn6RQSEysRJzZHKYXt7LjiDcrs96HNjs
7m7fu1jh6rOng1anPKZf+GM1985tYJDDVILgTDbtOxBp4/S0EXS3yQz9pK/4ZtX5
l1EnmnNo53VZERuJFaMVBRK2YT1VG5cpmMWu0fspjh4RWq07xyoYJb4sgLdTGrZV
5kekHnbui2EDKvttYriPgcDFxyUhwMHvfP6MeBisIu/DIeUBp0WGdoXlMug0Nubc
0fWeVueZ6IrPmtM1P7GKXTP82mlo7E9or/RGd4rGBNXLzPKdqD7M1t5A7jJSxipT
aKhD2/xGzoLfwfjhTUR0AwRb0ABDjC8+pf6PvgpNYi9yDdm3o6Kj1OXz9e/Yp8kv
qDv2v+iVbZ3gba6UX21PD4Rq9YpZfGZpaXm6LKam94kQv0bVMLrYwHxGY8Dx6tyv
KwJeFi2nICnNLrhQyTXW1DJyhuC+foUUx+3keKuj7UYWPMdk3zuBalupM2RGyKf4
kSydc5f4SEjojUIToSHQEl1i0uBiaJZkwdIPmwpRXy5HcRnL344nF0vcSscrT5IM
6bhI6mldQvPbNOzWAXLD7aucZW9P0qc6SeAvS8EQ0QNUViTggmeJneHiWrs4l8p8
8OJrzo7zcaAwcuRVHEzWqnvS7p9nyUUauubk6om7W1AIBr4RfuGPaa2e7/+L4O5C
6Y03I+CpkoKoHQW40unrZmW/TmAKPJUhJgV1SotMVKLFYQnmR6OpmC+2HZx77jCl
gnkRMhPOqzNHb7/b0Plo/OA6Xd52tIzQbv87mD6yz8FQXAsnrKyE8EoJT+VYxyxc
+8l/uvcLPr6JlfItIXRv7kCoQs9CNaa3bpC4YCX+Qzskk+E8clZ2UbZEeDJp0ibJ
xbgxshNPX8hr3gRmqW0FhRxAR28O7j9DvSWrSytR9azRpGhWdb41fyh3haZRK30Y
Ql20skp24rDmwtODjOSl1il3106u80yYntr2lA0DH7IJ1Nzbc8t8IAIcbEYbso5+
eJSGxKujIIYbwSvpyg90kgvVLtKhOR1vGzZl1jDdz4OZN6eJTqMPUfgV5DvCr7q4
7TtWAy7vxRWVSUkeaf4anKCKxrpnwON8Ho6qyaEpcIGoKNNqjBO1NrwJErmyk6By
eRc1wz+av1C3bIH0GP++m+3e9jVXjmYBzucj1L1jWNJ3l/BsBOvsxCmFf2pwFc1J
U0eXeF82pCirDb/BWUPLAjINQpRGKfzQTzSJjzHlARHd1Jr/KYaQiJG2CXZbDfQz
tRFy/3yEPlScEN7TjbJ2VbrD0UKZAPfbix/vqirdugtTqkru1wIke6pmzAhats69
OFaKf4iTAG8ATLyABaAqrlZlp+mpyT5GrFHhZUQ9CMMK6kz9YMtUcYG+rD9KiTHx
jC7AYwSnalmmjJn13rGAAazP2XfUb5/IwUv16GqeduGhsTYxHRPkxjbSrtM+b2Eg
ED0aBLJ4VT+QNfjVHIwnE5/8GBWnEU0T91I4vTrLVJSaV2V5QhCe0ZX8n+nRSsH2
qsqOkVqynMv64XMuLkAkfOkRtFtt+EHUWWDpcQLGOY99BAyKRfezrFQ0ZFmrwW7v
Q/SJCsdtrHPF6a4yDQbD0o1wRAJcCABJGDXjQ25WpvJI1PCltMa4ht8AGFPVBXSI
9OR/UGaXWUFCl7EWXC7fyT7CiCZSpe9l808kgNkM955wWdTxQHDq9y/pWOM6q1e/
avNI3+RGojTEYoIzGGtCIuTqPxtfYGm/GLWkjODtrrNhkSyYdSyoZnsKnRa6j/E8
6FznAbCPX82sMt02wF+i8nVaVipH+HA5MMMHd5DUzpq1fg33a7tTnUjiDBWolxpd
xmVwqVxpDZmxZEypUA6C4LKJfWKpNqP8rTMTmKPP4VQVBNpMlRPSv6Fv78waCK4u
9wqesuPtKUZZvlnZ2K1336vyQxjqYTU620gukwYGPOGpzDGgpfolvKAEGsPb+F5k
Wj7dq6FDiXa04KyeaGzWn34tqSHp9NuQ/6LGm/wH39dhGhavqdQic5UgVonspEOA
9KyWwWKEF8tbDy3YW1OrGFNU09JqYDtoA9ltjKEXZskczTbnx0HnFB1NuydEWz6h
u48XjxJLC5ewkQpz421i7xZaHXv4DKoVef7iQ+L5S27p+Kp+MTTFOxAQ6Wn4+zYb
xQqspZXN+VwH+9EQisXYd7Z2gbDckq3ly/z/mrdaBmOuljhUl7YX4f9XOJ4CRGjT
tj3+DIfcI8eDb3gUXs2wLdcqpL1VGdC+JZnn5QM6cnNnpH+lWai4Be45CmO4V14a
wr0C3nUddX7SUjRxm0nTSM6rwdNG3KZjyfwW7kUP7eUmVH3H0OCOduykl2ezgIjY
aMFQJ53NvDd+rEct/IaB9S9VAx42lJ0zsokgHqXUuCCwjMo4YZ+0CMOdimns2TxM
fJJPl6xaDC+F/cyS0I6+b07jARVQT5f9GbLGA6dO78ZTMsoHabY3vjwSrnGwKhsx
ONP4wDdI57BL9GTB85sBLSG/NMusjWSXL04SM6CkhoYvLQx88MB55xb/+qe8JKsQ
1BAQ2c2o7P2oHYkCS/cIGGwicv34aSGfohDiRI20Y5FnJ6cOLO2YJxki6ppe4n3/
V/QFeynqpVFxUE8x2asE8c37SJVMUm1AML1xuQPQxaTMklt6mXapMZ5z9X/q9bdX
LwxK0FYQeONRbeDR6CsiyQkAAVg4oG3Ezvj8ZF5VNM57aNQkEb75uGWilyOCSZez
6dMGsmtFC1nsASmtFyKpo2Qalvvz1k7WtTxLsWiOGvpDYib/6w5BGNXtsR9aDeDR
pJPOnDFmlb2zYUxw0JpIsW1uJ8clNeN4iKLwNQ6KzCNhImKMo/TAs6luyogNpLEo
13IXiQEFUiy1AMcHtpNX/2lsnVoGG+cnxzLP4o1x0W8Xjn9LUvJPocKhBD7zffDy
aG7pM3fwTkRPz+9xiyifbwrI8DBQfChwo5n/MTuh4WW7iEf0g+1vKlRbxaNb7Bzw
Oq7d2KkFXLuju4CxUCic3SP1e/WvZDHqdB+U6nz4sKU6dpyEzrWQJAKUG/q8X7oA
Rk0yjflAipyPdDllWQpABG/t+QTP/P2PWRn9ApwB1DlvvX9Yacob9LpcQWldqy5a
q7mH54J6U9dkuK3d6D8Yax/5ZvGm3CprjFGY5w5JwmGiwLXeAlIUjr3RluO4pLrR
44QQCeN7Qd4ZdXE8JtnwO+Z6nu8gb6YcGSzQMk5vi26EWhYN9k7cKTgsbsQwV4eU
qP61rEg9A4Bhle4Tm/2HcEQqveHCGmYAN3IheskcLBurPAxrVrhPnOxoRvdlk/rm
EGVAmHkEjtZ56nm84DI4LeK/ejT5WVJfxD82SpOOQqEiZLJQY+EKDpuqkJdiSVBV
b6Yq+Pmu9LXWFsdXjmxVE2jM0W2M5api/94XN4b06gln4d4YYz6K1MsCuQKhkEVD
vZNufppVCY/tpUpC4n26tQ6MOvvICYy5Mnbj6kWHofsjUGs/26idYeVZv5q3GILd
xJix/RZW8UJclnmP27Ru8zLKKvILFirr13XdTy5mTSha6fgkrZNgk5OBbP6uE5xi
QTJfPQOK9Yz78OWuNb5Nhd0RroWs5dl6W3vXPqzF8Ahv5L0UaPfW+KPfL2yJxfYQ
jzwy/ncnMkOvzZ9X/DHJuFULVjVgfb91fCSrhOvyx2BviFGNncoiuSJrGdWkK9hB
JXzZZrvjD3O2Fq4SSN9CqiE/9mbVjg3tNAMIhzvQlXHIL/U9IUa3xo0IeZibzJkg
2d7PjSGsw0wAltVtVCLjt7SGFiTDhBWqOqvy8nEzb1LYnAjLWuCgjc8Z05eC0U6r
ZdVPOJMqSitY/gfDdUTh2ofPfr7fs4DiroCDHypf2gOrYOBiQQrqe6o+4Mr1A7fp
muyASYjzrQOGBCGOiOlQCpjOO5szA01tLOz10tVCY5aSvJbbN/LrEsKLc3mMkJ2Z
xkDElr4kxQT3BSb/Nm+fRyE1tiqVdqCuh66V+7shPPP27WdI5CD6Xe7TJhv+vddO
AEbEm+kYMWF1YM8ya5K2qchhYUnorNqb979NPAfLXhYQy2loCPURJ6ZM6e8oQis6
P66BU70kzkpc26NrQ0C2sT1KuAeIXHkdAUuaiKCnSE7Bq34YVasindTH2LtHjEx6
hNa7G46cv4x5j64vNN0jpwxT5XwjXxBiC3mtpQxGddQjo8CagvqX2VpQ5/PO+PHX
dEhgAUAq0K9l4wlVmKE7cQ0HaNp2kY/uEGRzKt7/wiJ+jUs/alUKVSVHjsQrxEEW
ZwVi5WgsAMe0AcYIHWipw18w3W8tvwz05OAZuQRQlWTFVJzNfsz/eCK/UpgajyjW
tRML/Dp/CdQyM+HnURThZctL8TPgVozW9Pc23+svQayARMnHTpK3hJSF7e2R8/42
Mo5cRkkMu83G9veLnvHje17aHxv2DxC5rSvQuqOUkUhfMM/N7Ce8Szd4NkDbC54C
XOw4Y79OMH3m7vuxsTTjTRLgRNwejOcPuhRZFhe7ISSsS1bd1ZbhPRwLkLkgg/JB
SpHfqT6YEiEsZSVbSGzexL2ppPedKLdxz8NaeXNpjFX/o3J/qH5tjtVNnPw8j9Wq
YKBECVEzb/0w3k1rtyyKTPA2Jcxmfo7Ss93/B7itNU1SWSHyCDGVFYCL0EZibYAf
Z4Oged6sfSQz+HS8jj8D9pTEukAzkctQrLVlPnBmnTPun1bfTxp3A0+O3V/Xk7Za
pM9DIYVVk+HEfJpQG7tvmF7El57yJhE4l59fxmD4jv6Yf7iFR3guEbwWzV+KZPFQ
aeAXqx/lrE4Cg+9ledLu53ZukJYC+sZ1MAVk1+B54EtsfWlj1nV50JWMXwdsAowz
MG85ZZctm47nW1U+5R7OuiEYkSXHqJQMgaDh4Zk2c9I3HMfQfwjhaku1QYDpxf+/
XDBZW5P3VpRYevjFIpcCXfggXJUVRSZa/fblWLOa5Y2xMO6TuGyOPtXdCC3g/pP2
9aujkhSUH5MJyTk9bG2JsF+O86ElwnxY4/mkHZDQ5mxZUQIm79++UUxADLSIqGU7
3X6vH5vBySAgil160gCHGBdLMeOboR7B/t0r2HmV5FXb2VFSuudQptiXPwkhHXwV
j186yrRCykv9YFIr/m2z0PiYYy2G2/i2Pj1qPhggQJd2n33fPw+3KzAVncYfL+u6
QwbiOuC7WTxZUaohZoJPb9FE/rs4SdlGn7Ltkfb/4mS7opuG4nZkyOehuKHRBab+
VRU5MMn8QIjMRNputzdsVoxW7G2cKPEdB/VAjw2zJukdGK7qO/ApvO5iilBubhlP
SGhmyRWa+syh/wwCSL7BLH6R1xwJt04fC9EPWPIR8zKXzc11uryk9O9NK/N2Z5uA
G4JgkUUPTYEEgxICMuHUpuWE9zul1c1r7ZNPPIQ/TUldBsEjX9UaEHimObeoGojy
XLY6C40cQnJAerZvqBoEcjwOMEAbqZAq05y3CFbSgByv9V2QF+HxjjOiRiQjP1GE
zrsbhTCCTQk+KQS20j65EOtJe4mBEI8c3O04nA895oEo0rpyXIx+qm3w/+2JkcQI
CowtfzHwBD1pqKOfmminu6FVemKXd0PCx2WIIejBO02/VebDRKIywK6sOn1ewIrk
y3KERusi4BA9Mk/qwh/2rhc6g55BRsSt7B3PwTHnq32oXhpSDbPhMEG9/HNINUAs
3xxMEjBynOFLla+o3VGsgVhIwfZoF+ale02oSccIplqaaSytjXzslQtd6E5w1Ik+
/vOeA+4L8g6e6H/zDr7LckpJFrOYFEN6PT8PoRoPB6xcJ7ILXZWU3mTuTq56gfzf
awYsHRXouMownJsZ0f6Ue2FlYX8P7QwM48qYrTYT6qjqgaIBKKvi8Oygj0u7Lo+b
Rmpuzd3mNK0qedt+P/qf7upy87WvYf9GWhXFtKByTLeLn85COYlrGYcm3BOUqzMl
ikBJJaOrIGDVUSfvKLZsbmLB8lkGKfEr59t9m9uJTs9+rvcqUjAcY+WuC8K6l58J
u9/hk8rU90PKFXeO0pFR8sMcQuRtc7stJU0x4UF30AIhckVZRGmSE8DoQCsire7p
D9Q1rVAn1r+OWEQfpgL4+gpkTMtMhweA+WDqMvwA0RFlBIC/cpDLKU1zY+Rfamfu
HC5wCx8yzT5/eo0zDuDS5MECm4/SeVkyPLHGKnHbPk7c4PC8HCTPWEMMBEl0X0dk
tjzHVmXwtAaUP0m/PGFTBnIg0ww4LBva2aOKjLmMo2JzzwDfGUYC7xzPc81UY7tW
GIF7gpOEQ+WdJ9KWZrzRxqITyNBJjKIjC904OyruVmRRriJ3a6M+o0xCu+TWHeeh
yafF0PeQt/JscOhReLeBTQfFjCyuJziFlnC/N0l7A6yV18hdlQA6IKdRQaMAux5b
IK8sOrPX1QWgHcBIrWh1+qDzUiKXt1ely1E4FYOyQ+DIdcwe1p95FLaf48padF9P
heVndDQjcEkqGUaYA3HY+WSo/XY5Hw7rd9thNAy99vZ5dysagwj7Ht4EAG+P8+FS
96Luz7QVPi4VLDWiFFDifov6HaRfZqK45ZEgcN4jPBHPDLjOH7EkikKY/PbQFFOP
YfiwppsElZnVn/n6KTvyi9WaqWB0vfFNH9+Ip0y+dtevNz3x/cAlw8jGJzoQZKPQ
zlY8/Amp2D8TxPbmaSvcJ8pVm0Sd1uimopCzqtWvBAAzV3+1cy+HWEgM864oa67A
7WGzHWL6VD9NdB3XSJOtFsGKKrdxJHbiU3VDHr/075UQUBU37pV5nAlOf8OOXQKn
TrivXeu9fXeraT6x22aUYMCcQZry7PTxzU6sGiibAo+QwxPqFgJYizuR3r+Z6o5T
l8VtQruJqfj2wDCrnhPNSVWIGSxUM/1ZQLXDg7Klt855uu0Djzr+42E9nIlodbfW
XfwCOjl4Qj4jwQ4dG8jsjGZWi6Ay83D9pgYeo7XFI2fNoPjWkXB4MtOS5mihCzQT
zjvX6Y+hBeeemJMV/pZeTpsTfawtJWajacaCZGnEWaXKp7h1hySij9CANKROc4gk
H5605/019oXTLgaXl+70yAC3XRGu2b5d6B03Cm0mlVIVHnUiL8mmJifeHMNGkCTi
qc5mkcAQntMoH55pwiB9Q7Fvt8IrON0MFQoJwGpFg8oEhLjIUPIb7n0dMnJzHpMl
qmMWeDYE2b+b8rqdHI6//4RsQdwJHphFHLSyhy4eTVYbMcS4/9ktrAhsHWqqDh05
GIcW8ROEYcxe1xKbuIU0nw39SqvYmq1qFnG9f/7iIMbu957G5MyLmOVLVk+OBzOz
abnmH2NSUh1lcYaQ2L/08CT2hV8N7yNI04NWrmEQfxS330i950KdVF2fQRWQ2eWn
Rb+XQs8lFXH3Dyskb/XBgHGmyUZjFBuClWabM4rwH2/UhnOuKSfXQ9E5uNGUDmWX
DszfIhMVJstptp/X765pbWJrIXV8GI0lKP78XObeh1MK4tnkwTIODOVGfRH4s237
sDvJoDHO4uBTdAblHbm99J8ZHPAig1MxHpnocA2Ld+T3ULZ1Nks9rHDYHa74BkmE
Q8LH2N8OzkrLqRJ0eELyOWvHz6RSSsiOipRef4t0AipDFPI/Od2EIVbYw7sG4LUX
S6ccCY92ERVA2OUTSlA58savljdjcrOzoh6AzQOoy1OyRhFXq50X3JQm5sUGtjTe
9HNB3aSiht9TFvZmvp6tdceUl0mzSNZxnleMwuUGTlf5t+mwpSNp4P3syk0DNWAc
SyuNsSR8AsjWE+k0QsgvRv3X7+CTTFP6uNfFnYn3XR9O8o0LP0to3gfb+KRbar1o
mJkja5yCAITcrr6Nsj1JQnSxy3jKu/ddqxUG/cSnH9SAG34NT9vkc3LwwWbX8IJh
6nWaBiANUyzlKgA92Y6uKx/mmoJPxn2pzt6k8zgJ9+mCnGJOTUxYyJX3bo3mE2OM
/9pTazuuYxdpVmVdsszubfugG7CKhH5Yf5MXBSR1FT3FuJrNgH4YiPKS7HVoELf3
fvy/vXzqGZAzgR6lX7U3k3mGweCF/neY685R5Lvfc9sHWc6pAZs1SeEEcYCihO3V
/E7aXFwrRWePdJhp7NV3iO8NNwDFtQ45TWrDY70nal0Fm0gVcNs3v6kpp8m5Lelq
1dBo2qI5IPIbv9eLYIpjNple+OhIFKnLgjhpDq8nuqgFS1174F5OwiQuZR4Q1IqS
hB2W/OGBOwGk55Hstlh63tObnnPnm6F0sI4tIEhWiCz1tK5SCe+dr44hrUFB48PI
UczxEM8FFVG+eIegaC//Uly05qN5SUeP69XjoRkQ+8cy9GHD9awLcnx7GSoI8g4c
uUr+sWXs/nJN4wY343hma+oFaWQP8GtACUAkBX8JflTGLgXKA6T5S1NgUXDr7Dw/
rOSZwxSpBlZsMk10QhlXCQ5F1BsSt7F5i4isuNhauifgzT8Gg0zOrSHprODP6d11
k6AZrZfXW3Sb8qb9OZXLn0r3XA+/Rs78oAHJ3ET8E+6PxC2DS2DF0CPhUZxkzzqN
8BMWplaX/aVp2SsaZJ9cCHCbDYkb99+AqfHla290Ji2I3L+r9GwZeSSfGDFfelr+
asfrPI3cD9Ost+WMPHFybzQbhUJjyUIxrIfNs4Bt543VMQ81Afhoymi07mzwvFfZ
crsaiXvfboeZtHW9cm/jMWP/JE/MwAVP4IwM5riT3v3RZ8XY1Glk96r8NmHjVT8w
BZuN2Z4Zfsff+PEdYlHC5slc2DVQoO/4y21I0/Byi7C8TztQcZ03h9qUVsDqAkwG
F1QD6W5odT/utSOcHiur1FVvrUHto3LELjlhvq/bk4GpeEh4R7I0U6bwjkvLp8fc
LPZKvaFMS1JH7s8doNUMseprXhtVj4G7XyYCtxsEDcCcLhZrmJI8sK7Wl9P9/Ode
Vly5BaMPu4itLb/Xp7L6MlfKIHKQ3FIehBJB83kIQ4rbHBUzYhD1Uan69O02mhhH
++r58JsyELJ8ugcGFnBPsTv+DaOkYon4lwr+YYqw78JTF0lxkj3b4kiDFmloRR2A
0TBan/17T8FTSulz7hlh6f9QgkC2mba3sawiaVJR5O8SH86IymIIrXsgOz+ocsVw
XM0N8S4K1O5SbIYIDdQKr7wHyKhsl16ttaUZ7hmCrFYBVCOgrFFzsQb5sMJscA9G
Cer9XfQ7SXaGrjkp61W2Y08WZgXNy7xxeefvx3RO39JJ/SbPnv5MsfeirXDt8Jrs
Q85EhlVtWvWYWMCaN4L1ow3Ukz6j7gVpNGzji5BQwRzFBoC3a6Ru7l60Sashld46
/SPjBwExF8Ifa8GWp5xzCocntU6YIo92FXhMD1n9aiim2qWR1t19EUKhTmjZ0zYM
xBH+CNjur/rMAGBWiRtRd02O9rZfJOjMuuV8nQGCDbMhVGAf60D8UoPGMGr3VygX
k7opX5LsPvjdSzJdML/tE56GgPBML2x39B8menNorDJG9sgKCEsqGgQuqZrDdUef
NOOfnLli7y1UPrVR4YLvCdTsVEBqZejTlIFVRcoGBXSvU0EC4B3heJe3sDfbg0cM
1Xe8FXN/XXwjpc0ZOyUg1PeB3dboYcI02d7wzyv9GG8asQpDVaPM4MJsamMMK/n4
6p5z4hmrcC5BJAjRzpHb43/1afXFJ0m9dvd3A9UH93SJrZs7Zz2HW7SMyFsof8X5
O9wzlYTmwOU/hyE1IUSampJnanzq8cSmcxllUhw7+UGKTQy+Ojb8XLnn+4fbXqJF
FZgmSYVTo3f18PKZmO00lnclC/68NGn3cn08ZSr0bAbjB+8ylmd8vK5p+1Df+dYa
yRr4sk1D/JLOeU8RBDix94ZvRbYJt/wawMRaXLHpBXhYIyRfwNAyFEN76VnKZZOk
iUHlJWqaw/sZPfm7bQC2zpgFfaRrgpBKBfOpuRq5aqngW6FqqHPIofwgdCTj6p2/
W6YEXupyEMvxgcWEbltYrAcUzmqbQ39xkCN0f9QzzrX7dBQro32DVJ3gdRNz6ASh
648S0IpdtxWydJpkuMLg2QesiMrHYE1jfk5p1lFasZoYiArkHoQ0rdkBJY1xdgsm
09en/4VbA22zg/AM8UCGuGMsctLFVVujJmxnc4MXOiTbj6npCjYEorWGWExJdch+
HO4DwvWBFYT40Qt0G0HccYcXjo15KYamy1xR/BpmnJP5TTAELzhxkqLDA/hIm3Wg
S5yV8LeKJX4ORsYFYoSykxleiLVxXTQQJoV6fdoZFGKzRPX4k4h53CX+yEI1wczH
2jNWsf/DIw/cv+Sr/eUFL7ULos33eKiiZFgHAmiWezOJKnHe4HC4vp+Sx2CoX7WD
dkhMzIGE7u6979K+m6QjAAg+YXXMj2FDHzUdvANopXEASh4dlMv4yFwCur3yCzxU
xAi5xQcuTAcgEPRj3yWjwU1onzhTmQaqXvOwdCHXJ57izAag2YHPwNCkJOmiI4iV
16b49tdlfjkEGyDy37v+kqaYRH0+OksXyhkjS8xx211Wfjlh16Np6KYWUwrtHbmE
seD/C74k9YSI44qX62Yl3pJanw6raAHV4tFrhLTkjf3FoyRgjBrLuI5hFgsbAt0A
errAPt4WX7dJAvANxMPMmyxFbCLrEmz9aCxKj9qKpUp6nsxt8cDHSMyyCQd8qWuV
ySI5gYAxwkwcwJphG5TZdj/z3mxwAPMXldWJpVei2YtlgZEAgtAVZPY/+pZ3SNnf
sIztBruCqWkcZv+2Rr43TAWWhxcqg30xdg7izL3eueIcRCCBBLERMVVmThayZFg+
HhCYdFHmOUrbmt1kcqowLMgFCmkLOIpGTtdMBOqlC+rTJ9nnmhcvEneBNVdu08bR
2LM/yUls/6An0ds2JXj0V/QCnF3aiekPNQNgujEjdxCYq8xvxN6J18jsVDwrWqzA
xVrXIAcwt8DEJ4VGTccwARukDWYS45+sbUaB8OYI0ZSptWPTvptSwIKPLJwu+1U8
pQgmK8QG4jrk6cZvvYJfFCDH0IthYIEG7IewhPtGCb+0kgprbCILvOdyjPeB5uPC
2RaRqcbeHLdzN/uVcCFiFwH7vRPvIbtietG3/3YzV3nZEOOrNmBBAH2gJBFwcSXE
68X9GWnj1f6YLY0QOi2mbLb8EFFwRn9LpfNfN+HKJ+zIVDxSiodIaAdeXxwtbpOV
u/b8dZSiksJYBHkxNV8LJGVqsORUWGNhTLxOdo1mAHnJPG7rH7F6qEfXh5wIJvgT
oVbPklAY8cl7OZadJz3k3v10aTP5oJlhobwI5kjSe2kb7HQPC/u7BxQc2wZ38ON9
84DJ81fCIbwZ1gG8ZqidhowKjfqdKxsGa0LfaFwdqfJwt9V9MHnJQW4CUG0G9j86
bd/miZPRXHyJ3dBwBPmSj8viyJOhGtlrazfIoOr4v/mT9WtSPOvh2wQ6FN4jmo3W
i6daES8Z8JI2LdxKYeiuL42BKXkGKw9p5PgKbTc5uFLE3OiGF89WbcLquApw9hbD
YYsxYWKV9GokZK2/JmDOUmwc/PGH3WOr7UHI0ivaEReyrcfNaeLh8A5XdOewYPq/
3C4wlqHXepcyH5vVaNT5OFwhfJRojaxLr5mzgo+SvP0WsMMwqT97eoeVOT+d7fL4
EpUr7HpVCl6Tmw2zh4lauly0jhjjqKNqufxUvmmzAVe6IlNRydwJDuDvjOUQ3Fyv
jEmV/H2kJdOM7LMWUEA+5hI0udalD0WN4TNEq1plh17wKWxq7klN0tcReJdIE3JN
f9pkKKxZb7r9rP78Tbo1WG3gCm4LrytLA3A+nTEVmMshD78soveFEoGIFLVqfd7+
1+NW1LFS254IihKS2RMB89H3fB5A8qDQ7PlMUEBvT+Fjd/0QvHS6RRgwRolj4Cpf
PFFfXOOwFl6t5z/AelKd2ahgjt0c0gUijZLgv7gBrTO34P142bJ8nOGfrjvxxtw6
JFsZsRKwaF4JJur2JQMrDSXX1t78closS0OlufjDU/AL2MaoHmwb5ENxCaC5tI5D
Pv3rhuGI6ZkUx5pF0amrjudOCsB7Rw41HB9tSMXslhzereB3d9zwsC6nRZsovFFQ
kHGSjgbadcBMSy8yD0pmb9Go8c0FhfYKs6TIQikMtjmZ7vA/JdgJYoU0RpY4rejx
sxj8dS5J8F45z70v1oUDIZCjGUvhY+4zK2uN5mKFM0iERGhKoVhUKHp968DHMMsn
QIQNjCrxFUKmi2CbHhgbLsY3zvvo+r/UjyFtF3353k4j0QAyI5iTaFJWjoYfQxxy
CoL5oLknxjaFs9g+PTFwSAlvAVu3D9zQbhYUX/y9RYwZFmmMxzt4jO3qf18Qvnpz
FVmYwpkp2lyyMccPJwXPKL1EYByz6LZC+P01XM9/NYG6CBJUn1y2sqiDYm1v+Aaf
kzVBKfGMDogfAZgGXl6ujJROFGRufLncXxSL7T7KfMARy8oStrEQM2eQIJ4bCvW5
6c1XilHdhLA8PpHZFCN5BxP+a4WpxX/K9gNaG02UXrS8Kx56bLLodtAYn6lOMSDi
7Rn4+Tn+WDpOq3SfH8hXP/lmzg1ymY0Vddoeknja5VFH5Z5ztApGROae4UOjjdfw
shUqSwH5W2yWvHJBDjbqNUWHG1wwLP7eq9MdnvOPtTMdC82f8pzmS4fPBbuR7pAX
is1R6qaAMnAUAPi6cme0XiAWeFiATjWTKSjEvirk6Zrcjrf/qQjWIR4emlFiQMT2
VtfuxgkeJZun6h5jo9fkJby2IDHKb/Kj2M/E8q6gcuhNsw8RMJ0KbeQkhmONrIuV
Pl/Ii80U5Xwo8nGSlWVG/+qR/GczKrYFXFQ+mdN0DuqUvtj0N4fSZ3ktcL5Vdh2Y
MwbUKexymZMfmbKv9HJflXqOmtmfbVUfUBW73noF1bXHH54/EpmS/oqjpyww4Dpo
fQCpPFOeIckXI2P2VkDy/xYpzcFpJRJJob/EB+DDLC/U7ffaP9rPcrH9zAtq9nZK
qQlRX+U6eg0cdp7112ao1139r2+uA49PunsbBulDbC+kKoyZh/x7Jmywm7e6rxfD
15cZppnnHdjg8NRTxA0EAxfWPUPxbvXjQMA7mR2kfmdh/FdlHioeuCTR5HozGtrA
MpMuBhc2Do5xvSw4LoIDeoM8C/vtwgTKk1IB0s6XPPOwIGceA2/F2ypjUDPqxl+7
A1tNHMBJXfVPiC3MC3WSjiwwhdg54MW9zAkkWDW5CU2v8Cuvp4BNphOSiY8k0o45
j7zl4zYtOghP0KyrelfMdM6wtv15s9G4qrN0KYrRO06T6uyubl2qqMD4YExKU2oS
gbFgwR8TW0o/hGO5x/y7BlaeP7KYwjKz0CghHhEwNtqqW1kNNNJIUUkCBoaSOKCR
JE1eP4zU4kdAdod1Ulx4MADWysBXMPO3I5PF+EuH9jfbS6sbOWRdcK1LMZ7qQIvi
KupJn4CYgFmYfpF0CGsimDzKfOQ0IACJ01cssgDYvafZBXlkz8cAAp4gZjOwjVnW
OahcW4CbrSjIsFYsWsjCpNbvKhXAx8x6lw0kLrGkgreyi+UEcf1qvfDiwj4AWh5b
A8HISvd0JK7dhoE9G3QH5jHN+i4csaI+4ePpfBHmMJ8JCjgkNVClnHRUaM5i2EeW
hthkNpyvdXZasyUTTUXjoCO2hZmSJExc0ibg8pPBGFTJ5W86WgMyfOF6PueEeoTJ
EPrIyE3sAAcLC0TLkI9nplNuv9JA0uIrvY3J8OS1Z1j5WXmARY6reJQ/jnvI8MLj
nbAHDp6HWrJVSfvrWeSOKeDb9cRH6a4CYqmhdik1khMXMyvmFi5D82WiTaMFyF1G
/s8NU/5+2puoxTng1dfs1ki5mXsr/goP4hid9hTG+hVtZ67psBb5bR/6wQeho+O+
vOzEo8+tiJCKnw1o9uPho38Yz3Ahk6O2s3msr42J6ApZ46KPNeiTEKaKMbyx71mS
xUW05qyuHjzL7nK+sXhwpSZLb3pXnTUn2Asflu28cxrXfHe7k7ew3SdzGkG0WVj4
4WOqVX06LjdNDr/pjPqmvoF7JOFmNOsDRYUrGQMGKXf1EHHhQjHp9X57mXMfDZpr
7+Ju0OvdeBCLQhwIIDht4XiUVkwM8zsiscsoyguWq9xLhLb8Nzc/BMwzmYwgnZY9
mBhoprU5/0MRpdPzEd0eeOo8zI/wFgg8BUbIua7uwU1BGYZW8wfeRfrEUIYuX0Hv
GsPP+wwHe8FdKlAZV5nFrlZJ/nIKQdRJQ+psTOzRqrv0TS/F87qeg3qhvJzh0LNf
K5sBIxantVBB9dNtmvw1Oy6LE3OVBn3xXqMuuBhHrRgTd5EgsATGOPNrjDagyMWX
7osJFLaV/QjGyOzItspV1I99BG75eBsnxXSe9e5Txvb5aNwma59LCIt035QpgUxj
6vWwse3rRG/+lRTHUPVRCkw9cSfuA2kEI6JN3KkJuhOWvMoIZx9jrd1pFxiofh9E
9XiQPAbViS36b5TEvHuVyXpaD2sy1lz28eiS3O/gU6eiAcmfrMVOBUyI4rshjPSJ
WYql9l+SLnUcHxpr2R0GTq+77Xw+5/R+7oZ1Y3/xA5wNmIufvKNotkq2Z4OD4hk5
6Uw1Oa3GhIwSXIYjGA+Q73dT/xDnX+b2Wiu+Vl2/mxLqnZ+UoQ1nLz4eeoit1/tX
FyGO0Avxb78zLC+iYvUGwgsv7KiwxgvLL+OP5GdfYVE/iGcHMeOmiFLKAIK5N1DX
vDkguuAQdkTW8Np2SvyCue74J6AZnAifj3apHK/ksiXQ7n/2YkT/TyelHa5LbeC5
aIID8sCW6Yxp3BZBf3r9AEg2T2g8egZwaYpGyeK81Uf4JyYJfTiKDuYfmJDad0z1
9Tmv/kM3luVukPFgt/pjWByouf4rdZcr+xk8A5q2WCFEK5CPaURO8HPZ/jopDLDB
BrBAQ1OKo6rCQvgo7Qi384cE+TpbqpZ2+PDsicwzunyUrNX7bxWbZH+1Qjb2hEuY
2k8JEaa7NOoaqdYODSs8RwO6vtNjo2vrhKye6fipYqRjtawpdQxegTpUuE1zYdFt
UcuwgPMOVcHpDx49FPk3W9d+C/eM4FsL76ms34O3yuRpFHQCK5aRYFBHFp/2FfQ6
f0rn7ZtEfzbH7SbEKnYiaq/E8PYBXXjmLepoBP0qfUBihCPyzrurLzxitnAtGeku
wUKPmwcmLNvbvkk9JNJgX08ivmqSMVVCmHea74SvVInOLjZLo/yXn1XknMxkb5J3
r4JIyN0j8N6MA25OrNIPI2fLlvB+GX8griSPwb3fbl+jf7SmLYabkcJ4+WMEa0Qq
lJHuSpCyoeiPgutldB0udrvzj/asdTYLDTpn9Vb2xYmNWv2UREkTZ9tWMu89QOoT
rc77seTSnqc1GR0k6DN5b4/G56oS0qXPcItEwXLJz2pWYt265cDwFtJPNrIx0Dmc
DDMSXot3JQs3gZVPpjfEmLnEGVHD10/9Wj3Rlh7VLnWeOxN2SPNypgjMcDu8/XjJ
kK3COUtWIkuhKKTGPgj394SNvm6phXyMvCjhUbmd5rjJUNRxDvlGhBPqOc/K8Oa2
3E2FU/sEf8iC0A8D0FEkKD+nKgjgOxUdWg3Hjv7232A+cC7RdAcqg7LvuRsbVwU+
rC47J2I3zQ5rOz/a2ZtABKiloTDPFJzBBsBNeEPriSDjZYN1Ts0RLyKVdc/mkbY7
qiscZqqFKpvWrWtGsAhp0AWonvkFzrgWEEUvxBV3/MacSjpaOApsPhJ4+XhUQwNV
Io4toW2cEXmRu390/dQNkGKS3+776coImVC4lwPK294z9eivPyHnjEDzxZ26A8Cz
BSn395Ros+ggMV16qQbCMBiIKiZ2EKEX0zqDlPrjzd5GU9dGx3Q7QrRfO4xO0+Nx
JTk3JYBLbzqKjXVinfdSmHUX2ME/rlx/bI6shAXsXNwWTLN1azwKlOrziVSv98Qa
noEZ42jb31QOQoMRMndDqdKa2igDu8/qyp5qtJ9WahNsjEDYh+2y4S7nf6R6Em3O
YrH3X7hF+Hie6edxBa4dOZmNqxNZcNyokk0vaKJnGlUt8qiaba0OA7QbpteYXh6s
S4WYowsrS8H/vouyJac0Smf4S7JJHlm18CDK0lPlztkyVdytGh4UIxwnxZ7yTR63
18pj+djpKrU9zo5Wahc1fe1BaelOlN6SmIuJY18e0nzB7+z404XTYlrHVnMsSD9a
/dsEFDw4HBa9wc9EkBWubZvX3fdW1R0caPKiuxK4f8lyGQxPgYFvJqQAPB9T1sqY
pte0Jv/74TEB2IEG2ymMtnNhwV0uI9y1L/jzS4T3WPqq2wv9rw+Y9jNl2IR5ObAS
Fqx7EcNYaDLmtD22rcoo5FvvvIcEt0E3SuaXhFfe+/GRjYYXwAx5oiurXyUPtndN
U3Scq2Y/DY+EZVD4svclqhrsgWKP5sANHBwGqCClWuoSNT4AGlZCtUMhOxqrqd3G
/2b+Jcu0oAaFoExImpOg67ySZtIEHwQ/4u8jQh9ghGiuR4gBUQZEQCAfiM5rnW1r
SQWqZKQpCduQKI7AvK4W+Ofe4PMnfTXsil/5zX1ar9VwfmXZ3yyTLkAbu9xls+9p
F0T2+M1CcuYSrTuFzZ3A1Yjxa+mIatWuOqHHSGOIIQPltWR26xh/cA7HYPUCiX31
VvagM2RALzuHqSmQwwjYeZ5lD36jHqWUyPG6PWGscK/sHqYic7D5fYqZjx2eVo/c
F4yuHdLPDMuq3wWact8yIoA7bjGv/tQdAs3Y0Xeo6xwTWOWIE51Kd5bzwpOuncAn
27ARNll4+3AyxDI3DM1BGmeOg+1r2VDQqM78jRatdLKKCX9dHbB8MjRCTfCIo6V/
9Rc1ZPYJhLFCqdGea/PsyDPIY6UTUgh63RRmCHN+M5PT3JypuNMKrV2C7QWffVcQ
EdrApvZVFfCqqWSfqJejKo3kpVfwwce9qPzI5ew9kOuW0/w3p6GNWFuvJvf3h9cs
CMYpqjjpchlhjZhydBuxZVsNWIJSpBAzEtH8zoc64+BH+k0S/HmCu72Tj5hGfh77
4FCH+fNtiuuAH26MKJy6v2o0oNuLC/Y2kBnoo2gwmlNcKgUamni+rUEPGH/Tkvnz
oeg38ciNG04uSRQHRP8Jf3qA33IMvUrnwyQI5ngJFRGq4TedWbSJJyPjxXSllgeD
gR0fW2nid/a4jrbHQvig17my01ZB89NW77xbIKjQSBYj+yCih1J+8RMMLcAM4L8d
ncZV3RhpcepdyLTZb3mzGYg+oo2Cb7J6xrLsLLhGprhHkl5PXeUZMwz2RFpUTtp8
goP+QXiZjsMwb4abBcN61UnWQq/39Vl3kIGO5MjsNRaD34JgBoX9mHSdbE17LTLY
P2FdHV9YZ2oRYZaoehj5AOqv1Zg7aRCZAUqrGqh6tjX7CDR9xDRz+z7FVaWcQkWw
h4SIZGQCS5f1yCBRMvjtYKA775LBUbY+6oxpf5IygBN/Kjma0AGQInRfnVjgam6T
D2nKDh9bHqMGwT9C4yhDzPvULAlRlbp+nne4O+j/pnr0tmygaTgwC6+ioG7drA2C
8jpC5cHlVjoV45eMI3Q27J3zjWHlnxgb9fYAKHnCUMCuIsO0REwB28bKr1WUtm8+
tndgT2Zyk7DcD2uxogz58JdzrLoV70w7OBBtF1/RLJj0Kd7IUkuAu/QsFF75QxW+
4jeT1QcXMzwcaQFKj7HXpnGq/nqdT3LHzsyOT9pYSFp3T09VZ2g5rY9AcQvrswKT
vVs12zpOu0L8ePrJIuweUKX++nFm/cp9ITi4WkxG03oZTxSMtRjq9l2TtvXXHuA3
HqCqwTIvlWYfrWpshTIs4sF4nS2Qk9Nfdb8XnwmMxAd+XAPSFT9FXOYOVSj9TTBH
iKOw1kEFB17ctgyEnndRUrw/ToHhrGyRw2VkkoSVmJABH/VfqVn9EUTQPdgqV5W+
tsMThdNT0QQz5gJ775yK92G0f1uyY3KgVP+OQdGDivltV0Y5ZM1fZpWoEPx2P8N/
ybxsF4U3PxrWZrXMt10R9FOfuntOWiW5GKNG9rmEYdTc3d6H6Mmg0msvyMpMUWy6
WKqBRjd5AqKMzu61d+rMz1/KtlYbedyWxPFqvUq16LKET8ZmH//62zMfFKBUzQlK
pCuNTuMvP+504paPO8f2Y/F8ZxAk0wMV3bOtgeoUJUEC28zBVusD2ZT0TF8bm7hE
TWjvHnvv3FKJoBT+xzn/GllQXONac5oH5vQobbSDs8jV/yjEkE2MaP8WytASSszu
5OWQmrxDnj8ChfK84agrDvPhgIpJx9CZsMUY165g6YcjyL7G5kJXIvStzLO1itzb
U7XeZfGKAFcoIssqL5gCuCOKHvcfIv1V4atdy0hXR04enKjaYmeIL4k12g4IlUhF
e6L9lqC8vTDHrQmRM1G7WNqt4T63uTcRTwfrwbd6Zdsm/PkIJsfvqA8B7NwBBHuT
InEM1pBMtCLCVShXShbZJ4aonf1GvnGlRgoImIwy3DbjZxJE8wuEYcRJcN+1HrpB
KUj1hLU31zyl4lsRJSPAyggJTcNKaNidSsuUT1nAXztoCR9AWEPw3k8QufgSTLuZ
KX6y/zyIukOwWqCmO7lMKa5HqGUpbPnBM3KcqcaXJrspY8BVamtBys0NCvvTY5Uh
QOoOubCrDlQahOWHs188QhWAD9AmFFyOfNIyPCIZVulWYkP6FGIb9t07YY0ga1a4
n7SJ4vnDZB2/03Hi9gnPFZtHmcJGYwVPFqlJDvdaIqpTCtU4T9iZWp9RSMvo4UA7
eZJhjXGY0qm+txlJIQZFL1WeefD4pyimKzWjb4PNwVEKeSdc/OjMwQrqLX45tX78
Yi0mTHGywNp2Z0CLdvKmRqxyCA/YlSxhpiL0X1j4hYLZaFGkpXM6uIDTwx3LAUGx
0ZEFcSDE4HBpzqlVEBMrGR21XoMZUL6tRBNyBVp3EL/LigdB0Ps01GSK1c0TO0kM
IcsjV5eE6QkppRrI0H7ZcXoOF25VUuPf5X/yD7c/uehuQMA1Obkw/s6kNBwR/15s
YmkCJs5p43OB8bar0Tcc+qiYVxUxN6oVF9eObyHtzoQrAmf1kni4fo+SbmF+htWw
GmdCxz3x3WTSuIAfEapKVZd23mUO2bvOw4mBEJ/cpowdXjW2nMnWkYvgpKmtTD1J
8EJXM/MJux77al7EIkb6JwZt6s6ottmJq2WC2yDV/dMKmbZShnvL0Q69qL4KrDw/
ch7r6+9C8d/e/KSe3HPz/nwaLuW0vLOdiajA1wtvF2bE9yhNQaEhEdTcC8H47ZUL
nhkqJ1aiYd9qBQQaOx23+f9kDYdK+qesnwPboUIBCRUtnjBXx1pFfqx3YsS94PLw
s3TjaW9EymIqynpWqdpYePhCJYawj5EWVdUqP9ZH1w4MY6qhyLlvtN1FzdE0u2IT
T9m2ZQIQnXzjAmSEA3TQxkAoEH7TuUgX7Zq3KNuYjrUDSvNnWKA0R5CAUvyXJSIT
uDdKx5po2GHUcdLfOydt6X2QSbmCpx8lF+EwTrqs3Ofit2HOWPhJJlHLe07spOuc
O9d0kUvLNg6lOlDbZdL+ZMrnsciQhXhdiDbWfysSSV6sjagcSTaeJRXCDqyBnis7
COY1OMT99hlr/vZ7xlps04eUFnRL7JeeC49iIAef/izP6ui9zTlXXLRTm+lMk1Z7
ZOY9u/MUEE75HLddxgSMXMS/Nt1PGdyIt8f11ssxJE/4HXwW4gS7/e9v6p0p7tZh
AJ07VNK7p0/ej7/IZxfFZT3jeD6rOpqBySBrNstUv3KZWKiRQXdNi4ohePgG7E/p
H4JCSigxWY2wJ9arfq9uuyTUFne2FIWcRqzOsR1om/X6XKXcLrdhrsg+/CcPD/cf
nDAhXtv0LzBCmlrwPf7s7T1vBGO8W1uTV4ekzun/Ifc7oR8puEJi0jNi9dAzZ3XU
BIdwQ9nALQdAYgeRfl5QwNTcoQTRKZRdjO0kyhu+4OG6myIRSIYv6GYcv3JgKBdD
dAaHWS2pPC7HNfOzjbvlTdG2MewzrcrowyniZPmnsB3+ZjFGEanE+1oeoJqPpe6Q
/w+VFrFLRkHmiYdeCRNXw7S8TCkTyR95qfRnj8Bgijz2x8LvWqTML98Ecduoki8D
gq+i748+KuA953A5yFL/Lw9GqSn6qZfsw1jVLILWho6JSq1GeTHqyukUzFlZidyY
pXI7oYck/iEIHDwZD7KXnaYdxiKpdzn8ZNjS3Z0XnV6MRueK2likWagZCg1eE1ef
qsTExVpTQT7dCEFCeyJ1s0Nge1oke9tjEbsOqadfdEdEXEAJUJ9xLTB0ui5/xLJt
Z/2YDcqzlSDKbtrXhCNVvrza04q22ZUk2LoBZRokhTWhtWHAK+0LZ02OFsAt/Uph
nt3zqja9XW7YYeu4BqSbLh62f4tb1zmzl3plBoZt4r5kqg8SDHDuDQnGQ57hHQcT
GZf/Lz+/aHmWdwGxCrMm5/GgCx4uwQuvvWlIoyfDddJtFzWBLdBLptviiT04Y88L
IxQrrQWdZwAYjUdBLS2FXSHRhmvtYz76f9nbo69pIbHiywzo0eZW0SlropwzPhSF
Rg/yDiZq4e5HolcYH9I3cqbsZrDffRjGdU0Z4MwQ28RoZN0166rZraouP3L+tM90
fOBcjub1wKSR8+OZPrnPLqiT8hfbSTDrsXabfgCP4ckZi2xKXYL+td7wewApIJW8
mOAlexkg5JEYSaRyFR72IZWaaLe5shRuPe2IRe/PsR5a5A42z2ebWY1RsJQM5fqP
S/+fdmOtV2pZJnZQBQG4N5230cPFL1rMaGMRoFXsaKG+DK/0gtZRXZgFXM4TUPyc
xKfUBFJyGRPs97oD/cQCjXPMqpLJEkVjm4BReLkk2S58C7ECIFEKswq45iNosvPW
gvYYVZpQK7R85G3ntS4CTCfZUj1JEQo/0MhYdmjTblweFvQCrh1CwCxIltYS/9ic
uopLLgyva0B/bgw8nPB11IhLYzHqYRTWS5DOpkH0hXOHUdRTVOuJnbuBDbxxpUuV
xp7ShHmekG0d15GkC7oqy7DLbUurDWTFyacmR67KID+5tz7vyEeEt0Cuj8Qgq0pf
5dOe3W7Gw2+JQTj9bMkJ8Dft8IqPFSk1aKEk+PqSyB9cgtMmDq8WonZaZmV5XB19
uJPG65xpAOQ5vbOZtcO1LjjqgWmdb6Q3a4sQuzSh3bCRLwVrqMMYibCGamtUH6K9
GYzPSeWdStdbg/4yLE4RZYhrBy7bNOeE1P/2Ge2V1lk7bkqJFoz+9heSNBeKJLSX
IkvkW7q5NW7vFqMjfVqGlfkoxTt4Di0xmDHhXeoJfRF1Rjao1r1oMl+mFAfhffy6
vOLlf4JDAFFOHcGLRczpxifb7Ob3lgbiOUexUgbhwR9ZFFvQ7k81QFS9SGmshKf1
26e7LN+1p2n+NGAxmEale3sHdiagcuJmD9rN0U/+ef0tzgBAkkCJO6RDjmPc88tu
KTiIAD8NJusfBSmQP2cfyLKFRdxJn98CebXndvAdDFYwlIQiirSvwAePjLcp6C3Z
EIXon5H0EcF+eLkVJ08u9yKRFBKfw9wdvWXedpq1hRKRnl6Gil2s8knGAq2LWcW5
JgF4evrSueN060Ft5jNiCZ9V/HCpWVcTgECuh/IWiJKcDsmv/MtRD4pyspFVfL7U
Kt5jhlT6GXvZHsNTzIGnq6L8215Qz3lVhnwtHBTFPnlnBAd0paa63KpMZB6g9YHI
7nFTjbVfDD59dwdHEoTfuvlM+oxnEYkaV5vyIBqo9wTfsEV1k494VIhjaSPruM4X
1rCt/gEMwCFdlbR7jLH4s72cZoGPQFeIGhcQVYb7ghtW4j4khjIBlJbn0bU/bMXt
9m1xYtzCCzYrbgWWoWfokgS5RqrvdH92lqIkQI9Rz2G7dGvh9rj/K7IXmIvY/L9y
agr3D1tYkj02FGW88UDBXrARW6P4SUjPm50DTeu5DLP+r84hR/ezeLEmnB59FoLt
WzOmZafqegiOu0R3VOhrlNJlmEep3SgVL4vYdPPe8QsGOGq0WiGFMag0Ygt7wZww
/LiUCkKjHVJYi0vKeydlh7HI7TYWNDNdOHgmlt5DntiyKF+/v62CirAVrFcXgHC6
xSR7615U2aoPOoBLwnyfsuyRBkaAg4LLiiIn7pu4yn498O5gpgS739prtt3n3jhy
WoivVucoNa18ebVLRMwKrEQhIEUHoA5yl9xgTOt+qKKXx+fG9kk6K19UcAJeuQgt
w0BKJqVVsZVkzTl6T7K+sMF2arj3uL+/eHHAwMyhtKcnYKQ11/Am4+yxeV24xGSR
JO28fbYtMlDVuZQhpHuUpZTRz8lbFcUaBeBImV00/GjIJCN5lghqvoFpp5lGN5xo
UYGElnv+6Jwulu4FTS/T3iTPwVeS/Dv3YjaMLcZNpmHosFZXFtmwXnaeVOVKqzte
LHYcAredqiN8+lFxOZUuE4cFmQvFlP0Soq4YLxtyXUoVzkZYcrEd4PdVODN8fJI+
mOBo90AjXP3/MVi7tNXXgzi9RFTQvY+bmUi+/sn79dxZ51kLso2QdGHSl3dJmI3S
GXI0QPIO2EIlohJvVTIJAcx1maU5LBccbRZQoyokO1SrXiPvFtoEKIQhrm2DxGjA
mSi6nFHRGGCC+YIpz7dl+1WryHTSHAQoFCB7S58PNX/pS/gnKFbEPmePGJF+Gzgi
jE7Y4UrDg+QhMhMMxB2+F3b4Byoouwdaf+b26Cgi2HFv/lWVlliAwmkkx0voQHEc
XA9bDU0DXixULt1d2tks2V1CbwlYP+OwISsfal/+gJ+GogPn5XIITXW+sLu8Dxtc
XsGW+ubawlZ5ksB28DlxX2Iboq3gc/PvwEo8EOltqKYVQUPLMWVVM8LZLbGjX3g1
NMDMm0mjVVdRztfJ/3CBMhYp0el71C3bIEmdd3kEM0gyr9eQTUzayEUkLkS26i91
TP7k4VOWoGHsLUY2n5el+SewG0tdGN/vfjzxIKQs8jlYqzCBCq4+Aekex0O7WvnZ
NEzGefhsxf9KcBpSWf4GHxy9uMIYpK0ush7VOdf/9/PiBETJYu/+GTQ/zIYwO0m9
kspUBanFUru1uoAl88NGykoQuOZ5ciKHFNdmLe/9c/lxwJN89Myi0KLTbX4kwVvd
4p9NrOULxdRVM6RGH2luwVQ5fLgt9u/BChqM0XOPKsFXFBJU7dHfDKBSpqVInlb5
vg2FPDfPVLZtXvA/9E1CHbTe0KMRPegW+GMS2zWiaqOonasK3PpuS7l31zz6SXJp
l5ASMNZzCMpcqcIa1DMlVC6SJVwhaOYcqRIvJNcvGmepRTypq80jv9+Ika6gqMBx
76g6yzaRbL1IM8KQDPkiqgJNXeIxVywLwxALexmepnkHMpJli8z7UL4aemv1mqP9
FzUIS0r89e+liDsaXZAbfzz69VqX3lEujzqaTc/TQgjpM6DhSCItY2IlUW+nKN5m
UGmbb+XJAbGMxQOUTdCcUXGFotgMzk4G0wmiwh4TqUdqA2JSgzzQ70VHbSWcc5+N
0lgwWT3YM31oC9G+Ja25Neg9DvAsUqsar/cxhAMufpI2N8qI+4y39X1CI4eRUM+2
Puw8RcU/MaJ1UvrezWubiWKQB5d7l1TNjD4yaPRRHgExulQHYU9SEvc5nzx16fta
YwqiGM/9Hno21yh07gPH3ObOGaj/tPmzpGBhwnmlGI+rfC60uwWlcovPoEVQ3yre
n3BsaLcLbCS25oaPNa28di25GZJWTxQ59+e1/piMc08FHQrWiL+9lDy5ZdeLulWs
xckdqy52Z5pa9lKqs9GGkf1FHPDWY6+6KubGYQ9eGQcQFGqXp4XlK1dQGs9iT4mi
bVsZrEJSah6VcntYp4utORZoSJd/+iFfRykeFxHAGV6kRkf8cRlz3G28At8owiEL
wQ7VfHUDl3NrGInUpKrVTyUp8vouUKGQfnAlXAwmkh6liY4FV6LqJkQgYvgBXqxL
4CLFzmcn98k5x/7XlT1dIujW2b9v2aATMrRvnI+ooHsoJcXPqkrqDZVOnb0RyENx
pE/uvRENzhXPVo1uZiYCDfU/B3PvuyM74nkE2CiE+Z7MFfsvwFVdRQErFx/o2T/7
UsDDIHfYJ57PRNEO06UlRGKZ89VFE7KRwExe2rPIL7Z2KIcphY9Gl7DU9jyVrgBX
cmSjdYo0/IbpDzSBCO0EfJFzCYgPo4UKEGBtbHIwrYOfaqkHo3X7u05ly6lidjS3
nsCE7kiBFtwF5p7pal+E/h+A1GvPAdN1TKFiWKrv3ZwU2cLYU5B5uFOt1uBhloi7
TH+IEXccLGGZ/qmCeoeArHoCuHcte1VdTmSEoXg9FGr0rssK9e7UM4FNtuQ66Krk
8HZw2n1wbU2Sk2a9958kWcuQUcDHbiwsZnrBDA2MWtA1bv//s7xmYSP6KoFFqwnB
EsQ8FFRViKB5QQ1TtHFhv02Bw3/JTdrW6BWl9lNsewwCIR+I7edXUElIB0icAMgE
Jm3B9SxFLUrk0+/aXligsZC9mPJzRwQPaAY93kFKQa8IQXutgraz7DujsijNcwep
J2Od9lX1+xmUprWMtExgeD0FjDKutgmFFtdhlqlPrjTe5S5RxhLKl0pjsRanbdOo
uLDxa9aNuKpB01bSEOfbY0iOz+RgQnJqG7fgF44q4X/xtqbyT3+yvq+htOI2A5mk
Kcpp1VvJOtlzK7Uj4uTPrkmMJtxnnjryKKiTOSySFFhQ4DOFAJFywyBAe2gOJfcE
Fl9G4FcdgvTMRuyFgCK/S4+ThoXV3hLns/xnKY6ascR5QYoFzDgoV4g0aLTcrWwH
OWXqQ161utHERQzruwow73maZlkd44tPbG+wmMJHBdU+r18hu/WS1rvxI/7yFlhc
L9wVkRb5AO3chB22l+SA7MnlewMFM6Bo/xDSCf0gvUxc/NuhbxDF6/I0jNupVez2
GnAI6+NTSdmxeItXbBYVIefZXS/UACn+a8XYdpE6OM0qLTjerK5vG9hgQPovr2qS
jdDpJCGoYKMGK/ot2+g1y8MpNYOhRWoEkGYI3LD3Y0oWBYZq9Iag6HCNe3d1Krpr
s6f1BTD8bfz9JkrZyClY7gvFa4gznjT75L5CONhWSJft90A/zhmtlnuQ4PjeOZfw
T/a/EJAzxzv1KmD3uoQWabfqJj13vKrYazFHotC/zt9FWu91mMwdPBPzNbdx8McM
aST/BKOmZ2svUWuA2hf5ryohLe/h7OyuvUwlZP5F1PkjyBASvWBF7oObv87gNhKt
M2KrqS3vdsT3V9DOLMV3PHNFn0pqN/JorLwYSTLdfbQAe65x8jy1ZjcPf/Ae5U3X
bZUQqDDFpWKs/x5wngLAlyLSeasdEimt4avkjTGI4AvpaWkrwKOuUMESvWGKPtD/
4I4NYhuFjKM0rv9GQN1tr89Ekd1m7v/r3kS3ToQg4r//S0DZNeg+6IIR3iV2H1gV
xkRJbK2AGYL+1Cq0Ki7EHjaWSVuUILTQ1gfHCJDG1puUno3FF0/SnlClsQY4OEv/
QzYfn3yXAc3+gMm7V1AG2cX9gLyFMVecILofX7D1K06lP85QBaF+9ZsFBLILoLcU
DBxHZpxSHkGhLpprvrRcCTR7uhMiAOMa3jdESAjI7XBJKzum/LYqslQAgSBo4RzI
c0U9qc37pCs4bn/eKNmCuOhL8KkK05nREcyg7O6KPatreZE+JP3kx5WBNkyEVVKG
2Qr303hrkqMJgA14erGN5YW1k5II99OISg8sPPYcTeQJ2OZZgfAd89aH591Q5TMJ
cBGWu31wfMX0vE30lZk8lZBJiAaPUfBMa6Hb4ui2ZIH7EfN4PuxHnMaO/V4lLfTe
Bdhoq00uIUT1DaciNwOcnqQnLrwMyt1MLD6iT9w5VPBFNY2vguuNm5pCAKY8ZvWV
gJVf/jpcFHa9DLYsk6RH5WW0pcmYr5WaNlU8tWe1vX7Xn/9UOEtY8qgNXuSzz7l6
sjy36S3atmjaCKR0acBUbaS2Xs8PW27CcyW5/OB92CjUZEBXAoxIJ5vTaVJ36amx
r9tuJC7m/iP1pJLEBPqdpC6ebc+GN+du1uGtH2pkRzbW1jOjoUu3965aMrpgl8ij
nBL13UWgAOcC5zZ/4p15Y3et0uzWQ7+Y8b5Fk68YUPBsTulaebCMjsPS2jWH5S4N
MiNEkE8TSwRUggGFLhgfd4EO2b9a/23FwAQUa5zBsPtNmIqOytJwFvTH+BaSHqEN
4TuH3xovfZTGSnp/FO3P8FBuTGC1fKluXBwdmqmwBx3PAKmSHJ6bb45XQopF864v
zD/AWLhrEUodVPqHl7/SPxNBb3TkB7xQuXlxJJFl1AOFoUn8gPrPvRXfavVnpfkP
UQIm1VkqWOzo6Y3wsP4C+fmwkfl6jf9E8vliIa4YHarx/t9ryDyTMzn/szOQ3Vup
KmziCwMgaCEoxOHgDnR4YX30hzgETil2UdKyDFV5qkbxau/dzqo3bxhzDZWKQWzM
adfSApSMau0iG5oSvYWNbN2CH2Wc8vp400mJCoW7HAZ8De5Yh8WJ+gsu87PCOtjw
ZYAn6BJ7TNZ5wIHlxR7HnkNU2KZ0l2pp8jr7pttJJ9Yd/IIa1KrSWXCjwFjwCx/7
qJ4dPkPzpBViEhs3NPH0N0+5FDq1t6QSvySYdD6bI97iLLRBH/2hvFaKSiC1Y4pr
iizd2HBBTI2P0MDee97XR5SHWLMAx+6U5eWY7sXSRfg+1kO6pjZw1mHUby72IeNV
ZHgvVTTWZ9DSc/GoS9Jc5/tz6xNKZxHccgO8ByM9AVXfHbxGephDlaUv10SNDm09
2ull5/2BbGxQUXBzzyLlRfdo8zOmGHz1FIpNaeTADf497i9lt43H2Ij749dBZxvZ
F/lgj1aDJyRICEIAwO3TTWG1UepLrGYIf5u8f9ER1E6A6itLAVJ2HjpmogYlRSxY
A43pyhRj5fqqkbf0uABHoMVhbX8PsWdnMFV3zfG3C+k32PiBTIXtuTpIaAVffZHS
+yKBiycRdBT/mHEFE3OtnHi5BoihHIgi6FJfU1/trYZoBS3O4+LfoJLEcwcT+MSf
SuSan+VoNjN4ZvJzc0qbxWYMTKCAqIxAjfnPuJesCXluMqKbHiTvbo0MsNET7kLU
yalsQiv+oaBXRvwW0NTs0RbriWGfvVRlpBzJ9tXkfvbCODR1a/G5bW01wECvTSj8
jut0l4oVg3LFLC90ABE/Bm4BHArysWaNSibXAi6VWnJka7QjOfbrS04vRFm1XWRP
fivHCyzOK6ANhrbnyRVpuYFmpzV0/ejoWsnjxVN5L2uydUiwvTazCTUs9bbgB3T1
kMurHM4tniYqsCN+qThoVFIib2awqVb7knP1mO3pqWZ7OfoLsjpOeuXaxs9PZ4Ef
ny42N7rhXDKneaQDAfAjHIujsB0qB8z21ds1K4VctJ3xcvSVSahZtRG/rSWSr0Mi
ibyKIh0MzWTZJJtUdHe1xsj4N+UK1MaI+flKi1LjMXR/QgdLhUrc6I39AJwBP2YV
0fNL9f7zwR5BhDshE3HZ2kn3x5ufHGv6g5h77pPgvJ2emDC/uPFDr6fR0nzENfpW
Pc4H9k9Yi/e1ftfuHeZeDEXqa+3oux1P3UaEFQfMpi8rpBDzczBT8JY1pd8vylzd
zI0LgBSy9+8O17y2p3pxZcE9yxywP74Nbdz9+CmXLDMeIxpKxhbg04HvUYRO0nK5
Fowi5efNNlWV6HMQ4JeFYtdIxIr5SwJs8IF2BdKyqPi1AbkypL3IKAJuq6tYzBHN
qFchytl9xiSVD3yg3zbjbNk/BpSAkQVxv9doBz52GxBwnh4pQgn7TLMAwrPPUiGe
dN2AQ1oH8H3UkCbO3IJsmxPHqO4/08JBlrNZIDcLH05XCnt32HJNeWFTnREMO5u1
U/kV11eJabFUPSeEoH141wPOT9q595U6v6YeQeweivp/G5C52cHSceJ+3aICePqs
NEOm8NgM/cxLC87Y1Pd4HEXByMGCzXhMEH0UajNs+/+vS/mcY4CKJVDD3TbRV1sE
u9KKwkf12Apf4YayAioMoqv3+GUrc+Nj483jONYATOTgiOvW/BRV1vl2ts0OERi+
9fp9c65MeV1FwATMqY6TTccYsSDR+3ya00dommN4MCXM1JD6h+Pvhl+6sPO2yoTK
NNe7Q4/XbmWwBHhVgYOeCjAqcBR79iaXj0Jqwkxu6rNwu24Fnn6sIpxuXRmTqr7+
4FaPoZ4HEhrLB6pMWPMiDEaaPCiYD+RasrR8OGXAVbUI0sAKvqxhmHTBFoBNwykq
X16ppNlgp+vXZbJYf2qKn/WGarNQvW5WBg1CSX80BxHY7yhjp49kVUZ928yb2JVE
cUi6rbKUJHVsPKlkVP3fjE85u3DGCeilrBq/+LvAJs+5eSATz2DsSskjurojSoOO
cEpH6gfzC8u3+mhuRhy/GfC/SrtHxVxCVjJ21Ry2RQNBCm3+PRRKrIgWFIZMYkSy
Ws7sF5kG23u/xhIvdIyfROxPsSvr4gw9PyNJtre0LbIKHb2fZtjqmK854r7vMJ5L
6KHwcJQiykI2duxPWyrkSeBHKi7ONMJ3XJ6P3CP/eTIrs7ECn5WXLMs6yWw1SZmm
exR889oHh0F7H+23Reh5pwyS+NYZORFzCfRH17fZl0RZA06A9WMkO6i5uPBeKQ8o
U14z6kQ+v8fUZFVnnO2u09Ih/TrKMH/INt8c2E5GwzoFJxmLaKcZA+Bx+kEeTcYM
dQQmVhvuIwI7LciNh+/RbiC+z5zZbP2YivQu8+bEGQbX3o5d50Ro6LAFn5K3YyvJ
sZMSlVU0UsUgoCZjl70fxIr+eaDt+Ob3VjkypueABOjkcljpaMqOjXXHVF1tsJCp
LoxBxflvpQbf39B9SG8/+uBa9kv6r0yg6cYgRQDE1gm8RGuDmO2k/wmVD3pw+y8g
8ELMamsacnragkoBi2wQzwkVKMGe2pen9byitZBriIRcERc8RnW01+8JfehH15Px
uePl6+kC9wufkQm4LEXFQh2qyn+azDGTDKPHd2OCP3h4Q546l/4Jhp6rc0FUt2W5
sKNMonSzLEPNSfwL4YamoYRFHHYXcKRQxemd4zGuuMCGYtEy8d+qgsNnfiKrecTU
4azoHJFkD9e8P6SMQjkZPlBSfR/NoxT5NZ5y8q28QgnrZg/yUaSrHI88658aKEE8
kS/c0tCaCdc6d/yO6GCOlYUfR2hVb7IF6xelXx9R/Kvm+0q6YgPganr1785IVmvs
/yMmKE8HDqM1cUiOHDLRyAG3kaPl3VsXyow1w82JQWFvfy8zxb++GZNSGgvHKpGB
ArvREJA7zqTIWOJ7+JIrFIKE5gHFU87gBGUuiRP1JgaL8ygGvhEHOaz+K1dfMi5w
ZjPiH3uCylxdFMi3H0/rXWKGBxur0y8Z5JVAEDKRry34VFiAE5nrNndwhJDKLSjx
qiT4ZOQNOUvTHmbRYF53Fc62zI0EyAEOD6EpkneTCD3aGw2HIHI9+hI5Wol3fyEp
Bb/2opDkylYVEQfeGv6jvLXTuayYtUO/ziYKvx7Co4VjExhOKp9yJtJyVqbjP1ux
TzgGdp/eRLqMz/yiSMknVM9v2/9mlmne4JVx9DiYC/ptPAQMHl/DmcK3KwjWrr8Q
EVqJwIlLiFm/bxXnzn/FtxFuWpHmyfO63/gXAgzP5otbMbhorLMHoV4QX0GRUkRX
q87mGXV+RV7JRhDshfFx2obPFAHbaMIp9kjNLZaOSLd9HcFaTvO/SdWFPSjJY2fu
hA4wWuqacmiR/FrBzczhD4MEENa8HIWFkz3WiaRs4vrfVnt9qKDtufKQISSAyBrf
ZuEjbIj52MNSXKfD0oZulUeYYZby6NpavoQ9FiXeuQ0yE2+7pyu7BWMailzDAbeg
G98VFTGyrMXGWWixUT7M+kmMlBURqWm+AbEuj4viDTjkNqsjol2K4ZEL8Y908vpD
byzf+C9qxd178bN5dtlDUgUrGJbAn2aGEsl7n0HIlVCf3FaIEmJEAIYHTvaYbzNM
PvP0zBwIInk+s0aa+7GpmmY4iRrKxSwQ+VyaUCYjHbuyNjAmqnJF3qvxsW1/77HV
08OfFw57EOcW3rvrhNhf0MPrtqTCpJVxhqJJkeQldiXf1n76RV/fbho1eFMNIIow
eJBlUIkL9tV3GB4NAMFas6NugAmydiTjDICQh5QuCd9HaUoRaPS2jymo1Y3xzrNT
KEJZexLTQg0I1CNsU1JW29bBhPTa1ytwDBuMHVJ6Vp6atYpBalBVdYSxDYvzXCQM
1utFT/FC5t1v0PdGRdBYbrk75s/oOuZRb3CtPP2eviCsNF3or2PaEDct7iTUuvaW
sg9Qdv8usIowF1hX1YGZeejNMFx1b6vbo1SD5pRpzTYqILk8OEV8tqO+D2ieXdZY
Q4eQ7xHX2Z1N+yw/4CYaAMoohfFA22bPQxVl3JWIhlBozr1zT3Tl98kXhm0MU/8d
ppCzqdrGUNwv/9LApdIcROAmKHz5HNVIEzbCMsHaLYpo8r6GhDWZlj3dSCk2SVua
JJrB/Mp3me80D/lGHDiO/fJR43hYmlvlNJyfrff1e3UBbLDscWAqjlQMzRc+P6Gp
XRer5rVaQvkTMMn1e9bBlN+b3kU4XyPX+tYzEc7mmr5Rm3c+nv/v0kqCXjt61xtP
Em4Sb6iJ9UMB9xOLKbwRs1mGbEsNMAPqqzEpa+yualxdOtk/uSP4aZmmC8ewQrnh
uv875144Qq/Acj+SEZXxJArEVb8yZlpxG8+q6lzA2hSPSdiUZ0NOjsfxhuAK2Exo
a2BLgsZZOYCzLR1l5U0ew7949xW1vgdtGekbi6iUPhRYulFAy6An5leyOEe1MeWJ
hiZTMjuATzOzFA4l5z6Zq+sxgcc9EAtemaG1B/hkl2Qpkx3LMazf8gX253GFVJk1
qIlWqag9X0jfFXbG6BR0g2XOFhS7dvLqO8fm0FOqcBWNLUM+s49NEr93WfkHTHsm
Z1Kb3CY9gX/DK1b5NTXF9lhRfQpxKFX94ZZ74pIBU3YoPbrD7j+5AceXLzYYnxZC
Tpw8DenYOd5qJXReJYVb3//vIR6GM+Cj/DFx1GXr1i5nZlD9oBvbyIjqPy8R4ecK
FoE2U2iuiMcUZhcU76Y+6iuxSEKj+mVoVvn9dvEYjXOr+XX8XDX2vghE2Z547l1r
bXDHhCWOHB+2MPElrxejJN1YWsPNbZrtrFjHn/PpthLGDMRuX55S9yQoVDKh8jfe
MBoFAcpu3b0ug0G+sZJo6DWUPpJ08JpZVOfHWu0CWs4SQKaMAR7PF4xjRYlSxiSr
riR4OWv1kXlwlWEPIl/KquWHFqJHGFIScmLcvT1JAyu0VG5CuR0kSJa6gax4E2V3
H0JJzcR4SAEVac+id0VOsfsoJtcV0l92FTGGMTnfYQFLncpHloVYMPKEMdJoJPuM
7aU640P59McaMRsyYI2dc0WRd8MUtOhzR+b96a/AZNWH59zhDpsOcnhYKez6znx3
6WaSK0eq6ZDrnNle1Wwi9aCO3G8+i1WpzILsiRUH080TO6k5vYObribiV2zT9Ibi
Ug9JTKOWrsn5AkvxtSG2kF7ialwWjjZHckyLobGNA5fLELQ47sbAJo84KK1b1wv7
m2ymlEOVvoehVuODJ5SXuoRb1FKFGmowGlI1MxtiBr5Xm9lY6J0/mxaqCeOXkf/S
QWYUa9ZH5Y1atOXL4oX+Fiee9pNLF5BznR746CU4tuK+vX6XamT8bBhNioNJKYGI
evkBvU/q+dSWgM3+3aqw8U3CB/wHKyWlsmzyT2ijq8a94gZFPD/bEfy6YNCwF3gu
fCls9OrGPFxkC3MEjIPJqFm//u+MHFwia7dVEP3GjDbvp3XojKtl323RPWhJucNl
Beh4rYdz5mlU0LkV5fUNQeOkjB7BHA5iDOojWBQ1o56P2wJ5BhewJWlww0Oo3Msc
e9HtNRvJFW24+eUxcFTI/rojHLUKS8btTSTNLB0Wf2A2JUdr2oWvHCkfs9i3KQYE
wvFSykgmGKT24/vXgCiat5WrAHHYE79vHehRaWWlflUMd1YZLxcgbFbNgyjKkEFx
J2J+AiviJJC561rBJEHwQwDu6jBR3SPexrjX5KUJ5zVE3qu5qMCK+mHCegwU6PLi
5gvLBV1mm339WhVVrJ2/11GtZxgM6cmgiUtPaR3eKdYZUZViF11SdVBHf5pQylNc
P1VhUNho+ii3o0LgytjhrKWGXYSK9z6ZVc5quxz3HtBIZUz+tY2FFlfsc3YPv3wa
wYg+7sV6vaRvU/E/OUyZ5unmu13UVSXaexM7kHa3I0zCHF+7gVUEtSezrCZNfmKe
OmPE3xEgxU0mGC5+ZL2FPaciP3meq64/JNTM81D/Okvo+bdbuPMI2HZaurF4pW6D
YSNTX6BTB8nYhp8i+p4lQMP+I4mohpJAQuV1HDawA+guUEqDqXilCRCWEq9Fgcr2
EerdKpfz/qHw8LZOwSH1u4le8MPZbbMq9baU8/AuhwAvpSm5aLyiVh0+BccChKhC
X316YbrXoPp+zXd0nojAKvPpVMwr2/1JrbNDKIn6RnB8zjjZLL+aJTscDfqz6iAV
0pQkebezE2SJnFR0qHJcu0lYo38X/OAff401nnbN3BKzB8PU6bu0jmbLPFVkoR6j
YIGTFmUYP+FvUJz8O4wGoOjLkyRnxR2xMxR7vrNtqug8BYzP+MINe7chMbWST2fP
KfZInk+8hKS5z5QqeETMYoW0VVKyXogO7q6cRLsjpVwOwLdVUEH6x54EyPULdozM
mmKx40Xq+CrZIxI+A6QaqbMSMg+/voleTid7XkX2chUOVttlg7D/D9erXfWDUOQW
VnJRIZaAJaUwWTEbepHPCKUujVs6KMHlJZJeBZO0M/r40axpq1PexnJg45b8TA8+
2GTwpiTlO0cMuLuYE4VQh8iZsm0somoWmIKVHn32eYVdacoXQAbukcLe5KeG0Esc
cHzV4c8S1xkR/2u7DnR+9MbjeMfbG5vVyvL1YkWrYJNZA4H0e0RMbxvo+PQzl3J1
3OIptq7YKKJI0WsI5jv544wBrTKNRIICr97l7aFtC7p1wY/vtPenG0iyNZ5gCZF5
ik1OxBPA6X1xiFklCsujwIbIo0iGf7dPSOfKzonAkyPs6fn6N6wFcdbmPmDKgT8A
I1GKxWIO+J33fPx6I3le5JrG99AbvYku7SRlZIYBwFdcHZcJ+ZFcC7Mw8BFDiVjw
jHodE/x5Kf9WPEdmjlAk+ghrNsJmEqQP+tL2PYrQMATY1fE4vtcN9yEsK52TvmpN
UsIqgHdH4Q4YXj1GO6afE4Bl1iYWWPcTu2R3Zv9W/tOIdcCfM9s5N2GyYm8bSr5N
8rHG3YoM959+uhFP+8tAyygVLlLTj3HHUpW7jzXtfw5zYIaRPt5lTPy5ba3ALo2z
tE4jEVer0AgIMMxmCmqfKORL/W6SlH2j+6Br9I+NBH3P2XRh/amSpDn5Rte9Mec7
5ii3tZ8g9Sf7Cf2WrVVy9kkc86ccS2wyQvwShFddpi8303d5sPxxhn8y/odIo4W9
diiXWKT2QzVnsl6aAi90rFZxV3hcfursbQNmZIvaITkmjMLtlNrjslb9NiyosW1d
s5A7/P6WYxeyyv/PpoOT+aeAYmya+aUZ8llVAymPv8sq5EumMlorJXtbyor/DaXV
bSXAk7WuIul/MZvAnQgRLjrZvXero3X6GemIO/E4Wjt43Z10huvs/l5G4QmUf4b1
CuJugIh00MzaqnvcsXwZ7ZNNBe5alO5NC/7ano6v+OxTT97rAfhAZl1yiy5E3Ws3
fVWxvZBOefXAlcex2j4qka6BsvSppeOjJaGfT409aEL+Ky0uE0okdwrI3JZygKft
obIFzPIqO4EsINAOe9/HqreidABOD97+G8d3l6FaAUbePuViTrVDZ6Ew/nuzCE+q
MtrgpONctA8TC8aw9hTCrWCUO2jmKphpjtIPGkJ3IJAHtIgHzObfxrTC0VTLS9gI
gMh3WfE/JkQjjrQ7P3VfgT1WpOIAr3oPm8Wsv8KDVF8yIskoeEdd8HIn6hcSGgWG
N+0JRPvuQr0/UyX1V9+HV4DMrdOPaLnf5BG4HrgsB9DlBIDYaAe8pf/avpcWcAkk
MmX0q5ymKJHrkjAFJCKr3MOgPkPFRiLhZFazNaH0zUrlmd2vp9U6mjfW6goXVMAN
fCT2qm1/3uYg29HtGKWPwyPJ8IbTXJQlfTzuzYRWETnVN37hh3D/RAx0i9qhzKuF
8Wl3PxHpmB8DZAOJA2PxVUv9lDlBHY4SG9mQXKm7pH5Epz60WnkreGgbRTyaFbkl
HMsrBQMcJiEu/+bYY5hVbQfs9dp2xvCpqE95QGAPhBuCJ78QOHqU5dPkus9tEuAr
bzGCyJHJP09j/ZP2j5QPP/L8YPmG4CZi379kbl9brfmHQbBB3ONhpfBJ9owzrocr
GNRqve7jLQzUiAffFTE2y+N8aNo/omn6XH3X+QSl+zXSBE4UkgOWmAN9W1ZdtOsN
740MhjdFy/WfQCPLbEgv1VOE0Rk3wan76b7cRfi+4LEYGrEFnRMG3rXYxUN9WRzj
Q3f8xehyeGwzuPhc8z50hVyuUkzE6GBfFLJNSy0fZ8JSh1CbDASF+gSaPQQYr5LH
dHz7QPyapctPRxkMFmKXmc0JLDsdnU/D2zLNvGysMvYa2OkgC1VwY2OwsfH8xOuv
C/vzCHPO1qVk5l03plHcJ+xEbmabAWqRKWiSR8xZChhEm2tcz+vefJUpxdH3bFwA
0cpP0BHZsFUnLRKVBLC+TwYMKvEduMaSxLWqp9X4DZmPxiVh5lpQf9BHFhkKf4u0
l7ZN6+Bawn+S46UMdXduuCY1F8P69ruxDGh2GqA/1Uwaxaml2ipfGoZnzT9oXphS
tm+aVGH70fI9cMrLdtYuUfNkLmVD3cXnoBGikUOmCa/2trvxYyd1Benn5ESRpTKY
p9lOH1nL1Q1cKAX4y7o7ABVaQ0TUWvMfcT3ezenjDgHh/DPZto/h/nshbSQUjBC8
XVMB5d5nKrNpubnqNnJl2EJ2Zv6H9yAb6bF07Zkepl5Oh/G7OdHEHlrCSzf5cBL2
fgOMlqwgzx7wwvVwQJUcsB5wT2OcHdqmL2EFTZ0GbWbULW7L+GKyOrqGTvkj+C7I
ASijh6rsei0IJATQ/5SvTHrP4TDgjECJ/HZEAReg75DCItONUUCDjsnpP34pEzOk
GEZcfnXEAeVkmyuELlQiHa1w+ebD/MjNpDtomUaSGmNVxxcDSgOL5dDLIvAGpfVy
hPa/mFoFkmeEDHvFAkCT8NjlFsxuITT5hdIxCXRQ8xI7pYN7RyMcJ5WvjZFjOKgU
ypNDWQEtj/3u3ndVn1eKjco3QK5x6V65J3uQdptHpQv005rqdZrEUNDmG01ay6p1
XqWowBokR3k0uYPRyR6MLf30Pz/O4KoXG0s46ONNX4bjGNNGICUxQ3j3mDssDNbc
49vb/19IcKi6VK3VGBzsvWnZHQ5IEf10KWZpwkvj3z2UGslk/KmBA8xcJq0AB1ME
iH1bqDQpPO17AXO+dXQX8GmAFwWM8WrRH+muI9tOpDtf5sPn7dq1/Fwx83OB8i2Y
9HSv2RHOVUQl/NDaD1PsHlG5BmHuiRGRn4IMXux9K1wr0FfL/dKIlCuOVk03vrmd
MPfbxhWdTRcATBWQXXm7ZKaS5Dl4VkCaom7IMOf1PLZGYyMhht4uLidhxtBkbQtB
exOUVJsn1VD9TWNTOiLUo/cknGx39bGJKw4R5lmJ83X8jY3nIhBAoRFfSCfqZgX4
e46G7xERAaWprVEl1EL3J2i4LFgFTS6Si4Z1xZmsTk2nmITOIwGkjBer8HhESMaV
kPj3fJOyd+haxNC328mN187Ou0jTjAw+94Tjl2wB273NGSuqEXrLtVtZmuIWbPbb
cTzwJG1TAL0DT8isVvaJGnBogPv4aQ58U4hytNumGplIpRkBClFD/W4Owguay559
3jH9vdDecqD435gQr18Y1Hl7jowu/eoBXd60YWRAsCOCER+Tt15u7UQ+drcT2KMD
HLa3GNcMxmxlL/IgPWNaIRXagjC6SX+0Qw1GYF4DEmPLUWtpIIPonINGLSoqt7fA
2zpPxWLfMnIrxFGjJ1waRWTDImGIfvGB5yxvSbUigsamgQoMFgY4jnGZTBR0mCV0
NoLtCWCN2Cpcw649CJNDZ2In/DIEZTXwfR601G0X9fyXnaA8OpZY3uBz9tWVNBsA
1OOgCf/A9HLp5JNTQnF8g/4wnUXKd3nPmyRG/Woobug57o3n4cwszn5tRJ44tQru
8zlwSYzRVnyewg1/TyQ3Uo1XdxWiZU3k/2DbFlP/sorYK3rTf1/Pidj/6wqbbP+s
zWlnu5Gr/JWBLhAfGMCcLhwc9yMt9ueJd+RfOCh4geFcweBUca044txt6F0LUdCh
0jIVLjZk12s57hY62KHRdRQ5kSgpDYIopGdFJ0Dek/x68bZ2WZ35OP8fsz7u2Sa5
aitzc0arQ/pJ2nqAR5IZveisCZdQ3OkwraEkdyA/eBKCbYE+4BjYEq6C/fxrRmhs
dLOtbFhaEs1koloDDHAiML8wC/ukOMqBeAn/Cpmw83uAYeDLSkBYMSjs5QgYP57D
QovYzVvEjdxt/3/xDSF4qM1BDtiWTw3FNFZYGKeEmY80DtTf0sfwWZrl4N+yxnQL
L2O0I89IjHVyadphRTv7rebfY8Ng4WmgTCmWGYDxqey8PDfsdtVBqtkeMGRqu6P9
vg0JXYyhAGBQqbSw66tGQMgkLMV5aVw+x9S1rHmVZaRV7Zuu7CojQD0i1xlKtTVm
vYrjjSxguZUWHqq6KahkNQ3uEuU2t/HwWcxHO+hfMsQDsOqOO3rlNWYLQolNPysn
9GDuiu8U7B9jaEzdcpi7q1H0Z39C7k/8MV8zfnc9CI556BS5U667jN4zz8w1GEx2
KmcysZKfkYdymqXg8HbzMJt3hPkrjAk9yyneG5xwINfFi+c7XKo02j6b3jyKdLXD
aJkfDEucVcvmOX/4zqRJptSereLbOr84k9sbxF40dR053uGFikcgo0xXJ9mIOjAq
8lAFdlfIJGKWGkvCYI0f6yinCN14OGNq5iSqC2buY9jDeTgfMCSeMhzfSFGFwLFx
LsP94pxlxpshgvVxTqBCFnNi9Qu3G2aVbXH64EjDcGcDNp5PDXv9l0NaKIodqera
VCXh+uph1jqRxFccwaHees7s1kK9YEeOJK/byR1C4JZCHKI3crkvAbZsoNJw3HVs
MvZzmBEY695hqR4n90QY51FGj9Rn8/M+K/rCSbT0c8R8wLOida5EVKvLuD/URglx
n3wp/dU/HdIpmgEW1h0ITL4t75KOq3krRP9TXkU/Tgz6iblxvvp4N9QKF1YOppPa
ESiXgDri+dgbZ1wNjpZpLs85mrUFJVpTIUH9D9RyPkIR3jnWeKHm4TLXDgvQr6LY
oIhfRvuMsK981xWKqt2ZDV9pbhV9fmFQJ5WNBljL9PqO9Dt4CaRuT4TXgamdMZOG
0+KXKOnbinetF3Bf6NqBfkWIES9DuXmjRq/cVg+/YgE0Zz3KDpbujhDJuZ2c/frT
5zYvOjuIn0ECT09PrSs4j4wUPCiA1/M1xCnSharQQrG44gtINF13lKOI23IxdJmw
rYGyWZoukfGXhbHSs5ozPgLrRo1ZrIs2rLLwDvHnQBs3HfcaKQTytD8aGYe6bBDu
S5PF13cSdNITog2ocnAsN2TSc4FdcNwH6LnKkLDcvYGSvUyf7a45MvJ++oUhUPZx
7sC9vP7ScHBdXC1n5Bvg1/LDBmq461cNxaCit2152ZWdCSjf9AS2lRZktuO1LyF8
h2wSOJpDZ/OyS4vjv7JHuIDQgrKIKdfHb6dNkSUQgD9GzgVD3HSszVuWrMgwyXh0
JtrqZas5TSH/JZX4lICZ+8jXVeaH/0xWnUa0oMUtb/RLr4bZP+7h7bEWx/waGmot
53OPBxKKo78KAc86FIwp/0RztqCZynw4ApBKXK5FIxCy0a0HslZmpp+NaXwrPC7c
gZLt/zEjJOJ4MAepCM6ULr2aGAHeg3YmCn7FaeZf1E4fRx+Tt0NKq6c4T6IX4syL
H/CfZ9GBEeV8HWrerH4sxKDTjfodNdgBnvDuB8DUvBhZoDBUWrfxQ8k+fN3z7KdJ
s9XxhaTVjYvygbciyYieTrzsVTpC9DCcBzJKr3DsR481qws+1a/YvPMrRE8xRHYU
LCWUqeZwL3MGI7NNv0pGYEG76gTzUVOHNL9BNKdy8Xjn4tpmBsdoI9l4p73eNE7J
bRwF3QmUiLFar/WpmANmOBgxiV7g4e9TDXAJNtCzEZGuYzXXK3taYwReHV/G0BRM
f0cDrV7qUaQjP9upzc5F+Xi6n32IFwwvBdXLRqL2jw9kf14RP+QDl1o0YKe8YIZr
2P4rmXAdGAj4uXCnaUh1WxpDWuyY1VeC7BLUtmDZaVNy56ZyPvemtcEgstLNEODQ
SxpKiXv9UI1MaYRrmxZ1sN9Z5lzpWzG7ubtZK/7Zn99YCC9E3FSpmvJM+IrrVDJy
Z5ogz7D/0jqLnEULEDKD3EFjRFD7V3X+4WXh8/j0oRUkAixDpffJ03mw9n1HgreS
9Qvx5WLfOBuzrMir2y3YupKIt0oplX5JUMmYztPslQ8q25Y8dXMpD7DVLAv/HKj9
VAX7+Zt+AEuaqPdt0j5M8iZ4RwlwsAx8BMVQ6jGF8r3o3HUN4vKmisb/TYnRZhlm
duudjVLwq9SlH60UVvmI7bwb27oaIyUxX+2HxO/RB43bPLZR1q+c4OgVEgMf+trc
rFuxXqQxHvcdG3BkLwzjaooK+qYEH/jRGJ0v9Qyxjqbdn1XgGIgZ4QQLjNRjs3I6
Yi7nuo+ZcSUKPKlMWoV3P1Anwzjc2HhkzZM+pb54U3Rl2QgulraKJnwylb0B4E9o
Bb1CftHzG1mSqlElRh0zO21/UKCyaOF4duCAKxmpkd+fceomuKkKzwG5fxzdg/4o
fmxk+uNbBG4lfW5V4OJCrYeD3Zf0aGLgm3nDwdXvCaYagpJtUjNAydCH8Jdz3I6q
BXOayzQeg23MAsflXPw9Bz/BC0AGOG/iboNdrFKD1kJjdqf2cwOJXv+dWdEDLX83
4+lGVTu9L33QLppHOfvjaVDHA4l75Y24xg9E3hYgOp4ZSm94fYSJ2FnBOSR5uWDd
MOVbyRlE9Q7Wyga8j/5mctByftAq2AVXkJK7SxQrseKYz4LbLpdwOMZHpIiWbHYo
I5ZI3j5SOZLFR6BcjqdKwL9SYSNzPmX68/GhbAdIIsvS9OqpHBsVFDzfkrxPykyu
oER713IXcAtkPhoY78hmebtkrZHYtnuAOJiHkPPKZKrmLd1WSNZYuZVm0jQz8aDS
h7yUHAl2jFx+L7sBaioxLzbMRqpEMhzE4e4+2iMPcPcjgpzWDKPJx1qp85a3x1gO
i1OoZzVcPn46/TJr9gThsPplDnz0UlzKPCPFSBqW8xfvWz0jWH0T9DFha/GXqnoB
1qa7CKOmQ4h1nuVRKonsmrI5ZRpd3P3EKsxryNptT4Qgpa6MKAk7OD5qPkwUEpc6
YKm5P/cvWaUnML9H+QV8iun5AkJfbIZD8kg1ALbP+ZwXnj311oZvmbc6pOI3YinG
rGGDdrwl5MK41PO76QzQLBp0UnGwSB5/1ES1e25m65uodg5z1OhCgew7GlKxdTV5
Egb5vG6N5iCZ4LPPW231Nk1As9JMBcGVjh8u3E+Xuwo/ZJMzyUGOzU3g5OaxKJmy
H8uGCM06EVDN3zL8RCdHL5vg+IaXdU4sIc7JB79aEQjewQMNvXABsh5aCQe1bxPt
bstryDgA+aOuZEia/E4qDQzXn+ArVrsYtVkFbGTCmUMNVaGF6/9YE67iunk4Yu3s
5ULUcFZUv9Nh5eUSqGkm8hefCFugAsv9er++WTRtUmSywprREqOmAe7pxnF9rxXf
RnsK9OTYKHM11gwaPcflaWw8aLFj7KVSiYQBooc/D0NufnB5i8Pyn4eweLbbSZI8
1e3jrajasCI9dqABmNr1BVn1Ub4uCrVAjf12wlD9xrpnPYbt4TkyDpPlyzaILIh3
c5Fhb2hsSAY/IucQKFVu5ldMODhPXBpUo/c7FDSkKWRxQMJ0tHycXG7bPIuXnkUI
qVi6eng/akhpfg8aQbof+GBbU1ttG+MfhE3HfcZ6DRiTsX1uXcJBr1Tq7eYmSKUc
yukJxC7FUWKUaERR0VMsKm8JsF5Plm9GaP+SgWQFcIJ6M/koVAYrZqFpDJ80w0BN
zsbMIkYs2iyIu4a6F/aaIsFqI9n2n28Bjld4GDkGBM8raw+ueFKBM1sB72MgYifp
Rou0GL+FhAR1Xor7USUB8lZ+u3KGH1MVXoPF6wQBp27JTq6FlzfTOTrjD5hX7a4A
r5/syfefFacOofKwYOJzxGaIKF3cZXcIojHcFzaUloHZo3gagyT+qTrZWXAyvexA
afB4rVpWE9rllIXbHZ+F3aMSURZ3LEJvAHuPocDq1F2vo12sUQYrOfQ4A8jSWHQY
y00yVqaKq5ZU9H76NJdQc9Q/CL6c/C+icyNSEgAWYWWi3q4tsKxK6MXUvAlR2eL8
/h0V+jtKfyFIjIaV/RkIYKnnfu7BuakB4ygToreLfDzlJuiyaKOiuUZNS/8le0ps
5cKuWNwmXIBaOMWhzygnx62GS/blh0BmtmNH4JEapnNPUPz1WONjYdWw86VlxeMF
oAv7DarQHw/PyXDtmzoblx/qy+pZa0YGJMqO7x/9g3c5TrX3k+SUXfiN31VH8r1I
F8z6iryrjdn4pDJ5RyMghh9m3Y/frEQxC/sWzulq/HOFk2kH+sYpF5sDB4XbcGPo
PG4ry3If/VJnTN7OL2Tss1re8OH6NpX6iD+kUpwLdkmawsBbUn0N8Lfa/j7VTq8Y
jHWISSDDVm1XN+o/36Q2QO1gGuS1dYq/yZ0u+NMsE57Zuht+AZ1+jgMn5RTu5Hh7
IjXBhNH03Bdm76n/jG6wK0mor9o+qFIanYIiQafEUx2w6G7GhD16F7XJWRtfrcsW
Fl9Vycz2zNcfo/w5jsgpWDHpgHnVV/XsTwPMfFHS5olF83E4l1HXQBxZwMR6/NCD
V4qMcXYT5OR2Ds87LlLL2ifiru3t+UrY215XB0jItZ/HEp1tB9ao7gY5hhUDB1Z0
rrqsp/zDDBbytcwlOWXVdkswMTZ4rwI4LE/B+kf6VYdYi2Uxa1lZI2kknn6KsB+0
EsMvNY0xvCh5k16S6VBBBgPrA4WtLpitFkrfnkofrRIrXTwxYN8afZNxsgnTPdxx
UIbsz3Tu878XzqkwuRlU/pg3ZJSr501T1VYARwar+fVQ/PEUrVr5RH+eVGM6CsYj
Z/KY2O3RN0BGVy10eAOrK6Y/a5RssjgWGdi5UXAYKqtY1vL9iI2pbO9x5cMXPWKu
Nh4E0TkojWgKXAIZ65CSfti3AhQxPl0NnbiQoVE7TTsqtsJmkK/AAlr/NVHuoe4D
z5/3dmv4uHBM1A8O2gC2QdO6EsJNIdS9BGpbWh3Zd7XIl9G+c+MWkv5FBIHGLwnI
aJ7obGxPh8/+bFAZTcTC3+IERLNb5DZsMQ21tg13ftBRpk1GFZZtPTinCuF6fTEY
xqVu31Z2q8bRnHjZg+P4VhHsHvTfz5pjhqBHTGwfYBhfp1c4duIAEW1enMmjoxpN
21PWo9pBgeTpaxFjkFXha89n39hruI/PaLlzhFe9XbvLKeT5JP3oquhVl/M4OGuL
yV/FDr3FBhbDN30cxpOwlBgpRzJS4ddFwm+L9neWJDAlmpxcdMy0LHeIIIWAL1iH
TGKmM290niZJJ7IiT4rOrmOKUjYBlguhw8XqK19j9QTVVO9xNAA3wbp0C2fCrtOa
xTPrul2lFg2DbQD933ZbLV+LHM8MnlPKRRkXIRkPEzFS6AS5+dn8RQGHmBIa7ed0
iKOieDExJFspRdf3+MqOs1P+1SszauKWfbDHplGsjNz0csFqkBCzq06WwaBSGXqK
xh3PgR0bln35fK1p7T+93im4RJlYIZWPsfRyB627C+dxetLzi4ig99ZSkGffcQ6o
wMjDcmRndTc7lJtqNjF58LL6nOpE0COpW7xUQr96YipSmcBDLMmA77BKMMl1Ef4C
5ePQN/t6c6Fw4GOsY0bbPaRbLvc/WIroFk+V54/rChKYXczzatsiAFVTmRzE5Hpv
rc0EqBMh597nXELrDUcZLX8+NVwHuvAQrWeVDc49t7E1JBjgKwB6qHaJfAX1xKvH
/BJW5ScnRmEhlE9VdLtY111wqpCHdr29w8l03EMHtvA8RlDNqx6cnMslIM/ftCS5
P/l54xaeIBKnHwSu1xqvDW04blJrGKLjz13v+QdfvDjhqGdoE1B+4ffOapNg77d7
v3rrpdLHAu2lnNreSoryrsXGnyrqe3AIOZbie30muKhsSNxmz9sDNSIi5I7CwhVi
eAZFMUzVE7u45oW+P3wYaQy/NPqOZXq/yL8WmI4oBnXe8pZi9iK5nTpoyqVQ9nrl
UBZ7ynn6mltAdCgDpueARX3anu6zk4afJQkD0GWWEXOMQhx3pMUpvj8rELYZJ/Xy
yCdSwpbulrw5ozdXh9NyqMfuPCL65m7fJITtfN2F/V5wvdNCJn/ljFb01vao0cg1
HDWy3V7vv/cVocPtVrOKAMpOs2MgKy0Wlh5ynrUODJEeDYuWzbcKfnous3FadD/6
Q5avUa0+ll16Cy2E9CR7/Nbfab4caJg+f+koVntYEdjFiKFPgzj0iHCAIkRlLw43
5FO0cq8ITnlJNQ4BxvDJd3ooeO15F9A23cpYz79zx0erfFziCrkmValS30jNm4Ba
yP/QV1q03hrzzZsxehGhv9xDAB2COyEu/w23jkinXcZlNSy1oOt9/y3p0x9NzR/b
6CwKjQYlAmk54nFi5DT4fArvq0FEgzsRWYTP5Z0MP2DwrdbP4VwsHqhftn7Fua6e
/o0ezDcqNNff4fLXVNdLe02/3h7kWKc2OIW3bHnUzS5+yu+U07uMg8rQYf1Xd8l0
fY8B5pMZ3vzPZbMMO1A9Ew9xQmREKDWGpIry2NdrvWrhTf970ZLPyEUnIq8FI8mu
fS/qmJawhjQV1Jkq/lfxkn8D/Sb3SgkLoAIgLuXU1R4Y4M6mhMmpTwCtQNdJ0HMy
/DCfJXhjJ4iT5oQOF+390G1ntrs/AXPmhYYiNUer8Nttv+ieDAD8phgvA5SNzSEu
hOo08Qr1UjOJp30VDMiRrHQSH263bQdAvog/tRsdpoMGav1M5ZT9ULtuwGkhVTp3
6SD11qbdZQXRJY6YX7hS73Og4KLotLSgbjazpuOIkLQpwJ3dNeCYlC8Kddi7RYhe
Ln0Myhdf3u4LH+R676mqK5O5XPzXaQmFfN/pIIbR65WfgcIC5hhuJZQR/aYdplyy
8a2wQ/PMx2+6XxuPsah2alJqEaWWqcqCMCv6AsnTLrRB1mmfX80lbmzyT2EH4qPN
92XzNKmyg2vwMpyr43qI36vd+GleoAsmcnVvh35GGuj7F95b/hCywLx4HkOTZqDW
adRhr7a6MPTUBneJ2e7OtuL4cvIS2knlHzICa2ybSpso3+9bn4b/RYUFLhCqYVFE
9h9grY0zBUW/Ayqn2lIv4MFdHzbmNDZ68rfZDEyWA6oUyqUVZTr3QK8R9jPv+FBk
0wcH09QR+4JwZu5INSkzk9r8dEDu6iM6dqbVN6Eu08psf5LcUsjKYWnH+mcX+sff
0LgkDwOL1KwT3Jg90gRznk1CJ9vHKRLslGSeWq89/sPKTQPYwvtNVSBBN2As1fuq
bYFt2oO/KbFvOFB4lpUDsfk2S3zmd9f/k43jjjjYnNhF3sp+a/jToJJ9FeJvyM7A
b0QtzLCf4ZOd4gdIjDnOEhNWvqehQybj98Bb+NZGvIzF4yEVvR3zAEJFgf/70jVV
srDV6yFKrRn6l2wlXTMdPw6HHboHy4V2PBgV5rQjdQZB8l/oWyfsqfmonKtGQA/N
3bK+E3hJxBOs0if9RpxUk42GegH4N+dWyEhcDHfIKrnv/LRgN1nUfz4NlJZcpti9
Vs0B+0sq5abP2Ke2lHKXxtp1EfKx/wb/NfFSyrcAFnpyH7vCACHKdoGMZRA7XQlN
bwC9Sn7ENw8JI0zVmM2IzpYW7UOG/6uO30UcB38RV/Mv5xX21L2HMBQy7ELGZgzx
+EhjjRLyCi1n7/V4pD2Ykb7r4bWQiPt5lQ01HK2X6qrR4svAnX4fX6JWuD/9ui7b
EO0FJkMtvfG2PDQsqrJTzw9G0P6RRnnSzCSVTiraK6gwANwzKpgT6pMzUh8X1Siy
dGeB66Lwa2+PMN5O20xXL+zOgE92rGy+ARieeQdEVJU6/TdLyuymUBOZP1Bh1L/w
Ce3vO38sTlUuEWk/ax20ZdvhLi28eT78xAXUMY6XbnD4q/bCw5FZ/Yc44dmGjcBA
n/g8PQVoEH7CHpspwckDyae+8HDXLQtU46wKg+ATzB2OobYqJL5hhPqEG5jF/I7v
7C0+LHoY0XWNJ5AjxLZU9o4dE0I22kRiQ+rKeSID8A8NUgI531ngHJF1JpvaKf3H
T/zQREinISVlsiIEIMR29+2xeVAKR2JpHX/cpwRCBdVModRINTZ3QKlz6MhAwr0v
SZibVp/2H7Z4esPJvhBEwI3ke/9Rju7r7nsRKUiLEu5G/dcJuGxs5JGvnKYBtR1G
PJvNGWqA/H6Dbc80lrjn7x2IaiDeAJ3YGYe0zRJ9c+Riyc76pJJjtyu+OTjVMr9j
FKfspcNsR7bKbD+DFbs+hTVkxfzbjPErfUCQYTqcTBkdJgkqjoc9mLZD31jFstDc
NHLbkPv97V6Y0w69prNLdFby5QW1n7yrY7cU6DzTCKVhD6Q3+jCZ+3LKxFD+nYCW
ZIRVKYNLYNIO3wgUjdNxspei/oO1x5LIJ+H0YMeypH6adRRA+2Pi9O2tHoq1frGd
t6lrWLqBkmHeHp3YLFPFkT/2C19R0QGLINqK6bQpne8WFOqevZ4ZdoKnvGwFUI0q
yWE3VMJqIkirZ3fLhPR+gJyHHalDSFeCzcL6YUTTax7bL+V2UXf5xFE3vUJ23rYC
kI3C5mjWOFooZJc3GWB2699deF2m2hffKwdtEzrWDW+4xVOdtk5yu4KAKj+mrZuE
HWvHaf2h4+W4QEaWskwp68at/e8AuEwcmp2S0KwzLBHCItRL7IjiuE5+N4aZEj4Y
8XNB7X8pIt40u+VIhnq3rb/EccIzSANxgO7LxoG8eBM1zC2xLJ3n8OPHttfFt0TM
eNTwKJ8UbjpNgQNqRsuzlcs0nT/az1ZrdU1q8QAP2SjgCZkr4P6HymiHtEETDsXy
hBb7x+kMgMCm/i7Dr6F0Z0HlISutBA7StYC/WIu23B/fJgja9WHdjTdzYgVG5TIN
AkvZDBAb0/pfwMS8iuT0PRllHULdn+i5/CMJ0J39Z/FWlZYYqxmtFCOR6ehU2VGK
5n1NYiBpX9jPEHjDnPZQrwo60mpzka3vP01xrMWTD6E1dkR0tBH2LLxWcYAQwNp4
0oKFSg6JxskiQMK56yzBzc9eN5xzN8riQs3d6oy7OaW/DUc9cswPQVX8PaTji0WJ
NdwhCBeO9h2e90zYxo1ETI1CHu5mWIiA0e/9Iv7YHw8+DjN94azlAP0UWW2eeRqL
W8X2oSiyZ86s9Pz59FYzFxZjKDzNFAYIweUCYP+kzruFDD3tujAuaEPu+YtFZwU2
euxFpdJ9/NbqP18ownaTrEblTgy3zAyJK2vahCTfNWyOSFLUiw7hymXsDfysoRZX
jqyBvqzomcvPx+JrMTyWCE/hpB6zL2RQ+RhUWWOvL6/5dLpdfL2YmSU0jjH8nl9T
+l+o8ppB4P2SpeqrP6FY5Dnl06AKPLPhjtZ3fSMlMEcT/SLF4P/210dOGaPcF+co
T5d+OAVRreI/KIAKdgrSCJ3Fz1Ezf+IrvAaekJZoAVPzrLONWXpg2oPfyK2XuAtu
Y/RW2BPWPHifdndoc4evzFu+8nvCl3L1uuK/L6naEEZoVbPbvyLzzaINMNgDV57m
ttfmvHKfT6P9A8zyWXVyC+yCPTMksIu3KYHz5QHR25pUjDULHV7glJA2jVgfU6f9
UGvP3LqnIurZ1NhB0+0qHEQM8/Fo4bqxVX9lOyINLtpTe/SiuEzyCbvD43DrtV4C
ClCkIkkYQH6wYpYwRw2uFDNcoAYjbZwoPLZQBQo2agdMuJcq+ZKRdEeo7TG/bODY
hgjJEMX/Iaw5Th7tdnsAVRj4T+rupt3kM7ZtT0lzpz5XcCaZE/+7y6E0eI5yYuyk
417OVfScOq2pwqfCAG4Lb7i5S6JyU3J+cFVKl8AtPWsZrSjPiFDzS4LEoj7UuB9U
YJcR/ulWzTMtdB+aCB2WebKxTafwbQLP9rlqYKJIjzbAAB4qjkbmRo4IhCpBsRuj
J9/sqLfEaC1yBwQzIMC/VByNIalw5IxUzx4RvkFIWMubopyORYSxbbxclw1RFp9o
h3AE02sS3zaXo710ETBRiebrDEqbPrx1yvWISr/ault1glR8QuzskuCB10yQvdp+
z+kCuizIyL7IP5WmmpI3iwzHLgyeSJ1v6dPOOtbA8Srb1/DsO7IenKZJOfWsZTmX
y+0NK+rZnrn7vtXsiK429nzlabMZVH14ai1Saqcz8A70ImOAryXNJ9D/ndgV1T8R
LveEWaQqaqO06RWVD2hKS5tjuNWY5iI0J1vORLVySIivFJxBrsc5Noq5zlc9/4dP
k4bOXUXCnkPAVDDAzIQG/FziLkxZw6Gwxk37dHCn52moUlb0ZaFE1auqNezob6cO
y1VFGA0itgmHeZ35l4Ot/eNP/VPT5o/2lXCTWemziPv8KWvjk/4mjtt2rFj4d6R7
cBeC0NVsGC9/ZxudNH350bcNfoqtBj88bqQhrTzul+CTlR+khg6TC9W2uRIJRFQr
09Xl4jsKLkoJ5StH8g/sxW3H9FYkfbGVWXbbH6kiRTfAE97GOKDkRnnPJRmPi9EA
1MAi3+k0WMQtwVGP2Hnra0xswDsNVPct2UTzSFDVaIb85/cN/KNt2+KATaL7DjSS
P78g05uySmvZrynCI883ghqFtZ3P0S9OkeoQz58VVZIwVZdSeSBJAdrYUtmhMTWW
k/6DUCFUZb6Qr39FgPiK0KcSMW9Q7PdtYihgz2a9hZUIukCUIFDE0HNHSuobCI4S
5IIipPn9Vj2UY2+UMJAMq64b0ABGHQ9OhzHpD4ZXvSg2eShcC9fUBcz4b3tvPT1h
+zC3fMcOuv0KYk7pKrxKnjVdEMlelEZvw0B48yzy/QdblqtpyNVXh7YBbltfkX+x
rvqGxenvfYS0hCTaLUcqvSUn8/bVp12epAok3DmEdewieAbPtSUcYIPMSPati7dK
KahGqLdBP2cHY/BLZ0YmOQj+irV1gvfvVbKg3o0HJcRcGIXnXn/VW6Picz0AantY
klOMHU21vyybIHI8kdqz4HbrXwnNRxBSzGsyfycK6a3ioblWatAOq8ELR+GHmmuz
d413FT5N4Ha1su5eaklv+dohfNs84a+EOESnSJie5np6zEdXcu6F+RyeTgrvMuSH
om+lteAAD18p42zBmNPpOzLWzy13bB4+DjvVAjZKOSt3F0i+KAcR0ckBqyh5LAez
pZwqPf8TeOy5c7jbfsXDAJTzOLaubfPdOmuc+01XeO7F0qWUtUuC2KmCB+ZssCIe
/g1TzB1AnjBOFmXqhLLrzAEwHRObiLCQjrUMadAnckAsdCYo6oxVJ0OKS80S4HFR
5ectSf9x3xCS8gDkVaQbsgA6V/CEo+TZ8/QwimK71cdys0chXSaP1+N852EE14yb
DYWWUxspZq4xIMfAVWeqRSxNktGaRAwn1dx+9lBFyNLgt//nziIH1nmL/m4T8NAn
gaSorJgM+o9EGhTLTPlIIYErVqmkkdzdzarXVP/j6f7siDt2g7zgIMA0sgeMGf22
XP53AxTbGYHL7SoT9rNeTDRY2T5CvyE19ecMZ/Nb0ySg7dFK9ABJlwAkK8T4ma+s
hYPkpi8WwkcinE5JBaMHolzgdjlABmQbiVMdOrBndBzY0h+/QAfHBad6HFzxTFa3
s79+uKZ7/tSXh5LLuY4sJoRopqqGvBGSNDqoZ1sf+qdjXsqc1r7wfb2KHaqNZ/fX
h78jFf0V5Zs1fzlnF+VYNs1N4KZGALL0uJ8rKIHupzVUvNxi7vS4N+8r4wPe19f2
EA2N9y/Drotl/qQwBNSDSF9bJg7wyKe8Nf7NX5BjODHSepD+jidKbZxJadAf7UzR
NBfykA2QPPNKxHAmH0i4FueAtVr5qv5s0DgZIAdt4Z6GHEd7uryVp+d11mKmwt75
2rtJlSNLxnnrTC/p3AJXF1pDNyZI05IFv9fM4vhcK/E8q00jPYTQ7RKESZ9K+AYp
5wllUwl3skQwPp9svrhWKkYcK+BDGGAvhZeEcRllOfN5B+7DoWO3qjqb0fRF9x5S
8O04SGeuoy+Xy0FqKYsPIcGUaOFfXJChyVh180aV9Uly4HQHxsqugVvd0s/6+sfO
db2scl7C5dKL8sU6WIxiyT86QXjBdaGfiy/6QY3QO/TsumPrCv5nHLubb3hjymi6
mzj7aO5m/NhhGvBk9+hSc/wfS3oY4GAeft9wOwPrae/WpnYVCY2Z+3oa+De27VH9
AIoub0KKoFYUbgURxT2+zZ9rCbXlesJ8aDbBFeeRKjEFEZn7lhJ28JEjX9tT5sKI
dmckpVeTugzgu3a3vwI0EvSXHZk1UbM+oLyZnZ0akAURxwzNCF1XZ9qHihAQoZs5
Ma9mChyimLJBbC0bNTmzuoZ/ivOK629SxkFtMB3DU9QwZPKH/IaXgJ2cMqVfy/O1
T6iYX8oXms3T2S1e0XDdPjt7wsE7NlOnYXqGao3wFfX8Ac6KlzuF3erKpigLEX23
4ficKXJ3umQP4kQGp3Gq0f4obOKqMUMKf8eZXLBZJ3ryZRFOJJc9yMDK32hyxvi/
AJx+Jrc0S/NF5NXcxpue6036tFXNWWTFO1tzzxm2WjootWzIk38Gh//nOlztoT/F
p5kun6Kl3ETkLflqfecjs1cTJsTyoAmbxb5OVTZQtr25/VIXE7d4gAj5X+aoRigx
saFofG5i1D1lbS5+a1YXoEvMH+5jwL3BEBNqhNjfbSMkeQ+mA8tX/7HlE4veaO4W
0qiM82VOjiWMNcKww5KVKG+LN0inW1r59t5BjGPxFK54OKCBwaTNvcZInuLGvSvV
LXfT1tsDTyLJW37QHOEVt5Pw4gsRFRXXBdkwzUJJ6zyqrf/VaZzb/JDZZD+nS/8m
XxViAnKEnMpvE95LkjpLaFeIEwRy9hDNTfuRT3RYR704UESKPYPTWVgKgyPJ81dR
5Z0KgJgsDXaW4YcxN0c4u3ehMyiQ8k58YK8fBh0jwGtsB5AMoA01nZ+SmHZKb9NQ
no+q6g04+EYkaGoT4m4WvRBwstZkcX88kdvxUm/e+Jeo2oI9Xpgj7NoZAILwkJSX
nX2Bue0FP74ZNRrBqLzXvrwMQks5bQ1FpABoV0siTQ7F7/lKQWuOQKT6LYGr8S3Y
imDH+FjZC0WiqeLmPUidPFkCQKNwPmNnW9Nk/kSKGIihSfDdUwSZV11i0Ts7iLZg
tFy54bfbt/1aLV7qUh6/BPSEyQxvok4Qapy2gsrrnmZGnZSuhM/lrgpKXP+3QbmY
FahVMkH5FjU4n1zrzgBy7/62qLpIgjui3VZmHVu6QbJsrwbXAJymehK+xiAzDddi
FL/oG7IBambB83lCcDR+r+W7CGZjN8Nx22UwvHrfYrPI9BwQNQ7iEl0WYHX6dAfJ
tz/SeSHrZ5I/iD10LzK3hiG42kFeNmk/OeKXAhgZ4e2jCxPvuU3rAY044xtkIT0f
5PWJhf4Fxf36ypWsNZaBwtHQNZAXRQ1OlDxNx/RQ/AZ31IWKJOlzJPz+zRfLy7JP
gkNA43PE0bKrTjZ8l79CYdGSrmTDdd0ET3er65Qwb3cGvqCNvA0gZP0TZCv8R6Mt
NF3A6iD7lmplmYdE+tpSMAXfBjsu0I/qnzfpvZn3lsT4n2i/3uLC8Vhpu5weMgpX
Qhq1gMy/xIu0pRwiTSJeQvWDjDjQje0baIibpk69x8YzS0ZInBOS2jECQDFDX4P0
nsRqWhnDW3ciJ9PhgJdzSjGBHU+hDhmrQLDhPhxt1tUPRxGmNRZqJPSZ8tW9230m
Ht74S90ymtQxRMuhg6QbeExV+5a7spaCAKBDFRJ+zuDi0Kfh4GZhYyVFj6ujGV7X
OpIKkgOAFWU+DXrszC/IXQpXJhJoyUz6lC+rofeM9scLQOZoMjOWWMWnrhxp/X2z
8dkT79C72IU7RSTo1GeglviQ5hIVywFXsI7iMUVPsCj6/xsdQejn3kzAqfZm3bny
op+ovySUkiJvtwxGXDOh5JlEvhP9vBW+4tconKdQHjRlybqDbb2co8zvx7litwxE
B1pQ2O9Wm+W07A5IXF0tkES93plKiOo+IKMFVuWSH0G7zAHDW+y2iJWsE6kcVF4C
OZmS47BGLEgNr5XP2RBjxBPBo1X5A/jL4OKbSQzB/jkpKKQ7H6fbycYcoorl7RTz
fBjtyVYkupWZeV5DmwiAj5GEVb4VoCKzGEhPhcXlKgKZORcv0hqm9BBnNtlSU50N
bWo3PNf8VfidfHtKGdCrCKLPpvwSw0ExH0sl/m7Q6tCW7FfCTsM326cclMX1cDSg
JdcX22MJLIfybcsN3LQAkkwcfcA/Ks+2vikr2gDxCsO2Otg1cT1CG80E9zsAjxWv
htON9cEy4pJNaA47ATDtjjODyMQqaEXQzAcMnU1X9nlHkhHrGB1IQKiOjbX5Wa8C
PmOnmbMQPmjfuJ+sWtpp68/XMkvArMG8rWIq825Ov1oTenGWROUd+NQEpmsmgxwd
AZmoGrYtEWevVDdx+awX41zYj/Ec9CNYEbaF0nq9sQRPa0v8Y43g6gmMSZuWXjEh
kTzTmxq+9cz6PApprw3kW4tqgTqKBAH5fFsWL9/RjIcjbpVFgbec38Q5f7zPk47d
zmGQZczQmSXPreb7+W5LK7Nx4gsyV3XgdlFzGwsmO/Pauu2gQeCQ3JzuNswNTRPs
+yj3cgHGUHEWhZkLyjxuIJmUrbMM10eO/ClkM+CH+CpmwiA2Lmigw4WXHrskb4VS
1xBa/ihOyNIWLxoW8UMNthTEJBhcB7PfyaHF4V/4O4GuoZRUMdHEZObE05xGyXZR
WO0ch7un3k6urepU06Y6Xg3qGoBjvCWcu37w8jPrj1mboLIj8VT2iByrXSyjoIYo
p64/TH7hU0oFTcXjBJUINyWNYvyKA6zjqlD/NcZChaQdmjqTRZEc64utMCiLax+D
izCZm0nHAY8NmeNOsuc80+zEfyfqIEX8CT6c9pg2YS+V39hw/tPlkQZW7NDEXH/1
X8hBEjN+LfWJJhamHUB2QUEbUIZWTI1XDZJxiSfEJMiVS/jG4osfKhn/SpN3uysy
to9v6PFphhmDeSD3+TA5SLTTVVCnds9wMVdso5n04NqvxkCMONbR7ZrEl09lkzR4
Kxu61h9Q4KxnUL7T9NBVm5Oi6JskB0KYIhhDfBSOJd+UjsXn+gSODcwnSAz9Bx0X
nQcL+b1RC90m4m4RHox3Rb5he+XWfSaRBVZ4gt+MyndG8HPJ3KgyTxTgepbDSJnS
wo5AcIViXnjkelmvVseGlYxZMDSGLi6eu/f1bkfyLjshvPLF1MQgfTAypGLpJ2qc
P+hKs9TDUS7ZPu+9XK6Qq9RF0QRCkCNOq6Hpqi9xRQIh3D48gTWc7nkAjdhBGS+v
bq0jh4IOHv9U+IQ5D7/Ihv423JYKqYNQSaAYb/H+tXu/mpNbN35cCaNFHR8LIdJY
+3Q0aL6UsUJjj19Maat/ygQyMrrO2QycLETj+KupLkXrgY5lA4H6weMUd2OJciXf
q8RuDd/5kxxNVAFFQlNqSAFRVVQDB2QzjQiC2AL+5+mUsx0Il4QcQMkwcy7ngN0q
Ft9LAw66Jvz+4dk9iHSEUvGYAerAaNXMUkYGXiGzfpvAOmFRgLwwDIOamQ67G3Wb
cdThb+m2vSrbnh0vzUWl7uzvUlMc3tFSrAgjoQqlcCPOj+7pafT87njl/CrhLXB3
53r1/W2NEQyPbh6X+UjbFoB6+E2NCAoe2HcIs7OgGml9reN1rBDELmubc2eIwxo+
I/H1PV47nc2gy1QdjeIiOh3rJxzSF1XwNPEHPvtzUC8WWF9Ve2UEzcfZOpEDyZKr
CAamP/UjHD80QzGzqf6ERXJklzD3esotQXjJCDbWjSJlHOgBzct7MMXbcCndj5aG
1/F44aBKOKf0CJOX+ZGnJ6HxN6sJZpO8i9xKlWm2WiAiQ2yjNEe7LgS7ssTP11wG
J5knkXmVwNYxcsP2P6DIbwkCybHfbfAnMbp+Mss06nCcLHQTtX7hJ0UC8dG2+uwA
IKL4rnKqY49Chb7cfCDXiwWceIEKmLtfYa+uBACOJZAqAaIGFZfzXLEGwBNuubDe
3G1lK6Bwvfwr6VU6iRZa9I30eA7YojQ5vMMX5wcDJ0v8ZIqvHGBdOFEc1H7VM9td
7bzoMpTZRx8KYfPl31LAZVJHEeH7bijMzEKTVIWtTXIyE97+bgIXL1it2KgZI1h8
lxOxqktp55vr6vyTqg6eXGMLwJ+uWOC0PO0KWYwFrZBJIkfdO6+Lv0RLVD2aa0hr
C4mFUqU9qt5CdcGm5jkkR6be4nIfIEwBaJ0OFH9WDCdIOI4+QwtLyhXDEk0M8OBy
VmDXH9tEwNhFtxyO2OkkMEu9LibklvDMJFtOBbZOr589JtbqdX7ninZEK3v92L8r
+WhOL7osNsOhozSg3ybJSDzHtP/EPe6Eqid2p4eybOkYoYa5nsSzvVHlFoboyzFn
pzS0vb9kwpHIYGG1wjdzac/H/mGDH/X/n3QU8mcBOwOmGTO+ZHT/KwUEgNzypEVx
1z3zHF1TkD2XA8FVA8B9ridlcSSEYTHJkaaEd+hvdSWjIL/T8SW7k5VwGI0axM2C
ftAReMWl1VSXsK1tp1KYneF1IbS4+7N+EHvGtj13lvhfALtcsn2XxV2Y5Ccpvf6c
pXJJHEZHrzhG8liIMJGZ8mKRdeidqDpvdCgS1yMQ7ySAfkPdvPBlKcEo/afU1aUg
K0mn8OXQ+bHXAHM+ZLaPGFlZUYAdov8GA1HgmZ3Rw69lFAewDduvIQM4Yx1Eww8f
JkwUVon3A32LMS4MCwd6oUyB8MQtZnGFglDryVDlxWNT7laUFIJ8/zi19Pyr7/ud
6bQ6HCmYsNv/cKkyxg71dQunSOH6JMGB43VRALoxNdS5KqFmWUKFoUc1ywbUpUx6
wlVAowPmoO7MLDkqU270X7aFwMlRaVq5LE61BXHSMtawyO1+3EIUem/AaDHCq4fe
tUZ3ZMoljqXLeqt913Vd8bHkQInAFgILfCZ3lW7/5xvD/FrwuDCMHVoQdGYeNdfw
8BRZGPdNpRH31oh7KSo3gksNAPgojLox4FvZfI6YDmzb+Smhly+9PaPnVfL1y2JZ
hMNuwd6rmia9gz8PlTDZQ1XCdJPnLFYQ5Wc+mdpejrM8xybK7D87lVyE/Q0rntro
FddCgTU5W++yoRYYzIkhRvZp2hR23BhzFujCdZpEgq79Im/nNCvHKXoAELHXjHCY
7himy65Hw6pexzUgVtOMdTgEeEVe9WrAxhTIfAywBP9S/B91gpx2ajB7m4BdROZJ
eQJLSmOLgoXlssT+TWR7/B3vdR2/FSCKf92zW4bzgWxItYMR42YEa3MloD7+/29W
NWH58UqwjGhKuc98y1PUlR8mzwLRQZQMb+TlYyBfvFkUXJGT/FAJuderML/+fksj
26gRTBU9sySxKSZUtFboQHDJfkuHVK/dkOhA4IvGQX3YRPhHHU/uh5tQvgVBggYe
NmAB8H7OwiWOYsxa1oiA5XP4rVOQezfe6UyrTXcz/++vC2lfCxzm24dX0vIu1ers
vLzJxKb0YudS/gKwcQFF1OMrWYgZ5ohtZbQ38BmAJBZ7B9F3++BV2p139xq8Lvo8
jz/2O54hdiz+Hev+Hdfy6+/gMI4UlseUOB12U2PhHVtBNmIu3a842VhEZIVVzBzg
5yerm9fmqsfRHdgZCYLqF1oZ6PJuOZIs2ZDkKo3hdjqXBCVvyyZUtqZehAhRZJg/
k6IWby4/e2LPffSVVsfSa4jqBeprXhYiavqLwvMtV9Q8NHVbyUVVoy1p59ogtRvx
RGIY+UPpNnIucuXYXslYkgnrLszPNg3aRAmwCBz6KmJgpgf8/W+zLWh4g/9m084Z
/UTMGuRjAmvxJpGCScHO6u4DCeegXpPFp9n/iy9jsxq7OMz6paf8ybIxDoMVmqhg
SFdYGxkNe/9RRCL4Gx33/mwGxFge4ID+duLA7STul7fAT8fGFhEWNeG1cHOubvld
+KxuuiYnfrA2DpfX21XD4z1Dgk9TbV6jaZil080Nyqb84yi0yhHRaZ3uPOKHw4qU
g0/6/nBEC5chvphlc33OZ+NOwvTNkc0RclCtLdfAih+nT78ovANOtyxZdtBnLeWi
b8JgTU+ZIFEoy+ZT4Map9RqB/1N+/avW6mdgnGZjOXwCXKfJxFHcYVrGo/gxrU/g
QzshEzHNZf7uj33UwQuDd88vWefJaQApbxTa/o55Rk87txxX9NOubweg17mWgNIx
5o2RCNbV2rCBwiHIH/xGvSigCm1QnXFmZmZqr5qFN/C4rH0fWV7ise+haY99eZJH
g7VUoFuAyKVIr/HQuHUXrcqgASCik2FUuTZNlptzXIKHm4/GL1iAcP1Y8wIjqezi
XyLsRlawXcjtzU3LA0csxMamDPUMY85yCgKG8ibXrgv2SED7Eb0u5wFV5SN/fvE6
YsuXQCjAQrK5/RBnzDipDifrim1Vp5s7s3bxU6tQSIHd6km1DK7VN02u+co5lIWh
Kr1bWnjissWXoarhLJdUY0Y34q1xr3jYGQFMDwInUSeSRYNQw3ka2mScuFqZAZeg
yUJmOrSsy5a/nPQDZd2hO3VMDWOeASa09YApvOFoSc3i+QxRcExnVNfz52rGYvto
sYo7LCHOm/S8jUYl07F0lDLVnKKC9smdwHNmrtdTwnCTCioeiafULF5WLpDUhum9
genw0BCyDKZG0CM6w0WGeepbI28FO3VZEJXt68pfhP2Vf0pGy5doJuohxIGtgQuU
T2laB6BUyuFaEm2nqEz86sMOyq7Xx+3P1Mqwp6OCypYHEFksVSDhJV6zfLG+I6PM
DavS9uK0Vufda+dePPRfc/wY4vEvIRB/uZo6v5kux2aX1u7SbnNW4HH57SEqxokR
fX8HPNJnj6OUitwZlX2Qg0EKXMnHcr+0DyRhKS8g7+aDgjLwEzlwsRigfF8OF+vW
5Smus3k048SdlWekqtt/ySKEarN3x1pb7hvRbv1+QecIdQivwHizQ0xGxIjckl7e
4wpxLm0jreFXEjJ+exaTQtdZ04WapVtFva/1pnfA+IIX3MgXZ8q8XjTKjmH4Q9OH
ERWv+R2QI8aPeS+YO4SAvdomRLKFpo49XVOPqNsfZ4w6ttYf4SUjkFsKUGwbFlwP
05e6xCH/2l49GMrenD/9s5DNpJn9ZKH3rRpiklKcTKacpnqXxpkxycvJmL2Tcapd
9vSBkAe4gQeAF4Yu66qSXvk5THX8WqiCEs4crFy3qQk/SMfkIOQXJrv31cygFsJI
85o0tYwCHXohFYLHe3o+dlH97PjOgr1tdXfH+F0fxNEK3aA2SuLeQwv4X96avn7e
v+e1tsLW3sk6ytEeNCr9BurvSwI26kcmH/woWHnu4g6gVH4yQzifBs5vULHM/sIy
14zjRcmZnzenppP8BXJP9TNzxL8dmhKKMkkquIUTKWXIYuKdzpIcw15WICNTswuO
irXZIltGQogngC972ThI8gpiJuPcXHbpxy+3rofOW826ZY7xZYstzuZf4QbUyJTa
jN4r869evjhXB71Ve2MMPyppzPA2WhvOecVh30ai+niulU2tz6Qq9YNX4Edq5d5L
SYLEqeuuxfHDRj0hPPr8voly3qwhSZDFX5mrnPAfPh2wMA0YW2uSFWeSIlbvNKLe
RLcw7bvzzlRbCnZkPl9MOCd7dljIcQRkymQgV/sJvfpFWC6HPp00EtR5uf1r/JAx
R15lxFbImdTwTNRwyKmel7rn9T886Ozcf5Upqx16I+p5+72SKvYmfCKT88mBAvKo
KJmoinvrRPgpioqEMnJKDjTS7dwqw+uSNO68nJlC/68dMl7Gx9kbnmpaGf6lSOcG
OHqe9CkAp94hM9Q9Gp1sY2rrKiUYJaE6ojUD5wYY4441MlXxsr8Qg3whrwHxzOZD
NRtQ0f02xAZpRrDV8J7dUQsp3Qek68ENvArWm/rLGOiV70lAjSbY1BnXbSwnvNf/
xZVMHfZ2WXloiItBrZz0R6rAQvT5lfEZGx+jBRFErRKp0aeCwwvVGej98QOVW04z
YyCUojCfPDKC37wBRhhjjYaDYgL1PLJ7xB/NkHx4eiUJCyOJcPcXyNJF+ElflGHX
yU94aLUGYAvhnZoQHqUgIEDMI1EGOMx8vDjvydm/5RXPOGeZ6DqGfGSmUT9HxDms
HLqM5qGBPzzS2JglfzZPVspWQhGAzCTaoqNf6ABqmox4dRjAIbBJKMk1wgTsLtDQ
QbOM+abdqb7N9K9BsSbYbIDvCcOq6EI+UorX4vznqQx4GP8oEh+cZDH4KK5Uwwwn
GLRqbQ6UE7TzFIG7fIqRIX67zYFg+R5J+ZofeJiMfD+o1d1zZSpWlycRAyTFVlf0
lrXn9X6OJZVRsyNUgNQ4MPIbRRZXGw3gYjQzolwIRYBEyPdZaCM450vgO5/EaSBH
TdrXCr++a2ksYuZRsdZp/PA39ZppomGeoUSatC7mQ8Ksjaxo+OUu8nDMGvv2xNkb
6vIL3hXgU67gnLVagd3bi9nQmgFXEeBVlJ/wYqadoM4L7SBa+52YqjBmt1fjjli6
gvUfygMzvC23u8axLXgfmFFTfSRCPsPPHxUkAVVpj95brTBHrO4IkCTLYlQJWy3S
jy7dXfjFAoST3iEtPbMLSsINvqmD3QQ3N/wUGcCJknurCSQFCsmNsXHBaCxze8cG
qjy5QVy4a6jYu1G76/xSkbU8X2qFKeMSg7sfy1M2L2ADQRi5DFMJRrBEVfuseIey
tDuRQCoGB+PPkwSFd+cYON1EkuJlBCl8CmcN6CFil4pnJH9T3dT25OyOFxvT7tkS
vcSlvMKj0IBQ/UpvWTFL4OpdZ1zJyBkpqyIF27e9I/xT9kv0WSnE88bAJtx9WR5e
rbh7rLONG8lX/6VyehohW52CTavevERrsh1HJRup6f16XFyZta37a9W9v2XJK5lu
FTioH9ATmdSquDYovMqBk01PmYznHfp+xohZHyzhZchK+vvt+AlKKit7nFF/Yll/
LyhDnFAlyjkCXjRxLSNBqXnIXSUuOgIvVYSa9YEtvbIVGOdQBm31SJxok6t8Tp/8
EK6J1blqPkg2Cx0QoK+H2JG53jttLCJ6Hx+PWiKqZ8Cx3WaeL6RcfST34fmgqG+f
Yx0j2N3BZyjr1y+sSYXucKCBOnRNxsfOMaWK8i2rjQeGMBwpu5KXHy/IbDS1Yhzl
bLIygHZfrGqE2dl3bgt8knJ9pK7rqogGmHgyZ2fL4SRXidGW1OvUREnOZ+ChjKPB
Yl28WU/2zkznDCUCWiANbm8OraFYp9+mZ+4aMpOz6mAj2p6ILMo9f2MV+1LgbsFY
L/Wd1egp+O665KuUmG4p17eaDKxSv1th3tv2jDm9mm/2wFMuXu0duQtaDjujqfN6
bCkWISGMXSgccc+gNtXahmJJg0cAfPbcrZPW0PhU1mSsNlSF+8yENM36L3hwoDGF
uCDcUfR/HnRH03QECbwt7OEgDYr07lKBy+pfY3jvr1X9d7ZzCMKqVHIbX74d5iKK
MiIcYvqSaCYjHSt5ZaIUrMxAZT2Bv7IaHsKGxF1Ubcnl6pXrbia/m9Pcdim3sxlV
R7tKLrxOhl2D/AriYKdyXOIaA+24cgdC1lzqF4c1gp37WpgVWMJD49UNSbXoOETM
9hIQFtAmW2eHQMrs/YI827cJhrvV/U+jAs5kipV0VEXZk9ORwa2v4W69eTOLL8Yi
nMBhvfIfQBIgVuddi0mZtUzNaNEzWTnkTiS5fp7ARZcZ6s4cUmMLFmsEPd1HA4RU
cYt2zVujDRpnImx6IljvOtu4IjxM/VLE8Ej/dNIm/Mks1vuKDMKZSkG6o6JwLitE
pXfq6Ni4F76zgrFYlPz4iZ+sc/Lw/OgHJ5TX9LlWVEtbtn3I46tIQs01FpQ/Z2/i
+ciydPO2MTQeic9PN6gh7+UOcthYl1OG1UXOLqv6z8zNmq9dK1uqf+WJRQ21HbLU
6TJe7vs22NhXvpxBrqSWzBtcBuvvwIaJCWQeruvO9/qvD2r0a8Mp1gLjcev7NpJn
ngNogookY6Akel9r7EF/GqegWhPHt7e96mOA0MAqBIjwGqAYkKd0dAwB99UscZ9W
YWiNeYVXQ8KYVQkLtK06PIAT+06ySAPYWL7ksg27kII/U9fIQpy8iBDQ5aR7CwQh
F1nE3Kbg3pICDs3Mwnert4nZVuD+VQVesGbKupTnGRl88mUHrNZGZyVh5v4NlfMJ
6waURxmHEQOYeT5GUPRRyK8/TAbbv8sjMR/SSlyahW57CDnaS4bOLW2TQK1Nyt2O
bI40KhGd8FNW69K/tHfWJnS0Cnh0hXI8PASHMyW/gqoeLJDsvKk71+QDkaEIyvFG
9pF2jgZrjKU6YQr3OpbIkoaGzLscxfvjS3hJInWN2/BduzaR7NHe9gEMfaUu2iJC
7i/dEN0swBOsKWr+BwRBL8yV7HJihmIkE++JLemwT/ZT3vLIyrjdNR4E8xwvQ2g0
3Qv9G+PbJl5IPBMUD4axnDpvHINopCEswyahr7qcGEgZewfGJ/RghuShthX637D9
1s39GuwyDfoNCfAA39rKdy+ZlQB2hdP7yUueAZM6VroQfwjDQ0wXHnYeQrTgtCS8
hZLS/DWaHUxOF9d2lIWA20lxPHXaUGzqw5c9sBLMM0SW70lMd3rj3/YvCU70JurR
20+ItWaDr6h53S0DoLymhh1IJIblkJx/5xBiqXqUgaMvJA83Fb+9SRgAkFm70Htp
1F5AtRzlX8R0TWPzvvpK+pt5HJpgNaKAcNUPQc3ozgOk1ICl7EvF6mrQ0xzwownM
HgD2kEFJEkKZ3IWMgVCxQCg+KDT3PKVRKJ/BFhJr1tVxXDHqwQe85ZBDl2gAjLv9
T7cahcKaTNYxQKnL+6NAKS/TIOcVeyh8TEMfbTVLuzFRO3yVCyRpmywhbdxz9zhX
xTNrOd2tZUco91XDg3gzHxrqCi0MA3H5tD0HLjjdFfykaoKDjMALlD2lRTA0X03T
ksaPtCbcJLZ4d05rdKZ8zQkuCzRlu5m7RrR0ym7LYlqj5yb6Ogkym0Yb1fHpIDvN
G8iWVHHiTTkxJ4JwrxFfAh+DNQsLtHAvrjx6T6or6OZlCilzp8Y2uq5c669BOx1T
P2iP5JtqSnxQIcxSyCofVG5UAMJwybEozvd4hApNnKUSAcsfJhSCguJuRq+LjcLa
8v3t4sIcJ4EJWwVKWXwOZWBXRVow7N/Wi2kDK9xhTfyKDnIvn4oKMjWD2O7c8l1b
AHCaHd3yk4c4pW60QgA3GYN44dRitqg3Km4lgQszEJMnYdwAnnq0pxJNgnR7BkqM
zRdS7qaeGqu/p9eLNiXy49AHOtE+x1B1W5hnrT2+QhCRjUo4c2vmabFBr5rXg/0y
IJFOc0la2DVnjhGwWPI51w3e5IfC0P7CFWCuxInKXJ3ptp8QdM9wulG7RWE8rGpp
49MSgd+lG+szXcohDqtmcFrnFQTi+ClLMbrN6KB2YxflQbstRwB3QNWmHqrOzNy1
Tb7R6BvvUuR1+/JBqV7JcDaTSHz+WBO72UJh4aP/JeLH7S92O+vr+KC05dMMw2ZP
Czl8NEYJjPDdZbe3BhjB7pAg1gzQxMsuaoKNQB9VvPpMjPA0bD4YAstdQU6iz/zq
SKBNbISBmi1Ygg68SJXAGwEYHeTveJARwH65Ks/JKHbuyHtQaglIZlMpjagmUAX7
NrFfMORCEhDWIwKjxcLgf3MEA/QKmmH8lun6Wxk/c7tm+XpcAqqQvCoMcyF2FhWH
J07w0o3NjRWZLIL3dRV87PnEOvE5IYP6BwCpZoFD20pr/ulR9Tsa1aull0oLWd1m
waZB+EnpYDkHlvtczXzaKaOcy6KAHnqkbBaXoeJDRCSJv6u3WTlsHLQoZuAaufjQ
kg30NWe1z2F27LnmoOm4V5V3ahpGqE/BN9CR5uuA1iZCyf3IkOIEyjKatyovov46
SQrPM6jt9nd+LOaAdb6Y09mEwKRFcf4Lb1UC/9OtKUFCPQBLXM39drkzBSc8Lryv
4YxobGKCVJj0sbrB1oX8P/i3Uufwjm7vV2gSZxJqeeSXna689hbAqinFFOKxoohu
8SyNWe4uaRur+wWtz1L0WNKtjlE7wGqj41OzhsxmvX/SMGB+YAiy7F+2e+yB9YAt
vHYOKLeQMu6/0NEgYdY2oVJq7I5KCp0KokfCPc+ltobJy4bv45Oi5QzV2vLAfXnG
4oqNPAD3Oj9oYQYbYIZfcaVjs92nHn9s9Fce5aETYZNGB5echDKUI705novshzQa
6qr2EidRApDPweAeOEoXETygzEMlyVI+1ww0mvuFx4GH4MFz71dUDCbQCs/ArpJk
nFRwEmLqZYh5vmXRms3/HqMg93CPZqDVH553yuLbIiROYsab2aC5qsYhpbLTNzRH
t179jnDv+Qv+KQunIr/riHTbTKqjZCf9qdKLGO84gldjH5tEHM9kIBS9N3RvcVDu
xQWHHaaqhquffKJYVyekDk6arbL1iw+woOPxKTdgzaoeh3iLmxp56pSwKqS4qy89
tPOSkTEi5n5bQnOs5XaFp6g6FtP+I12f5d7/NHycov0bNsaOyGfUNZ5H7X37clMt
Lvhvh3cK1QAPRw3NUkDRywFQ1J+cfMCn3zII1mcFtOaZ7Sdi3kdX+aO8CTI+O2Fm
pCjjTbHzW6gSb79Xkbyqvs2TUPaX0x6RXkKyLpeSaZO4xI1onD+Z8i252nubi13u
UBjC8KfTzPN7Vl0ef9h+ZRTK8sA1sX54+gO/WfnEldwMr/vLv09cvt4TDn/7DEeJ
k7IVr4Y7RRiM2Fpc83bjorU6CZKS1IuURb8xUsZd2llLnbKpYMWWp6rKSxChqhiB
TK5SVy3dkVV/cE810kYwKS8HPg3XcSomVnn7Fcaz2UFaey3g9lJnU//JzLg6xSOz
ybNfG+QnHhzZNoehvikbxUs9eWby5p0WbteXBfjCON7G39fN7hrL4sSOCP7gIJhj
4dbUj8n8XQOyJmEi5/l2CIOtUBNhsbHrW40qQ/2uDES1p6l3rjAX7I3lFGti7dwS
A5fWfGR3kS5b1mSyOgG5iFD2Onsp4qPQ4X40d3BTeRh/Onh+3UI5VsP0NEqRmSQr
bAIO1buuTQyLl7Ap4YXovG2wLb53f0t+CoEYFjfBpcv7YWlO4sd6x3cXrWtYM+zx
RMjQZVrLMI2/m3O4hsY3Je9W9ljfPLoHuxtdBM3AXEI25HG8qZ1BTrUi3jSnO9R0
+WX0jiv1w34HG8e05Dm8N6jOMw/8TcScqQnpiTZaRpotEa3kqA5X6MAcI3AVO6cv
wtuoke7oWxCREQegMCsQ/MCYJvuifsDAck6kwV5wPCUW5cgYJoBZEPNzeX3a+bGu
rgBsFU8oAY+IN7CZ15MNjwkN0RLQ1hlrxPjzpI40S7OMBr+mA1aykMn9tP6JHNPX
lr7JYs7Mzf8PDoFPcoXTBOWtLfSCky1IJxcLZcby/yqyJG+/CENXdadeCqk37m5d
7h+Yiin828faK/6F4AM4gwYkm5du9LpFj68FiEoXz8y3NIriyr6f8GdtpyYjAfon
RD/VHyKe3w311lKcmzCnJdwT6QdB6/orP+2aN1aenEkUdklsTZUKh25iVVwXb5G4
qmFx8maEm/ZwMHWYpCXORb5N7fmG59gmjDi59O9gd891iln5/v3qRshmByBYjOHv
BZAm/NvThn0FesEl1CXw3qlreMPlmK2oEFYCin5G0/vFQ57I7yJlYIsFTz6oSE2V
w6QDW+ww8Ve60gVHPM0f58xqnUTOkdiGRu1GomUQyDzmXQ3noAdtJrb1Femr5zxo
kmAEUF27rjPdac8bxadTi6cwFzoPPcS3U8FLeH00z3+6kAnNRqUll/kXGzDvYy01
Mx83WtOAq9Sy9P4TseAsbehw6VZTSTzFVzQ1ukw6mtN6s/21GZq0H65fmxMlT0/w
J6apP1NoPpri3u1tMdOfaYHY3HnSu33/04PUeFe+rytadK3xqbieTB4aZkgzKHDC
9SeY728pv3W3UFWzt5MZczwafEujaidUs+DiS6zhyDjBKpk2t6oaBUMj93h7Bpuy
yJFBuEGPsduMGyPVI04QmxNN6mlu7wSjPnLPc+CLUOdKaGRvrE22eJzHxQzFk+9m
RGvnXv4o7IOtL/R2SA9wXOIUF5B2Bh2SYoDHG06IlRBJfEjWmosFhBZ5n3Lqw6+s
C+bVGm0a+XaVlg8M3iKvd0luy99VsKuSw3/jzMjdk88ZfPBKDIGM8dk9mnIXunxF
aYIuorHyNp1iSjQWBcTTumlLJS/c1amTo5nWn94/2urcbiRa7vQaeKMXxlWr/fvr
6QP5V05JsStS8YCR5Gp2vZjimOXJSSHDFYxxBKEx1BlsbQcPZAPfaNK+gYYWn4r/
XWvRu2e8R8QzNYRhWcWevvrMWgHHBbawg3q6VNThASxKlNp4xey83Jy5+GDzPUBB
bUvZLoION8OkVP6Gr2N7JCb27RxfpX/CS5gkAy9UJLxOpjHjb+lnIcfeBuP4hI+c
92SXztYjbc8DOfZggZaWsAWQKF58qMbrVXxu0npcqLXLVi0373t7OFwdSPJINklF
0z1jqPFNjiJPe4pR7ih7CkTFPthy/ByOQ68Um8SPO7+b7JegayYOrPJCz6IIDPzm
cwemiav4If7oectG1TKrKYSHpzEu+gHgIQ8/zQm9Z4X+HXBtLNu4p652hcNOkTGl
4VMepor6/8wU/n/HsFI5u6qF7FgqmK3e2w2srReN/yDabc9HAzJfo6Y5i/z+Qq0L
Vl2YjzmAackSeN69SyRVoal+y7n7i5aBlhyyz2KwVdJGp8ahCRHRlOvax05xboHu
6Z7/derWWfCGBlb4pvVZ8uMHsbyQLBx12JnUTaWSKKEkxYNarrxalbTpegIYgLXM
dpGHwh1NJpyPYkjvDoEAB0mbbbYVJDg7GwYZEqBx5wkYMEP9ANv0HDWhcFQIeteP
0XFwCueIoQqbyod6O9a+nVTIyMmA3yy/2ncL9T8vHDcyJsW4E/D1tQrj5hHegNXX
QCwiGOPKtvLq9G8MpcR/OD+EQz91Q7NpMISfrPw92+Rd141BWEq6ssrPvmYk05WW
Uq/Tkl3WUG6g0poGHUqeF+5BRovXRjxEcusxzuKyCqReEDhnwIQpakl3SxwFtaUU
sQiVtLMVE8FhYVbXGhqHXBkif43oCHyX/vHDjPvU6D2PLsjo7K1mz2Hqke1t8HQa
TscyBYWgjPQqGSMZ/Ki4S6u9IcsixbeX5EEFtArmmSTuLiqnw0pjeTYIqbzKct35
bRIbccu+5uKYB7+1wQpbrKhN6rmwNcEsJKt+HE4Ku6Q49nlLQC51AfipXEM55VVP
c5C5/sZvfStW53w1V39UE/9yPGYZCUj0+Wg95CZ0DR9/WrwTFaG3+iB63yd7xT34
f+SNKBI7Q1IxVCflK4MzvemIFyngni9MAi2j0vcPqwkOQEh9J0R6sg0RHrNWeuBC
CFS2L+I87ogKWJlw7y74cRfI7JVijCZ3KfheMr0guVhqU5aD6m7gtTTCqpO2Frxv
3yQE3YfVI/ryb58czhB57MnPs1Nr5LX42Z5oP2/xwiI/EOkduKm8Lvr+X4gxCGym
KV/rTX5KVZAbQcKNCxM77JEW7LpGZZDCd7cOCN7a8go0ZH24GX06v3UZszocNAFP
gBsPM/nOOEubFSSW43qFqtYnXPo4PpU1GG40sVuay7H+2ZAtAjW2C3JLAwumorqv
Kxn+QFx/Jcqwh5N3YiEOyvbG+3RbRa6PWiTtP3KDuh63rguSeCytDCu3qgeVUqUH
t2UU8lpngNTHgW+0ctauLVHpE1yFl9wZEXBVEo/JbLBxnzKlLKxdHVA/CUijNkiu
uxC0uw6l/9Fc0Lq9e6mqWsjH9Cjs7djsHIXyzvmmhI5+FGf7uOxeZzLYEtpxK0fk
IR5kTLvUvYnEO2RH2mxYVSz695B9XxRUBKxH7U5JV1eSusgJUGqb63tAaVHCTFUr
TWCb5Y999SkslGZv5dVkEZJD/QrnlEAq1QFJnw9Eobt31x3dFM8CcoBDa5txPx//
I+YsgpQqkPI+jYIxu1bK0JGdvjfRWIm/VtpfpABUWGE+sz9Kot1BkQ+edf5drPOT
3gfnMtBTfxtoVahiz9QPXsRYxb/wr3sxFZBeW+pm8jnzhdoP4toiaXaxwrT1xBAS
E9KjNosGNCHZEkxB85f7fgkG6MgRlqDCdgy+CA6xXKmINHwmzmTKtaNudBSa3RdJ
cYZ+gYjs9nDN3l46zg2ONd4Lv4Mvpgh0S6PJTBTphkr1tfAz2RelkCC3ULHWLGi+
hB2iLkCNwlgn/XO0o/ABwZVdUeoOUTCr3g8wuXRDG/tjDuTalgrhhez82EKtqOUl
ihdz16sFYKYVZ4SdXdIcDvxg6I3BwVNbFtJbIxIJ6Pc4uWxAWmRapr9SgJPS+VHX
6B+lSzJdbwJvRxLmaJ8m/7u9hSOtu1Xxo5Y3ZmCK/HIlSl3qk3jcy0oCpbC7XbKU
/MwG9lcQaGLlbvmaE+uLdepo9dHBhRFv9viWMZeE/BrDuUhGh7EHNrmQgjX36k0o
oRxyn5hGATqxIdlG3KnDLr0w5fnH7KTgN3qjoAPOdVO2WUusaOuVUHAUJSGBlUa5
g8Bht/QInGdQOiKCaFOZ7Fry2U7yE27InlWy0Gv9TRDfoQEPSdD6wSYJc8j5e0gJ
6X/pBm+h74OZvlcy9W6zbAR6ENZl/l+mn4emWq2eSzuZ7++sOScaqmz8UQxWzjKo
lZ2Bw42CI0ssyRv2gVGr7VV2ISWU8ETkA2uEQRqxv1pUeZAnqOM+joHnWjyqzI4q
faZN8WyvqThUZnzEAlRcmBZ07RU4mQTqKUTDkUbuU37ehuRGVT2CvE96XDQVdrYy
apMDR4KVyhtnrdRYF2mnJ2iC4gkGRLsBMm3GRksFwcJos9zGaQxittTH0tuODdAA
De0oLeJryaAcv9GQMW9WQaaTYGalXm7PlBHdUvW0HnNUj9OFIY9n99WCerVfHVdl
HPquY9OimVYvIzUXXiHMt698vm1PF9Vo0fB4RmzeHZDS+JCei6nqL7eb2Ew17lgD
MFtT1ix9nEPaC8K4Pxsm2xZyaqXxfSFRsEJOGUNFl0mC+V16016pX64EuI94U+k6
DMN8EnGVFNKSRrltw8SHKax7riiYeINSZLKAR5tgoYGWCy19nGb9x0HgtlTuo+Jw
yEcckXlZ65cvk1PN+FizirEpq5ZANIu0i3vbpGHrcqdUEaOQ3XQ2eNVBxIi7Zuh0
SI+bJfS/6hH1ATwDSjK5NnoSkH3y6rbuSRs0c2LI0Kc3ecEX2CY6SjZIvXkwXbvE
eFdOlNUAi0ofMC3+mpbmjyR6EVQrpFceAMCPlkLIMD6KLCzVa5ghmYWo3yHAoDln
Bkfbo+zU8/V0GIg2kMi0TP+IdI+O5hI+Ja/OkEATp7AD73VDYs7Hotcrgy9p9x7w
1yzXLWv6IKGSZIxa73Xqtbcw7zVLrdkTy9opQ4uKaR9V/LfX3zN2PZTqCRJCa5Fv
M4aVRectnGtMqwejxMN4JGOloli877wbIwn5o2O9ngAy3n6Xtc3qKg1qW5lpNeQV
qE8b91hixhJEELAMS6LYMQRwGs7tz6OoakdB8UJGTFSjrZ3hP0p4YtNOGgHE2rhw
sNR9Lpk9uw/QHBpSCCkCmm9rVKJaHpvPO5GpJlHfVQkEpsSx8bAWWWpNVDj9CcUW
swZhRFcNkCnyQA4F1TmuLBUYn7iDGq4TLxjoy0xX5OHD0uC3uM79nfqT1WqIcGQG
jRbOA2Ciovxx98zRB4NYODX7S/UUw1SLExCrDPU0semHez0fqzJWjeCCDkh3qgj9
23HFOaZbebUWBzY/U/GRq7WFhwcPOwhBbBo3oYdkzM59V87/KLEe0Bpzj4x+JHfD
dPAqzAMy6Og2F56mKKbNBXp6OgFOgXBWHIsYO+fG6LYKN6MCJabcLvuplaHyW330
c0SBnYVATucotBlnUULRgwYmqLbuIouEOXgJbLzEWYLTdt4MpOsJlHxyzWDy81of
DtkiCf1dFX4aBIXXNM195GSeM1wlXIy9BJvCdSaB/N6RqgDM3h+vnyW5QqPGolzp
QkHHVZ4sJ2cG7A9S4OKvk+5g1uIvluNxIJPNYoPzzHUZMali4gtn4MiEeiOdyHMg
X/eECV91sJNwP5ZG02MtdKND2oVtqqi4HHPXvT+1Cf8GY5PTyNWZxBH0ekttwiWU
CUWZRL9oYqYXE9UD5RFLPhoucnLAhFRNe1NWAPLCBmIMoTWqM+O0wSMtehnzvjws
rATX4iBfqEAs5/ev8xivQTR6Reh5eY9iACC4Od6Wyjt1tfUWzRPYLmsdFekJN+0x
haBisD8hKzGZbdf8CfRXjrOyqnIt6SFYSyyCDzZJZLu1M3ZdBVd+20502g2KV7Fy
h8+rgCCurwYeC3yQD/Qu80sc9NzRSmRjLcQum/TS7ghF5svf2DkkBqq6rFTUtj+L
yV6UFAxRPn9k5sD3l7qodMOWcc0/PEbVV63JtRwKwQdqXwcZ8PZRe+t4ABGw8EiJ
ILPtwUEUorF/IAkG52h0rsmQiXqmLGkup0JhK1z8HQOjuLSMF7QUH9wuMDmIeLTm
JvCqMxaBaP1+HzPYH9x3AvjHPXLCeBpMqiicTfRJS3G5GdsvmbQA0SunxP1UDAlI
KiR/ZuA3phGqoEHQkW9bXJMHoVd5Y/kVngFqCogV0WGvJHMy2XGyByGI53SFwGfA
PHmbSvQ0E71puntghOjsuoBWx72VQIKVHHgxR7NeuH5Ed7zK389gA5s1SX2UD9wN
D3th6NV1MPkWhQI5QiArkhD9fjbomIDKkI0avKuN3uLQAo0dG0k68X8fypDVP+6N
IOPrhunKWswC0bsSIh6oIPLVhWPi+wxEAQtjUFO8bF3pnAoK2e6il7hvg2+TetVy
tpbSZfJgj9hLgYsWFPdx9bl+EiBWGYei5f93paQScpxHi8o9O8lhVQPeVBpT7Rws
6A3+tFXYRfs/RDEfHvu64I1E75cy/4q+WlJ5A+9Bc4PNSKm2OlwHxfygfa+tGwbV
F5hq1+ClqAtRWjTlPht4S0UINAUo+QURQ70iQ47jYmszrPQXDI1r6QjvaZylHaS9
VLxShuAHr+vBjMDEahbEj1ewZ49wD4yq7DjkQ10Fht6NLA5Plb9RGmdlD8KCMuCb
hyWDARPjDNtPSdgfltY0hYqRrB4Ph/jij2LLgEmfvwN74I+to56/00SDVtX/SJYR
PFLKFOPc63e+xMuCtUrMz37eosc4fA6g1aDwhuRDbssY1RmBV89P0XOLnt4wTHIB
zxepVg6RHQTKanF9NhJysfIkaKh1Fsng35zwSewJGH5CpOrUo+IiXfC6J4PGzD5v
TLJbXQhZEVPNzhVEvxiC/fb2tqK6BNVkhafmEqLifj2l603l8uMcJAWU6PPSvxRp
OKPMWKq4eGW1NhH0aJrpQ4kWURTmobhEKjKSILpZADjTbmKG9ESF3rxEXA6rVSMV
eKKB4htX2LWD/izdmIkqbqGeR2Vg7rkBj1qZwElJXItk49Q5eHQ5Y2IOksX7ECM+
TxEvdg19EqcBidik6fWnOtd3qCN5syOJZ/F8cFVsG0wp4Mc33UrSG4LKUuMAuv/w
/FsGyGWMSvUddc0II6T5vrBHc8sNklqeHtL2zA3ugkUeAtB0ffyBg3DgnK4BGBxV
AHE+YHKt3Vk+ircfHcgBEzbjhV4EXyQss3Z4POpsR5bdM6JoG7XgzN0IEc22e67x
uYgVcnAPPEqe1BuSAvxTIOovlzjJY5JMspQbfOgRvMRL/xzyyzncaF4oiDBWzqPc
QmiyvR40A3e0moICrdYH5yfe5HcDlf3m2u/A38+WR/3Gt8wrdDYxrnO+NSRThJKW
XYrrk1n5pOn2nGLpPSgkE+BqYZ4QUkFgco4GSnfqZh3i7avuPjM/GrWKCeWy2kqz
AK19DaMVxAfUBbHaYbpKuZcxNOrIAQTQ0w5NdkSKT2/0JOGNpmQTeu3sTcmrqzvI
y7Doot1y1lB4mROUir8rzEy2GlnEtxHELm0fw+PtNyQxbpeChfgc2A/kG1G3erPi
x/m7x1q33LhQkZnM0Q88AXIkXPHbGLSiru5sOcwbnBTtUt/bk/aa1F1asH6wxIiX
CID9Tdnt4t+uMVkgLQD8UrouBEKXnhbOSlvigjCyV38RvYibU1k/KhU6DgaMne3+
+yYhvD/e7x9VCenxCpZLTSW6kS7V31bHYYZiFu4Aru1val1KAC5EKlhtxalB7lTw
wIKqzRZe3y/LpU6FTE0Wh6x0/A7Xq2LqtvLKrjzYmXRJePwkJIowg/J8p8OyZtxH
oWfY3uw7T4b4/9gi9cxxE6NBbGLvZnbzym2Xa7kuwVsyKmrHBbvWeqM3ZV7NmXhu
Q8f2d7SqK3Sn8Q51eIXr8O58oXMd8wiwU2kNCJTLR/BROVbOb5yrVWqO/wvkxwtz
Jg1Q8hhcR8BPI5/voMQs0w2NMET+DlRqPHjnwTSlRifG5G1mhojhGq4epPc2yEgN
H7CHD9MM06p6jkpM39X4gmSnMfQ7GpVRaDeJwnf+tLZN3QLZ+dUnMxBtlVoZ22t/
xiFYSyFh4VgTdGcSDmloCgZF706VDiE2rezAkc1v33HT/9UENaiAGEeBxXs4Ux0K
TliHsRndsSNePUm0pAxXu24a2S3/6Be3NYXsffVxYOQ12Vca7mum2bJo31dGtRye
xLNK0ko8w87texek/tCAoR/6JD48GmiF395AdgdUNduNxIpA92PwhVP49SSePPgL
5aAQqCP7FxpMi957WO2piOXFEKQVhXkLBliHSKCjD3nhtCEw/tA5VmyQYaf7w3It
MlaLLYNSlV35xmFnCHrDYgcn0POP/rLUBSDfN0zAZzlYuAnCDMJgESCU3xswvT8M
scBcFyiz0DMJ5O1vyL/Qei26R/xQ3TbEGKNx6UV3bKoIVYZz4Rjz0WYeLdu6nwko
bFlPWWhWtkaANMPFtU7leA+UTfy8R7qz2VQRdtk+51t5ABP6Yt6riZzcnMV4XvST
XEdaKw/+qlQfsWec8keiRAtfEtVEURWwfhjviS4aV8MOqE5AaVI4bSPnHJ8Fy77y
rXWEUibbq+1J+jaB8nPeFY8Sls3IVvVVQmiQbBNWZfiz29EvXCsRXto3/9jzhzm7
9ECT+WLn1kj3x4fbkUxJ3P7Fiw8MZkWLDbPWJ/Q7Y0oz1SUbY7tekQfc0mIsyKtU
ZnHO1H+x7OoZCPMsGv4Kgk/tV8+sjuyI40CPZ4wniHWQg5iH1Y45BE/9sk97ikd3
QCFOVRUaM31mo2Ef6Sh6zKXDLfdo/qPyYPuDL6Glk2Yg/OEPOeHQnkrMSlm2NA1k
vwxrujPcn5KwtI2IWS8Bbq+iQON2jFTWoJq1/f3ejbtUnzoicUJbM80NI76wqP/E
qOmnm7nNyDJ0jed1/jrCTp0bSfCV5KIj3CVRQeizWhmX3JWyV8pkI+1GjTF7bKk6
RGrFE7QBlXjHPb4QVdpSHxsR5O9tG6/wbWdQf7dnKuBuvWLTqcJCKlDizFAkSpl2
jLEvDifBEA8yKo8thRJbjr90BZYdanWydKXyV8finkeU4K0KTz5XTkP/G2SmaRby
NhiZHcMgGfjbU9EFq3ucQ5mQ/X5siqMwBowvO9dy1fCfcW6VnIjzVsfEWPWP+Cs0
3lUTaO6KoZCqUTwPmvsHjOK64ThZosvWnul27xd6Qrck/bir5xBcvw8DiZ0XmIFR
X3WG4yA+m9kocjEekVwDVH2wS4KuZxsvzl9NShL3XYyPLaHkuGcS2/gV6wEeourw
cLAgmVXAD/dLAhKLSdQ+eJP9/FILHLOwg+OhYA/SITuk7/zf4W71E6MltIbCNKx2
g5ICPu6Sw4L6DIqcd5yBWer4roSXfcNUqJQugwSNdknuL+kSjxNLnc7xp6DN6+RC
DgktQuvTGWVWj4ut+7FRXLxwnLMHP0gGu1Yqoh8W3xq9rzdR0P/7GzhofVZPhVxM
eV/HwCuL2/IYqu+u0mBdLbVc/JagQMijEiHDS5CtAtweVhJTD2Rs5R5zzZ3PAeV2
SKPk9nhNDPDRENXY4zidOhpY7EoGX3ulMjShRrje50OoVVKRWtm2pRQwEZCGt9iM
8X+R7ct3Gpue6hmAPpSg/ZMZHP6YUv5M09bDmyFND+og8PIr4xPXqRkFY+GgcKL/
9V7FzfXuLjKMWzZ7W5kCwklcv3vVSYN+Xk/OAdvDwUmXWVkd+Sogtd7KvIMJ+ya1
AFGgR/kGIgsl/uNXH9tdBBRrNRTjtQD+/n4pAY+lB/c0Hy+0djSc/slWRFaHWKvg
J2nhG7XGY0JhsMGogbSFQBD2cK5mEHrk1NA4Sd8LYEL1mLMGzVvGttWglljUbg9Q
ysJxq2vfLyrHgxdiLCPNhnb/Zd4O+sPjvH//XhdYRkGGzCUG7pY9u2XYP5uS81vD
IfGWyOv4VAk3Dv8T/TZVj6s2MeP+3KhxM8ij470FXidz2azudC0rEziG/FiiRyYc
roaQnPvCOh2+/qDjj5Oj2oCBIbVpfM568H2ybzE5gfzrYBjFoYyZzzfXqbsClVCD
Gs6NBiYP3neQPSkBHb7aDxWurvD1VUT8dUC3mTrNhxr+EDyDA2uDrgoWPe/v+k+6
egQ5rtDnqtjNhzs8BeQCF2npoVE/pcuHD+4FBukjTzhAY1UVK6jHmBX4hkMmCbeO
sh8Cb5jIjVbXnuKuNY1NEJLWaoHNXA7R1Gbg+ighCcKfGSDxWyKO0cgGbX1Kc3M3
knBt8S4rUqHUZmadGberKAS/2NBdHCMK1NSt8OUiRvChFII3OZ9CyrmWFvr7Qwol
Lu3vyfu8D0spodAL+QuCbR0Poame1GkbGaEbjCBiUM5r1Edm1KbGvxZZ+nWZ21VG
YQzmf0TTxLqvgKlwTZEPeQvDrfzDPcJids6BDgiRL4soM1wAkpdo1o4CuSC4wkhI
Ni427yfM26zTelpWusjm2SMKa1lWZTiy86PqoGV8kxM2JLMjo52+BpbPYcWBbrOf
J1V6J9qT+tsqi+K0fxwAf3eCSv3lt50Qs2brPh+iQXQC72D3Q6b6kyFrjfImI7rL
+3zXpL3YUbHIlxm8wzwQhGL98KlLPiAot/b+KnPwLN3DHuv3GrgzR85GSRGmzUK+
Y6UbZMt/mwUS4Qiavw4qcISQsVaSBeVUsJp+RIct6yE6xLaRf75h4C+ghOvUKNip
k3uPVsP8ZviVFyhLo7HzxmtKKHnqfZ8+LpDsbK+tB6igMqYb7BnwxGhAK5dY6eV4
rnOD+FnPNt6DX0iY8hFe7oSlBS3mfmxqqn+Lhxjl+8d308+Nu4FVLusAlvZBpTbM
75B8iL3Glt9Ff9r8VR8/Jm9hx6w7L9YuS2sLLmixees5k9Hp7EvUrtA0GE7XYzxD
+R5q7bNBihVtJ1vswfkZ0zD19MJmyDjm33b9D5ZjGSxMbDIIdhul8DSlFRj7+p/Y
pMQYlZLVLL0IaQIYY8g3nNkAF+3Gf+mZCPyY5E9cCIw9Xid3oNZMIazV96Ju6T2O
chxP9iJp8SopvDlwjDTjaIxvNgJpcN7BhNvUsrzL3McQfvCG4VMjlM0CJ9l9aYeF
bY/4S272PT9+qEVTRUYeV4Jryy42eYS37A1OuW5irXhdBuMg5yJgSF9oM3bn4ZbS
0QnyhEj9/XRGD2Cjf6/m72GjEsw0RF1zBbtnVBIWcX3uNjviXOsHgeLh/mNviWYt
WGhJVfoofhVwia2a1P0NpvWxI7P9k4BlEzLNw1QGUV+TljHzQFWAdnhCLglsbKv/
cyB4c79nsMCHdRNnhR7cFyBdkZqqXkbioUO6SQhIKrF7NgGjrKLSu+XQKmmv2z5w
bTYTXQ1wgYJOu2HrGQhzO0iD6ar+f6dhwSQK9PM8SgH29TrUa9VZOk7iLIGqa6vF
DHBXUEqYjYpOkAJGt7mbK5zOV3QmT2u+y/0uLrGGD8PRSxfki7QjjTnBQwvrhr4V
qZkjFjoGDxMmVdfb4XQlkMR1fUiKAKYdxbDwKzGpoC0TvpqRj0n3cAF5jdq1rjmG
T6WD/jMh5nLT93owLUJosjdxRDz0tHfupL2bDSPaafI1HvzASaZlWqK4oJlUxJo2
TDwUkWdWZ5YiJ4gE95u9In+aU/2nRELnVjql3DxNnIYzOAQt5L+HXj2L7iG8WNpm
NHkal+D7XTNxxpIl3U+HulZq89FttwYH3FA/u5LIehCJzBI7Xy3iHVLKNl3SOfxH
F0FPl2Dyx8KtXN6unHgZmY7a+f9mKqpJozLLu/rfohy7AruULg3FEDIKlUpgCjZA
yATgoTB3UIkbIo9Zc7lKIggdvZLjRFQQMgfjDz7au5c2uzpRrQgELm6uO3xg34DQ
oClHaVk9AtBvBAZ8/wSlIv/E2nFlC6m7idDwEDLpCvS33xQSAONohBnPxoT0AvZK
lFem7tesRfNXxx6d4YHWwAI/I7OxCRjd71uNMU3R9jCJ9qlRjczcewhPAjk+mNCv
+PvTxpmdkRFCIMFxaXqREage0EMhbZAknPutFzIreC0RnHwS1nMOOqDUWy5bDni3
BjnW9ks/Jmye2AFY6L8IfhokG+u2JVyFzTYyi0ly/w+n3apMZXTev1PgmA8rRRDh
xXFGsPZF5cDS9RyBQTJbkbBJ/kTDdqbjSdWUFKPzmqCDNPH6yVL2YIXTOGErZrfX
h86rQs3nTbpY+Tk3j+n0xHcK6f+dG6a3S+yR7Hz6cJd93AJhehLTqqVGK6dg5S1s
WRV+N7DfOzvIRUmiF410URR4ZD4F4NaKiZDCXRDV+u0K0gUrv/b3tobmHf0lNtUv
obkd3UqkeIbZs6li9riCJM0AT1VMU31Oj8cLRE08ee19zi8rbIij3/XuntcIhDf5
ArLI7hXxBIN9MuEMdhBG8Gn817m8QiNQZi8/XyEumDTSbX09GclcB/3v8XhSc+By
wYQM/Nf+4XOVjYDPINN01H2avLPdZYaCAgaYBsaTZM6MrJUDVKAjxxMakapA20Dx
3ayA5PNEEXcAv8i5CAxFfY/NHuYOy1H8/d27TXaowBjQ2HYlcaeYYWS9KZTfuiXr
fS5xTEmAbW0i3z82kenlwiz4akQwCJBYSp2yHIa5KAvj4tfpLUsTogVc1UnzGgLN
YXPt/q7sNpoLnn4Gr1fOcuTx95Z/Lk0lKiQpZtnm/8jhs7Lu7Hu/qvkp4DEXi1+L
mMGSgPoPCFJsBsgM6rCkHYJnzNgJECi1d5MiOLtB/YHFF5/mS0oWsVxBSF+I2Le/
W4WmsyExwKqHPhOOynpeXbix+kwEGLRVIkNcBHXveXSE6TAihsR6NSFRtQZ97A/e
2Y1AgoIBQzID/QO6i1klZkRWNbT5h2yqhYmNQP4UhjqWzskUOzU+FPKQ5ibvjt8l
/OPbQ0oVNgHT+i4cmdYPw5P5vZb8h70DPXpbQU6yx+hDPoHxmCIlbifCc8bgGX1D
jbwu9YdmZtvXhiY6IoCA0UJhz0TLAtdJP/OT+22/ufhRk5VpVnHTFEMViLHG3pwZ
iKhjLjXiE2E2QD3+kWJkHkLkN1qU1UsO0YZHmsGaYavHJXYJxIY8BDzPDQUacf06
BeMy0kcUgzzPsV9DXp9O1rHgHxbDecwEhY7QL8S+FL0RfoTDyakLlW+OJ4q9SZPV
/tR5MxrWwWN2nKvpNKjRyMVxEFGs0pqA4N6t/vmEPg+DIK/if8ydcCzwtmEszZtM
bKPCcyzKmrgdyZfLyO7pzRKSjsKLvBoevSvEUGy27HdkuYZaAi9uZP5ty/B0ytcm
WwrCWqlZcDvkJkpAXOCbFMY6Uu5l7lhMqADxj4h4rSmLz/NsUDBuPqk4m0JfOtIF
NAQK7TYLOMGWho+hg3507zeKpksoWxsDoXOeYxT8a4RQwQLG0OwKfh2SL3ijdUz3
46Pw3JvXQd8KpLQB/bnX0VuLdK7AqA/ExRA3WFpEEyit7D2eQS0dbQry8MS+CvXQ
tSbZrJAWFO4VDnTWh+frDMm3cr30dD5HAeUr/oVfVeEUxI4XDTt/8LqOxoZlwbio
2Ze0pFsppw/WRAUaZS9tJjBYLB7oxef1D8AdsLmwCxqRATbKSfxI5Xb4E3W4t8Mp
3vuUnOg9soxsQ5H2MXyMilP8mG6sf35IBwa31RcjJ2I+wAXFvlHKF1bEW0KMFyOz
am+hCzmXoNWe0zEPYeVXMgU37b3Dc8PH5dzX9ec4EfcZZ4vnYqfqHnWX8MUvrAd7
VxFSb9Hk8qX2mBoz428uMs8qpXO1Heu30VZMHdrVVq6R57izAdaI1Kr9K/ImRbP8
AU6f8k3HYfTK+nkqCZcM9TkXLjELmAVpfvYjpbjsnrXNoV52DVwIoZohUgDG8CiZ
txOhOnwfSBBUG8NuaY3XeKKiHhbE/OxgyOwUgiPF/+ECwVacjP+dQsbTF02gTdEQ
/0lnEPotAOipQ1340U0nRINK97CSvxSbQUORUUazgt/4kQsfr2RO9aKCjLJUpasW
zCa7A6Ll6wB5B2BgbQbks8Yx+0gvuLXmw4KTZ/khU+GzTQgYBZIgpGmvuu16huBg
+9Q0xIjpL+5nfjNMW8dEGscfys8JaI+iqxRCX4Kba5fZ0hM83m3oQFHuTKLXgztE
04x862utay8aIcRK/IYjG65ymOCG4GEt2Snij5VaA5kq4omtZwATxgBiJ8W6mUjx
/TUe/ES4c/hTP6kVyqhu+llPzYCl00K8C4nNHbrbDK4JrDn8697H3XDZpZPIfdJk
fL6jwG8DFieotHzjLcVMot4GMHh7ZUS+8z1V2CoO2MhsI74oAIjU35drd92iBnk0
BmvyZzlolWONqWnEcfoFt1DHZ7OFC90DQTU+RUmPgTcNN7AS1ndVAr135f/3z0ZC
A448EP81LM+1bCft5VTHCQdYtlW+se8lfY4yPVGfYbhr/R+HgaE4nC/lk75ofU3N
MGbVI8TUp6L25H5AqbRhWw6YBEyI1DQu3V/VgqMFMEYj9Q31P9HXdK79T89HwOF6
AfBPz9fkTT733wmH5hP1om0MYjYjZSRp3KKqL7m2EkzTVxFkfjfvnGpFcsznYYI2
dIjuhNpxSMbfff/hjG+NzZjmbb4y5L2y/OKzbhHItclZJGdYzmMVc4oxbbgMio2N
k4bquEkvcNqf0NB/yQ3pr7hrbXXcgAdR+0QE9K21JUTiQWAmQJ3Bdkm9fwORQFEU
Xia3uQ5R5kWVprzzbNkm0iXL0YfVCEgbEhFXPduZZU+iI4KeQhtquxLqlYZD5kNn
5/RrIDSMuYuOXEImCsxvF9eKmoEgFZdjIXK9axuRmUF+SmvwYPCbQOEEgPzyYdQR
KVASCv3+sSlyRGw2tTcC1UFfuN1BAVMW5Y+qb4tbYYjUeEHQUOMJWS8Vy2SkZMoD
UWz2O76H0cS23pPUTdxd7g8xNLg4HXyyLJsVeOG48dxPKpzdLSkKun2ge8rP7eDp
YWbK9DUeUr88jrl0e9mtRmf4L6MNdGXUMv6uPKjCOQ6xW4km7AMT4dcykA9Tsjiq
ApSdNXkJg5fpd281KugBrS8WQG9oCFNT/HDiIuXtxpuIq9J1IU0Jq1kr1V9QJQ6X
qh/JXAKs37mRhce0PYzNebo7R9BBhQIksmD+fiaGqML8N3jcqbPq5Nbp6htSG9NJ
hgvyWXzKYVwFC0dCN1UT5KqTCb0jIvOXL1XYoymDeadPGOWjwRbabzOp4jlfseFQ
Sl0fOmGE192Rsa4++GTnQdphbbtHzco0UjWqFymw0SJr8DJ4kvU3qYmC1ezR4BP8
JfS01XLxcNBJbngnieFoS1Op41UNpVlLQRgiNCiizKCXssol3oj/9/Dricfk/Ivt
RyChWNarlfYtm0UU52zHv5b7s/WN71lncgYpIT+oNU7C0WaFFLZ9AD/+glpYtwj2
ZBWfU19o4HZ1Su/7qWtOszwxqqGqTkEXVicHPcr4o/TosfT1nCVAUEHJK4pTH/DA
2cenvrKnIChao/ZOAQOFVfltdKgr//LkmdB02HlA3A4lR+/u8Oro5NMaL2GJaAQP
Ym3z8cf1CT5qf3vT4+qFSk5fPTLYC7tS6yHNKe/oBbLKhk1HShUODUHZ9CDbUzfF
/nmixeKbXIemgJGDlWrI8ffDR6+f10OBbRZFay6tjSAyoMTOe1AcVBX8tAFeopoa
QaTXoO6+Qo3UE9H1xGZm4s+ZfxD9UTkWdqSe2ABOYSr/TgOYWo7NYnDDWYCS9KEp
0ONqWZmLMlO/yl3B9gv2rH0uAxvGpsOmISO3UhGR0q1EDMyykkV7Y86dCQ5ijuie
2q4WQAnB2iQcZ89lrFIdy8YQUgT0yZgFR4IJWGZV18YME9IQXZwZTSrmxzaW5nz1
xWEZX6GXWadZUnMxZOekf8N+mr269qKbCQoifAYaz+jDCwtie9Koz2KO8oC6Ymu8
lCv47sjIgMDsr936VrTgM8Ig4V+Oqlm8MNxrfgQ7yJakqsjg40SaiCGYSaIIUGcn
mXOkgIAkL8GlNARKol3BoCJLMjRQLkHyBoz6my0BUxjWf55cPgXc9tj21HF1dhk5
O+wLQvkaEOHwhHOCv7INSlZ/XodacdNdLfnB6W9/c2dvVAOue/1lFvtr2DHUbpmC
JOxmug590rICK6SGRvP6RZFS8WspaFKOUdlPtiSBXQIHyyshh2pPrB0J29KU3mpK
bKd7DElzG3OgkXXXlf83tscmfH2kWjD1wRirny/XkpO834EP1V/toS1zCdG9fKjm
diFczPJnxDBwv+m7e+kguYKhp+XlVLqeCI3kCC3BSbHvADjUDdROBZ9RZG2z5N3I
SxdSG5PdiKulvPdePC2ogGzPVPSn0fsemdyRT30Kk6M3vQRGyas1cxELLyv/8oxV
NKb17px/I8rM2nU0D4mpt3X7+XdfPI/0nfgdsLxWEtYM68yXLx5XKWnC56uSrjUr
fREfPDTUESoH5jF0f2pilYHcHG1sc42vcWMN3VSmSjemXS8M7VjZntNNc0hqbHrp
2knKWYQWzGvT+9VpdisAqYl6vo+OfrQ7mj4jhIsBiYKb6VDyv+Ajd+yI+1Cmpy4r
EYlYdTugFp2HjFvwenJr9vUt/pC6rQcDMnibSvkj4m0kDcBzYN5JyIxNiipSnsk9
bvHdEYTAMPtA1ntp+Tsdip2CV0U9O90xrajS6fADsU76jpx2U8syLt226MYhCjy4
3B1g0cklKxO3axgNIgMxpyhCQqcuJc4Ifb/9GMh1ghqlGppCJWRSMCDqE6pT2t5Y
nATEcuQT2qhjib6dyvM7fCkfExFyO9mOPOjMlsKSCjLulFPkgV4LADm0AsNAYKWV
PhcDhIW5/nZI2d3BIl+PPOgm6SZSs0+t9md28EpXNuqRoPdlxib3q4IwAXkvGSUN
xqrkhrWyhTJox4liSg+Ot8EbthFRlpcF3HR8frJP4tGCaC6QRrvF1/Hh2Ly/9EtG
xTdzNwLBva6bncPvJVFi34QOKYf+6/RPob9GSm9ul5At5qruRFSQWm/Pjhj0YVFO
w6Rez15XEHIM2uPDTn8VploGeMfPhAhYKohdTz7dU2GViqAul1em1UMc6BKoxhSJ
rOvzn+5ZbQU+CNj49/5rKPiwF8SW6gqCB5b704lNyv2qi0Dp/Tn1c3aIVprWJuOx
Ao1Rqw5qQBititJl0OoaZiELHoQg1e1J6p6FY2foMNc9Af3Krq8Hzi9eliT/lBrn
UypVcJWdv96dKsTQYxzjpcwMJ9HjjOb0W0mWUE2YQviidoP3OwZasLqzPPrMWQjs
fuiE5FvYUDP27RVRBfp9VjI3kJsc3RL1SxseP5+EW2xaE/K+J4OSO3Js9SGNpIq5
xK9rIK9q2i9/cDSGcq1X5DOFMIMDtpa4J98lGyfLn+AMev/WKZf1z9MFkd1lWSm7
MYD2oaNAE16hhp8B1/VWEfDHRoHpwKEDPyrnrIKrIE9LGNxFtdQKF8oYL6CL7McN
Et6ZCAawDieL/9llmAFUq7gQL2EZ68Pc0piD7kDCWh0bsRvHizTjsLTl+kxS/qNe
TyfVXP5+9NjqNI+s2l/wMhBDQj0Gyow++spLcvjtceG87+v4f/oC4QTiOIWDXJQO
UoyQe5L0YcXkAK6gwIuyK+wHtYKkpmQ0fuZdyCaYvi9fq1xas67mwZ7M6vj/Y0gK
kY8kqVn0WrlMfKkBwRxOuAXaSOpaF3PLDOLrdhPWTAz/u9bUkoMYOQ9nn8Vfxssi
twOyufvRET7zy2u4iFX60ehK1n0KrrmZhfr1y9jozVIuBi57pv6vBOXbSb2eEO4u
FRmG8ZcQcfWW8BSzGECbDSnuydfbF8aWLM/BE+q85XXv8+x41KddkfQV7giJF0z+
hiImNifz0+SNb3tZXo96kA/5oNrS2zAKvgd0ZPb1GsrxEmaMBTAFv3NCQFxsOl/S
VOG9pdD8Bmc9+wSNSWM3CqskYBEPD3OoqZzOhxoZa0NFruqFk9z2vedb6WHk4LuO
6SV5+Hx7wRGHO/n6ISaA73oYiF4XP+mFq9tuzJvwHJyYb4t5JPAyVWMZkEWSc/gW
Dw3C0HfR8d+RjiX3Y4XqF2qGA3AnnbTSVYxlTkkJvfTjcyAsTNLCORRACfZ8mNxP
7Lp2d6vfK77mOTS0g7K39CTsX0+4/apF+DicTXk9wFAllVAle+TEoFtbXFj80hJ1
5fSlikIpff6g6/xAKScEIRle0clHjI3Q14Vwu4z7jAat/9Y8n3Lz2eWkkQULB3+U
OQR51O8fHlhp+FHWMT03YAP4oGHghhKSjVpBKUb+GfEkOI70mPuUbr1/FG2zPGAT
dr3xo7Of+/OZEG1SOL9jS22PLo4ZDJAhvtykKq0E0/Xp8yCbthDeEH38Hh4nVWoP
iBN7Y74qkhHlEpZmt4soRUTlPZMB9uOG93uwGEmYg2HdEj5nPbLAH7M2M9lthcvx
YF6+MHmEOUOJ3duHhDtN25LjkK9itmWWHXYI5dOrqGFhMk0Nj+XIUe+DOf73LMen
SzRQkYdr5Psz8CTvBCPvZrGufFGi+CeuIbPui9fJvfrSd669/VT7y4YYy3tzHeSc
++XtPetL3W27R2PbWEX0oQkbE1n0yJ3DCMm1F29GtNL09EPELFkiF1eNuFcvQ1Qw
Q5zPnek38h08ZgUoqLRHqdVGaOFhLEBZ8rshtN2hmqjpAPiC0btKIxq2059kTVt0
gXFPSPi/1gB9ZNF98UfHFy3SG8m8OwsqyL5XoxcqXdKsLqbuyb1pcK0q0U7GM99D
nfxwntGI4eObToa/nBXFbKOJh7KNYUpWD2C/85VZaRai0hHnn+DvKGm/M3pHbOjB
NC+1Gd4/P7u/1E1BLcMbJYTCNJltmJDsewbbo+a0/c/jT21trsPrYE65Q9BgpJJE
XaCmsMBCLKdhNhQuegoyN7iAq5A9H1dzqFA5AdEBwzyowPfimrlCtIqfnoAYsbI5
JL4zCnSiZlvgoB4LwQ9O9/arePW91rh/g+HoQ3JlT1/m08fQLRzHvuN0qLC14J+G
4VBuDeoLUWY8HyGvrjafq1nmm9LwTqqpiBt7Dc4vnHWEdKOeIiQ8ZLid3EK5hL+3
B5+jFrfKeEeqbaeqgzI8HoiGm0MFzt2l+zC0v/lQ3tHFPsx0J8bNfMbr0jgiUyVX
yFItuDRJokNAWGqFKfE0u/Rs+v3+dfdQbz4NpPEulsmOYAfUPS9M9lq6ZgkRxnxU
9bzUQWfGJdh+ce6uLUsnM0SgSHHehTzU5WqnyKvBcp7c+U5HCew+qSGOdzSfnrM0
QxU90HYmWThKj1EVMSy6EBQITTyPid+32/Sw/Zr1gducIQOIcBKSM1u2G94D/i3a
ZoIbvuuAQpr4/cI7jneBWhXp/zqWb6dY5hctSvW+dVtsOVKJHD5MupyMqCbKy8nV
Gz2E5oTjPfBXSrYrl4X8VcYFbbwHtrw4Z2saW7fWVsWy4sYqKqtvfDmjTgtOivVP
pmbE3vostoJxD5N6zrctNBNiOnmCFSnvMs0MjANlBCNJXeJzRh5tx8KG0EHjqIxg
6Y5ZeAiGKvdD752utGbfqxMUMA+V4+RBbJEStVKmJhy6nMm/uBqRQAJMb9Gv6ma2
6N/Vu9BQ7a2+T84NcrvZ15C8MAg/5oPoqMwA61niyZf9WZtRC+btG/HNjntq/kVw
f9aI1BZ4gq7QmOf2dlbT2ksUn+4uF5bPKk8Q6NLp0ACJhBIwWAh5ARobCVRoO6sy
r6xAkUMiNmaa/baA7Gmo5XMt8bHDZpVqEJAiWe1xny6VCy88N4rLt6yeF/NylBWG
fxzFVUgyaD+1ac0ELmR2FVkelwuaIv6XruxrzQQ3pzJoy879/1wTUK+rAh9UreX4
sxKkcf8jWcnG+bqQVPv1jz8r5Mwm3CXMRPz08t0rHpBHOWZUSmTwpfv7foREXj9M
dBPT6OPrPdY6r6GA+epjvsExHVth7A9Hl67XCVObRGQ2BkN0chdOYMJK8PCALEls
eiH3OnO+ytalwSR3Pr4KE/t65boNdmzWgx9cJmTP7ZzyrXu0kuRHW70luEUnXJZS
nIoOhFUhgqab5koEXQV04ZhV8m/Q/WV3FrpLCf1DGb27O252aJQZbREsaKJnyd7R
YZsPzRlm7pcAWjOMyLt9k4GuadyfmljCL3eeFY0QVN5FntOTjSvuCDurwEW2weOV
sTEDRlfMo0cd/EHnjNLvGyqP2M7Ay4luJbTuhk/+rgze1ZJb5tXIwNZ3H3NbYQf4
nG1nZU/2h/y93ZSR/SE+O+DlaykFreQxwCRFE3lMIhs11OKUaWy5c881K6ntpQaa
tfYSkW6RWIqBmm3cwGU4zuCQ5SNO0d2l5ckZSROjjpcm9s/lIn9UXFkTvHQfL1TJ
mXE1vtmqbgYy+nt06vag0zssNG7zgZHtmeeC9XyF9SJ103syB79x/ZREYOEUkVqY
7WhDSWwxk/cagFbEJZhFLAiBhqkFosmqRpq/bDYrn/AbSnwHf/yICAyn7Vl9+Dnd
1VYs7DRttn+dtIT3p0kbUXbNgfOBYhqR7SqnXaJyUJQfSN1Kydbf8efrLGW8gKfw
37PutFMMPG+/HbcwhEOIxxSXpVnhxva1o5aPX8osNbvenbmx+g0MNoM/ydVCAQBp
bTQnDGSDr2HZuxGk1kHKNNfaHRiDPu/BItCIp1dJQV7mctK3TXUICwYKTIT54NjO
SShitGtJmu5rZGkDObMkj1A5xOG5jp9rTX9maDjOu0s2rYZ1u3hmZQjvLz0i6GNm
S8slLNbiyTM7+SvigH/icejzTOVdtgViFOE3zMYxkwMGX08QW32FjIg9n64b/RvT
WwTIwqE2OElqPq+dctgc5c0LOhVbtpyL5HMYiTRF3bB9QY6OFPrD+fVDUQZbJcNp
DUup8pVdYj3UW7DNhCSXE6LTuA6pdnPP88Ve0y+fbECzmxmneCb715F3LoEUkE6R
yC9h+wr24kqZqQlceNcr7b2AkrtShWKqbOtw7iExKA7RpsV/bGplmckRMyPWN263
4awQrKbhoNOMBqCyUHm2UUICleQXttRIEVGSCwjlXmaIUsGQZgbGYnH8hVU4CPWh
CPzTqJtYUPmktWPMSjUb/klIIVWg1vf+UR2zCblh4DdmuuAYfppxXy6FNIxgeYsv
HBAsFT4pml0xZDTjbS6VNQKga7HJqy78yUySDeq0cxvkw5jehxrHCHWaHPE70/Ht
M5qoA9vHo0aFxzNrZ7bKovzTBbizdydypy04b8l7lzrvyMT/shqIxlJ8DZdY2jci
d2C+wL+TETjG8JjPqH2YZUHBQCDUTlCmdkhJibiFI5GiwPDSFoZNVopL+Wdj9j6/
F5dy2AqzKbdcO4vD6rx/j8RlMMMXB+lnRrZJm18QcFGkUpmAOo5uccJAgrcHa2B8
0IoEYFKg6RMUtLXjEtXyVeVBdbiKnvEhycg2xO96X7mzDUNxQ/BFMdpoiYhFUho0
bHOQaUI126/fjC2uUUmA2INEY84L7xZriqSrMohpdkWFIW0Hc6fcAnTCrJlISZOQ
s67cymMtUUk0BFT6XjboHNT8lwqy3txKS8oeXJfBTY8JIJLDD1ZQaOaF88qayvnZ
jH8g7EZ9TFPVQXjs+3eI0/O4g0lvhGqbqr2IHrjR51aYNnCUC1ZiSErBwSWyIDY9
SyZknt7PkEy6ubKRyzb1U4xi+dljv9muZoXOoqYBpn6UlCCEkTyxrRBSUN3xYOYo
xYVKUKvBXBFKAx2B/PXXphhvd4D9+ohnruK+mngirmM6RwCaCh7rtEViDeHR3ZOe
rkdyQpC2+MsSj3667XDDJh5BIej2c4CcsYB4ODfi0iUH7kboGdWNSxF+XgefITOU
pkpFL9UhYsraLlHRrbOGLULYs69LuMHGOLBdjWBA5WFEL7kqF8csk+0Hp50Jv9GI
hFBTxlZdFX2/BXPzCb09TNRwT4YtFkFRzI35rCGhm+EaNFzWv65C1/mx5oua9CWS
LgymKBEXzH70m/EtVNecMF0iC6Mh8+/m12XxZz7bSAAoKQfelDzHcr2vbSBu35Wj
ke9IlvALZvP0ha2PcLo+Fh7U1zWfn4wgVW2qKNOgkElh3AO/YTlbotQl/mmn9rZp
JP5mDLrdTdb2oksDT1Da7B8OGsxBHo/jYbXsXhYiOMS3JjERfc3e3buMbfLvVx6+
kmhvVIEccb3qrtsxqCJIYxwAC/7UnTAvIG55t/82FuFfeZtsiLaxl8cqm+JKMzxR
BirWjP3nDUcmyuibjz3fGBJU2zTAk0NoYuImczHKGn8zmq2CY/SLzu6a1y61sY03
Q6/aJEghp3NxDXwEmDB0luCGHheDSzmuWVB3AjHSOH8LbK/fP1BuqMwFL9WyUlCq
OfNGQSZ7RWsTO57UZNpYox6hTNZLlGQNE+p2Qs8EtvCA584CFtgmFpWyfHwgO5xs
gOpW4GJtWjLuu0oB1/b/WT+rE75Ep61pnKbPWpm6/Ntn9XkE8yCpU0TtOavvjYad
t/nxpkjpSs+oc0BKa2gQ/bZsMMbivWKExdIj5r8JZFA6T84pcAeHKvQcVC8s/j16
BVHdydv9ewTW9E3lZRYnBaFOuVDA1wvRhfJ3tKcHReH7/Vus7GqTtrQjYdGV2/dJ
n8dRCKYZ7NuA9MDpYFcFTeG8hW7hIdG9xKGKVIG5hJdquRWipMoOCjqh+w0XIY+k
BiFhTKGF8z1iun1jJ4dqLHb3Ox5WCg3KUxPovW/tz6TQqO1lcgbbd6Pe87dOSkaL
jeubS+/6iD7nGG4OZvUWg/A6y75/o/62QDFwkk+S/1+031mU5Gl+nAQcAo+41Cec
/9zkxsp9Q0k8EQTuLC6kvyANSRCNXiIaiPp7EOdAqMfBogsjbDOf8FkD57LKyEL0
k3YYl4L6S/Jl/HJQGsL69gWWKoNA4PdAo8XuXzwikBqoum7TKF1AYtcP3x9L6ik0
MxhhPtPaoRmj32ml7mN/uKmTj9pWjWPIiVs5FQ2qbq0RPeSNVG/nnZKHRfzBWkVe
y16BeAENg9ufsqzlHKeszZc4djwUiLT4XHbVKIOVQG9FRXKFE/OHA15xRwe6WWRM
dTqBgZKYh9yuISgAZf29EiLV49Pkynr2zSJSubTwSLcc7Sm75TU9TrB0dUTcrbQ1
dp0qJlyBoZif3pyJZZhPbTUp6bt8cQjY//AO1+oT0dMDnzfaOguRr2tlqIS2fNXo
5gagZ5Mry1vsa0gENM0leEXmMxbPV73j0ySUJLRVhdor73W7BY+4UWDptceHDTGP
+hRxL3f3iBFq9hDEGTOKcO2eg5cuql3PGMDqbkkZNNSr1YkTUPcOE0jqJe8feI65
1UExLcmYi9H3/x7VnH68PzugrtlGssimaY8GYxqiHkTr2MW+ENY+ZFOj89+CjMdn
3UKooDJb+qsDNbW/HpZ6IdQhJwBjJ8kCzFMFHdK4lN9fONzknujvojYYryHvEdk7
yyFqpJx/oMFzJOETzLaCKf7jRz2c3MD6bMArPtcpRO7cfFVpybQibJWLi6VYla9H
RS/tFEZSSGt5hgC2u9K4lw81q46UfMckHjT7lDxXTe62ICXyuub3o4FN68w1wOfc
UBgtj+PneqjdOznqQihOk9qiuEPL+OteuREX/kKQM8+HD46xHqrChc+aYM8PKEGn
RiOSXNGBHhEBGPtSp1vQ/szNL+WUTh07oNiGQJqmd2k8W74H0F96gtY0x3t/eW7H
/JeuBngOLvThJuG9ZBX5AE5t3qgIo4V1pYr5UmmoJr4p2WqWvHci8ba32xRiCMCv
iVy/i3OpjKA0M5KSphEkfmaB3mq2PmQ+anysn/O8S3zugXqrbCWPHnVNrh1T30QH
gPtr2ziQZdYGpPiR3dThCpqdF3EDmlbRfoi/W/LcT3CWWHDnNaqk8Prls4dSNNRJ
MatlNZYpPkYwmrSah/Bym5+fFSnFk1KzL+jQ4uR6V001Tkz2zDhIf2ih/CqcRReM
v1s0C8VMeq38UD12FY+K1PtYGRKvzatMY05QTTAd2WM39SUOsgGpreY91TCSlh3g
6WkCD2XtDnrYaTeV9i0JybW2PCq/seTs8cAy1Q3vFd3MYZ7qh8awqltCjC56nRm/
CYgt2qNofVMQpmkxAcuZSFfcAYLdxqGD9JOwAyzQho+JDeBj3BBACublTZ1AsznD
h2Mc5Wkkjz8LniE94vz6xZlRx1jVaRQO+WlYcQqG0uHVGnlkWeABvmFbGbYtCww0
X/cns09us0yuBg+MZjQzon7JqxdApP54OSXUzHbdKBtHG6TzAMghN0Yj7h2fan0I
QbFnnTFU9DSSeXEGt4mAB8Vn9EXaSCnwsuLM9c9Wg1AbXbSNSUQatLG3iE527Rle
V32mOjTgKTQv0KvfgXpIkrLbs8WnMThp3k3vJTuh0umQu7kcP97fxYJhh0xv1MZ9
jHJjw0OS9CV+uySJ3HdSessPGDjUhqwLwdp23If6TB0yWecTPyWOvxLEeic5k6Z9
yy2X4wMJ8IHE6ShFJz5Ei4/Y0K8kUInTwCS1Bv8XsCg3vWYg0OOIIZnlK8KmUIUb
A/LTiD8kbDQGV8YWOJA8SwOuC9Q6p7yFSg05iKdj9ULqKg9BYuST2XO7wUdPdyLm
0i2AeGPma/8re8affQLjhOEqfPWoxL98hJtqiicd2G05uokzpN23gzPs8zzuMu/9
4y2wPHG3JkaGq0Y1dNzTMLpqXMhlmRiEZkwADnhj9Y/6InMXFpfM3C95IySxuMoU
fV5INb6ib/glK3qvR2rG3LMfCJa8Tf0XaADhHOF38qlVxQo1P6KqOtK7bPPucbjg
ANo6J0pptIRc73VxYY6sd0Sej58+lI+ZiMydEFrg2UdNjSHAdMlZ9+N6a5gFhXEf
teeP+77H9b8yh/oG72ntjzNGYOJTbudDwE48MSdWnVvPhIHcjpUG0Fr29av3g/4/
syCY7U+dbT3cyxAD+USSYah/qA9NKSIcIi/u0pHH0VY5SnNxyYoCe3mjybcD7YKo
7R0dle6jdhuXvzP9bAMt5zlcm+e1hpfsWsuYgBHEjEdKzHqSpmDN9X4cqwDLI7kg
/xkucoLBswSG+93/vhUxjVqLNnedxt8SlJUW2n35it0TGt7IjKSiQBADbRhtQuD2
LNXFQvQD0x7Px61v5qJlB6os3va+O4fH6V8XAJmmf3Id22WEYqOycxNYQNapAFiR
0ojtSA001RjdzgZIdwy27tfmqarca52MsLHhVZbUpf8VW2CfVTYDJEzdtiSQjW8u
6aB7lJGSa2wXvSBS2gmX3jT/lvpONMjhLfdTZN4mUOZa0GYJABct9t4c46uRjwbz
iRXeJhDitgIlIAbGAoXNKJMdlNalxBb++qS3FR6nOF9ilQNdhTtQRmQc/2EYQLlm
Tst3RSVPCRcUTH7AjHyg3Mv9Hru9NCpfXmfvdTxXjSjPRog2bJPpXLmKpEGw/GFo
RQgHOub9GJ4uPVtFndghZj9Xyj/I7kyKz0XAOYfbIVyLk1l/LLzBEVXIfKts/316
tse7vCX5Bwc+qb/Ui+rRnHS7jVpWrA1CDpner+VOmh9NRQBp2yYKz/uKUeZbTCoZ
FtahDtnAgfEOC1pjcOyYoKCWVmofkM3SHN/gcGlUuIste5sp/HSzDYDCXhKS7JBZ
tqFlWtuT+gm8T3NosmXg607xZZu4NE1yjr35XZkuEc9TghRu3DR1I1iMnDSFWULx
DxMhuUf0ovlTzYa7dGVO1qnrBIYjSwUXUIJSpa5cLpgwCG4FhU9DNTbST/+qAByv
89myCKgmOdCLPipdY+WaAj+UTOwC7EqwOlgUseqQ2vNl5bk6BNl3mZpiZDXNQKvA
rCjOdA/z5c4P0Cn2u6bBttExLs7Gx49Q6cJNSZ5Bo8CC1UN4Zv4fAsQW4Nmss9DI
4SZYh0vMGW2yFUhofmVpCC6Aqffv54j4lhPB7gIJbokre2MIAyyhD2UeZxMZ70ZO
SlDnjbC+fgpZlIhvhdjSBM8hLX9qscNo8luJ8EsrWVbhx4B2gb2dxViYeeUt70S6
8GagvqPHRvOcDGS/E18I7weJRL4xQ2hu0QNmHoyAaPn33HSlgp4wjr7AvUgI/00U
tsuBjPBigT3p6oBGCCqqeKivfB8YnxHEVk09sUVGoh6CNBTgdvM7sqd+0aYgnf6Z
MsB0sx/6L8yk1urpVimQH+Gq+/myE32yWbaod6uH0V1Ek30hfIo6Q22WxU5R5ZDd
RaxvbtsYlO2j0WfUOLZcIcLhrK+PzjT6qKI4s+7fq0oh2gO8Xx9lGOULnLEhDoZJ
JQT1OPru0yBayA/hps/RLCDu3vgd01HcV2URPnnaACTIPwgbelvioQoX4nzDEX94
7TDNg+Q5pNwMqKUipYl88fbSafs+qi7TjPueKYvqzHzCNQfrx23F3/KA4q+PcurH
ilMie/JZe2BBP7Qwf+ObSX69o8Rqssm71mGH+Xl6NTmO6WS/rOAK6etwyKwW64mU
J3B5/z0VmNnBzxJILEN1ZDDchjJ8E/3d3fq0AQKOu/OEQPOW9bCvNTNjfI7sNEd6
psFDtRdAc+zMmRsSQGn4gVJuOvms1+SNbwdDuVCPtmEfJI8uewhJYWtHeS5JUyH/
GT6KMGDR8nTAb8HeSsbdCKuXW7npwTQeLC8BC2bQI3+HaLuCINWucY+1cSwSbD1q
t7/FwT7eT7TXFPM/bsd1K9sbbVMHOquAEjE655d3HD98ljpsi6JB1WpiEcAVcF1b
5IIf1GbUTHdX3HzGG8aaFrS0GVEdBuSxHdzemN35zSrTHSZO/kA0QnU48LbELuNd
TxLzlHSZhuPyaW2gjZqlBFHAEDrhxSQjhMRO42DVer4flb/5quSfQruwc8Nx0LUb
C5y5nu6lKQTOZnOBxac3vRvQPo5Yg0L1LHnGN+nrx6CvijcP+ggr2wCbZ2O2LUKh
XPXp2o80UKo9x+NZFLKtO86uOW6PTVAnXXPiNbfo9XmLqYnGOTlbwDTcNaEMJoGs
sRz8OTQH4BPH/O63ExqTp185xjY1whY7EvlUZffpPgiLeypjFrd8ZmGYwDiUqYri
JsIzaQr1zPDubsYjEpWsFTUrApdikr/SldgNwJIFSHtMVlcVnV40lLuzqxuVbTQW
9aMItRSYv9hp1d6gzjrZtbPGmqbQULq/TQP+ORWrPtcI1I6jnzHAICsLQYuX0OXN
9yq3TjA46/SfFHnhcm+XDOuYJjbFj4li06VkP0rKv4QP6I3jZ3UmicOtIDtk271A
MTK+8PL2Vx13OrJ+gJ1CV5n07U7dmp+mF4oyuzDMPESQvsEKDK/y4vHYYV18q/qC
G+D30K8DUsJmQbimM9POqtrQAULnCBShjpZiVaMTARtrmYpvDcoq5Wp0RlBfE/lr
A1m/TSgEUPbgkK1+qmL201ldTadNt+2j1z3DeJz/sr0+FfLWI4KAJoSZWbXNNSyP
6oMhFS31X6vqLGCXjLvostBaWRAYH9bwybhkQyXp0ogXiFFxyAGgUyYIIcc88LHN
ygU9SzFtjF7bXLTJhw4CXpG8RbQqd+oxQkgst6wiTL8D50ruGtFRtycddSTfBUZ+
2ngggJ8c6kQ8RoOomrH4lj/Hv5+dOPp+EEqAQwi5nSlExxdXalkJBajHjPPbYVDV
c/5s1vHwbrYbiGT0M/ayGhGCRnspy5e/bf7tyR0njj6K2HjXsDISCYAyTCcdF5eU
CbSz2ZOAE3VPUZsPAlEv/ZmF8D+QswSgWuUVWXtsxKmpEk6Zl3TqMhF5NoaCtoDE
j/DrmyReM0cPYi1BUITTIaEJZirwuOcRdmJtCauzzqlpBIhpdGIg6T/r8lW0rW3W
qp9Ki61y66MT1a5JAiYhwebE0UPwZiKxOvJcbo+6YgkQlcpj8Zmycw9Q9h0Se6Ny
Bjrfx8hf5jmi9Kn+lQxSco5tS9SIfNYb0CX2l/hOL+SFFM/tzZHYZgvJzZtM5YU+
SF8OfhdJz5dX/XkjTuwjhjbYkL/vF9bBiKNYXDqAeEeUA99U6XiURvIaxrV8o71Y
XwNG/vbeNHgrFIPTlHxR1MdcA/wKcANLKq6JoeHqU26IF7Ohpa0Tjbf6s/1GyqeJ
qS5hLBW1V1kwm81FYVsooYC923+2YG+/vM04lqO/H/fF6ENvdmT//6goRwCI1FPR
KZ7CD/US9XHYoDuRAGyf4l7N6FfyTuvlu/rotUMIVY4DF+At9ZkdySCzY3H7i6nN
Lf4zAsiAum/1k/8bT1RwiHHjr6kM/cuxAFOdMXjr8iuP8I4pyqwTcmMpPcSTM/sH
LzIKl4tnyut0VtbrHTXJ7Kwi1TZfMycAocZbaP5Ug8w0EPM8nwwcZDOkww9aWmOP
RidotPvPkHpRlOZufdby7mXPJdxZPFcs4RhvdMYQVGWeDKrcb6F+gXGtAQixDgiV
WO+znzDGQCiiyRDOtyvNicYyAQgJ4+BZCpuTiwjVf0i/cKCruXTQKsV1XmZ4IwbZ
/BTd+s1TnVHWKbM3BXAWq+/bftN3LrUG84DDasE6WwQlnp8QObcsD87SlzjAIIgY
r4MQujkZ1Xtk8JTutVym238qz/rtOGjlsOY/b3YpJKBcVQusnxa0weOfCC5hOpz3
+POvbphs4eZxr+Fo+75vt1EIKiKl5mTeO/7/WMk1angJ4X9YnyBsCcOoYu55eNDb
l8NMUNVm06O6EQEp2cmqzylWWWmqGIeEuYPe3awKMqX1B9+zCg2lA7d0BrURwJs7
UyzCd9XURfc/TdM9a3295sH6+jxczJzCCflzFBAIubJlZ/meczgwV+6L/UWyjxLL
ENxBKtK/TddWQ7vxzdfb5qJpg62/zYz9VtyyFhIqueZKBbxWXSGSh4OsEgP+bkJ7
u+2cH030VpWzzS2OW3E7HGMmOtAGHBFQ5sxnjjEfHPd2jlLyU94ZAsCeT1oM9Doo
Kewm16opl2UsNBZ+1s+QyuGOS0Z1fKwNpDZeabBlEhejWA9TmBrM2Lsif1QDF4Fs
7kQtLibcEj4YEdVeKEqJU/S8XivQcmzM0SXQOgmGR5A9gIFBpWA8JJ0twfZ9qyGZ
7hXNPldt3kYzpliFvtPTrxiiCJxLnB1hlJ31EX8mg2MqY8jzD0TC/s2VWYJoUH9x
v+HY7prqX9H9ZDTtwhrGa8jSzq4pViZigatVZQgZp00/Tl62ftI3ZAb/GUeCy5s5
T1nd/6qsyVPWuQi5+KcbsHOqO96bKUlNisW/ej4QQGptMMPO+/QTs9yk1el7w2yZ
XJ7MNiJZTTCsCbKN5BD8wGBM5dId70W9aQbgGUeYumhAk5EdB1cqX7pQRVN5+TJ1
Vty+Om3wI8ny1pdRZiZ2bZKb9HjcJa85HaNW01GkWQCCWkFASghONJeF6FKGtGt5
8r00Xv8We07eys6vsM8fY5JDLtB2bMHuLE728BXaw1u/lv8SSdmty0v8MOV0ay/Z
lHTg5X1nRYZoNPYryRg1ctOotc/SGAwGjdoVSnu9Gxu69MjSsF0IHa9FLcM7EnNT
Udo/KomVBY0VORj9Ly0I9ZSbJLmidSMx9SzX8fpmhNWMA7KKnUjyFeXRHoUA2vKS
2wrAG0ji/05EXMv612mAkGEq7L+729rOpuV3x86kJO7ko3h0wEn2S0m9hliH9IxX
vE9taHd+rzhi8gGLqQcueGp1nISSOfdKGVZtZmXryuUxI88Kb38D68yzgJofd08B
oBm/wcSMR0CEEfqpI3tae58Hn/QczIHb04WfNEZsztqCmKvbU5gdOblm2Zqmqdvi
w44j7Qtj64rlFZ26dOiWBKcopPprqL+kfCjqrMR22aMHehMui/7Cc6BQSrH9/15C
2Zhl/phsKyovwRiDUz0ZB11aO+nf6c0+Q6+fPxPsBWKafFz6erMVLaady/ruzszZ
xHtIo3/GDjix/MBtlcTPkBUT2RKExZ3LIrd2SnaWd+Du184x5evHEhY93qBmwqz8
5ge3TAuZyHCAu7egqlgxIlhOfOgKP5KDsU1PCt8jb3k1MqN674EOTEoTsNRfVp2Q
BNQczhIjkaEWSbhPfXgmjIqRElusQBS8rELQS3oODZdvzulAFXpi4A+Vl7uuD/GW
wugoATjEhVxj1yPJW0rGEX3quzuwCwJOr6GOGdXjpemdzeQOku2YJpLR1L45/bMI
ud6pzMQCH7MkJQ5jGt5HXKQWxNlaDAQvNuLMslwq+xT+ulDiX74AGCftEYriCDxq
YNstIVf36vQnX6cSREbgkFUPdhIgSUBERlTkSSiXJ8TgOPXN8dsArIb02aCs05QG
lGEYkl87e1vIYGf4PMz6B79Mc48bXT2XR4LopOH7gQFP+L+1KGi7cQOXKBB+8fFi
k5/0jpZ7nAReJVcG3oO5Q2SdSMCXA4cxQcfL/PNBexNMxD1jyQRoeVlrHz8qPO5r
oELbTNRIYZOffWtOpzchfxTy1Bfc0p2NQdcLUlUvuag+ykMpPJFvPB/AsvXItweB
UKMRfzguD0ZZ0e9k1U5b6YZSY+X1yyhrq/FhcOJxbZfwQg6CoLdsE7B/6+LvqIJq
wij+fwRQzUZ9dNzQamSVyUlBrL6H13Ig9uH1nG5wJTu8a0MBemqgFz5MgEu+ONMJ
cZd8B529xcTk71t/xKuJn5Y6qTJTTB2PKZzqyBi0pqXR0OZYa9cvGUyZPfwOrIly
Vy198aVk2FB4NDddwnuKwxk99MkEi2uWcAyBlFtM0UDRp5IjezmvZfHDJutltNPy
3A9qz7cRaCOrYKenlKDWPaLnFvMvAptKTkJnJWIiRnoez/6T4vWESkZ5XsNuWMdH
5pFlylce210AbOPf5sxeMOpy/WzkNdKAVlV3HK81XLhe9PPX608N0Q3MMiRzJm1G
vDiLFehjB18eSBLCAOiR2YuJley5vy72tCNnTn6fbIQdS/pFCbTcZxf/pb2EnEvv
yVomzx1+dXxHpeltBhFhr38pteFY0PTQhQAEZQNPxUzPNv/dp94v772fsycrSjH+
iLelZdsHk45+rxwpAwjQHszz0gVkXxGY27TK2sr3HWWiSTuxrKUkRjAKQZCd5i/c
+O+RqJWk6C4ct19j4+e4z6uPMcZ/V+sGqbKze0XPYQVPQJXUVmfZnBlEetBSogBB
Vep8mS7Bm6c8f/SWuWX7CsStWC49lk9oN7CFE72O65LrAA+/fjuSAM6EGtm/z0UA
hOnwKhNXEotgmEeUb+C3HHYjsw7E3ah9h7RonEH5UoNGLzvxd9gmEhD88qLQebOa
ym9UhQonD3SZ90rCVE6Y0Z/dXplmKurmTVZfzHDAftk90ERN7x/jNdZytBiViZDB
2pXmfQHCj86u/VwOPuPXN6FuOr3ni7BRggqxRUOXpxYmkARbKYqRW4ZKKEpz3Avc
Vtie/BuYji8NCcOeQlk1/wWN32eCKzgjtRtJqRi14l/NiIMv+/3fPSD9j0qz/Nwf
k/8x5cI4CmgfC7ImP0kjHavD6Vle2L2xEmGpI7kmYmsyb2RtpaGYO6ysf5hTmxdo
D9TVWtUdIEFGQ5FJnwI7+FSA5CL2zyCsSAPNWFa+AcCtm+fkgdF4duUkWQVbf3Pi
mmPyaMLrkQ4881fo7mkWIdaShOvXaGntr2i0EwVxpEbw9QTWOQrinZq9+zAEDALg
fy7vQaUVeCw08YJLpjVGf2T48oSdOFe6RbN0T1SxGEuhZQEAqg8I8pRxWfmCQgH1
w+e+pJ+QtEPUwwjKGLj6jHjhk3Tyf7bw8b2GMmURrugl5Jyxm3YzS+DG1QOA1gxy
jLwE2hhe8Say0W+sVlcYsr28o35H0VpDQUIDtgwwa1GYqFrBdHBMXwOcPi9f2eZk
h8LChSqTntULpbGwqAPsPhkZp2MHycgJNwXG3XKs5/tHKDuF1GOcWONuJLBgadNe
jhqFBwilpz3lHhIVyRYBh0aqemC0RC9RGmgMfep26bQNyxl5mLMSCblHEeqqw3ZH
vocC6TjGqUu7Vz24FjOm2x8cbzCicEpwRuAoq8qHvgGZxjl/SDQKfHFTic9XGXOB
W8sJYLFsqBy9Xp/2PXDfhXerobQ5VhpG6HEQs5IQDFqUzw1PeSYqcqLYH6ZkFWW4
ackiQyaBdmCmA5Ha3ng6Y0ogs5cXQnMkksf0RfEeKefr6x+PG5gPtJoZayqInRFP
1i/6o2RCqVWTDPPObqWuRvKhCG+Yw7UX2ThcAkBk5qgDZbIm6RK0LMmwr0L7zoXQ
WiNFWq8jPDq2uGYEV3Y35QAJBjfL8TNOqC4bgridq6TbD8HfWPjYnLmXfzFlKyUb
/vSkpQ7aPmFEJrB93fsIRl1I/ksLUuVSkKCu2rrwKzC90ukY7Inj9+z5Lcbjs+Vd
fqpsLTrKmFYtdnxupEHVxalulHbCpPzjaUaxZ1smB3bqrBBMo8hJ0ekd7gN1RIjW
AM2tY2YZN9R3V+B14+ZgYQFrDOGnze5n9JPuBn+ewLXX2vqKMfotPLHC5aGZJz3W
yncZRiZjvWd60G23Q8p5xM2f5/rN/DYlqZfiBClslLJ9+W6DWviVT+UKXjlYhF30
fz2ofkXM5UkClhtg4x4J6uXwjl2pyxykaQUMbLz69zMnymajYODoVrqtdYqxeJ1s
8rd9r0gDqCWNm3aNXBbk3idt6InR0CGu6+9gP/LNLZvqLHOjJgDeXljU0dn8jziY
Tmj5ZpdmkcEGqxtDVeRaYVhQNuu29+f7PqnzfVDs0PhJn6X9+0rvfHKg7LX+vA0w
C7/T/7zEGqmrYE5dF+vr6yUCokYmuFN5oRtQn/MFh7Q75+CqYK9+sVIQGznwlLib
iqLZmCpWglL6dK2+JccZrlQsWy2VOffvKVY7bUEpLV+Pbb7GcOwfBNselVMmn8VT
qRbGe2TkL/Ip0EtxYYWyY0i7F0Iw2hQFKX+1WlMtlurJKdThy+Z80w80jc0VpsCc
VkM1sgaMe7iLTSJ1rTOqoYNyTPARzDL0rK7CFytnxHbne1YIwzp/tXsOomtqFkFc
Sow0Vp7bfvowNDYDqL+JNkvYXCAtU89iXq5XyohfdoingzA8p3sbxaqz3wzjfhMt
iSy6e7ayhkQhOckanGBDMENVRFhu1cbw7EAG1aolVEDEsj6UIXGUua6bvroinf8G
zMoFcWEdsZM+a7RUh1ke2n/+re0u4j7B9GLggJoA2QZzTZ+zrW0O0c36GvzRBgkl
ibkSdz3VoiE9Rjmjd11a9v+DZ2BJmmr/1PbCzI9i6fIthTdpj657El0niKiVYLjV
ChdshPD5jz5WRTQa51TqBBKCEkxiYhi2IMm1wM+XK0+oKj7nMbyViYkliX8NVyOS
ozoYzZRqt1GhVisNvVjgxE/JgqYjRlFKoDgZo3aD4KnE1cc/ELSmHjZrNw8OoqdB
LRVgDrI6161kgHE2v8h9w8OqVXqF4FZpw3sLCaLJyxkw/6fF1y/BYEzmdzDoS0NB
0uMHwMzis8OxMkDVPsKM3Tim5NXRcPuPt1tO7IuVk1uicwzpXHjW8SXYVHzd3VNw
54UxRvQImErBheDE2kpaHn8HtXSEzRWyJZCx5l65iNfWl3Jz8FJ4jDVDoM2u/AYr
o4V69+cro/qgLg/DXOcWTVdCTAHK+kYNmb8PiRSs6FhWLtSuCVcvowcDngW8h/YB
J8AYK/vimy+cB7p8gYTmTbbFuyW8VE9FOx/BZy4aCeUofR5Sa17c/0ecnX62T1PZ
Ghub0HbOkk26EAW1z1zNYeyuPYOl0LmYFOo8to/hK2czbVJO0qsoIzulsqgPiRGh
L4u6gOgWllz+/3vN7o9rCoK5jFgcPlMsKQKTAZCSSZ/FGjNMvFAUKvIBtYhD7HAq
spzrhYO20LS+vuPmWkT9u7TZmeBKeXL4QlDLlyjmafFvrTVqVtxoVIlBg3vyTNJ8
oCAQvUJjAZXPozlC2SYZFekQOW7HNaIQx9HcjcSBKgGW+b9X3qMyAQHU4kSCo1sZ
xorRJq5XOH1vICb0HAII0h02kkpXwgrbJgVKnlisQBz5P6ax4f4bbwR1aY9SJDRF
KaaGLU0UzBWcgpHeD1NRV3GAeZm31GsaS2Y2nArWPH0aWpDnlnIw3JiRgoBMZss0
B109+Ql1NlL/Ue98y2+kiQSrCAC6kAkkA6LfDw/MTqtvCf6FJwkDiOP9aKzdiUq0
8gx+sZy92z4b1shLwqNIYLWmR7RlI661RgdurZaeu/RSZ4a8a9nOz43IOIfXkWY6
V39qQ+0Nv3+wD2g0OdD7G/jVg4A1AgWbWmPWSkUhoi72aJuGYKHM3QLu1KZ0ZoQ1
vROdr2ifysU6pf5TN5Hd0rL+15lF9wU+Din59bcifKYT7CzdHegNX3rCaxTo2U3x
O+tOymQJg8jIUGNQgs81nFidY5QQ/raGlbTU49j9DrtL9CXcgkLqg8IeKlWcvsoN
Bm0zkyoYkp5XPYLA57hl6yKdF2IhR83g8DdX4X9JKIyRoBvZnxw5Dpgm/Rx+vEQl
GpN9mHoGwWdSwKRA+JG5GOGMgEc2WkD2P91NbinHhk89XcBcdcSU/vljAFe16aK0
OiKCF9vSXbzu5Gwm8A14xhA2xLWzxn7wiTF69gt0YFx5Nur+9PsET6xES8Tm29u3
MkI61gVbckui2kmWbK28135E7TrmkBYstzpCJIcuk94pu5fqG1s2gh7mOBTvrIsi
Bexyu/QtUyNjtQHt86TXfI4ExlctzoBO+PAMai1ShL6kAidGGwVq1TPsNtZ7YEdx
Qgh/yjwg42SReetf2l8fO58UkkTASin77TyZbt9tMl2f0xWQiPpnM7wlb56fQr5L
zU3jIFGzDw6LAtp2PpKhaWNnpvZHKIovHs3XRv8MoOAKPnAB1h85wKSpfcgtdH45
+2Qe2g+h2sq3lzfmVIzgihOJmfRdnbRE9kNWR2V2kSzKKISANsY7nrI8s/t3gLfS
UrPDJW3jF2E73krn3xJwoPt83ItcH10BKOBiC1tBhAJhJTep10csS6llAhKBDMGj
KVUUGEwhnyDU8Wf5O1XNpz7tqtvLemGrd5uldkp/YZkzoM+0Y3g+UF88tw3nahgu
vTnXOCuYQkcykvb2L2Bo03F0hdyxd3wyI+WIFfMAfzLGXm34zLRf/6HUTBDU709S
QircDbS0wLFMx2F6br//vjIlNa9S3r8i97Rc1/qm29aJ2UfPJdVezgsWa7ayBCv8
eV45IQssZfzPlNBPcjFq0zhmUWtEjlmzhCnedcSjJzEh2QCU0pI9qRBLVkRm0OFz
tlP+3ViG0tRkSqWVIQy09Ndq79Jkc8NOSZTrNRGQvHNeuseS7AYSvFj+DIosSJtH
UwoWgB8UuLuw5dcF4Z8Zkzg4LiOliqXLmMdZcgACXwXBR/HK7RpLqMt7vBPKuwhu
YqrdeS7I2lgTxlDM4Ptb7Rh/ySYt2f9o5yiZbEWqs5pPCF5BVZR3849GVwaNCMFU
0C36IlgQiroCMPjtq6gqxEAOtc+4LBuBYnCLuWQcie2M/tqYBDzSXIGWoo4WsML9
xYkvA5ffiyqwF8V5EvZakfl175WKoHfcwZWfaObGdURBj23aM4W6N4MEq8+a/AyY
6bce9r6uleUwVvgPvP8zpc8hpiA0K8e4QT9HvKIkig0nz/U4zuqd+wcGbaZNt7K6
YflKRp6Nv9XhtAbZFRPDqZgPWPxa9NAgmqpWYrPRX/7Eq1cSnZE7ZdNLz/Z7bk34
E5hhrB+c40aigyIffimYItZeT2ZnAWBkWLGmcF2NsyL0Cfn3sNc5pIsi2rOUiCni
0g5dO44PWUDf30xJOym56FLNe06psr/UKz8x2Q5aVxrH1I2zyr10meFztJCLKfLH
J4Sw6LFQQPsXHtQ/XZag2hFOVS3CWA8bGdygX4FXmUPlXUn1heRRv8Gzg4on794G
bEfrAzRy5mEJ+tzLFEO8k+2jV0hndy5TS+oFL8eNpsZqkj9cMkCVqgE71iexyfIm
ifqzk3rFG31X107cgFkxa2aJNKqS4h4O3UOfrM1UIDGuhGIAQTxI8jf3quuINYdS
+znDuLTuwxjfjYTM3Er6o1HHGdST0EUWE/av2uzflgqrlp7tZoTmXSpDzja27B0U
RPIjslEM7XzMQ+1Mc7DTOY/TTHelKwlYrZrrsR/YqKJH8h+RP9zjDJ/vDxYQPn1n
VKQTL0d8kl2I6MNUS46zCWAqSnqWEdo5jzwN1WKWM4rMEeGBprF42dc/p4v/oR77
4K5lvLqLtPivFys7cA/G8N9XF5sNU7KgOWVaeuDOk4I7AGLcR4e2xkB+aUpVL26q
9DVho0Z7hU3ov9zFuDOPbaz8dIOThyrBNSwswLdQs60oz9Wlel/KWq8lenRId+ta
I6yUJBFq6V25duSw3TRtTKL64jOES9py0n95cenBLfByk2Ae/jhlbykDxIvWObWx
fwqiuYSu+JTW1htU3HNgwTWgYlI1PSLcEowf6T+A6Z/4FkQzyYZBlYYp2ftJfRr0
AbEdVOS0Ro2/Uj6evrxy8OjWU/XH5VYbE0lnnyUtWE3OatvWmIgDf0NF/SzYqYcq
akzsb9RKvBI/5RT48FtxSwBkobiM4VU6wIEZH00buw+bwpKv/HS3i1CyIQw5NbVt
bdYPe34jESbkNAusalH+AEC+QnVfNtxzZf5p9UcO7febUL3gsb9GWpP8Y3mMaXuS
jxWo6LHSPQE0ZW8ECcxhP36LUMY57b46eGGXE6gDXxS1TJa86lsf43tmLz6bBwMH
137ANwVwd9RPbE6Vo6eV4V0Uqv9V9KDT1mk7qBLOxrGMyvxf6ctK1hTgRpQ5vahH
h7f6SQSAcpTwdiGEJFybm4Gbhxau/f2RYQ8xcNhf1hZ73Cl6y/qT6MbzvSVC93ME
c757TJR8d1HwRIb9yMxKT3JayQKxzDoOhPb7zNH2mUzTUG9v3e734q5euX0r28mW
0SfOT+zoTcCZdkfit0ReEHWge6Gk7mZM1FnWW2VyntFDKte4Yfmu8QUWOXgGVmGL
+aBx0h9PJPMOevJ0cOWRnQnRlEAZvtxTEJha5pxjfS06lN6IdEGl+JJ/6ddr5V5L
o2p2oWsCvj2SQezbNjyafoDg2YSbHFBJqTDQBCr53/sMilM/Ry4RNUoAkgCanDAI
EfoqjauqaYdsoZdoaOaI49Uy0O4xIsU+fEMFwUKH99q1D3y/zTZx7A18a6J6mHsR
PVNwwLsqCsM+B9BQjdOWucS3517UVo22AJHcDUEGMNCdoChKX4mynV+TwlaqybKd
44pDnRb/g/L2GcnIE8DY69ysALGp1gHvsYU2xmsufpRCrlxB61qtnafw31OeNNJz
YLBp05jZmkCwuWOe7smTDWEbGUJgZF1lJaSwcHMGyUvxwelqoUo4Mtwyb0N5Ucj+
6S95j0pJ/QXlK0SdYHb6oC+8efCDGU4VfduDkjBk2TpOtauzGAh9592XCy3K/58n
bnxT4XRRNF2o++D5qiUTYPyhqRU8sbvPpTvyFWbMqtK9+U44NGigAGgiEA7EX+nd
7VOZuwXcmC7Cn5OyIwWY55JDmLEskmWrPke277rCTMFMQVhgGJzOUe98z1sDvump
nOOJvhfjHmAd5Vfnqudoy3i1KIvW6UWXWZaZTHXAUZUoQvFBWCSIEaLI1mPmr+sB
RqmIhqaEXo0MYo88r+St85aXaOTap0g04fRVargcCtxeo/7Xqp9YU319GivQLkuV
8S8GtmCcyiXueIh9QrzKknm0vlxHo34YrorJLQs7rjdXazVcmYKujV60oHMiFZv4
LbnNEr+YFXuuMZqD2xd9wU9pbQveWp/UOiWCDrDGV+jhb/3NpiyYNRg7Ql4LDfWR
vsx9GP6GlWjdojDQoqXysPTiS8J9gVTWsHFhMmCLM/ySpDwhjZnlbhyjXzfWH/tG
AmspR3pPuxM/pRsbPehH/Q8l+nPgTPtvoh33tOREX9NaDEi3c4fJdAb8ivA8ZfcH
5Y0rRCh45+L79CZ7/62CqANc6iXdv9PfS39O+7VgeCE+yeAfHK6G0ute1l95l3vH
EGkoaRqQ6T+7ZHyaKusfiZkcfU4qsJLmPX8Q4hufaUNNnz9nvs0daszl1KETLrTM
iQuVEF29P5/d/DcC2TC2ZPbWX7dUJ3i7qZggvxGOSV442Ilypf0tB1Ew42B+JiTi
n74bi8DtVGDmI8/DqCwfAX4aOwJWf/1y3hbhvjZ370KFTNr+mhSlmrhOn29qRG0q
YhiTB0WcBKqBaXhxa9LwSE7gpdTyVJIdP+rOYGKa9X0MR2HzzVL0q8xXSi+eART7
VvaeIz+MfK4T75Rj1OY6ByveEUERgmE5zIqjsZgQTJrUlTz6JLDxxjm1QUS/Rnzp
pYUeLi9xXWie0NvyrZX5HVKq+olnQpjD1Ol6e0+7yYqWFdIHBbHnuuP3Q4+0ZfKY
fdTOi3e+pSMhIWM/oI5HmokawNibsz79LXVz40np+8ktuX3iqJfDMb4KwAj/Re3o
r3Fy00JhrUv977wbd2U50RkncIQIbWH+Ms0gLR5xF4YS61Z4svFTVX/c5rErTg3p
8tIVexiQR8Ti2mLDOzf2NSd1b/tJSpjJ2szBhIOnZxd04aQFp4ARRYOXIiGHqt5S
rBEqRs+g7Q4lHZpWBKqD8fRS5s3JADQgMpiJZ780m0Q3XpyE7tICiIfWu8C8JZR9
tVRY9+PhuC20ohaTd25t0VXTH1iy7LDB1ZI6GQm7X6kE0FfrDzk5J48UuJqgV4/W
29ubwggpGwiu82PVKuN9wTc504ALpLED2iExe9t08RS2kRLP5qIaUG+IAodkBGl9
GgMtr5a2/eTAqps+T5K2yQSzJ8M1cnPOkXfTDi0EsR8odl59XpZTJyJF4/sRLzOs
N2WFRMoVovMI6NBRj/lwUS+TpG48cEk/c+ShCYpwZ86jRa4auIoI4tTqC3U+i+9g
MT9jzEhDvq9I+79H+bB+BLNaaNMl542BhCNAsMrWLOgveIk3kVf3n6oRNLaGxNxi
/zP+jU1tyAp14OrjSufTgVG3baiZhMCcYSJ3vpr9NebGOLI7rFMUmPiULYiVMJFL
R707dtf7nOl86h2vfJp0+yjSVEPV+fNYUBs1iEt5CCruslR3nmaXDefEzK7iqPWO
Xzjea0N41+nV9fuU0vv/u4u3nTqM0WAYSijMNSFB9dy2YpnDxDbQdYA9jC7mCz+/
4n5XZr9pVxp3g4SEOcRDQQrdKm2inKUzst96Mw/7SUIZSrzsRKBFSil0s4TQXfAl
LMVIM4l0M4cVkLapHJUk8Y2q6mbw+q8K5HmwXOeeupBJ01nSCr3gaLzCPwJx8/oY
q5uvru/W6318KDJ1vQFw/jApTlPflpsMHUPbe3ibTDAmonfmzAByPgkqPPE+ufW6
EsCu6eaIbhWO5ZbR0eAb8pZBoy/buDX4TbzR4DPum7kKaeAmSnqAHztOCc00+R21
9ED7bUzOeGL4xq0zebdobWwA2MgimxaWRWrm4PnTveJLB2axAKu2fdq3q5C1wn3K
MdA2BvWXvuu8g6zXHERvPdXjexSseNXDQTSMLT0dzXnHkilKyqSlrrpjOcQ9tQOm
4oi9+KIXxFtf9hbBTFjgAXAD6ed3P2j/Np44TdGuk4J3Vp61rKPGWC32UE12PPuU
6KAnOVNL4L6nUCEN6iJzj/mkvayNpn2i3l4o4bjxmt0axUCoxQHcZ/P1gebCkMH1
TmuOSBbn3/I7Qru1XPQOMtcnFrQ/VfJ/gFW92IN/hvht76zjRK1SSta3xrho3wry
B2tZR/Pm0jI7MtXNDIPxW81H/9+R9/eCY4GZ4cGt1zus7e1Qyvnv8S7Rh+xATXen
V6Z/Sdzqif+Mn6RhTQnpP8xqPodD1ByJEk73kznADsmnSzwyvMWO0RN82jfs5yKD
oLl2bw8T55zZLTy75Lv8GXPpN4P0bmwhoNA3Kuflyq2UPVe2Mk6KemUJKImo52LG
Ivqq9HSFBXkj9qqf5ZcANcSW3bD2CgipVncI/oSxLld7Rp4N2LFtACDFSeVUF4iT
zsrazP4rExqj/CyhX0NI7N1VB/16anw/djmUYJlahG7Uh60AGPVt/rWWoFVsmkSy
Pz8R/JCzN5dkGe8XFvbNqa4bh/pts2ww/CG426LcBDQm5tWGqsFGC3WZ18dCU9tA
Zn/tGG8sE3oM0lxBgaVOPzDHPZitMoI303BEoNDjHg+zxT9iYNkqSdBKvWHTpQ3A
2ju3ohg8mTe9jXet/B5D/ep/IIlQRju0gDiPhvIapcIP9IfWj/KjE+dZT6IFMN+a
Ov1z6PBRoIj4KPZpMOGo6a0/38NMhGk8pRM/xpWlH0iwXLrRejPJWrLPXm8pZSeC
f6uksAqnjlwClOebiKvf2dlWZm8r8NPfaFoVF+5fZUsxHpNkDNbwvLPcyUzMO2zD
sL416a99k3Ld7eSPWE2vTSGs3pOTexL7OmdzDW7BK2rKd6Cz6oDqnH+n2mJ7QSH9
c5oSeACc1jeYTtQ6TTW1/iiRul2nbMrLsaJ4TeXrk8ubIxqJhLKyWyD8lpYzbf7i
sCfV7KAqFxoPsaR3RBGj/fiurkWaKpb2dNEJtY6OhkaVEMo6GBTDAUAKwStjA7fv
3AxMil6vwIrND32LEOO9WM3uMzhdLVfpXNQX7L9J0Usl6TWZF3KqAhx5UfmJvfLe
0lPtqRc1FaESPGs0OdEb1IdbcOiSThTT4SNLln97nB75Wwyp1SiJNaBR4u10++UK
qiChFGp15qZ2gj01eV5Yp0lmRkGqWNA33YUFv2N3SPrstpFq0w8bMuW39AzdNgFV
/OQBGLhjnqTlepjm3DeMb57EEWT1/p5w9Tp42Ts+8iVsHjcBDyxEUNeF56BaWbIe
DLJN3DihBqud+mPMzB6AffU5Wy5CcrrqjJQoC8yBD5ESCoo5jxEmgnjIyWuXgi8W
Avk8XpOT5xurTEm1BbEG6tsu5yXIvfkFy/HE6NeOKquFH5yUZN04N0757x9EfTMV
i0JXAgII2p4WJXfa06xEaTcmUwqycZfATubwY4sUjbg0C+Hw7FjfkHNM3gUefYUQ
tAKu7RyAL0qUvQwZqtxnbWm9diJGGVxJG7c56YYUvsNoD85DKEZG9lSS9hM482Gq
mRcc1ynO+FiqtWEPfAIxR4xT5OO3Q6woDlWlUHpZt8n0fZmjsnoZtgJBgmb1ZW8o
3yWis08CZOw8PRjLesBJ1C7ivmwGNTs7jA1fCgxY18rH+se3MbimI8OYSHzYN8o1
lmZxsgWERsWddjDnfZZZSFW9jYSLAi3/C25XnR/etMhm1T1NuFMmicfspDLkqeOI
1CHaV/mpP6+v3xLs5CEMLE3WrMGnsp5SY9pqLPwqJOWghskDeNDhTTCARQWs0CXm
sjdRheX3w7fcx+IYZzUWTWWeyniuON/h7uhSu4AfjFHrBDfcYbPYRo8AGu+8TYGN
blfGvD6EcJt3kZMdWzmAXrWFww0ewZxuza4jpiaIV4IBCuJOyVg8oLWBkn0+B3Nf
YNOq8y0g24/3vUKnUJiT6PE0ZBZln/VG5Si0TXn2Jw5nifn7NF4j8mt9gG5TFFby
cpgON5C1OBS/JHkM0nfjydNYaKeVU0t/fFhlnsr0GAycodUe8egfF/6Bzu2V5d47
8f5iG2HcB/HakywcNHfWmr13Nstf539cGtxQlpd6TTiXeg8clbSvEn+xcMiX9IQr
68mE6zhXZNCWXeby2NAMAC3jltH2HQZh4D4fCZjkEW6tndKVi6KNudqj1M/TY/iN
B32nxy+sHI+S/0J9ITh3lhWePParSZSnV9fQWgY/oFFnc5WYHyFEDuGE5TJjC9Vd
jqkbPDUl06Ovl59ofOoLtWa03/QcAgWeVm5LMWOJRepODGUKZ+CTHPV7CYE9Ac3B
Yz1A1PsOuontbKckeK+xZ2ekugztEGEINTObFbAWwD0OPmjyCoxO/+jGKoV55mVK
QzMzAvbFAH3PoU18TLKeFO2IqI3z4gJPJfj4j9cnRvT9nhxc3G3+B/ZRc1GT383c
44kS+YVClMuXvSSjRKrB1Xc5nnJqr3KKf/MtPbS3OXfCvE5DcPNMFGP3ioQpGDrn
s3Z3clgWrodqyLNcMFjpvw0u5GlPX3ybM4zx9ldGIaaHJ7ipedcL38aN7LuAKlS1
4CNDfSY6Wyk2IMMba8L8/uNUDqCa7OzE11KM0cezpvucq3GylDGIgQrB0YJwQARW
fYdT4mkdcMlLZr9iaK74XQVZGPLBdsTgznSbrrBY3ndvsMTFSw5dCx2H1T50qewo
OFZrHeJhBbiCp74ci864gKHh2107w+Yjf2IXBzBtI/bwPITSMyMCftlChx8JdIPj
hBy0x/k6EU9V4umu2Uv/ivaC5p6cb93XfFv1GIgeOhJRm8AAVGoMs/JxYAEsEhCh
OJwFPeu1i8zzRNDxNT9xVi7kIBoSHnfuWt3z7nMf9AsQNxCFca+0/PwQvkr2B5Mb
VIBr5fRl1W7W2+pLOaukgxCgPpjn4cVOQ3wLHBMcwt2Z9rY3y6Efkz0WqEwraRuZ
NcQU9NQ6st8lFkBIrO5vgYvQhfjxKoPLNEWpP5v5rRGH259JMYvwpEBuhpS5OhWE
VSSn7DxxheAuBIcroaZ3AAHUiF0LE+UqU+xPMp34NH+UxZAkvRz8asmebRvZmdOk
boEfEWHGbHYFmntM8MSpO1By7iXr3rp24Po4dr4UrTH7wS+w3xLf86y7Xtlpf3Qm
yJhqPYEDqK8uOBiZCVF1F88UCiKuKUoNAnQIGRY3vlE27cMUqpNT9xbn8Mww7qs9
gjS9/yJUiQq7NMuBkKAKKIjxD7og28gpbN0V8t7wevjMb2FZXQwIG/n4Yaxj+0Fx
rK7N0EWqvangQ6FGyxzmPVB5jENKEfmvOBc0YRxyv840c9CA1VGuqejtqNvo5arX
WJBY3GDn988ivnr7ZvmaqvOLSCzLc2Ha9eVO+HmRWuYkThM66jhiXL1JkteJlULA
ECKS3jwjMSqcUelcgIdbM/GowTPLOi49S2shnZ+F5HSQXJUwpJeEXrdOVP3gKrUA
PeUnSzpZMHPC1t5u7L8b0EeHVMDMW3P8R9P9Hf6Lvm4lNv3X3DAdfVnj+72UCj4Y
2/Np5AilNqqptljPX+YWbN6Fy/+Yq7oUBYy7T645nu86c534+ng/+mKk59CbIax3
UpxOL/h3/3ec1lmXzZtYBTrRu01xrQvKSN4wvqQTmAht3TlGIE/p7/jhrQOs3gz5
Csx9pZzqs9o14wGtfZ0ApItLteDK+9OY1LLSC7orw2v5fquv14QV3t3MYZoHsx4w
By9fvCjEtZlaCYc5J4XdRzG5FQTN+U+SYtS8fhhPxqc26jn4FAmZZypPfiQKGne6
CGdAGSvTowYxlpEjuFF6GJVfeSSkd+se4NTGqbAoVEFKEqvg/t7Lo9AciwIHbsFb
tvY+yUMWRV55/zwkMkXEsbQwPw68y1yl+ile1kLQHLUSwArP0lFI+6RMhJBcvkxH
QWyGI8cHBvndThZVUgBwuyDbwigeLHIpvB74hiLvggM37023NjcuT9JGlf7BO1zP
tx19gqItMpyZe0wUYY4kQKTgKG1+fShipslSOqXq5qhHk/H+HZ12B0VjmAnlJBOM
9epOXXKaDH3UswTMZVBIuNuJJnRI5jbJpV1KM8fL5dDalQ84rGQw+AgXEceqT2u3
RS+PnrAuEt4b2z8ItITV3d+u67AgNYviNIf/5WzTTAR4jpFwU4utSOLOsZ9REU80
RSrdYYV2S4Qz3NCvJfzeIdA5W3rvr5Pv+O650cZpqYwCFe9vWUZNgpJxIiZoldry
chO3ADr80MumN90HVVQduVjZCWttxByTCx4MKV/Mxp+peJGv7BLVpi2I/hZ1/mCh
3C01rRCczWrYM/ATssw23V3tK8PXKGEsR/5Lokt/dyGiB5SEe/Md8cENAZXiHlDf
1+Yjikc+QY0moKNH8NXBSvS52VpbTzEvmzNt2u66qiWftLQ70S3lgysTPuAlU318
gumRyK7qyDvsxO/TYzd1MGgIEfuhccP1MKiEFwUWX8vKSyvHHukN8+4c/YKHIBgT
PiEZsuC4rCXASH9l585KzZpWrMF8pj6WqfT4ahkbGZLDWx3U+WxL8E0GmAVIfxBq
WykNa7KLQ9UqvekpiexVRmBlxe+7tXW3eKPDHMi+7+HqXf5waFLiPeDrKFNVcu8p
nnQ+QWxXUtg37YQZj7OQT6OsWCjZKjmFk6QllvNtxDm1iB7GFug30LesaA0inOWZ
vC2SaToPAi64K0NQhWMgvNWeZU2Sc5DH5crWxz5klHquDCm6nZTac8XRFN/j1a9B
gdV6iGeRP9/nef4nGPpgJWmWcyZgLCkBP+zR0DB5q9IH/gr8Ajl4BdBeFXcwkmfq
42ElZ3RXukVh1HBDZOuZzDzf2OI4+Qk9KvpFu54tjxtnEB3l/YMjyccU/vFqsYEL
YioTjUftcvakieFn0rDKWaAWtXOwglp9yDj5vfoeulApqVEiw1dwIWrPKACDYfU/
1rFdk5k5aPgR4net0fLTA+4bC8quiiyOkx5ytNZoPpzkklIINgoKhRxT273/JftL
6aenSXNzd1p7hF9GxX7bjNo7UdXMfsIJAwtq9bBFgf4gN5IUTKKLsOD9Jd2LLdLA
Kt8j7xQkbkBVbPfiWPwMliWsjjD6saJF4yA756jRRbz9q5Ha+eDrcOcnAs0cRUQF
aTVr70HbL2ydEQXDEtsGHvDvte1BhaH5Xo3knoH3WJHtxIjohSrBHIJGUzRzVagO
yVoScBLIScIPhsOUPJzm5F8mOzFDcdsqd8Uh/GuQFeArrG16mD3mXtEiWewAef1D
Luk8gnvOwk7wfIsQcXuFheKyFUJc5qPD2N2URTyksHkdd+yuRPTekCpyQ5k0weKx
EfSo+XIlUO7vu4XcQAF3NM0kh1mByyLeY62L0hkupAdrd+/si5Zp3awQ1+s3lJsn
2j/50/FJntH31E1blb47QpdRBMjsbY7GLmECr/YQyySlE3x3VE0xWokzMTmJ+6Tx
897pNEikfC97m84vgWroYwKbz/if0q6jrZxUofyIi4gNyc/hoFSn5j3dkLizk27q
exHQMVhZPxXfRqyxH9jGU62vmYeHWnVdShmjIetJj+vTTiIu84grd9/rggtbWn+k
ayyKAmQogfhHoX1ZcOxwxi1vNwFB7s21NbtrX++XnsHYZxHKrE4dls+QV1uHPYYM
TwGgVS+DKB8f5RGSo//mRCD6GSpq9SLVXVI2hrx2KvG8qZVfsinqxvpkjxUvJdRm
8OTJ1daAhu0aQ7rmqSw+y/eZlPDmxUumjdWnHPL4pK3CwbkX3ZtS51p5r6B4dJsG
U5Rib2PgA4H2ADV1MW5ZIV/k9Pihg+bMBDj9nEWaw0i5bA0Wc2L1uNJVGtbIUSaH
OmaqE2Ptt4ujRyYTu/l9vA2Kxcqw15ovRvGo01SGMx4plDViRtzG/AS9JVAHtfoH
/TBGa0aJWbpZryoEhyodQFEL/AljBiLW/7Vku/BycAvEx8nmvf6yQ/hmW3BXKmvD
M3E477Y0OuXmKbQ9t9pg7zCgldBOx6MYVik32dQujV2s6UcN91LBbgxypWvT1fOd
H9KgvlKETRdzOgnDtN5OXvf9qZupFaMDSMwOmzfNGAd+Vmo/ybZRPw7zywa6zq20
n8Q4u4wto3qEbKHnQf075cx25AliPLY1Rhy7BA0RJ84D/bXGYlMIBnCexldCoxID
si7m3P3JwMYZ3kywzVm5BMOWL6qkMIzR66qcQ6S6DOL2ZCB6wtP3Z3dp8RWeKPOS
t1cAIhf5TGLCwuo1CO3yUZv6WhyKI78umtT57YUkCuRmm1SgqvrUsf4xpplb/lFJ
r8TuIm3Skz/egBK2vb8ddv0tuMf2UYzIsmQrHkYHZlI1k0mG6E7+EVcAkro01GWn
7jLLv2Xjt14KhNJFboHtNySol/70CPQ6C7MUfsQr1340ar8rfnZ7wCffLOx9G6T6
okdYRqW3wKoDUz9pxSOZflx3j223L0XHaxzMH8qZqdS0+yVn9z8xGSY+fNe3dA8S
5QFs1yk611iWlPSFEl/3ZAzGUdZXyufpI6J4hOH6eH0bkt5/e2f50DvftJLNP95s
oRSG/qisg56tdqhw3PclQBcgsRrV5H1hemLgK8NZVQKcTqU4TXS/oyvg3qsbf3Nv
0SmCHf1Wz4hPlRHHglEgpc+KT/zAAljHmUo5oGTumxEv/MN6AREWA4GCCLLZaaAu
yySM5FqVU+Bwk4Vcv6wAqhea4SGCQ9qcO0x2Yb1xHI30erhMISpNxwRywlt3xrRT
qecWPOchSqId4LjqP5FxfVchC2ZXC8D3zqWncqMmBCl1OvqKSBT0F7wH/GCMdg7h
LaSwAgzsojlHCN9g9hzA8BjK5DdOeoR56TWzkzcj833093LGLIfcFACZkRPp9HmF
bD1erXcP0ZzrVNp/GKLeaMOr79ZSv1uKCfBcDJCqYblielJ/S4ji6U4hqWWCptIa
P2gyzEHVIuSjA79I9OPHDTIYl+906lPci3vW5vZAzhKTMiNpY2jWUKAVSpiJvl3/
ty+50YOnOqrrkTAkJqwDpJcWajz8EBl5PZhdF6nWQJckNc0GLvkhBlk2PPacuBWz
8GYPIHL7FdFu+u5iX8w9qnocSLtdThOqwU/tqW4UcHeOd2/6PG8iO6cTIFD322uv
A8CAud0miOPpuZi9mnRrnUSUAlpL1eOwPcJIN/eKTqqE4McPX22fVQ6BEkGpmQm3
Dg1NG4PWAmSAxhRFfJ5klfl7WwKqwMZz/51PRAzd/7IMgfccH6u4IdBySvaUuMNY
uColVDwUGC+3QW88sBxyyl4lRsIcPl9zD1JieJ+vtlTaHToIUfET5kqEbkYVAEoM
zTltcmwNavqBZ8nONSObWp/ZVbzWl2GBulV9vYAF7lhnTuF+MhzTeQa7oMveXkYC
031w8AOWxmA4DSxyO06iY4JJeqdGMQz4A9HvhxcNMRSKXaZDhgqnsAqooUVecuFq
58AL/dGRnYIyqSoS7gccrgteH/anb3EmemVLMkWTjwt5BoBc1k9y0xVXeeGl13T/
V1Ma/HkupGI33aUq9GcKNg0wZtt/Pel6Z+O+TgKmw5eJukPsJo20k21+ex/JaHno
25piVDpuzcDytEw9S3LFJ2v5XZ26SOxZgfOOP3jPARwSXdgZCboZxrgxeu6vAQzd
DkbG1m4ifIxAAtsmFDvPue151R/6V59ZrWyjg2mxXMe6ZD+Boq64UhCu/Xbbt9Q4
rKxFEi5pOr2vzNkRN+doM6iil2uu/6ikbAcPBsuf9JxxPFHIA2Q6i/v0tvrRL3Jb
8oEB3po41YglfuozhapnLZubiTDuxkir9gstkyPQ8uCHAN4SiAT28n0FZIPW0Ueu
19H/zq78stsJQDu3TRqJ9Hn1/0E+Udom4dj5YXawrJttjb6cL+A2XtqqxCN525rl
kkFl3zOEw+O1hCtsAeiiAwed0CY+NrqPcvFo0ll0y+6kyHOB6xCS6INyev75nVbg
nHhJwnTfTcijp9YLqDM0o4dn4rpGdSxoLq88xQIODtnQxmQUyV0sAeXF4QFbRu+4
0pf8cvaTIRD/7Tn4NpJSmkugUKS19GeB8EZNH+iYl7QaZDL+hj5tFslpHHc4ZYF5
XwvfgbTmmvOaupkgmFCNMna9dintNFyF9WZb578FqZ5v8sdoBBcpHRKm0JC5JeZo
FSujIuyiveQXNOkiV1vczFLUUVpG/x5+W0anU1kitrzhT4128duSOZO6NSMea/y8
j/V++WmYjH6MHho/DmhOsLHOSCKyZBhL/uQMEY9WZsHYrzZlXwfRTB0MsVVTI71e
jxOxTePlF4EVILvDUiPKL8EuULxIq8x9eP9KwFU3yewMWprmtsndidNv/cpehoR7
TXYoZmE9AxcDCHdnNWufAONe+qlIpHyFHchfQKg5vkxg5onDYRIMpSrUbPKHP1OI
RpG4j9hV9/m76Of87M18DHuDPhH6qLVmWO0MT5NwMm0rEG7B1hpf5qecBAXlFHaP
6jxFc8NL2/1FEluw7z6DV44IaIAfRbQ12zMxYHbiTtoXmB75b4Gl2SpMiiD5BN9z
j8gyUF0dIF2I85S79el4989BwGjJuz1ZzWzK2Gg3e8thsitRbNi64cb0PnnCLbjU
w13FYrUUS5YamYu9X+EDwNKcJcZyiAwc7v9w0Hz9pZvx2dXvisPeICMKAEGPxSBz
JsaeKPGkE3tkPx7GThLyruL6ewWsofItCV5p1q8192UsNO2HbGp0k8O4d3N5T2+V
ARGhpP7B3yZ9uFyugaElczQcYf5QyAUrvHqpnpySqzEx4eKzBYquxSyZpbbGec6L
Zk++TyMeQsAi/Z+Bd6+ZAtC/iM1GFOqMlhOzsGbF6/zERuCvvuErFiqYBGt28+MN
0oUlKkabiDvXgvHEvnCGd3UEQXqiUhco6uUS/ng0K4/kg2B8fDaP70oe3fN2USTF
QmItEK+5GCM0+TV0QMWOHvH2MdREw6l/9FPUfK82aRHwSFq1NDaBJr17l5M3gTvU
+ikGAohLO2lNb3PVbgfTTJ6qOp7FSfkoJinYrOp+TQCVqnD5uA/FPGfpFmJ7DSm+
448HlWd8J//636WV1NfJ8+p6ALhUk/ZPZYAxfTmDy3iLXdqhXEOswCkfgyJ8Ru9G
UbckP11heYECvXOVrkzL4U+qJ5WgvewLCmjxnGzd6k43VZJl3YdwBPxkBSQr8Cyn
dsiSmgq08pMsSjTB1Dr2pD+SPpvcrAdk1gZBeq9pB3Su2hu605z7ay3jQLSSXyQ9
nUXuQXF1Y/Fh1JaoUmYMs9It3G490m1wIdJF1smMv9lZ32YofKuXLH4FamtDAhCq
4jdseJvRfAIfPHLzSsGvFCB3Noh+dXUzWQLZaXnDjcgSg9mcIV6kdjJ90ESositn
f0TZ/zx6/WNeerFXanU+uMcOyzxEWUtHhwsTfGVSD+yEOnzqzLGy9S56vocAyCev
FOl1DeD1jyR0YS4J/YGhh3jej0A30A57dSVfYBXCnA7EjCTLZU2j2se3yKEt+9ab
+wZOZm1CkrLs2fjrATk/e+KRca0iCGmbkEilFa2hMy/eufgNzj/5P9WenzXBDCiZ
0B7ukC0Hk07rlhy0ymvNQSa0Ey1D3yJZRDAX2umdBrVaCEvn9RNn0j3LdABE2l32
fDWyhn0hLZKJu9JPGpjP5akWkMx5hcfs/j9JOF7Fx7lZx/ZBAcfmfaKN1So1xcRN
ZhIGksFvc5e2uu7dEkGcEcyWCZMVMKojQs2FL8vH1R+jQYK7m4RPRq1iZMLh/exn
32ikOQWWf/DY/KSpcQc9xKqRR41glJ2XrIMbMj3PB4vNsmJ0sZZ0cnVG4gDzgh/M
aHSB03CI1fB+yq3jFfE+wvTHyPFj66SO58raxnIhLVAMcW2c3JGBUnC3uz7gu1HM
PJa9GQbOQzBY6/EgUjPXJ8Uj6Ur//GZcyTDOZ+gDbVb+FMZVpTarFFX8H27APEWW
OoskRTUJgxDc3BBkS7wjVsmPB7SSNBd1VFgI09nf/pF2B/NdFMd1z3igwNZdKxwk
6YHG5vFRTz/3KJw4EYsm8zC+VCRB3xInhhACSYpLVcvrehcZkIeuiOHuA2OsSpjX
QTHRUunkooC1WYrs8TkAF06O+usvhvegjPV5NsvGTEP650F0aZ1A6HUu0LZpJx2H
7HTkR0JKnKKbbmppXDjzGk9cP02hZaPP3ErGm8LpZengAZwCp39eqG236Ootcvwx
sLx0RAj+P73v/zK49ntGgvMa7+Sz9lWmrQVeZlvJPKrXan+rX1f5HwXqendwgrV+
AddDEIsPvM3a24FUU1lNm9GKX/YDUwe0EiLGLFNnxRTYSPtNDPf4fzX5qjhwXW+D
z5ETPFxgOvV6d2qPfLowbdGRDvPpX4Z3CD/1cUcq9tAt8BupxvROzpe7Jr0+vstz
P3X+esH1hsEiU5CY6OMVnw0dQUB5WhQNLYkhDK7RI47BMvblqeT3E4IGQ1SMd4Qm
ompOM8M2knMTbEEJyoCsgWzOU6q7DevMt9WvOtIwEVCBtRhjjMEuxlYb69wfNrua
z/S9PPjP1KWhlMkpCChkGmTcJZ2CSNJugu4VmB4/6IcHQ8EHIsaefuThjSBeLNiV
PzxrrkWLpwUqWVDvlbgza+reKoBWM56YTmx4emxW9YpPyY/xrTMGPYy5QsWRfyR/
JVIDItHursgyiwTtHI/itsCtTj14KkEa8SDpYUE3dvDLcdktCPRgc9lqc70MaFYV
Lef7NxwQDv7GhMoAJT7byHIFEySDGa/ZLu4HU/3J/JCN5EKmTeZym6XZJ13OBCur
F3j0T1u3WQdAwk0wZUXbroq31qLuMo/aYuBKTsH+pAryuV+9noHAHesgLHS8+WoU
CMvC7GBZYE3DD4K4lyh/UWWNbArlVyFM2w3KdxMllvSDgwOmFYqQsrG2+VKnKlNB
4j2hEGPKuX0st7sHVrqfnzrRf5UjDFgXsbDFPcKrXEqWr1BvWqN+dVBFVQNm7Vcl
JiQ74kos4sHq7jAjYO5+/ci16rUpBOUueQd2IKUyyyQUWt1xfHAg/OOCwWBUt9Dy
FM4pNk5MaQtBrVWjD+xdrugo+9v/Nb4CzdmpyqJrc5NAdNlJE2QUmQU7BqM4FDrm
UbitjyCZthIuU9op3Sboe3Nhir/OsYCpoRHNmEhYqiJs5F0nhf4hM0ivucqhMs6h
XAZdwH2sfx+txd2027OxOT62vocb2i4oVA9XrYj9mgPKEg5tU7gPW6PuPY2AT2e5
0YTDb3zZpvZsZfcKFu4041XkR1L8IPHO/q3NKSviEpwJ2qNKEtyS+GoSY+Lnpgkq
2pO/bYQvmJLvo6zemvU0aFf/ZRA0JArzWc2TBypnxeXE9n5E8q1vz8WfvBbuCC4B
/5Tk5GQ1nssoW0X9SFl8LjYYVRcEEiB5q8Ka/8lqNHUyp2Ru5Z2/3HnlFEWJN2n2
MuhJ1OwaqAmDwSxqlnsXApn6nWX8fZZfAIVpiND7cENcwP6Dc0E/6BTO/uw5SHLg
DVXi1fyoffLU7w9qX4emENdcA7p6y5YUdBL0ABJ0Tm6xcLk8YPjEdGSvXcqWL6bz
hfztBA09aZHOsNgZToy5Je3Rb/ye2tWfiIInpgfWOUsWw0yZXhLkPG2qySatJ9X+
lK3BXZ5mghV+XfZqyHIagV4Js1BvmxfO+vkF+T1DXBozhVtiwaoAbm9rHaqhw8tK
jIYDZf+opzMFH5FHj9yh/n+qYvBsJwd+kohSmzBUW/mwkTQRabOoxCSuBXg4obZz
v+5IF36yMW0JSVKQim/hKZj1eGhMSrvLK10cPkynexjRwkqFmK8EM98kOErzOjh2
StBbNVE5UbzmCN5ppi0EKq7M0OSKrdkbtBPtNSdn5EnzOPm3lQEdaW8JXdCD794c
6QCa2ZiElzAlZC7KwD1AuNnQuCLwrqFuy8tBuj353dt/DXrJyLXb8Fkpz9J5kTDg
7D1zHyZrAQWlkSNaPY0kNbbs6Nf0K9367dOY703scOmBYVsT0uFMiA0dJiWd3tXr
7NVOmN314u8qyehkjbLfi5cDdqLKeciH1eOuod6j7TebMOXlJ4zhXkxoFtn+y9pf
/e6aZkP+GTiewWEZ2omO1FJDxcIdA9KqC0MU+bxR3caxT4hii9tZ/jyEgxA4Z+sO
zVmyBrVya1kPNIADnZEk0wNlvAFWfJiQ1t5onYRkoDaLOYp/obPU5OynXoL4au+F
ixB/IEmSNW3NcbeQDRLgl8MGelcgpwsFsJU0YcNmyv4gEr49h95k4RP3p+k33D5R
cstLtqlR+39+R7hvM4aQwtC2kqwvW3bg6CpXGs82yFMsYoyuJev9afLfDnMS3WQk
mU1pxrTKROsQzDlhNLn41LbIDVBPCOOEKcvrWKobw8hSq/8UkQ5t6yDqe8A3FN3y
GPG9r3fcC01l0goHTNrMGtbwcEnE52ZlOTvhIbDBoEt2irKepLlCR0+WTP7GU+CD
z6544RnKc4oK6mIy/OBiQ2JTYBdoIbIJRIPA+LQcDx+Ug8JEqow1ziAKaFpJggNg
/PaC4BVhwAEX5thqMC7kOLnKzgOPs5ZIcxlsxi55GZy7kIPHOXfSeolEioYqgg1B
aOndVg5EY0U+sPN4jrOrUjlJMFCcVpdIkLrV2Kqg53DP1P7p8OVbSu17ExaWBQ73
AKV4bGeqI/fMkxgO1AXkM+RVjs3JcqaiSwCc4yXEps20uoiLaj+m8zCPK7zB98Pn
2qLz3sftZav2QkGMdzJJldW64gswIEeaxRsI8w6rqUWp2CkntiQ93C8o5WtOnC0Y
bH5QCv3rr1n/VECE/tzWhKK7d3QOWbquKAkE0U+i86RSQByoLWer8o5Zh31QlJP9
FpnEHv+DznBv8pbWkrIaf2dr1LFs12xbeRq1mkhU1Jm4yCUfjz+0oBIjs/1F5M0O
M30wzZwosVmh2lwehVvePDnZP11wRNwtR+h8wWTQT6xKQMx8j3dCmyurb4QX7RD7
vMZYIe91SqUGW3Ytboy/4y1MYnL12o3sVaE6ZlQrgjN52I4Ao9Hxgi8mi93Q0jtD
EIWepjJprQpwwZKcJ6RIPOszMgtpawdR7Ejfv75kN6H4edOQ5+LCfVEHAnOrvaDj
F8I1VUk/J9cq/M5hUp+bp/PKO5Eisr0NqihSKh7Ze6j/CeIf+hSX0XmyrY1uK1fz
A68aF6aD8kEAPuteum1RTkJ3fMz8s01XmHqS5Mfeoz3R9m4/TtHMKkb4J1tWLWKO
0HGzY7X7uzknKenHGgaq9pAB+fxsdwlqEHRi9NZ3/VVwDOiOKfuTjdNTLS6rLhkT
/e5mhreCQaguIkW/+bQQ8N4oJn3g53DtsadJXJ1+MaZ1jzbj3FnH55HMVImsIdlG
I3I0J0Limgn2dP38xITsqaQP4W+ThJZIQaliF09TuQhHGJnx50VH5KdpitPWZ8Gz
UvFYaS9PW8mTWLX+dT+rrirBFdFTNYyNkv+QkKLLezQU7cY/pJJUFlYxdd05dv94
PHSGS+hL2aNTFFSmBSiqw8z0mSyfTvpAiZQTRQ1RwcHUayfSsY9Un4aKNPLyGrcN
GGt1UA3wRqowcXqzxMXK3VvvmDE5Hbuak9ReGQQKZhreNiwg53JaM6wnSmuR6o5f
6eEqT8QxHZqig8x5p7+8Nc+N4/8U7YmhZO5ioXLxWWbuc+QhtkZru0H1/urvW31C
UhWdPHMO9pvTjtGVPJkMUmGILN3E7hZuVNAbKuCuCjs4X5oDaygwoh1HKAA22LpB
l3xhM50E1wP8/wWmCYdFYsHBrSnFahWRzmZmQkpn24bJG7y7bQTnzvuKxBtXI9MV
qpy6KqyJLt88hVJjunoCdX1SaHGh/UZn76Qzc31SLieaahr8g/y9X2j1MVevDGuK
sI316ItswK71z1Rc4CgWxDa3vx/Jbb+2P4SMBpveoKLFZlQhzraQoC01GpJnY7EO
EJt93cYM5OU9x0vBAngdNabvcd1C+N4UfzcTk5MUvmIxHvs3JQffaH6hBvKxT4no
p25vjWG32kAOT2lDHu1oNY6LeFS0u5SZpAPZf3vCVV84/j5S7YRJAlM0uoozljAC
kclDZOWuJ/slVwQxU1kzB/rJJWxztLgZtq8GHiVkcxYhMbH3fYezoaduFDJj+5DB
5KuIvZmo4L/YhgjzoUZ7fHHUVnLGqUL2DPKlwH+kG1u4cYJWW5dOSF/iGzq4Lroj
mF+EjHcgbXWBneYZ2j29d4wvW6xCGg13194r7nc8AUnBSL6dcbDv36d32QLTiSxY
rHGoljB+fnTQQnqExX+w7+TD1RvpHmLWXxl7PxszIOGKyjqVmQcRGkmviJ63PAT0
JPmuGOnKA3yS+zche3TpneI2f9qej9pLFAykCMHlW09vEI5KWtYCrjdQs5BtWk71
OI7MpJVVa0YKGR7dPt0A0iFbct/RWx6TxarSPi/6xfDF24+4Xj2PaS6roEHR4gSi
Ws6XEo2gquM0fvuk2irUD0IPXpolmsbJqVp9GVyU6cOWfn1KUnbkrrh1iaQcaLGe
XU+MhI3445oqArFH3HPFzOWeK/Oli+ioKAbEepw9dDplWKCK+IN6f8xoBsLziPWa
LLeWajCgFfbQbei7Ec2Bvv1dP9+bka7NcpNVZXY1wwLlFIcyi0p9KN3PLx2s1sww
ri7QWJGUPMeBuncXl6UJzadk1x37xR9ultDAlbu0g3e3EHBSF3UHdorwf1ST9PEI
4HH3CLsVP3Z6CV44pQik+hDHqShHBS+qHn1nmLk+ftX1nC+imQ7ZmuEiJ7y3dtL2
NG714Aemkq518xh3YmRwi1xTv6S03R0x+5PqbbsIHQdxJzid5p9C2Y5fk9/awpVc
kZjv0Q4tRWS+OAug4k/oyVMlJ0gfgmTwy89kxNiCWMBKZAMdNPy0iOQTVN9U+6G1
ZvCy0871ZBpHqT/A+F/YvYUTgC4BSI6niAwBFc//8zUp6z4ZaYg2CGsRDwMLAOlH
g+ZmwMX84Zi+7+1liQePbzP/eS6UlxWROkZmyYXAkly9ad36KhlL62uGx5asEUAE
V1xP/zVRWrBvU4evb0Y688MZecfATqkzGKBBH/jpTWPpV+EGrb8/39OLR3nT8fLi
Qt90NCev/jHWbmwZuPFuqNWAPHJETr1FKZPEnKK4sR36mBYmZuhuvDnejIwwMc9d
bhnLtQvZthOJkXQxxpDY/M4xX7wRDIW+drPDcz/GqlXGdOPwwnW0U72M+sH5fKlv
mLMoxCM9p9WHOfdnetrJeX0497au5tkoGiLJM5KqY4X5HIHknXzANYB8Hy/p/37K
k1NXI8SDOhcDBasTtwLGw5aym3nOtz/y3Zi1c4fknnJtEyzBUCp3iPMZ9Xi/tSze
R0TZ2yzY8xtgFcwyd5DQVVQzxj2BQ1OuURNWrGQhFAsuPWzI0gKiogaYP4iP+JjH
yo9rh9VXA3Vwob+xOmPxmJ+JvyTH6BMLM0U95+mzh1nNZv0HVf5/kO0d49ZeBN86
Meq7gxDMmk/G3puhKQHcsHhmD8N1KDOBW1GiZZqp0fmVJPx9EGnAfrMp2TcBSxJ0
4C+SpdF1rFkgN6q4KvWJ7msOOx/sD2gHrnOaRtGEIhtds0AkJKZTobFGlkBhgsvl
zFk4Ts8mTWqFJPkIUcuy+fmETCfDmUOel10inGNY7l0rRIS3EcuBCTUDvCKqpPq6
cch2ctu1FUugO8tjiOg6ZWic5Mu7Em5ckkGVzw2xVtL9Xu+gYfubGOz2je1ejkJu
IHxKw1XFICcZQ+etysQW8bvm15F1gbwlIx/PQHeAv41vp7PD0nvh4NvLB4nTUlG+
LL/SnBzenTtQJvP0bANrDBdJe/Fdkcky0gpYrqbV1VgfQ85DiwzlrZEPtZifxT5h
ZKtDEgVGqlz1UDDqdnmMoYL14/Dr4VZNrtY9sHQujD4GUU9FLedu9AQQ2gXxGzk+
ReiE+1x3Jbf6jmI02UVSOL2+Xp2B62hp22cQvslZvxQVM1QsqZfK6dSyCXrjE+6/
M3AyDjwHqYkCcjM6GMgTgKVv3xvSCt1x3RneG7KKkj1Mrbit8q+P/5oUqNlbdiYw
ueeQ1/kqF2/L8vx1xUFNwCMlVHiynk9v95ihBz7yvHdAS071vC8ubktyfkAM6SvC
G587KoOOb1ZnGAVhbs/9haZbUvBTF6w82U4k3kQSkWbyNNvU5Yht23iMjiEnR41P
h67W7ZDwOkKOkp30UGKbCjH7bYxh4QzpImYyPcpUnByC+9o/QzoSgFMuYP3l1NG3
mNMxPdDsL68910Af8S8ckOjJMgIASIRdLk8ZUyNK+SiIOvNM2vrfZNyccq1Y1/4R
1qoe9pAo8FPNDjbQN6jXBRICc9jnKXrS7Lc8sqZJmziD9sXV2IWt6qVih8Cz8lxH
ORffIQS3ve/M5S029LlPqjfQkmQ+Q0TVicfsK1AxL/ESm9+krR8RpNG487WMJ4ix
eBGu7dHOt9Fp6pm/4PiMhiCdFvTS/t6QC6p/2ewlVO73YavZhix8VpmENh9eIgwh
lh/X94F3QvSAD8IpHJAnjYWNj1OwLLKz74WCTC3/aCFwoYrp0BfvXi1JRu1f5ANH
J/4e/M0JF2gMsltXVMo9HVt0qJWwkX9ZN/Y9C/gf2qR0mCv30yeAX6WPZ1ahWTLV
zjlSIodLVZYXHLRKOu6/uENqsFpnBfWFPUrOmI8yKzWVDMuGy5hC3RwbyykFQQXU
utl34OXXogWPf/USOIYYF7DFJxJFr/1H6AZexWNDaPy5E+w2Rf1ija6djHB4JAGa
ZaoCUvb2BtDqANmwJA1II1Afrsi0fhOjRBpH4eNzOqYIovpwF2kQR15O0TA0dgsg
S4Zy1gtowXfXKtFubrPycYdPAl0WyfcpoFrGWYCnWG7KLhcZhzNJNdckRRvqDAEM
NimJ/hsjX2qtmKNMPRoo8CAkXZQXt9LyNHU4/GaTUdz6C8AeosmAE1j13zFc0rBl
VHOzKtwnKp2cWgDVkUGEDvnX8sloD5zybCzTwvmv7DPTtJTrgYbQ9Wio2y3K9at9
jY4RyEcLiTk0R2LC8eJ+B12GVPNlLcUeoHY4C5LQiqqfoXJp4WagdRWCRbxTb9tX
HxCL/FbAVkWex34mQCGh1V4q9pugJvJGaqIB8hDYlnWX6DUN33SNQnWkHoQAWyaa
v7UkvZ/KPzVV6JImapJvvfLxVNC668JywsoXejfX9yqBb9d/ERQnm3QkyLTUD1nh
FNhpqE+fvAY0gz7GFF0nfhDr35XxtLn044mqDP8RV8+oVDgNEEpvU4P7EmWb2T9L
pWgIEgQPiVAsTwuGVBLgo76NiwMqEUxBDUy1rIPlpbM3OUS7ZSvka044G2HBPLP8
XC+Hs2Frr0kkHupdaj1iATm7M3l4rR3ToTfMvSj0Z3ktoN7pPZ7v0cq9Y8OonMfl
CVStvOmmDIut4D58Y3u6JVCTMB87nM+jkIMGGUyutrv3fRrvNyQdbHgaotzUFyut
jHNiCuJRkMvFwlRNF3SRf0dfF4XjqQCPpFCLC2LJ7hZmox9vQHbXiNRHDJqbJMX6
WIg2POUcbmsO6hYJ8Xw/x2M0DqU9GFDFGEgkKxgirXzgeLQLREE+YoI4zJimrZwi
udIqXTfizSS/t/AGRA0A8DI5f357GrvOHyZOMRAOyChLZhcjXZ6Pv4G+R6+XBX/H
euJQ0tlI7xr1fmFDbEwwQxC5tB3pzX+wTKDFbNagNSIlAv8kfMvWP4Lh0YB5Acdb
DBq6mqZZVjRXlryfn6XuWbm9XxXis+YSPve+ug08BBi1FsLz7g9ong8SyTimx4bN
XBJwit5tLVybhr+8E3BELoq9MmSthuqfv67g/p8MU2VsNloK4aqG5vtFGleRtTPf
twEfK+QGkSppF/D2grGY/RBTtChtBgSfMWiJM0tvgLUSVTa+QwKi87U7AlewS27a
EtdkT0cj/SUySLczRHYXhZOmt/TjMqjma8mjZebRSHMhkbVyzWePQDqGYiFEfCAo
ho8NXbgaS3vvoHCLf+wV5ELhBBmh7Ye7JCnJv3La0rNgJFZPrgq7a2xsHFMopLng
sNSVkfUGIp4pgwtqMvyXTvA638JOsydW3OtUm6aIuUhsQoH0z73mhE1/NHW/VEfk
fuklss1yqMjQF2WWBQAyhkJWmhd2mnW9cliMwHfod6QzDeYMi06C4Xcaj7/QWfQe
cTqpHoIWNKiNStzBHllx6Cwyoye4NHxDuKhCSCz7yUR2WAYE9lyjwTwu8JE5e96b
QGhvYr3lNRqM6RJdD2WauZKPkLWLoRA8o+n+NnoGl+MzDH51Z0eFxZk+G6CZdTqH
4cMwrX8cIxFDwwTU6poj/m3X+foG+IEwSzfcWxe3FVpFbeJXMdxZwmmABRR6vzbh
pLbszQW7s+7P6OlShduoRhibkqY/5EYe9EGH+zOn+PVh6xKxu4yFxI41/DpUf4HB
mir9i533pYvsoiXwD7LFINcV+6mSr5161MZlztpqt+p1eSy3UrMb4Mz0sTDsyEYw
n4dih+kpNLG8rAbPVEm6wXATuc3j4b4paLNRtFiZYEIPImHqbyyrIrhzKd96kN6N
R37ynifgztT8EUSbSm21dGv3u1X56U0DoWoApG9VmBVqxMlVWnMUqCCDJyXOD8YN
+ukz/U045/rY/Y6UPEmL8HtaXqkyDb2ev/QvG6IhZczaGtP2l0bfwOQ/aLpdq6mv
VssL8h5JGBRiXuR8GpwHahueW7enc/U9c+zDnxQ2j/91wVwLhiY/8qTf0xiPrzXl
5ujKvZ8kMRixj6x5moZ/Djd/fI+nzr3jbVDwAa/NZxgkEfUx5aGAcoLBjJ6sFspX
CpuLnZjeTSb6Rpx6+Rvy3XPTe+dCW3Y8uLD3nNouDzL9uyrZ9bWJX+fMuLaFHE8c
DbuK7FsG2EkwjCI5MS5bD0gqSLE14Gx+ovPtUnwjoqMwjwJXZr3CmrSOtkidPSMd
EZqHYuxUGOPggZCX6PK6xp965nwHbRQ3axmGevlhdRF+qnit2Fp2o5lbjQQsKOWT
yhOLRJ1AXEk99v1Xo7Az4YOMhRuM3XniaT/rgGyuVAq6HMU81oIeEA/9KR47ruUr
gZrUmg6LSUU89NTUPA+i06ljbkQgu5IvxVrwdIBKrZJW31JNeEfBifL1naLj6Bgo
bzXde13Awq/bwDEVz3JL2+v8eoyT/1u3SZUFaEnmyIInadxpw5flgVW2hUI8r/hm
mLu3nNTFiZ22JZO8sz3HQ4AkuGsImYYiKE15t/QQoR4tnWBtWE1B9uForOfEZc8g
PsYeVYe6vEoILHRTn85u18vZqZx+1OtPmKNr0eIaXmgx+oHSP5/mSsYUJHMB1lJO
E/7cCQxZcw7KQ8r9WyooqtjPhQc1eIe3QbyoytSgQr4EUQeAM86IGb+cUvIqOm6v
bBZk/90mK3UF0pDE+/KN4RRulxxhmbakWb2bcrDewcnwRDdeG5sy03UJTZpyJ9Mr
4lKWDc1ZUou3YC3TcPg27L6RYzZcqQxFiB+4kPZETAPu8hsjgF+mKk28c/afxEgs
cq9UJVCZbBNfK5dBO/g2SY/u4QzRE8xXWs+ZmVz+7L5OSztnkmpwUU2wAJBfZRbp
0Ugnlj2GuYE5M2PlfXR5kmgZL5tpv4xK4AiWXvjeZJcM8e9idc09nnfz2hTPe1th
JiFMXLnU5AbVG80rKofvQLaZSZ6PLsJ45zrLmTKjbHGZT50zfATy091YIaHFYSMJ
OHUKEKrK1SIy+YSv2Y+wRl1Qjt0ADNpogJF8dY+/mb3o3pWhobA7d7ywvkQ6xog4
bdKPV0oKaqwCziT3kOWbNtAPtPh/1EtztAC7663IF631yB1lU/JY1rohbrrm0wbJ
YRuOs8QKNKmEmGvWq/l25vsSgKf74wVk1LxRrZqtit/nnFw/05t5itUM8acnGX9E
Q4xDULD7z0zyjn+8Cajs70bvrV2QgInxrW6bYUYkKv17+qAvuePJiOYooqkf/T1J
fG0sPJ/1RrxBFTntZfgUKzaHVXd/w9Ez7Z4xn7KxUDEA7omQgycXFbReZfOanxIG
PgzUAoQ8bzmN6VsZqKvvJKNm+IjxVDDyC5QyavPzaCuLSTMOpkxj/5Q9rYCceUB0
BYmg5n+wjuCx4P4Ex4+Hlx5G2iSA0wJrEiMW/v+OTSRBwA6qMsor0IIyYwLiIfwn
zk6Pza47hSkLwv5nih7MMMG/5TKRo48UrxXhrSsXjpNrPmUa9CEr5WUbCXYvycvj
ZmW1PB2cR87/SbeB+/I4uGvQ8l3IBZ+fO56PDeo90FHWfDg8s4XQZopb0ROuVx2k
eOAAXyTVLxk4KAFiE0NRJDcKUZoCbvBA9/PooCymSfHEIb3MfClOzf17JsQkpjzA
mJskXjjXVsneyyqLRVk+jyv062eAU4tAxqmbngH1NHdTr9gNrzyMO19vJ0H4byfM
xkHc+ZmrqulTWQs9jrdsxn/mUMHusIb/1i0e0vmidvULWqSbaojDMz3l/W9u6rKD
X3q4Ks1qXrlrZO8pa8DdHyvIiyUpnf59jepIs3fsVa6KE09wIPGKbaGwg/cw2eOO
GwlC8vn6PGXk28xuOF4gxESQIekZBHnEt5nGkeCnrVPOsiMsRHKo6V+qBtfZweni
AWL2t8YzXfWlTIix1G6TBlKf4so4uvJtqRXkFdWVlRPQh0pbGfegT2aVLLGf4NY7
qObo7YkyVccH2wGaHz36WnyGBMC0AbYVuwzqCti9ZygC3Axo3WmJS/YO1Fl86nc0
X6jj9Le4QO5kzpm+Lg0BbplfOxRidEbDNeVVqU285rjlj/6JIpuOh4yoyHAyTQZi
M3lGV6FRvXg32e5u+hea1c77/p6D+KYpHGOTPK7uMgip+2usWH7BbCl2KqTgnMi5
vMjdgg6D1LBlE8I2RyvNqNSSlX7e5/6dxCK3dxlnjIKzsBSbvq2LjJdWFJQG+RLZ
swTIYe7vxdt1KV6FQx+xyo4I178AFL9hq29yN61D627tzJVkYmMBtr6sJOH4FhYQ
2ocu4X7a4rCn/UM7HyPqPbwR9MYu1cdmTowmTJRxDOcjQJ2VlbIJdXfxdj2n+tfA
3clmKO3jmcW6Z961o2klZdOFb7vJzngs2UAY+t8ooNSPTWoWMpPHA/980UJDLfOn
vNEHA78+/KypsmdgXTk6UvPsgMPVu7pwIYuCGqw4Xq8jkun441MPLH02Z6wJCKad
+PFrr4V5JMvVv0g4SSwJxnw//notimEv+rhjyW3s5ptuJcvtqUCiOglLBglrWXz0
MGQT6WXf4z0kuCNN9BHElb7ednyV1siJvY3YqUbBhnpWRmwCIuV5/3RusH91TaKd
8zO/tVe1jfsoLkSBWE1owZSE6vUGNUByvEEO2tDsrUZGxi5xh64raWLFfDqV2Des
P/ypWHIcov2qDnP1SXOJNrCPxqe7J+KwSfoPaoxI0Y3IiC7k3QOm0/DVio6zoIzS
vmiptzNWjVTbjm6/lmr7cTW0YfNO1t78opQkDPRfZHPESqea0/WuCenPHp6jiRiI
TgxmFWVsybOwXQW4FlLR/1EQS5MeHBMXiSc79cI7SCff8iz+us2p7Tq8OKPhHyjs
gbPus/miqwHGgHQRE444OntemQtVaKmIFIyLX5TT0qy1gLWlK+RuQejoMHYUvZ4x
obm534YvnuGZa1lARihuV/n1/Nnqap+caIKKF1fhVmq9yn1M8b/alDuFEwFMSP4p
6j7NXonz6GM0KeCgP52Xoz04VadpCxWRM+n3chaqodDLG3R6k/1eg32qtX71GtOM
Ax8Z8KEDQbC0jRV3/xOghkkC/VvqlMcZqpLi2oMo8wIu/MayosimxlNVIRTGLw0H
x43GL3dLF6O9GlKqrXcne+m5auiA/VtpIV4rfU1x2z2vN81wiyIreyOGZaFFrgq7
ng7rxeFCOMxSIelbskIQKuHv4y9ru3QUG3jJESeFXKRYXlpMH97gCgLPTt0nH8rX
AMSP9++1ZzA/gq7dgpCDcya3H+E1BZdSkx8C3Idvo1o8DChm2SUeiZkjXCjcF0ct
1qkGw/hYJVeURo9EmcvKi5bdkHwDTMaejK6ijGqUHaskSspRhcS42EpfxviVJvAE
lENUZy+t6F5BOPhLDGADlHxvSoq4XW2OtYnW5fsHLOwVB3RlWx8D5XkxsYp5eerJ
a8QWK1ouuU8qv8bOlZ39p09MCTFPClZxqJL24XhlAGYEntSTfZMhmbYlO7glipYU
iTeI703boHntGLz31zrcC5I/XQi/xMc9zWYRvNyKadRSZH0ZOrCt8ymgTqeK3tJR
a13vGlcrZ7pRmx1QFkQxQ33I00j71B1sAneya5H52C2EKN8m+WbEWXnPgDU8d08R
DauTCqCclao6J/NiWxgcaiXAzFOul89yOUqPQBQDTs3sQbi/tS0RbwNeWIQm4CBa
Tkd9yFhcRcsSNj3tHDTtaNhxp7wknSf+UeAiAY1M/Th/cpNZHohrwxkoXE9Kqgr0
fboouZnE0ua9oeA/Z1Ev8YzhUF1rZw3jN3vNAufMw4/DvX4iKoOG+Dexqkc7d6Q6
4zKH+QZVauVH9jfnkR0kUcVGtgrrtUQnlqrvMDIqDs5iNDxRQ5/EuZbQhZO/smxF
WsAoW0Vdvg3ChMWcgB4WS5s3u6+hQzUQQ9K2Ygm56KgnTrAQYzJR8mGM087nWqzI
AzKBwHKYUjRXttcffLlg4+Be7wAhcaJCyTaropIqhXQe33XZMozs0GJQmHZFEb2D
+Gorbay0q1cjsAJ0SObwL4dIcdhP7v00yx2QbwlCCZgFzKym6lkDnjwcZAUVbUxP
PqjnE+7i4TCN8FYAH1w+blnxC+ni6ZmBgVBfcvXn8sqthFjBe9eYMZhtTN4DkAqB
86tUrcrJplRoOKFllPVe/kRZ4zw6foId8ngn91UPRlEQoI4vKQzTPRh3C4tHxgjQ
wG2jyYyoofF6eXcO6Y1nJThG04Gyhb7lCLurShTOaw8jN/Lrjr8ZDDBXCo7V1n/9
yglU3qDHXz+s1EhTlhOgnv9H/Vb87Gle0TU/tG2Ej6kHUpq0WB+8rfPmBtR23yhQ
/QE6w5VSk8Z+MQ6cbfEc6nMi5E7FdylgE11RwV2/QBoa4fMj3NzIdKz18KYgVA9m
Q07hdLz1PS7O7iQ8Ztl/bwvjmmPTp6GHXQaBfVTx2py4P9ITGS9E237chnrBuQOd
3vThT7CjeEc1XLN0F95JKAqjlZ/K5J2t8z4cf/llvZEp/kaRxVPU8R74dfFBFGyE
Wt0SxLcN3+1mJPqFagxCsuHrHPkzPpL0tzls+waXzVYaKoHlUv4yytJIG8RkyoQ4
excI2nMWm1TdSh+ET7Wlf5hnJ+QF+1NbZ/MJmwfqeIB0wskQD4yCDAAF8PyyDB9c
l3cIw2kh27OQvdj8SauX55Np1STYFI1r9fq9D7EPUNK/HtWWy5e+opr0xByq2PxV
lpqX9dEBhR27cMpXFemEQQu6MjKnROB74uJCv730eZ0FdN5gWkt3/HfYP0YArqkF
os+b5qgbq2IAzqH6mHWNuLo0/1JIjEgM1Xp+UB+zcpe39Q4REmpbjCk8msq5r/zO
FlGiNBV1+r/k5gXv/hgn8yXB5LBowJrVkU3yBQijpO8CDArG6jQzoU1JHszHfaPG
pE3JYrSG1CHWwWqyRFvn1UJdLSLUWkG3UwR4XWfnNafyhk7tQSAZHVmrip64PCNV
m2ehg3uPT4xditvq8yWXm+ZT65zEpGfFUUTIqYWg6chAoNp5pYuQ5XE3sJeMi/ho
qbkkK6/dKxvc7BASdBkl7IKs6HM+7PoeVK6+GaeJtjHAr0sN8E4D6FsZEAdFttZa
vbI224omhRrKl2xVBGi8G2z8svVpVP5reDn6nnWmFz42Z8h2dCe80l+qNnCiYOzl
oHp0pPUbuVa+ssHKwWjzqfi6Wx0hpar91+HZVPe8a9S5KqqRT6l5ee9LEtwnCIgl
Km4gIZK3fTLvb7upVUwLCyKuA8gaID7waZNlh3lHzWqQAcQvEJuEKVmbhwNAUhzP
DTtK7SoX149iDoNrcjtG3hcB+B8hTRAbo0qK13EOn1hBvIRe4l/6AU2UaKxovUH8
COfG0101bPFhHro0j4RpgTGtQ1x9oOD2lbu63QcyZ2tE4hjL9h0/wxjSosefJDji
CVAoyJauqziLi/fxkedggEnrsEaWJRv48zZrpI7P3BGnDtAP5/xoOsDp+JPdGFMc
GQ/SehmJmDQTOs/7zA2m5oIdjBBZ/V9Qk/kxVwlz9GuSgOgrgWsf8qThi3nHY73M
fZMhKYoICGDBYlBcnWpO0/wm8e3i8xJfFMlIoeoq1ZGhIhJbOr6eesrVrtR7ouvf
0uU27I1qAw3y9Ehj5GTOrxqodXdwtruwwwmRxsLy99b4ZzDbdirw2RB8o2+rPzfl
wXA+ldW9Woqi8H1LSconG0Fr5fdArsFzeJQBI9vEK3L7OUsegj4EKH5eiBpduy6M
NpyrPrTnusDX8Lo5WjS05ap6HT5pt3SYMFcvFcbLEDrTdMNLYCud6QrC2dFfLsHZ
PiFTghFpkkMvy9wdvjb0qA/hWNmk9rcKIGPN/S9wKJuAfXU1MuGGhE1FsLzHC7OO
2+WIAgM1Vrgs9FG4O3VfYuTCoX3zgU+y/DW/0iayLsiwr+IWe1QZ95nmgdz90KTI
dMj1CexIy47zx3fQomNNYOuOJoG/ioyUQHqzUYrZZnmiGnjnsWnd0J/6s269BkyY
l4jKNZeXBvAFyQqOVqTtVNvicJ28ARMlk9e+EtUUY2ref8EfVsZ9Uwb8YrDTd93w
EToRHlW2rkjwSIJisD0ZnBIkNPEJcnmH8v+o3ywWDDYGTixeJxsIgrcAF0BxRUP0
cocSB+G/O8jtA6UBposiZLJZ5rP/Zhw2Z4H+YZYWoaoMBpxY7ghnucs5eB8tIJbD
G6a6c4XtRv3etypFxPcjd5jKiBPHAubzhnNeTS2gSOJYtHPhHB5O9Oeb0b+lj8eo
szQVxS2fk4eiongdKkXHcnHIGVFL7Tv6uqtazTk4k89tuKIooyy0WSnQvaHDgQ5P
RnCVSiAxibc9pWuqIaLV86eKXHJGL+zS32eWmxZ7ibpRYPUdIskMnmjifh7rhTZB
aB/VZkiiInHQscFdUaF/50Y7JUDBM+a4T8n6JWpbkcMa8L9DKll3+n4LfAR3Sxqw
mlGFAicVCc559HKel/VSKZ5TBh4NPr/+IYY2v9vwCjDq5CtcjtqL8M6Jq3SOU/im
2KYjp1gi/nZmKpD2PtTrjfvhuGICsOgUWMRTmoCn1799APIqVSxlPfvk180jC0Y7
55F1ny6nfRI/W0phSjXV/x8KGlg8WGRlkvKgADsa2jbriMZ4td0j7pypAQPhT243
d3LAfJRWr/rd49d3h8WC3TZa4ZNlS7jZXfPrSiHIgM7k9a1EkMkCS1FKk9t48PIV
u04iqRQveoomjE1Jh7DQJbc0Frwrr2vsY0GIZLxaZ0+o7J/uXmAGrIlhoLE9mmYo
WlS0FwZWj7BaSI/qFORgE5hU1K9v0/+dKdca7DqfY0n7SzHAk5QtIduA4XPtefBo
iTTBeISMMH2jSZ2krpVN1lBAZEBzIFm00lLDoTSF6qKjBjwLEI1gGhQatWBasFAK
HogBfC80afgmM58/zIPPuw3ud5DxMLleH4SKqZzjiU1gOTplz9keLVOLLcaHTptn
MyjNLWkXdp40Lu07h1CjhP3VNS2+yrMI4l4152TXIHrvZ7ffuQNQBvocIvmlnVO6
aG37HLrsTbmle/QsTMoiYPTU/EJm1gfbM8Jd16fPbjn92akJ0lHS0blxEwmoIeV1
aOMQDWxa5X1pMqsEAlnGtW0Y/xJjK4Z4i+HvfHE3yFS5m8XwxaSMyCoi4lp52O0c
OFXjBaCWTgs2yJ0KfP2eyR6VYfQ70j4Gp5YXrUkBhAyhB9S9DdAlKOF+ujWhA2O+
uksaiEI0sP1Kg0YOHxuAqJlIps+3j3l0UqmklBeasDp7yS1X1sXFKOvu9bKNM5Mc
T5zHVW1qEzhMZAGy8nZFBNHSUdL8BlB5pKqeLx0haZrJYAJ/8k+eWrSeqZsezOn2
A4QgA4ITyGe6WzvmaJcGF9AA/K3Bf1+lvZR8mj872dZxEtGESc9vkuO4n5fG/edr
IdY8Z7lOBDh2PzvMNC7PvaUFDFPXvOJRX9/SkNE8TE+YpO1kCzuZ5SY8PfNjwTIk
lLaxXwuE64WRc+oBSKAkdBK90YLQ18JyExNkFBW765pH/67DtRJKdhXbpUc78HKT
HA73D7XAvSAX8p2FSdNaSXUbXNRGPGiaJhvnjzA+6TbrgZN8+sdq5NqvdLWBQSEQ
ragMReYxKoomZ6d1K1hpNcbwb8duVCjcny7vjmkljTZ1lxiv4iketmZRIg8HqJh6
w7lYS5E0d1SApAZ9HL5Y8fxDaFcDAFeseEsmNC11LpstkG29os+0eJz3k60u9YfD
2J3SQiqATWyqwwoSJH2otsMPa0hHPVCI51K5M7W9MgDSQKzTh7gaIbrJ5c7YgrKf
4TMRQ7GYk8pBEE1YEIbmgJmIA21cEzwuASDqlKRo6dXHiD4DIjH4bWW1gKUnFbXT
6veS0XFvm6fCZIxf8FL4i0gdUowv27s2DfMBdpAc+lTsW9OJFoTiQISOmsz5+tZE
Czqv1uTnCztIqQk0u4TVEnPcQ5Vs6dnCrLVPPtDFKp0YZQ2ybmMzH90/UQHPbvlt
48WhCC/DFtIDMC51UfWxX70VRJxyfWRErnjIS7FdM4JY85lPfhejuI9uhoXuOgyX
MPBMkdteNN3EKF67FWyrq17Du2HGF/Pp2vT0pX6nZ0tSIQLTek6CJQmM5awhxs/9
QEtELUPOF1ayl96XiKUYbktUEF+pAyqac5OQSBs+3jEP6w2PFZgSFxJkgXR4BXiT
jihmUNbp9+5MBY066Ozi/r7nP+aQcD8DyDJO18Zfo0xVyM90MHjWKuVw8g+WlnIT
XUTHvqksBXv49R0fcE00sSNE1lV/9wlzVwUl66nVOLSYyR4wYKM9dFil41AhKTF0
S2InqLwHuQmNTR2jrRnSc0ifsth4o3mcINo7YWOp5Ie5zbuhUSOhCzFZ3Eo+rXvP
r+VphDpOGv6pU219uMDD7rh8tSHEiHDMuqqDT2kX0lYLLUNrtt4Nvy1qjWOgkvQh
grfSUpgaktS8O9BftLZXheqgFLR60OF+H3vvAeQN5kqwtCiEGfSdUZnwn/6WotMr
Ko7ECkZDu3aEzXnsDJFITNPs7/UGcGpCT7p7G7Mip/nKG1JUpmAm7ANfa3D4q5b9
sjECw4WYeyh91p8A5D6KImd5LGMVVyv5GEadCBNjWFTSf6Mx9iM8vzZmpdagu8NQ
dZ45k0dUOFaG/EHD04yu80Zf6wVwE9Ag4tGJkyQK6VuH9Bv2rXxcjUAAhaHMeZ7F
q3rqqrb4kAK1LPNvnuBeM66l5evqlpTKKVzyHHreNl/tq2d5WimrgVwungUrRykR
vFu1ywbyCOjL9gs2st0z8BNWHKQoUPbZicPxJXSA1UJGjxHym6OCRwkFocwfcCTd
QwIDMjgCItEaDMBzOcH5KdEsniLMg1ib4rh8UUcSGPPam6/p4/D4z5e5ElZfWV+r
CxDsSweIQF7OjuNQaZWS4M9gaaVzVJePJ22AWot3X4/M6QZLedFQydZ5GO30NeDP
Jy/hbfDnD6w+WiQeDi2o9PaReLaZqpnnrW/cEdM59oMOUaQpWoIJOH5rqFZY4q9Q
ZzYc5lUs9iB4+L7+Uc/Qp2ogdQ40uPD+hKzC0mMkBcJ2ynZ5Esv590rUo41sKjRt
jtbL/dYRZ9m1aXqYnP0Skp0o5Ggl41tUSb9u5lMVLRqCvOpUbG9JxYH8BHp81py4
zR9ef0ML+LTYwPXGxhpMUdJl4RuH9DjoDJO4itG9O9Pc+hPeEhJHh5UdfcxxI5QC
6FjOa5iPO47thW7hDKPs8Q+A3g7Xq4dPd0FaUpbZ3Unu7EBvkHbVr2j4OSKDPM6V
fxmfhrPb1nlBZcK8IQeHZ0kUT57zcOgIqNPInW9Ich0ojRdhetoQ8WyiWVDn80AQ
rD0azQqMwkARaH4mfvbEfRIe5HQu4Jr4R11FqNpth2MGtcF2/GJf/whumXIHJtp8
zmzKwoRC5QTHtc0MSFPtx6YKnBXAY5wqeOD4F2gVjh2liIeAEYjjOp48qU4Ols/L
hLPueY7KScfI44nF0B2gluuGB7iZ5c7ZGlO9atbfCb7XlqluGtZ/3b+T/dw5W2Ts
MlBKUi9k3mtpgfmVpWtxMiP3B+GmzPBmvL+KZesTXujnm7XXX0Sj0fr3+ydLrCPt
JKskXnVoZIu8KQvM5mJn1Zq2mLxDdKVEvvhN51/GXL7dSFaPfhgZPuV5xBAO+Alz
0QfpaEwzFBJwOZuW4R8RcHKwuLS7erIMy4sicsCDbJ3Z9R2snKqWUZNAmnh4vSQM
C+MADbfusA9UJKdqBnY0pti7/0nWW9jrKCINeb3KaZ4YdZU+vwk5JkFBI1D4yUcf
Rd68hD+GJh3Ewn2JTmS1kl/+R3jgq8+peEARWai2Ykt/HA1IXdzUX8CLQdz/QwiB
54Ronrs+rVVBZzH0mXEKVop5UkRPNF4i71/L4Hmwy0/43h9qvWHpU57m+t2hwBbA
Q2/YNvO1LVP4AgwGz+VS0UkIunKj2+iDMXj+cFq7ap+khhW21zAzaTO+hRSjlBtU
vZqvhyuAWswJ0XuGTAUHecpSsyecNVuTUge6kG6gj4K5Mw7f9JYDaSEL6piBlws2
sCyXBstHERjCJHr10nSQcP58kcVAY90IL5ptIZ9TSNstB9R9j0fLHeGdhgM3hD7Y
SsGXwfJLmUZ2Jb9rss+guETNUoZM+kj6nZiMRX/XsbWaRZJTTaPX5aTzxgvw3cn0
mwGEfvjUUh/K/seMcRbkQiDGtiau+NqqDqZ7RMdlowvBf4wG0ZhCebDaUL00vRR7
MqNrIpLfgH9SKdGCN3JD578zW3M/SkVdBprzOZEcvHuqkS3gpusX1ybGzwwSMd7M
NAD4RuIeovuIf6g+dRyHDaZYKuXYuvGWswMuoWmkNIRJT8hsCrThM/pdEoicGJhV
lzPb1rmkaI3dsyRGNLe4MX8v1RwPJYVQbv6A1Revnq5VsUScZ0YIDAQx+3l0WfeZ
bOomM/cxVK4gxr7pJJCaoFCkz7M9wU9hR5bpYBhyVv1qQEFkuI1lV4ojN6Mwuhi4
DfvbprQSdbm8skfRMNZ/kLABWL87IKJmqE8n2J2tHbWY+0TWySxGqT5RyZELVmZj
0rNnnTgLHWnK8CIVtyzdR+HtJ7oFNHzSwfiZsPM1QPR3A+tDXcVDRz3cT4iJMZKh
2997EUraf5sTAXIU21M4SicbJeNr990SeRR3VgGAFkeFB+zkVR218d2auIFfPr2l
e4xZjF27LCmJUw69IUwwtolm7W6QOWoMKWOGuzxMYv3DLIrQnn84k2+TkllICHsG
YwLLJcMvZFUe1MaYJ2I2Ttg3exrQWblU0gcJcd/eJ09ee9q09ayAC8irpiQoMyzo
dd7WtiSV7kzpWCt0KQ/bd5Jl2wGCZkaY9mQx37xW9y5MF9KK6EBmr1GM6aKkPiBQ
sFlljpCO4w/P18m2ypNwwsv+jlF6ckRKNjy758QwF2EVUPiksAYFFA8WxJO6J+px
dtoOZ4RwjJqz2Q1gGR68Q2q8qf4qW3XeD7C8KuVpE/Jf1CnNNVhyqqr2qgOrGxOz
43TSn4cU2Vr1wNLFBOpawbEu59s6zU8PbDc7oq5NTmKijmJo+LIXvExwwJf9d08q
g4KSuiFwHVYpdaKHgfLlcnUu5g2l+/afVbzrgzjKiRghqVrwT2RTK1+JYc+vMo+e
5DoLh5WcMviSXYNjvAm1sIeiIWxnA7AktFsNPqRJk4aoPfSnfuQS4YAa+1Hmze+5
mKcoKWDha2KPSiPeZZVn7xr3lFjp86tgTiNVQHYH+j83YCvM0oU+ch4FvAqvrYUX
k2uig6hjLbmd/pvBduV3rLOzydQdFffD7jAxjGRemVuef1t4BmK99BeiPe8i1kDP
M2OS+ln8AmSaz7ztMLjPKcUfzsHsKW39K3BxNTHu1K8Q6VS2E8/pFCe788MpT45/
/ppxDPRWjSNGrgdG0TApsHK8RK/itEjlELfHdbo6kMWQvgnGbsjOJ7Qw/BDyl+Tk
Af0OZyWgdtErop48YR9m3xgS6hEyrlgOuiD2wq90i4PwHHYbqrQa3kEap6EcVdt2
/pkBE+Iy4R9+PjAXsvkpfDSwfjs2zEPTLdEcZvoyjju+WNUioNnMMowdWHzoKHL5
FTaw5drQzzw7iKj99eiyFNDbj0sGktdx4jGFdlTcjZSEfUHFLK6bd48AIxFzWI19
5ogsokXYkoCYlpE8HUo90A147ixxdfjD9z3RKze1cMXCa1kpimN0iSm4QSs6qe4V
6GdQxoqDYF70hV+TmNKiIcCCJLTZvY+BGZNidbq+ZjWVMi1pQTpNIPzT8v3M9HIU
TChRUQDgLamzPAVd4Fs+nxd3djnJzJ1i2wCyVQ5L8Kmi3hkNHRJWJsGgOCGwImqX
jR24mZuSZfALKLCf84CgeiKgB+njPtdB6bW+Vq6dtq1EXt2jazyt+/CsCjStAsKN
Nem0ZKJzkWTkq1uHUW674ROF2/TKJC8GVEvGOKjq+/3ccPT17DfXArk25ZbiNY7P
gz/nCkRrUaLNSsGj9x30JM8JgeXOSAqU3VSy+hlGo9y/b9REFmZSCHACynee3j/D
m24DNuqV3dWgLHtkeF1CkMEXIJ2ltuhzEVrqXl2lp7quX9UnsqCs93beR104jDFt
s3C07+FOj1N1K02g9LdwP2Xechnm3g5AKkgqnmIgQ6pZuz6Ek/ymTXLgJAl2PdVY
qjOnSZIombMrcjNQ0SoIjojlBABDB6+zW9YTqD2GPv+bO256ZqZcT/vXm6P/Ew8e
vikSmIwyVkwirbU6p/Yn3XL7fVvM9L6J9D33lc5Fvowjm03ToQYFJtVRiItvsmYS
s0Y/tmjni390EHNCgZz2n1PtNCD165P3f8/drTyBPOvXe05C3Ue9YC4U9qmbsrbD
QwTwNnidQ8pKw8NvvXxEmnQTwAH/QkVLVwXUC6TnB5GA7/JivtLlV2WPjD6IZZiG
JRVb6dACWw+WXmb7q6zx1ApA+gvoW/4FU/0Xvkikcj92GnhXxmrxm1GCbauWC1ac
D0ma42t4c8qcWoyEXtxhJsH8Aw8MTgTfZaXd++dqJooUmBN+bzj2Pq+yaGlmhAl2
kDQ28msDmbV4Km/tY2Xxn7gZDEDqXtRj+sCqQ8Lxi+vxYG1QOGh4MBC+ASR1fuUt
hzjzVpe0h4cbl3AmgeOVOZCnxTzKyff3OULyPI7PUf69zCEyCXvS7iowxuGDlcEO
GLHH35DPH33EE9/3uXFWqhxrycihbrFdm2z3d7wtYyC419xGZZX2pOU0y8JFlm5I
7ElhsFtqFL1llerNXYToj4jDtHCGzGHH5/5EfrzRguzyiDWLhdUG+VlkAfdjfTdd
bCXuzfmhzSNTyRej6oKVIIO2lcetv2jAMKeLHfRu2TmiNIISJ6NoPokTLvKxYmq/
jDrFYiFRpc+ocvBQHjoykFAkv0x7piQDPQyVLkEFt/CESdNoQuQCU+ku8WkH45GH
ewfnx6x/+k2wK9MIJAzLhhc5kcTV4+vqYQQuLFF5t/glia9lqBAqz9PhjfmjGifi
9B9HL2T68ryw8DxzgzGs+Vtky3HjolrtLMdwk0D5+QHZu5Dlv5ZeWKVuYkmAk42z
bnZRaFbrn8lojTVBm4TkH5n8faGKU++9ZG4DTH7bZG6cynHF1Wim+ZiEoOOiJFpt
FlmtH+Bh4zHqDjiO0BKOaw51l2AqGRUOQ5p/y9RDu37wRDXStg+aPoRS2ORJb49r
tzbtVDo1UdoKfUXVIu860pkzRJ7yQH7dcrvXfjojw/Kwpw0Wu5I5WfFal5UhnbUE
+opHwJZNKiM2eEvUBRcyRaBDX2rrtHYDzR800LYyiWYvooR9ncBK0FY1bTf+HU0J
nvyR6wOtI4GxQqWZlPN4KUG+88/Jt/NGVOPPVJEKnpH3V+r4agXO7aY0TovXt/Cv
aRi4v0CCwRohTJNYN5ggcq7SGzVzmAMy4brEtX7ugldFAEpe38j4XpD3suOmHrh2
uugBRjtqfLYyDyVJ66mOZWcfh6gsmWKOs7YY03Y30oUexEksJk5UrHqeRqNUTGNP
HptiTE1uO4GOVFvxQqj0DmQ8CNxmDkl4J9V+jDIOdFtSxtl6r4pgtFf9twT7utJs
8T4ZYUDVd8PU30ILWtRyTdNGUwxB2ynwuY628CsJtgvwBvisj/y1TVLflQVCfE7d
OGbniwuCDUdn74HalgFIKdWULBiKD1eQnXo+b5B/d3M2KF0iUXPQYA89VJyopsCl
m4ONIcVx2zMbXK0a/sPiUXJnxzN+nKHzfN1lPXFojX/HRPZ1spLAdihWF0Y/aRPt
stlX+NSYvloIoS+HdahwikW/kkq3BZYpVfjT2vOetK0QSSiroENYZKkFxsNpfkUZ
b8prjksh8zCPwZ2x6Dq0cB3dzU0yk2YRNP2v36hHhphqh1TK8UgTFKthIZB5BGN9
E55lMlaBSFveIGDaPEtKm09++ZEobWpiz0zqZe09lbSjxZet1qbnI48CdHANwUlS
W/hnTsoBgW2FBpw2DuGw0ZHvhtiZObBGt1/yg5O9vvehoEo+iYmdX2R7SLCEKO1g
z/p27m3Yao0q0xlgyAGBlZ79q1xAcOSNmS1TeknU1bBxfI+np9TrHv6zf6Oh9WnI
SxfZ7XELHFvN48KyGJkoWOtkdh/71Jiph43UEjIiYLgBy4g/lnuC4EehzcDYoTBu
sSWa1aNEmkCyKBKfwSMiSXlMn98NUggoIeMgzQ/IhKPcxj8jArLr55KFUpmTxfUd
A0eXytTNO577Rka4/Vmd/GzqgLWC4wZxZU0aEk/CHhg4zRUi26+vp2X9AY5mUAnb
xJlt9nPS82YY26Iddt+kL7mXSPICRAkaY+qLjds3Dn3emrSRy60byOQKf1x7dB04
z+MBJrRRA91hvAEuKTkdhSU89LCXpZSVobgZOu1SWuWzimAwV4E+zOHRsG9M3MAA
eTjU/qQuQ3YfTRTb3lbXj1UGhVa81WvC8Np04PWHQu+MRn3/KzZK+4A9byFMCRwZ
who1LKZtBKeXiUXD8OWr2C4F95/uoPmUsQOoLVz46HVwOhR8lRxXz2Injc6AVbFE
3S12MglUtMp1D+1dMhhef6fuqwxgnlfuEsqrUYiQEMERN3ku8Wrhg1HgtlcFU9GM
qcPM+a/bqdzcA6hVJ2G1qHsYQ4PTa55aIo4f1/ItM/+dgBX2x/ReKA6yCW5J2SQQ
IbJjmC7ZGEk4iAgHnq46R3qqMoBaT9daJhL/oE3hTEw89tyR/k/f8tjzUXWGRaqB
N/SB+uqt4rUVJo1y862ciI5ZBNoJWMrRr0voMkvdNpazOBlOjyrtEgs6qcm/pFLy
xVJnNLAngIU63EOlf/TgpkW/69AnVDe8jTlowYJONck5S/7MCnXC3R4TYritMWgy
YTdnenWcq7JmFfJ6snswetIds++OmVWi6d+tnJram2LZ+kbqnaBCj17oNs1M2rPU
CshjMe1tKfHlbD9dXi2NBKu/5+kbmkCT/gvLgHzTd5WFy0G+krBvjfMPkEHx+R5n
yU5rtwREuV20HqFPYfQwH1+aaZXC1ULPEMl4GORmSVPkrNy9zlIoTTMJVG02AvRc
apNNgG+FblbA8lkCRl3OorISJ+zsH5tYiALnoVIJthYA6fBHQ3QQUwBl83Ma73B4
iZ/3lwJBrwPnk4Avmh3zS+HExi5xqozVPDv7cvSG7BOCTVvp+ddrnfBOHdOIT0FT
uyMUuwpVxDw/F95THR+EiRxu9DmaShiqulR8B6BsSy68IEgDHmtei8U3/ZTz1oL4
8dZA6SQB6KeYk4OfEIT9uOfXH85AV9sjH3/FF9xC2bu+VG6QCTpQevdlD5hPAG7G
H6PaMWnW8R8Yu38qQuFIGtl//AXaRjAaiDOQLb3cda4NzuiPKMUETyQ/LbeFNLyD
EU1AXLjhnTszHJCBI3/v2fsGq/YbogtXrHVo1k+umyXHiz5hls229mwA2kmON7wh
JngOlVPx+W7gqytNfjkpZFZDgke2uG1kwis8Diz0m9VyK/bGjHXn5P2XCC2zgH4G
uU0t8nVGEsWpsEcWXU8PdpN67htWOFtWG4+mdfgQviYZAijEytQ16YWsJ4hzFy2f
nvYD/kQSN8glwb7XEfhwpXzkVYS7Sx0D7ahpmTMbk+rTkOQnE/WnWEQ2FxPlttZM
gbbftulkgfGT11vaXMImrqsPoaJ9FrZPOEKEHUluahN/doHsHVEuypjqJGeALJ4c
fRQTm5NXffqveiBbtvUhidQD45+ZOZYsqSFvwiDSUj/Po2doHLfFi2iZMHfQzCcL
7444I+3s3F/saBjPc8g0ZN0g/J20IeLmLLxjyxSt7gazKmgjNw0H2Dp6RlOcdDQK
YlcY6d0Wa2mtTRNb+I9xUxVsmby4EYj4gZ1+mySJzBlymKXvXat5uvBuc2f/ml2g
0Zpk73J05jPm8XT7zmICN7tAQkieUx6aJa5rOtAat4DDsBwiMgaHZQkUAa+iwcjU
LVVMaOubKPjJwN5HJmyPOh3f/J/NiS7U/gsX8ImuBx1RDMjt3Wmi71wckLpyNuqi
VG8rfHY2nZs8Qd3peMa5xG9ZiqFIzCRPtduExa9vp8FVncBj4MbysgzPFMmuaYJy
TfqXz5sF/KimqXZeeMyp4v0E6AVhLZ3P9XRkVJAaNaRGLoQn5yiISm9UBU15GYLW
5IpzLyM/J7zPHjhCyj935M48q/QqWBzZlWpNZiL8jDODFntWQ3iszrAVUaPQOa5V
SZfPv2GslFmi6s3GRoGxBDIL9I95ceYqZnvbBvuOBhHAueuOTsYd1IsJbmmm6YME
0nvzH47/hTRRNV1isvVYsDpxN03KDHPWr/bDj/hF6beTY9HLhVHO7nmT/jObNhK8
2D+UFfeoMFlBFqaxvJK9jWSSiPEtf8cKiFCL7RkgopY38eIFRZ1bezlUu087floQ
q+n+Gw0cEHyHdbTWTlZZnbpxgHfg/VQtbe6qbSUav/m0qqFgjnIjJAwR3X0IN6Jc
E20+6B4u5+Dgfv8ujiXwx14AT5fBbinbtkECLWvE9TP4fyoSAqg1fXAoeEGHJhcN
ZDBLCIlM3YaxgDp9HmZrH+CeTRXfhCkp4I16t6E7LsM2kJvYVR28nftU4+h57F3O
p7zezfuyHdewyz60eWMb6eu7S/pyAfvwbMJi+Ri8RmQ9dnP7X8RnNY7Dq0VEf65L
z+jM6VqhTiV4L2pmaSJliIVldQtvu6qzN+0yH/bSTQHwitCW5HG9qev8ut+LbID/
3l/6qpph/OREIazoTuaBFh0d2RFV/CkaL4JCVVxA0l3LJkCZjMthJ7vJN59p4d4w
0JRul9KLho3Xf5R/zXGcrnHlGq++7QGBPgzf3qQ6cauTmivS/yXGLXXfxcE8mn2S
xStQWrVH1D/CxT7bK6PxEKfjp7DwvHPhgjZSASOABxUvpnnOz9IIgOwGPFk6UVuq
sAZT4SiBn9dWAoqSgD2M/rfM2lnxFMDUx2K0SejUzKcQTdc9mI6wiEg4ztOxM+nv
MDkORn7pFgJG/vVqOza3/6YPXNrlmX9iq9OTEBND9tyJxYaDtZ+SOu6sNEBwjPxv
R7YYLbduLXZe4k4ZQB3JT8i5XMKRxz83ZSIrXO8yVv33ECLYwwQ3woar95nNGzQ6
i9zDGFjPKl9Py8fHgcXxm5sEYO9wmVTBZpbowEaX/Rz4M4nGzeKe+84zgiKG4p+/
FUj42b5YjxfXIuBSJpnTVdeLWwDBXCkRi6tV1Qp6t6aqeluwi72d2gYgmLg8iWTX
hKGP7pRRwiRHWq+zWMpqCY90wLMnLQ0j9V4RsVLdUihNqFEr0+b6HmnPTZT+atuZ
Lyev65Czlia0LXg80HN3Np8hqYx1fZ9GBhpY2ghMLzAgzkpk3oma/YEY82q01Um4
DXSfrwm3f0EaskRgvrMv7gz1Vuc5lADO6sD70JLaZelI9LbOA2moTEppNgRvcJaJ
E3AFzhpr6KeUHGuzMpfqj2kawVJDnw9uD4qu8LV5p0jt7OJ46wqGZAgogl0bikhb
G4P/S6aIX3FgpbYeRwGH+06FzZlV//qJ4bH15cXAShb9VPGfR87O5/loOa6i+V81
EunP/ncuXgplpNObOwwVmQNckl+JRxl9vPxMx7VOp27hfh93QsA+oPI9onY/84BZ
6Y0qV+O9zEjMxBdBBHd8S3hkUtXusdKp+7nHl+5oYDr0zoFFqoAkTeuMz3v61FkD
2OdvqgoR4IyllR5/P7vF5gLrqb8COy2PhI3HI8vDlC2/j2grDCgF+1y0UGc04SvV
sbB/V58GwwsFhKRYKKw52TlMiI0DQmYtPMbL7kekpgUbIf3dky1DbBk9Q+92qZ9+
Nb5CNhxAO10O+4ahXof1Y8uz02gD8eACjrrUTQTIWTpbrzG3GUoTg+LME4H1SnUC
jszxm8q8yM8LksWZYfoJOtPHDu1770TRHjxeqW1z5/mhhboAbGEWdcs6XzYAJq4V
rU8oRUS+n8GOI3vRIxPF+PXEIrryVGdEVDHFedadudSxClcCUBOmITLM0BJNT6W4
xvtK02cVgWAPENL/41Sshcy5U00G8EpRMqeET7kQZQYG6s3BoplwacP1PpeIyx+T
avTKT/+EofvEeNbS9pGT4A2ZVIfIZ/8kxARszTAFBCKygzK7yPsUPnROY4KVWsf/
hZmKmS8M0gzddlymfrwKS/gAqQ2cohetjxZDRYDEAEJgRNJPtQcT5z7X/QB67uuJ
WwyDLi3xXFwhv6VV94XgDtzfnbn44i1XegSy/jzFPgC+D97E7ec7539LkLbRS7K0
LewKiXzn85BH4D+Bj7ZBE0jytZ6yaaz8hsp6CHfCTIUTZsDCkYj5bJ0hqWV2p2nH
Dgoon+WLhgYWrPB7Rgh1KEt7wa7lpXMQ3+nkH43aqqv/dzBjP0amYDfHWuc4xoQW
W+zM3Jq9dqz2TpJdAwYrxA4iOpsMa9oLtmF3xgTnP+dtdL1HrKBhtEfaHGGTpsjA
BzjLpsU/wjx1MLxN6nMcidf7xGZ1ntnvi2Iic0pFfctCb327ZK07PJisDLuJKzHj
IVm+CpcWbqO+sMas2mzmjuIiXpJZWyV1/6vA7v/9Cw32lbNR3ekJHhtGP/42HVqH
+e+8kCsB3lOXg22yGQJat0oZub0lgoOgPbpIC3CjBZ7ljH93+6wKfyYuAt7lBhgv
pxgbhfS54YSvGpkmE4AxoNAXl6yUYLbGoXmFIbyQeLiBOYkg5CQxjsN7oddJiJ7G
3kYmWEY0PvsZ79O7QJqHD8Ngea9MKXaCNb0U5ZVKJJ3EtSbYpOjiiJjkPTCOgkU+
s7y5KVa4wXWG8O4OYIg7JrEDjShBnKwXhgmoRlXhnWnAkQhHEhN0ExpNyp9NeMYr
mQVsNLK1gKt8b82dSVfOn/IEkZfZaQJCZ2Y4x9VvfQs+DzFkADJJEOB1TL7+MXr6
ErKh5NACsj4omyrQh8IkroQbPla4j3lJY/6hbRXiPPTbrfwLPfXUrSxOOI7ShQ8d
88pVoUPlg64az/4nwQ33f33Eoj/+v7yxMVwt6xS7rJfUtS4/OFSWzRW0FkUiR1fV
v9bieCpFk6nD5b//mpZrNNYZepmxEuv4X2fwqTZISAL8/R1ivr4/ZZYw1uza/gHM
lSGQzAwj1voJZdmEFK+kF2vWaLau5yZqbUy/K/FEFCfILjaG1YKRps1Fp00o8i1x
yjlkk7UfPYZLFI47OH6T1nnDoN63++5OxUOC573Ut/FwWNlrUpptZH37fgHSW3/U
o8LywH2RBHzibC3AQolHBOlzLE+XDUrqmgYOpgo+xQXkFeelTVEiJKfx12jaby5b
/lobyIQwW75c9XoHBp4kgVd9IXhbzYZukLDb3OLbMbWd4xFH2SjT+VduHZZEZicr
qZtR35Ocda2ybRlBh6g51laxQGUwyX3AeOQ/Eik+C6pyyxtRFawGuekKYsrIehV6
ATOmZXJuLQjzqaX3dffmM60niZkGSD5H957SiDz8jvl3gjKjhby8b5D1ZhQLTIc7
SjAfBDDikdUjvjmj+AWhFNJrvzpWIFGJaUW7VNdzu2umIkcV/Gk8ETaqhBkgbMGD
AKPNoneb6S9SfcanTNLGxhAzWwHlb6g4OMBpZQ/xOQEw2djKeYVPp1rki2jtStVK
oC2e/A5gNZCP7XhWB2sTWZr6isiuJ3tHr0evBAUAFAmp/IO2fkEpO7Bw9lKFAT+N
AcvPyiTj/2cpkwIE7goiRBhKkI+NetyvYO+Q/ToTkZNNsKU2lb2D4b+qfrSdgb0h
RNn9qgO6VO5smZv+tvaBkOzhM1fJ4qr681Z6qjchvU1j2VYiVsIgRK1CfRJpgQzj
YFDgZGXKSLNu3K1dkiDpOtA6Uz7xbjDnr0MeUR4HoCDnSai04xYxy7uXo2zwyW1Z
r9Q+4h2a8Q/G8cUAQ5vEgAnOlCQnmL1KEifiJ5Rvydxp/z14TCAm99uFMVfvD0VB
hQk7TtmSLauGQA0qnt9bfedOJZPhmdkwSW+sYEIyhlK4wKr3XpEFlK5z8Y1daFX5
jYtd0LUkeSrgUs+F6od2EQk9I7qDFkfz0oT3hmbH4uzdUnqCc9LcH3TWuKynjYMF
Ob1GnPf+Tj6NXc/tNcFki7p9IQx6Ik7bXfUzTqbSV0V3kWCFTJBHaJDuFryWThv4
jA0VLnCqZr0FX66UC+o1fMgLZxoY+RxENbgT8RPan7ZVK6h2TxANvML8d7qPaDsE
NFcYjhoeYdEXthNRTq2FGAvUyLe13NckItm82VHvkes3eKgWtfGh0RuxiuA0yIQG
BDxp5YLMiWhQawT2VnkCtwqe5Ughyo3tqtCNfzyk4cDdpPRg6YCz6jETcQOg19/J
prnWTvv7YG4RrLwE0c/Fm1GQTgYcUnGPzUYtpuFNUPs4FS8+hCJ04CRFVvamdc0x
xQDCpqov2vjrK1IzSLRUxHKKPCnH2D81L304VAFg20sguZRCaiSxeQ1QQZS6CK0S
d3mzELyaN0DwOfVZiLKYo1kyzz33C4OBzryRoig0OFY24DqJ+lxJAXz1n1lMPd4V
SzysEs7XJ2EfNhKcmgA6bZyDmmfPqlYhyL2WBvWLYI0NxYUFxGQEISNeNvTkjzFS
BjnL5gEVASRbnMjJuE4bb2F2TOBHCnlpAG8cfwgXcGlql7kOYqQjz00FbzbV04Ur
iKlRdDLWafJ/i3iPB77X8SRZuZQB56TQXlQQnJVlstdgjABKnQBNDKx6gB/tTEEY
NPZLNkSSAFLoilwtqHBKfxfKqHGDqgQRiF+hW9/iEnan9XDiaU+RKGlgw5yuUhwI
zy7/ZwZBz/3iwO4SNgsijbdVqlH8/yr+H9fe6HFybmMjVg2HeRIljG7kx8UtNv/5
KXBbrESz7sns+QraaL2KDsWIEAQ7Ae4tByIXelbvDBL4yRcV0kjZkU/xw8lKOQid
4KCRmy37hT+vb8DizX/OWhU3vP/SMYY7Gnx7nDKnP5uaGfLLBEgdJuRllZknIqER
oxayFe79rHClMLC3Yax/7bbBlXAkZSeOUOaepCi9UCZ/nm9b0U/CRSx0E9vHMbI7
4T9HonsdBusW2dXDPInh6KdWit6W/EcA/0IERd/aqP1R3miAYt27qzOe2F1ARGOJ
vZ+0SUhuraIgrPAO0U3bVtgRqOFYyi75to+dMDeqe3+0rtxytUISp0h8PFlO7XJC
wYILwFLeM0q4Fx84pa1SeSXPlkModbLzM6wTBPBWNl9PrdCo7+vc/FrUHndc44jV
OK8cUf7d6F8ZCc1ug3Fu3q/wnvlmiPQW2b24jqzNKdT9dq4f4rPhmwOat8J8Nm0V
D+xBrMFG2V96YgjfXrow2mqQSVMNyV2rZ5bCu10DJ8AkXgVjh5O8y4hb/yR5uDvV
/3gVSKFBFi88Yw9TFoilZm0Ry4apKT52PCDRloN2t0DXLzIIujjtmXBMP3xQfMQz
KzmX1A4ALqK7lhX5xZdck8EKOBcLIP1kJfQCycN4E39Nn5LiG+0slv3PjL9Oluyq
Da1d45etiIC8bTh3GY2n71dEh+LDwtG35xI32dp/Neup5BAjQNmRLkGFCwQdPvYD
wlJ4QZ0WQKbciRqnGrhT2uV01VzYOUEzWqVosC8e7Og8lMqEkRwgonqLEMPnQq/q
Ai6ZCZn+VolR5HBTjRzy+VuEySKp9m0xrnYlPNC2vZtb+xm+Fz5XfpMq+CmJnz42
fEu/vZueRUMOH7ZeZOKOL6Cmz6ESuPWzmQsg1SRwCy0olLtZFMZh1oc/AQBVlTB0
9BhfF0NYlpM51ZR2hk7Vi4rwQP2KfXQQIex4rtWKQsVXNPx2pMtf17ynPouCxBlU
7McfbLTptYITiXrEJq3nCD4FdiRz9Uo8rkxJ07Kkn80D97BtPxRSIs9yOTYiouED
eV2jM4xLO6750+J+fO6ntTqKoS715qY8GDDriVQUBECWAW4l1yLrgyBPz4aDvALC
UzRVRyVaUvSahqIE+VoZJA51SrDeMiS9gNsmOtOZpBkhHGDhvNUMZ0UUJoJv9/jP
BBeN83Ue5LjtVqHvOlfM9Jq04xtDUtwhFv8AzDUr9sFLLlO8YA3bx3xcJoYK2NFs
wpCA8y9K+D4KXji7SU/Jq5f769+67zilwLsG0UELbXQe6Bvlopu4dq9InI2kO+fL
blf/gJzfZ59iE0thFFhYUVLf62GeCuUOmzgC+IcnsFjrpFK4t4R/D5PS8ZxfVYdj
zMQbrwnauK+4wk/eaZ2C3Dm6MtUaOQu9EgtKu30vUGfDWx5fezpYr8y6Lx2YJ7/H
UMV6ejI2hkfsYqztwM98itEqAOYspA8A3Pv0eMnx2oUfKqQW5DpfzXz8/umTNu6z
6RwIlZF4SvebBzsWizOLDi5B9tt2Ue2UsdpnTTxjeZSmEiDF8pcIWuP6Fr+nJG1D
nOOj+w/tj1CJnZn6Y+lxc4xBuXBDZiRM5jXlUAD5dtBy2VUv5+pb924Z6QvyEpjW
6LQoT9v9nFHGPuKF4FL631vQbaRZicMuhcGLLfGVjhufw0ojgdCtYNpAXjA37WRg
4GQOpXp6DNArIQ55PRnJGfyXtP7sNEaMZRrulxj4pJhbVsp9r+p2+71WLG40C1EH
Yf1cN3dqe/qPQ/7CGm+gfOUXImNtcT9Fpdh3S+lLZwx4Pm0OO4A23YZflqrvgxHK
wanNmcCqdyBAH532hUgStTHxrWgZ9s2oqzNyax003tePjuRY89FRFk+G8SM1Dmvn
V4z9qG5cXcZSA39awrLpdFOqmmoL8hEz4DeD1Tczj/u1KR5akxHOfSa29ct3pD+s
oZboyfcp+DFSiS2xacWEuOhrSE1z8tSq+IPXIkhqyRwjZ9ObPL3t00XT2m2cqrsR
GTb8NGAvqFj3JUsRnmIYXA8GRBxPP3YxwRNPa4Yalhl4v1vEcJuenBI1U2PqQ0w/
3EGARnhKDl2fmWNF+Fj4t6H4uy8uXO2Va7bJblUsaDNycxggSmTmvTt0Zj9ulVGC
ZzxvBZOXlI7wSpsBINaPc0foOJVQKXZrLq5sTA38bejYSQfTaGnt2SYqBJCQwKP5
GG2xkwZhwBhc6JIavtpv3IdFWTdtWU3MgNG5cJRooBfRn4pggfyHIZk474Vyitw7
MTOeIyKyLyrocZ6kFhXtJHFYgHpEmtB84lkQ/1SXeO4KgxCvHxaodAejhCV7Lg6r
jzfmPo8BzVyiOahhJHSQ/yROMlQaArdEcUh2ZOSDOqr/8R247Dp0/fXbj/2mFCQW
0Lr0Hy9LuFppNeZgxeTwjKWzZfhbLxgmCLAZmxUgBXLhV/TBirAdZEIrYr1ArLbT
PZY6MfPU5zKLT779n5/jPpC6dJhizQAkB2JVETS3bK2L2vwR+0IE01pFA4qN4Dw5
bYgpqT/l1MKfphgHSSpDOC70fT0z3G6edxhgbqqz7c4DXnizS3Vvk42y3KoibaV5
f+SEqziIM0bG/xaN3MZ+zrfw35PaBZ5+8ws6uZCOnMAP62qZPaXNCqxC1bhFAN8D
4K9SVQQ9A5LqqNTpGgTE2h9HPmGXMphwOljUWfYgv3lNNkkbWqXeG3JB5EZ+JVh2
2pDXMa/vponmvM+SwZ55fMTCjqa7/jWo+bVRv96A4lZ1Uw/lLvnYgw6VNfIlP52H
y/FVjzCAdW07w9kTsbE+EKGfxn6l84/FFBYq2KEvYZHZyNJEu+KBJVr/qtrgq7Sr
6+BIb1VP6QBRb6+m3l5Jep1UZEAvyHLztFFkxzlkkvm8jZwi4Ms7zC1qQd3F+lfB
i+dHUJPtizjKjlCsRG6JvdVqwNY97/GfXBZSMAI3wQqfT9yt33FutsChj7gI7+OB
tEph1NB2CsGMXVxk7kqXELjuSNAXEekYaHO0Wdxry/QdVCRYTHobaQtgkYdYBzJt
1R8sP4XvGaigIK7KRkTf80Yns1H66Sq3/GUdUVQn8QLP+CuGg6Fc2ODu3uiZZ7Vk
Apm3P23JrtVvr24KGzDjYlAyAYKgrj+fJ0tW1+oHO19PPffuA7AN5iNL++xihu45
DgXIMJKW6LXAWWQuee6ODCbpzD4WcW8vGrpSAD6ioQBcOU3SpMTBZQXXHHVZmYHn
qI+wZjwticw24aMYNeCmrnzQ4113jcOW7FrKxB2iLJ4HJB80uRF36TVecKsuIlRV
10ezfeIhExfpJ8jqeDAPaUtWlvalQNf6BtT6q4jTYnM6MbeZUiqVj2KCvDYA0XkN
CwJybdYY57pmQ6MQiQ3IVFF+Fx2HoEfBzIEeBlaUrMTrPaS57YadORn3GKuzaWn3
JTesXoBQ4N+rF2n7FNbRW1FASckc00QLSvTrJw+HLnJzJZ8qvyBTRyCA94ogcAn3
umpTdFhwfyMvkGrMC3JXf8O4/dpy3rFbWfF4vBrvQ/oT8A7Le120QhcI+vfda0qC
EigRubgNfgANQTnoWQOQmc7TGLn0DExLFAlIPFk7wXIs4eq3KPpWyPkv6Ku3A7gQ
kwYOv57FzLkYkd1iMf3ndeUTJqfnKlKP7o163W+5NbwT4L1VtyWhcPHR0cmtzLYB
yn++R0Zfq6InnaAz7+ga1i58yJ1AgxNGs2iI+/ooLaa2rz4+1AfbhJCvZXSitnag
25/cuS1Ei5i+WNALezqNuRTZv+sZTV8sKRE4COtub7vRLhBz+l9wN/sGCMJkvrHa
EVnPI5kv7EBVp6PtgqAm9QWTjCHdiLBqJTFFUtCUEHtHCnOiHBWNPu76IePb7NqI
uNariwVorsHiymwZoe/aJeNFJhYU7iC8JNa1MeNriVrCwrjIY2D4wIlh2T99PQx0
ZOW6o/uHZMXfiaQIq1QInkJMUvNoIDsjr73zu8X3PgA2cMctdNRO0TnI6iyk8DqA
6bVWsAnKYzZuIyayZuroHDUmfxqu8JFWt2YJRJaudmiUni2CSC66Zu1f0bYruQIM
t6g8M8NBXsQLxU/Ep2qGHxGimimfCuDsOxZ++vpp3E/4I7f3DI3k8Q41zHcSNSxg
0V4gGyHJWr0YxucVOPXTfDSXE07Et2JRN0uC49i4qSFniSetTGUZaOGPDjB7fO4g
Gj8w9WR2044lhUYmo7IupApnl9WCwz8yA7/8iLppFJ+NDvrlCCwU38F93HcGAgR1
r5FVbbq5obpmD411+qKCbartRlGqulcCY4QoWghI0CUsRHNyIIsGNYeBfA2ylA0U
Uks+w9omtupgHFZwlKexiRcXMqugxvzLDtiAJD61kKrd8pMeDmM25kC6bkARaXzo
jY2wyFo/S8fGFZjbwG059SawevWRrynB+cP+NtpPtmS1dDnldCgDFsvT6sY+mLwD
0egYHyJernqJk7gvuASdkqi5WeFpvR2wjIuLpWhn4LuoaJFPLJX9/LInDGxGRw2+
rKiGMztvQO5wMdvz4vsSXMVKrPlIvcHruTPGNBMAAFAoPCrBMwRq1crcplsTT12v
HWKW/h0h6RlxqjZr3GtUIft1JVli65V7CmKVh5fsJ72pAmkXax2LibImhZmoRng2
NZ/s1csTf3kaAEnEN0x2O3/8uaJvqxog4Wb0bAmvZQNJDkSGPSIERvCB4sqR6WLD
Whooj8wfRBX2+cNlGemffJqRsU28o2MyoifOcsdBWOixSbFn3P6aM/9P9T7e6cp3
m2oNNowTMArczw8kFA0h4HqNrOy+TB7vhLz1wX2MXQzHoy/rMhINsOJxhrNcCeV1
OhC4ScmRLFRSS5jR4rstnH6re88d8Hq5dBQNXPbK8pgYrfiQVe1L40kyTOmkUj0S
jQ4GPgK4bmIvTzgqzelvUn1/RslTZ1MhP9BA2kDm1rhvAuqa/8J12N6Q+wz7pbc9
Qa2EqDEK9UPCZw5skrw27jzXM3OVVTBULFy5t8Hx5nAenPTkILh81el2g8ZiAldK
eOVTF6fWqZPsgrHP8I92ZA/qOAq5KI1hzh0tttqBobBMHluQSUtdp8FqZxPaFK/K
gPHf+IAtRdLq5SiFtD7PJifQabz0g89ALtmuZYuHuuDJDZm7Dk3I6AbaUe7HMUSD
8yt/Iwpq94ZjfaIzoBTW1Z/kVJWu03Z2UPR3TK15LchCEkV/HHCJSC624hsIPh9D
nGYZNESAhHiTT4RBDTssvLKp0KlNt1E8nEvXQ1pD7OEOFVFVS2al+X4alr4dU4yU
iWHxLojjK7A2enWpNHk3E/uwDz7cBnmLRArfYdR5Mz5TL9sbuF68U4oPJNkCGb86
z5gHfTClt5RY4hMhQ1wxo3TXq1yDITybloL6TBj5Mjhs6azde3jQ0oL8n3/sPRHZ
MTXh+gcVTNW6CH0wAycVUfuK9MqxGLuGUEYQbK69m6KZhjpaXmQq4LRVmdOQ+NI5
v0h+hyJMT4JvFUrecC1bOyYovYvwHxHzayFec+Qazi5+pq+rv1mTcS1TK2tkHFV8
OxLDjCYz9EjxyV4AtZlQOeDDEtjBhvOxiwWoh5QG5oL9TQCKry8lGcSgbzyJICCW
njcmQXPXQZCHA+Gqgb3+TxMyxImf0I4B6phkwupEIbDjVcdkT46zQgTmxseqad5Y
wDP727xrKyUwJMcAaMRSiOXFU1QX3QdkD5fJH66Ug9j4r2IjgL4ciMdq8FuWApDC
NnPVNENIM3CSDDu1RBk1QIbVEM8/gn4EPDIJ2Q4MGMz2G7/NtamPruKIsWSc/gi0
z0gnUcIOnc/lcD6cWj3njT/20qOkok4GynH9FP1Rb7b0ny1ml8A59o6wZNYG1s5F
6FCVPknBaNxozjP/tVCkh4OEArbplJZIxtuYCU7Gz2hVckHf8hnmYExre83fNLHm
7AEBLGL/TfjG4sND7yMC6GUUjltj8F/oUA9XNnJXyTXujx3JL3wvCow2Ngz0y0GO
TtDw8KfH09h6/461ZXyn5npLbze3bxNHj7s2gefGoNS2IxZz1+l56YS3d1TQnsZQ
Z3Fdsl5G5BDMYnCm4jy7XAW+RdaqdGRzr2JuqEnWgFLm7KyYGijcXb/YPArCmfI0
xxE1Es32gO8w+SJVtAmh8xYGLYcqnAeSfaE7RKe1bGxJI9NjV5+gYHurKG/5njME
BJJVEsQEB+T1Z9+urwKmolUdXBhZLlv0uRFZOyK2LHSCMYukzk3oG2xRJ+B4ijnt
1Yf4UcJZP1Eerr+uVCNh4ark0c/+znlZVG+yGX9LFFR5Pc8qrngN5pj2OtMazh7d
2kggMKdrIyMzNATHEtQuSopVA9+FeL25HOk82xN86CJrA1gO3SYjfkE+04l0UhQ4
Av1TuRtY5VJHsDQBLS90yUHYAthZnxLLl5T+KhSRhteez1bgCAdXw+B+TxcpCqnt
FsXDMNfobm0vzg9PsTEXV0cC9WmtX7oj81T7i16svav7/Mhp1iWFTn5059vHo2VX
xvnoZUSeKA+0lHdWNybJVsQEUrivY0kMalVOED95Rk+rvYaxym2JpraTyX+R1ufC
H7+OxbKEHvxg/uu48wiFFVhv+dbSy8H2OJtuzujkP8UfqlxeAxkSljPlSgXEjAQ0
VxmLq9iB+W+SiQUEd6GQo6arfNZ1ZLzl21Qg4fnpCGL4b9pNbJHc2oj9yvHkPF2R
UXLU1cu4zIAidpUhEgB5UwxqCprbPlpHLjbo4yyCzu1Y8GR5n8qDXEzYblJZ+Emh
dHcBJTPJ2MiR5fpqPUMKz0n14wdZI8QApo3VpEddpr5e1B3rGWqUKpjc/c3U8G+g
MlJ8OHqQ9xSV9ecwsVI/qo0B4VqlOM1mP66SO3enYG+f9d2PmzpSXalhBsn1L6nF
UwEQGv6+mf7hs43bzW0tRv14KTyb1rNb+9IeQDFMxrp0A0+PO2wYMQthzaX+bjag
9xIWZCwcl/VThemWnbVpu2vmyAPxGxMFVllQDFup/+9zQ4R3D3St2aYFUipvfrLP
3x99eAWL3xiV681D3D3xguBbDwgCkbVCNE4Ls7T5jhHW57OxzX+n5WppOqD+RsN2
muD84EHBti4Zm+JuaMS7KyH/WSh74Cjj3x77eboX/7zOc3SJnDayKjp2CA+AN9Mx
D6SubqDOD9PDD/bTvjwmI5Qq+CvdxkAkzG5wOUyJ5eHu7F2XZ6LUPwAWdLOK1o/t
HPMhpxa+a2dSsYO0G7FjuVG98qL5CH45avo9yTjL6jRQKurJzMSdA+otFKlSS595
0u+HW064KtApJ7ya86w93qD6txXdW0NVqEl5zgqciKqvkmfCm5jJ0349DVTAF0lT
5wvLQ5fmJtBmiqyZwLpNgi2rlubty7k7MuIqYHXTgvhVVPDmJvbrEtA5w7zlb5ZU
fIOSAHQnbtiwqi44jj7448e8BIaYXeodstyvugBroliRNU7jhfVb8q1pLszDjKVu
xR40yXX54Zxz5/vKY9BHVic5oVOIKpXP7fCBe2YzWCpyPrQkSGAoUGswb5611v9X
OWEqMhhoxMfkBPdF3Pj4hO62OLIp7LRV18lU6hNbTLoto/F7b94qcjNy1q3kKa5D
FWLuM1AsTt24chE47bgCJlqVM8yZdKaZrUfAUb/nrSELuZwFgYZpImfRqnPR4Ap5
9jZv5DjhkG+AhYGSj2cLseAfgcTzEo1y+OpNsTbBerlVaRBfr1q7/vqZJA1ZuJi9
6pyXyirWlONRBqJDNtsOLFA7W6l3iW8lZ8jGSU4BjfZQkLVWbipJoFIlONMsVa6/
W7eCGxk/QKOcKt9x4gLMUOdlfxDfmlnUY2forxMfDgo3tLkGm5a7IjjPE68zj6WS
KanudBQ3Es1C7qh2SuFWFr0M4HOwKqC3ejyOAqyoqjRhK2JBpx3iiSAR+DipUYDx
7mD6roRQjFcDWFaPIrxv+EWM4LocX1zRiOx2qJVofiU98KYu4zzHzjp1G2SdxGwt
KIclHyWQ/rbhYmpSjbE4yysEJPtTAAeta8ubtkDOOcJ8wxbgc+2ICJz3DEstwAxO
8Roh1Rxj8UlgFqquK7L0HaH9OcVCL02b+56lOpk9N2ThBsSmPtChVu0U0z0i/Zmg
G870X9eZdD2KIU815pJhgvngXvRnVLpw2u7ipg+XmZ8C7Yq1lP3U83rI/Gh3+4/b
K7K/FKIPlwJ4HhhQ31KBa3CIHSkfkAu6nIZoLj8M+DZnRYDkha0VY/wAYzPI4lsU
WamZPcalIelqJQLRsGWGOj7foFmnpogrj2BAYSHET7GsB88BaHYq4mKcFQd3UrFT
g9ZLC2Rcn7Tssz1m/SXAHqp+PtOCwpouByJ8A5c5Nl2ZnPvmvOiWTxTwQI+D8N87
//snGXN2UGGzRioGkMF0rzZg3TfE2IUGXZDMjuYCChnu6fswLJ56TU758VLQrZ0q
GNoajJxGEfFJlVw1Nbcn0vHlxrqrM6OKyaLtHK13FWGh1qjIGEXf9toSdR4+K+93
bKHipw1lNbP8HmlMqBYCXAjX+kTxlzut9TylWnX5PkfdoMazL8U5sVHU8dIQnMrz
SKQHjT2a3XiaOicAsuAI3FbUi4mSEExZsybtmGaX/fVN7mZkw/yMxpY/2hb0B/hG
BTYPvj79oKurcdg05a7CwkpgM8H2abU10a9A/Ip7eYIFuwbkn1CiKrwURomyJpmB
k7QzxdOSZmvG3EP0/tJJ+x2sBTUPIpBXfaSsOb4EXRhJ64TT+cAVJ9r1Cg5MTaJi
XwM6xZz7DRQPSIYJt03CpfDZ52ngNXQb3mvnHDtbO2nIJ2uSZNxE7UdhpEnujdYg
TPGoV01PkJ9YB0L57rS/H6BxOkkvM8/1j5WNHMynxGVDrG6wpzJG3GDf9xt3h2qn
3+PBt65WOz/xZr6EUc27pOzXecc7hoCv0Ewp4b5ZGPpUZC10fAYC87EYklqgSyU7
yqtwSbKcyaAKy8bKwiyrXR7UVGmQWeal7oB6YQ9rp/EXsVAWmBYi2qZ78G/MNAsN
FTGVLH/FSedryQ1TcPLN9NTwInlLovGTUNzHp/O4E4dPglC6cIY+AACp8aOmIrNG
S4HK5HLD7JUMxatT6HatlTmAhUpVSd7tCGVww6s8sUJYr91IwFEoOsdNUR/Q7w1a
+zplprw5vkwllee6l0IMNeEG9L0YjwuabfTy67ZSOEZAnjULlXBeJp2q8rOSW+0P
bJ2TyAgnqNftDJLaTeyP+pPMgSxDBjaAcuHNP7LBZDXkhidGPEyg82KlwRAcbNOw
ObSsFKGh12PWKZ6r/1pBxCcotOYAmTpm16voxE0AWLvp5MPoff0+dDQqkxowBDCI
7t40+pJ17Q0g5KeVYOO/IevFirSgfyJEi6317ZzcjqYkxi6zshnYwrIY+tUa7PwW
ILi2D1mcVS8t6ym5kXknVYIV6qQOY9zu+csBAGhZ9qyEIAodFprwZKE0FAGTYGOF
sATMOOnPvaicZKB871thl0UKRvQzalKqSJEg0LzTIzVsyUUD+J1+Y8Vmm1ufGt7G
e+m7Tb1vbPAsEvJzYR2cmiRDJs1Eu3HpaVF9OT/zRlC7QYZ6HWu5INWZQ5U8s1OY
sHFFVwJxSXtkll0rRjhE+MT5cwTFyTuua0OzcgaUGc5yiYpsUNiuVDw7Q0h0BarV
ctTE12DgSZNkmt3X02Aw3KY7hpp28jUxaC17u7b4SqrAhZ5dFlTlkhSTjms6ChKn
qtFgZt+zmjVihzZ2G8KlmRes1jUzFe8jQoRbvMfbOSV+H+sC+t6rIBGQV6xqYkxG
cub4LaphNCZu306SDwzL8CXkLXKXMFHK8eJCz6RZrtr+zferRjk+N9K+h83xfAPY
HV8EHBNTRcBBvfoG/FMPDXXS7FNiw1gIQhGU78Wi50Ye2tICHE3rkKhNUSc+SBzj
wzqXK9UTyjXenQTBqzNHswvoJkd48FP81e7EXAGpJr4N+8TwUJlRvYPheopoTM00
ClcyxblcWuAUufmQhHPlS0pq/1fpzLTLOUp+OaLhOuduINh6OO/cFPmvC6eEWFGG
cjC5Z6D70KCGKQl7xW26Vp6kwuOwPqLGfZGT9pI1ngVrFc7I2AYNHQxWkrzrtGCn
Z3zaUiBshleLuJTSKLzIC8TQ2/KonBFDFR7ifq2/Nyd0lu59WGzX++YjuzuZa56S
DXoinBLsYmyq3nyH2yz6pu3xhnJ8FmKwkkZ8F0livnAA5ZsOnQHMAJd9C9O03dD/
T1v0HoZuit7Y/a1M56znYHARn2BhrQmDkOsUrR6+uUUXN9/WEqDJAs65WJEy6GhU
vRhYA2oC2SiJM4QNilbm4lCsqO11OWq6a0uwjJa2uJmYdYxS7hlfTU+zQGi4MMGo
fZr+inj0XVGRxBdkRUpV5ca8y5KvYT3Hr95chjUFdb50x5EFTzN3T/Qt2ZpfeKfa
AVDO8i/RjRaQtlXZFa6w8eOmsj3zjJfuAJ8Y0+EwvcmJ5bP0G9vCdgvUVRZz4+AN
aDG9W+v2FeNxUzH+Uu+uCrCKhfQEc5rZSLlSbZtxkEfzbOHQjGGvDWq5+pcsERjF
VkSbwMMI+3zLTFpbnSwgUQ5yqaZG29N6mL2Q99cQcDPEHM/xnonzCjC92ZPOpYEX
iujxm54yBwe99W4fDohoLji9gugFZ1vuIcjNM73pH0igUXLuZ9xwtK5TmHpfstyj
Xh6hF8iC0AcTQoVc15C57elhRcy1z7+LF30nPWTr7zTkSJQoA5kngiJ4TVR+G932
XOkklmOtUCnjv1KA0hm+VJbNX+1I40P+VhD8F5UTAfPEiY5Oe0cO6nOu9/TfQmti
03hzl0/cHtO82yDW1d2UrI56woKqknWK73+13OZcwKCQVqlGfkcIf3h5yxZiTkG/
HZlg02UjjOJCa1bKue4H5fkPwWEqTxPtQHlQ7yW4WWOwZz6LwlwkbBn1t7PjJJsa
3moZ5Ib+4rrRvhxb3upO9O7RVrvRbaKqU0lIH38xJHfq2C6eGjcT7EjrpehsV8F5
Wrhq9X63SMQOLVcYMUskGb2NI/9AfBt/JftJSeREcre2mWodjB/FGx05IH6zm0Ql
bMuS8sp6qEyTmgDyQ0NwwjYs6WBvUKeaEGAasQ+jG7LTgZszdpIRaycw+T7HXQGI
B7GCeqArZBpQe37E2QwdcoA/lu5R/GRj8nsEc4dG9tNEoPrGrjyWQMwGts9eXNf6
2sEC/ms+y3Czkk/pbIvU3O8MVf0r4kkconxehH6RAKmJ5yhBKciyTyNQzC2Q9NoV
E8O5hgX7iIWWwlCmX8GLS8hSaIW43Y7ZNx0s02qXXRjjo3z1ftVkI1mj81qgp8Bb
thAtdhaVfAYMmFudazSv92+ZC3H7TqW1+NI97JVli7IvW9l1xbx8DBR8ERDuWMFG
Y1rY+bFO3NliT05bUpq4QjIos3xyEq500U2p7tqGZmIN9Nc19c9gLbehmo36Xi1z
yezhf5hhuJ8+VGClFbWJ1JlEvx3cS/zk8mck6HfwN4gMhB7nlSYO0aEM+bhgaQUu
kxDPzyNewPPKvu7KTL19CM4culVVYFQxNBLfXhM+bxtdYB3fI5aV/yxJDfHCt9XT
dzpRm6u42hzOLyXlEJcNT2geCZv9Q42uKd5pOEFJom8RVFlPRVWrSJEE6IYDK+QF
nsMYP79A5ZHrQdOdXG1PrLV1ba6y3rm3EYw8BdxfbITsNr1R0zcOlsUdx79I8r+B
MlKl/bQfepgrv0JUJNged/r8euzc9wbY04o8J9/9y973cqrNrrr2Q1jGuRjaxFv1
UtIAtQz97zKfcDmIrGkh/zXk8hApogaP48mpacj+24JUr9R6zrLXmTC1eLJUCywI
tqzulYgCnyzpaXRFwj6CBoQ0lUSGiCwa0ptdD5glnES6m4c4HmmFWy3HpzcLe0Z9
ldStsy+3DuHj1vWFkNB6eSFs0I/NoA8uDnv644S0rYmaDdgshmHbK3QTxUX3D2m1
BWWg+jxvNbLr9mo1prq3+usvmnz7LvF/I0w1mL1Ez2CLLq8qKYF+/HvLdfGAUYeP
QQh57KDmciu5bc1zSJ2N2l5Yt6KYdjMbSXfP/Wjy1k9ffrldwLNBnMQ/Z8zAfTbM
hwtGduCRKURppbGO1JZ6La552qQCAVPPNNputSGH5RDfrLA71ib130n+iMz3FePE
uQHUX65bSr4tTKgt+u89zFzmcVwH55IwDQPzc9rEY7g3HReKWJEXrROFnH11MW8E
qo5yRRAbnMRcfQZBaJ6LcqFqRQ03XPnYHGw7p2+vaddbFZB334VEtuXvqDF2a6PJ
r0rLnBPenh435YkksvLrQXsZrxhZk/SlBaro2NQ49zgi7DpMeSWalIptnS2MA4bU
n0IIcZ1+kuKZ4iJacqJvA1DUHXFM3H2DCr0NX8niAaFIadew++WLy0sAjQFkVaw0
8SRFx8u/2V6h8BAdPK3T3kRIyhBiovEzxJYKSJ92CJrCFy5Gop6Pxhvfh4MnnSLy
9KeRZjYap/Xaj5Nu09qAzWNi7CMr9EszrWFiQbEN2qKljvbCVAz8Mnvt2SEeFEYH
/DNSVzF/8HwITzOHddJQMi2Zi3Q2Z8VZ3M9bmC7KjvZqBTsIRETo8Ff1ZxLRFmhx
zuKJfSBnyLePHqFe6MQZaZD43YNMuXxVxRKAFxD2rlLlBrrjI3JEvGDZCEMDmzm2
1Obo+pyVo4x1QMarI/drvSoBJHVDb6jC7B5HocHAd9MBuHX972jfVWpiZ7dJOfuA
+UTm/IDOCyT+6HW2dg7YJroupiTPw55RuuQFZICJUv7BXaybxEtUENGTu6P7DHxE
n4k4Z2xMqyIzB0eyDcm6SFjTlsIuByYeteFP0jQd64lbXNr0JnuR97kCmDH2Ib+h
HVT585kZyC6D42O2QbPeMAowK/QuC1oPv6difdG5bKfUqLXEuyKRTP/n2DdsDH6x
t1BtBS2Fhj6XGIFgwjYy0zvoXQcIylmM9mQOO+vyAy+LtqKq03yCWHRhtxTyVdWz
47G2FO90xo+50D9wpwTvmLXyhCE04f4ugBObkQ2Ge5VoMw1jNt0+YhnnRvktqBZv
aoQe96McJ3eW6lj5wpiOXaWRRBmkRMi4ZbsUeGV5PYO2Ad3IXaGiBnExIm+L2Fe0
bf4tO7PYX0Lyj4H32JXn8rj+j80ws59b+bCARFIrbZ3hUbh6mA3Sa0irJv3U4QLw
ZKP5HoIm4DQp/CZHu7CzoMfiU3yTRMF4kDb5k581+sWd3vJzS0Rg+rxhg31Vptim
v3PW8nkFYAppq9BtOKLKMpmdZnLK4nidFzj/dw9IvVAAVB72rIltzCqeeP5d+KHB
SMCcbWkUOU324ucefyySZpdgqT/hITaXWFJID4sEqbA44x8tp24GAwqLVzOEG6aN
jnrmDjr4sMyxn6l6b5bDq8tKSgK9JyRrFZBYGtxWAHrX9wfyY2AWk0gthaebIbye
cwX8VmOAopAC+0oDYrNahDKZTUFkRjBGZu8cnM+FnppIu7dbuoa2w5PX3seZracS
ARbIUpE+15jQoiMqJoQ6RObjIZW1CVzbW0Cqi3depyILyjTzP2tByK8wkaddaS0n
LRp437KzaKS/a5h8II/55YlwFQRFKOvwdO5yj7HCPHJiPD4O26anVeFi85T56xGM
BI/IGi4Y24nJmIEG6VQNrjXDfLaDsfKinBfh1QTeVF+F/ALPwFa5XLJCu2bnJuLo
lzSPX2bNr0uR40UQKd7EBHzHOiHbMvTJzYx/Abqp6nw0GsVw7V+8n8KQ6Ma/Gw5J
V4f6CDMKTGSwMQBF1g5BJm9q1syESIMrHttOSzgjDwodjeWW04TO7z7UbSzqYSVa
oWlBOrj8mukeqCdamFB9ma1i4bKzEtdkdQ7huxhF6SvXhTS37rbJ7Jy1HtgR5pgJ
LPu2KRjxiVCqXlsMgS7EPU2PRWE28tzbZ3wI9ad55KN8hKY6w+uzvrgQ11mW1OCZ
i91TL1b1WREzYKs6KEb5sUVtdOp4U6nNzQmKJBp9s/A1ZPG7L6GQv3lL7h9neoQ+
0+n8CWO3+DSyZtJxdv8GanRXiTltVWn5WLHYe83GATceTHjYSROunEXE9RHyW9pW
2VojURFm6e2r9hhPvIiLkhg0SagZbLiMO5zmqZbVeq6NR7003I5G9ZYeIZ/He2Pq
dtHW5a/fVqvBVLwB2xxYFlJCTQ8DLdwHyV6tav/tQM1PwfBX/WYfsHPQZZGERk/L
/tIbwc4XcTYoj/konjVQyluL1ur02ueiT8W5XmnI1svOv1P26IvL1cXQRWVks1Za
JL+tVpUAdBAacXSfEl2vZfWvG6EzwBSBDBFFj2LJe6c5tsbgsQBKBVoGUWGmDeTZ
6YtZrYtTLktvr1SyY0H4/i/cuHBJQk1nMuk9cBPhB6yEDuf/j9ZRaKljYDDEm1AE
VXcFGnB7GAulRcFG9j6Bt4MceCIj0yz9x3uKpcr/KSKdpSIdbHCTLP4vUfAIo/gc
wE5tP9fxuJqFEqSutK4EaDuTpMiVDoipkS0VfmVJrHSfD6MvNaveqIC9e28HQYb/
KxwshUlCwk5B0Ag4TsXw9R7nJ5M65+ZJYXxwSIXDXC3IiOH+g+rmIJK6tR7OysBF
my4jadQvqh7t//2MPyX6qjmOmgwaWDTLqUPig5NDV78hBTdkcc+aSysKFj6AlTCV
OQDLlP3wdvUmXY5fuC98BxKUqASQYxNNX8k82P6QgrBjQzxexjFKWBv1Kx9XbntA
9q1wvuDrvqbYx2TODmD9geVYPkXN2/z6sN1rcKlIwks+ZBitWEUbpoIr82h0PgeQ
PcN/SqTaWm6F5L3M1kkwzEhnL42fT3HSXwacc2Q5TzVl8/4u20XJAJhcM7hAK3MV
DUoriV9MfDhTq/2HLV2BkPSLCdX+Vg+GNlX/M7l3KnuEBFrn3nN2APFVEqeFXIll
UhOgEMqFa0Kk0/wBMWKEIvnmsGWZvPh7ywQGOUtw+gv7FI7nR62mOncowS+jVU+w
Sp+mSVTGgOqV5aLP08RUCO4VgMsJBJWnz8yH301kgzQsY5ggd7TlragwbmNjiVdk
pr70vPs3cGaWHNCpAU3GK3hbPZ5kl+FND3/0+/rgfpSXjh3xe6A3VmF8ChY1wWig
yFRaWNI3ZPbLcqL45oVvWy+igeDRdk1LkK0WF0y59ndYjlSM5r83niwiv4w2Pj7z
cMM7gs3050vAfu9nIKKkhxMcy+B7RhKggQMjvPo9WsJct1llPyw8Zu8HJb3Sx4LF
RkAH/9zUoKQdmQdkeXZ075+smAPKzCfaemrZgeroxR4Jb5RsbtteTOQAgUimXxMe
6aCWeTShiYvTJN6VeD9ZsKwPVP9nk19ZSBgFaXJc3sWgRuzIznFF1iIKHn2xn7wq
/mEyye1uuSv1uy+VWB5U69kCAw1rxSUB3Mk1Mt5wppus6inXBuzubYNnklT+5vur
/PT+LKrAyb8Cq/hGlj8Pso+aEWORS9GdEtbOMWbvnWmGeNgxiwOQMKqiHTiiJeno
S8MaA7M6pvpR17YttdbwXxqCG/ZwK1ptC03Io1Y5w0KP81E2ULAAyn566kHYjMB0
9wqd7Y9ewrH3dfLbh2Nm8jk3hNZfboQSWh6dSBrjOORQ4VyXzRXV6yaHU/pMv0qS
DfC6ML8ZKCnvS6lqRYZMwLxZ2RgWz8kqDIMpWSr4CkjdTNK7JaHOTuG+Zhq//u3j
OzX5oZjjyIgMV5sinwgRsSHAUmvrPVAaGOQHM2DZKz8AAA83CBAP5f3tjBojdiHy
QccNEQdD0Qfx85Ejzygm2vqhhDz+Hx3mJWObNhrF3Fimd0DVx1yC1asLQYoiGjMl
xLFsvo2PU+Td6U4mvlctTtuRYfsuLAhF0+EkATJYjTQUM5HAojm7XVw1JitNO49B
qM52JEoj3qo+o+gBJICddUPea10gO0laoc3lGdiFZv95J0AhhC5EzwxIl/20daN2
UMDNNw/n5z5q5XezSK+KY/08V1n1n4RCZH2MCSA/zwTjo/ZdT00c+/wwqUYA4rJQ
blFhZtfEL9tlGgzAlxIEz6bsP6XcldooIRWZwVAuoSS9m7JrcdfLw6F/VntIPgcj
LhQbU+MNnSbkBPQycpAI8D8Sg694JLNXBEVKGgmv9/6ByNJUvzkzigvomzjLiH+/
Q4w3vlrj519r93kcrrojjlY06mECW4x7coHAXvaQBY4ywIqEfzjhfms/aoe7RnNR
l49b63HxBcVePuUoP4NbqdgaDzpEWUAf3YM5wXNOPYKa+ATWY7FH+6I2PSS5W8S5
J3c3/hiuKVOGwwwKnPHNWvX6ApsEWKfGP+elHkxviKTxsYiK+uUcshKUCA5Uxw8H
MDTZ4adRNBB6UYPO9/uS9NYNIXwDkhP86K2dN44AtbxM3fK8w9BP27mUGevIKXWK
AtZzcR+HFgRwZfd9R/RcGnJvBXXkJeXxRooYOxI+QaJLe88b/LGDSbsE2oNuIKQm
bGRLtvjG02DL6DdMtkU5SnALzlMDaVNpcmgvIneZ8k7gnrz+OfYl9nbVN1rLT0UB
AVbY6Pwe2VbLCEOaKqKZmNIUHscdQOl7ZWhNbp07D2jmCG7igEKuNvcO74fwiHIU
+5U+DcVs5QpTXrdFVb+OsO/QqO5coFnyqXT0W44f8Tp1QloVDLKhOKaL8lkvjotm
4ReqBMZbkKTtStkR7ETX/aWyGU/Vwn2PvkpWQsyHtsG9NvpikPAaOECkfWF2Mf6d
R7MTPnckYjgVbwOOPmElm0CON93IESpg4PZJYg5cE0Ug1LvqIR8BmTntsZ9yS5V8
Fu9VWv/AGeZkX4eY1BZbmY2n20XSuCCytEuwbhmySw6sf3aXXfm+YUihDYj5GCeB
ixMno81xisTu0S62Mf0ggD7d13FmmRJQfe4QAnaEJe3l2ykBip5QiTLWJaVHAIen
7u3Da6ncwKYyTPK7lWKkCs+s/YfmP751GiBes3E/N2zgmipDmykqIhHA0jwqgdPE
qtdzk1B9jPSNk6UpuM90zaSV3BVcKnaYmNxal9r83rDdsbDuVDOPCDXFK/BXHKSI
2ekom9zo+Hdf+fxRp/FoWTzG4j44o6DHkpl3cvDJNChVgF8RoX0rvrngiznXqm+C
vKlGCb4autIN1vYtvTsFizMzFGUR3dyf4dGBa/AYx9f42D6KwgEYFVUX5TLaW1pw
eQel1YWouWK94wmF5ga2dr5ufJpvpumPz+dyeZikTLhJvH7NFTIzeFTQiFc2VbVW
HMaXpu1sZu8cyUsz0FiHEO+kVsKX8w+nyxaay4GngVMUYUDJ4jNVAfkHPk4SQTbh
UoGZA/RvGpcbR0ya5LyWjJlxi8jjK2aIPa8epDYgm7Pwouo3xc99AOUEHYcx7d5r
SLxStsE5wr8alkjI4mFHQ7JUZUpuCCCT65Nmz+nQ7lFLmfoPrY6EBlQ5lTafTno9
Kjd0+FYS891sKFUZxMkyZoGVA+xfxHJRuWs1gDpk8xbm7/r3vECERch5SUFbydhU
ndUbyQjDOzFn/IqPkwKmkAGSaBhBLynUr9ksjYbzMt4rBNQJ/HM+RmUzHleWmvTc
c7znSspehPa7fpFHXzmAuC8F0LP7BY4nQqJs2yqrw95FBdqZ8aEHLF1YEtAXlV/R
OJx0y9Ki127L6vNJ77F3fU2dLel9cAzjkimBN7lmXLnyD1ni5IYq/W7O/9t8v0/O
O7CpQh994sUfJiQ0qKzke47yAXtOsKkwdP7HiJZzO4ULiJp8zuXcM1CdkohROyin
IKmONL/tWefMna/LEPcW2mLt9ktO9VB8IvPMfatCtofFfSZ8H7l71c0t5vND8Vkd
i8qr5XZvbg4IkultEpUCCQLCFmHhP4l7zMVlVAoNPMDyJfFsIl+Pv1Yd3CchPNN4
8D1PA5ZVnsmXfWr5sheqsvsXpJIgIJHQlseosDJIgCiXQM06siVpXTawugpc2e1R
XEnQ1aYXxDOFoyxl631u6Yn/e4ahMxXVGtjhKA3BlrYrhecPHQ8E9luTHzk50i1F
dyy0xzqia7b4tLXOnL2MmK6GUDOvB6/ZuyUpTBmaOXsPO9KZ/Xa9FdbeCpjJz5ks
FkYkKfcNN4BSDJRxkAENuxAFpl+JdHHwVEBg7/aJoAdZu+waBXdI4+5tDqWc7NHP
f9h1GdGsDKgBzMcAlMEcmCbf8ZhjDn8f6HsDFKSsaqCqYCZqlFs7KeMosTASmLlZ
30txovAbXOss/fnHynkJ6EWLeHhMv7556pdJnvL7hnpecp62hUusBKO2O8jk1FyG
aGSk1Nac34uVRSb27YazWD5rxQMulOnAbhVxMZAXi9fl4UjlLZi3tKqO3K1ZC+Kn
JhMetHqEO2xnj4I1sSmXwylr0wqkCos8+jRjpyclU7pwdasIiw4h2EhGLmaMuSyk
MeMVNgqccYyHIevuGF0aTTJm8AC3ygXaGUUN9DRrIVzyc6WdYnpTQcr/NgxJ7qok
Rd8lzUKfsgzVI5K9lT3MjlJVnhPdgN742zfxVFfZEN7r8g9k1HzYUbE7ayEj2kXm
DQFSi4KXgc1JQky+epk24Dg9MLH9Antyhhf8WvQiJyTr1XzBoYG382kfd/AjK+vA
aNHo86DdqiPUfe293MO2K6iRXLT3EcVnEFV2gU/x19kDuULb5VYiCE2HIID4oyhU
gKy1BM9HsY4HfMH3Ypf3i2XwMmzQuM5DE2I/btt1l/6E2UzY3QxqZxRwfmDIIegv
d0agwOi3RchRX3fEsfQHl3hWXhe7IJRVwzHQoCHAJdyCLrEmYMTaGKm23OENeRV4
FWuaNzxGDfBZZK31yPrnbouoT/Q8bSm+HaKHUMAjN2iF3z7RuYSWooWtDnhK62sy
4/ClcsRZKPdp9fxsfxf1KHQ4St1i+A587JqOuZRy8KemjSU2AmwHT1Vlkr20kDjp
5ZAfKX1fFcvvbUmnrKP8gB3bJHZ14/omJQf9T5sGk1OIlZ7WajpTk+/KIv6hPKhr
Bw27q0v7p3u/wHmbeEOi136zKPIjZP4i70w0mSWJeHz7mQNGCTNaMNQTlUcgonC9
OlpWEsSTyViIQz80pdTJy4k9X4gAfcQJLl4AxkLj4jV6tWTAwDLVoykaRx75tGsI
nEPox+vHt+lshpc09fhO9nNb8lAHo9XXK/rlUKMFtkmjG6xGWzMX9bScgCch+cVP
ZRmN2XDdh8GatYQF2/v5YOJgpiJmOoIIoP7JaqNpBB1S/n8JcYH/K9GhIoGd/6WF
kfjXqhbDio7P44OuRUmE781oKn/0xc02BwVVzkFy8t4VGvkrfMKAUom+HH7g5ONO
EE0Dwr+BM6qwXc2xM5p/3rQL8GX+luFbyv1levnpcnsyEuPpWri4wpR6se+VAWVH
8+8a5Z2UVqIdL02p9s2hZtPoyuTpIKbfzsf412lZDuLeUR8GrWrCUGK/zYPG147M
aq+pWfO2PDyznbYj4cFcKDvdFCbfpnmoXYTJ/tfddfQqYheuSYMZ32l1BfkVIpX4
dx7IcgDOW2li908dwxtwxhqrfRXPn5SRuGN9YMTgzmlAC9t3q708M24Go2CfQ/a3
/sJuFki45V3koH1vYJK7zVDarc41FLirNxhe0fW7tNadqaPXp4Z9yFD/5pVP+/O7
QBfbWC7YQLvm5hGNjIa7ioaBXmRauOjh8zX5DnmMEKe2SUMf70m8bEd7PVfq/3qD
K6aagBpolUf5FaVT0X8wvpRLQdzk/cikLlvVG7pwg/PPxbYQq/pb7eKBCacl2XU2
tyHs29gtOjHnrLlXVPCpZ0yNAxcVpFGhHyLGYIYp+zAug4ON3t2qOZELVFjy93UW
t6IZe1hKIWANb8CDe+pnVzjGmpC/T7boUX9yLmHkFv/DcRJv78ohcDGuZ0lgx5nf
aIYxFrD48jKDRRce9WawbRiaFuP7JvmDgR5BfKuaytN9buYUIZJHvW3S8O9+1Dp7
8aKuNKhpKRK4nfzGIKP6mXuwtU26ti3IGfBMgK6L2KdNEl3xxoTzqo0RAH1rAF+A
zKkHyI6rZLQ9G4C1JXIQQP8HSXzcXm0FAAdUN88Of8oBKnTxjq1W9C2/XADXGwnG
P3qFmOHJWzmAgqOEqqz5iWMlF3fGWFkSsUCG8ICoip9X/yO5y4wqjoRPXp5kR+Ko
fO8m8izaWz+ArP0YNEw7bG6aZ7b+v6wD81re0OaXCKKl/UsopO2QGhQyNSugdFbi
6k6RUPO0PQV2/bK5Toxf8rpzRIWUAJOMdvkeSFj2qnmlUSIqRWGg6OWIIou2XrxJ
5EH1j6KsVkJaueYhJgkMfkOBwgN4jRlTjG6VPh+1KIFw3ESPVZpugZtmKyPThU+L
W0NP0bBIalJwHWPX1HplRBcvpVC+r1/7Ge6GF2jmlEgMEwk1djvqz+5NF2VaJfUp
dF6/K+u+0J0BKaOJ0FLEl41gWGzfZTDlIAK1NjI/Xb/v6ZDhUv5+P3qZzKO6U6nq
ZYfBdRcvGMNtmzSLpiYgSF/grlkeovSP45q7TmC3W8PM144xWafT8GQwvsJV1gJT
RtPzpjs86+NFGSCf+dG4oP832OOuoHE9xlrT1f1mT+A+L65KIKUMbEkZlNV7/92l
u/ghFOoUNQw8T10gZILzNUDXOtuYJRGO6//6hcMjkjd9iL9LgSrmzeDKqm92g6Tu
agFgML5jgChVD2oSWSVZ+wpl4r82+p8iPCtAtd8kCJPbuw2TCf7YE9hdGi3x+OEZ
LpjEgU2HSzrzF9FNimJND+JYhddUOwVxf7zGlimWFIDXTj6kQ6EOONEgeUznIWK3
HBZvx7hgGeNwtQLbS6JhCAonL5Z8krOvYddH4W2dAsGJwQTxqzhmRdfnedwZHldi
fONvbt8H9IcR6IKLVQN+XS013RZ11J9TPBUWoOLPMLUMTcqBBPGKkbnCOKx25K9/
VWWUxfHqycj00hbvC3tSJjK/nCH6yKZSUUdmPol3rGrZijnOb8xJIe+Vn7vdaGJM
lwhjv+mCjvO0OXDewVnlrv6ZdhwSAToUkw5UJ0va80rctRE79B5fUwXw5byqfpPZ
gF0S3fY4e4QGTR1ShjEKtuZmzXs8+2q6Kf0pyigMwjKVna0SrWKlLNFnLmJYNyh+
l5LCA0MaQjxe9SGj7NFsBMBdywx3yGaiqwUGmAHLLZPaLr36ohwcWKURNfiOAEp1
oXtKcWo73iHJ1jxxfgQ8/0D9YzD6bAqYk7dmbSmyGmgmPIKRf5U7wVLZHs8IySNQ
krR06N/5KzustgQXTuKep6MbTvDdQjFlhthuk9tXD/fWmg3fcD50SsLXu4SihY/a
xTTrPgxptklIWaNUS0gJo8TfGRxD/Cy4qo5Tyk5R20XqCBnw0Zn0k847wD9+Lx6n
IfejLXlTNovwoyBhyxd3PM8xrMvEu9nj5sFeb2V7yPZswXKUg+l+rQtTtoMhOisx
QTN+dvNwOHWkKjp8SI13LR8NI2oCa82eRTcT/LIDqlswDyhBjBzTfnYTJmB0/gEP
iuQQN+vyM9RMc36Sk7VlfAUeOsCqCYT6HZlQ9h8QcoipxaOMZTqND967zaIBj6Y5
s+YL2XW//3IxqAZEd/nePNezqasMZenBSwnDIDFB3NcFKz7jH9QKK5mGqWQHxafe
qLPjEaoJrpKtCAxuTqd3civTn7myn9d8kSJgOGKanT5aZvvI0gJAZOOXYMhWbqz6
/JxcWAhZoCp3MI6rbiI9axLDp/t6wItozDzpFbfrpX5ln59B66opGe0MOrC8I3rT
ip1+zYOzbR1pH4sIMwVshQZYzpCV0lED7OhffMgt8K2xmju5Sd8keUfXKxALDZ+/
lex+Dk3/SQ8bh2F4NJrTdHtoNvh2tsRQvr8XlFTR2tNLT6wSE0SXTlBrXsywLBdk
7xiFCJRCs/BsdUURcqhjUR+G/L1AzjMXJ9v+7as2ookk17q18/DkUD2xSJEKII0J
pTvhQ8t7kAcSs8RfNoshr12Eiy+Z7HuWJALIiuhTTDaxlOU5iD30CexzO2h3hgRt
jbL+sejXTLFPYJIVZIuw/VjEYs8DooGLFhDnogY04L/bqx/bP6n9cssXPKbghzPb
3ONridQ0HW+6YIhKe+JXM3QvJ6GK64sKuMJic4yywk5xlWqXkB406G4wcGSmaJCa
DOWv2+0RsaMuV8aUAVrp8C8EZbbGk0m6YedCCuMcz5hUnZAXqmOX1U3XPvuD6P2X
rgqyd1vZTcpBXu7ISqnpFjwVg61cpySAxQzCdwt24JKgxF4onH8F7XCJSn4hcDGq
l9dB9OqsGGaujo2iE5d+/9YfM1qVi5DTCgES4R+SDfE5j61UW9U1FdRQMZAio/4Q
V8VeZ1GXDZjmYL3o98Ku4HMB6aYg3TMrUMpkO8hHUx1uiRP4hIiTaS1fWi0bKRRw
BtzOlU4TJ5/jxIi4CoPWPrCEnLFJyAuSCuUPUo1ysy9ORiaLwO+gtsX8ihRTIJai
YSwYFd6geg1PWoPvaLZuYvMpWsfQOodLD03n2JPVOY6xYFf0voSkgjO50EwY9/3M
wtVsLiS2GSUzdslBI21Dfx9SbPyPrNkZSYWI5imN1Y89ZRlgxF/7nbc+9DxnAyQo
UTH5GouSb16CA2uwvWLJtIJD63xR06JcCw+Wrzg0dtEgdPseDSuKQaJcSTSx8wfF
tqZCr2z31mOwPyq+2MziCTWsQpss/W3mCuutzRvyV23PER7T1V1BzLylytdVH6rl
rjEc5iy1gAT4DQNEVAJ/NpVqv9A3C99SyJ0bWqQT8YqiMxp9QF/jn3fJWFfAO/sj
el0M5IsJjSHBweqk0JQzDwJ4d8bB6CrHHTfFf69zhJ1+tAVJHasSy8aIak9cMJz1
hPXc1Wsu03sEDpRMmZ7u2be3jAt6UBzx/RPFJDE1AUeKVjNUVQTxkcasccIuIPBR
72M/n+DBa/QYfQteRwh3dxUgSlAoaGsfus7Fi6fQPbuodr+G7LPx7+D1xw8xfjRW
la+oulNCFCtpFF/2HgXd7j2Xuv4j8NqFM8FSIL0l0FrA5i1PpJxZE/QjEvBDZsnF
Y+AkbJz9qwpQmNzG+BN2bOobM+IuEaryfw0XD4Bd/qOkwrcXga1AsMCXOcI3/WJ1
37jg9wmwj2zLqZi3y4cJDduNOsSViNBKc0I4e7CsnQgfsdXUnmshhBDxsHXc3XfL
ImQ38zza/lA99LwffnC0tV18JSp6vP7xDeupcMF3uWdP7Gc5iZUuzI75YBjKvFut
5q8xrDndghxNEi7r34EVMKNc44tR9SAkBT4FLZVVWTjK/KhylMPgMRvGSnY5kLr5
0vkd1pdcDB8r1o0giPr8ScK8jQosbnefXHWAQ4+B3N6cdhKXLR9cP5yC0Sa+xpc9
gKbR3qAhjNXf47KgghPOSD0RhggMCp1PHbJMPjo2YLAkSlxbTVclcoXnW+PfhucL
XVY7Q9AH77uA1w0TuuoOPoGetoavh8T/+rhDe+7IEiYiIk8GGTJ+zvzJz/VF/9Pr
EG3JtKcEU21QG3c4MTjHEAaUNS/11d38Jy+ez1gVCcCezEXtl7f1i/rpKOLVN7x4
SVaWPBoX3i+HzLI5gUXaALA/jqoUG6L8FJJBkQColIBwmZ8QSs78ErY6aXA0fcoF
vDosx2JsNP21AMJT2q+kPreGgLGMwUhB0i7S5818vF6nUcmngiZtlMWAfj4XYtE8
An8bRK8cSbBQp2IqPXqTmRKp33IQ/iYb1RhA/SKhoY776/bAWBV4aG7CODB8KxbV
dbKVyEwO4aYDWD7nJKpUCcGe604uvPCyk0Uitc/MajHkkztztAhJBDJN48mbrYIq
DdlSiUQjiFBQI3LIYDFFrV5p6WUvpgXjGTYrwDpNTANo9sioDtiUmHOjnfSCLDaA
+Z11TW1xpanRCSg5HU9y3q7wZQSuk/Msb3i2vq55vQUoT11uVoYdDtjQXRNm+LgA
MvQTlWWxvxEaSXtMyBSgmkgOXdhHWYGJWJOZ4sdSiRIjXkSwz9BbdvmSPMhU1hT/
bdF6RDN9Bt6tNjjzs79z84z0ZdX77uOvaw1UYh6cC+2F/e6cnzJu8NjaDEsak9NA
WMYliHbccIL8vAJXq3+amaim3DtPu0drU7dDTfODaxp3cumKbgritrjerHbqX5qP
tCZYOjj+BAQII4DBLH3N9g4+SS+1NDaIpQ01EeiKVAnNq7WKMFhuMRtG4z8vGE1H
OIv4cI5t8WuzJ/HUXDbh8sn1lFXhtyRLOz/E+z+7JBp5g0j5NDYVD+QOzFUgp9Ju
MP+A5YNvcQ2gXcIdrras5YbLx7TNix8bmdInmrkkNDDWu3+33cUTrVlDd8cAUusO
D57o8qrOGtxeBqXwyRZfY5Ezla3UZiSTaCHAysRtHA5ZpY82ms0AKmVcCWxPhlqK
2CD6ORbvlJsCmjJKkoKPy+SG8EUEGWZ2Okn6fQG2yWbahHZdwFvMKmDd/hWobDt9
t7pB40K8WmVsfyVy4cKI7o/7+A1927npHBCjgfO11HwSTxcKtj3V+YU9073VQA4Z
IFG1ZRcp3XaXrYjEeKVxyCKS3qfBO85XMmrZqkXlA0V8hBf09d5H2xxVYPtlcTTY
NlA9fjxRjMoYNvYnuxFGo3WsbCbzj/9H8X66tKW7AJTThlMGzuF6BlVN7M59U4wk
EwVmOResVOLlkugdSGApniMkTbMHRWgoAnwLVSR2I8McsS5TSw5VFibvRsLKXB46
eKzb3fL9fO/fH3GCs+R7QvJOBspLI1oZFMnE3yxl2Lo7u3kR1m4jqsnPrVaBb0kV
T5+v/ws5bhUSeK7vBpvlxJKK9tDgyXk2/340bTG5loqdNsrldLQM19dlMikm4Lvo
FAcRM4ANhXfD/HoEaDgYWtpN55VU/+SH9kHyqxvREJWr8LcZqnNl65Piz2kjMwW8
qU8ZJZNgccM2xpnUR1bvX2SQUHcJ2kFLPJNTC40X9WktQTdAZldlbnV3SQZ8/141
m2LDdmzgDKI5kh6e2g5pv+H7LtRIP153azavPy1IEip2ktk4ZMRSfa3WxkJYODmn
3pG5JyDyO3cK9Co/JOLPOKMsQqX1DTBKq+IBusjw98gcuakfNYDtLWwlcX5YSU+e
1XH9KYu8qK+31qzuiYGYKeD6P9Y4KBpBrHtyU6ARK6dTIRTuaMNJi2RneWpC+w5k
wl9gLPzNGN0tUdYR9bH5nb0nD1vhPTSLJS4DUSDL3/1jtXX897f4EVlu9102UNJm
ZNLu6VMbiUfIPPrxdLnn7TVChgriXYV8zL21gvlQoOous7Bi9F+gCfu0P1JUBzcA
EPDjfJhfr9J3GkUcWpKSe6aiT6JX6McSnxSYBisF7hcwtcr+QsDGKR1ObPhoznAq
xAH905DG3YN/hOU6pMADz/oJSyTpil8Oxm/OxO8B48Dxukt44AEUk7wTw2lM5DoJ
AngrkGFyC/E3gvNJQ/LLPoUNDaydMszE4peECLx8hKXPG6we+sLuq2dbYmn4EZ8K
WXrawsMXg+WJ6km5gPBG9siSJfvSB0Xk6GexdGh3FhiOkZO5LVme23HTgQ0cMQ45
6l8Vg/6kJsDoHA0kLbgaBSIRnUdaJNCe9KILYK3yNW7dxMpc4dAXfn7UtTb1+uqx
G7cp6PgFK1+AAIKOYIHz+irDGjYvTEL5PCGQALTJII3E7p/+goDST01sSbA8z9He
ppcsq5cOpy1hCuwhWQ8velU9qqon8MA+PnH2tfHloCR6+/hCZXPAXPbjFgUarOjV
hKLEPygtAESa8nHqmaD47BM3Qh9LRON6q9waEnoE3BX3+u3FFed1i47iWfRxINzk
0T7ZLeciE87w4n688M1ibyS9MipNiWYSdXZK1dsaOCSJAnR4/XSi+drpt+mQmDwV
IPsUsjvjElIGZ0Fw/Iuz5+ZiQPG6qXevcr8uYD6N0C9rNMrCG/WY7DKWAD2brlay
eGhtoS1ztPvn4HI2jIrfyDJAyRyn+EtDtD5WFCWcRGyoDbRRID6ju2wM0KewA1HB
6S10ZZ8Mn4o3dPRUUsu4xfybLKlOY50JRv3DaDJmDTx5o4NWGdYFrWlelp1W1SPz
YcIYtGs05EEhuWFQy7ysYbBvGoF/w8BblhMMaJzI+xzUcBlqpfZx/clBUiTtH/7c
b2El/ohL5Ynxs84i+WiZ8JA1K5dBD9Vq9hFHI+SoxFhmQVLKziSCA9dwENXIIk8t
uHHoCG8wUbK7euq5eSAfQm0f2Rj2kF7EKwtWn2hjMkkHc/ktUz13i+MZI7TEjYM/
t7iM/Kf7pme4SpAN1cq4osBBsf7ajLSFPLL33S/kMzVLVsiOayfCXQXaLZOYt+8U
+4GwhwNnlthPXL7feoFNT5BqHNLLRQ53J/2MicTKPbolTOpSkIFWcsWLq327lJyG
AHYQVb0AbPjBk0juSwWKaS4ndqX3WT8aOiB0nEy6PLz5R6YxN4PbZmbUCte+4yTf
Zk7EF85Nwl3GbFeiRCpJdUOt4HuYITz/7rUInIwWWOPgfmKjc2ASEyvhSWm0NBHJ
DPDHXud4m/bstO8T4RcxLQAg+dxYCjYh6oj7yiMJ0QjEaQxdRO3Usy7kaL3KSZL8
Vo9ts5YkpjENy6aQ4nXukt7FCeilml/7hMkLGFo845Xz6lp+9Shlmc9/62NWh91m
Xnvd3MQOQvCOIB3SR8iRjDUBYhsk/yNkdvVQH8lY2MipPdkchJX4klQRFiBQerol
4TPf25dCp7fcMUUnH3MiFD10xzJSJObzfPfQQFeqa/61FJ4VbxPcO32uigFHFU/J
VyPxZFOce/6TYcincuHiUZx6AF2c6REvZHIexbK7cRQEPngLx8WTq9Puv6eQPYSy
9vgZehqDV/db+p38bFZAUOIpdIm6rsgLO7ZoSqHULrg02IhCErxemUKrOV/rxFVZ
3P0E5o01q6vrBTFDdcaVMUkX+aoN4hig31b2VRNCUhy+ugGScWqv1ZPTDjPpz+34
+Tr4oQ77bRLiR0SfijEAp2tjk82Y6pg4/4wLO6FkF2EGNWOrmosTumBvut16CKac
vXmCtYstGf6jMtn02T2Sw2rFed8cbN+1A+V8kQ3r0A0egSi5kcDVnI1+DwklP4Li
nQ1/4nktNrF+t6BS1t0pKAr1hLTAQJeC2WMHj0gXcLrox4tAW62kJy3pZBGCgUN4
XtipexP3D2FymXbKwYOWQkVpHhGGenreJGU0Hjde+SUjbVz775pCWUPP6EtO5FeB
Npih4WS/mVFEyTtx0gTsbx9abm2B4VF1o81A3NW4FhkgIBBsL2njFa7FeLgdLqy1
ol4Ja3GcFUVmeboa2j/qK9kynHDZHSCrrzRuM2yZ5Mv8bzE9EcMJPqghbn6IdZfd
bZFk6ElLsSou9ZAQLULCGRl7g2QbbfxB+HlKbNWq6pzMqb61tFMGWjkLJvg2f8uU
UVZ1VjIWxwH2I/RWK1OAR9a6Cg2f6pQzGXICq2cFYnNFbkWTQEa1FNM436gqPtI9
fHtG9+25r0xdBYs/EaPuXc5G3oAxgh+PJbqe6kadXthChbUJh3DYNNAQCY1PdqyH
fPiEIqubWmc1d7mG4Z1KXFNrwF/aPeHyLJbeO4llt5R/kKSkx+aWtOpVzYlwLqJw
pvndVyREhsXesi+AqqMLHFkSGaFzWGbye8Due07TQyWUg7fMdZb3qqek1FbXaAKp
lkx+CHhDZ5somLuh3veIPH1f+oq2qI/MCLhTNuCmPoRd6xNuZd0iIQklwmO6IOrM
tM1d77FW6Go7vOwiAY0I/P7BCDsGe88nHGHp5MdoE4BPDc9uay1hefv+bnIdOnNJ
j7fJX9G+YLPAUu35+aRbkg5JGen8vPebTYwTtnp6HCW9SFo6wGy7qSTE+Jg0Q+Kc
RWDF6tp5DsUyHpRumpBHXBH5+MsbiJeaSrdcjC3npJZIvfjgsZdTDJhOy/n6Ah8t
LTkl4xdzXCdznbklPu0FJbRN3Yczs/9qncspCvI+kQrx+6nIgwzHXxvXe3X95pwH
86pOJ7Su6XmEAlgpqKtsbWFOzd2PoPvTlkuIMuk39eeni3eQ9A18RNuJisoAe/8+
xw9vgF4190WDiKuEOkljzuz5uy5QD0RY2ZFBhA6ZyFKrY7EH8um19Ju3PHv/4IR7
11F82qfUMBxhnsJ1Prgq+mGF8z/RlCP/rWs9P7U0bkm0Gv8qiUT47niFMqh6y7BE
p8vjZdX7/zUunrakZ1OzXbHlWvA0SPEYzwB/yiPIOL37KeKZhfJTTXgm12JPhOob
kAXjTdPFGZgmqrSRC4RoWBzQysRXFtVxWR7kTPlqGaLkqse7JcsF0tX75b5QkO1s
m17Nh9lPLmlUv1zKcWtLxRyQcjEGNnJjKgVUvdnTigC628qwWRnlqsMuM5TVtK89
6yYRzrVQcPpl3N+MwgL0jewQ1xEd67hX5JYDTLe7UdpFCFMxiepdKCzrFbg6vUs8
4esuL26M3MVvGN5buQdirw/928BJjCe7dEYyM1Yalwe3O1evr/Y0Jz8cm5j55LB+
sOMkt/EfcYeF8VNPwkwGUn+pTLLxPP8aR6TEkoTYHsZ3RFF6uYtVCSeZSjv8LHpq
aC4TkGRy8LUr187nORYY9D1ybHf/rOoNI9gD1R6DXm/Jx4ZHQlYfqxqhnUHG4KvG
Vq25d3xAcf4jvzTOHc8j7Ca5MK7WSWSq38NROMkwu9eklmvdTu2Aa1SiIqTUak2T
lB6W8n6ubqiKv5laxEOAM+D9Goa4JINT+svFgmKFWW4YUR9ca6SsulmL+O9PYO/R
YKs2XRUMj6a644/ZBTbX5+7ED5i6lCOKqmKT1Q+N5bSAtvRXflx9qyFOpxoEsHLQ
Vq39qvCGOCBNw223ISvLEjFYgCdJyn0nwp4nhxzMMfj6Lm1CC3Cz/k2ewMY0tYQs
5pxeMkZh/tIBmIad3nT08a0IUuyHUcmqe4bIfZBo5ysXWs7oAzHQRMoVBrma50p9
97WVEegImaXLreb/CNGpNaSkRNeaR30V/VRJeOGOgYkf0zO72MchGSa/BHfuSniZ
SkCPsbyRNsly4gAsG1vF2L+J2vPSU7FdArT7ArkSGEuKr9Zr/5UYxkjD3PtlXMIR
MwnK9JPtOyxZP5xLl3nrpbBH68n3b+HKCtarvtotrRuJbNWPqgEq8JzF8q5lGcBX
OKabGy1H7Q1f1DdvtmqvZg/x0lOGG3lpaqb7pemap6jGdHHat8t0Sr09oy+kFYSs
3yT+dc9MJMmvSCIcpsebv92NAijOFWHXsCo8r9ZVbIRu+5UYCHk2QszeeYEvqgmD
vFfhJHkWHhql00Sw3wEgP5DEmX8LRieMHni9GhCxqeBp0dZ1u+QYPO5GsBvcVcXt
luiqjqFkMwvx2Sqt+IhnMmDzj84IJEMWUKNAcQz233Blyoq+vj6joOWaUJreVrbM
rit75N6qIbrywKDDFbmZDSNLfHvp4T1jv12NMhwT+Juf9uRCb1ij9eQqNKELdmyH
9oF3W6Z68+mG4US/tTRxd97RhjYS3zUttdZ09trY7qpa3EUVS1VVrfvb2wRXg9iV
3s0UtMUlmWj4mOHrgKLcwURak2Lpo6nNlEvxURklEkACw5tS1BoAoQVU5go2LrpY
/on1gWnLxKdlGjioMTuD/PB49xt8vkBbp0jSk4irOtDJKAEzHZashE2wFTrohxQo
Qr9NYvNB899rqmioM9xgewsTujFpFO7AG7v/r25i1fYtX/3vTuLNnoQysiXzuapd
czhkggZDsaGzBzah33nyIBLUNyBAwEwi0h0AhW+r1KX/6hJx5ylIol4lhxf/CYpS
yRmuwi7cr9OljQ/nZURLzG8qQ5elG/flKcYH0AdTCYEdwvb4JphJCS87C0Ylft7k
+/r3Zg6VSkT/o5NkVv5Ctic5ECOUdQMkaVYn4+Wcg/wPx1mBaMH6JaQnJcTzbrP3
Kdet4ueVkvNB66gA7DksD0zx3qnVGaZI4X+jSkNNoAF9PDPOHF/+5GA7ZSNS8hlQ
g3pMSrIjQqKyUxs8vWSWgZYneerbgDKAx5FPPmFoqeWI+Rk/WiLj3GFbzi0zbhv8
/qr4fk86JJBCnIKp+7Q5UHVJMxeh4DODULCRMWrfGXAvHLtmoolx54+S4VZMMvNt
KIzs/9vyJ4bdsbn7v7tqxTFVx2AcDm0vLqWEI0G4QXQ/4w7djvIwg+aC+sm9Ml3v
VfDa/1gwggRHH9urHOFu3mD6QDuoEhGiLrPpS4VXLvvU8lH4b7P27PNBXP2eTE5/
JVrjJKL2yw6bkiSySdK+g9ysZ2iDb+GxKwDrRGxy+FNesZcZRA/kW9AzLmAMkvuX
rNnAIiXGJgbP+PUeEGFloBVAbijfKL8MLZPHDPhEsH5aVvg2VMi5BnWRNlGfj8TI
UFI/Qq9RvTHSMxIauA6Jsv77wxvh0P7emh9+1Ym2dVJTUQwdbmsXEeVZdfweM7E+
x5YVOk0TNY641Mo1hD0/jHq3Di6KSZCrPpiAUh94jkS3IexEdxwOYKuhF9YKHfjJ
zrKd3HqV+MUHqkmaY308F/Jx/yeWMZ24XBSIUUru9Fp90CdgIaHfKPQSf54ooDPO
D8lQM1SwWDtn/dp52Gg0+FSPwwCteyAYWDuhKrBuUsnQcHpaufu6pd20Ug/OhFL5
ymY+nj9PURW9jduTzUJ2C/3ikBDp48GKbRy1I1BJzX3GAPTsBLZLAGA3//nXvRcS
fmLx6IbyYYI2AhTW17yhiggsA2Q7wglc0zMzRgmTGvMP1geRI11qdgIEOiw99TTK
uKudKPUfcdnFY+opF6RR5tSYvWUMYgVE7mZwfhe0wVJTYilXxh69jUmkg8svpXDW
TMc6f/ASxb1fy1fWgDCXHWrey6EfnANG2Zcf9/+tEfnAnGl/URZ8uvWa1lgXzWr6
ZNHjOgoKtCVOz7kNW7zPYP8JdIQttvBembBHgdPEpBvQ8sG8sYtZjVldflQK7z3e
oj/x1GykcMcbsCSii3x9V3Gz9PEE2iGyZc1h3w5ymFyBGqMCZODvB0oVY9e/7jv/
SIXagIITJ2EHi5m2VdMKksUCRD4yEGvPSBW1kxunBa2MJVAr6XyJSC1O2x2hEUeG
DW+GkCQ5iW3sP9cqppxqdtOjSaREro/AhwMFRoMIlL8E2fI0YZIbAVS2qBTO1sR+
JN3Gbsfeq4xl2VXvS7CazxOWCeZeJTGywJAlmq1pXTTGWGIUuvjZXycOifZzqUVE
fIv4D3NbufPWPtJaLtE5614+fWRbrIHYpglmIWdtI6rP1dMU6KZx1cthLT0lpYV3
FMgVKtFYZ2r2wr/hprdPD3PEI1L9/RP0xvZ18ScPxftLndV9f48LdGqXVkwBYzjW
4KNJnGEXAF7R9moyKTmgBQ12cntLMN4J9pyrIKKQX61sgqF+Tb1l4tVPrpTjAGU3
5gn7bCHgg9/XoRusNx3QSXlILO56dS2n/YopDf+7Qvf9Rx5T7dJeT8iNYBf1eiLi
jG4ahDAmzVUNzdKgdDAAS2ohIIoQsHPh+oXHBk2EY05tcR+v9hGJGU6nEdASgQ4S
3SkFzynXmeqWIfvZlFHlRew1Xh6F6CyjMANxlZ7ctW/npfbl0KJteyNitL0wJaAs
nEPKKcr7T1HlS62d1bVU4b9LnOpPZn0IC9WnGS8x7s75rQoUTT1E9DFu0GCLhFGX
hvqVx7BE69dm72tVmu2M5pPsx4O0Ju4V9bCb+v9gpcvf6hemtRwMKlvF7fL7zBPN
HZ3yEPcJItNTkJ0n1hQyjHKDzY8SCubj8fAOJY8RbfWiHB9aM2Dvp7oAWdAcUyjb
nsDaPegACSuX0EPlexopXtoMjnzc34iePnJBvrWzt8OSoIW0fa5dcjRqDhkmYDGs
eQtIpTEhnwr2lBpQVrWssssBRXFDa/kYgRWSs7F20i8XD70BtR0pxYdyRbnDl7WV
k2fnrGP4cWBgKtUxVUSFU9omZQzQTMvzT23TOmqpKBxFFfsDY5SDYmr1cMutBHV2
bQoHOm3k33HM8fyNgnP7SmAgcjdD6RqjmaO/w4kiUxYDpSks1Ntj10szZILzw+Dg
/QhR79Nu1cldq7APU7y4nq4NlWw+5SxbZDG/5vgsFnu37vpfH0eT7Qd5MWlzOVk9
FoX03d5H2YFu563INW4h04nYaySLcXCDMrQGFFBXtYf6B1Z0/Euu4+5L0UriRKEt
ib7y8YAjd0+a+KH3gfgMfTMW8a/QtZVp1K0kUv7aQ2QVA2IN5eMaO5PNub/3A9xW
PUEUzLmQrZCiRb8SPEXSKfCl5HbCHsxM19gfwHQNTQ1/ClEKVsomTDa06bgOZJq3
81MDpPF0Jjd2jHRGkZiDFzDS+BDM6DLtLvXrYI32yVfbOESkZdMr8NkfFzf1Awf3
kxlyIQ/95Pd7Ngaw5MaUG43NscuB7U24zYPEMoXjpcb/5C5Fotm2JMe8WNA4eLAd
hLoZdeuPlEwLBF+gCscDp68wX0iELYuOH2KeeKtE36RyTOuA7FIxFX9d9LyLO6kB
ByMPXXPt1S2rmdxhJ5gEKqj97vxJWUE5f9IUUbmpiW0oGABKPUndmx8XmeBfdbgt
uP8hSFID35Ykake+FONh/UJcuOQ67RucpmxUEEPM84IRiTbksp51n3ZHP98tv71k
anKEBZNadh3b+9dyx4rffSxIGZaL8IcmS7pwvjd4PnYGo+S9PWN4emShK4aOeuPC
7Vh4/AGsJztl+YRNhVSFNH8AgcW5z8GmeVloUCEypbkn9UAfnFM2gsGKnMM2zswF
Lk/qCfp7JLCFjQdwAaRc/p+Z11kf1DMxWpLLc+FfsgiUG9qe4arohZj5py+vApVP
gIoqj3LKocuLcUNzoFKS2gpZZwKjVoiG0DkF1d6cX7BZIAA2uiIK68KoUmZDlpjG
uafPDnf4slWwhVRXa+bMPnnFkUwQN0L2tyx4EKJhTwKYfRFM/+4srBD9fpQmf8LG
45i33A0h8qhoeWbM8+QDujM+zEHXIKupi/zW7stBxbEj2qc4emAnA50RzHsFA60c
MKP3yytfDsh3eW1n+a10f+LEUDWxyeyFkdYHP1VZNAQRWq4wSy9FL0INf31mD9nF
6hODzuTy9ktcjxlZvRyXgyVcs5J2OvF/EmUzDkGtAiMfUk1VlS9NmqCmDvdDmq1s
VNsQQx3zQylWTZf7gjtIXTB1h+2IYO5LJrh0UF2l+92Z2ZW6xT/Ccuak32BqWF3D
53IGkPRaAOXS4IafCVZ5RD/GT1n+XGa9AAGAY+zHQG6VMWREmSVjYG0d6azEeH1w
D/MsCCmnNFiKSeQoIXsqXNxRThrQnNcKqY1lUVFKG7xo+eQk/d0mtYlO5fQWSAFS
yT6CgEZE6cALXu9HE9D3oyCuyEp/7cJz4AC8X450sb1ja4fQYsCgHSbB59Yh4f8D
rBausovDhkP30x9MyCLbZT8pIz5Br6+/AAavGyesIIouTA6Fs6LPKTQPhSIGDXBQ
5GG+h6I14R4u8ZQlnl/tKqv7hSYu7ENHP3echiuuH2JGG3O9+rc8puFPGsNUksG9
k49FzAmZUgqCN4H1IqoPXOtz2Rsgh3tT3DgefAEENCUHvU9L81CQeC2sy/xRf0Lx
EL93cQrGuqU+QvoBPInHhMy/qn0L/YRuQBFzy56ru3kNYbJZANYYWDG8veXtRhcc
g1lpWEqa/zBVhk+pHkPpBMPHOuBJfqfzs8TGC3wb/79kR6CatyvP4aMlJv+DA2RS
tWUDaaKxeDzxumadoziZij2kUvrcQw7KuCed7mrQ9rU0zZRwRPD0theZu89hgZyT
y9334OHC4LP7/kmSrRxTnL3BtBez+agoP9QuwldPb+XT54hDVqqGMK7hRbI0lcAP
qakZhx4MArg5qC8dvss+1vIO8TgEvGjYIDuJuv+lRHNzMwCsJA93u5Yt5jwUW162
Gfg7DGR/cey2d71YT0epWXg/gpDtNuLzQrWoflcprGIqT6lhh5fKX2ei55tP8ruC
PPpVR0RCaGQTyoJStFNFAllgVSAuK1ck3YJdWNh67F2O1+TTWdVjI2DdzgcF4ZyF
nka91zbVZJLb7IhcONwh22X0MfgCxOgJNt/HK+xnWz1ZC800HURtrzYhNXKm1X24
hkgFO8lLS8GWDVMLretasrkjqU0ABQ8gy7dX+okcHYcqs+4L4THNJ5YGStv5g+dV
xKqEilstiLEjm+5GV37iuPsLCwOjhz4B7cniig6v8iVrhPhwnQvGbhFIxBuWHEE1
4Pnwx5fqh0ni25daf+b/7Au1GxZvs8Lk8brqojUDzDiX4fjonAAd65btapg7HRqS
0TfQx4+WqVAzpAOlNHdsWQsDIQ1P6xump1A65I1zz+vYRGg2B4Q9QcBfWA+KZeqW
SPPkWIXDmaxkjBs1soBgjUv1ebDSXwPVR/Qvf39eQ/z32xSANQ/ETzxf5kTpHdvD
vV052cY4I8rUpHSsb9wmuA0EzMVTv0yLt4mEetwH8E7Xb9w6Zvh4Bgrq+Pme4++u
5LvMm6cK+bNO/ClH7jPSjoqHVXjJ+YYph+wI/NffIuBN5KI8JrtgcBl8/G5LBuTm
0zmgy+PJS4w4B89bxg9OsuW4wCnsbBn+buLWD2QbW9JzDPy+nbxhrDPuA/WEHSka
w2ZL0p547dWxNhkjogkGghSwhRubcGMSQ6GA+iITUMWUECkBtOUfG6gw8Ejtl1Ls
V7hHH+Cb5MpR8gTXPaXeXcLvctZS0j49kxh60aBkHHwZNVDrCl8u/VNOfaI5qM1T
gxR0Cb5wdBJBr8rqOkGd4a+7hPLrAm0OqzP2J/LlNRgytb0y4GsRQmSetk+ms3wx
2yBGHfEECqmyAookC9L2SjvjbYhIxnDtzxKAAzl7plu8J1Qthd1rjwi6hjjiOCDc
n8AY6ovcz1WKJVvQ7uaWx17K7xVz8UDjGafFLg+0+G73aozH92ZVF8XL9UZEQ1OG
y9OO80gWM4u9ZxGyO/dECpydPbcw8C14pO1WJJVogsSOLAF1iQwwj6qBrTzEfGRm
XXCmTjO8/PyOpNIfmE54RIdAjuC/yv/7XqkRSpcijV77zdFdQ3Bx1b0TN0rKSSL7
dfLSHIXGj+ad7QZdO5KA8cjMe9ubZ2R8jJPm/YB5Qn78ifvWM5bFvbQLMsvIBSVq
GUM8IBdDHkm8yQAQgFm8CGIuSpu/ihlb3iObuTNdCA5zQUS/Z2ULQoV+PAB9KRvB
TVmgZHiHINUDwsnlmdie48IzfpLK20/f8tG+4VHPiD8TtM9XWWqzLltq84/THGT1
971TWVgW+yttFnW+7z2Mp6xPR0n3ZAH68ITnP5ZK8Cyr+totTkwa1Tif8i8ZveOH
fNjB2s07tL3+nejYSM1f4HXmg1Xte5A2KjLuWGR3J81YRCc7M32qsa9eMWRsZuAX
N6yqGq35WN/VDbEyGHDL+Iy5Q5rMYk6Iy5xUmsAaR3u8plL3jUWagnGQQiY+oRAM
biZ2y8bJFPpCmXH/iN+Lejwd5n0syi/vny2zCeB5u5275xtbzFaXW4+iT1vl44i+
IE7TePrZTPfjBBHWOxaIfwdjpMza6VQVu5JlKxb8H5Qf9AB1frNghl87oYZv5zFT
vfRxhDTUlP3sMcrJkf41tT4uBkRH3Vmy9vR3HaTIZsVN5EeMhJuQmERV5MSItb5s
hvKlP+NgBd38pA+TvfeLiDGlzVlABq+/U12YssTN/KjLJq2DC3DFLBwik/yHhV4t
rPS8gt/rBGHLdgm7NRc5Fm7zRzo1LSC17FLUH5OpYbt2RyxYzjDc/R6S6Gu6aajA
q5ZurHZH2YVfAsQZFhgUhY5pg6xf5EqYP6g5Ochpv6+lPWGsCAsFoGAHhjg1xSgl
yqwybELhU6tdkEsXNWF53zC9M8OOUE8k3hK1zgjyHrMi9cSbzC9C68qb07C+uqkm
mRxwYfpw6kQDxQwvb2hCODhPE/FhQ4lgpI5Nj3TervLkrdOWMncSsdmm4iwiV6SR
DXRRY8DZWgT0flfQXIaBAb1FNl6LeQMklBdIQe03FpbjdfkeGYV265bAmiEUENx6
+M5/RuvuFr3lJRFRFE4tD74W0DCs5FpnoW6mCds8NlA/uhJFlaXswy2yF3oA8yDb
SyH6ZDnAq+uKFqLlzk0Fx1hlMt30M7Ov1ON67Lebu/k8cAx1zn/kKapsQD8CgC9d
Mhlz6H0xawOFewWz4cKChLwu7eOhLfGVLNbjlvPVWzx2drYzfG2xuqf8HT3Prd53
CbAWQ2qJVJRSGaQyFHdiprHbfxBBiUF8vWNp+6wBWsBkUK8tEDZleHUdHHCUPiTN
BY9sd9UHNCAp6/l6D5JxJYPJJYuEsQ9T92yjN+UEP6wwY73MoBewYZcxZjKTrlYe
PYJ33XS55vh3ObP/Urp7USVEFBxdlO0PZaKCjmkvcd1tjVUKFzjLFFyBHPBqvhMc
+skS/Av2aIyLfIHaxpYHAqCsakdi++y9gyfLT+EcHn/a4GhzcdgcdlfdLLA2hs8q
6vkyKE+m6Dc41slOhyLCsfxnLRUmlhRMeq0h5F5D4M3x8GCFBxZptqgrC103ON3W
tSGJJz6TSDsJhuZAJz6Uj6PYj5Hdgp3VXKfXDrxPIhlV3aqGn+bziW0hJ8bHDAN0
Jrx4qHq3CdXrNEKjyLAN8ZKZX+A5A/CDU2ncpqNjpvcV4N6BkfwbER7gs1Dgw/mL
bg/uO09lJGEMSjXDoXwrM2QbcZbISEjzevRjw1Nox0UAl3awSe0pJ+Xw1qK30aEB
ydYi6/6RJmQRQT7sNOCSqRH1ArQal/Ns5usjM1Qo90eJQhnvzMzhk5Q4AJji4JwY
dmV2K/lW2ZeNfDflYz804FPioejEJeBzk2IGSWtKy2DZUxvWvk4L+X7H9S5uRXwu
OfVFgDkvcC5Jv8qDkvU+3ipuZ2B7jhVy12++BQtIuBNkhRXjVe933pTlYYhBJaJ/
W7Taj+Pv40sbNZNpWESwj9cjx+9gCMpeDptzPHDcQoRTfXsMqEnGKH1NTMLlFViH
156JV09+vVrmUL+KMv6zW4SgNmeXjIV+QQOAMr0ll8togdydzF67Oj3gf2zNqXlU
WpriDDHuUvVUnM1eYealL7M+soOGdfLmB0VUYj6Fi7RvrAvYL2K6XrMye8tFw3t+
+JQ2TwMNAd+YZvp9gvpD2wqgAq1OEDZupAor99msazbFM34/pXE4zZOmA9gt0BdC
C7SeDyogsN+I1HL2EZ6uSWCy6M0UmtOzIEo33qHGTWy0+Zm/kTU38u87YM1+RD5M
4x807sIkM31pWPvnHZNMt4qE+fOMI5hoa1tFo6f4P95IO34fLcyjri74toFL4HJv
8BssdXn098BZqwxoHvetrERyEWbzgi0a+7ieoibvcSnJDwntgS0FP8PfS07uzu97
QJwe8/LAZxA8d4gEO//tyfi9AdETnizORREc3Pcqn/vBeEpzwk8rSQsFKc95yT1K
eI78BYJq2jlFle9pAQz/oFR/f6alCxu5SjVDiOJt2VWEb/ZZ5qAROzLTTZxLe703
5+atHv2OVsLCLNxZ63PQM4XA8fl/OYBHquzB7aZHdKZPSS+1DHmx5RTA+3+Y8/m2
K1GmJQO2mLPELqGdbhkA4KXzGDbatf94VLqZi93OU2WZh9yrQRbgesnMtZIVpXAL
Oiidpnm3L77UfrCC7tcFDu4z+mHTRNsqguaXlvDaBA7bYxxXKp2gg95iYz1US4IY
ZS+mGtQj4782QOdKM6ArzMtfP2XAjbvy+xHu0XqM7HSd++DMh7jOw9LTy9SvLoyo
lM2GwC/CyRW7z5XNBrDYJt2evvXOBMByujvqZbLYeiQuwn4PR2w5tS4dYpk+sleq
X7+MkpWQkGq30qOq6QEAVQe4FsCLSdRYqoe/cu1sy51eRl4VSvJRHHyX/M+jKWYv
exgrykSsDUp1ZyhMCoHw7xdpJ0LYiSYEXDQdXQZ5SRoiesC71sfPT9hlXoJK6O0h
P6YuVU71wAaq/uJFd/cVnW/z321I/UxDxIvlS8Ya6boVpkoL6pe5kQVlXBvGl8Up
xhpJrC0x+0g6vowlP8k9c4cJti9afh/4vGw3T88wpT+S91QjnYOnuUNiS4M2tH0Q
PHgHumXbvYR2K3WStsO+2Lvz28VpeFKv+fGxLg44/eMbOGrlEI+u8bQRZDseJOyh
KmqzrWsd2rPkJE7kMUQ9INtTxethMu1myBRe7nJUuJS0yKYFE+SGtvz2AARYVXG5
oY1QNbL+K4PNucFgTaLK8S/725uUUER2veFs5UYhOG6ihn0fYpHKTMQUJ/kMQzmx
/LGGZPgIQnAj2A62maYT1WyuVdjofFVBcR66FkAN5f3ftNdxB396fxnZgTdiiO19
puwytVGaECHDcPPl+H7SX0mj+YCQqfArmgNGKME40W0qTbfre/lQx0ocYu1UpEni
7Tuuf71K6ssNpb/E7PO1psEHVgTSrcwagzSLr1pcb/tRwAXf+VAGY8J5L/OOA8/x
7H+e21yw09TZAeLeWVU2IGHe+IzjbUsWOGj56FId7pwu3kipJxQ3y5UXmtsV7snD
HFUOxtij/0TdFhL11i4ERDm9vWF2pTELdEsXzDz+5C+bN+Hl88TfmrN6O/Mxp7A0
GUB6kr+LhvMY5cnnhL44edRDGXVKdyg1Vnn1YBdtaGZUMEn71wWKNiE0xGU8DYsY
VWXvl27Nh9NtFYfVg+bVtpkTKkjZ8XPZdekF6m00VpdDpL8o2pUqQ6PJ94ICXE4j
mlVeFTjp/Ilr8wB5YvTq00d8BfugFu30jKh2zVwOl9ylyRn3Bau+X+htu9FEoR5C
7iuSe23k8SvRNyeN+Xp+3fbH4/gyBzGezFcVzx88EDpM7HCiIelkHQqpJxw996CO
x31R4jfpXlUBcbJYEXuyBessrFf2VS1vc+S7Bsjwb/Z26rYdDyEHlXt7ApZ6PZJv
GGiPujiLttaT3XYtkMBuu/XQc+t0jnXbZG+/b4bNy0dXTJCEnjZWwgcA31kIK0NU
1Q/LmqJDjT2Rm3/i6yjhpc+MbXeylQyJhQeEavRTnIzKtc210+mnIJva1fvnsU3D
6Kp/ubprdEDiDTTleoRJHISgS52sLDUBXDzYHstJ6Jcn8FiZDANE46pKjSyYHU1H
/fXzDiJiAoLVJHfvrhNl31tb1FKr+XymmhD5+hdIEw5PQyX+Tj64qZ4qdRI4dvDu
usjciVQK0cWYy5eE30fneju2im/sarqOU8MKnGeXJT7qaXCnwUwueUCzdhgFz/La
P89Ti3BbTOdKqKynHMbJeGm6gAurpLv4LFu4ybmRO7/3tgmio+V3leFxOohC1eFP
6O1W+4n/ifcC/yaijfJTnYkMvOJITpxXHd/BBwjl5EIpe72MiqaA9SMj6P6mQh3t
gNuICUWC4UQuwdIZmpSSmuvR8SARKr5f+tvd12fReHW1jBYZxUTSy8vjxr5i2+Bv
pR0vLoXgRrs/bbzJymJJ8wfkWtwAyYiY86Fh2GbcOGiTE/BHy+vVCITIYeJLYHBr
eVeRS6thyIFtITr118kyaRVHcD7bXIKcpMGweQtNDFZrfTSARVe8uGlrDBLX6NF8
+IJjcTk+b00v9aai2EmeSo8jF0ZS0RVcOdT+NR9MA31cwWbVGwLHvHAlu/sWdCiq
2ExJrwkdKVGil0+neLavjvibrtox/bn0R8JrkLS9J98ToKmL8g7k4+zdFUXELELg
tipwHnvRLopZYOlA+ry4XeJ0FaY4zXXNUUw1UReWVQIQGvns+20liFk9eDqbRPDB
036skwV5GzM8Oa10Z0QVR0soaFhsQEjCriTBYorak6dw3+KxHJpXWT1udxouFRWz
4++Gjrd+yMUaJl3s9n8vf00JXqrCyyOPvlvdGmEmYMX0hiBrepUMs2gKSojewJTP
+3Z66YPU3U9USs40i3YB15toJDVAhZEDXfa1lCsdXMgdqCa67LQ35GL9DTh81oOQ
lJeT9ucWKol0pEHjgoLnjWeevicf2HtPseeDjLxFGjYatCbgqPm7YmkLNf5dcPG0
z168FmmY3RzQmFWsnLqRvwqAWsHIryUpD2ptUp4EoQU3/OWr+h7BVFwUv50Kl8cw
y7WJqu53QrvSUiuMa5IgVT6lpWoPLRko+bx9fPbZdcfHuwyXCROx1E4SuL9zZwoe
szol3PtA5ClGf4gpFIV0kp8tW7P4oKyTaD7pHweZrssIc2l8jpCM3vyaPml1S/x2
yCqw46LplsVKVgTZ4plUA6KE2j5+iorzgjPEEaBtpfHmBBYDO7kRb+eLJsYTK9FV
pxQDG0EEoSy86+U7xkEotspl7Mmo0hNfbzMb6QTw9U2WAYgzqauyw3u0Ngpie8PY
SwP2TDIdw5QN6x5x/+H/jRwSCAasbJ4OxyI9sD+H4c6WXWQ1lxjfVY7MYUgYnlfZ
tFHgvJWXZHG0Rv2XjUZtrVIIe9ckD7Lmr0nMpsguAmLb8VmSxYMsT2D6NDT1BFRE
raopNeaInNk1srXUvn6zB4fFqJn0HUq9drpT2HqstSegJBqwxJQh0d9098O208ak
rSQ6TWY9Vcm0R7zMghkwsQv52YYBv8cFqRDmcPoW8myAxjsUktorHaEY+Ojte7cJ
qCPvLuz6McOCVk+9840mwz0E11Bbs3DmBDqfJ6E8munaI3W1ibyAiRgxhgMb5PGf
L838XFbwYT9tZxE7N+pZTYEVDegXenYGJen+2FB9Mi7SPDUcyemJXaALVZFdFAgp
fFKiuN83JYFE7DiNhk205+5TLtBSdGDUS3asrYN39xLjSvOaG6d4vMisNgGnhv/F
V3X23jBSchMJtgHMczVajhjidn8RYJVwI4QPnvHMpIc7Y4QR2tzDfnuCmqpJb/SO
HhVp79q1pKHesNfdAMF46V8zL5Qg4G8wOfoz4uOTbRWkYSC9cWyONNF1UUrU7kpm
eJj2DrUZx7aaQyw5CYZNuPyQi2YNl/vjMVPpMmGUdgggUeU3EYNpIG9O4+WIJCQy
GGjisX9cQO2CIB5DycB4kyrS+fRB3Nnx3cHlZi7NTmMNQlXRTrx7cl6znH8PN32y
Y1eN+QFMQFf8k4ClGEaUBVgyHoroXPpd3hieh83pIG7uL6CPbq0/PH7tjBa8GZ9F
tpTVWoqx/S3k6V7MfkOYVe+meatqqHqM0zyeiuuNLQUuREmtO+y1Q8mmwlfdBKG9
FColz3D+3LuljglmvbkJOCdknuJURv4cUUB7e3NxwDX3ONYIVPnwZVSRz1LPNKSr
uhI4HnMLQA6EPkJ5J+3CEfpjT/pppIPu+JbdeOD+l0VcI1RtwgagUUH5vPeZZFv1
bxWyOU3uWxjhQg1R5ZQPdQGSNTS34CfHW/YTo1UO5ZbFcKvQey074HQv/VU+EeBZ
VvEjSKPxLHdzMQC8ks68K9nWpIPzUag0PK2Nm2YTpUJy19h46eBw6JMPH5PnzOAD
Pi1tfytHZABYH1lR66ph6pHE6h5fq5zqzgK6bJm5yl63nKc0G/W8I8L8OnnUqKGv
pHZ6OcM8eOj26+chWZrGdMxo6Qu/1UACWiFJP3XnzOrZOPXoqENm7FzWUlTetV+y
g9JNpY25hSLFoI+owX6BSr7GzQWW/+d648aY2zrth0V71xa/JpQKsC5gZVusTXcQ
ppuDtw0ZRUrjswka218itKVCfftdzfKSa/OKN4AQk3ZmsyGNk4E5qFBjb+kTmMoY
BUuZPwAVojQe4ZMYMYgbblzOzaqE3wxmc3I6UwRPHPQHZO9wQm5Q6i8fliIZP6MN
ujc2dNZG5ZZ93OSwuLzbVWfOZ11v+qVw4nzQkP5Zo6cAUv5accYncWO8tp7oC6uI
enVfyY3/pZXb3e5hoqgLPGfKgnay3kMM4vKyqHHCewNs14bqibWr8YUJEVckhLU2
68WiwnDohYGENr1ABSR6v2dLOxT4Pu/RAiprcVVQaVn7yciBiCf5HGaNyM2vK15Y
RpWu5tWBVjWgilq2rOkWdBY6sB9L5R36TPBuswTXJ6fr9oY92iXqdOldpDb/9w4h
SN3QAYSRz0LAdrHB7ysWPsF2McFndpzVnALJFDVL7N3CCArSDXmMqtcuRxs/3Ezl
2PdmA7TYl9jpSJDuiQkF6JdxW9iNjfGCbTK/QTgK3kBEJc2iKZsFy8lUvNs3mG5e
l24uu5QlJx23qvnpL6PbkkvfSI/qLgMZsnzHfhSl6v46QIGb8mjCGsQS/uedTdbR
tsWX2eMYxiDA2Ugykblc4IrKvh7yw9p/hrwYdAf1GNkkEzYEO+XGgth1Yq+G7VPd
VPBI95oHIR7p/UDK7GO5GqgUc3RTHuOQqHc0eRZYsHYfdTOBqf986x7U21jmneqX
lyKQAv19KA11Ns7ANTxR/oD8sk3cUuMf1xSK72qpujwyT7t92cBlzn2jqa7vcqEE
UIkj1IWxiFfb/q8Id0ZLXgtsS91gUTpP5R4VdKYHNVHgMc9I8PSeWO7oDsRgY0+M
uK8KHnuoMhIQXSHB2ldX6RyKGU98bF3yAyTq6JCQcCYQLlnOUUU6Rhmh5xPs+Xl7
E2OJMOtT3VE96r1mQXALPspeS7uSGMaFsYoStbVVV6AjsgUy1e7BJcEDoLi6Ueid
/FxF1f5U2qhjaqyrDi0gXxaedk8W67CytaoegtMit3nXa1WEvu6lQj2S3EKs9iuV
SBdNo0ctuUPsmAnURShoWVH6OQA18amygD/ocmKCAxuSMOV+DdffvhPK5NDdk0p0
Gx8xPRZSQdr5hC5slMebY7pJqIlXR/vAmRfwrsJUM317yNeIIMOVNEapJrlEC21y
9TqNna4V1RTaQcQ2qXJmrnToyRq6lBh0kj9cPM+/R4xTloBD+Xa5OhWwQFa6/6Ey
xO16a6jF2qjwNiOAGZs/kd3AnWR29Rv2yY/3HisjvlfL0cqXuwWcQyZy47UWfHdO
r0//5WAChyaq6aUM4hjC2I/SrULSbNflPD+sOq20W1YDZtU0umTwqMC+LkWWlpVi
zEC4tI+5zKwawjhMWJz41r2oL4Sq+ysXZeHxAcZix2tWU7oGdCUSKW6TwHrRZEAb
qFHcriTUORNOPz+/YpLCJqiTRN+8n4XHxn+rmKOQQ89u/PadBjST06IHfALKayZv
lsFmk/RbTjortzm7dxjaX5tWj39zYnRZgnCb6hbJ6ZDzTMdp0NKD5RdUWVQz3ato
79pioxYA1COHxOuffQ79aYak3uzGzzsDY1ZUNTxLAWlF7B5bbTYZYhMypph0Wini
qMgyztrPwZZNgAWWMc4t8ull913BvgTIq2frMxLfcWCiwabvcwpwMv35tNqSHm7C
1M4Db5I5uY52EdH7VovykU3DMan90q9+WdAlGKn54VS2F0dnKLjXAVBefmqkFe9I
SMAY+ALMRtdxkOL0ie2JGloC47y1RdUoSqm9bpCQkx8/1l063pXtGEYOLfScHGVS
0qh+5/EGDRbzt1Zcw/JhZ2Ju+yK2iBwAFALze5Lu1FQ0uvvPGz5FCJCOyiUQw7BD
ixUgc9XyrD2T2RUAwMr7uauJeaFBUx3KFPDuDyXXrmo76zjA51aFc6cjMSFFrt36
8PVfqP+2rY3d/n7h5y61dNyKEmE+UMWsmhxjKYH1efc4Mb8oGxIzSy9uu/4kT6Jp
oQKn0UXWVIhTn4+Min3F19jYPazrXJ2th7EiTuQlf54yFLMaDbwfUikdYGsXW5BS
sJFf88wMXfo8NEcMcuA4wtjqGbNhv6t6o9ULG6B3C/t684jXAV+cCDgBW47f2GYY
4/md5JxwjId7eXDsZq6AOMxYpfeDD1PnncZdLI3jNEGJcfyC6+lALPEfCLCf/lC7
GKt65cTXD8NdGPlCGdpaBzxE9jypC+C/t+QyH+PE+khwLOk81YyRub6q84ZMzld1
LbJ0DOJLasUkZsxnCsu2CK1cybXgbGVi79t3Qkmcdrv3pLxCBbndCwMXiM4sv2sI
e4vavPjOUi6BxfheuddHuBJa59MzEHfvHUmTm9G6oTKTrytU0czgYnTJeXPdPj9d
+e01DGcGd4M1l1X3AazFz7rbepyF8ECV1CksmgP06tr9w/OJiVAGYF9jtyHGtbrN
TzJoKMYTlQ9EpXyZHHDAdHd9ke+QBHpLB9dLhSCJFHgYjEvvjOm/xwNt5glebC1T
+iq6upeqDtuY8c4MFyi4sw5Xs7ceb88jptR5ki4U35qwh2vHLl4Hn21dEcvQ05jN
NzQlAWMhL2I6UOF9gw8jOkXVxMq/eOgl9B5keLviJn2ogRQHwnAwnBEHO7laW+Yb
N0sbRS/5iNEkkvulBjsPvckHHLQFekKK1bKZ500ENjUklsgw/ZWjJ0ko6JmIkYR1
QPpeMNJrDwadgrBYxkZx+HZzth++4mcwoL+775BnR5Pw/CAdct5vuE3zC1r4imE6
pmVXOTWV5b4rvSGLvec2i9dswXe1b9c1DMzdi67Cs3LpmxIhG0yP/obTAuidfLHu
Tr3MVG5SVh6T16PWqnqGyHysJzaKtsT8c7mkcVhegsKGqya8loOtTjcdE/TzprBc
35CLup3oBG5O06xYf6+gWCWPFv0cs0Ta9PZAMZrsagJC3CVNIvbx0uqH8nyl1Bfl
pSlYt90ngJ93/KFs/inHhrEQwEXkmq1zG1w9RGx3DzdMq87HbGooEcmLp5rYL4Eb
vOYl9J2cZNRGKZ73V89eIzDvZLQPa0Fqi+SbWKYVJW9rORSLatTyQcBZkwc3xoc0
ox+9xznbDs+/MxjLum7JYZCMWPAfFw7s7DQhIyb8ifojHnfDcMcwA0YI4r5onMmA
lUlZm40cAeJ2iNZPTFHOflg38ggFe3uwDonR08FjY7XdBsjK189UEcxWbECRKTFC
Pv+2Wco91AA3u7CrOExpKXTSpQkgdDOsAkxSokjcWYnmQbZa/zPVvywgNbv5ys2t
x2ft9NP2+UPM7AaEW82cXDrqrW8Q123X11L/XyGCnNOFG57SNgqWqnGmeDAVl1/y
agwiB0NC6D7QCPV4YQxgDqdhuozNnVc4YsVEe4Y0dG1iS0JcxpMhaXF60R2IFMp1
WXvKroob1JWRzWaIMZIp426smhVk6IHFb9Vn0gZJV9xiKmCjIpph+MxYJjPm9VEU
8Q7+pOamWtJU9ys1cae1kxZ52HG8oV0QB0aDuO2hEWr43KiVa84wj8y9ZHCPH/zH
Mu6mTXxE7vUSrmRp2TBMmyVpTPo+B9DdRikKndhH4R4J8gJBcwP7SPYvqoyJg3Ld
Tvnr4DpzVvOrUhTaUqwQpbmRFc61eHBrwB7XrlDHX2pgUiPrHX72XDhTVCGybdOq
C10q0pZYmQmyQiF3b2BzgrXR5te/30CFdjNNgs3PJYEGgK4QJnGTSb/8ofr4UCLx
AHtGCfb3Jw0G3kMaTdg+vk0qudxhnp0XN53I25oTkZyFT8AuBC1hOaLQ2jeV+5+c
hGn+fVre0wLW2rKRyhiyh1V1DVX6rhR7EihQlIkicaJhLEqh/WBwB8TAt9XMJXGF
Dfx1vI/cF5xzg4vbHRRzVLv0y4qnl7TkoUSYl/esYCs3rABP9D7hxFJoVbXPtKXa
k0ee9TxqjDH4uS9TVzaeMc+NvGRHAM9oTaIMcY2U6d7yOhf6T86dg1JnQvdk3bxY
kjVYm3RGOhRwnV4m1rw0g0zXvcr9VwefZ+SB9xBfiUuMKDe9hnhQ5LaOhFIHdNnM
AJuZw/vAGzOJpjgYrpQ4bzAkfGR476Uw8932hH+UTLmFZDoH6Loe0I6B1WEcBAug
TWHRbXuk9AQZHRnCTtgwfjJBeUzG9gX3bFpp+b4eSwElqFfcnez/TJtkyS/RhBoK
OLr71/rMe8+HFGSlYbBnHo+iQpdVWAZSxtsp49KtH6psY7q1UFZmgvHpwxuoW1Y6
7a+8F5oY2ojIIlip+kG1U3uXeecjC0h9jLJcHnsbMq2cEX85ySSobjAxIwTQx2Xn
i6NdRW0b2PrGm8DX7Nr+KdaIbWn/Tv7D/16IvFM3OrOvCJehnYYeyCyNQK+prItW
McLIjvDoG26KIqgPKEgMzsaAl3mtY5gtL0OpEgnXLch/4Ur/9Cs1vUOCr8TPgIpQ
iDw9xlhaG3P4b+SqTwlkdvd4kZXDz2vUoL8Q9nRuFqXUXpE3qqv8V1dZC7JJ1N7D
ldXdmiNVI9n9aGd/Ll7US1FVlQM3xYL2FItokrz8sqfE2+AuUz8KFbf2pRudUCim
zxo3Fl8Gz4TDbrdo9AzWjAkZZTXQermy9lFjamK3zb7eEYrVB/zdypKN9LrNl8ZS
eQgYxvEj5kWG9//ehXKn8zXjloKRIGNRksfcO+6WsOkDp/Vhv1EK8TZ41w1ut52o
Bp3MJwD552B+pbtPJpCkIC1/uUi8ZHEvzUzToBcCKbWlhWuV0EOyl1cF9+RQoQcW
+/KXnwjwJFbjePqW9YUS6vSIn4LXeXpu/MNgiakHNqrbQl6D4R8CWpSkdORPwyHQ
c4viMy0yfgSXNEEVihRwOln7dbY+Jg+URNrWlbAaDxVvVsGYORJ5//Juti6D2q5Z
FPoRj15hJH83yIaKJ4yO3WEekv8xlWsjb2XFifMcc0B/mrc1LOeHAR2S/OC5A43K
qQEhH1gOBrb1ivU+w9dYnvbl4gudKDekaEhoRLmiBVq8cZ9LYwsPYZovFswghn9B
gvB9H5yMu/VdAdeDpBHHe/NeNQqp0eGhDVTq3DKt4Rfd9e+hGx43EsTH8huxtxA/
OSXNcSN0lGP5FvkpRnOPVTZP+Bb4zbIhMo9iMvjsclSw/DBY9g80jxRPyRJJWJMz
7bBCoQUDn1Amu1Z5s5v5HJzwoqrKzHR7kV+86EYosn0BPmeBbz10yd93AT6Mgzl5
OZaNdkCBKpqY1+2qWZMnM9wr401NaIJ4v+G0+I/WxqtrBkT8RbPjg6BkfDjSEasR
KyHGeGkW2a+P1rd4zR0S1s6HShdKzsekxY9La1D53G1+tfGvhbbJ4KitwtQVEONt
j0xQZa5ofUEtlI+ZjIQyKMow+pyROvEctWkxBRrMOZXIamU2Kvx6jGLUzMcmyw/U
JRT57C9L0+ZgdYcFc27RcX4uzSLuk99gGs0n2/jeHLzRuizs7fbCHFIBDdcdWc/S
3ynd0TPJVJUUInu/TuHzYl7BdAPmFXEz96aaw2rZuSP1FStSw1IKaOhT7hVetagJ
PBYgvbE/8oniRIma+d9SszTXFbyCUpVhi+CSDzPxp95AiBF4hZo3VcQZsvj8jkmO
tuBJ6+crUWO/Wd1m29oPbj5ssDa9KhcfhUA0buzMB/Jt4d14wkAZ2oThDafISDFR
H0qhejtElbCH+EzDCMmsandfEIxARDdRsG/PX8nxFt/doSveo+zQuhhF5oJxESKm
3S5YFVFKAv6WEEasp05Ezsb+q8UfBQOuzAihppqtusC+I7Vt1R6qvw1t1sXcs6iW
EtmFCRYNgIhwcp2xX56FYn7eKy3bVw1JKjtkq3WC2PZikUTnYmGHfXfo5Jpp1y0j
GzDVERe7kCuqtwbL3n6+dbOWGtFb8YGfkgpweoH7vGP/1G4u8vpIDvNEHCJikmZ+
iC1GcgrhhWY+gELWgYJeSTHGirs9BHdxPrzgL8nPAhSCVtRN7b0vUFyHbzWy+fCR
IyIqMLdDO3BrDRuVBgf57tdnGnJIHAiana5jEDkDl56dUz50h8eANJnL5N0D+9YD
Ucww4iPigUAxLonMcsfuD/55BrunA7q72lSVewKfWeiPaBSB9Dm+jezSj3F/jtYu
SB5I5bwoRXOVtmKQ7BU78GsNpuoIb0k5LCljBzStxRFeTZcqJnk8IECF9sZ7h2z0
dgBhQlLNLin7jGDQKaenwHIYsmNTw0z9DfmUKqmYKxeAEyiQGDPIakb9agM956HY
QgvUhZusgHWZ8t5KMijYI2uG5vwopy2RFBcJpQDlEvR69ZYSR/g/xUVf/Qls3G1t
RnKgYN9/TwQEyWlgPiTtT9GCO0iQ0SAa57RcWIg+2J+bSHgWVHY6I1DMrlyFI/QD
TKtGE15x+cSWlBKRpv+MJSCKLc+wGtxh/m80AwB2frOrgGa9dyTx60xRFbh1tSWg
XTp6cl/8U6XnEplBBd266Le3Il9KLHxmR2/tnUhpQ8Bc62qW7p8SvfNx+HzJiAuY
BEZGV9AcXuL3faeSV9YGbp6jZ+yaFp/za/C/iQ6W8efSWpgbHjlhvynu0SqjXdrv
DcpCpsIh4U2kMHrrzetXff0BO2ownhLeoFPQufCT/ifQaLpwpKJQ8gWjBtz/jokv
t2cQNbXLKj8M16eeCIldaxkUZfWRgLy2GemG09S1ZqD8B6v9Tkw5uBCKB25hjDQR
T2vQOO3Hp6H7KZWC62eGXtGbODrft8wJTKlMP9Fz6WOUgACgB6noevyWdH+MkG09
0r9Y0TDEjGuQkRtWHxMDc7WaJZjcWxCrOKCGUk4N0Uc/5/CajzVrrZj383tCyRqO
jY7cjAIcBNoPZlAhbfxi7PB4T+FMA/qPY6QQ1ul8JL969S97qmjZiS0UvaWNfILL
dNxAZRf+0FNO4sZ51rzMGLDQBoA+a5AMJg/s9drz7siHWtv9AAtq/wnNHA7bDWRk
y1kbBkZQllgw7Yh5g+90R48IxY0E+UeguF46TcAZKEMpv9UQB+NsS/u3g0vgbOmu
BngYh4ZScIlVUGH8ziCfNgP4TA0udFHbOvpbcrHzaQAHve1Gn5bfRtxQsrC+R1lv
cL5aI4A7R++vvNmH0SClt3/1I0lboZ7v2IvsVmxBpv9NEdEnLY+ElKhbZ7M/uOAW
N4yfqc+aiJyt8+NJfnvSZEyRWfXamkkJqaVoTc92A6SdOZkVrgZE6Ig/Nl0HKlEZ
bCwdhUwYE4GSIVie2ofrZjY6b9zul41kuOyIw8mfVecGQxX17pf/P0016TTNApiw
32FKpqAtg012gI63pJi4VCNzQtFrtwr/i4/GmMwGrBseaDvMQH403rhzImv+/B0U
oJNyAPvQ4FxOxbIdyHJ/uXJEYm7hIh1CM6Ig3fRpL2Cq0jX11bL35cMgmnfZi+My
Lq2NChrfBNvaCXJDSu3m2rEavpq9wDZATkjnMKe2ccJRAPoGzf17lsE0ZhMKc9Cb
7XGfXCxQYkdfmK8JUpUmRgetF7A/g7lsw7vWTro8UrynilUvbngQrpiTOkbMhJzV
qC1oDyNffGP6lJtRjKqA12LNh+cFnIADJHcIkKnb2P7xmj/mvrUZJ3LEEtrFAQR7
WC7/VhzJE7cQ0ZnJ5DEj7kGpvfVdn/mcpKWXjkLahwu7BioWyg9lpcYskqMRGem7
/MyV0xBzfVsLkSzOOqWWzVd6ijpeje0Wm2Ti0AH/fMOXoupY4DolSa2hpbfAqQWP
4/ghENHnP+QkrMb6wpYLx7gwHrwgxqWHpsx+6qjr1lYNl+Jdhh3d26nSBR/yihNC
AYjZY4O7kbeY0+WekcFbrNTZOljRzoFR+X09QycWjeZKo9rBwAIzwPGdZ656yMBE
gtegl/LRc5uLBSmX2xS0aN5M4ofnJGavyAeuPoTg4HSVV0MrcyaMkAttEsQhMvrj
Pkvyyd+7GftJ7MtGb7lUd7GJqrwU9hUzstbNNJ2PUq7iHO/P9gQLHjqEPcbQOFwk
EHwW5IM5DNSK2KylzMtb5Vd+cmCAP9lFQN6MsJe5Q9vcgjIWwPH/Ov3n+l6qkQJz
ELcoWPKS21QoHmwpkoRK1RD5/vTcJ6OJukxcIn3WebFBBjuRdcOlSRI2bJZ6gUgt
OBfJk3vCLR7KmfS7nvsXpzq6JLne0F7mtGCLYEWbFrvMtnjlXS4fnzKlR2wNkzM7
SR0s2inY8DovkjOeD6etA5VoYxEwHX9AQnjHGe4va+t0D5xcDrfYt83Mk343Q4Ds
FOLppRNo9qALnIsFzxW3SX41RK6bQWyU6S60YGhK7Av9FACEqnXrCUy3CXgbHXpo
xA9HauaNS+cn5f3FzAU+mD4NXE+I4DtS58pV+AQBRqeUx2elFCxZAxvAR/TnQcIY
YysaSN83fJPJata1br64++sQ7DeoMJAuSC0R9YWmbS8+z3OycIfzSJfwHeuTC/b3
X5/qFCTNQPig70np702Jlu3N5mOW83XJs+9465U7H0wyZoE0y25IdLYetp1sWpt2
osvYDBvrY/DH4cXCyQiJI+J1JYKmbNAo7mtKLu434jjcx1Y89vos05moEw1Korri
r2V4i5AU/PbCEcn+aXOdqJ9WQULqeCuo/DprxGmkmwrVJCzQZ/FYDb9Op385Zowu
pFd+U98M3ADizfWIhtwPLlWzj0Oon1CnVdy0O+1jzrEjDVoGlVDXV2y7Lqz2Wfmj
973NBiKm6An6foeQqIQsi6iv0Co1S5YS3JNlvZga+6giBjfbjfis13llNczCAqAh
2J3VsOSbH4tiMn7WGLnXxCjJHmAEr1ogZTqxlcZpe7Q02JJyTHjn3ZxI0Vq+CXdE
9iLQIG5c6kIbDfEvbyv0uKZGoBlHtcfO/vHhNVWAnqAP0Qgzm7PsAXFTcvNFzzbL
fCPSYC6XXfPD+8QH1KocjmCwW244HQLO3TcnXsSfeNCtOwf6eJUrUvfm4n93c78u
B8mDU9CnNYwTiNiwDk0BVMHDj1yWYYeyRs2XOHY2ApX7AWQ4L8ByWgxIe2nnrKaV
2LakzUF2ij2Ve2+tuorrLnrZ/JsHhiEzuCOLQxZSOMuCMuE9919FuUulWn6/PE3a
eQ99K5TNojQeH54GgVPHlWGqsjZTuJNg/QsDibi/4pzfp5Ts5pz2CQ00sAB45b5i
+VcAtG/djTBmEda3rdAF79YmYLsE1d+nEkbXFSN7+Ylv12/5YVVudF8ovVdD22E4
9fqjiGbvbZhhRR+JvbTrwz5y+ClWOasGyCAsPwBBysjRUbTFcabac2Ou1ti0sl2z
J13hDGHajQwlR71+M/4lMhve5wgIJTGYMmSwnULHRQjQ4H55djfxqsnybdox/SCF
UlEZaXcPoCk4z/ehVo4QfSPCgaozWrlnfJRfb1aAcf7ox+QUpjjjOatcVIrcSs5W
FiTVw85jrhYY8gDnh+KDK1hYsandJYI0JemY7ObXH+diZObaUYNwvMP8NeNed0cm
jxFH6k2P7M/gNuaOPRcU7JPUM15Fgpu9xTk1Az0BsSHXKZs5/CvbavwXyCleyTOy
CpUbhocvR48X31lNCayIt0T/5VD3q1Y15oIb7O+NKK8Ouqk60fYCpfHfQN0Gvgpd
sjS5I49sUoE3ODLapVKIePFwo2BhuAUzrLLkNFUuPGRLp4pOUVz9GHW7Vt/CqGuz
1eHlH3dXq9xiqccyUCSA32IhhO1QCFXW2Js4xSOFJjBEnzxgvwgYdlNKvt+WUOfg
4CVxDY5bpqTpzfxPCwAlomekombU3b6j9kT0wXv4KORxMRsnBSMd8j9PKGQiRgZ5
Gd23fcWvPjJDcApVjcP8Km0fZU8lDkoJtAQyF/Ut//pMHa/8ib20IJ+BmpL9dwk0
5i109k5TjPMX9Bm4CrJlvtgx67k8H1LQ5jaoKaeUmU2ZBeEO/07IpzlRyFzoFTfj
Rd+CmQ8Nfy254oWOmy1LXkkM2+77IX+bZt+kvbusW7Gk+stjKxle2UvgWj7fQsDq
fhFbGVgxJdrvEADAW/OmCMaikFNk58OqpI1tBL5Nx54QBfmsjwYCk3AnOduy2gbl
pe6iKRLmzzygym0UJTDMKHyZ97vW+zyBAxrvPojEY8HaW8za/3aJHWKL+1lPXALf
E504uNNdQxuWRMEzwk5hkUzWRjviGAKM/YxgSIWPbVWDAvHHUhH7KeTdxEbasyS8
DCp1DoS9gynQYyEIzBlQeu+UVwhEu5VaXJDNCas5PfaArJ9T7se/DsqRTv5qm9K4
x849v+7iKCfH67dFzJDnoqPGZTnRIR+iOyrV+LcdyA4CkDZLRcWW129L46roY4zW
AVyE904IEZv6CheDLpGZiV1fs25YsBYqdNRJEnIGKfxafKl8Bq96h9MhSoMMoM2F
+HhLZ6xd/V0wIwD47ZnWzwaNMTB2ZsUvZCCcYOzaWcOva+smRa70hgTxNtsrkbje
AeTu1Xjv33KB00kpNddXwCOE8CdYN/hj6Tn8piWz9QGNv42ALTEvJ1XvvhI8AkbD
TVMTW2O9iRSSfQoOzJ3Mu0NEZkZknG6nmUH1K7kR1KSrIWRscJ5/lx1qO2YpXKsK
FFT44eQDJt08HI0vG3pQXzFXWwF7RdGWaC6STwt+D7Fv6eQ+C87XLtf51abB+so2
16/nagFpaRlvSgmI/+tg0tlutsLhe3OcR3NHDRS7afJNNZ3Vd/yFECnWtB/Os2K4
9wpO4m1fapGo2BQyIYsRlSOfItnwBwDUxM+YEfSkt7kPuqxOqI2TivNtZRiGlgNj
i1Mtz9lJYjjBwlucwG6fsx+8alrLsAPR8sRcvrOBSFE1Y/2G9IsHZVFkT2FcIVXd
h8wy5wKBe2xt0AcSPEjzpP97T2RdC7XWKxG6lwRyQIuaHEFku1ktCI3pfbVxqbR9
o3YM4t/R6f0OTiF2OmOdSBtgEBymd/H+dBNnHEIcDq5yOuQxpzhv6gnx2FeIIW7B
yLnHi6JGyRzjBpaipD9rS44mLqDvGCD0bFa41Y5GlafjtJE/Cnq33sF0KIROnOnV
1wk0wTWT0Kalz2yXMeDwYBuCuw+4trSivxkJR9oj4YChxGxfsKai5An7XNYuypjN
KEmqKIrs0jYG1eeCHomu9q+mEoXw3uhPxhMSe435Z6T6otEq/evEYwYhVAZO9MUe
DCSFATl4JVDViM0XNIAzvmM18zvQR7edcNAYOrE5VgZX7eJfcxIbAE6j58YsN+E3
cBYJ4A44XUnuZk7MEEKB4w3GNpAsEqXSZJc61mtxAPVivhpBISUWp/Yw6kM0uxad
+muq59saLa+V0/OYL96yJlS1FA948GN8V0/unHsMXZHxoi9JyaXYq941KsxMSw2R
pToP/EzNWV+6TiGaIjFTAEDfsocwojhMklJMUSXM2V+9gQzRGVJtww8wIRwSzAgB
WgrHegcOStZm76r+VMO/xWetTtB3bESXzcF9biVe9fL3/64f8k+A28lKmKna4y/S
ko5HvRNIhbKYByh9BQ1EINTBoG0dcNxQKbHT5GmyntKk+sZ2VKoLCLg/tgtBCyMJ
f0TzFQnqhatyDYrpWWRF+ELXFlUQzAbJg/wcykmORP9eGydThld8vqGjuIx2390+
Ez1rRQvgTDCSIhL6gKajXcU1aVk0+6geefnBTDSnRG3oQMQr03J43CYJ8LYwyku3
3HIWppWJEoESs+bfUeEdfK5u/s5KpOktJGAphT1RxNX2PbJg2DfynPizCkSXMZJd
VbASdutXhu+/BGts2W62aOO365vU99/S629gnyUvXVlPz8Dq6vltpQLn6W1u70GP
8lU15LV2Jqwgvdl37F7gGSyoWherDOKUxYQdJip6wT0cWlrKuk5RQMDvgvizWnKs
244pq+CTgyzLsY78MKXvv6y8NG7IAV4ehCHYGEHIdK37mzGaWLjPMlhFHx3KkYKc
uF6bgVxHLFuAJcg/b7ufskPoCklG8peT9e215kSZpIlo2OHLsL5IxtT5vKFsEsV9
EMieg8rNgPIcIpkE6ZTuJiNz0yi9jwWVAohJRes8nplyXDOSL9blVc4HAxqi/Jt1
z6rBhWbQhPlRisAqaXiBPigprSG58O/fdvFsKmjX2ss9JMq7DQ3/z4mVdAroM1Ud
6yUxJff4DZLvOLRNOLNBx1zDMjCmpBLytp7DTnPk26osKndtPUY3i4fYa+5W72JX
Ta7rMDwGlrsAuNPymZm+QJ6qwDM4OkCH8AglQXXcEtHVqjGsvy2XPYkDmbuUU4t4
f/ZGeb/vlOjPDgWe0Eyk2NeUxoygNa5dnrViKYkKWmpu8rOjbTqngoet3R6hEkIO
/Y1dwO+J8pBWb41a7aE9iadw9YpAxAE/fzb1RkDKXHjQUlkJ5xFiergrO2GGqIo1
8kp4G2J7ZpPY/QqyiWQipjwM0O7flci+E4TauXgiylYxISoD2+eksjXoi2fp2o0f
RllFrUjR0VDhWjVuMgCdCtiUBiOt2kfodGf0QtKdrgHxrsWnbH6CXz1Ka3jdIVt8
/NjGNJzjNn0eI/hHLbozwlxYADTcmecaAgGjKupIw9Rn7eAt3FTSjl6lfDU4SQh0
HLxdblQEe7MqvtRIYmlCsCO3BazE34myGU1AxSS1px1Y83IGLDwU8WTpAgwO6muu
47p2Rkf3oZoXoLmHAdSv25eS0jLqLA0+Bsl5IItTeVq09Iq0TGuubOR7fRsLk2zG
7D2iZHR6g02MTfW0dbafnQIOrNSm5b7KWDX/nX6JL8QIBD2XWuBeqKJIVMqlP/BA
XtrlO4vLjpiSV7q0s5cDkT9mtfeLenxEknlLxKruNtx4DRgQ6IYxyisYVokONNZh
8GXNrYO9oaJ0wjnA2PxynPxcSOn5uDWGFUz/XjvgGUtp2NcVB+IOqCWU4UbLYHKV
CotAx+sJnBaHj0IUESF69S0LshsE8yzcNKzyyBPP4VFMEmwYeCB8rt+/Bk6OKIT1
LV3+xfCBBdnvKVIqClpqRqcGxHuuvHl1G9awHT7IXICeE4xANzlQvm767OFmyQhm
cLDqsjNx7z6V8Fv5oG2E49Uep5udm1rd/l+YZ7lcTXDrYFZZRYOoKAQE+PsxlTzU
Cj2eBQPZSMnApCZxka91urVKgRnEiyCktDyRIIAHedpFyMAJUHtA06JRM8iCGR2b
DlfR7oTWNAzhrqpDSzct1C4/ZVN7BfbZc8mb+N94l3FvoRHWpx8PMtoIG9YqxF46
d4038omtWmbyB4p9G81rB7m1N8ghomXjYHg8u0UAYrPdz34hqh8Shr+asUY5OFwl
HAZtaL84UOR6yQj3Nzz0nF23A37zOKwzzmzsQh/+mw+TPQ7Xjo1UFC8kd6UxmDkf
hTPfFHf1HJlC/n0f4Zq2sJChwgdOjm7lcHhGWzkwJCGwrkyklbDtT3zTbvNYoYEF
7LmjHnKsUJ47xnoiZrrRgnCsqjcuaQAhh6d9KyjvwM/zUBFiGtOLzoeYp7mRqW3V
UQqmQu0ko3nXAq4WOP5xP9NyeQ1yOv8oWeoFTaDZEH2zbzgs1QbiVcYxdl+jgJmy
kKUZAR7S+QX1HDz0fhzSjAW9G0sQFgeOkwwz3OrEiSX0Su1eErZq610OMorY/4HO
zePTcTf9qXdWh9MrQ29xVoXqh6B7cTAvr8O4YgAwLT190gK/f8rSzVU1yk+y/sVo
L34du+PYDlWUs1BDDynDV50HZj/f8S5a76WyhKelMTks/31p/BYsH3+r4EvFWt7Y
V2wGM4US3tIPFQ0vxvQkGJCJ00Ka6+/tqS9kbvZr7n6qGzNjV/AvqcJ3uC9ww9G+
4CMCV8udNlaPzCa5PYJKS10wtJndfXmOq8t7YkiSvzCBntPNxVgsZPyvpb6X1jJH
v6YKkYrsuDCRBV/zgfJzZuHcEJsiPKaAA5/4zsczLzgpCfRSZER8/zVNI3BdjYUV
wInw+F5gjcsUT/txmuevAxhOtgHkz01VRlOLUEYBaJq47Xq+6QodiLSnlceUIX9p
0Et+zRAzi8gjgVgAINyXsAnrclMDZv6whnLyfGZnvm4ojWTAHQ9d64CBkaIANUqZ
yIFZJQzBsS7OpuCn61R1DsPEQJE/6YNhiUczKgCsiDApyJ4jt7lyFFPiUxdmMasx
y0eOTD9nYm3VzjrJdJPqPfERapcqTAh+l+B7qO1VaDqRUWQ0NqvMiUbWna2g3Dij
EHetEudtJgatYK82xV/tBfekRqDw8ENtQuCHn1Y3X0Ejnlbjv5oHFgUZ2jctXmi/
vydSyDA795Ewnum9ReX3Uzf1iyu6oWLRRwyJ5pXAzz7lLzgX703RI62dpa9lrMnQ
HpcSJEb71FELlQLZJIasG4k5+5I1dVZvg/rzsVmILPYgsFoK4n2ZWl0egxN6b/gv
fUHD3AH2dTY4+cxcd8d3tyEMxwF3/jQmj66ZQae+64incfyKC1fXwFEKpkmJKIpP
W4VR0ZarLF9K1FYbYj0oQ+ONcw2xdwfTz6W3uymx04qcszfQTOL6inKoAB5Igz/q
3mW1A1jucuNM6O+O/a5fT1WEydvRaaB35Gsvryd5QN+03Pqswd6z5zqHW/dmcPti
jffs1L47eArq164vbfFS5TCxdwRofFCaiUasK2qSQ4Uyw+RWBTZVKQ9BeB+u7DQe
QXeFjQsSlYD2GO0mRNwOgX+tB8wh1JeNSV7l2cVLDilJQoTteyJUWyTwzMclE3Bg
ufSQqdToSmw1W3zFxw3Ohqeo+cgfLctRBuOkQYgzAaLQPRRmWptcrF7N7lg5bcqj
7MUKL2VI+BoF/DQq0aEkO1ahGfDDkYRXvZZPV2KdkHpTCF1Nq7ijOdtBvv0CJt8L
Mm3S7Z3oRqdQWT/Gp2vWfPJK9+5bPMkJMfkHeLYsMhwamL9L5UvR3Q21ERRjG+ea
qpcvU7emvGFma1rYCLjhv5r0J1cHttBdojpFFWxOVnqEI6xo6qsL0ktu/N4oI7nk
xu2mJ69v/6MPgJuvXFk2IVRy5GjkxHg28c2MYF0rs7k11hMcfnpAzj5diKd5skQh
KL4/eh78f9r2d9LWNMi8CeP6CI1j/dPEudR9/ctacXZTjwPDI+N5pIu7wRV6EDTO
sehZnPA96/AqSbGi8lmrWkB+y4gv7HF2w9vWpHQvfRx8uswMwNeNmpV2qpjC5K09
fNcSA4Ipn9QAzvLYJBToiH4xl+fIqbk5GBPA0CtTcYa8fyTsdOL0EtoHaGOrxLd7
VtO6dAvhQemolpt1gPe6duspXOodhpS0S7tjq+plzhiWKd1DgoVB76akmdM6bMcY
8iFi4koX9p9q1oAF/XMU7ZhBikZ0dl1Q8oDDV9ZxFXZDAbRX8UqPKLTa6ETmwRAm
IBXBe/fP3k8UsHnt18NMXlkTOxGaEsZb5Q3KTCkaeQlAPB3q5rj6q3yvuPHzZ8Z/
aJSx0M5sCGye3JLWMFnQg4XiPDWYdS1LEH7Tn40rlfJqKrvJYLvDIURI36Szi7IF
eqxQZyaonvPR6IkJEf1Y+fiLvzSt1uCI4ENF/3rFfhddKUAiZa67elGh23EzDURI
yh8zTsguVBeLDMG0Nb5QyTJbrmZSpZDa8eSp2vrNHSCQw1U2yFLQzt/zijTpw9hk
D/IF+7gZtjdgrnDoji/DXtW5sk6UF+aoJO9DkInVkCVRt1qJqvJj+OcBH0IszNX3
nsc0Nu52yUSuroyN05TbLEPkkUcSw6gJStLj7tl2baJyOc4h6/Xl1bkQGfJfF7Mf
Fk5VzY+pc2Ap78ecnyRnMnY/y2TsOrMQMUDxmQ1/7gRqp45UTTqR86s3ZEqfqPaC
rnJLynsT+djhF3p/201BqrUgO7S0jDYKBZAYab/lfswk5yxFiquoEYfVBx7Pp+NY
St32AHB0iqM6E5kAw/BiwVYowXZYGQ3wRnOWfqOUKmHH8xIwne4wDKRiDb4CYrXq
mMUHh7+8Y5nBgwQaTjzXUWpU997B7jSSb1RZjlNIya1Rm/K4fqXNkXGSYvUqu+2n
+QoWmCMp/XU/hVQCZJO5YJEkO4YaLqO2oHOxjERIEY4B8uvB5LQaUA5Zpm5H9q36
q5jDN7cLjoVthiKqYJC5b4ZglMFzN1pXUjihGz78D2lJEfLqZmoQ8W6XlCFlLX9O
851bJgEetIAFqy8JvacM1Hvs3j/Fp9uJiD0VY0bBVvO8s0pg7xoFaDgx4eWaQKjO
AjpWnHKIaTLGgUVw4yD/EO0Q/TdBLwQIjpJ26YnNkr0m68nsiZkJQyIsBodAGE+h
6/dCZy/O383fZEbi3krF2aw2u8vEKk5brkyA/55FnrJ6eawJJFTLIojGBMvzvdmo
C0mbOY+DMWL9/l5hbmBN8r/Xd48sLpf4fCQ9pkkqcMsXj7ZS2pbL8jWvnmeLztjb
v2XrjboJ0VCu0bTdOwLj/gmp6hLhNuYoNcURZowarfsEuC8+vMBvTacKherRmTq7
ETUbq6HCLylnigE42f/+f6IPWu6YcwuAePpg8VprmdVPncCAdsv1b7vAjqGjryto
yQf2+Eos4dzmrx8PCvimBtXpJCDS3MElvyUHak27cv1Xse/RwJfcaZ7dXjCkmrrv
QEz5mSTK8SfH8lPTcyA/wTyPduJuOHBTEfKnwOaYOy0jRsVtSOGXxUdTnhDeCfCg
QRjCb1v4RgUxwSd3g/vBNC2yZbyxi7e8Edgx93MyB4XDfl8tB7Gv7TT7hrNpPZgw
z/y6X611i9MZECLa9sUaY+Vmk8AXJIGsVM36f6L5Folg+Z+3z+0ZIYmR7qX3VX6j
c7Pb0lXfnmAWQ58mgdjTBOiIvIsg+eqgyaCI8U2uWNhdjTR8+Ht0QbhdzXIIExaj
uE8gp7dooJm85vFliTF2EAsuQv+q2sA8DsOv3Qwyj9cWeAqNMR+KbbIOvCJfQ8QY
WUIXTSwab9XOGJqqMj2RadMv/e6nfppF3Gk32SBPK4OI16NonBHbDK8Ene0Anqch
oUZDHcoEqF4eOl/b0w2QAcp8fs5UsKC+H56156/ohaVw/nfto0P1dDzs2AicloZ2
BoOTFvAlsQ93YMUFCUjYFbXTjTjPapBYO3sl3mONDdqaBX//NgkJV3IejZU4Nixh
AWHmF7ekmN2L6HMTDOZDmMUM32HtQmkOociyX8vIbLvPubLsd2D5cmnuz5Q0Ronu
MrLtjxrW6PqpJHrxi+izp8KilB+HBZZ4OVgtJax7GJNBGF/knYFsS3tCL2eyob11
2VW3+Yn9HZzp7y7WPSrnt6ea9ZrpUM0r8OWcd/G0CxdyqaDho377B+dJS/DVvuLp
jfbP5+y8wLHjM2NK7kEHTgF2BiSjTTlodQS5BPY81n27QnEB7lhpl9j79TxtErfC
Ezsr+M+V0wpQFa67YbkZ99NKzR70fWto6cCaVycGftsfZK6LXUXb8dc2gbV5XNCi
NvsEvRDD3l8IEaxWUqwYso8VL7ivBjlNSNplf76AasayVehnErdmQShHiSJRvpqo
WOcXAdmdFNln4grTxkk62xd209KQA9szWM6nLe8bxl8iT9LeYVBU5He3R5wmvO65
qc6gchDjgWB44Dj8cBE4vfKm7GPfvQsuORq6tOAroqxtZaKaqIAKk5kj5IVRswhw
HdIuP7mr0HRNXp8O78rkPKPs1P4Hv2nHlI2deDHSOiaTJYV8Gxnjds3mwrpJm3Ee
iOVU3HYcY5jlRFv10GE/6oDMEiu72wbFeEf6OILcl72/e2BKVpsjtlNEvr0nb+pk
L9Eju4ObaMYRR5QiHZzHCghgqb1uO7ahmpGMH3XcfGgdmMjJ+X0DHv/dW+mCqc0d
kXFedZ/hIzG7IWpmJ+qGtUyMzUZ/gGDoqZOlU6RS3XFy+eNz1i5CFM0Ug2tET+8b
c11o8p43csm6nFL/Ql8voBHQ3FK3yhntrzfBfofnNpDJpEucdK+J/P8XnYYKVnfi
ME9A+DeF4hHYN307SiL7yptkpxx82K1JSfRjMeQCCNs3JezjKzbBmqETD7UpGBaa
ygRj2ZA1k8RAIBzgCdUabhAf5Uqn3/wm7kdVSUbBmnA5GOHxpB1PlRFto2Wruw/l
K721+HEoZUjqHQ9HYXQ+0i6hp0NISlSYWYzi1XwfbN+KyQ2njWrp7kvJEs83XWdq
JVj+JEtF/7t2Vm17klcDpedUK4Jrp46lWU0617YFlBWHRB+owY2vSJ8ABCP+C/B9
B2Wsqv+ex/DJOIgHo+8OvoB9gWtiW7hokOd3srWQ164okX2ZWZO6+u7I/rrOjf+w
a60hRSahwHsV4keIS2+XY+84Y5Q+Uk1jZhlyp/w+oU11JG/nzLMxON4yaoBeNnKa
G86d/HOhgn2oMzWZKGj2y28/HyUSbJ9vGNxhkjZBwWa159PfBHsPZM4Aq/bAzrs9
FknPWmZnU2lG9b3lNXNAGon8iadTHZBM1ElmqV6V2HXEyhzFIJ+lVVE5dOkxuFnj
Q9rk7uLvLZqSCCshIE0yCRcXXxFKwqpS4//rHhvlJ/4yHToFOhXmLErjcuwjlfKC
LU9I+sOB3+Ut94AW/GVovSQaBFoHIilXDb5eMxJn7JJWDbjPHwRtkQL2onXQGXKk
Qe42f+LYcGyu9yCYAKcXU22GPUSGosvP8LpWjeYmmNNijudmRz0/V6hQXYr9Ff6Y
HO3u6mFhHdH5qi4MADmIlKCebbAQuq0mk7f1g2wfs5Syk0K6cw+/aalWOS9lx7k/
CDChJaXhV/BooAt7jl8BMGI84rh6jLUAmDg1cf1pepAoirRUTMp5MoWMWmAdXtZX
TYEYp0enKwA02UxVWoe1OBP5X9QPF1zDQRpabyECK/YbJCXRiNpBiX1ajwkNJWKw
IoVJY1+Ek/N3ibsG2gW6BjkFKPwZnbTTVJ3BITS1vWyUz866wXjrOIFlqDC8tLi3
EKkDbrOPPUi3fUErtVqA+I0WrWzB4pTkJK5f4I4Fe6WOSjhp3eHkxzk/Ota6bWJI
CadjCiI76f1F/9NvihrzjTLt+jxK595scUsjQTLUJ7eDz90bPdivF/q4o5TueOWw
Bq7iEDDUtal7ZbGbwM3UIcvEV4qB12zH+hINl88DCFZvOku55ZkPqoFJLqWkLr0E
su4qHwKFKrtwlWRqMFAqsfVhVYjeLe0IBaWOW5QZs07ppTV4MDeOVD0CDCX2JbTg
UUo0gaLWkoY7az24wgidYm0Z43Lpktp70nTNxOdeJLNJGLDJokAJllmAzr+9eCl8
vpbBfm7UNWUmB3r+FCVsxsTjAmuQ0cMddgTNwHSYomdit84UrwXQQzBb+Fl9TcJ9
0JPHgaSllvKwFIxkWFztHqBL0tlPEz/iwifz1yLsHCC8bW+7qSt4T+GWNSeKGIUH
VJw9oIHIcxsMYBhEo3eDh+388Gjv82HBprRb3o/56oQlm8DniXoskFb2jf/Rx5vT
dVbHpuBMktSmC9psIQ2l1xT6BaQOcdbM/Rlm3Prtv10gSwVMraGmEXwi7SYpNYmc
4c8qk2BZGPJmd/7RlQtWcAb9g7FORJnFdRMpkVMZ/SAfkUFGWnFDWbavAKzyJE+f
eaA4Zf7gGFEBgTPtL8UQ9gWVRmvDgybHZFiA4+81t27HoSQI3wzswtifAEDQjsPB
L8lb6UdF706D4m4A4ywa1CKcG+uU5cuh7ijFGTx4Llp0yNd9YjxPfwoLI7gaT+zM
BjH88XJL2z9dvH0w21phDCUbGE0q5//v6Jy0z19F5ga0ubQa1lBaPlon8itZGeis
stSG0LU1sLrcfQbhOeeg6Tyu1gt7K5DCA3LDTJ1TP6p+67Nctwm/L+kEpwdA+me4
WmkcEaMBBsVFYYVORMmhvOYKaxYXEKOvEjgZQin6rUEew/bbbJgYVSk1nIvW1NuB
QMYZMzSMMHRF1K1TaNC/DpEW/82mIjDUSM9zi/1tLiRP2mv54nnt6szdnSErzw0q
wZJY9GUb3Fqs0R/AqPOiuu1sWrol14ca0fafvY4E1yRbFNmC2i/Fiyin2+KoqH0O
jhrmzGqbHRskUpUxLviJzcKX6IushJqQrTjJm4+gCjnlRIRztBGvmb/BRuydAbuG
O61JoQhxyysGi4O/+1lObgbXjxApRlE6q6AodpRZCP0FKwcurMTyl3ovVQeg3a4c
6WxaMfildUZAEsujqBQkKpjcgLy0PPyQafdH7iZwiPUXh0y74U2kWvXHzoEOwu4+
bVlw5IrF13ONpJ93mgHd4oUk85OoLucY6h9KWsDZVoCFaKdVqms33RA2ZLi2KjaB
+5KHo6Lnf4gYQQ8uYj5z5UG/MmktmzQLPP1rTBo7t79G8YGP7HnuGlTORFdo79hC
nTcp8tecV/kLnB+aHQbw9wSL77ukWkllxpAj2zxqcSoyyV4tECXleaAIMRfZ2wYn
yq4QO+ZU1sSdJluN3YEK9q8/RCELlzTloaYi+8fTY70kWgwzEOOy3QMhv+RK9usE
Tok8a9GcdYEphG5yLKSyYl7d23w20dwQ/i5A7/AWpFyIrbhN9fPfdvqrt2w3f8Jj
FmNYPvg8aAPoRT8kU1IJZwxy4qc9W2veTY2amTu3MJLaudUulYwI/Q7MKNkNSHyh
VeqJgdhrb4X7B8l4O/lvTZbFED8yktZV7WzgLwjySF2hPEw6Lx/MRQmenewOlGWq
LwcQ0uMKac3RKixA+52YLzak2rQjM5V5teON/uATV1tWxekmcM7YOrzYJsUY9JMB
kfH06Xe63yrBpQJl+sVPikoGaEJNyYZ81VkzeuSNBvc4h14MAf4KP2nhKENjylMA
MQ0UKVSzjywBhxUJ80Npj8vM/FEQ2PXkTMqizshIOmSnreAFPm6o1cN1xnceVZDB
HjVXbqH7UTNs3H3NRAzr8z7QnVfh5cXlV7KvHhywkvGpkrEwv25bUxI2UR9EJyGl
ICEwuDtGYzrcvCEhPByXO6DxaQULo5IR15lNkoEnNgY0HgX4z1/sd2/9a4C+g6Kt
eTXJ6135EEis+KzVKT97OAA9X+e8i5o58Zkch1IIpO6Mh4Z/5RM2Ct5Romhp/to4
4mIZ9p+wR31tvn3HiexrZh53nzaK8eRhxkl15PcDfk+Vx/R4kilUfZWJ/PYC5K4t
aXgRla5bRfT/a/yTAYPjWBnOX3M7Auhl5NjwZPSw2JDfBTXIFBTbrOrOQL89K97i
ONioccaqjviK+/H1AI9MKoNd06TENOUCXGpCTq9P7TKx6DFb5qVRgzB+C/cdzfn+
KoYo5WcXEUVxMoUSHdMx/8FYnaNKX/eK0/bvFPdkKO7VvxmSfGyE+HBg3rgga0qB
DzMoh1+ef82ASZFLlfR5t2fxgFxUIxvTGW6Y/V8Rc54Dn2idtBERQZ4qgk41Aq0K
vIeEbnv7z/fyqC/1ZYRqivMrQs7/y6aaPBva2A1eBQMtVYdKGKLG/PYx6+3tGSFV
UMH/T7/v42dWh43TGPQsVtTwUPifgf+k7mCT2PvEOo5OlH4/BFsdZRkmZoVXuMpR
YT1c8+/kjv67LTmUMLqW3MA5zEwOA8FrnVJD2D51/Cq7PxwYNs1i1CsFZQsOQDWG
KFzX8b9VUxeGEaUiCCxULrDKMbhSAy8ku17HKj6NvFptsziJ1ofHfN2E2RQ63tVH
mz6dBTcwfZysBHjYvzjZHqwRspLWbgi8mIv1q6uBoCajl7liusvOjVMkob9l/dPQ
+Bn1GOiakrZNoN3BwKDFZexii8RHr1G2JeU8ZVDWmdfcylEUOzyfO1lCkZ/TVpQk
hK1yT5h2JwbafwaY5G21zCH1e/be/FwIXjj0+oZ8ADTUOba7QX9Mqw2eTSNgXfd5
FgAFH5ElNwpaWb8bhPV0VIqwaGfBDtRDzHSaX0KHBBzaJHxZKV07NPTjkioRXorw
B58/FEhW2HUiPPz/uR58SGneBI/BCYsZj7zdue/r0GKitTEu/Bs4kMXBvylryIPI
7m1xPITTfFZHFi2zRQh/3I2pnLovVgqkobPL0mo53Map7EOOmjSmKdleRu+WBwGn
eiJsIkoN4DpTrDWmesxOP39F5DF1mDAgGntomg8T1G1TQwCs2KpGx3DcSTknqMVT
tV6pgUrABUv2a0yutEOgYFpOYIZwtVmTjanmSuQaHQmtmrRvabL1rHWxrm1aShcQ
BZZJ/wOrsqoeF1q1dt/VVeYcUUJIWCuUWRhsRtIMsWybBVFny0moyWzmGn1GnObZ
l0G0K/HHYRzAzJzhsu+bC9Y55h2RsV4USYXInsNM2sAGVSlp8tV0O8ehYgXaWvSM
p1TQ9CbamaQRPfz458w+BbQ4BbF4+YAAIuxNRCXqUHzojcfvHH1Mx8KMbR13yXI7
vTcify0n+alUaWnJD6fRz6174reH3DJXA4GAQ1jZTsR0qwwJbgcbxX5SGnbmqtqM
Tgfvx/Kn4059WZYRQ9jnqqxqH9XHgwPg4GiwpOZ+zbv80GhWIHyys/svHD9hnW80
3CIYpuBlTelcytBVIQSL87AII6+DO2PLDgmI/rBEfszoFnMZGQwJBgdzJ1TC5LTz
bxncN+oseC2xW3zPDvSMWO2GsU8OsgXSjyA+xquK08GxKg7NT8Q5GlIfMESDS0c7
kzWzywVYcapCiuhpT0fsTMv0Bo10cngICAbTP2ca1oBOsSQVFyu8P4vuJbFo4HVW
2ND8l3lcQc51NuYeT4REc5sz4hNfdhgInz0QTkk1lwJhZyB5UBI0Bw0oy7GYcA1p
nuiVHOp5IB5UmVqgjqQLj0xZ3MnAFImSnC8/HNPSlcZzJwDmpUaMYfPeOeyw4D4g
TUrlK6lpUl5t8PxGmdm6K64eIJryqtK/qslIeeAiS5exExDS+Lx06Ot/nQmujg55
yuTL/egc57ClsZX6c1J27aFDsc6Oqp7qjPB5s0aMgyOGfaw0W2XWm83FX70OBNn5
G0pa9YAlwHD2LgydijkFirA5wfhc9M3Q64ovupUCRPmfA36MVUz03mVRVUiz5MvU
63xe398rxnuFLp8lUIK/8/+oAmHAoOozmR1prjIPTPsf57+iTDl4O9brak+gJw2V
Qsgx0k3YvoMzC983Q9HMMTTRb3OH8AyCLXY94zKz9/4uGCk62O8O+/FUNLsIOFrj
5OrLcfhakgu2OR9hcOwSiSW0ofBDzUml6cHtTC9JtJtp74Y1ICoxR0cfDbQW6KAc
5GRLTqnMQtrepi1aMPFyIG+0+1PCfdfTCFvjYGc7160/ApqIms4v0IMh7KddyXWA
pczdG/ftDRLLYIdRfH8SDW7dbkIho8y33SdbMhcAcApfrAZFeVljxjNPRp4GcCSR
dP7lPU0LYkWGILPkoAAQYt29cPDD43fUdYNY60yXi9hgIAYyJGXqVzQcx4jtwX/8
ghmVkEOE7nJMjJ0rK5YdwijeG2sdKv2BNk7WoQqin1tdLm6KY3FsiQKpOKqGhVKT
AHLI9e0UI+2iT1CAkx4nKGulN/xjniR1PdEqGH7HHThArL/FWQdEIh2K3wIl//WM
L7GsLi10bKvwhcPJT6fzqs/QnK0iEU+Ub5HrIDfgXhlIrtQIlU4AJfKTZtWOn92X
lRBO7Up1pdp0s1hfiNdrQZW3c8lt6NWzoHAhBYeVGhKgGLOnufUxmfvDUD2PhYOG
rYL0/yNipq9E0SYpNW/i0NZCICuaDsg0REXUFcclIk8GO35ng3/iNuk2S5ndur46
Fta+wV+p5kaSHN57EfhdunrXdkyrFQg4h9qd+UGmMp67x0ZmiRuoTJKzs0h7c4wr
RTCnebb9cf1cheVccS0hwxUAm2C9/D1n0BWdZAMc42EiDS+Smf+cz9s3+JQXNIMn
hneDkFRHk8okQVfGSGTvb/8yhcfic25VDi6S7hFn/KLX5vGO7w6ZaHBj63LPeeVY
1Blbf2lkALnzNR4bkrzrHyX6IFgz0j+mHV/GAgE3xbIf7ehOGT/5tcD8KzvHe4jb
3ux7cfxg+ZQwo0ZI1HKEdDg/Xtpso0Hyq3wJgo/gFj6pqKP+kSLadQeU88r0xIA9
c1VTKGNhiLSBLVUGKmdySD4l8mOGwCOOjPfc2XeaHjJNPHdXGx4frraptQTmfhdj
8+mpDJKvIHYkYHttkYKo84ebp3Va14mJ8bIQasJzPw4wnHuHMQ3PPiEKs4W1Ck/f
Yt/aY4L3VIttOgL5Qif1xq4h1VrkbGls5wo4alOZGJLPMqM91dfHrNyXV/p3frOD
9hZhudaKCfQTaSB41JhrXMnSFARG1XfyiFTlHWRWqUd8GyjuWCKeQgmbBaq6J2MQ
5/DeHsXCiNflA3ag73v1CfOsgJFc7Rmvu2ZQ3YXCMsMuqXRddkVe4vQfxC/kpLZ6
Dz4sxnnHh9rdRqSG3LLOuRIyEUIp8kMOulXK8pA33Us3AEYZvEwR3Tzivi14XbNq
tz9kMqdO2TYlivwI1233vOCPyQ5VlKiwOst2QjYodgPjPXRGUrOoVa4nkhzKfp7b
dyAEXfaNyRA/rgvGiurcXSI7hpTHB4Rcblb08+kv4LdA1tU+M+udvt2OKBIE11Zf
tKbslVdJP6wMquU11pMubCyZ+NWhzWgXrgk9Dfgymt3jAvFFYbht7Q1cuWW6HqAB
UT5twb0E4iBgfnsRlzThNsyoPaJgCSLr87VGN4DdcB529P3gfaoEqi8mewpBsT/O
TUcd4hpK5U0sfp0NcB1xu4MU1+3gg/F1PDOu6WhxAdfjn5gepw8N54RqRoPWDjk6
JaClh87PtHSzXRaC/buPLqpndF5iLVd8xWW5s6CZ9AL5S49qPN9lJng3a1B0UN9K
H2GpzR9BYazHmkmL1ZFdL5IxxmIaxToK1nG2YiwcwezJi7WWgQj5VuBIY83s1NZi
gcKC12ZBzynTKGNa/NLjjQ3LWGpdqaM2CR1JQJPhsKl+r2/EWlnTkUchSmrEE20O
12NPsNgIAiKu8xsCcHOOkuyWl6l6QuJCswfCa5mJGjZrTuqOjdGxW2mhuFMSZGoN
5JNkwxI0OXIh+dxWl4AciA0urUkTbJYLFZkvZUCtURakhzbHoq023baO0unZ29FC
vsJ7L0tzNTX5Pfsr2Qr7Mp4F6GegRBwh1MGxlMSEs9T/i1m4mHtm8oqjtGLVflzO
VqOTj+YuEvDylgVmQxhKRxUcvN+ciG5Tnmew8uq6PFzoQmPkwM69FGy7GF445w1r
229si58AxanCPMxTFt4CXl4x3D/UcEPmBXB5sVz1CxOYCnVIHrAUf26z1EmJFGh3
S4pDwH4/5CPFbiCa8aF9RuQHRARQvNFcQ3pezEkJ1H2T/bAcW40GcW3LQ7NfihDL
5JSM2hP2t3a6iwVdVxpjUu33MobSLyipKPe/qyXtBIuaCQe2/Un4/aGT4yG80v4q
raD6ETs9Zg+Ow80svOFsY62uwuucDlChMw4id8mQGS99p/SbTJtSFm+mwJ5ITQyG
pDSRsF2FCtl3ZZcmiCMdaDvNju4woaIxYXyQ4RNFvW/qeb0VEeK3MO0EH76+bPKn
mjcIajJePEZ2g/02/RszT+kEtt3xlbT07buauXjAcbeElkMm5avLaW5RlqOqW3qm
3RsTw54pdCrLHyKwbnbDmks0VjwciLWUlgddgUKu/pS78LRkW+ltwQnJuxfuUJWP
PGszx/sFhF005mWJS9Yrz6q+a4JuYoz5/oJoYzVeelhtHvuaQJ0PtSD8CzgbBccC
BVADOl+gFE0Fv6sZzNLVBNHELV9sUA10XWlNzsUiKI6DH6S/MZDQrIHKqjDcXKVC
altR1EBJOpYBYUrTPpQSJMK0vXf3uAmNmtc7VfsjNImFMkkL3kl7UvTT7Lb/N6nx
T2qFCFwaPBgGR42Iq0V6OwWxdSkEd14sqDu8f/fZ2VFAjk1WSnumX93s3usyWp13
WL1Kr17yZzrELMTye+xQ478G93Bwk/bfePj3E1OfiMfVG91kJ9L0sYJ/mUfhKhf0
gWk5VwpEtq7Cd6SQ0hWXZ1pVo8NDwV7h+SM0V88Aj7+/jjNEgPvDt0D48Rbpi6SS
ugwDOoiXXWvvfZuTkDvts72pLaerlpzlkgQdSf3qMwANDqlQkQ/oMeftHnm+cq/I
YXuvKFUgnkFN2DfiAAwxMfQsQYMmeLjXjEJhbTQCyyT2ZjaABlXBIaELhuSecwXO
hu9MJNOJ0y/b4xaVDgCpev0dsy05L2OsrNZGVXpCiFXG6NhN2pdOY2x/Etc9nxxk
uJBQ53axaCyjidz2+G7sT8YHoHRsWSTvC1q0hsBLN8NXcVh+LPZfT1TviYcouDiv
iBl36W7BCDXzIg1dv5p0vsUmLNV0LDOsT9SIxB4JOb51VdIsiJ/TBvEybwnH37VA
2zEFVGn8xuGYg9A0rNtHj+6lGrV+t6wuXv0AWgRGEvl4hMBu+G0GCMGrwKHy2ugJ
UgwOziYbqvqCwEvvHdeJRYSx1/vz23DrftATVFS627i21exy9FzTDSCmA1hQfFUO
ZF4/wbC6VuagOjKWUcs1WftMYR+EOzfiBOx10cX4RADuEF6sBjQBdpVMDDl605vg
SReQw+DHk+WD5MxwDWDoaj8R/sR1a1L0Uo1xtrEyL/UUDPOGslkbskR+Ew5FLs8X
hL/pnrSSGGorvZ11/M3Bq5bjxe7sfm0K92Y7uhcnRD7C3hLlqJccSWZ+j71EevIN
Gqbi0Ds3NBwfFEMRqzzdVYh6VwdBv6Xb0HrrpAdJLHqaYJGP3+9nciThbTpg8Jv5
VRy0n9lqFrqgaEqJahDUIiNeKFPHejhHiwIXAvy1eth0oIr5mZVqs9Vo3n22PjMB
EL2CoBcsCfBAHfgh00j7fqEabvzwfDiCwbYDF9sQNjicw8YjOibhpsWDJi9Ei6GF
XWhjk+oGJDlwtAfE/mTbIv1xl+PY3pIfoo2OBqtQA1sjUO0q2mBSmqigRQRMxX/B
j1rCljYRboFH+viBvmkW6ApswfqK2b96gXhFSZh2TKvhY4vP2ZR+SLdCAyuWaQ2l
elu1VNDqOB35z5V1LfZC7rMWCWo3XayP5hsG1fsKSB/SWz2CKXnJpEgK66aKv5Mz
v7LcFWJDPzz2FyMdtJyZmr4lfmPS6hI/d35A1p1F/sTgRPUAuc6FABoZhjiJQ5D0
/LpU4Q07agm63GlMhdJ5ogAUFKRMXYpZhLHPmdTT4+Bb9zgLi3FRZKAI7M+H6KaA
xECwE3pjSxSfdPTK4F8x8zUyfJ/Sdhbq+kJzhWTGq2O/tzPx4VZjeSGrl+bsPop+
U3Txfu26pxygUiU9HQNc4p2IIyUJYm8nj62xf8X2Ialn+NcfUbzFRNOG+TC+3zoM
VPuZmMlRgJH8tTfhbxtcV0LIwhXCzWUbZXntHYRpMb23OPs970hVVqKqHBStnzhh
M2hCApJLOr8131pOfN0V69O/jiuNrUGSYvloIX7n10zYC2g55eEevMYrjnB4et+p
IH1Fzxk8LdsY6pc0sYoMBpAmHrue0njnaF8obIHNIjhLsKiFTRtDv4/b8TqcR8yk
AZNA9x+b/5FsbFm0g+u+jkHbxSLIyvrsfwqMHcTg9xwQSMqbP2rMhCCdEkTiUPvd
I7sVuXoTs8Dpa66G0KhUF0BO4XkrRkfAz0VplqlVByhDY731Jiqk7uKlf8U41Ta0
ZLsK2jXiokNrNRqgARXILa/sk1xwx2RNyZzfMdBV+2wRTYztbHh0fXQe6RS9IQIC
2RbF9yGuYnRLvfFXGLbh7krFcUKsENN4Kr4Zh+fTq7nAhd2Xk9siTT/kUa2JbABa
G8J5SiI5UMQvzoRVKcjRJC+9S3zhgbvtQZw4Jc0uEo06p36HYMZ+2UrJry5MxLq+
15gy86ToAh+fo4WRrdiStVHqFQ45uAfrpdPAZq+PYhr82GpCn/QbNSS01u7N6mAF
l3Wx4w59QQxoH88eEsbG3MDvQrQD8KoqMy3HIacmFn45HRN1qRDTUDQkn2Fp9mF8
68xGCeZZdlHhbSEn1G+Sr9HJDxpBwkhe+En6YD0A3j3PvIbdxlMfZ9FIdLDIvm/d
tQthj2O/Yh1sFCoJDmKg6UcxYhTCKUULR8y7O5OsLrrGz5e5EbujIn5sexjUf6EU
HQL69Vj+T+ggXiYrUUGUUw1aryGdJb/r/3OSPuYY/VLbx7+QcC5Og/cjNgC/rwDj
S+CdExYQSsNmnTM5R1ODNNP20e9gC9Nby/4Z5drDwY9EkdR6VUrevqfKbpi5VHmf
SQ1B1V7nkRIHaXN1N/0VhuPv8HMa3ccBQ9bXABMiRilNnP94VRPxjnv4XDnWQBSa
JyrMBd2g2XgTrPBET57Gf4ssN+LfuS3DGktqGjXqKicvYZ8dbbzJtkR2PxrP3L9b
TrCSZhkSELbm0kP1PU9k8iux1r6H2bQGXz0DTqu0dHDh07T4tpUwQvcSz6q3zwB4
ZsrDkn3LoipcSoeoMNaa4SOwUb1jmD6QFM4OqqDjiebb7AriZ4kI/S2+8ehFTWI5
zEz3ydvgpla9zYuYTfmHaMCP5TGsRsAx7M9ne7i89MeJU7eu0p7qvHzADch3ZU/0
TkEM3If/1xAxoIO/ilKIyUISKdG7BqtiK/+18YkDnk1JdwbB6ZtHEhY3bkeP65eZ
2diN+KUQD1FshNdq701I5AYf/kRH+XIHyE2ZRL3VX1GV8WQnwp1VdeSUyswb/kUp
osuTnK0dxZ70jukGXNjyhXwWEkEkPN+RqX2RoxVEQfGKTv/D5609k5Zb0Ur/qh8u
EKHhLy8uBC3R+62H6Ozxq500kJ8HI2DOLfuGvMw3MRZ61ue0HBCcuhGsNaLQi16w
Oal1GRDKyUIWF31Eg9/h+LDreohyDWGgCkXjtS7mf2M61lf6NMutfOa6igk46gmn
qEJnQ637gZ2L5nHjQlqWoiAIMMWZfz1DgVWO6vDb5DW9XVR5zFwMCdkRq64xsTAp
TDgCzPrVDigWL+jmeWTw+ngx/FoBRC+ib7mpy1WbLJqy+TE6/E1C3E+ps4TARrKK
XqKMBVa0bpe+LEanT6qO2SdA8+MFv/Ks4D0czv2Q/ftv0xAoV5vwBqjTq58Axl8I
CplDA9yaMLJvvTUYFdQUCY1urLrXDWh7a+Sd5Jbs7JHj1lojTv1QzKKfzIfmEkCA
kc5qKKu/jb41k5FB4lCTBLtlrzOi3R/zShe3Ltz3zObCBW8McBX63F5I5hGRrlsS
AXreWWhK91bstrZcEIl/AYG5PE0wOesvy0zBxLkPlxZU679sjOvAi/OKM/zprqBc
8pJlHUe+VbEmbE9wQ0JF1OmPhr+MeZ1rYz2s31ncgWkf3/oyy2+/6wZ3tzyRgJ4k
I90g0QPNMifa6tqwu/HOBYbXLC0Adqkq3Cbh6Z5kx6XPJY/901dojFs3HUEmAgY3
oPkLtgijbODYttHaOAMzfd7xx4VucjxAFnkSlVZ1gWw8e0+NH6HQOSgdl0cmy8mB
1Bp6u75zLvn1mY34W8hfbL7zaTyrd42wJnD/HMCnpcN7lfKymUdXLXUziZsx65OE
zlvDiNTgYkjMDYcDgOJdzyQa6masUV0UNXr0Ok/BgzKy0smmhrdnKgD2f1sicB4m
jB+mRCsJbgRXsEdLTKQI08gMvVBacJlnVibzKizm7Sn44Qrc7x61PRHlnp9orlef
IUozeFokwh/l7O9K57v8x66IDOa760vkIjZpgyeNWj82iTYN6GMPrHWY3ZTSyOFy
0PBThO4uCEcNxdiTg9FaUu+wD2YPK/IuA4OTT4nUv1MR9JiWsbSyOUzwUs+18AYp
zb3gciGSanXhLJ8UzjcG3tIhnTAQDhs+Q0Z9i9ycej7hGnvxE/gnnuaMYJtnNOye
pyg3T9ruEc6HjQdkj7HiT6ZgBwjVWmN38SZHYGPnQxSoJqb3PWygKC6mNzdSQwPG
QMn3zcyt6UpQpdEFSua4ZuGXsPZFfuP1U7tbQS7ka8Do/jXFEHr6g/kuvo2xHDMX
D+VNpKGXKcJJtraywByCGRf3WaGYuRhtSz6A+smMOgTLhFxYGGHkw8q14jHnxeqo
xdLXNPqaJPOHhY9CkaVNJbWFdPu7cx9XOuiTK/U3kLRiFyH0X5QLHZ3BWGHfzirF
DToIewXYWPjzn8yJhQ4MbAsEL9Omb4EpzQYwgeY6Ne+0oxVNCWDx94jcnOJSg/hU
zRgbs/9kz4Hg8SiOMFdPfRBNUJP2HHd01vPMQJj05hVYd7Tf8HdJE9Iy5o5UvjyD
vUz/e/WqysqOfO9wVM3FzJcKGUGPu3bE14Lh83KVjGZPZK1LGIQad9wRYg51/++t
kHzq3JwcAt/nSpaobqOdQC1ttsuF1GjAdvuhHBziVk0JNmxiWXJ/3B0x2SgNurTl
INJyO9AAaG7b+HZtM9ToYzeax3j9mVBvcNzt4jQWs9M0U0U3pJjm1kuCbGFZTNSs
e+C50pGHXcaJw13dsjExp9v/koGqVoFk5VCPWNUQYs4q6QADIfQ6x/spUFWhSbVK
PcJ1OqESRw44gtL7XiVC++rUrG3Hk/sGD19MY03aBJPI9Pb5QUMfHslz6Sxfx/lY
u1KUXQZhtHXzwHSU8ajYVQRqM+ipyuHRBKcbjE8M391uAhCu9gDo3PMXSzRVAWXx
EFlEHpWoocrboS4fDEmRNmNJqD0He8ECIHV1m2c7q9nP20UbxDiZEpoilSRErDNx
GeW5JT1LvH8CNRYFGJA2pf8rTsfLWwIi+fMQ7+ryftLRRyRl7ezgLZYpghDS8W9X
t+QZiAIwuReYyvtYng6ousR0NE8my+J2sQohnMwDQ+6g5kPyAgAB3P5FCfbfkpG2
N/XAWvgEGXD5F4MVbQRLkkEiRgYA1/kcDVL3xXh+hEa0/I0ejBDv5nVsamQHR+VU
7kbGkZbfgM1bwUiqSCWimxqWMW1qOc4ed5J7JHz/7ZVKQimIudpw7/KZDYg03hyN
2IR4gpgxEMz9oXekp0Ud8DT1oc9LVTPqrwX1tdBB9rEmyKvBynrcwJvOZsG1NQB0
iopSMnkDQPxcgKryGCIeclXKSYUIoD2B2DBQ2XGDG10fqyUum0lZPJFL/6PYwjrD
yv8Oj5ONBYiizJWSEUhpBNwnr0yMtRHHi3WsD/c5mCNDV8u6KpSBdJMCbXs8CwK3
uj15EuWfeX5aZvRGpnObTyvzPg3V1/hjXGPrZ3PKbctp71B31/IQ0Fxam00omq5L
O62ZR7jhLveqlrQiWlYyudqoRen4368x0ScrvotrWFA9ZNZXW+5wGoLPZxFrNJwq
3BcQDCdbTWQFYox4Jj7HIYtxoRO7AJLjK+yan4UPLQiJY6P37pJyU8eLJHZuMgUv
sYTqbGrRBcb/QvZIPiiQumxcAw8XSLaWkWJ8XK9A7VB/8OvveW5+T2tn3MnYFyKe
4vuTAlDC8xV1zPwqm6mW4B4DL0YxS62IjiybVmGi+oxiETxsLOX8POb0wBbBj0gj
HIu9TMSkKdz78iFJ3ccC/xp0TVaQJHkglfxHXOZgwAwSYwSeBiWi9jKeyPhY0xi+
/A+N2HlP8bSl6d0itccSFO5e85At0yJJUyP0DCEb9JDRjnXYdx3zeiSYaQxga5Dk
CDegJPbiztdm0ijdYJm09ruEZrE06QTrWKFtBeorIkXoIAT7xdunEtoc3X4Z9Ljb
6s+1xVvZMpz1pgxMQxWio809J1uhInXDLfvM6Xt3unABIKEyEgJXNGF6CjGW4PT2
NNLR57iA72XLOsHe5VE/caNPENFryU3W4J6eRGV44WX5rc2AwFvNB0NzBtwRwtlw
XfNAtlvUOF1lvE0xOiW9HS9BF9RZyIxceOGyYYspeO0oFtXVoEsp2E/xmvKCehN5
k3hGdBEDJPzJh2DJTw0Ea98//mJ1K4PoLqfbH34Xu7L0fKDMaNG93AUuHSKy23WF
o09p+QhyIqR7/sz7KSeWMYRdSc/NqyK32DobgMJGXoJbPH09bH6jsZxMAiEnTdlK
T/0w2UIrH5/GYnC8FDp5xuK7pe9Fylm5AfwRdJZpUaOIsKt7qKnp78yIDJcKofEW
7ZqDcmnC1USq+lNynWvbQw1Vg/8dAIsz8ivyVJyOwfMl4yfBIJXN/EZOCtmf5Qm6
B7Ch4AYF6sUNyBl5K4zllgO6WMxmPEWIBO6UgtHroy36NgWE/LprAjI2ONB584O8
+NMicSckJN76wz5STdC0b3c58IarCfwLS0OlIOifYhtUdYfWrpqr+thDlPIbKN1u
Qgp6B2fCutI1/Gt33iqDbArZnBxesPP2LnA/d5j2qmH80gNf024XB39slwI463Te
4MCoK9RCyY5S1e46JTJPZs5H8vXLD8R18r/IPZ7kI0laG1PTotmOE5bY+jmZvdGl
jcghR35Oh5B52bRg1eNWRgrTyJ4D7z+zTRb+wJZiaCWRhuJJ6hFz4zsLWECMEBZY
2HQutfVOhvexy2+ezitSWeYMU3Ogqhbl28EDlEy+aOv1wNmgvNDuqFy+paE6uu+9
zVkPteODB+mtPfzMlomfCgBLuwUYOWSGDS1G7fZCGMGaNUlUhGlBGsWmQ1FMID9g
Km3VjJ5NKMzlCPsLizORKKoLWXwt/4h16dAyrcJygsOKrOj5O9QV0eGe4BG8rxeX
QVOtKVVHGx0vCku9Y+OFXRQEWucFQMj57HmS0iFfQ77dCq9Z3s9eMa0X0YB8eDKY
yXBXByuHuUeedMwqElM7P7YdbXirS1G03yra7OO1EGFpgVtvIQlpDswsMgHIYeO/
94lAICQLJpq1nwgAy+hbd4Y7G8StxezK1alKZDU/Ja49csIrt5djRLB3u8J/eGVn
zbVa4hhId2kd/vp04q9Zy24j6gguBvCDapqVp8myKpvEkMzcWA2CSbqaoSzgMPt5
Or1baKpPRPsx8ecen2sks1cxCayPUkvPjgazQ5F3a6UyFS2s70xVP8+DnocI2WWd
Irr02uxxsnNTn+3QDG6WBhoGgPj/VKxPUN2famFHSrpdsoKqWpJfmwRmkYUuY22M
AAr6QoIzsf7xAnkGrxrcFCjf1nStBa3Aa6z/KTCOmfUTjGo35vavoHW4BEg29Ky9
IYjhyZTmmbK3P0PH6ttc+/SjgK79iaJ4vZPkCFQN/EVFlmyob5xnBEUa5wCQqLYw
vDui8szM7vDCzk9FKGEo/kzwUxZoAYvOmdcQJOokYZtLBkPLDr9B/unzdF6avFTu
vvr8XZz9AlkpvomgcDlXtgjmlxlcxJa8O8pc99qD5eVdDvda01M82CT5zx9Vzvce
eUKhZlQwyWAslHZIjT66SgMEI5efR6UU+OMtEtHvsIOyDxs2h0n58zlls2XDLB4g
3ahoh7hgPA5eXxfbsqgNYiyaSrFWVko4D+QMVYErUsDWK3/VWN66XR3TmO9KJwKK
I/K0dAjBOikT6f242kuxheTVp+BHiIXMtJQQ92KZq7WKeETVNNj5fwxY2Z0IkEsd
C0wMoivyAvWEohMiKQUdqEiKtTSCFipqIFk8m6VBjyhfi/MFPlfFmDafR07t2Aqb
3YMsFyqAtO1zRId3UiihWgc0fEfkjIP1MidK4lOeVyaTiv1/xDLseF3Y/fIIybyx
113gPc0TcYhA4La1rxzKtNpNeaCJze5TUbwMFYwFhRpzOzPuUw7TS/oqolUsIn/i
OO8xhxpsOXg0S/+xdWHjPOHgTrzkamxDwy9cEmpn/sQeaMebotVet0vv+ShkRDWS
krqYTDQU+wvD699C35QdcbISiGgx4E5xy0Ob7vFMIGZcl9tCMUmqBkGeRMR3tIon
IKz6RGRWi0aVEarco6PqvPNvT++i8xW9+oZlwkCLzPvu3rtGKNP8i6Q7t6LK1dCd
Hp6xTgnkwIDdQ+2mIRP2ih/r+9ehkPICTlc3snjmqJnVsXumH+0RqQn3vNnoGL31
b9f2HnsvzAKn0eTwXdMjNnyfDPxShfY66XhG5qPVe62qNj4tZm54uaW/IPg9T6kO
Ko4daSp98Tgf7R2KNAmFZAGfJgPfaPPvvSJ6roXqE+bYE7WJaRYIxAuTiWebJ1SY
DFMO5koFVqpXnHalaepVHCfeh7R9hmEBbtVQ1bna52WeS6fXz7pvPELdHhdMJ+l7
FSWSNrBGD6uHH2mLg6Efz/qu3W20J4daifI9ntD91AMUhyMKouznw5/AYl2QMZv5
KWO1WkvjeeX3lfA7nO1g0HkU46+mXdv8TRqB9kIBJYsZsyUuYcaFh7/xpl5Eo8xA
7wr1kqcnZIhs/cqz9apnUxw2vY8hRqKw7UTAVCBdYNtXVubS2sjL8aYDmtfrKHDV
pNIKAaBaN8sU+2gIlgC+rbqfLDkpGtswPxJ+MRi7pi85pRW1+eStH0oRgJIgq/s/
8BkeNxJKz1mexo+LJZ48dtwihga8D1QwJTMUfs1ui0CTjgBWnGEpjot3NtLtcyHm
A8DvRsKwtjk2q5HXf2r3VHCDmW4N75DkU2aP7jT83I2NUQ3HDJbqfTWqp0+kP1uZ
8SV97RXBQ3FiPyjheG19AVyVFs+CdMQS8J1dXRn2B8z139DDruCD0OQnRLxcCODa
qaWMQPRaZBK0eKGvKkMae2/O8q0Exk1PYSQopNaA2gC5/BVZvmWDP1od8RFJEU+w
NnGGcKM26jEgaeX/AHOovQfgtHZBWPBtu3ZunaaHcX9o1mmVeQhz5WGoSnZ9lfIn
xCBU7p+hdzjx1ku1TeNNm+Q9ACxE2IxlLwBdYuE6g1FEMk/0EvOTCQsmOB3uUNxg
tkfzwl4x84yfzu/B8IwwaglsauGq3Bc7qGjeC8kgFAcsKcdsaqTDpyahB/7NhG6r
fb1pTYxaVRVUyHYHMTgkCEMbVU2PuBoeE119j3pIYhcbcwQpUOfFksvkQphkC9qZ
dSLeourpqWEJlvgrQp+k2bis78RgmZ0mnf42XigPAcclb1w1cQnsFoLS6QVpMck+
ljHkbUa8k/bLcRawFLuFgAvz3lNfiPNdNELpMU9bBCIO5Frs5ylGkXjN+yDirvPB
5eEKH7c3BKpWPV9pst7TZ5BKBDMcPDqqypWoV6shaqTyS84Mtur8+IU8ECq/gnQ2
Qn71Jr6a8jLOHXcV6KLD3SI6SkdyHeVj7Fxods5Ls3U5BwT1VrbGal7Zk2mCG+ea
SqkhcpJR+pILzad+hdiNJh0pc17dC3C18aG75Eh4R42r2hVTq1FenU20Z/zpLvV4
Cr8RU+ad9+r5nbZGQi3DEpY8tbma+GAsC0UWskva74ff1cIztSRED9erehlnxJfC
1JM+0uqubGcU6dOW0925kqptKuMo5j4hWlrVv9WuTBUI2AdcfukonC46uOhOsLlN
sBQRAvTQpG0bkyO0rSw1QZuZ5QFmeYoJA0U99H74QUbX4Pt4rRHHizN2D67dQWdG
ooTAq5DIj3g+xwJxzvdhXlzkUhT2QohC+seiozZU+rPYG7Y6ozjirdzgOOPBIXa4
YvGgUkzU63917x6uDSEPSvZaIrz+GMd1b5LaMnTVspQIWVyssMr9nPJM1iRr0ll1
pFQinidnBeCDJ95f4bAPtxFLBHf50dsO9MbZe6loyln1EmGHcYCQ8+c7OGznK2bS
YVo+rwLiAWGc7T6ZE1lMnb7LxrqRBGzvM1ln+cgJiTeN5wOx9vAFIRN4diFu3iK/
8qeGqsyFswM8r9M0P7ut/kZqr4tUbUpBV5nnsW36asGtzogz5EBC1ult1nv8mJrB
BiYJgVng0DImQaJUgbvsu3YL5CyC/t+IXqx3cgCropdAkyfIwa9uAMf6b7W+vTYf
5iE3XabN+9AtIUN2FAdj7W1T+PV9Mlrlh8w7OIwnKbh4vWPGfaCltx71nxhQwLms
Ywov1huFcQ4sZWCL6rWMcpAXHrimn4PaY5IdktEN41vycuRlg+6QGhZdYR8ondTr
GFKLWbC/f3old8G89beSRHl08GQXypRpxbWzBDN+dLNkCJ9AR7K7GGexmaELyKSQ
IvVNxaMY5pMyLNu6AjTcrtkejWZUX5s7ZDvl68ZoghaXIWZofV5Er4qBLcRDiffS
/8cAQjkfkxB5IH5l11Upy4DG4tWTjiy/Ux0ySXii7ghJqfL8MDh/eusjHoC51cwc
51yCO/y/ipNoK+N+iW2GT34ksJc7Re0aRkRaCQxTVsaACWEYzCNWfBXxQZBAsDA2
YZy3bFFL52VkbQe031divGSLnt86xR73SZY3QCuhl1I2JPIqc5Cj3KuM0pmprWyu
15fXj6wFzBRdaREcVEn6osP1ydwYkCld3N7A9P/H4UkEoSo6JiIMsq+wwmJ7Dk6h
OOt4rTfwlUmTauKq8Es3EhU85LY+61HaL+mziy1h6dFYa6fxArxnx4/Wokbhi8h3
MqMTCV4H52zHxa/nw4WyNt7DrZdhGWQ+SogHAn9kDKxCskkgSXhS7DgN1roAO8JH
OEty/Ktl67yoZBkucKKziwPOjA4Ot8fc1FA4RgK4w27EJ/WEFppbiIGlHyFkkZYt
H6c0H2gjk3r41ak53UEIa3iDe7aLPMQNE755TWaWWTDcZQn3GtVsU8vyH8O40RoV
aKX39qyuWj/WWt90afCkHBkyIxxA6KsGxDoKR51Nbtd9e3SMoTNXcPBDPLPYvFLe
oNXc3tSBCBtsxeUaeMIa1GJ65ft4kfh/xyEghcYvcUSuDh2G/JZJyM9oFxKx0+f/
Jcy2Z17yMCGGCmfqtY38kDR789L7+14zc4J8nNKjGneKVWjCUwcY2ynUChS+7aJk
n4eOirXByDn2FuGY8WD5a65Ho5PszgmupJbQvckCIQm+6hvDVofgZY+S4ZW98sn6
lFkhDou/6JCW47IZf8QG9+il7VsKhKhKGqMrsu3J0QQ25ZBRqnLvjHz8EsM3o8Ax
PrTiiXb+r9AffIR8RSuWf1FtllfG3HSk7tjhTIo658B06srbHR/xMEaz7XWubRox
D4J8wPDvKnXJ+L3YWsP4ooiEiXZgBC+CVwPKNUmBaanQpH+KiP3fSCL8FN+ogx1D
C2ba6iGFtTPMfoYYwUn38/wPO4FJXDFrWYonlwwqNhMVBNAwHsS+GqwygfDeb/Sm
Rwy9ASPj2fDzjKHg9Y6SFs4G+jYcFAupXiP9B20SUW33Z4GS3C14ye0pXHGCsnSx
s9IepJ7g75J6/6hzyAtfD/Ywe03UuJKXs8IlnV7UxKNPfJRhHSzRPvyoCroYPvWj
gJFXTWTCtPyKfofXpOZo8sPuPw/X0q15IlOiKQciMkG61mBSNZrNs0thOTgYkyDv
WhdTasvdMdFDZb5b+t7yMLbhQWYaGBYaoPK2BZKWg+dYoa/rsiYWmiOXTU5F7FwR
ZsOMrOTCQnbUjfOBVwJF2xbyMLFCQwXhFJ6YO3k3xBpwpLOeUPc6xu0hcueCqhu0
EYaqyJfQWMPfl1Cs4cIFY1rD1CXhI8/+G1xfbCdvFtgZALCS9Np1/WGi3xTTwWtX
DVAvAwYWAvyI7fhSbZB3Hk1DVWbRiILuKboATA7pXwyPIJJ45eOaCOtHOUCNvSGR
5VQc/uQd7sawc2nm5wBuhhDfjzPAiXu98RuGKq1bcV5Zog24YEro/6rtuTh1OgoE
4bpCTzu6WtjtQzkzWDEZ1nNbCFHQ+IHoeMYk5b9NKNF3ief/kK/vP0oNMep7TuPN
N88o/eNY2fhA+MkCdi1p7DsyRZfUlNZDulcEd5KrI5a42ganID9Leu73jAXpSr8M
sDfWZPnD5RFXz4Fh4vZmo1OTEMGU/xvVHrudNpwQsvNYka+NCd3kmoCY/dyRY1PQ
P6Rc9nUjRYWHsyI/u0Y6lTrhgMKI85G4/n0+3b64Uo18d9iM3ZwCE7xJfFm5Oa6F
itblicu5vusIGejlURKbhu/tJTZF1TPTiiCFxG8mlo5+zPZ55skhoYzMQU/oB4/f
kh3g+Tf3rg2sg7plXx55XiaEUggA5h+SeKxkyRacEhpRoPvSPV73WMjvNCtyEYnW
YXqee6OhPdEZ2pofjPwnZbDdS8GfntKqneShnik4e4E1jD1qKLgbWicsoG3hZkfA
UdaD+lgpyt0S9YknwmYP1pjlSXesbr7vfEP3RJv65LLsMgGHKo5ky5NrFoSeO6t3
hY74haVwjdt/r/jM6810CDSZ0FRx0qWTex5KzXjSVWpXwU9RQXgTDYgOlI6Sw1sO
hiwj5zPi/6xDFOCQivXnT6O34wZkkkdFzW2nMQIKNlj+52ozrX6IC2YTYdn4V6R+
RjfaUrewJmwxbCunJOtenxTL3tjPgLD6AXQLsOvGYa19dvoTu3WwXVb/My0AAxA7
RCNLJ34TgNlZt1j8hJDbhJIX866/4nogQASMEwvHAuhX6qPec3efzVLQNcsBtWFo
pkeKUkBNTE2nyr4YV8QBrPjLaURlpjtxfKFxiNnjrcBSSyqr84ib7afSxQxCFYzX
wV2xqyRyRJgtMD+8n5WogOwoiblP7SqrU1Tl64u1dkFgINy08PNeSdfWaHgUHKqU
IEzThmUW4z4DD+Hy4481qQQzuch9bK4ukkLfWP47Dd/4chsm+i/yK0B1GwQlomPR
/RggNpsJviT987ZzwiLiHCeOCk6W6UsDhVFqa0xg91qFJyEt3Oq+gHww2udEUchM
S52UlGTBCKldtSeTRq8IpU0UqSv5Fj+pQ9znkg1B2GpRYMwLZEeNSgZz1mq+uvPY
lsAwkasgFY39THl9yBfLXGjn8KUsfh2wQH80hKe3kQ/SJIe+1/rtL0ST2clIhxue
wYou+lMAgux6v6P9Gt6ElNikfr3xXPjQzZFE6RgywFHkB9j/wsVWw5Bp8ppaKuGg
gt2ynwI9QkBoolWnHpUPUbFJp30MJwgyha1u7gWnAvwx1/CncyCgz79PRqXwLU/7
RzYwUgqJhsmnCuvYUrp4JPnxXg5EReHFzaCbNxtjmgBe7mFAYk6Ugrx2gDZ+2GVa
l2sCPcXdMAoRjUV1tXiOiUs7SgsACJg06mxeAliITYMxvLm7S9+mR0BS4MYVdrUi
PfXZfTHZ7Lw3f/jkKsi0x68XuWj8+gi7HDncsZLygsCR8CrYAv3A9s7/DQcNjQ7S
dcDDn1IidiSXI1vNNi/rKxCCe5Slas1K8EcltQj482X6KY4CbKgMATZ9D96dHzG5
rAlYBa3DOkjozWKF9WAJ14GegZuzy4j4QMbWbFBBTOhHopP5xnwUrmcM+T4UlNsF
lssuqdP4b+Yg8oKj1G3sRBx29VBygkue7ZvLXGVDw23F5wWJ5kyo7J+nOgXuBMS2
4RYblv1FGX2zB4MKZ3yzHKLe14CuZB2esfsUImkp5rNpHYq38HCfWWCrloiVXyMn
f1NgwAx2SXldKRno8POK16+52N5lKqin3DeAOixHvGyS1CPaQ6fmjWa/S/zVtVFN
E82i+2vlBEMT5PEqCjIk7YJASMwbsaFgn4y3L+AlroiRvR05Me5CI9P+ox0NbDj3
LHx86qgmQV2aiODMu9zKt7ExxUCbl6+5512/A9XwLz9T+7oecTk6Db+qnL1n45zD
OHVusfYdgR0YQkrQLB5hhcSr9X5bd2IyDYlR1TA78DCWeI5U7/QW107AyE8diFzH
tPaZrRkHD1zkI5fTlVLBuS878xxXzOOJRzTYrBTVQWrSyvwuZBfkUht3XN0Raw+M
H1ddoD4XIcQbuYsywhFyciBuO0Ae3aqk+sR9uDdSwc4+7f17WvhABAsYz6NhArEm
ycQr/A5bpxqDRNvo+iY5954oB5uhlPkOkMyPZdEbOySCGylC2qTad7aRcZ6Znlx4
34jD8Jl9JzYLptG16d583UCF/wKg+GEAV2DR9cp8XQ43vLLms6R8QXipikD/hrjK
8bn+aJMwcPtdM01PUxVAv9YAEIn8E03o4a/OaASli6CIybzEIBRuyNGrNm8AUFq0
lCtOT1fNa16AXmUdNZCyptNeYMtqeSZ5t2uV5G5vBJT96ydMdtg/+OsH0gHf19H4
5T4B1iFF+9zSXfCa/WKlkyELpUR/sTDJV1wK4HCo5hewTg3B8UEmcJbu/gtH4gat
JLN5cANHdzXP5HYm+nJ0C2eKkfodcwy1VWHkaQdxMQwlVOlI7V9Q5x/DyN6+K/5+
60ACXvwyXVcggFetY1pTyPwstlw+y4n+Np1sQLXkqOlT/JxERlOBhzCAfXgRGqWW
uXwmv0yQos/jd4sApeZLBQzyQoC7TQXrhBfnshccjiBzlR5XVx6/LMTEQrQySSYX
sQOvaThhew/1szc0QW2foqWdHhPPb/1gUph6H9ySGiH9pTvoDgqFCfjcwiuC8Mq9
DkywTZU6Hz7IqN1NwqU2RMv4Uz+PuU7nI0S8SRJcwfSFEwByes+73FcwAwWKe0TO
SP2uvM/ILyvoMkTGJyqwDzUYC5aG2nXYGAQ0v0qJ7+ewLZ31zLNyFG40LHIqQQTR
I03kwIAZGu2Pfwq4/WNenXmO9LhRRuPQBiqCBCkUfED2hdIcILp9j/bB/Lti90Lq
pJkdpMp0U/NB6OCxunjSmyc5iuXBscJlUtQUUIvjCdme5TxerKLBCwqc+n7UpYps
c1uYrk+K0+RAc1DtlAh95mH1lr4FZv6b392NBMFIVHYpoTvNZk+UPxrJ5kC+1J+0
lfUiTnBni6trhY1QxWACoI9rhHqGJTv3AKI7XadDwahL9Hi1XDfQry96QwiCht1t
+gfgD9k7j4Z1dKpPUxoNo6JNWVktcw4ItjIyOlXMSxP0dmO8nDfbO0JpK7Y+MsLZ
hV+B/sdbyDPECrWGS7e1tEpznN1xGflcly8EXoTGbPLyP8ViWWISh/tMLMqZ+VPB
N1X9AJIirNxdkBzwEnFtwNfD9KFxx2ck6X0ENYdFyeakMagf4XEPC89j9i/cQIPj
DRHiMkcRSbmNzbSDWZnle0rQQtaCClbZvIou142Kxwsuvo3sjpz+fYne8XW4lrGP
RmnAIcv9JaKA3gWkaT1cD/uFe6KbqHgQroBj51URW9UJDiLLJEaeeydl2XLFBnq9
KVpiqwid/6pjb98zvdC2gKrcRixvZB6pTbXj1zyDC3y5vsEqk1n7zzO9mhkgaO2j
IiAGHlFEkOB1+Zk3imyvfnfmrDC1iqrE/PIx/xJn3wTZ+f+TPEihwmmIekSKF3XH
wCMwX9mjqBlzWyBgPERDFKDdh6subv6ui6QXP88yjE7wYO5dRWGkVJaStxDQgfJv
hZmPzZHVmU3kbY0nU3Lv2bkJnw+JEOyXBzHUwF6youSOyVuPQHykt/IfDMsWYBsM
YxjHM+75BmEFSBMW1UagljG3IcSZxibhPkfc2jY391pqzAreoi2+A+KLQAt8UOPH
KvEYMyMRqjJVc8TIqWbrmfsoc1HSpqac2X4GQvrNMqXi3dCiTxUUmqPH+rQBTHmC
VzksCIF0n8iWvDkhBIus815qQtaMUm5sn05mPi3P402XezHTgzXo/7lBw8/kiSjC
h4uoA1qVGnPWoAssArJtFd7JZ/N+C0OuTEu0PwBv5/qwYMulltIfuqIhF+C+oyno
0zOL6oLaSsJ5ohuxKEDY6CBdZpImNz+D9c0zFzPe8YPDNW4uTfPiyGQqlPJaPMIW
K9r9JkFA6swf4QlifRA5N96gH4vdG1qaxN2YrNslG/8TBHTuCsxNsNCuJcV+W0Bi
b89XP3ZOcd/4STIt1ksTe1abm4yA3SnHGeinnGYCZUu8grVUS+UH4D9fbAZTSCWE
7mAhW+CWhDIHuMZnmAQKLMgicR/yxTk0C5X1KzX/+oDDQCHapw73EtNnkiE1cz6u
KMQNRzoK7MT2obUdfsE72HiOVVEg3DfeyATBuhyJn/AHqbmbBoFViQnrPPJ7QaPh
nY5pXEcp73GMHadwX1fnWb3VFL5LIv6pmPxWOEB9GYHRj0hlSfCdfnEyocoS4SU1
9AVlk7BrRExiWlv0sA1ET1XE+FUGxWKIBjErzFVedaOSfJzjQLYGYR4WDKNwe0Qb
3vGObZvifhxcbisBJVKkpRCzCfkGRs0hYAIft/6JVvPT/cwDgloyQd21/sIlbVUE
iAeLS262PWFgBMZq8pQTnPNaLOxXkQsFKw90eD6bdXNFk4p+qL9RaTKgFk/e6whJ
40lojVz62pMZe17RKDU0b1TFYyAjsS17bE94sAirGs/9znWy+7Fto1MJZSeVaqH0
JfUz4r7m5WP10t5+1Maoqc8bGOj4LOnCbaEzxmA90URhoV1YIHWSUhoDT4Vpscty
2o+bJzPtku0JYk4ASpbWWzdBUdDWrWajWeaSbUZBpCvt4ryfV9J0MjaR63x7W+LO
KyxUHWAL5tYQOblHQ/Ulr6TpTOSF3571EgnX+Mwsc4HQvheYY+4crSocLQ4O6Rc5
bcqo4KLIs0cbtr9F9fV6QpV7CvqAJSLgBtEUuLah7wGPKcII5e5pJKiaAptxx0Ng
7Vo66n8jc1UX5Sx+TEjYZYrJVU4r+hSwABYGFWxiTE4ET4sZjdyobDx8n5jaJjXy
ABmVZA1hZXEPMwtmQkoNHgoiUPzhOC0/RyUYkEXTpdQaqf+KIJFqDSR/Uq9WN8Ko
NrpPo5sn0axTqLRaOPw9T3lWfOZWLYc4TXPw9xJmOBuYz65WCo4esU5+ZtD206vI
lsrj+iNy67bSwR2y00XVrP/G3SpzrCInT6XAzr8YfzVvc0u9z/WZ9GPA+2Zo/4Cy
imvRJVaabRsNUdjEssqVTWU2rZkf8bl3yVkdxBM/pZgJdWGdUy/uUCL5PCfOylnf
G3dYW4DFDa0aR3WWvYDdyT8JxOyfHXoAaub3bj25xEO8kvMQxLUxk0TusCakXYKy
e8cgZCQPaH+9kazFt4iC+ywNdUKcpzMjUJukqVOZIFYh1hiSfF6BxSuK1040vAZb
Qm+OeiVFl9KQLu9rb9MS6pw2+qstvjHvkcnrWkCXREmaJGEqM9cfwJbyq58zP1MK
8QWT9nDOKSaeiSgbAXBMi5/9C254gMDbBZVLoMlprWVEKvF6S99D6tBi9fjVmwKn
++gY7A8wXr2Vh6rnuLKnQi65vsUi9De4S1kEI55llENCW82xY7x9nV1K7mx4Z2N7
b+CaHok7HenOHRAQGCfOCMVSkVFBFtVP5Z8yVD1eFwRZGbANvjoNj9TtjwkT0oVs
QvvRIL2IZfEZEhQIBXETB1fP+S4rFhzLFMqVayNx5ValcbMtag9YFCWbUXboBz4I
+URLvrCSX1O/8S1NHEdfNl+gTJic5NJSFipLLNVS+yFYeGY/uBoPC3bseRxj7bOU
MNbLososeidFPUNtw6ZiJwdlSsS/rklLkZj21T5W7pBEQGFC9+gzFTALonNIbRv9
p+YKl9/Uagvz0jFJmAuIsLhQ38QQRy+1olFJsR557Ce4EvDMXLlMsBzURowt14W0
YLsbQT8iThN20dFxWv9/XRTWBVJCj7IJ+yh+woUNQ3C4SgwAP4XJMhGYvpGeP4YC
g0k2nw+xWZYOk3sfwoxPm/MrjXgYtT5mhph6BxFBfTRkVuqk1jpZlWFq4l8OEOo1
NzNO1nqkQeF/9ApjM6tqZo+ZuI1/etMrLO8nzsYigkGW4khwD/aVffSZZrcboSwz
5Wk12MhwF/KHMomQBGoacRcf0gSZdUTHD+7+GVXZ8FPNdh9Wot6MSIMVj/2/THuZ
1mbZW60n9GIbuadeNqQWcCYjZBNXUXosVyn9Q21d/koAZHptdpsyFOnjNuKUEY3w
mFDti3ZDMSCHArJBnLjvcKzaDZuPpxNwMER9K1pkFM8gtvjDE1U/I3KAlplmQ1oO
b4oUHjAfyjhnraKcYBvq6scPoTHTgdbnCuhvJP1ldwUp6qmRmFjhIM/mJZUIrTTh
a+nxR0hSYwEhfs1PD+nW6eZXQMvME7ZWONGahX6zPbCmNMVpBiviRBZ4lY95S/6R
pfm9dInk6VR0hhtwnx+HfazQZQPlCA2dvZvvHs21nJ7GSBswQTHbSsxvNbi3Lo1Z
ZJABVrZeJ7hoO6T/eLGoAd386KfQh9EQhV994am4kS6ZMjsnfdQg9VKW7TuP9Y+p
9glJ7Ga7DO+vm0KKpKXXAZOpTWpT08ImQDQQJ+etEL9JC1q3fXvGu5TyqjJJ4hQC
czoUIcFTq49BYBPYws4e2VyXdosS0svnGaLMWiTvUm6sik+++fiZoUbxkK+WEABm
3GcTcYP1R/DPXXgEPsfmBSGA/kxIWVmyOHDwJNIwfqC8nfVYQib1/VY/KYl56IGP
RTmm1jDnEDWxR4cJeYzMgzCzk0LyQqK6RTECOufke4shrsC92avVui4aXvZjbZZT
sg1e7O2wo2IZzIsKSEvjyWBJunGmWXMxVeb8SC8VuQhJyiZ70w2DYLZBs0SuU8Km
v+tK+A8GYNWJj07K0Kg3Yci3t5PX4iN7R/Te0aby2egmkIGheLhh5jczGfBnt1hK
hewix0Seq5exK3iTlfitIH5C15vRzsaDWjBxgUao1hAgFtg+mss/Nw00gTWSpogp
/dnbn6ARSHETphLi223qgm2PHzhW468QNtJtsaaTTfdPs0FSPGbnuG/L2DjGPjJ0
tMmVR8+2Rj3TXhOPLNglftbvxJTTuQxvZU6f1uekfAdn7VQX76QYxTRhdAtDWHIl
zxOx1+zsCn0ndELgbefEcqNFqNxgUmqteB2zjb4+psgFuTwg/kQFibxdkbSYpllq
t9gUN8FO4a1EdMZquBG9HXlttdaioINA+GVDEOXlaYPyLj4u/ACU0R8aGY7zAifL
3UR0tYbb02krxETM3gru+ybJmAtdiw/wdaNU71gWgPkYlZnM1vixMC63JqoNLJCu
uaR1njATjMTWohpJPHim4Ulw0o7eArPN18jh+ZbQCX1kqmxZIufU9h6a5gsxF3bd
qqidLWaIKgCJ65HrUfLdRTb6Uj4AgVQGKKfKTGtrXoXKninCZCVmfzh/bK4DxBc8
zZMCGd3FFi7hHzPgpK4TVU0TNgl+VEw6BhS9qY5F98uY5Ix96fh5ZxB1XT6k1wi7
Ufx75SOWnNH4kFvc+hydAzfMkra9DG2U0PCB3HGpNRONDbYNubWY3IfGT//Y76k1
6p+z6YTQguMzoJc+hm5rRGVCk3RsPRny80j4KNe4iMpEVdY9PLUqDew9dKPM1etx
AVZ6gkd9s9RNhOyHzhllXUZFGuXl2qtUDV+tCE8H7TQfgYBeJenDj/v40RB1kug5
wBRhUvCQrdDVG+I8NSmM4oPB5kBGdsNZbL5nFfuLFoxnNyEPaoPnO8TKoOq80fl7
w/Aymq7fFqCfVeZn+B8lt7rtDWY/GcXd+UX0C+tHPDuMK+TA6dBLnyrc/vbfiP6F
WYlPhmWJHLtNWOwiTDBOORinjzj7uPcfLTM/mtfGrWfTjakaUpgBYO3JLnxKyUXG
Sy/4OxIdOh7zI6LY+z8pe6eEQWdetsHLHOtjaDRyUrXSktpc8WqMsbXuWZEk1D0O
ZhCg3T/Z5hVlAmZQhR7DMFXBneqBPbPE2TC+ufA5o4ULcw1xr1TN3FVLaTvi41A6
2uxRezoenH7vH0ptm34M8Xc2Pvzul3TGo4QBAJBn5Z10JGIre2vNk5ZpLWdPP1iM
yQxqIIrwN6NZO+sbVzIteUlfo4uBx7gTIAsueojjLfvXxpHbV/1f9F7FmRbdTf/Y
A2vrCCod8ss3m+UW1e2z66cpMzh08CKxIJ8nI7f6nYpakOa3yjpgz6lvtz3M0I90
LZcr/O8TWAZCJBhzEydLAchGdZ+h2MTUn//Z7LVSJvRLnoKN83hxsR1vGKitR9e3
I8szjmrdlpAOl66U9xrIWcag7D8M16Buv2y6sgMtl0HHNic89V/rzgl/qXrYB4sb
HL3w12/wDoeIsOflYxYeANSOlq+LCX3vZRRD9EMz3EJ4bJm4x6vvYmRdiEvpHUpF
gxumWgAbHZmTur7PNj0utNDlF105gd6cJu6XIDxedkgs0SeaAMFcCmJABbwl8xyQ
LXg2t4CRBI29sZurTPqrdYVY07fBQNebBnQUS65QMBG2iAJSf3NgzFKt952IcZwZ
dfuUqstMkH0zr19vwassQRXKo7jgNp8RBe5Li2sSw52LkyUpdLr2HE1jt5sL9mW0
K3fU9NaoCSV+1MQQS1Wjbw8RWW8lcOY28LCMTGCJrjtF8VhNV2Vao3GgFtdMc9Ua
qCEKHnZpz+JcQXdLkDxG0gGKiEhHOHxfALMTcObCvHSDsXCqviQ1CBOUWb9NNmau
jL4WPIQNXU627sSX2IE0jHeCcB8ciuBWrTjB3j2tWrZDfSPHlmsifv6wMbEJdspM
cQD01alZqNeRto8IlgcWmBwX0H7+0fVWr8IJZKRyCG0rQ2aIoeDBrcjfNowmVozE
b/AvlGsSE+VdYknYtRC/Q8eUZMKb78SvMK4iXBH4NcX4N4HcBB1lyCDTeEEfFqzq
BVgsaXKZTEq+DFy/EkkVhZ99cLIXQs6/HdoHQQuTALy48ryI4/3V2zvRyBkxXM+W
0XGYzHWFLbqjHMtLIkb26+hZ/Gr60ZBeyM+VRvsjgTN9eSBln/EYFWIg4yN+2g8I
NR90eU92UDNMHmv453RmKoj+4HxgxtGpjoQOnDOva3eC+WTkb5hypM1f72na/gbb
QEwz5J2T5ecu1FzzJ20RclGGENZPXdrMSbrs4m7jnFHrH5zqu3BBk8T831ec1oYg
YxahKhInjJb5oqXUCUtVFTfJbrr00DeYDU1w32H1qCFE92pUa05S0R/rvioXqNJS
sL7YJDoUqOEjpE2CBIcZ/EE7TGgTWMuw1BXz16rwUga6dt4FzjJD54CKYI/XWMYP
FkwedpwMX92rjk9L1cvsCZeBcFMAR8vF4ZP8rWe1Fy+FB7wB7WjEmQe3Zj3250Bg
1n6WSyCFkX85+D/XTRuyNFObOYaEvOpVledqN8VssLE1kni9TlmIAxqzdYk4DVnh
cXZ27CL931pzJHErmCxidLvrbpx0E1Pmv8FglbQXqFG91uB/KoxZxUn2SiPPYfnT
DCpUlJPga0BCXKnqwQhgJOZbV2WSYnEdAn/+OnRvup72YeefnBACsy6CDNRayxYM
cNlbm3YKSPlPK0FepiMUKELis7AdX7tkKZ+5OE47M3iITgAhrQC9tMDy7A7LiEeS
Z4FOhGVXU+ACer8Q6aLcGr/4eYrD0JBUAYxdmE1jvF+Zp6IUpiDNvaYcq4PqZiG1
38lN+qozdaEHnAuhndcUbmbli+RtRdHf/mygshasGUK00b7mezuCb0xWOl+SGERi
69aGo8FMQSOfbkKIWLwf23/MExvS5iHnZmKWwOe43QyEIkL9UYuvI/oYC+91xyDZ
3lfGSfIag4fq9QwIWwFatrpjE10fhoG3d9jW1ejU4xSENEmKJl84kT57V+J3MqyZ
YH+s8gD0UP6Uqx+GKeJw5SuY0heKrBTNJakKq29FCJACxlt/pBLfEsCaVJZ4wmOZ
hXSuwV/zQWP6eQh3LQyBr9YkEyHZv+QptaLW84pedGSzo/IZahD72VFUAsje24Tv
JcoC7yg9Xnxx4gxrMCYIOr6uT76QWMC0ul2zytaEbJ6dymCc/Pl4Hui+fpqz6io7
cUNwYjUOrGBT+7kr5a0s0A31fRGuKBUWogRkyFdbC/mATHnVcz7cKZwcOuT6vP/F
6TR0qWKlFL4G5e6iN+BGQebdCC4wW2RD9DslbnI4JHNDEx3c3Zt8iEh0vEqQeUa9
RpB7gEZXuXZxM/MS0qB2q4s1Vz54wO+jWpUkU0sX/4L6toKa3w+8VYlLkQ6cnjps
vwJyhrULiX6d9JF1hgmV5vn3Rn+DSCyJe5fRsz832EkAxv+/9gCUJSHrt0+yOJEc
Iwl18GCp3fUK6rSXwGZfy2upItiafSN675t8l846IhT87diyKqQ4WP0O83X+mdLH
AfSyZdc/temMQQ4a718jIsCbdb/YvK4FwebFkN35mA7lK768dqHJSYVIZmREsY/z
3oLn6BG4AYJ3+5Fy4jpve/yYA/4n7qnipD/iU3Dkow9GbyITkH6uvza9pQKkhP7o
fKDiGpZOV3F785a7UE+X2KPyNkaOGZRUqdqknOYeUt8kgkgbyDUoxR92lH1Y1zde
lh5ozf+zAKiqJ5Y24T8bK18Ms94AdCMV6ErljoOOIxgEvQYF070wNJkR6G1HoMcN
ianJDbwWN7EiqdcHfQ58ENQBnQIqgu+nIv3PG6mWWPhxgpuIQWBrLB9q9sJcJSL1
hswjD+BIYb+ywHCb6TY/5WbRH8HPeH+DniabM4T1/Q0lAX9QxvlZwVZJDpB9kDa8
t6dcUy0Kxqmw/iIArMLMsGbh6XATMW9GPkOPskRme2qwXFRfLw9j8VUvK+uDKoL/
IfPL61KAkdB/R6zBa7Jq4NJExA3Aol4K8gqD51pDMv8+cxLXdXYTT/inS902SRfX
sdNo7K7Z/g8xRKsvkbzL3UUlowccooKlZLUSZcKj/qbtF0Q+RDXkehcBpzfMeL8S
T4X5Ka9jHBGcQATlbOLGYJ52UlimHRbBy4kidcMn70Rz5mgGn7gSddI+dcdGQwag
8iDQ1KfMVxhkS/p6M08XgkSuvpUT0L8aSO6IiBl1tqDWklKeXXogq0/DJraGw/lj
fafpT96lLwW0Z/PQOtguS797k5pSx2OKPbhDDwimHDlTfjSg3lbHchoP1a8UM2VM
UR6glWmpngnlW6jNadxCzYVzjVw4+N2V65ehAEcnQneW/tBWC6ZWcT5QOkq7UDtK
NfTFr+LRiRqVTXY59CuIr3MbPpkQwSRp+t163QzjbHrrD5YB+c1rUfWPCiUbmLZL
bxRqh6rvUTCaKfPL3bTp6oiaMB+l14DM4gXlkE5BpqQjqzOnjOQqDJpc3+jMbNFX
O3Oa5m7y9pYYptat4IUjOzjUMsLL7HOD6kbU0u5tfZ3WTCELCWZRijNz6CcPTS4+
TRMFSmAExb3NHb+vpPUlG13pNdKjXLxPSjB79+VdFTy5uhqqXNOZ7vgTKS+4W06p
voR4GauzqHdLi+0jjnectplhj67h1C5McSOxgUkgN8IzHeTJyAdDUSvspgaAtNVj
wj7hyfZNQEgm6WtMhFdJ4X60K74cBUOMjBF5DdHdonjbm5Uy/rK+xdPAnHDEzzSW
3/JnkDsR5tXWCfEydNZygxyAwhr1oDC8yRMFCkyWaH7y6vG1fZS0+1VJGI2/k7D7
WdueACV0N4A79toqkDdR9trlQZ5HRFqv3l0/P6WF2okzN7QuYfj3zMGIHioBqVcV
2JgXNLxQuBEoFy8M0Mw5ADu4c7HJAKSH4+IpFvv45FdWUEOuFMAei2PTMo3W7SFg
7IYqCmZw2FbhN6cUw80WUAE4UYrqH9LgaGodRBVU3DsAywYveySboZzpaA0YrTue
5GahTY1LE6X1JkQ6dbEj17s6dfX01onITaO4DmadJZEAhQ8u2BJmkDlECCcwtk4a
fGm/UmSyoM11CMenyfteH0Cd5YRKrZwrjwWBkL5+Bkf4UgzHtZvA0kem+AR1Nu5g
7unPIAb3t21IT5O12cbNqsFHUpkSXtK5VhsMENKG9DeZTz1YRW2n+D4AhuHC6uid
DuXOHE7TwTocd6jVnH2XrFA1ug4wa8QK5Mj4vu5d3Xbq0PRZMqyVmZrf0HD1KHuV
OaBf4Ko+d345KIKtaqI66yapy9XOOJy2elMIEr/cXL+xFBYekRkLjxmScjGvmCsE
pykgtEEheYy3WonTeD11kGnf5IfiB/kDycsSy/nEVwFkH6viDo9Cnsq+tLsCYg01
VnZBe/k43nkXrlKQQuVihV0ZulKCrdbMX1yViVk5wcybFc21A/gAIyQrrCsP1DEZ
OATogFrfHINkUTiqPkzcULZgYs5JniL094mgTW0Q+0wcGHTA4tjcoCh3TpVAI1OX
VyliBonAiix41ZacPuUvn5HBqLaRLQFrmmDfq28J+os0HUEaPcLHQyvkrz3+Y85G
EEf3r1pIwH020OOcG+HtnO9r2tIwhMdOC1iPB954u1izcAauOVECq2zOC02jJlZI
J21j53lqxMTe6uOsLsm5uUkizUYjeAH07QKG1vNrtSpNnXXTUEoN7y8zt0Y18wRt
6lNzjMQh7wxBqJXw+LB3eZEPixMMzbrXanxdKE6mRffrXq1PKyiFl6B86mfTQDEy
FeaaHEX38NNLreyllItAGO0Rv9vuMtZQSye3scN0Bqn3qqFmOog3Lc+82fXWl1+M
s5gYB6ubB+jzW8noX7t1o9P0mKm+Qd/iHmDFhah8Jq6Ml9uSy3DApuq9yQEj8FkH
6o8+FwHCfrEnJ86oyNkJvaNSSRPsT23x6ZOH1rvenORoX2S3QmzZc8WR1jBUC4wQ
XhEPlOOOotVrMXB3oPIsowxq5YS8s5MCh1/iW4We4GKXY0qHaEbpM+bbXbsPMPrZ
8edLN0mRylXezplvfKQgF3XxAb6CqZrS5XpY4tcUe102GRrHNyWtsaFhS6jwNL4j
FCPCLL+VDK3ruQyKSbw0yd3huzXeLiIcQV02ecmUbWuFXCNfgh/ZMgvDSEhvHv5N
BFRNt/VLwfNW7p+JbrcSM5S/VfLesiPEGEYi69D5qKsAInS1+XUD5Jqigcoi7Zrj
HL3W2Iws5nmuYtnVKODZtfHnCGy34j08vGsdRady6VzHe6EabJXb5AVd5pjWD1lR
Ej+UK+uc7/VB+fmzZD/hLHquwISoaJN+pWFWvWWupunEId2GNGLvZwbskJjuITTn
dp9eKhrgTuNab+XjTlQclHkV+lD5AVDIln12xAlNFyQ4JZyPars8cAWXGm58KYHn
LDdkftPjJftYjSvox6RDeINNBzPrUsaD1qjqkOMDz9JFqmi+WUOir2H2kzbyNWtB
S6XLOMhtbmirZe9R6XmEUlCguxnHuqIChrRsvBcuMQRL6OxzeQY6cWDMEYMGmRmM
LO2/tEz7GQYu4cZ8uapt7yzPCE+89oskXd7KiZctHR1UwLxXIbmxWFb2YFYUUz65
XDRcUacezQrAfGeQJDyPG7iHfoZJAtfmiFve8Akn7+mWo8096P7UJDYRl88F1x9x
f/jdcUnc9wiX2OQLJWWQU/s9BGfmPSrIFMXnHA0j03xRacKpdiEG98V9QwzFW4n0
dqZDLsO5wFSvmW5lFq6VdlR1U7ncwkAfESkje00XX9Znv6AMTwMRCrvaQojAz9qx
HGdGrevFvGvrQQtW4LSTGAVBW9aYzXwnsNNT9x38CuDqLacmBQ1A+T0pd0aHRUWu
kMesr6UIAt1d3FjK/jjN5jJFll4ipEZ34oMhCWBAp1mHFjPSb1440fg/E9ndndn4
r2zwaSU1NQzkabQzHPVhMsQSbsawuzxHD8qlHwzaeYgAuIRZoKvsNLR+S/a4036l
efSfBANF2EH7HpECMvgupKntiBSpxJyMmfkL0ALv89Ofn101RmSSF4/U13w3xYuz
Mj6ITj30ZeKCadrOdt5mRYhr8mMR1gm8w9jTrVkPFpO2zEU/aMQYu67NSDDnBZzz
hFAAB1Yut78E2AEi+a2VhEYBs78mLuK+lIIJ4i3zT+RzcZSlMFyVH2qoX4Ymj3Ha
tsBigMfxr7+JJ9PzXspQQ+/Ll4eg5mGVB+da3MQZaiKa4la6I6lKDzbznZD5AlJo
9xhtcP48gog2tBgjzK9dRlq5s3fQi3jVW6NXy9CojKlgUgJJsrJ4nGPjFnlYy7lJ
1k0KkehwC/GzzJi6fhlDGIrM6wu/Cnsf/z/keYm1f4Dp671xCbsvHs/swSArWZqG
PNG/BCJxXoxm97LoyglCPEwrwwO/UtOxjAg5DHLaqrktW32SZP2Q5neXd4pqZvtd
rlfwYzth6fHmdjPE0mwBj6isqP8Pnd+BfIyIMejGQtKsAYE1WFiyoV72gtoLVpPG
djhFCSCJJf7wTfBYPfq5KsSdnOUrbv2WNKdAs9miUz9TxGT7RRHxfHCj5zQnBrSC
8v2EjSjgEDpabJmhjO5IggNxaVXbQTHK3NpINizlNu1WNVECI8JH+XlH+umPJh9g
7Poq/V56UxIBnBMqbDO+rUlCrlnw7rprbRgTg2rk3JqYiNsIVsrtnHBgsVDExo8w
rbj6duilWlZChnyrNe6iXKbrbOM3nyUpqaE/VNJGqtqP1AXYQfidDr4xeTfvPe8t
5C6wN0tBQNgEAiMsXBlXlX35grzRuYfVy2qq9qFVGBwFxn//e5dOvKvxeJTGmPTw
EcyXf2nN/nkNytwTr3Eo/MpD7MO7f6i6hLh4oXPGfYBEh39WF786CLlEalB9Xp3H
36TEne/pdBodrYx66fW2tft5sgG0A89p+6uygMU2qvM4haVTI0Oqkj+k37vu6ZQY
DJYEd53+KorxiUWNrUGDyOVe+IuxDRW7EcYjD80mdjlQEM7FzvfUl/lzw+VoosHF
DlMpABUxJFbQ3aefjI8yc5QS9uDHUA7+Rz9BsUQDHi7zmvHug1N9iYY2IVGpZDNG
PHN0toOcME/t30XAHulDwha1qzzfFJg2qmbnLWGIg+ef2BOQnK6N4OVEgxiTZSeG
vCjqOzxv2GeVxzQeRFYi6N6/B+iP/XiQwivVCkKx+bCgNg9IaBKFO05dUV3y1kNR
W9hK2vASHfaZj3F6/13bSfARlQ1VoT/9xyl1FBPccq4oczdkGk8SesTYrU1ufq0j
lmgKBm8zrBBroqq1BXKa3h/RVWhboBkbLHeWEF0P5lvXoKvzNruDBXoCxZ1taGbZ
Nde/jJ3N4bNX1iS9ketiPuKVIFlmA645ejE0x9XHNQrJZlgl6jsjE/jsM4Hd6LGq
IaCT6f9aB0gX92+DyRSTjgcexyXbfsGNYttbPPGMZVSh1cL3yuIpjn0OZ9JYNc22
05Utd3lf1MgO/bWu1gs71O68YMEBs1lUIsa1mXLeI0BxgamLXbacp2WzxOLG8mjy
NNbIObN713leDNBRTwCW1mj8HX+Mf0du3wpItNsvbGYlz1u9xsOE3bfnXrtUDL8f
fw6GVp5K4I+1xmCwCfQRiMQS+G871S0emdrAQ/C5J4hErU6E5IoAwaQLKr6LK6+E
QVzMMkKGQwafOU7tUjcagFYP8J7ULQyCw12J4I6iQmFBTWZreQZvccJphqGtPAfr
OTD4f/PMiV3mJcfuIwojXDAblZKl/874buHNPRT34/AFfrwKNhoTEFqrMxiYVAZx
p3fXQgNdo7Awngmd9wSR2epQ8elIiIjBBQFV9vQFM4FebFQD8LQdJSZueQCiYkiP
pF8wdpwECN42UMxgjQmC9fQyoDeLsqLWtH6xsq1AFABF/sPXRPFIlW9Dk5CqP74N
V0MzRphFYWYbZ8pql9tT5lAH5UerqEWQhULy7pdx+2otndmKXi5Pa+qqqe1R6//S
COV2DjBjv5C3IYwKEmoDckOSrGxLvzU73CbmSlcVRta9OEh+USb8vUPduGs7KQjZ
uwjsSxCkONvrCpOfbWzEHZtHWfwqQUD55DirEklih+M8yiOP8uH+jq2/iduvR/1B
coANKP/wpgU1HQocI/oYu7S5Ewh5bFi2n1W7dkdiQTDyHNP75eKwzqWe0KceGFNY
YpaDMr19298ECv4f0sJZ8IpuZiGiQSCNNAafrhn2zkd3PzXFZWXTZqAkRXtEgCis
gYNMQhTHR1uokjf5hUP/YXGantgSK/uFnZRK+BUXSn9JbBLrHs6LMyu/S01VOX1J
QhOCL+e/BEItyF5QhPcrqpBFE1iSGpZwS6+2mmJvsheuj9Lk9UwtTCSCHwzVlpmJ
RrOaV3n4N+4e1WpfzuoNwYnuxWcvoWxg8imVYgFW2QmMmPrRYG7v2+6X9GTbJ+We
CcFa5ncT1qg7aIK2YD7nTlBufwTIAFnI26X+8bxd0bVJtVICSQkjsu5SAy/IUJ8M
7coMDHOspHbQc/TVhUPMkzpCWQtJI/bI45rZYFdcpWEjqEjZEFZsKJFILlswkPqS
H+sxZ45Excapm1T5QXnQlDlYpwKMCiP5Ti0dfGX8/M/46RT9kt1aUpeDxIi+9C+v
KKOKWtvEpbAZSzyEaPAtMekO971K6aqMYZmvfPPgkaFmxUHAVBZ30u1i1mpNqu54
PSmg6myZp+4sTaNWvD48Cy6BQ0nO35kS7iV5ogSfccAYkSaMErunLTiACVpG/hnV
cWNA+f4WTh3UWtA9uPdU1eGGXxMKUwf3YnPIo8XR0DxK1+UrRhYmzjHVzzvjd8Qu
byfjDHuD/pPkeQkAoc/BWe2lQEm2zZF9OBCJbLAqzEpjUAv/CSsc3pdRD0IaVUpu
erMCSKLrKhI+sndq3InEstrHXaaaFPGCuQKYaLi4Bg9XCfdJa3hFQGLHBmNTDUPz
86BztiPVM/z/TIwM9gopHeknlmPlnQYQa9R1EkuM+pWMXIsLrWPMMS3RXrufraPC
CqgqjHeuUyZWODyJ4oay9GkGzuUfDdDSJL6gDJoR39bZrSY+8wnBmtc77O8lfMtK
AZ4eoB1MR1z9RogbdDjSL3xP1S02l4p23447i11i1D3XKXK/zSiElQeNLmb+pGlr
rC1MslewLmNZu9Ll/vEWJb+wpxIwh0M9yaBVQQyVEC9CSeL4FCWO31Bh3w6uYMTD
xIg88NbKpermXJqy+OMq7JL+N+gHQcK3tEZwlj0skk95/AKAU9aL7rAJoPHKQ1NQ
FHqvNDUMyGOaeQf8s+kllOtd7fPjEb7tDOVWrSCpDTgNvN0q/zGaCEgWA6ZwJWPI
pRsajCCBLWV8CN/GMgbY/caqjoSL0FO4rSfH8LGXYEo2CfX2eJb9vy7FF6zlgMvs
YtnyDrR5c9s9CiveC9eS0LC9CNZf/Fsv0/hqNLU2+X4ZcoivSkYb5NDWnFJ19bCg
N0O9lYPXtuJW0sV/LCP7+R0b2KFpC9NOwr8ONdQmLk0I+IeXhhvxiHfi1qK83vzm
6RYwa52ms6sTzo60lH4M+u0k5F/LNepDNeSwQF9kPXWlJ/ZNZpFl9wR4Tv56pwI0
182JvZkBf52L2FH33l8iqDlo0R6rZP2wdzvHuY8tCC4hYDVOLbK0NjdWTZbpapJk
GMrnN3gqToFdaVngalI8I4BEYB2976TRdw4ziKDDtaRD6yvA4CHjMhzxrF+a1P9O
uAodlkAuJJSt8ong1gciivLMtDM+cdHJuR8nBs98ljVaSzsVYv3mwY33ibgvzhAb
tQTXahmn/GYjnD8sf+JPEUC3q8MMxy1odPypAbfgDQM3nRwNSgHArCs3LkHhOAAk
BD0b0HrtrxWoKHavl7JavOEWKjdqpiWcSRqxSJVtXlcISowR5uq/k4vpSmbbU9iU
0t3oL+/Gk/mcv6zmuJT1/mmryAcmkYuUNXoNWMZ/Pg6XhRpJuQSrcI383DdN/crl
RvbK0UfLJHi5/id7uqJX25+eeszVrlNQIJIFxM4MQQtrxcuNBCnPZAyfmd2kS8JA
aRjHdQdPCaY8KCTKiPGPsERCNJTeDHroBPnEZO45u6qbscYqGy7J9RD4EnWple6s
OemKZWxnHrIjZ9XZbWUj2VM1m2wje2lrWfX9zOVtpCz6zLUajpyp+zITJsqp4iDB
+6ZcUAIrhI/PRGwdvWroIZ4OGzJ3IbEeMrwBgawdUEFwDQIsG6N7EoXhK6dUyf+9
BsPv6504f3MRzNvNqvFXcv8ZGTOb0x97BtpBx0/+Leqz+S65OM7suvltrk0/66dw
2p0oy3pVraCYF+HyZnnndkSFyxMs8kXhNAi7p5Fr5xxlnIM5szb71nuWm7BTtw5/
HAhTAtjGvZEmOZLodDci7EV2oN4sogJKwjJ8Wy5Vu3x31aqtn3pthEMfeO788BiM
Ell2nBgJKqqYt9oYbYZH1PZcmEtHUq/KHt3TqkxOxBQpV3LCyXalhc9xPUR/NCLV
CELRuqiC3KJ651W44NOx3zeOxKhBDgm8c3s7rkNQ6Fwls6lmpAbbpFph+GjC0IwL
rL3pIOiJNH2V7IJufcBfAbPAAdTe0cWwJD34BHe9VGlk7FeEN3CltHFnIynTFNPg
A9rzxZglDWagsdSsdeq6YijcfJj183eHqpb6YDSC+mskftzKzUhQFQ5CDKfOq2Ei
hy770FjUGcArDjSWVXu2SBw6FR32pr/rHJsyUjQGukLU4Yxyas8o8A8eIM8I4oia
EIEhgw/4iFE6PlczYhMePfl9K3hS7rKHexK6i8EoPpW6fKHMlp/t0HwOpk6g6krc
vu7B4QUHY9fOiOq0NwWj7LUiPuZduR5IPVxUi6Ha34ICBbXG94ZcEg/iZvjKE3Zn
TuEa7+RnTuz2tO9hrh1exHRBBl3PAmg5YdKH9GNdV+7mFA33Lvewirnd3u7kmKkA
i5VaHqxBKNA+zkGkeXy8MfdP/A+3LmkbiEOLfRgGfcFNjOM91cZNk8ovwLjfPkZW
h3kdjRceZybOrshLGId7UVMdAgKw+fkKyRl1RiXtVeudyMtgM42m4kVNty6XMp3o
lTvqsND5Q1f+Fsb50G0N2hw3Txbs1b6pQTCfO9I8+gYS7VKjMG57A2UUF7syIoLr
kg7QQr6Z6sAnVHzAKGhQKA1GkCve8maUYvoQkcVUdUB7odCDZGB9u0JD53KBFI7j
ZcF208TbsohykhFMYYjLSc+b0yttZjQbfamBXu0VOjDDIO26nN1OfBh/2QLAgAhK
hrNpL1jP+IcTT2kuDY8Ltp4wTWY6ljYEZ+hFWMJrDGDJfBNdscjp0PVW7DYro7c0
jHruiIjXbBqQKgJIpn/j1bcarthM+pci3DHj66Xi/rgCXIWx6IPuBJmb3yQdZWAG
aKWjtHKSij3niLcF3joz3y+zWyHite2d+GT3OXOj7O6Cyj1eNWGV7J+sqL61nInx
/GhSNSDAK8SVAF5XFqkktbdRplOt0JrMBNobsdQI7AAPTZ5kGkSRFFRX5hLqtk5s
ku762bEBr8us0VNKil5bIXvsjM6Y4mKv1c9lLDquK8Uuk2yAnJI3wbDvS0F2+hU2
Tpv6gjtZoyygedowHh5mRtCYvSvzsyxMKe7A6TAFsahgSg3H31ntfyQ1HOhuEBj5
B4uchfx32YneeKX4Owpk39wCpYf/84zZt7yDWqy/OUft5LyBtrBSlbbk7GBRL6JI
mSOldV6Nb3XqfueYgYqAS6RJaVDAFP1WsZRnQ0QvIDYi6YoP3/jm/IO93cE8J1tZ
bdXDNFUW5666NDBJFx3zQznqm99bDIYeSxjctneCRgrWdLEOJho4R3yIO7+5BV0z
2myHAEzcIi8PpCKi3uFuwLoKBp/rihk5a6tNoRm9PoAWfAsAkJRanU2dlGdUDdGD
h2csug6//oghTdpcINf0jxAE7ePuxKuFVs97qZUXzYyt6KZ9ZrInOMlnZdbMpDIE
Ui3dUb9cEx3tBPoFzlmaPpP29SiOOUlVjkb8lMHslcKhSqr2xv1TcEITGtRccihx
zp0GarRtI+kXOgZsJMbbJQwBpq9n3UVtWzHl51YVGno43OBMa+ZoGACSS5XXzMX5
fJL2nueWhnHxzzCjKsybJMxcYCuRmVjtx1TB2UvBCyGxgmyR+vQWheWWOY8fcRBz
rR3ClCqVyZrJQVky7FijvaLQVdSIq0Acvbag0nYykBdvxku8bk5qVv/hzozllHEJ
eIPmZrWzfss7gewFQIWDzUBoBikEnlazi3Ar5hN1bYSdE5ijK2jeM8NuNelLDUx8
AfjB+UOGat0tulYiB08PfDwFex9KKgd+AFaEVf+gy7KS3uVNHOy7alUh7IHrNDge
O+HBjv1ycStcKuxFTG6qdWPLYHGmmWIHuJUPxjKjYXYBtWQOTfjuPBxnyfpY718i
rLwBz3kvs8g4BJSTXaqKME1z2BNTaoXM32QlczZL3fQtS+Afn/WmmOPQ8+siFfnw
AItKqbvLwdedLu0T16SZM5A1w3dKLXzrxCFkCzExK3wFqjIu3OkQGRy0GQFekx+J
mSFnV/7Z4lCPK1Az+XBQ7ORzApczyVnrqo/oZm/TCUuMRUIFWTFnpuGzFeMMfADs
Do8AwvTa+2kibPW1Zc7BOBiullDS/NchOIB+Xz39F3/trz3v+GT9DIKP900qH95P
702mgp7FB2t3dvdHkGSLweCW3s0wYC52EQN/Se33zZnNsRnLY5bGPmaoxjGwjQXg
lPi4rMaE3jSUuiM5yPv9su8/75fqRE95H4SiGkcg9DCbqTlczgOR5FhrYE2TWY+c
mHuBxI3clXFejlAmbmoZTwvPqfzhrFPijhmkR1Pt6Wo146brcs6IdMeW30zyWMuo
Pi2l9riCBR/89+F4rOmIJE6ail1sLSB0+0duAC5rzkxHL+F6zfFhgJkUhf9tTI5E
Q5z0jdK2oSI41AWL6E++6eSOvafxtdz+ad01sEaadls7ibfpkSa0ZZ9AOFQA861l
UTYVomRZ3eIkqOLbu4jkTqpzWA6aZGpthuaRvHzfRs1IVMgtosUsWj3ncW2C1EE8
YZTtKrejfPs95rDAvHcZxuR7lFpww2lMlwh/7ytVkF9N22FupLNrbYwIH0OOY3LM
OioNQmUTT4L4M3u4m9Z5HLgS2X4EiQAZNxwfmsSHqtpP1s4MRU4UBep+agMsmHzC
Axx5xNSnIsFJ2MsVDkmkB5ImFMN/Y9LaBuEMRu+MqhZD3/fz32npc7REMgP1m8qh
H7z+AO+h9f3tj+H8ysEHCq8WzrdK7z44Y/5mblB8vv+uwfib/pWNgt24bxNruPRS
9z22TF9v5OTfEvA+gghAA02gLwhQg6P65Wi+4dGmVJz5+lJkbXeToDn8R2tSwoxF
P3fXKJZCahJ1ErSJlNAgDVJxHgo54Si8G5wJwjBY9MYnwv8AQolkNcs9VB7tca5g
lLZoG/Kio5mL8lQOqo/wNJyDGQmbPCwdOmrns8clP5S5YMSMHGn+rS35D4JOxNNR
Yna8RrJmEmZQv+WIZ+f6XOdFdfMqjWH2OqsKFB0G4tnnSVjBjatiH3drr74CvPYS
EAn6v4UL4hz2MqlZ6DqJtoDS/uwufylv0EJdBca+I7cJd0NkH+Af6Qw06ixsFnpU
JHh3+tTQEt/ccNp9dqsMN4gMxfY4CZQa8xHTpP5S8VbK+mzpG/QO2XOodm+4SIBT
9ym2SxgbfW4eMnseSS02PTRaCCl6j3orvx9ibWvEuW9XYEEHE+q924LvS4VtD4TN
i7Tm3jdXplLsk+IAE8erdBjTrl7uTKOAOlg9kRl41fjH93ZBO0YEb3I6cEwYL5Wq
yNfqZXwXSxmBXd5VHGkiPUSO2lbuowywxaRLd1MZ56er+Z289iq9SP+bZd301TzA
z+LwktdlfVKT4+b5O5qBryxG/u0822vpsScojm2DA+kudOBLymGVtZzuW08Gt2wv
pjpCgVSZnJoP7p4NMI2RMa4uQA82VMseUNTrLSLrlC+pdRc/pfSmx/1r7moFO9WA
MKsIaGRSb33Yo9OYTbYXo7lnO5nLmLREdoF61kHYRjsDSgRtBcVVr+8xGObYNvTd
vpw+dmLYXilVhq4wcz6Wc6FNAVQDYWuY6wD8PbXvLQ/OO6XgbDIeOwMFQ0TCRB/K
gt0YGLuV7AkAeHVC42j2G7M14Q0cAuqA/O5f3ty0cYxqe17SrvoX3lg4A/PfOg+/
xXO0J6b6lN6iahbM7i8+lFSpNn6Mb0fV6U8Ue48qx70fuYkbUPCv8h4n4/WYH5ru
UcX+kG3DQX2QcZjlz4y3s0xgcOGg7eXbkX2unx4+NIsSa39M+DhHe5eslyiVaqfb
L6dHwyitOp+uq1J1xKWDvSkJCvUWmxToRZDWtAW6TJd+4O/ELn66ggagNgEcBUvQ
RWdp+5xnK9PE0nfUTSE9o9CZboyLQ1JAFbO3uCapI8gJGtWfmfO1zcPtUVQvDHvZ
ObjtgxQeqT8zBh5HxV4mMshKbgeyOwOgsrQjWQuPlMTyokH2BH76IaGEyizwNk6t
0A0/q0o1TZka0d749eGEiYAl0zangYY/QNx1WPgXDpBVsExUMw/SqD7/CS7RPzjF
StV+Gwyv0s93a6XfMA2WbfLQ882srLxJA64pbPXzwcCS7cde5W6BSvqJJeV/x5sL
KvxDtcm7YehRX3w9kYmqTd676vb9IFtudwv1a0b3leroyBhiXD0CXiWcQjDscaOo
JaNTkNgxSgXNst/XdZQQP5HfOxlkv2flFVi1a8dXGh7nC3lgOC5TbsY+7Q9NP+vq
82b139w6AurDyn8eTHfB1skl8RZsfw4tSHyundgiPuPFDPNkYkLrqZ6kymk3gUVC
DOLiubImLw/+xnLFTkzOjl1OeZtd7MyJC4SlM2GmsSjciFNwGb2N9cCiSWU+XZLt
/KBx5wobeDrU1YlQIJGfVuAtGqbvNrh1ypMa041zceQcXbjnMMUBQXD/iH5JOjKY
Iw4iM7aTceTKB9MYS70BM2zvOEvH94tqn898f2Pw2D/jfnfN3DfsVJL7kGpXFIBX
uuyuHSNyjim4wZdBiJML58cbqCSVh3Xkw4RRLvIAmIXfwGSpS9yrSdl5zJ1zmegt
MKbHchvmdfwbFrAZjYpbZeHMW2owmDYkHtA8lAGfpDPtRYnuVIVRkMPRG94wFkvJ
65DFnXC25fmHv0E1NUOU2/8M+oEyc0GR2fghtvgyngLtFeBfcbMMYerETxXs0+vL
QZRKcv51fbvNmkAZH9Y6zTuCnma/CZzq6+j5csW2VzhtVB6gXFYazjZyt24cxfKz
9LwbJP60tk/MBtfyX2Son7ZowTB2xzKVkk0zxwMBRoMZRxk0mRLN5u9QlmKmdzTu
GA6wtRFQW+a1BdupxYsbZaGW1doaUyZ/Wn6iec6WGS0BaYCd0Nu8Z0gQ1ZgYUaLk
edJJgDtiDq8PbJ8X+e5ho0TmEc0X3jRtr3bbibryxS7rIPS7+TNTXO0qv8wJe43I
hX8iUqHXy+iPbH2Lx44kpRncucXUNTN66gWHgyuseATfbayOEE9GbWt1PwtFAnGJ
YlzZaTL3i8dCTPbjeeNbMeLnB+r2VFksViAceI5OVk9jjrxcLqiLD0DgTAEf2HMS
cfJ6Yft0zrP5zzi8WaUO4Wfw/GeXmG0sLTCiSMKYSD1kmQeporxpbX0xSYfhq1kC
NWjS7marznyaP3acyudWrcYePcqoa+aMsw05AF4C4jlKjXRfyi7e8AMf3MvD/i4C
tEMxxcvN02fiKfVroi7X+edx9i/exF0mPXaUXHf1+LDj4B0wY80+zkS6bZYTC1B3
YQLG6IaGkrjDBszWCb+56AJ5uqhUjPfFrK2XEY9WbbaqMAKl01P8DXdhUBK7Hhm2
ZBRbTHrPlgEemBt8JZdC7R0Bj/t+UzGuboharf1qblkiNDL1NRtzOCMarvozeEIe
+V400BrEZgNaq0Sd/KIbnj7wultf5An+5SqfC8zycOQlhF5bAUWjQX44ED/XELFR
9ahbp0oXf5D1QsZZgbRgFwvhmMLfle3nEaLKMVmQqJOxIdcOs6dRnQSGU2iprht9
rxGota06hWsmpyUWUDoz18vGG7XYa+ChNXXSDHRAafADMDA+p3bjNcA0FnBFxHMl
iQc2A1AxR4AUOeAle8P2X/uRDOntWgx4rVfENC1xZRDj0fJQ3kjmwmkqPE3yXjtx
ggzto69SOzvBk6xrOqkmfjgXCdcrxIq2JdCUs5w21/P7s2Um8/fKBdQXRqn1P648
eNWMWAuCjzXBHTMLdqtKHkVuYGyCEyVEdQdq4WZxpDpN5bAn9WZbVCCfRjkD3QF/
AQbnWkzORO8FfyLVNHu+WWity6iEQTbF4Ev/fpu4xemDJU1IfZjrnqkdt0h4Rjqk
d6EQoPflIwNYzNUJPxrV7uI9kM4BFZcZHkPt9RGfdb9ZH9qKmnif+B9KSVVPc4ss
/oYSopifbY/bU/7o43fGJrLMLbLmohTGb1yuGh0ND1ctKinEERA9RaH3lskQr9xd
8FwGBIx8mbZoSbv84RoylqrgtvxcNemDNGFthZ7S/Q0ywg3HuUGGhc1AhMVasITr
Mj+qMSdDohUn/XVv9cpfzHw0lW9k+t3nxZhKHwj/E0sGZuU0J0TYoYf6UJF80u1m
fQ3se7r2S5PrW2vdg/pTRMmQI5UE3idgx8vaJbcbuLngCRbw5HNjNWm/4auNlqB+
820Jt/6VdhCKxO5+0KTz0YtWow1uFs853h2CHjOKFhtK9WOZFfOmNf9Lwnd7vxiD
PIVdPHnBV4oMvJ/4m1SZcWAdKe0vi+aXz0U4NQdb09QUzFYVvgJTV67KFv+X2b8t
tcDGX+PP3zMZ1R9iN76q2FFdKq64CtApnR6GeoK3K9Cv4o5BBQKknX0HgVMR2uZe
IKA+NuO5LmVZ5Orq5iJfZSpLwGt3PSIFcxi2R2iyT62UIj7rUJcCjVJ49XDB6U88
0iT9ySWiIlNJm0588WHLaKrAUmxxUQ3r2DmX3GrE6KEcDQ5K7SM3DxQT5eZ7Ioqw
JPZOmTxFiqzynX5Y7etdJgJQXXALBOL4OW++oEQG9c99qHsMf799DpwmGlYPDI7d
DFsTcA49sc/BRPEBaDuqylvUr8NsYbiGL11Z6WjFbv72HLJEdHXaHEqDLcH/MXTc
UjoejrSpkH1qaMndOwRVal/6nUXNHbakL930x4Flf4q2ddPs58udvyot8Ra+txk8
tUAWzGfYkYngsZLP/bQVBBrzEkcM5CFesYTDSem5hnR5Fw2I+FlAGn52bzDh3ILz
U6ek6XzLpAiJ0uJLKQUazbKyAEoe8yYrY476pTlbQoiq75AiJELvRFionTW/xxIT
LFTSlpXoi+8mugIDY82y4yG3IMESKKKwSZgaFJToT/LAqnm5P+bQMyJVTqJOg7z6
x1lxMzBvdgBKit2st/EL0YQqsDBaInXjQLoyklhhDARDBayAohY4DuCJ2qXRO2zd
+ZLv8G62e6bPKs3OhzreRrvPyZHa/cw+aq2NvjoKC3II0EIN16vq6dxi+VoI37SG
AXANi5Tm20HJc1N6f2glTBJ1F+2Bh6hjc2PA3kAXF0l/arz0jrwS0wVVAbUOUIwM
jxBH+Xn3vWp+4O2YruiFpfxhIkIGQbAtSd5D6laUiUT5zIupdSv4QJhcgk+lWt1L
o6uP0my898K5BU/MlNVqntVzvW555JOUfZrmqLhaG72SW01FD3SpYlCrl+z0pUPk
EuRoacv0NMC0m6DijscVZjkRg+hc4NBc4x148RFdHRpOeVXWUiFoLpXYK8fxqkKz
1SJVHCFhTGxJpjrLn/853i8DmUF/oWEPD7lW8o/tDt2Oaz7oXfTL3xT/Vs4mIfcB
QXmSeTyZ1nevH0YaPTboZFGIsoxfEABMC+igYfEUpm/4cfJlzV2FiW8GFziE8KOK
BRcasQxnwWy86vvEJywX3J9rGe4H6/AdyCkDn7FyL1wtZ/TIBuQcDgzP4/Xvk1vy
DnfHjq8uvTKv9eiskpoijRguPx1q0/7uOvxH9zpJOvybdz3bdxRUVRww4FxVTd9u
qM/nBuYkV4i9miz8V/t56Weu/w4dakrNkSRu2Z2++Vu4YcYXAYal0JVq0ryp+xtp
i3iIPzRRdDPD4Qn8/fSLMdNTVYGCpnAGRwsrf+FfNcorJCGu6ayijn4h0oEdxgoo
Tct20sakNUHsZ3o7yuc8BX6UP3xtGSP64L5/gRm0Ycs8SZZInPKtwCt8DlXqbyps
bZISqMz6zS2u+nF7gDtgTAOfACVkW3DUGyoUFC9/kAMZlX9ppm3yaxb1068mbL/7
tU6EnkcWiakwdLG8TY8n7qRzs/W+ImFZKlwm74e3Kte3jdpsqdtHpIVSp39Ka+Q5
qMUA2K6bk09de4WiJGAe3h8d33+wmHiuGZsNHolvk0I6lcBBHs3+NXS5pCDAYUbr
PyMwrZ/kFg/0ESNWj82n3pBJ5FpSEvo9N+Q2khZQ+GT5ZLml8sfpVaHqLUjxfIb6
kSMce039HqL3lr6LCy27ht3KrOQF/14K/R1uCPmcZRrfkwbGT+3CBMVWgHoBlP7q
JKDE++aZfmQpc2yLaxws1r4SiDTebRVopmLXoPOoMff2LqWKTly6Zt+YAxw3I7jM
iRf4Lr4Hg1ee8MHFww3DGlkJioCdAAarpiBO+8QNbKhmd9/EbT8RQ9+QvtnOhFuZ
kGLACNoxtmL/qBeOMcRtugU74cQ5EWRSXIUBnzae7lDd9R4WHEP3gTRd82RYIiqh
kicns8SAYyjpL+NnkN7RiwHla0K6F0N7NcPkIp6gCaUC5rtmtNNFDbmFDoRsYb2E
GC2lvffvFFAXqojCvguQyprFrm7xvejp8BKudBsWV798HmZcMJBg2/a4Il+moGKy
/youkUlhTVHcPpbZAbDUk4L3YTrluvAygWezkBs3RCjsPLcNaXRw3gHvLXkH6+75
DDKYKc+jIpYZrPPmPB+bS8zIt0r0aKZp2ud7aBKVWRDx8ST0t+jPZ6YkMJSw0dGM
/5A0wCZAgOFKsMpW7Msizxy4BIAhWEy77oNn0OJKGANNL/f2fQZNbwfQEemvEM7/
j8a9ZtHyNYcolOfdGo2eZyQ8M6fESEs2w+pbUtnKjIn5PVQxufWAIFQrWVrf5oOa
FgnzgxyBijCWJPW/EXI7wKtE/1UOsG+h+0pRzhfOTWk7iettd51Mb1fCbEgYlHZi
7LgqI7Ve/f1V3wecGRtkeKvvrjEWpLe/gWEITetqJ46E67vcdulBWYAt4UOUlIBG
O1UNpgJCtIKa9KaTXw54U5anNmamZEpVh5yfSja/R/b9r0zpvFwomrEhZ0n2DtoL
YnZ7rP013VaTpaddKYK1jzWFdbyTyjkCwphgh9GsHXKnfNS21YhU3XBtHe9RzYOd
N6Kl4uc1xnjzT6Xr/Fvj4xT38Qc46lHEP6V9slsC4iS7C01Sd08Q+RRpxP1dSp5g
9JXKatwXJomhQj9vgZIdkxYIloapXyITJJUZkMe3Gd4hlFvyg59Zqo+OM3HAvr/M
xZWXxA5D0G7eQ/CLQIg8WpHuACeugkiZy0YtlvFUOs1rpTmGhhBXp+QP2WbKqYuI
f9LDP6Bwy6W5i8nim23yNmtIPZPVV3HNlqE52wS1JcDI+sutfVJlZFnjwpeCDssf
afusEjN9E9usZcuxyArGyupA5mttlJOWTGEcSJ+9Bawg5ipSt3Un8asFDtq4KmJK
3qmwywZRBguWYboZrGQ/E63sQcqybO04gbDxMnvJaQS6Lfrnd9eWtqZNyMB2hAlr
FbWuy06ZENjl/7V5ZjpYLuZuk7Lzzu6JQfXDTpAULIVJcASCtbwV5lsqESrSpeMX
tHkuaIxz98C9wtfU+UhhXfHlbv5/l5M02W3Vd9CS8umnRg4ahT/v+LCs1Gy5Oh7s
Z3LWSLB58o/H/gQ4WX68ES073USeXc2bEsafNK+BKTFZWB7tOoIQUNV9cPkd2yPg
1D7mq7qQ8fUMpDJoBKeiQSoKQmc1eAyWfyVHCpu/Sede3sGAo9BGFw8xF8wj7rW8
KE11m+jUZP2xANwwhzptTQoTSQeUtIPr3EVThT9/W0tg4mWHFgs6+pGqoGESNph+
ao5KxCWMIyQX5wd8nLEJ3S27tSNxQQXxXISrvi6z94wCb91snC24pqZ3utm61258
/2q7iyZq9e21hTUYKVCCrH+F2Pi+kv3qD3GgqDs6A+7JSXDbfWz/r5Ur1+ZHrd/7
bUvqG7t5UXhDAeTtkr4j04e5EepKDJLqAUP3QAIY2H8DETWSBJGrkH10MwYR1M1l
JFITBHvhYbWydTBC9AUrmHMlgBB8Q8MgP0r0NzaN590uMhQpUU730KA19LWaVcZ9
p3jx/rYWTgUwCBCzjOuLZqkFdssmDT/8Kk+wC57a6pagUr7nkBzLvAF44w8V3wOy
IAJJqLpmUoEkIfnYqTZajHSMc7YFvMXgXfXOYog7DjkEB0YW80RiM1JA6KIIorcY
W5FaKcWQVeqiaBY0bBva0Ja57fxu423avVkdKMK82uBv2WN7T+55s3GcukDCnWJ5
tN9A/WYwVIwpw9qCFi28wiU2bOH5dXmVLLJbySvmRf1Lg9+QEyGO7394J4JAP07H
Iw1Qu4NiDUh90ibDEG4nz937u60g2DU2f9Al2dxzPHQBAYkWX1yz4+ZKgyM25KPz
YwrtuTsNhzQOQc4aYC0IRnM5iwPX2rKB8AcZPKwcQehMbG4maLfKycbjSdo64ZiI
esOrFik9jhiIkDFuqXI8ubjSjA9letyF2Y1nPYZHcbgfN40KDgImDFy5witRMR9V
z8Ugybfwvp5u89AYuPNwghPP5e5AJliSufA2CZpenppY+GKhUJDi2FwZh1qGYFAN
c0rnbpm/vJQUHyoStJ2UavgksIggimmZmvXdKfZBdnzvrfNQibw9n8HpSrUHRo1n
Jl8KqKn7ZN95dGXivKrubrozOXoRaG+xCSeCZZM8fOcb0oozorkAAXNI5UBssEUD
S/dhWlK1g14NFhTO1gxqvzmuP0yf76X9l2jrbZT7KsSgWHq/VpXJXEUZF42/VPGM
Wf/49NvDNh65HmOEMEuEW8z3k4bTKS5X6vDLSIpsMBvYj3/Qq9H5F15KymqzDnC4
J4cDOQk+Nw97lpgRDNZJGd0BKB8KEYm+WYCk2Q3vcl6Pyyyp9m0oFuiYbZC7l+h+
pa5OC8jmZfdBRUd3fNVbVoKhWNWBbvjkZMwU9uebmeQkwsDB5v6aPp/Vkb2RVdhY
2/eKJDN3CFcB6S+CurI3W3iVcAyIyX6PP4LqBvm+3wlpdpNjByLJEfX2ckdxjaeg
+LnAmt/Kvo3PqfmFP+5X6Q72B7Tu/VX1+xV3smXyB9I19ficZlYTGJluQ75jurpu
vb9fUjJTYOnYxZeqGdNKCW1hLkM2sPAXn9P+7tO36WJ82a/U3r3VwagYL2j25jZk
2BKoeS0y4dB+ZVoTm1M8uzOFAlboCootKEon8nc2y0/fVir3iIHMi/SawscMPx2Q
Oi+YCK5aYEfBcykP1Cwndn3yzzBkC8vQKhzK/hkBA1HHJaaBeNSdohqSRnOk3PT7
onv7Wi5QZ5E98ybsKq3hpTm3H396ZGDMqyvuLlMMuROPQp7s6VXWdumX1ODdP7fR
wzb2ZzSstR01opPAgXZfJtMLZ4IIXPtnp7ljTtRVdRmrEhwodfW9CZN28Sq+xAcH
Z+ruXCyKDeJn/I8sYga6iFhAjwxWokYMdrwdeES2mBZPbixGMmcShEWBnMeEQigJ
p7YC1DFTY6kHZQoSj+Nm5wFdyHF/ZheGciKcmfffn+YYihYyZ8NbwYoX3hrsL1Yk
yHVoDuu6UVxRPW+4lrBa7NqH2i0Irh0zzbhP5Chc0z9cG5V+FMVtmattaymSAUBo
fzJWB6aoGqcvbjqFXmVF/Rzd0JBR/NR12xO8SOJ89FONJ+KetRQ3dt8Dk8KgCDUB
nldD7C2Dn58PecKwIS4I6dDhxrvDjOwKkwi3F8IeMzIciJBrReybM17MGRf0tBeO
RLghc8UkP90FIIB7bqpt+CT3nlErWD5O4b8bmT2mojByePNc50/yBaae/pAe86zo
Mo38TkZvF2DrxGgp2xYB5uyxrdWQnr4Z+4eF9a+vl5ffetS3KgRlYFDRUlwPTG8/
MtZ42cNa0Gs9K8pUvod9YKzRjXc2FAz2Y2n7TxLgWFe19gA4TthDNNChSxlgLcLM
wXprlFNeurv7wNc274vC2/qLX+ymp7LI+kRnzrE/Ro6ph+r1GRpHHaA7n7TBOiPH
m2r0I61IOqjuK2V+O2OWnh2PI4A6deW/dIAFgjMYJPtSEObRi0JmPEyK32hyvYhJ
NS2p6pTN7Om7+dpevjnCAW8d+xywhADsm8n6L3qHDrbDxe+O/BTH0XOFUXk9jZNK
HLyMUMOLW6v41u9dW5/d5kx5zIEb/8vjSS62P9k4ZpfTDXGtQsCVKhLzYdyewrts
Jog0U9bd69aI2VpYEkvQrD/+7NFT8dArbMf+LYe8k9Qqmg0zsyd9FI/jaiQVpABz
zkdwzeXomtcVyBKMNruM4WqhO59juIXYxPM+vZT2n1tboYl6gdwfT2EGxs2ib3Qr
ucsXv2jeSNxzbAqIY2EBTMJvYwj5gLqFhxM7v7ByuhTguO9W4iCnLNF8m3OExSBU
YyBWRHXUGVz2futhQBbJWDjXcAFrBEofj24AixbU99zL7w9FeU1+RSq0PxhTaeUi
xUuk/I1pDLkRytKzUAn3znJoj1SgkcqntFvpnJ1UkbjO2MWmMfkPvXPRybHP+oBw
GXbRZT/ujabMkYuatOmDTrOu8e49KKB/yElyKEkzqqsId47Hn/cikp7psUSYRG3D
eVrr8RQjig/JeqQgzMXGlHWGQ+1jUPaEF3qjv5uGriS9oTDVTGkSzmYrTuLrkt61
DfxrrPHfOEhQCAr2yNJz6wwq0/Us81COXUUTF0cT8LwrEy5disXy0+YT1ZVNK4I0
X3otfuocUjo+wSmxyiOncOKscpq8gqT1zNugK7vS8GnOYnoQpV1+i1tYAAgyonYU
gopR7thRgIv2f7C80Jj7AtH69311dCD0hQNeR8B6AFV+w5GU2tjJ9NDZwHkSisrq
7AjIk+Gmp6yhrAExbByCLAjASilpRnbJCu0bg/9puICSbpsocJMDNpv0GvUJpbLS
tqXBdCJwdxVlrv8OIXHO+KW0g0qxPunBlv+S562qPjO7NFTv1UCsFDIbuS8G59XF
BhTAxG5g415RjS4iJQ55REx+fylA25Mo29aV/Ly84Mvs/ZNPlMqts5EK9L581DAv
CCBF9DfI2xNuKjhhGt0pvXcTxQDa0XwsyomLka5rgXBl0gPM9UW37CtsSeLQInPp
tshZXgoQJ+/l/x1XvNZm138BgrYuNCpgP8iJShfyqVlsRQq5o8s+cY4CWnyx/onj
SA2pqorXJzV7WWew2wdEncsKhZLT3jwutpKSNs/wRr0G6tcjbgXwVdq00kRyvOvB
Mn8XKVwOJZdDMy+54q11vajO5K0+n4Ts3VcYZOU6gFHVxl2xnxbu2qxuK9NEgKgJ
9At+IO2TE2rCxFtja0+7ZI8RZuWP+5Sf9fjm11LSnSdD03fcSrerep+EfxNMxr/T
gKFlICLnPd5QaFrqwWAKPKmhmhZu/v85AK8dLvwXbvip7gAXeRk6DOb5Y7E+ItLq
rI8K4UKebDy2xgiNPAB13rKGL5HPx3V68rsNbbiBwWS6Dg6sJu+MC21amr/GTgrD
o6zh+gioKKrsvypNkDvZ7v7kwvbCI3Lh06wDyE6KRXAKPInLgp/SwNUr7VjT+J9V
rFY1yTyI0NRgyjk2Xg9xPufFDp1PXhN91vZP+SVrPo4afy7rINhs07Hb93gDRe/e
5IxMDTn5lfvyQo8N/HvivOMGEg1Ac+J6fmHj9OjGhxpaoGdBn5m+41Je7v5G9nNq
CL80VJQX6itMCcl91jatNFbJ9H8a6zvEDhBpF95tjW08RrGfHPW1RHSsjjVnbqqG
JgI45GuFixHgdXjtBFf0E5Z5RrmbAlH0jEQC86nvPpMpf8jj4KIyP1EbRpisG6Q0
VKMo5wv2UEHuc8gujGsu+Qee0DPynWc7BjeQC1/f2+EYTVfaiguMn69WE71YtVSF
AyvowSmZNRckfk9lWWq+1RIM0m+WF2Q7jUvocYtSrVM6O1sstTK/DXZSAeU8gODM
V/wfPluVWPHSLeH4JuS147JcdjDna2zQ9bRPX7KuFQYWixIkaVyhE9d2PiHbmGGR
KLMQAnNjEDrBiofRMXmm14uQClDvFl6fXfJosrLObRw41c20YI/M5Xql8f2myg5i
B43YCz6Eln+6I0/stq6FRxBebxAoC1Ym0yjcF+E17HKo5rYhv4XEHQaR1JZuX0Cd
mtiBOJIpcVYi0FvdycCJUnsTZ1QbtsNDjJgPhOIHI3oc5JTA3h3UaDn6tBxX0tOs
xcEc9DrkLfUDLS7aaU/gIjgnnDHMMw1dvWpYJNAK5BjKKIbulNF6CJeMNvlGSOAW
G7PPtqfJfqN72GqJwbg0csyHoVmokbIqg0CBB6BgI04IYQdRz+mnWHTuu8WRIjek
guVx7nl/N00sv3COCxk3dRgDYDe0pt9iHiX0Th0SMihZWxMlIBMingy/vt4nRDu+
GIzaLLSQMlykiYuvnoShblHeYXXfxESMxMwz28PbIASVFsY0f2OVMHgIsPfIvU8Z
6zfBbGTyVcKeJmTG0Tuhz7G9Dm9AwW9C/q815q9w7JzOk0EdH50YvA0Apui2xKjJ
XLYdjbX7H68mrr08zt26ZLF5fNx4hlrhjX4VMMfboKnWQQZj4cPzrZGyEWTzqAH1
XLbzHvc9HinRW6UX1T6up035zvt4FbNoKN1uxPijiyegHvEMrmVpznJDZCHgxbva
n67E//T5kO7bRGtIxLByvCM0mY9H0cQ389l8hJMaacamPPOFBpVFL0rdFi7OEXh/
iNF57lygAdYdKjtq3SZMjYRoi3uT+xfB4tFIsfC5w8TP9mfsjnMTuEnKS4xSP+Oi
XqyDHuzbwjJZj9xmBHBocL4o6jKjmVz5FCVO67AWJ3Wn5Er81TLJcI410paAK5L7
2O0hF6KRM7+Kp4fKqLkE5Dh+fR2hcADaQzSZ8qHvgRoJcB+Y3dYJKAUvYBwyTuRu
CVCo+3TTBX+DUikcf5TxZyiu0EEZDHcPzyhcT593pbIEUxDCVeiQztOLg5AjooWh
MhpIunuFDSev45qSL/dmX1c4itpgKm8vYwlTxG96D/7SH63Dt0Iw+vPGumOMvPr8
d89jZZVZ4aPicS+nssHciQQRq3onWRyJknnJhKT2gEIUWzADxCeq4rJ4LBoJQbYU
yO0liftnPwP35v1Dio1S7ks8/wH2gzRu6/6b2nnhYD8U3ip4hR0WYpfU+ETyh7OX
Tu8Q9a2R7quv7xTxm5AI5F3ForPlvChHtM6JjUFEg9U4fM65WBOvMrCvYroJVpmK
xBGB8YVbMhoEdAx3U3eW+si+2QPwayouLjX2ZxFpi1you1JaMEctfkmMZBvBcGSN
w8raljNHlvwUFlgtH4sit37+clzbSGHVeGkbetyskpJukykaOQ/rPJZ5AHpPDJIT
syXytY7NV+U+Hx3yczW7zWoPwY2H1jOEu8bNLtwOM/+6AnCh1uX/Lm0JC7Xl28fF
W6/rfoVT7Syt/5CM15iy4idqQY8+bH2hBy5XIHNKgZPi85scLh6yHhw12JtqwwQQ
PIxwTqqV6NcdBcZxK5eEe9saFu7OjfJg2SizLmymeajqvtCclYgTkq+dyfF4ndLW
uKAmi5w5mpD1qDGwT4EM9L3eyPbwvX5yUS95iF4cpEP8VLodkojpQyT0BtZST8d9
Z+fbZMBn28inR2vsCMSSby4WZffzC86KUSBAlO+83URIp9zErOcI6HVgQi1ElH6P
l4WE6TujfJTshTuAW8jn6lReJHtwGCDuIWiUTQEYh9asFYv7nRHdBJpsvABPZ4po
oq6HLVQmscpAGx8e2hsBKuhAASamFe8KurAjvQFwwUCbwtC2bTFNa8ZMron/VzMh
J6AbNIMAM2RZgoflfgoVZCqCPDwgDNo3vnPe6M2eEp9l1XcEvAubC0F4WnRxbyZ/
RS+mo0aWOBHfMxd815Z3vfQ9qXF5FytmOCgrPoLXk+OCbuhqzyeaUIPglZ5On32S
xX0kkbCFmM5G2dvXKU56YeHnSmYGDfeqNvPDWkN/JSdIV/fbxX5AneWab3cBYq60
AIvjk11I7z8N91RbaR9kr/zouA9rdLJ+LSEV4X2uxEWwBigBlMoZ6jr6gKKEm5zS
rqYv6NpYjoddmYlLt/mjXSoq3NSGgIGh112oktYLeqJyhnayH0SZW7wpYVyNGvez
RlcumFRbSl8ERnU6TZ/8ELlvXwwzmJlUqu9d1NIKL74ejW1pXybunABwbZI3F88Z
EzLufdtFtwFbJfGE1mmCU6HB6+z80u44ToxWvZzZ//K/Su/28gT1wSpAgLz//am+
QyeSa+5gOQH/SxeuVZchwJLoTX1Kf2/GGI2KISU7lcllNsgtuxrOxF6DgZ4zpPOe
siqmijqlR3e04KTLE6G0AqOOLMVzOEWAqBggHPd8CilLIGno6V8/h43K9rj5XZ4E
g1ECsBgA0rYQvSV4LXqffW9Q1lr8FnmOE0K907+HRoZNkpp9uS3BmLAzsIIbgO7y
sh21Pw/EfZoFBCqzqxkdlI5ovqnIdS2WCViTSPBBe32mobf6Ji7gUyZsTL8tngm9
fljPJ6TOl07XBimbWT3YtG2heKxZmuiDF5VGLzK8il96kZlfrYo6PWxaJHhI8Ndp
Q6cdrk74NkhpagqB/lCrIuPtzE85B7YHbqKctV+9v7EeoAHK7tgcs1TYUN60x3jl
YX8NvnTmGhXgUR7EgyrhkCKQI328RxU1mA1rgE2O6Fy2JqWW14eVffp8HuKkxXT5
YO3un6PL6OK+Mz2EVsmP9YpTblXEuq3uIzytjYJmA/tCLqlG5fA+0/RhNAFBiZG4
yPytLQqJxxSy0ix71xVWcGY3Db2/UycqOFtS7nbWl/BTqscii0NIejjBIhRu4PH8
Uum0C1LhVOo2vX1GCp4W6ASee1criFSY1NvvwW78E/4lLM7Y4NXJURgOANxaqjdJ
cOneXSchRql9EWS93oulISIE51W8b2s0jtU+BS45Bntn9jiQw0Lj80Ubk0RAnpa4
XXQYwSyMRfZHUUt+HvDbX6idE1+RG6Ytkm+zt0wyqFO++PVdd5ADoEquXv7BeKau
MCQXc71VNv1HeazfpqjoclB+pJB4AvKOjII322zH4091Hncek5tOqNDegW5yBMsm
zWvKypGfRJ0iGfjhZdkdnifZXvO8iDv3jx4uFe67jLw3+f4h+GiVa76T2D5gkIIe
+OArr1LfKjeLVOK4OwA0nlvB+Kg0+62ons3iXKBSpLyOyT/d3mdY1OTtLM4AH0HY
bbDALYBN1Ukdsh8EywK17tQm4MHS1I0QFfo+LOUJ1wV316rceGhRZq6sa89D6l7C
6B1BceGKoyMRMDqJ5OiJ+Mm9Wu2Sf84OU46O1LoB1bBC58OLI2XLBjpyxB2oazwK
+TgTIadS5+szXaSNPHhWqb9+tCAucImwIEu14/EVwp+JnyVV1e+8pqz/yYhZhI3O
lA58RP6ckIYYzAzwGdodcJTp6eF6jeyBedGJlc9D6Xg8XjtGpU6NTT+wuhd9tv5b
AatrslmrzPimG2eZoKsM/DoB4zHEAhvLExIoE5D5Fx5gzoEXpthZaqgao+SwYjOq
CVfY+LUe+BorkltphndxWC7dCucmtVAaz/igObdVEBoWlejiHZRTwAZrVyo3LD7O
WCvI2xXuR/UwnHlRXFpBXVTUfwphVVK/+YFA9h0mZ7ERFhcMuQeddaj6nO+KZfph
VjVGUQ5PNFhF39R1G20JfFbu/aT2/c0oHC2EOKkbn2j62Wf13rOdeXml5onidt2k
VV4AYldWo5Ew+/ucE8Tx4KwT/JHmyaJ145dfLASDZxYFTRaT5fnf4mRPELlTfKS8
bdOGV4UNsMotvZL0T9m067CKtD8QdT0ZOU2xwgYbY+r/QHmO6FT17Y2hgSEl8qbo
tMPoRLzQnJhJe5t0wuC8iYa2PZ5tq/Sgy38gO1trKANy9nt6Qn5N2yljEVsrcH9m
nsA5Jkj37TKxQOfvWm1nShzsbHbOQ+cFxIgB0elb/iQaY3VZbmQGxsIX8IV6dTV5
iqMP5o4RbKg0iK7TPLz5jiL9w5UoNhB5r5jP3QKFeouZQeOOi3oumHiwEe/WxBYn
czHYcCLwgtRTlvBTWs7mgeK6gbucabkQttz1AyhNdux4RVo0l6djzFqpBQE6Feho
+xiIlz7I5TMakeQ8Zv9vTRz/EW6NqLBj3tGq8HE6vtfqNEoGXrCvFmZEGHF5ticf
OthVwgF0LxlEZQfA8qptdy6Q9B4VtwEIv4SDQ1JJLY/JOSH4l1YkP7RswN50d1Au
R9y3Nz69nq+a029aU24ohPPPUClvO+1urYaEA5ZWyucIZVkusEwXVgV/L/Yf7mZy
CHMj0KffdB80eP7i6Aos7hjXqVVZ0ax5n2SAuQe81ZDjftU0Qz1SoTCOARmZgFBb
WxLlUn3W/CkSgcbzzaUz1DL+oJ2tbaObdFUP4yw61gRAIMIHCEPg6nPnTEJhhvCy
wyrefyAASjIL8qZa3E8jUnRnhJ0PGmhPSpDPCBE+hZ3OnegLz0LN/qFBQW0OpLSf
k+qjYuAs8PWKASmS4q2FHivNJRpVYNL5LHcf4T8A/kRbxVonHbo+dR/ORgCz+sVR
D6oYnraIuWrgd12+amf4O0MKqWP4kHedmutLGQpSva7BFa07wbJGX5V5PJfGcZho
poeKC62pNJVC9PPEpjGdxChU2+oVmn8616CiHuu+EuU9YnxzmUJbIC4dvLck/NE4
VlCowmyTulZozIq/ca3YAnyjiW65fQeL1N7YXhCx5Tl55BoIIsdcp4Xxdk7E/VNd
UqIdyB/n/gyEsfbiO2mUcXRllqoV+wXU6Ll1m84Jc8MCnoQ5WSg9xXmZ9aADio09
piNvy5OTK31g5nt30nqItpLMWN4W13xSVt3AlwtyrSJ1SD/jhgr0i0S0v9eTE2g7
7IrKuNHnZRnEfjqJfzk81bg8S7qil0vyf89x7Inwy1dexIY+FhDT2ju5q9vmyaDi
UmeXRykiRbwzr1whcnvh0W5DsNz3yiUDsk/dvxuCIjW4sEDIxzeS484NiKLmV2SM
ReZ9QNr7T1qz3rWthsw+Qp03Snw1xDvdl9vEDUEfcorZPCHkDaOGw9pX4jfuH1D7
h7BMmRENYSawTdJ+4QhEXioTed6cgn77D3aMFZhyvc6AxOQ6lc7UMehp+nRgqof6
eFhvumeeAxfEhAyGsQNTmJ1/hLgrvLkBbdhE7t8bEFTShTWo2EfkErZ+vNe0Qn/N
h0v6SxTeQk+1FUfSEg6mHQcfCK5pFGkSSy+BClUurw3MkfJYeTaxxRBvkxc8FNdO
HzG9G/m7PWNYeRsiGIuFAk3gembV2rfAv0hv59l0OEObap5w2UHOi1TQB/HPRz7P
tKBciRwWb7wxsgzlDN85YGEy+f6xJ/rzibfR0bqBUddq1RX1/qIBFC+EXYISRzyq
vkgOgm5+x38/6jz0olHZA9lay+s/GSiiflgW2Bdz07KMqOYjj/A0cL5UyStOXGhG
YrOz9L1/Rj34EVoSdcDCPozh0SvPZJHXLV/Y14Yl8TO/hsMI6J6rAjvVPdB6koPl
K/NT2B7JuRKc96mJK7Ja9r+8p39AVubBJw+TaENJ7NyS0nnmUE3+QpIPm6Gy2UOe
6uJwYgYOR9ce0lEy/y87THNXrqYyrfR6MSPky527Ud01Gcxe4y8bxqJ9DSG7qgax
nN/E2zvpPBrzkOTtyQQ0/+Jj7zMeraf3mKrrQSlsc5CH/gMAGl1n4ZAFRKrjws8a
86IWysbeDZTKsewG592kwAJz1Fyf9LkRDxZxD0T0JGX7WwmIxC5enHLHHETN/N2h
e20HCKkXHoP8C3M/OniAxRtpVRUNOofAQ9176v2hRUzXXibpT1MRktAQRo5w6sRn
Zufv4VnC+tJNH5Bzbtc83osdjkhIXnTn4uERJP7E6byK7OC1uEm+2WE3zmMW+N8M
cVhRvFkH42NboL1UN6YjkjZ7pfZQ6NvxlCkhq5SqQzqY9MYzFHfidEuhA3WktwtO
jTnAxomvJ45FIEE7odK+L4oKv3FvkNqzFeYiURvJ3Hj1sYjCvF/B3DdhmpoialRR
oSBDWqM/gG0VXHHXIkSY9HHzv7BHqzO8zd+Le4M/KkYBlpTh0H//jFx7QeZZBcyf
k8rBfEPLbi6MNMpQANe0rkL1pEok/2Usewk2G4eYnfUvKkpwhG0aHyLnKbGMVItm
cgGGl80PdiD/6B2+sNDhjyR2SzfC0QCPSYpV9HoGR8h55Baveb56ZfgXA+w3wFgS
zGXYUx/Nwl974mtzOEPARsr0PPhT//gVm8pXEpgTlFvHVfp/xSdkCJMRxzTsDsBR
AxtI7NV9wQal5gtknR4Da2vni7aA+4jjHJbWmfPBL+/53a7gO8wZM7LYX91of/5t
4b9oMQGhwWO40W9RS+IHZLQt0xBIZX4sa3nAl/DJl2cFkH/QWKG/Up02ZZ82eTZR
DZYbXNBpbFHnVO/miykYNq7J+RAnzXgtox7ZSwePkkF1uwOmfNwjOVqgr7Pw9Ht+
BUnwtxMMt4bd6pvulCGgnV/X6ILpESLyRJ9sbE2VEEpJL5LkMhwP7y8oUXWWvic/
fDx6DylP9HgzKmXOFrxlhfdFQb4Xl1nnOn3g1ZhUsx5rF+mdKKCzTLwbzGZsJP/R
DCrrG6JSYLLbRN7jJjLJgp7OAijBvhFCFDGVgEwYL8FHlDP9arV5rtRIx8ShlfSz
rBbP6Y0sgyym/oJ5yRcLkWDwQJY60bYksPxaFgQP0czpNe795kf6HV2mEaFGGna5
zlKkyZPUzHZA4xYkW6Sggt0tsDGa3OxtBUuytoKj9WWtWZJw+eHxIpiJQaKG3Ddm
1hr2sMVozqI2B9LvGS42FBrqKMJZDJ2vP7t0xcIEdv71Pq5mWaXMozZ2iq9GlGcK
unsMjuRsPrvzJKpizaqhf8pe35YOD7DADGhY1OzE/ultRouMDpQkqZt4FiW5uOtN
n2y0AUe8u7CuNPJS+d5ZcvNIz3Cgkk1XGVC6QmY1ss4W1mB4WQm101/3hVYAeIlI
sj/UuRGaF0CPWDtjuYaVyvWsfGCUgBD3RsisYx8WtMI8WOG6iY2b0mZOCucX8YC3
gLmt8ol5Z5IXqbZnTrBALgepR1a5RecSOvsqy9zKSS7qHySHT/91Bj+U8BohLKQr
70wT3CYIiHCrnUfMpeIoG/KEp0huPY8bxuJDOpR8Fb8dD6Z5ddhiav6KKUnPKwAi
OxBURs75AnE4mx6nLz9vUv8cn+QBkOLiEAMh6YdAvkpeNTLrFzUwvcgzDM0lGe7U
revOxpiloJ8znW/gVEEe+L9vuqFvtiwsqBKY1BHnAYc/6ItbCDaMexM7SWME41V6
wndHk7SASPQ+gMXbChnIgjKaM9mZ5C0D0Kmq5nviqfBVxenulRokE+5SVLYFw/Hy
Oix09q0VHu/006CR9jiJM9z2i8pwHEGe0FWYi7116mALGUjb2++5NOq2fPPZuwWx
o8WeNyF7dhtkDtsXNpgzkGUuhqHaeT/mSsDLxvaAsMUrArddbdwMFOg4vPA4vW7U
L8tW/38NPKKhOhuxz3duE4EbUccDjSY2vlB+jVkcBobbp+OcYnGDhz+52uhXqGWo
laKGKghgy6rxC0C17USIoVoqayfXfcWdtsXOpVSANZsXiQiwRRj0wjBss97FJHBP
0djA5dQt2z8bfqjdcHkL30ZJxl0QxwXCLDTemJPn9PHG/y6qcNGxrQlJzB6s3M/h
PS5fCgKxjQg/s7Lps7lq5TOAloR6hplMzWBCXtrvAlpbhwTR0/e4DRM41UFVGsAh
F4DpQmmAnpP6EVPFtzMqiVr/6D/VNZRZ3z9+iECTYxjV2XN41ZYHT/HTtiwQIsY4
ALryd4pztbEhfytE/qrsy3mhQWsZ5Dj0jdoQO5FrijkwdrENHynG1OL35pUc6nQ6
A3DMevP8kt1YhKr57mOLzJbfAnoon5z5dMD5zT7BpP2xuDDT2t4de5hR4VhsUQK0
zQbhfgRf92j4ECv7eH78veo2o1mUXYUCRCJZN2q14vQgKk/ud1ncJpYt9kcLYf5e
pKbP5aNpycar1KMXsGx+gs/AlFACviRK1d5tiJT0LibM91HC/A4yxwK4OBs8lKfM
wiMg+xrto7ymza6uIFgRR3ikh0opQ02CIsQhOO0D0YuHuhne1NtlCn//lNBnhWxd
F6B4xwdEoKlG7ndiFmg32gyXqsi8/s8NbQbG7vow+GhzBM2B3AV5Xze/7Pyaa6iv
ZxBCSHKa6Lj7RjVr2BcLDshrf1hPOuoDkmM60DD48OnFOWkjJR63mhS78UOSYVYl
iF/B96+rVeR3oBu/4UT5tBCcTqqqknWrHHFrhf3C5/rYwa3SrFGwCWg+an6SECcH
uFznrz3YzvOZ4Df7hE2TA23sn6NwfZ5ct4MgZRDEu00GfhdxmSFX23o5rki1FK4/
JOeBuEFynY8RTAOBaUGvNpoENn1wOgcJFEl1tV94IkXTUX5TSNwf+ggAgAbXpquO
bV+sdHIdDHSmZehmMorPBzQs24UQazJT7LIITcFzRvIylObzsYHOiXkdXjPiKw5w
LCQBM4ctn7p3RXvfQRmFvmcgU3tJth5rO8NLdLTlhhrbNL+Lo7LGpRe4bbRWlapQ
OPOTkwZ73sFKZ2Jz9/pbvh9LqdtsvxecqY0ycYprN7XEXV1atuRk60z3AEqs1OQV
qiPaxR2f3VbQLJ84dv6POgrOK1Mfgx3mjVFlasZRFqwTAtkCDbyn9a0eZIAPKtnm
WiZHa33x85AUproAwaWzoCewbA6hP21C+WYsEaqbw1+VamDUiUfJwtaBUtlktzI8
KV6J+ic+9g74Ggdu/GAufX0mtZdFUaTZG16xK+hPWGbSKIzNbfBXyDeObulgPIKd
7uQfJh7Ko23B1s9TcEwTKN6IN9UQscioMSV7siuB362UDqMO08pnSnFrtDRqQHT1
/OX6kHXsocI8WexSUubNR2/C23eJD8q1f2LSA3PC3Z41dLGkM59NftUpwKA1ayPm
JbrDw63fx2cRv634XuYQtSDxb1xUY/6udy6IfdcLyHw3iSucU3mGW4di4+fCAoUF
6GRKZrl9+W+c2u8pGHLC9hvpcx66FFJC9f81G0LzOpS6+nTAGje2Ca2cmZiRg5m3
Ux9A862p82tPIWa6zXbokI6xK9damYmf3NWIdd/58ms76VMZmL431pPDEg8bQ0pn
LDfzEYCxAzQ4Q7jnIcllv/xygI57bsGDJKl2KszcaXqdxGjsAQbh79W1NbNGDLMF
QX0PDCF+aKCTKCzCwB+1lZMpEaT8PYF00cTN2ZZTIxvJIstnp6STJgHoM+ARtvHu
d/j+E1Aj3LKZcNv0j93HOaF/cmEz1jtmzUKsbRNtwUKBja/Xr4bCLHiHcZel6fAg
n9Yzwg6dRQrLyax5Kl+oNZscbBUSR2Lpy/c246niIGcFV7+y01+h0yoRbrgWTXui
t1ldG60tRT3BX03FHIaNMY8CNd9FxPanFg2tKoJ0SMvC/74BkQ7drmT+rx7ZfyGW
94uH4ruRYF2QQcqZLbVSCpHedmhjl1/7E4B8Pdj7GXr4yxWIuELBkr10uQ+po/Yv
sHUOTteAzX7fQVNyyoBfiuDA8UA2IfvkT3grbim0UUD9qYME6AEdU2JCk4gJ77O5
Qw9v8Ci4datkupEgOEGoe12//RY6hx3ntArLSIc7/okY5yJ83NDuKeupUfPjlrfY
+xxGyDfKy7mUtWHelDjPtxvZgrdb5Otb2EWj0ZUO05SjCAUBsZ4II7Sl0hGA5XhP
7z5Lt2uXlU868HgZRv43QjBRRhePFa4bvQ76udtAnSE2lJU87tdrcTjKzsZjA3w2
lIQuaAfQXYAcL5ug1sAi/AbTVvI+h9Hh5FDGs2hK8+Pr5P+JcGspLLIG7m24dwAV
85YweTtrXqzVehZ/cYirtEHbv8XAH/hHydAyrKEmcrqhAd5/AHvP9PJB6ohQQ3GW
4z2wmkXZQcOBrNbVqjx0bpuPkYAb3Iw+44F5ifOkXHm56sl5Rxo6ZYGlciMxJ8xr
yeedguKXe6dGnvAp38uAK0wf+IS/10VQJF4krKd1/fAf1HTeq3JGehoQDHrgwPMs
8IlF2EOvTCrgONlyGvdOnNWtbIKYExCP32PjEq13WdX+j4GVj6Rv/7xaR5TkKNk0
OvYkHQrTy+I8/hEw9nv5W+wvdw0BysxyFzNGRobS37gMeBhz+oX/Cf+iRcFXYyVC
bLB0y4XNc4PQvJdrRtPLCnXHYYhizFZALSE3vuu5xH3Z3PJYB6UzA9vatHUpzBwE
05Lm4S33qEYG9iEw4vh7AlWKAAcDVgN9iCTe0r+8TIe74dWqkpemPdvTWfzAWg2u
Hog2+1uTMmU3Ei6m9Skc/e6ZDbucPjxOq6waPHnMpIp3SO4U7G3DDkufN3z/NsS1
DY7s8fEh8h4ACxgt6DayyBX55MizbYYm6/mp4fvD2/Oepmm4o2YTS9co4ZXCqxdj
wrZyTB953BRk1JgpZOVzSkL13OloZJV12rrFNM5GytH/AZ7SyOvAicPH28H2SqhD
Vtt4nIYDUkR/Zffq3dn982Q2HKUP9+ognxBDF/nWTBubEUxGN/b5d8+TDekDI8SM
9g8w4y80S+6CuU7bh3QwnzCraJNxX/fmW7+gKTa2CQvq5JjvP5RdfCEaVSqyQsxx
elVbNNGJMsqY+0k4C3f4FgHHIcRjwWgAJkTh7iZ4MieE+e+UppY/QJQNCpPg/Swz
V57uxtjhJjP/oqeyo+Sb48eT/SzssUbbzvlcYEdGDOnwbI3eHFah7DNN4ZnqniZz
FBAsDcO8JAVKMUiC6fjbCL5bcLiB6VkOKY3jeQdgtoXjnkVgHajAwVpeUMP7Psd8
vHQxLcnzwbRhIo7sUkD1U1bon69c0kgM8/bg2EH87/hHOPevhhFiEHR7SnvEAEZC
eb45QGpL2o0d2qguxPxswFLTt6U9vAA+yhjTZLjQWTuiMCHTJU8GXY7YR1O96hdn
EryrXr0ziSYurH/NA+lASzaomEaFAS4JQWv8uiVKiZIAzx2/U6UYevBDqPdtScWd
+GsNqQqOz3UjhgB3vkCqT56QdYDi7+5pUHrQ94b5EhAC2lq5GudzRozKBVcBNeQm
IgODeTkNaT40sB4YDdJ3+Cx5QbhhyB9um0PJh7fwaEkqtf6ijwcHpQMPVvFKuddx
SDUAspp784q3iV+URgSxHRSlvO2Vtj9DHKTNX/lwIuXrJ8H72Vty2SsqbrkEOy4W
PTzGHK55bjZd+219aD3Csy7Uzc9FnLizJruwMQq0tT8Wz5uGpdHRApudlBVB2slB
bEJCgukj3NmxfKGWSMvVujNlYI9H/dUZWajRWuUUOD/Pa+U6MddLSeXj4N2Y7cNz
2hOJ9MtkyTDWm4aRzvugfiONb3BapxqUC9LJJUdSy8w7PgH/qAecsvV2ieuTxLbh
SbhJlACvm1IowfeOv3pOm61bKUUhRrzzodvpHEYLww9JbU+fmj5d/03muJoWHxMd
FxTaZNkqPLVPgSXQoedSST6mdICpjilvhiplYpMFZT5f5mTCb0Y+zskeqklLRevj
CVW4VyL0OVAT9CU7izZ76mRw7o4mFQqPCvusaAE6cb36W5alnEDx/upInxRIU305
Xl+8hRZqVRosfQaFUOgAH5/rraXNeJKZkpVMOtLc0dGuktBtz3leG9P5gbBmEKlw
GwqnRrU9hSUTP7C/aVkqLxEDmgrvs2Ko2ZJu/CD82BAzcwRqQdFQJ5fSVCk4yLns
818LQLI/izM9CVYhJQ2pGMO1XKVTxC+KeyS5I4V0kNNupgWmoiOlNCNsOzXP87Oq
bNPWDyxzKigTMjNJQsTPhz5TFnEUQgFAVf5DuDUJiv6OgAIIAYY45ZinArJG1ys2
MRps7rFCBPGrSjbRQUcluLwafQb9Auk36AYRjJrhH9gWxrps84XG8+IOYAo+ED2E
vVQ/ZAmH7rvBK1MFkKI98lFVH5PZXy2Ymy2mgiVqFOjmIObIPy2zOCkm5yRvw+yv
RcYUGDu+7vsx7atG+C7rpBdXCQOlXAVb3R94Fb7utMAXVujei+g8SgHQVLrXb52i
CPKy9Mg/BfB6kPYzCc9gInjDVVRnm/VfI1p3PJIi74T00SaUJGwDP79SaCuQX+Lc
ZCueZVXgF/QTOZkeQkRrzGOpMZPWkqIyU91MgwNy4GRFSw4KTtitNJHQXh1VLVKF
5fWLK8rln37OL/HrwNDhoKtDQQE8nqOkauoCqb8ZLxKP1MMhRRMWcYCuHCNm3dCn
rr355c2MQUB0AelG4TR4bz2M58JpkkeeGoei7msERNGKGZ4ogseFsu6apkC5WAEm
FWRehbxPr6gIixbZohik2WCywRwZnfXtCF5yLixKw8qBczw3GCViArvNjqxsoevk
KQErSUGlxdMRKQe/zmw8Q1TlAqFcqKeHpO5TNt46zHhj6+wxIf0XXpAek9JMWu8E
fyfcd8RxzM07buJ1ozCsUSv8rEvcgwkUznWaJiep8JxlVHdkXwW47V23HO1lKVcq
zM3LwllRFHYnjJvrej88oKpFvkalWlWhBiD5MQkmNMq2tHEcU284gmWYl5cJXJfM
l0jPtwXqcAF1aQ1GwJg1UWijeax+QhCWDHKvb5I/GWdcWez6eje8mT01wz/7hR0A
JlRpFqvixxJeeGvchXT2JNwtkPyLJzzFzfy4mlJgg2jG10QuXx92wjeRODFYXqPR
4d2DqtHsRFmeEknTdElWC0ea6a+gHzkd20QyBfICt/LVvihWdrvK7lLPatEw/d1M
Qo2/oK3Dbd+TqbW1tnasEV9CV4fmjVweTFdENz9F5q0xX+IVreWnAMZVMvc/CUFK
WSp99fOiGYnuTZcc6/CHtQfQOjJbWsZ5qLRjwEPVu+fOoQIWOkOl68+Dgj+2jTWb
ITMRXjysgKopB8EUY6o/Yt1u5sZEkcE1dHwGyszN9wXnH4F8xrFir6imzFtoogMe
9gkKfY+X49jTmsH1eF+0HWTndWeUQ7Eqc49EHpdFiZwyc5rABuoeYVQBb4oq+Sa3
uOz37J8cNnjy+LGQYy/UgzNAYMwz8P4/kfsDokOaxN3359qcVEH3/vupTrMtbntM
K/HsatFILbERVCy+bfaKb/VgXud8+zj2uiIW/8uWrkmioOZCXhTaJa2b9lTjHNNs
hsWofhy9M7CwYFjkrdb+4uhV7qg4kh++cqMSlHhPm2p6tmUbjHLKWSF0Kv7g7lv5
XnhIpuzqmUjRgSxF+hhZko/kwqctUzOwMeLOsLz+yK5dpjy0bnAmftDy8A0jiWVN
ob1dF96jDCh0cevpdiZXwlvBhLi3aQUz4eFe0eFLaENN0ROPdw0eiLwB3i7SMNU8
XXw2Z8D/FE4YuFoli5hvz/Ulm2YelqJVbtguryKd5XpMxW0NCZjB5EYC8aDlMgX/
Zt0kwNGHdSxGI6nipEq/aS+LQXTmL7o4S+ahXNCXT62IdSj466mU1S3Dv4nWnIjr
qADVSZWGJExtEdi4NlSZ7SiYmZu14AjS+AimPdWd8XzHRc2/YORejdQh3rVY6tQM
zfE+xV8a4nm1dP60me2SHhG/spON4wMz2at5K+Rg1POW1YLF3HEpO22mX6rmKE4U
uBYr5+QFCoih9gMCD3EX+641bjS5LZ6QL8sVdP/PeMg+D4TpDcozGpZilWkGAYhy
LrP6xBJPR73qufGkOfwXrrPBTTWynLRlsIIzHQJwzsy/GkoV/jLN7WEa0GJ9EzO3
W6COmzDasOi6qZV2UPTJ5zMJX3bnvG5NAyNnY44toS+YKffhtShCoAUqKakxDffJ
3nr9VPweCrV07MM0jQQVsptr3NEyDuzrTNd/YJP3ky0d1/O/6S7G4Ax6u10tzg0K
Ze3nWxuNIh7RuCo99JQFo2WQK8bmOykalazbHToo4g9Xr9KICtm5FbWC2RFgxWQo
gGPR5TmBS7FXKpo7+zY/onq1AF7/Gr6lofOMeiYqRHabhrF86sToGabsmr6LLB55
EoFsnNElgawuj2ojKs4NmBhAnbDFMNgMiwmCayXJss6N/ONxnSXSs8pmBqLnkJqC
dgvCbljZcTW32tjTlA3rZ8y6cDB8P/i7bdzaSiRRUlVoL+plhcBfFVC3bHfFa70N
7e+ui55GFUS/AVv6yiba7vR0FjewDWwnYv7fPH8vh1BAzfpL5O1XUMXQZG52w3GY
NLcr8Mvvuy8Ug3Gv7CofqxQpISLBGPaI/nZ3W0E9kl+sbZWOuqCtW6SFfAAoVE2C
K3sSQUINZq4NbngrvrDrdy9HXsEwuUAhrHaeUgj0ewYQRwx6ca9cagN6ZZyUOmdh
8KMjuha4Tka9YnsFMRxIjqSieomDBxQHzFOvW1vyg/av8wZzbto47KHAj0OLSDaa
S/eJ3gQox5zSqAVo6g8njfPVrRbn4OWSkOWW/HesCDyI4E26qxy8f5oJezat4rHo
NS8UXhOAnQ0/Bcxei7XGkwLNuQDzuBKdoBUj16IHzVezzFUBG93rP20DLq3tNsts
P/acd2sQnzTkhBkp0y616InuwX5Y+j+mpmbhXAO2O2jW6ZWshl1NT2DyKHzKyzCX
VLbsEw26a7FMnJSHWJk8lkwO7XhWuRwWf89f+YzQKsJQ/AjBpGKwNA8Edhsw49nt
H8PdSEN56lyyL4Zz4v5obpAoaz/OpVO1Td/meKnfMB1ciIbLSnggOy6k2t6XHy9Z
spJyASP1amVflTl6+JVV6cnP8fneeYBy5chwJ7YNTu7gMOo//eBjr3T51y+MtLhV
x2G56WyExbmH6g+x5VMf1VBTtiBv7O4DwB3LS9tjDI3Tyel/ruL8Ah0ENzlMV0fE
piPZijLEeJ6SpskrBnL7N/YvWeaENFHM38a/F/Oq0uypMcIrZDeH8b3dPFRzfV0I
NJaEtowr/Agyj/UXs/Mwcv1JgOu8z/biGUR0DvJV2H3COoomSUBdA0ll/WF1C9zs
LDgySkeW8xkY4wwTATcnvBVYMaL5CRr6MmOa5PgGFh3RLgfrb1JFM2isB1GppEbp
fB6+02n6W+yf9xgqnSM3Vi94H5ZULoYQNbh3BimM8/08nM2tV9UjGAT5/29PSEq8
hKNs/W0fw66nkq1n4Hkwi/mTqwf7EL/+CZlXv+OQgz5gVBGDMIDqhwdFR0IA9DHd
JN6a4jjusmHByOAdw2pEQJsZeSwdVBgRV/pA08ebdn7DCY8PdjzsAF1keHUynGR5
+fwEHGbRWnTumof6iQ+62M7Wydnh+22k/a1eGREQFTu3VFAsODj2MSLIijmAyNhm
f4G6+S0mxw3DHeHTbNvN+oXlFBeCj1CfUpv/f6u/5tEazRV+CRwidVzQGls589uh
ltjSIDVhj0cKcSEsiYmVRR92Fn92pOOCg1iAX14l8ow+Io4uuNIzXzjn4pRx12FZ
9CvEan0sDgH5U+GJfIHtOIJdNqLTHS2CocGOgCnJEf5eTseK3rCOH7MXeuCnzzeh
t8cOYPOKbHLewjYrJ8zJtCegLia5e+2scyG5f3mmTQTAJ1LEzjUcePQVOM5VBK/0
vIoz6zHfjR5qVcN1/jKUioV63ZJXdQ6olmwTrdrRoLikKFsEAQ9nEahii/uAvrrc
do2cs/BmgF9qSzkGliM9WZ2tcxA0qbwTyyp6aoitvHHj9s5QpiZ0BKggCzKLGcDK
QQ3MroEnYJAHCBteHbqy/P83wNt+axP5f2/WkfcQPd1tmoB5nKmMRNRIwKYL9duJ
0RH2xkYWRE8Z9RthKMoykyLNBL67sgIxv4eamcs+9SMGO/KFQJrJ/bptf2ehnvD7
eIK0jVOuoZaFon2+CQUreJgMmjkQnZtaJ4rpdJf1zPku1ehuIUHyr0qo1fLeit7Q
QzMGfx2FkVXKhf+I72yZPiQgzLJnO04Kn8MOw73SrRsDLTUztqOu03i1iLmnkhRu
99x5sps6bXIJkgwYtJbvEvPBUFvkf8LNym4AF3L7bOYbbdl0xz7KQiErFkWAyPRf
0ww783DOikLRywOrjpAy91OxcDYZmW1LwRPImj7WJ5YoTeaYtVwcalXa4rWnzU9d
FDK59PdvvjHhQU2D1Z/jpfPoWvIifXUTjJ60V17IqRHSJexcz5PGt7dFmpooKIdq
Bu9RXPnVTfba4yOQv6fZH8n70Mz/sbhzNHg2CmOT0KUQ6wn7olSbWwEcDT6FRPSS
SMPiV5fFiWkWUSsI7PwJMAWpV/ncEP7BiOWN/bahJyqjoHjq+ErlrexKo+ecU7hJ
LWggc7BGLj/Cd/DVLpWkySp+5RHqTG7pZYPwKde296B8WdGPmqg3cBvwAfCLMejF
IjF+7BNWEnOIpc/7KNhWE/XsPwKptu7FUug2tk7gMRj7EVv9Ch6BQDiradur+1/D
BCWsYXYmKcwffv9UryBZ3IKVHVouucWFbHhpdW42+cUpsvW7pt17bR9lz4mazRZ/
hI2mivDr69U1BimN2Ugyru8id7X+zADPETLP/jnC4tSHoTzfgWr7tOtJXkLRzNdV
u7VW7PAAcgeCwI8W5A6K4t7n9WHmxTjLfKthyiJjBEZG7nDcfsGYM6f6ps6mBou0
AZKseJRTgbS3FiG6N27PKHA4DqXs+XEjaMhd0tlyGNl7j4zlyZEoDDUpeLJrcuS0
5ZiGAZo+Ml4XtCcndcXIfo2mNzZyFuOPpgMQ+FvOXVqkHuz/xb+NQV+14mcj/jzR
QBQH4Yj2IWsVAo5jjLtk2S9W7ETupy4lhMzef31volDlFV4w4LEhlyHWzm6r0FX0
3EHPEzYx+acq/CCvfdshTvn8/zX42tMVmNWo3czH9yTyjCkTz2V/sbCPqUzlbfTF
+qmMAkit6hzQYKGQOhzKGhT+LAsnyoDht0H7OY2SCJhK76tSdLOnOBGh2ndDoxSD
/CA3BunPinil3ytBSk0unW34j97+SEAGKa+AzNcHoK3C9Yz4FtoszWi8fdnE6SPN
aVo8GT19oFtJksjB+Qn7sSnp/ucgtBDdvpUXhnpRWzUmvHFIlBwOXnV/qeafYgSN
bHahO7YXq+oLFe/5pPC7TquC05IvxlmSIn1oP/XsDaUHY4jWtRqXsxXXhKf/s5jc
9Spo0Ia0DPSAuNgvF6PTahLekubbY2Pc4RakaCM5ewOlcJXlkLprakTmSzFDm0wT
GUfgNBpKPr0yupts/UCwRmteanhQ6peSCLJvVpjry0+0bJ4dlXf7Xh8bU8+JmILK
7Z3LafpYuWlvT6qCvuWUuN2T0bRswV3EnkOvHo4pRewtYzdMjpfeNvqryCZwdzd9
gP9izA9QbynkgLaIpcxyaA3Sv++V2JK9r4QZbUZWeby+S+j3vpESKKV0hRu77ku6
NAL7nAIe3QrecI8WI1SkE9X58aX19lul7IfFF8vXh0ZSK9oRkO1dmoTjh3rno80E
sO6VG65zjUrWTQl/6vpZVAIKJQ2bA5z2cxdcIz5PR6UN3Hi0pdnWACVoZnVo08ng
x0znG813tbUhD8iq604DlFgvCvq4R+5JqlseAAPbulmbpQDczTPuvJLStG+DL3Xw
HSaot/kwgpqNU0QjWMZDsZW9JqcLMqBRJs/xkuN67naoCMDay71XoOaNLDRzNoHn
7oyU9XCiRZRdHue5tAmaQ/P1dg7o/3t0K5J1LxNg09jPOWuDhJFBcpQuXhSn9zOP
s/BVDWY5d7Fd+kuZdAQQ9aa1idC8E3SEGuLpjlFKUNbBTE9V11/wjIs7sZ/ap7IN
+g2A4ErkA7kZBhg74J+LcRBetf8CGg3qdTlgacWYAbgsVUb7DuYzS3raXFuD4+Jt
JeroYLjnT1MiHC5oY+pi9b4Hm68aD8hzUZc+5LlC93wmTc+gFmJ0kz4ndiIkg4QG
iJjiL1qLfq5iINcXCXzf/2+2XnRGJtURLxJoKy/HNLOrfQLFDfGVucK3wDSFSwiz
zlASyzMqypL+Q3NZnHPMnG2uFL/ChbcZqL8+GzFumbRx6NL+63aJdnestyLr6/S3
MJU3Nxx2vIE+xoHe+8PFc2o+CXuDNa2s6+MsuRrYZdyJXxmxHbZO8BBBvBrpuqLu
aAXED21s9RX8r1EI9fxmV4ftUFhEIXUn0FY+YH5uDr3y6nSRiK1TXXo6dvO3iWfF
jEHZKQIkhm5X2BTGtjfPeCLl42iIVtUFloEx6TltpMnMTQhpCxQeSExOZ0MRJkQ+
w2U4T102USb3L/t/nsf2yzQtK/3i69Q0gP+0FZ/ai0ICv1BKkSKiJIY+3piVskFO
i8BZeRQh801rJKFAXRYoO0FbwuOhu37+GuCjTPnxo3Fsg8ZDtVHxuaGQQpG+M7UQ
NpNLw8pCy5+4P85EGuwyuf5fK4XtF5j4L6N+G381fFaYBOxLnlEfI0ptFtF4adKw
jmlHejTBtYKkUXKqPeiGvk+y6WVjAJ7WTcpbyrbtxKa8I5IUh7jU6X3pRKLFf6rk
q25WzTyHooCWCucJzlFBiGe5t2HwRcBdXtnvjr43MAUnW2FcLVtOSbGTD4NVmCeU
nCUbJOa0sLV3n52gbGS77EnJOOhkQC/U8tMbaq76RIg9WlId1HbqVsZCwViopl/f
t1YexP0Xs09Yb1Urfuo1eCX6IFlqG9hceXbwya3kE+R6WR+FLqK6flwwpqk+yNz2
ELejjM0s20DGz6ksbd3H+fAwgDVBYAf1336IRuRm92W7LpuP5jrmBVr7hXBY4dbA
z9hL4s1gB8g3epuuCQEqHCBlmJIqZuDRfUnKuuRzFnV1AOACMweNfrJvTrIM9ZqG
cmHdCXuDKaE0Rne+nQgsxFte5oKOjKZVZ6j9FW2wcYN4dJRPAQfCsOKrY7nFXMC/
vuefucpC0/2M9ndzmesK6ON4Wg0KhGfu9xdiQtvdkKjPK0tbB2V1PpZhJdNCWMGz
3ROm+J7UjVrimHQnOX2cVoTZDfYtxeMp0iptrYsCzvUUcTDOKtSMX/CQi0r4qszz
5n7o3w6d8FgbQeFwHrv8hCCODCkiXTLYSuyA5zQTR86sHoj1TvEVoc9gs4cpABcn
1EX3e/5sEBSU2tJ0US+l4qecgS3pYBk/vErpt1h3/T+tdp6EEg6tOe682rXpGWYI
q6FklRu2FhynQPmHXDR6w/0yZMaSfNZBTutZ/CndiLtuocyy8dDq1q3NZzA0wXi3
nlnYLIH0ASyDQfod76xk9crB9cWNa9bYBvrlLeNPOjbXA9PMyy1UW3upqYs4jAKZ
11DCkikQNYsY8NR/+g+j/rzMdQmJ4+PAGuf8vCZ5QGGTjBWu/JRIhpnorzAY0ZXH
m45BlwzXRFAzA07HwvLLJxqOi5jxBfgLlro6q3k3DCGv23+kyq8q1u+uWW7+IvfU
uonVPP4zrWm15PxrP+st08IrhrEz5/6pP2645jt19IkfiSd5zZpkD0h962DjEdgX
kQOYFWeUgOYw82qmKd39lFUfE06knRPnOqvMAE6p0qjGsxi+N7j5JpObzcK8SS3X
mpZ3ygh2WJPyDb93VOxHMNfkp7fLXfFZCqdirurj3usi8LR0IP+OkRdPue+1g658
oevagx7plXX2VxTJVJulDLWK9FvHrIn3O0rFTR2VI+9lb5NJSRdjiB2e/wTFdKMi
n6gcXVtbvsZO/gI2c29aolelHxNN2+4tCcw3J6YcjH41Pk01GvgVp8gAMm0T9jnh
w9uOlS9HnXxvezkyfo3Iaiq+9eLAnMcbtZ00TdqmVwG67ulic3mPG7iZuRkX0dA2
2JjQiyZxxOro7M/af+ZtkagF8UskYtrK4asaqPQnvvdseXcbDaNZMEckthtQ2fzQ
OSRQivVoFTVlzPUL2h5mvGTI2fZhFqskBI+sBqz7GYIPomrk3j/o9LqisZjKi22y
PJmuYPGRHmk87JHs7blH9b1E/I9HavoLgZkzRpoGuSO0p5PRiWjBjlHM2pmPNIhS
6DMLWdJ/dAi1GAj9JA3fcdKiSmjMMBUn7DqJ6VzQMTOD6yIPsFw7Sdoc0RFZCes2
9oEjq+4DKtJirf7ch7la/AWLhKbR2Y7va3NE6imgJQopkO2tajTcEKooFN9dYuao
tetwb/1KENJM19loY2A1Yc7N2cOuaK9XT1F+i6mgugzaEV8ehy1B3TSeBPF6HB+p
Pfo51qUdoImxziqMOrdsZnqsdHspKqZH+5pLarE6CpwkISYPeEPefwJs24gvz6f6
boPls8EwmyHwjGgVOwVB7T6DPFgdqAS0flkEgOh3uRBUIomXJtqYGL5HyQJUzwI7
kxIrBnV8NIYt3Ec+Kfo6NOwhTA5XoCjLKeK2PlkbtsMd1qIaG5Zlecs/1qf+DycA
2ITn4cxLllyoZLxLI/KoI5q60nHLWciLeRADPcLs9tOAGxaQT/zoRznA3n8c5ZmZ
KLaWueud8ki5Z8U5iczMm7kNY4rdaNz1rcvi5SyBtgoIRATVJgTfSpi414hfo93B
NA6k4SPDiJGnESx8K/dGLgV4cQ569JX3MKOo5yQ/hZgB5clh31YlictxWKlkXGF7
4m30nZ7kYFfgb86Ob/6dtcVy9qGXtZzf/jrv1kaQliHzQugEsagJ35iHHLD14fTt
JLESHi0iDs4oM2DcBLIdQ8sdqnPf1cWTqsdlpPIb8jMVTBTViu4fa+iLAQ9Pji/F
4kjKDdOjYqeQNywB8d5FiORh1mvzhgsROJ0IrbLRRo/xwyBL0KFL/xpRE5VeRL5q
1HxhnBsoHuQsnQurbuQbaXDlW1IUKglH869tpWC6Y36d5wN09SfnUnn/aK2DVJWo
s8EMEEACykOT8PEkOqOgn5jO5uASR7YGuQwu68WWYPWGBQ5ESRo3H9vbUHmra5vG
XFR34gcsEtUybZrZz75tPwClmx0cfWIJHNLfLf2oMriFvdFY1aTRVKpt6x8v8o01
9KC1nSTss4F3NnmnLiG8PGESACn8eiDjW0zd05sVCg8Ucheon1mMAm0rJ3yF3pWg
xFRFqBLSm3BWYP9d3lyGzqqzWtf1liuR/cKe3gDX8SLwVWIXrKwQfoquGKK8Jh8V
2+jkcVD++1E8p4erXQ5Gf7IL6aqkxZfhA0aWRYq4+R1bKKcVzSY9mn+VRz1e6kR1
/Qa8L8aPa7akRY6rOiA6yPDXnPza0EnxF5tDplM2XMm4flPHFi7w2A+/aOIaj8bo
6v9+GQFHFii9FRVKPiqRSklIt0+aEC4tbA5Pj1aqTvvcazi4goUhD9r7bsFZ6PfX
4xmETA4nmTUQgxq2jFgSLR1O0CTwnKHik1HgguPM3ADzp0j4YiHm+TzPqfP5Dg5d
RVtXK/iFzSo0PAbezboP25jwaAGv01VIcCjoO6hYTwtSm1B7RAqke+3BKFIH7SS3
lFE6NcV9gmVYcYW1JAfdEfdBmJudv/CKGqNWs5EenSP85WgsGuS0iMmH3EI8TAgg
AHVCn1u32d1oP+qwWkDyQcB5NALHokdj1CDv6I2/FAczRDOBBYXXVOroIw/QAlFg
SdoSVIMajdu0nU7LblpI2haDqFgMD4I9JMK3Mj1KdKlGsfmcXhN4ypGEpXO6T4ey
hYvbdVZSc88nEYiLZ0Jsga7gXedNtkY25JCFCT7lRlNXn/dJbTtZ75ZFEmzGfi1g
jy5kUncP/YvBE054W6T/b1XgSJJRO5y1K3aqREkunZG/cPBwAxT8EMcPjykNoAjA
vkgh4ZalHbjbCFuZGs09uKWe32u6dCCqVF702LnNjISvYm9BDKSZBA/pSMGKGPRe
b3H6q6WM6D6mmw+bZyerHYxTm0ivUZdRWg2ClPr2K3lQ/ay9LGWaGQ+3355tKvBY
AH7VwOsktPZd0ffxOivO7Tc3/6TG75LPOunkbkGDMPt8yGS1Fzx2AW1cxWmGlisd
GKlM3fOxmB7aCnXcDKHLtw912lj1qcJwp4GJ28ushoR7uHxrL809XYE5xgAtOkoU
sRPnuZRXc4xh6R0VeukqRpnv+KD6MUaXbhPYaUHNGCEwbFGJrxINtFyr37ZsWYzI
A3BXWsSSUz/Ml+c9vbdo1elap1J92jet5aG3RTc9xJRsktLWureW1Ki3QZYvPKrI
gC1yz6rQiZme1wI9j+rtfeoJV1PwFkfe/Z1pq1jCEB+l/qhOWhAEqdmXNgN5vKma
tbvk3fXm8dLfPzIb12Rtj3ZmlEYqbEFG+GXbkZcWDbvo3HMpl0jI6rC+qU59yen2
DwhKLXRHcUcFgW6KGOjCJOUWsMh77l98wHDsj54icY5OJmJK210c0o9kcAFnVlfP
li74uLsZMn44k0bXw9WzYgIQd25ZwXLfYnMKQCv21W8+E/d2m7JpOSev+4qVLDqr
ViaAeyGBKQ51pfcGOu5R9VKkNCltC6dpDAlRYUeFy2CyY1LN2cqGvNB2R36LdpJ7
1x3sOKkt3tGhnJkaCifW4LkS4LwycuG6zViD3p8K9CQ8HnatBM0pQgDAnQYLeWmk
S6dlr3zOTq1yuMYmLDrRD6QM0Q/tAV/KUPebEN3ctzLv/LbfJja88b4dOmvHcWbV
0jQwvYnU0E38mYubTXBn/Mr+uqId7UtzcdH0D/CjujYRqVKEpdee/IzWcL3OgXPi
vrq9Iw11bwsnY2mcUNg3nBD0TDHvzdQJpOwWac005NLQb+u2Ga+KIAK9IjXnN3PD
3miEMC19Xr0USUB5oEdUTMIaYrLXex5/4TJr3p2lyGOTZHHX698mr79ZADdLbGCz
gvWVzmgwB/3kcgnCgjAfhA26aqmys/VFWcmRhQSS6lJhsctzxSiYLZHgOaEh875d
XlK9e6KFBrAdQKhQyCzCj9aYwNS4Odl02CV8xCajw0f0IIOhYKu5pBsIDfanQ9Tg
orcCbsCaR2aFHJASqXh6uTWZ6NpV8tH2hfxT9sQsalmPau8C5Jm2igLLtcz+5Rqy
0AKer3ZtoLvtrmN2mFbxW3yvO5CBRgo5xBbWm29nObj4u6zvY+78cJ9xFM6ynUms
1mnhUW+0wUwT40KkCRM1GhvgAC+mgH/7WRjWI5Q3pPvCA0NmAur/ViYZH3Tos2iI
3heRyo3hh/zbois8VeGjEGT/Aj5LycBJWnEAt0TIwxMu5jGgmh0LgD8Gm4Xh6rEj
buYOpd810W0bPY7XQ3z5Nu/6k+s8427AtQyCmnDgYnqtelvB11zBObRtPvcGZ80c
ADaBRU2tWhEpdMnioBv2qEQAai6/rzxhOIwJ45VfuoRS/+C4kKAYnbfhmDC3KKNc
T+PlU3B+ywPCR3LppkBK6ksBmIEHr9seynZONcoMUTfe77RPKl6NL9FZ8a8VVA5u
HdQvTfvYr3BhyI9gGaXRSFVKAr9bKoERK0zn8qgoezQh3btfxDafs72QIcTr7gHU
g0Dz8EqDjvooYWfz4dbRAa8Ra1oNeIebMQbu/VEYpESb2Ny7jaSM7hDJ3gvMTn48
5481CsTk0suVYY0MQ30oK6MQHk0M/XfaQq+k8APH7xGt4zf/fXTaL3TovwKojFj2
qwkxjnJQt4yE6mrSWOGbNa1y6172WJR0aqxuoNu8+dBEUN0dIIhBXbQX+V7fCwj3
gsso2TCZAcuS8ovpRQxfAT4nMb8TxavF8phXzASAx6V7O1ZCqI/Xikyl1EFZWv7u
+1Eh8ctkgsZ1zXHjaa5Zhq3QfTqwGv8zi+3Dm1ND22VdhuuK38Qf84jrx1IiWfqd
9k8c6O2IhBxS2PMBP8bXUrd4IsGrtlq04Y3WW33crU48qzKapEFqkKY+M47nWXGN
5moRlDYFLpHz5AB0Y14EHNIA+Bhe17QZUpK2a3sbsKvFOuuj3rfZ1lINU62BPYFO
xs0UMgda8XnlkbHuwQmOXuOhqC/+jtlo8zh0jeuDL/z0NdPsI+ruYHKYIZEh4rtq
hkLYaLc8eSbtUcxVL6GFXsaycm8mA8Dx2PE62OpSPyoFBMrQMHXMgrWMZM3j+5Mx
+FqQDIs077H7LyUaYYUviAeF9SQ7JDMjFW22dRzVv/TB8VnCrcZ8jjhIQA8BIzTa
Y+cbT0yJBEBHozod7p46qrO76Cg85A4/lxnq8OI+s2+gvM7OotrlZqBGEo4qisMr
I/lVFflHVQniGBPwhtnLKm6XqmKy3H9fD6pU8rnYqlMWW1/ITDdQZaMDIOMVGZnE
T3hmmVLPa5dbkouQ6lgMK8F0VUEVVGcsiFnxk5zICs6+WMNW+B9cVyeGf1+mMoIy
5UifymyajgIvQSrG693v5ia541WL/VAu3Jc6RH2D2ofOy05Qev0FoYVuiDTIF48o
5EtrELeuMD7K/Zhfk6ewP5BcSVBPcHVRMdd0513cfl1SI6NculsHlKxVvshtOOyw
Povtp4Kwp0oTW75QXkAxU8/JvRYdYwfuakdKLGJPk/WkyhKfr4hTdtkXT4B8xBEt
FaZn/JSC7oOM4LfPGu+BW6LptDoHAOZ/iKfbbVZNb7EwNwSvamJ4NPS3F1idniOX
Hiyy6B8Z5tjNk/mH/8t9jSgq+ukjctIxPhGMYLr9VDRfVIWTWEw8AFpBer3rUSC9
Prx6sqltb1bptSgcXeg0oRlLw6SehGL54bpsFXW7sUAIyIj40/jCDG2f06ZKoIJZ
F2/KH3ueoJulD93DMrugXMaN8RzVGNgn4VFS9Cg0it8dH/pHyQ2W4VPvMxD7SHOl
+jpihGjILdWOyG3AQIrwxcM3WHmzCk2egdoHAVhzwYe8mKFJXRkKnnh0RKrQFOTZ
YFoQVmjsh0dBRF9ajY0vtN+IZpBwCinbS+8/Oav21w7bu+Uko3nJGvQcaZfXI47e
f2fm3C6KwP6u6/Od8JTKUMyUafC3zY+DobD3YanAOOMl1dqSihHf4hmgJvVTTS/m
Ri/deqHl3evp+6/JYCbxzgL44boktS2UbiHBFyabp/gJlrM5oHemmG7g8mw3jiKE
M3JU9yQb8MHKIwDrekq7YQQTKMYxlBtmb4N1bUmhKbTw/r92RVanBYr5aymD6Yyz
vfN80dGK/56/SLj18RVOS5ZX+0gf1XusuhvwZ1AHI3JsvpGd3yP7sobbPEkP/31o
xHOwXD9yZx1AHH4X4yc6IYquAdUluWSzYbF9i19CKOAG/N7lW05aHE+uuNdHtPgh
PG+v8MKu1b8t8rFoA4YovahtXZom1hAFWhPJc2w/OYzszc+lYPL7vxt6Ack9Jt11
YoP0XpALXeprOV+SG95LF9ZitLazVw9QtY92EeecPw2PpoLG9v8mFTzrQGWwnluR
KpnjhYETP4a2zVoDSDEGRINhr1chiWRLA5F3+q0w/SQGo+ceenG0IOVfmzEFmy8I
sH5vujCFUUwJBFDRH5irjJ+8KjmOUkun38Z/Ee1tVm8RCqDA0cHS9SE2VsPEoO6e
LY0VT730921iN/AYY2QSoP9HSxQR524IG1gQFMhzDmQ5SByTbASExoQ36entdCfI
APxbmeGDvgOiGgu/Z0O0qQEpQAmeD+0qJJUMxF+SuhtvfpRo7nR3LWowI/E8ZIF+
l/ghpLJDrQ5qWSg08J/gdwB1Qou08RIFjqkIXzFuKpUu+hqObvSkF7j4GtVU4KR3
l2c5sB25xQlSoR0GtuJsODc7VSMn9VyMseK/yNXNjdRh1O5RdwEzl9BctaTWe3TA
8LTgtSa6lIgbjyIVUwLxtdl7SGwUvy4u8xJVyFp0RFYrEVRxdvc+3I1iwMAF1rQN
tclvwUwniSxjQh4kerFz0IiFcr5ArSjaABkTNxdbORYiRBz4Yp0MSXVGYaR2RcpF
Z6GWLhF9ubsM+5bO1OTsDZ4yJvPQSjDPmwMjyNKuz2DmI0+2OgO2ivIQD5rUCL4R
Pv64zTSygF2vYWFN/pJ6F7u+181O0CVPjU3sEJV/gic1+TZrFcEtxLg1GIhliKVX
urchOEaL+dItXR11pXh9wInLHuwj6mKftelpVuePBH1vhqVyWeKXdYTpdJ5Ff1c9
+BYh1Vn1sAscdY7qmPtmbpUVcsVRmCefc03Ii3RixxWfYdJz0eF0xXPk0ZBIDTTS
XRZ0fNGiWb0MMZDWMtQVZXfDHAygH9rVJuNBcI37Q85/W5f0sLc+mjIWyfONYzbz
T1rlPEgsYPYRVHPlF1zxbnEyz1h1B47gKERPnFNOXx4JO+bzbIhsUyeXihVGyIj4
YfLwjcEz+iU1t+RA+1EbgT56Lp/VqIpyN38mRM6Lj+OGH03iQT9sII9gsFkg2IPH
udqvfD3HHkU5I06ISMjynkSUxnq8plr+HhCPCqWlwFw4ABHKfq8qUnBDVaTnk+X9
0OeLXRl1CODUrXmo3PLBp/0PMX+X+cSEgmM09XZOEgUlKA78or2x+TD+fP1S+izR
wv2eBl8kB20Dy3DQ3GdOxnMQqy47svEXkfPMLZPPgqlL3F9Nyb0g92CUXZldj/W8
3fQse2dCrK+Rms+UWNH1XI0LwCRTyhhLetTK83sjhcaHTCwkA/EX5q3O9L5yP3og
hzYmCO6/z5RE/abaq55T/cmqCpK15TJIJeLc9k4hz3CBYMm6p74Hzy6iRfTBCzSB
DcvX1BX+qDPX0Xq4tbTExzWAMc/wF/dkmRLnZCT59vPOiql7Lfc0AFr1cnrjhIrM
UoeeOFK0CLAYkjuUUuf56AH2xTopE+pCVKTnbSS2jTumlyZKegB0jG/IO4WxfPE7
ncugEmB6NvtUXq95KwDcPbJm4nAf/hh/Wqv+l4V9hxIqCiUV/1nYCj9bCcn8lFLP
L30p78PRZSxlKbpLlCRGsZUL26SisyFDBlVVz9s5PvoK78F7aNorLfxWOQsHtXlo
HUyC9UwoI2pHHFTaO4k6Lz5hE5AiTM4eYAWepAbKSKnEbAUB3cYDtKPRuO8q04T3
QY+L7PCXMiUGcSjRMfSg5GrHBLs1SbuQEZXN5KxHXREg+usPU/zzSbahqVEuPYNU
ZsQJkBJqkJA/i5vyhDUU+OZyfg6hFeFR6wydvfuQvQR3hwXnWLn7h64Q9t0miWjq
jMQ11T7B0TulP8aE9ZzxeRxPAuBb2XjUb1plGmJt/b+0cmqlNLfJMzHSvSmPLgD1
L64fwttG4jZlokMCOgRdbKJOwxBSVCCrmpkdqvmlam5rQiDvD6sNoSi+gCdPGZBF
3Kri8i8ssnn+r1lRCWX142dsROsnKu5Spdyd3W+N76gyuVANA8vEYra5C2nuKPJu
aeiGRb+W2n98OIx0R9Iu4iQs3Ksz+uSjb0pGgVSKUWnbeyTXkCwgP/Xt/v0E1VFb
XBWfLbCu2ccJeKwdGm3vLpe1xxF+ZfqpDy42GRUsUWEQY2LeyljcDBmlv4UhE6kS
OGq9LZIzBNFEuZf/v+8WbeNYx6vA4ARhKsoteCA/ncpVweJyXyqF1NFOZFjFMrtj
/LJqt8Eakpiz19ElUNzIrqzVQNn8uY9FRQriTM+BrTvuaKhZn/EJvHZ5qPiL361v
SFGLYwfrH3jsDaJDgt0pjuLoVd2bDWlPemPr8gQ+gTCgp0QPq0JSPM27WI/9AanY
i9DtMKpQQFeMLCT1Tz7DIVYszKdEy4+IzjPY630tu3THIqVS09+NRJ9xnjyJAUH9
0YjomghqXxYC/f6rdB3kYhBWlXfnyyr/WY8w8qMwrGGKg+hpJaTA2y45L/REy1Kl
bOMbKAoU03uzYOGUfZb88VpBDT7zuYZmUc5IfvCckRKG2HO7HR+7hRM9h5N1Omww
0HKWwRTYrnq9P/em3wxYiDnKFvttC3WK8QP3b1UxQWYk7v8eZiZLPEUvb0gAlklr
YH/vO7CIbTw5WrmCW4DJY4VI+nLJ1/hNeTA1cAR3bnkKr2yHcDYaM/Mvfs4pPVld
1z8JiUKzj1FZn6zUbxA7GPTP/ChDHjRta676cKz9VdGzR21jCYZNsLMJ5jq6lgWD
JgUf9wqtmAgcG/CXwn3lgB74AgyorBCD/NLUb90gl5vBLI0jOuuG1pFy53BJdeeE
8LBKH77nZ6RvVXWRm0gPD2QHYEwVqB/enyjhXpU/Y7Rz/wEQ9qaC+anitW+8CRe2
aFUMZyLoU0X7Sf5wDjOsoE63eE/AylU/UUu6WWPeabgmBgcL8rRB3Fxt5731Z3+g
1F1bs0if804xzthNEzMhriYtruyR6Aeh+uDQlQKMutNVtr8gsv6qhga++VGqUmbC
PV3Vki9Et8FA8hmN8PpqrH2lMXaRfSxDX7jHnYzsyyIRtWXMbrQwBJEQ5X5jtXWl
SR8+KTKQ42UZrPbDdKwf8YgclvWlkiO41+kRUU8rc2UlppSFCAjphvRD94h7nEuE
YvLIrm1Z6Z3jCfKySq9m8pKHHPBbme/I3TMUO9yFDSNJXPnce0gq0RacqHg89MZJ
TZSoCzH3iahVrxD8Wh3Bn993PxS5mOPsjqTWxwdAeSwoNt4xjIsTw4jGvqjYdNAm
ewtZMuYF4hIjsWSf4FB82loAq0ntLU5CaEMpJ5VYImnG3Uj04MGIZOJwvm0fLlwp
dL/WMptkwxQmNY7fVPApAMsArOjfnSRLuYJ18zOBRdalTTG4D28JZHXa74dWza8m
FuEBDi6wkcFwhhy9e3xAVsDQffj4XpMAHh9bw2tNvBTuoqF+pfIFM415jE6D8HeW
YFl0GdYJlI7+O1lnk/cxlrtjwYSdzTrM26l/MqXxBDIf9bjfPVlFf78PWTmbREnm
NkbWArkxi55TG3Rw7QFr8qvdZ3sdMHRr4qEmLZqIuRURAXNLpa6u79a6Gb4W5xj0
jwyOFr/Z3vvo+Lmh1QndVho8vb9zbtTnDW/blCt1aNm5nzm+4WDSVXT+4EQfGa3u
UGICqzqeNhHY3IobLPr744dK/Z8O8iOAHMWKAYaS0/MnzY4EPUV9Qlfhz5o6FKJ/
6J2fxIrczb+vuv8sakxYDfEKa5NyvLIy3HuInBo8mFjZcHEXdj92HiSFQ9Ba5XE7
OORbafl+PIfpXnVS3fXzk9b053Ux5zmPm7FSX5WPsmve+J5pcxBdmUes0f9YdUBj
BuV4rb72wycvx00A04BFj1pkTjC7qkjvnqUmdU/sHGpDPFiNb5tUuQcZBqgodlqN
iXPWjloVTaubbPVnWc6hLJspnqLfp4oaO3ICd5VyWZV4T+6dM+ABexmq1V4Jddb+
vBZLzttk1T4y0pHmtAKi6V3QMQfTPxJlvOOI8TN66ib65QW7xUpbbikuRTEc2ulu
dI/rn5U6b98k5yrrZXRNCb+mvUkaa3y7d6QjiWfoOSPX+Kx2Pax3840c1zSUSH90
Jblu9c7PEjNCXL7gq9/8QqKOcV2Ik0PzDlD0Lzhr3j8dktMPTvCbVUFbK5gAHACm
skgTy+mbYjAOrJ8otsC9Ltz8gqiFF3OTg8z6fs23rxPO3g5rXS7iAxSJZeeCgP+b
qPvT9lNAKS3wWSBSmuxWJfpl/M/QnJTaIxV+9hF8MC8UA4HyldVOI1f7x7JBHyqT
7Z+b/PVF1lWsI0jRe88nqzrQigEX8DuTcDMiJ/zAavJBySTqF0duJB76of6dGwkn
gcBs2LODP1F+4Lg89j1Iiikv42T+aaG47C4oJJICBu6bmC3yCbfW3yDEsUyxoDD+
CyfCaN8TQQAAb5X3zUJXjl47zFfeh7h/Tqs/Ku748ujA36n98yruB5YaRzf+hcrQ
TM42Goxxs8aMcH4ZgNy6LHDMqD2j6+5L0l83vAwqLV8l6l6S0mj8Mja7XslKTTUZ
JX4nG8v848ctd5XZTAbGvAmDQ0LcwoL+rtACMGoW0NCIeKk93cjor6CZ9DtRWqnJ
IqsDStUfymm/E19wPnvn5gBKDabiEOUWoQU9e2J8Oa7UTVoI3FdoITOJWIDBLpod
/pS5M+gI1QxZxCiv/WE/NqM0YavkOe3U3BEtJeiyLB1OCInxaIftDzKKHy859GkS
CNEJUNgfemzj/JItI9GMT3r9CtGRDuFc/uUtYtA/8WKRMqv2ngY2QAbnuO5cOxaF
p1FdQ2C5CLVfwyf5VaJUrG3Y+OdPdTJiqWzKUjGQYWyeMrDbmLKHR6YYOtdXdCPk
rvh9WdDWXbnjus6FsW3YwYeW9pm1FRwrKSees265DdXXmqbMBxbN25hZZkDTgAtC
6UxXdnz/dtpB6oBPcBCYnuoqgM2i0UfUBc4MoJwxTZfd3qVQLg2A9SUoMOoARqUn
JN6KdAUt7QLq3+ryWQamFt4kUQ3DzC+Z3bVDyDESRnVFz2rDkvef6v61PjQl/xr7
dHtNJnXCsOz3t1RWWjxTYOvZkvxECj8SQQ2ot8acd+yVTe/VBhzfGBXErLlcPaVf
QPhhBCOoS7ym/+Avj9IzujFqxT+qhRPZLzEDIIOyspwQOo7eCZp6VuHFFdJjgPcg
Pz8tuA2H2jC14VbeN/nx4NzbKQxkv9Ctfvtt24IyvOmU2a8qolGFG1g4n8SsN3Q0
p1N0m5X7Q+sWe9FXkklal5qD44RYdxiW8sCGNnGXNyq0JD7MzX6gIWSOUsh60dMj
RYh8uqB6RlUQSnJfJmYbyPu0dQBaYcSBmFPc3D4T1wAfaPzNybNrPKYek7SUcfbW
AJgcVIH5YNslIbNsLz2q8gLrkD0UVS5ojUvqT61vW/M+5ztlxgFry09q0jwqoCMe
b+V7dZRGGTo60LMz7yjvk9PIYfFY/xG2ghqmxXYGNKkK4M7cYe3eolxhjIUqA5sF
XSYSLOG8GIhdtqFW/AnwgaQDyCScq7T4t5El02Gtbx68zyJMNWCCxP+ddW9pDPAv
j9+zYEhsozb2Og3VylfrQNj7CdkjCeHq/8HSkXlV2JswlIGCVUMsJl7PGm7jQyfe
1A8dQqPc0dMJhHR0vUcybz6omci5cXzV5bVQ289rwDVU9P31mEjt9M43gel52ig+
wfe+xfOwGMd7bO6KemPiuk4em9HN0Hbrh/CVXBkSVrC7Yunwbrg5jzoow5hthtM2
NbU8+H71v0zdSQ3GI2vsHtyFB/GehC5Me6OvXKXp/0+VOPRQqyrlp5xm36AqjuB1
4xwu+V0HBoCYoDmhb7aeYCPqm6MRCL28KnQpIq/TG8G3j44BCRWBW0iVXyugc6GA
0FxwfQGHslHqNUOcG+9rClF1/+rbIKwQnK3qjbSRPN/Zcq/lCQW6n+H5Udy4Qjut
oz/j5+731TGanVxXvl/EcNQGDidLMuEwI3HEYpoeyRDndMY7xLi5eQ0IcqWJpAuv
1QTsKax00IyUAqk4wbXci4zEHc+Dbu0ql6E34SV2Oh78nDP4dW3l11t9ci3gIIdU
oUqCqjD9oLT1OYFUtgPUy3PesTWOcaPgnA/Wi8UxRalN1VEMLYbYOtWpPNP/VqQm
pSNYAkG3HSLY/R4rSAxEzMcFN44Kiid5tqWVBg/0ApTfRlmJtphGDIP8CjwMhSOX
QVFrD0N443t/luEyoZ+95AfXdqaof0XmvoFM5BHU1mn7/HkR123WCRbNOV98Ablc
ikaHeD1KMDa0z5gQFYqxkj4ymDBsBWiqQ7W+J+LRpsLmMI82xusu1GsYl7RnEqjP
JfAz9N0rXTgRBNpFn9zL4uEAMysyPz4HFgrasd1yF8tXOhy0d6Anv7DGakBmR0Pa
O+KEHPAtyCaAMO00/JgzGxXJNb5otyq/CS1naplhpUKhMvNUMcQcYQgFZwV057kg
GeBiKmRoTeFEdp0icf/vEmqYKM9zZ9WnwcY/B48ChE4eoUbjaMnlOk3B0NIgKyEd
RD1WGkwg8QIUdQI75ug+0jNl7fL67nNhsEV5v9Vfs1qxyXxJH6VSTENNV9KN8qMR
gQV/LArPFVM+USWrK33x1whofG4GYFkUYHUpUemoKOFcmI6FL5K4ix82NFaXaUp5
BMdgAK6SOovrnyq8R9I9LI3xkoqzD7qTjd5wsg4oatniGbar/b1kfCTI8PLfUJ1X
AqG0ApGSU5bP0kuKOzTEJrwFR0yOMYl0C4ASK0BMUGM7v9JvLjj9SPBCQeBXxLs/
3mvWb4TmXuKVpYFLNtRvSgbKe8BojPcwP5t9fG5sKKa1PcCYpfIEE/ZGDk0D5CnU
0zY7a/15lNo5o6aFW2Y66dlMchMmKYQiBCUVMrbNXW8aV5zhMOx5TYPhpSUMTrYL
XDW2/7Zq3AMQG3UW85NfSiRhoXjOi7aBlrOnGScJm9N1CNzHQeQSlWsPS6jyfpr+
03jUWH1phypgV51P9bdB84au4orQNnYtG4qZDgOo2Kj66JVFOorWBYA2BFJdLrHw
GB3wllonC9CSwD+IGkoSZkdsKsHVEQUzMJN8VZum9VueGLrVdR70ABmbZuky+F9r
5KXgYxrgAnUXq4M1z+XrDFbPv1lrfk3wfbp2kVdpcsFheSzUsZ8gRK8S71fxGqtY
NomquDVy1lh0RWkdxtnlKivXxwo+DJN7YSfxQzAuJFpunj+VJZ2U8YfXQp1u8pIK
3w7f8EXHbbmaAS70Tk7vdWzMDI0uzVLwB2SM/pR2IcHHjgshpR85Pi7rp9wo1IEC
XYZE8xBeJAARYSRJIdWVx96w80nbKdAs13mkej++EgFHuUjNE+Wg3jcYbHPcNJI6
fi2OpGZjqRjzpstjKQ9Hjq4OPiN8MarlZYNjl6/uOEMSCCYjU5kY8JXA7uTLibaM
3FV0FznVquS4aUj9ZS4X561XfeNo8ODGjayD+5938R/9ouzxVdu9hGe6xFjpmEGp
8OFtSvYXie9Q5BsV9RZ4OPIqQusHJw4+Ua07yAv4WxMs49xdKg9HVdy5NO5aNpc7
mM3q5a634hv5rf2/wYoA8aRJ+v/g9/AGNjiqMr4KhO8SSxez5CA5FmFtGmsJRBn3
fT+z7+dSIFTDJUtxfAIABU4/0xJbtRSU7N3rd4bTnLoTCcdsNjf2OVoouFJ0lQ38
RXh2PTB3dhoZVeR+13zKc4LOidXEAmYq2XlTPLdW3Z+1iWWakqyk/+kGjL744if4
iJXrQfccyiLjii4HrNq4A8/P/xjGwNsWBnP3R59ktrerpul/Klw8eusb/Q2hoZ+R
9SUat/pG7NVpeMkdk+qrZ93/7lttw6yI8At2Q3BzGC6QSlZ794EVZGg1bXy0uegu
gFhy/6HcpmHpr2K2b01AjsuzjH7J+ROhifIxKoOvRH8Ym7bi1Xv4HcB2fKeGT6cS
bKx0J30jePD/NendAW9AFt7MZifa69zey4EbThtCMrUv11OqwJyRS7f2966r0uXj
VGN6dCeCgmxEo8khPNbUrMEfV6J3s1hqyJP3OxVddgagev4znMd7VBmO+BYTC8Gl
3v/MMOXYbKYPxMdoHZ7tq9lbwcYrk4sOiVGaaa863j/0hO2KyiJGR3AhV5B0uVne
9TBdCwj2V6g1c3wGd//h/Bl78vV/vBteypeYQWuSH57NzTh1aA9dP0XWkN35F8NX
4xlowPNrr6Am7rtuCsGQB1ToRMddKO2z/g4ZUqu5jP90fm1kIp2tuI9/qG77x7+Z
m/Vf8F5XNurvSWW/g4KKxy/Wofp9824WQSgDEjpVOk6EYMAfBRBlpSFHQNdqUO5l
vMcr3hSg/YWkwYPrtIfa3Jst1rxj5BAMQoPUMByC+OBZirbuk510jOVbDSp8gzJF
OmTu0IX8wQRlrnnb/Lt6CX7ySDi7VKLzmbBK1gDiX1sWrA0yI8Ln5iSeqQUm3kuJ
n2UlGL4q80z6SsXoc1Ardx/drwIiPjYFJQ5xnJWY1RPYtA3NP7RnS+q/5kQkE3Bg
Euyx1l7zkU0JldkWQEI5Iu5PTc6m2cpmNj9nq6Ua8bOabzXb612XKKYRMztXUnPV
kXIeE0QVoD4g33xWNAzjXFORVEa/JcEXmPEU+YzIR+FoBWsLNxr0k0hZcxKY7Z1G
T+EoTEU3gyoBVd17RushohEdNDwfIy6iye4ct8Jk59GFq8nrnTh/9sStH/6jSSWk
2JhV3Z3C+vCKdZcTLfTF5r6mHrj7+6bJyOpdTuC78s83l5nyZgaIjilH+bR105bH
N05DgZIGmciC2qSUs/ASY0/hgbrMqaPTSZkq82AlaYuk+Mgw3h6JANLPS58+uTeH
6hQyjOf5MB/cJ9PzOH9+MxkS4+/9XXvpDiGC253JSk9RiOptX+gtiAk5od/PTrTg
ORky0o4BqBdmrm6P+cEQakMciHsk4LRacp1GKgO9wBpPnsyBdejiChbOqdkhfFhc
S2637l/Ys+whpTPEPkQMi6UFTAPQKyBdeai56Q/PO3PUj0U3z/WkOIaBDWgwEn8Q
5TC5EswqZFBzEShkInRgCyNLaMmlohQANlxY29b9n0EuL86Gt7PAYXpv9UM0y3/4
/BSKO8hbMfQMYY8HlDdOfjSt9eS3Sp0QopG6qr3YjQuuxnV5S2puyorlH+dRd1RU
H0wWd22osM0NJ0OVT8tVdkDwiUuLnai9On4euUw5RtXgozGKob5yJtPknOpBL8Jw
ThTRetZRoVCnXAnEufQ2VdBXzWsaz6dlJCGRVyWvjsxcyU0ofF8AyHXIfRhEGruK
9X3/dB3UMcqtGmWUTbO1FFji9HXn88sGcdd2PqRDgBSDeXI/ZxJHQ1nVBTXqpiSr
l8Tz1yXceEqCDP+QXOgrdFAKodbLJgM58CRow9InkowVqlxHZqQRUdBsxRqy8a07
TF58IADH9qjWmWbnhlmI2EiTQbaEZy3qnjBHASwSI64RiR4A76e/m0AHu9Rf7Egi
hwuE5Z1qSwzR4dS2s33oZFjkSiknK4n8LkR6v1PDupFyhq4G1+UNfb0lJmLeIkA6
7sMb+wECCwgceK5I3/0CaZajv8rrrkElGT84PlYuS+PZEXmDQTvl4X3ZrEggK6/H
wtis1aKLO51aDbG9B7p+IcuueNV17Wj9oT6AQ/CESiOrqj7qJ9njx2Ukt+48tNWT
NyTr/DOveT3/IauKEZfEQvZnFvmegv6Bl/pl6+bhC7dQbKV90vA728JO/FfwsqhD
H3jfIF0cPSDWl7z9qhd0r6vGGW8WdBUHLMzd8ICDvTSrp6KNFMBoal/WZA2lMAVR
uKpQCBvVNgv1nL/l7rRQG2bCzMKoVJgc5iiVRoIdi5cuV6kVUpOS4TL31Y1ea5nF
VYeZcenuOkSFz+4luixEdcEck3MOnJOUuP5YocQ/ZUCc/xP9zi8aYRR38hC1vhG/
pVUlzwpy6toxinPlxhb9Wjx9PGxXGThWpcqeVqNE4yUR/9B6TmcCUQiXawsY6+ks
fgooeiN6NV6SrJxRHlTiIJrTvyGUztVfmBBYVMb8MkEyyMDkeqcCVHoK9E1BpytM
EJtQTgm+GXcL9bEgAFiVFGE9lmDJlgPJLl6kA7k6Zqx/hgUIaTy15iuU/15mG2yC
MS9l8l3yQE8DC5pxUgoN09rTfjnbwehFjRx7Fpf66Jvh8CLB+lian9AzzFWrwJtK
drFKjLbbNnVr9x6qT2cxEeL7KdLpc6fONBBtVD1PrD5gWVksOLTWY++SdbN22K82
Fs4+uoVlkxdUh6tmRmDh8JR8aU6XEOs0cQy/YeyxOoRU45zPVwF9b+QyuSfHHVaz
Vs0HDB1Ncn0s8Jy5j0R1H8UUtnfopLJo+ftKvpoYoEZaOZH7GKuAPWLQ0oDLhjay
fuJCdkSK8tGbqPZ49h0EbzAzwv6Env5tTcfzV7/LSZDnIziirAXH+zTdueGtvE8a
0jhxRCGegkHZZxlMqxauT+Q8vxQUnDVDDnp0AQw1sg70pTUpjWOPPXz50sNnzQaB
S9+LPnnOBCCSEwKqs5pCcc5M/sJFDNDIf8Mk3T/5OlXtv6MTPd9guBzOfdh6XSzG
JtRR0gxqxHvYsfMHbTJuJ9QYSQsPMRddCgxt3ht9tcyW2qlPkPdFPMbCo0+o5iys
yHdwtrNDTm8QnKChSKVGhFT+m/DTAlTwOHUgyW8nu5ukf7Thuib4dGH2d0Evw4k6
3t7Y3I5co0UKufuOYi0tdWujeeDh/6ONoivM8/g+4cg9O0/O3qiAadsT373mlhUI
s6qFVc7gSH0BWO4a2x7aQdpWg7He7y1sd2PZi6mCxHcKoCu/0fPJd3nedLgwMegi
gW9OC161yTsoMoHoRhwoqNxnVm+Bj3i1RbDyXz7/DSVr4qIhDhktQOIKhM2h/I4F
Ujyynn15K9l486hF733/95DpQkwOqmKqxG249fRdh8d5125/ZVKWcqO+yTrxf7BV
q1z7Nuh9i7dHg/Jj8W7aJjlBui6kTYOV2HtKjWPCSsuNXZJICdLUGv64sboKIupZ
xKJeXfFXfUYkqtC022pZAmWS/6NWnLBozhOR6UKE18uloaTd8cg6fGmHRHREyTKJ
AaobSHZ552hb4E9j8uZLGK0NERbw0nlbMH8LTv9AjajsTiAtblRyL6LjKdoxSZVt
SEG507f2jFgc+VSgxk+RWNtPSXSwkCF6Ca6u1khTgcih3tiU+/5UfG/CQMxdr0u+
x7R7vW5acwX50fwTsGrR9Yb2LuGth/WDiesbdZLar/Y5VhuQShTBqFNTpPPq4aib
4pXJ+aES66BS4W5aWw+7ovaU+CPb1KyVqPhoe5sNTqHUD+s43DQ4FkT107KF/Qz1
LmWfnQ8q0kDfxK4+gAj5cqqHck+sSTvPEy0ak8nrjduqxiFkftM63Pw7aRRY+HRn
EP3LPiLhcNBIn7VypHceGkY8ie/x7pWZ38a7HlaAK6I6UQ+d+iHWXv+WjkHTG8wY
2HZD5OeqINHhU3Me8/BqQSH9exTQR2iLEnZ8a2XQHv4r1o9UDtwIbjHP6su3ka4y
OEwW9nOOjnhQ4XZSKEPca0s7r01Iyh/+xEZoDW1OuWAnB8VpBVG8dbXuOBFz3dEv
svXOV47L8ZuSBnD9OHU8uQh4ZDwgl0mc8Q+E8lYyTx/AqkpdGflbqfe/pwErrZOa
gfO1B/4KDnr10CxEe9RPZU6K0hqjz8q22VPj4N1Bj7c/yNdAHIEBOR3hFqsc4RIl
nljWZLgx4NShffYiCmJ8C1NWnPOhBvSw6RMr1xx+4QW6hN7MmP+CJB8A6Almc/u3
R7IenXoBo7PGX0doyMxDLZrHlOa/liUVI42QFHhan51+ibRWS59e4O1mzqiJnh6e
BzmO4HSPjay8aO40RXZvRcIaGz4J3/z/1zgzKFdclgTRxNqmX4cKoefUzOq93MTO
zr4U/Hw3qhYyVS4k8DblIeifR8jRfhBfIRxvaG32Eom4vUF7Jm9xHUWPAcUVpFuB
QaelKUZ+WI6ZO+CsjJBM9VtFHEmTr0JE4K2FV50e6AQeNy6aOBLk6tbRdhGj/7dx
/rm022QOwPX+Ce2qSZaMU8gY9EmDbBkLv0dj9S2vNxwTI0YrE9Tti8mGD1Noq4py
IRBdFcmzpMV1zHuF48I87L+wQzWwYqvVylUSC0WbTGGCji8qHepVmHsSxPDt/p2d
BziTYZQ5uruyDa475jh1uMYNpSNgUYbXXv4SFGh8vJJiqMLIi4XqHJL5ac3AOOUk
2BCnqNsxf5muF+zlltI2hPeniGOuI0KDlyCXW7nJ+7t38o9lMiONQuSJtcokhvK/
4a8GgTCXc0q9wNun3xIP19o99l13Wob2iVSFYwhMeZ25JguKr5lmx4ZMzbZB78+i
VmKuh7P8wDzXYwZQCqHGDFEsUZz+hdIahzf0E0KTwqgfcS7mtHZT9i02ocEiu1gd
2js/SXj2z6LzaUzhrIpgyQIA+WtrrebKMefRCobdo4BQoXQBJ3Q/3ZFxxCVZ+k/H
VucAR74kctv25wBKkkq636uF5m1E317sRcIi0AyKMlOKMNEYTX5CEGTLSE/PSxB+
Dk0Pn447uCzTBHDat3hCUQL6VOX5yB04UCqRVLXb1p4VxHO0H0PjKSj7De5BxqfI
wxp2olskK+KVHYlq7qlzgrMLt8ReieC9NFnXWuSPWbGErcF8g5gRBCCPcKiD8Eeh
XzJhoWBKry1rhy9JWk+KiBBEqsI9yOXPq15B2f00RbBsjsmYnbbiPfmNfqw9hQ4y
2zol9WjZuU3tKHQQ8dw1Un5C3977E3siBJw19Dm8csW8RabTgwnz33NZL2q9wQA5
xvTgTNUqmrXYzULln7rSxjpP544thtv2dUF56EBhu/yv7VciAOUtjT8cToxNzocU
O+Aovr4Qd7zDi15AsxM4XNZ72ayEmotVd+IslQ30hTwCqMVOktZn+8BkIioS9Jxn
FXpZzaMfat4fgdmnRh+6U72exu/XFWCaM/MzsXMgIGhC8KJ1hACr7h2ohrDwW7Yd
lob5Abu7RAszUZBrylc1mSdUPlGbUNYw2lZqSWUD0wGtGilumKLBwjV/NqicWBy8
BLcH6klyXSRLKijdnCMm+A6XQvphasjrTao2eYJPXcCuiaxmwm2DMJgL12b/n9vZ
C3j8bpeXwWt9nkapMPuiGh8LfYbFSbMGdL+sWBLSFxiXB6gjhvtPNTCCFH3TklZe
MmhU7I9JcLWTbJYHtFHoMpjyDNdVr5Raj+ZMDdjYK9foYldZoqJpjibAioyDyomu
E7NZWjaX9/Rmz1aVx2POcVF1KHY9fwrlr9m76rTcuxFkAnU6lW/Xq/JgCa+3tu41
FZrJTUH6rhVf15WkRhQMA/uP4hbsAP9YGKB4frI5wSIdzrn42fI12pXcuB35d7aW
RP0VR+O0H2vu3mxbJBRIGOk05x2BxZL1DZwfDTUuRnkGNm9SPJohyMd2dk78C2wS
XJj9HFk16WP9HYuIrcMdfE6XJ1ldxOMX6NUo2QN9fAzHbA+Z7N6F4jtPbX7uqWLT
YXxSraBZoiDB9SD4OdxBWU4AcyHY/2DPdonAmZk9bJUQUHPxvBusqji96MtC+CWo
oiTg7QPlkeHsxjSEgrTVRwdWvdUDmHDWCOqkv+Rv8/5VvJD4QO+opeNVGReCF/1T
ixBcUGA6pyya/ZBR7T2oqyBWtaSloGRkTgYYNYAb1r8UwwSPTREGXHiWaknpTsez
yA1ZSjHLRc7f/zhQDAB5XuMrfOlkpw3wl0O8W0mkH60QVxPLh0HLTxt2kZoSB41+
cfi5RLi3MGZe8SKfq+29LbpmeqmjaEX/mG4MWC6Bi+SLBTSkjOM8YZO75O5cuj3D
CIkogBCBWgf5idRMgaTSiYwoUVk+/1uTbTtNmHTJXKdejHjTdu97oTi2KqTHgHO7
DRQCtg1rdjZrSNakUR/VP/ygjShX9ZhHCLWMO6OKUEiEhh7/knfFsQjpI7FQvQmk
6mKHI7+1gHRT4KRPaQN9hOGpK25oXGQ8hk1xn+526msU2FDw9uOtjzOg0Pjuq1k7
viwqGsqOHFlbIhLDd8RA52XNXSLNyrytoNpfE/kViAmVxW3Q5lNsTMKZT//4je4W
K4Kc9hQyb0L3OOTy6lWypG8CGS3KBR5BEZzHgXOKMtbNMl4ZALyj9eRO7/o1teiv
5Z1yubwB3NxZfPMYc/fFbOMrzhjtB75dp9zYA3rum3OvwaV0eGbCcu3gjGEXNclG
Un2TaA+vP6SmJmrxHog5b8hoxadzszCmFbFernhb62umcDnm6EQsGXuqdcczZsm7
ODhOHbA2f5FkVKZjIBvlNjD31xE8yP9Rq6tT8pq4bMoE8yEsCz5t1y1uRoTMtu6Z
eUi3q8h9SM2jz9QEA/jDZ4bIy6FgO/0qb33jSwaKL4Flhw/oT6ukegr6f9+XEVWm
CGvBAP10CPnkpVPmDC6aQRcq25f72vpeK2rJiffC/6cL/1FRFaU5KbTGrJ5L/rSs
4nfFCvbENHEhnUXwVye3tOjma9K2OJUb50irkY7F3lfjTFsvkjEyIWCepDyAOXaJ
vXQp4J0dV3UO0+haVDymyMhALcNf5x91nEldyLDcSNAstC+NLGwyKWDpHAnDEfwj
XgrRDOrs6ZPsUO5YJDYapUqQnMbwId6r4X44PmvAQQ+y7UBO3BrJdwuxpEBDsC5S
33Xm65u/bsmizYfXI94bsColAjXkEjFFDMJn67Mn151AjjESbq3MU0tgQtLcOb19
O5wDI883ck2rRyhKaP2tkMzbMCz4RR9xLrz5oerhkb4CpbZ3v0pR8EJN1V3okxx5
xZAuvUZjnHTFltYH/C9eRMUiSuZ0q7N9I5ORZN9Y8ba3od46HskSoYU6W1f6/eg6
pG6KLYOWm4LFjwx8S1J6bieYLIIBraVqnNieCqR9EPHFgsC9pNJ8ylfb94sI8XrB
tmQbOIH8vPyTXj/v6Ub9A2Hda5Ba9TtxudEE6mXezP06kNDMsqbdywtuQmnpB7jk
IltlVAO16+8nYgdlTdYni4YAmdTbOa//G9CWn+0S3nwn7EXSpDiJJlaqKT+/J+Ml
0bPmrXQZpFqxPMrOrY1FzhP+EmvKp045IOwyxEOdqv9qwn0GOVTb0PS+UD+4YjN9
uXtNj5Do00uyC769fQB9YdoF4LI2cOAQ/A3x12RrXL5YIdvzfIJgLEoP4Fa76hPv
ptjifbN34ibjAWehTl9cUdGyoSgm+GcwWQN/ofimoijp36NVD4fNJNjtiTyrFtd2
Mha7D+V/Q+sSSOyQ40xn2hQp0VlxEPeJ+tJESrvUdljG7gPaGIkwFJ+IVOWhvbfQ
AjDI+pqSY2CeESxG6n01czl5QdULJSRxd7Vx2U0Q9vY93C2mlLJTjnynxeE2r/w/
1s3XaxvoAp6w24CG7f7gACPAt4vM/0KOYg/ApITs8N8KjuvqSn4cIpmVXRgSjNe4
6/S78n0qQdrrCj4DuT8CAe608/ZGasS36iyrjHbOK4uylpACT3luiiAR5KNTvz+W
JoHXRQMp4bHgT2JVvb59naNpUgQyKao/xr+XB/FAGHucnLpq9MuJcqfAEkiPaKM5
SjabGW5/CVLtgDFlXBMiUbsrzyZOZSrj5Hb+UI8axGhrZQPu4Dulq1cDjF6FT4cj
fGM8KGx2+cizuCSrqPZ3tF1Y6miZmmYKKDPAkIzx3CPTH9hh8hbCVH+XUkPpV58F
UjfbKLDmEdeIxj8hVlDNCcgOmF5AaXoREe10fibgRrwt0kC4gQOWQ3bYlHbhBWIq
08Y5fRHR/SP1b1blodIHkUQ0F2QdYMMpasnxlClSzLwMUBeDS6p1P3+NpPE5nt3X
z/ixax/5VSCMY23meJdjkYM/ISSdUbYXPLVBjXIwLvt3lxTABWuBy6EAbekScf/D
dlW5vPJDRvUliG4FoWCQe8MQuUwfcr9HxQ1yU7GXB2vkA+C4EnnsKqsSrJ9rmrrI
g5Yl99zVxBgGcRE7yjKWes2mzlcTYtUuqV53oKp3A/XYPYHPBN4EVqqOWjHEj24F
ywxLodAzBork7ArIw0XVSb/lkWO0WBz9c47mCH6uS27+S16Yk1VxRkVjTyUdwgvF
Og8JzFqTkgK5qUqKxFZZOgIbOMcec8v9x7O1s4NBgirmpknaFnA4Zwc+BQi93NoF
GObF76ZXPhUiXbPB+QbfOT0G0LfHTVYQLdxbq+YKy/H9782vj3h0C9f6gr10v6+O
5w5z/j4ga5znjmnqADLGIjPkWS1eHz8DdNZnBmk4UwYQBDLWEzW+85kSGgWAuEUy
5x86CjYSrbVqO5yXPEpUW8rBXQ7SVq7BfNZ+M4tKYXL7mwi/IqOfgOAGdjU2lN1H
R6ITGP1nsefxGwikHyXCY8v0RFbJRfMSVV+O2cKfXWoSGE8zaazootFSF51bnVY1
nahjP1a5OfDSZm67/5yEVP2eihXnLCXi75Ge7XppLzu22LHA7KxigevySyFTgknd
gaUlqvYft/uniOLjDs2aS3Txywla7J8B3U2XPrrGNeVxTiqp5d+pLAIBK/X2Mk0t
Ii9JtfdavQ4SsoOTCUYG7yzqnUzHfAXfJsek2+nOTLzGNs0uACtgu23Qxj1B+egh
ix/pomqiWWVlsH8eHQC1VY0EWR0oYN6oHRKzQXly2f1WhX/YtciyqjxSw5eKKW2b
PsnRJqrgJH6VxDgvSDMIPdNZ15mzJT8LmFNwxjBFcAskmLOBU0+QrkTRD1Cgyghj
vYRryNRNnSFNurN3sjacMjbAtFEZENKw+CHczpFtOdoxjTx5MdTluoDi1PQfQmHo
MYAfeZFXAGDp29YhXloiAA0YEj1GB1hx1o995RFvCT1rkat23c8n5uZQ5g9Qp5ni
gBNifnj376R0HZFE5DjOPfyCqvQV22IuSt0V2V7jrBtkN79DpGjEFfv0gojWbEVO
qwV/E2rXelp4YuwuuGmMl5KvkLxTqJe3ZekVjKMmn6SjUgWlHJY5fQhvc5EUEzgr
nIiaPFhlsEG6rBrwvnKn3ovu/zzpsWIN8t49FjuY9eHsOSjeKjD1tpips4ChOLJu
QbqhkLK/28S8T0TSFtIYDnylEElwIUdMpp5uyKyn3mEze0GhjsttqpvZ/00m/x1F
+AjT34H/hl/mCWKtKSkhtwn2I+vZQrU1PvqnMLfvASxXWI2TwpOONvzQp0RqL8Lu
9nrSc0guUF9OtqiC2j8tcbujUtaeBHN+sGKShf5jXyrJ9Dr4tM2bL4MBaBAymr4h
JXRmIHc1KkpbYG7QghDMxmTbsHI/DRZMpJjrOcrS54HTGiyH147X7NUii/PcKaHL
ncUTP3Tmi+gWwAcLtMlwsUKWg9Pj2IpPXH4yC1TfjiQw2frc3cG74LYrBDLdiNHH
mdHEMCTJjLq9sGNOTxDImw9WljlD7niRtNsmMW06PLgFeFZs/Az/Pl0nfuO6mq7y
u40pmGFrT1eGtJwHjBttyaZSzl9cZnShXd2Kf1R1lxYKMngwLZzHHnDK/34enVZ0
GT+ppZSszL7Gajoeugu44+OzrBDgpgxkRSyu0Etj4EuST9dq0ZmgFE8R++o8yvvd
hBycDfA42MIwnTDAvSDnH7cQpamu/z8IzEfpIF6uC48U+JdGhDy9TDJZtVTjQ+4b
w8IPuATrJBgyhyhV0zkx5/NEiE4RHgJ2J2fYKZOOBf7L9BtoshRGIkDtfva1PYs1
kcDw46um0plRWHT5ZaRqTI7k2SDc+o3PnJhwYn7PbjWWszk69UzVpSUWJ5cIh+cg
gT71UnF+CDMkt1SVG31jVy/pvriOPghQCBrEKfDweiSs5cgwd5tkPWCrnNiRqPh8
dMkV7nhSxWZwmh9GiWbpff3JAYt0wcm1pz5bruto9Pej602HTnEdJSS9wCxsMYLB
GCVasyUUZ+TXFgiwok11fpX0ILBjXKO3cySri3QX1STkTqmu/Tt9lCC+gGv+1Ltv
EJ6y7XjYUkfcCeu2dXxWhTiztUvRn3fn0WrfAEl/5holje4wJn6WumLFTPk3bspC
417Sc+0cBoAZ4AugxQwdFRtuYHiYDavzlG29ifhW7/T21AZq/frRE2zKrBiNo48/
a3APEPu06JUEqYL9wpbhPEfDqj8YaWkl/IJLDxCIm2X74Ju2DlGboNvj3jxS5F56
nX26CdmtzrC/lqrZAS2DYkFEbsQOtuW/83alIe4PWO1SXbWBkLXtr+UMc7noMO+t
BD7Ity+/5ySi1QgfTpjZcG64S5dHDDNYUOvFwmiiH2KAmsSdYQRwTvzvkbWdjL77
PEScD1/bbsWnJdMSp64KD2YhK2kv/vUGTxNxXBWpHpCMl51O+4+bK6CmJ/cfEC8b
dop1lExsmCxbQDrNd5DD7fTM0hrM/8VzuItG+OfXHFMx7pZR1aiW6r0n2UBJ5qmB
o4+rqEVUlUSchYLhBnNZfsBMp94hKGspq9Ed56AopvTFhd3yOY2ydWznrvEzquhM
UxeDYDtZhz46MaUAVAaIoYprm7X/Httot58QZRyAfc15GNxl6t5HuGvPj8TzrVj8
oC7QEe+Sah1NvXPEwEtRZMZpZ49WOSImsreljKlQr0VeH+Pw+LSF1XvTC3JxTy1s
8ctGYoix8PI+e9yvaemUWNJY0yZ5ZbX8h6SwohF6GUBqKPYaj8GZU70OJv868bUa
mQj6K2cCwmmTPmUyCLj5cS5ZFi0kyrKmhx7OpmEEMGCDmXYFVa2STh2cT3bbyDi+
G1yXmnj3cfBvoszeshaBGhMwF8ql6yi0nbVNTxSWhVl1LLDD8jNT7HtoCP4YtCGy
kIx+3M9r2WWWRPPPmKuvXvD/lUutjcbnh2je9EhczQoJsuyI80iKsHGDKsAUktJC
d31Mib8SFuzsQygnbbqAnulOb1M/saSy8ZyvMX4M0EMo7RlDSzlTqOY+vuvXSwmF
l7zwgtWUFYzEKcre6pz4VSelSwkBhLxZet6iCyQv/pnBLNLocKw4h4gNYeS2qW4Z
ckGz66+yXmDrv31ZkRqsywH9Bwmf1GkGYNHLok6gdMEjLfh7iMhUSqbG+M2wcgOW
LoBsTNs9SLEoLHjrha2F1KMCHzdXvzs5ZHu8o0pnsEpTHnQvndUKKh7+wyTYvI1j
XWuoV2fMXP43H2n1sHbHHt0gqHf7PB37Z0rS+dmyF79/FBh2UWPTQicjV/5guNkf
O0hFRoDOtZPuz77jL3Tpkk8Rdw8Nr6UIpgGN4vG/3FNNrdqPJ36JP/LBKvY2P0Lz
77EUfli5K6QIyP/5KUY41eQwajywwKvQShWnCvHoLdpIQ0qiwvoM+256Eu+xkxPL
nPha9e8b2cp8ybvhLPpFv+qMuTXoN1r2mZ5TmMo4ehevVJ0ruLihIOqkXMLxfan+
KtF7omyG13RKgn1ZCD4Yrc77A3Fnb51P5EZXvur0AfuW3GiRx3yjV3uP/EzmwoyM
Ul9kFe9j5ctSeHW/ue1mnQXSx8PYT+tCIecIYVZbSb0oMFDJS0UV4DiqkvQVwVOJ
0VvJUCTR6l8jZuKKZw7tJha7yQbwwBK4286Qmt3suLQkx3wOmdFOXqWMur+jPY/G
EPw52yysJgxgVzJE56eYdd4wzE8ihMvCIsBif9Sw1gUXdt+ofwI4V90ALt4XvQMa
Y5L9rBV0NdwjwumsHc7+rYF1K8TfDdthXuLjZ5UrF7NDpfPl6ghSThAEEZbl4X+j
y/5A0EsBbx6pFSyAk4PsJOGCRcHiKjBz77re91cMFgR6POmdkcR1dAwYAJxiV1Qu
epH34xWelUpkGkWR65h2yAEfD6U7jFzvI2EYTHf8/0UKGejCXx0cubcSfEhUZF0D
5ScgOgDVvXTLECsFWS5KO9sn5r2goM5ps0PqXQABE1wL07+br7+f1ScjA5SBnznI
Q8CJZ05bfOKY0CQwNqpoty4T3iLjCyhNPPI9jy2KYFB//9qjP+QROQEj1SeYapXO
4rntuAHPXc8ZZ/ntovPRVQY8XORZKBIZEw99ZFgxMG602rhJpeejMSuEF53ReTF8
48M+xSnyWF1jdVwvzfuzOEoVGTfo+FL2sZHV9UEJtG22CROsRNc9WDdG7Dvf0ipM
thlnyjQN2QbSsqLFhTmebU5RZ1FL5gHPNhUrpvoOFbuAmj9kl1vrnPmhAKfjS+WZ
TYkcaOe+FUm/U7NZLqpLHFeiEc+Hlvp2+s9tf5Wt+Ony9+0QdcRjzZ9T7WZLRvKS
JmjC2Z1vGxQbhRU+egX466Y3CONu4y0RhWANeKoPI1cTQq4iUmNzTFjrxOZjoYKX
FU3wAEZ+63vxV8yLHzqIJc+8prISkCyUPvHwIsuITx3EHFCOIFFeOOhRWxlDDtzj
K6n0bgl+YGbIayNaZLjGCsTnvYvz5TcwjyZs4tugpvL5DszjObkxb1cn7dULZNiy
pM4Jxeyw+INIoaQagxSnIqvyJRcV6bTSUt2YTmoqxTFAqb9NRYAkZO0shpV/7Npp
7Mu2tK6Dr2xtaDszPc0jvDjz3czqISSh0PjSPjlPGvnhecZJCo93aBAIR4p5f2KO
oneNnXLQZryyBLGXOxft1mB2xI2usI24tIr5SdHVtaweb0c9tHnHDFf0IxglOmRe
P7vmXqM8YzWvEjjWxB829azstP8BoJsSu+T4g7zWinfsStIBme+cQA4l3d4HhtVS
120NJlF3ZTavJLWSQXp8t5PF8Ylnaom3IrcmHunqwf8/7xaMUGtI8XubOOQndTOO
LhypsZYWKVijQ2pV4ayeI0xZgoFGvzXMvVyP41FyN4liV6sLQXx2KeVdjErxc49M
oSvd5taujPh2EHB8cmdwbDXkYPcCNEOSeTyJ6vFCHU2600vXsEi5nHZyQFOebapB
laSkmouc1S+Px1TwmpSKlrQi1MG9ZQ9jvnbrR6Lzfa8j4U4xFFR5MdWBbJHZYHfS
6/WL4cItrC07mvlbo72ZFOBzH9rkgYU5XpS7kZLeTDiqO360aJO/BgXRaeb5Skpn
EYpgWA93kmXpBGFN8BvqF7EDVGmazJhLQh4zMybdUrpVun1P4cV9UYfV0odpHm5c
RQgU4GY8LWlwRFdbgWIkiGMVm1u2UbtTsVX07ANtvuRDMaeRltF0KXuuq6dCoK9J
jRr1I5boaD4Vq5sZEvmxQ8EDxQ6FalD+qAqKeev8HA0zLoL3JFxYC0qUOPzWphCW
tgub/rRrBH2gvcthA7SQPrk2G8HA3CdwCENFpm7Y+4xxPcWq1C9LpiL6zInQUn2+
HOaTcHKnS6PstALEcHPB1F2PS5dt22IREPm5rNH/HurhD8PMkoaEliYBLzrMaomh
BXKRZ0l+upnEpKnoR9iXIb7Z1laJetbgUVGFVCMHiyoZvNQaGAfchNpzpuVn5tVP
RRpP1z+b2yMgCHZrUYf3mj1iJgwFlhGsPguUhBtFurRWDov1ocTPkmvmnZh7pHNa
mdZS2W2lH3dIj59p1qCRI4AbRc7le6+cLJnZZZ6JrblL+uEO/gnbLIfCkomekuza
+etvhGMALBHW1YqIYsOHVhmXEJh6qTz4dGJdo8jLarN6Y3EcgzAWB5ekKYWDNS6l
Imdfn1dZATkDiGovqpR8Y3XuNNiQmOS2pTuv74HkOJsB7tFO03jvrPvsIzFLSp7r
XY6YFQFRG2jDXCoKter9tteEfKDU/kHoYi26dpzWDXo+fisPdRvl2jwsJOriqFDd
gbuPqqobEY7V3XTA/Jg4WAklqOg9gc/xTIdGhUz43A+HE+YntgMuU3ezncfw7Jnp
YjZBHxVvSF54pcBYIViyv/G8IEfV6/8bCgbHGvqiu9pTfYERzWElil3YDlH3iSxT
cpkqKUw+0+Uq+p1tpvHA8KGEtn63ZkkLaiKM9L/j6enesEU2t78YndLh4ISnu726
9YbfssxHPt+EfVSQOY+rvKPospPWe6Cg4fgFX7CaIzgEH57rGYkhU+pMJrvrDiEC
T1cCUbgczsuSmDPtVXOmBiWJTX0ohIvyA8ovDPmHvynndFDCa6GFFn2xGzpnqGa6
5Mi6mwyrItwNZUzcdyivWNBMt8iN/KcH/BZBPLmjCsfqfeJcLggLLEALQfHKVjxE
g80+nd8ROVlcMwtl43HDmHMTBBh+/k3jlRA880tlPK2Y44gAH+temXHthqD3mlM6
aMhQ5o1epvuB9Qrnx/HVhheU5olwwUZppyEksmfKnSS5ahBS5+/syNvuj4zFBT2H
iYvVxEeyCj0fbicK/IxMVcHX4pLC84myZIkPOkosQyFWE3TGWWvTBba2lammCw8f
R2xAc1ez7p2yN0xZOUY1ULPuchqDmWejVcX3bfdDNz0IKZLx263B/1qjZchDWHkq
Lppbyu0s3yqQBA/g6SnJqLW5kZbc6X/0TFqYAqFhjWOfUNkKDHGKH5Fh0sv/4FYB
6kE5cM4WZjIKKkjYpmkJz36yXuIEXDwPy81v1QuL6PaUMkudbejOIE2O4fmJ5+Ob
hcBvoaEe53MHdv0DBAYkLE+XthYq4p2bEmTj8/LosEhJfhAA0AomGeAQGfMY4aXF
a058zn3rS7YPbWJ+j503HO2doAyv62FvZrER76fx0OjW+V4Zq91aD/R4SzlBdy3z
J73t3o8E65FLPEfaMfJfWcC06BfLRTKKShuSjsWKEuOCajSmXxnQa6XPqUaUBJsw
4EZZ07tGJApIPnjeILCeGtM+wWE11HNjUtbekfrfS5erBHiiAo7YUB+iTUGpSe46
chqMnie3C5/Gd0sA8OTuqAA3C9skS7bmHyhQ/QjJpqzQJ5mDPdXMpUzoh8QqCgxJ
YlAoU6O87WVG1mrv01vunLT7naPgQyVa9pZ/KYw94xuVnYB/woI4GdWB1iRs3+3C
CJ+mkZZx37UQBaARGP7Kjf1dzyCsIhzyPDaCn138ZhgjeoRsuFQXZ/kO8q6eifQz
qrhVpla/FXLWzGLrRh/GWPMZis4Zjyez4wb9sKXtE5WuoZ8WQhNBeTbd18x6nWwv
8gip8BcnI+TI8RqJJW+1YFTVJWK+NPZGMSlWohxLvnsTrhPOjIyCajePe4uGymSl
7scofnlNj+MA7BlgOcXmaeD7qVnVcI0hlrz//P1sPX2Zmv8XfTUJ3UOvP/V2/LnR
VLKuKDeKyv7FjPbb1oi7K0w+yEWEHKAA6e/K9YYaqi8G0cduwg5RKcKpJm1SXgpO
bHigAoTYDx671+txDG1aejSjwIGmJX1cq6Vz/Fa+nlbD1Pe1W50qCHzTubhDTx+x
hWYiKZ+2Gc7pFcYcpPe1WJL8yUU2rEqR115Sv744LgcFtbMJdg+LezdUZkVlUAL+
Vqz7P2pKsqJORMDFQrReAESR5fWoIL0zUmbxhOt8yOidnvHVEeJH1Z2Gs95pxUDS
6Tqnpj7CUAh+PTpAK/LIFSOvGGDgb9TLWRqY2PJyvY8m3SC2yO3DQIO8QhxTeC3G
6dLoIOtxzX5JiKGxHLUS1AyMTKxJAD5kKi8O+mDnJq3GCjGa/M2ffEnlfTZR/WTV
sK4ixZPOedX1FoZ6RYsh7pAn143vwADJvwOyh288mRgc/V8mye8U+bLZP0nx610z
ALQbqG490dpDYDhxTsOm9WaTy3dD/Ame5CAaH1lJyfbIW3SdiyD5k/K4YzwU7w9u
iydqUtfvejOgT/87q3ob6u3nRubVYxxB4vheY5xf5NBp7hJyglqR/FR6ekYm+Kc9
+gFSF+MtzjkdUWlXvLVR9dcqUiSiSZA1OJx/iLGwri5UHkRA2KhR/xEbXLTImv8J
C0vztuH/TzECsVHO77alqOKQTng2SQJ+LQxOVG2B3UoPg2UlaDj4WSlW9zRDd0Jm
cDF/mqc2l6WLIqF+kGMY7x/l7N4DAtrniwExpJGcpz+dlgmtbMTRVdYd59eKzN1Z
wfSes+/Eqi0+813sDbUqQ7MAy6X+G0Km0++lkQdAqPQm5czpk36v+PirehkvJleY
4PGqmV4xLFrshozydboXDCYJra0MGoQRqEPl+iQftWKhUh4tgWVnMnzZR9zRxpwh
vSmUzWIu2gq/yGf8GIcENLSqGKKPFFXUFWY0OGpTEsSNz2UtY4S1pa3B7ycm+RkA
mXT90CyXCAB+M11SOFCYDevawKdlzockkR6/xtByFLiF5x3Yg0Q1EVsfSF2gXznn
21YX7YTqyaoDVfnX9+eQKuvSiomweDtl8VCu25sdnuy6U7aQlt89pYaNwXLUMn5U
rErddhRYMPIh6SxL86UDqwrAr3lhZQLrXn/8hiDHTc7XDqld2TBtgciMry+WuH69
HJ1MQNRrvrGbyvUVxC5ryRwgqPVIw8Me4ztKbzJTpgP7Z12QsFyAN+25PM1ldkeE
Ya1pgctqYg4DKugd+czyvlyXeqHXwpYt3Toii1OSqP6ZqfWS8TZ8BzBB2Pn5wiAl
3/aQ4i8xJHYn7u+sj5SNIxPtJ8GTI7/nAtzOVfyFW0S4TEBWN4dz7G9Ev/TISRY/
5Xb8Ozfuv6gSfczDgzSUmyaDKFymcTtEQNUBNWuNLXsWNttw2fvYYJFUfHhMU7bc
V13lBkL6edXYC3rjWCUz+tYWEBNfoIetUZgbfupG9+vUnkA7mxjRUtY20uY3vHzK
edn2DpS/VJlT+Ac/RsOHjTlsUFm+/LWLTdlbW2zpDA9LY8NizoihI4hTY9WDUqez
vCWbNwlAIFrczieF85ZsSUiZYjEitugfzaOrvlWFtvAQVR7MKTJGG3lUgJjE3JSO
iJHh1Du/ckUHKiuZgv/jteYFZTdiPELSjNPwh/AM5tw7ifD2gcPu8nNXENtpVV3D
KQPjZmURlhipWKUAXswPkl/DrN7eIJiB/2B+hM3PuO+rVGV3b7J1q5z1+EXiCj1f
irswaWqRfHEVU0XpfSB04nUm6N5hgEgFMgXfPMtRyET+mvlDGwObOjH7V0JumHUs
qd39XLN3B7UFJ8SJbT6WeOcugnyQawe7zHPxzfMJpurrzrw86dO/JBFxdOoXbOGw
Np1vEyPAdw4/NzGIqxVHeZytrn2GGdIkgyWfKxsSRH4hS1dYYU10M08ZuXgE3OEM
w7GqoJhfAAUzPljM9t0Qm1lVaWHLXDFUARjp1JY3MUChKX5300cIugI3nAVuTBbg
jdU/TqolfsEJ3JGytRHURJTiW5nyQ4Bv5LeNXnCZLcYaHoGvEu+QaMy4GGz2AhJG
CpZ5LGW1UbJtE/6LY/KW3E+OEc+TthUHpoQa+lmaVmsdMuvgRXcT7qXoru+BO9aJ
NYOkKHc1gv8tJeQ8YpXTgquAyK+zFwLeVZ14AJwmk5nKhpRFXfuJ2+vihwaU8SVA
7XclUMPMwDz4VzW9jblNsBhS4XD+RcnO9fUP7YHCD0oy0Vxt0b+xeNX5eAGuoXSg
MBrbSUTFqGW9fwASXYIHqz2LnGEP8+FgxukvNAJ2+3vWW5ax7F/H/In8UO07XkXc
TA/fYrG+HBrj21wSyKcJNcUECUU46Wn0yrU1j4W+Sx8WaME2pHl6bptOKzeSqgYT
YjjWZXUu8EKYCZa8byJ9KLan4YRSfGeNAxdqNCNEtqZ+eZu7eVd2Szo7ktgZSCBW
/22Je0+hCXVyMjeSMq0+RioYj8HXIAj26oIzAE8vQHSwXI9nGzuJ3Sh6sN1aXvrr
ZpVaE9wPP/lKuDSxM6KEqFye2TDmfHBm3ng6oDHlnUaRQJKsIY+6fSzJ4es3Zy/5
jSnDxI0qamJS+ZjTGgPN2QnRwm3DkAqb2UCb0QCY79DKpYXjM20P8UNN9mrE2xbp
7xZlN20gB2nNWcFCUT2reV9pFgbNp/f769RE3jZ3t9upIDK+Bqe4e3DcgkcCJbmZ
MqUQS6DQXU/68l50mQusitFrcsDu7NnW0pmOEwZC6KiZk5r1cRPAT7Ad2GyICB2Z
biOUSpmVOPmjioJTDkzbBRqoxWesayO64dZq1YhQYLSMkfIX7MrJwVJq/jRxYTEw
+UghTmGrYJHabUvxrXXOnvjbzzzxBkrUZ8etCOO9QWko3DJkg8BfHd53tlqeqdaN
GFeEdCF8X47pJSzzgqV1lsYn001fnI4KdOtIWRGtZNP+OkBTjlqur+dNujXe5Zxb
GBY+/ASCjzE/wktNfCFILtvpCs/gcs1WjFaRyQkACLQzT5C+MNHUWwQdoQjH6inD
F9fshwCpZls3ATrs4oMOSz3cyGuHZI9h8R7orCtWGmE0WKlyynh7+uSG6o4nCgZr
cWhEr9II/8CbSRCLaJpQ1vwN5qlqtZkVbFd0q4/OuXE81E40OWQxVHd86OaYUo36
pSHN9N1P/LjgADakBv4JlfkVmOblP1syU2lDdkMsjeG5QtlAJGNLO0iNG+i6kyRz
K3Ifa7QBMxX5WKTUYhlkeHl5gE+x0aa1MI67EAsnjMZVLtdck5dcwbtqAK2u4rGo
t86fvCFLWINaOvp7JUDazvkKxCRXCkCfwGwG1vo5PuBTnlwrtrJwH8rHmILOr9W8
eWlciOv97glsO6BH911A15ey1KTZ5FQ8ky2k68BakN78eL+4nnzNNMHMQvp+5Utx
BAqCJjMoiFZMBqaipdZ7RXfZ0sIxQ6gbLwnkOqJtyUP4qzxb9jtfPS6j3xr/u2Xq
RHX/saJMov6hOJYF9shqQwPmmraBgAjcNbtgwgykSqYJu3n4v6S+WeGZgZxyLZks
FXwIu7ucd5ZPfZ0GWhAC5VNAGGWVtwBozvuw3Y7CqQtXagiY+u291B22gvwLsOUs
fl+E75HV7hbRUlC+vxyUuh6AoUEXqmXcuztTu8aDKpYDsR6zL89w1DU/8Pyxwlfb
hDK2ZT3zEAhaRGcsY5bqhJeafUzoGY1COY+SLrBigpbMiuysC0C1Y+MKaqhGxVCG
45MJ7DHs7Ht4MgWOFKiwu4/+o3ql9LYD8k5bzOjuZn9jIPllWq46eBiYDPKQ02Cm
jhoXutmPF6rT7ZXzvQMrBF0SmhWto6mM4ePt5u/gjkZYePLWP+mVpPxrTs2utjLI
ZWuga4RUlZYmQxV7XZ96kgooS8UcWXplspQqCUZPHAQ9VuPem5Hce9NZG/MNC1TP
yRoVP/e5WJ8iN6J15Du+3kq18VfyBjT3D3oHyOAif+k+D8UhDkrowiuql44otB4W
7mOqaIWqaZGs5s+DniKwEtPh6RzFuEMsQ/vQzXXzmZRsi0byLzmxqAuiUMvGCAPH
pM6sjiGCqqHI69QZcBgixxqJHvp+AU1f6AwFevL5C54TFp78bwg5j1j/1T23niDX
wYpuLRnwcOdnUg2tAMD5C/yiTGlzg3vvEQsNRvcxoVAlD3ecPVI8wCT3kYNX3pRM
sLKT5XmzjGbwkatNZR6l5uptU68Aw3Y+aucl2UZ41J2Ds9OQZsfhMIbZShCzMsNe
+fSgUrTMzwoMCEZq5YykRTYtZd2DBP2Sxc5b03nxlE8sdSxuICTXc9FN7r3Fdk3r
Ma60K1oCaYnmLiYQiN4OMmQeXMR0OkNWAixNgUrraAFDDhH/dJL7jOTN9IsgeaB1
/lA/Zh8/n9Zo5XRDYMJH/mdyfIu8hlAyKvBAOxM8XCBpmqfV116jobdsnM3azD73
57cLYR+PY/vxoCiYLbwm1/9fR3//g6P0HRWfCcowk5h9gWKV24vkYCsuty8+MVxg
f88ZcTGtfVCXfjCc8eH3UAOvMWBZ8yPZ32sYPWjolMDtNzApsfSXFwQctegXuZ+r
PMG/LandxmLQ9Ad1B80I4ufSdr3Vij/402f4Iol16m6vWP9Zv9AIX1R5HCO4i7Dv
R4eCSsSF78YwwfJvw1w10yYekGLSSfWtUEGj+IrZgAxr6ki0/M1zTuvJHypGG6Ck
N/7Fr9aFqELaRLAnJAc1GUPr0ACC+J0Qka5dH5jJ/dAFpKSLpoJoLuQLyFWOEZTH
V9XacbOWwFrWSeX65wPnt+maiFydvFXe8KZVhMobBaDxg7cvOlGa6YKNwuYH+TZ7
IZjWaYTwMxDxqp7iKBEm/SAn48iqEKd8lDjBZ9bGWLnL89q5++FcWP+6iauY8MsY
zHzKuJmU4RzBK4znRsS6LBzCpZQniJxTbhqyGoZExq5dN4H3W9zdaIC+3+qkUiUv
KW8pUo4uiwf0egv49631+7AFPoYqLmj4AbIINZZUvyUV0/WhPH0z6XJccUFqFnHg
eSMLyKbR1TK3nSsh5O81PuurNDcmDc9rkVfrdgeDrzF+EgFXeRRyMN8gV3rduKlG
n6qq5pFSd/dctN6/yv3QBHtXk2DMVZbW4UiluU6kwvmWwIVA1GMTw2/IilsmsHa1
Yr8nL5RRDsVA2+tlT2tH0PdkuSy7arWVqlPv0FCWdiWrQ2wJrYX8/C/6UsORRjAL
4ycpYK2axLB35UWl+DgCLMnySlzw31D5OH93eSRPgnZfSinu5AaQO1P634y6QWiG
Kgw/09yoN1UjyqWs/xnPyL9Z8I+B0DC0vsOoObS/egPxsj5nlWAOQNPyjtq9CT6c
HAbjaDTGhac0dexD86kfBGBAX/UleFvm3oK+UwOJ89WgjaNip5SkKbmgBLyIQKKC
ydijysQ31v6RZzgScSMG8WM1ISeIH7AonsR3almGVcCteE9DszQwRgAphTrfPmD9
ncmTIzkHZzURo8UlCWSWLastahg8QyJ31gaU9GyXlvQGXDSN805X8LVR7oi6LXmU
NaOLk7x77opnTsYOWzl2ekgmrhgwEc5daB3PapiZC+0Vs5mH0OjFWwozlCCYnF5K
mehmpDBQaAVcqz3Nne6bx1H0/93lRUSufGYa6lgPI41Th57CKNiOTdFKDI+v3/X3
S3voOVeQo+PxJR88Xcyy4Y0G4HIehuQRj5CxsptDX4O9TecfbmmfDqEjnfSGfBps
nHbe0fF1+VS2VByitR7b3RR+YzywUG2SyH3HNH2gcZlPzhmfs8lBf4zzrRhopZlf
xU4Sm6djw/rPr7/zrVcozNtkllDkYG5OKpy+fmvYhRi5nKUTUvCOP6a7B9VRZ8Kq
97XRZClIM+aLLmzCk6W+L1Vh72xP6d3WOsoSt8aWyelDa45bfc3xbPE+SWV47ac/
KSS4djiFdL8iPUNhNOfP5RPK7xL3IqyG5LI3boCWNS9T5qT0RPkMB8t0rQvLbRVQ
wX1Z2jKFDDLuo2j3wU77F5X0tUgurH24kWYXqc+wa0/pQaoHS//BV1xbbDjuZlK2
QRNekgPV1dU1B9GzGmu333ZluYjDZxkKrf2Zwn6zU84PGHiXU5dhetr2WJyX/kQu
U8xJ19VujEw6LkwwghsXJ4g3Ohqjl0DaX29TaYgaEDa73fhl65vTF/8KBzjKKsmQ
MREyWxwt83gBZ+CZOkXzf7PowLAPmcNVsYjHgXGR7zxTOwKGEIPEmaeAh6XM7p71
JFr2uGVQo8eCohseP4JkL1nwsgv2zsWT89epvCiEJ7hdda8bMU4LMaa/Ah/2k8R0
bDeGEVLrf3LdD/V/oTQo+BEW2Rks7+3vrv6yE6v1HJdKiqNnynT7mykF1OIxb+GE
3/23SEqAwZ7zXsr5fiYb+HJsMb974Y4dlAtepqu0azmldQKPbHTQo4M5ho9Uv1DH
79Y9uJKCLmpMoJnKHzujEPlFS//f3JhNTwpMZB25kjHO8uq+cCjaUcCLcoBZ5VS4
ZRCoqZzns4wOTEqtT6CqMGWR9TMwR9UQbGSNjbMajFwMuZOk+FGly+/gNCoHSmWD
aeqNXsK1SGH8C0MVniCg6BWsfrbooNfVHyS5WHAMzcE7v+blmLWzqo84F9cZYD8E
/TcwZ6MhUCF2PEpxqCRvzNcBNiBQofqId6EjuIq4FQpoiSL+BFvNrYPtRd8yjfqH
O72yumqwsvecXNKmHFlzzn3Uf2GZGL09tZK7Zt53o7aWXF3viSfr3vglLlwa9TjX
OM1ptPJiMHQZ9q3yiMQcAg9f19LdAhjb9eSOLDUqEuWAf30SS9lQRr/Ycatpgh3I
A7EOkyJUrsQ4++ITiKb65N62qZGeDOGl9AR7g/Y/GtEtrFrGevPVZ3Vah46NnLXl
sMbPl7PPxEWKhJp7842/1Fz7BItrfBbg9s8OjHgajD2b5mMxGwTv5ukco55PhHC2
C5KKpwm4oNZawtPNJWd93YL6OKXleBuosBVWjSDp2dum+xzJANTleG5b/8G5gxIE
lweULvXEAM1EG/RBS2UxKCvRoxh3G3QIkar3PbIGO1h3K3efL6O+gp0ETiD3Wos3
w8g1GlK8Z475p7rjqikfic+FRgeHVGItM23Dt7LK+OCwtF6L+lign1Ev/ZI81xQU
t9syJYB2wVRiyZU4ENmNhugL9WyzL25K15HN79wZHxfqyl22SrIPXYnc6cvcTOSC
aDiWiAToJBiErFBdKyW4duZJpUZjNEHidH98KQpj4FEHSlQkXRMruZpzBDpu6Del
pSVgHqnMUjezVRoYDjC5TrKumF/Fifv/B50AFZz+5liZCxcT6HzFy+ze9TXAqmXD
pHzQ9C3j/KNdj5FEuhnyzWL0kak5jf4URi4N5uCcY9+UCckn5N8T1k9GCODtw6vP
yl+Nn7WRHL65W56jc7lfuKhM2yXIN9lK4ldY+FeFPy71F5dGsV+lOa+X/9Xt8JKD
m6fVJJINqDNpKx4TuQGLaNJl3XlHU4jXAhjXRLTtKPOaBbZSoN+W+jt2nlG/f66T
/BwX+7jzVI4u7tC6y7hGUMS/WUOUt4P8DRN9blGObr5OGa4DCw0G+JU0y2B3v+xg
CLZDGs8AeyV39Td17ddYE5Q3M3r1BpO6N6LeZKwxeIQnCOcjVqNWaSc/IGz+g8Xp
Pi5PAIjl71lEWCaAB16ZpSxCQFysx7gJmJUJEzg+aiPQwpAl9IlpwIepaPUMD+pg
bA3I3fEfGWVDPyKQkcE4ll6Y4EbhBkYBe26lCjWEsEU7Vsfr1q97uGPlR/ZvouSx
Gw9jkGAsesiUPziqKrMfMMKtXvd4xHC0oMtt0uH078zbOLuL9MOD+ymX63kYSpdT
tbKMUtVSSttuzRmlqGQ6JWmIhJIjS8N/zrnWeGmVjRswqZccn45Xsr+lMX//06+s
N0AHRLMfPTWVa4DoVwtrMXeZLt9XHNh+wFeF25JJNfR2p3C0RObYe9aPELQEL5IJ
o2EPfl7fpjSyP+qDbopP4QHw7Rl4iids3QtLcxqA5h5IIgByH4lZg+Z/wTk6o5ox
tBcsdks2BV1pU6iiSNdGKPtXq8MbWZ+3D9zKn7uwJakJkQhHGf5Iqp58v99Uis2j
GHERQkNhQrIlJi41ElJ+LsMId0Dv4yXYAQnrMuzT5hiHKUqYuVKC5fFVItbTRcBh
SQ9Y5mEUDYcf+rcCyUv8InIA3Bt7XDsxxLwUCsG9pPS4NV7T5Fu/7VGa6toBayc9
OP6lNUSml2kbkqwkQQGHLGU3Nr0vHDmFjekFQ8LOPDuugtQ6niEktojccrIyHA17
jtU71G7lpIeuLSVWE9Z/6d6N1QqoxtFSoaMw7RMi++FMROtHOfD44000LCJD0EZI
iu7R+NgHQhRy0tBXEgBLtzfFNiSt5DVdYsan3Xh5aVanLTaWcm6fiRD+v4K50JPt
p6s+ZkIN7VuK8ogGk+I2SBTDpSYwinRgpdooy8oFM9eChY/HTd4+v5H4ObnkPodi
8GTLZMJG4Sy6R6t7Jp62qhAENXtG4/Ji8WymOf60aazJo4ro4a2yN0ThwbjtPlUx
t65x3/8n84BNoOkKOJCXBV2DI7PBrguvkgjL3RwVazG5i16V9ZySBXzmGzuHTQhh
EUZprfQ5jzi22baPiFdsYYeV/N6iWrMOTBDbPWT0GywXLM3VoDCAxDuf+mM2dfQd
/wpqCMc8bDkpp3OZ6XlFsg/0YLGNOa6TsclRaX4Z5JQWx0TqJFQvQoiH8oPvLID6
EqK8lFn6bPbsQrRdaoo2tqprgJBTOSeTnV7nN+VlpxWd4+7rtQ7KJCIrz8vXW0P8
jilU/BdfM5dR0SpW7Bsx7doEwG7vvxruBhcuFFiHa9+T0rtdC9uBNzQec+9MujiC
EOqd6rWIpP9t0g4yQJSSVLD6F/coKcN0TYgUGbw0+BC9n3TlUnzT/H01UD6pLOW/
v/S8NNw7uhBFBb2lAVmX2f8GyBtSfulgFWfaJ0jH1vupK0b6igPBU3NdgTz+UFro
8hK3APr9yUKsclZRMfUx9aEGWxBQ9zMSmoypBiHOM6Iltz1RWY5tlpTv20QAo5m/
hwDIeX8/ZIMuE607We5hu7CJVpDJTA56sen++TlXISl4Ebo/xdzqD9EUKEBAeneD
fiiaAvi9st8ubE2r8A2Zjoi8/9bTcEZG9ziDpdahIL4mwFXafQKd4xvybpLnV8tc
SA2Rlxw6Gmc0tkn++kry9mPaaNWJ2UUaNjSuEbEzjEttNFCDfzVocX6lcAwGWyW9
30R8UamQ4h/OcBSRTn0Q2S/S3PUxRlHbMO2VWHKN6YoNXxCX+z+PKO9WQuPl843H
4HSS8iI5hT3Ey3hz7/TGHtGMzqjDHyZe+tAFPRsjnjDmuLN1kN8N88g8tFcAHCCM
QUi10bzB7QndeRD8u826S+zkiU+7Zu5SidQ9ZbZVSsOZgQnHtZ6Nq1VsHhJ3X/G6
XZhBnqReHvDJ9dIoPFOhnGZCqo54ABh703X8rBo7v5CixxpIfMD01fwOW8C3uBl7
S9WOgtSW/+1/Oe76gUf0kcDKda/6LdS95CNlwrIPwDnLllN1z9MZ06+ZDr+MhlAs
p55oq4No3FUSCHZlcmyU9rgdOvaMGG1BsQ6B/gCtmHHg+0UhQPq3DHN47ykWAkqg
0xLHjyHRFzKKmSK09XCbRyQarm+rsV6s/8umGK4s6ZxZ3SKWob8ybRoItUGjfsi0
WnpRCrXm0lEQHgDT8yhjugaxVXEiNGugmSnI/srQZnhaec29yiav0iaGEj2tIxme
x2jiSN/Es6fJ36cm+fNIQPDKFIyqXz2dn3EMs4SgLG7xeiBeU8iZONNDpgSIIHiy
sIcMJt7zzWHN4553pH+BIY7ksoaZVVW5V/5Ww6oNgTDbr9Amtn0m8jjrkFXwoj+W
oZsjI7eDbCv1piBvedsKhdJ8LyrwOfSrVeQzpJWNowv1ZYV+RbfH0DxfSuKWQx15
TlkHv8V/DIEAKaJlkqXagy/LPpSjPoQCHmKSRMGBlF8mENRQsQZ9vAI/zhrqP3Qg
LmZ533zxkqi/inZzN+/gpq3T/c0aBGAERHpCnfRmMY4vnMTa1nfOIaZO5RFpz8Fz
AiSzxxuE3B4D4BxYAMYDtsEZirG6ieTQCkYJVmACPlMJ1HMYyzo9N9ASmrZ4dq/z
umkU66HNtm2bgC7J1LEQLJrA4hiaJykcI6J5pk9+2igr82jKXnQwuDi6vRlcoiLY
vN4EddKEkn9tnwRSzHtRhMUJMFor3YvUcz7nVlNNm4sLywlvL5KdCXrCv5bPYPxC
lmFyHA/2dko8UuTIK0RRFk5gHrCyylGeKlQ1bdfJdFBzLUNvQqCIFP47hWuXXBsu
HoNEZ8CwyRRmZGA3YokP3k7m7jFVcuDvY1oOPo5a5ClBDZtunbsLKJN+f029n0VG
wBQTzz/OdoELG213YZHTxIBlmspMhN9oDHdoTuoawNF4fD/LOwGZSsbWuGYKKXVf
dnIFt3nKHi3kJL+jeAepF4KLIrY/MWWyHJwKSAtxwRSMPogmExdQ59a6+DfJsGwA
9Jv9dMiRZ7uBuQzZKldFB87DX8wvKdE4+hNsmAnfbgl4StCIQXosETcemAqvf9hE
D2C0MNVAYlaoR8DMTAh9o6KUZp2yYw9jIky3AZUczrzAE4o5IwTQBqJi1aXtVM6m
WzmoNJnUPI9fF+ZiG9PQehZEkDyFaN5GjIyzRe2y4nOvZJJUjxJwSUY9OJyTxjFI
J8Hl77cvhPkQn/Adk4rI+Q/dgI7nvb6WnsEUxhXlYRlOf9joIBIZYeEwdgFjKba/
J2glSSek2yiEdecSfT/5QTCLKiyicMdEe4icM8Q934pGGNFD8nt3aSZp0RcSe3fa
sR/0TbkJu9IS7BO71PRHbpWSqbvwXxuC/kOV4gOnxg6nR5wkveWGX7HtfEYfuiLv
WUNeOlDOKnyA61Bpn3jEM7PIasWU54a350n7+XtqBx6mbuXAGIF8kBocFbGyN6zL
CHYk6Ayh4/womBChqPvJ88gVhRPklYQupQskbZEb+HCskkpKs/orhD+ldm8Rrhy0
1IxE6/+edKIxua9QDXHC5miTmKRfYjdhqZ135M3IGT/VEqA94yY5FNPpe8AsPleD
o1gwVlXJbB2AX9Wow6VLN72at90C59ghsxQoyLSAyNBDyyU0NTr3S2GD9V4FjRqh
74BT6yU45TlkbzHCkS59eWkw2Dn+MsQG3D7IbdrF0mGNy2LWZ9cR2vUFegf4Ypso
fVAKV0ShPb/Z8yOWE7ZHIPMra/Rv0DyPRMfydHpmi/D62qUWHZ7B36+7bqNhGbkV
lAVpeFmt/wJOtUIkUzff3s1Rrhr+UoKwPTtgPqMzle9Kze+S/ibfILAF0fbQj33f
2TH5CFn+1/viMWRXDHKJT88AI8HATKcyL7632GrCd34+akxuyZ/EAlDHQODLp0lO
5A+vNfayP9X4GvewL5wtRJLIZS/+/mpRMbtV7YC1m7iwJONY5q2edlOLsPF7vV2W
REoy9ft/zcO6w+vMjx/3zhBV1f4lgmZGD9L+bMDQ4BU+iSE2pjwQnVuRkcRODHcJ
rLF2vqOfYDZURLsAOxh9qWxQ7fgJwdGDyqF/iSozQFHp3RE3FIIoi6iH/dtfzGrB
+DDrLfyUselePGJgRHSu72Het9nbWrFqfRpycMAmPlXdCu0h1BXQBXuCN3hrfAqO
gMSMxyLZAEvHdRwCFbtd2PxCkV3Q6K5m4Q7pzgMoDg9s5YK7DBkyxE7uogYbXF1N
S2PyMJPWCp/TWE0KQu4GreKkPOPMiSy8C/8fatYLdflAx0Gs5zTaS42RaSK3Nrak
s8P43EaPoAFttl/VGH1kBMpY40r9BMYETb/sgRu23ha1XXh/+B7PtCPEJhrjCq7I
AwP6VFQk+7XL58yreAWQ6rdnxCEFosfc2Lngl8aA5dnnzFwxXnrNe7vhAgsUiuri
UeoitJVL6o8B2hHTnlNEI+KNOEA6Ze+NQX3XSC6FYoui1c/sKx1YFjz+O0wVw/YO
QPHkXY+UrNuTbuIlTvHo7yXrh97A/YDoY5UeDMa/tT1/tDFN8X17lpXOXrMyoxGi
MpZKdP6ErosZWxC9/FaZi0W1s+G/M2jmjJCX+XtJM2arGnVTzdTYPhkuYbCrDvS+
R2cA+ukU6mu95SRlo9e40bcg2yD6qL5Xel6Y+7B58/79ZMe+iR9n9FZDFtAzMr+d
Z5zEI6hTGP55ROevWAQzZKlV1Fhqcs1DR5/WEImIXgjvJjjOM4qf6/s1ecVpvmWG
VLPrhdbVmcf45buWP9U7oQXNHDZLcA49KTq2JyS8DkeJ6X+PzGUMrGyoekQ/McKR
3910VMjBl5wvE4PyGljs1H5QyzfMDKmj5tVbBEpHZfh8KlfkLTG9eFt2DRYA548P
0+LvkyIrtWhX4dFNm+f+GmL2qU40L1nta7Kxx7J+SLeJgpZD9lsVYwwNmDtvbJwR
GBKFHVpu5cTgPGCEeREiDIZ3Z5Nne8aTp7+uoHWCzoEEew8788tiG+0VQYgsMzej
CdApjAYSqBuBVAFaEM+nLYZWjLeNcawe+Nb10sHWcRZkDni4fW1qMak7/s8P93I5
LjhDdgWEpK8F2xM8sr9MDJNqh7/dhyKEOgd6wRhXAqBnrhc5Alfk5T03EWbFX+F8
GWbmIFyXlggELU7zw5TBD7iK+bbucCTuEOX/hG7hoL3xDplzVnnLH39s1k2YRorR
b8JTZ8rj6OZnmq/K9mL64UUjYOp0P0VUs+o6HiAK/LQP6O02n+5+uwqzVC71o+9O
p3ep5NEBGTlGZFny4BurSthOEooVRfRk37Pl9KOXSw4pD5hEsf3ioLwHy4vSySnM
H81c+KF93R2060C8G4vZ8SQupVFnJXDz1pwVbzmdTiG1Y7Cy+z1AkqCcZrofyZ0Q
hEwtpydhhC6FK9Se4O9NFxVQ0b1jBp2l+psQoIOx7Ktv7FIQexwy6UO4Jy6Yn63+
LK+KdloeXRFd/PR38/eVx8Z5Vbn5l+IAgNEdNc7xDYXv7lsgIi30w3QeOmn+prVf
S56s9BaIT0TNaCV2ys3feMEErXWUiieMjndePWbUqGouDEGQBOQEBSU7JdnGFReM
38XMETJrasS5e73yb1BAEX+HdNvs3rIIIug0lFWnh6M0Ja1ZqvpKbK+H9oDDGpb9
VjGb8oVVx5t/8nXNKQt+CgnExuENRLy3cU8em05rK7R2FGR07d9Ke8xpX6gonJKP
VkCHN/uRjhc0QciXsZs+qwpTQ/Z4gB1WLwBsg208kooONq4EyCqtQzJiD7oaE1XQ
WHIjmztxvnFxpiFjOlvNot7F354I7qnGhifcKyyXUc5R6yLGe2IQo8bMqI9kXwKT
L15Tt+JWrhqeajmc50hstWN1CCyaBwLv4Awr4BwJptEEbvfqGBYREnyGuTMhHsJH
skN0gu8tOx5AQlGuEkw0cUGADNfT4x+wijtiAFcsj3GjDq0ZY7r8BH1xetf3kk2J
GL5d5MkqM0kmuA9jLOgtlEnWncWXGqs5iKYzUywlc7FemTxI9jPpkUNWDKK08ie+
SG/LJTeVtTZiP9hdJyVK32OaZYuwi7wLaeqSQm0P/VDpHZp4eGpPvQbEBriXzV7g
kLKWcPxR714St3Nd3zof2G5Q5T6OGHZe+nZvBXq3Z4uhxSjYWJquqdg8PAksNPBi
MdojGAJKLa3PvChYqFYSPH1/rqqqZrolHGnNs2IXPjvj2aFVeETdXen21hiYSsQ3
/4FqhlU+lvqdFg/4oc9XWTpRzsTMXTZjI4YWJUfL88FO1Bc0Fh8fjZhZQfMJ9Sdm
S0RG4t9HTU13SFeNYr6Oo3xnnehPdG5X7HAWpsQT4X6SmOkZTcA0lV5IHWhJdh6f
FmMCKu5yxMHXwpFSYyl+bIPuLJ7MS38Upy/OOHLl8cIPlHpljdkgrCQdyQL7Wrdm
FosvdQkPQZwK4fo/VInbbZXG5qUGtkqXQ1FLtM6WfkodsP5xP3Lab6JsXPtdjfZP
JZG54AX9H6VQ8ftn23cqYAhxXKiZtrqluA4ISMPhS57bp7kPH2affVAIqmkKzC2G
NpptuwEGsxQZ7+lIrPha2YF6ckodgHyxt78BjIULCXR5qgYHcj/z+sb9NEueSzWF
sq6+4vuPqDJT+LnQuTusKlteR5WRXMLemnR+d8sgWxMeODeJRj71dbwEWVvjQJ2f
b3xkGyvDvxed8iCAW1Gi9ARCzBTj/0wtVLy19PMPmVHxgOTH6QLgfHhkaNaz7vQ0
R5CSfOpMd8pLVU6s+YVkVZ44Xl4k+CrJ6hWRfK42Qv1u8ReQD/OU1/LX6I7rg+by
xki5aBWWBZiM7T7C9czUcoTFBU3yS6hzDxA2lJpa8hRU56HxY9+3VvlPx3EeKqvD
QWloy3Dlp8vqbZ2XeDc2djLhso1oNvaSjqQR3WPo+Hjo8OZzRnEZV1HzH3kJ0tnJ
jAuq4hfyqdRxU8HiC/7OSXshaXxkjYOuDWcU2hkr2rzgc8vWxMSNkSLR5xC2LJP6
BimGVb2/XxDEaNwxByZlYgesmP7LQXgE2LpWohFDHi/z4bRLbgTkSGWUR3WychGm
UntaRXiXPcfazBk8TCD9GUixroBFD1eDZKQaVH59Of7N/U5/xw5Jxs/5VqJbFgcr
2cMUkkjlmqRW/S4Z00WsQ4nIunkDJY+YKG0bs5hoSPEpIfQkFoyZ0kPQiXKaU6fR
sf27S0wgItjfM9sZ0ocGcxQFrMu4Er0EwYzqmETCwsTz58II8qa0welzymeAY2up
sGhciatibwDebJAk2G8WA0gOiCsAUVmNb6jUTPaswK/E8/FmidSeVGMardhfrMSC
oRa3mhH8JBnTfNQ4+1Tid5tdU5VmET/VVJWPLC0SVuxdDXkexwOKbWCGJtmAUFoy
h8h83SQkCmNMEAHlc6J4xQJ054rlON0eIyt8JKYKQsSuxVQOopxMyKlqubnj67SX
UHSzC9q/+3pQZbQuSmAK5H+dA0C9we+jy43jRysgVYV1TbSYbJdDrWCl2wyrKfZu
LdFgLpu7eGcF3vmiie6a82KNlIV7jOHLmLH3/QGMyCNRg+TrtnPyrvLzK+Xv+a8X
cgJFyT4cyFr12cxCEwsAF7da66SkjhfabvhsV02CG3ym2GA3y0NAPxvcaoXO/qNH
Or6tMhm6yxgLMACPtM0RgsO95t2GvLR8d3F8BE8RxeEYrn30V18zoHX9tVeVDb2o
lCRSlTJf2B+HiQ3vwf+y9GB5Ezf2ZyF7K9mGJN52uYBkCmkk6D9urQqKkRNKgkPW
dMLAtycwL5wj+tWxC805KFd5WYnARbQgwKm5eZV26LNB8yBISm9MlS3gkr7nZpO+
sHStzxuzZw5yNtPSMlfn6mQq39NZzjAWz0EWzUvWISunUtiEluCRNLeGG1oATKdN
FKfn3YuU6vTVXd9M7/N9yHvyuJp9JrmIKKRHAo5cQKvxYcpsmXeyv3VpKPffEcxz
Huz+4Fl6CYJ/HVyAkHisLorC7tBC87a5m8ivVETl1GNoK1p1VyQVC9tIuRNljG8F
sW5uxUAOKiQSgqno4SKU8cFCvk8cznRjNGCmeT2DlbgoVyGCye4E8Dx4CNrDMcaP
CVIaeVFClprHHg2h67663csKvOHQSTuNQvBxk2AQFliR3nNpGIV1GOfEDts46WqP
TwVDWTO67Gw6q2zfLk1FmkZDE0HjWCiAjc2gNSO0FwXBZMDa41jbh5eN5F5Ft+Gv
m/P+avCwvOJIIazEGopseSGjmUQBEpSdti1NmFVfuPwYQcvdsizqZO5F0NB6VavR
tn6NgHzgnFh32jEyUZFtJ13SyH8rJIKhupdVra7LUAnhH7lonVGBvAQNt7evBmDs
/SfOnj07l93ROr2MdPWDiqRPs6Yy0XtAkB301wC5A8KU8w3Usm/4WlIMT9b/SXYz
5ewYp4bsLq8q7qpQOpnwRzVZ9uBtPgmA1Cl3rSPf83nXivH6Z145QwFqOev0lQKT
c6axaOm0IdxbLv/oHB48UlVl5BwqOrdqOL2a7QpGUvRsfGgaADC7eepy7eqCtq9R
rhQO/YTVXvJ0dhYV7sGnLume3KqakIDCdxK04/VUQC+t3+I1DCQI7bfn7DOFJsNN
ah+in15kTdC1VhIwyfVWtsgVroJZWK2vEEnwFis6LG99wt9VtolIKcKdknvS+nXY
3hn2JIt2h+gjdVMYwhOfEzZcsd1Yr9RPPVUCJT4NMduBBPlKgsJqK0f+vE4MRpxS
K4Zhba2KTahASfxY1O9Rl1V3UIPuxn5eKYCBNiY74VPtvu6uEWyerLeje5AQhnjR
cM/zfZOxP4Ao3AC6ic0rS2iigdTN2TOAmdcrquWRYvTjt+NNavP8ib9gfZRq8EGL
lKPZpaqmeiB8d2h6zDLQq3laDrzNCt0JvqMhNm0qtPxrXQTll4p2BC+GVhJoyizR
irjaQNyQvB7+HHdmjGMUdECOvgfN7omC77qxnPhDNjswZkkf9EWQ+od4rDe16de2
sRz5vuZuPcMPuJsulVmMW2/OYMpdQaVkS6BjznnfcMCM6vPuZH5fg+JiW1QZtuA3
yJgJQWrDHdBSRZFWOAn33TYgqMR2ayHNQCOmnHhtR1WKUuLWtqBPzlvo2RZG+HCQ
tCKSPmnkS2zBsYL2kD8mgDRRga5lY09qU1y0no72Qw9mnRURsUlCiHx1fP2BCAmD
Qa+l+H05syTmSA4gl9FkOidORsLmtvizymnPnckLldVrotS1/H7P3Az0xX1MwjUI
6tAr7XOdlqL3GxoEgb3uQsX9oxecVpnQGlPrWkpX3Su0Xd1o4bFXv8Oxobpt+bbF
cxUnraNJb78/J1rq24S6XEf8I702UST5cPL3Vvhwqv2Vj4NEjHsvuGcW2tPJBo93
VRexZmA2LNFLL8+zbIC+yU1FpwSS7K0WggAIQGVaknoMBtMJFtU5n9NcjG7zl9N3
Gn2yATJcUbM/WOf1YmuDW1dyd0E5dGekaapORE8P5U+Pg08Lcpnxvd04yksLjVLP
+20fJrpdYPfEOhOC6DoWWSCSJb9jHSv4VnQbDWxY8YFm3WqxRr2iufIbfy7dLhKX
fdq5oLGGy5VceNK30YQlteVSBtVyA3Bz79JLYm/DvDRpCxTixnB16SpqqsaKsJp7
EiVNZv1vpY+9i1VE7/24KaoPJ2/Kpt/nJVwZ+LsGBYxVhADZskj+OuWY2pmS19xK
ZKOnhdPFH+UZjgtCJFy3XLHs9RKX016rHuaoCUxW/k0i8eVKB2PRKfNxlZ0Mmb7O
5W1Y+0sjewOidOJuFlNSggi1QwOUcdUbzNgiv1lPYJ5+cxok/1PA9miB0ZcY0gUz
mSmQBkv2s4qm+F2bJfOuFr/yUF83g/YYsPfNoiIw6Q5MpPWExP6+EBmb7Kyb7ABZ
XkCkSW/RvK9g3HYSQych3znwKy2/PMWLXqXV7roDyfYoIDvjcr0lwYt5+L444dLG
As360STtn1k4Jy0j0kntWO64gbe28o8+c1GgNKysme1Gghp7mmusqRkhrj6zBIHj
Y1llPjAENjidG67pCYOLwvipewvjQl4ZDJg8ofidHEAbL7wFScUeXJYtziPj55UY
B73oLu4v9qYRQVMfrNhGHevT0RKqkoOGw40h11xCTDunFigwcd9YAsNjSrRLaXUp
gqYibF4KzwSbh3z8hsnRXPeJTVnghdCcaiYjSAYRB0n/bNfbeisr8KyFvXVtKry9
iQ/9ObfrwHKPsPBLagBCfLkGhwYGQTUDrpLtxomznA2N/1o1y7555yCXVknzmXVl
mKhLurg7XNTTCYbzdlC9sEvIYI/6/nfnwNxCoEVJIFfJRq88iH+4CP9WsnXDpnuj
Xe4SA7aDm8BFLWUeqKNxZBXaRiHfIroMgADIWoumwAOuUkmgHtjgOTq7aXI/DS6e
cOedaONeCwhXgsiwLVxUaM63CZPHBKR3b2yG3CHsJVfJ83oFrreI6O9oYExEEa9z
zkmJkJ6VI9FWA7NEhhxA8yun/Ng0KrBsiY4dwsIHxvgPwpwOUBeGZ0yxooEgx+wd
hjlsQV9YBFNL3oLnj0/yjVoDSS5iKjuOFEXfAUFmo1WX+cxoEdBdpj9mGaemeYoR
jGuQkKvmekS2CPzdx441LFoBs5HFPU9wwwCY9n+WU1GPtvIf/1ReQwGeei1zYK1U
Ewp7AnsiiNzv96U/aRkWJllwX0f3L8y2YacsLjcPeqM/7S/DRdt2zBCyP6RM1tll
iOvN+uWt/nkR09uMXOd6je5zPnlI7yFbO2Y7I14NElac4j/FpEC2lEEDWQIT8VLu
Ld+bUK8SAHbtqcH7jZnxW13UAJqQSszAwzje9V4IV/05gXfQtVhQWigK1yErhVtA
YxkbXKj4K5w+DQIzb4Q1wUyhNzIwzr5ClI0jKUFJgu8EFU0u3cBPoG60uEZ1hAx5
qHSwbEccMLOQL7UwUJTnv5fpcnwYeJH/3kNrcmIX65WgMZIJg8aUYeOhVUeXgjJB
inFhU1nlFh25vuiT94OOJOMzZgRXnWxbN2vYAspaUb9NgIyX/wQasluENfBnyEYl
E7QqdUiibr1h5dncx4rHt9iwA8Pvz3SiiGrsbPZ0T/f3rsvOsHGjfpK7gtC7M6Kl
nT5p7+oHubzctWBE/HvSZTuFY+oWkygJ3B5eYsGERypzIZcJMKKEwXE8yn9i92D7
MePxHfm/+KQ1JfmVelf5b9ViCW2pwrDLSEyvCUA7Zvjq3BaUaoaDm4aIeSRRfpOl
HbkoXamtZrYI5JbrcpIkR5CTaXnPlCPQaONo41+RCGsdzIEM0VWBMzU6NAR01e6i
v5Ij5WbkdSCrX9RE1FtAVDKSntWR3VxoPVQZtCBJ1vXL0PV7eIRfFnzdmAHxO32M
7aTSxiuogujWWWv36/qFh9R/uVxRXRQudyiAuWMQkjHlhD80kXXuW2s7VGDiZ6hf
QNQjzwteKodB0AMCoaarkoYx/b7I45Ak29m8gneZFeaKfAGku49ZgEEHZAMf7oIf
3YThDOrUBDSX94qmD7PkRCuBtLLSBps4+fS+RQ57WtE/6kdXgd7JQ0jwc0ijnt2g
iodAImMSaFUUgLhhGRnP9wEVYNxijotiyAYeTzVjFWeWPQXlhdyxWRXszvcI0uwD
sBAJiXD/gpEh0QWHHT2P8H8F6RDs/bxRHANshddBpH8CKZJiXWopK3/ae8GyjyIM
TVWffFp97VkfK8735brgog+M0aC2wH9Ckso+rTp7yrlOz+FIoV8zldvCquYgvIZQ
nAtLD0cpfnwf6038KR3zdRxRQLL57zEIFn9SlKF+/UGZaqDH8EN02tMtDNa/CGze
d2NViw9Nkavp3jXPO6454+UZMlKeGXc71v2jichqFFUsjiqXRF1+xbHRNBcoVVDZ
/7mMSYCTpwMwcr+yYdQOt9OyXqNYbhTeN0f2pTrt0gM4+GELf3tU84AMLREajCPh
H7ujWjPpw80hmJfKreighI/GRypQgT/49yzqNbk/xfyGzcACxeHHUr3LXP7ZOR6+
YZiP/nIEWA1gaaspbgqNTD/lprNWg6nGfIA4F9vQoPsXWcXHuVFYUkL2pebdYDM+
wz9Ss67Xj89+XAdAU4Bj0Y67rIz+o3iaS4Uf+bH6aMUzRIg9oHLMG83OJhtN6gNW
U9rYTT4FuMlrhRz6CIKzl6DJ2Sw92/roLRgywNPRaup73F+iPoUDvV3ZBFsRpXfx
2HEAGjwtyz/B7OOJNgIP/1J2groyc3nVT0GSy78X938U7vF8/G/DOus+V4Oq8ew0
W58mMtJsndeVY6la5T1g466ttVEiKEtMBPKxx0qKjjHnujL76cojiKYsPUnAlaK9
Kf7voL1XvsysD6INw1yAf0JXO1BXqnCUPh5MNPI1vRnL3V+Oa+90ZiueIqFYY1D7
hggFI6cCEzZjbCp0bTKAJLn6eleSNTyJ4iHFDoaKbIfRbuM2q8HygPqbZJSq/d+n
vdIyYMz7Q4AOiYpf753kO7z0I7FmSZeKWmz+j+h8JamTJfQtm6PVJ+rH22HUwzFv
5mtXWCQY0g39Gg9jJ8SCxvmujM0q9wQqHQ01VgYx1O/nYiQeWP+huhee9aIfoleL
5Y0Rvc1jMjGgEOaChoPsT3x/dEsN7Y/WSzTnB8zJ00yyAA2LhTRWdjVgZNgf3kKq
bgqd68nlwh2s8nVF6K6rwzjLncm0+04pfsptXOwv/OQ1cEKVXloy5mNjyKjFAuz8
LbZt/qEMgZavxBnPnHqHQ3MxmOta95Az6pqt7W7DvhWbXdNn9c7kfcSrhYxJ/7zd
IHsiQozHVo5FY4pHA1RNFXARxPSHGOiUarzeFKGUvwtdEQBfefzA6orOuIdtumz5
iZjZNq7SENbFORhBWpGh0S+ssuggg/HNnfT/dxWsI0HtBIYuv5aDSYHlAxoalCNO
7C2wtA21x0jVV5bNN/OGBZwvTstobVQYtregu5o6w3g3Fncqkc2UxbHJ4fajom1v
tjOT4nNgmqbKVmPyp6u+OeOemHyhjyQP3g+Eq9/8zAND3VTQz30hK7EwdEtes2Rl
mG8GlUg6DbFyENIOP67StJsFyPX7cTIQKHflPoIYSpyv9z4JWwMVrbA7nXH3t8nD
EMWrfSoJDDb9HWd96yqoX5mXUMpvzhNoet4GbTViOAecInmiJFYx6xx0wYStNcq0
tQdCjWtmTB84j8RpEVLLNXmSrMfm0yNQR0rsI2XF/S9M6ea6Mwat/mEQJ0PsR2it
f13Q1r2CKy9ki6lrwqG1QA8kOuY5SF0m0An3uhz+aqOH5MtiWnpbIrn3zXL9ITvR
xcC3SHrDcoCnRpXFl+zKYL0eFcXe++jnoq/Ni6AvDJr1AlCIKhrwOCZt3wetxziU
8/YjZB9GpG87Pl1KSB0M0A36FfpiMh7Ppk2c8+51Xi/BN102HWYJwxho/9Ud9GPs
ReTx+ZE47XbNDMVgvzT1pVVPy7nRORQ9NJbwMwgxgsAXFD63w34WyJqW/r4aEAcc
p8/A5XR874D2stnxCbBE+cjt9Z+QCESZmXhPzMhV+HkztRMpaQFzacLEamYN9CnJ
7bhluXyXb0isWP234j19g4HbpqXF/B6T3ExGJWffg5WCRsvjFkQMgkMjLSpNWE/3
lrXVeoPsj0Nd3iLHV3/ByPfHx06kJLDGhyoovNqH5jkGJnoZCTA0o3eWypRjRV7W
u7ahbYQP4K+Re8J0M9FnKyxf9SE05+1FexepOlSVOe2hEXyGvsF4hLup/naQHY8+
QdnyrTZRk0n25W2lfnIm71I56o3ro0RV2UICny6/EImdCzA1UUl6MxXBYVURv8/M
HSgocy9qXkHhlq5AHKtFXcCFJrsGzDimsILH8A93EFvUyw6mB+V27pq8kd1mUDS9
hEvbstkuJzKJCSu58F30UaN0/SgsucDO97dHPMfavydCC3vvX4e08O35h8eMEKxm
v2ovSFs5ih1QX5ixUbnmbJS0DejyzSoANvmVDOwcdZEsTdPQrWCk0aWxqaDBkiOE
8ZWPXe3Ruxx+MCAxhwIBmQ/Oe7Cy0y7/6GOBdJ/6r+SsNpQmXsNjrcDtsZXEmJOI
xTcqE7jAflixXxrldlkTbfd4amRZT/BZE/aVVM6iiUkeSyJXssu1AJkRviwI3l6H
EZmbx7Pu2mlSt+XRUzEbxtZl7ckyeKiwljhXNcL7tDmmAlO/cK5lkyHfwiHiAHw7
p9mBKlJ4cEQl6pQM+8IuXgaobjZjeg6VVBSuR9n9nlQefvq2hgpsCb1M4QKUkk1J
Jhyof/3nS33U9uK1A1ONszlRy489wmZUYiCeteRR+S6AC5qO2bzLZ4y34CFbTV/W
YVs4wGi/VyT+DN3IpDDpIdIB0XNB6bkyOl2lw2iSthYC3r2esgMFsMqjmxDvFqAK
9hB1kcsRZ4lbkVx5UyXpKoRF+pLEy4AesgK3xP9fa5WWZm/Jbmb1qnW3h3ZaX0RS
yqiNU2s1GHPq0Ll7u8ccqxDfO/9gZIClTaNpRjpv1SxbtJga0UhCLBJD3nmRKc6F
a2OV7OKYRsdkCdXCUi4KXCltO1+N9Ipi1ltdFya+8eFojqQe7MovS2SbCR9QW+4a
cRwUo/xiggYEIze3tuLew9wQFNT0BJeIogh+b1XqkPP4FGuNc3gSr4ruo30FWWgd
54r3ItfU77npKaoXoBMHOVL2ZulCHLq5t3gEb1APB8UjejKU/jJyZVLrD584nNvx
Au5tBNIknCh3CMysYVjPNEvEFoY5YI3cqoA9zVM78S7vN89Kf9wcEd/lr0D4SFY/
UD6bthaf9bwXFxlxfdk+BtRc9jpeeH6nVD5YhhfKO5em1d7wyh80d+/PTKJgHh1h
11jFtyxPFRV8E/4QQzzk2YBiqsJ6JuGoQ9lZKSVQo/jMXqoYbltyhv38n55j9SHP
ytIKJH9iK+9CiKSQq5EIx85l0ZRmBQIK/JOTS73BtYCcao06Au/K2HynepP/x+MF
z8NXQEEWCUkJ5feFsQ4s+YA2IwluNL0QXsOP6wX8yCiEntugTuTFZeSlgE8Ec/4J
c1/iqNBfbSPnq1bAwGPHQ4zHEHh2Z6RgpnUOXWcJJRomH0scIY8XVBQvcwKl6rqw
PZoIH+adMTZzhVeRE7wkd2uzy+gSWD86KYL54GzGOvfZkQQj/3nvSpl7VqAwoiC7
Ad8Rn8kPD55iAM0khbLxNLPOWkJ86feajr0NxSjmvHqp5WpEiFbNArdFi9Lg/5Qr
s/I1w8isVb5yOte+vSH+mwx9uZ3/ty+uXoXcmGRlCj6JFnBcyiSHpyjDEBQFAeNT
LekSFFMhDfyR/QIOCO7R3rq6OjmJlz0OBqCYy3NAbQElQx2pEhiDz7xEphFIsh4s
TUu30Q70E7h4ZG1SmcWsk6BE7nahmxOUEKj9Uxs4j1Y4h80iCn47SEEi90goEYXB
eZZe+nAFwEfXD9lCxutWqfsQ2G2gR4dLFx0xp4OikcoM8XlOu/hta9sXcSQI7RY7
3gJIH2vSfxjhYK3m/1sTF1DcWHxC3UhhpYTMoWwg+dwHqKcRv2RqlOgLAKVrR8AQ
X7fjwlQtw+DDcjXhxlRRJhisJK2gTY6BrmzCFz/ijR5BX5GmB7UHa2pvS3KD5qpo
70k5iiIhl61fB69hMj/cPCfHR7x+WPXsUk3hhcPESGc2JZEELGgkMp94w+KDlLSl
hCpV7XVJ5ybyXIKtI08TQy8vCWdRFNdMpKsYJdpo4DXGenMrxnIOi4/HK7Ym73Mn
Gc2OdR1GC+zqLLb7/3J+uH0SbdI1n7/Rl3OczInvCTdWznMfXRlPARsZKslMH+BO
YsmwvKml5tm3lzaIrvy3Rm9mVOI9taKBMNF4axzCXJIBqKVYMSqDtSP/hcwH/dhJ
aoZ/O54XAHBYyRBnZYzn5xipBr00X/ok0GkmRbdub2rF08WkRpm1P6JQ7BK/4mLz
srEOa+5l8bTk/JJ+4on3HuvWXZDBBZKKsBTZOGgGeqLfnvkZ9DS3/M6j8vNmYvew
7MUf5qcOf42PnmFEGZDx67iSgJ2oCHvB/WT5/G9K/RawUsiXD+43s8B8nsfeW0rW
GwNG3H+olRUvKE9PpvI+I3uQe/UQYt3ufGjmNlSS6M3+f9/E3AWmv3kBGl08M6NI
gfZXK4SjId5ALLXXFs7WHprMtMZgbXgbTd9ADSfmp08qIHFkAdqfqm6wfMx9wIMy
46OHwEVnvjVDHxoGFcdPnRN2uf+6nD5Ue2dicxcZ3jfdetSbc2TuCTZmHBvingEH
tZN2bfAV4GxAfnjtEaKUj/5GBEF8cc2ps9Ri4JIBPpoBO+kX+hqxs4nhej0KBwTE
NgLrRH70EXdZR0JF/oBd7KMkJXtGcrm+t3LthIH6yjFEMjqu5YK0zn1T8mDRb630
21c7MnN2hktkED1i4Ii872vWMm8NV5zWBQwjQaQeHlU2ZRrR4rwUBRrS/GS5VgdN
ojv4FyjDDuCUWecdu1YbqVqhXg0LjoIooHYqET89YhgY6t2WURUbRfp7uK9bb54K
CGs1pCjtPAEYjw431Pa7BXlb/NreCL9/XCz+2RdvsMOcDNfDqQJppaMFS01Dhqwg
DUl1qkTziJ+tO7jra9fnaNyAmvjVweHOULg4rotuiXjloE4TaQWx2BleTQ1RE8UZ
ee62my6ny+wm5ZGiHj8Kcag2M8k8OEER5QiomKKnzpkjgPQq5weAseuZ3wci5T/u
qMMSNZHB+TmQk+WTNVJXKjt+tqNKCGEEVUNdcX5SbOn5ipSnuQMPY5F2JsJ03SEb
Olxz2Nnx0KEQjRF6hslEo5HYMy9pyhCkhG1UDEm9asY4jIpzb/brwuMzicfXBLwZ
ub2u+uoWllLMg1/VE8t08gmKcETFcejTOn4Lq35Mgm1Bq5C6PVL2VmIr4HUybnNq
dY29pVpwrgbWZA0sJJRA7dZVGWu1r/JJQnnA8PBsc+CK1IepYclOhARvvSpaYSoh
K+L/edjjdWNQh8HtUPcfVrc7iA8JLsmIX+Yk1ivbWdu0f1q/4fpyLic8rHDSH0Fa
u43dD7TFf0Lu0a8W8qy8mWJq7/Jg9Saetb7Oz2lM5RDy8UWgbhdH5zTeCko6rNBe
OBic2V1ldcBhBRv8LZYyupnRkJ2GhbmlACef6eqylzBnRXX4XJaHa6LIXDQtROsm
7Sq36N17OxLpCKNH3x5Awd3D8Z7jC5Pd4LPG+/VRGQBMhbUd9No97Fro8fd1PZXh
x0Ls36JwV2H7F0wuJisjvw/6m84EuBxbb4LVy/S0aR6RDX3Vf1h6CetrySDC3t2F
47ylNli/y2PPfFTuUAKN80xonk3cV4/yPiovFlh8Tv4+nCoBUGffvPEA9aTkOUqZ
O39kFnLgE+DTA0AcKovKpE2GXWtgfBGDRmt9bY4bkdx6Vt0NqStBoiJ0pNtv2xnq
oElkKUX1tb7J3T90ff2cO2+xxkvKoySDCDlBsAkh9CnGBDCewKLd3em9odbXeynT
AaMZ7wm4dUgTYsmcfT8MCPDPKYu3HsZbeh9HxPRS9DAgxnIVq/5W1FtWd732/FEy
C8h/Z4sZSCkwVIAIbPhkAxdm44zwgotKk2e50IWbHbpFFYK+5crfA4/KpZRYo/S7
OfkE6JaSBDqCE+VafFB+aINuWIDxPl/QxwgMBYKT2TJ4tE59c74JN47AZjlWoIJb
TGspgJ8nx2H6AQCblZ+iZI0YLGqGPXBnLpMCjw9SPDoNiZ/rxOO970W9Q1vDjWpM
UgMrR6wYweT8Q5ydF8+64GLMX3S3VK+fF5uDeP1OhAZiSnuEIbIOq1mpXpY9C1+A
ymcvaQVYYjs6WN9g6N3s487altSpcsedokapKbJfdghYNtqkGlcdlXvdpLQBinFP
1dGjxn6G1/rat3SHCfmxSg5K2pFgjsEcHiHpTCOUhbdF2eRwIqDV3GMq3+oGax6I
Bw/LEY4AFDhf2ShNeckF/n67WLeIAQn9uMfL8xw5b6ObPGQQUBeEYfKoubcofnlI
aNsrb8kyzezqC3x1XkjdEyehng8791e4kG6Gyfx4H9jGrKOFknuzFQ54fuKayMCN
ZQZLxpE3ewc7E76QwBFOdNBZOb+doco26+6tfMQ09PTr1aSJgPzpCTBu0uWHyI3j
q2FjcO8dkqNtGxPxCP0nXVRpqbuB7tWk7K9+3rPf1Kzm+YS6z4mD+wVH+Qpoq37e
JpPBGLzFrtetWc1vhV6TIs9GyvNrddwoNGHPx57mwaFKrt5xsg0zG7ynCZf0k4/o
OQ8RuLYZ73McyMXojASMlNjjdhL3zO/jr2mrlfCVHj5edpykp1NeapA24+rfFcuR
bdrpWGPAACnzDfNZoa+L1G0tyjWqFVqn3SXhO7GU2QPH+PJyS92Z17Z3sWrd34ad
PghqVifdqyKjl98vrJW6JfZWePUCbGjEGTbtskYeUO6atnNu+fWk9XGV6vaBUv3Q
AAGh6XULldmrZj+ic7ntb3ziTBEDSeP9t4NwvXSxLqjrZAqHQ3fCGDfZv76y22YR
SDJDMV7znQ4YGGzR8YE7br9NFqfBMduw4ZQgdA4AtNZBVTwbCTfQqLtVNtcaDpS7
5L4ikK8xBahdB4CPT406ArJ2hzDB4b5QNn9X6Ce4wl3C8D3vWiQ4KWnMVkZKoT2i
qwlLa54IFWaLan2vbhzlcoKYUeZ7A1+7BuobNZuu4bZQ191ktntFuZIhqzau6irY
ajrw19PSUF3cfqM9R2iS7/aFQiM/pojGXj5KJuxLgDlIJXgUhO9g2qIk8TWTENg5
VNgqJ1V05S+Su8t3aB5T9z3hGlWIPsi7efZdGCe5RsEcmbqG3ZLM/Vomrcqh8iL8
e0psFQ8tbLPxTSr5yOX00/ikCUxDLBRMHlS4siHY7Ywpc0a042G4ZL0QKycRdBrP
t2HhkeJrfsamdpLW/nRvXcpKo6VPZiEiWYtZHDt/nUIS7I1/vZLoDwOW/qlSsE5k
gCUrGrbM//YhWW8BY/BKX+3tw14ur//l6Y26CRkWQLjgSx8L96b+eIo4BnIm1tqr
y8tm9wt9fnPxpVZZOHXVgF4PeHnTfE+PaGDvAhL4JoHkfIkozfGVBr++LTU3rPis
84DAtVTx+xWliPQb6VMtKBaFf63938jlTFZ/hk6E8ANVgGWJsTtaXHrTMIsE+1sj
aOnhscPXknunstW1Hj4o7guIGL9Yhww7NkJPblOa1XklG4gdTgEtIw3GgsBIe44j
jZqsja4bxuj+6nbHB+qCPgsnC8kA726G6OdwNjvED4DnsuE7Eyg6HdUme2I0uaq6
3OyTJ3hLDdFh2YaQoxMgda2t0Rx/D8VDQn6YCWeQJ66e2OEpZtnZZ7ccdwslDKUz
aUHdsEeTs3XqabqjVbnayZbIoOQBLuoJrcxOUxKBPVG/v870NxiQ4aLFRqftGJFX
hWHHiUuHkLgRTZ6PfCwBirvNeGQpuWEC4BFnVQxiCp0IH/Y3sdxguZfPaZ7qqZaU
NosFhmlaf7BimZkw0cf6cSqbgkkiKlWmrhL5sPOqykEg/saXwEsamAL2QiSgWDvx
1lcojPdcJ/1SX4gkpd2+Yfq7QckJ3vqkYl23uMdriSGtaAI1nLi5OcYTPvWrxKGI
4wLcIwwFILk+Fd6EMaTyEw7dvZA6ZlksL5GYgIjr6gAkVWV7ALmWW5EE0DJykqDJ
Iwn8ABLYpbs5HhnGXeCiPC64ay+94hPmALjwrcsYDp9MPsPivOoBZPGR0FHOCBww
He1vEJOoMdYk9sT/VKtXviHYC1t831APpfT7kz1/l5lsgqKMoFDY4vj2ebxefB8i
yU/ofysnU6yYhCXBwq/bP4ukCcSx1lgVMUqF4Cm/zFSobP5jaXFQHmtx/synMQgl
qJ1GWMYJ8101EDAAij0FQoLDucqx23I6udueX9wtmPENNXTz7b4YRnsVbG/e87V+
n7TBEENPm9wNAx/CMPRNACsHz03uHioK+WvvtxFHN4NCMS/z7N8MGkzI/InD+Jmz
7uhLnsNzXLyXfU7XNxIpTAOYILhlQ+OPC6THWSkOAmjF5gz3phlQphKx/2mdY+rs
EwMyT0UXQrveYklZecY0LmIScyd9nFWEX0Mp29dfj9p0aNrFb+KtkWRikEMd5rj1
5u9F1QSpk6EOEyA2ioLw3mzmqfCnivENFke4Do258Ur1NAhdXugKN2X89eqyIa7w
XrfAUKflluT5bHaZ9VJSiN3L1rJo/HOvQr/t6/Cbu9BpLOL/DCGUZARRQW9n0Dto
N7m/O+FTTiHM5ih7350g43iK2hONF7Sh3ulAarqeGTwTZEJgsHaGGQA7bW1jT+Ll
KdsxSt6QN5J2pedpkLqzX7AMWg1RF2P8vFHvz2FXy87h8ulAzG9amksdEwDSATzt
kg2BPUfxhC4iVxOUCjB8ldU4gSaFZzqNEDhR5WEsCc+zmjA1QGrYF22O5OV+2jam
hDHMhC0sXP3WHZSIY4wrFfB73mZi8RNbfEt01xERmYbyBtIxAL8idiKUh8QUsPx9
iwD0OxpGSnsfzbrjP5S9pTKdAawA4Gu2QEK2kE977aTNZBW6OuZdL9UP83F3jr02
Zv8gUN2Rn2suvuDo9POhYiaMiXSCJKi3x9yDjYDqD2DRQefxHnlwABoBxQJGtTMQ
8yG74unjZq99o79x/f+pGI/SpZcBT8Xano9CsxmR8Jnu9AhX8Osr5fBsnZuBhHla
3ehF4437fPSsXGxJCyE/yP8ZLMMu2LOB9CFWdFiaNZ5HvVxwt33vRlmcwgUF7nGj
LjRoHJdPXXq7JAd+i+YV9+m3rlhQ9/3Wkgzz0DFtIRix7DQddayKiULcRrSKtncI
mYUaVOuN+EquKkUL1IjS9Rt9qeRdN31GE4pozFej4PAiesua+umfN8Ubsu589E4w
dB3BKnv1GvQLkUOAu6cOjRKHBEB6M39WX4ec8sm+qcm3rg5zMj8EHtwZ5bIIklnC
YGqJaOczAdv2d9E49KfD3uxVZMuTf6X+Ty/KQS1qCDZiFknEt+udEChbSEc4Kh2j
ONTQ0tGlVuRGDh3S3z/+EFlHVV0DOn+0ljcfHym4yMAYX08dU1AznboIw45dKIJ9
rcWraSTvnu9+6qO5zRg8N6n0oly9wz4bcXBiFJuH+MpLbXUucFZ9QuzVOQ56baoX
oq9nDz1z8j2XKecDhGbBM0w0aEkbt9hPLpClFvmbI23pACLc1dKU16knoysbJheQ
XD95hjIg3wqblUE1u9Qus/KvzAcEj28H2d3D46gX4ec9ZZIh3lDRvpcXBYZdQXh7
mjP4I5BnORvWqCTPSwZffS/HENzPYG6E7rdw+lPbOHJMEOGsETm1DX3NVBU4Yy0i
wOQRzIyCl1KBrE24/lYAdDvDoYWc3WeY3A8YIKrh9/p01C/wGIr/KkZBZq8yTQiu
PAShAMoa07wUyOR5rnvs15ey4UIXz1g++8Gmyf/XcQD//wiMGAnbMiezxpqyEQUy
+L8HylrBsjLZ2QsMKxvbqBmmb5YuQNa/ejlZC2NaB7ziLCLzzbr+rJGW5b9WW/dB
iFch35aHcZEO6pYVbfRsvW+PY+YjWa84PPYF0M++bZ3+2wFhR6XT170uDQ9mvMMT
np5v6CSFDoenTeJobMtQUd/NiBXcTBeshOuImJe9GJWibIyFvjRBIKQtGs3u361Y
W5r00k0MNwMR5HdNEijauGFEM+yzeBx6p3EY4HAP+tILkbqC26suG1u+kcZwZvjf
YIPOGjTUHGS9eb9sPgore1XEPF4GBRyWYbQgYQkQuVddWpDH2i2sslaLuB9vcl9Y
W249VxZUm4uvQ3y6ce9IeSeBZMrBBNKkLvRGOD4Vgkm98DeLixIj1I1DmgGJ9hct
SRIJ861thXUz2g44OWtDNZ9aTMJ87hGT94vlONedzo62eZyyZ8bJy+8kyO4LUI0L
NofskheI31nQVP3u4+2ft2Tq40yqvn27sB6CqMLM4zhUV2EZURUE5rDOh1r08Uni
e1Trecp7IgTZ6PerffK1KjWKsg9VETZLV971h5OVZxlX8LpwC7sH/ztB2uM/HL6N
DBdMiLOuzigetxngCBtqe7B9/Fyqg9KhIZfyO1g1NbT6G4b2Q0QJCSG4ttD76AzK
HyxIFm85E6p46nNWkLCFjGE0my84sWBBODelBHlZjHjmu/pfnCd2khXqW6TzlWUU
uTRr02nOXtLbwOKoi3a4Phaagh/8PvTwo8Sb2L+EIQAsfHnwf+ZJWjnVlXZjqWnn
4aDgLwSlYpIc+I8s2TsehJGDVxD8iAgnsAGQ1UCzsx6UXYXvEkN0vv46XXhRIFFH
W5WVSJb9tcPcaigoaoFpPEDToeRVMZTTOZbyx/TM0OkkANxr/Mw+HW0e0pk7nX/Z
QpB8mtA0eNfi3Lxlh34Sm2vouVO7KPjc1ObHUhrepZCAX7Zyps+KswssVL8Jsma4
zFjbNM7e+misuJB0crih+Bd5Tpu7Wipbxxtwl5OEloq8CykTVgS3HqS01Z785zJX
OWjiLDdJquiRwN3SX/TQ9OG8Oj22YPY4WrMcjcxBpstC8VoT87xW0tRZ2108V/th
dGHM3kJplP6HDte5Uvt6b6F1d/sv4UES0qJJY2huBqLFp92BMsmGCQdLWwplsN9w
W9qo3F9Cl5lONR2pR1XlXPTMka6DpejWcjyxD/8D3ipAPmu2KMnpGfL59DySujny
Wk+W+XZoAruYshaQytQ3y9jc1aEpmr/ux/pWO1gryEU2BNKxxyyIV/OLjSM8Hqd3
v+kySUSdanNc5pLvvdAsXJ/3QC08cq1npcTPBDZORexic7QnUeDU6DPaODyJqsKc
87IM+9ebagQCHeyalZtGJwP5Ad0/t6p/qo8gXq0IoWbpvr321gjan7+f02/RvVAH
uIk0fuviz7XBIKewJCqwOBDZIgWNM8RT9owJceLHkxZNfEJKBttEysoBjcURVSAT
Dt4xlwHyDqbiAQ9xTcnPCgzrWbibtt4F7O3KQ+C324og/7HlxkAmBrq5C7s0h31k
bZJ4xsx5iOUkkzPJSQ4OM8Bn1KybO0R1Cx0ePyo26+UkCf1wGhmwHa9XP/LMdHUk
Oc0/JP8iBmGxC4efL5Bn6Ywv/lAikOyDQdqG4183pRg/YmbN7dZJZZ+5sOatFcg3
IeiF0xXaHWSTOSwOjouns39nUaxCsMqha0Hd7GsAOWHWBq5I9FwwVEIHlOxthEcH
J7/XWsnBfth4BgUjFK3uvZDscCiZ/UedJnLNdL5rsWpQVdZZGmXBLMI+qbtgIEvI
E8paLx5ZvGfTMlDxTKcQ/vmzPhP1mRm9TAvd4tedPyCry0lVq9Y32MSO+7ed38rU
tBwKzdzFmVDOlyEi1jJ37r+hPPldVZhcM+0B8kYYcPIJaXGGIVWudUfFlN4OKOkq
eRqQCmOMD96Lw61kc7hRlXbJdCHPUhQlfGUeg9g35zDH9dUdg4lOJ8BrIirMlM8u
T3mz5QTsDPJIAfaZ8xLfRShAB+oLAVKTIfvQLdUUUgh6XFjPIozZDh+oU76jnRZB
zDxlUKGqFSamD6WbOHPshtBOqz1m4RliLJxDIzPK9qYt9GeCD/eafjDTBFIyY02X
g1f/sYLgAHEYRpJ7//Sh/7rkU8xUOah3KWLe0QyT1I8CjhCQcyRdrp+IcjHp/4iv
x4oJSEUzFq+EUOKZ/dX1PqWv9M6XYDK6oV39gD3QvCzg0kqye07lIGAQ3qA12p7X
yCCzegIbdVzI/hnEugMQXuiAAtTPQX49yRzJ4hlgG4V0sPPychkpp47tempsQBX/
/CLYuW1Lkgx/yAAzJRANYIRvcOFmDeYhNXJDgK6xfjG+MQod0BdJfJZFazPJSP+j
VBDUzSPOGR9lAAvzuNCRpwV0tSFZ1QXbpE1xxtp04i7PdTE1QCLvqTG0OBstQSMd
g3PIk48ImzX7c+u0vdKP3CC8MOjR4G37kmsTGHPB715I4sa8axAF0RcFYLFH26od
qt5cKuagSUGCpB5fATc5xq/a5vHMOH1ZBMgZmYn3+BwW91QmgGKT3s7EdFQZIYLd
t+0xLnpvoToBGF+2V5EqU/Qt5d1efNkAqgMaEyjonp034WbCOuNTHAsAKKUyJxAc
Qe3XbDSpY8OAGZaTz7JpUh4x3cJFf2BGG8UQ1+1hyyVLsoxeVpG1UlucgEEQq7pU
hzoet4ee53NbHQHiSQFEe9pLXdK79FPkh9XfOjFRUakaJ2h3unh4fvbHl3AJ+hBs
Zp08byXQpRfINdfynxiS8qWcJ2zSFSKqFhmPDBc61BSXQNhFjXOpBHpAuZjsujEQ
ZDZMJOM3R7vKEsZ/6jZW9BNWxl+biMxQ9kxzeht90vb7DnDe2ARlHdAEQ0B4n+EZ
DcSnsPFJEb/Ro0Q8PgtashpefinbvHy8U1bJuEnjkH6yqpCkh50BJeMo8lJdsZKu
AK4vpS/VxmJEj08yOHpQC0yh1J+z/NBJzi4KoUgkC+3ZKoVoMrp5HMKyMZLrST2V
ZtjVAk4eLsMUhZss4+y+q3198xUyqwtSU7+ABdQ3Ms0fuMPC4XtYg2Vml3sS1asX
MpJUmdGqVnwdIsYjwA1kCjdVkGtBAo9lC6jX0/Lo+nS2Ctx9vTulVIkngBQdo9DM
eXO2A5hU/ULj5FG7xdIAxHfNukVNy5A9nOkJlfakxalMiXNFgguhESad1mQXzBK7
P02Xl2sghHky9oSFaNQwWgzOqEzZQiCp0noYtNKZHGPcHrVkVFtEe8MKmfE36tNU
jXs5bhpBI47+ikGXQGnVZ7/AjkF+9znut/e482/ebDx7ig66k+VKmTQmI+uvfy4K
CMdQTziIhBQxsbT37wzXsGw2eEBj+gRBUiZKh8lW5d2hbhWZ1zxq8kdSePh0omp8
uZYIaYoQoWA5O/iAQZ0zCq26NchbzFBT6Ht/wIXR1EyGqTRzcFgGGFtQXwD0CEG0
/Q7dg7QKuy2SQ8nKblNTOtcMMGGoav/TfW9HShRx4sVDorQSmyoS2+bgYc4z9Kz3
J+lo6Lg1sLoIPQ+pVu5qOmqDncMK8h2wVlAa3dx44XefqvbCcYNFRAHFTrdeA3MS
eqrrZhb9f7q71LB7ZlRcz+viG2DXoEWCkggzeIg98v5/du6wg1Oj8A/yn9h2+CfU
8ika74y5p3DMaR0GBfPMw3uvF52OyLb7BflQ1wOth91ZTFvfnji/VcvDgNK1aUyl
0IgFgtN6NQ9E0QFP4TTT8WNHGBwZtHYnLro2sW+1NoY/sh0rHKZnyGimjzG8zSu1
6TidKVyvw8Ez1pTXLQArLhXvDT68qC7m5oOjAuWPGwnJO1Ep11qV0wRfNpOp4XoA
xe6phDAHFf5bd6bNABZY1lOjr9NqEEHguMBhZNxbYy8uVJpxeDjltW4g35gH4/CS
7PTOMKuzEG1fS3lxqnZcJlR9GpYA9tF860bFjTsHun/bxuTsXXzfQ9nQmYBkUVr9
EQr7rTSvNX8w6ABSeUtiKJddz9is5jTFjGPJ93DVysVZMp7Nei6fq7H+0kkIg2Jp
LqmIoXxBClTduJKj7YN1pIf7wEW3JyjPbzAr4r2+6zP8pfth8gGJz0uFSnng3tlv
WEQ1mWVqO1HHk6d5txPhDEIrt71yJXU4Q/m8jU/gk4ENdiZInGwycKLMpmiJvnoj
QTl5dooGmo00460XbGonFzyC+QTqmlnR/PIKH8h+WLjPO2GBlkt0QAWbvtdVRD31
i0x/LoLOuRHRgLzpH07ytR4kOpZ5xY3QYEqf84qZ5gs1lbNULNxASHCSgk8CG8CE
0aZqT7arOki/movB49zZbz3LnhfVAGvM00iT4B7VW4uvRoh/ZoZu/ikrQsbsxUWf
BNNDcgLRqacIxU5W20AxKQgW6azBED/fM74yixpXb6Gp4FGlD28rexuOUvTA0bGV
qF3m1/M5n5SqSFFBd+hF1INatQ9Ss/SJYUIs/3Oow9FW8HFx7zXbgpt0szKbWswr
Comh0XHLgsp5qL8ReAa5xDU2QQ+tl5AggYXu9jfrPJ5wZ2xB6nXTz9sCnrw8VjHz
HRu91FXVz/3GULKbnHUM+QeoCSRebusZPLNmoCY6oM6GdCTUhzftwkT5vKAptCwc
E+8KBWQ0/hYaIm4ikDFSle0sYqJArSGNDU9t9gSwMRDhBkJY8o1oAlf4o05VrKGQ
2PByPSZe/eeOpKySfmH1FcvgHDE6qaQkNg7B8ApKCkg7xBsYMEdKoV+UiwgFPTjl
0skrzR1TdihvGHZc70z8//FOI3nqI5dFey2/ROQkf809SpL6QLvfEg6jYUbaScgH
BY8A4h32GElaYkibdgRjb2rywum1QpQDwoJUmzaC6uKOt/HGU3ByZjZgAvbjNPvz
wBaU5R1eCzjUIeg4aijUr/6x2R2tb72OEIWGz6nSFLBu82NNL3fcT3frH8/+SWjc
5j4kA9TEL+S35h1gpm1QsEuE05OpH4rJY6W/RTaoqopa7sSbgzrNLljIYRFJR/N8
vM9iM6VvcYviz/y5NqZOFnLxjq+mNA9wbJw6XZ4MXa4t14NgEVsGJ717gdI0J1eL
//A0tzxyfSW9JNaTj2XPqnsDGPPRqeA5wwFZqPHoG5FU6jPq8x7lLlu+WQAGLgMJ
8u6Gcm+3Sh9rfhvFIL+wiTD3alGul9252xfUZV0m/K6+c0E2pcTg7ktGPo2i55P1
/eiweIM4wGChHGCTJa6pcJmM9ic6sYlE/gCiTrQWoROJeX+Rk9NvwRJTtnrZJp3c
4+Qylf/9r4cHtaESFr1AzaO13HMtqmEKaKOqBmqhYMsO8zTDt3pFnIFog/tm3ZH0
4GVKcJxPnt4XJT+fpRq+imyz+oq2WbLGOGLHuX6PoIYCXhNGC0nG/bt9MoCcEljw
T1pxdA4qm0Lk8LPw6R8O4N1/6qpyvW3NYT+EANQY5zYD7K1PDUO4ArPBsFPIDZt6
LBw0KVerIeoX/TN5rTZIGPjn30Z/901Hw+XhpfO02QCjtpMZo7S0nmQkfInYMCY9
zpmM+E2nXHiFZcVOs6mxLG7pOUN+R97iRijh+VtgFORDSVhI2NGmB7vx6HZRZ1q1
Qw0bl0YlYMkUt2cbgFZX/YvcqQza7rPtEpVrEU5TM0QY6hPZWU+Qat9Las/jk6yP
+4gLQm0+qcLVtrfy2jITIwiUX/7eWXsxjDeP00c2bNHD/WqIf6aSGusQRNHYoEBY
BzqL1OpXZXy9hzY+GsQFbKWAEaI2kKPjvmQqBDtGlA3dd+ZiZN2Y/PTMmwf5CojV
JZLYV9s+dgkHQZTJHwUVtjwHpasNA96Tu6YmjUAlxfHkdNPQBLEQJZ2A97HA4XK3
Sf73MUrLGs3ISksVY7toipraGixk7RA3vtscOez/8WXBqmuZIxpnFsM3GLkEoPOf
EYm82GhJ4WKrI61UjnbST3kKeazXIqLb75G7ee0Tu5h8JIM/tg1bSCdmRRmmpL+I
Pb3jc7F81GqZMIikDPw9+YwtllhKM2ALMMMvYJwPXdSAYxLN22ap5Mv5N6MBKaJZ
T1b3IYmkNByhQUv5ZyXE0AiVh35Dms5cWL0OX344/o7nnGHXQuM9XDP0ct/naeij
wA9xvTy99nFGQ96raq0Jr49j6MkGedU3cWfnMFAbn+slcDou2VNDGhf3RCJa9WP5
ChXfjeC78OCQKtoarwzjs18+27FyyD2B49nX7HnmglYVwnAZ+ONnKis9B5lmLWL1
e0nf9niz4j663TxDxTmbkt0E037tfqd+tLThgjg32vMRVF4ujI4WQKO5n1a8taRV
+ngfm/qq+ZzKGp+1Nd4lJp+V4x+rYutrYhj/Yy0jK/CMmswirx9LxtE9eilrp9LQ
sWqd20SKSBz0DidtCFj+PqiYamQSCqMMWSYhlAGf3dTsY+NXzoomIqROkp1bkRF9
ls2RJKDBvD9S6Xu7GxndWcsJjqo1KTddEMEfTMG8VQwbqrVEfHuXltiYpkvaNcK5
E+fenAbUbd6VQLZNTLZbXO1RlAbv/vNPbLNAn17/iYz1ZTtRabh3JJb5aYUK2Duo
I8iFdIPo9KBEHn5e72onu6HnaONuJgS1SVDT0+MDNqNPTUYDRUT0CGpozcraXJoT
a1pft9IIuoKXJkSdMN/yZ4EdcPHGCKe5wk1EWTiHJDH7aGu+TTM3luTqh//emKff
aF946kwOweiDIe1cw8XkfVu3qOB4YBx+tnrBN5KbJ7ursHI3xa25qttA4CvQGq68
27KuaFPE+2WaBzi4ppbYiiJ96fJ8TubaSGY3iUOb/lIZrlGya6/Kx09pZdGcTr92
Mnjf2OB6xPZdM1r6FzzAELzXSZXSnIwNEqb8SvZB1B7Rm7ZdVVAGVTHysO3zqL8t
A8F/6dXEtlJI2lHh2uujNdZKQ+sJUWimnWKxReK0DSki5ML5V2TdtUQsCW35Ohy1
6xHbhllbXM8Bf/NnN3UK5Yt6HnZ4/ulDClf8gvGBrW7A0mK1q4FyrkebR7OjsTev
hvVrpTyOgyBNzPZyBv5OPsDnmuY4Qcdmoczi+z5NIHxqAcuuFtJEEidEIQaJlEAx
yolHLLGOFj/OSMykczlZu7vTZXomlcBPO523K6nT9KUmYxgDxC1xn/PtjoL4HyJB
4EpWdI40a9vEC3JNQGoAVvrRdOPQYpkUlx2gLAdouj8e2NIEiX6XIPtbFPuTynut
sXt6ei8F0nXWdmbCBiqVmcHIesdjsGFTGTkqh1OojpfmDUaWa247UOJ0QHwcsPRX
h4s+3oQmLSrV9oP9ZfnU/o2N/0X4lnI0NVJk56AV7Pl6lI0kJxTt1D++kQhU9u1r
m6z1jl0o/R0llTkJQxppXdOMKbBRWPuDdK6iOjyq1HBpn4/3LiUZvTxq/VaZ1+m1
ozniEDOlSX+s34PID3EizDjmffjGay+i5peQfn2naqRrUrhTwMzjLgrMBFnvWwWJ
U2bT+rAWdL7V2kpBKfOevqpJfUJED23Rqv344qOhdoeCMldkyXcB5biXSLi+hKWW
pya0KEzQOO/9/QYPITDpypqnKMqoQrouKRdre4/BTr15Ts2Koy4BpNmsQvsSzjjp
Xn2AXuwRMRh0FxCL9xcaxiHyuDqyVc4Y11Ri5ZxFByrjG8WaQAXQ37z/RzH0pMJF
ikCmfi0fqK3jJdkhsvKGkD20FNvM24/4AexB9LZ8NehcCjNGl53JyGNRCpc7A6G7
D+013k8xfP83B+ab3tONtD3Y43gjPwlTEgt+2Hve1UAD0HRVmyZyEn/KVjfNmF+o
TYy8uQ2Z/SnNnFPer3B4kBUYRNfQpJq7Wo9d1d475snBgvKyfB6m1YPodp2ozcHu
Vr2pku/cVACv6M07e61nCLE72e0miEMZhTSnoVnQNjm+QoTBPhKiFZFVMi08QGe6
OdqlGXUPvnsB1YwRYtm1ST6dtcrIEe68AvnBd8ntaRQj2JoEW6c2JYN3DV4TBFcF
szS6b1VILROg0c3iSfeDode3z2a4Jm5d0k/pp2XlGWOSk+TXv3sZ9J3oSuwY+M8u
uPs5zmlISVot2g0u3gQPjUG2Ztj4mnuToaJ2lDKpA5y42Kp0Pz7Q9DN1prHr20nl
VrGHXq5Xk4e8DKHlfDJB3EbfGvSIQmf+PPBtXsVrRPVj71o92+szRnXLDUz9RjYh
TmoHHY3AVIkcW4td3BtsFeQ9cBt6PoizpHgZdUbwsPL5c1CmMtAC048xAzb96fvw
QGmFoH+w1QI6tzOi8jaVePXHwL9E1JuQycBI/ItikijmW0pzOc5YHkSGfcooVeWG
gsuvn+ccEtzYbLPs8ZnuYOjlkQWcPWcsE4lCzmNfgl8ni1MHhwk4lcEzau3r8Yqm
1s7rY8UzlFBc0EzP0z4KeCkT3GfzI4oizqJgsa/Eb7a0KpSicIfECF0SSRSQd9aa
pyN8s1uAUjuuCXpwhWTSeqD5BSIwQWzwSJn54YU/SF9Y9rXCHjV+JKTV8hDGYVeZ
EseizO/Jlts3wqHF45lWA+XRWZzyL/gSzDF62r6kT76xLl8B63WykXnu6dXUNAeH
fTY7yb+PmRWNv1WNBCgX3W7ooRrNVgkEVlGvrUq6jDFbz8Z34/588a2/nvUjavjc
Tg3lUxvh6y623VvogpYbS8UtooH7pSc5QzNtyUmco/GSb+KdPkiBgdIIsFPfu6/K
YIsvYI17M0WXHMP0g50OiZSZwisgcd6fAKe1bIbDW2yCfHi6tzhA15KXdIPfu9Vu
tm20DPTKN6pQtTcbeVwkLVCWiYXhsf0ZNdX89G+EvKpwutisaGGLW8xfrJ57AfTG
Nnh1oZssTZ0AE/cKd7jfTYpgR1y1cU3Lt2hXtyEimuGKW3wu8Prq+NMg/aKqIpTy
OT8yTSQI/jrEGXnjlpJqgL7ao/J30MH1U19JFE7IuKvRkIVwLAc6D+WYPYhi6aHX
7sGv7McNvQ3YAZWAAEvOftWpMx8WkYaYydX1GgY2g4A3923utQUVpIYpLpOjsMhg
p5IBARIoaUVPGjbIbLdmupZpkhMHAXmCNERarc+QMrr2jrCr7u2ewhfodcPrCdlr
/KOhan2ZdyzXAa/q3Ggn2x8Kkx0ahME4R24N8yOVMq1LfJyeTjeGrQvYjoRar1OG
ESl0eRUExh3z1yJdQGCx8+hLkB8rRwmtvR8/6Uk1lnvCvSe+FNZkJD1EyQq5D+GH
kKX/SbhSUtmMd2lYzqi3AKspWqD1AZK14YhlTCyLSzxnQTB2Kfh5oDnbJdZdlzU5
CgATsEDLTWNcHgXkj5QZQq8TRi0LZk4/DkCIP24m1IMctNXHchZDkUCIgwUCumHZ
3wtvIr8z208mmRNNg+XDh1NB7svcSgakE3a626Oxd0C2nWaAK2oo4kz/p99nN/8e
5lDAy2PNM2R2TGDtC1ZQ1AaytBC2etdq2QFONKijFIzTvvSnGtJv8xm//ywseoW5
G5KSnli8oKCoaFVX5BjlpYkj0pKfxQrC32Dbh1x8xO/tR6BukrRg6GXDln0M3Guz
tZikx2dWUZk9mxZVjDPz1mF/cYSS+mTybULSR05W+Gj3jDQ9MhL3pd6MapUUurpQ
6i7MgPMZvgSqwP2bxqmISsLDYf9c1Dsm3kaveyLS3Ha51bnmaPsaL732DAPnzZgY
IGM7rkKnNPPm2wjTITV6G7Q0gldpQjhL4a2BE0N25Aq7B76zmTwMSJqQYYYin8QS
8gnEWCnfW7+zi9pDM15Zq7zsFAq/S6kWTZiua+9G9xIcwxROOGTEjc31UN2tBvF4
feSkBPJeiPGEIFNJZUl8RxofLsiP2A1UeUWif9c8sHgU/nGVkRiDvPYB3Atrg5XU
VxuJpRHb/hF07UwryGWp5Cvl8MJsd6u3ofO+Ej0aeFuamwiRpUIdvbci0Mxc/Zt0
qEjx5YAU+Kc0J8dKgBikfhi6vZOnxVm7nZkY5cVhP17BzITzwLENQwQg/7f3OaIQ
XrIwk39K/wMc+Ag77rz+NraVSHu2NneMPpYYx5jOEl0Hm7vnenEs+xKQZZ/HyQzK
7AdnOF5LXuEJteQsSjmDtL+K0Y1+rtXFIxL5pt48MQdNpUoa4A2ykoBj7+/JTzSv
c1+k2/KuElXVU2YxSZ1dFG/ztu6PGsuFHz/hAfXxycwXPr7eRtCSYKC+j5jrBHx7
+B7FnBn2J+V2K7KsdRUyqjj2zOQoSLFUfYaPhiETHz5m90e+hZ1u/3JGIFvJ0J4a
fUh1jII4S7x6XovK1+5lqU4av7yOrdPJAss10IlZ3SgWGxX3GC0FHS9CkrswtrwW
JoGLvVNVyfIeZLWXKre6a2vgHxvJZoYKlSrC5uuHi+C/OQKf8J1oV7Vfak8G4cYj
XUAtC1a6EXTOm7wwVTT6wkAFGwB3LEznKuPIcyMB/QzaMYX1CRMdxf7oP48XSYzm
Fj7Tsl1ig9M1Ws2lJBdI6cGVBmVoJqUyhLHu3n5FbdxlZrK+ZM/V2gCdGEKNVyGo
4ZU7qMzJcGd/5Z3b3Oy3cimPf3yqudemLjWnughryfbUN2TgEDppVsFqAAHc7s2g
aOTRvWw4lBycicFnxVWwkLDAuR0t0o8b18wogsDA1whJtuySwpDPHJ0sLgSVrxeV
/plxQK3QHbmbPO66tGiKSEpW2odPzUWN3wy6YDZBXAFHtR9KRIXqT+yrZwBCxWZ8
MOf/1WP3LAJ1JTG5tuIaI4DaxFMzirokPMEmLWdap7daJMD0UVILCOime1DGJo9v
WaGpinu6kjFIGI0whds+JKhioM8UQVhu0Ef5vqndrlwJ7qHMcu90LtZ6t+RX+hH0
0mdPL9+vAPUMVkGWG83PCKIKnFbCiTSqDeyGiwtQ9owWs6ZXgRCOq/bwTPGCHOZ0
BYRWV0haymGhxw7ck7ACUjconQhzyR57o+ZIqcSMmjvS32q6Kb6NHOG6rEnNqaTz
Do/VBgNCAP643zhfgKfZMCH+M3qos+qS6AZcQkDRvgE9PUU9cLXxu7wEZNuRalla
hv8MVtWb4IJPu5KtKxKuSXoJmBDTvviNmC5jdqN7ykhZXWD/lY2GodG36OWataqf
UMLwVzYxMBpHBK32emuScVj+4B/GLSVXuqXgSVP/vNr/JKtXFRE7nd9Pfpn8SwbR
E6ArFWgCZCLghD7B/PlTRa5as39yUIMOX4tQou26TJX118B2ffp/+OhYUKUsRrX9
JnsmX8Vxf2e07wEQjMpd+VhM7scvzoivF6NjZJYJcUaLScLtE2T7GY8SBp6SvPTL
ZnW0lvbGgSchwmQ5xmEz5MEiY7+5PHWtXccq0k0aPlQPaLngThwCgdCqhZbP9euo
UFmrlyFDk9jfVYLz8bkVDCqa2iPM8OYKWOMCm9qfVEsAQGNGRkFGMdo0+RVb81gG
fFOzY2diwTf+58vXxQ0khETNlcS33x0plq9yg6d+fY4Udfuj7/mTJ+fQLgrGMsUH
R7PodiJMCyXrSb6/n0UvB17xOt+K85a2fzRqFMGqozmudMjzR82SP8h7ogWqPkY7
riAuB1dzkeLZ7zUD9RzXbYvGPw4kn+7kGcXiARski1L7Re6Hx45QCD6rRkc+wT1r
/v+CVkfAyMJaDzxQ08Aft3NenVN2btK4hi6Oy7D2MwcGsZo3ngdzXyuu/glwOkBx
e5ttBhYAwN31JrsPsJXRltwQZd37qIF2b/ZxfJuDqUrQ36neNr7yJDggBZMdhUlm
GvUxv9P+IOM3NS/JasrFd7bRkqmMjFqTtzh4+Hrx7XV8S31h2SFvaeac2PjEIl75
ivDmEki0oErcYnCEu1SjTaaASmCTq8lVS262yC+uOJz+sKWYG5JUMEYRgtNAYJbe
IxNDxsTQ/VT0PtD7RBa7tZKiaINISW8mkajuJLQ54PIbH/0a7ouEvwYELDVQTizG
1WCTs4hqur7zSkiT+OuNf/CtupvFxBqj6XOwnv7rghKvBWjVwPvjWWtRvRIvjugi
YlJhR+DqebAhYhejOet9jDGG5ncf5wjeg+N6pTGU1Abbe+OE8War2zKKqXF/sPGt
heHomH07otppYb8sMBBGHk6nybAMr063G9qg9t0qpqdyZE0VnmejdLOtWcyHWHYD
+mCDUqEfGPK45e8GErmTHsoFNwUtkr4UM3OXWEpEEfPrVCw1rGA2CLLDUejk4uzR
k6TFYFEejgQvOizegt4LDGwDizDKi0/E0uks1CcyqA91tGjAycd4SlL0ukshmeVw
JiMIc0tASR7UBIwXPw5p3zNRRsJ5YG5gUtvi1aOcI8mmVDb1nfJPap1/Tc6VKkYT
8eQ5edf5pm1TCFIumtQXW3H8bzxVuISzSxe6roz7L4zMjEicyRHskaUsarToBzPO
kRGYtj9XnaJurv37jnwkYxiCTGkjjhp0qN8Mwc34OCwS9ZWTAlL4zQHwkfWxmQ8p
5Tu0aGb4Y8AMoBetQN2Q3EAWr8uiTjk7sLaeq+5rSxqsmAU9nppvJb7u7KNy8OpN
pOkC3uMgdpBiGb0yAyjNq6sKhM7of7mdsHuak7GCeTBVd1S8BN4xP/uyrSJ79GDQ
UlGhgLCSk+kmj/cvsPG+qvA01QuyHOYWcwEyxtgxOD/SXVgw9A/ppp3lnoU1cwCd
veUuBxDoh++7ISbXbQr9/DQIAjF5i2XKynav7NTJFFftnvIx2PYAK6oDJgd5V3lw
5Q2R309B3XeUyyi2zstiloeopSe3i3tTl2AwTDJKoTStRcWseIYHUw174stNoTu4
bWgy/iptmmPH5ig5onNT3jkR6izTvGS5ZTT+mXZSm9UKVg1PWoiBcWqSCh1RmBXg
cDLsi1amLfBsUV+xuZO6iWUkbSvfLGQxxqHGgT+MlovEvX3ZdCifKTwp6HospZtP
zD33q4NEo7esy/s2qpBK/oltyo3U4uo8xfhd9B6jYvY1sLbyTlwxsaZGH76tw8zD
c3MO/48xDXPdGRiLTyVvDL/ModWbbZ2P6HzTXqivxT3CrMNVOkyvqOsF/jBualQc
3vFUr29HdMONY8ApGS8amYGZEFw0Gh65i1XUnD5xWCJ7F6ErZvCrgVZr3p36Unyx
DSG5yyNUVV2vny7u55C+7z/gAjRF+7jkANJydRi7vYGnbzHT36ARE7M5CpZDvRGH
nfnhyn6xX0LsE5kTOCO9B/YDyZKNomKwxBng2QuBpg6KwdhqOpd4h1cvLu7eRqoG
b8ztvkIxF1mTe5BCD5+zp0XP5vZM6jbf9OT7faPmXRdTpkL8iv1vxExnXW8RuQtG
Xo+isyLTQp2LA4HQ6+buqTPhnVFxdECeBBR9RlKDGFtnkFRttgRLtHpNAha0MOYK
gYCRBjfu/jTStrXmJTTlozKe5pUFJ4BarsJWbFD15BqM9oL7yDHCl1YnSYxrEeeC
tQxDLhxrR28Pvd+lF7yO1mZu9Mz0peNSYyY8Mwj5vs6BRh6idVelJZOGFbG3ZyGC
yypNsIMEOBT2MAWTx6H3bfK0lp4+e9X8YSwmrvPNZwpkkVWB2qJS5wCr1DCpPVFV
bfgC/1rHHWCgoYv2eqeMPlN0dgQyY9+gbZ99PjspM+qjeL9kfpS3LsvDnXVMRh1o
ub4svUQdMsKgc4xi1bLG90ldvLkhkzHtxndbelL1CnIMYCgeis/tCDd/G2EK75KP
nj2KWKHlsGMIyaCa//QAnglkodB+4M8wMzXzcHPmKFg/PtnACA0VvtsACjnkix6E
vE/l5JZeFkSgHsMzckybdN5SEOMB/0unwqOb7Wvz1gghIn/HAowpDr2AOYX7oqWX
bSI5JSKPFK0Xo1Ltmyei8Zkt/Ft0vs+hqUE3YypWjbpWzlSMBwgiBGEjjBamtOx6
x1YPUzHkm63lQF/1DKxldM+NZHTfjgFTFaBCpfuEIFdMhimQcNhRMvxVA5Ziu9AJ
DporitjZtAKBpOlpe6bZkJQZG6rzimANrjdenpJJHk9l8S1pqwzqChp0/wv0oNuP
uGEl6FcMKJpIg81OVx8yHAvIfof0U3lYYC+pz5zcYuKOl6UAWg+babmtVCZcdtDo
ECGlRyaPdamWV3ZOihxUxXliJkb9M3QCez5LFoQJOet9hyEpBoYT4OiILa3rcReS
X2HDyjA3uLop5T0941nWXrOWNrWGbHZRFjZrKmRK2QezD9yuRuLcVFHgkEs6LtkX
PiOXqzlZszYaFELNLGwfsEXF68qh409wk+vzEo9Hgk4irL3NZavHdEgC5h/ACWtK
OwbCvl7V6TvAvAgqiKgUnpzOE+/q43Ebo9u9b8EsplY7+h2yT7HlZfrI26MI2bB/
MyBtMJtj5VwyU+yuztODew8/3qgZo55jByTHUts4KvaPpWbRfEwDN48R3+LSGbJb
U03fTJpP3DFcdgPX9meXiLNnH0pQCoAOUvxM1zz81BExJMS3qNWexhfRXmpGEIoK
L2JqDVmgRbrrmBEE624VddNv/5AjHLzJ4+BUWKwSOajp28ksGKs/eKsSw/iLoTu1
8YPfAHthzTLKgXHcCZNA1T9yk7A1AwxpepXayi8+Uw7PuoMbkMYLwjgKhoYgesFw
Vq6if70B+78hOcQh3kPML7pZ35hm4tK2WsNVk5aN9gWVjtSQzQWmINLfzhKyVaU0
/FV1bHB5AUxf54/CoKlfP+4L2fhc1H1lAJ5jH10P2DTu/E17g6RRahJpFZAkbifj
oHb3Dg9Bn+X8weX0+Pe52fdB4bTjePwZQQPG8EUwuSLiBH6iq3Q8rPCoo3tTCmn+
eiX/RV0R/guOPIudiT7cMXJsmcs7Rb6fYZPwusGWfVt3lNqilkxOvzaoEenxNQoq
13REhsPrfjGu40++MO35oAbM937U95kXK4wV74wtQ7I8YHSHohjPvW6S0iFlI4su
ojMq8Ds+9cfMLBwIYEUYmStJyUo6TOZ7Y/G7MmIhiprrSkc5B6YKQpb5c9h2VN0O
IlVl/B31h9sgJsjbP+i7W+MtK+MA6VOPgcwxN7f5+zQLCd6I0L28miYEmk/UV4s1
/IHD/X7hgHoZv9AvjuPAblecTGESUw1z8HBw7LugyQn/JxlgvX80RVvscNL8TbP8
on2b7YtOPBE2/x6G+X+ch7fOmHYZv2WwOfKASYqoEbC2ZgJp6tRt4kW8y+Vt39Yr
W/lQsxC2F8BHtqRHPIkKdCXNqaBO5+jEGdJsiDtmOcQgR6+xff2cupuopFhocmC0
eLJQjB1Vr3cNVAN9gFzhAaQav7aGlDKIi9kZ7pa9GF4Fecaqt70Gns4kmR4YRjqi
4jJw8cHc4SUptie4E9EwmWMDLfgi0CbUuN6FeEf63nph4ZjkB+6B0N5lzYIDIycM
MmFWjNb4g74/tX6ZvEdG8ojb1WcQnbsNTTb5ruInuhjptzLC5qRXk59oWg04YRXW
DNNpXT3MBaw2mHf8so1vkk9vhJ+Wsm8T0tqhQS/PdlT9bS8CGF3vTate9AQJXDSP
2w7L5kpLHNhhXf072GwFB9XtM8VHFlazQCmKUTA812OKYu3e0jNy4Cyg/vLdbMAg
VPzN52lwT2nPeKX1/W6GCLZWjLBMBYyqCo76hZ5plCuHNTYvAJTbKgWZ4TuEBk4t
T+pDlsh6xRqfoTveelqCFBgqS1l3iNpJulST1+BGyLkcMntfqIHmgVr2liPR+eNb
n4KtxYBN5sQtzIDRPDAKNd8KVgmEQtRL9mfCeYFVyDCtrCt3e+u4s++MREXMlyDK
AICwChOZr3Yk7cdyti+velXi3lcU5dqwlj1zjoWCaatd95kSuW61gl71fHjAJ9V8
zuIxiKSevJS1aN7oaIPmyuo46cBqYZWiMKV0l7NRbdbu+5zGIQqQbtI1yD2ekP6C
ZemKjo3+RwSpsP57KOlRflnq6xc5qKxHEh2iz0CXDqGPrSekvc+tXa/EMPgFSEru
IUDJ7216yFQyCSav77VFkK5tiPVj26A0PhaUAaPTPEQTHtrBOfT6wlUad/LueEv6
SUOU+cBos1J3Bp4FL/JwFGZoes52UX41to4ErKPpkqvaPZzPtC6ZWh/pEbCp0ugs
kcpjCYC46A+Lux2ReLI7Ya3VUuY9kI5tqnZ3+uyWKCMvDHc5Wmwk9BejYDWAuWcq
J00RBp/HkTqmNyw4nMEO+Eqpxx0tN+JNWwFUFOXBtmXQGXSYUC9+omD6kdiVEnJh
FnV6cKAUZqP628oTczMDWa651sO1/eh3/+CclcVrXHerBoeMRd4ueR1W2Ab0P4+N
oCmHbsLR1kN0V4LwVjK+xHITcz1sddMAw7654dk0tDQXIhQa9XlgijRoD1w0IB1A
z87DT0ij5vX+kMPGp8KJZG1widkUVstLjUJsiwg5OSkgtf6wJxuu7xw4b2Wgskb9
stS7bxsnSUdmncPnRHtJ4Xc+nXnHP+tpePJmND8M+/8EF/MbaMuDOLi5tH/Wx6TC
3aGn5Uw60edCfNgZJ90mm1TqK0Xio32FpGMUS8v509qZtMBKTW0nAC18KiG5yuSN
9G5kQjX9L8hq6d89FCM+i+IyzE0j4s7PRUtfYyH0ZxbgHSqsVPKZyqHJZWN5LbuD
0A5KubycNpHqlla+rSOZi4mQhVYlDAx5BNLS7AlG+l5Obu4+H3BHUHD/Vsqz5f9b
rGMNrEsKIOOJ6KsHH5v1W7re3A/TbEY4xV/RG40AcCN4ZySPpLqSfRNySt4w5zvC
BTeKyZESvD1NlKerB31RcdfEDfdmko5TEwRKE7DKlEJVhh6X3vE1g5o3M8iiDVR+
BUy1pEzL2g7Z09XBSuptcGFjrlReeidRGKtxCydpeoRXiIcqu1A3nZOWAQysVaVt
T4A3xYYkgXKcE/Yc0Za8uRuCwcVktckGV10JPpsj5UbBrvJCtyMiEEfSlZ+xkHDX
bYpVSgxSXaPx7yPYRulG9S0VHfg/+Qx7VrqkW/vwAskCVLNqSnCKWpxWBd4f6Wj6
Xx7EEvuA7lwenvP4rebgQR4iw8ij9QTnQln8ePPxH6NittyiWvgL1lOWq8aIR94H
Fg7TC7dR/nTVbKNu6G4Ni1aHPafIJGhilD7WjuDXhZriyEmB9egFHBLnsVI1ncAE
rzTAZ9MXNn0aUtoLCOt63ULETLoMbxb5rSLoEA90z1nCYlUbBMzSX1MiqClJJ6jk
9VZX5ZVaknipMKb1WfMZvpo0Xdu3CLWiWTHNwUWNjWx2luy/OqE9qGiFIqtCmQCF
XRM1bUI3iEzSAfv3wO2cAgoNwZB+dpnHFeo9fVSbo936D38shFRXQVe9aAmvHy4h
snY40qZLmONV/ojWUnyHICjbD2/El5MA8LOn647waPFaAWSRsjSzGbeIGSh3AuYt
pLvvB3g+xNCkXQxG9/J82NLNtZzAnCjqgmAifr5vLfk8p3RQOHabTLlHngSYejni
RHMeTeWaz4VXT0fAnZQIwRqAgzntCbxs+IEztjLtzvCVclXpEsej3vAhQyLrWzLL
YSId4VkxdBx+lJXxhuapMhR6UaYatngMBh4ZlZEuaJ4kc3R3NBrsOVYby4sHy+ut
Qk7Amk77sZWqRcKi3P1SDnO/0jAq6I5SMlT0xTDgWucd7Xe+4irYpOu/ELhF8xJd
Oug6vx/s7G8jtUlQ/YZd9C3MSvmkAf1uUcO0Pssd6KMNwmfeOala3KzZEcXMfrbZ
6JzT0mJ+l63vW91w5PhE80HqzMkPRm9/ivUaVAfbRauB6J76SS13HgDdS7AH9WMp
9iuJfyBxrz0ndN0xf3K0ct9wtAEMyocQrPfFIh7Xtf81cPs4yR6NMC2npyI4Fuw1
HHH8KYrEAfXcZ7qtMPjjIWsre2YAueqKkSU+tajCsmrEMsemK9Eb3osTKgBs/t/6
MX+wTYAFGBxYyPJAJ5r5LYaUtZ3mcMS/r8XZ3STW0ZCgPcZd4Mph55M9W/P8vd42
27leXCcLg2S5lwjrF85FHEJKuWcgUUumRPoBtL37pvSikqeDIj9gbYyc0VJEaHc/
vwUj2pj+U1+yzZMCU+1DBSV5+XAPwiZgfDQzuCV49mA28ABpcVh8z51PDDVKSbye
p9csTpkdu68x0LNaV2NyFr7ZbRLwgG4PCI4VMLh7lS8u3Ov61su4p/nx/UEe/blj
Qv7eGalAJ7Mot+z0ebtbulF/Fc0zZz+lcAey9EGLgkFwueoIwT+2alnDhc/yh64k
ywifpFANkUPqGqf3rpJcxB09W2xiwS4mdE7BZwyglWceNNMcnDS+/Zp9w9XBfYKb
stpwsrErZ1UkSSd8fzJzttgLzTVAXnzBefqhBjctOlP0jJhXxBIGwkfQlGgIixgo
1r4Zqzeh7RdGDVowtg5fr00Ql1zwSM/6dIDSmmsy0ZI5OZNYRdR0zemfv2zY8bGx
1Ct0HNbE9sV+foK2cOFEcaaUH18+lPZzQDvx/sIW64YpStJejH1uL5tievDDR745
eYvlry5CCNk2nlIraxdHKzBY+QKmcXSLZbfjBqVT+fi9Q83ZuqTvdsxyOMLugh8Z
m10vdvcs1cjO6qQrtLsgVxDI+DsKce8dc/jwVsp8KOOSv8hIBeFq5UTGkGANMaxd
KW0VcHflQxpSuQK/gnYu3b8dfIRQBPau0YZUJ+PpudWXPeJjdthRxwzZc7d+UFHL
zwFP0tgFQJeqN3IOChdqsOGK0DWG0uwOvb65VQYSpLJb6O6Wf6dXCbABcStpPE6Z
iYFO/NliULYi/rR62ETgtFAHnWryAuP+cPSj0A1gAz1bPJl/0Ozfne3VAsIiqe8q
wvs1Ab73sYGnN3ZmswKXNI3YCwXBAxy/joCG79p7vgF/fbJ3l5iaJ2jVjKrwrjiU
MO6ULj5YtkoXOMf8cMdLhCPtzeUc1Ms+B8OINedoEVAAEjwmwl38jxX1rEnU+zab
aS6I31wuy09c73rcwjegvTdMRIizIpzLdEt0DOiBbMUWqY4FRC5nticB+ctf8S6i
tV6WGaVZ27NKm16Iluh1/CJkm352nLMU70nBx3h9KoJ96zqFg9/exdflJQCpmxCd
JbgFUnnirv73nVtOcTmoTTllhYj/1d+sxtkdkYbFqd1W6oIvnwcurrrqMrCLB/rl
URggzVUjhI2MatXcUVynZlZ3odX42PUiBpo3DZ2SC+lccfOb7SoNZ23cGf737Zje
+QdKFSsg+KtBhzX4SPjJfNuAJR6aEzUztQQFmAKiBGf10g66R8jKuEGYisC7f6rz
3zb2Z8hpYVEVvZAMmpUXG8PQ1XvUf9b4Wm7/oUWxlcBEaifGygHoovqnNN3Q4nlY
OzM0IVrPM5Gh/Phvwh0+exFH4dZampS7IY+Ljf282e8p80Gpmd9mU04CD8K1+NM9
HrWK0rE/vxq6jskAkBX+ByTN6KUOmCU5jkC677vgmJdgMz24jTnXhoqT3gLezj90
WqH2wtT6iJby48LZfG3A0uaxd3xeYxMvVHUUfSSe+CcwKr+YLcXZDc7FOrHFBHHH
vDqeM1phij3nrVktGfs0kZVK4jg/ghraPLy9qSmygNKxOKZcRs3gtngxRZNCycjR
8l3Ehb2eWGU/5ja6BEoZakEyRb6Ccepxs7vWinXDTYCh+N/0RojXTTXnN3wIYE/L
9azez5Wfmgd1zyXmQJoXNs+2APUdn0hYaz7eX8HcLMxEGHxE6MxNdxDJosGgrJVj
TbL5KhcVkQjt7LvGmuW7bJx+jRrio6Ase7KDg29RWDMLEX+BtCgJ/n8u8yyj/Spd
m6u7uZiirMLTZmPSdjF3NKpNZnUhnJemcC32QzaZR+1Nc4Nc3n6VWgAM0x1X81iT
YWDPqBbjRZ6iFqoDbBPLFt642gSMIA3QchGrDVDEZWepMS0xb4KD5kGxiiLtIgrE
DL4OuQRipexgLde5DW8UUDj36kqlLn9qS8OaV8a5hreQTcv+ub0UJxvqncPLDjAC
PZnsqUDIEgzkt/5V9d8EJvZEorVFUZZY4TgXR7vJBW3WV6CftYtGLX1alhdIZU5G
ujRCZJEy4YRU489dPrHurODWTn5CwS15WVT++AE3Qxpg8HqODECOQ4pazp0UsI3A
SeOlsHWfYALySPtzHKiMOBX5kvpNuBRx7LW/I4t1jLjUqtuSvpftZTtix/PkDHaP
pZHtRDpDGLa+QAiyeF+EEzFAwFg9Sm/63nVb0I4WCqEEtiPTpI96v/pQE1M0EIkw
9cYb9K8S1GKr1r/osTdNHVN0sr+uHfiUWhTnm+2OWC+NzdjXnCD0qTLFql5+KVlC
CCarsz4pIWQeAeDq+EVmpg43KNrbT2GTbfQTqybvTFqIsAgpd0zByNywlz82LfrV
FiOQQV7Qth5yeA4Q2Byl7alxzRZmEQVCx1aXABVVt2UMnH34wN9VY9xK/jYSaJhM
U+PRtKg/ULnGesjCkyD3za712jZC9uN+NSVwxMfUSTnDzc6p225s0/dX5NUk4+2a
Ggg7HNbcsm2/2NFK4y+gMUSt3Wttz5aWxT2oE2gzp+IlUkfaQNuy1m05HGtRxAiP
M7ip44K8fuF5apjGljqOA5sKZSfs9xjoly1rGem10c44tahTTgyWQ/whe0SA86Gi
Ll0mfO3hoOFOJhWLNnVjEB2PeyfeU8+6l07IpwkIOexhCGH6jWapMdPEUZDuOEDN
04svXCc/Ob4/QmbC2y5FwDqGRke+r5fpbbEzm0iHTiQ59ESCHthl3blekQRzbYho
4byzCQE/DBiaGrp2Ci5ojkb39ESUR/2dKAN+Tlj9g/Hlvrr7wBi6tN7Q3s/0BwYH
L+nNLxHZMh2lN8Vl1BQWPduTfyNmQzQuXZ52OHoJVCJSE94DK+LQ1P5mPul4AOEf
mKaFpmjlFGXbZbD/cswKO9r1KK9wtRvPmkRP/wf2lfK8IdYl6FsPjc7OyAChpMEM
6cgyV38HoZt472WJRadWjpL3z4iLQeQgn1UeVoortEL2l2IFhsx7ORQTgfrtrH/e
otUGQTu54n5F7RF4IpwGuSoPOMTm0zDsQUsrRkQ7u75yPzHNmxLx+JcHWOtd0Q2S
nsLqbaKk2AsXnhZF4cNXoD5z142vhF4MTLST2X3wcPz0kplhWQV/Br/eIH6HyPYQ
yZ5ZJWiEzmcw8aLZeBc7tKj7SeLbdbEF62tLwQoNzCM+S9LZ/QaJNy0mGuN5f+rU
iA9oBk3pyMCX9Nvu4wm2e7MeQPrNKTjCVL1VJEPSEtKCU9Fe16EcWeyPpIW+99qp
12hPUobeJfWJqrmdmW9HF5ciuH64GGm2e167KeyqG9ADUw0pSfw1ofCOFVIVkIpA
1MuX9kFPTgl2XuArJoOQEgbbEeU1KIInXWWU81/7m4730BYpchnNBGhmzu8zBfRM
ki2PRMuVn7FKlwJu+oP2WoIwSg0AHtXzXw4G4ydBbg6HJZHPQE2jKlnqLIHBCu+s
rTiyS/fNqPK3vgWbsuPycbk+Q2ynIeTH6NP57dvpzRe8ReaTGtacpNGkE6N6DplH
nGhtJ70eM3M2QiyMGfWsz5EeMujwOcItnxPGvnYY6fHGQ2AzlnhJZJWWf8jqkA/I
rjRBjd/8z7Db7ixaJUozG0jHjfpkiPjpi+jGSiapbNttpbawgILl+Xb4bNW4HjM/
bgHqrZluzBx884DCwd7DXQDE6ruCh7D1XA92atCm/2yqYYtHJbdXFYIAODBYt6A2
Q/7FoUlTHJ3YerGFDKLuMwkbzRBQGw/DNFkUExUtbQhDYn67N7Y6D/y21BSrFbUO
ThnBc5kyZJZgHb00GeNg2oJObN9AuN0wmW8S+JV9n+YASl7w74uoRc6TM0R8FA2M
GWWPmHRFUn/Kgedt+pCXoLiYihL6KXNoN3J4MugkY7/EOKQKUQm+5hP8ks31OLuf
e12grxMKhBZUXeoC7B0L62xCR5duqFy1JnR2tV/CRjhD69FF86GxtN2wIzhvc6v0
q+8gNyWP2ZZOCuwRDm4N1pIggsFWwRFCZE+b23g2j91v54pEl889ZQjhkLu0zdHQ
UYLifRDouudroAkwfDi8YbmZXDCH6c96Qugz77uf6rjQtK290R2t/WO8uKwTSUV7
UKpiDPw1Z1ucd4fi+4rRzlo9xYFnSvKRHwPXYeDVxOWKYDUGmoSXmrJUMaQf+oxe
NjN43EwYckyIB7C96w4PMq3GZlNP28WX0rGuss6oWQwssEn6r6WwV6ypbreU8TVp
Xc0B4Tj8SCpWJBMjM5X3H7GprQYEchT4BQbItXVrDrnFHgiEtNsuVCQT8IuYA9Kj
xhRtuLOsloOLVkDmH+P3pLJtzFNDjik9lft3LdQdY/y5GWoThmeqg2mYAy3BE3J4
Hlnm52nslOpEsjYmV0Jq/6aLBCjqU81IGMN6kae0XueCpxBor0w/EeL281u0pwB/
gx3Ep7Ajprxu+pQo+OizyB/No32Ozfrvx9d0/c3yV+PS8NHI5jYs7DD4zIfIWPGW
eFWmMx4tYAUqadpqpi3u8o6y6l2+wsk/rcMJyHzXkq2oUSNxTTUjsCNoVRE2drzy
1Qpz+vDOY3lIjC0aS1N0VBbDA/AnEOHm+uQoL4Tr9qGJRYCadQe3i8qRcgNRQvdv
gLJaFpL6dm783rsPNwPU1GLlGU2TquZ569EQvF7oFAZA7vmxhAoc+ju1nel8Hi0z
cVHAwHYZxNkIzQwu2kiRk06ClRI8V+AhM+A/QnMfbE3E4EZ6cXjj8QbuJga9MrrR
gRPeKNtnzqJmM0UgznZEGzba50I1FUZtok+cr5Z7EJarVj2iK6r1zxeiOKnLrfUm
bqIDhmqy732pFdeuUe+7ryLSpiZKXI0wh9erUyvwI2AEsYLnv2oTJW1sNlBSCfaE
VJYkqgRdvzAZxsTWVglsmwPc9muG3fK/6I9fixd+/pp0fZu1vfxdgCkyS7R+AdK1
twWWLhyGRONc4z79SMttMP+FawJ3SIllNborcx2V/iKUzPG9QytNIY9+OU/DQD51
BZ7XKP5+JKwCmclXEywfHFPrmiQUSLaDy6Ysa2hRvsoDyp1dbI4mrVZ1R9Pk0dBQ
ASrM4LSrnjBtaUlyl9e1JI8egRrszWiP4CNBcEJ6n3nPCDgQ7u+ngP0x/Huwm/XB
7RtM1gs5NHkdIBG5toJFEcVDV5xoQW5yInDGT37O3oRKR6vPm3DKSZTUV1v6hFOK
+RhpIGyxu6gEk6wp/Xrkz6ZJJSQfvU9mxAgFZozq+y/PqFehfXjlBpqAyzUsFViH
HafAjJUIFhNd4WRBsDjnzeidBxSZe5oRe2TspTBxdv5IN9EVnzanjf7JGBpx5TOf
B6tznahiVtntXQrN4HqNP168pW2XqFMniC4fWKDXlIXnTXRqeRVtrrlkYmYp7kH1
jbOzrjWyKZLaFKWjrF86e2ttdeNKXXdbxQmBs46uSTBu4OEod8w2O3FvKNAXTNkG
1mLlnjYuh5+w2dPMbpDPfmv2JlZQKD5osaNZWuelVMKGJqD3a4no2h4i2SnExUSc
ZGtXymRgJlIhoRaF8UNLPLkyf4tjS/S/iOisFqJuulPwAOSAuI/d+L2IDghCuQAs
IyLUxO7HRscDSuS9NZEu9pc2qLTY9fMiKF8vaDkoAcFrLIm4YroIHCqFZtntWxS4
bWf8zXRz4xy+wgMbU83FA1nYKuXSGI0hZqe6OMAOiTBb+Yjg6A76Zv3UJutCBJHn
8P6BWdBf8YGKchb3k9NvSIf+tQa17S9BYqOp8p15T+/s2qLKed3tlWoUrnN9MZby
eqFssw6b9MrbSWOtxJs3N4YoNUeDwZsexeH/BJankZ1xoEiXNKqy1drpm5HKzJbv
qnc9lafLx3xzwoEu8bH7LafTweaWqkGNjMwqT0PYmQ4vTYpKnSK8zhtDUigDOsLW
1NDX6G6SrTivKZYGH7BeVEAZdrqjksfrJuWAtZRQO+PSuB7IHuO6ApHjBWQ+dsrP
ARWxgD0sJRYZ/H21NfoRmBA3e3P3McjnmknfR5O5/bhBmnGRGd9N0q+mes/4aidD
vaCq1Aax9w2JQhoEBcLp6QGG3t7jIvtpkCvYuuCMSbIXm/pRRRh0ksh83woxKqn9
XLP9KZVhY0VtuEFDTVa5oq4fPxpTKAMHkn7+64gDK3MJ66CyHr2Qv4r+ijNunYYN
eK0JZ1vglH74OAo+BsrQYLyByZpFbOTAX5BTEO432gaLw5IYkhtrJ+82dYlwr3GP
G1C3GD2NUmwfQJxWM57lvkcl9r/qjZFT5hBhhw0RYBoci/JHJ6lJBhUwhvEoAmzE
RmIi7i0K+mDqt0RQqnyIKusiYPt7+bMCAnG8z78aOp2MNyYbWQLXbVrCm0NQ6LIk
uCYauLIaVKcWBeZgfaaR87e0k4WG0v56eemW/86nrG6vCElF6IgQEmYdZ0JYmD7D
uBY6a8YvWwDxowbHlHzrJEg+O6d+57xtyAQYXFO1UgxeDKmKV3wykxvPjPka7Vfr
TN28jTRY0r3/nVmCUo7UEkq14Fy52sb4Xmh4da0vYaj1/cV6XKIOoV174Ngbz1LM
d/DC7Ndj/vlqTeme3nxCfU19KAlQJX1UtxAGAn2XRjGiMudHm4mVHJVgEoGjBDoY
prbeZetgsC2x/qjqY4VO37Pyj/qEjqPDGr+5UZ0U8NJC0p18JMM79iNfZa88ZfEo
8z/YnCoPHBk8k7SEnJ5ArMr7YU2Cke4bxBGtImARVJxbzQ4sqF/R6BBiWqnfQXbY
Q6ZnduJCuAZIGMpjEDmrs3vmPhNsIYrCmJROreFVthBUtrvjYnajRMGiLijj7S1W
i9eaqAdCBrTsVYCnK9jE+e9wemdZMyMDdZiD/F4quHP4nSbD28VdELwB/GGYOcdz
J/355ZiIOjmBCmeH9XeZIKO8kVgA/2BcK50PlcS8eiN/X3h+XlTgJD/xd2xpSFg8
K9to+nY1JVpiKOybWplbwJq7LKx2c1pPJx/Nhlb/nAwqw86qaAi+V8IGAni0Gdua
ZBgrg7RXoegq7lvxIpZ+jDDQd9v0ziJrkDhLsF9q2aS3Dd0DQcQBpy3AkZzjZ8he
5EJbde8ArIdCIWdKfmRlUbvyvhT4x1JQWlRnuLd0IzCWPfIjC+5/bjs7nln/ZJ0o
SB3fa0QljqCshztWPszmFYUWlGk/Kho2MOm7Yr5fTgW9UI6PE7kopFSGtBKV1Jh8
uDazQoJkxj7D0j5K2TCcIixfg8bJvgDejuiWNf4jVNZBTwJyftCAUlytaZxieiXv
Dw9kVrcNwFB6TqpestePAFM9dQiSI+QWRBzzynBiAwC6cfb2IEuockgn/Ns7sbAd
2QMI6jV/8VhrSzHlCBQ/APGhUDf34AnUT4Ur+yPPAdqvP57gZSXN7dWp6GCejpCm
/OneQAChtGWlrK5bf1T1wFBBysf/3hgYu174x16a0/4vaCdPeEGeWpxWU9E9okPK
rKNf7mBAvfNBmr9wIRwyzLshIkDO1ezZi4H/9H0CrANKCLZaPEACAa9tj5ji5TiM
4L7VudBwzuZNaZmWJaPs7L0/MG+a8QXWj1G/642jAsekWmGhEZIkJFP/cpOHETqF
Q5f2en9WZAnI5lLMGZzVIB8UUrQVxaWQhMdWdkO9hyH66d4y11w9vDuMA6khUkmH
izEhZX5/ablwNgfcK5I5YiNyxJA2NUAE4Zt58TLdVFSAUbQ6PU9DFDXoc3+/Pwlm
uSw9/jNcaD7zOdfTbrtZzryFF7vC+9uSFJQW21c+hg1/3HwWEw60WVOYX0C7t0kO
iZAVfWr6bHxKGVkaD3rDfkiLbC7PqF2qYzwBlyBhzIgh6/oPLMSvxmVRoGunAdo1
NfViblsVrR+u77exWVYDkTnBEI6/5pcwCdBzuYz4Aorz4NEzK975RNb59ZpWmUg/
4+0ZG/1cphPPu8i4f/aHkuUdJ4kZvFljgQYdurXAbKWPe4F13XBJ9BL3zUfPtZHf
JA2vw2SVwxjBDC5mpmDsvA1RQTbYhrDJR0NcNFu1QdFoKw/m5Wy1Wr1A37EnLYy/
aOdDP1bYhUuUrFBFN60hmlDXWmcK3moqqwT9WyZ2WIEy1Br5jHBAOqJWqj3Qolkj
vCDKAeXVydGifNo3fzHOIMyxfAvTZmPEHHVMl/8Znw5unU9P0Q9YSNamEGwa/IaE
um2LQZTCaOBWOLdfnxm8thzsKReqy6kxO2tD9+mmhU2xWURLerqLUdIF0khGY+Jg
Y20Tv4bzkJiQuWKrzTl5aSQHhW4Eex0d8oY6Bk6CpyiZIDchqmoM9tCQHrZPc3qU
d3DsMYtygFHj9SEnKhHXQvFrYOB/ao656+ElSFHu3F6lcOa2Hcl8DByPyNkUTkTJ
Mm1B/c2akzkfP1QP/J7ZoGl6UCO7Rlmx2rJaNWxroFLghSUpD2l7FB86B2dYv8eZ
k9wzqOrydBxjOlLm4MhNHk2hNM1LbG46B+Zu6qCNyhkWQHqrz/D4YYKHa1eG1lpK
w60aYueuQ62PWNlTp93K5wKMcOpwdid9kxehONKgJS8k7X4t1lLme0adnYTqXymN
2fdT4lGHox/JeZQg7RT1gV4uvduJW2Vx6D3Z0S/DTjIo5A8HzhENQqzFlWwr+OWw
Y2fnAV1bLh0FHdZgx45/UgbWt3PQS7YxjYKwtKk8bQ6s+HlDAYX427FR2S5lBmAV
a9CFiEXeT47yNRqwPDTF4n+Ql5bHACEbertLxdYSH4P0G57N/p7WvMBTOoXndKoK
XjCPcyYWAMMht1+Ho+R2NAE9RA7Pxjsvep2M8ABtQCZkTydBVuaA1uPyyVrYVnLB
TurzM/tpU94VXedA+29DqiBQmPOuQSdNQgG316bQDws3XjrxmqTBDLr7xqCoYoqS
7CfnRmJvyn1bVLylYNtmv9c0C1tBvz+HagL3varpBRe1fQLQrV8DBwZfUCf6XU+Q
tJoyVcWKbOFxoguBJePrEouTYNEFwv6VSgmBBc9fJTqgG9f3X20qumrQepznr5U2
yVYuDziJX4CP6c+bFQ+7DDcn3atNGewmaZcNS8eFhTdyTG1tfGPBO/mEf0m4iLps
dEau6NZVfB67/ygxVG+i5iLi8IDd2zjXbmLHcS5a7KvNxQP5BxlVNecB2euixXt/
lEIyYdJenH+vjRnsPXQKk7v7R3Fx3bZlRy7aO6JIGhN93DP9+qFiyshronK7wqR/
97qs7xjs6+1j9vYIWUhPyi58MO9wp+EtuhGrvzRX/VWsTINS3gWxYb6aqv8t0h/+
zOhcjUQzJttB4QkT2KZ+Rql6vilgOYUa313CGeQcAy59fmqBuDgw3jAsN83QkMRo
pJBc+3KRNv3wOYh8mlM5CAUf6rf895EeUg7qCm5hoWB8u95cbJUtIampnFGrpDne
4SaCm4WCsOBPAbMxcKpMOZS7UUfVYLH+N2rpvixGk7aYnhmSFpVSt35ZP9JxSxbv
qRSdQYYVqbm4YE9B2bDzSXijCFuWdTdXy1WLI66PHjV+W3F1kZE35zDoYa/x5EYJ
d+XPzf2PnZ8Csnzaelzxqlo0iA1iMofnEAs0FSj7jGVqkZfe9q65I6iOjd9zq7xw
xHcmDfvDwqzUDdhZvOtXHWu8lVcAQus4dHBaKPaY2uNihtV3eiPcSE/3C33bQFQK
L4xAEmR6Mm2TSPJmY4fzhfhzJmGRloce0VdONha8heGL5Ajk41OPBk5eb6AvJXPg
NlaTMwWnm/afQ4EFvo+cL7wzDwbQtN5giW/GkfkJvzBZqSQWgja9KvSRGj/kJ5Pz
l8VFiJJLCrzTgC6PgQLpUNm+sHmMqO7YCqDczaNnjUrRQ4wmDhWSTKVnUM9+yqNe
orgUpBOSDnrg7eSkMLEH9r3nWMwnjAnNYFOvw9ZBd6Rhz/6cfh2vQIlKVnypHEmd
LppE4FFJiJoDzlwrqsuF3I2acEClkw2RmH8JFWjt6dz3HNIeBwe7WLwG5hBGE5/t
K0evOdBe5Rh+vFT4wv2wvQQ7QQyaWjQnzMsKzPQQRtX1fR/XzaabfLey1mVmyT3H
RNqaYwxcvyw/98f2FrCQJSRnR9pOOkjcSwWHyMrETstVTTh70JVVcRN/+ajwrJNi
/g9cm1HFFQCrXIKZtXd6/MO6k5ox/S9/K62ceL7Q5RGqxMBztZtaJHLvg4882v+P
lvxaPnUrF69M/od+YUw+O9ua7J6zAjLsdTZZrEy3zWfV60oEfrBnR3Y3URKE9P3Y
xmU/9f2KGzDNl7UHrnULM+qJOUxDlnPvXolskofVE8saA+7N2orx7DbRb9uW3RYK
GR5fB9CSAiIbFAYE7pUQEk1mEekDMuYY8LtPqGTQqBylx443CW8g3+0qg6OQoNqH
EwZQCHi4ainVBrnyqqVaGtSEcgNOB4QLgKcEKZ1dlKbrib8th7ORUJvKNy1Q/EFz
jwtHuWmWbMwzsNZM85VCgcIVY+oOI4frTb+RoBKlXOwANxo9TRPEbwP8ko+K47G3
bx7wfVRVCSqgVd/szA5hmZ4zKaR1Q5TZGAYffX8wnogsoUxRbDM/egMi329rAbek
OK7qiu+2TZ5d6hB22Q0Emv2npCh3kLMHNqizjNKpT2wnSAoGZd4XmC35xoEO6WNg
JMGeQFc31EQoFPdG74UWzb9i1C5vR/X+rRUietNJ21Kl29sX1NsAMt7LGR7AAorB
0cEvn1CVDR0bUb4encfkXhjYo5zSJ7RwmL3kmhzn1gddCB44/kEUfjtU+jnbHNAW
QZf/8D4oqyt/s7D1sq3FdSs0lyWYQphwLd+hlz+991rF8HbPKRWGSY7dWY1lkCog
O9h0mLH5xK8jZ36XnZ/3liVECECS4VGDk0ibKexoIQ4mBbHdcEAQijeqjGcLGbGW
FhW4aOfmb9QaTpRuqRZQq0j1TtjPpIO05R6nkfZ63ouGIzmzj3ty5k+PoeQaOYrZ
jadieVZhImuiFyb8AjN2BJrSF5nMRvQIdDHm2J+omDCWZC+5Y6By3X13VJRAi2aE
qr3Zsw0IQL47RSIY+EbO0R/jE6HImFB67AMyCPS9GzlC7gRZCuAi0J5os5+Xebq4
7r9+KlNyS1y6TzQBCgkHsYKAfnfaoG3+lBLM6Z8tSxG0pycE+2mBlD2yvvKRJrHh
Y0FWJud+KaKG8fC60WjWj2CfAvdEDiIKeWCbCQZjYxRyI2w+1JoJKhLkNmRsvonx
jXiag12VIYAnsZUNrIZ2lbyreriNwm5ZiEWavhAXAD8fustYk5f7SwwAxsBctVzo
6IgQWZ+J9unRKnbjWSwgHTx3ygmVSVu+mowkHZ72XHrFXfCwG13t0fc0b+yDItRd
iMmKBjn3NawG1oJ2zHrDu0yq39jkBVw7r9DIeZpNX2U+huQMppw7c423dlPtjuRV
S1tSIm/6V8gM21YdeWBxQCi1GWZMReQ4Y2nfUnkC1SflFJaxWuavF9z0Y9kFGi13
CsYnVFN/Gaw46nrsqp6JqMWD0Zn1H4eb4QErM2XFprPDPiz1DF7oCAZmpjCY+8uI
vm/qAzIFP8bN/+gfl6sWT67f9UhhaZwyqi26XXvnQX3JJHYapRehrg5MFQQyvR3m
TJG4n62qeT9HQIIdiDTCASo7W7c+kM325rLKDmCLWlC1zudS4i1EzihuMctNLOrG
bSZ4nP7VHGA8d9bsBo1mPWOYOAF2N/xNZka3ApzDpUy+J7LJ+WKG5B5dcKWpEar9
rBW4bejIPJvbdSetXWttouH6pyi6wHgsW3CjlgRKmAJ3vFfafmq6bHtiP28/JT++
j1/8YuWrS8PVqs7yMZVihB160HMctcutLhuL3wsy68ZXaOENr9HlE66LirOwSOYW
GXe09xqoI6W8S4I1h+rCWqQgIfrPmB7Weg3et3HTZoxrjiEjoTXQBgIQ9CQwhECC
YRW8Ee7wCKzC7xsojvPqMihpizT90OeJ5fQL1v5WPlyZHOzyDGnickjKtOeTFGws
y+Ei2Dxg9wMDHGOQTx8n2DxGDSSQji/Ux2/x5Lq3vNPJR9wWUeGFUq3Y65N/5UZ/
3clkSYrvAJ+lPwpfypz6XxAVeZuuo9yX64BeeJQG7q5lRDuT6yHdxGBMDP8t7h+2
0d1LrM77zHe7BlJ7jvVoESNKWKzdUYB9BqxgX/k3Elh4/BQnjHVCyT32e7Dew+z4
3qieRXf6HMBmFYaJvhR7H5edEreg+HZzmFm8qN9X/AVBkBjDNg3Sisce+XM1YBmQ
IkTeKko/S3U3ds3QcxJrI4SODvtMFx9HcWb3xweFBYnoug60RyqmLPFAGvW6HUt/
xKz0Gu8tFRSD+eTvsbOnndGNJ2lvw6NRE8VeVvPXVGAuItT6J1nJ+j34C1DKHG0p
aFjqF68ZNfdhDpafDGg01ZJKBx5lpp86ptzmBurjMZ4F03dooso5FfIfXWrP19nN
kg1NEo/I/T4PLb5e8ypinjKHiYDEr5vayUcjntBrxYyqSTZ0tq40sDEfJIwPHyMz
FZ66htLSdKO3pvzFRMbuPsotkO5nyp3Afrl5Ay2c+t4YeZBEcqceOOFItE8dPzHo
/I41gd+apirRQM8VB5hiDSlLCC1/CoYF5TxrZ1jqx9DeBaYla0Jgs5zKDEF8FXAx
EYeGqT7FaMUZMLEdoJ8KrgDzKicMFx68LPkEnoPbPq0Yki8YOiideSNQ9tgkNmUg
xiw9DRp/R3gVcAo0JQRfpVN41rY6i0xuv0oUI5bZqRwanUjusvKAhMc20f/iS4Jb
wcfkwa01dH558I4xYA+2kpRlvEgHxWfDnFyHWohVkrfzCSF28RCDpo/x6zqDHhr7
l19GoDC3riR0fHcBUzhAUAUJHW4hI4azgodOg6XIqHOZ3OP4PdJXGcrVXPkwxOOA
BE9RV6HW+/jRtgY2W+AbTBXAwreAY2/NlI3th4pq7d2pSjrThvRK0ZEibcbhdmLS
fu+q5a6/lBn+CdU4ZpTeSh/EWkbMSr13Vpef3rIhks4ILMh2GfdZLS0FWTOSakbl
ShaD7Ri17JODD7Fo9Qf3EVW3NGhZeApEwVZMM0E77xGYUp0iN57ZpwSAJifZqVMf
FPY9LkbCyUVGeSdXHl4BnnE8qnVyd0xH7VX5G47nPJSP7Z3DI/kePyt8PoyYaTuD
ZDRofmKYQii+QwwIEZtgwybDfqsQDYh7egNvJ6vcC0Mn9ZsK80xaF156aS9gAk0z
76UNZo9EX5zd9LUhR2ey2gtMJeWejYUnUsUWL9Az4DQg2gIWKoPsg/BQEoyRbDp3
CuSD/QbnM/v7HVKanZXGg/br7U/J/VvbCZLSkwcsqmp9jW7eK73hwWCVAET/8Isg
JaSDPu4Tmk87yQI9EV61z29IUggOaKtws/ccyn99P2zzPMrGJJ2lmZ19AbDDkpBv
ohcHWX9G9imWdn7paIxPrm2rJkVMqgn5xoDfAcsUDI1EKe7owpw30t4LUjWU4y+N
sp08CC3XkLmiPfaSoS3W1Q7V7p/kBsE1ZsudkvalFOdH3ubOA+FFngMJQQJJZ+0w
ukafRn8Sc3gNX2U0GBOcFQpuKhtiNPYS6Ah4rdoJ1tr30AeZ+W3ALCh+fgRgeQus
K3cdjbqSGnEuB0M6CAYj6ofJZuCvPnr6Uvey4IwB0raQa0fVC60KjT+sxwiot53k
kHY3mcOkL8Pb1mcrSNXyRd0Ym2Qkt0nxnDjipNrkH+VFk68xpo9TdAuXqmEyszfh
g7Gng6/YiGWMblY1dzZCrgNkP9JRjzGB5SiX47gOedlvtsszul/1fiwmmcfhUGFi
LsjcnzpJqOiPWEOx5N6/bm/aSJ9uLD/iuU0ybmLCcuNzxvnLGdEvxaukn3JT0lK+
OZUKAYqw0ktMweDFmS+ZVwF1RnaAzRrmKMN48IKABmHjgXFYC8VvQTHutfFPW5QV
x8KCUv8HFnf3GMuonE4UbR55JoH5Wegk8j5A65Dca+Rq4AhxEvXbfOhF5KacRO9v
9VqLF7TOwD4qlTG9rxNGc92tZextASIA1vv/KWDT22EaFmF2cF+5UjLWQKjN6IOG
3ILst3Bp/gGUcrNEOf2oq8vBbtIk8JEG7S21pMsuHYAzC5bUte/XGbWSD8WDNe4w
FXwqMDtAVVo2vO9eyMOemJl0zYWHzkYVFYbd41qpwAuyxcAbYzmwBpj6/19bbso6
fbubNjjDy2a1pjKlq19C9YW4u04zfZ8mYTYXEySeW82hAoJXG5upDWL9Y6oCLyHQ
cTm+yFvSaP1TMS8OG5M4MNDUHkxCzpmMArX3MkHxeDwyLQf7O06Czx/bsYKikI40
qUIXLFcXKIgp39Lxy1nJ0+CfhkdgUdSC8TinsqV9mmyvkjU8g4n1WTUvvhI9NUKu
sMqPCJNcq7BUa4s91BGud6eTOR5biFmTMjpn7iMj5eE5ciD1K8HWyX80+gzItDxr
wB2gzN2cbX133juyLT2GCKf1WYVcNLHSgf3xFrONAmk5XrzYme5PP8TDDOCoRhpb
4DKcPOG5mq7QogDiL/1zmgDyX2blLIK/ISCmzNmPTZm7Hfbl77LO8NLx7xKi8Iti
2Af3dg/Odh44VORZKBIq+V5j6GD+JAITt9/0mGAQbuUtJJ3tuq3oL8XLBsvRgXIp
kBq2u7KJwYUJvyukE8rkySBNIu/NTyDAYvXIhPyFm56OSnpffHg1zx5gdkDVn8mq
0W2I/UiKT4BJXNn4NIdoJZH91a9PJpFF012UQZYsMqDH2cxzg4ej/xTuWP4EoRTb
0n1/G275IH8dBb/mCJihV/ebQbXd070zU+b2K5Gaj0vk1Qk4i4YcHqpZV49mADsA
AkQMGIATPyvhCI620J+D8eoVxnR/OH0/aBHyORgbLWD4bPs9zhec6/iSin8hie6E
MoUO8FtX5zmO+f8q9HilUuujJwvKae9eW908L81nVjDABaXeYLZTG2RUdYxBRljg
JaU2F+RoD/4AZpJiFk7YDIrcQOO5ngR21eheupJOqXYCy/MXrgIursP8zFIvdwc/
MGW+6DqP34jp9e+mFYMvdoRLK5UDszVEbOjPipAR8n8In9knEsugXKFf8R8Ospvt
xsztSXSRfJo2vBKDDVvBIXFL+OMn3t6Ap8VPws+wqb4dVKX2ZOxDbiHN6E0z3A03
X/SLv1mJq9AdYjAbqgcV5kxN+1LW+3JevEa+7qcqXhtUbFlpEFnvKJrMghialTl7
Q/xyWxalxanyu4KXc2U7Fa4lJOdUeAO60AvJN3hC9pRsgA3cv/+cpOd4Il0X6iHk
zySxSA/nstQcabK3e711COiMsUxGW5czZV7RizTgfIstroehQV89bMAqj1+Wb/AZ
plxz9ebsw7hwGmhQyA4aUNEvPYA1aoz8yOrFfB6l1phzij7Jl+rpyZhbzaO10N5u
8fb45ssMkuOw/fAnVxCEL2GoN1FJikOB6Y56Am/RfEN1VmMwzXQeiWl0sYeMNGeD
Ioj79zHVtQWCOMoTizm/hhDg4d9nol0Ws7GDSatZlv8SI0ye/YBawYw+euhhjn00
1HCY7FtoSTaeLH6xd7LaFRbQNs8v5Kon0J7esqdZhRKryHqJ3tMyFRGedM/i9eN2
eo5sn5RMOk9iLNv+mmek7ZeHIQP8ANnkN/ji37ogBVnfvKULce+ilmElP9SYmEwz
PCyeqacIhe0ddnqLYQr9W++jqeZOHOs7vfTe9ouNNulYhcVws9HuWS+MRn8udGvM
qyTL5whj95b6rmQkWYDOfvMIdAxQ8wMucDRD+xGzCfd7Oog49lwq8DcQoqp7bdUl
wyQrpQynUpuSds5prOPqRAllJ4nS9nsINfhdqTW+R0XqQxLHFSjT5B+XSORVNOvd
J5HiHPKKdRamiLOaSaqEBBHsRw4fCzVL8b1VPEkRm8g5fsCdixGWKDxJSUTY4P3o
ngSFHOQwGP4X7iwBi1xYxbUD3jWSAgT+kjEXhqjttUaS5xICv1ms5hyt1t9TMtEQ
fGyqZyd9Jw1nctnT+M3sw7UhNX3s81BgiT2NN2ioX0jU4K/s6OrqJf0fguQ65RSn
fhT/+AXd406IEEBHFCT9oQryT+rbJIJc/m23ftW8QtMuW6nht55yXF5/KAbmwKgg
UgOagCTbdgqhaLoDK+UruMUnJBM/2ohpR7xLqrL7Sl3f1+7ppgbPpeYPouA54ods
/ZQkFo1aLw1p3oan8GVkP2bSP3F7bw3hcNvp5L4uzBF2JmUZCRAfNCVChGseFPF0
AXyXZwvGyflfwPypLVqUK1klMjf2JYHGl/95xVI2sO0QEA2wmHCvXyTZXxLM0rHU
o0q6Ibqh+9UJP6l3TNCfkrbBap3uyakrBSSsMOHHhOyAF40r+jrpOAfpyfzg3utg
T2iD843nqGtMins5YY6SUuGxByvrUR7UFnacfVD8O5z/7g5IdzIUuIRIIC8SHbZT
Ff/l6aas1QaWddWfomZms35sFIPK9hGtBv1SZWZkKlPS0YEFKruvpZWGJ3yNIerL
GXqeiIbWxHLYIGg0X57dQRlLKoCUd9LZ3q8OqXsLmqq044SF5X1ld9mGyOclXAQG
UX/eC2W7OBYi1D0eVxQH60qMVyxFaVBICJJKt6aooHOAc4pt9xG8n7ZmJskaJjNI
OMLKPblQS11lnKo6kBsYiD+vAVly11vMU/ijDrX+CF4bCuCqJTiz8FDVQLGN603L
Ze46kr5lXmopwz5Ru2KJYLLV84injbpsxrrSLN4bDEbmxEGEZb2Ghyvluge7cEYW
1iIS8NmJaNQTGaw6qqpOt1iGdsA/n8ZytkRk6iUV1BT6Mnh0PDzB++UZXk64IM3O
6ufg/s2g75y+f8S6+sHnV3ud7CCElAVEMPpEt8oeCOnxhRgaFIy/z2Qfa5x1nFpW
eWxJmyM2eoxOpUdxuLP1LMFPZDM6BHXwhOWOg4m41KHpAwiPplwTO8eSRp2tpxZD
E2eElw56OnAqoK+/BeasnM3N+PfN0SfBTshACBRlU+K5tm1+a3orAkCkHfvn1eGI
iFcHfnQ70Y2DUxn1sqoE3vbCxygM5bHGYeU9zRuXagabydCFhwLq7bkRthY5iH/3
2Qw8pNmnGFqEd7ekYtq4H1pHw0cN+K2Vs0T8b9lZ8EK0QIHG+KHLy22Ncp1YuCE7
x2WdmWFWxwFtZNSqBz/eCFwa88I6GqqTjS9IXfdNYji1QbqZ2d5fun/a+VbKfOJl
wL/xn1HfhQiVT7+rn3ZDiaQ9o2vORxc5ao/GWGEbR5caBmD6dG0a86h4WEw/KEQ0
d46tc9Y2N2CwZ/YICKjDhymR3wq9uuL5GOWQmwr4vYh7V8A9UaIlemWBfnG8Fm8V
vP+dwAr6xZVYK35sxEd3Hlw2I/huoruk6UxTew1URUyiaAARHOS/LdxjKwCwkbuC
Qsd3/nB40LzG+zjrBR+XHAJXyiyfvMiOVt52WAGQXmIcJkxf09F+uslgNao6n6Q/
fMqTPmQBJX8FuuQB17JdfCFjz8X+XZcKnWbHB86GpMYnqn8MJk9hTalZBthx0dTo
ot5d+SvlbrPvzcfBs+CwmknVLAd5slYJsJbNOoAlQ1363buF1/rboUZ+TyE5smZS
kZHKnKpBZILMBPwpbNGv+ODn9O/Vw2/rVdX2bOw2muljh0XcMamCPnBaAab3qaQ5
DG5z5Z2LYDwO8HBUXkLUbH5+oEGTtXpd8snVSkptnsRvH37g4Euiwbl3jhygNxTl
DyDNW6hqT5siKuix+Kt5i0DnhxtnBif2SFS6iTHUs8uV8dAp8C94LfeKhQVMXq5r
aFOmedEtyMr67EVcU4KMd62VR7J5GOjOi6BJWZggD9vF7JfDNdnwloQoK15x2ZmT
yVPJbJ/OBiPo0ydvyvSwPH51/7NMrapLMJ/08ZzOh4Ffer2uykCSoT8Ltxc6tbiW
9xHbVv7tValBynRIdKSm7M+BihJY/ulEOwsBxmc2QZ2BoFKYP6yFUhUSoB7rpjVB
kzxTcwgek+buDnt+stN5VhFdr+msAqWUHBnwsTW6mQCH8eCuKUg7DsoeGsEqEyPK
1UwkwagowuroSNrEaLPEh0j5sQVlizoZV92SaEAH9BsemoEuapqS+oVYI5m62VSw
u7I6pnZlMz+ltsEt0jh/dDFWyQ5pctrbsaJQJaMwljiKvPWZvgPCiFHtMUr1EjSb
CAy69lzKFcixEDYGVrtBJWaQ3f6061EzF5ywTInxU6vzEI9yzvpJ+0ztOzA+Utfe
DVS0XAbs7lUrBDoSZ+nP0ofz2M13vME+9g2YrKLLFnlEz03uTdHcwAJJW2LT0SiJ
i5it3DDHYPTcrsNQRjAkt23vCuFY7TcyjZOGzH6kFAGGEx8FBx3bunPhslch04p8
wvRBKp//vXXb4zxG71xCZuA7y1mceeKzzKpo2Pv0TS3PLafQRX3bIh+98zPWmbVb
e/9ZxxTkr7QXd/rYoanIkmTT4DG74poxMDeW4J0m+WrnfNeusj1Hdwt23CCWuVEl
qOTbMLJhxjbxG+aoJZSN/xLrN+0DaSxesZrTB/SB/1g4t3PMMaRmvOALd+S/ieY+
W/d/iPqmtI3q79WXMwq325DCK1mDWWKKY2LUhT4InQmmbLX1+gdAQR7ReJGIcUPb
v8uY35xlYzdhc288v2YjgnNGa1rxJwowyK2Ctrv1m74eFgKMNwcrozzJa+ru7wVi
SIP4ROgcHljRRu6zjVax72L+CB57+rsrUtuK7PMuk6Snljppkx/v4oPls0DLdMRe
y9Ku52+K2gTOOeovr3Ie4gUvR7P3c7ab70T0jzUY/nu6MxCZIUos64/9sR4pT2W8
LKOwGHTzprVI6clvii9xJf4nOpyy/4p5Dra754vxCTb6uTWdlE+uoGIOaruVypWC
MSMNeNtk4ACIS9S0kBd0EWv7ee+2r3Y33pZNl7ebLEDz5wbt8mM/v9Y6ERf4zBqm
IL3qyN5e0dSTDP3JtFPSd+jRJMoJUwAQEt4e983JLb/nf9se+DLJw7QwbvIvZidQ
disA7U1oUYNgUWHy7ywu2eWeJljdwXvI7rq17N1Pr7QLkMhmc22BDm1An1oWEeTa
xrrw0kkQPr4xvaxr0Gyms19iOfF3BcTqUMwcSfHviHczTZ3DmL/EbdvPInQ0y1jK
LTn17JYnHDtlGl2MH6cLxH3ce7NuoEdc882LNJezdUM7ATpqUYEWahKyWwh6aVjY
OCJzmemKHq6iYyBt56y2O8SxMtV70czYoT9l5EI/2rZz8L9ii8XutJMUv/T/qHA1
OsQQO3o0iqeQjP2e94MLxsLUh/GvxILcg5tRf3ZLe5zNEXjMlen9hbZjIh9Kuf/l
lDmaBepJkPPFwJEcV/yiRl0qx21gB2Go79NYOFhoLDBmUnONkgzIXxqg0NKDAB3u
8ZjZNaC4WGXaRVFprrMjhxmuc9Ds/6nIPgnxxgRHqC8E6sPfM04GR6Spcb2+Kjb1
NLNy3t/JcpMLnRAeMu3I79C/w4v+j1XkquBaZdzotbHjNEvSqtmCkCOaZHsO2mRg
NeQZa0tax2UKSejmILJpng4W3q657+kLetmwDcZAaRc+EXjShl66fuzNQRQVpj72
19KYjf8POqiYdmfxbj6yUmcY2PppypVlQ3fvRtMbzwlhX6YHiR3ZJtLobLCovVnM
YBOG0RG0LdYvMoHzwGPmZNj4tltkw2ZktzWgXF/F+IsNofittqlsbL/7ybV8bG/7
rsxMiMw1xJZeO5keXZ9QxKRNHR8KXViHEHifjBOGXLGMqJFnIxVFYFmEACEtk0gD
u/2opmopwB5IRmbNFUz4gD1CA6ABtyfikgyiIEXAvpD43tYoLbn9W3k1bo+adjgk
K0778jevDjSQ5DCxw8e4gxk+u7IqBw1pp8PDY6NqPyysUPznln2bMXk8hEs+QgTb
b5fxMZpCZa0gCTT4SY9+MucPzi/LhRNcBMQxoLJyLdX38pIqquApPvRQVQA4Sgrk
C7r5HERi1QjgLXvpOXFSRXIOUTPdl1AmLv9eMz5Ij3R6KvSrops1UQ//4LzMZKnZ
/vUF0NUfwc1pELzJW9LF91Yt1FO71ki3SutA24Puo61UwslT3pDHV44TQoqRsfid
F9NgWn5YW7BArxYgtbPNcMHKmSBwxj/6+53g8+HnZatL5vO0taC3ZVdG1ulzQyGw
21wippXdgpG3d4G3zedLxA13T4QvnbSFa5Psw3F5QrZ1K46Yy9FRIu2ZEEwNe8NU
mUFvnlWddERuFLjM0kIA719ASsnz4zKdqZvrEmNcau0azwfYTH6LUTZgrCHFv5lX
yRR6A7y65si7AnYKHEqlccs8WLWCLGCXlfm66ShKzsgo49k38BZVYsBZgEUNX/LW
gZlrL2+015vSiZWHuH5lLaA29tKcMq3nqkgcM+CsWw8W8U7px0PlEcZ0n07VEV3J
qpdj3UwesvM5nTnYMqYUOD9zH+n8rnKWJTjpuUNb9FNEAcrRtFfRdbOmw61hNvyC
NnWmFD3iOFuFvA7ALWIYRIN0MIhlk2+prZXFPemoZDhevunfTASjMYeioF0sbgc7
19aWGQ2cTPydgYfT7u6iZMRxhyJTR+5SPLl07hGxHpFxMKwjmGp5CtHUCD78M3Dp
EVOhvSKJ7v05whOhQadqEfRf5IzI+cxrdlhHFoxipBvWBJT0/j37g//j22vpOQWe
Qc9yRl3Qxk2Y0TFbjlUVNK6XKQvL4je8N32zll7QqUUOGwaz+5qAtr/jaCBT2egC
/mw6x8+/nOTz8BCJoZtA/QkasQBJarLwocRN0FJStPk0Gjs0U9hfScee8ISPGGuW
YTqZ6MvJfxwkyQHd4BKhvTzN7Ua+NMqhMFfwqubhJp8hd4QJLmQ+6yeMMVp52GXz
8s3ieyak4Psec5hoHXGhuE2sV5ExIg9VvHJhF0ljMx6ktTJIHhra8C0b6yNyV9bj
GuB9/dAwykMrkWwiDQxyr661eiuo8/5tsfxgpha1fyKz5n6RixT4o4LjnYgvxT73
pDZrSx5Z1fCZ3XztaUh9mpcrc7FakfRIaxO/I7Tiob+Geb0hkcJ3IJ7gUx4agUDE
oGjmB9/Ca6M3jfEpObrc7b94eRlDLPJhCWlRH9Tgd3yERMuFiARSL6YEtL6XaARX
5eYHe8IAdMy1vEBAkwlVVXlmLMtkGQBRItXYVckqeV9E5DrnJrCrHxdvje8ZiKT7
FcSIqsZSF2+8dhyO/FdsoRLJOqq/f8A3Ty340//O5t41iRSCYxsplR934AynGmI8
jt15Uv+8ZboMunl0zTX7Gt/MxJVdPrzFrSBeaTfBLEEPcYo5p3M9C5zmZqI9mLe5
huXTFnDNmwpg9s3nPp1vuQecEz1n8OSea5ANyn/06qYaBxsvJFPHsiY7hasb6SaE
BgVnyUeqeExGW2atSs8ojyYOavTgBrON9/4BCm4DcFvw5LYXfSqO9OTDJtU57dEz
vcJkjBQXkZ0G+IDK83RtEcoyrsVtdae9oZoSAXlGXgM4he1i8OAmGre+YQCZpmbZ
tc5SxcTCWWmdNgZcQ6vuy+2wjw0mPEtSVvQHqm5j3ku5pD6lVFUDIdb1PuVfcEys
DLNLSR+EVQ5tWEYUmunWhpoJmxFBvXHMDOmsONoEAt3+qc+XESP54U8wqbBNCXxM
hn4ez54CEmjgAfPFu20AbcWb/48FojPjUu16c+6SGYq+2/cKIgOZ7WX4Vll273ZV
k66twigaTSBncIjqA9STwfbue9SsB+xLVoDG8vjJ55PWxQ24Txpy8Dj+m6uWT26S
QX3NODZsBc9pmrAoli4OWvsuL1Kk2034+oCzdaXVmYQZ6W4Im+6F4wZ0DOovI08X
G/3GDwD8ohi1b2fFBLngHTsl/9+f49Fr/QrB7Z0jFnQjdeoiLmzI8CeRVMGy/vL2
tz3LxWMO7mSZHc5IAvAx8IPx5WNvWjtmkBIK8iELuFzLLbh1eso7t9RAzEEIz9ol
zIQSU00aU6lvoqny51s2TpwWmaKy6bPk8OSubqtrK7q4dN4KfBa+nY40Qt87EEVv
lpNJKZpgRRmpaml6Tze6I9IFrw1/Cz7pOoDdUZD/oQ1JL9G6iAbmsAdinMspeS+e
LKqNboXQhvWL6wVTtcRBl+0JznX4IuFcSqO7myvRfO07XStwGbCHZjBP7XTU7tPh
7ldcaJ899Vu54vViDqKvWT24KgzAozzJuaNHdiIL7XhGCZI/XB7GYNn7D/MbKtzq
uTco2bXcsyNJgF0WCGYgxJxYrZJUVCJsir4VhDCFL4p24Kjjy67mmtqdmivKuqU6
FQwv3IVY5S0R3R+sFYdNTqHfdpNNjGwPz5Ns6gItvtanE/YTfvXYFtLfV50y7ZHc
cvc6ko7qxGNq+3AzUhVx+h3VSq1MpG5UQ93tKAmINaT/3iODA+k026oGlevZre3q
64hKQWcMS6Y800mETIJ/mC+e+ZlOIaqg//617uEPxcZ8Hagd/kYURJrudIuSbFZv
Sh7Fr3/bUELLjplaX5bd1wMh2qZ34QvkiAc9qxF46g80j84XaAcKnHcwNJYxzhR3
Wyr12yfaPKpjTjA/150WwUQonpooAWSrGq5S1oB5iM3mD0OFBG2C75Ra0QBwg1Ts
4PMCIunaXf62v40t2KvWyMIREo8YpLacF0DCe6WGE1PVQgN900WHneNa0MNOFrJY
J+bQs1WE51UAnmDITAxYUl0lXt6USGurPmnPHxTe0XybH4IOd+SGvAfIPfVB5NHO
ZtWrsGegyG/It76YWdwvOX5qeJGiF+1U1/BsNIayGjxvuW5LK7PM3FJ/e3xhzZF/
NzOtsK76Mwte8YdQNbG6UswaH/5lzHT3G0P2gvFY6nENOFwUu7X6dQ+GFXjLO4f8
GGh768T0cAM/ReDy4UW0qbsMx1QfQnWdMkivjRQneIfcNyEtuYtFt8OFVRd3ZgZc
UIxS6/9zbKf0a1f7OvQkIylHXhkxC6hIW+mqiMOBOXENcjjf8CZg7FOPvbLAfyyW
1I3RQOT0iJ9ZLQoLepHMIu9yJt8/Ysz32P9x6BoADgNk6RMBZ6rJLl5x6d+cS6wl
LdY6NXmvAW6stkkoXFtDc52os1r+ubAjoETMF3YakKj3FeSyOQ6A4XZV4gExj5bN
Yo9zxpeiBoixIfx6tO6C1DgovquW0xUD/8Lp1UQJkR0T0+5jsliFbVgZIgbdLq/0
CeLZBqKZqmyprP4Hgkk25YFLXpV0qXs1NGdSG2wRQgRxffe2OTmSL1e7BUKp11cq
FGS3fdqBJx31YVdrlxKMoya5VwVVZK+UsIQDTbUe2tLDJis7mPlT4d30pHsNtYHv
LeIXuRCMcXAYHeLGk6wqKQUKSZN2sqa88uISjcKxuEKjpndEfILcWRLj/nlX3NtT
lskBOaJCsf4M0a3oMmfukzQxj96iXNNKmK97DfyjMwHkIau8fNOIyyoGTO5n2Mr7
r9Dk4sDbq3C5gUvNnPl6xP8IQ/kY1tLEP3+ZhInKudJF1FbjFBKsOejJ0ksPAYJ1
B7UR4eMoyY4VYIj3vIUxSHt4GyfoQKAqqpdUaYiD3kRYyceM5xyiDIoxewnLWdoV
l97pVTZ/1ZR9qFKfsenF/m8DUlhRQUwb8+iAqfgEDQS/RCcvrcUebNf1IGO94h69
cIfpNY9K4kvI+XINYJSgz2UHC15qBzQGEJ1R6wh2tSF12Z6NUTZAV6LGvTzMO9SQ
AK4q2f4irRTg45k5mIOSR2BqUD1XANVuObHokA0Aj+ZF+9ttkINRNZyymIOCetYJ
5FEAJSlI4kg+BUbJtMffODbv/LW1M1Ihvpq0RwEkh5h206H3/btkIT1KhkwlnYcf
hpcPQI4MRvQajsgBOy1uC3nkGxc9jgrBE/HhNliZ6aN5LVvP02Vs0m7KNAWEAVxI
92qVzobbpw5Xr9dw2kDx2PZhoz+a3b5W/CclmWuLg3PkNt44cUXGlhM1xAurClCH
xjj1VB1xkWgTZ7BQkmfQsfEe067GIbEkTbHCHIxCZA8YqR73g7EV7u2BaqrIYr+7
7ZGdvAvvJf/BMKmXJoN619lYS2ktBmLD4f6GFNtN6lUgU29nSTzfDYTPlXooo2bi
q5J3+769kjervhv6BE8cRSv4nRDedrHm3HZlnPeMT0BcPUzGWS5iEvHQm+lmntQd
uATyl6yTo8iQFQJE75ID+oAWO7CVZor8+ZjJqoaKqgPs+68RcIWSCJkBjk5RLxmV
Yn3uikplQDAJEzRHWV+dMHGbMi9XmIEd/SGB3OtahP+6lhDEP/q/QzH/t3V7RrMy
21mK2INYNFnvoD1lGbXeO8G2djSCBeq6yk4LdRxJJKgxL32oFgeCs31Pf8ghxbOP
4fQ0Xj6yQIMrodDcWIPSSWDIG6gNRdjutybRWafaJDvsfXWQbEPyFrVis2WPt/DZ
mR0JwDe+2x5qzog344yloriCkqBegk/Ji97EKacMLEUR878JRiBlLWxXaiZ+kkP6
moWRZSifZbrbJjRPb7dooXIfqUNtoXl1/InqK0AHeHBTNNFEmyr5xh6Z17dJdCRR
QKecJGrMvIR+ICMiujpkLjDlvBhrxKiC8MK3/ypo6IlIhNaDXVjZFF10xo1UNOwO
rOm7SONroZ6k5cqnMPu0z8Jw6uaOv7Zcsu3vEDBtD+qIKYJK1TPNXyUKYsDoECWt
5VfGNk1vi5NhyZcrm9QAoSOWhAttBoU5VVtA5CIAdx0ZQ9S+H+wL2QDQusK5KoH4
FFt9bU1WzLHjJFMZRG1hshdlTk6CEYj71vhk0LkKx12Z6BYUgpXNzeKDnRzYyfc+
sE2BGtHMYa6I+CxS8ZN+X+4VaWi6usU/UdHATZCZdmvBLl7IwKed6IrpTiFzV1G7
2So+QhvJS4eS8Znl5rTvC08fSeGXSl3JZkHwimGuv3QrhM90X76nLUz40+E1tWFM
oPRzpxDnIBnI2ZB7JIwCeAKiKbiCoxiBUnhTfCZxUPS5GSDUOy+c+0Rqyq37AiP3
3rhIMJpV69Z4kA0MJDRT3/sZj5cDN1WPQFFbPzAR+lVyGhT7Kum318cF1SU2rCVu
yVQuRy9lYW47hVAmP+ev/YTEwsENEYtiycYo5wIhHvrBzIOYD1/60gefBCz7evzR
qdE6rWueBFaTxk1+HIgh4sHNUJkt4cCgiHN4Z+HFHKinrO4iPSd0N8IqAtznX3Yt
uKlcA+CyXqQrIhyWAi04jRg/amle3m+Btj2SAHCK05V+Rcfq9J5ILVbqZ+6p/Nxo
eDh9wOg+62+Znwmdw+FLBuyt6zOdbvN+JX2EnyeCSlWSvukiml6oGzJrUgbDIvAr
CIcCvJbp6AW+yEk+WR/d+4z4Fo4UH4n3zHMsvewHnfqZjvCtZWI9Wz0cKrGk01gh
BgxcX94hgCW03/f3uX+SiHWncWlK8g5agHZApE9M0Vn81rSUxhS94K6FOoqcUzpv
/LR79a5IfjCzdWAG2bmFHyyHckOSsItDvTTfUtrYKz5fmgDfzgS5jZj7Nm+t1pAI
tDgEkLf6iWlpA/8eBuSZhoGJMZRmsmB3QW+/0sf9HVKz1/jOSmSYldqScoyck6Wb
hYJsHxAM5WOa4dFD8TMvlKW3Dd2QUmDYlYJTBjpggviXlflNA8I+GRGr4ihDnoZ8
hXFWX0kQUe0qUyk66GVCPDQhxiXox6SkBtL/mdblsfahbMrXtxUuMdnrZh/VKESl
gbY4xwFnW1zFuO0glUuztreEjvI8mvW+khD2ZJFJL2dSsB4eB2T3+sLtvRl8NKsu
nLCmmqw7XB7uQFf5HN53xC0n2DCZEr0TNfUHlI8ZuV8sgA2I4aUlQRBnxjh6DFmW
ALEHi3ywOh+hIUcCPlPB6pc20PALMcfvMSRLA3zBOVJdPdhN0tvyIRU9yxKk6zVb
JjloTHp44ioOCSmofTuvQDyVXbcbBDE8uXXS+tuneG2j4Pomv9DEMaBngfw6cWBl
wvaR8PayhoUuHgS6TnsJqPfNjXZpzTlAQgeOCmPI/xRKc4RSFgjPefpacBh6o3I9
EGQSmUe7/HoIE/XDQ3k8xCm6OTlcPUfd9KYLdwd6PK7w8ma2YrYoKn1lB2wPH0Fv
EOOVRuUxz4VNGx8t14NMzI2G8dqkKMvajiM2jMH3EB91Ync8MM4aRkI5JBTpsTce
QUOp7lx10U1o7JbuCl2XEvCyqbtaDQHaC2EVC5kLyz6FcEabr7l3TteiX+nYVZw0
EaTKJp1GGRIUZCY9E3HMqzcxE4p1OUc2IGuRsgskscwRPqm5aT1k/NRATZLemvNS
0Dy8h0nYinWZ0SncEVe6EbdXyS7JHV9nd3mkLSkDxMRS5QkUCVLC1OzgXQFhgeRB
Dr01rgwj49+F93Kmvl4UFiIO7LwvvW7RMPBl8SjdNc3wQI5XLMkPKqd/vwRRaIpX
Pd333NgmjJJryaOFybNAdaWWn5Ci15B7qH+kdspQzqiCG5CbLnclqHg2u47kWsCD
Tna7npP51BWRg5HTk0Y7IeLhHWrQA9tUNoi+3maJX7Qr13tB7khjM1+vphbkYHj+
2GGE/0UnHC8oyjbvpx1z2xSgyrRq8nlKDnrtBHviCD590NMflhHo12uDJx98EPl5
qZpjfkfBrATsV/WHOT3G7yRTR4R2Yhdi4f3csBTq3FYHJQwOwia/yxeF0afssuJp
wenkkO/CrCqKNfpA+VV6561L4Yc01vf2p8uBF4QBp2jWF3aO4PttVqMmJ6VUT/bL
VrC/0QFwqctjg9iEjk3VejZ4UzeqssFJPamg/sMgn1QestATp775WZ8upC7RS9OD
Z2q6VO9rUOibAFPyCoCY3/1k6MxpLOgHOgFsXbfjiwtoCZ+JFEOEpfu3WJo2pPpP
13yN7a0y4+KGUcOJ4zfSEGf3ZICNEsxNGUhNiqkVVBwATfzQ/WHok59wOLw1Mt4v
8LScI3wdWkMnrSbgBRQLzKOB69OobeNk+EnZe3kXNY0bPiaoH6NH3O4eVvfRVtrz
S/nCqrcZjj9SfK9fpVqEOwbT8aB01ITHB3X5oZCg94w6K8UeBJkA/o9WDcJzAz2W
diNDIYNiUWH76bmWNAvTbOtOQWdsDxeyuhOlYmJHOrFt4Jdvasgl85jHpDXBOYC6
iWj02atxmDYPGkq1rRKBJAxQEOLrx9lsH6MVtafpbSH7kVX6d8ieJsUX8gPaLJS5
HHPaR700o+NyNmL2GPNmOKX/I8GaUVmw/QRBvDVT1w8qbh5CxQld5kbK7s8ArAL8
TOM54PGVhSkQ20wYlAYyV/CQoxYkQb9l96uCTpNdMeXgpvQivzMKMk5nW2hZouvO
GVUUiS/nQZFmJqvmtQvFZ0bNnwQvkJnQHtZkrRBnebAHMmnIFiPeRqxh/xJSHDKa
/b2YIJnckT6rNDBwMV9K7r3dV6VV8OI3Ryqh9s7NBNbCBrvRjf3mgqAmLS3Mznjp
seUGKcKF+VG9D9lRNpBOBjuIhhUEP3pPNztCfpa584F6EFO9IS9JcBhha9IZNxjr
JzKHJhJHHGheOTTJs1snyPBq6JEQBkuW3iQ/azYCI31qh52yeopJx2PWQ419QK2o
qFhUi1S/ZgFhdcZCsS6UBjo9ligU49GRnhq3AOeGjW0rBqufjsrObLuAY/1F9L0h
qMYiEyGHO+ijh0Z01yvZngkI8XLEnSsy7oGzoWl6yyp41nI4FqU/D9naFI1uBWiV
MNFq/hLOTFFAt1lU/NpxnnyRccUeViFPnEtxxurRwhNpUZI7Hv8lpE/c0WVElaYK
xFPHPNEDUrGYLoEYiBDWqKDpTZEuSpl7p9EDLN55B01XwdDq4YL0IBFUvtcAAMHP
AR51aRV/hu53AQKkkk2kWdfxApzKe6Zv2SAcKK6foR63HGSOsrvYsnesWEX9jZmx
EzPEUfMwomsR2TeGaxyJ4V9ZSn3gSyQaLa5rmKcLMHR2DedwSlA0aBFL/S1YI3Id
VsAgsqdSe7/sL42x7XKtjhW8UF4LX8YvpEvRcO6S6QI6Nh2MUmw25i9JK6qX4fkT
V27cVzESwaPaSUMJVKAYWwoyYzK7bzavVL74QcwsyTop/VUmg6I1KqDtAvJ8hNnf
cOKsofHKIFmzdmtF2VsfGNLokVUBwx1ruWXkBJGEgmcQJdR3sNATpUdTeCwnTY9j
ZvmJGJ3Bzkf1Y1X1UNTfL01I44XDxUa7pyfwKTcmm9Dy8QVSdSLSvkK+qAdioX0Z
L7l4BwwLF3Mdn0Og7KSOGCKkrY5+zZbxF/dBpu8++eP7MLaUoVCl+7Wif2GZOtTk
DyIRtX5aC2hCNJPHNQ6yywp9HDdJt52PGkLAOXOQHtqzeL9GxkAaZiOKthJ0Io1z
LnthWIeHGeEF0W1oLRxnlY4I3odNLtbgKMlzgswQIF+ijdeEtxesHc417ccYbrrr
hanK2UxFbm4PXfi8QBrEqVWnymDB/udGeqoNF10EZLUNdNyJZzeCtaHLCOyDWhae
22Hy/tr4/EyLRBwG3umzST7IZ/cVU5q68n7OtWJ+rcbZTDlLYq7dbEhejBngksiP
D6Y11TNiuJj7VcVjcjDw6+QfUMzF5PKiDJ2Uxzk1hhGPxY9Q06Bu1ODGXY955qdo
c9+XIuytAfMvN5zCS8qGvIVFQuF4wVqe0M4HfTj69fIgyisYl7JvOiy4QngXYTs7
e4i0s1NyvQZ4Vy3j3HL5jtbZj0J1W8Sp9H/Pz2PX3Y7ZUl2RWQcjpLAszlTVeoZu
Pn8XBI4ku1Crq8dJzCeID3WF3bupKh9zuQXDlFi0t1yI6xwEaK/ffG7fc1S4ZlLF
MkjHSKR+0QdtuHFYnJHmQPcYwgjZYdFYBPSBlOmAuAxmE2nWPY0/E+Ynmb4YkG76
xXPChn6qSrmgA1FywgK0CkdgzIUPnXKhmqTyNTBnO/qvwr3l8da8cbZjVjz2nNnW
dg0+WnPUOBkATEZ+qvpyIrFlukuB/MadhyYXn/8T+TjzNKCTAgoI+L4ixvtFh7I3
aglrGU5kLlRl0C5g1AgiaYhG0w854XgF1O43JZOCtVOg8uMM9oORUQqmGUqjSUfL
VuY6dgbRXg7zUctj28I4gPLSJ3YOrrW2O2piUkudagZHP6ChpU/c7RE29nct8eJS
shXwpU/wN4JDcz2kMAF/nuG3AJZkojKVIzrphWtBzHJbVazLqNya7Xbfv/wqPp/R
FvK81DePuP1dIjyNJUWSPtSvu2ANhg7i6T/VIqppyqNMqXnd80Xh4FI1cWUHZ70e
BpPkFHci1bWhgEFIWSMJNdT5ZsQON3TJN2El2qEhHXMHJdTYfdPNW/i+BrB2qhSN
3QkDicuoZwCjOe/ERuUuxQFDMKwo+glktfyblUwaW1+OiAQfqce5xNDHjuMx3LRt
PB2ZEiGJwhjUPHHDYIECB2namAx6aklZDZRHiagQuRf22ZxjMJ9CRimczYyB7wBC
IRkgmUhRqaYXUpWfqdrki2df0aQnrlDbd1LHJKI6jpXaVNvdxjx67EiSPdHgba9c
mELf3QnSPwJ+NyxPNSCff+xKI/u8cKhKs1hqydBDcC42UYBHDmZR3CKTu2k2WvmZ
P1V7ygRdWVmsH3RKgMPCHWbb9v316NCrvL6D1TWjmxbJZ3F/Pv7HWnEzddJBeRyZ
3qwj/3KgiGH103xPdNLhfRAiH6urs6nLxKXgHgXNwR5nHQCqT0rYUM4UaAxab4lk
10XXW0T8TYn3VCjJgYUNn6n+eU2blM2fnZgJRVCjIzxQ9NUKJsz3r9H4sOlv3q8f
KIqdEFE37rtcUpjkhj1A31mSIl+LL6vH6odIhOvvWTeXa2u6fWDylVbUJJ9Di5bM
50SBTpJWZrxZmLFaezcipk7J9IiQheTROlBoGutUlBg0losylTRRxgDz9iyLyw+n
zTSVpZL7EbU7BuQST704CkJmuqRsWi6RkJ2o9VUA/+POlYoVoyVEcXeYSuF7ZUnT
+t4Ps8Md01vJvRY4VST52lEuhFPs8be2disBTuv+VdSqp3AmTsoDxyrPINEk7cDt
5Z9XXioAiS3mrOd6UP5T2rQJegzNTmfExZdJZxtMrnLmmuxRa0eMgT6n2HCGJQkw
Q/EWAl64U/hKja581dmzwwrX/JPObD+Jvh8lgSnP+hMLKQfjoudKthaPfe0icj95
qlPejt8BKA5e/vVNBaQmKpVI1zKAa+5vElNLyjIZxzt9kJ0bvdt2KoiB+28T/5o5
nVCQR+2k6tGhIx3EgtoVDs6iL621soSrsYqagm+Acxtu4a990WOfnyoipDJBi39/
QtGZylpnzUe4szYhe+K2CtONbtywhtYjbVEc1OqkHJoNqE5xDONYWQDubpNbO0b7
5owAU1BEvruuw2H05WZMY5oDFl/DND2docnLK/2Rbb2f/VwhNxNzews+dbznFRVm
vFi75+F+ay0/HcicZa/Wz/RKTyNXMB+vzFA881pYbuwZ0fgEzL2P268bXeYfinNK
AFezASKGRFPVFrEoGH+SdSUy5/CANvgsu/hcAk6QgUUjAy//CvgXLNEyecu3gbHs
5J2VPLAh0Nm+R9NOCzYTEt7esf+aSYmwKlw/SrNPynaYFwQivNGTGM9Q7UQW8Era
9Kz8Nk1X354S/xoceHUHfohp3JiT2+O7m/Tafsu3nALGpwm+TsOeb/KQgBMqh0GG
J86IyL71ewzP5fqdM2UZyV1jz990OCgfdFcvvIsAA2c72TYXLTKAUUTiQVkP+8UB
OmpDlngIAU64D3Y4ZQcJ3558S7KmfZoxancUf7aXKktqMmZsez+6ME28nWHt6kiQ
j6om/r20FAIGU93bjAS5ma/RFsylIHdWX8+tq0PWFLCXBbkuJ4rd20zhNb9GyZUT
XMsgQ1h4tRb5Xj5kqLabYIbFSMJLGCNBpM1+BYD8TfFktCnDYmejdbG/59sDmrTX
dcZxkSJTJY92xuzIkCmq+8Cb7JA5cBClQgKOZDgTNqdZFv/2ohGGtacMiOj8FoMS
uuvVpNT4nDMWTKCkv0gzG12GXeFuMIGKWGLEdjEa+YKtg8jIoZ03IIohJ+z+P2Su
4+mZM+26gcRjaqbJ/b7QpD/ibWbXtI/Mm5+qNJm+6j5Az+CNLd0qG7vcwfj8pr1B
zhmTgF9479CIrHrszLYhQK8cwVA2w1ld2efmt7j7w4nN+t6AyC9BmzWGLEObvUtD
7LSzcwR0L9ZK+7QlP2mT+OGUls3EfpaL9jbY8/PG7OIH9MckayEcKaBLpGjdt7kW
D1A+XQ8kNM0iL0rv/f0M/a4xcRSTXYl4d4U6RS/VdUXQD+tCzxS5nOPdiAja6yHL
uOzrfZWNCxN+nKH4qjIY1rPbscpjWxlMlW1ZnVQ3ENnJxGT60NqxF3GEJHMBpn7g
+zxrkODh8DWUcPUhnFAoGUudn3TolnRsbew7BXof15RtkreqHBUJkhErR4ma1oru
EfQSnOAhbcT8NVuEUb04Mmra6NZcuEDWlFdo1dwCZ1bK/0CiynAbuebqraQgh+ck
WgjikfadlqMNYPuHnLnmHde02n0bAZuqhOTjBGb/2J0oBmsSKLSsMEFJxF7L0oRo
sA1Oc++PrtPrucmJf0KxO+/nbNxTY+BGFPvCBF9X3wxAKdO1+vLNwjFHeqOGTxih
owYtixtjche3ZEr4nw2u9nNuq84WMnf1k5D3LP3JmZAnr8GLbdV1fKojhyZ0EdnB
mdQgODR+aDZo3izXHyZEa/Avj2YcjKSYQrt4KD/3WEM4FjTFWJwsfkmoSS3XKAO4
SEME5rXiXamBQCkcmBtpU3+siaRMRt91TtJGrPtnwGlCu6XOph4omHdCrnwXq9nq
w5NBlw+ZUMRgjLokQdsBrIDzq0UTJpoVlWCX31mSJqWlDnPXXDJpZuEclfCBNlTH
TbTejgSWRd22rjAzQsyQGsaQXtJdRvLngyhNsWOFByoBiY0GZ+7FKFLKQ6g5yHJv
sAtIdTOlrQbg8qWwe5j4h5CSdj3Q3T/+RrzqrVzmUTsqkQusmAyVIQ7l0o6JdRMh
PyyQlwSxoS+ziB6aFS+nfYUnvoszEwJbg424Ga4nifSs6at5k1FvkyWYplkOj6dv
J2OfbGbFHFsVcEYHls51xVtL2024HIMvMOuHL5N22a6BO1j0jRN8IKc4ruwzm98a
hQFQ4cTovIQsa17AbDGloM+4qbe2kcGppaNQKy7/qG+Azu6U+WeWj6nY1UZa8Wiy
Ni4BcmPZ3V/lA6BlxmTVy+F51myJCkRY8tMK/Lh+aLsrh2Wlms0McNuq/E3cSI3l
1Jtx2angKX8q4y5jtd86KCFlZIFZTB32O+IUKFamkpRiJCRid6x0vZYeKMCyYcpa
MKGa298QfHXNjSF1CP25ck12lcMfbvqq3JIlSKyuoLBRVTmjLIJRHLzXK/e9uEXU
N3+cRm0hnWhNkCesqrWt7gwCkG4QChucSvYzCh25SgEMhlXbS3Rd2AE+wh2I275H
mWfnYLoV/qmR8s0n2aTTln/xhaybM0D7KvKnaV7BFPX3R26aUl074eEPhQPeDRTR
6tZe2drFF5fSMjb+rzlWrQmr8BicRGB5fMSVcMvYWdBetejzRSYi0cBCII+Et8LS
LK7dz/SimlJosJSD/Z/BMHQuJJGibLQvk3coOhJTCXQnxU8xAbuWQVibS0WHczKG
wjKmYzln9k4hhYx3Dr1+rToQgyX2J486VfQ2nuQceqscsxQGGC/Tych2IQ75JfMe
dJfKPc0K/WfWr8po/Hq7IQzDqH2wr77aZzz3uUZL+3CPtHHbeMOnOwFFShejzD8a
iGGbIRMRdva89FvmNmfrj8D9YLsGNKreizv6Z8nUnUVq2B/HoEc9fM5pajyN8nz6
bLLZGPHaq9gNTcCZ0o/34UK1VEQ4Dk4PDsA22R0fSaS95xfHFESKqmbiT+Mr4TtU
e+nqPetsG9LlzFn/glVns1e1W+7EGfcm81R8Ju8w+9SbBfapwKq0alPA53LhlOVG
BC2ybewczLMrARxcZfkdZ7jnCffJlViZyhWmVuHBbefcVdb1IeAzMvJQivPnysgT
1LbCyVMsbs5kpi7Nvq3MC4IxRJPJGtpQmT6KdoGr01XFMcIPgqO8FAhk77SjtLG2
crBRxtbEJjnrYaYEwTgfA3iv7pfi656PZ0sXROLqXoFJufK7yyJhaPrL4jxl0g9y
QIcniP+ZvtyhDxQx7kxesU1kuYMnOUgIeQrtBrNRV0OHCd4z4DsSEOREZ0XzUc4D
1b/uUffnxNX5i3s4rm2Kg/MXbqgucah8Edp0EcrZ+TjF24yMJ4FBrMGtfscQQQfu
rvX7KuXWpXPrm9hiWxkU7VA/C5j/Z/o7unPDhzvL8wMpiCOy5LJM7t4cNia+W0Ws
nqNN6wAw9Et8UZ/B1SxkUgGf13Ycl4eg1gDKOy11XxvMPIqI56ETtyve+pzK/Bde
9qwrYUHIjPTvsQSco9FgRqAV05Juce4tFn0fpiGh7ir0cucwAPu6UZroCDvBgrST
F4de8srM2aLpq1ZbtWysLEJ6wEwGyo0255kUxS1upq8+RxKHmlkjAk+uvKhx3Bqd
cfoRnKkuQUMTUKCMCJ+4pLrP6OoYkJu0tTk5My3kAgIjGUYmHN/YyTpU0rT90ogw
M++EI3O4pnch7y6S4Kk91Nx367ViThtupi7TqoX+faqIbYprUQeSpqizWmogvWNY
jdTFCfMTuqdrUynSWHyuHxC+rKwigx19C7GRSA++h+WJJwXGaMh+tmM0Mj85zIhm
2qnuELpe3/fvbIxTCcJpzPMnxqAEUjbP7p+LhBo4MDB4y0hr/M+l5OBCU+jQ2OHT
wpXJ0NXVu5vzy+5uHp0DItBtPEnjKw7dJHya7WiabGy7YfDGhElIaEEsKPIMPb05
6BtZdP5p8z61koyyx0vr+o5sHfxQC9veexZ1sMtzqf6tRz3tCy2mSJAc4kpEgDUw
+05mCGoUe7Byxzbvc5kV4plTSve0E6JnnshQzp7T/I6ypUAElIQ88SxwMXzVLGDE
VSjEwe6yUbvSnDn8/YnUeXG1Q0cXWlJ6cKAXBhMLWVD8HZG5wcjknUcpdFQrRuZX
mNvIMPhfn9uTD7J09d7Kcv61s2ej/YGht44AykofWWiPzMD5vHx5CQXkUe0MQBgY
8Bu2V/2C7zjdC2d7so9TdG4xlmUNGINJa42mVIO/9Iu2+DO6Vp3wh++wJ+EoSz6i
OCU7eDzBeaWVDbu4MAlXtJU4fbCltDNQ/YBgNJnkq8n2Q+XIPEuoyM083bFygZqk
/uHwSoIzsJONQysUfkZphHfikcuGpO2WXbvnOh8awTV5/nz1zhcW9E2HxpmsXHMZ
CA4nlAnMj+9ZtqUIRJQdvfVYybH6yCuZVREZ9fOC9pkGr6R1igTan0rSVGPthnsN
XPjK2vn/aaVQkE6UjwFvQC4PC8PBV7FE61GPiXm24opDbbsvG+AUzHqdkbGl1kt5
tYOX6u5BnNCleagI6YazdN/c/Y2zpIUdA2VAlbAC5AuNMUC1xo/gmqXEbw3iLnTt
lmNGCCP0JFLvPKiza2YafeV+3jR61J+niE4xqkncxmjHBMKtsS2T8amBFy0JECP8
eEFEJ1YRpvizHGbITC3+AKTDYce9F29OQtH7CMHwF/6SDWegv7Wi7TUyfwcTj6Zk
wet8O6twAVGC0V/cBYQwJtE2UoQSkksnE0C76Iw0+7k7Ydp5fNQVn16C1pKIQKYK
o4L2NFq8iK5Kri+r8DXOEooTKE9paqsr41FiTDZ+YoW5r9L7Vh5p1dxLZSRVBGDU
OCUgOebj+Az35HanK0DaUWoZ7/5oSKqtAhc1Kfd4wGCK2fMcDDtSymSx5H+shkNz
zolxXKoZbHYDYKqBnPfbzmVnwTz+sCtgLetYVpgYA680Oc4ZG8mH+zWJwbDq5DVX
1PSVkqopo2COC8mBtne/Pzuk0f0JAYo43+IxwdaFP0qGmSIMLrT/8OdlN5+mANIy
HBKIZzE8bM3K0RLjXqc1qx/3rYK8Z8EA+l8MUAP4LTsKyijDqgGP2llaubmk0OoD
A3+nNopSX066h4NiAde2uIzldZJzNA6ih4czPqBkg2I2wM6dg81IGTaWZ7iigtCS
FpEM+6gtSAX+ZdDlAAGHAz7DnnIK8JhqAM9fdvprmadnwwoBeGmLl9v2b3HIAMi1
MPys9oMAK8V2RgmfqmPCbbsyCUVHMW4eCrbMX+yalIy/Pp3dBYDllM2GjY6IWCO1
CmqB7MMnaw88llgAyeaJr5sIuVUJ4SQvFHbo7Hvp3epuotmyd2/29h5FRKvMVr1N
qEkSqHGEJ7fjkXorguCUciAz7CG4v0gqwYolbFjo6eeXJCeOiHSVCozzmTzbQNky
tA21NJj4b5wN6znNKefoS8I7g+1YvFDfeDVGTZ/dR2glJZIHv4+n6EcESeJE/GdD
xy5WIZBKzqezW1LDDhzu5Sxo5bLiLhB4k75z4o3ql+9pDU1KskKrj08cTDwiTHt3
NIt0R5FXPCpjqopXuyLRnsgJcr69PKumVn+0Gu9PFQSCVmsGnRagM8h04jIk9lj8
9u/ekmr7qEGTQgFAhG0SppB0sYSKHiqkm/fhcf5zyM4CSqCsJbq+TBl3gsgbceVa
rVzz5Wz0+ptxLXNiRVf0mrX1/nPkUOfCFb5ftvFBLUifMBYtPae7nYlkZeBw0qdi
ox5uK3fHy2jLYmyEGUljEwo+/0OaXj0HVrWCWFOa/59pd/dvy28Imuw9k20ZqU2V
8wy02V/QWo8ZwZSxfZ44Mv/yX3TElfl5DQLo7RuLvEncnkpt1Bip5R+UpJI6EhhF
ivjx0GgLQE0DHiSgy93QMYtovanznvb9nAB/3zxhY7tUACHxkMc74jCW0ZWhOExj
RVfd7xflQHi2pSy+Yn/szmF4HFWnuCtRTWZCRUIpdgloS4WyStucsNmm7rXDRL7e
VXkXf5ddu9B2ZPvAqs29+iZVAXamDuyMSPMY2KYX35KVhQSIVhUcDrvMP/bkG8F/
oc9Fe3SrkcHnR/sNFwC/rEodC4X3cTVRPh3VmRbnM/t3qXHHVLTBAtggDmAEEdCw
TIRfM/f7pkwBCCML8DNlpfwC+5zwRGe9mCUWb1Ve/NyEzw0sYo6K1TWfIqFTbi5R
wXUeDu/6CJQuzRz8Vx9NUpprUBtorDqnPjFYhIHxPLRy7Scd/i9II6rbJAqr0+Hr
H4cVESaReZfdduDGgH5S4jYrn9gJzTcDHy73eieV4azYRA1u8NCX1PiLVgj9SDq4
eLG0pT014ZG6epl9WVtTJSDKTtaaNPNny3eOEFev/I4gaNjsoAXvkf6kuF+GZxbR
U+bASAn53VTaLw4HDnikLmIKBqTrtiCImzNJZQeOk6f5lRFJKwqHL6sOda4LLF2K
kuS1CKjB098Uo2sVm90vHIOhXR1uYuPVJa+IQ4UmFQ5woCOIOBMeloKI3EH6injU
H55WhUoXRoMbD62kp5OtrYB4KcxY+p0rHIJG9qRFADMmJWWLCU6imgenaz7kzedi
FVi2cJgLaZqiDErAaSqZDDtQrWn3/YUnYRKzoihdWJth1ZlmudYbzjbfXi4bDfaj
ut1GGWbz1ff85TZ+6r7WCL2FkMtVIieeFSi2ChjVhBMAIjq4I/Sf3NuUlS8tD4BR
p9NS5roYaAyDlr5tV+oE7+6MyoFLlwTnud5WD//XnAuB0e++my70+kw4K8O7GmVS
mAq2UfPD1j68Xojs3TNir15ArQ/4hlEO/TQ97YBna25+NAWg6ThQe4YHRtYrrbYx
2mfAYr72L/8jmHF+aW3YxGskEPXvHZAnuicF9y0EbAvRak19av4bXdh4YydeYVpI
ouscmPEK9dYGvZRza0ac632P3Napo5voSJ7HTHpugRjpJ0Y2VsyVl82S6ChSZJ5K
JQ0uregZiLRIBhqG/qd6KXsvtO8zpbsQW0HFFJn0eTViaucG3LudwAvJC+Rsvu3d
Vn14ZDs3FjRYcV07Ic/fZR6TwoK924OnoRGEQAj1bG0wWEKTHqFZ7HY3ifCGxlK6
Ay9Nn5WYnmOuU6jy86pOebDfEIMwcbGtZYoUIxgpEGv1QIwqwVI0DSjKj22abUcP
+S+nbGfcJOR2hIHfPoLsAueq5UE5esutjbsyFh2/yBylxmlJNKLxmWKHKlvuuK3x
/F63ab23f+O7RViVgDVHe8L5z0crM0VNtJBkG7M59LfM9hw4PN5eD9iG1wHwSLaZ
/aFH/f4zFffk64TUIJ2xxfStfFvl67ajxBFbweB3vuQNA3bcnXcqndbAYUStX5Q6
pjngMoTkMH+jr78//y05IAW79Jo49OJbhU022evJwFOI5Wo64MFYwxXeDtXGmgBy
G4pOj7OVHMXrXspmAU/CU/XajATzGmADVgf6irabVxbObzLrcOVqJ/yC+xg6dkaS
d/ZS5MGD5e6rl2pwyHNFt9/AFI8zowgqdlojmMnrPLMnXCryQtGub6yWpy05rNEd
5c9A4SScOFxgl/y0ie8xveyOdLaw5CZ0eIGtTJnfBDH8cZCdCsE0fw+WRkWIr0BS
LjYR0pA1md8V6s+ZxvVL6T+LgsrwKuTlN8Vn6Ab88vQWJYxyh30LlMnqTOaU78ph
STnDdEtsUsdnYLmkaq2rnKTNC+Ssq3CeXR9yB4m8MoRLoInY4jsCOSY1zqwkcd0c
COfcPAqA2sAVPj+kUchvazDlzGKKXL/rW3XklPUHQxMihLhUHDaA56p0uXcYYMxE
2tWNkd7CJsb04AHWkS12m6zAJ+NkCXwsi406E0GuAnZ+e1Ucb3r0j+CDAKX7rAKq
/k0QjGstT/7ZBGVL7U/1rLTAb91Z2ypG6vIExiLPk3hR7/DdruYKNUf90PX233G4
eaTkQL6EC4L2H/hUhv+5x6m05tFI26hxhd1eKaDJWAEyGxnq6A09jaGrGwSl3sjR
gWbnAd8rGDAV+cqD//Rbktn1iwnqk3uQZu3hdUaqxmqagOCntK4kB+kWacAz/LNz
6E1RRF2vnE9TLn3GsbWwS1asRyYF04YnGdjfJBgbvpX5E0oFAm1goc5kSlcFQxEq
FfZ9RTHMiDNiGG09WXJ9okesY1atHfTDtOzzGSOBta0HWP/iez9AtM9sOo19MUAu
6FKus0mhUnzUcAwWM80RH3rXJkfJhuUWPDPeYNUOM6U3uSbm0u4NfQeIrvdPfu/r
o3SLyhYOh7on6n2YRfx7dqKlpZEmaU+1n/nMeSAxoA/E6v648Qp3RBoi4NTf60Jv
DjymsQJDSlOe+5uwtROhvWUo8EsMTxx6/pcMuruN7VztzAvPy51dD0+FM/x9EwZf
aTa1MeybiCLd7Ru3GsGUesvs2XAaFldLiBNOI/UGVasR08jPYUpHMgA4k6q6apLI
qeczGXkDJuusbcGeka0SXw0G8oF4llfajuj70auGd4KpqHM7LsVC1UN54mBJu7n4
OXhUHg0iQikBYq8xBlcF9gwNPzY6tD0Bq1hPfqcm/hf31BxLiu2WR2cbEJsuWnJ5
aYjXqBaNmJ6QoAGqwX3xPsLScKEGDs9b0Y7kEW4I86s8am5PoHQ+AC5RrcQlsGqg
PD0A2+tU97h56rfHJx71nw6fIw+iipy+aENu8tvwgNKoo//GhIdl1U3VX2Yi356v
Zk3cDrEvWu8POqFQ+hRDyQwHQvJyCO2PaEA0pjWIm70BV+4tTbWLpgvjGCKvGTB/
CpZrujfX9UiwsK0fudmW+kRioGjONqTnHevbQOQ6uimluXKZaBdvLsJJnJdkUR0R
Dx3kjJVX3cTFu3wwQwcN7sOgwEdTFqt9/atK/L/yxHP9ZNhZx7FxQB2ZFYjB45Dc
mo6X91VH2d9kag4e+r0PPRyxGDU44VL3b2e9L6fMSAYRPF5wino2u6ztsnmaEbBm
HrvWp0OlyVMJMRZT6tqJiq0GzOMPwhjH8PCKSx/eVp5kHzXuH9JQ8Z+Vyqx9Epi3
6n1n7Gbd5qQ7BCz4JO+0eCwqk5WxiAOJr+9qKNwsac0DwQVIIJv+BZJSo2Bza9es
J/PvkPObkie+OUvOW0Pt6XZDQelit3XeIvLpuix8OJ/C7i4Wv+0Buaxy3SJx3MPQ
BjHaLsvddIhdtD+ZEuHEzA0JYkBz4JtuteukufC9WogtTkBDIYxbx10O2Me69nvL
C5KzqY5IqRnn3pegG3xB9j6pOd/Zb1SfO/OgyRxXCcy/aONxlrNbTPJU77kAheru
0TiGAeuQEINNUpx9/MjqycmE3AYykUR4YuCe2gh4fPlx8CiOh8f0BMwVf84t9t1Y
N2M/g4fNRSpHgAtT09G1vSE5ft9izdgyMNDlGyYivOb70KT31suQufHBBmH3aJ5T
19Iflum/fUjLixXdo07KVF6OXwiyr8CoqFDxxK+RqLSUjFl8LU773SJIK9DkGI/u
3iRexmPK2WL2nWc/oqNldrsaqn2YJzjUTnL+pwEg2YHU8QixU/HTmctrZzwuW2jM
zYuqTuAm0KpmE4p4RSP3rFxhbEzriUYOWqCcQYRdIimYCdstfVIC9S8PXbo6pPUQ
15Rc7xHiz0tF37lGZGkKU6mYvLOMAW2whR/g8/FeWelSZFmp5rQ+fOXePcVsBvfL
Vx4/z8nCe/BabmT1pSw8IQ80T3toV5sXE+0nTK91QhIkGzufLce4pbtXzni2a9Xq
GzdfgVeXkNjs2wcAspqTN2+AhPTJl+YJ4fleq4wns+C5ggWHvHxnnjpEiP7NUQ4W
fjtVBn08xG/gtIAJwGVl5i9T+KhtanTQjFBmx9RcRkI1aU9qmUUEPG0MFrv3BJZ0
7W/z3urtG0FtXQR2INm7wFE7p+UcqDv3nNCuGVA/hEVqz+C7nEUVLPQxbslEDBV1
pqiyE+mey1B2dtHDtTqbA66LZJy4NpTrpzTQhU1ZtTGWpGP6V/RgRt/2dGWFpKDN
LzoLFw7wSw3BRzzBWKueeazu3cKVNO4DtbfAwsP47iEwf6gcaj+iSjmdAJjvveik
FkL/xVG9Qo1E0uORgI6/Cazgy+bclf3N8SN8G3s0M6X3lUI3pvz9iktdev5SW2br
fXzb5trQ7A6VG5kK2r6WxeI09AjzSf05tpwajEdNN0d2GAbskYOuVoFUGxj9hZM7
EdKUP3oD7Qz1pCo4oQH4D//Y0QzvyZul86XoEQWB7XdcjgXuaxwQN8qTag8XN/bL
WekFt4+Nimk69ApghTIkHMKWzrRPiAwm+CNEfp0WyecT9nzB+KwB3kuFlBgubExi
+CEMuip8COIG0UFhOvqR/3hooA0dY9Brsck0NYXuyBDqiAzdgvyDmEaxQPS9aCGs
nqNQUzv4eGGZP6Do9HKqp5Iopctsptoqs9lcMcK7VZJmY0atKfvMtWWkgekqw7De
xxIes8mIGiZCtpsKJICQCUAI047rKWCJtWJPz6NrNrnWhdfLmTrf0ksOIctgV60d
9T4MyDY8X2uDE0lAmTCIkj8fXcS0Jau4vGm7D2Cuz5aZybuQbgJrt3jw28ak5KLf
k3jpxh1BHKHXjHo8YoWDhZihFXFNM55XO0MF3egRonRPIFU8Yy5YmBooXQIYd+o8
RtKPg+0XWwsdcUWAtuyMcwEV4m1kHm5JMZ/OGE0S/GCXT3aukulo8HCX54iGO5cq
YjrIsYu7RNZdkKo5X1l4k1pr6uTFs7k+cciHV4D0EMXMykgEteKOCZ7x/JagRmk3
HDqYFNBzd7lyrsH8epoBRtAShXHQ3QI1u5MhP1E3ZPYTwg4gHl6eedl5t30FtZpr
HrLHq2rxdq8qohixDse46cJpv7lmqJcEHmQCxFT0xk5yZYxVbpL9q+tyUdYA5BSh
68nGYTQxVdAb2Gr6WGreRFQd8Hdd/TVaPpwKAXOUSS6hw7EpC1mFloohtlkQH17S
8t2rpNVqLyuM1LZVr01zNBeQK/UEIs6xT+LUFdhQShW9ak/Wqw4zstyWRqM5RIhF
diRd1bMoK5lFCS6X5ohtSnbza+0rOSbetZ8l2isxLZ/Co083nPgFOyKIwJ1p7fkz
Iftu5DaXGDvHcA8rm2hbptvuwVZvWJdMLzm2w0/UY93QoDT9S9JD8VEkFbjxofae
ZDNgN5/ioxpntg28bEXg0mZzjURirg7zrxSGn2SS+dqj81iU2pAFQy73Lsy9p3LS
62JC1ytFlZRufzXdnwwZcA8/Qs6iot7djidFmxd2NjOEpi3LfCqMbeLcnKJ5ouay
u9TJH2RO/pqcpXj5bs5V/x4AjNMtaPLaA0T0qAmdc+DuOy0Bgutmq6wmAwkG1kHT
kJp2tRExJOqTeKjBzXpDoYBTNzEcG8H3FzverrOOiY5m6RIyuRbwfowtosfzHADc
IPMhzOd/A+7LqWMkOLs4rVDaAc/0QlUaH3gSUYqtgilZFxtuqCDPomzCHz28Ly6U
EunS5LkaFJZW9KCJyn6ifI06rDGip1PSPcAIhgy6hrXET72pB7wR1wEdAHHJM1ib
nFkuv7ErSdPh3nPaWpfvzn70k1ZLEhd8F1yvpPkRhkGKGeyM9Rx4G8knLK2nigdp
ikQEKQ2HaETgpEzXLUJa0FQX7Q5O+8kOz+/a4urcIW1mxnfUuNch/pMVfrqLS0JC
LzCowmOnZVvOV/oCbwCKE9WJZ1gYLYUP7FsnZ/ljlZ45Hh02NbHXzw83gXB7/oBf
8Jwatfrnf2xDII3VSOMtATEhx+Z6ALc/yUW9ASsj+KcRgSc2QtdMh4pdWD7gBfX0
nGZbWpm/RXZ4TBrZ2Rq3mV5S3CyFXkHhc9Z+4sZAuuvC2FAnxrcMG57+baGsLSnP
gIsnD6GsmyCTZyNLPwrKvL/xcxfn4TDCg5tO+LvVah2cHLOWlZ0fUA26XNvV0vr6
bFxdjArCcIyTyV/i8689Oyk/j6zLcEamrm6bij1K7VrmOHVCK5vshHmGF7DLu5Gy
Mhp+eRiRtjuGuD2W63iCmfMsj/z6XG+r7MKZQcgFjYHeh1GjoiUmWf9gwC1rHQ5W
tF9MAVb3/TJMEHoH3AkonBkliSLfVOWaDvU+sFjBxf/x02ceWyUM2mOH5uVpc9HJ
a1/A8FM/MLs+zPbjVR9wDv50ikHdO7fdHanMmcJXr4nXcrBwWZpWerzOeomM5hTS
N8WOrsp/MmSBeglLWHaPmlnDrtPQgFqPjN8000p3sY9Tz3EjJi6I4sofoQ5BNGBt
4Bc8B4hHDeEzKDQbeG+1hMXhzqfGtbpKTpKMKfDmIcyOES83j7hWOHDZL9nV7bLw
9Kjuwabo+nNfdk9A9F4EuziFvXz67Gecq/1F38dexmVRFp5tKbe6BlzGTNUlmfbm
gSWW6BjVYfeH/LGjNT5gWgjQvrvf3ovFH53cUPHAltawI40FBUIcT67X11XnjhDz
QnRda+9HucDE+AcEu758m4cJTk8fekZMnvIMnM+YP/7bRexBDsQryG9h0km/lArR
unnPyhcbcp3Bp4pqzJoaGDNQEa2JbeGxf7X+ITrZc/UXb006ucK0pNaihgGnrqpF
vxEKsqsXgtDBXeY2aNDmAkVRsl8Ki1urR9tpTM2YTcihDNs347BvF5o1fnBVfkrX
h/BgFSfBK2pu9ZjLcDuPm1hYPFdYfCWTF/2gOJO/5w2dupfgHV0DUz34ckQO8gkd
Kt+dWruuYJ86lisiQsXMhZef59cRBMbgElFyyvXhhZeoy3OBs/rg8+7UT2bxmOmL
AU3m8XcTEh1o0/D76ZsUTyX+b20GmAKD+EM3shvRTGQK4x6An3nipjaitlRBawh0
WLLFVZL3GNVmf+222JgOa71ZgcyLwvR8LEpqn8VUmqhYTu6mtBUQ52FW2qsJA/z2
V61MDxAdbXJZxunXspgNKKFjA5jB8mS/rGPq2xCmtk0SoOAl4G+rHgu1ZNcuUXRx
F0Q4sDWSxx0J/3OfznvW52jvmGSYMCCzAfIWwHV91HpsoLtOfjy0Bd8kkKTYByfd
EwM1//EiioosVr8zRLWQDRqQNYrxYUtyyqWjya8sSU2COeGKIaFxxILZwZVoAwbN
hVNcE7G3VbB47nh24lMilSTTpNAiT80Taj0adW+oBcNCqRChTHdbF99fVVl+G5nv
9Mo4lreADXsUkepDaB6ZQvPdp5Q4QXM3n3M3arbuxfI4KgIYOaUs/SKUWVDvYXzw
/kOoBQlItvOI1B0N/UmanlEz9gdQA2D87p87Lny95A6huaE5fm9FZ5slMLAoqKu6
duHrhV5t9hAdLytgcKjvV+1Yh3ViCRRp9AE2X1w2Ho5z5byRQ5t06wMIxtWsvkis
3N9/K9ueDngp9DFmgI25/TZNfiYK/60o5f+nOOsrGqHIVTqR0eAuH5FaA3XYefu2
UidYOrdc3Lcg2FG5AnlQKQE96rEn/t1RDbqQ91jGSvHlbBPvq4vKjv6/FHzcYpvQ
2Q/Q+A36ZQlbrTmQ2Yi+1wM4FffArSdtzeaxJrFYEs/l46lyHi/zaTQr/XErBM1t
/BVymcOySLHnQ4hq8qkO2GkbBTkMcaqLDZiXNsk3/fDjQVxBT3z83PpLU4h4/4RZ
ias235ArtsZSGWueD4GBXmyI1D3MHSHo0kzbnsDhIXmHkIqDItTHH/PM5DGQrtj3
k0FehEVTiELO10dqfwfSMfLShl2QEyyb423LhHpGDgvP/r5sCbqJhudh2xhXrBEo
Z+Ihn4korc7tItUYv8paJ2KGHHFUpDcgkTlGk9sI6sqrfOhC05+cmshD0Cs1Qi8M
ZMYZBc4ZxrsJFeCJPo/VvsRM9vOYPox0vu7CnV+UeVVSxCnn5+KcEdi5KytHffgy
kYWV8aZEpEtwjXK2+OaQM4lRbc57xjY6ceqQuv7UDCuhjwoMND3VXva9nLEMnZJK
T2TRGE4Ty+DTxKsZnpypSJk1iaQZU5vRAcOwpsU+j0TVKDUbFZXLXiBVrrRniLbj
oQr0BnWFkE+EDdgpDsKdiiA5ZK45gt6gg6SsfGCLtdw7hkG25GAIH18mb9y8FNsr
1nd4NTZQOeMxnTWLgUsjx+l+GmWZUK4rsQGtWl1QJ0xkIHDe6DeM9s7z1Dm0vzyY
+qYKoj1ED0DOPrjLJFizbN3lvt5DGELfsNOBWUsJKLfHfViVBRcQkGKe3EJ3XyOl
1UT4yiIFKe7r+rOg7wIgleEKkGMTv35kncBZTS6c0tb66blydfzMKie+3i2zuQa6
M/DfAFjHcxHD+hdTV82ocIjVkjeZ75E/szUDalZi05nOBmJYgyfY2GW1Qnvv8Xsi
2+Wg+6ZLY0xw3/T0AGzUklbp/yIjKqsrZppjfRIVPx7tDTXtqSsCvUDULbQza1tz
jc9zSYHvOim0Hd++odOk02CHOm6jo83MZEhFgccsP3qiggsnGM/aUyzjEg5D90Aq
shzaX2X3close3TSxpyNj3PMEvQS0cdnrFOQYmX28HixyEoNuLaKrDeYh4wuGXqR
bEVH8EI/272sOlJGS/jDLoXtHTbHLx9Dg28XjoMi02Tv935mEjgyg8aX+TAJ0wF0
0uGpulQZlewK0E8w789AfT+pdpK85rTGU11GsZPQh793Z/CJxv0JtlZFaHbWRrcf
ed1hfT1iEFCFzS64lhfwJJhMmxsGV14YiWXsgneLYrPKvIyKND4Fea89nAq3VTsA
U59R5vJbwN/WY7a/dgywLxW4UKAWse3xyOv5o6Wm+P6nSQrDbZuCA2ZOwZEnNbCA
XTbZ3/6/ZLtCCb0dNw9E8+RABY+K/xDjHzsNl+p0uvWtrewnzmgPVvnqIZpnFD02
GfbEmfzhHsxgfQh5WcKJ0n5rxR7Xqy2FED636J/JjsPfmhj/ZGwa5vT5f1e+Byl1
N2uJxxgqHibHY8b0SxbpyftKAs3ClWZmZhWF+cwnx1hzfC3tVTuqpc9oq8lKdTGI
5kevaCiJEss+p3p38xvLJjTux6ZfBOmyIjjOdKdFxUU6sYeLj1a76IBgllNa95KK
uXCT05qqPLCvY8S1N4w7vKF1zu81DU5RWjNFVsr6K4caOeVgBH19Xyt0dTKOGRAs
eZI1zeqlUOeW4rlQt1M9TZQyFRcq+WPCXf+NN7fjZ/IsiU1+kdjm3OB68nBA33JI
AJ4leIXDBpTUVrja3VEGAjQg+jdp9OHAH8GUqHrZ7xsJdaDduUAHU9cf32mWTSfA
og8Pfz1Azi8mQybgf8I0/gDzY/atmo1sXwm7QDT/WulRdKgT+uPOeYpEasJ5V+f6
zE2y9k83tEd+pWLvFIaSskMGulP3feo+cG9U3ENVFFw1t1i7g5syuDO/z9nvP23z
Bjo9L90kJV9wP26H9vxAAAo3oSSjDT5YHwyTh0sqjzDtnf1+7DxHOWmRo9iGMGYv
cD3wvfZtTG/xEb/ioHPah/pMKfRPSGd8wUnFKhclAZ23qiEtlsngujFKoDoygnpi
mkUnNNu6IbMlWC3a551jbChcv3WPRg1k8QyWoLe7OC7cs5mGWekA9uD99xzdZE4G
a4JymXQVvAe0X1x0uPnE2xSr1llb40oDMawBmXNtC3zCXJfmSEuOKrKg6GThBkol
uUp2QjX5mViKpj8/BQQp/66oMmxI8TCOY0nNbImM9O3ZkCJFYhcSA8t04RlstNzb
Q54KgcaWjum1dPyUXc7PNRNLbx7mKh4j4oXV+h3kSfwLYqJQ2m894UaI9a2+AfQQ
LDYZ657uFF63YjiBJ4Y+mGOywKnJqstMpq1UavEYdcvFnkQitSCg2GyiJmUvOp77
E03pa85qQ9/MYFuzwpwjrBA46MRTMxfAkBXDAe1g3868rTJJnJkuDITnYiIzvu4e
azJ93GWOMh6TUOl8kPSeaZlldRz1nqkLie/DFk1At74p6QVOE0TzvlNk8U4/E6jH
ITxjjE3Eo//bbTeWESQDW7xNDUMBpo2hi4o71fWxkEif1hDwYS7TDnnwdfwCKXok
KDipYoXS5fHwxoXHv4WJsVMmNx/h3WTayAbjq/DivJXbnoBavEr/FSIGnZ6HkJdc
XuQBhcjhBpYjluvSKaqid8DuvgjtoJBwtEufT6FZ7sJwe5Y1lSmGkAX3xfy5M/Gy
PFWOEPqqxDzjwuddgPJiMBVdNV2IfpXTY9ICqTo2W1DZC843EWCiEJ75I6Ek6mg+
ytGAEwNT4tyhGBfH54ILjZJa9pMOoILOil1zbTaxCmtnm2ISlFJKdaRPY4RcbW/q
5sMfsM6lqr/MZUEiBuWy77Y9CGgCo5DyDO2yEGyAxxk4xHTMKpiSgQCwiG7VyE84
mXeZgH07ZyJ1N2ukGc5t0zfPqUs+oYVyohlA/XH0rHp3SOQtP8wyHCB1bZ+mwaqm
4CdNnUIXOWFaT6xxYSTfh0TP+CqYbdlDN7+/I8nsxtqDzOziVqxLWVsCe5Jx+Flg
pFqzNSc1lX9DQMToIOn/nEMHmo71sI1yFAz7cAOttEvPWgDtnNp6QJ2heWissQaS
oFBOl8cXKkCJ3agAbrHK9dBq8efi3JESQ6sDwyN9GGN336DcsGXc0+t2JLJlN/+z
Mk041yYYBVFeyhTZl2yKM3V/uPIt6JO+2+Cc5q+H+1TuIpgMzBVE45osPuGLNflQ
KTDbb2+TdVIOXY6okKZGUNx9hhcbaOUvhW/i8iA2NhxdazMedox9lEYxidGFfpg6
hFwPYWpe0fSOptBv9J+WXpWDs+DOVBUT63qs8koslwE5eQSaNwqtNOMr0S+6J/ET
0UxS2ILQVPYlTWUptcmTSES+JeKWhuWbIdG0iecJ/N5uDBrop1BhBZzW4n+HJgNn
0aYOCMIvx1LrxV8KQzY+ZKsOPeOGLPWEpdfxVFs7sqLqdfyXGVZYErTmLaWF5RGY
+UEancxUMSwARB0b/ZojJ5J7fuudOgCKii86vmKUeNYCMZKHsnCS6q29fuL/bETz
RmrtOh1Fa2vz2NDFcyfZELs3XLHCeNohYhIsU4x2SvMErMWuqShN8wG7peI5aDRu
UrCBt2FUHK4tBHwQKWp8RnZ0bYgDUNpAlFL4ltpMGkegrNAE5RY1NWkEZoGSwiCD
R5a67ueUspJiQRPJz1oAnVMr75LKIuR3w7tY+6tQb8NIpqJNHH8DDo0+Qs/M/rhE
X6hGqWY144QzzQEOqXAiAX9xfnHzQG3UGJjDajq78+OwI+nGVKoFZR4ZbZqsr2Ak
9T1TlYgnHQNNsK69qDLDTKSkc+cx8AaEyHd4FGY9f7+mGSDKul6u9HonJeE6sUwM
md/ftgy99xBP0AwpMpHM4Ja9LhlCML0TJoqcsDZ62M4NllXREgqfMZUC/HiodiC9
Rij7bC1CFxGUozcrYfIywUTq41ITK3LWAhsKSn7S5ADdWr5GXMVhtKzItah/0p1f
h7EQAHgMoRTTohxskh8LSsXasXSJqEHyIMpGXAQVFdvjAiq+VFcsY3kQ7pq4zaI8
BX6CQWfOU1Ry4ErSh1WuXHxVSZyJ8TZV8ZShB8NJmkvV61piRRBjxxUgTcrwy9ZI
Fv8dhScik8IKt20g0xzBKl8CJruciZP2PEpP2piVxzLdX/jWIw3ut9Mt5ua5hkoK
k3I08aibZktFGsylek3EySwRJiN/RWNyDgatC/wDITbjJ6UEdVrcp4SSJnOeJE5v
udmN+fLFnzQx54vLO1G7xX0gYH3uR2eYkK9XJF6ZhC5ppsruFP7aP1XaFftO9Zd/
vxvqRWv68emm6GI+CFjmlbrDU/9FGdTfGE2Om2zQXFnCDShFhf8F+D2ZFZM4oGVB
XMfW5cPBwrx0Yhjaccm2AKd/eeaxk/CDW0pLil0x/1IB65qB/u0DnHcmzrELg3Nc
FOm6llyfiIg5URtPUQFRJ3+TG4ICo5DmbP1oSz+iN5JDQw7BW+guopHALqVJtt8f
4KDnbU7Ea0Cl9jS6VskARc5Yghn8QzIP/DMZUgfWEDBI+p/lnavEzg6JL3/b/lbq
gHTuDdkJDSXCc0PIcVRzqw428YyNTF3CeLM5mvInJJ3gG85+ycKUS1aluvEugrYI
A4VEn7zWjx47bSFFOdl6l8BprjcxmFvJwahjRoftX2pogQdRTIJCZ9SA0xR1j0/a
D5Ht0K81ml/GuDuvYnhwGgXZtNM1yQHY3Clvv5ytp4x/muAD3nOISJod/KORwuhm
YHUPdW4j4dA7dztCG6smrrObKeDTqxr/u0bGZvuAtXFWgSgsqMTUhNLVQOjKV90o
sIU705k+SqhQ1zUJ0zhQE+qiukXxZBHntfCbtKSA6moYQh5yUQlXWaw+UTQYf37v
eyCK6TSYWEVu4RO++IbELAXxN40jqLq83f3tPy/2b1yjaxGKganHpKOZ0/58wQwi
Z/A/zWIKjIeYfs5U+egqvpHlZwYrS4YQxoTpxJVj0OpG3FtT0KoWHDPCemHWmAT7
p55IWXFEQevoicPMMAcWbKaFYaYayjwooX3Y1j2jSG3nTqRm4feMMFa5xJw6c0GP
4utsmIZ/fQgJQN6Fv5Kezghb/w7TFUewtgas9+8kG9lQCDGM+96OWwscSe3k+Hg6
57hpgvmisQKrSgzcl0ClQPsxNpIyNkoUDmDYINLCZjCsZ5602kXvERdQRYMRXeAN
lC4bTQcOj/GqEzLnveSH/8RmICNR6s4dTEno0+1kP0XtQc/w4iMxLxXNz4rwmuph
bj8Nn4YW5IwnTPYFAMUUX/3K+OiaKJ3uW1OkyRANLQGsCyEuK9zyXNkWaFkLzuPU
zraS9XAtxVJwApvf5bOkARg/oP/MM/CeZjvlYJYdMKjHLOmRaKleTOXm3/tZnLUO
bCWnh1amKof6mOGoQ7RmLmet0te6nuDWp6PjPqOtYN2p3ptpAu3te35neAYkiuY+
WigODmoL35i4CoeL9rs4etyvlCKLlej6kJxHP5CrKMRGehdy4tsjVhwwoGcBepvT
ZTOhYlj/axmXxQ/c3F5CLZKqG1ZM1zpq+eDA25STN+++ocAamkBXwudH8LX3wOoV
/nUqxl4SkZ3LRFhqhwE3s0EErmW53I3OVTto3A6feNdUEwu1dUIZO1psrrgg72Wq
UixGdt7x2++lAZY9XI9MDhDK2Mg1EXZ//+famhihpj7ycZw82muc5z1Q5ksCbRcG
hZts/nEEGyUwRollY6EJsfrxox1t8HpmXNK+l+eEokjgruTCZDyJaOUnMtwQtz+1
bQ2T7j14iswHzzXcTBzYnHtCa4IKN77c1mvxKLKzxDmDCaufu+kvQKAeooQcjDHr
r3QJgC8i8M9oXsBd8mF0VZOIgMdH6LOT+MOPw7QO05G/HSFjcj0pD/XrlbhumsZe
dNE/A1IfIK1Q+L1DgUeRN/FqVmXrwfSMTQkqkbH56UcuUm9t5H4kiZ/PxILpFZRB
JH0bLz+02BYr13q3mlN742VCYz8gQ50g6zsUUe2MUQgs7Zj3OUQdkaSIXTeuak2x
Hg1gjdEgMzx7POrOrG1ZfFU6sD3B94v5tLJhN292HvqTED2YBvQId8HvB9R+uQGV
cAScEuXgE6OE0scSoPfr4s7EVkla4gEtFJ+v3Ks+r1zWaEkfqLSGTebOEkqndGcv
JJfr8WzSmbfmerBbv0n0cV1lzQE15X3dRqZ92Oz6jQgeyLnolkSRTLDu41Bk2oXV
MFRIoQXfg42eskP2oUC9TCa8sYfJCwwjYL6LJ0+kvsNdfFr3hhI41/HjZgmL5U0t
DCnvk51tfgqJPZdv9Zp3dajmVwGmF3n6+MRHOQCs8hAlhPYoOi4vANaFZduQcUUD
fjVY1YN0XaMnBsdd8RiqLUoyrkLcfiqCR3D3oc52pnDsPFuVKQd7+RLKhW465qBI
Npbz6J5A4PtlcAvavdcjCxQhXEeMFce6K+EsZifZbbU7zoJ6shmPqH0gNeoGVa1F
LCzDYxfHOAYrGaZ5UtB1/ZWfBR5WYwraEzP5OkJLExQfyjhjAHT6r6jBDMamwCUH
7vwDCGgyhFR57H3U4UT+JivVuHEyAJ8HsG+l71YUOxjzgAh898Vs6TGcIExB2Lc0
BPImmcQ8zdh/YEbKpk6oLVdUfbeiNyUeWM7XxUuo9DXVGah+vQJ37ArRHNWouJF0
8ttcGV6kb9w7P2w2gOtAja7d9+9iJXjAf6dPSJaNl0IfEyDGUB+K3yIYv70FepV4
rIWmkhmVDfpQkZHA+jxGgu5AsmpI5/w7LWVLkRcrZeli2DcXVWr30p1rpxZWWho+
SHIpHPT2+2lXrHCKGBLlI5oDtfniYj4y7ndM36+YH+YBwJStYQmYbQdV7+8KXY3n
SFAxjLyFomOTOoVZ934oz/Som0RiBkIgMZ0XJtEjrr5S+JgzE28GNLLwoksgVunf
bTWsqfSMHZPdzd9nudCIKM4ykTvKZPhHikQSrmpWhiPRyXub7vX5VP7CvdkdxE80
SrCnr1Tr1NwWhZNjs1kyVnUivSsJ840zykdP5LVQ0vqIXGwt5BD47/gD9a3E3JEo
utmXedLdcEe2lPu5O8CqqfwPcIUm+n1eWi4R6uYlhO1OAwZ/KK8mphFXeqU+FXVd
UwKYrRbASt8VxBj39C348F+OrQ8wsfQDzhb0w7M+i/XtH3ErIYT2shJVXR52UdQW
wpYY0neha5x2nyX731Laa26C9xQgVTag2ma4sPdCWVfJZwXThsKi/d4d2ch+jnqX
xCzdHbuwwytPIQnB7Vn3+4g0Okx+yiQFcDJgNa7zTdxlU9Xk/lKDh3FsLSsPQ+cB
SQQN1/qBD4xTTpF59Sh4WedkGvZvATVJ77plinq/kWOZwg+gUBNSpOKcrojP99bG
YBCmQ9Ikv2dtNMRxkIno50qyWARID0Ge2SsZ//i4Fv2+qKOps1nPKuGWNyjscUFO
HPI0lGlY+RqeTWr8Hpwa9Gi7NfFhFkFtveCwBgADz1E4EJnj8MbR1AQ5bMbBJrVe
65IiGwvetzJ1ofxbMCYz02g4enfmaDWPM808GNfsfCWTRzY+4zegYQtdZjz1vsjU
z740v5+ZHAubhSAejXWqcuBzH9hOMjKpczC/rmbj3Mk/Es3z5mUwKoZYmapFL7N9
oo+gU3MssaAUy79mF3beV5fRI91rORkAABG5XlLpy42iJ6jPkucyrMgwr8ucN71s
2/CeaUXBWi3q68/aqr8SbKks/g/R5p3megLzrYk1Ve4Fith8i+bs1dSBGjd8bXNO
tvBXKM06Z3lfDgdi883nPb5FdFL/C8YDn9UUkm+p5QdjCOzlyImf4XcxK/Wp+3oe
SpEGfwkWXPt5M+DoN6YKxGZ3ft6IKWUFJ83cF6R9rJjnRSx06c/MgRq5TGG9GxfD
NV7VAzJfC962wZyCzxK3Za/P3+vQ8TEwO8Wg2yNNulCZMsyJ7DCRczg8XxSXeev9
q2Q3A+uE7Fklv/UrsmhgkHfUh57NWT6slqx/1x0fco2GyPUv2erRjc4HivPCdeVc
lNTi8oq+7lGY2pjlSILuN1GT76Z6wR8tPMrvNvdnL/taySWUiCnMEqrqpyOcDeuF
rsQPg98wy/mklUJlf1YHkLXr4mTM0A4DeIxgL6GTLo9+KdZIZ5WBG7+22i+ilcM8
qyKbnhBOiwrZzDiV6IJexENiPFS8lxQQCgT7e33mBH0forh+QkKz3R89ghtZ01LJ
q1vGFZKhimJ/O87RqL2sMFtmIHMjvTxzcf4DgCMgzIctdkBiC7hSC/NaL6UzT6kI
KMDXzYK+FX8Lgk0b7oYeCW0+Rq7iIqgBNlYcmoe+qxYEpZoxq0Hc/rDnK9Mv1U0d
a5zH+C7wdRkrAUQ+1pNZlTi9qGfN8G1eFXoTWLsn+wLa0tCXaUB7/bAbJMOs4++o
up+BN5aofbvyv+kRdI3wJCV+5LgqTCq7uaR2dvxR6EsEmfUSeFwH/KwQ4naCu+9i
W47qbDvc82JFZP1tyUQGddKWvyMh1H7XigZohJmG0Dr3laiLvjXeg2EHk44AN9c6
D+6PrsSZqeqI/Phaqece3TrBgQQ3H18lImEqhnbLLibSHq222oIpBdWlX18J5e3N
I0kcLC30XaWdfDaN+XBhrjGDt4jl6bSy5YMZXPknoCakQvth/saxo1CC3DZmnYDE
pPtKlCIliuEinPTN1y0bofjE8bzkgzzWlJYdc863TwB/D7lfMLeNxiA84KzZ3pO0
Bl/GVXsvrhhzQCiI2fTns+3V9kWUh5DgN7RLNENWi/IrSm+n65Ga5Y466Lx/xQcf
I3+U90rT2yUS9Z1fvZ1a1TSZRuDWaFl6QoEziU8vSh6Ko/LZbXqtMHy92nGinqVV
JsCEd658LzjZmfdfPy6mm0Hh9cNO/VNrZO9zBSrk+uBx0G4HdAgkgwa/APyiYbnL
psT72vnyBeajXwqZ2KKA1tv4fyKism10SbwFhkT+3zeyQhLJsQPSe3BrjkodravI
plkQSiy8EbAh/GGpGkGNP/50jTrdnCcua7OqG70v/sq2c8L9sUYnWFMUGtA80Z0n
dJf1rQE1CfaNhcH0Rz6q/I2BNtAz/G40bD4/PSJeYgQtVseCP/Jz+A7/Sf0q2ePm
0/OerI89WpndrVakc320KtR4F4J8JdySJeyokEvZL0X+Qe9jjo5cbIYQwM8MIaIb
AsO/ETRlQsllB0YD9VUNRR2M2cToc4tZlVh4o2GnYE9xVaEGHXV55Ls6epoLzE7A
PHxMbDeUli4VkScgMNx+5MJ0ZNo2R4PUGc1OPHJotVHC6Vy2vfQ/fL+ilo7zN3ZT
Iag2BTayt1pxucsYAkDOmBwS7RTqRLH3DWivglmxhZDj3poK3tib7vHk5nOf7swL
fZ5pa7NRDmirwPW3I/5j+IQAJXFnHeoas90hVYde7cLchrt3p6S1q0MLTxVXsrSf
BqvkedSK3drqnD2kCthAO9BCP7FqojGHraQLdfYkSNXkpqwepzJyCPsPcMjcHUXX
0VMkYWpI/FB1Z7k1pCvVIf+kdATyFTs1aL4ULOq8a707NZXr7u/bufTdSqEoA/S4
hYIhCMFcNKG531M1zfkYEm2hIZm+0LOI89CmNITRjLwsHvpsZTxInI2ytQw7MhB7
1AOx6xBnHn/IGo810ilXoco3W6BzQGnOCXLxVGLLjDzBxbBFCkix5Q+6eMUBgmST
ve5LdFHdL7QHcPjA6iyXomVJNg9QGymPOBuVpf4ATSlPkV8c+4gy7nSmw+sflXKv
z7AZgHSsbo7pBj7o/ZR/EwKgvJ4+F32x3wFxKCdlzTE/u3xWLoUxYA8Xb9sMZ+vA
/dHNyhxQs2dyP1xTWASVcKUofZiOT1la6+UWX6KUzRJxCP3QcCbaep5EokoX72oH
SJYk+KFWNcFEFs+mQdbByaQYX247K1qJ4DnmOQ1DPId2S2zPlJgOSVjLaDahktSQ
CsMKFV9TgONzMPMiyRolDC4naebLTEJr0xOpqXg2z5ISZwcBEvKypW0ZDN83rcWK
bxllrzAZZA1HuYRhtWjYApVQo8iaglEumG2VuF5RFAk8bxEf2/l8o5JLDP6mugFP
WYh3uE7kdsHJyug4P9CW8QgUBLFDvINATjvctV+oKnfEW9wlpbDlpwBxPM8Gd5ZQ
SVyv+ltcr7tDRa/AzJYM1wYFnZvcx7x3WgHXsamUL2lHwYvCE4S7+4Ql+dK8HET+
/qhmBHnCCDlDqy1NgiLomE0qZS5vwaOgvDpHKvaBjpM6DMfLCv9RPc8nVKZPxQGC
DEwwY2AH3U/BucubxL/GOxnDQ1OsVqzzqcQ0WpD5oDpu0rdo5BS1VYDFYGdWZepi
kXhKxF/KwRSiRGvaWz8BgikMtMhYIsyNA4ZZd4nJ2n33fygY6J/OWIay2NFPPqN+
C8AOgzvZ+iCPjmE6eWKBKGw7JdQczBn+CFBzLCLtFbfr4nsKL4OROAPQk645EAiQ
BbgfDe/zILEgrGBjRkNwH8h1O7gn21pesXnVhcW1R5ByIDqgY+LBX/tViEmm41kI
e/ab+NZ3IsRAlzBWK38bgwTJypnop1Vq8G2IYy99yoHwDtL3Ix9bE3tjmNwQQtVW
Q6D+Blom6Y9w592NLoDOvbuQUzsD7aQUuhXsSjTuNffaWMVnTgChxR2R9WE+VCj+
joTOZhrDhjUiYxc4zZVPpQ9gjm/ANWs35tAtM4J2qrluRmMg7jvTlNTvSfrwuhcc
vyJ9pF++m0k8VLnJQNkznLcq5GrvipcvwHXOTxDwocSw4rP2m0VZo4HlbHOyec9T
mq7NtJ7nkEd6OnuGxrrkNImP3JjmBD3QWbxZ5/nXwRtNTxMOmJWCcaKEME62PA5h
9cRLnmfCmBfbH/yBdrXGNg6FaYQdn+wChYfALjxWKmUg4/BqEKeTWvKnD3465Muu
wH9br8YsFvYdfRwmoNCSmQSXmoFTTrbLAAU+uqNESGhIkWThay0xjRLdeaGGfC2h
UvQPGBn+RIkdDuwbNhkJv+xfwcyrC4UuJylEad/imvKmk7xb60tdos2qNx5+di97
vb5GRDw+Av2ECcjTXx3st5fsf4x9Rg2nirJ0/mali312Rmv6QEdFmt41enLVcmNL
n9oZk0airBjpszlGHtte4a88C5oReVV1Jg5e678HAwwFu0G/tr1x9jcfD8Far/s+
5W3tZ1lVwfuEETD5EJ/TbByuyoyU37f+Qqc+K8GM4tJJQosK7Cm8ZIyTeyHOO5RQ
p9lUXIIDSHzLrussR87ZCzvMVXpNPvWY7/u7h7mzC2i88Uujc7SsNrHhCeHMxGsM
HPVjqinQQhmetIBvsPotlSUQdlBqQgysefr4Yp6HHJYU9thUDOZsJjbXZ+tZcSx7
JtvW6jOGkuE4GQI8aXtsGygQvgUo9qHQn/TYL1t7ol6EPpCwyY1WiLPluoI+G9FD
hzrP5VfVqdg6VicIAfKmxW5vh9sEM6kntSp5adjk7sJYfP64NZ1g47mdD4VWC5TA
UgIbF4bORSUW8hK8bE7x3d+iH4U3gQQ5GE8aqUY1rFgoagxdy8CfRSS8670wRpZd
JxaOnYjEu5UZKbsUcwa1QEzVk/EKF09/OlkgcCgofQEUaPDN78WsMK83jBShX161
BeWauJ2epNIXCN5bXQiIPsCz/7Un4iN147JqX1bvgdHBbkhBx/32J9IKKdtuD7Gg
NXd6+GtnKYUIroxf8YechsK3ti9/hk2c7/Ijxz26rasOVn6cAf8610flgRdNGn41
mfPDjh97XXWchH0vXwo4645xKv3jxdJYd8xfQfurrpS6oAf2y77WrJfEur5smqxp
7/mVo31rCMKJ0ETdOL92w1zjtyi+UdOw9Kk69U1DHzQbRyuQq+Dq1qGu2FtYQu6L
D7GnG6w+xJNOTBwEHZ4UR8vBVWTbyb/AfuzY7x2BF4tx/hgZCFYvQ0VneDSFOyMS
HKdrY4ZDZ5gWQUN8cPWf5yS//umNT3rg+jH/+9ALX2T6ufswPbCvEL4B+oLLqM/3
OsmFCUiCM/FXD274EEOjfb91BbeukF2u+hI3Z7kobnAbiHmARRLYYLP7zPF6Wd4Q
bojqiYqcU2WAEkgteuz0tJAlqryQ12Bq6gLywtZyyr9L0DzMWGmBjqiYYUtst7Hu
TEvqUJH1W6zu9EkoEaLqbH+cNBIbFBFtJF+f2QxOPZnZs6TIE8FCo844diyGAxyn
7r8DVjwYUn0sZiweeShvdzs3p6doaIiuDdYkoHEugEEk5gsm3DiHNJ6KHoKYbbsn
MR+OEGv3MBzNlenWMC0080Yyefc15y+IvtS49q70BlVP7coxWTxtA07YCv+IFtXF
xeHAPzmiHmtb9EtMvoE83XbzoQJo2bTFZqNB3f3Y7ho8ekokETAfoOSai3Ofhilj
s7f+Kl1T0amT5WzIoSbx/p2zDn389arKcD04FgfZ91qLB2bkke8lsLSdv60rPDnE
X/AvpZkytooDVeeoafwm4JH8PS3L5CYZ9x0+c3M7wwbgbRB8cKvgYu0Aq9hsRdC1
x3i6G3+VaBHQzAxRkKyripjvBRO39B/devKo7ofOiuhPUJZP/+gnw5ku/BJSb8dx
7XskuHhNCetswM30gigp1CzTeWnzB+Ofx9z/EGb0RvgCgrKO7Xdi3GDqduli+NBe
h9T8mrKLP6qmX45ed5AR6sdoLG24PPiSTogq8XLmS15EU7FIzXUcOj5emfuH0aiQ
bSqKTsA+KnZXd/mLm0BxzpxkTQTlVVIg+Tt5dWaSRyTwPnzNKcBoC0rJ4iXO54Ce
Qz5wIu/tyT5WcUw+kkTOU/+h4YBT/F9yPUnxfS0sHVZFnY1nen/wFz9J3pFawW8C
HFYUJUqW70R03tbfEmDFPiJyxcNAM3N1pxS3LwYXJh1pArKZsO8dbmkNyE4BRAfn
1asXtS0+jf0WiItIrKbuaUAGyP3UlpN9fUjwlLOqJxqStZMwqQOQhaEMkqsSH+n+
jjYdXHYBD6tbZ+bkAFtAoquBbsTIWtDCzDucFAcZyfiF3HykGAbOadTfIzs/G8UQ
bVM823L0pk/q2kyzwSV8751l/mn7/JMPnklJcWEoas1zTaJWsMm3W5UQi9Q16gZG
a3VdmHVO8oF4EYYsYLFOyL4mMsPXMfdg/iFPZlx4PNpOMI1oVLgNoxB51Jr4HehR
s9Rxt3DjyPBi7FM22Poqj9Zy6bgXXv0DAGafa/b9QOhMHPTBNwa+HEznXC8x/QqR
/gq3rHHJXmgGhuEsjCeG8ucqFXYmWG9LRcSkwBpy/p4Q24Ney0Fn8rndA7S1PpzI
FWo2EOEtu8/TtwYeL8jfEE6LQMTbjhuu3eyrMuXQxOIYPtezkVtiC+eLgX14VgSR
NVXdZNYOKc9g9NC3r9fEJ8ipKBacN2xoQ858/dyuW8/Jsk/82XXwp9z65OrK7OBe
vh+Dtjc5+qkBcyTcekATdLVa8H7P8+qp4wRB/YchOCdFpi67Mndzvr/snV8W7PTr
wOVPG4VDQs6vlsjuzSoQ0KuBzzJOlGoOddEc+unJzqrcyxyisrIx5Eq2kSbDjPe5
hVNDcO50zGqcTTRoOoBRfW4Bv01622H5Euy+rpTNprzU7/eBlfUPmF1JB1iVukVQ
q1lZfVhHcW31jvJnpjme+4bn675QrA4yrFcSkhRPLU7p8Z6pNEv2+8Nw6N8zf4XN
vzw68lYpBeG1G76eXxiXVP73sKvC7XYtJC9A01A4aEg0EP05/3RSlKPx1BeH0tLK
vMV6ZAQGxFwmESVKPSYrtQpunWF2tWtarTYWNOzCDUTD72mKroCo0NQjjvNCPxOz
3J8lMwaNlj88J79+mvmIUm5G5Rht96+5UquddjW/1/eY886Q55HwPrcmSSl+c4vN
MSKWTisQB/hnLaleQWqywh9R3AkxYJbWfb2JO8FMWWayxu5/h2aTGhA3Fgg1Kzps
5LlxrDUdMgkqp7K8sYidKzahkB2i+wSiK2q0qFmb4tYgSl+JVWM0HcmqvQ3FuH2j
ysdHJU7WyFd3QuIQ58ThRiHESBaIr1EaWRqKS6dpCyZqwZumhqjh8eTod705tcXq
d3VPllfLWDHLVxm6/txCkjre2TAgCqDow/8H5n3k/RAUqX4sl99gQbSvlXM4P+e6
subs1JB7tUmlb+a+r4AApo6BtsB+jNc4GdL36fQwZjg6PLfkm04zcRBRBEYI/tn7
uPC8EcLNoaj3sS912utinAubnMYa+7N4xES+sZWEHNYIAk6LWc1UrvhJFppLfuBM
TNDKNz1zrrh96MXE/aBAwFoQihjTtpAs3yRxF1u4upikz4j9zkDjU7EthqTfg4LS
v5j36S9Gp9OkMyCy9Hge4XCKEp0gq3gL9Ng8prR3T8MluYXZLF9VZgTJseAcwzFV
WattkiFa/At8+sZGe7SGqDKzS4XRk3Yu+Od/Kkg+7FsWLxWut+31ndCpDNTyNxkV
xEoGbRsq8EeEDGGlbQ/JbBBIuTPvbdY1bBjv4BSUY9UTjO4sfbLg26A1Z2PbfpUG
6pdo5FYe6oVZVYEtfQ3jj+5oPhEUwralwXqAiFTMZLJ8l6Brp2Mgh3NVAcc+X6hr
6oWvyJwhiOI/jT4NhImj1COa3HqgsHU2cEi7zin4SqnAXdXhsk0sIl9wSfMuMLpQ
DqDIQSD+rMs6FLB3QjdwExxM9VkVFD2Pw45oEUMNbrntmg8LK2EKXter2C7u8dPu
g8HExogXIIov8bdHWStiSdQKwB5na1gajxBY38atCERJ8/br4uybjCBgooc1sDSN
TeVi4VbLBxAVHbDunz63HTC0OoapeNqc/WkojOrQ+I+0NJUvIjTKIHGzCrTygqT1
8pWKc/6z/vRpkGANJQIr2jsTX8l/ha1ww/wfqD7lDy7ZTEjQeKlOToNv1b8riQfj
PRLAzenBPAQ9XHBCkxproI+8YsqOHnCis0qPjmuIzE+PWni5Qe7ftBBQqGVJJd2Q
WYZkdjB3IhmpfEpqnJkqL0dsKZmCCHl45pIA+F71H9mDRMPLiev3/SFE79FOzpyi
GorfMko+8q8/8KPUVWeUL7kk8pncn8257Spl8XCoELL0w7Tz1pagi5jN6016aeXp
FUScGCY1H57ANJRHomPukja/0CrhztQa6zMijhlmVU3q9RL09b+SoakaGbCO56xC
+wZV/Ia5KipV0+ibBFN1svOO6Uct8RFs/0mTs3Xs0cpv2dgY9U9J3BLuxYY41tDo
XySgSxgi7fJ2ni82XQ1HF7BIK+Bw/T036gctSVVZQO+dxFiq3xfw/bjXOMs/pqrp
fBNLtDifRuLg+ipHYr7+nNHOfn6qJtr+WGVRBBfobUGM71RX3YT+INrVwCQ/LG55
D/X6HDArqg5x/8PGcOCmShhRz76v0ruyhWxnQw4jTBfJ9OuBY9QN28acuDV2Uqfe
HYe6kJAUNBpIOgVqyzhyQsCR2fx0VAieQcOj/XM1JQfEsbiGkJ5jtedRXCmvVw35
KKMdHwObVKw12GxvKFvd//MdCJfaeqyjNirPkOlamhsMSlcVLSzXJCd3pOtCIqVP
T6jS8xDGqQxJLnUHDwsFRg89fPv9TAbSxsV9EB6ktr0m5zDzaTs75T2qzcq9rv5v
OrAHSg7oyGvZvI8o23FhNVTRNGg413z2J0DNyDe7duh3JzCc6d+sFx3aZZxsC8Hi
PCfFUsZRKILHP58iq+J7zgTfsxv/soKit+vvOU/kLnsCJtMkCvrx6Vqo/gX3Xkj+
S8Os0dbpYpjp5mCykSZIL/qKGnjUWirH+HJnITLBBXyQOu4a/b9zj5qEUw0PhNEW
K+4+SfSkk+FwPk5zc+jM8QnIOQDQRwFzsFYCaXT262PSITIXazarGS1OCQ/EMJe9
e9fmxo8QAWi1Apts+I4Dm+6OE//OdPLroF1V/W6aln60QglK1i5JruJ08Ov0xzAD
+8o7OBBChxPo9LFCxDdUazueC/dlrfN/U2Dci4iSlon9vhb7nPBwSNr/qLzIVN1J
t0iRjJ7g+uQsAA+8kgn2HihylDVj5OonwD3O9BMrB9I2Z9/hXBwpO7KE6hNOjJNn
M3MMA31tCxSgiQaG1e013qxZQv/JS4BvPnHfyp80uVs4Y+M3352FLtstvFH9pvtV
10tCYROhdVDHPQLaXNjucmhyyPUQUSa1KOxrAOeD1Fd2RUyA6kDxlYiYW4EjHPhA
ZDu0WwN7s4T3StOrJyLUmHRIGnODPjDCIomfKO3cet2N3tKGcCxevIntWOpdBDnU
gNQiaKSiPEvI2v5umdTUMKl6kst30I4Gv77M3VoMMdLG+946XEg4i+o6WDIWRY9m
tsGtndYQtQ6UodAz6BF4T2AyYAjvHpk4Y6fqPIy/4DBgLKg2z0say82YmsiHqEi4
ynV4RN9sjrWfZwvywobzsihwwd1GkfEFoDkW1O2B+Y/Q86w9AsAcFG6DbhE0ZqHv
SsM11LDwJII6cjb4mW3gYVmsBKWCxangeoCyqa0N0xxvSu9VdpIDgrHTmIlvzTUq
imIryEjVHg/dUhqtiudmPB2hQV1ylbb0uEVFXdcA0M3TMtJMB+j8Rio+nJVjcbep
uym86p8mTT0Z5m3aDMInrDVLi/FpxH1fxhVkYgA4jVzTO0XeEXEqSV6GRj0b/uVN
ymh8rPdvtfhzayYQTXu5zDw+29SH2S+scEiMtCqTG1nUNibDWl73U2GL12XS/zOJ
ca8gwDfA+Mj0iHHgfOG6mccLV2ykbgoQGYptyLo+4/5RUDcUKEpQj3GG9p6AnF6j
ktAzyIa/u3h5ij01BpoXN4U+wT/8F5EWKS2kHRMcsA1mEbABN/81/f7be4nXubFd
KG2lvqxg1tc4pBHahklTH0RYrBzT6sUjLAGZMONhX8H9uINk5qYoeauExqwk3iql
9mQSjCcbG291JLkHooqdVncyybu2aDlC0MiWnzMkgF2z7kO5y23rGl/ykPF8GELX
UNq9AIe7SHZKByXKiC/NxFx43t0qdPIGUSrfeDzY13v4TdXxUL0hPNFiQ1heSGBI
YKjhNRa0qcVkTf6+Y5ish3AbYwUR0XT0EImtIJUj2jsERQ7Mz8Gi5BEWtULqVjOR
RIHtF51vN5NN/srq34vjAZzBhE23eDEj5UzEzIgq2Ntu64PQjbSFFF/YxVP+L7d1
tVHdKRPAE+cNvpvOzfWfsLZU04ScWL+Z9dYJ/Lh0sYINhG3aN1TjtILxFd210nik
DTLbRgRPmOHxpLCPvRWlgRT3h9SL9NdnX1OI5gWLFdeIuEXEp7VSYZYKZCtVLRNu
KkPqERPrTc2MCwe6QKI0HBEQovBzQesXzbcTFdGu7ceN0ccPb4cBFCA51WqC/rUF
HMX8PvZo3/KSpv9HDzgWqAxDhVzb7kH8lGx0d3s84geST+w+zB53KIfmq5cIEsij
ocFYTNot8pF41ke4XhAnko+LtAhh1iV2boURTG5a2mKgTyvDvcEPlysQzyFAGr4t
SI/zfpJUI4iz4Njx0E8Ih2Xk9ne19TIJJ4i93h4YZ+bzURPI65PY1UtT+HnURaoX
7+6C9MRX5li1/wfMTlqlmigYpgCG7W7SP+g/DCtkaDO33CBIalpVpf6uGJ3LkzCl
49MM5rAQGs/M+LKcpHg6DpjQTndTZGKHgphYOGilLXiWwG+RFqtsUoQdnIVUmD4N
zLVTxPJvU92gwTTXb79v6sra/unaPoedZp4fnz93OxCfLS/TI/WSNhlva80XuqZ4
naN4zRVc5ETJnXMeWJKJ+KxPal3IriJDifS33D+inyutGpfCwjn5dlp7kzhcuCfv
HSXx1pB5kxWMbuZ6pDxVXX4jxDcfaJbwRWrGFYn1n+Krilvw6TKkyuawRsSTeBDX
Ek0RRvtPobAVgW4Qxzepodi5j7n8azrCpuDheSddvelphnJG88m5R7Mnx2rl2G4u
mrqvGi0SWEfQs2QQqb8gXYIeq5bHfEmPDC4QRF3LwfZzZ9LprX9fpSqOvukDmkkW
K7PXoZfb5+GA5Cmi5l2Zb+FzAmvszar3SyfklCiIsoWH5CWbd5kJXcNYO2MteK55
vbCUvu6PxtRUvBVnUsgUdkFUHeNjQtpJNle4TwaLnhB7NQS9N72wo2e3Whu/m4sK
ekwMj7CgCqCwhfBAFgglf2E2Mc5ABvFKWsOT9jDcmRGSie7K9dz4E+AVDfvwu1kl
DBJYNMoImKhWvb913uQ8LxZAdDsqt9N0yTaBkotHMB6u5UV63i1Sw3Uvl4P6aD90
uc3niNIU0byvQGSWQr0IOHEn6kwmfmyIBYkDcgo9+hCWDLp9QXykFEyrEMv40qsY
8ybT09dIVcdq1QaU3LoPJ6F4hKsUgPvqw1UQm8IoiS2G7rRcdhYAqhd42Z9JV8H6
JPn/P89G+cYUKayu841wy0NoQnJVO511Wkz62My+zo+4lqKApD+fjMLbkh54cslc
5W7rUqVw+bGOkMkyYZCGhpORtku708MoCcjegJiCwoHJqCLiYt48No70nFGYEfl6
3EfIWmDDVB2PMWfbLBen0C8komPDwAypxfrrRghqS+zGGbzk42vhmeWf8VHUo8b1
DwcMd0FB2zmCv3EeXmfm35Gzk1cZOAIKftp5HqilAOhzTBbNBu+RPYtvcvgO+87r
iAE0J5816/tsFKJnjn8L05FjVaa+Sj+rxyh7pF4bSBtCZ6IQK4s5DjSjGbweaUNP
rGyq0iEIBTEeCWkjQEqVhj4s3Iq7G4R8FqMp1SfWQ73AFhL79YRLl8UnGUvPvnu0
MHqxAdFVjt+w7jRtd925kEdBiCOkxsr4i2HzJORln0vMVd+0eYnmkW3sRINGbRtP
9+ql4AhZtbezRkbAZBahgIIoX9uz8TVZ9zVHSGEKn2PaMBK9HzjtSNKlAMOBkRKq
oG14qXZ1CPCb7Ofcw2pPNVqyECBaffOEJgnMTF8EsVsHArvgOFmT9aqXTbi1gZ8i
+mSrDb6sS3r7BKpyKXdEVwNDaQTcfm+a3+maX7vI8iClOkg6b5qDMuXsaGBdkjPK
rR6kNhV2HrgECA6ZUrUL8VEFK8NWR06ZMI4OjP3b4PxWcrNZef2UtvsKfvVvPXwH
TnXiVfC+Gi+59Pk3j8lX5X3QSp90Qp26tQ5paondSGWlO5y4r5EvLOfAdlEwTN9J
Gv8DamL9s2uyiR5AHcKWN69jD4u0FcOUGJh57Zxi5X04dC8xv0p6GRQY3RTqSaor
qjUi2RjSf9KYHyGSzd2qKgGcqEEmWqevBQZrgOpFymLor+vEJ3s3taDN5qYyQpZt
0yr41D4TsVi4/EK99JeS7b1o5W1l8I65tTPDBRXpNcEIsPr1/tyYAe0oP9TMJXNt
CwJwrW9AvCYhA6L4yKH7ZzrQ6HgeminGNwcJ4avHd+vBsVyEctrkbEsGF8k9pfq7
Xyui2I2iIpcrJuF/ArdH++9Db5/Hjwnz1e1iC+x3Vw6/3yMhj4q9rsHUZsp19A2o
vbq1dhDjysCBbuUiZ6iuHebNc/+waUwevCaEkaOmSNaPOtjNijq4Fcay6XFGKIn9
3V/tsyoF0LalsTjtk63XNJy9X90dMj0FFybeLRam1eLJqE398eLhG+0rVgNlOgG0
qn4rhLO/mQqlalU91jzJ3pQi3B0fWvCzKHYAR0gmWObGAQOgwaoDSpP0+4jlV6po
sbtQfq5wwxlYvaY5+7P4wpvi5A9c6Guj/LZh+WBStdA+vdf5S2lbD/ZgOdjWf3sx
HykYiPiG4hhtKWy4i4VfYhKXXawOTcWi0kIUkzdHFf4ut8cKdKfDqORYg841uD8/
Kkp6FewoSML4VWJRG9mg/318aP/KEHGa2GqYTWZJISjoJcp+HewvdTvamtWa0f16
QfovbJF7jBsA5euvvK+3rLT5Qhz73+EgzhnIt4tb5ieFf6duLT0m/3NCrPVZzlB3
aR3Icq2sbE82ihfWek8qibUnjV8hGTcrQSWlkxT9SKSnuWYCtWHlgMsXzkKCOOfU
OpUw9aZnMPbwukygnRqwBCry5RCg0Z8/0QM4fu9L9wE0z7qr/Ps2pIE9w0ix9vEN
CEbQJ3pWzSVQ27P2Z/5wAYXjDtu7/vnB+njiH6vjc1LCboP4CP5BcPPm3O99CPdo
dHkSZy2K2nkymsqiHKfvRyC7Y0MU7Hg2UuKOujPEqh6XVZjPWayFYRI3SeO9NbBo
THCCTQWsNWCMbgJ3BeP2PZ+pB/BisZYbLjjTBXFVJ7YL6cdUC5KVIwDgKB3Wze/m
UjDLXZVGY+Uq3vKwnlA9KTncJ+uS/nFmM09cp6bMpVBpQEv19rmf1l+I2Fxc+g16
QSqVPJu/sfI3gWLyMYgRg9rtD7N3oXaY3uJuRIpjk1XcSqAOU2JKacJQtHQJH9Yh
j/VpNtlUjLalwf8DdvUXeZdVxahUFYo7mQrWOsCE1vg/IVU7POLlPwVeu0ufDlE8
JagG/dgfIZuIPd7IP1rFG4qLhepT3BOKrdWPYeVUVKveyyJwYEbsPdFYlrS9T1jM
DHsmSG9SGavwo/gcf8F9KLpM3lzYaC8aGtFoPCd20OTwAoHB2mp3RSXeXdG2YC9B
3p4L32TBSXbpMv8DQQ89QVw8a5DLqoShj40tFMlylFFr7CbXiMa8xGuiB24/mdvl
ZC0EaLFqgUc0Kvqqnce1NA7LC5QrAWu+JpF5XRiwiU3DdJUBEE+uGaP/6RgMBIVA
f7LjEcvbMNkAvWLoa4srBEzFKTwHgfOaKIrUOTCqzn/BF2scJg30WwIWrRN4Eb6p
hi1GdfIYgdhcv708mLq9l5NKofdU9ERu/sUTGGEtS0ybSFwBkxZb/h+1gHXM9uA1
UyBbvBDhEjz3WbroxmNazhpTZCM76gbHYL0YtnDh4RVvjYCSjRd4Ls/bOfaiyk9D
y1mxk3XdovUx0x9+M0NdYomMeQu4Oa+LNKQxkY5Q/U9GiiOWIVD0EgSfpx27Lwbz
k7LZkXHHIilJDPD4o9Uqku6+ZWOMtrrD6mudF+bR5GIKXZgAigNDkWGt/6hGQt7X
p0Rs2fztBJSlfVDrBjqslTQMHj0prBCK+QWeuhBrPrEcIunT+p0nAd+VNZXgeMCz
BfZ5s6RXLNk/mFyZWj+0TzdIGbn4y+zDBxb9uqMnbLECUmNasdIYjXKjf2lqSxKQ
ODY/ztfQOuzjgl60BekDIbGSP+J3nFu9JT0iPBXrNdZlMbi6aDSZZ/kJ9PM4gXSJ
/B1WCG5ns8MBlIWF0HkJIf10oYvzMHhwvSmckPXUiZqBMDrwjiRJakvEznYY+UcT
O2bV0XxubSRH2ZG0zBfuRCcXMBvc6Sa1vJ314HkgdkvKImqNEj/yPL3hKEyDfwql
WAFaOpRkUCnhEUlsxTS95KR3ueQzwsJGPlXZL5m+vHjZtOzMNKOeNK0sAQf81jm4
stppqevJ3lN5W4d+TS+wJxC8JA2f2DyvBFFoZEdkQssR9TJ0uBMTSUdXE8Syr+GN
WTze47WZ7ct/j7sLeu/FwSwZTgjeRmBbYmvQQoUlOB4i8Ty7fbi3edaqwNUoECRo
bxO99kDh83eTiQg05+/ZZm8OVwB8QPolqqAjwrfZgIN0NkEdJi+zOIPy2Lb8J/2c
1nGpmo0pq4xiJDaRv101hhsgVm/bNcpvOvYYvIxsFkNF/8/8Y3pRqidUl93zULN1
EzFqqHrRv4YQgF1mDOTkdyi088ETlmtxmD+LBRp7Qsg6l+wAvwJ0WqoJ0oVN9xYl
MojOMkxHGUyZFbZfSrKHEu+dwok0Iwav0Fhw3WP+7pDN1Wv2KNkuNg7Lu6SFmGLi
hWV6eAOyzPSqVccNFd9S7r+4YHfB88YbRaZkeYegv2G/uh+qGfkirkCEBe+LK8M0
H+4MX1KBu77TZBH08at2K6suw4I4Ls4/UqU37MkSINHpyNdS6Sn6J5HOfixneHQy
zByyVH02j7qRoVXwlWNuWDclMeByclJLcPdo+o/gmPUL1NlmeLoDulhwgCbhyXnT
mhtIyL4uMmoEjIxqb30348zCrYnAWwsipgZ8fLTiYxD8MKfOFmrxN4QlvbwZsved
ow5Xa5Il9DT6Kezzst7wlsn1OVPgXefSpUNa4j54vMhjtqNtqrCcgn0FHYLgsBW9
xdZT+hSZxqkWbdVwOxbKBtDzU+ag00BKBVQ0Q5Bgk2K70dlqpluvO7mvyCqQLPcb
oWtt+Ld8ef5/veB9eQHyp7dJyXwyPpNlN8BHZZ1gcVGzY7MHGERaoHyqcSWsznkF
TChbaWMPoh3BwYJ/uicGMwgCNPaQod87SDebZApJJvjFiXyOWO1Sbv2Bi9ER3KWi
ampVXxYZeziC07n6XoHcszKHTuZ371u1ahu2R890ccbCWFTCPM7a2y2mjtXmvvXE
PgtS6SJpb++vQQX7CNBmt+68wzXYeWL8H5mwbb0T9iXBoe4z4kbhMMQY0VvFXcmY
4m614fUS4CqXWMf7cUHScCEs/rtIxFIbV0Tn52QG1SJJZVip+AVuTwcDw+vtPzs6
4LLIVbNzXDLNJ7wo802aPWePnqUpfJ6bybZjxXTcTBQpI7X7qFB14b1K7L+iy4Hw
EQwo5RDvcMyHCfKxCfZROHZCfG6wHLgac6pljb9gMtCM6yYrrGmyMc1JWXdfoC9J
+kVBLpZs6RoQbK8bb7v1uEVRXg4akV9PGNjw5LzgaDtIVE5DySwsE14EyUkM38yj
d06rPLvIU102miMzvf39nvzV4xZ5tVMUhAzWU6ciyvdUyX4I9/EXdLnO+x8duaSn
qphZAyHlxoAEHPS93KODln+16lqRDOkBP2C9ktBHDhczcObZKTEnyLTmaSrWHwCA
CdXxn6NQstUefghbOD6/t3Ido6rLvbvyfczdQ4T2AMg+nJ8d/oz+KjExoWuC+0kb
LvBGHvIBFn8EvG4cW8N9Jk/VGQRX92tY660r4vV8zowfS78Oysvz9r8rp+KYZdH9
ARMgyrRHggE9vNSkh/Md+WDAQVRU82/EFqpcjlthqQvedFOlhRJzFJoPVHJoqJ2G
OPmnCngvQO/wVq5lo2O+xZDB+oTtwS8UQNHeDakGTKFU2j/NVLNAB9ngjgvhdciD
mXxlxWBGE08jLIGJ7MvG6DnyxXNNOhvNGGXFB1SR2OV+63MHA6eWHXzjCm7aAJDV
mOzS7sZBntAMeaEnWdncUN7aXDUAaX/AeF7wx96uNskluyAywN7XxeZIloQIExoQ
hEyVq8CKsZs5zZh/rSyIcfkOGIi1/8AgwZDikzENmBcVlX9pqzaR5+I2S8vMsa3J
fPULSgJ0uM4CA70ANMip1g0VIYSuwIuHjW6pS1mUs6rKlYNmG8EjksQb/mTcX+GQ
I5QE6vjGV1eAPbAkfMN1sDAUgopi9AWUsBocYoSvo2PYMm5cno7f0+YokMm+VNsz
iGHg/r5mdXByWpji7YOGazu3n6zU/NhmNaL86s4wG9CQmZ6dpG6MxtdVfG8/5781
Y3b6YvpkTAA+iOJx/cmVAQxk2rLwW8eORWnHrYxc3mwSvBud6l6Kb0Id3a7Y6ri9
3KjZCm5kJgSDAavi0eG9NT3VJs0dNe6BQXf4EmrDBCjg/f+0rlGrSSRjZqWgK3pf
JA08bS6gwPCXi8IKbt7byfAz1kqeCqS/K1b6fxUAb59R6rbg+UVdbzh1guX1k7hT
HPgJFiqePjjPXcPDm5dang1PiHEEe4vkbGca37P7QSLFD/xZBTvQAXFxnIYow6jl
iezvmpUUvhbQ036g+iVZx62ZAaNyoqRBqIb3UTYp29rUwY9GE7cUDp/mT3ra3LG+
9xpioRlpapQPRApI0eu58OUKF1LlQ5YE3lTVYI8ar1c/mEbKtKnRC0OGR+hsAe4K
ib4pbFzrK4ENnXzbvnyiDCc4cvVdvR1+wCO5kgCh/LvxgYNsYZzGQuJ73imfbFiz
564xOan/uJopPXIsFILppjmYWxFbU9URtxBm4SLwoH13G4jHjznIa1qZe/3gAoQU
bTNl6xg8HUgpd6SA9vsCZ0xbuXaB6FgcE26vARteNGeugNzxdfXyc5I4UkmqFfQW
uAG+AL4KosBQyqZQJ8YYeH/ITTJ0jws58oCJc73ykciG5rXcnFYhBjhi1Y3WJIOf
/W/6OcRs8/SwZbydTvoBMkZMjjQnbFldnsC5cQN7jZmZvhfc6TaVuXbJkdaMAd5D
kzFMQwyUA/my8d7WSYm7ZBc4YpNNDzrQ3dQOiltIPSi/i6tXqXRpaJvdE+s3HdrN
7EReoUuN5gBzOt19ZKeifcRZloxwDB/FXMkI+Zr1KQO3TeJpiefWH81HrFpQ6d2O
QgwbZ3X9zwdATkBR7Tf0NthyHWuUJ+RBpyHaRjs95VkK+fzmB+buIf+HkghnWyIw
3lxriv148QQz2urN5uSKwxL6P1YcHoFjBQ+vMhNlMAaTdeuMxl2GMK7YvDHC0ynx
KY0dju9ZcLl1PkD5p4F++HT3C06uwRSDSebUU+IRFEZKVqNyvsY+inXRgKVWAdK6
3XPEYv/H3Ml1/PAU9UTQjreDhWA4FP2GqqhFc9vRGoDKbdrP2U6+0CxmRdL3bn7u
LJoqD3clqUCRb2naxEibFtRMi4DLq88bAqVSgvNS/8K24F7+JX7SZpjdW89CNC2q
OuEtEQTUc1jhm+4kypkqrIEygicv/J9wko2FflNdTFXfxoJSeyzcNZYmu9PKmUib
elhf4HkN3JQk5heGxraVkNAoTKYVQK9hh+S7fPQWJjwgjm+FUoDB9pV+2fgTFHR7
ABpkoPSb9K5QE4tdOWdiFnWrcdUako7uYQbOgzHkzV7hriEkKCk3TcAITtujZZs1
aqRrDOFxXVBhhEHCEwkwTKLgbkfbsSYqw84+hq/iq0z9v8GT6yUlACwbrbXVb3PK
nBrxk5EC6mn5SJ+HCoxxWWzT/w+1rF9PNQRVHp0b5f1Ou8Tq0SZlab6ElbZNpgzW
cxYrZTh2Jg7Mwg58d602zrCVC+ST6ri4ZTBF5edzQQ1vjxkE5cbltrFliPbhtQsw
WUb2xUBSxgicA1zYlkpcyrLJVSybivUeeNRrM5nTT51Bupofvzj2nEiVETlFKzLM
eFJb/NMYs4n52TG3/hjXqvD5g/NIJ8bydQKCr49G1qESX8a8zitojFDdQe+SQHjY
XsO12PMk8y3fu/LQh4OXt3GOEqC0dGdK9Py5QAPUl0WF8i/kuHVnW+IXi5h0QiRL
DFaWfmhNOQdd9KO4YWYVhBvA/W939QxzquYqsiF8ER+D7jnakLf2q9cpuTt6ysHy
PnCgng/UUES+54VPjPR2Gi9GM4VCGB35yAOfRZDXJesOUxNIF+PRjA1EbQwbS9hi
u+uVQyY94hgTgVPMX5gftdmF7riKiaui4SYgBmWz7balQWulDIQns0R823LkyeSU
O9p7QR6At6dMZ0A9qLb7TLViiBImOM1lGP/7TWtL3yUSUhAEe1SdkP94Z/nrSA4p
ZzjWbQ1sR5XcyU0jhvahBvQYx1wVwd0466Z+BewJH3NlXiCJmd3+tEmvQdx6LwH5
nHMxsuuWjU4WmL6hUQL1VwMiNCnhkVIGFs6AJztH9HGpE3r1Hu/AdG5CG70HjFaZ
QTKSOM5lMz1NCuy6aAxQDsp/rYDksVKrFqUv1yrWRFQr+lIZDX5KwoYWoeGKOfkI
6Q51zb4r71uuRVyTsGUIWXOLEnGvvDyksbiJ2iWOF4MPYXnAeeBHcefqydF/aujo
4U2O5fTgA71cBcvNgWvWjdGXAVcjMYRppkt8sPgzQs5WX631IMOC2nd6izgA+I2M
KVzyQH51j2MIkqB+AE+ZI3L4EdOTM03CA0XRj6URwGlHEKR2jGXqmSxm4S8Jr48B
r2ZqO1MRbyZ+pKsUo/1pR4gHjtKI7vjQ0gKRMzmg5EnDDdNAttwTtY16U6Xds5KH
G6ztoi+qzjPJfaIK63Is92AuoikPqfo55Slv5pr+0UsTf9chhw/mCPO8OYVSdKyx
q3jiZg4IRyEYrTolVNOZLgpsElfuW3u2vLvpto9Z/4b5+SoK6kUuQHrzDsn7PJwi
7HYoblOLwP0qkdbDDoaCVCmbqxHAahUWgE9sPn/CakI+qiUMOpNDtDsdHtQbinlR
X6QuijLEdaBvPCRDVrAKMpcRBygfoSnjnauhWbWLbJvyWc69fL/8TEGMFF2B3pp6
RWEKwZLy1rKTmTlj+J8WhZpJcsjdx1UFbG7xA9Fw4cTaiSdptB0LP2NTdDWkqs3m
Y+56gZwBdDlWsH5nvGhxVJDRW8ICdS9i1HDSA7FLm7e6OyB7FdIhoXJ/m8G9283q
qYLj7nn5d4wQ4F/qCKmDaLv8Z0//3nKrkC70G8XDwDI1auABuFT8JEAQQsr3gOlC
O5/PziuOezHncc4zw6YNdfFKo0Xq7FOMNZOXY3/gsn8rB4DTQXd+IwPY3eqN5YxV
51/KwS7k3J4qWi9mMYXl6pzUvUpneaHSWAxkL79ItgIhJ/5h8Fx7f6esDPXuSmC1
eaKSfBrIK1XQGuMXc5DEizAdZdCYlSBo6qmKlIHPmSKn53so8yV4UV7A0XPMShTQ
9nPKzDwAH+Uik75fNaNJ/M/Izh0TKkIHg/7Wa8hPOsvHkBbxAWpgz8jWl93g4sqy
QD296+1Sj49ayNAjOx92OnLCmcDBPFIOnZCGWJuIIwPqNoqUhJbl60bR6/pClKRz
U5aDFp2X1jyvHtZNQnOrsczNYDMn5gR4aaDftl8HJfaQqB0wfqRUpRg1j4XpPOTl
U5hevKRiVCM4ISSTTK3g0CAYmUuCztzptmQWgPMV8CH30ljw+PKjKsZLqn+oj50f
DHxOZy/Y9DiGTyl37ybcbRkhNvbYxnQIJ1Y84CxuxwOrgdyjYatxNU/vWqW2o+of
UTf8TYtOvtllCgwbSuYwAhS5WdfitqoH0axnxaH1dvcb5woFjkrwGwE68bWC6sKG
GXGDz2rBswwKSSNpIcoJxgHW7wUOkKRYVj/LcK88fimHWebI63CVg/AmkagOsEL5
KClZAzHsX7hLQ9k8q7kWlwUPNp0CL3JaXif+bsYCuvuNILT2gjRUfeHdpSbLJ75Q
wrf+BN94Jl8GAnb50bC9G9+HDL1dCaOowyXlD7rzGicErt+iX6cTFGuRG/QQaqLg
EN2NhRTC7tsrXnhaGoBUgVZQ2RB+WBdF44sTK4lGVgC7HLaxFIz3SS2pPbkJuWyy
Fcjr0Aq3SLAzq3UU9rd6ShnJaCsScuutW98fTP2kkUqmD9HT1JkvTy1JbCFGJet5
f1rBRK/7Inciza53QLg9GXon4W2g0Ddp8HNeZCuQQFW6hxEcVQfDttLNYP4BxJ1y
Wzp9JwdevnY9LbrmWNYN6b14Pb6SkKAoi03UBKxqBQpA0aQxut6+wNmICeisX9Q1
rjVbxHqzYFFMGPqahj32vhyu/prpBqsUooKlRDAWMVYuvwqrB7b82OcrdPqPlmDV
EIHJaePuo9FLmshfiMy0szejSuVEVdqIS4gDUci6+sPmdvYF8qhFqDag+kM5j4Rm
NkEcjYtZ47cGzlcksHGH9UY4uOSku5HHx7hGuiF0kDmE0zgVh3LKcCZIja2b8b3V
B+lQS8iqARRnEsxdSlx3WGGI8NQez/rJ3lNVo+n6XVnGcvqfU/mgJrZ0ZeQFdywC
2HUR8G1n/hKj86+pxtlye8UxG+I7KebedOnzE+EzKO1+J0eN2OzH4e1qrW9m85oU
O0IVh2QEtm6CuWQP2nit6kId+HX3D5cEC16TFDUzWQTwrBK7SSkU1gxX+0DSdihx
mH2Bm8iResK27PccDOZfsjyEQBHrOPhF/es3HqsoJmDjfMHAdINBb9xwxQDctnXR
3Gy8mi9E4bbWk6sRfaveKsIS/WrSb7KdJMOaJ6DQ2W2Tmrpea7f6fSzmSgLqZYi3
lb5hx2oUvlWSsx/GOEU7M8duZ1RooqVO9SwDJQQzfnEYJb0r0sjeCagHGehnE1la
Iv1Rl73UGQ+LGwl6lE8H+FQ5Dp3enjtFXU0N3WV+v11z5DvUhJ1dnbM1MtLA1hEV
sOj06lqrdpsF6haa3Rxsn/KTTCc3Mzg7hWC7FR17WaOdVgPrKi59SGUv1cX1effP
Il42ydI6dtVN4WSoEnfNf0jjUrmdI1PIdqGgVuKMp9SdUZVd+SmcRUdpvVqs7Pg8
T0h0SLy4nTJROucnQoAabf1HyeEl4/pr3PE2lm87RU3ZGYQd/HBClZWUmQmZ4/Ui
qci/4gGNkQ3uerU1blTjXlwXzOLw0pWbiJQaU2d0CKvMvndhUdT5XJ6Q3PGaoG43
fmthR2WMR/SafNFFtx4WS2AmON1tIWBIC/Nf4y7pMcTEziCSvYJnB40ph+OKWWnf
qg1iYSMWE8ajHJKK88AYCkTwVlsaaRcHM/JcNQuyuICW8vfs0/Yd9txdgemIKhFq
eSq4dqqjXniXSekTjV1Qcatu/6YyYTg2L1aV8MQZEpz7BgSBMD6f/vS+vvfIrY1u
XUluRF6ijCsoa6XH6ffcLQ9zSmHfn0eVM9fEhIRAiuksyNPV5/tcY/6do95nI3sk
5GsGXswKyIQNxMBhYZvR/mSNRDzTB42vbiGTIoCazC+fCbDcIX2sq6ety/dkhG25
CysyK395jHz4Aw5IsuKlvflnzWEvbqCUum36UjSMBflG9lAtx00JT19keTph0b1M
+v/0ftP0YzAvOaHp7plzoOCGkuNPCJF0TPdBFqo/OC2j+onuBEmg8J8R2crWJd0C
icE3arpjr/PLRfKB9vUk2y5ZJ5AM4GhgTiCJA0rNTCcTRQAw3Z6Q8E+jumYUdxFM
RQmoJ+urEsDoGpOphrkvGFVf8qSCAw+7C74IY/ILXR4+bQNbeFm3/6XOjaFgJWZY
Hbr+kfqDxFwBoGcI4h0oMu2puDJPX0J2xHgHito1gT918X98QyH0lOuBoCJ+2ZiV
2W6tAowovR09814hqOL/IUzj3eNiv4bre44NxjkmZicffGjtL+HQ+VYmdZ6piquf
12nwsR07WgKEjiUBQqdOflrIxSntmPLgYKZmwaWX5zGcQA7SSQ525GQ1R7O3HF9H
/6UJnFmgZcdCEi4M0Y5cPMjFFi4DzhSDpPkiFyb+k7w14o70nZzE+/NT9PUJRin8
L0zJe5fj5fecLMK9YZnkulnSdri15ig5mhQsCbZSFnMwzyGySAcw/MvJ8royr6b1
qPaTm1VJJrZmXiLg/O0AEz0zW8yZHjZIqTjigbOj4WKNQYvSU5FhI6VwYOI1SYCH
NabsysGyWNglM/nc0tT5UNNCu8x15JG5pUvADQajwxU48Qn+0nDnRcW2QjZPw8Bf
dngpxo6aoEwkh1ylvqH1UMfmYIf7e5AiZIdRu/clfTIlTXqU+SlinlFp2XOYxSts
2GTCI7Ptn15v/vAKXQ0QQLvLJO+N1Qz0jxxtgiaFsOBfVbIQzXnZtooOtbKsBVYS
jY8SnEkvg0zvQ6v3zEDa3+H0E/XA/snnvfjOqH7QEheMaZt4QpVnqs6tKqs6Pr/u
Szxq2JlOTcm/SdY2n9Bk9aqZBDWyYkSr8SYojCDPIIzD96ZLszPiLmONeyYUhpIO
eY1lpDiMSNrbgSgNkwe1fbgmi9VHMnVsTCnKIhYPVAwLeHAkovDWn774YgwyCqaY
w9ItDfJ3mPHXejhImE+pPZiDP5LlqlsmLspOsM46ZaakqmXzYLLnk9VYYRlQ3XWD
HB+qy0NWB2KcNoazi2z9ySd1lpQymtpaZB8VVbcu7fGW5b2EaNWOkkmzU/9qJsTi
nRpDmZFQfkN1aDRkhMN/6zVITtKxlrmIGtD6u1q4fvVM5AT0UwDSwR3n9IyKv6h3
gMLNWpqCjiyGFp/qPSdWX5raktr6FXY18JIwyGDj2o82u82xgkHDI0cfvgsjwUhy
aiAhJGUM8Tj9ni0h9nmkaCzHXI19i0Fo/jQAJTOPCz4bomgl4Pd+MXQtNoOnDfAf
uBwLt83i5vX48ic2/3/kwR0y7qoR2k2EkTiQBvRSmgrFo58hHgx9IT+Vq8T/yUEN
/lMH+VBPEkY0vV+oQBCwyz+feLMDnjc/njGQsX2ON7ls54MQvOEeIInhKu1vy2fW
a9n6jyYamZZkrskzqcljQd2mGH0JFaaSahP3fXkZ69Natf74cPXftGvQgOK4p6MZ
8YYba66mgkKC1cQO2kXIOvZ36hw1YtLXcJME2UedYzb7MJna7H9lzNxMMM5T+9Qu
VouT8nMeGVZNCH7Zyr3ACgSpEo6X2VSxd37751Kg//Py0BhPbLW3sWtp9o/DWyZh
aemAY53E+3bEUQ1eaWs/1uyTPJGJrKnXLCgic/vFlWyH8xNVTYa/hbj9bYSs5xeL
JIUXe7+dwBhO/RJtlHD1ELBu9PrdMPnCH1XUw503OgjYQk/cbI1Py3znxA5vq3f9
FXaz8KDuARosPfzzs5fuFpAx9uBpvwWZV4qbZLlcIDsVvSnLT7m+I0AJlNYuejmn
LrReNpcV6eM/lop2HXPsGISRdqB0gLJU6ho8w0q1rnGQ9EGHPK/75QAE+oiCwZGN
yPJUKK41GgEv8y/A18M9V4/CiziWJLDradEd22wWMVYDISm9Gbgx5+e7xtLrm2iN
Zm7hejaMxhzmiD7bA8zNQH03Y0ZIvvPIfhm+TsckBaB0fq+RwIJFsNcubuAKt0GS
D670Ns5vjLLQ6XYnWm0uWIBI3g8FHK1blk16thqwZi+9lGDqG3vuSoal/hDPip+N
PFiwDQ/2/w0RCWx0QZCmu+GXaOiCIVdJnNx6z8r3cGehmAzwgj0ecre/bRkGkv0Q
khUY6NxC8CgyN7wxpaZRw2VJCWwmU1cRwiITdQNmzT8+ho7O71Zhi6VJ4fWCpXBI
0seBkiuWyDjlJbXr/Qm+Y9S66CfCsCxKe3OpLi9r9NpuvB32YBG8341gB6I3bUCq
EmH7/eUk5W3a4I6E0VxhrA75tqsWBrM/Pw5fNOD2I120KA9lRB1k1Brnfi0VbMcB
P4ZfMz2dBcArotM+/vqXSPJmBIye1jvTI3CbcK7t0+yS6CvPKRkFDcVfWSuTV/Ut
pk85cjcgOCPJBKbh4Slb5bGgEXHzCAvKfpXiJGwveUvzPvBHpJJEQ+JkCpEq1L+z
4xzXEH19zzt/7oK3ILgy1zxJxuYZXMBoynlIOm7LP7ar2DFCif1m1EIeBWcI7f/K
ZPrW9yeQHXld1eKpMUMV0hB6SaMFIl3oXwsI2xvLKfC9XKaeM+8J10k+9mDo3+a6
KafkfHGzI+pEQuYQmBdf0g2/63aecXR+GYdbBsKJmdaIeol5+3FN2dTp4BgeFwD+
z/ubAvsh4TMapz0GBhHNZfCAY7S0MJe882wuBHIfs7gFiZLRNqElUka8KJX6CDPR
62s/hJAh/eXdJfCM4/6GWn8k8kSOB+tpkYB32EWnpDLfC61OLrBSX6/2wka3BT3x
G9414Ai4sBvuX9gXZhr56iOnwSbzeq2G9MGUkROregchmh0k5lrpTtrZogbwCj7W
rxnsAsjeS/KQS1O0OD5QYlI3VBZlWI/jeMlcRluvC9pd7mNaoWeiW67dSh4gyDu4
lDyLJG/Nkkj4fyCBnNuCVoVaMz2mSNFojKUHFX1WUKu38FDc/72e2tLOG8kf4YDR
aWf/OgP6eZVcj8JJDfwHpd/7887pz2IXVto9ML+Wf9xhdyrA8ltYqRvsj5d/4xQF
Vitxzr5HXfcH+efY6S4OHuTngGEmF9cuzKMsrXIwIL+WGAb1Nz9/AgbWNL7AhVXf
JhdOiA7oLLv+A5AvL1aMgEarNZUPR2DZRJigv3PFcIRWXsTL6qq4c/ywVx2DoeGU
GqzIumjOByTBqGll2hVewktQwhY5hgfQ29S77uqgs6U1/D7p9KGFmiRgKFKtvoN3
3d5vab7US3534xEgHFdlnf07Kp2hCIt67J9gk4xt+4SwHDmA3hPcthqt9LQYeFKB
WgQAHHXTN87kCN4Fqa3MpxL99ZuewswB9NA+preWhSr+JuR/vlvhfXiAuSPbUZP2
4TBSb8J1nzm3rCo4plB7ZAl6o2ven/KDpEVc9aI7O80s/pWMkC3U1FVKXINchRh3
Jgawr9WevaMh95ncEOmOJY2kZ+TFW5j0wj2Qsxe7jMHgGlXk/NepmrJXMoAI+3r+
Izx2eVLtzwx+QEuFiRiVUu2OHnuDRvjThqAORJWJgYzD1XCfPSl2oYHdsXkspiPC
F8LngW1cLULl+Wo8xOateijL0lAjYI3TXTzrpjWwGF+ttdFhm+rHAFqRY1EQL1Kp
UGRmHCFgXZfZgwMEFvnoRUdd9n7p108EI23dA2LlUnh1LF4U/RaLVtBmYo3FfXlH
GMAfDD8nlCohKaH06jX7oqvzmuvg4EfDt0GSxENNReS6vNVJp9+e226rFBZwUSxr
gMLe9sDkmsAFWXwgDrWqBUVBLhWnQVG7eLenpk5I4Q9GkxwIqziNmvMd6hw0zQ3k
Jao4N8Hyibl3cMzLPOAItrx/hMiz+m4T7P72Sn6ZsJKLEGHeOGDVdPkDJ3GyK5e/
N+YqpG0yJH/OwZ6DDioS7AxeD0JJcWYO6oymzgQXMLqVQXP5vJWn0CLHcfAxO+1l
HUZBEtX+qhXAp3TFEIrBpUVHCXX5hE4vtNhBlx8hvt9T08TsBuXLa8qxvGQg+FHw
r9311nc1w6Kwh2NhvBDNQWV882OXJLmh9DafkwUHE8981gEYFa0YBkj860bcF8pP
6HPY51QmqAjpUxHrnu179EKyZR+1P8weseBTYhPDMGNYQkIQEB7oC3aAsMNhOSK4
t7KPhOqlvKq72q4oaGCr83V1tr6BYaL1LxZY/vOBS1//6dnA//Msuv4yUNnlGqX9
Z8b9rMspoeMqPlRlKd2A/K6/2qvocE/WH+btVYzz5v3gXW7C8htL/laWU0bEJPxA
9ETzeNm3Mkn8uccaDAyGe+bC/2kdD11mi0UYbC8ejNvdkgbITEVW0THBWX0SKZvi
AYkBAgAB3XuBeBLU4P4Jy6Gzu/tMy05BP+8b2Y2lh0/eSRk2CqJasOk6QayLyY0W
69aQNLwFzbywrJCgo8wtmOEuTIcJ155sD1UXxYGIl35Vexb2+7hiAwZG+WDgZqYC
zS+VT5un20tTBr7xGtlm6urdL3WniHiVSYhJ81XqUozQV5kiIV6eAopaS40YbHdX
I1onGba8Ku4VGAilBO5a9BnojHsJXGU1myYbBYFf8tR6TOkisAECmApmR54ycr4k
QJB/qaGZLNGLPn/CeWshtznS7u4evW7A5vlT+8nrduGS8jm82rvz+yJ9CBIJDiq9
ohrqrYLrkY2poUCX5WaHS2KsdatCZfvD0DFMdj2yhG1xUVPPOq3NGpkl0IWXvLxV
xKDBUF170Wmby4qgwi40zZapu7bp0AE04cXKxKFXPXMt+v+AghjL6Nc2VEaY4ZLg
1c1HOlTUkBq20St7kEP3z0sEkpJD4c562hwBM4/GsgcBu5w0GmcrpH+NE1TbMv4E
aUDldJKMktzESu9fI2rz1wzRgIX0qJPIzyZ+EB1o1/81cYUI9x/QSIoHfz++9tYN
El9MmzIugQQ51Zc7MM8AlN/2wESkaIXnaeA1pbtUF3W8TYpyKALvNr3s7QFPIND5
WkFBZub0eSNPj102VKoVqVzP47GJi1iFUeY0ZMyKyZ2/HmeMxBEGeJ5KI0bbuVvW
dzK5TF+jQzSF+pCTjZphuyGGbwaprbEkznsh97NKCA7YVlUlXFtQP2xb5deNbTEJ
52RGVOfCTsNwGHoWtEms1AgDkoWCPPgcsontAe6z7pn+1WB1Gbh/6FVUwHQIqjrn
m1jYL+daJf46NPCm5aef+f8QqzxQixyjD98dKppg+kz98REsQ8UK8h7lLqJEjp5d
AjMGYG+0X2rg9ILkskkW7KyCxEj8oak2rwDnsbRBExR9x7cHyUZVNdOTN/yfTil5
rWmineh8iWGq6LTeqx1EvXzSdWD45ko82bywd4fJ6yq5jJ2yx+kvuSYa3ipkvbvZ
f9fujAHgRqIRZp1TWbzrrhpg7aUGICt/QCPt+L7iHLOfNIqL43yCcY3mxWcVIe72
lhO+70EPF1MY8lQRP1C+DvfgqusaAnm5HXj1CtN94DZc5upMxA3P6ZcOLDfXf6Rb
INnfdN8aBE6wgCSv9UuffLXeqF5H/KLzBnHLxoNCQFOmoL05ScSSIVpsD8dnDAOc
aMLFiNngduT2QJEzG9j0osRG+iuSa2IJru0P45GAnZQuCvKKzJPJbmv3BJuBVOuN
6imphiKxmZhuh93GISE8YMUUVy7BX2AycutIWtmlppU4vkf4pRG1xWypmeRPz0I5
S/Zp40k2vjrxKbJLdTjrS4lRMMH72/CdLIeReO4P9X2VjjCtgeIfT4hpQGnfdu7S
s3Bns7ovZwONp3P0WadOSfuSZIi/f7ntWxg4+7PzFg67Ta6FxEbNotuziDAbUjLj
GNVyLBzxML/6SamMks3p+7KiCIHed05yMgdF2dQTw0F3TDpIqmiW7QSb2usw2y4T
8UdNjDO+CEdi+c3twyuxFe3XYVzdqGNpHPWZ46lYqLHSF8NLvjdt+rOgFRnllGUn
M52Q76zCYbFux9syPCpAdq4tXaUrP86FNEbiIPaF1YEOXGjx7cv261JLQuiCtn4q
SUj1sBfksxrfpKHHylnwnXpmrFDRBlE7uM2ttWiGQs6HjKHqyEy5Ks250Lc8BRwA
Yz4mzVtLqvylDdnJwpeUycv9bGpDUSNAId0uXlMj1q+AhetG2Ea7zvFiny6uUDvn
VB/YBmvmjJtCYxNfw4GHZXMogz/IEAoiZ9M/5U02LD2Jy3+D7YyDnKygcb3aVFYE
6tcWIddfPHIuYWAEodEzNyznA3QIga5Y6UYm1vTY1uz/FcW6xGt7rR2RoHas1Cqx
kxZTysWqiKkUFie+b+tLjjGsvygVayb5wFpeUPM9QZF14MCE+Fm84IwrE5AZK+wO
MimRrAa6aYNDbh6i3UNQ79HrxINU6CXk1EFQ04/OTQidqQY6BQ7WV4ybjqzYyRDd
APkgt1IIDYXSlluvTXDd2DJSgtDBukofZcEjeKBrYF/XzsRk39oRThQ4Kg41Thr7
QGVRwS4U0WOUwad3MaTxq644Cvc1RfI/jS325XJfTcQ6pozff8/U56tmAQ2SYTgZ
e1D4+Uio+N+GYdq56k0LhyV24J1Iy2NIQ3LXRu2FY1FKm6ec8Dloeu1znvCGKNUl
nZhBQdBtRNMfp9Oyp7Br9GRIChheumwCClVpViYvqioaoxI+U1PdeRoQcMUY34RT
JAfBec8LHNhe4oa/IKd/q62VzZ5jqUPBTzQbeAP+YYlFudZga6YlW3zkc4lPWe+P
FjkYUHU0falAdPUD0oe9l3t3nNtLUVKb7dsct0/Pp5hhInQnbYCu9ZLeI14q4HUd
Fii83Kb8qjAfy0O4rr4FZkPhYgAyFxtTIQPPDZ7orBzZb1j6iA/OUFwvUQDFA6OA
exSFtmKcOkTAEwqKXRWzrfOOyjk2lAd8oS2Vfh7nQUVv+Vat9U893z+GRodOlMqg
8GLTsUEYU6XdfhEoMIxyZa+GZ3ULy81SapqHIY+cqnRbES4olrJFElxaEl9I06nm
339+PUvsB7+XomJe2Vp00RXhjnN9CnXu8oGFmhrgzT7gJ/aIn8X2xNxX8k9mLiEE
/MqR8AM1R0S3hgH3hOTGQLikGhpAfPdRZBAI/BZbsnWoxvGMAPFgh9LaDAGvJ7G0
d85eUSu97O2Jv4CVzf59HKHLmrlhdSezxy1XSrxgw3f9bELihTWIZ+yiK7CXGWfK
sOBb8i6h3LNaBMQvHt/DZiZGTh6sHrnYbYL2DR28Dtz/HrM1p2mWr5TVd+7RF9Le
R6W6gSjygI27127QNKjjGw31mkC/ssBsAySSQdF+Q9zNzWKJay4Y2JAGf2JH3iDe
iMIRbe4oOE9sdiz8wOJhxOJZZwnKKg8u7nZMvsJkvE9ydHo2UciK3LksdThqF10y
M3GtNRaOPXFU39H+EXNLQ8fd2+mGI8Ea6sY2ONJ7BGhwtlAoCJTSU8UBZLVNqL8q
fxVWo24iciUt6eTUIAEjcKmKjf+FRgHO5IKppVUJO2yeT6yqdwMe6U1713j2wvmc
jWx0DUhxThbcywRdm7eD6PPATK91M6SoJrNIcDs6djOU198AZHeAjbD/F0S2V29t
vWHz9NT6r/RDBaTcohLScVjuVVxYsknjxR6sWBdxxfATrdKe0bMcK4oC+KvXHf6V
F7rM+2H8g6pGkLzGeKkE+IQ8wbPxPfjj5Ojjd3G/Phl+ReaASaa99gT4OIB0H5WK
aJ6nrjwxVSNqQr5oRDZpkA1wGdleewC06XQeP8fXFBLIphptwetczeDFk4//slXt
7DZTMruBoeo5DvFM6iYk6PsjiCAwYiN3XY+o9VT1FFiWGWqoopvTwtWWz1nus45H
jDUqX95wP3qi6nY4ibBxsz0SsUscMLB2EUm1MfTKbPhDDiKNFlGAq8ef8o1MtnV+
WBWh63N1pzUnhCv/ZUtC4Oc/P+FY4mHPtbBW+RbevTA9Zr5Abqs4zk8bPt9XYFl0
Mmk5gBZ3C5HnwyCbN8jGvB/X3MRqwWI9JOztvSJuchcTkDFtvFGWUtVjUE9CWZ/P
fs4kPzcO85O0S4scjddiiL9tmrQsvLPvj4bl8Lc/Rd4uxp17AjhM/kiN/TblwK3c
WfUk9o1yQG6XPKGf36ecd9uJ6QnGP5CFAKeCEFC8HP60JGad5ScZYPuDrTmITeiZ
3Wecqvtf1hXdajN9DKbB/TTLdSGOguOBnGoByijihn5sSG/meIFAYaqPhGHT3Jaj
NjGuu9nq3OyonuV6Kh4xyElLGDkneQgX3o/ON478yp5p5yFQbqfGDQ5Jj5SbocRT
xq4C5rW5NfyaS/NLfzF/1F0x6pcDMbQP2k/KF6xJsYMXxG6O2m36RjceAJNizib/
Zg3wPpS8ubLrWB5MLxlQ/iYrNMENdfNmexdqlh7f/F9BI1vDbLllsFOF5M5xDfU6
QfmsM79YkGP9dDSaSeJU38TvnCYloFOQKd4/nxRjWmMpAEmrSBE44jUtx65AWJLj
tOKOFKZmRofwFhNy+SaeVtGHE+tmlIDZmYouitrFt3Qe3pvMsoQ4dGRMr/WGuLJ4
jXtEo8RimgqkZI00otNPXvzrb1udnh6lt0uH+RYd8zPQn08qb4HUPq5Uw/uMw7Eq
9qKJCO9onr8jzuz5JszwLWjyMIWBTI3BlF8piF29BNsUF2xLneHFV7zfGFE7GeJ5
La658mmgpD64MyrdVLC3PuMrdkwye08QaiDpE6vIrlV2r8yhKakpJd3MsJzS7rcZ
O7c9hIpwInSlpaeqINMhRn/kd9y7mo55s12sUMqZvOJgiWW2xd1ENhnEXA8m/cX6
vjVgTveP/rCGtwnbAG4uP/2edwwmfx+O1e/h9kx61zfcqktWa1Wd1O7Ag+rur7Fk
xH5opqM6Tv3QPiAY+ATwP5UJtZBwXRZrZrYmcZkzztqyGymSI53EBd4DHOlR2v9i
kavjg6JHCy9RDgPQnWE/2q19QHiP6b0dmOWU22ty8vIk3PrInGrganVJmPZsyue2
Nf5ZejbLQ/F9zhqClGDPGA1OuhpWlLDzAtMeocSyef0eD6kJ1poresrbNE3BI8QB
H5wOK0KffDrnAbWpKrVRYRSxh3gotOInRIuTVhmDnEqCI3XnVAXlURcgZYDVjxEO
HLZI0RVUSOF7wbl4YNw7ByY53qgHoV0XREonWNae5qVlpNVAG1BDAdGJnb0L00jB
9kH3u69GHeCJaUU2qSk+CjOuNqc/0UZFl1P8V0xcgVW4Mxpe3gc1f1MOdGw5Su3t
ChB5DoMzk1ihIzGGL1U8vymiQLIlssM1zT4ahej+XNDNcDKvBTVp8k3nd6MOqlAf
SPYEt8gO1WxsxiNdlBA6l7/Qd4mXzlBSg2Evxg3X2ytAOUZmFsiVBtjppvH659mJ
o+TQo7PjdiATtjboZ4K3/C0V1TrlfwuAxlH7iGB1bQa4AzYk1NHHl2I8NuH9hffU
J1wvyfcAcdFTffOllOjlsqkp1P6OyIehVyuyLnssdQby4BN+x+4pU0/cbBiW3cZ+
K7aCi7UarjO6P+u22YC/xnZACbdEEAYj/8LAPEdS1TaWbqTO7n+JxnS3qq57otCJ
6H9wZqhVsBTcDrZCtM/vy8U+mMhtFm1DqjVL/rBvE+pWKTRyJyTL7dTZx6i+lMeL
FyEYfkuMqmGD7ep8WsffCbWip4x+iVuJQLCbMSio6gfc7k5MR9o44HS++NYGwEEP
CzvC8px6k4iTLvIa89z1frX6I0sJI+pjcuIihVwy4lPq88Vh/FzB0BrXDOm/Ju7H
z+gVwi4RWArocb5eqJf5+mWmci/u3XjHnijdjykSM//cew701aDTYeCvMH1uqLxT
icNptQSQI3hus+op2kPRVv5Sj9HL9PaAeUIFbGdGc/jiTxdwkLjDjvtNWEm+gsOc
mtGawM+T4bcR/hDDovU/h15uwh/1tgQVDa5/UpXB4z1nza25QjfDaWNurTP+oXqi
ryrGlSqVxVdlpy8lTVg07JJ7PQk5gSdYBn+v+FH0/CrQc2yu02iuIoUswy6Qb3WL
xTt3b3n8Vrmos2daXBSY2TKW9AA5KzQQfb66Y25B8jLdZmt0n4neBohe/E/n+0dE
cyxlfcCX7U4RLRe3NGN6C+D0KWO6rXB2q9kdFuSvCxOTJJSjRLvD3JNB2JhBVBhf
dxk6EiSBgF5tG1m8B8yurBTjl6LvRJLITtmsmPPezruFL/cnT+8S4ViaETeQ2Xug
dU//UJHBlNqmGZKMxj/jDXXV/BkTB4GC0/uiE2ivmlmDws0HDLtDgQ4Zs+PRz5f3
IktPEbVP9DIjeOiL/JYSfcG9ZrLT4pXQysQD2khsrVjb40MdDCL2yW9vhwBQE9dQ
w6rW5rdA2npEDYHqAWe/4vyskt4eROpGDZ+rKtXhtpL1n6UFWlSOrxiHVPyGPoPW
F9u6RA7uvrQ0XZTeHhAsYo9LnJ0XXdrukCJKUgSPeq2+vgNdZjEzA+n3JYsRvNuJ
fz25QoYsV8n2yH6mA/19aWG4DBj68yTVv2NjVS/kyzkxPjtr4P/+PgXQWLiZIwkw
RqmnnGNDbQmLQF91XHUm4gzaq1T/FOkQlbOgmRoQ7yCJo8A49WCuvz+8KSKzphkW
1pN3rIRj19c/AYiDiaKXz9uZ4l0yncgMLel/6miLkZ1NB/pnCib2z2hjaKnC836r
qBI7v9UCRehTQ4FEUshWu7QrS+66rb8+zom+F6FyC3ttFxEceo1o3cIZSzLhHzg/
jNdax8NBlNHzb1c8wJXmCGkmK6pco/eR1nFP8F9JTR6/ZwSToaoIijswSgxmDNiI
67hnkhp5wTT+MpmVJCSIzWTTb0TL7Sw8V9FJleNkP+IVvp3+eAfd9u9Yhsgs5A2A
2EsXCNrPAc+7Q6PR2U0u4i0soWmmNgstLnUTm7dtpYcaZr0BNVzpud90pckgtKUN
whpbb9eu/x2S47uwukm/jTXWEBFjtPu9/OLPF+Qeq0Xn8/m4W0LT35/CveM8hRDb
1nxMNrNtA5b3AYMkt00JJR9Q13I6797OS7ViVFv3NlZKId+oXCB00zjRK8ovKsYM
NaXwv32mk2HJ6FoX2/+S5CTvVj8mb1lU/fK3YMgzuyEGXYBeA/NgRKfVw/KxKoAM
WDs8J1uL+RZ0GoINmIV8rHpVjZLhJ4Ei/EIiqCkR4HUPZOMTBJLD8Nxy8XEOMkwE
WfPP3ucMRvG+B9tIZUyzliYTlf0BBrbLSV2rDyspTtGPXZgqV/bJTVA9r1LIT8Yh
D8HoKa2dKJkk/eH2s+MfOpM6X7Q86X+ZZzbZthmDPcgEK6DxxYYXr16IO7e7pxFl
i7e5IcbNmdHShwa92ggc5Bagj2ioW57QnexqGexIcSUXwWet8J+VBIV7xmC7v2UJ
SERNVX3fB9pnZwuZ3NQ3zT+j8BtAjyb3A41YjM0hIh7TsXcxmUChNMd2OMLosYG9
XQbEeWpiVW9BGRC9y0baVsFYRqzZuWAoP/1z9Nt5obMa187J9sQkxVj8IT5+Mqqy
yKaz8f/RdEs851RSXX8aEbyJJcnHVuK8oivV4laGmb0wTkYyE8ASHgGI4ndS333q
ZdllsR3ulCmw3uWnaxjgxyxe1VdSON9sDTwl1o4IaGSgt/mHp3GfN8aGjDKwx5jf
KDTU/wsXQaUgaeSOOMsguan2fkY8l9RawWpv/d8nAARTPLjPJ2YL4oM+ISHOmaQ0
Ptz2PBp0UUgw1RPW+D7hyCs1U62ncLko7LM2vTepoI4UD6I0JhCeW44vIPcxyEXv
+onB0KIG5L3vV9ovUAhLRJrZmE0T6wKV2mN/MEVjp3M4j3SorF65famn78BX2XYL
r+81G9gmm8qtvHMDBBpiW2FPHXDcqK5YuAa8HVV4Tt4l2mAGn3EGTQOO2VktcJAY
ycaWYaxUhGG3WITyp0el+DHs4GujRBC6oIx8/11G8Dbkg5vgPx+aHJwmWu2lLPv2
s6DmRkOwjf74LijKqobkoOPUd6nIdBE/NdmrQVfmqpN5Oy6dDFfXgayVEm/C2beV
FSdwx+twwfKMyR6l/E6U1tpDicrK3tXpa6i4LeRENVJDRmrRT40grl1E3cWQas0m
AQFVMSwSIpNGS0z9LDbmdAvPTjCsj0KPUPZwbD1kMW9STu/Uo8om32BbxStjKQoq
rR70IORh6o/UUORbmu3jLIVZ+vuGcNjhps5lO6ZbRGS22vqEHQ6ipA/ucRPHJgY3
HzAhVltxNoaLj44nmoKyK5DXVdoMa+HWi972uvWZRlzeabevK0wCAAZNEhI0Y4o3
3jqKosdqe8q7OPcP1k25KZu5osoWdcjkh/+bvR7QmCKSfUFWqT2Qqr5VWn8yFNRp
6xzhi6f7tE9vh31URoTqACc4QcAuw+BbrOoyFr0wpR2v05ud7+53np3CRGKFRHRD
rBAS0D9BtMBtarLjYRl5xaCJE6KlYnA4FS7y1ChUGKCAnZ8znnY/Twm0ZDvZ4PYE
Q9854cLrEHT1WsrP9JMiZYsjtCftwSCYU9RdgnW1Tb+b6C2av664UN2vkwsyD65j
Wmf5I1uUXIEXEOjPO7voE5227GaWbw633mftgAHH1EdpEKJUrvkaLsXuXwAH/8Is
GlU+EAhw2sxv31d6o/+faGgqUjkUArmBzexSflJku6mxwMcxjKvsybGmO0CLN1ZC
znOtMAkzIqMGfbWeMevoerg0Uz9n8YOUTZfSFxxwvhvGWuwHG8TgM8RS2N6LcZkP
ZVN6HP+39PNp/Iyxnxbt8W8ris70roSpRhpo2DTlO4kghp/5qTCUUSbfAhDmtzz4
dw8QNUK/j+jqHNGYnpzFGzwhz5U75r3HLNyt/arbnPd6XR5YMonmu/Osn6gVsxsK
tSm4n2p6RIa8Z+eiPkKP5GRUrX7RuUKklEm5lCkqQws+BMUCnTY5l/WS+Oml1a1q
EHZZY5xAa+YQLAeiXTgg0g6Yq5vL63KFcou58AWY+tFtIHJu9Qe7ZzO3jDCf2MYv
CRSFwSyx+efjy8peQagWhdXj4xg8ajP/zmRKacH/jhx1GOe7d0xXRErWxZTLYKCf
0zcfDrIJMxHZ+hvDOfQvIFb5utR76DtrxzXOBtCVH7ryRJsL69r6FX59oEjOFpp+
jExuKuI68QTqqKAjsPmRec9NAg7FucVyCNf7BRbw06eVtBXmTPxEgmlhwGH0Wevp
bV4zP40nP+TcDO2xL5X6CyszTIRwUE3ED3eaBDHf0BjlnrnIbHe/Bf7j0VPelQ+O
NqQkMvaP3ghBKQ6LcnTUL/MIgsWplmzugnYivl34m+9UiTRjvvkH5o/XK8FqG9qX
CuGcYlAWHFkJiFw3tAWox0gXp0n610DFEHrYq0STZUUfsYc/a69I9Sgut5uOpdqj
SPs5SnTbywLF0RFOiPy/++QStiv8dWDORetch52wC8Sm21QEg7k9Kh3ZBYlG6bhq
4HEI6Lma0qUW+E/6thezgvzpLl0uSUhtcW0L0lifmDHVIowAA0YphF8BUufy0f+z
2R5NONNmVx1tI/xBeeknJLAlwPIujJI8bGk4AfHmEBKEkYyCu6Y5rdVem31dcFer
Ke8nkWAuAh0n+S6EWF5ZKIclhEHIJC5Y0yIuXXBVlAb445Nr2HNkzMACvCJ2QEGn
pfv75uG8/eptEaJwHV7/c1pmequRtann3ruuzSA/+cNQCVat8a/5yXTCC3LJDjae
9rzLKkUg2LKbTsJs68G2ByMz2lCUHLlp9e8+i+VqLvsODIi2jtjMQmogUAoLZ6FY
Jr64/R20wVxrkY6Wet4pynI4XPOv8fbaPYy1NyH5ujGXc432xMz7QHZfTZSZln3h
yrZb94u7xrnNb1J9NqjWZyRd82sFBuLPVptbKXD931JIK2o6e6D5/bgYHBBHyMwT
VkDngwi0aK3vIEkVmlilqUYvgQwsPiOMms3+nj4u1Oy6bV8XCf1QlDo/DaAU26fq
U+dDLPAhUBu4K0meR74zajsFDR8s3++C4/xmgRg9V2lxHz8Ul7tRjAeZNd7gdTBa
mR98vw0LM3J/q7vO+rJhPnqmXmSgxZ3iuk/CJn9eDYhBXfGKkKcG1wM35bIIKQe/
aamPIMJ0DhADCI+qfyd1cPJAr+YkCLAN9XQKoWB9i/hnc8X6PJdePvJg7Q7NDju3
w46R0uSvHhpGW12Oq9ZIrmNS+Qac+fuwM76OOhVxkQcV6YuB4KAWXC5PIX0UHht5
2h5Zn/BIDmZYw9RBVZv4Thh7y7An48znCSqHSDe//yIlB/YpFVgwzvcVrL4RHJsO
puZkJm5gUrMQDAUkxxji326d9BG6KX3RkW0yLaNCgKyGFpdSBOc8gvp8JhukoECe
kc0tcn85WxGo3WZR9WB+rjZrt6JXC/mGiBnIMRq0VWrovzi6Z5vfUZQH1bDy+Vg+
dHkwGDPNR9/mCBDp5NeMuvbXV7xb4+xqaXHRYOjC9Sc7aPeohHm/DlH9mEbdVumk
8qDogQdF24jse2nDqbucQabJnEhsVJ64gtv4rOygYlPRBqurBH7KKt2kI3fsxLtX
+s1mUDeSEmt4f+v9s6+htIbsVpDHV+hTulTuodqE+Hfhg2A9JmqWLvN2boiaTtgn
kBIepsi47pJj7Ch7vDOghQUi2cYszClMOBdf1D5+hkfkwOJVQiXcjdqI3dVUcAcB
/QHKXXGjJMJ2aEaU8raDcZpdhBqkehO+rV6ghhhb8xbIVOpLdT4LKrEURlJgZBFU
04EJZ6Ee2mUVHklYDR0i8ZvcqVzIZN1dOxr33Vmzg0ppB805KK6REeFTo3Q3obcl
OEh21GwK5WrWvtNDaYn2PEWSBkQnYdcI3PDqszfEuBCv2RLIY4JW/fQaJL7q3OUV
Py5R2GzEDfqKt7MQOhcBii3D9dUIg+rKBJXfJPz24C8xXRtwovs3GSynsZkj5nJs
o3W4wifF16wuxpqz+n0RRN8RHVtwlzOajSbG7FLzfmeYu/4Ku9DUahzkvCBR+ZuE
1RNjSIPVQ5oBI706NhFXgHuebUN6VLF1d/HGN4u1vIpOTT8JWKUAOkqk60YEWTXa
Lo66zqGtMQQj66u/NYRGl05ZBusbEiIrOqhRt8UBSvCq1GeC45son84Oc0P43Tb9
Jyg8GhK3EQ+nO72VYjvuV7hoIjiImdehA2HYgOMudDiN7GcIQYPQ1d3ryBJ5Wi7v
Ubffmi7nSK5VTWncyBA5l0PLzNh3cLKMjifMQNy+TS7U7iWCSieUxvyFERyN5mmb
qowF1unWVTWnu/7uKZhTmNDl0Du7ufra0hqco1PMkMYtwifjSu3BrCuIUzkf+XQS
MhR0vsaZwjTpkJNym776H/HJ8ZzN3V/8Mni5MLkrBmn41hrssCUkU3YaZBfswATh
ukLSP5GFS6p10272H4weAtA2u5mlf3zfJgKS98wRaWiN/7PoHZVxW4WfCNrAGank
tHQ0zrXUgs36PSz0lbfAFlX5ULPGClTOLLBFjKFonZM8Oqd3rtPgGa1980XhAiKs
mMOVkIwzKwL45WcEPilI4Gst2Wwg6A3eJubcw2mhRjclQyABvBhv+OJgavOxGXuc
alqZ18Cj9o4CCvIoQEd8dMU16sf7sW+Z/hxcpciPDZPQ9KXvIufHpa0s/k9m5x2F
dk2a3NIQydQFBAfsA5Ais7FAnALm+sWSe2TifdOSuTdN26L0QoQL7XovTxkSXSPg
Uxp78YnAniKISzKf07wFbFl7W71xheb3St1Hqtu+QFtfujaGHEFBliECDLjnXwBV
yEMcf/zWpzUuJWu0CqNtUkEnDuFnjDSfM43uYn7d1DUiItD6VHgcog64OO9lBOUy
0KlYEFjiiH8VEwRmx3Cj6CJPbSLARkmESQcHCYPa+dqzz8rGLIIGhw1PvHBB60ao
YKvchhGfvUshJkPtu+uZDyeYNsWq0x2g6cY2yxW4EnFggrdi62CzEe4YuPAdzrxd
+8LTw4sGmup8E7+qyX7EWjL9o/n3oale+F+3jAFXNd1LeEaq3d2b/VLghytVOD6C
5sxJ6gmCV5Pk3kUwMJn59e5c3Es81byRolUCOP8U/mHE05m/aVrEgKxGP25gL8bq
BRNliXug9Qsdp4r4QnAg+PjwLH25T95Op6UIjmhd9xGdCBAdzJyuW/gMGJsBUI5Q
/nEl4ySdz97yPB1mBXVGnqNh5J1yD5PQuuOSvMXzCpMWC5gwq0P0DrC6UTc6OF6c
zAXseyKTNA2d/aqkOsqVBScnUHkRLwyB9lImwDzthUv8VDtFfHBJ0mn/MW9d5q48
o0lkmt8OpzyoADw0aCHjvsJR1+GpI0fDXNZV1G4Ntg5oWKfGkZuUHA21AbT84Pw5
ABYDlKFMpIgXP8RrMDzxSCMdZhBONetzyBalygJYT24a4vRGrn79O2+yOq0tiD6M
k1xCbjAbO7FwF8N3sALdibNe+nThYcswLubBfuS+ChvCZFAh7DLeDOmnnxAWR4qi
VnCiUuy9SxRUBt45jIhL0T0eh8LniLzITBJ4+2v0/jCTMXwMMees/gjaQKpqWFm/
sRp07BP0ig0UVweyIxjKG8+l5pQvkRU5midRALXf+SogqEMFSpvfPfrvM5DIBCBz
garWTp5dNQWyBMfoHJwzZx1WyQOrKNoFL6+OWd75pBqjvTBN8/NAtoQPBm6a2ne9
2sDI7hf4UkwpRKHXfgSnoi1MpQijca0XymjlGfSRMeGIMC5ehXO6QDhFWugr2NoP
yJYJIoQAYynylGzkRvw1FBJoQvWEoTO85xT2mMS9BqbfQkI+xEqYIXi0fOycqEw4
ybKIlcLLlPNPiZdzlH326smnVb0xf7XakZrID6Doy6C1qhaTtzeBIcEi0Bu69TDZ
ljWejovwtgywJWNf/WHPvkEjSGBc5sdot1wB5NHiFy0rToHpnW2rImkCv0k+wGcU
Gw3XxeHSfonsXtBel2YIYV1YS/WZ7doDFodOYkue8diIyTWBzXuXynpIqjgXKp/k
eh19Sy67/lU87MbtVc6VhZrGYziWtXZlShd67HFrova0kiWiDwdQoi7d+MHaKR/q
vmrf4Jt4CV96/wBU+gQzdjNaCf+1zKEhIdFJ622XM7KXdVNGCeyOmrT+18hCAUeW
d4J8hGgJMF0ODTSokzzYc3vnWtlkl2YRm/IBGXECxv82bCEjG2glL2NmwtveK5EZ
pcizwvz322ivFRZTEUet5gEhD50DdSKeeVw54vqROn8pRgnLAM0IpyUx1p/wVj3T
u1nr1FAZTBpK4T9ZhgTO0BFAOnn+15jxn5VBogAso55Ue+xN5x0FRkebdgnMqQa5
cXAXP/ewMjLvI74QvLYOpH3PGtk3LTMdmrpfziK0s/hdiL+gCx94FPNEtZnjIq/p
Dj8ri1vB+es0G+cWoNQbh3w+33hRpHwHWDgu/fwhXLnLb/cQUVPx+8NB2Lnu93I0
oe7ZT8BAzKOcuS96a5XZ5Ucfogo1smpui02N6VUoN5IEUCX/iXtsdk0ZJf1p9xqG
DUL0z2CEA0dYoGVskWdZj0mNYW4zb/t28pjckX3GMXS2gX9qfJjvjon+OpNaR1+i
J+4wWNHrZ5AK5VkYH8OMQMhCrZRZK9bK475PwE2ahK31tOYorLJp5/UKKaYDoJvY
UPRsSIxzvsWOl4TCGwOQMo6ERzCDdS0haVG8buMtuNYmVDgUsXuKI7JqC5lrkJ2r
6jm7sjNjNGmfikQV+c09v4swhLP8f5iWscd2GxOiBS+cNYUCD6kS+SCtT3A/xsg6
ksET9WYNSATebRn5SsypiLXcHSAGt3JS0CsYimIVm0iRgHv3zJRT8V4TV5LrGyb+
mS9f4ZFzVgjklZMDAH+GwK5TVU7QgSVwpRdUgUDDzrjPGDZJDEC767FmWjOLdmi/
670VdeOjGdYd/fL4zoFz1iCKOSaKsLUjqweX1FnV4bWWuPKrMh0HnREykLfe/nYJ
0MS9pHM90SIiJWBCb+IGUhI63tqnVbn5kfkdMzuEoDc7BQtukFOHjZn2eLccc5r/
Jp4rEqEj80DIT4O60mC4YbMCaB54UPLX7+TpG7J2pqjy6o9nMgwzEbbBsRg1LzPq
Qcx6YC1Pqi1qKJ7jcj0LajhRhKBoHS1GLLmUeTXbpWBvONReqN6mjHHX/jABAebw
KFLAZE5tDylW7XeMXUKmazH4DotbnrW3zIEIPM3urRZJC/bjIBHGBY1moxJnqlJc
/ViX9YQaAdywebBgepGe8PV4eykPcjy3Ih2vB3ZtCJpzwII7YF7Wr6MgrFkXj8wE
b7mAXaq6ilQuSm96D/fs7Nvf2Y2uEbT0pldEAR/P9jYifV4n9CsNQlo9b6uRDAjL
j6o+BDIcvepxhubd4zX/VB7vLD3i9uRjtag1OcmXpymNJEwtTw3/deDLpX6cpY9P
MKd4FMbVVc7rl9jTOAIIpoHOlLRmqqDSWjDqVkhRqDrZHg+FrZHt1jdZ3Vx9u2Zm
xIeNKhWf7hdO3DvHZcdlfQFixTNa5qExM3RRhSBf8le6JCUXCdye3GwCHAMZFJYy
BX+3EK3SEYxUMOPzANgQAMzKKqBIr+0n6DhezVg+PiTHEgu4WfG29Ba6mpxgDNcN
ECDrJhx9cLhHkhXAD3GrLCN7L05KrzzE+gxXabShGQ4BPmQuPnMW2DHI9TMOMUP0
yOyYhaxBUquImNHIstc6F7/h9h+A5Wdw5ZYONaIWsi/cksK/Vudof9WkLUqsw9oa
jD4D0/3+r1Bl0w2EIIqMIBYfv/o6irvVvluSu14HxgNo8lgr2SDQ6vs6whcEN60Y
0/dk03c54guhQEA1d0Epi9uAuewwM+dFoK+pzZ+A76sDimu9Va/vLtZxBTtmov23
oIuZPl1iphhcdwTWQ86gxSifWE1BpowF9/w7dCNsS0Rh6kR5VhppDEWKnTS/ctAH
ndMoBJ9M5B+DpGcPeQivNI7a1vvPcyQrpX6yPKvly/9YyQj5p1hQdZQDTu0MGbrO
7HERN9FbtGJldTIKK6es/V8gJxF0sbkJvIMQ8UnJ1jgSSpXj/WYSSO66l5AESLw0
YHgIlZA66rq3V92995RkMdogVfb1+WoOlc7CW6g4pNdS7JP+PpzamJW3K5RHWbpy
L2np5W0mcCMPVrIIk+KUZYI/Opg20IkZMx8x07R0hI5bO67v0/kuRySMKhpIuAup
zkjxRaSkcYqbWJH4P/GI/f3qapJZnMG1FokPaxRtP6poUMkq4GehQOwc5py7LEkE
B7VctmC/VI5JRE0VD021VuqqzIr5jxCkVOhiu3sNKUqZHRvUYlDCuHf1WxlYVyn9
SDbpJArAY+8kuAq0OFz62klUnZpEgsJK6yY/1Xd0ZFtv6dNsZJTpRACGLqrXGEBb
IVCQdApMjqJZtmxP4gm7IxpCKnD5z7MmgKr8RY/Y6Zw2jGw3aRR50WzCqXhDh6k7
WeK7htdKN/sT3xQMV3dCzM0zg9J51O6MwUTlMWB6rTsMmNTUu8Tg76Zt/kZz53sf
925ZfP5Fj9oDpgvPxA+Bqn5v5TAiC4BSsbVfdXXjhWNxJptNhAiy1R0M2HefjG/v
1hDMlGRW+1y5y4gd5AVYZZ/9chQiZR6K7yZSgWSUOSzSRRSvofXTbhVqila2MyWy
IW+mHSOTZwOxSXFi2/1wiV/3cQ6r0uDYI8DKTAY6r+S7BeS8yD3hwYQQDLDzNj40
GMVtyfeFERgpk85iTifs3Gfxf3OgtaAlC+g4F5AS6ENffBvTxi5BMwb6s3k5qqP8
Gg3GJRJqMDECA6NvqNdxY+ZKEtUQ4x1vhmJaf/o/xotpYxu79/eTSlxEQZW67I9X
g5k3Qd/yg2NR0p2jXPnFfAgdJKSSsmbQb5qLfwuAVl7kV+0uSsaMEJhKisvKc9rV
3thfV8/war7Vydu0VMlErGRCQXzAMOCjF23ppqsDziz+5ZH6lE5wFw+/evjp7Mhl
2bwCrFpmS5Wr+bAyTh+4zSnLiQEHvoH+Xj46P1OVMRIMD4mEiJU5KiLJUGhc0qH7
WtIqoDi1drdbtT6nukLOIGrTn6p1TzL6dPMxIToxJj36Qm4DzhJ/Hq+cMjGRg3Jo
t16XaQrZdWo0snHZuhdn1GLraPuA+nAbtxZpd9/ZBnvSBD+DYwVP3TtYY8t0K3V+
MiPAS78uGKstk2vWyLPrdjJ5Aw4knSJWXHyVLPzZDuCdnq+hh6jHc2Qj6apnYNPp
JbU8YRZvula6b59SOLGkAuHC9e5/JX9c+kwb6wV+yLRyQvFa4nNyPj4myOWFJMoW
z6tAOS+QMerbOJsrc7UtFeZZ4qSmCOQaLKCXHdNCJY2IBNjmn7Va25Gm52LJ6LJo
IgSuN1bT1mMEOCrGO11q5LtspRpKbX6QHIQmikbglgh2owG7VKQ6H0RTPeF/LCkZ
YzjKZvCMwgne5vbwTQWAjze7HWy6F3rjGHKp/VrqnXGbXmYPAqUcIztFm2ujCFmz
S2Z+xlmXYkiu4WruaSutA8AP58wHoHK8xGOUz/Ai5UbfKzmPYJ9m8/pPlly2ApJS
RbW+MrakLNYKaOxIXBdqJenCAiUa77+tzMEdlAlf/qJRQ0HPRD70AyC7rzXDo76m
JgbFJxcaqahPRSf82Qk2NLQ3ZT/sTSywkEafcKCK30ThH1yU218bhUDBxT+Rv3sa
Eo3d1B0tLJUb4MVZMjuWP+ppYOrsD3JVHImFmB8AiFSaPG3czydxXP5Rv8hl9+s7
6ZmZszWaOffTU22UH4egEqYrPtjjq+P0reCvCk0vcTfkT2bwv2aag+HgXDS6qfyz
uJ+S+OQHk1P7BpY0A3pleX4WiKDe8qJEo3P8MqHZfeMfZjP371ciu31dNpgbjNs2
qKI0LgybP8k+au6gC9CSi2uZjXxMgSi9qvBy3S5J9HhNiIqJ3IMKujmXXKzzNIzH
mAhUCwy3B8zIrrB/ADMxxibHOAy75vPAt70QZhta+9hy/fl0oRdTei530G+XfLZq
7Tn12vDwkljEFREj76t754cqDLXBXXOJ4d5yEA3X3q88FO8TgT/rvbdFc5XxOGsT
s6GrImcyj5kpNO74oZ+K4+3gpQkfLVR91RnndxOY4Es93Uz40ju69z2EsRtOMr79
LUeB1sqMTnTY+3ePagCz/LjDoVYdqoG0OO/l9MqFEkQR1DiQEJsJBfn77lyhXuu5
cEcdmYykeE8855p+BcCrJp1CbP3SuuMppt+RUTnno8mry9+Q2mRU2pPv6D4XtpE9
jHMCybX9Pz0vYNDfhZ3O+KcgKdd67gjmHo2be6bkTMRnKtcA5+w0Rx1poLWsWo3q
sqmxDdZObPCGW7L2MceR2RY1qFpCofcEZdzyhnIwtMM/DGC8y+C4WoW7VwSYRBeg
j3UJBQH7ZDsQxXomZhgfMwlI2MzzVMjHElMgO42QI1+rjfXM6LowZ+kezY1yKNbz
AbtFYhtRUEtN+lI70e02JKrSZu/S63iCroN6FyQvutC7x6Js5nws5tSUecq4kywV
TMz3j13UOPLNL5vLKEYqBywrR+585iWabHXWTvpidTXvg4OgizEX/N0c7mO28+fP
aciFAi6A2t3JZgu4fzYAU0ern+2Qw1GkVof2U0H36YDUIULrFnDufWfCGWabB/OE
2qf7Z80/0IeBty3jgA6A2oyr/4+0X3HZxhGHYQGTrpglPV77/uQSKJS/yAPvO6cz
mszPVwKo13Yh6Nxk8fLa5N2Y5hsp1ljszYtV+vIbxGL1Zq7aeAFNiaMG+PT/g+bF
t1ngu39c9dteCrhRlIJeFQbvSKXhOf0jro64OLJAuIvdajHJkavCmbqJq45gTaYl
GVLqGtD/LzWafOaUKwwJ1U3ENH3ZsVMI2z/AQBvOED7x55pwXwvLTd9EAoocmPPc
EmK6FmxgHkUj28uCPDKwr2w602ea5iwrWN6HxIY+YYQtJjpJL36c2umw+l6zDvYY
NU2xefSYF4y8t+MSL4mfc19lbpjH+FKVpN1tSHKJ11aWRssKul3h/tg1VjfoNrbj
xzm3Nee4WDAdx299xDwG219nwt/qr5qZSpe9MYxICju5RZo+CVupR0ZQ1XdrdZNf
HMR8lpu40sEuageFp5E2fgXI8B7bqpL+4GEEkb7mXQecrMTNj2zUaNx/3xZsoKzv
iGIzq6dRDk06qReoMsEO8ff5saSbyLu2MLOHGDniXP+qsdL/GkLoFNSWDNvQuuyI
otAm3Q67P/KiiDN1morK+yIm9s63lhM8UTG1Vxjnbx8jK0m8AjjbJoyMgmYaK+23
wfkhPyHVznrXG1pFegJvaH9IAaehSATcBKK8+c7Pe3xDkNAsefH+gDkxZsIgvONk
73gUaYG9phdAqgpns5/nibajyL2awjsFFWbiy2l02DW6s0hTB+4APzkJ7d8/LD/Y
ZdzsMfaFUEE5vLgtmPUFRkHxiHZfluyNDn1Y1uuhbmLVJQyNbrjqEEDXT88nMruO
1lHR5xtE2AGx1q3qdNSkpGCSihGPhmxIONIOf9blA/+hW0WMfOTMpo+ydi5wTkr7
PZj74zZOuxfF6WJE1P9b8NF7BhASIJTxcsPQH+xAp6pDwKohxZ3WMgmHQRDPVrib
Q+8wCjSce/AQWEE0agiZFRyTf8NpKBeKBv7Ze6lrnpywDumfsOtWPQaYwcuGqDga
u/EARVcCrUKcxyNDrju+/O0hJqYqHRKMhOMbQ/zS1hSBDyuSN+HqFLeDYgK1b4Ib
TouYTr6ShcebvrEdsu1d+loDoWL8m+6mlE9XKXCMGWQtXTqYjO36nEkId5wuF9Vs
sh44P8xLRXm/v9fBQMyjo8rLCo0JXAQMexfvhRF0/Xw1cEG7WVMJJMBjaNMUACaP
7CZnB8Gq2kqlcg9eeptz058wm0zb4TXO0tDmaDI0UT2gCDgzti9EkOHBYcIpl0p/
cX1uTBH3lTF4GFLgEDf4oP9+u/4MxpNI8iK/m48iepLOL2Pi2g/iPQr39YdqhMVd
3rEzBMoMPvVvp/bA9Sp8ikfceFnIXT7M409EezpyM3X6a9Rv2j07asuAuAdVbzpn
EH7Lsu+QI5KmLpS/nokotgKCiZA9dH2W9YbFVfid3P6XnVaHwvX5cJO8v7sCSK36
yhXuATRs6PWNnC4k+TAptJc5d2P+2SqN7IItvHDmO23qQel++a7St7RjbuJ9v2Ag
nd2I43vbEqvgWa2fKxTmiJjFqrd7sTZ/qRcSqKBNg6mYS0ENIP38Tuvt6EsFRrKt
N+9FQuS90e+P/W9ucUtwPlS0nBw7TNej3vNDnB7WC2KGEQIf1/pcy91Arghv4bvt
exRguBBHNspz/HSnDi2wKSTf30wLnICRTCQwH81IgOfVFO7Vsngq1qbgbKiGMOcX
3z7XJHtYHZ8BfH5tFogUEn9/1+dMcvRiW9xsE2Sjyyo5HoSAEYmD+cXKwXLMZrp7
mNVO0fHoYC4ZwLglv+R1ZKo+VeWMPTYCnmdNcEKgofCkcfB6YstHr4AhFd85hi6t
mGhyyGr/PBdso1zkFAlENIeaXPyttkSwW+BzrYKHOWXjA7yz+bHOgUMZT+WOEG7f
Xz6+sSwPGwbOaY2UX/v5zyTwZqwk6+JClJPSqUlRJ3hdbovbmEfoQqCc5JR47ycF
OhW78jtba1aRDSiXxL5wlbUj8qmqlphy0+Vi5uJHOHQCjrtyf525V0rADSWLveIt
LbGo1ZVQL3xq6ZKwvlohyeRIl/3cLePKeQSqNoU9uif2ZJeHUwBwKNHqCbSkrb5E
nuQp1Bijb+OCeeBN0os1Y2PWaFpERa82e9TqiMiyrXQSBDrB8g0cGX/KSBwFVNaU
cIL4KBa5/nvcE6GheO04QutCGe4+e63HGUKcGPXFOtbFCdZgMpYK36qwspXHG4ve
DKBH7l3tILwz/j1uPmE6arKnK7xT3u/NNXfUkj7yZlnVOVLwhG+xZSatRO33CLiZ
yChJmwsxQL0l14ZKRhBKC7xQXEVBRTqjjSTz4gqATudTjBJWS6oQo0co+1TF29mW
SInP6iLaKtWbujRwj1Cas78aLPEb71UMoFk5d6cEQ0vsxTLTyGx+/rSnuFmFCzw6
z+hCIkSApp/aoAEgnepgA6vZ8BJuqKw6DZfh6T+af5j0zKBMVOKOc1gwmIzeiabG
zsZo+VRlOwaLihoMtbOnujbSU2PFb2T+/6o14uTP8wm0x9ZetDwCRMF3nsKCd50f
rF4L0Ve5b19tDfvp7CeszqxVql03hdbhWnZb4WloHDTZor1ctJ2Fr3v0CPdxW3su
RKHjXCvopDXjFgaCEfeN6FSNah11xI3kKn5M34zLWnUPrSVbtBsJRYWH7ehydhup
6Tt+8+/stsHxaQy6FFQqm2xk9JGoo/bOMNEnq7xyMmfIOKZ/l9yKc57VDINFcnsr
vzR3+4EglwHZ8kAPXZC351ZlPcxf9a9fxKCFyfIGZ2EwFDTNKjNCuhov38XDU2hv
Kf9G5U8xiHMhEowA5Wk8z/ArH6Vxecuqkva9/mfxb/CGCsdZ7foOMW59IjnDbuyJ
OfSELsZTHb+KTtrr8w4teYGC7fUrGZgnVAf56Lo9chZ3A+PTNW851nvr+Yd1y+gu
B4EPSP3ntf8lNKg5v4plmJAj2WuzAbGP4wrHPrDUWj3oLhOU+BL9BZdWCJpPu8wm
gE1qT+EE50ua7LLe8gq1vc5FJRp6mCg1MwVAraZjBOslXcU9yGPxwPNhuqgIUV+T
atAkEJ/dwKBksve5jzLgHXfQt+YZ1iSlNGXPF6EEIBQQ9sqRiKf1zXy0TIU5u0eT
2yUX9rVa/aWH6qNpY8rxYbc1CDgLDM3MSwnh7TupURRLqUJ+WopU1oqdwsXhykR3
xTekiZhBFy8/+IV/RRTYPoBIvrpuU5VHAsgtjtx1OK/xykTT8uq2a/fNR6Zi1RNm
wCjChPk0guyineN/D0Ospf7u+QMqo9X6pCA0VQ5QVMDvNzYFvE7gLinHOENHyYap
eWblSnfX8j4Ux8O62AV5R6lZNEMFHb+bTaPn8smQVZ577zRAPt46zLLS5cxVJS6H
yCxHXOnsQK59RMk8+aMYhLJgCXNPLclGUVeuxIvKZwrwFWKxd92MmJjTIHju5QsW
CwF6REq93RBdz09VI+Ausc30+Eg7b7dd9sjyp6SW6CXGSQ+GWUj09grH0nngqXDn
mnioaGJ4v1SoVmv9PuAhAtOrgvU8Nqm0dC+FSXeCvdjaR/+4hkVzhRZo2VE/uqCt
z0Fjlime+CtF9z2utHSGR2tAR+8NgCYaz0DV6kXf1jsYQL3glyFPmz1wNeyLNQ6Q
Oc2Utu5KFVPmrukEzIy/CpAwMNGmcOcqJyCYKd7EjBZTGVGB/z+EuPjaRRwCWqTv
mXASmGesJJCJLDZj878C+/DO3SqKFohUK4ut49EQQkLqHTKQffCZg62IFzWHQc/j
vXkE7rqp2wQwJNtf2Upb2rh1ieIySVEt7en/KcxLEKA3D+SEteG7krVbeRPX9rBa
7GwDTDPX1ybFJkqTxnxg+OgKVVhJ/FgP8NGGtMZUIyD83/HuHNyy+cWlL4xkv2P+
WQ/g5tI1Y9k+I+wBAe74lf6UEPQK/6cun18zSkJuzqojvdrQaWmYIALgFG0T6Fqs
vLCzz56CohZgIs+ar7+ecDVnv2km7T7/jgv7v9DOACp/5rLL9vIg+Z9/uFpL3oVu
D9zm4/d4HNgFog8Hg1m8RXs5cZaEzq07KUcBxSEfiYxmFXdKzggc4penS4RJRZ/0
4ExdDVMmTvNtdUHptZspaiogpKbpJik2YbThHVK4S/YUv82IxV4VJ7xravtofBCB
DHqfyH5yUy59FUVXjg/HEnrCXylUxA3NC8X5A00wQQCinC51GhAcq10Hm/yOcNHH
g6mZzHH2iMfqAhluVxqfFWun91dDb7elVY1wKS2wpck0KK/BGJkZVhXPO1HD84fu
NpKrHQryNdiK+Wp3pDaSaT8viLB093wS+t27o8h9Y6fKUEW+aU2jZMfE2/HsKH7L
js8opydldzH2XtNAFTFACYgSfdaGnD//H77reWZrXG/Q9XvewNI8/XhM0x3E5G3q
psMrH5aQgV998vS8l5GGnvbHF/rW7TMSD7kwwHxaWRZG8Y0tJ00a0ddVKBPNkkpX
STyMsDh1p3lJT4Z2qOiCbrdhQhSlDtClminNq9kx3FMmiS3o9vNV6ifmWBDNffAB
uDyqlysC9mTGlREKg3RX5Fqe/aq2SeKHnKy9bFlcjoYMXC9RJzNpx6nQcAR/lKxE
niMAh+y9rabPy6KAEkP9M/cDDqeF/ctm7i7G7XiqvDrX0h4+BQ680g5/SdS1+AsL
H23FMVUcL8szAaoxBXB88Fvk50u6EbzIoL+s24AJ93cNf2d0jVRpRiDnqc1O/soP
8iPCXKPOFvR3+kqvkKGZWe03iRIu8Y+gYBa4cWgLwA/ey4eRoFhLsmo0JBNLOo21
A3YA+MPojL33nIJoN5OYYJS5scS+OxO/f79/qhn/ocxehjMBEnPt8/OO9317+gcF
GyjRIzzShrBmTPC8BWXvglsDP0yINTkzd8oUABF829juIH4fQ3mMaj3wQRaLrn5K
sR1w71Uwoo+bVCdw2rn7FGQPvvqaMU3vkoTzcQTXbIp3jXa28lGmyRHIXNcLHnAM
OieVwo2egbHeVJh7+AP+3u9OqMjH00OCgBxiZeEBbb2oZjUAVdLLRoKKcj7L4+bX
J08WdGcjMP08lnbyEUfF8GPHO2HBFAKJq4T9UQYwW9Z+ES4g7KpRKrRpnPFlXQIa
e1duAMFdmW0No7AARhlytBT5Yjvur5NCNRxgn2kVyzmDj6j2mMUPECCq3Klhb2WV
zi07XPvyOwi1ceZUdmI/AAzZSCe53LtlyJ7hDWKIDrZRqw+d+gUUJ0vY1qCBGorS
cOyYf3dFtP3B161xeqXnSqASQTpSpviwyMimdkKHpaft6O7/F5dj5aIG6K8Qjc7D
AmPGlp+IOrEDULbijSxuW1hqSDx9HWsqH6gZAYVCSJrL7Lebpata0Yo9qc0UCP7d
E0pD5a7GA7a/3pyVqSXJ3v0VqBWbKrNfay/T+9a9ceW8WB/Rcx93DLLi55XZPtzl
3eK575en3xVh2nkzKdloxadie1Zb34h2IZvxYNAEBSIMI100NlnIfy2EkXYwj79u
AQRvO6URX1cKH92mz1pPqrvPr0NjR6HndTzs5u7lvsTfkAR+7WQ3HbWuL5gf2meZ
IYdGFxbJ5xb3vHBb9prvo8Vyza26prjRj/GopvkVwIKDjsTqiARslpu9JtUUAPXZ
uUYnZ2dMSZ/bwRYzVGhGE93IlFQEvQT6CbutyMul/S8Cpy6U38tQ0Oixb2h+72HO
AUI+cGaJB7mv+16/k0Ol2k4z4r3oBZo49W0lrED3kcGQcjANEyt6WaznMjg6de8q
MeO/I9l7pD9Zjj0fSs/HpgNPybzVVd6rkq9jSrxnnBlpHD8whGSz64ecPtPmy8CX
5I7kl+JHgVa1R+ayDf2XzmrS3jz4Qfj66pVRLYmEvm1vaSDQ0rTJWc4BCxcZ+M1u
2TeLrzfnJmDMXmm4VMEjTVrI9e/SqrvuuP6UcMVeLXA4+nqYW7RfGyA6mLRhlBXj
1tnUYwWae5vSlHUuRkHIl4Wk37iQ6zNafFPgWtWlALAZXtQiFyMU+vqnE3K2B6pB
+5cJsswSvmoswZITe1w1lrZV/1mLCbiGZq2HUY3oBhC0t0IWZGbA85iUmsz1qGBn
uMSH6VGq+gBN2MzPdxnYJbVUzQo2eRwy+GfB0jWctyaOi5nThbKaW2lHwNK5hvj4
52b5lGfYKLk/vzdwPsr9KlAiq9SlFwnbuP++6y7MOS43JcqR80TUSBjz0Fj1+9fw
YT/Zxm842cimsZsXExTFA8tDoSLSODY1AxLatk1jwy2cyGlIrVWTrpalOrVie2yv
2/AgN1AQr5htXlgNtUgY3/ztCGTDb3igZWaDAh1HlIxO7a9f5z/WdoLkQdgtpggt
8QnwqXuOVSrCoWvja4ZenpQ/DyV6jJ+swG3UqiZuhTH5svxndnnbW/CW+Al8XCgS
wH8Jb5vVkhJ6CE9XEbUA2ns7/v+8zwibpY4A5AYN+uSBWzHceCWqYl+Qxdo11MJm
RLHYR/lGu5H13xQjwL3/OKwfMdcuoz6VM/PF+gdImac3C6UhVHR5fGiwj86Q1emZ
nR+pIZw5SLC1+8MhPLaNT8xLgb2Xo/CNt/M4hZbKssrgEWN177T1TLJZqVGflAMa
JsTXyNhbBPIHE8sBs4OdNiuN6CgqKDR72F7ju4xy3CTN8QhUXly/4owLP5b2+E/N
H3JKA46MUhKsYmLyfgSXF808YOk92UJeYYt0tVWr+8OcHZpiEe8yyrQIHSsSnw69
EviMXdWINpSVjymmHa8nUVp9Bweryp1OkJS+yOHBYaNHg2YL0IbICIU4EI2fzLer
VfFhdjGD9DV02bw+RpVSs1SxkrfIp39JxhGjyVjQ2nyw5y9nP1tmWhfOf/q09NGl
nNRkQH0dgsej4drF4M2MXv+vc92JAVbgMMlF773YuM4ccDoQ8wvAApxc/JePJxo/
vvte0vzBV9VQsTZkX3uweS0CIWsbuRkttF/Qpj6depXl95jQS7zq1ucapt5tt9nK
YDwfgI0WDyxQTslTSr9k+ATLNC/KbBAK/ANPWgWWj7omuRxlrXwppgOvzDaCbG4Z
HrP2Uqr5fqPSL9jvGpRGAbKSz1qI9PsykqS0gJcVjrkH7Kio5G9U4My2fVCLkbgb
C8rJmDQFQR1EYWJsPUXnx42kdlSxpH9WUWnppvRqGgCyijGTScyPaR9AsBHBhs1y
+AU5/XwuTYvl+8r4yBa9ZwRvXrPZpHqv6Qj2OHGBALGK0GruHHX52jtZh6ZOYsbk
iIJ9f29OLUPeKnUfh7RBIJ3wU1v0YFFzznLasA8gJ6pgLu40NVC2yEGbmXw6SuTr
5t+SDITUvK+3OONZoHr3ANxNwtKLsDKR8rrqX27J5aPVT4XNS6Nl0ojBnYyftCyN
p3pB06MkAnFHsNnWsOuUW9tF4pwZQ97x+2t7UOp78ZRGFLGXOkOD7Kea3kpJ/sY/
qRrBGFlC5TfrfRjbWJGLZOiR4yLCLanIi2lUnfft2PA5MpnibJ/cmxaNUjcXyhce
oKErK608J4LKknaSMS5T89Zox2cgUD6XlIUdIpjLyDhSeCONUgIjeCfVHT7Krqkc
plc+E4eQLAWCFwhXDWo8K2wb5kOeGZpq/UnFYZortGZTMrSPx288F8Hwym/ukhKv
SFvfV77sDjuwmti6Z3MOY4x75wwPIi8g6Gzyj2G8CbgHIOSZvXSCskhwerjxqhCb
nBId07ZaSiaDXBUeh1QdMH078lEsKGO42htkTzn1bkiE8NGiwahQNSrWbYEVNFLd
De/bpupc3OIATCzPk0rlJ3V3K8/tYA32YjPlNXYHRYf2GWOOXUdZmU4P4nA/3fTq
K9VxF1wN2X1Ga5+mWMX89Ug4//lVGc1vQ86jK3b9siSKDQwCwtvzdGhATAgTmtvj
3JiKpeG6qWX0GjqQxZ0B1OrGkWK+BgbH+kgyAsCa/N8mQR4Me26/TZVQxxDw95++
3xaDoA7etP6txVsb5QPzRRZi1x0juIfcpzim1hukCuI8ZUEI/LwJ2UjnS9hpUyVF
MqH/MnpINISQLvfXyaGMCbxPPWIjm+rA1Tpe/h8CeNUeCAB33h5MI+uvZwUBWAaJ
ICpbyYTh9/CcIp+tezigxc4N67p6QEhOgGBtYUrgqwMOOLnvJkEAZ46BvwT856qc
IjvjOafaEkz1aPffA2py2CqJ8AuI9vfRJFPWD8DQKWJCGzPNt0fQfmiCyl2FqKWN
d5jiK8ccBs8AQf9hhy76VIsyiZM87pI5j+uOT+n00gxUG9FDjl9EbbUjcSr5xIh9
Szg85kpPaG6tveY2RALwDRLCDIYYsbNtmRkk7LiDHVuLaO0yPQdZq/UZGbuRZyFU
GQT6L9WJf/Ns/VKwl2iewUGPQl/DlKrxQruKiRd0qmHLt5ut6XpFPSx8Zeqlx41w
tasAV3csQvUglxzXZj8VFsOH3e7+wGQYXDcyo7HPI2mDuLMMTcSSabDoybsBjSof
V5t+LAAzjTKilCMD8Q5AuMlwXeamUWSJWqcorWhG/ODblfFk/mhwMvPiEugt39fo
P0BpMnpFOakLFZh5rtmrAxhiN+NRj0hFQReaRhgHwkMtERkCEHstEjQRAClwmIGL
1wwD6jVpAUNl4zDPEQWyPt5kNtCodaLH/aXnXwZNgqNNaWyolJ0bLpTe6zOWZHyH
Vp9OBGt4So3I8NkXl9yFEZAvnDamZw3r9Dpa17NqZ+b51VzgD5gIhdtq6ACF6aKV
4dZlQIkeVuCRSFupwQiolqLad2pn8AFOR58+ZgAsdzs6qqUJ0Y5HriH6wA45TRhY
B7UoXKEXTmP8E5nVGBUlowU+vtHdQdXmXvrmtW2r1eIKx6uryjymk0X7lMnnab4d
EgxmEUDbEqI7Y+OJ3xVf0VX0Ed8LvuzJqnpuasZKJL15+GpzA2dQpLnMbjC606O2
oVZPzWpgk0ZNoCYaLLAfPYQTwjKmoIovm26GBuogwzq+k5ku85gGM6Q0TJUhA1oW
k8tYWnr6nBtp6aE5wNi963SfvaVZg2+9sMARRXUrK8fRUiDNsgC/VwvISuVueC+7
8UYh2WI3ZVUviNg3S+8t+dCbloFhVMfVENk1jSxNxRg7L1RUZmn6JK6OdSvrPI8j
/yAiQCE8kNUhOGytVLYxoxSWjt+o9GlxhSqPJthMPGL6aiNhkg6jUk8uEWsPYDBx
xNm3l+LNXSl85IPgWwMlmfjHizCZiTYSBD/rqWnP9+EVNUpNLcwZYcRAWvT7XQ5D
8nZPiQnm3RNkwtsWpr7VFm3OKtTJOyZ24ZlsPHY0pfbJibqNH88JhC9Vyd4m98Wj
M+UB7jE5q0VSC6wh1JKLkto7bGeDE23CIbBfzv7NVeyDDGRs6ZevwPMlSju2/0rF
8jjdb3F6E/oT1xWeHSQJj62tjJyFQ/OTOuwOfvjEVHwtk/Gwne46PenTR/Mtn/B9
mKv2Exr2/YhjPSgEd0bVg+j9d33PhyDMRb3az3+RVZlMoZxyiuXjYGAYPq59P2hy
679YHzCL9n7EFS1MDjvk4LEWzfuHO8d++P5M7FANeSL4GaznWOgEMg7WUHIdU4Rl
UiUo6vMPZT5upcDF5P/3zG9Du21jA8rOKsxG8FXpYKrtcJyZZKcQ9o4z9o7qRwJs
uinUopYyXOfhhNEyl3+3B+PpPP/mt2QGqYVOgFkqhsYxUrToFDT3eAoJTaFaCyxw
vjB0B9jE2IGgvpfTIR15hHCcXUy9pSf+5cb87ccUKJqN7N8rxt2Z3g3ZKb//yCYB
o781ZkG/cFWygOTF89ib/V3FIPzTDUdRXfwIT0pzfh9AfJHYhVzbqxJAg+V8NXCR
41INEUVLvpsX6Pl3S8H6/ETXhHdpqgxGXVolrJzVHbN/M9kvKMOGTDmozu0IVK3u
UL4ekH4JTGwOyOtWPg2Vdkw9Dn5DNARs5cP8jNwhhydwG+TsMl+Z7VlOoGVtttn6
Ha5UmnAQsKjFUzjN/l3ZodEZJNwiQOX7cn/HoubCcTpidVWxvFE4wOJGpNgVzjk4
p/KAjnzaBwuijefoRx0IcSgtgwNF3pw2n0sLtEgO2Mn52V/y/DDnsUUTI4QzTIoa
36yCj4TsNb+DxlcGur0g3IDZR8gbhu+MWOhlYAtiUGwfBlDSwjd7G8OBcbMJq268
UL/Sgc+P61FsnP39OQVELAnOu1GIwjsufWOjSdNb1DEBky8PKyxsC7LspostqZ7c
OBXvIDRMhOXl9q7Bn9L6ZPHcfj6dfGMmnbpp1aYhgXRFeKCIdXNGpcOWpwTFyyrw
XyVeGuoh2Uvkuq8j+dQhCKUpN7SxbX64DghibFoj8WAWhhdmqw0J/aqK0gVud/EX
y/g2kojwJljBZtZX4Zeqjqel2eX4OLgERr7ulapQ/i6bhBlAA+j5iPwih+AMKxPJ
Fq540dGS5F8b7XJIRusxaxSxxiGGAyADviEQzo5yBgfk7I715oHZ6pgPPD8V+kmZ
1oAZKSudHYQ2cv7RIps9kXC3eSZf/dkpBYgm7WAuiw2as4kHAx6gl2Jrpva7xpE1
qrnCE+zPMZ8fEj2n9KkaQL9w7ycfREpfOki4EUsK4XMhwbe3NklvURvSDMlaLAI8
WVhQ6K9H50CgcJrhzayZuIRuhrfZ2j9nbAQ6M3qua1bBZ1FEQeyCdXNLmxa4lgt8
QLFgoSpudiFc64hfHy/bRMJIquB/qcGdTOxNNPUxk8wdmv1Cg8DQfaDbZj+DqKMh
81uOfaJ9PWyXlIaXZVgZ+LuIJpMHj3J6sa8QrPUB3kvbJmNuNHjccoboJZ7vS4A8
y/Rq8dIDOONlGVnfpsVMovnLo8rU+jIutRJeEmmxE0Lh0K8OQrnlmv0aKIn7Y1fG
p2O/5Fq1jabg0l5bEQnw1K0rdTVQOyHhnGt2H3eS+q50v+1c9e/LHIY7cpGP1XxC
E8LPicUtb6ZJZ6RTn2Oc9QdSHwOGECVOGHBOgIERZU/d+e7UyfakLCHgqj8lqPju
RskY5qDG9TznujZoIDQp7FZj+m4iWuqkIelhXNZHKO7AuOCB3Wg/tcjk26WlJocO
+UukNheIRI6rb5208AfnGbZjKsdwjtfgAkS6HC/8cLxXl9SqOV+yIa4f9r6la8Mo
va4SrYRM9mxWpsiW8c6+5xYWB1QZRoW7qZXlmuvZzqEtAC9ljRvRSwGEbv3+7mlA
b2vdIGplTucIUxdy5tYBaMm/Ctv3rSQVRD7Iu9Tv1VevI56EdmSNQffMdCCqIAHy
QSXJ85Kqn34PvdLhxsojmC4nv+Dhz2pYoF7Dt4dF0Y7z/mkFT/ArHWTljIFl+bYN
Ru83qf2hr6v2P2+QeLoae/CXAvGDT0FLGa219K+THtu8dsTHFlPf7qjVvPvQZMUQ
55LqiDJmpW9dKAuXwdUh2wMIgJseQftm07HNTXXRHM2qalEyq/AP2FSDSspyoEG3
7zdKwmG/v4kce22w4dfaRL7tO1lS1BShrqFskvsAw96MDNNlCTJBoZ4sabjaoJH1
NEMoEKGvOEnDeRMNtYAFQVPLQFdOWBc9M0Rm5Xnzfdxl++Ws6QzQeYsnmC3wNc3U
KIUP1Zxz7Qf83Tf3sw7GZsY1lWsSBojWaJXwat+C3EALwCnxiPNfBtaQ731Ohj1u
CntizRH9xgtrJjiaDv0N6Cy22pSXzpCOO9bUtUvoiftJZo0hHZjB6xM7XEFML3Sh
O07o+dFbDcBooEGLW1aFK+eKP+M7+/RPrFcdWtZ98q0Gvp0FfE9GjsUSN04XUK+V
2PIetIHUArmMC+qUIO42O61qLO+jdoPuivaQoMqyQ+ogHghptrJwRslEKlN19MzD
Wd8JMJEyodAkERG81smPpTzK+VrbB1oOuUWKJ4GsID33tlWN9ZUfcMy8/ni2SmWV
JxfK+ghzqAViP5UR92lQpleOBdmqpHVgq3dQCpEZnOPJ6ZH5MvIeDW3j7lzmhhGi
tVwt3TKIxItjbxeJTXdgT/dTg0Ay3vivmkFGC4WLIcxWuAtbF6czJvzrq03U9UwJ
VMUc5BR8EfJy8H10i4cQG+6V8VVYA1TYFY2HPGqgF0v6bxIWebL9vtT7yr+a8CFx
1hRkuNstUeFwg/YvZwUURZL0WulmPP83bgr94wW4RHUWMQp1Z9rXXd1rU6Ua9FND
ZskAiqAq9xbIpv5hrJiPAOkPbm2NIzTSfQXzBZ64AJ9c+ATwTbqHhy00ZVvFBsyY
jUCU00QkhY9P29bDx7U0nEYw4Ri7/mrj1/VjEO9SLHeAb5FlDuCELfLD1AuOnAkl
Hi6eTAfED7i+4TvtzgZHLmCPkIbzWe4Ta6kvWbE5wkz6yqauRQW/hPKlcr5Bfmf9
qc0WcH7RNfkIIR1sYXdZq2zvdhwwrvjcHvs+YoHdrj7ZM7DmxjfFvwD42DabP7NS
6xZT0d0qYbUwKxjLy0O113Rkwi2qUQJRUmp5CVvEKPSPhpb5c/wbFl/FtrQRhqRZ
FEzmT49gYwZ3IpSwXKsBCYEW0zDG9X7BNk5/SzUCCbGIAFU30ryr6G/fIgMoX2RY
+6iz1GrA2C6NcJuGpjnE2/VjrQd9icv6fqBW6Zr+QkdMTVXxuwict5mVdaIqi344
DW3irpVe7mQQ49iBzAf5giVjwLM2n0DE5wd0yZ8vW9WKC3jKE412tG12G+H8uWO9
Zh+H/ba2IMjmqW3KVJmqhOP8pkQ4f3d2OLcaZVtiMG8bMEXV8X2GHWxEkFcv23Mt
qmVrPPgivRkX5Rb73JB2g0VcUhWKVtJlm96WAwIGa9+r/CpWyr8dgJuGaHmxDXh1
M13Qe29nfQQ816wJHwm5341kQu6OCnjbARtk/11D4yGz5lNWDX0B9NEz8cF6GfAO
sBkfIyeK+WdISZmXyZU706LGb4bFQVxd+9k7pOh6/A3zRtwXh0slAv2TWAZjwJaE
yM3+6MQuYhse/YcYHJOy/J/8lHK6UgDxzTvuTS8ltdHGF6EmNBlPh6PAi70Vccq1
tRATaH6ivUFOE7BL+5xGQUquUFYmgeUkoBMedNANE0BoZHNXO73epfvEJhJsMnOl
DSv0/4KK96lP8F7Y/iurPao6N6BVJmSf+biK+G4HuO0F5U7RdFSKKhjYaL4QEngZ
uWjXcXJNiWWLcLwX6Ah1n+1mcFjNkk0H3etUYK7IRWKkKVonqjTLmWddD8r1l74Q
FYWV37irRC1uTOT7XKVFw6nSvJEbHXR/I5DbGEQVYBXwBmT8F5C+r1UxXis3nfGf
fyV8jFaTkxXxas0Z2SqVOSFEy1RTjqKMbpmspd+lN7qRgosEixotTXVF8HaCwoi6
n7/GPBBUj8rq95DxRbndeBbmZVTAfpkqXYhBF00teE5OuSqL7eDV8kewR0a4CIz7
2qIwl6J5CVhYdcUo9Iguys8YzWI45GdNMuiyY5GoCsgV29/L1K0F+a93S4ELQHtK
gNxQaY2ZkNvJHEPyHeqbXB7h7suL+g8yeuJCDmarWG4A04cUSN7+enTUAEXdpCmd
CcXxd9UQOuJN1ISA26yQFe2kPVbE+NnqaYrM2JN9zDb3XPJMRudtowc3+ZImvw1X
WqvoMWuQvJlspgr4XLH9vcpOPZtMY1nNgzXCWveTptDJocctUZQ8cSjoU35hADN/
LpSAm+RSPMD2dshrcdOqF1syEwrwUmsvziYX7L4lG50ZwICHk9yvnCuHsEyskOAa
Hrf5rQcO797k+nO/ky0bcBoPzZOiK2aCDviyM7aWDmHQIOtdlFu1oom7U8uy6Jh5
0iZKd5evxEPi6/VpQgWQ/NsKgBP+7eMsZk5Dgwt6zI2Ozgvyy0nq1hj9zw4tnXU3
zRkAklHENr9Uy3l1Maw2p7BZjpMAsmMkc0dctvuDSnoBkd7tWinBZO5yyaBvioiZ
kxXGoDwhtvTGwf0PzHU7L5OizFwIjwXYMu5QpUJUpbGftRg+qLmfTE1VamN43OS0
eL9PDH1ETLonSaYOaN6z6xc2ULKWLUqjDHACRlJJpwaVCAnxBdlPz4Kyu60K3qza
fXr7DQgZU5s3obNt8nnOFCsk82jAL7EuVVEKs3RV+991wY6uZqYEdjKkZPqwYV3l
qigCK2PIzgVuodRKx1+a5Rp0zAnAK0X+PUv0g2iIT0+Hza3pKD09sT9q+vGQS8iF
eNRVl+UNUQk1Hc4cExiy+9qKVCQhSH2ObNZR4uPWWJMbJm4MiWkkfYt8XMxgwCW4
HLIWh/Z3dn5NPVXJdgYHIm+CunuD4p/g5HjZi7g/6dIO388gkQ4vJATPMf5OVUXd
W/J/UdTBGmtS1y+4ixc3zP9VqY5Nm3DEd1qxyPLIipKPmDX53WIyM2CCMArLcHUF
lgCwCjEinypD4GdyPKv5xX0KH5prtyQWx6nWk2ZAtyC6vdyEwinL2k9HC0wlVTVC
UdTXNdIBUFWZZkAUYkilHeEGF++h7nvs8RhpdAQfbgP873YFNgbSxRtxdQuEXlYw
FnMXeyuI40qvU+MoA8EoJgK/ez8jyfi6B77P+lNLPHhRJy3nbkKKecHHgPJP215I
XIZO+LNDzdrbW5OlXQhMSLp0zYS+0LowJkZUidjm5M7TEmneUSPb/hqVlsFT0Usa
BrWfB7M9iJu+8RouacSlunbW/1X5VaOEp1HlLVwrfskvey2kpoIbYPbiFVP8M2vl
+9VuAig8d9s2FgVew93hIBH+q12EM1us3qDyMu8fHbAnBwdJS2A+hZ7SyO/g+xnb
OgOq1quXRC8OjGmr702MvBToDAd4qe+STCiPAvKG68JYxOuY9bEXMFT4gJHLDpis
riF08n0XFCbhC2hZlHRnI+AKGNdMbTFthC/0Qd51yhYjJqIHqi5KgVhiwtSvXU8t
KTxXp7f2h+glHytmj2fiLgPU0KfN21LMlxcLkiWx6XJiF2rdq4G3F9jSz8oUIlpf
niVxaJtggTzYxoq79sn07x9HFHZS3VnigGu8mTg26kr9azR+R8K/milXgYVKacd5
NmJ2NmF6NYx7TwBwBqeA5LxKWZ4dc4q/vx6jSIPWbL6CSjquGmvo3Ii1bITdF5nc
owE+jWZ2oW3wTJkmj5L39j8CI50yNVy+/5ZFs7dRbZ0hIcXcEfznMoPlmov0R8jH
NTcAzyTwKcpmL1YM4Af058+f0iaCmwsedzD7Zhh4CRepQIl80kl8wI6y7RNlen3a
ttOaiGdCNgjYcbA23+zaPolvrzqBNNMWZ6xDpromqlmkqfu13qdFbTLhMfbNerPQ
4wXRdVXH4pyFjMJ7lukpeCSyUge1QwA/E2Wy4LU1Ty74IktFEV19bRW169oWFsCb
knhwluYaxftsEcqKrqYvWQAQMwdneuyFUZQH1YGdKrLthODpa5p9S+Iu000sA4/s
d81L8vCA3EFfN9OBb6iKAcJifSp3FbBEgStaSYicniwhFj5XJKm4ZUv38kZ//XPv
xtJ94kOILrFHYakJfyRy2+y/PdczQ6e1rSoWxj681l3795o7rnvtRwBOkdBqCPIv
TuOqqV7c4svyrX9SkFnavYC1MqyGeeLJOYYUvRfWYhTotTHARMN4kQNbhSdoVcSs
s2AQtgaxlOQAd8VbWBqHuXB7dBgkb9O5oi5k9AVYaamvQKWpsc2n/q4jFYY5twmd
cmT6tRwYEq+n0gvS6Ycii6yqUaYDT9JHogTNZNYTsWaudMQ9CaQW2rNAh5Z6nwZA
oB8UrU4jAw/t5/n+WqdNdv/9Yj1aBu+9PDC1T8Q9me0FYTCvP27hQCN0DmRv4pF/
gvxAeGCI6/j5kFmqnNdled9ZwHA7lMuelo+QzJxhYg9zjnWDKJUk5sfG54Dh2ZvS
zec+/fhydAPy6Kj/AG8+zI1Oei7+Twlu7tylJ+BJS4su7/ge3JSOt2TK69Bqe/wk
D4BYfnUevb4A+BPOWyDliDRmGnMqAFkNRloQTfEH9ihq8uL7Ymo9QB70KC8NaDI6
UzV3gNjeIqr2WnHzQN2Bu/3UlgE3bFlvo0jyLLmq4HEKeRdSr1OazV6ifZuNOlsd
HcNtbDUA4hToOjU2UpRQesHSQu57lorjKA5bZ22VjWgHfzWPCUdmm0dzu4CBmfFo
YyR1e3b1vVnJLgfgLjYz9WjNjPVR1hM+0afydKvtNOLeqhiqP2NAtIPBl3d2VEYI
NIZLYjLmrqcKy8TVgz6+CyQa+QkinDX3T8edJe2XosT6FD6U17Ohthw3/jF+vpu3
jjuE09lrwCVLFZgcWKb2bRiPdmKjTLQR/PLaARirdmrlmDuAzmz82xJxbFk4Wl5Q
Z/plhKlfOEPD/M77O/1DgYJOK1FhihvGJC7RtRyuLWVZ0MVd6o3mrzhriO5Fsi1i
0+BFbUeoCi48Nm0ag7PNBpL5gOGHOfSTyFQATBxaNtPwZWWaR5FHGloKtKV+G+Ka
Sv3DA2vdkDHqAvBXUc5Izv+uwArLjo9tgHV6XbyRcOfCEiNYdP5B0VLJxV1dmKnr
8MSIYcabaquiurh+vMtQyP8EmMphs72qz11L5FoJZMY6L1MtxXloFMU9NT+vvjmF
jIdP+QCNfprI0rhsxiaDC1BJJioOqeO0D7jZfpjX2XJRW2HtM1s+NsrLld1mk0B+
5NrQAuko9ZQb6wo33FMyBG36N4WvY5WlLal1oFilREqqvbtizqU4DRGDulEzhoT1
3gTd73I2NcxPbSo5ORx0Y/V+lqnFO0eYkDUYIDRlbL9K3wM3sBOA5HMWCp5ARDE5
xNIpsH1qVHuyWg0X+JyT0fMKfNClo8qwy6fQpe/yZc8ZzICbfBahQCsgC+5pFVIl
O2Lvs9CbFyXthDV9r/T6koxP7Dozb9yGzNm+Qt+Fbr/5X9GqUOoDQP+hZVaQf8wW
qsoIlrsLLQUK1Q9U+eC+GICuL8QFJS7QFMbeMbRuWyWfJFA6BXrXOgoKAAuqaNCN
fVICrHLvcHn+1LOgu23hj5lwklA1w4NUhnlVDetUfax6rVCqOAxQ5FsFYX/lS/bA
t0ZSWFqJHNtpzN8xOVu1syUej3Ap1KMhm+VL4tZoO4NStWKkXkUYwSkHo7P7iVI3
xKgnmhi3OJB506xUYUOSDcB3BqN/s8hnEe18o0mRlfauhbzhxNWX6aT3D4OA7iHV
hoKDLx53fp3UKsmaCuhV8tq4YPLUFbmR+zMC2HJHGiRF5xnlUTSJuCiwCVT3ff+B
OMtyTIAiaAuGVvJsuUtFiuVsWnxl/KB0IonjOQn3jiySHfN/KkC+WFJjVyKISR+/
QcPeGXeFz9O8NWbUOt0qXdUQVl+SsoCaOYcMbLuIJ2d1QeahFK1N0x8QIhyWd2El
4Cbpr06FeBQt7uTDmn2i3E6MxlKPFX9Ptln/tPXLMuLM4eBC/PZ9Hau3llA3SG7A
x5TpW2ZcCvyDBcid/Hg/TT/33G5+4mmjMSy2d4gbso2bz5MSm5LmEb2S9ll8Te8h
hX+5ZE8JYZ7Lz2Im3PCmYDST7kbPp2bOzaE9JFQ1x1aFoaOCsHv/mFV0T7tguyMU
zLWawFCp7oNt452Zr7Uqu7plssCbTgCjUBhTEq8EyFiwkm9debxvTDXAbD0WLuP2
5SxeHTYNEp1yXeos2DRgDuMy+KqPAUpyo4TDO7LcwQ/ODrQdvgGPc0uMVZL67KJx
0BN8B5hPapvUtNQfQmqLvq8rgstBPUEVNn7+Y3ZUnMd0Hz57Q57D5iUFNGdpn+8C
bhBjoxXZzFW2y3M01yEOyYtvAfrFoOFENajIh2eo3ga/0GKJqo/n2AzYzRZP11lj
W0i+uYjm4wRW/v17nBiZF/twZr7h2c5p2P2pSn1jzYgC0UXKRdIDL4W6bgeILiVv
fIJzR9UHtQfpV3yPUNGQA6m0Y/pFeWT+PewlO3EPnzROdACuZ8gw+8JHhkWzUS5E
SF8Crh37kp3xocVh0yTxAowzx3/vMDMglfbt+tjzGpL7mKUXuZwZzzFP8OepqyFS
y3DJnkqypVDRBCmkN2Gn++tpZB5tTceZg4o+8Sn8jmcwCeEGMuQ2HwqnV4IV9x2/
j9tfR2YCJZ7onPuwGaI+XqKGtwMgRh7hCL41bqbt4g2oO74V+0jEpCK6Nduv05XO
dop6nqZnYXHY8RoZEkPqh0NYNwGb6ekk2oX6HNNUnpdF6yqEjEp+Vpfe9Mjceoc3
s5XdxPphACWNaSvh5bd3VK5zBJE28wiEkdge1zppE8ImA9FPioo2xKaNILk6yc8i
ZaQGnT1csjn4OHflExV40oei8uCcGC9058wMeP8/Dmil4kXIYdBBda5eQQhHkCnH
hHYF1LtOp+/N89p06hKcvagz5FEwRoseovw16UubWDNuqmo0epVT+6DjwB+3dXq8
cD+nU1TW46DPxKDPvc+pZQuf+4oIl0+4TamSl13Jzt6oEgTymPUhx3zuwwN2DfV5
Nf3/8Mbsg1Rq/DUur7bJwQ7PaZ3pIo9+8R7fDBOiFMYuVZv3g40xCkkSBpZwmzWr
9ITlYCy98woDKyTUKy147HPqjxzt/YaqVG3ga7Ioxkd/GmUgrHY4LEVGfdmMMYs2
KpXSZIkSSBYPTlvT80wLc8w0wz9gZaOVDZjWgjZwMvovJ7yNTcbc+jBsZWMtZBle
WknacW9/FeSgsCgRsQTS4V10NDhjIPkWWY/0BBAe3Du1g8xEYc1cl9QQxNh5ShUI
TdXyH6Znv8BYQAdxMPUGdUjtNfGmiH+RP6q+FAuItXwTAJ/ZfLbJqaV3smlfO6my
jukM0m3mwjLljIBNnLjH5Jh3DzZNxN5f5ZuUOxvPpi8x52LQO8GwpNf87gGWLIgy
0U+BJg3TZFzYsSx9Zttab6YNYZkl/9Jryi312DvkrLrM9qI40IyWK4CUABG+nL2k
NGinsA85LpTYfjHsjyqHHBFhve1k45bh26AkZuVEr8Ma2mZBg/8T0OGAqPQVSyF/
3RZNtzxkasg4H7DoZ44nzklnseBV+V8KK+/k9DJh9xDFGIZJW72nEGDgkr9mmJOz
jnUhZy0JsbD4pUtIKk5TrpwDe9IeMgDq5/UyVKTCVVJ+//AsSIHgPCX6BhhdoGsn
W4FUfPiSFEogLnjOx1hCQ1bzfitdgqSFPRqrEesdWA0r8DDeNLFX/nYIlDKWW8ld
tvM7aVeWxjIMDrGOE79tEYapHNaSEQt89gG7sjeFMd6LRiV5cYih5DwQAxBTk0LD
+uMpB6orZnySJWIkshmHylVzyjErIfMrf2/tR58LqC4d4KFBVEgMsuJgcF9d67cz
SomxjJpHp2aLLfqAXbIYV4PQtI7zjROCY+Tf4cKYc2+DpoosDtAKzDYngDwTJK8K
ZzIt8NTTYyUx3TFhuwvmiVNU86K3THLROVE36gAX9iAWGVrqL18POb9AYxSw/skJ
pLJNOhLfNyfiUuA5xI5QGxCIKMq9ojaxVKInBOjy2pWSRhKhlo+362/7GG5+mZSq
BMTU9X/Z8lfc9Aodu+odLjwE6W68FzJBP8jvTMvqG4+Z5XiZgowATzC77feAQUaD
y6dVsWk91wqmeUuic0qOqzpuxIsDWXHX8EwrOWJc6zXnBJcSn8TwnuKP/VtLuQyJ
dbFABMihqVkLdaHcE3sD+pJDcRk2Bdg3ehj1pTYbKS4VMVWRsEj1zoJERZm3T9RB
ejDo8Vrie/HtwKdiVk57n6QQ1KkGBjn6if0BxrENsYBXxCDAw3XZoWgmqLKsb4FF
nSPVl5rK9DxV8RxgTsZND+U/D+bLvZVcYwypYuf1e9axGPZprxPmlVZ0MBY/4uEi
UjToLva1hLTv8YpireMu1e0W1+27ExWtV2WbKrPPfxdA3M2BLGVI0vk58RJZVTXS
yQIv8DJcMso++XW3gAvmRUO60ewvNQjyfj62KRotfIxp88KKhEPXBKJ5XEhi9/UV
VV3lupkG20LvAjtpaQR5XY4FkNRDiUR0ydK5S+2EvizvP/IF/Ftz8831QMTerQKV
HAnPZlI5Dn9X9eEJ23uy1YxkC8XKTln1UZVMgk5qCnCnhcjmTi7gPEeMZyWmux8h
AlQoxjyb9zBaukkIpEtQArRTxgIOBFMAQVCnEG1xZdI+xaZiUwmkX1SfyAYYklFS
VHRsckghjSqwsy9Z2FSu/WgPkol9IPz2tVCiZF0CMfMBbgcNUb7+qjGi3RLhJ0+z
uyq//wB+cWIYMBlBJsM7G+Vrqu87p8qJYfQiPZBYwGKZoi6k7JgsJi+fYPRnGoFK
X+43Ie/sS1Lcd+2MmItd0ycBJN1xVIbpcXhdKn9GmEOpHn8r8S9f5qKa7krm/2H5
MbbSacdhH4N7iDmVc8WX11i6ATu9tqctwZu+w8PIio78w4Q4c7qhe/H04X94s0gi
AHD5Vi6pqCiYinCF7zRrm8hVCIKyl7x9iLU+7C4v3FpL1mpDG9+sQvVDV8AwkxNE
urTHnZcc5wJH8z3aZfdXtfjGtF6mJ+bxZU2DErdE80bm15a3PXTon1XNM8/oQp3t
NkRhh4bJvbIDUlgVQcKcFeidsTPDf6hsNqJFcZlUkzINq2Krjt+BnqlsCzklxBZV
oRSYbt4CvwbxahGj/WXU2Zyekys8M2eU7GYrgGZMk9cNY+53NEtVFk6p85riyFEe
74rCE4FdTHzKt0/ZFv3zgRHJplnDmKuFiMM0FS/vTKeCTSLtoZRbJq79DT7jYXxV
CvI/Xsjn6kimCaxN3U4CS1u1wg2/hTSecKKxd1w9zierJIn13etuz9VOCPR8/XiG
usIZg4YxIrX42W1CC1lTBZHHfsoXE4joKxJG8fZpjBQp6156jkZDaXFD44NARyXy
Pu8X06dwjKFRe5NXCl0FM7kYRgaRDWtvVnKyDrqX+Z51q1J9/GhqAfk4Maqmd9i7
NFzOIMfkvNMxn3HGkGKBbCQmRGNYMZD1o6eF5Ik/iziS2hdLMxVbLAcojbnx3hw2
+XlPlB/B9M0QAxwTltrcwIxI+MDCrW6k8RZ/Chuu91I10mefIGjfp22diYMNKidv
5XmSE8Iv8I6Yan7sDv9RjzoTFssvOFl8IrasAFVWQsy2vNz8smswTNpk5Yp9Te7s
QCed+k2FqnfvaC0GDVWNnwRqw+Xiv0Ql9zjDIUHL0bZwZc+t2rmVs0uKQwg3jbvi
+CQ1Yj7brd8inB3lAEbdJwV+cOIFl9kgT+FOazmRy6pHMpQCklnnUHciBKpB+uHZ
bkYwoimE5w6c5EENeI8iBZhGK2rvR1p+UxdPhBgo5Gv6yjeZZsIXJG6pYivuMM1R
MkdwEnJLWQIJC70PHCk8OaLePANlb5Jhs2m7D4llTGF9lOI6jx8Y51nIP8mTxR6h
FD0+nrSFPdgB3fN9fq2Df3uCte2SmHnYSQVgOqwnIlL0wncnBpzfx6sZIEw7Mnp3
5vzxE02lBQ4AgZz7+wrZSy78pRdHF5tgD15UmR0bjFgR1m83HWcpIiEY2LhD3S3H
vxobCgj8bxAkoSh4lsd5IRS88gxD9pLVN+VIUZ3Kals83OCOlatWDDKTsHYJOwWs
yy/tUhCrrfBSh3uXg9ET4vmZMJNrd+hVxyLr5v7WzC2VYLneJ15RMC/k8YThxR7m
f7DDVl1he+FGEktr33GqZV0AyLqXNO7tM4d/2KoAVLPJaTeeOLtJp2IfJusqj/CY
YsLxqhuheMCLeS2c6cDO+UTWSEYLmW5kl+OcHNntaFb1oMDJjKnS97dQVo1Yr5Dx
uXfDDkctIHxVSb3b/scWByM0LcBQ3iFjMIosyRKEgXtRjm+mMrIi7hiwtJ6jGS/I
wHK2oJVEy1z4lKZqBs3rQw+OmMMPb8BYPhPsojoOafOMsuTUxA5wVEl+m+wbxCbd
3Hmo8nq8ZZEGrTbmczxk0qmk8jDKs42ww929SJSS9XwZ5RC7M3oUnWO4G8GKJmZc
aXuCemYIQuVjV97A1CdJKp3mbGSjZKh7byEVwzuoBWcYT/ir1pIYR9uLbl26/bPW
SOF4TRc6jMnMjcvD65Oghg2F7423qlhbF0x5v2P3zvVlYkfgjiOhzGx9GdPs3LFh
Pm4Iw9q1v/EDSDZnJJUTX1YSwH/ncM149hQ5fE1FAlxaudXJs+N6DfI/hBjHW+o5
MxhE8rJSMDfVuGleZeo9Bit03VQhnFjM7mwpVc97AXXTbJVXOVejUL39sNBzq1Ib
hOY7oqavU3GeBgL25YwNQ/xZ1Cq51lB34oHOqCUmnniO1yhTr9q4P9JwyWPlAE+K
6y1NcRvGyrxlUcU50oIZ3sGkBWhMqhx8Dolnu9mRAcQHjVYqUyRMbsVAfOYTNsEX
ubbLik4h9HrncicYL2pS1UwFHmLmtP7Phe3DoXXtfCfwhw4kuk6Vmo4fx+3aitDH
BykmVQuWTlY79oo6LTVxhlDmPepAzls8iRuvJ5BVDmK06DQDi3HuKq8YwATEb620
4VWPW6KCy3uoHqDVYHJjmuy5EWOvm10cRL9ky+8OIHbzCYLKHk2mc39UQRXh18wO
DzkmkxKN1CrOWUNum091Ly1CFYNJ30V6U0moWXjh1k+CTcPInFPUFdGHZCBMBqIW
peSqseaLno/x+jybzItvXPxOzTkuAAcxrrYs/Ln6AiqNbL1UO4N7xiUUGYFEgPz9
eacgVaY7LYVdtU2SK/QJ2mOVjEmmqfrAKRcYQIiT2j7wnh+L6N9oyxP2OtQ2AhXZ
JSK3HUFC3jT1pjMD6bPTz/uszNTmXEvI5v4tpIrWyv0AtO7x+bzNNezJi3Sq6kYb
P2aN8ShdQdoqtC5XYmJCM04mtyyDyj6E7wQOhPqahozDGwVlMbjsdSuOMLHoyYkG
B7unF09iqDHbesGB0s6s6JklC2Q0Uht6yZQoMFdo/82Lki+TsBdIvddMy5EPoH4D
E9NhgtuJ+UkCRCoFPuyK9GZrATOX9/+8r0s/SWtIBzwOljJW8Po4ZOWaVkjROgm8
XeNXVWHfK4b55KbsD6mChyCy7EH3Gk962t/eTV0X8Gyyoplfajir27+ZQfDtccNz
QYO+Lx4i+v9bEBjalkL9yGvYyZl+G2JeH4ATaWmr3DQRbwsAFbx+++AYBGnMnakv
ssfOG8Ua27mY+LbrExVWnVe+pmypdF9wkhIhAigB5sDNQnn7WVg8+qypS6kXfI4A
O8aQ1VOeyuLVZV0qXSHbyHgz49QhqExImK4YfI0ymcmvV2vnyefERYxsg5dKPVbD
Pk+ys87gox00Q20hh6AV8LAtvab1Y5OVYIKYXd2s5DzZeoULFl4pFg8ret6g/Gh6
55N1orBpNbIGrSsISds56B4RydgX/klbrEsEJF4cr2wSlFNcsv1xvgsRVlCdtgbZ
DapSIvTOwHTbYrJWz+0sDbKCYEkLv+EBeY+h/HIE2LiCMr4Gbrh1zLG4BWKJN6dn
wIT/HhTKD034OTpsQNeD4phCyONyXbSBTNqmU6XnJ11p8GoXQffPE0BgqgF+aKXw
Jw6Oc+BpzVLqt7N5HO2z3+QIp86eO9Ll/Dz6M2Xl4smTWkBLb/vnek7WodpwgnCV
+N3xLShqUN/IwmC73Ya4A+Q0E9jSse4MTPfimTwf1AJB2pmzcXSzDrNftX2aknel
nrbmMwSjVZ0GZQ8VS7+Ame52q3vY3ZWccDwnF2yc8JO9Zu7SajpP9lOh8slkuqCA
eSMFE+ELreeBG/SUmLBzOt66i439JldzhIU/K0O4JE8a0rm8JV4L9qVAlm0kfuWq
BUXfZaGZmeR7jSbo6XTEPrlLG1qpdx8v/PUXCtN4ddr17SIkPmN3dQssbNCgDhJ1
UUnx4nGvgLN6BSeZt0/pkBRCb/t1yUvEEE8LnNd8TT/WZI8bdx4nKd3BSYE3iYO0
W0Oc0Cn1sR7JN8POEnTcaHqON7t4lqm0Ai7MmHQd7sDYzsLmz+oD+qz3BphnAWI5
/wnM5KfXounILgWcMWfnxcR44dYKdO4a23lagJX+8rIF+66izFKjvUs0YiEwx0Fu
8ppIns8SbnNgMVvtpsUDHvCxG/+UuM8AeydxwX1dURmK0VvESQD/eLwxtVbVYMvO
MAFi4wMFsnjkZOYHuf/IbchUBOYQrknKK+uutdu/3A5d/8epEpGHV3xlMOqtZTZ5
67zEOXxqRzZ5qh+tAb3hHKtFCIvGwL7uA4KnCtsvogIaXAlUCsHcDWMl3UOeqwbA
UWlF6eKqU2X2J1EhtARNgi8kn8dgL1SAn1c3twfABBPF8YMXtI76Ysn5Rnw63JG6
MHCboIGYJ+twkwlXwi21m3T1sfIYPt3TfCRRkKWrQsOOmXkD7X2Wp5dbIf6h8Xyh
P3E+IVwauLlrlIpjFTohBqy96D1FXHyF+8K3p7lyaRW7jaC+siN5hiO3fZjkL5ND
Ovvm0MlaSEFnERdo03tYNgSX1dGtZ8HQdnrQ5X6nnUcBlLiS5pitla3gvkHJm11o
B4sC5av2egPk0lr7W0rnfrFJymNI4Lm987jdbOqjvZlbzE5vBQsGT/u+cx//AQAi
xQwjEbYtRBVAWMN3Hrh7YWDCC7LHg3x4ia48+lRnErWYRhT74tyzxR4fKCT8fSAn
7yGs/L1t4zx6RAZmzIQNfMi0DaQ2NtQspapJI9UWwvebmArPScArxDjPfuY3nMcu
2sToLkexokCsDmpjACkqPhYLmFft2XvYOJP7Hx7VLCWHLOZAQKmaXro1gSdSPxR8
jjUznGRBZjsKyxArAo7ucvhMMdbYQi/an6ZEM7AJ35Me68DHwI+YDWjF8GbZApvW
pxm7qiq8hkN7w3JLTEHtZYTi/ZGuUNU+jfSfoast5OpN4AfilS8+XfERrWkEkIVf
wiJdMIzC6fsy7tmsSYruGXadkx3QW3Aeso/+94pGNrbKHqvZuniWcxJxs3/X6wlY
gY1zNR+SCg/+pnh6UG8x1VQ9+aiQneXR8d2l8GkGUOTSq6KBWGj+Cw/TVTd4AwSq
Ad9XHdmu13Jj9G34Orm6/AUDrjOTAzdeEVsAo58vUlL4245iQ5OQMjHKygsBpkIE
Sl+SAqTwxaN0Hq/J9zvVHbWUoHpcf3SwWbnry0DVbW+yF9JJRtTmmUaRxYyN1bYq
dcYhj0qTFsH48V5wGdKmjIUBi3cb0O5FRGvtdJMzVu3DhYWd14ptO5lqcoXQmyNB
FYdeDbPHukzXFKK/ecb8iTFyaaSPsIm3Ze4P6q42/kMbwuTadzH3QAV4knNhT1th
+T9FC8uHjYJRXysDuz30/uI3LOfvkgki1MSnLSjPWzICsmRgwh/OWbvFXAqK/4rv
CBZzQIiRmmGsr0YCLhH200neb5SPG4uCGpuvgPYY7F8YEzbossWF3gb5T9da+VfM
+dZTaNn2V2KgJhhmpqUr8PvYhr8n5x9NrQmu52YW/hIC2rwZdG6aJHpC6M2vaApL
qaHHCOnzq47V+F/ZFIqCmsZnI6i0UhMDeu/D9xFu2X2wVmWdnFIyiauqmuEmbPpA
RwlHFP+XImQHy+1e2qXIh+kIe6SFsSedZpsIQc4H9oOj6VbJgmCeEbDqWT3cKZHt
ADevKvKaGv5oDo42T6EXvGJzoKmhbDqDpBuv3N5pFa5m+8CFWd4/xvrRl/KfmES+
BHEnsipr0btlLp7+kOWbCNXYTBjH4LlVT15GRF3dtnCQkxjkfapEAxbs2eY6J/Ci
X2fIa+DOoV+r+NKC7ZPyd02BIiaKXFTjAOyqe1dCaLAx6xs5VqFXkLRHnn5JYF36
VRa7e61OKyAxwQLl1vNZdAmVXBFU10R4A/+PT7ZuGFUKM0FAozRGG/ICsg4czu3A
CtdQNStmL5gXOibJ130atA3uEPwAVc0HTW8w/o83dJBCwvzyBNLP3PGeSmRd1fO+
k1PY3fAbBoUcaJVCW8ngXFVGTPjm3lvgcIC2eumE3gLPU1/QA58mjDemrKzBLu7i
goE+NglPSPOjIMjplNip+7fhJfCMOMFXGO/zQ6QCUpiQM95OygbsyGJyKmhe8rtM
yr0MYN2JVjueIKYE9vlp+SIHQNbSkk6WTwVfJteU6CIKb9/oyuCbH7HEWCuM8ws0
AkJXmVfgUBEIdSy9dI9PwV/R8jgZVy1od9DX7yUuBu/4f4SMMC7cXhd0SFPTklrg
nx8GXb4T16tidEkgox/VLWf9+pCe/tKLqSLKjSIM/22nUmE+WO1yR+U1Hp5dJR5n
PxVj8VYVxp4qBnN7EKULaG8DWQSDEhIwBro/v6kG1drUl4bK/jE4bhSTXBwh6oPB
1+SBgr1fzaOPW8E90qu+5BmT7AKUmVMarQrO9S0fxgZE20qNRq7KreIIeLUeK1UW
Gs24TeA7o0sVfaL9W1ZdMmQ96WoM+BUSFQVssGuj/IGf6m602nXPJy47sJ+y3zcf
aJ55inQMDUI8m3mxTAkz/4LURC7hl3TgG9na8DQMI50mZEwLaY+G+lxDzENrenJ1
yyPBJ7EERLUgeh2zzdmBwrl/oRDrqqxSLwyOP1wmc0dVprWwgB9i8QvMfMtSz2d0
WFuNUorc6gMMiq9DvJdyvMPwy6JB6808p8vIls4kbWlm/UbJl624tcnmOq1XenYX
HuYSUeODW9gf4HzaODGgF4uIopxvxr04rQlqaO94EZn7yOTMetZE0sFJpnCKN5Rb
34X8r09DCX14sq7IUsTBxNUQOjJQhmpgwrU88LN6TIYlE5qG/N2VFPpsraqUysF4
WTiYmMLxc4yaupMParOW1iVWlX6he2kAn/0mqnIpbHixdDj/lObg5Y7gk2untRDi
eDoLhjcTQ36F03ymJP4P2sOHDuwrvMxr7N8YIwL36BDQl3t2bg2l7pcU8/IyOKv+
3PTqS0BynJuDgjc2MQgYeHMXGpU1uHrPTa9hrY+VkFLoZrWq3H3bpVSsE6w49J+p
56gYKMzsClUQuCidl3rmNQMdiTyZJibBoukNWktENy6LFfSR0Dy/OfAsQ3LLwk1c
OPShb/Xwu8p2OHfaxjcsPY9imHv0cVK6YwzhZ2N85h5VorQEt458Y70vLmDV8rpu
6if/NA3LAwuk91Nc3IM9zcDmdQ+Lta6mNAN58iENUMdECR9JeAhW6nRTnoJesalX
Bq1eBf/ua7QHfxZJXtK/D4snfCOx6zazzTv2W36L/Deq2nXOAX1YLyvKT25bAM86
xz/PwPwfDKflFfOkPTWkhX7pjRGYdsTH2VlvsayoFo9r3EwArYJ35wOMstFyEOqJ
hZTXZZ40BgUKK/70kQ2uozBvcnezgPbph1E6imQFG+nJaqn0v1bmBHQNRDzwBKVz
RVHcT1/10PCEaUPjAyxLGfIE8LSjnm9JA7uSzJpVbobGeljK0L9m/nqzTDBCMGue
Ee9QdX3Ow3MAgZ1WuFr4AgdEGaIkFD0KyvxhbpxK/MtHlsu/jWSKuiStvEvDdK70
48f7px88K6a5BPHxdgFBpJ6GvPXc/AyeYGLdW79yf2woMZ5ArcndLoNY7p4wIAMU
B+fyNngSkpUJfE4efE2oLJTQ3n53cpFBfNh0Xs6OqPrPNaDhpMdFgeYJsVmDP6eH
QBSrOVCyvVPBLlAFRS9C4su9m76nekf1pBvQU7/XeBGu8CFHThykVoT+UDsMLfh3
VbB0+UiEM68r9Z3SsCSBAhBnRf3GFzpKjmNeWWhg+VgPJMysRtvritYBIQSTrfox
9+SK7nuhuDai2bxBHBmcPrWrq2VTtu4W4+/gT/Y0zwQiTngw3H0NW+NhST6mGOij
TofTyCiiIa4qSFbJlp2FApqtDFJeNM7NUHW/Uy/aVb4rWCRhcB6oyCPyvpUenvaA
l/34h2n7w4KCJNRtzDSEocfMYzhxDGG28Tm0YiKnZDj37qK/KfaFfwdhhDG0De15
fIRKycZ6hs5n43c3NewTi14XJXE5T0PJxCXjzoqhHIhR3TBp9C5HqReYXensdTmu
sWtafxtRa2Xc3MRwx/Y7ZnIAZEIcqb2xk8VaOaIRcQAPjw15kAAYQkSZvsgm7H5S
ZRtd9+kxHMG8SwNjlWz7jFP6BWrCFqSf69TYcjljP+A4kziqW/n76rpnzi+LlLXN
IXFHOrbs78I08vMwuM1on7NaSEFvpZ6VygYs+WtXlbIEVwcr7e7g7TMwvZx8wBIh
X44kblQ8ZEd/s36c6LnaBVNC1RmKE49awssbuaeQlvxDVC+LnEojZZAN5Er5pRv6
N3bxveVy2k8dLyVIWkZyp7vFOqxa6idfOJfWNIHfQ8ZbKsnCtu8n+2tyTxELMTwd
HI/dzwiBL/j+6M5gb1uzQF+D4IekRQYwVva+84Z5YneYAoHyKOBaz6O2EWkmxE+4
Oo0Yj2x4CIhiS44JeT47SCqxmQ3FZk7vAvxfl5E1v2GU8whgJVuDVFQX12KkWp5y
IgLw54YAv/eurFskkjP1xAiNRlA1S5QBKZJZ4gqpb86oohNe2BA4CSB2RODr4LYN
/S3Z2YaUPZheCsOPtyknRzvnO8oK4a9yPVUD0X2cTWnXixZvqkv8VFrr5x4WAauH
+hHap3xHxrR7Tbslu/uJrJl5R9NcrGtSGxF3tXWPmcNF144SfwCJlaaESI88Onr2
fHg6Fq0ezWpdo7F0pTY0BHwiJOjuGyW7OCOy8TxVKeskjItHY76UCYd+crTBZjXW
Wt8okDp3T+/7qrMz1AkUTZ5fkqTlxhRs8EHzif/AdeaWOG4q3fOmnZYEF6fOJQ2b
A+pIrCjDH/+7JxGuOtbI9oq/CD9uT09dkRYYYE0r1HZ8odOYC7+FQM0lFF80iLqi
ErvJH3MNL9Zmxju/u4FmBYWSz7NhAWVQkG8//SD3lZw5DBHjbm7OgotrDbcwRQHI
n6VBDofiYo1RA6zs1XFs6m2SHFd1gukFhuZIYhPdkFDdyCAPXEN/jGAPBamrlO79
xav+0qYsXJC/ySwOmGQuusSWyg9u+NR6tDt59Bfe7GbhFZWCPZDAdJRnWNSA30bt
pG3UiStlxHwjowclJl0elnwOeiYokGUqJR95H10LxR6GpoJRdkbUmCGpe5DJiuqn
L41wZj1FMlRITHi+SwrSxcXnHub0Ygh5mr5Qe/Hiq4V9hB3sYYb640S6WhLtUngj
s/qYtB3ctwxmd1t2H1iXuzwq/P13893Pa598g+LPq2DafdvEHRyH141oDpxGaizr
LA+jFtzAvxYbWTe1FD0hyluQ7yCuhNW1eASjSv040RCweSm5u0JX6VJ7rYl8h0Qs
6RCpZn4FNJfLQt93pGqas4vtN3KNpVr8k2CAwzwUKEZOdvXjkmfEueCpGCQc7k5A
lh4JUlgorw1toTll3awyfM6YOMwtYiCFgslDDT8VLBCJgqBy3A5hn0UEVxSjvXq8
QyoxjdidlAi2NIbBnZb4G6Scya3nf6BTniNw3iXd3HFjm8lZkhqs0GXDFLYeXe7e
Z8DPXp3u73mkVnVEB2wzpcidCOkNceHFocgyhTrUPPZbURTGB4pqsBCLbehQjwTf
hZ2hI/bADnuevUpjXgm0EKd17GBIDt4vMxiVr7kIj0I7o7R/bTING+Vb/OERWlhe
6JPEjQlg5YeKoPSwSmbNxTxa+XdfKy7Cak+NMjG0o1nXjA9uvCszvYZa+B+o+SKH
dqhsZWlTj8um9awKDqOM+aPKECOiq6K72n1AD3AupRUOV/FqaWrO5mdQz7d/nHjZ
F1Deah3gsKub8t3ZvsT+SkHSwHOKkg6uhDK+WZRO4GDWvDs1qpbsxIfLgIAgdYcP
XqMOVIHptOw0lTKNPuPpzZ/vuJFUQX3fxX+tQizv6b/JYcvVrD8YcXeY5SeoiMl5
khzayKP3bppJsJcHC9PmN08ehjQ723a2Z7f9Xnl5tJYkRT/vMqIKiPHX1fhBJPcA
XD8i7/UB2Uf0jXGiLHOK3/01XLyiZVmIe5y+/SIrkjD2iWzwK9Rfk9lX4If4TRWM
H3J5UAJ5F/5QYE136tyAAGuyAk1jk6NPfVdupYBxwTkmwYKmYTEnj+1coA/A+RIi
25mkVvb9yI3T+Ac3ng72jvU2J5I4E2GOcnzE0uLgSGS303DiYlXKn5tmpsi16pF1
2H9eqMW4v8kdtvCOD5ybxltF/vNEgeDPyoE4FyMC3NpRqdKNgFrxsbEd7IlygmK/
tWjVMdS7KPSW/ANXSSHZILMHg4UFnQ1/xfgJsMzEQ2IqbVfv2w30/GjbhEU925+L
cnoMIyqO0XflFkwgUC+rieogieFiUKiAD8x5/9jbAM9L47es1CwCwxsqzeV4FFaX
sQgA+ZqKSrXmzd9OcgW5QR1xrV4mLaFMpA2hKKiDKVhul7LmfXkUkyaI2Je0Cc8j
8MM8RSmGHS8ftmiwHVH9DsIUrObNZb0+kufGez8Z+whMfpG2udmeoQwkh0Ft7i/S
Dmx/20dHtKH0J2oE9f9K3uRxvFG1AG7eNkmLSaFQ5rxaTbHqPVQBjbb+gN/SRcwj
YZY9ynIRy4aFyeWuIkxVni7hK51qyUoNOA6gkjhKXTIo8MSXYBYwIth/PGEDCXd/
Te4+czXoVjU+jB9dnjQnL5Ah55268nziXqpawLNKjN94Qg8dNRbXIezyuRfUQdBS
rgjKxj56z5JUpgqPUbOdnUUtc7xko3vHXwAG9ZBgwtP0pEOZSCeP4fK5VZs002vR
JQsDQGxKoT+L9NI6CUKJgFLiQK5DE1CryAdiUehwZPN/P04RPK7mNv9pJh6r3Ptf
dRIcbIJnPi1sEML4zz3v5sylOQmijZp4s61Poy5r4Xt7BIZc+zYNPnV87cFzl52p
GciJ6/lgGBv9BSot9bZrLx1y6sXRIMjgql8FYDWUN3u3iaW0KsSv6vdiI3euFfn8
VPCHBz1gCiVQPbBAw+wOT5zRAnKP0s4lkWEq65AkdBL0wAVOI0eY5zVEC08845E3
6iZ9VL71KMaVD9YcPFxidGSkGksaSiAsPhrUbxW4ZqEMLxReqsmZNPD7Y60+tadE
mpKTL6A3UgI/ZuQhbIiXyV+Ke9WCDdZzd9GoeV0OqxB/fPgJkp574y31s8cf4klh
QRlMGsaxPFfyaZ+D8e0pYjybhWnvqewJvybeJ8t1bFWhR/saDCuq0W7P70JWSVIS
6Qv9pLnf0DdmfERti0l857Tasv2/RLYW68aOMQ1yDzYKLxAAZDLo5Y1JteOBFtku
NM++v9KnASNH2xSLO4cUZ/XKsi/csT5cXWxXttoyDWbHVCubeGzlgONG+eh9vsRn
WiXzKaNW0e/wttOEvmoQ5zf2X7DtM2dkg7nF/EKWR/oxlNyK3aPIJtQmsy7ULIbd
3+ckjqc4gWfP084SzY+l9IzKZILAB1eKg7CGf3qn71jt2fOIi3fWFqALI/qL6cld
lpKiuDQvDL4HrbYO8ZKBEeYGv2fijboqJ0rkqxONU4WXtz1rwfP1BaFi/pqZ09Nn
QxzANA3a5MXf2AXLQpFvzeN6Na1L32VfHSAWncFyFBgIyuWfG6OiPFsoKHTnnKsQ
cufAH8L+ujT19H8TJR7H37Uvqyg/FkFNjZJ/H686JUnEWVX98qZIIM/Tr6S7rf6N
C+4ZOrsuQzsrXW8L0+VrOJuxc31quNqHVdP71bM9plskFwXJ0AkyYI2+w3+j4khE
UKnJol8uyX7h3iS9j/WNXfxJvASlFr2zw5zqsPsxO4NJYh/iWra1ueqHUOfatY2S
6kzkt7bcsF4CVdr+mc2izxBSJEJcPAn79yH6sNwv9kKMk48ostzUUd3Jhe3f0RYa
LSOJL14cJT3IP8ltaCokABVGiEbY+dnkU+bcyGPMNatV4axJCFfk/wXlvhAx8h9e
rHrLpgOXgSZ/pIO2SehZZiWwyYmm8oLb8SbftnMsbgDDD1aOlkr1ROGIGoxpjb4v
KShFjVjFrU5UW1JNaVP9qlkz94ktCW8smtwaXASrDzFBS6ZxFhpU9oTdnDLapDpP
Qesak0Q439iAuAkJr0Qkd3c4oRDXQ7D4rUPimCDizfeBort8vCvINQ8XzftlvdBT
VG80Vx3XZ8fV28hRSz7RPOhFECvGWgHWDTIuBLiNBWenUBfusKTWwUNZgHR5+Xkv
64N0+VRd5lvK7zrLRlOiXqYcagbesGoce85P8R3sBjyZHCjWhB5/g5BfBWMCLGI9
XNJjcIWR8+TLCO0bzr28IU1Q2FVgN0816wktfyFY5eWmq09CLujjcLWCIw6dWcB+
2Y6N4Q3juiPq7xFzJeRPNCxpwh2FosXhsw+DwVSJ5DZFhb9lbknr0Uu2a8PDzdET
TF/tVkFMnUs7yx79BRvBbySalkBBEvdJuN3rx2YOLhzqSMRo/FAlQaw1CjK/7SHf
m26DI6gSNdYmQN2dd8/2pIbNq4Q3u3FP3diM8xYH7K6zs2icojmvSllqDezR9TMb
CZApSuCl9b/6oF01WZTE72Xn1mXC9AZwQOUdE21VdgzikOMJNqG5oSByqFhpuU3b
Qyw0m8gdDsTf98AGYuvyXPAzC8865X61ROUg7l+e7XNewKkNhseDghDFcM0tzMsT
mCsNp/r1JKSh8Vng2qhzQE6bZLUePsPD5KDztVYgdv4kYP/d+wL1MppUlXJYMScP
xx0I2SCV7kQ0KJ0JXCbw+MZ51D5yQgeyQgOGHiPCYIxvmJgvXYrK03FIN38g5n/n
cF3Do/24PBggFO8G+y8IHf7Hy/gj8lFUYZvvIZJ3Mf4u17aEHejHvsT4/3hgIsQz
VzbIpKL/CLCHsOJl53KUCoWK+/bb8lgbk33LZhTUERFFg7+XaojcBlReBMcigM1K
f/sfO1alwad2oVYauihdWRLlZhXlsMut7OzhcD9UFXfBnOC9bRKWG0Gl00urCymx
v14D9zzDajHJct9lzIyeGzXMinYkJk/51ELaVjzK6rTzgGs2IjTmNuhJbxsAkn/I
acmODzjZ4rR0ZRZ9Nv7Tf1OF88rNtcxT00/szSz1MwbYDy5C1Y+LEgGGNBfSkJhN
qQ4q8NU0OqUK7VC2FoXisjw8LJ0b3ZXxPpbdYwQps7HYYXwPokH0amZR097rDFl7
o8QCzRSe+lvs72ITRHHmksmnLx3+1ANVh7VfnDLggmF4GWuZxJOQVeeaw9BFn5Ds
3i10djsktkaIGKpJFcsGDNBz3tSFNlXs+DqTT6FVS7srESu+BwuWAgNi99/A0Ksk
0EVPssVZAfif0OXtFjdcVXlaay27/OOtXPJJMl/bqH7/laIZ96StI0oQnlR9vjJm
5gwqX9H+MK2YdgU/Y8PIoR+Td1IaEYXdk6nmekVqMsB0rtpUcMVs+6/Vdp1c546M
WIPgHG9qU+8VlK8Abk6VG+ZPbuRO6FINrafOC2SWpIwzNkgjnhw+EE0J9VFy65Pw
dvYwGufUoh6zzsr9D8TAwcfw2mletAp73yb9WlwcvOp69A2BF3RVj6ogBSxRZYzK
yUkkLXzmKEwXtoPG0s9DoqMDl+vzzc4Eh+YCL196d3lTwY7N7VXTrFVN9Wckx0U9
VJFa/E2jE867V5AoCi/wQqvQJvaI5P/ibJkwO2Adz7gK8H3KxaEG7+hMI5A8tVfC
866zdr6M3fp2YcAPCmrMStMRfvxDyEXOx03eNqpp4HW029fLmJG27MulyGoqESZA
cokD2QCuxZbQzo2Xu4OaprssUDgDP1TCdgt0sxUHuTmu4Xo/eWuhwWGsgIIaFz3v
9huuvahCOS9a8NMsnccmAgoCGOP1/nDoU994fY1ggTpIwxBzWT3e9dxfty6VvGZ2
baKwImIv8eK+lgwjI9UpZSGbI4+jXho4elfa5eCsFL386BSXxnGVpt+OqRC7ZP8Y
kujjZeqQsozWnPXmF+MfFnnlg/o7Ey9mB62QRxyWRfXFANeEXIkbSFypEbyVqjI8
pgDo6kEEzuG+H+gaYD8qokPqW0AFzV51qqePuoVWNN6HCdLhGnxBrjxynfySgsVQ
3jH9YcrQz1u/is+traYPUKA6GOjvXBW3rno8a+6IhPEnFr8J2WxhtKr65knaMRG+
pcZlAeeZLGB89aCsupBaQbdLEhELVeQ9KizSP1QQvfQ3qUxfpo9Q3BUDRfU1T1q7
P863+GnO96DKrXnhc/yIkfWf2KIBA1PcqEbruuzRT4ZwSWPDQmHfhTEzyBk2tX41
yF4YmYRirDJEgLfazvcbPSSdT76+AKaCQeAaNZz409/OXr83jisqTy5JQVOFyKpQ
aVAaEkevvp3778XEg24F7IVHwjrl/9FcjrHP3exmh1uSks7NqLI+o0Os+kelqi+1
MWilyCaAsgQqIY7Mvj4IH5Sf343n/BsxIah65Avfg/QHh9J++g24zJ4RQZJ/7Qi6
s8UUECQKYDqH7xTAS1WiOThN/ZqzMwIfxNCo95BhfRDrX5vssYQZIg8fa+HE06Yh
7hO6AJpFrRj+ExXUzFabiDMtQcj11YFJmOjET+MGhv61OZH65Mez3b2r32rch4we
PDQpVXtURiIbMzkFoPgmTuuUZjROUSGEFE5kFjZcJTsrfxheF/O6G9NVmfr+teZw
NVZrS/0OOxStpRa1hqi+hEVYsGDLVWpLeTpzUEUDB1O8wCEk45XfSxfAeL+650G+
nazxImBQxpa3YZ5iXFIuDhrLHE+YASqt5enLHXKEuSMaOF9+ak35TRX+OmB5SC4f
l44Y0gfXyAgbTcCAIjd7LSVsbLwjnZzS6FRkOIlObyps2RqTGn0oOToJ/7FJPwvb
hmp7xdHemRa2qpBzqeGLpq120XNLt81ND3IJv4xOTQdQNuEBt3YTfOKUgA6xXZpd
TEpCbexi0mFEBwhKII7vfZjICQ/2ZmouROVX2C4imsCs2gdxxrX6TPftAtK4a5pm
Xyc7c8MFAD8rLnwBDwt1laSY7m/OlnBCImiy4EUjoP9dRygRcEKJ5v2pc5x6F3vT
xdsA7FP7C93ufv1RYcyqqaBSlSytJC7jwEA44Is30UNYx+Bj0ra7B5B8OF4NOS6q
fh0c9nlmXWZZekpur7vHFfEg6nxl+DS8B/U3bu1RIYDvd5RIEayogPMCKt1K6iAu
DSYrxIPCq0IK2pp2pqXfPybA9y325izcm2IbbLxN7YSO6naZHE8Y+jAfPz8YXM6G
KOyZrDAWV6QNgDg02sng5GjXAZP58gvP8LfZeQDD0MUfs3+N+S9wOmX2C0QEGjxc
le/dEPqy5kaHJ7Omd7y5uzX5sDclZSywzRiWubutzbBYhuwhbi1KZZfwsX5LoPKP
OzsGrH4aKABTwZ3kII4ecEjCN64/KWRYm6aXi8fPOOXl9hbU/kwqf6GewtvxgqTH
25QMzN+GIcqJBtr+8HpAr4YYWes/ss0hY8RTLJCebYOpN7I/n8BGNFdyzZJCqLCb
1NspydQe+JD3KlNrDIWIdwhdrnA67+Jjd5OIkH6zTtrrLFeGi3Hh8ZVw9GGTlwQe
BVh/oPvV9or+PNqoxGt0bKC4jwVzqY4jvEKjZ9CtMWXbkyVEhhlXBlylPZS5tB3w
Qr2Xoxnk/zI16fOHNockMHgszEcNIj26kajiNOM3cR7zuEpj4fqO3Pd5pFn4ecSs
9rtn0ONPN2BTOeyPk2In7SKdbR1MXEqF3/Hgorwrmz2SmBXetnQM1j9BEGfOIvNT
sGpT6YY+o/RBKjA6hgOCCMCHJXIp1Rdjkhc92fNuX1P2bGoPpnYazMYgvy7Wd+Yh
6wkMd6Zhsm/2NTUOMUaPOzH89j3fPQvOs8G51sEbWQeSfSx44UzGffMVcz/CqXqK
vRiFebOvuLkl5xBParkusbQAJhAlfanuH79fTYQRhUL0D7DUpPPQiNr5ubdzIRec
OLv79znbCotDAPN48qlCOowUev2479/zWFhqqLnbfJW4aQgdxu/lF6dws3E3GoeE
fgs6u/H/9EpV3koeACMbcs4VPsVGfF0obbjhNS7BsV6YyCGw8x1PDijqFMn3GlAW
f0FxM1Lp606K2QpuyECyVV3zNVx8tJNIGqI892jV55Sj5k5KZN2+Pz+J2xzk6UDk
wdvSMZAxAJwJEoZzypMNwWuEw9QgpY8MxSDmr1YO5p0o+DohSmdpXgVOq/Nb83Kj
2Y8W54DMlbj7zWETjq/sK7SCFU636NKOP0lpxvWpiUaATqUEoB/oy5KALcUHO0A2
lwh0e86MfcDJT3h8X8HzmN6ctm7iTQIwWmdKSq57d6epaXBAW/AzQtaPEh5Nm2SI
hrlo0IMP5wbDrLtVus7rzQmC2xV+o5uInF89S4njeTZiF3DMiuaRwZ9uXusWrK8I
0xygKAJxfTDvBmLH/xrwVuLAAEY3lPIx26Ykw0H1CqEvH+AYTfEBorKwh2BjZ5Xt
pzWaHd90/a/MMgVjk5XhnNS4AkruRg7K7BiqNRp9pJLX0rSJyfEPoZwYF8lDtpmZ
DW0NhFvlv3DpQPsMD5OkUlCrRoQRHiDGgpfH0rZMY7IJpPuDQgK+woKFLyXIoUad
78127zWtN0w44aopdCGt2TGz2D6s8dlPShXOc7iQ7AfAFKYK5dXInWBbSHROsYMC
pJdQEmhXT0sNXSAVaT/P7BTfG8dDicVeEDDUHA1kja8yz3Fopqy4kOXo0PH3mDFB
y4uWi4GJOtNtsXmxubcp5iG85/+ZfTzZ4OlHzz/DWdbYNXeJwEK96WAyGQcGNIiE
KczxAFkVpaPjkeN6eCsOrG1FMPzTewrVVggzDMyd0ycsDD6LxPJMOqBgm5oeOiFt
0eyAZEJiQtYgmkVe2h5H5Kx7VCHHPWvQZgWsS4BwAM8tfRJd8g4RtOQ8qDfqEqeY
oOBkvm6yVEtSXmiMZyB4RA2L3Q14yFSiBGizzO+Z6jIeibP8fEzyIUvluYM88Pt7
SSdVOqKaza6XjbV10c3+ExGsI4Vcodp7grVw89qziToYsK15nxXzRnIWur9fEXnW
Hkoazrtu/LID9602FEjDv5xbCGrcvbQzlf6VrR/+0wby3hVZkmk9XmZr61aHZDfc
Ewrqgynx+/xHNa8puPHzQao9ExBQpaieliAaj6wWPMxIlkVXKPW0UkJlcGgu6++/
RjWkmx5sfO+CT0wOVOHQNkZ+HQfqQX9Fhb07EiHg3KJuoie/09IFcMUtABJ0B5fj
Cl9reg9Sf2j+Iv33EnLrN2duWO21w2nWVfI9vmbPQLIG4rImCSW0pQ75XPgUgD2a
nIxYSwg5f0RmN/pwLHv8T23k9LZJaKRNmaAP6OsmiZd0vCdM+fqAzknK0bWX/SqQ
gy2PA8cKZ6oFPXz9w6/hkmHFL+8/NMndt7m3oDUWkZ67XvzihRwL9VdVgrBYQXRP
0AOj0WnOwe+KBBNXk0/SdJAZLTjjdw0w3TFMlgg3E3saDi5frnzj5CnvbElJ9cgn
w4YevUUlDumRgXtciDlTSUKdyQ42lYVtvhnYoQ29mPkPiMpVYW4bRjjftwvV56BK
36oLhGEazHOABdpjDhRSXfXz+CKxBP80JcyeDGVXXGb24IsfGGG53LW9l3mI7hJh
wi7KxHdW/7r+HHUUweoHVzDGgJiq4Foq1t76fF+czMAhZ8Q9kSm2iXAzcr7oFrgZ
mB/jm7OiF7XKY6BFCwix38Dpjvat1rCS4QvWszuW0B9CGsTYrjD5uJ5Xtg0Cbh1s
dyDdzmkYka+1S7TTpD608hOk2jHjH3o113BiVdoqSVLTvQUQ1bk3VXNaOsrQXMpO
k8nNDHfmalHuqdz6AHJ4dNQax/zN1aq2WSEc59eMwAVbWgOT8uam4an+bv/fnD9N
kZk/0bxcvyneYNKl1kSgqqKjimJb9vUwfpY58uSJIB+qkHETeJirLjhpLHbOoWVv
JYyOECsRudY2G9D4SWl5zh+uh+Xqksh9NAHOrgFvMupcd57+n5qFMhdob+DNAalY
5ZsJlXwPH0bOFtmV0NfGIS7+QP4ITucik4tVHMnE4LCuYVsXvb6Bl9zOnSoyoEXe
TXC3ATz8A7ffHi8P4RfTBupe499fe88zyN8tOmQotG9grcWGnQu2LOCqCJ76rL1Y
BBsgKLw0q5pVXWsY648vANCuQGXgOYLhwAsVrbPGpO1Tz/YPheOQNYVb4fqgrnxl
Uug4BqyT+zmuY6smWZX2A+7fqbZJWQ8tQ2CVPIx5PFMtVTImywL78AjjI4gYv12b
2jbENmQrnIYNZbH+yuby3yR+AnTphexwXTbgUVvYep3ezYYlABFmwbt9KKVwEJDc
v7o2E/cZO4t9+zqvNLSSzWwzCvtvuzWUQttuK7/x8W+9U8PEdl0d6BA6q7unvkaP
BHaJWoONbyycJYNNEmhPdrz7FmbW109IMsQ9ImgWORri7eAxCl9v5whrYqjQn5aK
GiflHBP+uDnrJ7fSnCkk9iSEYwaYvgIqAL1vA8afRPZKQ1XVp2iNtbKe5sDA9u/G
r+DgWaEfuwzB6A5Ub2nlpiS6egpJnUvQaPhOiaA9fcTY4nmkYnf2nnc+bQMdAX1/
cjZqOZ9WHzK1wtOP42W1AJbp9BzREJJwZgKQ+SRx6OVL875zCH5ttGLpHi8IiglG
0S+WbPetbSSSc3SiISQ31a4sLiK2CH5jYa0C4ziUgP127nOvkKjVC+lPy6DmJxJ7
zT86E1E1rhu4Uft2VTOsFzFzUbe31vonKzqyQV3eiT+meqN6Zb/S52YnnjR680L8
jfYA3/BTIPdoCywBcg6lkRa8S78LLvZk/SfDqIKE9Si0I9HwubGeXgzlhCq9/WYH
k6TtPDVWmH0uMQ2akBIAmF1AfbgQfpoCo0FN5lr+YVH6bHBiOzWjDpAscqaNVg2n
AXWNU78pfUWIQUzDoTJQe29F6G8BXEUR7OdAlf1cWnv04x1u4hpbvNTR+9OVK7Of
TU4YfbFe1xmgUoNarNX2SdkJZGfawabJjfc9nwqfrgUIPKA+uOiRuE+Qn6PQ0YR3
trGUvhZVsXMy61hYzQ4L1Ig823fvPfBu13ftJMJPgTCphv0E9Pyx8QdIa8kSQOqH
VbX4PhN75tmRaAY2Rb5mCjMKuHXe71EiodMhXkvShkfYwP28LkFvYAziUBFFCa8d
0K8Qha9YhlebhIiLpeYTDk56Vq/Tk8TeFZLscZ9jITWJHNyhlb9LdsDxZwAZU+xm
FnAxuQwag7w4kqCPNCzWER3p7FwFRuFRW4m/YL9gjBzDB851pHMs68qduLQ3P61f
8s9OkiHCHH9s+xhuD4IRDPl3Ez/OjPcQ8+xMJhM2W7rx+qhoUdmdC10pvil1TfGA
FYXFdC4IASDpGJg43SlYYspdp0G7Pv+lWX1UdsWqoK4iNCY3JfkrpHr+kMvIZCN8
ZsH9kNvbNnAxAoJwkSn6si83lQF2J7YwrGcrDDrtp+/IixP3lKHvObzv64gKu9jY
WNFHNxyj915PEjaqMXOYEOsvSkNSpbMnwsiuiK0tgL6pQwNagsn2IBYqGYN2Yf7r
PxqsSC/nTMiHo9/QAt5HlPaPkFtbvfBa4j09C3FkEbAUait+TibXqwAPZ8+OmiEN
3E5fikOBKUucaXqSEkZo5vX+ttMhRgwjG1P+2+dNUyOYPHmXvSvufpiBNiXdT7GF
L2Hx1TvaX8/9akjPwp35Uq+2dc145UsaBw9vVHIFT8l5CObHThjys8SboLu2CcIO
fATNTCLaBWd78jg/3kI7vhw1DfhCHdMz56RUmHVm3tffWvczC6AgJwepXi0gin56
g8ONW31Wol3qKQqGp6psbhE5FmRj5DhZQSmz653q1D8eog98UivvHcuwDuZG78WJ
CplH5/s8fsZnph+j7s++2otXSGv2WUQnkinAlJdxLd9LfNvdmiK6ZE/jyx0S4Trw
qIdyL8ew2Q1afjw9Mt8YPlr/WKqTrOh7zW6muUpcMGL5j+8BXbVh3hggp0ruOfaF
iiXUJWpWHL7kq9wm4F1oYgdiqsToxDD6X84kic8G3rsUroYsjZzfvi7PgJCpwf/p
1gNxCmdn6E1+PegANfmbl+3wLmzmU/97RzQnVEflrA+uT5u/Zfss/ejKJLUW+2ci
uCUBVpnFy2aUK6FTU77puK/6bfHrHaepzEiOgNmLeVYcgPWS9iRsnKCVJGNIo7kl
dMgZ/+JlncBAV6ciZF17DdWElxvKx5r6eQaIqea4bZsrnr0wKmpPoB7kLi7w78Ao
sMcZfP8J+pQZXko15kHh8N1uxSB6C9aCBO+Ofj/H/oP/jI0gnPqNwfIacXRUzFpW
m5H9uBBFMzJvd9naz6+ThSvDP2RV6ANvEumdCd3V8Ik6JTCnzn/XrVNYvwt/X2wg
UIFD5F9X128j6SGQXjwORrXYeASP90iy8Z9sXWDVk+mWlncRCJh/v2r/xvaXwvoj
AwpPZ9Dk3HOYUvdFLxjq2qlFZql8DL7w9Esw2FF3F0Tn9B/gFnIrO0yASslp0L/8
5PBgAyW4+/oP4/TKrOwUjMeCf2Z9omxr7Ny5HS2kTlbPGJAeggiV+I8lR+pj4cYe
v3q5WGb+bk/hCIYcp8UeZCqdZuoFDCRivW8y+OSlWiZ+AYb3wKciXqeEeJk59ht8
4cqhtLMFFExDMw5W/lgoKFcAEp3vzV9GOkr+0Hhjgq0S8i+yvbaRK43lYvE7rPeU
UMQXdIMk14c8Un/WTXpIZwH1e200Nsi1crDeVl148FIhdT1LcPm2amabT7jBdvop
AKBOZHCFgY90CnHa2QfrtlkGjeQ6VXKXi5aMXaqT6395xFab5YJh1tjH9CbSyqfv
Yko+T+jp4iURxHHjAkVQQ4nh5RChyaRW3RM7FkLtH1S7YKGuIsxLWDPUeCn1mmUK
i6mqFqJN0Mw1/YpaxhUJGxTVe2cCbVeS+swXn+nOz8PtQQ1dNwZajWWrmJoyPnF7
cdKF6fxEblZM/3AVzhstTyFEsoL1QoDNaKjjWIxKzEKqK0qCygrcz+TVGU4MGbsT
Zs+lMVf/MVKZHfgjIgSZjMl/uYb4b5buczSJWVOk8b6gV48ag1WKcyXD3yxrsfG0
fF02vos0Xf2kXuCgLulMFKkXmaUbjxbg98/1zzsmrwiqn8OhAdaMTcjLMLVu9gRg
JGNbsKNXkPuNblJ4kVK4I55nqO8T8AHWQkNxASmyMoJgAHlb2zRln/K9nC7E3lxb
E15l3CZzeWQzIQxBBSt3bcpmvMcANkTc8BXAPULJq/dFNfVEPDG1dEsqDHD/dI0P
r6UO3rTjbEFmcakEkO7hRjZ6a4HjMDLtjoPypReeo0XMmFdh6FRPuF9APWTelnqq
M8zDMas+2LDrkUkyeLsaIifkS7/m/sQ4zkBcP5qlLNnBKz4IhqfdO7jksxqPFP6r
VJyEoS0VhCEXAtWUtONyGopo8bTR1uR0XAD8iWFXScpSIeTxnAs2v0S9BXvR2s3W
6vJd3BFkLH6bIHSyHE8c0gQZody9XO5aG3Krdf18+NWed5KPdT/zMTy+m1sJh60/
6y01iCKZxm4qDKZYhb3xNe20pomFYu5NiKdceDflPkH2nRuauk1rfIuSS+eS9NrQ
k/e/mamhhJkGMUtyBH1Tg5kJ2hst7T+1QE9M328tYVzmlGnX2bro06cSuPf8idfb
Y2c/OWB0fE/7l1vqn2bPx7TC5P7qVzdbHq2j6de1C46xXE6w6m9jSRkfZ4kExeAc
R6YjFYPMJ18pxTfne4rT9co1E4QBdB9E+Z9J/Uor5kVkyUMf5TS9WqRtMsFgLXzf
HAwzPP3+NkIIIDguKF07egotHXr47iwyn4qS67hR6i2NXuViOsn7+VdkTiSfL41L
AXfSvDZRmHbpmRgq/fQG1v/FinQ4mSappqDTzWUpAztTbRRXE19hc+oJgD3DZBGI
LNRa/vhpSM1g92g4RetB/UOmi6kM2XWd027Q0jT5kwqorrN3gDFYXk25+KZJMlji
gRETn9VTjSy3PLjjvLsbGZtz9FDGu/ayiW2KPMhurHEMrDj8EX41ylshZkaQ2eLU
9VJMcjCzkuUQKmuQv7pkNLAtzXYE5tkVQp3x/u+OEyEXjXxCVs8UFoN2dNQsqqPc
X+OgPzRDZGRQPawGoRjp8Q0wgfyBW05ICV/UHpPgrTOFXtlcOUfeN+oEy6dwcqio
jhh4S1eOaGc2yBdN8f3T0bn9NjmTafAHRsmz4PoysQHayNMhb0MgSZFu7aIDnn5x
P1TTulCmU+P/QYXEGCk8O+c3dZviqp1FUVYma9WritXOH7nTZrAQ271/TF1xycnf
azkwfOsxy+r6HHfCo5ShJXTXp+P1gk0gWXTWeJGk37qTsMZMSwKJ2dgKPHAQ+3Rg
E5q1tEY0KBNuhMCyKYRQEiMDQJs94Y97B0iAai04nHY9rQPpSeBoyo93tE/THCga
O9KEemvZjrkJOGtviyq6j6kaL7SRCM4L1eehkKvu46bE8W4AFCf6OBfoZjV5unXU
95adJw6F/ghxMesCRTMBYB/NN07kb0HeYrAJxu0kcCHGXjDhUmeNpjUTy6uLeCQQ
NjKZuervfKcvpVmkVJRPqWF8VKcdg3uJWrjqle4L7gdnDGAZJ570Nhumip+yZ/Mp
CNTYnVv8Bz/hO8Maxmc/etKJ/NKPMd48txXSGk6s/xmWqtKsO2/BQ/3iZ46JLEvz
GUFgRV/GiGP6zN/ZyfedNOAt+acO69KzalCRFEQf82s/FkZ6GDr8XLJU690TRjiL
ATIGv/iWJehjfXjgMgwflk1eXvOqV1d1f5QdL+gApnBq41S8Fttya5weW5pfnJuz
XXQUX1cbLO5MjpvXN6kGLZdJIPP2ktuVUv+WuJ2Y2VBufhLIFRtgn0dyfUPA5gvv
v20bn4t8JhG0HexslfODq6OOvfzLZiVUGLyFO4F1LGKQRSzJpatDW4IytTQmNe3x
Kw6AiaOSbdIDUPw04lgxKfNraHiTAVFNuvvUqOGS9s3j93NVB1sjtTYpeyJNrpOH
WZ618Si/OlrIJJTeRer1jTZr2VvURxeukd/bhf3tqjZTs34Dbf/ZD+7AUUAFNCxM
Dq+OQdvPa3j6zWcRbXyqxDfxg4SsF1/lXxA/FVQAsBFInbLA7G5WlzK2+K6X244H
tGtHScepbX1MG5MaScz1gHmD2Q09py473hUxE9C0H2+9TaQWXeFnp1bS51ehkgmE
YAfSTpamKyDGOeITBBpp/VYaPi0hfufN/KCY/kUlEdi4AMjd+gi/hC24ZmKF6CVL
9UEgodBSEdhNhw2IfQ5k/xPMco0iwTeoYpcx/yYb1rUpGmx6F1frxWmOXhhJHTLW
TiPjJaNVey2TiPRJ+MygZkMEgk7Dq0n7wn9P/27+2oiXBr9HTrUuyW97v2XfTOVv
c88EGn0unOHJ4MqDGF0mr2eern9fXOmpfSHPFoDm1DYRRehondzK0ejdVbCPIcyk
BzoKn0spo1ay9H47GQbMu96pfB4D+IV5zZFeUlpE39XSlTDSOd6EDLNN1b2LAbyz
jl5V7ZQLb1QD7KSfs9MnpvT6wjggHzbdH6gKjv4iTR0LqpMXq93t9UsCPURutFg7
hrNwGfAPLULEUYKZrMKNSH7E8a5W4EYaklhpH+p9KAVgd1IqJG9OYdEKOfSGT27b
aboqvmBBkHc1JG1jIeDTcp9wZYlbnT1VNTSTI5BySkpceIzMU5dKMs+fNUe6cKwo
NKLe9OrTDh3Sj+yvuiF5/SeVDtT1Tuy7HL+vt5TZFndlokc3oVwM/4wq/JlCJPtt
WzCGY7J6PFj63Ts+Woj/PYfa9WIWuOWgft4muypwCW72IurTD+JFTtLR0ghDH/ch
yuMQ0ZkeEnrWHPCFK5kHaDAk5/E6Rf4qSpP3QuPaTeDrkY1InTNFlGWIPWHmKD4l
EovDFkWkbQMxVVqNIKqvzGkBUvCJZGoM3lZFxKycwL3BywPLUmlyG5ZVabWshclP
YFeuGCCD9ebo6c0b4YFUrmFCzOnJUWWFUkxuqQnMN59QsBwJk/ka7g0lhtRgc/HL
FD+td9JCsxXEepBYgpb+BldFDDiAAzdPKErSF75x75Q2z9RTKVEEJkw6P65M6fDj
CjbJe5bFrNbVLjm8qOYaaxKY8OuxPzXTxMlAfNFOwq3VhUp7LChsX8DEMBSsr9OA
ZnzdGmYb+Cvc8QbGeWVNPC8ZVDaRXdqrPLhxrvXtOUKtIN8cAPidxVzzhXpuxYFE
MD7lXQDWi/Av+HgjsoPLplBmw/7DU3LuIPO//fPlab3OOC24n4r72u33t6NV/Z9R
rs1D+bEf/CB6YThpz4hT3MarGB2L44Cnm4Szzx2bjgVqAMNHvrHMOD9qyPPjUsDG
XaJETciH7XudrVa7X4IEsf01Bj/qK2mQysTJpL/qg3ONrE8toSdRdXukSAkLPbeP
6SqEH4nIQM5Q4tEnN8zUEPlxuzf4HijD9dyO8BtRHOpbvSqmTGkipLcbdqlbYerK
pCqaEfJTftnyVduC2gchTpDl9o5VxIxpHPRqPTd8pjlrrgtmlUxkmcWlmpI7T3Zn
uBMBZIKhfRyqC7PhAjlx2QGm9OQhnQmXodHdp8QPg9ZGdonRNa2OSM6tbD88Mcd5
dY9lStZa1GFiWbopzrguK+nWdHM2IcPLQwmdEaLJsNMUUnvwP+YXr6QeUHBAUsQ+
q65Ncfo5YZGOp/qNV3rEfeaFZsK3oBISS1gVVTt3oHWb88eoPUNymE+6BKE6km29
W1jsJdlPlplG6LU5greFwKRwDlr7WFyyWUyX1X7AzNu/iaLUrVJe6Q3o9F0B3gxg
gsjv5pgbefMwCeOTR/aJuuXIr7Bx9Yfl65XxgMeloU3DXbIn13vs3E/6EPO7FYLp
2PwWulpwnoPgAuN5pwbu1UW9Xm2QOhB869ajC4OWpr/DE/SIxNRK+XOt1vs2UNVn
4aYFG0IoW68K7Lpcz4+9P45VucI1mvupq2WVFFZWY9uVAyqSYoKEUrK0+gXCQsG0
GE8ZMvUBBMdOYHcEFHxhuXbcA2NTCw53SPytVnDuzKVOoEuOI/upYRkFSt6pI7ag
PKLdBPLoH+4nwcMMsKivyWNRhtCLsOJdH/ARag9HGaJJ9RVXKBcP9FLjbQuyd2Un
U5PIgd/YKRlQl1DsOFQQ/EvaamVdt17JBS3ugruqqNrZ05S+lMwBrLmQy2Uq3UTt
ezRPYe15BjmaxRlfpFugK1qpicE/Uge9F+24nhxwiJ/FAcztekJ3hPxgDSA4u6IP
Mre1wF4yC86f9di4ojAiU8rTQqmocLtZQKZo08IN15q1QOJ27H0IQ/HymBP4ueL7
xrloZmosozx/kw1s2IOo30FQwAYLcJL/B2sbsNcmL5Mye4HA35aT+aFXTZJ9xNri
6lPkSr0BhSWtnHcdGY3EsLynGDAx8iIeCHOglITtQa5GjwBQt3FL62pOEnewwjyx
9l31FyGfvpLmJ+WDI8S/WxULkS42xKuqq/OOs8GZ0EwBElpjunw1T7JnGoX2czp0
KBlEDbNwOuQAu6iefLaBgxgTvty4CwB2mY/qJ49OOFCytJHvaMVC9e9XyZX6BkkE
En+AgLA8lcFVd9P9MlIAPjwph/C/SDHtCuzU6yZaxsxp+38ur+hGsj6qfK/84/Ht
5vXK/6YDKgSQj4vZ5rx5HUbTnaOVSB8QB9Bd1aqkvoyzkHkv9br+4zUSe1GClGpc
Jghv1zeftYHl9JIND4ILrYNrxEOhn2eyB6cVT9BdmPheb+mQd2qTSFzq+2H1kqGf
u/LjoiZbEO3Fufe31beN3w2ZGmqxI6yMr3mujIsD5h3+zVxdn7YFV1GoLEAWba+a
yz2K01fZdfIaWJuasOuVEsZ/kKUuLvJrnl66LLKg9c+jvpfyWQ5M14O6qBCwh1VZ
Z67Cps7qzZjOuvLW7xOyAjwCjSvND4EI/Z5RKMe8dRj4XNQrpsFshLaTHiLxH3wG
Oc4Z8e97XkqE8aSTuVgJ6P86CuVME8b+ogz1z04DYG1X1U08eF1BCpY8WNUPX9Bh
m1oLgoR4q20Ti5y+99wsTebC3gVAlUa8OYRlfJLmKQnODfNj5hvKpia9vcgwYufe
tD7VgTz+2jRAE6NRg2IqT/Iay+qiA/dBNzMi8y8yDUvPm3ER11rebjE7pxqURqj9
4WQocJiNhE/1GXBf+BM9DWTtIU8iwLfiY3wlJOzZ2yV1dnGIQTPW5uLL5xTGq45X
LivcZwMtKu2IDpEToHkFs6R/RtcMG8ZVrtE9Hwhr51+JkotfbPNPqRooTyExE2fA
nsHjm2QxfGNu0B/86sGCUvdKHfkDzD2imkWtPiWEqK9ftYFJxJUTEIvvk4d2+mYA
0ciIix5MOUaTqUMmdLpgjVDHlxJ43xCHhoNzAxlB7jE/z/UqlBDZDAnZZaXhA4CY
LtHbVxzeNfpYGT7sdrvauxj7AYFbnRZewO//41Ku+KNCKSlWYNo+fsd/MaOz5XAk
uQY+aD4Nxzr3WjSCdi/hsF+2SUwChuai4gbBdCt6JrE9JOE5hGMUSKXaVth6dg60
pszZ/dxC18Q1/i1k7en45VSN2SqvtY1tKFQk+9DsFq61BUw5S2RSuqNNr12X8TJy
4lG64ddnSCvxHXm3rEWakZmn6umXWaiYfMR0rNtj/z1ZfvjUKvmxuPbISEaCx9h8
vyd1Ovxe1DLhfCRSasrt/eT4pas7WlM01E8Phx4OUXRfX/nMXSJwQ1/fYuc4zA3r
u8KsZRY5k6tUnMCzzReF3WsBZBc+H3icDaIHaM2OhVUo1KP2JL51ZdGl4yRcKyq+
9Xq3iNNtv7l1lDUU38212U5JS+Cf5YFd81RvbGG+0bF5WukIMQrzMCqXe+reuMzV
cA95Cap5lNwRfopxh6oQTN+gbkjfZmRedc0fmdQGduA+VDnU43dTBJeb1/c23Adp
iEJqH+in46m9ZV0apmwnV3MybqByiZKovTbCGJoocpoXZhPJlOAHH1oNmewZK77f
jsSgN8a3HGX8x8ihCPBtQI2StLrLjrOswO1ehOM4woKDoxlwJHO8puoSsmJNaIo3
CwJh2bIXsPUYam8HNvi0jElKf6ByTKw8sDRe/QuD1489QdDa+mbtXShCgxrqU8x6
m3F7zSDfpyw2CGp2RE10YzJ2lxLiWFnNi7kfeJcZ5VyYRRxJO12I6y9Fg4Rpwot7
yzH4FEG4D+naAYWMgIifJBRGZTr5h0j5wvRqZqHye2ZyM7aDV+vnX09wzHKCTwvZ
+rjCRcj3BGgofWareegKfpx7Ww2+aMpsLUtPplQGuWmJPHV5U1iNRDOgKoFbqkcJ
iBQlWlHbK+/sNqNBolQjaa/oi68cRs/YBAceWHKg+1gZNK9hpr+2JzkHoe2S4L7z
VX2kd7gScviCT5EqMsa8SJyNHZJnu8ov1DWccBj9EDPFMd406Z78UTzL3iMb6MVm
Uz11B2jBtgmI55l6YG0gIjlbYbC+9dlY2TE8S6B6xnYxmF0l1i/vny0gjdjSKkMa
zAyuhrwtzVyaCplcU5BMZMlxuctrFiV92PrbFNuG50arAckrdFuv6+b5K9oR1u/P
Mt5otkp3EXYui+qmzc7DlQX/GN44WsbH2hKlvQipavxYaqK38M9vro0L3hdE3cDj
u+P09b2B7AocKzHHpmjVfZrP8Mmf9uSRvpJLwYp31k+n2iXqdwVtsVDSMToF8Ear
Ho7jzwzcB3L0zaWkHxejkrCl7i8cvkzsvvJprHUxA6xZ+/BOpgFdZKN8DeaxTk6h
Zbv93gP5S7fmqB3E8R3GCyPKg5xitJi0rKlITy7HTdcgBYZ7jtofhWPie9nfx5xy
xDifKMPHMrW0D2suNgBM0eY69Tu1KmgkaIGaXi7MI3TLRDUThuid3vyoGEhjotmk
NbC8AnPOAa+7SiijKBSfkvOYDjeAEXKRpzCkR//ZqItGrtm1j6hpp5AycVqQhazc
6gn66hAouVL0mpvxaT/HwtUBXTmqarxoXdcw5oOFId5qEQtqE28TBOjzplm4NBBD
aUEQwiJ0nERqslTqcR7hCcqiGVXtDAl1If3vecOpfOxwyQ30NhtPbeiqtzHseGZA
KriajvRWkiuObcEvoIKhgucH+KBcoP7cl0OH5+j+2kBuQXxAUv0jetMUiOu9AK+S
O+mQ5rdw42cnI55iLUm2v9LZsWYQMsD3vd01isDb7ceedkgQJoF+5EiYm8f/BaZw
00IhvfCxa68Hoi3YGLTKJpKN+ddjlvVcFU3REjVNP3sZIggPNXxZbDqKKI/6NTud
DpEgxxIVY1iYrc7Iql0wrMq4oHgT8Jl0b/Xyx6JaSqYIDqPXuS6AgPcSjILKSDLu
zTrvlRgXBeysGl3fG6m16aJrd0FTwQ3rukJNf/YLw1Qw6waK5YzTD9p9P86zdvl7
HShBuSyGgO74KSki6QnB+fe4Df5jSBxO9+rKigIDHUpkDlksKDtDZnYnB+IF9mK2
OKy+Vdmg4Mbu25x+uxpPvrIIy73XYbedQ3IBVgEb+rvKXatdRps5+06jLFIWLZHU
TQa/6w+tnPIM6JttvBOajrpjQcUYhNsAlKoowD0My2rfzm0qdQifINnItQsBgZMy
h1WulZWiMNN4jp+LLHdnrBKwb62oZCd08bleMDaa6+Vxo5944EAYMqyITARZSPjq
fXiCZs+79S5pxcvfeP+XHYPS9whqjw04CjY8V3oVxH3wskEnt5x1m8Syvgz1vmkz
k2dxcBtf4th8dDvPmYCyt4ylofY2/eYTUvFetR93EluQzt6ZdL4LcIQfU9tSGM5F
lNIoAYjGBmv2S9cDyo+5r0IMPrYyRYcsx0kGYrS/vM5KdMPa2awytYU1ud1toLSm
Q2sxpjYZTNsuMPl2iScdZfFe/Qe5UkwAN58oaMpHGZWJeXBH1gxNPiy9p4ucZjRL
KhW34GT1ZkTBspqseMACzQirBj0cfFSKqWHEIH+w9uQq3r8lvTQuC39cBpsZukn+
XQWvE6xk/hJ610A0s89fvZEYNvfKfoOYNMgAsCmtgJkqbkrUae3U+QcX53+2U6Wt
OzVEiccB/5gUPP1R16AG02AOR52uKJLYgY8OKe349UwvVl/wDHDmNa9zyC7J+tHx
aP9Oz9CeNwWbJOkK9kO7KAqsKmnxqXOf6EqlV3EE/3AVCHPt60fpIts7QaXv5guH
Lz8+2N+1l5rq/FVujDMkbIV5TgyeGj2YQx1m1xeCSr1zY5OuBhaOU2ZyRt0ZyaiG
wKs4//rtz+hKygDQKgykr25ku5382Ppv6oIR0Va/qeXwctG67yzbzVOQWIpZI5mJ
1ImUSJDNYhSeyXgHOXzi8Po2cudR8SOMtoji6HNpiJlmXB2DSNbd1+mCpk1kBt4E
FwVQq8fwfbzW64aZAJdJmV0TJGlA3h+DTV2lXiLaNl37q/oTWGLIVZ45+kFfUL0N
igl11/EyWSjXAQ0uFc6AlyLV1YmISs+nl2jqc473oIF6GnGqFcbNyv+aSq00KqJW
Dj2nQq/jidyHZ7wys34WD8vJB0I8vjKsAbP+LQv2fiEcrrzWJyzk5/wSe8TrjSW0
24SWOXNLYBYLW+XuH1idyagsfmqRGI8EjujMfpgBXmT2Am9q9JjJSdqtvFrb7suW
L2IarIdNqZtUtTBiDi98BzvSs45RG4p8qkPdEfatf6EG6B2uVOJivIzPWsxuL15n
8eCJFkgN6DtPzuds3FNpC0l37xZjp2fzyAsxrxQDi3MyEpBS8Ci9gbqL74zuKq4t
nTJv7/K1PKvSOyiMS0MfAgH1kKBPpfewaKnT2r1w7nseUEQI4UQhOGlcPhgL+ezF
LDmehZoqtoXTGaidesH2x5rhzWCZqxvP8G9jcSesPmQA81GleDtVZbEirkda1Yc9
wwssrRTUS9XZEF1JpYf9E/azwbgJxloM/tH0O6QcY8KlbFvLptiOZbi0qInjWSAv
RzQms7ia3fEKRnUtOmIp0vVY/CO+0QXuiu8nnEf61Ugt2nqNGKagjlDc1P54ZP7A
WhSt405ZaNZ9lHRxSlohCPe0l+85xkspWbdmSdtNBr7jBGwULPJvRNvCt2qXCjE2
KGDePGjlAQCWSzldXlSUTe/c6Tym6y+GNmvD7e1Q16z1bZ6hdJ8abHQ7E/aQSnaz
h+BMfd7QgVqdcPtGFLtODELlOprgcfCJ4f2cYVaTfK/fK6+ghh9hhG3d2gO/REW7
VDq9HpCIGjGYmEEjLhhRrNhyJOf/KnYAWrh/LJXoxNICFGtibSRi2kPxox2rUj99
JuWKlAG2aAtbjq8zGcadJZMzbrrZ1oOKJ5lGfkEbKEmajGT7USE8rEdw2cRgvM/K
j1Mlwni1RVhF8StGbcrPHoyWl9WMQQEAPAqP8SJL7OIVmukNxe8h+Mo+n/4/eXQk
KVVc1EUcdX3h2F36QHwdkIxk42MhOm1r6FP9/Z5UpnT9GKHB/bIsOq5YTxPPqo9G
BNnZJNUBO9hnqk7rtLFEFEfnNEowiyW4KxTXhH/ZK2kz5rTI8IFRTNMmSUE2CQX0
+hJ87VHsKPSnySy/EnK/UiBJe2ZdS/OuFY3s6JKUCZ6+5uWMeNow6N4qKhWCGfmA
FYQzwLjL3IQnbWCAsbAN84z89YF272H1PFhtVTh/7HQ+9T/UTmZF82A+0cWXmE1D
bHeSBB0A2Jy/9esvM02Ilt+E73B8bP1J5yMoSZ7Rk5stzmp0TmHa5KGJPRltjwUF
uVA7YKCOCpwGzNihls2oanBHzURYHdRPZGb82rK5l/EzAfrXhbv0eARxCk6HHl0z
NoVcqoof0+uo9HdaNz35zjBnngDyWVznStDO1H7O8NBJmQTav2rIT/s9H0racEFZ
31hYAveIWVsVvd2lkQgODCzW6K5oz/RqFvPaeJUjIoLo/WslfFGS5MjFykoKoA3d
uFJvStOn0r3ANIgoaBYIzrEvALmm6UjwgOWvIH1pBGpCbfz6lefSyg/9L/g7O6B7
Wjlkdrcq7NutD40fIlDD3fuO13SjOCYBLYM1uWey9kax5zlkuBuBeoXD5bg3E7+0
qxA/cxRFky+r6ojRd41PVFLJQfotKnq7/u/sgu6GYf9cjsStgFeXNzdwQ4M+pwhE
cpxgKx2nsIesZYkRe0jzmySN3v6ZY6vd+8YXB0k7dKkNMkLUG9HsHhbIyUwtIpXc
qnlB9DNocYeIMsSWZZ/jNz0OwT8d73vp8usf/EkbeLXdiTvQGgnsVMBWL0+0aDtj
NUViZRn932qe5bppqAfbigosqknpECprA3zzDLqSUP6SYfR8SGvTT1ifgv8MAvMq
WqYdTvPhOdYbl5LmH5hkeYQySCm7WG/mvz8UQAgL/BJ3cxJ2CVwhtahOxHoRX3y7
Np/jqYhUxeFEH8M0o0arJpGGMCNI67qi2CgIykmJXfEZydOnDWrp3+jUcdlaKSN3
ccZ2zHaMRmKhFjqOO2NqCyXmhCGnL92IooMoC0BNL82D/ZCokpriKo8oWUHoYit9
6FsRGTS1EQnz1QA9BF0SWDCjak6xEaKVtNLJ5nbyHB4mhw+qvBJ8+E5nzOIKNzkd
V5fra5SeFmlCZHve0IWob5uP2gquxuOz+MV8ydayX/c4TSnAp0tLxZu2dZrjtiGT
czUc8WKM386PCK43ZwZfbk3+ktfhcKf4lcxtr3P+Dwrz6xpfrXCoY7As0jtOH8zN
O/jQgfdPANiclTUU9QyH5+pyKJ/Xf457CgjTk34d3yjZOQRcwlJTqD/tFErv+umf
1G9YXIvmBK/DQM5SStyeFjsUcRO5ZBn4yGuCC6pq/v6S/uaAvNi2CIxU6GhJ5V97
N/N5blO3RDVLciK1zmmpYxJVtitZ0VrGgCNuflJJGD+k5XSov76oUohkzOCmcXDm
zHeZuoHrDMu15qcKd1tUTrjMjtdkMA6M7Vvc4o47j7qUNxZQAG7Icede4lUGDUwL
fW2gRANIs1SucHQa3zKYaV09gelWFNPrRf2ijOB7p34/QnXsAUw/7HoiXxFpzDTH
7T7e2JtapBTQHih2HtEU0e5mVKeg+a3jZ8P3kIWgFXzqWImkQRuHIByBBtJC+XlK
XqwvgttwyUiL0wSYZKY6ypeyqGGXq2jFOEYAkW7ZTX7rQ5cemTnShjg+ep/fmS/A
EslDaT9SN7yYJFAkDy1ne9tM5dd0Xy6tD1/AEo1g5sQ7DaOBk6Z/ag9iq8ZHlBks
7EQuqfafnNs53yHhId4KBjvPZdsF15jodeAxVOkNbOzlRxxmSEbaYeUtR3WBLPdN
CTs2fqogKb3CK6duAyDOGE9UAafgw6S+Nzx/KxAgaNzlBWIj1To4CXM10fCfyqev
M4O2pFL8dvS9Cpz/iG1ABx7EYAtvbgzMbxDxRRKjjH5H13FFShM1sAkVniVYGeSv
2YfWgETsdTGtnQdp5bw7wVl/+ShP1TUPnZUZSA9hcD2rQsvOaumvPXaTmx5rwWKi
o1QbA6KiPwBei5anqSMrnyvOiE36ltPoXMLTnSmKE4JBioDwRFkgnpbXMLfd+qdP
rqk2ic9ZLMrdYxK2cDccFgAArVjs690vnwm6wOAb1LNBVq+SqAXsHQGtJMvxkngM
ICFhatDHlZ8bc5goZKZ6KN9FVZYgY+gORYQP3fue+rIeU5EwnnAM3pYjxVFoJAFI
58/4YxvfayzNaeO/FHiB+faqzAcaVwO7SdB5RLFfM6ogDEgeSfLa6v1wAT05K7YW
HkdoJR3eEdvMFaqiGOeKNP6GXeHQ/HbpHUQnqNm6qU4fZ1PIieYEwTyA0qnNWUeL
NVcT76kvnor2y7/VfXFrkhLRNqwNvyix5RRPl1gEpngXlmn1Cz1jVeeImFDqJ9su
Wqp7WBQPN2WXLETnGCggDnDjSU9X/ISXrskV+ACMbsy8YQOatp4q75uoVIhNgs+l
E3WpV5Pifc8CMCoro077sBLoagCJo3clA9EC5AdOv19RwaDwoUrxNsm3LsrKV9dj
Dqvq4csLw36aseXbiLOrAP4RZxh7a07qv82ILz52vGYW1NHCwa1MoKe2GFBL+LuS
hnIxKpyQgXQ8YYok56MpvtBiYfKMKyL3Gw2qfUSbnz5Lmij610o1QtCaieVN5dbK
CDbOJeTkdH57V9Amamd1Jq5sbhGXBWQU7WxnWdr9xComu05HkORtrpiTX91J079T
ErT6ZJc1Ukew5SwVpQexhNuc65ypgh++palqVc/D9fNq2ehyp9j+pZxg/G//hwTk
YA7Yygdg7XKdFbIfCWmLUKSqLe6sLv8+zTUG1kh1hIgOZRsQKKm6wsOj4VljFHUZ
uHUL6PidMLDyJiqXCldmMQuXuaSskOQRIV1LS4MU7puUJNLm0DA+eQZxCL/tDGrR
BAvqU/mHgwbp/m+Bppy5BG+CZV5ps8NtWomdeRf078ORBbBP8a3YNRHjSRqLFQyY
Dt3RCR/kxpv2PQiJ3WTlUiuh4jNY09Quvzb0QOAQJXDcB72R64X9d4cVw779OL0W
KVXLooL8nuPI13ty59DKuOcOgz0cq7jQsTN6N3s/gd32fvmaP+jiBf8fGWYKoaJw
LeQB04x/qocU+QfoujS78VeQm0sbSxPaZxXfsw4ccRZAzu61opcyPrO8qQwWnmcI
ErvDKSTNTF6vbjEZr4CsAfrTvyxWwIaxH33bMMMXNea9WmXWeRthW/bHohekuI0D
xiQ8Hwr8sQYydR0y9LsEwO2eLQLOcA6XCuUf63VK81sYdBNp89EhVVg6oA3ZyQN2
AYAFDY5bo74LNkJRxmMIsYQocJTVrhGet/p+Pm84SWF/IEUQ2gONlOMaQttc/y+R
Mrkxqj+vURxcBKvTC7Jk8oooOxbZHLEh0g6DLjjN++ezEotU0x+gY31S/EBY4NoV
TVxQGLmeiOff+214dGGwigWXPBh/BQLlExyZE6IOyBT6bogGj4Xe5lnK7TJ7TbI7
0yZ5QpOWqDMic5LPVq0FYgXtpgqqNkgv64IBWsXcYkUozGFERrK2yWC/Qr/yY6np
BTPb2iz0FytooI4rXNRL3v5Xo5FrIvdSASSPOm/VYRjzAtg0DKPY4gSuQUvc/jQc
LB4XNhpOzuDHM/10pjF8P6vJmpE17pM9y1A9QyYnGHAq5d4HDzyF3ECHEoKR4yR6
P2yeWOJ3ryWY0X0F69Bj0cF6zxV7D+FhqMW8ecSP17/94e1y+yJDzD7mv8I23bHd
eP3cKtdUcW9p9titn8D4BIQDRqmwCLelf0Q/XFDCl5Bj5NaD42+Y7rt7H1XY45Z/
8D4J4LqVBKpB46o+GF/FZNQviSoAKlT/xSOYCVHyj6s5AfolcjgryFKUHw9n62TD
OHSHvtRhcRuGlY7enAHudzgRv79EIQl889h12onPOWJk+xPXSmEwsUD/7kFJACoz
bfrUYHNvDBk7dzZl9dfipSsi1DOTvbw0N46Yx2Aax3mP0jKQtPmVuq6ZVITjQXTd
tM/v4LYjUU15oczx3/M98pzyJQuhyhGB1CqDapSJ5NVbHEIFVQw8sXaSmALoKzfv
w7o3vTYDd3eKugCKy0SeH1eeeFMOsGcc6ono/rSuIYB1NoIWiHM4z1EnWsobf5A6
g0sXg3IQonqImNT4YBn5XKfPAmgVSFBJm8FCERUVWbQeMKfpSPaEW+E6MRpJIYcd
E1bFz31F8eak/AOAZcWf27NZfoG7W3cBSMaZWqa0AjsoU9/ndalLuN6USWGAUoYx
7fnly6Ja0jzYoE67O5nOilMCZXa+CpiqxB+PKGKXmqWgSyG3EWjj3eN2QGtNhXsE
8rGpwnaBW0EvWKTMnf+gFao+sWkMoiPwinGSxCBfU8TOG7iNsgHpgjYglcsc/jgS
rcBPLsL8mfwvBpn6qyqtCNjNX+zoWtsClk/8VzunUBkezqXbXYc5jOrJdH3mSmqz
SqVKXNQVwKmUwHiqan4toq8AYlIz7zTtRoviVcpR5De9V0Et9xcHJyv5NWF9vSXo
b9iXDyNcLiA8b7eE6AbqnJdqdM83P+yWQ721smuBIkUiuD5K6gBQcBISWgjqHOTr
UMw4Jjdk+NvgU5zp2kLVM7td1iOPpwhxuyvAtjzLlYGPqqLkCIn7tmd99Sqx4o94
6l1yTi1eqlXkxmYVaRkAACjD/o8wH5cFqXC24NQyVftyPArdkI8L8UB4bcUtvxSD
4pIN/DrLWXS0+VHxd7YVx3A1MvWZHYUvT+FZsqAxhwXcrh0WJMTsA/MfOqfkrc2j
7SFx6g7jvhEwUc7k3Z/ACM0RJRkvLAsrHaVGhWrh+FjX3O3Ffbz+0IrGZSM1yqq7
EPiThInsQAybljepJ/5+jGmyk+S4PIbzQ0elPKfRSl3bdBsV5c1h1YbMXWpmFAfc
sB21hNYFXxIwSE780JRT64d57hi+SGTEqKuB8QJHez+EE2BFSHaI+PVFNLYY2476
EGryPe7Z4MXcs8jZ5KLOMPpq0PQv2V7LmjHOUuM86nXDnCzltN1Z/ZEwztSpu89i
pXDXunJkuGkZ+yG2zydbT8F7WPrm2zd9NXGS8a1vXDzp28VD4zkx0sJwznkyNmHY
2MAfVBJqAu4+RjVUA5kSkIkKzfkwVAlan6m06VCemz4+jITKD2Qtb1eZGblvEiaK
XqH30Omtr60l5QZ316L+2Wmg3D4ZKO3XK8+McOoTTlVbfIX/871IOpS1bkammTbF
zHQxE8sMT0YEbq0zwdD9UIG27GxQW8Khx+9opU3DV/wwQgPfexB7PvsJ46jX+uav
I83nDobzs1fqi/bgDV6cuaGIMzvKfCVEhpcnEwE8cWXLTrqqIlCXYpLjfX9+iK8M
WEmMJFMmjRIyT4S53gPe6jpj3OMoAdwHVVIrDnKKtOxjrEJrVjDcQVl1OQppkAUk
dpy+pYSmykyS7BVrKd2pFfm3CtEqxOylXje62OJSsCgmflPc5Q/AnqhWXrfkQ/A5
jXnRE/9VRM5i3qwdmlS1OOUEbUA0J2rrFmIJrKZGfgiaYFJxmAw1aqW1LZLPFwsL
ywdpuVOIUVU9031bdimjYJBOpF5OV/sfXlYa26ekg1GOhgO21sdNqJzpKGQGjCiF
rZjR6x2c0G1ON0MnA6DXBfj8K9wtpTeUVHbOFufIr3BH1V75x1PK6XkOeo9pNIi6
woCGFkq806F5PdWKiU4GaKWJL7Dp1poraRY5OiD7rzx5yiwHB9T+ivdsvzQZ5+EV
0JAAEDNboGYMIa69NnpnNoIUEmDqVb9LaEAxDCSLe+66kIUULGdR9c8TQRw+48qJ
7wXg8Fx7Z31TVHtuEI1Gnlijh85NKXOmCyCG+7azE85SdP1zQAUX/Z8kF7ZM0VE+
MvhS/5XfadorO/qL9SVZjUhgHA0D61z0Y52VNxcV4WBsSfQccu9UwM7e5sFp2Qgv
ZsPckAXOIaZTihAWb557T5O5G7hxYVgazmg3+zrGxXSA9mZKzwB+Sx3fJcUAq4Fq
Hxo3RwpC+kGgfL091e+ZIIuo99PDYtBHeIF2dsPwTN5vQUVtRSt+wKoWDkCUwRgQ
Hu527cw7ZPvmJhRP4u3ZCqOd+eue8D4rrH4DG13FqiJ1QdSWM1EJpu4Dxbajl8bM
Q8ESa3bT6xYACybDhyGihqlYz9qatxMKv9cfzhlR4DRRIpLOg9fEGvYux2RkcyfW
oKltszDv8x38XbnfviJfNYNRBHyNhJJwXQgP+TbuvmxIjHM6ZA5UZZHDxy720B+T
yd+As4hqsq4gaBYzJqQcwPBolgoTcc3GAmWGvbE3kBhanMDSP+sO/49HCx39rdYC
p6aIFLU5mysI0w/Gz9DGYMsgKBbeHqHSJo9xMRtCLEjx/eHKtthfE/wtq+nTuv6m
H09CINsx116bKM2azn7Svm0sNw6moRTuvIDp2pZP/oJLl26g3+UZMHp8aMVVdDEY
csAdZnalll87Oq7NtOfwWtsaWOHgYnSWZmJXE8XgSGD96ROCymIQ46OeI9InqMbG
hIAYolUCFUyik+Yp+UnMMWN9/BCmsu6TJwMxUGkxN+kijECykHZjIYytTqK7rpa1
USZuvwyZ6rSCZzm24C5yj12OtMohUG+J6SJePxUMnad6i++hs/Ud/aiHoH/vjKt3
pnMtM/z0jIlOlKZNRf6QlPqDFGu+bQyjtaNt+YoXYv1J5dAjWRv42atd/b/7luGq
Dj3298Nd9vgMrpZVIII1VXenvXM6GOwLKlh4gX8iRUBpGLykT0yVsKTvC7IUvJnP
+3G/pLIx/+hnT1AgIs13tALRY+sKeLVUprpEsoW8MT912/cZ0aDdCpGfx8SwdY84
ZJYSKcprQtBVtXTKvUKw1k2FOP14dCda14YlFwsIXvuDG9CWa8FuB440xMCucGuQ
iNEd9AMesCIMOB1WSWn6CCbvpBuVwWq/lSu/PoLGuTN2CpFmpXjrNhZkAMcOWdpz
Tr4Xj5LF4ZDhfiZ2tSMxERtuDQtW0ErCWHyuI0xzYZkL9RpaRdH6BT4NX5L83wA+
rir9M1lQymSG5scgNHkB9R1lO6U2Dgtyo6OMVMaRrkxEdTGj7BfFAPPR+7+Kk2W/
/igZh/6/YrMBkcnJtkFljwFFK5uR3qLpsrNLm+k309tTkvjOIF5pM+TdLf/RwmJv
/VL5D1pbKNf8DXhcX+dP1lN9BsbFjCTp0SlyOQNVBQaGs7JzzmPx25m3XzLFWIMe
3A+Pfw9ILc6Qik2d02LJj2RZtUzHoYQn8/KkSMCThk56aq5h0OQEfFBJzcENeRkj
1UzcMj8oveD4DYaK3SQ0S2FKxwXJc931RXLF8fCUcc0Jc5qX5Fs0LIwx/2lQojQy
JM862dWiExKPKL6F4PgfiX4mkxhPx5cr0yE05TB2ITO+g5+YROHxZxJvGQ5KZTq4
Lnl8AFm5cN/bH6a5lUyHtU69BZ5dtNwfecxGICj4lcWrZzWUydnsqrAoDC9errsp
1fVTbkmjLPzQ/T7TnXjcFmRRqcJLJGLbFbQ8k281mEZm60COpXeIGHZV9I/HTaKx
ribZcJchDhZWM/we6+X+JrNGXbsNM7EwGolrvMAs4lLsiP3Hr1J7cL8GX/tStqO0
HVLMBiwanZVYpYbZGx8CYCWMEi7mJVy3bBPaFWPn3nRr99yyw9dJfAFL/rHcGq+p
Mz8N1Dkq9m5x1rcAyrx20CTdl8gvTEGTBFvbzxoBVD2ah2RWrdeiZsAU7lN24Yh5
bzOBRbH2IZCY1qPwGJXXPFSZ9qlvt45kNmCCxFS1Cr8kVyP6gCgiIvlyttTIPb/1
lefDr3QaDkzqTXx+w5THCZS/+BMjV3wzQJcguyN6+Mp7xezARuNXw3Njlci5XZIT
N9I7uT+JyOJd/7pbWEUIKyVWAV2AzlKzpLOnKIPIxkCAh4IBE+7PDM8mVxPMr2PA
S3gYP386RVZK4WHnXd5eoqoK3HUV8OSjN54PvaUWGAEOe/DBVUrAcyoOJ4Ct+T7G
5Ag04pC9R0ovitvc7IL+PV3danBozn0HpL3bi4L6nNzPOvEmNrm6VDrNIlL1yt7m
z3IpMNt/cNp2Qo/A5GW5e2bg2JxqKo7JbpiksRpnthsnbH/6GDCRMHMvTbZU5q9d
Qk2H5unxfG/NM0Kzm1lRSRKSVIf7fBbCMkWvdXd+9o7KcEVzv2XdTsGnRIj/S7vY
9cO4FusDoBrrZ/IXSgpWcajrXrVj6qjiznF2jD4lNT74NCitqmSm5f+DuIqHuKuf
DZYZAA0CCIuy8xCQluQoy5Y+Z/ocwCJolYyzgWHz0Fzwu0raLE41mB9QVrPEaCIz
eSY2t2vu9nuPD+otxy8CbpDGrS2A/dlRYWGUMiXOcyOYae980Z+AlrYPMHvRzCfb
g6Nf5d4Guh+V03ZkEXxzz9Ym+sGYMU80hb4EqUACeW7QNAwMTKxm9eKJe3AUzrK8
uC/JodU0HXkzOs8bEh+WU3Qik523tV+ihc/5MxQQdbXGZM+ZvNjncX4UifKW42Oh
ndcFO1Ggg/j9cLdgfGSi48XxTpFrprfwiGKJGj+5gPBjdGF2LUFQCDKtAYzohIhA
HYXrp1B4CHRrPFTNWVL3maDXCbAdroEGoKFrS3INDHFonkvTG8OpM9RyzSPlER3i
rU9g5kWQZmgUMt9W+5ik0HZd12vshjTFdTLk3eGtW/ZEf15tlQP2d5eMbh8J6ZrF
nVPoEgyVkX3JIiL9UFDQSJaIBVDxbLDtg1nsY7E+P+ImjZzsrlJArIYM5U0dRlMM
HLsg2hjSKnKjUIzfCqKKYsainDjexBdWl5Nt6GMmlbycXLUaolT9OhMAaqbe0IN6
lMSRTLgqvNeAed0NJoklgVLj9imoLu2/XmOy0PURzKwpeYDExv3TXYnbSMmLsgD3
aQQNJY9dFHjtS/RnfLxD/MzMGQwm6/HHX4SRXOxhubHvc6FPyb2Ck6yR8pBY3GFN
ZkFRr0ud5cknS6gRATPFEL/QfAFpYCwkXEk7gbP8m/ShXSxRJRc/Jq9iFK35v+Dv
53UJaRTXKpp/fu3uFGhipyeaOorbKgSLzymrFrl/swMIvl9viF0ub5st8DlMbEE4
GUaNCKF9eL/jpJiqdDVYA17mRhtgBfDgrbCK8uDsbVTw/n7FHcehejPhoKmhvQ56
azFhF6hdp6LDleEDuZgF6Ee43CLob0zE5HZcbjHFamvEAnOt9LUJ5Yh6BTkchcSq
ppYNqX3H/ttXnzdTJFtOay8s13q7OhFTsqAnqC4OeoMM1gup7/faLd383xQu8PO7
dyXXsRR4h9BDgujmeScmTFLwkdbCDovnuvpxcyBffzHM/LH0BxdwZsAF3I8BoaEq
EPdauCg6/Ifweco3lXhO6HI9qBQXOqvbupM9PFiG8tvAWeIufIyKIQIBFpk3kP4Q
cPFINLCG2Yug49o0bLPK2gpuqXgKqMD9fyIjsvMdSt0QFtl7aSPTtbtaN8QxaqYf
7HXboKezRmnwgtXaA2aQK7GxxojiN6FtD4P7+1WGVvYpaIPW1S2oC2NtfLIRzlcM
iv2WFNyCi67ZwChjXj46C/3c5lklgAv2MxTr1KFkttDJ+wZLPFn/cmNxCKDTQvT0
VktXG3a52xN2KyqlSOz5fIqO3Ups7HO+nD4Dg7niNHJrHP/R19K/sotr9eT8wsBs
R36evJMFOdp6dS38ACN0Jtb59oHQrzzwpOgh5hYPmF0KfwKPZhXAQxlPYcUrchNj
REj8IILGFfNxCvFPElLfZSLm8xM2UNk9QLt3T4erZwunwnxOC/Q5iT3myyGVXcMK
DjEZGaZTSQn6cUXSKlsYDuAmG48AsUGaEwbjZlJjCsfG681URTyvgLBBXGZ/x2wK
g7HY7GvBu2XLDP4+X/IeCJraWwYi19LG8vtYknRJVkJcRjWhmeyZdGYUCl7HlduB
wtlejf71U9LfkzFFS8Lz5iwGTW7CuYwPCL7J1LbZ892WGJQtqP7+EbLIiKZ6vPVk
c5ULr90rJPZKNNUNclZmmqMEPv79J72FYXrslqRfJ4gZ5/cL/e+8eGyWl9m17khm
LjVA8rfcl+12lAONwIg/gIIPUjqfZ6qb4RAPy8XJu0hPHMC5/SVf159zh1GZoYM8
MgxM/xyvr8baHTftZO/zZKmQLT/hTv+D3TEGIFqctGGMtEHqQEMtUACvfn1EhLap
jsnV8MqRfja7uNSmy52byeK3rF4/+ZslNoDWtOUXvNRN0dRzTsRTZ+AVvjxGG00q
VHuXRq9d+1/bBr/LNhimcq+/wjJ1gUy/rtC65Jn8RSW9iifA82wNlQ02N3/zPPsr
URged+FZGVsVV4PrdKmL+c/KM/9VaVxFGBYW3c/JfI0p0SoWLGNM83K3rZAaFVoF
VBcS8Kku9YJC1SUcwpFJ39z3IK9r9rndP7LXUAj/318VqxADde/zwZ34HMrO7K4+
sGhlE7wiE/kd6YuSZz0e19NGnh59kaTU09rbFJnYLBVLOozhy0Zbk824nmuuoHXe
DUZM7MAQajRnD+sNF40racO3W/c2DCtmSNfTLnXD9At+V9rj/ZGOqzF2+L9LS/dL
EvL/sM2GqUGobwNOQyqJ2IuH8wggbJz2GtfitTVwu/7VK9Q07ixO8LNLG5sMujBd
SvseLO8mtOW3mF+EnMTfGt8Pqsw1cL8sxRnKr0OB0nI87AAO9nolV0UC8aglgSfA
/i2ZconRN33WjMOxg6iFcUkYxi7zQ5Wo0vt7sif5Ywb3EMu0EW8QH3WISjacW/6f
irpJaT0Yx6Bn+Dmx8UTPo54m0bkPq/zAxH0IXrVARC8lYm77ykX1hfwsE1hMXuYs
BPdtVim45MvI7t0JZumg9X/1K5Z3ufOIFOi1Mm0AgnzvAd4+S+Cild462nOg+Kij
02UL9UYWeLg7ZmqLsUl22KUwtt2sME4pTl9F///K9YpIFqe44SqFrK2eReu7xowc
dW5PoGoGrQ8F5h+iQgcK+Ffj6V/oGk0ASxumhrkEXvi0DPagkuBxcU2diWqaPMok
p/8dh3kwXz1ud6HSYrRfIp3NzC8CxnXX6X9wR0Azy15Lgy5/Rt2ccITORU0j8LVy
Mk4xa9eepw1cdPQGNAgDXAnBp19b93MyN2vb9uPQYFfSoEh3kcMTXRUQmTW4iFN3
K1rRGaas88aKdfO/vUPepDPWuByUrdTf+qugMMq8r4IMjK51CJi+ySViouHF63Bq
KSNc/cEsDEB3bBGaeIbsluzZHVkLNoXn77CFlfYg6cLj689c16ERwjX9UoXvWSCa
8Mg4ilEznTMauhhnbaG0H2ZarZLBodwhX357kOW2MXOXVCqGXwCe5oksEdnwxmG1
AEE6tuGmwgyujiG4lxAahC+kXXWUan83wh5bKltunwKm/1dUGTFS/Di1sB7qj1Y/
tQCxjwgUe+z9IRnmcqdVjnzS5iyhLhMDV3XnyWxg4BD2cUTJGOG265s6G+VFsnlL
hQSl4DnRaNUw18+LfP2pbknZ8+1rBjddhSHOXEEFtly41gJessaE+Bgacn/9Cqho
ukiAqeA/4bQIvG8jMB/MG55p1/upJWvSNKmG/XSqYHXCxgcmsLsMcbeS3Fs84sTW
PuxGXmpqtm3HA+KBzdPGzzpRIS8WMhruEVYxyQDz26s+cBydgqcJzMY/+pRrzU2K
v/ZVdag24ph7NmTR5RoKz3/OTPq7VeYvFCEiw5MHmOu1xzGsGWrrdqgOren5amOd
I8EkVzyVEilx5H1JkSZUNnQYWcwVirz4nbVNZ0VCmCCD8fOXenZ3sezjo7lJmwog
TtXqQB60NG0V0C50E6Jn/Uakq3A8A/+lyHPnVJXQZx5ooArDQnAN6DXNjKmwKgNU
8OUmgM4XLK3Qu1ISM+9WtoMKJkk6mem0DqEJHfwmbZmt4lIwlf3j9jVgHKQNP87G
8AFtSom7mv8MeKGgoqpl03BFSgNa5Mt/TJSPZCVUblFK+W9qI6whoiQr1vBOXzHz
KU8lLdd6D/CD+WKMa9jhlRkjPzkDwl6T53Yw7odGHiLMUapdWFCEL26KgJ+IjDH5
AZ+DssrtzMAJQ+/eBSgOJude0JpsDtNNOIu5WwlouwloardaPXIyE7XSn9uN0sgy
ZyV566W3VcvJhpO5nLL15VzJTrnhZJG9gDrZPARFzTDBsH/fkA3xw240Ko6xaYKp
lQi3yTj/pjFIMymJf2RuzuE8Z51Jplrgb30xtsiPGglIP5fEQeIztzqhwT2RbddH
aD30pW9n1YDm246II3/n6VUA3XujNiqeblFlz98Mpy5iSRHNiskK2YukgpQXL35y
dV2mvJPORdUQGPGeSBSrsc8Uq5AvrXNsX9v3WIYzLMx+acd7fDpAuzbZxhyyAkhQ
x1cOCTFfJ2G4HQKnDGrAEQvgWX/oLN8WzRTL04dozE8Byh5DX5DgcDwnB8hzioYI
YjpvmajwMmRFdrW098aQ+SWM/jhvqgnsuTmESDRoiJvrAIJ69qe9VgSIqrqLIuB7
eQvQ39Zv7Ac8xzz1Yozmc5GqvRrx0UyQdoLBOye14I2ptcJZethf8/W5O2A9YsT2
L/DQ6VhCT679MZOgWSBX80FG9uzfIQm2/eFy6y48LU7Z8hw2VUFjq181iQwTlX10
Zxt5VGAuCitJqPD6qROIwDbKT8Og1EtyUmute4QEZVUPHXBMBdJ2iiPRkOEpV04C
W2+aHHNMabgxEnaZcv5JSxNrlpSuov35T9AvgL+oa8kj2TZeiK3hJJDFpaCzz+Sa
xzT7dDV1b073VzEK7faLtIQ1i1TiDb+oUTVh6P0FjOcxKFAygy2ylWomKQRkwUPm
jRgXpbcyP+v+BrtglbHjH9bLcudMbBbF84wZxUesi5zKer+hLwOI5klhHbKnxH4i
iyo73pTqM8YA2Ik86zB65ZjJ995hrxdDn+c+GLFIYIufQh3WeEzDPduWpphTcLyz
YfLUOgeWrSoVc+cma0239uCdN+30dNkyzVnt6CEcZTDjFZbcfk8dvcJjHHbUnLmG
rpi117XLe7Zkzj4TZBGBgGE4VVqUq7UfFbM5SzkKRhkrpRx/YHVhmockWeVhiLqv
czbTCGQvlSFZjoIttvCcqE1Z0J4yD+WMTeqJdkOt6ufDq44U2w7qG/l1HD6RQOgJ
fWhMTIkU+FFs08fDgBXJ0Vi0rLxQpyu5nk6Y88reW8csh1uAYK4v3ys3RJduhen4
nKvPOR+1LZ1simuhB1N/G5oqyAie0+Aruiopprz9N5THFbyeKBGgzK2asfPzenly
EU5yzd0L6STha/aR7fz+jGoU5ojW326FnvnVXB3bu2cSd5rY+8bYa3vGugolXVyN
umPtlKSFX+Jbj9FchaYrPzCJEKFRjDWR7TtEFyyeBbj2NBsCa3oMYKas/0y/RSyc
HBJWQdbhBgP2z+j+RcEqgr4YLSTqW7A239nz+mTHPwa2maIQivP4+g9p5tKSFLkl
QFqB+2VqvRcMiRqF/gUmCD8qO/N1g7Wv/jslGukTOnOLfZWGa86p34s7PRcatEIO
QfDkEAc3omeU+V8iMNSEOZw3new87i6wJPsc4Cvy/+EOanK4gfhGGU+ZmXIm3MWX
ZdiPQv6rxRWgoaV9AvnXwSX7wA80OfWqmx7MbOdeWWt0tBZQF1lMgl5NdJpr6DFE
7cpDygYmrmtqK0tQfpVrlbaXWVsOUy5eZ23hOF2BlDmrmVkfs1Fy0wGcDApkf9ju
8nJxqVrjDKTyjzpTn6+csKgA0y3aeIrc3eKg3jgMb50PuRPaC9ajlgrez0fdO1PI
0RU3TaUlQGMonQ3/qiFHT8SkhrLLM9ybY5gHv1r3EndqGGWzhtQHdIhnSp4606I3
20UKI4S4rvnrZnq7s2GUVwJnF4hkCrrfb3zogGkUaB1sno+8GSLC4Bfjng53MW8n
FdmnHfW0A8sE4ayiPfnSOje0/cPUpQFeB5MwiEooeyLBQOBK644J4gvtVUGGRzOa
Oup8eyRFzh02Z+CeURJWGSYawp7d5V3MeI3s21TeWXOGBGQWKBpo+lOE+T0IxFYT
uli8xFsoZWHg2CmTXZW0mvgalgY4Ls/3qilVSIACM8bcW1jLqXzv5sBV5B7MQZJ/
qxLVv0igKt1t8nJ9i+EDANUUP2Hb5kUWLdi68T/r1X7wlq1+K4M4x5Y4Jm/YrXSX
jaYx+HH8LNMQp86Cr+Cy7+uicOZslo3zkwrYeMGppJb7nvRshZEDa4CfnNKzoIvv
KTEfkV3l6FzxDKDmGB0wS1+xM/mvp/0VJeTAZpsyykGfzBO6C9uCpIEry78teeQ+
SjkPwqnFDM8JNpc42ICVBakWBNUuFUvOJi4Q9TObtIGAHeWXwB5ImKQ6DZAsOE0H
uzZexiMVGJidr+Lagnp1fcVXHi0e2IneKbngXBciPX34n9VvRnlYsmeljDOCXIff
IFLzpUkSQnxTumrCE2iPwQizpW62n1mBhFT+PjiWda/hhVDqnlXggPG5Z+gxRRXs
VO558QpVfG0fyPhzTDeoXoWH0wu+PmwilaqC+9DpMHHxf7lKAoTc/W9F0MJ3Hldo
yCP0soNsMaKUfc0Y5IXYxAXwbdO8YeOxdej3nIjYb5QM8H0Ji0vAZhN0wrnkcQic
SwNv/kzdGEJjV8hH3U6DAV5lLl7UfYFgxxuqI1eiFZGBPgyVuibjEc+iiI0XI1IF
wFqJcG7x2TVPg9UfN7IKE8xO7PO95Cum2dXJA/lKcROzTDpRViK7qEbE3RBwxm8J
oksqGl6/pF90KqsCIrT+tX3WQySiF+D+n0S4EuPTp4ag6pHspsHqZOHFQqS8fMoX
KML//vSwm+/Op/9lv9yuTPbRgAExhDnipQi1Ss41K/sA9XleMR0umPQOvbryOT6Q
O1oZk7FElotMuFqHM81IL7mpgMWp17qCH/3zKqOF3E4nNOhDT7Pxyngsscs/JV0x
WG7AyMEB6AGp/de7TnPKDtgjK1/800HaQFKgrFTJXyQpSbEbRK3yjfoY060+QPrm
c+gb3SRATMvuq2/yIDNJBr5vRgo3Bvg6PQGNilI+zLCNXJic/mx9m4gDm7jdmg2p
eoCM4ivI1ORgex8ixMJQuM/5NQowz6zS3rPde7tLseZlftoSLi/SusyCbESTKdjm
e9x8epv1EUUL+0BSh2X/vZ6DXx4XMgbcIjXTN+o1QqRKMm12aW28igPn7z9wRhWE
5MCfTGeLRcfRFFVtFCn/cb9auy0DOi8Y2MQ3KF7p64DpoFci0H8vY6yo6TRMS01q
hBtZ+zGz/H0zGQUcnyp/9oyBEQo1wwIJAJHuk+8es0sRFsl+cYHneQCIbMmxeLgc
LhwcZ70DBHuIvX1/UUZdcxPZWUjIM5u1pmIRqkSxqUHl8bucytZemeAvTL4mTNAK
SlPpQNByAw0KwR9KrUZzhoZPmJ6icoC0CkgPCplpRqr61Suu5+L1Je793oUMfm7G
2ATfxTZjuW3Cpa/pzzsoA7EbKMZm1GT4G8wByQxZT3ON+EqI3jcKlz+IdbzSvMyb
xTbCCM++5SaO5E6Cwd49iFpZzUzEHuSQUlKN/Ej7f9/dpA5MdIXef+PSCtPActwg
Pw+8Rk/stwF/kXkaTl38v9AHc0rHifzr6OcK6X1ciw95HjPU450qTPI4dFmPlZMg
5RfOE7e/H6z72ZXOwRAvPSCiVOIbkb8R5Hnl2OdciLdJfpxaJn8ELbaqgdx7W6bm
Z6fEYE8ZDAn5MYcs1VnTABDh+STLX29x304/rnU++6q3Hw4fe2B6v3+JXxNDW1E9
npPYUDHylKL4Jjzh8KTkidMDmY3GNmm011rG4LRguKefGXd9fzWeudlQ73rLac5O
gtYFrpiKk2dHApHbicwgLbPUDksz1bEgW3DZvBGoiyrBVjtEzLQV/3DxtmuMRJy9
uQeATL8LHT5wQ60dbAKx8KTY8tUi9OZE1oYPf9aGFFkOB4vRlIpBL9uKhQqP8d3+
quCg0EtWOvref8y8NXQxd5V61hbNBEPPDfT7ZKdUTlEqvcDeJg1J4kZa3EyS/GD8
LO3HSH7pKG/UYjnpbs+e84IrIb5S2iBH0QXTIyNAVF+2zBiP9xHTqefzXDzpgPVu
oWVlxuJC5GozASC07aH3umnSLeV5GRMSzjhprVd0NBPXqChQIAOI47MAN/utheOg
FYnanKijluEx2csBNQXwsVgGwDkQWaWrkzwa1DMJmRiVDErbmZnTc9nEOlNws572
gesQCTLwxjKOlx9XDoWh6G4fOYyz7PU5e85WFoOlcJf5p2T4matTbUzNREdDtG2p
ebYi0vUz/sSLryNW/1BIbPMcr59Z8jK2fZuVB2PunTnrsJgWVMNecLU7I9cRuEbz
40f+S31u93XZ/k0pqoWS1By5Sqz2ah27DsjYYdBM4ATaVmcBeVyH2XSsvAcFAx7V
ldBCKhTLvaFBdx47mATI5DWm78U4CIRrl4v5IfHZ/BbqOQRAcvuKvXHUM+kMdQd6
0ltWr4RtJSXVQ44WTrtI7y/ncWw4/G+XMCRtgJEXhtzbRDfRxKTLayo20Eczoop+
uTPsrK0xoHgw8fqxj4NxmDfn1dD2sy3ZXWPpTrLPSGsOI2QtdjDVzxnNgZAF/coW
Yg6ZLMRUkUL0jY0I8J0VrQH0RAXgh3VnrB8cO1EYyAmOBylEYVjwo6eOjw8mrTsx
dq91tk7/Tf2PbhE9VJnkSdoA00iqjIW8sRvx+S3iZFyxEBvJWEnxOTgEiRqsODSp
8JPzJqccnESm5as8c5hkkHov49mmdgyjD68RKpaBlSEi1f9F2b3FVr/jppZKyPIl
FDYWB7Rb8JRmcriQaZnPZuTOvigaR8M+/s3+r5ib/InGCUHkh8r+Dl31wk7IhYVw
fDMKJMgO4iXNju7saTtV5USmHLX7WGh2Ipyd2JCdcf9CEi+PnL8kC1Du9HpfgKL5
Ekve8vkZk7iUIICInhdcOKozPUsyLCA9lbj36kTfENA/iLKFsOY5v3PUxvfB1iR1
E2+EblYVdYSmXcrO1BjRpIJaExW/eGDIwRXaJUoDHEd36MytwtPBZAz8Yba0H2Vg
ye4sgvPmnEqWwk9qKcwKr5sBP9wUu6i6XTKnZ+TysWNos5ULjd/TAhAbMKdtDjsa
2GIJtXPDzkkTKj8Yle3Yi2wTrAMIOejQmqpjOmWpnUPAMwfEReuUpK4IMlkf7iaw
MZELGiTGIrbC2bbGfLY3r4COhojrMt6milmkR7z6RcNHbexGR+8U9l2DmDXhUG6E
SWQzMjUUsz3K5zcEoZvmmORU9eicRmsuP1J2h/f+TqIigkDmntahriDYrsIuDCf2
fZm9wW48V6pcMzV9xEtNuW941KzmLiW4QeNM0oUwQ2ZbYiz7DpvU8uLueZ+TzmlU
Vi9fhwhjbUg3glK2ZUfyh8nivmFVbO1WNdxVWnPXBcBhuESSlBzg9DIN5FcIDAGi
JmgT/pAzFJcEpvDUZiiaCH7lRNIuQYjpGVtELsKZ6j1yrUPmln+kVu0P7ny2f5sx
3+roo/ZXREYcI2vc8wsVtPD+SX4mXpl78KMivLYT5plwfKrf35W9R0wBiUFOl2iF
Tm4iu1llubouMBoEdhgGxmjqhbANKvwdnBKjuNSg2bY11t9u83m6SMAVtAvrDL82
r0dHx0k+sFUDV5vgAm8h2jNTFjX9iougucEXfSLD2Twh2ox2eSZZ6MLN0PnX4eV7
wj1dDt+51QxfKyY7T4VGLalYfEiEZE36rJrUtsFYBh99r0vPMhECl68h5LWPgWK0
U/3yL3fNXlY0F+6LZkqzm+5SOde5j0R6p057N1MOJgZ16Vr1H4uwZNYsiiJ5v/4X
fEoxqDdzm/5Q0SNEjWiKmrE+zymjMGd7+RUJccDGnL6WO+wp1oZCbklLrCX18N2E
mOehpQM5Cd0ZjPM2Uxkj8JfqRrLQZKOeRElWGalMLuwjCKEo6sg83cYHBkDa0IwE
GbT1XX8ejN7pel2eoh/MXpm7AqURxtG++THR4PHxcokYpR3y57rfxjCShXcfPM66
MXBzKzfNK4Koo7Ya9lRu8Z/4M4r5qkcIbYDt9t+8EYcpwksE1a1UACrZiOBBlxmP
93OLTUi9Pg0dFFJJ/aAQ6xuUgowGIBE9p1yHqBoHPzPfxWFiXf0defw2o+HDkzFU
LaHx32OJLC6IkxaMyDL4gKa5Y4bb6SUv5FllexVEGf/vKldlRxLQ+ZYJS2AydZQH
am93KrvfEpC0VohGl0n3JPvDECBmW8av9N59cDR/VXXDp8OZDRi/C14gq7iLU4cP
Y6LBmAUBm4fm8hCY7iBxhVrHFDYxi62Q4n3N3YW9Yy1HGPWGgyER7ekMDP904S43
pCfgeWgKZv8IhvbJMxdnJONBX92MsN18NKWvR+mqrjwln2MUrE29RK76r0Gotxa3
Cr3fAYPGqaiSPvq8dA7QRWdjJ9zHj+hgYSCnqbO6r8ZTWkF0rc0QNyVagbq8Oa0U
6zlFyisVgKOHdtLLKFr7vFRFIAoZcK3rAY7tHYjNxnBr9AWLIEqUPeHHCtYCAMLr
F1oQ/VA8lTf662kS6oPY3gO0LyS5dcuYOO3kEnN1sL/DMOJD8VGTqZClZHgp2IVW
5uYu3pcG7H0+d/gpn3dyEd8BjdG1sFqejJ5H/I/yH9IxsMlFy7zYbos4GytwI+FW
tD4Af0zf8RW+ize+effgybRlq8W4fXZ6tnABIUqO8Rp8BiJZdITksz4ZqPf3dem0
trTA+HvT69JbYybWNmjvVJDIbHRXaxyfMBoxW8VWv1fG/euCzKbW9/ebgSAMUgtc
jXL+ALczKEQvLkArH9zv5U6OP/quBEdJuWsR0gzqvXBGNivoQPVRAhBCwoUUUZJX
2VWfN7w3rMLbnCdTn3DsEQUe48XP9D2yirPeFJnaVYlDogzOIWcDl9vlwlfGZrpt
M3dpKtbM+6gkhbNlwg1YKSU0NzGlBniQDJy1u2EXCigHUEjeXAdLcBU9wdwN2YeQ
UgsNj2kLlyrM82ZThtU72d9Si6pR3pNjbC5hUlnyIyhHy/nKzjyny5Q6ZO2vcrkF
PN1AV+i/TyakYfwAjBwTTpt1uUxlzRzhZA94MowqOKd+Pf5XUZNT6YyBsS3enctb
NpHucLanyaW+CrT0Zfxno1qRRg0q9JSMArPljKWRiMH1ZcI7AzViPvZOh9qaEhg+
DgECHv8UL2tLK4l2sct4X6o4ZXtrEDzF/exmmYUJdKV2T6FVgnliV7BLUUGYysFx
JTDKnZkrrr4n3OdsF+JW510Z/6V5SVRNouK3zhJko6vzod0CFCj2c7TCkDYabUG4
1fsQDjFskN7O5E/BHcBd235MijjrbGIRD/3QMu4mIcH39s7UZnHx2rRB27p9YI+i
lPXcuqnz3FWNLcYmSwXQgxYuZ0nokYBBX6GQGt6CnMPHZMBUjjbzqEc2bfEQaqw3
2YChkg8Fht5MMWLeX1/kL/jGH0mX4gGqGm2eU0mVuedFKpa/7p/Dg0WihqOzI/K0
V3prZO6/Z+GF1c0DmUDb+GdlqpX7dcMyd7h0T3JtYwLw3hyMmR+os57I19e9FB8Z
Oi09VlocFU195ZN65a1zzR6GKaDeTIfjGusIT9Wq//+CnPEniqwmjDUSD189qgyk
y9kIZp+Tu81hGKAbQzeSDR30BsOR9Z8gp2xQLfHsk8BC+KjTiq5t424Yx9933m0q
wWLEQ+ijO7/1FvmbAFQOT2gtFynuvMlKW3GK3hKNhEO0lvTehqAKVsjxmlm6Wxkt
8RYKa3KjLzTDC1t5xXxDVOyzakhpFwo5ocXcwY4Z1LxK/Q8e/cvEjxyQFUaoDbWf
2ZVDst9HrS0LmLjN4jlmIDkUXpJ4T6bGQRrYGlDraEibJL3Nl02jvx0knEp8MeUD
HhIRQ16hjhWsk/xv2iIOlhG6QMcJLG+XIq5wGGhiOPCxv0q6a5QMPoUJWzRXxu1k
PgtHbXVia9ah5YVJqlbNmDH5xqDpp+za+lULlZgOwb9W6V/hPIHfjhaHYcrGmhZ7
c6q/dBUICgV7VBTv9sSIEUy9511wmlha4c2S3vnrMuVXKxL7Kx3QZ1COr8Y5h7ep
IWASkfuDz076HLXFxL9d5xQ7V+5Ok59WgbqHWsPMh3XH8g6uBydj3bIwG/ZEDR4/
gjGmp7Ne7gMaP/rtskVzjfjAmj3wZS9lSIUTTFL+PEP6IO5mKySyS7MGwC2qn8he
8ypB3j4LkgwFuKL+tXDqA3WXA0NybB5pJCZNvkDCWWP+Ehc1NBTHrZStGzsUghng
4FcYOTbKs3fg2zsoUBFRd+ya9ic/lJLrNiKThN0ukuep694+QmkFjxbHw0reV9My
D+XQmFheQIeXDYceXTRHFIICzYHucvNTctPTWOxcgDIoqwUQloSfybbbFmnLBTKC
khBeWX4Er+BBxIlnb0GlPZJTXPGtDy5LiHOhA345YaOlnvRMD3j5VKJiFIQY7IOQ
JeU7o7RfZ0ztxPBIRCa4G/zVMEykH6bqLj00g61OdgCsInr/Aos2RGrtsmvrxQlh
a5f6ztrnYHFxOgAxgD8tFNubQHBQ3ShGxdtTHms3qMVZdr94Hz6uqaoiHD0RxJgK
OsQ/cCIOdWvMT3FCWCrhohDpN5mIq/jcfb0o5lLA6ctrBOMIlK2ea0PGc6Xz6PtN
Gm5HPXrwjEh/nB4F0SYq1wyo5gtqmGqfKpK/Ukj8c+UvuhiMqG/k03blTbprhPSg
aCxtS1vFmxDax9k9PiWXs8ebhlQc/r4BaOAiH/PuorHmxBwh7emZc80MvMq7H1U4
i68v40UkjDXkToeYE7fUTCHaqkKuzIpbeA6CgxMH1453UnCo+pi0154M3m6llIiH
0HWPD2R5i1MFvcuLyiU3tbA7wH2L6T5h0DUikqWZtOZ2PKpwh40gqoP9p9lcXWeQ
5XKNO9B62n38yq4DWCPmjkrpfhbeaS2JbkTJOhh/ne361t+gyTyS7aAcRN3CloyE
MNn+D2aN9CLKY9xE+dsv5/zWyS1pdgZng+PWbUjDpD+B3nUIRx6hfiBwrewsRXxd
jyXkM3agWae8/rPXFYGzCB7Yh44QTGcZh1YfGV19FYQykT9mJD/7RMxx+EvURzgR
ZPzE62i//OTMF8fKU2f/T4bq/lHAG/PbFT4LeeMepOmtm1gA6D1Mjo9U1aFOsitb
Tlo+TJPDf+5MmxwF5GUX8FxjZqgg164uqpI4KETU3l0re46tPfTNMWo/bJ6e9AP+
FW5PijGh6Cqu0jrF5U94AbyJjXeZIbh3Aa/8Rg1d5DlqDJBDBCviKVlRQ/RvUA6Q
jO7PS4sSUfd1uevpmZxlX7LPO1vYBUwoSAtmnhaxkDDo4O8z3rN0Za0ZC03iV5g3
t3Zf/9DiNBh4+FPg8u/CHSgR29HYwnvMpG9YWYuhmJWhOk63yePl+Fk/t4gCJQP6
rXY06/XM6TJ+zJZ0bwJrFIsJoeSGElo6t/BlHm3FBZZqKzF/YBZZ8s6x39EfhSZU
eYBeXr4yXEXdK+HxdzJ8/5uWjr0ku10V0N1cTFkVoBfIspv1wo32fYI/JlksIvTz
XBljmbLLDEaCdlIpsBxIPs/1nlrIyLTUukvUcXaue5INtWDA0YcRyFAKyXTzKq9N
pNm2mArdIRBTyWzp0PZ9AcCUY0w9Sj4aVLf6fx5NEaULpk8ourTbbtcNgIermFI0
1ZP0njGf2ANCoN/YmobwGpADRiSmRL4YYDR5rQ1fL8tOLXbUaaPdljtSK4SNQ28R
UaoW4sVhJfqV8nAR7RMJRHMiA3uXbucUODZCxtlJm+AbKPJlip4KXWn5ZXuAS2eb
ZxC8jnoPAxyT3/WoNyg5jtLEkLLlq0P/RAFeT7a9mUIccKcC+hJkVYbJiDN3YuTK
scrarpbq3P3jWYvy4S/gBwlclJsVxRV0zPyr/HGnM7ommcsgGWNvVjcBgbwZk9JF
zJJzRU4ECBDsGxr78Nc0b3qkC5n36zVluVsFMs+f0hS/0hoQnluvXvKIhrh5EZM7
5MIcw/Uwg8LxsnhhpKuM+/Sf/Dq+fKsM19nRr72+rtJ+mIxwwCzOHw50WU/HUH5L
F/4XylJkpZWFxFRUtc1ZlcfUw1uF4ZeAbUeW/yTOvY74y8ill+vi/rCNwjIoSRBO
N4CQxzSRcGJVa9Jd6+IpanrnqahH8kKw1i84KaIp+vBZ8t+6HE2CnmMh9ee32WFC
HvuKq4Y04Jbi1vn2bG2g1rLnluCFXmmkLkCADcrhziULdQSH1+2lFSfi/bKVKZ3P
JBvDXMg2EuQVsmK1wEgEw71+JkPKPAnMFYS0HSEOpMQymS2VOFm2FQZX8f6ZHjjf
8ZRaTBzsJ33LR3HLaAci36ZI/xsNwiS7E9S3e2cmluDtd31K8bfMcHZe/3p/9ism
XryOjmLIU0w9nFXO+FGyj/PnpLuBQC+uqcjz03AxZFjQsy46ZJ0BkxnJRsy64m9i
HRZNZENI4jdGYz7tvdaMyx/9Qnw1+Qzg3+SKxUjq77txmS2if2qmt4U6zqI2I1oA
hdr070Hm2tp7lK16dPMI4Xg8HpmJihzWMSpVfyj3d5+PFtt6ZADQNJYcW2Vlt9s+
gFmPbvBrdj8wpkKinznifXplX0VDVvON3U3FlLBj7v8oqTT2AnhyEqh/AMlytyO6
3WyXVvZ/gZt4GFEOS0wfnRWWJ+dCMslbyrmPpw9+Q1LHUm7ysIA6zdQAQYEyAwI5
Hjqd8/cjNtuYKZTbbtabonGzy0DJLh84h63JeFT8/WuguBvqfQr/siFbtFbeU8qH
ZUcQIZiwA+/pU/XEiZSltlz9dqAL94XO119g7nhW9dlU8ZmAih+Ii4V+Ycl1xfCY
swM7YtFRtYssbOlT1zgYJqRZJSv/VwqGq2BSSi6o6iMlR0ecmHTpcd4W4W7Rr7zR
dxBCKDUkwsTxJCyx48ua5kgwUeDSvDQOGOUVvW/TpXbXBH/yDHJPItVjShleAUG+
Fi3e0Inz/Mnp0wic6Zmg4xjhtpz9ziKFRa10z0YMwxbdyhYsS5/GlGz1kTwkaC63
gbEUpbvh0CFYMwBw+R3mhppiLRsHk0Dghm9bDSfYTGi4tSQsimt4ELJGiFsnec4X
HtOQebz3oPkQvvNFcHmv6LX2dsg22qyFERgD+bYcIWN3/4HY8MQ+bl9aosCnkx6a
a5ejJdsanqatl4PdwVKMuwMjhNaR54iVFzmK0XuoqmQojbsGvcgZbrBVKxzXydFJ
0ek/8hltMSh++lhXh4IrcCKiXiHbW17MPNOmRPaglFfmrsPI2VqaJSL4NEjiJaTU
QjdgDsAya0TSH/riffSRimECLUdNmk0is9dBWTXoxmn+P69qYs9PVtKgjSnlT4oP
InX4yM54cr2XQk92dxhF4RS52L5TmjyPNwzAJX6i771fg+GbfIIeydCT2kunMUF2
0f6tKZGuIEmHCdLjXQ9uQriRDUIAktJ6sWY2al38xgzrzamyW2rt5daSjRfIuolf
LJvjlgQan9S74Y4MUkWa5Q3eaMoESRQxwgszT2/3V85aleTZL2fBpcMEz60qbLqq
bFrpCUDAcIb6b90dp1jV1VI0NxW9H+cAnBXlWeuDLuiY7ZuQy1e8mq2kKCxmkXCI
NPkLp1MLtjGaL+4oYumjh9ogFOIWnvHg5STComO+UlhMHQ3LueqcXzKZ/NOWFiQw
yKwLM3z4mbNNqk/rJT3/0//MwsDZuyEPksc+LTGlhYdphHKZK2BHAADvYn98tMAm
7Zn21cN6yoGFKpiRpMsmFBM5aUHWK7LKzTgGRPUR1PAaOIJV8y8ur603HYX1lyOd
CkezBKrhfDwJd7IdvZn/3N36v6JEfI1/YFDwTIFgnoojyGi4yUhZihcNzQpEmv54
/lnJ4PAigTBY8Ox3AxlL6KdrGccktrllQD+U7SnpBjZSVhqxKxTGk7+srOpsSscm
gHKvd+CpBoID+IdIgoBUQ2QidNR/ccjrdlOGpuVxnTgq+Jg6YrTDft8iHIoYNCc3
x3dT+ULxNVhoUpPj7iLZTmVwtWXA3Hb8DbEIMiV9YBeJe0H8oDGCpY1g2RkFDQ4k
O8q5BPedsvWUHs8P/aCOI23y4T2wkXYxgbvHGBqIY7+8cKZtILRbnV4jCummWHXg
XPOuqfilU6Ti0tYleoaGfMgC9ASRjAL7zequIPrUDu5XpIfh3wBPi2otiIt+/YNC
7YtjwknukRE/HJfKvQp/GzlRboyi7+Z39gWK0hopT1wO5v+l5dFwegPA3GMF0OmY
KlvI2IprB5jWKB5MO78b+n0hrZfsW5BrvTKY3AISkS/Ieix/tjMc2Zn83xdAMA2G
fWxmCOOBf5NRn06gnSPIK61ul1mCbBdfQdcCWLLGzR9bxJMsgRVZXPF9TSnviGt3
tLk0ph46o83s/ThJ+jqI0VmIEqDIf562vjgTk+RNzWR/YzEQMzAJmB8SPtIUGbOv
ZlZGbbHwIWS0nYZ2SGNcV7lkOzVbPkl5mTkiiJt9y46ymL3WFB4AEfcTaq4JFbo/
23CU9mg1J0ho4MnbIY1y5GurNlnXlzfW7Ti5AfSFie5UihSxIJHe2OHCh+JDEhdG
/QqEZbWoC3z0JH4X6ll/WkhyKwckuGPX4rcMiEUj1MJ9ZIEjyEGbXXwso5qczTKQ
YQ9NWBpY/QoU+z13KZk61+EUkEyvclytXHvl9d/L/obSXzcHpWRTYFyYu7J607hM
G2kuEH0xmaaHHp6NLRODfrFiSuzp3qKTzYDQdnZbrMZ8yjSdRnoHcJqvI2+RmJfT
4eyj1YTLkKlSRwZR49PUai21rTHwizQy7VM+5K8C4/DQgHvNrnzLcyZ/97nHD4Pd
ZDFnBEO/TNRoSng66kD4TTZnDUAT3tPC1DDR9O6788NpuDUQ+7p37VvBKRTD80cB
sOwhcFwnW77AvKltHaIdK8grEE7NmTTPXVNEQCGd45mK8EC4aER8P8mSdhsFC028
aypVaIjdAw8mjN8oByNuSKD1c9XZq8gi63Uzol6/9pdPOEoY+QqzGbOVGGQIluv0
YS3hqqtfzOfKP7BTsTmjqfazwu7C3Z/9Lfm2aoq5zJWc22KPTDLjN3vG89dNx2qc
okUooeUF3xJqq9noETKjvjXJc/AxWp63UNxXVEunbnzVWpOXjjiKDff9ojma92lw
CMPXreD6/j44XMFOSKJICssa9SHK4s9oz/Xq59fMwRSyzqHAgeZ9hSzpkTpvEHvZ
Z9tHbM2LNpr2uE//w5T9+21xTKUhnnTk4fkDjaQb+DDXBJ6rWRvLaVD/kHBc6BvD
MdI2MYtpy5Tqlg0irUN14QCP82p5MzF8Xssim45l7IsNtqnE7vo0MOCOR+OkI1/Z
uXX96t1sIA/WTfdQ74vXhDcHmv2abaXG8+EO/twl1ik51b59fI30bxRRrurt6YTp
tpxVdEvlVMLLpL6UlwtXvz6/EAvqzKXAhAtpEatCXtnJ1iu1lyxFDDfkqp7Pb3jq
HNJpiyLiusUfYDXxI2DG7XMNW/h0l1u3rFdVvM8hOMWTNDy36IJ6rX3fnK9vL+N0
lkk61GDQiFL2AP5WdmawgNWlp5GevAl3k1In3IDQHHZnRVFg200drree6sVfkBI7
m6ji7r0nI9Q1wQkLRZFAKlPrm1KrMnNYpQPGQVg5ZXDUjkF0TMookUaWfJocpLos
+JnExZ9svyysy2kTNqMRPZ8Rsu/4RGmP1QOWhx44M/UpMkj+fJqoNHUaAa0wFCJk
2yv37DpQ2bdZ24LbuQccs/DUdIdy/osXawLaQOeA+isLDGDmiyQaLaejzgr2qexq
53rDxyvcFT2/sZS4hSpU87YR1kWms2t+C2iYRVh/JlAeiLKa0FEznQfzpEZjuv31
jYq4XKCj4XLXxEQeqZKpeV3hvIUlVjRaTKhJ0cvN/l16yVGiRnFIntBSUQ8lNtBg
WDbSnes7KzE4ax3SmzTe6y3TJkT5DuLL3D7+lOtj6RuR8vbMyxSxl4H0VCRIe8+x
DeIOieHnwXncIMWysQZa2OeUlCQcn3Er3nYcuKC+sPV5d5zcJ4Cf7KfFIfxLc6di
ReuzPuwU/N8yXQ/IFGpVK/0d+A1DxC2sGnbNCrxIzZpRJyXy9GkON1y9vdaj69Iy
X/RXnSIyrfarQYva2pRwHhwe1M05B+rzpfH38wmzebaSdhYpd8nyilFeDIweVvJb
cLK6OIilrdwQohT00RUZtJLlo+ARhXG1O1m2BzcHySw3PCjaKqFqeSD3R6ETyxhq
kHM+2MnWj1JOVd8e97NM3tr1D54Z/4UveStyoyQk7dIyxxwJgIeGZSF4i31TbmTh
ty5xHJPGA9A41tV/i7zOkXgX1kB+TtZjBMu6YxlHe0lJXIalwfNHugno6EX2qxb+
QRRtMgq1v4Dv/zGJr2q+lS/mL+M1/WY6IVjzABaioBp/Oj5rLlOLADoPijVsDThT
uPo0nsJNifDHrudPLhVKH1tYCVJn8sE1PjVsgwRrTZC2cZQXJVx4XmEyBPukB4s3
vitcQcR/eTgp5b1i3KoPSQ4rKeLoFDZfwbMD0h3YH7J9tU3mWMbQrxHOtDgDb4Wo
FhwNIpgyJUNiw0709F4AWCOU8dZ/lqHPoRF+rv9cwY54FiSqhzP+TdNiheekTdzz
5+Vc3a2Au8U6yWcxuUtbDgqe+ZJUcw3UKU42PUcJK1Kn9PpKIFqfsLGJzWNS2gQD
MRbKPOPAME+SWOBmR+jjmWS/iZfAcqJDuh1ctXbhUeEBZfc1fFUhm8+Ylskr/LDQ
zF+Y07cWLcm0Kfw8uO3okVAc+jKmwOKQLxF8UUHZVc5VWKM7Oke/RooCoJaGDpSK
+SVov+IPoNdRpjOofoKsibtOmlf11gzzXPMYHxRPFfq8lkvNgz+VZXRw+0vP0GPQ
PUtJFfZuUwGBm6Rlb1lwT6vZbJ9EL3Q90TLJsPfDSjNv8KKWyiC9GsrBHYcFwJS4
ewKT0B7Ng4LIasJkdfUS0Gy8ecnpQID7+Ax1OCrtq1wUvO0O1EmWx8bO5J7bCkbW
H4BneMreBTJCWJbEo2kYxbYkawNx7Yg1mD2t5qin/Jz87S7XNxeCFBWyzfZcsGRP
rySE4/w6rNtJaNqJWB8UuIZ9KsELMBbgHQsGibZvUmrsXFtvetVhEJsYN6j2jJwP
7s8QNeq5xLreeN5yDEj2e2/2u4F3zM2Q+Hz526Bb7H3c8v3RW/Qrri51alplPu60
D45rUrF1pvhf9fkTx5fyQBAdC3xJ8Rsrk4iYNVWsmTbAY3fhRRvec2wltTAMeREk
4d4iNg2/HRgHSgeSaJL8HOXEaweRPS5NDG55G6p63mOMELr+H7lGzMrAZeNfJ7+I
M07Yaq2BCtDGX6vRi8EW8FjYuvRCiHwr8JXj90DG3E2eaE5lcrdUYjshpmql/5SP
UZHeMz5jZbvC8+6zpQ+bxwZC8hoMvbD2KwO1HmiIqa7HHoQovQlU33/TyC3PXcOX
+WpQMxAqv4Uc5L0v+nUa2iBqO5a18mXdGszqOnxjIrnEtiFf46jIhiftI0I3GCze
hmQT7Pf7G9Xi5kI8l5wWSpVbEKWK4SUZEGGBv/dtXVsX4DV90ZOoqu3PbUl6sb+n
C6D10UzrRrLndx9jOgwxAVKfM2fTek6JDObYiCYTBBZAVfrRPHhUjm/scHbbGOwm
cNUYkLyDhcJTUCuR5MhgmLKRE9WrIRSGVR6DhQFZSe6ISy/0LJ0Ihi7nYfCE0R3Q
xCnV2i9a6cy0fQIjpI7AzpFrNH75b5LGFHzy90ZKETEam5oIYFXp5K2y+Rt1qqhU
oru+Z2gDnPOZ4P5mOiJ9/A3T9es2DD9mDSUGBDsBGaIO8GfGDT9Q7fDJMY9Yp0il
ACovfyzvtxDrwO808P2mOz9x516DZFQYjQW+dN00HvOullPaw3hZ8z4zoOhwZpml
+kx9xiXfHP0/TW8oaogGGedr3WhJU33Hcd7pyVtRUbj0P4Wx9l4Q5u4JxA8XCmC5
S62kk+OFIVfAup0AOyFKIv/AsIKUr+1/XYNcSfVmDA39gNCq6o6iGxLIGqbmWhkO
tzChZHks/aVksl7njRoCaYviR/sl7s5TOg/7BMYiUdB075L5ElE+dkQYWvK9/B2k
IMND7h++KZ/56wDlJYesCsRXPcpIF4tscTYWxnAeOFRMKfxkA1ZtdAicTxLWW9f0
pX+JRUGy+rLSnof1gyIrT5EGsR9+AiTqIaFmj8F3+prk6CTLDFLr1yloItHpZR/g
AODNEibaIrk4TKyiabstfMRFdiJGQjgcDPOyrTt55ddru8w+a6N4yzP7EOfGue2P
SNEpVBy/mGHZdm/Hd5x+jb5Yg39HPZvC1Y33j18TA2gS2tbuBilX0iXbRVjFen4V
CTUiRLyNMg/q/eY/nXYDzrJTxs2E9BVe8DmZXzBkuynrhmhY3PJnWOnZKdIPJgBs
k+eYIn4Betfwl/ZgHYlgRB6VG+L3JSc0Gqcj0uPIQJmDaooKJotmTZY7TsFgY+8h
DGmx3m+voCysGHzAOwjyESm2g9OOq27xBf0d73BtC9yxW2AFmBy0Qh/5XoqIsM6i
IaaUBWHxrxNkTaqysGisbB4/YsAs7/pk85ZuIFQUk2gWqGVXjId4IdCIJepNRQOL
T/tlXFS53E7lIGjItmzI70urP2syNekpsKpFlGfKOePJyMdKf6W9nISPmc4cvpAb
5EiMlxc8ZSFu6upgiHLVMJJGELwFgUyr7td4t0mSnX3x6Wu9JYlAaSsGyrP6TuZb
BSfOUs9oVd+Xk6f8HDF3XItKhO+NdKi4i6kRUq5PMV/3GawzkPKrIxvHDZO7BkX9
GAnDV+KyK9lOMcGyFRCaBeDKhH32e46yCeANv9+EKVdMKNFQNcrjLyVYrkkocZK0
XvT1tkrKwWQFFx0boByw+pdHlNBCxSp+WXbynzXpP70I+9zFODkfebrb2meu9xYl
IEYedp5zCqJ86GmEBmAdQAWTvTrdQBw5iDHPD73bdhFWq29q56AEzLgdmhDSCkAq
HF8knGcoGagDH19R13C+RwhpF0d1ndmGnTmBhJqYs41ABrKG4oXiw2527hog/5f8
7ogk3INuNfOxGHAZ9iAiWA+ENWee9q0vtnECshXnQ/ud7XLVK1mBNxaKj9B+wy6Y
JmRy3RLmsteMjMsDqBW9JCmytszdO8e4hGz5g23CB75x8Z2l/erCpybFEuZfMybg
apedCEM0WQmuJlrewKJQboDy/gmX6zO/7ncmVou7rFp5f9gh4IIpCriQy/+s7MoR
bhFloOPHrajX8NGGUS2FHFpPL6WSdjjJCN2mcjR9ZIV8+cDvJu4nTGBP/2opJOej
rZfqKOCCd0QMwVkCdiyIn9mNaN9gnhVkIJfHaLFhC9a8z7Jyd99S/p+9Ipk6xNoh
tSKDKtDxguo1LOyO0+P9yRDFF6ADNedTV4JIA5Pc/+Mbh5hqXcxzFQdEGX4zrWu+
ocxDWx6pp1BfT+8Fb7n2Nv4dQBrClLhfJ3mo8hQW0AlmvCRXV8aIMljZs01gUJ29
AuQdiGQw7jNlTeeNY2y77NCmp/TdfPF1ce3R6rLbgbiEDG6NHjZR0XpobfwF7etI
btAJVF9BFx8aOw67CeI17WhnLYZp6x3DgEPn2W8H/UqHg28JEIgXWeDYU8YLLG6q
1XajHptmc8p66C/PtgAxz7kmDGg6oMqWBjqEK1H0QSZzHodlXtpNndlzUJ7vVqB/
A6RyGFx7m6uD7qU439Ys74cXPurf/xtBhqbyB93ixsC1NUi6RCb889UMQfftmdGT
6akfpK+kIxAYb+WnY0fQCJFhLBV2DTxaU7Ewpy00y9Q3+KPatR9VJMVI+B//IKW2
mfOFjDunsmKzRfQcmDHiQ8mCrJKjS728egJNxz5HSr/useZG2mRcuGMYbnmbsxn0
iyk+Pxs2Zx2OXuKiYApx0fsrUD+Y/bDcCiRU4SFfCWVZYGtqCEs+8seZ9DM7dIZD
9YdH+h/dNfY71QUOLVTw76u96w7Kf+02jwm/oF2GeDcMWMSZVVa0ny/IsMSMeOGs
x9t7UIUxsj3LboAL0RuYRnVEP/QbwZf3RrggZ3KrqsXDIZ56ZOawuFDFiesoXqY6
iF03X8hgXIkDxeksRyXzg2IfLj8G2RtBCRllg7C4A77OJEHCPdfaFP7amxJBaCjc
oLaz0poB9KX4BOogjzolh4aa96wxoFRh6vzymb7etDCnla47clhLsN8Qn59XguWK
DTyWybTJpzbwiLIrq1B/YR1gfSCagNHwaYD1YDJBEsHM9EINuz1HfJOdCCgLSKNM
rkJYWcL3IcYkovPuhQ7DUAcFFcgVi4YXHgeV5UPDqj5s3evR+zGNQfQadkgorOtW
ftIrblqra9xFKfePMzS/uzyiw9gfboK22OmbSbTFZVMxf2gjPyTBCXItfM5gNFeI
NeuFBZB0cmWIlLFB+uxEbLniw7onuk+1GYroIW67MT/FSW2nuyHSmAUP7xa7JjHe
kF1CWTXrX1hmXileGvATu/DRvHsJdq6J3gpgQ82nRfkghcgCXjCDGmhciRjFwLn9
oYTWDHEyYpkKP7LjjUiqlHtBClo3lUCgk0bQ85H3a2nK2L8Vnq8gylOsuJ6A+rlN
7Qt4c0VHTh9+N0S5S99JJs85XDQhLx4ysaAlX47SgaogJsgIYfHsggHl+BI4b2Tk
EYxw1cTHD/44omiQZeLi8pzKf/yk/orR4MDOLmREhndNouQpQe6LvhivuezHW7ew
93t/LvmaYMqYuSibhHhkl0h6J/MndE6Kp9zrHth0/mPKAPlSK0ob89PagMUBJwvz
ujYwEQXXhshSn2MVdRYMeNxiCzUxIh7k/LTzpj4xdfAsgAgELEomVaVyg+usT/Wx
MVt42DNT7XodkRxeGpOwcZ37SqD2HvUpWzc/1opqu5Q3tEWOeJfAlAZTDMaiDxdQ
ol1qngtxzk/IZwIXEPdZ3XlVeKhRYmX6i+9xeiV79R7NGy5JW0yYLw/B7V1kAqKw
4aDZFtx7Vh1YL3CFw/ttzz8/C0ydk8TD3cuEcMnpBEzI/5j37Y1y7Y7DOIcLb/aa
bNLCZWmCfHNufBW52XRgQl4BYYvnNOhCF02Di/4TB5fQeF+ZOPdMToZrF69XGgOy
vHOuUKOWRM2yqzCec5ACgsxPVEsvHbCH2MDj4m0voljoJD4A7kMdql2IVg7MZpTF
xfcEE6nSmVdr54ornnpL3d6qyZkM0f6Xtz5RSvxoTxgIXRVOBCJIazprnSubfk5K
AQMCdE7VOQZA4I3HbD6w/mfV3XPlsOvgFtWY/cZeKP/1vB8KPXnKRJlf00p/51Ts
3h652idZlTbwCeiAT6zn4HlgyNiHYnbJ3M+XJVWAo+vQr7rwT5FPzh4F8+Pus+3T
qczfBl1BkFeuXrUkWjCnt/JD6LeOkUNTW2x5fCIDexCaUdeFwA2IN2VfDvTfgLX7
6jEEmy6ih8Yw51nX9MyTOgVvf0JbIuqBsbyErDfU62jJT168DBfZKwRqXnKSmtHi
ub0iZR+2civyS9NzZk1uFVcrQtEw8u6X+cFhNM5bXt4qKrGf08Ye+ZMcZKANekVg
AiT//xjmH8SNFj+n6LU6gq5gegCL2sRLjNG/zFeee1EHReRWSD1xbqVz8Cm05k5Q
jEH2+h5AljI6WMZz0tQsf/6fvbCzdOuQyrfsafDrIA5FjH1dSkmro+AfSfHasGNq
jQ/7k1KgkP14kAaZopmYQWkNfiRupNutpC4kz3oK6xDzlVxIpoR9jGewpD82dmZz
UKp6w9yVg3utplRmgrOGYfnzbrD6uZrq5BUnzEKmDiMbwaayHIeagQbSMu8ejwoH
gcrZN1meKi0e8OuHVZI54rIsCn+oYf82Xsu6IxHwOJQW8g/iQxdJXOpRj31C5zS0
vBqM6wRgoLgwjlGERqftguN7lDoCZR0/53MZh6WpYEIYLmjk8L16hCZBK2WBbWpd
o+kqHzFCAKKFwAKt4ndzaTEtOVr3TVrMFKc1bokW1Nh0o33tqMx0c02Ki2d77ear
Eetd2Dj93+zCIv2bTSTm0I/1boM5CI+iV9RFvwzPsxkO/dquR1dsdVdq+SB8eb95
mHRe1BQdADVWK7zMoi6ryVeni94310Qax1RQZYenNl7IjmJ6ZZDFDIdt907+JUGH
2rAavpasUjJTvk6m4wNYyEvVTVk2Nfzr1iWncBhqQQLGoOtQ1RlQf+8lnudFMbyH
UgOUNB3uSROVqW6VUHEiXV7+GoTg9vBIqlFhKAlsmfuenSKl8FByilEg+c1fwsmo
64vjywn32xezmiornP2rBZ2nzYN5X0zwybG4ctKANHGjHYvf+9dUN6ip/SRd6tV/
TzD/om37HGrHK6ODc0i17yzdWXWvdwXIaUtReiwSSc5nKwZ5XPg/2y3IhaT1nqUi
E/jdzTnzTL7OFUl+2S379ZyOhoV/SOxH+oppxwdee+mxLh1rBXBrAR/M2EHhgNA7
0Aa2kldJQyiqF8NEnO9f18wtfs/M+NjFX5aDxrZPFRtgBQTTH7UTB3Hqzxut0fRc
YiCLe6whYjXSa+dKtCzwxLm/kf/K971lK7xriiaJ0kIqNSr+kYTFkjR5zFXK9z9m
NKePtUKziEpG2GTjjglHlu2Fmk/AgFQ0t0RZ/E/rhfaASOpBZ+B5fk63AGuGQOyg
Gh32/ilgLOt9QfU07a+AplGaqRAwkuWptTG0wcvQR4wuosaS6x3mY3GODfscduej
AevREU/iLTL/n64lYXb6N83yV3CwwprAxaO85qvsbbu1XmH66LzP7WqGCbcjJzg1
SSgUMJi5Su0baFn5YUMEvGNxNL2GEsBxFja4wZEB3mp8siYYyhBlngrg8ghpVWC5
NmE0ClMwR9zZMXYnI28cM/bY3f5IfsS3fLXzX5VKkKm9vKavDnv4CI7GDWesXhEu
hFQpjsUOC/S9+6tN3xAYaXOx1YjV4AMAINetg9QZs3KOj/cahnGsTKtr4JeUmMSA
wbmWYTRQIdSjP+QsU2y+20O2GiNXQiOVa6IC6CfEVbSVfB7G/t8AA6J6PqRRYDCz
As94W/fqolnBTxAcbmNEPiUeYgyKGI7Cx7OojMzi8WIyHrtEMFW5OoG/WKRO90Oz
crqvqc92/A8Pcuaov5utTrE0jlDX6lPMw66cPm1txIbWwkpRpefL75KxFW3EZ0qH
0+nB+UAnnf2RYeKk1yW3+L2Ju++fZA0uFJ31rUQfHV/w6p6RefVULyD3gg9isx8V
YylheWoEKz5mcAlkEq7JPM4vOac9kXLEWD6aq9T/L0zSurf5kNXsXamBEts5un+I
2vuAHq27y7I4QtrC6k9qWZnRzFQgY5vbZgzzezx53Hk1HyETrNThEC9YF2Yn7Zwm
jDVNHKIh7ZpmrflPzomduz9nukIn5QO8sZUIa1nyPvbKEi+4ijOAn3+FXg1uWhai
UwJULkhstNW3HOu0rZLuS3+fZBEp8tS1qiHPFGx+XgUEH6rafTwq3hZmUVj/ECxt
7CdpGrrMqDc4bWBQ0P0tOKmdroUSTJxhO1lgGk+6Ts5DFMH6VsTi+/lJoNox2wmo
GBTsBLP+2Gu5QoPU6LeyA00sy200JOnBE3LRRCoxgxBxsQ6zJV909dRs0ZFX3i29
xjhQkVRkZfU3bu4sPlNFcmnsGQiWoU7eHskUOcbSJ4MaoRBypa/JJlZrGRlVzltf
owCBdpOpya/USFafHEdBbAHz8HhYXxpZK8ZPLSjKHhJvNMJGPM2iv/W5mzLC1cEz
HqtWUZNXzeZAq3PY5DhVExJagQxdhZuESsGbrMt4y+dpmYYDeO3xXNK/Wv/e2vII
LHrE34eW2TpjkJbG5X/DYQgRDJwJKhRXVmATKGcgiRVQRoc/kurdsffx4mb2KTrm
OmMfewZJm357ML5wKdglQZaXReaUnmfuCnHCm5/CzSPgDu3XIjdCVF7fqETL1I0b
X3MoiReBtTwIkzi7O0r3poHm7dyJs4xVp4ZNj/O4dUdwAPWS77eDj+rNlqJOMUH+
6ajR9dqbHsXh7n6qhvWXttatzdno1MGOSQSaZx/CguELQ5mj56L4xMBOxiW3rxVU
30TI5HCb9nl0Elf5ecByIMTMDfJS6sNCKOPAXhZZYscdeuh0/8IVSxDjLrh5ibKz
4BF2xGJ2rHnnMtew9n7hDYr5ZB1VhjcqT/zzDM95hWbaewrwl8DWaKxZjsf4jnKI
C8DYKefSHYExiV/D8wqvnPLcms6+++uGKK62JhQTGZ8dwWfoGiyoxzmpe87yuJN1
+Lf02SABfZOp1KxtEnS/LZljxGMIZZgblDPpHO++qbJ7OweO5MSe1fz82VWxpY6I
BRiUYcGdqqe0wTLLZOag8gIXVxqai/qtofjuzILSBBAgRLeq0lNM5qfiac4hrnnN
FYS5Mb6JZp+QglZig4ntP5kNkALJCsG128uePl3aa6H1cNB7e25+ywCKPGvpzUNB
f9vEnAkNqJhnQmiQboF+kJDppr02jVJqAMGd+4W3R8C59xk64Qw6RR0BInaHgHsL
ESbX0KnTgPu2pXPzOTIn6umKXzAtdVCh2S/8ZQIIYExTaOA0GzAKs4LdutLx+JFk
ScI+bMtgtDzM2EYpj7hFQDx7V+RqyELxee0kDkd2ajccTjYCMX+diwVkWdQHnMyz
wNYe6B1/83mwdy0cJrwA6GCl4Za91ScviOKHDFk3eIy/Zzul4V4lmLvLoTyNcRIG
5SZgbKcs3HSRuB+Sj2IZtcrjO3kz5cDjtQjBQXTPNnshc7KkJBG6/CQ+Dg3/X+sq
5XXoWZ8IksFZTLsgS292YvVipgPvC9XDNKYzqA6DlvazXzTcQ0LODJwD1pwuiLBf
aKKjhzHo4rxjlSP8I8V3gpbcpf2D5u/lkxbG9ec2+dsJy9rc5Ozmk1ANpzNW1m5K
v3CCbJpml9Xd1xi9P8aAvth4JASqhZcKywLPKoPedLwdALbjDQ4XN0e1k2VjVFuL
SvzeiIXgS+FbG/VckJubLvSh4k7aeFLYWThFnR4NUDO/gxXDAQBLl16RU+Am0rGN
xmj9jqEU48YQ13o7YqZyHb0gIX1yLHmtGhuPP/GLv12kg/4cyJrbVyTTVzqzGDoD
/1bpk5QnkA5+d6bCs+/fAXugwM1OULaJ/XuKJHWvuznJgHHVObVqU5wEhDRY18er
3uZ8OJjB7t2Ukcuq+d/cWZUHRF08dLDZ63jDy+O+tYpt011aHvsHNQFz8kTZ8Nt6
ww9Y9Fn9UqVvpm1fGXIr+Ex/xvXP4+LEVmqGbg0KuXds3DiDZlnH7ImevjmmIDrM
98xxBiNQMU41maAUOvFdc/IuD0vhc/GJy7hbaH9iEfwoaB69ZgROWF8/FPDjP+7o
8OHEx/+8BD8U6/qi1+J5NBqpx38RwxIfs42EFBf+uRcGc4aeKqfMBaM7s87BgDps
Y52rH6sEDuOIbMCpwCBoD4TgQWOx2+K0mG2e4YUgcgPX2lcUx3ALfgc7ngFdvT+7
ZKiRt/91ygADbHNKP8NjrjPI94oN8DvmSpkqM9vW0QOI8saAzrsP/4jxO29nzI/X
a0MvHXFBcpQeBo6lQ5WYNVJS8U60fX6HSUvrbo6/fHZsc+VE4MvGjYvfJu5KDp8k
8GOjPTxwq0TSdfm/8GHRHyUYnTrRT48JK1Ir87OinMrIEERSjbwnbBeHc+ouFZiy
0BnOjgaGks4gMAWZM6sfYs7M/G6eCO+wCVS6lMwwg0eCYgfLYpJLtmkgwnh5KeQf
RMC73VyAtuNokstx8glYFlDnTjYN9DK5ZpHBxCmmlT3BQ6SXFMqDtR83A2QrZa2m
sZxTggAY9p/IN/vrjnoF7YpNBg0rnSmufokMvEjIfiHY2gfkBIBQsR0RcUkbnaQI
Si5zuJtQsGCQQgh4VBSi+B4J0kxB19bxBy9kWUUkwQohDvKygkETPWKwtm3E8gwC
xRtP48mwNuH8uLkAhXB7mQZs0It3/tQQJbCe9jSZCbsD+ftPfcjI0g0yDoNJVGp6
jFgAKRb6bwQ4hIBSi041+OKt6IlGQxnMr2iislpb3Wk2Qym8gj1lrj8Y4ndX6HI6
2tAC9rhCCRTaEpsBQPXpJEKPDj+NiCbUgG5dXWbde0qxzXMRGdWYilkoR51Elp0J
4itfObdqu1sra6e0ecS9WS5TuQbJYpiywqbMdraCs2o6UNAfjt3iEKkmDEGmryHQ
R8lH8z7YLW3fIPFxt8hJKandXA/IJI1th1ZzkK9e4XluyjEE0186ew5QRAYL28RB
8/6LfisoyuqSIRcOjnrMrXU/1Qbu7quz78M3C78dkelWREZ8BEwnCudUwkdAbzIc
5Ga7h1QxwE1PEWis5oMya99ccGu7q+SHA9DkgrSVJ1GiFBSUZIxGxjw+Xp4C3zU8
6FKxm9kGpy3sglduzD+VZX1bQ6zV2zfrK56n0wdOnPZFNt205D8NsyUFpVa2p1nf
nWuGM/Z1fBlwUo8V85aeYvj1qLecQidR6Qr4xB9+H7jVd75K9/qw926wY5V4HwJs
iA+fmD0AxDKEI3R3cDJ9MCY81RVtgUEeQo8/OI9orm/BjWhB1K7ehY09/VGi2Idv
NLWUnOzjOQq8aVx3Ka7Re+yt+vCsIvwgBxlZ+IGrBgNZ8UtRd3v5/o/u/JLn5Amd
TJWoJK3wr7XT4Gvrp9aeIoGUROhiUG7ANZTJq26lOcMgP+/Xk9Z+QcqysKDcuW4O
1EjMo5rfSYvqhHLtKdJegrEOo3rQDfQUqmq/G2ERLES8A3JlH+BzLGOi5YA9btRw
gFl5a8TQSOmk3AQkFqCUDJDBBT8FjHXg5nBRfVgMmt+bckDVb9xUzPwlzUz00KhQ
W55paeSmkqGeANTz1ZV7Lwlbd4eBDtMwyYOYCBFCufF38RUBAi4i8vel2Q6ZjRj8
9inPQsSVPOXF4afiWfFbGovBQfNCMfBNmmLO2U3wPpjAdNmhJM1FAhN7qygNTgmr
rSRgAZxhH6L6kK/djI1l3MNtErW/p+ATxJm8G4Tq0XrYGcM9qDadbCMQkzORKmwn
htpYlD6TDh+tD3bnCkqvR3l6+F0TqYF0A9EBqAUYbIOzWe7Wbkcbv0lSA4P2Ig/m
/jb8sxA/nIlX8FZgsaN4LyIwuzHXkr/TnmkHlRUbtWQVL0sWRunQEAhVm8KeeN6E
8hIfB5EvpKj7VtSeM1Ut2kBfATfOy2+8479G7BipWkNf/MsOomDttHP7GKlrJce5
mf5pUpljQAPAp8WLQevhoSmsW2I82rvxbpNrPjulZJlnEKsOepX4+gL2CW08uGsc
swmzhT0bONWdmLlMRMhaceLMiA85xLzB+ekLcqDeeEv9EU9zwVIVzbyQF7Wk/6LD
GXZgPVKTvuityqy2wpxHUyL8hCcTaCH52juLZ1PrdMR0DGadeVNpYNQuH7eNznDg
cSgp4F3qAJYQY0v4wsRt3/HPZZX6wtSQWAg0B4dlP8mhl16iG69cU2+U9XmIrEjH
MSrPjqLSgYBN53mPHfGW4Zv5UrkcXbVey+ypsT1deSVF/LZh0tcZoZz6y2EhklEN
jSCQWOkkgwMCSr2OF7IFHl//yelU9/9k3Qvi+ezogzrYk8t4wndTOlAJ0mmtzBiE
BQ1R54FnG0EolmARX3NltN8MNpEM8EvPjmoAg44VFco500Vp4RY+O6GC+BCKrmIW
4aTDDYseSFEFL+b8H61IA1nR+3dYCpoEU81Tfkmmr0Eb5MhcGQSApeph7O0Hfv2B
xFP88Ft7bVzoGdJJzSrGaeMNVdHhUjY3K7YkadUJEKw25Euhp68hByRT634mIkg1
hDGZ7ncZ60fqGKIPiQWQONpmh+/MVDmRIU/+YwCCLbUIkJcg2Vi9aEST6+TBKzs4
2jTiL3uNKKHFrqLsjLHcE86txAFj2zjh6JuJ1OkGxK8d9xwNo0/qiG9aNSfJRbdE
Rfm7sReQk5fot+G335ePDFvrgiHXBsfb8EA2YG+bu0M3q1e1HNtOGAUfm4tcw0Ac
fZ7KF8lZC9wZs4BnAuEiWHJ4bB+Yi0ZS/oTRdeL1wN0G5WnqiUjrjwKsbabu/OjH
2Phvlmv6mDm487p6sItiEj6qcuZ55fwfcKmcp0DnpsESTASgZRtqO3lkD2yQLExu
EdrOjDFrjAxm0J47uv5QI3xjvaBpTYE92h8PlQSZcYy8FwukpdsPkBxc8/PmMyEk
V3maCCevGqeXNT0gJgyG5WSexNn0vADrab0au29IrVriLVVugY7UMk7h44HM955x
+TAlgns8q3jPTi7bvvKhlDuTmtpu3EESC7jOeHa4FnlTlAuHaP9qN0l7JUtGHp1Z
B4mo/NMPcyEggtUSOwM+EyIQtF0UWLNFLhrKz/Nu5DgyULQA150aD0fch946zVl6
I8Iy2GaOEaW44KEmtIAwpRs/dubRQ8Bp0O+rzfObrTRulwdqGKJS1LQUqFCIORtr
ywyf/ebyJZjccF+og7Ip+A9fOgBR+y5GdIrvM5oh+CIQhcVTObEfr3lsajQ585wB
W29+6chAhNwfUdLj0wqmVnn1BlAowKpridCjrjaANQ30EwpHNRiEpSnly0IptCMn
+RF9GfakRCvThw4gtca9UzNQ0X+To9fljGmPzIYkx6pCUD5pXkylxeCHW43Ls2vE
4j/bRM0sq1VWsyKA04s/sgXzkEm/rkCBsiFfvi+igfvo/RSirmaCpUzzhXSiy6PY
PNVGHMFsmmRC8JNQNTlgJSs1ZZYY39afW14oobsiJ3G8lYDtDxvtTxL4CywK8R2Q
7xpxPv4ny78H3vujrByZ94YDWmi5zdEwLBduuzPZGWRiE0MU8bKJos4fPf8nTSp6
rVIkRrcH7GdLmT5+eoNARvRh60teYzxChxeaGNiJh7J7x6d4QWj1ElGvtVh5zhOG
jIQ6idbwSokrh0t6hVqVl9OXngihXalsupAB7z+C4HKWIRO578JhDbHP0t+f2Tzl
q8DEuiRPj2I6Qd2VcdO2Zsx8mFP+VrRINxzTMpvlydW3B0W+G2SOE4b7yFyZCpud
B9iNmjBQQBcbPXvaJZ0J3Mfn7nG3eQq7oZv0UK23Rx1gJkwjxptS9G5C2CNFmNgH
VhGM5/fy95ishyQu1tpgpt/z8g2Yu5M/6DZmupLHKtB5fs9xm6FAY5iyeODCGVpf
QPb5ymnzBp2sWxwdflOSW7ZHIhYUuWGqDU90eE1bjxiEUwbGKcgRBYx2BeibweNy
Grlqxhd7V2WSKXrCdluy4kgXPu84ye8UExnsT8dETXajS0DTj8Z8l9WEXx8myIsO
BHQuSGu53yJby3tNCnUb63L/bIxax6iGXZ4hNFJo04MWg9h3mGsQShM/b3FPBPc8
1iQC78TUmow+1bidCe0BHodvCEkuAU87QqUk4zHjUFvwxAPwoWBNjoA3F43ib+b/
efoqJLKHW5Ppizq14dLYocgS2Q+iSFX75tubaAEvn/3fP4R6RFV9gYq5+tCvnbM2
C73EbKyaatPNzZoXJshDwRYFPYXV4xosmYAjf6DOUcP/woFZ9+JiEMqKqt52r3gR
X8g1IOOHktd3LUq7Qq0fxwUmFYDnvFRE1vDZ7hkl+qHdZwhqmUbqNRfUHUur4w73
nMuyWb0Qpb9NoHHagtU1C/6DZki4g4spaG+rDna5z3vimjKBWMUAiLRK8RLRp5H6
B2D6DUA83G37NioZ/BSK1vpXqTpHXHN9E3gyhVhV84FN3DTT+FoIwUukpQ4GddHb
xFBI8Ditl54LlZ1VtSBKrYm3xf/i0t9N5PSTi0Ttbc1puQ0lsxUssH1YbDenANVm
n5dL99sb1PvpdEOkTTmu9eb1bvOycOB9RZzpuYGxtuC9NffzT5tUznaPPoIv0EE8
utTiX0rmdHCDBwkhzpNCBkGe3G+z4+V8yGaWhQTRBFNbV2Vt3dopiqz42/qX57g8
ug2pd65xx1Xa12WpUQ5UVNsO23DUcMOiOJn1BMftYdbXB/zujJad+YEwRrI+VWfk
0oG6OA4R4FYq+t8B/5aoYB9uj0R0u3P1OM7MsupK9oQOpg//Gu/+M/kkwQdSTNlA
8YF9OIOpB0eo3S7NkqLtKoxMq0Ntjmi6iuPCXRKiWvevFKf9dqW+UbZYZ2GdX2GU
B9Uiv+w8HKl7TBhV7HWifzZVV0N/3yGcTLTzUOIc4FUz0+HtcwqySWABVhFU4piQ
1uFLuNwbiZ7e3tavchUg8rEZ8Np0+EOBKxnK6f1c2Gk/hwKPj33XCtnvrUwWNceA
rrTRAOXf+E3Aeu/CuqcADvWZuA7UtdB8Mqnv7bE4VHjVDCRRaqmxYRYZo/a+83mY
U18xyaDEkJjU/lgtUZrnZNsS1aIru1bI/rwdEpWH5N37qTM41u6HpMN0mUHBEph9
iuuFSls408TEMUReg8OVCCU9zj/eRzG25UxzPPCv4KxZoq7IRcN/Hg6dZL9i5+6Y
t63VdY+dg/EDmG4SgQgSkATzGJLXnwMq2lAg9lwbQZ1StMACPeNQFFS2Nszu5pTi
ujwogrHSJ8Sv0LD6Y0aBB2TqBQFJp0hJqOBIzbG225bkWRvLoHhJmYpzYBKweJRg
f7FnPt6XJYhgZbsg+XFtGNqCXCgBR/8ZI53u8VyytHOPtA6ips/zWoipiEzeLRVV
2izvPKiIHAAhev4fJIekFkGthMBWKyTdeBi6ydYKMloDAe0sJZPP1BsUqEGxgNM/
9x4mNEi5qhN2LBSIVviIm3auKbRRF90lW4Wvvyk/4cbF73lJXkJ3O4X07xdLLAmb
INJbukWxb1zjHzHs5PW6okV8+nZ5K/N6+H7YPpiyu1vzsGosmd+2uJJMr3hQayb0
Q6c+fPIY1mXJ//oW6Wz5XEXrKbPTEMbNiAwxVHvvblJF4/0o5qzRmOmIYkjB3M39
Ot1gvEu8SSZ/qNmlAb6H6Mt8mIPNKYUecMjGuIZc/hSlBK4epjFEQvzJpSHu5yRn
MX2sZ/IoSSa/Aw6OmvrcLFp/9ZdkczA6Oyr0JC7UH/KangMlM5vrYXeD/oE2QiUx
/rbVjntp4/GGR+L6NZcKXXtsloLRGwWeNgBZHkqvV9roNmKB1SK+nfUgffjomvTO
Uri+QiT1ionb/YIbk2CYVXidSmcC/rRjz2vDAZN75K1RQbwzVGhQ3iTb+l+NGVTO
1/XBMu0+XhTxpvwQUNpIDXUMTFraRTWn9Lgj0XES3b45OC3wzrJofFkypJZjmFzn
wHWzmn8IDYOOYRt5Vq2pXbaGS5ptaT4PTOA1lTNuzQVjeoXdZ498dtbNgFgZ5eLS
ErqDZoIIH9sMY6JkwhGWsSz48REaosRdyODrMfCFd91agvCvywP9go24GTrmGQb3
F++SH5SwPiNtPVGXrXcQW65tIKd6yr+tSGw/TN0/suIs8djwPd8a+2sTufdoEj/e
CHNu3p694m65Gft5Cop1hQJSnvh0nQ2eYAKQcUuB/qARpnTNPKEGklCXZVD5jPfo
Sb+PjyfdgoMEcZPLyzoUWannvvUpe6f4n7oYyRJGky0jdQDmYe7dTFfAhuGYY58P
kZHYvKmIhN1h3p61D3nhsVOjU5Xr4ByEVF31MaOH+NSrRWgU2Csuw/EtLz3LUOYC
qpF2JuOp1bJGkhV30/mfiAggfbDsMfels4NZePrJDNq6qNg4jdDHpz1nAMZ1vn0h
e12hG0c1QF9j9HK5csBd/swMtt03WKYz4CMkGgy/r+2VmFEd1kwk75mn8aoHsgZT
0L6kj0qnS6OTnzHxJg4jFkuAzC1hcjefQwMCpNCMaf5hNcXuMJ0aDsoWbjmGcY6O
FFWNEegp9e9YZ1on0LnhDVdSAcl/erCmk10ECUQ3MELmNUDl3Av1vwvfFL8qvwI/
COVeBTwPSpBIeCArwDOqxxxDAJhK3ZCsZAfWTScI+wzd6YYjmUMmdELedlRLLMFd
WyZhPdn7TLM0m4Je2++R9ibgoBM2ptKeg4AAsOKkrufO3Pm97W49er7ulIO3ofEn
rnOUeQYnaiXjWgq636jslCi/jpugLEXUn87yA9hSWKXheX5ocz5AFbu5qLXlrUKh
hcHHTngi1jylfgWtPYPQbZECkHuI7xTWAQro3oJi0m0tOaiMV9OQR26UBWgSbujS
orx/5Q+OPekzTZiNoq7iCtsAvguWYNGwPssFuhKfrUKemNlYFtVvWfgqG9Ph3drj
Y0eqN3CN3jl05AuOo3AWVfjcNcXBvqjpjol67I6n1gIkh8KYU9kRDwbCQrj/3hCD
UdRlfJw/hCVtj9aGKmwxpKVPqFFghS3HWYIu3GtFs+Gv1odp4dXYdkIA0OQfvBOL
L69w0ZDqBY+yNV125gqZ55v1rDidvklHPhJhrgJcgsB1+dPj1Vrk8KREIR+ARXh6
SwzRIWgEtvTUJZNTQOpVS0y0aMF6MoRUwwO2J0TLUhUK91QWrcLvcmfGOjaqi9mw
AecYfiWQ1Pzchr5/+mvqqlMTaCBWRELaZKptW/uLYzeRQiKWgpti0RWaQKKSDkDP
mhvjGYhRBsmCmzHYhDflbn/Ozj0Vy5zQTAXD5QzsCmAZBbGkXpmX/eyVTxIyVzfW
/xx3NnEfYlRAM//DbzrX6WxZ5h5OZY+Th7WGIIVH3UD5BGoCYyFSveVfwmhK8LS7
bI0BpAGt7SbdHMYQQbcU0kecZ9i92rjg4/iUPyT4M6fpufIOoBaDhds3Rp4Y8Vqy
sY8o+vX56vJYU6PO/VCpPyrhEd2om9o+MrSkpCegijtQDlKTXX0Z1gaO0ehot4i/
FAtOhrmFAzaoKGoemJX5IqduRn/zwOSm4r4K/KeINM/fzNENm27d7qyoTIiOQN+v
LeQxiKcLKArWnx8+aWzgOWcNHYTVMc3C7RzUYmE4FZXxLvdSjRxtpR2/IT4+FkKJ
I4SOuUp3oE7QSdHFAkQmmtZA6OsAZNv50NwBMK9ZrvUQY7BLlYENGzG4KJLtWysm
h7d/oBIMZkLb3UxF6WFocP3OyGqMyLsh9BLEuqOzTinUy4QFEVNWEGoYNIxoifDC
7Sx7weoMN66lQ40hehigX13H3UCM6lCX5oNHEQDiLYLZnV5npi7t9B2D4UDThA8r
HzHyHKbhJdTZIE+fOSrErwb8fbnxfxDZqHLNrODeNqf7JMU4XOQb2E5f7X8WDJqM
Px8C/NfWI11XWR0Cfjo9a3Bi6Efy8EIt2eoD5i9ZLYLJYDf0pPQ2eWMxN/6h+1bw
/6c0zzQQZR5zCUYEaiHbDUAPOUGOOyixZdfEl6HUJOnaFK8+fQYO9eNDz0ANT7Mh
p1jfvFZsFKxaJtqMEv/vp2gUVsF+URcBiTUS7hPMErUd3tvNzOQWVmgjfcypXdvO
VyHOFKvPx2RrUR/S4CQwQ+igTIbozr5koQtf72jFna4sHkKhX8HdYNkaxTZB6gn1
xpphDWjtY7JIYvKfUJ79ZOpS/qazTFMeTtRiln74qQqz68k42Rij8Gc++m+Pgf69
DAXr6CzjzRWkE8g3o9gt6UN+W41c7KNztgFjkidxqmQGwp5O5otPBTmQy/m2yf1G
pzjrNmVivDjk4GLzr/cnCMcTOpM84tqMJJTylVNm6gVlLbODo0Vg4aHMaMqSykb7
sNhvr0W2ANBbC+7cjZ5tjH11UfBpsu3+ifL8s/c0Mk6mCgLjlIen92SRoyNCzKkv
2iOoWw1s4nN+47KYSND/AUN4yqcjXLsy+4j2LPMr8RxsyoY/33KGFdIqT95qqk1u
7UnVXXsIaDs3wDIvp45uIAKEy8C2pncNJyD9gXKh4SJyY1EZpNfM/m7Ux1Fghc/3
YLE9VXvsJaTd6b2cjGkfYX7vV794m+LHtPBZw0q6d++/bCvnZFliQdWS9j/4vaZE
hcTOUgywiutKjy6eBypdVtsdh0nIWbuknQAGnC6R1Gms+uc0oLWfh3rdHffpWYkf
7wOmagbxTk+hMG6GkHMqknEJK9zihuO1fEdpXe/lLfOf2UQZ0pX9A5w8Fy0Hl4r6
lHLTpeE8BYGqy16tOSzNjvc7gA2c5quXBhkXzJntf6/Sr5up5hUG358L4dzhVnma
vOqjfNjXex2hXaSyLksfxYCbzccG+rBcQTY/knlv4LxnZ2EPA1odlSA+5ms/lILS
pmc5NiCrQ9MfJVOo+8LcVJIh2aDCQcuCzhMtkCM1m4gP1TnxkicUDXnn4pkUGHr8
ZHe7FPW2JFBvrXJ3+or0lTG9T8rjm0DR2GysW8uC5iV0hOOb00MmnDrIGEKHu2od
jA9cMaIdPqn0kbjAFFpGgCPvcz6S4E6kmaVACcZTverjbXPmtHC/qQMMSi74Bjmh
2MvmbHo8kV0UYjpnWpJNxf2pILUVeVg6CIvJS8vhfZHOK6IpomRnuJybbxUuW8VV
KaiO9ejJQV2cPdlHVCIUOCJwURcHNcWfzIGgd3xDo50F9ftRmH+yRuA/cUx8QhH7
iA0XUrMGk+2IxB5pgCU2TZC1zFeDcE/Xt6WwXg4lE5oHHNod5yyPv3OS/k4Y3jm2
K8G0IF5xVRvF0tyQRf+sPL1S+rjtq6VqFkgNLcdMFXidZqyMieoDV463D9jNW6db
eRu/fUL/V+wXzn6Qzy//79QtgF0+1YBK5Iwgv8NuAsjcfQnTmtsTtubi7+VVYZP/
q9jc6M4MCf66du0zET0CPMscwlDukDcaRxDJEvaAlmuwwXJevEOJGlx2PNWOyD7C
Aa5Zv7FhaV/EbZ0S5MTOrVrjp8616V+HAGDMXMr8Wc/CKd+q5jw/fU8rQm40KzYy
L3jgMjnh3GErYkUcGycF0lq/eMVHW4JhOFsaGwxsUWDOFjs79o9h8FsFCKZt9oH4
0824637Ch4JBu2ffIIm7bdO2YcdIwu5Iw4nX+p7Md1zmhpeAhIrCRjTCaXbIL+7K
JBzzdZ+IXoU5SyKjzFpRvsx6ecQ7k+Pmf3E9aP3/CJU48oZQvZ3IJGiL2LmeJ3Fe
8/FdzG6nzQLa7K+AwtfKjTAU2oCPo39ElLX66adKjh01rwmK4DX1u8MAqfovUUv+
xpbnccxfOhxULexx0txDGDvx12MtZVR+88m+pBZXN73wcjwYsd3CZtLIerRA8ZjG
ESNZg8Qx1vZRBPTNQhlgg1xYdPe/GL+8JjiBKcWB56xiOVw8Q82zYjuXxq7iBCKU
MxtBaqdyf3UcP6i3aTvDwQh1X4IYRMuq7puRZf4O2KvLbQRzqDdFXs59OQcQqnuW
k4KfKijAsLPGvDXE/xKdME8VhyQ5b+OiuYNpe9v0mk4zBZortiedhVlzgayHToJQ
nBqWpFcFbTrnKfzU7aszgCgssdcecq8SeGk/9P3KOW4gDDJ4vrrlTx6jCpymBRIQ
osmsZYHwF42cQoo+xolaIVAkew84V1Be4pY8WSnGydgLnhrHLzgFJ0+mUZJSQokh
TX7qy6QazVfaQM6auPpGj7Uq/PsBCHKLYWqzBwNnaHlnxzppbL1I+Bdz8Gd4rq0f
/5f8bAwp009i22jb2gxzHSoaBsAG1eyMb3BB2BckG3bnr5nZBL5jDV/vBpL71BU1
NMmsfK+q9zW+nqRPiQ2YFqbdL+zkGGRDn/vTlk226bpAnG3BFp2ZGdSLAd/C+egE
7lpQYyOegbIhQI+9venA8btn6W3byLQmS13zaWGW0QaEI0Wejy6JfGo+dYEqSTsd
QVVmTq+HDTU0NYyyQwNJV2j9NAR9NLWqK9Qo0L3o0EaJBpdVmcV6nH0ZcX4+gODy
zXTxfMF19WUQZH1kqNT3FgoQDeJs/7ePVBl/Z6LfE46upFq0MmdlH+wbxmsIzAvm
k2Jxf79MrTNeUzlBtMh4EDcGZVAOBZQCYSiGNhWbQ0GUqaI1qHIMGBCGit94z2Wd
+6rsfEwv4dyA9gAFq36WrBee6x1fPOe2jNuKzwqKrw2BgcgxXbIrbB4yua5Wl0KR
I49EUj30tG9XgOfxRy3KXTp7Z3ehqFS3v5mU8aE73geqWJjSxtNkHANFFO33L7GZ
CCBAv6s4h9vftqdoVLOdRk2rhnSDb6naG5namoAiFwa/Ct2UU7UtY5EFWw9R/qqJ
jMLwDPCcq8Bu9Ucr2+L3xRCw1sD8dNnYAX/SLFUhxvYH9gOIckSwrU7vLL1637/f
p33hs5V7zFueN9nGF5diHZJz0UuwKz8FbdSZjnGuCfpShmzVmwwizMqeTAAmwXkd
WcXHQ0ULQavKkyVLBWWoU1LXeJM3LwdBDk1bMriuBARZFN1gNK0VhG6DphMmzMKw
KZBZZpQBR5Vt2EfzkryCn7Dx8ZjDznMBscyyVuZxsqilvWWm7ZCvZ8efDp0rqPZK
gABItgxvZ7uE4rKZigk+62Wleaa0thxrHzJc3UR4Lke+E5Wqf750ai8jfP0OfH+e
r6fCZz0lw4uONjKm2LzQy+WQSn7caQcjnbyblQOiY8utyxVRI7CYPbfqqM7SQExX
TLyj0G0GaIMg0c2gxx6u4kzx3Oo4jQU5gQraxpiiIFhP1VO9QVut9gIApCd29Xy/
JO/0t2YwaEg1YfsGjNK2c7US3PCQK6ae6aufDWztvs1IKQLRuOGyQhZmYbYEdaUG
gdJX8xSReDxVyVqKyUIphv51BgUjY/DtkPxkYaZJ0PB8MFvo6sxEyr5Bf2sFlUk+
WpzT9SsWTPGGqBY/f+EitLAJTSjj/d5WteAE0RhVe77x6M5POIFonZRPZ5RYbDZ5
kWQmd7NEqaJ/oW/lpebanTv8nLFjx/3wlfOiJ7npdyWOVm9yhRRvbdHw8MZbXbZ6
sZHcQqe6grHSRgcEsd89I3C5Mt63BCZE42hUZcGq2ZVVfXW/FkqTYqYzb5pg2sOz
jGvRIJgqXYIbZeuXXzSKS2Q5LqhYlUqDVJWF6+8NRJV3sRkwyEN5bMzhp0QSRUWf
Rdi/cGD49Ssj/18awM+BX3GKEaIudOZseyuKKeBaCT21uYmXIqtYuRO6OPfXNJK/
QrzZ/eKhUiB+Sj9VnB+Y8BaYEDIbrGvSRlmn3vcUcw4qCTOH3wXTyqGi9yroKMGU
WKraM9NsDUoL8nZ3Ov4w5RBlLs1Nz2xW4BDtVxnqUb2MhtwfN1v7uJc54T1Y2iL+
bqAvUwrVU0Eiqo6WAaWdj6U3myKVmZ/4XEpLoef88H9qvdEIcIf6CiJZjDFh4OQQ
jvcV7nYSuYgP+IKPrZGgt/RW5mz4JJKiU8ayfOqF1ET8ES/Rz1lVXQnkpGjSi+Tx
zDl3W6w0VQTUFyQ/MICQS+yiJfTiOj+1VrhNaGtZ2pOtTTSLXU6fwmkQuTAlRLWN
TuaJ2qLEolud0HaAofi1DtbUuWEBgL6yQ3pvdLsEWxN6RKeiOsrgDklzhLPb/cJR
kaBGvLwMcHO+4imhyfUZvPcgWq/jgKaExoXexcjpTYWQdgr7ZJPLesjYInk4AvNs
hW/OL3oZNgOK3TVg8g7/FJR03TjBLXMXXMHOO6k8WkTDQ/asS9O0qwUZqZodIHYK
Ar5Glii1GaHCSzJyhqqQyhMgl/kYoojt61syrt2jolla8vOjCm0vJeilanDVoWv1
nV7PSnpiIxKQc3YtNduYtWgDzwUVIDaFXVgaDauCOl6cf1DwufVFV0oGaTwJ4275
jJyXTryNwqMpoUJ+2HKiLDDMJYU4lEizE2cDnhepTBim24tZSA2kP4gzk1wyip7W
tpKcofqk1c9tIoWMGgbvnhj0ReM5RAqza9adQIclOsjCXDW53qW2BIdbUUF5RVgC
C8VsaVJpXPwpAJEDyg9BA+muax/FRo5Po3/XntXqbq00SKztrH5kyUSn1gYEkeEJ
8xw/8tqoVJKkIJLw+w/90vbAORa5v4ebDs9YU4Dc08uzcQSSDO8bhtgb8Hsy7ZP0
jJs2dAlBnt5DYkWPfAJzvaOlpRfSiZDyFOic44iQUsmysOgEFDSSPAJHABlGDhSx
bVWzWOTG3MxN+kyTXP1dEduvSIU3gpt/Y603s4cuHoN7VJafnO2QG1JD1UaBAEUk
xOd1dqlvK4HZOeKSithsaVdgNW2zRtVbI7437E4FpZSXSqw0gZ0sE7TjAl3vb1oZ
mEnqDgxHq1XaADikYl0/dOL7Y7Kp6FYA+mgwv8MGVvlEcMhOjV3j/bX8NWDmqRH8
T5QzAJQPJZa6KY4+RpF6wMtbB68mf/dNSTPy4iFaxAjoYtqhN2DuHvK95XiSSwgr
H8/zF7xXtQyY9ngsFd+gEDz7MNhcBmlY2njFRnKsvUwkdSYNuGiryLcmA8y3Ugui
BUfzWg7CEv8CwkydOEJJJkFDw6YYwNqh/jiErBXiqhPUxN150udeGIwXeFPpxR2q
pGmmKcVvhKjYSeltmt72DS2iift1XUKzpMQR2f28IEzwrWAoMbR7D27dqMsvcQd1
KK9jW/7qMjJbqLmrYSgmETSpPgN1fXmYYvU12baDxImYsMIExc4WvAVoBNyZq8sH
7VJk342FlZMmrNpjvYKy5a89XplPGCQdT+uXuzwdd6l1n8mTXKINRLsLW7OL31hc
ujG0drcBYRxPbnTHEdsEGTQ8i+GSMkLj5Bqyj6P8V0mAmhp3v1xAqkUkibr4y4EJ
zed5OkAmhYyWUxHbqYnGf5d+SAPTBmEMIhsgkUeewgyuODR9q14obwgV7Q4/WnFq
5SU4CIwvltxmK1lkUFyfYxmObsKeBEKa8/qYnwEBiq+FJRTaM9GmdOqF3u4WUX8f
aAkZmPEjtHrKLKmS2T8DvFbULeiuSMZiivsMNC0IFIYIlSEIfwjaRxwY+fF95L7X
Z7vUpyH4gvmL5hcgcD9kfhrM+SKogXuhX9Q304ZdLBONHOqTup8KOS+QBcc0/hJL
NxcKP6jkrwS7XWMDwKBsZGZXTBGlxksAn9ZAvIJv/4vB1Dfj7IEHfSBgO7hpOcSl
gLLpF8AQSMzP11I3jfbfaBj9Gu1d3jSEgCvdY+WNYXsQ9n3MYprL88tsFK/U6pRj
syZaNaAjRQGsgYfued6tOj1Aj+GJ1ilTImM8RJthRCHebU/TZHjAp5wln+w5B3zf
PBZJxiI8QvXG8dWnYU5FVAN67+QR6vqwarVqyrbx9wKHsArzm3qFHLniY1VNOLsz
LsThWI0gULi0uGIFPvudRD2wrYDnF3ZnIdSiREf/9nLTRdbXNPnutyr7n7Vki+u+
V+68FSGlkj1BrDSvwu8rMiIBRzIY5pZTFtKuaLhZ+qZzwQm0xfg5eakY9j1X2ISb
rqn42JIrtXQpp72JfYR59a8jOvbzpXp+WK3SrHBs8XhnWDjJkLfsN1NYZCkGGn4W
Xxa7CDDf2jcWbvHZKACcm0F+GtTOWI0Lqvby7viA+8vljGHLKP28fEIjyn8Yr/xm
BvH6zQ4/BdF1Ski/nREf1+RUrO1MSdgYzFMHVcBxue/SuJ3fHa6fqtjEUY4b+S3a
q29BkcYuqyFRhcCDP0FCqMQcfw5merAI05b7bIOrhOBHinLZ66cL40fZFHhLbXk3
zEtqfEiu0WTb8BsJKOnimB65iAsgfe7LwcrCK8OsOwR/tLp2bYkJlvyRInysK/Qt
PJtNIkFNeBf0WNOdZ80MEHYGgT/8hW9Iec0YHz3lVJZ/LwL3LoXsb4sk2fAx7GVk
FQtNK4DlW7J4H8rwuve4Vc96MrENUFxGes+5DVuyylRqfapQRXp1Gjc0g1FFlmwu
UEeR5tCkFzY4ucfpoFThXkUbcbEbYfeVNweBvNoFx2efEA1dLieUlyAiBmXQCU87
8zuJaPWAGshB+vI9fMKkxPjZUvq+bu4Pt2lVNwT33Iqi1oueMjCQFS3uk3/FN7Gj
RZ1lR2YbVpykZVN960vMdpCyxeSPPdYYLpHOKXfzy0pg6AgJCLbEBnfeZRqGmlBJ
iPhKr1EftE/Wq0AP6EHCCOV02fvwcPxBlHsJgxpq9MTT3PxrNXqdZ1PD7a9oexUz
rCqJ1I27M5re660c8H9RtCJfX0uZCWUMnPc6oWOwbMGpdAi6B/JKE20X0J7QmFbt
1Ki9anfU9it2NOmRN7YrpN6zOxyfrjWVlQMuq4DwYWXKYK7CRiecPRPf9p6Kv6xt
Lg5sj3A25CPXN9/Tk1xlJjyW91eC+/MS/Zvmrt8aJC0rHB6iSPA2nCtQgFsVvSp4
6/unmJ/mt6qj/w9WydR4l6xMuzEeLlfEgzUTwpH7nBrbkIT+vq+0VaWYV2KmEswc
8rJMlrjcloX0g0a7uN49Lj93u4QDBfK4TYNk/M8GzHpPqbwxG6z8aeOICv+Fb03v
m4zYU57uqQmK04AKqV97vtu+Ks+vG5S4UH968ssj2YEWWxmJXGvf1Zhgq+NUvt9H
6xrgr2Kyuy9GcXZU01eRTqu90FJNky0mUBhNUqz8jCjnINm2br5t8HVUmP7R5i6D
2vJhZbr6pMBeGjNKEa6llQ9PnLaSKxvWk61XTfb4cfB+xo3CotICpo2Ilj8a9HRv
nheQPZQBc9JoJBaBqOYA0LH+ipkMp7gAzTIG/F7FUZpRecVTvAEtIwIiPWkPy2T9
k2JK2UaERybcXw5Pc26tLvSHm1Y4p2sYR9p2pclwKE+Ik/yRmOmYSzY4hNBIgO4B
XDvUQJUgsC84JsMEC2vk4LWh0e7zc8mUs//8wlATLg6o7jTvB9VMXX9R96PxAyfQ
gUbVxo8eQ9HDHllZAtaMww1dinVQXOqtO/rZK/YT4tY1A8srqv3e6uqX/g8bPJsd
SzRaG/Z4ACXvuDq2gqYysZw0XPAGdSj49QR5bb5BgNGG4lctAYaGUzg4WxJtxcOt
aQv9Q2cb0GxmIot4rhJZb+3YLCajpLOxTbXW+Gr+EF+jiHBYvfK7j+36fz35MCE2
LOrwvRhQbvi7Hairrvhkey03GAnNNiwST+i2YqaKZobwrKELYE7ZsylPrtWgABe4
PkoJkvy8chh7ckGGSjggsXeBai2SXkzLuo6Fgsw15E+3o+dHCd4oHAK5TxDLsVHy
DvI1gA2wR5FvuyevZAwmS//sEeFXCClhR9q461iMCXxGXE87UuCm3WqRm3gdu6fU
CvMfuOAqmIVjebqvXckFAOVGF3o+bQFUxyFpvu+NRx62lOj98WNZFmjyypWaQN/c
cZ3FgKF4rzQnYEiT0A+QFov6jpaMaJH43v33NkqmOPw7LyYNxUSjBlezV4t3iXmd
RzLx2L8yUDMIhU+tOxa2dQDyLjk3H+9or6VOYDmOHIyTplsGZC79piOMMIThR8fh
AohNQ1365IK6LTrpAelrEhwnya8k7tOXFuTKhL3UG+vmF14IK7EVd28gqulzT+Td
15PHJD3AzuVBb5Baz36rjFjLPCOeoFs5u7qJcJfri3l8rsU9UNeZYeE9Tj9D4X2L
/mSChMdVziMll42gsiQ5uuLzqPHFClkibWYses1qUerOpJLqN83bAZOXJu3DMkuA
BMlph5NfWjVSD+84o7uuSthqG/yRizeTvbnp2oqzQJwm3lXZ0DyvcEcyAWIXDv/P
qNJxQ+1Mlwv3d+IcqaryfedRNYCbh/nea1RA1vG6c95dnyLVJF4t3OqpB70NGWJs
s1S4jDDvOttSEZ5/p3oYSUfKpLpo4gi0N1IfsdWVbL8ZgG+Ju1ZPiYre4lo8Z8Ot
Sq6MlEIiddgwzcxcudPMP8Rzil54bgCopbeMCZCp8a0Wno6ELRDA+e4+HoCVuTCY
R/nSth0zkwpE3aPxy4yLR9UK9iQW7/IF8h0LokX+pt5Uf92jpiD99yHxAnVth664
wSuuYn+dCffIeh+jQy0G0SqinfRrpc87eXof0MfZnEmKTGnvxpyfiVOTvAFh0v8x
ZZH77rbw0vRm2tElIESD5gDqAm8ocRo6z61ZZJuX0kJfSITBzxq9IJ6YFLhYR09s
MYsBYFCzjPlTa9zvQMBoVC/vY5en4EkvVLl+fyJf/XvCsft8InARD/lefhYL3pYZ
aOW6ErlRUABCY3nNPOnbNRReGcQecFZcU3ux8ygmZeSabiUlLEQCF/GyOeIS1+vU
WgSxH1No4kpibWwwZr433kzaaoeHSGZIbcWLOAIe33BZy87l3+YyBDZnogj+38OK
CuDGG0pGU+KFFLS3J4pGRM22VpGkR9I+L+sWMitqTiRe1f1zfKr913YN7vdMQj2a
KR6BnvPqvEyVWDqS8U33Ch153hrH4iBg5HW6pPJLQcrt+VpjgIgEDJqZ81favnD2
nMDJoQ4GwBREGmBQBQyr091hZHp2O7H+CgdcIkbGDRUh7q6s0+tZzYzMnhN14jcG
brfeuIzNaUNhT2mHocszLgHP5NYvXsfdE5MSTM+mxq3gLHeI+Xn3Gh7g2sCovWSb
alGy5ocfAO+xei5Qv6m8Huka4WJASSkihrrb6AaUWkn4wnDVL+EfE9unpwUhlUGM
2wl/kob55rv2gm9mBWeaeaAIJL0tLEiszTyCRJO1o71gbsmpy3hSsiJX18Pooz7u
OIqNXswXKoNtDtPd1uCXogPRg5+fXVRWh+IcBNtax96N/qTLVse5W4IpnLd7cmQz
xYvQhwlDSWtKm5poblrAeAFOXUfBgdRW7bufv6nD3pTVbkoGhXFz8q7VnM0fXCPO
PyzzrTgmNdCERKvffj4Ua9HVoUimLEh5KLomNN47rlv6VMVAjsr+9KnOxjddTACU
22dy0nAP75VHSLouj2Q4Oih6RD2XNUuolvngtmLNRqWTYbIx0PtfIG0zw9pT3YW8
3B+HRP3JYyT6UxiGwW2/79fPW7RQGWeLfhZaDlWg+tl8KynKSTQ2ePmOdllDCya4
hdXrMleTqY/IhWO5njBKYcMzNl/UZpzLfj8Zu1gN9f7diC/W+xGpwrXMOL0RHjWp
9yS6gRSP5oNIeme1GTHVTFh0s/0Ql3v/cBo2VUvg6EuF27H5yoMPTQ8et9qkazNY
eifDvZhm3AqQydcb5ExLvtqQ/HLXJBDCEMwAj3LVbkbaWYcemaEEipd3f7unmhxx
dvNKBvU0lwA6cbpwCjMAixngiN3zJw0Acc/E+oFYoAjs1nnQHsakDlrj3Czvvbku
eL/o4DjOKo/xITJdQ/QdYys6IjwaDVeBnao9gBcJmJLoShNcg5Y89nXWMIUjH/WA
JHDtHOBXl2R+gviOpKucbIkJmufld3WTzDUczsLAMp+i8/8V4f0NQ/er2XAEPlUa
kWXuk1t4GwGfmxv4wrEYQuiT8dYtWbCW6/GmBak8YuKf1tVkepuuKl3hO4QjhDt7
sbNn3rCfiOtPYfHmN7DgCwXDBaVtEdvb8PdZXgvAPh87KdVZDzrynsb3bxxEzNE2
MbWwNsxb+IWiTxKpUdnVRpOzMbX+SopJZinFO+R2ULoQZodosHf3q6DckRScvK1Q
oI82F0Qsc+xpAIjKjUKAnYe5bpkTLC0xD2V44tQnA+8EmulVx/3eVJZZ/yAeUD+5
LoKfDR1UktZKduzIDGb4HrtsFhgbUj+U+od81LKCelIwhpFjuTy9XUN2dMyJ+unJ
ViIQrgFopORNaWSREquI0TaZuTQj71a+3+GG9dH2MV8HYWaBGmub8EYHINDxH665
120Y1/JRQmHXm/VNnuWDb2eFgWlqrR7GquGO7WCBjmIuC0gHiK5EuOK7RtimrP1R
WYZAI2H30Gb70YjGuBsfJV3EuGtAQT4LoKk9cAtiydHGT4drLU8fT7/XuxcBV0oV
byvAE7ONNWgt2mnjZUTJyJQNFma1MjIAwqdHooeVEUkfBQ2VPKaiT/+OhIQjzu/x
XNURJqFXlHmQtBLkyvyRHYfgwlk/joq+37Xe1uGWISSApirmOpPBjeADO22YBDTh
6rcrkj+0pQNCaBM8RH/Z4dUpPkWf4EAAnS+mYFhaSRqQ4JIboU0UEbebo2iijXW9
rqBd/jhiDkBivCTq/F5lvEhRXA3DncCLVpSEOruusrqmg0Z8rJkTWOo+nniRR9DZ
sFMZWPcFlLxznxw17F/CkCkGm6PsvuXdR27ontIbabpwDDukd6JVE0LfBOcbM+MM
DE9cl2PCamwkONE+A2odrorMiRCyWiAJqSt0KFhkx17hboeX5ZTcFG86JroRasq/
Q2eNBLiaZs7Af2RoicIDkhybgMNdUuNABTTXnf0NY03CVvrypcBvW2tayXgSVT+Z
vchNJjbWyVm/GlWaN1Dc5rEMKn4prLHZzbRBULdo6CTgazp2Vw7Pa6c568PrWRgk
pIiHtHwhXiK5dFqmtMFOivBE5hG/JNLGcy3Iki/p2SHXMOjvvAmHBNfPIpUXe6T4
J+AUEBQ3jYOJFjPTn85yiQ1oY3pJLUKsLjKf3LCm9lmEo9LouxjU4NrPssMn2iYo
Vsle83XIF4nI2lcTfWKnbHPl1AUec1e0N9mkSh+cgGS5D8/l5PSOG9Prx0lfvyJW
t8aaoWkftFWvbod2q/YhAWGe3G3LWeKwDF5vLIPR864t9mHMGqjuXBNw5tZDQuUb
kac+y+SdbaR/iQqm/32Hxeumg4H/QlkRW7FwiOe6NFQ5nMoZHavJcEzeGJudyqAK
dqnjSa7R45o9FLzYyOVfur/gtTFRmNbztD7alvzbODDuIbh7BwPuNBzLzcOgZK3u
Sz9ZVpI6pck5a9qMv5RzorriiVlAll3Wa+yaXzejMEZa8gJUSQvSdkZZr1mgvvKI
QRxVYieXyx4/cwbXQRZwXS/EOBOUb7qsWLWR5nj+TX9cHYDWkGrliZ/2guLL76a4
SToVDXrPhaczEL2ya7f/37LkHBHif60yFhMPT8YnJ4S6uZ/G/tYNcMbXs087gbpO
iCGBrDroao/IysWbwQ5cdbECETog/422a/Dx313HTzgYSvKVAMWzy7ogcAKVUql4
jOByPz/SOm+/4bJL00uOPY+DO7AdU1sazrRs/oSsqWV+KEVMkg5ffsf9C/KhWEhT
HrcS+ggxej+FQ3pIg4b6JioWob8l2wb4oK8Vjh+20ai0u5avdQd2M1C76bJOaO3T
2DKrq4+eHoGIZvl09Y2vMX1lSN0YE2wNx5ngpWuP+SEvnT/4uSaGlgZN6PSSrskr
jmMwTdd0EQW0QQc9TdqmP92MWuzsXod7vvP5lyas+6at0FB6ZmV4bhktEA9Gd9l6
ZwMHn71pGySKqxltolmSZ+baEhzSYnifUe+rv/xI73ZNG7rZesHGVfbeWCjOhMh5
ix6VoaAX8ImYdoVMApzD+TjmGckI2F21Q/DHBvoJXEuh0NoWElHzIme3RC9J8T67
CGk4DGBYjlycx/g/qN4Oa9wxtDTsRn3RYNSuzY6Hv7iNmbYhHzohRf2K/Qq2JFID
l47mGnaBqxtXOyAmojFzu9hxGdNmkk8BPZ0VWr5FPvYaI6Muq5cTZdTKn7d/KQVf
Dvi62/PBHOr/PGdKX5oHy8Ib9/vduy1wIGz9Fmb62GViSZaquFL6g6+hvBBEEwhX
e3j+bxxdbH9fqDowtRp9y6dGcbbrg5F7P/wbIwi/LgoZLwWpGPdGQsPYzb122MAY
QGHuN+H4mz/Zdr0E92wU2y/0cC+CHyScApX13fmSP2xZ0dfeKxLFOTrXT1pYrt/i
3kkVQiaq1hye2Igj5ji4LK5t2JWkst5o47nA5FPOrP/WTGYjIsPFlNb43gFn99hE
WcbC/Gy2y+LVgxbCV1bv7tNiUnipF+H+75AIDy082BC2HrMb9lvsVHcNa9dyBFgj
UG+1F9smfiJLpfF8ZddEf0EuM3QzpeoYkaETsc8WuSsGhCvgitQmRkZLl1S1AJAx
HG/M1NZnvX2XPqieuOL1RaiLQH/ZFknl4k9xFi912A2o+FDvwfjfl+KcqWuUwJVp
l0PMsveL9x3EFHiNeRmKncC+nCzXfRrgFN7HvttYXUN0SWxwxRe1WnvXJd6DOT6f
yliQaTFYmH7bqeo0+kLydUAb7zbk9XTa9bV4TnkB6VLqG3RjPb9MhEuA0bHhXh5s
AbxY6dnmaC7dn2PB2zuYdwinGV1xmiM75465dlYjlBk2+HLdKz45geyIqshDU2bU
zDIRaiiV/cAHDSCz55Rp0RzfbnBoaT3t+BPnZVTnyO0KMMz2enK88idIA67mjdh/
YjdTmyF1LtPGx1O3phNEKO1waWRqdGHLiLvplbOmLPGsQrZML65Aa3YEZi/u0w3t
0yxGxkbkn5ZFfTJxNPFeFdUz2rI3frZTeDbLeOc4GmocYIbJAsexxR+W9sXus5NB
rFHAwASTa/PfgtGXBJA8NWLMlXMhRuY+9NBnb0Gh/U08HFsNAwJnyuTCp/yRwirr
GO5JQwSJDU6Vwsb9nsi9Crq3JdwT3d+ND1ck6xRMPCWl4TspENLkC3GTNlXnwLTl
z7ScHtHKyTerBh9RfYSWGyT9+NS+dRpRVqzuTU0Jj+jojQzHBir992ywVJAKN2lU
k+e6xusGjZJ9h5TGPbwIISMZdIZtXNNs0hAbRQ4dzBrPmw9cuDU3PuD5b5aKTDOu
ae/fM6ae5qZTWo3BigWfOaQfkyUUk6eQwwu/n7LQrmszuN6snVPy4htr1czIpcoG
jydHyc86SFLtJ9P0wpZWVyaZsSfX5X6bHWmBGpeO/VmprAUEVRoVxghTVygXBfqN
Q5lv6gWc+hefiF7UA5bKJoh4dzjy5mQRXnoES19Wxrf5tjolrjfPGHKUBmASLTGb
75GuKEb2HtXv5qsK6JG+iv5+PHSIz6kdTZnNYmmEcHGi4Blw4784RThmlF0gqw8Z
iR+Qh0Mtr7monnle16YP3eFnFm/fJ5XG247vSHLDryd7Ey+V17WSYoW82bafqrH2
Z5PHUmDAlWkfGXfkUF8mypVmEPFaVohjvwiwUoyUS2ZjBeIY8tmTcubNO5N9IGty
Ka7NKTYeQ8cyiqiilq+sgN3e1Fc4ydkmL6jOsnKYdhnUQ34CYs10rePRMipMxrMl
RXjmb+88APEqIHTxx29FXGsKmWbnILRTOnP5K/BF/fqwk8IXGm0LNQbtwGoBTp4s
xlFfxN7szpjQTFce5cB1hNL7bNhzMIdsXEiQlaJD+QWRHqma5sLAB8fYiJiHuBuo
rKYvMflvKdJPHOYq/JcSx2RyEC5TAnc5RQQW66n7oPIxYOenNIsGKSgLUCJifXSN
ZQSMl1Kci4TisbxoCIje1n8TvrceNT41SpconverFKsVXRJ4hTAXKXkDWdjts6Yq
r+2QwBogbsntakyPFzrUvbJb+THpZ+0kTG9B28C06Tf+6rTH2sOMqEsEmICCAP90
e1FXT8HhXBiy4dW2npVYxXW9S3G0gXLY5nIpt69DlN8R6pY4j1gdIFUkQyIRfBkd
+90tESi6cFiY6qGkLiGxKO4sPewRf7dGKn3wC1OYU3pMiNra7Qnaa/3Ev+FPffXo
c/pI4KbSF3V08XtYGUD3gCO9ObnXM6ieiA9G173hMhTC8euEK5ipb3aZyCb8gbrF
1GdQVDGiGi95npg4xTGxOI6aIRF8wdPm1zq6rMYIczATBLtftAaQOxdOiDWwbty7
4Kjj/SPbpMYZB9GDU6OaHu6jmzaYaz8OqEhL01c/k1oPDpqOnQhF56N979gFPWQO
xMD0oFlCe3n0w7muPIPZZK6SiBwI/IpQqp5IGUXUwKc8taz4KA5XVzKBKbMBLN68
G9QjsL+rKzDXBC03QuY0JFL20MKEPO1pbkIiECbhTdBxcIUJKk8Z582ShGZvZYCb
PhCsKJYi4j8d4cXDMSCrXUBdbqDYnOo56/wTTVLbajWRT0l1M737bP3vrd++d4vQ
6AZEF0kGUu3/VRpPSRX00duY1ayucqMwQb/8omaZFyjTB5YNfwLCEjjrG3M/79WL
Awchj8RtWGfF5eTDyjaFMF1w2QdQPP+aHH5w6mG4o65dtK6pxOSG0kW27Ejqhquw
7AhyYJfMrUpo8I/o5JABUlDieOQtOfkHDe+0ga3UM6SY2ZLD6q68Z1Hq78J2PHS8
LRS2Q71ACeLdChDBIiMApsxr9X8ifENjNzLKCFWShcFW5kULhnGBrQI+7BIBIyPm
qrAfhy57C+PkdvPbu1jB3bm64cFmZ80ANcc7qSgzn5ZCu6FSliTNc6hn22f+zy7D
vnTBf/f1GOdRnUKc1fzqsdISxAuIYmX7ag2/w/140r85twZll+RWuPBXzIsnRLyC
aWWv/Bdbo2qLqH+BS0L+srbqGZa9s7HD5Xr4qohSFIXnTAMIN8inwwpPNBDfcSAx
GP03HAOkbevC4FSZ4vIC5fHezB4OhP5lmfHnVe6P8QPVgITcIsxY0TTh8DibSDCC
XcD4pwVyvigbPANG5UieMLvexQSO+MkmcdZPFfUJQWOgA9tlmyfK9j6bmk89lXsb
J4pTXDkRIIZEbmsR6W/yfgM9D/bVo7DzVT/3e3lOO5e/zYMAcxAs4/sBRwiWmjcY
u4ugtD83GbqJMjttvPkznojW7H8IHg+9Xl/lNoExNMLDRGAf8OCmNYDS+SQBqs14
hvpJlbiW+7To7VlmhWC8VLhzGN8xtSKVr8WBQwBeP1vK+1rtIYP8L8S5vYFIi46N
eZnkiEC7YYUrbbCBkuiLLyIWNy4VogImyfMI8RZPXbFz5Le2aLYkzKYfnsWB6D1M
U6vBo5+ettGlELFEDRYCPaam2S/mTIVxWmPIUcuFPkt83PaHvwyux+62k0sA9/PO
50mDEny1C4qF0k4Ve6QzoUM6Cwlv+ntzeX/bK0CLsCxNmdzadbdzGPegh8AvgC5X
2Y+eqqrprW5l3hA1fRvFtbfpUK9i/puUckNjv+ZTqIMlP2J0KkhsjuY9uZ36obEK
Y67lh9YDbFlUdpUhHk5CjD2NE2qo2KL15Cqy+BPxTPe+Luwgt2Pxx/vmjd4glvun
XNgWUBl7q95/NFr3yNnBu5HLucxIM/Ixm8xrDHsQ/S5/EWIjD3DXZkQTCAaXz9op
GS07x+q46YPBVzEhv+CvmK0TerMcr0vbgtIwq03Ax1LSQyHuafdyUw/DSJCNX4jT
q6UlakayloJ4weS8IdDtIetZDVv9olUBcoYhAaoT60hM8bzKhlCmj3QQsniJYNbD
1fKfn4F/2f4hnR+wCjuwip/rJLZcWbA85ngaF9GMxnooheSAjReLHK96cZmn8Exx
ho9dvQi8NSd7bNnoZSD0BrXcx31yzaBMomVUDmKCgoA8Ds4Q/4lrrNxrF7GcA4Pw
krOrQkMgIYKJsAgj1NDKRWSKfERpY/oXkNksWMs1A0ftBp4obWC8KHE/Qs5UhjZb
ulW7CPg5y7prCC8vzXm5DTwzu4jz2Oq/lXvIXxmEUowVXoX0cysF3usDi/jv5MNT
DJNnnrAo7vsW5C7uDcAU7Y94I5DPl+n9XuKJoVnpFq6iWKq414dKNexX3NIguhk5
87J4QZ2gi5QjzhN2/yTuwTXT8hst+QWG9umUnec2j5LYLJvVeh6fZ36EkDO4wMH9
WaE7CHEWMCY/SuoiRvZMleB9p53L7mCux0CJtNqS41R7dGZutGc7hKIF7KPT+VST
hW5A3qY4cIb3diPws16iua4MJHDT5QJzlU0u4TF1lD0Dpsi4rAGU0FaYcfB1XORL
DY2jWJqCDWcFPukdgiqBCj8GAJtPUX0zg6yiAky0nWElmaidyAAa4+wjcNP+Ulgw
dqtXmk39xIstqEzUmQmeDGXDfZ1sBwQBfP2jVQ2Se5WEbEQEq7wWrNHN0QfsOW3k
SiSZfKQxrKGXe5dgxBsGDuOWyoXb+lEe54b2jtoRarZ4P2n832g5HIvcEYpKV+Wr
CX3etGPbdwVzgmC7KyXSLIcZRBJNRt7TKeo+MIxzDAIwt8xgCuz4554qpKr4Lu+7
R8bd9HDxV/HL9MSENBIe6VmmjCfbl67/5ScAGgJKnd/Q7u45nHdy04q3IIUSBum8
LlMKrc4lEi7q1nYHyCpiRwSaxWkdeVDX7s2UdXIHEDrdQJl9vPeswh0zzFnsGVww
NEVCwL/ILKnTRdvscDwuuaAcrBxSH1sStBtnVWJvOI0IMXcMDilEpTvTKl/7eEPj
N45SeDqkRXHd0U48h82QWIxW4oz5HSfK7t+8DdKHLn/bosBSX5VgGoGTbKnrM5c4
KPQwXC94IxPOuFV0R2+kDCVZH7QvvZyq7xyu5yN9LMcNUrD4A4E+8D23xm7ulpU+
hQ0AjigDHLl6arJwooFa3pg0dnRbIn9wBJ6XFR6PO03v8YiQMDjT1rWgP1ooFpYO
U0RROIgAgCmCn+uJydxFbEFu6kfOUJHKT8yZ8YIS6NPibHuf5QvW5LB3IsiE5dx5
gxqPEdF+LoGBY/+5PWSC1FfTyoD2eyfG7Ypv2csG4jYWcUWs2L/Gr5Gf0m7c4ak0
7mRxGcgZbhc76O2mPrE9p+iAEtT+OmB+AXzlDXhh9Dnm/xC6+rf1Jvm+rm6Z3S6p
SgEw1X4P6x1cN+cRgZd8qGdHBTHB1rcidKyZO175QpupxVdXPqivkELsr3xsyflX
qYs/S/5P06f2QMnSVv+Kzk7b1M36JT4ZYdp19/uh+PpUZafEz7XnDLfztyixdt9r
E0Yntlz5PmpjiWdkoV+iKs4HcfXXAh+5mYnfjUNRCANfCdgJJYQOteuGXr7XCWYA
cXI8D37EhLSbkwAJtSMiefolDA1DTW8QezP1TTcSMwrD+MBDjGD99nVUrskb+r9S
mj8CjacXtHLTs/8vBvYH7I+uq9MWK9QckP778q4vYLXw35c+PBPFuQkwIgbG6Ear
937DEJNJzCR/U9uMzQDfT4DkBh78vnVwmHFW+ooraXowj7kmY+bSsq8T4wkOUabZ
1Z/l1VnpUx9vl8x1Z5tNaExo401azoYamSPQTjWB3wLAF7dTOBJvK/DFiQex/Hcn
kyYnLOwMFosEkQL5REPRujXuvY5PruIygKRZjrEg9nzvssLYBKMlECxrF/24+5N8
MRscQy2y9YEcrof3ENDDSdVEjGB/c2JdESsUGShxOKIHsZ9qg6wqVQ69SxsqEcWc
z6HDf/K9RYR1iOxzl0LXyuCkWciI5yzS7itXifPEnq8i0Vfsyl/czW3k7fnhOj8t
Y8MVnpDNuVHL+tYZUCGHx56gcuWNHj4H3AQCX3E6H0Uci6UK+mkt0uJ8duLb6Zaw
dB5JJ8nB5tGKrf/AFCHHpAZd6DXKdRvsRFTjx4ohuQvDnThhPE6WKcKLcFa3RlJu
MFex5J/Am1Me2erGPuZn/75xjXe53QFU/wWYQZS+srsH4R6Yf2ROKFDwlIY1YkZu
+OV0yXxdZVr5F3zXjgG+dix4kll47wvVwlbgN+yBR1RE841nOp7/Aelfb91tj0ku
3chi4pqondya0fRF1E7VN8cHkrBDG/Mk2xAWoEnh+Mc2Hm/UyYURTYuhQiUIaBQq
efhSUTMM8FgVYDrQdlrpJhwZCDCsROSpRMUfBCsUZHu5rNsx9+ABUyXWUVeClipn
AR1OGac+Wo4hBQ9m1AX23dWqNgHJeFxDodfc0DoOWp9O6Ubz7neQwD/nwL4BuKeF
eAPLE78RbJxGMCNTkwcTHUqJeJMN6PBqfyIwHfTf9FMsrJfcjpBoUqF1muoTMIxD
rURgosppWaoBRPtSJvQgzjK67kCFnSWvzY1fgY3r9o2exsHhwP3ootVRWD7az0Hh
jiDrHL+99rId2CMxyTiJTkHOhZLBTnKdl+otbb0hC/3E8QFE2wiucGcZXyqkPzh5
S4Us4KkiY+miCBjLjwteyuGtb2mjLA4hRCjK3T+jlChmkZauM0TimoEtvB3Qq8Ia
r6UXiTg0XrrOWFYoDXEaauNg5LsrvddRY2AkowFHklLr+1uBt8WyEDWiO7h01013
qb9S6RRgT+Qiwkbx1fLjzLsykdqT3R875h0zx3OLbHoUP2WTblssZVWIErJC2MZw
cRQmcaopJy/QbjOvMg4BshmuqCmX7PYqClkpP0OskcPGi7XfUsw39ZUJ5UNZMsjm
cMHz0dVJrx3NbNF6PIMPJTAr2iiWCE1U1LcZNv0Gx1tfVl6WUBthYTUWSrZzkq2q
76q3AXm+ZJ95qprIB1T3hwWDST0cs6QuKEuaccCdIbfuc90WyIx5SQvu5/ipb0Nz
Ng6sS/tH0oW3P/mtMq8YMo+gXoV/yLrnz7xFTLeWe88T09oaPEuDmELlGhJsGp5y
Nwc+FgqCKHyMuCzXIl1OBgunNQKyrQAsOOZoicILLTIhIRiNg/XE0w6p+L46oGKf
RdoVkmWoZUiruuAny0MwTUhZv2GIcgj7meuxi7LC+0gfcMWYLjc0eVjTQjgKBo/3
SgWwWlGbgqrJQ2YgfrhAXWLo8PgYNF3TVXzW0v+Y6EhdgdhFv6WrxuFESvhKyHBn
Cnwxu6c/ujrIsoE1ATMvEAp0qguEgr7w56xdwUqgKciJPtrkCDXiu4Qt1/IzOG8o
1LKH6A/pyQ0OwYWRYVIX+k1gFd7GMvOfru0lZxUUfFP7b+mfyRplRWbrUJdzxBaX
ekTswm27YCCScYlL5W1R6FE55gnZV/7Bfi08Y/10YjmA3uHoAG3luT9DQ27Ol8UN
QLVveWQD4IhEwaugo1UsznVq1bNFlHnxm2H7l4jZBGENjQ3fMSU1y66mjV4K9UM2
PzrJ1qrukmNoHCJtmyU3istCowR2nmyrxWCvU1nPiNhKwglYt+UeSvuBfPEHoXHR
9+TrtPmqkrYlc3v7NAHtBts7ToGFFxDXCUTCKwiRnkXc7wHY5LWREyPemdqVWQTD
j58fuYAI9bB6UeCJck07UagkwHK+1NEjtamVAEIIlBCrCYPvYsUn2rs1hCeSspRA
EHCWXTcbao5oEwibAoowI1Zgv3XhibEZ8EJdK58812Qop56LEuMv2F3i9lVhOPN3
CgeqmajC+3dNUJmaFqAVH6TpSPaCZ9radFpWmomdUipvV9r6CePWmhQiJwpHryuS
POg4qcFxRweihjB5xP0zRCYUFIqoMkXQD9DX8ruLmFoVrZQc0uUxZ3L+odUFAKPR
w9vqcCnLw39iIci5U4kuB8+mU9bLlitFv/W226fkupTPxz1M9T3FF4b4JjQbeuha
lENkCDcPRVXKAEGj7uh8t194jRRUvXgSY5FVShxVDs8qXNx/vwdvAX4Nvu5DfLaK
we8ivnyxALdLfZSr3s2W2oqvJUy8kuJaVKlsiYZUB9HlmJm+q9Us5c6v2peCPByX
GC2X4ghvKdo9pXVG4FuOQKwh2fi2VgUVAI22i+qEKaOUnj+OWb2IpFVGx3ATzCnf
8ukv/GMNxmyuK3qCNCihHUFbXGDne3VG+bqr3DXwej6CDScNQtPUAbImF3zgZikt
MGAdimrD9vIV0XjvUOmAfqGfGIjDF2tEUySy07AIJagaFRnwznrC0PU1IUb91Q1x
78QufO2rf1Xkzegr6i9ZgUnwezbtPyjGtNpZu2J6ijeI0ETQoj1R12AxX9JiNc4i
j4/VxRRASVb3fkYsf37edPGdFopVL4TjtFqBeMlZ1odJKZssMOuZC4W8hEiqjBry
zhxwSdVUT3OmXj6uwEJQbQECJJQn3qm2QTQGP5UDvCPowqKWZV+zHY4Fh52KBsgz
ooKVKx0+8/1ltXhqeM2TrVEvUsQeJYBgcIG9+PlFxecjj3/lDtVodurNR0M4hPju
KdBoGzHzLLxqUnIxRGnKHx8nsnCYE9ynESCw7USfx8yDKbyw0A1JMCgUDZRTyoGA
TII3pLxKa5frZLPmgWcKTDeq4E0LfBI4kOlDkO8gkDptYT0iktgxyNZt2kfbJwIK
UX2SJZ4MSo6hSZ5LgoIQywK/3m88hF8CwA69UlM8ayCjuy1eq6Q1BC0Q18ETAaW7
jKq0+/d/av2lD0mYJpr65SEWlXwk0CScgOocDH/2E0RTQppi7uM1APzRVC+ikPbD
eW+0O1qWoUchvz4VCgKXVYrGln7ReuM556y8Mm8+YdK5a1bb0+WrQWBLY0qBhafQ
84hLTgAIEYczYOs3VGL5cMIrFs5/ORVOoBpVMslS87aziIyDbPrTJKd4zjrUKaOh
zUdf/pfh/sOiCm26S2BGZCSqUdHRK/+pU1MKusUkSADCIKNzb50xu50A0TJTwry3
oFDszjuculN+tFriLXU5Px/osDDqLPH2pBHe+aI8W8bjes0OqIKXyu/+Zj7Bfxrk
MDBGmfQU99pElcjVoqnNlb/XWRlrA0uXbJj1ogIAbkIEB4SJEJcF18WZzkvgEsGv
ErI9aNucsECV+qWyCZG2d/nmYR1XqSloliQoRF3hGkqzQFunKuUA8DDSarz752zE
otN58FUzCnatnoPQNBZzAmJlAAs+Oju8esLDz08xAODzzbOdb7nhvTBpWUOem+rq
D3kALq3n7M1EyaVTY01/wZUI/vADK3iqHFNbBg2mQbFbcipdfZqUcvWwck2eIH22
kuyDWsIUaRezNTcKuIDkYb3OTLkQOD+dcqP4LdmOshs4qAvadBIHRCJ3ywc4R5dj
Lx6GjscgKJPouKzcHSgYXFc9GqF2d+ESVnVVScHoy1kHPGdS5uvKbD8GZ8m/2lnd
EP+l8HoBXQ4KFz8xVbSc9NjJ7LGKlIBJgVahDYw2L67foYHZe9C6vTVCSlIOIesr
Qq0xojI4Q4JyK5GrVVhgEOOb3uWG5gteNozzwUhFBOT42R1hibOeT5x/x2Xz4EEW
ARma6hg1eJ1A0xKDS2WFHxgeinvk00+zmr6dQa9dIc/fAxHt7TXxtUDvEAow9WPs
SgMgO+uLrJz5sCVicV0xJ0eZ3iGYY/EJIPY731cgFBUxvdzJeNK+CZCKh2NmH+wA
xOQ12QLFX0MF/hy+yM2Z/SE9u0XGa1J1ZzCWdnYLW7zM5aSy2x03w4vhxCG2Zbjb
JIzM5Pv2y5z2DDrx+iLp8vkT7pTBG4wskb3E12gvhlrUYDu+e+8dPSFKwteEeVuR
5VZbmKSTuPMnAQ714aCjMmRbttNUZG7MZWKqSgZdWPaJWLZmBB9Q6ZCgAUXV90Jz
q+AvXbEF62l0dGTReV1BVnA1G7iM9Iuagr3Q7JS3Fo686Pn+z1f0guwTFvzFVOwV
WMJl+AE6+V1p1kzcjyvc3anixBy26L0minrgKTM4kADOB/TPohfv0vFR7vnKLxuN
Rk4MS9CjWPMmW4/GSf+xJjQgaWwk0qSBR84hXCzTmUSv+U/C7Ptzp09qYvSesrcp
oXfHP6ioOpjnZA+F2kO+zB83cZYyibxSY9fvAVTuO6T8vDG9RxUADGKtL17SYSuK
vD0uYJBJLzzVGSxz02/Dn35+LoOnZ3/lR1EWa7Pgk/j6M72lug3mRgGeRj1gV3OV
sxO2XbDdYM54ixyfFq5VBWldtQVcVOvMxHMOW4hMuAVPfE5ZzBlg2gylSJ+61g5j
QjZuZdrsQ4XcxKkClASReqeIhHTEOzH3VOoKTc4uJt2R13LD6ImjCL168l2ACaAi
5pU69uAfr/jBFo5bj03cEuPSONnx0J4dTUbjBvopZeI4IHMyZBfTOVAImRiI1lzt
S9EmbvOW6/2sMrb8CDTNJgzUX5u5DfHI6/QogC7tC8b59KNwQrSx2jTVR/j9Gp6W
I0PBJpAao0vxofYokXAKw/+ejrRHDnUds1LpNN+ey13PCa00sRK0reoBCzwMhWf0
imVI8Q5aC+nXiezeD90Lc2pY+8gItBLjPOHuMCbby0xTPXq4Hdhu3xeG3+Ov97Rz
EQRNdl+zBxp+V1K86ylT2P5YhEe6N/bd37c5Z0JN5qsXTyZbHhXiLT65l6O2duR5
H8ETSjLq2Mc5soYphITWFw798Z/fb4MQFSL9z1gZoPLh4hKDaDo5qF4VV0k9YSAh
r5bn45GbhFZrDqrmF0t4wWElPfvtfp063VrOfTRk+emvFzEuF0FO6Ec6OC/775Dh
fCqIc0J31vVK2/oNRIlSfw3rQNl8brYY+fR87M/SyJoXVx0e5WJEU8Gk6HwY0LOk
RF4mpsgQv5DoAAQaumxkz+R+/ERlygsvgnotBvNaTRiLrp7kSBu59poCQ+gfOx4C
CheONjvwVZHJC7784kvrEUbAMzeFwhPx4nclTalMt3FCo6pWpj0Ru6G293ZGtiOX
d77spAMiKOq15Qy0QZgo266a2kso7qQjqoAfpdBACc0lCpJEcMf57FIwDzkoPKuK
mGPJuw7eN7u5+3ft5TtrhedTxb7cBnRWArzjxfCweYYU45V1/lGnKKPSZRUzWhDx
chky74qXZ4EQmwgJeMmLUDSVeMYBONg9oZLszCZrI6W13Zp1jSom/JZCTeD+CAb/
cNdYwbvzHTiCRIdiULEEdPz8tPKx9FiGs7W8SW+nesQEPNnRIMe1WY8sat+r+EQZ
cZqpRJzVrHnZx0fz63jS/iOMY3J8KyWOaubkqxWk/dMUATp7eicSUXHARc8PacFU
NDiy3Kk3TaebzJOSQHNDabi7I0k2h8RJ3SGhhFEHkHpc3nfDpgoXtgF3Ov9m7OUG
stg8Vyi5jdFsV03m+9ZNy1XSzGpdsDDI3YWHotqKXmBKjZrHMf74Rh27r6wlmW7w
yeyVPsklPDdE6EzKYtLJoQ5pBgtP0uL9I+b6tbXjB4qtmreIHmPOi3H2Hwxqg3YR
Mc+Vj5bsArHMTqkUaU4mSaRiH905Ga+qQdJQ4z3A5iTX7ucyltgJNMPT+Oy9XMN5
I1vOe9K6p5ie5EUPiohnwh1gj8PWwgvWNBwtvOf5cPGw0eDcjq8clExMZdqG+pBW
SkfcQCB7kxHJ0JO37ybkL6xveDtzm/YEKYA1nZz5HsN/2xTxyMLItYhawm81ujSL
yl9KmcDsddWy5kyBIGZ4MYHSM3ETImw0RVjx4OJ6dr2+SZ7c/eAH1fAS4vuJ4v5y
Q74FA54d59qch9Arut8tsfZEpusyDA/Xq7qwd4LJJrHLD1IXrCH3QY40/7bFs918
kmI/4pr+03fELTQKDiMh43gFBk/v9/0+cnSFlJa2jpVF7iTfsnL7utOBG0dsZC1v
MZvVq3mWS1L+SrZgwJjMWIZb/WgJIt/VWKjbGxVKelkw1RUR63HTuynhA2iN4EkO
1bS7lXhOTLG+bqnwl81NilTeyY8ViGPV2yXDkp0/uGo6Ogaog9x0cLEb5d+c1VqB
Td+H0XRVCDLkl6XNgboF4n0yZuYZ1xxSo3/BjHs8cePGeBlJXOwIcdb4iIrcCAf8
kG742y6DsLfPwDXwjxvdYWCICFKcEoyceTZEOttohcgUIojweHuzDFCohs8csfpo
9l77/i1PL8z+I/4C78+ERvZNn8MjtycJVEA71Wn3Cox7KnlNI0CIt4YaQhON0raZ
m26xCQ+WOP+r9TkYYVYvPG99CHVJNBZjBw2hlx/KIkETKTjphj+qEVPN2tMB1JuH
hMvYDXYh2IKnQCjmbXiL+P8Ek5MQIF5E1mqewtkcAbLrmFhjB3fSQOgrABCNp8Oq
zWJNykFYNGxKirPcD2EeJ1SFXtdoerWVaqIW0FixU1vdVzG6F3Vnmn3C0trtEa3E
5q+2d8Vs25clamCtC62+mBOyf7H9AMpn5vkvkml7Jz27ZBpDsPo35+BIXuyMM2QC
sncAMaPzSoL9RJ3mldMV7L+6sXxQ+tixXko1lRzkTkARPtfUcYuCm/WGm2v+S7E8
d11fh69PAgCiIVPFV5dRtD3bg7WJjEqTAN6e3dRku22Q8fomNg4K5p2rBtP3/yhT
ZAhwRVivjSGVympZ1XBDeA2DA++zFv7i/AXBdBBIh2s/6NPeTi2ZnDnjMIlGAOrq
d5DOGVYb9dXbKgXuE7XGtu/huT7hT7rX/GoQw+OZV9TEae/7EEXQ02Ks3PyaDHzG
4y5wBhwIFKgQoNGWXDFCq0P3Ef+YgWbutPJ3fIwGXJoSkg5VDyZ4eGAscR5NMK8r
UrT3SRXCnDqT4idwMjdWO/wkGVdpgDLLEiHddIsxPj0ZRv/wJXFBbJkauiIf8oE9
wQoATQW6canIQYCHSgZ7ENVGTGbEBHzsohiloK+dQIhvW/xYA0beEgDOr8bvvJuu
0w+wrUe4nt1nBJt3U4rR20lFM0vf+1dLtLeUzzpc3nKuzYpQY+0vlrRdYMbMWUV5
kjTbp+1gVwdyh1T1UwRbTGbdGqdw+upf95SawQp08zAC1TGv0iahg/VMqGB4dBzH
cxE7pFMB8PY9ImK0Riri3Dpw423otVxJ5TzLqNCUEoRyV8Gn6Cu+9IfnfS4aDq1S
auUa9mLMsnmAJFsRPR6x7I+cya7tfo9cjT9ZBZW42tAHanQHa/5bTVzqPbpl7Dy9
NKEmKpQei4NiiqrWOxF/QmmA4Eimo2SYEnECJAF4qKCkHhQfqFNluHoBOemgWmAo
axjSF5NPogQxUfV/DsjRgS6hHhlQgV/283q5ha6cIgP9US2P/8xlywCXSg+bWc3o
3+A+TbUwrCOS05g7AHlMw9HxbEFJa8wDKIi+lpsedUSHaA2ULabyxKAVSL7lOEpk
6kvc/uRUSlq60xTHCdxHnXQdKZ5HYyFVve43SUkPy0e0BhEhWWeMW0hoTZ6d3L0x
g6J+2ikt/w1SNeFQgGO4ZGSQAL4eKb2onQNEwtl5L1WPyi47/LS3O2MJINS/mb6E
dRhPEYnGeZRCeO6xXNFy7shktp7BwnCPdWcKoWgGUOix/xfpl9QwWTQ22UEID5Ih
TalJgA/djZOY4zXPYu5voDpSsU2yfujOAoBfaG0q81vJHw/ris2rcHCVuG+bx7b6
v/SycxVkZML7s7xdI3iGCtHDgrUDoXpUtScN5fB2wi2KOCB7ouBLioN9xAZaGnXs
V35o69WEopcoOtWkBg2uIeFeHGdwqKPhsriF9cf6UomOmzldcr/ll+sOfgeDMtfD
qmiQ3Tb9MgaPTChHB72kIMurhROtKTwG5VqpjAXboDvwDTCpimCtPoMaqzoWOK/a
B3Qj+vrSAudxUHdyJgvPTNAHngkUW9IAmTbnvzKXBEToW5Yyr9DJmt+lqY0ByCwH
L5uM6bGZWEIQS9Uh79bKASokRNj/CEU/vWtGrr5ul1CLs66WjuodFL3ElJcCFhWY
iocxhoaiaam1RXiejk26Y4skWihtvcUCj1r+uuQifJyExjnKLwjOzq5F/xQPlVAT
fbRRL6Am4xuoNlZCjTjza0Ty/EqpiqaobdyPGyCicEB8le9zUihJmz7lSHguiYgI
dWSq9f0LQkxLmgg4bPQuHeE8ogZwIJ2WrF0FA616VSEbVKXjQUHgu8V2gXHLp5uU
g5jjPLeX6UgHvfxdIDVsEbbQME5GQhjMtuoTLOIZFJP5b8rVTmSb0F6dwSnlb4ml
OpmPtRr5+0EnNqi6bDMg4xgzUq1CpJCHnUaEq7HQ6h/YG349aS8/Wo2OV8aM6v/F
rgVnjvJJ8HSUpqb7fOm0TkQy73Yy82VR5oRJ74/I8aFf638qRz/6UVRatl1fJYv7
Ux0ETYgkqvM4UxXnw0D8qEUkrsXZmgklFRtCj0ks1E/SP2mL1owp1LtB3nMxHHcI
TM4Qib8G6qLXooY9nRWRz6FXqU3OZlTDwHblGLTsN9chbPiuL/SyIjQgOd3D+3I/
bmTz/Xfe/27QAxn9c9QmqLmGqBWspIrqConn3+DpjUULaaj19nSX6MefEljKu+YC
/zjlh4+XQj4BtifO+eAN/zLss9iDV5ET4a0mtusl33dm7CXVertQ2rKGVxgt00wx
CzokSp/fY/n8OrHZu7jd4TsCRiq6pE5oRxTgW1bY8o0kIh42I9HycysOORIL+ynK
8dgD9TA1JHZH0gX84nU2jsxHcfFqOCNnMzRXEk7q50mroFEe9Qm01ySlc81qwUwE
AU9UUyEbgh2et2Gni6Eh3lHvf758EkSTEfkRm0WGSxbpCtsPohgbwSp87a3BiEbT
jkTiDxF5pmcmjGxjQNRZt0MDR3h39ZYlpZqmkliP4i2jRMlfGVQUeWSSCUTMdNv8
dk1LcjKVnOR+M7LXyLlKRP/H/JYjx6s2imcECCdnlvu/sdJGhCiicNGiXwRD6jm9
GOhbF4AF2PiARv1P3iymewSUMYpwWZ7A6atcUTTJ7AUwpolt/n2rx5oGoufp4L9D
zB5t1XbBXcH56xWmTaPwUy/FF+Q2cMIrFUXj82xVH5ZN/4ee2VNj7Rk5bqLXZ7ME
K4dcy/3R1fkOkF7/xZsZsrcAC+q/lmNB6rTkyMjFdRpyKV/W3GMlJW+Lp7Js0GZk
vewgk6RoHuhsjOCxbGs6N3Tnt0X2kAfrXAh9GXWJBXC/KV119Rlird5f9m+B5tD6
DdFgjFukrSZ0urBAX+GRgOISVhlwxWyBphhGbTSi0AdpVV64el5Q0Jtgv+kwpqWC
/mZIgYvI5BuovTyeF1MGqofowsCSfMgKlaYWb9ajZqOQwmAkH0F+qiUG6MCt51U7
jEwA25d0oj6RGVNqrxDAduWnpOePkFZONwZYR8xja0Dq68MmxIs5QMQEWBi5lQCa
TX7azYEryVu6TXDzOVTD4F/SZda8f1+e7S9Pd0NIKJ471SjefXPXrrWOUdwayG8e
jgPYWhTrKqFMa8xGhPN+qDgyqtdytTc4BMpmaGECHb3d3UZqThKq73G4WtmHlc5F
7cJlTHU0JlQ4LQTGODVMSIkOnLAu0ZUYNft/VCwMaoempTP5awWG3jLDb3T4UQox
aa37c+R4bOyDq3guZeXuDh8Z9Y9f8pji4vw324Z/oMU3wQ0xPVyNoBClPQuydACn
p1bTNeUoRdB3qpv1ED9YI9LNbtX1EB4H278s8+m0LFuq3xjCMYLk576RGurnBhJ+
cuJvjGShsvBPor4h3Sy+hTI/AzoC8ckGbKMtargP+w3QTWRu3WZ5PXIiRC3xcKoi
7HT626iXqPk1b+mDC4EjJtseiX7qiPLcNKx/pOL39hdk2Z5tjPKVDkOkrUXdiakb
VNPyBuE0y3NnLvfecMFwm24YyGWgRpbFzdQxWsPeu/HfXfVNabdxNo8Yhe9RXbnr
rAOhQtjwp+kBBVfP66UmHCXTkayezB93dwD1GSbZzN71I27PJxXTJMtHSf5lzTPM
Fg6sxdapfwPqW1HxCc3tE8oaLuly9DCzyc+A+2GaUmvNmlBZ5Qv4rqakMAboOR1N
jYrvPRqAdJZFFq5uzza5uHZItiiFJOlrSs4iqVK7KNqTEVObpmIJK24FJiXz724y
ir14dXwp1xmUNXfYwql63x/pGvKhMYD1lNu8wKSPK2FETz4WPHXot+CjlAHJdZ3P
NtF49TxlP7E5zC5+fQF6ne30RPtyhiivTTIftheVM7vy8rgLMhPVpr2AqSiPevx9
vjzkrB05wmpsjSPziZ49/kbYc0w9lXWynPZqmOSuNHbz1q8RG5XyucFvKBaJJFvw
7WEQ4ojEdsV98/olQn3lNSk+1oUUJGaD9fSlUgpoNlDoDzRqGrSGciokl3AzLpc0
g4wyEAPV5JEW1dr8QQqbM1In9AjFvQHkGj4fB9Ngkz41SBR/4LTJsmNQNX9IhcKo
aiB86U2DOv/+S8Qq7cEJf/pxuTsx2ZtgS7mRbT/km/Xhm6dnocaa/8bzQHFeCNvl
TKbpC2po5q/vA2qeY1/CkIh+t+wKvTxez5YVUP+f2dy8ahOy9rB7ED0W6Ig2FdrD
0VxthEe64OVQDHTPM/SjdrX78mMBmqbNOgK4MzfTug5TVtiOTe1kmCHvYKpHlFH1
YHLKUAEs7eCYOkzxOP3w2+UdIFGg8BI9UNGDv9r4NTEhzf36XGVDU/OZnAGUZKYM
WvwmbC2GpQNWUfqBnb1wwEbgP64kqdLlKwKISGRdZkuBaytUT8eNwokpSJAdMHxA
4LrgVxoDFuiGAjJTuAfBWzVo5eL22atXn/vaoxCBd6Ou10CFYiQvCp8sJ9lbhF2W
HRe5sEGGHPTtJFwLPqlrUxqpCApjMEGJYVW+Vs1+HZ84rmQQXcv36yKFuluBmHKt
onDfM5SSNywQg8ExP15AB0KbGCXMf+zRC01PidEawqndnG0KPglFkKQJcPQlnf3a
BuWqwg0bOknbmkT3dlNQuznsyvAbwqjMN0s9HjKmI//vovKHnnZaVqFiBPzRfrSe
KMe5Q5TO2jwLgzFOI3M4qBi2B0+2/4LTidBGoe+8Sjm1ePvj3linReb21d1OziCQ
1WkEfSJLvrpctyz9wNw0OSFerngBZLVqirAblx+9L4eW2JPNHqDBwN5dwCLCywfy
Hwcl+lhbk0be9/V/mHVQrDhSEcPF4J5U+lhJT8uLms73VTpzcV6wv8cK8TBqnG4Q
tT19ddvVsXQya3/eKMHJtGfaZnzqet+D8oVW7/o/Jo9Vj3HAc3XPcMlAkGp/FrAF
L1YX5B/qwmRojDCqxuy0XV6241cReqFW8Fsuuq6VVSCEvxLEm2JeQgFIIlXfDSey
WoTdof6lAcc5CVQWYiWoUrdrEplnQwzoBjBDV0qbXnkBzRGzI3x21qXa6T15xfwI
26TFtDchu9T0ALhDgoN+wf6IE3wvukYpLP8w+1lodL4g5zlKWezpCP0fQXr18yxk
eA4thRRtv2C8aplCL+YXuBTIByoRTv0MQXMfJJhDf7lHL7BwiLOQB3jvQIg0vJTH
CtYOeuxxeZdEdGnzYkHRohI9zyLMr377B4faWcvx1ig/cmanKXBG9p6kaXjxYF8w
7xfqqCp+ldth7rWPco6tatFGB4+ec3/gLhNqcYsJ/vfkTag5wBaiv2C2ksdp7Fya
HSf2YTJZ/qO0nTQsutFw0UR4EUKVS8pJRytC73c32isLM5u06zBRdu6Nbs12Rc2M
+f3SHXVpEOHDCOsW3AbRB+HobFhgxe5F9xUJVypg+JZEidHOFeZsyBxVrAB8go1d
IQeKR4qCsjiYVYK9Wc/Z1Yu1AchUjkqLTcM6aBc7MgY11MCLkz06QzCVuLIpAFKf
gas737CbGn0WE56tMZDRpiDE4uJj6tNFr/2UOIZ31ntP9L+GZixGL0FHFs4q/9sI
6FDeXM7nwRWxQqoSkhbxX+KirORYuHXxmbvrrMZSz5Ao5sHZ/Eqc8T/16t914fbe
4RJKsp/H9dEPzFNjSewcyXWdHwAmB7BjlBKF/Zo4A+D95RB1QZAPwEXDJhKkS9ur
o89k9x8G1uLwGjRjiGx8RCTSV45+OkdKo4MlrwbPlEQuE9G+Unc8pno+KkQGUiOb
sgCLua8ycEnOoL1pcqI31sY3M6WqVv4Pkgky9+Az48XCkO/Inzl3lBRitY2oyU3E
iBbLIjUBsob2Q2FTsW7Xs0DhLsKo+lv3hO7PguYpZhvZJyFIJ1PbN5ZS3y9U0kIY
2Pvm5Ld5KEDjlX5f10Gh6yD/PDyIQ0nOJztHo1aDuvgjaUb900QjI6+LrdZPKFCt
uH2J/GCwUjSnArDXeEz8rO6o8bbRS9T77DDJ0PXEaGOJluwRWG0rhv5Lhd/1OJ8S
fK+nnGSVGrHEgXNZyqnkMm3WKw9i5sQrESNA/a3idunL3VCoGXEMIblcPkT3LoiE
Kr5k26z3xGKgRUuBtVqlbz7QliKwoptag84ZVQNj+O6T5Ia/7TonjS9/LM7GbZHb
lwtU3nAFs/QdnwUB/gvWt9pRCQAqcXgOh5xog7Y3QYXhHFyL+FiP1d2NYY9efs6D
/42KKyrlUs0VrCcyeZ1O0/rhEzk6r+syemLVmUL20F1NyAVS8FdNNBpomz+gRY2Q
W3aDPuFgwdmuyRYgjiJT81FwM0SGlPK85YXyr7KOAVbPGyd4N+gRqXhVUtJIMV/0
yM5FTYgCnGqboPs19IPEiqugqargZ0AiEIjgAw9Zdz2z0jVbESIKSxMjrBpzvX8+
H+cZOQeUk2inwXkZMhqg4pIAbO8fYfbObvv2VYigI5ZWbd83IroQ5yTj86YObeGg
Yp3Zhp+tcuvuHzZiQYmVgjvO/FSVAmZtq21e7gj3unAD/Nq89Hb8o9kM/kL+Nzdn
9CuJ9IRdoqMObAPCFVMR2iRJxYIyh55SHHur1mWs3bwuanlGhvJR6DTawBRBo6U6
DhCt6nQvPRv1xCaMAxbEsQIrEKG5vNAf2emQiZboZUxPVis3Z81+XwmeUj1AifOU
RZQQfyml52Ftrd0GhqQh1oD4loIj4i/l8DoQ7HowA7xUp41eP5X6FnucFrXbrmMR
0iOqA6gyyY6wICPOR1r7lzhpIdtlA+rEU7ghr+1z2DIRbp7jvUlb5YAHK99Rnx3e
Rf3wJ4zH2bWh6IDtMvsd4SSekrexZuxSPLhmYhRpxFLySNPj6jlwrI/s4dKxMuod
VvVzZxI/sPWJ3jnK/8KtEcM4q1Mqd9F4Ncyt07RYz/yOZLxMhiKTn+4djb04VtTL
zrxV2igLWPnFAI3gszVaI1UIBXEWtGM+RWFlq/uton0LQ8VT3qyrnDgoPwhmSYI1
w4kFn95HuL05rcDFw9mUG8+RQHyv6ubP6CarfBlQOzWs0ZdX2TwAXVGDOzjSkXee
11O7JEM4laL21Br8nenvBylvWqQB+uEcwVdcjaROmUILHIQqDqTE5VrLkYfVB5CT
j6I0t65xxsBnvJQtUf0T7Oa7r3FHc7DJ9okcxizZuaBbtFIJs015QZJBgXfPAqwu
pSHrZlvw98KgjNwTp972L/uL7KNpPs9KDN5r8PnT/3OmSCJwMVoGfUSfXFYGiuLt
Jlli4leAuRqQvUIryg1LoQdYBWCEbS683/MegcwSOh8opAnMxmsV0/FwV7igS0Z0
YauqpQtYku831+XoL2I4SkPynSKbqTeBCKv+dPr6Xgokx/qkjIMrp6G56xdOi/hB
RnvNErc7UFBnEZNMk/PXubsD3TnUay+JstQeq113W5os9E34ZJoPuSvbo01CsyFa
DA4XCaRqtiMijwGb5x+EWlueUaF/WbBe3IWPQGcQ9pitUkE/3robjFsyp85ak/I6
pcfQn57kzr4b4clEwNxM7FuNXrN82yxoPvlPZHzdrJzdkxH6ZavdUol9emSopuUd
LG6DQcFT5H6JMmeBVRVR6tz3nOQkjY4GkjygbPL8W+3UgoGDPTBsuJHToNI/7cZI
Bif70+ec5ysjhqeRsWbnsa3j/nArrWo+gZqKkAL5Cz3K6rNuszCJ66YxoK7IECGO
9j3OxzNYyUhFQaeG2A9bLT4DZOsizJwuT6wfSviqauEq373CH+TWQgb5CBS4mmsr
MUamozXz6NYyUUZ0Pc0QCGJxRCEM1BbprACShi1k60jYX3Mciot75OlzYkqxg6jt
WJEFwMOcvi16fn/vm6D5SAuOCWN+6d6ZagUzG3bscIfJFUtjlfQ1iAp9gWu38WBR
xEjoxj3mxodWWrEP6QHn1CQLVzS/4LwUfOJDw0rwjUeO/gcXHzkbco6i7QTdo3BE
LEIGlUCcWEaCJJjs3vYWpCQ6QmHd6hz1yPtSDuDYYLzdlfps9qBXZlWGqQoTPl8R
SotvnkCtjHUfFEGPVofP5+mBwjBjTFq7QCZcfNeMKc3j433YK2mMPBMDzgddHllM
z2YpIuNtYnCMTOSpOyUhERDsbgFHxgtI+SkJORfdcRWv34VvuYHFVXjNgpkofr4y
w5qAZ7+Y24WpEIXCRFeCEIpnlgRLdM1PtdfpLIhdcZZOJc/0u9ekrCVUv++g3eyf
asDwBuXD/vo9VOatZ5rdueyc5KHDxo3mZUwh8mrIw+mEkZ2v8RzVfQQm844QbCBX
7NdAm+VKlx14Wx/3dIl6g2/9FaD5Ma/9fsLALQMQZrEKT5TFgPWmYrS9rdojXnjI
gKC841QeFWGeBE6ZkLaNjx7f5uOFiHE6GQ9vlaJhbI0uVE+fvin8ssevAazKPSmw
EsRe8XI3Cx1/mtrDiXLQS+D2425eD8c+3jcJmCSOJ791MJZT8XQonE+5jwQmVcfV
AEtHnbCRHt8xkPlYK6YHy9baFn04P9ApKDwoFDShi1i28Vgv5uRxLWYhrknUeeQJ
GYahDB4jJP+t0HpaziLDlG6UE4JG8T+BoV7V0wsdWnKYgT+UamGqEqjWwk5eeopx
77jVPW+ss/YEpz34Ma/hPayiurpe7WHlqm29eMXwLNLBaBG/UCTPtsg06G/kkn6R
tTx4myIWDDCFumNhrYMid5gUlm2iA4O6G8egBIzr0UQ49NvMU+Pbz6DegluFeMXq
6wM6EScqSbVRPmiaVRZz0e+OK+Q/F3Bpw4RxgzBWNVSGXyse66pCfD8s+Trz22bj
wHZV3EHZQpj5PbB0Ou5MGG4/He0Xvy0in7O0E2L9Egws9c1bFbe8fSMGARqovU9E
6Fiz0Yr1V8X3hNuwBm5LlmMmMbRP/edAfLn73KjLJIgApX6m1ajUHUts6ye5/puQ
CKf8KGG3xZArfzqeWo+OhZPPS4RxhARonP/hgy1UyfCsEdVmVWiv/iuKB9wGyeg8
Z8zKZEdzDehn7QWd9ljOF8hOA3ZIBIKbKG8+ExsWLe3gRKE5EXtNpo2/kyGMrPeO
hsNqwM/4GIdjGm0txjKvHd0p+DJjQ7V1BkFDwhcK4QfUtMr0dDLQ9BufQGTmmi/v
/5U2BW3BskS2garo53WQOFS/TWtj8bUQxy77d5ru1HeP4luba/hny15tF8U1wfW1
O3RaeJODn0oQZr09yYFzt20mrzduV8qF+cANmCNU2eLOh8xBIzERl3MhusHn9NYw
kOqXTAuVF5I/WY+wF2T/KK8xqepz+4CxFO5iL4BGNo6j1+Voc7lX9SLjWbkYZLUP
k9druoOB7CcY0xsiwy/FbiGObVNqiRDEp/vxTnvhJV6WYSe0q3wSGId36CsGNa2G
LFW9L4qonC1UZSE8pmzPHNglQrY7As4o77NxYQuwHACNVF+dLxTz49bzrMvUmSfM
RID40n5ZcMDoPYv3dGzpqBf6XBp1XZZ0pr1rnm2JCXhqvHZUpGWlllYH43wb9WB8
EzLEI+DcPsi+gQ2mbjgFO71bqrFtaNHZJfaAoJzjlMVsHJzveyrP2wm44DP117fU
Q+os6QiEUA/t/+RREoljdmgIADEtyCslZb8rn2h+/FH6wG7/T6uXnyWs3Kenh09B
91yOYrJukPVZBYb0EOW11iVewhppU2SMWF9nmC6mLQmfu+hXb7pu5zA0m818VYH1
JweAqxj0F6WQBiQ+4M/e1xFZvcWgzqXa/eULNTh0wVBVrzcAk6UxfuFtlc5MsY/e
ntGPni8GoYrNJjMPRACypxda7kqvCP98wRYGCzpPfabSiBFCqG1dIqLahjlq/YRb
Jwb8Ka8aGebxDixKDWahlTp9s0szGfZPP7NYm3CslpG0xttLszgvSg82Vt17VTUJ
dU45Ky78BbI4fFz7cRj4agVNGYAxMd2EvozwsUm0oC7Boj5yrk1pf+tG/y/vhG25
YHMjeT/lE0V7x3uQzftmOGP3EfBi8QnXg8D07SnaDfC6o5c4YuKjoynaLLVl8G1S
rV6LehJnTTeIxa/6rtly9OWAH07wS9Qd4Z96FdqXOLqFS597G1a1a/6lyTK3xF8P
VxpoXxMbPGXDS/15i8hGd7DpIMwPOpGxl9yJnVfdiP/XbnqArDbFapXyqa3SaPgj
7sqNFzeKIcqqfWqcJuKcqty3LlBmDn8ovto7hHrF4SXnb9K0C4msVnALSU/p/xHK
+Y48u6ArVwZcCosrR2oZ8xs0c1T7qAzAxTTEq4DKGKDc19uOuUDvKfQ4DpdQ+QGC
w4bmCOpkQz+j8fm9HMf38TtWbKr5urbHwSMyM1E8bTFiZ+EX5gCi5OOmTfTSyQMC
CDlt7KmPOi1lXklyhwjxWmLv7GstNCHOTeBQBb/nqw9qxtE4DdkkcN/V/i0j3SmQ
klGkKxdoJBGTlksQLq0JLd2LAK+FBe95gJ92kw9Fc/rlk8QYHGK8yTqSfd/2X0fW
U5bWMoQTodqOa6kHnAZquubj/hTTzf19hxjGNrev8exDddXDt3SdkoHiDM67/dvE
CMybxO4927D45yjIh/LnV+Uc1IJ5gcy3EOYHNMiDuOQg8+PlDyFnnHc0oBv/Sis3
5LYn8i//NgniJD0g7ytxSbbE81ZBz8qf3Au9UgQguBKbvJLAvGl7eMflheb4og5e
72bwUXHpqb9oS53LttO+e4r6o6IdAfHfw0ssnDrCOGQim85mR8PF3Z1uHSMo8Lld
U0tAxwchQPH/x3qQrRNY5u84vDfAQOE0D+koiv96ArSEfpGej35SxRGXDA1qZ3jZ
WX0c0eBebjy+yRdg4eqL4pAyO0z9sP/D7naAhATzVZb2Dc7NfaoSBSQvOT+BbPvL
CuiKi7mh4r3c9togBAK9IbtWr/iGAKcfzN0KrORAwqyGqHz3pYSpEbdRiG/E+Cxh
8xnnNggfBSVwibrjpKP+1F2wSNhzR3aF/4puhfktJ0BGtTANatZS+IgWXhKK3Nlp
tWgBM9cNW0lM028c6jcxRlEP0e9Ebja7Ba+5T0Ew05VdPI9nYdzucP+n0LUD67Bv
zd8tJ7J5A4Urn/Tpm69an5saJ9mT0ZnsBp1fG+M6Mtg+b3Gzan8qLn3mgbowzWpZ
DZ3m5oOc5a72ORGgL54IuOmlOKf+TJAsfGNVJILFINCPIZlCp6AtwjhyKvvsXNrr
OggnKKHjnFwWs7KsvxsmWYnQU3u33taDCbR/hqkbaOkTkSi2Wfml4Gr9FfAhUqKs
uDp7XtP3YhV2l/H+GFRRcak1Mo4bmb0Ki3+dqXACEwAoary/juWLypukRyoNfnVM
+EKnZdtKa8sQhiAv464sIbst4ufdthw66gUAqVe3eiaaqcqASo+0/ccXemWzsSDx
kk0o3C4hUS68xiqLCp8yij5cTzCTDy4GHloICNkGwCqYp3m3YY99F2U9dvA+H1ak
afH6Kf3GuwY6Q4q1OTvDwNvgZCGTtr2rfe7aXiZ24w4+8Koggp4hxMm84RrB9Ure
DP1R5miQZkokyYYHBNcg3iVbkNf1c1jppqFUOxc/nx+gAfa7kp9Eq56V5be5ElDE
SvzO6KPsXP8vFR+TpjXOXPS9EUqawWIsFwQop6gIezxiFnB8PP+VwEiRpS4Y59cD
bB69mH2K9kkD8avUh5eK7rmkooBzBROyFODcOaht7HiIub4HryQX1nz+jHxhO3co
SR6Ap5WC2HBa8LSKQAtTBNM9v9Dmv7RMAMaKs5pylKW3/TUUnQBQKJhrb3A9jTCD
qASeCravdjtQWIq4Uo5JE5tslEsxBrauz3NjyrRA+BSsxAHwwA7yw9NctdLXpFi7
geKOrRCuFEZaFE3oC8/sTouD4jHcY3fGBsXQXXx4+HvKjVusICWZLLYl8LIhWFe5
peu/vzwyRJTMNsIjJb6HmnWwMUW2pYcJ718f4ZYmEoU0mRLpH8ZTMpu3036Zzi6z
JiH4FSlNcjsDT9tAmtRG8tkDGrVstL+9izDxM1xI7lYoU8SDjFS/WnHLPz7pacWE
suOFOsRYVpefkQ3xlB4TOqHqBm6Epqx8QKKei9vAwPGMH0Dm5U6AMG/+QLcK36Yu
61Ztcvb2JUBjql3wL0uVZdtEq+dJR0DZIwKDPQaZq56nxHG0tlV8K20JjsLJXCyj
sfCy0gi5Pl2JJdPMtXYew0cKSUJS5zO+p83OkHxoRh5Q2iWRaUTc23VqCndXIkKt
Q6cwsnhFpR7etjgQwZ1vK839LbxK8/T5WMNTdKnlH/zHVGhZ/M6/4b+uCX1/9pjF
77cmXGrlEDate+HaRmgwtuncJNbvTdmisGWy6714U8I3Pxsbz+tnWfL0onZiZorz
rZKtH5XCyuJUd6I5rXp4VuGE62i//usC78w5sv89MI27deV20yf923+wKNAyC+zV
xLNg+CDEhr1boPL/7SbZQGydoSQxeNf5iZmNJ/n035G6FXtO65+Ar+7OTdM3Gt0V
0ea96qgWXjE4zzLBLkLa6U52RQ6lNJ/DHzxLooErx90/4TeGuHeaPBKyqSEqCyrE
mWZrjXk39H2JblAoEW9i6cHns66xbYSnvdqLHgyWZTNFPAh2XN6Hvx4DLpMZuV76
iyoFJ8Vv49rEfB0mxgyTqrI65N8wB42Q2QDq6RP4giDfkminHpNH6W86PXMzHG3J
vM44S7Ila4mrwgYAq86mY+98WyV2ymzH8poi3HW7FLSBHbdfTFFye6mKNcWJ5F23
MUfd3CM5lz8yts2Qbqf2USTuWtDx7/ciBpXIdx5Tw1iiMWw1ovVoIcQw91AARygS
5bRiPHgOZSRDReItNj4JsGnNqKYRYY28NjHccRNnVKK11WSw74jRPvJS5OQqAEon
W/DIFHSzgl9AHHfJJPGOd4/rrZQwLiE99qRBrGoRcWo6YZsSipRSMSRkSx3k5NAk
/uy5fA4i30G4ydJTczeFtJLm5DnmF8C7SY2u8NCmbTnI3sN6BwVUP2DyOkEwWQZf
U/sI3LAkRXjESLTjIpiTaoBr5dS8X09SRvbwTeaituDsLnhEBqRz42+nL1S76ck/
qOPxF0Z0ktTVeN+lXrb46/F94iubE789RVTQ/n/pJMSakz2gAvNDs9W5SWO89JDd
pMCNvt/QVC6TPmerUEZJs2OuO2eY3i0RDZLFymdydfWtBmzo0WVVMx1r6AeY/BGb
lz5E9ycWleJoTmZcVnOBtFNXa+jWUtULF+G7XKEPsC7FqettXFEmoBExJs5TCrCC
zjAU/pQhlV7cp9NoyXg45be/jfwQjLgZYs1qy3QltAi0zaf+555IBaLV7amqToaT
EvcC3H0Iz9wlsDbBSCX8nJ89MRGBYZRy+LY1/j3RPnrX5H7EnxZ0JRNIXUjP/XOT
K1cApn3UFbwIH/xB5hjLyJK6Ri5oBfvvk8RyeqCjSK9vaVPvi5jfAPsfB4s1L6B1
TNGkYntjXu3lpRAtVK8U9+ox5+0e3pqfSE9in71nkLfJ9VQ0l5LwDBlP1rCKeKFV
Qa0IP4YeHT9i0faA67eeWh2L8WORIFyoX7hEU6jyCe6ljy+UwqFTEyvuhuhRgX/f
rEUvfrIUR0I0HZkaIke9YmmdaZDKnyEXmD9cUkFosL+9wWC5GHeMz3nT42N7wW00
tZXxBezlmb20BHOzIowYoBLI1QtPQU4wFZqDghPthcdhmRf3QBkPcqIdG21tbD5z
XzKmcidkTT2UkUqgqJBncetAUkujAco2FwpcntBLxgzaR2rTiUsC201nN7juL5Zp
cUWECdtVtkZ3bdPFiD25f/BL2irdX9P+W/VDaIQt/4mj+6Dl7M7/3aLKbmkuJyrO
KLZtNsx0gWe7UKsuhMO9DJoUBbS4KxzhgKG1cM7Ubick0Pv3BR3UuacmJxXzsHq5
VJtHBllRAIhpZnFcE4dDg1I4kqz2j400+HyN+P62CwOg7KrCBkUw/mvUikZdzDwD
CHMYd4o6zj8gYFGqPsE2L7T88PspJ/reJwKsuA+4kzKaQ469NlsNT4YYaQ8+QCIs
eLkdNu8SYnq/lYAQrgsh5hLKlLMPf+51r5Ys9NPALH3tcxHztSn71W4hqrjrErCt
EKpwOUhr6mRsD0dujTb3+veq9VMKTyOooeGcTiqQVAPxkVKdGN2awreMXPiJFygk
+UZHnzbORAuekEdNQcmS77OutDQfGyCycgx/Q+QbZnEh+UbYs82iWhEihPm6EgX5
5AhVtEpvT9284qpQcfo6RJTNqQS6f2eHhTVnki0WN+ZZVSOZ3uHW/l8gjjLDA4OC
2MREYi4+9XfDX37BNCDNqhpBLiYfE5txVCORKhj0spXF4hrzhg4jrfaTLsQmq16X
m5Ld2aOd2MHyj6V22x/tIQkYY9mYrySNmrENOPoumc/GATsOzFoRHV6tTztWxCgz
rdXhc0VE4VEHTafao55RnXvpugOZOkLxamB3nwBZxyeXoUZUMyjzFXVTwSwWrlZx
pBjTGA4p85BVxYytvsEcHq+MAxG3rgI9FEYLZyQ8YeIm7oOTTQ3+N9gtlTZDr6jg
51qn4cG6Rh5x9tP9OG15665n99q2sBpEeocgKg9ZTrRHs3ympetXRo9e15IDmr3o
kSKrqmy8w4ldpIXPPFAbDzl0LVg5Irq1vX9fONw4CxmsK+7/ngNnruM+R9iL6FXE
kS8eftCVo1BUlFvZsjg90DDaEizsGjmbcy1rrnUWUWJhlQ21wNrNS45YU9M0PMyK
w289FqyN6Lj9tVcCMZcEC7hN5ucF7sQu9pKiGGZD8X378nUaYd2gpqlf+ZMm58bw
O5lBQiuBus4MAdQ8iotx75EB/JPFHWV04QYJu4Lqc5N2oCeBzk6KeYoYVugIA3gD
bmZcSz+OH1du5ebuWUj/wnrA6zzVxYGXCggB3o6p5PYFtR2qzvSW9dg9DqMHRasS
o2lspbOsZJN9fbugB8MS4wV2aNh7kU25A7XCgHT4aR6JqbsofE4aUq0D8BFlC/i4
mgVaw4B0fCofPMGV+FEQtdLXucCQ/qZK9yJRthZN3w1DapNPYMqeu+Xo/dDyZz6G
ZZHOTZ59lGrmNAQMLF+JJTgxTR/cC5rzVKaEFyq1+w0vgEuBx6E+2cUOhpOpwtMl
+zlQEEdLbfmY81lP5VC74/FtNNdjYE8NqmQWzov/dXfHFar7al4pmvOoLY0CHj24
qWFGpGGGdQpCqHE1M7daBmsV3XfK9qSLpUQor1Lw5iEOq+z7lU3roz3YHGdUPt2O
WvtZouUXwjMXOlSChOwWs1o5ekRIu3Ov9b02y2BDz3b/m/o6n/BBYpGlOj6NORF2
Ue1QsvKTQBujNf5f5i8uZV/V0hrye+iAyUJRZv9iZUbQGCelASKYZ0VVMMWHyKma
/vYP+bp3WZaRdyqrqbQefxvT8svAKtz2xFylobSHYzy0+7ZhMfDU+boHrWuEaJcC
iMalYcayKDPnL1CTJjV6CAm/fYN6FB2wWtzdb+ZOro7UbechqEC4xJttpCLfxI1K
E8MNls/hAi4fb0bKA5RE7fbctxGKCWv9ndFaWqmUviyYiIRcF1Y8htKejTeA61Bc
WdnF41gnDaJeDPqozr16v1mUnkwru+k720Qglu88/+f7Fzzv8EWvtocpehF2YZW5
F2EZIBI8NNc3TqkD8/fVlXOidJh00uVyH8Gsox8hUkBnwbBDVpxpnxTfhLJnpNAC
47iBn0lG3FmLBqHHfGDRxo2VJ8ezo5w9gRx1zyUieB/cME+WDr3MjaDEe2VbBwSd
DO85DBum81JpSSTy7XQK3s2NE9hTv93jq4a80qF/UFyrvd6o/MZQUvNUeUZaQ4So
Mz0N8Rs2b9DsrPz1hseFYmMpSlAQOebC9W3FMwC91bGdkVDuHY4jl3UBetYdQHJS
hDkJ5tWmiYbo4vo/wH0jkh/YRQ9P67eOGLVCX6rjTt6VjMuqc/lpmnAfBIzyhoEA
hFJDLlRrvfOOZkJLjYR44Uupt2A2Dg2JAkfoVw5sA9ioqu0IVxy68DLU/wJI5Na9
l7YInXvCeNb9s6reWoUMPCQUGH6a5dn37L0EgIPw+lidwWqxUDekoMVtk8zbK/vT
ngE+3848b0OqTCP49g5XEWesetE4p2SkT9ODUWMPZbgpu25WnzQR5oqCtMfiDxJh
3sE7IaoHctbNG52f6gyEj6XFaAfjOE61ui5GZeBXhZowYYzhgBe5J0bvIdppxYR5
YUhvWFQoFhbtqmJK1pinSzwyECUy8jXke40MqGef79tfhA+9I5kcR6mnZ88LcTjX
Q76NpRvOlkDL0ISreZBoUjtPSuu2G3ShElo9yF917bL2OR36/eOKC8s1OPSLrfQT
HPDps4ifDH31f4MI0bcRzuwDHmzeRyzFJcAxK/2piftvy89UMTuG9S1h8DzmEuvL
lVFXEluNZgvmdJAGZ6nRLWIdrEmfzE7MbnKMz+inEmgkL7qESwTv7if8jM2PChSl
oLG7Ps9NPODW7vRlR067OG5lM4IOonicNIHo/3jza6F2Z5weq73S9O0a215bofdX
+UMTmFLHAYayQRS/CFk4y+qiufdTqKKvtDJAv2WElIeJCMyN8+WHExb4fCmY10h7
4s2dFtfbCUhQuwWO1zL24gqoq0xiWaz5kR7fM1ZYeF/DVTJY4EaZy2tFbujfaErC
RDNMKKiCgKcGSdxTOYaBLPglYU1CKoGzK94U0QmVKpn7H3yD8LuDYVnANgstJjNk
L7jfSvhORK9PaX07aMY82ooaXsvnMDPcHjz8rcqBUJ817413UR2rybipn0xVdWHf
n7JTTSc9I/JKPb+oa0gzBEyQc3DQ3MmV0UBjjPkq2/HoiXPHizqwKJWlk8kjKpoC
0f291fTbid8Uv6tw7g18QO0YS2iT7rRgWk9vQLAzzsV6AUwHMqDRa435jEbbOlPw
HO4h/d8R5KxAeHsGljeDDO76uYtPybQE/T6V/tuo8xb/a9bNv00hmzN07nUHCOoU
OS9zfxr2wDsfNp7wnDvpsuzYjAF1y2QrG8Unxrng7PoAdt/imK0kPYxcG0O8wr13
6LXcSn2Mn4VfrjhYi33QTX+7Wc1/lmUOCigslno3Is8no7VT6O0P4loqx77yFcJi
Zbg01LUIZ6xUrGPWjKB6Bs6jpr792NvF79s7tDFcMd4KyYJ3/Fc9Ia1k5PUcoLo/
ja0IJOICZQ6mt2ciBdwysHWLWx/BZPZj+rT6MZTyOxrdvtTtQHpfLdsVkuAAvRYE
ziXhnGFdzGCxGHaRFCZ4+4fTGKPYc9OUDsM7cSOpOMppHucYcfFaSkQNcldX09ue
hy1e8ww5ACHQbz40XDkaoSdWvltnkOVp4T1umdA+UwEBHq5kxhc/DEs0e7dgGT2M
tCNTQQ/C/fL7E97heGNtdAzBU9TlQZFXx85GjQGl3msu7m2WEl39DbOWr6pyK9/u
lKePvUcxlcwlyjUs8uIDzTeSEhYbAYEyM8MM8a7g9mz1jD2MfT/I5+5epzSciBgv
Y2M/cnjVFUvCM3BmZnqvOFLLTFmRo84jvAfncQtIE/w3WuCeKi3zAKK+JnZVJy4f
n0XnbVJt8rY2CyM1MxKBHVzEoaIM0OB397wCcp6Gt7QML2SSOY42KG4QESh6YRuR
LFJmOswLoj53TOb5lHOAbeIB2ZJ4Ia835EKVoUoh5dWp7kj4OXqQ3tQfPUkHQfDH
vpMbN/apRsLyJF3zA1PmdG3IHbmjzgBl5DUxEzHh/Z4K9/AaUwMdU0IMaks/u6Du
MC7k6d7SBMsXiqCWIMUkxlD+2qMsMuDG/HtD08/paeLuy1kcjVlrqTdsm4TelCW+
738WDefpq+JpeNPbUm3EMIrH2q/Z1jyTyGfH61umZBH02vT4If3ZU6abYDurN7cw
n/ExoHc/psPzR6H/yaPvsGn9DLwGvmyHITLoGZ3kpKm2znkqR9ToLYyV9Q0HPekr
Doi7bEjBcFPVdqr48UMi46aJ274f8qn7w7KkahrNH8wsGPh/rmYpiDS4WOMGJkQZ
9WXahAiDjt0vC7W1bURf1EIsllzxd6Us+jkXU+lJ/M/TECAZVfUdnzOHQSotEOS3
IpEABkDRtdF6QnnlM4arDOxUoZlY2YOLXXAJtNXQf08nNGkkT9yd7pYUIsr3k1Qc
41WQTTJ1BqKqi1SdI9Z5P/K02GAb/plFsCHoEVXvmdAzyNvCVFczhkRs8upC+YrM
qk9/BlcKKb5avsLMebo07KLathqesz9DOwxRgODyHc6n5p/pwr9jteHHmUteupKx
Yn3zxuNci0+QdC7uKl1g8jur5zyObBBtkQm5P4G61mhMb8Ttgyhm2IMyD01WYJL3
78JUfaG3F3t1d7/E7m/lG1/QZB9lnboRLWubCH7ZMUph9oSl02rpT5wigurb9du8
laZ2+97qakwEv5zU1SIsYZCJ8KDVFv9fBRE2ebvvaOQSukFQfgyRHxsZQG2L8dtx
yyUl2H4Ju4ve3NJCt98zWAmQNRfNa2zDTdDh+DJifkp7bICNYd4powYb4/MV3P81
PqNEKOYGeBiH7F3Fi9b0n68lT1OstEdUuq2uMBex/shT6eGAmesGsK/vGKtuQS94
X/7p6thy6esG8ImHrvRViCCjBdpSzf5RvACKIEIYJYmOTGBGU2nsTXPibh2XFubI
f1ktYo/2wS0dTluBpgPnthCLuhFi5N/oPmUXEOxCTUhg/KO6RX1L53qdAXyYubG3
7N+0S+z3IGO+HeKJQlAQF9ywN5yS/eklec0MaMZWCOuDbBiAUWqnSuMGmvsNSoDi
ygKio9dxwyo3dezTzDnXQdU58Vhei0lHscExrKPLyj/P9SOlhmXmR7n5sficUwjt
exdbKoMRG4zUQTnfKYqPiurYACv2NLBWZdEUSPFNwNQQ0YiLUoyTLbmI546IF/AX
j0rYjyrtkp8YloRtdR5Z3JnySqWSD1MbyWhoNU1ifgAPnl0La65a0BaBbZze8MHO
Qb3ndJd9Gm978fcyBe1v6OsnLIqKaRkQ/LEegh+L/pVLPvJP53FN+FDbcvDXxkml
V39BLcayx/FGq0Tw8/UGXOc+pW6+v5ajqv+gELuiuHwgwcve/pTrLttdZTqdrHqH
9ij2QRbN8UiLSfdr7dRIhnis6COaQMy1ygL0rmYFfdCRtTC8Y1iHS9qI/l5iChKI
X0TEmkZr7jWtV4z1E6YLo6tl/1MGb2OmnWUeV62+Vly9xGCP6WDmuS5jOiZfviZP
RSUS5E0IcR+OtvEaPed2SP9QGGu+e18tM7PUXsk8dorjv13wVHXepzDilt9ZokcO
imzG9AR5ErsmersVf2Q57c0O7/Yr8woXcf7EUvWJ52pY1uHnGUxf56NA9OvdV++P
EqJ0G/YbKy3F8BWIegGIJPNTz9LCnyXMdUuagLB5faKvmTheTWWE2yVnCum0x0fM
b0T23My9qvlKeXFWxQu4TF7KXMLqQQ5jyjUcn5XgvoG0dzM0rcPicDgaoMG+LR6Y
JcTBZO0lA/qmEdmW18dz1C++9k5C4y4LrelVSU3f+Yw85KoW0Sh08EFIgsz7E/Mz
fZfOrfUEwgBQ1FiE+AD97V7vg9CYeTmQFQ3KV2eC/nOKeqQ25DWcYTe/fhmK9WZ+
ipHxV2X6vnW9dax77SnpE8fnAcQA66MSF5hdWJnt0b0ZK/gykb0vPz4dgLxVbId6
8Z8pz3zDCMwzjUgJ7T7RnK/68vrXplF9vLunGXzNiGQ+AgMDUCRbgiMH+gP3WiEI
8DssbwvVbDy4/mP52cP+7u1+jt6TlEZJS+fPXE11yUn8g1do3YyRqEAxQCNWnZla
3cmMLXZXPZCM+sl069nkuxMl3he/D20CyaxIhNlVkBgmImU5vTfEDSRSO8XFJnO6
GNBGcSB/AAvNiK9NnwXnNuTnH8v6j7PFttqr2b0aQ8KNaht+IzsEJvlPG2d+HVdF
5wSQEr1nZvvCKerY25eWobnwpkyJ+mEcQSfZ3DKiAr55vHyw3DH4z4aohbKRWdaF
1TVo9BFvPOIYMXaxpDHLK9u98Rra2522Bs35oY4dq3+PNxmkeBSr4plHjYyzdzK6
1yXrG7Ykdm/ttTyibMJmZ0uew1L/uPA7e9mqPil7EV8C+5uZi+ibxq/VIjXKMBFX
B/h9v8y+o+uwyMIpvziT9UlD28iIjq9xC/CHCQM0Zlq61yFGznr3WGnr7uPzje5V
7AHr119AM5XXxeXn6FNYBp33v/7hVTMDioYfdHwUDvVNlSyrOV6qk3aaS0/+99cw
eQYpxHIk/vyHMpdhX85YR8rXtcS1bsKN7x6WZEXLWWwa1wpH6quOeXszsNOo3JFB
mZ2bIX9viPBY0DA0AZMXbHGTBCv5XRqfncN8M/kCfRdumQ9k2swzyNxTB6xqtNc/
aFlxPATUpY9ngdYqa+EK8buuvmtKh8Ui/QggNwyMVJkMOfFdMl8FpHGFUXYmQwEf
ir85/4bkFALIPOTymkfUfxkWk8YNcsO8wz2xetlQJyTHE4MxXpYTu+I63KVZMp+A
dzSLVAPPtqz/eS+Ypn/mi5GdL1UmRtaUqcq/r9PlI2g7v2TeHCBPwMqppf2DmBWW
bzXQyHSLHy1uQfc/oX3JD7ApS8hjlaOIKodGiB/q8/U9L0fUZrFIYzLEtUWLEb6o
hkEGRXONzUeNcw6NEPrU1YaK4vO7Ts9Gk9akE6JT0+C9VilVuJ57BvvUkrsstTS/
ZuUWgbnpj1cutUL2bd8p0KYkS9f7dpEnBpduTsboxDmtkPhw1xMP5qCFb7icn+Mt
NfHJsL3eZQqOdvOnJoOhFicvKzTH5HeAFhTxRyrvcZsJb6kVAALOlC7rhB5lfuXv
qWr5w7Dn5hbGPA5Dws30/SDzXi2MZqmYklrID3aFQpytn1NqtCthyRBgQUMC7vsH
5LwXriyvMmNprh3XuzZqp63TPM/kqjuKuRgj2JQ7bLcPbEJ7i12Ec5+6fIUDnzQo
ZhQtmFjFFPp9gHlais8MptTHs4p3cAmF7dUvcwUt5cqnM5rGW3+F2ykPpTYKsVZ7
yg8fsDLUkAe95/zAm/EZ3QrtkbB09Q5Ho6ETx6hBQlhAXrnhgVMujCrxaX+7nLwh
uAkz2wI1umlGZR6CkIS99cqS5zvqftXcRHmnL0qcYTTLhogCfmcuAd1dIYygu3Gx
Da5Ze5BKsT0B/aKPTw1KCuxtCkUikEaNa088MEJNB5/+JrXsUHylgCz2e8SDs2um
VS/VLyJ8mHEwq3gSEE4hhz/QIcwEIP7uCMlNvdZaIoydMaxuU+hRMisTAa38GC88
pOU15fHLDKwbH4fGylLzEyElMkDhlnZ3YyORGJo6GSAvV/7r7Y+exDHWmMH2iQI6
g9mn4LksTZN6pRDlo3CJ5Gdq4K8+5dCClVPMTJsw6naPqnmtKSar45ZyjISI6XfK
RMDB/eAZQRlGVUMxe5nEFMUtfluZuGs+lGoPE/NuYcmraLn5Zxoi9SP4Ggo6r4lY
6uNwDdhwO+dDrvKA0Hc7bqvYMy+zVC23tNFv7C/+c7RMXJofrYw52yLwioFyDXp9
ypBjlzcOcjkpgTxyooJPxWR8iSU06XnbPhtTNJw0GnQOrmq85tAmJfoOdXCTu0Ff
xWornz2AAAm24AFuPR2FcrCwYRxNiIi4Zn2CZVxNvS+UdnOwX9TeamaISvmodrAh
JobyNCD/1o9TYDLklvEV9PFZ0WLCdzZI+pz1WY35MMHJ58vPmMVDW1MS07TpbIrc
TIxfQaDKLpaFH6DuklmrgQt808vmsxozyzmM8ngL04B+PIcVWRjgMGHwxlZcAVrP
HyCKnT+LW8BxPs8IZddFt8eKuVrHXtBWs9zML1zJCLvDhyc2oO3hg+Wq3FtLQSn+
3naMhbuvxVqwnNfC8HujzD8Q6KfkZ8WYMpDDRGb4/1DIsqgsAggFVv0u1DUdjmFd
53DNE0U3ssDWh1NXttfRiKPOZUO7c5/wDJ7HcV+oD8VFA6mDSXo62qzhf0qVjiK3
z5Iy17pD712GJrvukc/UVAXggcSVBmp1UiQRo3mejEQMWtqR0kEyctb25kz1nWB2
uIdEJLEbJ0k8/7AekbEjDK/1Ohm/nJKR1nOqgu6+bY701nGlyJ0Pp+4V9a7MXXKg
yyahOKnFV1hOvJrx9YVCIS+6Ww48GSm4TziEgCTNsUwUkmSDTicPw+e9JFcm9haS
ji7V5MUbAEYMeB2WRh8c8UPJJ3ceFt81g2X0n5HqPrMshf2bHoRbWvNGWwKMsTEw
vShLca33+jPLiJz2QRdjn8lZ2D+0tWqsOBXKPizenQLsSSAs1lqa5pxt9WBot5SS
yjxfi3ovvAfBSq+yGNcGteuXP/rxjZbF8bfzCSw7OqrBJuNSTrUQECiz+ghxhJ30
e3hZcIGavD6Qr13ImVSOoAWiNVfvelE/wwervCpSL+rmhieq/pG5ZZyleE9MneSR
5IM2JEDHuwvVat+scXK8iEf33ARu5tioXzrVdWNSUSYtlOgT6qEA2XkuqLf6qHPu
EON7swu6EVXUNwGiQqaYigMnSo5TW5SBt0MvVV8nm1J0UWNM7s3/swYtntQ1jpZW
Zhuvebijtb9hR83SWeEQp6mZCndUTxTL/cIlB1fRcDCUcoGp+g6h9feFjzintw2x
b9qggP/gyIgjK5UcY6ij+mgaqjJ7CSqhbrxW3QDABZ+3siLOniJQy6ga4JsKtHtr
JRJQbB5ou4B8iyHpj/VJLOGpGhLUm/PriKuu19ppbgqjmPrptDTQ0N4+XC4bOpOo
+5GQgSVMyaGOSebHc4KD/v9U/qKJ+AkjpcigoW/5d9b1+XxzWl55IR/OXitVvk7w
TZlq4TWMzATA018zr8yKZZosMboDdO7Mq2DyeRYOg+MvXLmB24i/g0iqMWyWzlne
E8jKiA+e4ImiqaybsmiH06hYl7oNOTb1EkdtQDz3mJVNm3n09DcSPTUrbJcL9YoT
x6yrD/M1r4SFejE5AH+a7JJTVn2SZqKsAVgdUb48A5X2+LH/SSMn7vRMDHprMRLH
Y8OsZfocOM/VGS/sHsvkuFm3SYP+Dv27OHYI/CwPLXrH/rrE0Xbu7RJwaRlFCJos
vxCUyuxvPeaG/PE4t5y22FcaXIUDCf/q6Y4nvKZsVo0tGDHY1yH/o2E+1OSu4QFn
pCqKjyOU0OwVYjyh5wH2a7De1Zs4EEc+Dy6YsWEtMjdUSHI9DznBfAwAhdp5BwJD
Mf37o+gaT1XTztve7QKGCxu8Wp7+RfN05HCO0vWLQIwpwTQJZXoJ0Tlt5SZJYdqw
yLR7J9nXoua1kqNzMnSF5t2OY/y3CnfijlzfIbpluo6DJ7NQcNswgF4/bmabN7u1
q+JacISC5UeF6/9RIJsa/ATImSzSkC1rXrEVRC+AVKYruWSZRiq5o6HW/wElW+gN
8nFojh4A6WI4z+SEgBf4ixApp352xnsd+pBf/QVIbwExXzqCQjsBFolao0IKqnLf
QLYtE+BdCTekSimsfmEsf4gTgHTXB2ynO74REBeW0ifwQ1hLgmbAjnuPeDqagejL
Uv6msd481anrLgcEKwTy2jXcPXDCdRzyVQG/2HJK3FIpUKKuw+rQn+bMg5LTtd9K
gFmWkoG7iXdJrTe9GjrXXwz5sKsfsHWowSR2RuIPoICduhIch8xZQkS6iAPqRMEh
iDSx92G408G8BcWPMUnLiMoEou9BGlWyviTIedelr+vfn3/7v76XpsEzNrXOi1Hu
KLazZNqllDR8ZaJS/9/cK77T7yD/c2iZKEfr6GdDrzI6QI2K6IgVjrJdRzS5gqjj
J0W/I8UGASCv1KrWLvzAKNckRcBkuJTvE2m2eNfZNYy5qSxdIPQCO5uSVrkjJWPC
2ecx7sBEMJNDSz/iTZP/jb++gV/xVZvkB2XPJZOjKEiJe4NRpI5g7HSawjFPpL4C
0+JridE64zj5V74kbwiQs4+uDWmylXc0DFSK017zaOOtAxp/9MVbLbidXs19ynwK
VGQ/q+0ZhUBQeeppVNn8jQlk+laRTLwNhaBh17fbivcIoXa5VRSUjzySA/pyu4nF
FsmvvjfWPbs43I0yyK26/QPpPKLO7kMlEap9CkrWlUuzWiyHMUhepQGK/TgT2Uag
js0hnNQhXp8HH644CCnip/XlLC55L/r872uVT3l7dGr8gdBJFuYB07L5X+95jGtY
1UrW52MRjt0wWkp3MGxctlAIx2jiwOAPFIyvlL6VasH02WKhRYcCJBBEEZI2speR
t6E/seoIxdnrOqypSvwGDI9+cTEYioRAkQRC1ZI7XP3vVcxeFlIJYWfVHAWTJVPS
UY7L/LKJMuTsX8+pFzCYT9R2AQNxY9ZzGI4v0Ct5ybyNCuvZ2y4+SiWFQ9JG9B+X
Yr4in8HAHgn/3d2AC31SFW573avEXf5Xz3GjF3exTBWHWeJIcycTJhsp0LnjKyY9
Y8JfslO9MEDE6meeRRTGVxWnzOP3OwzH7y2yWhCqiF1pPlUclMpevWAA+SPgYaq8
B8WOYNT42EGrsMsfJwIVv+B4q4acT3ZPjFr6bQQoFErAEmEGdV910t/i4y8ByiT8
ODaraWFToyFNia5iyt/IsGfFVDme0f4anMcn/CTbUKODbUdsrp+wyEowO3xE8Aup
UpGsroePBOn3HdgntzTkE+T0v8vnAocpQWH+51D8e2odd+HBUdbCavtt5P4CrOne
xSWpj6kUSwbQtWUojiI5BrHQ4CG8cjaPjlzARXmqtP1JKargHC8s6xe4bIS5Ysv0
X1CCt7fnJOzweGRVaJIUu6FGZQxIFgQCUNs4B9kwQEE3l6WyM2T4yWdYWXJJ+nms
kFi+gs9ur9Ncgta9cpvm3e9qMkohXtRL5ceWLuUyGt9bx7JG9AiFsN3BNq7KMygB
KHPad9ilmiJC3YsO46EMwR1rztHMwkC+2z9sWNy5ku3pgsEBf9K3YEFdVUjTYGkQ
io+X5MQfBfYVXN23fK0w60OuvSUQkZg1I5M5XLnSW6hwHIGEq/ldUFFJaB/X4Gwb
LwQ2AOgXT3mJe+0joR0gqMGetRi9m2hURAfZiK6UemPcFwYo4sDLYbR0sC4eiHHz
0RPMuvjw1fKTypjpoF5lHcZftzxudzQuZOXLg6eKeFtaDcvSfVael4QfQ3fg6Bz+
D4LYW207xK6tZ20PoFTVNnmxIuUvJkyBlCBz6cwRNrOu9zlZhbQ3OnUlH8AW644z
aY+IqoAm3xbhSaumdxmllAnL9TIvdyiA6tWBDnvOkCfCvrAoKbummZMwvF1dQzUp
9DuYaWdPVTs3BagQreHACTCzc73ybqDSeu4R4jUd09SPAIMBjCDK2+NEdaxG4SUB
Qmkr7fqTYiFGzGGubK7PruXQDtHxxtzmNyC9EwWk/quUekvOBfVPywS3i+Vcg/WX
/Fn8svZcGZLbX5uzMEQuAQlzw7m1+agI4GOk0Eo2OmEBGxOPMFsoJjjykGzTozPJ
fMXsOCthQYtMqZ2lid05Xt/mAf4K9ZUUpCGEDzD8iR2e4cFSxB3wzlkiEwb86z2F
icsa7BhPNFPC2OtiY8fjU44noUN7EHcME6iD4Nh0On+of6dgm9ufPS9ZfWwIPlL1
mzSSWbmYLNZ6ckmf3HsjvEfmL0+pFj2XTaGwfekBiQRQKekLo+6D5O62F2964wba
ShJ1glldllmPimKnVDd5YgP54wki1ISQL0GU3xLofG96penifkx/6uEY9QdjyCux
L7gwExWa7h32zKcEjDwzL+WDRKbcnEXc5TasSJXBUMstTjxx1SLkp42IndNDAOQ3
o1nZXHrJ1ftBJnKIIDCbuuD0ik2lw73+77bvTOjui2T5x0/GcXiSBN1DBY3U+Cgv
MOIDk96k8wJOgXvcqsr3UwosbS8W/9a+Sw5MpLYEVSlEedlU01lLtw1I1Tzqhp3M
cgpIApkXz812RzkcWyjK+C36g6kJSU2OAnTXRyL7rpIiw9WoesQa0HS98dV00y7q
noL60WtVR7cWmLHsKnfaH6Q6UjYxtwpwtDvmyw/6aT+H9SUh+x+JR0qafLgX6kpO
jIKv/cbtdhnzdzxhycrT9ZUa9sOMTS7xA5chbYIB+mAZhr1xGfvnaq0KWFEO3kqz
RY6lt8Gpla6Lsgeoj31S8bGZGMuQfL9I9UWz6C1I1ZpoKsq0KxZGumWh9Jq17o3m
OzWiNPs7NLfog9cZXrEurnpYDs72GRmmhAWsWlUTSX0ibSn5B5qqh24PwTc/7dKD
/q2fYHzi8KKi2WE9HdfIZPfpSEW0YExZDSSIa1HJpB5lu9L0caFDiafyl+NX3t8i
XEUhstGQgMlbh+73VvVvuSTwyOQhCKLxNNjGg8Pt5joFWQgYH0ckZVux5ch+5EuZ
fz7ojYYodkeSOehzAMyxEfvPMC2bO9f/9GdR40D+D9eT7RjiEuo69QLywRlHMcCq
OEW5o7HQHIQqHxzQRWnVkzLjNDGjsUZEj/M4sK722zcPpze0H1HNrp5ksKNUB5W0
f+wLH16rCG3Pk5FF54hPTzFgkXvSu4KYrMdUOY06XH1/KEPI10Zlf5gQ5jLxu16C
cZzeYaPv4fKx97PHKHwKsqRAK/TDIzDbUZb4UY7SAoOB5oDLou92QBH+PH7hcxNY
6bOO7R/12D1CoTm8QU/3Id63JP6+8q1gXB4eCcsT8H8ydTlpyZVG1IV/0Qqejh3W
lK4B1qtWPcA/EzQQ992oW5DvoLOO4UMXck58pCYMMlgh7txoH7srEHaqB2mHKpFt
KAvbUMln70rEK4TdE++9rXC2hfJ/2NgNuMG9oQf+pCDPiO48JbGNiH0YJc55B/KI
9NzemXBwegQhiOVTeLWwAOfuJfQTwpKmjH2il7T8FLHswL3CyWDk6vv7uF8oiUxZ
ijGR+gH5SAN2iT8qOmH0ULuprmSUE9q6MzrjWPfZ2zzpGLoPdhLL4pzIwBJZlLiS
LXWaRP7jjOQAae5RNnZ56GuUcm12Vpjn/lYNoWzx7eDd1Or62miTaBHvUShCf1dL
ES30buO+wI0idrq4F69acz/1ZMNHgTV1iC2k9k7YOL/3WhMukrYhZveTVRBdnHVR
30ySmeN2CSynCw30lEnBZ43Zpv4oeIMqGmTM54VwAQALN696YWrneL5tx6q4q1uI
Jt5jqabd/tjVL4tKnG5h06D9QbSn685jajFErcRNOD1tG1+XOcPSFKeIKl3fFmTG
4rYGsk4+FaLWsMSTFB8n6naz3/It4j1XQtbGPqdQO1rdVSQEWBz6gZqeMNpqSOSA
QLmXfqJ4UKN4P3u9Gs2O3iNShDNV2UJ1OEpHC41sp6sCKjH0P8T4A6LNmEXD1A6S
S8L30/v7uKll0YH5yU6Un5go3wpumoYwAibYpWS2wKDTeopJHTqX66xnNyVmkIrO
w2Sw0651ocdc50v2tdwLiWk/Dt1S2607Vs+4WiP5vArI3THVwrTDFsGaGUZ937Lm
ZuwNMLliHMga3q5Bx2LhWJe3mOhrg1pzHZ8/utKqKReZfrbDX+8LY6hIrtCv0lff
nWyH0KS7WSiNLAwqZmpnBFxNnFX6CvIotlyQteJPt60td1odofEdT9Xl9LVyFA0G
+MHCrX0DD+dPLrdxFL+zvwNQ0sMxpcgC/LQGuEetcHgAuf9ytloUvdOkGWGQXzX6
JtmnMYZNP+7CIyCe40S5l1ywkdUWnlnmN7wXWqX0Hn1H12Pnc8/Gxatbab/A0Z40
jfAdE069hj1yV8zbGcSv4fffD65dQz4RCSQjBq4x+zxJKcd/afQVnLdcHpztYSni
aLE9cgketTWPTNaUIfOsjnbl5jijfuDoPxtguyELMyA/JJ5rThJyHp88ue0dkL9l
D9Ns1368Np6vTRusT00FCWsbRRs1/Oa8w2YpKXx7gdcK9Bhb9hODltALfMVNQMEI
SlnYdoR6ch3zYfV8sd9+mBDG7CopXqW+CZRA1X4t2oNnLGICIAqrNj7I4hqFueok
7eU/cDaO2c5kN/H/bGiSWWO8jgNDoYlBJ3qpPjZSqanbtPfC20p8og2JW7o9ytno
srD8S3G8eaAD7ckBROOMlCMcoDHoVpcjYg7QLWfZnrlh0TSu8Axn8L6ZUMWvvYPW
/5RZdqUe4JNLTL9AFCab/YMXQvrwf1D/2FEjNGETu7snNbqskix7iSMtKTFTLYHQ
GnruDZUyhdMBFqNjTM+FZ6uXd5SbNZr1UIYWsD71WepTl2bhvknWQWIBLa1fL4cG
B301ffHYQ5n7PBpgxBsqJe9IQb5baR1q+mkuMK92auCJycVZzIJcqKMp9gIAWQQu
QAlFDtkvBz844llEYRlkVpFogKT6TJ6ZWtXv7Zu5RelY+35+l+XIEQnQHRgxOmAP
dQu/usB1XtNUSOdw6cGNE7ZeELpeL6+AKEhjoa7jS4Z7yoIiniuuzYnkuhVUTDjv
gis6Pv9ahpJ0L21t/pO/00oI15+zkHk6qd2KU1G+RpZ0XEcXnMJSPdYYJVxwzpnl
p2doaMMl/RJsoWzrxswsnM/WH+3kuKoGVxcH5gBPJBOfMmybCZ53F30Yxgk1Ey+E
VRRXKy9m7GQNUPNUqS909twUWDVPWNgy8L5RKJfPqrUdME8usSfslAFHyqQcGMOs
2Z5aTh2q3APDC0LN0qDybEOoDk2t14gFxPxCMwRidE3YcNmEVs3DYOhVunZ2SUeZ
g0dOmGoUXNJfuButWtUtOoricJ6rrxmpOWq/Nme9AuuGuXmIIzkH1xQatHRzduI2
RIIFWfHQ7Qwg0p/M3aDhh5/9BsO2cNd7/1zttNw/P8mTKlpyNE9vx43V7p2Ncqff
S2/mttQScCngR/3n0hMsmhj+fiGY2FR2C+6qxOUAcwNyKZAS7LHzbH+XUAtgtejh
BUxRR6bbjsV4if9ioDstNT6NWs21kd8YopoaPzManVeaQcW6zwR7N3NHW7bNsNLh
n0vcqZ2gJcCG3tMvN98KnUVvc9kRSHq2w2I7VlVUaKkX2YygMsuNY7lylS7F+Yn6
1gLpLHhhdy5IH2z4+HsFePvPrGzlICAIOiDHelOPC1k01aA4wrAuZL1EmrFKkrtj
dG+/hNDI5z9JrnNYgbyn2jfzb6iCPrPIcxMYed0BzMJtf1ayc/7yi6PZ4pDiBw4Y
fZ03cRuRpR8GYDKpSGnEZnKHPfmYpOPjafc0xk/H9jEIgDfOyi0NyR6PsthRmjNa
OlDFjOjJkOOzO2BpybWQB3OiiWAE58JNJV3m2agQHrZqgyFlkBLEKXlR1mjpspzC
INS309MCPc7qxeP1xZDaKll95SNmppykN3zXmU2oOdzUtnyOOsrDqkaWKys+whBG
0XdAtI/doTFqd5NbilFHMojL7sPhxK2bUaMxGVz2VKAaYgNza+i2aBTlUoOzuHmq
M11bQ0pOPj5FMfb9TZb5VI9KQ1+M2tQtraJfT64SXIfgiqQRWVEjcLRQJAGBT2Zh
fyL5xBY61HW6oGx0OL5+im8kchosz1+pIer4Dad0milnocaEMEaLzVRRVmdXGfKf
bocZVNoINIHkc2AqdxPq2Tc0yxQEAqM+RUexG2zkpjYPhtJAzcPfneWv7toVGG/9
e/TU9xBWqlv5APnnu1kYKUOglr3yMV9XZJvkhxTyzVrYJQ8VMKQ68JX/P+/274WM
yWGTm0+l0mOqBvLsm1hGSnA9tuwvtaGinXXjRSpQQt53L6vmVfojwc0BB7cTwqgT
XhlXoL4JKhfa0jIBLk4ewnNz6WftlXHXrzpqA8QRZxdF6vn5FGZinNPv8AaUbT+o
Pof2rVsubUlVcpERVSwGH5w2x3DfJx15c7b6alKiUgg01+OP/B5coMfsxMib/YSf
zH0PcqjXZLz0eQ7nX3Uk8c37Siydv/AERlZw8tqQu9k/zK2aVPQ+Bj8kpjS2kHgQ
J389jWnNtjFHvLDhd3/R07RkIKJcFIJflHYvmP2lxBNJMMXP4lyk9fcUNnTbcBUa
Ke5fLBswBB9lHtt507daI3kwugRdHm0+MYEHiuOwfF68ICqEtMmxNmsrTdjnrsbU
kgK1nlKbGdyEYgA/6JSYjdDPC2l4G17ZduNdy2bEV021VscC9JOVVX5YoFGb1UyS
HOEf0moj6tjUMOXn/9Iwkxbx/0mMs5GyX9idySstiwHJTbPS4lDiMXS5xn39xKZb
RVVc+YBCuJyQtJ3zhxXE352DtYqzEqBG6YmV5WtBNGgC4ypxgXERvJSMgMz4DN/O
hebru1lzl2pKmBiGcGVcbR/vR4bOS9YUA5AjGhjIozXeE2/sU5UAH0qnzarZPvJv
Iy51VD6UOw05Ts9c8g+QPdMXB+LFbf96xbwdWua+ZTdiLi+xNomZFI1G00oQlLrO
oB1kOW9NUajPD87/TiR/036yWf8AGRT0EE8XfOs9dWzmA33f6cjtDGKaK3CfWIry
EvjVatCmqUuUIsspiPfMfm12xcyXgBzm92Dwej5uBzxCJd6IuJHGeJXQWZ3hGAL6
1rPfj4K1ru2T2ao9wTQuAIF3KICZBPS8asxTiNVBAwZuk01iEtrW8JnKv5BlJe/z
oZaR6rUYfYl6RG2UOU2Eptw9lQZL/GTtrDQaNgx6gaqfqoT95zIghVKhGf0O/uJY
SvS1E5VJL16wH+IqGdr4PSosjyt2ADlXM7dfATlGGwIMsHfxn3zTtvYCjj8TiLwi
fpEBuNssc01hj+N43KlrWknEeDca+81Yplr3I6v+MQCjwHjxdx1ljzZrsvsZZ0oA
gl9rJoUv36hrH20Itfk6Gn3p9MJoRuR5n9wP+4RSck6RP9kYHl1oqUil+O/NAmvc
9t9GjwH9752SG1pOf7ihsq72jpLNxVeNnY74TQqQ/O88IHuO3Ang9eLLzWvcXx/0
Ml6MF0XriT3QQ83tOTRgskER0Y7DCh7O20l0IsftJ66wS1l/Uy4JpO+N1yv8uTjq
xiME7VKLAFgY+OW3gkTqeDDqn76kVbTrfeYiy5U+wc64gf9IN4oA3TKFVYg5ryIf
Y66LVdYZXUh1GhPUxvxuT2L2/1nw8PK9HGD+nX9Lo7OOO6ywZEAFDUmxFLu2+LzE
j+2PXOyplD73OUO6sDzTaUD3We9Xz304WaMqsT0nJWpt+aROo9f/2Bo84Q9ugsNv
20bpKqCX1eJHrUhbO8Fopr82GAm38m6PtsVUAfR5gW6LMVJBbgLNvaISM3Kh4uYR
/zA0S0HjsZk8DJHvkPWvJjDvX6NZcYF50MyRRfrEwU8yQNVr3uiCmV7g2oicbZ7K
Ppe4mrMw2VqCzU4ZKMvRLtxu36jIktB5qbWw7H0rrMr0rNbhbvfYvqXhmOSiwHak
/no9Y70Kbm1AMuoP/1SqWK9pzj93Rvogumf67K4vd9Cz207LFmoH2Y01wmPJIOUn
N2lMCnV6QII2V+tO0PYoL+6O5zuC3Gnt9RSCvwBvm8J+Y255lpRnNlEbij0gebVg
hiCowPYNgsCqchafGsnobLBmhbfw1suq3qoIE/FiX2AI7WkQrIN7Kq/bOXSSub5e
WaKvcpn2R335aVzxlIPCJOr/nYR9ZkcX7Og5jmyGvwD67IpKQAVUdOLSqq6mH9Tw
9WNiPD0lundlvx7ZgAxysqbDNR27J9YQPI7LEaxuVx4KfzP7kC8y4IOvu430dMrH
/48ZjrALjjr94Y8td7kRLfkNMOrJJKRnGp7U5kCoMPNV5XOuZgvwRkSp9kAOXLEK
gZINjW9LcRiFjCXxYfNwr+4GAnFI+IbKHsORdK1WT1VJnGA10jva3Vqh8Uio11/n
YXOjCOoCGDcmbyfZaTzT7pPn4VBGdmnF+8awm3HIyyCY/YcjuyrKs3wnKTDmJ0pl
ISv7bmEf/kSj1Eo4OITlfJco2Xmp7jv2HJbksCxXxcV4RQbOf7Md9WjsMPMONfAy
fQ7EQOJ8KC+Do3BD3WpPDtdv0YhE0MehX8+YVA/qgJv647vRc42TbMQshuin12zv
EmlT8JjeNYjhjxO1/7kel4R1rBRCSt18GIEqmgKXcVhnqboSZWgTcznInuDJrS8A
2gJmy58pLdsLV+oLXEZhLTYPFM+6ekAEyPxns6xFd+wITgAf/DG1kWVWLXYquqPM
OXRVn2ShzqGQyGMXRpX/mUjylryrASeEanXbm/vyPZ83bY0rFR5q+JPqGtFFzMOA
xyiPjpqHfhguAuI8xHXIm8UODkvVOxkZzX2rQCvgQfL7ut+9h9Np4a+4mKz5RX4/
9QmLXf6p8+aUX6sKsOparmUcN599uj2+Ch1OGnwEbuRtsj6kn7+b8+05ivk8uL0C
7Os9ntMhLe1kFliigysSqW2UxWpqmtkFKL76S/+NhodsTNKHOKbM5IOC4CBLg3ur
IMyayqct6XK2gypSnqeBsYz+2mlZmZVcWuczfl6dnD5p/8Popzn+lIrQfZGCE7Y7
Q80RSCUH61ixclRvfIGqwZXJMbkJgn4+mFUDBUWOA8mKZq6pBYRhVNohfpyJbJFq
1Hu08W0Hv3obvO/A+oWSESgD8dWmyY+3rUcjPIoCeXmiJ4CZc/Gsxux2C/qdB2mS
8zN7zPXsMWDOfCIEWiV/KIGYb6RPSgoD+QIM5483+zJTjaZDVRPcuYZxm704wURm
p8GO7K5mJfwzUPIW50VdTcfYAPUPex8NDXuurCZG9Mirk605ii2tyxni19cEKbQf
YIy02PLmyZxE63yBiELE65QmWN0m1HHzXqHWXLEbhrd7RO9t40+H92zLbHPWnVLL
yz+1tu0psahj4SUoSY6UtPvVhpySeCNvC+0ydqell55BufMPqomtBlCZmRNo3TRs
T05my6eRr499DFNEKJHl1kQ7sp2rOqNJXAda3i8GKwYW05vEsf6/G9YVK/w9U6EA
1ZS3+HcIrGrRUA7c9gNyjI2XqVzY5aUArkLidvScXBm61IkxwXCKfwwNxbZ0QTju
mP0OIzDArf+gghCJasI557gg3RZSBLvSKDYmGMnTsCahOZa2xTXkD5OvS9Umuuzx
8slEoQ4HkVHRSj7zEc39Mhgvjw4qA5O7rWT0wCqnKaw+vPhpG0wPDzFzrGmO6+YB
N5dm+rNuxmX2uCxCjR9TQ4p91bBZNg23OmQPbCgia2ANu9COYiTMpcVtJfq28zcG
5eZy2szOwUEWLq0EVuFXPyuRESWMRLEhDcAFpCfJy1fRIVB0eQDYdcsJPJSwajMb
gHZVurR3Rv1VtI13pVydU1GnXsvmCf5sSY8liUVJJfFoi34YtPomyjuY9d60/fqm
Hdz+kbZLv9iCbnqzj5YE3bOJQkLZ0ITKvefPfZHfxOt+TrYvvBHYpOackSFbi3eH
0mrZn0yeKhqGS0LDMtr4yX1/P6xUZlETRdjtq8mpwOTouqDdMcsdMJCRQ09E9twv
yuBimAYpoJnFPmXDYjw78YYVObJjn+G/78+t0faWbzTAa1OJ+c2F6gG5pI8uuDFa
q6cFWOrLu0gngCVfuFl0+l929j2dddf5rM/4ILB5gavp+WfQLaShU6pA5g27jae3
UIymqNqrCajRZyZjYnVM7lOGjZgCccPTiTZvmk/NJVH0PyBxsdysHTbsBtpettBN
cANA5Y3q+EzRjwYiqEPZOdRcfjD126dZhKqxAQ9fwMlYGEpAoA/04kjGPnECLGA+
ng9p9r8aBOQQ5J7jI3PRHEIHRYvru+AUP92BEj+cVErIN/4vuHdL25dsXAP6Xc8S
Z0f4ooIYbK9eT3uvOPnTku06ALcznFugrbOP5G/7odaE6rs9WCfl4caqfV8zL6r5
dPnikxn+fSJ+CyKPixUOYfUFqbN602RK2uIa+lyttNV7yJfihC+g3Sstn1M4XvDK
tebrw4tTe8mfNdlSennklIAfPZ8n4gbayjNCDhDgIKEYgwU5ZOVrawdjAeRY2E2G
CohS1RqFztlS5DW1GuCo/lO0GEn0qH9Waqx4NsXrHdD4lmlIw8WlS+/WseMRpGtn
o7UswwzGZsl2Z6EspMaHEJlPXb1z1I8MfQXQp4oXelAS64prE0i7wDjMeO8F7HLw
290jh5ZP5HvPoMPerYJgzXyXy+ZktIbjnOa7YHHAbruxti9LUId6rISSBmzZ1Dnj
ABMsrsEz+2Acu6uj5iIFhGR2oKju70B21UqdhCdp25K742FcO3o1ay3bg832q2U5
RiTaojDLJRP7jkYZZnK5fWgm5tZJqTkZEGSu4lYbIiBHKZYd1zFyMK0YbEC21tVM
pdwEdkputIkp5PvFD26S9hZfbhzjFH4LfLW6H9o5yU/O2J6f5CcfdtnqoTsoD3fd
Fmiw7Je3SgkpPJlU98mUCQdAsGb7IhL2I9NtbeDpOT6VWrXoMDR8b5bCrhPK6f8z
BBPkO1vS+FERSVn+R1UYRea0d0iFtO6lpnccTf50LCKXUlsy7sIRiRKxxxmMtfas
jpyjRDi5OC67uJMGFYkbt12SMMddPyzDxYmwkRO2p41yFu7xCu8hw13kDcan2dLn
FScgH49lOzwwKVNTmnpLOU3oqcNKrnoMxlZl8tBEVOWicXjW+1gGbczQWpC4Amb8
630Pf3KvwkS/JcTX6DnzpbORQJmH3G3Nbq9SkmRExXsz26Pznx+aMdFXGUuK3f4G
dhjl1nA2nsGJ0igcuGPyRUEbHEJu4DlefJO8iYZASsToK5BYw/bYxGgDswfMzRXN
UVgUJJOoj6zYeLEmTlMGjZrROZPcL/14Pp77LbmbDLFri9S07kTvZ/tO2VD0KLHu
ACrYGWMHo5rVVWsg6CjV5FCeaG96yHJ4hxRPagPp6n49h6fx7cTyL7+dnau6ngcr
aq6O6uKoxmVGcGStlR60du7mOrXHq4bK+/oOyiDQYfUMEwPzpx+Xditf63fdliAx
hqQQDKgWkXxNvaCielpgDmkh8VrK70kRuwpJvRoVf5JEtTGDr8HMJOJeINZ3G23y
F/oRPHi0TScK/1gzZ4nj9Tw/D/XhDIJ2n1opBsi8kcCosCp9TgStz7TfedGat22z
oE6Po4u0UxemLnD5ZMLTCvre7fNjrC/LGa79lSdOI64Ti+SVivpzLX0uaQoD3kEQ
GTwtyjqLgbFMOBhFza6cyLt+HMTDdbaIZAb/QGVh22MLKffDrDSXi2clSeKl26ld
aGyaMcHg2vajclY1CtFBgMnPaIwH0hrh6vzWcWGbOQSjVbUcklDaF0gW29waL/nH
XRtQLGVppyFyY8g6noMOe2A6GDN6wS+6VGm5mmcCJu0XsGh+XG1ABw2bKJDhFCxq
W2Fid2DiWFUPS09YyTtYGc1G/3z7mdAx/4abev7x45MUB1UIqAA9KAx4vasMmA65
DBNDExDU32kIMoe6c0m1wCEq535XpPCOF7vGQdCKBFwbi1pcJ8dnFL01wP2VnsUG
HkGJ/E1c22y0IXYn3VE2L0naftcBf92oNvW0khpovtc9XAgVx5XswRIe7m6BvEgn
iHhBm9AiE0vRGsOsdBXcN9brPkcCK0erHffA3dVjOCR9bTS8tlNcE8sQyqdW87fm
wZIp1DcQPZqGrIdsstCAXgxnUhaM4wbLaqBn5FUtnk4bxcCzBr4VRShVggxEaC/t
4Vb03nrPSpQdowodaPKsvcnzwzHy3vKIsSdwjc4/K0qbE2meiUB7zfi+LOW+0bDF
w//0ogSvFpi9x7I3UXFNbYoH1A9ELIIROCFK3eeEnA1CDbhVE0Mi52wOJlKlxmR3
bunR3QNoYI1EzVhiVtCZVc/6grbhqNe1O5y31FmsogtxrIj5U3SvxACxHkvCHqnM
G56pq8sqoxFurNIWevE0LwECvUGHzBxX85J4FB2JrLGgL/NLVkk0qblUdbB2vdRO
Kjyi8QdS/q3VAa5MLkfNH8EnSnwZXQ10BX5MI70l6WbI4bIlepjf/9wmvfp4TUU+
fO08UiabrAL3O9DkSoyXHMdHgIDN5+BOxpIlRY7OK1vWHQXptAGwcV3Ls+IrxdF1
nMRQS4faNjg5oIt1ysQvSWyX/jmnJXgfLdjdpnomZNZRMYYiEe/F2uB0/HEQIf+x
svXjBhuPgRWGploMxxG8EGdBI+cGpeJqOLKbqRxsUT40QpmUa2FBOP40TElqBc71
foOI00Tk3iiTVBa4axKXQid8qcQd+SQSq6S9YV9SgOKRNAPbFhYpQo05IGTAgzyz
uXMGF2xdPdhA+lXMKkgiooZOmyalue0P/oWqQS9p2iUtWrujWY4sxQvtdYGdaEjw
b27Cmfv3JujfYdBBdKk2esUx8XOs+L49V95O+Ty9RseyMbCSFDazWfXUY8biLUc6
iaYfmwIDqAwnsZMvQ/jZpNR61dRQObtkozo98JB7ofYj+yF+aWw4SYacji2ZHQV2
+zQOcgrDqhuJDrcMzpv/jI9967L6QpFB4CZiNSWSF7VtI67oorz7qC8IkbxIbvQ2
3K6mwXn/LrOSR366pcbikwmu+6Yx5GU0zJzGpJEwlR6ulAInqPUrZ2t7MdYf03vz
wARZO3uyOp3zMA0QgQICSQBcpf/VHsF8sB3yj2yhk/WQzdXZpnh9ck4ikCJonhsb
Uz2/rscirw8KNN+ovbyFuJbHxw3ErkLpWDNm7mcNViPYGrXMvWTpp7fB4h8fph3X
zFLuLKWF8cGlBkf+kkTL7ARR7hltAhOL3sBz0axVMssq8pXugjUwrlFd/bm5m2Oc
EgZnlpOqh/k64fClVxHecEhzmCilyLKmmnR9iLO+OJMW3kzxyijjeBpfUEpxrYJF
RUnUB+6PB/ehN6dnMphdRlvks5nbzIfVfXmvFuyGo+6QX8jdyWZ+Rj3MMgLgBjX2
g+EtJaj1tTPWU8T4irLA+05WrAgSqajjswNTTzQWXB2pbTwreHjxBL9vAiWHc6JU
8QFPSd5xwrOa7T3uAd4wdXSfTXp5PiDzwiiZjFnR1WWGxnhwwGNHsEjh8omZEPPG
yUG1cjKHeLftGqsnAO13J7IvEpeSSMdpCaf1S3WOdJwAPoVK6LPN32CRqYssui7W
IhskqlSmoKvdSc3/cxct5/A2INXvdimYvZajwaAA2hShF3yZiG5TPpdYHbKtidx1
PspqK1M338Bv9RFDSWCMA+zmF+yKuaYIDK7yUNq5bsSfoUx7gNYvVsYPq/eZnL8U
Q2az9zScr3m0qfcKoY0Vs+W3Vz4FOSTV6mwj5++GdtRX7xs11jxH/cyxdUUTd6OS
s7WgyKybrrikHpYtHuTyM5o7C88pDvnN0xurpkNvWNxJOR8grJuaRqad1w4Jabbr
6V1d8lTbgmKxDIQ02srNKFsSpGKQS8sNEAmX+SkczHrBAarIKVZsuJqG5SAqTlBZ
KI5SqW8beFBva3DoJ3eERKX2N2QQE+OdFCYUHO8TBYwtN46YZbUm1Gu2BNF8oNMU
62+VIbI0KOU+I1o8IwmnvLMoyn0vu3nhNeUGGCR4zAr9mSTWw4KU24JnacF9EVSp
c5hbVXdmsrU0QZCGS4elPDce+0UncoLAkg6KWLamWeP4clC9ZAWv5HesXUifybqk
M3T/AOOHeWZQUluQ5hntTHxWGR0R3bJ9KkE7WlD/XDbgUH1iTaP6Xog+eihAn607
zexK1/CYrlscxKuGzagiZFkunnfBVpEL7ZUrDYU/Q/9ancmcHfV9OinhovjmqjWn
hiUuLG35gCJOtGmpW6Gk7w31AUvtSiU4AtOKmrp6BLIiuIT7hJ2Q0NPgeEuMm3Pi
ezyGLeViW2LgitT9NYybUkGFqaB1wUvW6DeNbVrxfrTYlJJufEam+6egpXX0bndb
/6p+SIow3iFM9tnXMhraWh3ibH01HzA+Ak7OgJUYKm31LO2sCkOWyj136dU2SP3V
UuCbT8hLD1FDgijrpDqUvKceFtDPl0eG1FIk+hlQZNLM8X+QfuwWMFnwRXQxMVvw
6Yl2GmJg83rQ1IpGNVoJ3AaqIQakUQtzXRSLnoytU1S01QMzIFqIdm8M1GqSOGbt
0aZn7+O7/PtpLx2N3DXld/40AIz6POJwN2jftgW5jvo/bRTsSHkKj5uIYjqcQ0BE
5BlhIJciVeuDnD5/bcrww5uBJ1stWtuDfAbgImjM1JE8xKVFouQWa3UMec1cuNT1
Q2+lRUW8y5tpkkNWvseUgjyqaD0UPjiNF6MQDsKzidFLjnwC5oFx+fbc7cLUqE20
eS1bzUcPd2Z4Tifk+S1LbFwsF/LIjET0wh7uz7L6+y2RwzLOLrMfALTfIrOWZezw
cYo3cXhfnBb8lO1Gp91L54djlvERoqqLntliqrx4XPG+8TdwNSkT2jGmaYCv9hTM
709bjkE8xANPOuBzMQWZPHOyyKZ1+7zaSV/SI4JgX5+bAYtO/+2sJvH1xcPFe9Rd
4GkZlIwTPUwP+gIimrqrYoTJTJDoQmHsRyPpn2NDarhf6k4Uxa69y/nC+jjtu9LV
BjVx28ObaJ8NCdxVjb2uypP5qdt2halBoNpugs2re1DG0wdMuI7j6411XjMkymAV
EBvJzyWj/Y022NEkuR7xsHTqwHnfYAyvlZq8mfcORqFnntq//ECZJUW8nqxw7pS2
zIpcySSIS6TCd8ZFUZKZSzeZoQ21ro2r9/ypXDpAKGkGLHqHW6eq9eh3vkGLgs/P
yo2iV3MDLeLmlbuQpd1I97slGvo0DciYkN7s4woxA9eF5XDNhzFxgIw2u5jKTcaT
SyIL9wBGfKaBdMn86JYe8FjiFVkhLRdbuSnYaMLI6Bfe3ZBNPoXLwDmlFySM0+yJ
j3yvRuXYLIDdXGWgAzovQxR7oUNqh4Qtu8ZKH8PkVFo5YkMrashWgYz85620maOU
5I0pew8FIU9RCIvbed3Dz2NQ/9iYgvE9Z8HKkKkezhDC78N0hDZkS3j/VxJbm7ez
u2dpapkB2OW6VDVbSaqDf1aZPr6e7dEJh/eVozTzCpbOgfjhOp9E6wmTzEnvU2vU
a4MpuXdPtwn0E3lQmvTOdhygtxY89LJrs1N9gyb+U72L58OnBlckFqcwHLaAy7AY
c9pppjI84bPPw6uoPSMqfuNgN8nq+Mdt7EvQq+W2WsFhVMUbejcCTNWzFZQdE3Bu
AtudPPB46CLr5AlaVaZV/QZBnWzVadteH6aveY5w+JQgrhxDRSC4rHpgunwSDi1V
0ePyQETVb8fz7epvwdfSVQ99SvCy6jDPlFiycHz+jmVv+fvxqM4VQHQMLW3JEzfY
s5oSbO/wZXOi8Tkrek0oFFXGTZd2AgwX/r4pdCZR3cikoFrOQpbLt4/zauVKk+AK
wwfsrM3lKBjmpo7NfyoAbSZer8sxmks8J6LZQbPP4JpcLvkbk6EH33PzYsFMjIJ1
NasDBnGMQY0fAopzq9MPBb8iJSbtiPYQoaG4HKUNLi+yXE+JTFCOnkqkcvsnjUPf
JXRUVGEoLCPaW/JlPRsdk331WgmMFoHs+lcqGIZTs78zsrjaMT2T+4MkT5frvUQF
mMqCuf+AfcCU0/UDmb1tHS4rEHLQA2Gd16eXbV3fU0hnqcEkiOS+4OqhwkhFq5pE
9tgdqAkbstD8bGW4zSljpQlUgIdhqJOCjQmGUNk4ba2XKY22bixkD8euu0lDSQcP
Gma/Gbp0cjFIe49Os74jX4PR4bp9OYaATVY1+7sU4qSZ0WxulVPkzDD6hNZc48uJ
ADTG0mnoH2K+g9LPUwqIHYceYZzwMKOrXOVVD9Zya43oxkL12iwgytOGt5t1p0lu
jnoXWwMTVTYDz5y5QjBE21FXxoCZfF9IKnA2QecM5nlUBmpQuu+0aPzubSCY3Ys/
cV4/oPIXcYNmdLhbmE2yXts3kFnA/JAtrckdUuiUjxg5flPFiJK0DNCEkSTgt1MD
XrBVhkEs7Zrut3Lfe77h+E7OONZAgSRLjirWIy4cyP/gL2W+kzJN7yzPKkZvmo8y
pdi6FlrxtlPFLkmFJHBHn3kU5W9+ASJxltOIYaQyS1pFlTya2XtwiumoGRcs7zDd
5w53WnmJhoNza6IGNhZkMyjUtWjkwBymSCWVhQp3Lli2AtDx6ERipSea5xG0knnG
L3zvFKKEbDnUlW77nIbV6FCkbrtcgTqcsVg0Rky4mdDg+MGX6lPrTFEH/ArM4Hlw
CoDOs0bDEQDkHJGO3ZrnvabG8kx0oLYI5MOi8T6X5gH4W0BDEENM3BkyXoueeAAA
3Ab5sHHphzhnOBTVnU5zSJknqz3UkAcCbylYGLGsVHCdMsggP5fbkZ2fCIlAuhQK
HhiAapxW/p8c9KyNzKBN/lOTRP1HmW3O4PE9Ux0/FmjxDO27JRxoVa0TaP63L9Uy
ZV5D7nLi9mzVcRJC1Dloh9oSNbmIMF0L6zgDKdc7OYhRRJon6YsTLNpJizlroitI
MMZ0CR0B8xgPWegMmtdYJUzsmkRBRAp8Ii4NwPMSdWl7tRMeI1Dt5pybXkW/sKst
fWmhqc9l9e9bA20WhoGmskeWrTSQ0YnTUsK6F++yDyz3PMXlbixQzt2dyC38VFWk
8n61HhVSVPCXAE7wVFQcaFCgF/31OpFJQgxrEJR8Z6l+hKVQciF29t8ZvVEP5oBP
r+gsUFCZpB2KvFDFjWIZLkXXj5XE+QrtzSr0n5Ed/9Tk/4MC8fLzqaBsxT1k0h4H
v+YF5yP9HB1zvYZuNRcYFBGiirsBiTU2BZiZcwqvKGxSfphSRJ7s2f890i8DzIk4
on9tI0qJJfv6PvJAs+YdWWzCvVinPJ49O04Ttddrpmx4idliwcozBQ9RFTaP7NsR
NUflP/b2tkPANOh9BDcE2llgm0ROT9fx3TMeK1JeNCMwDUrJUtxO0q8lu5kpvwFy
Sj033P8S8be41vhMEf5v2Ya/F3vZsmNUw1ZBPSpkYq+h8lJVLViHFmvjFUl+dhv/
m5RiWMK4/ZTYK7mPow/NUPTQPld87y5pqRHkd/dtVp0OCLPayPqQFpMb7+Hqroni
6IkSwq5QINF4GRjcfZdCM12r41huLbcM7cF3OP4muOGGy15z1TNViP2IuTUGex3i
sD+zMGh5KV2RSeoUSEh6rW00Sz7Yzmr28YNccGsz2RlzoJKaH8ST99PTEW09ZY75
ZujcZo09VDao3TlvuQGMpID8VV1Pid2L5Qz+Ds5kXPi7lfe/CkQcl3S0ZQjM04pl
kLo5mYjgQ/Qf2W69keUn0g+juiB1RPBgqI/lP7Jypk2to3dSK6Qwig3EcDDYHEG+
xeQRBHyoe2jS4kAk5G5fh4eNoRmv14B4W5WG+QTj9ftxw2WTAgPEPTHfUcnQx+pn
rwR5qcVEb0RX95J+RCDN8LTQG+ddS6/QuP4vL6yPSA3c3cpvq6oDXNdEgrARUlrg
UP2XUX0k2xInu8GMOQiPhB3InYzfm7KkPNKS0M6XLmmGJV5O6eAJ1KSDYIyqIoPr
+hxzRfuV/1VDvRxL8Nli1y1Rn7wb5FXkfaoD/s7FPLeS6b/g1XYO7yyWgj83KFMc
wy3O375aQIRNgfR5SnpcGvFFCDZr62AAO9kkk7/aMyro57AJZMcT08gG4teUK6qh
rr9uovH0D7+dJRyc4ZSLVGv6R6ooaWZx4o2MAtSmTBdZRLVBONPBv+/nWR36Q+XQ
mcBlKocDssfCV0R6T4Fx4ql4k05838hFdaDoZtDx6bwcY4nF22iGkp6WrgmkcynV
zIfiHNKerusmvMUVx/JS71tJecQ863a0/I9qE0oCRDDgI+z2wdYT6mHIfA1cTTw/
W/7E+fr4179RdLGP+cXRCnwc8j+jyMFZ4CqPSr+HUuOd92oLRW4gnejVR6xSdAyW
wr2tEeV1tFgKh2Wbb/2bRcLYz9pmPuzWGm3v+3daCNaMfoB16j9BLkb1dewAINYe
mobVq4sxm7yib4Zkze+VpqhjH8lA84rIRhAYg2S3D0T3fq4Io+SMfyQJtzrBvHtm
bTpJQD0zXwTcDJRPcE/Mokvupdjoqke+/cZwpvuaHzXZfpuTk1MwT+zgDVymttrP
w/45H0nd7VQo/BRIwxoMS/zmBcvsZy1ngZji9BiZMHPMxpnrDRCvIk0/ncmE/BkQ
IQf9nXF7E0vdHL78fK2GZgXTX2pRGAxqYNVkIGnY7TWyuH2hpRvbs7hH3pEH2l/h
/XbG12TaWWqMeOqEIK+cy/zhSdkDLB9w34G46ov3T4XoTOk1vo7kl4UM/Z9duymZ
+Nk0qYrhoqhoMZySVYwiGK+Oto17cKuSFUnHIPhlZIV/lfP9reaGNi6gyvY8tkFR
AX3aS+yd7q+VGhWPwYWkYZHc/viNeSM4/SbDjwGuiXu5Ym8qw53la9HKS0fv+T0w
TeMvJTTjqqHoTTv3rEFpc5JbCcBSHoPW9cHszfxTZHF4hBAqBb1k7WgLFFXrSB7Q
XOfD0bNoo3tZiCSzLUCkEIx0xul5559AIx+V+GdUUfP1EvY8wg/aOEXL0xleNLku
zrVAbIVc+4mekREDs0xbzRwYzewqBC/fvSA502qPgVKXZv3XuVof8RrlEIzJOpzW
jbWTvxicYzd+hoffmhYnuxvZfdRQ5I9hq7N6YJ3U9Blif6gGJT3VzvwVxK377XZq
T7/qq8du3bimxxepMeObEAKiXyhdcJ4HLLT6a6iOkroRhtCNd6wpzu+7jOdsaImZ
MDVFVDY8murWD1U0wg3IYeZYEJI/9bC0DdyTUkKycZNTQjLR0SbEws0d+UMXl/cy
2r0icTiXN+gzR5uKenmzyNFElzfIj6hrFUyocuMmJcqLBt4cXrtqBt3qjm2MUOd2
r9kbGGJpe0XIiX5TL74daLWipEtF+sMAU/bpPKhuVn8TaILhoJbwAoOvRsY0Qw5/
igKU13WLJ9Zs21bwb5lIyN0Us3jnfd4+xERAOfxinonRbVpqTfIp1fwrbuWBh0VA
m0poJTDlE2fWof37sHqvMdlLK94wd/TFLzLlTVUfooA9d2kE7cycTxwLBobghVCh
5oEM9+UjkcQ5WmSoIHL5RXVlSzjs7SxdYgNCXcTRgUFu86hwCyOytUQdOkNc/kuX
ggORy10g3IvYY37K9krV+87VzbsLq0Bbdt6Av1DZ1bH7odgM6rWIhodCGahA5zCM
QPZsTcHlqoXVejVuFB3bQjsTc2LXcdMOI+hcMos/Qxtyp4WFb3nhJaEGf044Nz2c
mR5fXuIzlI039RobhovSu0Rkz2cBwifA/C/eTUpf8GhbvFSdp6sSr9o4s48QL0l0
O9Sf+LHa2USpPxtzKNVicofIOm9oux/ILkwTUb/9xD+/wqTxqP/Ba2SkSJ+dDsfk
ykOxbEKNwWXzZctmdPl3UZRQnrHQo2yjYZ88WYAGD23H2Y6EDNI20Avgs6BTDOZm
lj91GWGenVZBkXDyzZ7ca7SRRhHhRqiWUNae7hqSZvBIKz3kAw7KpsW/xT59Zujo
g9ATVkJqkfxll8cFulfE+SA/MaZlRcuiH2TBf44hvrAyGbt/2lVCn4Ik1T6fsaih
H9AluubQa7gun3jBVpjTCN8C4uwdlqzoFfA7Q5/JU3lBkryLo3vT5HD/03nKPoMJ
hl8j09mCmTTMPI/lygYVHI86p333gLualS4+tvOzuDCtyTnXu35GmSUMhjlePNd+
eiOnqyjmiJEMtIt5au2YhBkCQvHyafpZrDoj9WHUXjSn8MkiO+aAjEC81oKqhUiM
bPU/vhgWZOPjRrL2vy6xBg8QnDg/GYO/HlBvnPH/5atTfdfN9yLpmsbJB0GRVi7S
E1H4PsRsPi99XjgOElJI5EHCiPgOiANHEwbKl0F1t8anc5PT501z/bA6vNMDEhDO
RAmDZJzonpz+Lfj+7ZU98FkgQmRjqWPJAuYqKMGpljXEjvpaxNA90p6J96cNEDRm
9nL5+u30qjndR2UMSC5Dg7k+M/FcoVOb7HqtySEqOzNQQyHSdAU6XYxcEQCBsB8K
iEL5MMjnGn4zA9H2DDXdMB0yU4A+FjrjhpJdIPTwHrIHrgPdQpSMiWYVhiWh41bY
0j8ugZOtV7EddT3dCM6mrEjuqSdDp+oCpNE12OePiEvbwiGFkWpr9RHuMljwFjYR
ZmWuOBhwVIVdAY91rzde6dP2UW4CuyWlMoUQlG/rtz5hSWJEXyt7eDQjFftt15iS
xlOau70rySZcjMg2liyAoIGXyb2SjaDH0Vg1vFqf/KutBF0gN1366sMcqQmPVZVv
8XnkcfHyTQj3zDdfIVaktn5FJanvUaTyKbsC6EQjgneFz9GMCT7eYWS0tFMUSfOa
qv/UhW/NvMzjf+WGKhjibOXx2GmWNbLAxhA7Jj70FAuoUWbBjenoq1ZRT7cN4K5f
mqatTBuqo6ncKJnN3tj4+dMFavo5VQWwpNBPGTh9vNqDfojEJON3KpN8a+iz2T+W
T/LlxkdXkXsqkAAI5I7hubrN1wLVr0qBOLCVI6nCYvhiyZErj+uSKB7GHNKq26IP
pKqlZZvFU7uQ+p8KPRvt8lBN1JgPFfTqwZBB21kYETfKSCAU48bJyzZvfQjXsCJm
3e2HT5coI06149TGI4qEHnwNd/7QgwRjyScgx80YDEPieJaD1AxLRBsS0uwqyN38
xMRZMYn5zWXL8px6dKqkharX4IpCBfpQ5o5D+f8VV+26hNx5+SI2fSrMHkupbhAm
gKKsP6tlLq47hZxoaaSAPfOBQpzfGfcCcOQYmliCicONr2dqQeYt7CAicxtF1wxw
pyK3EprKPUVctpzDBgZ/vDKCqHrp+cn96v5UjWNGgFxh0HE44a0n3Mtu9CNaZ/on
PmSlapzEQZ67vlBBzVbZdezjvWRVoz0yH7CSmMWLwACXR1yU+4+k6dKCedPkIUME
98Yamnlvg48hOjmlG3r5H8mU8fEXXSpOvconKSrxNgY6n5aLKw08zs4ofrgomo8X
Y0R2U+CSJKbTWaUqgj040cpsrHjac3So+Wx86Url3XBEUnxYWB/ruDwmCLDZ9Cg5
ezGcz4l13ml0GRpq0/uUrwtN0n9wvV7NcAUYSuscIEGc+uASLh875VaSiYMKfMYf
zWZptHbfaWajkMY0XSexHtnT9n1KPKOH6YiKwZMwlZeT/u0iehU3cTnIePJTtcO7
sHxWdIl76Mt3KIFu1snkrj2WnbJZnOoU9WI8AxVA45SfF2f2XB8opVtFq6kQDxzB
NcJb/LcCQIb96j331JIHn2Q/xJGr8oYZCsgm86zTnNnq4QjLqcr/avgJPKY+rV8O
cTGwaEp3UDK5pn3zb/oRXm7byHKyqCd11dl7r3/JeCTKcDGMslxm/+rsYYCnWkQZ
gKBa37uD0DN+U7xPwmqGnUP+AqeEulN4tMYVYEASaQ3AbEi4KPB4iQMEUX6y7tn/
59KShyUc6a3rTpNZcYjJ2LkPb3gGnZmdPMlgDKBmiKSXfnir4Y5wyshWsEt4Ry34
SKTxzBYLVXBgXSQbmhW+KUOhviI85rGdd7v+X+Xt6ouUfNlB6dyZvKbLYcG9wsS1
2qOdWQ2oXof2oNb0eiqCmEANgXDy617O4vCOED1Kcg0EhuSMiuXa7Ekmv1vGRcU3
xK8NEVkVsFiuEvFLWYx71AWMzBkpUvTQCdX61rnuEa2AYGEGX13oplD9xEw2aozR
UfO1WD9VYiyGbcSXVX/WmuXgpf1lFW+tQWSZ8EGjSywQV7XFs56M8amMzYbecjHJ
zacqVrbcZGXyJ7j6n1m/CqwTVvbDp4J5lZiVLqbH6aQCLXBEBvJcYVzhj0P2CIqu
dH9pAT6nK2lUTn31IDd+UikXwcci6hjqQCqXA95m8sCRjSMEuvkb4jl60WIN2VG6
Q2Y+jkuzrDwnHGKvDZbclp9Zj8S+orZ6jTKJkbunH1RIApz4soMYxzhE8PBJLcZy
cSiyV0ZjN99OAIqqzJYE1NLzXIiNhKHcYq6ci/itwnabRMMgaJz0k7YOySNuhxmb
PKk+3ZljzB/u9WJG1VFigaNZ2Xslv+qa6Wm9i8sUZYrkgJWji/TZcmKGOZiY2q5a
crl8vSSADoh3cRjC0chYjtVPgHaoEHa9d9jsycCOk7OYMaS8mQPMoC/JMvSR9ZAy
B2wXf/A5lu66clcvUqNmkW6v2xU+rZIynibHGwzJEI0VxqK6s78FY6Lm279vZJpr
CojrFNy+Ugp1PEWiEHExBKvQDnRX0t30Bzyk0oafi6ehktWOoKxp92gv1f6yAFwK
1bL8MS1r6H/3dhSXWygj17JjmRMDQBJu4YwD43fFW1V2h+uxhyP96P72/o2l7wvt
xtCuA7SgTn6vTychhNt67vqdMtl1F9R8RqLVgZYjhjaq/rrF4YIIgdbnPZZ9Wzec
W89sVQpvBMuV6ir5H18LR2xhBWRLo2wYYNk3j7RD041BEECGwvmzIc9bTNvcpZMZ
dorafbslM4cOjgDcnrkw0r0bsRLGPFZDBtxIeJ+8E5RTEPWVEQcKo9I63usCKMgO
MDf234yk3ZvaMKWiD4RwlURewmJi1hvSMzhR2dxlIzfGlVEgshTHCObLspHDbuK8
AHeC6RpTn7qZ9cNgL03PVJ+8gKUyOSH3rdSQG/VbkJ1x2tioVZ6oMOFl+zOTP+qc
BUBNABICVo0uSANPWMJ4m72AVEy0xLtzbpWcbpoJXWHfbYqkLvSUqpujUAimM45y
WePngzl1Tw2h39dMo71rFCAwUlz37Eo9J30F/lwj4adABYpp1/7ode587spxTbnK
0e5Zksw2ecA7/iQIeobTZf45PNrTBYjcHFiz7TmcjP1HlYEod88H8q+cqADekxJZ
205tshxqdih48v8Idb/ExGJR6JygIxR6G9/FcuW5t35TSy7l+ho1CxmB+LcFS8lM
jEVjdsEPKs4aFQE4Ujb2sNa3hCJO6bTECj5fn2o2nvKg72E6/I8CJZBov9vxH3CR
NBvVBeKgf7pCuPsjwiYYVkFzCgk/wWOy71YsDsC60CEbUHf+IYUdybGb1HoNQ7DC
O1ZY0rks2coqlQg+E2QgzegdedntA3FUis5gj+7ekU6h0VxTq5TAaXlJou7JO/bd
WV5bB2iV6UtUWNPta5l9K5Ybf8wwbQp9gxPKp8ZMQjb25hLjJnoK6oxfai8HU2YK
hisa2G0LK8pYPddlrqhW+mhL0WeBO0t5uQe2+mSZtWkwnuYdIGze21iucm9CeJ5a
z1vAtlT0WvFKXtSyYIUh3KkJLmUAWYORJQAJgmjxgpoMrH1L5xKBEJl5ccsg8aLZ
dGSb8T/49SXF2yeKrpbE5O8cooOhROovN55v8zKzo2Y6Vp+wbIP6mE8m2dGM1MIZ
PiE5LQTmnPm+Bdn2cGSAd6GfC1Pfygr9ghcVCORIwiCGjnVsK/P82GYbzbARzHsj
gqS++6gAjUbQUIxIXWTJ2FniYt9ILUfJ+px9gnk5mD1+lC2DvI9dfiNM+PMwwC+H
sQo/867rHrzuPVShKl3aT7jLtDukkc1Sm5dWaJFsuJpzwCI+LLMBWlmPF7QFb1Tt
za20+tuDq0L5Zi4TX9N6iiV41BEDHfGkJ1q/xPqggSM4VyfHHk6vrC2VRZ5l3mhj
am8xiH3cjcllsbTobY8kJ3OcH4rrTIJbwv43DTKZulLtFfHAw1B0ER/hj48KMzeG
vKECcr4DC5jBgO55p3FDKRxf2wrf1LZXqBgxovcnlK9nl2cy2ztt+G9L4MolYbmk
nQ5wfIAZw2IQ5E99q6/ymBq7QV2qkmGCMzjI+4JYPiRgufO53GyREqkdnrElu8/2
T9ccreOvdW9mVdJ6dtlJ7b8mqfDcH13qFQ9hGCVgmXCm37RBl3Jg4Fu7mF7EyuY6
Ge+8BdztdxwuU1yHKUb7pJxtwv7u5aW+eBo/hv83fz6BsgFM7sCVmjE6J4Y8xGBe
/xSJNeh1XHvS8fIO7HDD2LCiaUQMBABwj0LMQ+uADDQ8E1KQb3ZnN7mc8RqdhJAZ
KPhSP7ByTb2HNU4bvwG9WxpLhIrxHNX2KMPIOsUGYqPyeLp9UzylPivUACo4YY+t
JCNfwTpAoooSWnSCR4m2Oj7kR7udl5M/yIKnCSVisb6oL0jlesEQFvJL0oAjMb0E
iHoIbWBXTIxshr8Q6wOoIScJUJdeRiH51xF4xvIHaSKCias6b20iPYYqWgrK/4bA
7hViLAmR/IuloeWdjvLwb2OswAO87IdkMhaCzFxtY4SQOxkMT5MvLT5PCsLsYuMf
Yf8HzX54gwbW6Bee2NtQAYu7/02RqqWTtpbFBGave1KtlMVX6oU4/6IBTtYiJXSE
lTMQlQmcHAvniRki8w0nhiFQA1sKnIyvf2B7neP/aOjkm63dKkWAi71q5NVHR5Hr
x2/KyIS5Q7Z92J4qLK+nEBVwAmqqq3FPfiHnIIofV0B4Nxp5UhiTCxAWhb2I41Zd
2WguNmQ8yN//8GlJPvg/DIRMl0AVIC0/vxK3GgYJxlGvCujZQ9gcQQUVxNIxXc/n
FVUQ9nSPaaZv45HRw2yXTOJWH7gibuhtGnT2MmCP2815gJt7GIHORKLijgtrPZ6Q
txyT3i9JHC9PnxcMsbIVpLUVIZLPdVtvuy1aQWZmD+Ar7Avr8tDGMb7jPzDNGaeH
2AMiObCUqbpFKxeq7R67fTvncJRHg5pY/LmKGT6hzndBJ8lhApWlarnYEgZAP/j4
xJIZ0KwNbrHULsSdKokZT9ky5TwjsD1vfT+deAUcZLnYr+kHvijUzd5RiBEvXzC6
KwGPASw0DDparxH+k3lCARcAx7nrdr+Y8CbCBKPd3sxzZ3VEiiuvi06S7TEyNYCj
hyHiOh2xgwoVjKYYWmBNNfgNfx97fiqeqvJY/gZuQceH1wFFENutDpcolA+HFK4f
AHRPdXxFv4Me0Wr6gGW5Ood4u58JBxJDrNG7E2t3T9vMQkkvB2ZLwi/RRjnUOySM
bbZWeSp9mvoNQ7o+5OdkgYCcKKJ1dtn5urQSxUaUtyaED3BHA1o/7TERKHWScr34
3ccArvlQr49wJYjbKnJDZ97p56l9yNgdHjkPJXxMptG4Q1jPAZunvp9D6+plDI6s
den22rO/YFzjJ7aKweokT+H7HE8E3N78yiZtuNzUiEkO5L0A3cyDCtyhaGU99Mzm
dsRwj1o+gztFz/XKOOfR7yfvWBSCPD5LgeBl8omA5WHVR8CRZ9Yf/0FFxLxWG7/9
4v/ipNtIGfsikTLOANXTkbUVlaGNeSbKwwrGdqf8CVCPw9IUNd1KiTOx04C/6UJd
vBbOLV1jDbblDT7VKrot6fj3gfJALkhwJCELA3a4A2hxpvjlOLP2cijqBxAec6O6
QvTr+D4voSTEqvAdy0hqNWT2O4N7hb7UF1Rs+Qvs7pMMRZwxY3XkMzwHt+hoFyZ4
d3t0w1M7PgGMLQo46KqDmBhy3qRYZb/BHaKFyIeOc+jPZte1l+YOqkq1izuso2o7
W+7qexWKhWM0VGm24p0IJ30NVW1xruwWHTBhArMnkiQZ6a8dcUO+teCjKl2SffxU
dl9FOk7aI8FXr7yIKXCwySqn9XDl/91m4v/IDAONcW7BUd6dhZXGGY8+Z4SggLdD
Ukbl/QqW/cKAnSIc2D6fT//4frccyMEzhkwV934Y2/qHqu3MPvzFOAPsMNUvFR/p
OjKYshk9aCQzUqTb1Lyj9zGXK6XKJJKeJWrYQEX+IV/+UVBQV0GSo3CL+gJPAw1F
rMQlUzeyqKRmaZtShfEtLmFeWDrZIj5nZVvMkTYU11gbJBAnJqHc9srHaUUSvhSd
rJYSgExib1hI4P9zyAAyOGFVDbgLKW2/fc5xQieTt6ttxCvcXA4JnHEOaDId3+r0
yZPwsW+ff/M5gAPJtRcU1B7rp0ccU1HK0Oc/k9nZ3Vq2KM2CTMzdHIp5T91skVr6
vWgIOfqB9ga2aNcy+++4NarEkKAJbiN8nYFOaPYQ6o8Gtat0mDEtlcToYofjIkdM
tZbrVi+DTaotYrUKXtAjfVYcLZO4eybRyZkuFYEBjEf23EaGtdhEnBtU3SYtUtNr
4gVmBWsx5UFm0+4zNiFnWxnkvfioiJ3bYrxVUqcNN9wKa0KW9ulHC0mxdh/16nFs
pRJZFnWaqnkuSs7sgKyVgAz1Nf5J+4K2ayFOeMKfFSMvE2yJK3z97b0Lbq82khZe
jpK/8v3c7sU/2fLjduenbx0H9c2deObbrdj8ox3TbGXAHFOs40Iu8Hn8XjEIQ5qX
cmooN2aIzxWHtbXfH1q/FnSDWSzexX00nQ16WIDRZ1jyV/2K1/yJ6rhQpDh8YzyD
uLmwAW95DuU4iOEGMaGK7QJ+30xACZu93Q3jjhdKB/oSiVxV3F1vgAJOr384wlZL
xQS6TAjgJM0S29ragXYA/Vp7pzLjdEPsUnJwamnq/ub95Quw0dN9LGQX4hKvM12l
hrkxIdNhLLs88LEWDx+aSTSM4bLsAO1DWlxS3rnkorex626rjl0NXhRHdDEJvN8U
yJVyYJcWEr3+mdFYo4Q80a+7im+6bF5fX3HSgPZ8nFSMqbvW5uLq1uWyKG+uk7k9
WSd44ayzlUHfoQoA3vEpxfp4iEaKMRDSGsYYro434nF5CqQSPWtAVxXru0PVpkyi
lFFWdPo+uMYC4OVDpiGeG3zMLCTomy3i0TgpySyferAYjWiMhkAEkH144XvHqu5O
ij7hauIZBUxoJVGMFtbGRdoWABDE3gZRL2LdejaDi5SjkJD8YujetRZTDRlmVnVk
Hgw71QhtltA66TF8a0WqWY64vMvA7MfaxJDLuGKUJhXOwdAKPVuaWrlczYtd544u
GZN/y1MLsrEO/Fucv3NYtf8dvh5Lc/9GGqM+umX46kt9gHe55b5v61fglRcWu2NY
zsL394tNrwovu92dEVouzbH3qEuVNszGs58kGT9FsdjakSfntg9Lj3kgAzW+EXS2
r0ahXgvdJBoNHRM7VTePj3mCXSi8Q/2xQXF8w7fZD3NOIEXDo0wGfgiv7ruCR+dI
gDCbrLZccz3/c43Xzyg8BMlqKBu3Y9mArr299r630or+MXzv+KVnrAe57i+sFe+j
g7EHi6uLXE2S3SY6qcr56YkCsQbIxa/K58KC1Py0JwL53D34wIp4ewE+42izMt+d
Zx7Fas8XEt164crgL/pXkPPeFo3Wex+AtcRtgkJq3A+sUDK1d6BviPtSrgZo2hv0
Pr3ucZxU9A1CGvXccbavkuExh3nXI6TovDCjsouW6/dyxH2YcnIy+M3u6npH8cma
3b7q9+MsM04oPswx6EqlEqy0oXK7TnZzjWEO6pa6mh9dgz2m/0gPa2K9hfUH3K+O
Wa+ozRxSziKmAGB8VrDprnjKYJ/PdYP4gtDBCMwYI2N8xk+9473jdOs2BPZ8wxms
ttTdgADH7EyyLNNZM9Q8fdOWfgh97t6mcbjIKZ5622NP8kPTXwrYgjGcBHGgyOrr
7Jh0dB8xDYI92JIMJsatwtD+jEGO7fs394JgLMf83VXfrZ/kzTWGpwlAsuVY/FTx
l2gXJncxmPdgyMZiQLFy/QjrDtQr5pakP4dW8djKo9rH5GBW3TvKi0yHeq30jSpm
Rfr3ZfxWeeYCpZgdyEP678h5kYXwasIKyTlI5TXRMFH8q50Oki/W+Bc79HbTsk6u
FnPim3EVJI/en1kesf8dSVekumzzlx+xlIL5VjqmHRmJigUM36/6B8c/SU0iDY72
UAl5nVGJxGvR+QxGR2dc8j/oTtr4eJ0asSu4Vvd1v4JnkAgA+MqPcb9rrYuMBJw/
yZ9zuYzAiybdB6zv5d7/cJuFTETyap4tfe1Yicwfg6zvuQEL0348fEgA60DNNaeW
3kTkGCsZP7hxoJHAQw52thvNtWAwSGtsixPtwF5cWqNdXVdBKKlW8tYbEblXzqNd
JHzL+93sk/cBoLta3KbDFsYj56vcvxTG9H2x0GbG6xmYy174U/MIomwBA+dAHLe6
70yYoWIBFsaBU7lHzEtcgniJlZB4zSmSB2H6k7icSTihcSSxPkxXc8aXBcxOZQuR
Qbs+ifytGM4z7xR7U0kDpzgzNlaOAVtrtB2toaPE16//sqSy7hMrC7IZ+2ClM1uP
+YU8f2IOpmCjjPgR9kvqqn5PrtmdPXR8UMwnz8sC2ZhPLphT7oWyQJG+T6OHOhjm
Y59Br663XOupqNS7RnS7spRevkFzN2/MY+fckiwIP1jQ0IhLyaUA5KB7QGSHTcdQ
6uwAFG4b+FIgXfU+KRHN6IE3YTJW79T/OPF5+DyIldT/sLb3p2VPpGCtNChnU9bM
PWfUtcHvGstowcFz7gP5z7qt5Pcfzu06pqrCLF1RWgXr/1VkT0LMjdgEjjhRuL2B
mya6YpO8znPTZld97asaQtJeoYN0QnOI8jg6sUmdcl0dFbqhnJFprGBUnK0prUMr
hR5XarXUo90wIkv4uLMteZzEyjy/e36uXZ6q5yZ3b9SNSvnS8L/aQJQyQ/zVNBij
EpUCHMtWpAnLxSawdp4186lYCU/9JA3KAHKf7eb0eNXSiv7+JksbY/5L1Qx9j0lh
FXCUkpO/PniFtN71batbSVuZV4KxV2wzCSVmeTUgvXoUnA0Gg6w4zGwgzbeUo/0d
gN2dcKdHxc6e85dhoXv9sSAS6wcrXfShbaEdzwIb5hQMj6IEpjdOqn2L0eLzZ8Ix
L3BGU5ZgP8wOq8Sy1v8ASd4LIVbWFG9V5MTS51CksW1Ks0HsCzpZn1KMRl0qT9n0
yz3OzPU0q+5O5px5a0q7qjwHgKORwHwkYEVpDGR5Tg/ZiZJ1PkWh15jMrYmEbtp0
yCIaRFFUCVk573H2aV3gDLwpixSamG4I3b9MdfDWc3Sp3wmxC2G3azDqax27FnXn
rHtQoKGf5+YOYSVoUSgpP3TO4GHJzsvuoGxIyOTThkuEG6+gg0sZeyn7MUDXY8jw
d0Oc4wtyIBAa0m/0GC4nqq7Cy0IMsMYfqdM5HqDOClMKjuJsLh4fnOzCu0elkWXk
sj2al/BgmXdkRo4fK0lArLaZR7oO2Kj6zg3QMx7zgzYCC7MoNUc3v1DVjRoLw+gr
K9H+MtD52s6NQvKQY+POmZ/AUzFq3G0TGenSwzm+m+1pK4VgNHBl8Cha7mykMjr6
/ZCnQaYVUWHFK/KpsL+jt/ZtI8E7yAb8iF3wN+5pIVyCOLCPV9L3N69Y9mBVI+IK
GGP0ZJbGTBetzfGb1N/neYtxLd/lCQvmLhe9i1+Yk9DR2uBWGoSoIRyrxtQlmVyh
MNF0UABidGQVErBs8GsOVqcspFOXlgFc+NmyWEVAthGeGhfrFtuZ9ixvC6AD1rOr
Z1BrUUvQlw2CYnOTPeNqY26r8SBdR6AgdbDjic16Sk0rZBqnAB1rSg3K8J8Mags5
+PLvJePAgbFbVZwwYjeXw5MWzqk0mji4t3D5KnW8UyYlOGPkAV+QhE0cu3VlOfRe
L6MtAshn/Pnhz/VOKwtDMzjwxozbrNoC1wSHwvrtHKsc2h+A8jmPiU0XJgVCNoJS
n9fd17M4lVyZDCe1nOCb0K6aBJg1JViXRCE8UBqbS21EzVg0ilu7jGr/y6TFu8EG
Co6obExwf2i58cA5AlZN5GShrt7Vtf1WoRU3KmzurgYfS+N5g7ywXPZCSsFf8HkP
CAEGS/ekRlhPRvBbO9pcO09EPdumq3lDizY0QL8aFqaXNjVSGt2IwaF9PqzxW94Q
kgcWQNqtJK4SYhm3eAKToqAf55mFLf/pQRx2Mj1XTyHsUcZ0PoP7HrZhi4DyXkCR
BPb+oD/c7VTATL22LOVoAWXzFq7oBkC5FO6f8PEHsQhQAEuu7o0jGzk1UOYNEWzo
PevJunGPUwkjv7ILWCsLCWwiYXyQxOhk38APwOSZwEcypzBVzQU2gBzdN//JWa39
gfPLO+2lo5bBPiTMrgA++5FipIsjBEazWm/byMg2d2rcc7qK6Livhaz5TtVHpCYQ
CAWAEcUwrsVDiKqzeRcWRPZ8iS03TZ5Vz2IK9JUpoWtxQuRswih992J4NGGoLbuN
1m280q89VhKnchbmOpJ2yFXyJJ1eqVP39bvxiSuFbnfYDFqwjfJflcsTJzP71EWA
xibYYO6MP2+h73SHJNv6UkKExv5BJ9rWoEj1l+pVjYOGq1pTuV2P03FwgcdBsYue
PXvwmgNXL1q6HbsbLKqDXExO/iM9IoIHTm3bNIFFNy7417w9kdhe5dwXqJa8RIkg
nhrTIO1PRnNR6HV5W278OJQyUtx1LZhBsrorE7AQjvce0o/c/GaBtamu/08L0A99
GWU+UcwpNEHq60tiKR/QlhEEE1Nd8JRnipId3OyD9If9X6PQAqGXtwtIKo5vRHYO
vPpeYlY6nJvK/+CbIpZb5EVTBzzFh6WNjw9WAXHlURNrMSy/gBdqLNNnvGdGUczA
avlgHD/SRyKvI6zlD2LlnxuDt69yp+kYvKZ85vM0sz6OkFVi/WSgRFUVbFrhRsw3
0A57iXYBMKvPPKiYi/WtTE/AxOS2+At6hk0ILkwk42Vi/1Zd/wMFFpZS2PixIy06
zM8z+8ukhbjRHO9iptTLXORhPOVasLqmkSXe7FLi+vV7oQFOWpNAVtK34DQf0Xo5
bI0VmNpph4PClZmoXG9r/AISdY82a9tR38nWPTeD0aWsa2SaAwbCZawJofEQ3YPg
j7CfDWtIsJrD53J5aQNWPDgqYDZpV/BlLunh2mzUVeCgFenCENilOQujV5HdmfNN
YAD/KkM3ta/lGerUB3eIhBjL8yfjMVVAdGoKfMrrana81mgDjEhcMAw861gsB/Y/
HreR2ATH85b2OFc44F0R+6PhW6ihH68i7GSwqdPwhLekDsv0vm1wVxRTVpcFBqUJ
+3gTSH76khSuHqMCBCeXAizwNlE6ean34f5VizKGSIXPgV9IFih+o6OSsW1Zw8h6
Q4KmJrMQjjoM7nzoxguvo9IXs+KICjRtkWXaooykHhJhtA6Uo/SYHLDi8Lbu5VtR
OtU9F3hMZrkxJRAD21apoY1S9GrMeUeEX2o9TGH+cCblRvXQfc+gc7CFawitTvMW
+UlOhv/k034cqe8mc+oeOUa2eSKrvRYKlRr1Sq2CKYFP6D08dEoCjs7ngXrr5X7N
7EarOI0qdqvaypjcVebe5Q+5qtjQ2SK7KR322w2mbw0w/OCELgHfuRpWYlZJ1T+8
IxZTFTkUVzcNrl4Rhwnr1GtJ8tVR6Cn2U2Vr7qgnj28kC53VzBSYcasDtH36AxTg
4FqX+jXiz/3WXcA97bNDkd0JAv1ZJw0pKU+YiTYFp4wGyAlAGnFcQpyIUBsyIELV
FfF0awJwGhO7XjFQKfp1AAxdCeCE/eMsac9ZZZEJN6y6PsUxm5cZx3UYj8X9SuiT
yRqJwT8iAKoVHoqKk7FnA1JNiRoDcz3JbK2LS9gUqJap7mUPyUBVrcySvU0UGB2J
fKo4pYPd54gb1EGSatlrVZl2zhdJeyOITiTQvRJ626v7OR31f/Ns6YBZXLuFHVDf
n4XfZIZiQpUPN17aoWNRobGS85MnqDOWlJmtY0PR2OW3UR3MD3UEYcpwr3mHIBl6
6mAqxM88rUP2N3SW+LaNc4eI33sl8bYfsmxIoi4H/+StowoTMASK47s9Sg/t2uTx
MjWqbrghcWbNYd1bkuGy46KyUBQRJIUF1+1WswsTHmzfQAl+yXmNjj20jP/Xyv8h
3/gTZlozoJ5jlQMC9dcst7tXEGM0yvW2vmEMiy3ZPJ0W92CeidpiwffAHiVFfuWH
g/OMmxxWp6vrr+Mx7HXhTCz7k9zrOPVsz8h0w44H5UKnX+DA29tiMeHAZFE9x322
orIyV9ngEXa+llU7e/rcSJ7JBR+Vz6HlWR9D6nxNvGecNk5QSTchYBtJythl+a+W
XCkCzhpd+GCegNLnbfyG82mk7Dklq+llMmfGFS5PhuXPMT8rWz2iHDJiwvNyEy9O
BmY18jzIJJgOyNDRvVIU4JsFSO/2hTQHe4TggGo2n2FFKwppju9Yf2K935GPFhNu
lF9BL4GwOpeGTtCwNEPU19gbLasZzHseQWYeXqeS7ctOFDZ/Vv/qLGUk/wyJhGtY
c/4vubb0vHK6/NxYKHH16CeWEGEHo1M/tG2aXIehMebQ5fbT1adTaYZK7KDquJdy
MsnONdyIEyCeoPB8m7o5lpDYjJtjnvSOHMZ/NTYvRLLUreE7fuZpryR+Gvz7MIbG
UsLEjIz4sXUIQy0+AZ0uIg264RLTXZQ8Pi66i0c8FVtfFjAlMlW1yDOMwXoZckfR
QgE1+bfDl9gftU7SzrO8UM9A4lcWzgzChkvCgynvtlvHGt/q49ttlRYQ6kyPQKay
gJ1orcLOTyFDFttxps4mer3ldJ0KbXhVXF7AHMeECRCgj0gQyCDzNDo14jURUj/R
HHD6Ddlkd6DsPy70Vvxj7mz4bgQ7LM7lJ1kZSaPPUjrtzhZNQHV2U1vEgLklPuOk
xE4t5vjN8Qppq05IAjnE9VToxq9wuqP0YzOG05gtJFGITZO1+ONs7yxIruUMMtXa
dQN0VHrDPExXMFxhgvwxHP0CkOrtEiL0g30vmrtZlNZ7U2QAnkE/5OxT8pZvR0M0
GeSbFwNJtxLQ0TO8XSGvc7OEWIrPnEc9ywGS8IxN7TaWOMRm9dU3YXfIiHJaeg+1
LqchaW9CQ8UdVpCKd0bOgr6mK9QdvClbtgdCITMbajYIp2T8p8B//LlmL6IZBTPR
DEarrTgEmxzd/PlQCxCQ6uuezQU5vBqd82TDWBbDfAac4LnQ7q1oKkp/KypZzSYh
xeR6cfxDDnGHnIkjVSjicdOAUrC+/Hx3LovQm+KsZ3SaZquF9CjYnrM65ynFrnVs
z1vl+m0jaNVuxlMG8RFIlXZxk7pF3XlVqf+J51NuCI9JylUAsSLAEJC8Zn6gZfet
xtlC3bUayjxXK3A5RvP1nk4X0SBkpSSFUV+wXrxOAw71VvHAPh+e+A8rQ7/0pcY/
QqTjPBoMVGYEfLRx4jBzqu+l7b7AzBx7Q0nPXkjOp5qrDd/hPsWHi9Td9LYusTeB
RkI+wAQJPXl7MtEVD6jehv12TYthU4Ns94CeYe+s57354VTksPGUY+iXIwA0Hpe/
5AqL1egidobVW6hXhlen5IslT0PtxYAMjqV9t0w3zgIvX1wGz6lg7qEqMNZZf/cP
/kKWej8J8zg7L8HFVgKBRcuUBt1buWndsTcLKZKzRyL3XrhW0nNEBnraENvKLioh
K6jg4RgU19ndgjGcCXK7PnLnLnXwzijuL9OcHX8Zv+KzJJqRcFDSZHV0u23m7Z2l
8ID90S/tkts29uW7rG3KQ+kR6SBH12p1plPmGK7dmpTabFGQL9iml3rWz9UPQHL1
X3dvK6OGhZnljQTc9knMPG2wSzHsrADkw5HU+WCjz6Mj1XaA8NcNyefr0yPOwJvy
wV2B1RYywxLjurZUlVEhsc8+S0oCd5y6a0RZM/mM2E7okwwptweHdFmAMrABEcAz
Oh4x7Om4a8o1SRrYZAxG5q0xY8Ugttrn4UGbDkUzYunTewM2L1Akyb8qMQs0fTs4
SOaN3jXoIUTsUpH2yJIcMzZM7g9EsodUfkO3AsiPiRZ0y83bfPcPdOY0KonkuxSg
Vj0VlimM+V/7YjORqVGK490OiWKcq8XyZtd9L3MAsUsMBoEqThxRdy541iwNDlYi
RMWiem2oQIv+raUurt537i78qOjrKz9LaH3ZRtELn7R20Pm9CcJz+ct54mpZYnB0
fNft4Zb7ohkR0FZQ5nHghIurFFtJCt/71iS9BwCi3wl3tpzSMRafxxW2rRjRk6Ul
TvBh/qlWLP69wQwM7sNnv8VkHykgG5wotDU99dmx2KmrPCLtM7hK0/UVknLGb9KJ
xJ54Fz1GMs2imdOzJ1eFHmpiNADjiVATENxihXLABIx5lYe1vtmFYEm83zZvlfjH
UYXy6GDG1phYnoaHnLehK88WcJTXVKFypyqE9UdV8DmCi0gfkp4ofPZf5VXxQCIp
yjC1LPUnOzVxxug+4SDuUJm4uAXxDYNBPE3yySGce15q6lV/f2PGIh+kFNlYv61V
/bCdoTRxDIHBpd5xG2T8deyYTV4qAdAuIUjAPxiVgYHRlMqy+8Fr0u/Xc/5FC7YE
Ul9PS7fsdIShkW6GDaOhqDSoQ4N/lLEaPTMoZseVqspk6Y4GgcCTIrGtcCDP/3Ef
VoS/oL644J5UrkU4bY0UZnMXNjUJ5nqA/civN+luc7jL0K2q1DJylwFd4xyrJRxh
BgeFru47wgoMslIkVV4t704mCPnbZ+tNysNiAThBTng70M4ToXfpXJm7kpDiB528
Wntahr79UaeroEwsdjn1nnK/vrYc6Q4CwXyxFZloR1C4oAmsTCo2feN6mHUK1hxs
cGdRbbs4UqV2AbAFu3GyBY5usGgwCf5Q8qkVBN9sxd4ZL1+t3IlFB3G30bFyiWIt
zJMdZDQnIgyfy0AfdvJv/drfr7AUS4Xur3lEgR4a0mj63JACTAekCHV2OjWYGiu0
d/XSu6RS7DJjp9TACQ+ZC8qQqDVg3U3EOo5fRBRsE/SR3yI+BeCybvsLNvPYloIn
j51LyMdhReF0o8L67GIVY88A6FjDeSKkNmhiqHrLhCVbE1hEt1eCJyOoA2FANo2+
zwjWpPOvAje12ffDc5MQuFh9t3nxueHKWCXbKvgZaElLz2rLyiWj5xzBqG+wWrIq
WWzWoqFX3HJCi2AbWIeVFqPS3oDK31CJx0+gQmBFR1qQTlbce4b8O82+o8ucYxRl
l02vt4UJBKAxst78ZamPyGZafqRekkGGDKr9AL7f+ZXugIPVTrQxyDgmxvmAp1Sm
r/PN/tn1taSJjKV2dg5NKOQKS/ajPYKSQaMkkdMiPaFMfYTDDcHr7eKWo2Pd8g/v
i7HtJMZ9C9eSi7IW2dyn7Uq9xWx+EdNaPbvflBw2TZM96fL//ry6ihlyG2+y/1ee
H9DFDHtlITQH8G4tAMsQ80ChOfpO3/vdnK8/UU7OIQ8lIVyUH3gE3oHLNmNflMgS
cPgMExbE192p+L2oGbyH2Tc7kKvjqnd8MC7ZzuwdEQK4tEbKUY+UFf/SEkHOGPok
WrSiv9Dkf1Q2BmCBep2Fbp2w+3P5ApmWpvdb54JnRrdyfuSID/IDAeVxgD3pMQlj
wJ5JoCw8VLzYyMeqRYm8GD7zdwh+w+IVsfmfuKmpRHiUfvPiUhCAHIA8v8M8+mJk
MRZS/eiNTbPTCjLqmFnWsyT9MPZgLpwEkmfhWfBqpzk7NJH24fLgfxRpSYvWeQBB
tpIDvBIX0qobt/ss9sJ6duYCvhs/5NCmfPk6JE7viILVC2JRGxGvMDT/Sb64E5Ww
luknUlSKAYldz71372Tysy0huTF8CCPAZV8fTJLuHWC2aDRaWzqflK7fOzQTywzy
tddKi3/Ly+OppqYenKgcW804NouyrQH0r4zcWs27POmRhHh8DyaGojzC8gDK113B
NUiTmesZZAaneALbW3z0BnSzGXGQMS+Pvo1bsCWh98DkdNEQQk4y8rz9CnktT8I4
7MTojDgJtoUhe/FD3ZRrAlok/Ivam2Q5juYP7xc7GsxG8PER6OWLbamRTETIEd2e
9ID7Re0ELBZIAwk3xG29dBptYcQkSDSYT3Sx01qbL0sCpp0e2NFzfQCh1G+Pr80N
UYh2DM0RrllcpPK+pYtrBl2WpugLeEb3/PFyYHFzqIOGF6INPmLn2IAZBByAu734
+QzrF2NwytcFR80IDJ3yD5dtxA2177GG43uEjdtb8cke0qGocrjpNgJp7d9CVR/+
O/bug0k4+pqOCgWk1+KYCrqUCa7wUcKoJTrAiVVc9r/gngLqiIILSm0o+KYdVVhk
e7p2Nazl46Cn57smAXngoJfpqWYEvoWs3db4bDWeYHMPCQXaRvJAjHe0+d8eqVTP
LF6sheDRHaXMk+pmlznN5mdvW5GcVe7i8/s5khkHPC4DG+iZ+HQBp85iBVkfh1+f
MbtaKHpgXZi1Wn5muz5L+qv8reLBbyEMYeb8VBbEs99YKag62niTBtUgwaP17iTz
Uo+i4kOCb6htfIYQiyJQ8SyHxDDr6pFBJPVAZi+JPi4ryJSKPksh2SN2R1nUBtFX
rPA2QEqXY8b57Cf7NqIDUyfCH+gJue9/AjcrCynPivLs4GUHnyyUF8aIWx3BkHY0
hBFWCYMblwHM+tDWIFQcZX5bEUM2fNxSUDoGxYIqjfiV0tB3jT9qlgy9h6UILahk
z2GwETJEwEsJbwwhLBiDWD7pN6vZEpissegyW8J3zQbkBpKkUUV0mn5URUUzmofk
i9Grjv1JqkOjg0bbMO9ACXuSjP2D69Qa0jVx3qZgyhW+xbPoawzX+5tCu/kPoyHD
O5WM5j5LhWh6yrnc+khonbErJBdgu5qR7k6p/MwfwXFo5AtreMMNk1PGCvTVZcNp
qwMUV5kWZIn5Ie6q1qlAwnVSvfe0jxvkxHyG1UkISlvEn9ji/ZJdP1euyMiM4viH
YwDPx+qkjwTzCE32AJHLWFF9SPQE/CrggclqB2QhiMiAFtBFhguYeWwdHImL9lad
eTNRp75K5Fo6ywOYla5gDXi66eFu5vd1kE1/snInm9JqeevKhNHrQsfccXTPAU07
+LTb14n2A+kS4yjP1eeiWxPut+BOUX79oeSpSgOOY9PxVDJEeWNGpqF0E+giFieG
K2hl7kovWSyajDaE9ARxkYlGt5LV07oXCeYUaJeWFMeyCw8y4oMZLSG/QCzjGDTZ
dWl8cx4iJJdTs0Lj4+Ai9K6HbUxKjNgvn49QzVfK9wdRC77xx0nbsmFlGZ+n03Xk
UC8JQmAdIDeoL3fmzLAUjduK/smInfftTTviTO4E9orC8kFhrgrk9Y4AonqSrAGc
t4aFgov+ufVzyWkJscZp3V2dcvd+5H3F84mehPIU62xrwbNnRCnacKG8rNq58w8s
pFhJ7m+3qeWh9CN856Kd/eb/IoNSM0fiFoAVyHgU0TislnJ5/o+AWSuly131qzLO
uK4tcO3r+g4X3SRNNaf6j96SVSdHTV6ZlfhqhworCeCU0wZK7Sv1qUof9RQHIALj
m9kzOr0J4s9qJE4UGIvem7T820KMUD+NIhFkRuOKTqzcT6ChSRKJymf5xrYnVcrx
o6MCDDSiwXUbP2u6IfQ06qneSzJyjEcUz6zueqFV1dWCdXK2dJal2oXC46VjMUaY
MrzY54siE9lk1GVdrms0o2A/lCh2UPbqDwM9HEZyJfmcw1qKU/x5U9/M60l0FpYF
3YUitgD+EYLR4S0tPbgHMWe+VeDplghvkHezyKiDIgedVg/xQDnRxuycZR2D6Q2p
9L7eiGXQFP+uPPBNlfDKo77bOaI9Js5F53cDkXDtWe99eyMKKVSqxHDijEuWHt0e
xTweo0RUnaZDN1nm2OTATdOPuHSr5RvZ8QEKX/GF6SEVisqfHAKonamD4f0ClU/q
O9JkSYYQ8WYzHWHgbZQ7AOdQZSF7+QX4kZtLrFyCXfn5ODd7je93MBq38Z4zPaJ0
IsN2hax9sN0T0C1gsY9GtnhcckK+y4eySDqU82ZZjGmblOu3PgrSTZh0GWrPPEgN
Ae7iBBOxliBo0ON7v0+zTryJI+qjLlgzdZb42RvvThvtQzXYGL2XyN8fs3WDHdm/
4I0gI8z0T7xDakVnrisIWCGbZX3YtNaKjz64CrsSd3ZGsQ8lA+UQVoZ7JZQSWFYs
T5+VoyjEkAOFhGwtqrP0K8Co+KBWBSzgiRXnWbnMxUSA4K6m12BhXtWi708+k1o5
vUE6NzOp6rhzh6ljLEqijUkHsx+ShDLKAf3UY/6sQkTLyHsC+DpCpRsM2GKL0Bnt
HR5lQCjLQqYlW4r5QX0hGuvR6LPOJUyFFcp9mvFVoidApVVJWm9MZ1pHhnuoHWW5
ax03aQ4O/RS4qB2gk2xkLx7eCX+wv7D9t8+zXh5tJQbq/quEQigsbAL5PX2HxGGQ
guB3sCmfqAvHEiniJ7OjKd4BNdnH3P3fgTwSK5MWGR5uYNFpO10ZJputEKT61ghJ
fgCwHLav0pOlwSd1Dbsq/UxCaichkSFo78KYXvgDO0HeZurKAxQ2fNMvlqrKSKDN
cljZ6RMNAVNIr60GhdIzmeVEzk1sRjVybCofTycoMy3FybCaE2pOGXZSDrdOEml5
6x4mf8JWJLlXy3Dy4ksmAcftFlcNf2qKgpZmKiv/J2AxgsVdugzXzJ2vlppLfVIf
50WnPHvayC7KcVUK6sqz+aEwyCFEpdxc8/xmKdbfuFMTGzCnpWh8wQoNRAorXI2j
5QNhQJLr6279Z4TvITPfdu8n7X/EHumyE5eiPtXLSBo296IMmcjJcErgaebc7GRw
7Ym+Jf8y2pFnYdOUHEGDePiICbz1oOKEGWjDTHaSGuo3oMNMgBgv8sYz0Rg9SIMu
7UcrGVqdYD5rJ9SkqXQQsf5Q+KVwSiNOpQDvv5X8VprFtATq9ShHf2gbwNk+ZSsu
ETzB/1TOMpChRLvc0jW/dGSgMKxEE9uoGxgU0WLfx/Lb7Uhx+JM9v5pCIMjOKdmB
czmLEHAl6738vxeVdnBS10JqjhKOSp0Jn99i78I/p9ny0js5MejUNG7qOIXXLkl1
VsXDMwSJonDqUbDx3PXHak/zVhbHK5liuz0sK2m76oKKfBs9W0I6ju7F+zXOw3m0
vNiaL5NCV6mLjY+bjP29+mzm15uzNbMdJoYQG5Fc5IDshx1RCnvoybv/gZJEWgAo
hrl6ihcPYGiTB/Aib1SqfmquBatGJ6Il5teqxihw8JMd8ZTbX23qrMaMFRhAP1cT
5BmqcePiYb2Sx1treaSKZBdtWthJDXS69T4GyBBRxH+phaSEiDdx15d96hPMEx4A
Rc8gz/FKEt3hVphX9qU4VCEUwY0COO1MSSxPl6KIoZRclWliGsU/RvnKfdHSipTQ
GsAkaS9xVpxDxfIm0fQDiu7wiZi51RO+uNgthKRstI+NHiclrst2gRodNmP/lHJH
X7ERcDjiXN722OsyNbdNtcjCqrkLZO0pti5+KoNWD2QAO5EoWuT2TyhdAkstCEuK
8U1Vod+likn9fSy6816xfqWhuSC65hxm4rwpnIYeTJUkmMU7mXUuzHyejEX9QEvg
eygvI75k7t9ubVERXYgtGb43aggR9YoonVmxGu/QrDTBB5QUwmeGWzc220kUMYfw
g+QcvIgg8MVXZYhhrvz+RrcgxuyEPx96eGknfg5SE67GZcwKs8SXU/hQHwOgSCOq
K2nlWGxyrq7kbyQehn+9fvjRMAqscTnfANQGXe7lMzeK8T0wfYXV9/q1Bx6evhzc
H3b65sGxPvuVT+jeafUYQTExDpqylXTbIbs6hKGmCwDT1T4Sp6bC3PLfD0AxNy0V
AUTfcBujJmb4EEqFrIxwFjqUV7pzC8zz3wI4zHgWkvy/Yy6fF8M4oAY/M9xOWIld
pDeT4/fsfYx4dvNaTJk21iIoIDHDZq2QqeIKsq3TT4xvH1Kh1XIiSaQR2Jk47lVD
+k6woi+uHvLEuEkuHBbA8c6i/xnVD8YA519T6QiY/Ci9aw6k8yI3tSu65zjCQBjq
7/UQ0aERW8u4kV/PgcodZCEC+HGkFjUYXhb7M+8yzU62HsUPH46JF1AMK7V1pISX
fNi9vPEbjMKqKQIFwcSoymF2G28d1AxXdRbVheM8pFaObJCJgj6wKX/3oS6xjpC4
PjyvboXnY4Wk1L5zmJkI2OtdvAnZQoDrFMiPFG/DFT1/o0A0fIv0QqtIYXjiX260
wt1dZqkxX4ibyf6ejavq7yv8S463b493DQ+DQCKlh0gQZLHZCxFC6JtNPJVDY6DH
RjeyZYHrOZheFaXowV5o7/mPypEXm/qYzDHJdXqVG4Bnj5XE3fUe+5O9tDfOOB0h
4+LFmnVcEbReY/ICd2S+t9PSZ1Ept46fRwYWcGyfCZjMHszpa9hbUgOInkBauJGW
gfqZFcoyPYzYgN87GuH3oRu4kiw7QTJhxXAjJR2NPoqagGF0uFFtNv45X7KFMaNd
ejKFBhR091viQYupX+pWqvaEfgdJO3i7iBxTutJFZP6NniFzYyeujcBuMDYXWfRA
3ge76Rvp1xZYi1qnVjj/a7r66yk5WqST9kllz3QxYATZuJJKnBjYMql+T+RxmCR5
cHjBDiPsKct3kagivs/0MCQWY8SUOo68PigESDhbw0a3wYl1uV1vsMyWtVP7ffdn
qJMg9PhUy3QmDB52kP54IEqDoJyb+0xWMEb5F8jJAuISciAEHZyLT2cza7QdEvtv
eLvis89wCfr+yK6pi5BZyWvuJp7TC+tVb9eAYMG8a+QbxQ59fu1NGNzOsgyctNBs
RXU3+VoOwbTI87vRgunv/qdI26Pixg4XsJDXj9z6MqOYf25/n3rkASMUJsJONydj
myTSeSBViX2pNRYPzu3fQOUfn7eKKBWp95mMTcIIWp25MwqJOluWwlWlZ1nmPWuW
lKFWMqOYq9VV10r/bLw3pN/cZGwFVXcwztb8IqkWIHyNdscmcyZxR4jQqO0dTZiZ
2iyudDiv6udFzTBuI2nMTNg6bwvXEWzRUF2rafw6xBgiZl57y9NxDF76qQRq4tOY
najslof4fFj/R6dvG9IzMDqiAdqx8m8Fgr/XzYBgzOVCX5s9nq8A+JBVELSygvLv
kvO2VDuTV5EzBfv9OBT1WqPDA4HzdbJow0FYOFy+RH8wzU6jc9OctSpY1cG/eGGL
xsOdppYNshjELUdu30GX5AEPdtg/NaR11fI5vU+8+7P6jyGEo92gZoN3cHfV5997
I5U58oTcz3POhQPa5QxuabPKLUGBk6aWtPPCYLfYDDOqwrrIUUg5GU6snUpn3cTk
eRDH2kQCQwaFPciHoLx5dnRWK1vxO4O8yaUkbrPebjsAU3R67PRwmcBmKC7IYxcw
2ZbywNy8Qx9kdzLu3rUVVhXQXHEPD9WPLIGIYt9nZlXrs45bvUDVTNynHxMYO3BB
S0ZL/UaBvJBrqyBEpIh8pILfHdB73nTVgqT7baUcddRzWpjs5yAazwzvXe4WDrzC
aiHsGKWRZy9ggxM0ogeDpcAWkFgIf0X1bBhD2gIJEr0dWj+lXYOfEL4OimlBi443
Ig0+w05ZZ044sYBFsfOvUB61mx7gxvs8eOvnvZnQIEE4COQC+Wtn4Hv4RH7JYeMI
ppowONQ7jPTKp3zVuLr8nZsogbUFIjTudzA47TyUDH967SNwtzzX+nBR+5eHR3vm
v3gz+sXqj+yeg+LiKgHuViKyhOh/fnXHtgjC0YtslMEVBI08cq7oebGvHLLpjRIx
J6zBNtrFkkiIBtCrcyFcm9dllp2mEnqtSIL3tgznn+Uz9xH7XOgzRWMgZ2svKg8g
E6tv8OF8yuPKFKjXUBXWWB//Fi36xQxZlt+CYRJWkDOw4iqeAcClIM/1h+svGd7g
MnsLOTvi00TfL0aMYo+cK7bd4uVy1L+4gUSc8uQcvX5YW+LbZdYeZBykoeuSz8o+
gbvBLZDfoD3y5DhyMWh3ZgtyiHfKn6rGZ8ZsJfjwE7eJAigjkg3GmhKiLy6eqV+K
OD0NVuJHi6BXT4uOEYiulalIUi1f9j7qEIrwaqGSIZDgw5pIwFKdpvblU4zxGh3P
9tcOrFh7MAzXhKOGhV9cq9UvNPsgc5CW/UQ27tnD6EJE00G9DkucHyBHy1+N86O2
3JY2Dci7IOl72MteD3tZmqwdHowJx5rCaBj0PnPXEJQGqYddOmYeJ5zK9sXw4Vq0
Dhj8eKb7U36tHIuM2gBLouT+zJVxZyZmGJdyaMWSgYMh4ttlxfiUuYKLI3pd8Clj
n9RvmQ0xFGTbW9xeQfBGi2breCe16lFnoW9ShqP8iQiUEbaGza0KuHblu8lh+JF+
DtoBFXT2i35NjLFY6C8GZNXk58IvAdSNIZhOt7DqmsaEW68+Z8OsNBHsufObMniM
VQwNu4mV8T0cX/3vN288zp3pFD9x35W+TjaTqY0BnbrvUcQrONq7/DYalUEtXaGY
Cy4cHEM0gPdXOty2qV90Z2E4TeC114E0fCvovTk6g3SVs0HvhZhOStHeKFnFwnna
pbzjO58HYKholnznIetbyu+4Cz/ejdluVBXRbTwtCkJL3WejwJkaCMxQht8Txfrv
BIxg8ixaX+t8Eb+ttn81OdVDaCCserZ9SLnbLbf1WayFV1eCiJciqg10wfkMgR3w
HHyrqTvHqwO0eByo0CVYFg2FThHm/6MlLctQeoFTTanPnrMHzUyxGys9B+GU8Oui
kt2k8MMwFev5FLuE4JnxVJur5mkDJJqVg5XBJaQrFbElwff2Yvdt3hKE7WLUKYZJ
O1YCwbxsC6nqiJFAiRU6tPriYA1ZAzdgmpl14wTxfZ3GelUbXPuPBW8whOrkp4/U
axdNBNTLyH3VLITuIw8K2iRy5fAadPNo1twMThbjuX3lMIRAh/GHlev+vjffzudr
5Pzg1lxHw/DxgYJ8LFHNHHMTF8OFrBPZbHNUMhOYXEL8S2IXTFnZYOEWnPPaYN3O
NbTwfBE4CSlX4Mth/af36StpvVveyXVuDrDkRc5CwqJ4SthryVGo92Ci6yyShlzg
Yxi3iqKBgWXSvJxNexZheABmcSehEmHxj4EntEX4ud+PQx4+RZndCWSTCjM8aumz
OOIDfZj7HiMnZSFUcQFa04eYhA3o2G5+qYmjZN7DnyFidb7RiX8vUzCIet9PT3d0
IgExZ4ladtNG1TTOLiMpYjeiZcR5IdBAOUGZYxSQ4Oj4IGI1QfDC7SCeSzeEyy61
ZHsVCxOiL7xDxpu++6EBrTsv81IZkRxAkLv/KhdouSKhRRMOp98vcJoOYYjo2r4o
WBKzZoZl/sW/SzxVtrSU//534/jxUTdxsiUkgaa5a3HCl+aMaFTNT5lxNW5qtMhh
pelfGPEqBvIWTX3rGe9jhuBuKyI+EpjL/c5HXLs+YaYbMMplKMAiZHz7tWtVGIAe
bE2Cvd+T1uPLoSDNfMY92V4CRglGKfI8IUHNhXWpRyJapeM9doi3gQVuBJuxV6UJ
vPIBHD+vHU3XqhMWNCXDwQCnlBkqgu9flq+WuHSVFOFCl6Ny/f+0bVlSSxM8GgoB
JHpNyZ9BNReeMHov49SO26Du2VlEqvuxK4BklY9LOMqqKXcBGLtv18dwEMMg6k6T
G4VjcKMzZXABQ9OezJ98hw10JMg5y+xxS3ZBnF3LRHOHesGIWkvgG17h4LV0iyUx
4R/IFYbyTL0qljjw/BqyCevoth4rUGbdc74rAobD2x/cMVICEANfmhKz1dUnP/Uz
pjnN8pUzflkI3w9sxvaU+e+T1eyKSjkqrPADKPu0tLc5Lk2LPXAh5M/4w9+4FW7P
/0/g0azbDXTqi/AUqymivBq6bp0volacUkC6JBZJG0n8Q83Y2lsILq++P8i36hVr
iwedJUgr0o9uTAbm6s79UTlyCTrq3mRH9I7csFlHfpgKLAu2gTNwakt7GvCQiE2c
Kp9oocS6ibmuSqh/6Qu1z/hRbjFMMp0mvcYApAjuAyg7HzIjsTWDlfNAxySDpsLF
7gAMgymU/bY2QSPLOW/T+PkoJG2YSALNXejgKcz9Wyu+iUR5zguG/gbI4NxUiA6O
YV9x8DwPVw1oNBvp0MOerEKxkjNxKFZPuEkm/CMBtXnFSiuahTBtYUqgsxseFIDr
SQlCtH5S37RNMdf2i/XWbdwOnpZu1A7J0R8F/ITC3fhT/wlyP78+4oLXh0OLLXCZ
lQQ+FLh1f78HpcTmsT4+2M6vAdpxlElvSCc1+v3MwIzzwCyLKbRLk1Rw7CcyfFd5
7VgBbFPxe3R4zXFcDoF7798/S+4Brpqd9wZMauTaj2ClUjYxGVNKOkwkV1H4CPD3
kSu0NGd7opo9Y9ylrFsyO9osyUbUc4qtzkPHuFPIKKMTf7uNwg0BGzQlMWMJKq59
edJZpWxvfhI1384p6IA7eVHKd08r6tsDru9xncoG9AdZ2/WJmFzCFGVaHFckDHz8
pEEV5wlc6l3MinAYmDwT5qZXt/SyCcy+S97OQZIEnbU6e8o0zafAmo8rN3bOJmFa
K7C5pss2dvnbdPfBgTLdx0leUHnJRU7Yu1JaC+pwvVL18TLBz5T6KbGK5de3yGLd
6XqtLRSp1u4mJoOQVYJrLx2j3TGYEwsTG4TC+m+3R0ZrP12Plnj9yjThuCOAai+o
mfwT/EWWn8WxlQj+gDrTw9A/k2h2ZTxqhkndMzjLFPQBlnBviQSdoxuaD4j+/Qu/
h7dy93+eV3jrQTdXChUVF9DN66Pi7s1PizFZ/ms/FqKOpUWlWVIm5+JzPtUVRMGK
cvcvgepL/PbSs7lMqNYFvBKy+vxih2B9cnjfrrexUdymbfRm7xjCjZSKswqpvD9f
LMu/vOWNKUjQ4qzgED8+7RPPxBIWsj3c/i0/L9PQJ1nkdBMiHSgkdvk9mAe/yJtC
QtZ6F9RgJD/6uinIsoyfRYELR/5Cn1bxo/9UKdpfkaRr6jUlBEnUXDgCezxFcsA5
01PKQXS+Iyqh/sTAd3qXeJyMartL2sHFQbwFfZAbRczVCZcfpgSpnjdAbg2J9iR6
Ru98OclqkGrTxyC/zYXM9tIFs9b3Jq4CEdCBsNS0uioMMAVt/2PdxzOLkXcUWwUZ
udGcmrMCge+6IIhtPAuLvS4nJaHbqW3DWP/vXs6vr6LkJ7FMY+i2b9VBQIQWu0VX
weBZaJx6t4/a/O97/kKXiPc//ORPys3GPKnIKs4ol6fmQWzPEoJ4eZDpTp5rNKVz
ghlfQNqSmCsfwTdskoKe6i4uKEcvaz6b5ctZJDQl6awH4VWJQRu34IguL6RqbsVs
gwPCzZck4NSPu3SYteOgFdoWvreHyY99eUYfE86SabD6vwO3D5VWi2QZKnDPD/Rw
xBxVqf1/nF4AKqPso2lmW8ESd8p6hfy3XquxMHiKIv1jZ8gb5Xp84xWpx5cg696l
aGHMuyDgrf3EyW7GXyvdCHhKJQNCDGN7dRpTXHjN1XEoXvvv2vLzu4p/3555Nxgc
z906TUGFPtw9jwuw5YRkOzvwjjgc8Aa84Pt4fA1Z3xrCoM7UentUb9ywQNFpaEq9
swd1yo7wQVw0HXmo/ceQCOHYHo7sVWgfGlUYjD64xMqF9H582mKwyWA+ax4h6Lfe
IxhPwlQ21FBTRuhQSROMPbEDjMNlJ+UFFJrV3Qz5fjan4EnIieuomhXMXznYgtng
Q4YOhErR/c8fY5tbb7fvuuhIv6ooBMGjtsf+qTtt4RFMRH8yB2UZ6wRQlbNm9+NJ
GFAhcug4D3LeDb+YhS9OhaINIPMwXnEFr8dBv07BGY4olPRte34ZqbQpzhREvYDH
t1QJDp4M3DxBvaTq/4OWV3qoRPcQqXWQb2B3aICjmKfrUhNmzSz1tfo9y6vEWZga
fGXnVKy0djD/MNRFzrqkF7+TpdfrVW8ztCikt1tpNtp+evfti9WEPBo2SUSppTrv
Fs2QmfYNYC4k3045LM2s67/JJROE3pj4PS/U5O/MS9iiWTQDf0GmVq9NCqWWsi/g
+mwy6QFo5w9uGi8NevEjh5PEUpuk8VaH9HD2NXZdG3b6z0Rw/PHn4dQUWWHOhUPK
tPiLcV5FCnr1r7geCj9vxssx6bn8CNn/SAgQxWubjzhdeaZuKlfaFbccKbb3Ap7c
NyvDzMNciNUEWEfuvb+MnmwevLzRRNoXRgitCQJu40EKt44Pb78DUKgJ4wfrObdw
WisbMrwNt+BlVAwnnO6VxP3Yl5UrLvF0oFyFAWf99KUl1Zxfm994ebktzdI42yy2
E+tj53EOGXNbCya8Rk0Vtw2UemLNgyVrgvUjK6p5WpxeIMmWUo8A2ojgrl3sMJCN
adBKXVi4+JZc+q5MfOkm12AwQGFgPLVcrSIGjSRMVMzgbbpsJbpEFJgdSyZDTrtZ
LVwAoGpWVUSHCeJl8+CT8rKxyf/eDqmMqlPT21nNKVq8vsIsubw5Cb4zUVgruiIj
mACYgZ3Smk8LWQpHYO6QgD+TXEdjQdAnGc06a9MBw5enRdPhcntWH0o/Iszwg67w
4zOMFb8/Pdl02Cq00XmAUbO6ifzZTuooGs1vU2eDbJPSomO2n167cpIkLdzWKtTs
4ekeBMt3TEl//4Dj1dIuH3F1u43GGXV6bAHb17kcFaNon+XrfI4T4NPioj1IUh/Y
zqLx31sUSbqIzU49WNkga10/PvIvFqCEgndhlvYfCzY91Y0CJo+5L08XiulugbCt
+BW8EGP9L2ZmzM3dlQIMDere788hXjqxREzALqoopdpJsOckhsYt7X6ObWDxy/p6
5WgKUv/OCisR+EdiXsjrypPrwiWpBtwbHXbfOcz+b2/nY7WY5gwHIB6bno6O/Fja
EanWD38zKl5QzV7AJ41Av9HGyl4tuXLDVBpXGE4kSXe9oNKTfhxK3Oa9ej9EnY2C
TWynAkcqii0ZrhU6MVDNfW3tuPUMHnnHpPQY5Hs3sPqq7csr7tXR4WdkzEsj4qpn
WHrcWQh1tF0iM3pIW7oQBtObSrTLx83NVa3byIr+9PIQFFDWegBuK0M7P/P5xwrW
aST5rStzEXAqoZmaGB3bs4Y+P7fvrc+ZFy8x7SpQSvgrSZ2sov/g7Lf/+oTSNfMq
aJaaMuVii4Y1mX7E0vIaeKH6zJjpKuuuITYaIo/7hIXtnECSk5G7oywiez+kYK6Y
7I9Gh3dAFxFHuBqrh45sHvEMArnvEf9xl4CZXqaN7a1HHBYhZm6q13HJrZvgHuFL
dTn4gkZFZKgzd4XN23YmnhSJUocn2Oo2DeghmpeF13rzlh/LtnogCJnIjLfXFB5o
MayoZ0ZkPCErQUVg95LlPt7irHuwcZZACsyxqDeqHnz2kQCCbznc4ylwqSxtcuyf
ln99YmV5nYkGm9mjYq/OwGWoBUHWDRFrUy+dEgpsEAq7XpGHz6Md7UyEp/0No/oT
xD5lSkOi0g5pX80Aeqk4/T484obmgmzdHhrOpunicho/mf0dNQ++SJN134nMe+Cj
QdQp0VwveTat96Lu2RJFgECecoveTVsP5GF78wnKtIqL4+JXRx3F/tRGypcXkZRZ
0x+PwnXc3gtt5Ux9uvcIRZMLmsQDX/W29TmJ3RZQ0sNdNs2p5FsJFp3ElSApXsVX
w8rKzG2W4cC90d+lnI0R5kslby0dkRI9UIghs6XKlYBcozhD/zRNSxsQPKjxJ+KZ
bIPBdyu152y6L0K7+PQH3rku7V9s14PbfCCSsEgjSu7+ceog7grlEyoVrvJt2Yhr
iuLz1IvkIagZ9LPjaPhL6sv9z4oNyTiQojTO30DXmggiPtIPgSlcrOfvSBxU1QqO
2cUWcrOFgbwrbFo7AcessTyBBhPWTuoLaKr4tLk3IacqxV+jpmjmblqmt0V5ZI4c
9wmMxRTezmq1vt2tGM75URgaWkpWsVRxMCRkessjYSg3yZt3Xbaz3d5yOzHpjs6G
/kTESRhF9ws03lfbywVi6edHvui4+GzmTaJj53kaEWHT/cDTdt3F5CAwbLK+1srI
qsLk+zVdFg8WDx2APVa5SDlJoSkBSCCYE4ZNPuJ8QhkeC+cR1Z8kOMyWGZLjIF7y
lZ9tRN4kzGc4ytHGlglu37SCVtOe8B5iHPtKrY1pJTWHJluWzyNRW06wS9IQNRVw
Lm0SiwINkpRhx7MfnApEEcNca/s6MehLtZPzSbddn9dHAuhEEmY2Kj42sbXw5gGE
yPFMxGbdBrPeoyatXKl6BsGiBL30AGcjshg9UF3O/PlMu5+S6DYcMZs2ElPDTSoS
zVnX4MrXg0A45Oysftw1EAYlxFv0w1DuLTFq4+4dm6Cszhs0WJrVZBAMf9bbSSVH
V1DG8m4P0OqAoafFeYEiKSXT1W6TTEzSQ54iuJYxUhhEzpjk2UyCRN8PsWy/QkGD
cafgghj3BSCNWllyanNqz/J7NjdG4HkzyYfliWdcr3XdQQlSYdk6aoHYgSCoi4Ec
ao76Ozc+fVmy4eFi46v85TwaWue1MCJuQrODoKf7sFrt0Vi2Rl3EWBOvvs6t77YZ
3gwCO3D9XDNiLe/f+En8Ao0fOnnDZ9BrGKHYLtLb/5WRJ6s1/vMfO5dsRTtuheTQ
9XY08Jx7Ii99Qo6VboAcyTVRp+1o4vj7Ge/LH4e8HgA24nzt9r6TGwU8GFwwng0r
me34chMgUzPJhzQQHUDgRTPwwcynI0vaGHfflYoKy9mVMoh8tq2zK/7JiNCCKUG9
TWwxU70ozKUplkvMJXsQDxWTWWv5nhuVAkM03m21r6HuLUV1PWQmAhZ28rqiWPQt
AWpRBwstPSYDRj2Q3YAoTzNzyqvTIzlgk4SwOvTe81fZYxPy9KDf2Da7jvl4HVzZ
9C/BKq43tHzHvZdRE12958h7Rsuq+HTqkw0ZCmbyQFtlZC63qAQJ0UO1VZgeK3Cq
C7mfnFswJ6Y7YphkwWnEsW37dfEhv3SXmq6c9YJbBJbQy6bumYQh9cgztGj1LoqR
JD2Bs+Bf1baMLyDWQ2QkNncPzzAVMux2GDiQCCxygdpofc/DVz1TNmLaTY232oN1
lebC/xH6MPUXeM/zUlJzhjgrOtIerQCEvTu6e1YLwgxYwYfBAIZBRTK6bMCgMQ6U
7Ic35WNE8sAXqL71ULyRq7fmttP1m5BGLCnsyaeuoMOyOFu7DP/NhULfKaek9qm3
K7FdmiSO9U5/CMw5infNg42EoiL1kAzPIyNrVpJ6+fUDP25zdECl0obY+915tCPt
HUWY2PO2OAoN8sx8KpLNCohyKplsHg9boiV1csk5lhnlYFE3FM94piTSIcdk9/2e
QnnlL2SkW1Q7y832YkjckndWvrGSVuzuG8uEtHrqvniraVXJmeBxaEt1kWZg45Nc
X5qUusUmNv2jcDrjrMRGSwcq1VNYYdiLsq3Hhp2nk50mjJmo28e41GGW6p9qlCyA
yFfBqZ2gWCIxLHGXgUCs5J8N9qAGssMn7Tq2O3/rh6F1PHZY8VntPf+5dzd8oUd6
1MiDVATz3tsGvWvG9ZHnJwwYFj4Z1ucBnXCedgNa/qevQE/bzTJUdhKtAMDioyyI
SNgUpEFr7cKm0RHx9e9WcRRXHd7JRKzrK+4cVxLIWwibGT74dGGT3ixQMKrASE1G
JxuwNai5j90XFE/+9R9QlG5J0PP4Z2CScV0vlEE5qxWJSd9nN29kGU9Ks2r5szaD
iAXM281HBlTOPdo/CzPyVnLtLGJY9MQ7nMerptmHROy4w44QJJYSlMQW93JkeHoW
tSKrbD3l1gDPIiDDeBRfFP0dS9OSjJEi4ZqLR46yzNygHK4mrs8V7RsuStEqq1eZ
6yMqKJ1L+Iw5U91E08a1DNzU6uBxzDAGXSA1De6Dgb2J9McHo15YN3P2auY1PEEN
ll7OX9FtdrtHGUj6T6pqC8G0NTlRj6gzpZumUSAcD6I4Dmv12XKBxG25RuttIgTS
rr+CokMa2uK1eM2PXvjk8jfXgVbFkyLeoxlY57X5pYatuQ6pW/DoYyKE+Ya+qeN0
ZRK+kkuAPv85K4xc0VQMcCs34u79mqqAbdSRZWF1rqur0zh+HAcxMbEA84gl0FPq
mf1R99I+qyJ5UbyLmP+ucHX55I8rLnlyXR21fhOe9N38Wc22K3fkhTAhJnqplQ9I
iMnGes9G61j+OrTX3o2ru3GvUTyV7SWWV63lGDpvJT/2f9PaYHChdjnOb1sAH9AX
nXEup6kVYHWiAYThTZJubI0xmK8WE/aMLwjil9/33KqA6gxr+GlHHKdhHWwwVYbF
GUxqcHv7UOP2mt8FYKa2ldJLLLgOEMtwdUsdQAV0jUx6KDOzqu3sNmrkcXc1rO/u
VuVZt9Xk3e1bB0TouyFfZqmmbCY/z1v+fJW36BtXaV7u04EaXRA7Xu3QOSJs6Q3Y
FWFQzFmdAEt39VXKEQTEewGhMPqy1EhlKPkPP5UHlEze1wgim3DQBRDlJzN3RwD/
DhUsJX1R4oDIM5gj7CC+nRYKsUPoE+d+WHhRVxpe7tITHfzYI48/fL6RewXBJhG5
6pmvh0RXnHN6w4Nb5MRixWIkBPSKuVZNU5c7aj2gO7T2En4b0m2jrU/L4YNblEu8
lVgeHqcYSJb6ya9/yj+tBvUT4/l/BYv7GvL5ksHmQcgjGCeNdaeniRn0U6m4rXVt
FFf+NBLJTOHAHjwdZ9djcMQ8K8ss4j4RDPS4g2YyvMUxvvd5QYiFhr2KHF5n4Cbc
RFJ4DBURJ2bYWn5iV5EmALdNe/43+s1Iz6XJrKdNntmDrgk+YQOt6moRVCmuWo9I
bYDkqgFWA0s6dahe++op9xY/pitS+jenN99Bn8UI2DPGetGhcRdRB7dC8814YSX5
G4guDSqMBIa4udf+/xDdxFlsdXMDUM3TIrRU8upQgY8rbX0VlielnbApoSidANwt
E01PO9DoXBbJFnbYoxOiKxbNhKXTF9WpayTlrt9NVauDYHHXnpCm861MlCI02YMr
N2djovk9CfIgEtdgzv3QLroXgz8BskKurlO/t2m+l+mWSTEu09Mmma99xZ+cZNSS
8Z4tSAugtIh9MnM+nW8fBAwR/cCgalJxt/XXFDuilowDc97hCBczzr+bfkKlXIIZ
/CWmDOPu2A4ZhVq0oV0OiSOBuqrYLxW3MvOvF+GWZ9u82UkfSldk1C7eyGFyEWMs
xOzyBQVbuUNJJ3KMYN9uA9u9NYj8hMFHhs3I5s5F4Kq34i1FdSAyeiF0n0kb1c/v
kx20r0/pKpfynxQrXiNyacTumMGEiSAXKgtAQMbwc6kF0Bux7TtAmnywfz2eELMB
Y7+tv1xU/lXhEchP7xOtuCKwji3h6mHjFM1kF7837F6uBB/xlnBJEBkWyJpbnCoj
IQP7V9/M95Hb6nojl/vn99AAr8G3/DfTHAtHk+lC7wxeleclDnRRtC0VOixUwNEX
Lu4Gnu46IdmEwJjJkQyOrSi/QeMSOG+jet3s6WK2ji4N6qyLm7lM/zqAh80KuSYH
cLHSxHL0o7vVIT33dA8qlYQJ1D1KfpQqjjgZisWXpgoWnVzoCZbL6WvFVSPgcFVV
mY6eZFndIX1TUlouW5mLCkaeqv1ci1qZ9nHH6E+lKFYMALDY2wj1jl5N6J2VO4/L
4zWz/HS8kamCJH2uQmFLgSb//qXUlJYjisOsDt9WkZ9VwTHger0v4IU+d1u4Bzix
dg6AL8q0N2VuPWqRANL3avE6tS6QO+Gg0bmziCFdLc6YrdJ4LgpSuC14gvhiVVXJ
wRrMZ+6R1L91P71XjhPIOOObikTxgzgVCteGdQvUaahI1bnzKcMos5XneJIEuUD8
alcDqcSwMyGvIvBuWfcke1aNsl1XBi1Y2PQXmHIRQYzFNy1s5WqGcEgq0EvabWXY
RiZeDYiraStXAC7mC8WSk25TTJD8RAxKVBYKtFEABacbBxbOICEIL/jm1qHsnwCK
sVDSDqCSVFr5o2KFaBJrZElvilPiP6sMy+8SeRLsD0bVJ3xDJe7t1VEBhvmfvDyT
Uec1SbQiXuT14ibIYj8UQA/JVCnxQDqTCd+Lume+/WV6K893lhZihucGYIxXLnIz
b/7A9t/ug/4+3iI9QL83lBxfPT7bcR08r2fVAUWcWcVZ2Nx+0RVE1ew9kjelO9/R
98p5ez3GSBLDrrs7D0nzWTk1RbD0GdYwWy7nKZCpT1UZOpHbTLLsRi+qlDEK0HDE
iXemaO9tdtynYBA4ZIfgrjRJ0zbWuN1AOlu3dSTHNGjClHkSJZVj9y5zoL8QuIFs
9CJpuXtTKpHYTQX17/L2cMTEj5Zmve2JriD4nGy2cJno0po9AlxcPbBTkBgAWXWI
P4/34d+/ySa87tY1MXAd4QvKHsb+kanPvfUhC9jweaoV94HDZ7yXdGmAReAufYuP
11/q0O+Z4FofRsqJ2GQ8Q1M+AH7mNcV4l+wqvUyCHSm9OJClo8ennn5j2JWc8IUT
Bs7Ko8NVVYyp45JpoO5UexkfaZ/lfSK98/POtSP6lZNvqmupiUx4CLK11ZH/G3Z3
G/3+QL1rA2BFJE1X/VFr3aeXsimY3Ps/fr+H6qw6b6OxcvSHHT9nHYtaJCFSD4lK
XC1SlY1PB15mMa8qA9KY4ZqGtLUFXPxsJo2JapYZcgRODz6/cOo6RkYIICkhD43g
LhR/b2H9foDyZd7ZwDd9Yr/pjpBPJSSiywihcFdhSqh3IJp4dBGqj6v1JLxkzUgM
PyYBUZSY7kF4xCThSNg001WYyhRc54ykS5JXURgiPYVrBj+M208OuaL/DHCW/Fol
eAAi+La0p3/QyoSw2cS1W/obR2DWK49v5c9b8Z1FAcPdLKz1S2zg665diPVt4jvE
XxKijrSs0qlYwpflWQ1aRUNQcFYs549KzczqFFAefkmmueu8O9mpmj9TG8rVoOQT
aoJuuWEdl+wi8m4Hh5MNTBKg5QdMax8Snu8ufLFso4LQla/YNGGqh0FxUxsYmfNq
UieX4OhihBdVjoMcP1rn3KI7g6IObwhKwSDVMYDKADLgq1oLWCxQBXWbgoQTMuKW
3Dbsq+mg8GbCyef7ooOfbpF1fejX/1PS3ng4P/YzZVHOj8xhHkL1yDxaV+6B2wpM
DwtYrm/ryaovxwDcgpYobRJl8v0qmn2y6aKm9B2W+QXhF6DX8jLu6NYP4NopYVl2
L3k5alftyzbZ4SUNmKYYgu/tQ3u5nnv97kdGE8KX7qPz8T8W9sT/I0iSCIGeQL9J
ZmenayWQpAl2eCGya2hNikV1LP4MOVd+jWK/jk3WGsmTpZUEF4/hs4bZAMgeLfZv
5jFWtl6CPyUdK5042rRV1Gw7q5wmbIDMdf1qyadlJ6h7NwApjIYSD1e+JCnlJ46u
wlXSRoHI1XvEFA9NlWbQ6smBOsa5m6a1PgJIdn+eDEfDBXrPusgtX2NFVGg5BBjG
hs1pcMRDuVnSh1vrjnGDaCrWmUIbS7nz2OF43F4GHj81fsWtoiAoZi/s9l1ciGnv
86hH1ZtoH0fCobNPcIBKaCuUNitoU6vUfqlClw+eA9I5f89FLPuzaNoXJalRUXdr
BLY2gXG8tzUsJH1NHi9e39qXS+LBLGzyJPtuqdiSULCX32HsZHV8nNJ6T3/eCBOc
SXTd0iUDpOtJd5IwkFQ7bMuOlWP6jwF48V/DPMi32gcwr9jsjKISPjefDl3xeEkK
XcG4QM4tIX0rbvZrLobm7HgcEC+2ZUcWVfQHfSPSnBn5LVHh1uGMf5X50Yi1Qa1m
sbDidT4s1lpnc14A0sQkfYwHYgj+LRPb8ifBGt2kxrV1H8plAX7gDYNuZyx1ELnm
zga3YZN+bmUpHJDoDsNVphNPTeaLZ5e8br/pM6E9Sxep/PR7Uwr03FlQIXalznfp
VQcCj+UToEvZV1pBjDIgA7jhJQ+UsuJOBcrVyqXX+2th+ypKi0pSJ3WOJ0Khfqnk
iX4mE2+qWoK1L+2T+0FAm1h/9+C28fCKqk9YmpCQG8k1kYpwe5PWKFqm1REFu2nU
lY3tRj+qPoze5upxdNXl2NVUozDCJz9XFzygcyTeXS+F4bG9MRFVt3u82etfteCu
hZJ0iBcif4cobZ71gapNfLv4ZskOkfUCtlPDN06lr+eyb+s8pr72GPFJPFmPovSc
WH6c8KiwvDQVtt8iFYUS2XVkwtY+6mYBa8gcjc/DQ4H147A3uyq06PWbiH8GIPYa
yd+01NyS/RnJ2gPL7ZOjWX3HZxXvIscgbQWHt5ZfUVlkQiZnyXomFrClbHIIcbqc
WGevbkiwcF0SA00Z1yPcsmgZa1+sQ9GlqlS8rKPZ4pkNStaKP1DyVW9yxnxExq0n
q1Im7Uv2fVUP3BSVQbkOcSyDoyFm48CU2y7khSeQsCn1VpD7RWxTvFGikqRAlCUh
KKB2F24n+1+HANXvMR26IHuF/HpNIhterFsumB3ycdeanMEaGg4yv4eLg+UmlntU
9b81NHjk/9LwX6ssv6a2wewbW0XmZ1XLlHYhwvSh2jMxYho08CxpMmwLzFSBwQ9Y
0r2rhyVGIXF7rm7dSt8bQKJkhwmkacM1OU7lmK38A8obgR0qXxUxcf+uaKqlCXpT
UfRuDmnaLouKF+0VM8lO5CAdipqowrPe5d1ZGsA3l+kXEI+ScmGuT7rZkt9Y4wyR
FIBKti3LojDzwziTt4rOOEBakp+A6N+vsj2kZHKhPRFVRmeW79G1IC59jX56voIM
xtvYAdmT112o6MxJt65QtTkrolkQ60GRVkqq1IeBlN8ifBEilH87p9xAcIY93M5w
euk9uFdvdXH+9FFgLEHy9hZkOm1At/C50S6kmv2JkpFcwgUkGNaaA1BoqY4YtLpY
e7KBtu4w9ECehM4NXCRJZfyLygZVL41/PJlfTak0/bObwNNkAbHLP/XBIQ8KpASt
5jpC6f8X5PTTK2NWcmgCwHX7uQ3ZfZGJLYUc0vJNSQ8LXWuGA4GSpJnHPAzwVKA6
MKc0tpiOWhwatE5AWoW4iDIeBe+uhQOrZT5CtYxLSxdrqmnOPuI1Fjs7rvV3MMab
ATdvSIMsfs3Cn7OdyKRjzKDxPLVAOrSyp0pxYGYE5o5GibNfpezEcujRAySUA/Nm
xLojGtkGdTsx2Sut2ewgVO3EMJ6xtwAvtRjXmF1iA4AFazhRFb6A3sdjLlGKshQa
pUfhheUCn0v5p0z9+UR0JW7ZYyfNN3KpEoaQYo1AygXU6cmxTZxFjk2rXllDnMY2
QPYY1kdW0lP8ZKDwpOM1jGJXJMNZ992Voe2u0v9AAieNyxFs1kJwj43yGyYEuvvF
G4EH7rafbjwTvdME957oi78IiOPu0rswpHjbV7YffwEZQe0hZd0caI+yheWkEOIs
bscmNHm71dw+IwiIXEGvEB4cuUwWv0zho6xbhKy2Sa940BxmcawwUe+hRrLGOOoc
FUz94yd1zYus9DZkwFVnnO5oaUhtKagzsCXwnND+eqWawNIxYfC5OFCWrXG7gE7j
jlq5u4pj3FeeGF8wOUo+2Wvg/Q1p0DVH2SCghBwP3IN1EAWTK8YO7f9/cKxGMyr/
A+wbqgP6KUOybNuvbxxOHRORAxQZ42Yuy6LnhVMkydN1mip4IovU/BjO7CNMTnjK
3iGkWaradXQvkYxw26ds4ePNCvwE/3iGFWrKV6pzW3UonzO2ek0IZpMN251ZRRFD
R/o1A9O53oQh9ujNXaj6yc42J+Ad9/mfDBmtXH/ia4Qz9U4EpLyWZCRMugnSl4U8
9BzqQUFel9aaViWpxj8/IDGXXsRE5w0FGWsR4T7QKZlQ7VB0CaKm9axKNnOLp+8x
2LK3o196l9Qjwk1DYr/KGOl4Hcv6b4VIYdwT7ffWaoc5flyLrQrKglGNZzD/3+F/
mv6rVfK63KvCFZHDZS1ADDkn/wRYOgqbxqwncVC/c0l6Fnu5iJPI80I7mbh9XBgO
Fzi+nJg4oiSYJK8N0u6lZVA7bR8MB0PyszMTOW+8sYhNMB4PR13Smsqoh7Q96qsh
K3BHZm0BSpP2BiWjbrFjLMv03TzOIDOHp6PLmvN6K4cP2xRKRqvoDW+Ub10yn5qH
+pfIDCL/KPWN2WcZItV7aAjOhIEOqIjuuXqjFnNmg4sFuG7M7BgQxZcv01DxQsiR
ccAM4LbClVPHaF0Z9sEpFw1/duPsuwhqhphrynTER8t3KQCvIyULXysB+yYN44l0
OZ5slfY3JeRK9D8yDk/+IKG+ORd8Z/tVzxyuB/xD3SKKb9FWtSuOH88bpzHoBykO
rqG2kRpGts0KR9f5iMrwxlFDfZu6B+npeJl0OGYSpUagW6T3UWbDBZ9InxlNH9h/
41jyALoxbuFftGVTj65t/pq25E08pCgfsBK4bez9rCgFqy5qOAJ4a8qh7pjsfDpA
+5Iygpb1CaFnycfew+2s00efH/7/btqkgL8fL1cfT03QhlM0NFOANJxE7KvImb4r
RKNhlKPP7VN5AavfIEtw70V7BS2yGi0kAHxZnIwUkWpr7fogOxpEF+GJn3VD4GJ2
MHvuNHtNbP1KTsa8cB5EzZ0+Hkm1JJbkdtUYxov4er/073tg3rRmqjesaZxUTPwr
5TIlM5FshiabqxOt61uzbtQX0BzcL/fBO5bRnVZC6YjfbnRDnx3Jm6ACaumpZHuJ
wIAD1/QJ2y9IrEy4aOhXAq/XuQFu929rt4Drf4Km8JrVZ1mC91BmUBIvTwQTfzEp
LfahcgARa2630zQZIXYoc0waiBYUBeQhmqdTLZLz9mr6gHS9TSjSdEajAhCeKJVg
0SlL2KdJj1p1FfIVxAQY4Jezo+4IfEVZRJ54ONDMyxXSqzgKC/2+2SI/S7wdbHUO
Q8FXApKaazgkDor33htqcIEx93rnqKK6vEbzX5UH0vhpP4oO3gz/9G99MkcWHpD4
10TrnhoU7i10kRXosN8EViJJNvGk4nYo4o+Ve3crYDD43LkRYLE0ufziutotc576
6UmiJ3bDFoI/B6ZMpR5czQhl6id9mshUTrNRtOLOliUqxYyvtk3dhlJT6n/nC9LE
LxLSuL7+QqvBROy3maN0nkqStp250ZLIXyLnGtThLNo2asyL7EI8WwwcVsvUelau
Uo9qUdyTb63DxM4vpz93YbQeKpPeFL4/aPjGOHRZBg66o5RWGS4CWZdctdfU0t/Q
1lI9z0L30Epp37IXg/RY9jNAv+h7NeDlHqFXud7T/Fpthi6GfyDmGex4Sym9PGlN
Krl9bKbgOvmj8LPiUL9BDlyK4g7JNSjT4OA4kbgEsOdtNcMomQcBRTk2r3M3d1GT
7cPmhZlmbFwz09TaEv3PBOwm+8Ez5oD7xEQ7BTbRyRZAckqM0N5gcjSTD2r/oB7R
DtXAypcUlldOevRST/1weUJTVlkro4ocJnRrHLjyrebNfFx6lf6+f0Eps0VIT1Ra
f+L4QiusRwsdFCRRvMeWVFiBR9fmFiJY0g66CIPhrkFy/yYt1/uUn7eK/sjfv1Tx
/AxwxRftAH5UZ5k9bhhFjpViY2+PsOaTf8glD/NXoQgean4FDymVYcXkfFJmPQn2
Iw9X1KsqCjBBIEn+pg04NO1mQy8r7VE+SxfHIhA+W/U1OpP30usHkj8auT816xrH
lC4Occ25IOYsZo21fc+bRW42YSIx5G1V3RuQ9QsVybPL3Yvc6YYcn0OvKcIGLxWd
NdGTGNg9JWhwyqQu9L1JKj+uo3y2rtMOvxQNAuthke1okG5Gbe+X2/LYduxswIvK
oy1/ZrXEROLkYlYaRm8AxYmfqp+AZUJxrhxog1VaGL7CMk2IjLEyk/pafJSxkbGi
Z6KjIgNb0bng/ytN9plqZtbTYs6Sb89iD3LWVpFLSW4LJG9tsrqj5Vvnc0DZFv7Y
6tCX15L5zgIbd0kqF197sXt4DASg/xWgaYwW7180HAXfraK6XbIW+WQv7ad4xVsu
R3xk8eG2lgD11aUbvsJuYftSS7wcU6Z6Pz3GIQhvHAyzLUHSLD06m3ZoC4cxaHPS
kpxuvOipHqpC0VZh2uEknsxo8PQ4sEkoIG4PDdc11NcwTTfdAYIAH1dXCu3dS3nW
Q0orXCqtKOg69ocUG+BCI8vBaP/AcihZbbmeQINZW+tZJTMvyMDzykHQRoYF5sX0
HmwBtHm2taM6H6QfjSgKk3iUswWWKjNVItdJ2/TY/IOA6oduJ1H8O5z4K4JUF/7g
NB9zYT307GaOc2TPepp+L7aSJ2MNKgiwR0QDRYr7uBtVyObfRn1J2LtLnRfHoEPv
7xLFm1trISF8Ok5Q9hjvXJQeuNCjatAbbe/umM+taT0xdrjWuGhHQ4RftGSo8h8c
vvvpvmPjRAAxnuBqq10pG5Gd2FRiBRt3iDJ4/cwil5iZpqsCeTSMyRUc+z7SC1OO
aWVolargqNwbN2x254h3zU8shuaxlziUYO/0Qk4PVF1I9jigFUk36ot6fmpWZXrE
w0D0qk2XUZyjsLjW+5XrcfK8CF3ur02kTpFMSUEb2JsogECJRjm05rrWvU1+z0oS
j7WSLTvKS8nJnAsFIHNbvsTuqOzUkX45BpdFvhCWvOpa2O6qXJzg89t1JFRalaQ9
uCY9sBkndgr3CcD4EBE0mVEBxc3XKZxRrf9ktUT0SjmXvc5R0yxY0/o7hMpXCB8W
FuokvTh3kB4/kabmnlalGZ75Y2y11qI0evMS48km8zrrhGyigg3C7kxiI6RaJ0ia
HY1571QuP33N8aGIo6QWRJNDIw6LN2eue+Y05PBHE3LS3TvP6RG5PcP5t+rh8PYD
mA+fooh5ofMigkEXZl1c144Nf6tWfwK9q0FK/geBMq8mYyxvGX9NAFbc4Q0W8dHS
OlRyzcPMq2jebsW09if8UKwdkXbeekbY68hLZeOwcfwTsCN4xNQ6mGPRjoNgg7/x
bcEnLqEY96EhXX9tLZNDI3cHEBm42VHTd5U/cHKEfe7Jy2Dc6SqJPoqxznR3Zllz
D85YdZ3qTFEA1Gn5+fNDsrhdTYi583gWlI1f3N8csLeNKIN3cY53aajjekMIwWa1
HnEclJqyoxHxAjq+UG4r/x29GZU/szRht7P9MrFmSJd90R5H4TbmOFeDAzcdF4Ai
avBkOnylJkr0hH99gQY3jywG3HqY9zi6NxpIjtBOMpc3ibqCNOYJgHMuIBS/7O1D
k9gWjmOwgIpKUC7Xi0SZLllrCDgbhRJobl2EIDVEcwuGRPsKijxTpEtUJLYva0bI
KIu1zWAakITaIrGiYZnDDq1fyzrEZjUnhZjEs/UwJKGhZOXT9no3GrODm+e0uNiw
z3sGTnmERVNmg44kGJ84VpK+9PMwDjt7Gg5ADmehsu82rIX4+xMgBkMdOHwZlHrp
ETYJmyKoNSduK3hkMzSNzaro8FcgZyV03zuuQvSry/y4oricWoVrgllJUDRdh/y+
v76MaxdUjo332CqTeMqLkZ8e4nj/TQ0mIxTO0Edk1UmGASmSmdGbqMIDVBSxVMjS
nbnttIyEEBD5IkALI8JV7cM8v3jle9ePnZyCw1OzW5+0GX2Cv6xoTLs//KememqV
k++IYG1Yqp4Wr1WZ1lyc9In6i/jmUdoUpTLWpFBP5eJx5LfLb3gnbsyPtRB+PjKZ
X20XMna1WpeUchp3yICAgbPnYzlHdiYB1wRMXt0cfpMmvmnscvjIuRGSV4Uo4vOY
OB1Oq2kWlHFAQ4M8xXPKYfXoC/rOK6uYnK+g1UqALv3iIAp1IWi1S1b01Ujpj0O/
5DG1y8eXF9FDNtCu3iC4/VoVtwYwuUBHPbPczme/AGZ83b96DeiVIJdkBXYvulRU
YYtocZoP5nIde8YnxPcZu7LwKOZzqK3qogc/s/nw1Dmnj7QK4YD4n4YfGvGHnlj+
RUSmDEpNkh8nTn3B9Ti4QV4fc70d9CuB22kVHvMd9CrYUg3EjNCQuUxmRv0di9SC
dF/kVg4qJEkn6BZ6rpy4p1idW8F9O+5c18ViPt+Bz3uVFXsihLCiKeO0/XTpBNhf
nav/EGbHIcC8SozgeDZxEtWNctcqbBg3H0eAqwsWJDxV2T8KPAls0Qpg/B7mvjmL
vIA3iMzyOxhzAlcFXUYTFx89Vx3JHzygd8EhQGWBVg3scEoyqJGlk/fY+5w/OmsA
GwJRRs/DzHctc5aqEZ0Q6ZCaIrF3MHGqcpLmM6IZnIoRvE6ocge91XdT5z2Mb7dX
tDCSFJ+AvmU9eLjoN72mAyCug7iUr2/m4l98h9QQ5+oUYPVq2OSjqZsjHyLilYJt
Ln9Z+Ys+2U2z45u+lvAxDw+VkREtcLsliITQnxpyNkEaSaINmQBHGbwiMnPfCD3y
y3qwDS7ESjoqO0jfKIXRfaOfRgLdNwwR4sTN5VROl2ju1EK5z8gblz8Q7TATyQa0
q4og26apvZ/b7lQzg+NuOA1IHjmb2kZq5l+HsXloSKb34nwx00LvwGeKmdY/lfi8
K9ztLE0cNzmRwj5Bx2Q65KJMq0bLsJMprlFRHAzF3uZ3VgOj8Td1hNvcl5Pw/haD
OZC/UpwHpKpTAsAgw1xCfwtdl7wJxAxOeyK6D0Sq7BAC7RW7JSxXZAa50za2nnx6
GaVnJUfSNi7XJPMb6Flgwtp2Yny1x8hV4iwHgVSmVnTSp4xyP94CZ8NruJ6m8HYd
rjnacC3ZVoLSydQthgvtdyQF+L1SqW72Un3J8CjEjbeLvkSBlctiCqTXPkKMtkb/
cbTLRrTsbQhuo223FtLOhfo25F8l01WVdGxhk1DTHCKxfoh83jwv1HUrhv5UxMnJ
uIBDpgmuV1eSs0Ov9z2DRNZKYbRNXeuH1EU2mTbKArWk4+hCepgpaYr+oQG/Z8Iq
AtxQ0fvDfYAtRhG5TPXGTb9vDIzBFAzuwlgKc+S8bkE1uqC/ZUjSL8OAP3wfEapG
GSY9MmT+9CwaOprfMBXqguV4dz5LWjw7Ux1japjkq0l0EtaDFrUczFnTPAt4sJ3V
jD+IOyJ9aJs667M1dIJGteXQpAyYUTsZ8JrHNJETqHiKT72eAlU/dQpDKchy0oNS
7J8jecZZtsBGHDDQdgPBBxpwcn5PmGd7f2Z4ZRscxXDKrnRFFusuTX3x4RNQs4Dq
KX6QMocM5EQnhMl6iKlgNbTVLC/+BXeBrYn0VuM1vuJ6zWsN6QHdg4fvwmWYnNGo
CVY5cTzOGjgXLkbQEa+XFVO0WNR9udkvvb7e4Ndm4U0vWGJkedo+mixxI4QGB9Fg
WjTGOFYH+JFA8tix52puKoF4jz+lMDwO+5Jwhad8QMwjlzu9FoXch1swO7sADg9u
2u9r99gFBVgqu+LrIZ93w72i7ar43GalXlCbpJNZfd2sjI/VoPtxpRsDnAcZMh9b
aVg9rf+ZNbLox/fLYpLqSkCqdXdgNiF0x2uEJrzzXCtHdKJzDXZsvEYF2gRbmGeb
lmMUb3WA2hP9Ffdx/W4OKzTPOfWKQoBMBqA6E4YVm+DNS0mkjYI0YVOrwae6RcaN
I8eDzwLUrzSnfZw29Rg4RKJsx7al8hmcP0Pg7yDnAJIxNM5KRd+wjrB0lGhg4QEm
FpNi2SQsTBFRIuyCag2e6qIf/rprkTir2vEWMd3qrQnnqm8GOBQPKk/ceZiOQMOD
t1kuU+wIbLj7T8w67w97VVPg6gTFvwK+iu3Po8SXtk6GBSS7lmTkrjOx2YSA+F3F
UVjYwNkeiG29viuT2eT+6FJFlVhGC06+OfOCR5f9U4LFE0HAPSfEOZO9waW/6Ug4
p33RRacAgrGY3GyXNXuAgGFE3B2PV/dBdxl1t5Gb49rNq7VXhOwObBYDWHghSAjX
20Wky95R0+U9fWZZywbYp3aRwZkMpAPQ7fwLIhWzTcf8i0fGKhyWzo3V3k9oq8ob
gb0/VdosgjDenMc6MfB0rNXU4pWrFXXATe8j03MZua88IiDG2Rj07WUkoxJMQMnn
hueD1wXupIUTDYIYThJ+EVTwUa5y9ahMlfq3UVCRiZZ6KC2RlLeys9d+qH/1BjkU
eTBAIRGGiTVCgca+SlcUUFfdP/SwkkpiyVttxWjzxftxMEipugvchmKerO21Jm3u
8QG8AGoqSeDFMqJZ2SHnDCC+oeAvugy6lqYY/KNGhPp1RET8dju3kB5RSLGMSke3
8xqks5xYYlVsurnKwGGS0Jup1xP3HdYSMtbraX/N18zNd+Eq9cxDyMmAUJ2tgNjX
v+ySrGRlTbEgOQ1y795xweF2DtItArOES0sC1CLfJCcXHkxFoPK4S8511V1RhoI2
pN77RHLpbnKZbqg/gbHmhLGHdDf5aGdGc9ab0X6SY/nYHaf8Shv+tmpZ+UqNEYLu
04DXH2EZ3gBJc1kEDim5kfaJ3IiAC38+2VaKfut51HKbmSWg4ZBZL6xsuqx2hurg
+15FPxd9cc+42CPxeTLyXF/NZ2L+4F/EIeL4m86/Mv2FONDn/nnB5wF5P/oj8I77
Pl9dd8jGHrxvs3XOxAFicmu43Cc2eSaNJvo/EDVVmgyWX33YhX0PH/NWamc6vZCD
2TiWaJDBY51av9C6lCkeAZpdy+QCZk8KeeoQ+czjOwrc+BI/WJ9tSzOcII3b3nGv
HU1JCsg2EzdIRCmm2A6nH4SyirMH8B9iNl6rl/XZuc8Vl9AySN9lSyIBB2Ny8xE+
oUHo7d0ZjgeEFPxOC2lN9wi+wDjOQZeZNS95zqoap90EBl7V8npsPIwTCe3owvPT
sZLL/yeZS4RT/RwbYrAiGGBtLe9OxynFg5svxuugp4fITvaIeJA7ROQ5F4mhNVBC
dRi/U9/GSprQYMpRNtpgTh1BGSwbhjpLI8tqWU2vQNsFeB6OyO15VKlHrQBaGYZD
RF32g9K8ybTjtA3Eu5hcAAfaRvJ5evN5JasMRO/FxR+01f5BdWIdiXw/wQ0fHbeo
vq/Yc6I7YYvLnx6udcyK0k+j4tmiyiy+6iw8OAPZY2xsihhEMw6ZPjLEWAMRTmkI
Le0AkBOpVBMoZLDzpu4piL+IOllxN+UGFL4kUHISkAUGYGAk09sCmNF+JWOlMW+Z
bygKseHu8MC/k4lAkBU1x5wEPJuqrJEa5Y+AkvIURu8MYDBerqT26rt4alVwciw8
Xcsb3+/1qkAZGyB01yD1STo3h/Is8ah7nAoaOnRTSyxEvhg5n8m1/bpVLUmhK9qO
3owIjp3iF3+djxQaXRYbxgQo8xT5i+HiYy+mhIKYUtLMUCNm6zFoG0q9P8ZBOBGC
WZ419P59Abrmx9hqBvxgMIW3v0Z9r2Qrk1bdFTZo/bmllxApoXD8O6TKxCKraAgC
2fr67Ms47Ej8U+j9wIcfdoouH/Tj3u0Afpt2Vj76i0iNO5nDfOo5rJoJCBc3LIrG
RU44AtLQMdIBqapvOVMU6t8TmjH6YPTO3ZssCVv95UDryBs57ETyuY7EDrbGwWWv
FqMXDWQVUlpUiaKVS7myJLKmFAP90Xsz/NWS3cm8Wf4486Ur67Uebp9Jeiu1YXq+
rr6YmI57onGKzf09CK9HTpLbkanfgYw+C9NKLADTeIXnMtsKFv72Racc+i9aBnM+
uDFhRxAWeEeiw49Sa4vLbfZ/uHw77RWvQH+ju45OtvR94N6KH7j4mo+1xzcYixrz
s6pPZsHyavqIsCZiak2ic3fMgyxKSbZdUg5JJmvQ2FilAPVuPgj6yMdpBL2Ouy1D
naFB+093/T/+6LCVcMWSzTlbNZuFx7sSQoGXW4wYfxDlbQfl+SZXaU+InO/I0Umw
OGNqvIT53HhpUY9TaUCiTMLWU0V82dCFjef3LtuHTIqMdsB7ugGVEDLG55mDUuNO
DPWZi6QbOVn90beyYDhyx0yfqdWsEuEilyARWdTw+hk9/SF5F1LonFiJu5bg1K4/
/FbZYTCsqFIHqkfwjOnEiL/O5qeDoNI/bFV+6c7upcWoQtqnb0nNW2hbqwkZZkEY
5hDJRj6PlyRmgy01kIaVklXkb0riJwlMA9NMoiEHTZOso1CFu1tUgAw4qbJgA13D
++6UKFralTcQDfjZjWiSyhalTZ+FOQEn1vNbuQU15SZg5srEMjHWKSX7TmEpWjzN
JldTqiJWjHc/KI7XYAsUfv8fwKmzefxh3nh2vQxGTlfIPwmUyv6Kc9B7epRfVEkK
aV1r3reEx9l7R+uG70N14scvXclQffeoRNpLjx+7cwOqV3eORVe3guHcp78rNPsV
SmQDWE9Du1OxsKW1KOcuAvS5E3qG81Vcw5ah6nMzGy7+jaWqDk3KJhmQncQEDwsb
iVsROm4jKBVKsbgz5pD+i8XJ/UsucQLvYXWqi8OX7S881YgTXn2+pFmWRROZbpRN
ujaZuT9XNiTGmPkDAjK+vUBbSaenbLTkRCOlBDzrCoZVQn7kQt8kQv0MLfct7RGB
BLvf0pOxkIjqJmGP75lSqSySsWa5cGufHy8oFEjyAStDTNbiTYA0ZRoxP8tgMwNC
U2xwSlScMx/8V/wAdzL+fnwlFliYwXx8MRF0UMbt8/YwS9E9tQz0lF/xlEvNs0Ln
JmTHE6uEQBaAfmrKdrXhIBhkQUoC5AK+f8oq4R0AP4JCoA3tNKDj8eKSzDnuAlTt
RAbN/C22dkXbKOz4XhZcNAai75RChWhXpD0D6ZC70dYloeAz2YiB3AHZBMA+Txye
lSdwxAiXrAlfEa3e5mZzJpZKGWYlg/YjE9YNXnRoikohymC8UI9wkEsC602HmTpR
WYbZNGyTj/u3naS96kPXiK84EYlPCYlOrmh/DHAaA0sZ3hJ/KRxozujgnCcexf3M
cVOtWYnhF9LQwLwMivcfSMp3FexVNpXexvd3KiiEOXwYXXGP1HrbZiwx5eoPOkR4
RySLAgMkMmhH5cbmdzwr2RkGUv01/MyNS52eGHO7K0CcLltZNPaK2TTpFDp8ko7t
Akw/QMH/c2TfRq44TDfRGWScsAYB4EZb6eQaH9vnujkKOeS8rMHoPBZt4Y3YEo4p
242Tfg+nrjnQe4FatoKijbAiKOkx45yzlxu9BqyFdjrotvunUUJ+KRrr8Ko+LSHC
FiMLhxGs6T0eT+Qf3fLSx692RwAw0gIaJVNYoOYrV17QdyMp2u6c2z/uxIeHFkrR
aovc2fYzxkqkH2PcHrFUZ30hKp05uMca6KhuM9hpyaGgoksSJRuRAeVgAbFgGMNt
6IsPigYnyMVY9mVAlpFJMMDI3zTqKjWwfsfo65af+dErxXDvFDxdtdgaV7yu7Mgn
c4cmLfygZaK+akJwB1lTO10CZ5JBCJhl3d2mgG9yWhw1G5iL0l/8xq7PukcJlH/m
ntAb/vvuZt+inr3zucUwy89Opfl3noMy7DYsaAuYcA6QKY8d/g0vI6eDW6vGK6cH
/4TKv2jPL6stsQ9EIt74cpPpk/hRH5o8zAxoZmT4nqDnz4VbNDfG3MTvnDa3MCQ2
WuBWCxHxySX9APoVAuBkDzouqKU1QqGmZjM2PnzEZB90rqpZd/de2OiuklKccmy4
4qJqlEO6z5H+tsEmPsmHwXYonoWrBTiV9DgVfE/vWWj+9zeLgbvPpbGe3eB54E7h
NeXhWLtk4/bv9k9R/2orRFrXskT5JlsoW42YfU2O8VAAL1Qye+tKgNf9JT28DW0i
xs2TJ6BiDaVAvGob7ghlhY2PE2Wx0KOHksIpCPVu2ZI2bhNtZEPTD+cpyEH1NP+b
V/bz6UUCjDYS2MLIKwVqEV6vsfNZ1Z6HLpBwWqibhpUNqQlL7JajPhrTiNjjj9Ww
ol1GkTdr3h+ClwG15LNvA2IR8Hsb9jobl7NydqzJVYtl+MUZC3tsrNLQfWH3Xik0
TyPyjtpMj1U8vq7bUkGVPaDKStlInVBHMfNJtAbNqZ4F3YQoQHkWJSLtxA8CKiFS
IFBDRokLWS1VGJ88obMS6ZqzDxBy5B/uuihSEqA7LowU/SsHe5o23oExpsY8Z51K
uVw8c+ESDoTbBnm2zsmfJcgJ8/bmC8etONWe/ftmGyzjDZbsgFANCA+mQS7Hu84y
+p+bHqwbbKIFE5K4569qFq0Wt7ZdlvXp8KnriJpi+qVsISekHeRa/Zae3KwnJotH
ef++qfzp23E5JBeuulqnDj495WFywV4nsTz9MrMSxvFcSCzeed59/N9E1KV5ldkS
7q0oJ4f/t9/HRrfILZggC7+9Bfulyr28G5uHp7a1/iCvmvQ6IWilMeQNJd/Senu/
8gRi8sa80XxPywB5BufX8MxiGwKlo0G2Owx6p9rRtfSZGG8HmAZzJQuhaVNslsmu
/rRUO/unCyhYRS9JpxJ+Mu5iEE0xif/5GImrhpz0K69up1HhoFPc0o0VAGqDAdWN
p3Dp6Dt2iFxP6dXJJ899hy58StL3HWiURZmcbId3xjgsq/F6PPzPY5CQhqgW548f
lT/9WbACh/10KoOs/VGDmOBmjEw+VvOwBhzcrUazB0Gw+AUbfPtXE0Cdr6KaZFBK
HjqBJftbfqDkxrDC6awGw1xIL6a+/vyDTcn8b6SowIGG6g+SwMu1TsudKUfdo/iD
aKSDcOOmvrerOb3HcuwTqqx9IsozC/R2uZzYSwCTZPIB0WLVRoMFzAeAK1RdzKu7
bNvFpom+WmdQWUxCvyJWud67P9qC27mC4BDj8PgfOMw1ZM8b4Ow8I6nXICog3M+P
8ORec4Z3gZOb3EwoiBfpO+WTkYGhf+blyZ0KIzxxSZGH0/2kHTcTdr3zvcMIN4y7
zgUWP8mqAFxy4zLXzyeMKTVqFf/74taSCVHi7qn4lEeB9I6Lb+1CCrYJ6sZu3JRh
ZKFwmpYQUxdxeSZsrK7m2B6VCoDD/Boa78LANTuJkcNoPlNrUNMOm0dRj0L1utNZ
+EueX7TsdRsBU+ad/uB6i5gaK00BaRgskjmu6hNd9C8huDuB4Y8AQsCW0edFbG6w
oJCOMpgpxglGZEdTB1z6V+lgSGoubaUcCeEP303MQgp+03Psgrz3JnTKpHDrnb4W
qcnH4BI30J7gJnsSgWh4dxh9unref0C0v7kCTeZ863gP5T4RndfK8LA2HXCBmGwR
05GANHOEXbA49xPLbC7dU6D/xhXdfNTs4Kgp5+WFhQGM/NLwzy907lXOpf8u32q2
hox/KMRQyYK7XFrRxB4BukOU5vcs2fFwNy2lu5IhS/W4QjKO9DRp8vk6MIfScXyP
YmHH9C6yt8qgz+6DgZGb71G8awmjd9s4i+Zna+0oqwjLvAZwTPF+TaxJJ8CXRsYC
hLADm44HtOrm7wv+DY+0nvI/YZTON3RzEgQaKTb1KwxTBeZyZH56VnlBWZuJcumc
WmZGVZMeRf52g6L5rcaFxNPK1dBDa/wMkSqYrb9RWpCBFBfl5WydKf1zKzkH9s4t
5IS2gSJuWUR7EdMoaRKAw6JxmH0dvHjuyESY1Haah0f2TbTPm7LDk/v/PXhUZhB6
NllcPz39gS30vmpR2R/BeN8J4YluaywCwH9wm79I8by73+sYaKxJ6EEE3tOJpcue
JVrGJbhCw5e/HsrVq/Pw6NSzPLPMVIC+bKg3KqegxMfA20STUJgZbTGC6IACJhVj
QT/BeoYdzHUTeYMd24rZ+L8+bePTnU0E/WA/sLu/6mxXIubiqUDygK6pWlDd7ghP
EFW2PYFwSepdz/4Oj5/VijE0QUiehHE93LByQas87QLw+roV1PugsDUvqyAgntbs
QRQwoMS2XB9nj4v+Fio9tBfxZ5CFJoylw0axmXmyW8WdRZ+tQ4qXm08V0rabjFL2
sH57x22dG8JMSJ7I+5VvpDKXGMfREftfXIW4Cs5eA14uH8j2BtdTZpusv/Idzl6/
n6N2Tbd7GTOBKSdWgcPbFhUKbF05+iGXXU2tlewxz1haRMt1cOAWi7vVgHeuEMlm
Di9wx6IXYz7ZKry7VlBH9g0W6+jjqrql8+B0TDXFQnPRL5/nXpgrWTlR+Sw6bxIf
5zgqVfCQ1ahb6bGv8zjdORe3N6O5sYbQRTRy1a67YZDH1I8zti3bc3Qz6r28n3R2
je/5U0BTLBa2PzBz2sCHctOBwJgoyMSsRecBLhCm6wTMlA1CPpMjt3AyXIATgin4
LLXs1DtPEN4CxvX/SgHhmVQsbyqn9Qf3LV3QmOALk0eg9gY8XN7Cz/bnr8dD0Lpi
Jyqhd8zxUJ5uMmZ5LQv7pQrR0PJ43QfnZijVjLkxmskHs3pbnoCOx0SlNEDvuXU1
/FbNuPXGcw5niYwS7GvpfGQ2OdayM2KeiJ5RFeaKaGza4gzKALUATzihsi1K1WNV
vSL5gylHprV625IHAf6bvanHntiTTjmawGr8zpxygdkCnC6YBuHw7uDVrACY82Ef
FfDyjontHybYP41/SQ5gmL1WBSG8hfMeYrIRaV28TNn+7P80GNKP82UduhsBjVZ2
VcX1tuZaUv8goRP0X9FObkZHDoxJCRcsr+R4mgtx9ZmjxgGIiTBGBg30iye8DYgq
HSKvEoD1bk5cQKLaSDplzDvCNDUcKrLGuu6G2WcLESrGbeFKE5bYTeGOSgXqO4FV
0nldTUZL1mei6goY7hjacQ+90Xh71gfUUImbrOYMc/ELF3boIltrQVfpygOvoTvb
WRRxqqW+G5RjP5grePiq8ikXMjXJXrlqX9fEc5C+yuruJdajNYPRGTZss5654F1X
B5vmP8TCRI16TN2LYZeAEToH4jlIkIYTMdjzSPEDlyYccJUP4CP56Zc9RNTeKGP/
9fFYhBHgekpOQqGyHjsuJu/Qvs8vAi7o8yYsesMuvmZIIbQWd1ze0g4dOsmDuY6v
8QbZg+KnSlwEThf4QGaBECkJrX7bI2RgbtA6iZW4T1lmwG0yUeGhkDn2RSl50M/M
JIEIPqCvX7/VdDX3ml7UMmpz2qaAAQKmcwxCYYuNkleqz62hzy3Hck5S3nHePO80
Ud1deW3c9yhu2QANQY/dQujByVBU228s/pyAHdlzSwXmfcvca57Fx1C8+WbGYn0l
CuOSldtIINziJ+S61gHL8tSUrk224I3pkNdw/H454uh9UJb8eNT7TfxmELRWm7UV
p+WAmyNYJj7QSpvd8mX+ZFOylGJSkqjL8B6jFYScii7UCNhvz8A/G4Q4+G4e0f9j
OeH4azuud8KFX+Zwz+Eh4ByRDCh9/YJqJWXabTfwt5GAURfff0HsnPTv0ZuWntg/
v8qFRJtSHWaCtM2UPapWd/rA9Wu5pj3sCZHLOYft4yM8LPt6IEaAgT05c7q1qOS3
cTGF2sH9bkN3apDawiijZEVqmBukScJw3UaVCOxa6TfrdaBiL+xLqaUibqTmYXEF
HQ2DKKSlfx1dp7MDfX64l4WTTowpBTFR1MAI8eJmeIl1SPfA+7YCdYiuui86IFsZ
mWIAcEITGBKd6/FZEhk0lanPSwrv1SuF3bni8XCXCSuhq+IcHgkncXQXwbgtfZE5
wvXcDkdeNQXQz85b8aRp1IGnG9gKaZuPIutjv5hkSsjdoqqv+hG23AYxtrrlFozT
UVNFTIcXJxGp6oF6lzgAfEurgEmyuETC3rCX2PvOWxt7uYR37Ic4Gs/rIhKPAUDu
py3njNpifI88rCca7AwuDkogWKJa74Zx9aNkyTEZA2RXfOqtH0eUdp2oQTM5roMG
RGDsc/s29kMYd+dDAGnqG3ER0XUtcBPF/35AqemSBmf5W9WUUw4Md5DgtBMBuAM6
0Bx3PJtq6C2ZuJ5hEKl7fglISKv//lFjeDTH8wQZQjuwYssqvwk6hJ/KANyZC3iP
ULLZq8uvNRNY7L8AfZjDmhY+WDI6m4qLkHnniuDtsIkZlqQkuEjbq54tBB1T0Nc9
Qe/ymga+iNhGnmy2yCzcaVNO10WG/E2fmnc9afAfAF3E0uqcxQD40lgHUuBCtitZ
kbWfgxlwOPkTlXgMrohyzmQ+vGarQ8rFPCwoobecbzl4C1hlc704OQp2/Pz634P8
LQF7H9CnIQBmwDj/Iv7h6DcDmR9Y4hye1vGdXNqLI6itsIZzKD3bJj1eobGLIleT
CJ0NpUDsLukFJMhiZbcxQKb7G3oCqr7dJU+FSneuYIIlO57S4YbqcZRJSFIXd6H1
SkfnfSzJ59ThFZ8DNQYuuXNhTSTWebt7MG4qitkgQS6LsE5eMBoiqf6ah87gFQOP
45byGoQ8ucDIuvZYqbd0sDIw1b4Y3HJEbCYuQ3CYZly+2SJjKHuYJ7uCz+I7XHaC
Sw+A3GEP/xWw2yeoil8PYX2jeIp1ay+mLIh8drNmoIVxafnUFL6E4Xp4quPFb0PH
dgt72so15Zf9DV6jwlYLE6T16xFFc4b7XsED097SeTqzKIspJwozxKv10yrwfIl6
dkabE4nNr+VR5IeWTl/gvImYpAxJLiZ+c00Xf+1lPnYe1qufjHjFYXu39g/ogtaq
5Cou9E17F2OvsdttNsque0sOw6gSbBRk5p9BiBSJdc5cuJDhqGHkeSD7yFqld/4g
6Gnz0fDkUop73JN6xZuSWzPncfNeokuBGYG8kZa3gQwqb/kE0zh445C9KKfYfh2e
96ejHjx0Zh83EFGlyp6yZzb7HTiK/ASzAmdXzJdnUlFlJavL0fA5fb9uwuigq+1N
G7FB/hNPPFgmkhoKQk/iS2agIUqZISXJVhSU0DId3p8eQAqrci+xx3vKDH+4rHOI
q0wVTNDCc4h3ZUH2iTpwAlWKSSqmCAA0BvzBVwR9gFytoa70DrGbVW1B9VqFLbnG
j7myhtVT7O2YB5h53DpZx36PFde6UhAN6Byhw3Q4UTQ2ol9MnRUWFhtE6aZoE7lS
vis8C0cA8/bDVkO7eRMxww3MlygrBgUNwaudXeHxb2dExCxc0+LcbAI3HuSaruiC
SZ45v/twhsY1zIjWheCJCa0sQcUiGp1938HVsJK1cv1p/Lpqmrinz9FoRTXuZGHY
tgG3azGpe3rN1RxmHkBphQQuR2GHRvwiOaUp5sSpYyC04ukahhCkCzaxYA8jHqdF
EB9TOxTW1l9S040B51OMj6h86bzmxK4IpajYOA1gsLGGgi+RyeJ6mvab7DAd55rD
mgWXiTa0OkQMhvymmKiL6dZhTVhyWY8ftxj697euFzMcp7JG5ic4AOiO0+nqADXf
31dqsizR5h/+USIibcDZ14o7UR/b/RVP5yd5dcbggF/3tCIyX6u0cbL7WQsRn2IG
F1tZ4pDRz6Dp9yOQ9SEb821fEr5ypLmWDqx/0N+SjUuDuUIU3rr4gSes4hQgdX8y
zww5TjW3EHIigU2gkNmJO6ofmIgU5t3sqFygtrmLyoK2yu+kQvMkTwEmbf85mEv+
qALlX6/cOjVMYRS4VsYUtvXjZkSSC+ikq/60BW/PWU8w0uo9izwhE+kmcm+swkRa
wEvW5PB9A12RNCREIMzLLtJ72k972kZTai2n35IKM9aj8OWjNiN0zr+tXcTIEwc1
jjPc6YMxUVRCCGyRpAcGsjY6f7YPBG/TdS59sNV7i2IR81iZrMMX2OIsMNeJeNkS
YTC+wvEBxcAtiz36IvMku1HEay6uO8D8q2n6f1in7+9qBZ/oKDqKcz7c9/11ekHy
1XzqaDKLEwd8Sk2OUeLIxqFlwBy6UmDDzCnlmnWcHQZAoMrDAScHcg31Dux+7zZn
YBSE7XgjnZ74YnRpmx6hCiUD9N3jh8eEobKHKOFmrYwZVDZxlzfyIRDulWdONrhr
+KlpXmNFKqnUSgCcMRBCV0ldtP0OrwmYy95s3o1vLSI7fSdvxH8HikS/0msX6R0+
3Ofjo5CsBlriXYcWMVOCz4oKu53++oNvYgD0UrxLmtPCGNCBzaJ8CQcHAFZJsbAv
RaCN1c1t8YH6fAlGkmU3f2Jq8P3aFLPAzLj8BcQMcqkiEGIKMQAvrsfeO8HO7rbn
+uDuqOD30x7su0AjG8EMmkLk2DbbaMxuyaWskt+jXSpqJaKrhW9rkh2tsncRIlae
NULo6DwIUC45NbuSttjMYeao0hiXOaMWDVI3/N4aHHgtuMXcxercjth/ny80mq24
n7EFEv93Fd04eZCqjpYTHHWYaUfOSsccQEC9FCTj44qQqMRnSo3Z5qzsJNdZkGvi
gpMkUPKgXY3pAJLPbxZqnr0EJLwMPKUIteJgAFGetXoI5Wl5GD5K6VFH9IDzYBLN
SyxU2bur7027UtvjBGygoj5CP4hlQnZfejkkuK6f4u4sAXX3C9TZQoysqKhjafZI
mJFmr84HzmXCs758lYS3DpYlWUqowsU5uoiRrKkcTZev/xvqMs1Kp2Ktmb5TtslV
vxhJRVSFzLcTQcpjYh7TkFnFiJVubeeSBtz+Nf09fQNS5bYtxhG0h+fRB7GfsOWJ
JfdYUp1USq5Z6rzUaeuP+/RTkgqY2pgBshZSMvUnfs4P8o88BBk55yj8dRR3NpaT
Jo8949BtzkJZTlp1tfJuWmoS6hyUcnwLdpYIih1AuxbNP1Er62v9iznaYJ/grSeE
qRefObOe1rmojECfGr7q2peVHStjqh/uBjGQfPJ0/imQcwWeMAnX7jS4KNKrnCQr
JtDq8ojlmoj+ubICLzvAzDTLRAcSO74qNvUbCbYlwaJeJdhe+ghx+vFU9kMT8cYZ
Ff/Q+IpsuH9ha56NrNsCiHs7dP7l9hv9Ss64jdhkv1xgEo3E7siuWkfkm8XVGWUR
BsiTzy3HK39hMLWA29KAVVq5ZLJ17C/+zgXgaoO1ImwnfpM6LTPHpY3F9xfJMFlk
ztm4jqj1jw2bl/3/cNeDTgeh9v6zGbRaQl8+5IhieJJB26o6tMhS0a3GJ9HoOoxH
b3CLcJdW2X9BWk7vDrMlpY1OHJcwLAeAFAr9B8OlYwnPzIsjBENIohRCmsJjeczv
wOrtlrS/3mkbjxYN6geGio46oet5q4a0/6tVxn2lACK+VgEAGyJyNoL/WDfujbif
/dgL0iiSn6QAqGp+Bgd668B3nHMG738GE9qu4PqGu7YoLQHX3HUhTN0dxjtwNPRi
yQhguLKc91FlKXGg9pGkkM5B2sYXWmS5oX9wGqpqKsvNv/o7yt6+dXg7JopF08jE
x1eJnY0WwxqZw4tV42AScUTqq2rfKMne29Zg/eYbrfRa/TwbEdF9aO0/2AHUiOFR
KjkoURpKuVgqfa2YHQtuvqclhhPM3vuuyN+GuA5jijHyQCAal/0u5OQ0y7AKQSf5
idIHHu3j6tRlpqMoYjWWU8LI7pJS/zPoHPJHQaFKFwZFGST1h+qeHNcHaTK6TaLF
i6No4wXPJMFmUaSabFOBclXYvUtYIyNOxPzhrMyCnzT+4HPN1T8APM2tTlBtjATw
WQBpzK6/Fz2xLDgNeKhbpRO3SVRcu6hgFrg8OgQ33Rdld/f+coAnuVg/fjJ+xUvl
I+ONPlECsNaCchm6458sZi/HeDa3TIt1CpWyU1ssABGLlelPJM0u2iZ07rcxOpBk
U8Xj3G0mJHB5lvCGK89wK7N5ODcQsyYgs3CVmyARflHHFDzptnogfl/iAIsOY3A6
V59cRFiS8tT1CH3Lvvu2YHrMQbB+bnDvO/svLP12r4Rfo6DKaKF/aBpX5nyEE8lF
KcAVuYYEyoNjoEOuFw0okFxgrR9QsOpiyEXs0UFGUDzudhCTNv+swPQlusNKdWkd
FSX+KvgUUFDFjYWoPMPJeXDI32NQ6Pj3VM9NdsFhcqn9InZwtbKu1h62/oewmkiy
jkVyMQoOykx3PB714mrWiuUnmriVgdls3wXq62NgLAG5ICBNqopr4KclJNhcVfZc
TTCkEJPWlQFW9/jaHzX4Dd+0joJVdx+1aLVcsxC5XWOKAmyZs4dtlfVuHYg05d5r
w82aRJcJlDc3FD1Krb0+MKbQUCYCN+EZLJ1+e79huCUJ4zP6srIAzGtreJpZ4475
D1J6xNHsh7+XUqy63xEPtaNBkGztryCCWJXfQE09INhyJ2YeAaEDTMS5pFDJ0wvy
6/qH4MJt27xP3UUZZgBYsCy6w0NTpNRrreXy46lT5JY5QPaTl4k17fqjHXGSQCFE
5wFipa9v93FiDu65kaGBluZ0BG5Qht+HtF2xUJig62AyVCQjT8uTcOlYcvYSLRyy
6aci5yvKMEiXcFwKvlmwOlD46eh9yVU5uIttZRJ6TYNlhEnqMUYvaK7X5Uxt+LLt
niIJKQrMmWSd4yUBVb4WWxw2hzaI9DCMbqgHzzGFWi1V3eMY9ri4HFiOU/WLrpSd
zrR/KTHT5SRBRaq13WhpQJCRbRCBnCcwugrTCnVvp5xPwkjy8imZzIFF7r7dPLd1
xmvhw6Pg1U4Dz3ebqwA9reoQTJsChmnx3Xb3uAdOokL/Np5pIaSRJ9XhJtHAy3Ih
+jnZLq9HyQxHFf/GRRxy1bGgOvGdXiIAGm7kZmLbFkvVx7PDmHNSijsVOM2v2S76
9wOeRt8D2wGsZ1Qynre4v6oX/Uejtwp6hcJs9g4tzcUnqYv6HVnKHSIp8SGpgrRJ
zOiY57gOKMZbziNGbrExi0gLdjiIyIu5VtY8A1zhM3Na9pX9l2C/CFSp1quFDw2/
izQMVi2I72igE0bFdOh6LsecTjaB3HVWSId1Om5aa83lTyUyr2pTovipAEMhll3M
3JJYT/tdVhNtJP/RbJbcFQKOnI92A+SyLffhCeYQTHz1inJQeem8Rcep8aM3PbxV
ydwHMveyxu4cu7+bZZH4znYE/BXra6jSNyhrTYJIk3YStZW8o+9L1qzTyVFVF/19
TLXfldtp8Yn1wOb1cOOhb+ZQ6Pdgj12c/hS+u3dr+o3mI0r6x7zrsNiChvDjZ529
/4QR0wv4aT8MO98e/K584OwFcfghs3nA6P8n7pJqsRU+V1IIKRKiN1WEptVBZ0sN
9CDy4OX9Nhi0LztvRE6KmVYm/f3kjfdejfarkAA6hLWhpOpXEuxxZw9doO4evfYW
FOHxTjDn+wIl7ETJtuuyGIgYmOjwfjfArRtFMzeM26nmx17gAlcLuhn+WBpLSSuv
CCMnUMz494vND//DOeonYA6NYvfcq3QRCuTcGrimK4PUIBBsDfDsLWKcYVNHwtWj
E999XIH7yBBf0ePg0aV4GRXbMPDJ03lPoJdzNRdZftFIIjqZJzieTmI/47XEgQI2
/+fyzrwa4DZHyAaulGfoKoOmZkVEYrq9f7d5EPX4yWpWYWTGjdnBF0wm6i0R55qN
k9D0at+Br3+o2s5bBOD35X/xiHPy+e21E6xexcr9oe9NXe+WnUURl8Hz9IIWE7d2
nD97wxvtPshuUabeXbnCAW6DuACMfNHP50axNceTWNb8f3LyUJk3S25Q8UvEqMlW
5tMLOsGbAxo4ZEYpnTtCMW8LXJcYFIDfwMbN8ou9tMIIt3fZn3S3mU/3/4njy2UL
LwvITPqYwFErqMW3HLlbGqgsUGLKSRATPr5BIgu71g30ulB9QXEp0eacKEf3qxvJ
munoJW6DMghr6pCnTP6+GgZ+4AJgMQOIfN+uo35ZhR+rHFYGuVvh2hNhFp6tyf6k
RYZuxWv3Hc8IEu6o1UFDj9yZKAZy/O/PDdY4N9+aggZuHpBMFuKpVfXyycd8+Cqz
Mh6o63N5M0/Acw759KFn5e9DvpablyOfkLl/r8VaxQj/yzT9ExZgn/ols01dz1iy
LRAaLyoKJlToiRguCqGr2dW/wjGdoFVf3gnZgItfVWSal5WLehcuSoz0auOshHb/
WsJGODC0iXexuk+qYb/JKbOi7jMC/R0YZ9jqflezjzX2eN1erAZacYS8rkKbOxtk
v5jxXQPGt2Iwq+066DqhdCqop/3Ha15LcSkljCh71rZPER7Kn+3A6/hENeQUDOWI
f+7W7R3gY44ArISQIK+nduXT/5YBG7jUlMLjN1hO6TOaerdkXli5Lg+Oskzql+qY
Qz8NBBoNMskGZgG78sOOOyTn8HZdtgzOAl3co5nAAbdQ2FwFyo8g0EI0ZkC/7K1D
WFM7UZTjab/nr6AGA+CcjASPwPCQmRlE/LexOMC45iejQTyZ+/XQCiHjf5ngs0kR
js01MbzETDNKyifv6xrs0zxqrnZu7Iip7LE7JJfMHK0OVFHpUARZqaW1z9RgGgzx
2D5HTrFZmkfp/ee398PNGcE5QRFXvTX1nFABbWlWvxj8ikKIc6/VZs310A4fssg4
z/gKSQO22bgsDjBs0G+oVgILqmyRQz1zUJHqn/fPrt4mXpxFTY3ckqgv/ZFkJIh7
Y+RxUNvCq3wzCXg/0z095RDd1Bx/7y98z/4qkMr8LjfaG6ScC7Roc69t/j6A4af8
HobboNJAN5rXBxkh5g7HYI38mdLh88sUmF1hXwDKT1pmaiRAdUYUis0Y/s9sTBYZ
95ICJUZJeOEelxyRHgD1U8PWjz7N0xuC37Q+6c2PMCqeVM7rhTfOYcE5WRuCZ35D
03Rb9TxWFQ/bkj/bKRW/Lgs4Yrg6C1CMVRReTY+I9YNMcgBpS94ozxinSV/FUyeZ
sHTPF5YypnzMFfAyvRxmnCWqko8ptWnFI6L4obTNml5CFBetRuFKAXQecfpVpwCu
augvaonG20NtpuL6K+XK90XkhDeyDsIKhz3Z99Bh6HFo7/1YJJy+Yj7aQh13k1Vr
w0dBunt16JHPPBUpbmAQMzmYRtOiDJtkTQaeaq5Ky4kzJogd1W1Y7xNUFhXuum69
46VYgiVIOfNcoqxep9BcFSziBLT9fdRcNQhmAd5qvBlFQthb8/M2owD2aDkhqIxy
G5mqDxpNoZvYE9Ww6+5XmzaRC8zk6u11uIRuMBcVb960psuKvnYtbc2xJ3sWIbd0
+00pWXFqOEJG2UWhXS54DMJD6b5s7Bv6wgoprcjjwwPWZgiXZTFNdJbS7DKu4Fez
jSeWOL5DT9W3WajD/i2H5UwvPH3wEpTXmbhRJHlsGpniY91K+sCu8RwFzKzPNmxJ
dcGYaZzCnduL01/xoZahjJahWLuCYZGUX9+81g3xVHLkfmSwRax/ukOKHdBLvNIS
JnPer7P6c1mguqDQCs/EsDLE0IOnDV1nDccqVoWlu06B08rZ2LHQz6/p26HQ8yjM
uhSFq0Kymic590L6AFrsmrFRtgsK4UBzZOEVx8rT8/Ya8K+PsGqb49rmfFIE5vmk
iAZEJli7jxxDhdBDh4JTr3oYv30PFhQtYDGUCge+rdz6VbCVoWEgQ+Z3UTlEeaF8
eBhAhui0aorqTh9vVb00X3rrxz00tDdDNl42f1Ehpt4atE/OafqlBThLSEmuxOYX
b8VPIJclrWhpYz/PTKOMDDrk7LaFxrweVrJz+/JY+2tRH/H7HbvU9TmuAwJYwRcZ
2ZipkA8pM7J+66Tj9Y5tMkZJ78y0gvrzDfvoCsDYfbEWF/zredkVIyy8dDC74uRV
cE4z1OFEDHT5d+y816s+J9f25UlJJUfVbnGSsrGVxy3yfaP2onLgnOfYyC/QXsMu
mP5rCU8llEzikmSYsOcgaEj3LXIT73FL9FFp1uLkR7cVLbpAApxz9tbER0eaXmml
ajSbWiRmAXz5FBREubP3w4ukb1pSnTjk49us8SE/3ZLzwrOrPMeZ1mYH3b/0eFM7
9f++LIvYt6N09PNxarxZHbl/nO1jCFakh3/xYZwkZ61nI/14REQeP66cJL5hyl/z
h5rfZ/guggNtgz+QVJAPnFdngY2yMUowvllq33GGaCkKQOVJVeEiNzfzGrLWRHqP
378zRxAtr/hXcxvl9TXyWFIw5XyQQRQzpaP+GD52KzTQQzGjua4sWuwddA9OixCk
tC/rUoq6sECVxHSRGLmMLhmhUKqvfx6qv9cLA+TihXnsgLEfdLxxuShPi4K6ojvt
MfwbAHt16VonoqVJLLb76l4qPrbVm2ESYvZQ39UXnmuU4gT02KWSuJl+UFQxCLj9
kwmGHrN4ezBOlt3V+i0dTMnsphd7zldg4TEL6BEywCli22kJFewqvtPTsf4R17GV
G63DgKbQcdUVVy/nB2rWHRs8FP5cemEnb/lk1ZdOTxrd2nbTWCdK58bieFDs6Lw1
MXqznBcfngx6P1AqzvpjYw4K8gTxaHFE6m+l9iX9NUfKhzqhB9IztQ9vIwBpEH1L
Z8KoLLlRJy07t1TRYmPCWKkHgm2RFloKfC5i9DtjVsXdE+mST3KarfWFvYHPBBh2
ms87mRZ24ZQ7YyNoS0sDALhzd6irmFbm7z00jm3aMdWKAIGc8KrlywPgxvC2Y12S
mwKuE2xIOoB8Q76forB9urHWK3wRnEAFhF7kg/B8FApj4q1ygPr6XEbxqfUCyDDM
gYBBDc8noq7WfYeM818KrTCwckR0PsYzBVkrZyNw/kSevdivqVMQxWEQz81X/EWd
WsV1oZbtPq0QRklf4X6eH7Ez/FXMEpG61m2uc1wnKWJm8XbyQkRAuqxj7+04+dQn
7LvgPPtC+OaOtUoMr9UTYs8ZS2U9cRwgk+1fZ2r1+t9ZDDhTKnd7YINnAS1rtN0Y
04cCRqj4OTgauLq5MoXUCDS/tw8txTR44dSmkPeL313auB/Nwuj93jOkguvycC47
vcU0c5nIcFBG8jL+XaNZjXfV+NGIm/JhX1xUaxj/axjznQnqdXU/+oMnWzgSgvt7
YbYdudIgNeb66AYqkLiHT1PbEwGtI50/o4dh9vsDhafaBIC7NJ5EBz2NNYOMtsgl
VZo4gitckIKnC3HuLsWsizyBnSJOeUUOOui+2keUkpzyEvi45Yq5hiVAjRlBP8CK
L770w+hRirpZifoZQNnkP7HdbGbp+j6Ywsol4tO2h8xCJze5AUq8L/0Sx0mczhwI
ypihKzH1Hw1wwgtOYzrKb7AFTdoGIVnahYln61DJlk/EMjUDp5re25zgb5CMP4PF
SFG/QVQ3N6u7T1K5nzOeUWNdqKbXfNq7FGxkPG3j7zzGigKWSkUeUmb7hBqRRCCb
sTqMXh0pCJRZnEnnzjLHUX/CJd7hReDO0u1fIgAxfnlQf9BT369443wV5rcUecEq
gHQSej4iwGSBoZS8zFlZ28AeNBIpLV+5PRbTs4l2E89Pk8ggEKn/8jyD3y7aRDtm
VU+od6lTLrTdsyb6LakK7mbt1P1GTzBJnkfAQuaOLaYA8/Hdb9hhWcQctGhzm4LG
zIo5UCcnqFqgnPJdEVLUfICmrNgGp9BsY4xXPfnC9r2Nr9gd+tJhOUfG0Fkkup26
gMlS33vcE8K1Os21llUoWfgxEYT7mJ7caZQpth2L8ER70j9hkW69K3LLsme7UwSK
Is21QQH0LgOjpEHmQEbLk/fdZEV/ZrFl5skS/iT49zu0bhcIwIstyV6An545dfqk
62wMfEnmFOVveyR9xjC5S+zsdykV8Dao99hN/rTkYB8SAxG6PqlLtDKrxOkC/P/6
ADyu5+SIkLDvx9JbRDzTn7tA3uDZhNiwor1f2h/1eNuUZ2VKWGNygIfs2616flRa
zFebwyQ3wqsbeYnaNNawo0z/zJct3VjJ3bNMZy324KUfKr2SqrMZVGDjWklwBHKJ
CwsPypC/1ebvKxkdybjwp4NI3/3wBciZV175Za+t8JbS2GAwJ2GfOg+cbR9oyBXj
ouBBJhgEu99eHYZ6lP5gip1z1aZCNC4g2AG6ZU/UEtZ4rxW8hoOBGxYbS8tCbcYE
oajuXniNUhbk2PeY8tevljevS037oCWTDixCoucd4OXSO+QbBYCKuE4TOMXdVrCJ
dvqYe8m6GgeOL5EQq2AoVP4otPl5Waqrgwq0HwNoYsajVLWs7R7jhMRbAW5V4mFz
IiWANE3tv782ONFQgChtFk6HvR2nQXbL41dKuOt47EhibsiPQD4WEzQid9G4OjVB
LhhjfzILt5qal60LVsIuCVnayQWDlZbs4GPpdjpk1PLPa0IgX3BtwrI2WOc7bPB/
HRKf+9c3G1pdwv8FwqeCrOR9VoS7r/B74ViTtJYq4U8hOvDiWeX8GGZgVMvuQ8de
OoHwPo4W9VEyRasaqORB74T7s5Zky4Ue+3sJIvwUtXOVdzqX54Dl5Sb9YN/TpGEh
GfjhLFNax66BHO3oo6xldi3uZFCLMOUh1MnVtFBPze3E7nd2hS0dNF7/Tq/ajfvU
fhqsxvBMAa3Jrl2A5jfT+z0J5/z5JmItW/GfjpgFWTFQojDG7FG3wSLA9wU6nc4Z
n5LVlcdASLrpQYpNrHA+WbM8kF5sOlgAfwkSsvj5OD7BQazhEPfdJ18HRIhAAbF4
h4aX0M5n1/TBYKu88alFwqe/IyqxCLuUkB437DT1YTm2H60OMgHjuHpeGd53uUON
MnJ6rULFPafNkmsgv/snIasqxstNqxH9gA9Tr8EBVyBtHxo1JTLDN3FUqWi96Ym0
Osw505ii9OahM/Rggxsif5XzRq3EQsS18gP2XLQF8+S6JCXlT20tGf0NkfDORmmo
qtC2DtLVyHKU3oeMfnZH+RulO3rnsEsIb2k+lvB9Y6v8gqunNyqfH3+njWSo6meU
BXFNsWft7AG0pIGuIofXRKggvcqH/Vr7Rc0LJMAiu8wsLPYnoEdlgrCNX4sa13wb
Vr36T0w3o5dwyd+UnRzXYKY5nM/qQCsTFb42/rxTHorRlRAWc0p4uSno27eeKaaj
WTo+LCCRtLwSEdGB33ZQM+iEj4FfUg0OvUZDEmSaxDsA62U9y4fNHzEGmTHR0u1f
ox7kd8Lv9MUJ7+HzuRVxjjvOOS4BSbZ7lBWyPiFIv8fD7ZSR1aXlK0zuzQP76Vea
y6RQ8fzd7DGLGqhLiinoLRZAMpozJYajjunYPZShViAK2k3qveKa2ZLZXa2LFetI
KTtARhjKnYouvz8jjLMVXPJzKlSVVwAJ50t2e/VIDFTj9bTL28GozC+ie2TG/3rW
1FM3Ye7pg61gYJcAch3PQLwCEs5YGKXa43ES99mDtiX1OV4ZBMOGuFMmXL5pd+Xp
uZ76seE6nElhsvoyF84/dHbk98TXSyET+1EHkl7y3jyJbYXfOYaQLYZqqKg+nwMd
k2m8ImYaArdWj3g9Vdx+XCC7fEH1twU8xq1haVpm4P1FShB2TzuNI5A4w9JYZS3Z
cEQ37vWEqSG0kskLVJtoXS0Y/XxBIlYk0A2eQ0hAD5Vu/iA3hvHAKfL+UJMmSNSH
1TXuqxKnqOTAi+1yIWUNnp16BI8KynLpWFKYhB9iDapehDjxpR+CvB9n74SPBfeL
N4eiDf1RKpNSlcRj+xBO19dsTy0QZveQN/hwj0iV174Itb7Vma7r3pn9dTmIhoFr
QaDjc4kAFhgbMv9R5CB8eTZ8eU/9cYyeOXm/ijU+twPJ1/xO/QDBQUPemQVEHwei
+ZM0zh8wULRBEh1/NEzhvluVH3BjJ+TR41OZ/hjVsbPsu9ndaK2q/dw4sYWl9jqu
bqq3YsS9UlWN9Ggc/DIia6Pr3uECpJhtRVSJHOX1lXKUb7nL2Hf+1/ttFDJg3eHS
CYv29yEJPuPy5hu4Od8kxx48zTeYTucdnOIFKDv0kHY0Pq2Efje8Kv9SqVSyZnhI
S7UakpVjV4e7+lfZVwgXYOox1FKf+ixdkE9Z6Hsf15ptERc7Z0t703VYSq7nS1LP
5aEoQFaDm06Uyx/YKUFBt8GSRQuesUNjouGMBrjcxweNOBnRbZo7Y+S1J/74Vry8
ZfTRT0UppTPOVY9yqnx6J6URXUK9lf1XSCKmmR3gaHh33vpzLxyv/7wnkpRhdEou
Gh5gjV7QR7/WQdumjQj444FDnucJBGtDCeziIcbI++qYipdIjtAu2j0/myA+OldH
rNt3NBiflBr0THf8/FsEwX367jLq9Ajkn/nIWJyJOuXTpu4eGNjtPWVZBoeFTIYA
kHT9HEfm6/YrhfK04o0q+U+sdu39exV2gwATsDw/yBzgXFOFd3YkGhnodm//3rS4
eWfjfFh3n0z4P00YECURVOG2HsmEbmZ6PMq/BQNklZ6+OSa3XMuRDdLciOfyScl9
tgoqGtlBjpIRFCSF9rlmYF+JMPjDmHZWG+d/E5Tf3/6LuqYVhqcvNIB8spidRH58
EWMe3vMVydNFliL5yk+U+0fMFhTHj6vsCFblEvCSXAz3eAIADxp8mHi+1Z0l6nOx
P7NYWuBNIBzi0TDSNEn+wZqh63IIQmYqNTVEQruJ2YYXS7q/CQR/+pk3oreNu1EI
04I2nFp7BPSoUy69QT1rMayVnn/XOOAbTlEyHiZhEhkB/EV9GDxESUxHMEyu0qAK
MxJsUlv/CraWOTmBziTIDB6x1kiu3DAaazsIUq1bEgRMnUeCEr8ultm7CNOigpXO
ewszGidigq6+9GLAg7wWR46Sdi07VeV+vdhX9XgnAyzSgUl0M4v7fHuBaO+i3KOc
kJJxfqr6Z4rr6IFg2SqbW+fU36M2QF3lH326Aa/uABM1deok9DtXlUZZ4mlbxOI0
TI/3/kfyrERFjaLHurN16caAwWTgx2ymN3JhJe7rrXOnoMjuinKS5zDSVwJ5I2aU
7aAnajVlHJMtdJ+orSkQSHn4cv2J9VxhEeFci/WSnWbv/8AOKYCbD7ijfuT9Ci8p
Xlv8zgsZp+QQGOG1ihplrgb92+q8yMEsav6Gka3TrzhJeSMhnXN2yi7EXqjL0mCu
TbFbWDA5xlQSgv+RjJCPQZ3F9meZerd2gUEWsAoQ7Eb/FfbiHTe6hU/gxYM5PDMr
GvMSQOFYf9drthhHzXCGwCFlr8E6KpyfelyH9DxTVheAYpLJZdWIT/b/+qq26Mm8
RlORJ5vXIvARocfyd/jLeiHpl2bHzLKx+P/LRu9Lrt090g487K0tNHrWznwXnKdp
5P3zoxFxot+qD/VcORVJyJbgw4t95C6Pfk4NyHkwrZn2sJaE6jQqGKnXiCTXvxW1
dZiLxr6zSIxPAq5e4YBxqmbQ98Qkgt4aS7lDUi6fg0Va4uLNMEc3tIZv+sQSZNeQ
Gz0WFkzWohcCk0NgOKr4SxfdJzmQnHKLXpmEOtPl9yyR6X8PKDjACJfeTtNzdTF4
f3OPpeEQ/PNQDjmHqLHC7BlSDR98l7mkYiKEpVdE/HQ+cuCvyr0AAmMGBStX8TeR
1bF5puwJmKGAyQn37nFJmnbUtbqSunQl2yUsVvJUttD3jgmz8hiw+lP86039i4Dw
votrUqu+UzZWm9g8BrHqhX7FTb70b8dNi5WV9V1OKUVVPCuYLBNUd6mlmPynfJRt
ObUlXeyBskibExzofqhgqoNmBib6BSJXfgRWmgn+F8lRKCvfgbdzP3Cs8k0K2VTg
wAnJAhRVh/FiWKH2AQTm9hU6bzN9tcUy7s6QclGAneKo7aYKTfDSR3Pv8hhgYo8P
b2kebaDfszRdYWSO7kg6N6gZpZGqqxu/l+5fqU57MIRx1FqGGPWLccSzvz+tsIj2
jCsVvWEJe1TNoy9qbGlk10eOSw2iP3XL0Ik8zQx0vlDRaST4UnYbqIimuR5unL/w
lhgsBOySuo2AEE4jgHFCN7P2OVWu1e+AJHXGKC8E9xpB/MQ3w6mKGSgaoAh3Ig5Z
BGvs0pZBhzuve77McpzHl9Pzxs419U/e1sPWbeNxfoIx5aIty0ez+ec1yNENaYN5
3Ae5Ku/6zg7lO54Fo4Q01oGlJYYFGgzSHFRGW7TGBFa3yWUiEsWstQRrNDGe7bsY
XqWC//Vs/dPwND7mnIJhV7JYiEFQveot3CgBR/UzxW5TqyjYGXPjC4UnACUc4Qru
P8moiodJNJs34iI17Nc80c+S67o57jr70+BpDEXa7lzf1OKbuuQb8AVLVrj16MFg
FjXOWmqeog0mzhg6OXczmIWNEpdGMaxwGrvUXYxIYCmbslpsac7CekxQLw0yNc0d
NxdmQc/m9HeUXqeuHOSizgVxN/LuzDq5Ws7Hxa3GRX7IXQ6Vpv5uhs1zuaUnMDZd
zC5tQ0qVN7AH684ArjQEwp+OKk3R2b0Z3bB03+T4lzFroDVy8UIfq36eLxLAUGNE
UEn+9H4/qoQNZE8EjmWi+BG/wT9ZU7+4uAQH4UVA64iw6v36kpvA62KWXimfddTB
yUoTsjyEbWx699716VgTmJMIyM7bJG1RHqG3tukZ7X4vsuKLEcll3mclefWsS57/
avRJhtDPFU6VMR1d51GZGVci0Jwesc4GI0cg6p80TDbUKFmVgIfU43z/TFQVp0W/
LZzxt4uuy1PUC6EOxW9AOrbK+nv4wN/JN940DEP7y78sa2S5XHacymhP/rvejeH7
bHIxKKbsf6LtpvEqoJpgbL9igh7srw5lIj8t5o7geRS8Zm8n9AM/E1C68yhl4SyN
5tYpZpSlOewYmq0Alsw/XSfrrlEyEndwt2mlWcl+bqpB6K2flBWz8M01aJCVZAZE
2W5huJmAbZ/OVSnEfcSMwj2H71T7gOwfLb87v0db3eoQBhUFsTgTupTgkV+oAXmk
tE7y4g6v8owtX5VBqcA+p3d1n+TNUzGcm1vw7kMq1+Fymx2O0Xx7IZN8CR7JRrtt
mfppY5aFiBw6RGDlkTa2noKgCp6aP3RIdeDnv/HCZQGiNQh/Z2/GQ2+/yYO7RWQL
hsULVWhBkfOl+f3MR7ann1+XUwLOq7qLo5vOd+YogEJvN+plAahMKq8IH3Z/Yut2
vMmzIbXZljK5HGmtt6rhYW2j9+AUzCCJgsO1Ds5ueYzQRW3/sTpIIMknOPJi345P
AATpLr5nzmV9lHHPHNgQ7KFywwTrszRCTxqXmvHUeMsNGQFAnVrGUziCN9SEG3mV
FlJ3XMQGjcaWrJitDsDt/KOGMnxtzsnagf75LiFGaagXV6oRsE7/1kK0xtHt7DSA
JfWPV1bAGGB8X7SzQ1ZJvKQvzTqFOZCKJ58J0OylhMGergCMg0eP/ujnsfVF7mZQ
a4PCm4G+rxGEaJqoMXN4BAcOXyLNBUakxFxQ08RxUfLfyrhVcDckYwFiSI+ylAXr
gMZ+3Pzw1QQlG4+SsjU1LNiYMSt3TfNEOxcUAZIL8Qx0jJQ+iTGJ9V1wq0w3frtl
m4HoR5pXQj8nzGFUTsvUJGfgcgHZFwGYWMq+2YavVxdoRJvttz5Qn6FA46r0THkx
O4MNrv8mqPEDZIawK5qCfpTal1JtKCajWcFoMpakvM2pW2JyjeN1Hw1c41UTTk2l
p76RXt3HZTOJxAjWNA9oUp+s08Ea9DA2yrxsocTXVQtg84joIj2WXm7wi5aIiW+h
eK+DHMC/Z10pcfziPsTxMnLtA3znbvjvLJWjv6U+ZCx0XASd9/wVclLcQ0tvhrvf
hkwJF/APbfMs1ZMiS8c/YV5dPZB/MDiCQVeYEwT9kOmLbIgQJlGGDoi1PvtEn7VB
QyYabAlOzDDRhGBxlSUzm1EKN9VaUJAygeqb8cORMpeUzDBZ04vKwNLIKicjvu9j
KeR0cOFaDYg33UQPIhBBFo2QfgyoHKLKS9EI9/KVqyeuuQkzG+mYjk0Rg3MUsu5O
rthJW/IQ20wPFT9q6PhNAd868tIhvNcgf0T88IJswwLjaWfm5BJ3w7A6l4Y5tRSp
nS2bHrNAA38ZQ++GoKe7X2jr7Bk8IQudMezJ3CuZU/T9/7uGPmZ2YkLoTwP5n8ok
jJhlCWPFgwC4QKidkWZEGaTQDys0pVhpwb9NwHUp1Z/KGs5sWnR52jHlyGE2bJjH
BVmz7Tktiwn1h+0EqOI+T34lF6I9FH3+q3Nb7vFmXoqbUHm92VnTYATf9PyxQ9ZJ
b141aXNa6AF/yOJcrIj6kC8U3LFDRyzSSnd2rsAM8Xih1rHV55Rs9wFmIu+sy9pA
BWkyOGF0nDibP9J0omVHFsRE0Cf1t+cUSBLLWhFugiu+lViPuAHHGGuK5xUtv6HE
4WgDsXYdMMCBlekLYaqGNYizLu6ZP/kLVUBFuF46IEJnE5tM4b/SUp0YPTVDRsNJ
OSewRLag9V/QTIe3Y2ZX7kE4OAxKOa7IYFyAej/n+Y2BfoUerUTuMzHVPLgTbieT
/mWpO4H5VzSvBz4JIx/+FUXBPRn0fc0cKS7yLzPLRr/GJvMNJdvlJnAww27LF4mP
smxQnuwim3D9dRvrVVitCjb4o1vbNGLquMuXsf8jyF7xZ3PTQX/x4nWPeQqfhL2+
NYxXA16HDrpLpuifZc+6PIPh6mku8Rg4rUyFUCsPKf8zZmv7f/u7dAa+oxNvgBVe
E0A6qoMX+jUL4ENJodLvuWAqvHI75r0MyyH0SCEturSIa43khVIY0qFuy+Lv1Bwo
FWC7VX2R/r/8cyxo5tddzgap6eqcbtL+G6TVfzUJdICFyVBMzEYOMxNbjhcHx2MC
zSu54oqeM9rGS1mDlgVJNbEUlIEJiIGQnjmk4rb+VAW6vooW1OT4SiUkVDxPbw7Y
doTuFwbyjQ2s+jp0T2ehYJlk/pDM/u8QBTc16DwYyzBp+s854d4CV3zXnxX8bLIN
kxnnPr/crgI4kbHST0p9lwG+FBU2El4WugMmGiZL5sTP9Yq4HayMXDp62Sefiwxg
Q6iB67QXR+a22rp2dfw3jcD8Kh+TvXdY4uMK5t25EGeEDR/hypVAFTt6fXCZ8bxL
WgBcJ1tVO4NG+x8+jzcTQWHZjNmcU/1dhH2zVcZrlXpIJ+oORjFnexBc+szKN4vA
JbIxtlRAefrXS3KxYY4JkzVYmUceu7D8R9Ho5DLdtO+16NtGg6K9LBQBefsmw8iC
YvcP5EVvDNgKPwiwKAIeV0k7XGRZzkseK5scQ4hL+nuhLr56tSe9gg9LWSE5ah2R
GqJ18SoWNPEASyHxVO2r5RqAOwnGbKyw/ZsX0L80ntkBRN5LTdN4wWj/F5cNStyv
x8Gd3yC69qTTnsz5mt075GIOKsv4gFqBXna/ZV35XCp57uFBjzFJILHJghJMTZM3
tK6vSwIDZmQ6SDPBIcTjdrFuPL2p2ot2eho9k70Kay/uYVp1SrzLUdqVypgmbW6o
JxbwE5ifMBBRfOhQc+u3KSxi4YPt/jZwkspFvMHZnnoOmsS5dBaTHkq9XVVXKw4/
/QO9+3N2l4vxSjKpLB7zV2NGP911hnaaoHiMX3IpvlGQhVUf9sawkqj3BmIe3YpH
L7CGKOVnBGWCV56Q3v8nJCIaX5qpJsjN/Sszw474IEM0l8OBiT2UkA1qVlCjTiCn
6CTYpnvKGf1n6zZXyq4n2KS3SCNy8x9dz+O1Y+XzYlrJImcpzUtY79UYBsOhKJ7/
FEfmJ/eCOBBxobghhYiSqhEU/92gjOIfbaK2Qc+pg02CAqVqDHNaUipiEvtS+jf9
S5TKfYEBBXGWu3qwPaGHVfkL/lWWXOc/NJMPTwc2vYwIsPPbkBEAnQ6rG/Ojdk29
tax8mKpsuTAyDMwVSuAZ4+mg436fUJBlcmlFYT/eotURvIK8FyACPokMzpFyiUkP
YlNSlGI+n6U59dfrxXN1CwgUJUmYD3cHZXa4ifIYt1h/+2kuJV2HMzeRODs6Mn07
Y4LQ9Z4RTGPXZvA0uoRyXboYQw1YmOkfIRfj7dHlqCxu/fcZA8cSuajRTZBCzv6R
ZdR04hVZw0kO17hceIIzd4c3o7529S/Wrjcp1lAqllZlNM/Y+8iiaTlOtUQXNI3E
H1BzoRt9Gt4oOjoLHjsl1ERLudXcSLhWWDTn4/ZskxeuUX+AXn73wH3Ro/IiTSeG
o3MpPQlc520dinLAjkM0paUvfBIS4R1ZgAN5c9CktCXdZ2ZZmvA9EpBvfHS2qqFV
u5dksr4ABJQ8ey0f8H/JXmGmvL71QvrodFJrjv6gzR/4xfC7/F/auVgOCuUEIHmk
eyRaZXTiZlEVb2wf6W1HVfckqFmIRPHGBmE01lUbCITAX7alTOEqnwPqHuRyIBKF
8h6MbNYH2oHKID0RZsuv9SI6hFpOzuOvPQQyG5B/0gZM5BZ6xR0Rvzq3o1kHreYk
ARVRtQUCAvRQA0+2Z0svZjGfvqV1dVKOWDlZhtRRtL3TYRjhVNtZKSoCnyoYBzzm
KJGM8jHKzYeaSBqSvA+lg/+Lyd6+3mLVxgUeexM1JcwxvYpcz0BsZdN/sb6lhjSf
c8gfxmxzCJX0WyN2i2miC7ZEtfeFIusE5CBwXLMiQgDNMVrL5DpgvrlXkFwRRPiH
+bZL92F+T7mYW2cHp+vF0QgKFl/zjcaPcvL8HBOyWxM5ICxF+99zdaUTkyU3Bknh
PBFEvIkl4e+M40LGkd7sTipdi1zrAUeCteapxPHleh+Og8cGiU6cOXgIDT8xqZB1
FYOPHkks2zd1EynkWV0jd//0gMnZLJZarcYwJoc7lEFbfn4fq3dEIjBqvAKmKNZx
vAuPRj5CHlX5L8u1iFTK15DlRX80Y/Apcy5CP07XcL+vQ/t2+bCBSziPGLLBrimV
mWBAzw0wK8fAsVfH5wIk8vSLT7++cT8ExTvEoLzk29GeFd4Xzj7jbgHAF7gDR3/M
dfqxFSYux5hvNiRP/KJX/6Nwkub0DkAYzvY9hcHgat6qeBM4F01F7bw/FcSQz5JF
nqgWccSGJM+aaBVm8+XTxTaPIYvXb6hO27owJFKtCPfoViPGiVjoaXPd3PvxVCZx
zN0UToteIfh+b0mFltm0FcVrs9P18O82wiqD4idjZH2nlhed28sggyVOoAdTB5WR
07aYbT1YdzPHw3xl0riJh3Tu2u7kDq6f6Bg6wx4JXchZsZg10bn1HCGWAN78ak5P
8oo2fXeJjAW+wN+HUlGoHhRUVQWTul8kSDNLsPMYo5z05NRKHgVr8mPHJh+k+YRc
GLm6+WPYTFm4GnsRkL5scZ2HjIfj9avQeRqtTkU0VvqHJtvJx3FeWrd1RlgSZ9lV
7Fe8hCtiEa/tY77NtdVeJDQUc3LdYC5A1uUrhyaKWZcXvnQcFyZL9oMwIp8Qbijc
5dOghLk1CGlO6lHA2XEqBS3nv6MzzMa3IeaY0VG+Op7o4wGmGM6fjwYUmn1qrDWB
pMObUCJEu/qKwDo8DkJdYj7Di4HtpUGGt46XJ+ThJrjSnrOCKMeZY4JFXSEoYWK2
W6YwDoh9ST0O8jzO49Nf0a6isnZUROk69JIQDpcX0O33Qh3x8P+K9cSMzOhi1Kdf
QbWZtCiYmjDdHy8cGvnfFcMwaCfGh4a+T1w12WXdq5QKsjaWQ8NE2htfPpDE5xzF
1gelPsJZN88lkgIpteCMhL8U914ZR05+rF6/B/3FJkLaQoP9qkoz3jh5sIyB6BAY
uj2QhdLwf8gtCMqkyFAvTY5ohjWIqZofyt+ZrTa+H1ZjdMBhqJ+qyUJ2wLY+OhD+
MYdEr1YpxMj+At7KodOYl/V+8Nvt8nHIFrdGrTk7yLj79rBxO69Hsv5x7KJ8AcAb
i8iNXDzRZjsV33n71k02K5AKEw8XowGNQQXguIvmM6PjQQrjKTli3a3bzEYiIbUi
SmqpVYhckR5uSmushL7LVFKusfVEoF1ZKscV6652Rn0jozh8zvGJ5VxcbwTUzUWc
1WMuMJ3QXmjpvyFYEn6rZ0vp5N25lHwJk6WJCWcR4WVR7Byadkawhb8Utm9MYzrd
GNGPvnahBex2ef/8AwtJzJaDrbsfj7byI/+UoS2IQfKwSaQ+qcEx2Pt/TrNlclOa
vl/zwMqqqof1O7b384nbpfv2hCCG/clWZepniFVpNUBD+O0uQsKpPDcMaNoiO2MB
Iec/QZegFqO/13XVySTLola3dFtS2U6Xcsm7Mhg1Ah4F/7oIs6GCBVdCF0gsFmfY
FaXB7Jr5OlTicN+QQeIZybf6cqQDQKG+HyrNJgYz5lJ+LMQtxazBDQIx2o9In/xE
hJLe4oJqR07hRuXByScNKt2wY3mrY9gCS15A4euYsxHzUEnWXM1Zjk/ObgmrSACb
6uwC1aJgH0LK1bjtjf7rR772ZHGI065640OmtuWvTOoslyWD+ABFPQjJ2qrQYI6D
XXhBAg/HHR7lRlzzd3No+kLF8NkTF8WU4kLLTg2xi/TWSrB98TyJ9btDmVoPdnr/
378cqT9ZoF0mFvi1MWMvB8W36w7Tei3IIVljcQ6Rqmxd3eS2odlZuTkfzJiFTBmo
XKn89Tcy9Z2iui85rXK6ood3HFFzWspD3+ZuBTtSWtgUbiABpZNIWjiEkZa8UJuH
uF0mEZ/owrU1bVJtLwKq98HXBPQBD5+8ckiP8Ccgczr9raNKS+wffCsXxn2peVuI
vFGwpIl6xohd0BoUTL+OpE3DpUEjwIt8ly+ShXPawn/eYpJFhEYwLRaF+lQwpfsn
B+cRVBEGDxkhYXVepYWibm3yMwSK8zV415nhArSjevqYV6ntD2vTsqHb9RhmIvHz
UDpn6zE4ZqfA8b4y+eqdtVCfpsDw0BsG4JFpd66/26u/YoF1DlpQ+Mcnw01ceEhe
0ORZuGsFUWQHgFW2vxam/ITslNdDbYyWMUQ+EbGiqbIiJkxXiuLovB4hqlQzOiT1
RZgyPtp7BpsBsJFQ97co1fEdD1yRpz9qSVXxOVU9MgCpwpZOlekQIRXnzE02vxa0
kI/ZxyyeQIcJ43LIal26OkfYTQrczP5IQKg8x6pNZ53lDrmTxvGn6IQ5w6nuy9Gz
htt+FMSNDoINWbl/of/i3qgiTl4IvkFIRTUJE4wEh+VOVyl+1CXmzt4CT2Whxl0Z
pSgOf8X4oOYDQyv/BDRssbZqdOONwANE5b0y87wOYBANHr2J+B6qtMyplzG51y/N
yiYGlNdRVCSLGVmgffz/ELp197oon5Y4QCZmxQ8Qda3W/8zM1iudnzdMkIwBrPxG
nIKT1yz33JzkcwDLhmWJIh7Cv6XMjIZ1Avs6TQQyAfmBsVRTDC25+Bb+A90pPVFW
rC1dcCXIix1qq7rDn8cf2rutdYReUUjcGftHYiEYea7pncg8zyL6xicOKq6R6hxz
KmzALZd5a0bwjeBPFsNOx08nyannkoP6KM4jH2LNqD0oNclLMZyk6iEzHeaaNsiY
x+7m35CVIGxtmCWF1hRyaknpLwEX6J8IKFu14ovNehaZWHGA4UtP1EwfrBzSMk61
M6fRboWv5w2TNrVtWadd2f6v1ywhj8JcPkYiC4LK+l6NNijmS7oXM/jZlbXynF1D
aND+vo+7GUWEGe0PiEV5IPZW2fJku1HXQkkgCLaZGtUXAEQwKvoCY2blEAHNsWTm
XpZMe9DErJsuytOcldryvCC8d/Gyr2PbA/FZmhAt8CBqMT5M0pWE0dHc5hmAa2Jk
rOgwKT9wk5gX6IrTLwbZjTwzk0ML6IwLaVVFbtOUICTmHFWpqnucz1HVUhoOoStP
uPe9fE6T01GAKYE6o3Gmv2GOYdmqJijWl0ElpLIeD9jtrUdKHrtdqMDn9brsLegu
Z4mL7HA98Dhx1y4/oicKrCOijloEO5hd7KkSn7lvS2Y3AAwkMI/FQdSOxyUGOvBY
FbMcqKClV6tr5uxllxKgiw9tsB+HfkSDro4Rt6+fzhr7PyjjdEQ9mFZRGc9iYSiX
/01ba4Mn37Krby7nSd2dypHtr7nL3mn99mSotzFui5kdvi0w4OXYLXJBCUHiFA0H
1wHL/xi0xKUsSNWJNNkTm79jKiK1Q4Xhr82yz3QohaBGjUx+BWkbgRz5e1LOVDjI
3yd0K3SLTitV1i86efUEZlTtkLnAV02H2KlpbZ6gCxXvKm0B/K/AUzG61/Q1c2PU
GbghMzYH9dlLKsLfFzErx4Evg+3iuSkVfSx269qRIP+jrwn6sQJj1GaQziwTwgAX
cEeYkCfUhqkco7zP/e9eZyGnyXTtk3CjQUcSck348P040vBb0WhBsiDAVipmH4w2
nzNI8booJ41Y14Lk9yyi8ZC3hhp/Fmpz+yJSZjcs9TBU9JEHeTVogcdDD1TABNsS
AyQK1WBl7n90z1n9rIsSLv22ujuitE/SJKuqYWXyxZVS5Or9+jP1OhG4O8ckHw1z
DPJuJa/MeipRwjxrrASxMEyPtqRH633phhLysYXMMw6mFgfKfzE1D2WYNOLWtRCh
Gox/AA5BLa/wzI2ALz4cUoE6WWf5QMYs+2BDM9xjLysT6F6pds4oDHzP/jJd5xAs
vFyRJJizJfm960GcX+SRM13kU8SNq3STi2Fp9ENjZ9+CCfnVHscRdF30Xy75cnt+
D0gntL6101aCP/JhutkOZdKzMNHcGImMg1QF+u1N6h9t4tfrVSIu8vxbcIBpaOOW
qd6I8m8D5kPocMknARv+21c5vjZ5LFXNP+BEG1IhbjR4PPrzz/mz0tJl/h2uokoy
Yh1I8mEcwgqarff2EWXJpXB1TllkT4D/6VXHZOyixs/IXX9fARmdo/TsLqIUcZ2O
pH+QHrUzZv2Kqk2XzrQhu4o39NOEiqfXP32OTPayAQeltPZ/a+xWglYrsBFegxLp
rrNNJNUHI0Irm4Vp4ryUm8yUUnECJEIydE2ls1mjZDkpwASCMB1RL8SU4hXEcksQ
lN+iEIHQzT9oWSLZQ34wYRv/I9UYLifOQugH7rVtOg6+IxRWIPw1YjTP3YaBiKcJ
XejiAUqKNFb/h3HEzNF9Cmia61t8ICOPjseLvxint6fTh9f9AHy0kJuIL/Zbpiuu
EukjYFtzgrIOrYI1HwmvLMXTDssYKBcXRHwmSTK655qSIb6//N3654PiV7VFEkRG
kaV9y0B06ko3mRiah4yHERYX+KAvIKvVSD5KTtO90N+X9RbsWHNVNN/jURymLcOp
nXvjdFW6JCW6a4X9urLBIBA5yRHhQxiGyzrcQqxnwH+SSZ+QQ1ehA9xxc0dCByTs
Ri1pLCKvnb5BwYCwZY5ArnlQINV7h30uKGYIYXPW6RQXuFh7TKz9SW3B3fYaSpJq
lEtyyTPdDTLqTU9vhkbNGzRDf6luBJDSRjoNJ1kFo2QzPOuceU8wVIdcYrDcXpHO
WZBZac9yh1ixi9wnamvACony1pKABfFAb7CzuMkvCWe5YA1oLHv0BkeN+WAUe2he
0QaPs8EtMyWFl03voKIvx521fwkoxis1lHV61FdU3ylMDaf3w4sNAKEY+B53rNok
Jp0Yg7F9UkAoUAAWWkqon5GnQ/9awnIiqH4Gljk0TKZwt/88xG5zQeeaHPmx6+Cz
Oi+hko8HmjEkqbP3ERRS01BTwbFN72lgY410WkPcPTwCzrH+4BltXwYP4MFTMH6E
LGtq/+ICPVXHOXpqOjZ7IeDr4bDu3A6CALk+2HOz2N3fj+p1uW2Rq7XVnMmEHzUU
Fa44v3Jx+GRlPmvS3yjJjpNAZHukQBeiBleataYDyXkWfVTMYn4V8NqZtRsTsoPT
yFscGieV86/IJjwWnnYC+wHBwX9cuqnjEyx0cryDJPp9AAe26QDBl7+UjSUYRwop
XHR+jcEvBRhbOuBMh2wGQDC9FtfxVoT77EX1cXDp+PCqdz3stgDMy8Xlp3Pd9HeG
7v23JgqRSBT+qVvIpN/9HfezRG+aVGjQySti0nPXw1cnlD5/E8LzEG9ujY+RSbKN
/o/pVSXA5y6vMzspXcuFzdzLCFw4yFIW4g5bD8QApxJf2H0n5YzT8DW6vPtBlu3L
BpPU9tmGo9n9X4eOtoQOH0JdX9NZSCXv+WY8F0E36YsS3VufAWAvWFsvxzxnPvpv
MZMIQEYhwzHwTvb6lOVWfosqXdVykarSz7RlkH8xolmuVDMhpuu403NQrOiZkDtl
tJtSpT4jx1UtCmLsX2qfJRr0zVG1/8NW5h+n5MOIb01SK/WxehTeeFIGqMXsbyYp
OK+TluJmuszTCtFkGUZfgiw1dy6dfaxPHi6/r8JgN6OyUoJhnwc4gRZ5Wlh0k4dM
X5URSZhlvXIHsPVn40UMza6jCsTISE7g4w4D8wxWptE+akZYawKBzoVNolIcIPZB
qqjcACSpCGBSoNBXM1ZqLrZAlDw4PVpbeYsweujIvAXwZrtWOwG46pDaAOr2597z
KOpBCLy4MD1QtC1Iflbj1rdIoSAud86+uTWpzvbcKoD7+zahzX0osqibxl4Pa3LK
I63akAT1cX4VU0B5Yk/Vc2UxXIRUwBIu8TQbjjyVMM0qsaFhFS/xwiwf1Qs2/KJb
PIf3HyaV/RUeTMJh38iHl//Aq0Xp9LOe4ITj0RsWt/414xknzC1Z6FVwuebq2ikr
p2pg7UBD0IXaaMouEeVnNxvPE8HGYoWD4pL+r5/AyxGoqoHyrt8Wa4T0T+yhEJz6
rD72vyUE6yLfDav32lPA/Tkpauxty/sEoDWkGhIZnu77aTBqC7gdofFmYylrvnHp
/Yeuu3I8gV5S+LSTg2GIY7qHx5HsmBjUn5NJ4sHZApx/e3RsWjvBTtYfFjNyFJ8c
kgdE2uVlydY1X9bCrFvsu49d0F0FFY6tISR9GsvVIgjElBv3SHXbMy7exoM4hi+N
aOZ7VbYrJto9COrJcXKPRSB3FcjElKENdKQ901UlZFa4u6WrsVVkRpTRbWVTQswE
KWPVy0itxhMEh1fRu5Yol+vIZBntmmlZDfn87WxfPGe3uKQqRasxynyqtAgVucZp
YJ3v+K8hOlit7cni64zo/n2BwcxaH+dw+Lpb66PqdsbunEm8ENCBBn6KYq+IkuSh
B6PLBie1mv5fgEUDhQv9x5Ilow7BfVTfaFi1+QvAM8N20a6bj7ZmoxMf/a5xqR0D
49wxRbEnsw+DmSIr9jLhOfasfDvWgEK0aLKPg5io3AYa86ed6hPT+9gbrlAc9OJO
53a+khMe2LfzcVDKKTykEXB7OtXSKr4UmcjSd2RzUhAT912A36MtuQ+hbqnO2iIr
eOE5aKh8381lakpQtRjG7GeGL5OS82mOh7XJ/9QwTzTqk+mcmH/3k9zTVzuuRfLP
8WBgNeNpcVVBLXBnYIPFr4TTkX+m7nXWKkE9J2rDm4tOUNyOhKlM737SBALuX3LO
cYyb6hOfQ8qodr2cSVazV7aEE/ImfxM/r8ZVNNLc4XepraYTK/vXzBNhW0Bxzv4x
/SINy/CxQVd3uH5CpSIjzs5b/0DnwKa6kwCvHnpjsgOQXAIK5Ebf+zdBP71/QX6X
A7Zl8kmiyCeEdn9vTfdDxf9kexHnWKoJra9yaw/i5JpKHBfEMGYswZXz+fRZBQed
VU2eo8cc98gqspdM8qAPTC1fssoOCI/9NkufAPwRyM7Ie5GR0d4EinOuJ4fqUhZb
Jc1NuvYFXNmU3ZhgWv95MPtj4VtUpXzaZCs91FCaULFMsxe1NAEG4yEzJIuxF8AF
yMuXMaYLYNL3ySyEiBBLntpZVI2zWnSQjjUb4Ek94UN9NNFvP6JSuFrR81fh8t7L
0B1vU8HjHsy/nUDB5+ahgzCaL7G2sFyOQn1VDtwr3NMWbPoncKqsH7T3m/82lYEh
Ya133Yx5uBq7mpY2SGyAyzQoZKai1OJeRfmbUv7FeAFCigXizQI0P6pJHf0uV3vD
0tSP5YRED9qs+BKhYwE9Gly1/l/VPZUAIs5lvskD2idCyAYbjrtCUdSa4oHpFI/C
WF42WyowK0dZZdlACxvTxWn4Nyo6Dx67alNzfLd6KZhswaVVx7viwbtGvYFB+4cC
KGH9n4hxNXiewUvKY2ooeR8VWOjTzUulBqBhoLc2YfSZ0hIEmqBCiGJcps/b4XMf
IQ5tnlvqW4IjaWwxCAfzYTFfYNSfnZw/czDkWWg8OOarnDLqG039/tNwro27rc8+
WKDt0MmZpwJVZGCVQ9P4csQKcYgyFN5GYnNz+Rx42sQw+rvzGkT7fCYszX+YLaCe
4paIkAOPwRhXzev6eDa3wAjSZ0uuCR2+j8mrlPqI464ALVyVpU5DPcvmaIYd+43b
tS85ewP8J6pHlh+awXLw1wJkLew5NJNAiW2K+vN2YxCYnx/mQfd80S17t7LZsFJq
Vy/IDKDF+qHuuZ8DaFVnzzRFFcsvy4xZF8LK29RfrA4FSLbQCPOey+8mzEt1Vxzn
/PsSKvR1IzfL4sgQT1AyDDFMWmOv5Iv00GBCcmhCNNTIkBO2d4fl5fGdH+C3BjYJ
EEJcEfpQj8q8DR261hpYH7J6w2iZde+8c5O3xveM99Nv6w9JxunhghYbGzbxKd3f
hSnpL4RxK0oUegLDdVNBNGcT/CvLDShygd+oA5zmtsQiJ9YoLiVgvrjU2LPdIQ5/
9ooN0ZwbDFqngygGaceYQea0qA7Q3rTXA7Vm8YGuUAeNxWaszGjsD133IRAec3Mf
KLr+gcPgFZ1CSjv8oZEWkX7kppvS/SatvdDQsSQN1LT97etIci6p94VbGfKS3LVS
6HkH7I//J5xu7ASERBd4jtlRmBQwfqF3kceGpJ0ekMrSxVoDbp/1fyc4ygg86Dna
NXoqV+lkyx92cK9EGNBamJc46zZAsmDxALAEZh4JnC8qlLsYmM7zIoRcTgeG3awl
x+VzB2g8wq9aWnpLpzw5sPrgXepxrdsoEA9QyjJda0Voq+ImsOxQiAUyUxF/WVlM
LmJtrKbMnPytk5tt3NlnhYh/E9DHcIpcdkdXGzLkgw7lZGWVAW3wKOw5Jm8HoUpZ
yZ50c5sy794Yi9N3GnkYL42iKj3MAbEH7MuQWybWKvJONIzJxSyxKuTmbzAsB41i
FeMFmvt4PSHQewTYgoeX6btrQj868N6tjZ6fEPDLyoVNJPWryaInmx48exTqPRj6
/SBoFrNuIMNop4jeP7KgfLQl/8DQzS1fw/RIb1zQjDCw74sFfNoulTVgDmDfmaXx
/mWuh3XpkdKTMJqr7F6JCicc7Ufr3w1LvHRL11dNF1/HaPOUNP2UR3+vS212EWP0
1ewIaHUobiZn98hGHGPzgx56xsHg+w4spRK9UKx+6sJ0OMnXaOJU4Zl/VO2QSwdP
BbHd1wwu3NtSnna89RDLPtOwfckGx+tLrpuzr2926kPNC8PBQVLKcLe8a26qJv8m
yWa0K1gjDfs/sSELrKOv692MBYP9ccyWUfZXBh7ZAU0X9TPT/Fef+f9MYEgIgH0V
5FxDbkR7PfLMGtCmyuHctQW0f3wAeo+tACiIBh4KLbKQHiXa+FR5ajqz9jkNnfv7
KpLC7566282w9ZALyMJUYTYixBOM1gloXeb/tdF+nW//HRJWrnq3jZVXC1yVQGhi
F+1nI+2Sni25zvqc3sZdB328af6nimwqEyc8/iBpwXLMmEttZCLAjGpYWItbInIe
PoH1YbBap/INlI1P9smO7pYePovDFU2p0vA9xVAw9AZs9HZRtz95wdbt8HRqnCZI
ppqi1nqUpM3wY++z8S4sLk5KQj7utOrq+6rspC3SopbuCWwQp5uciWdRhhIeQqJ/
nZk1l+bhIhkJis1Z0I1I0fy8agF+grwF1MhYn3D8PRyj+IZVztkXT0QJjF4oJzl7
FF/4gQZ4RMjUdvp6iP2p6ES8TS0P1afwLEZVFNUEYLAiGrDwH+Eeh0fOolyOcT3p
Mcq9jaKBt2lNxVNVAALCel+4Je4Q/oBTRPuUlD8Ndo24tNPPlFjh3WZNr/xncy3n
s9BFdyR85RXOYw6GuDbd0MIbCht1gzPpNeyZ+7EOVEsJYS6yTW2NJ7Upx2MPkPO6
VqNi3UzM6T/7lume9yzUSA5DCUDWR2Ae/sv4rljF3cyVgR9khAr1buQQtQ/4abzq
Tn0ceS1rcTYJlYBdgQmJ8TtDEFyrKV8zgOeS46t696CqCGXRgG4P0p64n6gr1o5g
OQOHoDPyVm0I9OQZkjVyiqDnhPvZ3Ie1pTqtZTNH83tPMb+DydxmnPfvS9qGSeIX
EB82jF8nhLOf1r6nQmcNhmWvoWzQu6O/FD3VEchngxJ7nYEPAfwi/OitID6JvUn4
4Xv1VVlYc907sSWdWxKmdd5qZQ5sjIHCYygQ5aF7bovV3w91nXv+HJ2/2P/msy/R
q602Nt6s17XdDP1vnbrfDjjb9QWifTQ5Dk5SRoPZblKTJeVozn6vXcPzfUKhcK5I
/rQLomFmNzqCYmQpyM3Pg4g0kOUt0mcGFMLAXf4KTEOvyX5iKHLkzmjpUk5jdWop
fF+hC7zIWUZoSgn0+5QMnLjTmp3FkA2SuPilmXMATf8uKftB7efSgLHKWD0f5SvI
dWtC2QGk13YwFQJnDi6pM/nFtz/6LCqIo35P1tbb5EYPAPdChlcfRcmXi2YMJ1Qe
0otM3TNQTSNhH1Acr4YB347H4FqPky/G72Lw+94aI8EFMvrdidf7pbrgFnTCoyFH
gbbcSb5jY1XYR4qnPHlYPmonuORaqjaxd/kKFrX8uxcoOgo+bE4rUaj9URj4R7aD
aBWcQNvXrg5BIVrsEbnDjWdkRuXBc4rjQ7MJq7RE25U8fUiQc/zJhbfZsmsq0kWc
Hhx4sge9EBfwxq6VRepaNzc1w+nUQxEVmVyDP/25EmfLCxzF6ujfPZh3qlAB7gAc
d9EGocXHzLLShLeMyVWTuqmOVa/qS5oqHPJCncYwOKA2u3yP9nb71k9B7dIHIIJb
+IMfIBBCvIDUZTt7Y7o8AbW4qiJ8tDLVtUqoHG8GGCz4E9n6ZwFX0J4UcSDBbeuZ
DonqHFcw2r9mUNG7/I6/BYiklgPZZaXOvVSyy+E/fdpgxbE5CvdrxyNr9+qf3x89
WUbqfRbNlxBq4c+De+8vjY8SW157T/TsmYoxdxQ0+Fo108db2W7L8GMzQ4s7TOwm
hcbLkiYPxdCINweEUXNhEVOvpBV0Vdk+9EFzJH5wgft++PIKt2oBvSECGoWJMs+/
SfC1wgV4y6kaZl1Az5FkLlj4m7KgmxFpyD9vUhZutihrpGHeBDJQ6QNSSVF9i0T9
Cl2tRsvw+732vNXFs3yQTVgmr+l6jGhcUdKnMNzHM9vBkkURNMltXrDYXKTGfiCe
bAq0DkDwveaPNRhNaTFwUHpjIWYdhDc05DxcbKI9bxgtMHjPm3Cd9QOVSUa1gRWD
WqzTPwMBVgDTurjoTCzgKQo70FkssK6vlfUa/6/N8b/gAYiJow5gwR8DWpuTNVEk
/w7AoDr2j5VvYjcmf6wnQo3Q1YA4lycWsqxWhqI/+n3DrH6kMU5j5IHrF/ozhsRN
Wky3z2JTM6oc1ydql/i9ibOPtHxjrA+3mazY1jXZr+QCdfqCwwsYN4OTCTztQXR3
jpyRvF2yKBhsBg8FjY0ki80zKgd8lsiVDcTTVSbTRUgY17AqSUC9V5Ex/TehrmFc
GVMFgyDRWhbLoup2/ZUDCCDAGNF3rqxHVSN3BvK+D4nLMgGIqzer/todnurv4BzT
fvstjylae016gAdgo1joduXYq44nSeSbrOcUg4m7ZCAtUvUOZnlYyBxnGZATizcH
CngnNxb1cF8OiaB0/JqGxwFR6ftfOictLxD2FRygDaeyE7woEJMdYRU7a3q6ZlzT
ZSlizGGyfrvA6bOXfmAj9UX/9xiC760fxjNOz+e0Br+YfQkDo4Y63uYpUhX3ZZmf
ByMbw/xUNQKG+yULNZAbEI0nq7UHHOmmjFPUmOH5JLUSl8VLG6WIjT8u+UQj1YuJ
IEOXzogqo1XUe5Fd5ObPzcEM24DnZr40zhl9YEEFjdzs6GayOE+BKre9qb/yvCeh
vHoVDN1GHoE7a2IOKVPHMJSmnidYeIPoAgYn6c6BeRYGmrsJpSHVwDQ9TANZsKNV
JV8ravJ0sAW/sQ58lb0RezpqKKwlqW/lCqGkQcgbGtRL+ssZ+dRaTYDRNkm81tHf
RaumR9UvM2UkXkis1cO57PYc4sxHxebnbeg6vnlUYWVulJVMsbbkzDen7I9fRmrV
NCtq6jMuWCZ39pX4XqzJ3pGfIqGjXYHtrAVDYaC0pmD3PA6oExBylRE26K+8cb2L
Uylki8r+bd0P9emSP0iZmTheBeSiLjx5fL4431kES+1xT+AkvWUqXv3ngziFoDvq
IMEccZplqrHxXt29MnJXPi37sDce+y4BcmSn0MB2ApLPNWxLfhZopF+uf117BRSu
G+mIz/VOnBI9IS+t289abRYOQpO6JuIpRAUX40cWOX2dtYoDp1/9U0pA14xqRuA1
1rg+xKjSnumxxW8GWS43oEt8nM69psFa+Za9fR22wI4ij+5LmejABblE9GPx5KBe
YB6AMOLov0h3DgtjeLI6mb/DWzuNmEGeYWEn1GMzzfUOzeT+l1rlH8G3Q/3c9EYt
iLU58rcNN67Pg4gOss36KvGMy4OtLU4HN43cYAQeeUBX93OpPTT0dH6k9x13/I1z
TM3PKXUu96CVQTV5V3Nvn+cMMv7YTwL7lBT1OOsMdI/NpTvvo2CgQ99+Qq8/Il1h
ygsJjLJARFeXhKCsL3NQOyQMtw+mB+l0goglOoN7m7ChL9ZBkm8TdPHi6XweQrHm
t509bQ0xNK17Q6zZz9EcG9iaYFhWoPrVS/D5aoJ4/9Mm0R1/mACmcJ1QfI0g7OXP
+BdTe4ffoHY81SzlNk2IR9Vt4NorNaeKDFBtuGqMMmkomrYEp4/QpGRKraEY0+1W
/3KDpWKXqmkjAuGbzfLisM/VU/dIIJi3s9IMMYgERLYYbhLuZ7bBMDzrCHnwyiEc
HBtrWiQS03YYWDUZuPNWBxrGLEPXSzjpoORyvx9UjZ5b9IZPqL60H0wToEIX2Ym1
+kmweKVeOlH6rarcwLzfKc9OB1sBxLaMC1VYgB9jev2WhBTR4YakcEnneVg0VsQE
u1or9TliPVEURXmqxP7AOdkUu5bl3d+tDIbAGPU2pMkc6r25pIJ1WFIvLW28A4wF
FLuf8fr0S5hCvICb/5qUvceBrxUUwok5e6JkZmmGU4rAh7gl+SfoPL48bi61o6Iv
q9Qc5xDT11k/M4/PDb4OszuwEj08finAjad3dOzWF7/uWaXM5GsnVr3dhikLgalE
R76fZCkLhDBtZKQoaaEiSC9voMTEw/wvOZjJg2E0OWFwBxLtUeEOlB8eMUmBj+6N
yVEoAbG1ERhq2Rq0d6o4DGBBMVCSBwCTilHBzA4D9ztpbyDDtswR1jB5xYHOfQpD
qlWZxbndY4OIDu2aj4pbZmwN43eWmLcztCJV3cOaaj3AYrnRC0PdcI01KF7MJAUf
C3o8LB3pD+opT4XVWUA3WrTcMbICzc+gaj0zFHL3GDTCpwZFDw5dfhkiFANH1OX9
I/pY1Yp/6C1KIhWgEcD2ZkiDcA6Bh3/xkeqwBvX1FumVyNdcxzoR3nz4HeRes6SV
5vIMousN89lHmV1Rx4i4tEeeLTLmLG2aysCRdMJmw2MBbXOf3QSig/DTzesX2c/Z
oAthpZCN3BrkkODR4cB/FD7pxK2s0Db+kASxijKLQ6iC7ll6psCDvMlW7H+hCIn2
DKQAtltfVjUyDRTKD5Jk5/miH1g7l+jN5pSswNpz7gS8TDkVXxU54NX+bVBGQJQ1
Zpvv+U6mU3NvJrVbCUoyt/wXiuZlRgYwdYxQdQxF+iVgpqWrXGy1u2sPCMoAI3Yw
+ykrzXQRnpSrQVpHyxPTadc6uFKugF4XS7KnkLF9dz0zXiiCWVDhG8GjYU88WaOr
xmr0eXvaozQ88/bdepn6SJm/aqpTAe3z+LiZMPUZ6uOCuOqc1qsld95LyeDctWEr
IKx1fxH31kz4+y5QOADIumK/NV3XYdSNtI0THPhVwqKYbZYPgv2NJ/P6QkX55q+O
GOo8VDiM87stUWZ+WPpIWGh5kLynmpO7heY7JstieFCjp/lw870St9n7YEjuqxLS
4zujcqnZXq8/sA7hnxKSnbu9CzysgF/ukvTecTGTS1eSylj7muZOZCy1rCnA8U1J
bvE94me5rkh1ir0UAU2pbP775oaRHywrinf302bYfyAFraU+MDsZnSXPl4FlZST8
dnAo6GPaBLRin23R17tdB61GNtCDTkcMA7EVOeKGwcXZwN2apNmYdX3LZd3dtdbp
9ogEZb9h1uAS9GsmkhSoQ7G8MZRFoiXXkpCKlYjZszMSPqwPNZeKnrOf8x1Cb4Hf
RLwcQqdRYM4VdcV1q/JW3g/pTT/nyedPjEfqdKPPIDBAP8sKkL6jXXSoM/mc/75k
/+E+JIjRFe/5y3xijKsVqm96TFhKC7uTTY5tq7pXRiTDTKrDhdLsYfotoI5dPTcW
28/jm5JXyhbYSuDJ7Bly2drH50G21A4seDDBof4Ph1tF5IAFvmL8IH6ls0ch3jkS
ehHNmyrhrydvXRauGbiKmajepIqpcnRUq9mDgPWbvBpj4LmYNKXj/k/NS/4TAfDS
4fQnuCKlqk6SbUx7N8xIQUhbJymAAZnW5DJL/MyxzTz8zeoi2AcY03kAXHXrVoZt
WhHnkyN48QWUZ6FI0TwXNdDkt/xp9mooYqlqKU8fpAJZBWVkfZJMVahlEXoA7liQ
oa/ZE8R5p2UaCG1Z30Eyj6S9CXW+BGvMf1CKwmcorOzUf/Zdlj4xSfTqIfDeaaEY
5sxGzLO4ZShwOCePuFRtyg0KO2dTt8X/QjIVZ976OeJ/xQmsGBz1hoQhtRsKi7GS
HhTCareY8FZ0S6aYBObFiqU2M/3sBRn+0YTH/7NMMmnfdCxw2M1BHPksZGJDPKKA
dL/3C77HJmwVwo0uTDCEFO0GO4F0FfTy+mCQkT+fX0uVi43nb9mtdHQMtAMTaLUA
eKQjAbjG6igbeoUQxKUCY4U1NQ6XOXuOXg5b5rA953YSSDUpc6NyeKKpTsKdYq7P
n6FFC/xn/g7AIaIURwgH90L18aVEf12X6Uar7UduSXTQYCwtVjziAcrCltiM3Btg
vb/k3Ls5JIovtWTWFtZPMXBw+XPUe12Ib1n19tnQY4sDwUnEboagbu7SAWmYUNNl
DN3Z4KKyMuiD7iH54aYY9dWB9KJwDhW0mwYSCgxT86X+RihUI9AdGxPwAa+DdYSP
cw4e6nkMJC77HNWVQEXcm6qHoLaXx6Y3r6oLpHCA6HZ6uHuvDEOrK6AjW7Yx8Bmo
nehNQR4cXnfgKSQzHEgx152Dj7GSjUC14iIt8KNnKcI9OgVPqiMUkAxNLGukRXVF
HaWndS6yIU2NBTzUKWTIa1tlnuhsRIPh9PrroEmB/OZaGVrJi0bnOkLn9VWiw7po
wy3atEfox+7Rag6jqF4Z3hBxlCmXoSMwDoQvGfdtpfk7UbOhXoaNgZiZ8I5OwkuS
ZmiAVex9PXMuKcW5FSpDJknIjXg0A5m5FJXoQtD79mJxMblRcMBquLk5vOB6bCGH
JLZHqZK2PBsJezpKJO9gJZ/ZmeY/etMz9V5RpotQW3Wl70kqrlr8h+q5ougW81WB
3t2tuE1Z34Z50JGDssNXDCU0MKm24vLJeLUH2tP0JYzn5zzmfAU1EEb1J05hmGs+
4DdwQREhbUSAK0Df/d2yxie+wt6zz68b5eiX6BGaIVFoDlDwM4oL5XSeJG7RpScr
De7JYt8HArUJFY2YkZmf3aUh/qp9GTtedmm35V4yH2MAUzTMPSCNHAcLzQHH0QLO
dUxnaajiKqlyGauclzGWIt875sY5U6f0uEbpZUFHzs2XTEFw9wrzYq1E5yE7No5w
tgGVeEpf/9tCrmSLbs4PPCpRUiam3cet1kRTRAQyzx5rWkhWw/tCsdAnlcLguFuT
v8DmpFrU/2fKWiIsZfajfBaJaQHJmgARNgbrpaj3Nwqd+SlR1Zz81lpaHWfzwFMx
iJox9nScxijMUC9DOBKiBs60vSjgQhYTwDqw8XTeoGnBI5EFfjjZZQ0Po2VaPAO4
3T7846U7Cvji4zHz0P/+3WQD8eqnPRmK5iZwLFL3B3LzjL2C6SSG5d7/9g6ke1Dk
2ayCRBBBOJmilNKVWGLXohOG+fZIAUShieVFZKPGxChnFYYO9ye9McTgPX0cPf6c
cd8glNLSY2KhFPGYcZZ0NsmAuMTqpXThrWoP+Ae2tpRF7ONPjjqlnFG14Zr9QhMq
hrojx4oW2wBTp6sER+k1DiuWUO1a1zxZN4yydUqzGUu+r1EfxDBhbMDBykwKUOhn
3Mz+Ia5wbc29RMhExXkf8Q937wnKTCrp9WLBBTVqztAWE1NLWvNxDo0bnC1DhGyx
y3lu6XwQeyk/bn4v1rzgzZUb83Qn811P95vFatpcP9PIunQvJg8biSLMqQ32So2I
qfUkVxyEDHx+hpLyABtGjDJqPghzGPsO2O6Tyav3s66Z7NO3xoGkvFWcxnIyRuGZ
i0dVlTnKjzNyEOxItuz2bbwEzUxsbduNsZ9xdnDLt6IZFuFl18sVv8ajHOdoGe6C
0xlQ+6R61S8Q5+mlGxAHXkmsUNaKWwBqZ/d1MilKsn4yMBRq6fmCpsVWK6Vso1UZ
qGGtU1drDu1uNfM+4SlIgeBt212KhWBFrZcvxu6a8a5QAKsYm7KeUmqWM7xrpaZQ
ql7qOn+0av8P+qdSzg/jhxebhDsvu0Orqj1sL4baLkMpQIr0hMtMxei1ZTz1Mtfy
b03HgIhA2b65eBLhxSxgW8bYjn1Uh92FQQvmn1qgNXJhV0RxfbGlsh2NMz+cjSMi
qFrmNNmtLxmieJIk9uo6Zfwh6bZYE5yUH2C4PTd4HypXMuXSgst+r3n+SDOVJxGO
Yc57wAXSCTITGv8XHITUegDVwC1o5/ptKIdU9XTIeAQ6eVfCTadCiSbdiREj05KX
6bffVOOnKbBnfpA4gQEa8ojBIX+WFa3h/WQ60oPvkwfVpepmkjtnosaZ6N82tMZ5
7Eb6VZtuqp2zQboIKtlb6ZkYnYHiY01VzhkxMwdxKt/F7jcgjG0YPUfiowf6mT9t
FpFOX3idkymgqq1oYyXXjxeLn6NRVBLFLNh3mgbm8t02DO/gON06I6THa9GtC7NN
7wrIOQ/XdG5bcgWRr8rcpMwjcH1HHXHWItOKIBqGrxcgoa4djhwSweWQ3Col6hmN
YVXczsH/LZ5cH8RRHWkXQgOcwEpH950I5yXrnp7oraWd0Jz4VJ7e7oUb5uiXD+wO
h4wVLg+z6UAUFZ4iJ+wQadOUdAEjQO4qBWdhhCzCUmxNfe7YigEX8OR7dOCS9vsI
Wq5B7KjlE6U4pTrw2se+ZsNBud8ISCKWm70xVKG9Ugg7CoGoBmrrpOMkofZPeov4
Q/khG5NNYPCTDjXuD3yf37m5TgosDTfGKkjAq4Y8movx6oSniRIlhVhRVRoos0JV
G+VkK++k86KrQuEdLuRKM7x6I/IkXiUUT/kBitRh7GCFIa3ovB7r1RPXIdJd36wC
f55TzZxcy5L0Dtn/1sBdgYA+9kDCpd9uZ9UJjAIIMTEdBJAOso5KPsvIJCiuhyOQ
6ww3Zs+m7SA2TYBSJRWv0acgzf08T0uVJ8++Rk4+lY0FvCCmO58cJmh4p7UvHNir
PN0gluZ1cRf/gfLLmCih5b/PIeP2zlm7gO5TfZxZDkuawiCWcQZ7BnKuoWb9bJ2Q
ylMNuMDefd5CU766U7fjGxCTejHSvrZ0iDpbyBAcFeX2ozCCUrR5GpShiI7iws7w
Yy6dVo05zFOnLjhfxNpJ5DDrEtaBAw4Jbz2qM+rFI3dlTF2759LHWsgZyof9kFkt
9dV6JJ/piUk7U0K/GyUkZY3IwsrrbFPRBL6qNEUl6nGjBqgRTlP5zyQYFH0qlJEt
HOof6R3ZzB6ttlNPIQFuSiqiGAYNvez9kGnUozcxz46pMwf7zvopxmN1Vda/ZigK
pwOttdn3P6+a6Pwbzy9rOERq6tiVG9nCkqihI3HwrXArR+cYE/WHc9VckXyOgM3f
CxL5zdcZ4Cq+OcrfPRWiASf5XkTOGqHqHw3rRF4W3fvIlqMQi7LhDjQK6+wU/Kod
cKWIa5dM+9kFWGjNXvBxWHnNioxq8aINvAhDLu5SMnA19ChpjsFAYaJ60nyh60l5
2lLDTmg9YJpSrVXoH1gaDdKpZUQ9yDL1l0qI3a97sg0MT1HBOzqYOaGE5XVuHR6u
JAHM/We4UwvotI7uLnZGTC+NneMEnT4DL5ckUKGL9478o2HyOuC8TAJwbXBHdT9e
Bpg+PKVBlA48GA9F6fgm5rCy7sRA650cWzdAPe2szlJRKO80ZIV3MoTbofDhV874
ZdW61f9uRbMY1CWBgk81755cClQJLyBjENbKZaZ9pm/aEDIC5eL58yCArXeqJ4hQ
1i15WIgXpxzNjBMBQQnvezq4Rri2TsXzox6PqJY1vm+1qpyVFTeUy2gBdHuL1Dil
SzU8BAcaJHXSkYUUkLJ3Rtu4RSJmje698JqXTeIRopuccux7gviGpwZRaBW2d3EO
v65PzvYHmE6OTqRrHBflNx7JDuamrh7huRvTpE5y5uZ0oEXtGvuQwuvqMlhmD95Q
PorQuYbn4SgSUqBWB4vnLDdE7lObI7aFDs9ILJGaD2nTURi4NGEaZpmRh0Ar3lRG
qvLUJj3AZQeZUPrx2XRmPw7qfmzZ4gTSs57SFsALVfOdREx4tB9ObPkDM8pb6jKr
AJUyaFhpKKVCSpvs7Ee/6xm4JGYryiZqYGn3v6Ap6WoVxKznycr2U4tUbmk9yKzA
gW2llQbK10pfAla4eZooxEP1OWJ+MOJjtE/8xOHkrc9I1iyE21dnn0Prz0ZX5+dK
EfLyhlEAuErSZb4otK27/OLggpU4DOUiUhQyexqKmQaGADtNX9kkijoYGU37CaqP
eJEnU3JcZV45d1NolbV4yz4seq/9p5QLVlhH5lZlcFKRjN/JBKfPtXjZbYESi1r/
kK/yeJP67RgCnKDV3Ku+houMxY6qKVBgaN4ioxmSe8wLlV/4pcexFv3XiKZgR8QD
4TFM/tbFIRziRTJeY5MRKguk/QqgOZFU4IKsO0GSKqs8LgW5oCiN7pnJupqhpbEx
NbiA5K89lpgqBN57MB1qOI20IDgPuX+DCNl1NkM7taoVbkeRm3Qc/1Yii6q5RA4u
QrPzI1vhaek0WPIEwbW7FD5fJkgEeTrUDrdCfgR4R09olBbL8owMwY+q/ZONoeFH
csIsop8gFbE7A0+NInXLjN+Wf/ssNMUuhuRn7ecp7TZI+YU+P8WXOOhI2T4S0w6J
wDDhbnBNhm4DgmCy2tpSwqeaoBHPOLXC9ofiaAGVoeEn1WOMHw0BFBIsF3FMEJtH
ST2BHs5WqtoNtVEA/wR7hgx2AGQRCZGYESkj4TY9S+Ltjr1QMhcCGvYBD+gxV36i
u4vRk2b9v5LrLdQTPUS+tHaxN9hrnbr3BFZ5IicTAzHVoGpjWt0SPo64yYHi+9ki
9U+iTNkEh+U5084BexbeSBxMAne7VIPH6Ms4b1v/jgvEgHSgPlzCFX+e75wEjL0G
XCTnaoRW/wXxqB9IgO7//uewgFR75uFweXJJEekG7OWbfHcKgalwNw7C+ll8eDg/
oaEUgI222zrPKqgr4PxCqqhf4xpbJvaB9E6bnR+qD7UrzSqHRyG6AMGk+6j4n9MM
6YIxYvsgDwIfMQDftObAiPstsOGIRqzimCxRdK+hzAjpHYATfns13CrqrfEdUUrY
LLZtTCt9yOpfaQVO9vGIQS8AhDVSQNU6A6rt89eDERnPGI4L5U28O3oy2bYym1B8
azvHXo0/OBzrQpMGgqL67PUoU4yoAV/ChtyDL9viQqwK4KpMTAtlsdKnnjbeefB7
LJIIX8cR5QBO7mCxvXY5LpASwTLLJdZeyfmyKF0Y6uTGgfxQX+ggFnHmstagEZjm
PeeBVnyqCxnesb6CejlK8J2CIMHm+hZTs3Uw5qgviBNi0glSEbtFfLTKXJiB2Hqj
5lvs/+/HrnaVE3bWHj9TrVGwTKj3FGPFgtvzovf0U8xPfweeOI6JoCEo/51LhVnd
OVrISO6BmJ7HAgBNmurfeTqYpz5DcjecHSh+hqI6VB8ntvHG8OgFsjKyAVzF/A7v
GwIPOlL4nhwNqV6d/PT78r0V0DQQp86Dw3MRR/5Tc2pVWc3/F43ogPIQjFe+63Rq
7SbBwzdDDcWQPzNAz9w3QrwEijX5ikM4mrl7xD97/x2DpWW3p/caxzR/Uij7jBPX
VFp+NYqGO3vCxhio3g5t97c3Vrk6qKXHI4UxnU2ucgSuOArkYqwBuplRFhvRBXhC
ruopHwO51FUGXLTmaFjRnPXU7R+PzrAtCVedkWpmlbzLM2h1GE2Tnff7uF+i8HN7
3ObG9Fptfs2OndM9J1Pcna9OpxQS763WUGg3eOyqMl8vdV62rKKL+2cbBrnZiuQv
TvHGr5gH5BQeymTDXeqacB6U6Q9tJu8sE+dnaqbEF+14+Vp70H9XdjfeHpb5rtQx
5jll9gVj6oeXKbNnnUKZo9roAeDfahlbXnJ7UGkfxRkd99Vj8dVH1oX4Tx8AD7Xj
wJHuj9sTOFX4Hrh3rBJ3O6DwPioQNj3CQhr/k0lLvRoPTkuxsKLYBeYHVr7HlsRp
p3eA0+dOkPXdhE6hknJ44Ar52YFKyconVzjyqiZHjtSaaq6bgrPvqqp2ShSnguPw
ghsp8/hver6EnsBQUMJ+3WVKpj2ucj8WEszFNAuSttcrwZ5ifQM6z2tt0tub7dk5
3gFQWCe20nQNTgK+RllF/NQB9yBmhwCOIEU7iYe65bpjRxTuWgPKgFYbIi2ImEeo
d9p0jTz4EGCJO2S+65r8GrGynoaBzkULP5B4WESa+QrV1NODtjB7YMSXxHU0kikk
wvMBnoS6yjxkQiAqr2u+80NN2ytKdMJKUSxDHwcygkMjfibikX7knx6/h5egYR/1
plbE1HNm6kXoUSSD53VnbS4X0aS9LTiL47PuP8zuxqLYfPlmkZyP8GpYOd/TluwK
hn8yPX4jn8D0cSHi5RXc+ZaChCGIbn5oQG6SqsEqiqtMHzn6L7PDEyQ+CCZ/UgJs
3d/xeNBOvLzk5WgTFEDM+lzdMA1OawlXLpFdgm1+JuUGLn00XOEtx5iwUrAXU+q6
jPtezUoHoOEuH53XAACgIJklUHitBBR2I1WUpoAe8/qdRrbinT14AfZLfRxzypwr
yzQWu61cEvjhXd6wO7HmRdCt1UMd5RFNZigN/GI9JqksPSQLNBVcVKgMguOviteL
SJqIS/DMFFqUtbxZfbZoWdPq3D5GnluRnrCcL+0+V71DbFzT1/GHxXDjeBQ58T92
wyXS0MdCIDVZcCf0aTPr7tcsJEC06WwW8EtF/McyI3jSdnY33Yy1Ql3XnODu9I4A
XdP2SYCLsEhCM/IAeVCVXX1HN7npCI6ydjnU3lO5QCqxDAufPKloVA08cOKxKjeM
hI2ghHQRanW6wrtvqDonFh8I03G6LqQFRdjtzUqwuqol6xMgfvf/TGwT9l075SUC
1dsPxcLH/vidkOwWg97zN48xgS+Hg18CYIAEN60uoUQ7GqQd1SOZgJSlj3ioA0/+
sHsK8xn43HJpJhJjaqerJ5nORei8g/G+ZyscCBE0N0gCRGzDlcWH2S7JFm27+gr4
RUr/Wq0ARc8JzwWFBe7O8RqZP+b0TBL8V5w9r1uVOIc1toFsqIrTJox8OL5DjDuF
771L76h2/FAVEcC0NCbUDx1rLSsl52KCT8ZdXCrX7008r3lVWV9Yxc/LhNOXUkwI
JNDHNL44IBL96vCUDr3gmXgbWb3lfEP0Jfu0giWpQ6FE/h+HPl9IVJ16GEzR1nUu
tS3StAL1Ry42mK12nJyPUdzxuchaBjEzdb3wVTAqkKx/UnJY9pKs0rXlZrRVG3L2
ecwzRb17UAAOhzIf+8TTMQnA/CDZrbmk3qHxbBSSUCP5P3s1XWEHMsKlvz6ELUGf
+3J9kXhxVgOsQ4r45PUWP3aioRNgxk/gu0wjtdvjWgyso94O77tNg2YaHTMZU4P5
8exSxMEpOCXXFUyacfvVnwyTRjf/K3U3FHr0ppoxQJOpYVT7Fv/zrOKY361sW4IB
TKFzxScgS7fny9xV/ui6vUIi4+BF53TzsXD0cnObkAgDVOGS3C7YFgHi6X0ROuBK
5xgH+c1wYNfjI+HBIqb+Qh3WQ6Kn1XzaJiYpHgcP4W3rHuscQ6+9Bq3svKOKLSTk
5zokuKcxga19f12anqvf0xFibAE9v5PCl6Su9bZnATy5Liq9gQ69P+N+1algvIJg
Qm7oelT+/5ZtuQF5fs3OgBAKxfTMaGoqMIJaL6OTIdMBAtLUMnfKX3ftszsKndlK
Pi0nzo5uH+08hU6MlzuAdVCf13S9giNvu7nqSG1+soUC6VDG65uo97G4BgHVdsnD
OKAIS25wRfZr6R5Awf/uF77yUbzyHQKFbVe1aqswYAY8bfjpmVWBa8aQYkh7Z4aS
6MQVzv6jq3a5iKa5vZ09wuRLf8551O6NWowfgeWuJgUR4ARR0aAwLLN7Zw+3ZTEy
2StCa5+VkeAqZUwSCkViGVDeSmUHCjzQNKB9FH5Z11y/ee4dwsbgh52LnILOb/XN
TR8bBONV1qiKGij3QUYjJ2ei0PzCbtcMWNm8wmSEDTw05l1GIUUb9PvQLU2WXtw7
Hj+/iRiZpZ7ZLAVE4cX3PwRPYxlzs91bi2itVelouAiRljULPjD2/6xFDC3cSFtJ
p87j4L+aONX73cyuVDqj+WwiTGxFpf7i5eocNnjvUdLZ0mRVsshWHUtQpXLGgss+
Pmqm1ccr9cKNq/5wUQC+k8J9tZWwOFEDy17MD8LjxfkDZ//P7vEyKR3iZ8tLVJey
oeRIhuogy4Ngi8LCDFJUzdAvRvkJPzpHGW9WBKef1Xuk5rm9TWhLODP2n4BnMAVl
JgG0d6iBoRUh7AWJ3jZrru/3LEeaAeIgY90ij9Ov7noK1DVUeIH/tqSTlUE8G6IK
zWW/nJf1rbBGS9c2QwXs1vJcMffLqt7GaBYiytmat1bwimXUQWFvwhQkm1apHGjF
xdJZ28aDhfkqBGIycQ9fhN7xeJaJwTlmcW54DAoBQpCO3m36ZGHv+ly95dA+/yso
w2E9LTLivCOL3pK2RTfs/j5VDsUMvav49RbT6xlBUcGWN0CDyOvJ4DGoaeEd2ngu
ZZzY9umJ/SvnG6F2qbj0g2qnzDkb0w0U/pSmEpBBDVFFW7jDRA5zgteQ/9d/2eQn
zw7snc9Ab46CGiHFBZ8FQmgWyBFHqN/AjJsbCKs/k91QilSj+Q3+fGA3nOr+wFZB
Eqr2Kb6VVoOC8G+C/g5ntorMIhMmqzrHXHyirytF9N6x/m02mm1N+S0pBczbQkab
m8vwknRKnTT0RxVtuQsufkfrEBfDX4+FF2feS7R8rJFnQMybRawzcVhq0bQCpdgo
zLSGx/RJmAfe4ANbCh4M+L4i0CWgHyMSTuOhVY0s5YzPOFSMcct6CGb0UbIBG6oD
HN2VQV8S7bJ+5vshf3zxZGkpbJb+/oihGNVviPu9lPxEOmlDaiROMlNLTSQGXkC/
Fo4FttjiGU5XJ3rzM9qOx4BLrLfIFZgOC+v8MAPYFpNLj6A1ZB9gxNq6N+cHoKdT
IlrMfgyo0aMpl+SmwqnymrCswccukWBXO8FMhuTU8owQMD7Qb7lKn18KxUwP86qZ
SUtbVKyscJbznqKgvPs7OXBxl+yRTFG+4Cmf7IqTpeLVCEELXkDDLLMy9rkIYUXn
rOlxKWDRRleMSJp1le1Fpg9vfl54hkcSulAw3HSK8FfdDo3jHHChBWfZXdwmycu3
1Hovo0ili/OZPiNkF24y1VrAkMIi5WKp3g+lM/EH/7H0h0BL1NsBPlexYGpBgNMn
xIVbk29u9LeuACeS+EibXwe2Ctz0QXe0Ntf/VxLRRWT4BVO/1E8agpP1CzqabETv
7hsBZNBMI2Ul2qutRw1OUol7JQ0BgTZTli17DHbvOwhCdAqtZDvMi7jqv1hZJ2oE
GFmWNejjPYR1h5Aw3JWiK/f01ZBux9ech2AAv3KHPkF4iTwNW6a+oP7n5yGHgeV8
n2+WepO4Vbf/HuyUksXr7v2a+GSfK8jbK4JhxWfT7gocyMwBJSe4FdZDmdSn64TG
j1G5/KZex/2mRXdjvgyxkDyfohju6qwv1duFRxyg3AQ1yhxFSgL/xa9+i1E2H6io
VaYoeiy8IN7GqbCEdxbk/C2wgxnyj/jX7jbQcHxucAn99dPxQqHfdpud/od/hCBu
EhcXkhiWWZy3J+D8jSsl4GvIilWp3c3pFQQYmyfd0tkyIj46+loMGEl/I/RGtdrV
3idBK3+MJJsX/6zcNLCFwXbBtwJ7wqpCYayqQvyfca9YkOUiUOtayDkxzvyOZ5Uq
M0XMYwebCN0SDLk2wZ9Idjv5Hn7BNLpWpMopWYxAGDyQnQjzLxYBA46Wsgtfb4eg
g9EcYE/n9WCwiODFDZyXEjGzl6+cScU+9X6tUzje5CYwNQFxUdVY442/Mbt+Cic+
IRJ/2BWq8wNQqDWuZmrVFyRajTip5quReNuzQMrMwzekTvYZ7uY4a6bdeLoKQuvc
1S9KX1FaCivEOl+5MrQm/z1jF2xFZgsX28F2M3wpcjFnBrfYC/adD1PBFl5IZq1g
qYvptTd+RxkPC46ZEt5CxHrsensYSCguu0FtDh0EVguKK/0OjXdlT8fAvp2mNNHd
2qhN6601zZY/u5vsZBMjBT0T9gpYLP+kiA1nDXs6kvHtoFKwIIym3Cr9Nx6NBZZ4
pvWMJ9i3wsrC261P5sq8A/T+6PMI8afO/fWw5SMyNyIwejlY1YU+KGaPE1LFNWsz
stapyxYU59mHlqvTRWe67W4F9zOkCozQbqu1ecr0HIfTLNbVWe24JHEMV29yMji/
1tiYmECBNuv7Q2B1KKq5TEk77F2PL7RpRd8AQfQ3gNycyUaxmrnTuEXxns8wzBdm
4ImvcEpW8c/TdSxF5RBv07CtnKcWVnPPqWcAM6dR0z7PeCFe1HuAwkhk6P4d0IXc
MYLvCU3tXsD4hJnPAePw8Q6FbYXnCeSJR0yJ6S+2jour9vuhCSqbm8EFDf/LFDRw
Ms0jCruoTehH7sEdGrwtvc0R2ab/1j6QkA3MkDFsG30fapWjPYyz3vdLvKUMQq2w
C0NsGxlAFMp+KzcyBCOP9gfOTFZJYdMpathN2oLe2lV7abKnaCywHyvFMjq4ne32
P00srBJaPu6c2AOSuB1dtG3NIpSz9PPg0ZBxMvmnbKKoFqWCrfmwmN3fJciwv9Fv
QqamWqaELVJWULRoeoQKcs0q1tEc2aQjlXvtuUpBBvYGbMWKZQmCkGrZ18Bf+R/L
lBtAR1Xe3DKUlXaD30YACtqCkrAwEGS7DvVYhf/acFUf5RVj6k+Up5rlafwIWKcc
dwavm+rELdk/VSZ6Xkt1kjbvD+iqsmNKBm1gJTCm5mqSzMio2w47GET7ymDH2yQC
jV4bBLfojc6/gLyqeTmAANz19GNLg0nVp8DzjMqkO8OPMFL3HC6Y548XhGLdM0DG
imoodOXdWE4fOE0uwn8/FuGdzbN1OSw39s2frBevhh+Ti9L+Nnu2pfxRp55N3RdO
IgscYgzvBdo5kgv2/lV+tyog1FTj/7cOzMXaSkl9ZucKT+Jr7CyxjZ25cU+tGewv
IHumo/2avFsT97e4wFaEQbkZVAI5+S9qe1JS48VoedRFEkd3AQ+ldHJ0DGZ/FaEM
zk8aA73NqiyD16YDbSigSNoj2f9PGpqHBPoVWLe9+/GqLV8s4C/aYOprKTERSt8q
a+XASbF6eDyOUDZEVnMyNOc/70u9ezXzef+T7nZ+NDaoyvByQqcHzAzL6Gjf3wFd
Drrkbgk0ZMWPJP9dJfpgo71h2C5Uc+D0Z4z7huKbysWrypT6FeQ/4IbvRemhjET8
w8kDDN3p8Ah68Kbl0fOpyfCeFszahHkI2FwJCjNjeKCr34CqT2BIt8RGgKPnfH+l
xf21gTlbRp+YbFGPeWndf+P7LlZ5LTg5GywbsxESnO9bNb/bWupSrKK0rexxLV6W
1bOyouIeHlG0VtUHcVHpQcLvnNbm/uIiv2twGkm/DE4/5kj+Jol7BlpeUWVxyuct
ddVr1yL8xpGS420Kx8lCRw7hvi4DLUM2jMDlwCtsr08baCyghJXCKZI2J3iWe3Bi
oh348c8r9C4W20Tmc416IP1h04UKr4VovC3K7Vo3kUimktNM+E1KQ6YGyLkf6+nJ
WRkccvOyr1Xo6xqR7rui7JKZMsiqs3QD3l4mwoRPJi0u8Df/TMgKKQseEJMEEio/
BZTLIryM0Gv9vwxKAWaBZOUlERucJ0oAWyy14nngEp4DuYhaG8cD7BXblFbtKXrG
hlKLMD4+Z84NXtbm81lUmqyDJxOjhXws05Nmv4ASnFH85gj/d6nebw8zeSYaygEC
Rx4Zcr4TgO5xT4yW7OZo91COWmJtKhMHxpNL5bMd/PNhVoPysfK9myh/QNv9CnCn
V4jpbrIKs85SJWak1cQcpiNPafT77t/f0L/cxTdeAf5EokKepHzv0qsJDR7MRxDy
wV1CRYZVHaTikoUlrKLYWewsYYpEStoOE8M/3AlOH/UK6MXhiMRd/lyuvraG4J9B
rMj9iGEzgWA9VAVzJHVk7cJxmNg/BZCpEtEvJFXj/ufpg3enspei97aqR61lUXjx
EDvOeZYYdO8D725F4X4kADoqHCQ4dpxrBVT7KraemIhPMdwWLFHF9AFPcIbcA/Bm
wrZb70v/RbjvUbdzF8Ry1rClHG9s7A91PyQ/ygj7XaEIDlWEDMmE0y6E5qeQJ1AF
V9KzA0/lVMhVNvW95o1J5pOz29K++RWDB1bP5UqnbQ/0dhFHf9qiSI7GnlofPwf/
Merj53kLeo2St013tm/+Ewdd5Ds2izxE0tQR7LtDEB9EFvr//OAquObwthE+O0pu
M0tEOGT/65aUJ7kHkLVb3R5PbR3oVK0lwcle40TJvX+nga0isUp4I1e4/OLxgRcO
psrN/zEpD1s5heyYLA10kje5jkAAjJOT/WYbpVNmUDNtUj2MIU22PWNpYh7Es7aM
GBS7fwchT7KDxoAUY5g/j7gLye0F4c0aeisWFh45hSmV1JgEwm/hGiBwXt9IZIoP
1cL5Ar8ryB485A4s93puaUrT/toXR3XnfqJvXXYjjhntpvIVncdBx5Vl7oF11vRR
qbMfw0odbnwACmFqFeumGQZFg0bofi++IzsZG2V7jMW6X8uPa5gYawbNPS7hGlTA
HkI1HcN3G8GrBERMFnmCWdIsH9NvLZXurVIg9xIgKXbcJR7/Z6r9qZdRodeRLiCq
ZOLx3k6NMuSfKp+ehGNVY2i+oKVVYKtOizBJk7I0lPUjTmolGe9WhLLZKEJ+aPiD
lHZ0Pc7848tV7eyQhu0Di7LUqUQcy5qAooOejJcMkg5LjM3T20KX/n6etuCgc9P6
OtSGIGRBPKjJG+1Qxm7/gFzJKcseb8ROmjh1ltrc3ucDDQf32dbsJ7JXtPOTgKTf
MHey+uWPjyZBsi3Xd2b4qr2N6DYtnFjysojEEZe88TJ+UhsgAJVojRCbi3gYgX6l
BkWn9/vdM2TagtarG3tCqmEzXHAke6D3paXI+BW4Y+nQgRi9vISo1PG0RwsKTZ/P
FBfli1glzw1DQnliI/03PeSdFLwDDfIFZpM23UQ+Fm+Ad23HxJy/nOJZiBm0S5UM
P9+AQAHLWxIkpkSlOpW68dmmnLELYJd7n1RmCVwmf7oqbUBCM1DjbETbjiRdjTyw
KjPxaFKsUm8VXDNIX1XN8NujIw+YOl5JV8sKqAtuQlusP5PdXYxbRs9PjvLo5KbU
Gr6lYy9a5gkvSCy6wNITIqEhqZAQ1w9t6PuqQOuYyu9faLN96pGUQC3ZqwRHMRQW
0C8xnpBEz44qi8yqYcsKXu0msNjA2Jkkn3ZGRv7s0HDEiS2PrqrP3lLw++13bKBj
TnjzSJAGGALPG14k66IxPx1CfsyPVXuGwUbRVshmHsDRfB1AzovGtLT5VYu3ti8j
AaVie4scVu6QI2p0EoldB94Sq1/woXdyi2tbiqjIWwZWqVHWfwPGzv0mWH2KrGb8
UPQwHEeT/QUnjEnINC1W6ZUT/OI7unykIlveU2Bfhg3FEXZEDC95A3X6lWER/VXH
mpe5tIKb1OFYhu2EK+BgJWqJQzZvwbK8aQESbPYh2Q8cnyzSL+O1ClN5sm5p3u26
nCMybn6pDXiv+KTiNEEFwv3GPQeFCoCRT5uMN40RrRNgFa55+umUKNHvEqQWlUyO
vjEzf6k923cLp3IBgvmkvMSBGeK0KQGfknWA6Wy8sX/C+Q+Suf+RDsq0tD7o0sU5
DRw2hoJ6KXZ+Xrch3NrlLOqXt0fTS7t4C0Y0PGXKk080wvBJqYMiFRCEin3t7fgD
yWF/dQ7n4lCP0+x5DM9UWsLxSTI6095CxAZlchQ6fBatsrppim7ZmlcaMMqEMPAM
auS5ggJvCTz8vEWLRast3SjG3Au9UUhu5B8bN5B/5/g5je4rezqChuIhsIkK3ScP
NsxUyo21trs1H+6nVCUzn/XlCf7aceBhrD5Tiw9ZmTlK1gI9fqZYy/ljrhYGln+v
C204h1b2z2q+2f1hymEjnhUfY5y9qYT99tVVVrXkYdB2w7tKfOgSdMSilXIuzEQU
ONujW1nG928ZEJxq4BEMwYGMa45j88J9g+c717ne+U+sXoaGBHJFWcFT0TO+pLzd
OM/OUXksvAQaIOePeh4zJjOWa3d++YjRbgeoMbQohgN4tNb2itGsMA+G+Gdmh4Sa
kXpaZGtGcEpUWcj1HsR6BwSf8kQO3T/0raKmG6Q6XbvyabKgSFYTv50k0mnwA+sN
iTa0HcKyYt5zdbCRWPtNF3JbRe5yXKKMVu0vbXX6WCL/rDBendkgVsde3R7uT8WD
ma/qC0zGAxfUWIYeQoSZpLtH6J4QWrmmwPcTQuQ1pdNmVMrm25sqjpit9xJMS5pl
BBpr8zFs6xdgAKGUn16nel+xtnELHGyeLYmzhd9x6LKNHVB9d+iZtUkYK4iD/1Pg
FCBPswvGJL5R0+JWhPTGdq3FPO8fZZn7RrvYgngH1bWl40qVd7m0tpi0Em65jvD0
aeuCIFHraWoN+4nw4wmWw7zzAGWrZy+ZADgevK3HIK5hHDTbJ0atthEcz4Ga1Twq
ZRFWJk3oImyrS+isBuyKgivdhEGsxzp5yks5wVGiwGmlzP1YBCuECkUcSNKRhNOY
fZ0L+29WeqCBvt8vdGjI/wnmEbvdff/0SrHDD8zwkB04uzrrcM3YbEpTj2t5K2P1
2BSse8Ni4YitxYuwYykMZM85y+aA5KxVBItTROx+CvmqiJylRU37E4hKtROHyqRk
WePRzfRNQLPGsU3jXHl18CNcJfETXcSUcUqz4rii55Y4xnl1kVviiSfo3J1pHiZh
YgsN9l4k1/LdUIrpdq9eUQLpYtAnIEI6uPE5DpZgu3tYzgGBK22Jeiy3AJ4uWCnt
iSAk1VPnOCDdDZS1Eqs4i68nU99picGLoT0tKINL3WtQ7VRjgg62d5878w14Dix6
Tk4gqrs434VKJG557tlQmmGF2cV0nhE7DrK/YjwziaOepdV4MBjGrnkkaiydn3YD
5D2fF7G9t3oWaog4wgFruLym6KPJkfw95iA96jOZrpgmzhSEtrOqsKAG2wi5NNi9
EaElljEZ1pd6GRjsr4DG/EMlGVtSGTB8Jj+mY/45KmFnK5bSn5G5eQHb90/xhOpK
eEeFi1Bmy6xHTehJklINZwSaCbtaTTZd+IzaACKEgeWi16nQVs6+zCsy4AYmvO6B
noZ73/5bslY0GtxLPFuZIK1oHlr7YPMXUohPHhyZh2JLSU3zQGYlzbdAryFH8WR3
T8IBS/UYb4JKFTEy9HzfE6fyt06H1HNkb9fLS9BA51ZwAQ7Bv/OMJ3Wy3oNUHkPb
tOQbzDQyQhhnBozNEM1tdUtO/Da7+SE1mUXephsF9GNds3gVa+EeU7ngDmTviEDT
C9Y59ahJp/AQeSmAWBnIZNTnrGpJ9wnElQduOctd6fOBhB/sqtdCW7vfB1kVsQ14
SYCj6fAEI461m7UySGdkwjX8OIEshc7PO/KmOoMQqRdqykGXguWk3IbkrCQYH1mM
c4T4uCt395ksIpeAf3LrO0Lb/VlBtHM4pDGOl9x9+P3SwtvfhR8/ISC0YQNEGj5L
XR4GcQxhTvWGYOpt0KriCDKa+Un/VwXDVeqSJRTBcB4UalStS5i/tFcnrlz9DltM
jcdtUlecmwaqGWZg/rqgnq6PbURP68IsEAGKe5wlCh2uSJ4BkOmJwKw61CuT7Ae3
Qt2Mm/rmsTgA9X/Du2buNLyNWWfchUg4cTZkty4QnrrMT8wTG3O9bbOlyAvPnOAt
jhhOt4xLqlPBSOrsPrymtprEoXxumiKiRY34T2rZnx4PkYphO9MIkX16GVR4cYWG
UEJdPRCVKDGyGrIaGJW5k9+TaqtaPzPYnl7bcKKwxKKBU4Po3Ne7hAgNCJ53b/cE
s4oEoV875Cza/PgLBRzqZ3k3LMJHWUNrKBgEkfT9GReHRccKNksiN+Bjfrsa7E3K
qKDNqinmtB/c6HPUfRr1zoD0b07V6W73VBnPDq4cBHiWxZeiDdr8a4r0ASScKU/+
3DGxf4+rzDyOlZfFSDB3YAvN8ZlCK445WPyEZxpFN9oeeTzai4UMiAgg2pg/OF3R
zRx1mX7pYW4PkaZ69z7GmgMGmf9IfwK6kY0+bhuPg3Mw1td27bo63cX7Fta68erg
w1l3EfW6AmXGd9bkhlFJgnJ/K2DE88SHzPVE7tN+9HoJQ84qmc2P6tpg47tlc3Du
8JH+GaXli4esD7Xb3GI7AQ5I0vn/v6bOD8mjpCjUR+TluuLENNJsoFlyBefbaSzl
nelS13NIKSUKJejoxRDmA5624VeWrPghZXRzOcuyqicHvpwH7+0h/HkY9wGzRIif
bQ2Hp686wEs4doKjSK6+uErjfyft0PEq/DYw/kfotG3VYAEKFWNXdTDgn82Uq8sF
epW98wtSNC2DEv2oBFmWfj+CK4mI+HqUiQLdRk+hxEcmuiwvFfN3htRPmnrIv+Lj
7ge2Ulors6vC9IRyDt5mYcarU2IGRRbnQ9YQ7xW/nC6lIVwiK2uhlldoW9x0d6rH
/8pNkiwyiFugOhI7HhhRbWz9XgrFc405KH1jf772k3HB8m6RESJCeYEcuViyj4WJ
waZ39xOsAjSr1aEN6ZCU9dyfi8LSJW7VfoexBrrF23Zq2rQ+OSeyAPX1FxvqxdP4
yXvknfbTBn/GDLnWwnxJtmXJ2NQsNtKmr0oeFM7Sc8o8Ae0d+b0/xR+sKKa8iJJJ
Oc0g5GZw3D5lR2scgRAQ9781gDDAnnqF3LK69CDa/VX3bEeJkejF9UOBDzxyNv0A
7t/Co/F8rC7hgnSfEWopyKKmINuhp5AF1y+weeYppRhanfIWyt+TxnJBKLLyyccn
CRVGGzvJYMu35TqzdnwIWXK7XWFzKIw8kDChxsbGeDl2lcuZ9INLV66N0j9duPM7
VsunJoNIGhBZZjLvRVeXzSCdGDQAzApyjKfozV8ipM/k81pxwGXBEqNMUQBeD1mn
5VoBhp4Syz+fXVN1t+CsQzXOKuj63XOpeVZlKAXGUvHEm9mjugw57IdCxq5mIOs+
y/1QgnWVDatI9VKlgAWF2z5cwMKB1Bne21om95OtyDxBnADH2/8+bpklFTOSoaDz
hqftd+0x4v7KmdHwbkhYEJ1cROil875xAqnu/hI0CyN5h6Y+askFjAUy++DhlVsE
K5y3dZJeHnJh4pd0EYJr1lP+NmiCqGnYxmL5OK0pNZOyX4bAL6AzTEdFUIZoulev
O4j66tfQ5H5vEUyxqbV35ns6r1sjcZWHN2+p7i5WyybNaFCdmibKNvXmBPsHJRhw
k+HH8zO+LAz9B+dr0sawTMB7h33GDgQbyQzo1KP2wqOl6K5RftrFGyhYxq2vZqNT
vYAqp7Svu9Orv8IFPHPiR5ivGL8aLsENgtCt84tb1DPVAslJCPj34eo2lBmpwJyl
zUJmG4Tip3nwOxfXuFu0k+rzMe1+fIdKCbzlTVEtjoleYgRk1E90QchriXyqLMkb
gK/yyU47qXFNCbJSGYpwW6Ov43xgt2+ThZeh7/k+vOoweo/1rk9sbZvKNrHYZbQX
5BjMuoQxIlUOb7T/eqLfW2e4pwIdDIMi2V7zM1MbJY1firwzuen8RT38+d4iNGDp
eg4G6v7XLxM3LU86kEI3lVINL7RQO1ab5M6Yc49bYYWJrZUoLYIbWjJW3PPfmvid
ibTywcezvxmdf6Iuz/Q8M08UQf3WfZqN7H5ZUdNbDfAZeIC/AnLMBMhK+aJTIuoa
XviELb2/4jYNa5lS8oHd5JmQ5rQC2kwQ81uO8Qa01D+HiS6+nV/61XqApuqJFrgW
NxRuUAj45eUzBtSKWprde/7rp+Rd38e/zaROKKoA0u8uCCN2V7RF8fX6TxVS11F8
k2QMtASwGNAo2EYHFJ11RuIXHsOZbpMUU88asZKni6w/tiyOC+8FQwzwKYzeInpf
iZ07xEYvbmZeHb1doO/6mEHuEXabzh4DMpJ0yQGYwr6+IcYhG4F+cucCGXhs599C
mknnHhgSIBYl//XYt0mSJzE57Zf/Ry5V9aCkI5yVHxG2uzozDIuvYpYO7r9S6kvO
GrYYg7f86tnISA9mI2jeNXt9dsLTkPwPGKL+reFqKOouB2GdeELETw1dKsChVtaW
snjZJLZDY+Pi0Btmg4+7GQQHFAdGOpiQamjFhweA/wTtEuSbaDYKZ8b/FkewPLUx
egxlR3LfxF8zWfYGjR9ViECwfUcz/B+cZbpe+zc7EmjyEDzr8Dtt7OPVvMNsASDO
aKo/ouPZc7jtp0K6g8dLXVQzaETkKSRFDqGP5vQ/KonVeLJ9/QxjB5edqHNPKY5I
WC0kJCBfKslSX69ibbve9gzr5HIcYUWP25I8k9jcgTtt8pyix4oOwXAKnIaZChK5
h6EPmS+HkACwG0wtA3XZ2AsTXHSEIPjUuEVuyRPwMVJBsLCKmWSg1HIvtEcbp2aY
nUlSN5PvRO0x3/GjO/cAXP6QOqJtjPk7ilQ1r10Gaa6Mc/UQUBWgeaj5b0uddBzN
9X0QksJ/6KvbhbLcIrKwKdrcAR96fbK2YR8phHTSgDA0+UBqzMxsRhjHjNtEvAzS
2xblFaqJ2lojxMMuvXhfIP9Q0IeHy8fEC+xmS1DHbpZPkVIwWz0LsIaLXr9uowl4
2vCcPokFTLPGJkFs7cuYqKe4BH/jqflP7Zt1zYuI3O9lpgVHhR4ootqZs/bjKNU0
0arm0o0nTl86RnxhvUsMlVoW2HU3ybTGtuXFtlC8fFeJTffOryKj0rBJ0gV1l7Z1
lfcFI/xjORsQv5E+jq8+QnIrXFsFbF7LxhsrSVCrX+f0EL/dTX5hojiyZqXqBX6+
cvu7biMJ2GWxtZ561Yw1LKzE0BmC7qQ5ILbLByFug8hcpiX0hPSU8oiGNUvLyQa0
7qUuBpHFKc25qxySlacGSt6YiKqA0Q3TuDDfhtDCC8aC2v3gaGtrvUr5Rp96O9Ne
C0AF/ib4s+/TJBsdqRmwkcrturLmzuIiN8gBjXGVb54kq7b1keKiQgGgD1P6Nghb
Y4cGudwDqtX51TyPU/zvgLwOTBSVHIqXdlPCWxn5e++nN0yGf8snQ/D20638K0KO
HQ6rmePow3s6yVxo693tkDgUmmVM1SAo3ECUcuxFob5C/WfCsHoZvMFG55QRROEw
KOFYnxtB9oHs9EtqZJosSfkXKmsXf69KmpDITX0ObAPo650A33N/wzYzmUunEY/Z
EHOiDpciznnEB0BMW3lLLOfTGqMJIP1u37WSw0uHB/zbxb1eDWnvUU9ke2Sv6OWp
LLt619huljssRrS7kdNtyWrbKXWeYaqFAOYLUcVZy2z36AMhl4vD1sJnWPxSOhZb
DaNdJ2r2xQQ7d2mVW2wQVVelpSHWhXNeLDDeZCzFg9TmH882IGHiHJM/aUkSWWkl
HZUzQK6XU9duCvWZI+I1nDO5xImDLrpnKhcWO7lbE9z7k1hTgGsWd2Ea0CQ3EQRO
Z2B/FwE6/r3ph3WDrJ+V1BSNYcE+QIZcJOGg97Ojxxm17l7aU/bWqW7rGNDkg3ix
XgwOT+VR/5+PAeebcPGcEjKWt3dpUCwwbldWJzFc3YVg4UFKxZ8FSt3oG77srDPl
SyJkta04bctaIsfLFzsRUGmqUGUVkLAfTFKQabK603dcxhb6vDWzcmrYhrUN1a7Y
kghtXL5kY/IcpCxopeiM1U5zT4ePAQDlZ8nbuT0C8FSwVGKU2PHlLJAQe1xhQcaf
t2vcnMx9f4/UvDfgt/9I5eHsO4l/A0tngWcnEb7I5HQEN97SI1sA9CWa3oI/OaoF
b3bpySh6z3+/t6f06hDuYQbRRrFB6a/shbmWALTYQHgf8WEAMoP4uqa9uOCT4DLJ
hP7HPJ/LMJ3vcbICbjdgvzV0QxQyeota3TignsCr1shGeiYj+lHAmVsjs9XW11Qd
ESo4KCRgg9dZoj4gTvajKh+TSZPASOK9Um+T+HRyES5m/Z/m+LmDQIiGuPxRhSyI
yacqTNvOLw780g53wxO207zkKWbpS0MFkIeFP1B2E+1BedblUTWteHdO8cfv/aP3
RhzWy4PFyL8BeM5L4/iiEYdg8LeQ8CX9SfGp1CG9QTz5590tCT4N7oDwtLGbOHb+
OquCVfS6afA/YYt14rliVGhcUHGdvhNMJzaW749wGOa/kStLE7OF9MLds/Rg8ut9
oqb10xx6pNrS1i/exhTZxpGGKcfzOnyUTpp5IwQ3zS/eLJBMn4DhWsdTyVBT5t+o
MrJoazMbQjXYndxkIAPIpy1Hg4DufqYZ9qtlAq/hTsc7Gf52wHOl0tekgX6NhHeQ
+Lsh/uQ149fawIrrtPoEUTpsQ5BLuG8nbZN4BVKSkSJBrCw656sSn2jyscqTWtKx
xigTT9U4oj9DohACtVDPogbEsaYhbhsUL2FAKTVD4MxOZ3SMV+0vgfW062jvg0ux
u/Hn1FvD2jvypAyHVRb4KOa+PQlL0GAnEEdrz2sUNbtYc9o5WKOQoLDkaUN2bu+u
CORgIJ6qpO5HZMyaIEneAfZeX2098mPP7h1ChxBU2j1IJlh+WZVCmATSHP8RF4Vq
XqFowVJHxkifjyBR2RkKQu5f10Jyxc+JItz3t2dNluuL+5uAv0ItIIfC4ffyrbPG
btQcDn2Xxl5Rzb1xo9HxICW5JCkoit1pjFHO6xh/wmcAJ0PvywxURYWKYcF8fqVl
2bAassGTHNK4fOmrK6p43UNsZ08amWC88rI9qzGLGq8E4d34kXJiDzWTOpmffD/4
VTrdWzZmlkEcPwxOFbcN53q67S8JTmRFpv0u0wMHiPyJ+VyvxN/YCYBwa3NTwyxE
OH3yuZj26EJH+M4duzffC/d2aObwYMhPXZydMTRmVhOf8x0+JRGb2CQ4Ur9pLHP6
c/LOIfvQTh1s+ECBL0sgPcJsPLswKdHbjVnu+REF6TvQfTslxnRvitN3KulAO9UV
SLT0gXuJQY7N7S+kflUe9Y/g3cE0g7uzNuSgLNaZ0o/jryTzYQgW1Z3R4wxnQ278
b5PKb3L4qU9gILETI6JfqA07mLokzJuLkXW9EjW9LddfTcmVfAtPkaw/s4jy4aYg
z8PPCEBgWqngOGZ9Pu76LAuUdtaHY4dakdmvqeMFT0AwQr6hD8bJ4XRo/5RTce/g
uow+G/aOWZV7mP6Gf8E2ObIOwRNGQ2toCMPYrddzacLZW7rTeYhwtN6xJuRBhrOV
co8vedY0qKd4F6U2mdY2M/hjtj9MRmOskFQ0HTEIfJzBs+NDKDzQnRTV2Od4CzR6
BaWuxpA9wREFa9h8POf1Hpl638lP46IzNkscG3qsmcQAW7+eRhJiUazX3EgS0JWD
PaygXPQbtztHFF4C29u08QMH1fUQD9kit7ft/Pf17G9AI78oPooOiRq2AINedGci
4bB2xp5+7Wm1DYeXYFUAp3q6FHk0JLQIFtsOjrLmfz0MSkej7TxBmce4PN2gFFvd
BLN7l53Grz7BINZeeKBR9k+SG/MLSjQ7ZdkbSUUr9pOiZadp6KbRgBKF7nM4b6uY
UQZZae6wA1QJDjj4DbvTyUqXJxVKhIRO6WBd5lI70xcrz2mVsPiFkzN1m7rVd5dF
MTkWzgHemgRONjgwC5YQ5l0qRIIl2xMzfzOPp3MHNKui1oAW4fSYa7o+OmpaeM61
mOLGX0vCVOLGbpZ3oxZgCQtPhNCu8/YnW8juBFlvS9TshPvdDs7vD4qpFcy0d3av
82eWasPZ2m19tf86V7aZ5AAHE1V3GDnbSw9mYO6kErXFKsKJQk+pE8Y+cVrDLLA9
JPxfqNEEBtPMQa4JRA/RW+E/kiSIZknDs7iJ+N8femVUUssTperPtE2xrvxVDO/0
/VIdDwCzuMjYt5Z5itNv58Y4781C6fqJ5z+dxR+/OWIDltyKhXlyD9LNZcbIixly
8oJPzrg3MCsrIF1UvBaYVt7LMJkn5JUlvRUxutwWCdZsIb/rlnt5PI9OdZ9M4wNM
5aSvAk46FBt0kOcgaL4m2JZQv8M6XUsqZUDrDRozcH0RyAsZAYmFi82sGsjFeNAh
6rUwIyQ8+98tLwHQQDhzwEiAwpJTxgLVu3xM9R38aYws0Dvx7t+//1gAJ4aRFB/W
8zf10WFbSewfq5ejMezwQF4xhgszPd1IHga/7uuT85jCliyHJbdqZ+YZOtaPeTO0
Zdmpy6wr1Xko7xR3mjb2zoMXSc8L+OAYksxwgCbzeesrzjzQc7pyxVkaQjP6AcuW
U6OjYGuZ8XRf5ZbE5JTyTNl8Dc/0LmRiZhawQv3cAiohxzkl3mSUZOGm4JzjzoVd
U+Yp48rdW6xT7PYtBg9v+ipSGmNzfUXB816WbXWzOKfQDrQmW4UiBKxjpKgjhE21
3Kv9N8hgzgniMcX9tqT/JtPSt0fG4heN56vx4lQzGdF3x6Aa6Tt+idzAvxTSSSmD
xpZkiOJBEeOTwiITjrJzKr3QJSWUrv5qr84HMsWzUJLTa3WRIj4hq3aaeeYCw20C
B2XamDOGg3oop1zoNBXkHcoq8Q4SMmIJ8Z4BCgwnjgPMtJw4M834zR7zCNN5UEEb
Lk21BfIFu9SVrxaSNrVMWladIOIww9AoLBJu0ouLA12ncqwy1x+xPENxSkwciexD
AZPeKoe2lNDLlBxRa5eM3YqB5rdP2IJWm0KS9jUKYd9zU5iOHp8Kq2MmGXiwaISh
N/XLxLiO7lUg0bSPlP3nYRlFHpAuYa/hj4Qb5dUZOFGsYJNIAXyuNWGbdQmS6pEW
f5/PstpMv2RaKBhBZgGUiY2yYbG9vcVmeNQvuI3qG9M7+RBHOMwV5GbaHR637ZS3
0GFLYtsuQ9P4Vr6AXmC/bSc8eH/05ig0o8XWmOcoEBlQwa4mlPp2EhhgdMyUmyZE
oopMw22j05fEeu/y6KLm8GVQgHdFpnNYOGPpM0TZoJF3EgB4Q6NbBPKSosATe9rH
E8uO9jrcecpbKfVe/RMC5bHQ5nifYXv/zlYuZUg3SMAdp5JpbuNfng8EKeh4ThHx
rtoBASd7ZC7SGuPLrKYpAKDbkgEk8bINhE+Plb6F/SunlzycTPUPxo3mloqU0QHe
jEWYg56J3KgRaumkUdah1jMHFDrjLlixeAOiRCq2l3Q5xajB5JKpZomPSNhCDKwJ
jhNPbKAA+r23uaKvBYuNXbuFBPd4Ktkrf94BEH8I1fT+97Qn8+mWkZUENhVB89sE
jnfUdObJ0hh8OnnrPSdy9lB7j2oyUqVUBCoMLA3fg2FAIboAtxBO7qhoV0lSTVjL
kRk7uXqgeq/sTWcMm0eb8vudupzcWy0ED6WkR66jGGzWcJ+o/EvHAxMW56FeE6Kf
K2FGgglla9mi96s0vLwmfLTdO8fbGA5lN9/4ZiFFOPV/4NXSQVVg6rqgg/CGwVqn
CMz70urLb0n5vNReu4Kh+LtRStl8c8/XRXeq0wO2behzsdJQHyFSoBCY9P3H4h1K
yc+8AuVL5dp664L/Gc06E2MIhPDQTgUNuwk86z/DZLE6gD1+QrYj85bxhz4rKDK1
lVlbttlxAnOsiYMgTXa1x1hHyRV6TpGYbmfQl1haVskj4fJ+3HGdVkPgnKRkCLv5
CP9/Y1g74WD3QM9QqeEAdGWs8i1rly5B+TvhQpALNYtkUFkg6N07cJz0EjayC2fK
T9vTQPnZqsZQDhtlhIMS8VRkTDdlmhkg6uLtpbqrmHo0XKlZpXrTEs1X1yMFnYH+
dGWxdGZxQQ6V52MSFngmL3DNjJ8W2ZH210kW3ZRlLvp0iblugUs+l5gGd4Rt9qrd
U+g29CMFFLssgwH/OUriCljLwZzyjqrkKf1X45VES1JCTxe8vKdFgq6tZNsSuJ5g
BNrAJk2xjiIK3wsdLSqVlb067Hgeu7qbMMW/nyKPfKRe8bsLGFlKkwmlzZ2c1OtM
uPOaVr8v9RHWrmBdfIKd531D5ngIy6lQ0Bn7nupDy0r07hqqBV2EtbdFnsDUMun5
zGvORYyncBeqF6b1Du0OM3ung7C9jtJ+rsL+5u/5TCDpOH/OzFg9LrIYv+ouckGG
iYqXMoaKQHemjAOskeTSrzOOr1dtwASgmXR9nXVJU5t0i5KJaapgqkDoxjMtt5ga
m+K4hEBaaeg3msQd2OeRq8O5KerWloXF84wxD7O7dRNE8YG4VjNw0SFcGH5tCcm5
s7oZyQH7VefYmNtmCMXXcJtgy9tqIfXLgwXurC0ZMvzjwlZoKNDg8RMmYCyvmi29
z/AH3yyQN6HfXhBOBGl6Wkm8M+uJpKb6Rg2EVnd+jQfLLQNwgcUHpEX/xzzFFqIk
nhQ0fKjtyuEUB/BzlA5mOqoT1lEqHiq1xt8T4SxoFo3fT4YiDoogLzpbV1bwJi7h
xlBdiXqOps6JDs6QnkI3bRYD4iBGjwqbfInRCFojmV4zBh3+EhP9JcEpndmGHoF3
E5ta7625zA9R1srpNA+KZpwKqzvu9M126I5Pk9Bu0D2MNMmO/A5PQDJupovckAvp
Lz2dU6JeUXvI1ilhj+dm+9UHnqcraTVndt1gbuyTafhvRUYrIaZKWnzIHRCsrwwB
pzFC7JTngn0y73XP7G/Tk+A4njXXQUyqcVQ3FybhX1KNYmhWMOxkw5RXbBRtXYwy
uv6Ng1JSMh5B6k6fG1jBxxMvkHiGWAyT+TT8tPsPddeOVpbV6mFwiZs9Nxk1yPkT
AeC/7kfuCbXDapKHmcZoxEqJFCG8W5F8zc0QZv5Ck6VmUUKcLrGI0VrWV9YAeTER
mLov8IUCUyTewxdhYSlw2k6y9Jom6x5Hn6ygv+fKzSIIDcvC70eBrzi1wRganJId
xCQBJ/Rqsm9rTxiK3ag2gOPIpotd3CIQffg+8lJaJQBOnrzIHrtGORXA+JycSy0Q
7shkS/IA/MvteYOoL0XOb5DJ2qhAKU8tyM80KHyE+mN17fmuqsnH0SxR2fuaWbr7
pQD66sbOW0rQSrYscqAdL19y/xybJPlskSr7QgLxopC8Eww0dorjerIWzQzLPYiB
fuujxyxNdKM37vk39eQ4v+R/gxoXA08MyCqcERG6E5FNr8G+tiGoTQcjmnMJ1cIb
Y48BL+VuK2enb43pFFfcy4mtQgdYrM9sx7JSbf2oXGbHcOR6O2O6vdGhMWpGLji5
DMlnFs2qG49M7GlNq01aiBFOmdnFmlw4Dxjcd7pqA8NiS8oqzTSVBtMdGznTp2TD
oXIvR4T7afIRcBEPp7UIkWW1gESeCq9oHdj1vFETRUcs8ACsXnqbbOlpWI9AAx0B
/hk67gPD1J43c8gFGKghVouGCQEQYvdGG1rlmjBtp3yTzgTzrGoByEgXjRhYYG5G
LYs3bU2N/yjrZ/cw/ty8MOze2+iOOHa/9vvG4+cPjvYxcZKlSVejsTZdUEco7ZUh
9yCPxDBdU46ENu90f5kgOu2No40MHeVUA1q0Yfgj4EPQBNlzsOV8TD/1aDo4iQ5r
RwVzKBvnZOtsRPTAV7dsbO0An9k62v9qV0+Xn4r/QTXnUodNCJubOIt0+LqOwthT
V4uH1cG2psISJD5xKT5Mk6SHS49t12dPBENV4segvdn2OTpRz0ffi6SJ9hb60eRC
bamR+JHGkp6mTKqD45UybEDLG4VThYpHn+04RnpysSwi7QvrLKR+8thyuu52dpjK
iJjE7onItNX4GnE2MdvDnGoPyVApT/lE/8npSPvvbVs9l7ra+WGXYbAn1RgGqyyN
LZ5rbu56Kk6MsqoMfZXpuJr9amV/REk6DZEkjbuvnfhAgGNmtjL7e8DouB26oXjX
i2cZER32DrZinDSfg5WGKysfCjoA9mukcHYnkfVbIx0lSMUrVDgJWYxAWNnObLGN
IN3ODWZbtZIWogws4/ST5kn7iX6Evt4skkF08lhg4o8aayc3jo/UHVi44xqyn1SX
tTJobS/OZQNUI38etXWGjTgTCDVSQUpXGOB8B02QvmBqVwCkXhuDMg5F7i4zk9n7
Z9C+JUZLBVlLMEZZZ4gWZ4JKlwgAR4YRKtybc11xboskxrKXxhxsglzGBsky1mRL
XlmwZuMfkbVYHSUa0ymyBwEguUmV2hpzk2uZ6xLm3INm1mkrMLDGwnBVG+hdKO9p
jf7GSwyLYfdGx1G2SNL6mQja/XPLzPW3kR6c0cGfkoQtVQCKhUOeQXMU9jo4Ftlk
MQBCGO6EqNl5aYGm5KrGvy+r7jJfEgFGlXMkRtR48JDzCkbVp5rrCd23W/UbJ5fZ
tE6YW0rFYwM211HAPxqP5+guyZiZwTbDFijrIweEHp8LsQvqE4o+r6SsNuom2QcO
Wnp3XUTt7fWYb473nWAO+GPAY3mZVSu76oU9j6p5ldZMmXZvDlnPu7f90nV+5xiw
6KX3yyu1fz6D8XyEnjiQXF6h+nnkyZ2YHXHZ4sws0hEdViixypx62wOBEArBuL5s
nbatooBOt4ZxHIXnvO6dKDyt09LoveSYL8HwFgysubsx2I1bSW9u9JUvYIFAKu8c
WHETtUYc6ZsS/Sv2P6KmhUMfNclGv20mqChV/k+IaKln60f6VCTUaZqk4LBLhWw4
rOkXLPmGsSy1opRdkZWtsEKsDaXn5uSoUK6V94wy5iPAMIseJ2fJ67I0ialD3nvH
/ywtNM3CCFQh/ldPeyOkD7a24bl8rzRopdrozmaWUmovtY182VTN4gADLD5dmDX/
VjahBv5IEXSXf10Hg+PrGhg0C7z3XDhDnvF64a9HyFV1MpNH0lkragpDdR6eGfY4
ZBO4pAmyn/RMhcwoeuP9KpwNh/MuC4lGv/iCGsX8ijlFIdxnVfmAs2iDKJmw40ks
+mEMySDWqvUnbMR0JxU4YtAuAMFwk05HOIo9X5DV5tO22vqdr5c7oNxYnBSyvZNy
7UqJ5Lt8X5fKnxfuOoRjn7oPssqsNa5YlQe0KJpGRbQfMlpn/7YUMFCE/7NP4cmC
pxAtZQvbMNs6Q4B7wIW2bwQa9N6fEYJvPI+pxIlc0mHXdwN8MYeN5QEhWNwIYI7V
vNOu0gdloRMoKnm4SyIapqgJz6pfUw6MZSSWsOxKUTfk5u+IyNhgt58T11eA+6Sw
6pixWaKZGoCpxX5s/vtuo89bmGIyuITJRgAHtm+nY6Kf2xx89vlebIbR0f5nXsLe
W0isryAh6UOnskW2YgEs9YqpKEnpCUHdNHy5HWQIYrmDgfnVl/PaVzmzzDoZlZpJ
tsSG3lKJLI1n8i9D2FrTvjlLHqWGVzHwzyVpveTY2YSHyqVYQc52SPEg3ptuPfeU
eZxLllvA7STXt8SS7fneChm+uyz1L5QWQY2XgHUGQzeDaWljd8RPw1yoau5Hgijk
g026YFfYCnhXB81Zx9UVMWAgzc5UsHpG/tSXUPpoQfMCiHNNA95Qv+AiuYnT43n5
eoHban9V3pCfUfKc4/3L9FAiGRuzW8pvf6d7Oy0C1OLWT7PWBZn1jcJ/mzQHvgfA
0W20NlkF6rhesziYcqjiCdb7HJYJXN+aZQmOgTCHO3BV+X33OXVFM/bkK0vk+mAJ
gMiKpGpmT43hMjy6p/VxNCi5fbQCRFUWdilmqe/WUGRALZUjct0azxqR1QCAupgW
bzflUaBZfAjHd5J+DzU8l/IQzR7xqZEop3dBIP4aZ0Km4qWDXxfJJULRoVSBuovL
sTZNmJmHbZGddXISQJVZrGiAaVExtxhv+/6/3wVDr4eBRktfMlcQNnTTdcOjJ7fl
Xr90jQrunHzSDI+OrcWkhZhOrfjE8UiIE5FZjKzyXnMfS9TjMtlODOrJTqGOBofc
9nQe64upVQuWcCZy5cgsdvev/R5smaHvIT0hoTVTkOdeHK7FbTr41L6Gl5jRWU09
Wm1bos6OVuuiW594oJgU6gzPIONuYKXgICHyptHARcqHYspNAQypps8ERg1iDDKD
Rq3c40hlKpQ8sYR0Irsi5xtbm7GC+7zb/ViMdFpQ6+68uxj6C121KP1A5BkOVe4Z
ysU7bzpCGXjottU7lGJPg3hvVQV78uC9cPjU1W138MFKnVmG0/06eWx/IA657YAL
Yayv6DdgVJlBseUKZRHd6pL9xGzyfsQ1aFovgyJUzno9w/F3MmtaZu67mn9o3EvC
Vrjo09By01wzsI2E3pWpbPPiRhuB/LhcdPQf6tvIKWWWCpeqBGISxVNx3FzHpGiP
LN+XH0C1dXB8v2/uy00cT2P2wgdloe2S3E8PD+aLm2LmsHVIc3eLNWGPw2Pl20lE
P1S0T7YqTE3bUXfNhroUq2o4mYHnHyNRe/CvT9w7NdLfDftZA0XkFBQHDQjbIZGC
Af5GRKvMP+o3kSWnuYkNnSwLG3P9xgRAMzheVm992f13P2YgDI6XxNVpjjnR43JC
Z0u/7BKkwXUZ84kFFeDOPrgX3Nr7pA9WLJcj3GUNJzgZLDznv4SU4lpJEohz9JIf
Yen0cP5zrIuanvKbZ0lo6J1BfaUUqTZc6pEHLXnmu8oKDSxVnln5pLC4v8+JUoPe
oAZNPZ6jhie9M05DhFzmjk5oTNRwChLt0eKkbbWaMJ0jOPvhU5AEtpSPutdAbGet
Po1+HnhpfYI6Vbf6nzNY2/CjInQjcFvMbnvTbWXPIKznUFF7BPS5FhM5OvGxKxV/
GKlel7p7nZxq1WEEs0j9v2VHIbtg5/MDqFbXSfYHFb5dMOKKZJl3n1ndWk3IFUnM
FQ10N7k13mpqbBZ0RVcynMZzemnQEIXJIxvwzR0It9o4Ly+b6u6FmoOcUzzMMjNi
fTEWnXO8Hy7HkZwLBbhMec6gx28FDg8ZRJAdWUcet58A9CP/WmUrpQ2Qjpsqz/pS
MATJwtswUZoSZLb2K+6vcK4iyYw1Pot593hEj21LpPJvVpOyQ5O/FIHr9Fcj0UNa
F3XjlMrlcYRn3XJ/HYRjQtG9gzKXp3FyXcMt7v6G1FJaaDpM6drB3Ym48NDejZxH
LhCT9WD86aEwYRxN1zHnF+EIKEoQwDj5FzjLmVam+RLHqgnXs7mxfDFPN9Y3ijom
OIvKEeMY4K2GK9HgypB9x5Iq6EXIDuogyZf2DdzEVdtqdmZ/UIiRZC6rVEr0Fslb
5/M0EnSfkd+O8lF+puy16BGonV3YaG2KjEbDp86ADjRRloQvlq+43l34x0Wri3n9
YpC0PCMDr2f4KfHOjJHEanK7poEpfzMMFtI2WXseR+W5zVNDlUN2RAkc2MdK9JZX
yh+pUVmbjPfQubXMlGB+zoCrdHtncS2mep3x37Dui96pEYf74Z1kSgVk1iunqD20
UxMX+3FmiKZzuyXDwBEpsUJaJ6NEvDpTJamLCyifykZwkqF9vvyAC7Jca8TIz6YB
3R/749vXyhMP3ueT3tQhaSed0NJ43nXaLNscCpWpmj7QE7n/4SRvbDHijMnhBtjs
coIyAKWeg1hmCHCmgIaDKOmnfX4hE9Nzhalu47E+hvah/gFH7J/V922e/m4J1JzB
1rEqPpy01P1a7iQAo5VJRQxxWkYbHG1ZucfjIAyP7W5hupYEWuQLCYxhOHLYe3pF
/TiLzBH9IYZKIAqONnlLw1trk7yVuNfa+siq+7x7L0KZv0WW4Tp6ExFM2IbIR6ib
Kuvahv58ZiD7s/SpOPDhYAqhNdhF3ef5AD/oLCH9h0lMBE+zu0umFPC9PX6skcH6
TI1yIWSTWCH00WrlJhKTtP3y1Ja+qNwthCwMQxIHqFEiiLHhZ0QfHQDQPbIo8kS/
6QYOdw3JFMaIpvPDF09IgUeRWVjryjO8/GU18ExoePIwSSIlCo0rOIN8qsXrPvFX
ftLq4krvwT4Z7od52SR/6+B9quMN4BuEVlDxAaA/P/yV++wbCZShDURaGx/2CoiB
vpTs2lCadTwQ5+ZqQlvKfj9Yb1i9xswk89l0aMHzIfzplNgrlN5FnZoIcjmUV5RL
Uiq+dfxyYAqnz1FPFlPq3i1qqKZnmqyk7btTuyBmfe6TK6Owp5Bpbw31zV0EYDYh
lrSZzBf2eio/OtRBa0M+lV8i543h6qsDQPdu1On3RyX29N3xbnMU3ERXlhf8WtAp
F10JPPS+Wf/YxP1ltgDS9vRsRNn1OMEDMOGU/COHhSiTW4R20aV+l1oU7T7Rkhj7
LA2gMxSSy/3lORxTLFbSjFrJd+rjqLqgjRNxoV+9PYmr8mLdygWTc2sItEpkopnu
2D4aeRW6L6loxhBhSzc7ihct43j8mkLo8I0kWuR/udPYSiZdzlF5FK7iQpwA8Njc
Tv3PZsWKiXeBvf+wYaFLhqzbnevH7TYOeHdLMFp+Hz9FTIT4wZMkPmXAAbsnyjCx
THMTtEbnsjVs05+qYXyk2PY9BxLt898C4Fo3f9u2VFQf6gvyXioZ4SIpA9EfjuH+
stW1BDgbQ7BD1Y6F1lxGFqOZWfAXHLPHNrmGgW9ywk1qlMIya3yWMBq6r9cA+SZU
E7hRlNpLMUx8qS4GhLM9SzlN8Yr7m8YqbqlhLc3TieSbsTfUeujntCHznBflo9d1
admpOo13GOQmj3OkxxsbWXMF+wSZE0wvQJcAxzeV+qhV0HlxpQssxiPAnCnkWGQ5
h7sAE9boig6Jt5vHZcQqNGcNe4TBlSr23Cl0Fy0VZu6bGeuUwdEaPQJWxkSX+Una
zIhC5cKu6KLjaSjOu1xLbJstO6CCUZViTYbE02dKQpnhUOIjkx9t8MAYTTvA1k4J
4qEnHaC9FMFvmOi9bJYprQm2cT9FLfLdS5eiH2zVb3Zcn5Mi4NJ7gO19DJW3VKet
fFtlWzWV0UZUr8Dd9OzJ6H09JsJfsnJ52j62jrAwJ5S81W8s5WIswu2KzJ91F9UW
4pjo/yZhkse2CTSPTRVUIa3uCoYWhSyhuZOuGi9J/MWGG2YZyHkNoD6ocRgFhuZw
CzoW5fHWbW8CiiB+JKfcOLjZSY8sANQiKZCetFZdb0RC+fR/TQLlTd8Xc4Yijuq+
Hp35p1l1bApBpQp24/PElOSe/HJk9NLavFukBHhDH/9mICdjvlAV2XiIebIzIO08
c1WXn+cxC/kD6rwIkCWTbnaNGOsiiMWIk0v3wqw3o5tuh5SUmc2omy0RwWcNh98z
7effEPlehIBlirW6tYRrAWBQspti448PZakFtbm0Jj49kNhby238qj+MJg4cI5Dm
nR7KTKmR/FR6S45qzx2lw0l5EROHOq/CGcFmygf3W7KWOi24OeuIA36PYUqr1ugd
9C2u3mMove0OHssNmEOYxNcsd043QAweb44AfuKHQb+zAT3p8Fmw6EDtSsmVfmR/
8v5GNz2Rotq8Dx/tIVJneojeLfUDD9AjvOcyPcv9B12e2lqgQm6NAqZh9cYaPiZA
97ro+2tsHPIdSDit7UBntz8Wh4F6lokOs8RvMqgtXYbPY4lFeamYx1SNPtHLkV6L
3rn4r72/TEjhXBbykFfCFh1RMCKRw3DMXJGUMBbdlWBmSSFKB1hC4bPNbdhcfd1h
SuINAZ+qU/3a7ppqCtMpjAVqzr0oLFTusW2m0x/jOrdb6V4R7WO/X3ghH7/8sryf
oTBIOUOQIklUMpirVh/5u51On+6DOYUV/cCuZbBuvsK6eAeR6hgpnqXc7bNIOA2a
CShyZ8xYpLYWD1NLkyLGW95LIAjIyZxzAVUqfj3/VxPY1ThBtdpthETaa4d3iPVd
3YF4u9lQiUdZ4uAaF5wPkSjufPsn4CxfxSXoHrpepoW5o+JmixFI1egfuaWuVQcu
cr//zMOVcJE/LgxmFCqVBf3yUjNDwCeNG0KIdymH8gPluJ58UL1RHmvvuMlBDH0i
oAd7yd2i3xxpDx5GLQkdhSWYs1fOufGyi91a+dBlqEDOva817X0BFKkGWKuszmWS
odlqyjIYwd3F9UhhBBOW3xJIkiROzO/N9REcIrssNR/eDzlHdne9k66GGxf16Vzj
jiCTJg7KgwHkkdvQ5wduJHFOMl9EmwnnPyTreFdbIJ1tR72sPEMWbHWzdlkf5nNV
TJYaEepWYcbTRMJLQtJFABgyICkTX9s+DzPaove6210Wgk0a0ln7Qw/1jf5En6n1
1NtObRtw2eITOMLGnqSN1Y+nZi/SrGLkvSVCRaWU+mmzko7DzSokJdQPllradk1X
DEc5btnciyepglZJ3EOY9rOsi9ilzN4G84i6eyaFRvXwbUnr8GTYnrGa+v4waPIj
fMSoVlDa+loIcPf7Gf3Sb9Si0EcBu1Z+yQZdg0/pyKSYk1952tGZrfI48mPZ38X4
fC6V8t5fRlfsmCRRivV/QhEg/0OpfODO92aJForKOa3infRQjnAr+gr2NjYQyAF9
q4t/vN4mdgAvWXBhXAdXiFEsvlK8bRqrsHgHYD0P/tYZ/oIU2Tm5kxqf4uAlFFFH
huQ3khm+S+G00TXunLiQJ0KPiMKWALWnaiKqz30x/YVXrXeg7HS2XZgkFTJ4pUgX
UqadbSmfsaOYjmycstIilCyFxRAXRj2/0pZcsLYEXDybj3eRvQfnJ3rG9qoRS5pp
TFmZOMkQgmyEXdTq9BfFMa70VjfHry2teZhscbCihwYv21ThEZvwLwXYkhtivJD7
yFYDTddA0mbuxJxjTXeI5MGjds9EUa+qckqOS5V/MnvjLL8f2iVqDZ5TuC85Dqik
ZC0tQLCrMEITJR3wOGGAtzezL5HgX/6NhJxF9/BU2g1ALcJdgwVZxMrJVdvZtHUI
SdfoWNEIqYHxInZAMtl7kTIJFzt7PChPlIUUvI61rVX8H1sNE9KMpjk1Dfmm9IKx
++ighc1tEjP5IDc5PNFEuND1LHbfaprbqyBxVBQYqnoggiU1kEqw6Vsk7PVvw9P1
FpUxqky236gr3i/aLhTeQ5ORWaPaH9k+4xeO0mWsQjIGD138KlqtWyvld13/ZTnb
l/JNUQmgQQ/qKDQbU8sOIxxt7+FoXGEVEXCmOmrCnwR+c1qKKyy6gj09OcUrlVNW
7vWyPS9yXaGecgehW7MFFWjg4iuNyXG7OLkg7zEnk/zaYz73amcNGMEEHtECgINM
30xyK5JG7Ft21D2USqXSP7kTV+9LlJpD8geRSSJt8C/WaZA5JMeIEZ55DLQyjIdZ
EDQgiozlKAkORmaOijzfl7nbC3aiFiGSkoHde/sx2B4aamJgWvqiEpRqmSFILHLs
uOxvCfpdE53qhLS0UEyvP/hdLQA5vNRfN5ZJLlBZHXqoT5KLQIAiJYZXCq987AIS
e7sMRKE02zUPyNC4BGPR1alKrUu9j7F9H1SRh7RJbRF5oVUmwI83JVeC1utXnE6J
Si+BhmCgUWP/TP5aMtsj69wN3hEyYMKbaU6C88CJUtJOHEUkFVNZ0zRZabgFLLYu
Hh7PvIS9nCxWgorv87fdWEzqeFUN99J7afiXo2MJFsNuG51gTenO1fQ4Nx/0ta7i
xsnaOe2oyhnhmQ2sl+ZNREpvX12UPLCouVJJKgVRYt9QrJaAjr1k+ZDDMnoIo+QT
LTO2NjQUyXTecE2MwdXA6TH/S3ELnaywtf+Gev08GtcbgLQOkGvrXwFt/nQ9D6XJ
1/52ECSWGwdqg0EGE/9pX7RGaVpTF8uNlDs/ZEin5TyCer3Ku5W11ZufSIJVCkhI
jqOL9M0s3NZFf0Tuj50SpYx4Xs2A5EFkJrDvwIdgWeeO55yU7kTs3VFyxcNBo9L1
8XwoWxHuo9u9+jrF8j5sVInkOX/0D6eRcykEpAaGwZTIMEglz3YZ108y4N6cOBDC
/uxshRsljF28cve1E81Q8KgPjELr30Jk81blWlcWibyp3PaSRe8INfOj3E1qA85P
st0i2f5agf69zjzwoSXQi9Rm13iMjMD6sFHzVRw66GbGEMQfXCLiy9kf57+JyF0E
oFNa2xuf70v1zpmMRVw9wNINnvEtUvRn3gQaV5g68Jp315CWTGt+JmBWCQ5spxtU
fC/YyCVI25dE16sVNRDbtiQYCqzFJEN5xZdy4IOS5MYFPdjg2I65kDMAQ85py+T6
sDLwvZdnv2AQJ+VMu/kE+qmj32nyhAal7U3RCGfG2Xl00stARiJwKqssaL894b+W
UlSrR7xyJpKVP2knoCQ//E/IimsRkyy9yE5yEOqOARfju4QUlZ71DWID6x+3ozmp
yAbopxEwP1+OBPmMAtMQ9pN55vcmDgxXaa3Sw7pEnMHqB5daTt6wuTGtxRbIItw8
E9rnsfspBBr1vV0rWgA25gzNEUCfwqshj0WCVQdYT629si6F/2KRKPdiKctcOkFg
OPCih2Q5MNz6DVtx38zKqBtUAn9BlE3YXdjdA+hyUY4/rK4yxDaCAoFT2m+gnMHj
uGTThtQ5XfmKdnZ8/eglDsA7Q+RTZNHxqL7QuSs9HjVb+lGc5+TcqjdaRk5ZdI1m
f4ngHgX2of4tVix1j2R7sCFcytLA20gn9fWVeCnpmebSaUR0dQOAJIp/EqRpsCd2
0Ujkqnm8rpnG1wjrT3kT0b8cMdzqEumpMFo2o78n/xwDCR3bBTXsysAqo+urEG1I
NoJzAgRV7q+4xD4iJUD0pm5oJIRk4+ICDReOwyuY1Meb8IrNQVpZkM57AnU17klZ
WiEmTHkCo5I+TpBl2m0mQS5wI2MDzKzEbGd+VI9nY6lUInJzg4V7ZTtADFrQ0g2o
FFgDYlSsJqOT9dfuyCBKynK06GQfbVRYiepLEo6DUHInNsFV0qSqM9KWeZoQ9GBz
Z2U58JdcM63dq9xlwhgadH7WyznpSqRKp1WWXv0CQgbVgb++mObep/+QoIAOKhiX
VGFeJ1+xeQ2qoZxKVMtm6BifSJi+4Jh8BMdBPHwc2W6hUghLub0JolVYg/0R1q1q
BBiYM5oIUrZZc2x2NPt/M1LYYz/Vyt8XeqJDMt/3YHNtlMgYpxMfLv9U9GzOlxMN
WugdvAGlW3sokiUmcLCf5OWOm0Ddc5xpO9VxvPml9Q3GXGWUb2OfbUMAsZ6unWih
/nl4W6thyTxovgDdKT+f7EHG9r27F/Ufz0cpMqpUeDQ87Gv37OQGg2kKC5ipjhny
UVdv9kIIrqLqvmOwrenP2lEsSRLLondFwjcCJYFK9jie3mo7tCVcaHeTRiUeY4BD
xwJyr16HNW3DYyxOKtrOAi7GW8LLF4BloNkaMXjS0z2PMIm2pBUS7xLdEZCfIm0m
+H9cWhT6bJ9nFUYiCOY+FQR7hbEOkSBsJKeMfQfHCqMqItMsJTfaCvNiqJr9j1Bw
o5f0OfhdA0VVN4x4jf/jLrABb4c4gFkYwq2+IixF0AEEbZ+aIgtXVPxb4Qsku2tP
KhOQh8OSKfB4NC+4cjewJlKDOmLauLICrhn+5HlPXeTlnM7jqEWr9/td6dOP5MVE
uJiDzUnHqocFkQK+g0GIr6hAuFH/UWAGBkQlI7G/M9zX0zYMfdiLg2sPju3YITlF
hDB2KKR5gKA+dNgHIm/hibmBNkObiYNpM56MbRfI/v/dLdjL+H9RhfSyhVdpC07T
53lbSy4f8z+JTjrlf/avttlWKmyrD5RK/Tl5tQU6tubq7OQ/yEUkRBxVIs7OkOfY
eWGi3cRdsYWVMNM4rlTTo31n8Y1oRwmaMbfOxMLT4RKLiq7Gw4Gvo/B4MLTQYaJZ
4zy4naXE65OqJXViu9dfUgQvDywJ9bHj38dG0nd0EinF6smZ3qCa1cNQPd42JcmH
8qirw3Y2F++dFFUl6IEUQrZX3NvyxsJtS9kAJnyz7rXXVH9YpsA97Z7n1lzagua4
qsMIP/PyMi7mbzw3FNs7ae/kwDmqjuwzI1G033LIwCOSFcMETU3gCo0mvdljhrD4
5wK4a08F8LyCQnkvoF5YFgjeCC9aILoidCzcjkuuiM1tGKjCSbK12rLXl3Dn6qBZ
TA05LdhSU0wz5cGMY6wuFiwtpxhFJStkVT7stz04XLQXUGgMuoRvUmQXGJdSpkid
civ3cPsGf4C3cyU9xHgROqeDYSu7LzJUeHYqK07+4gW7q4t0aFIDgPEW39y4EnIZ
WglH8cOmWOQmPQc/mryL7t1/gcOnJwUJbTI349yrDseWsDQm4p+OkMXzzT0YVbB4
/6Xix4JXuFjWk8pvRIponNd3G3rL+EMWEVN9AKNZwtmzgoj17lfQj+/eNw6koINI
XlXdk3jzVClyTsdHXshopkNv4j6s0AmzyuV71QyX+xenGzPDFFkNHlwXpwj7PPJA
CH2/M1fmUCD3jl0C/m/qZ9xwWRD1zm9hsO9lunxYMjexY81bH0osWPh96tWnwa7l
b16PXPb/auMKDzDpUBiFlSA4lFMMJsgvaEA2O3mdO15+9lxIAs7u/FbYXa+mYqCH
+TtJIcWYFg5bkycKhY7eQdeRhEz7XRHxMqRtLtiBKV9uQmlTUPXmgvhbNkSYLu04
WWsKj3xzD5AM8PLAP1WQqMtz0XvWTxWTZojN8ZyvFmn2XRjTrTkBPWWD+HMfoCdS
WCbncIiu7L1vxEAuvpZCFvSQBxGsnmr9zSvhloMAd4T97Grf54iwpHsCeVja2hp0
44j815R5WGt1VkczMOIBd1EBmQ6mcXgj6gYfQG6I2A0UqXgboOqctr1fzL7A2lXH
8uF2dDt0K0DRFPYxgMOS69sdSDIOo7U+Z5nqvCtwC+d/uA6VGPX5xDgHg1Q9MaiW
5+uNOw3suEWavvvlMvENF9UIqFMVr9Hl1k14tPYAfPGhwsoDCe83rh3/jyvpS3Fp
cJuH6RcvgD6VJG9nn13kg7YLhxTsroxHoiTeyP+0vQZAAk7wwNoK+FCLr9TzfrC5
XlaYosiXd32gUq2lQPTV2rzCX/hCzAFcg8zW9xwOzIW0G99g71syO0eZFelO9QXk
6pJLUb0NwAg2tWlytqHwPbXn1Zbdgy8No+7HXgDMEO2vKZsUTprvUys7NvbRXO24
9NPPWTaz5h+mWDmZGJa8QbJlyx3SRPyNmOEGdWPaNZ8CadWqm+u+urIXH9z3jSz7
yHsaLln49kJSA4cR7SczeUyTe8x2xuPn0O8pEFXgo/QFVs7nmFFBkkT8hl6ZT5Ru
lgyBdX7RxMAZrAEu19eZwquol9ixToazJyTiNyzO2W6mZOF6YY6vOQ8vpLCkipRG
/ss9HjeayN2MyBO6Lf+TH0UXjVLVl4bvvUyZEfOAskl21Gh0HzqrUVel6+BflJAN
tIpBma0pat/1Md/Xj2l0WKbl6sht6NK3xd+P6uqFMHovRXeL7z6m82iNwqjKtnDU
T3QClqrJz52tUi1JsrNRV8LLnBjiabXhfuTRQEQZOeIdwOP8mn/AZ7F51LUcLmXR
S94KmQ2f7wPrPz3aBIPZRQk1isYqDBLARhxqs4bnoX75Zo3q3eEcIV6lrhYoCvlD
pIalc4nAgrcePGi/kLBIUnjAKSsKsEJVqOqmIvExXL7cah3wOVLm2dSYOaEI6fia
nh/Gv96m9EQHJwKFzanyBPHadgSzHmmIW9W+dSAGP7Sbhky7xW3q2aVXTYkqb2BY
Z4HNIHYvatjQK+geImVuQDPM//85HjxkYvJTCpItPRV23GZTTzDFctnFB1NKRG9l
aD+zE+XS3QhjmjjPIQpFjy0t+nrhNtcw5R19pZjrecWXwk7Ll+zb9hIigawRroSH
6UIncRyRVRpnDXM8evhmTADOhaipvEdRr72xQCbf+UXu2QrNBaVBH9PO9XuTEmgG
Rg6QiVja95UlzPeMU13rfhpUcAVBe/VRkz3wZ297cbEwo3w0ZdujKbt+6PIf+TIy
HJwcuTjDP85gr0GtGlxEFIUdlDQMBn4COv7V3KknIz/AU3L6M/wKZVK9IRDppM0l
0pIroa/N9OMbBAB7QD/OXV2a7lDpXMawkrLt5MwennbVOOl68vltjlBQ+0IAmKZZ
loxLbdqoNt5iM/O2UbYZlRsafcBrZtDUeoYGzCUYE5kFAgLwBSt6z5/sos+O+98A
0lNS5WeuuCoWgHOoJHcBT1n0aei93J9PHob2h4d6sNOE8jvYg9IJYjdRictPqyEL
8/Nfw/ZJzC5vbP5OySytR9vrQuKf6WWtUPGIf81Ln1nTGuCusoHbM0el5D+qETzw
Qw/Py9shGrz14gsbHLXtw7ff9LnEFVJdEmLELfDgkFZIIib3lw2V5TYcrGQ2/7zq
TNgEAnvqI8Doan9oBV24q9Ael8V/yFZPmV81zKfpVYLpS5wH3K9KfltWLDU9jPxE
pjIcYZWoXguXAdA7ueVsf1PKngjH1pubNt+8ZVOiOjkE0upeVKNfhFx+IRGLgfBn
vMuUHNwTglU774lyGfqLltiG4PJdHtOjDwKVZIT26Lt55xkcoTwR+lI1P9nPtYyW
ezNfZYJNtD2Pf2sr95WSVBdzGW9lO4KycoEOQRZdG0V4NH5s6JO5U8w2lqUH2DF4
Vyk7iWlZRvkV+esmBkt7ZqXKwbZWOAjeQ3Ok092AVeecMykYWrWVkDX+a1z2/COF
1neyHRwrF99J7NgOEgvBonh9pStUWCXWESEIvT10YlZasdIhwwYJaF/+ap9LhXPc
trYUHoldQFovZ9rKoWBtzSKjMkIgq+0RkeH5uu0LhjQwlwUJdFTXFQ/2kkrCmLgp
jiHC44RhAEvPtE9f9qrAIVnsowXhre58NpZlwccjE/HKzkJmhUU/BQ5DlHiPHZdx
M2Awwuvkhe4Hl5Lznn8PoGyVPvj9l8ZBiawTRO4hVjMY+N0BEvRcKw2AqHf1hZ/Q
yxyAfHIknISPjeSWNVki+VqTftbz9sscCRJ4aNuGB8HZC/m2+zgogScsRMYdlzCT
f7ypeCNSGu7ZCYrspAHFiHanoS0waIqR3w+GAqYQ45zsweBk2YVZI89G3WNxHOO6
h5LsARfl6TG8+hzVoqCzxht1zLjSiB5qq9M82dTD7A8moWEtQx1n5OIhsgib4XQx
TxgKTy6bgfxVN3zQRfYTnxkfTnfdnJt/CVD3boI1tUEeO32lS5x6ObCHKq9Lm+8o
Awe6OZSfY6voPWb2/etopfQ9DnqOeRWzkyjCC4kCJCFwdNWQ+fM9LGYk+QWmZffW
IaPzXFGkAO+MkELoTiJch9C5620WUpcZSS6CsZmHZEihHkCF/9R4ZWxoLXh17haL
rMnvQBbpTTy27yDdfvw+bRJP3vrKHrHhSxFaxf+Jjii9qBg92/hJbcZc79driZGY
Zt8uITJIpPeweGI57Jey416rJvi0i87nuP7++ndtRhcj0NKYgpaf+7wLartqjVOR
/gZoFfskH10hQ13OABCyDgXEVAedPkVbNEulMuDjfgHhbZsLFsLmXxe935Zvjoy3
YEs8NofLanip770BSLuB/1iIDMBQyITuBuDOYhW4MMLi3f2F1MJ5FrDJr/d8ugSI
7Z3ZyoMQHGQX0+MgC0q7L6/hnQFNxZPhgetvsxjCGBjchmDxZJ/tRh73+wfADSWu
iwoPk9GORWMP9g20eNMVN7/ABSiteIz0UQSVj0t/EP/W4nc43iyNl9i2YKtFwLAB
egNMmXC4UirueeULdE22dnYmGFFY8sfA53bPdT/MD16jFkSKkB7iq9EkDB/DQRFO
hsNbCA9QB+3EWUFkV3MLlLF/obTjq+pouOQPKh/w5onzOliXoEAkIL+XsDlmjfYz
fIY6D7aayoRnLPVErRdnujI+a9ad+9PPT0o8RBMYkRuWtX1c7ld4X0U2fQUuU4ul
ALFVQl1eO4aulRhGsmJELR+/H7lzgphMCHqCHYaxU8VUbOcIveDZdtzdwxcTXxjT
qVv8wY4UYW5Ke7jgWG8M8odbZ3YJtFz5DQU9fmYON4iw/DXhc5hLLsNJrs7zMB07
FIcy5ARiPqcFHk7fSBHNyntaG82MBMFJOjPeBG+LsrBKvXAmVGy19HfCYEnB2yXX
+Ob0IhD5fJXYC4zgdnOhsvWG/Twjf65UXqiYyBW8F1haJi2n7BwpSvOE+FU3rslB
11WcGzdPY4Epz5yaUZlEH+QW9KU9uDUP+RaHEolssOXZ4FRCheWcAmcR82mS79Zg
GLgM+RxRWz/n9aeHix5MYuDjRTlvbVmRxPOr98y67xMPlqoQCsGlvzRjjMpzlRHM
f2Ts3n4sQxgMcvDlkWr5gpKEhp63YSdDI9RL/vTDgvio4MifI+bas+AjLr7M8uWb
bXPMOMYnsLZK9hyxD2GRZgLNqnVtR/Rdm+/2feNwPwoLlwTKDl5jAULSDoGNi1mq
J1xdHRrXY+E4DMygz44YtpzyQXStQ51xQiuUHvgtgPb4J8bkpF6ChkSqDmxG6AB+
p9IvgKWAT7PFR/Vb/qAUpf886IAauPFDP1eReIgCjOmYjJNYzNidyvAHhEQWv+T0
AtVv1aiWt/bRdSe3rlK5dJwTlno29sDff1CJnCWhA39UKhbboecdGb5RFRm7ePsj
jflE5t57yd3AYZUzwlZX+3C0sZzrWNnRXu0nnChLkTHTBQV72mYFWyQkA8lFcESo
fa218C4U5x5NYLhKsz5Vtd7I00i1bvH8Wy1G0P+YiVD/jWcF9w7y2ferJ+gjfT8G
Jjtz79aGx/985P3cATh8jjCCagn9PXrKKXZg3Pb/YFE2tkE1LC50jAk2e404f7/H
Kk5ObRL/w5BC396CBH7SGNCOHLUhTF1PvfE+3xndueGTmufMWq3ecHQYzE90EAsC
474cwERoxvG27lphe6YGT0jXTeRwfQfzqzy5MF5bAQYYj8EhbRfFhov9UMtWRVIu
6F6L9zlC2GhY/hL2876JL8I0DBziTdW6c+UkM+kWQGgHEGCtKDEYKMZSQij5T9DE
v3TShBVN3AGm+HafxM1XeOkXSAQmdkKfopx2cDAlBWmzxotGDxM8ssL11UclS7sT
heJgm9AJhWZkw23PmB3rk/P4qSczUzzzUe5SdEDK1zFThgGGKR3v5QdsT7SbfJUx
ipt77tN91pK/Ln75AwY7yXkVbP4eVZGZkuH3wTRPDrWz3dhGJFCJYWX2WM4K7lbH
2mscSGFnpadKykb9RZ4FYJ68bldCTFQpfnmEXrOYfdLn0sB1+frERmMgPoEqyP4Q
Ka8wHQoaC2XfG0eQ7n67wCQYmU15u4CgrZlUgxRIstdsHUY/w03MT4smrPQ+kP6a
kzjn3hHLF9rMm9Ru1PPtYrVNpzs8OXDBV3tkvBkOi91NUGqy2KywF3AZ8XsZzcSA
kRf5pnEOD6pE0GxoU2FaQ5DIvPDc1EAP7THeyRuW8c8no9UrcRdkZ/HXwcgGZ1QM
weDjmPlRa6km25+ZfACT9nlnF8ExDg3bicReYEcnuGAShZwa0KBFoDDoXyrh2420
2sccv+u1hWp3/wv6tn3oeCsWuhwWN9BbKN10ZB1xs2cYa7jFm2IHsXIGQg5+gS5b
RNfSdDHgQi4AIQqQb8H1LTwO59PiO0jeqtX3svrm5B9jcP11eNg4o2PH3stnKTca
K3kjXbBGJF6FKU4KzJMe3+JIit4ZQ4XL+q43iGpwxNXse3Z6MESUIABQa3t41mMI
w2fNFLnt2izUzxSRqAuMFYGsnFTGlVi4fbj3EUo/QgJpv/icntCD4OlNj8SmgDrF
ROKY1GEX6welnuNZ16zFoQBzvCikuqJSoM49nKpsWIVab6pPgkDzafHf1831+XYN
k7Vggf7RR81VTu1AX0B0w1og/RNeG1Y4ub7B1zdjdTndsd/fua8U6NChy09iaXl3
UmKEINlkBNZlOKV3s9RHBuGj2WuFhPikowCuYxDCDy142Ck/3XzCJve5jE5O9JKc
FQwRf5uuM0glakSc+xDFaV6nHp1iLIUM45ji1dQYCxiTl0+m45jReSjTHQOtYeWG
tqu3oiCseJo9YoRnVZGcBoEQ3iaRTCSBXSGkzw/8eZQyhM12A8nT32p143yRN/s5
ogCKkjmQbQYhQFf1H8k6xn1ni7ExioOEbA63PE/X8O63ZzYeFFwHrZ3GyUU8vFtj
8uYN2elhBoIQPlyf4YWJqsWpbZ4f+Sj0shnT21hNbUSrhbgILW53lMJKSdeSBLFz
MvvHNGva2wuTS4xwiOn6WP7PqBTyYYfe0L7jt8bi5wa7Uxc5kitLZFyXoSeyv7Mq
xllsKz9MWUe/JduflQlR6VndZ1P10c5HeatIJ5ISO0iGoiq+ESlxSQVb3mp145KU
AOd8Kn41vnnaOcggHNErLIzr0TO6gPedwnzRPdBWDYASWri2vujShiCJHkbj5zzQ
a7idfMI8cYOL7f4u2anV90hyACxcyAp07VAcqT6807DoojcJx5YS2jdNNEqmOPdL
256NDjaCop3bLwIvz/Zau3wGmbY77zXxypld6/7SVpINkhCyVUkZASb0u8Tts4+6
gkHD71rZrmTvxCoEn1VScr6BhISwFKX/7UJt6zao/O6tuJm+6zrdGkjh4zHj1EXc
lo5PAExp5Wf9Sfvb6JHRY7aUOHFMncaXkf2iNEic/rmRDAh2gtfoayGUxG8A8+Il
fJdNZ3O3+C0fDifM09FMBOpm79reT1P2/2gqgohALFhdlm+B6yFxjVLF1jTXzsTD
ZcZj2pgM8d1u4aBlRdXMvKy6LP4CgA0eP+9dm/wLT6jz3jTaYCgHPEeEJoPc02UX
EvGvhH53Rh1Le/xyJSKy5UE7ol6imu1hWQTUZwFOVBqU++yhA26RCVYwhT+QE1yq
54jYKZpmw3HREKJv09XKQ5T0px++mvECw4PzTrDlFktBLOtX5zYoYj5OvQoqkpDQ
KagsKJET9BhJttBie/ExCeG9x8/m/QHBGYpl5SqxPr2FNZGLdB/zRYS8QYckw5QH
zLYODdtwjUECsyJq1X2TmmVO9zl/vLL3Of03ISVG4CQZqFWAq80TXdP/GkBVX0Oe
/FcjgFn2SFOTvivn9ow7cjX8RpbxzeIgunZf5b8qTUp91A9GEP+0qoOi67hqedG4
xA1k37z1af2ISCXuEDs2wP3+bd3494jEl34+aMa/dX2urn6uk2i2twxs/DtV/n3S
HOhkqJg1dZfzR9Y/lWHz/j6ROybV+OoxSWI8NZEe3U0un6U9Xq2bpn1hxpIFgx0q
nq/hUMGemGWtE8V9Jyf0nGrAK39D+7trtGwQbGopqD/FNLiiWryczbg+bP94oW/d
pbhljLgPOJPtsdXV/kFJAg20QoyKm1apO6tHhua+YnNSF7a1jSzf7orTCCCvoQo+
bKwgsmrUM7xYHtWjxtBuHN5SqzNn9p/xX51roRa2TkHYtNC1TIhrFVSUNc2rdfd/
xtbxyl6w6pcOMlkNSfbIH/idXnEK22nuFk296b97VjKCdNRsGa0W9gTYbWqbSgBo
pzjOD/FhKph9MmzZWMmygjI9nTKAWrQzE1Ia/HOwSiJpYoU452T/dmGpe8v1OuWQ
9FtT+5uiyXYuJ7wn4Q1VnQqoU/f1698wDnjASdwqx+TekFjugVA1uowpuJCw5A4a
I85CqJB3xhRbUSgb2Hq+ejo5QyQjOE6tNJLyQC/y7+uczLI47aWmK2VGxWiP99py
dnYd/V1FrwguOvK7g1KSoeetPwvqezm6LHoqFemXtiZlXvJKuySK70lAlTtTnf5o
BHRCAjEIw/rVKJ2iAXLWGZLSaNNC3uYdtexjJZJBO8koSoW6GIfWk9Tdx6qSeuA4
n/sbtuxmIzLvVWnoSkbYhi6sjmGdnXnSyfZxwVqb5uxxwtSADBkmwpYBhI/WkQPe
iLLnIEf/u4zYiPjYc7J/fWdWaeqagTAiVlphEDBDywHUKhNhhxtlBcMlqQrlywr1
fMThtAJSvfnwa71r18UN6JRfiGHTzOiOBQ/uuxvd/pzqp4A9yB61F0Jl8SZUzElm
lwxPxiYA6QwqlV7lIsR5R7g/OTcQNhPj0Wd+ptVYzJ0r7YkH//enfjNFe+0jY/wV
pE8ikOJ8/oi9T7Yfl9c5creQR/m6oLgA5yuvqKPwTgXhxjkP8+8wjqx9wyM6PERg
jrJa/Hdg21FGxtlgqJ0fqU8y3nBgt9U/QyT2JGCRcg8oHAqR0UILKrZsct4NTT7e
HTKUw3E3FjSTyVfB4fAh8on5CysWQoy9xLs5sUsHZkaK3YNl6t36IUpRfjPScsLI
Up8Cbs8J8IZsHtmHebYRFKsR47WZDtOB7c4dOSo/Tcs0ucAk69xpVmhkmtY3TDrj
HX/YyQ74RE7oUllNemSBLa4BwIvaW66hz9lm2sRrtSNvWs3K5ctw2xyQ0wbv7+lb
Q6ymP3IuCB5EKAZAglhhaHc7/uud0EXd3ybe8YSzCZwe2b09qofc4w6p/cpg0EfO
txuESFAXPL5CfhpB/luLHT/DtNEnAN6u5nbGGiIyJtPemv7JMBWqWOe+gxrQ4L1M
R/Expzy5JXtD8OHC3yrXIsk/sIU7RPsE2gMxvnC7GzPXAgLr0+xgTmQ5fWDE41V1
3bwA8Pb0zhI8ZH4NiiOpqzksk8dH45Kf8I/xh2BaGSKvvNczEN9bgzHIxO1CyLAa
MnpXdp4H0H90OMYAS2i5MPbpStdQfp+x59lu8manWDfml6netZXc3oukbN7YTouG
2igZVoPUw8Tf1yJjkEOXrZwqyxkIN40P6UgetmipMq1N8/7MlSrN4qrDsQgBG2sn
EG29DR6o8puk01br0wCJj7oBZ5a99e9K3js5dlGHRUExwEeiA1UuCBCwuiHqxhwW
Z3ebl1hKdgP8JXoP8fdtY+8rpsdzguaGWiEaKMfbrYeqx4k5Wwh8zyGXeDo/VPuP
KBpMU95EKJ52BxdlCmah9FF3thWSvn2yQjsBSAvGjTZ++fRusBEGksNPmcTzMvWE
pmIvHZYUawt6CGOe7qexxGiPC//+rYUtqzs8Ge3zvhniujtAE+JsOrX+HY1cVAE8
/4dvmST6Hz8t4OFbwexbRxEdKx/BhzwfNOEwfavJIdNkK4Pwfp6FSgteRh51/4Z2
1rgsCcQMs+3ZwM+vXxMck2zswH/TbcGWAgzJ4rA+kfId5NzOrc8y30yTEXV281kI
WTeNT91UHPfSQ8HB3RdGiS/2Ju1jmQFKmD8xyNoDTIoc+/dUdtk//z7kGEiHYYoQ
4pY1+ClKvVAypeHPFnMnUSgmh2zq20pqT6fU+pq5gh0MZS76g0P3Ik05mF4RMFG7
uqcLsZmsfdjcYi3E9IGmynO63QMc5uDtCV+hNcpuMbsTC4a9hSwgBh8nqF8JZT/b
ybnYEsEMiM6RC0gJM02p+b+GlvMqVGkc/9wPMunrbmS85k+ZB+FXmziWLoJBZ8cP
H2HOHEejCfHT6d5FitL2No4QKlw+hOV/ZyYOOw6GnaTqR/C26b4vRIkOqs3Whjgq
qYh1Jm3OvugYyZbF6FIJ4hz9FkXXGPDuS5A3hne3JIlNVnqnpLtJ+TThR8v5h/L2
LuL3/3f9XhFzp6aS636UIQMHBAze2G5KxMxW/C/Kg9lbugKvUD7weeWSFdmZ1vjS
AYcfNYfRggb7MyETVL5a3zytzyUjzwQ4IeelN59jG8gcDZbnQ4dswLX3g+9Ot5au
u12L96ZtXMBIWhS22leDbXr6t/5VrS4eaOYeh2KktHZhHf3PEnu45v6HWZp0AsAg
7Y5ck02AvC6LB4mN5IFBKG77jpH1Insp3fEdtu1DWftjpnQSRM6h4x102SieftKO
a8Z5g/WYFZcO7Seiy7cP49YktQ5iWAksRurSwyWXOlkA3Nqsc+rIqtqKBZabE0jO
B5WxFydBGuDXrNDNy7o5OCfKNEk6wDE5YJxJrYkWRg6yFiUBK9qQS42c/60UlOQW
km2taWsVhhZfi28RRrKMiO5Ds5/Wg0kQ86O1kVAVPGWaWq+KKTepRNKXz3cc5CJF
uf8Mb44K0iTm5rde0oUrKm6pfuDbsl4BNDv+Ou/imWVBjNKMuue1QjwMlJw2Gtpy
tqUP+Dw3En5sgMmkqK9hkN6CC9sCocIESrENwAUTgdbaK2YAJo4XLE22WL5wL8nY
dFT/XtRCpec6IDFMQgq2dqRX8Z3wZFC+vB0F8TeM18pwoY7nZOvE+fEFFi92omyE
exvdZsVG6dnbINPqACSfZhoM+2OE5rAEGMKipC6yG9vHTLPhCaCYSqw3V36SvsI5
TTA9mstf7nIZo7bSI/+VzSQsZ7IojiWYSZHmw4nAVAERwto6q2Cop0Ss3uwI6iBS
Mq+A8EfGxIJPV1HbwOOhNIZoAKTculLs+ccdI/VoiTEb1FlH+O6AD1TvJ/5I9/kB
8MJHjZDIl4snxvHHD9roake0CfcywDOSb7wKk4y0f4W6r4AI/owazQlSN5s39btP
IpYpPuODEM8p68gN2o218GdTwA/2vMs/ZpzMhtFczx8eQ57dTGjU9i9KuwsJht7n
9v8Aa9l3dpLXonjCErYZhohHoUa6sCbGPVQ8DHAH7OEPN/JhhO0KZga3wtpVOLy7
uw5awL6dke6p4EB1MLKhTyryCxKjqUSbtCvWWJPPakcOhWL+SIokjvF6Yu/Ae0mj
MRsXeO7UES1bqS/EEKYcGZy0MPvkmaZK9pVd2Gv23UVNDwah706G44GRSIVostUi
DMxhcgYo9D1iBXEAldjIlDgo61Gmeyc3+kavg54kZNsAgPaGpIy6vspt8GD+W8RS
XxW40MVP8Og34bwGKuyBCNwsB802Ety0cJZalHJwTlbhHhMPb5xEBjtM0KABv/F3
QXR5eG07vuLxYany9lmzHdoeN5wdmpOwQHtPVeAOrvp3XjlJwGMKmN/VI8rdaefk
zGEkuwU/0GLxPNliDtX3c7zXwAOrdeYrlOGYCF4uPBgPmk6+W5gAKVC31xQeMX3d
L2fnU2c+cWo+w++Ay4CQioVRnY7MwxqHO+dMNPQMLLnzanwZ2FqTOW4bA/uvY0yR
drowy0de7ifJxlSq7631nuoRkTzu5aU2eYVKViZcwIDEf2J/UBI09SlUj3lOEMsM
YYC1zG/ANJppSBVlUxrt+r04EG5IAeqAZ1BpWyFmb38tUdwcnYjzbINiuMOuOytx
1mRLgxULKK3VSDjbrgPwcI2MvBp+JCfo6d0C3UYTkHKHdOzn3P/rLDlofU2XWuDy
i2faeBuGTIIZEh3jk/u4ORw6U8UslOLt74A6Dee9G++MwLu7RE+phcw8ma49mMFT
K6w7becIqav+nklKUpIe8MlP6c0vZNNlMCerF1wAal7gdRONzYTPyl7GPiptGk6v
PAbYz57yVMsgFa2XlZZkYzuZzjVayNJGzf8BmaKoV7z/1H8V62XtZnMVds3S0rav
31pYIE2ox9i1xY3eY8PUoEdb/kSwGk7Jto2QnxfhkVmVI936HxT9ML0LyNeoaQrR
3i2MF1VQpVJGXTFaVTjGCvJunCI7anQDVaz5N+FGEz870KlFMWQ9X/l2JPh8tIRB
/6xWagRUxUG7AdLX58e/qh8fDhEvnvqZsu1AoZ3ljSh/eqJfALLJnITDlccvTxKA
hf9UPa7z9Nv7V4tV7p3JEvnEcoEyL16JAyHO16DhRkyaoeiLrkAur4Qie+a8DeXV
o6gRW2xbydK5kKgXQaWEqi97aZo/1hDhISf/P4/rYVWzmMt+MIXh+z1qVBa+QsMI
OgTbOmjr5pSgt+KZcfUuUVFaVxgPoem+U+8aTT18ATka3zWpWE/WfwkD0xw+smfF
RHGN7TmHZh/nE2k6lWrbiFL4wsmJ+f6bPVvz1uBhV74IE47X0FPxbvL8NSMoyTzR
NTfj5yARK5nKJnjuO70pXTNUvCPLidH818nz4eyMH3JoKofVtzMO2n3+tOZtz8/9
RSn+s2asB8ApShyEyAVKEsBp9dJd/T08rTlEC4749qttHb+ywY/LcLI19VwKVDB+
BNcfJclFGbxi8OLPYLj2kxJiQNj/pFuBZs/uFqHwquw8S8+/SebSO+IumlQNucM4
Fji0YoB6OozVYhimVl/4N6Z7l9Hx8t6pDHhF5cU8UFBfakKkJUFlauYRrLwLU71B
sgu2SRAEkl1BxN0kxKAM/tYj+/g8UkrtvhIJ5EB3fpW5hU7B93s1dtoM8Wk+cFBF
X8uOIwb4SSvlqEILAWiKZQqXWd1N6m3D917GHYFtVcWfcN8JsmQ3bI7dbtXGEwl9
6P2CR9v9Jywyr6WjYFjwEd1t4Ftdl0YrcUalfVHgfIa4PCOoksG8FNBxZBrPnskR
XzfJTdSfvOjqrSIOswmMIbMFwUuVVsd7Tqq7CI+noSJhh5/ZensqWqsij2aP+AQo
f5RUgUlIIWtDfFfspVwDCoW5h9tug0gtjAYi7t3eQykiIuTcs8U+Fl49/6Y9lqTd
sHUk/gOTh631zAkcTWSzmk3xiBBqyiMGNV6dE5rdjqQ975PMz5aL8Ac3VWzwSi81
/2ITxUBHMPk9xJpTdGiGVjtNy6Wc64w8/ZvnCrqyuI/8Z6mC/wpmWcPZkMpEnqMm
jlhOdmG2Y6I4E0NRkKoG0xHK8KqE2njIuK9ipI/PA/lqVfq/1L3DOlNbS+3btcRB
qLKKrALBv99q2fWZu+6X7R+PFBrHSnpyqcUsVLnhP7cyAzgK6Id746RZ0seF91D/
L2t5Q5xnWs8wAMlRlDJJPBPP493yaZlicGbXl7b6GAXvp5WWf9BEIKWRwO2xldby
o7bmCshn5SDWSoTxnjlWZsse1Z6oxY8lyk+PHqeyXGxMRz3/++rsroaU6EeZsqoF
BF2gbOREHeDixiV+02dCFfHLMzVAHQyCKByrvysyzTqLeA7XpYtcvp58py3unavC
74Shu6Ey02yQzB3PBrbRURCY5/SCZcMiJmmgkb0apEnk2MlQ1/Jm0dP4GI3TDFDf
L3kmatva68mqw9NLWp1WW8Vtc3wNoX8av0Y6PXuaTyZjmoIdtQiBdbElTVSlSrfU
lqjMigylV5qDPzgdO6g/sDHoBT1vo0Bod5w/tbIOl3PYCasrCo4LbDMw/Uf8SDS8
ln5VlWdkm2LFm8kgUx9PnH4IyhgXWIaFYOQXo+6zI350vO7ox54Wlh24nhgOYU4c
nEIf35zskAvM77x36gn73YYliD2vFlwvF4P98ywLXDhFXGYEqhh00+Uh8Qsm2z8M
oapOtM99AxUIikRdC1xmKyRzYYS5b53geU/CAXaWYUV1lRjCcgunfMMpnt0mwcsL
/A/EbSgMKeUFWQKjz7+UsNtoeg2thy6xyFTqaw1ge1xiKyOZkQANj3PMYJoq0HNs
IfTJIYK8qGzEZfxcLfwrJwTB1oR1o9S5LaRWiKSiT4KH9j55RvuMKamMECjJc9DI
ZyuDMTlYQ0tNUw9bNXWhA3Ted3kijnKBhkGyHZ3U6EFK8oZqyQkAozR/DPOqmo5L
zKaZW3Y3jzEJM1gTKtyAB0R28ZCXRpghI4ZSl/zOe7ZZvA4ArwjRnkID/eDX4ZED
14SUDpn841prHl27kaygZAzkP5PLVloolnjL/YYb733w67G06PPUutLq4xAMw33d
7E59klKPxdmBfXPhOa46FeaHusW1f/uhj67AWgSEqC16YDBbzCWMswIC5Q/EA7V0
hLMwo4GG4W0GWKqtGFygLNKOe7OLCQl98DY0b+zVdvk19UPwZZueTHTCNKRQD/Qx
zM1Hn4Ihx/STOHbQD7a6Eujy61YxtZVx3TylFWwznAjUqYWciI9voeJTVrRs6+v7
EMl6h1ZG5DfA87cu5b+lsSc8ylvSaG0852C6z2ZvQzwASPOOUFnOAJTbDjVEg612
95IIgDcMDzghPU2AxozEw0FvcFAQOa+nGuVYKFF7JMfwhhBIj0pWEwlEZpUUcTLy
M3StdTT2JlBiI3zpprwWOBBllz4c6ZpyGThgkzRpE3kNxPNt6pT8x53ONBXAo5xO
3QZixKZCQKaNPZ7v2iu6RIbrcUs+Tg0AxoV0ifRYcoTYWFeVcBpKtz1VuxHyP+mK
mqBszmwgtiqidItGbYWXRguWrmkTe6uA+RlfL09tA+FoRHvfrqHTrdW9Ti4DLr9U
su2dmImrzzJHdZV3zn2j0en3qP5XABUmKqIsr2lmRGEsLUlxQVfQ0Qf0XowS+asT
nChPGHkpduVBlaKJE2iro0bcEyG/ifl6U+bKLXmqW9q/7rj7syVDHT0uflRjWaur
GG2CgCvlvOyCULow37HlFgOWV09kSmQGkfiVUKBpCyS1PkL3lDTaZEWxy1nQA63X
ajwez9dSYLIlcvznXsgx8Rv+LB+j3maxBf68FpKtNMDiCSc+mKk8lHDhF8mtub8i
0ihV12qrCB8cN/t2xY3KvXyuLAhcHUCPSyxNGCbCgE1BnXAkvEtrw87hm3qDEatD
F0rBTvczKqzWxYOZTz+pRIRP4gI9iLlQrnp3EsYG0LPeBRoda/V4M9rvNtzKwcBr
lLrFDVny7j738z9VbzZTo+WCBPEwHtBXZjaUPLJ/dscoOgkMYaNF0BGsAMq9ey/z
p1mPRJWI4l3eoX/aao7bOPNHB5rXY4lBUCu3kLsdzH6LZYgkWdu+xdZ+0d5fR5lR
yCWEuFNPDl8StR1L14nUWYdbtOD5m9D4YIjTDIOH33P0u5SyO9zXBSeKqJoFw1Mw
xmH1mfGDiL3txK0pGNePZ9B5PGE7RHvExSkrBULFwUtpzSaYxo86eyZozOTo5Rk5
pbsZBKxDSc5lOT8u8mq4qip9qcciermsEVtPVQJeRfdPwDv6GkIiHEYQRiS5v/3B
JU/Jnz6ArqWZaEBQ3ubHw4JD0jZLRjmIbim91SSwYGUYmL1DNRQtx6teBLPtxuCY
K+EBakl3aHIiGAYCbj8Ac8fbphiBMzk/b1RwXdqIa4QfrpS130oIjcDGvqW+LaPN
TCT1JkBaS7gVpihd33EWXh+nJigOIAGvq3emI1YcC3nIV5KQUeYug+dT5TAd26f5
13TsdBv1yyVS0uYOfSXNuzxv0VQ7ll4JmeZSCgrtkC7NTiPuSZJLtKeyYjB2RvOB
bLU6wKsNnI8p2xhgqgdMd7lWtWJdFq2yGfLUbxJw00B2T+lyVU76gao4QghnFTle
mFZ86dAhy75SG30/2tgTcdbFlJNXWL0A2FCaljiKsw+I1MYkfoZB7PgSrZPZpnj4
v93RiLq4A5jkdjiolt+md+LRyMGGb7Vg8tXzrudHEvJRZJXszXBxl8Rf55U+Z2Je
oQVfMX63Ci1wRkxKZpVgLKym9HpTPB9OsqSbe+hE5NsMK6DeUAOdzqxdfCKw2VP/
zpsqhi5GRpkjtbt3/UoiM/DPLWtHOyWl6ROXsAjOC4+trYy80cpJN7KHF8IGEXnz
LUTnbRFVg82zb+iMDfNn0oYmR2wIyTefFrojkF4rcd+xLAfeNCGx4+H38feAkCiJ
1mPW184xtBqpi4JgYr3phpLycZkpX6B5FBWbBS4nCuD+whCRdmx+l399AzKW44I0
ZHTwkzS8Xxpz6s4uhIJAE3FendVZ+I/qhNbE9Qcoj60SMvm8OfOy6DPq37QhbqlW
D1K6FI5HULqiKuNs/ANht9wRPd8zEqKSgAHIEvX3nvMtu+v1eXaHpvl/tDH8UkwS
3LjtYE/L1nNFDxaM7RM7HM9bLPIeCFP9DEA37GaUEl9ajDM8M4PMiKXISK3g6SJF
BUGbYChz1xxHbpgzhwXOxeaCJEouW9LLJDFTVboBSL1a+cGBWH8zCcnm7jBPTB73
01kTIu2GabhAHaWJX3mKvNHqsz4i004ptPmsXKZb/YOpG4gQ00JeiRIX9rSwybOI
pDipK+XxeDrZYgbenQDAsPRMbVf0pu1MlF2UvXEzkWycjTEj8P9OAgyUtZ8cIBHV
npZ//ujfZwof1RJLhHhX7r3CA9nk9NbDIirrNxCmYiqBmMvS7FZB8kWRCsoV+Wax
7G7+Pz7/Mcowfq4kI1ztrOuZpAL3BHBITViR1gLyUqbvvck9iMivREwW/gnr2Q+N
V7XY0CnX7zQw2wPjnaIW8uNNaMRpb+mhUFg6KAiDOOlgZmZH9qmhQXZnzvx1IMwA
OtziRrcfp8P2QjKj2tShANrwL6/gfGCBRgdjJZtHw7i+QDZ8gtsUmGDK/meMg2iH
X747bBzALcZtbyKwl3Pg79NWBoXq5dYy7XWTlzLgE25KlqXrYE+Ck96YxrydmerT
wgCJYxFGolpliZjAFP81kp3cpZHx4Wmps/9/SIk0lR7Xwy3KuSZsp+gnriBdxSQG
uVSWLI5cIsaVD974x9zoXbDArOoWQ1bGQo1q6qphN88UOMHw6RUqrjmLqzmOxO+r
LbvsvmE9zAfDulxI0uAWDjTNFNJ/RK1uw8/Pa7aT+tXMpjqUe9fNcupL9EEng+d8
Lj/v2UWOZ/ohCpw4TpP+5HJfMR4FCnzWiuB4Yy8LOcnNb+CtBY7XwktgMAehXv47
y/TrhG8llmEsDb2L8XKMhCKY8Vyao4bidMKxnxMaFZrqazdmjLK8Q/JIuP265qgT
8Q5soxN6k2oWzTVPJ8T5hibwrlPEXhlcChoQBV0DPOr6iOj87nM/a2RS3LigkOc2
Y1gU4+ZAvD3Hn3mz5SvhdBYyh6bwAcg8tEtzYJ8lNlIvwZubgEgoHSXyhGxFF6/0
rT516HwV8q8SxULcFvsSNkUBXdhQOKhQnXkau5Jhoc4KcXoDBLlbCrmTxdcq8EhQ
dM/XuxJ1xgXn8gwCdX7IT3ZpTrgP1tsi5nAX0FMtJlbj8Z4LNqeMHkBnZ0nqrQPy
IkayjxJ6Pok0UdbUXwjZw6OfU4kVWzhsTb1XohEmEFkF1RLi4B27ew/AtTcU95c1
thJyw3L6oQ/9KsTnTfeAC8qj0OAweFg1wO8qC4KzGfekdXxWUYS4jKXKQo97Nml9
CUhIdoWb4AVpv9edHtbSKzTZgfHveuYVj3sjijIEPcC90JrNcF3YZejFFMUDr+eE
yhzCQ5WzhLNa+fUWI6FbrcXTjZ5dbqQqs52+irLJNgBtE4u3knVcGcR2Y2cI2Rso
N+0+AqOw83tZ2VzBpbM7C1fX0ESTTrLPfhTB1hmeTDXukCo+oo2qavRLyRMLgNPM
UYVNzO5n8PpM67+VgU2RJipHc8yCT1bdyh7pBPKJDBLL11QLT0O5oNDtpdY3d+62
dukDR6DjU6qRpF/XR7vyYvigYd31Z2ZIyDY7GgBrXgxcB1EVze48iPYvYdm7cA9V
eH1zDEQNMmmQ3mHwSzz0WMFCfB9VPlo3Fotno5DZH8mi+ygC5AfCNCw1bivIRnaO
SprLxnNFwJFCgzdFAmNEMBb49veQOS1vs4FWyclr/kMyUVHnXWLBQo2pxmNZ15s1
Mh8R27tMhvEtsQPGbWpjnvZnKuQspAnhXnB/0w+zVki9VPHQTx4Bq1e3RWt4Treu
H4Wp7+P6VTVi6civrYM0typXVkAMI+EeW9uo6MrjHp1y6rm94Pa4gTqVrMSrpm4b
P+jZD+dFf4REJsDfmpZr0mN6Ynn+gEhrjn8yP9j0Q0lwP94nNK8Q8VnbEFUjk1QQ
wNxrNZP01YxQE9l9E9rtCdUJ7Ye8Lvd/A1qxFLBU4xsPvYoYhcffd9tAiuVIxau2
KO5VaLcdiN4o5fCPDCKRIpUXXzpmZVPU6AWTvzNUQ1dMZQ5/0i1D5iCR99qNLyGk
90EQhachcb0lDd6+UrTQMA29p5/VGLseaTIRtg3jCn7yXcPlUU/g1WN4bRNWwDnh
xGiinUy8w91qE6J7UmADLhTs9sMRwRLaWqtoWwxI2eB0FIEs/gISXG5oBTtqV+u5
iGa8lazzVYdnyIDSsaDU95FabnBpqfl206zWU2otODLtn/Kk9VDUk0LGP6ZjcLDz
Hw2xgn85wsHd4YJyZtZds1vcbe2qMSb5ezT8NSObc6Ivvx+q7kP6PLUuSIjWiNC1
bJKvgVIGdYw7w9v5LwCOZOl/CVmg8slMFLsq8GuR9tzeUkWR0OChoJtZ+nKFeEaM
qrE7l9kdjclJ8qVpzQFe4gMeRP29UbTpjiUkAln8W+CCkvHhqG6r9k7wfaz3pxsv
jj2TjJjtiKEThtCO1LkkmsdJWCu01wXD6BarVWIf6PGR+XrSc914142lLuy8cwZN
6VZ5eBPeP1tah1CKou24U8nGIa1KzZgkClnvjUNuqNEiGT77GspVC9EWxGg/gcB5
j8vmSk9I3rEbiRdMq8j/qxQR0LiJak8h8eSJnGQt2YuCyBI5p03w/FTbXWPE5Inl
3f1JOoAvR1t3Ftbn2KA1gBN/bEomC3o8bqvVHWWVdnM6bt/l4LPun3tlUMJQjUEs
zkktSwNbI5BL2W/mPFPd02c6dAhnA9jJ48J7vkYDyneScvieT3hmjT5AccjmRGh5
XPcN0aIRxIyrrsn2nCuEddlVJ6ITCz8lYFRG17xbVQCSK/E0bLma5rQr+Ph0XrTy
tr6oOZ+9G38Q+Y4RadtKZ8+ZYvSKORBSgkOexpzxawjt3hsYid/+lzkmTfRylHBC
v+AZ2OBLzVU3XOYNoG2fLjS/ljz3imOBHrWppHzq0Ng2F0fRZosVq23XQF8g9KUr
gzxqMtXhkmbnvwqDOsIrU5Dk4n7fZgnLn8b5d5B0H2KyVDeT/u5eDlD9RLRfHlhS
EqLd2Wu006iEGilFS506RFeGxvc9KJ/DU5PPmZ+aAQHA+1VF87mDsrIICHRF/YRl
MuclRQP+pdjxQJQC+e0czAKiRBnYAskIlC7Ct9BCq8/7uIfaU3s5XDxceHCbUF+a
oCpzYIYM6QWz87yINRS5MviUi8R+pZVC4mraIOSc/pa8lxevpR2f1Nu68F+p5Svr
weMWt0UT/DaU45LtJrn95H7VZ5GVJtOruyqxdJWJWJ09fSpL4+RiLGSSzGdhn8PB
oQ1/kYQafpnYR9+QffOtGOT8Qs9C0aBlEBdStuu8k6nRUokpfiQE0FXGRV/tReeG
i6wVDe7YI1ks44PuIqvGESPkRtW9X1IylW5Qbpz68naU55aOa8JSALZDOoGI3bp9
IQghUgwmAxPZRWxUvBlE3ULD5zb/6CJbWalhR/n7MrHKoKXQwStuZBn/chNevgoo
9P68k+/V94EwDid47iAGlZTsJTuyiaBZ6HhKFIjYVmQkPqlYncdBvN0jfrqedAo+
ZTAe2OH2X/1De1vZtgDkOT4EpnWgLLBFuUFX4cNbrK2x2zb88JE0MCcfU5BKSZOI
VkjO2BS0girxMUY9tuVb9xAd4UEe7jf2kFoSOy9oj2q8HCnDwT7WLxThOg+Af620
fnbgugu2lBoLdOgovcuirbHURi4wnAOc/OkAqXZ1NruwLxsgBrv/eiKuyuwuBK2U
3kXCRFrftSgWY0lDOy9pk7T4hb3wzOJiiRNGxtiXQ9AsFDBv9+mgyZRWmvz7xGdJ
Ib5C4T4qPhbzz1dtOXwPSw2T3ZsCzvsr1KIASbLtbjlKJjFS5InP75SAJsTWGOVO
/A9c5xDzzmga4w5YNIuVqyAucwIACJYgjkmaj9//qslpWYqjCpvVsre+PxbtfUGN
UPaTBAPrSpkMUOZyfHdnww7b92/LP0y/y5PMmShczOg5ZWzlZYayaAvVrvQXKtF/
SBFjzeFA2KOcuzSZTAlRmbIMuwLi4IrZk+6Fneiha697O6s4P2NO3kuQmbm0I83G
/7bVw3ctjc5URdAXZT+OdQl8JZDoQlmPxLMrNXWR9DAa9JCH7enCNteX4jpJBK3C
zSswHl+3w9VGIb/P3+k5mc8L6XwT5k0wk9MlVlJ/MOwhyX5JI8qiDU1dcVSWiSwx
4d1Q9IlQ+qdHez/QgwQhfIwMsPpAVn/cNyes3FljjLv2mOgcqePca3G4uDPi+CM7
du67U52YaFjB+BhGIaGie2MMxCUkumkVgaCwiCtnx0esH/tO3sO1RWrWglJF0AaM
Geqxi3bqfZY43iYeGIz0+w6kmN6HPulPnNT7lcMhwKjYXVFQQBzvW00lZkIDezkW
c8/3CM4nOxAy25FTdRCYifEL3j/Jwi2aBlcmrPRjsvgHEl2um0rpMuQ4mZz1LxjF
602fiwVFpRZ3+PLxTMaaYCosyS+pzTB5FjJNqxNxU1g93GqWwYg14C+5PmM5Y7kN
gcTZRfn8mHN4COxGJZs+tNnHrZSeADWLINqogAwjk7WjZyBiTC7DI647PdbmkZSv
sieRaFdgtgF9mTcT3vNtRPYiPOgKMfq9vdlHN0uGr//85EWMygcRgDIcGcBwszhr
RKX0qR7sIzDJZvwcoqxkrXlDe+aU0rPPNsavkKJrNTFR/bVREPc1KGBGa3mqJlpZ
l27WJ2YO4emJkq+KZxThKH5D1o6fOTS5/AQUXsSB4cJWgxF6zR0URCKKWIgLI0ap
yAON4whi3H/G6YGgXSh7YTU3rkV5sYqfFfIUXblhglzJN4tb8XfP0hhvvYKH2tSj
sWmDbvsquVxIcqwTtuEsPAaQiVD0LAkhDHiDHf0gyU+jxkAsagIrIQcuW8Ub7Aw0
zacwfAPh6klXJoI8RdNFJgHMxB0kWhYWEinQqe463hyhDR6Ex+DKf5o7qi5ij43r
xcvvIJSpCZfpQkjCYBn5fqIe50++as9RrClmLdJaQExC0qdg0huugCA+56kB6Wc2
Z1ZoYvqnzSf1R5k2ILY3wIcuSyQtwrdWImhY+VYTtANqtKcvMSPx+24niBaxUhLb
ttYB5AuES/HGvMUK4tVSIoF/sQOPBYqDsitTwOKCokb1Q2whQPIFQcGInDMbU7Kx
Vn6DL7mEyjBtSOrNgar6vQTEhJ+JrfgbhPyr85+0/RvjqUrJzjYSykMA2YKs2Og7
BDTAj8hlIYVd2ysR1RwYeKpCVcjzqV0I4NpPVUSxStcy7kRgdhLiaB/xy13tlrWO
gYtSn5ElEYB/W23Bx7txP4kfWU4hZ52pUYHxslT1ejgP+v5SH3PvZo+VQaLAgei2
nOccv+qwjJfLGT4ngdmQarEDke7YXM46KX8uTrBn9vzF8DXslmExYdCQNxWXJ6gX
5LeVMRuAzH0mvFOq65xR4y1g/Erj28sUw1B07jCUlevmG+zrov9qt4a2eUdmal4H
94vzNJRfOvVc+ZC/9aDLixoySt+dhxu8pDDoGdq8qbsRYfsw2YIKlN5ZyVjX5FKk
et2FxnxktVO75xm/Mt6y/zzB6hL1Kt2JxuHnOUjttZnjJKzFSd8bPVi9pEPrtMAk
MmBcVUXRZHb/E+gusgioQAIwwMowx5YBhq+VK7UGs/w0LhiA/gIlOxA3PUldQcHY
zIFLA1oLxn/7VvY+VrWy8KuUnMCITlmouh1U8IgeZa05pRN6Cdbnx7GfApEorcEx
nV2dlBNwkQV+2qbqb3NQCRWwf155SLMfbkPy7AHGGDWfOpHdHBijTh11KuBwl29O
nsW0QGWZdU6h+8mDndk/oDHyNbBXh+3f3mWmT9ZRCm01HcjgJzxm49GxIO5g7oPP
BiSYXvmcrDK+0I3Qdylqaj11uBaXmNAXHS/PRgXai6Tr3FtIKirwl7FlcREuHhpe
ezjalm/A/X8OITRSVf810YvkJXZYKvv/RX0mV+3waFpX3qtfgLQSxyAt/UxpPKrx
a/CUdZwvGvXfSyMKsCM1wtLGnheSYrl8hMHjbznGiHMbI/jvBQqG3khyr3zKz9LQ
gNeu19Defh9tp5X6pf6G3JdOl3ahf14v4s2V+HCRuiMPUvUK+/mtU3h5n1AgX3WN
JPshm1AbchA7Pg4a+9KsE9IMiuyds+wCEbg7zzEI8pdtMGDXN9b1iREAU23iK1IO
4ok+V72YQt+4KPcyf89scLdW9Z7gJrYgwzgr6bUT0vQGceVczilKQqpu37cvuIye
dVnAdnIyEMaf+Xzoyi/NcP5pTPB6HeYkcYOo+IVpaDBWIf7OVZo48WzID+Dxl10X
6xrA4+/3G3ghFTIW+qyCILyIfi+IQM6yyL61GX5/l9xF+yLVGbtw2YZaKhnwYRK3
K8b/DvXzF8lLXqb4RHdrSv0zMs3Hbv0RMaaeAlC1bY2QM4cE5FQCqL6DJMKRztX0
88BntfXMgcRZiNbX7P8OOohIPeoSr1A4sW3oN4XNaSdxeU8nH0WE/jD2R+tCj0Gm
4Ci1rkovApTXDt0U2xWdkHQCl5H76WoIk09iKozDwd4CI8ifRD8rZ7MGW6Um3TOk
8Rczc2+uAuJfeNHr1jnurAyOph/AE6j7i7oqfPebLDuhzLz+nMCWiCeWjvkjijOX
Yq4NcaD200jfUBtZEJIKeehmh56bk5FVJSn5KTfOZnJoR5WO6Xy1aupQL6AdGzjt
WAxOHFYpmog11sok78/Kr5VGTvVshZ0t2M6hObLbC8+qcfjZZIS9NXgPtob+D6o2
Lbwmmfaqz4RqtJa1QapBeFqnqt7+A5twiV7D4JCVhtkciICE4BoFo64otXXDbMFR
eUtmstmh26ZyTDatUKQmrR0b1hQFTIz/R0pTwIXqf0xuGZkkNat9E1y+KY6crJlv
z64+M+dTJpSB8wYGTP5hhGbWxPZxzT2hgSCtwunO8bLupVdg7akxLP4rlIlj499S
bm+j4m3nSM6cVnh8XelokeocimWQDLKsbmzYm5brKcBEGwy4pz45YNrYDU7vLdrX
0/zOKFQXyckrG12ycQ83J6VMnkHcrIw1is+6OvpgwTUS2J30s4Ty24KkdMRhSTqW
orkLGPvpBQtcTG2RCf/FRfm7KEqG3EYagEKzNmkbvXlAmPvg2lOdoOc6wfBR3ttD
ps/NJ4zFBUU2t/golJLMJFXEMj+CdwbvMEgX9XRqV7vB3cH3oLhmReHgOl3TvFQS
Amh+QauL5vdGI+iwKLCsgSdiz0gLh+fE5B7FoefVKGn5BQNi4IRq1PXNtag3YZjR
wgUrT+Xv2g2dCgQBRmEzGobyKBvh2gf5gjSvisTfmsnSBNnRep2EiSJcW8yXfppE
MT5p4zlzBWmsSvZeJwcndyAMFBziJb9yLiac4zloETv/NoSIrQcFbKpzTFhAOLXJ
FzgHd9NoiopRdkrKBldrmnZucn6Tlul5n8qgpoyCRXbOTQ9DyS/CnfVpD399+e78
OjSd1xdnQCpAPW2nbTG2Of0CDIZnCy8w1vOd26nGl1jaqQgE7XQ/MJhyvw5TW2zk
xsr4ymFZnZ+6vUhgUT6YwV9JJj/WgUC4GPxZxo7eY6RwPPY2vMMG7lwa6EgCFyZe
isMZoVRvhuhzq4t/OXwn/49XCKpnq/SQvJ4Emdrt1JkvAC6P2LbZbtKTud9Sd99A
RZb68z2HHSKTpSH0CLtCdRYHbmk9U75hGQG4q50wYidLukBBiaKr0oHFzGp7f/0I
VKSofnVBW7WTkEpITwZtF/S+U6VYqyhBDmMgYNsdt8xDIA0e+pnCBJQ5l9WbwlMB
wwGvVMsdpMx8mXuW0dG5dwsSo5E9s5sYrzKsrEyl5m9QnxTRFeJMzhOHZ8Y/wNsD
t/J7HoFgE9odeHxbY0lOn6NHfCRe6oCcWwKfGXGTB0QMFWgRXixVgmPI27LbtV5Q
b8LFuKM67NfILBkj9aN58UfjAGCLoHo8qVtogf/Bl3K1PK7QcNH3NKkglY/GW7bb
8X2SsKtfAJHoBSXy/EHh6h8ViuzFtbg3GaWg8xQNqQnJJMVpYKFlae90/8/iufmF
xG0SMh1XAMISj9moJNNZ08e9iqWR4n3OEUbIqh359yxtjhxrWByQHnU/hj+vHiGo
i7Fk1mOC0qXBR5RakOnJHdeo16R96ullT6bhx+Zhxivej8UQwNnWwZrR1UrilmhP
vJOBUF6KGVi9XfrpMcp6a2jyzP3wSQ82hJ//aersI1Fsc0pal2FiEX+TiyCXYZGQ
yDgDs1pK4lByS75/8F2Ra3SVU4/q8VcREah7ximEQ+vOd+2JHXDZ0PosAXnU3S9N
bw2N2aa+aOtqM3EysJGYbwV6wtoRSgidk8J3/wje8hvNzwHywea2EYqRR8ZazjHt
GqlUvRDkl6/wrgDHVj4afM4Zn9i3I7cENIb3qviFW325ADK1sgV6BFErnTviIQdY
dbhNxC6G5ZLlvjaT7U/k77qncRGM3z3UVrGqyFHaH8Vn5+ZCB0qaqrgJbKxUVvlC
AEOr5Ake596VOPYt922jDeCYRZAuCrIvSOG9sm5aVirUWjuKahdXva+qveMZAQHb
joStrJd8ZqAvPRhpoDTN0Bt/O8mlMJOefiwuT6BeKb9Pjw5mMluhHX7u/8x4f5U1
6EtSNauveEDnO1xa33skdHHFTn4AWyzpL4hFq3L3QNyCKqJl01Ao2Wo9THH6HmvX
ui2afDDvqtuuKCbG3LNFb3w+41YN5zzpd92W7e2ONcTnwLa/ifOOnqQnEiTVox4Y
dpCqQPOqOD+QLMtZ9+sZL4gp/+oyk3/hLks0i1pRX4paT4poBqSmXUlfnaTfkRY1
1rFuxMbItHCj8txWJEYLBiLpPOuc8Fd0M3KqeoOK4bN1gPHahdukiYhTXWpIwZtC
cbuEMCzzWDi4UjdYSezM1EdvyfdgIwqzbAs0Cpnfo9X7zoYul/6I7K+YoR8F3gna
QfgM7H5gnFxP4IRmFc/VZr7OeMWzT6e8+o7EBE48ZZkvGTSIAp5z7CVmBkphiZ2d
0hxH1rbaPFOCrwe2KCjow7r1UPewKr6ME0wo8NRviit2aO6Xfca9CxeOqvrCsH0S
kQAcPhiUiN0Slr/aM3qlFI2n5Nvr4jq2F2Dl9vlHCf1KJNGHXmfvjwJOOLdBHk1g
ookBUS6PMW0FMhWKMNXqoPcZPgBfWUQly1TETTXfamK000ME7ARGDR5fpUN0rnNu
UIwu4IrMdun3iWzM6MZdM0o0EKzxN+9cL1HY2KMqvlCylVB4LG0ye/VLwwbFpMFu
3K6EPaFxYbkNCGEOrpSWORn6k4UWw41RRB169MT+AL+9AoU8rsJ8r3WUcACK4CKP
QIWATgyA2vtQ/Tc+w7/STj4mxAV0pKrY58vvI0Nt1fHm6VT+fW4KHRQCRR93lIKf
YY83ieaQM8NW/CjDNTmLTmJ7qC2Yu2CFo3Hxux0VgryKkIJEzYQWnj03UGqkjhRG
1vnrJ5SRHm4BNBcErJUfClG3X6dDv92lOOxJM9ZKLNldkoCPrQXNxEbWVdi8SZGz
aF9eSaRH2xUmw6BIozIwYzPkc4ez1/Rx/a5AMpQv8Ey8DsTVVCOq/f7nDu3n/zPy
o4VFsthBkXoVJ8vTFW/aVGoat+dS0YT2QidWIBqIwX+LQ4NO9oCEkiCMJPwTlCxz
AMSaB6P13ZqBGp48WMHczM5fS3a8LamogEDQ5mIfcLXdwzYmKHLJxNXj+gr0kt49
SHAWcWUZGuznj5m4x3bSbIEiw/sxe31o13obQDqDGnMjC0sG1JUpgY0dvzPPNqqD
i2Pbf3yPN6/nfl9z1SUFv8t6q31eMgmLYfr4Nr9UdkgXcmchJwlt246CoNyR/86E
NHJeezSU4/qMlEAXKR5L7JVsojfV72C4fwl3/VvhA45AcpakJBwKCTrrMKnwm5wL
PD5P/cBodgWM+4hPymX5VoMkRTXs+aZDl9DaeNja1WMs8HPAZn1WJOC5lrAu4w5C
AMQOboObqyaiiK9QvOAtNIexzYCG+zKYXaQU3EMQGU+XwB/iJDcgKgaBP7o6rYXl
n2F6y4lSxX0CLma4f6Y0xtm50cfdqbDD4XN2i1Cux0tAKbFmdR3TtfXVf/IUmruT
E9PI+WfSbH8mGmrnfYFQy9S2VArEppffNntYeWE4G3WrU3K+obIISNCCjqKUSjhZ
mPrm1XBPHMwLRJSFG4yaEVfZP8HOPA0WqI4YuQnwSEiyyeaXKZVP3/TtJRW+OyN/
baE5mCzoxgnwoPo1U5yjih5JahGx1s7ITwU+uGkCtvfGomYOA7z+RHsk5iFx359J
1sA48W+D16KpqgOCgBvT6Qjqblh4l/2qP4DJIHR+keMKMfo9Q4VFlBqZaYyJllI+
WAW21Tbv5qiBq6bbR2ON9BNpd3TLZDfvOz374ki2rTszKVTK0ILxDE0LOcvYalPK
/vMiA51SqRS3ARhznYxrQBnUAJv7uF1j+Y8HL6EgOJe7TFvRAlTjQE9vH9nPMNdF
qAg5LSeaG5EvywTn91MOByO0TI+Sahh0hmU9ryPobLjCAo4b+PLQX/Q1pDz5aR7r
KO7vRFbJktkzRQ3G6+JMNNY1E6VO8my3cY4elx+bjUq8o8LU2Xd2xO7yXeoIkxmd
m0sXqIrO7uBsT9hCNWT+Mmiz21rIswGx86w/BtBznM6JwUJBtPGHV7t6K+hbVJAc
rCLwyLUl0L6aJnCeW/K4zu37TKtrGgS5srVnC3XPj08vxXGnyLdI/qYQhwxxq0eF
SgrPeTlWRblKMuZf3s84fRibDmXZ+oUF7WgGnDfK3Lx/OT+ULDKquNuORhlI+iWd
iAXdYmjaGc+7NHJXcbcez6wHEvYb7DLtJqawWmsTJal60iB27YJ2zIQp16v41mau
pATr2yPqm+RYPMu5kRUvPMsQPpYHEF138QDZibWlbgDSR+SA++ektucM3wwj+Su0
Ttqj7H4pX+eeBWNH43n0i/d1kLWhBibQKRTaG0wA0M33yRdBE219ZgACwGlB0Ftf
aW0gc9iDZatcywX2IgU/NWrty9SDJ/8TUDSZ0TaHvOfmci/RbUt/396jInP74CD8
t6xcFkmYQuaWrMfroP20wRx2HXiRlOhee2QXP98n2wMlhtF0IDegGqbgzZFcSAm+
dEQ6fHkKSlGwIBDUS5aaqv7Ez9wOHkiCnWMX4u2eSlRO1hNib790gdTIz2fS7dcT
C2oxEKstXBMutNYqxEUTFHVxy+sTp0qPwQk57CY96e/hRkSbaWvocTQpwPw+VMQ3
0Ct2yeYcwA0mROq6C6TwzXFxum2P7NNNXUijMkiq0srRjvtyevhqAU9kNa9ZLLP4
DUOcnPDvi3gzNG9yftzUPIGJ0gtDARUmgbpbE8T6EgnjnG5buSj7JygjsPcyslw9
eDL0Zbnimha3CgWqeSGNQ8bJvKUlH12BVbsV8vBusD6uuyScs0UZlHmHtleS8L2u
pV/KEcVyDB2uDnPGLNrDz2Jzr0zDnAopDbFl3Sp9utqWN5tcqmV6QY0Cz0qB+fsa
iEk1+6C4KlAps6iM35zm/RvPd417yZLk1yHaA+z5467Ut7C+VcHFHjWsTomNKuNP
gX4aNXaFY+ezrK8iPcbKz35btN3m6KTB0WjgL5u1lnaUcLADBqMYJ4+lr/ZGVjxI
+gwU7QNA/DOClOWyb21sR0WrKc/W4a7SiwR01M4ZgGqiIXEm/HdiGbwPiZn5daX1
WPI6zMg1WtouDmZiJGUXWae+eYs8CPtxbLeHGxgtib0xTBFEXnZtiUx0Kf6KIYq3
SmiI97OfeNs3MocE0AkrK3ENKgI+49H5XKdcMdY7q5kMQi0oeYWaoLUwBK5amAug
sU0XjPIgMbFo/7QtmZu/qz5tRaTn0TNxBBQJ+I+Um+ph3r8Rnq5UNKL/1y+jYW1F
6Jm0otW2t7kT+igTFt7R6S62easXqY78cA1QTSn+3D0amLsBWE8eKJKl5d/IkuCM
XszYEz2rnFQ3f3P+TysCkl7FYGe+yBJMuCrjjs3C5D6qaS8lRdvOTe1M5edwbUv+
Omn+bExdewBtxp+VWIp2SNn2yeb9nuYSyx69+REVIBns/IVejirtoRLqLnUN0EeK
jz+EhDJzzCOJNxrrg7RP0cF9KVSWYxIFm3DT5u1oooa6sUodnGM4UvJtJIUjoAyd
+o6UipvxMpGSj7UPg1i5xZkFymnkIPjzhvgCINZ3xIoMTKQI25nL+uOI+pDq0hXT
xVTe/T31g8N7amqfKnbgEjln7QVAlrIhxjlFYBX4kFSaaekb5foNjTS05Ko2rg+u
CwB1lQGxwbEq7sE9EtkX9HFXM+Q3DCHD/7oY4KWOCBHIVZLDXYCkDQuDsB4ua4iH
K2pvvJ2iI5LoQ1saPrT26zuXcu1S+0QOoHKGzQxjTnGuBkM7BCJDFaeswaKM510T
JY3KuHhmjP6xJShSYefBsksMst5CeM//3prwxl3zQYjwHY9r8PdOJYjWxmjyF2f1
FO9+asPtGF0TVh6n5ifaSaWfwu/0dPcLuvSSmVQIqX0WGD5+HMK3HqBp8IBz6IYl
ppbhXiNuMhq0dc3L4xo7Gls3SnX3gA5VrxxUHArytmGS7dzSZSs0WamGZFDNBYp7
bwx6dXNkSY4nIp40wmjpSk6+EVXRqiD6WtxYBhsbI2kUK9n86jpOionnGh5qZ6ZT
dsJjdsyEyOmo4L6BmPP2KKEv0YUCzVwXMxfYIo/C/cXeFEuQsHcMb5VGIiNQMXE5
3JubBBx23jhh0qPySPC5rBuvp8+LGUbmalpHSl1bYXSTT5UnJKUOs22K+oYmpnFY
z7WFAFVduePvORffwXDrM5DE7ywGcsKKRq8ogbRK1mXKazFEPYXNK5lNGEq8mBdb
FOGkPeHifC2ZtRJkBPbJq4lfQWRERwiOgMdvxzFukUbgSzvPt4EVqe8KcWvB7oRC
vFmuD2lrSwumJ6P3D2xKMLS7+LGAp7kjG74p4b5v0fSxeyvpFosQfWis8Lvwo0FE
rw8NgrPAjWkle8wpaiDgBNukGqfzC1ZoYR3gFkX+iggHw8GtkljyUYjpC/hAGLgh
WTh5t31yCAN4vq0t9pT+PRGZC86R9TZUzRgUvi1b3TNp592wtWtzcJF9Rj50hXh4
nyzY5IcyNQji6hSnTb7gPDeR6Ya7DJx7VQK51rvJlm8a9pU62AdVlr5grSlYsRQT
JHqVlHPihJyRblOSVlvo+4swPHi28pK/LJHxlrGbEF+Dky7t1dcsneEtyK+DN1IO
SdN6jvLmr57kHvt9KtUp7Ix5/v3K/BTWv7oiyxudQaPZeom723ZGmrvrmWgGgsTJ
4qGouZXp/7GQQ/ITIMg/sJb9yBKWh3Hzo+IaFvahX26no9vY7CZZviqwL8ojsgbI
P5kUEkGC+crfLz/VmYWHc85CQaanyZkQbSoHd5ikPw2GPVfw/e9+EbKQfnv7qeYh
OTqCG/cdCiGHh9MFTold/xOgnCuQxxltG7bEFdM1GFSPNt2f8YtOEyiRbuogiJGe
PVX71Rx790nbNtNzGleRX6ypPH6qCgEZfeIvCoGJe2/HMUBqigBlUq1X4nUC57TE
/yY+dgbIvyxDAAUBskXH/do59wo+mzjSjV+oiH8fOqdGgcIeZakKBTnZ2vPpfefj
aHl8wymGfQQClf0hnycNNDSTXjti8TJ/aPbiCdZ+EZ9oJ369UN2vScrJzAjO2ugo
hgiXyteRZGP8gMCYZEWPW+vzd3b1NzT65BuApiCmOJgE6SISKA+VHCEsUCxEZKAC
FylD8+wQPKW0yKmj/ZZgelXLvGChJFQHRJPdB3R0JpWBEirgdyIEbIf185XCGrR+
UWbh/8hcy51QCnkH4dil4gg9aNhYZfj4BlcjBtnq4rHsR/iKCcX2e+c6vE/S0xSm
E3Vos5uC0uERCfjhxHpsC6W7McVLccRAb39q/u5MvQ03FdJ74ASMic/bwsLc5hYI
lgxjZcd6mqahuQRVZF/LBAt3wHVwevMKn/MdvtJkyTn5rVe9T5szk4S6lihkpGdo
8R9S35IzgHXYQV1ySvMJ1C+zW1nmBrwzvGRHeA3opoHoS4ilAQZJ6KIw0+eL7qMc
h5OnC7CPmSPL9CkuIKjk7AQM4QhFhaY2SuXMzN2H9+zLqVBJrCq9h3EtrENoVqzL
CQaV47aJjtZB4yiv0QAtmSd/V5io50yeHT484jYYBWgn0XptTRBRdb5zSUmeS4+L
n9fEJOOHwBy1Y7IXRjn2ZYj3K6ihHqSRbJjcFWwLsX8ZMQUUaWcVnB1s6yYQFhP1
S/fC9jVMrf08dSnKJ05Zp/FSrsUzl85p5OzdURFfEfIjmlRhiGzlFppPIq5Gokq3
JM0hGPVoEL4jwLyZzzPpqO4N/qlZsbq1YHI8/zL1amKfC4J5q2mQxsxBpPKcMlfw
FAtU6bGpnjONRHyWDmxfbEyrmhNtEgGu1p2KdvRaAKdgsLoTUOWJoaLbg8uDttKD
1MvevVi8mlbH1kIdcRWhol8AMw+C0GQP79F8Hd7ODJODbTyKIbv3Yg+erHT6zWCB
zqC1t+X0Ssa+RzCGRcpkQNUPm/ZfcmN/3asDag+bpe6jn2sB2w4fGIUmWuRkoaiZ
fYcQCUdmJl8gtFiwWlEEqqTu5HkwgSGxP/Z2rI2vXg5prF+RbKkzYYqaQyYY7HUa
9JSqfavFocqnAxTkF6dJLKcPmLmBHr6EiVJpfQ2/pIhGeEEIcmlkg56nSI9RVnca
jrx2A+pSa12sxw9xStbhpN13nt3zrOoSSsE1Oa7DrFOJgvQDXMY+ifYeTsYDqqdj
VoWD5EvhUv0FQPbUpHbscWPdTDS8/MEEZBOGjC83a9NBTrTSVdmXVY+z7T7YZgyF
PaFh1L7AX0w+Qn/haQH/aKi5GtZKiSgRyabw5CgM3R7dUrQc/XlLDoV6Puan9qSW
2xusaEBnlSPcRGlP8QePnXUVJdxu5DCOnyKPirE0+L5jCWQ0mQg0ZBX3o7FfL7o2
2oIWLtRjHi7fvFyOS8lsCPY81golJWAe+44/yqRtyXEYRajCUCdw8020N57fnixx
G6GdKiMf0C0oqOKyJsDZKu20gBZOt3Rw7DkNXnAoXIATOdGT2QgSq5be+t5pS0Cx
Z3CgExh9pEnKne1uPHinE72/Y2guTxkM0jkpsSk2l4icpS0NYwktH3TbCt5I/nvL
a2GZElJgBQlJR1KIhwukDfwVYgWIjZzEsHLo0GEizu/tKv7b4gd2RuoNvlHGgnrj
KDC2irU9Nt3qC/R3nqNcLUatFAV8IEuKEXNCBrOStsCwNfTEZJOEvYDI+5jjt2+U
PFXPjOihniudymW9hWLa/iBJfChX20NDbbKGtKTOmbaRqkfn0g4tp9pXkty2oVDc
R6EwppqRz/mEqNVJj17KEh9NZTx0o4hdK/gIqBwQhM7u+5icwrKDhZeQhcoj9Itp
6rbbNF//wvzh2xx5vmIXhRC9i29sRl+BPG037LJDNQ/kJb8uzU1nCX9e0ujDg2Ac
nHWtX7Tj6pNRpwsBZ3lNhW6BK2QQcWaRtKQMVXGdQGUeXi5xANBUbxC6/p+ug5qb
fn9H6hWAWjFgIWO232ZYMhgZH3eqvhn6xfvx/DJ4RUlMTTKnVEu1Jp+Kt9YGacY7
150kkc1QW21Q74iN/eUuSPHblxybmQt21D4BdQc0oCbQJHuZuSwwBdzW0yww6/YQ
NzYsRmbOvYFETs9c9bdZP1P7lwBZMmgI/NAfDCpOFUplJbvcWFoyb2Ly3kQorJON
eQRsrXBYrV8ZrC5QrZmnx2XRYsMOlL5S/6V7hbDZo52WgodCmTLM1BAyHsS050sM
wNpTZyDMn89JjrvCrG/JuLVbz7WKW3kk5ZCgRpwGKf6Glm65mF0yB14Gj/rL0vXp
Z+WjzMDLKjO6y1nUdqmnwkxQRqn8j/cyM2PaQ2zVrlfDu0qDQo7dGVDPqoZ5RIVV
Le35vVS3z5ZSD/VfvdYEY4FNrNQ5ORhBpXkv2ccZv4FZMHJcF87sposrkyB3W/Yd
ubWy36E+gKUaU/YgcUmGYeBcsrcmXOu4ydofFyctNFnMjoTMMKAwJdLTtLDhfnni
eM6BvWXHdXNrfYlQf5IrpBL70E0S0jlAHvNidaAPsCIZMNLbkWQfG3j4zrD9YKsV
pWEuiPOLiKjVJd9bUIN9spel2UqqrK2QjqCsuLouogxLymiBkWCJX+jgka7tBaaa
wHtWAloFgvOy8t01fXxdEwmyhw5XNaa/+UqwVQXRjDdiWqCS+f6EklXzI6vasjqG
iLbvWTfJslu7Gg0K/2WOo5LlnPlv8eLq2Sw4jQKQo74Lb93WT9v+N8VEb6oXQodF
DDU5m1E0GAptHxgq7TeGNXFMsuz/DCgCMwOdbdpPkpGs0/Ah91m1LUsHmgHwaarn
4+PKX+L/DvaLK+hTdRptuBXdJoE/kvlTW4R7GDlS6RiSmE5+4Ss+s6uCAPvZovD7
CERiqKpmDt+2lA8kaniJjKQb8nQAZ3238dBrz4ahOf7a3cIcAvtmPMeGs21KKEd5
TlWBHdRzV7jshAKxuwsgJYr0E9jX1gzQIN1qs21cUApynd1xqUoXarXtFWgAbaa7
BwK81yV/NMBkd2FjqC1KvZ9UzbInx2XdyNb9S+GfxzkpSfj5vPaNZlDUh4Bv5WSZ
b4BHsImSkfhsFRe+8vwgBSlt6VDEvjumyCR4NOJJCUyeassbOtlDASoghSn9xAOc
GwjFfnClzGn4S6Hj0qmdgZgb7zf8rvmoyILBOc9EQM+KKZ9mIe3Gv6Xpxqffj9aV
iJLixNuarpZdOfazUN30T5PtsIUjVxrSNDmbV464ixDrjzMm9It0sqJXrv+ZGzYg
FhUm9YWXvqHq3lMMyaqZ3Iu9SD6PQmhxpJihlF6GyOgMI4hk7JltzABbwBuQgdNE
ehZOq9fTtsj+I/GNOyIJM7QCHu3oEpfYBBA70ibhvXcEjTSTXm1lqdqEud99U0do
F4FI6AFFdMsY9QnT6fgrjBfLEqle+8dejkc8ciS78y8GAzL1Y7nzraR34U+9hiZ8
QWToHkUZtVuPS68zOnKL5Bjs6CjAKuxSAftIuKSD+cpEukzXlEHZNiriSEahOjsz
gV0pyqfsehOwTM57B+giW9Juv816w1UdHcM9rNTxJy7vprHA/gNWUZTkLnrXv7M1
8D222j1xzyjmruRqPwNjihoR+/HXYlUsu+1LzFSNhknPPSi8+AHcBZhyNu7eWNsy
pQ9jHawYQeFIv6hdyoan+Z3nxwtZu7GhoKAEcvyZf0AIoeGxG5epdsveydIV6Bki
dG9KQa8NbGCAYf8p2xXKRRwMtilwW/27NW2+CtGLrqEq3pVGEzh7TFjz/ZCmznJe
Vkbi8noRSkz1tdf/KV5+ERIrIu4luWiMRZygBWd95KZTR/jU+nmraC+rSew/JEKL
hX1WRkuRqlznNQxBPBxE1BgrWiUN/p5JQrZXrJfVqbSujxjHTpO692+bdVjV4T5q
4OUpfCC0zwgqQLR4VFTYZMyF7kHaVm+b3yOvqihV7AA7IC5KKUMKiOACM53Km+yL
DDc7EQR8MDp3gZIr66q9zQXgxn+44pHTvN7G/LVctPlJEnQmLblmhG8cuUg+vrl8
HDpcuTAcajYGCn5PRGS5c7CSehBaqTVpAjqycvten2fa3K3fioWXAZPHGaJRcpBk
tY4zubPlAnRILrvf9Ig4SDhrvA2B69O1x3AfPurj8a/bDUPyxQsOEiVw2eInFr4I
aRWpDfN3UviRvEgScXfFt8TahUugvu+WfL/obxBv4UyW2iOX8b00qkMEI+XuzMfF
Ch/CUwC3af+pgTXSvg7N4oRo02voTn5VUkvZqdfaHrBM9Hm4Qhehz1tt4uMh2iJU
P2MRMK1gHZFMKTIIN8+Rs5FEZmhcyCb9jiWX+0LgLsLhyCdKSNkJHxTSb/nkC1Jn
g6h2pcj4s6gJJ9q+457+/pW2E0zYV5JDdT0heLm9aZmVAa39JAP89E40PyqN0Dim
beGHuVW7N1E84GTErIzg2uTPbeTPc4XXKKrWjco5GvoE10s9AJb04EfZOvVOOrWJ
h4YC4oGZ4iF/dYm0gJ8xAVV7r0nDc5lVq99AVZ++JIOJCciM1aHqDpe0bcSTzKqg
XFUedn8eHaGY1Cq81lsE4jf98TWgBY4QfI/UK/0fvCWp8fjX9nnNl3IKOWpNO1ri
1sTO3GwU1S1TFzBMqrek9aBIEyxP40aq1WRYSM80b559rOa2ePJEDjNNxgoIMeNr
WZ3zsiGHzJZZXe/hRVeAFNhb/G8sFWRSwrIFu8DngnReQ38mVX69RjlN9W3HUALE
OdnD9soW5a+rCSdv9oyS81wWEFTgqls36b1wIv3jrbqfSxoKHkI1zOb56psASwI/
V8DW03nkYj9rvqK/PcNCwKLQf5B8f944BD/KAch3m5gxpfKT1eYvW0K6/CaJJIfZ
UOIk4Hht0gY8mLywUglHPOqvylayPvQ8mHhh+6WwJNI3l9+ZIXNSdf35Hu0btIrW
MYJToC9LODQPIfsOaDhdmM3AZhzuHCAc2fRoadCEbKO6jnuihI9/k3A5HHZAqpZJ
Bx9tPKAYu6Ii3WjQ06MQ7MNIaq9Q8/je6skHqHaUU1GT4daC1kSEuQGCSYhBmPvI
tBOPJxpS1mjkyKehHLtorEecdofZ6ed/1fohojG57RU5atGSJlO9VglNVCKHcn06
5SzqNnw7PRXZ0+fg6HZW9/z4OcmwuvIhnEWGGn1p5mhHCpvJTf0l9yd7Ox4PbM2g
DjFv/WKj7Js4Mj68JCQF+tM/pXXaawe5jds7nHfi79ezUWMrTDG/5Y/iQPDpK3fT
hCnpnCGyihkeW5hqE1mHI/WHdjAWXSH9dlaugA0RDYmEiycKjPPRHNdXfmq+Rn+l
NDOxlpXEzTV5ucwLhdLNOtpu46xwISTrfmnJvzS+Fw9VBvwPYuOt2mNOZt2OMeCQ
GfOJRC+DwAjk+JgB99vnzUZWY0cIA8rbJjm6CrTSlN4i5422Qq6SYNYrVW9PIjXe
8qer1zjDPyfaV5702JXLi+8pIN2NojofZlysWjDJOZgsjIg8MIwkt58MWCkC7l5d
NzVusYQshjQ4PfcskljqYHCzzpiuSE8U4WRKfwADu8rH/E9jolpfxbevKvI2BE9t
QHKpsOLRCNwX1sUWPe8U9ljqmj8Xta6dUvfibjdwynyZtQjWVGfTKz09mGhQ1KSc
6mjQmIcEKrOJI7vZOgJK8PVAOdaTauTzoky2z171aF2XR3pNLb3NpBa/reqB7R8L
jaZ/iHON8dr0dz/bAME74wUioY6fRSx/Mv6/QhnNkBOe4aF5rL6WKduaergl+9od
PuGByPD9eDw6Okqnb5OwpmVC/ucbatpnKnkw6o5+UydmslkALJH+J9rGQvNt1ITr
19Rha1Y9GDj78z8F0CJmwTF3anf0g3tgpK83j7Cz9McMd/nDgvGaDf/cDOoUc+G/
hjFX6lPMwCCWh2nhTfhHoFzFTaQ+nIlapVga8qVjfD6I/DUk2fOgTouPny7MkNYs
iaNCEiyKc3kiyQhtMV/LaurnwRE95CsCLzWUFUmnW+6WhGwPHird3tyXdK9r9J2U
uHf/vn9kedSXgx47bqGHbd5thZr+thiWKfeMo0Vk7zPz4qKzRF++Y3INXLDZJ7zB
15Upq6fOHi/AMA4ijx67ofwpy8ArsD8nv4gexTPx3YTje9Rh6iXfE/olGA7/ec08
i2/2yQbQq7VFROFLctxyMY7Jy6AFCeO/nG15SzUoeynya2XlgI/OHx7aEjX3vDtI
J0VfQn9LgUsR2ZNC6Bi0jC8hGlXMzvaHKlZPr54mzmrrh44dBsffUYpWsbbGWN+9
83/ZWhJCAjhthPj/mKqsoVWTMHb8t+2rRLeI5CvmF2n3LLJ5v5aYBNhEYQCC97iK
0VZNhBRhM0LZ54PxVLQMd2aWTKmZvlmZhcyIMIFufuu7p6WoFvgI5PwAuAYfdeRh
OyKoh4BAEKKFPCUSxeMGbULiEo6NE9VBzUFxVmLYg6BdNgXcNaEz0uOQUujDdI/8
NfciH6U61CqjIsybpP/MQc7KXnYbt+7iIJPhOL6nwrPWOLtlzDS+Q7mYjjQIUd+u
hQ03Syz4U+IAPf1zd8twt3jSWytr1SKoE+f7/S1xGAXhl20LxcjBps02ClE5kLw7
yXk+Czm9t/5pOxiL6iwcnUqnm/hChWXBQUz/GyMVpzFFbiseEszec+62m8zOlbPz
O7HX/yhBbCjqh3yRvWkdlZjEAJxg2Q2q5wrKr3gBelyBUeuarpn/JU1vRNr7eS0h
YPIZVV+++r3vhdNTMYy0IStBxmW61Z4wBj9xqV8GPT3Q3TyloRgrSmM5NeKbVIId
czhj3/76Ff96NzUvTuSYIVtDImJiBTkWTVgoTv/AHvB/y7vrIvIrYa0McfsFljKV
0mx2nmLiSdznYS2o8YOzV87Lx3IJSx+c0IcUCHP3eNA6VhM5T38TGXPYy8JckSro
UY69YCgq3RqYL0lc8o6cSVwKnDx2Vo/SQ4FgdrE1tTDGIxJ1M3Pq0viQwmzeTSfj
gh3xNENO9ynCT+pj4bY3BunnhbXI/1YA7WtQPeBhp/KLpHmuuIKnKjU9iiS3PkJv
2jPjDdvTeZRbi5whlsn3HrHLGmnhyvoer1OC3ZI10JzPE/gHXizu0IZQF0fshGLx
CV6xvBUolAUuSH5EpasL2Y062eQH7xuw/Oyu4kgg41kWcY/mNNqXBVaX7pkJr72n
Fqo9Km+ErkNV1bJNHpk+FUIoVnDvvISkcw2aQRyOyFrOP50j23HtYrlAWFHDo8lq
NaU+a3GK40dtTPTemfKQwbJAkpVfA2uUiJMnEWpyFhn8qI2lba0NbVBqUB8apNHZ
xlR+OHN3w/FwVjLFqs0Z2s2JBKEcYFCJaX7STM66iJSrqxPYunlrBpeJMhXmr/kl
CMVmEwCWkExq+PkUfpyJ0U4Vjv4PTSK7i/ZUKHnRze9bxzcozNZncGflMAzNI8hS
PDrh5yic8fTcdRE1X3HKKeP7KVUK+rmti5sP7/ZF5TstZ0WbZPdtvUVNmPWziXze
/20DUtHIjbo8rxYf4+u/fYuGv6Jssl6fy4JE2SFXxSyD8jZ9+HL/e4wmiDygfo8a
sjtNsGt+fCMbKBaSmI2fq9RCbME2x2ylMGbFR/QKKly015iC/3uFLETahIjVvaYR
HG5ULINK9wRUd5QreTyCt0uS4wBz01Fz5vT0pTmCqGmMsBVlIYKfrwzz/pZ0lkv/
xx6YbuxAPsgyf8RF0SWA4Bz/be4dlxO6oAGUxPEDwxfmyKeBGeocpgw4MleIyhUq
GDXXP6n5C3HE2ruv2RHTkHpahSQAs0ptc6LnxZF3kc137QkOCCy37xLu7goOq52x
Zn9QKsQRMIPth0JHXtTTNQ4BQnmR/Z4VVohEKlXmhrapD16kSb7I61ux0c8391rK
M0Kn3UuV7kAfhYpRyto0s+kS6by+L47uSHEMJcKlVzj0AEI2n5qz5nDTZvRHYm+M
o4GzJWTevP+LK5HUzK9WWVALwUtHsjQ3RHVL1UjCgzpSR8OaBJkR/OApJJ8P9Fds
n6aWadMjO6KWpN+VXvpGJP8i/4OtA+D1qZATrQF81Ruhdlv1J90MJpx1AT7owJq2
N6Dxs+wySHNpKEbclXsw22w48BynnHjR1ESILsZaP6nmExczKFZQMRIBXvuVv5Qd
9mU5rJ9/NANLQxLxnI20IbbeXVSve4ctlKs+OgyVxjC7/ZPxQhsYUPWlvYFrXCY2
piPh+8YeDpDv0OUPwe2401/hD9e0Z2XJs1klUDmAoL5st8TA0P8xIJ9KtBQoeSB4
4tMd+E3wQBRLcJoyESKmq0VoNmXbyjRYsjw+1Cf8cJHdfXvOwUI1MeIJAYKJ5c5P
Ddjejx1oPEHEXqWGmzH4C1Xe/OvF4LmwBnyO3U/4AgVUQe3DAiedl/U0JHAlbmnd
8c1cdZmYfWExNHDFCBZXSAvwsbHQrvvbxSdO+EHJKNTfpPMtmLQd0/XcNUK2uMRb
vTT+MScwJzCIsgFNCW0Wofw31GhyTweMAVmS5iPyfmBG5Hfwn+SwUfIquJ2KR2r7
3ly6Zj+oTNX/Vfl5/rxYNrRJFb0+7A0oRxyf9NvMoGX9mTPZGG7gSfWScfaCJs+P
Q+QzuCVft8VmLMA9CZTNWv+UFfjA2YvEREzTG/mDpQoTDqEq2KEPB0Z5vb6ZO1PY
iwe47jbzSgMM7paDe9pbIR3OCkTTxjAJHuz2kET5mK6T+IZIhQAMt1/xxOrwvOox
O182KPQAfv9qapkLytOLZu4vxigiJA9Wa305PcqCHbOzkm6RN117Us54Cb7BDdqA
vOVlnRos35bp1WolXbayKu1edArysyzL3OKF/T0zCn0+H7J+qw2medLHCGv22LCN
KjAv4YcdQGbcQaEiwrWIj4te6mIS7xgDbCcNrej3XQyf/ppqZIeSvkY6Z46IGgVB
tkbTQvdmcZC2mFM/gcfVBEY6sH9vgUh0aDPhkmVsYXxwwSbQTp0l5Hk6TnuFKUh+
xqWWPWDXaCUBYIdlIOhq4JrZGMJqQE8IuJJSdw3lrmyqqg9sinIKS/DCZXpKOjfA
FkIhvX5nroq9sU2VWf1N7JruVqT9m9l3g5npB1EUba8G+rSb4zA3CdATt0d8Gmuw
dVs4yvdjzb2hacOoULqE9d7IBAPBD8LFxJCYXVgu2unDxn9KpXk3MBabQx6yPz59
0+bNDMaQbJQTDG/qJZ2TS2qlfBclnveFOXFCWxvj14SXLcuzp1+Xvauw/a7R4oxj
1qQrB4uRRYrPpg0/0N8tfAjKnHPrXayr/Ad2cmdyGaK1svjm8h+nENtMWDLhhq7F
6/2EZ8EdCYv34Hfys7pKwvc7m2Rik3g/CffYO6dSa+FtSeuWov0+2FbnkS9rXfGw
w6vv4r8nDzT+uMZMbkM+PnqOUV7/NB1hfM5KPcyX7Alxihw/ZBkx48svscdxk0QS
wLO1RfzMjvF4oDMZtk8MYHaiq6iZzZZAvQrQfzah3WsPTLw8SUlByuEu+9qnOnjq
qufxPxTMDuTiVvrmykK+8X5Fg+e8Vfk27Cvot1YTs25Cr3tHHqlIeRSNzrJlWLw5
75Pr1DKZDVPA4N6e/BW0LKdEpbHlol8w5IEdmsuW6D5kFjrGuUdA4zV3YoIoX7uX
Z7Gc+zQvdx70WUbBz3K52vpbKqVEkN+e4fClPscYwJAWDqmBMRuBGzxFTH0OKAW0
dflNg0gOAHv39jjaBNeFOCAs4+avTrgXcAoHG3lgtSPnEeYNIU2M2oksonFTZ7hi
BmomtcLq0GcPRyUd1AJDg6ehzbLQd+BcSylStvTibJH6qLYtknzYFHS+nhe2qilH
fOE9Jgh6Qy85fqY+TxCp4JzObwPbpldJipJ3TET/WBAe8IP8aWTOJAGAGkY4l1FN
7DzWFDa1awUUP/eREftiPHVytWTHcGJiOC1caDoA8Eb4xAdjPOuSxbmqgBR3yHZO
Gj8VEVQ2x6dqQ9HQQmnJYFwLUFWFVn83X4rzlWPMozQ=
`pragma protect end_protected

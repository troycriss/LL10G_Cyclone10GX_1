`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
pJ9IUhmVe8kbtXpLN96AdxZ4jESy3lWuNeG+lCGNWz67YNFRhvn0wH3a3NU0nzDz
eer9iORosVhoGexj6wdL3ePB9WbNluKGDWLOdE3EbPg+OCFX/VkAOLlYFFo0xdrB
kVCGqntXytUH8/QpRT8VlKchiTWZ8q8MjrXBq3GhUjQ=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 36992), data_block
RtdMSr8IV21lnzqq679lvF8lOyiHLM17E/kyIwhtb9/MUxjpNMZVcqwCv4eL4GlI
JsYpYF5NHZstTPA9YFx96/4U84uqs7eHh/Xjqor6XG5MpctFLSGCHk2C0RVp2+99
qzmPhYSse9akHwPBgbeTV331kDUkcNUq9Jiem2KTtFILXapK9rZ9vOEaO5zVh2qM
fWP86gNg2FxCSEfmRGXhdzx2lyrPrxW/F380+U6qGw2ADuLRshLFBAVUtya0MODG
LhFJxDVKJ5Ihl9f1gX2z6WHw2iUfNW1vqB/akW8BQJjIEQBFT46VyEnH1p/DSpkh
SJluN2G+48Z5ptfCe1wHiWpngn53Tjw5zeIY0rz/wkNNeQSisX4f5W8lS+2DfcpM
DwTGzG7KKa3gp93sYInmXs29W8B3KeR36eIy19p3/Cru5Aije9kRhmGdLHmqoCBx
xWXGByekT6S6LfbYrWg9US6sJd10sBozUzHKvvCzQVhUtsf20BtqWnvEameg1I62
xwi5hQa9dPJ8EK65wz2skmo8VvhvneNoEzZfwKQX8O9Z2v5FSQhDBpanyLvs4NeY
8b0FoGyvLhdLWwLvazqaCMbrcFyR2MdlCH3+fLPmEoLy7VXe1etLPWo58oTITCI0
VW33bJJBi4GmpsmzQzjMOZlpTn9nVN9tdAdk7cWWZW9KfGkL89GA+JolYLZPOz7j
4ZQwnIbovv9aq7lsWxWgmKo0e2HP1WomS9T1+2kFpKCFL2arDdDCD4s3ZfuEwohi
PFNXfChL8VdiQc3W5HFw18Y4U/vhvVemGi+O84WlmNbzkQCMVtmEE5CWl6D/a6mh
hOLDi17uzzfF6H1JXUSHsYUrq3GBFW8+uNOHKVzpbslowqPdrjXqAJ0XVsRCRp6a
iJrF7qPU7mOu0Dx/XM2Tl8QRuSvTa2i1RoPmAJIbaVuIvXAidjEnF6u1iTw0SnB8
tDaL2rJeOk4kDlbAmHXcYRq2D/Zbt+6y6O8punJWxxJvZ0cBVpbE73K70mgdY2me
uZOXczS7msPMa8pWb1IXWfqFJc484oX0Txm8FvHGztKxGbtywvHTsO5/CcQj5Sn7
23PSRnRe3f9N1tYqtOl+JWAA8yqhWSiH6s6BiW3AmiZqpPLQZlVcuiavy73LBgim
3+0jEXFLRVBrJUh01rAvfvmvzDXrmkPk7Sy7U7Od/0AUG5+sQUgAeSw9JzBE0Iim
us+CVKLjArjFiVj4tspXfBp/QyF9FiyQn4KoH2WvK0bSjXuOW0LWNN2AnKHfk6JY
g+MhRJrRUVWcDTPjZQ+MYALHcl4DuLYeVzgpChvBlNV1AKz0uPs6ZpXBU3sYojWV
TmH4fwx4c7bHZ2IzKN/6CxsVcNvW/4ciVXTA30soh+WXYSbm5yHcay47ZLW6TAQ2
0qfY5+M3py5ffbpac+7h8jHl1R6V5otCAj2KPJL26RD8t352WZw5OVkqwyRqFFHc
q6n1i3xaluOuid96Xtgzbc3+KQrPessq0BPaY0bkOl7PPtbOXJ8IE2kHDo+iSyz1
euTZgDctqUTGBv+iC/k+xFrNq0A/BALDxkA7r9CSku8aHn29vMtFYjR0LsRp3aXV
KBoj0H+OJkna3cGj+8Su8J1mI344mAXrOZo2S2QSBmTTJPDJ5ZLl/QugdEC4xFZ8
rifP4Iqz4IA9JJTm5Vg4/7ccQBZadWP0DzH9dZIRXUIZjBd25IGBcs2SL5kBMgvT
TgX6iYGbdktClpE5Itrav9GtduJFQ+H0F5xrWGGwX5kUROIbtMnGKgV5SAhWU9IT
V831SnqOJEcFmSUB0W1TNErZOdBDzA12h+fcTbf1KIYLO5QkkCsvFeQeEFLIUjbK
BUzs7Bdy3ozvt2yklxch7pA6T6jIPRKHFWcWp15ihFOKoQx/SLk91NWI1CW6FlET
uu1s/aC+xv5ZQNBwvu6f2hnBISXYA57Gu3XSlF3BGeKyIOAOMK/mauDg14EbRon8
hVBu+/p6xfiHwo/god+lC8l4Tfhu6Q0oGqd60/AIM54SlYLD5z4z1JQnhCxHolGr
6Yn9XsS8aRqoS6dMlauvXBV6eOmYuxrPzu47202aEVJ8a49NJTQCKzDUBfaRP1xu
K18yJvn526911ZWPqV3XYw9yyYWnnVQY28R4lij70dFWsu9lYzymFrMHRPnDs+ja
qpcDK9fTHwFzU3N+Y1jIqiFr8RAtL/23J2gWsTe3YIsrGMroSMirE/+7OctCHyqp
xbtATRm1mwTjL3mIw0fK0skrIm8avg+lF+y/OxN74gzX0pqVbC2uIFFKeUF2MbO5
Pf6py9/sdLlEOPXlJwJHuVy+vZ0fXDVtnGv8vm6t8a8LzST42ZYEbFjUCAkaijv3
wzgm5axK3S0R02wlHYIz+If1qWckRpPmIlp6HvSBZis5yV5AHas2iddELUgW2zz6
JptGhwjfvAZZNcgtDCX6huvug0IwilTIAyZVQck/hBe7J99+Z44kKLFMy8mztV+D
9kU3myGT0HYWqTboYRpI07RjVZ2YVgIXxPxUURit4t0DcMIE2oBIH+rif7UwtzHF
SYJ82nd6pp9vIQlqSNzYcxm9l48kX19nXNCqTNpgQ0hgPfvH2AxuEMrxVZ+Twft6
gaOOaPpok39kCvd6+gy+JIm2MPYeMd6AOGpCn9FCubbXUm0PGyP5MEwYK2aYq8Gb
ssDX5V4cHtXVB0CkCwg5I0OVAzK0+Yuks1U8q55oPRNCscQo24NVtdivDyohoq53
k80gqVwnyIIii8wGuCxM0as5ML91OtSoE4ZYqn06RXtDWN9BWIrBFJ07aoWDG3HR
CPTJainQB66tWBBzScaFz4OFPP++omZxrQ/tplgFYm+9koPY3Onxr3qIABtNu/0j
QKNqG03fcoYumRtQRau0mCEd83uy46GWMnXCqKxV3nsvO2TbNi92ZpyyoNOibJsO
03UHjIGqR6NjiD1GhNV5XvphBbCQiI+OKRDHzC154d3GZEIz7+9RE1xbbJ3qbvJn
I29/E5RRWi00cBz4mTEKjbkJ/lPM0SMChGEe1BJCml2CUecncMmxu6mA9PZEKANK
RMvkSlCY6YnIicHBBWViK0c6jMe53/yGIHwdZzCASncQt2RrEwKfOWS5BD+zHb9i
+Tx4nXdpF6jWTXAvEYSI15mldA6nIl/JVM//X1uo88SxaFHthgkzHvHKu4Omon8T
lpoib3YW3q8sF2HtxSatgTDIt+r5IsEgFs+RunwDvrNLkXLo5ZPQbLZ/gH5cQgcs
jq+N4ODtBN/jNNCGiaGHELU8/wEvLKTl80ojf+Y+8e5KDKI62ol7r2vGBbncKBcy
y6g/qHa5zxQ+LM8HQ1sXaQEK4xGIaJwedG+Rt44FheeDODLbjW7ahMwHyLlRQGum
fqiVbgzK6wYFrSOQEqbNus6osliViW/RoJqg5GVLOzi7NNYL1fGSGx5RJdDTyUmC
Gnpw3m82KHp4ueSsvQLhulkq/PPHB8w54yjEeFBhNLUVKvQUU/QlOjB+mnIJTDuv
d3f76ejsNwPQIQAs8MN4r44bbx3rHjCGcOExq87QpB6FRNHJSFIMbphs3L4sH4eW
P0iybjiOn/H/a14yT0U+zvXeFawYWdH2Xyx1dAeFoqnSbCcZ+y5U/2F1XIqAKuXB
nQB/5rimH3e3JOkSnwYSBQgEVaz1taah5A+g/4jHRBvGVXaZCQXe9LgxMJTDDmYZ
D8bfcEzhzZNHqnMyL2TFyj+Y66z1q2tWIgMbTaLP64uZnWhIrNvEQg9xt1m5qEkL
9n7eXavqKeqsMUKi+IrfDXHz4yH/Gxag/srqxzpKg+Ddz2u5tOUnV/oa//W2ySmm
OaQQG8cNaH7ttmLRE6VmzGWBdpqDITGUCp+/+yXm3YzsgiH6A31k9aDjvDa+e645
V6/qr0AXGCEmyL0xmVifXopPuqH0CvQCZp/MInwiJ8/eitHq/L2vV5e7gZvssyyc
17cU2WRHyPfAf3GM8H0uECRaf6XaDUyXdwOuvJY0G/mFHjV6NEdH1VzTqvvF2byp
mbUQiqhvW2iEf8EL/Ad48uaUmxO8Jq3nOVsnknznFuqHDYNWhnRFxNd9RFjLNCW8
9EaxuaULGUmGGfGkP1jQPOY/rs6CRNXZL/P5RQJH6VsWE4PHlKFkKHFA/69qlfwa
EhA4Rd2CoIPKYq+dOtEKf2Wnt0mcncG4KdBlwqK1/A+aLpW2fqY/QbCSf84mpgfP
x31qDBkecdY6UIspcviohxMy9UN1hVmw7xiv84YfecYDZl3tlOA9M185nQyc/X/R
KDaPYRWdmyqNB8YkaorVHmIVl/j4ZAdwYGuccMPzC/MZ1NgfisRMwtzdLA5ep9iT
AING4vxXEq8ieWcSOSRUu7Y9UrQXhSAXgAcyY4vjdk20QtwIxzoPX7NZfNE2g+Vi
fylSiwg7r/i5+1hlNeUWjnFLx16glE2Axz+Hv+Dj/TKmccxL4AztnWj/S+xTqiM+
iO3H46C0D5ar/hn5Z7Bc/KqJSi+WIB0XwuSxnJ0zThVcemPiW8etna2y4BbFNuKN
CNhinv6TRvelO9WZPp2zjcFS9n0yMSMGh2IgNECOq19rVgLuJ6lAIXKeMFqrepPd
A/RTm4kUB8pYH1yFYfvbxjdTg7p0BDSeeEOQhF/d/jhTPWo1ml3yL/u3ocFfCizX
iP/9Tfa3J6FqjnuFNIal09xcNyeWIUlKgE8nHOQQR89G5kvHRawzKEFwjT/pQ/s9
/FH+z1om0Q6gmel7V7PxhoP/hwodLozGFxTuff/JYYTq2fgY0KMP+hWVziDvdYOe
S4UndzX3yBouhMYtcGfn3GJ3lCv7WCsYxrej7ST+Ezv51fUU3VndH4x1KHkegqNa
bhjN7SFbcoQ0K89Qy54mdoLli4UjzdqrjyGQt+9ephPdOHE1BGVr+usgcngyRA/B
8zh1m8fjLBfRUYZUiQ+b+/tHn7R7wEeVqkHhQdZXxzDsK3ZGz+yJVpDebYI7mcek
EBZP78aBd08jxoQ2LMlKnxhrIsS4Avq466eLpuV2Q5lTXYSIOZm2SjEB04p13BH2
pl84FQkaPCG9pV0hGGRHe8y5eGNNZx7ftQ7kq33sgvdKr7K/NnScbyHP5REil5M+
9qon/k/tX3eGDQ1b7WUtTYBZNw5XoChHJDv+APvv/E38gVjrWDhG9BfrzUO2jnLb
tJnsWfJyicWrjgkms2DmMR9v7Bs3FRiSund6TnPQANiKyQaBtlU1O54GMsj772fo
oweGoQOs6rpt2t8ihuXbTqGBWd4s9h2lslUzxblDgSMTA3xXa9tQu39CbihhvZ4y
T9ECAeRBwHeaiWEDdWP647Iufy/FllnA7RcxAK6KlI7H06Q9WapUSwIOEIl7YZHi
/bJig6qWTYp+JKV/nIY114DT4qAqr/mOyzoh7NazRZvBzvEQMlAChp07JFfniCCp
IN4hhpKmY1YfXqR2ONRMkfKUIYy09GNqGYijnEJioDJJPHKMvOAu+TkavEC7on6S
WTORxmvNodUguFnoAkS3/qRr2VK/z/CTwJ/ysr47lrLunEE4Ttzg51Iip/u7KHvr
lfPkkTDsx3eMJvDUv8PMdBsmIKeMbRYpaOABbLQ75VPYlA3qZzDf0FuaexMrwPs9
TibGS8dGV8L3sfy/L59vjFgIi+lPdRegJCCge/qlsxF3cVpECAVRLok8q8tDGZXk
05IFf06FPs6FgA9Las7X50zRYF7tuqJQRIrTWFuDvC3iOFnaGs8Q15zF9xg/WXJx
XDuqZ1AskXtHlvkgyGSukJCiTtBHe1S9vfQ0S8I61qL7QCLprvhZVlxei2GQEdp5
oXu5Eec05BQNLvjxiylSr6gf6Fw0HVPLhWe2mE+g6XydtLAwwjEAo6KI55KIv6m2
aS2g+I0HYizQzEpIBoXOEXzC8XchJ6uC8iH8hoGrC+duB7DupfuKN1+HAbOQeitW
rmL2T5hXukOr9wjyDX9ONsytCNDYx6wW+l1nB9jDq1nh4JQIkyc4NJbFkgTNqRAk
2Z0McZtVAMRrCxRNl0To3PNbtrNI6W1qam78NZRFxEih1v97Y9LoIejjqu6D6Ptz
h8yusSAAd8y1h/GmAt7sgckZygW9IGK8/SX12MZvofKi2v30hDTwBpvIfh20uiF7
+aW1F4m+JvzB78V6pjQ0ekYAf2y8ejfCHEn+crchMbu8D+zNk1LGPy1RZeJiuY8F
OV4MireNLAe16IAJmQgi9kLhKFVOAHUe2N38/6wtYyrIrtChb+sXy1BiFL+lvVSg
+uu3NHmGSC+fDfSohmFXUdBkutTHsBnUQsFCaordqIr5E0uxvEdQVGlQtWl7B0pY
ZCuzUq3oQ2EqPIpYFkussEanjlja+lkQDkhtkaLlSSHTyVwJQ919WOTj7QFck4LR
RyCRli5Z4+l3b/k9bCFeFOvNmDYP/2YAr69n5R/sr1BDEDfsOLs1NOVSxthq+9qg
gteTjsU7iUO9p5w0wZB+A0S/JLd5FGif+9ihNhBx5DmGwIuhcD6iO7VgND4R5wmj
v39aaokRGiYn4R/57VEP2OSniyzyL1OM5GdOOMhvX5R0DrRDpOf9VGXHxzoOhm53
ApmdHhX1AWBBMRbFpmdmfB431Ktxh+BQoNZiAB99QtjOMXBXZqSaMWFKg06O/p5A
c5RUxeFSxNZALuVAvPfNsFICDz8BxgGtFYfo/6f41dZV9Ijwpdo7bfqXuRP4k6ao
3PxOxAPrpBdu/2DlamM7ZQ7J36R30Hu6ig2uyur67oVesckPjfvSnt5eo7/lv9G8
vU5tK8Xsr+YxqDkrX+NSiN+Z+Rb/mf3VllqQJ0Oo9om5Uqt+iHzY3IjC6YD1jM0W
jDbp6niQFu91wEchgp4qHoXmcX+QRG5snZKpESSxf+rpkULkFoNGm1YQuTZ2CwCP
GF4qstosAwp7I9DnaPUc3J/6oo35ra5FO8gDmw84GM/WiAyeFLECOQ/1PStUHSvC
o1oSc3Wn5ejjy+mF6Z5oZn6HO0DC+FqqwoX7R7gMEA7LkL0BJLL8tOWdb3ZnBjI7
/dG/YM1tzbO485RX8kMscqpMCJLmDlxSyEihi8tT+n/O3500sDQIktjZUN06R9d4
cC1r4B1IQWIrHO07hEeh7MqSIs1Ja1jS1GOpNg/2w0crXXBdghfmsc1hkHnj3Hda
8o7HqRWPNZ0S/JcxwrOA3baUioBS14j7iPxEMkKourfksTaqu9MKZ4LUJYeRBAF7
HX2ER5aKPxUjUiBbef3goAu9cP+z+X4g4GSk98ib98IqyDuPQkp8muQKESyt4h5R
/6lHR574bc2W27ilCFS0mhqrYbG9FLlzECsCmcp2x8k8ckNmWBb2pRxoV40l77zr
y/ku96Cw3ogewJErr6Rr13rltPu5ukrzFfyUGhMTAB9RNdENfF/o98+97C0KDY2b
cXAS1YsGOLxKBSeDTEXeuYjeNiuzkYHFn7yuxsYj7tCufmB19TZWsu/aqsX+kvE4
DvGyDSXfpWAQJNGnsQVSbXJXcHKQDSb5dATzIzZCmi9/bWLzgtBj8jzR4xAzgs2L
fYQ56TpYBATp4U2mmUVR3gsAggq+B/fLRk/OWH1ftez/Dk0kn1TsjblG3qtCVJPu
Dt9wTQv4mjHJ+3BqPbodj+r+a1ySlRa9gPZxaXqUJSZzJAetBXfYoDi6NmirQILi
hejX7Kr1+53ID4yFCJFL4N1MkcD6vv58N7tIhM1VHvUlZsRlgPvblr3Bm3A9xybm
ZKZP1IKM56hdYEugJFXbeQf9GiuisN7Q1Ovy+snNOp/SgQ+Pb/4gdIP86Oq2vR6j
agBx/3UOov9cCsJGOxkLNI20qGLGgBOf8X/+IblKy0L73ivXgne190N+XD97hOm6
EcXtqXWub+ZztpUURddYhBcLmoVc/473d70wH6xz0UMpbtSXAkhr1euxnC52w261
xuaKzWAoXeuPK2bRGwvslsETTJ8fj63UhB1Ngm1oX5z6zUy/ekfccM66CU9ak2WP
GYT0h998Qnvctzvi9ZSkFF1ppwpgqQ6bratzaCQUXB661zyrxftoAClruLsUZYsn
J68RwgdgcBmtjNgSFqmy4XBcULCnehnLMt87+dnCyqVywg37/lKuEv+6rx38tBVj
BsvtuxbV6AlVoyYmjvpU977afJOVP5UFvoZm1YGdhIYAEb1QtD5sAIeSdx52IEOR
aTdDfG9ayZi5MO0W3ARe/DdcGAYmRag6lHwEPZPg8oD0DfNdjI1TQiMj4lFiZkcI
CcHYK+eA/Rlhk9cd8TnMoi2Ukx1xt0LszBnfm4/zAI60jcfu6aQ0I+NACr9eCQMs
zkOKzF5vD2RjowcQTTlF+mV8cz+bCNZJFQUG+Bmax6R5t/4ILY+xaiN7NvjDVORc
Zdvu6RAfAzUn0CN1Ley786RVBZxxgfG6HCVMLUNNFHJrE/Rprik2pAYWZbpsduf4
Exd8FqOf1Fd3jdHQ+foFAIWmxTNcNVg0unvRdKwb6r1FEs3Q/Kc6pjQ0fFa68O+j
qeHjLZloZG1fTLTO4LpCWdGCxxfZuE0iygHGbPLwWYIww8kqBLuRAlPD8fXPgt5Y
5q72RqrmuzwgnlWcl5JBcudNyrqneQvRKjxt2OtsZdkMD2Hl8/xhK6TrLp7cDAYs
M4Sg26FDfnrUtzlZjPCDzx3VcD5fTODxHAUDk3pcQvvhBQfrhW62jEPK+wwzTEwQ
9NuBQC0hsLOvK7a6GUpsRXPzkYfCKub0RGEb+tyG9LXzo8pnuzCbc06dVw+U/IHZ
JBg1gqH2q6nbuguRLNYNJPsRWab+9s+oSq8bjSr4JoYuw4hqf8R2BWhl4E+Uv4f+
Aq3743gRlzVWzcb+duvFtzxG3h5z/J8JZ/LaIUFS2nDRPMsfnjh7xKlGehGnfw6D
luw4dJNf/cl8+aQh1E+nsKwgAKg3nxzVpqyO5L3eWd2a3sKXauiieiPDHc3EIPdD
MkPHDEi+Am6meiEyc05AfwV/QUb2rDkQ9d01XixK2hb5wRe14ubAlxy0J3OtWpRi
Bc7L884/e1s7oAC+vAzy6ZBwQ35xKcXmacKKxvGTVDYad/TFqXZLrR4CkkjqrC6H
yZTFv27i4WawjBr0E8p5u6JK6hJdjvqrbOR/c4xsxnTB3Yi4tjPC2sVPgIz4jSZK
kpGGy71Xvhc2BTBTRlbT13O172S1Yskd3k8+TuJWRFar0DrBn52xJ6WJ8Asx/pch
iYVGzbaEmUPyhSb1vIUeL091d/mehX01IKU5wjhpWfXoc/shuWnKX856+XQNExBz
BZKcpQBV+ekQVpbUUven/SHXJvcUr8kMDJ9n9/T/7TbfQj5LBmzd0PZ+yqJ/aIJI
U3IPqcQs/acoTyL2/DwBCinSQq4XKhgds4FY/hJlMR5KBYVF2C5w1v3ru0W7WGem
Xy34FtZqASMvTBG+AtFNn2HuYGQjhgD31HzDpD3sr7ED4hpJj+DNm7BngejGogaw
VJXf+ZQHryTjQvE6QH6KSkwbXWbprg/AY6hX72m86uKvoPrY2KZqAYC+bW8geb7E
uTDU5MkVz0Xi2MZ0+5xyMdEqMaG6MaQuxJIhZR0oYYLJYfgIxJNGiOafEbRQVPco
Xc3jxOusK739A+qguRhYoUZWnU2jKrDZly0g2kOIOfxHV19H17Hr7Xsst8svJ16r
5J1DU//VOS73t6Xco6hfFMcCuDvUT8yTwjUQZHF4xQYyY2ZlxnTR33/Y5jqHaZls
BWOQAE4ppumxK2N2zyDpaEgbL0x4gzLIcuklqHAN16D52UzPlt1Ega/9yxBzNLDN
SHKhPburTHfQrp+2AhGWrcTnLJWCfcLd5i2F2ZeqZq0huBTwWRkplU2on1kh+Z4z
T620fDcpmK0sWopkNH/iJ0g4rpf+PUpnI3mQIXChrOwgFHKD4PO05dBHOC4hjYo8
yMAAoBm7clKnnb0sOusC041R3JI5c2ZlMD0/byLc6nVFEUYu0i2gMjLh8o4sIPCL
0nJSusc4zwu2oZoX00X1i2teq/OLNj3oO7CA9D2anW6GVG5BEIiMTmGfJvmora2X
63uglzkxpi0zLWIQAcBT0KKM0+OVMmo/4xHXlYkzGVzAjwGXH+LLfJDsswT5PojV
vQTpH6WvodbZ39GpPB7Uf83Bc5dYB9ARTaW3Ep3aRYDEIZ31/wMa55lR9sc+asR6
FsauYeHxqP9iB6UadqDuQcRzv4Tbz3PpRTkok9zFcumXeFecTutmScaGXmCRdoNM
YCa83QLFRiZemlvwW8YWnSWxl1yosZkvzB1/8ftdGJfByf0PsehsLT89gDntc4CU
iEv+GDpJTiQi9TX5REcHvXnbZ8MZg9Y9mhKKGzWSV8pDg+DgleDPjbS1CbwZoMfO
VYaoLw1X6RH9d102zv974BwxzPxP4pY+HucKWLjz1Hg6l16YHbwRGY+A0xpsTtQC
AoW1B67ziohr4T1RBQL1gBBQObYxnWxHjIF3Lc9/HqV3OLzq5Q4ulVHDowME4yhI
baoeuJ3EBtTo9iZzY1TpPXKoUlKdHMMTd2J12WHsD9cge2J/gRzwir8xnsW8cCb7
Cohk1k2UrKvICsgCSHcjtTxFmwBEfjqSisnfZ31hBLS5cBx505MlZd3Hp5ZKwVxH
GDCgHsUHePTzgVKBCOfDkLy2/T/vA5OUQmpV1AvJ0qnm28LmmIZSVYpva0Uox5GJ
pL/pfpNFOvjseGq79gd233MEqxwnZIfNpsH0La5uO30nUHvzsuQUbCKMkeI558Jh
tgF0sbXPXWPvAGGelBidNq+IDlLfnF+TgFKA+J/Ifenchl0OMcWPEyLPHKPqhydf
/HCD31UP18YQB9IafPffJ4VZ4MLVOqnJJr+DwKvyKMArO4QqDEfrxO9SaCWAmaPz
nY2ZsTyk1EzlMFkivOPzc1m55j3SWAXUSGWT2hy3xyitWp4B77uCAsLNFeeHFiDm
4y4367WfDbemDj+w5eRXk0alx2vIuSA4+861wSR2ZGVq386JXEQcoz2KLdFJsCO8
xgsYMndB2YUo6iQUchmFNQNiZs/bcpw1b7kVAhR8Yi7WNWfZ7XKP5pj8DvyD5kMP
NkADRGELZrq1y0L+exPQ/L/A+VlKsLWCA7ZQWiF3IJQv6cp8NaYOJ6Wn+AfsdMbS
0mmdAc1b+E3JwKxjkTdeQNJaaibBag1Q5+O4hjl7wkgEkHhPwJGdbWRQuWaDBOf5
Csn2fR5JxcaB+p+J5QL6yXa733RrORdX9L+wTQ3bjZJgH225zYd/qvgEUnhcV86P
90z+/CcfPRdhE8h+l8dCz0WSUOBmSkiXXym1s+2FljeD6CWYySnNwpExMuZqlQWn
4NjXTJ1DvVKYUeIL7GIRgHifZuJRHu3mRyMQX8hFOMc6OQcPBEQjiSBQFtRflriT
qjFaLwUFrm6hhwfH8xFFOa/5BJnNdnJ5eKb2AXSf/XWj1ICHn1JlCJpKaZTBZDcv
W6C5K47K8ZfhLksYXFRVHIJEUe7zBYyOnQBR+D7kgCOxDNYF+qeZQDhBR+0/tARS
UxFYeR9cWQ2K4SSpv0dy8OG44OKj+NpvCa8NIezZeiz7BDMXlO623xNKtU03HHEX
9aEjf9ooRBf6UO8ATQPuRFkC1aw6dHypi0WDXAhGEuhEyOXKEQFR54wtrgOWpDbj
lXPVcE7xHfyK6DTmImy1lXkXDOkGvn0YSBhcwsBy6ClsaaGGBRlSVUJMLN4PGO5w
x0HDkG6FbrBnEybe0I7EziTLYNYrggTh+RusmhvdJGNX8KhZ78euUafKuK1ka9zv
UK67P73pmcPuknR7fGeGMbwhJezyYxklM/UWqkSmsR+xcjE3T41ZjYMydS035dWc
+B88JHgXRqOmpOo0MAPo6/4YXwqEfAn4wXPFJxperqXJQNTRFTY++AYpkiRqdQgg
NISrF/phZOLtMQq+5Gyj+IIA3lKT/lK9nBmnIBK0Uk/yG2vT+mVEReG+yfVT3ORK
wUJRx1u5xwdnGhIbyQa+BcV05hhw0pljKP8XJ4HiPdIQic0BAyV1exO3PsgAVyrX
Q40Pc+s2EsZXSHkaW89qOmY58zhRyqt/tPOwud0MfCvd73VSkrI+HDtsLARGYx+Q
/O3oljw50EjkAxdGW+qxZrSDiArLFewkafsOrCW+b34/pI8Ym84B3qfGZK6G1HD1
avyZa1ATTGIehIzz0w+DFMKJAAZifkTlwkknAb0PDbjrgDoTBgYeFeT9ymaP0SyF
SJSG9o4XM9Az2FTiq21UMOUt2VLBbqTePKE6PU4yKD8HUOgJeZlNBzJQPSErgLLj
Cp/J22yveYuQrMfznAxPv8G6sPzNagE+XlSOs4GTRKk6PCxthnQvT5INeUNsuQGV
FTsbGeSW3jI/NnZKdQGgXonSKzk9qXxNdIfUKqtxZ8v+wBjaeLzoRv5z6FE5cf9Y
EQhrr5XwN1T8Crgmi7nMzE6z4ztg7wEY31yyJC/PMLM/Mc2KTplvzVFab56fmFWh
m9HGXvPQ7pD7Zk7/pjW5EY7WIt19XJWmUflgXUgEuOrjk3UVWLf7/Qg1H+4W0lX0
WbJwGxfsiDcFQIF3PGLkJhZbokxmnvAgUxuhvMHzQqcy67YPOvxEPtdVYFWpl5YP
T/n6rwGrDuitCo+scN7Ojd4dlDMwhBqWJ0V0bzUklahuu3UYuli3IoqhWG4orqhe
m6QHFrECzwysX5n3iJKS/jH7Jo+0UNSFaG924dtpaz/H6MmtWk9y69K0V7hqbKCx
R5KQK9maProDKsjH4Y8T5gwNkX2ECe+9rzWZnwwQOQumZowWVG5+Re7VaG9IU02e
GCVycZCgvYfbU1fGpDgHw8VVvPda+kWCyTIZRDvdIhYcoi2dKSx6xRywxuIm0Vus
bNphpRq/MHekR60fJbHqrFW7y1lJGxzpFgLBilH88Kbh34/BldhP9UK/04Jmfsqa
sRigkl3vEorogEm/IX7y1VucT8pgZdUX3LPrybZhlNQFoJjwY0qUj2d3mBZzqbbU
oVwTlMlNVokUnSbnGyyfgyQ+VckqaweWZox6ETtxfVgw81LEQmL4SIs4Lhdb+Yua
eKnEG07/JssJABMeZF0Bv61si+/MRqaQIuTNi9FglCWL+wOAYv87w/0pWidqsfnT
BZNHac0ehFvqXxs9lsOqqWj/Z2xRvVe3e4yiNh0a6UdcnfSbW3dQbH/TJ4mhjwFJ
QS/P/q5cMitZimJ8xyOZhSmGlRoiNpn+iZ87zyShNxijuadFaiSBVAA7WeJw7r9L
5v05MXz2KydusAi84iTr6CQTh3ANPHG4eRnw+4MduqRqVoZ1QswC33VR+NpiyHYB
1cLwJUaYu5Y1LWkCtjkT1EFRiLZcVgThHsZscXlwrgf791mt9bfWlVkpPRyEXRmN
KpMRYSip+F02FocmomFWPEFVIcta06U9Q2hwY9KfoMipmVKIV7YGy/XunH/cqmz+
d1n+A0CfJfWWwsFc6EwTeWiS1Sw5Pv60CB7YTsAngqsU1iKZCkvj6XsbxDk6TFPW
glnKgj9vEZij8L6ZOo4JgZt55bbnEnA9Up080gKlj9kZEHe4GmMYh9r/AopWyEnB
0ru3OIAvNWWrlW2HV8QwaLSVppXRsmub9waLDo7BfjCYChNP74iHkqZoJK+VKubI
B4s1Zo48NE0DZmqDR/JAWrP7ATtCpwyE/RR6uU874Rbix2CN95K5mx1SemPKIPgo
/ubQxVXAq2zKUBq8ttKhtMO/r3EtP6UG53po7hc/orJI4yI224nQp6HPo4sQ/Ntp
IcXKDwzi5SXne/E7N62JbB9OoB9MnlylMb8i4yVPq/Vex2xqlAYz5hIoB7oO9AT7
TRHNisEkimJ98PeriNbObPMQeHnI7Eb98ppMtWwoY3icJJ8Aw7fCGZC6ph1kB0Z9
EF3dTFS5GE5swBoDcT6iTBamLd7zUwWPcv6D4Zx7mCtTtBhFu9q8Y3D7hSIxcliq
Ws70SRCzgbGiMb+nm5U4AruDVDDtZCxHccxm74PIjw0/5st6hHJhXLS/hwpro2zE
5yeNVkDYklfcF1PXosSQe8T23zDcXwUQ5W55gB0WjU8nPh995qHgdL9HtUQlztCh
TLjJ2iaQv/uTLguSk7cx9m+atwLUDNu1VHqF6/AnKCYL4A6cAhwaXnFXMEwTm9Ci
PEoQKTzGX8LHurcIHhLszSuc7qccCC1tbR6KDAFhFbKK5awLhHEhXHIahvFr0uPh
L7JXfY5chhhV0va1PU+KAID24Eq/hUVqz7zd+wyqCa1UEetUKD/jguALJc0L+6Kb
h2aYuARXuZSvYoj8NZtj0GdIpC8d//zumpyVCoVbINJ+JcpW6ztYL9oTjiZX5F/Y
DYCL2Xo5pwBVEEdDdtwJYMcv/JaaVoTUWhgqN2KXDKn+V1qrPlJ99KWvJyGbs7W4
hLGywwLavmy9u19AYYFTf0rS/+8bv9ML+S68qSUaeeZNmAHQgqiBaZWvYE1E/QVX
8Qti/wrAPSe9yKBMQM9/bN/wGnE6R1xEXuJ8CZ1nYpwIsiDqn4TRI03jHf88vahO
Ic+KOkxxFTFu6aW5BYSmznTEw9p3gY22OixGkWpZhokXGO9JtwgvAAGjO8r7Fk14
X0w3qR3wwbvKFVgWAw6tf6oAGLCrnWvLDkOt/0sf3ji2tiKzQtbFPDjoEoUhSSqq
EHSD6+OLbSuDDTm1hxYiA9P28K8z8+YXI7iBnNd4btY/M/w/yXdl8jI6w8xBqJ4f
F6ax3XmZqrTwr3bkdWp1aFo4bReiGPLe0C/FYyqCvXu7omJVdNroMu5WIBa/La9b
txGxVPVe6/8Tlg9vaVoXZJIrye/POBnZY0TJpd8o+cx6UtcjnCh5TIXxfUkAGqw4
ypQb1DGpklLx2+5vu9k7H/8mjDDIR74JbGrOJGB0+BpZf97LnMbS0UB+SRoHt3GM
7AqI0GDcsGAvSAPQ6Wis5Pi7m5e1d9gPlCKWi+FQ0i0LLmhMwDNfIMtkhXURegXf
RttHx8v7Wnf53dn4dRdTieI04M/jT0GenOZUvF1lohJ1n1drDpf4zi5QRaW//9+O
DTT4VNl5Y9nX3mPCJofefU5+n2cIQb5bxMmpnCO5UOnp7NvAaLtIZSGRXQArtvEy
tG0n/6B4+fBxccOgZXenw8zNnGvJnnQaM0aujGN6C8JTMBvjQQKfVm4xprc3wvSl
bgcIkNpa+qeQJshyi8vGuArzMYBwOTaLpfptt/qgRmTkaxRqW2ctUP6cRMyJmHrV
T7DrW7B2jT6S21y1w23Y3YbJbrYp1oTA1M33wgeFJ4epvfw/ScdsmfgA2HfWtohZ
TC3IR/5HxkmB2SldK3LZ9UnTxTGEJJPQNwYC7gHWr3TeZ7lRgdon1Lar9GGMDPJs
ojgjcHcpOBlOd0HHOtSIT38fuedJryMIAz+UHTkHV3YMFJh3caPdll7AE1h6/+je
jhBqKnmuQ93RTloYjbUbnk9EYwS9X3uPv0LDeymQX0TpVKzaSU4BIL6i57hGN4hz
28inyfu2nbjlL7DbhqFwSpRFngLMQVDiaUL0XlV/HnPP/koS6WTXvQrxUjuouy4m
Mc5Nxsd1BRhdJ5jtq8xlx9x1uud3/QAMrGh5SBN9UJh2jtsOFEBp6hZ5PTMBvJ3U
VSuUmAw/SRBzrRIQBQc9dlBsaiSMKTdeLTZ71Q0MMwcrIUeQd1LJ/GvipjJfu+gB
dAyDrrC9c2ZSaAD/vJFA4IxRZE1Pg8lNrwLUndbpEWT+1NUl6PThCTn8BXLxn4pc
KzoA6Xh+xv3Exof957+TL48Thr0Niq6hT+lm8qgVGh3kT2JJQDg/gEjqkeOype4L
sPiPsy45jDP9+6snY9ahML3XDlejL9drgvqtBNJLXlhgJFJ3rpsOgLry7NMtp1uV
REPnGKxHWfbK256tyaK17T8E6UQmpiF1MlqOVAZtzDJHkd/mWJeuC/7Pj+dchx8c
fAQAFpxDa1gpQX4m0PTyhcyV4A287EaGqlmKIDg8/bN9cLeqJMTNyrzZPJVgFEBI
cMUQ63gquPDhGaJWAIdMMljMqVqi06hRGYjQvGR1Zv+85dSjryKcs5lgJjSqODEE
tzEsRvqiaU+TOWnxYYAERbltCkQfJigSH2U6bKhX8GWZf2LVDZvfcnAh72ZW7YRu
ZQtZDg3fmVMGf2XEj6KIdNG76N/aBWlwRDDIOOnlw53MfWsGp0xjA20H92iDLcBx
eHiQsS4x/iUV27GzF69mwk/qU2teXOXPSSEu586FiwXjic8Duvu1ajHGfcqHjO08
4ZCezLcgZ/0Pj7lyIjik9qniHMfBDNykpuNU49SESrrUt97+W8IndWQYDIiLuRrf
PihaAnoY7tYBMJGSpSocHbplTrbkSfdJ/+7InqM6/b5DaC0lE02t5n/xKE2IYd0k
0BFgByWQnTORTMD3rJKmjy9k4kszxn1/mnvQwzXPi5bBwRb0KYDxC/na9U26hRfz
f8ZR8tWsP3Of3nUwFMh6ncaWTjWstSKr6tX+8e7WrZHO0ei8Hngt12DRpAnWEtX2
MR5tN1GSL0A33G/8BMRsUntml0faiVJ47y3P3kD3r0bAlnKbY6CIl5NpIbINdm+9
3qf5iwUEJ9T9zDSVd9nV22muLdTFWXq+baIFpiXUTbMzlL2NNwxHo2FD/1n9ROpU
3KT7DKfHrstcDlaaQ69Zob69iWFnhKyKAg7zFv/Pn4p+TcDX3K1Ly20mTqbEGD8i
dgab5kXVQ3vRUZMJtZirFxXakycN2rdAwcEbdMftMOzAqjJwjLpQSNRnfeFd/OsQ
q75+KQ1ngcA3efP7qGmqnWJuNGHKR3DEY+HDiDA5x2MTI8GfV7RA7pRppuszjfQB
uR6RMTwFWgUPoTlq5S+a+bBOVG8DcKu1pTWZWKOahDfbbdV9P78gkLD6A0ROzZBx
Wt45Kh7XRzMg5xTYftfyYK1fAa02cKqDN9M9/4EvogLcS3m/J3i1VTTbcTgA8O1J
qQfZIa+uniuG9rP2yCNcKtBadyIEJ4fT0kxAdRShYnMe+m9ucxPqE4s6R3RO4Mlx
YISArfGwBYAY06lPMDJQ0Ev4V5jaAg3B41g5Te9rAIVfnsISScUXXQNajVY57gzu
YKV56uHm+PFroxGFjEb0zyuBVzuGgg8ZVsAL5fRd8dldbpHT9s50CwCAj6Tf7F4z
2lEzWYjo0LZr/2TQv7XoI7odUIeN3hjpPsaT+T47nnDWUhpsJRYo1/5c4e6O5ICa
59JpBgZS+Xaamcu8OcJSbKW/9+15DBOi9XFEXlW4tF3ynlK9uFXT3n+ekdAB/ZAG
EuIKa1Dxiwtqlhth7o0048zL9272QXwNJSeNuL4e3o5Mna1e1pecIDDenBSh1eLK
5TV39yrADL5yk03jZ4HXeJiM5gnlUuxeXe8FnleMQn5DrQRfZOHdFenr0fiS54oZ
aC+7kweP9HpAtLu/FuHdmm6rT/LhihbSdmIQFFVo2+qkDK6sVpSC/5PHa2krp2kL
GKcgU+vU4d/nzMG522yooXkn8n+DL+hmlTalI/fYCxv3wgZ3aZkqzSkA5qbpQ5fk
SAmXU5/kV0i81hJMt4ei3r41CffcRpc6OF008lwJN04Wjq8N51D+TTPT3iEFcqh6
/q7JeNEa3/8L5d/0mA8svghKNYrGp9qvVpyAxlPp7ZBgdpDdeRpPBgDpWvYD6tx7
N7oZPPw3wxZnx1a7kCkZR5ncnaNZ/KM9pwdUrQJvhb9svh5XzrEwrGiEMSvEl79a
Q3AhSfm9p0DG5yr5ERpwPyHiI/SpI1bh1PAZKPZHLjfkVc3Dh4mr/9GjKVbOV1XG
dLS92H2SvmXni7i/0Sa+G2338ZlYbNK8RoNtUStVbwdoU6cV8W8GP8uSJZKlud2j
yWP7PFEomDWsExabLk34rN9oi9V+65oibyeyLswUW0/PZT/k58vEkZRxfGeKGpw1
VR0Rp0iDy/ogAhRIE4QXQqL7o38HwUo40DDjv3GaH/L7WlJfZBhCAVgl7wJYPuTX
lV1nckgDwoAQO2jtlMUq5YTg/W6+YrGLyYVcwtqY6EhBK43iEtviJtXQN6HtJdrH
SZ+NDn8VjgTJxlA2yNzh0jYNlo5Xhbuu/bI5QBGS/+kO507N6QoFDAleiyZJgDFe
3ev+T5tB7kNHmLmNTK8WYTcgHmBYdUYAUEeMaFLU9RDOd7edpwMStwKjPxatinjh
zaHnV1bJm/+owvYWbBvcu8BMAH1zvJ0Dutgfod/uInV4tPirqtP/TikdSZRJEGH2
tKAGEueTIWsAK6GGUVi3TNQ/6wQQu4VlCwJFvxoXNqpSfUbAIc/EkRLk666GcPMi
391+bg+gZCdQzgErpUvB/WzN5XOsy5o7wv9Rws7GNoEZxNf/HtlUCiG9qbcB9mJm
WvlHKST4+RBbuvnI371xxojeVEGU2nxKJ/VYGa/aAfY4kJeIslHxrJyirz9rHoOs
WJrVjMFkX9i/9Y2axXniW6SqAUEKaNbVAouQHP4i18aBPt3uawtHJaWr9iWDVCtM
OWsYSQDELGRmZBli9O5E6+KdvGnoX56cL9oujNjoyLwmywmQB1MOqST+jYdbqmAj
Ex80QyOjk+/PIYKG+85pKnsDiEgjMUCp72krCBziES/MOpTmHjNbLmS78NKQBjDa
Q0IH6iJBd5U/mKFNh+n376m1NODd7K2pzNnhghknzBHM9zgIWWYp1Focc51ZtRjG
/ZnGVv/6fDuJ1V+wmZKNRgO6s/9+jjW32oFe0tQ0j/vkr831Bt8NmQNCzzo7dlBW
lwRh1PQ9HiwaC+x20Ka5elx0TsIn2hqmure0hOOyfWPSvOEHd/p/30rDt41pXyhQ
BUXFAUvFMLsXCUHpSlUIQjl9XhqnKRgGn4MHT2/ba0zszjqBXHKBXVJza5fePObg
2ls4o0fBjWB0JezygXRjuGE+RJVeQAPGtninnFJ7QMy4MZ8RLhCvLMB1lUJsAnnz
3GbdJeSAy3h72TWk3gsV2uzoJ9v9xXbHJ9fp7TXbrLyuIGFWTrUcYk2Tlk6anv+y
pm+vYr5iDGInIxmNtxma6L/kfRiday1uY2z4l/j2wVE7PKtwkBzZfovIQIqb06PL
XfypRlwUhkb99jRsFeErBTxbfWhpZIe+BxKBPyS+z02ULDzSp0fXj/4DTjvwTnBu
Phxl3V1xG8lrAxKPaZafwAKABGXo9eISTdWgbG1MVdxAk6mOt8y9fy4yldGScS/0
dcmEnS01zP2VhjQU3/MC+8WvFFUh25aggo9fyP3Z8DuP3BD0p+TWNVUwgzEyccjt
AyCAxoLS2i3RstozwFZyFAQJ4xDJWDZO5zsrB0OmKMrVf+j6D/XixgW3/U6y1IEE
DNbJknBS3/8GgtXw5dYvnnSPJotdnmZhD9lCPtMKLV/xfz0WhGucvL3BP+/CSflj
1dRFCfnFcUGfKRRh9SkQ7VJljOdlgMouWAKGjvHFE1LR6O8j4tfk0g/8HNHOIU/9
1fhkei9RDxtNxFtdUnNhu6CrQfpX8dhSmJF8btqkbHK1SI7xjcXHMGMr/zsjZxgA
GKTUaettjgArhDPxdDvxdJhGP1GTgHsI/DJk/Vb7C6letbWmrN3fumDffUBiHirX
4EXlWTHjYDAquZsiAFRi5iZrTlQl/tyzZdlU12RMGu9GGSiNytVBZSI4TuwmIsUa
ukdGOdGZVzY92qE7LUGsvS177hSixGljVeTmx8ubsJohC7HpcdBot8xXqtj49i5c
BDwGrPMj5jGnU1c8wEWv9NGL2Y7WnNAHZy6RK+jlQbDxQKBCMDFi+GhgprDlJXSC
uW/9paESPTjSuJuzJrGRlPAURX1E/NJsACfk92zximzgaSnVNDAmm+WZ25BKIUpt
oNDNIPjKLk488g1aSpWZWCJMK2LA6j0fOJ62yrsrqmtv9Vdlin7r0J/zl3IAdRnb
j9N4MhpOjR+V5oX9HlglBfMH2A6mCrd34AA3p3CpA6neaeIl/jmgOpT6T+jvVDaz
hJdczX9TvnqPOrF1xB5/ERjNlqzJm0X2JCRTPtUqOlEmutOhATK5wWO1vmomLFb4
4JJY19AfLBf/Ks9lBdBMAxsDs8QOU50KMcMjFhup7Fycd2LJ8El/HUPW3E8ZXuqk
D2oM7BecwUGV/t4B5y363dKgEgYKeTdje0v4NMUsG9N43x7LzUx1Bbe54Gq53W7W
putHmIJwVG1nP2Ag00rNY1N3BVqgo+hkCWH/N6absKfjWRGB8xZtrso7DP1QaRCM
iOjrSlsGy+/ijShdpY51wo+VCBXfwIYLKb7+/tGNr3oEWcw2EwyteqLwmF4BWpj+
JyH6yZUDgp/seZ/jYjPekmKQIwxDWxyaX6H8jdkuUbicOzwtTOjr013FjPNAgQDm
u2jtKK9csdTZ6TSv8t50Pv2HsXubG/2Rp2KD4FRug1OJ3kXlRQIMZ86pY7v4qq6l
6FabTCxCAivPXHkQEA0FM7okKv9GceP0YUKjCA3Le3nhanW8RYz05WdHmr/2YooW
UcMga3V8+XyS1gfyInSekVcyPnemabuWsWV8tEorlQWat2D2sbTT1Mbvgjm86Z92
p+tEOMfQl7RNXi9eTjygnRf2/f9fjzpoSY+JR4DkIIWftXv594tE7PB0yXEvmYbX
vzpQ8gE4bJVjGLDqFSk2NBWYI77lSrepi0bBDQ5qNJ7Wxvt+38R7IOxxy22o17S8
CPMUJ/FfDLTKkrsupSmOBq0+IRaHzHkbH6gGMww+NITET5tuegJYadkwf4u/RDG9
kasvtvXdf+Uw/TCnl/jjBBxPCo+pE1flzuxtkAYwa/f0ONV948mSj0+bzWd10tjE
YLD4Sk02R7IdqMEIhf5rTapcRm5XZUu4xUjFB8MulLtpSMEgZKRsTsukRJZuXLRf
lsk0vmFrYsinkGHDZpmlQ41yTi4TeaDossLdX5qxtIL7fX4GdFE003fcsn4fGLbV
/Vdu3HZ8iR1Q1pc8LQEz+NC2ZSFbHy+odp6s7CnzfimGOxXmlfOphaRWBvfZ+9cN
N5qJUT5nramzD61F8pkwyXNZINfs0WaGzo7VU7sjbHSoARxEIWA0LrkIho+GMXBS
q34zH2BuPCE+wJyYUTvrthqzNElZ3p83exc5o9IWcmUzwTzLhrKntk0x8imTW9E0
BaqOyzLneCpUusKP3sMVeuK7aOX8d2+yz7y4vmQHdd0nb4rYgJ16HgGK5mnbah9X
2CVLrS2/Oz8oa1+hZI4bo5DRUd+2P/880ve8EMZKh2AXB1Z334s63qxeo0U86a8u
hNtdS6AgcQy6wjdObcSRJTcLpKfq7Hu2qMDh3dXEWh02zaaHGww5fYFsPaqhvv6n
1W5kM0qiyPAsOHt8CzMQP7qx3PQ+Qnu0iQjrlTro1G8k9yYyGStnHCmzsPYaQqiO
NZpWzYX3mlon8ymXVTfEOooACNymk++scpZGevarkP3KGYLYGX3UpjpJx2u5lvBo
Zp/Hx4Z3vkjQlSk0iF858qp3EBwruyA9Z+U/gPVprIlO/ujK3VZ3xV+0Zl7A/kSj
5Uujym2Glq/1GDGmZz08qc7g/XDw5y7PRRwVJM0IFGrJasaaJYPgkHHAtu/HQbdF
vp0XDz/u87HtFvBwSOWQaPwDv1uSFRGQew0LH7VjiWPX0nv7Ak9uEYWUZ9u/ycJB
slf1aGRfDt+l7YXtm0PSCb11GE9j9oeqzceDvptjR9J+J+f8MF0pz5dCsfaXZrW5
1UDejCabdp7ss69d4mK1uhpdpwQe3InxFXGsqVVmwuySRm+NLMUbw+GGhvCAdqYD
9SaTUvzRDWs0FVXl5uVOWNihIq1wnkPhkJRzt53icsEVtMOnMrN1EnRBka3acPl9
eVG5nSL0wziUJ5yOG7a0gdrN3FuKWdlW34B8p7ER9dj0ydfOx8DtY1o7GJpqxOPJ
r3qtSoQovLcK67I5bApIPo7oEdQh8PrzqBNCv2DIK3u/fB4ZuhwP6XmSQHxbWgoy
b7OVe8vN27WjOs7Z7ikOwQKAFRJRyTxHfH62vZ+I/l7FDSMRjorqiXm0TR5s4Dvb
ELoURk4Wpj7gqo4DSjcgpOz7RndvMhiPrm9vODTNMKDrJpq0We+pjcX+ZGXdPywo
gCVzvvOHdy2WvVX3d0RszVm3Hg0nty56whF/KBzKr9CP4cMLZABZSATzQjOGhfKL
QAfgTU+hUkDtU5T+zLd6VgjYJOqzooMxtPlL8FNwiEUW9dzhcovKjLpcLCxklcop
8GmLyk8dbec3ZhiJISLUjoUlPgN6Rbji5AzS6zhyTtEqFajXY2Jpeh3zXM5x7Zvr
L5+h8qPA6LrfKK/WSGFXMrGxpq57T7UDTP1hBTlTs1NmxL0ajW7M+fIhgBjsutQc
mEGD3wDihHoYCKqMmmxK/0ghXDtkHENokLrmKq7lmR8OXJUnr8+btU6AT74aliH1
FjILMoUO8eInnc4suibZFj7tCiQ6y7PgNZHgBGzoJL1746sE3FxxVnx1ozro7Phm
dVfJAlM2keKF5kcF4RBzBZDpco+qdbIUo9kYu+afG7/KpQxsAkxVlwRuHnm6/Wf6
2gprd9GSnUk+3EtKFMv22XNM7EP5I99XkpAVqztnSt0ZHM58IN3JKrN9mfhzz6hr
+kcPHXp2g3iqaG8IiL23yyY9jnvdWKGZjYZAKXOxscgBB38zNiAWNRNxCEH5OEPj
LqSvuA7DQ4WjsqXcqAA+rb4xNQwPur3BxzHlDho/lkzD97Bd/sd+fbPtncc3TQYm
O+MfqP/6UXIsmPq5APP5AZRkDF9mDMUIAn7CiTE2mCzhdyb1kjTU1Q4cxaKrx5D3
uN711Z6MA4wOcxVu6aJyTRz/u63NQAlMp3P+8NqXjOb+Qqqce+qKg18BE5hU1nqs
9nVXFJ8oE3rA95YnE9cbUZH+gzvvFVwUTU8TGp+xTmJielcUFgBC8LFlVbkaX2BY
pFhEjOJuvECFMU9KcgEA8l8dLDQ57iM7Pua1BkiaAigMKsq1cNGKSOqgeBaH5SEK
JJedtOtR8EJgZ5mx7UVYtzbczM9jXkngroSpMVTJC0L8LbL2DZDjLyMCRE15jRND
4TDlpJB/wmgUwax/IOd0N9EBc7nNyyfGjFLIjKlILZj64pUmiXFdBcONKkize630
1StW6LR9NDvFKw5Gc7MOPLrBZLyjj7J4ghx9SQqDA8NUBDSbCVe5EIRysbuu4hHm
be/1LX1ehOoJVgyKYMaCxCZmGdo1j3Ay9sANpjvwVoEGTpEpjMLBJ1wo6XPWz6w7
82yT16lXBR1i2hThIeZOOpbjf9W6qYAxqGuTIvAqEo7vVInTvV7DqnMK1zVKnO2a
aOCyZTgcvdbs+Gw+p/VRR6Na5RnxMMp8W7fuwjycbT7GFjhzDstGH2wVe5H/i8z3
RmZOuOYNyI0QcaUvg9efED6jsxSOmHBn5zbGK5F5cDm9+xdg0x8wnv4eGQn53980
fqNwowcR0XnC/YTtOQK0XL5nXc/WPn3M2iOUATN1ssqD6eBWVYW9l4Vp0eltROpl
MZIeX6eRa0kn10p5nvk/QnFJ8QG5XYQh6B7ry3e3xP88XewHGfnVBK+ofD8Od7GA
A9wICLBlF+4MXQPa5SemtMgfTtJy5aRp4zZsf+J+ExVge0+0bYkrZ72C0Boka1hF
BWEKYQGpSKkyDS1Hv0woEsEkftCZ/o7tV3+Bwmz+4S+dKCmNx66o/sbIaAGXFaw6
iHD/J2IOsCuZdURe2RHHjrvAGgbnGSFpOio5v7iUrjP/0R1bQjGeVqCHUTWJvvWr
r2+qEH3ZpNcZlTzhFVM3lPjo0yX63b3vkocdmQrzZ/3uO2lNgTscUvZgbD8Slr/P
RPJ4T+PRSDUL4Y7VL9ZSgKIsf/rcvuCFOXK1aK1yhoNffyBlqus7SSercCWPeF+T
BDDsqcyOXnPaRqk0VJN9s7s35kSwa5yZxz50tHDH6YhMpjlPAz/IdwFmpRZP6387
B0M5BpyqSA3SO8Milt+o5fYPBjuxlMKgpThx+04wvQ5PJRRA03mnA0zxQzEenICF
P/91FwJxu4ASjJdqLWGAi0F3XmfL77VwwrSDjayuu7Zxvkl75/Yvrl0XsoswMmqU
J9uzjy09Sh8IZqncIp9tFmOxXth4cVi2v5Pag0WMGrKww8EDlBfFWnRSQLaUK6mM
7oZH+60WSioP05s58kv5qJYgVJBuEGKNF2L87p5qgkekMyDLTzpQ5IwwtNUjRE/M
16YNZVhuqwNwpd4uh95adfdow2S3yM/trP6kfyWBhgYzXl3BW6IYLmfaVja8xCK8
cKQSlaABeQlK7K+jv/6Igc7eB89UgWbfg1dXw5P/TXMo1RMqDLbW0PP+0BnzqeUp
qHhcnoa5lN7ReQ92teTCiECLsHI5spMXyrTEz47eQFecDI6w5giDvY8jymILdmz+
RmvIsJCW4gyqiJEBeB8qvwgvOrGhq6t855sD07XddwwSuTM0C2muWBN3+9zsZ/F/
3w+OStkcMNviS7OiTpq7aPq9f0vQtzSRK/WwqiyfsQ6Wtl/HuON2lbTIgXQ5PdCJ
nFRx2MJ4BxNlPCXAu6YDS4mgj8tbRq0Lu+1TPjayK+BX11oZ6J/ziFT6QS1FTlLH
ix3RFZrf5A6OGG/kO7O4hfT/D6NL4MqRXqRQAsQ7KEvGpMnu9xIO2eWEPDII75rF
xpoyWz5qkMR5i0k4uglxWjKOT+qlVCDVkjZIAV7Frr5+5P23YZNO+oHsIpfDjxPm
yJjv4awG97V2XrIjlmymJPwcnoF4foqY7QTgDnbM7JxFK97xeBJ1c0cuA47GNR75
TPWo9499/8DClw2n2DmoBrF6baKaINLkC5ICVZJEEXxi+aVeEubFX8Eg4Ht1bkrY
kcTtWWMSccrPB27JwdkXf3Lgg5QO+fCQ2Xus8lUMgkFA9gEv617TXMBr5aNv0xvu
ia9xJiozpST7VhdoZKN36mz1+39iVbfNbqUIlt57mJS79/0eWDgK2z92sftlVUQS
cBtdUjYVs/O3zMBTGiVpzu2BiW1zP0r1zrs9Hl9OfBUfN64wgWaQcoKB2j6tu3u9
kQNAI+BF7AmVu09dlJCu4WFaWVV0aAfj9dVGzC0yWH4lF7d22Q1ZhQ8Z3kbwhgoc
hS92R9LXN2MAzNZsrC32Jq+iai+HpUp5l+OMcrh9ZbzKNAjwpVG299yXfgv6+IA/
w9GlIlRoLbEaodPomcE4inCuvXvIiO01fxL04hwL7RwYS6F7Z9Smx6UkjihwRje2
Iklqpef8yAyzpfQgYGZFUkpq/F/ILqiloSeUfGrS5XpuNsEqJF/EXWYS0FtPsjni
gSg4k3mO0UPFKFrtNOa9S8t6L+lRFtQHOu1576q8KwQrsI2evBKzDVrL104JfM4B
N1LglZjehZwMBk4yrw/z0eYYV1icwzWtYyvRfKun5/Luo6F1qUUaOl7HzQO/KuR7
4S4GWLtk6tjcs5nixFeL7NB6Ft9bdXCRE2Olj8tcnyLfzzM+gtxwbiGsnb8beuYC
idSK94GGOShp2p9N2X6b+BJeTX6nNGw2sZQHKIG3jJ1YgvK2Q7HPRC8WB+p1kueH
IZyGZnNElhGpudtm6V3OmnJu0eRMU2cRx3hJLF345FfXUGnfCxqDckV/Zm81NhN1
jWzX8d55JLNMfCci1jyOj7Pyvnwb9NuqMr4ESc9xFHeRhJj2DOw2Z3eqUDCakFAH
Wwb+HimnaAzvR4JUVNcMuJE9B4Jny/egGTNe66koDCCB28fhyincZA6QtjXHlNZO
dfrJMuTydpueRg4XQQiYrRZXftlysMZxme1tbUzZLR7KHXjNz/6TCptAy4tUi/Yk
SWr45Hvf+1Mqc8CETOES6SpDs6We85ltKBJoIYuAdRtiyBfs3gog4ZJdzH8tQhD/
lH7YBm5l9uxDVMUSQsnTT83ILhJXRQYC6T/1Ph7HIuWTXrfj3GIRDznlZO/op7zx
fKN/ekLSpU8IdRKQZKYtsK+Yyz8umd9+mfmvGs529svLyyRtEU+4Pe4PmsZp1Nhy
rb5SjSgsFLGXeGedR6fhiN8GoUSMTzbHfJpte6Rn5RExp4Qco9JTgLa4XaDYxP97
CLO/stBSKI/G6xRtbbOdAHOWy50eEDEI+wFFkJPy9rgQcGGrsDHJJPoFiErVZyhj
LzniqcX9y9wP5vMX7eSXMcxcUl9Km6e51kSGAGA2U0KaH2y/Zvb8HA7creNxVVLM
YgbhU4lwNpO7XYW/Fwg7qXGQkBBw5SB/ek8Pts0vcGj/QbYj0/bNuq/0Q1oQIvit
oTSk1HKAb+xn7pAeGmfvxHTK3Tb6woAknCyR3lOuE2A5OVssU0Rm4x7Zmtm68kdy
gHOpSnHuGOTfFhwyc3nIOR5X2gXQIGmWFHvFiBlEMWSiLmBshFDXpJbkjIsVa5WT
P9nP2tu4u5jJ/PcZ0iIYGQIE8hhEW/PORkZZ9KsLTymV18Un5ZXOnoIoC+t71f+z
tNHb4yipqsHpaFgQMDdojnSieGJW8idMbNc+BkfRx/qFGO+I13GuxIhfDhM418p9
yaqHdCt643mUk7YxHvwr0wcMCPGrcmecqOtz1dIurMbBcA5glA6FXyDQvEZ/yG3y
1W6SRohGoRGvKn+L8zsj8PDDMkQd0fa6kFCRtyk0LYFltHDjDUmYMQcwWSZoTDtj
PQpnCMKFjvC/khV+Fw2ZwR3f0pAfHIcRQVaeSJ+Me4QKMkC524zgdBa/ZFFWHANi
EKaf/I+WZji3mj6Ww65K4y4js7e4pMWyS/IGFMFngnTL6wOBzaQ8OxWohOVJW60e
YYClAcQDX+Ht/FlmOVf2IKRz8hGO+FXW8bsstBlpeoVF6opkSm9fTxI9IqCIaDik
u70T5mD67X6AguTgpXxYhBxgSRiHiVh6ueLNbQlPc3hieM+9jkpeP2Mi+3JClNRR
8h+br+A7ZyTXd6uVM93J6wzvMXuWvrXj3om1tHpaDO0KOeb3WDu94eZoJwjUAsdn
d/YE3AmzFZ8TTPuepl73LqsWI9MPVyDoLoeys8jo4Byqx7YhpoWMX4UtHu88KJOO
zuppOe5Wyn4deyKSTcCSPEjP/BP3H3ymHq8SQK9e2syePAM7eC+fkx+csGB3NUpy
03drD5LtG7V73od1AVD5a1vE04XvtUPFrBO/9iRN+JCU46yjROGoB+3xry6VDC8a
FFas5gWTK+Hi4vRXMSTuMrE0YZeIEbSiqaohpdDuv0UyKXKQq9DcXHnVLgMbyrML
7qMIbebMVJSH1G3zBQgTXEWJnOSrxgsmW/88vLHoBaIlgJCcnSLQkTHionCTt44G
/E9XXF1F4rAlTtFtVR9iY+v43zcJnIsiwLn6hEFC7RQXXf/jihT4XJori3jLBXJZ
SASMPnBa9jgaRdtIwZTzJTsFfmYEC429jHGsAm/YIlNUFjiP6+SJUa9Z3EZpnQwK
JIsEQWyWZ/rbqHoTtU/S1mQRIQ0OGnVnNLmVLPejTjDTH//ocYaxCTK8e/QFtdV1
v1NpV36LnsutVJhz8ItrJ56V/mOuNuKN5Peo1kGfICtmoOCXFV/92EZjyObUFsSf
05NlrHFd0399oAq7oJRJqJonGPqeEf4kXAdsLCSIegc3ZxYOMMCeYB3QplDUs2SJ
UJzn+f26IoPS4HhShXLcbGz9/qYv6cO69ahaijrZIYonfNGUfegWDQ+ClL+JXU+D
mP+CAePtlRaNFdAw4QJKsBm7YIr63NunT2hpACSvh+/liD62ZdbUj6CJcM+Bu2wP
MRI3544/iGCpNo7YKzy8hnKC+no7lgwa8s28RMUcLvvWQXgQ5d1REiu4J+PrCo/q
ElbdjSXHL03vPIdiPmT+lsNWDsKK6NU8XgUsGuJt5yWZItoBl/uiheMK/H5vG/cv
WdvOnVK6Z2FKiZomYh7sMKSyVKf9VAGyqNzSy2kfLz5bFrD4C3nKqu9RnNY3h73L
G2qcxF7QAO0xMLTLZ/tp9Cs31EKYQnkkWy+fQTEW1Cn4GiPk8uP1Ge1FkD72YRhO
NwPX9qxUa6VNY38wmrW0O/sc6HtN9NyPB15iO8FXFx12hv3g4zZM8l5Bmmq80guD
vcnrzrl94gjj8kPf8MLEuGiu+z7f2Kxl5bZdq1rNwS7dVjRsSuANXFiGEjOSpmV1
08cg66K6urVJ/kxl2N/Rbe1LDEm3+or7B+uGoa++XpjlHyCnZkUoDGzqU4jPDRKU
c/Gk1B5mPZELPZeDZfIAhe+lq2P+ZsJ/S+lVUWhu8WK0+2QoYJMt9t+K06G9tEmg
ucSEUQYQvISqlwd4CFGMrvZUjs9jzOPIgFHd5nrFJQGv/11zwNO73H3yp1Ws72mt
ioTxge5hT5BIcynMFRiRURlky2zN007N87/IUhrw7l8E9HWB4HIbzIucl6SdYWnh
mRASsJ2iMCHShlrIndGs+NBFLhzb+lcvwyZAgx5TMScnEHI8XNfWtRP79ujQfxnI
GdyczcVDQ4wbgj55MAVxWY5ZYClCTaV29czfEB3VOku51kTKuD97BMdzLRGA0HrI
oatiYV0o3TpzRLea6xIdo45BhRoPZbQhN+oW8+pMPkniVY3xh/hE56hzT7VnxSAv
e2JCWjd91LbMKhMwG+6MGJbgYsVWHN+7VeSXJ8IfXypidg9uNjNXq/fLmyaIc7ya
M1JXen/BAT/unoNrw48x4EJW1EPEgpZ0zYa+xH66OgW5hTPmmZot5OOYqnlIiLlf
eabYh0xiasiEE0cPHl2BqREjdJS4vcopyBWKtQ6OmXevfr9p5CN67wxoNj9bCa8a
gAWLOJTShJY1pIsX6WjmBO61fAxi2rflqSZgAVJJesXvkbOa35Difs18xj8b9Afw
9zvKpgniNWlTCnWze4SOQIgPR1GvvLwbzPJZ0Cbe1um8RJvUsPxO5lJWwCw2W/x6
syPgsP0gP+LHKaTNG/tjQmbvqlaNbkKtYlA3ZN/3G0SNellr+yorM5pZ9vHHPShj
koJSmnjxV8K63QxgXL63EL80YAF+1EQpSnMZF0PGuTIe37ntnuuEimRi4sg5dGrE
O4gD/X8Imnpfg3Njz183jimXdXQq/IijgX9OPO2iQI/j90ZL4J7ZACrannBHySW/
TBqCkl9yBM4r/k5SSQJ0bV3RB00QBH3jOXA6MrKJI9p3obcP3XoUxRjWp0HpdUaW
wac1TEPc1xDoVZhpLlOjUL6Ioo6AtMvP8GJZyMCpfJNtuIHlNHLjFhjTthjw5D0z
jGuz+NNFlLQLKM1cyao7rQk/+fjjUdccRQhSBAz7ZtYx5oSkTPY8XcgDVYejZnxi
78BI51Aux3rk6iA/CY+Lefh5+J4sF6aWyzfbJeTFPh8WA1tZcYvpGf5s+ktrBlZ2
ghuLFHNRDbuuNnq9XXWzeiukytTMEU5zq/7XXrpIEA4+hga6OhakbBo7RbsPWe/F
wYDD/LnJaYCXAnQXQxj2Olq2Qiu0/caB4kNJw/nCpnO5nRKUEE8HShnHEBw/+5g3
6cGV2NOFUr3M1dMn0LIvyiAIqbNn9RV3eb7FB3zeKCTt1vX2SJyhoAo2HUELQtMo
CggKF82bykL9Ye267JEBwnsTOrO5JL6EXN8D/1lDqDR+vCkmO+tLp1WbICkOYryd
E0Am0WGJYGNezYuY3hsYp2QTD8j9X1cFrHH7v+WkdZ5oYSEMnXSvhoNi+Z0G95PA
hdQW6aq4ImxzWSO1UwHCksuX3PeZFzcBkzqsG4jTJy7Vi6gLW050iwZ6q+fStNCu
5yWJMK4hLIpO4i+hToIv2LUN9dhv10e7FkkGNtKUJ3CwyOyvQucs2/4M1Xu1Gs1y
tIyFvjIsO06mFU+b82/7xW6d9pAuLyxOk537A7/7t3JRI6YS2DvzXTKTaQoUUg1v
flIUPhnnsdfg8m36Q3yYOH4PEHv4QWlsPtYnMX/s0h+lJPvDFX/ImT5+1JwFNYqV
lptFg8el+7Lm3aIUiC0JuYCZpCZzVCe5PEV6GqxXrcxrBNwgoWivjdRPvb79jOwz
5EHPlO3lWO+3l/y3+Kn7lAVDDq2/hACTc5PXERxPpD592fLINokYns7bBF2QTxqx
5hftnijnDNCXVFuH+Pb10XfeyInNVzG5iFeSWgwn7mSfs6G+h27MHdSv+cVbcFuJ
CVHQiTF0cvbqkqq/XvARtg8I6YRUiSnWk7VUnY7pW8b+H4CTkSIHwiBS/xioOM4o
1+t9OnfSVqB84z/nICRcz84TJffhzIJiKZmAGeasjp2DEe0Cwm/X0EpQHqCh0Dgs
Wv/mbcHTrWmRFBTFNKw1caL4g45v0immYrHJSP8Nl8ET9BuQWAM0J2lZHV10at5J
ezPOGO1aKTfSLQHix0T3o4zoYMBTGsgLRZQvSxU8/jlGBaMkJ6vz9bhc34FLDPoQ
/7VUsf9uOfeF0e0IVP9PH2y9UQ5a3s+LiGCOlpWtkY4yQbgRPZQ3lVDAWPacZLln
00uDwS4x74Q/T9dMg4tghSrBUz9NteJatYusmQmHvAZcb6+dqjVrbliLL2sJ0Bml
Agdk7LZBbfgofe2ukxuXCo18noAg6SU22YFSS6ZtOJkpYb9GbAk1BMRefeBtssYI
9OUD3T3bP+RJsBR7U2GO2mLtPzUpG2pbkw86DkbeXGMnBqUYJWOaKK7bz5KHEr2U
NXvQd8HvwvcRAQJgyspt/JYyDT+Z/yjUKqdUKN8mwjd62oZ0DA1uLXzF9FcDeff6
JL4lBRo5vDWO0TCMtHqGLeGItpepdmNSOu1nLxSr9D/kg/4t5Co9ILjkbWFfMCU4
iDEcq29LW3GVu8k000WqxtpfRen2y4CoPozZZ2d5bm7sc0mVt8uvldvFkLJS9O89
STJ/n/NX8GyNjOLFe6XSBa15cs60UPIYpaEztgL7GLJQlD25DYwcMIKzpULuKsTh
5fm4ZDOkUFAwybFvRMxhCmS3l3o+/PuWXnYNGVG1YOPrXKPW0soS9TUYrie+KbRK
73aKOY8E10vtvP2mCYpYYkyC/jx39QEgcsm64lR26i6p9/cc7QXZm0bqrozh/W8y
Qm7bboGnOnCKfGNIOgV+vNgrG4h6kM1m2TJmeTH2IXt6K/15IqLhm1LvDlQbU50y
oDvBcaqHQ/BWXI7FoE6JlpA9yiVAKEu7NcDuJ83jfhWvPYoryVH8U7hulfb7gFSJ
qRxCMHzfbJb+KPBY4vCY7s7kRg/c5cbpWw9cJHAFlDgvAXdVTPBDyzRgQiAxJELO
pVMteTv3EdHLrYmGZ+kun7dMkxtdJRxkEnyQRkenF0oHdez94mSDQmY+t8VvX29v
3ZHeYjVhlnQFpKrpmctvkCOYD0NQsPyYBwTkN7orWVA/kj3Utu2xlOIpckXcndLn
0kejs+kHAIMlImxs1eeCRdIulrqpRs6a8FyXI9Is/WSYHd8eIXTvRjImGh4hKlMd
8AzynvHB2f0KM0EoQXiuwoAIAS94+ibkw2kNbSKT5INXDjpxTErhMaKrWcqIB/Cj
DvHPckZDT1MGJjYLGgyVbBFaIuwtlNBnqF16xd8cR+6qR+F71oCNn1/EzL7/lc+X
WERN1QfuVKgvPGjo6S3iAzMlBV2bGuhsAcjem/wPIbynAoA0CnD4xb9pTt2WbScD
zaHaBWBrOawrmgdbP2vRV2RHGwJ4pOMp2/p/9VbyfcD1HyzQpFTZmaHBA1zorTgp
yN38hZcXFO7ZttNFgr+uCu3uojjR27UbwbE4ZXkiN4kQCPM/7luC0yUOanoN1Fhd
DsXyGRf7t08UcNv9GPCi9vwIP8LQaBIc+L2u28rQmVXMvOIjy+SNIoqlbyyCPYBT
PDt6Vmu992FXcggDWWOjzeVGKrV4jLkQK22pNEOn7wIx28SWK/yWu+AIP7DIsjIu
GdYTZXa41AjrDMKHBg3LuSwR8UseGGCBQVHBl1SnZVddzQumkclt8XrCY6JcSyfA
9IMxnfTept1WYbTQOH+kxC3RsqOS0FYkWnBlJbekm/7NqHxA252LSo3MrhEBpnWS
2gI+fXPYW+WZyWnib51tBis4peoIb0yQPR/wXxomUtEIK1BIb5+r3Q+I3P01B+ad
lk0eM6biJCmwAA0Hq9GpCDokTUcm2Tw88TnTGLc+npBbwtVafxwV3Wfk6laiOndr
736RgOBjmDUDqWxIDYq1YhdqFnoVGfpQ7f1Agsj1SQsJ7zXPNc0ERL9qv/s7C/j9
yv0YmEZ243Gwjzo/TqwDMKEM9osbys6yhR30XpZYK6j7odpCTVZ+kSi8RbaT52w0
dRSfljgOJ/by66KdAYmlCvf2dAyZy97Q54fUJ4+lrBfF1eGpmVgGl9oXAytvb3A1
8BMmHAzWMRlGXp7WA4eRAujgW/Mz/Vpj2LZJCYTPTrCEJCmNlNEojGaZ3g/0hlNC
HmiSuzjTGPfk6+67moAQ6K3CDrNdZKEO0x26QHiBvLWHcRAs97rPa0/EZacsPXs4
8I/qZozlPeL3qj/qPrIQg/eAZTdNxNM+Ol8RRCWM7YH1cPREXqXhYPOMVGNpYOyk
1ypPhVk98PkbkkarnwIrZbSGDlHVTX7zpemU/ci5+U2wLZCK1vUhIX6PRVgtH3wG
yO0aPOabcR0kNCROdB59e/6zihga4YZ5agonum6vtfqzT7GGYuzpVgj2VUC2YCKz
nSHPAOeKjVxvnoDkeipoHkl/EgbEZJIwRCQHuQA1ds1H2V2F66F7+IYLIP2VHtL8
7+4eHOAHg2X+QOahmPdN1f4ySeioYqqsq/3n/pJPZJhhB5skZB2FVZZjbYIwJAQT
S58ivCANix+r1Sini1RssiO7vL+/kk/Z+WOJn7yU4dupTAuWY97FkVa6a77fqnA7
nJaav77alJPuslwGXK3q7vVsupn/wBb8XikBXcXOXFY1j6l3KgVkemZ46aOM/nXv
IW/6OuhDrutty8m4lL8BkjD1fip5CUDBd5VomsYaTYJvDxrW/fdHKB9HWFvFNN0e
Vydss9cabJNwsOPRwhglBqMRL2OaKjdE2oXr6kQj/Ksg6bt1K6+YxpdFhGCncUtw
yWmrRoP4MI/R43rtsdydfdy8UpMKtqaPHpD/GhXNLZkcwVgDAt75hXG2Q/lp9vO8
HbK3Kr0jeMoust+QR9vcclDmhWO9CcqeP8r1YXWXiIwu9ko72nJOwbcJVOmWMk9K
t1dAb8okoqtxDkJUa8Vq7dfkLBTq4DL1x4u0v3Z/SPAuE8+az636f0ESwDcZD3pC
e1dciX7Ktdra6al4ZRg/CcTCbIbPuaoLneCKkeBbE616Ks1u/ko4w8RL+OHURqMo
dmRJues17EtCaTpOTXE5GGuroXt+Dw3UdBA7712sU61dljl40mmXBZVuW5ChxgUP
dqCCtqkeffmoYF73dTkcstUzj4Z+p2EgYHvlbU5VF7qQsH4Pmz8DOmFEw6Fzvxed
qTuvTD625Z8/nC4tIEFIVPlyNOm8Rp8/EfS1QhVZ6/vhDXLJsPA4HtvX8fQtDJwD
VyY0BgOtL2DRONygeWEX6TLckZEtWoREvt1xOTE/KSFPzHlqjjqKLBAV/zYG7WDA
WRHAX7w78qEGYcRvK5x+6T+qP5pejQ9K1Lojvc1uyDyUJ/AOinJrJK1TQRxwhJSd
LFIL5NVw1V1irRAPMB3nj9ClSm+SWx0m257zVda6WBBS0b8EX5luRJruy0LCJ0VZ
4v1lvGd68+LfCjIYqv/YBbZ3X0FtHqTH0FCHJM7TkhSFa9XtxjJWfIbeTen7edqM
F6swIencFVOSwsdqppTwVzjM0aMnIDgXhL5S4QVQRK5wupF6CdbPX1GuPn2HG3+2
gXXZ6vzht4QmZNDYCZ5dLTf9Rf7V6ieumutoF8w4JFsu+S9hFRzI7D2s4Tbr1maW
HU7uhlz4/B101Wyop0Ca7+IrKW8r8z3FbHiOT+0/abQz/xla+IFiLQqj3OwiBuO0
7zAJbM8ciuVYCKEkjT54R7qdN4INIhSBDGsrI2W62aHaSChpZ6gWVLhv79phk0P6
GPxCu4FlUngayOVo6TTusW8OIoOQ/2iTEtNYrkIdzBGe8Tg8wE0I2LVkcVgZtAH2
02ZHxnHaDbwynp8UJSib8vKoWP4INYNT02v57b9N/0ZgrphQnU/WO4t8XmtaSBVQ
iI4nkYnt3qfMAkSevD06rpWiFVPv2GI54x9UrE/oLNqdwjtix6efhJairW7JLSFr
QsQRI4S3l887RnMyaA+QAuctCOKYjn01iSofZ62BxNCTmq2Grzh2dahY4pLS8/8G
D1237+UFZ72cva1GDMptQ5CJz4/PQ4fVifZaQEQq5hRmU11d5TK9BKs3QyY3qiHM
M985qoglYwos8A2BrESUdB6XxO8NKCkD+8u+y60/JmdKgQvDmA0nPmVtEXNadoG8
jJVWJq6VcR+Udz+zMQKplFNPmnSgb/DALI8NN144G/FoKVtBBxp/FxBxtNagq01w
2zVHgpavhZJVtOIoLfB2NeU++Rv3iX8banb3BlM5zaholiHHbFkSEiigtCBHJi2R
B9Z6JiTGukz/+nxlhwA6fGasUKSz9FdOpuiSqplStJeRnB5eXFAmpXmmJ7x/Iy35
Lpnvgep2q8tEi07Ai/l3AgxT5wGkkb1C2NsU1zHWQNuvJexGIBhewB6HoqAx6xAU
Si9/PnIPBlOY5aAHl7mRkUYfJdiasSxKdlQ+9OHPQoZhJn6Gu0Y7I74HciLAWVRl
ctl5oLiwbejlXwkDGAGe+YCwKya6DHL0yxsXdY6oU2/hmtvgFXI6OesJomJsJ2Ny
FteisSIyk0fFqRjK/LNInRCJGojj7/iRIiQtrSvW/eT/Kx+OpsoyLgUjNItEXn/G
gCJbKsrDaz2R8gdrVEvcMM0XiP0T9JEnUdhlNB20SRX8c7mynD6rgSLMTXfLw7qG
R8eW/C84Lh6TYqgpwbAEAOavYwPEUBWDZwznk4sTeFZzEoJzvsLNAKtX1C7kTXDG
d+02xifRlzhEpf5uRij5U6AMKuInEvaPENpgiZEFFSTIKyojrY1iefuJWHqJhYMz
7EWXiiVctFIpqxFxuEo6yxRhXSoGNUa8vqmKoVt2Iy8eTM/P7JoQ6+96LBlOdV/j
pNc2Vm7N8aR/UJTdVX9U/Gi5+Dl54KXe9yTaJRJaRz4Aktovv3dkyYNF9zmhtBis
xgCiaE7XXpf5t0jRyODNUUpkZh35pEFlIu7k7Hlir1EPEggGI4LhqS9ITFXOZLFk
2DSalZbv/zictj01YRa8FpDr/d7VfxmZ4ZYNMGbKjCW/rx9aGwRLIj74RFOvMO7p
9O0NSS/5zd8LnHZiSUK5utPV1ZEcTkjyMgH1H64Fpiv8Vi5/O5kOHnvTal+Op31b
dqdQ4F7GLINdD4tSsjunXBTHG+YO2JnmPRYOKbtsfTGNHZz8XFIv41MTFml08nwW
uuspyP5y3r/53k0J1QiMf5c5IwictjkKvIrcD8OYmMLeuvs+lAWKnyBis1LYij9O
79F8FuYyGpu1z6bPn0nVg6en2zT3UEtFknjfAdvk1fYuKrkI4vKSP5hO83taGKy9
0Q8RLJt4yU3enlKQafl/Wai7gynljdWqwm2a+GqeH+Rp3blHbdiIt5c8RLTwrCvM
inq/YN8ECEl3u+fSSqdai8xWVCOvBIHeDk1lGklFKsBkWqvgjSjtsE9J2kgCzLKD
ppq4NSA3lLl0qrMj9xsRai4hmEW6V6iXmaso5v6OS3cPM1E6UpK8mHVrPTZqHJGr
VuBymPWk+t/39k7qnZHyxqSKjQdOORhOfX7GgNxwyZRNRe2S+kIwe0IBeLcqt3BF
Nq/x+B+eeZkv9YhokmhGNve4K+D9mRGkRSaInUDnCX1vEuk8JGxW3RrLItBRw8K/
ExiNDNcelhRs8Z8kRGUFs2EKtqsrXyKLwK0XkMy5Bw5lfMFh6ATKeDNF6Q/KwZJa
n2fJmWlKEC12A9saUSRi71hHMpvHrzrxo3ZVmazxJSVurnIpQ9pgUNeiLh+Sbw7M
RHQGaZzwXLQZ3Bgynw6ihPGzEmOdCV1fUIHNuXgHqWb3r9P1YGMfnB27rSiU0GLc
vlzT3lbqsgF482hHM+Fz6zCqTNVwRZ1hreb3JOCDqbK+Ln1OR4I/wI26OQAAwPxF
kLoq5Jv4Ac6y7wVc/jas9Qw3tP/1e9DNNP6+jtNmIPMxRqBig3CYLdhLheyFdfM4
7ffnJTQr/rruAJ72NN+72zb+m0Uq4hwCuHiravkYDiJ+U1XiLLxuoetvZOMAJ1FZ
SX/B8H8T/o736Q58ZzGfqxDs5h6xa7WpPDk1mcIt9KJuo2WAkj5qfVdC2lxrdhc2
rur0VipR6c1KaMVbPDteu3Fvho7WgH+WeLkiQ4cHiSLQto5Je2u1tb0K8pVFAYDv
IGdQfSKraK3sw8EjzeF7Oyj6OVUtzz4q2DtzTuPrJluH/mlWZU220a2RpYIw64nR
WDwbqXYKvaW1ZPrS7GAWj81E2hxUaE+h2yPHEowSeCxrFIemzvndYidiiNa2H3Za
FWDEeOGjIrGGcVR4E9TvRrnK16Zytmug/tKLiS4f2roxYlDiV4PdSZU3zACZNQdy
i+riwuRN8hBz/7LcJNDiOaa0qjRmyMcncoOCyeDS0K5d9JfBsq/tufo5BSxIJn4l
xLpHMRhVU/xQYRO13YTVnpcPkhVl8f6J4BeuzSzZwT+kuEGMsxMl4evROKEhQYLl
I0odj4HZFHwWrrI8h1MOcQJkaKHfkQSTeS+gZqSRl1A6YVrkpZ7zTWib+z7rQ5jR
3dSipo7CpZQfc0rspf6WQpzNN6zVBfBX5+g949g52efKHn/qfMMJ1SlHWU1+Hb4q
4jYhqRZh5tkCaN4PxSMinMJievDhX/LJn0xzfR4JuqApeqJZGL8vlfSFNsU6gqW6
E7u08WA8Pg2YmChEjzX+58qp220bHRYXbgVVXqpgpd5/POVn1d/kSqbJX1HwLVCT
KTatcwuKVp/ygU5uxa6b16awiEMpWotMU9cJ5owXmH6R/m0P4C2L8ZpnrIB7J8Wq
TJVFl1QlSYhL68Gat0b5RjcHW3GR8yPXCfAtr3+cxBQ3mFQP5ZQBAbw3WC9yPe09
cCK4jtE47Eiq6+N3o7NZ6gl7sE649F36vXgow0IS4VL05CyBG8qgsGYSORLBmh2s
xDQ8cDntxdSUrQMUL0+SXkP+j85xnXzpu4a1eNonXY4Xmn610Dfhrw8VciLRsDGQ
NsacvVCf6PD7PTCMFKKkQqnI88PHbqCvLVjsvTdI1LBze9ccBuh2STwclo6RGBlV
eatOW2BWIShz9a9M7Dp37o3NPvjKVFcgibPfi9CxzbYvNrHnki4BsgPYZTTFhfLd
AgFJFkm5JOoKeYQyy03/v/lEhanxXK6o42RntEVAYCoASl0H5b390tUZEQWUO4G+
K7koJlonovPBCJxKcU9Br2ASc5oBKftt8dpA0pzxpE09farhZArsmGEmEjXW5Ex6
P96/aF8UiOPmIDMHs8Zyne/83UdT3Gt3DJO9mU3qpggUuda0MVajOK/qKxT9CDEQ
EsUyEJRJKxrY7IrBth+8gcZ4Nau5ujFPX/zK71cyXnLLbP4kDgG+hAlcmcAjfQzq
tfyz12D3U7jRZC8exDDrClCFDW1iuSMYpEeo7LuQcKVXXwSh8s4v4hFt4mmLpbBE
XBfnUjdOJdOIbvM2zzoQroIMCPVqIYxTin1mxqiYc5LI/LAtCM5XBnqN2zrf0iiD
d60HhUFJJ8Y9AvnvAVNYmulEP22dNp7lYEkr7A9L5gJzF74uxLw3wh43mUTYwp9/
1Nzj6Tsyh37yxlka6vC0VvXO1tUIqGyKwcr73347UWjCH+v9/jnPrSe6st5JeJlq
coCUrkLRa/gB1Co/1xGOJ65m2qHBBmOoqlw0XhYy4QBukqERHKq5DmWmX0kgLl8U
3DsBKIBVXFgnGz4JhxkAhFy/K503FBLBNeGRbrYMIaUNRlBXj8nlDeLjTBPDcvzI
YggSNnf5WHPlhIneY2nlbba5Z8lFvVXz9UGPxuQnnqBRE5kcZWtcebSapJc5qtDn
3doTCtk1EyJG8/R6+2cRrHvAORHLX/3JVs1MdSIRUCQIfTm7l36h0jCLqd2v7YIB
g0WHFI2JyFfJHeFdMxxuh0kkkgXvV7IYJ8p9jMKYPZUV3+lkkuDzFH3pi0IEK9rg
+ZM7QIyALyTCY7gNfaI9u6sz2H1aXCD1a6BoD8RbaQ1ON48S2KVJKE8u8rc0JUc1
Z/QYZsDpRhK4aL4pyyXdej+rL6zI/U4UkEJk7KSQ/fOHY0jFmLYlq53CDcX1iTaj
IKBegYIOU4TZmWSYd4C6mi2VOE2WdwFAg2jrSDsGAz8FQS8KzeSYZ3kMbXUnLUml
dsXOSPGQ6G5yKJB6JX/6/BL/P4bQD1z8O4GKYw/vfXjVKEh8otAVR/O3cCRRdf4O
ZWqAlfPfxwgk662fcP6ifl5cgGNBDDZ17nJlCFwJk4rNyYrKZ9yPOvuhyeoYKVvu
fsxXghlfY4NQAWij9FMnGY37K9i6kTxYQG2KCLwRQHU+2EyB2mj0C3gnIrCmegis
XgtUbZrWAC5WQmhuGYtN2zaW/Rm5MYzjZ+eaG8Wp07e3+CePRwwSe6y+3/h1vb1H
ZLM0yASWOUCm7+xfQRLs4h2/w+1sLftKt5a53mUBDz2ACLPxQDE9iQoZ3OGujhyW
6dHCKch38yzuCJVxOVSFy2k2zDxD8sQ44i+LAxRxbJk2tLIwXuf46+iq1UrH6the
ag9Esr5vbOesCwsNPkVTtAsUXTgYmD4RcjLKvfcC438AeM6+DcZD4D1koMaY9emv
tifLMFG9Y/8XP1ec73pGxB5mB0rEsJPVXfts0RWFAklBhEC5YFhk5pRFC/vH5YZE
rUT2wNY9+JGU2/Aav7Vc7iwVeemCyqUpsXpgDbunL4VjmHJm0WwjeU8qji0Cjtjo
y+RhpkPdhcZ9tPBGz7b/Q9VI57nTGwc5I0NTFSSOszldCKFO5OdmUM0OG3Gmcbwl
RLgam8j23Vs6gaidq/Osk/dEQGwPmVpO+0pgZ5qNSoxZ1NtLplXS9ZNkeNbja+oM
GHagN2iSAdKO2Vj4ijZXmwARG08QbjZCer2Zl5RtuWim5i/JXg6QRF4oKin/jMHP
H/YA66B6sPnVljlsvH3/AywileajQacpiH6uETbLsULEOIOAWde0/H9HUJ3gwKk/
JBYKaBELQ3sdinEVhIc1jS4kX3aZfdmiuucHflBatu1jHvSsbD0BnVJahLMTl0HK
iBuVfuU1CHI+lQUhmZ98kzFZgJO2pZ0SxWhRIPAZ9iqu3iN19jXRh/elQHmVQsKD
sWR4LYHyc3ijx2kfZOR470HIMYRvZMz2sWpM20JbUYSw4/XtudGG+BTeApCK9lvq
vxqe4akbB4AwX+4VYn+Qd1T2HIdJf8stJ3/GLq9mKiqjFlg3OMOFQA2M31GtUPRN
+8J/4g7dXjaMZtrtx6tNwEo3EjDEuOeTuJRYEndRx6+MZRzNQZXo1cwZQRHSR1DF
DLDOolfw6wQv7DqHL2AmlGi1NXzkrXolXCggWIk3jbtZfzoiQNwoINtICVGMGBqo
tdBzCXAwLGUBvycZtlY93UsOVE7DIEvx8GMS/pJRtu5y/QsY+9dioDUaGlOE3IkY
JQfNiOmnfzC/uaVD/6jhACGM+PfzGZuJ0JoOubOKbF3K1xekkUJ5iDQ6zTQ22L2x
eXnsY6qQ+0N0g2tQlSRdYBg29mfj7UT6OeunOzwVLuOv0VjGlDx702tEkKQYTdXz
ADkOVBcVwvPE5Cdk6OdatB3n2cCFSQYghh+E6p77bHH70ZZC+rtQ6Cidvsin3/+z
bcjrZuNaqsPFuP6z6KQsF7pwzIJR0IDTM1pmvEiTHm+Q65Eo8T2lTjthnRONTjhL
obXv35pLs4o4iW1/NuxQWGwjLTHT5A/ib6lpW98+cV/RQgoIFFl5RqoNKHyXJNkj
PCbWGyYiw3g8cmmweFAOQ2etkQ+wTW+VckeHeWo2kxSfj8RjGUiSROtg7dEkaRQU
GdDFWb1HMDldjf/aFQTQCLkU4TQrYr49N/w0UTOf8l3uWldRdBFANOm5ReGH0bg9
3KibfIxDkF5GJBQgEif5g0piZhM5/uo4+rzF7YQGFucUMK1Mzigv7LSjJ6Ama0Fy
nL/LobSM+IVTMnM2n3x6SoAW8D78BQCHWALBJ0ZG4vy1sMjVRY5aPkm3QgvrSra6
bblK1AhSuz8ycwv6kTcX7RIGksxNf/f0L6elxjNG1kmMdFs6N2iYjER8DbpbMdyz
1tvqLp1DN/pw1SpRreLLD5NWD6g0UfnS4Du5b6hpXYjUmFXKiNgqdjcAPd0I9GIr
tXiHlD/1R076VoO9rwVcmgzvtFE643+20WJCCoBnFpKkqY7MaUx1EynedKcaXN+f
kGJgkzGkZDen54H/6+xePk7LsfDudgN4S7kWKUVkJULhQKhoqpai7vAzeffr3w1c
7MB03BaR/JA1DeGiGJNuqz5rL1z1mhJRvYuKlHNHrOI3drAO1iGLhHKvfxN+FV0r
3zLotLMOc9LsG+k5u25LVtQGabYfxCWwNkTILLW2YpsgBVaySyozci9fwomYzW6D
+TJ45RuXptFsVxJ5Yg9u89grXt9sIzLZ5nnBXtiTrczR4bo3W4xr+ilcQqcDEPgL
q7pkAOaru/NtZdFm8LQ3uROgJekyOriBWiOesZPZmycRftQ8iGohG36nJtfmx1b7
Qom810H5UTGGo0Jx1DbyZUdQHINZyueSIyNQatUHnzWM9rRqb16ZGhweyGLIM0Sk
0hluZBJKrwkH8/YSRRV+AUff0r3yA3xOri4zK+uGKAeawAw5sMr+L4LF1FHox9zY
jOctJ1jtWB12zEhHeXOfQGZxEXprpXHaTB3i1gV/fcw3CkzZRPcFdhWb/I1HzvOR
yzvIQ/2NK6ee3xPrUcV7n2tU/cYg0sl+umYtqMmodXJS7IyS/318csyad8bh+SG+
DsbYK5e37avYH8RLVMXTJHExPAJLh175kDKFecq+Nh3EibrXCqiC16BCuAcl8sp6
2dpbjulaS+YKXMpEWXpX5CjGybsVbdk3bz1I4WmrRo+YbwOxVt04JGyWEJfzyS6c
E25UFdjXn7f+AIeT34aU6Gsl/6lXCcJwG6NJprq/LRQvD5iNOvH1VfqBMm2J3MaQ
t1EXdVzEuTEGUVtzIUinB8dmYfW0GVT9riuh/vZK4SYg/oOKisbFgaGnTYTqoc+N
lz3uOGUqaWFOIIdKbQCgauh00WqnNz1Oshm/I7jDUjBolVJdHuZ/uXwSpqi3F4fM
0hRJtdcxX021bQe17UBZJcIB86CZ+aMvsFB8mhs5mrZueR10ix9qmnADfxbrRFlH
AiAVmlJq9KgLeDGbea/+9FZ5VG5geTn/YFw+bGol4xbg0O0x5uiDOlge+9XO0KRF
G54oKiSRjGiLGADW/pfdF2obYjPDK8w8An/mYp0XYPq9iaeOp1xe93aDf75WcNtC
JSoFBL7QV2vm13CguXXEs1NlP21cksRKx5ewiKcrFBl6syFPGpSmE2fuPrriss1l
UU4xl9XgzfSNyvSWkFNFoHspqL6twswl7PHMhAdeFS/w9QWM8JfQnwHZK9hjqFdk
MHskUHpkj7Nmgyz50JDCYlNYOfc6C8pEkFvW4DSxaV16BTMYmUNlABjeiTax7nDr
LlXAAcnDayaFT8+4sOPbmlmzq21sBd53ZfvCtk5J8uUUpZ60VTzTIFa3YtDTqLzE
vVAq8Eezqmdn4ekjuqL1szcG7OSLlKbSZPxF4WlifkKpjKp8NkgMcJGzJF9D9hdn
lLCmophuWJJDbMijruiCzasiS1SAd/0bh/dx46pWsjftE14xLP9Vrpxf60CGkCkd
n3e44P9IeqG6CL8umhatkQDC13f9JQ8cetZuIyrmiqNuKwwDZMlWLbyxmLLmzf3b
xa/PWq4zzCPz4PCK3Hng/DufMy0CdUbJov2IBgwxSgSss41pt+1G6pP38EB79p31
ALGA8hT21R4VVVZDIk1qsrVhSDm9CVFApFi5k77Bcha1v/mePb5FMzC6QUo1oku3
/uKTK6xUvdoItz9GC8Vs0vcdy6Z4XI3r6VvzFZpenryYwgiwIq0kw3lg8CwYeMaU
eR9PMljjNX/+U6IKdflsAAW7y+zbj1pYQrzsyuzXf/+9COMTRZow+uopumo6iFde
LKLc4epeBouTQh8UpOQib90/ebTzRmRmGujB4pmTdlJCidGOXRlEATNIk0GRsiew
DnplFmSq2vlyO9ji8dzfOqow2wrsRk/EUKoUqOsTDkbpCkCYqzwaH95AKGke8sl2
/s0sxLvCwpndCZ65iHj5YJ4FqzAmUHYzfEFAInrMZ1MPAo1rjl/U+tDnuzWhaHjF
HLftt5HCUFQpT6phhtC0yUL0OzlNg8UDyN8peJjbTAUs7i+SkgVHNFYVBfm5NHp7
oGLmxqp96daE/0dTTgkV7FxC5x2IwjM4CGrbiparyGh1lY4EsW834qVo/TRVoXnM
Q3+u30wui4i0T1h3HCC3j2ayuNCPAQPtmG0+zjd+TBHN/ogEHyfHD9ZEocYxYIQS
+ya1dsVctDGDYt6WJkdyGPekM2rpdEN+bqNMYFYjn71gi35LaBFFyHVuYwbC1027
DfxcYmuT/FECMRudi1KD7E2sFA28HXO8koysbEv+EQjoYT5M0gbq6FhYM9lVAFG9
Lj+ry0fOCqqJ/gqC9qI/PDZZdcDVP7Y2ga+EHtpytlPGP06X4hXIQ2JSt3IlagQu
CCM0o4j1HeuXezm7BjikuQQVbDzdLfRd6cV0bQac5HFSpDCUs17W8XoDsW12pIcD
m/CgQNEt95K4ePrw31D2BdZAEcj7hfwsGgvze/FZn54JEdDEEszyMfQvvbeibHc4
we7oJsWlTB28lm8YUz5ExLysfDnLlIUXBa2N+3rxtr5H7VxbAtPzh6atiANGg6AF
2cLoHaMekpYlRzWahz1QiS6WusMksOu++3KwPts04nOH5HfshCxjhnkZb2vVBwzn
1YhKyuw9NooR6wXj8UVFlbjKiz6w7ax14EybzSXkm5yy2Jbe2UNDX62ksnxFnKf+
qc8zgqWtGyf1vo53SLm3DHxWUuR/4kMWi+F1hi8qlYeqWDVXwhS4l8XqCO4ow+/g
xgzt/S5GqWnKO2vNglPb8ziLmijr3+/Pcd20RvhHJ7ASX6DXIy7+MWd6I35yam1M
mFU/SqLy2qhFwWlpCnK1LETwHGu/pckE2XkceIbiBBLVIHcJwHr55+bNeo7/542n
drg7IgDAvSfz2ozHLKTbfOkXdWCYNoihtU6Q3CTQVwyrZbbTclTFeVd59TjY/hD3
7IRlZO7aSMba3JaAe/rLk0dfPh8xjtASl//ZO/WzgAbnLcHwUnPFAuiOt8+xg2le
vJooA53xoQPZCkL/TYmnAeM1Fl5IwvJED7sgT6HdxgJHieCnbg+kA+CGJJN47Uf4
RPtamYG2d4K5wsPlogrZZ9F6r/2rJaH6pVdjuSi2z9KlcvV9VFTzQ5owbFgz53Pd
ly8yXNOKfLB5WBsbUSqw9nQIXQQyUqM+04hRwAwGCu1zCClpp4PN1B3TYkbctoFC
/IwCveMGYDbZJSaBCyd9737AelQsnnVh/SIlwdLF2anDJnp9BulvZDEYutv3ImML
8kbpuEYt/E0/F4ykyR9GttDj3AIM1RLkC/6kUkxMsesdUsjC/Ywuv7+/xAwAaIL1
jQ659yyZOguXIIUXW1O/5oudWYwNrFdX719kt6Mk5yTv6FFlQB0I3nrclVqttL+4
dBHcAAbmFi3H66zVcRrGH2kGRLYqri4Xv+tJgDXTOIlmc8+C/QJBxJWwFRrEk38B
rwOFjtJZ296HT2reXF+CKy5i1Z5bDnozkjZFo+xTooBIAQKiowM+78J8Wh5fN5ax
CrQNOMiq49ZSmxDAB8YCb2AdXcbEuS7gUXNUkxKGCypiPPG4iNnIyiBq0f4g0has
UJEYgP0iQuPd7GzEqsUiTbgGzHrSgJFY0swtm8eiQA60XOP/7q09WZP/vuAQ23eX
zIfCbaD6DrpZLJBGEvCniRP2RorBpGj7/GPhaEx8ESpk5bHIT7z+TD7Dge97Olfg
9+M2qPsZ9l5lrylVIulefe0LEcEDnCmiX+Dtu12T/kMDy+cLq5b9TEnLI3Ua4c/r
FbJgQs/PbcN5ymte8fLWlgx0OYNFrd/k1skTpGbeFaWyTcnu80gKx2xEOldSPyem
v/j57E6DaGmi99SiO/tzgG0iNlpT50hfpBj5dCne/kRD1saQqTqhdei/ScZWsDTO
3RVXwVMlrppgdLdHYTIoJ8U42EpiL5fjOciSdNxnb7+MpMuduUZ9ck0ot4LheM1N
pjLFit+1p1EG3SEEpKNeFvO51ZAKvxyHV3gsoiblFxScSADYW9nIKzzdkmwnEPaQ
118RLnoJ4xXIp2qNshMeAUgyPjsKnBtE4w0VrbpXjVx68Bm+6cZSSIMHaHwqoZSR
OaL5+2TK2uVLmOlYagxyI8gZdrEffBYsVKxsoZvIBzAtVyoffabYxHJKxJpmqMwY
jVReTBKSiOmycPKrLLapQo9v54N0K5nvZbuh4UKIzVHtwYOljAVq8W6GdVvGW0it
KULQfFf1MGjMyirmiO6/uAbyMFR0OGlnzWclhtgw9bse/qQzA9OEMq6DoYy+REee
kZXpttYcz/Lv0lSNLBAfZzz+I85G/NEz4VgkEJl8e1W1FS0O4tXCeqzLDCLXA9KF
+Gb4fV39WhQZ3tTAVzx9UwFNZ70aL0xh+mRDYpd08vuXV6W6HaJHeEJ7C3ikvuZf
E0zisheWAdduNTJH+0HweRakNlIZ/r8cWXRimd8YMKnq4JV8A5vOiyn4ceHd064p
8skGtVe8ZdBxpQ6NHXDI1aN1cvTvDYtINsFu0phoaAEhnYw98ki7rnb+VdRLiIg5
GlF3HAFKntGhB+vj3Tafm3NbLskyUKHx6VdIOsttrX/w31p0h166jTNN0XLnFuH7
Q7JKKBj1jatlSVg0DU0w1OKTs4jlxlzDreTl1HnfDIeyCaoaInJ9yYZgNNJ3HHoW
KqM8BtvMVIvpnfqUbAb6HLD+bj2L4IFyWvVJzPCeu/XHwznWHo+zAGQNCE/R6W0o
B++qEu6U7sJZYtarM4ykP0QFciiIYP23Nq9PnY9u1EBGHm8kRGyfWGlJ2QrNhhYv
EY1YKZ3l9T3geG5V5dwQqvrp97rakZ2vIjyWms9T5CDzu44LP8j2Q6HNojHUihb4
n1anhFizXYJYJ9nVVs22kphTrBrZAFHSNVbob7itOMzkTDhCKm8Q1pET8UwKAFn/
c477SFCyhjVJvLzxh4HJYoEpyw8E38U4p3rEU8fPoYxuGfSFSzBnjN8MLLwRUpnk
QFsXr1ag1YpGSzJaF/jwYStMc4c10Z6ywr5htQ9WNl/n9CQsQ5dHXGVtHEyJj611
KDxegYPbLqeSwkIi4jkTPoxTFSWAKv11MN95g+tol90FTa4niV/zUHg2qZyk3sSi
kayxm/HMyyjEwG5oHOZg57TqE7jYQ+K0Hnb/3/jz3LacqRMYT9LEz5Rnd4E73RPA
nIQUwa5mVCq3ihcYFcVZJ7/pPgL3qVIKd6F6uld1Fuq3LF3a/PYWIzutbvlHmhTB
Mfy6T4CG0dKg2K6liNkpEhgawmOq6h5RjW4QkxV2tIDwBdzF6tmg7xSm5ahHZK+a
Tyjaa7emsJPsEM8F82gz4ykhJm9NSZNn6tt7c81K7irwAEDqfbQNiQgLoky86L4s
Ha1yYaaOQeSo18fk5dJ6GFNRF5xPZsh+DvVZ4jk6fnIXRKUZcz0Urj8YLJwngan6
xUIsXlRVKOcJo0hIgYgMQWyu+Ndmw0fHEWhVa5OrWWNoJBVGFTKXElIGB1EDZJ07
vRilzMtqY5SoVJ+kBkTwEoXyJHtUU/CTUwEP1LwOVC5sJngoDcgoWPwF4NPKhp2K
TWkE8sxUgIuCltIV7IAdjMFL5PMdOLUPnhCTSu19K/bf66ynVg7oA6Gt5xufLeSg
lpOz7sNCMDaBGEuvPaORnmV/LnEyFBrXGc1T5ioTBw5VGQVv0LkVMF/TNmdUIYZS
ja9BrUu74IllW0MOaWjH//iggtFsgyzlL/pqQb4Ch1LU5704RQZyZv9ppj4hYyfF
v7cTvddnCTot9z93oa06lQM/+JIxqSufUThBUsfu3VZsElZ65wxr+/8ZJHwwLzH8
zC8r1z4gDhpTMeu6ggg+dOSM1Nes6wzxbfCjCLCmvIFLxa+9QM+63056rsOd1qpG
zD6rfJc+U93GnGoUYHY8lnVoGJVMpRIwVQ9YqR5QtZ4sER3BcMrDN8Z70BBBIw7/
g3Zeade40tZhHcIVPIOZvicb5jjDymEsCJeTZegBkjffzcfABDqjAEY7C1I6hAp4
ptgOQtyPk9sLnSYFloBV0Sc3t9nPybsMonerInMVpolCQYdsCC0P2U/RWBh8x6VH
W1UPnnz+b91c7C7OVKrpBnNNRBYZJOjKGUrEdebBkZ+uxkNvy0k0RCD4jeYT2USE
62zYrpfAwF5HTlvOBHukyo7P2DBCc9HL2tywYhPSjZuyI/76SdLFxHn4a4dkDPTm
sAfkx9FVTkcaMAFixrLnpIv8NV8gYxvOQ5B+jeTBucW4eUxk3H4HJ+seyAjkjh9m
QEbh+RDSRW2h+tZGJ5E00T8yvGY3ffEakXknmlKeQqMlFNOCvG7Fdp/Y7000HplI
LyIW3r7wU9A+CQm90Qr5dHWH+eF4XiQmVBm+lLqjQt469Z4K93pVPXtOu2KZrgco
1zqxGvkwR0mruqZeJjPZVKK8sqxATY/77riAKIIFeOO1vEuZ7rWJUo/W5gv8VNI2
aoJwUKnfql6yVPO8aX+Dj0Dmo9KH4TJ8V0ezOTsfoDIlzE+e7kpW4NiJp8s7mdct
E9r7LvO3gqUG4KjryxAzNuJp6YM6hC9ha6jB6sQ8iBGS1Kd/fvcaEcMZwC27afNC
w8KkPtHMsbQNO4BTvNiyEO7ppHzNDmQkdrPsomA0F1QfddMli6SZ14adTQgrWgwu
wJTwCvjQnIpkyNrYk2yrGZbj2argP891TegNPmVCbhi/beTTTME0ya88NHWY3KIL
N/nsgNC687NrBGd4DLxkDKlO8WvAPICD4g5ib6dgkLlY/jb0NoZlh4FcLW/wJVYj
APzxhC2CHFW9aTxFnc4jmWQ1TnthOxIvKlbomgOvmDHtLj+louH/rnlkiW2UIr33
UnN1H3tH2MmqUi8bPZ1XVwQ4zcV/mt0GXBiIXOzTX/TybT5L+rwnn1+CvXhIZJO1
1wqVUkD/rmLHOSTJ91S5I1KRs21EZ363GMibxHhOWMW6zUbMV0IlCpUbCDsKYkJm
yj52TVqycYPiD9z4Vt18tE+vesvMQPjbTVuPLV5JDgcvQpEJ8VNEXRTpEPqkTGjA
8xSL2Y3yitReQWy611AMAfZNIgn7CF2EHdtaqEPRUDFctB0C04xLkf2fO2856Cmj
0Ew6K2/pddcTOmn2BU7vxbBc7uXx7yixg6iFDlwB9qIiMtFD9ur1euYoXdW3adpC
kkKLCe8EP48MYGmY99hShx1VpHUZhWLO7MLSyT7eeCg5fNhpS6T/duWzvFF2P3s7
a2K7/pKodYV/6QAN85cJ3R4gqwT0oCTU7ezM25kS9SRGZsX5qql6IzUKvydsXJe4
YDkzRP7yXmetYyJfvzhE0HqyxS/jTTWrQvqEdAnlQvB6vF8yD1gK6mAvKfKm1XXc
FfG/61oUvDucuN8oa2Ec67TbOF2gW0Ojwd4N4wxJeEAtyLFTWCOFnvzmzo5EzrPi
8VqbOkBrcd7ApkdO+7TVBL0XzzKYnb58D1WWZxMd3M+3+/DOXn/BvkQG0YMC9Y0Z
EKH8XDluv+XqoeGUnSoMS12WE/DKOC9wZQuQYnBM46Rm2Uyhuno5IL6Rby5Z1wA4
L6OELqJiPLFIFQkwzk7G+6vjhgc5wL762krNcwWwOBWYn6ID9xGKFNDwKBl3qEzl
8nbGA0e3WHwa772ejMvYUd9IMF9VPqm29Y1iz36XxiIX8UtIp4dbRdDh0dC6c27N
gJpdUELtqh7ioRkCAzWCfo5oF/1wcZ6VNU4T2K2aQ0Wlh8BimTJ2RN4IJvBDvaSV
PY/QWT2rMfP+DYgy56fA68Smf3XMfzwkxLE//wm8o/YNCrfXy56bBuffekrwIXBf
wAmRJ15Xjl/2dIdy9Inkh2U51OsBdP/Ic8Ia6ebwCTM38lVU5DascBR9oOV2n8UW
0VXKPItb1W4IGSSySzgdaxmE4n8vG4C7sHXJ6yuUIR0dMSuO9hXUXdmgWCei+DxB
qVKQYEWO6wgH86K/sDeR7QjsRiqNJ6bz4Al89LokLBGZuJvjutKslSTIJI3bsH+S
DHucKJmy7Xo7plW7ZNT2Ak5FzBhSJ3I6HGfSX+ZgfkO6hwwXmx0pZ/VTPt6OfPFU
fWZoSjYvx8jh0VXMHcSdueJh63227oBDtyHFZkc8f2cvEK2+XFTL9cRaJeLVQDod
BgauYrjZTLF7FVbSDhSgmeaqSlMVpcrojIj+foVoJn0p/Dz9aUWxH2k4LsjFbkZ7
7x37LkM6MeY8oc6y31QpbWu97Y+jIJvhi8bnfXJtmhTSpWzJgyFH9jc6dNZRBxcY
o1Sy3rMXJrkRjezNf3mSD+P7HnuXTDjF2vgmkyd0HGd4/W1psOaDUloTrFX/jAeH
KQ2M/UIvY3pB4e1Q9JzBuHbhpUxks2+xvEsYFyq7hkLxgJrXzNW4PFURe0wbXRZ5
mqK62HYGHONf8qTIRrDMRV3GhybrLnPesq1nKpjOm4jq7hxa3hIDs7XJn0G1FMp4
ClwCJoZsHyPjJRMQetNov+HrQc2t3j0QpJwW+Q64cXrjwzqic2A/fjpY6m6XzJbi
3YM4aG5FDdTZq+2gNy57wI61L8+ApNjwTyGJjbJNjpJSYDWqFZ+xUWqkYvA70ZWl
SwJ+e6PtdWrJFaZeMNtjaDUibxskRpdFk57vOO2wQ12Uh3/dT+w+BgrPR4k7UNIC
nq+E4z2xCGoxXBp+gb4j/Sf4JiVHRTMJPfNLaTU16ypXcKg2Vpfx1AxCC402SQv+
DqtYYvqOcDUstjBdbBFfI9JPMBsOUS2K1gRg16o87QP6PWdQ6pmtv2o+vYqOKyhl
tz58Hf84qfJAd5gwKEPlMv5mxOpeiyacml3t27KZ3dg8Y12MPaw+rE5nLwNkUwhH
OJJLBEHeJNbpooSinc/0rnTLRrqcRPp5eQU+6jIUb8+g4GFMCKb7qsTCD3eV+qFB
fKnQKXfd/fGop3FC0x9T/MJnhk5C9qdtd/nlptxgNOSspYDj/cJ4/FwA8mYKFgrP
sjqgWECtGLGD4ziwQM15hCWBkOxhNOXji74ty/O6ObM=
`pragma protect end_protected

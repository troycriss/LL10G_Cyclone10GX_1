`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
To+tQnp20XRQyYJZF7Ah0CB62gF3x2bOLXgHaeAoDFKNskWPVNX3lXUHeTENb8D2
UBBxf4om7gvaZaPkeaUCaDn/9k5BgOwc+/LG/qxtdo6uZBxHvzaR+Vh1s229WxFw
HQ2pIfRBJmsPSgb7pVaKcouyZ0TWS1oG5FR7zKFiJ4E=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 6336), data_block
1PIKUy3bLHU+FD5RAKUGcaVYOo7sHatOu7Vhz1odNioIEL32RO9tPCf5yjxUm7zs
JSwDDEvV5rQ0G9nHA1DxaPZZExtFR9PlvpnjrxrRr18mvxrehFltpnM2xpB5v1s+
g+mlGV+OgCqz//ik+r3GGx/vGwiuXZBe0iQ/D9CtmhqBk5rKCB0PPFCVxeVLQJwE
P0j8RM9lwi5nSVNwf7K74P5xRl0zr1zIHgNSefi2ZowPZGMYCljg3pzR5IceSjbr
wDbLOxbx+QT2ZdA+AgV0p418aj1RP97yx4Lqdr+aPW6Z6L8X5ZUZJKyn8R2XuIRP
YN9eJMK9FY49eTZjaH5n8KTml2w/o590D5iJieS+Y0DGV9B4m8NUvtRT7rQymtq2
txL7fcjFmfnMqoSQwliIDrSEHUkPBLUbg0i0RwY1sNxmq+2l36U4LSW9FMqdeMrw
8GIVGXl5o+A5WOGcfXSh8YnAIJhanVFczbXRiGJSLwF+zudZUAnfW+lU4gXJhwQp
B1odkpl/dKcrEHD7QxigujVFlxX77si6xYBPd4xq0VyKttR2t9Tbb4EgB8Kp7YHR
s9Vc0hDoZ1nZoXDU/d3Dink511Vv3N0PUs+WeRSLSSOf68BBAp+GOlFL+A39V+R9
3rb3URXtq8qGqDF3e/geabGS3Yk6w+VhuIC85BhcP4N3GEU25nAK7nAwuIdrM9ak
DTWbnVJi5ULvw1pL0ICgGmvRAALRpbcdtn29EeCULWvegrd0pnjPHig4BjHec/xS
ScyKB7O2M1oFGnOAnBq8aNrYAJ7ujqSwk2h/uK3NCN8ex0AEH8CeNfoWJvwuK4qG
7vpLNcz26l8PM/flahbf9be27dIy7MaqcAFAeSsACXyNG/HBA1UHKq9cX7bxxQfM
AThMf+4xQCED6ZnXXS2OqMyH9T8TRxF9pzvrNlP+yq0zBSZBzQJcIa/czCzlkZJo
3oC6Sx4YYq7hZulWl2KOvzSedyL2y2W+NzSY8o5FlF3pezHrDR2HBzCdF1CKZhUf
2kPn3wHFfNhcx+oAjaGxEeSom1iVMht0yJZCtvi4BxVQDiP65natbzmwMmY6r5MQ
50l2KqS6gXZI7lU2+0bkJOzHN84wqKwXLxvhlTxoKjjqhWTKmtApa+1maY6X23gD
uY0e7uP0CsSXWwVZLEhs4Z3GgMpRhd+fs55YWdjTRvgKQwHw4gCzFI55/xk+EyB0
BsaPwaSaQQVAuBu02R+nYCnnRc/bpOo2rZnhv72vgSZFCEs5TVrusGNQnMaCQAWO
jZlBtsQNjBXZVJJvYYmh25sV09FvnED1Vkp9wFrvy8IqefJSKrCthA6D2IESHYWw
XFR5lu5b+C523Fw9M1AH0fhHObOaLRYwg87F5Rf5VZSGCRzQaaoALyTX2g4K2QGr
ZWSYcwFK9sSa5pZgcAFyGVKUa88zXkIvaSYs7byBna4tEs/3sybFg2obPXyONqZF
G9/K2+uG3s50euc764SWVjBixZTPfROBhO1afDfM/U5CX7jLMybvGMcSQGChYdFM
rQD0nLBDHg/JpITPzsryedktR+bXyzWTgUWMngpzdG57GkyE676z92jzOFZkrjBO
iRCcIFpBfPWhhqnt/SO1Wz4ZwW9VAUpyAE3sbD5e5xovfVDULKsjeiZ7aMmmpr1h
WU/q/nfNueFQYbzP247+nLsXmbsX7HLwucv6BlC0NICQQOIGYyDyRMZVo+KqE+Gv
2Ltttpba3UdnrwS7+JbJuZ7h8b79261yXfmwLqcDFGg2FLRYheN28nRfDgR84Jm0
MVZiwtqbIwdezBto3KE2H5iEQC23QnxER6YO/kSrmM93u3rsRC+ewWbv9We4wYnt
WKforfGrnJqFOw0b9VkEhYl9Yjetxx2+e7tbAzp5F/I9cMNhp6+EgkF1IEKd0sXh
DNwcgdwxuGigNA/ju/wG2YdEj6TxDAQ26OMqbhxCOQit7m1rNCML/WaeQsbZCSuq
defQAu4ph8jVAaaas2rK63YZUW1YUjaiaMsieGP3cHjydfvV23gjpq+K2DCmWTQ4
hb7xIt5DynNwJwCIYc+OtkiV8sfOIfSaSJamRnlyis+1YXi9AHzsS4QfgANoaERp
NgzuXO2p/eXazB/s/Yi/i7qGEN7PsCk1XXshpazYRXcN3xT/Y5tGeqZPGT1orMSU
8tSkIm4+gstlGmJLWNysjdghqK9t0uNJ/scf3p+Io2CVNasedYJKOi9dDi84Favn
97S1qYpN6K6FFRnO7bQ7HX+d8AkjJy745gEoeEEv1mRNuftqyWNaH7Xc4fCTOGfI
aBKb+vLWiExm2osILMSod3IXyKb6rnCnricRvjl1+W98Y/YnGYv9SiP0pXwZE+0L
OLEIwGdi+riGE97HejLtbodj16dpDDp2mWdl/l6nL91nTDRZplrEJtgYZabNYL9G
d0/+kk8n7u86aofnrJlkjpGhQnLq7aiZH8TXnqVoEhUwxHdyAdJLTO14enePoN99
6r4JcdFPkD70S0FNvyBt/UuSpd5vE1jm0GxwktPJjRk+pIyZgJo23H0PMvOmKXku
y8yIHPokZvaSRvpE0gxNTOg1CH96g8RO/uIvCJSb7NSCobnYsibOegQ3mxKPVT9l
btZnrn4PYz+yQobo/NcUIz9lfpwEz7eEGrUiQkdvZTCypM/Uq3O29g/JFc3OLBJP
z3+2BVC2bfJeAmcBDEmHUd9hicg0Ncjn6Y/PNuHAyryIclBXWCdDeayy4dGLv9M8
oepX4H1TgKQnTjvBLBS+3hKazXEW0UajhoNgF1BWHlS13DtpfyRpBYtql4OWOhgV
iWrbSEohD6ik0OOsA05LfqHFSJjZ6IEv/v7ywhTusQPSdSUv2lE7U4NnG2HsVCzI
CKD2DfZMb5jhrlZkW5fiEiozJCXwh6uLzJwFdbe1ROegJuxQN4EyT9ToSFcAB1zJ
x374CicMK25cdmGeVCFZWe8ZUyEn0sFcmJKn3NILzBcJHICIvAVmo1g53BQEvR5a
60T338eoVFZ2xhVQeR2RoY8E0jn4Xecyduyrys2PJSLDh1n4m/5/94UbhdDLH276
B8QGxXyK9sWBIi2a8QXCM61ns5TlqJgpHHcAZE4uKqc2zDNAKfQkZh+RgXweFlBq
++9GY8jSSnrBj5hZM9nc8G6l87Bxh8V1f76uueSg556gE3cEXMGpPM59wB9Y0Y6u
jJSdX2tSrBaHwlPPN9HPqMmg5+Nl9MK9XJZv+GfCe9/DA6JorjCxxKU8U38xqzk7
E/jQiHrXhogoGyp9UzRwe36C5vZyHjgjWeuHQ67THtC0aYtC9E3InR0N1KoJBwdK
8Br7bfEatEf9GtqJaKR50IQ1QCpufyzelunS9RMp1axEXH/Q8LjGOMyhtOGnxR+j
6ZfhYMMOMGjs0JFMlO3WvDklWEbuNH0JLmGAlDTTT2/c4Jvb7NjFaMsBfbxFZL9s
La7JXyWIMwlCkktA4dk+uXgrV7471blEA7l+NbeBi6FpcNELezDFZ27HPXALkVut
fchvFLw2mHB7c8YrimTUmd3KrrdR6220Dze6sGIFjqIkMnfS47eCKCA7RZypwN31
QjZV2Zq5gz5ig+Fdyw0zpNiqDl2RI8UcOoWNvX+hmDHv1wC7lrEtzu9Y1TPvLRKe
n+lhjecYWo+idBg+7Oe0QzelWQsDgswbZkQvetdU+cs1YHtG6IBWYwAfGqyq9EeT
v3y44800BXMSZ7dKL20WOva9oB0+QLXjbWmukaaZGYQvEDon8kXu8YkIlPWQXcR7
VT9Dxw73mUlelSwzMTOOT2ruxapZvhaRoN23rwk+cZhe8PQi9h8IBBQIfDSaM6Bf
LyIrF/m9F6lRYZgR2606mBk7xV3yViEOf92KLTtwi3je1DhkSLwfFU8GKGDiJRD4
oQGtjd0Za8+dR5853ahMdlpw+u2Oal5AbOIYzhCcQFu0KMaSLQFxpXvk0Ev4gHxK
ivesZVVOKC2uLxFwVGFopltW+/gBXeoaY/j8vvuhli5Uq+UPMG7FcW+W0y5ubH0K
AaZO7pq0XmDeXOYL8v2OL+0sfPRrWS26khboHAUXs5i0iOqRbH12tIZ7pR3zBwA+
Je1JCQ839QaPFa+sJ1NN7W+RCyojsLqr3bO71Z829Pi9TeOq0uvqMzo8ONPq9lFR
YSQBf8O3CfcXjxaOR5EIBncq2JluFiGqOwMEAfQk+gTKqaZIHsV0T0ZEiAf1vD8U
e46bPCRWmxJxLmalHGQ8Wp7MWOlmDKNxDztsvW7YiJ37KZCvHrxMj5h00cGdVrbG
cGeyoXCO4CchtfabX9twZkGrz8wD3/7rK+TI4zPLHbXKiCl7cdf8nRu2QWQrJ8Sa
aD9uvQk8T34njk6Cjp7tqvne7Fe92Dq+sqqvngoqvNicrq7dnBJW+yA5WiZnGsYR
sUqwPh6wFbymFCWLAYYS47cM7F7mxBQatNxNzfzF1Fg0DE1mF70DimXTl0WHbGQU
v96tNpnc/yKNSKHNSy6xsuvC4eYaSqGOQV5pvklb1bHQNflLb/yvGBzxqj3/3Bxi
aRjwwgi9gOqcqwWm6QXONKuvzvlQ+7ATWu4NHWbNDVa6lqPe8oFj2mJAxrn4hbsO
063HcvEx+KYJlajVi0k6DQCQx75bewPKzyZ7ROgCtKyyVdt4sqED51L7u3Lx07IC
/L8YGjkFMlPl8pt6w7Gd/JHfQIYR0yEYaIAVRLCuIAuJvbge2LwaSCLOnFdalv6L
ivDdGoSit9aOYuuAtVeZv3SEO3CC1vYFonbzoM3HSzoRvVQbGnWJLBkzmW5681bw
FYnccz+FhKrGDUJeiFHjnuQ/i1J4qFuu9AFpLM8WSYInKv66QhISXuH+ThApWOoN
GzLi14Ll956RB4s6q7s8rh7Ubt2G/TNGaOmoAICTR3/tGrTOv3FMCR5My6R7+pwQ
kQyfT4rJivSO972QEIN3MIMLh+ScaawIZUANoD3DNlmhZF152Up7xWJJQrn/STRX
i4X9y6as/2XshHcpgI2l+StTrvf6elqxKvD30uKmjX+zXcC3+LqFjlvGT5Pb712z
nzCHf2Bo2f5k+7r/CFu0xSDot20HpTsWctrG4ggiTvLeu2TkC9Aub/f2+kVmq1UJ
0QQEItfuHprLWyf3hQn+Nf8xz7qcxdgYx+H9xHCM9CwuSl9q8wy5wnfx9whSpWyn
EWX7neuinujtmwEk68sgj0m8A2pqocHoXKPrFpJT/JFCxrMCeJC7RNDazMRS8r3k
Z31xKYvr/uJUGeObOS0cjmJRGkJY3k1/UOsU1GcMyTNCp/VNNtjfLzsSV/+wk34/
qyHFNUyXWMravy01stbP+TEMNeuAML8Mvvp3ID2I0oo4VB0nKT6N8i6lKm4pohPM
L/6SLz72w7+6ih/FsryWwQ4v8oie6mcHmxjGRj9yNEuFnQ9B+8r5qF0xS/Ofe+WF
f7RI05ib/xvaLJC/DZhel6OHiUb5NeN3Do0/vWdfnDUU+ovQgVa/qEeEXiwR8Do7
YwHO2PfLZqUBad/Gp+gQadY2suQO9MEODNYWoQNO28jouwQl5OjKh+2gtEHq5xfR
mGm5Cqep/Ooq07VMFJ1wIo229KOBjWgedTaTa9db1ZtUrGKAwwhjqOu/Ef8eMuBk
2/jZsmesBaTplLhmnpjsuvaG8zH2Zfo25c6Z6p06PURTW24zGvGwuZ+4uytGAA28
Tt4Poa9WqVzX12pEON+ECx0JEoB79GxCHNiRgzpQFl8E48hAUocHxCn6wXiQkyfD
quK8/Aj9l8HLNQMQi35ADa1xy0ggTGqmqaofAKLrRNeeQWlH/W0ZRhjjBghni7GT
iuLg0+9PKxsBs3J9cJmUURNRXK91Md81FS0OHYMp1j/LAFN3xlrGEkQo2YeykefY
tY/7HAwLCTI5ANuBwy/zYZ3RM1tZ3QwWLuQHe09Is+64KkOBwdacaM2cDrD5q2ce
+vz+kaEKdcFaLR8SDCxxZk1iJ9kVW76t4ZSWNAS4WP0Lq4GjopItjnvovbqElqvJ
xa7D/Yq86seWp+NIDRa4QKzioXMHHqhC1UGBndcXlTopJICJseLfJ8safmleoEDD
4jZqdxsixhgPBadZ8fYY5sPu+T/6tF6BlOFGXxfQwc8gxzCISZTvupSpqYsvJl7Q
9agVXmmc2p2gEEK4ab//Z6I4oiW6pn5NTKf5TWzC5JQ3mgknWjoQu5lYO1UOr/B3
v/o7sr5GZdnRkgNn6CAj7TOoIUpQWHwYWeUTbewbtM7XdnjlZosFwv0sEDKiGuJB
zKkq/+4o1c+yJiFCqHxn3t0CPg0SuyYgzIhzSECtR5oYPnsMHYiRORmavyDr1vnV
fbM66TqC0n2Z8GIASHEyx+Os5yV67p+I0Lc8SBjCWo7hKAhbYzdWANpSpINNp/sM
eHtubGLm38OfJKm7TU3/WUvTKZVVMJjKZPmsIJruuHGDo6Ib9r3Ozeb4eYm7Of/f
DsTvRsGX2wS1Naa+5zemQYXsVRG9maR1bsc5ciI3wtpySXTzru4C94Qt4sSnqIJ3
wlzS0Hz+d/xX4KPFlid2t+2YpCoO8FgxgecJs5XWZW5W7oVXOKsxubDcBrRpXytR
5PMDCYqH5Nqk64NL3LipKLm3HoeDHNx25VdlHZ1cMzVsEqtPN5DGUB0yG+QI9pO3
+ovRlMft+holf3yK6FLY7F4IDpiQQgfo2HGCnSwjdv2zAQZdjDrd+LlOh2zsr3KK
8yLUSUWPea3Tr5J8qmDPHnAywRwKT1iAolDd27BbejLDxjqGWQ2bT0M6GksyQ4HM
2zxudkwv0JBq3JgFNNvNxVjiAjMcplJGjLLRrZ+/8IOJCuapJqOzNELwr9e5cj8G
L6iQ8W/Mjc0WbRYM49ilHwd6CYErl01Bu9SAV/T+RIqtA5ckbSm0H+oYb+lhQshb
94OlEyu60ZarR2QnmMVBcfdiiCO4foNoG8RKLZrJ58kdkI6Lu1M4OH76HKPLuSBF
I7Flf4AgjcDp4WCilmHeYDHzXGdHGYEvCZXoEj00t+gu7JVrQrIfNivMUcj2BGnH
zN3etmCuyUKL5+eyMBBTXo/OYWIVeX/hFs9GN58FAIstXzeOyqhpJOHbWVdZHPgl
dOO4uYM16u1glXFZNsxeKB+xqK2GwtiGlcREnKirVEcp2drkXju5xq5+gJfWaBiK
pc74Y7rr5DKO8pbfGiSV0kUuwi8oE4yvxTOBOFw7QF6b3gea+mZBQBFE7gcflfQt
LYV5uegcUhv6Feqj456XGk30TkdiKVzKwQAEewSUZUZl5CnuKBYMIbY4AJTahtyx
dDAooRSTuVF/yEFBw5hWmZo8JjyMQ6Y9qFs54bnWrWRaKLND1Y61Nwhi+tFcpogi
/SrDsyPojRXqBYR9fIFugHK1OybBAle2uxSNLR2F6hg6Vz6IYNS3duYgFam7mxZY
vfJxxIMGtzagBZGykwjfIYKYThAZLin9IqO1GWiZUmVCivpuVzJESZZjlrHQhjZB
Itecxuv/zkC+n4lqGTOULRu7r8JazVg/2ZMs36qUa6tZGvD5jtY8gazvlMAlgo09
zHZn8qi8Nx7CcL0QPsIY7hGQAloyoAl7xvbBT1v3942Hhl6cTVl8F7I8feT80tVg
28okzqlAuTgHemqjJALHvzszyo7LV3crxFR6e1EhBFjU/KNvpx1iDkRcOl+rlyT/
knUyEByNezg+/9pUgZGJMQxkR1F31TGt+zW048hLggCq1jz8eJx8JAxRvdNzJZQo
ov6QCtBXEiwSlDu20UaZRvg4uoywSDfTEyLdWN0fr1VTygoXzbZFPKGgmuxTjaB6
Y8tWZqmNxImii5cfuVFsl1yQZLTImDLvC098xIDPss3VQ1uTmcHsE22bkB3DtFUx
QhWTUtDSFaYKoOiN1v822PkKy6G18k6w3PRqOZXAlb3OuaciPhyDscp52Btaq9qe
MFF2Fqa3wey7C3hHLB5+UtxDAFyTlZUvhAJ/jcTXMhgdYUyewumIha48YDF1v7S6
x6V+lCcVdKUD1SF0AVxU6T26rztyu1ZnNZjaysDtHAskXAq1uLqsio5XZeTwtBfe
fBU1WQJO4iCkgssvMKx1SF7hNsRoO+sE6rHwrgRvjDVo5vWUIHQ+QHaqPfAyUDeG
tKU1E3fSWZVgFR9baVcWmXp6ti4IophhNMaAbxHrgpevd14JLlrBcXPrW+ln+HVP
szE85/VLMMs/LnqyJeFyggG1KYytjwSVi0jzo5TK7MJJf6cSV0s2AVP3gyipWKKT
GChOAFHzfaHNlJYbv+Vc3/8R23y3gXYmTEsc8/CAz9kQYYpARUdHgSGcXyZx5QO9
UG9AgKyjYiSl7h4qx80BxjnhgqE+8c8XTaT+fVmDetuJ8rKaYs0b2z29AfeOLAAe
ER4BSWcjOx3dR40wwnCNuY25wx1FCf70xn9n9nvyAHGRih708zoZlnX/sRujDPvX
`pragma protect end_protected

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
AS2h9+OUgyePC9u/7P5ff9Xli4yc3qUkEr2ZzL6r6vo90nO6F4g0T17rNJppMRmw
zGUG4aSpvT10BxpFCiUb7WTdA0hMOzuWhA9DkwrQ6HXguJs0AQTDn0VBHkkUfvAY
zyGtBpTuU6s9VfI4+0JC1nzbkj5UWz1Eiq+phocuBxw=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 21904), data_block
XI1s14iONAUdDzfwviMgN0yIFvCUUt7z75uGis5VADa76I8wHVJKkmtt6wHCsAgF
3o7rLjisJdrAib/bG+DecnylKmLdtWbEzhmaonwk8YkoYZJYkoYsBlgmk+NVu8bZ
J2z59mOMFbnIanFRFO7qKbXXlK5U2Wo9SgCJTLFN9/pSe7NM3PZHpBHZjyKXhYPD
NxMuA8aR8XeNpSioH5pBobYxqZO45OEF+eDKh7F183JbNeKnERmRAL1pv1uNircp
fvIN0W4NOCHjxDkfFE1ci0/VlPEdfhmIvhxyMyTc1TtmFIshhtgdq4UKNuoJQmte
j0n/xS23gcuDdrQN6//HpAq9o/qsXem7lfllvYw9Z3PLwOJBmxEgqVNwX69yzNRo
SPZM+H0XFeGXIhPwgtqGIFkfvSGzHTDu1+Jl02/b/aVEkz5nhIcQuT0XXMzj2Pop
zEWfDT5mCSsKfl0QPpbqn5aDvC2h0wg3XaPmIAdRK7Ou4xPHPCJrqOEgmqJIqk7p
NtHHHm/Z9Pm2y2L8XIeNd5k5aB/ekDTJUVp42l9VlMNW1JThOaF1zck3r0PBCiZg
eS6g/9sbYcyzUVW1ATcXSG/PLl7Ht1cHr7EHEq5Bk/zdRYJctPbCvuuB3L39xAlV
zGAbKuMzX/tDHfEXS9XPHGqvRlCyKzYknPOpoWIKMdaNsGgYAZ7e8JdLdUfgJY4o
hj20cxEQcrZYJ/XdHNQVp24RD/gP4iLiGM/gwj6z5GYwFr1EYlpEMVbx2IJGGc4z
8xftQI0xXxNylW1dFaktdX2qXLga3zsDoTPNjG3DLiiMp/hqT2c93iQzRMbIFhTV
q14JzMvIFUgcp+Y3CZRwjS75Yc4V8K4gDMzG+Q0PPwYh5XVl2iK5IYcRwHuSc189
r1AkYhcdRFHNFRKrwW/O/tQ0zGQtquadFpZj3XNfPgRW9wrLm6mHgAz8T8fuJTJF
P/e9Yza8oiLWXg7pNvJt2E2aXRR95L3kxUueh2F4f3K0Vo2k4dVafUDm7FVCW7Ql
qSUg2EoLcOmSREyII7ehBFI0UTed8SkGomu++LAciPHX5DWIbnPXguIZYYvDIr2X
1grqOH2m1wLdC1h4bAXurc+yea84M8I2jOpU2KIZxsKpaQuPfQngksG9OGejqnTW
3Lz9QNObbOwT0qdGq/muZNmRbb2vutvTzO7VuB0zZVPX5IY6Hh/RGPmIjoebwFvN
bOtrZnXk5mwJ8DYNjPHxSJy6lcOS8vBMozOzHx/cYTViny1xy+3xkb3ufEPdfHv+
Wk284p2SQDcM6l743mgoTKp0fHyixSiH097W875SU1ML1ahpmTB4S25U/hRpc6v2
TrVEOo8jAM10YT7qVaai0T7lEcS9smoolJkmJQwzPvtqVfBIs8uj6M96w47+Du4W
HQweysaFNcLuVRPsbdm/3+FxTl9sMhmbmzcKdDdK4ai8fD6WAjLdgpJK/4nE65WF
YEOhIOeD/43QXb3B3p9HFF5eZPRBBMBgjn2SMq/DO6oXZ/KkJnLVmq9FigSRqe1N
ZIIp3LN090lKZwjssmHecyCaED8hB0mgrPKsHEKreu22rkzKm51xjh8Vct8iBQ8Y
8GpN/xwtq/jRV1k78q2TWScO/1bKj9ngQoOw3RmjkncmJXsOqHZ+hCTGr87qZDQ7
kiVXdItZzAj8fd4+UtkyDmeugJwvnXNmoCFbmPWbljX4A3WV5BPj2U1X/EGjlSZp
vmPXh4hoJejGZV2o1kfvz+YkkIkfs9+HMlPLVIop7OZTSXerVInUsD7OHHLLRkx1
acu4vNK81UYodREhg3PCpqBMrdkIGqqfH/B6DA2EKGZwIWQddsCw0rqo7OCgyjai
1TYsebqXIWwWPtSA/UqJfym1epBAuDHgj0npT6UIiTHG5Ps2lrtdR5b2OuadLZL/
5gkDqSoScIBHn2QdTv7iAw9CVbaFvsV0Cm+mOzpHbJiTbROF1LRqVDtvCucz5Gsx
tXef5FY5qWplSRAagYjD8mLuzk5dNIa+VZrEfqpkrkiS4WoBGS/ntpHbyPLE0he7
TlYo1XE42TpmALx4IwEPz6elhGdPzWMs4/jspoRi1ISazVMPf0g00yS8JgWvgeCp
mAaIOvN+C8SciITut8swmZnbWegBnh9ckUNTXIpnubHsGRLUBMe19nac0EDEA4aT
pyUuMn1nMEYeeyDQL/n0johEvz7M3koifBWP3XeARX3OLeZbqUzCMi6A+8lGQ1YW
ViDU3JU0sX9mfpTSzXgqQxENEj1rscKdQoDLW91I8LoqmqSF9IQK92m/K9Lk4/l5
BsFA9XYHhXUAdeqyzcN4u7CaTrSdfTTAty1uA5EtsCXV6ERqyGrxxCnlyjiuVzDF
Hmjhs7el12Aq/WrSxEQYaCqg+i8EMVmvC3csjjosvs3jCXOl0xAvYKaMbhkxe7hL
8OldsuKWsbOs4QMV1xb7+9whDn61itC2SKjxKhm8Ngo2ItT7u45vVfzZ1ewANbNT
AE1803EeTBeffoL+IimHd3izp6I/Lu7lZzanHluSAWE6kp3KG8oTprJ7vPPpD189
XRZISRGoOaAeyzaTPlJiycDCtXWwqfXCWwWXeWcFPDXiN26EfdH+dIGBfsVqb2BZ
NhPwq0L73ejfe5JWXzwWwgPFsmgJn+Gek9NUzR3fxmeJFDZM3GeVUdgO2Vxkg+lY
HcTgZGVeR1YkeB3RzEbt4E+B0tEoUtXPb5e+a6uwl5d9IdzkCr9J3YbEpDJJK/pf
w1GNjOKTYIuDu5dgQH/wJd9mDvdNe8/fabdSvDye1XsqhizjlrCshDoHtgGKmrMF
Fm3A9l6yUL4PPO5UQ/ClIObT6q5ujv3iRokB002vyeRU4hxjeIhVjBe850paysMc
AOefzSEk2adaG642+4GLg0str6jQOesg5Y1NXcQjX4XakhjuREKBqyjJA5VQUEok
yko6tNPwLCHH0GePS8Ge6V2Lyev6vsP7Tu24/kPS94c5vDZKlod3kPdMku11dU35
rEWxkf49fkkUTwEu9OHJM2cQkz2ykTfjEENilTWit1MCPfjz3tTZX6vDJmJqZEgT
a6P9pCqzEYg/1ESDD3LP488XRFSAqQGbQU15L7vMTfy5X3JQPRfV6575eIQkDBcL
VwkgG2vsEZhkyLI49KvTNLW7NBskzThUffU0NZNdjdbRzEiuwPnffVfczdcFvpvu
pOy/EP3zfmwxPV2uXfw0QaPleJDiBHbaT8d7WOPQ8kaYzXAMDk7K2BafYtSkL2SB
+c+eykUqi5tnEG+tOon/X9Te/7oFxF4RaGlQu9cGMSGX2P9Wdms6sdjuxJhbBPhJ
dNTs9HelQ2MCpmtJqdbPIU2bER/+xXg3xKiZwm73ySkhprdSbzDI4pEVkLKNI9Cb
56Z7HRWSZ36ivrmNSW5AMnvkmPGHNPScz/5qyUlcmEmFMetuz8jOZJLXg7E5wFHW
LCOzrvocG6SgDJNPnyDmN8dI/lr0JwbAHoEKeA5KLbxxLKGeklvAmnTKmhNlY0/v
eJhQuwlHXlbW1Llcgp3eBHYirBVkiwxhpw+X85+DF82nmAwRXNatlFrdHsVKY5+j
wFUKny+SRztRZysiyb+pQrMMgFNJcjbE5TgjDPgrLM7B1vfIwcdvhcnpH2XT7X1y
z0/tR/jgRRxKawyvnJB9qr5LhfB0T5wk76NoG8fGiO+GtDZcEoRn6s6evlAlZHcR
OD4nc2ldW3Km4nsRZGr5fjQ9+GuChqmgt7OQ/T7mSKIO+8u9HWLKFej+RGTjuCiy
NHCJmlof0k6M6Qlrs9YBo/vFd3PKT/oUYqJh8fr14aDnRqIxFtYwTeH2tz5iJzG5
b2I0wa62Q+LuP42pJideDbDHp+JmEu7HSwuVXglTBlHdhB5fhlU+gcMHUzbtdfHf
s29JjF6wIRrz7DdNTPzlMQ0mrC2noDhTOujhoAD9Opnb7GFy+lw6xaTHHB7hx7xS
LNjn/t3h3GZNDozlR2EUE6QKJMbAPEWX0n7FICjm4VDHzl28ZiUcjNme4s9stCa1
cbo8DAAyDMwpkm+jgr5FfQWumd85ac4i3BsVFvF1FPA7lCCZjB0HXSnmF2odDLyI
xxnReSKIKQLJyhm34XRncN9Ihi6RfoLOLSRGYRLn4YUeQcnGU6tepJ4hplsELhRK
WKhj40CnJVOdDG4d0IvaL+ck+kpVny7DL/4abuaS5CGJLu1w0Zciz1k9NPKMCYg/
EqfeVI6mxH+PqayAPAgkf+BAvsuqqFPwIUgVNXZrbcnwUMhLSadiRaXYi16wfH30
k4SYO185XoM7F+4U7GdN/HIahr+gMpi8f3URsuYn35e+If03OD3jKulqRPJhCrKu
WYHsbaARGw0BiHcfUrx/kjJHpY91t0368yNqlhMz3EaTWCHPU/aCRU2cb5azxysM
WWc1Nr3Y5u3hqmDye8kVjozE09ago4LjhLXXtwLtqPXamgY7dLVem0cRNBC9lZ6O
bybK0HQ7bYT9xTSk33dcI8Jk/ElZP4W0abB87sFX0lUM3P/3ZtXlUhxjNInfJQHn
TheYoMOBswN2s2sLLjlbYdg2CcbrC9kKTHa+TkPsl4RnxwPww1jMJoSlJqvdEuXD
8+vLuoNCwKsQ6UUmZhMGGgs1kIgxNFA2AlVnAnuQAYXMbXrN1h7pf3jRicAB7/Q7
YST5SDimkMhhvQpWsG6JM7/rf7iVdy1S19zh4WtZ3hciBDAC9xU0Somge1q2gjW4
YhZSzLSWjc8LDt5YmWTSsCsruk800zDjoYO1RUp9x+FhfozS9K72eIKyxTJB1HLZ
hUybo7AgopFmsWYG4Gon9B2BX/x2clrWoatLUCXvMhUyTy51ERgsCAQPETsaaCj1
VvOeZdVd2Cm2+xvoM2ucIw7CPtFxJAPZKJbNo5BWx/HbbRFlnYAD7ugojdpaURxT
GewBVEK/x0XjY7CpJ3CqsdqJxCd+liLGoixLOQfzIU3WtM8gggzmBYMuHXNrxgcn
xeb+tN7SBOQ2gQsw4+NXJ3xcYmHc+pNWZDQF+Jr8w60ykCJ1uwqU0P8LXLXT2orC
IzQqeYsZrqa9dSAq/uUxxR7EX0CYEqRr4Rs6nk30xzpGJ9O9poooJ+jJcxu5bMbw
KJftGQcVsDYpVYwy5LjEA3b+mrOYGb3miUJqUnl8Ulmnf3VHtiG2Wd6KpeFpQ4Ep
HqE6sC7X23jpdfF6Xaqn9cNTTRzbqUlg7JgLJI1xikk9wXooGz/SMJbAOBDv1mA7
k1Nfu0pDiW7CbqmRHk53mTkVoxAv1iWAtMc+E7DNLqS3S4PJ9QNZgFzm2Nwst7jM
6a1fwsbJwv7FgsomyY5FevauQlP/QmjQSYRaW6fHJjmLxNbnhETp2ukqk4AhmdDW
O313ErYluuGnxmwysVkqxOHrL9eAcXVpvQKu5wIYdPvK4N9GpqZuNuEtF9mnAQ03
XCN2WQKoVorUpC2AK9BKH6yCOtNXpcju+2ZhJYhHTM2JtzqWWxsSCLbac37a9eXJ
JZuw9b3SiyzZtGPzsJl4Kd8qNft4J9Oq0wECQsar+wA27TZ7s/D1ugJvcliBzeuV
2XkrvWKM1zhXt0zfkzq5amMeoeK0iBwrtUVhVOwO5C4D7qOxB4vDmO+3eJXaubft
3lOvLS7+S3O5cnV6no2g/PUYgp7py1yG25UEUtyirjtGAbjms6K1C23QofHYqcUA
ngbRRmRyJwgMqLfb1j10DMN2uOfEqCq975hpnfcVubFtqwRtjCVJ/MorZn9G7Oth
6ysgBGaA3C4JyJDNMArhQe5Su3BBoNMI17ANaTRvlCjzzeSPSjiJqRwmrVTs0EH4
/wL8ANQQcUUQuQN4CsV6Kfx9+7mudRySHZ1IyEFtvofbvwrwhpnT21LUZDH/4YrD
Or+ZDqLo7v3o1NVm2TFADX5Bbcc0T+TbbkqHj9tfdH70uVKEzfRsUwbCVznfcO8z
tqFFehVh7YWGauPmKXCqSc1fTyM9Q9DqQIsFAkVkaiHdh7SM2ePBYLghu3pLKi1O
c7s4nwbCUX/yw56N+sdbd6J/rBmMyp3gTFEojrGmPZXrVeRKUOxejrzCpa6yCYnz
SRlEIcY5I1oVyw9gAA3A9mWNGN4EQB668ysNDexK0oIh/aNulSkDDcJfBNfIy/ET
hIU/p7N5h5WnYLFGsi23SDNALntUCM+37cswi36qS0KfZrRhvV86ohMnYxX0D1MP
LmGTXWSYphcHWr/jn2PRJtsEwqUZvJ80HVtflooP5iRaNP+1Bybo/3NXllmfX1qe
BnxMOdBqyZ4KZHtB63mmcxB57Li6zb52kpNz1ZL6ArMCv0NLQasDADsITcbOga+l
PEBr0QPpJobKULWRciiVMgMiZLJGywRR73R6JwmxFLmSOHIHI7xqsO1PFFbiYo5T
vhCQt5GUaiSsbxRtuSaoqEqmLKiw4t204FHAzHJNMbUpvLveR5F0rNg9DgwTlUkP
iIGl5vHHXw67EFylIkdxEG3lUwwAC9vc8xAik/I3oZjqlRTzUgpUtowL0ik99YXe
+fKTTF0Io00nNoaHAG9GH1KLxk0velSb9Nrw/cnRuMEbUbSRW2nLHYBGsdLfPUGa
orcXlQ3MbUPXkabPMrNthH7+UXfWvazKdB/5XspuYDJs4Kd52gtMN51bw1uzjB1U
nGLP79IqWRVDMYZvkzX66z1md/Zh50+Ey5RVdLj1WWNRq/pGV4BHXmaO5kqUNOkG
oTPpqQWnbm3Ky58fO5aNx4zsT8eFwkKrUAFgV+K0RF+A3T7kqNzyxMdwdQLbTQy2
VwC66vZhLcjpAVjki5Uu5VBmFGaZxghCcOcY1+a6FjPWbAu9JrcDiIpBngVqBSZC
RlNv9izaDgDBWjCmYhd8MRroN3jfYo6vkIDeDA8JVIrexWamlUSoyWluu4f3JsO9
6wCzCR3MFER7TXIvast/vHsShr1fhtDI6UaFGWvO+PHGZIPLkYUkT4P3YhC2mMY1
lWUWObgmEcGgvfiK+sRbYIS9xHFkn2euW7z1JUXvATLEJJxWzgD53rJj5q24lVLt
o6L8hu/XtFDg6UGNXbHwgbx868+5cG4eI4TLiLKd+FTVRouKHQTXcknu9Hfg7Rw+
IWu8GX5DdyInuUT74Y4sixImsJviWqp3NZ0wO57P56WxQarkVcompRoaRxYg4fsF
Hh/p2X5OYgJzJ2oBKbSdZ++s1GjlYzH3bZpeZi0pOt9VuS+vAh2fDFpCH6LQ45Mg
OgX5A8ZNb6Gyiga/ydxQsfQE3sNdRlnCHLHOqgmULhg3wZEN9Eg7JVpQoXf/XGJo
R8Uo4SAPxadzUfea+OhqdJUsWfDZeXM1XzvoAY1CdNY50h4SKRgkmTe2gZfsa7rf
Ebk27H5ppXNgU7H2mLklnWa/lAkTqMW4tuIg97YeF21qdzLlTqqUYEGBl7OzG/x0
wiBwVUSkVdeEvr8zAZf8rIZnzvvUfIhvzcyW7KLR+Q/GeYscBmDd3XkdvB7/bats
IeIewlcR+snP8V6vONbZJuB1zu60yAvayI1QxStrrDB2xCSX331gMcBalhYni4h7
4IEO6Sp5wX4HFxeEXp1EcdIp+DHTw8T6dUMLVe8yWi9cklCtchgnu3sib6dzSyNV
aIC1uIzoz2LedjXxTKSpc4Qw2fMAb+/bIPQ2/HMvkm5hkeLCXXbUoEt0DGL4BK6V
PiIEVdEtpKE78U31uRkfz61tbsXdfTPk8JE1p/m7NGAhhXVvurQ5I5570tq1eOT2
920NEoNKN1BEhAUI29WQVGKqrS2Fy6KYPLVKmaRUUoe6nLQMgJqjtciW3Pkykse6
BCoCey1gNYc3F6A8Mr00p19olJvAK0OqBgAV7xBiJc0WQaVEycyw/oH8f6DV/9l2
yImEdl+jSCuIkd4yj0H6nXQBT2cLGKnnzId6WVKoGZg4t2vKEZU2csa06Duaf4ch
qEDilyfojBRZYBf7N6UApnUt6KZ1IRSwvhGuDlhZxiSWlEew1a4Atabl0BznU65Q
7EC3lcuemZJhkObQwA2AxoB5fuLJ2UN1hzwNv/en1373+0hmYNFi1I4wR9jzscLX
9qDPRl/0HsHxWDO9dowlbWD0Qz0+cYVbWneH8tONTzikvAXHMUn3jAm6cLwv2ag8
LVCS7/YSJbpEWm9PvESeb+6OT8xovYd92jm7oyXXiEwyNqltGqJVyRy1iX1J8Au4
mxuMpTxA/6J6URGIk3t/SGJ8gxqxjSFN6rAx1rvyDodxTqM38Aa0ehApJzHcZApu
TH8etva5kTGFe/+3J9QpQRPsrIjGbJn9letS2LC4Us1UEN43xcLTcrT8aLQbVHuY
VzZxysObZZ/7yYbr/x8eFzuG3ttoFJNG5XSDc1FjA9brFm1L2pvLJUaRxtEQj7n4
OZDJovKQM+Wg9VK7cHui3qETLNtSunZJQnIXAM2CZnQscjklQePIgalAE685Cf84
zxct8deWTndKSyqZCF1qe0mnfmgJ/w7gjOkTp3wi036C4RiSa9XCpWDwrwJ7eumc
TcZ6/l4PHdXGxw3o9CXWPjQiidO6JIJxywAzp11t9kc6H19gTLhfJDDO+E7amroM
SDdGBfkXOmKq8nUOk4IMwWagNehjdYTR6OD+uQas6df2jfawzkKLtThQfUKsJZus
ezROI6RsSvMo5hEwPDRmrbAUuSFnFMDvu+RCiMXcnjyaiAnubJhUEVpxeZcEbzp/
VHLN3tvVczuTMQ70p76H8jjq1AcOESaMKnM+G5g0ITC05Nd39cuH3BhhUZ7EuUmP
dA3oGOTFsmYte8dxRGbbRkbjZHca0G+E+DPEgfKOxJro09DoRD8EupmmyjPRcLc4
Tn+ArHkyukj/KJWR+4ZrQxcrt3m8au5FuEjQL8E0sBPXKSH7ML8jfRKyfq6LDpKi
oEQXcIqPlAD0zFZNIsaTZQ4rgX4+x8GXdkqsHwc/PJf2pgL6vHyDlW3o8GIjADEM
5OUGvasMHD8TJKs02VucuE0/UlbtUmCZQIpyxAtm7cFH2ZtFVElMpb38X/J0eN8f
KsEbI38THFOqhoAJ4sLdyyDvzaI01f47v4ruskjmdW9lbzo43Yw3BKB+Hjfx8EKC
b4mQZv1eDChqnac8Xai2wTr2sST733U4ms21yRJpLNKT8lIaphIROhDOERIQ+FO8
OVYkTUgyzQysC1UREadMX6REYVjQ3g+vrJvy6A4xiKyVAiMCjkVQSCyRH+XOz1YL
YN1BNa+b8gK/Ai++8S4Zezhdyr2GgfEgJyZ6iUAaS3vZqAycJGH2xH6LqmJsijc4
ZFps03+ZGCOMlEq9ipE2xTwcNACepRaypzjnFE+7TZM/WtK5zi2PPNc2Vx0ubUXQ
aWFLLjJir1nZvzxpcijkbKl/pF9Spr/NxayzRG9E5A2NK2q4FDsmEJYglxvrOY7Y
9ztHKR7PQ+26NhAOwjnxd2elEXYCsgsFeByX3JRoIMeQrNL6Hy3+8BJFOE1jp3Gy
bR3TPtJqE8ecqJPOlERgBgUZZ15u8YBlxq/lndlD3hMQ5HDAUah2s5eSmGryIIKc
YpuAGTjXfusepbZ+TBdaN48zJLHXhEUZhrs95NYl5sIC/3Xx3farzbAwtOcAXsHe
XFOj2NYlox/tO9wwj0KxRMi+GIua+lyhMq4yp0hAhteDstVDx2OhPnYAH3k3MVFT
lF62TiZ53CXQmZLjmdNxK25OqJhWPCzL5HA4xKgXPWkph6R3SvH6QWT9hNFSSIfn
RPrYge37Fsfi4FHUW446Ta4B+YKgdFBmvCcqNSLqPJM5NthZWVs8Is5e79G03C0Y
u+dIFhf7oBfGvyttK9Mv8+7a72i6bj7kSCZ634Jp3w9dKrsmumKcIXF3AghiAkUh
7nf1pvNWJt8zyH7MhZnX7QuGZZ262oVRHRmaFCBN4RgQVa33JnU2SyNwegnioa/o
ld/MLiN6iCdJgE5QzgU/Rf7hXABJqeYCmpXsAxbMvJl2BGWuTUKnzj1DwqmMQ97v
bxpq+O4lBuUMydV7HeZqxeGluZ1PHB2ObDSPeM1fxN532Zjpgi+LxYxg5bRy4rtk
KqYcTyq5z6ZRUX8Mp7DyGMt7WbVVyCcqXOY1rATakcAW/Ox1EcwLzcQBT9Pda/Fm
QK/Kaj/5wWQsyjlcpSQPBlyHZkZJtrgPcdDMA2pL1pDwxJ7o+v30+UCr0HFUYoid
nI+MREpdvSZQ2X8B+Ono31UrH9o4YMtBHAEXbGWVw2xBXMUXnZEZ9vL4TaD1aBht
XRgQvQ7OpQKE1d7VZ7a4Hc/xfPl9wBxepdrf4AvCbu65scVYFPj9M59aMHY394q0
WaXYODEANcNlZLWMPWp9tqSgVNASCaxb7eazoy3Hz5kJ1RVtqao1ZCWAlr7LYyRA
Iyq38t/RRVyzZeX8XMvBfP242+EH1OePvZOx6xw8tpBGNmJqzv3YjhdSY+IQg+GZ
qAjuMdASXJgwTiE7NQ3U3Xdq9ss3ypf2OlAzurrITkAAjmmCntnK87+oaGFeQkLe
2/idY3yvEfLoyTA+d+f1kgGw38HyUf6UuoTyGmn+wqOX59s4OpxqW7tonIoTBCn/
74sXlY1d4ITDlzVQasofUn9rJwHzAK6u5246rgmLUFt5gWprEd9iwuXiL8h5zg26
YF9pPTL8H1fB6nUs0es77UxqFoJNDS1ScWkgAKzq1z9LozkNmi0u9JV2VK8XSc7g
ehPN0/TTCotMqAbYaSEU9oRmx+KR89BKBFpS4UlEw3bk8CJr3Ks06Qzi2ImVuf7c
PxQZtd6P1N2KL2dAg0yqdDwruc+uMRoCqYxExLqSoz0ZdsAXbwqwh5oKfv9lWCG/
HVE7H0HOaKwAOZwph0HMM9jh78tws9+ro2ZGj6j7x2Np27jIDtaG+YSI5mqRBtfi
u44+fvwkU1KR5WEifyVLBOzS4VOl74s1aJPhWphLt8CG8yzx1bpQfpXhEFCHBQi1
QPkSomXgc1Y6Yyu5S2D4Jcq5yMVMsnF63SX520k2mFc8jWvw+um52nmQdOgRzfIa
FGQMGvgk2H+p5HjcLUie+rMBhT7R0PYu5B88/muGXwy5pePtM21rli8Uuz2NOADp
7YfQyIuRTiud5DCKeIDKfwR3KtbTmUnt988uNoIPGxenc1ItQSFMmIzJ+P+WlMTZ
l9V+m6JS8zQegqe7VqcYoHbMCO6FWHb1pZs8tln/g1UOu1YPn7MjcX/7gVA2bs+e
dxV/5NRPyJX1wPvEx569ol1TtrgY2MSzXKRfSevruIrmZvyURQojc8MroDxDjllO
knMw5Ow44RvV7SaDwT/kY6J/IggtoA+j3yCZdvmBP2dJ1C0rEIaphsVNeyJ21CzC
/bO1m18cxkLPVMzZoks2zXQIuNT7JFBe2aV8RMg1N1+YQ9XiLKa7rEtHtFZhYnic
2l9ZcVaRl6Tpuqxvr2LuE9eFVqmFHU7VWo0G2/9VaizZXgZrFPg+SibLOplM4CnE
GTNMjL6k/NBCNuSNa+52TiTFfmk7URq6MWWNC9JIhFNDEDMG8xu09vIiL+1khSj0
vWATiNQAcVkwvPWnt7rovNCy5SSRAH2DLNGnd9FrrpcIF27ngi3UU1+Kyi4/Ad95
nE+od4tdm2lYSgzEfkGlgM2HfSQ6Z/ufkD6dFsnp4Ed5AbeAqmjt3Q7Hp5yidhXX
9rftlfettFheNYi0qQWy8yhQaf3qYeplz/l1WC608MjEUEjzOAnYakUgJ+Hp1GCU
sPfByj+nN0ejyjsJCaxpLxsJHSh6+Xfg/qi+Vt5IrCPEYXmYI7Amb3Qv+634B1U4
A3oVscU2Oo6A+RzQZ4eZJdIZVWgVDEuBLzQzYKDEiHPaaXB2Wc8hN4/QCk8EI37O
Edut81XV2j9RIVbfaDaHIM4YTuXhe9YXaT3tKHC6LE4//E72mM57nTSzpY6ymb6Q
jBvOXXLiegQCArzX8Cut8vnPO2W/G9dC5EjD8XpsP8gIbD4Qmk025kRCBx8h71GO
uf8y6v7CjhvzrqNVaisdF+xMKIXZEF6FzZfgRVdYLf+LYl6F6ZcBi7GIxFfNqJEG
xhCura4TMQ7my2HCsutZOrIweImf+SeUgWbbGw7BGOQUDtn3TerrMaG/EilQw7bS
1hwjYwY/qzJKh6OcCwieYAjAc8WOxtAzr4Al0flpXE3uwCGgWtoBGrpzukjdS0z0
8NG29b79iEgdhsD3mOZCvaAgd+euR08BnXWQ2YENPRgGP0nwKVqsX7JBRmQOnwJI
z/AdI4kFJVwnjL87OsVpURoXuiepshIWMzW7tY2yuRfedWilXMz53a+NaRVfEick
nugJqPTyfBzsYuukboAZD0lljSbWAFB1gAgzF3XqzWND966aMn4fH9N/17Fg8pRZ
NmOKGagMrzSB+n9TNgUm+rGTo6j7J6xuaRX9RyYLy0b4XbgEExrXepboP0B6Atjh
ChCSR/ovUMD5IYmuvr028JYv8xhARfYxTwp0hWarLLyKDLC0l2Vn4CjhNWHtj1P9
QP/8NL0zEEs+k4Hh0foR3ENGeDlineOneJSup6W8Kw+8txYNk7g5ZKibrXqT9vU9
5h2AXfYQ5Pn+nRn0oj0lj+ybAdwE0VtOSj8+H1G89cIchQ5Z+DZsIp97ouuGoNUE
+0YFIA4usy6nY3s2adMtHyCt61WzdSs9C4bSqJnhyiewXBiul9lPp8u/q0el2706
+u3ENTHBVw7ZnNHKROFnzvkj1t0wpqZSby7j4g3s+dkF+r/kfCZqATVKp1XtYYRv
3mtI0qXRvaXhKxhVOpmUJ3b4OTGqpNDNePxpmv9jZy2BhCjZzwjtAg/LqOL8TBRk
fWhKFb7C2EZPNUOEorgLNmKaIndYt/oOctEP6YNkctd5mhZ28qr0tdt66B+CYwT9
FOudqFAvJ5f/h1MpdYhvJzZT248+CdyZbkqKFlLq9uMbtQ2M+blL7cI1ULy/GmDf
gGuBMbl4oyP4Uj9YLHrLqwu9tzyn7S4sh27BPaRalAqP48fm9fUHaGjY766peVnT
x7KaD3chwsnNN4gApsHAuH1jityzB3SH1TwelEAAVoCZRheWMkYPn3eGPLMAD1jM
esZtmoXf6+ewEFi10qjWYf0xHK72rB1sZmwPVLzQN9TwIATclF2nYhqtMKuffJ3P
IA77+UyrumRuUd8i4EArEfqrJv8E6G0vWGxaQrOC5GTFjfKzxqEjCCOxIk2EDfp1
xd6T+q2UkMuq/UXbq6cJokgym8ytlOOo+RxjjJQdcMLBPqOU5k6rLYJt7UDsExVl
hVevxtn85Qh3AxiugnxGzUCdoCvqOm/XchNbWNPhbQ6g9QZw9chok8rCWXOB3P2X
2HIdrX09szCyVe2k3eWdDxt0u+n4Ta9NvXdHS5df1LNgDEbaYtEqUK2CSjMCJcWV
XdBpQoU6kay+cngxY8aD244LVkWX7tNk7lg8WvahXOQYbQNgZBGlotk0QGoO2gq8
p76wuCPFjd4/cqFJNDmH1X6Kf64ESysjqUYnv7hCZm11g1UrOjAsZlDTWa0BPw0F
23KU5PzT7d76DYQNRNJuqku57nFlKk9n6M/C3dETfa+I4OKXkRm6dHzyxcoWVFTB
1JdHWV0ASolCM86eg3PiL+zXoKBM3ha5OCE+uHcvy1w9/WCputpMKFoW73/r4W0b
nQl45T+FiHoCWwA9sCIZ5VJQVvgqu/c88Y9S7KAPn6F341lUtHAIp+KuRdV2+v2e
9iq62FbK0D0IMlYLrX8+nF8KJuGT/BTTPOHgoBPivDixvLuHYmpFHSqcgYu2kpw4
YkzvltB+5OMLsD6MNVXRePDXdmT+thQuMRfZbtGGaS+Pgeq/O0/idTyt/PoPCln5
5qFk7OLnPEN1SCDpJu5VTJVUQFQpxGU3YMCPz0GwR0v7+8KYcTAGDiC7mX4LrNKh
uiPT6HicRS0Xm5UWindzVxb6QF57BNb8DaDYcMzM4f8KOIAwLnK4Z47jJoSHBECo
J763365zoBRbkO0ECdJb0mXUOkps92zsX7LNnltM+ano9UOeASA7qXcZToznvc6q
aobFOQg8OJPdwX1NJWJ1QDRkbkSpfd4ui+R9JvCeshixN/Bj/T1a7wg7ANIptjgD
bfO1yD/AbF9Gs+ZcHwCOApXpa70mzRtryLFks+x8dLmZzXRMJxUVlNENqF+0zUzX
jxS0v3VnhHIuB73FFB1afQkboY7mZwUddLYBY2fuJ0C6WMDrqE6VcMeK6tILZqCr
irIVxpZheKM1MqTPNqzlzs8rKAQJzlu1d8rC5LjepBClMi1+gNEHORjr9HgsNmHB
7DlOcMNF5057C6p4aKxpMwihQsxu/YH26bCORSilDyhe8DGmJ5a/X8kCbdh5Td9G
Xk+B+XHdEoddjECO4gdTw8deqQuIpKywXLPsbFDvOD+14O+YBQrrTFtrmZCijLal
FT38BQ412QLKZKuPBg0ASWdjwdxMAoqZsOzfZe5s1DfJtQPNePiz5D+qvszx4e/r
0fGsIK3qkkPtjEdyNrSoS+7bUQYqOJ1GUjvleOMnNynjYMs5UZRAnbfzSFLZUWBW
FKYUaDLZHrgG3nl3zB3LM4gv/EGOmCrIbq/FO9qSOXiKT5pUQ+dPrBgzq4p2sVFG
WD4pd1gKv+T+fJgEe3FW/QqQ5RQqgsYa+9ajVYW+gpCxnpPPX1PY54qmtOz64aRZ
UZLmq472QKaDR/+L5l+dpexLukcoA/kLg5NjtDeLeh57Wlal78aGr5EJYp5FapJV
YAF3sgP8rIiJVLnRETQuOPnCX9Qx5ECub6oQhjJPUqOB/UsLfbfOQatvEs+vKCg3
cyg4ElegS+mTgZgs7TPnG6eK6kBSVxF3n+ha9gMZccTAyKpmemxVpSthK2CDRrbK
KI2v+qMMFkkXLM+aAzJ5rlNBAGH0hU47N4LrOFEq+t2TMA8il2v+yaIeio5y5N8m
n1uMkA3C3wnGmCHYV95f6KDuIrilYiqpauS89UQGDRxHyfR2aDdEALjTf090rO3I
qPhdMnzrns7r7ySVzNabTklWWTfVEe08p9jX788nWgrWsnHCMsPbsXbzk8JNMJSH
oOUKf5CvZyDz5uPSQPszwObIh1EOV50CtPnUapOjK5J0HfQO0qGI3a6S9y2DV1Tw
KUTpJDJTrdNOJP8tGzf2gvlCbN/O8GZIeUHJe5wl2R097JpRLyJ4k+Hj/lfto392
fFDxxZRhxVX1OSbNh/IaS6nU95WbwdaLWHIyrdQgpkiNazpjSDPbvwv29DTDCT6M
6Ew78OmwDePPDtXR7OeBkJ+tN4Es0ie6CxWjKsWo9gWyl/8qOuLLJXnLyVi2FFGI
aVvh6GNFXIznsbgTlxJoyRBUY2lGTP9VtSvi2tUS4m9M5kZchwcLsoF1B+kpE19o
DCT2RdjXVI5p2HqE5xnGUjtwzeIFTwlb0ZZ/fEPbsmNCzlDQAVikcn9q7qreN9V5
RzQioBPDHH8z0HDDB5N33VuFkRcRritt3AwfE9T2xToo4SPJ+QDx6KVGFUSPSxmB
4oG3RXkbnnhtf+0w44xuF+U7643PUdc5VGvWUFc/jGFeRTPc9I7mniFW19HEFtBh
RiSLBBaa0tORJ5p/yrpcCywSH8OJVSrYnhFUoQgAxcf1tlmg929KGYST/1rQ96ct
EaUWMRjGzp7eL2WXXaJn04fpaMEQs9TwreT5rvUkI3GBKzXh1sn9XfOOR0wltTWX
FUvfEH8WRt3b/fwMo8m0FwLYgQUULa+fUMmnnmONJm5HKLBib1fWUGLCdclla5lW
O12+aNsOiZPNLd6AlrCOFD2CiNf3yql+CykpgeVg5GGbRS+7aWgIWDojR32foB3+
KpTolf+jj5u2BWF2xKdrSprYdgzL8Ruw3b3KQcfBuvcZFlkYD4Uq+bDSpE2g9nbf
RDF8S63ujCHm6r3De/A/BgDxaeLIcVxkDMsJeOWwrEKqqqjxxq3rszhxOMXt6jnA
1yX/5xi7CCcU1UjGMG1i6rALWWfqc6UZ6BLcw8Cib2uDLiuKREYfl5z76sX//0kP
0I4dYvwusxO1/f/uOlFGqkzU+9LfIpLGzASyzzFUHhjNU/P7vfi5KGhguYfygIXf
jiRxuJVBI87JarFBl8UJ6kZxtx7f0zDwM8RAu9IfulgwM93Z//W25ZkMNNFdVNJe
0Ytgiuinwpi1n7D7sQ1+QjvLkXVqZMjXb7hgYRDLArVM8J3fW/vfOG4fzuqC0Hkq
1IPsdAQSauEE+cnT87W5vIHg23BuLWoSqkO8oijRwEBfgF81qorv787wiwUNwJmz
g24s/u62ybjL9cramQcXYSWVQir48xt5k/m96rSFiNbobBbBUvV6laK1wFCT2Vz+
i1gREHi+U8/lPNz62hEB4nVWNUUCXhLOXYt+KMROBMYET4aQfrFpN5H/7qgx/9B3
M9XodzWKRkVAC5PWLMVInwKVwv5OL4BB7xzVaF9nFlbPK9oNHlAEn9L7EzGV3t9E
HB/rtwGCocpwyUbdIkTN3EGx/DokFRq45Mw5QcqFavYuXDoSpbajyWE0WChRoWcN
VTNi+S82svgAuaI397gKAxHoLK2FnTJdrwPOPSuRQtLHL6dzBHN29BciKUjkcz19
niMQBbCDZV+1jMqm0o1XuRyWubf6D8CYR4zMMGYkcQYRddHjOqRzkHyM7KPnHbjT
642Is493fgktgp8re14qME8q2cK/3Sy19U/2mDOrbh5B0hnXc8EfW0CYwmInJwgy
IvYl1QFl1mTmRFEKWMFgXz48PaE+woNcLL3txqHb/XRpOhVspqhwaS9wQyEFWno6
DkKuB7g+2irgqKaV1cTUsSRhuHfrtysTULpmGfWpfO9iZMHAo0iEEcbQans0zMqB
4GRj0hqPydh6OdeLMWRK56F/zRfcz/EhwLFPwRcCkeTYNzdLF8w3/vKot9pEpRkJ
O9qiHvdV8+Rwp+zEkOoC9+Iyh9ujhqwtb9S0apag/uOfXDqIAa5I/mp347ymL2iY
pPUqI8m3MLclW0DIrphCIzUlAjuokqnAqfQ6esbSg9RCBGusUaLERdQoa+E3mk6X
7IgzYc3bYquVvC3KX5Jl63BVAIml5DWdmCPXfK8clWQo1ZBL00ZnG6NDFffdG1u7
+syq07H0hTG27WtMzQ4wukmv3R70WgSsw+t1CNloSq2xFYL0YQKMm7rzIKe2Wnt9
lFQrlR+pPicsiajdlOEfWtvYeIm/t5AbLr/ZyAKVfuDcksC03K6UnYG3j9M+aM/3
n6E3NvD7c0tjLEhRlLq3LqTA94Z95pTH//3GwNwZUVwnRwcWehsub4LEsvsD6kKh
4wlE1lKzvQk+O183MrQHG8MPN90sqvOCulZFpV4Y41PDFpD/dwjHbSy+q2vdfP7w
M/o4U+B5Adp5IPOfkY2OnTWhaJlCUSBiOfKb5DWU0N5piaHXyPEd/RDMqRlvcYR7
B++C/sAIXG6ta9Sb+Yf8177ZAo+qpXMGSXllyDCTLdlNheB5GhqMQptkxZwL9geT
UJp7fIaztR+d3fJ4fc9WXyJhOJEjsU7QxOjr8iBjC4Vk7ZJFz/UiTCFmqSs0wYTF
vz85JNKijXg24/h3K2SZvd4Tp1+WmHjxaLNMexCm9Is3F8U2FKQbTmdbqjN2+yf6
QhV7laavkILRnlWjRubrXsYSc7lq9XzNsnlBDHPZjZZDGB+/5TWHnzgRWlp2cLG/
AqfqEVBSY59bGpeTEOY2bFwm9rDB9UMeleK0KklKC7qJK8+Dmn+BBSJ2Hlb1zszi
SRYkbPD1YpcsX+mg2V4ydydqWS+ofNVNGcXgDcj3VycvM8aNhCOJwbU/Bt9Atpdj
xXZsh49Sf3DrMor4wpp2xOsSR0iZ82Yt7qU6f5oAxzt3wqN+LQJbCdHz4tEEzI8x
Oi/0glUGXKjSpxihIZWdRCdxZT1FIEyGlh99P1uukzqQ8/rG9+cljHoP7/uwxPUh
Fv2rN/aaxi0ZONz14vZTHHciqr/58easCxBLzMXuOmTb2T3c+IcsCCMv+ZbFUOPI
QRFyCQxjDWbFmAz7ACKBYTTjMOxPg9YBwFnjV5n2ZrZz1RnrHwG1Lo7N0FzPdA44
USLiFWJEFtjLCqQzzmf5XOnmnEnl5aHdEek5rMHsn2NAILS3tnf8/z4m5QuoDgeS
X/FEp0ovUj+m/xMvx6hm/2hyHAnjN98NyYix8TjKsV5JSWzkEnvswI8ZhJDMMsPK
dsKRYiBYnw4ZYOrn7k4X36IaMu6VoTMnM0jrhSg0ygXcV5gzkr/dTLobXZ7Zo8i1
jA36WygogpWvOWRtDaAsRfM1k41xEshFoAgAkH04B7g84sao3LQMrxCN/rOCS76t
s4tM4czPAF5z00+Q5NEkD0L0NzcRjmbUlUSiv9RY77HXztb7PQvtkoJLNE8ZcyTA
83hf2VYkP5QYpre5XiKckUu3PNuEUReI1pjXG/uUuddXyCnpLx4962cSpL/r4iqE
AW0Lmrm0b8aisIoBe8Z8VxWrfWuYRjx+QZYzwQ6LZpgmTqDkPG2c4bwJ/Mr6FwLz
xfcvXx/3jOO/Wh9z8mR4I0wAgOlUquKADk8q2pkjMXT9dkhZWj80ufFtlFKOqRtX
sBgqIgU5cSgaZNp6kdh4/zvhmp0QYJXk9tIBuIoiMdIVXAMyjlKYAGGkdAc1RauP
iHFkQOauWAavoSeNcKq9JuB7uG6m4a84HthO2KL0LcYhfPzr7eh1R0gFozCcLLhc
0J9sbqg/o8nuSfg5ddQtat14nfSdbuHGkwIZfM7H43LoaatNrEOXAWF3QdYl7Yvs
udN3tNzFSzgOsc7JTCR4VYi+Xj78Npcl+rGhhxzNWBPYWJiw48ISHui7mL5XmH++
oRfK1i3U4tZJMOnNmAfQp9r2NPwkDIYJs3R9QY9A5WPxe4m+HxsfVBSIkXE78/tb
RQYKdK11+caDDbJma/5OwTcqTY5j/WEwhTjfB5rjBSTOK6c7QlaLhm2GM5AFZ7N/
UdP0vp4cdskaeqObFztqbpKo1ayXJeDy8vaMWltEFwECOwCtpQzZQhx7fYevlE6P
Q1Q+3aHxiLcRYUiUiRd8mo880FOB3LbMjpRyMpIuRZR6NLpBla4c54RERkAXnm7f
wAJJ4FpkmFwurUDaBz8NGsK36YdifQ5lgXCT533XNFMSBocivaoKOFuZ+IEfyjfO
xuiPmS6rxoDy8wiL74H9cs/OWXtVKmXjhz0/cdGJw5RLJq7BoKYfhMgcH65P99NJ
q7SSeLlqzUwvgj0CIa79y8FTBjF5xGpv6yIEmEDNS5lVbsmkK1jdwlLPGlxCDQXr
ai4KWVz6UR4m0G8PJewQxdgU7b8lGJrFYi2yQUBGE9QqmR/Cy8Wl4NwONdFUE/up
273Oi3X/+djJY1C03Tk1JeiRolVKBp6QGeeTnLH5rAS6ByhHKDpiaopUUHIVYY43
8saESAIC0R0QOm2Vub8/Z9E9QTXJIk90LxI1cXP9Q7Ag8/6j1G5QjroyBc5mh9BU
qsjLx8D+H6sE96d1ZS0SThgL5BtqeAQStxfnS6V5/p1pHqz0QF5dsDls7Cs8Anzo
6lih4kCa9uZRfjnLowYz0SwV063jAjV9KUvLcx7sAeNh2YKmhVzEqa9Uae1pJLGU
RmAaWL29u8taagyAZm5dtxNY4L+WWwCnMxbRi5KRb2hUW1xq7nv9DetWH7j1mZ6p
H6Wj3JIcP6nA7JlHnQXxsb3Yv5brWhoS+yVRrWbBTa3hJgX1bC0lkNig4g+6gkrz
EzZBvvass0O0zdo9HLq38yzf4eUx9B+n98HpdReEu7sT959MCPKG5ry5BJB298Sv
JMuyUkDTgiMM+p/YxW6R/I8WzWj9rvNKKDbSWbbTsa6dkzB9dClKVFCyn8M6ShsV
yQZsvMRMC2T+R/sJnhAV1e5OTz7r6+umHLqebqqIzmB0/GvqVWUvdycvE041Ymwm
sIKMNakFaOHTEDyNTWf5bargSeCL0D8M9cK4c1PGr9xDBrRYku7BAKYHIc8scW80
32ys9Yq0EFD3J7kWfAjdz2//1Jwrc3qNC7186kRBq4FIzCQh4WdeIPDCziPs1tk3
85MU0aySEMlAMPZ+RoHzctvcrPNolQp1RvIpFIn3Yrinf8XqKz3Ar+6AFHDVhKiM
ZPA2TUrDKDREPN2wcpktvdEZxG3m2uS3VDAZ3tZKHh5FEa/+P7iY4ui26spzaay9
FWyixwLjsi6UKa/OLrC5QpCJ4gSp4cNbVWUpBZ4mgviIoV7RXtcj1KvhxFn7crGW
mfO2FjwOBMsnOQzbICQzup5JYu6KlDavQigRQqzXHkuEX2tes6GDce01LFYl885g
4I5ZOkceppMB8qDnDssYclxXeCaPpz54cCCgQJcf/KGV+C4IDdvf3HmbEu4kjE08
GTSkvSceCYwXkWWpov+4ML1zaZXE5Wu718wcIbBvwXTTRiSqsVCuQqpnWxx0nh6U
gJfCVFwVQifrd8CkMneOSBuOAOdoltdjSy3sjW97+DpCv7M0IRLRyU0uZCSOoN+8
F74aZ2vimolUc94UGGxyKmKJAJ2yhbrKEkvSNrEO4L8wTip0I+Kgk+3Lo8Gcalpq
zWWc0SLcC3sqyh6G3k9LDADz8GYLDjNufk+Tb7ODRYDw/Ifjjw7FgOzctMA3VlhR
cN++7LHPCs118kRD1BpGOZ0BEQcnRRkJhJjnkr0GUst7BFCcXjgGgO2wwVNsDZhe
X5ryIkRIRz2Icn9LApRZvSR0izUklpbZfHK0NbLbHhipGkAgcI9Hyry7m20AohBk
LnH62SgaLtC+sa0OEvyiN6DtSrFn/H0M17uYTtuVdGt3vuBTbP8H00OwGI6DUS/X
0QVncAee0fkB6LmHaDE4jIoKXALPOw/WucBV+Pw9Kf2TJrgcbbsaweVl4rZBNvR5
tekxZwj2UPB/FRdEm9WT53gaN9V8UsQ6Z4pyz91DebOMJRvn49Ax+1L9e1pqsdl4
HKw8cZN5iHl8MIQDPVzwWLoAohSuC8a2GzK94kyQOHFIwRiZU1o2L7Ag+BlJmH1M
VPHKGHqFJFvrufVvEwk8j1kXv5u0K1krjFWfMI6z2jRTmQvSWDmImYLKFrj/pjui
P2r0NbhIkfmoYUFSdLvy7X8izFEs+us2WCEwvhnhEPuKVOfT8rM7Fa3RULPN2Z7L
ynX9R/dR5GQtJRGMcz4sy5nYfgigIlMOy4n6Fnh47SDK3KIIWa5/xiwvAmjpbg0H
+91yupqWbQhi1JV1dmgYcG8X32W24REkuZmM40GjOYng7wnZPjgCfv/kN4A15c1X
NVGOc0/gJFOMa9jRukUDQAmLxvJb0sBEduDrJy6/zE4Vk6cvkK4TE3wUhJcraxcn
bUyljPvM1wDGQtq0J2yVcEIskF1ZN5JC+SZPl6GlTzFAf/UXbdMp+zJ668GdYmt6
ep5xv/61T8ZeWiJEkzI0KDiSmZ5Kn4+8fhBroeGwqtuMNAIpLNm2DAgy9U6kg7GB
/dMSdB8OgVCUJOTShZDfozfWl6J3hrj+hhl4VyssMxTVJeGGdwPQzoKtJg8JYAZ9
Krtly4J+Xi0bBUCzw8C4prKNBOV1rTdPcjnw+zdLDfeYdqfvybWAiZDxy2b46U9x
2pb7XLYmZae6bKTY+f/DRgHINgvX1+R7piha6HBca5JdG8wzMvagdRXlcF4AxtY2
K5sM47ml06LMgYHlcuZJz3MdmN/RHIJzG0ivQLdlQsTyjV/RPdFgSZGKxU0i/stU
+u//TCE8mIn7yyOEa2w+MvaXSyqBgSk9UURXdJvnXbJTP2ehD/Kw3p1IOeS9Ik7M
jPX3MjQUZrzZzAYqa0lowGQD6eyFIxXBB7VMVZZlPMiIoZNzc2mh1Xh6otvKp/N9
Qn64XsWsvlJEIIidHLLmSDhXQdvP9zb8HBp6mpycR6D1fcLr5l5XSQJlt2dKv+If
QwCT9YbKqMeZjzdsrzIAAQJIg/6VUZeVI9J6c1OgJdUgJV3U9/6WBL8B4PpXcI4e
0Dve/VhWCTbsHJ4cH2WSdNGoZdJ8OpOxBtiYic4ykQtyPj40eneIAPO/fCnx4+jC
g67pKfbC1aq8b3JYsgLEdaw85klYOsIth06wM36o97sFBUX/4SYoA0zNDzoluVJ2
rPTqy0zbVyXUSdwFoLn9Uetp3IGZ+WsJm49+0siBv/eYVX6UlCHPZIfsMYG6CWm6
wMB9+2FT5IxIHwMNDpPD5ABiDARerenlH09GTuz2S+nSTJbwS6kEqfZSSZOrVuuk
BEbUhoAE+sL5ZFTE7MVDcfozhhjTcVohZtPAgY6AS8Xy/vL+YimprIR2lroz51+S
T/n9n5BiVgtbI6r/hz3tPpfYkyaicDF6KCXJOWKGkISBcHw0IjWs0r57B0oNJPZY
AhaVRnmOMldhA1YCrrlfemIvzvNsT0sXa/XrzHGxxfxJBc/aup/7JOHjSMGFUNHW
TKYt3QhmtDoP6YkTqaf9tfDDq3cXl4DEh8BqXWDqB3qDRQaIm0oYFY9a6ZSPO5h0
onPULqdZfnFpyk/hbnT5pMTIaFR+bsrrxJInmBGpN38bk20TmK9CnP6ACxaAIEYa
dGPOpQn+aVnr4gljVLnzz15rT9m8vinYAePchawJ+UTk+fjaQxEJybzrFF5t9uCd
g1KI4sIxvEecbtSJTwS6naj4VewhMYCDkIgfUFG4grZVKFfBQpOIdn7IDrVBSmqp
aYLujlMl13kXHc2V6IhHC5bvK1BFpyB/gphffGNWRF6oQhITaxEyWMV1r3HOzRkN
6KgAmstLepg0u/xD2Bj01p7LCnjVrJleXBoDQhdl/ldVjFw6F4qDrxueVrAf0v2R
FA54r/0UDxfB9VxH6lTndD+Ustz9a00ff8c/n7knr54HxjlQVYVPFUyaxVjHFhmE
PhCG6JAjzYH4g3nBh1Gf3hCTjEJcq1mDt4qUVe9FsdEluB78FJDMjMBY5TzJ+8wh
hN4LSZyUJ6pBnJIqW3ZJ71McmfyHkI5cghfZVvB5ie5NmXbLFBbQBVXSbZLPU/4c
RvwwrpqqgIRwkgsBKhjyxNrJKewvetwOVLsg6477e8LCasW7FyA3wGx1EdWioB0/
cJU5jWbRDbulluuX1jx+77T04qyTVxk4v0yzIRnoTkHbsMccSRci47VnSyLzPVuE
8+tUZgQ2Y4fLBoKF/B7PyniuKUA+x7czqSsKeSwqy9DXWE8HWAU/EZhyGjplJHRT
NpmeMsa2icYR0hOmN0tn3OpQVOI7cs1xdfFxbfovoVAPPM7i8iHgBot6WJbPJRR9
SN28Ai/B98gjW1RDoxq2rIEhrrk6E5LBh8EuXHGwurH25xJDukXcrCnK+c9IFrZK
GzVtRWPMJpRKVaHqVJbv8y9S9f7rCH2vUaHC+UAj3agyppyOjhejyKqII056fAM3
NHfW/Jo6wvPue2vaDPoLs7dI7qeP+GLVjSKAnk4tHL4+pUg66ojhnr2CHzS9FUd3
Dw8wBJUCQI2HvfP4Jm3jzZQ4s+1fwCHy4dYjKoeEO0W6BTlPEWdKakLBQSNE9TWj
MWQWX+BRrPKr3dA0PN1x6zkVaVuMKgmmLnnfVr57e8HBtquZRjFEnIXxurgA51N/
U2aA5Cxq9VeI0B01jize6DMPq3mJ5OKSUBnvlmG5laNMzEBMHN+Qz0p/FTuWnMY4
a9cTeVEVDSLZFLUBRmFqlV5oJ8YiUT+kY3tdbJZX/quUAxtru2paKdpOZARWdFT8
dxaZH7alXGxmGmijkKOss7JuA7TuvF/rUYWu3JU5nhHKKpD77IJ29wXLlfw6f1WR
d8sytceV0F0Q0J/Jm+jjWVPi3MnGksCTH6sh8hYiUP9h5GFshf3z0+VREPjRwT/p
H3pCBXg8jsTdEjHmumEUvp9DQqFDNglcXdBe/J8g+L1g1ONpZb9QR1+KAY7tw3IX
JUDdr8KREb4bD7Z9LqRZGHq82XtHFCr7vL36fWJ52QAqcut1ozbu2d8cVo9Hjizo
B+9aFXIfLM56jA3H4zIx+gyGfOOKXBUXj5EF2Dg6bgDGSZIybGhWmbpBbqtAXBmZ
IIdvmP7SW6DEg9Zp3oxBq+j4QR1Dte7bK3+eC41PZM/KqSX0UbFhZEm+WALR6w/P
QxY6NP5/7iqfmsxsikdoITjOHo+/EFNOiI5brRNC+nJpmD7E6K8Lkrv4s416riB5
AEQsLQP9uQy12kt4l9sxH0HGCskvUiS10Wl9U23RKHUan1yQVw14/W1fKOs2UBoT
rZqy5NhOzN3yGuEXh6/k25anzAbFNFT6P+SaEBzx765dTcWhZLxOqu9DzZh8xFoK
c0mN6kR0dOo1y2Y8gUewPNKd7Lt8CPPELKt5cWo+u5kahbjC4WPbUIV2R9nxFr3G
WzFEJ4MX1nPT2PLNXLLFxuOg5WEylC+6E6QrrUWhD/6iahz0OcsyGOfkJZpkcfMw
6jjM8SKE0qa/s6hmQ9T3yWV9kuVsckWtSvVHk3zZ48sM4I0ETLbpNExJmaSPcko+
DO7KUVE17XTm+VL197tsjGaTTbf/jDUOie15SA5eicZFiPrq3LA593Ob8idIWfsh
JAO3B1XvN8Izr24yJlNSkKSPOXtD3ieFRBx/+st/CUXYHpbya7IazIDnpLpFKBk+
jCHmdndDbQ8jbz32f6QIrLNb2W3P28zJrVlbmsn+e1LbE9co0j/RlNYnBgQySpWa
lRGt8CoVsEfi/fMt90K67LtC+U2jZRCxL0Y+GPV+s/vuh1F5oF4DpeCC6mm238dW
QKmUF5uc9+GAg6+B7qjob7xmh8y+Uv/QlABUQOT60EHUlLgfl9apS5/luvbiCWd3
WT2mCmQTJDDm0yaZLFzgUsy4hD5jDmWs4NcOPPbaxbRgK21DUNkxJrxpXaMRrKb1
0JL3JkxLFWiXLB1373HVSpBvrqmUmm0pGR6C2JN6gzKD0Ka6fdrjlczfJHVw6Hs6
Ju2O4sOrCq3bX8kyTZBpHjyn2L4UaQYurvRQst2FJPJ8XiXFjxdxvtdeE937RAMi
WuHG42JdDheQFCk4gLIjRDM55WXDJcCmUx2PGFQ0MlwZz8zCyjV0qnLcRrbvEpc1
kdqdjfj55w0/m2YEJq3X2UoLbrKmNEVtuaV0s3JoFu7tl+dpUffvVa5N9xWZy5DN
lbephi2kbOeoU20HJbWrHJxVbor5eY+PwMsqrMzWGPoZba9+QU1wUd/jBtwnusUy
y3p3tJRpIoOJQrX2ohBoWnRodU3Pe4CQq6TbkQ18DyL65/72zfpg2EZS/0MzXXkl
8ILT0aLRhz1vY6CN7/h9Qy9COdMxg2qxqJvSTZmeAeZf8jMi5VO6o+ZtfyT/6vxS
mgvnPomh/HNXD3zDZcYa+8OfoFgJ5QuErMNECyJ0LH3l9qe2UYXRgRTdtrSDtAsO
p1Ci6VV2snSWFH7jBEis6JMNsBfG0jPs/D4sOIpdQX6t2kxC016ykZPsSDnKvjxq
4YtrXthc3op1tPWScjOonV6BhZTjFGoTF9VfrUJMtmxxUrcG2F1ldjRR11ss8eVZ
aDFAzPy5uMJdoJV16wWIimn0tAKhUlUlwEF45953FJsgvegeCMUoamtXtnygt+lk
iaL/cj9l3bHmrmYnmOfhD8ye3ruGbi5/4eC0csBwDRD0PoO0/HPKZ8dbDJ6bUFXm
zwctTi+RsM0Sf2vO6/DE4NhHLfPEnJoepAIgGnzo+H/PQXyHqt89KzhnVJGqoVvU
cx1BZ5OdFszuXLkykD6VGJdvdz2lzaQ14w/qztH9fEA4bWE4AqGLjSZPHk9TURFY
QUO/1tBdD2NqLjEzXMvQ964GD29JxF44u1d4OQ6CJrGh6Iz2rYSH54B1aijj4W1d
Apc7E3SG2xk1ydElt3+lH2hdmu7BsfXonqZifjUYUBSVXt1FVJ8ZRmwPuJTLj8fa
2mmvWwhOsg9Bp2JHQbbYb5uoFLh91PbLn9HvFCPYZn5js61GJt6WKQUmR17EMV+g
nbFwH8JMwXI8xmokG69p5uk7PRcBNHZ4wic6dEMSKit9DYwQSc14s2qLKTuhTXT1
iNd4peZQnjyBTkSpY9rXNAdS7alQDTxNykoShTxd27SomcFiAV8ZL76x++Sd013i
fhE7fbSDWIHDLleOTevO9RmyxS9Kgy0Ke/HZOV2JPz6ryg/TNFVKyYFUT92r5KXz
3nuW+iowmzTFHDWaMZP+9bW/p/YDzSCjsYMMiDN6DVpKwExLs34Kscz9ttHWTEkx
tus2FVI8V8DL89DBj3jcn5QAMdAZAVBeYX7vgId1XpbAxlCR5qHjZ3BmHXy5QOHN
cnQNRj1vtlDkMqHLxtD0F1RinNDJyl6I30OGvPMV0m5KLTAt4jkWf4MJxFcMgKjP
iQ6ruEDhuINXiJwk76c00VgvWtGyshmv65c9nHLN5Qar6KXe1X9unGS/jEm4N0u7
Dj5NzuXDvdm5HuYO6kA4UoK9OKfxDAz745/GJjNe1y19h/LGsyHaatqSFmuY5+p4
Lcx3eE6WgHr/TlW2Ubfu3BUBXJpUm6qzOQR0ga81JVpxQX8au7luxNc0TW0tu8RD
2M0iyzNKT6ReDfOSga66NVAVcIn3o2RofWH3Dk1t0vc2uOxJK7XuTQlYWkcjj/JP
ahE5gHDBtfDdCo6gOdHSr6fponxY2jf5SlyzTv9zug1+ysBId8ff9bSyZS2ICeS/
VFJT2cbZTFW5cfFMiH/hOq+M4p5qzwNddYKIHKQzNLQybweemPd8GaHxFbwjCEC+
o8BEaihNhOkqpUSCb4kcBZe/e899vrqRdrim2odrJBLXyKXLCp/Cmo8Tx+hekbzx
6oDtwRuuQ7TEWb1s85oBUidTxTrtH/PHkjsKgt1Mcuov0XuC7gKaA9c4uN80KsWb
uZUHPDzhIX/6TIDxQG80OaRfXZ3avfCQjCCo0oHJwrbwTos9j3JEKASgBH4kI+K3
ZZSq2ExNGmhGiIpapwRUdVIXFyXrCGPvsKP1o2kgBEv3FfiBxOeiFZZEDqetwEHG
qr3cn5B3+Vl1gsQtr0AUbC0TQaABerPwg7CnU5xiMRqQ6dAGoxbsvPP7aV53HhME
PSrjP4Qpzt7O/n8s4SXRZih/hWLId58mwIKoC/gTeqAcsSnVQPWF5HboLUui84Ti
YB+4H73JL3THYGccLD+9e8Fh8gS0/qWBK9dh9ifSgpsFbJf68pAS7LMWdc97xMe9
7cZ9LWS8CX6fwWGBuMc7HjLxRPDbRpYX04WJz6+gk+/GioBphep5/nXAWshW+VJW
DO21QpWmNelFg4r+q9tlpsh3CsJP3z+SCYUa4PREPsm0WtpPtPfDlA/HaLjsHl6I
e9GpDj4hC9xuooogIpDUYhm/MoTqn1qYaYtRzYMVt+3OqZbotK1y59kSlBdy991z
j/0D6MFFgdjI5nou60XOF3KfICaGYskwBsW2+6S7fGFRpbX+h/udzeOPcVsp8Gt2
j+eTYOqT2ae40Q/OwXYfj0EIyVzrcpI8DyYh2nkMXeMFnJBCZm0HrIF7y/6y8bXV
C9cpAHJHD+ohG0JWRKH+QOPXBPZ4dqmyMG3xpBO2U25Bo3QdR/I2Nb8dWiYNIaBJ
x+YNHoq9OGPmSvVe4Nr6CL7XJDzf6AdwaEAyDEAor1FyxLPvkc3KNFx9WqCVUfh7
5VMB4S9gSR4F1wgmIE5tIiGwBOsyvVJRVqIqfkHtCf+hvj3vz0EFAQdDoqQPe9Xm
ueN7Qf5ljNGW4mRkbd8gbQ3Z4mQ9TkNO7d1nAN2exB1j2vbFR4vrMxY8Koj1V+NY
VsjUfe30gRQxxkvm6fw5tdVrtr86dOryK2FGlQ5/AHhzTCoEHBqTz4oAKuCsocPT
JMbyRSdY3FDQvYn1DPrWIVyPjtfmzOzooc4LHdnRfh2SMojUuDKNeyJoaC9wcEuI
yTBTqjcEisj8Lm2y3JBjAirvkPlZmUwzCj9CdmaGHO1d0WUnZrzc3fqPo5NMJtBu
JyMR0kKq4tADx7Kw52SFbpnV69wgQDu6fOmw3NJrg0X6g3fxBuRICDhpvOVbEboX
hY7ZP1bm9qA13RG4CmB3jXO7xxfGJTILhVqG6lG+hwR5g5KmVZM7D03wPHMMW6sv
FVgKK3ka9yQtgXmyTNyCzhYRrhp5ibJx8M2UZOisoO/ogHbuX6ZsHHj9zamCL8ap
v3FThLHUVQpj862avoWKUgujUchNelr5GGxp+0HHqN1NEgQ3E77wDUYOMSO33SCF
Sk6asNygjy9ZImoAf0RJyy3sywJ39LJp1gi6CrMvFUZJh3HSx4Vacrf/ITgadHoh
e9kj/G8DKcCnAoN3v+25cGPQsihN94nMIG6APkoBZpddl8eOZonH7gYOguWi7V30
/moSj7P1O5MGApU3n3lrgaiPcq3YiOn25wZMVRDQ9ttMm5lFf9cQmT//a+2HsuXH
5Vqkb8IvpBKzMnivdW+BYreRZI7DMyuxhFthlJXOPUH6HF40aeCxmUMSsHdPTRcy
ZJecZdM54T5XMB9ND0ymHQMX9HI2y7JPDN+RBBcW6DaCRD/fO8gcRwde3RCQrMXj
QmRWEkxTnSUeGfHkgUOIbtYWXvIKCGrXnd3WVy4igrULlDijf4s7c9se9XHstxyX
PW5RYqZaDo87tLRXByQ7MfFWn0z+juinu45YqyowkhX1DhVyVlcFbbqynQwX4A2A
4h9xdbOJ4GGp6r/CFVXFhNzM7v/5dGj16QxR/HOrGPVUKeGv2XPIUcIDb98xLbEb
wQnnh15KyPbTbuHcIheZyn5KSV3rDWPfrKmorO9gXaDP1Aajr2/JriU9LSVU8wM9
zTlp9OKeL3RpQ7WuSkLqpBiRqrldmwcGhqstzlQu73B0glkNbPdnCR2dIS0Ys4R/
X26wxsinb8SaeHdh7g9OfahBJgNzPriRg4YTCdLpOTt1v+lBUcU9H0jl7Bv9TuGo
fwOPb/bFFibQkIRnbPjo3gsx24q/aZCXcYHhaAXdjsKb8FPqbOaXv+iJLKh9Ioxh
wC/4VQRKHo2daslHY8bqYpNsEs8BwoRUdsLLPDxXxHMwcv8LHMj5wBvioYOkLs/Q
l9XJ4FHSZzBYfje+IGeKPGvVZfwxZcO4Nyekcuq9R0Fg5sKTjEpG7mJy5GMf85nZ
C4F68kwF6uTMWN799wB/vz1gdkn3uEF4VQRTqrYlH1cFUbYsrGzOeAwAVd1r+07g
v6hrcjQjnqLFjhViPh0kkvl7H+0430WvZ7OEO3YUbmDPtiiL+3qM4KGSEstlC5/q
y6r2VpgN4pN9M/iAlvj3Mw==
`pragma protect end_protected

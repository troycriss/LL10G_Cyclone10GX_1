`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
U1jYDNstJEX2dKwIEnBcshhl9Vkdk0QYYH+K2CfPTg7ch2d41GgBS7SjMI2ZRUSf
tnz9CsEfansl3XMTOTRaC8aMvhrvyPt4O+JcGkR8NJXlgeD6pQz7R5T6HkqYPw4f
6PDG6vQYzCyt4kDMMVYgFmC8trRamSNWXb/C0eRMOu4=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 3072), data_block
6nFX5QvFKl/fctrWHPwJlXPZeNsbRm+Jf+SyTgdkDIr09FdBdnJ9uZH0T0XFI4mh
frHzovc+0JudiIXxSb3tbBWHygXulWLsCY27SfXAMjqvGt8/E28ymdLPy7QwI/z+
AHoQyTVGCZOI5NPIQT+BHh14FLDFTtGd4bu8kEq2Tvl/L8gpXt3NEX8WmAgDhVzj
oc4AYsJ7oGYzTQWYA4zB4hVf1Ud3gmZ8WQCQiiZT+iM/y+dJzuKpzr3xwtHOpsQ2
0lian/zYm3l5AtC8/Tpq8dGCd4whi47K0k7fH7ZY7254rWb2RTxn2HVUa2iknCEj
HV/CPeHnOStZOv2Y4bOkrWzcXXuqZhG7+p2uH4gb2W++fB4NI3eVgXg4IXWealLh
TzUYaOMJO/rGyIaLnaBHysY9kdD5pEqApNRmHGInGChsVzkQJ5jngYBedDCDvNj4
+Uz+9iaVsuWUTqiet49GN1xZg1tJmC35PCcoF7KgkTSF1nP60789pJx9GVdocgOv
vBY5iTxtPXX0x3f3bEHoWYrqsB1HNSrIc9dpVBCQRhEmuEEvltxicK20Q2i9j9GF
RVzosSd6L3zUQCEUCxqocWxlBX54u3aoTPIQUgODSBj4VCwoTDC6H8/eqpFwhVlh
2oZlqOqJRf5xLQ5unEe0d/xGOeuk1tHh6md78r1dW4OpxZr5uvsaAf74049fowRX
05R/5WiyN4dGq7rR9FIeWjRfKxgfZI7WdTFpdFpgu+LdssbpsdA/Aa70Dnv71ZKg
8OB6wg2rGPfvqM+OX+2c8rJkMwTqCKDPjYcT1yzSIBAsVCr/8JG6RCzxALqICmqI
ChYaNWhmTfrNeXZKnzbrN61Rsr6WCIe2/We2g4v3LdMvyyQdc/rHSnl1XL/1rI+k
Tt9Mj0jTjIQH/6/4BoyxNzaVdWGgmRl2Ln0n5GzmfqWU95W4vqVSpB2f7gFG2aI7
9GXB8/taj0jv2ionKDGAai5qlWIQHDjRLosyr2vA9D9dL9O5a5too1RgMbuwRUCm
zM/Z0rtN5xPNH1pXGhKKyenOgGFeIjItQE9xLgeQSLEKkl47B76RwF/udAw9ut3r
CG5P1MLo25GT7hIp8UYq88mVqoX24PIc+OPyj7WHF/A8cNgWccIUIpL92VnGF4LO
D+FaAAl9WX+mXXLXjxFAhoVVc+NA+QR3SgaQC1m7GQp1PWotp6M7yMQ8xZGXndgG
GNTbLYAXeiZvvhLqTJ+ogy9lWuk9QTKNx+j58RwEF0ptae6BJViQR+WnVpuF+hJr
+GdfK/fNLEqiKDDKyLteO8rWwlyjxdZwwQgVLzEN+KeGHKikcwUizSrX4ZRKp69X
SqgC8dl4PIgbKcr0UdpeIAlHeWekSIQt0Eiw2j89xGny3+buIxCMgJvQoG0hNPNg
S2L0qTmVPfusxMv2nlM8rYUHqlVH9fn0cyVz7kydk7gb1dnXGw257rNA2Zu/lHJE
+WN4iCtT6UG0VZjhff+cW6aR8oACQxxcTmsakpBSRPHUPlZQhfJJ2qXkup+njEXc
YJ6abcWPMXEGES1Sst9UYSnFnM9iLq59N5rMCkfdqKO6TRubPxcH1x0C17C6cNcl
lIYgNY4H87gjiLw8VPEmI8yuavdOYICgJw/HTINdDNu4DS2jnFMV4fLqb0hFjTse
nyZNWtdTyGnFcvHjubhMiKKsYY9VlGKGrEyNeJrcdrIWhWbPsZOPZioduzBnlv2V
pSIUXcr5G+qnMIHYTpXx5ieklffm38e5dKpcD6KdED2g0fj8rNQFevHnEGUFgPyH
M2Z8/b5LcmRFOPKChhQgsWpeHPX7W+G/eIhu/M8Qp350lOx8chpaDSQYApuQylBr
EgSri810xD8oiZyMn1UgGkGe2i7+G1GHiWKfrrQ8alo4V7o2+XWfQCBbXbceIDn0
yW2Fg6NIv+BmxBUmY27ZO0XzOe2iLfriJjSoILyMh4N/ollHq88tCGXQSImcGazU
acowQMpP+es70DSbZpVJefQjbNucNdUSBxM0X8X5InFO3UiJ55QyheiyDnsmkgjv
yt2udAOcH0WuHaP4zAJr98SfwOd2uNPU6nfwIN5rajNCYrgdzSQvQYQ7RTCFyZdt
elTR3vswzaIGkUA6gk1tIW0KK/Ey5US797/rFtd3acHjR4oU+/QK+rZw7iPLmsAj
iNLIfb+UubhX7qN4Q4/PWi7qsJB0s6N/54fFWgO+Y/szmzWYpUdsQ8ZDDhtXDxXZ
22UdFQPH5lFTVpdoqi+7pACCQBJ782bN8f7tpboUxfyo5TT8eOEHpF4I96mVda4W
PIJRJXXDbTzE0rNFnDOrzZNsu2BegGg1GnLd4IR74FvfloaPo9cbhZZKRvFDxOk2
Kn/GI7ggAkSPJo0vFpeENExCeqNYCh0fosbTpEVRw+9Cq66q+LGXi2eJRgT9Ufp2
ymXIJWcYAwHjpcE3ewZe8oNqy5Juoo/v0mCCdxhHWH6Krp+fDHiez4UebZqZp0Xw
e86sbdF2xdUfkKhRWMdULxUK5ObhOKHei4t61MUznPyJ63aD59yS7PfKatojkZjr
snXe3rEGrpcBG7TNoxVoZLg803H6v1GCzxH8MhRFenIcoVzlEokBTxenYqYZ6ATW
nT2siuWsDQLMtWD3MNkx84jrDYtaleR1yyD5vMtjQl51S5QzYc6SLPVFiQZpuPTM
1wOfiLcFsQhXf3mwJRoRF6tXtpr6+XNqjFFqmh9JDFNFQe/ieBvYMhIe1k8kCsOt
US4qB9gtUNbaj6amX+3Zwb/qvX870a/knlzm4Rt7neRnBBzFVCwexzCnx7MOYe4n
R5dXbyfMargi1dP2/f+xAtURnBVd/g60Jbes54mEnzESzVeJr8cP3cJuRDXBU816
2eSOoCcQ7xMtdG+5rZAPaT7yunIVtBMyoQpcVmZzD9HeF3JyqEIi+cjQtamsM+HN
ep4zy5Byf0SYffrxJQMKQpMmpE7giGQ9zjGGku/pW8dy9a5dU5i3sglfGROAF48D
jOY09lRDpsd/OWn6er+DvFCPZ52/eF/bafbYfkstbdnVTp2q0ap2d2tesPP7/Po+
Vd44jLSlPS73+q74d/Sof4vyHJ4K5Rf6e2kK7wGZdG+DVGpc59WST6qmXsgMccg6
sT0pmcPUj5+JHejc+gu3L4vRVMT6l+iCSqnf4kKsPlwrhZ0eWsfzD2smi4a2rptg
OQ0IJqqTwWznIwiUvQregD+FnknSNAxEDWhU7HHyFdJlykHIqoY5SRzwAtVn2OQp
p+vkM+yjdG09ZH9NcV5qiXga3dOHpiIQ1LB8kLECmzL844JY6u1uDasyXTcefBWX
A/45IQhpjF5aJG+dIlfyQdP7GRYWgYH6cUirjQ26wFZLLeUuKiGFI9VqkPmOWL8K
hBPkgE0nUl+6Hc9hhIdtTKqfyxmHgbDQQJYgi0bYF0laI+87Nyhwwmj74mihuVl4
oiLOJXOBxMBn/QJCLKIF1KysbkGhk0fYE/oKYEwy46PPrjQgrSJN9bVPkbjrlD0t
LZllIiJ5DhVe0U4cA+CUI+dBdbQlLUDCF1ilde8yhuLnCa/1JNF+iX4GgtotvQBb
JBQXDjeHEqx1l+sA5osqECvW7/zI7D5qZUYF+w48PHV2e8P8R+CfkR2wBhHRydy3
fLNfSBGt2HxnhGoXT6WD3PYMf/rxPFR2yBrrTKpZHiSY/hr/P/UaRnZe0e9vbzDq
GuMHHmVmEP0nC3RatZKFrL6YpEwfjAh/5i/6FoXZDlcBnArTnjUYo+hIWBe40XR0
QEJ7tCOT6rW6Meh6W7ZYcqY713EPWJvrFXxRq9FuT+lYaWleqfMTrdoBSdamq6K+
zrs1cRSRaVi0BPbCWTpI7p/R+IVmbcDnMg51Afq3eaWirbsLhsxnkquaiT7rPDBQ
o+o5Vo/Yl0X8KaC7Xl+75gT6Bj//4SACmCTiTLX1KFW2wS2u/mbnW5npAu5+0g8I
HWlOY2OpaW/yXXJ2OwQ0dXY28u+bDJJ5A13EeO7aBSmCp8urDtgqUSaoLEMwImed
8+nyjFwP+foVS9C+Ikbz010xu6NvcD0+V7amLTjpaOt66ayY6d4L6twFhZYbZNer
`pragma protect end_protected
